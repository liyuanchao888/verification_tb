
`ifndef GUARD_SVT_AXI_CHECKER_SV
`define GUARD_SVT_AXI_CHECKER_SV

/**
 * Class declaration of each of the error check stats instances using the 
 * `SVT_ERR_CHECK_STATS_COV_EXTENDED_CLASS_DECL(stats_name) MACRO.
 * 
 * Each call of the MACRO would declare an extended "svt_err_check_stats_cov.sv" class
 * named as "svt_err_check_stats_cov_<stats_name>".
 */
`ifndef SVT_VMM_TECHNOLOGY

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
E1PUUKDTbsy/5XsQebe4xBecP0vyAs8qab1iCitqmm3ixc5+TbXBsLn0vCVI+b4m
AlEaazI7s5xKxIcsDpXUb0q/rzvtMo6IV6V+nzFEyMpfCbHA76pxzBXf8gxUOBi3
O2qOR1iPZJOmWSYXyz23Yx2Fi0X+xMcFckntiEfJrXJXA9udAOYGoQ==
//pragma protect end_key_block
//pragma protect digest_block
DAvfhUWNveKIgbO2sxeANpFpHmU=
//pragma protect end_digest_block
//pragma protect data_block
xq78efh34MvLRbuPoNDFpHruXbCzZpoZul5fRPFH8mfIFbyqbn83jokWWQnhuYdE
XKJjy2mJnu68wVDi+9FJQkhdCl8IqN4U5lgjv0AKMhllBeQvWm31um85lE/leqRt
ClPlxuNkU5vn4t0sjsdwg1YPhAEZM53Owj3lc1oifHkOAc7UhtdyMTVuFcCZPG4X
4wNi7oEpsRfGsPyXDA7eJ6zTkcRVSy4wDPDVBoAOVo8Kw1ZN36rhPgp1yzjWvSKz
JLlbl/EQFxurx+busfzNz9aGSM0BdB62rWkFr4Bu7q9tyHmpR5sY6qXZ4HKHbWgN
071K/u//VZPw12rOEGwAAKV0H3nU5FH4fvAbg4WJwZxZy5lQGoY+g0fktElTGU1D
sgux+a4rX+4XcnyzIlqiM7Q81Q8VCOsV9n9JYu5kMXrMM5P0KAxED18jGxXrHkXm
eQZffm0Z+L7oyIsuZLBwI9SCe23ZcBdH7TQbfc8YHxekSh/QdT6D62DFrhOsU9D3
STMoTHQ1PuUAinXYC3RKqEDn205nbde9K/hId9rmORjLKHHJK0tPucJwc8djOlHU
hd8SSlsoMA3j5jOuhR6mDx7OpcE5FgHWs7DtJFd9nBhh1o1ch1beARcWEJ/KiU4e
xiaO+IpxT+v5SIPzm2hnHW632hGOSLiYgTBTywKHH+uutSuuFIH8txTlPVEMCl2I
nMyUZuB8RKjpWd6PkFicNPNpP64uYAISax7pcFEpXBRerchGSt6k6RAp4zZBZ5Rn
VGEDzPbCqiru6Bh0hRmFNtcv+QdjlwQZ+LHdU6Iu3UHnI3nuQs3dp41JS0OPmwi0
HUFEEHllLRCQ7wwAoSA23h0jbV572ArtF8d8AFIK+4sIMVNv53XpT/BmxmTWyr7A
SO/ShWdKcmZTYVfBesx9WLx6fDcswfr8yFoLbIPwdwlnN4kn6t5ZdsUU9IrRnkBq
vQpx5MdDUFnb3tfQslvhV5KF+KHsTdkVQb3gVhEQbHvbxeeAy20eiy7C97gMDMtV
Up5Eg8RSBKTCUst0dwIjP/zoIx+Hy9+H1Mzp6tlZizLT8u8G9jTevZNsa/1QzHtt
FbWz8MXAPTpFAI7egdVja1C9sZuXrgllY05AvncB8zBKid6QOR39UajyMRw4zOEf
s11/p4t0xnmxvewJMVrP9uWXC/yLh+RqXloiuBwxeceGNUoof+FVn3xknV32iI9/
53yDl3IIb2M3Cq5jia5Ugn7OFqcOXRy7Iak5i4Rq/Dm70wzK9Qt2oOWrp+ifK//p
qwIp9GHKDK7q1m/WSKG1HF8ituGeWgGnpIJ7YjmJcFxJl53R3UvpE21Ta1OfTxPx
qzzCjLb7OzXs76PfVFQV61LvIxKxCL31TAssvJ4p98oGAAKGS+3SnuTU4m1i5Coz
08WHTlAJOiu7SacR53SGiaWZ+asLgtvaYupCLhVnJNGAapwwnHXhGtkEZoqP6AtJ
//VF8x+1ih6aEt5xVavRwkJ25INsGvuAL0PTWZB7LkLgJt/eWIo3+dLafKGWKZNe
X1iTbk+ml2oYP3t8aFf5I/gNVveIKmv06ZKDxwUlXZJBBc2V2C8XFOaMvTHLCkMQ
50JZ7mMaeuTGZKARU/q1Gw9Y3SosZQr+uL0AiAAfWwjlS3odb1LAEEBffBXU2nRQ
L9GYMNI680hDfm9Wp0MzjwTAgHQSGJhrW+7c5sNLLCBdRbAwOmtViZlbMqRu3t0r
9l30ittkvuNw99/hiQxBpiEhcgYaIXKGWnDtezBCHsQY2YQYgd2jiICqT/lsCU7k
7BY13cUQhIZdkQWIG2avpaOi22y7y+Rgd3cHTxOHBPjnFccS3qsNuuxIdpbTLV4S
IP03n4hsm4onO2aw5bBZLqIpYIQUST5zAF6+h59LDWATzdTkDDE1M9pcPJe0m4vC
ixI3AnO5tdVKpXpap2Q77x3d2b+n8HqP24iG3r/1th5/MUcFINwbmRg37G2/GkYg
naedTztx5GTklfDSCwKCbHzaJtHOpgtvX3y6NGaOxUC1KCOtPtzOvmKRk17RqcRn
tI+h1c05o7CFqKKm/1yhmYBHiXE2EuzT1NQKTpNI2XyY07tPi4B6nmZHkbWIkoOi
xtfvpi/ubdzEyc4jv+K/z92LtJaKbxui3CRYxWGUeHXT4pZK3CE89Ldz5k1ib4oF
tqP/5RSL98yAs2wVEuIGcQFxv4aohIOLbA6XtWna+E5lqWRkcO4dj1uNQJO9eCBp
v1SuHqdv22PkP8TpZZ7mxCA9KjYtWRgVlejIgIxp+6qp8AKrd/v4vGjfWBZGdMOd
EWtFv938gqWoNgfPfe6RAqDRjMqKhU4Tx7V96/dWCWGMdxARZh7RVkraiVeBYf/a
PeX904YqoeqhotOOFFu77kqYmxcQdMDw/Vu52qK3LaIuXMQU1WlHewsfSCtKVVhf
tC/KYcm21wIfFOutkycu01HEC3Jn3f4Iczgkc2YK9IyEYN64M1xtoikzBdVDByMi
6WVJKNquehsUtfL9ffTvygecDDIRP521dPFhANbue1ljGL3C/VAeSlbN4XlR7ctG
LaAWyrg4r0YHZlbS7L1etoV5RqwwxBIi4b85lLnuwhwiwKWRDxgZ4p0djrRK8OCx
8WN0jXOHtXmOH7KUgozFCmIZtBny4JyqvrVex8itngkj1MYqzeSXLJ3+HhtKFprp
bSVfvBvK6ZbUE56ODslvbHpkagzxOyI3z78OtwMdo818tav4QjYwWEzoxUkOJbJi
8R0/nTSkxIelwxG1roW7bHUrbL+pzP6aNrOtqhimUuPJFYTSqQi2eqr3dES6LEna
uTXHkJAtV+gudl8m/aACqIMVHuoT+/D37JS8v7uM1J2WjL9qk/P0MwL1ROCiFHL6
am8TkuliSf/17MXkpj1paJHR5zfA0F/UsgNv1+Zbgp2HR9JXlhq3B17OEl4kCwaU
Zd1kIWWO5Y4Sc44ySIDRzKg12SO5VcKDBOu4OCBHdRuT19pwVhZkVnRUcWkeAynv
8JrrUYcSFTpux28gtIJl/M1NCklDg0XU+LKE+ioiCXp7DHsnsojsAT+uiNW6z6ZY
3iKzMMNw+N4NJeTNtl6O2GEKkXKncjJqsz+bhYcojSLLMRV/ztKteOvUpzZ4WZy4
kH6JoXP63yZhEYlvnU57TsRV6EC8mptPh/2X9BIfO/Fh4A4JHZ1EeAhEBBBIDE1D
uUmda7tqz8FKkcWlKzs7uYKendWbffzkH7roGB9xSWYQgw8x9wpA5vaSVnAkjqP5
b8rrPfwXjW56sUgH7CDF9Hc6cSvvJUOBBk6mvmiUNgmrMjZegf3ZEOjREi0GphLp
oRiPeMt9hWAA9BzEBNSNKjcAh/Cdj9f1nVupfC+Qg4cURh4igu9Khh3lca2OGxDX
hgqcPBkS3MoDOAF2Iu6jpYAcJn2MZJhW8kwSZK0op4XxXbzZskQD2oP2UDPta41r
eUy9tT0D6ZlQH7E/NF+jy9y5Whm1/bBUzDhlKC2LYGc5Sv5wEvfMoSaynQYAq+pL
M6noXCQchfd8XuXDFNsYhKy1G9VLT2Mxb1yFHqKakeaJrxgxpJVyyL9n+vA9dGjF
OAYrUYY0kOK8qPKRwbG0WLIKnyFnf8EpdcTy2LExs0HX6D7h6U/j2WFsHf2YqNXr
UK98/2RURcKqEpXhSGSYnqM84d1j0DHQ7lFRYU6G4bFOEJQi1NOGS4LI1oTS67wN
6dujq8pauwTP0cayNzvBibnwbadKaKCSRRteNvNvP/EEZsBiej0xKCYXyGDx52EG
4Yt99j3jukrer1wN/m8oNxz9v9Qa4o0kitsEDOGgH6/7iwlsdBPcf7uVcOrndEPz
wkNTgP3JTNXJUaSQIr8IO/qrJyU2FD4c+AN5KILtD2EE97864Rb/f/MXFjUVXT9Q
EcBh7znkbeoSUtgM0MPNucwHRWVlP/hy/9h7FoIaue3Qx5bA2AaLeTYMs6hDiz1E
fEkR+7QWZhO2DVRlcmVXZUCOLi8KUhph4aBL2tzYhFrlZszoKN3sY7MEvYMiI407
lYPvop+Up6SbXnjDDSCLTtZofBH2WIXe0aJ3TlrXniElLqYj7GUJwGoMAMHOdwiV
Du4viJT7PjfhtvTm++OJk6wJWeYxb+Wv+ww63aht948gXBxnok0zTYBMX72ow1oA
0Eo3A5H43550Iba1t9Wh8OcLkXynQMdquJiZjR/D/Atm+0eR7F9j5kwijnJDwo/Y
SjY/u5vljAIGQn83HFIauu9qJWWCQ6enWIAZ5Pv6hWcpQu24qqoBc2O6KqjbB9r5
QcJGBT4G8R0y9ox4MQne7ahLE92LMHb3WvWi20mlXRsSVj1GdSRYcKOlhF/Rs7Nj
c+JIQ+5A6t3UJCWpl8Af00B8UASyVMtDelC2vRCJDtOqRV4by0lxC84R9w6b7Rpd
cSud24jqWq1kxPpnzOEj9osrxVfQFZvnkmz3+G37ITzQwH0qMr1FKv2A2gUadst0
nMlYf36pia1RF1BKyIYTFbwmfjepJiD9YorNKDXzZO+46r4FvUIZuL3goXzSV5EN
dtdwyTBmq9SatJTm1qNaZIyy9BirCzDzc06V8rHPpAP5wowNnzcSchZfeLESTKyQ
c+MAVR/ofZTJ/fqE/oS6D+aXoyA886yYhmP2GEYOiozYasK3k5fgaJwJhfk7P9yY
N9iIhmcg2Dm4arVNWHKi5HsKEDgIChyd3HsmvldzmZIKWeto6vYWvdAtGPY3AOGU
tVvqsIcmzhlRaecaPnOKdqcjB/8hEUgbSd/+OvewTcd2eSXctnB2I9qT6mNTVP+S
6TUgiiE+87UGobPcrqOS4xAkuh3FhSuqWdNrC3qVR+IwfCh6+8RcgJl5wyTvoYkl
EFncJH7ByNxknh23uMnYin8LKqH6nwi4XewLLFCaj0itog0dkdmtKdUhIL3wqaHG
/z8/lFrlhPwByzLStlNwuvlG5b9+MfLTWXrlAu8EUcGtHPsFV6xGXEQyVCWbl5nG
rbs6e2DlpL/boJtdL6nZOotaJorwN+3/yMCCV9EwN3Ft+OvjUqAOPZCjbAMo+IQr
Wms9vNJFeNUZ9iW+ZXRIrjbfnGHI2I7EwWWU7M+7VEfuPZESCcjAlL5ckgVZVxML
6qZOLsTBv8NiH9ak02SDGjb2oUNkDCaCFsedSuz3JU2ja98WfTXOAMbtjk78WZWC
laklGMFRut08tGbD1alBsrZA9WgEMHMJ/qVj+O8yi5jVb90I7wNKjqv03201iKst
eTzE3gYidWZH28/iqss5BRa73yv1R7LA2CWFhWfWTVZQ/5JNVtDGW7LhGW5vnbcC
fzjHuaC+aQK5sGC0d2IEvTy4ETejGNiFKLhFxU+xx3aeFfG0MsXfZQYSTCVFX71h
+wtYnquJh7azPLmHnbMRRjgYBiLjAaDXsZqhexbV6sJ5YcEFd8E0FMs0qyE33Ubg
CfbqPI+eBR+a1PdwojFrJpAEVvVqg3M5udCj+ZYic/rpqy6PfLHnnvCCzVQXrL8z
W0V7I6ToEg8ubGxBmtwOM/iTNhbmCLdjUZR/1mjT4vBvYQpWl4GyLrvhNWkTX21w
565rS5nEFghYYZHM0819WL3RqHOlE3sr9xa5dEg1oZqLub4ywJvXqIerWyTjNz2G
INhen3XWhaM5mLh++vQLariJWMCH6kSqSb1KZ5SL4B3V9gwBbgXQlWYgQ5ZPH9oI
pglqW7vD0F8ziKMONQvPX3mmhOqrvQGrZA/uzX0tHiO0MrMIgj5pnMgLxaTSEN4r
tgnP3mfDdNH+6DkLL4YgJwWH7EsGnUpVf8Rr+Li51izD+0YgmA19ZMFtlGguV6TA
QO5wXBrsr7Q/Zb/QQ//yzWMK8e0oqRDDRrUsVCRrz5Z3AHO1YYxnuqRpRFcr7IRL
Lh83AF4a8MlnPCNyoQH/H0HXRVXH++vITKSvpP0RwhBICHrK54AMiBFKCZ1bwNnH
AH+CgS4c3uE/iFst1ODUL9Dtnb6d8mTUYJNSRypdR9aJOm7VSThB2B8rIdxpgVKW
JS9KEzIVxfnYEBzYFI8QTCl5oMc096Jf9lOCM/doO6cp8d+THfbvpp9r82l5ADki
Bdl5nouSDXWsZQBSyD3ZnIN4R/mCiuXV7xgTkLuW8TkkF9mpfSOUeGxLvJQpR6dm
1DTDznzL+XLFrLKHOonabYe5bJkuOK/6A+oXKABbHp4ZoFkcHV04xTu69oBy4bWb
lhUi/8/OLswazl3Ntg27yLRtskRIkxjOmGn+oXCyMy7glkpcmLUPOkwSzv9Ur+sj
9/e8WyxpxzE2TUNdsl6QxyS/cGy4MTVO9fDdJSQQpYEIt0b72nAUA0I1MABiiNIj
geleNi+IBd/7ez8WwGlrD9QNzr2uAzEm87Kxk+nCze4H5V0lryfD6zfW1f7khv6P
EzLNW1h1dHMIQ0VOzHhaHyyzCyMwmVQMEngaotPTwIOzMm/dU+xNt58t/3e40Eio
kB1jAzNDp0JyfmNG9b3e07hDI9HF1/HFjD4b5b2YlPZcdDcpchdkwTUHgJqsSbJs
QfMwYUuM2dHHthiiR+puhhSETtlHyO/46Lo3OXfnULGBz4CdSy728S7LNNi6Of/L
lrIroIsIKkXqNLbPGeNqMre3ZNokmCMc1atTZ6xXWiyoM+TIZYUYm7QMymrpJ2Ey
+uXBOy2lvI2cKxaaXrJtV4c6E7s60WTY4nKz+GmE9CelxcVdAr5QXFpAJMnGPRgv
gZEjo9hhNAdw6BrFXFQDyBVJr1dBxGLikcyCBkDzombAEA6VAyrD5w9U2q+1BNfi
NB6jAS0rTDaplI2vOS1mCK4hXk1VNw10vgYl8+CDmkRfvCURjLQ34B51nxAjRLmh
lkLcEksbRCCI4/4BBo9ELyOZODNkyDVp6+ob8JMKxZodogcvcM67fqbxt5fra1mt
m9LG2Ak92FWR7LGvmAVFKkQyigKiw2tKFrtNrmxFR8uTwY86yTLPdPxv+WJU/P1V
UIqxRV/MJzNg5qigJyh7rkOFMkzzAunjfe/V9g+Qmoxs7J4K3R2xsCr68k2HevHY
FJAKOVHOmq+kZVoy83Co3ZR1BWQ9WPyWCfDQ2mdOLT+cbBOHgnZm1vJkldrQU/BP
dAWrFpp1EtmnYARkUUk3cct5SEZekDEsl6ksYeFNUXJpg+rZu7DxaMnvUk12jTme
ff6YiLAX6Pvwzl6OrzIZ9a9wqI/MUIRPNoY3rxpSU7AKrMOBoxvNBhXTBqx0utLp
n3H8srBi0pMF7Fd69j5AFtZoB7S2ZWCdHBHOw0NLfRdX1StcfvqksHIXoq01jitz
wZoonu+E4RBW4XaHtP7C/aLrl8HiHfbCM5YZUI40iv8KtMgOLLdRuyT8TabdAJ0k
HlKaMDRZroo4n4QqhRVp+PafPQvzirXyxrrBkwBf+ODY0lYdVeKkYbC1YBnwbNHJ
IQdPoEYBa3mdfpf0rrUlSPKRaB4HlqueJycj9dYDYXO7WenfCROGoSYOHGjOVvGr
ZaHlOBrm+kyatVR+w91zyujhLqs+hMsMfykQNw667QuvmfXFwBD8YQ8IrRQpYZq+
qjVXwlh/O6P8z8eaEza4RCQbRdCc/En15VqJmVf2mrZ1X0fNexVU9kXAMc6Rc2D8
QzmQ+bANDZoU1bHaPiQvktkn7z4cXqxu7pdvytsX3vP0+k3Bxz/V98zuYEubDG38
X1mncKlkz+96RZFbA94AaPQzGQWnKrWZmovJQ/7spyDIEbRdsxpZcNR3TagQUJlO
TJ0oWXfGgIeQFPn6BBciIG6c745HB21HIJmtu8BZiryQAiYikKP9GWnF3Uju5G/2
PY8bG+xPVwfhveDuFUOc4U4mXbdRhHtcwvm0y0wnR4pO/1uiG5kuJ1PIz+5npp9Z
3TyeYw4pR6WCkal3sp+Qx7dGvfLBvubuPtGoFTv51rYvECUO76TuFI1kAE4O2Zye
OgAyaJTYZeYVNYkB5KB36fWIXjrpFksppjRpWnVl39keEEtF/QOVRBG42np7UODt
rB/nUeSiUB+Gdefaxk9+zn2ATqCQpVpoGxZ2U81u6tuqDUDU2u5a50fogAAy9hrA
OJoggOrBJ248BJ5eRplqhhOsXdIdejAFK4h2rCbtY/qHSCBAn9pq1ayrVH2EDtGl
7iUru+RaFSvri8GR0/74d25RrFv0EBqF7EFQd23IHuiXnz3fSkXSw+0IaS2cOmGx
dlRuUwzzNIMSXcmHobL1Hl9JmmhVN2Q27kcVqBDM0Ybq7Z8iYgbmdXj8Rcjh/DNZ
0tHr7NXJeMyn7AjWXi/tA72gKftNtBnTPpBuD3KyhaZn/bpZ+FkggpFS+3ig3hsC
cfCEIQgbKHTerqxZcr+j5RgcRcrZsyXdErAV9HJFZ7WBStvrc4hA6W3KbEInEYrl
uW7svikuLyxToKoSRoO1xsGxguMza8elBVjbWo0drK6a6uIOZbW4wipAXXZa42Zd
lAUPC2KK/VMe9of8NXoJKEpHqwwRipvkeogNsNtjwu95Dg9kLLAF/G6krZN6jd0/
Oj4v7XTdGZcoU1ns18kRMigll7XhaIC/eQEGXHaZoFN2/LuPbaYIqaZ0GLRATIj3
gSdRGEmoU8fqR6kEs3OQaY2l3I76lC/0Pg7wcJkwceHLhehaVKZNAt50rLUOpJ4e
/A1w4iBbCpcr3RzDTyZIQySI5RNlaRGIU3K3L0AATIAX0/NHCRc4tFkokkm/h31f
d9iMiicFr14T5obqceXdxR3QpPia8+w6uqF3rolV0TU7fPqRIA0PGGcBbjrksCD5
7W320F3lUyqBJpFZcX7opCvW/QTWDYZxlcmtkDzkzgw53k0QrOZTggqGkc/T9Pr1
4SVJKBjspxTC7YFh1rSmEA8kLCRXDHc+K5XEjZ53sbhjA9F7GL3fAOdFfL7F54Jz
7J5LOPsbBvSM3L19Oqa1bz+fZlDDEvH071N994G23Tv+wuoh3tb/RztpptZjgXRl
nI6ngZ1gcLspTzEltVpD8mzO96AFaz1i/W+d16Tze9IBRtoN7MeS6lCOAuZaBlbM
cICJxnEOfueprEPbVkUqMLxZmH6peUOHma96yZuhl+ijL3NN++MjIG9SLj+MarNA
ntlreF8yZT+ZimgyrU5QbTp8BrKvQ0VXQdhuh/AQXx/nBk4+bvjEdV/QXOzVJmOo
aUfdLIEq2J9TcqZcUUm162ikMNgJxjeZ8JO0DPF6dlfcoqaG+pluJKTHHVEOrvB4
32vsImBJEJkkzpL5NKvmzG8qOmu0JnUC5PVxFyy6l6GAAYUVIq8v091c8T7UFVNQ
YT8KwafFZPHkYSeS9ARsssB7DN1MO9gczaoLmm/FtG3BLfDRRfk10TpxfB7ebl0d
tx3TIwUjMUYfQ3CDDHZW66k+j4xENU+a0URCOpsfcFzu0rg5V8aMs6kxc85mt/Jc
0RHlqsrby3t0dG+AVKLNkr+DwLkMtILLXeZvCZaA9ucZX8DKXeOQ78ofLj3qfAAC
s4qqaycAuUlCPU0c4FLbY28+iWQTRc3Dofd+72vagTEsSDnojaam98DCV/1OV64Q
/nWMHBnriw3RMtvvAofhYV5oLFSNSYG4x2GIInO9nitUaINLXtrieg2Zrs5lTbyf
vKgX43+YpiZZh9mINvp124UAdZtN6Li6pmxTEJwEDSMzeDfDINGcUuWdzNFGIu2j
F1G/LcgSGwbf258iMejFzizKiIpFyEP0d5LwkqcBR1vgl9loV0BPB/JdEkbY1Bcf
JtlSqxMwBF1AT7oYcPbNw79Y0yWAaTgxCZHJPplKE86xBTSHwCpxlgJYCwdSKNHq
BIjTUrBf5VOa3U27Jzu2CC8iG75ih0xJtJy1WBAFqgU5i6HfTK+8fZJpqCZkL5s7
2jjKJKzszWSsd/RU6HnacM7eAeKq8BRjQfOqaLbqykANOb0ffmLSkoaYICQAq5xK
rGjpCfZVMcHHHGGallTcK2EBrjzoluD3wYv0XgtqP9+ZcgDbX0bACuuuDmKwSnwS
wRivpJXy+NYMKhVjsgf4AujZkoqY8sC17Aij7YGFWDG5Q+ChBzs4okSd63dQui3Z
F46R8RJBPr+92jYbwH+WC7Bg1ON/PoqZx2yc1uxjEZ27SIxeBbmD63Be1uVyoG09
b4tTaXq6+Xlfj2t/Xj/0oEH/L4cIo8RySZp2Gz+XtoEqyUSRvO0eEY15N6BY65/B
Yj9d02alqRlBYrrXlJQFSFz8QMo9bcgV5JvR4NoCpRm4/y8Rm/GTwRUIsbMe9Udn
bYfCIu7N8UDA2+7US0iy7/S96k+3kV6BqoaJEmOH6aqDwTwK20aPN9hJZi09PfEO
o1Y1Sr2xJjslrzB/G+qZvlcULaPXFtdFzEW41WP7Jd7kCaEyN98Zh+2+2lOQwTxS
ohwtX494odE9EiNFsdGxxInMaYk50KpTYKCQpwMwgfWQojlcOgNy2bwE0RgWkj7m
wAjU6QGLYFtCV/xCBxrF8BtEpzc+DrtsRKGVF6dQNyJBYEQFVZwejfiGHYKOlOMg
87i3BoveYfvt3G3bkhN/MlOofgoF3g2dQXjqWzcEuXH9MKxKa5alwPlWJMdv9sqv
orGu+5EZaZ9nOYmWIK4K+Afs0GiQwzOm/ENvMusG5cL1mtT/2ZNtQDo3w2G7Xv1y
jGlLrFAMLvm/jzDuKxU97Y5FhXY81FGcYrHvjdY8YIu8UVHPpg0FD44e48SvtyYe
EwFs9TSLU3/QYm1XastJuKzUSEGxOyu3za07VSuaUbgspvjSWRouZcR1qW7nstl5
0msO2kS3+3A8/+FsV+W3aoyHTCI5rZaLdl9QuDF/PaY/VBa3OliqV19tRhRtGs3Y
t74Yvnkja9DX97qLqj/rBN796h7A6O9NOOWDAyjKNDwChPwHFue60Oc1MXFlQ2Rf
FqKJBB2U8CuaVjR1sKv1GC+8jiD9/fWoMXzNGtG5/zSm+GL9tKOPnLe9an/yKFbb
I77uEHe2SzVu4FUU6Yhdv5JFFcV1OveHX6lct10kytHxqFf2/n2pKyL5138GZydj
95qz20x61gUWXb+MSN3ueBijPydwMovJntM4zxPdxHasW5t5laZShwfis+TJCSLa
sv7vmdvMIXaWsC/FIFXrHgjFXqjB08i06+1YbXx79ghIfjfum4SOBo/79hhWXiho
kqSSjQcsXLhknGJaH0YZRggpVLJrFSMys4R6vePky3tjRUy3VGKxGtVZiXwvoBKh
soh9xTKFBgxHZr+wDDhyVWbolh6D+Bf++SNX5RhA1TIZ26iwHPBLU2cLCyn8gV0j
/59oOBg7zhV5bPZ5aByxSXhgWJWXNo0GlZKjtAPjh4UfG+EECccKDh2pif8sWMkg
oEAKnRAx2ybsDkEr9FwokPdLZN+9NDGUVPLZUmlmu88H1Ldn0idXj/wD8AuWG45q
etQo+EoOJ4V5rVQtXioxuQsDfh8ZInS6glZjU8BLldSIOqnB1cOLrYVLfrIMvlxB
ph9PtqFh07ChvHLVS98wGzJ9HURLafVXBlUzbHhSKfZ6NDeZ5+3WySoqk3/CxdnD
G0DrbqBjg7m+r4XaOUzxblJ+k3bZaPJuoR8K7IBEYQUCF8Rkpnw1239DBzsG+e4F
flUu6ZESTvnKPs+vbHt53CjV0hGX6ELRw9mjWJkOMwzQt8U+vYXcdV8R8gryvnsx
N3PLV0pKyrOGeNT5XTHuO1OVHrsBQZgrGFauUDkJYoZ+GXjFBkQZ7Wk7FJG5TS6k
SZWud+cep1swxxCyMPD6JHayttmn4j5OQXaCKHGYq++pgrOVAJ/edCPEnLiFwEnf
Pl1ObqTVD7xyg48qSSL3zlNHikq3FCHSHgyFRWG6nagZPj35i8FGABcGsTEaYwt3
S6dZGHT2piXSmrCmCYkWaTyODd2AIyJIWGIP8zUddINsLL+r9lv0ur/UDz4pKG1T
k8w6Elu5rN4DVdhi1+G+jqRmmgsmjx7mk7eW4k6eo8JPMm46RY0vOaos61s4DGe1
po0a3lhLLx+5RSKzXLGnVhNW0i/fvjIelI1D9wJWo3YF634tTpezQu11LbDpJsYA
Q9aZ0rHQyS6CUc1LkH2x/XkVmrAD/poSasWhIIZ1m3S1KIPwHj5t7LQZWLtVpljP
aBAI34mLeMixZmNBVvPN+SIvFB5ZEXmJTLBIh0o5JD0YCpW3XjKs/HXMZf5Ol/dn
ES/fy/kZtydUi3Ca9a24HFencxWoE8QbDdJ1KCBYRN+nvT0uRa5JoZb4dj+aQxlt
5UVmtqdu7k/W8iIC3ArPAjE14AqEbW+rUsx0JU+ttIWvbnZh2F7scxFM6txT/tH0
0g/N+kVBAXVGdDvaepTDzBU1Nh+B7rzkiiLAocz6Dj1ssrwqpQ8Y+4eIK4Ivz+7D
OpPVcMF07XcFHyWjWf/daIvJm8MSMV5qEFSh+8SElS57UrVms4Ib8rosqqHMeHPo
wcuzV+84DrvF/u6UqdQaGZMQ1OHon0Dq/Oi+LZ6moQDZqIOcIQVUaupsynL+FbNo
RIqMcCq358WRqgctTLMVqMB3rvu2eqJCct3+ezKJdEr0tcyOavjEd1/z9d0e9KDd
Fc7jgekAZX7ZDH5gNuXt3Hqmf3OROzUezcDpOklEt8bZUUysdfe2VgKNO39CNvwz
Z5YYEHvCph97NlRAZzXtBAXN+UdrhfWikTB36GSSQPaJzIJIFnpd8Efe7j7va5d1
JtJ+yclY0e9vah32BmEFR10rQhzxzRN/Ug+1fPb4cy6s7sy51qJ4b9b+W6nurO77
u7rB3YyRAEiuGvhRj2zTbFzt8SHQ9vgYm/u+jivYaNeK4En/ycZGjstA/R+UsVe7
d5PIxYho4ipIQy851TPGDzpLX/eyOmKJMcbEop4h8N8a3XhA4bbYIG0Pq7MukPS5
pZnwxj4NQ34u4p6ViBfuktrtCvNGeiEDfz2dCgZcZLkihW8cv5iz5sF3683eZRvJ
Fj20o2YzGaH0c8VxVX5C/X80D+DL/9uLfM3rSXaHS4wclWyZhCmr9epsy15rKbk0
KITsWNGie4myF9JSGtrnAT2Q+BxC/Qc5LrZdvIZC/cYLWke9gzEn32RrtXwlKrhe
LwDHs+zBPctAX9BoPh0AWlbR3IQ9/sohgPJh46TfEZ+kE9qPHpsNl2JNDU3rWtzt
9nr0yq7aHyE1bsmURFKJiOOKO487TaKiJeSt22m3iWwEq1R+pFGzMedS+61i1Jyl
LvMGrIjNZ/EOksJojlKFRnAJeTzAbIlPN1nX0ZDrtQKPjm9FVkL63prS4ZMSaojt
QGTHZNn5cGFjGnEgUf6I79OhKy1QWGQP9WFvjHsqCesYMRmNKlLJqTKHZWGKhBcA
0+PGHwnbWuo6tkw+YgYnWj1LXrWVYRTat4CbKXcfjiDcDRhVHFbKE40i4spQ7qlw
D7CtQqjNZ02PES4rXVxEkEFiVNr9DwZucpjXNk1NNfmOQpy46R68SezoxZZ7DiAz
fm95iDbbINJ4mz6gXm1qaRhFN4mtDd5MpBSv9BGjQjNgu2L6ayjnP+Df8uwx+kt7
80utFJVXnqyCyTPtpTim+weVdPwo5L0XJCGLJEssPR5Bg96V3qqxW9LYPwVNDVsb
7CuKS+o97OTY1+lr6zbTqr0XmZc7j1ijGmnzGi6JgR5Vs1aP+wXx0EHnQEektKq/
N3DHW7ZiWqvH0f44jLldKGX/OkpY9LEEoAek1Sp8oiCZsQMgbEcxc45dfFjzfG7j
oB+L5CV7FVY7aD7XrO0TaPe2+3FHjmqqbszls0pwtAgnnhPU9fovrrpVeRrUlkqw
tsHuQB52T8WFM1yHP5/wU0iOWmA7/V7BJLVQXOPEA3AvyD60ggVtqGMS6ry8bxHY
nXsjxIJIYlF54zSbNrLG4jgL85SmN6vkF7IG4PGH+vP+G82KEnERVXjCYUshnkhG
b+UjAbw83tEq5l95I9BcFBmxLcgwfZSkoI1QJDnZwJGAtokr744kFnpDOg4BygKZ
w+7SfMW+yeTfn1aSxH7f1CrR/fxTEJYbVhyiKvUGrjU5dpyIOaGpmRtxMBPjP9go
u0YNlxSL2pP6BPC4YOCfD0nf/Gjsasyx5c5lqHsddQvAfRDiwGyhBC16wIhXsNyG
hmtQnmlA0MVCkdupOSQnP3suUNzgYq/m+mGjEmotWRvhxDZUut1bIqDRx6wzb330
CEBLRXmaLsHNE62gA/f1spDG2hn6dAgay+QXHTxcijFxVCr9KVNZvnfXj3EL72MH
VX5/dh0WNzJtLEqdsJKtbYaS3hFo2giB4zsCoAhUmUecP5qcj8Mk1wowBsUk2iii
hDnWQEPdKVnsOtV57Qm0Br1OCXFs/pbCC8vxIKfrUYKJM6suyplQGq3FSlz2dP4D
NcRgcr8T5RDTWlLFnrZ1zyDxZryUBE1dt3Zlbjj85KEMiAqqL72NBcru0HBEkikD
n7lmrQl9qq0d9bj+9dbnRUqW1Dw0xzL2RhYnzpptz7el3ZjPLITwKceTBFOLPquW
inC7xJPiVfwe3Ps1iedBaHGL9sZt9eozY0KtHx9ztmpTT4JWsuYSMJavaxmbOSoi
4wxp49i9kafuozAKQqHs0out+4MqgK9Y1KMBx92DDt9D28PhO6o9XBEb68Kr2Pzf
ydC2HEdF8E98AseElpfk57VhF6NuQlm9jjLsuSqBcHr6LVPpl0Tn/U/kFuH4EI+n
mizQIFcacCtDxn1uzHDyAH/Aapxu+PWXfuNj9yIOJCuSNAFPgop8PyIruxPe2Qkp
L1+9BgTdFzZtNE0b1MhRIUIcP85MN1vvBoiyrtXh7DR+4QDehfzxhF/MHh8TK2/L
+LTGnV/MFSQCPXOrVST2shUADDy2+z77fCOK/6zEfb19zPnFpqYbz7u4ctsfWQ6L
UmVaXcC1yFsrCwgDLZlIFHoHiUd7AH8ejRUDnXYB4YWDVPEbwsHkciUHKrGbVrN/
W8ufu2B7pYj0sFsWET+u8xuqcKYdqHmMSY7sExFDfUF7xadl8iMs8t534NHl1EM/
WF2ssikPo+J4UjHNXEeNjlb8mmtxTCghbqcveTAgGd8O9Tmm7SdNZCCvAtURcAoN
g4yPOwmgnsIIxmpbnka8tv89d8q10qbQqK95WK3oe8tL+LOJ8bnXoMqKUG1lm3+d
QaHXj6dgoGahK+n5aheuN4xmV6TF9eOTZF8ZiqqiRDR/OSuootGf1T7XOHtFEWHl
GpdhuBnCxs5YoPPMJbrzA6GcZ6us5N20aFSmBzt3e18DYRGzmuoZEhrqjsxj27Ut
4UNhgKek36Exlawq26JKI4BRePpuleiCXoeHD5pzM4kiaxFqmPU+8AH/dsSDiAGO
ppC8VI2IyOua6kxriK5Na0UZrEwrn9qPRIOrQF5juYOizqAzqd21H1vSFIanwpzV
xgDti00TqPQP1qZHHoH+UxbLdFaL1BGlxGR5dqoVvfRW3JDT/0u2efxC3QBk6xYA
ID7Kk61ygBQIcg6lP0gI1qLcGK0Fep9qmBUnmhVntGtyW/2SN5TDS9Z1jtmAnzRi
MPmrd+iSYSZJCQlSOC7vvQ0Ag4vcZho/gzmn3Kj/26otYRhir6yxeTdyBxP1mV4E
dP+OzrtYDrJy76SgymtOgwVw7A13uN/3poas/gC/2K0bO7RScPx+pz2k57Zt4zpo
Vh8FlGUV0Ryh3SfTWej9PWH14yhzPjdow4wAalRBxUb5k8KiutdHbs4cwKvdN55x
IVteN9bKgZhjq2mcpOMqNce6HdwFKczebz87GtHzmHbB9e82zOC+z5VsIgkorKYI
qFdFhbhDKKKZuKZT4qNTGe4U14A2y47ySmEF7whmtJ77VfyOAMWMs40vNasJg59I
yKiz3T9pMrBzkM8M1OvdQb60rGGGuEkHkY2zktkR6S6gfiYUbHFXCbRSzJHc6ZER
l0VUL6eJ2OVvaAhqvRnf6shmm7uWJo/pff3FJmtWAup52O8/bdVLMIwlbOydz5zF
rfVtbIcD8+7i16pc3K98U5T6SdmgOFaIurL7Udh4DeUIkC/aCZYi8mzsgYsm6kSG
irsILrI3nAxGKWj8HkKuUcx3M2b7qfWGLIzZSqKJ2hdiFxiKkKpml2qt8xmDnSBq
DazghhHhtTma1bhTL0dNvGMMxPdduEkDJHLmqgQx5y4lVS0J0i4RCZnTeKwUf5nE
HOcCSFRBN2Il9RYdglP4J9O0R2ygkyd93MH7ybwWcvROFJcBgI5asVzD8BaAxB3f
7dAVa9PY6iI3+JQmKOBMFbggVPiLBvKCpj7T0LL0MG9waUf93lM/GnVnz8h8kgCY
iNgSA9QqtjT5XMWmn2eMica4PTJZzT1t6kY9MXCHXOAQ+W8OsMqgcnubvbubBq1v
V/620H87KiStaMope9Rtfq19SWAnM4QA9J9zU0nwUMc19o93Nac45eu5Kr0KNtXT
H9LyCnTQB7NIvffEaJb9IuWmxAksyhd3ok9BViZebzl3c2xuGMQeWMQrEtXoU6pt
l/LC56dykffOonCvjpGcd7CZ+K2AgVOHEAx3Ry0skGcrl0h4dKPE9doRvRh4k3td
lzMae2LAE+rA/FcF3OajOULmjg3M/tNcz0dnY5bb8csjoQ0YzFqm2+OP2iBvDVGe
BIhoxVbd4B7BV4R1/jCsji8aRUPezcgKO3dBNkTE1tXxqXsxKYooAvO1NJpXs3+U
6OBs5KHP0k/s0n+6T+IciiH5/Ok8mpKmDFZrivbgjhuI95NbR2NjlNYCGHu+qA87
B/4CvQH9nmwjFAGjEM3dmUCzIiz8AxebgGzntqNDmBDIgFDEk9TSxSMhdPSQgE1L
QvNHe58Orzp2s2zai7RpPSkMM34M+TQOvLwZwsADGLGyqV9K/05XHOzKlsZv0zB1
akkhi60LxZKjI8RgQR50fbcaW+f/T1Smeumw+xtOSXxiYRr4gu5aMyWcbA0KwH8I
Mj7rsN7L/z9cXnlNH2C1rpoWaaTQB4lHEGfDyflPnqzNmhuomWleqhPI7BGNbxXR
qyozm149W/tysauzSHUfXUMZUen7P4hfdxKlEY524WlrHHRq06q4PanxxMWu0s+F
FfrGrjaVRdGtYObcauEx0lJd4KzVBhKcTaalldL75zIPaFqii3Li0ZYfbcQnnRoQ
Y6mbB3IpdBI2+38RyFw9OLQnAGvcQGxDeEeyNfozvaOLzZkbM3ZqSZnx8nOr+kPQ
yoj289RttEkzwBGW3ysQda9adpmVVTH2CLp9Vz5DU5blQl9iIf+3kI4hmGMZ1+TU
ucCw6koo1p1IFbdoqEn29akWoG0WUTQIWzbND5cCEnJadAVA0GOvPzgKRKxN4GgK
XrYeOHyjqwr6QJcdxrK1eNMdzLs98k2xR0dbSmEG+iHDg9Diq4/dj1smXwVUgVO8
isgJvEmBlUNg4tr6Lw270fY7eX9UgJnJUnSINAYeMBjfJBpGnLaNNzpx8sHZegje
2gvRd7qDz7cz+POj3ABYT/41ATvQfCxp6Hx0bl3WGPRf79wPZTbY+JdDBEj9rSaz
LuMkfP96LUuzbl8YzjtxA0dST6bJglhEnQQMu3thfn9+Hzq9JEMFKAUKBeNp/owu
gXN8i06p44NkDjaKzVhnMoqDck/CrfLQ+qa2uXdgYlUjc3uQ0MJcNsE/+CH6OmbB
SVjF/+YG5f5KNmFZKpPgjlpuXax1PNVxDtBd+XJRBF4tOeHj1QYYpZYLGgV8ELtT
EVv0vRemqg0kC8gRyodj3ulSKiHDCi9nzm11MmqI6h7k0vZcoQNByypPV5FBjqWP
NjgY57yrA7+sC51WsirmL6vjYdHY13RjOMKODg+Yv+sm0/yFKChfLiW2DBq2fBNz
MxABQdxHHdtB4Owvcke9YAzXoV/pJvY8CXtvRJ3f2sVFS1cDR2UA0cIIOMu4EOhy
hN0osNJt9Ez2fLLKsIevViimJpYeQEvefw6Q4eW6+9aQv4LUCMcHZSinZ/A+/AWU
TUhQu2s4A2YdSgGxSt8D8dbq+7PvWPjGiz5q6cwylq4WsCYKlrFbIm20GRlXf/Qp
qdmSkYdmOtWGGScfsuJSHn8D6fGDyYbCBiCql3t/AXCv44dQgz0k+kb+0+U/M51R
srYaliPG6anEAKTnpGsT0koKyWFvjerkJ6+RuqIube6m14jH2k0LRY4s7zODXv4t
YILWLIXJFrOfqBcOaAS22i2nBQUhlDj1tvTcg1dzoyWasvpUAQb5rD2El/WXCxA8
Sd+FCYEgR30Ia54eeIFB6AcZxAEEh9W3lA+UGsqFv69KcSzVCV5UEzq8uInyqdB2
bcxQDGVgNF/HjHUTQEqaLVf0Iw/y8qsSXw9bcVsDZvj4n8S8Bxu3vqNbcNvaaaU7
a0QqXy05HEv93KUEJAyWv/t4mtTimOagCjGA7GzlGO759JZ4umCIutZ39uA3Cf2h
tfKxNefxkYG6SOwV2+6TabuXhT1m0PsqV8T4+8sXO8av9NMRP1DEPkuSQ0YiLJKT
/nBzLKePqmHPdzId/lNWrVYifiG8hkwlKcehX1pHK3cOJkhTDeMMcqR634jLTwrH
3RNa69wKx4omCSKLoCJisZVvlKCN93FYB4FwPflo8so2ideGy3IKKIZDMf4LRcuB
/Drg8a+ffyoo31nQO2F9Gg7D4E22ruQNdsghmqz2hBZe3sPqyE2f+4Hv6/Eb/P5N
L94GexaJGz5FhMSka0p5gFCBTh7wVCrH55p1XNningILbOZtBmPfaW2JAkrNX7Da
vSF2H9TKuJ1qpHgByeSMzeqPAg2xIja4vYDZoVm6GjGpstcat2NoeoltjnxsU5PU
T57Y/y+TjPfNHwTAOjYga+dqiKOfYiNKogyZQSsZiBGO6dxSfOHF9ZnWdJdb6Big
ujQ9kIn8eaIrMqiFf4UHliTbMl+PmsKoQNU5e8kWVfHxJY4VFPKB73fauPpgHSsp
t+THZhXLKLI2zR5Hf5pTByvuaalHeViFT/+ygivkV+t8IYoTE+jaPh6Fkmf3XOe/
oQFbfgcV9ndXpB4ABp6yqmnEMNuTNR8YvDX/IT6KtTH34Zwq//15Y94osg83x0ia
BA7nnNSljOg2iXchrCqmB16LbHWxHk3Yu3Hn1YrxipW6H2NJ7O7p88v1YJvyAaYV
yu518cfMD7T0Iz3sKc8tFZGIfwr9YCIdORg/0wOgnu7Wtu9CU/hP2c2QOAKkr/0D
WUFdB5fjwVeJ6F51QpAGbBP2GqY9Y8RbXiLkvWb7jChCQIZwF+0D7jX56MMWt8Pn
C5DfKLbKdDAuH9zQzYGQB1c3qVN47tFk4YupOjtJbNd2HOUdxf+5iCnWlxNxtjpa
Hgysv72qBr6QvAa6oE9l9hF4692K9KN4xRJpCBsxJsyeBun6mzZd43eENt7icCN0
NPIybGjx71UOS5I6wF+VJYUu2vGwy2pZ0E8IIk3lutrUBpF7yyJTabgIxdfuS5PJ
N3bZWcKPAkvwsdhCoRQ0+D6k87UBxAMuY0oQKJsZ5KN69z99ucsavfSuaN66EHWB
Ol974sT5Wj+JjB8hQCDYdxYPJzONtlDg55VQAqDHlzFl1qEldQQLIklri8f/Ibj+
n4axfbsUPXScYWMYoaxbW0E2d7HZT2iYgLjPjbJe0StbqdinJTm24mnSwoJxG67+
lyPCCAOHfIQfMezcSyIJWT0tWdOdqYiz3s0JaTJqqoIzhXhTZMu3OgxsC9HFWzk3
vE8i7jVHMExHEg4SO/CRZ5i6uv6zuCw3IXPnIpWawYmA6fji7Yi8cK4rwqqzJh8Q
R/Ge17WgxBVXGRhe+L1hPFMaMZnXPS1G4TE576/vZwKIZLshmx+2QLh2pg3ufu/0
4VF5RjKkclF3ozy7j4Qa9hcg/gzJkoFjReU17NTv33+3jzMUxghheqVMrZ3VFr4P
sQV786jWG1qF3Eobj+hLhjfMyq1lYSUD8gHmiqiaGkPTdxzylgyH+zoU0eUaBik/
w5OEoGkseSoTzzxV/1m9cYwkNxQSRh/6KYLYJ5KH9cTInccJ4jOao7+3AR+kjRoM
t1ufv5pyxVniHHMv+wP3selkwf+OF+ZF30RRSKdonoFlCzm80TQiwjzv3sNI369R
x2Vp6CU8WCrWFltEL1hDeVOqWINaOkS1BF4DkN95C/WMAE0HnAdk2W1i4pp7qzGS
EVkd2LzFa8NTZNKmCaBk+R6XLwrZo06B4eQ4yeaDQ0iWJMmRFcrvOVvHkfeqHT8c
tWTIkZ034QlWFt5UI2cwL/sQNmGKKrdm0pnZktKM52lvufnAAjIcs5xKeLCrMI8A
25YtCTXOhi+NRGIi+v6MSq2o0Ol2UuJ2iqf4I8ldARD1D4T40dO/OkxlUJbVow7o
xKWYD0c1qiUZphAROsrHiudFP2+fPKofIpFeubsFJJ6XX6MBFHMnQw6k0wcOgIWc
cbgoy8ZD7owdZ839e9q56ExzRK/wWE0jIeR1eeVitZtbJ3zZELc5f4cSFFhnhx2c
3qBZPuOIDD/K/d7VCGYkLUmc5yyR08VOJ8LohKX8DXEXF6sCNSh+4vRvgg+LOysr
oXdFgWR8DEJ0fRN52QNT+R5G7WgfeN14y+l9VsJnW6O4vaoPvBt2uGPZfRRKuVX1
yvZC1LXYfD/zgoCgZgXWT7sO/UAUjPYVWQa00ots4y2ka/Ki2kae+JP510FWKeaM
bzt1uADXDYzTRQw9UUL5145EiEncygzaxjM1YcXPer/QG8fPOPhL1y/f8GEbyORN
8k175l3EF7T4WeQrY8GEyxJ9k5jJHmIrfyFacBrO/p1LPw8fPvK/7d875Sx6b5fS
mXyVzGYpnMrYfJxZ6myDafM6fIiv/nq5CXvGFxVag5ZzG194jjYSrR10hE4inTKx
s0Xvr+9hOIwbemK08KEVNipZAzRmB0rR2xMerwu5CQ0K7TKujKm/cxEO3oVewGP6
DaqWxsdOn1S1BJlrzG+rFCWKu1tbSNYrolp+znQ4HYNSyAuIURBAXdHoaCBLbtBV
LbWZFBYrKPH/t47xOAZZmgxXnMAmiVnXFJxsW9l6Uhv2fyb5BtteykN1gf+XcOUa
s7AK6h5DUH1oijG8tjlBRc60jWiZ24vth1TLbLNKPz6LGNrVGgHQLrp4PSd2WsH3
jELhSak7QIK5t2aQNYmfdv4CvOhkxi5sZ8NBbrthqWa2+nRwvU57ZYY5VGDIsB6a
eZ+OB4i6sTRIRR5SrDWIZzZ8p3gJQUZzk+he7gvzzGcZ+HDUG1Nk7mH0UF6BhwMx
8cUe6Z54LsFfLZGk/Lv6CY7LB6MoMrLbWY+SvRxokwOAMdcGNwWmaPhSjaZ3Jf//
za6ELLCMs0dlaUZYjcTfgGsURnlbUuqD0y7dxO0RpgUvnqJH+UFqZ9hr/tUYxPoh
cl2ph8928Uw0+IB+/qEfPFmkgYud/urq5tGNQgGORy+hWOGoh9u39XcWPbso+WgA
bowqxMdYlB99aD9Gc1I2Q3MOam6Av9YsIu9bebNDFv1qyKdO2HYmYYo6fznSVYxE
Zf8hQMihxHZhJH/SD+eA18airQWKRUO0U5XXZFNCnnibH8UrFfSSl4JpqAaerQ91
7XaOlOR37LZLDMt0blhrM8tdhVTBtplS2vPhbkF4ARylYmWGLytJ65aDB3fxaygD
FZvyRTMxWzI1qJPiV6TPxYYg71R1cosyiUKBg2j9FrS9nnaqLHiBStcqQip48ITN
IS6JOauQZi07gfie6BUHJQkLUtO59+byGwjLjGgacJG49Erbr9jl+zLpNAv6/InY
Tp97epqGiKF/79bItibiI+BNKpQwfiqBEfcJiigY8lz1Mp4/5vEg18z7riE6sTSj
GGY+korh2urDwXiu3r93EVv1O2JaPuNAqy9VZvT8SAQ/PV75A4GkIDZ7M/T8mAfD
sIS8REnYCga3RgzWT7+KpJMMnt4J2Lv2vHYqctSNOR5w0VTg5YkXzYuFrVMl9Lis
ZNAlYoisbYYX+Y2sHRKZGEAR9N6wZrxaHHU7WyjOj6R72PDI2NjVdn6KUQNvDXc3
g8pT6S/xFUmZM0P7bewlXgjUM60m+yLwrIGQfinU3phK61stPnISdPxTOjnkND1e
udX5TuacpdaOYH4P9vY3A3U54QVqFdr/FKTO1gacytpAM6xXowsRJ7IPvQFt4oke
of3gjH+S1YCUxnklfReTnPH6flslZyomIuoH7WfL0YUrd4kzwxncdZd6HSfZdXds
P5aavBTOt21rwA9b2B3n3H/58W29FQLwzJXSvndz4huRwUPQPHc4+0Y409+QXvkQ
AgjF7ujeHa+NTrhe0o696E7DXwTJgqifGoOLysny6edQubEdO2xdlL+IaBzud+8b
TtPZERQ6+CgAFkDlkXlBW6UkBXtS+EcrTAN9nZ+NXbKkJR4XuurRdqUvb8R9Jhpd
Twzz/QYlF7jIpFAKm9XrYaWzQV5yNEbGH0qMqksyT1tJiIMKzSdRryoLBEog05RR
ElI3crt6c43RrU1UDYzBLzII6XQvMe0KHqnqlnKW6wINz4Spv7in4ix3vQQ2/3/O
qgKaFK864yd55l5A0Mh0TSiGvnGT1N1MiAQDs9y00utPA6kfLlQgJvBHrnrNa9sv
wN4c1M57qQycoZ9oWTwJ328r+Y16u0p3eEAIVkzaUjelxkqeeptuA+tqZrjO8bJo
aQRxStE6HvywZyAip/EPqcdEggNENVzfolXnhpkIn00aNfQpcLamZGQepxGbK2pr
yBCXUBorbwiC//yU7bbepZrbb7GeIRBVrxQ6WbAfnd2tehSLRkXPY/8e+/fkC0mC
PgKHgQP0WMsjMUztLq/sf4R+16DGK20X4/T0oifBbquGmm785QSWzRAZc80XHVnJ
G0aZ5ZkYAVfENXLq61zumJZrwy37XGLeUjmUx85RnIdzSEIIswhS51Ag/m5/r810
pTtLRzVP5yThn+lTky5azAQRo6R+TwYSEnClzt1bFMM7cFudnJtmEWxZJ20uli1L
djqCkHAowBdkhveWErSt2yCXYaiUFktr6JbQc0xTHJ5Pdr3YJ/5CNDoBozCKoMYg
nI1iSYKmsAie0cbmg414jPu2MY6sYy1vnuieHrE4lLNJ/RpAlydGD99xMViE5KM/
tVZZqLkz+g7ZvcVS0AltD9gvp6oMFdTxTpI/nOlTr579bJqFwRIiCMLeNhPXSnrt
PnhveVXIrxovkakp+P/LIODlNhClRnT7+s8Or5NGO776kSjmS8WLwaz7fTiGhWB4
4pRfXV6j787UZYMp1u0shzdwawiELXW21L5va3I75Iig0RCapSiXDXT9HDENcbqx
aehKYnSO0fNqf71Y/m5efZMsxhGyksneqRoocSCoUOIa1LTjS7MqwU8BppbH1fSp
9eToDU4Lmui1Nj3mMJQlXep5NSrQFp5SUNR6Merz3CvJBmQoaoYhbpx+OdPqnTJX
pGCb1OhNeVm2coNbUA3Fh0joe9DU8yAqrKzbbmaftGAwhwWw1HXL07UybH91jL7t
CdxBM6zPvdgVtN0jQbZ98h6jmYBMVMl+8jWW+Jt661aNYH4D2uWvrhavbK0k8nFH
E+Hb9ajloSoUM0qZWw8kYTIrz6EmY0mMmA0Lz3YnbtboFS4Qd8+xO3WEglbBNk4v
vE7dUjRnYVF+57A6xkOKCwbr2IyBdNafO6xRiQUcDAOcoTKFimgQGCPhvcaIlqUC
0Zh3vKZmVVYxt8E7irqGyV5sjxqb107DZn2ts675FtaJzElxm6zhKGrK7D+6eYbE
Se1ntnIPDubhkECV4RiKDfrOS+PgPdH3AXDfysbakjTdyI4nefhWMeBEk6KANpcB
xhaMz7Bd6QhVAhhs3wSTfgcIiESRJWAFvBhMqWl8aZpnc59op8+ph9HXGE4LTm66
kVf1swTojwxJEIBHax55CdPYJbbhhmr9TzmHtiwSrQhAxEEjfg4XjAlPw3QdiECM
rkIzMz3sMDL6c1hVSeQWLxuiTORzUMhMaPjzlrSnEUX1UUvcQn0H8VPcYAL32NBr
3I0Ew4P8WbZm0y7jqDYjJIayY54TmolqwV4GUW17aAlrUCwUj2B66P0FojXj8SQ1
dya5YISQwLPbXGzzkyyVNQBXX+RLa+n1MQhJP1e8NlCUVPEhxNcSL4NFBVJIWsJe
OFx9LIPvMhoPe8YG2o/sXP3PkRnc0aoc4kMuVB7j9ym8tevh4fZAM6aT4XBYonEZ
P3mScD7y/K5pbZhonnmiG+FPmJ4Ke/LhDFNU1TcQyD4c97CZEu4YyeuQMqpKYt2n
CJ37E3cezMSr3y7ysUkq2Nenv+ADgX99/r35JObhQxZlzSabb6dJ7vfb8hg1+VnJ
Lfo0vyNRbF55G0D0GbQP8VABiLqeZ8WEmLNFGFFpo2fBNevkqyZ6IJXg765Hhq/v
UOkITDAiR1IorG7mqnpmXpKxgGYQV2oUxyep5qzdCRgRqHAMOPZI/cz5U01fpq4k
fzbYWTiX+z9SOg38XfLZg6fWAGY3ISU1pGqR+RllLqKbNHXwmRwSUygJaSS10OvM
nEk0XI5GMYxLQ6GLKkPyqraFKaBROljiQ8BPId2s2CYNTPNAwyRzfjbMZF7YV1Zn
cVZl3Bai488UWl27skWEPXmyz5+fyKGZtTRbg44yr/2Sq6z01EFWpiFqBne3rwX1
SBtUGv8Zgtn9FQblXuK+c/HFavW0dN6d4XwqHomLJ0NkhVRArpwWmsGR96er0C41
syS/WxIO/5ubZz6euSWLRBepQwL8CsLwcEYcEE22yEEhfbZW1fX67yMlxKw7b77k
hwMKdLn9i4GpyuOYzDDcqky/P+CFyhFlBbKmkW4y+0Y1yl/a7FV3C7/UhT9i15ZQ
nDba96RRSPsolcR42fjGwocil12HEHGeU5Re4fyemtHNTzIeEt6MbW/o8lLI0LCV
ppvJi0LkHY762K6aRQL/vhROFQMZpG8mhdIkrOG1eNXlaWqlfUQiU6lCM5cUuweR
wO+xSLgiH6y211Zbzc4s/y2swLKlJmAiT+REDCTRQ0ZFiCkdtZtBvuefUEsEguKo
LbEGiulFgkj5kEWubE6KyWqVOb/RhTOG1ATjSFQvFoaJMeZP/WaGsYaJ+SyGGSAt
1fvCYPSOXYOSYdLFmVcVYbKIbG4dr+Okd39GYDazrEkKR0zKXU9R8KD6Yv49Bhxg
gC0xA4UoSUxqvL4EFlHhQX3GwP2b3u5cXg+m0gEleE9IYQrbZDDAIeurxXN3W4Ov
om0zq5c+27aFBbecsQYWQAad0fuv1ibi3sQUir3uVfN4rXnYHDKB78ACKbOv+qPb
0dIA50mv15zF6lswUwXAcCiaXi18ubCPi8mtdwlzBCCl6WNkPC5lQKJihCb7ENDt
1DjqcKmwCzorTaMniDr1JaSf/qOYbLk1RqRAzil52afjKeGlqc/WVVrZpXwuoPkC
ftfZ+TnljmuzU+hdOLtSUncOaiGkBfL+rg+PPVuSP05K8eghN7RdJZA2PAXxbaAc
ZLGj4rp63M7GKpaAOyeyCzVSxmiiyNDTzNykujGKnTEawSa6WG4rKSW9pIMLEkeT
HPwh6xhcnuNOyJj2FJGYXAQaZkKUrVcBvnDZAfGLnZkL71h8GJDLOXfyZ8zm95Rt
eeODw43nWqh1dqOCgia9BXfyz7aBVr9xhx7HrySpjRPzqvXwvhoGNHhp6R6Z0tjG
mB8zk4HpBy18eSHNJ5EHsM43uQFLB0SlTt45Akmf9uJpgbI2gM8eT8UiBZWqJxFj
q/mP7UHFd7SuNDv2LBGLGKb1sI2Jf/1/iTV4YDz8HYvWWra+MND17mtOiWJ5IWGT
bU6xjSyhmoDC2yglaUxtdmaLmbASvQrT/XmCgrgdXwyD3vdNDfw1uml/lY01aW74
BTagy7dgZ+NEiGYJAmhcMAXqMdqoiLAr7H5MEXjlaPn32PhJS2/oa6B9HRHF4n2R
7aYJdtTo1wV1u1R/C1yNw5nugB3Q3lCVd+JlMQ29QMnugwuKiySv2IT8qgzDE03b
W9Bjf2uGn9USCXlFxXKNBsRkIKs5s7ATn81xYm0CZnxOkn850wtU6cs2KR2gq3hG
kEEZLCpAcyuQkApewTtye01hj/7mlZ9Jsl7POlQg96JLKfHxLKNy6Er5vlwH4wen
jJCMRHo81NmH156SKecdue1/OWEPclT7UAQSs/ltKTiQjNoqAdH3OfdenhHNwokL
GPZBC4N120JktioIOxKCmDTKfu+fkz11ggCFkduyWLv9Lavh8EKHY4p6ezfD4b8Y
vO0ana6DFL033dEeMS6DEOLKGmV86UiAZcJkKV3IRpDz/QWEZE4P6SveGJsPfUjT
pW3d556oh71LDWlDQrCmwYFR1mB3aqyfd6k5qpgYP96zz0ECSGFEAtLuqCbgZxUJ
EE8zqzd+Ggdg0tTuJSRX+z2mjZQYSiuTjoDOuhC9LYsvsObWLHTxlL7MA3yw/VyO
KuymH8fAQxorP5yAAkYP1TQGZrJcCANG7ZKjNHzTIFFyZsiq7r75d+Q99GmK03dW
IJad5gyouOEVDFSuB4KiZ6Ev0egnecRwzmApxqKR1qOcUeDLQ+7r+8YaazLQJHNO
IMqDj6w4csEgHeoAPWMza08vsdYTPSVHpM6acQphHDtlIAKHveoHUjdyVW+1VKb9
5TNMatwI5HbnSv7zLTG3iiXEU/sr7SLyra1N/8klxHf1NEmXaUhFAAF9E9POo8d3
ECX68HtHe2Io3WpeIbLla/jXskmUvFn8J2QxIeG6n/qq+O0mB04XYvWQs8rPB0hi
UoPpRM1rkJaOgVIMYX2UBcAmQZalbOD02MPa4rzZ4tw+MPfDgMnIaUDJijIDPqe5
7/ePuMO4h0Vt2y2ggu/M0lTAihBjnovwBt0IQIKLqD/STFrcWBD6vx5sjTo+AXtR
Jj/LwmCdh3Qi/RrCwFOzjg1ZQ+CvJgNiMmEaMspht+sFb7VQAk09yXRmgwzs0uja
Zd9ZgHYg4IGlb8T3De876J+4O+FK3My3jzNnrGSpCyRN2EMm68J8/yewCbaD5mtK
kDwELW76bTUL7IY0brQHKbNPPOxIOnvpc1nyb8bKLIHJO/AKoKt7Fv2O4Rs1ou0h
bM6EPgCKPuO0xBN7mrwbDFIqZBvRvIf+OnFOMRnS9JkqMDb8CHgKH9Q/mW4Q1Lt5
gdopusXWFyI3GhTz3YWXf4eWgOkj0a+rCukE1SyRXpfMD5B3MrLFy3n/eH1wFXXe
JXMpB8wKbo9dbnD/6JqYgWE1/P+FnDW6Ib1mntQSKX1MGjIWCytqpKRg1y8xrN7Y
asvfkW5gmyOWkf0L3pcuiq3jiRzYkBWeRyV4qDv5T6ry8qUVdr4HridxzA8q3WJB
Plkz645B129VDjkg8fLndBpmwkGZjnkJNtvx2Oxg5NF02v7i6+6B7aPsnPVk8eCE
UuNMJDhKivR7uvX3kR03vfq8oYPeHP0paiu1jVrhByOEyt6nAR4MEDt/zpHhYOYr
R7GIHx4bzVnJknH37JARsh5mUsukexAUMP7v/IpVfgzAHnZmnZ8YtotI3gvAp6qX
GkLHwjaYm+4g5yq5ph/xQlG6bEBnRk+hVNnWIdkVPrzD96LXgxWt+0O8dWzxp0Wn
JDCJ7yfmXdKzh9tJ0nX7m/aoMNq2lTFZSfhC19A7k10EQlgE6sLzZIH1TOYhyk3X
Quu2vTt2OYSKPRTJKu86cgeYdCZm04bhVp2eH3Lcxy54RMPsx8ngG7kW2LmIW0wJ
oqdZSoTVHfoo378cr0cmxiNH/DtNsX3U4gtZwiFHrlyqW3C3Z3RFwctw1yThRXuQ
CG4TeiLsozJrDrXPJyNFEeTq3Xghh2Qvn1nYmYOvk+BwsOsJgntBqTVOr1GVmCDj
4zcSBrinj1gqTcjH5Nbwue5TtFhTNYQqpsJDx6V/RD49ZHmHEDmj58wzV8ljQKMa
55m5F4hqhfNcgLpv7WKvzv5qdWUNWl7RDkxKZ7syPRc3gwr2TizHOqBZKelQAUEn
hv9eTYF6EY1dqgG1tJCy3iWlyFxrQX1sXtMVICMWfshEER5bvI+isOfCmiBDgxDk
UrSd/iqsuBdylgyZVeTTef+NOcRr9j0ggoufWaEbQGxmMHblDFsMoaLwhWF7DON/
UOLl52xN9YhS/+K35PS4nsFzUwdhMo/cnNl7a/8xelzpdflKarZFCLPoUB5jV6B4
XMXyIK56vZxf4RNZAKEDkMp5BohtP4QRJtwW2BGFNbUiw/vfhToP4+JV4I/tIYoC
DrTVQC2w5suyBUG/vYN2dSkLemJ0fkvkynH426wzTbhzUPgbNhQJI5OOlivEMWsk
m1mS23rgoQt8cSvRYrZeb6fCo+kFrPk0c6hhJYblf11Bk9EGA/UiuI+Qb/4WFOwA
Mne1wFDuSQUGcsk6SzMzqHK1GVGWc03NjmKUFuph0ApbmtcFCbRLIoa0SkQ47lsY
H4gKoFj2z3uFc5DzS5jZr0yCfk/b2b85AIZYmornorXk23Qv0mnaTzUJHJRPoAM2
z84KQzcVH8CD0Sat34CGZENfLk8fRMjLldcDAkW9ctW/MufJKomaBWPE16YUxhbr
iJUXkxRo+v/B9t1zdEami3v/3VD2rI/tXw63yPcS2/Ja5eTAEgn1YCWxn/BKP2Vm
iF8+fu7M96zCQ/3lWy/YPqo4xUB2lzRYNEpd6W6r16hTqgGIROwXunCGOX7yOk6Q
2aBJ+cXjX6lr7dGj3SvRf+e522zTjFF5oTAjo3N3cm0Kffu4ztz5MqSYBVTsxOjD
EdK7CE1coJZgzbMtawfJbliNwmJKm5OLGBoTEzZi7M9JkjEKZmsUGFl+RQlPMQ9b
H2gdQP/2qOI+aANoNgH9qWPosBHmpMKByU9p3kFCtVLT8mt+y+8ggbNbFacJB+n1
AnzqRDqdvAp1i1b/Nd88gDuyyxgFPUmWLSPvUqjOodYNPJGbhkvikDG8FoeCgUjC
ZOPaVQS686Z5EUyvKygEWae1isI/uf7GncG8BZNs+MtYTTjlJcLI9k11G06R0KvY
QesqXNauLbb7vtzk+ll3PrIxh0gZIBJSsUPfnJemuykTI2w31y6VcxtDSFC4v3Dj
j031NjJa/J1RvQRBKwoJtheXDV+Ku2bhCpUYDu9k7FNpNlhgp+5bKYtlnsTwy7T7
eLVerAyuvE9JTcj0ZFMDyVLG8e9COd91FlnIeFfBShmLP/EswrDcIJAzDgyz4O7b
cdJSlmlml/GiRjrBw3YNuR1DjVjrgP3esUMRmZISkxIBLbGda+OAGfZhCROLSsDp
HZTTYJVcLecqsPBMF/iSmkxcT8u94BCj8ie/qDMw2UZTuLl4OzryN6Z9OQWMkDg7
z1TKsItXUllFWeOq51Cyi7dX6VZMz6hnoOqOI2JZiZEu/FNn2b8EdJB0obFuUjY2
IJi2oiaYRizMAJr4LEeQRF7WT2vwzAO7CMxMPlM0M/cJJV07Zl+42EQNs0DqkKDV
kqCfSd5UXtLI3yJXJRxb7B/5rQocWFgDk4PudHOnWDCoqqkYSa6o0bK/bYE4HZqg
b2ZxLRX2d6COBWn8MmtEnSLPmdEuJU/hXe/iQfbSoEIAh0uZZYLlZHN74TMptE1e
sIk+km4N5hzVKLkZjpxvxQaT3q3ABJdSwZF07IgSXXA78Z6AL9Kp9FrEI/OqIZOV
nLzpAN/AcQHRbI07S1pRr9kTBtZbe1occhC34CZAv3phk+fa52blx1+SMCm0Mruz
+X2XlTb5XYBhME5GgPewMRzZf2NKQkve9GX4/gtnPOt/QXz6vrKYlHnyK6ClEyX4
qoNB0ZLzH3mlPb/eA6ASXO0RgtfR3SqynbtfpjNVy0OKVN54PuN08Txxp0s7QVxg
Oy8yhlyCtEkWBBKxYmIqNND3kOGyeJK0KyOmGNmuu8Xk/BQi6i7kuZOC6J1SQ+aK
RM/Tdiuwj3OjWj5PkPewTU1jO3rEIhNSTnTiNuRZhK8Q9PCuy/KDQC2kfp3hBbGj
dEFzQ3Lnc364Q2epmXCUXuIRaEUtjj6HIstLd03UcWej6gaokj4yD6VFr1a4zPQk
mvSxY150NXaBcBTbxKIyxWstlvucOkqFAF2/nhz4fsOGHatOwHTA0ZfPlKTZvUgd
YZmqhxFdYnY05QYFN6o1Vp2DX9Nemq6sd8MJPBGUuCiCMBV6eIqkk6ZmXcu0gGZm
lHiO1RHAAqo/EfoMl7xCgwOnwPYftDqre12LToINsbVvAGlypBD9ietLMgD7lUm+
sMlymBpapwpk7I68Xla10KYh3h/bLMnsaFsJeiSX+bcCwJyL6x9iLuLing/Zyg57
gNOwGQBr9Z9LgJke5QPATSm9cMUxvXw1ka4VkfvbzA+lmj0duPa6wOL1rCNtuDv7
qE1LRPCk5MZI2SthdhwCIaTb3JOQ0q5ol1hQA2Ia/WG+S2Q9EyHMfIwTqrB6dC53
Va48UjaupsPlyPBrlxvU/DKD9IS9CIpaCZBCIWCqvD79T7iwebrCxWySKCiBYDlG
7+7ykjdM7c7+eLJpLn8dh9oU01F3LWyOMSZJkSmkSPT5RfSqnjoFYBK26eDb0uE9
SdaV4VlIJq/LSGdtSEvitRqbVEmY3HkhEqLdNwuysq+J655rKEFwtxjQIbhLb+0k
Bg+SP9ynTSDQCP0dM423hvBASD+Y7lMQJ7yPyNYngD4EhE0xxOddifBTN2LkDAa/
W9aADSB9bWWH6bXA4O8aj+uQV8JOWq59VDQApfJ4vRTBx+MNiuv2W94MOF56LXsl
/eeThe8MmgpXKCjiy5KKCasTJYmF8lUmarejkfM7HR90oXVHqG0r80ZCWDY8+wcm
tT8AkJUuGFfDNGfbXDVgJ1Kn1p1SyJfS2rXPrxZah2ZTWfjWvDMDo5km7TAvp/FU
TuDXNZQeaNEcJT9wHgdTAGTSWAk9zc9BltHxEMkBiO85oT+PnsniOAupldFYmKZt
U6EdNY90/BqGcuo6GZF49ihLIyHqm7vevTA8n2yQx+i0IbDbGT4psTsE8Bo+pitO
dw6jQNKnvyz6exOu5g5/MkknN9nYK0kDwHRFzhpoGUZGGdbItEVoMXIW0SFdye1P
iW4ZCkQHUC8TvNaGFh4f5U3pN+XUo5irKfIin64H1j457T/EuCmtTHH/UFeE9NIw
oOw6Ch4mBRN27r3YQufwSw8/R6N87iwQAC487gmcad0y+Z0hpN32mQeiiBqieUru
cdjJaU3S+l14ADXz/mssqHCeB8ASPmRAae9iP/QK2fzg81u7JhNt8TEhWxmcAZxr
wBR2Ruor9uNZ0Fgm61wsdhaiHEdPjiDy3Waw35GcRqX5g9CZVJSLmIWwrEihcmiP
YImX+BEmAbWJwRgANFWx09IiJgs6/is6Ru3xqiFA7XtWhgbDQOTnudaGzjLj9pyy
VOltA3TS47nuT7ddpXGABu6vL/qakD+qUMlHpG6pXYhUuRxW1m2jurmDGi4CTx1Z
VON9BAIycw3lXbE4/FX8MUWEqzDbVJxoE/QChWZOZQ/oyksmk0we1VG2v1e0wGDG
k/xvE430F//L2Do5UqhLtBmrf7icyJ9L11udrYWuk+LQZkhyneQQ9kADXrAvKfPj
oawU/Pn0VALGjrNq546X+RdAvJEKasF42gr2nVAtuWFnMjP1AMghuVizJX515wUT
fBuQeI2rkwUaaX+8GXjvheoV76lP+qon4h0+iIp2o95jzPiI2PPRh/RlnYRPUbM4
W3+uOo5lgP6yq7bcxwe1diHaLeTwCYzhnL+YTq5C41Qf8w1GTqw8+ERSf7uCq0Tq
BISP2NN6YPpt0DEdamKj3/zecTvjlctUSXH9pIDcdNfEOvkcyqKBjuqJVtFOyFFG
JrBSAFad1HfkNwOOGfJrFG+tXT/Bjhd57g4BIFoHFFpa9ZQ9BLo7F5wqj2qdP2Xt
fK3bPJKCgiHJ6Px1sEzQb886wom3BdmIyPHc6p8AS10lzoCv+UszNzwmn9qqMqOm
s5wLyFr7Z8s+i9om0MipmjFSEq96b8qKy3aLXLSmgowFHluEOHUtGzRLlMqZsGgR
bY66JoO+brtU34TJX2inJwXNxt1yjNeXGMxF1hf2N0ZzoPXTrOWvOvKad/vWcSeI
i8cd5AJEdPxucy7pcV0dVU7Z46u4GQp1MicIxrkRmpZm+KZjT0CQxTQ+6gd+vcJ5
wgEQ4DdnUoxh3WVnfdAOxVqnR9FwJER762gF9VLDIrsa4QPxpdqiHp9MIlDE9nsD
MmqW88iA80Xayu9/l4OTJejYjbVQNaOycL6U8BCHnZyMJquT3zZOPR+Y5gV81z/V
tc7flDrt0iZqojnVi/+AHDh2sfAdJho35CqsZmCf3w03mAxpRMXWQf94rLVsjLzU
SnsPNt2hS0Qp6eZGboAD23iNrlI8vOrpoRd/A/NMmb3I3UhJRge3udgnqbmKBTRv
ByWR0FChpk77GwBQgTvBtgo4IZdm8w02YISBmK5AVuhFwGqVw/tN60GzN/kzzWgP
JW8jDKtjd1fo1I8L87T7BhbFei2SzaZ6hv4+bbKZohEjQxQLZ7YGEgsrPQo2k9pc
iaAyxAX1C6qnmphxSVVs3pfOsAex90Gvl9fRbpDh1eCc2ajtIsxbylkMWIsRL12G
mLY1SgsxQRdW4pFJi3SQ0Nn4vwawxxg4Tu2SNvMYzW4pqdaiLLCxgFlSJEeC/P0C
7Fk5UCg/67zNJttUvDIZ7uC4MNgJoSJUDDmJCavs8cZ4QqrizSU3N//dU/Me+Ft0
9JO5zFjyoPWkguwmcGqe+vDzwRm0cMhQUDPGdUbHjM5C+IWasZ1HQa+Fp1Sz43kz
IpTFqYznFHHyfifW4T5gntrW0uz5hDwwydSm1P+1v0EVpc9AXGuSOLHXtEmKrNfh
XpNnGVYuAB55DqpTxMKWXhEq7hZ3QWfhPcoLECTAZ4BHATg3JLK58CHxEekTwPcR
oGic0zD6X77JD5eXIsiNq0Pl59z5nIElR5RlwaoF4oLSg0wS2aVPgGtoHqNov4l3
d7s6mQJy3LOJv1z9DYjYWclqxbxC7TQ6RA0KzDisLeCqu+XsrEA/8XY7Em0b0X8g
SHZat3wL9mPkpejSg+eu8jSqkHwSY6E0t7DO+p30a6TkiQFhBYVDGPhhERRWDm+p
iem6VXSTr/8m3jk4yaqprhAnh8ne1e5frvHAHbsfsmeHyTO+sUc7iLZj8sg5iaI4
hJoyNEeLbaw4eMekVvERpT+2ymZ08g7WTrHv4GF+flkW+Mo9263njU4qmhTuPPAD
r83y/7fz6yUKFVpH093GliCC42pc5e6l1ZxH9VzHAnEUj8LoF/hknH8uaddx/+xa
mWcE4Gr8VBhe3iDhq21NiJBFqD5WuhtsRgxNNn8iDXW3X1gg12QjGYgDzx+MXv5D
OBhQzQE9d7coA7RY3OY35HvVb5Qx3jD+7TDRDx0FcQsJmby3JVTajiKd4KgWjD0g
I+AiHggx+ZTkL1MeZ2/MWdzC0XYE95vtqaaRl/YwmittvMRYZtU5nwP5SLhjuf23
PRHV6/nNRRUG4VX1fMeui01NxsdidFeyEYBb12IrhNnpJrUwpzoVB3CEb6BQAuFr
IitQkn0ivWl47HNp25S5dcsauMFm9c3o9o6Xiiv3jnk8hH5jUTPBznrODzxq7HKM
RU4YalVvpTS0VNUs4r8WLP/3dWIXtuP1gDZdt/H+nQDKDJAqoVjCnKDfEXir5iYk
Gx5lazT9XynP3cakID2+QEMoJyG+aKyn1FZ/1vb7aeTDM0PG9meLV8QSndyDXhGd
/cTmTvMagC4dzpf0MQIYn8pQgV7ab21VFhm8Y6DfnLg9Ds5+jD7bEsIeMEREuQYy
MBYPkpu6leG1IQeX5d65C8S/sqfr7CcZg3Bx/P+CPpq80H68lqDaAb1hl0mGJzNL
E3zgPZgfv10NAInyrRALEDCkxpEM7gSz2OwjYiG7PfGKZollpx1yBfnOrxHsGz4g
W+X2+M+6kmrfzm+sCIHhViYnnTsjCL2L9tyU1R66HnynPPoDFVpCY2953ooxR/OJ
w3X/YKTT2LSI/RQsMtLxOdw+WYHplGq2fPDUKahjmHFtjJ3C/HbbftMsjAlwN9wy
zGRd3T4ee74LvoVbUSdBFiPv7/KAtYEO/lnEu/kBMqMTOKTrOSMLzxBxCp18yObN
PlQZEGZxFFOEawRzcG3xZmzJib8m7DcKa4UReLure+ogPTqfIDnxVA66JiLWKRrk
2wZdz3bLINVInSTKhb0Lw3p2LPcASrI0/D1HTGt8+jTNaKLyNzYhCA6y1Un1u06T
TcnOuhCRZ3TPWnUYXI7oKJdWcxzhE+/YkZ04hjmAM1lYiA9wF8dr1s0d4vBgdElG
xbWLhBoSLBVhH5EHZl3LaLzTMGm38Vlg0768QczouccaqU1gSPnA+S4kt/rB0ABU
S9M5kjQFpOopKmWlBdQx3KQQRRPxFwZNCN4uKKCKVBWSm2sRALrrQvTSsy/H41yr
65Tup/rACz21IesyKt4+L8bvSZPsloP9+Xz3b7pp8YY5+xpPLvC+TNflbMV+++uf
QrSoFQUUsDM8X2S2+BlHD3JAZ1RuR0fsUdbZXhxPsSjN9lnKSfWhonyMZkuAB/2z
+PbtjTTxN2uJektlq647rvztX3HoAOJzmRSvICpZjc0HTKvXQ/DU87X91JjAfbUY
QgPMe8C9+f9+2eWfl+/P1vkbp0pGmoxtO6kx+hvzvWMr85vK1saRwX3Kpw7chVCR
QS/sFmzmhUIW+yHjjvzSd14hGM8VWcu1vkACUgm1xSRNRVXz0SpHmJxE6c1sTOJd
A6WduZ9iblsa6VPe7u4Fw6DlfEiUZRXpkCbYXqn7kg0aD4mVdfhLkteYvs098U43
Wx0wiHwjBrnsC2suU1ikWzArjkCczp0Gs/B0meQ1kmtwEnBRcXbFGL8C4vOVHqGY
D8ZDP0SSIchiGex+372u+ll49FOOkchCUKIMGiUBrnGgY5eMgH+p61YBuk8ig+Dp
jqOBHq4wgVqB/kgJB0YD1BYAAmHJKnhd1xsrAjBDeMgjpMckX8pZswuYE/PlWluF
VetDt1O9IyLuerDvz//y57jf1uq6vv5i4yu2AXQ5oepNskaD+uLM/hH3gPayqAgv
BQwQRD9k/u4rHX3fGtoABKqA7l+t4/5r5ekFWyhkuasOArtNxKbM+XiwlJZKNYlU
Bwaa2KeFxyaCh+5V9yvhYtkPRxIFOvn41l8VxCV0zm4kg8Sq7SbHSiVyaYRTXEMC
PCSs5+Z/5n6z2tmwfq0N1kcRQGyd37g9RHFXDmXA02MY94kOZsJ+gHM3zvHRTe90
pXQLnRNMm8A4Oq2k2d/Bv608tf2wh54ucvwPiLbabujeRr2u814m5xWhZm/YiF8a
6MQY0q9fZZG3YRxWrqcaoXsVA/Ux1Vb4SwkI43ztQwpHvtDcWmIpUEYxkwek+yNL
f90SuarUIr+VOmzRquKr+Eg7uVGMCiaUf8e07n+dHEryRjlYEg6cIah++9xcJjWO
pEmqOR/Y8dbPNdzx+2B0XtsMUOApFtY1SJhs2D0z4a++EzfTHRyeKnh6FQkjCrTh
gyeOptYJ4/MH0WT1YsG2ve8HXpKM+gTjv3jLJriN++iNcHezMrh32gOpG9J177Mn
PdEm1vptLKdOrHoIK93RSxD4e2pe61ANBCR6hFslkgsYuR7N8UEBC7IYLSNn5d4q
hbckSH8sL1cb2PzpM3MmnWAgz7dnhYsvF8cinLb6kEmAN6mezQqp62CH1Ug34NKn
j2COROYllx8JkcYAYF0yAFRY/xrSd6aaU8bzCKPCBQFCVnaKjq9bjQ6JineMUeND
f9y72X1GS3VFJHSsSA8ynJflGGmOi5rEU98fwF1r8uXfLfSG9/uAYhNwdKql9ssl
9TcMP59478B3bOat9Ov2ZXzyENh45TSJ5dSWm8gtBxqsozyJXuNRwfurIwVOeG78
6B1YMiB7GpXZJ40eU6l1GH88fQCuqGoqlAazAagniO5qbqNu1wwNiq8KWaaqJnDo
XCJ4pSLogeYzQSwr9Fk5JWHrPmsw/oJhY4/VtcY60B5PnPlHmnXVuOwe5kVb9eOL
/NIXbKLqwZWcADz+rYCw8ubnwCUy3wGHO/zvXnFl/gE3iy3UBZl4R+CYdjlswMVE
tbL0jpF+i5ZdAcm+fctpC7hbAmWQLsWsCeWw8/7VrCZ5PQ0EDCuyFULq5KmfNHO6
MlCfH3RmF4xX45qvMpyw9W07Yr4mxTES76bcdbJyte3kcTmO0fg89vpOkQzFukpO
DkSW2Oib7mqsj2nc7BXhbREZnCsI6IEhQ8+uyLuGMfBcDj4kLMFlvYGcVoaccMAN
W9dhHJlVqZOycylbdcyv67nDdBi1y7fAE6KlqRccQEXylc+Mu3wXUzWS6Rkr1tYZ
Qv4QTMjJOuHSyMkcR6dyuPld64M8yARNfKzg9dq0ZF4TVBKOcYnqrfCvRe9WVyni
P9rF4mDdm8lihLYqlO+uM16c2dUkuT6qsG6j03Rkk67an3ZXQmM3aQ/XX251VVOK
84x9GkMNu42kZ107vce2GVkOEiQ9uvsulcsYGyrHAwXeH07nUD9RgjhMZbR/K1Sh
JjyH0SYUR/tiiJC5Ujeo8lOhbhOJfuXd8VFyngKC1shsQgi3Dwei8wzkxOdDgnGn
4vl3DlmrR16bX0GGGrPj6+x/kWJ932qHscQDZxtkVLQ2mDe02v8nOLpky/TckSKF
JbFVPzuPgdeNQ58ReM1rHHfiDtYSI0oKCDYkRE2ZTEW9Rrn1sPJW4wkaRiQlIrzw
J9/VHTSw76ySsIxP4fMtDXCAUk7ZZi0dMJH9ae30bIwsYKNFlIr4rfvralkJoDBd
ncsae2t0YlZ8DQkqT+oTWhTXb63zQh7/6ZXGBfU3VbRYQlYrbYM8KXADnyfq7gjo
1c63XhM0HACG/pYXumVXashGlaK9p3QU2PPdZKRrTljLuIePoLB6+IKVfb1fWJCj
iwdaZpiK0ilz8nboar2n5IJwE163T0XFCjfUi3FkT7H33c9GTuStSAGTaUwj9Vbs
rqY27lqQFs7NHKj3+br4eVl+iIhegB/tpS/7WcxGcdK92SC8nZKQuklfgGQF0TOM
mqt6M63lBL8CeHPopTdmw8RfON7dAFAlWlOushakQ4as6bzjewfKOd53Bw4KD5Wq
UkqcVi7MVJmsyC2jb4REhZL+BjzB8AeBqM7MixZXcM8GS/C+ujbCIR8XB006NO05
0HacTSZ8SRcivg9QBLttAcByDlA7i5hMHAipRA3nM0cmqh+hA0vSu2aVQ+VKFnDH
xr0uFcrNGvfK+koK4CVg9TQpWyX5sL9IK20V96JGKXAI5Rueo4uYgpDV4PnB+hwB
FD2KmR/QnnlhxV1swaOPq7EVIzZWlJkFtRle87A7/uYQFzF7EYApbOOBvubZdhsG
h2ok8O907wOsvASJiIT0Dp8nlPtb/8L8adzphXXRQrA+qhWChrjjjnBNofshr3eS
7fYhC8dpu55Qj4UBYb0AbnmGASEMJfFO3gIOdyVx2Jd/3NR/kQ3qQoHhMLDMqnNT
XojfM43dn25YtL2SF+Gftnw7cXxDeuf9nb1MeqqUNtzU94xg+NFO6tqlbbwUAIqA
Pn4GnXLe/bMGhrcv9v2//PjHv68J6PYglNPGLd/9x/VNMuqurtSrX+FAVy7uNSGC
cLOv86cDX/vyxn27r+yM0o3KFaKYnMxdiMfnr6YMTyVpFef2mSJ0E40g/+2I4WIS
E7f8xf0Mhqlgwj/kdo+gdeNlU/LgOg/KjAynnX3XW4tdTYpFV16js+coGzbignEK
rSk7/cLNNjCBp2pKleTkIY51awt1iS/neC1iOn79J19gySRMKeq0NqomS3mi2Zi4
ict/j15wqjOZVj3UHMV4A3r9mqvc+ufXYQZdL7XF4RQtw4E8I24oNtvYBEabfZCQ
yGMvYAak6ae40Tea62JJ2MEwdbMlJa9EaxRcctxeVhfXYbsx36DPWAtLPC1NcHrs
C5KEsD9Dj5YLk8i21uD3xrr5FRsDqXqaaW83O3s4LVZ4/Dg0Nwtjp9ogxRSd9v+H
JIxck/v/bZZPnzuTiYwfHhHcbtyrx/Li3pXPqvB5y8s8TPipYo2xD5F3PvzvgFcH
Ng1Y/cGa18lowbZy+2bh6VI+rXvX7ixaAwOC4UAkO+9qZ9gRgoMeiuMCTNm2xYtu
yw+ZfiQWEommO0oDQ2vuNoPyMyYt1AW9bkrKMvWw5WmRzOjFGbcFQL9M6AvcL6oa
firuLLhw3nyLZnzQVe9sHkrWTJVzQX87Okjj0Pn/Ov0j81vLFyGIOSdW6uEtei2k
k/98pjuKoOwDRjR3VMPUd9x4jJe+oKVaGIGe04M+Sox6XrEbXDCb7ojBBxupOUOz
swZeLmqW7C7lY237JyJdW9F9ofA2iIvveRNM7CqE1LzLKc6VkSJAxDE8AqOEDub1
e5N7wFcEbWUTvrm3cKtMOq9DYvx4GatBeidSwNOpOrofOu6V7vnSd/QOmvK+HPz9
7feue5uWopJnIPymnft/oFL0vfMRvQZdkbCdrMTMJRb2uGsGye2Jz5JiBG1KfGSZ
UDEtp2KSE27vtvHXy0vQCgf0tSPA9cXdBtvwheAH43mcpXJPfUZkUVLOj686h+94
KhJUG4na7Scdo3AsENoStmoiaN0w+hzwkx29B/vDzCEkCxon8nrhPxXdIqBr+GSB
FdFLF20p8QcE/1ZX3qjN9kK+NssLABydm7wSo6VMyEqROO7NQu2oI96UgY+qQRC4
+YY/2MPPVQos9NJp1OlnBfi/j18pyTcBPjoMjNH78dZlp6tts1Ml8LES87l+i6F4
tzJsk9dfdhFknn6j9n67ZMRo2CU/lL4iKTV+DcIm+i2xbwV4uIQwrEo6PF5geRg+
TffNb5xxkNog7W4vBFvMS1+9yGDsQM9FEj8Bk5YWKA8B/qdRU58w17lntPYc0YU5
S8+5tLcXS7I9BpIbSw4srA6YnJJXWv1jaNRaAtIxpl65Q+qcWzNJGCuYtZlIzFCP
8z/mtr+TMeRnWNytvdIFVE0OQmZneQxWDXL3DD9ZECFmPo6wDTbno8tS1iRUyrB4
YKcMp1lzytuU6EHkvdI6ovDWRIs7IgSFJKMKnVaZuh6TJ3NZ7pSCEB9VYTylW2Id
9rkYCy2VUcBtVc/2FL5sJpK/8KDKIeHssqMITWBkE6Ab2N5t8Zeki4z3Xu/FpUKW
ClGD3AX6w9hDXp2+GEtqwSEeuIUjioAmmMSRn34Zsfz1Xe5dV1hoeg7LuvTKaon2
nAKui2jV1oGkmb+b9MK1QbwkyQ638f7JPrEsWPoBz5OAlt1NBD+eiMPPp9KEw/Si
s3DnaAcT71G/SfZFaq7nscyoi9lim13a9ONsO08O8oFLs00brg9zMg3DFfeP0Ttt
6cxdeI87vX9AjY0EV8fuDmasgGegnUoFEnXVtAjBekzZOFV0sDw2TDBzY6yXqKvW
OwFju6AOyJBH8OAf63v7CWlgK2Tx3XRzHBiEAwVONpKqSX/GLa1sRn22nyyBohh5
2BVJzMfzv9yMFSuwIb9euvHc9YZa3sCKZZy1jdiK7Wj6rbvYpJu0hSf+sbrwrbx5
ZWhPZzWIfktx0HDWVJxDGUZyZOEywAzlOCixF1QTu+5xDAW2gzqePbLLFHqOEVyw
QUnIFRQPKUNkuDFiEJnLMLXTKR0aPEHGZQNI2HQsY6Jk9BqE/9s8FWmLdxrWW4A4
Y10Jcpn4uUcF8jZ6PaYcmN9zhr2I7HSf0e7krnbIXI1Xp1P90HNJ0Ds0NuIqCPsf
J4FTyVPEpZlXZeVMlEWDbqu//yJjJAxqRiLxHF+tcSIhOcbV9yuJnrG74H+cmQEu
T1nkmOKdZzdNLHB7KN/mHgnPj3QzEtsK6HYgX2tfn6kJ0K5RRqaf0/DMp0Bgu7Bv
hyrMefp+xhJ1izibrlRdjZSgX17FkLge0PI7MSYd91oAfMp7V65g7GLBACSQ9ymT
RdYX9nrRGdZqAwJc3/H0RapXDUQGAvYHhhrRltIaXkLDbsGQOAtcsraIQg3T/cxP
qiznTVybHNzOkyALnydWy4PBHA1CQwF328kvoCpbc/uP9ZNI/7lt4LlQcY3C8Ja/
QlKdXlXCWiuqML2FWFDDzfncPQbj+3cOPYNKdAIb3oDmiwrt2QGxyf+0RmrnG0Up
Fl01hgpJj3wb6ZVA5JwKSl2LJPVuW0sAe3TdeGFmJtEYYHRnK7Kum1UBS5czDYaI
yTqyQ76nhotY+KPrdPb7mf+sr73pzqngovBznbj0IET4xV5XEg8WJDc46t4HUCJj
4kvzk5n3dUxavvbjtHifaa45zClIom6uHOWPqqk2JFcDzXZR+0piHBFL/Ht3mlWS
/Sy7pFhDMTm0haYXFgAcE2ewRN9JIgNFooCLn2v46u++do07EOqtvU13Pwiu4fJB
ERuXJWoj0WUJLr9THX7rAPC+qhFC2eIgajsJHdWc/61XbY47gO6xhK375g/v9WHz
EbEEEcz5EsH+PMFMgQptSLLPNVgUYYNLDDg+S39e7L/kCr41T7YDx8QsAU3m2wCV
w9i2skmFp6BZjTbsii9eA9l2XB6ueD5iV5dJ9nujZRh41GIcjCa9OY5S2dKIllRY
2dCxFCp19Q4qOA0Lxv19UErB0kzdRqm0CB3HMn3PRD0RBiHdUCLdqFFsYtm62jAK
lS+pSP6klmasps1amZ3Lof7BAFf/xTLIJ07/6ow1USlcPEPRqrov239mkZ68ZPHx
se5k6xZfk3nQ2ot0TbYCqqA+50J50FtsjnMWl501sCmZmVGo8eP9jt8H7QgGCp8w
FSryRbkQkWiv8OjolUXF6spKLIW228rq+dVpDEojoXxB2V5uh6Vkf6OyBdUFn1P6
nsBY2BnwL+JKLfZmkLsOGMhIM7xIsgKuf/nRrnYtQTmqMflIaCdZlGBtVPyeqUIH
t6p5o9RmyvcOAbBTt+IRMOoqI+tgMNJDSYNvEy7HgtE06x+YPHN40WG4i+qvVcv2
4BnhOtl4o1/LBSlaFBtiX1MDKmJOPajiKWf2H8dfhdAs9/h4xkRCcsOoEkcIAQ6l
8/yhSLtpohaHUvU20/GPdD/Kcx+0Lx/uYVvSSq0xsm9hC3LXtR4jnuFjD4DAtr80
LRUVeDgoYsy8bGFGNRf33ZYnujRrG4KIsi4Sh3UpTsAmX76T44ZMQxjy9nCiOiSi
YVVgI1qR4yNBuvgFWIe1E7GsuNwvWgZaALEYd/orCrT5fJYn74J5Dl49sYEsmn7h
NS3C14U4A5kFqsTL+80rFdLF/HzNugqz1SU/87i6YJzqA6Ybqxp28Mfci+lqS2i0
Tb/3efteTvpxwvIpb+65tyn4URe1SRAVpOudgRhMQF//g7A9LIvLgwdSPrtGajKm
8CVBqWqjQuTi+EIl5TRlYJM1EYen62Q2C3Em+yZJsA62s66GfivK86R527dZCjK8
7JziYaVC9Myafh2hhte4PCpYWc0ZzG3irqFWBL73vM4Hqmzi4+1PblA/d/SVGsL/
TcJTtj5GWbUwJfz/7dbLsl5mqMWOolYz1R9iNv1132cEsGxr0QS2Sq5KFSxr4fhV
91oTv0tf0zl9sHTkRfhNJAkXFEDx3JMJrFufS5PT8af80LqTDNKV3+AF+X9AhbeJ
M6m2i4LqB1qPMnh7UdCflaNa/KFrrdpgTq2PXI6tCU3csZeXfTLp8bgdxRXOKgcK
19sSjUu+lpRmWTR8ZKBqPRqeFFS19JzpEjVaZfRXlK/2/9aj2/7XRX5AoTf/7rKL
bHWMDd0OwdIuk9QHwWHU8uZSa3e4/LbrIESj6canlgswwYWn9jmva29n80HkMpvr
CVsdWB19ahf1E9EnIZEY0blThyxskZjeId1oElZ+Sg4lT7L9pz1yKHookTx2+99B
jVPL6YLx38zH1vMd5S+CL4cZN81/ZifMkzuSxdYID9FZL3VnPwv4EUTyteGj3h4N
LyzpLQz1F42pLMoHQhOVQZyNU1fjNjobX0pam5CB+ugG8901WKT9mNqMJZiJelOd
aHhLRyiGC22faCE/xdMtZitoIetGMgLuH1SY3v6Wo+tQF/G+HAc2G61QHSzDPHVz
ymJ49DH5IolUD/zoYL6QlBmjm8iVUM0JZMkYvFFRtxCp4SZ2cpq2hFMdK4UkJdUk
wZPU8C2HxUEXyV4wRynyPbGKi0twDbabx8ELojihTRhJJ281qIDhI/NVuGw9ugoj
KvZi+G5ETvLXtY4/1IYx13bd85VZHf/VJ9F1Monwh04AZ79PhwMW0u4Mrq2oEagS
CqGQ2GV/ywv8OySLdUak5EkjJVvOL+4DQRFqDTCUdF3/sLD5KUTna13xNaRhQKwM
hVa+grAXHrzGFdKZmfNullvd81eoEiPXSezP9oWa8VwjgpMdsUxEAsutfWppQkWm
Hsg+S2/5rdICFgBZ2ddNUPzOYMpczKnDTEtxbOooPmMGTWEgtOqGTjqDv9yD+TEd
nAnrCb2CXs/hknaJoeGumYZO0dALtZFTSTM68X6M6mJ6gz1hXoHh4aXy3ube8YJF
hYFWEZNIy23Jzy+gyEpNagXlejqOkyqfk+xODuNTT4QouVhvtajOcy8iA7O3JNa9
PuIZb+NUaz1MJ2x0wVr6hPLnw3ub+cRNFIsEJVbnvkCUz4ZldPHUhZ+8GNSRupRw
S+hYxmROVDPsv/O2aq4L9gGzNg7KKv9fzwsk4FbNyRlKFB8+5YmU5DAY62MrwL+v
g1xYJTHgoXvQxW9fhcw09hiWkUQhhXSvxPfjknoqTnvIKtG9hEZRhctA6yMLZewf
6+RKq6oo/ZnZTxj74uAPmD0y8Pe7N6OBIa0tGXd7NWUE/vpZnFtiR/KbTffGFW7+
kxYc6m+oEzcg912tRABy4q5Hfwpu1RH8IX0F6rY2ilefwdO5bcOxJKE/YJiV/nb3
oRh8qQY7HPZrnL51w5zbskol6kyHylGkeRHDws5BWjvxdD/Q1vTIS5TLAk8MNi6V
2p/7WIzwOp2YRd8zweOm/lbZHMgOEVlQIAfxV2U7PENLjwTLUI0yALczBvFNn5HE
AwZ+wMz/3hTDySPBT7vPh8DXZfCMez9NhGr1AXfpJ+WZPdHwVhXI01+9cuJmv5Ox
I1WzvWzmbxX92EzqPyEr53dhqOB+k/azi5mDBbPJOvtqDiPSAgVe30i3Bj0Ny9+c
RyWXIgQ4i80MEUg0hX3yqULIM/gYpIUheY4ShH5GvdxuQSBkjNISaPLb1TDRe2c0
BnEiMegeUmS1NXGRZmjUQjrUpeTOCnRt/YUt+pwmnM03L9zT0X++Pm7cKW77+vKB
2mtYWxI5sOm1MGDQHR4Qc1DrtFAB2Ywtzzd5rE3xXxYt/oHqnJIwDUSJ/oPPkU0L
V9pBb7C/RixglApUlG2IEsCsj5ujUo4yES+Lz9Cxh+8dZ/Qp9EpQ0q+ZA8ewjkKi
KrXWPIzj9kikQc2N5U6xwwPEuxxG7aDQzxiNtSqlCeo7sJxZPHNly8ts1/ha3N+H
ENwGCbysw+oW8y8ZyCpskO/T2n3obeuvGnYR7ObtJ+GptxE9Dxvfqkwf63TgYhzl
JkmZclOoh2Re24MNBG8K3sIKg5KjwLXKTdAzOtdS/sAvZrXMSoGpDSr1uI6tgxEi
O+Tt3WzhEl8bf6m52zgdfQ3kJF+k8ACOcECDjoa7mjQg24SOdOnhwNPA/kdRb4FM
FCHcvCDVdWLbpVp83BFq1attw26OGl2ulfO505jlqgAv7UcHKWxmW+dJNhYv9Q3r
Uu7OkwBiYKMSTx3TLKmqgtkl3NsCqt3EfyEwwOnS5vCimyGpVLKy2wxKf0JRZx/R
xnuXvWWtn5WAOJ5KEmYYRjb/kpebp2KUMbws7N+mN49UTx1VF3H0n3w50X3mWifH
u9q5ieCM6ukXnYfEYVeKQsIJXF9TaxM2biXS0kBiFun8MZ702fm05jVRqg5XRLv8
VqYaCYoa10eOj46kkRgIIH9igaUY+prVry6ZRJkbMUmrU0vAJdr2GrWJlVIpQfxE
n6EriDZT0ySI9lkozyW0CGOhWqZj3xKETFiKII641vFZiBwnXXkWuUBTO5TQGQQ/
jlJtPmvuhJSW4vhaT8EWHVbOJd3Mn9VWfTDb2iSagQC7in8PX8ukTSjtyzk0mZyl
qaQwWl4m5Zd7tKDAmsjMDhBxOwx1neZpIVcxWVZN/5eHcmhs/mE5+2B7XBXxsdrK
dU3dFUYwoGeFgB7HwxjJ+saa9DlG08Gl3DEmb6fS1zrkYLZplKdnNYVQOCSKqH7T
sW9HlqsgFPVcIDm+uDJBjoF3oMrc2C8+bYeb/z9GEoF7wwV+/hAIFIF6Wwet71zd
F2KNa6J3ba7t4wPmcwos2DVE5ZDUwArIpvCTFk61bHM8pfCmFv6wsXQK/0ci4+VI
4zott+auzzzqwRjjJKmIN2zMVF6UBvaCt3AZ1p8cFQodXVrriNxeUzbPOFk/g/oo
GwcTUGB1ORLIT3rwYnXLAnjD6/g1ytLhpOf0RV7USg8mk/CIHsri9/eOdWxhKvYj
Bo8pGxpjqjZGl/Uh0MhuxKqKy+1N2nyUynhMTk8BwdhpnUEwlZNUAR6zTv3kMM6A
JmZveiWLXd47RnNz+aYC7mOlsu87VFngHhnj8Ph93ytPorgzDZxAed8Nu5jvVSwH
Tp2tavXVNLYRYCUGJOj38D7umJXr85O+ktiG87ETeaRMq2g+X/LE7iSkM2oL+Kjn
6DUgITO9pMQUrvrsd7PQrTDfOILHJLXu6D/PueLOHYKZKo7viRhhWCasXNw19YVw
h8ScF+kyCk4V0+fv7DHuR6b/KUmWt6EU91U6+r8I+Vl8LA7noaORkVGFiAT8Nj2A
3NnWW6TXPKV0XIGtejL+Z2vjdxidV+wz5wxjwGPvnTtHCfKcdcoQB6GS1OLtiNQ0
8/d8BoIDZiogid07l2ReY/pFXhFpV9JsuTm/hJ+elfzkreCoRqZooNUKf0XwTk+k
Yat19/J/PGs74LyjQ17YXT6cgL21oBelz3nf2u1eyMrAZ0KyFchAlAFK5huF0h+b
MB8G8IMOyFrp9HLJIIxNdshI4TEFoHuCrpX80FTojnhyGk58gY3SkmE+ENZZ/XKF
gFQwhewnEcaMeZgv7RIgMDlO4i8fN1bbp5mgg1bI5X5roUos7rxVE+qtSQqbbJQ6
iEGK0XTbkAyDH8gvKVE/u0ez2SEt0D95vp/Ma4TEluUFm+CllUVi/HnBytWT29yK
SgUW8tpabaR61umFHcZKxr62LoOB2l9+N5vOAJJfRxh2V3ZmoYKZ2SixgdDQ/Qip
QxmmOu2nRT1ONVaceE5/9pF1O3Prc6zELk7r+49s46ziIDNXqdlG6mBQf0yPcQjw
Scq+c4CRG1yec2PPvtjwIK2+kdqheMcwVE6d8zfVdw1qEccDKF23EaUn0Zz+1nIq
SDMggvKfrV+0HAgur5d/iOlweBG+szd0gjT7+wZs0I38WXYWuwplPfUt9pgaFFpw
zUFJb/dMX7zyKhPMxeytvZKeYj5+ArH1p/XtWUi9drechkbMuXO4f61ssMYs9ujq
uzim59cm2DOeTIts4G+Jevas1Rvz5WKOUnJZQBrYeG1bBn2+moY3YZP4SrE4l/QN
hALH07R9wA7kEWGux6yR1e1trdFyl2cLlj1Ob3ZBDe3iqRWyPst81bMXNzv+iJ7S
4+6zQT26x8r9UPyijYG+y8Ev2k2XTclsuywUf9mAqfEMJ9GKVI9W5HvmBbmZR420
+67rQCM48ofTVsGmToKLz/0B89++kFnmJyZxeEiNXKunHUPB4eSizVwES7wew15T
ySj+LG69ORUWChzTffChN+D5GMbzQ4yT85JNYmD6O7ZnqOppLv2jxgGvbzCowINC
LpUOR0gQl+TWUaaG78B1QMMbpAfdM+jGTf8k8iRWEAA4HnoniGtaECJJsZsFW31O
qVR4pFFi9tnBoALBN5dcgZjjbDxXx5C8iNxDnYwEHrpf6lM9vPgKBgixPhpWJYV8
uquXecGPPvYJarAqQPZo6L/z7MCFqkjGGWXOsXDBJlwIl2bnsb9Q23jke/3yoHeg
YfDbRdQUkX2gbbqBoVl0lL3wZlxImvrt/mWA9cDhuutjJfBIPcTNkiUX7gMq0whb
xyVvDcuuvuFCXqEkCsTmnCaTec+ZAfniXTWEV4nGgfrQlLXmhNA23WOm771nwYY1
e1YydhlTTHHh5kokAyAiVhLP+vOMNqOCguxKYBWNWhuYGgVdU1Q6kgqU8Op2TpAn
l2wxM9ua3EG4fh1pXPTFFqYH2mXKYNFVL+j0UFcgcvJmLCVW4Q5lGu2BrZSd2ACw
aHboSSHE5SfOrO5yPEqU2dpl1XZRxOnuSClkNGDuQIMvGhnIIH8drEZEg6vbp5p3
Mj0bbsmZn+LxJM8kmJE3G3cKOONpnCbxG74/YWzMblcu3SvneN6SkmhwD95xsBU8
hYWNt7XEX9PoB5yCVpvtPqcx7H5J7/N7Ilz+7w36kglYWlnq5fsVCC3OV448bheM
gfMemD4SMaDUkGYKkpBgThs/9vdAh1bNeeSklKNJPZeaTgsnsvA6YqUXy7JNqW8/
r34KlX7D4gVt7FlxHmGy9TYAvWjBR0k7PG9KVVPyqvkagLYhQ8w6ZIlcvNQyBl9N
PFeEEqCqduxDskmwIlJNmyTkPuHyNO8WJU0DtSpCa8z+zP6KvPE9re+eveGCu22Q
Q75y0OM+fY7PehQFwtB84rNaIyVEjBMUKZHLWfwI8f0k667H71vkq85fp7RYtnbf
kNMQTisPgrDUPv4q3ZelFpEVxc7OCzPqnX5xljVZY/2ghMpwbFsiG9NqX8lzXGta
wijvfZDaxPtoF7ARk+sdCsxqFs6Dj/qFkgKr4FryEFtPoK7sNRXC1vVvwMYOugCe
E8TP666GdDwv0/acDlVpOwhaUIwNrztevFEyugDl/ECqZvaxzjkYsqbX/ovealcl
gKWwlw2BDjB4gcU84hEZydD5HUJSzZJ1Un26Z0DkUALOt4RUlSLjlO4S5rplwrLV
pmAXpztxqWO5P4Xontg5KmRxWf6tL5KiQ2I/KjxVMdt8mIJQHLJ/o5ftJusl2yQK
F4/1wtxKGCKLBIcmLPUmyND8fu5OmIbBIiByd8FBYM6UOHlppt4RMeVKHNaI+Kd+
OFSKF+rBmrjSqA8BSxrfP/PUNncX7DADQNymy8MShFFgSyXr+9LehkGfwoPe4ECg
X8p16cTeHZ+WoyMYPFGyccl8W9Dpy/LbvD54UK7z4kQpbPcmc42E4vBeIFcLZF0J
cQ4LN985GYt5oBpIdHO/OLuGNod7UFwjhWqi/L/xrDOwfr8ay3rtA6DctLfdm59W
BUwFs8UkD0OA0INrep65MrRYJvSniszKDlM95CSN3/soLWSiZ+DtKNxIdjqgHxTU
L67WCEdFmC6g68MZIgiAzCpygSEHwgXX7/4YKmBFWH9nqHFvwv/klwbWo913HpV/
Xc8omBKASaL5efUb36D0vwBlGX5LffNS6G3ZFbbQjBiqIcT+y1J+bCus60O4IVlh
7n84Vd4F5YT1W8nOtHsXr50Vj/4gpkDAuhUX7+fEBt9rxnYxdcXFWzGRf2hq2auC
BEwU3yWnu+55H2L+oZfxBUmQuNbx5L3AP23XsYlNbdieMU1CGLXaVK7X0sawdJpF
TB8LFYk6yCUNeizrEs3xQ3gi4mxQFyWpxBNSKtf5yrVavOQCzvQB05X0ZWbkHDDc
agpDPg1A6tR2Rd5X+USILHVT3jA/4Z03H6xNjhcRPQFBStnHFb611x5iMeD+Fg+Y
NVZS4KfbjaCoF4hh8kvpRm5B0n4Nv++l312wkQSQqarkwgeW9LMEFJiwByaxUNqh
0S5CgS4XuI1ysIXVwpIYNzeGGAfu41yUcW9YxFnji6Fd/3LJOgoZCKtdd9ICUg60
bUHS42GTkc70u+O3j3iLPUAoPjmguaYE4a9VPKhb4qV9WUedtQkZZAxACR9Hmmo2
sXMhar3XBQuELURKFzrDSW8C9xItswhhGb4SJikvV51jO/Gf0uc6emC6jWm/zTlx
YrbfZK1KWW85j7DZOa4zCIF1DwDRIywdH8jzMhNQX+izQ+n0hUn92V65MFklx1f/
D733udC2pScvOF09rXxuQtVcnlVGbLnljQJVKSXYtvsZdmVwqBsE85aA/fcibDp6
3NCzqSYd7a88f3GakKYvN+P9tTq5lc3iVxMlWZXJiDf9kyfQZd0xpSfZE9qVo9Sf
DzWJRHOHGhauh3qA7zOQGrzVKGf+Nz8wfwkG6NAChmAgGGdGS9w9k0oUDzFR19n2
RMoOddu3e2BpDXz8F+iJk4G00vF5tIKy7i7Okl6e7PY4TFbMR+/K9qxrGXGN2QsY
E43ouxpxQVjgNH8qxEyolhSgjGfjK5mPhoiIjUMVxZQMSeKqjyBLAKP6D0LweLLl
9znRNHTzfz8U+h93K5hHasqBuKOF9xOXCSewjJnBlzpyxfSRruQZqaOCjDurcIM3
Mb/notLFRBpW7yHx0/mOa6y4srcL5UMszIQqKlWXbw4Vq4sF+l/rZ59MrALsGYR2
64R75HBJSy92UiZsAvmktsib7EQUn+ek6/aKgUFi7vmcSgQzKovnh2CFlVDAg8UW
3GZHx6HtPsSZRWf2IwxqtbwSwu/z/2TqGKXCmJwdXUi2HjIjV8XalQuvx9ZxJO7h
R7qyGbqeSJRMRne6i/s3DYnYEhSMccqx8mQJS5kpFdqKphmOMjNerOFRVE07WxgV
TP7G6pWuPKHL0yKzAfYe7/MOEbF55GTiDj9JrzRa9xyWXpcimd8ViePXHS3p9uyN
NzA85mLu+ojzoFfTEHatV3Mz2knI91/6PwuwAZ3HrJmSsHZ7+c3d7HWN8MRtep82
9JTXWs03pC1RxjB7dCJzGf9Vv9WbtZkvAtmoGv7vCHp36U4yUn2ggYr8r2p4Qt67
5wOA1RVIklIl3xEtltf2dCsiBeJiUcnQcg5K9aOJPYhhCcpziu4lD36XHdtsF6Qg
lH/GEl5Ro5SVhIn2nauKEoneJhEh+zx1v5duuVRibZWv3uAq4VCuu4JGT3L5qA9r
s/bTb+j/Vzep7QfYL+hDtMvfRDmDaz388XfQKWxlNVQnK5XvPN/p53rj8WDdXjpM
I7s3LXjfYt2V8GnhEeC1X67rTDW5fNg2srNWLZRahvpF8I4VpwGX3QbWc6/GZ67B
RYgi2gslhp3WIvjVDaGIz/coFWjNnYBv8Sxcy88u/r/qEotnP5b7kFVHjwFOwmIO
0s8onmgN2TvX8nhT7fKf8e8QgpzHUCG+4o8GpirK7IPVfBYLXKZmkrsyy0pleue+
pCDZFW8SS35rnJTJStKQJbeqJHM5AmKMJTrqQLaTOaMtr3/XQ/DtfwCxvO4QISMN
GJNUj9aE6eofXwsNfwDHHT5r52Uw2VfRGvWF/tnvDQE12KcSl2KrFaqmPBT23fCN
QVE40fXQ7oqC4xag5YP+qLeugbkQw/Pi4lfiq7M5r3EaCLCXyzXcSySioj8KVR7I
sUXuxmo7NHVVYfaABDrJPe7o5HwVgiwHweQ8h+rE9UKSBrPrmjyeptspIzP/pLNP
QmV6zqFEaG6dPYHlPfESKxbXXiijoiTg4lni5CAqht1VDcFTzc0vTocFY7fHsoUt
T89vkcbjmpzokwyT2EIuRYDd20hl2EvP6ijOi0WIKcgcO9TUkl1xQutfx1hS1Ggn
mjzc6a+zh91OcBmIz8myRxod7JYjsOt2EWtWXj5PC17iQNevJXNZbnxhb8u8yGRw
jjGK2eS4dP72vPFGIan/QMuOlwQgtPNYGs0wLpWWmXodrc7rQDxJSv6tKS7kZps3
No8vCd3t+sbp8KHhUZY2d3X9R48EqMW1CMWkZfpDZHELsR+DozjRM36UkzPITIih
L1joov2F+crbH6KuPBADmbucVpVY1koFCvgbsS0+mkcmsDsJLxq8m+/uNaIybOYq
0RaVNaqoifSPzJ+BYSxpYLX4uG5U70lJq/6z6hTIWKfFUp2ZpLpW0VwfbZ9mRpU+
4xtMXXduTuG84pT6YUsrn0gHL+2qat6gPFtWrvzmARBxVaGyzK4r2GE9aM/Y6KCl
I313NmDjT5NS4QhGw8BwtM+axcfdT8tVjJiaX+F8n9vTjmAZ2VxkhxfCWNvVd5BU
odeu3GZwu7W/IWhksG/S/8WGqny9uG0CBGZHflHFdFRFZux1CgPmEFFg0rV6PbhG
wimvHu44yOQnHF06ZTsvYRL/v+4LL/8zqlRHodWdGZbVm1CCxH9QpKmprzATSGpw
ask8hTZeSpNw9yRwUwAMf2TzDEc5/qftIshpkYTyib2zVGXlnyCKPSyjPVug/djS
y2MpyhA24m+UsuTEb+ei8hwn789iVDXtxvZAzwyfANSsp4lMo2YPlZ30Z39dXJDg
nR7M4u3IdeDpZUx/YC5di5Rhr4AwfMH9nt4JJxJzBKU7MVNMJ0ByfkdTKGx0BVnE
o/SaBUux/HphArC3jSi9zoitGWfAaZHSh7+IVTAaH6cMvPY1UQtwX1TAb5HDJgSi
0KF5lRvs38cCyXPH5GWV/++DhvqWl/RkYxKN509cNzekUfnxj8pOORoh9VrX3JGZ
sPFhIoMMqiYlFdtVNR/ORk5py6hR2nrPVcIW0belJlg0cWsxQmHoBsg3OrKGl9cQ
0tXsjzOPe/LrzzvU3eMoeRoCPV5pN+6EW6AhpWvmDstlcjOnktqaXzHDsYexwXxd
ldXBe0Y15sdWHcwphiMSlYW9nwhfFDwR2h+ytV5FN2BCZyAMUbnqNNilUoEx/VEq
1HSW1nZAgwsuTCXvcFJmYiba6Fk+KyVlWRKUBs64aSMhzOAV39Ai5WaVQS2LJqQn
U9+EKTy0fLoTWbr0n/r2/SkkCt7CLyDUlyBHs/PFdepTs7Yl/bnX5uZvub5akIpE
J13+6UjJulFIef0OkTcYTfQGB6U4CVPYWDPutJyks6WLtFJoHHHQDrmdIn8X3BY6
kQcGjRQFsZY4adxQ+TjfBKIiv2aKbSZ/V9CoRohXlCj+oSgezZUMRZsJUMucu2nv
1QF/TJpL8M2io6XvFI+rm08Lki3ywMBwjFcX+w5A7fKC+7MkwoJYo1C7gnE4eBfe
5YQIA6Wat3u74EAdE11NUEK4ZaY03sYn2K9FBSVszqHwE435q3jseAKI9+xmTFQR
LXz6uG/6D4XNNQpM0rfYoFwDnrcGG+OpX6GaSISAPrXPU0ANQSbjMLKm9crw+7on
GFHPjitBNmVzKTbYg6DcxEBDDf7cqomDChW6rpVB2fAELtpUG/s+ovmyh9gN/DMi
8qP2aCdHp66d/03bRJ3KY7qT7P9Slba8KU4x3MJ4I/tRZivXlQII+eCCDJQoZmrW
X1sEkhRwsbsTJrtmac/JRddyxFih1yLzWdS8+8zAtbotgBz1IWN34szdakeiyGXb
nOKyzgxtUISypViYAP6uWhnJFGU1VZqVwhFdf63bi7VqSj5brgjEV7V9o30bRkOQ
ZxWmmpRO6uC8KXkoY8dteJU/LgrFg9Hg9ZlleICy6SuY1Q/ik6UqtscbRJ5fOPwG
qjfzGgZzkCi60GiqXKQXAMm7q0804mPI4ZAUNal58kUNHkoa4Ek6tvgCxDGL+w6N
039Nw+tQSG8vZHGTHiEGRdfGXyKOwtDo7oWLkNk7aQMvfqv2RofyuOAkUziQ8Mpb
JWOSy2Hp1zwXgwzUCTy002e/9/BSNGx9LLyogK+WIxyomdJbV+vXuNu9VBnU1Puf
810MILhSexFXKWAcJxE7xJDBM3HXHKF4sVg+UiTvXdd1cd9AtkSwlJijdHvb3ra3
nwSEbbNP2lYFH4e0jkzWkhKJMhKi9LN2lNLUkg7HHecLO3/PmrIY7+lGE8x2GK50
mdpon0n+54bceFbbefFpejpnb1kod/C802G7N+scDaDx3/HE2lf1gbd0XW0gDW60
u5elr/vt1h42go7bCXx0A7njybFcnZAtqmkW2+WdrlFP+ne7TidxHn2kMWfSs/6v
7jcPm5mWBKNuIsaFmgH/m8c9kTYMYlDZU+ezL5Ff1orLiPFGi1ofO5QIcwQh1Au1
wfKCDMHh+MznUhtABDKMthlR5gJ5MX4MpPnoGiqPznq6onzNvJknX+SkAtabXTGu
dNuz+Z68WWVKvzliYgCapnRPPkQJ21Xy31BKpyq/wqXnMNc488W4oa2k4ro0toak
bxit+GVV/klOA+prNTl28T3GQo6OhF9tXL4mwTDOIdlckpz70OyY29PIAwK/YlGY
Zqtjrq5/DV4PdfdLGA9+W1txQZPnAXPahvQFfHWd88rnNovP9S0e52BEfgjqaA1R
bK4Jjh+VJhRd3/bYeCYutFw6omiJYEd4960E179YBO2PgEIqFDkrAcHzOVJ4iKeO
6TeblI4R3OJ+BPy7fM96NvUDZ3HP6qs+1Zr2ZTbLJruM2z2GOP3lE0McBPaLNAFM
fNBHuyxoJteGPrOfFrH+uDvGsy7D0R382fkBAHPEGtnhAZXseFBmFDavMcMxn3FE
CDifX8iVMRpSg21CT/VxmEBmcBFrrqcGszDkv6ThkEubV1t7P5NdwQC9v47QSkqH
ipB2+Nz7c95X4+6i22/TcfGC8jaCCHVcPAo1zJyMRL//S3CmKKiNvcTISSY37aqY
5bz71VHJS9T0FZi5Q8KXESXoR1d5KIuHt0QjMABzM24FlWgi0YxNcNUi8LpO62fs
RU7hJArXW/ptr3LRYO9mYixngTh9Cs0beZoDOe1tHpRBSXGe/JX4OOeLuUnCB/QZ
9tvudFLj+yZK4PI92m1+Db4lYNDsbHlc/nkoHmXEis82sXEv1Qx3F2ndaFiiCxnh
bz2QoS4C6jtQNBEhqVNyWpAdHtCnAz54lgB8AuHe3pr10CBbP9pXoT8+y0y7fb4S
bqjX87HM4qCezGh4AkI8uHNwNY0uhaj6+BT4B91wogSlE8jOtw9m9h3ge5gbuG8G
XvIIDO0JaQR+PWxhVc0dVezl552s7aMU8NAVdzsD5uEXltbnFsSFRPLkg7TO1gpV
XSX1s6GTnZpyxwOFJ0yoCPXm47dZZhkB15atZ2p3mBTl1et1+1N9VpitcbPVRNDj
HaZCzS+7HmGhz7CKWZgorIzyZG3MF3E1WuWE0l5jl3vTKDXe8pwy7AteZYpKed31
vvLoXbzWAcKZVORBux8vzPDm9aFRghnmxthLHR4ltplo2qDRpzjP+xkD8Npud7fy
j4I6/LrvAeTPCsu2+22mQtskb/bAf+HUXkFe2Sjo4fVb4OckdOayRvxJD6lnJa3E
KrfqadxlvARoriZ+/j5N4lh2Q9n3ce6JwQZO9kFL7SkgatcehaWMCr3Zj2Rb1BVh
COLFBujHDDOJpn/M07BCNEk6IVgsltmv8wIS7yq2p9svPxvN+CwOs/SAtdiLKgu6
OE0t6rnq624csXLGHheniDJ/Hp/nzFfZRaPPxDUlM4eN4W8gQYSq2TvM9CKiQzNx
4BRHgiGyjU777elPH9x71MkUcfaAMQhj9LbWYtiClVX2Mjuhh3IGdp/xCIjGDl9J
rJXQZAxOqleh1n8bywT2mTLIOPZDXAiasjv1S71/YehbqmNqW98zY/WrfgxRjcey
193JU5zlH6QTQfYKqtTSXaBRxlUg/BkGlz5P7dYjSBdh0hGN+GR4cdFv2dbDE1Yu
WKW8do6EcachNQjcbnNIa1o/1u6V55/rmP2AkkhQJ3WFR+lhJOJFao72W44yW8+k
FLa68skSy9/80uJKphj2v7x6v0fW9+IlvCotOe0pWaSCclceRKDDT6/y7NLlrmN4
41Yfz14oalYB2cziooMif8r5VjovyindL53qCkcLRK1/jFvzor/njPbkve4KWCZL
mu88dtgTrQYHDBkc1m3xWnj6sTrF+evhuun3nWJ2mT1wBKa9BF9qaBU8IHrpPEJv
QUVR+XkpJ1AUx/zZuGvMOc4oz9wfn9+oWAFEUjKI40bhsZlIhg+Z6LVH/gNwcV35
rR8EVpYdryCrtAzNwJd3AtZP0zFGasUUb4UhsRXhjSfW0vVz47dqkqoi+awPBvic
FBmyxVvFE7A3PQQMTGIAdcovEyc2L7ppzHBODZ8DZB9NgRuDT1nn8+Tfs/ZyyQoS
ZPvsm/mlL8ifsUmFCqeeAkosa1zRr39prWLr8kTVY3aPTNXIIT7nk1IPmOzJz4WK
j0HM3wWRUmk94gaEW6jXkipXxLlfYuEbbU2RxgAc1FthGx8YN/rKsNmR1r0/X1WZ
BJ32QnYK0P05AIC/P7ET5jQunXRJlfWPC9Q06e6sOysuTaDy1DrbZ9PL+KkZ4c4U
ZEIJNYpvPMFkuRc+McfslylqBpPF1OFMxqcQ7K+eTYtqcuL2Cc09MF4+7SSo9ANY
rpQAAHBvesOM22MQyplLvFlMVsdQxOSYiZS632qhTNTHc5cvUMFeWsH5M3/QuDwt
APqGrDMKnIt/UdXBMLDDV2+g1rafdvuqs7SARxCvCDm2UZmcQlppLIab3Q6GVrJ9
pe90v5jl4u4hzoak4R9QCWQBVFen2nOGMs2g3Cwk4RTTWKC3II3ymRoEt1XzWxHv
D+RzWCGcGl/KJMORZvyzUSnl0dkfco664cM1TxGQ4dIcBmwYKxs3b6yV/aTXyqhP
l+Efr6Z1FacNF4+4zZU9SBvwAJRbvZwrT2KhurUqKWXCmjuNKm0BhFRC/TQxkK29
ZYCQuVjFhqTxf8cy2cF2lC7VRbWLUE8N2rNQXsDSLulqN7r8Sy0Kmbw4JfeA325J
mTi7hQXm0MQOge44GgTaWByrFZoNc4+wMj9dJaaI1pu1ldYduO5HiPLT8rSJ66si
0YEaWuFsxCI6LA2GWpzjjKYLDTv6E1uk2oKd6cWOQpOyplSljMjXkgjmhdu2IjhG
j0tnQ/tKsrkisM8tDiuVN7DDo1iCG1Zc3KV37DT9sl/HSZrq2s1AUY6Mg1OfXkHr
h6zNwuJ3KOaTkjKUKCWiHQI8wzafhasX9ywuYG+jlg9uh5TzEIAzrcsPyNQM4kEY
L8FbuNlh9/hzfKv1QO3OAYlmTK0P8lYJ90uSWsvo/VdblMyQUnFsfuU29uezas5Y
bae5TF7BNtU/M+VWSDbc1834QNMD7ENmnfWBhpLzx97TlNxaIQEIBSo7X/GxKvEg
HS/xXeqZU/yv2fO3MMBqndTZhihXBb6NyTfCrPgmUTuSOMP0AgaqkvVUZuQ4g3y3
y+Gv3QQVrirgnzHOqQo+lQ3LKaSfy72EeNt6Q1OMRRI11KmlDuQTVY3M3WjOhvFK
O50TgUzCl+b5QX6c+qbY7nk0HjAx6tzPB6mjlzSS+Xfnz2jEfr7FJ3n8YXR0ODB+
wyaW+/BKhyJfeh/Rl/Lf3FrGi6Gx9axjTfeNlfc5GSutHrvJoHScGxJxad3d0/HC
E9EanCWHjG6xDx6G3QYV2SOS8TGmTDfMMvfn76U2SuKhusDbIpk0suGYAuBCI1ov
QzXgZRED2g9zl+0bCsgqOxqJxWzEo/WlW6r0GI3l6BYLcEMFSjCxc4aZ0TJ2IW6W
lcpzQ92Gm1bsazdgmUmrvvEp+qj5Z2M56IKaRk/clKFMJjODPh5kHH9uu76863Bb
yNWOoBAMzGFUL3OvuJEXUw==
//pragma protect end_data_block
//pragma protect digest_block
h6eAl/Wnqt9FVDIKjAiOAcCYcYY=
//pragma protect end_digest_block
//pragma protect end_protected


`ifdef SVT_AXI_QVN_ENABLE

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
nvoQeT827SYp9zXZNILl2aP6gfVPKQL6zS6o05eOY5ropG+iMGoY7nQVTBZYVpXs
JTi5hCHJEoLbhZV1b5FuoJBZ+fMI/+ACV6/0cv7m2yYHlU635SUrdK2iAquWf4Qb
mPAm7paCb9U0OoQt3HAqXnj1SYxnX32J3tAy7tapMe2OJq2qnCxr3w==
//pragma protect end_key_block
//pragma protect digest_block
+y7Nuk+tvm3aLToUiY3gsPYOwn0=
//pragma protect end_digest_block
//pragma protect data_block
spyUO6yVx1P1ks0XdCT/V/pueWQ2fJRaxi400cedtyy2Ux3PnIL2IZgWBjLucttB
fgGfamUtudoUzfOZpDoExwb8ICBWPxZD0+RTo3Bq/M6haJOeG6pqKnQRbeps+CF7
rWMOZ0Jz0RlMbUxa3qpp/pvMJp70rf2YhOaU+sRLphL3jjpLWOY/797Fs7hVOj1q
OAfVzSOI5jhbokE1OvFD8zUctH2hyTJbyVw5H75f+55h1VeN6gtN3FUgHu+QwLF4
I7kI6tAL3+iMZYu3BqmCHwLvl1z84cPP2rK13HfGx9rrILuBTdiql5c/4kfuU1jC
YFUJAH+sJk+i0i0Gx/XERiTKw/41V2aLxozk4u4VeW6zah6xhIL6Zusl9UBa2ObB
HtUXGHOH0HNJAOjCWZDbOfC9QEo4b6AR/yjceZ1GWIeF2j7vk76bkLBDprREyoDg
073wBZMHHGg9CTIJPuRclSErIsbeO9gSFrSK3lHX6WoFYuB6WcNb+JkiKFz5+Y46
ax76jyPNitr4dA1P8jiPQBRFeLUXJrPX4XggE2/bHkfMwIMhg3vE58Ggg/9sVqdu
WfyTyvKnOUH2h0v+zVbGdZRJ4IimEaAJqWLe5UgUakRFtsUGNiF+MxNlo6y1fYRv
CyHpRuTncI8rxsFY1Z4R4kBGhww/ppbf/3wPKNRQRmTMIlm7T0gfAZSqGMWy2XQG
9A8WgqT9Dj5++1LB21z5E3WBpxVNW7PhcjG1sEschySUCnsLy07FQBSU2ZwU3wit
G+0plfJHiY1mZ5ck4l8ZLfw9MRbklwBcqyU8ay+3z2zG+QyoMpfFe8CW+MP0YgOs
J+D60aKaNldDtGwLQF2yO46qjlat8dULdfIZZc6cPDcxlQsWB1zf3VtkRwL3EpIH
2Xbs5jCb1OkzvE3JDaDd43F/H5mb+zuL5Vwx3RuLcozv8Jw40YM96rKMd70iiPf3
Jc6kdsydkbDvbkjL645vPMMfxhOZQ07oG0G0gLk7BFSPxTR0kBtxS64KXA0nvZrE
yr9emx/uFRNQmyEKN/pfRkRvy59jNEHVcE73p8FADLlqmgWTt5LAWWWUZ4yv/NuN
nPODfVX89EvYnqIJd034+tL8sbNhDLrmo89ohoEb1yKCjMB69ex8T7XcBEEWu7kW
SHOJaDSTIUeY8xCvd7HUJ88E4zyEvEpZ+uN2ZoR2UDWpxVSo4UGJE0HU3sRmTRMM
aCuoUvY6WGhaReHlGBOjbFKKuLAswqjsGOTxGl2mvGggQ5TkWoX9osaM/NGpAe3t
3D2TaCG7a7xNpwY4jEVTLapBUnhWVxDtM5PkdJ4NQLDJEs7hYk46F+rKTK2luT2e
7h/pYOvZRgWNFvcLu1Jtcv7zmKlq6vmRJ/WyKR8GkKxKcFCsBiB1C7k6tpcgzCbL
398wbKe17Ji5FXxwqGkmoF1zLrQME883xET8s8gkACBPyi+6i9iaJGUeF/Ny90Y1
a/uTBfGhWWFC5SjkxhqEiaWFXrDD3A3H7fCOC8L0kIXhRhTvH3Geaeh4gXA3z0gW
PZ/oUiv8SPJwse64pjNwvCrapUzl0+5yG0/6M62iUD0nwDOA7sGytmSHvwgf4ELy
TxAud8wT8xyzfqwIznAelYAJn7v610KM2Ve0SaEimC1IzCOOZS6M6rOKVxyavukJ
nHH6lumAg/eBbwEC3ofYdzBlUOUr14YvfE99J9JeZlRypVjXUNG8XRhjJSjysA9f
lhbw/SgR4Fg+m7p4UbpAACZAxtw7Wp5LMKPOBSZ/nJNg2sWhuBJ5JgUxtOgdLc52
t/crNhg7kpJ9VBwcBn4/IFs+wdj47YYMzopWaTF1wW5UJ6i0/3VXzR0szSseW/9X
04jLhvluOENUmK3yDAZoT04KVek1N7k4rVNy7vWGp+6DrpqnKPUJi99fIecq2ns0
DBxd1MJ1bu+NIFc8v24TOCpW7G5RN52hjrIsygEcjdnms3Md+dhmX/OhTKgkR3WU
+5uXb7GWEp4aeWMQl/FfqoF168Pf/KJfKnEJP8QQhyjFS+8DQK7gp5l2ARdMGHxC
1sdfUeD8eaSFO9OBw1bbLCaNOtXhc2AlnKMvH5/NpYbJp7c7g0hi5BgMYaPQywuX
2wvpnoj7YDXyhSywzR/Yt2CCaPUFI6ped49mKdW9lj0etV5H6pW91a/EZOVyecEF
3u6mTTw6RhhIbos4FsduLENxE6uWzwawu+XNlsrSYrh7+xtgKp+Y+GaFYaj2km9r
qJw7JNRsJSEyfj+5ITTm7lDyLHoWxAtHW8GJ0llFTviDae6WopLuFpQuJucGW86y
g10aWjDaQPBCABviDnL57wm8ZboiX/YaSZpJOdWpluh7J1lIc4+NMPHoSNFlEWrg
Cl4AyrSzWUkNK7ajO/Wq3gDmwPE14D9Znxpa7C8PuHCCj9Gem3fbXNlCdWumy0JP
ldO7Djf/MYVVMc/ZAPZP+4jC3BW1Elzy1RMUzGXtQhQKARbRwBI5SOGg1i3peHYH
8bIFmpBaAihvI0vKR3CfXhFKqjdct+p2fJ44/ulW1ITlgjKlqmMoU5kYgbi1WghV
/vkR+eKB6EEubzv1f0XRjEM996g9CE+tRF4DnOnIKqgM0Br+LwS+y1WyvMxLdIeL
Lmcq/zwyXM/o+DvnTXlNfxkYKTMTnaU14ZTL/cxkF2YYTIeKq8Oru3HqbcazNBfy
kbD08j4IHGD3Fo6Jc5lXI4ebJw0VaDTN1RN/y8tmiAp+Zw7/Q0R6QS2w8r0L3ejo
QAn8tAg0hqx4MYjeWqhPveWhz2hM4jseYG25Gb/s3BJsyJMk2aMLPxrxzxxbDm3D
y9/03NsGeXwEJOoano0eMPqIMflQJIExtFuW2ZdIgr+6LDUdx5eumQ4OXSlWrXhZ
r9HFkttoX1yrFgLTJ+zbAUeq+v7o4rodq0bHD58FYMTI3jMv50VK7DYVypd+Vt/I

//pragma protect end_data_block
//pragma protect digest_block
ws6jIBaukwuZuQGEKOW+C1icdyE=
//pragma protect end_digest_block
//pragma protect end_protected

`endif
`endif

class svt_axi_checker extends svt_err_check;

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ZiNrOH9skEokci7OCnuQAT9PmKODF0tW2ETY7mJVvSR7c98qdZGp4V62EG3BVk74
3HPm4rNZch0aZSJJkozl4Za0CLZ+ZSwYaai8TVX9a7xHW41RmlRF9DcHYzaV+8Zv
eJzRj2wthrde+/vLwyITsjIHdbBtcmRXMFWxaqEKueY2zicEdRNmFg==
//pragma protect end_key_block
//pragma protect digest_block
mL9VGmlVh9VcjTOm151ocFB7Nq0=
//pragma protect end_digest_block
//pragma protect data_block
7LvNrYM3j8XZgxx2o0hdei6utBt815WbLlnEY+cHv124aPgZPPHzmIUEFhOV8WMz
UVcS4GF67cXHUiORPtR4yyKKIHnq8ucF0K7MllBEZjr8W12FZcFJ5BTLLPRLRCgf
L0wZy9laOAVVR80PcCWz2lbFxB6332NKPQ/9dlJlycrgrwl9nCbFnUjcdBzqyE4j
fBz4/xF2T6fKbKFnrWm1crCxt2x6vnY5utRIY/xUEsxe6tm/F5Tw3E283zTUJMQ+
nrGWTrIWGOQZn4rdmWZsq8+xIhl/yFRotoowCtnB1KXaG0Ku6NDsaYnV3QdN4SBd
GCSQfGThVaU6cwILQSMs6navWxLqDYWZxdfLn532jch0ZzPf3XF7eCrZGfdzVNql
HNnaAUMYIdb7Gy6YojdnK5QuBVMMwYadRqUr/GM7Uv7hCRiXIoBrFwlVlR4Xg0Zg
zaME4WwssN0ORYN6UKE71gG34qyTTBUZcW55lZ0j52c=
//pragma protect end_data_block
//pragma protect digest_block
2cMBbusi566AhSztjHrwa+lqrLg=
//pragma protect end_digest_block
//pragma protect end_protected

  /**
    @grouphdr port_interleaving_check Port interleaving checks
    This group contains checks for port interleaving. 
    */

/**
    @grouphdr trace_tag_validity_check trace_tag related checks
    This group contains checks for trace_tag feature. 
    */


  typedef enum {LEGAL_TRANSITION,
                ILLEGAL_TRANSACTION_START_STATE,
                ILLEGAL_COHERENT_RESPONSE, 
                ILLEGAL_COHERENT_TRANSACTION,
                ILLEGAL_SNOOP_RESP_FOR_INITIAL_STATE,
                ILLEGAL_SNOOP_RESPONSE, 
                ILLEGAL_SNOOP_TRANSACTION
               } coherency_error_type_enum ;


  local svt_axi_port_configuration cfg;

  local svt_axi_transaction barrier_xact_queue[$];

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
yff2TGvx4UCB9yJRSBrNx+mw5MGGcrCmiEVM5yrXcFbN5RiPlsr6/PTEhoEZO/in
JMRSRnWo53La8KTuCHIUO0QBQEQoDJhY3xrJGTQB/1zsoZS3pARP4N70NHPkvAtB
eJ6kEsZ93SAIrc2OvWJTTYwnD9zOZ7XtK0/mEmrweHV3ResqKXirEg==
//pragma protect end_key_block
//pragma protect digest_block
Nrzh1DxwnFI+Eeh9KFVVdmQDPs8=
//pragma protect end_digest_block
//pragma protect data_block
j7vyo63ss7UKEZMY2bLdtErZ/iO4eHdDwKqpms+RgXlQODYpM8ENrarCFLkjQUkm
kRBFHKk8knIBCQhEA8ey6YWON+QTsVSw27zfDyIIDgx0Q0vUc2/S7D2Goj6f62sD
kZ7ULTvH6Mr6CWemEZI3AdLkf7Plo740052WvU/r2+OWTy8bVDzdUqVgHsFDoocj
SyLx7ESx5jbWypkXOxoHI4B8N4AbSOSHZhexSIUxoTbjC7CbNTLUYcDA/Y1j19Ji
rBI3opmAh99xodOcTAvIABhzXEt9gJUjgGCtmgcjby5uEPBJVYEM1ZGc4/NMkjlD
K+ALXXmAOdso3cS2YX+05KDpEXZnZU1uqTyNesuhIAWQntcHZc87oH8BB/5292VT

//pragma protect end_data_block
//pragma protect digest_block
CHr7D9AGPU32WiRkAHsMsRc0hks=
//pragma protect end_digest_block
//pragma protect end_protected
  local string group_name = "";

  local string sub_group_name = "";

  /** String used in macros */
  local string macro_str = "";
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
s+PNdA4yubhcvyRXQ3PhyRY4I/BJAX3M6lEuPx8czvpcnFTmDgItmcUSprKNAYVS
NkmIkmgZsnBsquT3hgFMGJ/w8De1FYIPqB/lBN2Vfhq8kCx4sCtUj6MCuVd4x4aQ
MOpGySj0fl58mAhQQyYFGXwGPOGrF6C9zaAYQzooeAw5IRZCvMvvEw==
//pragma protect end_key_block
//pragma protect digest_block
zXIY0/f+3NOm9z62G7hibdiLQfc=
//pragma protect end_digest_block
//pragma protect data_block
oD775LO8AhLSiOlUo2lC3STzBN/fk8tKgrSGFpRvRnKg1SMmhb7/YskSxoL9Dd1U
wwGK64vfKim2g0ytc0jzq6h8mbTB1YcLAmcBSNrh3R+DABYR0aeyGxG5RqXwPW8s
juN2kFxMjLPrZ3kqwpQKnlYjt9wCVoeSXCcKq0RvZ8z3gnOCFqVZhqFZ31tfl31U
GLB3NEXkDVHEMfcznVoCjn5k+BvOUGX80i1pA6DenTGaR6FwLZCZ3yQgKEQVbWAS
poyMnvmnHPEVbjqmBPpxSefGdlHvRjk0gQTE1JIdCCOUTT2XekOPeHHQFwi8gfvl
UoBikHTN763pfqq0lmRj4Pw3JV0PBniZik/BYvEf/uWP/pv+VXWGGuViSDlMoiEw
/UdKWyCQKeth0j9oWiReLd5FQtKIToYQTAfNKFoprlIDgMXJB4V/wHWt9umLf/lz
KoZjPwkf1B/zphj8L1dJbsmLiXA9g271+/y7b3okZCo5qZV8oL61JHZIGu/RVZLM
er3EnxxPCgIoAaEvm4k9t3UYsY5t6TfSPHBPVbSfpfi2dxg3l4zCD8d1Af3nrbrf
6oU3poQL1VknR/q6ch61aLkWpwcL6XDrmoiHJaH50x0UI/zsXTM+7CkqR7pQAi+Q
OblFhPXtss1MJxnTbARANg==
//pragma protect end_data_block
//pragma protect digest_block
lMdK5pWfVt7EUIi42vqbrqwPXc0=
//pragma protect end_digest_block
//pragma protect end_protected
  logic previous_reset = 1;

  /** Delay from ARVALID assertion to ARREADY assertion */
  local int arvalid_arready_delay = 0;
  
  /** Delay from ACVALID assertion to ACREADY assertion */
  local int acvalid_acready_delay = 0;
  
  /** Delay from ACVALID assertion to ACREADY assertion */
  local int cdvalid_cdready_delay = 0;
  
  /** Delay from CRVALID assertion to CRREADY assertion */
  local int crvalid_crready_delay = 0;

  /** Delay from TVALID assertion to TREADY assertion */
  local int tvalid_tready_delay = 0;

  /** Last sampled values in read address channel */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_arid;
  local logic[`SVT_AXI_MAX_ADDR_WIDTH-1:0] previous_araddr;
  local logic[`SVT_AXI_MAX_BURST_LENGTH_WIDTH-1:0] previous_arlen;
  local logic[`SVT_AXI_SIZE_WIDTH-1:0] previous_arsize;
  local logic[`SVT_AXI_BURST_WIDTH-1:0] previous_arburst;
  local logic[`SVT_AXI_LOCK_WIDTH-1:0] previous_arlock;
  local logic[`SVT_AXI_CACHE_WIDTH-1:0] previous_arcache;
  local logic[`SVT_AXI_PROT_WIDTH-1:0] previous_arprot;
  local logic[`SVT_AXI_QOS_WIDTH-1:0] previous_arqos;
  local logic[`SVT_AXI_REGION_WIDTH-1:0] previous_arregion;
  local logic[`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] previous_aruser;
  local logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] previous_ardomain;
  local logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] previous_arsnoop;
  local logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] previous_arbar;
`ifdef SVT_ACE5_ENABLE
  local logic  previous_archunken;
  local logic[`SVT_AXI_MAX_MPAM_WIDTH-1:0] previous_armpam;
`endif
  
  local logic[`SVT_AXI_ACE_SNOOP_RESP_WIDTH-1:0] previous_crresp;
  local logic[`SVT_AXI_ACE_SNOOP_DATA_WIDTH-1:0] previous_cddata;
  local logic[`SVT_AXI_ACE_SNOOP_ADDR_WIDTH-1:0] previous_acaddr;
  local logic[`SVT_AXI_ACE_SNOOP_TYPE_WIDTH-1:0] previous_acsnoop; 
  local logic[`SVT_AXI_ACE_SNOOP_PROT_WIDTH-1:0] previous_acprot;
  local logic previous_aridunq;
  local logic previous_cdlast;

  /** holds number of databeat transferred over snoop data channel for current snoop request */
  local int unsigned cddata_beat_count = 0;

  /** Delay from RVALID assertion to RREADY assertion */
  local int rvalid_rready_delay = 0;

  /** Last sampled value of RID */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_rid;

  /** Last sampled value of RIDUNQ */
  local logic previous_ridunq;

  /** Last sampled value of RRESP */
  local logic[`SVT_AXI_RESP_WIDTH-1:0] previous_rresp;

  /** Last sampled value of RDATA */
  local logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] previous_rdata;

  /** Last sampled value of RLAST */
  local logic previous_rlast;

  /** Last sampled value of RUSER */
  local logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] previous_ruser;

`ifdef SVT_ACE5_ENABLE
  /** Last sampled value of RCHUNKV */
  local logic  previous_rchunkv;

  /** Last sampled value of RCHUNKNUM */
  local logic [`SVT_AXI_MAX_CHUNK_NUM_WIDTH-1:0] previous_rchunknum;

  /** Last sampled value of RCHUNKSTRB */
  local logic [`SVT_AXI_MAX_CHUNK_STROBE_WIDTH-1:0] previous_rchunkstrb;
`endif 

  /** Delay from AWVALID assertion to AWREADY assertion */
  local int awvalid_awready_delay = 0;

  /** Last sampled values in write address channel */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_awid;
  local logic[`SVT_AXI_MAX_ADDR_WIDTH-1:0] previous_awaddr;
  local logic[`SVT_AXI_MAX_BURST_LENGTH_WIDTH-1:0] previous_awlen;
  local logic[`SVT_AXI_SIZE_WIDTH-1:0] previous_awsize;
  local logic[`SVT_AXI_BURST_WIDTH-1:0] previous_awburst;
  local logic[`SVT_AXI_LOCK_WIDTH-1:0] previous_awlock;
  local logic[`SVT_AXI_CACHE_WIDTH-1:0] previous_awcache;
  local logic[`SVT_AXI_PROT_WIDTH-1:0] previous_awprot;
  local logic[`SVT_AXI_QOS_WIDTH-1:0] previous_awqos;
  local logic[`SVT_AXI_REGION_WIDTH-1:0] previous_awregion;
  local logic[`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] previous_awuser;
  local logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] previous_awdomain;
  local logic[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] previous_awsnoop;
  local logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] previous_awbar;
  local logic[`SVT_AXI_MAX_MPAM_WIDTH-1:0] previous_awmpam;
  local logic previous_awunique;
  local logic previous_awidunq;

  /** Delay from WVALID assertion to WREADY assertion */
  local int wvalid_wready_delay = 0;

  /** Last sampled value of WID */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_wid;

  /** Last sampled value of WDATA */
  local logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] previous_wdata;

  /** Last sampled value of WSTRB */
  local logic[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] previous_wstrb;

  /** Last sampled value of WUSER */
  local logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] previous_wuser;

  /** Last sampled value of WLAST */
  local logic previous_wlast;

  /** Delay from BVALID assertion to BREADY assertion */
  local int bvalid_bready_delay = 0;

  /** Last sampled value of BID */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_bid;

  /** Last sampled value of BIDUNQ */
  local logic previous_bidunq;

  /** Last sampled value of BRESP */
  local logic[`SVT_AXI_RESP_WIDTH-1:0] previous_bresp;

  /** Last sampled value of BUSER */
  local logic[`SVT_AXI_MAX_BRESP_USER_WIDTH-1:0] previous_buser;

  local logic[`SVT_AXI_MAX_TDATA_WIDTH-1:0] previous_tdata;
  local logic[`SVT_AXI_TSTRB_WIDTH-1:0] previous_tstrb;
  local logic[`SVT_AXI_TKEEP_WIDTH-1:0] previous_tkeep;
  local logic previous_tlast;
  local logic[`SVT_AXI_MAX_TID_WIDTH-1:0] previous_tid;
  local logic[`SVT_AXI_MAX_TDEST_WIDTH-1:0] previous_tdest;
  local logic[`SVT_AXI_MAX_TUSER_WIDTH-1:0] previous_tuser;

  `ifdef SVT_AXI_QVN_ENABLE
  /** Variables used in QVN token handshake signal checks */  
  local bit is_varvalidvn_deassertion_check_en [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local bit is_varqosvn_valid_change_check_en  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];

  local bit is_vawvalidvn_deassertion_check_en [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local bit is_vawqosvn_valid_change_check_en  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];

  local bit is_vwvalidvn_deassertion_check_en  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];

  local int unsigned qvn_ar_token_request_ready_timeout_counter_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];
  local int unsigned qvn_aw_token_request_ready_timeout_counter_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];
  local int unsigned qvn_w_token_request_ready_timeout_counter_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];
 
  local logic previous_varvalidvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic [3:0] previous_varqosvnx [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic previous_varreadyvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0]; 
   
  local logic previous_vawvalidvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic [3:0] previous_vawqosvnx [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic previous_vawreadyvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0]; 
  
  local logic previous_vwvalidvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic previous_vwreadyvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0]; 

  `endif

  local svt_axi_snoop_transaction  multipart_dvm_snoop_xact;
  svt_axi_transaction multipart_dvm_coherent_xact;
  local svt_axi_transaction        active_multipart_dvm_coherent_q[svt_axi_transaction];
  local svt_axi_snoop_transaction  active_multipart_dvm_snoop_q[svt_axi_snoop_transaction];

  //local svt_axi_snoop_transaction  multipart_dvm_snoop_check_guard_xact;
  //local svt_axi_master_transaction multipart_dvm_coherent_check_guard_xact;
  local svt_axi_transaction        active_multipart_dvm_coherent_check_guard_q[svt_axi_transaction];
  local svt_axi_snoop_transaction  active_multipart_dvm_snoop_check_guard_q[svt_axi_snoop_transaction];

  /** Enables protocol check coverage provided it protocol_checks_coverage_enable is set
    * in the port configuration as well. If enable_pc_cov is 0, then protocol checks coverage
    * will not be enabled, even if it is set in configuration
    */
  local bit enable_pc_cov = 1;

  /** indicates if only partial ID bits are considered for exclusive transaction */
  local bit partial_exclusive_id = 0;
  

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
TixcyPsNnKO1ckrG8zDjYksxdVx/ioJo3l+aYilAfPsC4RObfwUrHQqTuH5pJPGT
cDmS4S0kc/jZf0cLpTbobjZW+okb2nqDcjRDB/53fowu7iFzkDNX4YDpZxjdrusF
/mTuTH9GNn8ktORkMhCiSWqfdlq6g3ikmYiT2JuQu5fCaNfO3xl0CA==
//pragma protect end_key_block
//pragma protect digest_block
iwRMHbqxq+/cKFkO8Q6C2Y34d3w=
//pragma protect end_digest_block
//pragma protect data_block
L+qHQwq3N2w7AIds5tjVWXTSzDQ8uwiuUvF4s13GWPmcIOWzgRhlkbDy9qiX/pIm
neq9qmRBxrMTBMnMjOcEbisCYDqi4do6d45+L22tBDFjvl4yHx/9Ip3PmSRKgVi8
9Cuf416uPU9KwL6+zJBRQafYmD5kclWxOl4cdFs/Jb74GK2yQ8JuPuJlcBXYIiOX
t72IuSRV0cA7EO3Lu4gZkl8UNK7Gp6ESihHrQoc/NXOL/WyXjlibaJPBz7eNpcDi
O5/vkcmkZWAZs/yssTddOVk7X1oj/UcDwkYTCN3XPEwvad1SxTWDOShxXrH9SHd6
UF6PMMti2G57HqHfnBfwTAEeclsKdZjkeGElGudIn4TJZTlQiwjnWq2k/QIY3vyk
AHupVEic7ZkquJcqzOscBwcGzwdoW1x5gPFKaEPBkd5NOkH7FUk3XUiMOzoSxi+/
KqsNTjE/IKKU5YgV8dgWsk0fU0C+H3eRyUOI3JMlDlM=
//pragma protect end_data_block
//pragma protect digest_block
MaoLsb840IEPXMpbQjF231yeF70=
//pragma protect end_digest_block
//pragma protect end_protected


  //--------------------------------------------------------------
  /** Checks that ARID is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arid_when_arvalid_high_check;

  /** Checks that ARADDR is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_araddr_when_arvalid_high_check;

  /** Checks that ARLEN is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arlen_when_arvalid_high_check;
  
  /** Checks that ARSIZE is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arsize_when_arvalid_high_check;
  
  /** Checks that ARLEN and ARSIZE are valid for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_arlen_arsize_check;
  
  /** Checks that ARCACHE is valid for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_arcache_check;
  
  /** Checks that address is aligned for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_read_addr_aligned_check;
  
  /** Checks that AWLEN and AWSIZE are valid for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_awlen_awsize_check;
  
  /** Checks that AWCACHE is valid for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_awcache_check;
  
  /** Checks that address is aligned for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_write_addr_aligned_check;

  /** Checks that address is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_addr_check;
  
  /** Checks that received write data is not interleaved beyond write_data_interleave_depth value
    * An error is issued if write data is interleaved beyond this value for Write data interleaving */
  svt_err_check_stats write_data_interleave_depth_check;
 
  /** Checks that the order in which a slave receives the first data item of each transaction must be the
    * same as the order in which it receives the addresses for the transactions for Write Data Interleaving 
    * transactions */
  svt_err_check_stats write_data_interleave_order_check;

 /** Checks that id is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_id_check;

  /** Checks that response generated for exclusive load accesss is correct */
  svt_err_check_stats exclusive_load_response_check;

  /** Checks that response generated for exclusive store accesss is correct */
  svt_err_check_stats exclusive_store_response_check;

  /** Checks that master does not permit an Exclusive Store transaction to be
    * in progress at the same time as any transaction that registers that it
    * is performing an Exclusive sequence
    */
  svt_err_check_stats exclusive_store_overlap_with_another_exclusive_sequence_check;

  /** Checks that, once a master receives successful exclusive store response EXOKAY
    * from interconnect, then no other master should be provided with EXOKAY response,
    * until current master acknowledges completing successful exclusive store by asserting RACK
    */
   svt_err_check_stats exokay_not_sent_until_successful_exclusive_store_rack_observed_check;
  
    /** Checks that READ_ONLY_INTERFACE supports only read transactions 
     * Applicable only for AXI4 VIP
     * Passive Master,Passive Slave and Active slave will perform this
     * check
     */
     svt_err_check_stats read_xact_on_read_only_interface_check;
   
    /** Checks that WRITE_ONLY_INTERFACE supports only write transactions 
     * Applicable only for AXI4 VIP
     * Passive Master,Passive Slave and Active slave will perform this
     * check
     */
     svt_err_check_stats write_xact_on_write_only_interface_check;
     
     /** Checks that READ_ONLY_INTERFACE does not support exclusive access  
     * Applicable only for AXI4 VIP
     * Passive Master,Passive Slave and Active slave will perform this 
     * check
     */
     svt_err_check_stats excl_access_on_read_only_interface_check;

      /** Checks that WRITE_ONLY_INTERFACE does not support exclusive access  
      * Applicable only for AXI4 VIP
      * Passive Master,Passive Slave and Active slave will perform this 
      * check
      */
      svt_err_check_stats excl_access_on_write_only_interface_check;
     
     /** Checks that burst length is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_burst_length_check;
  
  /** Checks that burst size is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_burst_size_check;
  
  /** Checks that burst type is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_burst_type_check;
  
  /** Checks that cache type is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_cache_type_check;
  
  /** Checks that protection type is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_prot_type_check;
  
  /** Checks that exclusive transaction sent on AXI_ACE interface are
   * only of WRITENOSNOOP, READNOSNOOP, READCLEAN, READSHARED and CLEANUNIQUE type */
  svt_err_check_stats exclusive_ace_transaction_type_check;

  /** Checks that ARADDR[2:0] for multipart dvm xact is not other than SBZ */
  svt_err_check_stats signal_araddr_multipart_dvm_xact_check;

  /** Checks that ARBURST is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arburst_when_arvalid_high_check;

  /** Checks that ARLOCK is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arlock_when_arvalid_high_check;

  /** Checks that ARCACHE is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arcache_when_arvalid_high_check;

  /** Checks that ARPROT is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arprot_when_arvalid_high_check;

  /** Checks that ARQOS is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arqos_when_arvalid_high_check;

  /** Checks that ARREGION is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arregion_when_arvalid_high_check;

  /** Checks that ARUSER is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_aruser_when_arvalid_high_check;
  
    /** Checks that ARDOMAIN is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_ardomain_when_arvalid_high_check;
  
  /** Checks that ARSNOOP is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arsnoop_when_arvalid_high_check;
  
  /** Checks that ARBAR is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arbar_when_arvalid_high_check;

  /** Checks that ARREADY is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arready_when_arvalid_high_check;

  /** Checks that AWDOMAIN is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awdomain_when_awvalid_high_check;
  
  /** Checks that AWSNOOP is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awsnoop_when_awvalid_high_check;
  
  /** Checks that AWBAR is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awbar_when_awvalid_high_check;
  //--------------------------------------------------------------
  /** Checks that ARID is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arid_when_arvalid_high_check;

  /** Checks that ARADDR is stable when ARVALID is high */
  svt_err_check_stats signal_stable_araddr_when_arvalid_high_check;

  /** Checks that RACK is asserted for a single cycle */
  svt_err_check_stats signal_rack_single_cycle_high_check;

  /** Checks that RACK signal must be asserted the cycle after the associated handshake or later */
  svt_err_check_stats signal_rack_after_handshake_check;

  /** Checks that WACK is asserted for a single cycle */
  svt_err_check_stats signal_wack_single_cycle_high_check;

  /** Checks that WACK signal must be asserted the cycle after the associated handshake or later */
  svt_err_check_stats signal_wack_after_handshake_check;

  /** Checks that ARLEN is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arlen_when_arvalid_high_check;
  
  /** Checks that ARSIZE is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arsize_when_arvalid_high_check;

  /** Checks that ARBURST is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arburst_when_arvalid_high_check;

  /** Checks that ARLOCK is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arlock_when_arvalid_high_check;

  /** Checks that ARCACHE is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arcache_when_arvalid_high_check;

  /** Checks that ARPROT is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arprot_when_arvalid_high_check;

  /** Checks that ARQOS is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arqos_when_arvalid_high_check;

  /** Checks that ARREGION is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arregion_when_arvalid_high_check;

  /** Checks that ARUSER is stable when ARVALID is high */
  svt_err_check_stats signal_stable_aruser_when_arvalid_high_check;
  
  /** Checks that ARDOMAIN is stable when ARVALID is high */
  svt_err_check_stats signal_stable_ardomain_when_arvalid_high_check;
  
  /** Checks that ARSNOOP is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arsnoop_when_arvalid_high_check;
  
  /** Checks that ARBAR is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arbar_when_arvalid_high_check;

  /** Checks that AWDOMAIN is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awdomain_when_awvalid_high_check;
  
  /** Checks that AWSNOOP is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awsnoop_when_awvalid_high_check;
  
  /** Checks that AWBAR is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awbar_when_awvalid_high_check;
  //--------------------------------------------------------------
  /** Checks that RID is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rid_when_rvalid_high_check;

  /** Checks that RDATA is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rdata_when_rvalid_high_check;

  /** Checks that RDATACHK is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rdatachk_when_rvalid_high_check;
 
  /** Checks that rpoison is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rpoison_when_rvalid_high_check;
 
  /** Checks that RUSER is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_ruser_when_rvalid_high_check;

  /** Checks that RRESP is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rresp_when_rvalid_high_check;

  /** Checks that RLAST is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rlast_when_rvalid_high_check;

  /** Checks that RREADY is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rready_when_rvalid_high_check;

  /** Checks that RID is stable when RVALID is high */
  svt_err_check_stats signal_stable_rid_when_rvalid_high_check;

  /** Checks that RUSER is stable when RVALID is high */
  svt_err_check_stats signal_stable_ruser_when_rvalid_high_check;

  /** Checks that RDATA is stable when RVALID is high */
  svt_err_check_stats signal_stable_rdata_when_rvalid_high_check;

  /** Checks that RRESP is stable when RVALID is high */
  svt_err_check_stats signal_stable_rresp_when_rvalid_high_check;

  /** Checks that RLAST is stable when RVALID is high */
  svt_err_check_stats signal_stable_rlast_when_rvalid_high_check;

  /** Checks that sample read data has associated address */
  svt_err_check_stats read_data_follows_addr_check;
  //--------------------------------------------------------------
  /** Checks that AWID is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awid_when_awvalid_high_check;

  /** Checks that valid write strobes are driven */
  svt_err_check_stats valid_write_strobe_check;

`ifdef SVT_ACE5_ENABLE 
  //--------------------------------------------------------------
 /** Checks that stash_nid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_stash_nid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that stash_lpid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_stash_lpid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that stash_nid_valid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_stash_nid_valid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that stash_lpid_valid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_stash_lpid_valid_when_awvalid_high_check;

  //--------------------------------------------------------------
 /** Checks that awmmusid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmusid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that awmmussid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmussid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that  is awmmusecsid not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmusecsid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that awmmussidv is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmussidv_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that awmmuatst is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmuatst_when_awvalid_high_check;

  //--------------------------------------------------------------
 /** Checks that armmusid is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmusid_when_arvalid_high_check;

 //--------------------------------------------------------------
/** Checks that armmussid is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmussid_when_arvalid_high_check;

 //--------------------------------------------------------------
/** Checks that  is armmusecsid not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmusecsid_when_arvalid_high_check;

 //--------------------------------------------------------------
/** Checks that armmussidv is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmussidv_when_arvalid_high_check;

 //--------------------------------------------------------------
/** Checks that armmuatst is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmuatst_when_arvalid_high_check;

 /** Checks that awatop is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awatop_when_awvalid_high_check;

 /** Checks that armpam is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armpam_when_arvalid_high_check;

 /** Checks that awmpam is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmpam_when_awvalid_high_check;

   /** Checks that AWMPAM is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awmpam_when_awvalid_high_check;

  /** Checks that ARMPAM is stable when ARVALID is high */
  svt_err_check_stats signal_stable_armpam_when_arvalid_high_check;
`endif

`ifdef SVT_ACE5_ENABLE 
//--------------------------------------------------------------
 /** Checks that ARIDUNQ is not X or Z when ARVALID is high*/
   svt_err_check_stats signal_valid_aridunq_when_arvalid_high_check;

 /** Checks that RIDUNQ is not X or Z when RVALID is high*/
   svt_err_check_stats signal_valid_ridunq_when_rvalid_high_check;

 /** Checks that AWIDUNQ is not X or Z when AWVALID is high*/
   svt_err_check_stats signal_valid_awidunq_when_awvalid_high_check;

 /** Checks that BIDUNQ is not X or Z when BVALID is high*/
   svt_err_check_stats signal_valid_bidunq_when_bvalid_high_check;
   
//--------------------------------------------------------------
/** Checks that ARIDUNQ is stable when ARVALID is high */
  svt_err_check_stats signal_stable_aridunq_when_arvalid_high_check;

/** Checks that RIDUNQ is stable when RVALID is high */
  svt_err_check_stats signal_stable_ridunq_when_rvalid_high_check;

/** Checks that AWIDUNQ is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awidunq_when_awvalid_high_check;

/** Checks that BIDUNQ is stable when BVALID is high */
  svt_err_check_stats signal_stable_bidunq_when_bvalid_high_check;

//--------------------------------------------------------------
  /** Checks that RIDUNQ asserted or deasserted when ARIDUNQ asserted or deasserted */
  //svt_err_check_stats ridunq_asserted_deasserted_check;

  /** Checks that BIDUNQ asserted or deasserted when AWIDUNQ asserted or deasserted*/
  //svt_err_check_stats bidunq_asserted_deasserted_check;
 
  /** Checks that there is no outstanding transaction with same arid */
  svt_err_check_stats no_outstanding_read_unique_transaction_with_same_arid;

  /** Checks that there is no outstanding transaction with same awid */
  svt_err_check_stats no_outstanding_write_unique_transaction_with_same_awid;
`endif

  /** Checks that AWADDR is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awaddr_when_awvalid_high_check;

  /** Checks that AWLEN is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awlen_when_awvalid_high_check;
  
  /** Checks that AWSIZE is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awsize_when_awvalid_high_check;

  /** Checks that AWBURST is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awburst_when_awvalid_high_check;

  /** Checks that AWLOCK is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awlock_when_awvalid_high_check;

  /** Checks that AWCACHE is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awcache_when_awvalid_high_check;

  /** Checks that AWPROT is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awprot_when_awvalid_high_check;

  /** Checks that AWREADY is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awready_when_awvalid_high_check;

  /** Checks that AWQOS is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awqos_when_awvalid_high_check;

  /** Checks that AWREGION is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awregion_when_awvalid_high_check;

  /** Checks that AWUNIQUE is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awunique_when_awvalid_high_check;

  /** Checks that AWUSER is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awuser_when_awvalid_high_check;
  //--------------------------------------------------------------
  /** Checks that AWID is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awid_when_awvalid_high_check;

  /** Checks that AWADDR is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awaddr_when_awvalid_high_check;

  /** Checks that AWLEN is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awlen_when_awvalid_high_check;
  
  /** Checks that AWSIZE is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awsize_when_awvalid_high_check;

  /** Checks that AWBURST is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awburst_when_awvalid_high_check;

  /** Checks that AWLOCK is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awlock_when_awvalid_high_check;

  /** Checks that AWCACHE is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awcache_when_awvalid_high_check;

  /** Checks that AWPROT is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awprot_when_awvalid_high_check;

  /** Checks that AWQOS is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awqos_when_awvalid_high_check;

  /** Checks that AWREGION is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awregion_when_awvalid_high_check;

  /** Checks that AWUNIQUE is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awunique_when_awvalid_high_check;

  /** Checks that AWUSER is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awuser_when_awvalid_high_check;

  //--------------------------------------------------------------

  /** Checks that WID is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wid_when_wvalid_high_check;

  /** Checks that WUSER is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wuser_when_wvalid_high_check;

  /** Checks that WDATA is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wdata_when_wvalid_high_check;

  /** Checks that WDATACHK is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wdatachk_when_wvalid_high_check;

 /** Checks that WPOISON is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wpoison_when_wvalid_high_check;

  /** Checks that WSTRB is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wstrb_when_wvalid_high_check;

  /** Checks that WLAST is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wlast_when_wvalid_high_check;

  /** Checks that WREADY is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wready_when_wvalid_high_check;

  /** Checks that WID is stable when WVALID is high */
  svt_err_check_stats signal_stable_wid_when_wvalid_high_check;

  /** Checks that WUSER is stable when WVALID is high */
  svt_err_check_stats signal_stable_wuser_when_wvalid_high_check;

  /** 
   * Checks that WDATA is stable when WVALID is high 
   * When svt_axi_port_configuration::check_valid_data_bytes_only_enable=1 ,
   * it considers only valid byte lanes of wdata based on wstrb. 
   * When svt_axi_port_configuration::check_valid_data_bytes_only_enable=0 ,
   * whole wdata as seen on the bus will be considered.
   */
  svt_err_check_stats signal_stable_wdata_when_wvalid_high_check;

  /** Checks that WSTRB is stable when WVALID is high */
  svt_err_check_stats signal_stable_wstrb_when_wvalid_high_check;

  /** Checks that WLAST is stable when WVALID is high */
  svt_err_check_stats signal_stable_wlast_when_wvalid_high_check;

  //--------------------------------------------------------------
  /** Checks that BID is not X or Z when BVALID is high */
  svt_err_check_stats signal_valid_bid_when_bvalid_high_check;

  /** Checks that BUSER is not X or Z when BVALID is high */
  svt_err_check_stats signal_valid_buser_when_bvalid_high_check;

  /** Checks that BRESP is not X or Z when BVALID is high */
  svt_err_check_stats signal_valid_bresp_when_bvalid_high_check;

  /** Checks that BREADY is not X or Z when BVALID is high */
  svt_err_check_stats signal_valid_bready_when_bvalid_high_check;

  /** Checks that BID is stable when BVALID is high */
  svt_err_check_stats signal_stable_bid_when_bvalid_high_check;

  /** Checks that BUSER is stable when BVALID is high */
  svt_err_check_stats signal_stable_buser_when_bvalid_high_check;

  /** Checks that BRESP is stable when BVALID is high */
  svt_err_check_stats signal_stable_bresp_when_bvalid_high_check;

  /** 
    * When a write response is sampled, checks that there is a 
    * transaction with corresponding ID whose data phase is complete 
    */
  svt_err_check_stats write_resp_follows_last_write_xfer_check;

  /** 
    * Checks that WLAST is asserted for the last beat of write data. 
    */
  svt_err_check_stats wlast_asserted_for_last_write_data_beat;

  //--------------------------------------------------------------
  // Checks that need to be executed externally (by monitor).
  /** Checks that ARVALID is not X or Z */
  svt_err_check_stats signal_valid_arvalid_check;

  /** Checks that RVALID is not X or Z */
  svt_err_check_stats signal_valid_rvalid_check;

  /** Checks that AWVALID is not X or Z */
  svt_err_check_stats signal_valid_awvalid_check;

  /** Checks that WVALID is not X or Z */
  svt_err_check_stats signal_valid_wvalid_check;

  /** Checks that BVALID is not X or Z */
  svt_err_check_stats signal_valid_bvalid_check;
  
  /** Checks that ACVALID is not X or Z */
  svt_err_check_stats signal_valid_acvalid_check;
  
  /** Checks that CDVALID is not X or Z */
  svt_err_check_stats signal_valid_cdvalid_check;
  
  /** Checks that CDVALID is not X or Z */
  svt_err_check_stats signal_valid_crvalid_check;

  /** Checks that ARVALID is not X or Z During Reset */
  svt_err_check_stats signal_valid_arvalid_check_during_reset;

  /** Checks that RVALID is not X or Z During Reset*/
  svt_err_check_stats signal_valid_rvalid_check_during_reset;

  /** Checks that AWVALID is not X or Z During Reset*/
  svt_err_check_stats signal_valid_awvalid_check_during_reset;

  /** Checks that WVALID is not X or Z During Reset*/
  svt_err_check_stats signal_valid_wvalid_check_during_reset;

  /** Checks that BVALID is not X or Z During Reset */
  svt_err_check_stats signal_valid_bvalid_check_during_reset;

  /** Checks if arvalid was interrupted before arready got asserted */
  svt_err_check_stats arvalid_interrupted_check;
  
  /** Checks if acvalid was interrupted before acready got asserted */
  svt_err_check_stats acvalid_interrupted_check;
  
  /** Checks if cdvalid was interrupted before cdrready got asserted */
  svt_err_check_stats cdvalid_interrupted_check;
  
  /** Checks if crvalid was interrupted before crready got asserted */
  svt_err_check_stats crvalid_interrupted_check;

  /** Checks if rvalid was interrupted before rready got asserted */
  svt_err_check_stats rvalid_interrupted_check;

  /** Checks if awvalid was interrupted before awready got asserted */
  svt_err_check_stats awvalid_interrupted_check;

  /** Checks if wvalid was interrupted before wready got asserted */
  svt_err_check_stats wvalid_interrupted_check;

  /** Checks if bvalid was interrupted before bready got asserted */
  svt_err_check_stats bvalid_interrupted_check;
  //--------------------------------------------------------------
  /** Checks if rvalid is low when reset is active */
  svt_err_check_stats rvalid_low_when_reset_is_active_check;

  /** Checks if bvalid is low when reset is active */
  svt_err_check_stats bvalid_low_when_reset_is_active_check;

  /** Checks if arvalid is low when reset is active */
  svt_err_check_stats arvalid_low_when_reset_is_active_check;

  /** Checks if acvalid is low when reset is active */
  svt_err_check_stats acvalid_low_when_reset_is_active_check;
  
  /** Checks if crvalid is low when reset is active */
  svt_err_check_stats crvalid_low_when_reset_is_active_check;
  
  /** Checks if cdvalid is low when reset is active */
  svt_err_check_stats cdvalid_low_when_reset_is_active_check;

  /** Checks if awvalid is low when reset is active */
  svt_err_check_stats awvalid_low_when_reset_is_active_check;

  /** Checks if wvalid is low when reset is active */
  svt_err_check_stats wvalid_low_when_reset_is_active_check;
  //--------------------------------------------------------------
  
  /** Checks if write burst cross a 4KB boundary */
  svt_err_check_stats awaddr_4k_boundary_cross_active_check;
  //--------------------------------------------------------------

  /** Checks if write burst of WRAP type has an aligned address*/
  svt_err_check_stats awaddr_wrap_aligned_active_check ;
  //--------------------------------------------------------------
  
  /** Checks if write burst of WRAP type has a valid length*/
  svt_err_check_stats awlen_wrap_active_check;
  //--------------------------------------------------------------

  /** Checks if size of write transfer exceeds the width of the data bus*/
  svt_err_check_stats awsize_data_width_active_check;
  //--------------------------------------------------------------
        
  /** Checks if the value of awburst=2'b11 when awvalid is high*/
  svt_err_check_stats awburst_reserved_val_check;
  //--------------------------------------------------------------
  
  /** Checks if the value of awcache[3:2]=2'b00 when awvalid is high and awcache[1] is also low*/
  svt_err_check_stats awvalid_awcache_active_check;
  //--------------------------------------------------------------

  
  /** Checks if read burst cross a 4KB boundary */
  svt_err_check_stats araddr_4k_boundary_cross_active_check;
  //--------------------------------------------------------------

  /** Checks if read  burst of WRAP type has an aligned address*/
  svt_err_check_stats araddr_wrap_aligned_active_check ;
  //--------------------------------------------------------------

  /** Checks if snoop address is aligned with snoop data width */
  svt_err_check_stats acaddr_aligned_to_cddata_width_valid_check ;
  //--------------------------------------------------------------

  /** Checks that a cached master does not initiate WriteUnique or WriteLineUnique
    * coherent write transaction while any WriteBack, WriteClean or WriteEvict transaction
    * is outstanding.
    */
  svt_err_check_stats complete_outstanding_memory_write_before_writeunique_writelineunique_check ;

  /** Checks that a cached master does not issue WriteBack, WriteClean or WriteEvict
    * transaction while any WriteUnique or WriteLineUnique coherent write transaction
    * is in progress.
    * It automatically checks second rule which says, Complete any incoming snoop 
    * transactions without the use of WriteBack, WriteClean, or WriteEvict
    * transactions while a WriteUnique or WriteLineUnique transaction is in progress.
    */
  svt_err_check_stats complete_outstanding_writeunique_writelineunique_before_memory_write_check ;


  /** Checks that CleanInvalid and MakeInvalid cache maintenance transactions are not 
    * initiated while any memory update or shareable transactions are outstanding. It
    * also checks that CleanShared cache maintenance transactions are not initiated 
    * while any memory update or any shareable transactions that can make the cacheline
    * dirty, are outstanding.
    */
  svt_err_check_stats cache_maintenance_outstanding_transaction_check ;

  /** Checks that WriteBack, WriteClean or any shareable transactions are not issued 
    * while cache maintenance transaction is in progress.
    */
  svt_err_check_stats no_memory_update_or_shareable_txn_during_cache_maintenance_check ;

  /** Monitor checks that when master initiates a CleanShared cache maintenance transaction, 
    * and receives any snoop transaction to the same cacheline, the initiating master must not
    * assert PassDirty snoop response. It also checks that when master initiates CleanInvalid
    * or MakeInvalid cache maintenance transactions, and receives any snoop transaction to the
    * same cacheline, the initiating master must not assert PassDirty, IsShared and DataTransfer
    * snoop responses.
    */
  svt_err_check_stats valid_snoop_response_during_cache_maintenance_check ;
  //--------------------------------------------------------------

  /** Checks if number of databeat transferred over snoop data channel is valid */
  svt_err_check_stats snoop_transaction_burst_length_check ;
  //--------------------------------------------------------------
  
  /** Checks if read burst of WRAP type has a valid length*/
  svt_err_check_stats arlen_wrap_active_check;
  //--------------------------------------------------------------

  /** Checks if size of read transfer exceeds the width of the data bus*/
  svt_err_check_stats arsize_data_width_active_check;
  //--------------------------------------------------------------
        
  /** Checks if the value of arburst=2'b11 when arvalid is high*/
  svt_err_check_stats arburst_reserved_val_check;
  //--------------------------------------------------------------
  
  /** Checks if the value of arcache[3:2]=2'b00 when arvalid is high and arcache[1] is also low*/
  svt_err_check_stats arvalid_arcache_active_check;
  //--------------------------------------------------------------
  
/** Checks if the number of write data items matches AWLEN for the corresponding address */
  svt_err_check_stats wdata_awlen_match_for_corresponding_awaddr_check;
  //--------------------------------------------------------------

/** Checks if the slave must only give a write response after the last write data item is transferred  */
  svt_err_check_stats write_resp_after_last_wdata_check;
  //--------------------------------------------------------------

/** Checks if  A slave must not give a write response before the write address */
  svt_err_check_stats write_resp_after_write_addr_check;
  //--------------------------------------------------------------

/** Checks if the number of read data items matches ARLEN for the corresponding address */
  svt_err_check_stats rdata_arlen_match_for_corresponding_araddr_check;
  //--------------------------------------------------------------

/** Checks if the number of read data items matches ARLEN for the corresponding address */
 svt_err_check_stats rlast_asserted_for_last_read_data_beat;
//ACE CHECKS//

  /** Checks that ACREADY is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_acready_when_arvalid_high_check;
  
  /** Checks that ACADDR is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_acaddr_when_acvalid_high_check;
  
  /** Checks that ACSNOOP is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_acsnoop_when_acvalid_high_check;
  
  /** Checks that ACPROT is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_acprot_when_acvalid_high_check;
  
  /** Checks that CDREADY is not X or Z when CDVALID is high */
  svt_err_check_stats signal_valid_cdready_when_cdvalid_high_check;
  
  /** Checks that CDDATA is not X or Z when CDVALID is high */
  svt_err_check_stats signal_valid_cddata_when_cdvalid_high_check;
  
  /** Checks that CDDATACHK is not X or Z when CDVALID is high */
  svt_err_check_stats signal_valid_cddatachk_when_cdvalid_high_check;
  
  /** Checks that CDPOISON is not X or Z when CDVALID is high */
  svt_err_check_stats signal_valid_cdpoison_when_cdvalid_high_check;

 /** Checks that ACREADY is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_cdlast_when_cdvalid_high_check;
  
  /** Checks that CRREADY is not X or Z when CRVALID is high */
  svt_err_check_stats signal_valid_crready_when_crvalid_high_check;
  
  /** Checks that CRRESP is not X or Z when CRVALID is high */
  svt_err_check_stats signal_valid_crresp_when_crvalid_high_check;

  /** Checks that ACADDR is stable when ARVALID is high */
  svt_err_check_stats signal_stable_acaddr_when_acvalid_high_check;
  
  /** Checks that ACSNOOP is stable when ARVALID is high */
  svt_err_check_stats signal_stable_acsnoop_when_acvalid_high_check;
  
  /** Checks that ACPROT is stable when ARVALID is high */
  svt_err_check_stats signal_stable_acprot_when_acvalid_high_check;

  /** Checks that CDDATA is stable when CDVALID is high */
  svt_err_check_stats signal_stable_cddata_when_cdvalid_high_check;
  
  /** Checks that ACREADY is stable when ARVALID is high */
  svt_err_check_stats signal_stable_cdlast_when_cdvalid_high_check;

  /** Checks that CRRESP is stable when CRVALID is high */
  svt_err_check_stats signal_stable_crresp_when_crvalid_high_check;
  
  
/**Checks if the Device transactions, as indicated by AxCACHE[1] = 0, must only use AxDOMAIN = 11.  */
 svt_err_check_stats axcache_axdomain_restriction_check;
  //--------------------------------------------------------------

/**Checks if the  AXCACHE and AXDOMAIN value are valid */
 svt_err_check_stats axcache_axdomain_invalid_value_check ;
  //--------------------------------------------------------------



/**Checks if the  AWSIZE is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_awsize_valid_value_check;
  //--------------------------------------------------------------
/**Checks if the  ARSIZE is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_arsize_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWLEN is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_awlen_valid_value_check;
  //--------------------------------------------------------------
/**Checks if the  ARLEN is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_arlen_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWSIZE is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_awsize_valid_check;
  //--------------------------------------------------------------

/**Checks if the  AWBURST is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_awburst_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  ARBURST is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_arburst_valid_value_check;
  //--------------------------------------------------------------

 /**Checks if the  ARSIZE is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_arsize_valid_check;
  //--------------------------------------------------------------

/**Checks if the  address is aligned for AWBURST in  Cache Line Size Transactions */
 svt_err_check_stats cache_line_awburst_wrap_addr_aligned_valid_check;
  //--------------------------------------------------------------
/**Checks if the  address is aligned for ARBURST in  Cache Line Size Transactions */
 svt_err_check_stats cache_line_arburst_wrap_addr_aligned_valid_check;
  //--------------------------------------------------------------
/**Checks if the  address is aligned for AWBURST in  Cache Line Size Transactions */
 svt_err_check_stats cache_line_awburst_incr_addr_aligned_valid_check;
  //--------------------------------------------------------------
/**Checks if the  address is aligned for ARBURST in  Cache Line Size Transactions */
 svt_err_check_stats cache_line_arburst_incr_addr_aligned_valid_check;
  //--------------------------------------------------------------

/**Checks if the  AWDOMAIN is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_awdomain_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  ARDOMAIN is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_ardomain_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWCACHE is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_awcache_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  AWLOCK is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_awlock_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  ARLOCK is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_arlock_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWCACHE is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_arcache_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  AxBAR is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_axbar_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  AxLEN is correctly indicated as per the Cache Line Size configured */
 svt_err_check_stats  cache_line_sz_eq_alen_asize_check ;
  //--------------------------------------------------------------

  /**Checks if CLEANSHARED transaction starts only from INVALID, UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats cleanshared_correct_start_state_check; 
  //--------------------------------------------------------------

  /**Checks if CLEANSHAREDPERSIST transaction starts only from INVALID, UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats cleansharedpersist_correct_start_state_check; 
  //--------------------------------------------------------------

  /**Checks if CLEANINVALID transaction starts only from INVALID state */
  svt_err_check_stats cleaninvalid_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if MAKEINVALID transaction starts only from INVALID state */
  svt_err_check_stats makeinvalid_correct_start_state_check; 
  //--------------------------------------------------------------

  /**Checks if WRITEUNIQUE transaction starts only from INVALID, UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats writeunique_correct_start_state_check; 
  //--------------------------------------------------------------

  /**Checks if WRITELINEUNIQUE transaction starts only from INVALID, UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats writelineunique_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if WRITEBACK transaction starts only from UNIQUEDIRTY or SHAREDDIRTY state */
  svt_err_check_stats writeback_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if WRITECLEAN transaction starts only from UNIQUEDIRTY or SHAREDDIRTY state */
  svt_err_check_stats writeclean_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if WRITEEVICT transaction starts only from UNIQUECLEAN state */
  svt_err_check_stats writeevict_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if EVICT transaction starts only from UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats evict_correct_start_state_check;         
  //--------------------------------------------------------------

  /**Checks if snoop response has data transfer bit set for cacheline in dirty state */
  svt_err_check_stats dirty_state_data_transfer_check;         
  //--------------------------------------------------------------

/**Checks if the  AWDOMAIN is valid for ReadOnce & WriteUnique Transactions */
 svt_err_check_stats  writeunique_awdomain_valid_value_check;
//------------------------------------------------------------------------

/**Checks if the  AWDOMAIN is valid for WriteUniquePtlstash Transactions */
 svt_err_check_stats  writeuniqueptlstash_awdomain_valid_value_check;

  //--------------------------------------------------------------
/**Checks if the  AWDOMAIN is valid for ReadOnce & WriteUnique Transactions */
 svt_err_check_stats  readonce_ardomain_valid_value_check;
  //--------------------------------------------------------------

 /**Checks if all transactions (other than ReadNoSnoop, ReadOnce, ReadOnceCleanInvalid, ReadOnceMakeInvalid, WriteNoSnoop, WriteUnique) are required to be a full cache line size */
 svt_err_check_stats  full_cache_line_size_check;

/**Checks if the  AWBURST is valid for ReadOnce & WriteUnique Transactions */
 svt_err_check_stats writeunique_awburst_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWBURST is valid for writeuniqueptlstash Transactions */
 svt_err_check_stats writeuniqueptlstash_awburst_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  ARBURST is valid for ReadOnce & WriteUnique  Transactions */
 svt_err_check_stats readonce_arburst_valid_value_check;


/**Checks if the  AWCACHE is valid for ReadOnce & WriteUnique  Transactions */
 svt_err_check_stats  writeunique_awcache_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWLOCK is valid for ReadOnce & WriteUnique  Transactions */
 svt_err_check_stats  writeunique_awlock_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWCACHE is valid for writeuniqueptlstash  Transactions */
 svt_err_check_stats  writeuniqueptlstash_awcache_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWLOCK is valid for writeuniqueptlstash  Transactions */
 svt_err_check_stats  writeuniqueptlstash_awlock_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  ARCACHE is valid for ReadOnce & WriteUnique   Transactions */
 svt_err_check_stats  readonce_arcache_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  ARLOCK is valid for ReadOnce & WriteUnique   Transactions */
 svt_err_check_stats  readonce_arlock_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWSIZE is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awsize_valid_value_check;
  //--------------------------------------------------------------


/**Checks if the  AWSIZE is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awlen_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWLEN for INCR is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awburst_awlen_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWLEN for INCR is valid for AXI Transactions */
 svt_err_check_stats awburst_awlen_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWBURST is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awburst_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWDOMAIN is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awdomain_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWCACHE is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awcache_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  Address aligned for WRAP is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awburst_incr_valid_check;
  //--------------------------------------------------------------

/**Checks if the AWSIZE x AWLEN  not exceed the cache line size  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awburst_wrap_valid_check;
//--------------------------------------------------------------

/**Checks if the ALOCK is 0 for WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awlock_valid_value_check;
//--------------------------------------------------------------
/** If a snooped master receives a snoop transaction when it is has an
 * outstanding WriteEvict transaction, then it is the responsibility of the
 * snooped master to ensure that no other master can update the same area of
 * main memory at the same time. The snooped master achieves this by delaying
 * the snoop response until the snooped master has completed the WriteEvict
 * transaction */
 svt_err_check_stats snoop_response_to_same_cacheline_during_writeevict_check;
//--------------------------------------------------------------
/** While a transaction is in progress which has the AWUNIQUE signal asserted,
 * the master must not give a snoop response that would allow another copy of
 * the line to be created, or an agent to consider that it has another Unique
 * copy of the line
 */
 svt_err_check_stats snoop_response_to_same_cacheline_during_xact_with_awunique_check;
//--------------------------------------------------------------
/** AWUNIQUE must be deasserted for WRITECLEAN transactions */
svt_err_check_stats writeclean_awunique_valid_value_check;
//--------------------------------------------------------------
/** AWUNIQUE must be asserted for WRITEEVICT transactions */
svt_err_check_stats writeevict_awunique_valid_value_check;
//--------------------------------------------------------------
/** Monitor check that all byte strobes are asserted for a WRITEEVICT transaction */
svt_err_check_stats writeevict_wstrb_valid_value_check;

//--------------------------------------------------------------
/** Monitor check that all byte strobes are asserted for a WRITELINEUNIQUE transaction */
svt_err_check_stats writelineunique_wstrb_valid_value_check;
//--------------------------------------------------------------

/** Monitor check that all byte strobes are asserted for a writeuniquefullstash transaction */
svt_err_check_stats writeuniquefullstash_wstrb_valid_value_check;
//--------------------------------------------------------------

//--------------------------------------------------------------
/**Checks the valid response of EXOKAY response is only for readnosnoop Transactions */
svt_err_check_stats exokay_resp_observed_only_for_exclusive_transactions_check;
//--------------------------------------------------------------
/**Checks that if cacheline is in invalid state then exclusive load transaction is issued only as READCLEAN or READSHARED */
svt_err_check_stats exclusive_load_from_valid_state_check;
//--------------------------------------------------------------
/**Checks that if cacheline is in invalid state then exclusive store transaction is not issued */
svt_err_check_stats exclusive_store_from_valid_state_check;
//--------------------------------------------------------------
/**Checks that if cacheline is in shared state then exclusive transaction is issued only as CLEANUNIQUE, READCLEAN or READSHARED*/
svt_err_check_stats exclusive_transaction_from_shared_state_check;
//--------------------------------------------------------------
/**Checks for no data transfer occurs for a CleanShared,Cleansharedpersist, CleanInvalid, CleanUnique, MakeUnique, MakeInvalid and Evict Transactions */
svt_err_check_stats perform_no_datatransfer_check;
  //--------------------------------------------------------------
/**Checks the valid response of  cleanshared Transactions */
svt_err_check_stats read_data_chan_cleanshared_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  cleansharedPersist Transactions */
svt_err_check_stats read_data_chan_cleansharedpersist_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of makeinvalid  Transactions */
svt_err_check_stats read_data_chan_makeinvalid_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  makeunique Transactions */
svt_err_check_stats read_data_chan_makeunique_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of cleaninvalid  Transactions */
svt_err_check_stats read_data_chan_cleaninvalid_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  cleanunique Transactions */
svt_err_check_stats read_data_chan_cleanunique_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  readunique Transactions */
svt_err_check_stats read_data_chan_readunique_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  readnotshareddirty Transactions */
svt_err_check_stats read_data_chan_readnotshareddirty_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  readclean Transactions */
svt_err_check_stats read_data_chan_readclean_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of readonce  Transactions */
svt_err_check_stats read_data_chan_readonce_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of readnosnoop  Transactions */
svt_err_check_stats read_data_chan_readnosnoop_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the CLEANUNIQUE, MAKEUNIQUE, CLEANSHARED,
  * CLEANINVALID,CLEANSHAREDPERSIST,
  * MAKEINVALID, READBARRIER, DVMCOMPLETE, DVMMESSAGE transactions
  * have only single read data channel transfer */
svt_err_check_stats coherent_single_read_data_transfer_valid_check;
  //--------------------------------------------------------------

/**Checks the valid response of readbarrier  Transactions */
svt_err_check_stats read_data_chan_readbarrier_resp_valid_check;
  //--------------------------------------------------------------

/**Checks the valid response of DVM Message Transactions */
svt_err_check_stats read_data_chan_dvmmessage_resp_valid_check;
  //--------------------------------------------------------------

/**Checks the valid response of DVM Complete Transactions */
svt_err_check_stats read_data_chan_dvmcomplete_resp_valid_check;

//--------------------------------------------------------------
/**Checks the valid snoop response of DVM Message Transactions */
svt_err_check_stats snoop_chan_dvmsync_resp_valid_check;
  //--------------------------------------------------------------

/**Checks the valid snoop response of DVM Complete Transactions */
svt_err_check_stats snoop_chan_dvmcomplete_resp_valid_check;

//--------------------------------------------------------------
/**Checks the ACSNOOP reserved values */
svt_err_check_stats acsnoop_reserved_value_check ;
 //--------------------------------------------------------------


/**Checks that for MakeInvalid transactions a data transfer is never required */
svt_err_check_stats snoop_resp_passdirty_datatransfer_check;
//--------------------------------------------------------------

/**If DataTransfer is asserted, a full cache line of data must be provided on the snoop data channel */
svt_err_check_stats full_cache_line_datatransfer_check;
//

/**Checks for readunique cleaninvalid makeinvalid illegal response  */
svt_err_check_stats snoop_response_channel_isshared_check;
//--------------------------------------------------------------

/** Checks that CDLAST signal is asserted during the final data transfer.
  *
  * protocol checks : port level 
  */
svt_err_check_stats cdlast_asserted_for_last_snoopread_data_beat;
//--------------------------------------------------------------

/**Checks that the FIXED burst type is not supported for shareable transactions */
svt_err_check_stats fixed_burst_type_valid;
//--------------------------------------------------------------

/**Checks that ACVALID and ACREADY to be asserted before asserting CRVALID */
svt_err_check_stats snoop_addr_snoop_resp_check;
//--------------------------------------------------------------
/**Checks that ACVALID and ACREADY to be asserted before asserting CDVALID */
svt_err_check_stats snoop_addr_snoop_data_check;
//--------------------------------------------------------------

//--------------------------------------------------------------
/**Checks the combinations of ARDOMAIN,ARSNOOP and ARBAR are valid and unreserved */
svt_err_check_stats arsnoop_ardomain_arbar_reserve_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWDOMAIN,AWSNOOP and AWBAR are valid and unreserved */
svt_err_check_stats awsnoop_awdomain_awbar_reserve_value_check;
//--------------------------------------------------------------

//Barrier Checks //
/**Checks the AWADDR is valid for AWBAR  */
svt_err_check_stats write_barrier_awaddr_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations AWBURST and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awburst_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWLEN and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awlen_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWSIZE and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awsize_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWCACHE and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awcache_type_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWSNOOP and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awsnoop_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWLOCK and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awlock_type_valid_value_check;
//--------------------------------------------------------------
/**Checks the valid value of AxUSER for write barrier transactions */
svt_err_check_stats barrier_transaction_user_valid_value_check;
//--------------------------------------------------------------

/**Checks the ARADDR is valid for ARBAR  */
svt_err_check_stats read_barrier_araddr_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations ARBURST and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arburst_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARLEN and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arlen_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARSIZE and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arsize_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARCACHE and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arcache_type_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARSNOOP and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arsnoop_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARLOCK and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arlock_type_valid_value_check;
//--------------------------------------------------------------
/** Checks the Barrier Id valid and unreserved.  */
svt_err_check_stats barrier_id_valid_value_check;
//--------------------------------------------------------------
/**Checks the Read Barrier valid response  */
svt_err_check_stats barrier_read_response_check ;
//--------------------------------------------------------------
/**Checks the Write Barrier valid response  */
svt_err_check_stats barrier_write_response_check ;
//--------------------------------------------------------------
/**Checks that both transactions in a barrier pair must have the same AxID, AxBAR, AxDOMAIN, and AxPROT values*/
svt_err_check_stats barrier_pair_cntrl_signals_check ;
//--------------------------------------------------------------
/**Checks that barrier pairs must be issued in the same sequence on the read address and write address channels*/
svt_err_check_stats barrier_pair_check ;
//--------------------------------------------------------------
/**Checks that ARADDR/AWADDR should always be aligned to Atomicity Size*/
svt_err_check_stats align_addr_atomicity_size_check ;

//--------------------------------------------------------------
/** Checks the RACK for valid response.  */
svt_err_check_stats rack_status_check;
//--------------------------------------------------------------
/** Checks the WACK for valid response.  */
svt_err_check_stats wack_status_check;
//-------------------------------------------------------------
/** Checks all snoop transactions are ordered. .
  */
svt_err_check_stats snoop_transaction_order_check;

//DVM CHECKS //
 /**Checks  For DVM ARBURST 'b01 Burst Type INCR. */
svt_err_check_stats dvm_message_arburst_valid_value_check;
//-------------------------------------------------------------
 /**Checks For DVM  ARLEN All zero */
svt_err_check_stats dvm_message_arlen_valid_value_check;
//-------------------------------------------------------------

 /**Checks for DVM ARSIZE Matches the data bus width */
svt_err_check_stats dvm_message_arsize_valid_value_check;
//-------------------------------------------------------------

 /**Checks for DVM ARCACHE 'b0010 Normal non-cacheable */
svt_err_check_stats dvm_message_arcache_type_valid_value_check;
//-------------------------------------------------------------

 /**Checks for DVM ARLOCK 'b0 Normal Access. */
svt_err_check_stats dvm_message_arlock_type_valid_value_check;
//-------------------------------------------------------------
 
/**Checks for DVM  ARDOMAIN  is Inner shareable or Outer shareable */ 
svt_err_check_stats dvm_message_ardomain_type_valid_value_check;
//-------------------------------------------------------------
/**Checks for DVM  ARBAR[0] is 1'b0 */ 
svt_err_check_stats dvm_message_arbar_valid_value_check;
//-------------------------------------------------------------
/** Checks for DVMCOMPLETE the valid value of  ARSNOOP */ 
svt_err_check_stats dvm_complete_arsnoop_valid_value_check;
//-------------------------------------------------------------
/** Checks for DVMSYNC, DVM Operation the valid value of  ARSNOOP */ 
svt_err_check_stats dvm_operation_dvm_sync_arsnoop_valid_value_check;
//-------------------------------------------------------------
/** Checks for DVMSYNC, DVM Operation the valid value of ARADDR[(n-1):32],[15],[11:0] bits */
svt_err_check_stats dvm_operation_dvm_sync_araddr_valid_value_check;
//-------------------------------------------------------------
/** Checks for DVMHINT, DVM Operation the valid value of ARADDR[15] */
svt_err_check_stats dvm_operation_dvm_hint_araddr_valid_value_check;
//-------------------------------------------------------------

/** Checks the value of  ACSNOOP for the DVM complete */ 
svt_err_check_stats dvm_complete_acsnoop_valid_value_check;
//-------------------------------------------------------------
/** Checks the value of  ACSNOOP for the DVM SYNC */ 
svt_err_check_stats dvm_operation_dvm_sync_acsnoop_valid_value_check;
//-------------------------------------------------------------

/** Checks For a DVM Complete message, ARADDR is defined to be all zeros */
svt_err_check_stats dvmcomplete_araddr_valid_value_check;
//-------------------------------------------------------------
/** Checks  For a DVM Complete message, ACADDR is defined to be all zeros */
svt_err_check_stats dvmcomplete_acaddr_valid_value_check;
//-------------------------------------------------------------


/** Checks  FOR DVM Message the value of reserve address bit should be zero  */
svt_err_check_stats dvmmessage_araddr_reserve_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[11:10] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_hypervisor_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[9:8] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_secure_nonsecure_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[6] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_vmid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[5] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_asid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[0] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[0] of DVM message type Branch Predictor Invalidate */
svt_err_check_stats dvmmessage_branch_predictor_invalidate_supported_message_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[9:8] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_physical_inst_cache_secure_nonsecure_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[6:5] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_physical_inst_cache_vid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[0] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_physical_inst_cache_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[11:10] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_invalidate_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[9:8] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_secure_nonsecure_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[6] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_vmid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[5] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_asid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[0] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_addr_specified_value_check;
//-------------------------------------------------------------


//DVM snoop

/** Checks  FOR DVM Message the value of reserve address bit should be zero  */
svt_err_check_stats dvmmessage_snoop_araddr_reserve_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[11:10] of DVM message type TLB Invalidate    */
svt_err_check_stats snoop_dvmmessage_tlb_hypervisor_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[9:8] of DVM message type TLB Invalidate    */
svt_err_check_stats snoop_dvmmessage_tlb_secure_nonsecure_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[6] of DVM message type TLB Invalidate    */
svt_err_check_stats snoop_dvmmessage_tlb_vmid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[5] of DVM message type TLB Invalidate    */
svt_err_check_stats snoop_dvmmessage_tlb_asid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[0] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_snoop_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[0] of DVM message type Branch Predictor Invalidate */
svt_err_check_stats snoop_dvmmessage_branch_predictor_invalidate_supported_message_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[9:8] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_physical_inst_cache_secure_nonsecure_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[6:5] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_physical_inst_cache_vid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[0] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_physical_inst_cache_snoop_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[11:10] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_virtual_inst_cache_invalidate_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[9:8] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_virtual_inst_cache_secure_nonsecure_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[6] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_virtual_inst_cache_vmid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[5] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_virtual_inst_cache_asid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[0] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_snoop_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks the overlapping AWID of Write Barrier transactions with any active Write transactions */
svt_err_check_stats writebarrier_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks the overlapping ARID of Read Barrier transactions with any active Read transactions */
svt_err_check_stats readbarrier_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks the overlapping ARID of DVM transactions with any active Read transactions */
svt_err_check_stats dvm_xact_id_overlap_check;

/** Checks the overlapping ARID of Non-DVM or Non-Device transactions with any active transactions */
svt_err_check_stats read_non_dvm_non_device_xact_id_overlap_check;

/** Checks the overlapping AWID of Non-DVM or Non-Device transactions with any active transactions*/
svt_err_check_stats write_non_dvm_non_device_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks that all transactions of multi-part DVM operation have same ID */
svt_err_check_stats multipart_dvm_coherent_same_id_check;
//-------------------------------------------------------------
/** Checks that all transactions of multi-part DVM operation have same coherent response */
svt_err_check_stats multipart_dvm_coherent_same_response_check;
//-------------------------------------------------------------
/** Checks that all coherent transactions of multi-part DVM operation are sent in successive manner 
    and no unrelated coherent transaction sent during multi-part DVM opearion over AR channel */
svt_err_check_stats multipart_dvm_coherent_successive_transaction_check;
//-------------------------------------------------------------
/** Checks that all transactions of multi-part DVM operation have same snoop response */
svt_err_check_stats multipart_dvm_snoop_same_response_check;
//-------------------------------------------------------------
/** Checks that all snoop transactions of multi-part DVM operation are sent in successive manner 
    and no unrelated snoop transaction sent during multi-part DVM opearion over AC channel */
svt_err_check_stats multipart_dvm_snoop_successive_transaction_check;
//-------------------------------------------------------------
/** Checks the overlapping ARID of Non-Barrier Non-DVM transactions with any active Barrier/DVM transactions */
svt_err_check_stats readbarrier_dvm_norm_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks the overlapping AWID of Non-Barrier Non-DVM transactions with any active Barrier/DVM transactions */
svt_err_check_stats writebarrier_norm_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks the receiverd RDATACHK is same as the parity calculated from RDATA in a read  transaction */
svt_err_check_stats rdatachk_parity_calculated_rdata_parity_check;
//-------------------------------------------------------------
/** Checks the receiverd parity is same as the parity calculated from respective signal in a transaction */
svt_err_check_stats received_parity_calculated_parity_check;
//-------------------------------------------------------------
/** Checks the receiverd WDATACHK is same as the parity calculated from WDATA in a write transaction */
svt_err_check_stats wdatachk_parity_calculated_wdata_parity_check;
//-------------------------------------------------------------
/** Checks the receiverd CDDATACHK is same as the parity calculated from CDDATA in a snoop transaction */
svt_err_check_stats cddatachk_parity_calculated_cddata_parity_check;
//-------------------------------------------------------------

// Checks on 'Sequencing Transactions'

/** Checks that Master does not receive a snoop transaction until 
  * any preceding transaction to the same cache line has completed
  */
svt_err_check_stats resp_to_same_cache_line_check;
//-------------------------------------------------------------
/** Checks that if received a snoop transaction, response to a transaction 
  * to the same cache line is not received , until snoop response is sent 
  */
svt_err_check_stats snoop_to_same_cache_line_check;
//-------------------------------------------------------------
/**
  * Checks that the if DataTransfer de-asserted then no data transfer will occur on the snoop data channel
  *  for this transaction DataTransfer, CRRESP[0]
  */
svt_err_check_stats cdvalid_high_no_data_transfer_check;
//-------------------------------------------------------------
// START OF LOCKED ACCESS CHECKS
/**
  * Checks that there are no pending transactions before a locked
  * sequence starts
  */
svt_err_check_stats no_pending_xacts_during_locked_xact_sequeunce_check;
//-------------------------------------------------------------

/**
  * Checks that all transactions of locked sequence have the same id
  */
svt_err_check_stats locked_sequeunce_id_check;
//-------------------------------------------------------------

/**
  * Checks that when a master does a lock transaction, it does not target subsequent transactions in the lock 
  * sequence to any slave other than the locked slave
  */

svt_err_check_stats locked_sequence_to_same_slave_check;
 //----------------------------------------------------------------
/**
  * Check that the master follows as per the recommendation from spec to  limit 2 transaction for the lock access
  */
   svt_err_check_stats locked_sequence_length_check;
//-------------------------------------------------------------

/**
  * Checks that there are no pending transactions of a locked sequeunce
  * when a normal transaction is received
  */
svt_err_check_stats no_pending_locked_xacts_before_normal_xacts_check;
// END OF LOCKED ACCESS CHECKS

/** 
  * Checks that AXI master and AXI slave are not exceeding the user 
  * configured maximum number of outstanding transactions (#num_outstanding_xact)
  * If #num_outstanding_xact = -1 then #num_outstanding_xact will not be considered , 
  * instead #num_read_outstanding_xact and #num_write_outstanding_xact will be considered for 
  * read and write transactions respectively.
  */
svt_err_check_stats max_num_outstanding_xacts_check ;

//-------------------------------------------------------------
// START OF PERFORMANCE CHECKS
/**
  * Checks that the latency of a write transaction is not greater than the
  * configured max value
  */
svt_err_check_stats perf_max_write_xact_latency_check;

/**
  * Checks that the latency of a write transaction is not lesser than the
  * configured min value
  */
svt_err_check_stats perf_min_write_xact_latency_check;

/**
  * Checks that the average latency of write transactions in a given interval
  * is not more than the configured max value
  */
svt_err_check_stats perf_avg_max_write_xact_latency_check;

/**
  * Checks that the average latency of write transactions in a given interval
  * is not less than the configured min value
  */
svt_err_check_stats perf_avg_min_write_xact_latency_check;

/**
  * Checks that the latency of a read transaction is not greater than the
  * configured max value
  */
svt_err_check_stats perf_max_read_xact_latency_check;

/**
  * Checks that the latency of a read transaction is not lesser than the
  * configured min value
  */
svt_err_check_stats perf_min_read_xact_latency_check;

/**
  * Checks that the average latency of read transactions in a given interval
  * is not more than the configured max value
  */
svt_err_check_stats perf_avg_max_read_xact_latency_check;

/**
  * Checks that the average latency of read transactions in a given interval
  * is not less than the configured min value
  */
svt_err_check_stats perf_avg_min_read_xact_latency_check;

/**
  * Checks that the throughput of read transactions in a given interval is
  * not more that the configured max value
  */
svt_err_check_stats perf_max_read_throughput_check;

/**
  * Checks that the throughput of read transactions in a given interval is
  * not less that the configured min value
  */
svt_err_check_stats perf_min_read_throughput_check;

/**
  * Checks that the throughput of write transactions in a given interval is
  * not more that the configured max value
  */
svt_err_check_stats perf_max_write_throughput_check;

/**
  * Checks that the throughput of write transactions in a given interval is
  * not less that the configured min value
  */
svt_err_check_stats perf_min_write_throughput_check;

/**
  * Checks that the bandwidth of read transactions in a given interval is
  * not more that the configured max value
  */
svt_err_check_stats perf_max_read_bandwidth_check;

/**
  * Checks that the bandwidth of read transactions in a given interval is
  * not less that the configured min value
  */
svt_err_check_stats perf_min_read_bandwidth_check;

/**
  * Checks that the bandwidth of write transactions in a given interval is
  * not more that the configured max value
  */
svt_err_check_stats perf_max_write_bandwidth_check;

/**
  * Checks that the bandwidth of write transactions in a given interval is
  * not less that the configured min value
  */
svt_err_check_stats perf_min_write_bandwidth_check;

// END OF PERFORMANCE CHECKS
//-------------------------------------------------------------
// START Of STREAM CHECKS

svt_err_check_stats signal_valid_tvalid_check;

/** Checks that TREADY is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tready_when_tvalid_high_check;

/** If tdata is enabled, checks that TDATA is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tdata_when_tvalid_high_check;

/** If tstrb is enabled, checks that TSTRB is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tstrb_when_tvalid_high_check;

/** If tkeep is enabled, checks that TKEEP is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tkeep_when_tvalid_high_check;

/** If tlast is enabled, checks that TLAST is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tlast_when_tvalid_high_check;

/** If tid is enabled, checks that TID is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tid_when_tvalid_high_check;

/** If tuser is enabled, checks that TUSER is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tuser_when_tvalid_high_check;

/** If tdest is enabled, checks that TDEST is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tdest_when_tvalid_high_check;

/** 
  * Checks that TDATA is stable when TVALID is high 
  * When svt_axi_port_configuration::check_valid_data_bytes_only_enable=1 ,
  * it considers only valid byte lanes of tdata based on tstrb. 
  * When svt_axi_port_configuration::check_valid_data_bytes_only_enable=0 ,
  * whole tdata as seen on the bus will be considered.
  */
svt_err_check_stats signal_stable_tdata_when_tvalid_high_check;

/** Checks that TSTRB is stable when TVALID is high */
svt_err_check_stats signal_stable_tstrb_when_tvalid_high_check;

/** Checks that TKEEP is stable when TVALID is high */
svt_err_check_stats signal_stable_tkeep_when_tvalid_high_check;

/** Checks that TLAST is stable when TVALID is high */
svt_err_check_stats signal_stable_tlast_when_tvalid_high_check;

/** Checks that TID is stable when TVALID is high */
svt_err_check_stats signal_stable_tid_when_tvalid_high_check;

/** Checks that TUSER is stable when TVALID is high */
svt_err_check_stats signal_stable_tuser_when_tvalid_high_check;

/** Checks that TDEST is stable when TVALID is high */
svt_err_check_stats signal_stable_tdest_when_tvalid_high_check;

/** Checks that TVALID is low when reset is active */
svt_err_check_stats tvalid_low_when_reset_is_active_check;

/** Checks if tvalid was interrupted before tready got asserted */
svt_err_check_stats tvalid_interrupted_check;

/** Checks that TSTRB is low if TKEEP is low */
svt_err_check_stats tstrb_low_when_tkeep_low_check;

/** Checks that received data stream is not interleaved beyond stream_interleave_depth
  * value. An error is issued if data stream is interleaved beyond this value. */
svt_err_check_stats stream_interleave_depth_check;

/** Checks that the burst length of received data stream is not exceeding the maximum
  * value allowed for stream_burst_length defined by `SVT_AXI_MAX_STREAM_BURST_LENGTH. */
svt_err_check_stats max_stream_burst_length_exceeded_check;

/** 
 * @groupname port_interleaving_check
 * @check_description   
 * - Checks if address does fall to correct interleaved port.
 * - Valid when port cfg port_interleaving_enable = 1.   
 * .
 * @end_check_description
 *
 * @check_pass
 * address does fall to correct interleaved port. 
 * @end_check_pass
 *
 * @check_fail
 * address does not fall to correct interleaved port. 
 * @end_check_fail
 *
 * @applicable_device_type
 * master & slave 
 * @end_applicable_device_type
 *
 * @check_additional_information
 * @end_check_additional_information   
 */
svt_err_check_stats port_interleaving_check;

/** 
 * @groupname trace_tag_validity_check
 * @check_description   
 * - Trace tag value on data channel or resposne channel should be valid as per the trace tag 
 * - value on the address channel. 
 * .
 * @end_check_description
 *
 * @check_pass
 * For Write transactions the check will pass if:
 * A slave that receives a write request with AWTRACE asserted should assert the BTRACE signal alongside
 * the write response.
 * For Read transactions the check will pass if:
 * A slave that receives a read request with the ARTRACE signal asserted should assert the RTRACE signal
 * alongside every beat of the read response.
 * For Snoop transactions the check will pass if:
 * A master that receives a snoop request with the ACTRACE signal asserted should assert the CRTRACE
 * signal alongside the snoop response.The master should also assert CDTRACE alongside every data beat of
 * the snoop data that is associated with the snoop transaction.
 * @end_check_pass
 * @check_fail
 * If trace_tag in the request packet is set to 1 and in the spawned response or data packet is set 
 * to 0.
 * @end_check_fail
 *
 * @applicable_device_type
 * @end_applicable_device_type
 *
 * @check_additional_information
 * @end_check_additional_information   
 */
svt_err_check_stats trace_tag_validity_check;


// END OF STREAM CHECKS
//-------------------------------------------------------------
  `ifdef SVT_AXI_QVN_ENABLE
// START OF QVN CHECKS    

/** Checks that VARVALIDVN* is not X or Z */
svt_err_check_stats signal_valid_varvalidvnx_check;

/** Checks the VARQOSVN* is valid when VARVALIDVN* is high */
svt_err_check_stats  signal_valid_varqosvnx_when_varvalidvnx_high_check;  
   
/** Checks that VARREADYVN* is not X or Z */
svt_err_check_stats signal_valid_varreadyvnx_check;

/** Checks that VAWVALIDVN* is not X or Z */
svt_err_check_stats signal_valid_vawvalidvnx_check;

/** Checks the VAWQOSVN* is valid when VAWVALIDVN* is high */
svt_err_check_stats  signal_valid_vawqosvnx_when_vawvalidvnx_high_check;  
   
/** Checks that VAWREADYVN* is not X or Z */
svt_err_check_stats signal_valid_vawreadyvnx_check;
   
/** Checks that VWVALIDVN* is not X or Z */
svt_err_check_stats signal_valid_vwvalidvnx_check;

/** Checks that VWREADYVN* is not X or Z */
svt_err_check_stats signal_valid_vwreadyvnx_check;
   
/** Checks that VARVALIDVN* when asserted, remains asserted till VARREADYVN* */   
svt_err_check_stats varvalidvn_deassertion_check;
   
/** When a master sets VARVALIDVNx high, it can change VARQOSVNx proir to the slave granting a token, but only if the value increase. */
svt_err_check_stats varqosvn_valid_change_check;

/** Checks that VAWVALIDVN* when asserted, remains asserted till VAWREADYVN* */   
svt_err_check_stats vawvalidvn_deassertion_check;
   
/** When a master sets VAWVALIDVNx high, it can change VAWQOSVNx proir to the slave granting a token, but only if the value increase. */
svt_err_check_stats vawqosvn_valid_change_check;
   
/** Checks that VWVALIDVN* when asserted, remains asserted till VWREADYVN* */   
svt_err_check_stats vwvalidvn_deassertion_check;

/** Check that master must only set ARVNET to values that correspond to a VN where the associated set of token request signals exist.*/
svt_err_check_stats arvnet_for_existing_vn_check;
   
/** Check that master must only set AWVNET to values that correspond to a VN where the associated set of token request signals exist.*/
svt_err_check_stats awvnet_for_existing_vn_check;

/** Check that master must only set WVNET to values that correspond to a VN where the associated set of token request signals exist.*/
svt_err_check_stats wvnet_for_existing_vn_check;

/** Check that master must have read address token for VN denote ARVNET, before it can send read address channel transfer (Except for a Barrier transaction).*/
svt_err_check_stats rd_addr_chan_vn_token_availability_check;
   
/** Check that master must have write address token for VN denote AWVNET, before it can send write address channel transfer (Except for a Barrier transaction).*/
svt_err_check_stats wr_addr_chan_vn_token_availability_check;
   
/** Check that master must have write data token for VN denote WVNET, before it can send a data beat. */
svt_err_check_stats wr_data_chan_vn_token_availability_check;

/** Check that transaction with the same AXI ID that are are sent on the same physical link must use the same VN.*/
svt_err_check_stats same_axi_id_over_single_vn_check;

/** Check Before entering a low-power or reset state, the component must have the same number of pre-allocated tokens that it had when it exited reset.*/
svt_err_check_stats pre_allocated_token_count_at_rst_check;

/** Check QVN token handshake signal are not asserted on unsupported VN.*/
svt_err_check_stats qvn_sig_asrt_on_unsupported_vn_check;

/** Check that slave component is not granting more outstanding token than its configured.*/
svt_err_check_stats slave_max_outstanding_token_check;
   
/** Check that token requested should be granted in a bounded time*/
svt_err_check_stats qvn_token_request_timeout_check;
   
//-------------------------------------------------------------
// END OF QVN CHECKS    
`endif

`ifdef SVT_ACE5_ENABLE

//--------------------------------------------------------------
/** Checks that ARCHUNKEN is not X or Z when ARVALID is high */
svt_err_check_stats signal_valid_archunken_when_arvalid_high_check;

//--------------------------------------------------------------
/** Checks that RCHUNKV is not X or Z when RVALID is high */
svt_err_check_stats signal_valid_rchunkv_when_rvalid_high_check;
  
/** Checks that RCHUNKNUM is not X or Z when RVALID and RCHUNKV are high */
svt_err_check_stats signal_valid_rchunknum_when_rvalid_rchunkv_high_check;

/** Checks that RCHUNKSTRB is not X or Z when RVALID and RCHUNKV are high */
svt_err_check_stats signal_valid_rchunkstrb_when_rvalid_rchunkv_high_check;


//--------------------------------------------------------------
/** Checks that ARCHUNKEN is stable when ARVALID is high */
svt_err_check_stats signal_stable_archunken_when_arvalid_high_check;

//--------------------------------------------------------------
/** Checks that RCHUNKV is stable when RVALID is high */
svt_err_check_stats signal_stable_rchunkv_when_rvalid_high_check;

/** Checks that RCHUNKNUM is stable when RVALID and RCHUNKV are high */
svt_err_check_stats signal_stable_rchunknum_when_rvalid_rchunkv_high_check;

/** Checks that RCHUNKSTRB is stable when RVALID and RCHUNKV are high */
svt_err_check_stats signal_stable_rchunkstrb_when_rvalid_rchunkv_high_check;


//--------------------------------------------------------------
/** Checks that ARSIZE is equal to the data bus width or ARLEN is one beat and
 * ARSIZE is 128 bits or larger for rdata chunking */
svt_err_check_stats rdata_chunking_arsize_valid_value_check;

/** Checks that ARADDR is aligned to 16 bytes for rdata chunking */
svt_err_check_stats rdata_chunking_araddr_aligned_check; 

/** Checks that ARBURST is INCR or WRAP for rdata chunking */
svt_err_check_stats rdata_chunking_arburst_type_check;

/**Checks that ARSNOOP is ReadNoSnoop, ReadOnce, ReadOnceCleanInvalid or 
 * ReadOnceMakeInvalid for rdata chunking */
svt_err_check_stats rdata_chunking_arsnoop_valid_value_check;

/** Checks that ARIDUNQ must be asserted for rdata chunking */
svt_err_check_stats rdata_chunking_aridunq_valid_value_check;

//--------------------------------------------------------------  
/**Checks that RCHUNKV is deasserted for all the transfers when ARCHUNKEN is
 * deasserted */
svt_err_check_stats rdata_chunking_rchunkv_zero_when_archunken_deasserted_check;

/**Checks that RCHUNKV must be the same for every response beat of a 
 * transaction */ 
svt_err_check_stats rdata_chunking_rchunkv_same_for_all_response_check;

/** Checks that RCHUNKNUM must be between zero and ARLEN when RVALID and
 * RCHUNKV are high*/
svt_err_check_stats rdata_chunking_rchunknum_valid_value_check;

/**Checks that RCHUNKSTRB must not be zero when RVALID and RCHUNKV are high */
svt_err_check_stats rdata_chunking_rchunkstrb_valid_value_check;

/**Checks that the number of bytes that are transferred through read data
 * chunking must be consistant with ARSIZE and ARLEN */
svt_err_check_stats rdata_chunking_num_bytes_transfer_check;

`endif

`ifdef SVT_UVM_TECHNOLOGY
  /** UVM report server passed in through the constructor */
  uvm_report_object reporter;
`elsif SVT_OVM_TECHNOLOGY
  /** OVM report server passed in through the constructor */
  ovm_report_object reporter;
`else
  /** VMM message service passed in through the constructor*/ 
  vmm_log  log;
`endif

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   */
  extern function new (string name, svt_axi_port_configuration cfg, uvm_report_object reporter, bit register_enable=1, bit enable_pc_cov = 1);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param reporter OVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   */
  extern function new (string name, svt_axi_port_configuration cfg, ovm_report_object reporter, bit register_enable=1, bit enable_pc_cov = 1);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param log VMM log instance used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (string name, svt_axi_port_configuration cfg, vmm_log log = null, bit register_enable=1, bit enable_pc_cov = 1);
`endif
  /** @cond PRIVATE */
  extern function void perform_excl_write_addr_chan_signal_level_checks(svt_axi_transaction xact, 
                       svt_axi_transaction excl_xact, output bit is_excl_wr_error);
 
  extern function void perform_read_addr_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_arid,
                                                       ref logic[`SVT_AXI_MAX_ADDR_WIDTH-1:0] observed_araddr,
                                                       ref logic[`SVT_AXI_MAX_BURST_LENGTH_WIDTH-1:0] observed_arlen,
                                                       ref logic[`SVT_AXI_SIZE_WIDTH-1:0] observed_arsize,
                                                       ref logic[`SVT_AXI_BURST_WIDTH-1:0] observed_arburst,
                                                       ref logic[`SVT_AXI_LOCK_WIDTH-1:0] observed_arlock,
                                                       ref logic[`SVT_AXI_CACHE_WIDTH-1:0] observed_arcache,
                                                       ref logic[`SVT_AXI_PROT_WIDTH-1:0] observed_arprot,
                                                       ref logic[`SVT_AXI_QOS_WIDTH-1:0] observed_arqos,
                                                       ref logic[`SVT_AXI_REGION_WIDTH-1:0] observed_arregion,
                                                       ref logic[`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] observed_aruser,
                                                       ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_ardomain,
                                                       ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop,
                                                       ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar,
                                                       ref logic observed_arready,
`ifdef SVT_ACE5_ENABLE
                                                       ref logic[`SVT_AXI_MAX_MMUSID_WIDTH-1:0]observed_stream_id,
                                                       ref logic[`SVT_AXI_MAX_MMUSSID_WIDTH-1:0]observed_sub_stream_id,
                                                       ref logic observed_secure_or_non_secure_stream,
                                                       ref logic observed_sub_stream_id_valid,
                                                       ref logic observed_addr_translated_from_pcie,
                                                       ref logic observed_aridunq, 
                                                       ref logic observed_archunken,
                                                       ref logic [`SVT_AXI_MAX_MPAM_WIDTH-1:0] observed_armpam,
                                                       output bit is_aridunq_valid, 
                                                       output bit is_archunken_valid,
                                                       output bit is_stream_id_valid,                              
                                                       output bit is_sub_stream_id_valid,                          
                                                       output bit is_secure_or_non_secure_stream_valid,                              
                                                       output bit is_sub_streamid_valid,                          
                                                       output bit is_addr_translated_from_pcie_valid,
                                                       output bit is_armpam_valid,     
 `endif
                                                       output bit is_arid_valid,
                                                       output bit is_araddr_valid,
                                                       output bit is_arlen_valid,
                                                       output bit is_arsize_valid,
                                                       output bit is_arburst_valid,
                                                       output bit is_arlock_valid,
                                                       output bit is_arcache_valid,
                                                       output bit is_arprot_valid,
                                                       output bit is_arqos_valid,
                                                       output bit is_arregion_valid,
                                                       output bit is_aruser_valid,
                                                       output bit is_ardomain_valid,
                                                       output bit is_arsnoop_valid,
                                                       output bit is_arbar_valid,
                                                       output bit is_arready_valid,
                                                       output bit excl_read_error
                                                     );
  extern function void perform_read_data_chan_signal_level_checks(
                                                      ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_rid,
                                                      ref logic[`SVT_AXI_RESP_WIDTH-1:0] observed_rresp,
                                                      ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] observed_rdata,
                                                      ref logic[`SVT_AXI_MAX_POISON_WIDTH-1:0] observed_rpoison,
                                                      ref logic observed_rlast,
                                                      ref logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] observed_ruser,
                                                      ref logic observed_rready,
 `ifdef SVT_ACE5_ENABLE
                                                      ref logic observed_ridunq, 
                                                      ref logic observed_rchunkv,
                                                      ref logic [`SVT_AXI_MAX_CHUNK_NUM_WIDTH-1:0] observed_rchunknum,
                                                      ref logic [`SVT_AXI_MAX_CHUNK_STROBE_WIDTH-1:0] observed_rchunkstrb,
                                                      output bit is_ridunq_valid, 
                                                      output bit is_rchunkv_valid,
                                                      output bit is_rchunknum_valid,
                                                      output bit is_rchunkstrb_valid,
 `endif
                                                      output bit is_rid_valid,
                                                      output bit is_rresp_valid,
                                                      output bit is_rdata_valid,
                                                      output bit is_rpoison_valid,
                                                      output bit is_rlast_valid,
                                                      output bit is_ruser_valid,
                                                      output bit is_rready_valid
                                                    );
  extern function void perform_write_addr_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_awid,
                                                       ref logic[`SVT_AXI_MAX_ADDR_WIDTH-1:0] observed_awaddr,
                                                       ref logic[`SVT_AXI_MAX_BURST_LENGTH_WIDTH-1:0] observed_awlen,
                                                       ref logic[`SVT_AXI_SIZE_WIDTH-1:0] observed_awsize,
                                                       ref logic[`SVT_AXI_BURST_WIDTH-1:0] observed_awburst,
                                                       ref logic[`SVT_AXI_LOCK_WIDTH-1:0] observed_awlock,
                                                       ref logic[`SVT_AXI_CACHE_WIDTH-1:0] observed_awcache,
                                                       ref logic[`SVT_AXI_PROT_WIDTH-1:0] observed_awprot,
                                                       ref logic[`SVT_AXI_QOS_WIDTH-1:0] observed_awqos,
                                                       ref logic[`SVT_AXI_REGION_WIDTH-1:0] observed_awregion,
                                                       ref logic[`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] observed_awuser,
                                                       ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_awdomain,
                                                       ref logic[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] observed_awsnoop,
                                                       ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_awbar,
`ifdef SVT_ACE5_ENABLE
                                                       ref logic[`SVT_AXI_STASH_NID_WIDTH-1:0]observed_stash_nid,
                                                       ref logic[`SVT_AXI_STASH_LPID_WIDTH-1:0]observed_stash_lpid,
                                                       ref logic observed_stash_nid_valid,
                                                       ref logic observed_stash_lpid_valid,
                                                       output bit is_stash_nid_valid,                              
                                                       output bit is_stash_lpid_valid,                          
                                                       output bit is_stashnid_valid,                              
                                                       output bit is_stashlpid_valid,                          
                                                       ref logic[`SVT_AXI_MAX_MMUSID_WIDTH-1:0]observed_stream_id,
                                                       ref logic[`SVT_AXI_MAX_MMUSSID_WIDTH-1:0]observed_sub_stream_id,
                                                       ref logic observed_secure_or_non_secure_stream,
                                                       ref logic observed_sub_stream_id_valid,
                                                       ref logic observed_addr_translated_from_pcie,
                                                       ref logic [`SVT_ACE5_ATOMIC_TYPE_WIDTH-1:0] observed_awatop,
                                                       ref logic [`SVT_AXI_MAX_MPAM_WIDTH-1:0] observed_awmpam,
                                                       output bit is_stream_id_valid,                              
                                                       output bit is_sub_stream_id_valid,                          
                                                       output bit is_secure_or_non_secure_stream_valid,                              
                                                       output bit is_sub_streamid_valid,                          
                                                       output bit is_addr_translated_from_pcie_valid,                          
                                                       output bit is_awatop_valid,
                                                       ref logic observed_awidunq,
                                                       output bit is_awidunq_valid,
                                                       output bit is_awmpam_valid,
`endif
                                                       ref logic observed_awready,
                                                       ref logic observed_awunique,
                                                       output bit is_awid_valid,
                                                       output bit is_awaddr_valid,
                                                       output bit is_awlen_valid,
                                                       output bit is_awsize_valid,
                                                       output bit is_awburst_valid,
                                                       output bit is_awlock_valid,
                                                       output bit is_awcache_valid,
                                                       output bit is_awprot_valid,
                                                       output bit is_awqos_valid,
                                                       output bit is_awregion_valid,
                                                       output bit is_awuser_valid,
                                                       output bit is_awdomain_valid,
                                                       output bit is_awsnoop_valid,
                                                       output bit is_awbar_valid,
                                                       output bit is_awready_valid,
                                                       output bit excl_write_error,
                                                       output bit is_awunique_valid
                                                     );
  extern function void perform_write_data_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_wid,
                                                       ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] observed_wdata,
                                                       ref logic[(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] observed_wdatachk,
                                                       ref logic[`SVT_AXI_MAX_POISON_WIDTH-1:0] observed_wpoison,
                                                       ref logic[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] observed_wstrb,
                                                       ref logic observed_wlast,
                                                       ref logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] observed_wuser,
                                                       ref logic observed_wready,
                                                       output bit is_wid_valid,
                                                       output bit is_wdata_valid,
                                                       output bit is_wdatachk_valid,
                                                       output bit is_wpoison_valid,
                                                       output bit is_wstrb_valid,
                                                       output bit is_wlast_valid,
                                                       output bit is_wuser_valid,
                                                       output bit is_wready_valid
                                                     );
  extern function void perform_write_resp_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_bid,
                                                       ref logic[`SVT_AXI_RESP_WIDTH-1:0] observed_bresp,
                                                       ref logic[`SVT_AXI_MAX_BRESP_USER_WIDTH-1:0] observed_buser,
                                                       ref logic observed_bready,
 `ifdef SVT_ACE5_ENABLE
                                                       ref logic observed_bidunq, 
                                                       output bit is_bidunq_valid, 
 `endif
                                                       output bit is_bid_valid,
                                                       output bit is_bresp_valid,
                                                       output bit is_buser_valid,
                                                       output bit is_bready_valid
                                                     );
  extern function void perform_data_stream_signal_level_checks(ref logic observed_tready,
                                                        logic[`SVT_AXI_MAX_TDATA_WIDTH-1:0] observed_tdata,
                                                        logic[`SVT_AXI_TSTRB_WIDTH-1:0] observed_tstrb,
                                                        logic[`SVT_AXI_TKEEP_WIDTH-1:0] observed_tkeep,
                                                        logic observed_tlast,
                                                        logic[`SVT_AXI_MAX_TID_WIDTH-1:0] observed_tid,
                                                        logic[`SVT_AXI_MAX_TDEST_WIDTH-1:0] observed_tdest,
                                                        logic[`SVT_AXI_MAX_TUSER_WIDTH-1:0] observed_tuser,
                                                        output bit is_tready_valid,
                                                        output bit is_tdata_valid,
                                                        output bit is_tstrb_valid,
                                                        output bit is_tkeep_valid,
                                                        output bit is_tlast_valid,
                                                        output bit is_tid_valid,
                                                        output bit is_tdest_valid,
                                                        output bit is_tuser_valid);

  extern function void perform_slave_reset_checks(logic observed_rvalid, logic observed_bvalid);
  extern function void perform_master_reset_checks(logic observed_arvalid, logic observed_awvalid, logic observed_wvalid);
  extern function void perform_master_reset_ace_checks(logic observed_crvalid, logic observed_cdvalid);
  extern function void perform_slave_reset_ace_checks(logic observed_acvalid);
  extern function void perform_master_reset_stream_checks(logic observed_tvalid);
  /** Performs checks on AWUNIQUE signal for WRITECLEAN and WRITEEVICT transactions */
  extern function void perform_awunique_checks(logic observed_awunique, svt_axi_transaction xact);
  /**
    * Performs check on WRITEEVICT transaction that all wstrb signals must be asserted
    * @param xact Transaction on which check is to be done
    * @param check_all_beats Indicates if check is to be done on current beat or on all beats
    */
  extern function void perform_coherent_xact_wstrb_check(svt_axi_transaction xact, bit check_all_beats);
  extern function void reset_internal_variables();

  extern function void perform_burst_4k_boundary_cross_check  (svt_axi_transaction xact);
  extern function void perform_burst_wrap_address_align_check (svt_axi_transaction xact);
  extern function void perform_burst_wrap_burst_length_check  (svt_axi_transaction xact);
  extern function void perform_burst_size_not_exceed_data_width_check(svt_axi_transaction xact);
  extern function void perform_write_burst_value_check  (ref logic observed_awvalid, ref logic[`SVT_AXI_BURST_WIDTH-1:0] observed_awburst);
  extern function void perform_write_valid_awcache_check(ref logic observed_awvalid,input svt_axi_transaction xact);
  extern function void perform_read_burst_value_check  (ref logic observed_arvalid, ref logic[`SVT_AXI_BURST_WIDTH-1:0] observed_arburwst);
  extern function void perform_read_valid_arcache_check(ref logic observed_arvalid, input svt_axi_transaction xact);
  extern function void perform_write_resp_write_data_check(svt_axi_transaction xact);
  extern function void perform_write_resp_write_address_check(svt_axi_transaction xact);

  extern function void perform_snoop_addr_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_ACE_SNOOP_ADDR_WIDTH-1:0] observed_acaddr,
                                                       ref logic[`SVT_AXI_ACE_SNOOP_TYPE_WIDTH-1:0] observed_acsnoop,
                                                       ref logic[`SVT_AXI_ACE_SNOOP_PROT_WIDTH-1:0] observed_acprot,
                                                       ref logic observed_acready,
                                                       output bit is_acaddr_valid,
                                                       output bit is_acsnoop_valid,
                                                       output bit is_acprot_valid,
                                                       output bit is_acready_valid
                                                     );
  extern function void perform_snoop_data_chan_signal_level_checks(
                                                      ref logic[`SVT_AXI_ACE_SNOOP_DATA_WIDTH-1:0] observed_cddata,
                                                      ref logic[(`SVT_AXI_ACE_SNOOP_DATA_WIDTH/8)-1:0] observed_cddatachk,
                                                      ref logic[`SVT_AXI_ACE_SNOOP_POISON_WIDTH-1:0] observed_cdpoison,
                                                      ref logic observed_cdlast,
                                                      ref logic observed_cdready,
                                                      output bit is_cddata_valid,
                                                      output bit is_cddatachk_valid,
                                                      output bit is_cdpoison_valid,
                                                      output bit is_cdlast_valid,
                                                      output bit is_cdready_valid
                                                    );
  extern function void perform_snoop_resp_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_ACE_SNOOP_RESP_WIDTH-1:0] observed_crresp,
                                                       ref logic observed_crready,
                                                       output bit is_crresp_valid,
                                                       output bit is_crready_valid
                                                     );
  extern function void perform_axcache_axdomain_restriction_check(svt_axi_transaction xact);
  extern function void perform_axcache_axdomain_invalid_value_check(svt_axi_transaction xact);
  extern function void perform_cache_line_size_transaction_constraint_check(svt_axi_transaction xact);
  extern function void perform_readonce_writeunique_transaction_check(svt_axi_transaction xact);
  extern function void perform_writeback_writeclean_transaction_check(svt_axi_transaction xact);
  extern function void perform_axi_transaction_check(svt_axi_transaction xact);
  extern function void perform_read_data_channel_signal_value_check(svt_axi_transaction xact);
  extern function void perform_write_response_channel_signal_value_check(svt_axi_transaction xact,ref logic[`SVT_AXI_RESP_WIDTH-1:0] observed_bresp);
  extern function void perform_dvm_snoop_response_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_acsnoop_reserved_value_check(ref logic [`SVT_AXI_ACE_SNOOP_TYPE_WIDTH-1:0] observed_acsnoop);
  extern function void perform_snoop_resp_passdirty_datatransfer_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_full_cache_line_datatransfer_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_cdvalid_high_no_data_transfer_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_snoop_response_channel_isshared_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_fixed_burst_type_valid_check(svt_axi_transaction xact);
  extern function void perform_snoop_addr_snoop_resp_check(svt_axi_snoop_transaction snoop_xact );
  extern function void perform_snoop_addr_snoop_data_check(svt_axi_snoop_transaction snoop_xact );

  extern function void perform_arsnoop_ardomain_arbar_reserve_value_check(ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop, 
  ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_ardomain, 
  ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar);

  extern function void perform_awsnoop_awdomain_awbar_reserve_value_check(ref logic[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] observed_awsnoop,
                                                                          ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_awdomain,
                                                                          ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_awbar);

//--- Barrier Checks --//
  extern function void perform_write_barrier_transaction_check (svt_axi_transaction xact,ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_awbar,
                                                                 ref logic[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] observed_awsnoop);
  extern function void  perform_read_barrier_transaction_check(svt_axi_transaction xact,ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar,
ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop);
  extern function void perform_barrier_id_check(svt_axi_transaction xact);
  extern function void perform_barrier_read_response_check(svt_axi_transaction xact, ref logic[1:0]  observed_rresp ,ref logic observed_rlast);
  extern function void perform_barrier_write_response_check(svt_axi_transaction xact, ref logic[1:0] observed_bresp);
  extern function void perform_rack_status_check(svt_axi_transaction xact, logic observed_ack );
  extern function void perform_wack_status_check(svt_axi_transaction xact, logic observed_ack );


//--- DVM Checks --//

  extern function void  perform_dvm_read_address_channel_check(svt_axi_transaction xact,ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar,
                                                       ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop,
                                                       ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_ardomain);

  extern function void  perform_dvm_arsnoop_read_address_channel_valid_check(svt_axi_transaction xact,
                                                                     ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop,
                                                                     ref logic[`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0] observed_araddr);
  extern function void  perform_dvm_acsnoop_snoop_address_channel_valid_check(svt_axi_snoop_transaction xact,
                                                                      ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_acsnoop,
                                                                      ref logic[`SVT_AXI_ACE_SNOOP_ADDR_WIDTH-1 : 0] observed_acaddr);
  extern function void perform_dvmcomplete_araddr_valid_value_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_araddr_reserve_value_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_tlb_invalidate_supported_message_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_branch_predictor_invalidate_supported_message_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_physical_inst_cache_invalidate_supported_message_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_virtual_inst_cache_invalidate_supported_message_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_snoop_araddr_reserve_value_check(svt_axi_snoop_transaction xact);
  extern function void perform_dvmcomplete_acaddr_valid_value_check(svt_axi_snoop_transaction xact);
  extern function void perform_snoop_dvmmessage_tlb_invalidate_supported_message_check(svt_axi_snoop_transaction xact);
  extern function void perform_snoop_dvmmessage_branch_predictor_invalidate_supported_message_check(svt_axi_snoop_transaction xact);
  extern function void perform_snoop_dvmmessage_physical_inst_cache_invalidate_supported_message_check(svt_axi_snoop_transaction xact);
  extern function void perform_snoop_dvmmessage_virtual_inst_cache_invalidate_supported_message_check(svt_axi_snoop_transaction xact);
  extern function svt_axi_transaction perform_barrier_dvm_normal_xact_id_overlap_check(svt_axi_transaction xact, svt_axi_transaction active_queue[$], bit execute_check=1);
  extern function void perform_barrier_pair_check(svt_axi_transaction xact);
  extern function void perform_atomicity_size_alignment_check(svt_axi_transaction xact);

`ifdef SVT_ACE5_ENABLE
//--- UNIQUE_ID - OUTSTANDING Checks --//
  extern function svt_axi_transaction perform_no_unique_id_outstanding_transaction_with_same_id(svt_axi_transaction xact, svt_axi_transaction active_queue[$]);
`endif 

//--- NON - DVM Checks --//
  extern function svt_axi_transaction perform_non_dvm_non_device_with_overlap_id_check(svt_axi_transaction xact, svt_axi_transaction active_queue[$]);

  `ifdef SVT_AXI_QVN_ENABLE
//--- QVN Checks --//   
  extern function void perform_qvn_wr_addr_token_handshake_checks(logic       observed_vawvalidvnx,
                  logic       observed_vawreadyvnx,
                  logic [3:0] observed_vawqosvnx,
                  logic [3:0] vnet_id);
   
  extern function void perform_qvn_wr_data_token_handshake_checks(logic       observed_vwvalidvnx,
                  logic       observed_vwreadyvnx,
                  logic [3:0] vnet_id);

  extern function void perform_qvn_wr_addr_chan_sig_assertion_on_unsupported_vn_check(logic       observed_vawvalidvnx,
                          logic     observed_vawreadyvnx,
                          logic [3:0] vnet_id);

  extern function void perform_qvn_wr_data_chan_sig_assertion_on_unsupported_vn_check(logic     observed_vwvalidvnx,
                          logic     observed_vwreadyvnx,
                          logic [3:0] vnet_id);

   extern function void perform_qvn_rd_addr_token_handshake_checks(logic       observed_varvalidvnx,
                   logic       observed_varreadyvnx,
                   logic [3:0] observed_varqosvnx,
                   logic [3:0] vnet_id);
   
   extern function void perform_qvn_rd_addr_chan_sig_assertion_on_unsupported_vn_check(logic       observed_varvalidvnx,
                           logic     observed_varreadyvnx,
                           logic [3:0] vnet_id);
  `endif
  extern function void set_default_pass_effect(svt_err_check_stats::fail_effect_enum default_pass_effect);
  extern function void execute(svt_err_check_stats check_stats, bit test_pass, string fail_msg="",
                               svt_err_check_stats::fail_effect_enum fail_effect=svt_err_check_stats::ERROR);

  extern function void register_err_checks(bit en = 1'b1);

  extern function void passive_cache_check_post_coherent(coherency_error_type_enum err_status, svt_axi_transaction xact, svt_axi_passive_cache_line::passive_state_enum initial_state);

  extern virtual function void passive_cache_check_post_snoop(coherency_error_type_enum err_status, svt_axi_snoop_transaction xact, svt_axi_passive_cache_line::passive_state_enum initial_state);

  extern virtual function void perform_multipart_dvm_coherent_start_check(svt_axi_transaction xact, bit drop_xact_if_error=0);

  extern virtual function void perform_multipart_dvm_coherent_response_check(svt_axi_transaction xact);

  extern virtual function void perform_multipart_dvm_snoop_start_check(svt_axi_snoop_transaction xact);

  extern virtual function void perform_multipart_dvm_snoop_response_check(svt_axi_snoop_transaction xact);

  extern virtual function void update_checks_on_reset(svt_axi_transaction xact = null);

  extern virtual function bit is_current_xact_multipart_dvm(svt_axi_transaction xact);
  extern virtual function bit is_snoop_xact_multipart_dvm(svt_axi_snoop_transaction xact);

  /** 
    * This task waits for the last transaction of a multipart DVM. 
    */
  extern task check_and_wait_for_last_multipart_coherent_dvm_xact();

  /** Returns 1 if only the first part of a multi-part dvm is received */
  extern function bit is_second_part_of_multipart_pending();

  extern virtual function void disable_ace_checks();

  extern virtual function void reset_multipart_dvm();

  extern virtual function void reset_barrier_checks();

`ifdef SVT_ACE5_ENABLE
  // E1.11.1 (IHI0022H) Constraints for rdata chunking for AXI Transaction
  extern virtual function void perform_rdata_chunking_check(svt_axi_transaction xact);
  extern virtual function void perform_rdata_chunking_num_bytes_transfer_check(svt_axi_transaction xact, logic observed_rchunkv, logic observed_rlast);
`endif
/** @endcond */

endclass

//----------------------------------------------------------------
/**
AXI  port monitor check description
*/

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
kaL0BWBflkZOlB4qhfltIVItI50H1EqrVbbFymPy/W+GrU31dR59rA/zllpg0cVQ
1S3nyldP3h6sBPVelALPeousJUOHfZQ9cj7QhVNWoUOqZaplDfio7QYin5wgTZU+
uaZNWcZi+A4tGE2YGG7/lA5hXt/z4OzpKyi+aWNaTlKYcTYWAe8t6g==
//pragma protect end_key_block
//pragma protect digest_block
5jvpVfgAxCPwExXLojT1kFSvsa4=
//pragma protect end_digest_block
//pragma protect data_block
47eHQ0J1Rel9vVroo53aHrt1CYDBHSZ6GjDoKVkXmVB36594IUyf0VizRsRJcluR
PhJ7VGmma3O9qpdkwvV1q1jwLFIXP8b3BVywDsxqI54Kpe56YQmda7SqRq/VbGqA
/2DiRdOfwzixhD00zHAqWysenreVxnE7vRvjtSE9DYzs+sbcMt1uTKLcuddB/qIN
rwhRpQedwRGOeaHx8rOgpuvrrU38mc7yK9MftadvaHaRf8PWMwyPu0BNZNua4pdC
E2Di/4Kl/++mrELNRZH2LUaio8ZvDIKHnvA5KxTxuyBbacs/TbE+1YP0gIhTlcVo
WiQYwvvDxMKsqRgbgT1SA0ndnBY8qGBejy1iirEzT8zOP7ZHEnP0OCEIRW6xQsaM
wAas6x+u7u+JmZwCuP7pQr3Ax8jS3isdvI94MnMkXUJAhHsDun3Pac+hgiBRT8hs
0ygpRAXiOppW2ZDYmHYeguE/myZZfGXGvDpCiiWHnG0jw+VqaI+wL5xuF9B4Oz4u
CjlfQMqhbPxITr2gXNMps4sHnQjwsTTwn3O8WSM7Nb4iErUD6ht3LeaBXqCiQhk2
6UP8XEdz+OUlev9NNYaU9zRSuCJY2J80h4+l/IOCPTEPOpL/IiEGfZtTpv0V/XsR
uZe9NH9AhDNvizNKXaW2h2i1zsGlBR5bglRGsSbX0jFaZZbQPzkNpLLuTt7xec47
1UbogmFYueZIEyUMNb9rW3GcfdR02Hfh+h7PDsj+UeSdLoIABNB7NQhW4ymkehZK
gB/0xSn9zuKQ0wTWUuiJpekUJ0qgrqFwf+o2I+L1zhkuuWuas0qr9pzRI0k8b+pk
bpSmWILm7fs4Li0Ik3QL/xvT1OcQiG5zaoy2I5SIJNPQ/oo/a+7V/Y0HHb2KrhjE
aY8+44agwtDMu4Y6crjjSix4XaEDGcG/Se+zxxyOr+bd7O5v7gTGroQT4SYnnoMg
Zd8EiiWU9TenbjDvu0YMJiNTXw6ZGEjV9+G0Qd/My0nadcK4++Kd+phreQrGBqRj
h6H8uIpOKnWAUwbF0JuGigJZUIkHnuuDuA9zD+MsyAzakzjlE78pSD2HYw+wK5xG
Mlmtmmd1UWoe0ydVTFdpvdirXmCiw9mD/jmULxIMv/ebRaQynRu0NdoFxBN+8iQ/
lkMVmWkxQijxCB0Jou/CkdVhqtDNfaia5kV9Ou33Yzr8gjWeaXMgH9JkAPDMClnG
TWOb5bAkRggLPTjOAiESqyfQj003tl8v7NVNENrVk+5UvgJcHt/7b2EDflTtBjOI
veX/jbLuYIPLXWuW4MFWNIYBAiKFHHVVRs1L88nix1loH96mSqOeCCpC1VUSFRTS
eOPFCZd37+l0/hcwjbfIDBlm1pClmUFWIMrHj5IuCTvSo/1t4T6YKPENOqPJ7y7U
4SeVDPWjWcRvmnvrPo4BSnNbRfDgtKHTQeuThuxHf9rSVo5kg52QGGrIrOlxcAbo
n8nfQX6TqGtnDKmhrDufKRxz0MasL975YbkZg6DVv+rtKFfb7dD+l0F1oDBy7Fj+
wkPZXT3thbegi0qr31SRLN1Znpkp6RebmckfGRT9/Xz8VB/hYmwOKU+fKyIzrmMi
HMcvTIrs7nxLKVw9VRk8wWOLmOJjowrKN8I+WynqXFKqOLhUlCTWdGSsnqXCJ9Es
IaXByrtNcQ3X8U0V/7p2fI7rVBO2fgVDwHsE1DG2US5W9Wzdbd4T9hf9EXJRLBts
8CYtYvTAVP/cGuM1MtFwK793OcwAWwbJ2FjofzZhgLfMaQMQK2OIlZasn57e5lDP
HwEV5B8YoSorxhYV+NLmvVE8UzedYLYshSGWLwH6ZrwI9jzAunDbQeCRsyX+5gd4
sI1imHBvZVQ/O5c8lAjRfHASU41H3LQiLVy1SHk/ZTmFFeGl49bjcVHbbnRXzIa3
+tz1tKbkFZ36KatdiAnIK0c40cN+INI6OTPKPH55GlsvAYHRTNDfJX1QgqLrFpTv
0/8PRLDWryBrN22n40SBh5NztbI94gvOzAgr/D82D6fHnYTt3UOwRqPIU0+r7MC/
7KPkGfT84yyq2cWxkwSYoYsPoqRElqL3H0c0QPYCgpX1slZEJG38mS6ETaq7T1wg
wAWDyJ5cQhkGP9e4JpE+mrDwErClz6+la/lQS+8LHRoHRMSmf6pVewRWDTXxxqbt
H/pyf4QxKiEkkhAQOc7D1dAWg3sdiJMu2VVEzA/TEQKqXF2FrhxTT69M+q0wSYG2
svM9MTWwBV2la0V6ByNO+TSWW69T5+Cvuz+nc9pYstKTUwLy5UHyf3tIwt8uoGKQ
cUkp0Ricrtm4k7s9ebHOMyVOqUd46tkzbxT6i5T0K7lTcWv3SvOPbCNrMP+PR+7e
RwgdqRqDY6v2c2w690wr4iP53Ze0d3XTRRfzvmZLTA/cJtqb1n8utonJIZOUPUkt
IYKsCGFfkpabL6ObU/tdFbcTV6obA0FW2kAvJbQoZZ1EvxIj2wHIsDXHEmxMRem9
VFl7MHF05wv56Fw/mB08rvk1qVcaqyB/Yt+9WtoeJjXCNS6IYsY8kqNI1F/HMFIy
FWbWWja4nscIMWlkqxWdbmiDH1WK/Zxvgb8Xei6UaTqyR0V706E+WogFGRDfKRNT
qZsnyx67aReSKyQiS0r/p0cv+rTH1Rypbfd5ZvMf+NJHfxXX/XTlk+C9hj1R/RI+
BN747sMLLlL+MyukLlfTs8kvj3aKUQz+ML4K3OQ/4ssvBYzxp8y9gY8yAbPT+CHa
6dmtIiUA4u18dVCgTfpq1L5L3oyEZgdeDw9wMdy00B1bPjpynhuLdlXQeTwlrD/Z
9acnw7V+UeSlyUql4pJoASfwvXLCdO47OWqih5jMxvKfbEF1lyeMVpYbWvXMm7qv
aLYSBdSuaWNZ5gWmSeGfvdKe8n7bsOVy/U4GfYmuR4dlW4j+T6jaLW3dJFL6q/fC
kARpjIc6x/+WZBd853pGttg9uydJZixQq/sFqgW2CVBwmbu8SNgzaSZW768ot7zA
ZwZ7vgBgPUuOdB4DrzmQSOvBjaseOhWeO7aZRuKs4MMMg61yIIHZz10lA7k2NR1G
qiXR+r1RkZ1KXltgsBMM4OtgO5iS4Ifae+xaWlwWzwWoGcR0hl7xdMvFemlC0haT
WvsinBVJl/4v1zp+1uLiFbMm6PcJDjmGyXdx1Ooe6zwkuRLt84w0RK5tgIeWu+de
Asxogim4btBOv3D8YlJDyFe91fGH2YN/cTrRxUtwDFAzUIrcOtNrmMPrF6+gAFBe
K2JIkblppjCxr42pY5iG0zeo4tKv9QuY5eHj3vrBZErgX978Jo1zvr3sn1L2sHWC
PrA8jAU+P0OWIaS2g5ydj8wPFTISQ5bnKCrsOBBX39HfmgZgUYXYnkWp4H0M9q6e
eqpLPTh6mtVB3wZ4w22rPuhRRDrn9G31F/PGpjTrJdwCmiVcVhh6ChB859J3SJlT
qR0vFOmlQcfeiEpbuoFWY0YXVrZXxPMvDhV0v7mHOh9jD0Dk0pBx9ktemRDC6F37
hNTJm4H9KniyADo7M4EZWE24Wu1AmorPK++dMhGkmILv1G2as5w1M7ijz0BcDcW+
P4qu+1Bmw3CoXKii1SrY+dGF+WoZ9MWUEZE2p1I8ig1H7z6mYdMXtVc1ruTug9GU
exOj0wWbMrJNq2oKS6G5AjS3LcWIVLaDPldhfr4Xj87NRTL7hD+Nf83AozzYgodi
F6bg6fjGkVXNpo1KDrGXW6DSSQJCSR47JKkDVLUafr7s3RzywaftIBDLone5bhlm
Jkf+JBigv2fTfqvpkmcfJ9blVAJ6wYtaLSSBTFGjpd1J4RGVS6Ei9Qo9/8n/UeMu
tdFbY36l7ra0BB5Zh6vkYksm252MBMpvMd81CMPdBUNIV+xDaoOx7WKLRxhg9u0a
wNrO2gzHrsKKcTfDbFHf6KuhUu2wPijOnu+JghwyyBBqhFx1LveyUGnssSBRyqTx
eTLuv1ImV7CBjQ4jkyEFtVQdpsSCnfCtPlWkSeYPG5HHznKA0nt2iTHSKvBgYH/2
fKruKkvtmcf8z/Shs76+oPaVp/bPi6zL3ie/UkuHoQNDUrZIIgdpmUEUZmqWZdc0
SzCN0czoQx06RYw+GKH2Q5QCVKsdmqYFPRZfQFHVgWBpui3J9sETlavwheAqEuZL
AJqO8VAFGyptlpxb6T7YTyKRcrq4TEnKc4I8jOQh8o+qxgQ1/lM31oIIL96WN7QX
ADafrZLsAwgvbfHug6YrMWf/4AgUkoeSC9/TGGjoDhvDcsugD9c+LZqEJyyefV5r
4YhcEbZ5kzITG6lrA+MItL7oZ5GF9zNUdY9MPFClBFOl5oRGlQV1tRmembMpqY4r
y8idOAaZvPQcka2jzNkW/fLB+9Hf2l+GH8NQ2nwU824fSsZHjQTn9pogfn6uQdiL
VN7zHfKWj4UO++uFtXXvuSfPyrwGbtCkb5SCe1ZoZL4i+p4Bm6ZkIiZseYupeaEw
Ef+xvTE63ndYekhM4kvaAUWql3vRmKSZ7GCxXf17yQFWsRvnxzUwTsuyNFUWKbj3
/mE3JECLM1VVYmXWhu9HW9zgtjYgL5zj6pv2Qz0/tlBZQEtceB7HLnD48Nk4faPA
Egl4Y1tet2thQMOIMncp+P4J/nqTid4BlJ+8m7ehopurJxSg4F1izrMpyk+q4kuA
8II/3MgL7taoILaMgWPKvEVhXP1hwqZCsWydjm6UnIZkag3WhaTGNzH1S2xBoi3C
MgeqDIWwOHJy4r2xyTO/Tt8weVrljwKI82G0wlxfZRnLMGRx5c8YD9khty2yeYjJ
i9DjO5u/ATL2qXpwOqVGPhla4eb/E0JMS3+LMKqFtOzU3ga96ZyR3e4IkzZ/RzBB
BGwx/YK7b65kDF1mhJFI9XPSh10AoqzJjqq+N1yXSOZnDv3f68lkD5LDI0VzA+BW
d6qguvEUMg8xoZMm5nbHzg271eI5WHKi+XAKaz1jPR3x6mygZQDPDoog0RhGC3f4
ylHvlteMZG0r9h1uq4hh6AfW3ZjlnTE6MBOkr8s907th0l2et2ZfIPr8/BC1ZgSu
rKnK/tUlOSRoQNtFVVjqUNT5ez9cpJ2vWwc8kvBM3Gz9N5Zp1oofkI10jqgRuPuD
xQvugiWtfZsW+sTnQF01O34lR2VjjTcR2pZde8g6jWy5WjUoT99WnuYHbdYDP687
yD3EZqX+ZW8iUpY318+ibVUgGsPwZNiIgWBrLbB8w61DyVYZaz/FU/gzcAHCTtXt
EY7HOxy//+71yJPoIStf279KSIDOGLVjcBX6sCwAcnkWuxK9eN6CWHpeNeAjWxwl
BS3z89C1t90xE/qzLvv7mCqtIz3QPD8/sWL3affSnWqUhmdF/58BIvairw74nenv
UBVDD8hz2FbHFog/mwhNRABsue3TvjJVJsl+s5T9U3cz23TKWZGA99eIpXI8brzS
++D8rWkAoX0W+piBRX9apboHF+V0hsdqHz+Ej8iSzyD9ELiVbO1VNfgUCcqA2qhc
hdsHHgYDe4cM3YQ/xZ9R6j7yj9NS+zAxnBPf6GSEUiFG/fYTiWbsy9Oq08ktpDvV
jdn6RVYACgOPi7D6V0IHVBrrP+bmqYbbQaYRDBpeGsqz3x8EoH4G/fu42bfkSyeY
DFKbQd7BgrJsbU9Rws1CjyE2DdbLA+LU6G/43Dsf5VkrDeiLWLVOrI8nCl2nBTCp
a5XKqmtvPBsJxOt1Jee0Q93h7cG/bnDqn7qoVBWDnOnSITgUb6WbSBeg1IjeFsIY
Y2fa7LakKxB+dQzWSM1X96nWFz65gg9/NWtbgje5lZWNifcC1kcp0PM03y+N3kUS
XzUUebEAMWrnafYDzQPB73or/tTNqQd0beFLYDiSWVTaWplrbJGZ03rg5AAuTT5p
sYmGV8rji1KJkcsbCBdjUSB8FxuqgPj1P6An8bJvF1mu3zMnNOJG6xj1qIsAKLj8
salJAYf4x3SOrzoQTeRmDVNs1U76U4bKpgjYfM7e3QvHfib77BulMfG8uxNlmlHQ
Iwf54T9o8F1KC/FGFSJhIQgTCN9RyhXAn+kIdFO6Uyp04YDaYMFFDvBJC56Jp57D
09uEmAP/ZVcnKmyuJbfR08T+t3wh5a3azGzZfkAivtzFsFtrxCIPt0k9yW0PNonB
efIEau5m9TCsa94fd9vvQLVIGmt/B5sHkBtDJy1JD9f6eodeY7rBEc2uNe4DsdDT
EHiIZk6eo5bPrRQQ2aij8nMJnDe5TTJcuQYnHck/AG2sC94X4TZVsdrErfCYHZ5n
QHylV65o3FqKjZWk23woyKWswEjxMH1tnmiuZjyV0XZcyoYPUGlNRU7JRlx9dxaL
ztoKJNw8CcwCqaqsQCwxO3eWnsfkuUMfoNF17ItUuMOChqQdQArhdI+40SPq0Ip1
dJYFnK3F/cKi1z4dDJq/J6Sh19+Cqs0A1GveytDpVl2E/9wIFjmqkpuUp2mNXH+G
wJrcTxQiLEFkWFt/RQXOVo0teCFy/1kgB5YVrgLqJzeM/fehMNM+psc/5eHr8Efl
ItUFaqT5w5Dpuzt5+nibO1/xnVJjllNhe8F2clh0EuBwx+jHW6eIaLatGoLd26wo
XPdHVzBg6OpifuMnJWLyGt4PbxMBE7pOZEY6D7ANPTZTR0U1uaLUD+6nr8EjYiPd
C47t8lu8X8F5F5vRWB3vYzfpu/qWg+lKnC6qyaXG3ck+9LzJrxCNhDZM5jcHOMWT
STKjnGAxK39jFyXjwN68Q0BVBLT8tqlysn2lRYxStdk8QAF0cFMvIKppUnPFIvJB
gIX67BBFvxDHKWuBXm5T3fwreVpmB3L2L68Yd4QQUWz6UDsc1/CxX6/e6AlSxkkO
4/GMUwluuXBetX99npKOlybGry+IFS1Ghv7H7yql/S7Svxu7Zt3cc3NI+lTlWpPg
srgbKynpMSTd5hFVfrY9b37J4oWCw4aIQf0cgOlPgCd9qJnWgTN6pVRe5f/cWvJu
RRm/vFVrrPC3Kms6qZEAOVm7GOtSBuk299brVQpLROjxUKVG0LVqv9irDBwabfIT
v/OYYjxYdWe6C4FNgzvtQg2ij4Um0GKBvwTLF2/7TDrO2DtzwKD6Rq8s1xshAjmA
V1FYF7NvnplPbDu0nCDma65lvJFLigkLCwxoo6A9dB2j++K6fJ+8X0D9g1Kn1GHJ
yWV1z+imXzgltteWO+UQcDdrWc9AloDfTV0nZIFiZ4DXcXTSnk56WCrXKktpWmnl
anpssEDj/3QQrly9J3+y2VAAstUDa2AtkojshXchNSZXUYwdJQbaub1fe1snBuKi
wezs1e5RfPOt2sk0Tfqldb+T5tUfjxSFn3bZyRV8rJTnP7EitQePglwzoXSdZktQ
DUWgRk2jK3IlVdlikFbz2WJ2T4tJmCV47dD5G9L0ahxn+x3m2HPNqRIIv/DbNaJj
q1CJfatoVbuwblzBWgq6mPgGZjeG55IwaDbEYVLucw4xlWHCfBlYe+nEUy8u93iQ
rA2NydmuhD+hnjM1FxoHI8Sr0SAho68n+uibAx2rZJMh/Qb5g9tqNDoYO209FASD
OOUwfB/RXdHUMCHKgtmURZ/UXo2jQbjMz6K7x2GAVDBBh2TJBAe50IOg1/yuSoit
F3JlRxqpPL9p7qLmtpXPwVJolvPX5guYv792VZr0HFa3Mb1eOQ7JxAD8vG6uskmB
0Kvtk4egCxE89YCw3H1SSqJzFmlSpM4RZSjWk9z9zTy7nGpREYpQ7NIYCWLPYTK8
ZYLvdd4GUxSJm8MxQRyH2CsOrsgR8rEzsquI9O8asJA3nFGqFjUvz0/kez0u+zp/
lZPRvStntaLiKP/rssKv2o+2NFaK/pu24xtY90mFzSFZFDblBHrQFTGU8ochZcNc
Y18x6QEOpjLeAAk4i9JCs7b1QDOryOHxbYqGcNWa1hHfDF+34++H6X8tJUH3DPw0
kGXJG00PM5ar3LJCPmS4N7LwADNtWRYp4iIi5ym0fo/S94NzTIwUJqkiFp02pad4
fsKWbv5VlCiiKDQVuiAboUieQpo5m1G+VLHw2XYN8QNfM7pUL0f6sdU4UTV5CyB5
6VCAmW/xl+g7Mgy/y3aCImLxEu7HDKxZ83Kua2FERpLperF/W5oVEnFXS1KJuZbP
/dcP1u0cSoikCsP71aENCUbmawyMvHprDlxWwt1IlmRY2ZLlwXCuY25s7Lesjiq3
JgDUtdnl5s6dPib1peopclyDdGm/5MlrslTaOuB+f3I8zL98R6ieMd+OIlEV+YnM
pxv4DtA46Eq5/o1dZcab3thwiPRrfS0pWpXLZwFp0Ki5FNE8iC4bIS4ShiCvVqEL
tSvhtwZsTAWa3O78hBBFy4iJegmf9G5z39ts0y+aR9WLYc7AA3oK7A9hVkSIoIwL
U73yMgNHo2TJn7AXfqhASjf5zcQN6SME+FN6rnYtiskihs4taxVHtuelVz9X0NTL
KCZ+uG3V6j+4k7SXOSpb0SY3UgdkRCygBk8XQJZi0U55fZPtLNdS96EqmW/4oYLM
16f/P4c0rsGT174vssQ4FQAD1q1AqKkuBgAwk+rJT/f5EuS747TXjaX4y1b+nUEU
HLevzMmh9aWWOCqdG/b43pEfZuflxUugspn9fzf7VFBGMQfH/ElrCVg6uL7f0a8k
Xrbk8ol0CJHP2UhagJJYZDIZ8OdsfrMguf7PQxnAEpZ4tzmbyfLgQi8IhtmBquMy
aAH2kKX5hpIiSw4yBL2Gbzc/0gK8LXsm3Cnz1Dj1TCypeB5DD1uE2sOVSGA7xhak
s5VwPZIZRA5IQFV+GULt9be/2+KGIuV+ZiD8qspVgjzi7sEB8dThVMNbL1so73QH
ouUOJUGBURGhzWhykHaCecSi096PwuXYUGxz86G+lzS4lJuS66+PRmjUlgyCNskl
40AvnT6ClmXaqhIVOMS8F2MNYK00WvXXQBFXQxvOh+L6611luA+T9xvbpI744Seh
FFxwcPk6PbD4wZMbcXXhiRuAogR97YpbWK7m2WGKEBQg5z4EuNYTArM26HKa5zQB
jcxXAa6DR0MvFCc8mXWuZctDKaSXd+fZNpoWmE1fG7Th+jRyBdBFXnxwYxWvya60

//pragma protect end_data_block
//pragma protect digest_block
vJxMPOuWIzZygEr9K4jPFs5DGRE=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
LeZMclF2wSSwYlDBGD0PxJEUut1rnarzDVxXpbWAljRnF16peArqgBqhU4n0Cmkj
M46gBxf1n0unfBCK+V6qEQXCx1yJK9BVO7nx/aTvpeFRDLPCgGacSGnYNb6TKERu
WUpFxJTzVqLGHrVSDcdExMDUxxpaaAd6z/ptGo5Uwcn6pDRtxHvsQg==
//pragma protect end_key_block
//pragma protect digest_block
pDZ3InyhK10/4Zkk+ayOYUhuZME=
//pragma protect end_digest_block
//pragma protect data_block
eSzpRfj5/fccdph12gGEuCoavb13nAw/Bm78sa8z9uQeHFD/SNf27CbkVsmF+XxT
VCqoS6njjy4Qe3kjazgzpCwkq8OqvplxhI49Rdct/98J9qbL7JzWDM12/ERfkmQJ
OWXbzkjpWCy5TFolCMukmXjQuyNu+93cgxUDnDfMAFWJdpsARpysWT1xo+8MA8O/
Aw6fkMmqIWAc9KHojq+mw5uCKH5nuVA1+7oMRepJwLxWcc1siX20AOkIMUggD7Fh
BzbXK1LKX4rfEOhYeIXRKR7j3BGTl3x2UXf1rMdyANBxanpbZ4OkT54GD4BcwpDF
Cxh83pRNEriuxi85BKyFb9IqIZ/LubaPp5QseFq7HCD3YSpjNfqnjmz97s45QO4A
2A+Fs9ac/kRRVPjggYlr9/qX9c28CvpaCUWU2H66bRWhNenWwmTsUm5g27uPYuml
wyIBfp6rrW792388t0jo2/yfotKilnfddQ0AG1DXAEoQ8y7JZBmOFwhuF/JeXHuc
ABGtB+mtAHLuF8doIpjvaD3iTVZj5MLTYILr/OlleyKTnbsHDNU3r6zJOLZvY8wB
6OlhhnXoMVc5ni9N694Ewm+pwiqE5PxRRzkvCKUTGU3usDRQgfx4+424aZycvXbG
JGpfn5wY6k6PcSmOv/866d+fBixXxT5zAqi3XJgrQf1uBmeJ5c/+071sM6xUiTFP
vz0y4iQhwQq4dA+SHNzJsMnels/mMm2LJwij18NowBmbVJWGPG5MRfG3G7CeAqWs
r2KTYI1jkV/Z8j6zSJfA/80YQSxBBZ3FFDLyW6CrQNNdUm6x7FKh7E4hz8f20OV6
KMZvk/3XBLCGxRmNa/eBuCcoqpJBKo5GkM8gsvovu/wvTERqsmZhQhn1wHSyf/y2
5mzYrZ/WOMJCu/cl6wFXFWqgFkZGzPUZ05dmxStCzk7CRaekjb0owU361SpT77gt
MF/0+Hf3CHyrIpyFvcrznZrbdQllz4hkwLkOO+VC9IU0MgVhR5Dj2M91I5bAFIHY
bsP+S2Is75pB+E4Hc3XtGGdKAnrsDQsBBlabtz2pjOJyUndABvVLjDqRTa2oT2l1
chpr6hsScqQWM3WG4Pwo1YbpI2Cbm6JPM4Uypl53I/zIkI1TW6UcK1lU6xYnOngl
MTm0zNQcOxg7GbOnZVVZU1KEzQpsm0ZZG7R5QiAZeMShsZ/njXNxPQEhRkKwDQL9
70Q5dmIyxRFUQmbVtgBCi746fmOpi7LBoTnOYfRM0GR4xQJrH7K90fRMT0iqB+Vs
DMbEIqCVpm99XHBaxE1P5eU+Ru5Nz3hthvvL5ExcMIK3etd19l6XxQqn7sMbcH3Y
vx/pY44W0SG2NAB6Mp9flx2bezUgqW8+7QIm4P2Re+vr5f+FURC+t/4pOpLCu0uh
+drbHWaV160rkinX7MJD8Kg7PxsOqL5xZp4tRV/b0OJd2gduxNHhVjoEqfJcdVBG
DdZyTc9vULuhK4kHia1lTQuYFENMYY/Gvx3JP63/vYMQ21GHix9qyiuyx0r7um2r
PCwWL033u7jN2yIwYKgo1PvYYD4W6gI202dwqqxqlVpiJzTqPedQw8xnwe9r0sdn
2OAp8WYZGPpoAxEsbUI6oghL+r4sJR/as2mVbAKwAJLAuVY8vlNUKVPcYTwgy+6B
hHbnT9RYhSlrX64n50uz3AkeIQL16pAR91rFFD1CY5Gds9RMQElzrpuC0DgBdSQj
XRq8f1njgEPlQe4Cy8XC0BiK1aK22EFA6FSNMvNjG2bANeDzqtsjgr+tPZY8ccKG
rA7/4fllWCQcJf5qKpG/122UeRfpZykjIECjeKQqepQhy5Dv786kMWQDbPVvgIpR
XtB7GHiwnpJCx4SizXwtz13UPtBAFMlckliiD6Kbra9HW57cb5WEmeyQaTFrDkxo
97cKJ0D+ywef3JgU/MqKGuPTOS9A+KlnmLlzSS9nx8qyQlxNJocU6fBAV3JVQoDK
w7Cd4tR+4uGr9tDjBeyHec6dqNjbGGizqCWidi10EGj30dMSdYwSuez+MaVW05kX
NVHcmKMq9JA+KMCVVP+nD2SETePKGJ0vsVUg6N71wTW2t3Qf8z+lXOQ0P4aPqrRZ
yp+nnwgLryHuYZJ78GYjDa0vItCxFTloKYWR4zKg0fGXVQn3K4vh5g1XlDROdcaU
xXyaC/wfeQzFEvX6djCEZtEWyLSjZG0WOzzxcP6Arr6dIubd7PB75Kyyf4RLR+A1
3IMjaL1tErX9asrA+cR2jqxRrddr/CRaz6Ttuhy/dX2jjHRE5dNPNOfi9q4q5pz7
E5gw9NKqOsqakU5DRwWOw7VvVb6pefnlncWjc+Nh1T5hzew0p2FgTEqnyk1/s3fe
MrdEP5XbxqyWEaTK/zrXzipHUynMnJcnLJ2PuFnaDTt1v0Sf8AeRmJvBU5UtgXX3
s+7JQM9KDtP+jcz5cUAIdGz6nZXopGSbbvFMhNcmTfnM+BZ7oZssXpVTKu4UqnG2
a0UUBJK1t1aGbxKYhS7kq0u75RCYpJtfGlHG2LNPe8mdz36H5YTQMGJ8yE7MwipI
4YD3SS2uA1uCGPB0s93klvTOQ/Tu8alABjDj/+bHzDqDI46/vlABHnz3+roAXXUy
6nFy0pWtfDpmusmzjeoZD/cc93Y08lKERbkfjHH/sG5J5QHlnPmznk39fMuZnPCR
r1zxQw/pdHW5BcynfOFCgMhzfwtVbnosw5AHB4j/M0ZrGchVC8nymLibqckmydKe
MrlC/+7uRlHyqGJCe7lCEQ+QVLtN0J0ztsAvRd9Id3Ak/Yk75lVWLvnRqMQVrvmW
tyNB9X7KNCu58r7tf838Dil2uYFJIpdetTYsQkhfSAiQYOtw/KT/Tl1foPLRILO6
T73siNV7tPKg+H+GxcjfPhNkW25IR52s14I31MzP0OZhf65C+VJf6Yqifji3jvel
jo17IGdOTD4WV0RDILgD4MVb2ycceZ5PdXmYbZeoapmKvaE3ET+4O60XSBWI5JJV
Z3rrUCO0CnGzAceM++o1C/rnjFe+360RTR1oo1Jsna0xARYx16YG0cqqtApV+LL8
bC8czKsNB2h/vUI8bH4+D6l/YUWg+46TNCx6ifjVkBdQvGxYGey8MeAnkF0tw9l1
+JRAcBYUqLq8Jj7kLTraAHdp/hYdnp/A6APX4595L9/yPGoizwViFXtgLsGGjzK1
8sdqMLGd6JzUBbHi5XL9NG2lIL0Bmmd8fK45Sbl+qXEpPJOOaGcy1lMfOCksqOEY
DBC9uBNTtn8vFrgbmWfBRD33Zj7WHdUlsa/gJg4Q3xVQZbR/Xt6AW+06+Vqk9KzP
tNS3amsYE7h/CoZgVoLNdajw9vlazJP3BLd8LJWdjPLZhuykR+jStY+f1E4zIvCi
FHWo/ka1u9vxcXHS767AUGEy8hJdB3sqzIdhStdLnodqD3oeqoblESLhhMOz2pOW
ICgL4HVs9Ms5l/esfQcVzqwLBHQi38VP0KmqV972hwdBKsL1rxG3cvx01LCYv8AW
go5zS72yGAx2LmlnzLiMXNGxfWbIcR0hhZ/+BZGpZ2omjppdUf4Q8oVFdgNRJJgt
ZSz/Vq5oY/oXm53U0qIUrLgSulNJqKTurB8gYq1zNTRGxDagA4x92Ya6ffLmuvcM
5adS0p83K1UF5xlGHvLWfyfCONrBE7zL5NAE5JQdxNjycBRhPI7hJ6bDf2ONU9df
6FaS0DVqzXXTwSvmvpS6XARVKtu1hc2dZc5nL8gvv+XFY1LmEKZEXDZ1m9Wg3nrj
rscAYcI+HODvLE+f2jb4Bi8og40U3F6geUZlX1cStI2Ag7ZhM+yTFAgJtRl7mGMD
rUaOE3KMOZmqiYtRswOJEzP5eMsH/pCL6NSuUzwMbs8J6CWUSWB8WJYXhW4dRmyy
ad/hGOpYj3oDh4iKOmPkAMXiWeB+vIW5zsZrIMZp/7mGDjUZjxD4vSXNjTLszpRa
ebgIiuvNZWm3e+AjDPLvHTzA9jZlnRA1958XjAMpu8zHBDFMdx1S/ACIHkBqlqFt
dSBefhQ3HSKRuELZrsFYRICOCld/3A86rzAwbt3h+TYRSzyqbklK3Vstu4duasBl
iTHix2jlb8DgqtF13sKJ0Z1N7yWEyoCbPNfWdMZUwXOLTJ9eRHIZuGFugG16of58
Ou21QHxKMgyynDOWf/1/59AOVck15k99/Jk5ZcIo9vMYT4iUIsH8bpO32m4/h25Y
3g+jjQ54jCz1m7pAFjZplAShcuiZq20+/i+Bg8pfQg5a9RveqJq4auFBDX6aGavi
FME9C16nGcltGcqkf+gvxgIJNhlfjgiA/ReJHe/EiXphbtemWfRjaHPzvGpETW45
f/IMDutpu2uiQ7vYfUPz5PpiNfIlvAnePK2Obs45alooBk7J05RupIJPxtQyXJgL
0EdlENBE+KRHKuuuTuTT2SDJJSaQAanPuOdlu3dJlm7T3uHVu5ID+x48mSyiFO1x
XOqDjX7xkwJ3OHfmh25UQe4Ed6OXCu43KlWOtvYY8Ex80FKi292g7+Gr+Mpr8vfF
rNnukgR+D3o92ZsveaBXA8XUVvCNlglz/Ql9idzdFY41XJmRhN1VpOQgufWanLN3
eqFB3rx/MHU86t2IZ3ASgpdid5qcDw2OZywn1qk67xonIX86iVrBxXXn+YRWwuDi
sPOiuGEHYkBL4/Lw38MXnrYVl/r7Rze1aOLeHhpveE87v08TQORkco1gBxD9cecp
Kl5Bmwi3bg05O35sHsmQk3mB4IhcCn8mBlpG9pFUus78L5B+D+armXOWomlnycJj
ZRuGrixlIWBMBSJQioCzVNUNUIDfW+8sURo8CbrzCGAXSkEjxEX4XBsULoJEX1wc
JF1MU9sLSL/Bv55PY7Zfwb+MU68i46q5NMJPQPrxRZQI6E7X0I3Dh9bpF9MBpR+l
HOykl9vB2ExNJqMzCPdFN4mm/pzEzivh1jut2/87LSXVUWtxEeITpxIdvgmjZqgI
643NdsORHAFR1VWmciSDfyyCzi9pG7hPm+loISCDp4a3JGtnmdQHOH30WsrTCdsQ
xvkSsq0r47NI4N/aiOL0ZFQsAPEOvpnOgeqiMxZCymdOK1JCMXackOCPyi8hl2j6
+utn+XZDMTfk9tyaULzBgRn5cQHIloMV9ESWykrYfhIuHbDX5vl8IYnr8RaCq3f9
bH5hvK26925gE98YAApFPpIvJy0sraY7nGMkVMgDjjNBQJsU1bvn1+EUAmiIyzUy
5hoXtxAaa2WpRfgMJetVu3mSiv9r6pK0vNFVZtSo70T+UuqHsKhJeosdqu6Qt/x9
vMup1CfImo5dolSSHqMEkly3/h/yPjRlpiU1sR6OBblAEIyZMD+7B5V7iFTsUiG6
vo+eODd6UlUVFBFaYVJDn7cz1RGk6cDOUA0vuALYcss1MbEmzNHiPOIZv6fsw9wt
9GJ/6o6QO0f4Q6VODLGwQknh//of5jOoepFnqZVH6uRN0rU/fh7ntgpy5mOcYH14
IbwtLeI9wRf+TRi/6y81cw3VN6uTKXDz2Gaux1FnBRzx2KGciiKBVGdM4SZYVq5o
SsgeBrnpWS1h860QuXmaCzIvZA0g1qs4TNH1AXRc6V7uxPRtvx6yar3BIC5AsSst
S4r2DPj1RSN3PKJASqQWVZ8xspG6h8X3V6FX8+PxWu6Z/FdFvmJNkUPSDFKuV0Y3
Ry/3L4xA+rZm4N2G7xDVi9GE1lj1jy/a7Jeg7iPe9xckeHiw9HBuMyZny8MpED69
SWT/HtkftmEyxjn1ky6kVxBixTKJsD3nWNAAJgeHtluYbFXFZbRvdJ4OJ0/aWRNM
HoEKrSaNHdZAbFaaazKxdBoRLj4XVPEzz5UDubwz8xSJg1btMnf9aRpPe05SEgQz
/Cy0A8JHo81XCVN7xMKgqkSF1I3p/S2jxjTzuRHbUtZkf3ncQPx0ZrZSA/xE+fC/
LeEQ2YMq6V+HQncFP/SxdcsXYM+aOTtIf/aUupACHNij7WfMF5y6IlzN6M5jpLnE
25TobSESwCMf+u7HVb8ODrJ3wtVeuMlote4k2pFom6pEfZ1Goc6tyStvJHoPqMhw
3FwnEpCn+YcQ3lQ8FBxJzS629JeaMfm9ILQYt2x5us+RPn42IpznvpAazvjY27t9
yH9CEaI2YrS8H3zmCX7vXQV3yn1QhSSXOz/OkqlyOImdZMyf3CEfzPkZ17ya/sZr
R/S4r8GEBzSLe1hMze5iTKTkGuzFOddnxC1ysCrOiD7K4qc2DQYFruOAa0dTMiHq
z5dfbP7uGxaFAFUNJmXiU/JDrdGcfxjl/4+vtJYmPYqsidvBvHQaDrUJ96LcELpb
HsjPJheMpCWBAarjRnmE0gYBhSlGU6vowrRhEJSEQmj6bsk2iKIl+cJecDATgBjg
/WOyjf/QidqMBZcrH94deJzWoLiPg0FcW1nVVH/Fj7MQSAucY9w6XLu7PlOrMK2x
N4YTY6PuQ1Hr7a6VY+EJuh3FZDWSqoIFRh2TqjasoNOxSWw57veQqwa7odA9l8Sk
F0uZK+SfYs4xZHD+kbX91NbjCmbc/H2sabw+fnrsogB0ppu/Nyy8DVGah/DmpWDj
1emRBJLjK29F8taAOxpCz0ldoOXNN6Gk42JtG6bm9znzeQS0OALk4kcdW/XymA4u
6swcG/+l0uTn8m4hDNrIPuWRS8wwZbnmXYtdgCKsxxbTpPHT+pl3+AIrSkDrhfbh
dAisMA3Etjvv/R9MbZmzfjs3k7vLsWrsBLb0QWJazHsO6ifbP0NAWPTfRvsTSo5l
FUZZB65yDyEXQGcurCglHoEA49A3h0wnm7xIZPpTNZPyy/Hnq1nSE7F1TgtWxdDg
W3BoJI68c7CoBGEyNYN3ktnyYmT5jkrX5c/+4Bnb2lfLOL7z9wZNWBANv32W+0ax
da1VqcKxDVU6lJvo0nUDaeZFI8A/Ws3YlELvvrt/5jyk164LCGaG/HGHUHmQG9QA
5+aqa2Dg05/I4gNmZsUA49nkwTJ0artiFodBTDIYLEcNhrZxsgMgDy7oKcuss5un
D8dE09UVvqWWlNz6NzzlqiBzCxBNkieohq5UNKeHkDU17c3TWT3DYC+nJLHmAZuq
+zuqfSzKIApq1ctPWM2UijGKUZxS46xtUsE0eF16yYwUMcE8S/47qSiuD9j0fuBV
JPPBCQQ5MW9zyYt4QQ+uITHFEhgjq2Bp/oK7w1mJ58qOneAErOGW8nPr6w9D06Zm
2eujTemcf7voAn6ADzCcslGWcm34qaqm/XfH5j3NcU94HuPBmnUzfFumRSLVcTbx
K9h/vSpQ6EXoY5CtJZpsUj/5KOrxF/mFP4nb++Qh2cDMEXnp9jqCaWfvgfee4q55
0/vh7eeMPigoYIfj2zUDtvRA/83qcYoLY0lxySkhpSyhCwWdzfqw9R1b12jSoUNr
LxpFIwCo51jc4egQguMbtcBDDSmEhJhAuqUcSZ55O8eoywtlxaUztdqMczZCE08U
TCLZ9ObLjU9zocdkSRsKUP9D9JD1WGmPewz9Riu+OT+/vWey1idwTOfUdOERwrPZ
x2Sl0DuvJV72AB4/IbJJMJPVb3fNLVrdQ6ilyzVlnd/GfDNrSReH/l7hYhUOnYh4
bA20BjjzDifia46Tnvl0nYVEGfqJf0EKSRnuGHwZW00pC4PsWAoLDrbb4YLd2E3L
6efrsGrVDj349VQMyzOoqkQyzgsIe3hfnNLGC0qYKDmWZ1HJAHgSD/XlVtMjF1Xk
a675/XhSOJ9pcyxK4DZswWSZbPH7QiDipT2XH+0XstCMaKjY8fGbnI7Qs8XRltCN
hTMkLx07rmKlM9ohxIlg/2R23EoB8dtzQpyrb7yU4mqXU0iOF5JXifWhV5TU8UUb
wnNyfRFnb56zwjDlCUw7UR2JHsn3M3PcQiq+1/JvziVUqmHPZ3BDSIU+MtyBX9Ja
RB5h4wNZyDBLmSEOg0/MIHtXA4M6Sq3M4L+eEr+S38KNpsbrlgOk+lXgHeH925fH
Rolv1NnKV0vhJeTHV9XOY+9grWYQCICSvjKNtQEHkBCikA/CkRWJUr4/2Ed4ydms
0vi+ER95VPuKRyVSZ1MkHYOfqoNHDyUvdLYHj/zsCur931nfYCc/vliOD0Bz1qNb
5DBjEAIuCXNlJdJgU15AKYsg6d9C/OUl0B8vZPZmiFE0+iLVzZ/dOr9HT7qJc2dJ
HUhCe0kIW2tfjpaunhimPFlpJdZAYWOdb05sK0xvENh4DWYw/LEBqdEYEU3xpCWW
L/HTlZl1SeQdJ0BvSRvWiFKz6+kjBLY3w8h3KtG3HrZBjKSV3uQbkxT6LvGZlC+b
qukhZnd5BsZ0jpvGc32HDz8p1E7B5UBQiJklwCZFXhPsEhovtAkOX4XlErVOqxux
GbQzK8k+CW+O+0OGhGigQQOefLKdJ3jysvWt7GjtDiLsjfXodUWhps6vsabRIXpY
QOZI3OwsQ49yehtossr8bQCK9dyQbO+asj5Ygu0bMtyCNJbfr4YR1L9sBTMX8XdP
L0yMxa3xCMxDSuIzJf8X1qJydkPkBIhPgrQEq0L/GUsatdRESy5/tXeCBRwPg3gQ
OquYKsW9QW++BGQA6tQcZI6PcxUUbzF3peGjRDc/vCdHKz+bIEAO2wv/b25VOkbC
dicRl9SPOs2vYT5LvUbqttPlF5bIMLVoLxUmmBo4vhpYZ5zpwUrSt4zWzB8P+taW
TMfKEWclyh3h61m6lpnpM1miCwP8oRHyVfa2dPMsCbiQPacIgIuB7tW4tvuyhska
8FL23aJF7nJCiI5H6kHOYiLEcO7QVXxTH+u6jxu3fGXhDwedN7k0C5Wqd+ce/EXu
FdjuypluJojzhep8Foq6pSxpMrRszn3DWVs8AJVCLV9LB4xo8W9V8dFd8QiSZUrX
Rm6RyG481RpAGLL2HDO07oH+zxPGlnyx1IpaX1Uw5BZnrx4JZv2Uelpg/mQ69b2N
h6P2fTQrGWOwrYVYnwwV64ZwN0lkji3MBvTnlX6N59/+MHnpHMMHYmP7cPyVmQyn
uZVHOc0s34ZP0LMPyfq+MG1kw3eWgUXBLQ7eJNPfxNsMiGmYuaGzdPutumAYcqnq
3LgL/TcJnMxUvyLypfgbO5MshrkeLYJeKqYZ461/CPAvaqDEsVjvA6JTg1GNDYVf
KFhPDU+dSZuYzLtuLtKN+/bzNbf4BiSwUb1gkrlF4oQghaYCrlyuQIAEqxry1vbi
1dRqvuHFL6aXw5rfurGd45JngQtMjeZ/ltMaGqPv/5sonWsbTCxxnDkyJ1V8nYf0
RcFpjhZbOMpTzT873yygZ2Kpo1kZopG41T3uZ+tOGbiVGC4LgNF9Y508U9OplZrA
sPLfuov6k5Y4ULf7WmzqebBDO4u8aHe+GyiL7M163CFRq5hVMe1huUA3oTaETGwF
9ExO0t51Wfqz8EsvEt5JbZ+OnpaEujowGpRz8uiAUef/ub8LV1g5wBROyLIa0gNa
U071dpS4DTMvTNfpJDY2G5fD6lWNVIa4QBbMN8oXK9pYIvuGdTCERvNep3GNLDWg
U8uJhKi0jhuq6mG5JpjgCb/MDPOF3NoNKXD3yAKd+mg3pHrY93TY1tz4RZ+ThnZ8
Dv306HxfoOI2Myc57XTO4a7bb/GsifwjhZaDpsySLV38SR6XBDwWBJvSPAfB9rGm
LUY4UfY07oYJ6evkXUsyysIMKtSxPlgTCvluYYPaZAcfkKM4ndeJR2z02Mnk94sw
TvOk4ghQQBh4vnxzfdgSA3BMd1MQjSW3xlkgcdX/Ur82gp+F8DnL9wFpf4C8KXde
KtTkwMfJV9UKI6zjvJl0DbF80792Rtyjal7Hkv+F20UfZNVzqiWnq+9a4nh5bWe6
9JfVx+oGyMUnBKYJCqYfJyl/QrQvHsdQRfUmkFpv3bqWjAiCOJSue3lplUfrvnIt
Z4EEMX6ZSdgS2xrBHqS8WcThrImyDgiB+u/UriaubtrK4Hbz9FLbUhxlL+HaslPn
21t/hgn5p6C+b+9PRe78ilLCOAyssjDfizVgR/pb5w4Gz6A6nWRMwr0TcY/izl82
xDYsz5boFDdudi3tRY3nImNJz8aQrX4Qu6+QuapSMFnib+0IGWWL+/DI1SIKOrq2
rMwS/aKW8kGyNrYEUfhuLkZ9fRSLM/ONNDNb5SXDA6h0PRA2aC3sNidd4Vi5N+q7
cP5VJU3Hu7E55L7zNOheDr8tZDbOz7K7sGsokrrKTvbYJB/E4u/VmAkMgAEettZZ
TYR1xXgdXNKXee4mgQs4HBqSMhvZCpvT6jc3H6++bSFCsnUmrSn5m/kozycZYABd
5b0Y7IGO6p1Dc+ZBpqF/pl91OCH1n8n7lXZAiWtmtaf5YNsU9lutpNv0lLDVSfm8
zvfVj3gc1zA+JvdE+bxj/lelht7yMIA0JwkjayEcXuS9E3hPtF+mvPtkDdr3m8gA
6u0Sox4ceuAzEi80DDINbuPf6mMJFjuJZ0sBGKqPspRBYFwcRb7xJg4e4gl2ClFs
pCsg4LvsiwRuyPgZubt08Y/LLge9N/bv8ZhHEJNPlSk4qwzkBN+7VlhY1vx8uZ4e
KIWVh6dXUmGZeLLn3LBi4o7n0x3639Vv6mViC/en386noMG8zK0NQ6rVNYFssVse
7FC2f8P+mrKYRfBB5KpJ/pLvty5nFRjtkG3qDa3GFiCkyQQ9meUY/2Bfsnx6H//f
22Et1oDKUppGmGdISTiyxvaT12cYsSOc7U/FmEi9A82ABvIs80o2/LNjx1xOQ+v1
jahWaKCOBhKWpPN/T6LOAcNYYjf3SybkE27S5Mz+VmKKEomEA2qa/U/ckYWXuB/i
hZJ2awqZVAkZGmM0hXo7XRc3wT/KYhIGeagSZ8gAB9a39V5PDJO2PaToYiDmN5R4
0dayR0EEsVr8mKEV/qlDNmT/xUnD2rV+KtHfUNJKGueFvcKf6AaB5P335gsj7TdU
vgZ2H58dkOz2BNXctFA56oPC6JAMo6EPlrs1Sv5onNIyY/Rsnv8z8k3QPDKwNyce
hV7ajJOnwHfolQEOOMWonyEr04E0jAzkKlMRlY7s1ObDJqhFAgDPhZ2GBUN3Gluc
s4agHOsBM9LyC+XkC3RTTQ0CGQMqUX4s5XDJLIwuZU8tdWXpyY6nncKhnooiBf21
/hspejf1GgulvGbaMZJEwn0+pZPaUdVmZSnuVjaO+QkWYGxjUoPNv3eLRhuDWEgj
RMumecmvo2a08gDgr74JG0zFs9UajtzI+WeNSq6IWNPdJIcTcbFJ2I6f/gpdtOns
omg7taETXJnl+dn50uj9L4B/pxs0d8yyU3XZTbXv3pcSRz4PoQyiW4QIYCKjaYkB
tFVLoyjyUOyj2EgBnSeOwca9cSddnfGemdoumrCYyXTALdtKcCMCgmMZ5aAJi/Gw
UHrV74S45BAfyJtrOopqodIQy+r+7hiSZtabfH4CjGBTIO4EMSoW2d72y3P3jvbE
5bq0qHRwdrMW6eJwPxwGPPYE33A/thniApxNP0dpgn/XVqxjWaY9tXSorcQLipZ+
ekIbWKuIN6db4eqKxWqcFouMPwYytM0cNZNUJqY/Y/rMzn6nd4t4Bw7f7iU2Em3b
vMI9JTf5vf2NwzbWVR1paivw5DNzn9/tZVS4ecIwmuAKtnaghC07Xr4gtLTd3XpI
tjYJNFNqSAEExQgztzpk6QwGdtARpI6aCoE2i1mVdfdZTDNxO6nlnyPI7RLnWjvn
Gjtxb3yoYFzYVvdYdBwDOOFGnNigAY+cVeD39Fs/09HK8MYYOtWawOZc4/zxbYst
/Sme295Gl/YxrZuq1hzKTI+FioOsXDPrnRjihthRUiJaqPcIt0DDR2IQI4dPOVX7
uAnHMk0dTZHOVdzhZfukP+nwloSwjoQgjwTo6zTEvdLmfcBOfeRlkSN3gULFO9I1
BtkCR+yncfbnNlX5FEUIPabW40MGUeUzyrS4ibrZw+9hS6HYia0k26O/WC1TcQ7S
9K7P4eHjf7K0G6MdHTJ1yjNWCgZWTjOmQJ0a1vphOkZYUThL97ki4M24yF7Jc7xj
AFuZKNSk7ByBv4D1goa4LpOPXk8OInaQk2frrW+OnWcctfOOFWRKRjWsV72YxfP1
tNsq8lbHFY6IVK3n+r2iITxs1eI8g5ATKnyyUSQGOMKE8GyZO2IrOF/RDZ5CoE+M
pWY2TvFTBqrCaN/7ZDGeZAn/wzYWRDYVZWVKuHZWCozywIvbVe4FP1PHl9KztsB8
Fu86CI8Lr5PqnspGb6NF9vu1xLEN8WQxx+b4xUwVyb6amvORuPH+bPgXhXNM/BoT
OQXARoElXiKiR0psDoavnQws0vGhmAegwf4a92TwIQQvr0CpWYkRkcYReSzmDThs
XmJbqPUwDEbu5G9wWkAnamM1fkCAD/h6ARsYJspsLqDNYLT1HooqpcnGYUHZwVZO
UnKY4H6UW4joWv1g8rHdLf/ogouEmij4GfwQMKwVVUlcw2EUuDQY6Wap1RK1o0/p
WsMLW3SOO4SgPRdAEbx7AvjnPHdj8VWadLLU3kim5GUKZyg83JTrSLBYdFX8iJkm
JYWFZF61AoaPkGvOXnIxDp6OQHhSHISO4FsgUAZ+7yIsH2DWMigUxpWF+G83ajwj
U927GE8g/WcPJlxw7jE4wMb1xdQi3h9sAq7aFoHLT7xv3LBouLl31rJYpNZWtdj6
ZtXQtdl5VjhMBUr5Xf3Mia/9DPMtd0/5ONlw8UtUWCYwIeHLTm1HDXXAcIe9niB1
Fxi4s4b9JAl/5mm/qgT1N3C0mZ9hQmC9KJfnJqneMm7/45THoTCG8jR864z7xxtz
n00zOgiKtemziIlG61bPCZ33VVa25daYTkQtUcUpA6LpaX8boY89TtvQ1U6dAcst
NETK3gOljxyDPr1K9B4tbIC7d9aNuwI3ivJrFpFI3BUpm8mGGECt4MtYF7fBt8ub
A4FGKLGQm5BcjtWG43/XF12rbGov/qshplsn8RgaEGY/DjSCVb6x5RRERptqMceS
vqok8MHxPlvWkh84xz8cuAz4W3yG+oy3z6FZTBqWGlx57ojeynqsfeTmC/HZ+8Fo
rJBaJ5l/9gWYfJbUTtcJkdrxxn3jgPvJl/dgdyL6Ipkt4E91RTzFbYh8sbQyXRd1
lCNkWE4lZbVij9fIvAqT/MlmI5E0y+eqYqqilfAzTQlp7l6XCepEceqS93Xy9ERc
itx3s0OM+0Mn5N3tdTaZdqKPEDZcaddDFg82JIfzf708ObqfzPhTWH5WKPcA6z0W
Pl/Z6KRyIDmxfg6hFXzdw50tNdDSMOAhwBPfV97zTfX8nZNHC1n8qcOFTU3TNg7p
4vvlYngdHddyIRmzO15lAtMelf3dDqRrinKLwvXHjiEAs+5yjmhXKCtVwid+Px3w
8P61WPR5VQLqzlR6a7X45eL+daF3Lphip7xp8VTm5SUQ0pUk169/hShzdklvaHbC
EKDZSGUiU65Bd0XeV6Rdc7UzdeZWp5C+dyKlA23lVUhNY1y8gZ+NRQy2Wz5WeY/9
U5vIdnBJqr2ZKmQ2vtkw/t1GeZctpcd6Cst0Ed/VtsRJhIhBCYmfhqab5KJpNmsL
5Qd6VuH7ARSfU3NDUu0KCtpdykimQcShtYk7ZoF90TDV6mEne8P4Qrqp/zIXp02e
QI8gOu3lOhUrgnLu/w2hCvnTd1hb4DtPayNDBcTjt1yC4rUJxySp+arthgOHUYrc
Z11zqBfJV51KlVMpH73O+k3f0EDLXaxWap6hnu4hXXWzP8rQkQGblSKxQlx26PtJ
IjiBLRSsnVf6hB1ZVGZAHAlDit8jLuBJowYst5zRCmnyzdWTWOzQhNxvGPtUJ3Nz
CJF+eYD/fPDaqE8U28hKTBtF8El8U4txKCyGR/PpkdNyH1nCW8WF2XRwB6F9lZvQ
sftc1fm9+5lmngTJAvtLfJ3K9sP1EJSfBkSpCGUj7NQN6GkitlwsSAxzzxofwXTD
sJGlMdPpeSc37an/rB7MaUmjHLy0LRV21W+tihMyofIFJRxLhWa+2w4vyK6WVSZL
I9I2pDMVpTpV23LCxWtTf9kU8wz7ijwKgjdfRIjzFBSKU1cCy74ncx0E9UZw+YWw
gXEF2Myu31rEgtipTU6+s2orm0vgDuas6zFwoW22Zkw7BdKf1xVf7cpGLCCGv/Kx
0ShzoQJ4Rpvf+vXivxTHPosrXkA/ROHF7n5uwJ7WG8tn8LiynsoQTH/wGH/Wwo7y
LDrFtzlwLXqxgD8WXRkgD9rfFTl20b7hBSS0cVPqMpgKNO5i4D1n+aRA6QoyMlOv
qGC9aOMOiKQDi5i9MzwerVbNpAPz7zzghOLhMePi9KTwlvC6mc1MJYHpRd0dx45e
CQ1vGyrm511O7Ka3oG6whznD14/2XkA5gVvW2yUbc4et433+HeV720BZpD4lU9Jb
zfjNntG0SYgQOYKwCI///6kzZsjhJvM05YUJTXk3KVRHRSW4c8nMyx/wcXVh24JK
ptp7YrtKTH5yaVH4yUdHW2CF4X0nNQJ4q+iLCvHT32VoWsGoRl2x3YRxbQiz3PXh
eQI+VBF/X1R+a4l/qsiU1xc98u9L+d0XHoc4xQkkVW1Q/EG9QbYc5mH01cVgWCXw
j/yIzEwqZKOAoESyXnlOtXZ/LkIofW3c8+FyJ9HzUyT7seUR2xc4cAaXHouWLQBK
Xb6IqJnlVVcKUfhQ2ytUM7LUPDVOdoT/qVlHztKV3XwDA/pmwTRP2nmnFLIjWXj5
HSb2GYX0MbLtOAx2+ok/N6PgthSel2yltdIn2/UuiCcMJ/GTd+FyTeTVWZInhpmt
uBtKgVC7hRV+zqCSzlJ8Ou1+sRkgKM6ZUsbh6qRYNnGtxMRHsxuvk69mvDsIU8Uh
KEouh1NHwXeo48H/L46bF+AZIhYdBjEFNSZ/fD12aonz3VXNh3nzOSP8VGlgR2kw
HK3eEmfV+Lrbbna9kY7k9BLVmT1OXfo4hGbuXCZEU+6AhfbCuFSzyWpj6m2PazlP
YXr/22XvP9V2XGb5ljOIDIHG6fXniDogT1h2BoIBqoP0LqBgC4Ejs17ZvkJoiDam
jpJ+jpyWq/Mr/hNG3tBVlptKBJ9rf5WKAT5gW4mAXwDhF0YqGIhC/qQxA7nucsuy
AeodOgbls0tutL++s9BGg1LAE6WQzhk4PKiGDGjk8c3xb5P/2B6EmBC9YZIkYJ1/
HxAckXjP8wRD23b7h93Pl7DvvZ/7Q/V7+MsQkzHKHZr+dyBgLbojcHULY6wSI1gN
/tGDSStcZDJaL7sUq+Xq/HVDR82yVMOVcti0PnIjU0Z5XNgRFjH7/yCv3HcQ58Ln
3hR4HcAFULyGgBLGdT2l91ndu0zns2EJP2OC/VtDiLiWwtghFVRov5sPwSEoBdyy
Lb67UJ7pVFL+k4381IM8wbGPUG8q02PLxsxg5R+HzGy63D/DQnfAS4eVpanejI1u
elo3yCpHxDRXpqx68ivE9Uj55hc6inW2ZUOurDb8Iwgpr02oPkre9jM7jr+rvQ+y
IUIshKSS6xjkUBB8yBTnt5cqxHRYfcD6YiojssgCQRussBMbo1D4pmBejx2tqJ1h
yPnog9KTVG7Rqycl/nHdZcfnCFjX+JE90fmKKphdoAuA3fE8mK3KozP+YEOG3xxl
ReOafg/f0xdgBcTFaIAptgzsgmcODzrwxjYVcIJ98+qEcXfvzbUIYN5o9/rbJ43W
wIjfe1KWpKpyQWJoJzN3FQ36pVqtT1cLgnXqYlmHDBQsn4aq3naBo/FAo+Cnxebm
1zNbJUxRB1SZbJ035Ddma9gA5ipzcKHtrtoppAR2T61409+8GHfkKQ2Cl0VQE8eN
iJyIIvOxU6JKusvb4OYSvln/WTtAxCDBWniUnHo0cX1OyYrsD/jVyJDzPmw5fwAl
xWEd0EUxiSxePiMK0vF/O5Kp6EHxB/wN0izGI/xlhcz9TQObxUtwTNbMapjPJS45
vT44xgymHGVb2qDxnG1ZtlShQ9qoZtKUd9sXZHncV5xM2nBNZwp8gNlBlqoaYb1G
arY+iazE0AxPE9JhEDdFUbWknaEk3Y3X/TiaP50Kqfr4K0k7EqZmPPguZdRHTSyx
jMUErmS0Cqd6KRD3dlbmM1Tl6HWdpIqbtOHubpOfA8GrMSbFuIv2oWYN3PC4oFwA
CTWV5m/JDBMPETwWjK3SDCvFs2RbxhV5m2/JiOp69cK69H/lDSmOb1OVY9rdjTpo
GTqeHKkNZVl0tiAoEN2CDclBrHfPXJye3KI2ohAQ6g5beshhtMiU+uVVUNJ7M9mg
1fOUmcTk679S9w+4EZENm0oPXs6Y0W2B8/Ocyt7KNfe4dFRJeebu7IkLbVbevrqD
hbhtapyrIx3Gt2JY7d0m6jRK3WEYQSW58FCXgNdbLSSikM+0sQLodoM/Dqed5jDX
Z6Bc1W5axVZjZsM2PhQhYij7KfEtiEKMeiirxR54ti54CYkFWrmmw7C5NHmB9OaI
eZbJnOdtvgnUaEMjmr2uIAbTKPBjuUGeGlB/RpjR7JXM3OrPZs2Kk5GGIazcHeVf
deg4fnahDlIOyOIXic3KDWLaJG7JbQbZSTGKwxLQzhOSQouvBWO37hnFALxHeMAC
F4BCfyrVBHeQ0x1MOzzIFJZ5v3HXQztoYENv+xgFaRNzyYp3uA8u99n+KOzXe20Q
ExZe+oH7zrZYzGeMEpjMS1K9gOS9rkMYTOw5MJu+qGsgDM/KFxSJlExygmVSUGQU
3neKfgbBbE8oNmwTihfHUm2r9gWcX95OU+R7QS/eoLrQ7ZQjaHLgkoIV4sXyTED3
p7ORhrJH7EBlqts/43VzEu2ndiZqIEHsPA/1oX3bhJzy7ZWSDGOt/MvgtppHOLVB
q977eGxaku4saxr60o/IDrqzwauvaPGR8UX1TkL/E3I5JWLZgOjWmU3i4kOVhQci
SEmMl7BbPef8TSKnp7FWRZ572KAvqC4Sdws1JzqtC1V/4yPkfDaFIW/HkrV9x8uX
VE11UFWsJ+uRor/s7mCfLx9pw05siVBNM/HKiOM5rK+V6AgjTaJL2mgYpKAt1p+e
2W8FGIDSVByqQyrZr7Plvw1pvsuPojfQ4V9OYzvCc6Z7WIj7PC2uRlDHqYF3rEPy
60dF+EqGDaKaXGLwiNWAQJ/8Wc4KJ31/roXKS3DPp5Hznf7k+3k3eYXlnW38eOWE
QqjD5sprUffiZToz7m8DDjeQXJJs/adsVoTb89bGpjCwdihhzH0Rby0CFxdkT+vT
iw1S0IIs0T2+HcdPcHL3ExMFOO3ZCFY+URo+xRHLrREOenWZRDy04OU5jjDp88n4
TAEzysp0OzQBeTQvl+slQz7yIBfC9IDvl3efqfpNjRV9ZX0/mNoGEBJjWc6IeKO3
8WH8g8IpYZjfq+s29lr79xhp3G892YhkJ0Slkr1NOpDXQq6GdXGLsYOgoRLu50q3
i38OzZy2VDLb49Ykv4Wjsm8LRj9zpe9FiEHr/bvEKI4PS9mXSqpkcN9EPqMY2i4U
VjaRH7yODHcXfd47TccY+v+Ns5tSh3VXlFGRnOCGEfbgop0zOYYVCJDV2qf0qZ/0
B4ClYXKzx6+MLFXCbLBCydlyqQQRRGKtEWC7WkmUnt8RM9jdk9GjY0vcu3fXM4L6
yeFf6wJES2ZfCiaDdFtjM0U8OikTCypuq21B2O6kSEd3f26hK/xt4pmMb9NCww1X
2fTalD8CQSyjrSDo81YqnE1iy5qDLAriMUOEH90J6ypkdu6AgMsmQydT5Ub5nEWu
eb4CrRcCGEkYFvFl9ZfuYHiAiiV4HnGHDD/c+lX8RYvfxDFZqaP8Rd7Li5rsciBY
CqZyoO3hlZTbZR9/PR2MB8uWsrRHRZMO2If+lcO3WY9e9A/q5eofhabaTxjXP1B2
/ih7EvXhGZMPXtEIuZCVCC2FLhDQh84Pv4xR1F20q+K3DcGIOA7z10t/hDKa2fL0
hmzSuJsS3hU44AMP0DQyAQn4lKD8Rbz5GT/X4dYPxpdVytoh4Aj7mnza4qpIVwCJ
I1kw9PQX6qPHC++F4eeCc7qsG9COQVgYaiM/u6+mlaRtj9J0buDe8E8k+hRVDYa+
52zK7X/kAaQV5J3d3LPUVmgBlZ7/psD9wXyTikookTVg7Z+VIXRKIywr8dJUK0Yy
lac3NQyhN02zM/Pe3G2gJ2ZLuuV5nnNs50X0QJgV4YocdEgS4bYZAupKQqkbGzME
sfzjtZjcjuSTKIDuEaayriS1JAuP4cMyIJBf7bdfuLUJNLTuGcJA+bBVJp66+SvV
dgAdlPlPq1NvwRaUP+8WB8LRd9+IhG3lRsZddhrYtA0ZlWIIQJqWjTWNjBAoMYIn
gXm2bOPuNUITYXRgyCoskPGm6t6cjGgZqYh3V7xI28W7X7xkPnsMIp98MExSVYa2
WA3ctjnnY3MDqE+o9c9/w/aW7z3V8DhRljDIXyhTKzWCK4o9It+MjbM3c35cheRL
uDikXHesUv0HX8ON9vYb6r5G8r1TcqhnBkz1LaYX9nLrVCa9JKiYts4t0p+rvkZ/
HsTnooKvv6KGByOtkyw5oJYItyGzQJmdPVw+Wc3iHqPUW5VqZuEZkZElBELVd1Tx
Wrj0nPx0IAd7yUj929yS+ZV/ZqyBWmYPDmE0oXCEtFHyk+lUgpuLOdt3+Oamp11P
b3tKPY5R+gK+iYI2ONPQey7d7AKWpJ6Px7Kli9E7hjPdUCOmxAukAc7lcLtrIffe
V//R+zkg5Ma+SnuKuoM7A0UR0lVAtmVfAzAH5jC0j7W4A1liHG0emsF8OX5EGr9p
Vs7msh6eR7CO7Okl0eFD+7Nzo8QQ6gu3e16ZVyWQb8hnktQjmuOgXRSdd5aJzGB8
s6fhUoqz3132kHaeX4qzvz+qvKzwvuUkepH36x1h2zb0HEHTVcqkXqBTvipLN6SE
mBEAkajDzCtSeGmEw2jn3iE0dr5NHgYcV0m8wRfOKxFuGTqHaL5WDcN5duvK47lm
uflBhBlvMdzd+AdazD9YJYlMsSzVU17b5N9R0ldUsD1IRzECLouTJUKVmtxYlFxa
4bNTyhr7gO4+RTbQPDHk7IL6F3yHuR9uSCdSdo80FlGpkP4r1UqYTDOhF0vUQ8qP
mnRmONIyz4+sC8v5eKKRRAHb2i7yDBGx6jvKVJi7fxEsF8pyXE3Un1v4xARsZFKD
sHY0c7H7YDE58WNE7WWOQHhm72nMSPaWBk4ha7ES0sFCoEf2xg3efBPV3KngPyGD
RnE1AOEMrFyt4bJsd1v8f/XdCKTkasF91eoedNfTBYxnQvsJTKAnV16ZKZZ6gz/u
A2QjRfmX1NQi+FBo4vFyDpdJqV+nsjFMS7ZxcwoSbmZ1v2uK+SjP6S7dAOxu7C+/
cqDVyb/fi1mHa9wZtLoWlKQzxfITBBxCU6/JNuA/wRsQKBW9L4KkdabSV1dXNztn
fLUa4e38USaEcEdfYmu9wKqFImOnnH29UoF3FNBPgtTDaH3hOCcdZhoI6RuNV/cy
UyZ3POGFx0yivX0cCDuVTsnlg5rJIrJi0ijVfwuRofJ+suX3wTJPfvqqgQgvOYrw
J5lzqa46UG3sp2kB2zUpQQhl3TLogHhGpK7Qnh7s3FBAzWr1hsSprNENEkYpmxLU
OwJVO4Gf34LpK80Y14nqUXSuAz4R6dMWiTM4iTTCGzcJ8WBO2iYHqebDNeEHiBs+
YCfpPzL9kRKLFotkaARB7P5uQaUdhPOZMtXjSRtPLpl2J08RI3bQryafpvhZSz5z
S0rhy5pUZxD7/bd+vSFz/RO18vQpmrGOBIvkK5zbP3gYc7850+DW11uQfk43n96s
LOIYdlp+gmLRKmPTuxonvvWKNNd9oFQHloXdi2yevao1t5ZUtzUKS/BopM3s3X3A
B1W7DFko3DU8SDMFEOTrJnMvWltimRuXr3QBBJ9w5paA5+6OEJCE+A26QHiDa8oS
ZLCX2qVUV3qUczXmiMV7zdTjPAWcdd3WTjTS0/tgyax/QTh+pmQ4Vo5ABoTzV7y1
8Wd4q1rwo0VzzkUZwG9k3L+jRGBDxZCeetjpn6ch78mrQclQbFf7xRMvPJjfExgt
pGX769lR93Dktq4KQOL5ZZGHkjnEtUVbQ05MDz6hUcc7NAUGEJ/WTQ7YwqeDuxPd
vbzpxCeRjSrCz9XTMxBdvDeqPF5JdUh5zTKRUUfqlts7I1bfGnE6EYhzSc8lDess
0LRIsGn2eUxK+dDLHc1qd41bWZ3b1n5SmGy7Hv8CR8dlx22QJ8vK8IaPVJvUmcUg
G70GD7b7fF9eV2pkycy4UHfblVMTkiWDbVzoRqXIkVrSmWV7RQR3uiC+/1YZRAUS
lr1Wz+DnfbKuw/+Xwd7Wy2oEQX02Gy2r89GA4nznQlBXh9OAiB1RUNEfRcV+WD1d
JA3uFoQ2HfdNUbMDapyEvNUk9R773PyVnFIOYIo7ldW/IswUv4A9UHwusPB8TtuI
jI9if94NPQxZ3uyddeIg+ifmdodsoW4Lagrl08J7rD9kLy4LjqAAv4788CrJukCg
zOvN2B1uYNt5+pw8OLDW4VVsrOrSy2AaIHdyC6t56Cz19GQh1Aw7N+YnVRhIhnEI
0aoBhzvV9aAuYhOPMWH8azZWGwBzcnpML3XPZGGcgT9lL1Q71Fb8X49eP8jioIb4
yJQXo7MujvCaMey0YapR9SalU+OISkohhi/Ts/rhWcA4z38q5gqjjiUVtqoZOhMo
69LpRnPQzYYHCh6dBzd3WlRFcR7nicyjUksRE2RQfYhcF1qlOa3sqS5VpYo+5zxH
Qaet2z3J/paVW7sL6cRXncFKnwG8ZmETp60uJ9PckoQ6yIFmmZiGJqt/M6hIN3zm
g5cJljg4chzHFLRF9XlSnXE7mrnbdzb5rOQJtEkzx0iKcwkZIJ1/xjpUZ//uxjsO
xiGfv/rNGeoiyXzGElNV9WVSxYVB62KIDoBIkPbBaC1YOcQDJ9L78jDRcwVsuuTc
NrUDlVDxABeBcX8fG3w891M4ti90XW8n4TSm7Wd6vMg0HB4UYxW0xFRbsMdr/ELK
23pddhL446bFOpEv35vi70G+a0gM6Kw3RDkftJXaAzF8fivJAUb5PzrcRf5hdmFc
94yzsc3HolMiUx+qv/N2cxV0lnWsbbYuT5rUXHk9xb8nQ2qcGa93QMDurxd91vIU
s+pyIVkUpW/On59Mr+xTJ6XNbCgvkb/oXu6g9ouyOC1TG1iiqFXc7E2VljA+D4OW
/ZqHCXX8p8OK6PDCaIajGPSEaoDp37dSSQcC3z3NrwSIxegCnoaEsqdT/b1A8Uqw
sSABUXJ/wUcX6WAN2jZB4+aNmRxT+cRNBaDFBTJ1Jk7wux8qDABhQnznirNoeT0j
XIXKLbUFTF1spP0pU9THH2kZakL3JQWy/JmJ9GSER5ubZzZ30M8ioD6yHOpHByLI
odjpJshH4FwxWT6qZba5ndeyIIwmlo6/ddeQmjidBTLuYF3zYKnxEoIV4OE7IhSU
ZJORXriYjAMFlIHoNswdofzsQXW4Ec+oLfJecBAibrep0leAYkTtk4HAvnI/9knO
gsw/H5m5sHATrjdOlxzX/Qtn1UCbXotAvOhN2NydliDUM2bVGMqHgXCfqDEByX2T
gsRCmFuBJ7Xiw4oua1LZl+C9CMT/35RSrrTuIf86tVGPSKQCIE+nuF7scQI+Pdbd
4HbffLY8Axb4pLt4WBwp8PWdMLCzKYn3a46WjRjnNRKXFR8UqMwTKUNcc5KkWwe5
XAN1d9bHhfYH0+e1sN3ENt7PZFZ/ZqWuIgo8h6v3uFZzWJ3Wi2I20XGsyiwOA2PR
36NS+gPVg/USlOkVjLX5Pu61nh14PNo/IyabuPnnKBGcvN6K73z+17TZ5Ur0/LCO
gNI9PFS58gLbmBlMtdzqjOAJM9NgoVaTi4aXeMRv/Hxgm/YdVt9RP8ni1mUJQQSf
uX72bAL9zJAdQiV//y7u4kp246PBjNSRR+QI5R2qWx8FroBprHV1Jn+RX+wm0XH3
v31+gREfBTujim04BEqIe9Moz+R/UeM6A3D6ZPqJqLcXBwFU78RfDl7geU+q9Ikz
CN1T86mHA5F1++azq4q55kb73eDatTErDdLYFww8GOY79zGOIXR5gkskDmRg5EGE
Reg4Qb6fbFwTzONYdCVsP5NbXC1UXXWA2Z0AJ8rg7B3LdhCt9OwxnfadZdV0Mnfa
6AnJM3tab0/fyFXajDoSOUwIw4umS8jUpVtVqbyab3Mt0NO48ekmsDE8McBPPsHl
hgJvrUA+W3SbFxiyFV2XPVZrVxY6b6UY9+5K0GJ1g+qhB2f6OspmMJfhNs7CBFfn
BzXE1wGZqxMajdi2sgV5jMtJr7vv1PGmNugn73dO+SfOXUeGi8rXVO/GM1yys+ER
coZlN9LJ6lMiX8pdpItVfdNDQ3w08Y4UcdVw7V/iL8OyY1h0cdaVGAOhqHg4b4ps
bsPhwK4AXnX+Ta+MUfSMdwbj5rZepWMdCjNHW5ifnnNIJVQbHCaZt4ZDOeRUXUV6
QjFJp/K38EDLi3eYFSCtDS0fTEAkrtkLvBOo7dDNYu1xMDlUYf7xeBLtrbYT+gLG
+qz16139VYDrivzfPbSw7wFYey4BbEYxIiwlgJie2pKngwAzMl0tklX0+aMgcVB2
dts9+5Y0USjGcvbdOmI5cxZZriLZD4QRRr7mnMRVsAg862tHcc1xMAf9yGxkpyHE
buDh3H9Y6lO0ryS1Kz3jK0blpV/aWFY2fLIefVQjf1+/Do+0FkgUZzWQJ/wv7A2D
nNHKlOc/IhhxPDci3J/bhjYLQQC+1EbI42tO8ut37b4UpkpETJjLr8u8L6GS1Tk5
hYkZlwj7Ya8/5YjtdKs5fO0xWPOiwWfjr9dDRAckR2t+m2LiuD5kOXHxowqfvxXx
Nhwy3UdnlGhS0uTU/tj+o7Pa4SPnO9BWDb7O3neDUwLaUr8L61X1tc8l34fEQTgP
3MBqaTFrgisjDKeSkC+ZSvL91z0DTn7o4wkXredUrdam+xT5AYZ+kGxK1mFCu2Ii
jWHZ0l9W7Wz3DLOQ7EwYROjTCPZ5pLZvpS12YT3BNF47Ker8sPpqOooTbDFi0xzs
2UXBB8pJ8gVoi8JDot6VJVzFdbyiARfXVKDDvdd1MloC61hRNd+kVxA5PrC/ck66
CqT9B3jslL7xz1OxSN2MJoLgbprDfY3VSRvia2ppU3S9ZGheMvNO/d+zX38kZNUS
bR8o8jgDKisQ0unD5XuaxS0PL6jZXDHo0+VYyueP/zr9PjFZ5tS9isTLrmGZbM9l
NLlefr/UvL+GQ2+KL3KMkefx3ORWB0Jyw/0K2UU1/wJU3UOMNeshvsm4PkBxifuV
gvF+eo6D8Zrz2DlQ4i47yB7hh7G8BWzwng38u/ORxcXpRh4JL/mQnl6oT6su+VL/
ee6Mm6Vt8M8C6eWU8IfFQWAOc44ElPbPxiuP3D+RUHZmWjfv8qjbexTk1FNlyYKO
CedwsN4E8ytwVP17GvrbN7xaijgH/+MEg5MCa57WsGxo9umGSD4CUMcZ4Eu1gOg1
xkncpsbsGa2abW1k/S3lPEvvQrySsL0uNvk++n7zz0UQ7Jml6WELG0lES1ttvpYK
4bql/VDzcNxX7MN3GPpADmnrryym94PxnRJRsyX6XcJl97UHcIVNf/Bm8rfnB7vI
B/Tm0WjaVdIzvoQE3zswwrp7hez5TfWtxRJRX8nz6pxGW5AEc5ZmpvZ5I+uTeZuw
eS2PJAqN6B5ah3RqaOsGat8RDHFo+v0Xgf/Rlp0O2fMaxiZWqcODUkyADlgIYyQ4
jzCOctehH/1fGjQa5SykRncYU0rKWpnZPumfx3zJU7GegFM0OZkbrSiuktd7Zh1m
gt0edQmhVnrKMapv0TQ3qCnm3NUZ0KxlS0FqTf/xwpFcGmpkKCaFqQgKF9Cl8Bqg
6I+FA/JGjZW1/vbRh2but7EZYD1/cqZCAbqttXSEQDV3FzP0KxV58BlCVxQ1VcgU
c4ogv1Wc7+FrSNARXhmxTunLZFsNb+yaNJ6i2Ys824BP7JROhux8M95pIwHLEMxw
gyP94wiK1YNQWHeBLAYrAG1Pnfdh8gxWvO/xCbV6ZqhVB1dXsjaj7oFpwvcEmSym
woPQHccCideK3cXgk1f9rfLfz4xsZQ6bGxK/JUAzTzcFzBh3owQBBF2f1zCYPxsm
YQLx6XG9IhsMIlrazgQaevMZNYJA7e4wad+xqibhlGkQO0U4sn6k0lIf7W9JXzTD
Dfkwn+RivPo2/ZpCRlfvLDdPFYPHc8jp45msx3LGw/XhugaD8op/FIlcEycj5tSY
X7khHF9VbflgeuMKpROeyT8RCg1YNQdW/gJqHoKoz+HCKDnOFh/EMl3gXwgdCnSX
27rEaxG6OZB5OAUIKdMtDWjloSrHHKtCBpwe/Ce0Zn4PBesHE32SiATHh132eh3s
r+2GlcfTMX0ar0mC+srb7kyA2WWyA9SuKj83FejTgeWjnMgQ5OyDSq2lDgGANMnT
vf2eDeSiLp+0LuMDlFxvtjloKYw5CW/Vq2sgEJcfj5GnLcjr1yaMlIMfZwCp2qK9
4sX1+D11cxoOyoT3qBpexBpkXDWt+p/1GJWd9B08BHmppOHsGG2Gi16SIEKPaCO7
y+5xykNxZVMO0uERQig9OYoS0R5C/it/d1PFKYZ/IzBGcNhZaqBvbKUkV2k0TJ51
T52I/1MAtfdsvdD8S1xeNw8VIo/HcDnx+HY77djOI9nWtzKVoH+t+qnrd1DxtlRr
aQyh/L2lq5Y4qJMttZQvU6pmsTzh+DfSqo6sZCmvUtQM1l2zSGsZPh0RwN/6atnZ
WsrzdCq6HaFuwD1zAmBOP4i9OG8yeWWNrdIoaYLrtxKaZVj4b0eLZYczKioNkhk+
Woh5Kna1q2S07xtZvv0hyRXjsPl0oVMG/gGPzqIcIkAjVF04l3bSHnml87b75UDm
ifIDOfdWLoXqzF/++8YuVOFupS08G8pj70SNTlHulIaXUni5snLUXcntiuBRul3q
8waMPzSY1YKhmyymrk0L2P2iJ9thigCQQZfQ8TPq+lZIoKab7FhYUttd0VI8JogD
4tW4POpKlABfcFyMSbi/mh8BkHDYmjwQyXLe/4MCrZqn83W8hRocyFc2ntKctBJ7
XZOrn8h4S6u97UXcd8DVSztMSxN+rYmTriL0hI8W+gfqF2FB5g11mvss8Tv9lrlP
3kqoGysxutPBshCBeed6VxesueUt74Ca8vrnuC4N/MeyehdBeDcv2Gi+8+hg8hQ9
/QKzvPyqtyUudQcuG1YYddWI3oGTZ+G4KTm3LgOe42ujvs46qilVJpeqfFyt7cxK
3B2JJoQxi5DDq41ubielpT0WFW9wK+vMh6JkLg7xQl0KhpPOcAErBT2QOSXcColn
rFbZQ19GWey9kBlT4+JJ3bT+0HvLbL7aO+zHmorYJVd9OCRK97RegUcnRmQj+SLy
Yh9g/9wHK+9NqiZeOCDWepXcM3Tlh52XU3TK1VBzQK5o6GaBtyEtmB8fU9Qprp81
48qNCpzBxQzwqy5WXpX01Ju0GuvVAf9zwP8wY/Em//fovuPSXbpWrmWuue4tVow2
dFmrr9M3f1HEyHzleDOQd0xb8kvjYQRwI4eACsx28L5z6L1L2OZcBAwxrsuN7U4F
wdDOWlyKmMd4N5L83gWqu6Enlkf9Iq4V6oKitJfUb/IpYgIiyk5KhgEJQdml1lyw
g+6dgJ14NwUzh/EdTaMXUrxgzJ/jw76Iyl1qXi/qeJujWx+vL0W76HGx2tYr0KFK
LmUtFiKTNq5lPN3pt4y7Jqcs0x6bWPvZk8LergE6RB8yTSH4/3/4B00lyZqWqvuc
f9cCO1vTLn/CvAAmZ1/JPzWooVNec5KLA0rt6Oc+yNFm/s7cQZ/z8U3P7JIm2PHi
oDbf2+4+i2sp1eYyhVLM+jtgcq6ZdaBFUygAOvho98KAH4Hzv33Wqlh0K35c63nd
JWAVXJNXYFNcWjh4wb7ue/H6oYC6x8i76m2oET4OaSFF5D72zBF9m8wJWb7ALrtx
06wvqSEsi9m5vOH7qPX9JDUpeIXKJ/eCFJHUNVt8Gue/xioN9uaUezi671I38LmK
lt4iNai2K+C0Y57Wx3jBLBDk8qWmUWcLszG1Ix0L8qY9NL4dNc8Ev0WwAj/jZcjA
TJac/fkpu0UQGFYF81mNoyPaxwBUfnLCmaY2979lJfIJ+KWpe/AFdOTHcBjsXPu2
P0nTU9UYi3XL/hSJbZQzhPi+F2OJQRwGqAoEMFnFg96506UA6x+aZuv9Vi5nLl+s
BxtGAB+DoHSkW8ihMFLUvNZEnE7qtgiTwdSnGE4jEp1BxY7Jjv7zfS+pu0KYsTH8
8PsvVgDTTtIqSPxFHZiR2gWAEVh7MAzmXAL8JD35mnWv5OKSDu6Hu7kcwCvvHg0L
UVzCmrLIhTiLliENwn0X9jHrRO3nHOG6crALq6XbiNgprzod0r9JLZYptDVaq2eQ
8XS16khFV/owDhD8otmlMs12v+bsYA82ImDKq1ZLaQU7YBscMjRg9OZIzo8qLqxo
maffawPJpj6mzQTYwOtch6zHLMa7OX3IffjIZ3bQS72aIBxodu539d/xy7bvJXYk
pV2MOi5OkM1hBcqs7+RrjUbP8OZJwXFfaQvFXSQeaXRck9/+G9+H4j0S1NgYrvJV
GdRSF6w8zn6d9ZlwqraJdTMEll6w8a/oJODwm1KAOGZ+AYbuj/+m8y95aHXgc80Q
JUpnSdDEO+t8iKE47EOL6egoqGaMj6JTmY37vF4SJ76B7Vha5cQBBEgLnXncgyHt
EWniojcIYZhog0Rv+D8FId2IvzEA/2jrExZRLWC/ZRjwcjmaLP8dBi9SxGnjMpcT
D0zxRnGC6CdKMyv16oS/tJSFZNQD+TIJWZk6lLaF6PXXoblqXHedDpvGzSRb5D5A
mAOHDMe1BG9YmS8sc1QgbwwUMi9LSVKWValRmQonUhoAjNw5T/XkDMYzFil3FLOz
kP7Sn+eJa8FvQOjaRo5RY/IM5NCFT63Ze0fnAdDXR4T6UgjInLtHePdPzoaKGIiH
RwEvBKWfM+xRPhzoSKzJfp52SmmIKtuIoW1oyw2zdTOwAKuICO/OJ2GLfMPjCYOv
DGVnzkbPxFL8AgGgMlTUmz7B6EjMBeAqEVpcRfxKc1gIwEecEUbq4kvVV0OMaKJv
QfJnZFUQl4W4izDn8lbo7L0S1erFW0Xexbr21aqhhYVHVZksi/ImMZn7b0KiD7Zw
hltcXS/1aVRZSiOm9mYPKFORtOy/vRG1fWWbffOCqA4Rp6Gm5U+XO/W8aBH6Lxce
5ck3ttABySkmFRwF9FHAZv/3PWw9zpoY8uB/Ap5uYgA+Z1/6hmxwuamLaVE8blo/
JZaAWFx0GRmV4pzzeNAz4cIS6PXOMRQM7uh1CtFPztQjl/jV+mjFjnSWq69Tpw0f
GJjc30vzpTKoCG/kILpASv4p+aS1kXAyvEZ/p1GDNzpexuXwEXoq2dsYi02vaWFI
cholAxGRwyQ+t2J8spoIVHLLPCweA/eYphn3ZkshrO6akObo608Td9y4W9l00LDH
eA8ACJ54UpEljgEqnd0OZUc4uOpgMh0Tn7WNpR207e36PggItfmpnObDWNNPPBMa
2DC/6k8kcCwgfFYjPIHuWJMKTOnzgTIQAc9lwGg8O3yGLdaQDi4l/ZEKQ9wE1Xjr
1V8sTyGkdQuN8WahOi94RJDfDFnh/62DChxmCNqz+bmu910n4cO9OUGfRPDylUCH
guN47ACJF9Pjg4Il67lqgI1CibjjXRACIvLFTG+820PVdDCEVJ8S5l1E4PHNap1o
jHMqou58z5TmL4cQO+W4V/rNpiwSKKVaqUqzvOkh3Qzq81XpFIHAZOiXwStqMJol
fjjRIE9WsWZFjyyy+bD3YwmYG3hRUl7cG3fMy5w6vyHkOFgETHAezY/WdGufUL8g
l/iaCxxe9M6bnDpSxhvkKBIRm29RBwKiLLEyzd+TqLF+9ndYBJzpNkPPsFlGIETA
jVC52GHL2hnYeWYku3CNJZlHBwD41XOH452/0uWYJHEOjEoRdV+cbuVK+QpAu/ot
QbobqLSa4Xlk+tp99zdTvVetIPPiWpter6ON1iB6W4hP77wdfc4WgMZm+KznDcUD
wipv9LXvWtPutr54Fr+89hOUU5RyyPIIfaijbrAwtlLVNR1Ow/QBdUhdVfB9B45Z
dbH0g18kChywtkaAUHN5CUXwQmGHL6Qqc3d1lxemAsAn3dOCl/Qk3G1OmUQWQEO9
FBqwhuwf6TQ8NbhwOUOuKG8Y2drFgd/8UdHyzS9lKqO0Bvo4uuUODrPo2H0dwzi9
TO95dQ3aJHurctbwFhcDuXxNOxCxfi5kcookx/kPA4MxuxpxEvAUQWsm9H5cPfdr
3pUarZa0HBnuxQVfEJVPUMoyxbTzFDKHOLSxBWLshmC7+1MOjDBCYNqEHUNzcYc2
7ctIKLNhn5dinF4lXgqG45LnwC0yt5r+3Qdvay/baEgepxT11pVTIqdCjGmtB6Gc
FDmhLVPETbHj6FILvMg9DcFGkQDlXzyquaQGJkkp/bfKVlLKgQr9xv4bYkIdLdf+
cfqQ+3HFCkzxW5Vo0BPHcgrjU2nH5N80O2BTIGLMYYFDJtqe0WtCJxhRqLDi+OUS
IRdyT1VF5G8f51MjiWVVopIg84E7OtrtoMXBYZ5SOCTcOxsyiQrbpgiLTM3aKfrO
Kzc39xh+ZKIIGKD5hBQhKNxLhoEt6dcUi9xsRYmx3HQnZHg6Ryzb6Sbxi+tETjxM
Wzf+yv2Mxxv7xl47DclW19suHOQjvOdtjmbtblmDutbmLengI21KYiyOlnYI6S19
7w0j0VIySr5GwRuZC+dmEudpseSGkwctrYUSieDLs6nIp6NnPzJCxexJwGqQYofn
9cNSb91EuMUIr9FqSoLW167uaV4ziByRbPxl7s5G1oFalpX5Vby/IJxQ1i6bwlFf
1M6Q2J4EnrpvQM9JSPA/CSIMmoUS7qdWHIknSSRyQoNEcq3XeDUALZB2g8WeMn9R
uS39pWCXv8CQY39sbqtN4Nsm542jWIEN7SiQ9PcijKUfzWyn+s2nb/nwg31FgQrJ
Tq0/NlQFd9MnLcYkYM9Qy0dHdY8LkahiBfEikEh0LrfaU/48he8uWuAD57TFI5gy
NbeUhYKOkjgCu+Wz0EpXo8g9u3BWBlLLQPuWUEva7ZJ7lj4ffworSQA3DxhcAfLN
+x8n+btYO63DQV7+Nu8wPa/PoJTJAr2DNQdHOCKwmhZjCsLEPfqOQ1Ap7TCFy/Z+
tXG61JUbe06fF3yKupuA06wVX+vMyoiO9ftpM9X953i5OkN6cYc9ullyjKXmfRn/
cLWugaTZtCQOFK3sUdYG0qBlU0FXS/As+LUHsTx5Gh8HJ+Be79BUztRtjYdcMMHY
Kw209edKIwYG0I/zR/qxb8N5hlsi/QhWkwaO2TRt/9gQaQtpSGz2ELnuETMpvG1h
65s6kaa0PKuLEbnMg8zCZdDoEBpT68NfU8bmOH50L4T6OVt/Zkcdwp8krryG1z5c
5VHBOctO793c8mj5MZ4LcthhzwYivv733g7Tj3zhc0LekC/LQOrSP/hHdUYKmxve
wbmk29KH97P+L3sWxpK4nG6G2bpdI2uK85tsfjytwNbVJeBBJJ44GJ7CFrQ6sNH4
qyord03RggV9ZbZZUUGsmai0BJydSW/fnSshkSIzISANiVW1c1zRZJnNw6viAfQ3
f0m1gRgz8WVoJXcDimBb7yVAEJEMWDjfglRnCPxj+mKX2vsAu2LqZf8Fl0JLZe6o
C/BIUgSaLYojpAmVJu/rFDwE9Xawf5/nS1iJqz8xLZHV6PEdwwrIyNzsq7iFetf+
RIGypvnMUsuAeaZX1ySGaZnZYy0gqp6HCsiZsYkObf1dRWlsefTFgLIGaWplwxt5
6X/U4Y48sBH8kYNSN/S8PB1R39LuPT+WSFbEBftSnjabHRR2mTXZsSUx+D8tj2vW
5jWJPapoPIgzuuDz8WLXiEEFwJAFPgBNKd0wKv5uP0ZLGEKHwsmb7ObUpRofflNy
RHduLQfCkhdDENZbrBBmjbS05wCTusWWot7TKKqRYVW0BT9XBSxheHw+X8iDGzFh
Pkec+ChVfadBkNrO5cF9CRycCym1dKmCmPckGRtty4yvNFJ87QoGIYuWpJlqOijO
+Zdfpigk6gQw2zNBwYKihA4nBAJf6bKA3xXHDEDG/5aEODJyVbx5YDtx2sxFNRV7
T6RgL5k24u3gqhBJJu8ItAuMjqgUw7ug6pGGS+15TxjWk2g6OKp1RfVTIATiWBYM
+zO0tEzT66On/125Ci6VOGwAvo2EmLVmNepVQc/ichl2SKa7e4wLV3/+ri4BS2Hb
nicoQFnyvfoRGdFmtBgsUcMm2cvVz6xKhhl61tjzRejqvFBq0t21bS/vt60lkl4a
jgTGoWoSSxAfPTJ7dwuEJiDlPChKNIxJTvn/TWVQqXMZk0O12zH6zL8xQfIN4TYA
SM+sPBdJPij9ZZBvREgdDAYOhMw4TDJOQKy37PRrnLiHmban9a/RSq7sgY7QrGy1
69XMWxCXJai53ujeTWHW1ub9dt2M6IOQf02oKuPm2geOJcFo66uM3nimUl8Ol36J
rsnqJ1ZV7igt5lNxZLZnj2pCCEVSwekln2kaYXXxF9KMDBlVDofe1RDBA0drYAUV
cqvL2vS7W3PPxcpfipsOTiuiqrEtb1X+EbdQqvEBEJgpNKP2MXAH2byPi0in80Ir
bM4dzMUEa2Eib3N9UuZeK3+bJ5LjcB43UgZUwaesV74W9kfrgStezaLodhHlRFMT
5s/Zghb3qea45O2yDtMj83vjaVPTo0GqE4jUy4tiYbzqAEDzmxehbRN9GTjNJipH
7tJ+G+m47sJ+ysDbBBcGkFNWbT1a1Mp1C+GZLjSg/OF6mBXEFCO9+952ANUq7uf4
xRq/lFE4Zy08XCfa0/INA9ji968p5028oh+8LWrm8FO09dQJUG4xb0X0EGJr0z8T
eOGwFa9BCVVuiwIvw1RctYsdLL1EmBJDRkFrEEM9xdbRQ8zzofis1PHInRrkZZ2f
7V6GnzYzZTLcAIxGY99IbPk3QoYjTeZAyMav1xjkui8bRY95xmKAmCF8OUKGL/Q3
GVUs8biagYvZJOtTWhhR4nedfiq+LVUeTwXq42oyMXgRb1UKlW2ESpoyedRUrQ/R
HNZpFCIr6tSQAfq1QzS7Ou3maEla0wHZhxUF6OlAycl8jmHb7sIzdgsX+gQgw1I3
gZFe0ItbvPr3hPtKQihEc8eKdkeRPetvcGdDjoUNrz3V/o6dQsx9gRiPREI6Dwmf
Eo6ok0asL+dCJx/aFSrS6dGNYtcx+ZOS4WJBEsihLSAnu7plWnP6RqYKbidBlcbg
kpKRVwGdEiCMZtxNaztQGz09E5O3a9/n0qg8+3oRV6nxYsAjWAcC/ribtBS3YvUr
+PTNk8GwO8ffI0nGx4am9in7i2M4YBJaknPyQlhcD+5oI4kkETRxCo88zIm/62bB
l+z933MBlmgNSha5tWdMS94gPjvUg/aiKGRVGRPWJqC80MM9xioiyLkWAxO0e7po
j73X3qjOBe5CKiW2PUPs4gXfAU9M3LQK4EtnoYRGUJywBqUEoXixKS3zTV0kUe8/
mbqVvGYst0V4XsWzqvlM8aVCuOOzOTYjvbocRJhu3IMsmGtbZGQWkWNvhvk7QAOq
fDcJ9i2t2Cdxkhr1tvwKj9ba0+kxI77CUWJG4kAcyrQI7spOKJ8rzcKpmy6Ww1FK
ez8HCelnM84PZhVzezEXnEQezrDMxWhIyE+T192YXPflPDURaVSZJkd7lHw/YzLb
ES6zH28iq8GmON4tmkfCiaW5bpfam19VKD5ml64ohJl/XNg7HOIFfoSKzBMv0VeT
OKPq/evJpTykRvIt9+CVo43VAtKSuMWwI5lS/uhydjHiTHAh9AbrMMgY00fATSmO
qX1zp+GrAcRnLJ5yB2Ne9UdiNRt0rN+K83HyTw9QNeDk/cjjoVtaJ4zn5V+KnGPp
gXL7pPFoaq5kczJJswM31rcJxQNB2d0nZd150bjn5qaakh03h2qPTy9r2P6kQ+CQ
ldzvWHLH8xSAu2d0tNNkQOPd7TIGzWY89GPrabf7dmq1DXHeUKoElmbF1dd/DZ9R
mj3mITYz69v960SupDFzbvycx07xqPoTj4lQdTKotXB+qykGwhDX34VOuRd6U8qk
FgR+p+LyIa8x901tgXiRavb84p7tpo52zHJs+TkVM/qSJiihh/KRBQIMYD36hVAx
/yBsjYxHwKxg8QtCuEBmy55dM5mrolZQVHjNSpw5LDa2KNBDfN6cWUGjW2BZdGT/
218ZGsuY3j/CORYJXxdZ2WvTcNGvbRh4J55kqLdktz6nLwpxCAANfSVfjrRFx1cE
2PPBxEnDVY+ueAny4UitaeSPC5cNoJRsX9DJeRzX/qm8AmEb3K1vqgqLHrC+dfum
W/ZeZk/1S6s56SvNPx3b+RG86pn3fdAKVLLO1VRjflmftrx54MGJDr/ZCqNbdntu
tYfaGzkld5pfK+XOrSHVMpgxeszPT0zSkAsg2ZuPVyZCFwBCP8TKz70huX3Ub3CY
5asjRwrdmDgFVRXY3IhXD2GG308Kwg3UAG0ABV7sMRbrp+MR69Ys23wL5OIjWaep
htRdAOaWtUwpVo3uczaGQ9PHx1HKwjVTaQP8vqUYSciyvJwNqOkQNJQg+Y4hr1VO
cXm5hIjTIbCwjU6Dc4Yi/BIR98QqrTqmxpnnjg8zw97/DfAofT20kJu5Nco7u+gE
Z2+o4phDgwbcZIDtGBtG/j9ujEdLvq4vf6Sk2fPxFcdil/GmhlnFiB4gWQ6uOgX3
qleaX0VkBJ+xlRqWaoErC2odi70CZzEf08Iswh6j1VFkD2lSb+OYZYy2M1wLGkwa
9+Z5Lv4Awcm/ygpRcCOdwgW4TpIGsuDYAT356+9BygDvRi0mrpg0/hEzG1aaxZWN
BjN2mrgiOt+ilDuEiSWnWoJPjrKXOkdekcC6VuN5TnIryoETopRkze7CQCgxCHhS
J4nIYNkXf3faYV9lzy78TBxr/8+Oo03xrByWz2v/GAedg9dXjAb5ZWD2OtmUVPhI
WgcMNIsq3VhdQ658fVXlB5U5YoLoYUq+1JcyN/Cg165SAyc9KosmzabvtjBJOy+k
9FnJADui+ujiQau/55bgqGMx8mHt4jxip2fSyjDK9FiXG/SgxKV2/Vfs/Ff40KBM
Y02X2MmxBbRHqYI5KIFOKh1VUHvI+98G8bHSuh7E/VynYzsmv4MQgOKfYepJK7DM
gUwFLQTczUy+jwS+aqovdxVjF0xPli5b5TzjvktBK+U5AnOxlj9Armd/UPflSlHL
lCSlArTA2Hk3O69N/Env3GnpFJd+TCwy0ZgqU6/lk/PND0AWYzoOxSfL/sCFwSyd
RuNyTbfyLXXpoRa4cM8RjoQjqLR+dsSD9muqqHjofHAc3U8vFsZgv2dmw+ocSvWi
srjzZKfx4VF6LxKQ/sgTuIAPcnmWwY0J6Dais8hc18QlEuZkBQxx/uEZ3w3ho1xm
l9ryLeka3Zy2I2XnLuQ62VISIFWr/Pp4l5FjQtdmZWZ0mRtP9MmILy++5U7D/XfY
QSo2mS3pCXLI04zXgc9+4qUG08tv45vaZkekai6AcfdF4+Bg3BfE+z9Vzlu9xWiU
qvzi1DxGaPQYA2hxyNEXgkqlHWKJqiEA3PTgzF6yGXKrd+k3qti3U56ObbtD1Des
6kvHZJlxP868Dq+GxTMIrxDKDku4ZdlzkQ0m5IVVMLB6bGHKct789m54F4MmKn0l
28ceRrnqUcssYOXJzHX/JLnNQ3Bid9ZemZDFS83o9vBma7KY01wsGxsj1MOwzOiP
4/GcliVQC8HTJhJC1BA0qqrwe+ZQyaZ5SI+TxKaW9hg0XbvY31MFKZ2ctRrdVjyT
BOxICDPAiV/bkwBs31OcTYxLuSf3I8JfhVj/eOs4oRH7xRwuTCxohO++i7QbSLXT
KR9+R5PH5RJds84u4/j1E/wD6hqnrk1FZ+QCvC8w5fdQzZTQ2Dhw5uI+suL5kf7U
HoTAuBe5uCg94uNculbKn9i2vEwBdXgAasb36vWgxhf0/WtMblSlpu5f8VW6hjs+
oNdmhk66au3KyLrn5fgDEwLcsivG3HG9rKiOWmWiVoMSNuhlK8H7usMrFkdhGPkQ
fHrcQxaPDsTfHw7ZLE5FaEA5t/cBd3T3hW5OmKilpwP17GlolwgE7EBl6HvPEWKd
7eoCDD2hFYDkvImwkx8JEQH+49EkU7cJUaSH3H/rm2TE9Ol9jgIpk5OGjnYbFdfz
sGbrPkyNGDF2EWA5gDamzjXPs0bcfQkYVppuhazKLaVzR1/qrwjKm+xNIzJVMwmI
o6d25iy9A8iYl8XupB6HyUe6o13taLNTQa9Ma0sVbifmzEtcc5bE5pH8wIwvbRen
cbbMSP/Tb1eUUdZddQDzAYxqiPZ6em8pv9nMLoiU1T2Vhg/M1rfujhWaK2ys/ZLU
CYCkSBOubGNovG6FStlfpzW586tP4IV2XH7RwmS11fVfCDWkZ+EHNEmXtxJX9Ttm
AEUTcIWyMZjOjL6hLTqru4xApl9PXjLKD5CCqjfXiyiOMAgvw2GVAt3N9eVpNccC
6o9L1uYoCgh18ASc1UJQFjcnQX0pqB/lfRtb03w0EcvWwpQ22Su7rMypyi8EELQ6
4YfTBZTN3MOcszM3WZYeo4d4SFVAQMIQOCu1kvzuqpR7qBuW4SWQm1an9bL9m6GF
Z6umXaXvlW3fbNQ8K93qoTF1CDEVPXOBEVIDUsRlaQKC1B8vGvwlp9nsQmZzOHy+
193tGipPjZeSZyVpSGAQjtHp5uARB3pKZjNHTPdtH+O0fkRG8hSizWCwVjdoYpFb
4krlEt01PhtKJHg4NqkaDmr4eCozE8o6qAiv3kxGJAhz7joCkmq9XMuCyR29qGWU
lVAGCehAoF5ySklqyp9FHd1NNbNET9HU3Hd/YMdtdr9ZSXQ0HCk4ltoP2Y0e4Vok
GZ9fzQlfP17JS2+/L8RWKMGjaHjWRu0h1Pbxb1lRau40ccUU+eHVeO6FoFhI/5/5
HQxn3h6W9wa/bjekULv+yWhx8GxNFhcib0/3C7cHePBhIN+wlzSJQePA0kme1dg7
PHWHcrzrnK3+T+GcH2519CvSBjSaXriK1HrjmsNrLIyy4If2uTkcGoTFke47nbCS
TSsAMJsnAOoSlqZ6IjXpWfOjuvhaxBr58kXfUxuMnoISr3rtsdjn5jlavzjoFU6j
UtX6NDAIG3FPdAGCCWxVzBO+HCXooGiiZpf8tDToDSvm9HGlbqpPbXNNC2+6tDfx
iu5Ea1wae1LZRBvJOuERMZUgi4jwHQiHRsekDlKLUFOKMXo0+NxTRavo4b3k0/Iv
T8UmZIRHU4g41SKSFkQKHhObYSDzJlSsc1D0n1R/ryBTjh2OBNmbAWiXo7ZILXt0
eB7QLnlfkvhDcm5N/8LYZ/8oeI+nva14O4OPQQ2YWO74H2pxRs4NdjWT8Wb+AZHY
SMo3b6WxitQ59LC7d47rzw6yvIL+0coNFFetnEj52u6audfIh+LsOMTuk0K6Gqr7
+qBPUkenKAFRTOeQbAfxc3QpmnSvSfodViCXg2O5veVsBgd9Qu0vPpLwgGvn6QDv
gscHBayMQbvflBTgIVd9zl58G5XKWsngZNdsuH908SzqsekL/gmqclsyxY4MGS5+
fA48nifHdIi0mPptMsTmeUQ7ltdGyib77pSkdvmHFfMtMgrrgZsg601LRoxgc0Ub
eIm+xzmcQyuDa9NeNSsRaXL5qnMkARX9I1Ix5+UYPxBzq+ztIspRO3hCxYWxWpFT
PURUK0NfpKK4FZQMyZZA4y199IMHuqAvklESyFxM2qoBGG07Hrf2OjPmg9al9dxo
TQfHRNuZ1E6ZhoJDvBYPMvYFsUCJNY8tR0KnibDctflKB0y8UYtWVBsW9mh+DjKd
ssVVgZ8ewMGQs1qoBgnqHf7PxoKUuDE9e7knQLC6NSgKD1Quxai4QCRDmWaE66Yt
yLq6AH4l+KMC2lMmnIrch/N7z08BGQPrI0I+zMXNpmH27AufLg/Th/ZzBIAwK0cP
787ZENAzKDMaVOo2rVrvrmtzOCTcV1l3urHa4T3vK0uD1wmZGB82alUWE6BaV/gf
A3K5IqJH23l4NJSItmyrVOPb7t+fMC1i90W4+cvP0cqh43RMckPGKtZadVjwdAQi
EV1doZDpzNIB9C6VXkeeCeJeBBOezwsW4VYTLD5ziwBA5sDjOfdM3v9rXYMumWU+
pOGFUCVfe9oAhUfKGYcTENshDR0TkNCP8ZWi4hSxiO/KEWJRIWZsVksj3aKLiCX7
Wr8S2YF38IhB4sQk7GEqmhBP4WhCWCKjOYXzgV1jgipYAebIRlElyZFmeBsJLmT9
kWTgjWA9qQ9hDuv4tW5L+4eP5daNxdCuc9xYsjNBXO6gmCXnCvGwB02ykQ3lNHY9
gtt+ayZKVaOTIYH8qw0OXk9Pn442qrWGiVRSZEWA82ON66LPky/vkt+3hnl9+zr2
dxoszbi/CzoAXltHmdw9v04C95vK0OL1BHdC+Qvn/yBJxJ/l30/sAN4XbOGCi4uD
JlppWFdkA4I7oX2t5heODUG2yNAyetdKoCRQxoaFg2e3b213wJFlb0pAhQz5SrxL
/6ocIh5JD4LEDj6ftMceIQqkiV+gbWDk3Ewx1hrv3lIS9M0kUyX+syABDvq9SydV
K+BMCNylgyRA++9+X1WFrtC+m04yIFhB1+ujcBgXM+x23D2hpSZwWXTLtyg4il8A
LVzhR0IUZ/lbC8iiQWsQaVjwDKMfSnpeL/mLoSh796TAJfA+4yOGtOBZid+MScx+
tu6/HOTxhU+y+1HlrLSEFv2Vf3nu34xd/n6L/UWh+SpUnmUN7MdnnTT21/SUK5WL
nLsSDO92dJ2FbTkSk8BSONdDJxcnlRBs0VGZ/oO72SEw3Zieuu76e+TyfMRaLl41
1BWUuibcBv+24317I7fyQ9+LB8XodwuC6AsHvHLzq2NDSZph0Hfrw3Wsa455P8Ic
fdEDhu00j7tWuMSjfyHdIncGGhLiCMOdLk6dknRXqGREVTbDxMxTHKGTuj2YCMrc
OFBfbZEaWNCTKxedv4+yB4z/jUQNXF/N4qil9Kcvj6jJFVgUDnZJQuRhSgVedFXF
hcSv/SAX6AYyI/EexqMDKkRLpKx43Cc3xaXiyAxlhUbjrc5YQQ7kKyUive3/Bvkv
ImuG27Z3HXu85BpBJpw5g5abTxBvYCExOzj8fEt5W1Bmb2JbvFQb5uomNCjONqqk
0laP2lAyE7tnt9ZRUiDnYRroMPEc6+okN0+qcmORjTprMG12IZkC5UBKzPcE2LPM
GXtAX5FNccOFYGd6y0aRN8N7xfZnEP0Seh7quIQ9aw5Tp7DOgTztofUNwOBhZCsY
ag6xu49i66tFwk7pxF43VUskPIGXFtd9628nWtjpXdWLlpmRkeNQWAeRJSA3ylbB
6jXSygue30/Seh9tMlgsyzXm/w67TeXNKlZRjEgQIuvKlG7PJDN0yo4qv+1sYxwm
Z01vMPLSxNm5Ci3TWO0Cf0OsNvJeuocXuE1uy7PD3Q1oKUit3AAGH6wNnqB4gIQp
L82SWdlC6Bfo/B+4XpBLzLHfabjp1BaY0s2CZc9Nm2yaSUGUFm1ipsot4//WkXQO
zFPIzNnZveKtIzFUkSFFPDzV9zKZmAgYynct2czuH6X3rrFFKS9q6pD6jfMfCKhP
kGxYCbFmr2RjtHBcKIO1dt6IsHTVYxsAi+LELdRjWxsQ3VDo12VoHXVLMDUuNE5Q
PDolgAHaFd5LQpm9SregXm821UjXH614RbweSRkCT0z3dLcW0u5FG5ai5D7birkU
ZjxKiWeR88fRxW67392YGKGOZBapcR7ylkANR6PSRUmiw62MUZciz2oUNTZGEibz
fYjatpn5pYqUm73PGQuTnmSKyhowUX8lHb1KbonOtmTX5k08Z+Ow09FGfHPtKBeq
W/amIE3AU0YfxlWvsFA4A23kukMoAqNf3hShD6P5WXluwWsMAefyTx7bT9rbQRx9
T96XSBUuohRjDF3PrzSE9Ikg7oq0lLdqwPmjZKbhE7kyD8e9azzQbMmSxTsMao1X
nhhLn3u/vmWqakTpS/g3VKyMsO5VuWaXq3ZOh3KOszCtxAaisLxTV123Vr6SZKKd
LKDvidb8iBqVJJJVji2b6/VisvsqNoTOgHxmE/Q+xz1X0JXeyhuHWnivgPsxKmw5
h1u3hRQ9oaXp7oeHhXYI5zyG0NQhKI5DveWSRmoTME+3KcIm4NTlniZLtaXF/Q7h
yboKml9GJkgLttr5MWA/29ml+vKNzMTld+JigfrhQohjD4+dL2LZJEaT9cC1TDFI
ibPxjgX0NHBfmQk3DRCU1IUcuTv8gz8c9msQ7SpgALw0JymWiTywfoTCplA91xRn
C3VoOQdQZO3hVrgj5XnMZ9O3kR9cndLdHyYLxzZi5KOLMBqDkFBgEOGa1nr2mpS+
3f6fohfhNeD0AVA9C6bnwEU8N+qehaTtdWHFDM0pYWX9lHIPAo0bB9fxWf8dCzwY
T/+jc69kVN6GoN7Hu9tGlppoMnQ9fJMDFqFdmXHM/zFHDVL5FEZ/8VNvS8LDv9mE
v7fiVKV6tRNnSf4vNoJSODdEzT5agr1HJkVD060+Ft0pqWZo+yaK2Y79fYtvWZEg
UDs00wFw/7ao6y4s1SGZUFI0bN3G+y/KdokRFlNCVujiyDjmS5Vw/rvUZkOZwMlA
oqlwBzq8ZnlvELmAzPvrA59JtrkpUc1aMwdETNX4xpSmBeRPQ3TRUJ+xMOQ5OTrU
LcA0p+S07nGH09X4hS77pb6a+KEk/jS5MOWq3jb/BwDT4G9u/yhCBbT/ut/sRYEM
kHShMICWfDozL6jo3cNdjNlVJDxLJLwgEBuOjfU0r6+VSuiDPQlcD2RivLN7Jg3T
I4e7AdArszCrY4T7dmgopjI9t0UZf+C2JCDPmaEZZpBiJnrm02zd0HeJxkAZNZMe
TGoPvXIuaC+2n2LKppVcHHMegAghfhsqEezg7y5xrxccQFE1FwVeiw0JnxRcyUA6
qrP/ImsdgU3jQU3iDBcju+cuoMEGBc3noeOVldvaabfTSLQaD9JOAbHaq4vCRp0a
BcS6lIEehA/PPQftTf5vKLKQ1qX+b2OMhcK/SANj1TFFQszi1aGmVqkHYXhlmjkx
/8+2Hb/S9fgQ31/uJXUVnflaLz3XEvKGqAUrR5laRHCMMkOiknfU2BQ3hFywUH6d
yFT9vfQ0atRK7f2W271oO+yS0aguWzI4BeXuW6ebsztabf/JcYt7MEnWOmLugrWc
82SoWVEOGsaUPcSsbBowg14zipLJCGV7Bux9rS4iQBolezIht0/fIMOYhqQjsPx9
5eBk8RPQW0mQhbLvpLYEbb7Cw4UWilcBIEqVS9MTw8NU/MI6shp7osFxt/3KJ7FQ
0Tlf7jtojuvmD4piFjpjD6GOIoDHwcJz5TBTTLpsAE13j7PV40XlkOZ8Bk8DvBjm
IFeeaRvhKlA+7CnPqCv7zIWIDSY4YZEPkXAve78t72Lxo9zj0LTThZ/flzzyCzqq
vfVLWEjLvr/KfVYOS8wn8JCHQvAVZxGIC1eCNzag6qJoPlISj13iiQNkb7HlrTay
c66rNZops244vaqTDDxi7PCK9WNPalRi34xiHeRR1aE8bDO7IeyxYuzHj+LF4m7R
X3v4emyR+jcFhNY1nchBW7q4NRF07h/MsNkAtMZ8XeeZVF04WgR/LWTV9Eg5uQXw
ANfhJoXulB0eop2/UbRNyr7NwMnTP4MWcKnVNmkAPX1HlJDKHas30MMzz/Thxi54
zWUA5w/Njfhhkesy17e67fyoXuqZfPo4frS4hgNsNCMYhzn5j9aen2BD+vgra0bY
iFjaUzuiY+YuCRuXZzezolHvxG61D+8ByZNqSplntkFaCxhasvYnY6CJvJd3L9nc
WFGemdPpZmYx6nFhCUUHuLm0LMPoyK1Cr3jor9zsoFSDPiRogIMsfK0IiYXmpzeq
krV5qh3RGvq2avRtGmecmFTA5YBlUG0c/Es16XFSDtNx7ZA1vYBaY+kP8u2zzf3W
FZ3x/JytrNfzXTNJ+qzSXgcosA74kjkOtDZI8AtT+sn8qbmoitxm8HlSADH1nj10
hvTYtFdrekT8Py+uAoKul3UtHqEwymZRMfU+UIOQ3wFhD1EMwTqzD2pkYij/wQOG
MD7xoTEPGcfE3t2vaW/Q59kP0lHDX0kZIMzokpgqHB5cq7CThhvJ/9XgjbHUaFGD
dUPUpdR1rKxswN3Wjw4YxyTALX4Hnm8NEPmgKgJV+OxuLjpcllZy7lK1UwtmMcJu
EgssrQWCH1Wxq2m33VWw6e8C2kHxrkxf+71+I1vBB9gCJ0pndEvy/Yvwz9KeIA72
gucpUJo2bDuBteOztY0G0mAOl2Gb1TNHQLItyLtY54yAfj21t2rzzd54PdvjK5pU
+tOOrMYefjTlhXDxXMtdHRQ1HLzJg1UdgwSBfL7ecMGTYIPLdUcgciG720bdXkzL
kao4BeaG5wS3mpBKvMoXDLdi4+YZo3+8iaeK5gyb72s4eWLWzwvdFgQgMZYSllzo
RcU5xBTo1SDXl4UP8ML5reaLRReYyho+n03yd53Qm5TUefh3zDWoCxj5fLr3ydu1
RKt7cMGkaSsfGMC4ak5zPn7UoyQKBm8yvInikh/LJDqEiI8LlnaJR/BM/j1eAHpZ
M5Q8xzdNDKtiEAA6JnqoJaqw4x5NDpvOh2hLsOsbe/HoYkpHqmFcFiuw/+tuPsQU
hCO2lKVHjfhtprwJsx1nOiVSJ5l428su+TqS5vFt9clKnP19Naw9b4tUPNg7gjrg
OYrkVg+6Ual2QdBiM0Mby1DFQr+E9HadrrJUJL9F6h/pfL5yfXRrYi0aRlv0UEun
p+U/p3UI4xBvvpc1oTYfk2cWrsqVTFb5hOuI49jKqdLuSQHVspLv/i8Zg+Bnd+OP
2E3nDGcfvnuig6ISHfooeaJrEGof1jX+E6bL6mNkxWvP4Y1DkQh2M07mSoV0W509
zlEv7KcR5CmkY3tpiO/gsaSRkZRqgXqCpfGwKgYfosdi6DgMNfNhwaU4o1JEFo/W
4YXpM2VdRZP47FIQFsq43M1SNr/Bc4TKWYKzorfiKTZs0BZqfxIb06UDYlq5SOQF
9Gs54abFrV3NbEAx3wFZFeSy0jf/R2L6jQHzKms/7Vs2YP2VWqzyNMZLbiE3gp6U
4+5uo+6dF14tgZaxHQpoRR+ozS0H4EcKbgKwfaLVouO9DhuDDFxLM3fAphPF3z2J
gVnhKoyGi458E5QdbaX6EBwsrU2jP+OZdoaWH/jxKJi0NT8ReYq0yRR1yVlCLC4s
kxzcJTPZ4RVY5ejhd+ikUPJ8kNbIDPxZPgUtsnohHoJcqmk1Ehk7a2vU2vIIUda1
QnrqEM3E5ePf5sARf3AHgLk+lvfHTVxz2wjLsv3vp80WSHu8F7FXNIwYjsM79wxJ
Hmxv1FaSTKvA5/kmGa+uTHT28yLMHXNYOZx05mddNY8mJL60Wvo+7oq477SwaMGK
prZFucCSp5oq9MKDuZiBffq6s5YS/sjFRH1UF5j5Ndshd1eG5Tw5Jxi8dTv+GtGo
pKDwP2r4JByVmco1IKL2Zr08HgqUHkd0DxrCKkwCoAmjM95IWbLO/C/Fc9BZuhkS
0SKPh9Ny7VqbS4oG8vyBgpIdJ6UiWaTZDAIbZeG1GP/BCiflWrfwtZtUN8J9H8jk
I0xL3YdMzXgwRD3SZSkDj9TfKRT48BhWq/1Tng5zdAWfexlkmqEWz2nwgvMBb4kR
ejB9xE0NatFfjURxOZEZQCfzTsy1VbbjPJ5LzF+PlMl1XHhKiVHOdBq0bvn6McEA
5rBtWUYwk8ubuk3cEra1V2jply/GiMvthJQy3EHBamxVSEIKg9k9gBeXbYndq7jl
qklnmiLEqMjCMu0PgXz9/NYPkpO4HW8m5lOrGYvRBFK7o2GdEsfaEyMu+Y43JyLV
SB2Xy9nCe20zMr4YDVwiIHntPrka3y/LG80sbU6IO9VW7bJFJuIO/5K7qYkct3P/
mz8cffVFN+UMDG8AR86Ahf6SQLjZ17lTwJMrpp3EOjhvH6A5G96XlOb3aUnG9VpK
XB25z4dvPC47/MvU5CH3hv0DnAAn6tgeerePmDqfdcLLpDWQoJRnHYaKqYp+/0pc
PZs8RUQFjMJ9sDm/6c6yBo24HdW8HUFsHz5uuRcwTcVaElJYQOJ5x13J4kAiBSBr
jLgHKLDp0IjoUqGlebTWEPZf6SS1YjWdUgvxsdcB59bNN/df3sNZwo9mjl/FfMtz
EW5UnZIPUdzfJICHgTHN6Hp/57FkdyMZ+ay43AI06Iy+rEMLuIlg+nFywVmy+lRJ
pGA3DaPTERZqV2W5nrprcsD/MZepLD5FjsDCQOxsm84ZSyONVwd1iaKEWMMKO2QQ
+EfAHNmgDlukr9ZkVomY3MUZZG+fyAQkozYCd81RFmd53MHje/JLNTQ4a8yLepf0
OjkXCqIA+KWD15y7XYafwmPsXuA2bFiq0jExtJylLv5ur/6X4G+EP65o5DGn/x8Y
w/Ackz6PoRrhGSy1K9Xve282ixnPSn3wkYLgD7yZa0WtV9C6R1D6hFmW134/d2ed
nulqDjIAnSI1CsyJemp21h2EFgT/doxDLo4cWJtTzlIkXW4EEVbqcbMwfro9jRcd
STvgk/Jo1iZhW28f7BLu4+rPbt+krvOQwXcf/Rg8oJuMWaJ8MQzBaIADsZooE9kv
4yYYF1Q4Lr0Iy/knzWqCgKACoBx7labxpGOpYfs2/cT9M4Eluk5XhJvUk0ZmAmpV
lN4qw/EieglNTGS7GbcvdTyxDMaj/Q0SQXcu/EiIMFgxmPk+yCy0bU8c8kV1E4Xe
k7To/5in9ACd4tkhQECdIzp3UdLOxttMxhDK4s1EF3bIqePQdwoMnmvWJw4RgzId
UQFFwgpGpuQ9ufKfLZH3lvNcRZTT6db1Bj1/9FiWe54AQX1bVpuC7VsGKOAPif/l
7ySC7emGe3VGT2hY2G4Lw1TzFD2NmeH9UCxR5Kl+SjzQgICjk+wiHkhGYGf1UyyP
S7sWbASmfreTem3RL/aq4Z6PGNzgpDdDieKPuysCXnX8jA5XWLaERwFkQkRdooXz
uwEpIOs1rW7sildeSjr2vKR6+NAidOQU0J5uBJ7rwvpKCn46gbRk+TcSu/Duujl6
wo2tvyZo4egCQLda/Lh5Pr/YgilykVsi1TcqSDfLz4zq9B2YDMn4RApJ/xLVHghm
Aq3CCV6fKb5w+9Ovd2j1N3SZ4ULuPuCQZrG1Sx8rPJR9GgXWbGfUsvmOXF2MHhrX
MzQl4xos6yfryIeHd2bHw0pu93us0Gn+16Z6XX4Pz5DWtLLffUKWZbfWR8aDQadU
+PlZpmfBHXo9xnKwtvwb7FJzSbi0tvSTM4WLHntqfPUCkZc7dv7h4mA6RI6DPHmZ
yxouZ3tTrkJvhdvY30JpQa5U/u8zDLLtcEs7r+FOQKjzdj12nBEVfik9pKB7fJn4
JoV94wuPyoQWDwhG0PY/pfQMT/GyVWAr25YughttV8iH64gJ8g7027jl0Zt49igH
HSW8DO8HsgQOJPgyPmDJWpzOC4ty/HuL7ECTW047sL+Mps8ElyDMpQv25avK1SYI
9paVe/EEAkKPjfw7CFsah8rEmq3O3+sQP+ZHNZGq1dGvoNOvYvZe6kf4vwnjb6V+
dqCjaY3yZ/Nk2iOgmljxsBFswQLTywLekAb94S64IRQfvbjvz4iYTPZecO74zRtN
eaXNCyB80//rf2Ehe4GKHFGcJSxlmjludlgzeK/rVQHXiKbp1A49JditTrp5aS2l
2oPVeYmOXaUXh1fHGlZhQw6SegsZ2xqroBQAY1Qm4PM1oFFS3aluqBliijOF0Xm6
qNCebhyISnp9H7sPh5TMjZkRtZ9oJ30YKDwH0kSyHx4TEEAryeC8Xd9kN5769O42
RdFfPVqLCu5mLMhHwvJwvsXNmRUunIsFri/0NEkCsOXgXEx6lHk35j2YcMD9FcHm
T3e+crq98v1HYwYwSNwmL8qV/mk3KSo25L87keP2rn7H04UnEDH0COF/7qEIySZ2
Uv3Dl9JzakPuZ11QHXR2oi5Fj7NErPC2OI1rs8cB0TcPObbHJzDNBUIO2ZEMsnAQ
I2iQVRzYcCDRxY+7+0hBY+FJRDbqWkoECFbOqfM9MioZUm0piNlvJI6vdorg6Ngb
g1iVJQlcnhak4xIAvgG1K26yBPyV0trUiOqqSEqG8JlGJEhs92Zq4nMfdI+htLRI
CZqG2Q3ygjDKbX+y7J4UHaOWf3k0Y5GuYN8GUyBLtLM4JlvHBY/3ZrgfrLPkynZn
MEF4ykhP/vp/o1AKCwBuieMXSVlebR35wlhdX2SK05KadnVpYHFG17DW4A4QWGNo
YZuGSQqp7/l//l83O1RbPDElS67oJByItQ1TBx3NzT50vS1hK56hL8MEzhrk8Vgf
yJrOlh2l832t0pu8m1/Cs/qCMqkcci9TveIxpWZuBviUiBuNNCAJw3Qi2oAbR/cA
rsBKnKPC+Ta+hV/IcStiTD1I73UgdNjCh3FvLzKr+usKyzfgT27nSQbI3sJstOdR
/W+4qRXJla7z+LiF2JLZrpjn9BQuJcw9bt+Sbpw61VP0UOiC5ybmRNEtaT/04onb
SvO+EHiItlRK1SEMkgE9WtIksymj+ETsu0lnwOmKMva7amYCJnssDG26fds85Z1L
yduMXNFb3Qf3mq27gkkntmLRmibXGIJKY7g8vR1Kvx5rIE0jUcSMicDdzOD8DwEn
TvGNe1shxa9xlaPqCY2bhT9h+FJHc0YSWchBCpxCBNORoJiHlMbWDTyFW97O5LdR
XDx9BCqmbb8SSxz9RX/qMtDhA2qmYYBoZWwTAKBqZBKgb1+pKReKcMWSM+L7Qvba
jde0Hw0PvLN9sZ3WcxWDod2QIMKqGWipzyu9a+GYmzFQ4aXpkY+3+NL8WW/7g+Qc
VlFIfEZeyRcY1vDPzBcmEfjZkyivYVTyIrjQBEb10Vq+u6t1UT+pP4OAdMvYu3nc
3bk/PsnoI/zOHp21TaXFZO0eoxVMjd9cyU5JE9HL5jdvta48F8/z+J/07Pn/RT3S
GgqNDg5sDWJWxV2OeCohWzv55eEq4KYYw0Zkk4OFDfWNO5qz774Qy3EtWqdiheZQ
rSbHJw5qd8A6MlY+15tKgH67myjZMI/dn20TLPYCdtJxMK4iLVOEkmhGA5a7zqJ9
HQITRcn1Rj4bhLoDypTkBXXUjkItFXDvoF93bH8fkayMg0p42y7UywgThAppimpO
DAMQUM6xiusNEflJeV9xkLxb1FBaeFteM4qNAbHjokYJ05Je1SFeZ/5ZeZYj5HVj
7CyFFx42k0sifIgVy4NR60wTe3H6bzIvsi1R8fao6gRMoGGb/0PybilgQ4v4E9dC
mXn4gfU8HFOiyEZqHnYNh/5ynhyf9etj1OeAQza1MsmrMzy/n6KqU/0RGyQC9gLN
CNSCMSlWLCmoLLztTvRGzXp7AnuNKRr/5Hx9x7dx5X2MZYUXcdvhVsnqcoegpLwj
W5cQcYJ7Nb4wWC2TJofpTO5YBhqIjuMIqZKjxHRpZGFM/M2/mk/WkUD67ItX5caC
2toJ0cOS2MorCR+zMzXylXBgmimbUW4w0aq199606eGCKn1Kms9N3pYI6shoPGgb
HIkHK7uXUub5KHc1hix/vVTvjh7jDN7RSZXCoVpU3V7X4EIso5AgO5QJ9qfBanlk
G5b3+9FMtYI+Z6lJeMEDRaO2KwDivekEUsQOHc6yyaOH6X3R42N7U08lC6sO/qWl
TftKLVA0C6hiQgcWVnaMVzq+34FpST+qk81fjeNrtQt+aPTKder80qBf73GGMhv3
EOk8gstLzmOSmNPKAAqt4NEiWJaTsZNqx5AJzGL8ZKNf0uz4n1Lb3a2TDmL8615+
Vh6lrD2UTlE2N4EMZtHQAo0c3e8EMLL4Trlv6iYCFeKvGVs9C9J8l3T5PGp/NkUa
MZoroI1ylxfAAPi9zDIMmz4ft8zwC9s0/2yAC0sXYHcvFs/8K779wzIocmiC3Vio
Oh5zFZpKl0DEc24bIKeMsF82Qp3tyYkMcTsvobW3zP50we6ViQn5YGnhjttVjViD
54gxZ+/eOsvfj8A+4IWwb3+nle1jDuDdG9vBAvwNHmSN86au9EzQD6j/1YOjQiAE
BvTau47lo+4uykSJTeDXyylnfD/Ka1fh/QnDkC/AUXoPYHeRSLHJCTexZh8X1V8C
emU0/XOKHuJ8w/dm4h3L7a5/J2TyifJ//7kJW/5gSqiZvtC0312ySAb9XfYr4QqB
bYSWl3pyz5Rj6ZvtFXaH67duKBt98OBbJcFlkjgQbj3OHjz+/K6n79IAeucNGW6M
zhNyjiNLifaNmfJXBFILenmhC/nf4ohOWDzposb+vedKigc/2Uiy1HIQ4ZyLsxc4
PzQHzum+EABG5nnm9Qp/Qa8qhBRy1GLSimqoiRIViGPWnV4UZrCrD0uVX8VwzzCr
dbUxTWJo/Spmk4ADyFVtEs5rgCit3lcz5+huzhxHqTuuWqdh0UAIUkXhPzWx1h8i
8iV8rsZEwklfe4zFs7vJf8L0lIL+FY2NKeG3aEFtnxrYiboFXtv7LFi21UgoRKQx
zHbLGslhcNnNWaN2gwepT1rn0YowKM6PfGjXNKsfHmL/tZ+mEoBp0IP/JWG3Pr2M
nBRms1+O8dD6gkjTNqYpQQqdazDm58ju80+tFEIe/wm956ulVpcJJVR7+3wmyauP
ScYpN0Ns1QVrSF/lNo3vRQ5Eya97MJzLn7r7Gnjwvtd8wI3j3arV86EyWURadEQ4
vScvptlxBbuhSzOxBg6H3GU/6QvqnB6cofsBpOIySVq4LALkD60DAgkGPezsQdvU
RkOQjsDilmUhrTdlEBl6wcENPJE2kqff/RMSHUTyYQR6BM9yAFvi30UrIZTjWtlp
pl3uBzV3x3Zp2UnVobL4URaL53K43NCLAC4hKaB16/0oDrJM1lXd8Unv+5fm+CGi
XRDu9BiOfC3s2xHaOUHk44/Zfb7M4R+L14uMcVjqKa2VmccYDGYSWFXQtQkt+AKR
/ePK2VJPUa25V3uI5GLKq+aF//pAKxlJ473R83dFCLj1odXZjeElqhymqNOUvbml
F97z+bqyNUetRBZaI1HDep9hS4sCDENa4W/fn+uo0UIdF0PRNgYlFHgvenzIr01n
cs8YuzCgkXUpJWQW7YMEg+5cdR1woQ1C5/dFOTTxnDgFzP1vxPxM+BXbvXEJa+Yt
G4Wq31QJBwEAwk5v5KjkXlteFtv194G0xUFq6Fzlm/xTaROrRe3yMC9eHdVanUbc
O40r81CvVePfaO17bRBvfHjPht4cOqOKKiuvSeE5mcfLbMsD1P2ZzfJ0ag14n68+
78j64046NZKyzZEe9eYvunhQ4avr6xQkOw1JaiW7kXor9Lwm/n1XLrI7/PHQEpuK
kgEcu8cCGNWJ+afnqw9Qs8LYHDWWhLzAS6fGTFGdo8l4QvmHueWgvfh59KO84zCe
/ZmMyA9vxCHv+IiWTcMlVQizgLL3BeHTPZfwbGBxZvhtUTJ7QCuQBLldDtq69ljD
OnKIhS95RvYYrtx+vfUOF/ki2xvgdzDXpsNqhDqlKvu91h1NDvcoLqJR4xyZ6NyQ
6HMDzvc71HlHPLoH6G1aagKSr0KjWPrMyRvaubB2nufLIK9+DrbetZTl/nEvUizr
QvJ6kuucAPAg4rbCu13LiHw4cl6IemJxDTF0l4KTqKDU8/CEGWt4KF1wj15+bt66
95cu7TUcyYKaiD4elIRHRXAD4GJSnf3611LhwoQF71dzHtYs+vXxhhxHbYq3gpRW
jx7kjVoLHaWGaBDGTVrb4OSBtEbeenqHsXwb8605X+ByzeS6hBlPGtn7wtpXGwAC
jft4mkNF3OpK2gMcvdoqy3kx1QBj8nDk/mu4TumVPf1q+vEgHSZYHa+fYdvqZcyf
zu/r/GT9T0gBjIXJJcC1lPwiOp1xr129bSpBS3D24dZuM2Y6PNWRJpzKcCkf70Nh
u4QvEaKkpRmGBozUje3VOm1jmu0p271UCr3d7iUu9P/oHifrpQieScccJH0PxNhZ
Vz8Hhj6mBLNyEoxfgHnfpAP2M8KeBRE0ZTHBjakCanSzwHKmVsKXJMF/IfgHjx0Y
TT4Nw8zgyOWxsmzNq793k5AoVvsbOiYX9CdyRsmBm6MN8DZ/kiPcJNl0Iu9O2BNa
bubEZGgX0uYk0yMzilCPUbvicluoScpckafgUC8gr0MatVFZ3LUpy+O6bopPbFz8
VSsxboJNjzVwsCfAiFkNO0+SKrf1fNzFxG/GOXE+vn7eXgcl6xGn9IQsrg0h3sqJ
arZ8GV7SwY9qVIrFbyF+6UOYppJ9hj9K0Hp/ZgwskpT8byzGh8M+Rn9QB8/WZqyZ
APlIyifj7IQ3vdnF49Oz+aA9E//QN2cTWG8pg7IWRol3D5hwSnNL0060wpK3tzHo
h6J0RUrUkkzfJKCsBnsyhl+7DaHkhKGVakZOPgpljx63W0QjteOukq0l/VcPLtY8
v6/WeHOGMq/6K73o7d65VDGwXrFqmI5Cnj/SNMuTbgb+kr/46dFp5j22PwMEumd5
Ddvz/Ivi1y91ok7bKjsQQpYUPxbbpT3WN/PCo3KIfS2si/N+oOqZt62bFyYUQ9Ns
bs47JnH7ehZNKUHqERHzZ1ya9G/z4LdlXbImhXySNcVZGmaWkppKiTbTojplWiea
+0lVDMl/BUYjqu3PEyXbm4tc8Q+ZoOTBK+R8Xok7Tkq4GXvgKq83e7NGTF59DZei
jXrh1rfmLyAi7r3rQdtzxXQtcz169F6xz3jwDIW7g9etE5VwCmmIoHHsr6wSFSTU
6ZucEC3Dktm3ns3DLJlOkS42xeCfBlGDJE0GLCjEksrWQ3Gr4SjUzVfU5CDIVaOo
UrRidks7Dy2GvArr7Km1EzN4PdHNvDqeAIiMKUydwSHEdw+QesuLFJW6bp3q22Z1
yAN+7hYpVBNc/85/bfKqHN55GWne1+s4DabF0PY8hJVHqltu3W6TTOJKRUtXIQD/
g5xBrZrG4J2TWoJPsv+Ptoo6sXqN2jAFdH2C6sgZkIaHDnTKNU0brTgCG5DvUCFh
jQpzVf+YITK7WpkTQZ1HUwmp9Co9rhnC0dzG9UBeCgHtlRaWeWxhYJBTEXtQz5GS
YTc2+or5TR0CNexjn+047Q2NIKzEmRcxy6ZxPMjXM9OhZgCKvPVtLawb//9p7RFI
KszO+tnifEVD6DH9/Xr+8NNBsAPi+1Q0YzNZINX3Aa1mE+xC22OkkCD6mo84JpWK
4X5iB808/j2z2DShJIBeTSb5d8dPqgwgPddhH0LMy/j28rqyOf82egM3LjmLubyD
oPGYZxdIqHN7lTiO0SVpvMIKiSaaWB6dk1/LYkz/M1H4YUVyZIG6PirsfJAnHAgN
uozdkz007awLYkRHaphbuyF/IcKxU3FWSyaBoTRfOYcz5h+ejCZdISFiuEtxDUmg
SBUZZWqL7pL+HDO0Efc1XWMPxWmBRBV5u6HlAH+fCtpAP5OjAamvSUbyJJoFy/Jx
is5tr/Ca5CuxKO0GOFPCNtKr1PywilTgjVs2sE0rAJgZwzLiK0QG7KkDwvJEudJT
B9bw4kw7CaGWZTylumqjr1PL19M0tV1ufQt4416VUKx9BYjyEBPgc8QY9sbjQsD7
XlEi7AMiV8IfpvYpLTSATkGEc/w1AXHQtNiDK9+vzsCd8vetEaZOX6PcN2fh7R0U
2LUF0Ys1OhqdPLYKIgzxzog5HZHzaG2NzlDXnH8BVmYtYhdBukjDa9a4ZCV15sgw
ICN440FpDJC275pi7+LjLlFxp/7kJEE0kv0Z9+D0GusXkK9EpnZNhZpYv8PB/Zq4
LUpZbwmAvGZwO4TuC5PirFVTO7nOyJU94QdLf1f3ausfPrsv+jb6vD7pDQxdA2Nm
TQI30mFwO/ktq4AA0TakPP9Ttp3z6FiPWBJGHDqA5fenjHXRwWXJ3wt0KKqqvjpn
4w8klq4ZtsNlfeWeMW/x75b58H6xR3EYBMxVCSHXnieGcuedzgEx/KFhJXVlioGa
BxN0yjyH+tLHzMmo4LHHLiw4Clrw6KiokttK1upWvDCQ5IiDDeW1NZ3RhhYTQSM4
Xfp1ED3fcXKgsjYugj/J9+DTYkSSFGzNwKvloAQceH0juGs42T2Vl9gyf30WHDDo
cgz8t1rnSYoyXrGvu5zlh7DllOB4dPulTWJD3iqkC8skjVkRD4n/dUOo6D5S3nP6
ABQ64H6lQRKWsKueAlJJvInfzaCu4vSag6sAlWUH4dSmNcVraUstI9AtIDIgeVjc
XeaHfi+uzKxopRCrBW4h/rwedsKLem/plLwfWD1NoVYHBBM6HXW2eB28h7I49a3G
lLw+KfjpVIc3KQ2ADdzFfzwBXjq4gL8MieKs7JOknxAEMAsNpV3YwiVBN5d7enGB
YEa+N9VCbtWYfAzoVjHKVUHtjL6hsrbc7bZBLUPwLJ0yprrv0ld6i5Nacvf/xAa4
K+sgwrQZNLO4WcI45FGliKSn0Nf8Ay9R5RiCYYKcUztMO9TpfBg1JbHF9MqiCKRQ
rZKaED7ZxHQ0zN16pIlYEz6Ci6sqkez5nK0MQUfecI34WQG4dOvukCFG482oC7Zg
3+usxCFRzY95YDasQC931LXk876IfBsJjwtQ6HqNXpc6iV2EgjIKYP0yGDmBTDH7
lJGr/wa3XJXClYL2EDa81NopvQ91xEWticgCuhuvnejqsUyD0DngaWzde2E4fpvd
teo5vHW/kiJ72NZWLPGV+xkuABjykmhjvtxZ7b0rDFkdqKeS/TgPmhkfU261+3ve
9CmRimWqVHNZAvoC1MqlnPIKzXG8Etkupoh4u95ofxGIBDw3/bs3aa+J0p5EXoru
d5p8NF5RAQXBDNLnr+l4y29ij39ymrgessjsrCpmj0JLd4ATnpq0C/smi0I7mnLa
+u69Q9He4axUAZyDlT65+ljQNRpctEYUDv+u3jEXfJ7BOdSuWFmHN2/PRUnjlsMW
3o/AEjULmoRSpcc5UmGdyLc3M2AjRf7KijxWxpoLb19VhQIma9fJ685u+RM8YUj3
0wuW9634OBRQpdmWVzKoMBirjdjS3KmIzFkbu6t81F7CZ+6MHmIKjgPuVboRyVtS
GFGJ6xT3Sk3qIwFcE8G3C9WOsJfuNZWhiGFJnVaTS7bQYqJWfhDxVp4EM3vEqQBz
1Jrw1988HJKFXavfMBpVsmv7S4fX1ixkz259rkKznVaTgd6vns9JvEo8B0MM1WYY
4TYWR5qJFSD1d14gQga74G1O5Ujy2+OZyNt4vfAFpxH7jeVqH4qaJHDlFtVLA0Bh
MEAJgfA/DD5bLOfANNCk2d89uhK3p0gJSr73om/yIE6+SS6F4TDnLM+dLFXRUxU9
bS24vZ3gKtJ9yvRjw8EDPy4ODmWKWS7laClY+Sb/71K0Hoakq1nWqrbjhYgnVPt5
VT2Ln5zquApSKxmOlGRkBeUmB++84hFzfw2IJDk9RTvZgFBSzXbI66fXhhgndxrl
grPHG53gcFIAl5of7wheS0LkfTwN1uA0rNw5e8smcVj4aKXkQHLYe7tITApKiJP6
6YX+XJFNAJuNgH9H/VbSdKAiOM+JyuuVhlN+V9d+MAg38P3wq5B2VUx1WS21Xper
YUcHON8Onbqq4dHAmndbZ4YVdyBdNm8BVppuhdhOSkAGmC7yfaLkcCLqQCv7xqrP
3vHcXnxrscpUrtVpX1Bjk+5PQS2QPRpUzH5V7aLstjtvgOTkNfy21MOCawfTS0HC
Yn2oGxpJ5f+5SdpZqzHXFssDpNx2qtBfnehbwE445esEB63OBKNqwBbls9i+5jJU
GLiKfbQDZg4oaueWzPFZXuUIqtj1JMcQ333JpChQgBNT3pCKqqjPn18AQrm1gyBF
WxR9RmtxlQGRSgzSSjn1SM5WQs+1QOo8pWaa2V0s7mL5txvsi0DtHUyngLDq4b66
z2DILkMP45/NxcGcIdg5Wy7kH7RA3WJLG/k5LXuQDJE/cHhVTnN7E/IyneCeibXf
dnJNfbGxs78APN1P6OZWEQypw3iG7IFLgHXV3Fa29laksPrRj+oDoR3bJ7zxU74A
g1NbDTCJ5Ili2gLcKNzMF4FB2Sw/o+jOJK7ApK/tYvGiEYb67YZBOLffJZx3XehO
xVOYzeg/25epZrK5g1za1E6zovW03mlT4or6VY9yMiaVzRjOAqav91q0j9tIDxL2
M0pDJBz9Qkv0AS0Y5Fn7/jqPbY6HBijTUNLRaMmY9ZG86KZuvHduMsbitAFrRFI0
4iw/25pk2AvOdYf2YRgv/cuYqoud/p8n27L44Fm5FqTKj4bu7P/V39W1+JqiOEND
a46phdzZCpbw3SzMBwRtTuZXw/KKFcDSDHAen6ppqaWKQXqWFyBamavjUpip2iPV
YvLI7aV3EKgk6Rt6h30PXCkktPJ1Dgjh+bhmQAbt6jNwltfl/DuJwr8YW4jZjyc5
v3yErXicdXU9oGfpzHCYcvbFQLE4gjI6c+cfhFb7s1EHi4aXKgqC9mATXM1iF/r5
7r+tWJwg8KQTPDmFQKfd8lL5Sn45DpKjyzXRoGf/TewDxljGkfLoy/trhs7hgGd9
KrSzT53tEeX/0x7BzhwKic5WJ9+k15GjAfMX8ZaqHZSaQn8u32BXpl/RWwQmw0km
F5l/Sxht2N3ma8C3/RtsaNDnzxZ0NqFJ2fHgy1N+n28tzTFgP2wL38q+5/83VXQw
/me4kWwmw/Ra9UN7yZGU+i59M3auDqCi44ee+zCCQP7y4rS1fm5tI5BJFZNaQb9r
QoNB6DYE53oGQXyL05bVcmDWnGaGbl074zsUsn4eqDWt9CRKPNC6Vl1i4E6lniyI
W7+s7PjKEcgx41xGn0PvxPx9629Wzsue0CcToAr3sfjmtUxBqy39AD8rhKZKPXGf
lZ9KCrxLO3zAfJoSTzdxfozFMYWWR/DzOcQn2H2ajSX1iQivx5XXgbt9R4Z1NCPy
G+AHl69+hKmS7/g7VVSm3GvnB/d8EIbHobBEOqWq+EE3HbLk07orX3hpQ/hJnPZj
48sDCYzvPg3UKh4INx5E8clg0+ZYTnJ1ZqS0bYrFvdqCeL3VYENZMvjB5hgOHnJQ
JiY6vMQkjDGdS5rJUX89rzNIWjBt3HlxRGKTd3OZvaTfVb+hX/0g6/R8gEzTch0B
yg1w4OL2suo/MOL7mqaOK54AgtdHfAlHOGoY7DEep19OcW/WhaO4YgCqK21+C2mv
fdzgbVZfx+iKp3jXM/fzzp08F5yspOZi6y6mwA3dYvXOc59JUc4bNImq1O3sNJjH
UTkcT71CV2zJrTSB7t0EozGcR7/NlwSmh2MKTGZ8EN+wEG8wI358AfbPCyehpA4Y
gi5oVhREbOEYefcKqjtHpDMVA5pLXtiTYvQvRk7nymd/HyAhMNF3KwgbeYYkiIX3
ZSlaBc6Dd1LnXCGcbAT6OH3ISF4WqNvbYoUhr0xeP9iFLYTZR0QMcE88UWNeNxOB
8BMMK15xeS8x6JrQM0ILj5thSmFbN2ky31iwAlFOS4VanMHoE95wId4lmWcN2sL1
noYVWdvunDlChrJoByCLOqyqMJTSBejM+4cqS8w+HK26F66ikWzw0Rjcv2xaRwW0
3mrs3/Y8VNgxq1ndcSwkWAq+KSf0AdZXm1Zu0jE5xs24JnZ+hJNTyW/g6WeR2pXb
wK9Ld2wxeq9xpvX9bZTP34aJUFgms29v5I1GFKYOG2nONqp3p9U92vEWyPFVFfjR
5IqJ6iW0+x7NCSsX5Zc8i+K7JEMUJYCxrlaYK/LQfYkqqsg7tyZpHog/rR9HH09I
MADEZDr3HmiDDKh19JbBdcBr7ofcSyO3ZgyOqF41oDXjisflIqCkXaYjjyZ/bVtX
i/BtYnApKMa6dsypiHv0lZuBYqAIjlCgHUvevFoPavhvtI1RlqE9OFHOBpjXcEGE
yOOT7NtAdM8Zj74YZmuNA6RcabqSZ/j7anhOL7mThl9dQkVlgBOIDxO//xIikq+/
WbXd+qrB2liu+d2l5SViOQtpy/tck9xTnb5q2bLiYx29mZv9PRg29HNezYytyv+E
c3cZz0jkjspU954lKl6rM3mh5w/7TyhRalY8cM1NGhB0OroXwXkQZh+V7LQCUD56
9KWb3tphD2Fi0dJ+PJIizz7+mU22hRQ8O69jl5Qx+FIdRBtyMx9nwMGSKixlhlJN
Ty9wkCF2nGqvW+2HcWv+kZ0eACkCpga2EEkoD7mpXVy48xYV7VxpJ1QLh+A2VViW
E8UoVoGB6lJ7EiEWJV6/Q6ACzsOGuFaBfq4lLCYdXQv2N/U5x+0zlagDl1V6nopS
tsAl2LqOc3uevwnLeWk3PiYeL9/t+5yq5qskRAz7aC42ZgXvMT0YX0gW0f3ej4yf
a09ZPKmVWSeF7awgFYoueNmwGkI/N6tmdkExSQF5S/gSJxEuBZAu2wo6wZHoIL1A
p/keEu5iVb9zCo+uTxbw+8Sh/8LSikhfPendJoTA62gHPHq4A+OotOVVScXEDq29
WZhdojythda+Eng3JR3mzUAF0ZM+w9e1v+dCKPcUEhNshQnuLHJTHpY2WQxEi8ai
bdlxwKCJ5c/0QXhWJNLUOW+mfuRcV6OEvypnaztp0emVMqwkm/v4H9dtrTBUgQrq
V5hkJ/QWxCLVmazpRvcu8YxQT6GbE+eth15UijzlU+spu8/7gy/ETFegQ7wQO9qY
aHDBWUVzKBCR8yNFjrckGzT5RjW62XIWZYtdApk73G2E8OP3kozFHdTj8AtFkI/Q
OU2eWLMl3gZnoqS1cZUKU9ThBY0/22OXw6me5CSjvT9Tj7F4cWi7IrwjZM0uw5oq
3lmLo2w6GeeE5+dI3/DcrkIr9Vf0w9JtY64v6xVBCQ8FBY39mGKSZFbrvigRQQgJ
ZaNDNo9w5NyigHwsqazAAlu5nGmQXcMGQyO8ISTQ643RAaMyZ0dl+2HqLjmrTzar
+xGSduMzC6ah/3AeBU98TPAp3tlWr+r+Hj3j1abZ58WHEu5yUeRIjg64FVFzNIT3
kM6FaiSPc87X8dc4vEEcU63SBTDtcv/gom0Ku5HoGMreKJ9YutkhWE1uZ/bMFxgh
UPcWj90mqYsO+6nUTDmGtKwBBlz+ZEpyu68av5EaWvekdYxnXVmZJ6OLlQ1cErfM
8uhlF3r0B8inChFmkyx8asFBk3WImpLdcL2nD5SBzRGLx2Wkst6JPmx6QPofTaxC
DNqe9845aB564oLi8QFWATK9zv5kozgjpBrb/COcYCN3OjLILq25HMHncFPzpMh+
cI+kRah+EpARtyp5MaWrZiKOESrz8ZTkNqoaIlbKv8A5h6tBTZnffkeZdA1qGgPr
mRDnc9EinhrQJdWX5hg1sm3XVpGcB/nYq+cT3IVQYQrifNBQNhkzQ/ZXlM2BFSbT
aaVxSKKp4xNwfQ6qv4X2I8gcMII6/yk3Wvr0b6W6J01sRGWcZpn5csTt6SycNW3g
Vcl1IHbrz8NEV5kZ8femu6Tqm3YBrT+Fs956OgccCDNVWWjA4rk9RQ4N5SDiL7Ur
xwazEFohi6+yaTH4l/cBoeJ06Z30P/MDZrH0N7A30JnmypEFmWdZLLlTX0p4WPg6
UJk/Wopujp5lFat7ba54qX+BEnUN+0LjNLUeDYzsayHW+wd3HOOWNepy890KvEkn
FZWOXjEpXRBk9qrdWm5ESK/r6DrSzMctBO00M6hjATkvs5JeTtZ8WC2Ox8Ud6Vw9
mh0HH5MH4DA5Kg+zlBaOFfhGKJ0IzQPzxoOORUjSrtv/XTZPi748K5C9k7sHTPhl
9fjznZIFTDps5aToWU+rxaOxXk3zP4JjZPAu3W6B5wl9oaX+BdXUqbcDOlsLfQd5
nkAzmbEBb1NdeV4otRCv5Pr9kxJxb8VSTPGJLlsbRVwZ3kzQsbci1ym1P+2lIrEh
hAE3YQIXB/HgkFuqn+kIDO+3lhnuWcD5IowEZyFoQSoVzUD0++xlYoV9RMw6JkTu
vGjhP05wX7hJNdryj/0QMY2MuzCIeN/4yecFlpVWcvOMemitWb9hI5Z7M0FmlmXt
vfzlFSoKhHwUObZSocKqsNlR2Kj+S9LX8fQFus7jiMxe7aGksIck+AMOBmMcOvFk
axyPBBkYy7o2r+YWhsSCovlLXGiKKIaKJuQY/WjcT4KYVRTrTnMywDYjLoH5ETsj
/T8kFy85v2MurNdhdnrRU5C7/kZ3gOUQD3e1Cu14N2zG14HVnugEkboc7q4kPqIA
HW/0P7pR3K8Y9qH5biL0jWpcKL9zWTkiPb37ekTgw5PalAlGVhGD7F7heOxXP/vW
2U/LqmLsLZgsN29ct6EttY5GsD25+WqCQij2kLVe9jwxZjS/s5gilS7HO4ivW6mI
8xYmbossekhOQH4YauBp9Z5wN22dHQ78lFDy3jqn0l5UFku38exnX2rieUd6Uydg
jRoMEJMl1fid4vCOyWCoKkfZjDUVEEKTE36y0oG7EjEdJH2wpONrP+i74kBB5ese
m3qevbMeasGK2IPibPxsP96g0UBn705kvNRW0vgLSBjEfr2hfaC7yieXw3PEZqBr
PIUGqK5HECO/CRP9sSQjY8lMwuMPKGSECvn3JI65Erw7bcY+InZUdnj+Tlp+21p5
jTvSutit/MAO0iG1ePuNobhs0QzGNBzrGdYtmMAr63y5l7gSAgbYu+onjysaKs2Y
LmOVKz7UvNXcJJ5vH0cS4jjboip/MS5u9YAt8J0E3Q4BPrk1H1htncE4ZalConLA
l0LHDxIzKctxcq05ysN3x6vauoBdxmkmFJ9sgtLH25qvb7oF/Wt7SEhSy2UAvD7B
oKWJtZb8olQkDMbuUmj8eGiYqC/snQkJ08AI6APTJE65guomlGIZbUb78/B4M4iX
2kTu6KesqJjhOyhJ6f/bt4QHjVkpCfFb7n3SQEXAqy4GR/r11DNegyrAH4CvAEs4
hyUmXrmN+E+JvC2sGXlX8gs68RLPfzuGFyXc2M+T1RXcu0+Y96PLDoh5y4fTIZjz
LO+OrvmdhlYweK1o/Ym4Yql94JL9rZPKTR2ubALZbkytjYxGeht+eQLeFNyb0joX
fGol9crQsSNbhjMlCKFc4IA4QKHauM0vaXCvM3+46H0j6pg6cnQ4hT/aFssYE/x1
UukCLaPFYIvEcXPuyAkJtXn9l26NKXSac1BkXlykm19JMiyxNh/kJ91aldgMAkv2
/qj4yBeNx0Ne8iYE5Fy2r+pWLOxFiAgk9bur4z4qILCPgbyRyXfgnipiIAH4I0+S
WSRNTmkiRtWIm0X+DGctzUHiAeGW0wHAmFyKpASWDic52xkB+7Dfrt7ReCcvaV9C
gxamX3zdK3PVe13wPvIZBkcpMOcDxm/S9j6P9ial5SGzo2RXikDOQMMSvYY1Tj0C
pm2isdMWgfhp1fWiB/0NRUMsp5FOSptx/MhadjBK7+k0K/PSCvafgrpSl9d/vEyH
4txgDtemKsYd5T5rtvRyeD+RbG8ihbgYm7JYkNed8H2sGRn7K/KNYQu0IM2NKqjt
QUEYPwdhQKILqYQtNUcFr0+nX369A8VQjAB2VQQSC0UyGEeEfwxuTGEPoIxJKp2K
2f8mH5FXi+I0S6se8QakYHyH+Rshx9T2b75eevdgOqI5MPfsNhEj/sx5aYXGtTCm
TWTqOkAFqPlDPR64wxjBWNdes9AxnTv0eB4Eu4lsgiosJkQyK5WDbjXOtbbuwup9
drTzahV3tQfUfR4D8NVuMoKmzFTcxjbvRgpUhli4s52YxRgt85XEvhS4nsiklmL9
KRLdoAlrTv+RMOyFyqBlSiwcNSx9KyM2P5ZeTbKqwCAo62S4+ZerBk/syYHsnSDW
mkcxK3sBVOdmJerywzTEGnIlWBjFdGE4tNO2yDLEdlgL2seqeELiEmEpcXn1JLR7
CPF0tqUve280AbxfckEgC0gPal59+a+ajaKEoZAyLwP/NPNfCd9xW2rkXmM+anJk
fUzd6I/t8PDVMIB3HDcuUdCAPQ9zAG9a+cLi7CssLPl06kVYnzyUYxOAB9FbZ1Yx
bxH4+4cvOKVqhVqLnsXGDUtyxXymD8jldl+jJDXVlPQshXDOvmEQLwxx/QCAFIYG
PeQF6w2XSkUW9QEtBS045GOy9cobLtWRybiUXBVvDQU/fwd1uYCW4c4lLFuy5vX+
jQRZpR4XKXenvMwPu6ILvTztr611PEJmLsRCVcehqC2YbAEbktQyU+7TzMs8+sHj
MAG9dMgbfbCLJdPR09JuS6tTsRbRbqEahE06fqRS949DJIPFZkGnvrkEWpxeTzCC
PmeJvBtWY5pR5RcH7WZSS4Zi8uI1WHfrxcBisDTKfy1qcmAKAjAyTP5jNYFSfTU7
+aj8Jc9lLUoqE5gC+1JFqTdP0uvWHoHj8I9lXgchtKC5O2Pz2dy4/eXaIc2S5CrQ
zjvWGjnWkU7tuvq7KGGYoHlNyJg/IbXwRKOQge3XOYKvjUqKIVpd2npY7Up3iDTU
NSbhibEVZ06z6Bktu53ii+NrNkkdDIBWbYPuYL+0P+Gfg8+umYZZWXhZybQ6+9Xh
J81q7QtBfv+nfjBiCaNxK/G50mM88jQEZLZamWKy0WGV1CKomRnq5rw+JKuwG8v5
KaYe42HlFJ5Y5/4ugpyCvR/ewfq79RG3SPPvoMO2jyxT9FaJcdjLbRz8lz5RdE76
NLdFGjPyLgSb7DxE2bF7vluXGctu8h33hf2PvZ3R5udW3SF+9UdshutoxGf/DbLg
gW6jSRUXXKpYpBZp7Koy149UETZ5lg1JHjjSjPy6SuG0pBelPaUX7jBOff9zYRuJ
aeHlBZb1j90M5olS4hZGVcM2GdO/XdkdlSzcXgOJYsL0eu+nCIm18xdS7GVjML6t
uA9yzdUSTQe9l2g5CkzQJPD7kVYtru708ekJqn5j21NGWbroRDnLpco5Xjrk+o4G
ZLWOohzSVSDtGQvIWlytjqGXjAscPaclAm1+MGnGgeeQhFIRGBpfmfZqrWu+Xjpu
BXVS0n9Y4ofHba9YyUobPFnEMDg2pfErBYOQ64xYgtcmFaba05tiXnYP/m9BxC/k
OWOPbKYKiTuScl8T3CftDnPkBwy4/zK6XB3zGyh516TgWhTUwIT8FVThzN2u2hDT
dKcoxI8hJY+hZgO22y8kD+1clBTDm38w0IBw+JL9vkJMrtia5rOcEYrjZRQdkcML
paRdsCJhcVtB8rPHA5biggU7rQLpeLxHzomnOhzBfVx17Af9gE1wB8oWldWLP7X+
0LadsimdxpAez3i7Atv5b46uoYXWZxrXFkmtYnYCwjFaaRBlshq7esevfQR2z3Ff
wIi9uDyf2bJNRNzn0JWQrQ9kVWrzpQEzAdRKumdjuupQOPiTkzw8kiebeg9Q/zmX
0cNyqUWjIrp5sJEwEe+8UrsohTvLIH/0xI20vaYO7uEa/W6GRX/ZITuuPsl5Mow3
GXRjmJSZrIhN6qA1/FZBZnpGsq+8RKFTrtnCELWz/VAvYNQFj092IDXAaTJSuEOK
gE7pFAPuSzij6AOt4Ni0BtQSvsAw8bbeh94zTqwnQMQIYWvPqBzxr0SY45Skt/f2
F0QgcQ8vdUL/upC9YJzG5xLDDNF9HOQjeP3JXJOr3+d44mSEmUSZ2phwZtqz8v7C
j8EOLykRPbXqHi9xDfohiLmm8TqBc1vvWuXGlZ9k1SMJrzTwP558PgIaQPgaEFMC
SdZ+purW48OSO/6ckao/+cC68h4DpwMtW02+tbz0tMpW28M9DXBXEEQDjtjztrIo
X3NvLB/DuxV+P2tx6hsFT1R8bT7nMgArUAz17vU3R/lNg92AUmOItC7fxr5RFS+F
3BM1reGzfLyo8Z93LKyPQG0NHd+Qedjoyz2agZtg8V2QS2mH/fHdONjqqL3wp/OR
VuN2zYe36cm4jXYQeVv3i9bXlf+CzLQ7W29ireoXdSd6dzI5bC98RcgB9KzjdOdZ
oRNQ4YeIFPh+LuzFR8edoXaDUS3BQhwCikz2O3+HyyH+CQFbEcs9OoDA+2ToLthw
W+c6h3VwbN177VNinpiPOb8jnuERsxdkt2/oZnQESXrMGInoad9VEJ8SOdN1B/gX
lopxyHpiUyAMIo15I2P4Yg/q/BJF4onHf+0p/gH38ha3PMHSrqOVNLDY0K2JFwZR
L+AXXUhc9ZIMx6YBTQit9R/xdqYps3ChcvwkykpE6SrkmeR63rG8qiGhZQQWLWBp
FWU/OwexvVBCzMw6RX+nuw5qVJhbGipYo0jL4hvawByOk904heOrYwh5t5kZdSuO
DSYZTxTTQWRbD88iwWqZPO90Qe1WmwrHezg9PmPTfCL2VtebCv679DOtYi7JIDF6
qygR7VKXwvlhKOe6EuVkryQc3xlU4mPhACB9VEeo1iK/AwGWPxapl22VM2H0pYrk
veUOCLlzj8WKhHmwcMs9NhOkbwEPTtKzVtFQ5lGHl1lpghYravWSDSzxlF9o//cB
GDWPi8xumbrdktbIbaCkAIGcXwWRmfAnyrbvbqUJzecgsxhPTOr5bfftyBILe9kt
PcDgcKfz1j03ndCkJ3RNK4i4uK9L/S0LT4cXuO94FxVgc3tVV2bqq0Ty+iOmNe81
BfZnWEe1qR6CJ9AyG+726RJd7lM31koq01gKHLPnsamYmyTB2mmvz2awgJ6ML5Io
Vtjzx05pVFUDak+WYG0IcmY9gYaIpw7n2Y8dUjhUUjwR9oJavY1pKRC8RjS2IeB/
BmvT6nYlhiMTeasJ5bXjJ3yb1YGwG+WzGcJYDHLkYLGkY46r8uyp8mBxSmwxg7l0
aYX4apLf0zluehZK9FurTdPuBKt7XvbcK3t5bbR7gfM41BnmKGMGhs58GGpzjrFT
IEgFyOqooMA3VaJhDp1JHStNs+5Rzxbcyn7jI8WOYM6S9wTPdtdbX5W+3xCs4UP5
FMEU98dN1KsmcjGivmQcUJzFzc1QqHMz8+FQIaGPdlSif42+B+31WyUXsQW2BqRY
lIudCVJ8mnxerLOUT00Jj4R7sPSbFalPig8JBfSyIc5FIENJUIORPafFiFkZCQKc
z8OI7pkGDnmIbp+uCs1S/vMVwXs2/CEp700MzJgGkMdCNjiUJWUAzeqo4X/Smcbx
y6tqPMY8vRd7T/RLsCqVpP8IEpnPr/fTZa0sL1QC65+ipPUsSZyjKM9LQZx6Rxij
xKUetUMZOBQmSxnBB6shixeFD52LBXfkGJbE6AkBpgDDszGNwjnidiWznyziB4Us
fTJbQXbm1VWqavHbqPMoLenYCIZ0BVlQyUJ8EbF3XtuSG/AOopMe+lTe61NoC8m0
I3CzVmErz0BgbcQNAeHYUYUAaARqUjnQCPOoP15rbdovkoqGUF04I9saF7G/FwY/
68idMkIwHnq6papqp0veSbYvEtgm4KjvLTxcXH/WtcHUD4o6ccVHLg9p0+W5ke2d
2VZUcIqNsQfuuApKWtFVC/MJAzwmhUeXMuE9rogeaBuwEA4t/40uq9rwbY1p+QnL
fss4fNMlCH23Z1EWwofklg5nAmDZAHD9PjuLVelFvVt1G7AJqJroeHN+dI34CJ1P
20jiQqER6UL0b0XMZsqxnIBdi7aoLaOTOP85Ye+FBKUyFL3EhSe+o3p5Ec3GUs0O
oaptbOpqxGBV6OyueTA7XyetiI/4RrhMGUP5wQbrLCO5uAOq/LyT2K4JvYqQMLml
AKXzLa/N+YAOarqgqw4kiBRt2r0LvzFSwdx4rzQxv7BqH8bQ3IEsx97wHE5IlAOr
tmq4v4GvWM8ITwwBJB7WaQZL/3Bwf9+BejpZfuKTrVRWaLAWgEWh5i2wMQBZq2cu
m1i5t9JDifLHYDr5u0plYg2lfw2F31Ub1eKcM0A/urLyrOZt03NZAnpnjHzI7LsS
2O2VfHyhMmlloAeiebq5h9X+azIWWMW5BZ5Yl51maKNa/Id/z8BTXE8KHba3Mub0
vY5c+T7GBFo21DpMvH4q2vvxT6refb7Btn4jVIO9+ictVUH/qbh4Mqc070HZN7TC
GkApZgqFNk2LUTUQsSkbyzfrVNwxWEC57oWfQ7pWTXCb7e8eQ9ETkMU00GOwgNrj
tFGdnEsbBRgVxuaUusK7zqJcopm7NZN8u14V+oF942IR+Scbyimpg0y1530WzxlM
BbVwaA6EDyPAUC8fjyBvPQC0J44RjhPtwkXtoj4yU4RDCzRIpGOVqax1bbtcikHg
Zm2a5vv9XhPbRNluHHYL4UeUOe87vtzWCJ1IVkmtIwLKv3GbSC1RGNd/BIP1p2Wi
vlIDlQ0UX3YFmWqRtS7vuyMQ8zWzrMQfYMQqsD4vTmj8jIR6unQSy9xEsKmhnH21
ZeWTa20NJ5JLVYIhy2dsLOHWdRdAK0/u6LvGRmCsP/X84Cx4bE17NzyDweOesJ9b
7HsSN1fEYplTea8QP530igKM/OnBadTpZyWOIqApiHixK/lMC0Xrw2cXQOHzzqYv
OyzJk0LDizVcDJDsDbzI1b1pozA1/s80wAs+jxDWl07Tf7sLm/NbQP4XGdR0b+bT
U/bWJHzCzCfL9HBgHUs3DeCoGQNZvpGhNWq4z+s/zyCcUZCxuQkaABI16TiXywcz
+lyrzLWL2eX89MfqhAp9eoaL1nqou/K5N2J+Znv8hxeN8eMSCMbBAjttunlwCuoL
rOUXs07hsMiGTiE79jeX7qaeE1wnFgbANSKSgcVc3f5Yc4e8BjDOZBVQmbmfdKP4
WnF/yExz0Opd60eKxfhXVAP/+4g++fBwrKq9oL1+4GdQbrRH6aZNU4kjaThGiDKm
Hkamk3tK0KurlXT68Zy6A8IT7HkaKDy9eBbrbQDzYRmLCoq6huJ87twhLViptW+g
YtTEWqVw8CVKk3+IaKW8GBZXRIBTW3q623/gaL02ddigSughGI/jFskdzPI9UUBJ
eBYfovEvEzmiwQgQXtvhgl4dJ9qgAaHOLgExa43c2x1c8vkmRbYBBTza6d+sfff6
hLqgQoYVm+3hL3oBli7Xsv0SlOhXJ3zFwmwDgJYXgEGwzF8VoLjvkpKGNNcAEYpg
IVFqH+NTJYnumwCj3YGcdoxJMs/YtBvaO7pO7H/ts4zkNHOMd8DgefKUaKNorgKF
Gpy+SclyOWqkgFmnra5duXE4E3/GevglaNzgYRkxFHx3r4QcXcGlndUoReTpUVsh
g2HBo8pb/70xaZPRYBq+EP7RBq8FTlrOTV3SQsN5SVDGuI1JQEKpWdKCN3yGHORW
aV2gdDTzAiTj9mTvUBsQg74s1gbHUCYrk5RyGWedxctKP3HIvp61iVaUUbP8Q2MC
PH2Rpy0u4qMMgxu2e4jFH4dvRzBrR3ESnMCY7++fqcXgkUOw/iI8TgB4YAF9IAkO
2m8BrmcMuhdbg0X5WYpWQxFcr35UhYbm4xgc9fFttj/xKv/d+lXXhfsFwlGmkT0f
5dv1R20eHCATC8BX1L3MJXqr55TjaiUviNVbXcAGu2K8tyba4ywP3RIBEMs5HApK
Zjs9kc/oEd8ws/kygbGxAjXjDN1JnieocHApeaDKba/PrBzfL+64CTSv2sFJMWFC
se84JsBQ3ZlLDlwJcUjK8nDRLIKgB0PEO3Uo4pyl1uHWeeVQDhkhAFqMw2TtZBs6
+NGAyYloUZKV10csYOTiePX/fTq+VrktJVahnfe4tNvsYD0wXNTy42//fNcvP/zW
mP+YmzCMycUj+jXXb05hr+bVnuM21/jJwv1in1vCv+QSQ7JqZIEfZybJoHSd9LAy
u2dgr93Y4qv14YB6CQhvcTG6ZmZr/edgPGJC3c3vXSlPyjEUpuOjsL5tAP5ePVJp
4RLwxI89ql9wtQsE5bIX+A2FRIw7d0xOdCaotzLOznKzS0bBTK+RdMQ9BspdffHG
vmT5MUTq6GE+RjKPGEuIFx4ZhHm8F3iWahSJ+qfxHvrtEVMxirhVwLLbsUzAN1fQ
IYCH3JCJQgak6PJTCCnUxDzfPp3SdHMMJMSJLp0jdRRbYWl7vfS739E3jTjzqhfw
yGYoOMgO6tPCaxZwa5np2dKQxL3NqzaEJ1TzFRT4AefatniB96/y90RglvwQHI+8
+ASB180JYi7vNBdDShhyFZ1zOIRH9jI4vxqPkkkgV/YYG7Sm28sfAsZSo0mZhfnS
/MHDAqU0zusX96QoayKjAKZmEwYtB9XnT/tzgpRzsUt+WRfre0BjXISb6vpDz58n
vCGoNawb0a2MxgEjJVRw5Idi5KmzU2w1UEGuvwfksXfoVFEGBgK+ep53xaCiHjnP
a/FAOzVXD4Hl2duPxLGU1lYHK447DoKxE6SMfLWP2XVDY5Xf/I6jxMYRLN1pzDil
44yyUYSZkpDo6wibsLaiN40W3lqNlDiHZPMxcKCb70j4yZpZsXaU0n6B9SuMtulg
rx7s9JCSnuKCg86VYqn9OwpDFQ06dmSnfiYFUplCmCsU8Iw0wQ43kl3TMpg7bzhx
jjdSOHxvMEt1CC8zXCZB/IeyUNnizKqAWY1YTBuoPwYEAu1wsRxsrDMg3PwgPIWW
HDj+/SyLmhz5zFajgzmwgD9xt6BFSmAg/t5yR2jsFpcNnln+fiidE5IrFM8Aw6DR
pNhIIZzs+2DaRcHINZZNmpqZhfXzjgyqor5f/mtuEU3/9+1o9oIjL47dpobGo1tQ
5oB/Q0ijGeyneBz7GgqUDGkW1G8/eEj6k0fEjxpVa21nfcXNb6hvAlzaiBGo5kZ6
QfLXYY7xaFhZUloMANE7mp7u/90xdov2ESINVy0c4Qb0GAlvalIiqGpzUBfQmvt5
sE1yQBjqLjWQLKKY8z5i9FlcXGonkoPXul5kfO9TatSWGPmkO6EKOTdKryLK7UYx
NxaHxtpDYvTZ09Ippl3BkTeJYI+lqV6w/VipCNA3eRRH5RrSKr5BXQCD1LflzZ0Y
vxpGo3l4gaEvPa4iiU7YEMF1QqNwccIq9nqMpvmchkdHKXllF95aG1pSQL5y0DkE
AcADbo14OUM6H8l9CptpAGCqPdPUYDiChrc8kCkNg7AhFSc4gyKdcI3aXGpYd6DW
q/FDQ2RPC5cXVJkvkRnTown7DbLUVcO4/IfF3bqAcMpXBNfeH/Ji5JMn0D2i4uwq
sLyI/ShkKo5sk8G6I9/6j518Rl+11SuU8NH6NQlab7Tjmm5oh8v4J7Os6i391Km3
S/CxyC3s6IeFphhBMqW7xQVXcRnrAkwCEdfwucT770IXq6a4/3NIMUQXTocrVIlW
K0TOek1TfWRhEiLYWpT7ryZ63JUoU1Om9WYWOUPg3xU9b/TWhgATkFbCk1hUxw/S
V5uXhRUIhhaC4KQWs/o6uB5oURrLaeuZG3HMfcSlsFhRyK9OFkU2X0mEiKA/K7i8
8rvotDKolsNmzSpenL2/ZOJWjNDNDBquk5PhaCzgRWh08ADEp+fDlYeP2wKIjfsm
b+1BSLj1qpdvj2nqJaVHjX2UEQyfJOOMHbQrrYr7K69JJwylylrweeZ28SLaDXVc
CuZInWckazPuoyu/8OismUTZGyhcxOXy268RAIvKO+0KkqttM7zbAqm4kPytyFhr
Qc7EivdrERtPFIn47ki/x7sQn704NyFbT6GH8tA+/y8Vlfeg4uOHP++rbUIBqOK3
xd+NhcRKY0QFbR1a47YT7eC/S7a2y/ayWUSUANppwg0qwShmanWTAwOOuYcNzIcA
topJbDx3ap+dhVGBcEdBHXXKU+cI3h/ZPgRiLo+pAw77xWWENzmoJuIinIk3VUCT
sTS++HKtvj06yhr93fJ8mLCNQYdHS9niAeThtiue1FjYDzwmGXvGFn9rCYTvlTdE
2UMU05ax5zIhUipMTehsXDnYg/CikDJ8xndHWiBCzNChrhGTIlerg/t0iOpn4YXi
Sw+8eVZV8DtAxBw/6RGNxSdJJb4GxUcxglED7LSpSlk/YlY9wbgOVH4bZl0IHLyV
Tk4TYXXBFS+LS8yREN94FiRMPNOuaC2LqLknpVt6EHsupnKeL6330G4B1RmC1X2r
vLf00hvHhXnH/IPB0ixAWf8wQFrZr2IuLNuloaHsh01/DFxQ4wANRdDio05RADSg
z4H+6tKsC5pvUh2xKtnA2SVILrl/+1GJGo394eiX9PNVdy6SMTL/xu0wHHEtIh+P
x5IhJlWtNddOpy4XCCHQKeWLwrlQtLBA4YXI+E4jOoEy4IP2C4glBxgFVuFBEXoG
T6sH85CKtmbt9/ywRmCPbSX1Zh3b+SJzajVJ0mffQwi5BUNmAgOvfBVqcOcRi2Pk
7hYP6Pdlsg28Id/GOxbyMIQd8kkJbZT/0bfQg24ciaJGVoonNH+O2u/o+aC89Rz8
yDC1cQ23MdE1HVtl3Zk9T96s3kUSe5BN4hrQwt1f4VAo1U+MSaMpOqPBKPsZSPT3
74DqJMrMEe2oTx+vDtWf8oB6oOgnF7PXmx+seMA5k3KS7nmnU+5twlz3cWt+vwpY
PbHAK4NpPn+5PJLGzpq9mn2h040RGvAl362hSLwpAiXs7HxPKvwgnMtCfsGx1Lyq
PRrRNfMV+wcq2WTc2oK7oj/3DJ3pgyEmfSNx7VF+CG907z3StBPikvIFvxrE2agn
drv3C5kLdIO4B48m2QNK3HwW/uXykoPOB9RRWFydtowZ7CWQltNR94H3wHxKtM+B
dBXtrcYtuYiQKoSmJc8FkWsxSH90SvoCZaxUtEO97oPOC0c7u7zzhd4xd7GVIWNn
wZ0fhd4sfEj3GyKz3tuogkO7dAROM5UKboHTZ4VXjikEhm0+W1/eudcU/o0APJRo
TN0priS9zwwTmwh250+WH7Jn7QFoZ5qTNID1vluXgmlRKQQBFe5epqKm2mHQkaii
g5ScahUZnuCwV98vBnQeWeFaHVxASGkRKAC4XL7sjDQqJUWFeAd+j2+njIHgPFXG
yr/DpVVxdvo89a3z6kLYAK2cKdt8mqfsnmT9C1sAodclpRLKGZyx7Ienm/uDGuTx
tFJMkf8oDrQffAdd7EeI0msYosSNZlygIw4sSEZSayRz17tCbNKbg+h/vJodhcCC
welHlBN9mxhwMpAWmdr3YCsvTzo4OGHnVUXJGIANPgwN1xlEz2VjAuuPnwEyCo8c
gK9FIdKCMmeKAPtFtZjV3FzQGL+M69SEj9Oh37NrBngaL1pY0G/AytKIC8TlwIDN
onQYU6MbWie6UDlPd1FTB7PbD8HIYVQCScyqPU3ASCeB53k+fU2qoaKpN6lWu6sm
rIhBbXWDa3aIRKz0ysMq3RmfoWT1pzgK9GYBB/7PvJbMqs228aqaj8iXM4e68RJS
r953ApGtBW/AjZ9shUnqGFcl2aTLH4Hq7vjVmPVBOaL+4IK65y8Tf+jvD8pRyKg9
R2TzVbU832QmjH0/TIvNsG8rrQFKgMv4TXeGkCB+K3Rq3olFDZn5fmqr5WFVMSVP
I0VqpZQCkuEbLXAGFVBXUB+SiZROVEFs5rxNOc5JFwy4VsoJ7iDMyOEz6kOgB3Dp
BTMrps6EGK5ihey7ptSxIlFX2lnp1BxcESuvgci72svSPQi3emjw467qsQwuN86e
2wfgqX92OJG9fCgGfl4SQmhd9/ez+JPuvyobZloxNrruoIbB8D9HvbFKhO8G4H4c
GaGrKAG+GfzhvxAN8zEixkuYXJy/kpV60Bi9sES6wQvXUcspnBIEzyPH22i8uRXF
cTtVvFXpkDx+E0/7gie8lIy+PXsuTCACG+8V5U5zCJjq1nekohafE6T/RKUogDFq
1uv/LR7eW5cR3SVIDOLLf05ntUipWGZdyXnWAdECfzn3+eq3tv5B27UxjOM9+VdY
TSZSEAiLIewbwNshjwTklP4YSZpzZuXt37CxYu/skutjQccU7NCJSAI7wj8iA1ml
9lSJmwGZ73A4Z9BsBu5C9EsmPvNzJQF+pLssVugpz7yv8cvNSl+E6NOaXaRUI6aq
Bqm/UpMQdZ7eL00ML6lwpJshbOwqjHq3J+/V0LhMMEg1KH6y5fkmEymm6E6lIEu+
07i5SHGl4bjCk8Q3qyHMgN5v+mMRMNNjdgndfQW/jWVvGWq2tFIjeusGP/v08ca3
/h1hqJ2TqoGPJlXxSgaxLLb0NyY1I/e7nF9475Ds84e0nVAPr2EYFbBXblQoGZeV
D5LQGJu9WpTZ4Mq/zAQyY37U8CiQLk5mPrVv/psfka1GLa7m49O4OnaZX1sVhDNC
S6uW8cX5cEF9SO9ielC4QBVzOwo/9rwg5KO7qZYfUmfaAQHBPgXmftSsfLPp+ztd
n/0IF551PNfpP4Cye0F0Vv6caItH6fWWGB/cHk7IKOJSZCBMURSxA+zVStmT1zUU
N/o4vHxiUFcsL9dzYRZsRUkJ9CieSSYj8wdRDw84JblEeDNv2lwXav31WB9hHQqO
SCv+Vta9gvLWNVCINIpYWmlSykN3nkb561u6hwshDN6s/R5WWh/J1AxADEkmyVMN
tSmUZ4myqvz5PjGP3rGv5leffOn9dQZdPN2DTuxSEGE5+DDUExnQU9ZZtKyCbUR7
756kLfOTDeRH2JMvCmpAagSTWQus5YnBrZ+kkEI+vxVm0TzRHKIg/6I6UHAjLI6d
ovX/IOqBefgXP5ZrU65e8nqRSvy7dEYnldFLkewsFPJCGwdiWoCkcdOfo+ilCxTd
28sG1F724gwzAgjuk/40ExyYhuTC9XIwL5a+GOY/R+ZQvrY8MO3Byvb1d4+F06gH
3lqbECpyNevoNkLFClD3SiaQrEk1yWjlCp6XLxf+wrRYxXU6jcXW/4VNR/I7tAGP
xxzgZsvUgP/AYYGJiIiLbdAW/Q1JcZgtauk7Fjwou74UbYSIR9X7kzrkoZXOjAkK
am5eLZaiq9gbaeW6rf97SgVsgFSuKgugVrI55Iek+mRu7u9sBmKMVfnpM/lYuHCx
i4SqHN3TicUZs+Gbp2+ui3eHgt1FctGiER/vik81+680zKaGDgX0gm+TcUmRYgA9
avpMKiBqx98SaY+wyRfYtk5/PfRguPrbfC9XpvZF3gx7UnmpfHJ8c+KZQh1AYKrk
O9gWc7ow8czdaaTSK2oc+cuimFsrXI60Or/6uoHUZtL06j7sD8yTX+ARpdX2S05M
5QGDkOa3RZwPoZEEMxuPqwmpfMtH2cWCS2ZTYKaiZgEbeDXxikXAT7lxDjCrImxj
/DXEISeiwLV8kg10n7WiKSZp6NhiCuoshhzUGurMbrNv+bK2dNbDAFbJu/Rn7i6i
cFrrTXDp0N2LnGyT6sW7llrW0Qh1Fmk9pKU38y0rOIoSVleUGi9UsQNDV1mpVSlW
KZAe9kz4p2ZgYp2aQaoOsRN2SvT/S419MoHI69Ig1zq+NZE0gBJeYMdAGyfz4chz
fvsjL5tTXLCPOM/4OS/CLscmr3zYlr2B7E9QuwnZbp306wlc1/yQ9dJw6cHGyUHC
td55EM8jGn5ozcr883+Js02+wwN4tNUCT7NmCIYn7QTyfpQOGQRf0fMNQu+L5ERB
pFCgLdWlOpbwBqn9yM1dfVZKtju8pqB92F1D+VgoXSEJR/2CV3IkoCMBlviSB7vo
VBI0DNN+4f50FJxlEQoSxE1V63L3Jvv4PE0QRnYKFIOlFOCh1Bq1lX9nQyXT1ZQ0
2ftkg3AWzGiDmmCaAUZBRdaXOQ3z+p4VA6aNV6neVzPc4N42JE62Hwlaq3NsiF2Q
a1ItlTiDlwlfIpRYbbyhlIAx3GnwpdfNtJcIdwe/mAm+vsPPFXO94rB61IrdELCK
e9q8KqLR6Raq1cXYRgfTC7/cKvvk4UeDe/MVA9d/EBvADYzSBr5cjw+BeTZOvY9m
w0PkuWgTqgtJDzJIIGyRqmHJRzZWxzXdf3HVsM4cOfA8mjhIH9xqa3bvzS5DVkLX
6H5wuzO+kOKgM/bZccB09LUrP+3wCoDUiMmrQZfKnABvIWLsSeatWa7a6hqBYW/N
yxwYY2eZLM9CqK7oIHNfMKVu0fNnje+VX9DCFuOqAVZwD+d+lN1A2T6nPoG0sbVe
q0Nez7epm70HxdPqtF039za/c8JCOmVkAZPwdGoNt3VdRQei8y7e+ZqGSHzkPvGN
jEKcf5SXpCkbKDDUfp/UUA9lPOB++C8wWg4oAGWYGAqFzLu7HPG1SXe8neJmuFbg
GvdSrnjjMR7Upnp6B/1KRmFcvvXVsRNBSqHQ38HfNNzgcgnS7APA8K9Gv8/b1Hp+
yky7e3FijycFPUs9fzGorREPORgWGg6TRM2l8UA0uN+E4nxpQzm87v7o/s7HO7ME
Oq15x/+Fj2YemRp3B1BfdEx/GYOC7BkQQxkesH5iQXiFRpAlHGND+fZ57XV3UGaM
GNtzUU8uA2hSf9yaWlAB76eOH9kIlfEeTIctsGGBQFnGhrQHEGuOVi3sdaiApfDG
evLcFNuD/FC1vnWrhAtOhFa1w4Xzq30j+jOEvzR6I7Gshvsb7yWaGmvg9ZodlT/e
wtHiznzgKr5WF42Iym+HTb492Cf0FynXFl7AlcuF5iC5nPBFHY11Is8/HOSUkFa/
ATYDY7f//GRQjuTAC39QT50wt6uwClIOLYCShdoTKf6Q5p7qrnHLVpEiak4FUcrO
ZzlCCDpButyfvY++JclziPghKm2LLMnojtfvgpabNYM96xa03JbHRkSPyCcVdNUa
J4ffrj0Fk/ghxIulaaTPGU49YOztgpn4ggSqrSq3jCH/VZ4BnxUZmVls+mE8kirl
rHpi+SKSyl2SMnxx7en6IIDPe5jLmevJ+cXTE99ugN9e+HDl8oWYpcf1K29I2nsB
AhL1nu7aGsJjMBBUlndhGxk87j42cJ+FAXlsCbOCfLtcTvu36vS5w0tI8llO1WPt
v9Ce5+0QhLlrsahcgJDLYqAy63g73fIiSXTAYZRCZqjaZuFSSQtPEfSx0QiowP6X
GXMwya9GlZhMgahU205rdQQdqlvDdoGKPciJ5uLe6g++YuHPj9I7iCFvWarTI9mr
o/xWieBfoeA7HiPBPbkykVPlZCZ+5yBMRBO07MdxekjeNYu2EJcVA+zzHIgJOoAg
K/YOa6w5ya6R2mEZ/fy+yUrHEijkW7Mn+5HWtoxTNOEj8VcrvmYTnI7fIblJj33A
hTm8sZwPBZtl4BRSGvUTpLRlqQmtg5BftpWppnGSTgSoB+vDcxGcDMGK+X8Zp+yd
IUrU1NDNIVGRqgBwZvv5dyoiNXCSZ34RNfHtDwv7RwfMSNEK2zLyyl+Y9t9FjckW
ab0frbVrqwsXBIy4IfKbGzl7wyG93+4HOMxelJl2ndlxl5Xiht7FixG/3fSXDQp8
AhhghBzkK/RjvHmyWWyPOSWWFeqnC72EkrYT4fclk3FWWLlxPYL8/KcM3GWZYzss
KPfAW5ICP+WlahUsqpinKkMJlOyLkGhV6jgoG9QWlYpLtcmYcQfj44HcJssq/hOt
scbtkLg8aS72zZlcm3ZDbTbM+OHenupT7ZbFKR9rQJNVWO4OwVFPrgPGQ/DGigf9
4pLMhulXJgHt5q+Fn0q8sQSOFieLRTohCbeshvpxv97JDcc+NVD5p/yOOhtfnmr+
woCSJUyfuucdjHyVeGRzVTw821jJnEYM/hFXnH7v+LOGjujGrUjwMz01omsV4NCa
gm/zQhg+XPpDf5QZAuf97a3hJ6YfHUio1NkegeQjdAlFTvRdqrgrDXqsE23JtQFJ
cM9k4GjLHxXqAgacjtaiwKkpgamm4TL9KoIN8DjKPnX92ocxHYnC/5r88QwqKvDr
P2eDZZ+Q2f8frMzpiGmv6nMykQ8aT0obDMTuh9ACiDNw3+2wV97oe9a2ATtww+hv
XNOWfnfY8oe2/Eu9OBYOh1kyWkiCa/ugOG097dimhzA54FKzFysUgn2t6haOnxK+
lE2VxVuXj3AksUgJy6D+Kr9kyDwPoz6Rj36qhv+Vgp2KwYMb9gAfo4smU1FHjOmS
JAJGtTL3Zp1P6JzTqEpZH+14gEeZHmnR4Vmto3lFzwOYHDyXKHz/fbePLyebRS2D
afqexDvfNPPIt5jkwyMLvy3fTiwLpI7IlrdfpsrvdSFsH8wnwg5m4bEEX99grBQC
CIPYUQG7w2KO2Ipa7hQKNYLKwu4MXLMATyDFgTFQsFQE7NNo7FxlhubpCFmPHRW9
EJDZ/YTK9fiRt8Qw2H0hTYs9zQrfES8LR+j9Lw2JdZ54x50WNsd706D92rEq0szH
XqrMMgTrKNAVj3Ifgps+0NZhwuUA16c56oz5wHkaXJNmpMjBvnIcR0iY41YasEtc
+OdRwpf3lBvneMi5diLYb0lr0LlwcQNKe/FingXtR/7QLAP8KfojXe3f4E5vrpI3
WT9T0Md9CFSAQojjAytW70iJaMo/VmBXof34NOOpvtqOKktPCWg1UZUMOFBbQJiC
6uK6rZAxAFDDr3FWUvfFQynpP7XYSeKIqrlzD+ea6Jr4c1NWhZ8af0s0qsaEwnEF
bmovifG0Kaqk0R+Wir7K3+Wxk3bC3WV1QU4/9jH7bCS4ZvbJnu6vHVJZBzDzGR02
D2bjcaoiCz8LMfvc/ZfxFAaE4eFFeCT17pZjYvdspETcZhctg8JOWr/aHSxILv+4
Wsx3v44LO8W4f8xjZYeEkWhANRfx5xw3Fou2nPkGMZrnUQPjspawINF1Qjrze1yR
t96Q0ESjWWcsiLZNyzgf9Yn6XxoI6lJXLnh6VrLkr2ZNLgv/uwMq8EjqvNDw4PUJ
1HiX0x5AS+PLrISxjOKNkMY1USUiObwJub46tVrqP4c+0NjTwWLLu/SdRjagICLs
WkBdvpw2rb0kj4b21BNESBTXcUusH0bSiU+6d2JAjSwYgqT/a08jeixzQQbXJvPp
rZkoiyQOHMcfEPc+q4ewrNF5xLYQygJ7IFQtEBMyvgzsznYdN6izoSM0bQJydWEs
cVfkspp67cO99ihPN5lX2u70PT7Wc8pND58suxeGGinwv2iYkitefDeSssrGV6X8
Wiq+PcGGPtpIrkJw1AF7PMfcFMHnjyyLAhsZxNpGARjYXyK3CECHuKHOY+wfqAgR
i/WkI3Vm4GM4O1Lh1mNlIRateZ3Qa05VOGXpCksyhFmbZwSixX03yRww0Hc/0cjp
TMUNikxJoqMc3qG9LupDMZVGqdAralrYDo8YrB8CbkmoE38gGfvnWwxRkqhEz/dG
OBMSX8XEfYd39124h7uxjjR3IFh+sqU7r7+wDK6QKm1HJ1kQBiVoLgCwJ3XwTFr6
cUaiy8GZlQJum9qeC2XLF/04YiUKbK4wwHZLLXSj0OULeTx/Bz1r/9oo4KjBROAy
4lEZoVKB01XNDhvc7yv71fNzfAbqtJ4O73F5WhB6Xi9+Ou3vH19eD5pwCs1iowWP
Nu0YFhGWw2B1J47Fc2uJM6KgwxVgW6afP+aFRd1S8QWvvY2ASUoH7CWWl8NK3YRz
qbAfayBdn4VhgYewx4yQYZBZZjOF+2Ndaj/bt0omyUWBOVFSbINnh0xfWuWaHDCp
VgJUNqzF7SFgHHWK1ztAxQtEP+97V/ZjckT1X/8l5d/iJWd8DAHJp4/UfdIXOs7x
nANj2Lo8bVY7CCeUz++L2ivMvrLLhM/LsXWC6k9Ap4GsAAQYfsRJ391VlamudkBR
xfVMCRPDNkVZig9QcaG0XVERnTX9IRWXX/7rLCOfEQzGpji+EUYZ0zE6WFMLKr7C
WxNKdXblX/juYXkwh4Kv1nIw9pZSx0wCJxC8SQYqkygnzrpXWNkSK72LQwDGW76j
asLFNdKy6n7gzJj2tX7Bv2jcGn9KkxsqNmkmVktMzfYjTchJCqwDHPhEAJqpw0sm
YHyNa+eQpVG4RIPc9z6k7P3lH4x+W5I1ivaBvsunkqEVkHqOP7vYyMQmUD+SEdEu
K2okEsZNfaSp+I4eVmnvLn+psxWmCVQJ1ijKWjru35hgruqhNRuhVpeEHaTiQo9C
VAs8qU8HegxDK+4ao7kQdIJKLQFrzctDEW+gVTR9hQKquhdQ+FydzqS8/PlFoTtz
0iFOC4+yWH0nJuEpJsqLOIQrEm2+bXvBCUGlu8ztYV5Tt+PAtfxK+/mfRhvK9fno
Z/w6D1NpqKW7AbdgYCuEWwbJpyMD1Mj8u51GRwOuqoEkhT2hsSiqfujgUADIkpGB
ubCMhZpJ1jsFLMf1w8aaXYUmODlBkri60jY4ZoeoiDxVt8TEuJZCz2GIZ/pV4EMz
DuxtVmRl8k+oIUalq0gkYbdmI8HEGaOHcl6x/cT4mCH+NkaNI2o2JM7H9rEnbxcf
FwRoZZnQpAXiw4Udo9wdgl1zjt6IdU/qWfXCtCWHrvMu0VQ4cHb26CicBNtKhEoJ
nvh/O0UfApv0axrA0I1oBxEjrtY5ZHoQ8EYhxBW8bQDKsFHHvhcU3j+3DUJylEAs
9oEPJok13b0C1y5H7TLFDgG/2tQNDYeUP4ohTetCTr070zbpFNmVMdbGC4eV7SH5
yioCH3OTIktZRrVVjkprba9Nk+xvKhkQzs29yy1ETyoziMfth9IXz4xiHQ+DD+b6
RrwT7ehnc1TuI6RgC2jIuQqb/KV/7pS8ALg0A6EGRKb3BeT4gSBFQfmPptb/I9+c
hBJFVFSsaep0cqBg/R3aSOXS+L/UFPIU1D/clhcopr89hPiTRopa1VORKuyxYCeu
x2xAeRgWrAeoA216HNFo7q68KjnIWBmxqOXJQiBHTmFjQToGtMxPF54hkn37rPJJ
kY2bxbXNAqI1UfaqFbuupi45sbfWyzksThy04wSImOpjNvIFU6cZVbEejNEAKOYh
VzZIBqwi+9IIkAuwRQv9y54B2fts6AE8/5Gqcfk2766zSMNv2H2aK/zlofvMY4Z4
RexgIE2Zm33OVKd/ucDrfYndau4XrIC0CScg+w9/6Q1J6De4SCgO8tOra0ndl8Vc
zkTkbDZ+P7gHFPYRCxszcxoHQ+p19D/TdBEwW8TaPCKtvX7LwBEEJgxcYoFVqmYo
Dk9N3yrm/o7Yy9kRYIxWD/wB2oaJgKkb9eHs88WdKzEvIn8lgcWe1Zb2/0qFBjRp
6wqEz9VheiQ7Nv4rZKanq3aDFMcQJwU+oXsLGlCjJCQzsJHTcAqL3NSdstFwYuLv
6y7urVB11fGFM5uMHOyp0bMRmEIz1QpC9IF2ICywntR7xnKJfsbGBFS2MRBGpY4t
RI4He4Fb2gA8D5ZhpByDcmbAPCZK2JaR9xnS3uPjC195XtfqZzpuoQxo2MR3Nxjy
22OVHEjd/T8NQuaimWZO75xi/JY+QPGI9kZziZquoFRF0LFA69Q1YA93+O5eYM+2
N5uQtePGiko1GFRG7xS6KJaZqUrYgS4uhhiNvjjzpIs1RfRwa7JdfKpPoOV6quuf
UDmuV0Gs9B9Vh9CRBdkB1i1xx7UMphgarcPIZjk32fopk+ZLalGxeSUQkRbSMmOt
0Ve/Nwyd6ld5rUyS8KZO+xrfcKxkDvEplEnfahtLJYj/zjIWIXTpb+8FDgC2WJ3N
mzU+1Xr35/0tEBu7Xwt/1jXlAWwqu3Av4NtiD5Jj0xkRnjRLS9Rfz9kvUSBHuW2A
i8wXsPbe8pasyK101gyl0WWwnzj/VtXeXL9NwdsBbBeoKoFiUZqcPa2uWrGoqYbP
/MVKyxgmj1ebBPDu8kPnXeLjIBjVumdST8/1Czha5DaFzYIAS9JbC6M2+6hb5Csj
7h96Ic2JutIlFHW5YVnfHpUhuIFUfu+qLZ2JwpQa7sOUEdjHndi5n/+5yM8qIKfp
MVy85pGdIhF6vUXd3pmM0NDnlt0mKUsdcah3CS454fB6CDMUSwSmVq9NK7rbCfzG
5P7apuSx7U1A5QAAERTJINyovv+VQHRzqDt2oaz1j1GpfUvoVkrDxUZ5NKb65gS+
8s+9kV8RSWXoMawhEuxOiAd0BrFzGTE22EdudosahgvLjgQCpQXleQx8W8NVIeX3
OZDQrP8gacaQhSAdM0/0BpY2O9EnG/ywpZC/d0CzfdTga++m3fv/y/Cgk18dltEh
WIS670XxeYTcwXPTdKH0j8997tDtA+TpjLJWIk1sxW10ozyrNJ9vyH1H8E6mGYm8
O4gbN2fkASx7m/Z+WHphgl3YDZNRh5/o6aw7+95zEqYsDPjldsu/fqPNP+rupRyx
FnEmAWi1bVguniQn30l6d6xImLR2rIhr5J4p2G5IErGKhzfrDTHEb5opUtF/ozBw
OQtbH84cDJQ2rPEnUFC0EtC74aNgWUf3B3PTZ993npIU1PV+SYd319ZAl3WbWPOD
OOJUAAlfi5ft6ln6QtI1tRt82ElXFJlYp6YzJE0f4Kpsk+XShRujaDdqcLJtRBh9
JcxdGkbn+15cu4v0DFv0JEYO6GJYHcxBjcxsotE9ZlqBQmBiKjhCPGDLbinBd1To
QbVE3qqYRlG9d9D9rXKqyCZ3iH9rjvWPbxPEs6IF7SZPjfU51e8Bi1f4Ccqg6G7g
PSvIHz2LvlOrS2IlkBH6Ft1RpXNzHWw7rjlp3MuBham8PjAkF+2y6sC6pk/uBi1M
qazXtW9sMSCuepF65LoWhygHiIs/eFPrkTodQmvYI8bQv4Cq+FeHU3XWQA1zg1v+
GDXvwDeXxWDaRFf9hm2BPdBIKftue0wy7yQ/uLauW8eiZ/imyDVDC+Rz5nxQ7o9D
JpdSL5JdyExVBjtbRcPyXFoz2MZSUzOiTrRTMQXmLjk5dyWeeMSAsQcsq8+/dq2F
Cwbp6DqcaSsZgZFiDbvPbxVjyaHvzWkgqQ1HvOFebwK32KSJ9IlLel0nR27C+Qs/
+YXcQFoOqp5fP9akPB0LDRFKsyEhmnS+VOu4oTO+didxyZARQq5dW/4ZY2+69bIT
tasJSzux2lcLfc1okcRuS5L/GwjTKmZzFi4uT7Br2HCRU8r2oxhqBhuIw06M6Awm
0doLWWEmeMmTtgj86NKuJ+nUObnA4KHhtUG7NF/grcD6svr5LnlDXYvez2JWFejC
llKkOeaMCRj7Emb8zOcxlyqt1Xg6DeVdlsM97u4DefW/qKfy0rLdxUlbT3YVcKjm
5eylad+KavoyQN3ePMOyLKWj9wT8NJmI3jltbw17bCSWYISpKLQY4k4njA547iP7
2gUzvnu1WwYshDbWPALAprz1n3g3LERp8BhEW0USk7gXQCkeG8mwefEGmqq2ZgJu
oErpxeXak0hUZ8P4H15JXcuLVwX6OCGIp7kpH1EcTUk6cy00CMtzD3waA3++IFgz
fFu6MklNY8LwOciwUdNG94JZYqGljPuOn7uKQpNLTRrchbqtHIWW2gfkzUrNir1T
j8lG+SH7j158wc4dj9bGhtd84pseue1DCU4F0L4exqjxZzRwv2YI7/OXoCAeLL/y
oD/wBIihPaxynMcHxu7Yu4mdkwStfcwVQMh2GGQtY5vugYSbdFQxA4/ukPdyN1yt
82NaY1ER9ogkxllq0wMqdPGUIsvOglNzAiC+5KpZ4VRjPeuc2TlMLyV04zmZ2Ytp
D2Ck6hG7W/KK9ZndTggyefwfJBEIN/YDr1PL79ll3SHy6Yt/5A4HW0UuFtgQm3ME
bj9gai7bbsZIhr4MjsLhO1lWBfykqg158lZVD54kuJmBEWXrxwVeSOJGWVYehwCP
vJSMIPXd/fAmtkorK4VReCjYWxC2gZOedW5E+nEEQpVFqEI5VghpMLCTrLB+G2OF
fucMhaXVxPHHUixHOB2qCpYv6cZleypqoO0G/8ex3mB/Kc4JAI2OqShINVfSzDTJ
xXVx1mp8YUziZrELIuIHjz9NDI72pfCa8aDFCi7k2gFFuC8qNHactXq14pmo+Ucx
EIxWngurZZMYH5b+Ci7SInZvP5j1DMg0jlCIb4nHt7rVd2SJOjLGdlIjigjz15ur
azIm8NkjSqfHCRsUKXz68FvTrteuU61uRpd2wzdFuZoXqm0oJWrFRqBjdOithniB
/20oVW4UhPdZZaD3IvhUm8O8RpAreRGZl7BdZjAyoJjHomqa2G/SOLu4SqfP+Q9D
ovYgpnx8xT9nAcGgamyMkjHLhZwW/AHVBBEgMi8G7yfgL6+pNSamQ+bhlng+li1z
YXUgKYjU45NfLawQbhSqViqs3sTdyGLlpioBoWyBKTq8+IarDbbRu1JD0L3VyDIp
KVOB6I0BGlqoxgn9agBMY8y+thHCuAcH9J87GZJwDRIqyYahLNd6QI9isMzLb+Ni
F27r2Nm/Z8AvL63lFEcbW3My/3F2ce+D0eNdD85j7sG/eXDjW/4IaRCNHbehz9Im
+Oz3CXQAFzHaxBowKNnaVmnsv/9Br/XjIOCD8yF4KPAwOTUKU9r2bCUKS6RtLVrW
o5eyuDrzU+wAAIhUNCK2yD+K5LUu8kXATHwOwIdRiC8hBer27AvKp29FE5TMkrYV
A2z7a0Mis+mU/ZA4axngTOa/aQkeQAf9pcwqKM9kJ+yYM4N+uh7SHugeKGdVwcSs
0BKJagmShzsrwh4o6T3cBQTaVB/ckLpnkqvlQYP+kGMQc2oBx8SKaHzrnPAr+u21
YGFUX3hucJE+6qnf6jRI2KQLYAMNGaIYhz+etGKpswJKuMi38dXlAAV2Qc5NU2W7
avOQaOgUNOlJ2nEcgP3zdcF/Au896qFHNi6y9+NJcI5nqfFqwunfO1NEpcUFv+wa
m8vmbBY169FM8xR+LixRsTJ4QsbulT/2LzoEvPPVtNqzwhawMYBa2DzkoHbUv7Bk
tRGhIDGOXAFx97bbPcPyIe2EzslT3VLJ3p8/gWXnKd2DYB/iyFpX7RKJ8ih/ST34
Xx8KoPrGfX0oTxc53OxMG8lq8rpO83y9jcTRSN1CDZgR4pzOvXSi+ytyE2KKTVIs
A+NAUzKnI071t0WZJ5pykqwtf7y6RdzL/YaqsX+enHhvn7KxolxiJtcZdweH95qC
nLn763sUNQDR7QzGoEPsOkC8xHtBCZYlRX6mzEyNfFpjxiqviXB4PVQpdszJKwfb
cbFMWVtWJg2s/zbfFC078JjVONKJ/kVWXz6LlTCgs2tGHBTMIP3EWmCXBF4mODeA
ewnu5VOIh73qF/yViKQkW7g6bsdoXKtoew3567hwxXH5V5qKfZ20vzbitv4uTCYC
739ZtOfiA4FDUan3aU8eVmB+d7OJI2BhCJA4vVGCHRO9KON/aRPHrto2MDVGf3n/
CDlTBsAC/lw/UE2hch3Z5BOPq3ZetyTu79+S9eAUS18WJgW7Y/b9fvOybzz67ioa
D8/rLfMJ2fM/eJUX7WG8MkQRR2tDMIPhykv7VrkdhJW19elADB3SVEw3V0KWtVC6
6YHJGoafuYS/vsGdbpmOaxzaSJzZwwqkKpyOzcUfegX/WUprWMjpWk993vP9ZbpW
6qcB1c4bpCM0E3pk96vTY5GRQ2PCovVBH67DQ89AyCEvoUGrjmHF4e60R4oEkwc8
gz+47Pq+/W6TCdjXqhDmECys3xJ4l2wVEb80sxGEeljd7VGPuCroiWtW0dqeTO+D
b6Vlf3IaicI/mZUUKAa/FD2HKmsUkn9rhuP2BYVteICJT8vMyIeE4l0xcm3iQ2j9
faipJjKxxK9OLJqL0ac+0AuVVN6XzrIoqew1PdQJ6qzFG09syNVGpkBwQZcktZkk
tp8eAfc2oLopESh6rDXHn8PxCWYniv/tnY/Ng0qcEeQqVgSHj+jXnHFjyzPBAH5Y
R1mqrSEFMJlD03rCPJXcpy3hgWCDB1djnkgm3aP5k1B8o5ajGYOxxdWulHAuyM2U
xWcS4uTZEgnJ/wa5lF0mXVajA6EWd2ETLkVUvnLrRMoLRNLlpjy/Mq/lT132yZs7
7NPK12TCwlOKbhHj9Uf9mnUxf9uCE7NhJ8Y4N40752V/53tEbq9oIehZicii/4lD
/ZcO9JXYQMpR5L6LpcG+FCpYxAfg3IQ/DHpgyHGlAfVanTCwzbxmnPHogJ3OCq+T
OJxb8qw84jtTE/7ye7nauopxH84HdmShIdeYhnJP167RkbM1PZHk0YcjyQ2ckwzn
55ySdFRznIQ1grFzluFIFwi1v3nkIdNvVqlr5zWbXVyLDBH6rEJYiL2HsCaVl28q
KO4zFvt4cRMzXi4758bsGOKtGgl6GHmudgCdEX5osFOBqqEGFcyVjhkj14sYrF7g
QHdrJMnXQOn0xNiJ+ZqBAcPFCZ+OQuWOsvewkblDzYC/zF6JeJj0bROSd0rxRCoM
kS3HBr1X9xtf2nEUZuwsOyB5OulXRYNM2aNYvcqUOb8BZPOs/ZddqsSCmRgURsQr
VkWYUFq1quwebGp6PoUUwKgyMhx104frh+4DCiDZZR8Sl+4JpzclQjM7onnKp+tY
jS+5OJ7YzOwSP+j1byAOC40n0VsLKNRXtlLwo2ebG7A9EispFxXcMAy0I1o8DUrp
e6wrXlBKvtlx2fWbhUG6Nc/CuvCEidGpNP9TWs2uH1yKfLqA1vOhhK7EvuAWroS8
AKVrdW0f4YgagsxmTz9m7AiFpCBoYkFkMdA6umDbIl7hCvOjqoqTbRnoUh8iooPx
0ecwXQUvGlAuFsUxp7JUIZEXTWRybQGUmU7avlvflKJYEBLy9ENbCjsfowXzCY32
cmqD7Mwt95m+8wzLYHC3ei3QGwucMxg3fUy78iu6OA0AoN2l44FdRjWm3t1aZ0xa
yoIkBsR/9iCT6bvSqb5L8qJOZJK4rqbQ1PeAQhIeUFApRqHR5SHFrn4X4Xy/bvxV
2tSy04nV1iB0ziS8eIiUaoxxnF+PHju4nSnKouYv8qQ+3cvB0p12/+S04aprKwoR
aRHUsYNFLKnHYj+RahrOtqpinqCeANtW5q6EplFi27+7+8DHS9TjBzv00g2+xfsA
VhO7Uf4n84/McM9GQqxpa26UPbPofINvmhCHIoO833i5I9GvCOMqDdkfmqE5D5Uk
6JR/Qymeod2gOfrz1oyZDbchcqvzAbPSUDrCTbz7blbjxsj+fjR1OxjwT/EYyErj
/9kud2bXKfO2LD4UEIWkDWvzNJrRgZufBMSArcbWPqK+S/mrg4Imfv9vJVhF6juR
o9m8kDpmSIJQyKRfbiqe4VkSffEp0Yfm4rBLjLBszC/6FefgPcmCFlZYH3PWVn4j
0LusT44fMCJUTFgQYZuf6gx4Os7+3lkahrHiwIXbOewcCevqxqWgH+NK5Fz83iJC
jU1oVbtMAiCYIDoyYGA8abudHzNVe9261RK0502dYEpQkHLQ3LUCMKEvechpEWIl
9fG7Dnp9Rp+Bn/VTkkqIHX3MbRG9cOCsPaBL4stO6wU5S2DA2dCGpf29hKRxrAMI
FnDScyf2dNelpXR+KmY/bDNTqJkSLDKcI5PyNwwz23ayYjZQdW05RmQKxUr8w3lV
itBo8AJNOiCvmw8U6F6kXg3eZrBEYjjcHeHqrHAJp6uyhC1k5ZoW/f2mGqlLqjzn
6nKV1mkxj7/Pws6fRflVlLYEMR/4TAvBiKZd5j/M5eBn0fysojGlsL0k3HTqvdrb
XWH9hXWsKMDG/NBaD8vb08R7tG/6DV+VAzff6OAPlBtZnkmJurw0iA5BG5q0nYCA
VVKIu6o0e40BL2ICaJhNZ/Xi5bcnpI6Bb+rFitdOhnA7wOFZ6jFKNCH0Yr2tNo3c
4LaqLFlhShaVAPL7gJDrwiRMyKP91sHkajnsrtUq2gPU5fmI52FsuUqgI7qgkNdU
VzYcEmBjHy0J0iqnCYJChVSlAVbeElpoXPsu4QgtNRZoeIpYlzfF22wMns1Snd1O
ci9+HxedVbY236wKVRu+ZuS9DWZxQyhrpK1u/KcVUCul/Nm8eMZMXNg4EtEJzaVw
mPcWamjebLedXhHsNBor48zl5gYCgB3pNtN8qA3zX+Ex4dKpqWP4pHZDtXXi+ee/
4aQk8xtj/pXRCK2pEXBhJhmG/edIQoI6ueUUL5kUD8nB3CyVKEa6eu6fES0JNCdR
6CBBVwD9kIRYUXh5pu7DAaKs02narysLHAKJV9ASgEieIzEy8jcyXruchtrLlVQK
9WZQk9lKTC+4BRGq55dHoTXYspP4GMqpX0XyCOh7xAIE8utPoemPl217Z5LDjVBW
ujJhwOJJlbQO0tggEFUvlQDQgOqj6ECDaDATB/yCcrERj0pKbp3GGgJBQPg2swOT
PaNIycfYjLNEKOz0mTo8s+j0UmOKuYcPBwTdWyvG01dgYuz4rr2xrOrei0og+u9Q
oR6pqJqDP2ws+Ieu1rqkZUK5TeIisXeH+XLg9JR0JY9v8zPFI1XfUefvS5bZXc7M
dxaH52G+8RpQ2iDLqIs0HA7sudoTi/D43/70QYGCZbxdH+pqW8unI/L/J/wwHBE6
CQplEdAONI03K8RDA598kuZLvtq5Nft+d9eE+zuKIcirDzu/6HugGA/tCUkn6hK3
wNN9kgPPvu8+AqKoadcrwnI20p89Z2O7JEK4VqjrVCIqpHrcNPb6pOv0mf2Tn5cW
lE/QuEBuZwKpTyDRt0kOa5BFWLlJgEy+58AROshIq275eO4/JQQeCozvXZOCw+cs
5549Bnu3IkmDr7Ln0jit3CGAjm7ugIFqLSxKqOu8p66fSFbAztYnAKjUedxJUUuD
4TTMEdSG8KpNcOtTJYgt3HXcw1XOIPceqexZsLDAZod9V+5IVG6AxeOGGN20J08y
1GfQQoMM3a6YdqBRa7wunQSadFok7Us58q5a9muliinKnyTo7OM4+tju8m6mCCyW
LlkIWWuErDlwxZFdrxaC5RhizEEPFKVmZlwy7R+pOBBsGIKYUPn/LdF5YCPjEbmr
UXO4Pi1ULmeXHZWKR8xEAWHUVRLeRzITxx0GhCfabToGuldG/6/LR+wOVo30ouN7
Ka2wYreQGtbh7xwu9MI/b1Va0QhlGUgUtKukjviIv3xKQ5irStmvM5UYROhsYPfn
ciKzY65QNr/NiryvJiqwxrU8XJ8F5Mhb1jMCTvgvynAGZqs+spp1XLwnWlGmNwjo
5vYRR1I7Ar1fxyOqOJzo5UzbFt01Lq9/x9qkf9UawxzjVUsYQ2bkHGFexwbRKvvk
HUbo+850AR5dUV6dTTejmneDYWXt5ryR4dMZIBYYrfkuC0MFnUpu7ZFLAmwH/wPA
lkrR1cfe0Sretvotg8ZGuL9D0+3COulnKrgMakN+8vg3ilyvRoIUN1jCIKiWMvIb
3qXpPSqmBZevjU7oD8c6smKBbhj5YRMEM5QqjoRc6s3x2HqVMb1INZw7RR/tJ0Le
nCni82svq8xoZUGSJq5Vp4xNxzPyIKnSd46WohUt0228zZRc0xuKBWLTZar5f0oO
c1iM4ZEvV3CISg6JCBnfEjqlpDGCfy/Qcpo3mkBQIbq0dwD0P69U5+Ii5ZfzrTcO
4MRrDiHXK4DPL+PR6hGAjj+w9ZdaiRM4hNkVjBWIUb8YG6a00eI5k+8822jkUWCY
sOEw7vlS+8sl3MuHPZ0grgwOgbV5RpWNN7atCkV93v7DhBmRsOxYZ7CVbQXFyC82
JSUc4PrtpTueLGuVJyppKUJ3ztl5ZfvqSH2SSAJmFmeMyj4Bx0FPb6h/K/dFeQwf
mzwOebSNetH5OCmw1w7RFpiHSRl4D9lJ50SjQ5yHILuS+fRaGKBVjK712l5PZFzF
F07kDlfvKY8Wk7+O3Kk9H1nQn7+ubszi9LajVtoMAgYQndf7OIL8cBNn1mgDQ6xB
Laby6CMCmHK7zdDTftZRyW66FtbBoM2Axpx7LeLsoZq0jDHRUoaqQAC+VdFdOkP7
Kh3L0q0JCmi4NGAq3jf7klDxOa3jMZoJAMydnpjUniSLojlR1D09/QdkhzlnKL0m
Ql8qdKwKp9SOxcw85FVqlFXAD5QZP/cq+o0p23aurZyb8e0gUvEDoEn4VXhclfLF
0sAWn20854EzWBYIPu9uKd22grFwWQOcQQG42ZU/XvXei4Ya0HVQd2PLh605AD3b
oFLKT/pPgpq2fVEtOom9NbhS1sQg1iaib4opcvZrpr6/MZTLYKcAeTqf4zHTSyc2
pjOSWUqrGySz2xV4tzJDPeYqXbjcifnU1VAaY/vQnAINuNrAhS759bQoY+u2DSe+
3qh7y9DVuAo7D3RZ+EpD+RvLUKl2+peSsmWrZuW6bTZTiTkfqPSGGeAFsHUlxmeC
VaeStgsHet6GLFlTFmqSHODQkNMYrqlNif1XgXFY5x6KHeiX2eGmbZcxCV05vlPv
GF1LHhWkkal6MAiJ8UaU4i5IX5e3+P/czmS4WNFhLWMs6cEq3bAS1gPwy0Ou1QOo
39fQUY74CdG+LMefIQxis3CgEU9cBBzRq5YxNf+shl/hpep9WVTCPc6O/Jblxg6u
QVk/XCNxHnvmZpISZ7Eel6OwDAm2wED+PdS0ybfqhDurFmupH16iE9Nw9vroFCPY
DfCssFQCZp+DsYeqIEneOaDiVOnJ6fOuwvAK5FA7P2xSv4Tox+O0MTnwLPie6yMi
jn3y9kMFhpiWEL52GjSJztnAMbVJV5NFzx4yG+CilzyDb3yFf3jlGmZ0k0nUstp0
QvIbER3YV+QU9WlpZu3g3k16j44hkAwC+8RO0Rhetzqy3fXkFwM52H7In3HBuAog
d1Q4e+aD2zKZ/t5sgXvDRzCooR7vWvnS5LDXxH0joENDW4kNq6UiKZ6MOcozZjvG
+gvj5j8CXaGHXgkSSzoUgQRMeNu7wFl+JwPCnd+0hqWga6wcVvjT082YZ2fkaFxS
S4G3RxMf4uzv/AhbOsfoAPLQacVX35jwbKuWa9QRCzvmU+VUB/bUCvKRsUkXZPe/
LEJOBStcuwV1cSA3aTBPsArldnSdQGm0uc7FxR1yawBtdil0qYq/VEtPXRPRTr6z
8/r/lzbMS3rNKeDPHwqnYMXiubP6mhQHNJuCcjTSlvRRqTS8o5h+q/GUlI39f4e6
nss6o28QznlD4437vPzqAKsre7XnBOe0Rte/VShjFfkztkhDKt1sgw9b9ofzmk6z
v5f7g/W3m6FnTaFvMwcp50wV7wYfHV2uAd0pQNILNcNazdzwpOhy9s1mCgpQmYzp
+wKhcSuXP5YyTRrCnrVR47+mGVlsM/RhN8cUsuvW+JX9r2w6NOd7qtq5r4K1pQGS
HRqAyH/6mKD4M+eFnUHkahLvNZfhAK/Y0YWzVv3yjxw0T6hA2UDLasD3/aCG0FGJ
iG8ZrwV3xXq3H03HnJm7q6bvYbltvu950/e6DoTy/VZmctB8oIO2P8CLXHXAOj0l
LD1a8UW8fd9bpU21HuQCUHOb3lxngPBu5jkE+sQkbJQqcGCiRl905//B9TC3ZqYo
xKLN9s1pQlyJEzSQb00zsXCcLFOQVMim6VIkoK9Q+cPOfuUj3WwIEk46Zs+yZ0s2
XssCUmIdDiuVHtu6ku5/WqqE4Vz9Fm7C2AFVBE3OvqKnFRZMtePScoobfnEq+bcw
9LTS16fQexbiOOsCKAir4teM+vMV0P4toa3pQrSIn650fVhGzDoOAGL4lu6BnwMY
Dr3lS6K/gc5UhrolAOUrFMNC1uNp6jZWwBP202Wx9JMLiDfrBtc0g5FspsHZDNoW
A1cOv/HMqgR6AmupFbwBX5V8rzK9nSG/NBCSFuhxOgorY0Z024LtJgMXbiz/CQsY
SWsKvyLjfkL6r4oyBve+6Sw9nQmTmh0Y8uLLCK8AgDjLwPgnpA/V7XWq2YtVHPp5
Jconu3ksSax0uRqcJxoQ/vUFebSgSiYCcxi3oOezfF0thZcpqFFrVhrt9OW46k7x
CIRk0C3aQ2xh6hDB091ZSQhLXxkWvKsfCvECcm0lWO3dmQ0VCXoK8t7ZIXCQOnPj
ONjH8uUtAmrkNhGSm9x3/mdP05ukjzm5IqoMMSbQFsf9fchR7/itK4DavF77J28M
6E0SzcE+kPkWsxMx7pCA/HZGOKMj9vxLR7XJ4J/fq3G1hnb0QXpd3lcJR/LkkODj
uE6vj9cxSFW2EC4WjA1FwM9/ZwCVvpDvN5/WcuOwMHa3OAXA37Xi7BVAYOEoPq+3
1n1+0imYoBjmVvA09xSLbtNE5TgSQNI8VC4gRLYltTrQUSrDF7XgsoHhEsOB3jal
OtapiejMRfPw67+mZeIMGEUF82G2F9ApYid8ax2kbcgr5dSQwjCvt75DqddZeAz8
yWCKEIK2cNrvFzjYJCskk9Q8h6khzRTaImng6ixe8IjOl2dYdejNicJunI2X3S+B
WavcUj/scqamUATNbXJYZgXz8atFPaFcbMCGlJsevfx4DEBJtjqSLUesOiF/vTJB
QFZk+2N99KFxkAU8e5u2mMQE21yIAvZwiARuJY+L62tss6d6E91ery5rBTWg2mvN
nZGGh1eCCmUkIGX2BozMpetfKcvz++Mimb6G5ZvHZ4NwSPFpkwWr1cn/tky3xBhn
ajbNs197HYgwCcXOO3JgAa07iru6d6lQ0LxdUWEEl08i6BVWOUT4HPfq77HScSMY
B4oSTzhL1VXgpGOqDloocGZgg9EyPFQ2L4HKRsF0uY2YjdAOkSseDQNq7UBL1CvT
1O9/Xb6nJe6jzL85DxZDy9Me5hiOqGTpw9DZ5DIFQXQneIyIiN6dEP8xzmoWWfqb
Tg+8HzDqVKa6XZlSWRd5WxOUvhXtjbUaRaZJSjl0VKEtNd1dnQYFLXjyMwdIY0+s
i5KxPMNQ6z3wO7ZYE9RxSZZsVoxNthgsOEgEfG+k1wHViiK16ftrWpeR+fWCz8CT
gF7M+OIpr+kq4Zor4Fs3nHWTDAtuOQAIhvgPV8IS+ykft4nxRmOtXzJnWAWG8Ikw
UXAXV5juSdOD8KBnHoXVbu+6ZxE01/ch3IgxymJylAfk0RbrLngqgEHgFqaHpRU1
E4oiI8VUyCfq6aYDzmvnWZWrjQcJt2+b1qBhIvdpm4eg7+iymRY4theMF5czHKMF
Yhu2DWiDi/IzWg26A4kFRd+zXUpfsveRLYvCp+Xi4XQuCV+pkISQOX4STbUvM1iz
gAoc8UsU1UrWA61/CCThb3jHzkDhiR6s+cQgXSypJzYU/WM0hZ+hcc9l2ElToZPJ
FKpPJaXh+9iMFmpljjnD2inh+895uMCsEuw81sKTG2zlbvgJh1sbPENAA4kFcFoc
oI0PavJgZFd8SrUV/nL8v8pnSTQhkg6IbCZNxH8r8Y4aZZYj5E99UxvgUdefYbDt
U5EtKaHZq/9eQ6GkC7JCX85jXHvkY0qkOE8hj81//hlS0ifvCNfWCmTgEBhAYRD9
omCzpzh8hKDXeF+yfry6OqKayE3EuvjURck6FwVXYhImAIyBeScq2IyUItsXDdC6
TNIO8e6fDLPwU/qLNQdqtS9Z7LE4+sObzQb2etETKIT0yzn8jN6GrO8z2aAfZ9sy
QrQT2o8LEH3dyM8zjP7lWtj4k54tU0ucGO+m0zw+r0uir93nIM/LaxVYrW1QB0MJ
FvzGp8lxklum8zU9JO7413mePKzIsTJQvujljmGEhtztEz3y56k26WbJf97enUds
Ba7sEHWNq1UV6ODbRUrn3gnxXoiTHbyfZd0UYWhpUdG4gB8+Sxg4hRe93U2Qv8XE
vp/ZXL1cJrRYJcsWmbvja7zIsTur9vcgpSYF/BnxAkESrINdFyBWzdnURXaHlmso
JQ9WYz1qo9Uf/TLuAT3itz+Vsx2jlRr/R3kgxrOmMgZH6QY27jnlaqWo+JC9C64V
mLKzhVfV8CU6jSHQBDd6nyM2v+tnlBczTKM4daeWH8BSEirVqRwfrZtCAMrj8Czd
Iu4QPCQO82YeEsw+NoxgdAiDVNYrqW2MLlRj5Cg25wsXksrdSayUVrwnjaRi4u4p
uxw19BLts1cBdKMF5UnFhTrtYcNQXJNrrByfTGfYYh1yeBWOmnpD8XrWd9bw4HK7
mmKE25eLRiA02cJUZqdu6NGRSlhvczKpLamLwL12vNx9nHGQUVIWszr52Y8t9fv6
WjuwDxI4+laf9bMDiV4C7nlzSF0M51CcPB9vSjB4ErnR66XenETLvyWB9luYchAB
iHrlAYoZfc+S9opyyLNw8ut428aKTlo9vJzcdvdUWIOg3IXjUjqbtq1KhgEQHkCm
QMcrhhJQ01bBMUE7y+y77kWWiKagjSxZ1RS181kydLr5fLUtV5LUco+pqMF1CvbP
CkxWC8dQKEO1FRQpkNhEDGzLTbxovQrRMx2rkDw+ASoaNemMCBx3G/thRNfhbSmS
2Ce59qpyuaVvYczhVowOr75kqju5VPkyYIzMrVlpLTxQQxPiULkn2l5tdaXluno7
RPqE1B/mpu+9FKIPMopzjkIvx+ibGvcMOGYQbm1tabTWqUhUXrC0yiD0orjxXwb0
W8N6UcJStX2LAFI1zczDk42yjPz1rkKIZzN0fWO2XQ56UgyzkrVeh5nV/mlLlVDm
FuJL/kaNyhPGb9qpe19hfphAfQFFaLGI5N2gzol/iwx79XyuBafHb1qdSbgw9ZLq
52KrFEiIvYgCiuUmWuQBmeX3+SqCJ6bs0C8x+MBtgBflEhj3v1/ujzk58yhHdBw6
bOHgCrwkj1wgOwPEAcLY5OTbYQG/IEbMzUzfvRv6erf0gLEeBN3x+GQUYs37RV0L
Eq9pBhYxJv2UImvXD4X8fvty1FhJ7UAgQvBBhUMeCT2ujMwn7o0P3Yfwdjv168Nu
nWc/z/a/FjO3R3yo+1w0NBoKfq8kriU5GxOWKEmzlX38H+uhyPTi7ymkLzkZlakR
dgwiggOBbIuFlxKhwJdOs+at2s2XhJrUOkkt66xngLDBw9uNS21xzHlmpXdKt9Fd
rvnO9JF8IZgR3cGkNbqfpDKm7q4eypOxAwI3geqI+grpkOdrh2m2ZzZ3mIICMSIS
cpsGrPVY00Z8JMi/hMuT7cZKIXKiEkFPMQxW0b+wSYLVLmAVi1APMz2Ldr+s7DTo
2x6ah4WvVcJPwaCIXHfK2eQNY16Mj10HulBM7ZM6/dEOxnCDvOAUSDKX6XCWBqj2
eXBUKXHLT1GylIHHp49IpdImU3qfs2bSNHZmCtbtGCHDMumbfJbDo4uPprB14yIR
pFaFwIGGbg31y5TNDwQ0x3nBNAicf6uJCDx1Wlwgr9FCWSuUcNyAusJTTcdndHTe
xCYc7FnvK/naAXjXCI9hPdnRm/1mnD8qNrMXu7QvHBaoVopPeEZkgejyBOK8WQQ9
/1sw8rwmsklBZWyT1Cmac9jlm+H686MHEPHSxGANSAPcsjPZBrZEHYSrJJ5IX6v2
IdAk6ujlI1tRNcpt0fNO8ttXK675alHgLlpSHeEws6Twpif5+sp9ID1Z61B0zD8T
5XESnnVi0PY+xf+HWs0SRgi197J21m6ciwRAAZV00w2SKypmF60d4aAXRqqaAMuD
615LPq4xAsF1+KNHkRfrQQMwbfOIZ9DrGM4hNdhxXzPewxB/AYZndKdfbb4/DdOq
VZK4SAz7XXxzpT+9apcHYD8CMCIi7OeIG+lg9Lq0z2/SsqkF6TKT1pm7DAty+56a
En8E2N0+IeAIRdk4BXufAD68k5nxe3yFMalcVdc1X2qo6dNMgsb7jfxTpUPlokrL
S0ZG5yXE+K5VNOGCxEDtMj/WJEl0XMqtPjkwTXzoVneZZ8k3d4xsDWHHgr6rrZBc
Sd277EfM/H8yG3ZqlGY4NEdkzCnHQh7RvI4NUUOFaGjXa4g23PhblixcsTkSvU7w
cNJde6Y3/EL+TCdCz99BJyzvFBFdv2XrzBscue4mQLbc5V4S+0t6nq5/+vJlDrB0
imG2XgbiIBSLJprDCUaGt/lgKLIZg6PUTuZqQymK9xhbaVmrYj4LKPPvMLK4tKmk
Q1VOj4/ckQVFPZttbkxJfNc9DmvdC2h1ROyqHfIflLIJ960RalKPuf707yQD2CWa
cAoCRw9WlVm6AVzqS3qlrmb3a40/PheUrf0Z4hIeemQ5GKbSDaljYNk1lHEvErYt
XcfyALzOt6PcPC1UA4Ace8sGx25EEeSGXhynSF7zIiynkXua7FwA5DpouFfaBjbz
l8bOBe2c37bu5lYAZO3m1jjdPW5VXchj13G59Z1m1cYj/e8PrRfTL/0suTOHT+qO
BO7eWSlZmRldSi4zJz9n1TmEHxf/27rU6ujl5BWh384EoOYM5CpfkPxoPhe4BD2n
7T6g591o81Y9V/6hrwBq+Wqe+RhE3JfCCAX179xiQJ6aKYlg9gj2Sw1QWEKf9GZ7
zD0ZzyTYymEaq9YmJNG8fmYbMSWOEcTdnfuHNfaO7VJe+CRoOcCyrxPR6T+JY9vg
n33B/HywdQzsdOfXMQN3yhb1fymCRfYRL66vxRdV3Q/D910/oVTRiV7zjstNc13u
K+Bdm56ba3uBM1eJ1WQVG6Q3AKHWaMqxZg16FYLtLO+3K6aN70Z17P2frN6czF12
aVrKKb5kKigZhsP1KjyGDvCJW3mHwDBdrtBZMQUV7rwHHBJPwA4NYz/E6PiK1OJu
2zx7GlBAp72wo7YtJtC3WcFyO61e6XdqMdYEyc7/tP/y6nNUZ/T0OGheAr9Z++4I
XuEMisumnbzXJOIAwu2QZxQHFrsf8eE0JKldcXkXXRLju5JfdwV6IMVzIMWjQOaX
E8wCXl95aqrib4MdNmx18CeFgy65HxoBoy605CA9UTPHKvjgJe2alP/qdrYfaQDO
ywbM6LvwaeV1drurnaT2xR7IiSv3AlKj4nGsGjP/5Fe2W/dWSrZHgmBe8l7WHUzJ
YO3Ic3AO2UvfhU1qgtCS4s9grezUQxXfnOZwYY+VJUchGeBNl03/UQYI5xjY7aAX
cflORr8S3STA2Hudj113KBehqn+jj0vPCPApWgZjbz5Hn7C2wSp6y7RO+eHYdGTi
2B++cHYEo8A3iRBvELMwne7NE5rNwo0baUdtZenZ41SztodOWBn/ErYLxEAk2xSC
blYufuBOse00dNIT/Vp4tum4WNNZDTH2mtdzyeijaUF+ZY0m//VBbbLlOMPYONfH
2btH20slO2men3VhsdCFPFG0sTQrNbQFS8RcZ7AEmtsJ/z4sMDNSPgXQeo+QIaWs
2GCXQrMYYicbL1WyoD0gGDfYqM8H6FCFYMT29QVND/XxhrXRhjQFERfAAOQXbu36
dhYO6KscglFd20UaJ88lAPiuX8mMhIAkKE3DkvASESE6anLAZi4hrF8zPJyYZOOD
uvyhfwnePuHgJqS69F6W2AzkHT5+NiD/UG4JDxaj8UOIfNzLJMs2skMYS1OMtUw+
PxDke56vPeLDLUcxgvtRNwBboSaOaLj3GXbSGFyaMc7eQj6ZIVvPIBORHL0Q7Nan
O5d4Eu/HJufaYEblALjnS/qkXNMR3Q8Zl4JVD+DS6tIJV7DJHyWorUqrOJY64D3B
VmDYVEJMpYCo+FhGXsK3+bLAyDMs6O6MstLZqt9Td2mxXv6/PXHbi+2Y9NSlGZh3
LQwCyUXYqqdhXLVjBEfLf2tm88a5rgBPxum6Hlf7GxHrotgIv9RNsMrSOYbRRyFb
tZTW9ziDAtFdUeN4as2AcIRpBcEmtuxMtGlhqJvhxAkX9NAchJCjac62rLf7zY/N
fMAihzAgPRqV989tY+E+B0DvjkOzUwoTingjlQgJiFZaBMNk2khWTadYprRf7wrK
08Sr0qsQ9tJP/WYIFYxLWk6gBwHhSeXhl1IB4/7uxWqyCv4OwjFKEhfc7Vh01V5A
rPd3UCKrhGGk5d/p7OmD6MD+FYK/Y1eq45aWNH4aFGMn+z7xIouMwHRad7PUQLYP
zZYJokbTQiHw9iVlNKmf1hw2RfJf9LEZhlJKsxdQVf/OqLf5rELjncVQKXKnvAWt
ivF4pkYEXFf7iHP5hYKUxVOCGl9we45325aj8nvsA/UO75b5M3Fy3TSoPzIdr8ek
CGJNimHPI1G3czG9P04VNgZxiIpCcd4EFyTz6c+QAhE8Fj7K9ubQ+7TkzIuW38cN
Mejzn37u0KoBauh0rI8qd8ylVCHWysEoD0yBOYmFw0x0sZ9fOcFOsWrNSe/0AaZi
XdJVwqgpdZuSVil9jQ75FSYPn2DxdImgi2wTAWdJr39RLvP2aWEb5Vfa5likEB4K
0+FwvCvodqZYHgurxd0t7kqVi/+6TwMwTGr/92KZg1d0kM1nhGzPqZcY7VfpoYsW
j9X+dJ4RhzE/TlTLBuwADxnSE8I91eHB3hpOTudpF079Eip6GMqBrqc27sXzPSyg
8Sm4PzUjX+k/kT1RQbPVbS/fyPWCDicaVZn0wGoV69PJOUFKUbn/CifCEAkTvNQ2
9f+eXRnxPcPthNgn7RjwnKK0W1RYiWC0Z+krI4XbmZai3WGjcL3rFZmK0XxOZEM/
idsuYBjGHkIpVfNo8vdHGzIWeIXBWOQZsQ7oh8FUd0LGws9AwzCYggma2wqkomHV
uoLpdgIJmgYLFFN7Mwe+0oDwWL2FdnUruoJ0vAkEUtR580s6W6UrZdXhXoURBSCs
h1aiHXiI8A6bdnmVZSfSi9yw5HcjzsR7TsO8FQOpmRUJBqjVkFyssZXLwHjV+GM8
06bx+iLRLM7vHJBZzpaSRdRo0HHUHGLwijm1GkJJS7PJy4iCulTs6Sf539yXqtii
yob9NxIXim+SwuFrmSmDNSviddYe12O0C/LnZ3kXyfzc9iITisQtEtphOoLbeF+i
Y4Dog6Q75GbN2myEcgY2d5T8f1EMWuDOjsDGSqqW+mnIsIW0+e4EJjyyCtsJ6pa4
fUGzJnxnuCNNQl+Xmgw5TebPXr2dDYZhUDpaG8XHSSx/24x2JX/iD212LCKUJjXf
Qis1WDUP0IMYRnQmHr2MwlGIdvg3l1G106WSfEHTNyHPc9U11GCUTNorB8TedIq7
BoVREcCeCV8ZSMlZcsPvP0qQA/q+mqoMotfuGY7TJNuXPWCPBHXomKTbfJIBH3io
QquJpwo2ApvJJ26cPfoxXNv6J4YHO5hi6o8ZFeC7hqkY/kGVlObk4l0cQPZz6HaZ
04dY2cZcNLkkipY+pncvHQsLTw7NLIVMi2goYPXK5a2d6ju8sK/kQnbmU3ILVg61
9yO5Q+Qbu+UzGQLBU9TSnP8WfTXzZep27rmB2wu1cxyGruUq1QfpC/HxghUXE49x
FiFjx+B0cFM9hC01ovz7I8/ftYt9qARbi85PJ137EudIdP2nscqWtf4777OJAlGs
Un6dlZzyb3LMOfIOgZ66Rp8oqOOrHiIkIi0fUBhlPglrWKHf8mhGqws2jhqxvvJR
MG8lcoxTekZf27SR1kqeoczpmWcaNUklhX6kW8i4mJzxYR9Z3Tgt7oXLcNIEDXow
m8EvfK6S19DmNh364tneNFnZzuP0yfeDBzPtj+5xu2wyuZY8O3cFXOKHVzxygvb6
KV1g721nklJa9xivwdSabPe4DvJDdGk9aqhF7xqNC5bEF+gZMKJpCIiq2wGYFxP2
GuwdYMefqCNIZZxf8kARwb/cZ3X9ZABMg8xZIOXTn7zReGks1EBdaTs5C1EW0+o3
pnuZYeU/qyjamx6jB6DouJnr37wNc9OZnZ30WvQmzn20HMkNO7uauYhaakUhuwqV
8mNvuFvLiuE0oUh+vQxe+RBDdCDvNr7jRwvOGPIQszHj2Crn4IlPLtGdjCA+6yrK
6k1sXC/90RDYVak4U1+n6lG92J9P/+GcIt08s0o0gb5dPbZIYt0nNwVOGHOAwR4N
E1kE4P1qmGhr2IzBkxPnKGtDCtjPySyDRoZHSGa9jIfjhxxWsdb3XGrXCXiCGOVb
Ht738EK0MaM+nAui9db7oc3heWjq1s8EtPDmICOP/f850vBC8cDqTIhdZcgwTIIy
dRv0ZZVzLCZidan1DR4mmk/BVIRBegNzCGxGxN43OsCbjBnaux/CYHDy5aTrLxIq
7TM7E/e0oIvlwS1ZPaWzNpt9ZGs1mopwxQlPsYrWH5wXqbY3oIdPXEfp1f/VOhMe
YB79iNmvMZoZ7a52AxCvkrlgNIy/wGIs5Qyqv1wB6gVx3vnD9IOIajfz6/6eOyJi
AwAvBfYO3oM07rvwMk2gBkRIzQ68rqYREuVSW0xVTlvN27SPolj7txEL25+EFSVH
7xLc8YSOSDfU1+p4HN5LHtnZv92wemtb9bsCbllr1jPKID+8R8ravxbSAFsisqIo
LC36xD51JfXXrlmJPj1rGI0xqcdAWZPNT7tGBot8CfJBIhsNY8T8QQwOUZc7U10B
zPomB6VSS0V/TFjTnSxgLwFkFv3AgoCZ3o/ZGxrWEStSDdnyJUSTOCXdir4Htunw
sFbQt5AJh8x4aAcVErUoFQzESUY2Y0x2gCYJjDen/VVUcWc2nQ31uXDuCfj3+EPS
xnJuE8AyU7eewIPTtJw4CTshe38ugqDV/R/SZw3/hkWyC/kDnHMPwbNTyOf+V+pg
xydLPN93aDx0E/o1dnBLNNxzh3os26FYYEzOJpXnyz1Yj4s3n24gVc/vAXOhRJFB
9pMVNUZy8Ulev7YT2J5eyNUiioGZgOo1hvwwJBnZPhH+L891p60k68i+8pakqv77
nTvc7cQSqKTSZBKHzGUWpa8wOmwGICxU165sRNFcl0Ni8zsV7HlZMqgKRNZIg8GC
m3GkWK6dLNCK30whhIUBBxzln/MgKYSFt8LSDMJT0JPrdn9KE+2jTn21qMZXxNPy
hATCkkZqkAmhxudAnuoOE0VZgl503V2OmjfQ3ox+iHTuZRsxrhnamKDAW50pfmIo
3IJzl7w6MRN23A/phzcj8GOxcGdhTBjD4w9Gt34X/cmptnLO/4c2smJAJzkhUl3m
fTo+aS54eoB8la4/oVH1WvCSK2fxDGCZYyLyDWefWViYJLw7ylt6Ax+h5FpTxAJZ
omFTbI7qSF0y89Nzl8fdpufoc4MUTtqAoG59LA/DQSWHBgVOJJz/rGbCbOSAqEq8
j8yGJvzTRkkq+Ax+4U2fBIAd0tpepfbMjrjLrIODP8XngHdCsa7i5F/3I+Sv2qsX
6Dkh7nEnKszjiaUHEqDucSrENF5oocn9wKKwS4ml9C5irz63F8l30RiphGENu8w8
j1dwPxw4U/wEPGfXB3dCTJarrzUiLEIauyHtvsGoYrZL6weQp9mmWS/mGEJpXZ3l
iOOWfXRwnv2FN54DIk06L+oAigrt3pww8tCW8/jGC814mz+bw7FoTo5loufOP6RN
sQddla3Y47v2DR82L+1Atx5//b9ZAjDmay3rgDZqAPWSS06woM3FBPMBqts1oclB
DUSDUrYiVwtHJGI3DpstxKv9nL4eidvOjCmBHj+RLx22IB6QjMTfNcWYNOzNBiKs
CRW6paelNfQyz428Tvx6wlVuYEkIz7y9R23UC3Qj/xD95Hf/VcIRFhlUiVEnbJFH
wWwypn43aj9SI8hZF7R6XoCH4YDxIqUBqKfFbA5kLVS6261A2SB1DZvPrbSdpPWT
0YvYg3PzZlkezDr7iNcR2/pulDP/wjUooKjQjunJuL1tk27FGIkU6/k2fuzeIhCu
1GYS1hgf0S5G5o6zx92Bugi4/l9dFtxN0LWPEVym8P/RgwAfjtpioLSJ0jtrZHul
uYqhc/TDpXnmFUmpvMJ7uQD14DpktmBXM3+yfRuR9lY6VwBTBhgP+Fib2gR1nhYf
cBoR8/cObgesDonoLEEIeEKpbg0aVTERJ1ix4t1Yw3QLCbfE6JUiPYCiQtG14xeA
b765F0lDNXETCu5YGJ4K3HZCmasJcnE1Twmhu/Vr9Cyf+NZYr9uonnjIguA6khu8
OIf1Vp/EfN/BLMlIjb7vRNgW2JqzcjKsWtIefX09EZW+xqB3JeSBW+5ZDNCk1GHZ
TagCjL1C7A4OFmAfXCPNw5pIpv79NMS6pjDMvqhevTSYZM9SpxEUfXgL0rNOZPDy
85s3ciZ6soXDV1OvntZknylbrTQTw/5q0OQ5O7zLlBZRqTWZijZPeqGnKJ0vFi7N
inGRws9L/BxA+EryaVqwQd2u2Gm/WsmIZCeIeg8M7828Uk2iPIcTAABhuyNq3gRR
IxpjYmA/Cjd3xljfWAsgiHyNhcmPfBaT9yO3cmPFzJkfJTgc5pQU2x4O78w8ZKib
B2834EnYzk0CarSjJ2VxN/vMWy6O0/TcN9xAfr9ojreEkwx4CPWdMM2Vr/WOsQpU
ccoCDUVe05MrxatfNCwG2qp00u28ySt83h+jjbr1u1+Wb+FVOuvhR9G0OBUUQBnl
pJ/SlCiLCqGWhrUcTYkhAjmkPoH+nEDHyiLI3M+NtSclqgxot7bSMw/C2iFgXC6X
4O245WL+kEufQBYuFyaxkZD9w0i9my3uCrDM3b+5Ygt2LIyP6wYyXL9vVs5Akiz/
ai2SeLSG++69zPCnG1PGhzLjS9UjrqV96OJuZUu8PzNoNctA+bhhxJK7DAWeO8fy
/Hp4dkHF2vNsM4hhfYy2XMhMjlOOpMH2nABIXEOuBThIkuM6POtuQjRyp42BXv6h
mGd0MBK/YJ+wPLwTQfG3P+kNst9lWE69dImt/niUIMnitxfxzJ7Vr0R93UP+ls25
CQV2eR2WvVc2nm1IhLIm5voehb1VWY+qQ0hsJlrQ48LsPm6jK2tPGUTMKKI5MqQF
REO77MJpf5uoCNhNLDA2jBij/t3x9/l8a7ZVdtTVAVBK7UkDg/v2uaxzcBee1xLf
lbZVv31B5FLbFP1Evxq7F847IAl29ptmJ96XMwLoXWYcw+OEDomxRvdCsrpJI5Sc
VvUZyjcyKtky3L7dk4PnhBScrBPxNxQm9rDLnhC1pNNnz+tXCbGKVPNV2elqSrJR
QjvIdHlDr8IzHTWcLhRyA4+L8sLxQ86+ev0hKeWyUBqHuVCl8TZGiidcOfDcraxF
Up/FlGaQYowTdmWjr7d7fv67sWlzNYNQ45oNJ4Ru1gtYl3LlnpdQEdlDgH6RcYU+
ah7WDwx9yPqgi5QbCmhQ521Cjj7snEYk8KtoajCLFcp4LTwKRa8IMVBp6N/paSzw
0TyhloKGsfxrTnJbW0cotdVJqvZp1OYWCmLf1ghtpBJC46A+kkfgDwMWc1sjZ95p
ZVYOw0Nz6OkDU9mdb+UMGc/ZG++RoPwQE6WLhhJwwhagTJmYLW9wJkCka8hRrEGC
zS0b1d6r4VJOIRBCaEd7x2lecCXl4kej6GcUP/eeC82qy+wGN328ozEBASwLToTV
aWB6urT5+zjZDzgTGMGXE0Kt2wqjcIDdc7wowHvOclFaZPbPDDDtIdWpnKfUZA2H
y5GDvrnK7oZkq0mMAZ1d3lNLWnpOrwXOowWcNaF8vhNrx8/2ESDGHAjElXlqF6Un
CkAA4K/QPKwBL6c2VgIZZ8lUbTYhaB5nD/M+Qq/qeVGZGiBMHu2fCNYmWeMt12vb
lIrEOrMTzkxpON+1dm4DcDcOqaAHVwCVqIhaIcyeDHVV4zMOkbZMtcDVXP19Eh2L
bQ3oO0WWkPWjo2eOjXR5K/kSq6YkZ4p4Nh3+2qkxKba0woosvVCUbo+rN/oVpW2Z
r+Hi6QeUpRKtFgwrE62nP/FY9yBezzPWEHTGLxZp7Ab9Fy2LjdA8ixtLmcCFPDeI
ROhSdP6xdZLEsOLtN76A2DuLvGX1lZ4a8IJ2a2LpR9OHhnGsRTlkuGEcHejy+Vkc
piCzWzQzZlXKR7D95xaEulvMp4fq62wwTG8tVY9eAEpygAUlN7ctWVz6EtyYh8IR
uRrN1769OdAzhipxFHWwVlHRduD3BsAvOdNGWASaER15pafnD6PXgdCBRRv/COdh
EqDiZCrblANSA/d9Gi4Mo/dzs/aaHTP7fpUrtFgAIfmJCroG9a7LxtjoIKYeExrK
CfFeWg142q9cf4n1C6y0YtUiW5XPOl07zDgnrdMI+fFMMixrr2LcWHZvGajijikj
Hi7MRKbfw1GEdg876/RIBv/pw7tOFcQErSP/I96MVYt2crueheJt1F6VFwFyhI9J
OQj+ELpduBOOBNZ2EHts/GqZZOlGI7cW9PHZz5mNiLjExSubh+woKUZyssrTsUh6
+wEtktPRQCXjdA8Mm6bCzLilba57xhSO2tj3LH5hCsXA1mJPFHwkiSxqgsgj2d4p
xOsGEJICAm37Eb0xZCOYuZMujdlcGOUj9lKus761Pm5Nzyi7fkdMIaHajApoW9zi
x/9kVvrLisjeKCPVo3XyvIPJ4PVvVJWvFIPdBjmkWKH7Jwwhm0GGkaLpDb4aqOON
zN1JE9V2gfoo9/Z6A9xqSVMl9nL4W5qIiqK601uHSJ/0c+czfWRagjaus4w1JNdY
gA/UT8EFBjrwOR3GCG4ZATsIA62OSbP1EhCSVSJdrBMNKEB1udddDGw0BE+Q4bAQ
A4HgIwJvR+7qEs23GHFF+sXXhQPn6mgMmn0DVTQubtyaD/9Tk63qRWwY684ko1g/
WtDWew37CaabeJNEXLwaz67AOlbOJGmwJ1F4VCi2+aacpRiP3POfTV64xwD24CE0
C/uOZS4iwsDMQXRLsczFbLiEaEKz1GU0Rwqn9/qZ3MUKip6bwNY1ZrJVBURBLHDi
Fcdz4UDuDGIiNWKfvIdAPoTplpmFUAZhmYZHFj0BCA6SWOucdUfNpieJV5MZLoCd
SB058Ims7kEaH7D8WMHbETeSpnvvhDxSMgKod99HynrVCOeyZTKMofBrVez76m/T
bSLN707Dgdt01OEHjCPLxS1SEMdfm26TIz8r9ykwWftvHGxjkjc8Ih+NfnRbNKsB
EPac+eqM6VLbl9qGqObVSF9syrqHPVPjgXTw/a4YLo2puO494yChmdWOXphyGKLy
Kq30UsU3d2mv9JV3AjmVdvo9PKwyW8Pnkg9jAx9TgbccHzIcJyv7VvtAG+av7/eu
qsfA6TMGGcFwdF7NQKoeZxyrV9qqTINW6HN/Hf6CPsZzGT1nxZTWKD2QhKGjTsuf
0Jb8yTwVfF4667CTNnknYDMpNVgWCbrpOYsod1svyPQFnneWGx0usxhOi5pOFG4H
gKGwu4FYMvgyk+BdGX+9yMnGITKC3taxvr5L+6afRMzg1O2yvds9cMJmShr1T0zp
9m9k7PdyTtgqAFHu7lDXhcMjknRIDF+non3hcOeiqh37yT5AplStMmzuysq76qiG
qt9ScXO9sAPhQaS64vxqWrs6JxsIu4TJ7GO4P3uD+WEMWSNl/I+3qC1CkrQnJTg7
PF5fuMIA7G7eLLi4KSEGuYtah94nKtATXEr6FIAsr+MtDcro2HGluUvMA0KAsAI9
Sfoji33xWDJlI9zePkCWUUT1dyeojsKdfRVeR8KDBceYdxLkyGYbR2yHwqGFaUbM
itZMGbjfyo8OiHNIkbCzCOU8RjcAixHiblGd72/4XxFHkZuNfFxoL+zPd2wnvd98
WX1dnXGhF3defgmbVXf2pWPik72ryo1uLRWl8wwZJrrhxB51XwjCYL0woTpOjNEV
ZzD/G5/Js5Vj0Wz5YJ3CSCl94r/bBudj80vQt9XZ/7ixm7/8iX/hrv67sWH4Oiwf
rVemQjSCLTZowUokZvOf0GOeTX9UNPIXDkHI+KMJu6j6ItK5/C4uGM3AvVw16kxZ
vZAOuKiVfDq57bIHUp4Y9cuSr08iaj3klFnQdUYR9mrR3SRwCYRm4B24FD5IwPLg
Jwh8P+MN3CPcnO0i9N2F60amWwy10GuCqvD94rFyeRQ0eqxPhAVILWJGLnPFsko5
EJcPpZ4ad9pcWj/S17SvbLbm1UBwkyZL8fQH1h4s+wYLH/Y/91J1lBRGs38Nqqtb
s1RIXvq7DaeiBg409ZirpY707hvjSgzXaFoHvrXNbsPuLBCIm2vYx/jJ2zmfk2Ho
myl81QIsbbYfZFMFC6QTBYqZG2bAagUrgNaVRJmc4/VNSxwC5MCLmR9iEGPksmK/
bduw1/P45FJw9ONEHox+9qdP/pLc5Q251jtzULF61IWemjnHuqCqBWBIA2lXPCr+
DouuEWirSJA4IneYtM66LdCH6u+ZU4lHmcEudM6AY0RWwPetMMQXTH1zmixbmh/j
qcboQPMlKOSeQxmFo6ZzWEgoXHR1MNxnuwv1OWEq1rlu3gPvpAa5hFfRaKo0PupT
folB5YmtSlf72tbJ/dS4qpHTWwDZnNt3bM9bH56Bnqhi0LXWxInP3tMogZycKs7T
x6mLPA+vYQEn4/zCYMJ29rOn1C7Dw7162XlxD7Q60GIANqyzPemkUpodF7UnjAbY
u9BfI/ziTxwYyJgfWYTQkDYXO5Mj2KEuMQtauUTr6t+nJOO3HmExkucJjHYvUX+p
140lrNPDJPSB30a51mY9z+9Kyi1s6CaNE7Ji+xdESe96fmlVx4pyhzBkvFJ0nbPv
dUiJksctu0rVPUA85n0wmzFr8GZTwoJpGH1Zo4jHjNzWmL9Ns5dlNshSTXPXdf56
U9xOXRWVe6k/oCZuGD3qQVF1TxKJbJHuD5TRN4bvIVicHdGwsLexzWIpaJ1XpSn1
MPAzfTiUHW3xlUW42mn1Y3+GTxPM8Z4jyFp9/mC74vEOHzQH0pj0pOqshkMmXj5t
BrscVlHoIRSKfnJ0o+OhibjonJwinM0qYqSTDi4yjLHn3/OaHcjVBT14ansVyVGj
bwQPxZp6iu0JAgvyVwIwnQLYpX0RscQBPfZxMCMKvkPFAFT2dQqHETHgRiyVYga3
8UkSgr0VV9hO+DXykWfL8V2sCBgIyDqKoMCXhNLHXqwN0gef4rj5At3G5ho8vlHQ
diX/0IoHsBkYw3cGd+RMWBnBUnXe/lszvVtYvTgj/Ae/iOa5aMboBD/3Xg+h2ZWL
D8lDjttSWN5iUdvrvM9Zo+A5F2g0eXPa/NHk/pqFRbVG4ygHBkYZeIFCiAWX0edm
a5YDTCNskXzhEcTQbW/PTNjMFdxpdsC1+BacaYMD1bOElSOBu4+ek/qhG9j7kUc0
ZvVpl5fGxN+fHVbrJdj/lk+moW/UZcXUoonAQQmohTcV/VBeu5xIhibUhy7EWgry
6CiiMFDXiuaRc5lr+030IhGWoVOWOJmEHzIOZr5LKU2z2wNkrQT6j73UEqZVW/Qu
WPj2EhntFQvineMNAZK5WZbBma5lhEPfNATXnVZql/DuWt+I6iyon02DnSo1u77m
zXDtr7JE2Of80tIeriOSHOY0hAks4svsBd8MMKY2eIHLGvDxRnpiF07RMiAxAl7R
dSBG2mnqaKCs4RkdI9PVEVUGvP7CCxllUZVok00PASGZYYHj2OHcYwkuFE6FxWs4
4+G99zCsGkikuN7Ghxredr+9JdMreiuJc3dCYRm0Fr0Rz499hH/bF8LdAruHfv2u
CJhh9Skue5Si9eKh8RzqKEbFIkK7pPVYG/GdoQZ8GlWzwYIwMD4PQE4s2shrtlaF
UEAEoxw+QtRKOMQidsRLtU8jofw09zzZO4pBSDDf07bywjIzM0ZscApnxb4ovZpo
1AwTcHngBGdXPNjPdeVf5fDOMrnL9NznfP9UxHvbuP5ZMfHEVi4myZdpBuf/5k9P
NxMxW1tKu25iwg6ZPbVCwacK381fHuBgcQpqcWxFHWCEP+pNMUhalFLb54zmnPrD
S1C917YwDeoNV/OsS2Xt33vkRGbYx/CQwr6Z3Z0raTMPexGIwpRjT4DNOKEmfFBo
Yild8FtfeEqFjbdS/ec6r7MyQr5stqfSgrRIVVDgNPS2WyIsK0qunBMUPObbLfmY
iNVhpcKbdPlZVqKZ1ruuFUq+9ridztndtMHQwOhMpbuLnOPhkKzRe7LnVeDHd78K
d0Q/5YJAp04DhO4WwyzH5UObcr3tQZI59PG/+JjAtVPu8+NL35ZMXCPmnVl1AKvN
5X1k04yR+emdGIHpmORRDP9T2kqDqDLcs5lqZm2GoxiXbrTJiOBtUOW/c6MvWJQm
k5RaJWKKWTIvKW1wjgap+cpHvnrqggb2SrntctZ/pWKJqA4+8TJCj9hUDDI7icoT
yWr9eRAW/A7G07dBBACeLYl5Qnvwoo5j4Ds+dh4Iv7zdtKbEC4iUbP4JKLb4JLye
kylv5wMH0V69BGDHcPHI5UfOrtSIFrOH1u6bsCu/6fwOeIU/I1uuGAz82O0j81ox
AnkfKVR0vgycbK9hxBptFvuH+7zZAdtlphJ/xA3W+1OxKTgChOpQ1JY9IbeWVdSg
V14edmNNjlRBuTEU/YxLPz+cUTacDM5ThOsDod5VuGysdv7JIpSJnqlE09z6UaZ/
xv2QpCrMAIkJZbfbk+fKRQjA6QpI7DVPgJrWTOMN969v5oyQ/AegpAiiiCJ6OXj6
TaYY3Zk+1iazxo0wPsH3zyccN82wJ9C5+raTlrCeAI2AEqvUfixsK3NZjMS2KhN5
eZMr+UXdicbS6AipjE6TqZubN4gZhBNaaab4jGvBLcDbTEwQCRvWzNi/Qt5X5e+3
W+hSIN+2QZQFmkgXKpuJ4tzGvM7jh9j3YahOU4m7zTXkULFgbin4iax0m7I1TvjJ
apSmI1VspG36MuJcdY7BVLlHH9KDYeEcjy6YaavCNGdFAB/rMyoNkoyW/gZ97+S0
g+YhTG0RaV0gL0KAIkGnlPxfxGuXX5vD9R7iq2n9zT/TOUSBom3P0ugRNuYSerYG
nsaQSRGT5TxZ49MFruDLypOObgEmdvbpdWbq4PP8iEV+OdsnsvLHCTVZuW181i6x
W5xDSxuyMErYR4ohgPjYmvPckv8gaxL9bU8h1p+W1ms86pFk9sttozLI0K6ihsmz
jdLB1jTS1ho9zYGU/kGjKhjPqZNjcUb0cKcHuS4U8tzDk9mx2xAc1bfxrQ4XgVZ5
6nKNmHh1lH98DRJFe/LcYcjBfaqWev1MLvDHb9tGYrwKyrTw3k6B8rChagrfl9fF
8O/lmM0pQPBn0NDRPp1jv3KctmxL21ilkN+NdkJG2I0fs9AcRSHqqH6fk9BnxIxS
RQ6nF+x+S3lTpxfiND8qJx82LOKaUd10M2uHvvMeoEsmjPS2Db+OcS0wULakXRPc
sngTF5eM6QCcQ1qDxKTg988tz6lNJ4h/5vKRUR6bkm+cvm5rqud5nt+s6Omc9zDg
x5VmvE8q34iwr4UOzqMucAaHTjyUOpiFzwK5lGoMXG+SlEDjFMUTe6TVLTlDsah5
8rPzQQV2Ny5Tqwc2n0xFxlc4jIO8Mlxs0DfmFTRFstX6L4hoEPG9CE3ZpkJF5bbB
jwXv+Nup3SeDvFMuMT3ePhvODTyvewikxLR88PxPSsnQDhP4ll8v2sDsMhUsPjX+
dRZcrasIUmoGG/q45+kNenqfqM3vJzqIeVWslxZVk6kUk4VLjLYsfHtKy9nDomHM
Ku9j/Hi6emuDExdg2kvWppqP/pCDa1EDpQLHGH5o9NRQFP1kwcbLByFKig3UCjOS
xqj/Tc8XYloF5VhbNIWmhv+5dSXm6LD56Y5189hI4ahbh4X3TcwQPg5mieV/Hrx9
03ubm20VpwgBS0Ad1xW7RHVmsQokRUubvwpSmxO/ezgXsJ9D/jVYjumRpo7K3m+f
eUUqxJFvUiwBybLecG+5El8BdtS+KoC68gN2aMCXhpexIKGOgwEefu3LEJlx7KHA
v43S3OjM3XjYdFnXzZfLe8SzFg1eue4WkjBDJCYDiUoiFMmYge0xkIboNsrFbx8i
mB++nnToickLLYpK8XAy4U2W0PVzYOFwcx71dGLStjVUM4XL1WW8SkQqjF0YBbuH
zjEtRhNYPR0rxjGC91KP1rm/e5BcpLfUNB2bdZ7VtEGh5koYIUPneBvA3vk9Fc5S
q05U8GLHLBMvZrDzrV19ZviINYSutKZn5iLzoBgGcx55rwSW4P+L0x6kpz2p1Ovn
ueeo9HOPo+Q+JG1qul0Vb5/dMkaqFPFDUcZY/jyhmUss2HfXTVkdYMpzIGP8egjZ
tUph9ZIy614ATctyw+JgPnD1wJBWa+5wDcc/PMFNXipLyqsOoX3Mjy/MRI5ije1K
O19gVoDtVk2IPETAK0wOX/7oEdmsE7TeiQIrdd2Nk+Ps0c5N09Sptx8253mQoE7m
DDlxG/zkab8CiZoec6it/1UNXk8yyjrm8R9pn8BN/pre9ayo7Dp4mAFl60yN83Mc
GwsQVFHhvdTK5u/p/Bl9YrEcknH/p78c4n+tbHHxDoj2k9SNzAbcVpyavo9jTgsF
um20sSflQ3a4i/QLgcS0hm0MdATVMwMDm2MtXzqtvd40UTTwsd3fGQeKbaL8v5DW
on1dC8oX4Vv6PUykwOOJX3/rNcSJ7569WCNMj0tespMHM7WMgIb76eyCb7QCXfFs
bcBy4UgHjjDcJwlRcGk/jCu2eUiPrrIJQyDMiXee7Aj2vzlo1QEMPDF85gO2e8uz
9QzE2IKahBb5RGdC8pkCrujRmkgxIdSEIXo0VkXJJ3BjNL+mlyxArizCWs/SXHXC
ktOPfqHMWYgr6ag63UoZO7I9we76CZLL4ZG8057BSAzzfR0sye0MQDDl1XVmHP5Q
w26rdPyRfCjzAVZ0TMYeEM/6ZKU0hGFvxRdIn83tB+Tv+uAo6v/bxyzAyWQ+07nW
Vuw/METCWBWEfVIJOnqPPqWV38DbNxDUFIjyjRFDCaH+598GeoaMwBHvCyudm1iL
cKsy5xo1+sG8dy8AsrWDZJRr6Qi8c4I0hjQBTBZV6X7h8FUDHmqSIyqYQb9R6qtB
r7cs8e2CpEnonds2exdYSpachXS9rFQBlsTZcwgiDMLDJgqSkuEIkmVen7eqx1e3
pu3Xny7y3V6fhcZ8UPBI3kZbwxcaIkCnu9NAMXSBw8r56r+AsYX7bNerx1qIoPke
muugJqtiotGMmB6LNIQwf6BNf4wboDqoY7q4P/NN2JFWCdmNjQPSnJd1O+HA/gjS
Wepc7m3rJn95f57SwiZfVOyQ5SqYe4sPo1fDSO9KV7wfnu1XSsmTne0s909STUPk
cYms8+4PG0xfIpCwa2ghmHbtPrxdUWeW+s+8PqzCuG43mb2dhYIKG9BeC7Z+n3pm
qx1Kv7kz6/CxQlbfstsRYYLrrgGy8ke+mSevXcIejIYjkZXfMUFyctOr8NBYU9Cq
eR8VqmzYl6RZY9gXp9OZ5gzTUG21XkltvKxoL/HKdVAT1d+qtZBLsrzqbIHnFm9X
ljuZkk3/4kEhi8V16WfnXAdRJV9KoqavxCO/7fgS6AFdG1DWaeO3qI+aSmC7EQTZ
ehFskbZHrNrNq1JrmVwaRxNwsNTHpNKjJl+IAWXeeX6snQQ2tte9GrgDq3avPDj7
RY+Cmkg4TDmfYk68j3LttL6Rj+yvz2mWVV9ujszPKBrTh/C047mz4Hwltk3BNTrL
FvjnkxooeB5iBM5YmsRHVNByBPCY7D1JLiEqvPM1Rvee07brLFIUP6+0idyXIIOt
aogxusgBl5P1G0M1uWbRSAAFbnc+T4E1Sr98LT52uir7UEFmYhx20ZhASnalAf0f
MneU39dIqoHH5taeowjL72TJeRRU84fTufg8VRgKpJLc3/vym0MsXnixcF0md6ey
kmN5aZ41+XJINqW2pvrmwEFsJMU9ztK37bNdUT0zkH9I++UgQYERwC8S9mBfM/vK
ZF1ejzwoFbGGTU4VB8R0kfEURWbRMnKYvb1IuIMnMx18mEt5jtCC36+J0bdQHzsk
9A1cUNjKQ3XayFArzqq7JylqTn8mId6Pwdn69iMV9glRmN8QgoHwm7kKoBRI2jOF
1/byRMm2bSjmYU6gnNl51wYhSd0mDP1LvWhAvnH9NtYziChWWqkX3jT+S25EN3T+
Xl0StHhMrneKhyPERGP32aGPogI4CTvs8Fyj+vvh1plcoGLSPc6bET9MuTGEq1/q
IIW+nm8fBDUY9YpdkVnDC9wBEuq8KPOSXCeTur5qYHlLP+DTJ0z3oo6Ux/YIlmXT
5MvC6T3bPP+kmaMlzhCBgFYtdRt0pMrVqQtcvr4QHjqnXGEl9dRm54Rr1yZUBOHX
keofv2q5ru01wlA22aLF9d89/ZJKzCg07KDCwTztZHOF3VKngTRqKwkZZ8wSoXpa
f5jNRpZcp9Fv7q8HQ6/QEnlfK9p+NIS5Z+AjdBspyhpemmD7DwOsSURtLQmyn41x
v62GVeY7rUfhci5J3zC6Ks30DriipkA9uoULrJGApBTYT76B9sVjwyjqiNvu+tMM
DBm6alc69AOvt06LgJ31tNqIQfcb3yGFFKxLCN4csuz0dfcIebwoOyH0pqg/fZr5
v5c3oMbOwpQie0NV1qDyfZCZuWy4pmEpwbuB7Pmcmc4s5x5I1/WSfnksF9sG7tnZ
g/sgUqGID4Okzm60oOAK060AuCf8k+e5TVHK6D8JhapBPJYmqsHeIhkOFm1Oaitp
h6bEYOME8ozD1POeb93PyVM866EVpLWV6K39ZHP0nyOmAMqnxOpNlmRTkzoceY5h
oM4kLNvkwwQqXQTOg5W4Tw98HAqXh+28TvEaMPzhMfBI8pzvhRLqAw0zYbMya6Y1
kyrPYpTX1GKFhEUFhajvhHNGMQYPX8JArwKEHOmE2XWp+DVBXmQGHyCHDtgmYnrt
Nf9rVehR9JN5GHgCMp/tnQ4nLSo+7n74zOiJ3vSYQ/A4Gmhiaw6+cc79/AxiwoPO
D8qkFQMOI9zq8rsMBj3RZwXvjDbRvou5PGP+zur/fQKgljgHYWaBRqHTL0xjBCt0
AZiEMrOQ8tzvreziOEHeZD/yCBiUlLscp6eU3C34qyBeo1giF49gHZaOMdu6wsA3
WTscj1tOdg82tQVIa/86jCnPOm4oCJlVfo9pnFrJOBw1mFICLheKAsf87dcQflDT
q4h7r1OZE2DaB25fEeErPdJyvrR97grqLg+zgAh3lkR+r1urNz/NpotWS9pwOJ+y
9B0jLvkhzrzTvuG2Ggw+bvYCc8GUXyEwApEpNYNgqpdk4/DgCxPhcJxRoKD7GHXX
ZfRBejrO4my0vlF/bvayWLwncVTjrFpF0oVa3uXeySp83f1op658ozwK/rHPbLMG
+GIE2d6KP7i8qMFsPm/oLL79jOJjfm3jfGtY8MTbzTLuuufonOhwkQL/qwg44OZ+
vn0UhER6WVNeIKFXJIditi7+eLLE6xUCLEWgWmuyHCEevTZmN2hrVVtg4rG0LP/x
luu5t3LMIMB8tOFL886LOyDimUi9a5cwq+8wvhcsd4apZkcM+0ooczLRr3NjYlx4
bTMjvsNb6wDBU+SqrklxHOvKu072zPpIdLy5y0eJH3r/RWHEmFjPLgzCWndnLxFD
spGulXqEq5nKJ4zsIMVc5x6HdDsGC4EvpKTkzHe7ReQTHJgmrj7S+BXSYpqHV6pH
gZczSUApQ2P8nhu1p+kG6fgFn8LGvuNOCzRuYay4DvOM1w2knUZhso4i28VxJeKg
A7F6QtvoFB5FRVKoja/G4cZk+MMuzLjEEDwiqere1x+RtMNp81fO34fPFv0F8PFI
OaUHi42eaSAe17ZhA5wwv9dup1X0FWY9vcVkVkWcapqn+ulJ8bDHVi3hMI2zUtzP
dqyUCxS/G+k+t2QOoFq5g5eTrGTGlY0iK0FX5o6o0ZqUBkSyZHC6NGKty0RfIhzc
EtVstv+aHSvj+pIz0BRPL2MAoOqA1MMYduuepEdGsf83K6YxAagKh3Dn/I/bxS8j
UkAnU30D/a/ktAsxXsSR2ruJQ0Zp09OwUdR/wd2dVQmppfbFxfZWN0QNCP+zD3O1
ZfEuzReXz3omn+EYBlcypNzxLWEaLg8V4oYlrx/aKo1jabGOLfDM5VScczJC2dkn
aCl7oHdXT/0xEogxxP5G5MM/T8VPgk8yeyZK4j71Ljn2R4Myarzs861JQtESjHnn
v2XQBzCy3ZmWNTqLMP5+cSrHpouNk1kgAKpszGjzukeYbOnEPHENWc+/4W3ey7AQ
nHzSvSjkysYWllcrRVv85BeIkoZl9enMz1j5fxmp2r4Yz0OMPrGCHht14o8onsSo
MPkxs3Dwc8Zb4q4LvjMSiv4WbFytPW7rnmU4uZFh9AGGA2YOFk9NH/X3lomaOhEI
17D3c0zvYnh51R6EGpHMinxpNxIeLLPJoCodbCBFEzh7KQBd8P/qCTMHGafsdDC/
kfrSIkp0t2GjqYg67A4vQzEfAOsdrrWu0YJ2Itv4EwxFmOdZEVQ0WJJIYNUbMQHO
8DGyKHCNkeYRnrakiAukOsz7aQF6CjPsJwQr5fqBClcxPlqi3UMLDAHIIRvFI3gA
1Aru115QwjPssyljZAJuvRCUwZT7pDNbbjX7PaaNxdHjGV5Mgceo8E4UmRWydFWE
hdTdmezukV4TorG72YqvE6v5LKFACN1WPO6GadDn51TuvQA74AIHQdPLyAxZzovE
nZ6Legsn6ncoygFcm7efTYOb9FZWAvh5FJslCrUFg6nL9QNAgbBWNZQyAQqFMotS
ZWdjSkC2zd1e7KfPig1qXdSKdvk0kRR+8u0rB/XzcKcvUV+ey8vt0807K4ZbBf+e
m5EfxcnV0pCNPjWBl6ImrmZYdrr0e4y7cl+GBWw4zsyOHzxV6FObSf0KqOwYx6Dx
i9Vcpf3GXtZS0KRa3CxWetoTQWUHQ/LqUuFFU0TQbGQzvS1Nbk0426/zPE0dDGNA
+eAR7HZLWdTbdoDdymVOmIg1LZV+OCF5dww76UoVPP/CWleOpuPxJ4xA427V1OV5
E/KlZwvMiWAzZHMSJVS3sKzE6Lit8rP4C7uW78zyx7tK0cEmI8/RPyOVXxIDg1Rr
ev5Lmx2rRX9j14sO2w9wmILmdUbr6KIx4HKcF8MQOhb/I0duvG5/1RJH9spXR4u8
adN4nyqqmPfefkv33GUqXuhyBGKJQJrul14lChKPWDUFEui/PL8rKmLk5SQfPEWx
a1MWK5zDQYr3R8GTi6mNPwFM18Y1zJEYt7+Ekv36Py0jft2J/aSk1tlg9sKT7PSl
mwH3fugP+KKrwsjWwMBB9P4ok6I9jzo++w12WiX0ncLVHzP9tIbEjRjEdFDj0kii
Kax8AQyiM+iDsTQE7RAmEHPI3Su59auAtIAEAfe3J0sRd85UcbDduwtcaOrb/h1f
uyTjSPhs3dfgE11pWzicHf2sga0hBqY+6Y4XwfPWZLCSPY4v7FJrUAtdXqPMyJR7
krfHEIUlVXREegw0rNcEFXreF9DNTOz5ohC+/NaW8pUrHSUYXhg5fF4FSjc3jscN
ISWprYO0gDEzbXGB7zUQM9uLVk2wtPB2Wf7n/1ZFqrRvZaUNVtyXTp/preDVuH9U
ch9FFIHF19VaZOQhlc6adz+8+X+eGxF5hBr4aO8j+3FkrQJtRLJTIHD+sRr530uE
xPtNA2mr46yoL9JwNE93we3XDuPJZ3tGTO/LbQTXomFD/aevcjZY3g3W/0SxABeG
savDJsxRc6wsJpwWK4+SP08o3VsSabPjiiWWvdZzY9I0fecjmWNl0pbLZ0AI7ffI
/UU+yzGi9Vtl6qvAiUHFe50TGOJQu+vRGrpLwG7YwflzDiD05b1O4ZNS8ovE53Pb
WmL7AgBYA3OgDXEoyHKp1CvKQwr3xxHOILPsl0wEm9Azw02B8DzXE6aUjY3VbItR
ztJlJl4N/k66WxJfWP7lZoCC1EQkUY4ZsyrGW2VEi4lWAhE4XL10XG/H8FXrreo7
sQCuI7AT2PBvz69cQW8Tzyt1gXOL84wL0LalOMVilYshYqC1bnWaW3Lnumm5KNjn
uTPwpEZnignXA2rwX1DK+S3vBij1kmaABSDL2wGefZv60zxTKf1RogeXZR9DRcIH
SdzhAZ58Vh/9v8ANzx/zIknKEn2joT+9RhVRP19hZ5Tbj7FnvGbBdcR+jrPUuw1C
GRWnIEx2uLn3sSrwr+uXrtWrwXhRJWLB1IHJIJMqBFk0sdH9RHWkP4lHzb1bahCd
W09uxs4BIBZjFtsxxX7yTqPjpus8pFTcbEJXEBf8Y2PqRPY76iKBCm0jga4CSibv
fCRdOMRNSJ71oXrmccd7ExLZBohPrQbwuQsYFXXYM3tXt8n6tLDgF2/QmiYMpc4u
KBpULR5dODhP5gdN1rD/twBybSbeZNUPtOUNq/ik9CNPQXD8v9G0IOexqT4JZf+T
83XEcpVxFyc/53q5snPJFfFfgRc05uTgjjtklxboGgQhrYO4e2c/dVQHlFNgU1Vn
FFTcFgRn05G8wOE4BjIIZ0cKvIcZk0KboxHhyuWhcc7uXIiYo6x3a8ZvN35RENWH
58MNHP+g7hmQGjIqTTAnmu9uuDgbkqxJ8vjuBTZcrZZCCpXDKwLezGSspKzoRQxM
Bo2QmKtW8MfH5hpkb75pixLwnBPsnf7mJQ994LBf435DzGLhEO0719DhbhbfWDcu
IUv1HISrkF+N03Ixj44Piu0uy5NB9jhhCblN1o/xJo75LnFGkuCSbYMyzeRsQY+m
yhI22jR0ITn5aR3itY4SeJlIEq7pkOGpMlUcp1xoNPa7zHi8IyTcKnWkEg2j55ht
67nV7dzjRRWDujN18j6FAyD2q7MB4q1PxVAkLY0qX9VdlxRYrrmdXmS8oOnZXOQX
RkPez8B+ybbt906g9PBuhU7Wy8G9s0gLHGzTXVFHLFNCuspVX7+5H0zWQXsd8SCH
yZZ4qLbFg9kWgMlpFVK8vqpP8pEAT6YLwSzgRUa5IUSREvQIOvNSOlKIrDDXAyzl
7kUhmAZwaESPZyDIMW/KHb63EqNAYZLV5w/9YPPPtHj3AXBL8qWGnUX74bXdZIrV
lntIBa6JAcvO+oz/+ikNpWj5rvLFHU35ggIN/eEgehfsC5aELZ3kShH2MUlJmPsB
TmPrTvcMprohMGSIC0VafuZ/rxjnCJBFHwDLauh3Wtr7vCjRzYwXe8AlIzdkj2rI
F0dMR3bETAY5oXRNVyrR0eG2ngL8Kp3Ey8bP6S378cRtuw04jguMQ4UbB737CbUK
dZmnRd9+0srJdVKqi15OBWrbzGQdfcagWwoIMtrdzkefSkOQCvswMtW1NsPYqRqb
fHSa1iWH3XIN8p9YCY0ifNnSVrlig66SkEFCIUH1fGI2RXlEPodjfXuT8mnczikr
DtoA5HgVQc2TVHGJ2c4XNgBBLVi/bOrPEDlQ56L2HMejlOm6jrVSj1AcCsqZe3Vt
x98gFgKhQBZXGTq/t4sGoL1INPwL+v5JPLunn+zQZzCf5O57uwdo9b5TUBdKM+eh
MxuIYUrvnDya07ySeiXHa3MOxSP/Q3QrtnM3Hoe/w3f/QVG4YDYS+/AlF7F7KZ7v
95gSaQ9w0V9Ihz7pifZesb9+4Z0zfyFko+wvGMlplQ7Z678QCdIJZdF/x+WilX2P
QBLNNMjcF6xF5L6x0gNXPfFRhihVIHLwnHwhiXpcrNZI5k4PfhzFYfZaw3FFLPeF
Udbxel9Aw2FQkc7a6oa4V/UIF+huey1xr0Om2w43o6SiGH0+4QHcUYGihFQkcMIv
cxD0xpkQgjQZFqWBZwKs2Vny14e+iu8mwBN/knnJyLgCIJr4AgNWKnqKyXtwOgxw
+iErEv/m1Rpcc42TKRfgkUVXMDyREVqCq5fplD0BpBryDtVzHcaWIFMP8Oy7298O
+1bGK2JGvBI2HjVtJwjpy4NFqyD0jwo5xd/yOCnByleAJMEArJymakgdi7n2yscs
ee9J3EbKtJSMqkNMfdymXseXRPwfawKqbd0bFYS18X/a/GA4S8Ux3Cx/4QL5LbWY
sOUeg4++IAlJ+DFMUhyv4LI4NltooeslwIUDaITVZCPLqSotneb932Tft5DCkqN3
thH3mfaiZPPiFLwtnhiv7raAHV3qVNoHbF/Ne7uOvxZbl05MN0OW38cizir/XuNs
2EcKRSLOR0Tq5zkk8oEbcuY9eREG7/5hY/4GfSZ9LlVeAD8qMYRmEzQ9UQs/k4Cd
2O5wdCjGrB42D3sOYyYo6072lS0gPEnkcxC6DdH5i8n6i8j0cKlA9zGTdvjar3xN
p+b3K9vM1N8Q7LG8WwYH2zChI0wnFnlkM1K6TXpt9wcjoLKmq7sDT6xgwfK/kDd7
urlAT3RD+flLa8vBRTLdPs02q2/14UoMW9JghR4lRhcp3DInoqJ2a+Lq2K4U2X5s
izz6bABTQLVZ20RqK4e5EkUpIamG3DaF+GR9nkR+7xq7cPslZur5q+HwCMfd6cGH
dUvTGNoqTnLQ/I+jexkdhQ9g5zE9ifU68aKs3JribIe6OnQ3iV24vPZUn20+Wdtc
sbmOHbXfGZRe+ScxGBSOaJTPEzxO+81a8NvfjBB3k+JuhracHEiN4jZ/DudwA8hf
fHg1wzb21w8MwnzoPOccr9x/Exyfemef1Z3IIq0CS8LIP+Sjw09OTbmOJuaTBWVs
REFpkU9XsV1X26wuPtL/Cyn5dODcU5Rr1JB9X67N3538OihczRiO5P8R59oY97ro
w2wjYUKEKbwY3dCdo5xwG5JmADJm5E5jsDEdK2PqMHxIL+SaiOAz5Bnc/vBgZ06Q
gkYXc4knIDWDCiVyLWtFOrW7ABEf4MMpsgRDLMZ4D7wlchT3tbxJM6s5wmnguIY5
qZo76juQ0lP85kVdNK0ss/b9oH+7RZgc2lYEVzFwK2/803OwHVpKkOqJeIguqGYL
freIqGN/rtfUXf3SJZ11BwAsa4QWygIObUB8QmuNdYNKIx1NlFB5Gx/R/TSKbBxR
QeGR6FYEVKLSDS+rBwXQv0k/6yakY+bAwFMPL0TqI5WwaxII1+z8Wtwmdaw26Ho2
ECFdFvbnx3CHxryKly4bWHPiuQUiAHF5EZME+7ag1FBbC4hd+XOTUyu00MfKV6kM
WgpvDMHxRkIZqE/5YlkM+KZoodGMZ1RHIQ9jg1Ek080Ic5Ej3Wz5O6ETexZ9KqOT
WMuDoEw5K1NpF5q353ftZYjDEGCt8+nNM6IEhU9C0UlGqfujcGmb6XMD8mhgHFMg
1fr+joO5F2fL39idWoPuEhi1W1V7FB4mIQZtoXZEhh7/V4kELgIODGnKeNkpxhvC
cBiyMHsfPjxBNcrnoYkeeXmUm6ghrJTvGh68fRUfLusmxn/QWjfzOKav+hi6CtOA
Z+hjj/VQiWceAVuI1+UouJhffdtk0H57NcDmPgi2wlys78RTKM1Fo+IYcDNowyym
PD3LDVgHwTU+FzXWD59qEQEOf84oAfHrYryZVv8cJqqxNKFAL8y+nWJRcgotslDx
uqx2ZUHey2flfDMNZyHDGKaNjn+FjGpffXmX2XE01gukW1ldHy3tkFpYEynuDRgP
le8k5DKivQ+HQnk+3vXZ0DM/J+imQ/ikpf0ztwcMGedjFkgXNMvkhhOaKoJxnV4e
YLyamySuwlssF5gSd0Bsc+ntCWbwtbasO41XrFxiLnz7s4ccsb1ZV6jVd8kucMMM
eYF451ajL06FaV/Tjsvzf/K8QO3jrRWY0v99bD/Q/5ymZqbERDTnksp3B3Ne7hf1
GzFpkocFPenVo/FcPzh20avp0A4pMIa2UfO9/Zd442I78XAZMDXzUwcOCp/2ibCT
REYzN6+hmLFCUFwppfoHg9Wt/cv+y4st/wEifebO6XSExuDCbsaKEipC0UcaPXr1
MmLnNg0BTy+8zBLR7nHmnzmv2gU+SZvmdPp0c5u/f8N+KSss3y3ICkAZZYKhaDTW
lQXLdYcEi1GnQfTOnMkM+Zz1tmKz1rUmtGG585OeBLV5xVEhwPvgovgiHjqTsggg
gstlgxj/tfJOYrExsb0uw4bK8VLrwvAH/BFBrM5FJxEeF4EzsJPa6lBdLlbElKWu
21qFQtICUzQOL7Db38ctbjNvnpseRJ2xM/V2lVnIcK9JlrXWaN5QkqSEuQtrOvGw
zYYtLEDOUANJTr/ZkyJ31OCQ3pKBM8iFbvuU8bvLJWmwl8IeCOJVDLAmxrpPzT3c
b56LEGoJvqaztVtmR9CZexrW81d1k/wJQsc2KwfW+oUdGbZ00Q9z43b+jOg8jO8c
+Dh1x7dEGgD/y6m15JK1Nzmd3K4JN3L2eBwwPMrgYLv0tWqN6eSzav1pB+kCxHMk
mdedPn8VBhwPU9bHa1R+XL1jU1qqbGOcsJX3p0IuNJrX52GFjqejhPIGe7pZ9zvT
dmbHAFgNLWagoa2H9hv6aUCtMYxs1ON1jhAsL5NPho/SP2yufox1EpeCdlTMCRAT
MwHMU8ETZSrf7XHtGTR8YE+bjPMSieFytqRv9VdTFnMbOWk/KScr61pL3HEqU8Qn
LlnAuQpnJwtirm8V1Ock5DvXUTnOr6cJ5jq59u0nhgP6jedd4qvGTx9nf08GnTgW
KSU8AmwvzZ2/uEXfP9sgFetILf0Qsd3v18Xc1ThQetTUZAv2/mhYl+5qm1tKlFPO
0EQdb9MlA5TTqA5j5n64bLnboG0siJYrrY2p3V/4+Q60O4FPmRSTDjpoQAusvjTm
4LQr365+q8Trh4BmYdgyFAulb/CAle0nkIyKTabn2c7qGTywwCUhU9lKk7xXh2C1
peGhAXJqYV5ATSe3pnYQOuH8yqkDqQNo41xcIufr0gobYs7rji+GIl6uMQQk2/qD
SbAMsUJN3LVE6zczYNPbt4ICqUR7fz8fqYjeDqQxyLIOEZ3V+xp8+JMyPjK6jUWd
QigVZcD8gZwcFRdurbC/EDlLNX///uND6nrxgsIb7HqtRzL53g7uwJeyN343pU0E
B53pYE6k8b2x/sVVHit2rFI7ArAfB8uf/YDPFZt/d+SLDk1QwssK61jG/zz0U+gU
qwlu51pN3xciIzIJhZcugplaWE3+PEVVyLN8/xvo8lhJYT2c9lCcYJN62pCeSJsJ
bjXlzy9hi1j8lrszWZVKbQvZ5VsVexwQhJfVATixTcQhG7XIlH+b3CLbeA/cvbM7
S3Qcbc9sYnnQLXTrVqGhrVxDr2HmPVSIyu0uXD3rvbbVuRSFzC0IGjfZZJXxWQF4
PqqhPwegpYgLRKKFlNMs8Np+iPsTDJEloIBnmJLsoYhMfh19/CH3Dhn2hog1XRby
z9sDzfJlbfQNCvcSuuOFGFpHogYX1WsUfrYjKlw9OSDbAKPj/lbvq6hko7r0xNsa
0ntEBkpY7241YGTMUrwjddXBfBttK71rLgsRcteJMhljNP0P+8zW7PPGNTH2N3LP
6LJJJa+KpMgmenFtIWxxyt1stTX1N0LGvJgoa/fCjklDEyk71XBhZPwP0OAv+aUS
qb07UG1B8b/pc7D1DWBjPM6wclGz287xDbn0QoJZwOFZA+9N6FgoK2JbE9d3RLRM
Wj5+c7WGp+g/TMVHJQsvC/c6PnO5wzM4/KlDvuNkiT6OxLKr8eKyclewHfCy0oI2
ar++0TXX/8Fv/PjY7IjwS32nYliP9XbK2/IMS/WBWtuqFXWPGCTopLSlJkuP93zI
W9IBj+9lHSghF0p0BJdEZY1iy06SNOn2Tz9UAgKI9M2HkYAxcsoJkNYjlmrBi4/a
C5n1PeXzCYekYAc4WWgDb0ssoz0JznFuQkuB8x2FMmlzusy5PabY6ZOENHxMFco6
wlyoo74VC+GVnTzP2jOuyYZJvC7un8b+c7eE6pQ4so5WukGi0ERErqYjEe1yeVVJ
OUY7CzC/q+XcUpmu7wq466LXegkT7B/OXW6k0pEMF6uI+bgklKEoLGWsSbPhUfsT
9ghU4Wic3+WR5VzBRXZkbd4bFFd7C2GdS8I6Ghu59/5pZexk3UQ4Sz/TB2HClM42
dKnTeA9WHBGofuu7fwbxV7POiGA9o+xnDV/OJfvQS17RuJGJ76BPzur8fELiIuiJ
DAf3aNjbWjZ+K+OuyXWDFrt5Imm2NT/U89zkgy1viwOHqYinW6aY6HaqxxNocb29
zkKYUqsBCscVp5A+TvD24n+vymsrYWU4yp9WtHzZlGLHsD3FM+0S8ErPECPwL8d8
i4WsJjCEWW8JqVg2M8uzAeEBe3ZtMeXHH5j4psAvkHWlp5VIzCoAp94KXVWtgPQY
hfGgK3jR9HoFuFUgNBl5juOGsuhFfxtL5a7WbX2SLMgHdIlZkDjCO6U7RhyH8uAo
cEOTmcOggDG4xlkg+ZOpp0d0I2Dm2RtoT/8pZm3GOlFQM0OrNgvxmbr1cPOypGwz
+M2q2juQ25cMtTujW0PZWv3LJvGvDwkFe8bZHIRjCBZhFqQr3buHmw0Jc1DpRGC0
icHf0LRViAlhHi3n7L42D8jjgScskgNkzUFvC4ttSzHwRDho2OZK+Od5umo8TKZf
679bvzjt/pBJwtoV+0ZBwdQGkZDyQqC55oN6QdUlLkZmWpoznk/JRWhO1OqoEb1u
vXI8RTvOG1NLJpW4V29pOK/wMiwHDcFNwZLBIn1NN7Vp1lExyQKRfgx9DxLRst8H
FErCWGr7qxzT+8EhD9eoiiB+QhkkMM12lgHLVllMm59Vt0dfNVeWEmHWlkj0N2kc
3mzzMPkqIKDcDg2pl2gzVXLcgbOathsoWa2R3xmuf+4sJsQiDlKl2PaYgHeluPnS
VPa+54NxU77juhnWkHSHjM+MabwvKAhA9ZUxH2Qfz+kG2ertRLLP835X9j+sglVd
D30cnvnby/wOSaDAPlEfwJ1zrEGHIHSlZTyONRsFAST0YMLM2Kk/RYzjaoXNIh2K
clPkBWPnAdFfp1VioJ/gS/VBokFVzheyOYUMW35mBOrfl4+uvqcozKAKBrI0YdYi
W8jzDmTpilutIBlBa9W9qwLBMcDPgIXpJx0xhr8la2f9Shyn58mbR/6QrdolbsqA
P8t1R7XHNSbFFD1VwdJaVR7XfE8zC61jV/dITRye/Zm/O/Gce1XHtCRfQYnE//HD
T0UogDvwlDmu+vWUpcDCgVvBkWivAt6aunfZ9wyDAcL8qfRBQDP/Ywj0Fo22gWpe
75WRhDZ3h7EwW0Mrp87ENKaCjNUYtqENiaVGyXxUDVq1UrNPnLXvgnR6GFsGFa6X
pPBT3qIXWoikcV/hwiDOVV7zVN9iEPNjFG229JGBMdJgs4olKbxC5+KjFaZgmHZm
LKot7ItP/aHPa94RksCmH6YkMAxKBwWS6X83dv5aqxv68AoZ/m9wGUNnGzRdunm1
Qifid9GKNUjFIXx341TNIAFvOhdBdPPKM3hhLCCuU2l1xkgY6r2nX89yGDi5BZlZ
bVOgrnjDekPyHj+l+cQmbIcdVqFYwwrItZcsTOnMLVLes9OAvZR77U20uqW7V38U
jhV79QaEh/QXVGkcGQrVXKEN9c224evfyrN1E+iWmxuDalTvhWI4xuJRzIJ91B19
v/EDlaO2FpEkX0VX+99NALKUVX4PzdOWnoLF8n4w9zLDlYqYmtEXeIHY0tTpa8aa
4PWReVOkwdcheSiOqp30/AbBjZ6CuM36ZlJewIn9irNqOA6afZ6ycfwUShlkbC5e
vdozSWMUEDgBm11nN4iumx/05DM6YBQW7zFcxTXxdx2mlKIECFSokVyDe1EENBjM
nfka7HD/ofqbfPWpwZcr0ppJKF9xGxZTUUZyCXzkTBtG+w0CdJIyYcil3LaCzgOi
sDfCqLiZjgDDXObfvLO6PwO1WsLGTTxywLcFOI4qBcvfsupjrrHxPi0t/czZWmcs
RWx7o7oa9mumhXD4FP9Sfqq5misTI8Fi6fCDFJQ0wBxXFCU0a6EwFXIh/2BO0EB4
yIEDap8uKtoT6SY7t2Z/VouuVRXmdJOC7Z74FUdFQfqCC07cxuKLF4Q7grwvkOpi
aX+BVoL1qU1xP+NAgwwpIZv1XY2EvvDFl1SS0gtZXmPXNzxBXeVzYiupJrt8QSnF
fexd6MXLEqG00HsmUO8F65LMJR64q0qZ8HicVaQti7c2i474SrYwDbU2qmSxbY3C
8gm/aYrDbox8JxEtbfnAgZlxX08os4a5UY6EaEChT9HQEEJktKgzt15pWNl7BxWc
YCfhQgB1p9d+4ut0vr6qVWDIesMEwnqAKwpxBpRAbxkqfBnaTSMK+ReE3HcYTZMr
UvhrjqfGJLwEQObAY/GdwG8QReGkMd1tEcLeB6LQ9nrckrmTiKpYVnU3046ddTFF
kGfo8JcDMMPboxLjxywx6/v0xmJVchVLcXCDhD8GVgrP8UH9d++VjaYkRKJnUUo7
iwo747fO8wYHMz01KChtCcArfBS3ZO6OvduRfwT6SFJCy4TmG2dgPa48X8D9a8g+
nIxKSk1h8iIwDNgUHO5AOUgy10sQanbDBLkOlEBq758a+XH9+b72U0PjKAkmA0sX
+GGvTsy5Ql3ePkt6bSnADFn7nCsn8eC7RM8tQikwrRJjWcpixZ0NbcWhPxbN9gqz
biA6LBHesfOXtCNyjocAHsZpAnk9RoovSDyf2be4cgN0w6kSwKgTFVR7PEeNA6Tb
r3nIyIp5zvSMix+kiXg+8GnO4Pw651IMo5TiuxgvzQmZ1Ot8uF80JcRxvwtU8KZq
JOxGtxXUs42FoGjCYrBXAp5E68DQP7F9Nh6rKPYuZax/OWQSsloRfIInrHSMGMTW
ciVxlbRFPplscaRQmo+tXabOKqgkvM8DvI4gS5HFC2tP23+GVhi+Ata6kUdfmYNI
2HpB6UwxvfDuY0vqbmkwO+4tOdJC1iO0SVjv2oT6Kzq0PUQS8dz3voDsG7/coVwl
WRd090cqnqTjMCq/5d4CaRvucwEeZ3DbTHizf/Jb7LCRQhe0xstS00jNr+Zm3U5n
EPqosdUKn5Lhey9ANW4vjRyEsTdCRiG0E8UXhvc5qeZy1sZHAiI56eJ6vT2RBaTK
iFK3mybHPe0pnmM2ry9Gna24Ra2QAcJRKfvMBGevdqweBt4Y5BeU7P/49m7tPcgw
JsA5fJnW1jFOAFe47X6Ada8ugmJg8fSAT4Ep5m/BC2FbMFTAn2Xh/uGKKvHHNkTn
eU+iT71CxKFpKts7aaVuY27xaUwYS3CsdJfFPncKsyoTIgZHjk6OEv7nXBQ095H4
osxD61jOqoEXd+XbE7N036oqQQ4b+MyRzbzbOFw9TvIePvu15+HH6yun5BOQoBWH
Mom9R9sXC1S7cy+c6XYOqY/wcIhX726AkD5/LJmp1qxtjV2aG/PYKZAyj1XTwIvy
kOEoXxbraCgYPnxwKnygCvtQEcYYZZYWRPz8bIZhax9cQReQsP4twL/a1hvwVBc4
l6SLPCcgwohjhz3VWzes6n+dXxkYCvr034NLCWB/UBldNa2IiD1eG7d+XaK0CgDV
00e9ZUZG2cgqHIW6joetF51lmT0vCzU/g/8PeCIiU/CQV7LfM7xGKDoaWlMBM9iB
/giOEnGCrq7aqNyKEOhpZNeQteO5qjd/cIXrXV/6wjLUzNnKz3PhHztZcKgslpQT
lsBV9FiCq0VrLJ57NAw3qtgDYYnqogGQB7eAkGIFjPPClDtuhVto/o6zBXBjoPCr
d5ySls9RuroWJlpc0ZHNyDGVJT/83QqnZS/2RPzaqSjekiWVxOgV/diLqvY5DORa
NS2ffehxSeuBVX9fx3uBBfckGqdwxxxHHQgyISKHDE6CBAIRmlYTV+DVjGqR9zpk
iivycnOrZM/+fry+q+swkWNigjgZXNMeDdbNBvZ1HWNf/ndAxdACG2j903Z1lOMg
lw3Qn4CMHgwwHbNmHQaCuonnf6ZMKKG7IsFNsWm//nDmVsHmEnaA44TOS8i/35JT
neZAm+kGWGnyd8kv1x48Et9sz/4A6XDVQeJEzUtgyxjmSskBcC4uWmzAOVRsbYK5
ssIuArFNxvOSUedgmibl+fdqpXYH5MqqwNRBfqY0eZF6c+s6dk5sirTpNeFHxcpC
61MrAIbhg7E1bI5Cmiy/x1ZRTEMKDmb9yORW58HlycwVfXZCF/2JR5pG57t3KIKn
+EA/WVnJpWY6W5ugpmuON/C4SulVQUVXt9MZc4qyqfSrGJc0sq8DP7hgIPrRzziY
tUNxJGpgKaOxI1Egf50Qsn60IO6nVyiemIEvhmPcrymfDYQr2yfFx3bfuGEyOCn2
UodvWI4Ql4LwtOnfWiqff+EFpuHGbi1VYXgTumRCQWEkX6W2OmExtWTqU/zvsBfi
uaHuG7RBMfybXl+DlyuKY+6JLitEkpAQeBseU5hyjba5NntsqpZsI2GYB4eimDzT
KFDFZ85uVxoLFKZsatOy3NaxBU09MYRC/5iyC2UNAFbwPHt76lto2bY8jVMBxAkr
tKHKlReRKHa2SPCJ9q+f2VU7I2uatvau3mRORRQrQPWXw6oSTnkHTAp8779rOAqQ
aOpoZkzzfVuRoCX/0aToEPsb2F5qRK1cG6kpCVL203/xKmlMv8+rNvOEHtB1U6Ka
BpGBLI55wT1Xl2W77CnUIsoJ/tUxStTNzbFoinddTU2cAZhwsyqDEdqnvhBrZRKw
JVUCLEtaQ1/VQnJn62vqfwv+o703sy9HOQBbRNxA0ofUXqi1a1MNNcBICo8TpHvd
Q1thobKmqpc8idy7gCm5qjIJ2WvY5Sq9GeBXz3KZf4QLBnzSvR/QCXKuJKKc+gEZ
UcO95l+roYG/F6TEqDlomOIv4WWWcaWEaOvMCZ1PP3v7zQ4MHN60oX0VOYDPMAAf
JH/8jDyEPXQOMY8bYEaRkxt02GST9mkcsQT7KR0LTR1ZvMrEQ5LOUye+JcuSJ1aU
8uaRavcCwtoefsWtF61RgTQRjhWbxkibe7NCtr3ndfp+xeCo3MPaJprabzGmwghK
g07NKKMDf95ssuytvV0r1XS0ADNJF92fIuellbk5krOtP7oVCeuHXenySvK58rMq
/wB0twycRuyGD9lX3vuqbhkavH9TyqGpDMFKQJ/p8Yg6LJlnLgvKYHcS8mG4q8/m
38rQmbx3m7NTeMkhql3ChFZrSdXzKgdZqe7aDA8SQBNLF/uh6EYkpoTIJw6aM67U
w8fWF39X6Xp8udPZj2La9ZpstuwBKV1FOL4l9mqS66atYGUwFHoy8W+V8Epe6aRd
Ac39kyhzdWrrfKMYXIs6FZS5gSGuQvM0xqcpjUb2YE0Pb2AThcWWXUAiEz1MXU8V
LveKPI+pOBnYdIPOvBcLvS5KrKtLDtljT6MBkSliO9OW+Wo9FDrdMNDi03eV32yJ
TFovsOBltSfgXkdphrluiAagdWBf9d4hAaUVDtPoDNjW257hiELEEh8mXhQZJ/0T
aQVOqQ87yz0XrPiA5TIhaHj9exeLFGgILAKoVWp5uByhfryAgTf5xrH7ww+Fl/ES
SH+z+POeTWWbgNRBtDhr6+kCxDBRChkqmMG+L2xoYMroOnzdCCIF+r68Ts2BeX/L
aqL0ho5ZJnS/chdnH5LqH+DmaSR17LakArdodgne2SqofL1Cgn43CCFCp6jnHnd5
km0G0EOumv2vWjy1r4/Nl1r8s/NeVkiNMeRoxBFwp0ijhbyg3gwYb4F4G4gH5+oI
jE0ZCdAvy9hy0Jnp2rY3vg1gkIPZvIJinFfCBSlKRilHAVATsmKL9HN70hrDppgO
ekZeAjrwSLl8ADlu0WZvONITGU6SycRnU2z9KaAPMl4s+y5+n1GoAXIoKqIj9lir
NqE46OV7paGtjWgA+Y0gLTap5q7hrXPf3PyDtwOvjJqfhWu/4YtauOz450qRFozU
bocdeZKPbnd7y/GQDnp6mnW8THWzKE7tF2fXvfWMRB4mdcdYsmUVtarcybiR0fDe
6AZZ9UUN6uDq9t8O9ZMcNIr1LTtRL8fJVV2cem+hMAhYUVhFijts2Cagjz2kimIm
6BixsWTes2IcUTMx9ebwzRorq1rkpfhu9DId/Xq9pLWg1oAmUQ1Xm1gHSerIGzVu
Exf6Kk/7HJjXeH39LQWCKJUGRrzNYOQQ5RIaYYyUU5/BOIECnHrn28g/5mXKcP4j
OCIaKGOwdA6QeSIAlSk55HiWX9I6zXeJ7FFSDDCp58aPj6qT34hwZK1zedRXBkuS
Zjq4KhPwH+/5LDkWJnUqvvoBuQXf+frPQXJ+pEol30auWSeKGfnyGzxRroQzJGiV
MzGXh+le/px042tDfPTCevpkFbHto947Z9pkVtYdjhGoWR7darE8vCARM0CrM5v0
m5uj6hu0B1iSbWCkJyqQDcaaSO/fjRzIM32nBXQUIGC9IlLQrqG/cWt9bgEs5k0R
6UE+e1hfFjLFAVALSnd2qCL0mnAEbrqD2t4uUfBls2VLdnrey9nNIBtLoJ3+1gUx
FLyi97DUjXDowEiSJA0K/RvYTsxtODFaQFusRXE+FeGC9SmJ3jkwtousclSf5nTU
hMUW22VTjkZUf/XN385Yw4dXeZyRp8BP2N4xpFTog2uYUkX0WhIRi/d/29ECeQyB
jzR3lBzRM+WVXyOOWdcM12Mg+hTN1GvNLJFUfW01h+YQ7nhRCsokc6UmebUIfTku
nA5WAr6hQ+ufXohHfyyOkNW1GyeXuJEH8smAtNo56XnxxGYC9RYK1PNVDtc0eRfe
Jb2FQzwwmjm9eQaUce8igAC7K4/uVaGXwLmbthgJr+y0IkLba3D3s7XiukcYQnJE
8ojuh3A9njytkHdfMHVC1BfcoKJQf+1Vfabkgkm10K2AD6B2yV2LDTieGUzhBUbI
4+36b4AHXaohiGSsZqZgYHWta1G++xu0szapAXTXgrjczq13X866RVHVrpy64RF5
pEDziFAD1qvuFMRCd4Y0Qrg5r1PpWqK6uHErHhmf4ubNXc8giyfAB/G6RlSyceZl
NFM/iaY6sQ2TVbRV+advnUEjLgvbBVo7fsfBN9Jzs3r4mH1crlH/3EH5SsNEvN3e
Oazw/S55/IqdzoSrdWRPw7wz6R7/1H9KXY9ukVzDTXMffzKKr8srV9Mx8guBW5Xc
tx7EttF2tBNF491E0f4mNdoWA0/VsmlxSv72LZYNQUMxpFXsjtOBi91tQkrdC2ke
S4rEKbVQpEoVZMIvjnc/WdA/GATJ6G+NyLqKfGXKZkCVzXGqQJFk/DxE9aPLclR4
zsH/QwPgOmyD6sKjYXYFt2OSpFnTOxR36W+Fk+ZBEnR9xP4wbo9Ut8cX3UkJ2IIs
5egZPl4yO4mZobWoa4zkfCjyd3g/4F5dY5IlruIfyZI6Cqi9Un5YiT4gfpyEYiif
BY62cy9gWh6buCaZ+9hfPlau8ZwcSzNzGuB/DrEfZquT5Cswk4+WrAYYl/WSPsu8
M6rt66Y1gOKmN3ec8tkaYtR1NIJ9+2/E9IIkjuNliP7O5Ry543gl69TKKRwnwKN4
8EcD2qQZrn95vTK9IERJn5XW570uIgC/+0DFkKdl4veL1YjognbQc9ut/5Pn0l5/
UK0VOWV/5kaMZhsNXqZA/9BJJz1kRQoihyryyxiu8jrG/63tZPUR83LGU/psmh4M
7x4OYo2u7Q/2Enb64FXpvCXPvBYiHr69hbSkhazyZ9lsU1JjEtJXM9tPMunpK25S
uhkIZxCO0YtBju+Tj/EyZ7dH72uK5I7NF1Cz5/3HOAr6BUW0sKFIvH6EFL3rnIUQ
0PTLVJ/77ToJ3dvfcs7M/NiAIVV4rTwbnfFkzMcFK7+q3UqpG5bGqX7hwsnAIYdc
sHCbwy+hL1etdCHqpUxUEFK9ETD8RL1zCh0rl7sSDVBkqaR0XaCttxTiNyBCBQOu
Ki3zxj2TD94eRtqqVaGd9L3tY1I+20utf6y5gedHrFyhKc7Z6SV7sXg5IJawYQ1I
VvrfqqW6O3+nXNR74hqLz7sRUQPLp9biAoWT25KJ7EY/lOFT371HPN+zXzsl5c/t
kr+nnRqgbdtDXv8VYsPaC3B/SUcC3aLs44hSJJAbfl4qqk0+M3iP992Fwa+LEbct
spmQENt0QKPnitqPNkaf+9pdwCSxiWdBKNVLXsEamoghITlbnmE8yT8AgQeRYLoi
cNHrTQOz1dH5FWvgV13LoXyD72apoKYGLXcRRvg7/dVAWMLQwNh1suzUciFP0KMe
u45kflNzPGiLBciiftPNVEHztPzkMbh4QWzYgxZf4FPYPdy21EgEwTwOkv+naKN6
BgdB1o+3PBe/nOBhJLkAZPojD57h7S9bSY3Fnf15ThwIto7SreiY1e8O6h2Ork+n
fuK/DSDpEtTcx9y5BNycFfSJgDvWmaFFfPAzWWPxcpUTjqnqz5/umY2LqTFlSw/4
pTdtt8ZcW8J1drnRyQAKoEQNi6tbZ/AHWniY+rTFZm5d9fPK9/6TqqbOPxX9VdWf
tQTgPBEDJOtphgDHi2rHJLaoKH3Zo/+Gjvwg/7AvaNqHao/jnaKJ9hIHAtJRXyeg
vHgVD60Pe9hiigniUkv1W0hxqm0KpnvMb1xGIMg/mMOPlLHTS3Z4doh+3nS177oB
PaJlmHIkFVyaa99obUsD9YbEpgd0Xa5IshdvaHTx7Kg20ZeCal3lY4SSy7jAVKzZ
kf29QHojodTWsGmvm+BMFhcXz9I8W9SdeuwJ7SXgXt9BjB7qrMECyTa5HjDAoDft
PW61Kk8WftwFYD5mqQt4sUwBALwCOF0eNk3B7oQud0BYrddHRrwJxZPA1+S5l4a5
mUMGLS6QqP/48r4kBVSEck5G37fYplb+O6+pIwzQz/9yBA/Jn/SoFBuZyTqnIUmT
/uyz0zvw5Z/ugpMxvCco44H2Ju82yRP7v68A6Xcy9P5hszM15xJesh0fdKlN3fRz
icXIxjKQGypbJj1O+esBPHmEElGkLQ+d4QQS1hFPdHXlxapntqt3bAYgPWLmfQd9
gmqiD6tGkVb++yTsllsaVl1JhVbZLFMZAky9XmA8nXaAlKKTvWUCrJskLPUGXF/W
LFJc4b4Aj+S23FUh+WNpKdySFH6HrXDwqqiHF4rJFPctiMoVN4UzprVfoQ5cMQPl
gRZCOndPQn8pFX7uVrHrnWPZrCyeB/UINFTla/e14yEX0Dp4oOzFxeyffbSoIXb0
EDCBfn1lEoksOvOJgVlDZJJmCOamNpWugN7SbnvzOR6Lv1kpkocCGrKNFsDgzjUg
arJt0pm3z1zh2/oEDpk20zng6AdH8/EHUISbrzOpUm9IsMGHwqU0NR00q6vcjWA2
5n3A6tSRAUOf/17Sqdi6oRVpCYhpor+yzxcp9McGXjmTUOD7tEfL8UOyuLtoRNsi
TR6QwLjx6M+M5+ptTX5wf444iHzYLWSoSeDoYL6rvvnrg3Vm2w0Rb0qGoN/wOuGd
yBIOrdAt42MUKXEA+2BQCpYp3kdLYUdDwNa9FMYP6MTfqY+fPx8mFLwMLjj+sOMC
r0pSxRdul1Ga5N6HgkxAbEoMlPFH6YC6Dcp9rIVXmBKj5atx3z6FcaO4UL5/deTH
eJhRKpFx5GsVnsn5TIHA483A095g16K+/O2uVuBeRt0ggNvz4qlUW6+spPToM9cZ
O7C1CpCiclMCI46+54kLdLouMM2GPbAR47KqFnbHz+TMDxN2kW/YxQo5otdezdRN
lP8/HQZKLe/xSHAbzFnWt6gXlwcwBcDAwWpyc/RuwK2eeQWC+UAZvlgqlfth2aD6
A9OhOrileMB/bmPl6mNeDELjNBTB9rB7c3uP+fvx7mo/BMEms6CAk/LxlNXq81iE
AZiB2QTU/mnRQdrdyMFSH/T3K5AAoTX/Likd3wPESsDO2p3uLuJcMcTBnTDwviVq
kf3pZNH712na6hQbNaloIOflYfMupkeEzdvgX8YVeym+GUyUXr3IlZTdmOnQ8f4g
+uwtbSif7XAAsvZ7Vn7ZxXU+g+LtkJ0lpOOBHsYoEaeiATI4vfjDpADSgZ167d61
LaW/a7KJOm97aX1045A6T29Ac7UlFaqmvmxkJo+1cRKW7FY89yGWVzggEJsPjF3t
Df6VHdLsBrvLfSNbHAIUs3wSovUtWsZptArEnuhB9n1goX6HETI38dTY2LPo6GvJ
t7dGPmQX5jDrw90B0Z4XwJlsCU0hAHfViPiTjLURMj2O3ncPmHedX6mEeUYKGdW4
lRiAzWYcudA3kHlNYT62Kzik1W4zn7LpoDjeFPh6jWwTkS7SvXULwkqrBGDnblq8
vCo8NV7LB4fuTee7EWLvOKbbLpxslkq7lbtEaN6O5BSHeLglelbf1OF6BKUR2SzM
0l6esi+Kv+keGHtscqLlK79bvZr0FMCU3rxGlCnJ3PoiRVevYUvJodsUM3H+yFej
MiE/nVcN/H+rJwav8qOvZ4LJG5BojrgZp5St18IXjfY1jxMvBuMlt8zj95qWtkrc
1cqMgMoBv2ISDfha8QVvKN8n3wixw7vKKwdxzdEHhA1D2S1oI2vgYTKsk9KZ7vnx
75T4NYIKmfDlHZJ5InJ/KjUwXI5tHcw0JCzWrRaKgh4xgil9FbgW6eu0PnZVHYNl
fv1Tmfa28mw3nyeq+4pxzuhbyh+1p1X+S4RRUxLE9ibzVmCt/pIOibSb6KzabKDe
1uA6Ohp9f9TRNB6ZsQAZsCKRNTf1bm6Ia3pJ6PfYVMawMUoG7TlTVJF49t0+OWBH
ss6Dq6aFgoylWPxwQrk+srGC5SiYGWRiepR5mwrF0kEVtMOD03g7NRpGN27CGlo7
KOtQFkeYVnSZFBiJiEO3LCTxx/AXCHcdt9khaDWhBO7x8cSIMak/fH9b7zKuHHl2
OygP+mAC+m3RVbGkhX5u3txKBsWEbolpO2fjU1rC222AGW449BxxNCasgF4fINSa
mGGb+udvYbij5YRQyIntvEgKrYvRm32ETC+MZyNyb4B5PJG1n20ALlamqmTNMxd7
jt/MxIDb3yopMTGthBw0QTSYdD/dFjDVlatNmFFzDU/bE+ie5xNKSGP3I8T1fDPG
ibCgOJYDUHefC2N+JVqtcw8Qb76fPMLtiNemxIRpG11PN+NlWIVBaqtUaDXE7dww
mJridITe0khHZud0/rfdp618IZUccO/2BYu+jzzFOeQOHc+KH68VdKispZggPBv1
dZYIx1wMZ+Co94ZI+v0noYcj2s64Rhma3ofxrlWJKsElc97/TwhZGCJkxLbOhtG7
QvWZHxdmeZN2qncV4UWNp3WFHo+njUdb6G9ekNwfyBVGTWyol+cXGq9Op0FP5W7h
LoQvbxJC6TetBaOk1+5AsEYebhkxUlP2BrOc1CEHBH8Q+g2/4RizYa1nvBNogERt
7zEzvj48/K1ki6s9Ujd6ixdvQp/plZqgmlpBA5QlApYAf3hwtCqk/u3GPQ6aiGtj
NrKGhvoxrAtuBcS2fdjMZDDtN6TB57pFMKOAaftF3X4iqulCdha8qj76fEkI4oil
+WtcXwIWOQwQEia6mk9MbVW3KWsCJJ7kh1Zgs+QPrmuTpjcbjuAkgRkLQJ5Vah7t
pwlXTI3kSfeHY/lfa/bocclPgBhAdGosaGsOOWNQZEU3dN9TD4X+0gv6A3J53+VW
gLg1OZ4gaNBozLO4Tkl/Zy7YqWFHOU2XsSa27C7u89+Lbf2Eo0qMd5e7K/QeM+rw
Hng7Er9LWuB1p4sfxffciRTS7cGNdlNv7+pbuA35MVkMYCMN6VEspXU3BYeUdRwG
Q0waCHTZ3Ea5+GRVuMLTHAHmMi1+uJW/ioc19zUfgHl+JWPnTlzuEJkh2FPRaEK1
OjxCLeDNRbkYfJXbt9IooKIERKyy3rEnKce71UBwrKuZFZl8tkrxO+sVUmHpLOUS
fAYptREcSnLPq5xkflMRw/vfHjrQVBjKXrZq9kl2+Xz8a8ti7YTVkcgHkYPbMypK
xSK2+B+w9BQ5lY73rPdGn3Vb1+frGakHF0PZG3BPXJPa58QQkNXcu4CUPFU+n7Xa
J4e3MwI1HOB83TWfRfZW5MFLPcKnYCDT9FDS6o41dRpyN2tfypPJpGi9itRRhlz9
rfqiErh0Vj416aoEWvg8PLgzGtRPlRmOmk7r+5RhweTTu8/q5aQtYxpyiSvJ8OT/
Qca6McPvB17d6lkzuv1dh8FHey7aWFRnazsvu5gT74GSdB7HqDYjNloPHvEnbitC
72v2kipQ5wOmhy5BSs4RfMXlZdvbrboyQm8AbmMjRQfzdwmVSNzwTQailEqicbbQ
5lwRrMzNGC8Fc4gEMKkelbh2KDrfor6QDTBGxr1A4lQ2T0p3LBl3Z2m8+f8TRPSz
kdz1WrgEzphC3SYB7JvxiY3zJ+qfR9xsJjnbKUl5xNA2hycUPA2q4ySvrZSEM1dn
2xNR1xP2lCr5ya7CyCncgCom0Wo+iZ4krbh89G90MG3fCWhHoCcYyajTSCV7yN3a
ipRywmIDtVC5VljVPk9C+fgLKR+G71GGHpw+AJcXv/J42QIZf37Ub6d1ZyWav4oE
3AC0KN1S76EetYovQKY7N6uu+OWKGGJyWoJogwy+4XZCX6bQOSEBK/kIEiOp0WK0
q+HGM6OcijAPjFD4Zm8jqwyDGCScwm2v95cpccvRarDmPQGEqqT10kDF/opiFisc
i21C6rSXhswgyT7edHXlKStXSJhZHEtxUoiH7FESM6+I+6+qVdDTGnIsa5Zduyh4
LGFhnUfUEwU2T6LxQb/BKWjqMZsVOomQcj/BotnOluW3ymqJGaHhPqnObuALpArC
q2aYQOgX3k3Cy7KhUIqNcGQUElp/joj8lghONi03Iz526LSzSB6FDj+o3mPiFAo1
KB74vt7rrnxdtTg5sXd5dhA5iwswvfPcrHmtes22RFt8xB2822aq6Trx+7hMFZ2u
PgOkSjdo2SRIPBoJXvQ39z2RhHdABynlMO/MFjIEYeAyifGFfMoO76q7IfC5J2LL
VK1JxmBR+QzJskMCq6hLWFlzkfrQkxZU0TCfHkY9hDookV/8RDjgtZelC9Jd8mGd
p4OjFieNQZLkzsyTcqkgrsJ2X5XhJUqb5qE/AgA8vcbBtVi0BFRL+XfAGyBS7650
w6p3S6nea/S60hLd15Q5FMSpG9k5eEnuMdP8m5Z78CaLEtAdLxE+UHLdSCIFSWFI
gmwScD3vVbOHjEyKJCnHtzUJeOwHB19fDh4sWS0ZrHGLdzZ30hutyoKbDiT1iZzp
kDTx6kVk7+fnLEwFQ4DgGjV4vZb9plZ41q9T38UmzrBQA8x1uq8sKwt/VkjE3S8B
g7kO9Y+zCbHdFn7OetsHJa3+WiFuf52/erj0RYcP+p++N8PpixmPAJimFesbDJVT
U8S4x0KicIZ0D/SFgIcdzJofe9DuAIHnyp9J632cMjD3P5iVAGA4wsU5/E85XTtQ
FrwqFSgnMaGE7Qz5hcqofON/7PYwTLvMJTw+sMEODcl1VUKfzVTavbzUjw0ApPmW
gF4DXxdCcLe3A8s5woQKbOt4FfSckHBGZ5kdlOyAJsVU50U6dIDs1lLZVFLYQAio
36+IJbSkXqCa0LBCd7vIX62ilk7kGM/kQuzEcBgrKYPaW+n6Zu4mjupe7S+VEVHe
Wd+LbZfw39kLkBaCJRWeDb0sXGaDiwhErdU/fNvcFpZDIoo4dbwsYuc+Aq+d6bJH
0QKrLvaLjj8KyKNmQt5AJIIDw9AE37bd6e6mSUIJ+J6x8KxqGKhcswRDtamNO4K4
LnxS2lxbyLRDLO9kutipySE+f3SyGo6+yGFzD+2QcIvplqW7kGJ7ytO3gLp0zbop
tkuHCgS5Xt25IIFQ+g0IoO0EnEvO7XK4B8Rzk6NsjhKjycr2aQE7SdH2azAzy/aw
wPv9IqdvHq2hyeUyGOyPyifsok5nXwpAGB4IJdyG0t27elm+DsuO1+KsO2t9Of0T
//KNV/KZNuAvqiBUl4Y5SNFwPikjAOaHi7/2Nl5DoY68kGufxeFEATSONwY9DDUI
XQ7D9dJvJHlBwTHcil/DS0sM7b4Gng/3MHpIRDVLJn74LiMZiMZgW1zOx6YGZrz9
BfkXh4pKVj3ge9hrdwV5dz4sF2BH3hm2huPeSHfg9MONJbNZTfbvau6OeoMaYKMq
lT7iFSJHruC9pf6TuD4MDNMWLXutf7JwLd2Xwl90iZ1/jk8K7/DlTKo0lhk4blRN
uv9XmshD/6jlUAC4LeGgCWjXSPudA4u5cnQEy1xaTxia5WABhZEkAuGsDHxdTL66
n9Kb6W+M/3TKRisovdPXyRyxs8cxQB2yciB9PZaFlcoVjRTJh+UhUhcUgBofUgfW
w7h4FTfW/eZ1mdJb2E9KItdsRM1bAlKeI39ZW3z4CWMJnq+GhYKFSea+IKcLk61g
y6qY2a6PUVYGhWWO9de638g40JvHwkErtmUpJakMt4kqyYB7RlvBcs2bxuThMfHu
abHwmTOTcJy/KNVwqelRrJvvODYi/+CSVL3/5mUiB2Au0usavGn0y3QXxqVKvtGf
OVRdS/qKVHjtIK+14zx3kd7IV/uPHhEGIUWxgsC/AHI09i2y8NDV6GGnB5FFcfiw
DRw8AnfVKPPdsDZvPZFQuOiBEQwN9Oj+N3Y7rmn9Kfvhk4S7mEZS8gZtAmIXLsLJ
jkoqIc+6CxghnzhOxO5R2PY8Wfyqyw9fWgRuhslyXdS11nrlMBEYSaOuyKi67Y7/
zOWq10xmto6ZEWVqeLtYOQv9PENrzHsOfD1q1s7bUQDdWT6mxCv1Rqz5uL9RUoov
k9viYVUX8nthMVWiypy/3X879u8K0T4zI7zksxXIMqS06RBjXAbwoOlosUL+3cx5
jR4+73MEMm/DVVon3OX3bpLa5pXzPMhu/Djrqq591J2icK7RmzPs7LqqIOGqqLNP
hc9dek8eRkP9J1pTpS2ofGZmcD826yqgxgyXuiA8PtN95D1cczX/v7WdVxIYyfD7
4jIM9191i/wcjdopKx1PqW9pBafPnjHln5w90AT6pCj9dmJIfMlDOqPmu8gtKGNq
f04Dizz5bcI1pltG8YtVJzCMLkJo2U1+yjOzDdyoPQLXIXY6Hi9t0fmIMGroJpr2
z08MCN7fhW7TJtaTayl4I+QaNbG0GGYFJYjCIz80gxciVgffclSaxeEWkBRSi7QO
tMFFSe7qd1h4pJEtZvAHGWrQm7+nQ0/oTJBq/ITxC64q80OILmd4Kq09WJFY2J3O
eM1a8HB7gJlbky8WCyA9NmlW1d/7n+4Kdkc78S8819cpiDnSgSfSuX82KjIqskye
9RUBZCU9Se/DghFwkt0/hkyE37H4yp1EIAC9yXenQekuLYyoNHHWydfyq8emgTAH
wGljrxv/wxTyXG1itzNn4XsSWf/C21+ltnlNPc0OXu65XVA3cEhhVx5o9z/cHJnw
tLaP2p2pZgj5hMF0htc6lp/s0dhtRjev1SZnnwUqodQ4oI/92e3fpzWjnZb+1mIa
FeTnFxgb/Klkpr1lcmRv8tmoCO0T+azrFqRypT/ES7LwLnHRBGkbi5PO7EU+0wjU
n4s89FBJI/Ghpg9Ef/e02AfKinXdFYr5xiVP7kOxzONtKFnffdbYyR+D5xPgzier
USy2NqqIyUA91xV+OiQIclkjMJOXyrSqTTNaGh6ArndI8AOHoLj4x0UCxS5xn4CJ
4mutPfHwe82N8Z2XO1a156I3akiuHxW0g9uoKt6gnr23NJD7ELn0QWJ3jQg8FKre
lk8g/U8AxHtwDokjt+apN6k8QZsiBl9Ais47vPA4ly9KcRbnwAmWcG4lcyY6rF+a
+LXZTJJiMe6WPA7nHrpjPRsTnEEra5uhCIE5GeXoWxyknp282llWECXj9nS4Lgqo
QhqoLYg8MAohOcZOnbfGfe+cGYLATdfLxU/itwIJHhdOAX21X8Ws5CzmZ4k9zLdD
ldQNmJHDDMo8H6kjoYi1DQ0oe1suIZbIqgcylqbEL1QyY84HP4/bFeSH1H5Zg+bn
V6VjLXV2JHORtKkONCSiNws073GBLRs2cYaUlEr1gC1VkMvIUv2GNl+HNprwZXbe
+3ruI59tcJwRS+gENf3KTBswZ3w4LL6zXd5t6We9+85eBKw2/SnwenRRag6I2QZd
qusxezo5+PIyMkbgVjDLlwdPtlTc1wvsYsz2iZNoCz+KE3mfVm29xSoKZ+q2f6W0
SkhKOmJkX3z2u87ftssdGPNBOGXBG9AP0933LmOd6vZYdoV5rII70U19o5EVmfTL
54iyKJm2g6yEupCyyoE5ChU0UsF2WRNm2/Hn0FQTlYRFpiBAH6wG50dFer0K9gvg
XPPJu1RdY4F3qVvk7fH6OyhygvGaZPl6mktJaVzJqVvFp71D5rZThWfN0MFV2tSP
YevkeJAdZyHbujhW/meVeepoBo7GyS4nS/H2dRID8lcF0C2ReBPwmXlu/+8E+Dry
TiH9kgVV0L2eqzR0u6K1EIfYjcSvuSker3hlOni2ZyYKjCJg577x8WPR/4YszEV/
7qlQauSm6uAjq/Cs5FeFHc18kr99c/TxDO9/FmJLUIlOykoMbk1DDqY2JgD7da/N
FjepkaN5qlPd4F11JZUUcqIXObR16asyo8cGaFrkopbOs9JGAwCT1rk4a3o6bh49
PqkYq0OCe4RbJQKBDUBMPbeWCdGcC745xD76KVymE8MD1LObET47sjsrAxvvtq1m
Lw0Lw93qjAtrfb3G9GJVkcdgUOP3DSogb/Iol26yY1jO+uO+YXqjsbNDtAvXZp7n
KMSgoug7UEhKKFkGSPAV8/RgO3tQzpH+YNEP8IQW0sInaP2b/4a3hDVtffa/aqM1
Sw1o6hqxqqa5LyEYdyQLyW2VytTLlzww73ZtmiiKAmdgWw1mnY4WLP0z7kTMpR2R
A04/X0+OGuYgR92YkxWxk43JjBNxmR0Uh/zfFbl9g2EzJAGCh+xyJqyM5bq/Xydx
tV80TKq3M6AOvO6hf4Irtrduu8+7eVyABMgpkFj0UOkvRbKACROTKhJYV2HXlHP6
lPzY0QrCsqSSnrITSp4xy4Te5wYrk2fVDVFD0dphn2nayxVp/CjiknrwTOeiVMsJ
n3Yx5Fty1uNjZQig1XdAfflqoLUFJxa3aE+Oe3uUBeTh8xyDt2DMrYYurIQTTplt
RAm6spP8FlFOcKOPIi7CS5aB/KyGXghzJlEDxQFPQnlTO+gXuo/Nf58VT/WRvlZJ
p0v0rjKTj6OqewwuEc3b6CjbLRfP8Dx5i5GDQLqwtvWu6BWSn2kMnhneV3eo1GSZ
jVVhc1ZVLdap08+gMwcMjdUH9QoYKWPPpJVGTgxGPYnf2Ya09BeJe1oJ04cf81oO
9HTAf5D/Au6cud7z79yGK18R1TZMrBp7tUeafHCk6gYcK45H/2tpelHYKYO/+X0n
gu6qowWHlQjAMV1YpzX4PagixKtpnJRmD9Ow40DO+4Z2S4PFVIO9bxUXHEGJ41R7
MqRSSJI6fkKmVpTbGyKYPt3xcRCYggcEh1PZ3kJj0qMOGp+rev2aU5obAjUhkwDL
MwqsSyRecyJ9/YP2lI0IAeV67nAtnzyv3HAaR8mKBLkbw8b3LKrNYC1dg19lyuk4
me9PJgtgJ/VFgdBVkHS12tfOOK7nCJAlnAWfXSNBnKCioZ30g/eGQlizK3tbpK4P
DWJBB0Bkr8v/C2B+mBu0Kj4R9CXhSS4WdRzCBnLnD4+8vHYKKvnLwKL1vw64l3Lw
8fYDw5fp/CEWruDHnaHuD4bSqR2YGWTwfnOESYnjjj+N9NC2RfNd5anuxXgCV/61
Z9RQrweXEqW4doPqQU6R8sgSavyIAqdcOvx6wXEJW4l5tNNENkA0+mFBpVuQ0uXr
16d6XCIQkeNtnSCXy1oI2wPJp36AvlHA2B8JC/RZ7vckQz2dLoEP3UlB6FqNhtdu
fLSKqPKNHqwcgV5tTLZNgQiL+aWL2jSC9mimKebGsWcoRplypHodfK3kJyZYuM2Z
YXxE/ZgHbp0Nk0Ftv/ZafBDomVmFfonRO2s/uIHw1vQstlZ5V4yKpSD4xkyCMow3
OuWEsT8Zank/Xmj9E00u+9EZ7NYhaklz2GJ9riZqhjTAmDrKreOMTDNXsRjNXh2Z
uONDrO6qsZSh8XyuChHq6PbzNLHMjCuSzt3D+k379jMFCoYjZhu8f2JzNtf3HBOo
XP9SAFi5KDNq4g4MHuG3lN8KgcPInbh1GbYtzlESmfqS4m1Pt/Nlj8cjzzRIdaDX
8zc4R5we6O+3oXXlwKLd3fDQVzjiVjP3LDWjf4hn4HrA7eBCVQRdxHXHDWG5qhZn
zZgUep3uV250+Nw7thLAX5609p4DGqw7DnBt9KB7bby+Q9eIx+JqXeLALdp/I85H
84lafHjBjNgagG4fqcI55O311wYHjuuJA0uGVILHGBtBF+i2rYPDSX35d1zYw+l2
MZZFw+55hIVxwtTQdV++TQwOnQZxCE6xVAOkR+7di3S67T8QqXeFAZL6ZrEfP0wv
o6kPlZYS8UQcBX7qy5Re7dMYb0mpKGelqlD+WGmcRseuPsGt2jIOGegQp6Xwlt40
aUGw7Jj99OoYkDEiCfzqWmgor0C1wpZtdm7Sg2Gq3cUFMpa7TEw2d7z8H2J0Ek2b
oxy6/olMz5FQZhiwTpPfpgM3jhbZLRrAkr1p+zvhxqDM7DwkSRSB8IQcQP5jEhlt
iJQy94uzWrIfyQWep4k5lgbsTDnWEBICE8cU+QM9CEWOF8HOoPCZyuK25UiLF7s6
twCDBsRZVGU1N77N/oWXWcY8PfIsO3c6bZsNHlTec3TvinV0r4birdzsR4bNAqsH
LYKMUr2ArutfNoCRNYLH9x8d2YSW2dGJOBB2CK89HZ/NXmBl/SMdJarbK3v2iDcs
brzSyWXT72C3UVzEpg1rYKYkHjIW+vRWm7anjmgklkx+dgRmVcYlwhrC2DjKBTHz
V3R0em0eVkYXTDI0qAcsDcFkqHwDwbLgYOOBMnKVXf1SGD0OY7TytmFo69vD/YdI
rghC9b5X+I6/l2xZ0971Nyg7gVxsiWaQkNCcNY/QP4AgM0N5H/SH5C0qdcVSTI+3
UrKb07tmkPnfVZ6M2EXtGPd+UxDhfgXH/BdswrO2Wa6Fj86KN51P8bxIS4gcCI14
Xf5pmObAcyQuZrj5Y8Pxi4ULfwM9s8E6J2JisSNuE6aUMUU0CmR5yT06zNq/VLUp
szVWoczIz/TCvejq9ySBu4l1l1R60NMe2mV5TmbS0AqtGZnZFN8Fo24IcLPmz6dG
KSZPOrJarw/aSX2fgIaXJT+S/kr/SHC2epETG2nKBpFQG9gM0E+Ca7/Xwqft14E8
82KSSeluS8lQ6oQsy9dbjkysON7/PSbqArVM48WzANnqFt36yoPDfYfqUIAfsKNL
7HhwU+FdgF2e0FwsxYiQtossnsB22Xq8o2POp6ZNQ9FVDVdP7LTrAVxr72MCXhTI
4tQuOiRVtu0H5DY2oRPwiUsNGuTAqAgdYsMo4MmoQXxeQERkPnUY4c51gL5sq+Zg
pBCQTITNcCpnyMh39aD/S6k4G3FO3CzqJUkxtGTnbZ2q2JikTkQn1TX9xjXCoC4L
kCjVz9hkJmMe0cDe+hYgVmOKc1WwDmX2TsOyK0Oy4G2k2Rxz0/u9DrnKBe+7A+R1
Xr6OlNjRJS85WFVf9wsgMgmE5Phps+OcL/I6F+8YYvqK9VzNoBhx5snrAUg8h8wS
n/0D0bcvknAxrei/W2GNF+ZB4MAewdi6qrVjMMJXEpmP+vHBQrXxp+ZGFGIMjA2P
VqOqu/sDeefoDAoIhecFTtXHJnMgeJzBMPQK8LfWJbbltkaBVXxQjNboVkdSsWK+
4ikZxhAWb5JLpC3jmGMooho+4svTJ8eDdxHt2pmvGMK4GGc9c82EcrxImEIZ380U
mDZX0/av0Tyn0+5AmSJRv4Ww6ZQwIJ4FaxkHe/doOZhMK2ccsMBpv0GyahnDg8w+
DV2f73Gqc4ki8TJkwqbq6bgDQMjNMC2YbbIZiNonR2sgAR0A8QpblxMAF9hqW+Uq
F1aZ6AHbuNIw3wKxz3lDWkEdaFYKwCC8FAk9BVm+Q4B2LIbUaihUDyl7R7m5tgcF
YvBgyC8BTxqAH3nKxyDjzDHL3KdhLK69djQk/UcA7wqVsmEQeZEckb9NxtFhQE3g
iJO/1Tl0BsIKFMEe1G9vdgHpk6LjTzi8i0iObzHkwp5hJz0YErwUJdKeDLVnsXGg
xW8DCTksUmV6qdTlIe5KYIBJDsyaeBT4U0ddCeeit3nOV0vyGPsRCT36F1iR5mQn
5nPuJ1b3Rmk+/l3CzAkgBLQcW93MRXxmrRlFf9UJQmkFqVwVSpX611LV4tgWcwuw
s8HlRzdaIA/LgfRtb0XHhtGwCs86trVGejFX8wnnM9VVbg9zoS57yPGgF668+Iiq
LNFVa+BxYZkk3twnNM6gfCbQCVhlRad7AljJzlkeahCMR84WUd/wfr9lBKxO/VQv
Jcf5MpwDxiTFAMXkiP+xg3GWSUI+vjqBR/lmKPtGn4IxeaMrXw8hGA7SandXVuE1
KsHIuC73qNHjT+c/hIu3I8OS2o2/saDJlYFr7G3njsY5Lk1g6mPSCdZZYijs0MPs
7o271Eh/x7GFEdxiDG8ABZaJYy6jBgc3qWa03XFw9Gt0vW37dNhky/QDJPexl6SC
4qE2ZYsHbu5frhWh+IHCWn87gNS6ho7PVf5wjqJOWff+GqmwCZ+375dEFst/4Rlm
i0JXm+8jdLTvbHiMAddWLMxyngfZYrbFHg+HB2SrCsXn1kOzBnxj2Jj0C5j5VJTy
RIF8HP/DgOxXxEAh+ouB3ew4Z4CP8gsc5IdzFHPAnpKUqMewxeX+244vWVvzFTex
FQ43JfyKwNYPhZ0aaV9l7u6orc/LxcwWwIo4nI+YXVsqPVFmj8Io1vwO3/nQnk1m
++l4riOxr/BXhylQDZ7aNbEdkXAmoY9+8Sb7fisQfpjerTQ4tcL6jjsiQ22VIwWe
3aZbnQeR/rJy1jaNqpPoO+pvIbePF99KRjH8sS7pcK3oaTqkRE7KkzLodri8eajH
yNnb7jzep8fyTLkpA/HCHN6zMJywLiiAVFJNRDU7MmdC7U1A5ZMiTa+dxX5hCv52
s12B2a0OKG/D/O+MdVn4vkE+IleRshDtPWY/Z/ntNT/4sKpQCt0hs974HipkHTOq
WFbEc0gNtPuzSB8Dktk2/WYzC1ugu0HrInmthMx4RVlo7dgg3BeamDpcJ0P6OfUs
4/r+GqkonPnCg66/rmJO2RmbPDM35JuKI0C+HzxY9umVPQpc5aZSzDhDzEzokc6W
Ia1Tfp/HebNTd+TTAWcCtVlSyKhozYXbnyYXwLBBNg+Qct8NW2AGxt7R0p+8fqT1
mkHa209uXi43NZr3xlw79O3GLZIAM2MU6JSIAqnNUGbmbbU5tNPXWFibcKCS97h7
d5MpBFr+Fxlm+DYhtUhveBVr3xUt5LSnqgcegbDYLh4GW8J6RqK95zhMIcPPPou2
IRKUSd9MtlvPZFvgxedu7sJysPvWiynRcMWNlAMDSuaVP6gihQNHn5yw1YvG8JHp
M0k6C9sQ83PslGYqaxzGKkv4G/KKmJwOqHUZZqGbTnaj2zM3tFbnEolZjHqK6LkW
tkjG0XD/MNCtrAkqRl6miJouOnIla4CNymAD2U4rZAjQtR0woSfGaBaJIyM/NzRZ
GCud3Le3mjWLsgkROeJ19TylTwiBPej9zsy3Y8YGHDcsqfxCWsTjPlcXqZd6umxi
OB5TuwUvLEllf2Lf1LE49J+ZI2/POPjbuWq/wR0AgEe/lfuEHyZxTXzpODjWevPl
Xa+7BElZVXfV26wW+FHF/2X2+8x/yo1uJird2nt+bgKSxuISirtGXF4p8C1QXEX+
DNbDHSTeciUscAR8OQCV0oo1+AQsynnZwaMy591H1d364bAatbg89U/RD8Ai8YUI
wlyQnj5LTm/qclJDRigfAUHfNp5xa9mBzB4stXvmRzH0LVocPmFesC/x7AgQeyrT
p9WL9jmwPVZiK0KtaFCVQZZ0N6XueYyA0nDGAZ1aXPJ9ljxuPQBbL8KdXAc0Ihlx
gD7VLwTzhX8uMuuFgYhW6G7hBS2W9Zz/fLP8EGXP2GdkONrLHiUIaO0VSu89/eWE
xDUS1rQxcLf0WT6dVmW/u5aekJghvHIJ1+s4IAbOmVVwbOS6peCLNHcSVVqA9ZK4
yF/iX1CDBomRujok++We7fMWvETqEWXzw8Fy8vq842DftPSB/PIZKrVa87rTK0AX
GkgCi4MLLK6triwHxu27jIE1c/elMPt0M/y/hfNNuZCWsSC8WutI/IYeUJf1qpUp
taRUIShczvOBZHnuGNr4DKQcRq8JDgYXkufwvAE6jsZV0JlRlnhXZd2HFyIYwNd8
0LRdIbWAnvb8LOHy1bb6APhQRm4gNeRJCN52qA0KPn0yUeLIU+6PVouM4j0SYdRl
2/+5dfZ06CvW/BbL8+0BZx3qyFmBCghHGIQQyBv5+a7pzZS0N/fjAsj/Pu91RLOc
mKVy03Z9bmbrfNlHOG40KQxU4CT8Pu2oMgli7Ns7aMPP6Z7psDdPny5T/Y0nnged
JQfqiISjMLKmlXIgKh/jnD86Eox6B+efBNkGRXJi5JUuQlQ/GZUgBdJuM/dwMVeP
4V6TWL2i23hJUgCNBi06TJRennwZrV3mftMJarVzoIYRv3k9X+OrF8tzwkGomv9y
rllBdQAcy9xv9S11yOGEwyk/XTsM0Dv9aL3HEeSOiQ45d3HPJ2UQmpvxNtpnvpLg
PdLDv1+18/C7bcz6lIr1sVpoQqMo4uFxZpjH3OiQMATPYM54hth1XaC/8lal+hLr
2zvs7awv6EcIAN+QOF+8hJkD3/Wi9k2JktgIGXvyKI7KnWkVRM8hY0ZzQADy0XXR
T81b239agWxoaSQ0wS1JI4s32LoJ5+sjK0jug+MDRIimzfB5pO1wHYwAeKO0EF9W
ADziUqBwXv6KG2jQ57zuUDLTDipcFuj6nMkpCsT9KGHbyBu2AVcjlzi3QoChCshL
G9H6P4epbAFwRBByBuzBoSz/KCvn6d/2TnBZ7sUSsquDT6TVX+UcxP9vQQdt+d8D
2YQtSkpmIAC8d+XA6CQVQVnwAyiIjU9Ag77YWVnPlKyeMyVGuf28zP7QD/WU1RMz
XESBNe/z8KaN6BQmbQS8qlZ3lIqX6W8KA5G7ZvaEWRZW1rFDbO9KCAK9u0Cfu9Id
nJPYZflALzMXgb8b4j0aMfTsto5aEH0nx5eGc4qHVi1o8VvPQ9Y0ngVOzP3XBAVG
yJdkU1breThJaC7o8+jXQFM2Too/c0a6Jdwj0VkgdtNdKsV58auXbKxT245tNLYJ
wWmfFl8Loucc7sn8OpqGywbvQ3dumVa1GRAaQs6SuaH+JWarSfj4wc8lYjNlW6pi
qNuU4LQvKdMpy8Vomg/gT2zvQ1N7gAkYfD80bUToJ3FF1bPhCA9v0z0IhH/weFk6
WNNxLGwJRCTpoxGVYwPX+Swdw4wgBMOFkTYUCE+Esjf+t7TaWnmFZ5Zuj45xyq0N
46Gck5fXFT34O3NME/3x8nA6ZkWmqs/8b4mY2XPqTvgcx0+Z1OjupD9PqBlsZUog
iJZ8FtyxdLySNl2NNAJmvfS4JOUgutko96eu/AitfNgkjDtwWpOjh4GtltET5XjD
piKEkbpCJ2BioquCUYCEERPsqY1GY9FdLlfXMv1wG9No9FyhFP1oOmEvRmYQY5e/
60HxiXa6N8ATFJ3Mapr8Lj5vcJ8d/CSVcZgeC1qNWMQbbTQmdWnv+RsE9GhPWUr/
4Bx/dQa/LcIn7UN3p50YWw0IZe32vYNM3+4NB3bkcvxoxAU6u+KHFCKXgGJFg+fv
3Rz0DuJJZxkyRBFHUHuwLh0mdMCJYDgVXGuufdyGfsAXMfmo1qXhR3WjEWjFgsub
QEnD5QdlmG1uJAFbUFQLcAtw6JZB9VlOuaII4ChSVPBYbwDgMSwMT7jUW22BJZhX
wT3RcJbISEumOmEgMJZCtOQ+b4qpsbbnGcCMSOxdjY45xFjUrZEKnLciVXnxpe91
I+nH+9w5/GBCKJ4AGvZrwbvCz17WLKWODFYEbGVkvhC6j/vhFF6D0dH4eJutr4Yc
j/w+AD0MzdqeiOjCG64ApVS53DftAUr5Jv/y7s/M50PXgMcWCRQLFBex7ExaCiNS
kDla4q59MTo6m9HoRr//BhQ05II4jNP86GPTYeeTCsscZcf4v85KqHdynkpjfKGG
5L0x3i7KbfUtf5RIGvCR2ukw6DKKvBjPSl68RpEXJBaNJGw1GinLnJItfe6Vqgsv
PTzpyCNGiHY4zlYEFI8eruAczt38uvyTu5BFUzzveExi6ZkOhwKyxmtNNwn2AQGB
rrDMttxpO1vWXnWPhf//JPvUZQUkvkcYayvV3IOUi9Omfi2G1uEs6diVa6enPMlg
pXmZgFIZ0S8j3VkmzMzSW+L2oxKGsaNwovm6e7BflfazbeMt+i16toEUwot4CPgO
tI38lib6xIoWw4x4JtLdnpSqAPYD4N+b89Q4KAE7U+iNxhNLIoHpdtAmWwLA9WQ7
TYwCbAtsfZB3+8yZRkUfZcbN9pyOCr/1GoVWhGLfsTK97GaVVeerkyn4mrbuhhEp
RCB7JjIbw1Z7xBWKYfa11yFEw+cxNRrwxm5x6Lt8YvVMrqGx7H+dQ5iRyD/ZhuXB
r57wqoYbe1DjTAHmlzMhw430vbMc7+Vb+NcN2YQlDqPXp/sOa11REmuqfCpKYvbp
/R6qacMK1d6hdirBkGRpHqWa7Qm7goM1K1B7q+ljVENIh1+77MhNPSjxyZlWq1OB
6K8GZHJbuYgtKVpNq2RcBk1eFUXriaKq8iwOhW0zWH9vbFFrmp/LGmTVgKJAj16C
KC/DTijDP/f5KY7afkJdugXfdGutQO5AsCUPzHy4squcgpWnDXmBWqyWceoea3VQ
HDQdrCEi7K9Co/RyPsQh81VW/cV5ZZWvrgzh9wRsQWKyGMCja7fbaxwxeIYwB31Z
g7puUzJu9Xa+2m9sKeOphLf55vi+iHKi2cVfsKb3Wz/PiUZY9c1K9wszhP5KyyZk
jBPFRKYgaRqKKZ52w6nqD6918p7AZr4wR+2tBhlr4fuozvxdKG81ogiKR1y6YwtI
0+qcfscrhULIppy8gOTl+gm6CRgd6Y8eXtcucyOeoP92dH910bdqxuCpeb2wzpuH
AUfqYfx5H2lKikBxYyHjEVU/CnEJgf6Io4xZsOfvTleJg9DlUNs7H3HXjDC8BlWT
PUjPq8Pb0rLyPyWaaFvcZubeUoJMlQSaHpj5Gl9qI+cp1fbdV4N6GIlfPOW9kZHD
u5w2V682m6nf52jdNLCUWQTizaMFYlaJrM+eRg70XylYEeGlpihLDeY5VqM1lSAE
CEZpRHj2v7zsOZnLm/Qo/kiOaaljStljx/1ztYiX//Ez1ibQ8VgldCGJbBh7j9a1
iZNsUUlAA1EQEOgeID9HqjABGAv0cl39LYNA1F+Wqb5Iwsgax/EEsMz8mELLLUkO
N38AjH2pr+ywCkAfMvtwl4bi26FKDuTIbxUlAeVHonMl05WPZ277SFLkEsMpUT9B
tBL6YitIrNKLGuvNDUqWXdrgDnytETLSVhv5Z+khhk77bhfinXwB/ow4QyUQGztL
QGX+VjUkOJx30otX+86WXUNtUfaz9zmaPTe1JQJj8hREWwYFFpy9iM6ksI8kaIRp
avzRM3x1fgyi6b0XEMWoxWO83bXkU++D3LFXIUzRD/OVYBLtvUkwAIQyZRSiv0Tl
TtqBs5wCO5GektGp5MluChl3gxxD4iZwcmSxrvPEcuq1oRRqtQx50XnmF5vCEh/0
tyIWkrxr9oHbrTRyS8Jff67mBaTe5NMmkUeOg9SaNU/ZvgUui5Mz9z39Fs5TR11X
oBLbTAHKM8X30b7YUFgowc6y3jd2zP0FL5zpgaU8LoYMEhIdtLfBe++8AP/dVbKY
4G32G8Oz0vP89yzNbPSaYVVfIMoI5fdAG+Lno/QXuUZIC85zxy4t3jomE+/ctAtE
JeYoasdNFV2036CSFmr2gqs3Fo5uYgrG70OgkZak0UQXdSq/wspIPO9d3vj0Fbz4
tfoJYWEDkt+Ce1tmyA3ALgR2UplAa3sQ+oa10IGoTMmgC4zUF3Rey7tX7QBMFIni
ImNdbiQSC0mnsSlgMF+ZkVsL/3OhR+PdSwh6OKvMaHogP0wJyhauS9TvR6Rr+xvk
OlOUn3wLaM329pEDntbLE6A0wyvFPPW/6KvRsV0K5ulpFQT26ipf6GJXJY0U3WZT
qJhPtbUuA0ZtYQAyP0KjkvcLAZKBZsKriM56vexpvMX0BslT9Y8lEgiB/oW8WsIF
66gFIOnJTM0hvYNX21GjMglOVHf9CK0+ancoGBaBZHe0mtt2OJ3IXU1+jDELO7GQ
vpXCZIIzC0V6Tfb7771pn8/IVbwMte7cUJkebaIxPCWlpQzNt2FbvS1+PVDzYl7m
j1qYd4TVYyxZO1vOk752R2ZhRnItskmq4avjdfCEEqzDtgiswgHsKRsR++k2a3ls
oSdW/iwUnWzuflsYF1FFLVLzMwHFi8fkumvOc9lp/rZMgfBDW9M/cn1xp1vva12K
tGPByVRT1QRypOVrfH/nJAWQTCDO5tFdEK9FWf5XGMamZgC0XwlYul4qzasfz7DA
lKXE4Av68aRMmr2q95hAYnAaG/R+0OOGuN8KuT+O2srZB1o4/EhdNnUShvRkk3TU
wAZT62LXRLRugFXHFbSGStbPEstxH2dbBpJc956Mm5+pefWJ6b4CikGApCMIMJYd
WMmSz9/wMxPS/wuRZOfg664DLXERlUhUcmgDHmLnuoPB0UPIKbpCTcXQOrUWknn4
BafFK9NlSpWsCDNAvkjJgD3JNpyqCAKwL/hCPZrmDeMh0rC5FYjHUicCzXisWMoR
HxwLg8f2v2DcMHnYC/ZPSfXRbpd+it1S+r/XwSNOmDRsx+dNksm22WwdcdhQY5Na
bRTWEYMvhb8aIU0dcLNo+wOxHETHu/WlShE/cTRZZ/G6IzvRVrEeJmVdMGWFf40J
fxzKLoPt2w5TQYZPDQ8I6fBHdKsGwShAUGyXzp2ySsM8ZqDgTG+le3cwe+YtL4vD
UfzrXKwbNejR1xVpo0lcvN9hPJSYV718WlivZIG2b2jMO0mnFke8qFAPa/QAZ+0x
t6N6n9GEEkAVttQ6XxzEzsaWgYPtYwF1NPZhq/yAJrtGLllHec+PRvbhc1gDVKhP
LbP3wjUtSqVrpc6hMHgwBQwKvmaGjSFNOwhjAS/4PdVGO7lmSR/jrdhfMTDgY8Nz
Et8pRWc1WZT/bACmcjrDASbMfbL2dA07ggley18TxARFbIVhnbKoE2Xn9u0Ziju+
qv9+MbE9HPEzd7ZqOEAm4FeG+LWa/Kx7QmQ3neU72VJbSR0s83fXPpVjJ/cDZ8wH
pMctyNGig97EzAKi3JHmD6ymRV6D1CNgvPKqSqdft6NDrYKHb7B/IPx1RHmN53ZC
IaSbmAggmjBReSmfkatCxpAC8KZprvjeUUo6hE3MyvnA0cKwqtZNVqKkgo6y9xMU
6HzdcZgx8hc/Inqz45oGPn2kUIiyrHP4uE+q86lZOHLMWcLjLdwiKMtqDPqLBr83
ZraVXeo9wkt1Mt3KIGVEG0tcB6fItJTc0r8bvWPKOOE/Ww/Gm/dvespzLFXBGWX6
HA+c2wa12pMGlv77rlFlS2m1DM5yhhJ7z/e2gLhTvaLggzSelHk6eHYyoVcXEgnr
Fam/+WH0bXq4f1fi0TfpT4+/TNys0dg1Xb+97ljAScq48tUP5Ta6jwvXc8HA2qsg
N9ap4tTy1ThrMa5E/BQt6uIRC3gWXBcvicz3Fbi3TCoBGAWsHjz8B+tsbrabWNRB
zAqpSPsTbebusmx5kRRnwR7fbEhFkCTk6Br1fypsX7zrpAd97SDw5bScAE5UI3XW
5hsue7PK+egOiJdtWOZHl6DqFHL4ZwDGah0pYgMaAd14Zxf1yDgQjjwH4qP6WbWG
0pGM8wtFAsel46OoVSpHzW4CznbMI6REdDnRGDgLeFfkRqSpY0M+Nzhj0vSwn9/r
SHGZBWLwyu44L2NUHl9r7JZarHfhjVd3cf/9gGw5qOzluSGcERLs7sXxDiHhNlK/
hTwFRwpx7tOaj9nTWmVt7Z/ADQfirbGwPSFKOqDijKjhdJgC/jmNmqErdP63ExBX
7ffZe4akNxhpJGdJ4Lzp7CJQZUjQ/+WAVycIjGSIi8T4pZ5iAo6l7Gd+2jSAd+T4
Cdrvy8MDDXbWJ2f9ZGDcrhLwucZjosKv9RtGi9amCShSBMgk4NfPWBLkkC6qp4Bw
DqGrDzL1PyQTF0JzS26nxpSwiTQIKOX1gqtrBQSA1RbCEUZEN10qHRToykplNwWA
KbzPKZA/V8p0xELxLCYAf9mPDY9V+FbeM3D+ZbQkcWuxiQT2jC0N//8P0WA5RZfK
aNu4XAC0Tr0wF6ZGEVoeZQDc3RcxMXUJil1lGQF8w0tpmafWW5L3P0/YczYpmmRt
C7UMnO1RwGRfrbtMWP5Kgtvh7WmpUa4QM393lFKAWQNBCrWYQsG0s1DEk4sr8FEr
NkWLBH8AqaqZIQofiIVhig+onsluICg7HmEy4skSNYZFWffn2MbBEWeoI4XCVaxw
Pau2xSyF13Zg7Pp6UzmgzFfn8jCFk4+T4gdZGq8TLLNKqN0xVKiJmv07Wkpi9DNa
cZt/a+hNXkShu9y6KL4elxbgQy5XgQ22GRf+uB6v0K2GSiCNapV7bd0pYx/RGrO0
oXJ8ggmQ4sOVfcElEVw/zdssvTt+pOAQKwMU5NGZkqkwcITCJfXiR+3hz3nf7TtL
WZdi01lPw7zu2SVbWQLBo5os76jZFE71DVotFzPMLeNBvk8n3VN1kAUIuCskD0qP
sz1uRNtQzjzzSui0DpWjb87rxFh+LoIAuWBsAm5IWhXvhqBbot023sN1zQ6UBenF
a8RyQuX8b5mRixRLX4Xicp8Gy9awu2j2MixKvQuH9/YzuJPgrVgpfnha1w11z9Un
2tJvxD2DZHfK4FFaNyBTiK/qIyPZE4e38xJeWf+isN0NsFGPOidRCRrJrn2cfEFd
N57skVpMbUaFCOtCMXXkbooUjbn4O7aKhodBgJqHhVM6oq0t/t9Agh+C0oFCCIL5
REl56bDyuN1fswpmeLEwAF0WB9g7ndtQ/w9t7crKyiNOC28KeKF/MBfzeEqZBmW9
Sy8gzUdgCzSy0Yd7Pvnbrim246mnO4yAzKxDFb6tE6W7oaVM14T/jAL4gb2q3YT9
fAa463WVkG8sebmkenQW5RLl6aON27tzk5KtS6S3KdjCdw/M2xi/d8JXoANUQhBV
wUO4z/QItAwiBcoRExRsllf7Zo81bj+bKvnnnom//1gXviQTKOJe7VRvp5KQ6acJ
hDQkqiiDworrky8/aF8t732mbh6Nr7Z2tVBQPzYBvbNAfvI1B7K+vywNbyGo0+8T
KBzjSEsEekcStDwuNYCFbb/SwF6npffIVgnQiXB+T51DcV7HwpW3iFrHoXJCHgOQ
sdsdswg+ifEo2J72Axnl1DUvOTzJhzL6PnGlaArff1IqOEoz/Vfe71X02Q2wF9Ql
9frPi2+EwB6QpYt5ZfFv9Oor5Glepjgh17NdvYcws77hpvAgmxCLcGe/QBQ7q1GS
+MmtfGlNBj9K22WaX/vDvKBS8z2u3iE4iYeFIn/aixM8Q1kSCUkjSJ45OOoSPscI
pfLIJ8n16FXCpR7oIueIsSBRU9RQZH4Fxy2BntNssOp+LsdR8XETifGEKbkL07Yy
wbv4/zSxIHAiKgHXrHzpZ98tYAZWOTcAS8QjncVC1iLgnSQcPoWvZQp9v/B7piLy
JfVscDhm690KEe0g+odP+0xuPwSfacuS2V9FGdlFq9gy79JpNKutZALvyLWAuqZ4
FvN7lR0MtR3K7lAOUYFB1PELN5u3C1bmbcBNfyhaCSy16ZMvlm0a9n1Q6j1Jn8WT
1rq0IWbGXl2GacOuNcO1CmmrZpuXZhuxeQzUPIX3vlajL6eomywWenmdlw6DqAaR
eFXbc1MgCooJnkCiCJwff9hSGyM2yVDC+7VWQwbr1VFkPYPXfkOVpg4bOt8nvnV8
t6XyR7ozE/Y46tJP3hOfkWEHUTg8tIaOxUJfGLOIJEar1qBYPuN4+E8ExaI+Xr30
zw8kYkBcWBVYb60gNAod4KBIjy4ZIWo2FAUYpVefU0GK344Q00JIXFM3fO6nyhHV
5MezW0ewK7fzjExE+pW/EQ+YvTt/YY7mVzQLh+8fY4lX3CPOajFL9h4tPc0hXSuB
onnBRsUm/zMX1QagSrvWtCDxzJQ0BnBI9zXjXZJ+sVRzDafw9D1xtqh1PWCGCSlt
86Wz1gN7Yd0O4ci/JiQEAkwHflNcSZgl/i8t3h+T6wRUBuKWgkoZnNNrhMV8y5/J
FRr5g1wIdcqjCwqxt74T/0tqfvvXeyJTY1LEeUMPyGk7JyoRLUypmbpzEM1dBWTA
fWVBmDfafkQczE9Avjkz4ACt1h3qqKKz5RN+pEKQfs9Ke8ZyWkqU2N56h0Y6b4ei
LC3GPTSX0bu96dgY70J7Ez3fw7FvxjzuXEk7f4IXakyQeuwGsDKGq8sDw7+Y2vbg
V+MobuQWvTGREGHyIM+D6nbBgRyvdIAht7eK1VfYstsRPiczJlmXEo1Tlxunw019
JH+J7Ag8aiXhgCENdwf1nsaggXp+60QhT95jU8S23ksaM9YEPPYAtkIacaXIRBay
ayOkTuI4Kr306lR2lXMieNds7hF8720hXdrIddo0TiCeFrGSz1YalmsD+Y9KQAIW
lgyxg5uNAyHM/47K8f4YLRrfSHDhwQ63P1oCBFH2zQGIebyH8+DNqf6Ct40+DZ1Y
REWwg7p8t2magZB4ceRWsSk4UCitxwWIHv+CPl25TjC9Zs60U6KyefQSvQtWUo7F
O7LIgJepgE7lLSl9xOqFICX66FNKS5SwEIln7BJ2xoRoFAO+rNXWPMiwUriaXUQH
sWZUaKdajlMQgazJlaJlNB/eJndq6CuAjTGTaHYDC6l55UqEr/GzLnCS5GoDoq+/
D6bAWrFiINosSiCRWMEjm0XNPV1h3DMN4iIAdhktTN2/gh2tFAV2Xn8RQHnS98Jd
VGPiYyzsCmJTdOnqim6e9sq5E6IR4FaCWvt/07o9y6iauEhhAV8kZueJlp/jo2L/
suqsBftfVr0iiGaxao98UWUDaIAlCuTwzgHoXQJUG/vCFoolaOoGwYiCpzvLqAAS
pnb+nFAM0SGmywAXiAh6gl0STi40B95rGv3c8+eBF3eJaVdtnMs61PCAGw1REAag
0aZHoMsOD5n0T6WwjNcYJVM6ItF2rWfqSHWY0zk5fH4xx/5VjXWvq7DC0FwRQESw
w/tTSu7O6is8iXbTlXJnovzKtm5gkhdCwANQa30oGwqJTtuH7FafIgsO8i3frYtr
P2ecI+dLUK22lHVvXmNB0RmSTKCC4GzmpfzP0LE0LSKbgajpqNVP4DZ0Ouw6oaEV
jHWVvMpVOEp0eMIJ9Q/WCcTMeoCT1deup6U0lHABji8owJXHIijul+3R+mQQh1yV
eTiZ1vTfV38JlT6twHYgAx4N+Sw0IYeIa6xSnyMHfeAKkkFr/9yaCsAtRsGzawnS
NH0vxVBn1MMpyrQw+HNZC9CK4zImIbMYRS5fdrERoYfbFiV9hwOdhGXaMwyS8Aas
aokz8seYJgT1heMeWzz4lAlcNxODdcum4ipqeUqXbCPpREKSlKQXhbtYLMaVKBNH
FJATJkSqkEmhfAdkeclk9iBoVvKiysF8COWSfMyXQCrsY4w3Eb2FTFtEnF6rIl5y
K2sth/4HEgyJ98oiHCGBnVCzYukDmBjcR0u/1Ti0B2k0/LLUjj5mmaQ2vmd8aHVY
McCN5RcIOVFPaRSNCRmNAzBaPA8m6wkeb8cY33mrmUrxF94bOzd8xuJJalTjIlGc
CFmzLHaYlBtVPxuunEQo2K8cVLkNHkLFunk2+pbofaXMKXDIPdnYHkufrDYlJP0g
lhZPSdIitRTUMefP/jt5K+QPP7HY1oHFlaH0Y4/5wuu32UCqmCcQ/PiPidphvmYG
SRFw4dyXEi61oKB/nRr2HbEKNq2ks5uIX71ShRDoDUSLP0f9NZDeM87mEWbskgL6
4LBAqS374H3J0yk/NJyTH1YhcUUNctixBIikbEZF5hMLHn3VzJ8XUpBpyirUrnkT
SL9+DM7qTrwRPPzQjUReG+Q4TNOEVs/BaGZ8WDswRNbL1LzykSES5zvcrXF5dMga
7P2UulIwxyVchd//preA1bPjLGWfW3L3sAp3VLYRhe5BiLTyh0gbjpEleZ9tvk0w
x/IWJfMrlgpSoYZPOfzdPCo6YLNqBQp9jy8nIh/2yCBZ0wSHmM0TSQoIO4NKNSk4
lVg8l/SxOxIWpWfZqfURHiJA07zf7Eoi2IyEiPsnUPJAIkuF/xcFBvt1evD1+tip
1uo309uFJ8sYPwHJueBtxTAB3lyaSoX91Jd3NISQ0z5pPEoIUlahXP9c8biHrRlF
V3sHg5VNgWWJd0fZl+wYdTcbWrKhGDw5+lc6Xo7JqeWyB05hWc+FncK86ozK/ia3
xMjehwHfsahG1kwicnGyWcf54O/VOB/IB76bwgTBKQkbu6+24yUKzRY87kriQAqq
ADj7pAldfJpWskvlHmjU32yUSg0Vn82FFddApKK/BPjuhkVQHAbl2hypBo9CjbXm
zEkNfKVQQxERGZJajqyHzArKct1DtpR2hSY3vxnZkHcULe82TVGRmiP9KO3EuJVH
xHhaR1F0idhcxMwH+cdjcVRz56DJcDBBqX6Qz+ggLcRiP4gzNGU1+8aSEoTiAXrD
aDfeaTv48Ft+UtFXep0hXgCb7uV+zuNCjJ+rt2DTtog0350yap1BhXpOcu5h+WaM
rh18w9HxnK//YAc9F7PoaHanjG/VgEtajicy5fSKmMj+HF3Pp1j6a3Or5Gj6EZWH
Oorx2ofomUnJY5qjQJeMIVxoTyteAHg5k2t3MfWzJUxdFibGPT0vI2zWB06MHzFg
aQdtKYe5JMGvL3GkrDg6vRbLDvR7owQPWIpDYvLkfFijTuvVhBZ87rPRc28fwqUo
56iRySofaWxM82q8pnxG9oE+A4dzrudyBJRmoU/NukJYBnAvv8h9NPuVWJDkNSRX
s7D7U/kW4wXvhre+PQk4xyJtXnUT37ZI7C4YrxurZPbASfIp6Shxge/vpHHNb8gl
4ctC74GVHbq78+66ykzIbtC892mHXKaNxrhjUyC/8OJl8XEmavzx74NktnFNPmvc
fVqUqE4sSm3gMJxegfNI/qLUniJ2NK2qj+fjl3Ch79FnfpM2lkZ66k70sqv2Kmyn
y3wcwhhS2bOcoJ7b+Em8RsQu0I/8BkAI0SqFIKcKyh/0s3lYm8hLB5DDGWVndGUz
629L00jTdzHHkRmQhHiqlZxyZxu/sFjp4QU44OetNXwYBZz2LVO290Z0zIyuq0lc
BGFiaqUfrBLQcrV92Mt8JSgNuIKa7a/2AZXcf1JkoKJXDbyfhsMMGeM/XaOawchQ
szCs4u11/DyXnQlmI/+SacOvSyzWslauVKvOh/HhA7xEO1fzPoD2uRAXc5O2rtNs
ayn0YU4EEvNWwRSZosEG2oy682eCswbSTCGwx5Vwo27LarauIEYjXCAYKYq/rcyI
8epHCQNoYoRbDoY9ehIph5rsFuJUss6fuYHggobRhN7jG0uV3vDymDhry0G55YLD
JoBEmOPEDwBUGxkgddQyN0ADJHLe+MbThTQdLZGpiXA5LR2ykG2cRUiR6YkW2VA0
BuGn5I+Eb0G5evV2XSxftuNNuBpCiK6zC03OqUTmzlyx3NY8P950xZZkKMR5fnx7
ZybLz2jkKfxt/XOV5aPcBRoor0/Q+X477BkOwVCiMRIVGI5NapX2JXqmnND4P8ER
yRZ/SZEwmC7NOi5n9CpO1rMOA17QpMHlGkthc0bOcBeV+rVvYmWz7f82mPBLm+L4
KNHfXDR8+OsDiRVB1unzYnXnRDA8AALugyE5QwJzVUT8XbpvWOOBOGjGjR2OSwQU
WLhkBChw0FX8Pj7us6kDB1LD8tqWuIhfSXB3j+4Kl3r5/TiBa+cp+FieErA6L+yj
O5rKTDRf4mptWRnZhxPXkgAuIqFpkAgc8jTn/fr59hdYQPJByPa0HcYFhKEQrH3A
oXnkH/VKVOXLxgMJAIbX9RC6buN2gy7qhtqVguuSSXgihh6NZlbSZmzeW5fiOPBh
NNABOQI/eCwLvSKr83lq1sJbVfTBkTFrT7BV51JOvhJkGCb60LWLo5IyV8VaniEM
fK8PpOupKo0Wpmu1WqpScMVfk5r6YLTLFP7ydlH2nyUuq9TDcVnEasZO6qg4VzPF
aJYbNheQXU3RkGuoXffYZpz0AeaypKxQewZSGX7lhPoi/bDo7QDX/oF0yx6gDIYH
KZ+9UeJF5eYzqwT2F7w8K/MpaZyY4AWtCqjD4r7e8fFK9aprrgSEEGhUVCgvENoQ
8XoLcB80Zg16LzaZjmWFhxMBd0FS1Peo9ip1LZVkdzPm56ETnCOersz+xgsX5uIU
BQ5qy6jZbs2ecCbjlfp57f1cnZjggNbbltI5dsWypHFcd5Xf5q3qUvFWIGPKuteD
VUY/UlWZtEPDiFsVxJsxjuvbqBHkwzdWrJaSvpityRh1Oqqnu9bT6Uc0vTivhx4a
VeYIZecgD1hPrtYQsQDKvBrYC290RqjXt3wwEGAsOk04oLrwLccCWWD57WEAykKC
ZP4dQDf7lCoovH82pUrMyoTETgcW5W+YNGRVoOw24tVXEVKzdqirzEyPR3gpoW33
a4jI7PVpjgc7m8qrcy2GatVaYnnDMbfPWLF1r4uFY91P9HXnDXTtYqkFpmnTo/JR
394uySSxeEu3W6yllvOhnfRcd8ZfEz1LS5h+JP2Pw6NrMzrFa0U6AUkIHQjuQldv
iyc5RqyjrOCneAo8yS3/DTquIecFrjNhGBQCN0PxZwSYCfaaztzea0iPaQ41UXmR
qXq5L6rdbcjHpYL5cxRCGyIw5IsJDCLdsV1sxgqswfJKAZBFimYagG2I/UhRN+KU
PEmHC4gjegMb5cZ9te5Fa6LdwjIW6zhWXSOAapYAuP1+F6xRubb7ogYlUcZZT1CT
Jm8GHp3bpvUElWC8b4j8P5/9VNRZXIExkuRMgNs+7ZA1MlAY+01sLanyJ2GwVEqv
UnuBlfurbphhGsEVVJIHrRHow3lYKnvDwF628cjBeT6+HhExv13gNZwOTR5/0Sxn
h1TVWEu4HmO+9o2fVj4zSRDx4Tn7zE0TAZhttmyDMYgcmCEQrDs3c+Y9cHLhOYwd
BChUtVsXAw/XKAvu2d+EEp0v8mvJDwgRhdA85Nw0jLcbsAHXe2PypKN9Mz5WBYN2
2yQSkt1f+cVbTl0geA7OemBpB8uKhEjdOH7Zhe6/1wW1word2wrGHq9W8yXGeHrd
zUvAbm3JNaic2jSIRRjSOPGg3Ho9Xl4V1A5ZHJHY5d5f63GKKcqjP0sg8gYQn6Fu
QwS2OIC1pt1DhS6TWqoXEsMCofxHeFZoy8HZFhDJI7la2BX+UArxAiEDCrdCIYjI
id2dQaV4SCwLXA0c3NZe2QgEhC2UzXiB1HaZ70oUwGEm07fqz//PN2GIY/fk+Sjg
7Aqk6NlpyRk8TFVTyhpnJjO2w0syDdLBOQY5W+WNYv+7LquWSsfU/K/5XKEUJT/k
k8m4HHl8kk6ARAcZ46zsdBzKwNvIFOkuHhs+btDXfHIdcmk4NHjtmWjo4mKXq192
Caf8RS2KdV3iqS31mdg50mT9SaTKVfZT6lPT2eZkyRZaLPtwQPNKk10g+MkzAH53
DiTFu0NdLqzsWemrONtAQyqnabJJ0f5gvi9My6aruV6isULomCQDCKy+zmQCwXKL
gev0IhJ+BzGC8IJuhsMEE8kJDFTSG1A/YMJ6mwYXfwLIl0PyunhvL7dTa8P5VXto
WvN/P8iAJxqgf8scYzCUl0v6SzwMLJg3wy3IXL1SWgM7GixHvX7hdmicmScuXJIw
C9ykHMREtl3y2XzXaZ6lELK9kP49ZX7pMEFqng3DIDQceMaZ+FfHrFlreMQ+NMuz
bWptpzLKwfJHizX2z7nhiLbCw9z6uykXslnv2Pk9PPJXuhqXg6C3hvYop2VsiSkE
9qByoHKy/qwFeOnsLE5bTpjaep0qdUFOqkJ7iGAOElRiFY+PozFGJ6oGBu17rnkw
dj4ZCduPtC0vBnF8r0n4MNwcmNPrnmTh5Z8VRTMvhSMVgA5FFXK7eF6iMXBng4aJ
fP1gtsWOhtmiqVn6BfIK7oRRpUkVucqo9zzfCSUtvNZvD/X2dZsif/cPVDL+eWRm
umIbjeTyJL8q0FNQeOAEYQtdZfgtuOg24th43umaEuMQWFUO3QFfEPtYXU1xEPKg
iNfV5kRtNYlZwqT90QaHarbfCO2+urahOPjz2Hh/YOleHz6GOG9j+a6S1rgDzEuy
wrq2pnJXMX4aCHcAxYtQh8SbXO6eYCRyPPrB2zI3oZfHxLixuwxtfni49rv624SY
c09g0NzLKsqj6n7JKAmMkCPIKa2IC/58mdSjwQ46X+pdaVGLVIqnBhrxqrKb1paJ
MU4hsW9KprlWhxUYkogIT7BokXzAWninY4bjgAUMy8kcThK2N11bfyWcnY99fuWp
fH7sTJAbbrS2Ai60dlYgCy1H8I25xJ7G0QLq4JJSKqaNnifFifNPecUsQg42qHfL
VhEe0MqFmmPNxDjxLOEmE2z7Z3bRCM/1nR3L74L8m2AeEoEz1knsqpHCMm96dNyF
YuA8BlNznX8ibhInmTUz/57qedVvk8YJ9PRiqqIQp+MdnaZp5IQXa6gDsfNuDPLh
Gir6XRqLhoknSEMNNpZqmiHlnjUo16qESQk0qh3M0Jz7LNJZ9eqSa2qo+I5m9qPN
/FvZGcey7Xj1UMaXPgygcNmtdvVgikMHGTw/4UjVpSlqMeM+k2cLuDWDxkdxErxb
+8Ltz5PXRHihKG2pEzRg4UjegltitJwYkU0tt5lb2+wmhN/ZR7GhP+X9Zxs+opwl
94iuYnoQljFmAQSbdGEQNZWXDicJ8CNbxViLcKMgt87mTWPk/5y6CNpWQeqg67JA
v6vv1Od0eSLL+VC/bAq07yk4Hhh9sUCabu3RN/ysVw1l1RSj97/rTsd8xwuXnPv9
rTC0wHWLKi8ec62B4d2om8gHddLBtEiMU7l/XJIUkwrvxbfe0oF6ACiaRryRPUUq
1iUb1IP17+GqnE13yf4KyliA0/kW8hod9V/kZa3uYP3+8RWdFP1777ed/96Ae5Jy
t5IVqDdhydTR4T2g66Bfx1ow0nWlNIdfbVO5fuhShPNsBHT/0ac7I+wz5xFo9IXF
0Yb/iiZlJAI6MpEse2/MpbcCKSPf9jGW27eor0effangq1dKxRNoA1TjoyjdyjJF
zuNQzdVl0H3UXXrxz/dP4qJDxjIX9GjolIBNWYmI73j0Q/Zyy7g6xZB9Q1O7NC0e
tXDzG3LAhUPgL2N1BzDP3jttjGhNYhmCko81jSWHLw2oaOZM2meDsRpoEzDOst8A
MxyGZgddx0kIfzc95vuPSfeFYNaJYC2LrDx62EOYy4yq21RwYGCrqK0yfSlbei6F
Fq9AQltR0S6176PPpdoIOr06zSD4W1WzzO+cl//VOdK/FJ/29WILPmob6D1wwN06
OpcgC4zJXd+yK8SIgAc/mA8Dbin60c+50F5JrVUrU29k1BtU0GsFPQeO8/hzDNUS
JDWd9eaUbhegtJtxBC9g/sgKmzVUkVRP2l5ADzFtjnFG8R+a+R9aqldvgdcDSePc
30aUDfDu7uw3u8YVuMeX/dFSQ5p8dD6blfoJCT2u4edvnYEB2d23CzpcbyyF6C61
7G48ezlUgGfhUXCkhbIPbVSdXkLjcgiC3i585kkd27IbQC4r0w5/Qeg1uT9rfAnf
K+ioBvhDWuhtJh4U51JA/kf+sGWHWLeqhn2leXZY3G5mJn86SQsCZvUT301Ciaxt
m6HnM/xbbh1vQtL8zyH9fTXZxAA3PTmOD/i0+vEi/SWoTUqjtWDLmhTsSpq6x7lW
h77KB54UfqfkSF7w21KX2OMETIzoCK5a+jVGJSY/tBLpeQzH3JQ18eE9PvoAq1sV
CnhpBbQKGbsHPeVyEu+osBdA32aJvk6ARxyBYA9N4iqafGjZRyd/I+frn9pGb8MS
Gyk54DTrMpa7cWbWZoXy0slcWV5pem+2mUSz9JsPd/SH+BF5HXbuPEQqEXQ6o5/i
6HhRaTKpMnoIqmK2huk/PyzdYn4Z49n7wHSBftNhibTvzeVHL5KvJ+LBliHnXyeO
PQg9cK3CosrMfkybnrRcb7T0v6481AJ44D68kSYKym9sR458jOT7pPjxbmwsDccv
5CEvoTfHMRj+umQNv1diNdzRYmLIvQLhwrbYDx5IQ0fHpvIyjw7MJF5E03Z+icWx
vpMdOboIVXWikqFF+OR5l1Ml4ArAT8tZGn7pmCUxi66tDfB3kQAApCd4Gz9gnalR
QfUeTb1JmPoGWmmVp1BkVzjXHychaIcTsjmdJ9Djpfs4BRypzbBKT1qmB6HHQZo4
Q5y373/HMsM2vS2HBqzf9C+pRqLK++pStjWaK553bmIeX6raH48EORgtKIa/g1NI
jMl5qLDrT+wDptOqDSaijeGDKH0hB6f+dHp3ZPa31Ru6av2/M6tfIYwtqt85/iiC
g6MmjfAX6eQ3TidcmI+JNrgUnL2v2C1mrN7d7QSPezhjbpDejBdLis74tLn5ciy0
Te+B5r/Rp/IXMkZ89NBG9EM9iconv6DhOE2PU8JztODMNx1jZXMQRrGYTSGF3Ppn
nZAGBtfk2eosJU0/QOuYqhd8x9+Nl5eyuOZrikU6BwW7FWmDc3aUM8RKV1b5NgnN
Qf+0D3ckX2t2AG4kAImozbvipeJo3MzOFDEleuteORKWPxhilEfoTqmilwJQiMp2
K/H1YioAS+TC4o9dpvv295LkjHSX/G85Nf7a/RBp4E7W2U0R60wk8uNwSbrnjdOS
BzViXD/pg2Dg2kKeFjCKr9sHSki75plLKIBDpGwcRoEepKa53kEsZgqEatKtzI4m
klUpeFA16b8Vf3wnt/1STbZphdhLrbzy8mWKjwhREBkuOnB3euDjRs/Fo4kIv3uu
nNEJhj4kX1dF7u/IufawH3+qf7aUTiLVYX+81je7BTfbyhfEdPzVHsuJOO7Gwc1L
Jzyw5VrmfW99cA9BbbRfxlyB+IBvBV4PxQ7WRRC7Oxdsg3U9rHMAOFezQ7o9+wfp
+Whbd/M9W718wxR4xmERm7HtEaVQ1BKznXVWc/ZlQL2uvgQZ27w+AsAOtuYsbxHF
CnBQIU/6BaKXqgnjKaREq6Kkmeq2Vr0LLo6feCEVeGXQs9SHWm2DNYqoBe3Y/Lnq
yeMzd+sGFgiyYw9dY1xuxFgD5rEUENptSjIaUrTNCTIglQUpl8a3C0ZzuFC13CI1
QS83vDBcK+Hjf2UFj8nzg7LgCLa2CL+CLPzbEOFDLVlfsEKxcEIdfPZn7CgjGUV3
Cod03+YI6Y9s1VmF6jlzqNMaE9pJWOkZj11G4EOJ6HJ355/Pttyi6Uh/UkFPZ2tZ
O8Kmt4pKe7LlhQJOrDgdxE9xImj7y45tsnE3Ry5QwDbDqE7ny7+JpG40H7nS/y4A
T/L7KNJjI7SwXzmp6iRHiX7BI8Ur0mQRuc4FGTotJbJ+5e+TJZoSw2Q5Ab8WuNsD
cpblb5J9aNiYkj41wNIRaNxw615oxjBBDpQO1RjBTjYKKu5bRlRPyEzH6LXPbG40
iEcAO9ZT4lrRp4Xw+WCsg9s/dT73eAmGF/eo6sVOOdjNAQjJqQZFVUQfjgmwBsVm
BZ9RyWVnD13EFwSZkP7H82lOopevFwZ/5QmUj2eauCdkpMbuRuzqe5czt4k0BqxD
w7OLW+7e2M6g46od6OkgJENXnMGxwu9O6MfCjlK4Viaw4DnHFmix8byPNqovPAOa
0bM4d4HX3CFqp6tjPQQfLTHYRW9v6H0AIq9YujuVFGiF6w4H6Ayw7nUBJvOiAeEZ
C1pLIS8CHePQj+/IYtHy07Zpi7Qoa3c1+dM4+JX6Qv/4caZYnObmGb0lhTyn5Pm/
j1uQalBzivUDZX4GPkBeM3HQ2jKpoZ6zX7b6X+qAidYkH3C8l7uqS+zQqi5VMIhM
lG3V5rkIjRQy/E6ZEFzCpNoTm/B/QM+CPmunoH8t8LLFfKnWhchpdMdtgMf9Jgej
XsWDoyZKVDR35FDFWGQsDfFM4uiCirotDxfaLjf7RE2AsSSBVNx7O2cbPMVHgERB
Hz7iPYy1U3zcd9yhWSP6SMyFazCpZueBLFFe3xPud4ilnQvgKRcUchhTl96aso+x
xckdMl/Ert4ZRo40SDRxzLi+DpVKXZS1VsuLZi1SLNf4LvD+7jUItRtg1RztGvGU
+jSel/8doyvfqzw3uJAu6lZLajvd/CfMCxq9w37BC+Lr76zydFl7Ha/rcrVAyev7
4eH4unaslzRdev2xrvRsjWoXHcBSkLN6Rff+5pWAwXKAoAx6m6RePq/4cO/K3cLS
DNrcWcxNVo6P6pzIrnWd15ejJw2zc6GHqUrJQQ+CkemMziX/5S8fceuH8Dxws3JR
vERpvvyE1dh7o+v2UPjSXME2gwytvrb6gP8QyhAIAhbX6+4i1E9MgAoJHTM8R0vV
nf7h2KPkrEC0HQQEodqte3CYkUpvvMohnU4RaiZ0MKftrIPeHq4MG1JNWUSVYI+1
+uLzt4KakfJ/X33YrFy9mGUdq5PXxGPUloSm914ugJXp7NwIG6M2XhfCMBtFhF1X
kMHoYbyGC4+wgpYwiTmbjf+05THFZ/Cohn4RH3u7+eG4P+/SlKLOrPZ2l03+6F4A
lX9rpDvMSYRtpWSeK0flsiJ13nO2h6dAMiTrgUzYG9Yq+5fTL7ueFEXnnSA97BkZ
TuBqpc0RrDOkKbAQuzu9XFT9wQMVYUiJoc+R5wo0Kd7LBc2sOeJNhTOXxbvbTQhL
qS9rRdk2Pr7HnjmDe1aS6RTOS4nYYzzCLIqYLbvuIqiaMLA3ejvChp5pwUto/MFI
lUG/mS3X6vLJ+K4fc1PZ3x+UViepwIcPiUuwI3Xq2iGV6ZfiUj6nmqalbLCv7GDw
n2bHG60zsFc/gWg6N4cs6cOL3XpS/Rv1MaivZP6i68Wm2uKYLgRHtgYA0Fsosc//
M7CblzeASPnmZBnpM7Lb7XDyF7/x3witnF+fO/Rx2NCFw2VkL2W7X9+j777FY2Kb
SrYvAs8TKk0zwq41zKKFqg+V9FQgtOLQdUqSZCwN4i6xEMLIK2L9hNHx6BeL4OQD
VRgBDdcfxI7DoxBAvW9q7Boyy1kriZddR3cRYnBa3Asf90SJ9ZONR1xPn5CoJ3rW
EgU24F2RqH1ZR8NtcDu+QWYYpXYk6BGYZdI1XQtYtC1f5ukRa7WO8fq339nHtypt
Q8vVSPu+P+tOhUb6L63a+vhdA1eENQVpqQSJGELlDK2MuWXuEpuNKh574U2OzxWi
gfX2U+ZkkJhdnNzb7XdylKGqrv2FcuoMWyvEH/N5w8tJY0A8dcN0+RN/0KzvPHW9
Gimu76FOJDcShC6FG6zoWOJmoDPxBNOszVGOsK70ZmgFJhhDHFaXJ845YWJe1xSZ
Iw5DN8Q/YHTvKAH3U7Eac0b1HhLoCL5ZBuLLUFGQ+as52J5h6DK5WxiFyUk2WIa8
fhztsKXNHlRywMMJ7G4nP6lmEiSuh7EEKNhzdYQTzYdrOoM+fDEVPXGZSPaXoh2l
l4rsW8OZnVttS3N78IDmco3/BGlljJ/ZfWWwOpsxkitLMFoDoHUoDnuKUlVt6xf2
floHMhK3/5M/cUBB9emaXfi0U0bLy8sV31t971R8Swn2pS9IGdjRa9nA77mG7xYw
VnoztiFovtguf04KEBIyM2O00K9Qhei/fM3zH0eS5rp3PcMK7DyvPQVkHd1iVI5p
A2QMG4IccAcuu+/4EHj06j56Q8hfnTRwoGr77jrPHaXtS4eqHe11Hmye0EONYKcR
392TkPtgCaqBnf6/H9ayIw3FBjfA+sh/U0xHOJznDigRQAE9nAnR6m3a/boRGJhO
1PNnrZcxBEP4EIxH9tL2gCDodf0gYZRN2yQSAUTUogZZ66+4P8Wo4GxGH+2WtNDG
DPAlyucORniqYcWAJJDnlKGlsekQ5jbcvBPYRzkOk+/gPlQIdT7M6xUN50azLfzt
73crzstf2Y7sXytqSGTQzPAVB7ikYFTW59Ocry1LvjnOx+9XYyVr1URFI9aRmhim
znc9xq3zTCJCJZ7ZlZBYX94BBqmTqjHtT4kOSD30bGlooorhkiIIRZIV1BbOCOaA
CJu10cYG1onhKTRqgz/dYVTdBUj8Jnmvf4514TjZTqjUuABq2xSPHYUx/uD3iaW+
/7Zq6+GA+ijIA8F/LNzJjtpjtday7nyUbvCjCUICbVs29NQR1cmybBpGiNW9sdUS
n38Ifh3nBa/iQxumNE4579stv4H6B0pmz1zmwnd1Tu6vF9qRoFHOvGJjh6cqLiG+
WITAGIQ80IRgIA2BDJNigxysDb1SSulYYHRygf+Le1MnJoV/tj1KEgp5Acw8aiEC
/wAox3s5NUpdrOz/Hk9k/x6V6HRQJBWAtWdqIzE95XAIsfnnNpE8W55X0gAMOuDO
17kbRYajFEQDJ/iEm7iL7RJ5ZaPUbtS5G5MoXgFJTrvEmb0R48Bws5/LbL1GKH6R
LWphnA2+fkH78sqpwnfBfNc9pfdfTbRpbjvoZswrzYCQWv+1tNyJ67aQEuF0SZZk
c25GBEYUL5qqbXH9IBTKzpuInILkLrCG2mCCRqwJCUbq9Nmg+x07bS+9JuFCJYCp
7IAVeM+hBlUT83/XbD9SB7MyOHbiLQ1YUrcVXn6RElqquJeDTahe1eTaPtFRJa/u
OLCvfRLkt6NmLkBSBvFKFDDIkJsB0THcTt4c2n71y2wgdzyEYC/k6TjMqxNiwd6y
8hsxTh5HLQtbNRS2NXdNC68GFuwV7+wnRcB7B2Y/L5IJt7iEMxQsyeLyMXBuSDZu
Zy0iJsKxSLnBdULQcUQANWjpiUEBbSCKELlpZOhm67TqILiL6TX+TQFMIOuwtiRG
HSq88IDbbBjtCU6PWIJEkQAPgWtoiDCnxjta6Ui8wYwvAf/MxgoXUtEsM81Qstro
iom5CFKI/TsEkP1YGHO0A3i/FQckoPT3U2F2yokc58JoHPW5gUvGW85pUUaUCxrY
CG0o96QsoKzXbwPOteEflO4JNwfIroIsNH/FBW3gwY0hhBv94MQhhAaFyWX+JKf5
VmvZbvTuUIy+Z2z6AVrFoHD6wH16s8p0//igtMeJEgyO6IDm77ri4ZcSfmL2HOR5
0KJr6zEJf0I7Sg/+FrbOQe8JHYKmx3RHfOB80g0+3UPBRdwpdm6irq+RwITyHqrR
e4MUuqsRz9K49zstOrpgWH2/WFtKp2g6mitE2qkiG2V2zuxnbezzb4SMzXsnkDsS
11PcD/JT/RMMWfUcmD3fpNlQqHZlxFzOJNDwuQBXvk3wg2PtKt7d6ZxaWGZ4R9LZ
H4mNT6++p/oSHOe4goWtuAh+AVQSRiTfI/qZJ5WQf6hdlktQriqDHF2+vJQ7mMVf
FVGpFIJ5PMcDfz1Og726KvxSZQJkrdWYDV0pc705IVrR2E/fOxTceWKWh3Y1y2Ze
gjPkp/WW/wJDVSX9rqBLTvbUgQ2aNcRW+B8VicpAeXsu0+L2mziwWuiSfRqNP5UP
CVJxc68D3pZnbnvzgcxi0B7SnJdKrcOZuz/lyekz/woNFCvUzrizKc5chsPnGYNO
aUvZMGGHEwgLq/QSqwVuZzWQJ7D5pHA35FYi7sno+gVJEzxweRxqISbdGAEB7aYs
5IyVe9Y5hBjYiTP8V3lomdpb2FF4AjEg2MDD+IMXs9EiSKMf+jWvnTLvvK3KTWBL
dtCvCGMoRBfWdMNyNRu02Sclkq1M7JuIBMH9lGSb/hTMajlLNCvoaVO/wT7if9Hm
UGMlR5nPQ7cx5UgLIIh1GmCHFND2I3ePH3njPhMZ0GI1E/FFtziFLXUm9+4q7yWM
f5v5MtL2KID0RzXJcHHN4FI5Lna5uZUbcNL20Vl9Mp0gKFeUJzCAm4VXiNnMV0f0
3xR8oAMT2SLwIySUejotXJXaZOToGNqKSILyvAUdCagBgq0/jMj1IVsz0oOB8kNT
yVnz907m6JD1koZVYx3vRZPsPQEeCT9mwlRV/LkMdfQ2h4APClnX6O+tlU2C/fW1
NI9MGiuCpYqgbfbYWMGBtqay4+Ms956usqQ5UwTABaDCs9o/5aqorCGSxZtbTU15
kOf3EjxC0kDlMgl9yGZNKFkjLZESI65MwY4Y2m37uSddxFv3BOPVoTTfmwlFPTZW
S8wBDQoNiNgRf17iqU00KXjT6PxY5d/pjkZgcDxwIzgPGjy0hBU4XIZhj6doph2V
4NDuKPoMaTBTUUO1WqHcQ5A0hhKewlMuA3+koR7nNMNcuiYiXOSg4hHonh1w7zuk
3fHXRq+cGq7gdMOE5qy5fPh7zOXM8ZAwS97P6uQ0cohzaj2z8vt86sjROrrzRT4I
3tTQ9BPRsVyi1l6fBKzDANxbJrVBlwIKkeUOhxU5brKU3kR2k9eAlIhFIbnX5qHg
25/xTSHHthVToxMdKC2yzQ93l8jYzUfpKgajtpKfl9OHH7qOgnAK39w6T6zzSbRr
EtoQGBeDX7AoMlpeHBU1DR4BHoVk3oqZ+ITef2jb6V2FBnRo/a8u5jswzJc/b49u
ehI7eU8JktUaug5yz2qnsxxPIYQPZO1sElf701cbiYtVvs39nusVn971pJpXkQGZ
AKYwoKZh6GfyQn4eo1h8Frtsk6S+1qDDB/ntyih9SfghIXUEnVvo3qZ2FF4Wd9oz
P7gWJKNL+MQ5v6UoWmUM6t6OGEz5Kap42/ITYb4FA8/28FlhLRYgHDrHwD2Fz2hb
wIcjhvna2VZIxyPGBm48UVLERQUyyBbxrfjqrfrFJdBeG+T8oqsRfKqzTTZal8G/
puT6XjH0wS32UkV9JP2WCzM8S02RTs253jSMfn8FvbVJ1wrvqv/U2+VsZHVfbkHU
1Z81v6smaPipA59FWppcR1QQ0gXDEd2o7c//j6A7T0kKFjYtK+Iy+Nt4Mvjd27ry
i5PutP1fgH7pAHltJUS1gc9BZOuAED+ja+qeXUlCLdXHUg1wXN+EjJWH6ETcdI5d
gd/rc3KaeRh76aWZoDu7NYNk9FUtQUD8g8wN8vQHDpEnhQQ65z+AEqWX9seO2RaO
9yhD8AUciJHmEjjWB99Z6D3EOWcoAjl4pWnA8Pgfi/63SchrXmqSCPYBqtB5Ju0H
qvPfrVTRSW3OHSNKVQYhAJtCX4vu+hFInkBv2Wa6Kn6keC2uXD7xBkI5L96pQmdl
aOagaq00uRVivYerTSIrzQtTzfBaNApPXGs8EcYnOx7q+MCd9hjwlh3nEzycfGdx
qDp8UOweUkkbdForuVoydNSe2O1lPu7Ybb1MGH3el5vF/pt/1w2HKfcZ2J7eaCtq
FsBQIbwYagPUKUOHP4CxMobDstn86qsSB+bQDPz7ZSF4DGuAIwwj02eqogcGiomj
sZXe92IKp89Tfgc0CvgvrDdFpystz1ywX4hlzfjvH6MpimUulTWUP7s3cLkBksW/
7OWlwdvwNnafSs0YZIp2HpOmbu22TvmO0tVXbt53Ob+TJpl+QnBWftNOSsjaANpW
oAdeY9xXIjE9+bhntTkU2/OCmH1ZXu99BK5Bric1fqQ7UAwEkihx+28zChwRGi7Y
qRizigJEjZQXwbHxDqXuFxRfUjTme2i1O4lsKj1OdizWmaLB5pleX7zxgB+7evd/
0GWF+4X1AYA0r6DNqq3TzmPL/k8Iw5bE/+/T+8BOr1bVjN4FP8IJFQg5SytxK8GQ
hplI9J3gIl5qdih5f0f2Vg7V9GAICX7gl/EH0gm4sfSJQ8jAXXpjMKxThyiokpM1
bBZ6VHucbHlFTYRLB+hz9vG7JObsrN0s6871tj5GeXNALYtJvLNbsGDSXaJGcp/+
k2HUmJpqM2ax/ZBv136COkd0BVzdVD/oGcLdmZQ9zmKUCUga+v8cLU7tDKVEh6N7
p04jFGTSBlGIIm8EhMKC2JjWbjRmxP2xCU8Bm6yipf4X5JDcaZnWIYCB68z1Y/o8
EXjzvwjE5J+o4zCmoFb521ZnWmmIyxiMrqW6younyL+GTpcRrvHBNS1//kz0lVDb
+RyOimWwc4rH9d51sSOsStvFkuwn6847W24vnlWffb2PP/pbDTcgjV7mGCX2VSod
TiXjaDzB763qUUe5ReRcgyq4ObMCl9OknwbL96R2rQmqF5tsNXQfkrBsvXVO7B6/
xKbVhSbQvjkiMMfdCL00SPIogckfwbK9tgaeyxwYvoXNG5DgXQh/qWuLx9iUuH6f
h941Vn/VWkbi8ViXA6iJCdzzJWtGOy6yDuAUQghnU8SOsrXbEsB4Hj0C3iFQD9jO
TUwZ68P13cDOl8bpunTImLcqdjAQZGO28g4eoclNMUfEUyMOliKtgOiQhiAnxI/4
USW9wxJ5eEHaVoWzMApCAFQB5cv6iXR41DDfUhfQaEuLW2QVEz+wk7qTjXcDOKG4
inT/5ew1kLhKN/9D9b6XUrrM81P/gyHbzVP8zGLS5JBC/h0ZeBttbebzb9tlAmPz
xqKJcf7Q6HAKXLDM1hl9BVkWz0oQLSdmGgCiz84F59WvmFciX2muYcjFAY6YyxTZ
02z9hBvahLnZeILh7J+iy5iE2OV1VERxCWfkRaGQRQymGWl1MECrPmBsMhrKoR+T
fXNT2YZ2qVJoiu6Qnq2woIqJ7rkcuct5lIZqVA81mcW3hsPSOyD5Ox4QU+2nLDME
pJcSEfyU3hDvW43Di2TZQ1la2ciqCZmKRxivUkcqhRCWo9gYBg3szzFmtJbjn5AG
91y4tSsnzwMdz9cHPgr8BZ8mvSpGFp46JZZh+kI2/3V5LXbZo+S+nQKRw0+W4cLM
9E7KZpIS0gEtL5jqirgZBZHkwUBw2xYiyl63KR3sd7ZT9MGhppk/icoqF4XeQiv2
OsWYDpXzN1AJRlr0WYDRsDZ0sBQSF9Hjz5aChS7YgrQKn0yUvoDf7Z8O+b3ZPIoe
jgnKPm8lsuCn+XHHe9trLtXRf7Bfdarw3cXwgZCzX1LYXFMc1mNYYSUjWpiJYm7T
e2jiAR6tt6kZVNZj4OuNEf83jIaGi/R7feEekafs3unGfI7iiDF1QAJZh4finQgH
Eg95tIW78P1x/e3AnkA82H9x1/ysAABkLeufg+YNX5tAMDKpVCk0ir2IfTKNHOvC
71hwq25ICxy34d8PL0m7UQIDQudyC5Wfo/35wIoS0oGhXcYaLAasinzzNr/lLg5b
2k0a7ILsw7I/zOoRfCDWPWyVujW6iRLyyK4GlbXz5ztBAUs1UWKwhEX55BAkA+gQ
DqlevZWItYIRk/SfLeENsa/Yiq2jrkSfFaz8spJO6l9ZM51VWLhvPGukIhNcp9UA
a6rytNzBmQzStq6w63LN5kqMy4/QWwbAB2hKCZeTK41ZrchyNe98dSXZUEH703e+
cSfYZzp79gnG33hsrPg+M5fD8syUQjzMH6/ZnreVQzz6c9fanyfqWKI3s4/jzRx6
OqN8k8u6yWVd0LL1kZXwubJASWkU5uGy5eyRQSnRE/4PwEF8sruz99foRQYxo1yd
Mz8zAOTyIyfdc/A4JVNNkuLMJEJr/w+lX7F2hRR4sqpry/LEnZKqyeMQPpuF4g5W
FaRqocbhSc8LSAwsWjaXxzuYTTnfq4iEuI5ipsYnA+TnoiLUsbQf7a19SfApuagj
Bcd4mAfLIK7NVqImM3bA0LXp8DtxvcF1I9ERYJ9oeH4rmry66LCZoYjw/tR0MJGr
ftA2fLm6NOyNgw9nakE71l578tGZLMtj1FX81pLls97gv1pOTTK5DeHRRKTw+R4o
hSIR9KcJa02sVQqdkiqTFLGqoSUfoxqrXiUZm5AYBNgf+Kw5PU6C2jbul/mcUxIl
GjE0wuSUvxYlu8kfg91+sKN2hy11Covft9QLZFmid9mgufZWzKAQ0f71BucNqjYy
lcXW5w6Jq6rLgUEOgvO3+jzlZPptEuHtQNqKnhl4Pr3h9ByfMcedsV0Aom0prprH
J2ie9vKx/u6IQMTjLLYB6g96Nv8jbv3sElSmuBp2hcp1Vxk4k0wbfjaAGDW4gUgp
E1XkwnWQ2Ios29FUWJUGhwIyNrjjSZN24Wku9zgMoXsGy9LHNuXjYyF0PlovIAkR
Lco2C8MgVyfMH/cfVMYQyWmHpZkcwE2l5C6dv8ocXabzj8CZKwkFx4n8zzXuMy3v
rMghHkKHFL6tPFUmb8MMZGOIHz/ITH0Beg14Qmzx7fm/+08W0fYktzhp7a9HPR5H
xJk47BcPvJjD4rF3XPulwJULxyUDMz6xXObzbE9zFfVPHRbnJomtQZsCEDuORoGd
rIj+641MvG03tZ6RZwL+0L6C2ClH25Zs++2c64707AK/hB9MnNsJfP0fr9xp77FX
m4SooOpjK/DxvJPrFKIQ1+3c5be4abqScS3n8D2Xc8EfHpeoHJZtLq1XFEdkrUyy
Bt8ehVRR2xNZhzdEDMmEXGwKtZajNu/h9wdJ4tVckYe9g1jIy9KuvHhUC64lwbC0
9Bou7f45kM1QpLJU3tIWEixZ02GG98Q4kjpVrWnT1+8hkPBFsqn9Q1wS4gVvqtaA
I+XfbwarzN1S73epIRiD0XjTWg4piCnIhi92FNFar26U233vPOu9ns/CAEL3X3Ab
7eZW21xOmBf+gBz3jd92x1nfadzuGKsGCvYOUuYvUTauv7BhbRZUpPuh3MJDZXmD
saElVFNOLxL0FcRm3zZsqwOOIzPItPSZsJWneUXfcC4NUzQdxEyiLkqIhyAySKl7
qvZYctdvDCx1BGW0U7L82X7/PN/UTMmQlo87XHUXOCNzC0/z8V4xfEmYBkCnsxWQ
TLi1BEMuCrv6Rb//9C5IQfII2hW5nKy7b2YHPwqrWe2xAV6HVd+64g3vlHSajbG7
4alRPj5iQ0kTf5Bgh5L4IFdt5WHxSYpXN5bWFbjc4l8C6LWiXIJxrtWBOVT/TRwd
xe1C0Tb8ltpx/gjvPjKsfZeKvcfZTNqaPDtIuyAIDMMQoa1VJKLhrLXg9X7YSloo
gK88sh4q4IZYKjssF4kQFDyfp83pr2neLVHw7qEfbi7xWKv0JqurO2R0yHTVmiHz
2rND1iNmll/vtmMGdCo6Q1bAjr0hpWe2QXCEykw8ZoV3L8v5lM3Ykqu7TwnUeO3Y
QcHNBodBBGJiZOfqJ/bCqxgZlSlgcoyZJL7xerMYNMgVTqZnOreThBgQYfByu00C
tEDEAHuZOUw3P1gS2WpKbYyMLtvYkKD6WkjBJSnztWnwQ5useVe9h30ucan5ZSjj
P8SCfpGQwAxczNB9AKjrW2e48+oSOlO8HuLETQvFXYYD6v6WkO/451Jg+CQb+XnA
UQciEuI7Xq7wqYA+33h2Wahpo8PkODbfWisMmnN2tF6sg33x7hNevY+9syL8MMuq
KGoK1fjqmsxlE+usmu+28DUC31Trk4HT9estqOM1XHdgaOi6mk240ZUeM6zn6edH
f1cPspxwNV55dxZKVTZRtM+dK0KIUChvSMUK59zsXP9uFbtcSb3hIbTI+3+1FqRu
ahWLw5FJ3A16fhCeiAKeV2OYDuTlX1dS67ch9RltwQFEKNy91oPyQIZM+rkL+2gN
8W/vQmadJGpnM2Ga1shn3AKa4TN2PWc50H0dm9lFGsIh4wu2qwVfvIHqaIadTA85
UfHdEG4GUaE2FO1PC96ZdKM8RWQP92wwlWTrRAJPOaQU8G8jzKIR5xzMshOG/+f8
zqAWQTRdk15R0XRKSwx9qcemU3YL/isGVNm5hwsFaX0q1m9WK5SoiK3sMnQxMPhi
madHz6FKmLH9JxvwhCfWCORxu6MujxVExWkOKir29R269YNK6U4M0U/uD0VzKQws
MYIHtYVjAKACQcqOibiwkgthcaGu/Ybr2r68jx3ASSWRuJoBko0PETNbuTKFFmCM
rX+nASnR+V0tiWswhAW6khnGwUn3hnN246I0ivanqm2z9nwUxuSB99f/1byf23qs
WNVuVG4Ch5doNHMHPVJyyADz55ouZqe/Rojzl7TcnvGcMwtRAWIFFVr90g2eROP9
XAaHNj4jEuBKNaIlT7VDI5N7ROL63Y/0nKYGoPss/QK7UzMA2EqLEgR5OLBDxhCF
4I3V6cdCpGoZmlRuU87PxrbIUB8cfuV1YYOU+wssboMUBexr5PEEkzIFMkQr0O7H
XF6WYlhytuVO8vhoHwwEQMrEUuK+eikFULKpnAXZIRnCIgXEu/swbgXAVkL9g+iu
jJ0tYNnKAvR+BXivZN1iEGr7EsL+dBI5yiUX9/aiicHD997gbnii8sNtbUXs3/7/
ESXdcyrdSmfE4uZyo/SGkAVNq/ZbQxk3+cv12KXqU26MkAdBfaoutJ93SvkbDC5X
UF9SK6DKwVV2W1i5d80KV35hQqFgARvDmA5Jvu3T+/0W3Hohpxa9OXQEqSP/WOeK
CqV2XRvK2syIo8IA3D7yFQrNrumMUlTiVfbR8qkamr9yyO8vGL94LIdA1Y9RTXLu
FcaLnrsE6qZ3neAv6P1paHDzx5OnnF8UsrDvUtxGi/hhFNfD9LCUAJM8latFJLVY
/8ZJYCDb9vDxWFIt/MA179KJPKHyT945FsMV7mxrnMDjNFZEd/6VrEi+a2HcFnGo
53AchIhCLcunnPXz+gOhQF4zaNnyEBqNnu86RDr3Acnz0s4hB/S46g7TEoUHcWxl
wHw3m6uF6aY2rTHNo8P5tvcoEK6f2WUhDCh0uPcQRpQvHflGF5OI5wPehSDsF/dX
VTS5vfvF5h4ppu7+1NVZ3lEv9CrYEorpj++Z8L0fLoGGPySuTAObkWmrIAUCMsoM
7Z52ur7z8RhoZlLBHwtYpNvQ456SIsmu6UqLLU/gsQTQCl3zl0CmB+4ra+DWzZy0
1Y0xf7bhurdaagz47i7nVsBjHzNoS9Ar8Ehf4uBo5y2B2hBcE6T5pMMoutSRivb1
xbtqM07QBRiJ/TQ0Ns41mfVMFfiWZ0jhRhPiQNRT4g1V8ZMYVQluiW7YI6a/Ls3A
YYymKcg+NgET3CsNqWdctJFWMhi2z6PBxCDzG+X4v+9CxaSAmKivUzI79Wb23yAX
xUbyj0fX+nBt40xDONmTF3aZEnKxlrD4tvqMc/w3a/rSKclwHQAHvTAU9qUqwAfw
XHCJOdA7IzdtZ66QETtJ+MHZMfqfThJA/lW+c3XnNZionbShJl3lGTmqDnRK/RBH
fsss/pR80tmA9YeVCPFP+cLUToS1x1lGZAolnr1qlUeqWhUw4CWGGgrrXkrunAIQ
Clu12h0CIp1EXei52YtrV/5zScPz7UytkJdysdtOhhQIBN9wnBkdbGeuiRZU7Qx9
2bnyGHEmaLlsCiy3plXfBf/1TSLisFijPaDl8YB/3vCvrd/TayHmeUVQN29wVIfZ
/S0quTWuUO4bdCHGMneGHm6V338b7Ob62qWSl2/3QAG34gkewYKb9q54jWO1KDsv
rVPtdONkLVOejk2E+9xYQ+itxX1HmIH4IlnJtcSLyrmlJusPjXWA2lcNa400r6vV
WGSc7fyNuaa0qWy7FNCXKI5h2mS8aU4m1XZMatZR4yPI56cu2i4bBBmWZSBWZmbP
m+Y+ZpJpl6ZibQyRfk//7Evd79IaAKTylb9wAIgYBcusDvMxQ+ShcbB2GdFqWQvC
OMUxTTYTk5tJQ1niMxE5C++5Ex21pLoDZ6cuICLbJgoF4X0UDixfDXP0eKeixO5i
6ATIyVkQEO2bG8bjCz6e6JPq6AH+OZfT6d6dR2XJkcwURZZ8PKZAnBQpmsRUpTOa
ru/8rx/RuhQJtCqu67IKSMZEuQIrqigbTWduL/5X1jSF7AMwLiunuuJRta3/lpQg
MvTf1YrERvR7ec5iWkqB1Kod3GDQEdGSlNcEjVD2ugux/YRalE7IWomJyDIYbarf
Icr6KdDRccmobqs3NlpxWrigKPDRTQEXJwwInbLuqTQOSTjE+Jxs4pmUzlXV9Fkm
d3s+YmA1SJ0DTrESOyNmPYxoo9DILRKG5XoRzW71dEwfGZDEQP+ExB2jWkg+3X6I
gpw2myOjKbm/z4zeth0aX9UCLIFEaT/RXBfGU/UrBjLvVA/ol7Z/a0PAYYU1BkSz
qGCcHVc9TopoNXkMP+YeYM8+4cU9vbMXnvIOdThJGvCl5GVulgfNWm9t+qRriVEu
CDa5wEZBlyQtIZVi/fxb+aNDTsCgT/HNZWl5OmR17dWEraEeoquzxqY7Ja8OEzrQ
xI/xSheKW8WtyowJLfKe4ftCyP3A2uaNJ968w+KaP+eNPQ00lk7PlEyGRaArVGBs
9nRBy1upyfLBals98UhoPanbd3G748r/G+RDSI17ScN++dLMHUngldMtpFgzA8LQ
3BvC8uNMwhHPrJC48+vcInm7zXEpTe/sjms6/0TdfJvSA9VdnwfUk3vWyLJM2eir
buwfHkoUGwfhNASOF54x2w9ik2TkCLaXZQ69FJlX8692/RXcCOhXhm8GY4zwtp5g
t5DId8Tv4YWrY6b7/idIiSAPhE231d3qjHqkGviMnEP+4/t2spJPtHtUJXKTRTB0
7b+/6X/UzGFqektxdAIFAFQUVfboVK6Omn3A2Q0jWNPhuqArCompw2VIcwQHPwkv
t1hkjjtAI3vUih4kzacWX/9yZDDYkWE/DyVQ8MS0YFJnt7diYYYG/hDsTt+hWXsH
6LrZQUTkuNOWGc2758FlnulsppoSWT7P2Q8z1hRWec3GxouSY95GTU2XeeH+Z07f
b4V4CQE9WX5YaoLhacdrc6rz7ehSarckODHheimVLndjC8q68ygTc06gE2+nUh13
F9zz96i9ThmRT+6To8xgA8gK98bHajhmx8B3CJ+GSm7Y1hZXY1YB3znVAp+Rrkxk
2xGwro7iM7UOvGKZ6J18yH9WKwZSi7KZ1FQy81k8hyBddEljEKt/yU+Sx0Z5eT/4
dqAm44kZdfXdX1Wr7ANVHoxf6sl53nCLD5xtYaemXk3fCSRNPw0b3Cm6poeHtv2K
gK3gDCWAfqV3KErWZxEPutlbOM6NVB9kXx1RRPjvJgd2K5XgycU98D3QkBii6nMG
sHMQd24pcWEKyAHDruqYqshEF8ek4n4hz01KA/V3GHArPE+S1mUE1rjoOkqJIjm+
beNUegKMTjri07bp300T3vHmjqFi/ogheE1xrAnzgQubE85jvYOZ2hHUAa2K/aRg
Q1Xi47vMZkzuG2ngxt/XmpYZ9G2cJOEjrGdczn3nVarabYirjU97xhhovG3VJ+yr
Be7hzhAg3j0FbQBjgAlNXh8X7BOWr5jd8Wsb4TGeE79W7M6d4/XtI27sMXuQT1Kf
anE7ErypUTZ2ZPVnjWgxgb5z/WU1jgvfxlbxwqKm91+RPLGpRxs5kWbdP42VLZWJ
V2t21mGnbGmsi0h+Pw+V/3BIJTR2gAO/UmYpWikErLsuSUaBkB+lAj/I/tMuFVGE
kJSbY0IbgMUH/48kQm2IsoeoYfFQ84twZiBitzpiFs4dFwm9IFy7fSbAZW1Q/+kI
imE+TR/vBW7UJ7V86/JSf7TKnZAXPaCRVqshAl8wRkuQRbMKdcsTEz15f9dU/3s5
LRMAAQjQ37OEO8WvsQ/yi3ET3OisYxqNKuDO+qBktHPuxfGmoIl9jf/EbrlwuRt0
taTG5Nbj+YP8T6++O8yJ9HKXOzr43dB0c+sqoz7nIc6z8Ttv1rLHeRrH0PGsqvjm
P2pt0wDV8Qy1yP78jEt6v+P4kjgdEZ0aHWNuk7RKTKPvGSLfivn5TX5ootDEFxIa
PyJ+4pXBqLSWMH12awgqhlb4sRKv4BNapYoPpBrEWn1Sp355+jD7uVKif3yXbWzp
NlJ9FAezzTjcGHhNodmLi4QDQ4GyCa5+e0B8YFnvHSsXlvvt+SgNX0CCN8fmcqeU
YL8WGG0axIK8kAxoRVKypo8ZB8BIq/IMk4IFOAdjpQx6HNUW9Wz1MfdO3dbX7nbt
kt7a3sP4ovp6WSMc/mZBG8D4AIWx0MrvMsDUXM9dNfeK9P6o0pGdW7zkH9WfkGat
N79a1lbgMZRaTvKk4Q39OEzMChtuY18g6RIKS+7efmsI5ysVFF+lF34cLlyZcANE
nanOOwrt3B4KYH7z7EjmmrPtoK0uTprhKRWDaM6rkrTJGTfkD8Tg3keVa5NMH1a1
RhCjvQnk1hezFPkF26mPIfFQuR6KKkTakt/Lm7joegXJMqDzg2nyeyqiqUCRIYiS
ghlId0+Tuc2mF6WShxt9CYqQzhtFwIeAE8yPk3OfUqjdCPcTLZzccFOY3D8QcIT7
tMUmgaeVJqB5MPiep8w7zo7WAUPPOrrrO2LtIZB0RR2dJzozW27cFPs11d1KLitL
hbIKFJoqxxNK8idkVaQYkfUVE0ePlWiEI3+2ndgByfyGTPJGLoI6OAOC+vnPu7vQ
XtkosRwxZU6o93MrLihztrDiZnpmW+CYj1vJ8atr1q2KeRAASaKmWEv2J6+0XVO8
C4ctMFvAJbulVxqWfErmT+Szk1wl0n2VvD0WXIKknr1QM0rnz64+bq53yf02eOmq
8jo7W9P5DwvHjrsfA0HEE7tXiLhpgoXUZoV2Ay0A7GcexIQ2nruyXu1/OBy2Hr22
Rx8b5skqx4YEY1TXtzwiNR6wSwM3yMAw1SLNfkFS1GXDvDAf8rB5aHWGLIE5Ymrc
5/4v3urtmQVYFjA2zTpWkqchzBw4HqmeRjMDvgG4UuXha30xs8XgDEyzuVpZ4c5H
Na3Pft6Nzj5k+IR9iuFhnkivJKDHPP4lNpJNkSpwk6P76BuIDxnu/J4jQoHI7BP8
FR9uEGX8S6W10UaaI0C59rS3PULFx2ty2sKB2qMBTyrEwxwykx5ENMpytJAv7wCw
nXCw/1MI1VREGAW0lobDEj4z4j228VCdkAM7jalW1jRD9UWKi99KYVi1ZmGXuEBd
fJ8oHZDPCLXOpcSddIRLAYfXH9pYkOJW+eU/KexJ7xkrDvuM/+Jl9/jbGTrt2KK+
Mmm2lnAr7M6AaF2tYkYLaBsyFHEL9m0qNkoo0eTgEZnzeFK0T5e/HQS5FAeyIukW
G6Fcqi5xOKpgK3WTzvvzDYSxLJ8dNAUbXh0+a8aRRD4ULJKr0pUFTh8Jiqtt2irz
rWeYFKbvdTZEjfoWUg0NvUxHWhKCbo4SsaoEUIBs2uWqqv0ZDyiFQyqucha10LlH
/O65mJ8AtJXviNZsaTLdD5aha7dRNSTWVkngu8piDDXmXwAlTD6h+bLRtoBGgD3D
9qGLuWShcEOK8aaMrFmOgRc4zsHneyYlaEWcoLGIzqgM0o+YRb+Uz5exlPmjCUPW
wzi+Wqi/W7MlPS5iEr86kyMI/UysSZQLe5AYKVCG7CnpFTXl/hwCotjaA+C2ryxF
3NLXGfORLoe278Ujs7Jtp3f2YA9V8kJAKqwcdTQOf5f93aO+O/jWqjaQgfTOqH+k
wPFJhnKpZSLP8PgtT3elAKVev4BNU9TZBsSEyhelvwTMUGFtZiHhLoiAkrGgTJX5
6tAn3k3fgIQ2LTwqYRe1OGnB6/V8PSVou0oSuWYiOwV/flrFCxXMYwmrteSMNUOQ
G3fKuthVSazNuAiP4FKjbjPpQ7ONrBd5Ot8Xk1MUt/gZJf4tw4dMT+0UjUHyi5ld
iGzVWGPI4Jx2V9CbJrHYYt926WPKMPUE9/bhKUaRCZdWuWzgsejdPHRB/mg/DMCg
hjm4e7LlTJn7kkc+Acufgo00ogOwFq3fQnA6mYzTJENOcxy71MZO+sltFTtpr1RJ
oNBC9pC1lBPdTciYP4qGoP47x4iJwJnfXQKjH9/3roV0dqqU4QAUX+e5X3Le+XVj
DYxNp7byzVZhc5NJ0NayE9sQNhFH7hpCRNz64xJe3HkNWTIjPDQ+gdcvKOm/MWN0
3uMhOUx0dagA+jMl6RDxUGDU89oOJ8DQPFboc9T+7q8TftZDsvfDH1Fl36mdaqy0
jN2JGj1UOu8yg5qNDLj1Wtb05TRZhKjdXAkidrkbsZ+eaOP/qWW6yGM7pIlDHz8M
Uu0QAKk9z2LE2/vhbJmRWiXiSxgwm6FqT7kBSqRiHic6+lxZ6z5GZfIOHZc+NbJz
5cuhzQvzUp0HliBtu63aCou4AIPzav8eJaKaLVfbmavHjhgNQOUhr1+GfU9N++zf
DIH+9GYosDke1ovayGpQIM9xoZ9ojRT/5BgdGQ88wSSEpeXkRXmFsagWkykpE4CN
EHKhyQzVmNNmtuGnTf5Otu15wq/yG421aAcbB4a0Npf+9qGt17LykYROlAdsx49a
QEYrqD/IZ64CRr7u9RCAJsLVxOPkj4qSEptTaH2uCAUMFg7UmZPUc45TchszcV9m
UERFDeEYBH2WhSOrSvoLe7BpUvqLikS0zLaEkSVaSHclKdwVP/ItKdcRaKDG+64S
L1QTyiwn2uEc4ksFTEhrUumXNRH17AqHMET01NV6h4AQPuYZqfGGbmsBC5rjZAVz
FM32B4T3Uv0eizsYnV0ay5Xs8qOlzmpSn8CZtGdRQbv8sOB63a2O8aHbT6t24h9W
sqosSpGAEUPc2EXdvllNbB/AiPyBFUKLgVLPsfjVczJDOw2Zmh49LdoNSosHNQG3
N+fANTxggf0lLmhn6yhJ0WHRCQkcAzVQDluWHlxHZ/q692WGbFq/CH+HBBjwC7HG
SEDIbIIXe+Hpp4Gx5EFWM1ouofyVANrskwG5Uwuf7HPlC7OOmg+4uuroF1h8owX7
+BauegJyGnTC0UNI3YWLz5t6TWSh//7c5OMA4Db1hir7UNGB+p5db48lrtElcoVw
MLo/831AHWr1m65NbCpBwmAc6cKEfQkUI9tyBCkwAHRLq5RD7rgK3fs4QMqUfJnT
sKFLWDh8PSBer+cMiu3Tg9SR3bp5W++lB2DS3dhrRj+hiMBeBTXpG5LYOyN89BgA
LuyFE+767TZ/pCvXJcndM4+TlOkgxmYrIiddSLapN3U6NcsshL0pm57imQKGdMjH
uBF+WBSMBMWnLvyHlU6ZXwM3O++lh+Ie2ZRG9be6z8pAuKYdf4S6tB+RDVAemz4z
Dpfd2/9dUs/ZV+wEa5gtJlzpOyt4cKOrj1rED2flq9wPthr9RbY806FhKmi7AVlK
eYh9Q/i3HT/0kWRioFhqvzfilyFHKTyFFoyV44cDuzFBavSYdZvyta80CvC/6cZv
W5l/DAi48JpWpIbq+sCq4XzJapstkwS93z2ns5VOByKA4ZZ9LSa0MXNJXAtCUzQJ
yHf6+zjPam/jjfsFflp2NhDUqRh5h0B96bjoVEqHsD0k10bdrixkyiCzH6FX9cJU
HFZ/xTjkzjcWvREW/0K8aFBRC19RCW3WtR+5guQQoRR4s8AHHPtlEgXB5PClsF3i
nCUtxyGfaL8FFV+vHckeYBZ1qIbizYtXJdRrs/WxDSb9mVjj4JCjAasfEi+Lgx+N
eHiP6C9PWoe4PSWB3sh5zI1sgCZNcQU3PHIHmsS0tmzjkNhefrzkGNBvKYZ7g9Uk
giQqV427Vs8tIchviPJNslSHHvoXl/BfdvPOV8ektcqltMCrr5rzEifXeZCb+ec4
Pp7ZujiLDRjoX9yGqqhAe0+rvs+ljc1FZzFryGuHrtOi/ZmwDRbk+CringwIevQD
uLhCWXqZjxOUzCEeGXWw7F3H8lEtMARSPx/hGZvwZpa522W3FlTQ47xBLlWcWvcJ
7R5xt4QbXE5k4Lmytmy4PbmQbVLtUSm8t1fDmh9j4qx377SrQABosq+JbDQ+KSKu
e3LHypC0nLXQ6OsiZllBipDcNTE0njiuJW2GzYlf/Caw+GDrEyzRPDvlUVaF4NrB
aWTSfoVEv3Tc4haLVGn5Y+1mijhtYamvq7RtqmWgYZXu5rS/WgpAU6ghCgrdrH7d
S07mWzPHRr08CBqVNduIg5mRcHMPhp98J8tD+dw9Z51vI1esOO4LpxzfkISN54KV
YzrriS/HTmVWTOwdpuCbWgMbZnAD8jjJo+2+klDTnQCw78FLuaHOgMhtQ8k1Cnnn
8HGM/pc6uWRo164vfcAlS8lUaBI/dkVQnFCYtlT+m44JrfHVPzs494NfALeN6GJn
JwCYyeLm2I27f8Q3qngyyZfJng7JHVsQb3z0vAS7VKIMN6faquN0ZHjvRSz++o2o
7pd7JmVWJ84VbhZCBlZLbUFC1wVSfAxMoMYVRRdhCcEFymWW0UwPh8dQcdPVWPY6
URQQ8QuviFufdlU04b1B5GPm/BccC1/cr78DpgC4RiRak+wPymm5C/WBvX9SEPCq
NRtsw4fNom3fmKfn4yd9QGiGKqBkqiK6E07ubON3QDF+rjc/STWtTd/bc6O/PVVM
Z6QaqLWGPJWXre5dWQGiY6kImAiWXU0HEhgBC4diI/CDW4cRemM4pbcMg+Rl0MgD
mfDYKwUDzdbm1sdZpTOimd73b6Cb2vGamUBYXa+a0WPW1sehCyj/llX/z2tV7Vvs
X8HVQ08l35WcMNL+h3GtwLcsgTfgHcN1YrwFXv6G+ZuVYT3tA5fP01YHjJfaN15I
PEW/N0zHqGxS1UwzsYZuhT5hnNDVuWcPgJSsCbdVr5ZHnfWbZk+LP7M8wLtJ9QTf
LQnbmHqnkL4+20XfxjlNBDcohgiCiHmc0WIirycDG0Cfm0l4qKKInzlYeZp9KgQ4
jB7eLdIyp4mzC2BJcWdTFpFUwstDPCmuuStx5TwRgagQcawz7Xw96BzRROo61STk
nd0ZeirST5vhoNwUQ+Zu4gsXabGQg7umFXc1QtWBRkq2puQQDhK4+/bNWCKmffhk
/3InrJAoY00M1O7pAgZFOtd7Ol7sehrgZx8GvAmo2SI7Gecyvb9vwVRiVoDbZ6RU
ly0esCmzzEtNUlwpHHMoBU359lsc0v2e7nAtJLhB507i6sk/ut3l2Cp7dZslsPKE
j593VS26nejfTcHx2cPdVgyYWUYQ1hfTrnxjHJTZUnwMzyzQIqcKI5WeKlDooAbO
a4sk8NAn4sSDTmIPP6yuQZx28DCFzzVZ8HDvLyeOj5mvpKRtoJU+0SAYqI4uKL8b
cU/u5tHX+zY99RcIvgrm2YHZudlBFfUNN6AnbZRHpK98GXCa6YTeNVUFMovFiSqv
PqBEyCfQJuJJPoqwj5Afr9fqyNnVMkEBt2kVI8mIlZtRJCcE/IMNLHBbsnOhfxp1
sj5XwJ2zs4rlHF1qiiuPMpA4mtRY8Jz/ZR7DNtAq5GtIV+qA5Q9oulyYqes/PYMR
DISnH8xaQtNz5rGT94D3A+sOiCeRy5D46vwcJVUAM89yZHd/U7VDPNcfCe+pO+7j
txr7mrsMt6Vpet7m05/UY0kHY7lOyqHZXI0VVWpl7QdeHogQ19DbXrJ8e5IE9yrr
j62yU7TnEnm5JY0/F2bGlsB+yQYfVxlc8T02R/syj1Pfgog0TwKw0lgLZ8cU7SiA
1aE2ZaEZUAF26HeA5jxVhVMK0B64YcDBVjXwZ7YY+ShoKVOwR3A6X2hmFt2xHc9g
JFMYdz4/PUMbIRHI5Lg2yEi0r0UNIegZKhR1Csw02hdZFXJduN6ONtYFnDC9eFZB
/PC4kMDBMSBKhPIqh9d+ThcJxZlGj5/uo63jUzk/mVs4m+QB5VNwPWzY+8htDWf7
mNm15fZ4T+yBp9qsnnjSN3L4u/Y4wJkCEE4tm4zmHd4x5pPtMpdAbjZQAvVGsK+i
1noNZRDYZaKM3fHDY9R2NvD9NpxEWjRlO/VgIVHhiYeyeaWjx9NSulNqrnUPqUug
t9mj2XB08F/2sTJedtoRQ9RDaGPOmP8nrYLkvDh+XdzqPlJica+I5wTa8HuTjKMY
o6SCPy7MB1zch0S2Jsgjf8f6msuCdedhSdSqV5iHmPhYnnfXDICUT2EfCnLVjG3V
lLkTDHJyv7q7nDrWpa4CpVG4195QI9zlhlrznVfYqA/SbGRIZryvPgJtV92mXVBY
3QAdjMpAFpB5AhuqDcbrhE4KcJC4Fb+YTtQO5779VPqDzjmchwp1nCwFpaEsuC8A
/Qun+XNxK7mRe+x9n0cLWyOY9a+TXXjumnk7CKjzPlRqcRSmvNxIJfFATRkJNeSp
FuUOwgeUyuHJzd9rgHmpefdtXncEoL/LvrvVUso+8gn4JuhIXgSHPAkkYiinvnbo
i1oKq4kCxssJId9rb4icsOiMxZmFMOvO6e2tugjih0fpkKbdnqzCX1d+fGWcokY3
o4jKazXZG4K1QPW55nNM1FSwDUGkytHP+ilCRvhZHQPMEdXHPCqABpQdS0xj/QKT
yHo3GB+xbWCEnaktR5aif9JvD3KYPgeXbVOSnJtgqropNpxoo7c6bhmORmfRlbh4
Yq+QsyDarN+u6YJPAaePrjkyaRqvrDNGIxgsveytoy32dwnvWBuNYXaT1ziBCpPb
P7X7zFlvdP5gurmHV/motnrWIL4tGxdQ5KKzRVe6vCI5yiQH6WDf3COPmB5tRtQX
/9kv2vnWpJFV7Ev7rB38cPI7jJ4zaqpnS6AJ0wB/4mDBztdohslNTDqCpw6AiVHN
2h5GqRbN2WwQZyDm8pqPdMFcqKOVN8cNOHNEyvWrBGZsKrDYU681HZbQm2fsqDvl
vCiX+npQDKb5HBrviqEvdmj6ndCYcyEmcbxIb8tGa6Bj/Eqg6orxLBNf1wfBpEHe
oplD/USyTKWfsoqiHgcIHee4oKr7kkERO6PGaITe3gY2ZWJ58NYeNUN+OaTC+T2K
w1qtnYh1djk/OAi1764FxS117moE5sLVzY93XZ03os1OOgYIJHur6GM/XEhBCGqv
+1XGrOcnKlBEYMGnz+HhX+GoN0y7RwbaBT0+jzgUkiyiv1AzKToh+WJdEp92/eUb
+Wb7nsHxMMxRp1zOOrk4YR8g9tiQj9wEPOc7TV/l6qlsQU7EDquQpzI9esLnccag
nwXbWAeBwdrWyPDWh3m2n4kGqEaPVUfL6PmoO1N+zmPLDKlAgbktRhIO3qseFxYi
RQI0/t4K3iBVmHjuBmTRe6KEPlYq72PyDIblc0FB+7kli8Ji8+/e/DxzK7IHwZIm
RzSTmzkS4fpXmivr3+u3pz6KiA5xkFT6wEI1thU15Bxnlt1h3toWNTRI0lQCYs06
DjjYY5KBKTueRRL28LZiQDRJPhnh6t3iucixQvsz2McVisbd8Na9Y5DZL5p28qHJ
k3UxfgGFwV3ZNk8QgBwpEm4m1kmTaPGqYWvJjGhiK9pKWFGxQxu8O05ltxMRdfi7
aBc96CQciD7KSwYWwYwPHYW7YwMc4jN2SSIF1coveqHXTK1dAZyCELafskTT5CdG
yRKYdRzjO+JE0GNfuTprRW8IgNPdHaNyxO8pkbksK3XyPcdMyC1QI89/ZMLA5BwH
uUqYbq6AwzYabLX/3i3RXS8BrY52baF8TUzBbH/TySOLwd/aPxDf6LULQywl6SLs
HJAdT2chLRrQEmt9x1OCLnAP5tkS4VN0hy2yNgYBvFdpqA1lOpeWVr6/HaTqSOOe
UTcKqUP/tUpR2wARMnriMjrGBGPfOjGTdyIMZRfokzq3u2zQiHSPyskg7AP7JKjV
9VfPVyafuAVGjTl9o7J3aJUYEZqRlZTNoQgRjiPXSqiaOJ0YLdAYXqgpumnQlY+T
dHlh5O65iulJKK3GAZv15ElSbLHRkrOg3gI0QuZ83ysthhGzcQX27buJglnIaPk3
KY5WhIk+Ppq4AumiXg8qE9803Ee3mNrISmq9BYFrFZFRyjXEDr2Qgl4IFphjOdQo
1lwC7tYjL8kvDMobYyi+Mz0feBtwtURABHDaX0vcoPYlRHhzt79JMdTwFiqZmpdA
eohnCC0BOJRaRsBl+TYR24Iyvc1HgOsrWdVFVXb+EGMrsOYpDE/k/B8L4SlFgn4V
JtvcMsbiDwCImRu+jv6ArEEu7YXyakQRqizqQDM76UZbCcg6SF+Ar8pvUirCuxQQ
6TX0uDZUpoJ+EfXs8XuY0LLhG1EwsZReK9RWUv/k9yw4ILtLZqE9PT4HoGPoqsi/
nP4bStdlEvne4+R3C8w1O/nkTRRskORbQU/yLBPJFtVcasBSK4BOWPdA0I+7ZtLW
73Z8LzfwCToG6gjfnC57w3tKd1s9mQh7FECZGl1wy521kTbe34wbYQLLbF2XxghX
nrfurHRAyQJT5ltYmax917mmxt/0ysIdK2NBNeR+r3QqcsuyoE+u2S16lFjrAMOI
AaxOqblz0rLaegNsAranH0InMFbuD1VLb2flbP10BiK26nhCvFzyzH8LhB9W+0Eu
jctfKrBIVolmLHkGaou0Zu4OJgN1QSX8iYpqFq/OBsEa1S8lA75W5XI3nyrp6jTA
9reciGxVTL1VwthkHEEZINFTFtFa85DTuVGKk+p6a0VV0UTnJp4W2EexD+Tzvkcx
jMiFM46KCGR5GrXJA0FoAQrCZRM4S2ypnqN7+io0FN9b6rGc5HU7mi3X2XRTilfJ
2PklkTNeVDONDNK13qXG2eEtFeQwvUX8iZofCpSPla1GjFk9PK6dL809jL0YDgpK
ryuS4KI8Kf/6dHxNGbRsjg3Bvt5sQm88DwxwEBLi4bqH1zmtKwRKuX9k4jS5IU1Q
ne1oOgZWcMu+D6xlv9BRLcAKhoxTP0lReIeP02ybvM2iAZrIfgF40MjqZPWFK/sq
yYKhaWj88AWd1KEvlDejrDEd8Z9u/7JbDMdl48XYcwvu8yUZQPmFzd3WbcufRQuh
Iu93QEIYXLx4xUUWFFktn3Q6PjyUWKp/qpnLe9xkhkYtuIeZsZEAimALuB8bpMSt
GTRYbOC5IRCSt7IsyYmpO74j5T09XlXcm+lfdPowCQMHLnWd8PFRkToDoSZTPL9P
0Zs99XIE/EES20/znHoHYb1mdZMb0LFUWSn4Xn+QL/wGcbCe2S5W21b8PU0waUqf
wtzWwWo4OYkUhoEx+oefjQvPd6wH1ezz4yIUmQTkCNPtGLsirUpQHExrrZnXu+BC
ignThuc0tPXuPrlzwL6BQFfGxfxiCS5RpP3LMVHUnesfDIlSFluz5n+8qhImA5P9
Jx6LZQXfv4oypi8OWeaw0Lk2d7KLSrzcUelRWtWK9gvwVh5rHSVcnQfxYF1C1UhM
rqHVX9q32Ts+5tocn4tkXDiSmMRYy+xWt7MGpbxaWRQDIg7IS7BixlRHpqo4Yorf
2r57hzOxakzL1LzdLEKLZXZ+eJIQ+K6XEkh7kJjmzQZeiVftzRc/cJmHgyw2AnVm
/2+ExVTx9mlbzDybTj2hnWl2BaqSsXjiQfh5VusYvBhtnyGUioAnhAy3yVL1Nd+U
HKqRqmxlO9DIyenasUj0E2NtI9mM8HRPchpJwlN11b/jyhxjjNrzUF+jiCaUvldc
3nHbZODTaybCSGjOLZ2jqXnuHdqELzfvREpyqP5z4n0ei+OkjhYoXj574YpsWlZw
3VdCw4TOKWPVe6EMsYGFq24ffU/i/SxlrqnksvSDjJLY8pK2aqw2Awj2dwlmpVrI
21w+W4tcvmM91v/oP//Id+RLxEN9/Sm1TPzENPU3FYaD1f+6AioPA5zpMebgzmM9
4PRkQfxONZSs85R8djzp9qwGWde6tsoYzrgEcyVvQMw6jL7tM+tv9Z7C07+Bdppe
uj0msPyQ+PbpS58qcrOFoe4gBhNj3l7PkQltyUsn0JH/yq2F8U7+NUa+/Eesvfhg
al29Aix1RTyN+UodNAU7qTFnX9rUtDJLf6a6aAXyY8kYXSPgjieztCR/kY2O9gOn
SqN2KxlEoNb9qlRS+eCfoGjBNSo3H/wrc4UCj81aAQf1gfljAcefipCcQngnFezh
39Ez4qgtLMkrU/8w4L1/dIJSVdPYxQjx1Y6cJ3heO2EI0+wHUWKj4Uk+rQc4wEO5
ofpy4KDPxnB665w9rRX5wY9D2GZ31Ynhw1GMo9acXIPDVYtiofGARJ0cFmDJAyf5
YKcsXGG8uD7RR6upUJYlYUr2CjXIMsFOngeZ4DYQNW21V45I6FTYw+ENMAr6s/xG
lbyFPcokyz5PLQO2ySgN/KN2Mjh6UZWgFn9YNxXbyUZCTRt6aAIa7c+M5OPhi/pY
oAhhphu0NgL967TgNAt8mEYwKv507ZpPHAzy+mAszzwIodcKtgpXIYdnjhlMxhgR
bjeJI/Mgqx58NPLyQz92tQqtIye6X0yMDCMYnNgjDgXVSD34tBjT0sLYJQb/9mWG
CJjyD2uvyguzV85OqF+6JiU9PGd9ilPEAuSl11HazFATNQ4G/1FPxX+1gkOnDxrZ
zVzZQZykXr5hX7OyuakwlnMBKlw8WNUjxjNL3xPxp/Ynj+gW91BjOtv9BqSLNZJF
R9CUHA/dCBZ5M4OBHEICmycqFzeZQNvHWJNpzMyRogzBmjenhGf38rvVxHvbuP8Q
iygdypzap2LLN+bakoBnMYRT38sL2lbFYdVxN2nCV3If0rFZ8dqNiIfl1apfpSy7
TfjW4QxMYzEpBvy3EWpWtF1xDpWSejVhs9hf6R/4xnocpCI0379yAPclYqRt8FDG
55YJOJM1xdVryUViPC6RTeVF1BLaNSFZ3ztx9MjZ4bvbag0keA2erTi5Z8CnEBvW
rTNXGhzq9WZhwT2GJb7ZePkiwGlj9ncqSkdylkzozdMwbw+U4eYjAvk6EJemyes1
2MisAnwd8Kmhs9sc95ziZoDNoK/h16HFqHTRWb4nLNSEi+3UU26DXOowLvwGmssu
D+B9aa7VDp2m1YRgkJ9ygzKJYv7qyjhPNrpOmKbUsHKP70OifFUJCFta9Se4HQY4
fVrSRkxST8jp66aAiFcrYrTicIeiTXjKMXt4h6Jw7XTHiNlpY17MXTlyUM/8ZxvU
gYjsW7eFG7GTzC0X246mOr/0hN6DQTO039Uam1deONeJYHhhizitXgeV8wQ9QrYv
gzOLWjMZkDAcE/DyIHdavCV5mrGtpPwprDy67SkRXNrwaX0PPb5OEmTr+E6hHOc5
ME1a05HUl3XgYN9YuFl8Gyn5GP4Y09aDd2Xw86ODI8Ew5zECEZMELVCOhCJoS5J0
8B/6/Zhfke6w2eOfkl/ZCPXXsFdcAw6DhWm0b/FHKou0mdW+HZW5IKZke/RDv4nn
QKkvMquxx7GZLqSKJo6dGHJ7bAvWxTcFGRK4nZIAhdkXUs/Fy80KCnC/Y+tOSKPl
8S2VpBtU3smS36LRjHqLV0Y4YcEG+5SC6SkY91JOrzMGG/HnESy9rmUI0grQZ1VQ
AgJEV5KuvxFW9M6ZBv/D77OONGCy77tf53Z5i/IBeYvd1kwRjaqgSneKeBti74Rl
OFGR+HBN79mwonzSjnM09JzbVWP6LtCtLQH5dbhfY9mcFQ6iadtniucCCvateCqI
a+wqzpaUge03ZbD2tI8sUqsUlLhggd+Z0KSO0lMVbceU+Rq3QMeBQ/3pxumiy4tz
qYI3wqAk+N3IwIC7OSogRP0FGDaaf2qxUnCK2ggyu3ENDvVSICbRWEWV9Exe7uEY
1nEAgFj6ploAjsVp2nqPCHsgXF4KnTRFtQpLUMMvc5pEO+R5N5j202BOZZY5ib4X
9ikQt279lZl0c3a9xiYakH1Yj+Mzr9srrnZRJVxbsmo85MPMjsGPHrYt44AC0DWy
nWV5okSPI82OidDwnXEVv/pi2RGIfeani4YlT/sqXWQEK60Kxg2iTo/BnU+I2dZX
iGHycY/XpmOhs9zGHR+B9ttXHBkAPzlNURvmyri1ZgVtil+ROc7drNSqNRDFEmrY
fkMnwDlbHfEWaowC8ogTyudfLws2lIifLyPpP4BqlzDB4ehCvW73O28aUVzmudAn
P4CgiEH1wOXALfcCnUDYuE177Se0xH5iRfAJx0pFkRy2vPmVR8rq8VU/tUNpfViv
vkSeqSDzN1FJzM/RzCo4GiD50k3VTZCBRCQkGH90cuchIpSRam9Ets9IOf/XOAtH
lRi6fUio55nsA6EdSIAmZSA58ezqmQnAEryep8RH8B0lzcPuhxwm+fXrSNQHBm9x
OzcxMcnvxLb46OFau3+rmbAJ427Ev0/BZeszUwkKmAAHhk0A912BAPFzlX4YtYgB
klOQCkI9f6gboh2gkAU7KM0xKldlJ6RtY4fv8E+QEcv+t7elu4KTvmz5owvXf85n
V6e4/j4VkxQQTdiHWLtejHq0mAyuK183SrPs45yjEmOz1kOaVoMKX/3/QWZLLxls
7nSPqriWl10OGhfCliPKrJ0AyI+nWagAVOJ74d+MOIS679ZjMwJOIod6JNBKyroq
yhbfv6tceCF5Qs34bcJZZAa9lIR54cC8BHYrSAHAFL6xfXZysKFi9ZBVUnOcGMEY
nVbiFuKm6ZzGhhsvOhqRWNzoaCeH3IZHjspZPCzfWZ1x+CGiX+6Nw+/uVpKvoQwa
jgCQPVTQW5EHY3qu1bUh/JjVT+xAVPyjsDKaxkYMmxOmXWo5X+ztEk1Od5dga+id
ljoIruwftn69QenUXXrmdDoIUew/JBQmF1MyLe4v/KyhAaFwzmGNX+8sDWOZaw4/
QllIvAmPjrIe7VyFnsN/WhWm63/KsM9CdaCrAdiqiR0DfOZwzUD45QkNHq34rWhQ
s8Vxu75cZSg7pe9arCHUYS3W+t62/UWRNhzMujEBwazrWtaMylCX4vlUH5kpHI3K
3j2u2H8ftDXElKCi4AEzTTX4iWcxfxm8RDGCuzZuKGfR/e00K/SnbwXhEIYLSxgw
W6SU+tP6S6Uc2xkimHi/x0z0ZQAHIESXgMU0qC/aJtyhAw7FuauIemsNsNBXRmvX
umE9WBhZsAZa9I5sR/pbBB8MXNatxNiZa0dswPQMPzGKWoB2Lh5v9knshy9q3JEH
GlXnBUNhOUJlBwNT5HQ9vsYrqwbBt7IM6Mz4ttts2ApkPU6B/Lm0gzNDm6VOkIIS
yM1zAQ0wtGAxpOgzLDgfhNhD3zp9iHRZzT1pg0v5dyCXoucojvaoozjJNGr6W4l3
018875baizkLz9CgdxsXqDng0pPIWNfp/hjYp7KrXPcKPlXT8xW3XrJ1J4HopxSD
+KIuJUsaDNBgAadAMBLZ9ki2mQK6k4H8dIRw2yOyk/LMpIlyieH4GggR1JQN0rGt
MjSB8SzB6E129FBj5MwSISJ72jpd8qCwdlMzCtApgKijTomKxE/nhWkEQ+i6UzeI
f2IL5vxbQ0XiRh06x87vvLoPdjz7SeUydnhB1fmU6C6EsorRh3zzXpI6S9AfNbAi
AtrNgzNN5R8KMgZjoRHt86P1OxtAW/WYeT3wzCLkTRUYh8EqAbvR7TZYcC0uwlPB
8bflQLivOhN/wa0z03FQwv1t+Vt/WIVYaeO79IFsyoliXTKvKG+uR612xH8Dx2n2
XVRaF6fpc8FbMlthIqJp0YKXVx20yjeVup9n0hBJmcnPYQdlxaQ9p9yPn838KAzQ
scKDd04Jh/g0urOh6lZRK4P4DP1Z7u4P0dLBSc32MXUWfKgzdBqPTwbnwJn7qkd5
wrOlkPW8z5JCjewbzbkEnaeMkzT3ocd2AuoJAqkOxBrrEqaxyzVv+V1MlszMcpTZ
o0ez/UFE+mJtYGNguWFffdKq9Iy7QFz9SffgjgPQ4LSkOR6L5QONRqGVIhwqq2mq
4VdqOc/N6vRQvZmwVa/anBt9fh1mmRxQncnq4UQ9ecuvmwR+nDM1EonGGT2rDg9k
VKZeuTJW96UCpjU6K9iUyN3PWyC9/XiTcmWITUnfDNzv0WN/kffwF+9QNenrJeRe
jlvMkz7BJxqzVvU5imJa0W7fvibjnPVCjXRplgoBHgA9xuuhWByudFr5HIclxcJf
yKj54GIc3IczON2PRNAbo3Tki3PYy1aibPP8DvuAc5y8oJu+f6Yz97QvdQ+Pw8du
atIkW9oJTZP1Gyovj8ADvEHkLCltZro7lQT0dr3uyzG0cTBOoGBh7Omt75STG27C
kLHJ8MG1DAb0LIn0lAz7VxtOXYThi//KWPY5j0HfPgHZ+Isel3Gf4enU5yM6NEib
BJxNavNAcS1lHne7ipklgI/N/6ENP32KhNaeIEX2HJ6zNqyU2TY+gxTZZWnl2UVL
M9IbytOL8MbC32TQfSpYkMIDch6uWx9xVE02m1q/cW9UG/27GrIn9LwewSTYkVHj
b+o9cFObU9oenllgNwyN2/pWehUqvtPXmOMOfaqLRYRNab8YZ/A4eHxyrq7r5C21
KfByfNjyVOy83emwy5mvr+xZHOTomaDFJMmvi4iZ4LOGWmjuVoEa7ikSBfvbA/Fd
YJ0utEVqpmz9lJ5CZivi6UZi0zfNQZeTCmURD0g04kwcYuSzvF0gP+XvMkCjL7pi
prwApZgF1tljUfmecdIkO71DRObCuzAIpnH3zY1Fnmt2rzTbKSscADPA4sAHWbGa
ZU5fUWTySoXbcG2IG4f0HynbwLKWHOHcfrWJDMn/nkWTB3w/Pc4Vr2cErtwwG7/n
xkVvGe7UMGfjO7NS/s4uA5aGwr+HrbXi9q+RXiW7FrtvlIYiG1sIzD0HHf2pvJOP
VcJ8YcucA6/TLuAQJSJr1Dw8ZQZ4rtvM1HB0z3BNDCC+4c/y0h5PKKJipUNxmc2x
oAp4aiyt0e+MgeFruQ4bLvBo848PXFP7bo/r7SAXH0TUxWsmq5PNNQdqvKIUrIvg
DXm4goazF+4JL81JTv0xm9CGYURuMXM0naCRFOkeumk5HOJGURERBdqlCA2wm78N
s9YvrkGTCrsueJSJcuHZGDdS3Ajz6ON6AXRiUcLsu8taIrXPZBc14T1SUOQdnXaF
DtnQgtJeQjCsAMGuwBt0wT1FA088vf3QzLVqTRoeEiTh8wfdBG9e3/zXlsq6dxnx
yULb0IqzAhL6LSuW8orjLzFk3jQEj2Fk29c/RAdAIwrtTlZSgux/OGt/TyLzm+sh
UQHn+weNFNbgZg9X8VSR8I9qr+xyiaFBCi9LBJFz+8BuOkVTO+x//pQ1RvYSo3ED
d8vEc38nbqjB1DS6nkpV0hiw7SCdD2eP8ZOxTCEgHIvuyDqYPuNZqAGt6MqzUcGN
xxSLlcywAp7VzUpoTRLk8cHe3QAoGE/2Y9Kzoo1o0MeMrfscd+XoOAWrpQ0de1u3
qKFQ6ytPF2uxpGfkPunXnG6paiKwhmFS3TVNvyq3gwjjIPxXg8lx/csxN6Cb1mxY
icbGe9UxHYroz4N+6GYxfL13s9Ns7d8m/gGfsWZI761dtcPdJwAlIT+NTni4N3sr
gey9iRdQulCbEXMTOuAhsEA0sZ4WNsGjlmrf9p/7/mk5r4h5D4ppL7/uq70iUqoV
VyPThX2VqOxttydb6zF6GwGJny0nXfwrbIhbrnVhPAX3PBvs6nSc8MYV/JKghVpd
JCsL6zV2FRn4nmbvQVdHBzhj5MZh5ECTH7m/8kl8sathmITNS+DqNm60FCCKSAhc
BK0A5ysSUaPAeAabKqbceod7310YHR30KxXyW3AedWMlcTHYmkgy0ok5h2XhOFFH
nUMAbaxjZvxBBFl7cG+1jIv3hUX3zYwYrXorg/vzMqH1sVwO1au7Q5FmQ5J+uLj6
tJnA9+d/axCzUG31/dvW3jPj11Iq7FShg2idLQQioiKn6X4czVmYF7nQA4jhmMAj
FMbW0JfeAwZJJyjI2rPU0ooUL4gDdbyVcaLiQmxD7eSTGvfkmp+apnBjsA3+MYwf
/PPg+84OPY6SWtGfMvSNI/0w5Dz6eUgPFuxqVQQbSrbIP0tJexyMGR24iQLwYQeq
2332YS7s4HckIF+PWjR2pttxx1pxXBMbu70/s0NTaDPSyhkTdAjJQUPTR0XMX4S4
AvLnsgxyQMwTLLUMO7CLm5mxNvOsC776lURGkp5Pbt0T4y8xmJsBRvL2Fq+FCER3
5o2OKCyOaUD7VTfTp6YcvXCC9/P/UKu02FCASIOmU5iT9nKcv1hXa3/0h7FHY/eV
RZBfYXMCWI4tmeZiMwzBYsDS/LrtID1Xw6JCzobZmbxyajt2gK63QVAgcxUWtf8s
XDip76Vh3NXaPn7cUTniGvJYDLYAHGZbAN/FX6KrSRHDn9ra5K58NmUENLff7rSP
nFleo2ZFLb5hYrwjRSsvv1m14c+MqnOuvnskirtjDEUCKi8FpIcD498IuZPkpnCY
WAbcw1TnXOS9KJPJgSH7tPS8oEToi5QTSdHkdtmITnsQ+xx/Emmo4mCIyM9E3TAY
moYivTTvZGQxWbe5RifntBaT4BvTuTG5x8pLe42UZzWkhVeinN63ClLo9tKPbBBf
oMPIZnLq5bi5kARDmX4niZVfPFwxj11drAPzcLADVWq0DkNLE2Ok9n/L0UVuzvfQ
BwfCm9mwKV2RqKuwG0Wy9RztKtl3mDUxngvGXFFhhaRik64c/HTFsnL4Q5T9gCQE
0mg+q0aKEFyJe4+EcNWxYW8/9sF2i3LvutSRUd1LZTwuELuGwaTjOr4jV2SwnIQF
tE0i4dk9LYVacP+OqDdLHSnr+MELEShPv2frfiZdIwbYrmtKk+OHKbD77YlWGT/3
xLZ82vBlfT/czwZMsIWTfr47nMR+B1kPihYf1ekdRXOoE9zek14wRQX3RhhxIoQq
SGL0KH0NlfqyGW1ra7kgq6sDuf8ElqH+JBik0MD/AKG8xTa3YCORXIsDZjoWgdJc
K3PCfF2IFn02ClcZDOikoE8+Re9C9aQ53sbdom+jFJGMlAIA7DpRh4Wc5OhvHO+Z
QBmyf60y3uAz6wknHetJRRyY/cnNTM90OwfKKUuII0cUTZTZ8y1Zoh7jiTKqS6MU
MpmLA+PSCILEmVN7S1XcPMsRoXF8321E6/mInGssvna2s/b2L8rBo4RS2MB+g9cS
xJSQPl3E7yRKfaefiGo6eY5xz90McAx+EtV9dVn3Nj35bBbHijsCBe1lrvOxMWzm
Hu+WxJ72c5k4F6aKqUz1ag+7r75BoKRm6df2UYiqrZqd4MtMipDBa+Z9tUMOVx3g
JY48C5tg1eR0GO78EOMtJb4E71DpE50LRBAK2UlhsOpN/OVoYvqmpNLvf81Jrh2K
cS62vISjYvHsiD1+/E7X+BblAyU3NDoH4aRIzHono2bz2STMmlKcNMb9O/sYjqbm
diRoF4EteAJG1d+v1D2r5VPCZaYg67n98zfdZ1q9lCiyu6BW+FT5UejInVsTpJOl
/d7ucO6jJ14e8oRXHlVBag2vjGh2CWTOl7PCNWWmfv2M4AI109BGWPMIizJrODS5
BITnXKhukwdr6wRI5m/buDC7zNoUg6QWMN3AE7wNRWTFWJNEjM1SDGbMqI3OTf/C
PglGAi6+oh21fi/AxGq8bjEVHSltDOWEZsPGDjFjuvyTCHmqDZ/+U5DcbNZUOunc
xtmzg51RLETEOYJqQS6Rz9Qz5wkHDpaWih3iY8oPRtZsD+ZDZBfaqDdNS5W023g6
9SVeoNt1llRNHk0ae2yJxQYbqHkDEtWLzb5bQlHISx8gvg+TXw5O/5BrsAsF8DR2
iyxcc49TFwvH1wMmDYMA/2iBIr+Id7BRhxGIApEz7Qaphd59E0C0Pta3KS2DeCUX
P2xWNeQ5PTDiYibuAXS8qYChzeqQNxxbnNsspD/l+IMbAfEUjkR1whQzgbkZtnMu
ohizC2tG04lVzIzwZwYr3nCp+P3tu5wi4egoIBdzVLTFgmGqlwmVV36MSmP7XGMg
Qlc26Qk8wqZRQ2EUWfDnMy14IerZJefvN0yNTVeRIhl8nk8NLoJJ1Xs+/3NHWo6c
+I1C8N6Li1TxffApNlmg5NXV0weCpylIBmW7aOpqpJNi5YqtPtHGa91MsqMtB/+I
voieub1QmYSEkeYLkENm4T3/+dpPI0f0OF+M/w/rLJIraQFBvWGaoDGANuFgu/rd
ted689Wa2JM0myPcOTQ5NIJghYZ94KbR99opNtJ9zrSkJmfvQIIJsC02DiGFrxrU
X7SmQ2tMROrdrLiLiaZI9ozolpkqbfSA9bNLP7exzqezdHT9kqQDfQ1jMc2PEvaG
uIUw96XVvTYNXyaoQyBUpGMZQj8CQEkdSMj9Hph69SiSZqTYOXxohYTOII9piNsE
pCnyRegR8oRw8IIVp6Q68ofXADmUT4rRjQ1BA824rdG3mkVSyXjor+YMXXffax4u
jU6vBietjjsNhPdHfPzcgS9Jc5wLMz+EJPs6KFvLr/fsuyriNDh2nvidRBUoBpmy
j7BwjIQANTDgmWY6n9KPshW15bLFKbwx2Nlu0tvG1WBMaYChYnMlzHEHXwM12EkH
0mIfJEcg3Qfq84NVzRmpZIAih6tA4XDZxO3Iuegt3WSbMSJNrHwVqa6QteuylcGa
U6hvR1XZijRZ+jl5tJpeEVXgb+M+7KoYWJV3eIAg9H890UTi9/yW+e1AUQoRKA/W
3aK5CUysL5DpB0jpaaoshswC1jAXLKUporhMT57fI9WW7LSo+OYI+9ZM6oLRdV0a
BhdpZRltpEiBhd6xBoERt9NXt1QKCMO6or0kulPUFJ2wCB5t2popjcJ9TNFqK2EC
HMDdHZR6E3P6tKAkywxtGkrb8bwgF9V2O/8UeyM+FDBLdK8WtMNPpnIURqkiAWmR
2raTlWFGhr+nmH26m9d/uGsW9hVtZqlRWx6AdVa547FAUFH7b2oY1LLiW3eQXjYM
CXf618YM/PlDoXkssCTIJjUWXICDFP4pFzlXYdTy+5IMp7qw5bIhCOHU9dDW/PXK
osYJ3+OTs+6D4Lrdi09cpVvzRYD+WlL71iuzuLjsbZo4mKdkVloGuKobTo4P5Lxr
0uOAJzbMz3vVMmDMcblmBRFjEDtq8yRFSn7LXdcHx/ru8waycjCbmA8BbMBL43cz
/ZHGsXKTavYwkAFuzvl7pvZ4gSO0xFRBphRnouCzZYYEXAfmJHTrTjua6Xeqz8T/
Vu3ZjHvVQ2jyjmmgXCECMfLdyI9AWbCxtIW0zvubLdjOlF3z1S2h83XSb4lh/Z1f
bzjEwuy7NnXYp9nRiPadeeC6cacNmj3xBwkhzjLPVytKZXWdbM+nBpBksIrdsqnB
0n8FKkvTM5cdtWY0YaVwPgX5xxBXZyDjozH1oEtICfMt3ex6qQ0xBMNlvc3F+tu2
64eDP1uDBJhsqNRxWUYwnhDC4ItK0Ajfy05z8z+StgAoz79dXywi51hIqTF970fv
dJhhZkqOEeOSSjguvqEpBEkfgZqvcICvbxm3hXyU41uLWljigOI1B9qgVWD92f/F
hxATr+zcVBYb9tRPPJ0xHjjZ5JWINlUOgJW5B7vaicuudDsXjDVaHbp6N4TPOJOr
x/1JoxqfLmLRVoYvvIRGtYMlbGUWvSPy6jYGf5LuhQ80U9HkTrhTAOYtPVT9k9bL
1PFFHZeI5944PM0X7yd4DhsdJELFuA4iiOV5Ht+ObpUNDSYqN257XRHh/g1urG2T
0ps59o5ix0K6cZiLvusxIbOf9/bzee1NJw4lnG9H7NIkaLdd0JHlkGtrrRfAMA7c
XGZQCZQFi70dSGvmH7m5CidZym58fcr9lkO762nUQ1qdQkyl6hYxk35pqpny65Xx
x8k/esrGRgnxJ0djgxd/aD6sm65GDX/720fDk1TCY55ZblKsGfR7PsCHyOeR2rEq
fGXn6FH9HQsb54Z4jgWWHrj28VOEnAb9wUVqoA6uT/ZjLikW4XT7I1BB49IrSrsj
ywu6tyIZAHsiGyX5KtVbvb04zewvjEsnh8ipekUplGwHxIihz+MNJKbbKvCXviWl
PPFrpYFN/4nESod19GBfT/zZ2PE2aQQ/4OfW545wNhwPV4tqh6nZQccC972R3gaZ
JXLjNyA/V9KBlcZ+mqEWiTyfbC5ttTops3RHtDY45+lhiCWF42zZzSRNAZ+FOkza
lfSeJ14NAyzLWIXidt3l/jjKE1I+D5NwkqyDnfv5ZPliZPxa797vx8xvo4+Csq+L
6uEQLhxrEaynHrmomT7tom7kb0KWvutI10Yr1JmaEPBedETyYNk6MzIsgrZpJMNp
sHpJqawsHUhmVAgxetn7HkNf2H2aBksHESa/iTFx5FS3AwfrIss/bcEKeNIis9xG
SPmnoLDnj1T/PWL4sEY8Rp+5BrmJ5ubFyu9FSwLTStrxtp4omAZJTZQ2QB5bUnp1
ESRS4APDVvWLZXW+yJlfgUBg/njbVnfPjpKlGzg4OJQ/C7bqaVQgOI5QLxYa6Kwe
Wf1sDJ7ng48PhP53nOuMc2YNwtfGwmB8tYZh2upDGPDrZBiPgiLQp9B9gDmMDqMQ
Gqhhwvhv1mF3FNhT2pTjG3aS2Sc1jbpp8j+es+CN9+7p0/qNPQpTqa3hhD7J2s8H
P5daGG2gVl7U0fsilkJAJqVLzRAzreyFwT86vKIRt282tJxJc6+5Mrga2PFM4rHl
cMx/WDJzM8/p3JZt1vKe3lxwWyKuNlPqQNviP4SY0xj4Kq7SwOa915Hcwbjq37xj
FwQOWHbUcvPlpCYv6ff+ltiekNMiyfa5Zx8R7ZiF9AosLi15Y0A1/mc2E8jl/u16
uuw6hb8rdUDjA7B5r0UAzhRmu3fG7En4S4szgoh9Ldt2IFHftZ4yILZfUsNVeDyf
Scr7xb1or+hk1ZeUuMyvaVoX4TSdlC0S/oDCoDgQu6JFQkuQOyPg9xZn1082RguW
gQ5FLL7wIsaRWlCTFpBL/nGehkTTTzHqacstVe11eIL+03zcj2mrrZBePR29u4hm
+r1bXLz/lV2Cl4EdVjEEfFoeSd/LAGnz1n4mHGaO03rxyc1vztoFLEh6Insrfp1M
YAAKDt5h/F3LDZe/VBnffxr4VznR0s3rBeRZaE5n6nOG4ndod3D5qnoGqUfg0lWv
JwLJYkxJVfRCeBuAzU+NEQkXPz7Wa528JrOkCv7OAYKpOWvDFiwokRozkjR13sVg
tP26Zr0CGXBem+t3xWCGvrm9y9nCPr8H0N2bivypHTsp0JusWLrOzaDkGsooTv0U
8wPJftrdMD7e7MNRjVCd+WNJrOFDT2zEOhKs7Z5IsxCWYuilMGvr4tjqGRKu1iPb
r9sbXOtnhhVRuQwPtiSPawQbAI8MgUTblIthFIQooSJcfZxcr3RG9KGfXZ8Hg/Bz
90IoEUcZI3jydbGVyQXrYdISQybLR7k2D2lP4cZ9QSSI6vRnXHJ6+7XvNDG1kmtJ
CptaMn0Mb7CEDvIBp8UYyrhqNw8dq0PR3frwW8fC6d/Bku4w6I8cwy+pt6R/dkwm
ZXHgiO1xYF0iNLfArUmeHFXkqIudNWSmFEiQQta76xU4GtCsAJ/1r3HkOJCddInd
t8XaFQEjdfeBlODNAy4iv+N/5dSBtB0jwCtOOaZdmX3WAtoo8TG0H0TNrQfDnVX4
DP7eED376Zsdha1M1iRam0XrVAtd1hyuNfGIKGtllCTI1jXrQdw0EL+tgbhqOlqI
1t+iyaxoDZsWV1AXRH5zjx1zM2uWRAePWtEsq0j43nVPNhgVcJ1N1nkhCywKg62F
rKi56YNSDKEEDTojGcO3EH0bVX+WS9gVjL0zDe3M8iSgDodxRHGrc5NQNxZjiZV3
jBl+98FSiaQ3KFjmCyx80tpLLKdO0iy+pDPLtDDWKG4ZnLoPCe9pXGZxy0NoqHzg
EInR8lsgls4ZAtZgHzkAGr6Hh6wX1U9Dn47vPx54u1TVe18ZMfSVm4MtEKLVc5m7
oM7K6ih3lRXRpvx6C78J4WKkTK9WEHtCSwiqH4Rnf+reLw/0ZS/zFV7QVKjL34cN
IlJSjYXnYlgmWxNTs/MYMtK01LJqy6ht4DG2lBw7aWn8sUc5LlNsv7AlG/8v5XKc
+g3ZmZ0uqVN4YeEOxz87QzRksTKLF+l+AZ2deKJGQfcaQNxKd9oyRI62Ic2vrDXy
tTyZmhCCgIgXArN1CFTYmrNF7P+6TeW4SPajepnDxn8SUfedb2VkDfZc+j6LpmGR
3SzUtJzgrF9uEWCjiuHFVzzTNjjVyNJzb3CkuElPRVilGQdlFxVlK6ZcBG1qgyWx
mwXOkbEhGQ5TEAypaFCS6XsD8hSLJJW+185LgZWvk2kua4xmMKgGUX+7iwJ8a6kD
JTUXfCC7pG1rynfdzeq+KivdPDzY21UJL4Hfa0xgkobNvf65+IDBtCDYLOOUiUnC
0tVtpHgTGdv0EhiGhTbHpXC1LoRKgWL48fXeQolGAE10xQNFvuyvzHgrWV7OuIyg
+OPDLg8d2bElUq6vqbILg8wx3j4Q3Skrt31hAgytQAoLg8CVRtcAa19I3GTrz75N
Mkpd0xDeTydgAa1cDUtLHJjzbnhg+cHM9g0f5A3LjSHpoQhGNW7GhgV96rP0f7Tk
Eb64K/vhj8SWgh1kw7fSYsW8iJJN6tk/ALmozDYlPdMXmRGAthbmcAfxfI6Aqvd7
8Hha50E4JNZOxDeGd1Ac0G+helIlwEBtsdTciW+F7oNzBystwH+IrxCQjcNVWmND
eb370xR9VuoEYxm1108nMruHYpVINXPqDOnHdp8txHNnhhrpxZqLc+syjDB1/fqC
FUxt4vXFR/FoMSeywreciGcbhF44WtTagWUkw+UW4hMwtgV1GhqsivGnyTiQpYPM
UJjFdRXw8VHJIaaauL9eEz9iUz/PwV/gyEzgybQwKcHanisNCrnYi/R9JdUvRFOv
w+Iq2Ahd4FKoKjOIuI1CR9/djoLCaAm4jbcevD+D9PdZVPP+wDu+GCl7pSUt92V2
m5WhK9MytL9p6C8J2+plIz4h6Bbc1Jp6qj5m2xAE73+smhh8d36dzTWi4BFrmqAe
do+4butEjUgJz7gsGChrcq4bDD/e/rwBfKQGJopZuVGG7xSI0sEFdH2fWdKDv2ez
0uF4b9GF50ptbhRRrVXnrMRk4KJwCcMI9zczcClDFi/Z04nSctkRJ59+d/o+S3ff
ePkpfx8s50tuR4WBPif9ArN0k7CWH4eEgQVHDijLXblB0f59aBohONwimPw684NM
g286wSpQBsVGPdUjR/JGkW5PsWfMTzUjqs3auY6cpOQWZnC8uVC+Yl/1h2r9Jhfj
fulE8KCtw0AOOgIncX633WYha1985M/nsyc6CJ6qVgOlvBY6ImmtiBnDfpH1NW8L
tArxwxvpkCJIE69CoJItU8BxSR2seEBAieksewckPl2fhPt+JSjKdMBdNNAj9WQC
cASc6ut3TSSlBqFPl4r0eISXmSx3IIFfFt+VgGwJGkI8BiBluO0WijFZRvdbg5xI
6XDCOOSkoQhdoD2+2xmPcIrlvx0h7UDDlmdk4dUH+sd7iO/1lAJ6SGU9zC+WK5CL
LXVJ3mOf07ubS8XzVCM37MkpqHcSJBNAffg80Ih5q3vll6FM9TlFbUA17lwXehJQ
Cqz1zyeAGvOXKdfyKLYaafje8g4pM4ATTPfI6F7dfldkSTmQvRKEQqJwxu9R29Jt
8aB2GHXgZdJ3xaYZ52X9+LUfbqW8gZBbYKJPMVQOPUE9QAZ39uZlaa6NhziEQ8eH
GApEIh9ajbSG0gziQN0JPs21O9YB2kEF61iYkuHHd3tXdgRBjQ6sMGz+PRouPWFX
+hIyHpGaZbGCLMfMg5wAON3OHyhq559yzHj37JrAyBhIPc7yW+q8yMBK9FbR8YWV
n8gkoXZb3SfLdBe+OD9Op99k8ua+aFBGPLCrUVwo9B+kcYQ+2exz0HBT36Deg3Qj
YMvEg6PLbvq0r0pTH0G8qRxvk1qgpwdK3O7CZ0j534OuWrX4Rr0uqGllp496SkzX
v5EWI4GCu28aE6ogU2IGyFTWzQZf/TEtPrAEbLZMGTUy1lonW3ergUFp8/l8EtdM
qHkS6phs7E+2w+6TiMV37OM0Tl7hl7a6SrB1e5tBkVg0dKxiSqDs7k0Dcun4x0Sm
MTeek2Bb5l9hweurwqUVpxyHDxWHUHEo2aqdojkq79ed4RCE3P6UNkfvnBqLuKin
WTGgQ/Zn25Io/lTfoZNR4rSf4LYmEpoVxWi61v8fGB4J6GGCQFzSXSVsEpgK2ugt
n0NH1AlOiuMRCGI1pqwKLkEPUjT6+Kc6MbuGpjs1dNE+Uqcf9l5S6FNfGwu0AVr3
TVhkGDTy/UaCsv0Y7PWQJuBuIFqGQw8B8yW9wQoBhtPcnjGxfDRDS41+B48NCWmR
DmktMxsyW16FqODTN/ZUxCT9QvPRNdfMQbrO8pfGeC2SDxVR+0XhgxFuHtb4DPIZ
9Zuxgpt4JDxYuL3YJ6ogjrId6UAbHiyWVzrz0Q27XofBAxENWzoiDvQm1yl32m7N
uZ5lbClDs4kW7bhxDs+kShOnQZxrN/sqtjMchsq4nGXXtY5DnYw3kwzuA9O3ll4o
KuEOi+yWV0OHx+zOLk8dfM0Ole7jc5lSXNAVm/CeI3Sy9GaF8vdGX7Oa6DhXcrWd
VGTLIxQ5yGMqsJ7goHLcenOZXH/LiKz83w/Iz7hxvOfhLzU+M+FiH0cb8dCz7wMK
IyDwQ12WZXApqve4cijRXReUmLn/nrve18AT8lAnP4tvJUbjnMKLy4py0HDl6yUL
Zh56aLS61bSoxmDTwws8WhZUQZrXsrkWCF5XIR9XmNrkbC0Zj7/GYjICeBqSa6mi
UznACVpB4QvogyoAOsXjMSED6yXarvfJPGrlQ5vkE5zK+HggU3sdQCUKuPWpc69z
+gFXeG5yPbUTUzf+2sb/P6ieFkaD9IjdWs0CDyQ7XB1e9CHhKvrvM2YhRKzPmhpB
BUjF/zQ+QUAaYsn5ByT/+MXoWrLVmQQ+4VO26iwoSOLPojfBp9hOGB2gFoUJYPC3
0VuNzGbuPgzsKtdwVPymKtHOCkJDJTkwS7gT1680quRdtG9Gcz9/Q6fUs/9mHy95
bOVYkgkMIMJTi13DuedwzAr+S8Fm8o4VpC+bBz1GnEyIFgL/+G97X9LM0X1jz3h2
viUQ93l3X7Lq/V247hmeH/5W5M2HxXZsy4jnPDjezaeWJCO0ekTQd9l/baHe8Voo
wJ5JLshK1oJkddDYSpVQ1EnEYYe79FIRODmAfryUJy5/m8yjd5QCz5A0o9scSs5y
k9Pro+fap/9OnsWuql6e+SH14vUtrmgNoosyScL71ZuGQxvOQgJiPtroaVpjCIuP
1mEu5hlHQwY48b5KbGpZKe4DyHuSc4I5pdwpL1TeUQWvrVKYZXEmQkEY3a4609q5
SSKZKvHP4L8pdr/fGRup7QzvFmBXO7W5VQxBVc5fQSXh011EifI81YSflYi5q4O1
cH+PGSX/T57/m/EA9ECGJSuKICFgxGzfXNLJYcDYAPhiD1ut7O7u7irO2eu3s+5m
XoJig2n1DU+7FO0yGcQbotK5LQmE5vpppOyURzP/UnvdKnl6jx162L0X0r/y9t//
rN7nAZ99Z80DHiX/oL4qgRp7VCY7tK7TToJp1SO7hs9Aa7LEi5uLIENoiNG6BbME
k/EKv7eIgQgfrm16VVLgb+oR7ROA8N+yt0vG/g02gIDPi7ZLWk+I+1NQtvvZCNro
lfu1vTanUiLoehU1HYtK+7CESHgeMslj+GuwVU468mvXmQPe10Xd03QpkeVqYy5T
b+97lsqM+w+t7ksuu77mLVp/ZF9MGt7mupJVDnhIA8EPbRrYqeJV9zq/Dtk34SJ0
fgtR0Phsp2IxNAhRQuyYTu6mTjrGfzKVelzzefs86x/6+Y6mzpZHdH7YM3LiQJhO
G+AVDO8Yc+2K4CkZvSx9MxIZ4OTCHL8YqvGbRx+q8Ufc8E2Mp0CNWn6GZBPtBWqS
N5Zlgnmln3CsFZuT/SxToqOWa1ZLKrU6KCtvZOsA6zsi4IXbyz0XlSIiMWS5Vqh/
6mER5m7B4EgQTTq6SsDAaVZu7BnY+QSUTrHdtgJ5FTnXCqvK09CDvVYbxfKVtRYc
S+iYdG/LuYh7sHC0w74u+Pv1bx3aieuj554mF8fUQkTIKvSd2K0Idljx67SGV/Ti
8OcCBOXL5e85IWnXQlL7f1u9dP+Uh2UvfhqU6USpfo6IjNRNflzKdfWQzdrZwASf
whRLFw8eslzth8H8mgbWbN8cn+0S4g2hRWVIByKzA7QkfVuHcvZQCNhFusTFbbgi
SZqBzrEPQ9e6HdRdOBk4KMUKHoYcvYZ6iUzyWjJyiT3QKkXHaP8CVSfIlL/4NqQw
90Z7Hhz6/bxvy+w4SsNsgkeMfms04ZTCdfQcIOMsXjx74G7YZgZBQK7T6o5EdSHg
FWROcV+3+F3VFJ/gG2jbmKROQJdaWgYQZcI/8pPCK5pBki30FDxHYL5BHm0Utny7
TPbBQNXNNEoka3DyRtnaYknJs3hfbBjyNLvpMBTjZ1BXjwNr2NAPyC0s8glBu3nk
zY0dJfYWWDUOT9yZfkR24jcjU7hl6TXvpmwQeZoOSICc2Ybz1P+8M0dIFUlFsfSY
jiK6bc02ApLz+p/JwTIok6ykngG6Uj6CHeCOq4AxJdGTswe6KCtagxJKoKqhbYpf
pPChu/ww9/xKDaaStiRvR/faM/Tkop5T0NdBCU7dz1ahhlfvbxdv41pAu/yEWy4Y
6Vq8j7euCsLDfreAxqSO7TzH5qH+7clxJj32QUwujxtgeKhnC7AFzb6EPqMwncMY
nadG/mwYR+V9CjgWboYGIv4GYrLpMoWboqNxFTn8ED7VrnZnHux5+cPCZ0MRXjKH
HWw067sZqixIcw2VDLUtEGlCjs5D56raVRJsO1MNphMOEQXGQRUw7UGCCtceNs+q
HHezpml5Guhm+KhUmLvev3+EDXl0DZNHbo044RmdUU5DdcngOsQ6Lzc4PWIIjlpQ
zvhgThFzAdM6er2RZ561lxnxDchwV3cxuHqw56k0mZZHjeG4GmGs88TnQf9x3xrL
SEHZYtQ1LMiO2Xollx3xE3fscZ2CQS40Q7VN5YwTveQnpuE1QVXrSY8OmyulIOHr
4QlFc3KtEgCh2C7q4FEWP8hcD3HsdPkanXQPllSd5EtqO94fuqjkbxJT0Kb8Ioi4
PhLjeGugyJ7wq9+n6QJ+/0edgIa1JO79kFCaYOQdMtUqHZ/Z2l6/AN43rSC05OA2
DJkBko2YMNF9FZo2XzFqkXxVZoLi7tT9o5szb1vETKk4b5crFnit6ZOOk2Zm+M04
SmwfOjVkykXHYeX7RbPkHd0C+/T1MiqSKCUF8iYUvbz4tfo3aRy+DfOJmf8p9D18
prqpMuPLObq9M8UMo/J1wRs9ygEbdkPGAvo+IAcULIdZfh15XiF053FKNFsOxDso
qRSvg/wkaGVg2X9Q/61dbxOF/y+C2lgZRasNEOJiShBsL00amuugeyNc4bcNZcon
seLawVuQN5ohnZ5QwePB7vS8CdBescbgixf/AWL5JYJTRkaoLiRWZ9wNPocUptS+
7tctULxE8JLJzlA2AMHqejD92JiHDTrRknqIxQiIQA1cK4/zaqxAs0JOJ4VdQcot
Fqm/CkUt8JSUWbt1CslMdy6aRMJYhDpPAA11wdAQWt6HRPakwCw4eDK5AzITHP6L
2YmhMv36WJMCxJA+euFEpjP/4D3NwTmkCT3ROkx1hGKv0KurbLvjkQ+NY7upu4oN
4M6i+aETXByIvZFS0EKrY0+EnzqRYe0VPM6RFJ0Ux1YOj9052xasxwcBHfAYvhif
mLSW+KaLEu13tpwPQDAAkM58o3/0ofXEjOD+dH5nTI1k0xnNxKblA9cZU8eM50Dh
Y2+NJP4+JdY4LXwk1RzJ6nz+XhrBsc2CcztlAI8EVIAfui6NQVHFX2jFo7ELyNBJ
zM/5l+EFdPj9+iF93yerHDuB2e4ZhmgqFJHcJnccriloLKzf1jc20yW670OpDRk5
GYCYRQJsQdZR3WWxsPZEhUDt1CWVqzOwWwaS9MwI7h4Y9TyQCdicwYMSL7I4ShgU
frwm3mz/9B1OUWQas4mgrgGrTY9XnPIAwsCFUmidfuHPXgwoab6v1DQtEhnaH7x4
r/4OSaNiTU3mdUv2k0UxksGyYuS3ciJkYewuiitfgnbTjwkMpZH1ZHn8XgG9XzJx
LwEsUFyS3AZGAOeCMOHLEdTGm1VUzsKv135l+gZd5fk8tNTgi5IDnSHR2I3zqnK5
X4wE9vk0MVSzeiBALNEnPqKao3IGEa7RxwgApTGN7F7vtFk5/a0/4QtfnIn7+Jh/
7+j2Fe4ofD5o3AyOLrkZSXb1Bhm6f1Fh2LOIdOdkLrFhxTi8w2ZkL1DZAvu0t4Je
VqhTUM5dZpOcKxMtb7uaCKo5uKJLyzJ083ePZKT/XCdrmZbc2yhgZEgCSaahX+n2
FJmPHWXMFuqnVQ2+x8Q2ViNPA8PfIcw2PvFgQUo94AUhGPcsBMM4DzS/96yCDRFJ
beoaXnPNxCggjYnCg7pCmlSAjjYu/lP7cAH0r+QigOPdQADPRPqn8nfeeYHO5Qrp
47ruYOdXjhRnwc+REmMI7GORmOnlGSsyEarI/92ylE4UimCKWFe7JEWc4CH+t4Q0
9po3AC/AbOjJgKJbwe6ALQ6/NSSJS+ikTEyF5uj6STa2Zlh/7Cydm0/DDID8Xa2e
6tDPPjBudDSYlb2hyFO9JlTcVIxj89lAY627GnQcZcddukahAUnVNPaSym2lLmE+
NjBZ2SZEXvR3rCQIYqRyMtOaBlFKV/kC8p7sHDQoTd5UoGq1v7qpkg7Gab6Gz+KY
CdS3CbPVMO4yUcdbkvMYdHHR9OznJSFMXEJnBRErRtWX+xHMi84pQUfO0Ny3LzFZ
1rDvag8OZRBpo20T7/bli7lxkKBNf5xs8n7LIe5e/aHEQrItUtt+M5i/rDqn0kG6
f0qnOCH6Egn7smH26TthFoDYB46rLtp3LXCqYcsUNlXGt1tt3EFwbMgg8mTuHZpB
ThFUy5VzdZ0n1F2Mfeo8JJJP1UXGogU2BsFTMbnAvuL/JOWdUq3RXFTSOSRSgZAW
lAeXG0KOFsNetko10dCttwurtpXbLBZviHdYo6APduQNLvdnvphgkiO6LO5rRZBF
n4eQzHuYPftRVQ/4JnnP8W2KyE/9g7liclHbEt94TCOnYz6IJfd/SbLtGIb7Ci2o
eGYM3DzFiXpIeWS93ctrkXlt2ZlcjX24MC1D+EW9u6PZ531kI+kIKic3NB6YfjFC
hf4xHhKXGSTyA/0chzW/jMWtmfkgMHoIobIvDsmaMlx2S9XM9ejHdraEW8tQlA0V
PVtjhMOovfZM2PErLuXEUnGi8ekmywHwfdTDWHVUTD2PvaylahOoI1QCH71NaR45
mUsTWQVcXX2wczuJK+vG1fOyY8MTUuSFC7mxxrDVZb6ubzaza4iB5eH+2GzWu62d
KSz2C7kKuqLqtQtU8Cmn13Qqli57+wcZXvxOTisQzZazOTSkNkmbJlzeouDqtDTc
Gf3AYpTMkzoxD6EruZaUlvR01NQWFUwjyG0o4H5t3+VeHo0ctOOwkGPhx2YgdS/8
FZlyGz37c/SVNELQxwyG2/S5JbCF7pKPb51gBVq7ELark+nThvWzJ/7ydP9GsGQZ
no5VKorvUwE1QJEky2BlS71McTbt1NseTZGWkO8AffkcNGOgaHGMTlIlWt+8T3VI
r1YRvK95xvdqSLo1jIlO/tMDBLGVuA1zy71rS4PXNofBihchR5ID/pJBVFJknanJ
+86cxxg1fURCi+tckQlP2uC7exmpjfpIURnhUohsdHbWOC+MBlnvFol3h3T7Ealj
oi6T4u/8/tkKYGD5lYBY3mERcP2cvqWLU8G2zH7MMhJeWyMk6qb+vxt9wA2mj+bb
ktk/I9cMXCWHiYM2hX7DkuwdTHYd8a+zB7yFcerOXs4DfXI4SOupeuXKpHQzl3fF
2xfMb0o5fyWfQHvh1o+sZzIc2PEZsdlouTbsO5uwqslzcU2fMthGv3ONOkz8hS5+
bChU3iOOdXPnB/lyzaqg+g+j5TmcAp8KV7WpkW4YqXqxg+ez3VbznyiUJRzmAh1+
ZevGGOfyFV6dCp2EA2nHSx05dRWkRF7TDjG1qjgE8ognUUFZ8WZ8UjIQfrabazOV
luoL3/45/MOW1AeDq6/00Jfw7Nv62XWupIK5JJb/bPHs2fNMQSkF2uwu7fuBYKtV
lRApnskhIYZaUnCeGZbh8Wlfd3NmlwXVlrp8hQRqcMyWmFua8fzf1xranBzRkYWO
K2e4tzpdrdCb1eQE7w40UcLOvTfWkYwsg7nryS67Da77L1xycKP0PeZdGL3nQtBa
X8+A3GorfGdDYi6RycwT50xWnsOH6QTvSVFfe21U2LcvoVREioZQFXzo2HIrcTyL
dtKHrLN9IdJENO8zxfCv5q/4G9A9B3HAVbCeln4vtelLyam5/wrHG22HmK16Piz1
IsyMbmm551jplmK28W7GEi+DBf1XXLZiAtqSX1sZ5m2QpXHQPhK9eZIhLW0N25Ux
6aHEFGZ6Ujvgr7Hzt3NJrGm23UzesjpO/HSShDOZxzL+ecq6LKOKD4FdsevsZubp
bPB/jn8FtLp1lSiZ7nktEio935PK1GfHmU/m4mSBBaqkg1omU1liXeMhNS9Q4ghT
xrzY5KgjkkfGXv1aPl4m0CATigkiUvLHNnWl8fOOXPK2oEoGJyJEtQ38HBfI2BEa
rev0vtcwL0APoeovBJ6QclWiWCEIrQ1aWHq+MyWtf7rUqIYRvQPnhPyclUS3/tnI
/ZXs1BqiSlgrBI7L7wCFkQNh9pyZMuaUZnM5agL5Br47rJfaxQjpmFofybsvmc1J
CMqtUKCjDbWtzSqBzTAbeWLzgH89YFQwxRUGqQN261G9KOHiH+N4TeEBdC+RxJgM
h49SsEiayRTnZ3BHr3Bn+w2vZL1GqMfsNc2FqyJGkmdRb4UgaF6zMRH1mk1J5gDx
rqVLMA45rc3TcMYgZxwWibhsb4eyJl8gbamafBAiWHxDl5wExmrfQerYjdhYGsUL
wYLcsIbwyPduTnmM/3bSA15AoiIdBIEEITbwjP07biHeuV0F9vvI27tO3WYJbFsi
xqQDR89ZjitLNWNnFn5EwKxxOnkdaqUdeZtxv4TGvJqgDklUWkzRCeVithvf7gG+
gw46Un8iddtJntqOVWk3xbcRtsI9bLtX1+YPb4Y2GwalqQjz40zM5MU7/7i0TZTi
n6Zn03y1cyy0jpAt1riZU/z7yRUIyB4+ADbk1qgogaHyadFxgazqPkz2x4DgpMCY
v+FUnxf5LUmhjpZkh5e/ikv9YBzeVZtyCSvAW7kdkDkf45re5ibmBSVlo3brjSeM
4riwLx3ci5YvJixDymkgNUka48CapswVhx/pUbPI8j0wqL6LSc7E2rEisSGF8bod
9OSfTqRSvIvEq4dnW7l9m1murpZP9jmrg+j/ei2BjoQlqTfC0kPPs5cxO9FVeU7G
5zG3sriUfHnvjEDL2IoMXwdNs++zf/Aqbh0UDVYUj1HE0FKSpP5f+tc7kQYn0xim
Srcwx+mtdoJp1FRGLeoqz9h1pmbYZrZsms0qyt1fNCA/pFRFKY75vOzW/CR8RqvZ
Zy9gt+7U4mj5veg25yXWQNQ3Bm0U0nJ4M/oSETgo9+cmpoZxizsG7ZuLFt0tTtTV
LQwX7HCJSyc5WX9RMrFarCkK9Du3miyNqDKW0gCbLBk8lYqLxCUPRBsG3DhRXS9V
npNAtpu9BMsthXXHqG78p12bzN4qjIjG8xu0VYVYp0+HOEwEtLHsxvol+YtnALqD
v8E8hPt7mKpL7x8FThpOvOgvYizvZar7IbhdOVmwZLl7lYoSCsXgp2/S61wZhKzl
KjjtoVJJZouIQEkJIGbAabyHELpChzxtm7TjDqdwc1b7IbhHSDykZWOh1q6HHN7N
4p3l2igVkPYVGQ4CKNAsw38pgU79LTFR2fGPFKEHSH2srlDcVBEntTZ2+dHkzMOu
hEL+fs0QzbsFPzzAWJ4htFnQBh6PN3ICTpszdxxIcsOzs8/kTa/vXe8Uqlob/SfC
k/oK6Gt1sIYLUs10KSPGPGJTn0KdglU8R9Byrse79Tpj2Rw90HQ4KUb4SwxtRZ3c
48nL18gx7Ypqlb6N2CIEXAYbO5ybN+gfFunXpJqOAnKt+nCSUe65SE3InR12g3j9
ssVoabMq/IVUIqgB20HXj84nKEQ9ssG6ZN8QCjQ0lht/lrxnowpLN8ZiXiEtHrJa
7N8xdxIfbsp+cXYEbDJxS0XJK1LM3IhOf/hz/UvB8/xIRJzfRbSqOeqTRojIE4Fz
HCCfwnqfYhsgsx0H1Om3KiHTHBOLJv+xnsOxLoerKlx3xkZFd/2H+8CYojEEJl99
gfD4cZxsUsVbGDFTMxFsgeiXAWMmmebRPjAg987RMiO8kEc7FYecH5is4+3kmi2B
IuhGvbChCWt/Eq1vJPozJQq2pDXClValBDyFFe3YvQ6d0r9dyI1RlbDSp10QxlBG
+JIjAg1hmyqQHDMdUkaQMnm671Fb4DR/4HqxD+K6iBDu/S9+aYJyEnWd5tfsuhqU
CRx1xXdTlrrLvHbQwMxJ9FGR4fqkHT6vK6PYuVhANbAP8p+LEiM1Uc9x/HziVq/7
FxuowRw9GUvm0pMdtw4+/3XgsDnrTEo8fUObm3uo17u5HVK1ghwoBS4ueJWIQXlC
7f+fLFIA4C/hT5ndfvWOWR4aRtxlGic1Ww6rpavxibxu0CKfieYNY2GLhQkZVjA8
CJZdBn3TnhY6KNbGIcDESlMDOBrhsdCwib5Teu19in91wxvZRH5HPDz74+wUpp6c
7RGW+CgEGwP1yx1BzPjNzrSEuRh3x1HbOuvzMBmy+PZj0WozWgk6ZyhPrGAyZjPu
IwHsJ6WV5zoXzwZd4lzkqV0vFtOu50pLpcxRKz+ryCUMQcMwic5Cv3gtiUDFaRcN
MjwGfZy8JU+EOrnrkbCUxqxpcqqdSrVRCXRKBtTv53rApJarDMzZFim++99+XnP1
kHcl/GPmgho/9WtneLbqaoAEjZzzHLvimVsIBHnzDgbN5VIgAeR/W1Hz7lMhvnK7
VFJ+QQPV1pc4J9I3psRSty6IS6q6LBtoa6Ud3eU+QBqxL3CtwaVONJ/dJw5c1kpX
RzRzL1BgX3bqdqdDnHQfCF0S9TGsP/1u82oCI8//4qU+fI0ueQUEYBA/fQUeoqHT
MgaLg/hFCtf/gUIcxJ2EQNESmM3zWpYFKCn0/N0x9ukfIkxPS0bBEfwpsnFWXoc+
bkAnc7FUE6oBroFSoFFM7OaUa+UW1+PmkpEitw0iJKGIAVSTA8wqPFLHuAaA3Lec
6gltx9ioE+ojhBjkMKTK8mP8meaQFqAAA8basCmzWCcGMYCRJFiVt/Bkppj+SEoH
LA/CRdSrUGjs3kkN8KcUYNnkpNt3P/H5+dz/6vlbQ0lsvf77DvtAeqV5mhb+da1P
CAEeaNFfd4a3YgTh0wRtI9VnK3uNFSn9bLz6nH3y6IEaBQ28cVPh4aV3PTPJME6P
tNEXYQDPOaOLsxXbHJPH5KvX9L5fZAemjXDng786gDwlAO7fQY5/kh0E/U6KC/nK
N2OLeUyB7s8BOjHUi4fO+vBlvXoyjMfRcp1sdmHidtFm4hZThIJbqGcsxbEZn1hE
qjXuHP4rhhlKnNYmevTOw1Xl0JqSis363i7vb5YO/MLysIRDoUUiS0OS0F92GMwS
g8YVEQJJxhZM9zLvpUKM6cED8aCnLu4tEBnFecQ7G4dsDqCpbLYT95DY2d5oxLBU
+F4BBZkCbFVY8SCgV1To++SgaMQ9vvjppX0Z2ErHXiBXko0IOPApLr9M/LvBam+4
+6BZivd+DrWs5T/2QK/mhfNZI9CrPCbsfsTMV2fMgrsOyrySj2ZzrKr8tMz+JVBL
pQ+prlVjiIPYpABIkCknbQL2ZfhQ+g8SQRLDxF6otYNPLpQ8JpNvtc5ie/rJhB4E
sH/IYYE4dVAs/kx5wnyWevPJTNL1MOD7tbOEzW41kRwnhYE0vWIE9fHTWxEUBWKl
O/r3lD+BfWEps4V6GRiyFyvFZai8Lc9TPscyUYy7EFy5MzA1mqD3cszqV8IUuY3V
Aa8fHldguU/mAhryE8DBqsZimA/V+2b00ux75pgx4kMq9LQFHypuU8jGqCB2QkXT
8M5492PJoAQfgD/kYE6c58VbqKkWcd8RShO1+JUkiydtqgM1/28WxZf+K2c/pNyZ
QTKvVGfhNh6/ERGdaLQphcO3ws7aJygLT3zoBnMRE7Az40xoXzW95kykEq1wPCkt
yfRPS/G2BHOfil5cNkQj0NnrByau16OMhXFu2yWLgTchlDs9RVkGxyByzZVskKCP
UaG9dOsX1NOmaUgEM1EVljvw78MF9xlF8z5QrakzC2uj9I31fh9stdXydJyqO0l4
u5NggEsd4reXHSJ79nrgPGIaZmGkgu6aC6KzMjKuLvbbM9N7iqQISRnRap4uJe3V
euog3xtn7Vt3DAtv5OXGG9WfnWqFUv0N2tnc5fLGsm8bW8FtZKBF19zwjn1Z0ROj
jiZhIQFJwA1K9RYwtqsiHoWKKRzoY85ejgrE3q8a2kcsHjJ0Q+1yzf3HTdIukaqH
LTakG234UDwD4eSXAEaK7K5L30XQgj+jrJ3GDc3Hm/HuqlOd+2T5Mjpzsmtt21l1
ffO2+VwJD+6CFmGHGmaLVAOJBGqdp61+iWvkw24Kiz7jDQOEFp4M+Tqiq81Eu+ys
Jt8MWYNUfHY4oewdbnJ2i3TxZ/IJ8yar5qQEN5/oVoxh32CjPlzwtiXg1M87B1Zs
Vna+1sFMsVwwwK/cbfrP9+EKN2juQM3fEYohVir/LU8VKIDRWywEA3ig2nm9MAqb
bIXMbhlMwNcG8L9WxiI/ZqjJOAPwzonCV8qc7Gve5JKRZg9ldlU5/Llrl+mTMj3m
kT+PIEbq6S05Npc50mX2LplnzccQsxteX6o7as1LawFUQUWqOhm/P59Ux202CcEM
z9365nphnyYASzjSa7A+KpXst01gqrw+VYSOIG5fbJyWYdYzHcS32d78gTFeLAbA
KBSemBs2UEa8Q425IH94kh0BeXds9IfD6gZbU9A86kfS10i6UzF48wVBeotXEvaC
QYfs+UVdgSNbFQB77Z++DiwpmfRwV2FlBwZJe1E/tASSPpSxzeQP2ObRGXMMBDKq
rGVVf+UhRJCOZgA2taHbftnSKahkTE6h6Ro3EV7jjNbarN5AVlBAEEb7tPQQNgYB
1ks3RrMeRsNVSCtU2uxS7shsJuXmAvj0wlN7GHl9952YM/Z4rtrUYysM6G5laIHZ
Rfn7/rfAHrtc0VyJY8xMLGWsdFcn64a+jdN8KLqlmw+5oZOow3AQeDvdWLU2FyPk
07Ox2pE5frfn5G7uUkzIaF6VIHUdnJ/KCTz0lizOrsFzmMA4oKPMyTfJ0NxFmJDD
K+NENdVON519Dms1fAFgFXI87qEoVU8kgqF/w81IpH4Dt0HOV5fYSHS7xgBpEOJM
kWSzmyofKGWiPC9FAFeIWaZZ/4v35SiN1hJDjbSmUQl7ghSK99eJaNdEox24gL0Y
rAkJDb5y+U0oWvL69ISYPuJUVpH/QYyy7F4As+WNiimK+uLL32N6LFEGt0U06WUt
sPHmSnv2HRTxXKh+0paJnAfnZnM7lzkH4ioKp8JYmTzmOtcNKyQrXpHQG9MdKlNV
Zw+FcNfNhp2Cl7E60Tg6R0h/bMYjxWjDbouKNSWTqdtnog9CiNJ1dy6hSBaTZ+dq
/XPGfbK6FOUP99Ptglcgn2R+0dEr2qFhJg+k9B2SsZJLLTvhGIYPo4iAzwFlSMR2
nt1DHjDxk9cVzKtQioPldBO3Dls+aGFyXDLddDbHjabPW1pkyKMFTgZNFfiVzIj5
F7O99RFNHmRcegTL3XGg6LKSziXRID4BbERw0rDbClmxxs2Z2z983+vkehIOo34A
H1Fdg6a0ogOMnAyrAiSXIUzfhYk2CNCAu8VdPTheAUsi01p2LrB+vDpWvBot1J51
XhtyrP0AtyOOTyCilbSOmuJBRRhmwof40YgcI/efg1WsAmCLoXbeN6fatG6mNRt7
KdzIFRcdPshAiOwFY0q2xLndC4QbVJl8ubmdw7I8emOfb22qeCiXQBX0oDuuXkId
fmNgPvakkYyd59jckrBEE4/vFUzqOkHzI2nkx9E/t69HkSOG89o/8rfk+U1l9HCf
UR0pk6+U24wWfCKRyyNBOI5OG5WkUy3pZSDC8Ef6GQdi/xRAG8NFxy2FByajyYfP
FWJw1VRP4FIp56HHUM2UpoPC7i9c9zLgTqv6/XkPM1PzxR9EU9RAc1iQFmVcbOxI
ztMvEUMVDkvb5G8uHerkYGQRSvR5sgnFsPGE2T1eKMGOxCmm2paUVdT5lKT61NC3
fJn7LCv82N8UurWasrl8T0+vstDMIshIodzhEPG2iX3l+PjNg8DURgZeUYvH40mi
udvjuT1uYkPOG86RwRgKMibwbCE7/Wm2b491Z1osPJlRT6ZawH4lAXeBApeuEnMO
+SHPRxMSfI4gEzkCWdGp9WOctcjiJCSt2uNuLq4W6MTkzXUJEx6+L1pNi4O/ZhDz
LjUzU+++ekRqJm+TIqCRdSIWtmpsGFUq9emhSMjhIQUgLKnaV5SyGOxPypaBhPlb
iP0SZlzs2W9XJ8Iycz+8JtKanTRM/z5dp86G56Jo2WBZfdf6Q1ePKEfyJc8P7G+O
3MGSpvdn0DyL4vA3sMLdDzLGpO1+51/fOcVH8NSpvO//phCZcwlKWgRL2pdjhwsK
RO0px5LIBI066jsYbM5lb/0BJ5Dk6wdLUO++L64R7LIlQtrmk0lzh1b8Fu2e7t/W
4c8HliBbvTxbl+SlIH+H3Z6uSZrIEkdBgCwqQ3u6o41+nRC27Y0e6iaSzoFqAijH
G3Kcc5WLJ3lhE5T0FTt/dQRBSh9+N28dYgJbcGd/1Kpct1WFII9PHVsnqHHjcgUa
mUUvSoTB3S43ceg8NbO9wSPZANVVrPEkfA/1Oj9S0wbpt+cx0j6b+a1DOiFHoeHg
xXiVOevggQ8i0L1twCDO4qpFAcpb4G3dPdCMmwAuhL4SsCPaovC23BG5cBRywX/B
Q3cOAnLtTY2EGmr3VomAp7Kl9hmep8Qi8UFMDRsIyZHpapKleNnTAecnMCtAx8JO
zcHZCaxatlUy9n/iJ2B5W6REX4R5+hAvlTaNv3GB7IhynZ7pXz8sb3ji8X6ZWssn
t6mAiPSDrPaiIu0EQaMSee9LdiZzYNR2KGysYVVj3NexvRm7VWReXkK1EFu5tIm+
QWJjHgcMoG/IwVPr5WIBR7hDdTZtTR/8L98YC0QR5EF4fui9I0V9/QTMVG3AhUfn
lKnBfjEC7U6GRH4D8Lt8azigsR3wJkZufPqrDXZNT4BFKIaDDbbDrZXEEkkByngn
D49oBhXZ13Yc1zYUwf0krUnkL8DgSjuiZUUMbOwdyYlbfZYIOhFV9XoTllH7zew9
tGNdFFB9Q6Us6KiKvarvCejtn8EHnltTOi+fTEomtB2jeGskS2RYcrQpLuIuwYOC
7pkIGHPi69d6XTUfSsbl49KUwaKC87HEP7r5+F/qbWtUu/Jee8988DtOQ9dAoCJw
IHZywFNgEJ2zx8XB9eiHStbkw9wJ9FpX/m5cUMkVZisGp/ljdTMXX70Xfo21wc7L
CVy9gpf6NynGHSlIkriY1GxRDFSaq19CJjdpmXE9qzA9WDfz71QohzypcixTpU9s
WS+BkrGzC7go5qP8zL7/A2vIMqfB7vNUX2FH5GRm9ZgcBV29YA4WCBZYu8dfZTAh
IQYTmQQnmwl77PYJ7wkwdIqluJRJ+8Whu3O4mknDjsensh0nSDE3UXZ3QKWZDhRA
tLPAtLERTU4/r+p97IrF/CA4MjhfpG+qD7igaSQQahsdUzPOnHqk0LKJ9kZB1kcR
ee2HE90gHLzHbc2ZI766mDQggMLJlSXJJ3BDE7jVye4Fwlfg1VPvuJoffX1k3Fjo
hXFMy0QGG0hJYfJz+0XEw7tgCnIqGxYCJGVXUtbTXeq+E7TK/Oi1g+D8gy3KVz6J
lX3NNBLfGwTZjW6/fEku8lq+XKeDNb0IRXcu/GhvKvrDegFMAGyvfotlVKsgqdU5
ebb4mEu7G5+c9F7U22ljc0+AEiyKQX3g5PJHHvhRS+3xyhekKFRrq+rMul3VfW/G
O0hh9uHATrz/uMF4UQryP/uU3cgLUz24uQxSBfEgyrJrA1jLU8MQ8BvPZXX8Yf42
wQja9hXxW00GIs2XjsVpUNQfrLdMTiuo34mhREEzIwPTDU2Axw50KQkWajaJ58z2
47/x0O/1LT+o1SHsID5vNscFAnvcp3W2idAcRpw7ve95SuHUUFhjBRhfGM5r8ezX
C0r2WcI2RVyb6hqM4InlI8qfR26nhiJOX3QenAGzhiAnsBhGmQRcbfGZwxK7hIu/
YO5KQVQH8e+cNTJQHf0CwlzWnvNx0J795WTuUO35JVCk/nPikRv5VbsRQmk6fqvR
P5mOMNU38fWatpJYEHiLGKyjMIr1t9jp8iEh+WCC2iytp+gyarTvJCD3IXDKLjxm
6wUbQLH06WAUCoqtM5OsDj+2DdWX2OiAeKSr4k5xWVZdcbPPpQud89E1wXwniXVT
sfFNuC0OD0BmetOyHvK6lR+nlYN2avU7w2Huqz9bLD9FE4Ld6J5ZHDXz9wpquZ4t
kdt+CY8A+EzYMhGkrD+Ima8z14mWdd+moiNxXf2xRArA8HVoAnK+OCtMLf18oS0N
TiQFNEAn+cpyC2uDePXWnHIJzOC4Yko3vN4XdJ1L6wMae9S3IgTJWTtfLO76T1lj
7TzOt7j9p41c8y+ReIKoG8P3T4n204XcuX0/uObSKerB70A1DwSbloJXaqfBY6gE
U+5VYDbiNrL5VygwUjrFUgkO8Nv5GWj9Nf99i7SDjJopTeec1XdGq9zBUYiBougL
9onKxsS86ZnAnGWs8D7ONBz6r3ucz7Nf0QfIU0JgNuZtqU6XAAGtxG0RsKTzmORz
Uf25MloBTFNQVyp9ka+3q9E07Fc7C5evUJiWpRI2SgmNmHFIUZwVbqZnKhbp7fBe
ra6fbWd//SlL1CRI3CUyMc5ip9NzpSnX9aDGwX4L7NBkyopCJVzdvzX2aUqw0dDE
cUR+QXRdgAAahMS1TcTUgkRXZbuReO+InOz4qgiWG6mI9JmQJTIkF1WSVCYStjyI
tV/PZWqVJGdXrSiVXmAnD9Fh3Z4X+M5X94s4S7aYtUMBSGAV5NYpxBGewCvDI6OB
B+rkm5aXcoL61HLed5gVCDcs/MRt/0tZVtSt+Hu0pnwybntwv3h1XY8y/2GNWh9j
bjP43s19oOJ4cu858aSiHXwjKY7NbrcpkKmnnylW0l2hwBuTTJUCvlCYPbIk98dJ
o/0clnZqBV64FNzdSji+JGiiSeXGrNYDKeg0P2JrTaFFjRa7ZxdRo6VupslqEb3b
jVjbdiWrE9IptPPwVHBNfhB+VhUS32ZbCp5qaDYn9eMs3py98N06um0I8ghNv9KN
uRkRhcpZYRzLEsZoObU5ndFSJp6eTRDZ2w0qXBXJeBtzsq/DbkbGcgfsLeizFF8z
hfo4FNb6uyidqvYo+JE9A/JSRu4hbKeeM5BKUTNrfDniQbVY8aXV2eSCY5IJ1QyU
JXLYRTjJF6KDP2rwf1KmvHbsRFWHMzy4djozcSsSzVDEFMwMdea97yt342VtB8vA
ydXvun9CmaZsNudHEbYQeZplMEK6N00oyvde1wkn7aeweWOYNpW96DQnes8YDMxk
l2AW71voZ5eYFA4Z8QXZRWjrRyllykxuIm4MNKru2oLT3LbnzqqJmzgptji1lcJW
TOMcdmzClgP6TUzKELrnTqA1LkZzJBgGBgLOj3RfsHYVJ+ZX1ARyvSPgj6ZF0R4B
jkA/00bXeLb/1AB5JSHFfFGvYfpvbSih9iJyDlI0zcWLBb8SvPnoyNQywrQDUftF
uSEpFRn+REzbfm9qJ0TcM8s0rb7XKzbvspg/l4lG3HqjTTX2ReEO2pYqsbtiglVZ
SrvWMwMXG5USo/+3OzmKCCYmgZMITIVuM6c2YcOoThcPzdMfJ6Bc1GhQ8aXu6h6f
pPFgMaWlnXEy8msBSeS9UKZYxaB0Tlhzky84tsGkhE6IZcFG0rdEuQ7Mi8E+CgJY
S9Sfaw8nSxphVgwjEGUlObSX+uIztsZpzaOgkiMCOF06KbDl37AXzMwflVmrj7NR
dARkJ062nWOgl4WUYldDdmdX2uE7+Br9/pcpXNnxMVoW7iomC9EbE1zPG3tvF/Rp
x3CJamj9RRjUxfVAkWgT6AjyDkbmm6mujhKjko18GWIFj+EJM5VupDmXo1lP8oqZ
DEwyMZkZbrLMGPujQ/lPaKlp9LACK64Nzm7ydv5isBiQ9zp3q/mc4ajAP76MpUox
FJ18cHGRpDPX2Fu53t5A2ohOWzHfpm4Nqio4qGlo37UXEZGIcYUXIjE0WX28jkaB
+jmDv6eKxKr2WLUCttyNEYzUyA5V7dyPxEwaz0JXRPakNI9IP6C+2mdmlxnulSdS
nRKrw2cCj1OrHHguDK55CjdGAIc4/Kt3pGGBGcQOWZJ/ZFCTwurD842VX/TPDFvf
Sbaq+2vsAVUQc6tXQTIwEvIDQCnTyA9/TE8SCWyW3rHj+SdoWYW20cLGhhXQ7eCY
YkZZ+2Il57KjMgPO2wtHHQIlrCuTAsvZyRJ/uld4hx46x5OeM/CfuBVXfmoD6/ky
6EfEazZlSx0KTn1+pbr+1jKkL7LTWO9YaUTPTGftVQVKkMhftj7P+YQXNaSxdbrq
RXHyy2qqetvYqwOse5z/404HCWs3dCY09oJ4Vb7VVhjz03/n6jWg1FUn3COjCcpn
Zxu17xHvSIuhzwShzUgc9kJOLR/SIMJUkUz3U1tHjhbut358vJ/Ao65HJ3DU+vTA
GE6MbMXRMy24aDZYcWRWyb6pHxSLyRDy6vgZtXs+je7k/KddKRh3DCCrKODkfCqk
PEipZbxhmR4di9qfj9vFJNd1PauwGh45uaVffUTnGZN/0H3NLrOE2+fUee6xxsWq
Zv2lLDlrVmagSHORyvuiQxcW/V10SJHNdJ36ut2e+i4MDapPOQTxWJTVKbnVajFJ
cAN2ixhPnvdI/x/BSp/R46q17/nYpa5zVdLQziID9wa8NgKBEjPYuuntC9EWgArp
KedKVrDM+I+Gbb8WXd4aS/A0tLzwNO0NavPacwNxoqkvjK4vzWiA+sszJ1w0ecOf
pZDG2ZpqDe6EKdQncmiGKIVKM66l9WjxCy+lo8VDJLJOItZMqTjHikDbhuyajvOf
osIsTMH7UWl7ThxokymGZ/Wl/amr6rCiShBHaHImf8TlYf9OC+a8I/9gwf0ETB+v
C2vKFx02o+HjqAwaGN3h3lqwjcUlqaiKemyczo/VzZegZ9PiAoxcTb5vjnDc43id
MShS5DcTsdbELetEFjXTq9b71eig9mvyhNCa0blkHfBFcbdaOZM6HY/MQZyhqz3A
967HcEI6qbyzuaifQPDqDCcVnzTqLFvpN+71hsN5n1mNW+VdKxiwMy5E55hTVuYJ
d2K6a21wXX27sZ/DNnpt6jReRGYE13qWsdsa20JPGco3Lx4xar1Dg3lj3PxNFhPC
g+YQvXv73Qo/dDPG0ZBzZToXzUKxoLqHCYd4swR4oO28gflAzGmcdwstC0YlwUDi
VBadf1I2oYeUxju/ugVx/oM6IOKp10h6i4kwbijwoW1VW32YQkxFa86mXxJu0F3y
Kkr0NKcdJ9V/IcxdmfLNCrH1eJMAe6tguKMSaUXAvOTbDH0GQ8qcihBTbXZVN/0p
b1jKks+Ii/hqzl8YGZNOjhaCRrTBBXT2g/Wy7VWBPJ2wpxC1xQ1wKXitxDtd/TAp
Cs8NJlPUhwQHNzB7mj/MKwemGHK5zca9eQVAgd3kCBs9ZA+RurbtAvbtJtqR3H4B
9Mo2KHEN0Z+Lm28vj1ecolWSriDHOs/Y/Ph6CJdxsx4gm/CvxkXGzbEwNQqHYqij
Yl8koBZQpO8JVUYkwuzC/aF7scJcVzgwYqIDuLV0TNFXIODVWigD0JTdFsUSJsOc
CEmQVm5WVy7VQHYqdKlhE0+MYzrkd42WfscVEYgljsoVqKOSxTWXM8PCr5VzrWYt
RYkwAKyqlgYWju4omnSWnFGZfhWbUiQEJXb6mS74qbj4axf/hdGY7XzJ74MxE8wB
l+TbGA5NZhjRwpSzpMAWr1U1709NInPPy9XPP1RTmmUlGVTOR/gXtmIo5JEQcv+F
ojY5WQkd7nKXGcc49L1h/kyO3C6rvohtbN35CRCXkmk0CrXMcGVGwwK7cJN9G99b
N+u7JEGtVHKxrjcTyZ+mQLuo3OaMZeU6Uz9ATJV8Ue6wUg9fSTh91xKEUsM9DogY
C4OLT3r5z+J6sX8BOAlKQihDI0KHY6/OBAnQi8LaD5ADUYR8CfHXPGe1Sal3rJ4o
a5e3Lnln4HGK8CVX0F4aB7vSnY2I6o/wsWs55EaBBrIOSpuBpZz/0pRTHGwWjBO0
a621VMbASk4ET4LpRoDRAqO+C2nkP9i3UWs7VlYNNXRHCCNMUCGCvBxX+wrz0YgU
wgavvoSWWu+a2ujP4XiHvSszHw6jpsDm7m3hwXCDxnRr8Eli8jML9TBpoUXvyYsq
J565BpudjuIHS5lmobPanqDh8G2QC6CKANWwFEUPRlAmHgTcrEYhMgE1xaIZXuLJ
REdAzvPQDvR2tmmZoSQWJREc3UXadbBs84LyrQYPYB4lntI0tVFh2laZecUt8U7q
iLWfWiut5M8ev+XbKmWAdQzuMvEDIoz3fWyNlU81jcaQPmyWBEGOe7wspcHNIHBJ
MSKYbTAIWRIt1sdgpbdlk8nsfAFS2jKHABTYOszl4GKJ9wdR7ZgEvSJuN8QcPumP
aCCTvjVj/CbTFA4QgEfMUPMgA7akeiA8Gy8fUVDXkl657k7Iwr4FyyJzag4//b7v
eWtsLOp/0G0TgaWsbz/ob0mWqMRHYTEOVtIKgJbBCkmUJFhyfw3z4+8rEIln3BJe
gf2B+flDfPynn+RQ8BtRsboI9pXR/04EKQEOTbaPGs4zCSivWMVQCA2vTEAZgY43
Wm8ns282gRBEXDkEZeN2ba7JfJ8VfR3AtaMyCWDYb3LBOr+1JG+2c7S1orQolzd2
5QJ2hZOihhsFOdDNMK77EV6o0gU52Zk6J64KBe1LswkCjV1shsQKGd+/qIgFhCpJ
R7YDMJ7HANkiLb1gw3SR/oDUqpvea1SbS2zYzozcas94ifyP5HG+mhGtWFCuqR2e
MWDgBpCIB2KEYvN7Fd2/Ypdzya+56cR5dsYPr8ypY9Ht3sHsyEGYVvC+NIx0+Rng
ivLrUJ0h1V/hyl522GfHAlTuq6JxHi8fUueWfkM38hIsaMy0p8LcLo67WFi0GI5M
MyvAm0poghAG1KSLYQ6oDiaeSSSTR6f+r90PiImOtPhjsdlOeQi5v66KPeQLJlg3
ZKlBBvFlUzMKeTzDmBT59KEi6tHBbPKINAQ2ESKuUIPCr7dQk8YCBe5IxuDwJeK9
Ry05hyDyQWtBalPbXHdM6HvFcYz4R9QnqfqmHe/ZvO3zc9Cz8YkYhQNKukP9LeJP
oiiqXjyyK1QI3dQImaVqgGCJDPlhr5P7jNco5Q4kOjICNbxkbC7+fRp1WdsCFFyW
ylawXyPQW3DY40zBNPlJbCnBpcFETmpWRnWwPQwabh3UnFRzkK8BuvK3MxhbaI60
P6jqWteQbwQwYRavVoo/wWsJtY1j+yMzYXfMEj4JlIw79iMeNg5GGuKwCZtU+LL1
GM1ZnZxry45Aa4eE4U2bs7ml+HdgnVsImt2XHkMnRAT1pU0hElYpzgYDkVBfvnLN
l8YrfLfJmPMHhlAYjadjnuCkC1EywsysX7vDjagqfEN3Q1OLQfv1UzqwhHWu8jfM
n39p9rtxyYLDWE7FhAMWUEquoeqInjKyP3vNNozhg+XEOU1rjYIKf4dyusLD4JHL
3VyoXQx1MaCGjUU0ADUM5V9hteggzT27usICphNFwoixs6cT075mHIyvidRRgVLg
551/2fuuiBWLJl/F6Z2ozgzWceFM/unH8mNvHT6Xjd0RWlNehHSzkSyl8ia0l6e5
RNx1hUmtzikNN5zowi3j0A==
//pragma protect end_data_block
//pragma protect digest_block
xtXaLL9+ujhqaYjycFNhkBqYMj0=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
v5wTCvz4FWYrBzAo0uEsiSrHr97nudLTfvZJN6cYybLjCqp16XCU++g/mtPi9rJF
Nu8FoiVhFLORqhoQQv3/cKoa/85wavTYSN5w0wofSz+qK8zzda6463mojRZl68Bw
Nv57h5MlWpnzUABC8H+LPT9HuvMpVsbEx4NpDN6IeZSPz0aOXmD7Bw==
//pragma protect end_key_block
//pragma protect digest_block
qgXyDxRuydUxAEehbXILz9CbcNI=
//pragma protect end_digest_block
//pragma protect data_block
xgETSaRuBQbrQD3t92X5dVhtNfMUroZ+8z2rBYoebXDft/7hs8PcttturMqwTFGu
CjuDFeuduFUOoFwQtllkNiigmLth8V8zeBT6PyOndanje8doeF6XLz6ftODuSdj/
iswIXPo9K66Wg9xACTn6SAX2RaTz+BYVELhzDZrZOkH/PYKwEMlwrQyVV6u4VvpJ
P5xned3oxT2OAQ9G7o3L7XW40q5JZ1lI/MSQhJptoPUx7cUA6BZlve7PihZ3FUnu
Y0rmZ+sM+if6p2Lgi2qJHmq6Xw1bKNnEr09ru6gxAzFkx/OlGHuLuNke1F9hRk62
+xOWdBTsLUBe6cDDOAihJb+Lf6yYbLIUTpzsOoXIi6X+vCk3qdvI18zR2G2sVJCg
1rJBziIizhNSBR574gV2iclPjA66f714ZpE7xek4BLh3kcFIcv7do6dGW9e5p7Ek
ms+XQGKbgjmC3j4d3LXBv4NmebYI9wxehJOrnHWnzwM=
//pragma protect end_data_block
//pragma protect digest_block
WFrgrgOxScNQwNdLTEzwnM4uEH0=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
GROCvo/i0AM5cSyuZvmyOzqe7y3mQjXMqbCkA4iWftSSwykysyAX0f+oNSGij0QC
VBHhL6nVnJ5zsUrhgzBA+rqyRtFx0tYF3oTQ42R65TaK1yiphyp/yA4aBJoufxOI
a6OA0XtfwX2I3kpW/IEY6j5QzA2+Po07jJdYkSVoNPFm1psS8F2cfg==
//pragma protect end_key_block
//pragma protect digest_block
xd2kZc7JWNxMfHUbzw7szUtQes0=
//pragma protect end_digest_block
//pragma protect data_block
N1YNYISf7rsqRfpcvxokqAmi5h/ja51O6tncfLdjijHKfaD2NnSnS6zehnxXXDCJ
2ufGzrf8mX9U8rsw2Np6lmNfYoVOBMF62Y4+/qn1cc8dN3ifJb9A2Y8ediXFC3re
mkvhzz0RpGaT8xHKqfzTcgiRUBTCW+63hrAMQEfEhRXKf0g+1/Oo1cB6VEANkSAG
303gZ0j6c9PGfM9G+YQwcY+kYh0Ll1PHI4uLYuZ45HSEuEz6uz2v9CFNo0AEv+DP
ASUc8KbtVEIdpip4ZXbIVwthmia+osCj4bISjpQoO09EV/cviDFclucRhq/SrXEL
3HJyi9rMe8zvOnIBqrZguf2OVGEK6TeU42oEMv+8GjJ3Czkst0AZT6kT5B7HW6Yq
A8RjG/s1AykVcti7WjF6x8OKxTwXpgeyND+3HCU4YTtfRAx8pZsGa4s2nRMLejeK
vLVwITENKGTzKbQdxsmNAcVN7vUWXf3VwoGLHjJRlU8cOVujPDRCMRqWdxeg7DBU
21GxvHG0DzJBe8TcNvhL6Tt3wDlCiipDW0oybiLb/Vkb2A6tBvMsv9pXDRELjhA0
cMrn4nMKuYpXtyl1O3TYx+m5MRLzJp+C5uS0REqzCuobDRyKaXH2G1HFOKSkAtQ/
8Z3pjGY3CeVyP7aTWNcgdPIgy31QoGARjQ+bzB5pqY782TIiUTlhJ97xR1Ulg4bA
pli2Mg6SSzntXB/KH03DQ+t5SR+5GVfuR76Jeb0h60bHQhrV7qgjALw8YRJdn3UT
lEC2Ypr/Sh9YjXDtRFYb/wmfzVrCRe5EZXw5fBwQuHwtf8EYMkCR7aPXvQd455Or
exYpmQ8WwmEPEAzCjS0wATuqIQiow/5KHXUtlUjc6RZrOn47nMXTxZoVUrFaZgez
kthipnZ2gkVXSEl68vXY3D23vYldfKMFdd1ASs2Oq+aNwrottqZlC+UafKxTuuHN
UlodYs55sI2OvLc4MO0L6NVr3ar6vBG2r+BdYcBkEXNegP3ZFSIC9wQUCFRYHlmb
jYcG7GE4FrTlo+CvGHJmy+yJTff9pwsCKvkiI1KNnb7xv4JEef3nv2OcCZ/HoaHq
SkeJ9RworM1k73Zij4ulO8pvVg4h2qF1k5gkJJ083UQh0k4nW+qKJaHWGMqKxjBF
NEGTadM/T1p8betP7cMKG993xoCGrB/vPOZmjincyWOnKlceNJH2ffZWMp1MCGqK
wWHyhs8rYGuQVEeou1Vx9sIQCNMXS1Pcv+03d6GlWkii1R3wHBawY2r9EOm9emLw
2EcIDNmNuaO59B9nggn7BOwUo5OITagExRUUjrq25hdJSRg+yqnzCA7CZk4OSsJc
9KUeJeA5TelGWlyxQ4omtobSnfJOqCWVf4Z1YIZRJTRRcQHKtFHRMW28WIT2M74H
Bui0tf3EyT51MCfb2nCCEy1pgiuO3s7HjlNyaq+FyqkSpFcGpPgeRPMZBtbR1Ftx
IlximSrAFRyoeQaqayGUWc35cI2+1Vf7pPKx158nBzcP/hPoBpTPgCKot5wyo3YG
FQ1BnjODzARYsRAfuUeycukQuwOxTKN2DA0Sgb0rCj6L1jzb75G3FuXFp3w/JS8P
uOH7348R0qIKvxF45S4Op8Wc4rWYsddu8I6pwYnkLWfceMbmpBM4IzvXOPrdzxo+
u1ZQLdkOlc7jLPDYsgC+k9x/dlQDEL8LokD4x5bHVuE+OGkHmhO1BOZXWyjNrWml
0Uh/Gb+2+YKsnmfyPqTZCyRzEDwVXQBhWkq91ql+CE7SGDlwFQ1i6rEXuPKSG+5r
5ITplj0lfrny1+lCNcNz7sSryT0v5iQb0ebhCsKZKK2im3BHooUf2FF23wHgvsb0
s3ci3UBT59pW3+SqlR4TO3Ur5NZefqMu1r1Oof9IMy/HmkA2RYiGycWx5nqHIFBa
V+pFY/0gxPkAGHu7oINuHXnjhVre6JPccoC8fIHoxpjeEZkm04MmVH+cKJiAvH6b
I3sCro5ipJ5z6tnPldZDPgRqh+jOJUlVWA3GvhlJj+ZPG8i28bgqpbFqrXBrgr81
6CeCC3Adn5AfyaMTQ7Xk6DRKC7rwNY5zuv3XPLaHl/ztnHr8kgQbxlHV8e+Rv07h
GwjX7zhM/Up7ecBZe2/4dg/nbn7eJAm/K3JIk4dOmlWQx6I167lrsStxuVemMZBA
LIp7PdsVbBISJqZvSRxz1nDMtuTD+9udfQEDN2S5qBWj2EvXFJvtBSmWw70ureUF
2GSH95UX81ngBjjctFmzNOUNR5xz41uVGmvrLiYBqEdxGzvYWjVkV/JRNH4rvoJw
pufG2vlSo3X3hbDagXkyayyQc26bPchM6u1/kB25Fmj1q1eYAgQGULIhSZNkPjQJ
s8pugCbKcoW7beClV39g4KKMrCH1DqzjBCs8/g+NzmsDgunFO9CoX5KmJGlazKyG
1PaZ2FgKMXrTVM7b12mkYA7DoWXHIRKUyLwEL5e+IWohWwFC3SQRKeFXtvdyyPId
THNiUhgseVldhrA0CB/QUJQx6hYqouAZj+6mQsGl6EQnSQrXS1R3KvdxvT7cb4Yx
a71EkuwIVbdL+5H1+4g6EEQPFlVq4YcVgV7h/gzp16CyaXH9am6NkO7sPW2bSELP
T3U2Fv4yfSpjlBZnanx0cg01DnK4Ct4JFFn7XrgJVakDJ6n3fI3i7PQwSmNqAeYb
Q/q4Fc0HkzcD+THJUnNajQ1QtgRkzqg77DD45JZMRKSQDsSKgLYgSMPA/qmQnhkE
+4PSxfax2Xu81oJcWnn2m8hQQB/2bcD9/b4TFR/IYwIy+T2byUqBf52u1Hix6z+8
dlDNUet3JCOAt8lOFo6EklvIi4GGIn9uXiV69O8XXNAYy8G0A/s2RdV/oXAwRjx6
kH0LKpuYIJyKrrmaP1JmJqEPHDW9z3y7FTlDgRv6x3YTQDSIOfNeXF1CQUQro9NJ
HiKulvoDkZ8RHF0EWdv7RHs9T+Ni4en9p9UwP9eANHE4OWhCbGTS4qaPTVwztwA3
O/WrbmmBgevWEaHMAY2V4USlA+IJ3hT8AsaJ1D365c50MSaK8vxQwX7ZvcGmxscz
Vp4pkQsUVhGuERfeeKwXCUkBBv2UPzs3Xwm4gqMEDrcqrDU/CYsnzGmTro0lVyYe
gAimAxN5EcWD+i+oG6602BxyiBBKQt8iMFBSKqIiUq20zEJo/YbQMli0bupr//QA
trz9YMWcbRbGL6eQzwYzK8gSbc/nQxoLPbxOnOzFAwVny0l4tEShse6sNxRdvn6B
2VlqExytEHDL+ufCvVp7HP3j3JQ41exe4/WhLE+WJCJ5CYiqUJaSe1j5nHOyCJDr
hvaReFsG4wJpczJ6U0kJ2563VfbP2aaCqXAiQmurlp4y/dljbhiIw6comI4CAPgQ
c9axRkiA4cDv61hxUmBWm58757x6OY7rxJmwo5CJjtoLPqq/6mUPdaaBGXSasmNb
qzfhemnylQGSEL91lwcRypzagzxeIBOsjN+61d/RO6TYVSPa02sPq5Nm95xrRvdb
SwIXZ9Cs/mFtDMcFWyRqSMD176XQKfKIzNd0qf/4n+JWdpR/ReJlCL3fGYtu7Qq1
9c2Zy2oayG1kKMhMUkZoebIoOBQa7qqr9Z1+x10NmoHpU7/CsofGF/LTA9n64wqL
Zl4nIoe+gMLfy4WGVuBY8RyUBbqx9XqYnJetFmFSNMpewlmH5SLlblzyv5XDtfQT
OpCETphuSBekTHBsEgccBkEXH5hyOWOq35goFDbVgxDUUvNlEpXWjzb+yCd9hj5n
TOfHoWMI8AdhaGmx3st3gU4NFVuJJFOZxTTrqi6/7jASyJ5JI/q4zv/jSAEXpYe0
8SD06kd7AfjiZ0uSw/HF3Z1a1Acy12qB+NFHP9uPh5Hkkv73v9KZTbjAUhcvm0FD
Ua7Yg+kqfDaHldyHLtlDu3713mGmGBHlQxy41JCZwMut9rcWqC5H/VdM2FhHf0O8
YSUvofDwOgU2bN3CuTDrVpGhEY3jtERs/RepBOdxEx8Clv87KhqroiQos0hKGxbh
Op/S1dEUOSJz1oAx+56y63G96mnRpKwJHv1fovZ6KsOr+Y/2TYZ4I0G3+OYq6+rF
51e0+C/9ZdaHEQFBCEgTOUpDaZHozgiI75il/yUKEepsLKdbiOm4yS5xpskoGdPJ
Tf3zp6Fa20bJntF5fovAZGXwIuENeaeUimUnlcEhH26MHGNQBUgy04nwRUE2ow31
yfiJF4U/5qpVmOVPm1DrTEoKICzxdV4Zjd69iSM8jIkFQc76h/iTSTwavzY20Ueb
RyJYwrJmbkkxUp2QDHK5RP8tS+i39NvUo4q6Wd451H4h49Rz9owRtzbEYp2Dkgnf
fUXwoQUbDH7yFQIWgj7Xe7kE1DlgrmZxnNul3fUs1bSaijVZfWw9zbPKlelLyUzu
J305HYQJZxMvqCjzQsDW1GcR65lyAR77uAR3FJqsgzLt4RrfRWwHjw2vMsh5FYe/
lG2h2kHqZPoVkIhkH2EuIGKKScg7yKi4u32O45BgNi3FWCH0d805NRZJ5BfLoHwt
U1BcsSjxFZhULXROlfIZx4iiKt41CX1Nw0J+c3J7RqO+9sNKaMzSbshBDWJiWN/8
Fc4r78k4XZzL8oPx26h+yg5Qkol3QdGfpX42lEX3+UQSrv18+ql7MEyu3j0vvFFT
BxkuFwNGSCWdchdI6PuJ1Bc8C+VPsWLb0rBY4KGr0rsbbqk3IjoUSsBmP8sqEILQ
HmPDRO1AEO+CLGEQGDok3F/6mlRHmczyJsHGFBrb8WdJtg1CN2+ez45NRwRdIhDj
NceyhrcFUz1tlPA/WTyWwPAcoZ691ZZw1W8wFRrIb4AmBLk1CKGfRVNIHTQCbc4Q
nLKArqVniDKd6XsrrTi0V7VqVezErb84IjDPxeTRbCkLpzmN9Aarr3FlnQMvxQ1m
2UYfBiv6iQbv2I7AuKIr44MeaObtuoghL1AiDMeJEKR7XqCTgNyC6uVSA9XPjkAg
vLdXfMdN4AdFq9BqYyWV4SK2FIqbweaw1fZaKsQBfUTw734g2vQSxC1azmmKrhAn
5iq3EnxzthQLraNj5Q18u2VSMb98Tb02TIl+7nA7VI0ftSQtas+dslw0fBPPt9uq
GhA0PjAZwlW6H6heHRwiu0SI/VM+U9YHs70jj8NoSsmLfwm2/3g5tsCgPvMcPV+N
l4/Z3SQQ6b6sEppzOBaZZLIC0O54gIU1agp8g8TsBz3ww/0w3aGulfoUjgh5OFG2
vHWT12pLtCWM2ZUARnVwQwTmf/NkNlj3205/7OQF2Je6ew+p37NMDgErNa+1CAKE
vNcu4B6d063AKija6oY5dsxF3kjhp0ztIXrkrQe+6kE3qGy0MK79mMhfV9KwHiGf
NPg0W+0STBOsY1kfWrKJFwQTfkYzT0mw/YLZh9O5gc86rA4o3S4OnAsYg/tao5hs
yUOHsmufwebmrT2UNx4lSxZtwyWNFk3MLhhQ5PjhixhOHJdCUqFnFZVsFOoz4EqH
AYW5lAW4LUrtgMr9DRG5stmHdx6k5ijgpYwMzpQsrBUs4nMjXWGkpmySMn2kbhZF
lA4Ba4gPwFQXkgQzIIai18LWG7CsdA6AnY7iOzLGgSyqtBNADYUVjev5Q9zAZ4RV
NIM3EA7DVI86FyfQOKU7geoL/J2ZkFwUxVXigHZaKnMbzL5qvI7SlC4xwIV8lWdk
bxTtMXH5jG98ZLQn3tGL4ni0PYS96xiKiMJaYbxubDbF3S8WFrcroAGHugH63mic
tUbxLk4hBrQpUu7+mEMPwigRczhZUvVGFQnZS63H4z5lIoz4fOa26iyMLyxB+cdt
frDF3dP3iBqM8Nn2zY4+KbPQ1uIlwZ9WS4cTIPaJ8psFlXJDP9oSdhXmHRUfzTjq
ghuLCFeDe0VZV2ax4ldjPld3xra1/18gq2T8tZ57kv8VwSjqXWdzFevrT8FIKSbN
R4Qh+8AFq1bR0wv2Z4wRhiRVpvVWCdjc2dfvfs7vGdpr5mUepY2ixC/aZ5HA7QxZ
cZqvI0qaYMprlgbtPFJHkeWbgkT09Tu1AXX0+h3A6SPln+FsS1RZ0dwW8lERGezB
AdirUQtfRe6upgKzcFPSJhvtqz0+osCxX0yPO/M0PRjCn/3ZHbozdh7KHGBoQWQs
8NtQ7smUF/NsC88ocTpl2FkA+E7KNuUUvE8wVXKKlE2yc0zdUQFHBBuhPUagj0VS
/tqBN7Y5dy83qQQmBTZSlxaM17nok7eZODWrzGCz1x13GmcevP32NbJnwFxL30lW
4HSeMDEiXtLussirVLRoWsY2TyrVL8d1YNmaUym6EZkknO/hw1tjQ99b/f/7wcsO
Qb3/sVwzQ25H9Lznoe7vA92BsNxF1AsOzqcIntHljgOUnwetZAFze5lWU03JSUrd
cwqJUoo4vGQv/WGSIZ4ez2nzSV0HdmeDEJA26v9Llz3myOa7lsmAgL+8CtHFQyZ4
xlhNutwmvx49v18Mr7ARmnsHOhX76OLE7kwo+7KVBtnb97Dw9zkIDrqDS8RyPIaJ
Hc9rkdWdjCbJ4JkTOiMncpMLrt+twk1Vdo2eFiU83H+rFw9yFbGah4nGnRzxmByJ
W+vmysm2yEBIZzjjgwEDSfCBHFuLJjM3xamJczW3r/ypCdDTPyPlnFhE3Mtsarlo
eLs5EQOw0faTetN85R7lulVVZiGdHLfB79jEI2/VaXe8nRGj/8oS4HWcE3ZbRzUw
e3OojlBTcXzJNuVyZ5YdL8EUwQuuq9IafEnkNaBCeiMuqmnMxVx7MjcjB8hl1hYL
ovmGh1bYqvLkDnlL7BFqtPHYHNuNXOURKjRQJTSleSTdCBliKkhI1Mr6ViIbPz4p
txhItwVslxl0S7lLyNGDumtECeq0MeyW98ei8dDJB1tyU0SSL9ujiDfPnmumhtp+
XrVdksKCmp6WMDMaN8XKXNODkkx6zn3etZmHGuBwj7+n7VVdtyEgxo2T+sXx5UuB
wlhzfYYo6LpeLZSN82N0SADEjsMWTCL+ORnmosVw8H5/2uCBC8q2ujrELNSngWE0
200hRm1AfU/ALN80xQ4FVhpzrqPQ8HZ+QGxtKbVFgr4yX3SI8XKzkvmyosm2yBNs
3bFz0osOAh2o/AyUrMO8R0BbXz0sWiNucpHY3Y5otCxMIEbgnpvurM2/gAGmvFtg
zmZxIMdfu8YfDV98wE0HdSM9Sl+uyE5lEZuy9DTPTJ00Iy2kPxj2r4GnmEMWWUzl
JyjVYdCPCVak8bmAsyrcsAitj1Rlg4EKc4elAavE0UfNbwa6zpBrgd3MFH9wzd+t
fzEhkqV+EhLiTbVnAR7BouwIjzewGWGbwXm0BRPuaDWuK2r5vspwnUhbuX/L8JID
QZClK7tRd88qNal0+8oVGSR/sKdKr8jjDNS24zrRQrmlSrMBpMdqE0ybnWpeI7Zl
olLNWvvy2q1dLAkQvtR5NP+Fznt9xPVL05kFvnjnw3IDRlkqclD+dqWAqSZg+z/k
a6+ouba1n/wwbcIkN29cfAJ/RC6S4/uu9ANnuCoKLQNnbsTDhVxiOswxMlH3DVCq
cljW9y8fp7VlPqkSEZNDwTcHTOb6jtTq8DZptX69/08O6DFzsmIslQ+h0qIqisdz
F6/aCaZOzrgqUXc67F5gLk4uPU30GfQp0FJHkxkFLzPAntf+Z/xy9PVNYeza0So/
s9o6YUGyRdm0oFLGQ9qFJAAHiXXPfI0Y6/KjZoCOsFSTqQIBgquuT0b6o1fpohlL
gONjwEXySBgf2eAyNG7EuS2EYP/XXN0zpUp/+hI6uNPJZvfdTxelZGBa82ciyhFf
NFzs1pr9UZINuvPMGKkaTDIvuen+45A11t3nvqYy/GTPfOMG9hZUn5p/jeEsiKPL
MYvmExTGvjuQL5eKtkjlYRDytA5vVuMi0C/Ncwm8uHpsTxMK95CKxpTk6et7QSZy
dTDie24rO72lRlDIou7UeRCEmKT8ZrGX27OCpJiHcG5rLN2WaIXgNvO9uNlS7F9s
pbrvkhaR9ah2RkruduluOGV+BnylmSAZoWijmi8D0qYxdysSAV2nLRsIl7mVZA7y
nZ1nCjRZaune+4IH/HvO8NUj7G3qfMXZRlHR4/XZ8diSbBpU+nPml1+3idAKugan
yQ5puVMmSzPxsal6X1ssniw84Wo+LnCDD5QP207FR2r8wtMIt8+itaCPTOpRgaAN
ErawkjC7yICVJfHGWf6Gjdcch9zXaeOboVIovc7orNjDy3dLfS27rUt3EZov7x28
VC56CV0Mqb3zmXfO01gtNyMT6wnXBgIFkBs2sIvmMQWBkPviXX9YWSiLgdzANAy4
4I+icw2JLDvB2NdsK/YDHdSd+PZjYFUA3j5z4l8BnmqRzfkqIF+L6AYCnGNIi4Yo
80cK/vJu3HlqLxIwJekikzM76lrHQp1OHTlNDcGmHg3YdkIrZR8xyXFTwZzfF40/
MQ4cBpjU7JPQZe0sbccDUSb53AUBJ9j6E9slHnMqRLTDzj/cTIAt/LHQ8StJkPbe
A2jetTowwYs/H52nWdGHbU5jaJeaK555Dot3ASXoEWYJPkhxen+QEoJEN2i14WwM
UOiLfyNNkBjTM895ZI6rm8Xg02JeTMat5sk+tv+I0he+HoD+QkJIY5IfxmzQPwqJ
inMLRLDL7jqoLOPSaNWrvPjXo1AfviZJJeBnuQEyQ8H4Kc1VCr4AgVH4GpFNSu1a
YxrQiS6M9xEHfAG2SQQQiQTcBkHU6Jd+5E7grJd/56um0NJqVfZbggJ6j8g1QC66
SRUUFwwxs94Snr7dmQ3rnj674LGDRYkSekpdF0BGqIZn+2orjHGfgucsVtvbTiMl
y9XN7MPwMbPDfmB1UndZ88I0u34PIjXO3kwa5nMLwXT7e5HwkOYPP5QE/78LXTmq
o1/VIO3hoNsZXMds0B45Kt7Sjh9Gj7h7fTZmsGnMWIyB9T97hkyvDnZ1s4XTb0iu
elMlzOfML/3uHef/CEF2x69y0mfGp7Mu48Zml5M1ma9oMOG24umjT8jwwG0wWyhI
OLH5bDhuw+UqVKsUq+Zdr1/Y/6FPPZQwXH88+5GG6NjJ+CLobHJfUw918s2tn1RL
WCUW9E8CAKHw3WW5RJdfbvpAnmCFOE6rmJQkccPFxO7QyK4sq11KR+Cy3jb6drXb
ZvOQ0IbZI4vXXfXXG6ahiqf0TttR/LtI7IYyO2JLZWTRT5IqCxyMemAsQfHaYctj
fl0Rjgw9KKOSoxNcRutDLWXGXZ2YIMO8JkQVbt3rwhzkioGNM4IAJ7JtE/GFG6ee
NT6QCjGXOSriAkC3VXW4TNuQa/RQqxaGcSSZ14MEmIilupKKs0JfMMDF5gFZiiGL
kwH93wruChK4cEGw85ucFfEOgOKdh80h3PLpoCZpI4FP+eXg8qKv8pSCmnIVccZo
w3GPx/8rmPIqj5TaeP6fUxhaKthiviFhBoq0YK8I6UUWhxJnsPajcVzXhBoozvJA
2UbsgmRLuAOIwqyxtYSfvPi0IfHv8XSWbwCUrxhIUX5H/4IL3owmDEwmkslSfEOg
7n0BuC4T6HUwuEIhqm6J/I/g3xesJc/GiXUb0TnDdALWOb/dHRy52WIVkx3VM6Ty
uEAbr/3nLI0kU0I9iYUy589fBB1uyW9Bt538LZBY9U0tyPoq54HeOQAZcvhzJmo9
boRG5LxAGIzTRnx97ir3ItaT9z4tlQZ6nNmq1NZ3Bewz9b5gsb2JQ1ulZ7x729L8
6YmK9zGXxhwmNyc2FGUPV+5k2JD0H2FqrwNX4o4o2ogtHfZDeeUstL2Y47+2MWTH
j4PEhQ1s6FP8wWWFIGIJYqphZOALAPfO6QnMtvv5EYCoTWrPmlizV9AkJn582/m5
yf2EgxbySv0SHw5zzn/q6+7eqQnHDp3piM0ProOaCyzdtjknp6eOwNSaQCbr3W6R
VfwhEKMV94vmJWCLzdpqgQmrZ+wWXQfrauevoK2n+kiAXpf+wWyV8y8zwFyS9KDz
+WxMr9vRCZ+76kDbVmtVI1isCgi8Vj7cITSN0ILbjIuY0zKy4K0g5zJrl5lyCpJR
Hk+QCXf/pXu8qD6EjauQNWk1cO70IIucSClRfD9CWLd+To1n7u3q3tN0tvEQlnkL
fYf2coHsDcTlNIIFvSgfqBeQT/+p021pSUHS8QLLXzzk+5sPybHk9QGVmg8F2khB
6w/5xxX+uipPBOyF/OWe8i+CIfH03Kn7WZO2UBN7IY0DhHRyRnc8/rF+pjxuu78v
oPahLGCBU5V69WPL0iWo59jFFNMJQoHP9d7zNmNaFZGLREuqKTKWB63o8UQpK/az
Xf4jTgReHo4UKyjdGzAuQr0iKsLjhuTyGHjCJd5G83rjpi2FDjJxZFeGkXUXF3Ph
SA73edT5iXlCQv4QD0VAk3zOOTUT7XNyxwhkwyLHn/27hyTyzSCFqCYvfFcmkPto
p6mkcQl4GVBsb4PKkErZ93h025VP7OVH+QIg0fGdSmByuX2ek8lShPL3NKXBROii
BhUrPCEyKFFWua03VFqjNOyD29SNqUOYAqa+aJqQ+B+kNYlvDtEi6R3ducClJ0iD
Ysd0ihLoElWM06uaHLtq5oX92dam8a2fqAoZk/OidXBswShhTSqE4cuOidpjX/rp
5qI1M6R8htgJ01UISkLcuN0Q6hCudBIlz5IjUmseZ/SR3I0/Mnlo1LYKP7vTLOZ+
USRmw6hlHY+8sc+eLHRdTq7c/F5BxFf2VTAhtfzCkkrqjgSzmJKh9nV0O+/KClkQ
Jhz1gi0EWqNOrtytLgGZUsl1xap+38pJ+M04bqEpiJw2RM+juKqdyCXgmb1J53ul
v/KzkzT6u0QXmf+frLKMREM/UL8cooyPj5N/x4z3/sU+FWGNIXeeAsV7Mm2lTRfU
iJDV+iK5TGPKE0aD/GRyZull8qMDSM7KrJ5/i7lIqVUZfeN2G37pt/3qRdYDOw8l
PaynkQWWTS9twerpU9+Dw+b4PVWoPRpny8kEFhagkoqEPvbc97r4u+UDTj24ZRm4
bBwqtI6sSANltDsji/Nus8Bnhe27iqQBXvROoLdEH074cQuIUx2QzDo3WWiB3PCY
LnglxBJLQS+kCP4HIyT5hPFb9U0oUhnZFTi+u2K/MFadrMHfBZk+11F6LoabB+NV
DApURBkdTsoN7aLHJTg0QTC7DiJriOrK6u0MiFxaquBviknej9a+qOaUfi2J0rLW
kBqldGXs8DDsYNRKVSqrsbQY1FXpxj5Fqbh0hMuGFugVVFozwhbyxWSv9vKa27fQ
QnzIb9avQuYuzFjCpuy1DHdXskDZMXcYqmmqzqfZJJnEANeh4PCUc4KTGmuwmBkk
U3xxTLX2AE9wZoRt9jZ2SN6nyDgqiYYvFqtZrYOol/EIsRwPuXFQ8NrVeMeTn2W1
bvva7fZ6rGAqO0qkHHNvgImhgSV/Vo9ESxq5ddNO//4EsfG/EMBnxpDI23ua9iRi
LaStzX32c9f7sEk2PDRJH+m4PiZWlbGGmUAoM77pN1dufb5d+IMwrZfS6LC7XRRM
jxZJN78ZohbCOoaWYgZQ8gLN/zAZuSXT3NAojAI7vPzgmgkyY2z8edME7ZH0fN1L
XFgiSi8EcCxVmcrbKaeGxog1EoshK0lUS8UHLqq29f2BZMVMdB+Z5xNJhhAyCPfA
TCyZaaEPNC3vEkhampM/TrFesHVJpK0Vg1V1H1vXvjq0pLeU8RU4oSP4Z+vnu+TC
bmhSjt1gecNRv+qSDlI2VSVZhc+4QKCLztEU8NG+gwMYCHGoGOEpYReuArig3Csi
I8ooWGtBuaCZVfgGvD/25LyAJYmn4uy//9k/DbV/qUzgeZklNewZQ4NAFWY2AUTe
XnLPOkBsqZriNpOwMr3FElnz9nisA5pT0QOPTA47id2hnJIPgHLgzkfHRBsVqKIK
0DgNo9NOXjjpx3Z6O5QCDt3LB2ehgNP7bUg/YirKr6q7T83MmEsNs12ZKs34kmzN
yOUEKEeTQ/UkY0gxfezA+74Eg76y8v6PgCFetKMrhrUefkUWCTYfpUU4VnWBJFKb
Zl5zBvTgdZBzec3Cgu9pkKSwzgRfFuKJORkQB1zN1GjZaiio2Cmnk36KocDsaFkl
o3eQZC153sMTzKdq2QjqVu/lCJXXZ9AkUS7g1sFv55r64Yh704HtU2UlsdURURSl
iyxjtleyb6VC93N7Dtiu5tQaoipOy9XiZlFmm1nQiOU1s8Tr5xg4ex15MuaXNnJQ
ThVnhP6xBgzYYUDi8khV1R4hCZGRnhgcTa+fiuHnuA0DqrvGwsaTXhYZgysEk+PN
UXIRXJiqD71/ISvBvI5fmv6XVLxdgU8kM2YMWHcZofEIkKcyQ4JfK2Uk896xsSua
QnedQxQX4JxVUvEll+0VQACaZyPtKbVZHkj5yNK8sNJ/PSf7tS9aZbJUUQOknWJB
9MedmVc2uFiy/Q06OD1qxf+8WxREPdLSuGRHmhAUMXvpqUk0OSSbFE7h5xzyzUeX
7vNUxNNiuOcSd5xYbS9YSg29X2lSnqvDI21qUz5xdrjtqscFASlbknsvYMEYfru/
0EHI0uFqiFLfB3MdPS2tS4KBUVKJK2Zm2YsuiZJ6Zwf4+zCSVWB1htolCN4irLYk
dNDbK8oPWw+fdrWq8vLG01iQBprjuRtWh6HGOvGgom5msXu3S7YmhWXTnfFdLspk
eYqgMJ8o7g6uD8y2idxjlh52c35R4wCZkUL+ifwJVMEkTWnTV45UhJ+pSptIFJPa
c+7Z/c1PYP7NRN9e2rBFyYDWeNegkyTj02DVEM/l8uY2Y7K1mNMVq01Q+iq8fwtE
PG+pKtnzupPHmYGS8276Jle00vfAAJtv2LWuwGhe9k6PdWBOxEoHw+AEvMNjk7DR
uJioC2BhnFlud5knPTOVlkCubTCSALRZeJAOrDCaZHeQ/4k7bO/MFzSXxWtlXyOS
mAsTVz1qM4x/zOg4N5UvJWZWmp1pZg1hULoPcx3yc/IHycwYXoRpGgcwY1IywQso
fo+/0oh8UIAxcck09waAvyGXqef+bnTL2ltRfh+qMHwi8TH4ypd8J4TuyBsySFew
QS/SCyhxJqfKxER8gCNv3z+llZDq94Sf0ocIDJlv9oPipCzv+qrgz1LJhbyuBi0D
vWqobrUvtW4vWJxEH3vJJxKIVeqlQrTP9kr0Twx44Dh7ydlUQFxWgoR8Z/7WE0l/
3DDQB2cwsol/K+ggb8RELRmdp14pUCySaXnACvmb4c6x1OEF/TGTFsSfGgMDl57C
4JBDDmr4udRVHEUH/xmUijW2SgAKgmlb+x1RcRb9Jc+B4xSyldWm/Y0S55FjStmb
y5e//TM1u+K++QwfbKKNgzf+o1k0211iGSQZiL8Ga+LiKkwvn8RgRBmLAoHT/Rlk
LaT9qIcbjx1bTh4rabqRMx2+ghxqUZDFLXcZCuulTN0Ooz+ZFSsKui1hJlK+hdI7
hCTRcR/47O+MImKQVcO9cGvoGzyw6ianLbWdpFejr+XlXbrmYiasN+2tsZX8IvGt
mbWYbSppDWh2WSG4K4471xhAVFUxNGbgtGP0cjkkY+dREKltJAc2XV3VfsUr3ajV
CrqRfhvl2QD2bQCdvwBNazHHCOS6FfuRjTNQ4W50Bu3I5dB7qYtZwBC5DFlP0sgw
4lhL43QKAzRq7gUGy9W3AVISLpiGp4tgkwGj1pNXRnguIRLpjYzF54+Yjy6Q5tJ9
UQpDLFCaLOTzKJNNfLZ7EMm4lssKpYkMDpkNoupZwux3cl6/tPzZHV6XKfKhGkYA
yZUdpAJHOVHJpen+c665Dn1RrBuX6bHYEPy1xdroCKMrv4q4auQRRvrZkG1mp4T4
f//doHsoyqY0Yfb0MnTzmYVfdDw8dE1NKYUFn8QK2QL3csbKcAlmr34gsVpuAu2l
K3lxUjUBAexPIBIFfXPdgHvrnm8bPy9oz4zuUrRvkcmvs7NOOppkvfleoNoxU0BJ
iyyBe1q8p13fbfRADLviQcBe9KJ9ZD7Kemt8Mz8ZXNV7uhGqb+7VJhByhVi++mFp
/eFit1wJt8nUqFaXk9wPu2dT1y18Jko73u71/jNmCzJbownRm/HCRLo43hf7J53W
souH0DVPFWhssOPz4dmweuLGQ1QS1pNovX7LpMegnhVyHjEbvh/WGpbxIEd+tHmX
WvDFoP4yXbU4UXvwQ+6BfqEG6SheeKcknicPw10tzKw9KdznBxtpSLJvJPTThl4r
bOG2EppFX2+stoowX3RY1Sdp/i8H3J+Dyhbs9nDqLp+PDwXLQlpByX61rTAb7t2y
9/sVX5SRnfQ132Dw2DToFzEF64oCxnwJhgusiDpf6AOPSaMs6GpZhuZ0RBiCT3/p
RwbpxahV/rTAYGFS17rWx389JC49BkxRM41AUK1/Kcj9a0Kpw8DDRONqVHWdBP0w
CE/XK6B5nL3JJIbXW73pCalSAB1OrnlzFuMXbc/h3V3umGPSWtrI1WKvC9u/iT5q
Us2VXKiXZb5Rqrz0jUkL9lO7ykniAja/CkgBZ5JL39324vMYnImQU46zzMpHN3/e
fkuQTfOtlp3VTTm13whdi7Lcc/BWPOiWuN53RUTieyWvtMLclAgjYivgoczgkHcd
HXxdvnWSZKYTdtHcAqHhmNEmOKD0RpQCrAy8IH7cU9YNJhwcBdkUk7xTR+YPgQ7I
OwHVqSpuBWJKU1z/ZG2jZK+PKv1q1NT74BQaWJMEfwoosNOBkfnnIl0tJAFPmtNB
R18eJ9AmCSJBeTHTuz6gcL5vxQgJ6kESEfZrCjk+yPuesk5kGUZxKjXN9Znl5lRX
Fn24DjCojFvHqvpy7K4fNrcqC7ESaWPRQQV4Zzj3fljXXZ5cwjJiZ9B+gYIu5FAm
uOffWThS62vVBC8D4ap/C0eEzdDQZ5HvUgYb/7LMSaP9r7yIrsNwjz37d2ig5Ky0
/mwuxVZvr5WRxmHhmy01FjajHk/ak1t4BKo9Nc5RmkAlNmtOud/KTI74QDcHCdpY
hipvHJfEtoj8gyR+6NF07dS9Mhc0SKpoApY3PvN0sjkDy2ggfiyxJjCprrNAMcb/
OghHHu6yip2O8MMDAcp+fRAkezOFGQcnrubck/Q9V4KIiIuF0IGe3wwQKCpRyHl9
jrOzdWItAnVue93/6VRbZSvZbQekCwFlQsqztDhJKwvFv5xZiGDpVRZjB2C8RSWA
gmMjNieQpyti9ph0w6ABP1+MaBa+T1Si/NZfGv/eFHj8UT4JKNr8qbl0EUpJmnMX
tQQ2nIbqTrItOVTSzYWiKWP7p3uq1srUPw591jYefDu6BaynJ1ARII1EWiJvd/8c
mHP2e/L76u3CJSRESsMkxxcwUkiAANz87PzXk3V+Ret3haW2+I7fCuLwn0WU3lGX
zSQawr1dw861ejL+v29d581BxGAGBhmGLAdUMqzedXEeJdrUaAW8JsXsKkXDjTq3
iRNClvGmnCWhVoL+HiCbtFw3+LXUEQho2DagJ44PSAkRfR07E+GKWmXPPRX0C2dO
glnVYIWaJAVuOyVzUnjRcxBcPPZTgy1jrjX9iFU5WfzRzJLu9UkdU0mks7y1kWw4
/K9F7jlwL+M7RCnrAvKgGSqlBhoALyI8HnGYLQSfpddooCAsv8Is5FtlW68S0OTx
UDF7MPGFMMHvzkf5PCADmUjMfpuvD8ZS7OrQB9Bv4xb3npr3PaecrpKl1qwT8+eX
Ip+IGnYSPwGxFBJ4RpiNa8u+NGV4uasWZxeN32wjX91h5Tv0DysbIfzfYC5hqKF6
Gor2hfuF+TsoUT9GYdS6uPeM7Hf5Gnmga3SqAUTSYwyDQLuh2t650tV3x79ajb5R
OTp/+M77MM97tOrs6u9g30PXBV0eqqi+z07Xgn4dGpXBZwKBNkiAdXAEDqzGD4IH
wP2LEwvm7iT6C3JN0HYiFt6cA4XRH/kytbQdzKgbvvg3yLfcTSdQV0i2T5xI8Oxy
p3n8g2XEYjoKr76mBX8xBjUkpc7mkvfFpdnDEzvj/LfkWNlXhY1MAVtKRtA0hvYL
TI+/kEbhbOrLrBx2SZ6pFi/0uc6SovAJlEcK72C8aSf3UGu5dFaKYZ8l9Qp3i4pS
fPKX8T8O988vFn2nNQDiCZ06sp0/ly4URUYwc4C8rw6WADeXihUKjoBfY2LYR9Le
nskADPl5OKiE5vmWaUPi/X7e3x0AlPxukeDjtNDgDKdNM5iuXHqRykxjfJlGW2D8
SBXQcxNSzmN3jvabu8nHpsCN3thKfPyzvaBeJVmdvekQDq2hhEtHNUaI7+1sy1Ri
D4aSCOlcZVqm4ptcnO2BxZch+kQoBjmyZzPrSIYhejvKXPJYmcfc0yLf3WIaLnA/
nRl9oJ2JB0w9J2qa1ndYFN9qSlsguy5vsbScUaoUnqkgyWgl/vRVS7l3TJuOD0wr
uHmU+uGUbhWncMfnehLctJ4j0/jPMXQH8ivHvPRHd6NQv9urap15fzgp9p+aCUGn
EL9NNFUASyALaJ0ZsU3H8oha56ZVwpGLxzIgaMPbobexVxMnpwxRkCX1tJZms9F1
VVPU8TC0HjpoVPBeTQhp5Q/ifD4vycUxGL01FcgzUVWJigVhQr/l6j5RB31IK4xe
VDA8Y/n9ccZQTkJhrj+aAclxsWrSyi9Lg9VojAvnNEDBlzcaDzkhnntKBwXFRmL0
PtXaROdY2OoEQxVPBY+RA2/L+bmJjpJ87wxkRrV5wrX+7trnAcYLKsxiUVdGtaVN
tBq3S+e1MmuE+AF0zfuR40/bf968Eik+KQkz7pBbjgZ85GlK78jQeRl6MddaZeQ7
AsfadIan3KOJ2IBgz3AkhHm9gwy86zRQiZzpGnWeawHgWHfa8jgMGcUOyU8yuPnw
1raMu0bYkB1Jung/WwPelO9J5AZM0pYnEBNeb52ix+uV2X0KR2d+4IjiaG/3f8Fv
XCa2bpB8Rxl8/YVPSCFryp0FChb+HXvUuKG0SIK/yjqbhnQMqH9zq4xKNS8/UgwU
uz/3xBhhVgr1Jv5IQ+AVtgPYHEHtcY7O/01RUEEqSQ3tgewMCq2WG4kYmVGKUJpG
+3wfojfjjgG90LKJJ0UapEJPtnxUCox9VsaGfZCN/BlcIarMZrsh8AAVF0H3ibGt
TapoVAxlFqERqfwG6zcjx8XlLDC3uUgS1zLa5+Ah38NDioIlERz/Z3gz3Ii+dg4F
DLRTg5qe1fhj5YL8dORWlyK5IM08rF71VU0LSZVrjBrF4+ULQs3J+v31R17lR7FS
b9axJFCFtSEw2B3XpoFN/bsHvH87T/VIhvvY8tRjWRbYyCFnFpw9Ww19cv5SkBKD
cD/H0J68AKzstnCd0bcspT5yFgLqW72mpYcSU7T9ykQfXwfX4GMI6hDg9dUWZKMj
8CA3HKXbm57IMZePdP23JoshXCeFaE1W0sxrRQ9H3rQsM/24Rdk6BtvKtge2JBia
FWbKJ/T3Yggr5uU8Kkmnk9hjNsepqhIq1y/jg1wSYvzAXb7kbjquyjNF/X70xl83
w2PHXECmbPfjY8vThFbTyTX33pROnFnsaTIr2OVe9tSqpPo4hbFFiYvzcseG+Eza
VaJFMO01CQ2i9o1l+OHwwYUJcE5WWB2Uz0xXgHqwJ+9FsKbZ9o/azcF66DxLImn2
GofUzUl40PRPzz4qUlwOGd1hC1vXHJH3xhMqbw+jlBTtTtbxl9zR9LQ5xixUx7cY
0DCqjmsNAZSGeKD5W/MxogJVVjDfBNG1yCKBRBclZDyV5Mg9YyeSD5V58uhBVrBF
Wkkjku7SHWx+O6dPFxn3JqI9zvTl0MD2b1Mx7LVSvE1mYN4xcUunoJ0zzAUZx7n7
sQtvtnx7moC7RzoClWTEX1Z4iZtpJaB92uqMSsp+oZkK+zn6Ap4VHUGtCScWQV8N
/ejYNz2hPanGPow36xCG0e0rU0quC4JVGcWNP1idymZf+gfdWDlsgPL38Bk/5KQt
Bh+2h0Bost/G+0z4qNeaE5u6EO9vFg3xJe8bkqU7LTA74KnFj3bUox+0EQvOCRBn
icWQLayOo18Rs2wJIhqWK57VlJPhau5kHnnLM129Aj0d96GVddLIgaVTFnbPqorQ
dhh5JXoupsbfci0Kk4WE67G7KSmPuJBP7/KfMLswDGbB2dwcB2IRfWntpoFZiXpt
PDOb79ngXde4Vzls+dadyiRSi8dUjyuLSbQPx1ig8Py0/XrlMZrja1qsJzaNF1O2
Qk+cfEpiiuLl2SuWvmkQbUNg9ZkqIWwMqQs0OUCHF/W/YDnAprjPiyBnpyQsEcGW
f/heVNg+IGxpntGXwFhvW6IKL2BKyIymyPfErIo+tOfYkIuFcidcVx84F9PWH0wR
KIp9ki7Kmo1y90drWdDAsuxNlLnF8SM7qU8XyRKDQp7ZuOCeyYDOf29Au0EXkq6C
g5udn6cQ9gdYWDeaRuzB4Rtvnmk6ANIPEIDH7y5S3nsbp87k7gJFp2CF/v0i7Psf
uWQT0CobRjgUazCYgYYOhK9ggr2yUzLjIuO1PTjxNppreCavHkWZP2qIxjB9m+e8
2g0UBCbd1sxhO8yul6tTt/WgffHaeyUGHSGo4Y0H3DNPT0m0IJLjAv6h1TN40xIN
XqzJyUGem4JSczxbSX52cOm5j5AHcrEPKc33DaBCNKRD6maLWTPG0Vlk8dUo2tT+
6VOm/GyOfGWx6YENdWyF6mzu4HPfwFuO7DvlOKasQxbUtfbta4Bnzn1ax1tzW62l
9clqvZGhLRoiTP1pe7DBS91R46wy1AzWi/hdbphKlKMHylYKXH5mKOjVjdpyRT+U
mhWnEc0DiP1ZuKad+V9f4RBCGVYmbLDnsjIT1ypC+ezSIrH9CTzYyqYLmTEMRoV5
4XW7VPTgLQ4DOWyPA8N70q+V9i+sghC5mg7JoxRsE7dx/BsTd06DT8pKPo4/1C8Y
j0WMsc/37Oz13HlmM1g0l9XsNOZETqK5uU2U042rzYP3K6OgPlQVDHPBSuukoJ3r
rjZQg0Gh9l3Bah/oLBh/x47ZuL0OweqWJYiKcgkGMHFjYyZkdoLi5f0ONSzgEDf2
54Jm+PM5JrTM8odhmuAYvFQl3upLtirNhjaHBHCktxla9z09zLoi6IpJ9GTLZCVU
eRB3rH5+8AEvdfujWk4d7zet2ZpbAJbe1vOGQIyiXQHWcrSDwkfRTupWUxJbX+gd
iY8fp8TjdQwbjuVAoRQ4esG3RmxUTMJw+3t5LoQmS8eVK7qptPPQCxu7J7t2qlD9
zuYIJ92DLgC4aDsBuciWnoL0W9UR/sfseEJjAoFb/YnrS9HmuzS+QIJgdkHKYe4w
BZktnGwWOdzXisiyYpydvNvSghfdnkkIqXfCImisO531+ymHvGQCdVjYSKNQuWUI
oCFSXZ6vhSZptMNBM58t+gyqIBTtRslxhkysKeCCvZuYqDbJf8ltxTG9Nvbboxkz
ll6FkkRyTu9LWySRRH4odr6DCeFWtv/YVTCsBrDvgv+55livF+AQINrIFASLSc0W
864ymmNy0bxaFiwEibgXwV2OcKkxXOpb9YW9xATYDNQBmm7HmPmTuePE1IppZpjt
YfMpOornXwBRslaPYYJIEXNn95x1Laigw9mWJbn7hZhT+1TD5J9aXb3pNCEY4p1F
Tn3nFG0MNQyoEq8W9PRLu4gArfxSuaww6GjUT5Q6WPSRxYdy3Zux+ADWoLCEqTQX
I26iG3vrjUwcJu5eylIwxS5ZW7C8UbKI+PkAUcoiqAiMIduuOl9TkQmPslabF4RJ
pjf7qi2VK3h1uKWZ6Bkaj6QsBLcO0y64nwebXQYMPdWkw7LH0CmYZ/O1x31vVmST
hVyKuK2ANIPPD9cXnzrx6dBUELczVP5iW17PmrwxvKBhvdRjsWJ8yODW+jxWD/Zm
2HZAGTsXgl9LNqixuEGQ+6iSLvu2u+V6B04TY73UdckETqvWfmnKmOzqsk7jITMV
6kmZKDMpHGWHg1tfNprULNy0036JEInT4jFsYqgZNCWfdTzmE7D/n8pgemVuLacJ
Ai/705GfUgSTyc/EwAGlLV5ALkRyT9gSXujOrpAQoasnk58QO7pqD17Kn+Yr2yfM
aP9mzJKRArD7qIKfunHRS4jT70lqHrSh79jUFmQfSHkZL2HfIq0ayzk3pLOy4Eb/
D6Er8gKnt8jqypRus2svNrYGYt9xMdrKKhCVhyc29FzTqs5sezvjn7Lq+t5vbD/t
NMgC/rhHzZ4x9sZtJ9I5O8+H8/mU7vwl47AegMCekiM/ZUJUSa33mKk7cftzXyM+
JrEzKdCuy+/IBif8h35GO+lzKEsnLJADlrJjck+Kpi6I5db+ufbQNKaGItc2wg6b
UXcwgRrAbHlYfu25Z/piwat+8vKpj1MtbV6TVzqr7f01ybdVbwPifHHx+DgkWbHF
oDUZd1jnVmRdQNbmp1B/BH5g4rsIM/2N7Vg4ZYduqqnF8D6Qn33bC++vpGWDX7sH
z8HwUoKBjoVOY1hoAkokveJtzW928Lt4wkJMQajFl4YQDv9YH6MSDpdHELZ5C68a
HwZQg+t8Ex8AiBvqjiHXeJALRmpUf46GU1hJyLFnQjtiXKdi9nNtCvUx/sJpOCXB
BW+1F8nAYOKDNgDc5HA7FSYYgnhstzd3/QfusOCB/eBDWGLUOcC5Bap/5vsnc0XJ
GCFzhc+NY9gepLmu5o0zr9/adFwQBi1Rh0OgiiB9AOhAy6/CMuvMR+aBIE3wpArR
vcdtOM6Jdr9ywWInbVqxqJRbGQCo3NBWisVo5XSJJrRy5v6mVdW0Gmnf+gfPeMby
2lF+4p4ycMYBnWkZV3xAlTaq2JjAb+03rR5BTSv+2IZhi/1QukG39UPUy2pT88LG
VppXCLJ0jM8dnZRySWPLyUoks7cqyaZyZSWTQqjl4ikzag0OyKQ8nrlTMX0Sc0Iv
UfEoQ4R+Fr9OYlaojss1dNwc2RUazp9o8jQpcmZjf8TwQmg6hhLYfwqlsl5vxxwY
4ioUvgCoGJiWU+oNnQ1/I2lJvqcnWJINCLc0JZFlREXzLTRTc1hWNNGeDr9+kUQ2
+/AsTeSl1Ve12K8xsL6ZFQIlXgNEG4uFVVWMtju+D15+dVlHsORXoXpDlx5P/rgB
7OqYAYjWThJxSRcYrNjQGRzUfLfJ4MkMh1rAsFTPPxeUWfXYDfTXTLLLTvZhv8Nx
HcXw6MXIEkMOWtLnuZS05gy7WRGkHpekI/zN28pvcJCmrD+V3D/iim+Byt7Lyd1/

//pragma protect end_data_block
//pragma protect digest_block
WB7ZmCkyg0p03kwREYD/KAycOA8=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Wm0RB+aEJ3rH+7Vxkstleb06v+tWxydBfM8Sy4mnYjbFD9Hcrv3B5PTnRG+YfAeA
61vEIPVdH2mookrbcQXWJ04+5zmnva1GUj/K6x8PWxmkgOumcYcU1U/lIGPeHZKx
bLwYkIsz3ura+ICsuS23YA8Ad3kIKV5Q/WL4iqMQPP0HnqT/YJKCIQ==
//pragma protect end_key_block
//pragma protect digest_block
zq/978CCnbeRz+Z68/qBMAco6vo=
//pragma protect end_digest_block
//pragma protect data_block
bXW+X1xYz/jTNzGvc139MjuQjLT7o5iQ2VI0+EuEzwT6y3qqGH7ohjO7qmVFaE+E
akMRPVbJY0pQaw8n6vr0qVo1Vsf5kyezQcgVYi1RHDFJiT8uJ+0xhhk5Yrl2m8qO
pZsbgUd2X5FYHK8Za086l8fMVy76+ewrzTqxxy+4H9DIpBFKif+CdDL6cQxkbIxt
ZBdWMwga9zWgsorujMq8aYno6Db2uo92OIvPhZz0MWSlvHOgzLE+8SRKt7i10OWS
Bog1EjU4CcH1DaApnW3UkbfGoC/x3lGHEqnaRXGjq9y/j6wKRj1CgB/Vj1dKGoGW
XbiU/JcwpJ0DPUUsPmOfygpRBsADTdpcHsmOwLMCfONYt8OSXAFXkUTZF12J53Sy
XyjBYzvPa6Zsuxum47JCAXyZGd+J9h+nJryRujylCDjbhBqg05ZegXTa01B/AzAi
y/lqgspctZ/LukPcQnSOiTgqfoHJS5a/Y7etXTWI53i+F5h1CCqT1W2kkJOGpIvL
/kemrd8UiOvvIyqi5tfLiXQrU/n5xpyGVHV6NEHsyHxHw3WCCSVCnfMtC5bX05EC
NHdwxpHWoBcFOn9CSrMqV4hekQ8aU8UMW8Z7i/ELmaL321zyphjHs+6E/UMHb6vV
Ejn40cVDifKlk5W9dbbHY3DuJ3hnbrulFn5e+R23/iR4rbshMPQxxCffYZpasuwz
Y28c7v50Nq4b1OPGT+gVNXcHhl1BEjB21UVD3H7YuRO3KBY9SDNXKeHSskou7IMJ
v6WVroaF6OZXRyQJBhPS25R/n1J38quzCHMFhkSo6gs86eUa+2kze1jCPDt1zVmL

//pragma protect end_data_block
//pragma protect digest_block
W+L0AuoMH/uLOG5LAkjJTsmcEsQ=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
xolh9mNyXeZfXcJNVkEBAFKLNIAaRud4qCFxkkoGEW0VuVsaFkj9QemqbT7x86oo
28ep2ZcWCYMLmbq1CEhw+W+EoCjmgezjeBzdVD3sTZA5U7klmDQUyEMk0jAVEXyk
fJXsaloc8YeaI2ZI132oxU/Qe0IOZC1Gt3ugtgorARHuaXKNMu8I7A==
//pragma protect end_key_block
//pragma protect digest_block
rOay9jSemdq9TBpVl0d8IBiBsXM=
//pragma protect end_digest_block
//pragma protect data_block
mnGJpi9n4kItboiKz1Ev85vnw8fGjEWYCZFp/jTas8LZvpu0PXjURjvhlR4ojrHt
XPJUKZ9SYU5GjJloToyKVP2oyR3ChXlW6xwamZfMfWm1gsGkrNjtGL/C4YhjzutC
p+CWLytXJNNskyuvadVP0V3hJsgWdYcgfCLraR2ONgzriDCRvFkBBZ/P42Jdde/G
8cgTc+eBMEUb3Fd5QLNH0QjnubppOS+1nSJK7t7iBgxyJTGLZ+DnTIDdTvcfj04K
4PEtoBVMFyWCNnyWRFrAWflV6o38nla2v11aSlkk+4P17ljuVljcv5P6WQ4A9sR7
3gOQP2K+vmxh1xl7APEcZxI1HQgeZAbzYRNVVwQFzn8juiGB9M1S0fFjh7Zha0mk
rlFvRSU3EngkBl9ucur1DVW4Fza8ZjDOjDPw8gKkO8XjOoMVsOkNo8DvRCCRRDgp
Za6Jue3++j2f543weRniWFXuBtmBJLETAbmDfY54gZlYhyA8/83hXb7GjJWkn+FK
4Bo23/M/qmUlZ9P1LdKo5GzSlH9IhsfkcYEDSpiOYUf9p4avFSFhgRLUOWheAPmi
oB5nPbKWcvt6OQxUq2aItlq3ur2L4cjllpICyw1ElMVWWBeQdHTfqRjhYJgkkUgT
PJ7jvYb6WrqGg+BX9JdLtvI78ukGbfJMGdAJfgegy99wSHa6AiS/3LSAzasiOq+k
WMWGM1pxJGScROyRgkk1a6SIuudhiUDcEnFJuz8amtvi352MxuA1VI65Iw6fBYU2
MKAUdUqr+21bQ6+KWYNzTqaOYpAM2JNR9t7OYKLQZCvu4YbnxNfs3Z4eLzcUbz0T
Lnwy/QDkv1bAbDENax7MHEKtkQfCtkNCeqBBx5cwoLkEhJ1AOmd4PLwrC0zdJJKX
0aeDiL/fEAJ7u5jRvcYUKyGxjcbo6m16xuJyXdYEwatpb4r15e91kaYi2jeSu3FZ
cR7YxRZ99CeF4bMlFHOdyzaDP5IPrETfeLKo9V5hhPW5jxd9xx2UcHGHZcrMolw+
kfJJ9Hzbvrq3u7GIfASgAM5VVkswg7mneMjfQrdqnIHFviS3mO4HWImlNZzy3bM+
iuYiQVOe8HsqF2NqU5JSe7aXa/pf+73aTp2Qb9VVPPAB0bMPsEOtWr7fybVWPMlM
h3miPQpZ0t87ZY9mtOZhc8xWJxl3WZ+/9ah7OGiWwePExK4+DxAl1Gsfa6TiBSsb
qTZAn3d8HoKdouWSXvYgwTbXEAhXcdeFg/nOBYH7d2ODS5bNkJ7EJDw9XHrc5EDn
iBOC4qRJojnIoMOmvmMMarx2b4Rsl8SULOpfq3cS/4Cu5uOgVRcijC0NV4JOkp7A
ii7O2N5lAsbkKPXM7ZdK9pGomPKVDWMOkTObtRYucXc1QhZ+Ihd8aAOQHozC+XEW
q1h9dQevrZAML0TjY/vCRUyIF9+HJCFsp/6Lm8My0pYpFZlHytt7TybSCidxyl0I
MK93Kj6aIR3aiF06Nm6ynx5XxQaiSNVxZHmIZZ/zG2dckHGLKdETWDYZdItyV4vs
LsvdWE6fGP4OOSoEHrLdB0dCwlw/MSZfTSbfqzruArqvoVK2nenN6GmDegnIVrqA
lSbxhRowY5OX6unOdQvNhyDX0NKn7uAleB3mg7/fyb+yg7Jn0bEOJEy5VIfUPM1R
lA+OeTaFdolwDaxE49qP8ZxzV1Yhv0OevpcMIzSqFDVs0S+y+espfZfmMmvAgpqW
VUwo64jhWOXIn1oYmeYw8SiavVpziRfvaUZEsIO+S/TSPh5VcoWgL/mGw5EoedTj
CJ55s/HP712OlgrRwYa0Y8bHectjWqai1t87IYrHBNLpJDWABJ/sP8CeXdr3J0V/
3CI04bhaHNYt1fXwbiMXW9B0t4Z6hFk/ztWoRZvx3N9WNZL+a7S2mPgu5eh6b040
lxiZJILDRfLh+BywseBCN7u5Jat4dJyUIsrsUZfbMD0InPtuksdq1Kw8HBy9CHuK
UDchFIxmRYIkEH3zUpkkfWa8a7JuAFFBsr2iHduK3D9Ufl22msc1f/3AvyLs8AHE
IqLooKP+SREsbzbaEBf0hUKHL66WoXAYZGQrha/zczJF1fEiK6L7P/dAH9hEnk58
NI15YXd1UCHZAPjUBE8aHCYxcAm5xyQ2RtruzNo5k1kP7ubcJLbQnd9MWIAnAKLr
6Y3TrTWsqdkllcXM9b8SJbj9TJNZJUbLVvE2o46yLwBl2TFb70JtzcXVqA0xUduw
vgerxS/6am3n7UmGjfh3Ah+20Eau8KjnnpFf4IRG/qdHBhSUj+LalLiUv74V2qQe
PVw6hyzCT7iBpewcudFMSMekKocLQz008yLN/WeWATiVbkCoIqqWaNVsCg7ExZnY
zRm77dK+q40m1k26MRQUmCyD091adI8O+CAxYvJo3V0/kxHRyd4EpAb3Xc+qN9u0
OLw3o8hlz/idMtowGnGgfUZSm1ZFVwFuKjKHXEUviy3bIvbiOvkGk/Sm+zxDAl6a
Rd0aJ83FzqCv0nbXe4A73aKzKShQXpN5mzRzurH25B3+sEgZaT2czZfR0OrzCWOs
MjX4SwvO0Nrp1g+HtMpJeU6GfwPltrbGvHCbND5isMHsn1iw8uPM9Jbyc8FbAtMI
Bvp5xTw+t/hVBUYXS9Xqo36WL3NMtZ8fhXrPwebSWBVmA9+TQhZPxPJyVT/Z8bp0
6sxrERDsmE9op24YKeyhWt7AGEmTKpQVNaW3vlRV0NHg/O9iF+LCVWFnzZzZl3Av
YbZU0/QsfXsaQX17NByPQnmUbmlc1Daybnrj7L+vDojcnK9MZAuRdmASrdpVf+eC
ljw0QE6Uq+xP/bFBBc1b8Xj5H1MEmIwmjb6ahwRC+9ry/XrRicvxRKrS6IgMs9gO
w8Hmw3so/s0mTrB6Ic1qUnXa0brzdAQy5n/abacSMY8sglJMxdVuzRFOmrgwv1yq
Rq7nd0tSNF77HQWCl6HNYHh0BuoaIEVe/q9gc3i1/yL3c1kZnGa0kSzIiAfhV4ey
OIYRc1A4XzeBW/nWW/EVIQ67aNV5Kx073PkLnrnq0C8l0US6MBzdkTP3rBdeRUcF
fhxBotDbl61SONZqg1oIfumWwJ6QSFJ4kmFQRyW+crSqYfKdAhxHg5eNYLHXtZa3
hSYSSai48+YjuWsa//Y/H4XRLsNzvZc2uC/POqjvr0IThplDz0dGawJDk/yNnCG+
ZAZZVDCJmw7Dhm/Xqfc62k85Qh8wXN52kwnyQ59ewel9jMEfjkI2qBL/w8gez32s
o8sDdw+0NHhnUQbLPjDlDRyEhkXJqS3Cqkcw96b/PzwWAdYXGD9+f9DvPkF+WuJN
jFPSb/xoRdGraf8sebDLsxyb0bWBUqCFua/XdVSzexS3ZnkakRdnd1pH4BABQuuL
u6mbzWQUIEgQzM29wfEB197sTH8Tg9dV48H/J62LO39bclhNzvskVqO7FNL9f2g2
AowmHvX/wz+cQa3g8u2wtRxIHwD9pBgs0QsC+DcN6NZzkjDZ76wEUAPd4idolTuz
78fzj4uYDJpZUp3STkJte8B/f7BWtRC2D0WuGooC1720FQEcv/6jjzVx/0h4deuk
dC/w9zX9AJIS8NS22VZRzzE1vzH6RTrg9sc0KyYbjrfYzv5cVAWo3NKxNoxuHYUi
AvgKmelg4/pe1LyhXQMOONyXV2NzffXgMz7NKpODnr4o6UNlrKIW4uf5HZT0IADy
P3icO/XDwUVjbmUvdz48XCqxMwV+v2RpgSkZNQ+0B+E1yIHWvju2G5P1lMIt/WUD
W7MYacCPZqrqsxYz/TlGO8q0gMBkpWcTgMaaGyz/anvy3SkXoIfDHNmlRL/d1mQj
aN2VkywfRJwVsRx2q3zPsfvdsasjF9Jy0kQ/ww9WwZ7o0bW/zJDNydrvVuoQPP6M
qKlfMSGFTyj5bCxHSJRaHNDGvjy+SXTxaD6FXveB7Ykb7b3t3eU/nRBUtCkZnJSw
HWiEZsQpnNsGJ2ACL20Ol8N8BtpBFSrfe1dpZTTklHcVqNssG97tyxMN/B9wPd7e
roMMbDmUEswfDR+dosjd6Pej1b3a7Nt9OSH+9ECjSQZceAubH/6FN1ge0WVpVJe5
z0qCzgzSNpI+YNdXH/FPE1ay4EvzXrM48p6T7ygjZfT+VU2OgfedCoTDRpD8gJQ8
ktzymSeWUEktsOlQUeK1D0g0nfx1D+lW6ilgKcKChoFYIOqnH72WN7rTyPYhB+uR
96mbYYYA+cMCEG1kc1bMlyLD7pkfcGQ0ojJmA4h28S21Xh9hqt/Z1BovKQgkZMU0
Cgfsf8QEdg8tg28/y7sTLBoo+1lxzAi2bya7bcK+Cw28nTvi+epl41X/b/orJYcM
bTH07PluOgYweR5ueMYJpAljNBmqinFIDtko2ULXDzYM7+Zn3H62u0MFKQeGGrP/
BS3PJqZrjsOZTqJX7GzwrjT+oXWqJ44Q1SXf9pOmiK15Jqtj0rZxZbo0hZGKlDUI
lt+ZsoT5QWiCTVVnwIlgwqVtHYXUwKnZDaqophCI3eBLmbp1nu66BjkzBQkBYtEp
k7HMVNl++3Ba/IRqQcZVNeW6YOScPCMt41JKIBTnuRvPwRUocrKtcpYkzozXTamn
JriSwKQxYrc6xYaW6NwpDeF6yJcdwsTBvf/aekRk2ube2WPAVB1We8leCOPkDE55
nRc5LzcJN50N3niyZFzPN5fsY+fg6cwm+juu2P/9CTiyi21EuxqeqbE6Zk4Qx3V1
QjCdmYfSUn+X5v/u3Ma2dzwyCPCaNT996R0WyIPDlXmGkrHUNpQR2lAoEFeQjG5W
Rw2MhFrVLjKeKSPSHRVUbOTVr+r6MDgauq8QbfNUlfWGDZuYaHiXmVJUmO1L0ms/
45rTc8hb1QOlbWOJa5ox56mLDoZKSSdlRvJ9oGCVhHci3FIWXBZT2gylNhBlEULU
K3+nfcC7hOLog8Vlk4o4X0vX+hviCMkPxKqm7llnjNyln/iqGu8DBRE3y/XbtA9R
19wodHvrCbefgdpvKTfMo8od/pQCB8vPECuK8idFMz/irndZOA3HLFgK4w7WTX9B
+kVCpPKflXdy112UcHGMuReCcXG5tVSc+ydII2zjP/koBGp+HuLBVu0c7EzqbYUu
fYLgIzjJv9ElslTKFbT7w4P7y7frtBXulx/xo2nZGRrJ//hBa0FLYMtiot8u7srb
4TgvC6wkMeICuUWztnbbRGoBdzGwPgApkhfZYbynH5EKGgNOSitJMZ3t2nBQt9hN
ASZ4VYgSOninxE6xJuKqpa/oVKexg+XMfhbKa3M8JQh1LXgdk1xGVbrtn2FeEc5W
dcAY/ZYA6wy33BEpRTqJWS+uV9LYxnT89vBjY0CUgBHYll5UUBSftSdvuZ16tG8a
Z3v+VciysqSX2ccMREIDjUptB5r4tWGYcicm9MZQRBiZfHhBtAEbeB0rA1eO8Lc4
UUCJ7eXwd/+iuiyfFlqO21L/2VkZuZLTL1ePDScfsXhuWKm4am4CHI/AjmBJZGcK
8I/cKxO21IV4Gg6Z2rpV5a3aNhf/7dEoBybTzS6eojOxtK4bR0r3lv6vpetcLXaN
BxEWYLxoxdnS3OP8pq75e5S81GpNstXlxGvfByZEmF8YzG9cnDD/cMVXTdziLa+r
EBsVc3QWzWEUuENGUOZy0/KrPE30D/zwtizeW7o+uH6njxTCTMJbIfP05hjUmQpM
1QCTnBZdxaa4FnqYh9odFX4Pl+tmvGn2MIfyTpeisRb030c2HAEnqlaLpTgDQ06I
4/CCH8LUt+dvO0H2VqizBNKqqUWc1Y0XpLuOY1knyhhobvZK+IBVpgKI4N095z56
VQbMpEwdc+pbaH6h6fAVab6IxLbQw1NY7szUp85478qgrb2S3mKRTo9b3JnYvckZ
hkyE02/5g6lJJ0fkvXU18S+TrqRZb3Bp920NQbWEzvcRrilWh1pBbeYMhXFIwp/o
4H74NoUlzvbEGW7mu4V4Uh1gL+NI4NSvarIc+E1WJomdUgRuWTHSUpRk5mfNQ+8Z
ossct5ZtViy3l867Hctn0B8lGyTUEDdaCUNxybDQqrTHYTLR1C1oMfNDAZfdEg1+
kuP+t8JCLs7K6+l6lLfU+UluI7hdRsWH0V9XvezcmE1AmWRRiCVgeBAkVimr9fdL
zngNM9HKvW7tXpEFN3JtE7yGdxoWvGDekO4nVaxgILaD1jugPt+ijCkSjNRnTe+n
nRhiY8z4D8AjOr6PTCCKFLpUzm84n1BI/xHsiHFZXLtGFKUVPdopnKQv/w7bmkH5
bwklh3TnM6vjtAgDBEUKR+9lYPZkLIhe5xR7HxhB8xaA9NMTOM8rdKWzDKb890da
2Ajt3zoCDjuqO8pxWod0FK/M6oyWerGz6Ws4OVW0vYoiRTsjH9/TKnbUsETBh+nb
MsR4Kb7bdpXhm+YH5FwXWv0mmeOzSdBZe2XwUuvjZYQ2arVWZvDHiKniQxtBQcBV
wkeAkQqwOimWTZcD2gMf1lW7EmbYJsw9okUFNGX63vbXmkthNEC+IZi6RM7NqDJg
fuywnSKa3obREdZAugylbo8qJn0ACt7i9tsB5Dy86B9NIJ6w26sCaRZxCan+4OXj
uCQ5jaLVyvZJ0o02Nwekm215QS5rh5bdCSFnfziK1moFUdiSDf7C7ThRZSY2Tw9u
pL1PUvd/4y2Lu6SP2bdpFGt5gCcJkzlnaf92PpEviNtcNC/d7ibv6nOgcGLYXwzH
h1ARTsQIxo6H9+VZvEKf7smPU1qq4HunJXncqRGi8vc3zFbO6PE12f8yoTOOLwBz
o/R7FfbC0I/3d9t48xdR0ldxjgtVKqpK0g8alym0iG2i7HbNIY7zOOnEK1Jk6yNz
zKhX0/JAvdqj+dMRLb1RDalp9fBnop8RuHNyjfy+bv4GnVAHRFBM9VQvdSZ8wsVz
xcw0kct8Zwox1NwI3EhrHPHUypWwE1SIQ8IQnTH1sSNAFyI8wfLJcNAa3jBHVIGM
SQRRpzmsv7baVQnlQ3Tz2FiDNCb8OvISpfuVvV7uUosblia+O+UWMTtnhFGDMpVy
Rp7tDtC1xahIa9A+a+zzlAVSWTweY8QHvC7MTqakApOLNDRqya65r9iP5wgNDx9l
YZIkf0LsCqlmV7Dmj7Yj+blaDDaV0dke05/Zi7rI2+3+FQ8UKqICKm1alQ9neatz
Sf/5GcmZwohz1LXSvA1hWjnBR/uljVEaQl6wizg0BRCVvHksB2XCt6KkSxyj7wgS
/ssubuY8yse9SU4QQd0yBH0SwT5m0rz1pYoJb4imS6TWL3DQ41Jx2RHoH4Ktu94T
YRq42tL22EucFWzVaHCIGFas04O9Wd+HASnhZrIMeDhKtF/z3HdUpW/WGqRvQ7h+
TLu51HCd1YORBzjdwRHCTcC1IXjRqKo+3AwO1DOMXb4qaAnww49rKIXhLVQ8Sl6H
UH2ofWVYkBujUc6OUET4zNMvqVB5uX7IkVC1tHAMEwX1DF4LQZhekIkLqu9FwwjI
xZBY7TgiVO9lq8xHrxiWVCMZWX93BAH9f/94jDNn1l6u1A/7TX567iv0O0ThbbYb
I2khZxGo9DISQ6QVqPvAgt+dYuqegGbv4yglk2+/bDA3/uODjCqqLuY12BL5pVl0
MxBaLrmnaEF1uy9iXyp7J22mEhfNVIsYvZWQDh/wi4iQAHTCaJqtUb2ZbLyf7TqM
njYZGRMyxQJFLmeN1CrCmqlylTWc/lDZ7cixON8HASmzDmevbGkxjmZQBmcZrzab
oqafLuWrwkYOUdNtQFWGRnRfBhLI0QIPvzNLDYFaEX76NzHAaXkKT6j10x1MmGoJ
+uYYq8fVtYFkMMCuMMjWxpKM/2DIOXBhg6UmDxDnkljhoh4RNZ5jYSU4o9O+4uVy
I7gguOxSsB+aaU56SIofkRnvqQwOsadzDhF7/mpy420W7rbpm1Kakx+UdQ6bkLVp
rPpEzyS7vGlEI9EFt43cOnjLSQ1YipStSNwAn94OjTHo/lLiHvGDRgXY6ZZuy8Vt
fxRK9ELy3MikgkpNoQTTgTyPsf38jPxWTiOH3CIS5RMCAJZRv9506KZoeGnR2Roc
mlruiQK3O5kKA8dbbjM2rTtMVvdzVUm965m5ApF1BNhFC44jDlepYpTJVgVZIPNh
GS8J3xHFTDsjH9Uuqc3MrayoReZ9zmSFBemEOp3e9JgXM+w3970sl/YK4GPLYUeZ
H73PBb7iwMz2H32u7kcnKiJ04v8ObMkgFyaamuaOnFXXCk2Ug79rHv3hz5RqAvpY
8bM3ZF5fBtxR1Pc4L2QR9GP21HAIUKr74WxdNN6FSC+LBjMj5BKrp+JAnInAAkVJ
db2A6c02LNjBRaES+mc6SbiO8CfG6ibfBHzSOcX/UU33w2qOoJLHUzZhIFrTteqO
4tUXLJEyh4KbNzDvBieIgILF+3NYkjFuGsrq+0Na+Iq1fxmoeRG+ioiKB8Hwtmdd
W/R4ONPyJy2oWXrvvA4vWrwxvYC3OZD23nrZUObIHsWGZtVx2F2/9w5t4Tv9mI0g
gIYgTsJCmDQXGGkt2xitbtT/NnxkxsTwrOdNVqXz7ZCRCRHb0glCYdVLFGhnifO3
4iQaVhKfQst7+wnNFMncbpm8ozwsQLpOKW4Me0wROGWAuwT9Cguo9O2fS8/n1l1y
faVNLRRfFnxQ9++VyUAECck+lTxM3rRMDG0OYmrTsg0uDMGOZH0dwsBgT7xTohwz
Uyz6OAIZRX+K1g6p/2cRiG8RrwLPPKdMD2Jain4ClIiuIx5yg1N8v6ap8TXC9zhs
sI5I1qVpFDD18Rblih8bpayL8eqR23JAEGeb2KkxqjKkWs43V9Ehwdby5NP3xWaF
N1ZhV2U+rHSrpv07ZlSHiQCjYmE25eXBlg9Q35Cql02akPdLXxzceHlPJ/K2DB4J
1Nh9+KVD4qyd7fY5abpgRwvgUDQ2DthcncGVpaJBZrUBZcmf1eA/jizpQzee3fkT
WqJpgmoCr8wCbgF/I4en4YgcjPXm1+g9rL3Q2aQJrx6VAO6X6Mw8zzbyYF59dVlq
BTtRLkIioYoC1UoQknhT/HM67uoTmo6lArvbpCWgHMAL3fUgj4cRgtidJHC52hkp
XNwNYloEkObiJ7qWfA3p9cUZYgnfHG07HGlL2Z1BX0/k/IYIxLxopMvcteAFYEGR
1Uh/a+uA5IDfHj0dCnab7h+tsaHH0VSFWVmzh6OCh9cmYFET+4yfwjEAA2c0pvgT
JluBIOM0hxeMtCZOn9uMsidus9NOD80hLNB5qxRG/mMtQLevOCQCqEgfKKqIIEU4
MH0rkhpdLyrPEK3CwlVLsZ3+XpIE+8GcIs703orrapa91acc4UrhiUu2WMnmpem5
Jetzn1fGaArUcop0hDMGMwrvO/tKH3QSWBbD5uTQdIpu6tlG7R8YZA6tB6M70hp9
JQpopOgksn4mP0u0SqljXWJnCcwlLOFr0mM71/MgOJmZzTNEmQS4mJuOUqhUx406
VvbW9yGbWeK8nqJaaLbc1dNCjQKcFrXP5i3sk3NqWmt895ZPHrTwqGXWdYFstZOu
6eUKXuqRUGviNmv3Pq5roSdfzgrexPYovCOPb366qU3FyuyV8SRoZFIXlGIoh9so
UwrYJDjiktkx9i2WH/EftF+A6cgoMZ5mNaoj+ywW2OLDvDXmArYjnQJ4ZCqBnTc4
EfKHQBjCR7oiL1IwRzr5aWUwIi2N/nOjf+O0Tnqr4jdH/WWPCG5winAjIKUwt9HA
efSVohB2kKmqa2vye4xmVoahgEaDERdWCTlQqXdKuB1d1N7Hthre886rCRE5izE/
mNXPIbdFG3vb0Pi7CwZZuNEqT2nkrjrG7qqEwC1SfY/E2Ssdyg2JSLJXqs3Z78Cj
4OCQgO+ngukCUMkPaDP8a2UqNevRt4IBOHZ+sUeQUfZf+joya8V6WjOEg2qyMupG
a4/SQ2zm+JoLj7cQb8TosI4hy3k6EF5fRf9/Vo8Lt0/4OYh7Q9xmLpjOVkzNJsSx
LBZnw/xlHQZvRYNUDVdVJGJ5isaT7lcdc3N08+s0PP34I+nV69a6YXaStbFgYn/s
mm5itn9DrRCSE7RUCYB/RX4NrsuHeieK6u5dafQ4yXFAViFXxAw9VsLXbXS/uMRe
PSwqE/QVgTTR1FTjBtNIC5wdZeGS+RY7rtWEpH4mlmxv6sjsUm9yPGeakqkKqAzj
iis+Werxl8ntzne+XfJ8FoR9/MX24srQQxbH9tnPYyIY6cBRIfUnjTTTyVxh3J2c
BY2N/W38vb0kqQbjwZinIQiaB/rmg1Y53Ih4hTS6QZsz18tAA/AYZVNQrrTd3FmH
PJIBkMgZY0IP+hV6qyGiuI/Lw/FINiBrSpiaO5+ZMEowTMYxecVkRxP4oxJNUf3S
0WdIutrHh9EXmFzrG3ICqZdFVXEZARsx94vsE4HTiv0segbnd9v5nEfbNAjC9KdE
DWGObgs8FshgybiB+y5AhCyWToDEdpe8gmhzwPydsCtXYEMirouB1bdgyxChG/97
Eyp1eP1RFZtkoVHCSKXFswMs6o0UOGwcdQtycKsXft7HN6NBmsNJF61dmlf2yxkN
UtxovN2DWv6ARYHVd7ovmwfiLF7xzdWZxJPHvyenD7Sb2T84gmXXKjlzku/3yuH7
/nVH7HG0VAzzdtIh9fCxHmG/utMUaH+0ZtpsPiUbRxNcjyMjaXDbmze0CsBe7AhG
lHBz9/iCBxBaTQg6MUnufsrjrZVLurl7dagtZDiUrTV5vZigYEkKJcgAOe8ThOUj
9CB6DhyVHXVtFq0cgcN7uW6BtxAgH5pr+WtcJuJ+hz3TbJvRdhlCXA6W4UoZhfh/
0HPcOuKmfBz/CJKNSdT0+MrAb4/AT/rd7oY1TIy+DUvf3JEGplxTEtjMz8U/KLcn
K45S81yXjn+RXZ5CVb/Z0dyLUihLdilRvF0bi1qWwwO9VsfoyjbiOZJ401KHk5IO
BPP52fvklDLRLlomZjSwIl/NNmldH+lbRfl5KYEwtHpPQvG5bm6aRCwwxfgEH+TS
sf4xf+sOF0Q/bGkd36Y18BKSqtzbjZgihDV4OUUZ+kASqWFuO+I1IzsUo0wuHv84
0td2d3UWbwtB1w9rDE/0Lg==
//pragma protect end_data_block
//pragma protect digest_block
enC6aOkBHaToSPs3Kz4ZB5493IM=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
XGDahoDVrCtxnnB1kX3iaTqL4Qb3DOM1g+3lDiMJjBCHP6SaNduVP14/LYtXwIdf
55XYflxQdAdvRw0YamudYqigLPILVc9fnUUZJuYrifHpW3TpRS739b1Hz74zUqeG
rsSNbmKKsNAUUjBwTUJQ5m+0V569Srcl27Q8QmvezHcifDGhmWxwZg==
//pragma protect end_key_block
//pragma protect digest_block
+3m+Y+A+TBr7flXlgiPeUY4h2WM=
//pragma protect end_digest_block
//pragma protect data_block
Kx33ehb8rEptJWtGJtNs4Av9g1sUvS6llZz5lpYoOF2wXVqqxlKvJJrytQfcXaQn
TNtn+nQWBKWSm+quETaUkL8CUL4JfvIESMua++mB6M3VMrmp94DyIOLfT+mj2ZZf
GwaIM1WMwHiho9F5IxDskVpHe9qlUNeS0fecQawt2Kh+mFdfiTidUAEGcdy6GVW0
0kF3JBq/FxvYGTerrq8CtosSKVyFmtqM5KZmgaBuk4IZXprjC8g9sL2RFJANqFk2
7rtYgxvEiboZdMvalHxBQp+47iBXTDu1nsU5JfWrtJ7RldfVLbzzB88OTLYe1VJK
AmR6v12KMtXBJ4WqYVWJrJlXN4gdbODP0hcRE/FDQoAzVCIrXjuRd1FsAKXZ8Wcn
hwoi+TKMtk7udH6b96Dq6g==
//pragma protect end_data_block
//pragma protect digest_block
a4pNMCRuTJPQrGwDkJYwF77g1qw=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
e8xYTuYuRuWEoDS3Qdk+pCoKKveVZ122GYXPuPSoFgkPg6IWjVmJ86qtZOiEFDrv
pUieRHepLquSrPY/4u0RJL2zbhjdAdyOL1FVlRrlen0wvRl7xDc+LpYGqN04ykm2
wwB5huljKCTrvsIcdOpuBHclZSk0FIWFeIAF6Gpix7nt6t+HXYAyTQ==
//pragma protect end_key_block
//pragma protect digest_block
+dI+Sqdpfo15FD/m6Ajjw8DY814=
//pragma protect end_digest_block
//pragma protect data_block
LvI5XDwEOJTVoX7Vm2R5uijAtSgAbbTB9cR+d0efz10Q3hstJSrgbaEmRDM679ar
hqEBq2ta1V3txG8B2kpCZz4VRXcRUcVx023hvaqe36CzdHr8hAnOkrdjc2tJXWh6
yyte21etr48aLvo3HmYIQLEHMdzkHjDYVQ7Z//VpDDxO4y7gqsgCDBu5sPRqGJtc
P8HsEX+SZFykhqn8sSPdy6ZavYtMXvS4wZAivg0cqhaX8aAar2ZRLxiOfupf9LCU
g1jc5DZknc9TwTOhD/huCT3y/9Vxo8mXOkOm6/+fVyn+IqTwh+W8yYHYjWWf5mcq
Jxy/O7i+jPfr0DMn4OIyvQuTfVb5cUU3bZTqILeawAD+P/ZguwdBvbBM09H+QgS2
4SihKMe2YaU6ujWVy3fO0iqhbzWlbuFAR2XoebM1izBplyy2ES297DCF1xOgSs5y
opRvSseXmCikFQIK1r0Hq/XiWlBHt8kp1Z4qgN4K6kVXLru93IhZFUw8TD8DqIW4
eZ6vUWxDLRdae56uy1FVoN87hDADogj+NFV+8Hub9BVfXaFhZEmqD1Y3yY0qkinU
UIHLdfJc7nbRKYtJbW+ZXqrGKvcAhVCoV3gD5lNxTpyjjmQxl01h+3Eo7DAt0Q1A
pe9C5yiD4rgZ76vbCxVSts0do/wvOwRViwzG0Rg+TrAodmw7Nz0Z2wIssYffTmtf
G4FbCtD7AhnVCRKRcB7UFQB7d4rqDGKv4YZRf8WUw9MDYKEU1C2xEJ4bt1bUcJuA
IE3AZkf6AzqhWy00peVuweRjNRjnvPlsagJJ4T2hiMqmJXe6dvj8/KZSUvESYslO
OGN+d0iMxUM3bh9XQbacDDsVGntZiBM0jpGrPxbKMO7rrSwL/dYELZvx7X5ebJ4p
Sfi9QAs2qUhpFhfzHHfgeG4AS0fqnK0o1zMZKiKZU5+2H3hTNC1WU9nCKudM3q0I
14Ojdob08AH9QBWbDH2hE4J5MT9hhlYC/W09cBFU0tIDXvAG94GnIHVTUzXtZeay
/rf7qQ0mVq6ZLeJPOb4kZG4nhhzcghDWttN1II71liWi0v44BGfHRU/QxO8RTqrf
M2qFWVSU1CrKPa9LWsFUc+xvyFu1faaZjAW3GJM7UvLZS/q2ijy26WEZ3ZHd7yCM
+nx/oqEBeYFJzMUcKM88dz6LnJpy8m32t2xLFXXVNGcoDTu9AqBALpCK8CTJVqOI
AfuGAW+LN910gq0AcNl9aZioT5UHbFTh4fWzsEWAaGLTBdksvAfrpfNd3sE9MMRX
wHaxt0yixnouDO+fDg8L0gNktlIjWauH/zwn/o5QgYwDrlpUpDAkwqFeB/GnZVJy
SGX0wzP5pghFpuYElhfHEWk2Tl8XkfHBtQUM1fzGHuVWY8a5p5OtKUhawc2Xxk3N
gT4c2Fa9GDaVibc9uNKrXRsA0027epEzkqM8y+F7pMsqy3PtEP6twkK9Qdn6YGTu
XZF2IJHRk/pJxMQ9DPoegK5Bqg4PzDjgZaT4/FVrzRkbVUAKrZ2xv1ZqQAChkEQd
1JX1ElKzahAXfpou+QtG3UXpmPCFhRW21Ro5TpnUb1zNiSwOkP9lJLOyGj5YWCF2
ncETfUfKQmaZBp39BlKxjyDiNHdCu9BRIMQ7Bu44Z4oQZ/CF+k816qH0UDF1d+7D
HPUtjeP39DjhZ6bq8VQDEOBCQsUQYrNvMtyHwsN9brNiRGgSDvSP53TU6kGLuWNh
YCxBlG9N2ziYHJjvS4fZTZZz/eFZ+V9Pc5dgFP1+1AATyN87i/4ujMUc48WbfZNq
DrMK+lOCx1fzzhN4bTE5msVe6mlaniCQwSiFNRLWrZePhujd3JMV3uDnAv5XPAXI
o7SoIiXVFeyP66Y3qcNnUmS40kCslXsB1PaGh7B0r7lddbXoqYaDsiNjdaLGusXM
0ljYJEAlN5XBZy3fVv3qE77VUDiqNdA8+8KEmE5nd4OPS4rVHSsPVR1fl5OEMstP
GKwzNCMfmJTotopbSyE+9mDDn7vfZu37v6atw9b8XiXv5wiRwkHL//Yu+2IOOshp
XX4kWc5wPahKohOwUNe6tNLr8vSv9VmFJR4DZBtsN15G5nUwyBiRk6DIx+dEnNav
ut5BfW7mMnp8JHLdqh/vjEQkFEvgZWsmwfOGGjTACjnQ4yHufV4S/B7S4Ox/svUA
FbtTEh45h8qEbrw2FgCniOZL1laqh3xvnfGHf+bx0e6Ql32ZMIbYRv8EG7yAq5xa
n70PO1rJNxZnU9WaM1r2/o1Z4yHuVqFZmPk8HBDxxKdIQaDU9ZeIJPnvUz9WFVqs
J5+okJCdyaoYSnGszXHjCN4PdE2uUHFFR9fAQp5h+PA0KvqFJnD0p/pmPuCsM7nq
D9kADMO4tsbRQrOGLfO+A/jhP16W4pD/JNNV3XEa3anM93q885+uZbf4OrSJnRXC
moyx40T4jiTI7k+Q+O4XXB9IAXaQGmipgVKWzJbcA5ogyr6KzsbQgxr8v8VguQcV
rRka2d/b4JA23uVbPzNDEdhsh/5TtM1q5WBtoTBWgH9Rh0udlfFaTf1o8dJUoMO1
xloOZoFivsYQYn1mSwtDxXfuRLg+qAWrQTzXIq/2bjVBWJ62SpR7Ua2W/GPbGiVt
zwnQMD+i8vy575VI123TkVoFQjkL9k6LQjWBFd2gFY1y9At1DE0ckVEhpvyFzWT8
MiMBcWMopMLhp4h8fgpIo+Be9aLM9ee0vljvIxjtHv2dC80fSw2cWId2avpALet2
3lWC8YChalBzaFiwabvqL2jKukZMcORIuQjJZTYwNnieVOU3DKI/QF1dLb4f/OZP
mnEkxUlH8nIg/Vt4awuOV6CBEsTbBK5cRVvEQTvfZrHIxXtBUZwzV5jOTu/mfHFu
vKnWJtdwpio/vj101M0mbuFqGwmZk++psmw9j/yZT6KolIlN4pvQjKd2cHnf5DYU
BNOnW5TS473+naYpsMUH09PhArDgBSyFDInYuiB9CRYyX+4yVI+3spUyqdsXu6T+
lg+l4FGuhNqkjWuyAzV61REFcjd1eujugPki2FsW4t2F7WLNkQb7jLokKE/OiQeV
/n1BZlncgHDvqLPx7pDraq7IQnH9G4P3+oDlyuPiuq6zbsZabNk3bnIrvDSVD33H
u75mO+8ScrSer4qfKZIcPZLPsPrCH0tHnvvuuEauRA5UhWcf8oRHait0QTINq/jS
8XG/mJXNHA2Z0Ov0p8ALYiiZ0gdlJYuPkCeV3lLiJyQGfndr79IS5Bd81clUR+A3
V3zFsznBP7cyRbRPlYQHspfvkYv0CTFpj6qPTh6/yhTBVbR6bPK0Yb06wGA3AKKQ
S/4iBKbEmkMXxddoKtwhGovUUIGiDDgK4BogpZqDlplcBuH+//GDQz0tsjoLJ2IE
r4vFJrTm4e6dR98NiQviZpF+Yj0ojZ1WyDu4H8+lwdkMSyok3JX+19x0CdF0EMDD
Llhpja3QSKph5vXW+snqWVVWHmSgVm8ZjJ2cs7FJD+xsNyEqn/cvCCJ26vHbf4S0
DZP6lrzsBE/ELCPtQ09d0nqaul+v4dn81atu1MHSU0MnJ4NCpo37D58T0edvMgm4
HEDonuCY4TJOI5NitwPo5dmvVQhKHjDZUs0RJ1o1oZPY6yYhRCGVlg5L33Qpp2qs
A528R95GimhatelMaAdpWRq8tPOpxwKjIhgcTGehJnEutB59JRlK5wkBiDlSz2dB
e26QpzDt0D2dqzBN/kq2sQD54GOI215WuE7/eU3qyY/wrrQttBWC5bNLtyYNR/vA
TQx9j5B+SlDxUc9MRxBWHUZfKp1mJjacSF/hOlzil8euX/C3P94IX18QhgjEHcP7
/L/JtUSdruXqE16zEiz0LpfldnZVl6FJVrVDCfHRfTeUtbpmzExEFKIEKO1q4Dz/
SBSK1dTj0uiMSnICX843olHrZL3SeqHbSjVMLQSvcfW8Om0iiuwOfLCU6PBuS3l/
yAej9Dkgxx2AQnWgslVxen6XdxxMQCpNqmmEpcpM1iq8zFR2apRscrPp5LYmDRFa
bM2+ExvkRFF/Jwg5TeJfoh9XwgUhEskqWoacb/EQ7um0GnGsIpM7uyXhfidTbHgk
zN6H02rJZiCaTIqEi98xVW1t4+5IfZP8eUumzu1LZrt9CL7zzp2NBlDGjoVwTRpn
cCqSSG92RUiiMk9U/0bh+BmIbZrQ6iNdNlwaqZPQwL6SLvdLAiXgaIjp5gcia5sh
fDpWwvmjkeKAKHfVaCQZkZZLDZESj3646b8hYWn3Ae5Fyqnm8+FegbdUOtP2b/+h
hPJ0QXj7vjVkYcMmKORW1itCwlbf6Yz/c1U4IcIer4O6IvdOq845awxIoLLtzh4r
6KwLwIve+n5h86qDwMvP3lvyeQe7AwQdSspMHRQVn9a0oNgXMczskX95qbzpGdjX
DEY0+RINVacxZKCH+EIW/vZCMtGKk2BQX4MPqoCmKQlRfZwXXLff9rDikVI1P6aP
0lPTGhrn/MZMMEzr85Ub/OEhHgIO7ZNk4u9Y2IlSkbEh1tE3yiBKVCUGcl0C3Sfh
P5F6JW0C9gZnA2BjEK2lHj0qESgSrI7CEpuxPGbPNyiuh3uTRDgiXoD9Kw6xVDtO
emkfhIFpTivxPr9h3oBznV3MWIX7BO/IQ9sDIFXkTKPfn06kuxoNqKt65UFbrf7w
QFaw3PwmGiHD87ukjWmuxuzq/H43kO/mVzVI6AvWSHaHRSclx7wyTyBCFyfatpPq
4lcuadENUsGxnszNs63QpZDiWFtoJT5M32OUX2mFZkww+JSsNm5Nl+yRfyONC1X6
0W8J9LY66zjYasV1O2XWf+w9dhoSwLfG+54HBCUDzr54Vb8i5EeMLbmguKd+ALEL
7yfgJlIcgTTBntnt7yD62CppVPpCR+Oj9y3BVMfGZM7BJgtrF9NYFLEvAD0dQ1y+
ycEibV+SCconafOAx3mPilIqwwyKW7w4Cnn+4aAYj4O21xLgIuARk5CvkBmQxidI
YE6I/5oSm+X0aQSGthiq1+MLRl5lUdkhPZQGRy4hOeLaI/ysBCoCX7fVSAHJGiJB
volzLFGVJLp0L3briU6dFbuNlIVi5QTnDHnrbGMQihqT6EDoERHfJjd3bau+yiRi
HVCSaEcekIDPh67mU+9qX55eKHp3Bgt7E3mol7GUPJQ/Hs5vmyr4EMPH5C0srcqH
6ZxbbgI7EZZLGz5Wq5CEBjQGaueDSi8yoOuwsUI8j3/MkEVqhYRXDR0T59CntRPq
IhYF8Zl5zBDf5HfsgiNRnnCGb50jrhsM3hXvWSiwOj9Ds83fmwjQc0zZBBuhQwHz
X6DtuyOAkoFBpinOm069ryloaUdn7VQvSE9ONFeZIl3g7iT1pXIHUAys//e2nc/G
648UeskwXQQAgqjpdfnFLYlFalNrIvRU4kBKwBgFmrYpXWBrG+g2qy0cKNjOBBot
O2L0NajaslwLOV6Ee1jZrgBrJDg+HQSVSETZerQrcA2EY3sf853IG6SvDQPiAJHg
Xzo8vHAXYGCRdi1jn+YY/m5lGVJveugov3b2CPmO/tzAMIfF3sfjZIKk1oA5peyT
gKU0b5T2NQaLgIHZLbWZYK44TIe1IVG5nDa5CiPycnjVf+KtV9BWGxTCT0vHqnAj
YFONrGUPX4Tc6IrD2hJiFlLrj9rQVzZzgxCifA/YAT4Nt8v9GCkqKzXtjmHhgvq6
7YOGULxnaOUMd93kOT4A4es98mipyYQC5t2EDp14WJhRuCpl6ZjJQWiv2mrM6jcV
RYg6X9BnDKzVOVIo4BSUSK9aEKetzKB8dOhNAjazHpvYsOmkC2bUzBSMEoZ8+FIG
awZAJC1sUwtlp/cLootmX2d8coPI/sQQPQo6pMPrx86sWX2+7HQNoCpLQjdr685f
S0R3fZ77jFQatIJAx4ajRshsghioRCFX96UmK4I5f3qEV6ErSCVleGh0Y+bp9TGd
dzHLaYZ9xRZveJ1adwhisE/iHWrX1mgLNFjzexP/9NgfFjaS2BUBGjoB95avUmuE
UkuBem74xXM7V3A3N7C78xhsZbftNOMUfLys6Fb8nTkJezrw0E35S7LWUN2T73XB
z2ElPC5BaixajFJN5uy4EaPHEaXESvIhU04zA/asOD2KeFTSCt7St1xyOXDmUWRE
BxH4cjApmdmYOr5fhj1hnXHvYPfmuEo2fYq7/yJQIhtCubz8fQGGtnjYsvL3WGC7
82tDlmB6zgUcXK1A9kPlJR8kk6ZjaKh+FjqgJ+dXWf5PGv059omzsrJOw5BhhyIj
tdgyDPSNYu8m+5syYnaYMp5jXg4I/V7DxrxCeetHXELrmmLHdLYt0vbV0UtReeRT
HdOxARHwsLctRrH1vcH4GIs8u/9wu48ESftRhZOei8xAA9gI52KXhnU4M0Zu5A4I
qOo6lIdvi9XW6MKWjpoStzgG4z0BrAl2XHPZvXcIEbw0OfXtfXpOzjb83/WDGNLm
3k8NxPKCi0xOPDAKVal/BMBMZfc5KZR9xDRIM07Qh8usQupfoFshsK7b7Gl3PpUM
hSW+JXfQdIb06Xlg2eYhP38AOebO9646yUXsUCEQktqWOANulkvqH3zd6l0FN/20
hqRvY8sRrI+vL3RVrYxdqSr162Ld9rfMlUffPO040XhVUFWukfo/qOank4GZyt4m
EwGfnIZl9pduR7AD4VXmEPrKHSTL+5EDBFTZM+mh8aBVLmtoKaXb+FtoXYE6Vd/j
HK0KEo+ybBRqQx5nSBr8S99WmFdlcJ1XJPnkkGAjY/RWinHWkrOLutK2SkNZYUMw
etSmkkpkdLtJGh7a2VmIKtlMWCaUZrj//VEU4/aMiWVHlY/LX6mpWGk0WU3VQVfB
pHli+keZhxrQU2qNWFNey8kpGW3MSr1Rhz+uHnvtGa/FffJsJqRcx8pwgZjSm5RJ
VcYeHC8aV4dn2UpkM7MWShnoFiCIcy6EqOrDuWZvQqHffH7aHi8niDKVOQPivOys
oAYFxDUV8Y3h0wPwh6cuSuNg+BtlwqCkTkDIq0oLqb6Z+g/04vyC9UAUFdTwMD0C
bjPXcapUAC52lecaIii8m7vLN0NXls8ITlITE5+WtBuGOljvg7FPm/NoTcdAcEj4
R/pLYMgqJYKE4RK6I5L0ZUKfHICDpCTIa99UuQAfmCx97YVk85LuflIMYgAf8ivC
lOu0+UtC3sTLiyA9XdFAaHrrx8Nl8jOAmIWAog/vvFxLJtB8ETvrSJC98xzFqUNW
zkilCzVE7wYNzo5zrzGYS80L/hT93aBgiZ2MD0azh3qbFOjlpkFPwz5KOaC+oC1U
ZCLEmuBeOwAxaSCVI5xPJNQCcI/Gjbw1xnUdzIpJIISz+wqkJVo7Zln1rVNXk6GY
ofO31ybTmylCLNTnhTjffQ0R9wa7wUGtgLLxrIZnC745Au9hHKLSAPT87QziLQGg
f1wIa2h3uExAuFd4CtgZwOdIBziebuY2c7WL8d9SGi/zep6jinV8zcUecqbqBSdW
7KXS/Cy4lHKvKeGvoIpmgdLE8QuwkcJVhNqKFh4c2Dm21x6LkRWBlx0eWd4spjC9
VuI6mM7R4cLQzmntoCXGkvDMOtu82m57/ESvySOirfQL1QN57HSoxL8x/Wk1N/be
AE+eZFSR2MUdoEt2O+WBinnapT1QrhXo9jMW3Gly8qaWh5IqShPWve1D6kSg0SAl
pFWNji3vXDaw496sRWkUkEwSJfxMkod/MHMzQ2phCjDI+R2oHpI0o6tYbitdY+CS
9wa9Do46r6K/5xi5lXtJMYck3crPuxwOJgNKcCDkDIDjFkaRvYHJMR5fyYkzhEFi
1M/RhzYP7hyKPh4DGCI4Lx47HoOFSp04D+XiwxK8U8T/57wcXQzDbnryXnW6oJn+
gItUtLf/uMHnd3Enr9NuA8KiwwgoZ8DR1aaMP+v5877/w9tzZ+lkZyBa/lOF7ym8
lienOYOPFMQ2u4G+xbhSWClIJ5SucrvsVqBGMJUkVNGTCPa+b5cmJaBSRBKXXoIi
O6lBOS3GI/Rm98ot7SlFWo9KXRqLsoc24Afz6ulBDhY5O8hqFNB9NksxNP8mqS/V
UWOyX3uAn1Aq5kuOdUDCpJf6N+Z6nElLHH7RKBRb5Og82AUU8W5/a5wud1h75x2b
2xkHQZpc9DynfJwbygrt+XizF8wfSwWmvhwEnDBOnJBqApC9rbGZ8YtndXXbVAIr
6e9G4zFM/raZdNPjuQwQhcHW2LjXPJSe+RRggU6dUaVEqnd0aHC4l7xbgJStIKZJ
1uRyzX4iuvud8medD8HIA0iE8vD2jG3kOEaZKXAiEVxnyS4kh4VV6NGrC756U9cn
W4qlauOFfeSnEKvI/+t2Pc8Lls8cVG5mw9nGXjGWLntLwEGUPTNRZmCrbdPeWLDC
K2m5TosAK+T5Qe/t+mQ2UlWB7+I2pI0RaNd4Zb/z25IBjIsXEvGMkgqrkF8D/omC
juH7tkAFShuMAzTHH6fVSfrWMkOfvgnPqpRsMpF2UHIk5ubVL3TSM7ai2FoT7Eea
gOFkm8ASr/JesqzJuAIbAJE08Qfy6WutUnQoSMl1O4+2ITRsYoxIsjTafVS0krMa
W3Lkk8waGFi2cm3Kc6WpujjuOrXZetG2ELJy+pTHwnS+eJojIW9L2BOEyIEXLS9r
nBvTbnlXA6JK7x6Dd4/09OLg6z5g19hO6wFzXUFoT3rPcync9Hr9C7A5nYBhIwpz
VF2CYx6Z7J6JP87CHye2jPaRP66xUrH4SDMbYhhl+10ePe5p64dQ3/uYJ96+Jp4n
PLC6VtkIC79xcfQlH2ZX2QAJW6MTDxcuzuYQgt9+ZyRSlD3jzw2/ONYWNXnjzNMX
OFBkZGPs3g+AL1A7e6o8/hzxOM/GyBCkmO36Ry1XTQhR11vQU8ZgavbPVQFqy0Bh
TN/qU5xUTJTUhVk3WW8V8h6Z2tJtiPU7yQrvns5yHHXgeK3v/4dw5S7qALxbjMey
eTHpshmHMgJUu+MgJeVoeI2rOdt8qOhxMWuiGGhmO0dTzX1d46+UVvwz9BWia97U
gYmo9uC5uSYj713YLOQEp/UjBSxR610yj/YXO90WMrSgMHap7J95J14vTWbJJxCd
oUD2/MV8PlRB3iyN4pHn8sy4X+bC+jZeeaC9+XNQrmRKBbdxIwiuM4wn4WWSuGBM
fJUszSHbmBbMa9UdggWRb1cCx5iIUs6jv3TOcG/f7MW2gRcu4FnLE56ZXN6VIQ4p
f6KP6/Cma9dpwogvBi058KZaaTeN5YySiQBW37jjy38IcDTJxx+Ppp259A3QSj2p
PHbEOODjE4Nrvz6FEcy0adqDVKY189I0fK8HmKVlSB7fHzvwT7rpgTbSa4uHxstd
4/726wbSg0gt7gOem5DWuvRnkV1Mf6ulnhvkYu4fOmWVVMZ4urVmlsx6PyrSfnRv
6x8PufKyOMpkb9LjljG4hoNbeN+td614mf7Uj9zkMwLXSJ8Yykqg2mjQn+9JU9pE
xKt0ZgASs6iU2Q3XARKu5RdAZ43Z9R7OXVAO+bcQM5kGjoGXrKAruFOCiomv0rOi
Qxpqtp8q+RcW8QPRRGYlq0CC3UIUwzeb7AJD/sfrxiX7pE70E2jZY8M+oLq76dhM
umbzZI+T4nYH56tnlZt49fHnEGfu1lXdo9h7EbNDslOdT1W1DvnLr3ijKH7VTSav
j0SZ3CEVZ3FLNc9JouCAedgDGYQcE5NVkSD0LhOHJSufU4AhrWpCbvibHowQdpvV
gqA50SCFXuXwxk7Qq5bg2mulgM3wjeBzQoYHBdCRRu/K8lbGk6kYMqalqEJtJlJN
XvAHX55tPAK3tsJrT5t6Adg6Uo6LWx301jSgXLtDIt1RGXdk2mxdgfXycfgn/13c
9V6n6mI1WcciGn64DyXZbOkpnX4GvDMM75sENJR/LTl+Js2URejvZL86xGHOa7EL
bfkYA25aS5lwWpEh9e0VGC17Sxs9Qrz0CbN8n7cQJl1yf8a77bCcGcQaFTFFf3A0
uGIVWiyKV/1cfQ8/TcQGL044YKygLsBjjvOSbYo3VBDbdl/qK9yLroJTes/Y4eqH
ZfI8Lk05srWxp/qpYiOQgBrZMFH3mm3LiM2CkN38b1mr7TO8/8YjZqppFmXSvF8w
5DL1gNU4oCxGcFgAQHPE9+bvJCrnNhwK0+l9XP1XHHVtk7YvzrSZqsBJJiuFpboZ
ddQMFEXHBt5edes8D1ThJMKo3a0ufmjsx/ttuS6xeOBY/c3v/YVveTs9s0g4uIXl
X7YdWNTL4f4CX9d7xel8Lewoagu/FxV2WDDlh8SLmvOsUY7WviW3OjQgqvrShDUQ
g6UyEzx1a0ssyMqfF/LMqPJt3BHCkhBEGxGjfaolIyLbkeswO5CtiEQ64odZY3Up
74X7iMVaYrF93yazMhia0FGRyyWMI16j5+qG0TLpApEDN4bgU+7pU2jNK9gmMKO/
3W3i6g+sl9azas5oQENEOSF/mrWg6Jo2JnbbTg0FzAWG2LLSn6h/v83Xo2cHdMoW
zkkiP1eYUCog251uH+v3ogbw+0Me02K0QYlhA/9PxWaA1/HufazqQu3yt1nFpSFb
mg7KlkUBBUUMhZikhF1S8V1fn9RB17Zxt3pCQayOd5mirKITWlrDAyZeHyzkuFIu
JyJyU3r8puacfQgcT/Y77JMA6XViDs7gpCUDBV+oje+sDcNYkc+16N0Ac9KzQoQE
qztJdiarkpfU7cFpQjoJ1rFzLTBmBfehTkRQY6oabal8HzrDKsFyc5w3kixtoX0u
U/XDuZo5QiN5FNKj8v9DsW+C2ANPOVDz4eA06Q0GN8GrjF/ZAFavHZrl95Sk0X+x
jR+NyT8o9KmCiZ+2lnRYMMQj47ZSV9NOJERtD1S6zalM5yIKx50If/INmgONC+6u
lQpHhBCZELH4jR58dx0r+81rIqncbNxq/U6f8uHp1xHGegBjxz7ekf2iuW0R387D
u0f1luML1NTPHEDKcrxgqEYV6Legp6lMAAjHRnXomlODkQNG4S6CDDQFM781kq27
jPSY0dwZ8sJEWckFQK1k2KHsNxjOiV2AW3YAsQPkPSpCtShqgh0sjUF5fx6ZvNwe
+OROUtHzqLeBU+AQrrbIihFGmrD6RrOzaIDFpo9SnPpYIElOtzvOmF9tBPlKxnvb
1oxAiBndPsPbWQCxSpzV4rR8MNihaXs10Z3DCQuDhfwZ5WgvhDWCXzwKLkQWoYQt
nwaVIF449UEIUqKqKOJNVwBaHSNErfO/FY4SOdxB0PKw+QrDyXAduWlG8/TM411B
bw/icoISY/z2i2BCeKhjh0lROhitfJR7/A8s7JlfX9/cyGA7eASjFsPeVL8ZqCqX
f9Itc1eWkzL3EYaMT5LA9iFMnz/OopxUMzI6Z36RpB//QKleEh9bvdAY63HPs747
9onwhFwfIpGJ1GUxmwJKyeF5tjNmlmJdNAGxuYScRGROZ6g7EHXo0iuuzVKlfq2Z
04e1AN/ZPPmxFlkSj7XJMypSTAN8eogK47H0hL253Q76lIVrsDr5/w4bLJCAkOZ0
jxnYh20/u5N7o7hWKY8X0uYEaDsuZEBs7ctcKkR5xbIVfNuS8Nx7FOb+I7VcLWRV
mJAmTPRQ/hKchNVA0F62N7fbizf5XEMQJrNMI2GNt1x/YxkyjYQxTAfe64B7Hp5B
WV//oeCdR1NiZwh0UTpxv+MP6rUL9ulXdY7huEK8E2flz/mThlp+Uk2Vf6XO8kZQ
zG0SZDQFluHFHf/kdAjYKO88Ej60G5RzTG/6GQpnHPqYjcfgAjnE2IaZTC03jBZM
mtLMXHFk/t+tuslFQ2+9yPS/WnbK+SUBopYXlnh2cEPnYG5dxIcG6PMmhl6rtKud
4QpUbLLcW/SpEMeTDScOOWXLn04IPfY5uSkxck9j/OvUV6MbYJfrdg8/VvbNSGwo
3FyVx0bKgq2Lz3DPfbNsz8R9BpN3R0ghIo/NY3jQLb5+1NFieotUpyi9x2tw5hY+
yoz4JI6tKzGKIL/8IpZL4uWx8RdMsIsgWlDga4TyV/ZL8L/w+WJ8P7V4eiKJsvIh
hd4mxQCicAb6sciK/jTRnVOSaiqUVGZNq14uCSG2QFhTXEjLldC7frqU2MOARig9
AvnIVuGRtaKqRB46nNpI6URGyBGDJ90JQlBUzJrUWo00ap0C5zpPnKVC/DS37xs0
AnfGiDNTI8ff2M0hsy8Y0oGnpDBbquQZV0+/xMuCWB3j9DCgmiCAGFmdSqHLHxXg
x1I1rCQGu8AK3a8HhfAU8MvtCSgTrmHe7DTQTw5D85omhHbFrBdxDQSMQfyXIMm0
/w6ZhBDfN4XFEV+aYJfqhcWRcsahsc8WWKCJNHm+/6T5TSEBCenkxKz4jfs76SbV
fiQX1yx2jwioVvWI11KCyxGT9h4gt3iTD7g/fEVrPpYQR0tI4XmZfTRwmEcj8Nwr
3UI9GYF7AcANDQmGFlV/uwMeP88d8t06felQqUEe4O+9CxG0QxDJXpGg3skAYTNY
XhdEaRaUU0WMuLlk5ByNCEVRZ31RJVp1nmfXvfgxOVW4SOjvMcmQ9kwuUWCsL1VX
wOdfsMxqsxsgDrfFpk0vhh/QzNXZsStdK9n2ZctxUfp60hv/blYewPRtxiXwZvnv
P+rJy2XncCAPDyWDrvMs9y7cFZPJHy7covL4YAkX1ti9+dQ1zwU/c7KnhQiOXhfg
HSS68QB1oApLoTqcqlXddtcSVuWj2FIPln6FaXDSrm805iux7/FSXEpt8FhUJ0ix
dSIm8DkbYZNLBMbJjfGG5Nm/5MZB2Yk6u4AsRgKf8BPgcc4IbV1CwN7Iqrx8wKax
Hs9Xu190Dssxd0i2XX/AXjRmBx1plaXix6vqAM2ad9jCUcIy5nyg6gseYdnTkxI4
PUePXI8NmWcAZXxiLAbm9EYpO7KMikBLvcMu5udW63LBbHgSGxPVr8PLCre/qP3+
InHo1axqvbQ2RFz1YIeeEgVNdjIh1YtVZtYiUW3LlYIMwAJkI1MNwyI+emLzfiQd
8L6dKyUmJF1a3hv07EpK8TwBSgMMEg7XQdh3KiQSEnoIzLenbVyAwkOUA/MMR5ch
KHY72QuDSDYoCmMycSfDPp6P3xlhBtQm+EWIeQgMKTfsJ43bTBFuOTvHZgRNQfQL
v5fdzxqJxc0mvnNDvd3fmTQ/Df0Hu28/tOI4jJxw3/e01ugWe2WYoVTsEWAoUV7j
ytFQciMS5zNr1uExj3lXTwVouxMwk+XxSj5j8lu/YoaueWoUgTtWN9uNSgk4vKR8
ZQrohQ5SB4EpXEqxf+L6YzJDXa1GoaRrbEWbganCtm9oeoxHkWTCi9lMYZ9M29Wj
rMw5UwwY1aypIukQgT4IKKjc76mKTmT83Kv7morXP6zP5ti1FWZlQsZNw1e60eHr
wKS1RaTiYMTwktYw6UkP0UhkTifzkGULhI2jUKbqT9HfqUBN98KqhH+mfYBrsIIy
zoBG4RIcObRraS35VKIPlVtDMYCjdWY6rq1nsqxc4itV4i0EosS6YgURyYBgWS+I
0DrF62IyPHnSuIR8IIYqdJuR1gDHbMtg5lUbpK/w8m48ez6xJyKeDarvhrVF6744
uBII56OtmwpT5NGNRzElya0pJF+Kmpp4kCl7CVM+3QnfyFBwdHjI/uEv4+6TrwLx
61CO3MoQm93xW9+JxLQma8TD8EHNAtq+CJK9zLV6dno0TkTEW2ioq3MPq0dxdCzs
BpKwTDjelUrGGlESki4K5WW0Zpz/xYuCH1QuDLNvlj5BOMiCuviF4dL/g1HWp0Jx
qIOFBwKvsiqHuU8j1fpg2Kb6D8gAbLJMDF4vY/1FZ5f6q36xh1ZI9o3avHI3saPe
JSL/8Eo2jwbG0ekrkIhWELpGS/MNPmp6cy5vdKRkmWQbY6FfEK21c5Y9htWSM9IN
kMoO7XuMke3dlbi5g6z67jp7eD2Cs7WPu5vYPZAhR+KoJO5h7ZaTikbcYJFj4aQM
ZVdnSTcOU+cyPgw2osIlfZRU5iqiZeKJp6kSQksnyZz+6woZ8/Yi1IIqUSj77ylS
dw7hMBIcY9i1C2s1FLuE6AhKQqiM7mve2NE23F8yxXwDbMyejgpj4x9f/GNbKdgL
TPRZGDomAVKErsw5tYJOxVB2uCZN7dqR6Z6L4aiLigcpuRcrtG+xM5QZ5obFUmxw
w2WWnGkFP1CYgYc0AIFDrug/ud7jGAfPv2eeXtMiWTwW+L+iffQb4z7NF4M8yN3k
CYh/8xnHLpH89eTQoZjU43kw1j/zsxoYKWvpUhgqRpTA6gFrsb4350x1nC1qEL4r
qZr+NRNjzntSboBVcHVheHzrGulTsYxmk6jdi0M7k3OvjSs2USsHQlhSy5Qe30GE
thrkV7xcojgOteyzDaSuWKKzvt/1LXgfJrd33xgv25A4P2aXkPDDysAcRAosIAZA
CfThCf35uGmmYvZ/gXpkgIxX12EAgvvS3CjpuPeuEoL7/8B9oKvgM4ol9jxvh4gU
2AUMvKWNVyVm4LJeNHXOJmp/+SpzRBs8MWy5GLd7Z5P6IiF4Sb6NpxS+5GGIxOJ8
KIF6DUZ6DObQrY89RWIKbgFIt/7k5wdTpx+26nCUlsY4PAN6q5kI6RvDf3I6yTGB
GKz/fYNjk6UWJMufkkLuFRCd7zmh/NsdQ1FNoRAZTFatvGTaCRWhxE/gMn7B2CrL
Szbw0rDoWJ8C7J4chlYJaZE4zo13slCEthI5DC6gNdpvmWbGpDGzez10aPJp57t5
pt3kE1Z7s/JgkUPVm3uQqZT8pEeu/ZpPcQG9W648b/EQxvT3xy12fe+hBcinckp4
mBgwwXsl8uflRFUP+VI+PUS7mgXzZQszlN/X7XG7G++k9KrP5msGEqkNKI/uoYXE
fdySC74WubsGmwqyguvHoTwaHfBO9LYGdZv2jf0dkfPv8iSecy8VHqybozGtfE9+
zbD3ckvXBiXuNkMDEGuYj/OUFP8Gz4sDYMt0T0Qwkmt/+9HSF8d/OYA9QouqfRsE
WOXV8zGPBX1UA6aqevBxZFkfd/n4YsqUXqymG//8YMduXG/zqwXWWD4QJOMDrh/d
OwlMYAqIIOCUJ2A1/EswWWNozPHVYK097qqwG6sSDYzp5PNAipp23zyx1MaS4HtY
GE9jvt62/ExE5o4ZPnG4VXI1MzE1HKj4+YjF2VaXz+PKV4yKz4CTXO87UooSnptA
6lh+ItSM6ru8x2b9Uz1va1u9utaqjJKkHgMT7xM+lxmO6hyqxwpCS1Lk/7Roorhl
7KVNEA/XM//lsruU/gAoc0CrC8sxsuiWNHn12oj/cwx4giQrqqmdkUcNKGi8rdDx
ZQ17TBhwfBOOpxY8DgDxCD0Ow3pvt6fzOY6ms5T+9OiIgbf1clvQ5sYJ/jcrDvFS
VxTb9BF/2PRgFTNGOb++J3uWCO42FMeJ4cw7Ghfl3ra0J6xHEVXTH86Hv0ayRkdu
47T+jp7MuOTvvlERTYDgvJ9JOOSZVADVVtyOvecMgOnbhTTKF7xAqhL0Wdz0Pva1
p0EnJ8FTaD5qRS8Xuz36I0e6PXIWzCr2e09Ttxj+FmqXvKEZntJbFlOarXjWfWlk
5AK7wRTm9qm8hEZ4E+yNn9Z9Gi8/R3ymPwXkfVzR2kty1tV/RNlhsMUwVCWmD0/2
jSZmbW1wjpvYl+hkiodxPPlBYX2WTayHutgcSK2eTts2Z1v7d61KQrYTwc5YZYo6
pVPP7otfMceAq3Uxy3fHx+isu/yF8T1OWzSEKNugoohrjy8MBjcUBFWiT1EZ2F1d
ddmni0JGR+SLMi/+R5Usy1s31Z4NZMlDZ35aUs6P2IOitlyKkK5K6a/WQWiRq1ks
QYpLn8nUpO/8NOroN8RxFFaG4tjf/gwVkz4Fk+zrGnveVRrDOH5VpyCsmMyoyJa0
KwrT6Qby5FHzqcjw8j+x88T5oadu3bTN5m/oTfPcNWU3nQeT61N3BHADbqbutnQT
/JfIZ2wQF0EMPpBvaI5Dc9NluZu/9rpZOIrn/BYUyPy0G6lKpO7M931i6h1PP2z8
LoS3kCI+tntTrIrHOs65ztw9L70L6oXOdk6lFDiNEZdFo+UsLQpSwzmFglrQljDE
9ThMmR3FA30RnlM7O6SKlFgYc+ATYe0q7pZROXbcyJSWqe14/lWqfgD3NXKyMnQy
RCFNwja8FY3Id7qrIZtTIR34bJJ+57wy2j4klA7Solcv+4qYHdKzCHFyaolGAXHi
vxDn/6EXbjOynqO3h0h8PKugu5+3ZgTH5P6jE3swhYnVPsEab1vx1EaEbZx9P0nU
4Ll7Hkp2hFIV2IuAoLJcu62DL4flMY+EAOs67ne7RSiX21RaKbGxiRYzl5A72RWb
NObEMyb8vHfwdFUF/l220qyNqdobHT5OGE3OugrIpbvIqLGskPCqMyAnWUZYXF1/
ju5IZag0afD6TNUL4Pt6IyuL1/Beg+zPYKxkC3wwnQ1tri/yDAeEvTFzojoirnj3
XFxJJ5yYQvL/4N/GFOmC32nihUZkv9a23s/+Y7ow0oqSJVwSQ5ldnYq0bjqk5Kz5
PoWIEb6cB6iUXd1e7v7zqcVHfsrEVUiz+wt7sX3PyXRTVys2n7Acw46bCCJZqYoK
ALO/uzZmmINxZmia6r+lLkSRI9RFcN9QqcmH7LxdcPsEHV7UmsQDHv1M8/FC7lFy
86lHuuLOxqicuQnPN/F3Ft5bIDrmugQvJ1jA7ggy+zIl2N9Rzhdy3+RjKhkIom1q
/iV84mznnDfS399HJoXmi1JWRDLnkxPKT5kqdrWTfondb7I8Q2e+w/DCuDPAv2yl
IF8MN3ciAnh3hWfnc1d4EvD9pOm0T3hH8qXtF4rDBt4LYKYG8QNHdQlHQ+Q888HL
DVFqBUuM8ohheLQK/PWxe4absnNFpKRrrLkFpIJlJGgy0ALlLfCAcVrOwe/lN/4H
xZxek+JiugFLugQMR7G/W8zTOexq0wuUUB3GvItQqNtd6rdEPUErxFtnr+ifz0yC
pntdf9S8q8ezrsr/T8oN8NoM480TBdgvbWbRRxjXY+JbIwOk7i70TfLlNlgoVIxB
hIPqIWeyPqCYY87XlCGOrKswg+DzgMN1HQw4V7ptbOCDyHGLlCwDhTg3aVTf0GCe
LAEXC5BAFYtA75v9/0Jll4lZyKbJDSFX/O0QS8e8ZdYSMrKdYf12lOpqzPlqMwxU
HWfX9GMYfFW+o/Kb+pHP7jpBmiaRUvFdu4OZ4s4lD4psmHX/GDWbU3KYIAHo2Y+d
bc75Uy+1fRfVys9JzBvRlmc6WjF3dNOpZIqqBNTu7JosqMzaZ+vyWKbcyvcXhR1q
uMzYnntpULzzJ3yTktoasShS6P1sDlIxefrdbVk2dNNP9hv7CfpN5W0cYguaz3PJ
KtHURRtgw5gshj1CUUy350Y+AvpPkYmWEpoknt68YumXKmTI7AmeAgTVJb4Kj4vR
Q6eyiph4ZXXbKr+WsmsfRMNwGI+XflUdP5INMXEabR0ycLlHrPNHcDmYrz5466cW
LKwavantrXYQQ5Ju91X3Hew4Cgimkbb+bVgoB6VdFX5PoPwYvOZzuC+A5mj70nWS
31ynuvihsFg/8YagWKPpN6ewRNH/o47JgsSADcRrxGruOD46xxC0jBR3gEjdZOJy
mnQ8Ob5YQY+cSc3/8U6SwyDb+MimwfMG6a/Joc9pAj+10FZrlf6PFQxja1W/Idub
wcJFrH6DGLtvzgscSBz4IR19cJsmPrUD5GrRESV5vGK4yFMdSQrYIxgir2yNBjSc
emrGE+enadl1tBHVyond490HEeK+SsEukKrt3R99kJMZMXGzfp49XJ+aE45qoplY
dqk8be+KPz52Mq77LUh+Bh3dO0VeLJkk5zAEcyF0atTQf/dVXG+98eBlx9Vc6m69
AT4QBj0a2CTz7nBVRtbzh7mQTjizqRPxLMbremf7vCrDtnQWFGKbmBfCGMI8IJc/
iruzT1uEaIfLT4i+agWUv7j3HPg/QLZmVEc+8//6Gd6i8vmrHzSrjdgwI8BJHZCz
U8Jad2w2729a0eJkxPnHUzuGT8+UNW/CZejvcAjz1iBNUByoFdr92GhtkEgIP4ne
ri1khGDyXQ1nUZxQELf1QjgG1lrrqpGEf+/KpNQy8b3uWHdN69aBwda7ouztBjcp
OX0V2Ofyc8ayG5Mr8aFwc3kfajCDhu5SLxkOkc4cXxeakGbNcmzkPa34Lk6VrjSS
in9jSOLLLb0IKqAi3hh44wsP0JgJ824cm0VevXoKJVsPFowDDgIZjMDy3JquCGQB
XKnHH/KVcNR0INGLmc+AYm0oA0iq/UWImdEVET8o2P0MIuIguh2UHR0te3UN+6qN
WqRk5RSvfrC2UI9BKx+Lk7oZTFCbm6NDmtKiAHI5eT7XqfrTGdRtz0XkVYAD65/u
BWuI1Cm+GhRuY9RQ8DwmNzK/2znOWHsddIE4I2xEMa3JWqZixisDLofq5fVsdXSA
V3QKrND2HLK0D6kBYC2IrrmPiTpAT1cZ0bg1nUCN/wwEyryUw3f8PTutOppgHggp
eqduYjIpw8RAM74pO2NbB/TRf2TjjoV4Lfkb6emUCozCumw9AkXAGJSqTjIzJo7e
TZrwNrio/1DNbv80R93hdyd7M8S72ukK9VK07CSmyrTxiJ2EiWbozAobRsRDN1SZ
sX0qQh4utmSSpFd3EbCArFkaVCXdAGNaQGF1EacfM9NvMw+584qLoaiW9nDWBleg
x+hTqJ6ZC01EAw/KNKFLiY7Q+BhLqe4YEbrf5EpvwhsxNOlKrfLaGWC0/l6oxnup
ujhsSTVU1xUl/NlgmU4VbQucsr/S4jSeiscFn/A2wHi3o2lBA1G4fSGhvMI7xKex
1pN8ZNlS6lt31291F/Qhw0ZH0TGiJCdOUUIF/KyoIDyvwVGqIHo6l5mkFvkTaFh8
Z3DC1Ix4WVBJvNcQk2fNDqdtuz7nlbit51D5e1yrg2hp7HgaYiI0PwX2phNCPEK1
szol1WH7shR4DDvhRUl2WaqVx6ebS/Fqd1upHwMTKhwXwaewtsnxIuCH57f8Zpox
n3jsiibx6UNWwLEkEN5DN2X8jpKLhdkkcpma9QiWZIqaqyeBDPfNSUFVW08LFdZ8
3upHcP6GR+ZlhprDpod79EYFMxyQ2KBKBTuxQQrNmVj1D9hUSggIIsPP8j5ZOaoO
1IJwhcKEWAK3bZ86qBu7Oyw/Y9nLEJBbLFGP2YUjjytjDdASiNJIbSFtBnmJ5sb1
C/QENE/ftWAT2IzXfLSLHLuRjTbrvQ2uSXY5F2TdPgMlQBvsdPiBZ+Hf+UwxNutQ
w78dv3JVv5kyBFJ6OkrwKzw0DRG5PVjODF+LrD1QyOLH/t4VW/9CzF0mnF/MbNZ1
ETsw2Cw7ju1hIlH0jgPFf5fBjSNYO5++xNxhMbJYSMaMcmdDl7UXIFR12V2KTY8x
GZpheij7XL0IEPOlFhDwbxKNYsAwhDuYWXaT0vZMSpY7LdTtTKQ+Mrroo5rMx7P7
Q2Or1Qv1pBewWWMijQSMXcRIAYm18aaG39s7b9+Q2nLoZEHxFYtqTRcBVk9yYav0
xImX6cpnwAxbanvEMTcX82FuD3tHb0WqljO7ApNrl9UzeZUrhv7Uh8BRhino9nfj
9WBpALTz1n7S/AMA1MRjaUlMVnX1Fq3RY/Gjuqrjv54x0Hemn4Ne3ma8zGzibPo6
djiv+irAdvJ4yNsHf2ZIXb43YH9wwm2bWxRZcACXO8Cx4Yvq2oNPnxcVNXmIIMVV
IrGCXXFr3ZqMmRe1xBBAoXC/2cL4wxqFX+OwvJxwtV7aXmoh6rY+e/nd2Pyb3PzT
T66ccAtR/EGr/GIADsIVGK+hEybiyhQLkmk+QclmjsWXEl7aqFyEMUROUVLPOF7T
w6azlZdy64H0bK8qvExC6kyKE4oC1lQyExGPxgCOGeF5o/x/bw+dgkdIndXScFOK
eMD7FsnJgyL/du3UNTmKnsYNUjM6DGfV8GZsLR2pWc4Z7gitx2g3fYY3MY85N2Kv
RHA0CEM7hX7PkVWVMDXVBzOxZWq2iQXCuWYqkkCWDrgLzQF4i3kbBMAt2PJH7cwD
2kfCWgzw6pShVeES1rK34qXYVrfZ1yFHOb7jwnPnMd69tpyrLLx0sZzMDVPb66Gh
5nTEA9Ugf+0gAVC/WX83+6GLPvOkITMv1ps/+I9heMcBVhoOypBwwVhH0YeYiATA
tckXahtISpqqhOGE+hqZLlIXm3eEuXI5+gXNKiBbyC+AfyPQV4FKsGgbsB8riINy
Sh/MqEffcGQSjThciulxQGlnFqEhBnnLd94w9cV9sL/CwTwJk2hV6Hr0+LvkF8SJ
JGQAr50AhaCeq7s+sZ2pd7ykhsUKGjFJVzUMhlQwRb0B3qcnuDIe8BkAnJeeJvgA
/2VlJ70m13mzybfjF7es22+vY2exPpJSjyO6aq2BtGtrTieTUrA7v/0ip9w+Ktvz
En3uM3TAdvRuh6pB+2pzVaggwMj84dVQl7odB44c2XIADqT6B6IltGtc7TC24MA5
ET0H7feg9UJJVp8Sl8OyWkZ15HiNVUagwHkw/5FOyrpoSWgZDDdBTtaoJS9TqYdC
nduFWJicuhjHVvcHZdpt8mM0bimedhVkqyQMLspDXWvtqY6Bdp47Zsyev/3n3Fzn
G5uf37t+UiLJIGWPhPP7Fa784LBNQ+rxE4J6b9jMmGNBHEAnM/BlzG/+7XeXWNdu
eZGwZVdHBevT5yzsNVfmcaYbeKZj8n5nFOAUPUXCR9eMRCJib6mn2kWtB8CqIr6p
Xhq3SBbf/8T2eVCOgOf8y9ANLj8m6O0ava+dpF5DXDBc/1W7kg881KD5EOIVU4Wl
uP5fURduh/looI/e3DnU+RAqmkIGTwI0xI/Gj4rAEv1EMmEvOMnxAkQCDEPJ2urx
7lm9MCDyyMQKn++j1vBVvHD9ECs0YELAxV6swEL5F3kdOGAy1djKTjbtkxImJtKV
FMpQApnhgMUpc46CiyhTFUrzQ3fo18TMt+jd5/XGWmSqG1F3NZIvDf5Y6W9hJoAw
TpwQw4BMc6UZ4rqtlMcnGTA88sZHidLwNiIxsq4ZFfjqopRooLOOvXtcS/Qi+uyY
jjrp/X09wp9vAgXIYJe77HrgMOQooCatiW7nViDaD+joGjqPRIp57Gvlk1b82FnA
BGYHwgjfjHRlH8sT8Kl4oHVXNqJJzcz1nTfYfnPyUgBeexJrEFYUnCv8kjRoNskM
hEbBa7UWEid6pWESMvxPc5LzqENqOsGQBIunLadFHu1hQJCUMIsiWkS/WGGb1klt
oJkoFzjF/LKhPiLqlQEpf+zVa1OvWn1XPXawEQKRwUDhugoHLd7F4aYI20EqNyXu
Kme/eEVC6A8a0F2eTrp6r9XWimDNBejlklA21sN9/a/zr5auzcUcSfvw8EEH1CVr
GSRIUOm76lB5FdErbGS0PKbGPWXGDqNtXgXWd2dNgXgfzVwMFIN/OdaD5GRBItA6
LsqW0GsRCRzrzFQeagrbML+VEKyJ2+5NFRrbkb8U9LinxTdB1uL+3sgwMThsqGMk
r7e6rnKl07GXE91J4oWtf44cB4LzvIKhYHqltsx5lNAG/d0MlKwC3GQco9SDOInJ
S0Ahn0eMnB5e8TyKVrP55iwFeerRsEvH2M1nCjxBJVFIB1TvRcjxBPT/S/fDUvnT
DAoHhcxDTnR4AdNC6nVvTYBz9E/RyoUkOEOrTHNflXWB1OZZqKS1evXtO34mhDY2
MgL9GhtEWBmVR9/FPOLYlqDhXhSyf3gvJ8TNsqxVupbdjgbIgORpPdRG4sPv7Gly
IkoVgoCylQELCHcHdsnGyx0Y17J669wyFGoeBqEXWPTshhZuq9QvoNHpscxuTZ6C
b08CPrzVQg/Fe+4n/d0ufdvodFI5Cqa1zmYcmLw0dNlxnmGRoFwrIIl5P40ENi/8
z7inbEwQEsIrKTHS+Bz+9zMzViM4Euk4A71qwiHcwl7Azvnf35NlQNi0JYRdRhrN
FzmhRF+X/Xi+ffLRGcVht0swKcB4a4iMsECLgIavh4XOKOzALDbFgDZWVMp6LPMh
H81/PhjzLTdw2VOh1u2FbP3YLc48upj2wG92Dej6ZiCjBcdsDGT01WNXLCewjOyW
DAVblu2zLNs2onIbyj+PJBdOrJy3MzEksp9RkkDOeLh3l8EG8VVmQ2fJenAZRB28
ihCNuLITGJExWIiFPLpqANQ4Fn2IQPuCbv8X3Fp6tME75nQVD9jGYpOKzFlg1AEo
mcb3CBuVrfE1Oc0qmekXklWO2obUQN8p+oGFR1dYpODsecjcdvwdBVCP+1VPaNwt
gcW5SWuQvxfqyy3zTmaIaaHQYdWctI/A3YTkXp/5t3R8j0cjVPvTZHI101v9oDOW
xAkcj2FsX/f3lv5qx2O5vwPqR9ESPCLV2RMRgNNuPooyRYpO8hjKlX8OxgZCD46v
DPN4m0HH9Sh3zj3leMN/49xYZ/xZQzcUaa/QQaXSrje7KhBsWxzrfciICxWl1Dti
MBhcRYRybmBEHcbDGOA25sGBxP4T2oip/Kejt/Fhy8TwAjJW690j8WHSlM0AlWOP
rxQ56ETY+unlovchYQp9RK+9tMqEW2Q4EErNuQ6XyboKa80tkCAStzSvyO53Fcsr
qqtlSSrl2GFofbuzTV1VIo7lMUxEXFoQyS0a1Y3ZklmDAasNwoKvxZ729NBCssOU
bA6R2yfe5KdJtZNkcOWQORSfn8eUw0PTqtX9UIuXYHJt+ZqLSSAyN7sMCocKap6M
7CcpMq2mZ48LjpZ6FByt8hRYtLBOUgDd03T/mm7mcNxLap77Kb6VhjGVt4nrlXR1
lbAZpwsYLYR5JODxM7O8i9QSH+catlSoGck1spig7Hc6pcZ3R1rmZVNuomNm5cJ0
85lmrWPUkGhGdbTFfvrTTu39eu2F7ScVfhyAiYE7Ab8mbaDmnd0fwLNBW9VX1YFP
TFiD8KqQIZ/8GBL0BQvuIqrso/Lu6kVhs4fLE8kgzWWAjK5LhfRd+TZC7tcEWVry
vY5dCUPaDOP6anT3vOo199VvcILNn/GSzW8xjlc5/jDSYxxaLX60hdQIgkKSF9VF
pSV3pRolpgRKER6CjXuh/Ysy9F8B+EVu+dgZxV12qKbrM1SKxJkpROBF5WhlWgoE
DzTGFp5mFnSDwjsLRxFnqXDgwFnJTXQX2YerTcIOApAkJbikHi3ps3gp0tybully
N0R31XCJpgFE2vvf6TAngdN7I23b2qKoBbnnXRebz1s99qTkL1aVAbA2xUnvbQPC
34UHm1iRaXZkD4w7q8ItJ/kkZVe6fnEAfFo52j5cdDYVf2EdQh67wMdM+efOuCPa
qXzqRFjMwOtuyeSmhrwjdr/RAPrD57KoWuXrh2u3p0LvRDCqF+y2fud/jN6Y76oZ
TObaOgKPmFYHEjtVYZXNu9uy4RkH65HlAnmb8LXf/EcoFD0SUOJSPhWbhS2dbLi8
uPcqVnvChfZ0TYh2mAUxa1rsOBpVlSZK2BTTyQsZRuKgvVcUEtiYeVsS0tGY/XVs
vFMD+SoJW1RIgr6UfOVhdhu8lFjgktpziCjOAvHbkO/uWf3XdPmnYW+Ny11Nv6ow
wnUTnxEX4RH+cmSixnMIeiwlRjFECRwdoL1tJ0wO99B/2K4CcrLQ0FnqaGQDia3U
AaB42rLwnyrunbAxFz/fQXM6Y9N2YQ1YnGpuZOQp7LVQRqqQnnaA5KQSMe5ZBX/Y
OmuSjcTPS958pRJ8rfkWXveER+K41KqH56p2VejmyK/nWP++3TJtsVlQDNkFO3fj
+ttEkkEab+sTjsckYtV1a/adCs1aiWVntWnJKwbME+4QDHtmc2z2s0PXFOi/5Ym+
5l+OHq80RwQmrttYlGP9vNWWScOYHv61VX1XIht6qKs/w6Shf/gBdB6jbnqV5Kk9
IiCMOpT62ta4euc3pk0acyGetf2qJyhVdgQo+H78wvFi2iZBfR1raAScz4pwJnyX
wWoPx3d9+v+sbACwS7s694JW8TEv9SHAh6GyNlyaAaDOqf1JHlf79ZFpS00l3w3D
TZ8U47mqkqdu5cXPF83bF19pxsoZEstWSlrv29QraXtk9Rg24WNAN36VLlYC56vS
hPU7i+zhIRg9bUhrvsa+ULYN4HnBE1DNHl0ak/MvgCZuMIbkdbsBqZXoH3KZR5e7
mVyOspFM5wbN3fZD2jGeCEH1SgR6RmiESP/dKyHgMZhgqr2Eoc1Rcj4cIiLOYLUC
gkUef4TAvT4DA/LBomxtPtR+roynHAp/d+Zot5FrVefSosuSr1OLxML4OV2Vs7vY
6xXzpatu90FzrNk3Ybg09zJbq0EwlemRr+zO7hSsEyJ9KGVLUqKp46y7oOu/m6LC
VaWXd5qOAdJ7oRqX3MiKtIS234CC+C48Gxf43yR9hVWx1V7n2L6STs7GslXmGNvU
LHt3Q09m9nb9y9QbFbAjKxGqZwVAAShm9onONhljh6wiFTjF20Pq1YLOnJ9EaHr/
HGld0q/zF8Si0M/eQ9EqKSrqiHyrSrZHmYopmhxrkUwrd6BhyD5JikWk9HMyXnDz
E4LlT/cZ4UfD31DqUbDiUpiJSoKGxeH1wBAlXpCx1yN0Zgqaf1WwYpO1fRWmAj6D
Twt8q+7SmFIP0zZ9AHM/tXADepLQNVp/toZNcbWoixg+84wE/O/ECnQHKpzN/LD/
fSPQPos8xvtjGY2YtJc/VZfVTtnwTO8MQR1FCd2QbALJr6o8Z0HDJUwO31WdUZ5D
oCtaN5mMIk2+vWeCYx05um4qHT3oZxN4BB97WPYMS1Drs9mdGC8HuMicMsGoT0ur
UxiKY0CTUzOw8arvmckF15S5Nco+SQ7f+TWe4gl1zKUnAzw8/BXtVELWqbfGRVTW
SJx6CBQmdMwMt2gr0xjgdAquIqvxQyTFzcbCu3BNG9S7aeMVa5rBK7Gj56aBIQNW
rozReNQjplRLXIsurhhrTRRu4cvtWHFWom9gi34j/B62zVNogiBJCLMLBrGRFMwU
XuK+xUqRkaNUCBCiXMzf9yNNptRKoz/OgMqWHhVTjPZ8Z1ijAa1VqSI4Jy8h1+hF
xO2ee75xU8h/KnFiHakoC1mwzB4NdULoY6A5cgb4zxCcDqqdSwrHTZ3B1JU8WV9h
NHNB2sT3kt0v8l3SI3OYsFTIhydMy3PpjIQVyluIiC0dpwmUewYbbNIopoHKkd6R
R0XRlYIAzKHbcZ03o3+k2Omxl3Y1XViljkhSlFWEguJAIJKfTgYJ3rqjdAQCQXfe
DEUsUrJi1CPq+7n6Erqv0c4lXL0Pv12HPfsU4BHyRr7Iiqx0/F8InTcUw59rQhgk
SRGpqPiGKg7kIobDDI/oemOpsw/7oUWnpRiglup/f/bYI7LD8nQOCbdfv8kJ0OME
woIEPA4jExglhBFsA+A/vJzJG/dpbxsidAh1AXUwNGrkXdipJLoxlxH8jhMPVyEs
6MxlJfVuDNwX7+4G4Jjjv18Vg2i4GZJZjpC4fEaUPxLH4Gkyoh7P4ndd4Mr7j3VC
or8+cqDRH/Yh6PgjcOtNngC4e3fy6ZvdrIorFqY6BKu6pgxuCfsBHAwXu4yMYcsW
+uPOUp2pJ7Ct1Rb1oA3ql6X0k0vABazwJzz1JI/KNBjmQtLTOH4tPf+DRO+lzN1A
DVgdpviJsmyaqD8htqiibOi3TvGeEYKzcD5rHV9Ydf+zDyu9ue1D5SURTxiHEnpd
j6rAMMT3SyyGvd/9lrxt01abnHozKn5neMzjoOWHqFcuH8kj+uADC8CDW8UFKTDv
44YvW7WMk9mQb0mVru1tYGmSfjT1fq9Rb2IETGLvRL/1Hpyz7qXx9C1MMELiST8i
oRnIbLTzC5m7D70SvySMG74SH3J/7ekkcy45j+LBW3td/vRX4MHOnJpT4xvJLKne
szK+BptB4ghtORPDE5Bxo5MiRTMWXLSmPjz6WobpAtzfiypoDBRKBXq0FKCAjXUO
hKq+x7fYmtD8Zoq/eIK0anMyrhZEp/8Cu0ZdLIF1ucNL6+GcU/KUAR48qU3Ey0eQ
vaOnsokzGohc9j2h3RUmUK/ZyplwW8AEG0FgBQ1gGE5UEKlisoEJAiIyod8tbspX
aRHev+Jyq9Pt5d8oKwFx1j5rA4/IoIRY1uNJZT4LDzXqMMazaWynD/ezt83WqQc/
KgENf2dLvJKbe8FpmJO1YpuPbhLZ8B6t9r8UMAXWb8Wz0923xGStlQ/1mHn5cpTD
FXxZ9snf0GR/Z2yAEY30P5sau+DeyVvO1zokIHkV/Kv4nRrnMss7mK2lXr1jZQo8
ttyCZrYJmuW8vwzVhb++1sAYKl7H5rSlTe5NuiMo6elVNgtU8QptK7HOlbf+OzWK
keAg9tSA3VMMSrvjvlWzGFjXnRrpSeUJ6nQEoVdMNnihSNuQmrWxTlYEUx8LiiBv
yTi9uUbZZsK17ZND6nTBNsOYALpfzSL2OgOf1o9Nr/Upd8JdlUjRvw0WGBvnlkOA
rlcBy5YGVzcKEASsHmoOYF8NZBmVpjUF8TnvvN/B0s33lbIT7ufQY6lnY2vPaTnL
NJC3BOM7ZS02i7H55lQ8Sx7dJ/QrLNucfEnbEJcNrsDLj+oYKtjyyIjGz7dtslCT
eQ3t9FSjzNN3ajle+LxbInvdjdSom48WNygGKhEaxYe4VPYwtc2mkgeBi2Cb+kAZ
sSQLcsEVG/fe5/KpQifOXebC9vUazfL9X4BFcB8SSpkDrx9AuIS2r+myH/gMpdF6
RA4urTjIMd8Kbv93fYCFulRvrZniZcV5qBUr8sscwBbicKd8DGKtzCkVUwBjtaHz
4Z1IU7383JjievIaSmiv6uaUDYuBQhWXl8qrrY7DwG842xYXQZxauaQfBwr/AITs
6IRgWNRJc9jxXtNfuSn/6I7B61bUdpdFb2eliwAvP3sC9AztheaLgqXnL+1ifXjh
Tv9Fs5uYRAEPX4TGTToUAlfHUvhIudjoTnOAu9PiW2u+sUN5ezScJloAJI4Zklbt
so8sAGSgKpjkNPKTxJvk8kL0S0KcdEs93BECU8+zMo6Yw9q4/TL+w7fjX61tku8V
hZilVp+u36yEd994N/I+9ei0TjYEvpbCej0CbBZjau0rCATzLlsQPlgPAlBOAfMj
ZRqX+y2wV27XGGx3LFg/KEe9IWmnVigQmlrmxmcb5Um0MLjDL9it6sTYxdZi9lXc
+fuJyjg3eTfFBZNn7K14mHAGPJ4GstJR7btM3uSIQRsoVloheR5njNcIkr4A6g8/
lDvrm6DLxKx/RbhhL4zfHvtUHKPQBdmayBoNaMxj3gl9iiHlKoj/ASh3F1VoxWud
DMa6NjALjylMRktoX0NU+aNoO4jRZBvTGcXxPU6fK3AB8HbmSKiqwcx+ZP+ngbMM
bS/PgaNi9L5NBFoZ9tf3wbWkUFV408GZ2C3K+wyq0KmgvoNumT6rZjlHAmvJd3CP
sMco+kshkx8HQvQxxlAwXMlyTMluyNGqUAEvQylDniLxEGGoRvxAhZp5F85B4vy0
qRK+VqQxU5KJD3/EvbQveIIn5jlUjWt1BzJbAdBDQ4I2P0KJzaoW333YGLZgLVwH
s9vGd/OO+s7DFWJdPJ2yYD1eil9/+XVGLjgZvKrOP5X1bWJsmJEcdpVJL235LhLv
kLkbpDPkcTwsT2Qzxtvlb+zjU21LwnN5fa9MuJJfnvMNToIuArL2Y0p+L47rbz1p
6VLv71DUdMauS8kafbB1NlSIHHaw3RBUQSaO98TVGfyMExiM+hxp9wnDOmS6Hg3X
rc1U1FAyG7RnkpGNLn5K93GC9ZezN0cCZt4CbgMQFUuUwlhavUjhmzOgRiXyOC0B
e+bm1DN+hxX7dfKpXpMfxvSYUKJjcvgzedxGFJdHZAWaTC2arKepov+5JW8EZJAj
PJ6EdrHzlIDpMgyPmt0LLLYvylpvu28xR4/oSsq/XMWefuf6AIWKr4fpGGplduY2
ErU2xblD9adyMk5ubNGmBPrR7gBw+eGtWwBFph3BAdVVZcVl1JWsrKO7AMVDLqKX
zw/SWm3dDT7YeZVTu0DU0bTzWAhuBJZ9dnASsDF0SZSvEjRP9q3QNKFGGRt6e6QL
/8T1Vjcin8KrzshyMd7jnoJXOmNeF2NE9yf5c0vICx5EDiuKiWy2O47v9jIr2bmB
OJlZe/qXo1N4zLo8QQ++IQhxHCGOM0gIThpstd1EuZ5GDOMt4cDqGXoJgD36j9Nm
MpuON9N81X/VrZc4bOeIqrXXd0i9yKLcViYnVEuqq21R5Qo4/138GlVpGMa90oaY
QI91ZdtQEGQBucgKLg7LVviZXzBTHdVE9uBMHyZA2/48yebRwhaZq2U5XPtpt0I7
5fk2uLWDzJKdWF2jYdyKOUi2mMYjDPsiP9ij9vfNw7bVcC7vuaewb240dmP+Lys1
5AXMzvwLsW6GHmVFx5668q/87k6DBjrk1ggsv2+9CcfuzGnGxawSdIAeH+j7W6Bm
slMLaCfXyE07m8QIY2evT8NTNOTurOR6jzta7Ig46cRVo9/vD8Q2NBFvzdVI3n8Z
FT8eDzRhH973P/SBkPv3psK2RCkGQlpBZWH64fgFdJX0bTvOohMoRpPoVEskGGDQ
yZz33VjAva5PyzTUtEzM903ejH3Y9LCTJnbuD2yy3CBq/1boi9JD7HmN25sfJ+ia
tlh780+oLGbCVmbXfd+oLygRwugRdB913aMcChgUgVSuc8oHoWYOCLQbsabozaii
zg//5vZQQzBeIaPpvN5aEslmmED8qsgXDc3XVW4dLXztMngbCSP0WjgYqFxrh0sA
N/tiPEFwkf7dopGEutrxfC/kXMiks1S5JcRNObSlcZju4wdqLjIoWGdAzwIfNcG3
vzz9Oo0Csqt28o4dhpzfLwSPNeLCdJJdawzmWdWi605uQCuFcvx2VPLFYu51bWwr
GFsLDkZC18jpgtfDbwWS8Vh8rNDYgycHCvRcURBdzGWOkQlEuyI8lTxGWCouUH/M
LMmzp5dMjEC9NFmVFuHOXjD0Kc78MlMP9Bj7RwIUX19plJ5vHHpbfPrRYZc5j3Jf
AaGiNc5yVynE4z842Sdu5I5U8yly3tAi73cp9bzXRwnGlXz1sEkazX7sYUztkTYT
QqHtKr5WPDoYT9nuTuYWBvxMrqLapkXYXjBZGwP0vXKeKRqVlaPbP5164/m65giq
h9ochk2nWMZXAi1Xfm25iPs80TYAJcI2AdTodMlkY55AofbmH6xR0Tl/uaByJP2K
Aa0UIKda5PQpxZ+1uNr6S+gj8l5t9t3eNLAJVaFedi1/cPohtKqm0b4tmbpDTajC
7fIHGclCaP6JIqINA7ZIlo+AoO0u3NKzXRl9YMJdoaRCc1QVgkbzTtd2uRR8jK2t
+KkTKe/7b/qy3DuYOvRAEE1Tn8yv8rvWwS002j6v7v4DP9w+TcFskJJPShcuXtli
2kF35IaHgaMLuH4ZF0dkV09mc1i5Bcp0iGKHUaZXdbCyVmLBmNCQRnoKc/SQL90Z
i7Heg8M1hZjoIqPLtfiY+DqNftJLFxpzU0yP9wDMaJuA7VOh2sdKioBML/sywC0T
Sxypsxzfz3BCFQ//InV3c5C1J3PC/Z1UGawOfCMQ0WE7xEUmuLL43cOqCp0Og8Hj
QmA8LcPtCSeHIAeDBZMVHvpziZh54HZVprg1tsYSNcKfSxfYhdWJ7GA9cspfngug
HzEL4dmmW04vRZta+8rw+1uyjJhPZW1rA0a08Koe3C2eBFcJaZV0B/3lmi8jY6J9
I0CCScPydYChxXCHNy/1t/FbKbJAIWqKHwrUCMDHEQQZufE6MHN2t4813aNKTPL0
P4gYXB8oows9gIxaxjyvbnOfNSiLVpyZ5pzQVUIckoeCz2d9cPrnHwECp75EdeS0
5ozi6704AwcLy6mNt5VA98PJq1+gPQa8D1ez7A8gHUPQHwgtWJGVr+7GC8owVDJj
0FVZeKPkidgM3csGQNzYhT7RZAZ1oX9OS7g+Y3Wzt5JAdrQF4FrCcmYqUwfu19P4
DDjco62u48OSwlbsQ2PBV3UuaWFT90Ef7mOsWr9sdarMEorSBkh80d52T8p1bVaT
yMZmpynibCVc3HSmxqqMU6xnZrJCvjV2fJ9r+gQc4NaQXdXMhFiX6TW273kozv4J
EJX9NtVKMPPFxWF4/DSttdHMSMv5YW8uQJDtfDPgoVC/TnPGZZUZpvpAOdbJyvmi
sgMkgSIdN8PT9527JBgMV0kFTGAe/GkR4iYVnankgjlssrEhhRUOfLwL6a4VgNx0
F4WL/yEk5ukIqwLG/3xhLhEW+OKfA354xeb7nLLQ6J7SLpeYSXqjuph73p5lNlBL
PGusL/0RKp7kddYmIc0P3vrplLPjwQppryV2VbgCO1MyliRNK/MwuDq8BwA81KfS
VAe2X3Q2OOZ2oOFVuPBkxUVl2fWY87WQxLvcVRrzoDWsJgim4aXWB+FevwdXnVZg
Jrwf301xCI/LW6Oe7WpOwutkFQOC039FrI1qqvciB+jbMnwJFbqfVfvRdZD1ZDEM
nX8YVDhw8Prpeo+m6QXD5rmfyjDxv+qp8ZORnn66h1/liwSDwrER3DT6j8sDE/Hm
0VIdp9AdBHThIe/P84FbnoIJVyp08mvW6hAC1fZ7QISTlu52T1KP9JX2bgFth/Ux
xuZWsNz08N/bHDWkhouAUWZNEteNamf7w6Q6mREyY7Exjxo4er/nCKbeGBfjNc+h
JKm0E4/Fx3B9H7XKdSeQz3uo3u9vBFONr/ezTutqW42XqJVPL7Psel2dwX36p8GS
YnCKBgt1r6//NP/MG4W5ByOtI2olXFr+mcQxn/q6dhOKsqMKHCSwBmYWk8CfB3tY
YWK6cbcRZsLBLwcGrK/VEnKcwFEQASEKNd24KAOG1BVAdbKFjOz/R8Cojm4DGGwz
p8klmYxMJyGS6iWenSawLxzV9s1cUZHqd8DL8QVEf5Ojmu6y8PG2kQF3d7yebzPh
9QD4Fgqv2qdCqgC1J5NBVTepdw1gEWyLEB4hKLd5c9NmqkFovrs7+JFDWhbWq3XL
N+cUFSjbQMdByVcAo4Jr5bUiENGycwykABE31mt1hAQU+TzgFtM/IYLqDeakjKxg
EQAeMmgGT6+vAu5zwGcSx69tzDIgaorIjHYY2Yojd7KQTQCBgUoLenjyy+1y9zEJ
nq2pGXOe7i47+wdHISWwlWk9k6kDFHm7hIQER4AH0teUSBdYL4dUQb7weRprt/CE
8R1335ZZ8xwiA/ApCCVTK7ebdzYP0RSTMt+QNAQoW9i8o+usI4IImFwqNXCqSXX8
KN8Zs7TP9fwTVjPup1LcnMCD+BuFAe7DkgMgKDURSi1fEyHbQr+0UByzOiKjPUbI
7VesjJBXY8YP0DchVkduQjxTqFYbWQJJ2idfIcyWkYab2LkdLjC7RXN/vzLSvNzR
Z4b8wEaTcOYKWQtJ5p/uv2VdYS893BUotAxgEnBmVkBxqLFyiKm7O2AA42McSiBG
s4LxbxGOgZzX53AoXC34D3UjeTXSc7Ma/SDJE/2sRvQBRZ3sB1HC3vwNYR7yyBCN
tBYuQpKjmqRU0JFS2ZgaQumqFxvw2DZ5hroJq4tDD4pBMV7DczD2wv08MsmNheIj
jQKr3sLA4lyMeNyVrXGmHBb6xicwJlUwHLzGcXqwkLLFeH/e470QaNhzDrJuOG1K
aiC2wGp7qaAYtt+rV8zScT2mRsETnPeevLcAXc370ZHNzD2q/coZZuTIYirf0bIL
QSkF/xwmnsLkzmcovT2I2zZY1ofrpnyPmb+TphWgwqzmEEUwLTVtK0/bij16RZft
fayY4LdW+tI2Yk19ina89NAE1RVITZ0+3q+hR3PdqQSnxrqA8Zm2Pfr/jJTU2hTz
Ny83ozNjyFwSVbF0Ad+9joSSr1zDF+C6LFlvwnqk07c0YDGY3evjWQA98iwSTlB9
aBXqdj4ubhXBt4v8hOVJ3TXUy86LueGafMHp04DQy3F7rm5IQgxjkAFE7pkjb4VA
au46Ye3euZSUdDD6XZRn/kW4BgJulN8hjMItfyG5eMg58NJ4c6PAX7UAFujxYv3S
obMhR3bEXrJKbrjR1hhRykydKyqcYIk5Nxq7PjhZ9uKW/s2V47yTp0Ghdk5iKnbb
TCwA7Cr3e+9NE3t6/Cs6myPoNKEJWUQhtYMXtKj+WBVVC5vuteE2zpSQ4B+maRJY
7tsvKbqoyy7tj9kA6bQhTMdRXd+OVu257Jm13mDrWuzL8FGLM68YlTseJ6L5r3+j
qFPJFQtk9A+P8QjEFjJryW4HVyVghVfgWhbtiWDNludQSArezBlm1tH31XobEkH9
87YxixBZwxpgoGeHd0j45DltlFkTD3AHJuaDSa9Hh8gVoSGCdiWZrfW1rBGV8iX3
gSIYmjQqCLRUirjeaHUV90K72ZMyf5+TMWNVVDb9g5K7K7I3Hz3svXpXIIB+CXU7
6IAPRki4OPJSKTUNfG18i2lwlSvfnYJ9sujqKmhspR5sQZaHbrUQk36Jf+0QtUSN
OS4uOi9we6FYNob3W8zu/rRFxaWuPvY74AAsm0IPH31trMbQv+DrVEmUn22zHXav
mVGfi4uT5umf83CgjbnaDWgJB1EYRyug9tvFbqjI2UH3342xaPSasVwMN1HeCUVW
v4Chbu/u1jCV6jUvNFnve1r+hMWrUXV7fO9BUJWzLuAw2BHXpCPNFAnrV1yuP6CI
uQNfp7B05Ux3apyUKENpFyXw7t1mb97V++Ncr755XeiYsm7zeYpPQWh9y+9bmmLY
xCve1cYyQxnt/JfCUOXHYyDhBmzzIUaR8v814X1aqPiGLXoZzlg+TU9+fH4kT7ES
jObeXLgLhSjv60ZYIjIm/ls1vd52P8Y+s4OGCdI9RzrNC2YOWcbIML7YfEEHtnHV
gjsoPS1RfpBfej9aWWXp2HBfcra5OPmeGUdmqyuLnjpqB7LqZFoxv2J/0BZTHRWd
zmIdC7HzLu88jiM5pOFwIJuzVbfp5xJ8v2nURM12O0wZ+THu7bgrsN/EV4hSIf9a
QrsaVsXPibrVKA0givmcpzMWvSg6hhRkXBwb98dEqPu5wNpJND+P/TVqowiy1XYw
0PJEV9QFw0Tm7hNN/fXXdz1bGTsQVeRHAPeyTwwp2VPO8Fu6R8HvvKjN5FS8ypa/
///ZwHwJfqxgq68lcYRps7Z632m230TCPuHq4JR6HE628pZfPjAjBO80DfUNwib2
FIiI8k4tlmTYhsfLR4Gx9w5AgEfX+DtqcyZZAGScyQUVkQUt5n5haY7yieoWSb6q
qKgs+pN3EGCUi3BOyAszCE83+ODjhUaZyaYhopDr9Fpvu1+fptJD0ia2ONwZDJR5
dGOInGGU7FPtu+rTtualn0xM12l7CXiU4Iq7xLC80599q9dHzSZeeJ20qo8NbafX
0VcF4ZHWOw+7S+3AvLm3fRf4UAdKhK7rV76PhtnWEfZAzAAA+3uYUsIrQBYxBdIy
G+1NHPtwjWs/BWgFvz4JmrpNYNJ9VMaqCqP9QUwFcxcIMwBtS+SbAyKYzwA/1cSV
iGJVsoaTwYBWHvW8kQONy4fYSYeUfKSEnweDR673dYtLlnPGF2JIYwUe7AQybLCP
LLjr8TjtexRpbzr13kjkx+OBcmU/qo2hL0+BmmviwQUyluODjoZ9prwT+qLKcyQE
ffDoNxZnWfijOW1lpNcrZ60bgGO7uxZnajoX8Bp24spHAeRV6zZnywdylEjdjp3n
8stmyXaF7zRHwiPKx1uYmO3cwC6jif4vuygYG1Sc/0CFlsMxni7Q6Ax5UEipuBQQ
loQew7MkajD7oP4yP8kLbiBUD3z/T5f0oeAi4Jvf/IekbSoMBJ1p17thKx3oKrIw
2kUsjIQGVg/BSGX3irFe6HD1ZjHuXYQ287W0Oj1bi79rxIPonejW+NUnXg/+mPQF
GQeREe6eoxHynCvu/MK6RLfmn1EvXqm7DOOIX1gHTj8Gvct9DKkwqSG2K0w869Gh
8Dt9OFDJRTsp9MNrSFYIgdS4aAgR9/y/Ru5by9KkuX1v80aHtKEqqz4j4nmU7N02
Ije/3E+QuAhsKR+YOiSqJBaI3p/3kNHwjmch3cVd+Bmtws4E4XhtPOn+vAAlWMEX
RhxUyvzsh44y4XrGSkPibLfE7aBvL9/R0mPzRyOsaCVrwoo9SB7OS00P+QbsOAKW
Ayg/RyrqxpCwZV3tcVDwitsAiwXOUrEVyLRxJC4dHLtcQGCLCGmB1pGFJVZBc8pe
qmXNKsS7eg7JzEX8uOkadk9q/Ta2UiyQddIb/gFQuH835YXmdqFj6RCWdg3FegTO
k1m0yuNQz5puExyD++EK2fLL9LwRHYm9s9EU3t0j4douTnmzFTHO8a3BLiQ9nTG+
BRbBGsr34yf9KMfuhmnqfB4oYIWHMLdYmTMlA2iqtmd78qEt4XH5SN8835bnANBq
Nso3rnxFqu3HotYHOR/Xn7Ixln1ueblhanFDtnpTtq9JRqD7/8OcmfiR2oUww5k1
yenfa2G430PzkxD4EANUxObqzkoBzWTM1HB8YHxR2y6HreSmaGRjZ04fsyqEf0Ry
mopXmXEroQPUJwCAA9Qo/3JgiPmYJWLMvzfm1U/RBw/uhoV2jc7Bjv++PQoWU8am
/8UjiJms4y74kWbzjkXxt+DJDXUE3sQlo0UPr7HKFg7dGkIZvPp9TfPKnFpXZEBx
txvvox6sBuu+65hTOXbw4SZk3OyI37+1zDYWq6aeS20RvGajKaE2ItXrGDCbtc2A
fHQTGyk9RxqaZVZiy3gaBYnHAoHtZcUgHHyC85NrR6a7yuGSw7Dr+zrDdb+2krpD
kl3KsGW/qjCXaMtJjcjdJ5g1Vr/WRQ3/IyDxVjRdVMdn9Jy6usfaHjUvF97ul7xR
+dUAKj9MuAKj66aW7ViV5nA0HMh+aq4yEHH31ZRWOSkweesG6LYn67W5+hF4hAt6
uijD+pVG91UEe/vTg33E0ECOdc8fcKvpqn9wLXmOPwkh0yWtulblypTgDuQCjTi4
PnUR6DVY2Yz6nD0wgflwXE38CxJt0/Qv+xpSXUfRFc/BRGM+xPpa4UvJCBetTfwo
4yOlQF6iV48TLlzpvGobQTBs16nTr4gq+GJ+Hhd2l5l8F87jdzJVP/VuCUduxUBA
XZHcoworWu/oIfKQb9IOrlm18dLaafJs0KB/PzWh84+zyszBBnHK9KSaSeRNpl/M
cq6OyQO5sdZoH4klPxY3FWhXgfml4a99Ov0LfDjBcGJeKWbUOsVkNFKL5JVWK2Pf
sbW/cRzA5Nh4HmSpZ13XMzUBF8kLjwZN9hs6stMdAFhgS1SAVIT1YTj1gGNYV3Wt
CYQaQLL/uXvhI1XZ//8BwApssMJo9xf4dz9o+f/v1K1wKrhDS9Mr/KKf6HwxEX4d
D/VpZpg5KfRm2zuBy7I6vnp1O+Cl0lecXE4YDZzfY2ROQ5Y1FFLeS3CmkaxO6Aza
vqw+S85TV2iXgFc43LdLpBpj9J1YMQZWOyhGpAOZueC/tkyMYzhS2X7bP44HtbPz
mTaUcrjsLcuwFgQ5+PoNkLuy2rdmlvrB60cKn9qMTB3GAyghqz6yPy6TZQ/xDYqP
f04p/MWLPcLRJX+0sod+daXlA5ZKQ75hFd62YWRuTIFRHiVQo3mEfIYoxOjJjLXf
ZGIqpATO/4muhz26CMVmW3Izf+i+9NTMxRDQOHnv2YGwLR0eyv//HykPPEpQuWLD
u4xxkU8pCCsYSHFTr0QI3jAr4J+jQvQCWzjnDr/+GE/JkTRM/psZPk1lEllBT+Z3
GMYx4en/pYNr0m5ilRFU/uNMSNUU175cfV76FtiEKSx78z5kY53MXXkGcfvGPQXn
vxw02g7oxaYRlxKHKAG3RVSxRcmbkAK4iJqwzYhZCGKLJ2yIzJ2Xf8DUm8LvaCAR
X9SbCBAf6mSzQr1nuwdKW/czEwv8MtWysEz48x9p8RjEJsIBB1fAJ3v4TIKCFidy
ifYKR99NnKVD22U8X0GPLwvwVk8l59ZMQeU/j3Dk6g/xo+2HZs7eybRKQIxqN+K3
/cQ1NjklzrPYofNNJ4pn3mqH7HE9+jTqBYQHeDslPapnMbEYihGdmRIOPcwMefWQ
g4myZXrzH8RdkI+uDM1e2jr4ADN8KG/sWNSDnqa2lht1nOmXHjGPJFB55shPFQRy
nelC8w+JxBQEfLUEXzleNTJhuCOvW3xZtrYNoihDiovXp6trFKXhTODpIW097g3P
Z5ZgtsZdRvZNU2ldZRmteH+A0SFeb/5eATHyoPrHeqmL/xwMwxgctifJltjjSrX4
6JG/5IUoQb1mXnudpdCeZIHnjaAv6kzoxvZf98ELNrEVm9ug0vtB5mnzlxJe5Aud
f6iFMeukLdWFhb0QImcgH7sL1ZTRAqvIu8kaKgxXzYOoFSO76AFJMEZxfwUg8C1N
KtHcgYo33AzTBUlP3wHD7c2ys+D61N4Ws8PsO9h0qOS7EVDoBUqmrhOC8nu9K+Wj
V9MbfdZ+nYmcR09BPfrgDNDvzZuQtVkJm8HGoAVdfHzZpY8hVn1OZIkFHIOBmWmc
yuEAKR9Gpxlsg0YcQgvv0IC8tyYiHjPgQ2Hkp/ziQv2/4AA+bYcYnRcEy6ujU9IN
F0Sf5Us7/z9h/lf1L4K/xl2yKdITf8RWu6s0+Mehi0fD+mfqb/XQY4n2eF/l42GG
3vpBCcUExCAYelxuskKfg/2Ydv6t6avcdR6HpqhO3YS+F3avYgCj56TQksIG88nj
xJzOBraaYJEsAZSKKXEPE33ueWGF8DYpgSgPLjqkSXQbje4r4SLYHl5lillVDSgo
B8QDxsL+1KDf0hW0ejhk1kdm+Qe0c5KSY72BGM/AOqhrxcRYP+0A67BR+Gs3lZpC
E9yorwnSDiO6bVhgcehAxJJbHXCJO2gIsp4xw2+fjf+9idP0gtWTJzRugKh16Nsd
AnPfWZQngotpm5HUx0QCaW6bihHB+5dd3wYVYwZLijtNUSxJqsRfdIaCkJb5uALy
X4WjN1NXgrWJdP9iI8lppSukf8P2YIdfQsZeOJ3CSe9Zm9UUMgVuKy13HK3t6hmc
qI9zVnFB8oIQiAYFlEi4lOPGGq9AjSzoPFwgSS7qXE5KlSFNEGbm7STjNa38EfZk
e+QLGNrKTm/YdRR+LO0a9iJKjljy30UH76Y8+yrZu4+7VUmnjWZkXc0n5B2X/zRq
WDFM6GQjY7Zb0ua0t/hv3dF8/3hDjo8MUb853W8QZzh1pNy/xxyOE79SpSm2sbne
MJnQeH2F1zLTztFkElCpGbjFXne8V/Fswiex3Jw5hOfrzPejAi36jHBj8x4tFYkx
oIWb7RO91mUpb9u0VN6HUJgLMdKyg0rqp1noPudihimgLlowPetpE8DKsSpo7MTP
EhJqGl7JZcgBhWDy3IK4Qe4nxCOpN2blVUFC/93+GqsAvm4gqsdgtgrnxHZi5Xxj
lJ07lOvCypq8YmVSfX+SWRxq7VSKrZoKhjG6igmrFi8ru/RTC0qbSoYropI67EV0
rpTJ3QOC4SfCPFaiRVzbSQDnef6S/dhT6D26ctdRAvtleftNXnBKe8k4BmoVi8rh
u4c30XNjmyByrOdT2ICY3httm0wFeT6AI7v7k9th3MI6oLXZ7I7z4IhfkjL3NLZx
EOglQ9cZw23RxrarWD7TM7RnGGda/KgsBs9UcEj4Cs51X1z361S+QqmuE/qooThS
xGVehF/6TesT4C1xdG9JuTj3P38nsAcHDpW+FgFahzO44n/5k2Un0kHYWDmLfhBr
yCAvc7UK6ySpszKR0uwE4st/imA6yP0eYXHcb2wWO91vRpkes4oUcbIJ98TL7Wdi
B2LcOpKrTnxk8ak3lz6WRUgn0y8UM60zga1qGW8tBN8MZDaiXSSTlcASwMo8IE13
k0xgaiTNUahzEi/zWcwmkE5jRh9GT7uLwDPLWcXS0U1crv/jRM8ZZ9s6u8+y6gJK
EJSwuDhWtNYi9BE1weliBeb6lQapGaw45Sn0p7c+PwwSEUAliKSFrVqjBYzMG+q1
0S639xA113TulLdlGoL8sybmPThal6VDd9NP94a14lMzDWWz0Ym/k3SMBDAzXc05
UV/2//7Aj3BHU4RSmTKDBTkKX2gkiF46kmgCNJKhMP6rtwgaPc/iVQV2G/ZqQNsv
pG3aYIthBlM6rSDRWKylK50lLV1GdS//qO1ZL5w12WFyxAU5gPNZCh/ClIlfSQAs
00dAWocCo8+Dd54IktLRW3aVvdQCEbaDFSBx/ouhsMlvaHtbeDzw7kY+y/rPej/z
nTZ4+u4AuG+R+M/mg1keOOgLQHJ9R9AMJqUJQZVNRUYFtZJNvclIvqmJMx4MNM1+
CIGcl4I/o31c49/z9iPne7CdkbeqCBijNRyBr06t1pV9tUNXtJ/q3usTttM41fn3
ZvfL9Pq5GxKpe5pHz1FGoJd4xCJwOzMYpPOOJ/ZiypO+nlo1S9VMK4Ri0K44F3ko
6p1Fa4mOO8DFLlibjof5EvVMiiexNvnvW2QJHS9QmQm76wMECZ2VoRx0MW0ES8dy
7t61Wt3FbnupCq//F+mVqSu6Bmt5ouFBOHVqBcXbcapulJSBDy9jPZc0TDPKG0I9
a2dumMz/W6sgJfMTbpzNBMrJL35jmukPzbAoHDSFyCP9Y2aDDULIx/03wqDP67rV
dFhe8stnsVUrvi8biaggSB6082SlNZcg5UWQNJ6QoVzXseMsG2citQ5VBKt1bo5T
21r2fUOs5bJG+6tIAhyac1hkNRVHEwfevbSFch4D4YIRb+scB+ye6539ErJ0AK+m
FYPPs+u/j73FZbx4VKZUKMDRD9sVyl500yDp+XxcA81N46uc0E3VO4T3IasiIjlh
ewo4Zsp2lbaT4n49ZsXXVfdYAFrSxxZoH3T+zKAeA/VIL4/wcaXyZ1ISsGjLmbhh
ackVnPAKUkGML7zeXTsIy0j+tZlbl/Ws94Po1XiaMMtCKFKsunM5Ypc54NQbCTNE
sdxrXI+cr30aI4rNlh8U1QnwLSyjSoh/tcQltbYGYXYlCVPc/4UGFZ5Ktopm8e1F
S4HJq8ggdVM8+k5adsW8yv9us0u+4eipDLWPDV/rlpSvMUfcPyWJjpEEaCAZSbXy
zQzCthxTRk+Lzqoh1vlx1uEi/iVgbrY7/sooHggDx2gms8Pjuo1ie1L0zDRi/IFo
jIGfAfClhDUWwECnifYjJY+A9UmwtTUPGScfwTWtnUmVRuGtM4tsV1RBJn9nD16r
JQSeoLeYwte8C+7IgGsU1IwrJmuwIoJCp8fAN9zLByyC3cXUNLUEzzZC0CWTOdQl
JPzDH9uNNetWe8/F/OM+UZKZnUXOVS/NuB5aMx/z7tOY+1AWAq8Ljd2Sh2er0tHO
dHiNgfXDp91gcljxFD9Ees0KSvDkdqGL5wBCfopA94jGO7bLyp/oPwph8b+zY26o
JN3R6ZtiOajRE8cCeyv/p/+E8LxddKSRGE+5weN15oa6CalErCwrf/gisRl55kpM
rl02nscYLKSKLlHxXEzuFyi+bH7W9koHfwudoCt0UoUjMGlucMmN+OcXzpQcibx3
dHA2ptRFYtPVz8e84/z9htUjWBoR0w2q1hj/ubaVepEF9FYYImI8Hya24oZli4Qw
MP0tBC/vdYdoJkv/YeIPJss5hOa5EkXkgQ14FC+FCJdJ9a+Pc7fwYkzdi9s6ik8I
htalWJ29Strw2EtMxY44qSJ93RxVbo81bAiCq+tutLXZHxDgVBSu9CxAukMpYLKL
8HUuxEIF2T2IhO2a8rGhSw+ktO9tUpKMZlhaITf0yzCo9HBwcX8KzSoHrpHtQRWa
uStEKlO26xlhiqS/GR1wFvsaUC4Tlz7ZVl+Xxi1QFTrAiJF9iwVpoGNVEUK8XE2H
yrp0wgwO14sltjouBID5yMwjlhS1t0FdMd7A8ZYHmQwhSYmTI17XSAdvBPym2Mjy
dVofFho+PIq0KKrSWS2IhIGShYVe0eH8pNK7ZhyG6f/ngScyU+02So8mjwDMXKSZ
wd5rPP9j2vy7uStec1/ic8sFpXE2bWPWr0E74dyC9YmiNH/rO7YkKwUlQ4Vo1mmX
hCUm8lTrhhTGqZDZZfBtfeEZYI/HZXVJ2osNUzvOO21GDvKTzGj9zCPAU9AqrdYW
wvVxP4hqRd0+HnBb890WX4V3NlVSfMzm2YZd1q0mRJo3dosYd+XaVzuVr+oFwjCi
hzm44gJlnaxQNeDFEcqm2z+CqBjDTWlXNfrIoPLiafGoN7CjhS8qqVa3ij9HAZ0I
zIvR2tUtlQhH0HJDH3L0GD+zhU+hcnYcKl4UHHiSpA3itVLpTR/zriteOjEYa/Ma
lS6jUXUZS3klySDdurzpPPNt/a5pY535YA1uJQqbSR06JKUNkuZWJ/DNGTETwrpF
31N8oUrQwRRrtkDPd0jb2OGb1VIvMtkMTwyg8iWIsAJe/klPdVOnZOs4zk0OTP7P
Rof4SToH8ZcFR2l+QCPJK5AxsuGNlga9ORo5aV5jdBrnrfbiNvVqAR4aGvp8wfkI
cnwVYwEH3rSvxdKXqBlLSAIHjBkZ5C8w2bL2auMqzlvkLendXbC2BoxTvGDUKDy+
uapDPHZo8gX2b1y/utV/dg0DgfZ+ojlof0dLK4oUJtwbMS0Zc0b7vZ9WXlL7hqP+
cc+c8ZXWe7XqEPTnpSxXvoRx5xCR37/F/BOTMtU6mlRoy8t5eUGjniHZJrQxf13E
bYGNrrlE/iceFtQQNiM+sAGRWrPee8DMcPLI1Fal1f5WQPNka5pfqZxtSNtl7dmQ
9UPQeRQ3w4RXNgKF2N2I/XV503SppFNmU6xUcsZHIOk6nVw3MyBcTXbHtNTHZmxU
hVuDutQttEwm0epWNS/6GvFFRObzCP9eV+XbjtlmG6jHGHTXtxq/MAWQi0nOKMLG
b/Vf9DIk4IbkeNpMXQQceD2m6n4EzsXe9uMPgz6B2eNJu/KlfcxGzQgvLv/Sfvgr
gj3xuhryj3/JinmP8ntl1iUdGAZvct+2HUXUkuZrPvWQCPd/+2YzrKTqKrLNtrOo
ILtvw3bjZPq8VaruOAD8ozQtOR0unnQLu1gAUYFMUfqEXsUxE0WHVDsNPC774noO
eHONWwF14YPevgVQFc+X9Ud7OM7HSCKN72H4TmCIWRtXN2KER2+e3UXLoYELKGt9
KIIYOhn9z/NSNe48weMckEyU2VF+I2otECO0hE5+hlYOj4GHPS3/t93U2sDXrsG3
LBKqdvp8fzNl8DRRmiAkmpTzpN9a1m5Tph6E5DwaUDnWUTsTtMid4dV7aZdTlOad
NftHgl8fE8i4aUsaO1IM1U05YQbVD+Hj08hVXfmDRLSND/JMKd7krFN2BfsL9pr7
qLKdWoRAELYslen5OXb44f5EOAzg4c51lbl1rLG2hyxrGbvhQaAjWWQmfr7NFXVh
E9lC3YdpzR0jZCaBEnHSVGjJtfYKdBsJF4G+GK0iYkn6dC1kjPsB94UGCviFdtaC
MJp8QlHu6E/dNTRsYB0NxFYa+BqEBB7lw86ju2Q2GQt7kjN5BOv0xIQeuyuC1T5Y
3lUXuRnI7Mviy+ofiyBL3w7scbnDwMvAQSFGG21WadBNMVB3rpO0up+2UhqlXtmq
SNcEhSrq/OTxJq3NEqrYr0XW9DzdEF75/sJFpreISRV69yR4YqQmJTQCAna1MuhX
ZAKTi5Eo76WVE4VxSR6rXnBRSFfYfnROMFICW8tUQLw449+T6HSkMXb7aou9XvQQ
giO07jDtcbcqO3hWYAJPB3ujaq0Nnqo1lfs1MSpO1mQdsK/ATJON3LcPwlvG6AGI
/ojZ+LhSQmrk/8lXvJdJyYWICX6CPoOl/c16cFeFLvEDc0ZJd1FE42QxxL7Qlf5O
jp8LQd07jEzrAl3TApeHdh5uXoWqwbver4/A7jtP7ULWq8J/pUr4Fz8JLd6zwA33
l/R8KnE6MGgjrXw46L+722YZ3HuCBw4ZWMk7N5hkk2LLo4CsgFX1uNemqyKwGEXg
aVrdEErpRUkGcNwRby7zM5RoPB0z9VDdRwUHnt/yr3/9a8E1pWHRWtkBYJquZjoW
nS2aE22CtUQnru/B30TX5f3L0njskQBcdZ478fDeWGvJjE96umxrglozpjwdtJYY
lor6cmb812t5qc2vUV9yc0Ccpx31yPwokIZpHwS1WCICTRDu0Eio0KSSaZ+lI+Zo
pTtQXplQydPbzyjPr54tsOb8NdEu7Lg73nTazn1he56W+khw3lr/aNSvgLXKmGCv
g93CVvZSHx3/KXhft2rZHA55NCUWYlYY5uoxJS1elw+sM67nLme7nd60Ltj8/IlJ
zul+BWFjRfZDBOggwdxXovy07joB0IplAyfUZWmpxQqpeJiVdO9TZE7pS4Ii1msE
w/ypNsiTqJpYXPHBvdTqLTG7tsOTE+cx/3TV4aXiGbBhKHlq+Cryp/9EQAVkP6Vq
e+tnB9nTaWXJjVmA1V4jGzTZA84C8bt/dXbWytJhX40ZPgzL936/et9idYlgJebN
aS2g2tRCaMOfVruqIhcA6yGpRRKWgZOSSjgIwLR/2eEfpRoqfS28duSePMjS/FrA
qkovqE3SQUU1eXAo+NGiD2N8o43xueFjmWQ1Pg7e6P64ZV7D0zyTk16djHN9DVS7
yxZADWESIo/A7DydQToI1xTlWe3xm3JAFscj/U0eYNUd6fADS/GMUVS5PtB43WwQ
gPboc1iqCymzveb69GB3ZKk1901IVtDILlMeTesnW+a2dQv95KeL6RaYaUagBNmz
Egskj/oEJTtdTED890rdWkoehueiucPcqRn+nQ4am+i+i25XQY4srWTn0klmwVKF
gKoEI/dB7ZkiUBDeemUGD8YTvxw3xvataVPBJGshviCqwZ64m/UXK3VFyrKTDcIP
bt/7gYG6BtF0am3Gb8Aqi5GBK97Ujx07KeT82PGyA0oJNFAaD+V5W2w0L8OXZAP0
HOy/zE6OX7CAaKOegSNiyHed1AaJtXgQHA9ZoAll6ZF3NKoM3342sOZmTo5S0n6m
eBytK17jDDUpuGrJO66/zoV6iXaQri/oUtTW+xeMmN3xwJbYG9Cdj2Lz+Z2GzUky
Vo/XADr71lXewaQK3J2cL7SGuqhnx+S+Yab5YAo4nhyntjryWhcRyWAaB1ZttLi8
5W6513v0sx+Sxjym/7r24whgBWj11a7sbrL/nGcIrj3pRy2UqfuFtphJrKvbftle
EVFokQe7SsFcaT32+0nqBAIJKU3/O5ly4yETgm6W2Zv3dH9WgStpXJABuUxTdbgj
6oHRuUZG1aDTXB+P1iFUbVoBBRF7dSrUWiNels9EmfN9pqFIHrgO2AYI0l2xiucx
p3TPlGmJGYhzWlqv5RQ1IiHDj85kUYYXLW8M4CYzwqoFWXDrYjbqqwWhMFckFJN3
SePLBgEw7kuna4der1H5NhkeDnNmmid4RwUBp4Wd29XNRw9nz7gOAVVfOVBl5D9j
XBLXFL5GkNjjQOHikXxhTfJt1KOrcks7HYlHzobKwWmrKOAVq2Oyjcdz7VdlDvZz
A9CDnsd7DWEp2BEUJlakBKoA3xcqhEA4dc7VcfFLvzlqkh7xIx76na0brOVR3vsJ
SQwYtlRkYtwo5jKTuY7HGEZlCgfrf54/rElPgdJU9Jqhj9k4T5whTWk+7+OZVyZp
yFpycQFpZiKCSjk/zy6M5azJCSZfsWkZfnBIY5YuyqJPQkrGUGLwmqCQJ1PMf11k
dqSg/kGpelJQ64Y4v9NMb4zopT6m6RGgropkFPaKjcjv1smvabTBsbTfhJZ+Rtkj
y1WMR4E5LLsMyAuDKIyqthrectDz1sU6C9yiTMXgmOfBzXYczPIAsPGq61Ir6uti
Q2bXMhaNTAMAoahLqigJqCtamT2fsjDLfGevVyE4r09bUtfPJCtRWb0jvI5f2NCl
wDiYzNP3hV5KFNd5KQ44eTZiIa9RfIKEOND0McRQ6IjbUchGooMkTbzr5JcDPjTM
Lj0DZUUJKOGwPDeD03qhPpQaCWwdOazvw+LzETofV1VoS9envR1FWnX2Z+eNHb40
k1V91bgcVl3TzrYkncfWSILi4frkUdBpzTwrltRZuECi3WZa7ftEmZM40wKseeuY
HJkkZJHWG4EU+Xs4X3sruyCvGSXJ3tDP5U77bBqHo0sMpZd7doC7lXrEMSRjEzXN
RABHBkX2vPxBXID+bQ5qJBt5sPWtTUjvRQQfcKlxuCJsxRVjw2HBLgEZpzz0NNE1
u06AuAOw8wYrtzXMuzXelY0p5bsC7lkgKsBzety5HFIdvNsCPHvQxK6We8fZUqpL
ImY7uLEHnXOmnGTFg7LoUDZ2NzvR7BWXtMFsZtKc07na2hwAR30PDz6vxzNCReKJ
89uwQ5FAy5/rnrld2d48EgUKeFlVvpc6mT+XjaeLuBiB4RECcym73H3zSr5rOzoQ
agC7JLbXYxDjt6AJ9C3CPrNsABUI9jXnCUOW7Kn6ywvTsuO8Fo7kzQpSLs0d4iz6
bQg0oZd6SFC8H3+7Bw6OuBOz3oyaeHgHdjj8ZnHymieULt8P+jNjEwl4H/zeGmhh
arwzQOQ1BOuhADu1gVT88njwQhs2HHcwMhnx/QC4t4znl5JIcf+vD13nclrFVyZu
tnsocx00Zla42WY/fGL4xOmhoJB0O9DVPAB8KKd60pZgyaDeMy6SH42KjpddDEK0
PySmtBUEUHlibsKb3DOm0+Pa5YbnbBJkGyHI5RK/dcmz7Ron8v9NNt6LS6ad/QA6
oF9u8s+hm1b0GQ2yRlCC4PD0OEgVh7ULK3slOh5SWkQSHvaVzPKxyS6hDpHWrOGB
H9l66IVtCA49cR6fr6RqAtq+a5JxNUyc6a0eEH08SvBAD2TdYg+hAHABiULZs171
jl+kNzrmWdO8pBJ3WI+E9o5XeiA+OYlTApHjzONdxC/ePwJmhr+7vXKcuWxMkfvR
1YjTCrBkpyIIym9mfEgZffDbJ2tVsn6xpM7hFYVIQJaY2nLV8YHNWB3lIE/PUUQQ
6n7oMznybS88dIFSGd6XdTPTjU+on485SpLUkvnZMkk6OaK3RSz9jhm0ucWPmzmt
8SOhee0m/wApI8KDORm3Qvra53mc861pBbHgurGtizFQ8qhxk16VZs9mAlMkGQuZ
+xdNQlaroPN3WTHSEspDfjisr3bqEeRqkM95ImLuS5zM0DLa8aDnwH7RRPjs7QJW
TIDXqFmQ2YBqkqM1ATqs1k9X/9IrF77RhD7IoJ9U6w3Guq6BTF6rc808YUi9Rc7C
Pe1Y6l3o9c5I30O8YtbSFm4K4qApPy7Potexd1RotXs8p9+P6ZLbNZhGKgARjtwC
YFfIlorMRTtYBwMnsdnn0/MQcLJLo+atFwf8iTP0Po9J/EKYOJ6wJHrs3gW/ufWA
ZkE8qiwomtlE0NyrtcEdJbJ9KMFOSVwtNF8m7xYN3m8yeZrI3dPBOwwVMnUfPIvS
USA2gyS4nTg8XF9dR7od9YjD9BtTXzjhCsz7z9d7U9SLNvh76MVc6eAR/hSBrl9q
yX0ev9K2Pb5KtHnqM8rD/cheJbXHXZUPUXufQQjZwcyWJ8KuMwMdi+L43f7e50h/
tjIN1EFgbL6eaHddKOh3gC6BCqdtdpgqwo1jskrhhAG/KcLgNU/wZjSVKxtZZfCx
bKjiz0Y9XZRdFeaWlzsF2J2Gfw+G7rflOG/WORHtLBMj+69CEh71x409z5Essyh9
2klLKee+9vTHU8IEik9etWWVL3zURUwwvbH6PEZHDUg=
//pragma protect end_data_block
//pragma protect digest_block
CWROFSpUw+PoFcIhIG1EL7WHmNY=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3l20QKImxLXceg9pMxuQxzgBCc3Nc8HRJr+SrYUWrPkn+yUQiokSPOHjPc9XElKk
aFUxs64Qe+gazS3Jz5xb44ffGGtEJNtd4osiwa/Er554HrtLTAwSr32ZBnvkE1UP
/fHwe4N8eViW0iL3Nggyb5s+nxC125lesgAZJfne7t8hXcjXAm4Sfg==
//pragma protect end_key_block
//pragma protect digest_block
cP/AhZ+Q7f12do6ShIcrmqwDAEA=
//pragma protect end_digest_block
//pragma protect data_block
ZPKfcfXWWfQu7NvfERF2VPMyS+SJYgiK8SG4tLmChNze1i9qrVTqJMGP5A98mbbH
w+F9L+EtMskth2FhcGLHX8X8UFSFDAMyrjtgReAityRkeyFJfS7kaF5Oxci/gEK0
yW5ib7KbnYxEnSwK/tnvZSfPkR9A32awDuiM4w49EFn3qbE5vLRRAMdN9M76wahh
hIFPuNffBZdHRxNuvpdM0fRiqozXt9D85Q0OgadcwZq+zIv78W51W2ttJuIM6LIQ
OM+uTOS30RSwqhy9nIfT9ndpCqr+wtg0mpVIsJlEaMm/V1K+sWS8wrnuaZ+XaBVp
ArP3MjDCG08GcfYFwgx9uDVyLxm3i/iSmZ7+WTmCfBwmgDztAekiVTFOh5hudlMP
Cif56SFz5GK+BeFizkGE2w==
//pragma protect end_data_block
//pragma protect digest_block
wub6QJVd/SuUuo6DMO606XFp4oA=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
zlmOqcLu6K8i/CTXh/RZC6fyFiHqrEPtiWSunHYJjivwX4jbLq2kXFcjqyplQKQA
PMNk7INC4PxEHFdei2l5jgM09UmkbVj/JhkL8HfYkx2B985iIWzbls6hKKk2/4ur
QOi5Tq/+cAx77Zfr15DbzicHc7C4UA36yZedLYEm+FnjPLIpGt44oA==
//pragma protect end_key_block
//pragma protect digest_block
68QU4PKHixS2D83zp1u/mfyggOQ=
//pragma protect end_digest_block
//pragma protect data_block
ubH/WbPaOYKyEwsz/14WLosKby2sChSemeoqsCnFFaRIjJjOj+xeFEHGCT8KuHYR
E3duJQK4BOcLtqOy7XpGao4CbhoaRU7+/qtgfRcRoETVyOMwUqD1SYPPra+4J+lH
WDvlS+DpDPTfdQxoAB8s1R1dnK5PdBVYt/k2HQUovgrniRlqw+j8qFHiBXrzzytp
WK4uTkZ+3UDC4DRq2oRT7jGuCv5inPcU2Az2eQrlivgnKoBVnmE0AtOo7N2/y6Gb
xdpLscuUWW1QM8ZmXyew5NloWrvXVZnuF87PkspQO9IonZLDf0oAdxm6N3AmKksb
v+m8KSslR9hT/LFmNLOFm9bQIiTod8+82NYAGv2OevwrWC9Q8YidmSP2SIwgv3JH
Nft17HFsA9UH2L6wy64POQJ4f8O3OW1XAKBxdHQTASnEy9S1bUZa7pvpc5HJg1MF
IE2CCRKC8kg7UzUXSoUOgywYA+srsLW1Ellhlmez1DCsh35i98VbEXstLmDk/Dt+
VvUD9iCMAgDoFHg/xvSV2PSFUs9hSfSmT16p2w4gKfEEMIeg1XCHt4xT9xRyKECV
mzx5G0OIhjqMgY/YQR5qb10cNcSMudUlT84juTOLPfpo8VJLVh/qYcVTNoFy2EXZ
0x8XJOY1KUQnkvgfi0BJpJx3taeppzvgeMcAl077sagxoUn0YGmopdPMhw2Gfedz
dUf+2GHMU6CSUooBrAyHxUmcw4st9JiDDiYS9TxtRzl9ovWt6KPO6lqaIhGe2qVX
t4vOaDWy2S2XTUANL4/xouUBbYLtW1uH7WVQUhouWvMYCX2P/DA5o9diCNuzh5te
TnSkLMbJwhsCmEa1XeCE7UBn7QrZKpGP5GZRolbIByzcEHKWSELa86eee3W3sP+w
Dw5D4pNrW5EPGqUmmSpy5sTFj4KhSaD1KKnPwblsoOAtKTimcXdcRlzyODiiUbHD
4dAb6TAIknsJrZs+z6NAo1Loh8Ycn3a+JwAZF5mEFkZnNasdIcdBKGLO2SIunHtc
SCxj05OYNPnBuMOlR+uMwsuIQ55102V7kExu6Ey1KLXe3ofmuJ5ZLxhXvJaQ1BDa
z0EffZ/X0v/pyZouKLKMlErzY2pynlhkXmtyBGU3qQDB9+azA2w8c1oJ3lIjHULR
PX7/luAUO+MBy7007gkyl3EOcWABpOhCQc4uKLuVzkOp8YfKpkwTxIovcjKVVPr2
8fXuoqrRvSojTwVJdK6VCepnnNTvw7etrXTInxkMv1M12DTf+sB2J4jSifVXSfg3
97wyCcgNdpAFjClHcYKqVQKDGU1mr4SaHuQ+0cXooToTDZJC5NYOUAHdvDADRYhB
lWEZpjLid2yGjqEw7wSRySEyWhAg+s901PyEBZF4uhAaz11Ohj8iZgvxcYfF8GzA
SuApiiCyj+i4lTDbVnF5Ngq0r7PwCG9PdPGBHIXwJFc0+UC1t5OchZ/OH4brJQjJ
mxRe/hYNFbPqdnQ0DvKqkZRgCAntJvkchtZ+RhXsq9OOdCzQoIY1I+ZoJnhQEXnY
sHFO65Es+WCgSHbO7I2bf14SHdkTVXPmfRuKvadgmgd7v2K2EZcI0RoUX/s9oinf
tLGZLdknjR2iH3wsi069bCDdJSPkN58EM/cnILy1Hf7cc684UhCQhPY7ipK1nOfZ
QNO6U349iQWV4Jl1i25+6KCgDlxCKGrKPVSyrHTgjwclB5x3BQkYmTY+5T8vKiQv
+kpISDfFCXvcMJPRGnpqi5LH4gxlE8ajPvGkdceFe26SJIYsdWT7azFk52Rhi1S+
CjKHjwf96A1TU0cPKSSCDbhfeAvcUUIVv3eYiz++r1RYzO9cU11iOEUFKGx6pA9P
y0ITUp9UccJl/tb8M1m6YN1KxEq1rpBJOwNZEvHEeCdMYFm6QLDoWiXTttVtMCLx
oUIn8kpmRkz7W5lKUUhMQVup225UVjScmmV6HzA/1Ar0rh8agIK3PClUM3I1S5vr
YP69HZSnHnHJ2csAcJFK/NleIGmxZHcHHvMheKdOW3PXo6PbyjKrMDOCVx2x6DyH
cKDzvyaq4j652xIn+OtCRRiMWsJ6riMBTwKEEW2Rj1IpgRg2m60GfZhbcxHfR7XV
HTkP6uwmojbobjQSRU3lu6fBV7jlqqiqhVrb21OEJDja9ded1qWgoVMqTJuGKUlF
vbKt04L0WKJG1ceNvAnTlcIreuk/b7pBej41qtvyLGJgoSPGhM6H2zYT20/GjE7a
Eb0jj1kbIuH3FsgibQvYYKyu9rRl24VODcQmQtKHRcQzry0tGgZqP7H/tYlT+jM5
WdX6ipuQ87yOW6wpq2hBLap4YyfAWE6iM5OU+KNC7D9nnxIIKsjnxGJNuGxG2kDO
VCbIBaLAeNqHk/6g/JbuebBNfIRa27Z3NLaJnjcS3xHPgXqFQcybMQuvfUMywJ31
NmIhCiT4kdo49Zt6awDXf9lKk+KhiAnzA+fsaM67uUm3+8awjN2TjrAwuUJpsy/S
c7bNLsjFNxVTqRj3+yAM4nz6iX+RWP+8dM2npRx+Xnw0kHeYNVSn1sOChNFQSvPZ
WD9fcqPv/paEMJAMYoAhuzX/6BsAtjel9LLBrqz0a2sgMXUWf6GKKM2xdDPFL1Zw
7EROelNLVwd06oBjfyLB4FsudyJQl7C9gNUggwJAST/pnz1lnhVzvEXeBBeUCpK4
M/gx+c0IyUu2xJunqxiebQ88d50AuLHF+pUXcYdCF1CvxLFXSYNk3H9gMnsYD5lJ
fnURcGE8f5qn1DPDvwVaptO5f/YKNAq/Q2LNvBqT2n4rWoUBPuWJ5v4YmE/++k8A
HUjeKmjMtn1aFehSrtigrEft91O6kulORtjDlyxRjV1QTJUIL0tDCaXzHHAsJqyg
PBtWYmPuMJtjO8+duW1rVXSHDxJuPTnKpB2LicfHIXc70+HPFX4auIAVMIJrwPU+
Y7kQkfiPUHPvrb/hWNQzQ1vSqbOY4ADoctI+C1PZiq8vMc3g9VjALRLK7af64E25
sHYaVgjX4/pjKUrnM9GM1VTRCP0jKUUlLckMJcMBHiwqP2S5y+gb7nR/LcZ0h7vG
dG+9N6s8FZLEPR7pFu+9Ivarzo9r9Gnc8YDOlGyoleZBdrHGQJNaKSBZPkxCg4Oa
N9zCNKA3iV8xDrhbQJesSWZFBX1Gx7TZN/IZDYfQfWzsXz3NOMjmab69vOxIusfQ
VkCKXvFOQakCnjwJoKXeWNLzumwiAXEOZbneWUHPHV6h+hIBlViKF1HpWJtwBoET
ojvMYnru0QlOrwSi5nmT/vq61CRa2etjGhHf1w4Panq5oDUDMHVLnx93HNWul3F6
DSTOyo2+1aJoxn4U3R8B+IQhcksSrUNJtFWQUBHxGkXvph3fmGMCQyr6yFZwx+jt
RwbmJUaaRr7l3BCQ0Y1xhyI9gw4FU35LyW+1gOp7Cfu5Q8uAiJV+Eu4R7hGVM4Nr
kuM+ADQIAbjruvbcTVB/hraPkLhVrQgXjN9ckTzVIUaWCqm/ipmQ6r2K3KAjIH3S
k0jYp3lVx6H+daKRJiGYqyXFdmnOdtueSubet2buHXZFKjriuS0Avt0F+L0oCQf/
09G5F9Nvqamocto4MqthVSVVbe3rruuEd6zh9Gw1xxfbcHEKSNiWrFrHbdOabL2r
ryZHELL9moyorvNWCrYUXrT8oBbb+YIR0Eewb0D1S+3XgvMUB5shJbQCEFse11IP
ru67WGhTsGDxwEkM7B6xTB9ZWxLJMxFw25jK2BhILt7/oy/AXfqUY3C4xx8VFqoH
ojiBVz8+nTNALcBLqtsrILeFDBZuvJkxSOpp0UCX94N//ih34Oj4Xn3SYs86qWbe
N6WWh/Z2Lgfjj64PO2yITXjry91sWra3UORZsTKwWwKTd5TmgxA2s4WG53MnwCQQ
B0NT279e3POuNUAopvpm6/RMbQQYge/kW6tynS+YwThcg7ACElOtAyt1gbwMqBWf
tkqfKNF9BQviQc5ziFDMj8BhQYpXxlS2mqvo9WXXKTFglRA9vdjhffl53Z29/Apm
ed9+OnJuVTg5jHEHdfqHNvUroosgAg3sUhw+RAtPt2rHhYYsjiPASBczkpwdhwyR
k4bZeX6oBBng5UiroTIkDSJ79Pq3QybBc5RCX1ttN02D4wSIJipBwZNYNuK5fMTD
cUljDXT4H94GLPIxEOBaOUQ2Ea7e8/X9nYIjx9o8BEt8TGQTB5IvenqdhFBM4lCs
0dQUnv3RIDGgdBTze1Tg3aoXc2qYSOr5oUa2PayeztGb8Rc8IMg4TSoBIHLfErr7
4c7rN7wGnT0ZaEx51gYQyapyYGGy9gnn8/fKibInxbFNQc95n4bPL7SuomFoNSe7
heO8XGmacKZmklqC7dSsZrk3ImIQVa6cy6Oh9zAV44igu6kQR+cmFLVC5iNe9uOR
b8NphbgfK/v791sKfw+14oTJk3n7NWMG0ZKewi5c5OhYcLRRh8B5if17nkpskLKx
JCovuTCmCLjmY04eKEg0vFX3L/bi1/JA06bPgJnJ/5DwwhyxGU2G+H9CFrDVFejV
kXe0aj4NBvbckn59rby57gJJbkKUu2/wBoTN0Xd76MJznVhgY1snxDRW9Mu+niPe
8/u3vIkymRupnnt/zjB+VaSgkzB92Hd8VNvW3Q1tATTxdqCSWfJHHOTCDhx+qjv6
bB3P2W9b3fr9lBuD1NAbFRGp20V3ioLQ1FW5Pn5THyQC3UkbcoED+/+urlapz12a
VR4xAzlYhs4BNF5owp9vkL2nTbH0UZIcpeiNNOYh3cVToZZpR/5vvvlYcoGaGIWc
YrTljd/et/EYvzlhrIkLTmqcy9G0kJJG7Bwt8IVBqFvUZ29ycEjOGOqG5UprR8Cq
D0QH3Zl+O0wBQrDKh+eB0KPKNeXtVlHqhnHvHgiCb1GLxLrGcaibdg0Dq/ZKXCl4
Rb18ja9AcuaQs6IAErYh6lPh1SthVlBaEQUjJInBm4yLA2ghb0pwtUDGGbsiZo3h
+zX2FqXHd46dJ5pnJaV3vs3X+8yP4qip7TxNZpJA1ExmjrIsy6Sje6CSvNSiHwuL
1G0W9nQIdIicU0Uf3FCMgBVcCtfPd2O+H5sSsUF9XpWHErNqUtGfjeWhs2qMdwjt
4n4WvsRqGiUssic+hR8Ggx+YUD7/38eoqaTBaD2P51e2TPTIUT1qEXYAKxpLgtfG
yBrO43fRXzqqcWBaSGNSjxQO9fuVoAtN+VCxzQ5bo6RAuxCtuzR09JZvlysKogHP
RFjV67L0UezmyCJiVCOQHUbqBQ6KT9NsqgLFxw08N7zjxAaEJr+vuvU75mELfz1G
6xcKzX67NZGSN4H5hOnXoH4StYJS3yBJ204AqWe0Tmb7+ZTge4eB9R6W4FMDeVqT
+pzSTpCce+LvHO793ouL8hCjn8GGT4pGnb+hthGhCCaNWVLvON84AH+kiaQ7z4zS
23TIxgo3fOeLL3kf2BfiXV6r3WAT4Vf1LDoCudlmX5xozEpkKiZi9dIyinXOq/5p
1lo72KVVQI1srReF9BzEg0QyJDr7RIoRpj/+8pFoqNKt0QY161Ix+NWyRHBAoEVl
3Bya/InRP2HjjiPQ7jZSO4qBtY26xYqUNgD+UdqqfBFr6Y/Qydl9y3N5bsReM8g+
bq3yHbCm4NBU6bchSSGMg4Cp+bGyyg7EzZc/6+uMbWg52fuKuPXQ0ViZKihxnVXX
Yt2wsAGnroQ9I7M7mtA9M6Ns7GBWEdKa9i7ElDQdNk3dXlL55ikjF310Iho9WBpT
K8H+Dr1wFs0g/unTHEWMK1w/B0GeNNNgAuh0YsVnUlBAuNKDq5TNBnzsa2oItgeL
DBfFUAhoXVTVQiZ341dkIPNx+PaySyEcZUFpaO/X+htoolcQym5qwtAwlkjrADWv
xldH6PLbedlB1sU6dSvKzBdSACsQO255lfTZhPoqEIIXLOQBft9Ib/2e26O3VDML
zDV+FRp7dA41hssmhxE+0QDna36siVV+Yv2uX/F6ik3hRv3Le2SnmXj+V2Xjvig9
h+UR3IjkVdGpAkpF/LA9KjnuX9Pt71Xy49wp/aDLTEB54zVAZP3JJ8jHKxZs2mTo
MW11VRSgK4s4VluS3Ym6s9pJotc8DimKF0dDKgDM8CnO8PqdJN46qnLeqkRhYvi4
vFgeQYr+1VkDTgC5bGGvxrGiczmcb2BpS4TCAY5+hsxhdqhoQtJbbNV++M6erm4x
VVXytdQR1oc/E1ssbQ2MwYdocsJOuQ2D4TNkQT5f2SbQ1sqbHs2R+dnMFwauDVU1
5TnqXpWxHufFdn5dZqFJ7T23hh/8C55QbQ9sCcMwOmsGn63DX/qCnS3RzYr+5oPR
ltebX71u2DO3M8NT9iNsZ9TuHM6C4CaUNtMdUSbk712EHvqLfNxw4UGfD2o53joU
1pxsPJMiqvHWK3zoC9CIqTPK4JH2KutyYabhX65Lp0vm2rkpF6bSRP6rYJjSx+tD
cgoCvxVCknzgd/KwRU6hVgKiEBwoyqnvdLlwPIkWEg7PO1m7VibPyUN86CpLq2Tb
50DWTMp6LsBv3ENTeaalHB8ieIALNjp8KZTS3S0H9CJdGDVuYTEomNX28kWMtOMj
d7jVZoPyxGzz+ZVCOVfoIR0NT0EFttZzT2qPN5373+gVh+34RQhsLAM0YKPe6fXs
nCZ5jgjZzNbLhQsJQBWkI1U2lk40BJsm/nGyp54sEr5FyjErmV7JNaMm7ZkyNBNg
XEhzTFtElzdedg38IjwZJECxjtR2Gehp1JE1l2jBCpAjwdgaceRoM7jB2Xd2gZpj
3YA8NsTVU7AHuUTpxtTyoigpB9Hl6gYKPq7sOJ36NgCAbocockzSqisrLmBdg8wk
Hza2M7AGh8j28jZGw+NmkZfXG6vOzbq8A6FtKY23QPvDeKVR2kJbAQ0d1rdsM8gR
oasvHhpW/r7oEj+HsapXyN5V6/cxdi2XF4JVIPYFLELAG4D1ck6PpNoCpXtm9MGt
NjceQLeYltKbE2jhBFpW2TX2zQFvGswcvK25Q2Ko5fVY35Z3DdotkWJZg/qhNOwm
l48M5wRyvyJi1dk5eEipPflGA2nbkICGGNaoymdexUtkT6wxXnR32cp2AQNOc41v
gnygeNfPUXuyfCiKJ5e7l0kXyriAfx3T7eIBhMYVt8FUS0RkBRgQRvGwDY2pMmZa
GxDlh4y7S+DoJJKbPpdJ+LwTBEvaVjc+PKHjSmpYrzG2cKb8TbwlOBxbFxESTC/y
JFno6+AufwEjTXqwVgrVJVj57ppKhCWvGWeLWDqb6SMV7+lJpFY5v/zafn84ywAA
2lEt5IRLiW8mmc7CwngnkDFBHSW4XZ36O4CS3xhkY0qmI+VOwrGS/8qQSdWs/V+P
vM5hGYdPljqk4PqZtJQiLsY0qL4foDz6bfo6OIVI/662W+LRqnbsYAidJ41NRfKG
xgDmfpHAwIsH4QEy2wZKH+b4WsYCqMxXv7yEYyQ+2hEWWNEry2BoXGCYAecy7sDl
/ja6/nOf/8t2BsbJNY6gczqmKAOxKHNcJjTbUOL7ZpWxPm1r33uZehBiqN2OFd8V
H+JpIcYkpr1uFzXAfCwOknBXafzV7V29ftF8kjLM6EM2KdMzyhkPChIudoH+YeLz
4GW7HojE15omaN+n7xEzCzDQUamyfYD94NMNrBoUEPRpH8UvwaPVTpGiYNGixc7T
AJWGflgB8Mh1kUE+Vyurws7cfYQGAbxS68RnZRY+LLNANm8r9XDFlZvH5TNJxKbI
avkD98i+ayjIkx6PiQJmsBd7Lkn+4Fl0jtSJ0+NWnuVR/5v1EVOPNe10Xvz9sB9o
eV5MWJ3/60iYIG3Nz4Ne4m9/bgealr+cVV6dW0Yx9lnFsc2sSPBPA1TfC74WrLsC
X8LTDfwFnMhtrZjmJkbCTfMcMA4lKIQND+a5+WYkNvYp8gk/8kOJ5ocNJWZzrpJ1
MVYgsfpR6s0Q8+pxwQ70tRmbSMzONu5xxLjNnDMIIM9MdxrzDrvEg0hnkPc5wVrb
Pj28DS73pulFP/ynbDXvAN6TFE/yt0F90ZrYbq/BWVyoOm1qCecIN9zmLWTDF9Zp
HwcRD1r0kISXl0MDh+AUFEkV4W9+OAM2VRithgjNDun3JjSp1EEBV63Nu8Q3JP6a
obHLL3T62Prodo7Rmj1f/n5p9M48xevzaGbpTH6Y0eNJnZvaatzsGV7XLjYv34MV
4GEAB9xwGEyrXJvG7G1WV9eQpWqVR23cc1T3velxfkuNuvz+ZrKeMy71t2yoa1p1
FxuB4HNxgefdU6cLhAr0eLAyfrN2HW1vd+7SYGVpkYxT4nO3UKpXRm4yUKPTjfWB
f7BPpyUO+U+XGNaoroG3J1QwKqmbSHtPvdRAGFUADAnAN4JgFJn4OBSfAAp4Lyys
157xWqDJV0qNf+WO0ZoQUmty9bOlFkNOUE2uELMcD8WGBkhBB3uukG4pHOmgV8QV
jVHTCG+M005yjUae5VvsKf+6jbUHE/cgMHf5uYhdq7+NnkPuynL6t2SjFpExp392
X1zTogxEM865nWnCuxU6oOsrBuBenzvwJ+GPCaEHolotyYEgwnsPbmoYpSAYD8Mn
IYBkYq6ll1QSfSyQlSkL/KCtg03+i8tePsRPiSDgv0Y4Yq17THJX6I+d/2wlrZ8c
MOs7+flOPmZQXYcCrB0Bs1SPoYLH2qxDk5ghSR8MOLVh4FTEFkSTIhiz/dTEvWvp
Pypt8EixED5aO+GZkmjAzYnYjwPGMS+FR2OV59t0/R5Seg0RrYiloKsAb6VhHsGs
sXq0uXzjaP8wNAlhB0Z7oOCGkGwAcbXju3KmkCLUbrLp3YKEj+osqLt3KaHhtsJr
6BiYxioGMwW66fQehzsjLfAaSmUxgf/Frl9BPLshA2mQh4JbiuBQMszJg2Yv4iCH
2ZRmMdfZbsuEJYc8AeqftMoX/aDTZV1zhQxOwir9ChIycfoh1zCFjkrmWzfGBHGQ
V8xb93L6LEoRTA/3T+K6NUrhmm/Phf9d+4lqLBXA6AdemjRZcHoDgQWX1vfhJegd
KlLHTE8otJdz5fgIWCCmz+yj3a37z9ltHHVfSPC88bDr0yO9AYorfRA78stFqQWO
UqXNGsqGLm0SSehKx5nNYfgbWITjTJpWOv1vBb5d8xYgDyoyYO5KIWSZHim7LsiW
7ALDBa6WsBib4FW1dfTmFnqpuOh+bAgVn53YF/Su/Ev8+jVFhC54KCJHwdUqvN9i
jwDEH83SjE2LszMRfTaOSYn59uCod5jU0vvsXYksNfINdNi3XeAr224mJNXcz0Yh
8wHyjxlM5gjmqSmZpPBXneoDZMWudM3F8pNY6UNerbXAoObyYxUS2xK1EVSVgI+r
ahc4usmK3EdOc9H3xJbuYYF9iV4MBUPj8OwLlYsWE/TpeNVAwVpjDhFbzMpXQo9j
UVF8Lm8MWPDY85EsY5NuvE61tbSFUPMvIq1aOioZ6DF/VkqtxfZgedompDKXD/Nu
ZO8SzE6QlL7TencCN266rBIGGdyUtcoR1MUTLyRJWuo7MDrPhYavrYG/qI02ceDQ
jJFrhXVZUh28zcp2L6NqTTwxIDQlGuF8TuB3YITWhOl1vias3O0cDm2ndunwldvM
Kq5YDYDkDjVYo1dMxFWoLJzm0zXW7wCStzBfAbyorlWikCzuKivjgo8XINE4CLzD
EwrNxgT+IqS0+RsC6HtFhsWywex4gs6UhMIXAlYZVZ9BJb01Xurv4c2ZdmLg2yXx
1ZkiMyMDqS1i3rfskTWp/8rJ5ZwXKcLyMwrfEeNfaWZVDMaM5bCAZYIsc5EKmeYs
pAHaT3i4GVoDgQ897CrVdL7xZw9u4TXK+1meZtjOnW0zf0kvm0RQd8top+ZgCe/4
8lU8b2xY6HIgAjBtGXUZ4wcfs2izuLHTJpIP4yddkIHPillueh63fQqDcmiz7kcZ
aZ5kP0xBcy3QJfjB4oaSRgrT8E2qtZ3QWAe1nbtvG+3Je/ys1/6JiY8RSC0QkfW+
EkbdiLX470TjAJee5wuacjoX0xWScJ4fQljmPX4zg7VaPmLhoCLO5Phjsw3+Ks5l
0kC5pQjNkH2BpMU5MXFHJdLzgud6knXnirYgzyPYuqe52Zec2zW5jqMtlghjWwRf
5YH7kKqTPUTDIiF1Na+IocImhdYMtgTR9ojZZILj4zaSOiuze85kJG/d3wq7p7QX
IumFUoZ3quBY98CSWy+C+gxPzoW+a72/6rH2YEBrP8eKZBDgDMYEZqt4TG+TXqjR
UyjEqCXU5WJ8v1MtflLO7h8WNsrGe8aVZeXYeSrHzRhxMpKmxE5BjDwCiB1D8Gbr
rv7M1i/H0rIi6I07N+d0Xygcyg20aua8gFcZpCUENNhA+F6qtGEatT8tlyIIHlHc
4uSRb7HEFyeXoyL76VVAayjfSt4pKyyMqbXW8d4CKVeb/FLrIThzOQ5NAQDZgcgO
D6x9tV9arg8J4edNCkHso+YvDZK69uZS8h96gitNmgg0L8I/IAQMt92j099xccZx
O+Rz7f8OLBBUbWiQBJTm/u1VdSXd5Sm8VWtGu3pnPkTyNR4tLYzNMks7/6aiFVGv
MJaS02O6F7yXNUrXO33b8e+wTN32N/Kvy/AUit2ONbEw9OC1PiWUthDDEJSpxkQt
hTuctFoMzrwkFKYm9ug8Bme6rzjusqXCxi8Ezf1IG2jgLWTzGCrJapZ5qvU9oU3L
v5+X5nRZ7yR430r2iBv/cxgGi+xuiutYnoDiZS/eAJHuZYr1M+o2NAyENp9DViJG

//pragma protect end_data_block
//pragma protect digest_block
LqyhO1516ye57lhlI9i0bTFqLn4=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Ix01KxkJNpqXloWgZEkEVYaaxFIuczGQjXtV9Ukztkj+p4Q5FDaPIDkESx84fyF4
6YZbnkpC9wWc1cmXCzhGTOCioEAYKbsMuRamx8XIxMPaYprSWocQbPz7BaFKl1+E
uNt0Di+JZYWeR7qRpiLCnJC6VaBZoGNDg1GRRmBnf/jYDUcMtnhV3Q==
//pragma protect end_key_block
//pragma protect digest_block
9GqzfxLjcsXtpC05rIJzZ1tAEOE=
//pragma protect end_digest_block
//pragma protect data_block
r3053Cs8iUGeRFVnqS6PcCR2ux7zVk7UHCS6uNuk23BRt5DlVcicV2ytdo143e0p
n8NnceSZzEvEBrrwSZbKYmT57T6j0pCBCDriEQy4PKNv+qITP8kClvGqB7WdrTxX
Uy6tkumWJv7mZPUhsC/JlflJ8CL4mp5fHtKvFDjJ41+35hTTEraMRdj36rPzL5RC
zvXygVRL21GAmhgUvajs8GaLlbjAdBVL2tgG/KqFFAoCjIKvxJ4mtS54BteStY36
zkeBF4bMvSHaqFr4we8vBA8HD7buqajB/tQ2MVH1sY7C/SJEfR2Y+V/zSJVcXXoD
l/jZClphFrL+pHxxAxiznz6g4q7RTZBiFfUhtSINzqEQSKjY8vg/t0W/Y52zlPTS
Pbd2DpQ2yO7Ephd6YyxMKar+V5drF3BirQGv66i99uSTH/WtR/V2k+84E7PwFGyl
laYgXk0D4BrVH+q5I3rM/4IJQ1XJ6sndAKCayMrGQR1kdFOSsQCDS6vR5I9Nt7Z1
jPsDvnyNrDdn3LAkd9BNpQ7QGJ/+i7NnlOjY9NRaVnJrEFarPOehSVGeIQGrUgWX
qHrGiLVp+QDU5LMDgz3wyL/+TpiOqsvSsGh7+PIyfq2JbDXqoRub69LljLewXtbQ
Pa9F4XPQqiSFjBedl1d5T8doJUolgK4Ot9l31PmSzTc=
//pragma protect end_data_block
//pragma protect digest_block
jubcizW/TERcY2jHUMDVAjB01Pw=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
shDZWKOdjbaip24+QX+S1kWBwXpxW031ZZdpm4vg4lNlWEV3pJnAAXP/wy5bQ8cg
Z2fUO1Jlo8A+VDoAVLHtY55CqUL0dk949eSp6SwlYOcEzju4UBWNfyKUWK5D4ys1
uwW9errqgfUm7pVGUTi2dX5CSo7F7Gs4B6Hy3eu9W1SoTWYwu2N8jw==
//pragma protect end_key_block
//pragma protect digest_block
OKCEqfFjDzSMW0/XEniqcWDTyLg=
//pragma protect end_digest_block
//pragma protect data_block
vtB0xlo+DlhoLridat1vuz1NI3PCck1eTLOcMBQOBZlKecVD/fCcY1J+ECQ9Zxnd
TbrcoSbRA3PODIzQQcYzTggdBphA/6xlHMVke2L3sANpoZgPeChF8TY0d6+fCXCs
53Uef6UPlOvYSCGsTFJqh79P4KFJQ5Cypn7Eae7ddy0LkcsGakXtp8af0tLdU+f0
cuK7ACxWd4NTrZx80BHg0rAooPKdyqIzHrTg3J7IH94USXgMGmrM/XdzQogQW+9P
2DYzEUIwGe5qqYp1OpmISbKBDoRB1ypyMUzB510EIEqSHloDfY5r/5myMn0j2CYU
ci3RSVrGukSo+dz4mhl2MxvPAloxcJeJrKWaWRp9f/xS9lt3K2kSC75TiO/p6zx2
cKTfJ3YiBb81vBjvlxs17YxK468qTofnTQG6vLPmkZ7njaT6DoCwtW9piIUqrB1A
liPYL9S/m6GUOqT+PVYVEj/GoTtaffY27I9bt2l+sMzAHQF03u/6RSd+ryTfBvjf
JGbiKwy6jWhXu2XRcUf/UHIDfZovnFwP4lsGfs459KHCAXdv5PMyPsLC4DNMpDlH
5zXZjtsIIXJCAh+nEqhaIANUyXs+IQpRutBrs5N15wyuGi4RkgENu2y52u2UloKD
NJRHaoPQvGGJKmWACdpIAgKU8cxwMiFUSBfZK/I1nJ6g8u11on2HmW8DojnfOZan
UP2a6oOI41ocOGiDlmU8voSNzurgeXFH5uhzyNcMzz5gdz/qXr6XHGHYMgtUsiqh
uD9LAvRRHHGlSdUtKUOwMFB+dezDnp85lx0wNMEW5uaiuPwkjh23JsqMKjY7hefV
+1c4D9Egbu47una5qmJJb+mk4PTPb2rlgMl1LYo3zP4QTJbfZfIT8Rr0e4xshOVD
WFGCFIUVk1Msb/klmDoJRO/X4Rt8XsY/J9VMWBruKe2ieVtxWWdIQFe7C/NCFKgF
jCXaJHNRDQFHGtPMTUZB+lWpZsNP5Wof9NXMWq5R0qzk7ohsETgP53+LrqYZNbeu
/MxkVntK2iD9V3fXrAUIE9+7gnZQ2CCE7mNfOe0XkbEYXj79vRgYOe2T/03DNu+S
TATqpMWVnhvsZTJovOnfVOOb6KR3ZvVul5t8TzwFEvINM1dMExAj5wYESDYyIPDH
O2n485PJE6eWiodN/FcD1TRsX1wpdLNU3GdeNuMhIbnT5/YYqdemBzQT3A28kvuV
G5IImN76zEPoUZTLJhzfRW2BO4IMukWKTBqHSsWkb0wj1ST+gAVrphu8xQFTs5Js
Te0VgKkEe1ndX7m6JHb+h75r72u4IYhxNN4VeAWMHsMBzXmpOYa9LQxQ7IPfQ2SN
UEuF72wlygKQPt1hGQetWkaak/kkDc9P1NdDtqSgLXnU4BABoNE43SQACkgCEfsM
i91hn5SU1C9u/cVeiXrJeRQbyl8qrg8VkJHfGSJdDTrGhe61nHf3UT+5EfsloZkT
5hMzOapJEsArYv+S6osOd3xUS0CwZo+J0mVMlCEflBVi100ljZM/z+eJC+uxLBIh
+bg5LElnP2tR1BwTDL4DSgYULoMs2kneMF4TAHhElsHyl81BY288FEC+eFMUFKj3
dv0pITWjFE8srDT2GUjJSi45uASE8iwaEfaRzRvjZpHuIai/UYviiKZkkYQtg263
QDOiPhp99CxUsJm/IVold0lTPsNp+07RXfy/Km2jUR7Dj4MylkHsSZCr/kGUmXsD
AcEq4LGdT5yLyn54vMofa085VGrgPExC5QzhN35tAQPHCKC4CD8eISmhlthlUNzN
ARpD/DhnlnZBTHr8Ehp6UsszwyW53X5PjkPhWkVbyD4euUq6MO5xgcEmy3K5oMY1
7uxqatOdogYEbyg1GbSHekXc1B+SPIofA1K9v9TDLKZeCqNkH4cfJO0IC+4NxH68
E9OmsfbMceqU1aOcEuHt+/6EzLWPAGgFgEXdLje4cORygRVh4t7osFJyCvyDgvBo
7NiqJQNaUCNBuTYR9PB8+O0nJI7vdHQFUIEkmW7nvJKTnoZMFku79Oh4JAERmN5D
ig3lNZrXKGQsvTUJYsOvqkavXhTJpWNHDEsBqqDJwCHqh9KxPPhHrg1ASOmXwLY8
kEhva+QWKItxWnO04Wt5q/1IVk44praAi2qK6YlQKAbuHp8BJG4yek4nO6lPb617
OpVm87RlqX47ptmItnKo3T0BT/cl949PAqRPvwJtRfW1le70IVAP23ovJHcpOo7h
Im4MblHZBUHuzKNoDJaYYSzNnEJCts7kh2BZTrFSkGQOrPEJ1LWo6Rt8Cp8D48Le
8x7ZIjbS5PetMhsifHDkmH8dIGLvGdL5TyWUsKqKcOvMnrmaY2Vi5GRFwzqCYX1C
1IcjGOxB7PW6Dzo3nD95GVnZRd/PMpOrKBmrHNHYWqCMsguBUcU+1Wt9TwSRnrhv
emwWfSsT6j1w/V30xQTyD37te1O16bJOXCePgY80k4ShNCbSj2i6lbh1eGex6DPj
mJExvGsDqFlbACkKsP2mlKkGYJvY8vrZ1pJ+Nvi3HYKtyu/Fgs1ajcPGlFoAw437
jR8dHraRmyFdRQNFKMXBb49qciwg6i/hS7s8ffoumJZzdCpAimAwIKLOfqPvEIVv
SvpWLqla9CwYypncDYQFUUgEl/1sDaQVXb2pUqAJTzJS66bLN8aoX1ZTbjrQEBdG
q8lTsrZq37MI2WS3JD3yiOd3AI4LYfS+U+dy3P6PshPpU1v6lQx7pflycM8+bA3d
TDUzNe7hjkYxgns1qBnvA5oLXen3dmQpAyE/xP0suAbL9rENDAadA4nSV78nnEiP
6h924Vm3Lp6ohpKDRaTCnz7zQ5pfi67SBSmB/wgSNiAxzvVKV+6asGiHYL5r4hfi
h0U9CI+iPSSYx3us+5DjIm6Mxr5vx7xIx+IU7A3WO/rPo+0wTgjGO50YfcDGUKxz
OUUAL9+NHPlGBlYQfJUnCgJql8K8CpE43fvMTpnnPf8fnH80qijKi8D8dPdjxmzu
XM6tMQAOS1Xk+Uq2ol6r+H/G+sXtBrTu6NuvdYOcOcZ+JOoc6wzylNADzuILjEl7
MXRsK1LrvQRZyoYg4oqdIIdiG03N7pbSDfQluJ7mpng9NmIw5B42lcnOZUmqvXSm
+dfsU9gWUBbk3gwW+MWNUmm1DDEOrNo9UrY5CIpQbOo2hy3/Y8a2kVfOd1gy9VKq
S6o+asu28DRET2GnKGW1vzFmSUI4XO+OpAkm2j4vx+lUC9FWd+zOOWQyDrztSoYH
pr/58AQjTuobj30+OZWjPLkEW0+rnUux7olQEgUZldW+Z9zotuhgd+MXqyattaiw
xuRVYEnkQVCb2hYUqcI8XwDkm2Mm3IQWmsEBOskXM1nBSchVFacHwRPjm8EF391k
MutZLBds1l7j4BDIZf/JjLGLm4Cwkm4Os0H+fZBLQAlf6rYWTXoAOWE1bajjlprA
cgFkxHvqw0zLOHcc5FyS9K64KPXMIar3NSh4DG9aSpiF25A/jyoSYBLpIxCDwnx5
3F1vLf6wT7jV09+hJD6qdzPiCPTAN+M+eXz0Gc8GGnjYC/4THjAkGM8fSilqk3hm
Se+mRZp/sjyeM8M+80PYYixyEsrrE8nZKRe4sRQawAbzeXMwQ6NiFqu/kANuQtj5
xXW45QMRn0G7ZomNoIOoCshE7DoOOjnQJgpCb009iVuErlyG5O2t/+8+UMK1z/jT
vf5NkahhY6FhiS1VeIrnvA1qpdAllecJtzg4nZMtWygB/7Ly4030TEj3R5LUw2Za
VZI7NIudWINFDw1BsuFh7Dtm3uwXZvqmJMVyYIZYhb1S20DGNvdnWc94y0OXYFNt
Ly2OI51sH0rAxWf+jhzECXWG8PCwhMQtxopXsWRgTMEoT8SrL+Jks1Erlwd+km7V
5kO78wq3EZCiqVQRjLm859tB8nxG8ZvwXxDO4qkA0ouBgIVsJpEpNBXmII9Kle37
5xCprZdy1jjZtlH+pm58EFJLkSi99PRPptoX5lawyAA5XfcJsq1SAPL3DP5fEVSE
j4++Xoc+JxnPxOF5sU00XhHx6uJBYP5r3Osr5qcW77Szo4WfEUSeo7K2gNyICYtK
BlU8MeW6fCixLKsLFWLUD+YD4ayd4A959juDsGpq4anegBbIRWii+QM6h+OWfCLo
EjD2rKeXuTvDM2ihWDl9G163XgQTZunJdpslp5YrAXuzWcajHrpUjtqEItoInYDU
TV2XY2cAdHRz59dR8uzFnNEjfE4tw9bzfw9pPd11Oeq0DKL3IzQ5NgbzwExs1k/i
bvfXi9AJNOweYjRvQvZl868O8ESZocWpjhX9/OPYm0JTRV0o/Fr++8z9YUBSdU0w
PNhCxGGZtQ3huZB8iu41LnEPiM3MqLYdAcyI/IatByUuCAkXvdm1eOhCLycVeodJ
dVudBT+S5yZH7mzgKXVb5jG42KVrArtSQ+ogGtqOeQyQV+yuX3g5ZCCIZyK62Wqz
YgnxXQZfVW9IFVmeI2QftVJ3QQnxVde/KvoTAKhP2wvZEA6/HpMAzHuT6USRmq+D
/kjwpMqkVdBV3xjY+LNDoqOd//oX+7wIVWmxFnfaXNxvoncAy/U599xCngiTuwPU
Zw1+nBVztFh+F0BdWEbsEz6kZWxYQIGorjDqtv6DdObX0idNTR+LzvqiqzFeWFE8
M+lJ5Ldbe7CaOhE8z+PZNo+l1JlGGeFFYYzJ9BRAOOqxgmwUD98JTzoiUbb4bB9I
fzrWJH13bidQ2Mmk9hg9kpu1MwbN42TVY1nGW9pXqjjYv3KuHBp3r0T/VM6VflU6
NDqRd4oxdrwpMN/Jd+wWaGU5OQFT02ABPLoUq/MI4JoOzQamFBTObJc4S8CsteQP
QMYrZfTiSvti8fES+jVtVIrOEu4E9C1n1cWffQc2RJKvWgwm0i/V8cxi1yIWAq7E
zXWplbz3oqoqy+W34UaiA8btCTPtR70eX4537PQ7l86VAhAagYMqklyM9pSz6DOK
SvqWpVjP4ZnJbnD9C+s9h6n2b4+lRlhWrLmn5i6RYGhmHHEsDgSANGnYxP5IksQn
PaiHSWBZz0VjUoeW6INOvUEjEHJvD1Qi6Qos4H0pooiNW7VSxvoUGO+bnjG5sbe2
AUE7ub6omlJ83ewFJ/8JDJSwrrnZVjuWnJEzYbbY6GWLuVkvzRkAttWr3zEwC1qb
p7tCfpa6VFE6jHU/RCR8Rhb982B8mwfOd2RZeRyR28njuftVfeBgNKR5mdyfSx+8
1ZiY65X87sZYbTC6FOaYLBsWSS2DBvWlo1v1OArgRxp3bBkgJCeXvevkbA1FGBT6
KzCsV4mAIGz8NhJCm+/+F2mPVyVEKseQdGXl9V+QBzJhYR1q558NURC311MpnfIZ
bbqKbzxkO7q1nHURQFYcSQKBc5JI/lv5Gt2nSANpHoiJMLJTvdSub1Psv1Twjg1l
EsASuCKJT+XeU+tRFPNFIqNDzylapVNPCUB915Ir8Ii1UrojQxZT+A2op31xLBUS
QQ2zStcgvZGZD1QSV2ysDQ7BsEo/5qrAGwMm5Y7CNgM6T+VsGVxFqHqcxT1027Z/
Lw1/N8Eb1eJpzwMgzyfaDzyBHyKTiY7vVOKrgbj9lOk7zJDZRv2g5PXStJndX160
rEPmYoqMatFlbI+FIgFHSaIcZ/Dz3H6JBPUwlWOrlLDQ9ozJjrqqvNXxh9AlQzFh
IIp1VaRk6v1c+Pk/6/l43uDMFXJxUAg4K9FaXvzHiCmv9Xt72ARdKveDLtPVMTDQ
xNFL/lyILYwhF5ryZCpdKI4Mhm56gJPykl9kePCW6PmXgxoxpabhWUjYuf9t+Ueu
LlfeGkt+K6MKljjbi305Cw7+O65fOLTDzQ/3fCdPZ6klbnHZe7yeHaxHxKiyFVyB
BTfkm5DYzMfqk42FR6OpKjO7ih0Gnmn2vYDMWlV65QFZNDpY/y/nWrrbppwyuhbx
I1Xrz2r+ggys4Da/ld/6GFCIypMRIRWMnAG0H+oTVP5c6zRtoawFXebC/OMIbsjM
6l9G3hvSf+tct/C3ZQs882zUHqgE39kwmV8pa52GBEVY/q7SgdnSg36WH3BWVjCT
UdhY4tnBLKLaKFDcUDKUdaSpLh5PQOYcpQu8x8YwQJwTdEDpn+wakhnZtJbFy/rr
J/UuyuwmF+ONfUsDkl+s7x8t7L+zFRbXY0SZPmlyk8Hif0j0ynCrIYzgaODC+h5R
Kk69zZarm8eDPcRHOGFSDwU62VXbD2Pk9OXLkowvNK58nTsz4yjoLXdfywEUXKdG
p3hzVqvUFdj636sjK+2IHP+5pavqTKd35cVkwGa8hFK3Q2Olwlr/rd3ttM4Eet8e
aEBybZY8XEVLJWgg1imn6aEMQyIuM434+jEMX9uuFSk7A6B6ANmKBw3Lsr6IJ2CZ
+C3WZpaYMZuPUJSR5YhN9bEpBXfY+irH47nsASVAJifmBZrBBagaK4zSKbRT/kXK
FLhDZc/h5bZGrM9OR1B58k2L8OCWxtkmgBqmWNH8w51m8vHGqhnKpxzdaBJZXmkh
gHh8vuDCk6VphcmfIPiBWDASlhaw4fNgQsxgQe1XBBw8mSs9QB/El8nVh+Cs6Dco
WJl7V2q7kKBlu0jnSN51pYNgGfNyvS6sthzlcAcnpmByQhHSeI/c1WdxN5SKlZnD
60EDj+k48YxIb+nEGA2eo7Arzabv1GXxK22LE6G+pCE6gQIW+vgyBG41f0O9YE1Q
OW5pO2tKUeVlnAqhRAQDlsbHsRGiln+zxjBPC+5vuRMxhZZbMOkuxpnVHcjU2URf
d6FUYj3llV2G1PhLCp0PpW99Inv3pyAk0GlyBgVQUafYrrWxUqV9smCNpvO6aFVG
9QSZckpdwAahdzPSO1FGG9YdYhIoxbtR19Z2ur9Kkt2FkwJ12Hh8HblJMlsgc4XL
sDrOD1UTzYvwt/Si7+2MvvapEAEwIuBvIBxe73rvf2xMteyq1An71/i2Szs3Qgco
T34oDiTZkagfhWorfrO3iandEMtpk5Vemj+pKSVFHcWRoj7tS4WjWevjIzaJ/vk7
E3hjJWkwo9NAcvPk8WDaPtBNkOygSaAUrgEZBbZD5+Y5UZB//5ugxS4fyomnHvHM
qb3HQ8g+vSEcwm/JGxzsMy1frv2ps81dccfv5HkLVgtGMtg6vX5SFj+/olO/9EOU
qB26rqiLfa1nFbcnXJ7uFyfwBeoDUiBv4+b9nZfhR0FHC8wUcZ2cPGLzeChqgHpj
a4OZijizQ2UXwJ3UURUURvFc3uVziMEOD5FHdcLFGz2FiTeeHcwW+4w16aptuGIC
h3I8jXQtnv4A8/LFZrExH70DVeKv0/jqvbzFCOgDzkq/lHpBYhYPDzeGvYtbmW7n
LfcyZdahYzFJAqGZH28nE61c6pENif/Lifv/jMBzWhf7HS9Qa9u7fwP8vzbWyqqw
WrkBUzM36XCWGs+xn/8SroxJrzHq9uypAToRU5PqDpGj07K6Ogj2po8ig6TO99/r
qyGz119tNTHKab6vIs7LazyyMK7Pa13P5E28lJxNO+BCnJ4kEm4dOeNetrz0ltf/
4+RVG0jUofwECTyyKLkXWUnwm27vQydXdQyzZjTE+N1TNk87eGQvpuzGC8Rei6s1
Y4ZxnU9BFINccyzhScTmnruyVVm7cZcPyQzolb3fCY0P0477Vs87HL3h5g8+JvOF
YaijEWGmuP75vdIUoDEWIMltNfCKobeLkAuB0X7uIWkBl/rVxK/z5NTkuVu9FuVG
FmrKMCtf+OO1lXpdq8hmuF1LX3T/bMWxNppSJjDaFUPJ+Hg4MHMY9N5zjxaElWYe
/mOOlIl+h5OHqi9zqSmrG7voIK5j4wQrZiKeKn7cZdKDAS/oT3qZX4FC1nkTC2kB
kjdyzUbBqoa07uEMq7qIgd5JnQ1MswyK+cvjtKFj6rET+fn8xjSbPhMyxkBPXIDq
RQQSA74oxDEIqE1r9mBDQqrpo2RClT/cp4FHie9bGhW6pvRRJayS0IG5bxSNnr5x
pxkgxBlZd0Y8A1PDCY3bdGx9PeCi0ss0NqTgVRkO8kDTo+ldL1chF8JeWae/2f8H
qxwJ5YrkFIvc2f0NAklRof5KrEclQMjQgdLNivD77VBHM1peYb60DuClhewsBFgL
SUlvCXhriyTNzccF63zSdRPENFN8w3IKBevtaLqsvGWhRorkTarLUIT+5y63NWd1
E1R+fs674Qy0eFhrP905a8bojyVKOGbXEN9mj4Q/yAT42eWURVjKmXT7zwx3cNuq
pHid7IRXVwfX0p0LN2wji5KCGCFI+Zv4Bm5YFr9r4aDN+NWEb4U1+L5wBcJtp5z9
qQbLUOhr3idNTDck4AgGJHVK2UyIgqjnraJvHyzIe5VrZsM9n9ypBOJxgmThZWYA
G0vWFc1dDTRDGhjaH2j/RRKam/PWiLG/jHK+wiXogoANICRQdkuJ9P1ZZUQb6cnN
c3ZCQe8J8/gc4+TxM+oEJN+zMpabMHLla/ZHGi9dLIRF4e8qpybnZn9CDhG1DqUc
XuO6xuLx4hAJZwgjVeT7KHlTzLrgZ54iL5NylVdXftu39rryAUusC0UztcQj8cZI
MBkbIUgHIddeUD5QH7a4SwNlU8nNt4pOlVDEgzv487zGgVF24c14y5KVUkr/FX37
TAQjc9P1PcKLpYfyctx/S2kSS552IScbewk/W/WryNYYkN8c9Jw/zhAvxdJ6R9C2
VPR2ur9T3KNMe6bCrHpTvbfBiWHlGTw2jMm9Wka+1x7rcb+PDmZWrT/lrCiXpW1U
wZ+BfFouSB9LCA55CPOLjucRhUc2DDB51lIEoD6E/kS7qFDLLygRqqGf2H9c0orl
dwHCxgQMYw2pKLIb4nTpSvo6ysym+KLTxRhDA4kqCYYo30WPy/4n6SbWYyPWf9I6
wTeY3X4zsQxEa5YGvvezeFZwz4PbkL+pr0HUGBp96FibsniWqEW5RZKU3Dq2Q6hQ
DJrPsvb66Bv1RkGiBJuKd/PwfBoOPa924Z82j1qTRWaHGXldwUyFbKotpK+rLGxZ
7riVyCDQx47t7Nr3UlkkM5HdSQzPIMbo4yKnxz/rMw7+avwZiG3Th/7Z+XQ4TX5p
WxIiqfXS3MVEgpjef7XNFVWe7fG4ty+0RPA+sqyB2Po4iy491zOSa20wKCdhSYlE
isMO0zIkDhGEFASWVVVL8wyfe7VAx6062jt02WqVu6etXU42YBtCSoaR+7M7qlkB
Aq17BgXAKPIoH4GKcZXKtjDlu4Vk7Z+ecR8iXg/ry6PmF2e3QGl+XI653JtwDHL2
bgAV00Md9/W+H94SnhN91n/AVe5mvKjSikEmLx0o/S6W0Ue1z5OJ7Xh8OjDoQn83
lGORD4vmJ4FbyGMtpHkozIK9oBPQQvOrEOTyGpW/B5GO9ahbNhVREq3IGmk8Cv+X
a4D6frDYe7WddWIMXGcm3HzF2f5MJd9TyJKTyHhhfsXeyRoAJRcXpF075vXgm+xt
ogIDxGWSc+07FxBxIzDVyp6z4Fq7ZJIyc/W6y1HhjYPrDj5bQFuj8hv++W5cDwIS
ASi7bBSVyDFF8/mFFER4eepZF2XNnMNehkLXs3f5wi56WhJIMg85lAVeSk7EH8Qf
v2SP/HfKCsFR1OaN2lze93sGMATAghcIQmeTGvvTzkEnmRS4cnQ3hm8lv73qBGBB
FVoCfEbml0MDMaD1+ZxAR5BmnSUIdTE0WruCfLC41WO9qzZB/zuapt+G5ZSoqvrR
A241Fyl5pU/U6hAvXEIUZE9wJoDmg+GbhtFE6MTOQ2HotX676Atfw3CGSUATk1iR
y3bIyLmcB8nTgblN14Y7J5/tCgMcDe6xzQknqrSbugugOWELu/3SrZmoti3EfZj5
F2k8szeKi+xnhEwibc4m6W8MUccto7XPwLT29NHQlVGU+3qReoFd2gqDU/1ix2aj
ul2keFzjJK1Z7v1wFjsUviQJOY+bqEZ/KT193+yhy6vhoBzDWs3PhA6fGoO2djP9
Whf3AB+cWlef2bnJ+fdOXX/2vwkh4p8zIbOmVYVfsGQeAgzAE3pr7IIDEiOIzj5k
oLBJGKSz4ePNi8lyGCPrB1b3cxIorF0TNRDQR8u71Acdhm0eq/SMSHuwyA+SuORF
62bqJm2HNmqih7Dxg920l+FQ91sa3WxT7bjlmI5+YRpCqp2qJQ0PNQSFpVgOLlFG
u/s4fKPs41eBfkPMYsqscd77fsaJFfLHE1KO0C8/PlQDZ5EessZzNRNsBaWc0r/N
9OLNKFJsa8w3ItKLyIrDyRWhVDhC5O1QOCxom5KUOB8ZrOh30ARu+39DJ1gmacW1
kIHuCt8qB74qBUoP1QVJMYjswCPDTgoQsgAzuypf89viryKaU4b1cbbbmF+fnuVy
wBzPf5G6IuVdlnyl2YwXppl4Oml5LVZFEXELZncwy8U0HVLEBiQCbg9q5jcFKlwB
fAyE3PwqhPU7BcaHJO1tnctSWZm82007Jh7ngdakJ4/3vKg0uaFwdj7P86NJ0Ofc
cEP0VyYlngH9sFXRFo4kASCmQUtp/RTIHTbKs0YV65S9rjnV8etcVd4dYT03O5TZ
XyIDAAFNXCQNjMHROv7sU+JSn2sPvSTxHm0qG5XNgftPhKLhFrvUvRCDkKzUWpDV
mq8Hdena0nWdlNfnsN+2BOBe6iagQ58HeKWb7MhTP04AWS+iFaKRR6TTrAWor+bP
WMrfcQmfT1MB96jbMGSoLlsVbNFwV2dCR8RsM4c12FCq236nruPwpdu8RsRmXUkX
5hnuGlVtFwIo0iycqz994wavagkTGtv8SC5QpzWFqb3XloCowk6M+ZGIRo0sxKBQ
8q0+ZB8E0GkZaed/cwJVFwDR5T1pIY8mpqQSlKeBmRoKtA41hzQ5bgzhs0whona4
177VFWK8YrYLj4vW/Wt+a8emDh+q2DL202QND49y4HrbzkahoN1m3Z+rP86qdVV1
79fDgEwoDd+RJpshd3d0BnATXeZu5vh/aAHrUPKRj1IiKXobpgJxZXOAzsdVz1U5
Ye64G3x2U4dUdNisbpYhxqnzxz5++6oXCER5BZY6+pmBQEAFku+PExnHZOMZ32IF
kECyCjabrcAu0BDZqQOnhztbDEKc69IeYLZTpKpb1zpnCce+XZk15jJFA+AkBlcH
D0jdKAcQFB2kqquJlTLqWSDzab064BhQkehxuRDa3lnd0RQU50cFzWUiSyCCQOoI
cJNRP9p6Aq2Jbv2nU1TUktuWm+fZ8+xPCWyDylwg5Ildkp6x4JLFKu2Kb8aAW5Hh
Rb64KvVtvhVqj3I7Fs+fq2Njd0T3d4xlKiFXJqotY6qxIvZvDDxRurU053i6O0Xa
va4K4pEaSe7dqzPcLrpQ5IvGW4ByaTxIBodvKaCES5XtJ1lPYVbYaD8uzc98tSgh
I5Z6j2EVr7x3GNZS2SDzarjeJEL2EIjdQ8WwIevpoX/NqHne87DDFqUqK502qYB+
vuU9q0+Z9vfZ7zwrplaEYIfDJ41LmrLIXDU/WZ581cvJnjpTBv8tt9KTEnbefPwl
4wh+MHFrne9kTivmIWBcbhz5BRYeO3MI732vFjyDtfZPJQ0p50ONieUC11yiuF8K
okzm+Uf+jWI72CuwwWR7EFAPrCQOhyEQehKUVZY517PxXpXn16RQPD7MPDelJxnb
nrcAmi2BkcqKErJRaB3qCX1iUj2jPov8mDIleMfafWbXOwSetTWFdPORObGdr87i
JQFTkIpXiDQWGLzb9CEZEg0D9BKkaaJBTiIlqphKTrSgtEHnfkSLIw+Qwlxoj6eo
QI+/105TcKM3jcblB/ioO0itfaSTi+jD+GUBwhMkVQvt3JRGrSLw09raG4/B6rWl
XLevaTd3nAstPnvoKJ78+n9puFBoHmSurmqYCmwY3ftEPeehFEvPmWaYvryd+ICT
SBGi8O3prazgm/WtKIopNY0N/b9L62T51Ky58QMy6kyZLryMUeNYxq3Q0wRUN7Mb
Hc2lapoYAVIzJZUe6vGMrbhrNKi/eELdPzODQeHvK2JFOd+Rs/Z8Cga/QJjIY2M3
+s0F3v/iYzbzZh+xCNOMaJ+4fIzZ9ui7EZ8klxV846C3KBIvHB3IcgQfvyzgJEWZ
qtF7kepDGr4e8UggzjuHH01NNIu93u8cYQAzjAbbDSRiRsgksCaLw89XcPAyzdYX
D4BY5acodzmgRCoIaEsx90rM67HzZy54Qh45IKteHjrZOtDgSDajUO087J1J9xh9
C/nSXILFbl0H435g5yU+y47hyJf4bENwMMYAYD5sq0rSWrezLu9vIHS/7xRpnRZW
Imc6sVTcbt+Ml1q7sQ5XECPAdhvt+o1kh2pPGqKYcqYoXW/9vucQREpiGcQc1aQL
FV4mgOr0ivwWaLlJqJD3yyAXIYZLDJObu/EWuUBJFWsEZPwzXqdarUOG9Q8vINgK
9cGR4RSgBjcBTErVi/2xkpqmCAPIR/j89UkZ+oyvg6/n8xrnIBBsys58Z0H1HLvy
eV/4xfTGXlAQXqh3BFahZ/KuF4GTKzt4EpsEuNelfgJTkWJF7p189Gv2vdEVVsf4
RvMsrVYXegZR65S9kdoFdZqBJxDYglj9SX88SmzgC7yjZTkk7qmEOFViPu45jZlf
pXAUPdVDQyhlU/FccrrxSbSfkR/1JB8u91wIkx5T6uYSbsKwPnYigt2Qs+uM3FZ/
ww7uA+/LcCCyhBwlR8eDffKzz+gyoAv+WEDL/cUd0p2SPtZPPvwLDGPw6z7T20sH
bNeQyJ6+S4wypYDGQKKV9piX0fmkkJdIY1XNoI2hRAKDgvYMinyDX4qydbbcvUjM
0zom2xBpB6kpqCebzMw8JPe6H1rrGyejKBqJvoXHYv5ZPQW2wj8+GAwM+k2nOULh
OS8OBppD8+4XbYiEMSjOlAqvt8xVMo0wBctq+PGRbzujDf9Y3ZdD7npLjzmaKH/P
N1vOGrX+21xNH5kv0NVB5+/y+ACIOSHG4zjYN1FaJUL5GhqUhWGXBMxkT5hqk/4+
ckhlgr6nX5jUs8EFJsOoeqLx/laGOL/yNbRfiHBgZbvC5dFA7d5G0DGSoSjNWQyN
5LXDSwANHQb5ZCVtiqeFhG57XlSX6Gwi0p/Ex1oJ87QAQXhprv1petddUeqIBgsa
EAwkw5kLy40F0+EuxBG34htAxVIWFDUb1Q9JinUzwmznziqFXKze87fl5bB20MzD
dUA2L6LBAYJnfINRFszVklk22kvSKIUPvPlBhyaurjuUT/Qp2wLh84VAB87tGyl0
bGBRtXXIxIfDS3CQOptLHGLCWucNbiIoF+jXFk05VzKOFvwDy4ppEbfdR858lERE
4/tO5fU9N2yNo2kgSRbRRl3hVY2yZ0Btxuku0VVI9QHk286G3ZNdjD1OOaFf4GzA
x9OqIits85+XsVpNEq+4mL9lMYT3WV3jjeIXdb/5y4HYb5JoiFeE+Rck98F5O4QX
IUIooq37PXnWqHKnwKo4UoPG9y+7/mdmh3gha5vctGnLvt3uI3EfMovLbBV1DT7d
3wDQ9QGnEQs3ykIWrheVqNcRGrcqkJ7jfkNg89yAbgitjZH2BNQDhNbRJ8ZqGgdD
viss3bxo2QojGV8Fvb91IzvCD64+73WDWV8HQ3aS7XjElYgVIxSL40oVPeGeRJNL
eVrqTGyVIYHodSlhIshdi02eNGgXn9UbVqTW7F92D1L4kcJHC917DlhOmapliZSZ
IMUo+4Q8Am/eKEIVS6myeyHWStK95LuJHFYyIlWVOrK/5JZ2Qxi5MduI2DCpvGOv
dK2wN7n0FGuev2//+mh4svRP757ju9M5YZ2HO7nbv6uresu2FkO+ior5fvZgDgag
+BQKDTswH+JGRvaMIsi9XeDk/wlT0rs2Tu6pqJi19sYP30fgDmMu5cTsR8bwbWVj
9zrSQQp0ZRe8vJ8ow4y3UtzfNocfvL8Xa9k+gne2JpSxt3t735u2W+dpIYq1IFGy
ausD30PboXnnlMiirPaG6B+9uwUHxZgOU7QQgIZzQyR82PdBHP0hjB3ozdiYJNfn
olc73pgaP0jo5AiFR+jCvD5yDLfo6Fun7KlERqjZSCmNTTiqO5cV9hUvwgKzBNeK
5KB3qzO8y6yoHGQ41IKXYVmNi9PO5+1RXHaLvMT05j9fvLP+8MLG8Jc9fHWvGKpW
itiGNIm+FluOVfCbycoc7XqnmtvJ/oMa0sI72kenaJGX0Q5dulYBArRWJwY08kif
eZALoEKLUzsksBH6lSNRcy5MufdEGG9O9MfRPDNrP96XdHfsAt7FVHQd1zY61uBQ
3wJQm1QwAjvN0n8Eb0PRkroSlasEpazxoFBNTVMHhql7gyLE2xbTZfFxo6Bukkij
UJGcpWN1CrQfozOuAOxtYhvNQhstzREwJ40ZyKstESx0vxXLIt5t11pOEFWTVBml
mbqgq7amGW+m0tczqyE+A8ovv5z1SDxfRq28S40x94dW/DsIoUGplqgfGczUek5b
jdo96KZ5UijpBPsUN08yL3Xsy5aDQ4kqI5LYTt+WCQ6RzweySwbOS2soKYTSRodc
Ly3C7ZEFkYfeXU667zys+NDfAYoPPixi5rqS+9AoCR+SM2z70VJEFmbGTHT76IDu
wBH/3UedKPuZbHIEOJ1ByxfDDdsc3MwRoOrdZ6tpBAZbU+yLDNVRH4zrnhynTeY8
irybJ5H/Hma/tN5/iwbJ8sX5MWBCq/xY7Rh9iclAudexOIzV2O0Ez76b4XqOtJQu
YMaFT4vt3eqECChlJUBuRRzAKgsPLPozJS+rnL7cZLuNnyW2VJaOysbePT6twNco
FYrbo0Yby4EW8maZzxB9xYds8FmS/mey3FDdPXhHudeWb0by8W5GXwQV7o0Brhgg
A0DdRieh8TaLFiGIt5VWlY+gO4poBFmfoWN6bw5owHSXgWJhuMaelJBDvkHTS3X3
jtbcl0WoWNlQxkwzJLj4PH8u8AH3y9s4QGpzXj7I/haY6zkt8TbBdRJhyGYm8F12
8hId4/U3qNpzMKyg+qb9lD+2w8Pso5WguTqc9ksm2iVxopJt6kC3u6AIgfee0Mj6
gKxfTmthYe3LU5gp/NEEzGt9SakT2tBvFKSIFrkIuQZeU2cqkucU55HTr4KRWJQ1
1JZRZyNqVQ/oTaH/6o0AfTczbAS9Ft+uWaOUjpS5e5g=
//pragma protect end_data_block
//pragma protect digest_block
9/IV+S/Ih27FhrCOalk+vUf023k=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Ho2alO2qX/30hZgbnzmFwK9ayZJWy0wzdvrkRFj8v5bnqPBci/tyX+KSwduqG4yQ
gN/z6lJnxXWFWwvDaWSpGtJAclxI52Ae2tYAg7q6p8Z4s/v6FqK4dY1QBrQpnJvD
lIb8Tk/2g/6kMFPYMDug9Ta/XI8DDUn3Cf3qlck1idGBGsxsNHT7NQ==
//pragma protect end_key_block
//pragma protect digest_block
MM3M95/ba/pJlKgYRTOHM/09CHA=
//pragma protect end_digest_block
//pragma protect data_block
9s0PbsSVQAw1FTfNdDpylI0lRp+FE4/JiPBJiCW7NIwcCkeYT5ETdtB6of13YuOM
D7vWf2Qm2LR/6v3CgjloFfhyLGHDQMlpuxbUdIPyp2/9nYmmUnPQTrKWuFheeaRK
QYKNCgBnJWko+8u9NhHOZ+riW+V/NEoksJVjo5UWPOfehFOjQIOn0DWV2U9fh88G
5mHUzgzavFZcArjchDwd7SourEGWotI9BnwfY6+SpyACkdnBJ3FF6aZZd4fdbbJ0
uQyjVCCUK/AoFWg54dPY6AVcYz3+6H3DmP8il2T2QwLGu7cUqNJR16ywXgSQSXqv
scQZyIfb7sj/dPoZhV8hta5ciaf9T/UOBeUEIDr9WnF6B4Rg+kRdlp38KC1eKs5M

//pragma protect end_data_block
//pragma protect digest_block
bOsOoJdIuYeexxRawJ+8Dyo+3kA=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
n0ekQ8WvAvIooNCMu06vL6bsxZt0BoGKOIYYw3/uWHjUVqRNg8qj/LNGyC/UeU3V
QE7fgNzqVdDyOwtW+Aw5GQnOY5MlSzDUSrV0p4xlhyFHxev+FrTiE4zTEIhrxwWe
C3zv00WVcshLM0LnvUyCFc8fybnqVuKIhlDsTs9flhi6EaVo8BNgMg==
//pragma protect end_key_block
//pragma protect digest_block
wUlQB6erBXGkdvEALQgEWjJDNcI=
//pragma protect end_digest_block
//pragma protect data_block
sA1YnRYTva47wVvxmsnZzdDXA6GRWLldg+jiF1Kh2GSXvHOedrGeOPPK/eh5eqax
jsuhL6K5NZ5YDjJWa6BIuGCKCjUJXP6DMfzCn63V8k9yHvUE49daEI4PI+SdRXCe
xVWYfJaOW9sjj601rVbECof8Ejdr3v2YmLWQe0vrSS/vJVXJj/0k28aDGj8CaF/V
8VxHzW9GHXu4Ot6hUzcSLxZ3yULxBmjA8TpKLqT5KHP6o4vbVf7Ptu5CLZF+041h
0ZrPku2WaTYYGHfCTEpThgQ/bD+zzB+RL/nFWUvKh23VFwprh/Vmmj5150bxzrao
JeRYapsJ1MsgWOXDvbs/dyS6xEv7phLz2C2ZIvQ6wkYwKsh83vszd/8Zg3nR3gqU
1DP39bycYf17HpL9wz8m4sInl49BASWw2clbdkHM4x057ySP+5d/p+ltZkVmVRq/
X1saxRncyDBNDDa2PXzhDFMQODVvWfuWoJdq6LabU5JM/pqMcZ4kHi3yohwD0ihv
7DZ7dtdm2cEzNdwuwOsRxN2/lzV6cGIMJotM0IOqfkHosdyZXnhfxY//vIkM0uwz
L87UkwBGWv89t+JEHTnSxdswYXRQAeZzEW2R4GeBhwTbWNLBmLyiUjNO7p9Yv05c
dbozCdQzPms4uSOinl9WKuZZIY01qdSJfep9oc1ZbGDyHVkto92bBwb4FD27ey0/
eaWYovqb53Ffo2fye4w/z7S7w1JF7N//HkrdAPusK2v9SVWQZRzB0tLzXh7m7ekc
WfBKfjGsraAXxgBJWzbIVTBUM+3sm8+66fe3/YZtl0Px1+02SZIrnas3PYlqkOPG
QEH1MEkGXl36jucX3NZG/+VcFGrvuf01aJ14qmEO9BDCqWSugELiVkxfn47vSw9p
b0wVntEF+TNhWYVesIRa8lRSuyoWgg/K7JjKSdy7BAIXQsbF3LSTILv/FH3tKwoD
6lszHNnq/ttgPMLjKqWus0vXauyMsx5u0UBl1bLKu4uCE+70/ohjmXUDksWAa3oH
BFIsqNT/KDodI2uh6+76pFFAiKTvOepnkiHo5lZFofwU93MWXztnxxNqEjWOcrmA
/0gr7On7RH5OvLzJ8UrOqMGIwaSYUWnzKwZYqPdYwAzj2whXlxamb4AhSWCYNT5p
bN2mdSOBjtL/Hi/CNUB3Q/yZi+DFeiZM8HxhGvqlqqviFa/dfDkTLnn1bga3zSS2
QQjVmOe81rmz892iKK8ZXuBJmEJ4Vxbxck6k71NK9f4kKuWImqZWtlrDluOq23ON
rnerBykzNTOUcFxMVLdQ8plFalus2cC1xAGm9ItW794ym3GJdckRIiL0Dsav6Pjh
IZYb9+OEN3vnppYIr9sUJKdRIpAwQfexGVOUbM1t5gsVcTayxhpo/zMtM0e8HrpC
8SSDS+IKVQoTJBXrva1WStOiK0cUtZBOQs0ljg5vXIMx1L58qfDx8Jq8gLyyA3IM
880i2MqiK/yN88D8cOU+3sGRXoNYYlHcHDNSR71vp+5KDKhCxx+zxPmpuzHImxEm
4/uLebT9H6lXKJvLNYGlxORh7lfq9h08vpXsh70AjCa1CJJc8NWhAcXEH+OWVO25
9daiVsjgIoXdaUAjj5zLR+JAts1rue8WoRQZWWzNvEOwCc1INPFnisBfovh6Ilwy
08lmpWfnMeaLZjnqzFQkjoUEygKqH+JlHZFe7gFclKmhoGte74i8aSwZhdsPfgaO
l/dHPwmDFfTvGLGf2A/RTQquPULPuuExmgQ2gCHnyeQqlylorJu/XSNn13BeHOgN
JKIAo8+XDwlnHc/DLhoUT6jT4c2j71FRrxvuhi2lprGFZNYKvKdbiPsCIVZwzpn4
Eag/M9YKgdLlmertUfrQGBvay/NKVbKy8dxVwzveXOIkDGbHWGdImGiWhngmWNSY
6HvcSOEYYQ8lFi/zG/8vuviuyzoApWNyQh/ZEtdQUl1BCXFTqUs85nxYAfpjJAO/
4tOST8eag0z70wnrH+hUGivsjzIKdHvbiKPHp5npUNQziTtkmtt0kDDlpRoMPaGz
sehemVqqVYsvARhBID5QQ1rbY/ZPrOnHDOBotle1zpnZRDYV/SPediz4Gv3O/osi
oOinFVZgN54pp60JpCPnleYgcQ+J1Y1M/rxfmWOFTHFvoR/uh5wc2LsJ/cQhFkpQ
CzgZsmv/6qTh+H3uiVIiMdc5AmwwQCgmu+ubNoVOT4YEopP0DfVWnyuW0dIecm1b
nk02prPTwSJW2DgyLNZgefj+ysG+4kj7I/7B9MATO7PfU91ZAmRV5dzc6c38Xp3H
I3M6s1SfkvTXwl0o2CvqyuqZRHKuAoKVy3y2Nm6+oYnPwNRwrvhYCDybj3hAPGLO
6b+PbFJXVKsS4yttngJeFPLrIk1RKb1hLSf0fmeTYqO67+APgo1Pm0EWBY4lrXfx
JiJuAO+/KblpOXEBiNPHPWXc1xHCtwVpMOxUKq4kRc+fzdSzpO4Nd0RZRdxy4wqg
IKA1FC0sj3GwNsmJrSe2ndOXe+w/RhPTvz3yT+4inCLyB7F9ZvijZClpCT7ap1VN
kKMcGLBx6oAkaYQnfJLNg5JnAjTSS+iowTcMwuyEsLxSynsA0oEQFEfzhmDTNua4
YC6QxheAd3bXNnEo5K7zPhnfk4+Leif/iMEXOmu46pbDwgjxQxQJV6RzDeA4LijJ
xuVfLaBggUxTxn7HFbfttoLj4DgxVOxDX7CDkuD4ax4j0LmO01bcJC1pZo/8tUaD
hcPt9LnWjQoR5y7WpZF5adaBUYEVnqsRH8E69T5ymU85AT2WV8Ea0f5fRxH8SCpQ
3JIGHq9JRKTsWeTIxlskwu3vqHY2u8BuY4D+yor0jRsxUapwOZEPcOFt7YtrAH7/
AaYL3l/CVvdyte25EBetPDLXAfQrmSkvsN5H5IME2LSDSe7cAga8KYpGFV01263X
nd2zsNuf3m3HRVClAPmae49qJX3G1tfV46eeMBr2RJmuP5y4YVDHHKm2zplAva2G
az7wnPamhT4Vii8LZq/G2jZVxt51MwkvUFnSA0qtqHK2MU/IIkGDgBdM2bW7iwnA
7nXTjvB+6QD6KL7TWzHldYPzGD33uJdjaZ9jmrysJ1v1Od2enhQWAr+7cqql8HR3
CqJwkAqnl+BWNBfzwjimk1qGyH9x9MRc9DZvOu+ngpH+YSyu/5hnIOg4ElpGcXCb
NfgUw7BpT/N3T0J0M1DVyCEk5MjoGHButLPXTQYAIFsTnSyP4Chts4iBkSSnGJ8v
X5lXl0jvMvB8GoYssVeH1FYLanqITj9hR0t6Bi6XS5EgPIWfz2mg4Y2N+G9H/xPP
UP//MustEJtxnj0fQOP7rfPSktMkQozyHKD3dgZ/vMR0aGFaa4K6gCA8LMpKmiz/
RniUN0Z7il4hCSRMlMlKoSeOijTfNrVmNbw2505QzjJvZhnfomZ8LB9TTjHjQ/yF
8qBFU4D+Sd8BVZbU8HIhbYl77Bq1XMy/FPa6EHqYUzzf7Lga1t/gxD8gUo0KWqZT
zXXBv4SAcp30oIIJFoGnOCFfLhnwnspj7LS5uplsKADmbimkXjvQEhz50nXqlRTn
E+pT055G1N/xuVPxi9ESWPMU2sdXC50lTRG8aRPYI6osu6LWV4SMbAgjPXVvUYHH
VF5ey4poANAsttrOxnmOWpDuXsctkGOaGu9qIIBO7+TIoTOszYWqPWDsvL0hhH5z
fRsQjMMRMbN/n9R6DnDuzms7K++phjhf1dIaR8XNiUqubcchtMbLkFAlqiJhLaXs
m9d2RPnUvFshTZdGF3mpj8ZfIZQUE0ga32nky/7RIIt+YcL61oD/b0VUt2Ggvyjr
eX+uAXZ7TDwnBz1BEaT3zZYBw6JOoMbkcZGQ8d7o8QWw+cqgofArkHHYlCMI4pjm
F2J+hk5hqFj1zDsPDWTa/Y1KKOn9bKHOq0Z3LGAqQMXw2JguDiSKkDre23wQv2Kz
Ekawd7KxlsqZT/fv4FKL89clDy0kxglMR+DAAjpjnzUXiLpkzW6RrvReRRgbXjd+
wIaK1QkHgWsHe0xBgkLDdQwD6X41bEV8MjE8jpIXo5mo/qsbVJUOD6LcT4+shHrN
LWCbVzfvvYW4ElVstzM4X6dWAgHHamQ/QxJhlDwuAqOCjhkdQ6JcyOKeQXtVg+4x
/O/gUkw9DyeY2QnBMithqR0/zyz8fBy4VsLtcO7LYhKtFs62NXt2mCgObTSpOuYX
glx5fUXBt5ac1UjYav/8fqZ+06su63wJYLaHPAwjAMrEIRQXvC0bfAlKDm7JPSUp
Rj1QdAKkUs/WOIsZ5CSu5cxrXYggyo801hXR80EZ6B4cKgK0/VB8U+2NYAmF2+EU
acTCoHVD5ZN+jspeMDFZsU7YjHI2C9pcl7dx3Zk2aO/eZeeNkdUnBGS2XKqIxaAk
iQLV43IOasmMbE+hNyhLGRU1I3XArHOn0szLjy6cCFj2GPJB9i9JMJ6a5CBAbtmh
bLbiMWMMbP+QjlJaKnUT6Nt3p9OBl5qX6JB+qt29SQ1dP3n8jLGDB/cQ1cqlxFdZ
zls7mL9dX6mgyTJfjO3vIvPiv2NQnjgqaL8Y/JnT1WHl/5zuqI8qIUAwoRa/L66f
1UvkEHUcef5C+n0CpfK4VE7Hc1Wh6R62oJSCkP4L9mNLqbKBuc28vgbvCxy7/D4l
NV2xSnuIrh0XBwtW460HrDmBJvZGPsy8l3PUrQjl8TG32l5DWKP1mzTb759eUwvJ
Fst3hYWZAXk9tbZUzRSSStvufRcTKvWyDav0O0KUwfhmaX8U46I7rOxIj4kxfbUP
pAS10nf0iT+RfxhtruN5+5PVhXF+JqKLNsX5LAGAaFQKWOeCEGaH5zhLuY2SQWT8
pvmW+whplWxd7/W/mVFc7hobHJaIa45gHuISedeOBUs+4JL8Zbtj12JHoSBVlcC0
QuKCuEtnWSe1oZl/l6ODjLHCFY3kICQkSOk475Nr2013/4eShLE8vJWY1QrR03un
IO+B8b6tpyr+kZf31IxtF1Eldi1gB+edRUKmfdXb7Ge36yxDqQL9JCeC4aGZQsWS
f51Rn1yOTSaMcwwy+UXBI7aNI/qCq9XrGlKjB141vgRxv+psQrH4QbCREC1xnOA9
ZGL1l+1KylNfmWskBb8rwVYOUzLbtOAZTTYtY+ez0ZrI9Yaej+QO9bBwQPJfFsIm
vjtJMVgisfCfqImMDsazko+JOeFjdhRwgaJV5S0fvmZpX8uHY8hZ+0EW8YHo4opW
Qk71+mpWIleT7/NOQTob/mXji6ktI+cgF5d+T5+iSoJZcnwX2XTBkrlSy3e+X8lZ
VzpCb6p1tVdQqL0tC9rfCFg6QU1fbt5IhtbgjxDbvxe3oCd2LRtstv0aXdlLMc2D
4mGxMURp0aelh4+l2619tlwjLOtEc4wjWx9OzX3Lho/SpKk46rwxOEAhcK0FN0Sv
kB1nMFqtPb++vzBVYuXKsl8PtnEIiab/BfrHVyuVlVrxaJZwYQxajRAyr+BVi99L
IKmEXvRjTxC5hjIOuVG2HC7xJcAnyNksHmEFWUZOX9dZZ+yqSZECqd0NlOdXCbgp
hRCbGilkc+5MrT5vejATOSWn6vU9eyCcNcKOZiK0Qy6RapevoLR+7lh56Acartk6
+XUXgxtwaHwhHWcr52JYiPfk416MY4G/60z/vnDCoMyP6R6BNCAlIb/+CLzYijS7
e8B3bIinmVybu/kqal1I8mD5nMsV2pMQlphuotreB7RabcV9sEgcTjTLjvru/RLH
AwYcP+H1LBkokkM7xWfpcDdi483oGcV9ISRB3fyi4JYujq9qW5te2id4mq0oncq/
zF1ZZ8qBjKVGsRmVjuFSSxe//url++HsELDZ2Q69w8cJ5Q/6V13UBK9/BpjAD9f0
84Zm0EuJxGL3r7kyLJ9NfoS+5l618UbTA4ZYAizvfROd++/aDykZ+Ii7pXriEADt
cV9uXo8REjrDqfh/v5SvUUxQSJeTmoMp75e/5kihfWg1t1Juxxxf1VRh49OO/x6K
tw3qo+yPRDmbi+VaMDPb4/1mztahsnrU9urRiFqUSrM5NpZAE8UmHkgZVp85p/i0
GJ3V6ehMrggXzNUgORl3K/lwbUVzYmZfukyH4kt9bBsSyyGca2mZ/1olFdPoODAT
eCEXk1mQBcvBl8sIiiw89aFUUOj/aCZ1rSdITf+y4RCsilVfKo1sAr7oztoOXby/
7icoK3G0sg6G/CxI2Lr8yj4eUMARJL53JwvXqFwocCedGb3as5kAZrulAzSLgPud
/Cqbn7Og3NTGeG4CQfwLVUmS8HV6S9dfnVnSpiZlBodf7BDL0/uJTYTz21Yrrur4
TmEwN7LJEvLcExE9qtH6UDOXOJbdf11aNT9PmdS+tFDz9EBPyOnAwYpGM7ul6BMC
Rf8cvGOjKZZ/HSp5c+dItsQ3NGwPFRew+R7VF57hDh8EIJE0L0prgpHioJavwthF
yCXiD6Fdcab3q1phYRPFQCdq0lDoZR8q+KXspcI1YfvOZJY+kTeuHrSFwBvRXRw6
vTnTSyskvMhn9XOryKY0iJKYWT35szY5YDHw2MvKD9hTVOKhsc0NNDYodyYwPTkl
VCnAK7YyIWCneRUkLiNRJPCJia62fBb0BRsBWpq3O/fzelWzUx/n+rcvWB3kpc4Q
qab4uCk4unf2fjcbdEtvZ7Wg+xcYBScMEBddOY9BtEdhnizVQCo5MmKDN4Df6fuv
jULf9MfmCr0TA5HHTyDSOTsPnglZ1kP1TfnWiRr+AFfttuqrYqeXtpYjchp6Gp2x
Bzp/QZVA8XH2wayQ9SZOJUMpbLW6BFdse32IZdHwR1wOQ1rbXvxhjG1MhRUYRmIY
Ye3RqpEgX2FAvZmqhEiCfg==
//pragma protect end_data_block
//pragma protect digest_block
eWMcWRUqpjdWNiVORETXd6hccFU=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Gugnbdk8fbGMphoTgcWceqEzDdSMro8PNqeANIkRa/Mm0WcQhadcPayDoy+YrlBM
FCZwdLt6E5Af5VJNDa+7/dPE42hedsvFJYYikzhUmRep2u0dLHnLHIJBjFA1QOMD
uXDAS4aF1rGCLCDa5RlRLbExdK9ZFqoCIY9mjBozNPCczN5SzAhhfg==
//pragma protect end_key_block
//pragma protect digest_block
aO6GDKas+46XLMN/goW+8o1bZSA=
//pragma protect end_digest_block
//pragma protect data_block
8e6Z9ut3wytYE9H1r6wGJQNCqSKEBFoXxpGWBSyuyNxr2jwm3/Wfo4vm9Iffd3iN
jxhRVPfFYb5zDsmjn1wZXfnXeDBwZGY5aMsu9gB5q9GZG7Keg9Vr2JrH6M20IIy7
oa4zp3C4PqRiPJW/YmZ1hVSVcVwp5DlR2pg2283+zfQ/DCuX9D/7VmCid9lDVV7Y
zXpfe1k/fb6N6RfBt8PQNfqdTTiJbOtNUiv/3M9D4K+sHhu96tyJy7fQhq3B8V6R
RruUt8UQxOO7Mo2UnBFXyCD/3nNjjv70rDHMPYige054b6kzuklFA1dA1lu5Aknf
sj2zad4OkovWO8vasYByDKj1QUQja/9v0Z6dw7IydTIreoMj8XiLki6w2U0+ZWZ+
BuvZ6+vmP2mYm7zXijvyRg==
//pragma protect end_data_block
//pragma protect digest_block
0t5heoKw/Jm2T/27ELjBL51NS2A=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
r2S1o/aoD9+ZEe/85TlqgFXw44KYsSpl4Z4mBH/4G4RiLTpKtYf1ZTBIbemj4dp+
i293NVFLpK/M6lV+j7Py1PhuHMu56xrhk0muTpGRNO8UZjDLHVbL21LV6y3w/1F0
VrIEG5DHKNBf/Lqmb+Y/jxttWTmSBp4cqyeGmG2/NCAwHbc4EZ9tvw==
//pragma protect end_key_block
//pragma protect digest_block
PCnLONm1nxaFTgKR0IliDwcZA/Q=
//pragma protect end_digest_block
//pragma protect data_block
ylzNGxnX4YS+OpScBMXTnJ25m1/JHEdjKfSN5dUgTN32s1e1XCPzk2s4lgcBPVYF
GIOmXen4zEG/ZLe3GZgdHwbBa0J+kWbCmPrvR1Vb6D0WmPCrQf13u2jWRt6FrXqO
1OZLVd3Gxcs1pRwKUA+ELk1ftz0vCfFofRz3C5EVqdI3Lk3FwKiaghBexiVEiSpg
F5hb2XH6GRDhV1GjD6kSgy3fxiAvNVhkFu1Z0oZdyLDkKVjFunuXai9nPuWYswVD
z0pMsDvP+am16TZ/48N8WdpGvBKiKgjp4k6ECTqMA01XkN4fvai24Vyl2heTO6kz
h9wUTiSI9ZrKCUYjSbndLWHC7LUHvWAUtlbpucVGVaFpavrr3XUJHfWtKzotblVw
W19w+YlpgSc17zHk4JFPprmgK+WKjolMnEWDnvac+6lismQYa+bbg34keJUN3JOP
xi5Av5Y9evWNPencEYtUbbLmx63WesoJAAUfsXoymJ5w/4mm76OcYvRKkNY1yCUr
pNaZzaiCaj7S6WCAHiql0GcUcgRPiMXIBxDFjzXvr6O2ZOOpstWYdvM9XXbbn/KJ
uTzhECPT2mC+KPHeyfxiM0e7sgY5iGRrI1g308opjCa3Tk5CO1P0lykv7nWCMccs
v4I5q/Mqg4SmGP8R+sj+BTPFgmLTZ3jakzQDtoiRclwJNe+po+rVwdYhjU4BOk9+
+5Wym4hsdPcURvUre4dMdT5U0rXYE70W7y851hfknXTqjU1NyH6blRfo2mZbC2RW
TJzNssO+jE/CIydp5h12cMybXQ4I9yFth6gP3foW6O6VzTq1f+n327mnDE1CL06a
43D4DgUGbt6WTjmbcIFotkpTpJfNUsema41Y1zGsJ8bRBiw3hsyyouN0wSvmqtKn
vO2kbyGpmU4S/x7d41Kbhy3HyP/ZyQ52X2GEMzWYEpSWBpjhEt9wuvDasyjWRywI
a5vA2dEYDuDatg0/rQq195MHOv2BNWqR9f+igKFd7VjEULYwCyymaQhSDVKdpEHU
rXtjtsJdWfjfBf24JJnUcRe5kp0rUjft03LV3BwPqLgkFaEr6SMBr+DSuLZykjz+
30AsdSy7FKkiZaSWXbBMEq+p6lLgJplmYqLskQIENlVsiVDXTnl0Hy7lLrkkR0rW
vpUIwGABER0+vRqbiGcQqyGzf4ODKsJSmihYnnyPdehSs1nEi9ppHeoAIgpRhS8F
LWao/t+17+/r1zeOPSCsvuWC51rEhKUes/gUGb7dbhg=
//pragma protect end_data_block
//pragma protect digest_block
3WGz9bPZAiCYV8vu9HEm9lI9edw=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
1sLegJYWfVsXZvzunrLJz5khfe1k1t5Y681Kz1h6jxTOIokOTv8NmQlVElyR85OU
ju0WgK6uueg6EivaForuAKoxxAg4K5dElXpiuZc7qrIKMj/p1bFuyULfDp2g8TMQ
Xl7QPxHPqYk1KN7AU5KyvvnAPvMRxpK72husu8DTgdr2qYxGJI3vsQ==
//pragma protect end_key_block
//pragma protect digest_block
/31hiJeCr5iOtRxEQO/3BhRFZ/k=
//pragma protect end_digest_block
//pragma protect data_block
cKGQ998O8COLjk0JYwFJKuDq91fIf0+QC466FMc4zPr4IbPPUeYKMUUU7izvFCXb
HK85qS1YR00MSiSxyrGDTAzRtbZaNYvzPhqvGFW4Og+dEeEe/0s+/G2CXpOPbqL9
E6XhsQ8bhDlB3UuIlZnwHbQoJrAL064u0ubrgPz02iiKLUs+sJfi4Hbr6T7vhFc7
nMo/2FSTbxpKeeQUGB+eg/ugSVpP5+7CKaQdUxYfPFfGaiuik0CDiYDb/Niinpky
f8ZQ7WSU0i3LQjIARYeq4g4bM/McYSzBAMkugFX8X0b3osQ2CkERwJE2A/uwf2+y
OP9dg3/y+q2AuIjMMvGSMvpxbJpnLlhxLtDF1yTr/LhGUE8mOvC4cZzbFNWtiLde
hgUCJNSSiXJsuzkLelgkcw==
//pragma protect end_data_block
//pragma protect digest_block
aENsyNkD2elFAsux5Uiy8Wuv91w=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
a51bempoCqJrrmVk0Pl07e3gdK/H2dq7bWJq5tKu8IJnKUm8Ua3XAZ3OyP3ByZBt
5j+OneSrun5AzGN3mG8TkPqBgV6w2gLWuVEDKKfv3l7w4LHPSF1z0DxjDpMarUVJ
wEY+Bvyrv2+/TMSvhP8RME0iocDGX1+1Et2db4/ciUHDblG7YTafaw==
//pragma protect end_key_block
//pragma protect digest_block
0yj03xYOCamf0sKi1IBAcGsX/RU=
//pragma protect end_digest_block
//pragma protect data_block
TF9RhRbogsa7ULx0AfKMmNlWBGUQlNZTFdSOmWX5inBBlRvTxdP9fc0oBRYPtTlx
gNffbEbjp8Cct83mcDMLVMeZDPxlebDBMxPdcoc79mMdGqLaTha3r/aftIZTUu+D
G4AZSukNmVzacDiKIazd0pjrZqKfMEIajsNM1CsssogR8b/VdKbBPavPgB7sqM++
vQ8dUk2RQ1ATh2LzKRJuTG3WdQDxvuaNqetmK75goWK5PLRCFfQGBjepJNQrbMtO
2hoSDqzfokNlpjBpNtNOz+wyspJYWvF8DOfC9KPMK1MEyQJVierbl41y/tPHPwrM
g41wJf3+XhZlSYc5gIkA+zXcs3AdpndQrOImSZuQzQpC2mlqzqO/dPPoGOI+BKfL
AU2g30uglJMxgfmcIUJci2MAAGSJHdTURqeJFqJQASfX2OSlU/8e+rgoDOPLO/Fg
gM029nLevvU6NpwxgXUs9vaW2V+S4TvYs6yi6d1QTMaWb10qn08e9y8UDsn0+7zb
5rsxVWzVdQafncEZXvsy+ujHFGn2yamDT5T5ccIX/1wgutKHc2I5Rn2Y/V9qe1y/
eAjYtMtXAfa+XiJ+LwM4NqHgcWH0p4/Uy6bbYZ2JKr1STn1MwT0vJWwMT6/RLO/r
bIUaRQxCNDWwhNnPsfUJGtKzFjjeubx6y8QQhU1PrLpxBEhn0FdyC2xBciYi1hDj
bwqjSqGoK/HbG3wpJRUqtYSNpcEtjar5kzsZc/Y9tLBG1NvQfzysvstL/M/o+H9q
ah6vUOQJ42Iof85wFLzkpetAwXKdBtycuDx4aj483s9wMNReaSC06L0Rx1d6IuNd
dEG4/ESEnOeFmoowf0HxjEaTTvtid5niJnRt7MyJmu/W1FALPRXdKgEAPCu/JKfC
PWItNoe05o+am6DJeotLwffWbKIUyt/WhZ4lYVmzdgWPVNUNc9IzDaHGYOxQTgTh
LpXIQ2ruZ2EVxg4q/IAeTshhc6LX7y2Xi8+EsD7bV6RYy5l0Q3IWXfmcyLxp5nYX
peToSFkPW5zCkrXLBhMAicEDcZ7L3G7iUPMTHdDpf02f3PpDmzC3z7RkMzK9Ug79
IPdy4jrC2bIyVebQGVvVObPTpfNu9Bt7dNqX7mWm65Y=
//pragma protect end_data_block
//pragma protect digest_block
BRHwpsxlfF1Y6vZXxEdDEYNdBEE=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
TGJAanIHHp8lImKf1B8qXThM9n6jClEAq7Xz5kj4jZIZJEPPNpjl7Bv9NNCFNnDs
R0e3CUOn7QVdOQPo9+fRX6+S7kIL9EXSMgld20G3LmtriduNosFnGhiQBWW2efBE
/2KXU7kTui0KPR5zbEjQ56Qc+esSJaFNT0u30xfU5lTQcJdcC5+3+A==
//pragma protect end_key_block
//pragma protect digest_block
sUg480JoZ52VMh7UWPFwQtuxAR0=
//pragma protect end_digest_block
//pragma protect data_block
Jtohn4p2T1o2+kvd14T1wLCkgYr4fjoHPlmDClHyDdcLYao41ibOAQ/sNrlzEQBw
LTp3t9bvvycd0BOzpU+LINC69rm8DzXCuGlgTWNSNp5Dm8IwW6BPV+um5BMvK/+f
DgwsiLkdwuh4QJL7x6Nzh5JOjNAulliKvpy3U5HWkCItYYxeeT745B5OFdFd7lGp
y9uA0hhYe6wXk/HHjh9aTNIfm1KPcSz6o61EQtP+qHGYDSeVXNHJcjxndUNo31HK
pL5LcU1W5+wu+Rnq6PUI/Z+KgC6nOQCFnEC07Ij8QaSHvqjG2IhcwaXV2lu6vwJD
ttBWuY++V5LBksVdFF7haeRpkAulwOcw7UTaRjEeJhv4h5Om2uG4nuLzOgwXadBc
RODfbleygq9AStH5C0cckg==
//pragma protect end_data_block
//pragma protect digest_block
1E19xdOHPhKbLSlIDei9a/VQLDk=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
IcftBpFoJQ6QwW6ls88TCygkAetmUNWtgMrgAcC9Jn9JZmd9yupphBAD9hzVpIWt
08WQfv1wEjf02BTHHdakUXebBym4QvbV/F4pYiBvI+b6xhvaxrOjmLPlvwjy56E9
30hNz/2MIh33yBoOk1VJ7UAPwSEJPLXwtRQ3Hj2S+d8LkSBR8RwkOA==
//pragma protect end_key_block
//pragma protect digest_block
pJ+TAMY7tGMsLepX4WYQIYeX4uQ=
//pragma protect end_digest_block
//pragma protect data_block
PdQdNAU+QkmNcsTLkkw0djbmjrWzFe6ZyHTrbLJpA84g+ph1HFZJOdira7Bu+Fbm
0/mWORSycPhOl06LLuYZ79lF3CrklRIbUce0zVODe/2F4KDfSY8hNaU6wFBK8wuf
MwIYP0huoSyi08CL3mmDknxV3ZZC8R62GNsCpm2zWIjmnl8QMpgUUnO5s2ZXWQXC
FK5FYdKiDhAFENLuSWxXG2S/qwGb+Af6wn/R5O8O7A+s+B1/H1mQC4Vo2ja95/5I
sxv37qFwl5tYNYsuhZZaUTtGW6c6GuAtVjNexZ7l9qTjuaDYQG+8xJCWhn9NaeIH
neBtTqKOn5Jd9fo7NIAjNaBB2r8x6GAfc3cKAzSxNtCP1BaSFUlozpk00amTI4l4
Rp81q5jDE0BRNurKyX8eMb7joAacHff/0HwowP441JfNs+g5fEmok68i8yKtSs3Z
FJ+C7ud45D4OzazuF8b2iMpvJ5fh9UGVVTN5SLBCXPTByRotYd4NeC5tVy/s7CEV
oHxt11FbA9ywahS666bvC7bfMHYHaN4M5YsD3SrIQymDP2UnAZDaYP5KEWmTzk7T
2svHIPZ1Xv3dViWJo6sHmNOXKamARDk3nrwU8XFIDLzaqgkytDutOY/iH0Q0kS41
zNG3lPRu1jS7T0B2nhxJkFvfr6Y2KHQtgW/Nu8hNKT+9Y4Eyp1UGSM+ttQ6dR9zN
RA6lq77JZzpOughg6pKh3G20Regodt7sgFD2umURMWDAE/6btuZO5njm7AXq9qAA
jjcZp+3F7/kx+fll5cZKrZx10UxYpW96BPB9tUDXrrJZKZ9kfqTM4rXPNu7Xg7dF
rworemP1VfTECb4y9gF+ilN2hVIG+jYJUeQ4ihSuZz6fFtEuuVHgOfmW3gbg8NrV
wk9aKpzSTmtGe/0WL37B2/8gs8jXkN38N2glJASnw7ygKckSrVHSaXrts6az3k9e
Dc5nHVeQpY1eeC9Fs4YQzUBSoGAf15M4m2A4FEPHf/BI34B4huDMJKuVwrtZ4fvH
l2LL+m+fMhmY2Zx/omL4vEe6OMK74mlTlTAwzWjyvhozlVSCC2n/CU5yLn2Hojp9
0cTxVLx+B3TrBtjyOHMETM/O/B7+Wijuu6Uh5aZec/3aK4wZo/Vy0UYx8n3+d6/s
R3wblqOkws6/VMgsgXLrE4kxDQvzsthLBO3NCYCm49bno/H1TSub26FyCwfHjrBU
dqwSvqifhTjEsPPlgihc0OQwM6CdVfqlJL6o7Waw18LrO4Sd04dfxPRonQP1whz5
dmlai2z63fKVoOuL3ACtDcM1/W+ALNXyP9FWeJ6fRHG+PgFczqdjHwIjEjEh2mDe
9vslHHPpv0J7cmrVSZgI865NjTn8+X4EZVfLDVStxNg2vsY6lNZSZS4GADBsS48o
a7zUXLOXwmHuT3x7PA1fNbA/iCr88cn5qZ9o6evFi9bWDr8hsoTN0Kv/R6MZ9Wh7
inXZxbrEsgmO/i4brzDYPm8lHwfeqM5a0GXppEXjqnrWePe4w+mO30PZHU6XqrHo
3mB1g1+Q/0b99LvrHPYYJpsEX/vxvKznUstnvP8sMy7lKvbHci7uOcZQ7xBvzZij
S20L7BafipBG5QWzVDEqxYoX0zHNN7XXYPA+Q6JbPJqlZcP8wFzfNuvNVK7letQx
HKdW+fD3DayeAj1lv15hB4+mcZMLOZhwE+o2JRAqiZRT/4fIyi32vOzSVRRBBkrS
k93rH83Z7i7xmQUSG0TQALq7UlvV+bVNXiEE1wJ1A30Q/eZbcrRLHRIR90VkV1uN
tgZ3VBGrUkw0etOKy/LDxI1jt81vMPXmwlX9lv6uvfWnfhktOkUBhZXyRwMY6LvD
a6yZKePxHXSUGsU9tWJFTGFx/F0JqK76upUfMHB8QC/8IF4JV8lsgMFM2pITPCIv
hWG+p1q01kRoBNTcg3SeGyNTrJwqGsxc+b9lkV2UFQ9r294Wb2TiaAJgmMypqtIw
VOId6AOw9VrYSZP6rSR0LmgtWWEfLMMX4/lRv/GtiaUYtSgoFIdsalNz9S4Btvcz
4JZiiNF0/7NKuSTve2v5pQHrx67iJWuNI0qcd07cNpMKplv1ttpJQIhR9Om6i4n4
dxgIaqo2yeoqsxyl/nIohYlH1rn1RVrMj/MfkW3teLIGeFEIx7lFpHJ+s+GdXgcy
J2hahvxE/uFRV3GKr/qrj55eku/G5mej6OWoVIZkepkt4Yc/rG5ySO0lo8ywyNnH
23hXQ3/rqPrLGUWbZHD4Bdal7Wo5/0IjY5mPL5PEoaOBiwUF0pnx81wmupIGeCf8
kL8rOmaXJhm+xUSQQa0YURpqN1mFfsyexJUWCqzDw69+jlE0rIA+E3dfFb4hFgL6
QjNLdZrEzU7JZ3rqBqvVl0pAQ+NczvXIl8MO7QPQWUXLN7nDHaitrXVvyJX9Iw0C
35kDANcrnm/zgoaYV1xy6F2wwK/0pn1V5CG42FEYdCESQ7wkg5KizGZMbHM/SiLw
VVy8OWe4twMZmv3zs+xJLa8i9eSwKQsvodYmu7O8LupVX5w/wtRfmZs/jvajIzRI
ZyvIIEW9L/R+PUynnhNdZ7ghcjKMu/0njq3/I3I6HruYui/CoocJ8S4i2UwQ0uMZ
bUh5prrGkyT8alRUusQg58ut3YK9cjEq3v2T26Q4Hgjbg3VyTzQEvbd07N5sLqxp
yvwUODp3VE8dLCvh3NGrymzevPKy3SGRRBZECewiAH9kGDKgwU35Ui++A4ei9mvi
A5hw8ud47XeY55XXsCHbQY980CAox+KyEEdTtOd0dMj1NSlHisXXxWa5Cnf5z8jM
FCUS3CPRK/GQlP32+v/LOWsRL/64ZWtVbUSCCTu3y4/v7m7/Cjgm+aY/B7HdrPcD
r5X71mxh9uXRQLGPctrjZ7iD88OwE6VTCJ70s1/Izg7kP+Lam9RT3gFf/Umqi5wo
8I8VNqBPOHBhRsU9RMK7b6Xry7m+Rpk/r6rKqTZsklJ92M2YoPPHFBg2EKZvXW+R
d1aycFa6kOZmtlHkMmdSseUqDsIjoi3AumQ0jhfowFUWj2Q7Vaef6+ldVDE8+C96
7PciSGt5UlB/he0fQsR49KqwWLzyi2PFC41V58P8ICZeOstRwXgZnnZ+ugyMoHlP
xl7rajzBOaF6MPCYJ7ERiKb+BB+YCw8mfrmuNq7dMQLjjBvx3TIhOcaucYLQwE45
UpL2MoCAPHaxER+P8KhQFR/kmlIeXxrkhH0Kevm/63+A8Ia9zN2Zw/rPeWXa9uDf
11f9zaZVNgYxb0HIaeJjbRL1NnFMugMwirgBUdLe4ix8M6rUSJYO+MShJV09kWBF
ov+OgWT/L1GffFtSn7FAFdaC2tmybEtMr/eWh/b1ICLEOMhCrjXXegUO21IyrxsL
HWmOKJUgSfpIHgpDctm8tytOxEB9zLVaLYC33wszlHgKBqn8rP/GcEKywWKcwB12
QVQS2KcY4JvaLKsbTIJLsKxWOSikZkQIex66whkYUhSnp5SJ0u4PvjnF9YO8RReH
Y1YwZq28RTniXnyvmjuoln7oI19tq6T30Gdn1WLLrX0SEwkvIdIu3YJtt31psZa2
tRCb/WZoVbWMtMKMPwCfPGoWRgVnZBpJsUREsUHskMqFmkOqFTwyD2aViyswlsbg
G+F4wC3um+T3xFbSbbFdTukg3NAuY2Ji8/CEUJrc3zrLy2mji+BY5cqaoXIflo0K
fYB0MgmUq0G/mKzfbIMzE+UUFVEi/Dv7kkWPRmT2EJ1ti4s/YsmDvzO9/Z742PQS
aFoELwHEEQhkvtaHkYWb0fMYLVBzuyrJVOp0ZzrBZVsz2l62IqvBSdIxGeBttCxx
6J7uHpWV03F5eBC8fgjm67PbkyEb0e02dFW98SXPqiX/YwR8CMXKcyhPKIt2cJlp
0ty8dZxJQas0PFdf8OdJ6rksd55aDVzipE0Z0i/AdN89+ZVXcXfvGLWgyDNv/iXt
QPdIffj+xTw9RCBIY5aKbFQ4D9vrLeknuh0rSwPwh9dV5JAfS9EfS9ctk3hF+C82
l8j4FXw/wxX9m/jrzwwXT2jKhYhWfTMrAzXaFFYfSVTOKMGc6KRM/PLzNb1RMhU3
aSNDHbmY5gCI3lh6yG39eu9yPQ/KkYgwYRpY4v9kNSPazgc0JUSYmKg1IVODBVL3
4+0aIWHsOs/cGBRimqupkAIJzs6KZGoIwDPlhJ3xhKFgWMQ8e2xUe7/DmRM4Hy34
japXXmShSRoEiY4dZ69RTFGxI3H7HN7EEH0I+XZ04xKY+HWwKaM/8qdSlH4u5Geu
6J03p2ZxnGdMoDJ4YYrCADibR/OdxNkhzgkNo24ki+nq63LlBBnTOF9yWUxqqb6M
e49R79466IZY4rhIOBLiQM5tyZ0xXOX8AYRBbW3QjUDH/AU41bVTCe669Ovaj1lg
MR4r5ZWb2FbpOQgcow/gZnuBlZ8OqsHEm61iKEU8etbmjcFj7henVias9Uc/+cET
SsqFC28CetyJzbrATxpPh+gl+/cF2rG2A+vLsHlY64xxQyuloZL8cu17Tpp0T5Kg
v0x3NN5LHRN1xF2h0Qf7928cZF05Xh3jxnCDHLv2GbN/RW6mHWsTgTN5V2JkS3Ky
drmwNRSVxsKwUtrGRjYZYkAhqBd/nJhUJZHK32+7jYeohRUUsWblw58Lom19NX38
lqkVy0W300gWYGmlv9p2hJt3uPVdELghwi6JrRVVpv/AqD/ZlPKyxjPodKt+eu1z
LkMry4DUvl394HM5axfMYs0bQNsAXUd5d6TUvPxB8Fw6vm44X624ovJUyMjQPMpp
imcudiqAz+zawpsTyQP1GmuOULg6PKn5Jfr/pZw4m3XXFoGO3CuQm4X+HMqdv348
I06XaDdlEKwoJNVpHyeX2NrZDZo3ZLLIkmERIhzFQgJZva+ZfCmKKn4r7j6E5Ej+
U41JWYP8/30nvElI2vAFwg2bxbdPWBq8viv2YMCNxDup2srHqz3CSBDMXOmJdHya
/uesAb2GkOzhlY+1K4j4sEYvyPs2X3uQu5wh9/hwV4DYMUNLzvkBMaQsHr2lI5Kb
VGI3F86D5GYKrUEaiVWFk5F6gTR6MEovWafPmlOBMhktsp1UZ+hJA3uPnyzG8P5N
i2MWmqaSMcJiEAbZP0z86NxNe0NQmOy93Rs6IYzLBWYUx2JNlMEdQAb2WaOkCUkp
+hAg9bjY7Ri+0Nax/0nLPMkMuU3RkY09BtbTCmTpTfgOLwBbVRsFz7o3cohEMAJS
9cwBlwaCGlruhG8+UMhuDpit4hvB/hQNovqaigV7F/yUd9pAzlii1whAAhHPKkE4
EDEf4zZ0sGOVXEi/zMkC5fnE4vKzxEI+E3gVgDqQOFzsj7AOJDjoVed6vUVV3dgE
m5NRR/N09C9fYu8PKWah+b7P+/aZvVOy+aeJXfaofNrvw+h2NjhoYw8IO9hE2IAL
TnFWFbvmd0plfMUPFpniWIGyY2rb+qOPc3dSrXd7Rz0BrLkWG4TNKD9YuYkl5ALf
poh9Fgt+AzYz3CVReEnJNrf6NyA3eETxUAEXkUv20yEftZkZWBiVvcWEysIVeEka
YT/nshVIzR5M9kaQBQZ0BUdU62kjmhk8f/PDopAgo9005UA53IhcoOjGE87A5oQU
qxjasThkQ/9Zp7y/gLWqEsaR34fQxLizTOr24l31z1rBC2Dhb5RE8wp2/s66R3LG
Q0dn61vfzn/OtqrCZn13jnSyl+LdLjB4inftcNTGB0IzES56cc0lE5itnReYn1lu
h7XrB+ZdCN5X2WhKNkCtaQtX0KqSt5m3YqPQr0/kdZW9psAWDLulEmiSiH1SH+BU
rRwpg7ALgo+gz39SkdpFHM/sUBUSt//O8aEEvkv19Jp3jMwoujUHU2s5FX0UBYpJ
tQvOsFIwInSRukS+TvC9LfFHnitlJkHoMLZMBxHydQGnnaGOwMTW0C1QZR9hqPCh
ZvrsOSuiFjyX2im2em0NT6VaYEQNzZ6rPhn57PI37Bsvh0oB+8uPcp84kNuIz6sz
/Cyui2ztRYp4ZBtFMy0gllOOCErtV8rvJ85TYr81lDQrs1HmrSwakGBPcx/aMInd
acqo6ZxKRom5rVI5wQdl7X+58R2A9e0KfM6Jd6amjvqK8yCcDNw4jue7laAhVbSM
hjXIgDgimjhmApQdTUjQrxFDsafrk9wGr6RNnDY6DvqyCJ4qSZy2DH2ZN33jrs4Z
Ajizsrut98+XYfTJowzrqX48P6LByIHneX0u10j7M97MzNJ0vWP9hv6rbcTiJDsi
s84rNNxLFhW1FcHF98ECSVZlXPFBpxDhshRhoXtigr6McufUZFSxG17D24cXEaVN
enQJo5uO6PFYRVvomANkX41rKBCKovOZjg0Hq7r3Iqwk37+KeACQpsvvZFywZtzb
DYrBlZV0Ez6G84u6ZSSYaYWqGy9sJ+BZ7c+r2DDlyjSPQN3MJhXqG+6Dst7UkJMl
cH8owTOUzGBxb+goWilOx+Ij7wLwO9/zVIO7o7wXbXG6ZrrhmQZZNkKdOgsjwbDF
rIU9gcSq7JlNVVjEjeOsYag2hdzCeAfO+L2rcvaiuXwkuHCKiKbd7cZ2D2orCUoA
wLEb+UKzRJDZyDEs4dQuZSLoMqMmTWNa8wFFhZd329vs/7IWsW36LrHZu1AVJf9Z
b2PuOuLDqRmWLciU7dTT/xh+x24iuoQRQxvaF++wvyJkc21Ov0IS6A6ys6UtaLop
iEMaHj9UAAzR+tniHZiRoBAjQPfZi1uG+1OXUdbrc8gc9j1tpgSBxp1l7CGNd2hH
Slqn0rC3fXk3PuZ7Dj3+Kvw1540KWNK5WaKh/NIcolNjaCOwfcKdcqg9Hy9g8Mr2
0iWg9LDKNuRkWogGjLLH2HIFpAmBUGaC7SqjjJGFOTO03QldPeAG+uD71fc+cdhX
dblOVrJ8qDN29VUr+jViUicKRG1AOJRDrQSdv8lLw+y4HxRth7ipdJ4Q4cmQcNiB
b+rZxlFhqRXS9y4bx9pQbYs1lUd2W0Hhp8tuHiS1OT53g1lQZLYaZ3ffo4zamEs0
FVP6TT59C8/U9yuDzsIqNWNc0ZbxkECC5BHfYsIvfa+CN8rtIbkAJPoLt3kH+egl
eGETLPkyA8NAsB35b6qEJ+F3S/kdqICF25qnlUg+ebMaBq2jOaOk7dXEIrhCaiJy
Zw9gYWmCIxGNB/x4l63Yzv2S2zDDfXopu/EBIA+R2iFhByIrUB4zbCj+JXxOQbhJ
y9qF12Q/VyZVYVK44+vsuKfFAq2MIaUtjAgAuPHhtgbS78Mah9beU3GS1gCOUNrL
2ZepGOpZONeUu/UfEcU+2OhAJYzZSTP8ZGduSU17+a/7Y3Xn4nnY4k9A7PaaW1t2
NrmbzImOdDdOYSeDN0vbQRi5UOsxZmLdUStKu3C3KPQdCph16kt84I+DY+VLTLh+
Wf/ASq0+VR8emWogDMwsYo1+/dORYXHZcDxt9D03y6uvc0X8Siy29NVRwxJ87Hpu
hG2E0BO8X0uiVtf8fSE/gGvTnQ/eKRJukNBBULGGX4162MVxa5wdlIPT4urSTV8+
43uSJBg+6PFYo0gRSxIwcSUCnIYn01/ZDrcbnldyTN5qojMHI1kfWN74yP51KmXw
673pPTl9dynE2lKooafHC6Z8uB7qJGKUV6DAIxK6JGHVh0B7xzVmjt2rdt0MIZlP
MdzsMTqT5WAL7T2lKDbZ+M2BJn1BHE/zum13voQqQ/qCJAbDIOS3zFCbbJjG1IUg
hhGHP0RcUe/UU9tJTyZW60NAovlGeWOvj7jzPQHmU7XgqxoJ1JML4jxxEhWQbDCU
sBGXVQwMrXjjgUWshfIWak5v2G37xloC7v9XViF5ESrNa8yu0yn4zq8OBtX1qyK1
R5vWAW+eIU89Zz0i3hu/WEy/uTXVBK50Dn83/ZY9nquQwcLaYxpddD/Wh8o8Ukki
qr6BAD13j+UPMGqASkEJ6NhmVGFrAQaUkMPno76ZfrsW/WOvslbO6SFcDI97T7xc
OYrLHqjgqesIJGzobpMG2uIWfylMHFKOIkdWesMwewM2ixAkyob7dmZC6WbZGllS
0dLAj8AanZGtAhq859epLA5aTSY0wULFPcTW5CJjTpo2HcBkWuEErQsHcXRnZId2
Q+kUgt7UldxvU3bYxm9Jzk09/0v4NPAGnUrZGJ6XnBzm3zy9Pr67kgaHdmJ10CZ6
1dfW+8xL3OZIU84234phWWX74xH87/y3QP5e2uNopqWOHit+3Lsz+jq0x/P/k8ut
QqJfPTv67mCMWd/0wZ4AzTkLh+YNdQzihNzyMODIX4cHhyZJARptVpGmQqOde+yF
iQ5/seSMZxoPc8+oAaNWhhtoxiRJ/k1Dx1J4Ft41Knz+ZpIbnIIEMka/SJhh3+Zl
kru5Ntmp7ByU1Zbr8SSHaBSZZNS+RJAnQIjUL+j79HrEWSPD/9DMVw0rNLR/FD7f
slIe+zQLqF0/krmNAnYzzkTBC+RW/fQ0DX0Vm8TpgS5ASu29Y4vTcxe1kbsLKmlU
g/7DXWhTTCw6/VTQ7ynQEsiNGijVJ7r3MpCYPW1ORrc4XmwpFi+NbzQTi5HtAE9Z
/d2sjrAraDdF8ZC5L1o5Cd/3GYsVsLO9rEDZC77XNPTFX28yVeLfuWtHKRmJY3fn
G+KY/qoDbplkW9CjzctJjzJojF9n8DqUyKDRCi+Yq/M5wtUU8POAYlLrcRg0Wo6q
2j+EKr77Dti84Ioo1PIQbbuuEyWIv7HtfFofRBlwOeR5bIQ+pfiXvtt2/s4ySLec
fj1y1ngIIicjt4JzKse95bgtr1sBjYccsfGpTERhBJ7hWFBNTPEZoCR+hg5Y9sqG
C/W6hsGcWdasc+Pb+xnF4dC3k+H9CymKHI/zgqzBx54BemH8hMe04fQDD++l6Nke
JZ6TXQTmfztOQTJltAOyDHaehQJs2HuQDJ77cQzJs+G9vuw7WZcmSnVAS6GbPIKo
xm99B9hfkMTGrAg2qAu2gGgfYT9cd4NYsKxt2q04U03/rFsL0oxqE7t7j+CC1v/q
+HCYx3k2m0rAgBQIezPnGfkgkrdWH9M0G3QDPOXAKaEqO3KyULjbw/cA9Io5CnFs
D/bSojC3/r/okSBZVnpKw5KuhDGrB0WkkeOoE7egbuefBQ0LwKUFkkCkp8fu2h7u
Vjw/DYLoEG0F61KAZ6UakHc44S2rSRXK8iV32FVb/gE/CF+5RGgV0KZ9jIOkgmgI
G6e4AmsCVZHbrDP9omiOYVUBhorRggyzPZYM/mpw0Fr9XJwcvbS6n0PFiZf6vzRi
3uzrkWckI8y7FreLWZK4AF4Ja1BLcbF3FNkg0vR/bpFSdeMXQiGjQXxP21FcFyS2
OecgnChkNXRKCGo4FZZfsKkjkHRhmc27Nn/PtcTqv99Wm9VFh+jJcrD0hEslevdl
/xJQJ3PAxScYo2r0UgMUx/oHwRPLXfPDgbGQSquemGFWZPIm01bWP2V9k1iN/sMw
2BIrNxxi0+q/WwmBDZDFgcvSTUwhrexQom1b5DlDRR2yNzaTpZYOG8zlmdjXdrpt
tn/LwxlLiFXct1MwSLozTAsv9x2I5YGw6xRjZ4COw8DmuqAHatcRtmc/yHmhhOnP
gcoiu6wT6DnvhRlodyF4Q1UvDwBf8Q/+Ooo0mAA4rrK9knytHoaJjTKjQSMBLicT
zYuceIM7DCuL9uwhEOqhaMuya6piqn4ziyFD39uiant5btLTew0fHO5A2xx2CTRj
j3RcLZDPaNRhM/QcJgWUd7q32eRFJGq8xXQy3p9WZDwd9cXpbtY/IYugnSf38lsT
bA8o40MlBEsH9Emww6zaACxtpvrmQcM/MNt4rDLSX87PsH17YdejhV9jUlBrZjc+
J96y2Xu0H7KufsKZpTfiCHqZn/3x5qf9Pnt9dqXWgNMM3Obh8Jy0rD5fzM/qGeAK
b4+5UbfLnSYXpjOxE8gVyA5GaltFGjOuE9z2FnDLCGkcnu076j56tw7t+f/qenTK
aYxBPjERJpWFN6cOchB9Hpaxre8CHDJvj+792s0hRpXZb4d5PwCy/TwqGhiyeWJF
vwvFUffsNly65y2fucVDKfUTlHjDVig4SUpA424tn1cUR8UHRRmCUcng9wG4LXPb
CtPl8m8cKp4a2wefexz5bzBYZv0ci5M+MfmnreqPdv8e3cFmkVsnKRJFu5W47YHU
nClaUTZziMW3SLnjFWQDCsQrq8G6+Rkh5drhX2uMPsbejNCExvVBO9zhpPwdKodv
vn9CS8FMWVDVFYZfyAjMvHbyOg35n9ZxBox47PlS0Jt390QzVO3qqdiWtymtZCc/
HmH6oCcxUw3NriwynttRbjgH/DOGiAKt9jdfXmyNE/lujxi0aeG3YWxmjnPAaRgs
rBObeEZui9UBI9uSRcJ5lokCWlbqS1kBEuGk7mouorhq99PoX3X8ZGtt0aAh+mWX
tJ+KzNy5g8aBD/dGGdjqKwyFXS78Gzxq3tvsEg9cK2oNpMriHDCIE4OWJTJOlRKc
NQAdpVRipgiA0hpFc1YMne11m67V75YnZrkcMqku87nB715G5tCgE9TlfqeAXC0R
dzkJcsStAI29KSbWHd8d6fvoLfPP0e0Uo7CApS+0Yu7aGYztagaUMKtnKg90IRXP
4bWz7BIHvbG/ILkYjaKk+IXmg2ufxvgk7arPPqMWO5FzHWCK9qOVLoE258BhLdbC
YedOuJeWeGFfV9BUVwpwk5BT0LYOfFV1ZFgtz66u+XLskS7GCIQ00nk0PBBOCSuZ
62ZpSb7lZksLu/AlFuK2DgpDuDYMXXYe/K/cnMT70wTJlzLaPSLIhTck7op7HGbl
up8PFLAefMn2vGQKVGKvtV5CO735F0iaTMiq6SGE0ZC43wcs2I0SsETOj+aj5Bki
A2rJC+XQ9RLs25DtaTQ8GtaYi0a+WGrQo93N0odH3l+WJJ7DEDjPFrfpB9CL3LXn
FqJed2tMwcBu0FPzO2ng+i+OdEg6LD7jiXZf6g0gYOYKDtvkjOtbp39CjIjwmVAw
AHBw4VhkIAhMbO/TGVl3ZUxN6c6XsOTK/6ZcvXA5BS4Bq8hbQjiiN8z/SBvKUPW6
RVwCWvOBs73DDl7WVZp9Fj9Acp2dED0qPJBY3IIVgoXKTsizeHewuWnxj09ZN/rs
Yu//iOr2qYqp4fdnuYGQfi459xV3jjLx3uJUdTAsYKYLi63NoWidkvv0bWK8VwYs
GHJeUnpxrZFeoNjOjRmRAUUjGKBWfa5VGIFepe7qo6tfrovx7sjZWJ8aUqIPd/Dw
F11ViQSYhGLKiKTtp7/cfGnxjZ6N7kukZxovrw/zZ/ojXNNf8UoTA14WlP683wcb
iuOxpSRJoSYGNszbsrO2dY7NgsPYz2B8A98w4lzQXQP9+1pVhsth835w7yu4n6HH
nuYftseN12UNXSu8yVhWGUYtUQffD9pVg+Q1IgYOBT5fVkXmph+MkvLimWdw0jyE
XKZln/CLWZ90rhTmUqJxdIF1vKH31v62B8mHoGl13A270iwI2huTUZeIb3EzmDJn
kZun8absue/Juv1a26N4wHuUOdOxljfQ36galI98Cs/VoXqW1ZiOSWt4NsWth1vK
VVQTuCYFaIKN41m3DMV6UNi+5c2NTAqSxAmYxM4jd80W0ZcCDA0gvE0VBr/KcA7Z
OqAYMigvms5cfLr7mqSPJQprtg9ssClKlZd1rtCrvdYoW47OxofZOWoeQ5QcioiZ
oo403ZfROzWRUrf6fDj/U+PmzzzaVSqV35NMmr/WkybLUBQtvQHmePgiWIXj8Nc4
XIVfo4g/bSQHoJyv/kIRnO2FGWhKoGoOvIE6tb+PdRhE3n2qcS4ZavZx5K7QRjLI
/3TGLs6M3ym5aDEHHCxfu+iHg/ooGdleoWNZWRO08L0z+taXtY8WPwQloqw4w5+R
AyRepV3lCsNLFOXIBqCSCO7oivaWFxbSS+wt+oxYkVIFyLe3ymHo+qmaVLVRj3yC
FoyEl3+aESUBRlMlDn0cpl2U0LFsI3zdmsMxEEypF70Qxr4lSkyQIe94njSWHAxy
TI2+dQM7FErmMBdKTegjqULSOWk0C2HPiUwovXg/4PutFChxl5622zk4TomXUTnL
HHTr82yxBhK+buF3ZULiZ+0F0Wn5HcEbdQzTPraqNq4JFOQ7abD4ZqfnLRr8jZum
ILbQhgOyDPV/fv3pURVQyHxh1lJFuu21GVRty18jCj5dFN5kLRpcgUGAzwtUZNL3
YTHeWEfZcN+q3zOqiJvsSCdNZp6gDzQacbdWcRAGJQzlAU+QZYRKmSUBKFV/P4qC
hWB3Z7Qj5DlqGMZDh2/cJNkAfJQ+d1Mq6tB6WJN072GS2wZR5KyYZzMHdvne//cU
A2mz902nqQNDdlUBA20e5y/+Ar2ZwYkUpun838gIVpPfNRWnB2hxwG8F3x2gn9Wh
O7S77B2a02gXo2ac6rEUMr4cRUtS+2wGhxvJnFRFs+K629o2/X4ew1ZmGolLde3P
uj6JLoCJULm0B+WKrXQmC0cx8hf0Ma9hRYh2TFYykT3y1ke4Jw7vPX1ANQd1AR/b
jQm1HICshrI/fqUshOTOw+M2jJrJyVpXkxFzlnG8fIn/KBDdk7/1HZ5Nd7jGRlLh
QWhIaYYgyLjHxhwF4ZMZrEAC2Z2rl5OnlICNMHQkYL2sB1ZYm2tYRuKqrN/LJIe2
LVpyk0hWRz8NVaZdXXvcerQh2tqljb6w3xGfKecqiPWAKuTZ/5j82faUZiUebEbR
sLoGpmVFxHyi2DEjWyyYle1lUaX8qE6WqRAtIUu0WQoZ5vOzlHOQXKbsN76DIpQj
ABY7CD01ZPNXA+02rMEZrJ6AAN4rJgYF7Fn1J601KMYZZXcEJS2JM+Q7ZO5LAKTi
SRq4BYEqoJpEG1bFNK6sHG6hfWC8N5QJ+UcUdaYlRNTB2+j2c69YhmiT/fMlQmSu
3upf7xOPP1CJ7xZ1krhlxgtIaOhEZ9E/sbgs8HmNPNJorWPkP3qeAndWYxXUxNLG
m8PygEMHfm4CyU2ybHOB1Rd4UEIZufk937isODxMpWDc7tRGcPnhzZsS7pr1tlZO
tN3X+6Emj1Vp2h8wPn0r1KLVHHXC4l2V7FSA3yn0yxgPlz3G+jHKOh45ZOxgno4b
eatAtRM7fDOUxl5OHdxRcTQ05M7ptteC6hJZiyRaNV8u14ZogQd4YfaiMuP34hut
a7Exi9UxUcUhnRwINbr/IAQW4zKxPcsi6wFjeBW3gqrUOJhs0t31tqILAnY8hvDB
sh9azmgnGEOz8Y2doSIcKzeS8+W1UdLmMqeOblSgM1uxBY9WZFaFSBV/tGnxUDrO
WNeSDZRtn2knQSA2l6SY23gfPc1+rLtJtri/Haur7Q5jvum8sk7YHeebVTV4wGCE
FHQHD1WGglB9nDUgTgtoqYf6CgjSrXur/AoLqivR7vxuvq6ZAZcQ4X8GcWr2abmx
3n+0MXj3WE1Ko7W5O+3WWWG9umfUR5pagTXh3mdvS0pQx4qbjrXTuIboCU0ipx9L
ceVcvi5lrG1GsVZtxqKJh9Yx2AfJl8puFy/cwDLBF4nyPklJbQQdZYYbcb084XAS
obCWhiKCNUBTQ+iWorXiMSc8C33e+v3HpLlnZ1Ayp9NZy5x1ZJJjKLZJqBEj4tyO
wjPNjvZYT2KG+7X76713RBBkEVPdhHLKbqwaqxl2SpGAzLFkzYYVpq4Uv6Gm92GP
zFDIW1aCU0eZn49ndGifm4q5NIbdUTpHCOcskfWYMP5L3blD5nM2g9/ioQKA+Lg9
9B4g+1mgxf81Qwy4Ho10One+fqcsCZRxdVQ1zLBuKMtEmi8uLCZEj5WgPdYhEAKP
fgwTWNZJlv/7waIl/6OFR8RRiiEaYyddKA1c5b6pSWcqFXmwBd+P0vOFQLW30lR0
zA7EDIvaavuQsdapEX808nAmhj/cycmTuLDDZi7xIkXllej4YIECl3GtAbs5XABR
hQie1jF6kBk7m1xfzLBA+nElp9Vkl05/gxsYXmXUcb9HpiQ9lVNS1golNp8O9dON
mMeHhF62I4wAIdmPY66KrOaMPAxA86aYDmwi/DMM5tJeQ0gh37pzneJM8NwvG2JW
R7K7XhOMQ02Zl8e/8d5NYdDKcxYBZyCpb1dR0EfrsWxEVlkr/8Vi0igE9aI0Ku0l
y94DOVUl3mKq/MfzGU0JRZDcdEa99pywqm3srIZLerEbNF90bLNEf78YDBLOyOSQ
pXc6d6me1pArIyOG5Se/vI+gQxkl02igPc3mBHF3CNqYvwK4v22H2DTuIX0LIUMs
qCgwZ0fCLQITXGDabrtDlFO/5ElbdULrKR0MRCokP+4Yzezy6Y0H33xIeXebQI6s
0KvNvG0IUyO8G/ccSjJZpj+JWvcBlh2MY9CTzEzjUB0EOafS4Id2be6k+4v39zrt
fvV8mk/e2ZqAbI/j7KBlxdKr8CsTMdnoKgZ9mpYC9kRTZWnfdP0dFm54XKVDtV2K
5dt9WOBtMF2Ck1NYF+WEvVwQ4IcmluTgbPXc6rt0lC+PpLO9k0gP7pISj8sipZBF
H7+1s0ARXLfXcwT2+eUmPvKk4LaIXB2YhLiarRzsqv1WXvaZu+qpJygriNH61s9p
0LivRKaWh5Bq+LLdKXM2pcNRKEDSxgZPnwXiRPr1b92NmpNQkwOhQx8lnyrBSlTD
zH79bFhEq5CsL4/t5eZ7Jyo1KfLuCj7FGp7Ex0nocCO7jEU9Q1pNU5GBeiWsraxq
BgksD1yIEkulIFeULREICkizHB0l3+QfDkxvjB0j7CDNZAEbo/mTG5/IhnGfpr8r
VxUcywa4VMnQuac5OiEcvp3xridPk1t8PufV/B2KDDkoV46j5W5k2Q7I2v4BuhM2
iCK0dqXktYIDN2CejGhIa0h/xFm9tt29qYHxKF+VtUenwBuQLgZrwi+uu/4GVP9g
mNZvv4VwQZfnVtmKdeWVUce3/btdbuJN5rcdmReTKwfWxk88OcgI+pFhvWXShPdV
iJLNB1uV65HQvWGaKwzOpxgnxNwWRftXFMg3ZbEjPWq2qB0nD9HWGiEg3yL+skHN
LXngbaLBRbhABcQNeKJxLMu5loJL8s8PxzmCOLi5VgDWmudmPQobMDLzD1dtj582
FHn91BFy5pzOXgLI1qV8gkT0S9wo+xGvAJrcp6l4ypWZox4lCEB6mHLnqiXPRucg
KbkRT6BaNFDciiN4SXP8zDBJKyBIv4sLqjd44uRdA2omNdrGF30beW523ZeczF0e
8XSeRYmbXnk3/dEuDBe0rdSQSJcE3O5AO6GayAiFZawmnC6Nx1P6AtwjEjEQBDQf
sjpLD6BK6o4ASBsNJBBA86DaXGc0yN9bzda+0Yf0BjHsuzkGnpJ8oOp63yUDiUMs
O1XKQ28PZw6w4ikou46DZzOOLQQu33aE79Q6OGhl8sroPd3eAhQ7h5jiAk8WhdSy
cFC/CwouaKASPPDmbCSdSw/Ytm+D4qKMZAQfTE/kGlqmgigJrmeaPVIr0D81fNFt
BQpIIfENhe20FLZYT8CFbe0dl/LcVrDKabdyDIstav+bbguLgNrWBgwZi1u+QLti
1DUp9We5vWQrqZwwVk5FWquwR71L9rw7LElW02l9+gy5/gC2AaRXnh55+wB0I8fO
q6galwvJYsPEZ2Fom5N7QFIXLV6EUpSSgH64cMNpHOi/F32/AtKXKi5/CNTbzxB5
EhH9ASVWk3iJMibFtCGpZO+AzjBjbevP8TY/mVdj6WFitl/+pNS7QUl1h0yG/4HN
vG54wTBlFq0LO1Gtm5LYFU3talSI67Bmc9gc4IA7fMlE9ScZbwrDJzZAv9OG6KSj
hCHXmSn6hSswup1rJNHksuM3DA1JL5njULSIBgAxj/yTdvJtp9FES1qv+36dl+ZI
LS7f1zak1uMV52nXlInyyXerrXKtiGc3zfs9+T/8RWQEUfcKBqVkU17k4VIjVhLK
bRw9asBobuquqQZ+oTdEqOPJmbsC8nP8pIEnXuEU9TY4ldRHbt4ToMeYf3pK0Ss9
Mdex/dW/kW54BTQeiVsRYBvEzCZd3FPNVdCUIq6VsIxHWNXT5aY/B0ZhwN/7dWhx
igwq98DJI0vpp6k3iaJCjFklT7ke+WBHdC/Mu0sfpmwdISoAW8szJf0IkNTsiWSU
PB0K5xEXXOeq+ugGZUCO0NXEsZs8BvZSOgvm9T0Y1uIU4l3/sYsN0a1oOEEOaF53
AaHdFID+syuWZQ5StpJh0Ji/JUiOYYdIR1ZW+Kl14EVqK4TX3SMCOaKm/mUSKL05
UyyiKVPGya9xlo5C4dv7etJNcLwkVKPnSgPoFbG154eSagshwwVs59vxNgVpwp8T
shdzK8SHmjiyiJSPdm2R9oU9Bw71IAXHQQDQSIqrcKAXcd5ouxM9muZO0EzNYzff
B283fHLk4tp/e2P+vSrr77GjlSyb/Zh84o46oxfqYtiJlL/Y/yvTqhLcfCARc5Fe
d81Hz6MHoa4rBNh9IXAJQ69Spj0/4nC99mjIAoxOuy6q7AO9f59A3zQuYUxQ215V
KlcZSrtVrERfwJLIZedJBu+E3wdQ54pdUZGSzee/lbgb3n8cmzZNtKbULyJqh9tb
XjSDpt+0GQKfgVFCwdrhh8AXPeWqBjIn6Mk5Qps3dcYqwjX/AYDbrgp/Ed8gFJbO
XOEyQBj18kEpC+CEtghOhgJDFObQcfCuaSDc06L8aMh27obLrP+riZFMu5rI2Pc/
XXOwbHf/XiKyzPYEvVKzbUiLsWsEXDalGbB39/STDpPC8SD6xym6TJ7ld2s6sNoH
+ocEHEDd9gCJmwNCHDpxmueP5e1VFHW/ESfB/6hOFI0=
//pragma protect end_data_block
//pragma protect digest_block
PVYN2Q2XMPeFQctXoXABqazHHU4=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
meRAHuelRECGKmQdOMkC2aJkBz3DwuRvZUnvSLumTjdrQB/L+ABvr7JqRG/KVkfV
hvD+vW8Jsu98GpweNgu//QPa6vg5cJtPXm0oPXEwARG0mhI9PbscIPBy8yo8plno
WyREf8rtuioGbpifbgKrxYWpNf+sa/sdEUoM3uzYDB2HjghMxXKhZg==
//pragma protect end_key_block
//pragma protect digest_block
SrjS/fqyG9pH3tbsnsoZEkCTvjQ=
//pragma protect end_digest_block
//pragma protect data_block
c8a05XT3xzVotDhumTcegz2/sayYpUQMi0oGQVhTC/G+yiZYhl85KyK0gU6WJP8k
hstQrp7qd6YNJo8n9lRiB7x/gfcKAlDYI/hvm67xYy7Twc19Qb+8p31qiMFe9BK1
utm3k4/SnkhkXhM6+zi3xp4VJxxGT8gtZPAKwTZFjbEQvoinHcdBQ4mZEd/5yR0u
5FETg3GaCCcE3k0LCqwdOmx7QrCBc+HTC8Uqb8DAagvDEeDNBilWdjAWHGuNJBxA
rT5l17f1nWsd+uymFTF9zgEkKDmLLdUtuMEsEq7bLwVxiXhrFI3CMk5eIqolZvH9
rVNlRl0GGdSQEJy5bqu8s+gswSUVpHdwFBQrQP7QlAjEETiA381ojbwqiQrXg5LL
cgipebQsE/5zWL0wBgeSTVZ5eeoo8oDpnqkHXb1J9tr8qnodied+pLTxw9Pik3dw
GjHNm7NdeYSQtw48mgSDm1UJnD2lWR1pm5ONXQVZdqniMjIgffwYOaHddlaj9CDM
vMF8LA57jrhBoiJ1zoqXYDV7UjCHZrP0Qd5g8i9jtNyIihVWNSDlDEFtbt2KU5iu
r5Cwnrm7I8c6yCxo/v55u8UZnnFiUg9iQEAnD2lVnYPU+ZJdx9juO3aPq41zW03K
FXzA28qJywjY3BGhwKaRC1NLY+3oJxC4z5R5oiWfTl8AzV3VrUL7MPJyjPrcgcyo

//pragma protect end_data_block
//pragma protect digest_block
8GyY483TT2tCAB/OA4oOP2v8Kr4=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
/E9j5UDq8mVMnZ065Xo+g7UPV5cRJqW7aCo4e63WLNz6q27pZ4fzDxTrY+DknW7y
DKJmYPsda2gt02V0Wi6zjYpNKLCIWY4dhU+W83AGfEFgN8E4Dh8aamuJ+o6+hvnf
d9Rq8cPyLa1+Iw2JEdm8e5abi9UegqXGUFJ+pfrmWBu0RrBeazvh3A==
//pragma protect end_key_block
//pragma protect digest_block
okOuPPn7ArDLLspMCJJSzkIQNAM=
//pragma protect end_digest_block
//pragma protect data_block
1/uDHrdw9r6XdMQ30MavgxfeZHJVsUsxqaucq7CT+I9YfUl9ZqmVoyT80cJ4aEZ8
ESWRP99BpOcjfeEPqBCoZvWt0yJWt9iRwM0rtOxB4cApD52TeiW4Bzf3i6JdSdqH
7eVVZukfE4WjnuDUX02B9vLgEC0umXje6q7z+di2YQ0Ue9vIiaJdgKFwJTUUL+ci
ljhJQNI1iqx026tik+AmC4seCmLm6xgITNwdy2Jntlx5r+JvRu4VANXiKkaKzjGv
HOeFNqjwx8tnUX5+EVr2LkZ4QVTzmqkGZFu7hJ+NNk4q48RNmrAyNcO520y8DLQn
b1yC0uoS33shDQOQUViE7FKwbR+lo5u5mIo52Ds7COBXSNV7fsJeYwcJc5/hbh9b
uaomrynDBy4ApkwEKz0DX/SPfk3VqntZyMWSDYEPzyRUKtoPO5+3NFM9pbmDYfjI
d4iMhhyOaPd0/bfCU15XS6djFYbmYWMMtOwtQoSMUpBmchAm8PrJPP321fQbMKdU
DqHIhI8aU0FHUMonzPfesYi0t9Ua1RhwVRLx/UKHbRJYqpQcM8/THB4ZEAcede/h
nXNT5/12owlLf0sehZFdi3DJULs56pj9fyCyxTYDLipegDdzqcAmt9Yc/2X44YUI
TT+z+POvTZKer70y/Tg58lUXi28XXtt6m7sTj9NdzfuvSw727aUq+i0Spd8GIRIW
k/3SqmK5QyVLJ9wgCNXp8qJKhS5b3USfZjU5DCcrqNBiDKA2LjHp38z0jUU9rZoq
Gw5dPUwo3MisuNZTj5eQb02X/NXbVgCzM5xO5+E7ggtqSH70CFwAKCNfNoAHDseW
VQykgz83gl0pNZjpXhcWJWbIuIx9bt0vUYttP5JkwbfKLdgUIXAAIASr+5sQyAt6
u7+wBVGXUOMjFjR+YHeBbOUIkpwtzup5eaK+o6R/ofoL73zbOXiYrh0JSjII2k/h
QZRhQXrl1/+HDoeP5wFBnIEUJCRn230vUw6N4Q/iPDX+UbTs5xz6XLNA3PMIpbaM
tGOZKOs41Y9UwpYn8zdH3PGOFQtgs0Z+TuFSuNq6QRSTklOjA8IbgHunR0rJDqeM
gcJd7i0shgOPfHehz9oNlIKukRTH3mFHDX6TwIBh7/ngEyFu/AhfsLnrLrhrLbCl
7UDqaEX55u6R9FoY33BtWGUh5AbREycLsDz8MfFWUFUDZoQAo1NZTyPvnd+aVAtH
mXSPSqbx8L5es/vThNUJdTQPv0t4CLio+k8FNt08NBJp5uWv6AhZlIFGulxgRA7F
HC0ELPmdjfbxL/psxyAzCbKFfU1VNKwkAReJladDOFlZcgORSvjhiOMPsjWpdNKE
yP6/VoLjfhaa75pVZk18L085kevltuttb5AOaX15h/11zrzhDT8AiUMSmoOvRUge
32x70dheNJ5x89cp6Frat0mOCQMWoiq5IyfF5RP/wiSY6BV8wIGObK3GghMMzcgg
fm2v7gjj/2gvv5/N+/NQY3MNpK+FcvPUc3orXzqbl3vyXn+Eu7sQW+UYS6AuhMb8
z/oSAnrl6nBR3ugAA6beORPLlUHcFb0MOkURXkLwIyw2p0rzdcNJNtqsXRACMyGp
M8k9Z24A/54xH6EUdrYSAD/14vJOlJBzekIIVgafMpbqrZkzCOPguy0iLtf3LFaH
Uzxt2nJTn+R53SoNwV3366nFA1B0zphU1vyl+T5MeAvaNpr6o6QALldA5NGsdtiR
1a4apy1ppIsxmZMWDrcZG5JhLaX3SYp1beFdAMyrSrrw+XwW5sWOa5X5P9SAgRpv
4J70uhBkTqV2ZbRVUSxEDn0yMu5KmO3H5IAl/wXceAV8b2Ftt0gnZnoYUfScpC2S
oqLhC5ILzj1y/PcqSB9amC+KSpVXnx8GqvmFJKrfWL3hDGeGgvBs1pk3BgtV39MB
QE9hr9aMNDptwvnGhKCP3/ATsdv4Wk8YD0EOIa2ADg9RQNeI6hDvdqEm09iqLdmw
ISU9dOhFa9zUGRj5ziN53Gzbg+ofMtfCiho6KarDlO8Wl5SmQ2VG4kN+Qq1NGyjA
8ed92Y4PFa0V6hx0ZvfpN5zqeowTgSs9q7mg2lWxWnDkduISNjRdiQ0OjNB449vS
OEIhbK6IYRQMfum9nRIqlrtKKMo+NQFLdst7M8YS75/Tp4zEW7L5uQUiiYARhmFC
Rld+tsEQnQEzxndqcVWjFt8A/uLt/ivButHt1/ENFToLidncfubAQuBVcthKkU29
15osPq6CHxiz+uORCdWnBCHW85hW8rRPfLPGTUjEev/U34tYRsM0O4Ow1GDINbCy
yY/YVHRalORKLDD3kXAriUpsFo7oLs4VidFS17uzyh/JCYV0CIJ0qeoI/LOYOxyJ
rqYnRkfYbNlE74KH/8HFmQE3xPm01mpR/Zh2y53/3BlsCxOOSowSWP9ba71wTZG2
ZmrfUnNjuI0Ypchwa0KYMZxEB9eX4HS0vdgrKiiJ34uND6HqnItM2meF14AQA3ly
iXyygIH4cW1AC5x7FnOPybztdJaiacCPb0Nr4ZfklibNemUovb8Ns3YkYpsydz/K
EbT680H246/zJVpucTuly8lJnjS3lfbmP62P1i6X5TLw2g3AOn/xaMVoMqLWl3EJ
7Ed9UXDxcl7mtFmxmvmIvGl3DAi4h5RDOQpAw7h6TeIlia5ClY1iznF4J0yivvrk
Ci8dcX3EBMK6DLq/fKfKNtTIvxRn8TPjNaNXU4c07GeM1yxJp/cZo6OOWV6gk+rI
NM8WrCQmlZtzMAuaTfOUi8p+vha42oFIYOJpJ66YaxQvV+yVb6MOAHaekmTyq0GF
hbPTn0BtVPujeaT1utcLPR5v4eO6LSMxUeJTizVk6/usjzrCL+1eZL2Y74qwUiqu
I457/0Ij+Zdb6QKIlqoMTzyDc5V5wNUt48i/fqQYA/NdgllXU4txadV723JB3vi+
UakKjFdLxkO8TZ8lcyIqrpCoVkzbJuUvdQEk4OBITYe5ZLLxzPAadIKfKXN+XquZ
aALhb8sSjD7RI6lKBgN1As/GHbyHXXj89X68HZBv+D6jPc0XLNgG2wvNlWq8UCkP
hn54w43Sxg2TzSmCYRd43GBG8GIa3+6YJss80WokUQMapbgLZfG1nE5dfc+UQDpA
t0I3Gx/8PGrvn9LuSKYPWJCGZRseWkWr8iLL5hvVbH0WnZSDAnVkuUoTLqkSpbCT
2ZUdv9BuZ0wZFOBuqz9cw+tkTnO2OxdlwZj/PHPuQCjoCS9tHDjSUsYOcL6I5w93
X3FATGqS3bkjWzOwXr8mlyLYgBjTVr4xpwzGJStZBWmBwZMhX8rco3D2PPhJ6tEp
oH5DbDI7VG96QaFit/VA4JKHm+q32F6nmOWqMSWW6HUEyHk+pabui2/x19FWPTyP
3E41tLyB1yjsBmr28CVJxSUxMcuNd633bVndr/4h+kW1gn9BNP+P99kD62QRkA+w
QGymza1Fg/nGb96tE/+Orup4Q42bK4w861EvfThJIaS9t2NM78UK5d2/jh0pAMAZ
taia0xmQ5tzSxBFvodcr36/O0NsxYND3WUhbP6AmQtk5yVTDos2SafCi0tzOCh/q
8pUx/0fgAEbUBh0fXOdFEnKH4xniY6sKKFjxmXDcFKedcT8oRqXWAlupWsdcHKtd
evygj6eSTFVfWJPFCInYfqqX/Ti1teWrgcO/P8GMFb8P5hF9O0Ahr4Sr1s0/ZebE
L/5wX+N+YQq6M1M4Q9arV4ulIfMdHj1X+/KrYJxnGFxhJRfXRomYrWYwScpXD4Zv
dOrY7qKop8jJIhrTNoTN6GIq93FtR1mjeY2TwhQKtSmTeVwa9BhjQyNP1sce1SF7
CpCdBqMuXHw3xssxdGrBtiaBXEtEUJpWqRxz0D29FBBcvLLqzU/lqkB6WydSLIxF
vENCclZ5wxUDmM10BKY+irPR6aA8TIccnnz2Y2l4cya4PYDnYjDxPva60e+dUtkJ
G1nZ5pYBR4QVsQAapByZzqx5ug2dZ2+h8+yfzoE20IHZsMaeDEFVYJBG19/M/3X5
mGXjIWWst/Bo3/wPl1WnX8JcexfU/16/554raRe4ZmD+DjLLaKTBDs9tb6FppqMl
ucajnrxgIS1+UGFBpFSNo0eKZth0CrMJmytUk+l37UDvyv5vgNEla4DAydaK2dm6
+BMEqgJimslhzb+O1iMSW1kwzSvXOEvIHODrIeiPogvxCVTe6Vu2ZPEeusI8No61
fQBoyg8B7ICNC4SfgjLHVUglUlXMDwaTstOBDoGK8hKx60wIBbzhkh3ovRaYILY7
0fChcyzyYf99Ii9xOiXOedqCH5z6XkEqZ4V15aoCpNoXDUfwc2Mid7AgvXoBReSf
jotAN+YTIymXw5DBL/R90eA9uK2hu6Ql34Gni3e0a9FnbqSVCbvv7JaFHAFcG4zE
c55Qeyv5KoXaiKavx/sKnbes9hPiEnm01zmCNrbK8D1V1wKaagUcynk9XEAgJkqd
KU9srPJTG5R0IeBGpz3esB/wor2O1DuwKDbyZ03BQKZbaD1W4SoGcAee0OtOIz0R
3gOT3KHixhszitFgVpNndp1KJ35foKe5m1GrmUUZ6zrX5JA4KkvNOpSLHykBMnYT
Ky7fuGD2tSXk+oc35Wy9KcvlBSymhg2PeMNV6x2otI4iE42cMaLh+y5XNzPajeL7
XX5aR3pn77uZ1z8GFHeFk726HVPXaQm5jFQo5IDcy7TkyDg5zoRePNBx5WbOZHqn
J5fsviLkS/2NiNL6lWs/cyDB/0raZ002AO3Jfcr+v5DdkCFmPprovVvEO6i2k1gr
ZVxe+gYZRkdPSKJe8NWXk6Q1UtZHQOpwh5YU0GuatTJgKVlAE69bBKjGRO3SAEJg
8Ccu/AhaLxNRZgvc3csz/ng+ahvsCmWzJ5Q/r5Aug9KeFAqEOvEJkqeGMcKSvyea
YynKiLMGdNDbKp2Sy3k+tOEAmMyPWCNciZ0kQHTU++LU6n71gA9neTmLmGpyHSMx
yo2Syx+FnrB23lPnl9bRI5pY03i0F8TTWHjtJdx/kKiEM6Falaq3pry3lGObaufU
3Q3brFOOZVTkJSWAyH1j3/TKtt3faDrISP/uoGqDmoIzOhuV3u464z02pNIjxAhi
7tizxAAqLDJrDcJHplANgyp7k54mSkHwMLJ4cLTl67CQnNBT3dYd3ONhtzSCblaP
TcDEPh3rlC4GafXjnsfH2RZFUGiWgEw78fAA+p464ttQPWiPFSHkKw9VmoSDVk9j
M5xMRHtf0qCuPD54fPUnMYubldJG4f9zcmu9AYncePlU1YR1Cbqr+bpqjUfuHvLQ
Ca9LZTwNFiF9aQ5QGlTlsqvlB2yxNzbopWo9fB71YI7XzCBmyU752A9tXrdeSygf
dI6bvS4BoExnlFBegU/KWx23vYzagUHS5lFZPLktJugSycbWKRKxAqV172Vj8SqV
eHIbdsnCMPn/Llt1FeOVzye/mSMKGW3Ovy//WOdVRnbNJiw/DkFsA8Yl+QnR9AEV
lipn27dKSTo4b8n9POHnzDfQYE9SP+PllSr3v3gT7VAlAVjTGzix3heJII6ghU+l
0DSgPK9ymS1JzHHR5v3t0QVdzTrAi9OA7fdKPtuxwiM0sHwcEge6LxWTgviKcL2s
ayAVkd5ieZLbLoZ5tYFIcjLqhDzbb4rOQ3zaBCzO18u7l9fCeHPaadKcVQnBGRbr
PG8Wwkpo+FjkOmXShex3NLnsgQkb+y0xAu9AeBq16YRTz/hW8LTCEsPD4Eop7yix
VH9NeX6ohTLJnHBwWnSCAX8rvPO75JucfSJqP8twz9BfBC5p4XAItjbEiC8J2SOB
ux5MBA+LAjnTaY2W440PTYf7lmrK1Ibv+dp8OtKa9yvWZ8aQNTMaWr1d8OTRrriI
hLUcqVqAHiEp00rOltchIDodL14QcNdXusWMk5tALsuuJoc4Mc0B1g3O+F92p+la
EFnVV+1sff/gVYDKsVjrDLMiLaGlo8zwSrBzm57C7JzWgfM0ab3A9nb8u1l1BtQx
8yrp4MaDaHtLuCGXSV1FGJYL0cAABOJ/48Rsb+6cpBMYDkA7lN+8Q4nn2i/QIaPr
qpMLNgWyL2IYf/K4pBqiPyevazlWl1ovy1qRxmvMSDP0T+iciPr9EYa6Y3E8IkaJ
aAhBZubOqZ7x0dEVN61fmtwakS4wHGufwCbh0pxCuvjvPLW7EjsIVpVeep2Eu1tb
UMlKNJS1omtwE7/45gYKIL2SY8xlLEapc2WDfBsRquot9E3ltyKwBLGBGfyei8mT
DGlbUO5vJMVhiMsoFYWfZUUJJbnA7OUOHSbTltmNjZxQ9RiFcNoPrJd5rlv89PVm
4NXKik8R2aH6Z9LuFsA06xA4RdgPeHiyBkn3f5cxazJ2zOdtxhgz3FOlwLkC72Fx
Cw6v+jlc0M16IBqF6vowESnqHSMi0AN342sCMrRXgcrtyySCzbsC5xf+11zTKWqm
Vl71+dZ9pn2mg4BaS59K0bf/+2+CL5hwMR8BLmJv2vNq+gVU2OuPy/RtstMFss+0
GTLDrs9e0hpeMIC51tgS9ktnQZOJw5oj0Yh0liLZpYw5/P7uoZNeYIJRdbq+l7Kh
mje+84yywwLfWrpsEgzmghiviF0Jk1NKmzoZTjsY4ep/1KfsLGsH7irHTpiaZyY0
ZcIBQ94TzpUJX4eoK+cbKoyC8W0eq0mEWIeMTZkq4TwCYJg9HFwPDE6fi7+8kL7x
e4tqv6EIvs1/jLeuROTkd1jPqNxMnldzanIlESn0d3W5qeXAW8YIEI2EZwdJ4o+3
hIEnGH5MfsxoYg6IqkJQJHyYj7oV/OUTltOK4QJHtZx0rcCttY2mNY6kWD7Uao+p
VYfkrvaW31BRdKUBWS/lBBqUgFdRu9eDN+33dz0erfQHMSlouW8ApX94xGQLZoP2
rbYdFW1qBDAaI5N/wiuC2HWeKhHhBGLTj3belQIke30OEjjnUBENtq1zPmDNI45r
0DX4fzW5rD2Dh0d0pBVbv9Hp5xqeUe8fRpUSVG/FTvU6MNZpeJdxJVPixS0kOR81
1/nuAp44XYYUcRCnY/hUHX/MEnqXiXOePS3N3QZdokmM9ft9O9t5K4c2/IPOdu+d
hZ0o9tXZ0njyhNrT7czGAFCqBMnspW52CQNBEAT4Ntg16WX4n0s+P7bBsyZ5X7ij
KRcfU+8CoXVIaZVuhKJK0moJPV8K+HItqT+LOeym6Nzl1V62xI+pbCGnWXG6COsp
b9gGK/dFV4ym4jMN47fsVXZ8EiYddQkZQr+WNX8KJLL288ZRilJ/vmnoVdKJ3C20
7Fd9C4bLMVaJjDXvjN69hC+XuSUQz+GJz1pu73gu8GSqjChuLDNDhl/V+HjlizGz
l1Qn7eGspmKLz/unHFifVfPGRXpgTY/3QTT2ji+PHfQLhaX4z40WPxwzhd6LxNhG
teWcTMFidOgHTNKZT2dA6XOUIDeOA7YkJ/DNESy2BPjGjpMyA0Wy1vGdMjreP8J8
Gx87kS0FZgKFfqm1nlIckkAAFsA0F/YALhqmrWGQLJ6WQ6jJKQns8yeaPaezhpHi
JbBH1x5dHpfnxHpIg+hvUma4pHHA0QGhuhzCA0frfrdS+x/4hoOL3en/kowhKvtm
hhfe008xltWF4cAELmawl/HonAvhb4pic34qkUy8aSHFLtc90NX0gLu+cS8DG+Se
pmJlEptLirdrs/iN5A1gjletmx/jbb5ZD6+9Ys62PO54hLqIzWulxj+5ssC0vR6H
zmrkI9RD2Rka1LXDQYxe8j1iUbm5fYPI3D2nVPx4jiAWd0IcsBkUGetn+AIpPQLS
CGOuNugptybqB4+AX4o3D0kTfdSnGVKUNIT96GIO+PZAh6urQc+C7o/mMA6LWadP
uxfTsq8UzE1gYX6Y6OZ6PQPys3tVuH45GFX4a0YrMOPEf1RwTyGt15g5yvUWV+Db
zZ7AcLfR74XfTU8yrY6QjuzAlos0vZeBauJf652s091RMeALhXGWhx1vE9Acq3Ub
cM8Fcbm0q1IXXOwZvnhof6oqHXHfA60wX6i2+OnWDHtmy2E3ZNOSb/v3yx2eSW+i
M3Rs3VmWtfnZxTy65rqr6SaXiAeAKnWIJlEdsCrFrmHZF8o48IUvlZaZ3DG0rcJR
QGfCij8iPVP5YqDo3lEl8jaDN4Rluau7aVRLWuun9i8dt94lynA+rqZdGLwg9F9y
09U7leK/66unAk8tzwhEkrn9ieYaS8A2QDL/+aDZqtxbwAUoEYwU2tbSANIfANnm
hsEjTxzHngJfU2QC9ITZR1Qyb0sMN3jsdEIEx9BQpztR/X/VPHlpF1Fp91kW6jxw
3e8hfMbg3mC6cqEUrCMIeMqR602EvjMMv5F8qpiCNDkFNJ0PadxuuQzymdk/w+p3
KfHiWbNAAjF9u4qgru87PZMesaaX2Uvbt4eA5XCfoolFmTAkc8fCoHdUSD3X1snF
5LqiVCzec9eRAXJuM1ek2vT1frha++StOUrqby24oZnAiWDp9cnIAuL113y7Niyf
/n/iKOuzl0b3dz5sbey7z0dWNarPyT2CX17EQsMprWdqM/NjYUxnj1xWreiBFsTG
jmXwQXsviEnmpqLQ5eDrU/27wwfCduG/q8cNCErTX4W2Jvl4iBnNVJVF2xA6Pu8f
SutmKu24c+bDwx/elLW7hl8L1yzB+QySWY48+UtLzmr4ivX3sx7vSoJoVqzyPOtO
+1Too2zZa2i97PRm8s/vsHDJONHtESDRX+FWS6I16wQTAjEdPaI0x5tWCLuXipjS
qCEIVIw1VTQfX5GMSsoY9puZtOdYBSGj44Em+NJwbBk7+YM1wpGEqIOezmF9R8Tp
zfKwrS2fJFMgC7knI0zLM1GSMWRXQvN2UeNUOYd5dGK4y/V2dbNt3ASJQNaw0d3O
almODh1GQBWHhx2IT/+zZTSx2GIfua0b8m4Qlht3WOqxr7WYhtIs06/bY4gh/JJe
JqZ1eMJQ8vAzui8Wt71vqZ2+FWXwqUwd9E9Hg2l9jXcuoqwGX08IvjTsLcK4n2I8
1rgW+xiONvX+Y6ToSvskM6NhP6/fQ4E3bC7wd65pokLSbU/mMvCcJEjUw11iX4rQ
ZEVfE6DdC7rlF+7sa2HhMTuXRdQYn1X7lr93PCCoBL1X+SBMPLKumguZaHjNAZlO
mw3G38Uh6Kuxo1QPH3WJD7UlvdoRfG6S/ocXsCyaHuv8uId1nlgd/TDzhlK+ZUcR
4US8zGVcNtoy9Vf9tklLdj9YC603cvrLtBTbJ0sT4M/3TNuDppWRecSnYdsF4Fi7
s0N7adzvMbyroOTeDLsnnYHf5uo+E0wouURhjKU87swhZkFt/jBrHO9P8zBayrf5
2AevVIaR4pSGdroDoLIF9nln1BrIITEQSNhTrLqKsN/3a8rDB0uGMpSpBoWA8G9F
+moyf5H/hy5UWJ2c2y/hBJExQgJj2vH1AQy2cg3J56KIgO7ZVNSd2MVqJ13V1iDH
BQeSR8qJknY2hmg1lTNWkjhqGpeLF6z/7P3QeAaZmmKQf2ezAESJme4aO8NrEleG
YZMXprpaeN+fFaLDGNmC3dCAwsjOhEOqQVsNBMb1ppoM678wcdDjuDi9pVpbSE6p
FjfsUubPKjbpdd0NgsTiovO19n2RS2mdqjNsOeuW5GXwfu6SGK/ht8gT1YahYO1X
X9Rl6Dsg+rGsNkJiZqs4Wqrl3Oljum5x6/UWhgvj6aWsOrrHWWcYGpbC9UacEMki
8nJ5pOtH1TbNgu/XUYnLfZ40yHCwvExQFKX6HSA/IiAoAZ5gwayKAvGjQl13OQnC
PsxNGVHYUz9vXdO86GDHgzxyJy2Uz9t9nXKCHDNjkEwV+Nb5liZGcGEMI/N3PoGq
RKHk3Q8QaHlxEdVCufX/PFqk5lia3JFhB3D0m2K6JzJOLpwrn5jYv0xzY4Q+cX6g
ycQzjpFZrRCGbBRuzf+XoDoAcpnSJ07ovOcyZY6P0ynBVJaXMkm5nGphM24eXHUq
rpIv/vAuOjpQUlSTFjMGlj55C9tMbOLkzsuiK+PoyoRSkwZmm4e/nj52mld6ZCKK
jFUbJa99JtqgcMgZ9MyW+EyR40ohjm8i3mS9W1D+Qq1J3KxiQUgLuSVlWJVld2TL
BGO2nmHqcIiyMvE6em2LonoJJ9VR7Xiy52p7NaD+xUcj7XpmP3epDDYU3Il7m4PU
IOT0QwLIJkxfRqKM145FPuEq81VPO48kkNCxVbzTK4ZoFS8unf5OMoqA32uuNUv+
VhPGUbURiq7FqRJnyGIgP+Whj8n2gb16oOGnKqR9o3lXzxOB7I8IPm51WjqeQ96z
WIzojnl6NVOPQdBRxey/WStFX+jgo/lg5za8EfUIe++1VrLCnsNPOANxBtD8Uc49
D2P+Tzjlkp42DASIaJVI4kQg7j5I3yLSPIMGoYF3DPfU3FbeE8wUjns0O8HGxWv6
r1/73+4whg6eRHyb0r5uYyr8sAzlQGNDynRfr0lhXmofKilxTqFcpzb0M88O1RrA
LxIV7jxWqmqoFwDAf6VNerVFys8E3LtG73DFWPg/NnExfyOZOSaQsHMziuoL2uEA
6zwsqLHBWBVT5K3nURGr8fIgOrMAKnT1eVSy8huvUdos/18Xw6KNtRETzE3JG+5f
2CyUNlPp9/SKwlielxQQjL2tfS9V9O6O+k3PSdnxqTgI0OasUOFg15wRoF+Lt/c6
8UI8O0F6DQjZCjWJQftIaOQFSdp4DWlVT4a7VBqZ7Jkh5ymXGdaXccK57M6cJsjm
HOHhELKc95cCRdY95Efa0mpMqBimHrapTDMPK/gI3rKH4QLZuRo4H3DfU+sgcLt7
SkZ9WrsEFxO2PnxKf89CqbNO57OxmM/cdyEzPducUUC5iAUWPyYm0S/DdFKedqSX
fX4eLZtu6ZfJ6KPcMlapdsSV74My8FOueb1JDwZ17bEu1wXem/DbhY7Z/QVrPyJt
7TOlWq+nWFvINNEqB4pyd63A9EPmxbMgnC879tGi5oz7Dz2fMCpzfTZbSL/NVhei
TFJde+RNK6/IPze7JfvYRfNeFYobF/XBoGDiJkwbXsor2OdUx3/TMSShmnOfMWSw
X2o6Oo5qAoMEKG1BrqD4DauyahxtVE+foGDJ+bC+Hs3lVbIsd1Zr68ZMJyIAiEM3
MAWagK1yUSj2YXb045HGbbACYMLJQ1OMlSrAr/RHGPGu6SPQDg/bF0oJPhf5G7tv
PWB0IfFlHlNl2kWKUpwjEidaPB1RXOmurEYHOzVE+9DP+y7EcmiBQ/biTbB/aIYh
wPJX3P5Q69cWZiLt4hHZcAcP3KSSqmuttJYI7gdTs/5dz95fdAMb02dUSG7Rc+8S
DwRL4YWBEjr1e1h0M+71IC6hNQdp1sgpxtJRVLdf66Q1FEABVGeDJG1qfe+U5qM3
v0S1/Si8dGSEfLDm82BeNlUdV9A9XrUw8bdgBIr8xqUpnIZWN146nS9rMpNs9tYv
KLbTdu8Us8UiKD+D0+DX1pNHYcZ7q0n1JKhk0+Tf1uGf5OTfr8IzSglKJELaPqFK
1aYNqLZPolHHmBRkpN3j0uZ4VTvSmCoSNcT1LOJ51utAuJYD6V310IuzXtZXyItu
b5/GnRJKEUFj73GQSvTV2iW4hueSNL/8ybtiLhlIn9W+noK4rer5zvCaW3fkBG7a
S1tCF6dT0h98CSjb99ODcMh8pUyc1Hf4Dl+q+5EP0kSBDOKnNr7+EPy1MFNXWZLN
ggd0kBQZTgv7U7Ptrbqi054/NQl4sf1pOoY2JLooR1is7OpNxybpnfrC8dYqDnB7
6lR+Zf3z5EBOUCt9i6IonQePrhLL2+1hYKPwvGqyfagbLXgmk5ch42FLofNs4L/H
5rtsukPiH1udxboUZqfxZRp2AC6rz/X5UxLz083tX+0ob6dF9sWCIFtAZYHIq3zS
w9W2aCTjaywPXU0cVusY1Dj2hrnCE097t+6de6qjpbVwzL9H5MJCldeq3DbdZrfZ
9t7B+hFaqg3t4xTkX2fbB6rIFwkJqn1MkZJCheBZ4C0E/jRlOEyw5PKGR9tL+ZFz
zt4FB6zvrZaT2JKpDcvoq6pTejxIZHVQ5GdyDckA9ZXEwWgZsSxcxEuOffWp1GYX
VkNt2ZfoD5nWZPl+l02W+hqSvyzRIxKoguLz0cpfMk17WZ0dUBZSBcuwz7ig8dN4
uIoHJ/r/dSPU1iYdCLY1xFFuc0BEJk0p7xh33tLnhVlebKI23SMg9TLX2m4yPCMk
TyhdIL7wtBbR/uvdTBbatkQUKCvwjMPwXr+cLbMS9/S6SaOQX05h4cEXpGN/3ZTT
yzy990bkwAasOkZnwevyXAz49P51Nx25Q4kV58brFtHY3vM8319ED71ttBN0F8+Y
85LMVTVK7ObtLbBiVRcSmlhSvyAOWn72m9WoNakFvlumtZSD9ZeOhhjRj3OhngRC
MGmsw14j8M1PdGPWeBDM4z2v7zuta4kAdQRxcdKsHo4KVC+umFLo5n/K0Cia3CqH
qQl8oeRy6RK3NjHyoE6UZ1ocTM12pb4NidkPb9NXu1I1erjPTmWpnXdWKlhvL7tg
AkcrEs+tgUgwxVtTOsghQtXQM3YQoVUzBn15nEn6byLASAQnkx/NOWp/ecw8H3wz
e/2atfQikwhQKBLC9Z49UwjZtEpRuTuK5TyH7T2IEE6u13i1ZyEOD6jELXuO72P2
xzSUmkx4lOwzWHFiRUKj4DAplK+6GTqbMgLImKxKz1bGcdI4agG6NsO8xdkyTGhp
+GKg3PmFO7MPm1eKkK1HnAHpBqsmj7xfyFiXtDqDKHfRyD1qGCoK8XdCcC+mSsUi
VgIUbXjHixfIhu7xg/3I6cMFhtl/56hl37u2FOcmmMSp+SU8ZCz0YoACn2q3NMFT
8CZ2/RyHU1+8CdHY9bVczyvWU1kORAzkO2beTtTj4PBBzHOUIiDodS7GXKzTOPua
UyA0CKJNgkV2fDYggykMEHLSTH+JznFdKaWQHp0ljkXMjKsc1yL+xCqaFzYTYIc5
yOiSjD5XO/9ZPsn6YxX12Pw9W7CcRbfPUGUbB3u3XguNmyx+wyj4TETEmvBKgOaH
/ai4/qKLfZiW6EewpFdTKsH90GGXmZPZa7679J3bXHVWIRaPMH9DnDornFod1LcK
5UO6Mc4KYDYoajr3ukpzH/sQ+CKTVjApxFxxxB8TAjDGYKbP6EbEYxCFmUWkc8Xl
mU3n+1yrtffopdh9qd+0YpZIbAEVLPxwhUFT47FMi9x07RhqQmwCohg/lvSW9yuz
h7FGCnXYYh8iWZ7TdyCggyEoYswdLC4yqMAibTrHJ8aCHYuBoka5J35wGWAYQwoG
V8MsfdFe9ZLrOLdrC52RjfjVMS1m66SIyjKAXruto3LIDSX8bS0nyjbyhKmn+j0c
e7QC4LCuwT6ama49OVDD0Fq5vXQKPCSQi4wFJsm0AjLMbKeRU1SsRIQkMIPW7ebn
CmmfEDD3VjMa7f+IwRE3a2y7omXT0n4VeWrKIfhsonSfT1e003KV6vA1HthSVVnz
kpSTsNs3Qi181vwLL7kkooJSBi/DegxaXZ3QEmuMP1qQ6UGS7d64QDfWxZTrtplE
JjaQaADaoz8O1/myCauuPF2Tb3Pom8+cJTCCdQD7bsEP9S3t/QKBg/0Y+OxO4uXk
5ByzKBA1iKZQKrQE9ZltpHyC/tCu2uWM4DkrIgms0ciedJfjSd2S/zgZ5S2Kevzp
hnWanX+TmW3V3hJLR+aGs3CUgM++jXtGwfsZa47zhJSsu05aXRBq4efxy9jvXGpz
IyRWJD2x0QyQ0UZAXAfBd/Kxsus7jLQtrqmlwSGPGXe8OLsBPfO3S578JdpOjDN5
rmFozWkuS/WkmJMwadMRhVooy22xKa8wUjBx8rqNkhWuQzcX/tp4Ag7zNiV6kNwu
X0x4UkgOfp8aJ8y/LnrpbswsBvd2kzAleKL9ei0xOhO6rbgRmJHQEoxpY7PYCpSl
MPy6NbBU5iSJOrHxWbwnAY4Ii6a5dsh+3M1jkEgcGwtLDJEnpM+qPRYX5jheDb2f
YWOEDBHPX4Cvtuf3Tj9GfSoy11ufEM+YCWpkMoJXZgilZITizqxqVx5SzNPKh1NP
WFWT9xIY71F1SwRYbpK0Q2i2kY6t0xJyEzanOLdTmulqu4CKPkV9iZ+RAZg3c50o
kOr0y5ubV6tq+IUIgPfnIlZj/JmyX09VJMtcjf0ZBYAHTQPYqldxVLjqAqmn9jJE
NCjOwXaaE9W+/H+h43NGSs2Eyvn07xsPirTByHU6unoOlX/5JN9QFl12zKOpclJf
iwejO1RMthUF4reHEsEePEN1a+r/HTZkZrh+lsWE3MDc43tyFGHEmuDUHpR13TH2
MirRkiHfVZR9UIzsBRDI21lwYCybroSRRAeJzYuZErlfA7BJdM7lhsaZDcLK3P0k
TkEot7d7OS1/D2N+TIFPnQNy2rJpbNp+csPfRmkvXmoExfDNwtvhTwowH6gqNQuD
5QU/GAiRRtb4N4wLsoyEf3tw8BBNot2YFTyWXHXVxWqSrYOH2MTJu0g0vEoD4Ce0
4ghPF4xhVLegyN/4oc+tRZyZCgWk5w14qrTnissidJcDHN5l1yQtX9PazfxSTIdq
TZt6Lr9n8XmPHWkHpUM2SMAyrNqvoIvRcfkaozKcuwCaZJEexl3Fe8dANxDUpovd
VcBxlAyAlod6VrGee+bPwvF30DEQ6IQS+2KQyBd13opnB9VVnlZXd6qrlGEEJz4b
D3xvt9MQznMP4nZhAl/IS3RMHZUU/T27PUlW5GZhVg1QLVe4SgTb5Z6S6FbiXklz
10EAdk+wL4pjiNKW3dsDCUFLtc6uR6OVRtMaLMHsF0mQ7kIp9j0XCv4bzeh2DaBp
0c93cejtFZZ4g0iDVmAyqw6r0K/ROfCqcJoChOryRXU6to0RqeCPjHtXWf6cxPtc
eoOMzxIfINuWuE4/+b/F+yzrEaryjvxh1rjkYydNHDfzkBskbMv4O0g1xy4/3WZt
JB6O5prSqGdzFheDmi2ufoywxU6nc5B8M4vvs1pmZmXSLO0Fs43UcMQ9EbKJs5lq
C4mgUmjQoGeloa5ykbHLdOIgnugtbjIlvpho5xxjAsevdETE37B24rQ+jPNwizXV
vOvBSpHyhiRqOMBEp68Ot0FIT2MUZ45OhiOSWvdNIqd8kz3MiPQPlP8uRSh4hQvV
6nsgOtj/ia4g7Jkz6CMXrw2UhcDSshNP+KpkYlGYIBkObjn6dHW7lOsEEJz6VmrM
ik02E+jMiBKAcr51XIRRj34oPWed2tUuoRUBLdHBonE7wAjgjXoIAUXgdilUYNVz
/DYivFyib1UeMTwwwApUdTA+yvFHurm+RHN0BLjqesvBdIsyI1IToiMjGqnSPvdf
fLHYCGAA3fvi0Hy71otM7+T51Z+87B3q0Z1aE3T+DeZAU1/5qbhA6A/H2KcC3g+q
IL3oCEzac5SoweH8wYkYCqoo3Ocs1N/c9In4Yiu+WX59CRfbWMt1UKdKMiayqeU7
ubv18x8XDs35Hb024bHHiciHzigORh5m/T5nzyNakd+uMIqbEbnoPHBibqRSj2Wi
QaQv3sclHpL2GiA6a7fpep+ff+8h+bR89ZFPFRPtcfOBr3OD3J5O7N5meABJ/3mD
kYwVN6NPz72lQfGRrcVAHIXTIJ9Hi/C7EvPgXWfwEHha3nSrGdSJcpZ6hRxx25sC
JrbsFi8k7WzFUg7AYnDj9jvnyULezu69sgEJd2zu4MIyYHbbZQ2MvKRPhlxAX3cj
WGsF19ZCZPuro7WgiVOJkqD9701ZPN2ktRD0lyYERHTaio++Mm7SPHDtlV9Dhvrn
XH+VfKT1B6itaOkYXzPis+Hca5gXtZ6EBNmPidI1ongHOPhVS0HpRgLRS8zvTybC
TA1t50q7MrEZgz7bqM2l8gkHIub2LWwNwuwqQgpDajtPqWOstjt2/pW8C3ZV7vI+
nhMMo78p0WUnxX8ok7dPpKY/JAVMBZrwAj4NIOjiQJ1MIwvVERlTYyB+/Ztjkifc
VVC2GnB8QYWWfdMijLzFDaCfUIX/r++pKRHhL710LTrGTKLGeq/I4wc32K+SJHrg
odH20K3fiXf33ngOBAQ68rR1Zy2XBLyyGXBYjpZ9GneeZEt0ROZCZjWOAkJW2bxZ
vJlei4stdaUNLkzYP4sN52ijOaPCEO/fZmzrzv9i1MlAwc6zRbs9bslM/Bl0HSEk
lyUO0ZmudP4nS2TX6wLej/GekKXLtYmkfrpgS5krHzD/4gDfxMJ112hos2gWY8pN
04DkMoqFSUxV3gRbmOcBqIfdgDwXT5Dy7jmnmpOPB+XfRRKDPogCmRG2bek8qzAH
6XBgTM/juzwlYq7I0GobmXu3/h+yQ4T1RQZHdz+EMqQvo/OQUh+8BX6+mwl8bVX+
llWdIEcjYS/9Nb+/fmvvxH/qWLVX+fPlTyI15e07fp3mNJJLSpHmnwf04e2jNDjv
bUeu7DGIDxrF5TLriDmwUAgIDmlee4/4nxtNY6HXgSsrW4ZOw9QajjGOqWKL5vSD
0XI+/Xd0WXYAz+d68RCUJCeHo6B6evDeaFQOj5x40mZPlHBcoODObsUekdkrkgTl
aXBoe5HMS7+4EYFIQPL+oIfWqJndLwrkd4K41jvVFpJzh1BN/J7IPHBPqY3V7jQS
pHwlD4fcoT3UiAEoSuVZeN9A5nzUtwdNbL0WsRdtZKtlsGH3YNJP7jMsHMijfx++
u6ErJ8kXjz7PSKhxahIJMc9gfqxUEEvK9onLCWJ9H0MNyaag+ROzOMpbcY0gcvQG
rlOTLCyJWQArYRfSPWuf3FOKtPFbVFp3UjXFzT6R7ubAI5yhN/7ANfsGaxtXuJsL
9tgRe6l2P2K7SaPfmqoXdldGzwpUm2aFb+gdHzcZfRAUjzAvxUXuqE0h4dZn3Piu
k8JrBtmgv3UIwUd1v2BnFhZF+J7FwZBhVPnisyp/uapjX3IGyTCkF7aYxUoU9zKR
77RFUgrnnp21jp/X9/f6MF39heL89YaaRDnPQvKXFepxsdRuxNnAYeOeF70qz5aP
8TxacpV6BTRYisYkI4xtnByiDiYTgybMab9OYURXSJHp9g8fiPSoD3T6p+A9eHXW
oo7Hs7P2upRLGiWW4C/OpfUBSdnmqkNWEsgdwd90u3v/vFBDdZqJpKi8HCNNguRe
hjt3mVDEfvH70MhSMyPTuZZJzBpUjdf6bc/a+Us2dw/Rom7zMgSDUiM7Mlp+z/UK
PInfgz1mo9B1DlOkEzpbK6yBaibOXbVCuZKFoGOR5IwX3X5CK40mJFiQHYyitZh/
+K6uRB+VGmt3PmdcZFk0qgEZgz61nSEsuGLIAaVl4xhE/RIZTQmkkwdDgOss116k
hAf7A6a67MgMbNwrxUfMOJrQVQ4csnNwQw0F1annF8Nbr6FG1RJMXHH1aLg4hDYi
5eTz0gtuC1J1wsQW7dFmn1xPaJCa9Iqdpu2NAKd2MojPNZDuxrNHMJrlqNQVbdWT
OO89WxkbRtydNL8NqfVVCjozX633ZkhlCuCIF/1+jXUGB9hVaFEqXYtbEqUG3q+w
6A5aHbLmN5Xuvxv7uTxEj1CwxNOU572Iwh41yV5G5Va6TvLCPRxXqj3hyOZUwZnA
gZM3gAZ7g3j8Jr5KwEo/DqxhVLJsLa7Vjz1T7gKks2V6Ltvg8bTbTCl9bnxdmn0k
1j7GzaqSNPwXNnmKj2BfBT2+GvxKbQ01BB6I33sMJIxWBvla6V2xFDZg6b5OD9Mg
Jhb6eoeYZblGG50QVLxd+7x/m2PeFBzwfk9ThvHS9m0uF26eBvmB5Wa8zigQ1ihs
BPEokOYKbnCcXV8jrP4A0dIQHqyHNb7k4KnpO8S+snK5ZdYOMYgo6DDsnTMl19aK
9DWIg3xDzN9DUlewCYapdS6cylrMy6+GQHSwOspl3TKe41ZG4w2CYjVdpN/QJWNR
VAzy1E60ixfrkr79eIZTewR2atABvY9zHBE1KsrxuqYcEFvhNwIDhuH/CcdxOq3w
lP6ysvHvJ78AkU6z86RybEDRKSKfgnPBlDqzyDgr4+pW5cMCBlcZhAQH3R2ZQ+2D
I189ELmuXzBhE5chRsDLy0i2T/2tOTzXbJlu5i/57jVHUfHTpMvWJQFVTvUOZLpy
OgvZQJcXGi+tt3N22+uNMlIWw/AlPL3DfT2V+5mb31rN9sO3TpVsnE7Htt+Xn9/2
ihwyxaWHaw2McHCR7YL8CCtEDfraPCAQ7OcxvYDABH7aQV1vYoThxN+2kW47ruOu
T9WW5nnt/2h94TA/aRx6fsmWkJTkAwRVfyMddGh57c3N1bxM2861tmH47GFqAAca
NOzt0PUmdLD/arcasOj6YXlWicVOloS2eu4W75V14Lo0+IdzInhZ6Oy2BU7wlJ8u
7P0bdbMyH7iQLq+1GGeFbGjOddIvNDtBTGwygpDnJVNxGaDvtJf9CgeFSYOMz19W
ZthTCPju8HAHFrQVZnlbnGV9e4iSixiQqqF5j3MDKukX3XgOLns5kFtJz3j4YS1B
T83glQFHbRPges+flXcy6moN7DXgadgWpHSg5LtnZC/mM9Q2wqn9HPeFfr5zDjUJ
8Htzh+nYgCvgImw+Rv+QhFv8JErwzS7XfBs/XCuVRFZeCHeqt/nyfD/Xc8+YwmkP
q2Zz2Yn4EVINAuXX1HeiyyP3nveXfAfq8R17B5KG8aNy5mW8XOW2lytvTNqxdmF+
1p7Wkuwf6QrMt5l2+GxZlgPAyClOn3TYdl9dpXfY+Ds8qP5HO27WMyBsaDoPuDpU
ecs5g5iJcwvBAkEcmv9QHwzk76nROTt/4/PRqm7mGxTO5STFDUSg7ATt14oYgi22
JQaknTzUjKaiX6YVOf6CHRTPVt8you/o0wYgwoIprZkj81FQ/1b6nFAzlL/f1tVS
/pCVNVO/XEYgx0yQQOvM+85NNzAvTwKAgYoGvvkviEFZVle358KKzN+jOMcLbFY1
mPCw5km4dKwZ3xn2ynaM73g6vBxxduQOBeKXhy9AZwwJmaEayGbwWeSvWdGiItUf
j2MRNQMnbvXUk6OH8UTR2ntfa3PlVFzrQzoRi6eyqHJmv8mhNbJ5R0MwSMsC3TuO
JbgTLBSZsONuTxmpeZutuM+kj2oqROxWCFP2RhXGngZ4NIeMRL8djyEErYSkOpX3
EgOsMT3+MgejBI0+Tf9OeeJKr3GWcszaMO/dULT9mbSWQP31v8iBYMRYPakOF4Lt
lTB+Fp5dWZMfPo6OihdPjlhd2eNDK+GSPAWDHmbDOVqLwxB+DdD4AZUKwTvvcdaR
kUt4mENfr77SRHc/pRSbOxf1o99hcb9z55rB1YoUe4p4jJjeYw8GNmQJf6ZXdbJo
XXoo+9CFMzyVmR9D1KB3GBnOpTfxKdxIYPfYrd+td25YP8cZIBjMt9vRPjXoXoBk
ABRHz6wbMairwG44+Sj3Vk85YdsnXJHU6EEguwfSQR+iBCly0GHVSbdkMI6unSVx
o4q3lM0g/GmcMhHUvcj+F0wSrRt2QNVHaW7COdP19CRqSr+vESHTuTm3ts7aWCVp
+JuAmyBMCVMSD/M2AqwxQcOzyZ41YE/RCGkR1YiOwfwkQ0/fzOucVfjLz7E6d/4p
ARJs5snmEP3dwQKpw6e/EHmPW+HFt6+GNYqvXPDvfSQZHNJh0K3tTO0CyLIkdG3F
BPuLp2z+OtIEvjstI38r3iF0v7/jlC0I3d4pKdhMIqtmFv6rnqP5M5aq8Aba5hMH
73hV0SRtvkeC2esDQTr57q0/IfXsq2rMq2Rp8xXXIJemnWJ5e097qX7vQ0VWCaSt
wfM+v1tsR8rdsVey13Iob2xtvecFN9xZwEcZxrM4fnFYrjN6gA72sSUFCfKvhGAq
fWvWvkcPh7mV0grEEFVYNn/20DpD0Ef32rMax+0cyUD+wJmEUH3Y2etgbW0OTrGI
NljSRDfxPjgeutZAr/wuck5zw99BtY5c8bCeBaGVApmua8GxAV2ypiAPyfZZFNGt
+mgf8/2UfUdAHO43RNhauymAuzWC2QXgipBpRIOV9fmqetBp61JKM6aGkySFCIuZ
fquZIsFAZ7W3JlgmFP3n/eij78uOSnudIRI799G++j5lRkID+5c6t8x0zp/xyU5w
c/ALVWsYPIkW2mEocV1Xtw/RCMZ3gSAjHCb35IzgHJZkImaFfNa7udX85TGrJng3
KymjNdLSernuqm4cRjmrptCgaApGf57Pou61IoDuzNqYKdIx13r6bXdKQIL/v9YL
V62W4huwnq4MuF9JlxvNSMbd07sWsReMahSJZf7ZTeU3olsLG6Udtbb683F46Pcf
FRIKgrd1ca/Lg5y3vLc885BuAbk4zKf3H+SyAf8Equ/G7o0ah/ubZXEVfEr1klyn
6qQRgXwTd4+oyHf1au4dR4D79pxwgG3mqJvf2EbZrtE2SLE3miIa+NmFpruFUFkw
2rpTSMf82tInSn1VPkWzZ0jQsnpsHHYbE0xyDJLud+YZUqf9DExkuWll88a9Q+Yb
W7sv+MoTDpyQWFOOQVekvH9hAyo52lDvN5oD3IRTdnWxoHSnsXhudgJ0h1+8yYAg
gphCSOKlCyJlLWd9kgAJ4sej/DkFapX6bGHThhT2KkLuJvojIvVzIWsmR7LZ7H4O
1hnzlnxV5yb4hmLe3xJ9I/zKeZM6TQ/8HFWmPO6VHN+OEDSMxWAmQLFMJOVuAYF1
/nFIRfDCNLPQ+3xWTWjMQ1sqAzoLW/sJ4g5Eqv0PKb663S/+5pIk/u7yuiYTh0Fv
qZgeruRxNF9HQE2dWEpd8x7yB8SK/fYEhTbs8GMp7lTfctKKSPZ2fIRnsg/TqlAm
CkcIBi/edqWo/uHbH9OOrYW4uKBfAK3WloNqBahrPFoqkueSwzphpK15BSObziok
pqrXp6PwBWOjqdPSiftCjTYltb7cFFF4xg95jq0RapNwkVUrhzZPKa7T+YLy1hS6
DnY1fMvXedHCG2bP+ftI+nxsKahAGwCgru8OJN2lxohSngZurv/BNlM2sfDk9xrh
t86VFj2B3v32LiC9gSzOa2r7I6OKzfH03xm+QDEMu0t12hbeAIUKeo0iU+FOpXkc
vURtmzli6J+p3Qglk55/wHKw7v7BS5Xvr9rfYo2Sohh59+4X6vTtQ3xmmq+jiA8t
ri2wwTX8l+ifu4KAn5MBd3kS/Uri0zLUHQ3FXKgzoB/odJhFrl/xCQEzOwTTtRa5
YBApWhr4fyVPjBUpKR4YOebfN1YGOrRge8ZqY6QzsWbiShAC4xdiqjBxGNIxIqQC
EBLB+UP8WobNRAED+T0AYJBVb7tM2AmOCnKbDS9BCJnIlmgl254iUK2Awnx7KyCk
+qj7v/P3+1D260GW0VYoHWXSWkEJ3Mq01IX4fzDUMkt4LntSw9xnBrZcXRJjsM97
8KYh2EHTcD0tz94jXqcMRUo3QOg9mWwaDMXpnDmXBxaeaD1Z+S4UYCXYx32GFfGY
shlRQA2ywwcLNnFH3F4gSmLWkRe80AouL2KYK6wpv1yXJRljS311QKzRzh1NXBAE
bS6RiTWF8XC1i76xryNffyq/UyEX3qWrdHmwU1xh8n/brnVQS3igZ3LyVQ8sZhjH
j3UcgpA7NvgLOhXC7Ete5bSDPRi18jLAmlOj/FlkG8HBTSdGcMpxTFNJEs4c6J9a
9NIQtKc22jNEToHHgizVFqsOd8+HU06LZ02k4RMSuaVndXtPJ9XyCOv2EMR1P1CB
02Mydqj2FLnupRlOPTipmSLliNF3qBMOU3f7DqU80/oFOBdTmoXHiB306CES2Ef2
6Id5nEVPMX0KKCBqeqvpKJxp+zHQFYrsBnGV8RqAOMjf/ASkmxiGAWsPfMSwMIOK
+3nyAO6RkB0mq6YnjP/KI8J3Bo1D0U0P95qxZrKICNE/9ZzPk9f6wZKnRcxB1+bC
B0QSBSJZ4GMVAdxWAbLwdfJhDzld02TDLKhUu4eeLKgapFVHO8evD1QesGeiMVSM
VFnYcFFi51jzk6VA//KQRV0Ld7SN2Fh1N53DY2szhHdx5jRM0F1rs9ZTRV/7dPHY
tQm+TpEJuvycKDT3DSnweYV1eke5SeNqi4tRQC3Z4ykJfF0raud6IvvpsjGE9rTS
Dn6lAhtD0MxanVY8riKOPgaSiUNWP7hQmkjoVWP3UlAUPlMawgqoEuUX7nac1nX9
VPD8ULiApquSdTmUEcIK6BtJGAFmZS08GkL05YWpz5aqIICbIH4yBpu0VQSeERkQ
izIYjyDvDrWVKES7v09bsGGjLPyJIuhphNuewn+sfmR1bvnDEoJQzmT3HWGLK86x
LTELiFXBU3WpfsWmcIBBw+gyAWCbvCMlfR/8SeKqVu14EoHj1ycjh1GwULHRtwiD
v72JP/z5f+EBHfZ/eSFn4bRchvXy0v2w+6MfwFke0wvJ/n4y9rsQwYdH7UqGxWm4
ZPoX48M7onGt7xuIMW7eXbaSELATgfr3thNXQzAjUJuwBO0Zi4GOVkh4vF1Xm1MM
tc6+1+MNULot7SE5a0FkzaiLll05bswl/VkaYgBw0a2OLeVygqbFGNoLx67TZtDJ
v0o53EIw1MOSgvpMs+Dc6TEgCjeji0eqsHLPz5/hO1B9zXutdMqMsllYVNs8z6qm
qM8bx6NXwVcbBQMSEddWadgjgdn00L5Z1vB0MgacBlYJhfuoudj1w8rwyuDP7mz2
q4yZouAXXlxkPH6QERUO5kTaXJJxhKUi0GtQ5dN9YZlj2Le30oImbOftOx+4HuEP
2bkpnNTfKp0SnZgF9RMqmBxcOwADRcTPvwC7SnWfJJ6SVI+WYrCf7fQusixjhq/g
FbmoZkMZ3HKuOfgydPXXNkUIJ4j4Ozw5IXMdkPDb44kk8I0hujxBoXKQja5IxhNR
nkRfjm25iDdk6L4n9/SUvHnChIXoDElPd1581fQWQScn4TIEWyrEzVQnGV/DeEwS
1+CyCBjVw3VtKu7jXz64VAsNMQeJ+zpTSKkPmGtOHW5w2UsvnkkHlODJ54U8ZfRb
m6fRRmSM49f3R2Vrb7b8CGXeb7iHUj3g1JKv3Oy8r5XGyHsEVdfBr5rNXKkMPxdx
z1oHtEpfQSCHC9IRhCcXKhtqj9RrPG+i6hloMwghgOdd0xXvM1Yo/CtM47LWoq2G
CRRrAmNzQfcLcRZFrmro3IITMqDMoR90ILkZ3M12hAoneYGzH6tAkgcaERyE9pRz
kzRi4+hcKlvK4nSXNQCkf+hVJRt0j8cLw9iAI4qe9QPP/p1kVtgIxCnrjAlv1KpE
jL0uIw+tDwbOmHH+aBo+f4RVX0+IwfO+q/ab8dwUbxyJ9HIss0Aqvm7ixqGLbnWp
6wx1wYhmbAJGGiXpCcWmb5G13oQYd9AhFmXLqX00y9HDFX/QnTpzUVXct/2m6JDY
FR6I7+ytxO5e8xVrwTk4EtfT67zqRfCdXMUgIMkETMrzVSpikB8Sc9h4WCVTWt0r
VD6dSOB0nBGhy+EiiuP+M3/i0qrJLxL5L+3g1wrcldw1+EeJqkuPlbNHjTmrJSd7
r+fu8x5BIjkGA+8ig4JF5ZH+9amPkmC0ytsy4CmupbrD9qo3Tz+YC7fqGq2xohG3
M1SjTKDU7hijMK+kNCa37IcjPp8CM52LMhlYvRUe1d8E9jhqNFg66Eho6pRFZkoM
1gf0H36bzHV8VAoR+C+zTx+m/sZYsTqlwwBHkze2FMEmUknRIPCzOGqvQMOeahA+
t9YQLf99uZ99XCClLpWEk+d4C2wTgVKYomw3cSmwjrARYB5/keMn0n8l54qqMKZ9
i4OkzvDuKKpSbx/ZZa5+0y1pWHiJx22qLTqlYIxDCGnzOCc8ugZL3CLkSxfjojh/
c+Kxgch+sFc1dMLqEXzkSjYpN+6o29Pewg6+G7pUwFrk8oaL9RdReGMniREcyfYV
MGy/fU4x0vXbaWG49esvJ1a5fQ0nKZ5B+hflnOiMdsLZosTxvT7X4Okx5oFrrPbc
yXlOCLxPqL0qW+9/D2Q2+5O5eH3aurAER2xUXpf1fJYHnutJMt68onW7bH1umsRL
+cn7VJamriyNoZJs/aYkyPt9WFerPaYfRTqx3qaPWhiljegwD4/6TKtqW0+QGHNT
yMfeFceVWncjx25ZOy9rp+4hKzRQ2lSuEvSXfo2A7Wat1VcD/KlN95YVEsKj2tYs
siHIzwIggTZKeXRyk3bLZbqOnkRT0hKLWFTJaJwh838f9HUeaWEh1WqhFBtEJY+x
phIKCsMsCatNByGxeSCPKojaY3yTlX7xyVgM3Mln8bxwnfrZR4i+AIjs8YToUHQv
euB5qcagu373y6Ptg0a6li3ceq9VfT9VRslTKY0xsG05TOiSZZKQOV38UqFIY+n+
pXTs562Fy1H5+r8zBjCGJ5ey6WaMPByVnUojg71ROnZyorJN0rdmcgr/3epL/lru
oFGXzvXCzZq8qj6fPJ+/mR2veXtDAm5X+RSh6W3fylFJv7GYxy5khWji/K3fcUXP
UbQvpa1XHPWKTZktseX41j7z5b1if71moRLQuOo2o2NVW+GK2ylQ4FktXGCsIRtU
FfJ8jc9OhK6CefTkexustgevtthIryQUyQesbTKS1YR7i2uvJCDDcl/PopUEi6Jp
0/9onzYEXlcVasb7kOBTDL1a4ZXT+xFYmnj9iBPh9cPscnhlmuHFEnvZqsQIlJ3o
RuPRvcHpVa3iXXppG77/J9Id0o76f/gWuuwWjwmC4kAKzh7wx8Hm5alFtH7cO14m
CTbFKK8+3fXYpoCI/6vZS92evxV4uCyp3/cKClQJDDdb0qpX9xuMQmtSqO8+nLDX
qGOF9iqeCGxm2gvaRwMew0hvSJPYSjyEUvHAjSQlcJflVv/+pAj9RVZwddMbcaRh
QaP/VtE8B441vuG6CAQrvCRp0cEhbDSNPV6DSJ4lBtaNtgCoFOxOsiKBYTF2mmE8
FYMrNxzylJ+4XtihWeGBaZNTSIv+CN5LNzMYucXPN9fWBdJbTydkhU8EcozDGl2x
qFE+kGJozb9GyKDz9F0ZVl8T0mGr/2SUwFtTDDe2U5pmHHXMj+ptPMHSApZ3Y6Rc
K++m9wRoubWbwp8LIg22UwAO+K2YfqOXV4dHM1Q5bbnG8GdJIFom4EZ+yqTGv7/I
j5Pwp0c9jQfZ+odiZ/KIBMnfs5knnde9Cg4pXV/mX+YdqHYPYvaUY3X7/eUhxMI7
HFyefIcQS+clq3rSArl5wNlx3wiTrKvIMYilSRYnnZy/JnvTleEvC9NvNI93/wuJ
Ys3pXBjqLMAPx/mtwGPHgOdyeJp6dexjOPlxztn4Ib8BcORftVEiVzTmsgHyKhRB
HhdF9IKPKsaJ00EXa/zlPeaMS/x3bEpULStCF6VF1BYH7Wc7spwAfnvJKJJ4bLvm
b5PufplDGgiERKkBDABnsk4A/GzACMWhJ0G8CiRPzdqDJnH8iUB6e1tVsYY7KxEK
049PpgyL4kZ2vTuGv8LYHwTGWlxZKD21fyaLV2R66YRIuLVVLK4btTIVjzkTpNxV
Eg3argQetb9gggkxHyyEzbrTorEMsljVTbKDctVYP+tVnqwtEf0StEQ6KPKspnP6
8f0nuYHz1hhDUl2OBbuZXXLWFp3LhK6JpyuqXgYGvj+cw5B9B+jj24M7BWJXhjBv
axaPcbvT86VYD3v9qlhjw58HPStBbz90J1v8KYfr9ouq0KA0m76A1fGxz9aHyU47
K+mvSn3i39yRI+6kX5q3wA7AGv20AtgAVyXWuN+Zc8h6mCoqucbg2+HRl2vyN5tc
a1GBLFNLiN6JRvZX5VcoYYd2GDtmqmdRgRKnJP2pE36hYhsgVShJRO7KWWCBk2L2
+U64jSKMUj7dcfG8c0vc6Lban75YqoTx6TLC5RDq//+Hm+yRz6oFl/nilokWf0Vn
NAq3iJTo9rseN7jZ+7iUTYHjHbS8VAr3R0+8CB6MxzKdeVGx23rlGBvJzyusW+bA
a+juxdhUvDMCsYsaV6mEjsbIQfVM2I0/2aDi3UweuPhO6umpsWvr58hKKjM0M9No
+RRzdJMmyf8Oqk24esvB5P8o2jF0TyL0miRK1dBW5yiMpvCHYkGbMduKK1LukMsM
0cHpGVGwHFFYrJxLbgMjgU0yrnq9K/HY1UQdhUQMk8AQgY4+cATmaRYlFqScmsot
gyWNu8Rqc9G8yDyaL6W+EO4t0X3wybEdIB3PmmlN/J1V5SPfRFAoW0HKkRvrm3et
eKWD1VgR/IOfMQfKSr3a8Fcks0vjqTPTDBKxGXemriI71fG//el+n3jlSQLthbNM
KQXRHdlXp9JYy3lmf7siEAKWlcbo9MZh+jBTSbl3+hs+Qf1/12bEe2eCndkSop7x
Vtcb/4qg1H9ovvw5OUpFo6i+BbnsrMjt/pq6ML4B6zMa3mp4DVo/5PwM+biWKxmd
4CPXnvT1/Hfqtt4J1gBXZ+e+8KspQCEtlyhG5ELogGMg+2kr8bC2LD/nQJ/C7nZS
e1zlq5bB+ikjHwvdznpzRlPnd39lanueS5jmIsWGtrrTCA1j6JA2VbJfwvBQ3F1I
0DJ+Gvz6GY9xzOCj6/yvYz8888z8vibvuINWJFAg56+/9SZC6lsNZGRf+99az3gJ
ggtyj7OPmkfkY1tkMLP6joJxhb548Hoz8l46wJMwqlgg0Q4fayAaS4SqeJRyVZnB
nvDTO9CUEDOosRAJjQMpUoNqaJbVhIkOIZI58/JJd2PcDjVn9uBph4Dl/tg5gBJ9
gEGsc6re/+wiJ+1Z2oOPTR+ZaiMeA/UrchoBUAPhZ3Gfckfk2zRGsnL2GHfTrwls
qTqRYxjdExAFjgJcJ75Kk1TMC21MY6KtyQO9BU3kTkvjE2OQBY5W/TbZJq5sVgYF
XfPsGpxykWsvBCTWcL3eA3PDIphdpkipz45Jc7zjHtPLb4dpTuNciX/sr8ZX6Dzp
6tyeYJRHNNsJ1ApKRVO4diMt+Xee/03AWPJJEdvJtOYzzrMxLlBkyX0pYf5XvcGk
8BdNudnMqXg6871Uogslbf1GueCakvQ9BgFhNWjgelALxdcpOJy96wMzHwu92UHK
PMj/Ze4gTYjj9NRKycUxQedRuXQ6LAYSIvWhEo3I3zyZOiEzU1gZAqKIaE1eVEMb
zmNWlMjKJn/zgRZvyYIj8ag2JUnyvN+z2UObLAc/2W3dBe66WbAzBnCc3sCaez60
zM6oqFP4EA4GIOJSFHVQRPYM38mYvzrs3KBGTK3Bdq4XjS8yEh36dXBFFLz2FD/c
EkuCgRwy8dUtU4+m28+H7VJJxB9l6oyr8r1NLjXhDOedU1vYbJt6OYKaX1PGcheB
VjmXwLJtltvv6KmeOrdw3u+JFNQlj0I/rxV4qHLyncymO+TBgGXJozqFWdNt/1d4
fpFAYNlPlHJNlB878aFOkZYsHCWwbp+paEZgKhByBj+6iHI1CixRoA9svlOJSWJ+
l5fl32AF33WH88k88KjcMjkpZXWphMGgK/1ky4dd/Gv8Ll2v/SYCiTQ3wCe27dQs
aoKjby5s6CaQF/PvKBg7PmFe2RTVGTeXC/GhrSroWQo3XdKOF8mwG72ODB1qWA4i
eXjatcaufcNnwqHG/02PQf82JZR6CILWIqJsWsdNpX8s9+ExVi42xYTh50aowEmx
m5AF880mQh53KPBvB/DbISapZQicxK+Pf9PF0xdWZ0Tify1HUlgsONzXmLo1uiF+
jaSTwJPbedqo2ivCIsGX/OCq+ip2enAJvCgZylR8MCn3TzxswDd7QfZhZahmSMHM
aHmwXeD+W/ySZ50aKN5GTZJ6SkvIVGTLIitad7BfsOSB53H9+/eg+Ovv0Lv796on
39ojbefQS6+hM1fBrouZU7SxuTTz9uxRpcS+0/ybf2U7nLF8jM/LsgANjjT/0SWw
TdlFNVGnObvhVbNIi9phuUDZ+a7RFAqYzEAkOk/kPDqsY0dhXLDyLVV5oyq/ocI3
U/oIqkbOiHAJQfTrpg2Nl+IWxkeYqPFmOHr3A17vvB/FOFvCDzwAOTQH7AUmu5P/
r3Zi5LXrNa1dSzo9QdwV47qyUWEfUAO8wH624tdEsHfFNChyK8a5DSwKayMkBBSo
XgQpOq63VmsKChMt/WqxEJNmkfBiD2nkZ8QkKrVD7HqBiNy0rNx03HfttzgU8NVb
8Jhgp7TsZOW+jSo38x5DJjMaIgqA4yQZTjAySOGXB2ko9R7PEIwPV2CrKC/T/TSG
qir58C3alZ4tXG+VHPlxHP9jv7c8MiASlvWLGzSDpf88YoTXWeUDr74Z3mppkWNv
GTc+2VKR46EVzjPaNi51MhfPZxS4dv3U+ocBq9AvN5UMxSUEGgOrvCn5ipgk3gFz
Xxa3/alpB6UCySz0Zm/lF4o/SJgNBaG1AICKwzmmN4GQHbpUe+og/h9FCJKorDzP
Gic7id6+miSiKXV4sgOFcSzec8IJOaSySQIGYTDby4mOcXpTveoqb/nQtkPllDYg
ZBmAWQ1uwOXDGqwUiLROTw4ec7ziZqBYb6B2eosKi9lbBIB+7L/IqC81F9jsTlV9
hKoNG9mEVF7wJtsa5Ft5zrBG/57RLIQLxWSRjxWCizwTBFViRMvkjL9ukRHklyWI
CoUz1o/d1Gm6x1TztA/v0InKOuB6N9dlaCRuxDFpIFzrJy4IxTjqeWmAiDUWqaDw
kUSjeKA6R/2NEfC+0ZSCaq1OF51GkxBhSDl/58/H9WJnTiJ5ugcX7lehg3srXfCG
xIpK8oTsGwxEnFuwuokBMj7Q48g/XoTyY2qNh2v2WrGGBIk0ez3njEnJ0k+TFhYH
9OeURVjcJhAhkO93/52S4ga6yrKPIw+FYQdn9EIg7Y0/2oC4jeHVHNLjFaLNEp44
5tSgF9ybMCIx3znBrtbi5Qx+q4zGGzOQgprVibFtY7eJmo2aE1PyeppkaILiHSoN
kpfue3EO0Ucq9tiqFKixFBz72ZtGFbr8i1Lz7rZBVOntAuLSn5UsEaDRzhiv/cQA
SEo5lRFYfEapMeA2YbvsxASBEtZXnL7szU/R2JDmux14I9iqG7BmqUmfNjq8RkT5
ywYMbm8DUYltWeTzgpkktZiICKwHnrrQ/ehPDw1gB7HXPZoI7dYgpaAzj1wKshZe
r0mmyzSn0FIZl1CypFqob6nXIszHZulv+G+fDBt/CyT9TrLt2M5WaVU5WEIO5sfa
1nxP32uL3DNqxlFSmpKZMuwei2CaxaDcYKHLASf0PTRqCLyVREtW1tgM5nwKGG6k
qlrAaPxs0sEFdMSrHUKa9RoZLbgWo8EXJoXDefqMT2K/wTtzTsIKlXoNGWI6nhY6
29qx5ALLMxHWlHLG76+IdyGROSdxiwe8sQLEdQFTORVPnxoRY0mu4wUqmG2BhkGJ
cMw6i5aA9sXG3Fo9x0LYM7V03S3MZQTwsijdGLqKpFaexTDJS96Xlf/DDWQ/0DYE
DBHglIJKGXo3xFQ2aaeh4Q/UwdNsp/HCSms/EA8hHfUDOkXDIlxbyy58BP7FFmLz
pUyJAZn1d/dy566rv91m47/PqbRHE4KZ75ssAsaLuE9VVcs1TXeA7x/vAX/s1qsi
0O7gxWikaDgpnz2OQSnAoE7JSlgSdgEH6d9HUFb85FvNOdNGNyLjf0SAQ5gTaZ7O
aONKwTcjLLoKhXJZ87zDcsRVMSzW1D1B6Fp5fgE5bjyZavJ4ufdKwDZWIyRNFFVw
G5YxrCCeaa6VWjSIPsK7L0e1ay00cvgsqZ7HI3TFE8zM840vVAlTEOGYsO3ma8Sq
JdOxu1SyA809POxznew8ekxHrwVibx8BvcyhKDs3I8FAAr/cV7ybCbu2P+6hhbqX
trIjKwyZ5usHVycEK5o3HYE/g3s4kRWB4W3NOgDyfOPfP1MyynQs/RZMj/NmV8Mz
GNSagTpaFW8rJgxkXbv/lGFy+8wgP0XC6IP7yIXFIgJQQ924xTwqBfDxoMzXDvPn
VnhJbDBpYjOgeFzmkPUImgg2jt8Xc0xZZflrX960lBWGG1DDMUMZgP6osabwRnZC
rzT4970A+hKe4VpnQXPTel29OWygRowDXOjmBz+8SNf6JoqBjoWk4vBT/VISmRAc
PDqzK1gjKFwlXKRFlEhkbXC12Qu9OYCRNdpyGr0nPEUtqdtkd86Pa4hROSfi/iO5
dLQI7WWvBkX3C/MgH+Tfigg/Y1whAXywPKMw6oLEzORSFGmPXDXEJi0Gin7tJin1
7xZDyYL0SScf0Y6a945BBgiKD8e+p+rfXG72hEtvUa3/Fb4r5PNAOV2iIuWKPyyk
RY150bSHlydjxmy7/UUxkVUPksTo3bsQWti1A9kxj8GBavwbrrWdJUaUBWWu/0wR
mU6lGo9TSmbjN1oUoGJ+aHKARJG4HWZ06buKu+QKnrvvPpLxQx1fVffO1FUxGXCL
gvzjjpW/dX1Ci2h/RRZAMij7DyRtuPpTNeNmwT41Zmra3UId1d9a79HVfeD2m5/I
x4SF7/74CUlYFmOgioFO7bXw0qHRo5WSaycMtzBQQ1wJc9chUOgxks1ekt+mynW7
unPiMh2d0Qv++Mf+ItG03zT5rSp6Tpb7LjZpe/CehmyCPVACjiqqnaC+ztpdkO97
MG+K77PDjhzF6f7KmwEQQDJvyeny2xzcmSMsmghtRytm3gsfzWN4xjNR5doBxFkS
hIXNULmosmZk8MljPHYURQMyhOK1axd3V3GcoPU7L8qoJnTnw40SAjbk2p8vtBdP
dYJc/IAJakpnuiczW1s/O7dkPAii6zEbi+NkMRaH/W1oGSHx83xhGrs9z677Efm3
e+5DLcKbLbCf7AmUtiEJgR0QOVOj6tT3ACwoe0vaC4QSyphRc70i/vLtb3d+Udv/
bO58jAxY1PqquS5uTEJkVOjvPivNzAGaS0vJJf4vo43TVbSf+M42rHU0ZYo07z+t
2VrNAQQpGbu0eWfmXqPOuPxpYu0yzWMA8Ij9gQYk7j4LWNsEmknotZ1LgqPENBYE
VgUTvAiFbhz2Cxb/Ty/X/e7bTIHTiFnNPqr962OEYKkzDB3Zacofu1Qrv8AULYr8
nDTGu+ypCIG6p+QDz9HXXQVyGQOIfm3nFaPuPXWaVkCu/6uAHcbeCOucgDyVbFrL
jOwlUqyidxBQRCPIqbUFDJA6oXElpc44Nf+mobAUsn3Gb6JjugoTBxMZjLfnroOu
AhbLIgRWha026Nt7tmcXBKbpZcUSAisIeaLzOUMTWT+0FWJBUy0awsYUb/KRCEg8
yZt7np3FSxNs/74WmIRm1XPHJxJLkhFovApTBJ9HbJAYfPRSO6khGKk+pkllQdYB
osbLJFkqTAfHVhB4TVWr1CLYixq7t+MmAbv6v4CBawp2AnqjUMM2Sluhj5tu7YKY
2/sTC90/fMkoLSOTfTxd8qs6jc6b21AE9iCPqJZvM/h4VRiAfR4w1WfnXjVwCIro
jvE2kXZQat00F8LaJOCROJ5isB5lbBejedQ7pAUOmxb++eP74W5Bo5wJ74JQF7Mu
96/LTJzSkrVOAyjqDf49ciOEdTXYTMpWGS+n1XZQZI3DTS7LZN2CEWrjwjPyuS5p
kaWsPIgffeziIkRkJ13g4ATDtfl8c/1+GbKsVTBVEotu7P+Se9NQ8GoZKld/zCa0
aIS+G2kBs0+wTdPydtO82kmyr10H8g5DFciPuJEKMSCej3D/e43Q0HgZ4OBzv4xv
uBa438yeMBgstniAqROv7A+79MvRspitNgPqwgnlAPN3gPf0FtWYhoQ92mDvBKIU
hG2NBOCqSVXMSuUyXacXZNTxG/6E5kHoglkShZ8YjWZ5JVQLhKBkBUIEuODplYOc
drORwGX5Gaido6cK9s4Up24NC9Y/2BAXPiadx1iPoGr0bi5HqxZEcBGI7XqN794G
jxSVQrbBvo8C+LRjFq20srLdemByArU9p2AqscEj7hR28ce6KxJ8cW/0SgqG7m5F
juXulFerwsbFfe+d017GIOMG0Kq9q8oXs2otZeq5XLsMCkF1R0R9KefJ5fcXuWcn
d8EysOraMv49HejGXH2SPtXJRaiIrh1IiNTwr2ha2jo9CORaU3AxLmmKJlEp1YJF
LlgcBLEvVXdYzUX0XrQuO/Bt3no5BxCBUFTHm4ZJVyMFqc2R/LZqgA98BSlEUyAK
HBiJi1e3QTJOby6Iiu22xskhyxRBoPnUZodqUThisHc6LGJNIzkrHnxVISUWUDZs
P+JUBjFUvjL9qGWp6UTeicbUaijKH7XKGWLzk2O9kjaka28M28xAIOM3bpKXI3fm
C1YJbf7ek0dyVDxGbZvLG4gB7Yi6phkNpzzrG7BOEZoCC/yFIWNI5306KW2G1KB7
xvn9iGriRt9+Xt1JSUMQQjdm1YZ57dcf7rdamabkB0Au+bYswBU5QGrh/+LSFG+v
/8JyPkj1OLqcLHoSs6Xti8XQQYoolI6WFnxybOk1oWDJRz9tG335s/Pqj+7r+f9t
B1FxDlVxLDQKW37lLztXvRCpk7hCDiAnAPTJyfZUSQCY9E96SGOF6n9Bb+IIwvmL
Lzfbdq4qMzbAwRIkNOjsCvutftnW3LnyEOrPgDcW3/E7H4urcLR4EEgIl66LpFTk
nzbMexwACjQo8LqpcV2CSYecKioP0uHqxSwSmS6KDyOlN8v3QRAJpI4Hp0WL3lzh
BgZMWofP1Vgqe/18nUa5DS7qu0laJzMpNW47AHg7E2aqheySfRDHa8IrrOAD7grN
NeBL4Mb84tB/zmTqcgQRvALQUkcA/d8ZHL805Se5LaB2us8MFUypMlv9amLhorY+
GFAvYi94qqR0VILdycYuzJZyxMJtNhWM4vLDpH/m8eaH+97X7RtTAe6494Ob4CzT
2UYkMzV24Golo8U31NkgGqTfvjUbpQ7sz76zl1Qfkg01i1ZGJq8F+YbO3pdH9kI3
A79K2c5rCqpYtluqhJxUrhh9wBp6tL2WNdfZ12ZVyiVNYXQtk5EIli4+xy/C9vpq
2JWDUjhwFHn88bAfWieLc91bn4YkWXOkZaaa5p3f/j5L2zXgk4vUOx3HrKxwiy9k
bdK9WYr38aTvy4DheYOy+AzRMWVHByH3QTyJobBQgBdJqB6t1y9W3mubDFdDUa2m
sB0nLyZPX35/qccUX62nAcgQjTTQ3ERbNQEdhzBvTh1+uOy4jT0spPMh6c3yxmzA
UwwPwtwBaIcnlBqSkxlLyjMlTcMHX6GsTCjdIDPrmiB8ctj/fNRmjjcMtxFz1Uux
TjuR7/fH+dhyxo7J5tjdTmMAIAAsHbFY8PkxKL/+hTiFdlzE2FvCPN3W7Pgowedu
8xRBDHljyBubrqK3ttB9AzX5GItfcpFfO6oq5KJm33jWzz4i1KWSk9bMSihA9Gx4
YbJo9eJyFJL+eLo56IwdJ+Ibc1a6uPtBsu0QGYOTj4D2+Thv6ZUzCi/G4EvTKKtH
V66j7Jz6lNJgkID350QyvaO7aR+Bf3Tg2QY8TPhrrPebVeREHqTV4YBabdGq0DMB
a+bmglMBK7j2agK7G1I41JbrA0vZM6p7alRzakh5lK0eijOVEndd6OzGjIO2/tnb
DVWVzT5osY3lYz0QMSvrkmVFUIWv2U6N3GIlgJM34PddU0sVihWs47sFG/LsiW6L
MT4DqZzEo9hMXjTCMM0Qu0HQVsUQYYjhv/58SPfJ3wnBm2AT0M+QO02zGq6A2w1i
5zOxuMs2zyYJN4GBUX6suerQVOg7jM53o3nlQJ6I9pZMHY/5uJsGEFWpOUpU/ErV
bPKasdrmVxfnv7rmjGkEEGokrqP11BeiitP8zGNubZz+p2AFH07z5ESiGwIFj3Cd
e/FKCnHZP+0+9UXD+92uoBOvUZrIQquHUIISIxflmJ3K5iS4Z2SftguZO6KxbCns
ZN14fjf3y0sq51EmEO4CZgMFtBF6fUili+U9IZwsgHuQzhNNUOD0eaU/vxUXIIMC
Q73f8/mGwXmjnfQ0TYh6yT9hmSxBPzcn+ughtAxaZiDsTeqK0u6vu5GfoorCaPxt
xJNA+zimnw2OE3k/Poaxtep6i/jOIszTjdcsVWKKyaJqzdSU4lW2szNQp1FaNyZe
qbC3TPXLX2d0m0Hl49NxSC2zZtmGWACj4RWLhqQ+J/wwwmYwCAUfATMfurId+XSE
UG6BkyZ6QJwKCqLzZNxgLSdJ4VX58JEhiA3ncfzz0pAt/COM2ojJl0nB5wXE6M5R
1FTun0PqsooPM/n5O+jupU6p+YM48fB/1rlzjmHw2pAdtlURDbCcARkeSDzKz3AS
IWdc6bRndnVbR5CPRpm9C5W4I5LzGzpIZZhh2YVxmyVIDXjMfl9qKzm8iAbpU/gD
Vyh8UnCVS6KEJScW1bfJCZ7ToYDD1SyvOnxyxq0Vbnm3eCGsSvczevCL4iXBYYS4
DZY5IXmWKpRKjGDcFKAQyvhB3GVQ9q7wLIZPK/EoiSf1P2nYne9JBvmF8RLkqQZ/
+XKnhoJsLU6r1M2CbixyLrG0srEPV2wHlMuxyEQ3ie/271ffGUSjTO4HrkGuufco
O7iIKcq1RrEXAyiYyMZTfatuqAn4KkLrioBvFUE/Jac511Z5WHSdy45INlD/GF0o
Q9V8/ffazrlfMaHGhxuOf7tmaXQmJbOGVlgMWF340k8MHFeaqEAH7Fz0HqEkpffC
1TPVYQkqCAz5+SG7xt858O4X514Z5vWnq3rYcbG8+7RAVigctmwZ32D+P7k4ko6e
7XOvZvuJnEse6JX9UbDbaLCqgh0oqbuZj+GZAZ2pkzSrnyxoTqAsgbLvPP5WUMrC
XzijWRBZxNYk1iCKmLRI0GihsrL2sTlbpgVixAjbbK3Oq3q73r23NZD+Uca58noV
2mxVn2NbDMY5QWhSVl5M77eG/pPQTVUj07lF3KW9i5pvEdN5D+FUOTDJ5KMHLcfO
xCoK2FAYTXT6apHoQONmuVYF6ayKhjnOMr9673W9+SOg/Oxv1114jKGKmze5TJQ4
VK2QCQMSbRdjdhjMxijBJhCBn31xZc8R8t0UlBNlgGfb2/Z/gtLauDg3hXwPSypk
2goZdsubyCtaA+N/IyF9/psUGTWtKt5Z1bmN7AxTthoVv1dd6siCWW/oXhouSYBL
waKSn5u+aVBfcLmTeC1sudVmtXrtA6RVBfgpkwDoOsmpo+OxhWhAT2QpTsfMhXGT
zoxYxMmRraB6QNlFgOy4mIKKQjRfI1KxMWqto4zNBMO3ji2QPqG/Ypk+yYqQLOpP
oCuTALIjgBGFoRoND8NGl+9re5upBYkU7Jc8JJPga3e+fY0B3q+vlNxghr6dBIj8
67hFQMhnDSJrKi0RWcatuLHrN2Vs0fKlqdbfEnVw56wd7cOYIKPjKZOWCVSIFDy/
e9EDsVH3eXSazIqnDm1SOyRHm2hc5YPFCHuZfGErFn1PR1NcTJW76sk2NYKYM98J
nACgYvceNIn0awU7XAj4DGm787NkiIoc3EjFMslr//Kf8bR3moR1Y4K2daF3BZ1o
R+81dDE2Um6NYPzpFz6gXXQFvBoJFLcmZGV7gmqphs24ofkaxAZXIFF5qxMExKTo
wOjk0ZDaHFAM1LK1sIdVb+spj4S6J81j+ujSEvszG3CfdUjFakj7FjoA87PHxa+G
Q+YsBEoEY2pAwhaTE14/kHsHt6j15OaqmmBqNjTj+l0VNq1x3m4zDbxL+3B7jrK0
Ub3J+hF0nNMDBKvBhuzUVAydbsxi034HJLUeMV1XRuznzVcfXsotOxYWMbrnhlgb
ZCBk6mLsaL07H5EReBzbo76KO3df2UxbxZW1YKWEbs4ZFTkAFhUEyC7pda3Pl8hv
L7gksgXdLPJSaDXjdw/7+7ehN+ku7riAUxMZixG12WKRgpCpPb3HnEXK6opMG5H2
gCX1RYAtwJrynEDmEJOtdjjLzZKiE3qHupT14WcZS9vf9Z6BCG3rUaiGQCXGiQ+9
GTXop858HYMsvMJ+zQl0J01lECEG+WhdmIV4CE2HkB0VA4BfvPQE7lc5hJW2SC+g
p19UQdw4MKyEvR/rYkCxAlGxeuXsgJz5tjH2AN2TVOFTgj5E3/0RXhsbUQf6rYRR
ggL8GerDUmbqQ74NzzXwf1O2B+1EVIohEgMa/eg5n2/gkKVe0jP5D0bNfDd/lcP8
ZNlla+9i2wICluKynlQAT/4GWVNx8bjX5ldMJjq6nI1kYiUroiniWNl/0gEb8LOK
I8oCZsQ6rQJqcJxI4RlecrW1zzX+hKcrefcy2IRUxFiuRbbnUQc3sp/x6nfJpE8X
BuNoKtKSR6z1kZIJAjwnnV/8j418Xx75Zk5Mnxe1VPvgG1x6epu7ynjXlyX1EBco
w/MYwGq0R6OJYxVeDpCRTyWUvES95K4DUqJ6Q8Xq4lzrJ4XTB9VjH9r4kLZv8an/
fr8/6yCsX73GI/2a+lBAhAPMnQSCT31Q2RWM4qnzT2MVl1qYd1PuKORzFALLp5cN
cQjecVnpRmv6witU7forfpET6mPfRCo7Hl1hDVeeI7c5pxqgxcZ6D7ZmiJVfDcan
oEHdSCEevNJs/Ch3fEeOcBPXuUchYys/THvN0bNfj6Q/pNqTiWvB1eCkUMthiJqp
dZ4UTwOlKfnKCm33puCCKN0KmnKIJsKUVDQkKiK5HHd/lJse41GHrOhbfdu1mXKq
EzJ//2y8pjO03gu8rY9Y7SFoNALTo1BhfkLk9VyqdpBiKRPlg5++pJjZtBV4qq5S
kMON2nqoLHaWORwOU8f9A8bagScaXbIzPRhUkJokZtnycqbe1LgmgawuAQQmcvwx
6MorZwFI8bsqzN3MZEfty+ZT1Ik8ZkYJMB70BxcodFSXIuQsFKLP0ciIA0PE2qfY
MT7cZ0TQnOTppxOGcc1h+MA2kn2FHDz3cdOg1S2FecFUZmuQL/Kp/cA/9haCifu/
wqMJACrd+Fcu7JAcq49FjarHtLcy/JLEdAjP6IG5CDdZuE09BTlFKhPFXIAnspLv
11/9X7FLKTzLTzDkJT7Ka11CliiOGxXkufc6Ics28vmObY+GEc6TqPWZBZrvhwUX
Odwsd8alDdSFLs7/iuO/wb70ME5pJuqeN/1ZCYr9AWqZrE4Lu61SeM01a94Ol7nv
9CEg59I6cRvGyPQAVBLx5nTlPb+jJYayuDx5iM1sjbEUOeqBwnbrNBUgB6cQg86G
X6QNzDpONcz/iV54gzeL/BP0oSom4RG7bpM/nHAijU0Aaga2Yjfry/T+L6r0npvx
azHdscln9DbJ3fKvHHcEl/TB1QXOFcXlOJHyh5c1D6vDwCuDZ7x/qQ23qlcn2iF8
kXQQ7OTxm0ZDmjRDLsrIYxpybjdoeLnMUicczP226ToKK/gyRzB8E7p1M4T95rSL
89znjgfmjIlwTh+Jz7m/dvWGxfwI1B4tppdHO+g3zJyzK4uVPahJ1drE1Klt8OqE
OXNLutp9oopxwS03Lx++5Zkacz1HmnmEiVCwnBxBtcirap4mN/EpQxTTaHBFPhhS
ZX4j9Zsox4d2InX0iDJPraI0U3sqn45iRr2WuRklIf+v6huyPlfK/1zi7IXTa2jG
pMvIRG3wiaiFRNqpJvbF5CCmr6vJ3Vvz3m9WMMySqZ6/4cG0CUkd+V0PTuaGB/p6
ZJroreMLhBvMySNunJ/sS1Fll2+my0y7J2qTW/x+kpV24JTB/2VY0eKHuMNK/j+A
7s55ko1YBPhvuhNm5ClZHcRmGD9nM1S0rnc2Nbs2LKh44e3ym2X8vR1eugJkod5K
yHTBpxVDykK3+pd+6uS8RI8CXbDAC1SQJ1FPHVTRHWqmWJopwMN78mqwylR5JUza
ctAic4+6Qz/TojYmQFAhq6eUAu0OGZPq5sbkTJQlahRKuWTuhMEF12vBn1r6snFS
0OYCVFtkHqIZ6Mck3UaOhC6N6zUq8mklmRmszttsuTXw/mWyKxsHzkIQ54lN2r4D
aVVBxrQwHKo3OiihCULgud6ZsQoQcN88T3G794kgu+snfI9MS2PJNGE9uDb327x7
qojYEAUn/yo/t3SviuvZOjLPmvHgSZWcdMikGYJEEXioudJPAV3IUzqySi02EW7l
gkQ50VO25eK2mFbqlNTwJNX3gpxopuMzUN12ruIHeUFDDDlfJyuyrWLciwAqBGuJ
5nZeKC4IswAoAxef4oDa+z9WmJ0BijJtpjK29SyDWhq7lhdKtcRmu6yRagdk2s3F
cQyin9DtOhMo/d6L8Tdram1jGclow7bnTynu7Q+h9Hv3UX07F1KiLTK2gb7OiC/9
AxeeJ9/47WjvAXwUalFkBWNmXpQyE6QNsFHhq/L8tkl45AR8gPM9/TCYfbh2ZBmC
5l3mQOulI3HEnoovCLacAHWReBQZ/pWfDUxDuDlSbtNgo2kqR3+9lNjNBytOHjnN
JEPqJvkZIS+d+fFZhTXef3d3O1wIviEJJG4ctWB3GQv2NQ6zrX30Ra07Xrizkkpy
fIy8CPG9WVLf//SxG99wpuIPVBpnvqseTlE8uR1l9er2xjgV77UCWD8Mc8/o5+0S
sJdsm3UGEb36rqpxEuXdEznZD2mt76rx+fJnDj6sMM8xLwjPx722Tu3WF93skOBe
9fGrMCUhmP/uFpak8z6XsXADwm5Oka3gUutkdIgbrWqAtEBAdkUlgGu8IogDgh9m
mKEKLw+uAZw/aQyDW5eS+mac3KjZ0Ne1qlVrFp2dL0nYq9rAUVAc6QJuqKb4ei0z
Xp2GBmCEr38djG+BLu17mYCG5qFJYkCTiJgCkaoRD3zkuuio2zN+4srUTl6SGXR9
673AMJFnqn78Iues9ugRJukEdRDpW9wUDNZi57VCatu8wrYV4KXAESmLAP0ZyXgM
yTf1X4EeYVrWsrsO85qZIr1+0EgM4xO+n2rGTrX48zZ1rI6z1c/m3hWjw/ktd6Lm
SCVhWO4ESd/3AWciLRtIiTnpONyaqF/OjkaB5G8PchZQz7G+73km20Zy59f4yO1a
ajPy/Wm2eqV80h8Zi8wVy9Dq3lu6EMOqIzTu746UIzG33ssLrCBnmQd0bUnmb+rj
OCM73Ol3kwZhuvNOi82ERENq+x9N0Gyn8skWJ6cMMQv5yhc5jdPCxbxt9sw58pA1
YTuF2gmMgiWIKWUg9RKfE19QitBsh5JBksmHySFVMLvMQZQwRTNbA3QIMEzxQn/V
BCWJDIjDkhNHQjVRp5oBSHr1qbtP8c7raHH3BNOL84zll6IaxvAUJlpvxugDmW8r
CjBLSMz9RpBKHcCUnF+vHjJfiFXqvc/Ttw4TdPeXVI+SmZWCVTXRlxgyL8QrIW9h
jILWEexl5+QM9f1bcaC8kGH+ZM0v4L5sOB5qGHRAPLa8OcO61KnNqhkbPD+AZ9Au
FXZZeR831O91WC+47JT2PFt/ZX7pSAv4Z2j7En5gI8sncSWixYAH0ubpnD563OAL
pmVufnqZAZZE0K3TvLNz91RKSA1alImhDfL106BVXzDit/SZBBYe2prdkcgsx/yp
BcolOfUuc0UhQ9nI6G97yWDri+6aiA3+QMb/WjQNpLXSKcjZb02Q25hXW5qK0E7D
M5BDlYXpkc7jkZtNulGEykyVlJy6TRGtGYvCLN6oBg9a209HlQUSSqz0HEtJFYvE
jhyNqgPhotXQBYh+kU5TwhQNq7+6NybBJangsS3GphOf++GeMNwFCB8xCYH5FSy1
BVl5zVZr12ugI7mvENSPjIkk1cVgIwHmwONwBXrNMVKD8IqwwWVeDCJ0NrcFnZRs
Iys3TZ/P08rvVn6VGceFV20KNeFTzBFVCFfO/7kNB1pUoVTQgdaA1aPr5oiIizEh
19et/0v7Z2pgyjg6hNlHroHBWpEJoeTApC113QXbt7OK/yeDVgE9XoI58Vi6hpAE
qn/o8HbrAmyJDErq9BChRJNuDKYMxeBUlNcRDPLCorNpj0xgYF8/F/NGxdtBcDmv
LKUjHFPZA1+6Nlo9TeVLPSF5OytHhZNRG1TKrXuWUwEryg8dDbSF/ylclUWs37DS
apT4Mwffw9VW4UaeH+9XxMtfRkIfk9S6MW1abZoYpB2O1wZM/vahMunU7abOSnCK
KaOZ4+J9raNtBaD9SqHzqwIxwjVMXi18Apr5uDBLLxkCuZZtYKAhvjG3Usp45sbC
M1EmeAzhVYkLv4izLQ73vOzLicr2c/TvdyeFq6etJCYZ62F15vf7iwBLFcBM9Sur
omokH60yELoKXL2wkgerdLnpo4EQOgms3QOgJdf1StdXuZ+ISnIJwiz7t8wK4LWA
FpqkGlbku2KJ3jarK4Cyv+4q1ltbSGGbgNS6lMmLKF3NJUO5ctyF7DhbmJ5b7F7d
fOeYW0TyOJpiYw1HeigNBgayhkVJahuSCZk2dU54Uk3GkXFxYmLSKlqAfXKBVTYB
SfhLlsFvTk5K0O7qXeWlguOglOrHAZ9DnwalK76cO63Io5ILda+SEoJdar295040
q3YrAf5qC/DKf1jRMviJWyzesHnWWyOT+1u/GKbL6ucnF2O4kYvE9uQ9SSLh7aDD
vuUIu7epIQ41vFuI5hqdIPcF+7wKji74ESdcN7Ou4TBKcdXx32cRszdfr9MuuwVs
nbXH6YH6ceiNzwFIr8zHabGkWdNVi/USQVZ9kL6hF1veK3J+Wj4SqCzJmLMWRd5t
gtcgbpZVOjzW7tM96AYJDBTCHFyzyHPAKodDkZF2gB3PVPu6f4dwsphCq7yl3FWs
BgAFqOiDSSfOCFaJKNIo0Gcw/1dEyWAirWqGs9VN6hONmhT1d7D2dr24F6zazML3
bryM6QnBDt2NmRvk6MGkEh3FcPTcjPJFKXk9f9ld1qFYR+m1Ed09k4w54bChhNhj
fJwP2i0x727rGUTSmFR79f4enZNZJi1Tbhx4chB8w6WOfQfNEpluIIWoHaENaDiv
uMA5kPyMf1j3/sUyio6SAUCSHZ3OxnDhEUNTgz0IIcFDwLb6PALf8a6EycMS2bko
NP9g7NqX7AtpDfUaL8FVIuCuoSGDuFXgIYfxWZlQkRLFVx7GgfahGDpCRhq1r55f
YKxmAIf9EL7cwA8frK7XgMiteKU7pMkdyEsZixu3JIfhLUvaATvdufQ+oH/cWxQm
VPwvMP765NCfuxPOZGFYkcXmbwF9E6AXcEml6MGQVQ+5K7yPm4+7+KhQWNyd5569
dbzLH5kNQRRgT1v1xCf3VtUS0g5mpqJclWu75mWkUTi2zjD419nLybVeQaaM5sNn
q2e386SV4eCD3N61LijG4Z5azxk6yas7Vz+mhHAOibLtfsVFd9HFZarH/q5p7BFA
9cp4BBdgb8TedOEB45PJEIm2mWPkfTAJBXJ+CqYKUGbPmD9Ix2kqv1Z1Q/xsuxeI
T+CWveo82hLHxtJlfuaG1HnWIUNCdLwK6SKUP3vhnRZLrfBOsKFoKkMTqgCqJyvG
htIY/jC3sxOdZo9zXeBCv/+JzqpDxIh9fQU1RBKd2n02s/a0JkxivZxsu8JEjXFv
nLkwJLd3HgfnpMvhPxlHrY7odsAVZkxflAftMw2DzGa+64qaFX9oDqPM32Da121l
b5OI4+ikMSJn1Gmxv2WCZntw64qNWEdga/4MieE8Fb523Mgc4R9mU+duYPGZ59iX
gB4Bbp11c8J13ch6/l8yCEBSCWytaapNZ/X+hAhygtYajkMqRhnnZvKK2zOkxobE
xayUWMrIE885b1JPJsdZMxTdEtPkQzlEjgW4K7FZ79wmAE9OgQNRpA4n7iCws6/j
vrfsR0Pp+3R61XBjOoILGz7vPmRVnChI0j7SZqNVR9Th6Y86aaP5QAblB1ZY/mrW
WDRUFjgsPkkphqo8n9uAfIRiB6kZCDcUBLqZTlPc4Pjl+saaKKS8eEZMlIk/ysu6
vGHpU1VWfMjxdhYyUy0jKIu50kp5maCjrS3C63jONHhlGj8cnScBnrTrDp2Khf3S
gvnzBTruxjvQn6jJQ3oC1ERbIAlvjfv+j6ponv0AZNCV3FOFsF9vmSoDVgOmSIN2
X8M5Xatv2RKQRQ34zlhyb9Aiq68lmQnlU7i3fhrThCtxuOQApNxo5H40/nQPRicB
+fgrJARE8nWhz3UrB9rwxQL2jv5KR9VNpMKoBdb5GqywOUYX8Lahiwn4MXrDqQHn
L/+5i5Z0XQrFsY8BaMAQpvBvxYNj7buEwWwErbrme3J1qxqfHqccSswwGhwG1XtW
NN6qiwvfNRuf88ud8Qo4aYSKnKP7mhDzRB4AFqj9lgec8gG/mi189OfZSrkc1Lgs
Lt8DDMrErRRKQkWCHqrXHMP3FP6C+cDn16jkM/y2Fe0UppTttqTiUJTPaxkEnisl
M8Eh8lCB/aJto13stFpmbUG/CY9mtKIMLqNjAppep5QLCPKB1tdiycShqcu79Fhf
aPiZcRu+/LIiycA5chdM/An9FM/oKfr/7Aw4508ThclWK5p688wZx/gkrKy0191z
LRzLdQXr1Um2VIBSjU3bydrSgNL0nq79LWiWPEzGtQqOIKGNATJ9A/kBx7aEgAO8
duS6F137iChfGeXRSyn7/6/CdW7zpKRf10qXLEcbHbjwRgSTLAUWE7NTRQKGdrdi
m+s9be00u3WVfZn4lDcT9bRXeF9gSQn/wyoD2S48nfQiSsuydKVvdX6aQuNuYMVZ
LVJjYFIv7SuBVdZEF0wxjqCcFsF/jCO7n0CXSScloizpOw6w0M3wI+rGMXg9XYkI
gDSnZt+turfKx2HD+moWLoTeC6SZcHiU8uSbQuxKn9Ur8cFzTkvg4ejsDgN7Jlgo
NtM5i0t6Xy4Q0ahfbAiUS9YxGszdKGh5CNWEGlIoqEe19HIGwXVqdpQa95tvbwQh
VYnuU22Mhh1VVPWnwFHnRXwxY8ScNNv+sSA1mpIWOpn6kyVKoM5JBm/6mi6+BDEx
Rir4oItmr89Unc5sYB9L3ZYmdgRBYf/krI36J2Sp6oY/jzQFlXc0KlTZPtAEqqI/
OEGHDYneFB2X/Svkqt3w9bn6mLJRbSsGPTb2nD26j2AX96NZkyU/bxm40AG+FYOk
3URevEshyUExa9kdb0ZqoezIevOJP/ArmIK47GQ2vKQpduBk6IFT0tdfzT/I3Eed
qg1UAZVFLOkDhXvArCmuLvcurdOhPNCP3KddvqTvsPHYLZpbj00Ljkm2uy4l91yb
8KIg7p/pPn4CDjNXCkMp4c9/LHVBXAHM4TvaIoEj0PLPd19qSc0oDPpVV93TS+PX
JRXHkCseRApprPBVMmtvvSXPN9eAIsDxVlgzk8NfjiVox9N/uMsZoCbEHTQkY9Ht
1gThEjNazHb44WuxKzuamTT2KUFH+gvRu1c231GMbUXl9R7O2fhSCv/TFYnb8v4E
6shp9NVzmoRPHMP1mEbT9b5yS1Ub2pS6uM+sw4RUMOAVqmhvCUqwFJ5jlHGOhiHG
gfO67LmWIfOCccqfr4HvCHjubiJ6C9l5EdAlAIBTDGjEitNPvrD2k3bQY4yF//Sm
RwFAMXYfKV1kG5B/wSlO7a5i52hoC1f3mUraHodvQ1OrACvA561UnDrcc7Fl7Ngs
Vw28JCmqcHRnAKDHyEn8vFQ6SywBP3dgjSq5SBBaPgoSpYaAlc6ODzR2nvInpC9l
qdS0BAEcO/csJfzDsGlR8DWyOb/L7hzaYDuC8Q39rdKkWx55OFWJqMjJNttyHFjH
DMvLCh0B6s2paq2O9MJqDJltH+9+jkV3tgu785J/WeoY9QZZOF345R2GGLNma8RM
TBKcekK7WidSaeaba6e/bNVxWpUloZSYHYeLPDPlyaKzD7RfqA7db83IVqihM8t0
0w8nPGQnLxcZWDW8BXQEa8FkVlIm5xAsOvW+RmkjMYQ5V19BrWU03aE2CCiM0DZS
kSehx9LVz1R6PTiSKaLPdeRtTSf9zPw3PbJGSUyQ/IOEGd7Yp+7hIidlvrUaAQ8O
BSOGWAK4YqD1VgbltW5B5dj+CsZ2DI7Ti6jVH3TaV/RXRpmaKluprPhbTptCd1K8
vH6oxOolJg6da2dd8WcTChgN/zeD5sigDxhvd2KJ8TJu4XFqiGMcIlR6Ozo2oRWi
dUOcI0uxzyXAt6njCIEfktgZHi0r/YNhaVysx0mK3RZQi9kDL4JyODjHQhXe33lU
zUsjI4+tQgsc3qM997W2O9qARwCnxY+rL9qXEKxb7C7PLIWViaqCuNB2VbaY6StL
q3ben78mGXRCXzVKB47V3J3CI+QL27zLWumMjl+jKYY5O9tQsztShAgD8L7LZavw
BUtyG2E9qarKTbclfKbFsjYHwebRjWivOBKO7qRbNJ0poJPOZSjST5MFYprURaqB
c7srSIkBtQj1i71j6hC/GSI7cjE3tdxzYv9lLuF0Hxsjn5dlGnFiLVNnu2uyUmIz
c2zMVs3GXUW90ObNw1jVOWcOJXN7NH379KBCRpAtHNp1AE1jJ4Ea53tyO3x8F/NF
3618TI5eVt+VoDmAs4JEjzbT890OAtgCMfOZEB/uYMTJdxf/a17NQQ2nr4afgDji
5qfilejGpk+WpNO5DaGEcJYD++LpZrjI+dvte0edr5tYPfjiJrbiVE61VMuojQyD
KZkiXAEZ1YDuldOm04aiwXkFiJoRe0W7m9yC5o5GNwsPJqwsBLOWchnKz27btYWF
PCny3Pd6sDbzaXeqT4lOwfbVbXkobdZ0DAaIrTJCZuokCqf2WVsiZdN67o7U/3d5
RlemenMsaN5jzI3TpS3ahBfp9L6Xwq5UpiHmCtXXgFWNmUl3TZzpPDZoa6f9x+1Q
5DDFRcNv9glm+eMeTO3TLTdZxENjlZk4F86J3DVDUvwhjVzljPI0iPUeQxA/2jI1
CBftw735GIx+ztoVu/UBT7ocUh/YJIPncOZlB/KX89ax793Jyt0yOWIVywOcc8QF
MgKG9O12KvuJcFyCRIJUTfYVZekGdZST+Fedt/TAkCF9/4bfkXBJL/UeZyfX3Wo7
jUqGLj6joFNoXOx2KhnQKv7/4U5nxmSAy6AgJ84bTJAgkEVbJ1LvSToUc3Rli+5x
rjn68R0xziRoQ/j0v2UxeP8Nyy2L2O8Y5i7YVEYJcUkoDI0D+kWnwGtsf+g2qgub
Ls0cfKBR0goF1MTwvBYTKaDvlz7C2DMXQht8xXRiHExunYYieHIj5/AfzUEf7kWG
EO++nww0H/GFUZMYQEYnpZtlRD274G0nqB/a3/ZD401RI3xDh6EBXolzjsDbqfjA
ZRxPASRLcnzGypkWc3+W75Q6p9nTnXrfVSR02TENuC/iL8DqKVWfdGm47SFiqehX
im5MF//L0o1nORggBfDzuZLB9lns/K2aASSpEGBama2FPNCE4MFv1HUGZdsabAKJ
TE1A0gjGepBzvvEqqPIYAd5oquNTbAg+0WEGxsRBTpnQUIlgkyZdC3PSY1vWQshw
lSnUHu8Yie1z60mcfBNb+Gga+IbpVau00j4qryjibv4IoeGgzJsnZ2GSe36N0ODp
41O5TA76QxMtLRdkS3kCgozuWMcIkNfnR7MbMWL+JtftIB4MobYC7e2C7w/bKJQT
TXolcxiwlBUi3l5CoXvtbojocniRNzT0QmAYk99eO2F5Se8IuXSmoI7lsgiqfeJA
wTcd0Dpt0AXx8/5Irb7HyCcuD+5vpRMxSwrbaDhIBSNStxGnHIbJFj2DxTzDk7CZ
1Zhf7Pa2+01cOfLqYzo7NlQxD9YXxChDN1crfEtHB5CYC+oYLRTC3CoN4ymrFBYm
uezlc8qbJeTmhI+MlxNI89FBeKbW7Mn9T8xoFDGWeLe/GnexeghxPCnZf46BGUVj
7K+Cj+RokDgxU27YM4tOCUIc//1uT8EMbzKBGYA1rn6FYDRU3TT275218hE9JCjk
I9yTJB97WIya/fWtZLMd7fx10XkV+x0UssKs1xLvm+/eZlKKQwsCdnmPDvpTfBWS
3bf+JD5V22pSr4KiawfVqsMXaQkSIjfDdr0sRMuwlOsuGd9NdQYtESxcT0bHLBjH
VWU9yVXM3uRQzoN4PYdKHn2Gt97ZDjqeqPJrN2/R5e8IIQ6cdmXg6BMQ+b4vOad8
Wv23CLqj35DR87zn6dsrDOsOjq7fZJL8P1hMgladhD92D47u9vQtMEwCSN3H9omu
dWxQmOxEMXza23wvND5aTOV15pRb4oTjbDoLRw6Y0pcis31LSoTNM1ZtFS0UTexS
ssrVYucYYLIhUK76v7jayxiNZYa/J6BtlDQPbLZwA6n0e5JuYxroMnznn4o7Ir0+
j+CVzmYYyum/uBRVLwx2eM0cpRKjBgdySeam1dj5DPgAFBMdHKFd5ew+f/VMyzU4
dA5xHyAi+ZhhdJUS0HMZc2Np9KaLOfUD7jYytonCCqlhZm8v05l+fEZ545foOuXR
qCeM8ZQEhllPHH3+p93EP72Lr0R5BXUKwB1XBpFkBwMmqpJslRUh/biETgqcdGTA
jrwqNYcALozBDO2xkKeJF1V84wRz5s+UN3hV820XXxj2P381pqzWdZJVuCK+pmcf
Mdlw3RDgv2lKHSTIEM+rNKn/VYguLCfI5mpC0Mp0JQ2/T2u2V1E85jZp3W/sLeEy
X0zZDOKQsAihk3mxKPxZmo59mrvE2d4ZRYHhAumTcVtt2ZrPKXe7Aa5S1y3DB7ty
N5alu2oy8OrR2LZSuCZGIDQJy4mWw9O/Ik3sVTfvcoDkDEJhsAt3SWuNEzEHlX64
Hn5Vcxm0v0DD3Wn6E7gTfRlvhNI0ZlgsBVfd+OeY0t9dAUm3jUPKoFzWSrPZmlMy
a47dNTdEYhXvjrwQd1cj3tWdCumQC8G/l50dveAifbxHKECaJf2EVfIk0s7ZaGJF
ckAO5n0CgDGbeqxaK2rk1P/38skoubt1aE8CI/rcfJkll7QYkMoSXMmr/84H0VNT
nFaR0l4sjDn4I4n0GxsStbdkE5Rg/yEpWPuRnAXmgBD+jnTLWGKyQe03SIebu8Me
fOmky8h6xl5WQkTu3eCmfqKbyXkKZEZ9v3jWaMsXYWbk6JM5zD6qOmVBkoxXN8ad
baOQtX5ZtkDUODqQBjtapkUiZQeviu6OK4CXHf0XCm+MMpY8Aa+aELKixQT2hdo1
KNcUpqIiAXmVTzN1aWdvW+vnzMTGEz8GUtwivTi1qUmIcBBg+tV+D/k7MIzAjmPi
8mFlKUpcbPAwLa6NPMXR6A3jT9wIoTmK2gjJ4wJfIXs7Me7yFw4Pn/SpIwFvkc/C
p4uu6JmmLYMENMS/7hfiW+W4qCL3aBEj3E2t/VfUdZ7NRhyxBM2VF+0EsYQUMaig
3e02Goo6Jj75RjtphXWvZM7rb50YEaXj/wFWP5KzGZjD6syA7oGdIj0gY+46HeMR
73FOBpUsrtGRpzIctAFQLNYQfaZmlBDEpwVhFo30gtDphPp7vO8uqWqXm83q8lNu
70Z0Q167JVYSfFdjndZqRsf7HikYvS/KoPWYH4KtdnP+sF/eEBHz8OtQs3gjhpFD
Bc4HGxCiZE0yXyWm/KVb6f+F7BFLaQZV517Jb0SjalApHph0igx7RjOv532lo3JE
CWj/hYoyvZYLMpWET9pAL7KCgO/ZN/vxe0U+vKoADuwjEogA5KLEhryuHV1SQzqm
IKJjm0dAZTCkLSoZ/4TQgT7UgFbUJQ1rbWltttr5/qSuz3Qce9vjgi3B4Q0uCtOe
8UCoeT52VCEkrw9SWVWlvn6BUwtNCMR7hYOrJ66R4JtU9PiL8lq76JyeEg5uL3e+
EuBAjy934SXwAXH3VPRtJtY1b6l+PcjOzpX9wSh7DIC0N6Qn+D/Jr2YpGBqocyZ0
qXpLmKlvdYAt92eUbb1sFokC33l2jAJQvXtJPfxdWC2KAyVLfHvYEcFxm95pNQyQ
ty3acCfWxmIMKC/YNt+48T/rHqfXeX5sSQS2qdzWvA6fhZ4NJewEFU8DpWHC07kX
QVXsr/Xxdls0tsdBYgMUHSBDn7bxratRXRtKHmmOngEwS/OP8PVJrAQcBj2laK06
lMd8ZlckNbRUz8jltvQ7SGhF18BMDo0if6ZC07myiFK+dwZK7ggy1vz2TTzMJoOZ
w4VAnuYXxulY2qyNFKBN6k+tG/WIfErSyPSav0EfAad2RJCmVyil6u5UFLkFM4Iw
80HNFyqAgnzqhGpUfKpgCMCRD+dhkAOfVrcxmZsPsmspHM9awb4zg8JNPIoEJco3
BCFsHJqWq4jnuSDEoPInSX0/0EYOp7QPzddTR2V8Cjgkfk7TDBs3kjK3CS7s1amF
jo+QFSa+aWIscO4KjWaD5T/8W6UBvESJ7o3CYyIvPMLd8v3snOY/v/KcTwaqDoHA
eJx9BEF+PG5+NwGBQ9mr4SaxUhUHy9ASGpvpe3GJ14s+E69uQS9ML6dI4THjyBlk
Ys0Bfme+mT+dHLTntvVULh4XETeBcPJIWamutzp6I5XYxG/O1+0KWAzTaS6g6hxl
uO7SVeQJo0Fua58XFfP8uwsTs0cpSSk+qg2LUJctMDbLHIvG4ZZzsFSGcjLO5n2q
nYgONbamOWDrxhLTAy384jRf3+CJq5oHx35/1VgWf1Nz3SRMsyU9sTTC4uZMtfXB
zvxo15atuNu4onWXLQ2IbMoUxMfAFGsFp0aXsK07OhMFkMf6pQ5x+T26qzTIFfk4
g9mmhYm4lxbIl6crDatYE+z3hdv/9NqikND24X4MQ98hqaNwEIif+e5X9DOAQYlA
cR+gxpZ/EuR5aQoL6LTjc036tMwScTUPWNsWuM+J6bma2gJVduhkWT6df0kIKr3T
q5C11LMn5OVsk522EFe6rie0p7fdVhNJSJmlY3+dTQceso6v+vW6hxqYYHBYsX0h
/fdIEO73j+bMf9GK+zeyWY/P7yERRfcJLF/vio1eop40xavSxkN1dN6se+QiBzGh
RhJdXBh/CXthNnnrLhd45vNHkyZ1D5DkSJkzoHUoHiX38kEwBa3epS5pI3gqI6Uo
1PUkKi2byuB9vu8zScWW/Hz0L+kB8kyMLFIEFmkN8WlOOggvRiTHgzXLpr6SwK5h
P5yelRs8N3Vhe+3gy/PmDZE9FquWIzmJzGKufgNaYi8jNIzCKIGQ/aLVgqpRDmPl
8yMkBY2ZPlprry0OIW2pFDHIrAJKcjCLg/V/9OsCV3wCCVpKL+tNRL2tVjFJuGQW
/PrGkaR7aKTs87OyXVgd48L5DcRCvQrvNlewRLgTdMfWXrxv29EdMnMxc0qDXTYV
x5C7hM9pbtaoxNwY504ZfuFb2iRPLJpcry12khSH2DlZHY+4LBHt2y/dpgTf1wUt
rjoyA9XAr5J7RyJoQMTAj4WU+p78jS0/ojlSmbxdgnAe2bel4U0CJwmGE8SMwVNg
jOutUzaxRUvnEW4ICskNIhjQbcj+3HMqisFoMdbm7YgVKizGF8eZik3oG0uzSQq/
zzGgOktZlBnSrP7a9GlX+vypSXN0SHQ/Qyllrw/Ual9c8aMPYV2cEl++TPVLAoxq
YVT0jpDB8gmpz+7gFfdDZYCWnP2u6yUARDmRWDwo74z/CVXyxGfwFuKS2RaxVm9R
fL+4HkiJCKY+yqnDOSnt/X6dYY8EXP76hbdjXjZEAE7lBsFibxntojVLXN3jJbC4
sK9/xheSeJOWlPDsTkgIqUNbhlZeceEhLAAbjcvzEu+e9vtBpacF2FAg8Uturgcm
xTBU4BUTtTrZSKU+NkVsL6bj80DG2iBJAKrBAwwfaivI85T5Agyv6zeUVR3hkD27
blsW10DKmCzwkH9aqH7VBtYm+pAqXGeepmvzEjJwWprfWc51ALbGbELUCpe8dBF5
6o6cO+fxah+1nCE0c9v9sHYAGkq5umoGdxwGa6+/INn6lx8aJvePFF93ElKBlaVg
vyd/30f9avyczKrx7P41kDnzOTOI2Cg0zNj84V0Q/oqt/Aw2nwpInf/zA5A3Airx
IJkuhRQchmHnYjzYuasqRFmIbH9B/YYjLe6Xyv8czh6C7YdmDKcT51Y2w/eZ1KsX
8+Seh7aHeGkLg6so4PgyvQPmlW5xWwceL/S//XeGkbOf43hqlECoDwM7v/M9eUzY
3BV098QhX+sD8JmELjtUjrrEf0iiNOKCA91gAHyQk64Lzk9OXxaEsQ08kK0yuzns
7r9kEn2KaJyi3QdF7FHQYo3BnlLkUkYX1bMLX332WdYbdCpImrtQHHYyyZwYIO2a
SaLJ3ZS5WW4GDh3l4HT/IjwMRVfp5C0QOyoNURlyDvgTqBRyLJGe0YVug02JxmP7
xpPjmi1ko+i9hbVhc5Xm96wa9cYyzTfBpTn/XaKqxjsVOr53C8FGL7keQQHtVVS1
SFEzGh/HP1hvTU+5gWl1V/gn/JMrQ1xrm7EicQF3gi4gub9+IyC0NFnRHWOYgDTw
trHhWgrPOLNn+Rg6rxb5XuPiD/rJOB3tgTkjmCJZZaTvI7wb9q8msRE5QEfO4c6A
aUGHZmkT0U223plhhwzjWBr8oP09JwBt+n/waz/AJpVXTzbreB0cewlHRl+WlIhl
Hsxch+PPD/i/qyDV0lCdPk8EiBCpk6UQ+BtjHjXxLpWtjIpA6yEYAcWCzk+DK/s7
QL78p6Gf3W8HOvY9RVPQsMToURRWMToRE6XU/ACotSsS+Bgk2+26ltnLqd/9WZ0l
UXUvbgurxikMVb8Nksq3nLGiJx/R4RhM9p9DuXTE03ucgqQsR6Ma3dYDI+kO4lfx
NjnRd03YMTpjULUvMqD3yqBt5D/GBSTd1LAdzuvK3GQDfI68+d6u3HS0dahhEqRT
h7RDdkvaxYerECiIvAPD8nx42x+6BboJHwmF5rPdU1DPtHN4DHRF7+IpVIi5YBj2
kxvpXbjaiNKHLJI042FXpgePTe6y7FUao2rDW+X3ew0lZLwciKI6Pq4+nwwSna5d
CUXuUDXhKZ/m6xjsDYwxifbgqnGypWZu/HoCygkmIn9cTltrzqYmzmgyD/1FSVyr
cqQieUvM8gKIEG2nkqngOsVoOKSMz1Sc1foiVnsFmk0/CVRhnnN+lL6eLnKwloRT
6975d15LJxKNXewSwzGgd5IDRvqeXkx+7gCu2qkBPbEBpdbr19ckO7oejKP+C5m9
ectBZd1Ry+28lzGcMSB8q9HbT4Z1/wpAWGQSnJtEQ1Rn9FLbK/D+RokNbQ80Pe9H
MOzEESOm5qt4J5t8SxXzhV7odheuoLCenoL5vi6f2TWvWgWHckB6PjtuhnCmFuWL
fAuZOrRDO/melQYYRlLK0zfiTtVExVjHW077VGT9tSRzqrXuJTx9X2rcJpqj8xbA
w45Rbwgwl5fi0z0PSUyCA+W1UvVvBCUGngDEH48fffTL/YdPZm7eWJZgYoMjpxeK
rvjg6pg2UDpKQ/BARHKBWgUCYnHCwFWZE39Ea7PGCY0LXnigXjutSW3v91DmpUKA
gTiWYakpIUNey3Cs7s5us2HnBONmdl8+FwKqTaqbzZSn1gYfYdZhOIEAfhs7Y/aU
Jm/MmVHBarbMA1I6jQleKJW0OedbyaYmvVHkEdcyZF8SaderLMF4Bck/KFxgYZq6
dwHqf/F9ivc5IwC9B7WxjclCmJ8C3r/kK6qj7SGIRpipP/wZ9z+n3Ssu9ZD1k2NN
6RxGYgwdUn4unzAP+GblHYPBRttRNTzP8b1L6ck1KWW9Jk+MR511UPDM9YB8++6y
d0a5E082x5+yCg9tqhsw6DsGyNYWxuJMAyX2kIdlqKg/hWreTepy+GuPKtpemPna
rSCRO2q9pXaysdjRDlqrlqH8USz0u0q2wAEh6uzIaFjuWfijAzop/KX3w2EEblYk
hGeXweD0NJLF7+sD7/mQWXJUET2Y7A9iSA+8g5XrKZi5HpFReFRtF76Iz3ac8LjZ
IwhnfItqVZ/jCsAh7E5gUUxiir2YPoEk92RhUZi5QrrPjRlOAoVUfwJmPtHpVlTw
lqb/tvWCMPcM8HixgDK0H2/yTlN/rC6DTEtZAR9bDCuakFoDXORqkUtEeLAslDZF
m/rbAmR4VMv8x7Cas5ggOrvP8kuv3ynNq+c0PVV1vrgskB1IjcVAHejSpSbLeVtv
9sBUlkhr+XhCfAXlq9cG5enW4zkQk29u30z5yGFwXxxA33mxZfI3FRK2b0TxxvBt
bvi/8v0PzpE9UxQvteLrIpBaicMr/zBtDm+wL6gAFBMGT42DT/zmf8SkgV21wJ9J
+yBRJ8Su6Dz3Ns2ylV+kmRmQs9EPj3Ty8KKrj16os4iS853Q5kV94QKu86eDiCK2
pXoO34lAA0G9d84UkyQNDpz28VjaOQTYBTXxklHtVq+KC9prPy1RDg6ag/BDcI3J
DZdwTW5mWidoSiFlgklbGy0XZ2VhoTUn77Xgbp8iYXKR8FEsQBGC7MrBTys22vi7
SZ6Nei1mccxRUCG4v8sem/fLZWvb0Sv8eTsnTXVA3cyEeZiIidSRz6Vq3Tzx7z4L
qRb7p+oJSwciLxB7j61ilD8j9kSR63FUKWYDeY/H+LZXLEypMCzkvPpTNRBXpP0Y
jHTK+tTPbmVNHr2ckRT/2cOxrezbY29OgZBUTXOun7Qh5GQN7ISUChpJHMwhQ/f1
pfu0IdlS3D9OVDoiJOnyZ6T8JQRj6AAQ+W1t/nsm8AFEu9prG9xUefqwyIgmwvAd
6yhxZTdUC++XpNHD26286UoyeYZbC0iM80x2HvnaAXyHUDZp3YjQbq+BJHjHNAmR
rY0UGvnkHqYM6wodNOUQD28wnM5QyIsjgaGF1F89fEETayUmw2ju50Rrrla+YUHl
zwbXBPCZOVAlWp9Or/HsAn/m1qaMJrHqJN9s0AIkx9K8FmP3rl8I+8zolMuYERsP
K8pRaqBLm3g1/VksYvD8vbHYqLfmGj/sw8IU1XiCU9ZzUOiKk+PFvEaJCVDFLHFT
ss/l8kOqPbvi4dauj0HdnF+dHbgeCv5oj96qK2dpraxehnapaNT3ANC/RapGQ/4c
lYjZ+QBoVbZeADcH04LHTxMU44Iq8mZsQWnKVFLoKiOiXi7TBgr2etQY0gDKQ5Ib
/SdMO+/n4pV8vscnDibjNtTUx2YpaX1c7QXZySmjNKnMVYYUUQ0p/WGe7lsuP5b+
9bl13/23oqxTmElzK3WADnHXagIpD+BXtfMUasFuUv2jjNuCRAZmrvpI47lvifJ6
8MURJPTNWsNj6jDDTjNGw7Ng94yBviVDIpsxScE1hd+bAUpye4SRKEL5lVFz2xTs
c/vKjJnmIBNwEa6JRxSnb3G6JmA7+V6od/BOqO6G/MiH7+l2N2VtUJMfm5OuVoYr
e+Xu7dqQTHR+epLji50Us/0q4EZ46s5AowJUuCWcSoJTd5QeIW+++boBd7HRPaiE
KmBVuBNVMoUzDmQhbdfYC8On7ZrxmS/S575/5HZsHS/0uYG9DSpjPA6uaCqn2SQ4
U5MY05NEkVfa3q2mLakOzY1AYV3wEKWYcc+piP45s3xL9zkW1wqHpDCH9enF3GVh
RN6hpuCdSd42qnFxU8w95pJaio8YS62uFTJKZQ8g2Yc53mJK5kVduRhlgX6uIShO
Jl1TwM4X/4uxSG+0cP1sHE4BNhQADLv/kkMGJRuyR7tq7Q8+rBG5Y4B35Wjza1Ro
8bwbsRFOcMVIWEGch2+h0bXEvPMKiDrIXuqUURs6+NcT3LuwC9dib8H8ANmsFdlf
Rj1DL5eZhrADF6VVcrY7GA820FJi0DE2czEIoX5EyZs3rL83/5eCGROaihgTJizx
7rAV92X8X/cZgf1BYE6z1xRAQ/l1u5ijyLqpknnZfizCa9ltIqLR/Gmd+/F5hjvB
PFRxNUbeEpCxXsw9wJZiJQla2X5m4HP/ninawnnSW0vbjBYM8nReSM5XGlwJNYUU
J/krgVj2q3BzJk82MAGEOe5Z6UD8CN2E4tv12xwIoFEC7+XFFoNSJJCV2R+Kxc9B
ktLKOkpJFWZFvxEySVxa78fgvQOJ1zTNpJ5pb2k4S3jyEOkrF0eVl5B92E1BtIyw
XAOvJg0IeaThg2hm3EgWYXrRPF9yfh0SByG3cPonmVM4Trcp7Li+YLvgzBirXaq0
+uixPtZxDONGunI/uwHjGD5golV5Q5IhK7BCZaLaG9sG51V0/9aet+FLrrBKgFVx
s0fhwJ3zczC9afFSl6H+bHy5mzkY/yEI+d7XcRwXku9jYUi1LyasXwRO8J13/RB/
0XGqN/ao3yy+mfXMus2mzVH98BEM7AIfdXY8A5yxFM+wGp4Ur1n2x3P4UgK56WEM
5WOC3WFAG63q7+cKPr/lcdAe9AbYZYXXrsDrf1ZtNeLI01bt2iAFW9S2qOzwtRf1
JRsZcjxlOLBt98xIT0+pIdL30LJ6IJu90mQjx0MfMQsqWElXTBAFunNTjupcKH9O
Dv3oumQ9C2mn+x7g4Gj6OFrEk31Jd3jpiZTBdrUeo50HHVeI1hRJEb0fnfRv3dN2
FCHFI7EAIvy0bPy1cu+W6+COs0MIm4gmYmpFzKTWW3T8xu075xlwr3B1OU/8zTbw
LfqSVxBGlpbA5c4GZRj1CdPiIB1qpFzzTDt5Ajl9XRxcrsczM7alVjALdpyioyuF
e27BJC/G0nZiAH1R/Sddolk0BJoLDgFA1/i7UyK4R8llZR5XkW5aRn+KwwITh/gc
6eo0IvJpt0bxI7NLp3dC2biD9Vm0p95SFz9wE2C+D1gYkDRn/pTJnoJzrDD4FPS5
6Ao54w1vC63FmYILLq1tcd7+ennJnvfD+iEGrl2nYAU1jfFDRu+4KED79EAsjIqZ
Lzeo4xZfwcTeFUDiQKFcAvvxAldRjE4hP5JKIoHBWRkfLzr392R51oyKmaYZbaN6
Sz6YQK+Abr1YZHeaC7RLO8Pb/wBF28zwqofmGbYsysk6SzRs+Wi6P/H0POe7h0s+
p0lJU5QneOrUsxD5INowX5VQwHneO625VPTgR46DuvBqDJ0XoOpSnoXJEw2ngKx7
W55PmAHYN4dYtahDFGSFuKEat73lKMqY4zg4YUEs5ky+vZFNaaBph1fl+qhwZ42m
So9o/sN73Mv9NflETy2Ie0aaayFqMcTQBrFbDYog276xoNZZx9A12wm1xf6uNQ9x
TmVDuo0eybVCCTAOENkhvuxgNJPslz7/RvaRxFeSElu7TJjimj4cnUOIiLQYblGw
kinUyjHlCaBVthDGNbx2839Lsa2yh5SLyrEzRNxzBK23gWGWbUU7lI4+a7PMSY3N
qyzK5qHiiCB3pJa/gmCnYNbOFzUP7TP6BuiSqcbLz4Qy75jpE2SimugRQteiwVtX
oNa2HPcqZbrb1bs+oCoWcLGyd9cb+R3pYeCVhUZhEqH0umDwMUyzrBb41opR7jTD
Xby/4L78DWhAimguYdP/Vo4S3y7tXVZlh5Ma8XDPYejKtdkPj6v2Syc/modrH7xF
EFfjwI1GoArpBYK/Y/cQcQ/yWFunxWN1VzVG/qQuiV3IyrA4x/DLGuy0c1e7eMYp
QmDNvZCY2KDezQ1y8wTNccl8cXaASYKToSQYoebysl4tWzKNQW/kXR8BH6q7ySM1
xzZDcVhJkv3HoNCpLNg7lpot6CwGd8Y6wYLAYyETGKLy8YZgfwsxXT7Ec6/WuuIv
9SLoFOXYf7PrdkUN97Pg0uWsPcl/x+l/cm9DjORwysLg7ywkEzcgwV8HLEjFIyKk
UKxiPDg4qIg/QKOmjHFtRUGei9+aFsR+kHeXgp16/CHl6Z829wj6t97TtS15sG7N
IRUtocogSDbOLirKp5ANMvhnwKBl6I8wkrn72lA+djXenybajovMbNG7u6C1G1gT
TfgI9kmt71G07dwUjrfKAIFYRXhXe8toT98T5hSdThrEyoSxLNtfmitgdokaaI72
+GnqemGvrXU7ls0p4UMmGdSP5O8IdOT+Tny+zfNNCA2qkmDcRozPV2371d0NTqAj
KHef8gScMY+ifNPnwoPyVjw5k58L1Ru2f4HC0BSnyDw4vUAWJmwlN3hY883w6+YA
bTQ5yphyLKJJm58S9Q8jXMjZUAxYbu9v2WavJcshDkZgKskjAWVvKZKftlrL8bu6
Ps3mi0FvI+/BYf/5pZ6JfFhDO2iWcixr4GOJRy25xUzALbxU6LYA9/S+jmMB90TX
1x8bhQpPFpf84/LaCQns3XCuAm5sccHVRH8Evulu58eNbBJdjrfAJ3U3pbptg9wz
B7IbndeU6CX7VlDMvlSl10cJeYusRkO+6yrJPCPVbDi6NfraAL5HjJCUeMt5E3XS
dWz+1DF95u+TDJpDz7NZQOELXPxEjcRqmokCd5jdpO03AB2UH/Vxyvh6Zlyt6ttD
rOOmc9tmGTGzmE/ZNl0gx7gWH0cjKX1dbGQdnApelu6l/cBvdsf32Xpu4NTq2hx5
wwMpxGQMO7YR4dqFJkOB7Pqn4ZAnejO01tee9ooUcyUNWNk2ZIzGg4S4gZSypSx4
R4bAhDHOUaGragmNzljrDVbeeU92vtUgovJs8VY+epP1GZvaPCi2bfcinl3lKPGy
KLOe+IgPpjED15DZbgVbVCZ2x5FcQ2vTo+uJy3vv0Btz2xENrhBkkSxPK/BBDUEv
cg+nl6syzZ6btsOtzU3BnLldvExNIQ/E1g2J+9de42stVj1TEpAkv+7enaOdO6Vr
103iVsgTPxuk9e8MaEe75sMEDq+HLOS6KNGQ2s0tGF/mYOQrW28b63ouwnzRptXO
5AL0IQwD5uVK0BdDZ7PHxUIJQmrblzgAHG5FIbIjzqgcdisJtbaHZ05HxkwigiBh
HqZcCXcppb4thIrJrcNMWy8+Ldlzi5MOIDxHKHluMppiLvAmSU9QrcemWiBKuuJA
unzjaIQPvh77JerT9bNVyq+7ExfZPSjBWQZoKkA1QIyo6Ge/iavAkI4ilHJzhUEB
23j+1zMqKtOG5w/3dnD3bcn8Q3IHzgOpcLvqM9BBj9dlcc3k3CkfarCo+kexCfzi
tU0JbCUdvry1CHzcTJtJWzZY35IQoZRvNBoskMm+jOKp00xQmgFIrpadshZUm1jR
SFWpIhsWg0zT9TzBeGJCZ0dx6DhUzW5GAuzjMn75u1cH8kKTwwS5VPiecBnAsw5O
LLDC+uuakggL+be9yfo4Sc+s1aElmd0Ydm3cWG7fQyZeJDungfS5QcuxWFMLF8uB
FTxwayHndpqTPDJKs7Td7sZT81MGD+46g7pZozm1JBE0kSqcNoF128jSeHnakYWt
K+6NzcOz1DO+niqJm6KO/REKJrt5RH7/rXSK3mmJmjaiIcTESRz4yIZdwoiIDykg
Ra70hsTdY7Qbd6NaYaEnQZx6WfI+Ry23pmJJo4cZnJLnGoLinsak+I9Wb5T3OFC/
mNYd6TMH99TovCo0xgMehqWtHOK6ufYXgPbcDLVik20OXCJy35o9ohPO325OThsW
3Kcl2cV2A78hbFYO/R/QcLhtM1uDEb9uMU4czpMgJ1wDrxstJ7NfdrtMQT2SRuKT
timIKwyXdXXjADUyg+5Nf+wWufaSF8Wm2k0VfzPWMsMsowgLORo4KXfqkWUtU0dH
RXmAZdqkEZkc7sHh260X9BM5lt27z6mNIQld/HNVa+A6FJDi3Yv07MeTS5aDb/o/
OnFB3P0vNuxdmFn0rs3WoY+4+X0rhNBcfWwPCkx5btwo/zKGTyjzdezJW5on+CLe
Ys+HEGn54riZZOn6K8DqB37sBIf3wq+hVighr0dtaCvn+WQkmoLUetBdZnQ8sAd+
M/E1hbzkqqUeNXK+CIsZi3GBmCT+iQEBek3cA7tRuQiKnwB1Y2FtO8fM53P8TlWD
ZC14yriKN+ryRqIL7l8jE4LRPeNmuw1b2bN4sjq9CmonNB3kanZD7jj52YkKABg0
eU9p+z52gCkjpSY175mi4vgpU7vzV28akym9O3aBWOy4cLN5KgGCD84X0JOLUnf0
cYcv8yJDqMsQCR3gJ3j52gDmRUqNs4ORpeFqYviCyCSMMw7KzPShWFg4Vd4UbckF
p+3NGPw9ZKSmE8dz17ljz1OaEdRAU/kY8i+IXrDYrc4nOkrjlAgJiSHJmLYx22OF
RplOv6Yi70oObiQylISJxHh5Qyl8iwRxhK+XAYq8lIGk/4nY574zUXAdAK/NQdG/
GQeUYQUeGhBj0dxc9bqFKf9BxShfsuADNW7hxxDGTT7NvBbX9rvlt5t9JXGDqjdt
HfIBh+GfZl/YahmfKBQlNQWjWnbq5ekROuxSgSP8tp1ITKn+nXrV7yszuVlMSoz0
ruku0ud1/ZGEoyrFLYSIMbEqpICyyIc7gmgdsBRj5z79YBJ/Czd0osWIpPVS702x
QLkshA5m5QYGBWxKhiYQfiIzwRESGmLpRq3KH9Vva0bj9ow72hBAYcl4dt7g/Wni
sjC9khMMTS5nEIwtAe91UMyLK8UEdHfXvySrW2mr8C6Z5KjMA2S07njSYrNRYCah
ym7ngwKmz8nIX4IRO9feWcAGAqv93qrsFz8Y4YMNiJqm+AuykLSxSFLYXI3ihUoB
2J6qI3SuK8TaF7moM2Iqy+A0pQ9qZfNLmZPxs82YiStHdizez3S9rVMTMA84jLx/
6HW9c/pofeyQIsEegUfVXFumHyfr/KupY6vOwDQGI4HJqRWy3qPae08RJzw41iRU
Wguj+RIPCyvk9qduoUaJR0eUpPMV5mvwvm0B91gv1TfLrJjorNaBqvrYlWAwtVnD
h3o3JFsvkwVtdYjj8yCOYokBrIjo5uvgenYVnGWPZKN4kJTbPPTLDjNTqdW2pmvW
ohCA1SJG1g4itOMLJpAzvEVIYL1C0shmbR6vX+tvHSh8zIUgZm6tEAxq4ZS5Liiz
wnZGvqePpnRZxX/T+g5b/JYjNta8zMKmXdkxapFqzBFVqHamkjD6v9bK6aXwhT9d
Ee7nn8eHchbyInhnQfUNZRh3zIyMSbbQynedZaOWKw8AdE/ViJSivdVC45IbIlDh
gTSlXtovH4JAV9pnS55PQwoxUQ6yNXY/tsz1F8GbPuvZjx2QuzHcGi025j4V6UjA
/tjPYFxqQTAx9/sXX3p8/w7PNSmWsKIXUVtxtHOX9I4s/TMFxVk4O4CUvjob27TW
B+geIhMfikyUp0KIr5NGfhZVja29EHC1l49MY4GJfuicuxdxxMCw0ar9o0Uzx4uI
L62ar/fbYKCfcosMjtsB0CMwOu8lRNClXJRY8DPBMqmckM8kg5/ewVIvlwdzw5kh
Z70bGZ70/Ku7Qo1HyybDr9h8ypApVt42urfWI2BwrsA9JVy5aZjRdcb5NLqaSuQF
RwJBA+/HSeVIFZRnoZlARJLEAinybyOJIPOel2zLmMSQQFh4S0OFZxAXGjROI9IH
x9GmY9Qx8hLw3oTygJycFA56NW9lne5Lk1DiwHwXZErOlPP/bJmUOi3tmS1fOZYQ
wmYvAJ4Oxp4R3ZF2tietxcdg+2yAZU26mqfVcpYTX5l8R9oUQCfb0jRu2d39FHgc
WFE14Z8SY/tzyJYAww/SU8+gRzhlrxEgJUjp9B1Z5gVpaNBzUOAgb8gKDrKN15Mh
NnvlZPK1h8G3TUb9gFVsrkt136Y78UaEP5KEB1d/WvIpmTufPaoIzzKcHiAvwUCK
hTbymkjTZF8zLY/GXfpZHwt3zgbK2WlH/HZUP91baWN4UHHjNFmx0NIpAqTqG4gK
U7zFV0+35/+O7c2ON5SdZY+BJtChek9qJFZBocpblb1jBMZ6FBgnLIOdJjjAlBWC
c/MBMd6fRgHi1oUe2c+jiQWw5LtfOnB3eMCFrnf/NSjKgUt7y6TFHjzyWiODfdkk
YWMgv1r4ELhPgbZRLJFkz2NZtBHkEvosuITx8haeqmWZiHlaU/36hXR9Ttlg0Idc
vRzBrjOmx3lGpF8WVivJH2iyU4KX+ER/Rld+eSkYpXnq7cFzxEc6tN3vV4pK8toN
jp5US89clpzcVy6TfZ+ojOfjjBpfL3H1pZhVqB/NyTD1+3vGE/JIHWNpi7LRtd6y
enhJJJGigMefGK49qVqIcBRAEdzrZaCn6gRsRuAjhTDc42XKPFHQb8KukK/c8XOp
wC6rGFhdauFKuFgFEXcIZ4R3RanyfWR8HWh9GJFWDvQUpjT9Kv8t3Tll3LzMXzlv
8DG63O5A1HYBmLt06nkMOvCo7u7bdWvv7MSXAsxdNyRmjrYD1lXaFCUGD/4EUVSE
bp+cwHdE5HLC6w6EbbYbXJqB00SUwVU0CP80tKKOlraEeq7ZBciApRC3YqE6JAhv
utCl/DxHB9R+ipRiSldzStpfaAD0EDe+9w3z0bsGL0DMOPsUaq94SF4YYw6JhuKo
RwUBEBZ9dvp4TH/E2OqTP1YKSeOwHU7ZQuccQcwwvHmqqCXYhrucYK+xKOHih9Ml
fHzjoePKfd8XIYtiDwfBQr4DQGLx7U+2azbH9vK93Xxj6FbACPt2fadaNE0M5HnU
Iwc0ShBnbVeWrl018lxiuFj1bPU2uo8fqPgy25YRoQPUL/cf4c7VhmOohCRGE6YA
/IMPe4xPjhmK+Q+lKNehwYH8KZsjSkaRGBzuWUE/zONp/8kMHanTkJWX5O6Ra5eH
pCSC9ChZhWJ98RzDaqjvSpEdxsnE/vwhMXzH2LJEAEnMrjFTgRoaANF5tB+UDiMg
LOrSmaRQYLD5mTQNHzSpYA70NbSkBGvMf5V2DCvM1qIDSvsi9rjmswxLD1tg2BBl
fmYfxCyplK+pwGaxRscLPbCNRhDQh1wqXO1tdg5gsd1v1kwE8d4m56a+TW2EHlyO
DbM6bMZtfVDoTwqO9Unw+HaBv9ZkhPzHPW5GLSQZHjJor+4qcoFYQml4oTSePCS7
/8UPSTJHA9OAGfTD0hDM2zyRJyJfjDp6+aWSYB49+W2zSVpdMloP4bnwIe5T6dAd
g4qY9g86n/BXg1gxYji+PtUUwsN7MWQBZe+C7NJ0iaYtQGY4PTasE53yaz9s3S+4
hms8K+g8eFfweEMncQ0KHg6WVgi5uwS+u1PWpzlNS2dMCAfY1soh18LhgCIo7wbv
JvaEnKhNzNOqeCm4HBzHqJJpvAmYXWd3CmOLhYgeNAzRNyX+qulKDInksC5MNX0k
BIaGdOhnnoNkY/AM+ui52fQ4o6tA9Dl/oNHMPZuRxIBedWHxBrQWSHVoXemMZ0DH
ZQHLShcQs2H2s+Lq12cE/38biDAd4VY/kqyfHC+b9UBEn6kHRwGgtX0omjYLme5B
/xnILCXf2N71inkncj0zVFlxWpxoSkMt8yZhhA7BuBL7GO6ieM1QIiha0e1FFNpI
RYsCpJafB9393mTqUHXx7bzcFLDg6CdD6gMYGGvWoYMX2yLHcwy9m7cAy1PtlIya
P5juzDAl5exUr4slXhh10DJMlaVWixuIxTLcyUshIw137XqN3ePGa0e+cvZ5Azvb
iIK2GshSjVq1jq8GmtjrJGbZNXD0G/GF3QVzv1eOQU2ecFYc4eFoHOZbkdOWg9vh
N8w6DMEPjqJBZN3uLk9MmCTfXeYcMe+ykWH/Vai3PEADUJYTINV1g1mGK0Dci6DC
fSGQFddnX7i5D47Cx13gDD8g7OCSr1emr+jIdQGml8lCeSXyJ/qTALqM0O/ybS6U
xzYo+YQdXbsAp8s0qQmiPGXXWdgsew2cw+6o1rq3iGoVTTMBiOxr3ZoPudGwvB7J
RzG3dz3TnroNhT6b+QkNwfj1WYenOGN2jKvT8tMGK25h5kkgA0Srpqe5xdrJQc8u
0RRAb894tcwSHJdSiUMPydpDXMmzabiXVNDr/yF9o9tJXunQ/VdafFtQUjVUdz4h
iBrNR0kdvwpsEs3M2SjOGWvFq5rTmARiVbRVNe/kvoNf7XpBvfKF+VfD+lUcqorP
Lzm6OSq5RTdEVwdJNO02+O4s0NKsPM7/7SPvtTynKUVa9SfBNa3xA42+YDiZozfg
J5OjiwZhqq67ZXDP/piP2T5UvKjDsTqBBOeNVD7PN5Uc0AHm8zXxInT8uYgQE2se
Re2A58f/deixj/CViC9NAg/BFtdJSSEOw9k7MB6f9OqL7QPNyaSCfOOKBVXzx4ze
O3oVNa/0ZIlpsc+fVZ9yg2Hqz26DERHDY9tzK/BrZ9EIGtzaYGE5mKtH6Hu+XuEB
Fw+QSqjGG2dCdZd5CFE6s2UgaC3bhgTbEs7X0vGyrsa/p4zTFGFFp+qgydcEe4t4
/kCfvBf9qzTqzePNK/TiZLcQrZAY/ki0843ZSQEX8UUWtGU13JNkgnuxYQtaH1p+
8h6oQ4bwysB/TRDjQFpl0zlOcw+MVk3dWJXdMWLnJ/Q40yQrx2GQie2TTsAM6pb6
4bOPN17B0XoH0Q6mPSxSjgRMWPk/EVEFjL36RJaBVi+1vG49s/z2STSjbKDTxKEu
3iTW8t42eZpT9UMbcG9unUg+UL80/84fMClbJOt+oiy5FNeHxGQtvnXruox1/AuN
fM0cxxIHKYmRB7igrrZeQlwkTX6XatxTyFrkNffT2QGGS3p6Ox0JQKP6w3rO0nm/
Lx/AE2ZFphqvBh6GX+u4SahyL4p8kKbv+GAFO1mWwKVwyCnG9boE6/by/uqCHL6T
VDSOHKGYa75NBjvKm2+6LCyDu/0BsR0ZEDVvHgUJhBC6pf5NRXvjFmUTIZ3xJOSl
X0KW1TyH5QCoc8buCa9MDbXSHcUXSe0VUqTn/Ei4psDsB7Nr+O6z8pcq0AmHaqYR
P8q498TBK4IQao2ckC2ibddXtoMPA6Vv+ZTdggTsszuq83wg80G8p0Fq/+dNWNxC
0l01BeqNzL0FvSVVgESkLfqLV0AyK86diWEI4zY3LkzDfjeujdnRyt5zg7Nfvq42
JIjyean6Y4PkJkBqqHQNGiGzuEYZZpPFMd2bIh9h+m+CnYFB9egSCOOWiZajyo3f
yNLk61FIU5JQboyg+c0j+qMqOFgnKod2CGpJ3PxPBUIeEiGrNIqHKuQ+B4/WtDAO
kM/KampwFgUH3GPZsVBZGrbG2Y62/69WuNKnjqI7s7btWWmoVvVboU+96Ccfsehn
Lot8LaaGpYSkQMeOb0b8neymZIqiZU9XEfz8n8HoNt1QORBAgtfVYNEALuAcDsWy
+Zb1o9WFXT9phQC8zQHtDcr/sf5mlzv707mvXqJtPfkeX4zhvE+u7VQhauk/suq2
p4XhBaKYP74DiQaMsNMwdYQWtZ540ZYUeRqpIhVd6pUBngbAQkhG/82lowyVjPE3
8QEWCAbcIRkuTqYXOhNzH1V5fAc9ifIiOZNn6SulBMl5VvXI/rZexyu2Zdp4H3em
PD8K+wEyQMo8HEKo2YCfxL2fxKVrMJvqu+KvNoqZQyEYAA7mfQZFUmxHs1uuI0yZ
bZzGSD3cWun9URPuwCfs8fWzD7Jfad68lCBdYxBU/Xua8mki5TZ5tXLtQEBH2gRW
DF4CFPCn6odV44v3sj5UKg851ejovWv5cF40P7tNVhtWF6MdBWvQpY7cVvnYTS6T
t5HtFFna+y9a2OXGTGNiKzxbBKKyk4KYmJmiDEmzCIknxb6ju82b9ibB2mwWvo+F
5rHl4iAP4sTrHaomPSt4K8fmtt7sqJpnimG8jFRG8LK+tre9NTz8116TR7OYas05
gjgRGKYBtW5FLYV12aWYkf0Dx3ph9DdUBSDnw3DicfjA5SW7OqpYMawruUWIVJhg
EiAHSHaEyLBx/u5GxqNEYQ3BRyfVLAfbI6XUxUsa4cscvsCLltGHcjhtTsxZA5gJ
TRsi+G6K3ckIkvlrSziPjLwdkEFE6RhvfJUe09UVyMv1ilIPHNx1SxYoowA/9n/r
+zP/v72ftMqD3feut5xf3j9cwZ8xxzFA3clP5H76BUhpnM3zu9iLR3juHvakCKu+
ecKAzPb5eVVmegbJqAln0mBMSQsULkdx9VMf1lU1cjgH9V4/3sRgLihK8D9KbDrT
IzcCm+ODAvnlMEWyUu0GFOb4B4Kr57T2eHs1YHX48N+nLLkZ0RIqgePd2wncphuY
pef1hDQE/FrB8oAaBnl/daMMHZawfqJBTuqdjaOIo0DDDYT7lS4B5XUms1woqCZb
TaB7+AC74dTfOLv5e36dyfGm3+nqIcge2JJIj9peIFItf39oFq0EUdmd+PCYvBbB
AeCw7RZmybxsXtUYNRxuBM7yyRDveS2dsteoMekpkgDFOOJMR4Ul/EK8D4U3+rSj
UPe99/3IdjYFjk08gxIRoylASI4MXSLslU9WDaImY3G3ocXMBssOBZAViGG9cmWs
RqKN+MzymqLwsWgsJfXzHTEMynYTiQmJX/PwJIdBXbMwk8B79YbZsplN/EqTfutr
D4x8k/Aag9tuzqD5VKUnxSjtZVwtU7w1lbVQ0RlPsBODQwSgCZ8/fB+jizkyqyuE
9a4my3mNA+eKFLL8ZYS7ammzyZndP0dKxhkX5XQC9N+JKG+FRNTH28E+3oWYivKp
ZRNFFoY47JYWNDHOSNeIGFJPftFEPgAXlHX3aVnjlf8oNzVvxWFE5fIYjyQKkHSK
VO3dbhPDWFWd57NLfgr1Ngp1rvM2XzpgMP/PLrmtJwH2EMtLr8JBnT1z8OQje/Wa
4IXv6vraWk2CbpB3kYWdzmUn730wZ8QMwliGlcraPuiuY+f3bbtmACl8Ig9WKoDv
W10x3RCzGrIia/M4PnCMWtF9SxMNq8N/5rwugQjJvgaFSwC1Xw/4QxMkFHJaT/dR
lk7JS2aFAEWLMYELT4DkVfKhAWwTo6bcf4xmzKfmErP5VnVQqkLcq4pU4VMo8MNL
rO0xKiiJGEPk8GyBfPUL9AIJhEy+9D7WNjGRrU8+R+rKGtkzL3szAxgbgMoUofGZ
HXQ5wzh6atmFrZ+NnZr+PN+N7UBmpg3/ehIK6btC4vyW2HpWEf3Zm5C5K3xfQ5DW
bNNC+ma2Q/sDSubV8NlYXukM0GPPrAECTH17c+0KHGy2NE206I2liI0IhYNNG5tO
N4DAoeM7ijJhRbxZoEoVS7prZIpVp5Le3HqzX3w0tk2j/nAErdRnng+/J8n2kr8o
EPMB+OJu60pdF4ttMmD7pUPTG3y3skqr4vxkpB++RJ1/n2knd7WmtzMxAzFZK/Ie
ronNuWVVR8Pz6yvypgBo1MJ6ICitsAyz2oZCPg3+SZLLTV2niNmoCXdvMAVHcAm5
Qo1f4SWrzV3EaOzjralKEhwV3+MKVUP+VL2Yzzwb+SpLQBuBbcl0eqW/PyWdcc3i
B2WZ42ZDI/kT6k1CbyDC8qt+JzARsKswGoA7k52rJu+GRio1CgME05jKT8OBR/51
gWUcz2bx/7iQhLOgEno52GVLqfvHB+pLgsnsd8pLZ6uhIf/xGArAnevVYVmceTUK
GRJtci8UH0OpC0+6I6QWvKS0XDoNaHrRk6lFmOyzJSx/B8J34AyNUlU3Ki/s+UQM
HwDfANKltQSreCvVxqrilHj0eeduSx5MLBqOKH83UG1eFi1Hm0vaN3BVV3454jGW
mDeaszUZ6BgDVyxm90RYuONshv+Z3lR9dxuXaSIuzbzbwVhpPMqpj9tkK9TnJBOF
FyPDvjIGbDFZ1Mpz2o1o7UMIC1LNzRArg3dZuwTxN1+A7iMduLXdazs+mlTBJsrz
gGhj8bah6HHVZuroWIFtBX3+K7bJWPRISCg3a1n/ybGJr3gjqB3I1UGAV4JZQw1K
UdO5Jix5McQMMMMOMZSl4GQJ9i9ZjD8Bj/ctjYa4lwgbxQVmPP49tF1V2dt3LbFB
E17ZXW66qjW18egmSE7I070oI21Yla3rfC0ZF/ADuPU2k6LdyDJGoNfSpKHpbjKj
UYdlZgvEaxjdmMVYv3LEzxubSvAmDd5fV2T9FO0M9xNnh8RvkBAa2oAJqvK5dM+J
LJ8y/JXJOuuR8UM/ZITFOugdLLFJ3j8HvQzPdEDyczIj3VdcRG6AqcrtaERAhup8
rC/q3Nq88bKeQnsxzAbsOOMrEowxk3uqWGatPhX6X8xKvnflB4IqFfkG+IpMMi79
7Nrz+MiZ+v3JeK7CSWiFPkWW6IadxNMKMwFPhjQVg0A4D3FE2EzLyFMWM81zGETb
TzClAbOIN3Nxu/p4ZD7XnZ6t113QmMLYJNcemB9+G69eI4MP+aMbBQugGg/d1XYe
brSQ6a2IrMm8xxmgxtctewoDWeTjn9/iXQc7Qh3KmdFpv8ovcLqxKyjL4Yng7miM
YhEDxlsWWbY6xrbC9C97PufM1PSwbflwlu3wraNTzGYB8TCAw8wj0whbp3+uGv3I
Zmsz5wJXf0cYO6FVZ3oMIYZjIqT3zd3XrJ/zf0Odqv9W8QmlYMyxPJxetjarF8t/
qHRFV88afUX7SYocw44TdXOsVNEKqVSzSjGhuaQyc90NKzlvTZ4zk57DzRIAJZfY
TU46ll90GTJupUiyMbyPVgNC/FQwg8i8HwMC9dAyXmLRnCmjR+UK/tRg7+RQcgQu
YNQPnJYqJXWaz7hdSrMJa0vguaIXrmTvj/PIUK8JZIzwZz91e+3wQokcJjQKhwMO
59CLkr4wjlYZXVxo4/UaOmbvMHQ4IJi2IlOrzXlLi7A6DfjHKfXKDt7cEkbkoUJg
v++qU8LPLx86mtCczZn1uYFm+/PnxZdLx1cgulpuXTdI0+/NhEJISEs4AHlli3hQ
vzXDxPSrVagvCAYvodKuLPD/IiT2UQV/mbPDIl3lEHNXeL78a7HJSbNeSYLdR789
DBN7dQvLu7RSrm0m5y6ld7iM7LzPhqvDPh8lW7EU8RXmzs/dLfXMbgoNsHRZx2Bz
XRvqfp4c59SRcJiuRDBfl8/DDu4tETFH2WU4BZEDW8xbrmungNYYb2dlTBcLDM7f
0F0W8ICXWZuv77OqPYdlvUaQAMiwmNtjQqqx6OXWrKulSfWNyP3fnaMU9ca039Tb
j0mMFcMwPU4rbrDm2wyzwsKnqh4MRctRU/pd6PxNJ7XM5rjcwTukNm36jj/mOFB1
5AqgI93Pdv2Ifn+Jiym6z2d1QlglcJHwo7sSHPr6ibogOxE8pVTh0NeKDca8+Ui0
JYNvXhOCe6qbfemtEIsUvATvXLmGR6caAf1MtRQ33LVxF4XwxmZFoo/HZt/xuQsH
6Cn6ToUA89HnrlmyzhuiQxvRD7uU8TOXnBPBk8CWE4lhpVCKKuJ9KyARs8rZbJR9
+6YasFPcmLXH0ZNm1HpTjzGpq1zjyfrhF7Z5FpKCRX+m5sRYocV/ImQrggP+DIZE
KYAUqAYxyGfd5TrnKzEyyomOsDhPePiZ/85GxsAmaCYBWony+VWUG3y42JeaOe8H
AGwfXksGz7+/pjgCjmrcjUID9+WWmLkahicywTAKq3zwxEwq8t6zx+S9BMK8NrEY
pGEDPIVsnjS4G8w6uS4T7DwnDtbzP5k5S+kCJmwfI/Uoxjvuud8edH5WikLRJ+eG
Pblrk4AKD+mnu9D77Gwnp8FWZsixz28GkQxZuNmhOwIihF6BkyZjwQWVbt5d1Wvo
WKSiKrAgo9IYVFE0b1NpZ8TA1WQOohs5c9/GptGLAPDno3qez6pGKKZ/NmXa0x07
+MoTP7kKTiilT69b6sAW56eqxO2h0BuuVdBUL0f/MQYXr/kmvch/2IckLH+mv0/G
EFM7ay7AhaxM7uX7cNETR8eG3UW1pJFsHTNuS3FCldnBF+k9xCJOgW8MKsgzR36A
mEf3MY8IgnV2uBuxdJ4Te2KjQ36wZwtZ/R0P6rZWZelWMDuwv8rB/OQwUB4NLObC
B8Mwxoux75qKd8Ia0vxWE370xLUWKEoB5+s22GLTA22Jsy6sfNztVuJus0QPG1uX
3Pl9omY8Lf+VRelYNEyrm7UyP5IlY2G46GIHu+5wDWGbwKcROLrSRncLjQD8V/NL
YfZYI61zgSH5DOA2gx2UVhLBBbBs1IGQtmKwdzWiVQxWCwiNeg7LBVoDNq4ZNfhT
OQdhLuMrgoJU375Zo2UZfgj9GLmymN+/NB5VM8pEONO0/FIed8cGAR2nPNa7Tf7S
rJIi9nmOFJD+WeOekpfR8tQ6B4SfomVOLzarIfM2opAhH5iX8OSNAx2BxLqsTalC
FJmJb8XsBC8bAxmqcEGwJY5WrhuPvWIeYex4QTcybsRw9h3/nEUN6XkM4YwrNrLg
GTAVXcWJXzXy6cFx2Qty6+9mUNqhA7xDklWFzVi0oCnERgBsQ0D8JHDnYiZYMiz8
EoIyuNH/ft/E22BTBkM4SZCAjFMx4FqT6RZmopQu8IdDP0TkYeqDeK+jReDP9VmM
9LALumqIgfy0T/e2+6LDEt1tFJlqwtEPbtwXlsSNxTnoQv4DYq3JOl1GCzcAirg/
f7AqdjOWUiIDLlmDdDdenQW2nNzZEU1JdVdRxA+v/Riu07xHa3GrJvadm7o01mUc
oEWaV14ZS645tBYA3cRSAtQyX9VpDPZqCwsFaJSui1v/96PXJRkh22rabVd09/oh
gOmA20swQbGZXqSazoe3RSQTaxMEAAUpo8NLbqcuTVsXbXCjUvB6WiaSasiWZ1Rx
ny2tLkR9OOeuNrItqXS0U0Keifc8xJqwXvZyqFB9yUc7wNW3uAJOUmTD0TUjLgDZ
8eyk0IJ3G/XG0BYbLyyxr2QzUAqIC5OctRwTI6Rh6p5zTNo1Bi4L4+2WYQ5gDGyt
p9Pii33dJIST8NStmQNdFlhPJYKkAV/We6MqDmPMZnm5knGmava748wtrIgP8DDn
oX5nWBhkzN4I50SW1onJ+OkA+tznInga0DxI/mDT5G/bsfCAlyL/SjGo6cnqibdX
LOl4xSFp2YEndvVF2508Lo6H4mALE7x3N+TEyI88LJZm/xWaT5XGKYFLuopld2Vq
hfYJrhFU0Vq3Zps64SM97Po24zg+31GQ7+csALoyt1YS1SP7LEdZH5KQK8wg/TIy
jssQhpHMn939A04NtIsd8w4UDUz9o1+O84dHTSo1cvFDFiSRvosK6LcrNpdILtoC
lsjJiGkLzwcBggULg8fvswaARw+jvvKnZkCwTLrOxxAEy/A4FFlEptsMc14vUqUM
k+oBu9gcVmg+8ooxYAWRpLfvSnO8lkRZRbf0qr+H0/HVuST0P/2WsleNXZC0zU7f
uEdtInSIpnZdjXVMwltBnlnYtBVe9+Jxs7VUcBe8hkroyNNIUdEXT/VIej7ARTnG
FBSCDisK0TK3MoAeyMZg7XE8uH7DIGp+WzzokhVJFZOBtX3nK/XjldC3Zu1SUoBn
W3DOqveBeBjFdV89rfCWVJlulAqzHKctyjkNrSkr6IrdU5nA8sQoxM3ovPHPqLyn
i2NB34rw+Ip8JGSxRUiYCZy7gqX6mmIyspv+zCewEJq670JasFtpG9iHRqVb3C0q
thVTDssNyoCc19f6Ee1Hyw8DV+dUt+e2vAki8+Jtxsz1fMd6ThZMkwAl9pUQ4iUu
vZTyPB8MGZjHewvRsxjePXV9j/znmtFvACjDqm+E7qfN+d4NNCxWfrtMbj/iq3XO
cdeJOp5fsjRLIrlqnwnKibjtdRKVWJx+VlVUx78JXQGcVzYcZjVKdDkLxaCBchLd
RZ4/QyU40IoRNUzvTxbwrLec5Xt+BktEJyng7O67nt9F1ZgdtdQKiG7qsjHwbTZW
VhgwQ3BrKjqgYXRDJU6vC2/IQfnO7NYZRm5JqXU+zA87OKNc1I3Y2oM7nGI4SbFP
R78iCeIDGYjtGkDHOj/poZ3wcpWrgiPv2eTMQe2MzqEX8kDDiINk+X0Jlffg/cP1
ei/uvlILVUcHDeWAoizEpXNLyxpu5Yiq9qhw/a12fUQ6aPFK43o32UjKZwqM46Rv
tTvSPUwOQwCjSwWxsWy+MTx6XMXNCLEM5uBObHiPV30A8WKopVKh54PF3+I6RTNS
mZICJyme+NTLhp8IZZro5OM61/N/lqkaVGeruDBsMu/d6WidF8b+b6wotmauvsqM
e3KZamhFu9tym9tXXKuTL7NQkSxWhL8LP8EFvUfFrwCWNJfOVGHy0yn6Btl4MJ8P
4+LpNBnmm/t/G3XRfGeXiD++YtgR4R389PcVcf9vWKF2WxQIe7E9mm3owKw+49Ym
MgylBNNCr/J+Pr/tGFKhbvB8Q5gJ+vQUFtfmkhDUz5Ckrp5X3nRWbDRsvPqkc70b
/g2XB8stxPxSEMOBI07nAHj1Rx3CAAAYBMSZzGqK0/HiIoARbdNV66PqYwOSW9xm
VfD+vschKXlQ8sAgeaiqlweiXIlKnV7MNByRkRlBfKjovIJayepptLewJ+y9yJmO
1OB61MvCDRB/R0d/3QaJfSjC+Vnu0m6ffCWPRdYZ4GDnNaPfMLRn4fyov+Da8RdW
MVsYOfDeP3t2iwQEAaKNBTXk4+bi33Ugg4m1aWVLLABXiRiFVuiPXNu+II+Ke90+
1cq6gGOU0wnd6ItslQlgjBFyA/D/wEue736+/PpPfWBCV5Y3Pn2HuyPcSyRwBRcs
/ZpIGHUs0nqR5aUpGYisux+9VMRAYS0Fctigy+NJ4rEaySvhmim30864mKmoumJx
e4xkT2nyU3m/yDDK6wdBuOZ1m2sgvSD08Vzww6/kuPyjgaMo/3ZTiHuha9ji7WTq
Cu0JXObHQLasiK3gLWpJjDtmQ1Y9nGE4BTkMNfOjDLp9T+9MTp0rEV6JMYxdGT5M
4ZFMC6CkmHF0zp7Jgz+AF4/smu0HsDp9GoKiPdoKl9PK0QqdP3Lvm/u67KYrO8hF
8uxmlt/KY1IHHQjJyh/ninA3r79SMCI8y7/V1AD9hXhFxoh5GbB6kgv5hbIjCrJX
VS1u5uIAC2MwoVuqrZi523IEuHOHb4edWZKWKOPEDz3jYyoaJw0jCZrxv/USgD3f
+/z+7AWwikexwjtQUiRsB6KRDMYq4Glb/oERBvjy1F4TH06af3l9D0aEHPuU8G46
bXED+1YpTp2D71SMU/u8YgelWVCX0obLJWBYgwas9A+/pOPCikmpuAsEFXENLcmu
7/ChMP2yTvTqM8e8D9NTD/ybDb74idC8R+jjDqCzWYi5tQx+oC3ZZg7O20b6GgUe
GOTD7ehMVVv3SiZbxrox+Xqee3HnSSo3rG5I3hPlv364DFaj2v7ctT70fCHn/0aM
lkaaQXI23fQLVMv3rNxev+z2Yooo+ype6YlXzNpS/6/szDO1fYOrdGY1bpdXGc9A
Jl60PmlJEE6lbhSmpfTqFp8NaPuf7ekc0hEOzP+JsJDpI0LLKS/Jlp+/ooEz19lT
+oJIImt82xNIDrLFz0se/TjKIYQ4qduipk5qa420Isl2aMBi9PsAob+oZVWANpaO
2FPLSt/Qq4RedTiCWPPBQIVhJqpIe9sLvb4cFpCrmrQBOLHglMhTdfid43sJb9eP
HW0aFGV2rAcDSI8Ndy8GU/KYPo/28fmk5NylOmM1u7USkUHhYPCYFAS1FBaL7kcG
nAkHj4S5xBysriEmF+d5VEkvDWUksn6VXgSv9RT/elXKTTs3EXdFN2ef2hV74PKX
oFym9/2vZPC07CAJoheloDccskzNXhRSGoZJAUybA9P87eA2gRiTtcO4pGmROs2O
Jk6YlCUZSMtHWsiqK64Cr5IjCW/ABXVpgspQtTmRhVkoQ5ZdeyEIZOuXRIbDKVvi
/XZ7lc4z0hh//wANOLZLlraoeqsEJcmvIO5DyW/P93IlBN+CqPtMy4Mt7FO63CoS
px0595WghkE2Gc3n6oUJTCF//u/tJMu83OK46YraH5tw1r2KWatTIL4R422ED7d9
r/rdJzjot+9quWAxtxSWX05FTbB2bmnQacDFGYD4Y5fZvUIbshygYLS4/4TJ5C1G
DnQ0qC6v4nW6uptOXgz5ycHN6FDTzTMYzg419SXhtO8vYdqrkDs48lVWFAHhzL65
FIj2v8jB8kkpt4cmReofU5/i2uxBZqzmvJ95v5aZCuj0UMe69+D4B+rIPLO31jvJ
/Kf6x4dxz9TIAs3D+s7jLEV4PNT2878Otqmc0dczIK3QvVm/QqnRK2mAP+pUuNgD
Bfx1su06v/pQ9P0SXWE7GyxDDPA2Y7BVItIyMStcOp/LmnrtGwej2IOb/Fi7TN/P
P65X4uMWqsMhkI8JVvFbhqJfxZaw+fNdsoUF4oeATd6U7awI1NSDhfilDZgnMhZC
QnhFD8wbBE7g/m88ptq5RjCeROVQVr05oYIaq+4ZCWqbcr9Ukkx949tMnaxLPlum
FFHmingjrxLKM7OSWWElVyH0Wm7ivq+eyXjj/MH/Ebogs+cnjYG3zDtJjnYPuWoF
LMpZ19zFSA1WYSBTNF21k8voGROXTs5IpsGBkzJokAryvC+EVst4MLZTJN4JOSSo
aQMZple3T7BqdVItzDCy5ru222n3afhJeOUoW7J5pbmKMZL15yU4+WUViSfHfns4
1ppVMsK+X4ChA2w81Znbg65FipXFTNxW/6h8HE6DVQ/2114VW7t3g/vrgN8qwfyc
ZMDzhLrC0Ibm17cTsaMArCfC9A7Vxg4qPz+PHDVoRN2OgUpud4dN8ndvGNQckm5/
EymdOuN9ANI0UejBClqzF+Si2yifAiWTnzyVVkYVtSsopzFCfWBU+8cM3KgxK2CL
FRucbncP3RUKLYMnn/EMUkCqjwyhh/9xCjvWhLTy+dFjWBylI4IU6dJFDKu+Yq+c
6dEVRh4hhO7z5hkvOzxpUE4qCKw1MntlEdE0ZLJN+88vOQlB8pIkb1hJrIPSNOgk
k0c0+mB7xqh6GK9C2BI10d4VS42PF8Ok2IDeaDSPkGYCQabyU3ngU+wOLvHyvmy5
LEDP0j88n0AaY1OJgFfmOQyvfBANCVBC5HyA+1PABccN6FFKEFX8gL4GrKVHwHm5
bPKDUaHaIm8MRsDKyAQpJPZXhM/M4Bw0WzRbukJ3DJ5T60vVskctNQRm3rvLeHbi
mZKSAF8xg9btoyvbUVs5SiLBVfcPRNiDE/Z92owu1B4wJosNMPNB3eRFnnMafCR3
bOvApRe5cA66L3kkI84RBtD0tpWKYr4VA2meaoBsF0uIlaaP8F4FJKtWBWXJfpfW
DDH7K9CmtuzbHVrcCE/NCpylBk59Jj+3sdpKMccn3XjHZfXXnHl9ubI18vSbrPKJ
SHkPmWHSof6H1KI9bz9cy9iu7/dxGF9V9yA2cjAsKO98Bxk/q92vUgWWa8B87fw7
9XBMpj1Nkglcr2BZI8RAlKm6pUepz0cExJxZbyI0oi5LFNkymBHDzAD5cPqlMB+3
fmBrwFl55tFxW4WLqUDYSNOumdhi6pM4UGNEmRqcWrVSwvAVi/vtKHVp3tU3zO6x
JMFIaS1tcaDqV3s0wjTCxOpJpw9t3yBUCZsCo13Ap4RqEfaMU7yMvXQWIjINaqwy
UNMorHD4RQTf88MczhzpPMDMWKMNRojDR/ecVSDA55/aoLzPeK6Dh0e+1uGJ2chF
TM3Z+kMMOH/2bD1UmTuc+9JG/3g5LMgBU1W17/FzVGg0SQa0yYYwEjhiyk2QsQex
RgCh53FyzwK2uZR0eyu8NSmlOOxd7WvJEuzHZ2cb8VJlh+ixsVolOwND6jmp8kdh
rLjbpouJLW8ZuNIOcgYdWzA1oqHFTxX0906L0hjqqYzSjbzhBeaBrHkzzirbYnsu
ewFeypXED5wejLNjQiH9bvn9PMZWMbdv2lRrrinrYHCdFIZrcGIkjuOnPVXBO3Ha
udImgfo60F/EbrbJznPvYs3H9uqpthakmcrlEFDaP5qSAr5ODn0DrqBcCkicg1B3
LNI8De7nihgybfNEOHjVKENSVMk/k8PpDclifwXerZmtSgc0ZXAq1zTjSqGp47pJ
5oZ+CagkyyhqLJp0IN7hv9EpCF3kVeRFSle4rVax2Vrlr+IbjzQoq09pUwO9fU69
VQwhtuPCduSQ+YynGLBgA4EjUu2mGUk6qf4L18kzIMHPerdE4vumWyQMBc1u+QrA
+F81sXuwYgdJbQHy6gYzwpochT+FD/Z2373iDa5LBy3ZEvYSXbXm7X17sow3+3MC
83zsKheuc0aJdmu/vKNohSsDaAWFk0zu3LsrI5cDagxuuVc8GDpBj9XxyvH1ki7z
m8j2GWy6LpL/B3gk5iDez10InCjo3WK36EJyMXXYQIMvJj3fDL1aMI5ay9rgJHOL
WF2HNyRxEMseYxR6y0I9CI91wpK6YL0zvKlQzmQtC1uqUa6ZUtMUeTTDKJycpigc
EJYUJSw72hCmR11S36dnfSAMwPBfTmcdiRxzKmWXtrcsr9nM7GwZYF7dcAP/oVLX
0lsOi9h+70p6sxILhZYrm0vr19yHokIWSimaQYNfigmaLWC+YJwXea/1fsantj8c
H77vuTmArcnVs0iilGoE+QcIJcMGZeWWsiMtlIv3rKlaL33KMgYtb7C3iBJNPSXW
5/cCDQeRPvUmvJ37zpYI8zTfSp+Q1y5+0LG/vgM8sCeku3VD/+rxQ5NgWcmpV/l6
uzFrMh2B73yvOj9yXGAHV4ANYs8rW9+TUi7HrHrMS4mFPzxMswzboHm/BnMxq+sN
rlrp240NNhmpasejF53+72kbE9xoC13cn6wJDV6OQE1WnXaHIsqOHIcuj/NwZ9TU
H847DG/QMaZdB1IeFNwYAzEc8PlhRU27JDJ6dhv/qnotdTGD5tXxT59z15Vaox/R
jMQskDzsqUPZW+96aH4b+1oGdXVwFZH73RSI2ccHn9Y6zYW5SCPkpa+m6yY/9LjC
UkXZYmX8h1jVkqITIC7mumpn7zKWqFmmebP6huJp29kXOYDTU2g3Ur+0urqsnjTu
r2ORXFHL7yVLm6rGtwMHTs1P8cAHVDJjnyHmDxx/Iyroc/3JcGpFSjjTu6IQWWJ7
d6tYk4XMu1IHkGT+pnKsQ3hSt+aLMkpLw9107AJCUWxeBzUkGWmq28kOMtHSRQm3
IYufcxzWq4RAPMmTN56jzkAxjs2AlTUIwqRDOvrXEm3zA+Q8ZSCI6Lo+FZvadBgQ
ek463xCQrqpEt9pxgKvyxVTcmhoeGXE8WOUWvGieMKYHiyBjzgmYaeyIF5bRiDat
c4vxMikBoOzgAcfgGN2ew8RSoq4CLszrZOGROUeR0QR/zW1nNdUXP6VLJINx6Zpr
niEV7xbi/atCl5BJjbxNqodcnmQfQA/VypxTq9/t2U0YVOFakn4F/pEf5UWJhD/9
FvkC/WT3isDBJENE0F/ia9JCEd7tAoZzpdwmcphhUCB/xK1eCuQwSZPJblqolEx3
c5B5xn1wwUrcL3RNHBjtFSF+BFhDcad9KSQiAbTqJOMIJwdEWybxhle90Y5neKC8
2wT8qYdbpFAwa6YVwSS118P/BM9oLuNvIGE4QkkpmvPoZg81BUO49FHRj8K6z5Ei
bO7YaSeNOm4LUtS7lYE97yMF2axBHEkDZaMj2VOq8vmzfpN4sKiMICQL+0ppfhZZ
gDLVHcgjcPUo6u3NLyPXhWs/OubjCn/8r7Dr8psqI9+yzRxPRh3dqV4rjmceGDJE
cI87x6OjZemBK7z6F+KancbWHOfD1tKmKEV9PaqhAk0vFoH6ylOM3LJodIZRNVn+
t5mjiJxle1n4za4NRw6tLZ6r7YoLaBSy6SENNbAVvXO2VavLtsbbJOXZ8BrieAPf
9BYjqoxLgVyZI+xC7WG/TqAKTVEQ6o49P75EQFm5xTJgoKTGrWiHlBqvT99m5b1b
BVeVUHajUdIx4uFbxF14iR+CojEAHJWXyQ2So83q8AECEl6ErGwzK5NhFVquZVUl
etMXCNmkDdN0RNj3Y+84JZ6MDAI+kspdO/kbxFl6WJfUGFggLuWntnNcv9yQ9LL2
hq60+uh7jfWSm8m5D5bh/kPb1gFtGprrbSGM9viSBGc4RVMkv/Cae45g51a8nOpV
iflehx3zUIaVl3dqF5nQdLA0m4FsDc53lI3FZMPPL2HkA6kDGXNBEatGKhcaXE6d
A5w7Crcw4hI3rFtVH6HsP9wzZJ3EtL6StwIzo8VSnyoCIIH4mD+Ag+hH7k2FTRn/

//pragma protect end_data_block
//pragma protect digest_block
0NAANkqwtFQiMoCSvBI6m4N6j4Q=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Z+8rHxTCyM0RePmgnoGE78eK55nHGOtI4DbNvUHzovFsoXzzDXEeiyHiL9bPOnGp
TaYnPVJd5xJ+ZwB8YdlTgJeWo8NMHstrurHp4uoV+Fc9ET3qN26S/+APK5oUkQct
8beiJdyBvlSOziAz1ONq4ATZPNxHVb8MenQMYld+grlqH8QnKqldAg==
//pragma protect end_key_block
//pragma protect digest_block
l6DsYac/nctKAg4W+0cjKFNO6Ls=
//pragma protect end_digest_block
//pragma protect data_block
x1qhrkVp76TqelldrkJ+AKRdxCejVGd/Mok7n2srLRGVYTMQN3A0Kvo+G4QvYCNK
i/dBqHb5R3ABo4VQH1bLC7INBsD+7hegP6t7p95FprcPPEuOqzCOWcFh+STSvitd
hRsThGCxoI45kFBUAvVA1UK1BZC998KDjlUK4cKPkMBDtRuIJDXzapi13nMne9va
TQ80P1pbIi6zTpX5PjAT8zHNM9Q1z01YVKdP3/5ZYTYoxoW4OjMBhT9IsroSmk0C
cHdsQyrrUso7Xk47e/zSl1FZ3cG+EFsixa6aoAA7iMZu1aqa25XfE2ML3+cvD8M3
PyP7IyZynzptEqKhCPwSLCtt7CHXSJKZuroBIX3w2v+emOiu39RMxrjss7IqGn04
Cv+WKY+xLeXHH6lW2NF5djFeTzAoM7YigHyuvY/VWBY0DhnZKPY9NJI65efelfBq
bkH/xlrN2Bi0sp+69CDIr3Vmh2nUlSMJ/Agurh1ZjqHh8uUyqJYNo9+UGGGIsdwi
zd3QeAofacOQjm/Gt852gXMCj2zOMqMRKC67i2J9o4uplLht22qT7207/S0CJLyY
0F7+1/JGqMB6c0safxCdkWlxV83JdACpdWo7aDLwEv2n9x3Dq8eEOTZ3HZ0J7CvR
yuuGNQNEaJuDAazNliEjdCoXOztl9k3GlBvhxQbz/hwual9q9TlXT5ETuk1JJ8Y7
E6b8tVUy6T4LU5BzbIFPtRT/cf76HIlhBI60P5jQID7afx1DFk6DYL6IW11cwjxZ
g+R9oHT4Az8yzBKZmN+L/pXTSXEDxFjwQEdUDjvJ7d+yRESnVIf0ONOJ+LLLO1pg
Co+QHaQomH4GF+RCpstHUJqTWGa95D8rQybi+p5bReZXvUC+OpcP/kkqV9sL/5jY
zU+0KoIanZyng067qNuWDsySN9mas1IxEB+WkHzRnCe+bpK27Rvi1cuSKs2F3K+E
SRvepwfme4cjXMgvqWi6MFloJNLC7ZgBRCzHZ/VMx9iF3qctG9hZT+KU9qkENzEY
eG9VAR3miekqsS0Hjtb3+pg5h8onirgL1lwK17qXaa7NXPhJtX9v7SJZ9M9+lMlZ
aiJbm9sgtrLak5GFK/Y7m3CUOViRfh40HZMU1jkUK7OAqOISi7O8IP2JpFuFw4fS
rdGD24ZS1NNokTY9AKtAKUYNRnBZpW0zP8kNrfFd7MkDadQj6siScAJ3UEQcxMGQ
XFmOULQrmoXhgKjBruq/sLQi0MQ4nh6Z2wWK6SsSanlc9d5Cck8Vh3qA13puMr8w
T0AwBtzSAsvv8lTMZgcjtM4cubJG8X/kMEYzDyUa8oIJSdJrKTHJwi+D8ESMaK/H
P2FI0yc2MXZjPiLx7wpX2ibT7klteOy//Ceqgls52XoDXW9aGqncK29FK/tHjta5
BXVJdYvtQRfY5d5Da0W2sQDiGAiiSXq65dokeR643WIczb0oTXyJnLLA4v553XyP
YyhJnk7AsSj06W9aLut85oKN+mGEX+1JzEd1LwaClWPQ5K20QYEwuXcTpfVvCBqc
G4SfeTeWLx0OC2d0/exORanO7WNxzpVCcbaxdQS4RBAgEBBhI/CEf6UPvpIoSu7G
0rseSaOaqk+uuwsAJIrpCSymZc0xjmyCIpcnfnrIx7UV75BOYlVOpSkSG08/3aE1
7DS7GKuNQFQ+9M/bgHgHYD1R2J8v0oGdYd8VF0AMt04=
//pragma protect end_data_block
//pragma protect digest_block
A1nikVaUwBikac0NSwO5zGjjZPM=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Tqplb8JzT6Ts5FHXxXWF/SAhzZlFa3QPJPkzR5Bc9wjj0kuQ/z3Bz6rtTvzcjxz1
WE6JkwlQ6E2X70P/uuT0gjrLA0oO3jBs8Vj6brVslMWxx8CtqtN1PLseiGeqeBgW
ymCkGzzk+XzunFupVfXVKEq5RpGBA/tjt0Uo5En1hpO1YEwD+IawJw==
//pragma protect end_key_block
//pragma protect digest_block
GoCDrK1JmlHiUQ2xqvhWpxX2WGE=
//pragma protect end_digest_block
//pragma protect data_block
uemJRUuPdlbbEjr0xQpe+6VP2OnouHZgjQV3DHv9yxgug37luCN+F9zdq39j2PqC
s6cQI10CG3kBd+jCl7CMZKdzVCOJU0f9U1Z3LxHeltfY/cccHjZKz0TwwsIFChC6
/Mw4KCW8N8yYc+U+wgJWk7uMtkTNA6kieqsFwIz3tBAac5ROfbCwbSFmbTMwPMYU
GOh7l728vUvvARbK7syxHV6Pkocn/ZrP+OLIxKX4F91FjtQMLGvINNyIOQWRqC1/
TCgdxL+7H+Ri9L3Vin/w6vPYzsrKmA3pTFkgWk8t0vxtvFn3sHEOduIKhO9sHQZA
+BHECR5qyRw1IBaFerolh+x30hHOCDh+3+5ntESPlTQbSV/ZYemFQRtrJOyHmZ2t
GxQ4u4YleLS+1cdVvtM3+TRyKbvkt+rRqz5IBIze1uufAat4U5ZjjXcPEjpU2v/z
2Avb0y/hWFNyEcp4ykU3zIs/P6jYnTZzlTdGxkexfbwD5LMSGv/64J+z2+m3aQdL
hsCh+L6/mFqiqgJbeF37hWaRD/nzsoaiCyIV8UhWoyUM5NDQHQxI+TVRt3Al3dqs
Y2U1oiIzSHXMKQlPoUnkbhjfzOp8u+c8LgEFEDUkiGKQxJALXYW77lzytGVnwSuI
r8DQuafYDajpc6IIRNvtbe0igKhPT80dLYX2Rdm9VQpXkk5QMcpCkYBww9uCxcXA
xW9adFZSH+Ab+QHdLuG/YM4c3of7TyTW9wMJD3PHtQ2BdbEG/yqkO3BsW7pV3skW
W9D5q9nHhVgnCy/bp5FasaKkp228GO7MWSxrwBWjkPFfmJ5aanD2ZzfCjD/qsOaN
YqfT//K+Do8e4hdHZVwOn0AWKIwUogKPvDzLOmmEKY7kzF9H16cU+WNr3r3xFDzk
+phmXYyqHc3PsnOjEJ3VA0x8NvsWN1zjcZOabL66NOniTv7Sl+7sZMrx3/qiQLvI
dRCbqvVN3GYWEdhEL/33+yeoHK5s8VBWmVEwgEcyauxLmK+E9wozn8Boa74qAVvv
mXvgJAXmnX0CWnqJkxsZexN201WSb9Cn1hXoTf1JSunTeA+5Kl2DLR6QuUs57LGJ
K0vnenoUpcbj4pPKFn3Lk1QAyWEB87ERFLZy/ngUK9xR/WGPLbXLYkR28y/Y+zBL
0wQdqa8NnFUH81+hnDdrVGJBEMpi+Sfauk9n6u/Ar3ImjrQZgUQhVjTB2+31i9fj
q8u4jTi8XBh9oFdXGcyJ289sPVGVkuN/3hFXhIeBYGQumEp8O8IKt/zQSqmBe33B
ZGoRBTXH/FTRb19oQ0VG94gfsRySmEzkNAV6H0EeKPRiw728FZupBWNIkF8ThxF5
E6Kx874u278gpAbmU17POar8qGhGjHm0wuWkp64XI66dfKyHgUW5YMaN93Y3zP4u
u4nGLUHsWp0IOAnyOuVwfEcYMZbxGUztyGjH7w8AkLrokHTijRIv1lFykwb9k7bg
GxemfR+3PD7iid+qJUYs0/hGBgqsgKGAvMVmhkBFDeZTvsHBk586xtlSjp0GZl5O
Xb66AJ1bm1CAgfNzRd9wAIpw2nEIINK+OU38MgKQdPdPzaRRGHW6lop3SZS8pQBo
oSVqrjvOhYi6QXT90BFmDT3kh26ZSqTExkaLRCE18ZtSUqGrxn7wG+HqAwRP37iQ
uHpsU9t1obHFzjx+L0QvwyERigeZaMhSQ6E4IdwWKgvZBv6WpFC5z7Wj0PiR6MWV
lZ7ni+i4SbLUgncaE6o7PP1QidSLw4BK2LzxadjftaX517G18EHvyI9uJRNlmoNk
IMpYrlyo5mE2+eTPlRfJcG9TsIcY8P38KSaS+ZfCvBHzDMiz9mT48qeeYtB0pP/S
abnx322rlw0XtVMUOwwDkYUXXTP0KIAJH8mT2CI7EasWXB2yyReGBtW5fjDbYvG+
5OQFiEMSquwnlE3v8uMxgXujhYcfRRCza1LviD1GFY7p9KhlflAiwKnBXO9LEqmh
TkaMK7vjMAjqNkEFy71C/qJwdwLc2WLbC7JgBXikfV+fnJgJyl1UOV9KkhZUkQD+
xAWpPqQdkZYfLvI49wEoB0T1IqnXdOiZOPO/sYcUxzGZVd/loEQJMEx6jUaptxsk
3jmQD1TygqQb/SonDtU8/nP8UoU0AD4eLGNoxFe2BiIOLA05FmzQVWcF7y3OhG5z
3L/wAgBiBf5Cu7WK3840+xcJn9Ym5P8jb+uGR0ddPyihnEO4wcvyiw8kRECiA5Kv
uiugjDawIJtfHHhtXzaffYLYwMbMBZuIIgCYA1bZggAVitg8zegtSJMRzk6YodyG
JYibB5noQhD0h8nsqctA5BaSIHe1/Y2R0QXigG9evh+FEIkF0LTVaqkCU+5hKiuJ
kQLe3eq+5vjTgSmPrNc7JqUrNT1CWG/yqVPKqLoOlUo5AnT4P8f0YB6kuxmsfTN2
KqeoMPWosM88yS6h1DNfDLGD2pVr3R3lXaLUNQ6NOtDb88Kdb3tgHqYtjwQRJgwd
0xIuXvIrEmpO7GxwZwGXHYEmWsrBtTG7ZX++0MgyUdPJE+BYomEq0I/vkDUpHJp9
9ttKyb60Mn5Gu2jDbJTkxNnqKT1zrzBM+Tk8mH4DAUvF5pCYqs1M/aSmI2hGZRzp
mRMPZRMhWlNA31R3aCYLpJXPdYEnX9u4L7PH4QS6RbVSDiLSeHGp8ZhVjpaYwdpU
+LLhmQegHRhvmG1x8IkP6HOlZO8L/TA0zwojqoSnJTeKJwKegbxPlrlOOkvzRG6d
y7nPgADUsNHqOQh5iPkZMZqKsXAbrJvQAkQOYcJRWdryQ0m1oje8dZLsk5vQ5HeP
6XiUD0PKZyg85IRhpVqS2ajxUaLORohBuaGwN2sSGtaitdr666NAesFxh6hHsNIt
NdDj1Wx7xgYodHpPhKxtNcfAG9bVaT8q3RxtVaT05DtaoM2GIQQvMdboLF+TlBVP
e9UfoZqAbbI+dZ/4hYAJhoavc6niLnsLX9AD7Kn3wASlXo0CCNHUN4UTv3dMZUsH
t4oHFhecQPEG0oHyECgKTgUCuGgfR+NBHafUZZVjJv3kOz+X0wYTO/cdQsUqYDMP
MCs7hHHo4eYAKMsVjkvgefHKeoulq0FOa8RVobt17j8n2SuctTv7MxUmQNrUeOtS
mcHv5qOc65L8Zzcsa9Vwy00Kqk3QA/yMTTGZO1rAtbeyNl5IiQ6t1oeXUIau3sqh
CCmELx9T2H4Gxm8lnMqKCV1HRHZHIneX8/ZfNnOTGdPvfk8rzgC0Rm3gxj4p//Sc
MiAfrgWz2K0QiYDFq2xJmJAJu2gHvElHaCXAL59WCkeqi/JqloZF8KwtnROfL1GP
hdMXevy56Rf4uTQ0j7U27SdEIa2iyvRl0h9FrRQxV8cu6E5OQJSbZHo3gTbuxL3c
7m5ZKo2MsW3qjYCylBs2foAPMQCz+8FfySqRaTOE0TkfnvzsqWRfXpebu28PZC/0
HZAU+aAxULf+/j52K2jCEOovJ7uSwFE4Rw08KxaLjP0OqHYs0Xhdzn2BzfjQvMe2
BwVI8MrCtCnLZpJ6gkzUo2wPhfz+s6oRt51br07JBknwrTv07NVIOo+qv3eLVgbu
9rF2ehW10NGmtVmk4GtiGP/YMd7OJqZ+uAcc4YKVB7lIaVYrtHOfa4nOutnPBbiN
ggofWUrxehieIcC8amJSJTHJ4oToT92vnD9eqcTyoFAf3p7rOeFlcgNhcfjPuKKw
/gL+SOqwz//XUEWJ1JGaImeslxWqzcNLY+Vrk35aYwqhJnBpGuviSn6Re8kq/0Yw
Xf2md2rnOpjaSYc++2Rbix2o2jtSfRJQ5oV1d+7e81IcCl7KkG3Oq1JAOP5GJM+0
XCpJzOFus41zuDrsc2GiQtCGzhmIz0hXv7l6j7Yo+9j8c9hvsnJ3pCoMg2TGvX95
BtiM/CvDNPfy9P+ALU+mWLYNkN20RMTCTZu0GUWn+oP67pNKrRXC/zOVAYrgvVIN
ZNA0BpPh6wl5RXVreVvqDg9w+9S4HWHvJUgr0/zPztfQWS6NmUvI0VjMMK86Z346
gVCY4KfUO3jPhcJ3pW8AjaSh+ZeFJOwursUJ9rAUk/onSRN6Pi0NRP1hJfObhKZZ
UW7oy12CkFOivSaVqVCRSoUNI8GTNtueYih4szv+GLWu1E1RPYho1F3prXwdrPCi
QCxXHdLVIQPjpWBmNTXjj0WcZ/PmnNxeTXGnYx3HXgQG2WCuyII8pfLK7ncqNJeK
h4iFpLFlRo9ZNvSnKPds2iicQgvyjMRpeUmuAQFL0Ux2AAec0RTBg8BLGhc1pEpC
MnqcCFLQbdgMO39js1Gw95JilSdkmvG2OLrx8TLzkRgT7qlsgh/1hdlK9s+I9hJD
cj3JPNiOBtZb7GXTnsHoFr8eG+4PEmnj1+3CCiCczlwxRbwMBzdTXrvKwoiXZ26Y
hK/Kc6FJcruFVxhoKuYXIWublCd6fIlLjR++osDQ7c8UcrHL7hmSnXkwpA+Y3iAd
BdbNg5OitXE5rtYbUOJ/DAuiZq5cLtziqD/L+mW+xUMz+z1p0kow7Zyd5hTGv1kL
HBbyRRratUCkW8u0Fu3yaBlz0VhJnCXA6Y9ah60ARXxKPBzNjpDsPzxeQVhGY+oV
MPudbRNLJZucxYkKaegHxUOnQRNCEn9M9RPGWeykMJTWtlDXhifzqt4DJ3zFEx9r
fsZyvQA0G1VSxXzVkwHUyxjsEGJ6B5gfGfb+c7qas30+iT+aAvfBBI/J/csqb2rB
Lrsk7WBwKVtQIb52FA1bCUNmpt51bfXe//OMhkm5JBsxogpxT9EVn8K4uoWN4yTL
Jd/d/UXjsVSGUcHc6F60lWh9idzsEzuIE+lGdnDe1ouDU9O7wkFfEF47p24yWSBG
H6BaDgvxdeJ0A+7DsZZzMZoLj0D5zO8xyM3QoZ3NQKumpCtRom3WDbKDO5bMkyWH
otnfD7ckj0vSJw7inuasor3z/IHlZyYWEXgZl4EpaCCiQXHHNan3vN2N8hA2Im0J
eIcG2MwKURH4JWgQWSdQ2LByu+5Yap2a3pa8tQ7g9oylJUgfknwNC7wZglwwsFcm
hp/3f4shUO+ESKJ43ME4iKWhKXHqWiB10pAKU16vBOybHorY5ILGVOBjjrCf3PaO
ba4gidA8icvb7oqsVS80mJJRDeQ/V/UKYuXqTzLdV5qO9OMat1hEY4Ooume8cJ32
CrmOzBGjmP9EF9C9Nj1wXNqMykHUag8FjxvNaaAFulEFRgJo1KWEEuW1CO8cbzsq
EXfIBog6OA2GWqpoTZP2tuQigFh8keldvdt7FcWFzFL4yViTUgUrzDFuAyj027MG
aCRIFUMpwchuC0z3PtUAp0rygAhClFJAHeDC4pDy2ywh/IfNSvSa2Te5EcGNYckq
LUqlOhT2QGU6mvTd3V0INALY7cINfMGjBn/pWgsv7pOiei5OB9DeSE9uQWts7FoZ
JSJUZnfDn9yxektFNUqwrNvT3fSz4JH+yhyNUPGdXlIFHWJy0F8a90z8VHq07Hpo
cOTDrTE/dY/8DVEHtcpMxG5pz1yEIbHe0XFnBA1XothSPJ4Wm8ITaM4NVTMsnqHX
ypPmHdgIUR5u+AbTSc5Z8RfQjt0l5fqzqecbbeTlnFFIFU0N8Aq/AEHakD3E2Ejr
sSQLoyZ/Rozz1fKN6PRukG616N2vkpr4B6FFSWIfdHiy2On9gFz/XO+87n/yYPiP
1qux8PnGHZRADKbyIxIV+WnT/3ZSSVeBZ1s8EZ2Dr+oEERsUOyE9jLYeT4bDpNgI
Zt9H3fKeCqawFZXKB5w5QTeHvP7aYTN9UdmvVtCL0zAZBZRTrqxsBoRUh6KaFLBl
WIy5pCT2604lqgYMGSlHysOcWCk0e5Qe5nF80kKY6a3Xe9JgBMx/t35uFh9LC/d4
e6cpYohJCE0akweQSp7CUb3AzvkLrRssifA4U/KJJ5GZCLJViyOHZddqfjqDZPmy
GEYDScsKPNcUllGiz6/iY5aq1FSasaHJffjP4wizGhH6P7TLlP/uaR+T/v5ma0tv
+T4/mrv8OtaVvU3C1wtQlYvimNLkfg5eyVIBxNZKD/wwQIvHNpFi2e2j7vF8zhsL
02/7zLBKBft1ZFBEmtBcfm4x9Gr3dwtMmNmV4oWCKZPictsw/HD16ciTYlmQ2o+8
qdpExiGKUzwQWWSw5YKIyC+n+krWaH3L4AncTynmD/ZTQL7cLUieR72F/hcWE2On
XnQY8gxg29510ZWuD55KDrx+vea+TKo8eitgsFlY1rk4QGTeqdLg7gsCgqRN1Mq+
b0tqbpxgwrARJGrS2CXmOyk3wchtZeB9GZLR5tZI+f+j4PVBbiiWnSxpmvbI6kYu
4sKjGogkJBQ/TMwZXBHmZIxn4lryp7gV75M64xt++4+gJoKdzgqFQ6BPYncnsI7k
rrbr4J2zeYwJjwM9XqJ6WKJkhOXiejf8YIA198zw+cLDq6g5er1hJi03nBfjWsHn
iZ+iXVlnpIhNcbRDLR/YJClOxfh/rhSi0PKCGMisIWL47ZVOolXVrAjze0glZcAd
La3XaJ6F8ChhGt1Jsxe1Acas6eRN8CR6fIoQlvfkWbSlCj2oGt5aUaCDfj+gPLtZ
rzr/TSrfuoCqFEhUMW2smbjreUJl/f1ux1PiU64LxgK2nmQgRlAvyUKY1NbtOpPn
6CUqFkJcL8FAjIM1Hi6y4CX2ft0w+V859bX+jZaxBHMqS/63kbORmS1+QZbjEAjp
Lr7p3jdx0ciBch9FEvGUu95o3n3xKILtUsPpGR/9x/XDtK9lUS3HVWTRlXv6S08e
QmUKGaeWS4umMMrOMrq5BDgYeWmeYox9wEmHCZVUOiL72dossRNwY+OGW9Xn4XXd
0nMdNQHweDlxOWEik49ddMDT33AR5rxW0FxXfxCqZkVKyHEM8fPcE9c01EFjMFWn
B9B48lzBfhY245zAZW6NJ3j+zjEsv6edeinznZ3BZudwczY6FO/DMwRXOadekIO9
2nw7+CFahMN+8eZ5Yuz7Er4vZ2dpD6R6F7G0O2tz76Qv9O0Wc4M+9ryIv8HGUh6k
8KoRgjDPhuRg382+rL9/hvbt6mlWYbNPpeIaFNQg2bKG/4b0ImMtP84fKyrp3X0V
ELdwqqS4rDL83LPbmIqlBWfoCf3un0GzMNnByAmSXda6q6fNLv2tJXvL0piQ00qF
FfdkA/gCJ80FHrwPHhNVowLPYcKmSfWk70nYiHqxzNXI5v6MdiiHFlb5CSsxwxgj
Qrk3zgSxr1R783JGYkPcoabhTwSUXVp0qS8M10nqVdYtT1VNDM7WKWYI0FbLBW0U
0/QwgXji3iaJaU0Blm6v/UGp4G5+NoVNC5yZ8MLxmnilb62mVPTB5+Yo7tmVs2UL
LNyvM9xAlviUB0WWRiENgFrp7YaHDQd/8KgqW+hc71t6QszRWJNsEApeUa8/aY+G
+cpDGZ5NkRgOwhFHoWaZhNhfGOpRuqMFidJHQC0U7sOXaaOiNwTIxtr9k9ikABzJ
d1LhEqRlG/HZcf/kdMusHK0HGY06SOfiLyiItE/d7gxbz2vppZQ0cwRGyY1rvME6
7xoLqilze3DlqGJ8USdahMrptz9uRkg4uPFfGD3pVHzJbCNfGBjlazbhuGYZ5DF5
267PmjTCyD9EPvebFrL2uqnOD60L6Fcf3b/p+ukC/L83bEAoI+RUpWTFOw/N4HAg
rhxs3nFRzFKdIc1nh6nk9kTEwCeSUdUDHoxbugtqcAWSNcjEJYs/ivJIBZ9ndg/r
qZTSEbSJwY9B2qc6IRrSVg33WKyAeQkIrX1L8HUPP0O07Hn6Iqu/efaeD8sV0OeY
TKf74jhL6o7kpo3DrIzW83Uj/na9cLtEsJELbijFZsT87ICqWRo/yVqXYaK/mI1B
oa4WJOp9ovJWCT50QPy4j0tW7tXF+zNcekXf21tdGun68j2YpuGjmaRJ7dS9l/6r
5rqCoBwjGvJGNPFgUqi6kHqKj4LI+zuXo6OuVgdF2z22FXZ9FwTtc+V4irSfmvAm
T/3gi2/e5zhxqVrqZgjfsJ3SoUvX3bTWHnb6mFp9x9RTQwIpUMP7c3qxQHug7AXv
VUTeYPajU2eOw2Jbge2tqZm9sppPP5U9NOErVRFwnjQRqA6FgUr+/HiRfl8CFG5I
zRaHVWUpTxRn41QCJZVP+u9XswyAxV75EvGfkNRkQQvT4LjOzbBRoKRYF2Lwtowz
TwXzeaUWZaEU1c99qZzy6q7Z9MKXtJbGFSvDOwZidAlC0heR9pyZgoDAHKEwroB7
fw4dGq8yMKwahS2OhBrNZc5LuRnU7sqmEhOfkbKeFIyXoX+hYzLfRWI3Cwy6bqRG
NSybo40xs200YiNPcIgALYLbhiL+cM/Ccs9Po58m6A1C+4xfKA/TlJZZSLtWZqpb
u3o2iD1cnn9NzEM+xSIJ/KnR1/hjVNCED6jhxKRIpNmN572aGlnGK8xc1DoHqoux
9DAJFX0cdTfVpnR1h1lffGoyZApn1kn74wSt2rjDEXuTznSsyx/tFAKCnKs2TD86
9Xa8wHvwXaWR70Tf2Ms3kXC8l+5Z409Lv7kdYq7elzQYuJbbjqA6oJ8X2cSDHnvR
w6x/R/pMnDzwkyuagZ5dAzOcENPxvfCHQP/8a/oQ17Sgti0MuH1z8Os+wUN1WT7a
8gyzm8aM2K/CiabgDuECe9l/pw+yKyWokxrJJkOyFsGB9Oermt4NtwDwEyJMktQZ
EQb67Z6zbPwwyPhjKhB950nKb94tZc2Oe62sgR9GXuJm3PIGA2qpw8fSGAnUGEx6
Y/8k3jHoRigrpMttnid0JL29yk6mJxwRnCr1VSH+uf1zVcSF2AlP83W+wnTrheDA
OL+j2kYg6LTf2Uo2Vjnx47FPUZPQoJ2Id0Cwx+Wne6BCO1C5Hkh6P8OJAZr8ks5N
Ky3mDoKXex1SqfNc++YG+DXMZ7LZ1HwvaMX6G5Py77m0LwZuSEMFrwnWV43WCopf
gxwnSZX92CvF7wXO5zwedfZjSHCgCQ2L9NZxqsytW65ISFLv6vjMOFsr1347597v
MqI32MU+fvbe+5CDCULWx4QBDf0thXKTHiNevH4t9WoXfMpiRVUpRMADL9kRSkMk
TUFrhdLgZkhN6qS/DfPEGPWENIsxRQBYvKouZFxK/9uIqkDf3Qx3iroVKCtPkFpf
xdpuzrRDUceXjR6n+QEQKMyLzziNlDOwTn9uO2T//MDf35Os1Byl2UwjwVotIaNS
6SZQFZ8pa/f+NqrHpKlppecyjcahF/m2AHiGHS4cPfEThrNWKd/vWQM2FsuTiAeQ
QQzheb4IGhL2NZPBm9vmxWoe+SemdcbwG7tqCylCB6hQqMvNE90Br8HxA2rGWBls
qpOmIdBFmSyZGhHhGJ7Sc/7r+H9Z72lPjil1j5JD/eyNtn+9APf4MjisyFrjAO+N
jXItSR1nGc2Ptc1JjYbeohDJic9K5l2bcWWzQUI5lINTy+jEfVM3HBxuU9UZElwk
vgUlaIijLUFRuYyKrwCkLhnvnbOfOK4edXEAsjnGXtJVyGlxQRTJQssLh8qTq0Ty
0xpYBHF+hnwmkS20boa7rDbboLFd3NaaQ+Fx+G7ubPdkftIYoVkBOpjrqeZsUHLg
/ao1leZqrT7+r5+AL5g7Xg+Vfpetj4U+wCibNfrZs8O1pi1I1k3XuxclxMY3x3Pt
aSM9ZM3sUUwA+u2yjK82oy7r0hNrL21pmrL8IqlcGKr/1IWrGJlEPv2rR4Zz3OKf
1fQRqj0wYZrOD1aPLGrJVIMYAj/sH4PhpawMb+Z4/tF/l4AUlUvn0tsyaGVU1iiR
pX87zOyZeGA3q8R+u5yJulj+m65RYlfgq1kNnVIR3As2x/M6unMdVNCPY9fRuzXz
Z+rQU0p4ixuVDUspxQ5eBpA40vxBos0lvINf+HIV9iSkMCK/tUUsE+HgsQvPxC6i
F3XG4NMr2CcjgZoqtzBbne8b+GW2scnnIM7uGsfnOtH0g7N/5RzGlDFpE2ZyUf2l
ZgRjJRHWwfPPaKHcahqT8FskbGMHO2Bo8kd8WmfT6aMekkBb/XbDhrMxeda2C49V
rRhf/7B2D7JyZZE3Xdm49p6yqzXQLlPxb2hgL8mUB3kqZn6PBnFfVKxSgQQMcD+c
1bY2j0fcWkytesuesLr+ZXXFdZWROrL4hJpnEcDrvXbL2sR0tj6FywvFNtaDhgQp
CkrkDYH35eOENsDKv5CH71b4LWeBdqyfwpFG3F082jgvGXWKVjh6u9B4e4fwIE+O
z/D3NbNdN+oQAs0gM2ZMOWxRWqPTt0K+chZVM04djkpz/FRKzhJhvIiVUCNdKGi9
Qowu2phhlccDqgglA8RavHeqIA6eNn2K82lok0GmsojiiEJfDYKMwOW3M9vR/SUv
Ws1rO/96uXVKuJncAyhj001YHfZIOpEsNTylKIS5UHP41QTdnXvv3xpaTkhxlw+i
GTf8+LyttMTt/PUUS1j8nJ0FBQy+ZB2MWMr5I47+Z5MLFGRcODda5lQ71uc/a8uF
9Ce656gGsoymhqlP8AHifAdVHyWhVLZhs5NT3E0nNyIUnthHdj9F+O0vWwuky0xq
hELdfRLgMPuTf32OBIjj5CrdyBwN1xmpxYAJas1fTH+wutSiHqx3Tz0rko5sffHt
7UejPa0UIvJqH28AF+1OkDXBCQBV0g/FpA5b14DZmVedmJGGoDDT7QQgVF+rU97W
ZiOaUgRkm6O1M9Bl73dcGpJTHs1iOBOWn3bSSVTADgQZSl4r7VchYvnIB81yxCK5
bIgLgBsDD6R1v6YdWrDPCx/mB3IwlX5c3U8RAhSxTH2nB2GlGmRxhuyMva8iv+xY
SyVnsszsw2dyTedQ+TKSr7wkwVNGHriLiADdI0Wo4z2OdtNaajUt/flcuoon6kHs
A3J+ruSabbNHg7wjVdgDF5o7l4bYMcyc8bSB/Qv8ai+noR84h3fOwn+Ama9Mceg7
XZAbGM7z6xetWwIHPAJsJkRh79qghSDw0hIea3xnKpWEJLj7tqzaBPic/u+FCATE
Pitq7kf2JriST3ItMq/Nj5Lj+RHFyqnPCqhpsH5tmLgHbIpqKqBxnnMQHZkbwhWA
YJ83+2jinp3/BetVr3ReEZl3a5RYgJ2zNk9tLNEF6esBsbcroKamG9yg9bOnillo
rn3Mb8FewQEaSyOag4gcgURg5xKJPedFE/+tpjMYDaFxtA6QezRVxm9Wr3XPxyUY
+s18BBKJA/g+Xrbr2zlak/jxLxYCcVZNI5NN6Cc3kL5AOG/RP10YulNTGkWnmOAP
QluB9pFbAfZG8832z4uDckq2jT3rVrmcdkhgcyeqGXGlJSwV5kktNeTgg0HR95+v
q6guIiqi4UuS8n8nfJn01Tw8dDCDIXvLqh0+rs0/i/DeuDEXY7KZ7zKb1BN4BQvz
1R7IZCKrSjmuqyD2km7xXxIxedKPOCTnuacqU3m/IzWOr+kONcdaadHrTtRGPgLT
0SAA/4SXqmi8JOCzgJ4GQjX6Vjh+uI088BqLruCzeX21i4UaA9DJqW/4NE6aaetN
O2VMUm/9XWjlk10WeNw6mMkT2wIoVWAkHcl0ZQORTA7jNWtLfrd4VNyv2O+qjNwG
Ge4pdl8R6Hufu740XkI4djqud8dXbY4a62mUb0N2OqUEuj64h0c6ekGdujgZjLZT
xpRSNjuZgcs3zZBa1dDhrdqRJDYtF5GOzIUtcmT9+4aVHFz1cL9JJx+3FwNhEkKc
P/+0N8dLb2oi6QkpqlxMWN1mGmYJF4oIs2oqVBwrD2BEbYp3a0LD7VH4kf8KbeJ9
L6+E9osfV3+5jGfR1ZC9fnaOUvMPdSzXm1IhtZlf0JUZ24pPld46nJzJpWdQlXvp
AGNxeRcnGAkBaaO8CYW9ILnIdxS9JRRUUy4OklQs/Z6H0p/GSl0bhjXRbSZ6tuRH
B/w5bdZ8IAj7uFsCmG6hFCh2alIAMHVAx1UUqGgtecgxJcfEFgWeRIAfiW6VLrOc
JruOB9IXYpM9Xr4IRI0frGF2mBG5XtKvng4nOSF1Z9iurmQKugjsrOloAVI5KHph
YaX+j0qSawRz6s6jdClM0LhI2+71eXsUzPYXGXOIB1XVaxpkxbaSesM0AgzF64Mc
2mt+YYJbKYCNjilA3z0rtCitpyOaQ6U9Sr4ksoXvrUtySeVkY3IDEezN7YJ7vRz7
xAbUjTszpXV6F4MgfnnDWyuQSYl+vAFXAiGGEYAajWL0ToNi9B+bV4TuJZjD1OeE
lGfS1bX2x1wfFH4hosR1DhwPw+LUXI9TGjjxG4ZgIUfRHyt9IY8Ll8jy83TtTXdA
Ct8hBqtauoXCQNg5PweybaLlaMa8pqhqcZaYcGrkKg60GNqoTg2yLi+dlx/5l66j
Q6oceGEE5peEz1NUaXZWREB0xec5TEOWrqm2uGlXJ9PYcmbkjXviTpUjd4Kc45vI
KJr1ZhSnikdJfis1qlOgTUJ9r2FWT9Hlf3UiS/C+LmWz1Bm4Y/D/pURrIrzmYy3K
bGihHwbnR9p/62CZ4OzMxJgMsWAjN2YCm6gZJ/qKumBlFV2u++ir3iIg4A734KXU
xk/KVFapQHQ8jrU0oFMzzqk8IbAQ3YtEo2n1g5A2bp/gX6Ojg+z/aFbArPvLsbbO
k5QfyDrt3HaGY9D4i9fBXje1Q/L/MYKnhQBTKn1pegKxP5rcjE6Osbf8Wv9qrTjE
89Me0IUCj1v+vMTGseFonVY5kKhiAcfCbts7LKy9ZY0yE2Sc3WI8saSJ8bjFjYUl
u3kVGRPD1G5kXLfHhyA/y4p7HWLYD7RAP4RfKTUNdpFYeobHRQkuAoAkno1+nj3F
m+Lm3gXHh7HMnS43xq5yIzXDoEEfaD9nUVryryXXW/WpmxJl99gIp2TFcU4Zt5mb
SKfKk4maQlvfgRzTVZeFDRzOKKw99NPfufCMc/9X1XJ5OdNV7A6q/z/VPJ7ATcwT
FglNOqBBE2YqVKcaAUbprOgkph35RxGUxf0QOMmLgEKVtGvuZxJeBSJ7A4x6bhND
w7Q3cYRW8SXvsqynXqlxyzKBgMCLL7pOEo6JEIe6Unos29i+NEt3y2axenO2dXrO
wXZDh0m3A4uaQGC/DTR0cn6EMArR84WddzrvexDTNogX32ac4ScC2scs3AUQ4Q7f
cvr2XTaL3FTLQdDsnd2iRA3I72bWSw2kFmghNE+XRcpEsCzAf6F8tP6V0f37ujji
dBA33TP6mRl+PwTLNU0i+GllMpiuKtSj+iOIn8FUXAdM/OiWsrUbF5f3vsEvlmQE
NeLZo05O0eaWLBLdoxPhwuw92LAH6/CS8Nz9SL3ijUzrrfJ41DISrb41y23Y95im
Lw8sAy2UHrQAWKy3zIRBartMmgyS5lve0e8lPFEE0xmVb9HWLGZUAmC8qNkmBjMy
8tF4G+B4VApLapdtMqp91FCKkyAIDWEv88efyWxugvUIlPX6me2Dvt2HjMSQ2aPF
XtkLZ6BGmvaLM33tX7Ie+T/3hiYNKzn74vmABu2guQ0oKllm2zBdTeYm3TGDOu0T
fYQUdgaMNkSXckmCY6gRwfbDMZx4GO9hHOhGHkt+OvisQbI0Zj7ImiFLIb+6MS8n
35IYexiEaGE5qFOyR8tw6tddeOqtc99ea2/MxwbdXFFV1euMZYkfSRbLu5L7zWA0
IDg7d3GuVFoc2SkMkmCYcjWy7ZoFRzjZLeuAfqcJK03oKDUjrMiYa5zgjrh00EvB
HJbI00H/fZUuul74QQ5X3hLYVt89yzPS+eSTsWSd0r2Gr+UJF9sUjhzmGd3B9BYM
TeQydxM4CBvFrMvglCDk4SWwWzyw4OE962SOQDthd3gBCNea1zzfJp9q4ZtcjbzQ
dM28C3lhlG3iaHqWPgdSClrpGrTg1fb160dUQQEF8EFpzoOc00itovSLeMrx7RGX
kjj3CetJukF+Ws6LNuKrZClGnvAh/RBCizserQvIuJnFao/B7YI+65qZgKyoRUF8
TuLWiNfDCdfCICd99/6RA9kQsO2VxUyIEhgJB6X15Csq1ddpgI6szzsHstUkTHFd
4Sej7IxCCTCa97t5x6brVlb17Zbw2mCEq5SiEODsRz3bvQUkBAv7B9/pt0sv1Kgl
UGcUBN9NSVpNhcGP6g9EPF+FUDKjc2dba1YOkdNDbjLeWGRcgvj2yfIE1zgWlE69
jyyStcG94F83oYebzqbfPilEwvw8VH/WMI/Ty0dcCDKoOQuLBhFFCRTpwX3gcXyE
J+mblWjcOE/v/wuOpCfXM61WcwThNX//KwXHLwDZmArY2xh+otX6L3ccgCRMpxYu
ypDMfgsT+hpry141G8QUufV77RsGMlxv0LOVGuY3jHEL/PgiTgHIt8kfzxEqWQd5
nxlQHUlBB5XyUwofbI04Cq8RDt/bEWiUvdyWC9XEY4cS7jxlN+EyqVAellHIVpQ7
1anO9Ofh9elfPa4pkvVpxZqWQOHbl4/cl7TATkovdMiMSzmHzBmvWWhocqGNKejQ
PEn3rX+pbI7u8UjGlDjg8lFBHCjW/kvvgEuXGVFs6gII9I69mOMdVQaRhqDxu/jz
fsIEx/KWi3+IbJanA4OdimEBPxoPB06Nvr5keSfrfgGeovZa1kJsqRD08n/LWjx4
XHidcaXfmhmNNQqkg+BlQFcCwLvahztBIe2n4bFKklyImBTllbCJQ/hXbOFlTTBU
76SyB3gYdCc0nD0UwWf5a1Dy0+xOir+Bw+9/Zr7BwDyb0WWz7/GTQi5L/zFkiMMp
pU1XGHMGXWi6A8BvHkLDgOzT+illm7/insdHkkhac9HnR93tPJdvZueHhg5GfdRs
669G5L7su5Nepz1veHFVXuEHSmkX2Wovqyi4eVbL/2n21oizpWUmdgwa+wFs3fr5
aQ/Q3douF3sMmtaEZu/cFFIcNsz8cw3rT/zP+AGAWVgFHgdUwc/JzZNL1RSeGiHV
YqShP4xPG/xZ6LSVuzGeFx2kAojAYv6CYk4CXwpcdeDpCtrkVWVekO+7HY1mu9xn
cmAjtDA8EIhX+jeCX8A3p2YH82HIAUgnruXq+vptXYe6No3dVhTB3DdLul4cw5bM
I55GYj8JAEVKUfvMQwz0oA008xl8QifL0TBivJE4pJfKkFvt7ArU4uAd+V68Zod+
13pY1qkmsqr0pzudCoXP0UOYuo7PIYiIRuAHpI33QI/4r8r+oXYoKIEGTtOTVX43
QCoNTSSI4rLBgjO9mQWvncgUZOJTmeMCX6Kd4EQSKZM3wMtvbNPpfA5FskZzIjAu
wzqINJkrquraDfk0vysxkUAOqNRbsDpmdTTtBsEKv6UMra/s4gI9azNSyXnMHjCX
DPpHgyXh64P/f8wpZFP+Qzq9bqDDZtzCrPIlPuq/aAB19aJbnBlBO25NahE2MluG
5dFySShRDEU2CdfAQlL6TVs0i+hpDBnDFB5ZSL80QJOYX6172yJURETqLy9Sa9wg
FGoDZFoUDLf3d6jhJQBdmrY2/L9ECkQ2WuvrChas2wI5YLNJ97V/yum0PsUlpK14
Rs+pkyRO7hdqvsbPQ24VtFsfHJTjOunnYKWWnP6sNfyDr7HmurwtqIRrVBJhKVn9
li0SMrv7MLWXFOoyvVYUZdEqpd1je4prcMdlxLCmfmixjrY3oAZwovqqxcr2JLBT
jH29nmqZzxvvHlSxvdIHcuaHkK1194c6ui1Vml9YP3OsQdo98oCi6Dn8EJWdiy6O
l2mEt3LYfALtLs0hmVZXF1bpL6efESYyhAA4fmyQSn7faoeh7NJ2OeCp7ctcRIrf
hY+WaMbEDu/hCAGHc825XjsPvH/CrbnnlUmTtFgLdKcwr99GqBAQYQOuujlMi7LJ
i1PDMVbx5MVMwcdlViQD7d18KDBUlsmPbIYSO7rTLHqekdF02sozTJ5uK8jrn393
JWB7Dyht7ul6+67pUIAPOBNVxuuHmBfq963Mftc7Dn8inSCmTp/4S4AZWj8ClJ15
sr5inbqXKkcB1+iq5v3i5uTYdJrpUzfz5TYxsLVWnfkXbAKsFuj7+iNVJZBQtcYZ
LHN6sKDDwvPIwymJw5dQvxp8M+33arDPjTUgZURAxMFMln1OwPioOL6hwKAOiUhd
/fpT7WKaSSfihkqctS66G8MVm66MtuIv8eemkSH7+KIFW7LkSlXQDhILl4ZXbKZt
6/dCzqsMHJmn749tW3yEGvNVmikt57GR1vZUufj+iv9RmpNyDQcpL73SfmDCnTsf
nL0f0U/0fpsqwl83KD/xWnKwNnW+sDUvnPeLBZGDVzWU9c4Nn93g83xqtj1xwRro
Z7kh5XlXAIpKXqV8Z89KtIot0ZCjK7Xcjz7tafcKrC51zp2VuLdSGu+UsNsGyM1T
Fyszv0P5OipLaYV9d+u/Sz2ar0YgN92UPx+fEOe3p2NOEdxyr8Az5Lux27pU33qs
YChWDGSyf5xg7O79gvjzfmpG79nipDth+0ed36/ekgfAf4s+NNk8OTZe5I5Q1jEu
Soyu6diaLO2LusCH8Ak2+XskMeb71U6GZlemE6G9tBSu1P347yOGJudP9Kf5QiDP
t7tgRZbFai4eO37VcG2zLNTqUuYtlCZiukReXKqfo8BXkR819LsXufeyqnRn0POi
cqQvp7WSHVAW0Oa3iAuc1j/BVF7uSzSnISfnd+bLweiTtt/B1bQ/DOR1ukCMoAC3
RvJsu7BMyMHojhDrvx75PWWNw3yGILOOvERMQEgKseATecMJ5G8O7tTE98oh06pZ
hNA8pqt9ZmY+GVSUts5seYOxJ4b3OEuT0wA0pGLIi8x+Br5899q+FGJoVce1RUMb
qJA7uC59v6gwymNpfqtiNo2MDTZhcb8u+etwF6eWK5GSBQ5WPD37VcVkjWCUqqJm

//pragma protect end_data_block
//pragma protect digest_block
CnO0tP0L5CI2g8Nb87xVoecu7tY=
//pragma protect end_digest_block
//pragma protect end_protected


//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
xHFSsrkAJOC3bDZDlSfuFL1/OGVVKk49ueOHpEDbpqBOvmNChJTKbvWB6qY+oVuY
GcdbADqMu7aVmVXeUI6mGtO7CC+TDlMdc3NN3xa8/7FdYZooVVHL6FQK7sxYbmrB
hoWELduE014kfYbnBBHZce0D5twT7YhbwbXgctlpnANYg/NY2+VH0w==
//pragma protect end_key_block
//pragma protect digest_block
GcbrlLKuix6YbtUgV4oV1wf2QJg=
//pragma protect end_digest_block
//pragma protect data_block
WWo1cf3xC6DFviTDt666WIQra9nDZY7XKO7/bQ9keeEtR8ah56UGQPjsocgwhRoB
ZQKJe/uDxD9VjVJVsLtLZSYaP2xR3CBUdnjRwU6uJ3nIJsV8gbpZaHmMDPNqzc1P
erASVVeHrR1l1jiLCafU/jRJBRu6Uf3IV5/SICo/SYdqYo/ehl/EfzUgC/SgX5g7
N1fcfJDgpcDScxj2h9JkomWMiYB9cCzGv+l79SKC/p6nD9vViq7xTBiYnOjXyEUS
XDAnmLzg4NgDWUazfdJ+Y+1+X0IC/PCuHtWFanAewL4JlXvQROA27tEpdXRyLnxm
1VbYq1/snQtiEfMKYWBNbChkcCcGp75H8gyTGdkKPcVuikSaWGPAl1UPH5DS5mKF

//pragma protect end_data_block
//pragma protect digest_block
qS2T481WuexXyWN51aXLudv8j2A=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
IsxntqbzXioCwfDWck2cYexSuPww8+00Tckn4LYvDP27L/ozA/xIng3s/yfmUGh9
uakz1V60Dj8ekXgjPbo9tUb6p/6HLJehFsXS5OOzCDfU8SydLPKsXPwDMMwTbeWz
Yd4PoN0M9J14v9xmK59Kb3XU7JVL89Q/K3thbQJ4FgSeMhTW19PDGQ==
//pragma protect end_key_block
//pragma protect digest_block
tGMnk21j0TBc0uX3XM9p3+fWl6I=
//pragma protect end_digest_block
//pragma protect data_block
t3UTHyxARTfe5ewE3jxWoK8EmC2YItkC2WX3aIB4F6NhR2arhAAl4UFHEJfZ4Wa6
Krl+h+Sg1DCqL1J1hzdGluNTOvo4mO35WSRDXrUJC+VWJeMA66jzyViZeGJkmYzQ
pkTNWrlMtF8Mi0o9xaDX+Fxq0/tMAB4Evrj14pbjFfbcuY8bQPPqLWyRjyBsUW6n
iJGYXmcDzUfMCJ5d6ehBoYBr5l2qSQHGb+e11QN4L5dIqPEEO5S0HiYc/dgTLocJ
QZofphPbGM0I5sSrfqbG0dYwDTtrBTgv213oYkDp7L+CpF70lklzSVUkIqm7y5Tt
VyC90LwMo1HVFodqnI/MxzWrxVV9JqYAJwC9cza/1QenPMtBgyozS1Oq9UIzkSBT
WUuBzo6DvX7EbUMf1qpchEf1Z0wr1JYDRKpbkuzECh0CXzgEfjcQZww8EzZ6k2HK
6Pev7eiS5+uQyC647MSRPqmCYnl7ca3TWA5te4q62fQZEwYi2aGL+NRnhEYV+rgd
Tq9O2j6MEcRWZgwjDQXpWynjYMMak9LmXr/gpMB3KXYv3IEiIw8xQTgpgUjsM6ey
S0PmJEqGaWbuECZeXYz2f2w3pop/sIESK/iqtegCWQnjDUyoqvzeJlV07V+aa4za
z4FmVN2of3Ov3dzYlzBSIbNWOSZY5O5gzyya+NOnBR2MlRoQTSY+iC1QP/wg5HcS
N1KXfMXBlAEGaVx9RgxAm7FxTqMaRLdBobg93h+yutPMPzdvWJ5LUsFTgpcN42J8
vG7LV+K20kFmZNYDRI7aJjGlEeU5bfLZ8lSr4WF/tuv7NZG9d74GelnwgKo0Qhs2
Ccf7Ssg3vo7XJIv6MNdrCNvZS8+BqUIdwf5QyJ1XMia5Hx/zPM1vX3GFKu8Cn3FW
npcWaB2PTMtscxwwZTqZ+tg6N2bQ1NKP8GASUymm+ZlazO8wLuaWzcjDdd0FGpnG
d6xPkV8R08Rl6Qt/Q0I2fDo63IPlEGmTW4Tak8k001LKF4iw26vbvhy3ES+y1nzq
po3EKQ+RjysisbLH46hvBAgRmfEHGDvLVDTh3rBATtcf3l0cdV+vO0/TQY4gq43d
9Kb4hIumEIp7WJPl9Rg1GjS4XtppqwqhEVDkhMvmnDnAYPCw/85/gtgCRBAptIiv
CjaXC/hcQBiOHA5o1tFIHR0wxRX3mhzMuYKbEcq87T8HiqURFvmftXPWJW72aW2o
8SMpjiLnbp/HPz21aXlAEVX0wCJDP12xz07PesMsWlRJCNdQQMByEVHXdxe77loi
sh2mNufPl4mOBAYI45MrE8+q9HbHJ2Hj6LsrDqPiuAdNqKXghAt8qaHvRtELimhu
LvwckVliYaWz/yOfxPoVSD6ZP5taqy8CwLmJ8vqrMOtuaDBXzTnSm9LDLumrA5b0
40GtxQlBT3ZaT09/E7ySuVOYuhv6qrfub9alXzY1Mub14skQ+vzHDWA43dPpxJNG
YfijVelGmU7Z/wP2ELFnIPucKecyjy+giXeGz3ndnBbctugMmBhHk7MKJFoLSZQC
RTrTO+uqmBOF1tS6ZgtS2LtkbhI7IEZqF1PHnobbiDpGtfRLHJmBilnI/EbCsbT9
xHW01e7g81xF6Eb5udZSYXgBzThNlzcZtInqK6S7eBsnPTW2pfalb6xadY+D71Aq
aD6ozgZJGugEJY3qoKTKsH2c/e7RtAT9bDl3jZUWQZnQG0zwEXwE9K363QK4LPga
UJVpQkmwSJUdl9K4MP0+2cPMWrxGaXVLhjKYh4oRBE7wSnMv3rJWbwKdwjdoPNyT
h5TfRG7Jg9X8xugq8wG1mdhx+bSsdANXA5r3eWrTJurEvMJkiiDru2W7c2LNGk4d
UfC6hN/zerrxyXWhEHSXGDuFN1T1gm91jAEj2ZXvu2y2N1vMUcOKdfDkbobnnxmi
++GHlsSlJxT+IZftPaUM40Qt81SoRgXB1thSVbXGhLlmLBwRSPCNJN+0C3umq0VD
yzdieYhP8D8LWt6tiHWEXV1CueqeN+9xLUwTZgNh5tK0V/URhNVZTtDgVV098pOA
ulS3GrJ15sGsziE515p1gt8t+EYhBT62Kbt/9tdHljLMtrh6KyJ0ZI5BM4CNpdmb
bpEUPEW5wGucGXvkM5oezyDYU+crcR1ZV+sXtEY217kMer5rj52L8UckV8KhcTBX
fHLTftUwzfKxSwdJTUNbBLZEyFd3tG247Hm+QdQ4pE6F3KD4yNmLQuLXRRwSjbmO
H4/OX/t4cyQBwFgLAxrIQLGSSpWPEIEGAZ3VddEI5ruIxPKdXlNVXA3+HNAbkdXP
AIvoRVCSJV3g7ZV94Dj/8yZydCXT6XfJc/3KzCj6s71SK3AQ8sO0YRrC3aaMd8pq
Oim+hUPMX3eXxvBt+n/Ok3BNY1rUlHK1Kvlq8Mf0mZBmhk0H207ZOasUdEEnnn/H
PBmwPAzw1Ti1YmYkT85LMecZOLz59Ettz3yysfNR/m/S7vlM56UJkub4RjNtWhRY
0+MWL6jNTY7kPkDWDJeiGnqH+BImglc82IRghN5NYt5zJAk6Gsn2D2DEx/Thmw3G
WyN3QA9k+rUSCYUlxpG1QY9hwluQVgJG/rN6o0g2TMzafxxU71jGCUPnDyiNfFnH
ZhuEA4uLG1gN1qhy9Zu33X4xNo5+PcqszudV9fWWWVH/ag3TYWo6OOYCglLNiDK+
k9QXOBpNsaUWWWrEJOjdOwFOcCZD1tgV0/JyDCiDpgme04isFkh0tZc2UprYQ/aG
kLf1mRRA2ybK5XXWSzsIAuThtV0NwE22N84vTmg5zoKvmAz4macMDK2SbnDOt97i
lhRSpXOy83DabJb1JUrtn/JC30YGvPs4cs0/DhVw7Y4wCTu+yAYtfDFMs4AuyTQ8
VcUMT0zW+VDyhP7qfdU1qGknIESXRtjEGHvB1Qp/KU02HxAcZkpt37g054LmkGQS
aYKyQH9cEo9w2+HmbwnnG533cfSXUUayGmch/OLgg+K7JrPpun9kiqNiDRW2GySO
mY74ppI6xzWFdURuSkNkv+PM84aKUy7ObHBkx4euLsTh0DdU2rib9hmZFw80++7B
Gi53jvtRBf3YTKKFJPcyAJdDUV7agaBIRnb52tavhODA+h7W9I1JlGyqGTVOWGiK
y+NlqM1qZ960+P8rMAUOlwXSPo5OSVZ1BbW388dvJv10nSy0261kDujAYFnaWh2e
rcgg5sqnHwPlrLWveK7x9Oxqi/oabj8M2r8NxYcwlMZs4LGik7ORLzXxUebjwFMa
JU9antdkaWYTdlenPuHfWvCn71sE0uWb95l2RJ49By7674zS4BYJLm7yDRZaMXgW
Tty9oEANWbj/rlpCqHfxVjU0P6GhkGcTgK/490sC61DY7FScjnwr1FpUhy3APs5U
rBDk1Bkc/S0rNwm+DKlAF12sn6iq44RMpf/LoX929btjKxPTmBplY7aLG7YB7s35
vdKGAAHJHPba8MiiwfGsweSHVDk2OttNLgOCv5Tnn9lIt6B1NSTSjgRo3aETtTv6
iUN9JMCUOJm451mEF3mSQqbnbAnJNoDfp8bAtaR0X9KrfI0QzdZR7K+stSPszdN/
28e+BDHbtKRWxXbQrwz3n3Qnkg8ce3GS91DpI6lgjod7uliXHNklMQzoTdQoh+mm
tfZBWGBqDTX7lez95jP47/SzLxrGmnJT7xY6zI3kQhypjcWMgQZ8hfeOrvJCxUxE
JEThzuBbypX22UPFoaFFCfHgnfSxnxRYjS2b/O4nDmZzIzCkJNi03Mbuyy0T4275
w90uAj2AmQKMxgvoefZY/Xy1Sm8rLs3U078WUXte0b/A72WfJkjOSK89XvLj5Ggs
vSppZZqga75/fgoyxqOrPj3sAhlqJXiKkd9ETsobT/9YnNABiU/YtYCCTgZpq6ov
De4oIIwYHOtIPXLJnhB5EYuEXT6IJhKgm6Xm8mKE8neWC9wn4C+NjxGKLHrb59+l
ko8X89Ho9sZx8Sfj2WRhqJRpjragpEqN0omqUBEWaEbBREryywWvngMSq9JuSlJ/
JroaWOHjgzNwUCSDH0jIPrTB7L3tAlNffA8GZbyZts1hhm9hGAeGjvRlv2JRno9R
Lp2eEoA+cu4tQDoKJYj4L6YGMmNNjFp1TsjP1zKuhQ0PySlL27b4lfSKLeycaYEY
A1HqJw92dvULYkZBC6GtMTR6mUI9dTw4ArCZkeFt9ASTcKxX4xVUMaKDRmCIvSyC
t5HspRk2ysDU6lZ7d0xF9/9cbzlZwO9VpA6ye+dTO/5fnel+wjk1unYSKk01gigL
+7wTy81qrOvE3qDNHewSprYOKw/CAcNpFXOHkMqMvBCvlbR24WZpmX1s/LkdIAU4
v/H95vr5fDcFoD3O8hMvR8YEZvLCVkkUKOGj7Tm8VfVwt6ayNH7nD8fkacGpTMGk
Gb73uiwRYPmsfX6Dz95O7uzz3esTHQZjaTebOqylPZOHYjUvqk8Ii5HXNM3q+Z5Y
LrfE6vWoZ6r+4Cbn199cV5Srv5p78cN4qFw4Lo2HFguBkuOTWkw/SQrodhF+NNaX
cFysxHnoWa7ToHTajtKR+2/+sGKI54+sT3XtdY1PUZToZNZ2Ednl3/tc5dUrkCt6
amRT5cXYObb2RMN6aztwM4/k5itYIDVW2/27cz00SfS1HMkbejfmd95FhFcGUZ53
PFfWemAb3p1dc9gog681DSQjWQdB98A8FmaBwF5R6zxORMIyMcf5V7rAxS1wX3Vu
ssPvNSwXqVKsEjE9z5quBkGeMRb+Dwz0exaxWYkhQNHgZQ9kGR8T+HqTn285I3sC
E959zDwdFBNdakga3XH+QkTuIGXXwUpZ7mMg733jhHJFti0jwFtFgrMojK7daYKT
qNPPAHis1vJ1WYRyBapjrqDAuOY8+sfD8LNAuoOTeQYhblGr3xEFEzyaQQefo1bV
zlGzZjJq6LZZ9gS4RCkAwXzmeZZDB+YhtpvAmG+HcjQEGWAJ2D2nOE4IMsGOzxgt
HiP2f3PFMd0KEuSnt97ami1v3JZ5J8twXwNHZbMkYCEtUMOhxmmXn1/zt8uisQqS
WrTmccBZy02UcsoP8utXsTDrBYbHbggVZzqUcYCkWak0K1MhpgSALaHFFctK5z+0
A2GMP4LPhxyJuYRZHKYRkAEhrC/Tj3Z2nMwAmz/kDHv9b9JG8TUUl/ghxbZEzuaV
bbm/eG15TcJKiuxu3cgTJPr6+u9+lyCO7C7wQtCEcXUmkZMh1hCRlETsze+aDzs9
85Zw4d00e0uazMi9x3LqPxAoLWftBBr+Lm/SCKyowAGXs9daVdCKYNudOXnIAbho
ED77/C7EIuswMvliMFqzWQZi4e/Qr3CZQFnGJteWfzerzlAsLsbEpyCsOrnO5noy
aIgTCgBmFKy4Anbso+oOMJERThl/OLzuVQ6y8XjshhXrNA+qkyCHyks9WN+I5RFx
Q4ShXrJT6BYTK4hCRV46W1Gyw0fMZC1LNZE/JztmBIQPJytnTda1MHA+0P92dBCy
COEzWzqhxAJYzGgBl2sXWWPENOCSQXVGUkPmaO6Fozp+UczaP8fgXd63KJXxAC1E
PGsdFgau4rFbDtRuco3raw9ciKk8UcIsqw9dwz2JH5MiAyr/KucZYI7gTexX+p0x
cJDn/M3PYTxh6/yo2OK+wZJiH3w4KI/hYfehakYzPLNkroaij89t2nu+VeD/A14b
X6ZqOFFjkKpY+qtBZjNCRw3rZteewMPSg2C+VYwyrfZn+/y5lMOvrKS0JGEDFLE0
GIXEXiimtAsYHV25dVLiYmUGK2l4MBWc88hTPTUwpZFtWeUrDDDdkE01ZAbIKP3B
FRfcJf9k/ZVrI4DWCRToRU9DkfTV76B1tEFEkzAiaLbYfNHfZ4BmaoE24OFuOCW5
ZzyCmMOHsedpvlwTDR1L2VjkvqyolNGguteJz1yz9qJsHtqwMWgjQc1ffyJ7gUav
+Qux9bHhK5/ADTt7JT87XINWToMzw8boR685t6G44qf8w2jUi7I4FXbSTIT5sqBr
3C+Wuir2IHinzbsFizOmG/ThUpl+F3SIfM2wt8KqarenP5Ev5Wj0BAuAZgpTcHI9
PakHSLTPdL7Wu0DYb8BLv4ZWVu3+7TAvBTVgSqEw+ywawSd5B+2L+GenOPPlNm9j
D3oKwRxxD3kwQnqvQXlrPwUIaxoT8hOw4V0WDCjlXKpOap2da4lDlk4vAZBQfQJi
BddwH4vcS8LEdQnRvhbQxKIYRZDt0S02kitLGUGX+G4z983LnklGu4okL2hNL+v1
4J+zb1BqSm/AQFOG1yXu0Z3vwvhzgNCPbd7Ae7OVWIB2WV9LygxNINZp/nCr64Ui
Y3UZjW9lDSGmHoPXzzcM5yWZWC7XVQhMkY7u0Z7qM0tI8H2IPbalrYnbo6G4I1LL
uH3wYdI6k1mTpWuTO5oCJQ86Dn5CcrKTcXKiRrpCjhKyGl+/kUbeLJMHfEOcYs0O
dX4WYgU/43z330tOIh+bIjVpa03KahNrqRsk+HZJBxgFqpq15yRz3mHzi36uSumi
KCjW2siwj1A4SphcFErVd8nVqKK+Y+ampaTqLjDGuepXlAEdGPt4LciyYGQ1GwE4
0jlOlotVzxkf6nAWRcoNQzUWG9aKYWrJiRCxd0fEKW82RQsyYIHAZfVXTnZVGZ2+
XhesJQkZBcLMYIjzFPJ6mM6J2g4aPu6xJ4lwWkQlzGG948kR7PI6Ebye/54YJ+Pa
3YBHimQ/y+f+Bq3JWxCkGG5ONr32xCTQnmMMSGVLNm0uYgegfEy0LCEJMYRp5v/4
BHJQ12uS+bTF1x+6/Hm/dI5Sja64bvdeCgJfN3YRi/dTIWjDaXPzC5wue9Am/moA
w5KTnTh2TjbAs6vyG311SVpmtkBRB1k2/t4323f7kLb3tQlAWnNAWyT/LBkFXw/w
gal7If1ro9vgSIg0PaNiYjbl34jnW5lVQX3+buKzl7aJBMY+CWpyNSZzdZ9ZHD1p
4W7hwmf4foL4QLmyJEpDYxpWpRs2gdbiF5oVsZX006ZBs1Hjzuk6Lj6+nUqM6tf+
ijWX99xasQgW7gOmEKMpx/3S73BCIRl3iXo0680a1upISuy8HL4MxWC/abJpLSnV
TBp1zwdSpZvz2XeAafSh4cOfHxGJkUZ2T498noG1yJ4rcsKmOmpgIh/tKMftlAEQ
RgsXAqgjhlmi6SrEkZtLcmORwyCCnk+nn/hurwDoMQcP6DJd9O3ihJpARSw22wjY
wJUK67i+9j5cndSG5gGsF+ryLD5H/aewbWLrAeOtXW56iq8dl5+Slvk2QXlvjf0+
9IFtuA7SrE6SoSMeJVGodS+D/g9hSN6nIrT720FtB7UVqD59mgh6Fgkzjgalolsw
E9ImQrQMLbrpCUQk6ShA+BHCR7+t2iY8/8vB4YEZd72DmePnW38v13A2NSJ+881A
3YM7yD1rJj1qWqFBO1cbxYPhgTv2Me8/g5RkrjYe0ZGPn6jEa2PogXS3wJXCVOjO
tJlSnIYqjz+Gj6wtzwMAvUsmdwgYllS8+KPBWNt3WubhvKjZhQmG7as7Ahzs50Gf
h1bl0XrqcR4rHtY2o1NDuCIV0XNEYls3bF2/dn2Bl5tjKjwuDDNBqsU0O/A3lnZ2
lF+TX0IinVKO4LlyybDkCI8lTdcY3p7TskuX+JNPbLVfvfoK6BtTLHFVV4XFcVEu
mWZdIoLsQUcF1U6xG+fQTS6EjcwIGqjEx6mjXMDa99QGpVHRtJ+kKg5d5F7q49oH
tR0AwR1SIFtNNcgrUGmGepvlOzOpdMvgA6jgoPOJC5ECc0dYDfm2+AFk28EXOb9Q
kyPjYqK9lSBWIoHnJHdHUf9aJZJeL1aL+FpLEtCXV3o59kOaJ7vAAWTqW6TPFdto
O4UcwolngjGlLDI9SPVgbaPKglvOvCEsZ1oVt8CXpnTtcPaoi2sDd8BmaM9VC15f
/cTKcorD0CDevGn7PDmi9Bn6uqoHGwqd8iR7c3Dy5P1IZQKfkqG8BP7Jb1g7Ha8N
wyWdaVLyqMj1EsM7DaYV+W9gmY8o/htbUpceerno2WRbeaNLGiqLspeBGJi+zwWd
AS+fJRKtb4EKiLQ763u+urG8uGwG44e79Vah6Ea1bG2l8eDwlZOSLxfjYi29VFDn
ZB7OceGvXaAOoE0u9SgTz5eTWQsKnNJU0cS/kZc/Oud6x3ch8B844i/UkWjY+9Mn
pcvxGu2AzAQlkfBxZI+eMRz2yfoVz89WTmBacKdjjFy+J4ON004QuWxkfCoInrae
6etuHCzyzOjZUYxUGjjmeWuByWbGeqxXpl783YKiAU2ftkh8U0rdms+jJYBnZOsI
c8fBt63txCMwbzSl06zgH6xv+QXuL+YPybItdlweq8ZTSnrttf5etLCSSbj83Ii5
Y2mc0YurSI2Rl2gmnP0HyLxK9aG3Rotyj5xQ5fh1blAEOuLxxISTXi9KYRkb/GIh
SlIOMOIj61soqMGkzJPSiMQIt2tWytnZVdNj2gtV2706GGU88T3LtVSJKblq0svu
C5iOqhyaqZjpCNE/PTvZkK1M+7MTynmL4UdtadtVv2ilUlPLLTu9hGsEgQV3DFjH
9nZlYZJxlNnFX9YPpNrzLiMmehkBXKKo8kVIFdTaNhRrd6/bLcDRzUWZKB15Nrdx
zG2GEciaFmERxqUHjPHdJ5v3SWyf6ElFHBb4yIy5HAewypCbFph0KJNqOvq1nhgO
LaS+PboghST2txjucG1CFncN3rNksfM/2HnhHAjY9c+ENOHpc5zR3FP9u6JMKAv5
OpaebRdMKwZCbKZE5DVbYiJFJYsddiTE2pm7TG5l3IRVRT/veUQZWdx12N4HXuzB
LO2Mb3/3tiMrQ4N4npRhuMZV8BvivS3IaP2QtyQDIKUW/uXcOHCc1FKJ/kUUPrTv
JUyiwbyZQrrxDuEOj5pDR8h9TmLHkvF8u2szvEC1rOvJ6J9fcdHhHfeAZFbrSWAm
f/Orbf9RTy+Mv2oqIgrki6vtIlTh69pRzJLvqXDS62Obg7HOpQZAiQ5ODoXwzVkV
8rAeln3R0XNYcd2g3rHLSBXl19GjpxdCZLLOLf22uYXpxkMpnXCyRMB4dgsn5I5X
qUDxd2lZUOUkPHRP42kiBbT7cbNNOrBPrxgkoxNEUiQxWIx0d3sV4CqOJuCb3Ex9
T4ty6zbKDWRZT9H7BSoiRf2ewlG7zWYeXw77xpRUG0FN4RvplMqdH0UN3A5TIIje
yhsTheY0mZOq1uJM1HFOC9lz7kIh0E0g+pU/z26NIeuKFtRi8ltLVV7PEimDUgwZ
Sb9nTeawXGj/zlQ7vCNnRYvE1MmDFjX1leO7Ir/SPeQV+yU6uB1abUtUdW7b06X/
2qkQcFoZ5ufCd4YaHFbzmvlzF/5M34pYrm+EFWGP3FWNm9tOTJpkyiPOda/u7zDf
6ACr6IwKLaTj4pzxKWr/3bYwQtlbM7G2AnxVhAgXhG4zJC8W7hjMEcL+EKF9S9qO
+WrHrFN3SCKe3lW9XZD+LmbCTKM0PwH4S5UWgNpQZ7DumSjZ6l2lQhK+eUUaBTP4
TAEK8sB3cuXP7enhSe+Ub7iDG6bteWVQUSC3Zn5CIHvL+SoqJnHIWPr9yeQLymeY
uAyyEQ6HgQ7O7+aruMfusYiVU1mslDORcbhzyU1PyN+bWX43Ez/btQHExqaRjoIl
tftY9lJkSptF20MfFuOni8KAlJAKzyQ4yDsWmh2hV9/1OlFosZ2ZK7IKp2iWu2RW
XrmBeUpZCnLuNS1Aa81l3rR64zBjyaBdlnbWq9JYHmq25D5JFfVVgGocm7Kp5vx1
WoI6HGz9e6F5Ly9jVU0zvaiTVdG7ugTGFLwnZmaF54OIrN6UaviHf0ZS9ZO9dlaa
h6w2YQrjRCYzyRpCl7wU3XcsqO7liv5bS9Q+9Ih+gH8VTvdswELPhjF28qmxc+yx
sDgy/D5Tl+sydbP8QTyjyU5xI4uXVsPIgz9jCWbIdQhwBFp98KpoAQBexTHTITXR
qqqUw4lWfJzIc+PNuLjLGIHkv0lHZMoEdBMBofTvdcUPHnCtmkiQsa+bAz8Y5Zg0
oUR8aJwFKUGf9r1bhbT3Sjr4hRrINt25L+1Lmx2JvwVRLeuBz7Z0Qfs+AHpnI01v
FoPNuZc1AAOGd+BsZ2l4Ik8AwIeutvc5R7qSumTn2JtI7LQXgnNNIT1h1OjsU0/p
wfcMH63USe7Z7EcrS45/nwxx/aL1+50YY0hQi8mTHwAqewIKQ/ICfuEbMGJwcFVE
EtW/EXULoBZTRt/4p/d4Che3r/rela83qIxd5hUUWVekQwpCa2YCW+21UJMMTtXk
sLzt4mVACuMdKPUM/+e2H1GHRQs+62ZWo9+l3avscHRRwACHkrO3ckwc/SIY/MCx
JoMIdpOYzN8guCkaBWIaQMNBp+FSz9YKOy+/RJGM8SzJdQYehFyksu2jpzvG71Bo
k5dJdmuVU0iq/l0tyB4PrNfS7AxpfzvB6WlOxJOxaOPoeZtb4/Sa2ItHkcgmp2lA
L3QyaYrXzebM1XzVVSxjQuI6lxlExM68KTBpfIyvEpCxGNpm83T+bdD8y3iM3UnJ
9kS8Q7PlgCZsrUVN9kWHhTn3dCrnXdM46Vc422KMQh3hBlCuMA6IFjvuxaZI2PnD
tU6n4HIViCVzJ3XD+fMI1Svc4/8pLuD6nzyH+qsQDt6E24fmIQWM+eiLmrAXKFbC
nIJtzJNeAVeJp+saqvwiwFpVYii2lCjTgXReGIvdi0fwMUn0mvwDNH+dDkmHEnrM
bTjmHQqbsE4EvqNtnYWy3F8tHyxN9w0uUiUFSp+DI7wX7weiXmK5rPM7OcqS70Nu
DWPAjK2N2DKcnl4rSG1rZ5Z2to7S/RWC/DeQRkGCsw1no2iiBj4Nm4necYxjVSod
b3MCP6KtIcy1nuEhjaJQdsWPYfJ/MVc7egTMUkv/8gDOaSmBGuU0ABF7z3uRdfoD
TjTx41ZURDjNqKzW4UzY+CBwu7iRm5TWlSeKzZubVa7BjleYYdmQ9+gN+BEDdokO
cnZCVJYI5XgqTlC1BpIhtVDSr/6OZvYLJHG7yFVl+CKlDmeVxW2J9o6Jd+gETzS7
7IutVhM9a7N1miDUrFYL5YQmjl3q7c+U3peO8B+0NjfPo7BcMfu7/ft6rOHd3cIl
FslE6NEPSCoEMi14w0HSkIiOvLSKVLssj9jh7ZRkV3kKzC5NqQSZ/9C5584cGs4H
CWRIkYBdHURvJl0il03orD2Pm+S/YxF+Mv4m+X+XHT/ybg0cppQBuTXuOfRZ8tit
XpA4SQNbFQ3Fn4MvPZn360oSWTALuvkSg3vg0SmDN/BR40Dl/2GWEqEbZSyIEMWK
pvghvl/0ebeZf5kpfTqUfG927ZI6ayPQ371PMdRdorobvkprx04trVWwLtz5rXEl
j2vua84OVIkjrh0Ouqv7HYbvR+uPfnNpqFeEFa4j/gf/pwU88mZ6e9Gk5cyVhE2l
ZpBHCwZv7c0p22a1+OaFSqhWixO0rySf6LuKhYHGhVk8vQe6b0/3GyM419SORDGA
sjCNdUC9fwYXDs8xtiozJiaFHV2yN8YdU0I6oTgv0ZgKeO4p/a3442XDfqBa1upt
LjeUGGXs1+B4hmwdFGjzcL449xLLfEvnccuqtwPkPPhofraPrW2B+wrmiFeSzbyM
Zcj9ZzN0LXJJyGjXrGhXjqjD0IZL5Ju2lWHyBMksfoez+roBdadegQsnVldrvFi+
uS1NU4xMXoP9Yf649gnX81c4wlu7DTbc8b6HJZCah+5GTsRkED+76vDgLKHHhXaV
+a4LUexhXoNa3e+sU7piYykDflik1g6KHFFCBLiU/j4HoMf0TiS3ruWz1BsBtKX0
d0EMAdSs+r7QboFoOwWk+8KnUcr1XNtJbn8xzuxBJrL4AMoLHfIBWJKaHacsS0/D
0RGmkMPjn9thsKN1vxuDJpoKdtuNRCJAXccOazTzYfV5rYyqOXwTwvvU2c4w37oY
rd2Q85kAq5wqv/aL4hQ/XedVX4Rt2HxvXdM/zm/mqBM59ppuRVlWzBbXGIENrWuh
qjuEiUU8R3e9rkg2TYV8nKVBwi/d99VzokP/wrwmbmAk3wJ5/zM+fskQNMeek3wp
wb7YGH0W4akLKOubNck3dIO0YAiK7aPAqOfH8c2x3Gl9nQ9HvgPpsPwdV2GwrYfc
bVth4fx7iGgekzBLUgFLW1NzZd3eNhyS7qBN5Mwc/6YLBWfusfST3rTCtUk/h9W3
Mk5igK+UqToab4dkvAJeaPrggSjNIoaJvNHwOsNQuS2MmVxPPIzaIcWxSpil4l9A
RhfpupKHI3CTADXm6iOwRFbdmsU26Hizncl20bvn6tP4eVk5QL2IvTBvTfkjMXsB
3gU9gB/Yi5d9jBF0ZNnDdowLGXFR2ERFuXMv2VjZEjWo8LM8M3n+v7pKeKIoFGA2
jszOD+9gdnf/pzI0J05qqQBTjrmDyI7MtwIMKff/MD+TKG0NFPftG6E9wydGXDf7
co9g/st7lrKOLkR3paYCVS2kHUm4o9HK0SBVxwl+aDmSG3zp2SVKO6Tjnsbkftu+
xrt9FEBqS6ElGornfoadeZST4DJ0DfBMKCZaVnUQwc5G2q3Fq/lQHXhAFUMbEdZS
b7pBop477yowsk/tcl46WRb50CUwPsmlbz5SJHc0twFfQdsTJCUZaY5MDSCRVTjo
AvuGGKPulzFzDvTuerWe5BMIyFyfUsNOmOe4bdc/4gez6empsX8rVGOymxWhY/Aa
f3YmJIqVQptuY02WaR8MNJ6oU0PuJmVUgOCH4JfZEToOxOh6a/TJP8ICzPa27NRf
NjwMt3gGE3sYzo3xLnfmCXmQgT/nTWy2TNpf/7xErnpUBbddXm/W2izL+cROE5cH
fDChBAFLAyoYz35nDsJQ3gkdVLsbfpJHyRvzSIoU7gzo9XARvNRjR039aMenyr3P
mXZKKWIX4Sl/u2YQ7iWBlkUEfO5U+1/rKXNYlejMMTH90g0mn7myMnP3Bwt3Laf+
CfxuP85tJBqVktrCwAWgDUezjxWjBagGH6nkwZPr3P75ip3iea6w8cNnogK1Qoon
tYg6wQZ/3dEC6mCxraONhvgxLJeWtez7PJUkchqk3JmTFz8sM704Shc5mbnz/BDm
kOjPBUn4jFKjo1Oz+Kk6FpEt763CpJgyOREN06TAVwgGUXMVlTYmCB4SwpqVxYds
Cqz93LiNHben06oNWt42sfBmNwImy/L09A34iDe/ly4STUVLXzgCsl27ErsiNRT3
5AyqVA5IleNX/jmBZAJlxByN5Dbx7F/QcaL5T/1CJu3GnvnW//+V4JRcCVMWSMU0
pGIgLFX6iVFsgdMSjLlSuqSMRta/gbaDgPhSrNjurRVrSzuFLX8Wu6O7/gq8JtIZ
pwKR5C/nH+9vtaHWQk300wQBkxvfkau6n7ta/EFgjPkUTKE+gVGLbyAddIja/H1t
3B+hh5I4OVUf6QVL65ruzUgx/UotzO94T6X+oItY8RO0u7379Qnqo20NnQGwgTsr
1ivks0kLROE9BhlGuAGtTRXCRezeJhZEi/DmnwVVixgY5Hzm3HTv6oBSMRtYCFCt
DerWa2aREQh6YKlPXABokWXE0oz6ZwZAvz02PknAQyZMCguIbEUqIfeuSAykm1qA
y3RTGzFS4cyg5HmTWmL8mhZtd1PuHaOCwRZjULw4J1C6PXJZ8GwyQQjpb4EZxFDD
354zDmIRFFjIHVLJpHNxCeLqso0AnvDIwUz+87qY2hOjWYtJDDVutvRoB9zgenm2
k8sOrSvWOO0pARcNZgPvrGzxeSsmjcDVYFIER2r901Gq15kAKG7xYUlUrxlFg92d
4AkYOseUUZ0Q9CX8JLXmbYE9v5zKgfpRvPdat4rPzzr71oXlx9Xzis+NYkf2cIH1
6uhT0GG4Ocb6mDSLdP0pvPUuqcfFe79UXDwT+AzueMnyVYbfzTLGtePddJqwdPwr
+b3YAfXrcUPP+JAcUReKZE0z1WGbF4fqr3I8Q94GWRIUsAawpokI5/JPfxQ3PfW8
Iaai1ok6JziInRQyoOzwZEhCVZoymA4geljEvpqnmzyZAAwfzMw2g+CS11HolDpy
4+M9T7GWSagbKAeCmMAgkhBQmudEUSh/PqPsiBXYVzeOQAWTR3ErnpsrCMEPOBQ0
JyQCviDwxnhqpjzfaF52yKviJOQoEoYB+w7pI3uEZSsZR0v/LPXxuuNuiPJk/v+U
RpL0fzNiE2eAdRHfK03idX/ZYhpaCusTejs0WSLadp79+dp3s5X3LTuZpPy5/qhK
TRpGjIez2G8dh2IkEIPKlXD/4g6wbpIjMRyfHGAGmcpBFh9pj90AzSvAPZgdpaNm
cQ5UtAXJeMv/+zyl2Q8Ov71+w25ba1e4tpUmDQxE/BTRzWIbRXuLaL3I4BoBUDh9
puNgyRQEppgXlL9sdAuZQw7JvoO2PCvuoUogsBckSLnDehUYL2/awpOmDrN+2wFv
ArOoGIxy5fqzfaOSGOvOr/hC4LKrcU+rmImIna706iiH6LVj4QIx+ImpuE/7LuYY
GJ5yMZ0ZEJO7x1HtiNNpw/i+L28nV202sM1PddeVt5YyIInYhXF4FL5/AoEGxklX
gKbBxWFZTdiSDCFCK7gO0LqFMMfBrLT+B9ZJMByIKK9Z9C6ziuBxo74I2BI+k2+c
xymSonQhdWOkcse0+9St26ZwhX0COM33r1/7hlLL/93+BOPsxMBR69zFM1PCinNn
sIUphTtfQQxxJS+wcf/9Noo6yxSGu9NG1Foej67HJ+4/+2TLUDNZc1QQiUSSq+u9
5jBl/Sz3d4VymvW4dpY7gIIFAPtdjeirEcNFbUtUiuImkeEpJf9EVBZKlSnNkMfI
gOFf2ixmttKM4b0p1hstbGgAHTHNo2f6TvxTUGyra/Bf7HRpXlj02XhusDFEgB1z
kxTsyo4jlIrDfiC1RglWZzNmPjAyNT8V3SZsAds0goqogYXXLRhTcqyA7a+QhmHC
psgMqsGQf2AdB2a1OR0MBrO2zxwqVrXYGTnXJfZCDs9FIzoRx0qkN9yFHNjxR4NA
eRyQH8UXcBEa2RfIxrikhfzYwz9BG4HxwRP1Dp9BIdsb473e6yOwSWdbUszEs8Uf
LDRrzWOQtN4WS0FUkq7j4kA92X1wggtm6YaWaMoiigcK1+M8/nnEuH9dkvUSLOXl
yv95Vudpo1arw5Xou1FWSVrjuo3KbQGgNFQqWchIqoc1uGLTySW1EaxR0hojBQn6
OVuYxG/jkn3pMy+JMVo8OPlVTcomcYTCq0jeI7qzAGe8fHXXiN9PLKbXS/Y2V3/N
qipEL/Qh1UiLHO8H4Rubq+JR3sWxovqMAXG77iLqaVuwOuBM+oD1EwGlwqulyMUv
IH73Ja6CxdGA5+g5Nqz7cF1ow8PNlTYYTWOu5X902A/Mq5ImocwIMgFASC30O/ju
CNvTCtRs838B06MWvBJoTcs0kSVCTLB5BF/FK6/IEuLQmdctCDcrxBOBMbFkySEZ
/1HvuMiIMMMnviyzKQyEs2zNhWXLxqttE13vovRyDXBx3pgTTgUafHD+7vdbAI2g
AqCO6uwhExqRVWOgVMIFMHi2PV0W1TRFIbhhAG2po/941zykrK74GInUM2MnquKp
9LcUptD3iaWZ8ShjRTcodNPDkcBEaJENJiPEeTYAmn+9TdpPXVyeCYZdPHOqm3RQ
EzY8wsmRaF2FdByLi/3CYt/ErtsbHUyd1sRHNG+MkNm6ewSSyWBmFB4JT6Ptmk5e
jBbePdMO+NW5wPeMV+mGNlOV9UIEOri2ukyq80v762fEcqrE/1XtpsWPiiepfjFa
V288CiCm90oJrDEzDfwb+AgtI+16Dk3AzPndymHy0px1dwPc9SNeh5z+OV62hDyB
7WlyN3VDjkUqP2s0YRR7zPc3OyZ7gTfiIp94QuWgVTqZguOSRKzatDmmXIFf/4Yr
VgGuCo+DdohsVDsEGvFpZbtlAx7yCwX0kVJROV6jY872y+L7c22XZPuwJUeq4Zf0
1rz0vq14wLlpNTNuDBQJuIK66RzDBJJqan+syRHiZBgIDSD97sDoI1wFj25na5mA
WzTk5Vm1Pz2WeX3icyfbwlxM2aId+n/ns9xECt1GbZkv0eO1iudNZzzuVPVrlT4/
LCpkXsE8KdTvzlQ3CZkc5V7LuGBJj3DLRxl3INc8T9Zvxs9w5e0ijC05HcaetaCp
u2J3fDpuvkrdiLE3NBsDsaBz50EajManxtO1jpn1Oy/qltNtABcUCbL0Di1z1y9I
2o0RnZEOIVuKSDdQaOL1+aIKc/tKVkbCjhQpBSgyI5Q6LKNK8AL7UEpSW3Qcgo4p
WkN/DU3NpKhSC9PmqychsgFYSzY6qfys6EeJfK27Vc29g+nhIO2AGVwhs5J6l/KT
B0AVkCeJFBW95JIJQlOaDCaiZb4/e6yZH1KMJIkZt750nxKzZ7UaWZoQ+vWGvDup
1hP583CaL3Fgi5/6+UhqTabIztVwWcSKii1MUzmd15KnZWbdraCu3n85iELb4KCT
OyeO9sRw8BO/Y+EEgCB/IC4QQ/rm1oQ4nrIGVASjrxjnBJmeZSMcdf1HbSUJeWsF
6jejDSVNVgtgL/beZ1fitWs8LW9KUSEIXsNUtAaM7/ZKw1CpqFft1OK+5ctVqflt
nZ+gyBU27pAqVoZNsJnprS6wLyOmGDJyvRNcvu6ZGWLp9v2vPtMbIgvq0s9FB1tO
6Cu5UA5cC/1xSUTjSwsxrsPvz6SUk0i3CRVcTxlEM4XyJDMqP/0dfoX6DxxRLKH5
oh4gDX14ndEOOThvtn7LQRVmUIoNyf9Y7zzPIEGevoVUT9cabMJZvqZpb2jbSqwO
pP24dzNTt4VfRCls5QA8X6rkrcjdqNoxZsowzs5zO5Umv1araLQWlaDYC+w1nTJ7
h3+klnaQw9ruUqNB2WltC77xry3MS7psp3d0OuyR68vHIvQsLZ6WyHhAXttNn4+8
GfEKVeAOuWB6C7JTgr4vXfn/FBhRxvYchld0j60RLYga+nY92FhMKpJY3tzIq5Oh
mPM7zYHSKkI1OcDvcowgYGo/HkYyxBNqUcC2vJYcMZisVcQLp0kB0TZ3sQ6tFkVF
OPKIerJ6HdxSEpr82qn/0dMA91SquuVVMt8wRKkvo8+G3/wd+CtfXPe1bBokJw5z
uRq63IBTxd4OrfQ+NWqV6cpiWetnt5HicPMCgm675vJ7Re98eU4L1plA9GWdXo0v
cA9Gvzw1SeZvfr1Y4oiLKLBHitPr7gbC+dAuyCMS5xjI6fCvzVKg/QCFvdV9NSTT
7rvmXU67KguCeE/IUgm2mWfF2jDhFgFeUM+s9VqGzlT1plshzV/dVQFh2RhwPeH5
/gn1mjCr3mQN2pjLSzmkMVg662H78DLLDxuyruFVsERhw50cq5A0MGEhn1QFJxqj
PG36uqafKb2OiiwqHymLtjvWcpuURkYpVlsUXL4WL/q8YelGh23BicJbn1dODTwr
aibm7U256bK6A4t/9AdKpBU+UQNirj8GYXUKbFThD2Nw5M/yCTU5S1JPoOAAKfIQ
rEYUjSIQXAidiuGjkIfh/VJ53LolnkPlQz4FqScrwy997udOLI6wLrCd3Apv+qRB
s4KWkfc/ngXLGxaQfzOKVvAuNM+B6UFEl8A9kv8BGzEr23LYbcYDmejkPAiR99XH
+pW6sny3tXbUB3aDxyoZ4jImBsISN8Gh01ZTI1ADnkBVQ56k5wppghDlXSeoe5PQ
EwRHs0aUiISEhCe2tEazsJZMk1N2updaDITrVYC+rkn1hn5pcoyOYsVT2lhztZIs
AzOBtlS+9Z91xaM/Ldz4eP/bq2wq3QKYSCiKjLKvnIaRSSjCkYYNokqdmRDWlywa
9NsA2Fs9u1iVYZyp97VPyptBsOylDx5WZIOdN0gYRVllSkdfKC05XdrhSbThumy+
ogn/0oia598cINYewbiD+Zs6B+3Fjx3/hJNyEhsR6TB3sZDgien0HgrF+ms5Uwer
R5pF+GqJjDhuHSnY0V7oWwhGV+xzMsIWMB2FK1ijSCwNE0KXfS9YZp554ciSS/av
FygoRb6TH5obSi4euMf4pM8EuGySD0acyLZMFtZW92hMvvitFgKqGOcL3EWTRiJK
LqUxkkikqSFCf7lMiDKkKXDHRmCdx4MBsN3YKWtF27ceCkU9kK5M9xLLB2JMqHHE
DXdAmjAgwzjQC77GOaoIlwQ7QQxxvppc7XM9NujsYgcCuZ9UOr2tUygR5UX2oM6A
TnFF8hKD5dBK0paA5GH9pdEK91JMAoqXvLIFBWMkwvfZ8ku0zR7/vv4O5SWnoCuZ
iJN6htLLltvmi0bmDnfrk3KH9grNKkIyiXVwWzUVEozNrH6L7BOmGT+zSCLav4mf
C2jNuKW/Lxe8yBINJVf9tg6nn5Q7RNNGiHNjsqBJISl8G0ahRv0j9O6SNHvCWQmT
4hdGdp2ikd2NLf41BqCkztF7IFXd2A2UmZMdbKQeKkf1JyX5M/ztt2S7wdHPLbIR
WsPkAQpqstY9ZawUTBh1K6rZIWhKrQbv6qHPiLQlb20ABhMQiXIkNYWxL1iDkvMq
IRHT7pn5oevEZHBDx6SW1dUCYrGJaede8VUpRMjeAsJAEgtt2sWYiUfCmioscQs2
mrrLUi00oqb8Bs4MXntY3eT++a5gSPQtKjvJllBlnCdjEIGZGRUzLYzAXX/q48qm
TEZ/hqX48yfI2yL4X+hgZVOUdKH8BpSF1/fECxOgRvV3ywIW/kEXY6Co38xorezA
PDp/k9swms8NSxb3hra7jyU3sf0GI3xU3w938t6jGt+iK849pZiYwRbJJ2Ea3jmW
6Wvfwf59O67dcRmO8yVINth+CikRj93keJUoUX5Wr0T3RqRv3ysI5sLiu73vOi31
xnmsbLukrdGUVOsk/4jp762kkEV1PE2LX7WFY40PRduisgEmTB5Aaxq4M3guF3IP
/7VgjCiPt1mBjAu840XvvIdXGjr3yMNIuaDpw5QpFwTDfbsjk+A02rLak4Ez4Ug1
YsO0S3MEZmL23SnQWRlJ8+N2DAKydnLYNXQKiyuv1snv9RJ7NutYLc5P/EFr5rsi
UeewUJmHWpeuD/j9OBZhhR4ex3Ln7CDsx6Dwt0WvP//MOl2TMbnAG7X2kSSS9O3r
AzwLlALlxfd6X7m8UQKg8plHd5IZgJ4+q0t84vVErRRtfhkqOa73apBmoyFw+8hx
W4cfKK/66MEkNxigVchgJJ8G3fFs2mkR+I0Ij1VK1hZyPysULGieuIDfreegfvX8
DrdiqFbxor1FHe7vGnPng2w7yG5HzbNa0KaiuqMHKKW7Z7SrSSI1KSuik1EuGeg4
Iq2ynJoQVxiUUA72HJWh8aJUzJ5790EhjoxtAFIuTBHQ43lLukT9QjT/dLBuLMPL
d0hr0wB8VufONzWFQQGk5eYP2igEE3g5s+4DdKpc4Pmv+2DvbuxOT4Yd9mMyF451
XhSXMWjD20bBc/5NY4mrNXOLwA/p8Hou4I46LnLwODdmergehVTUu7nIBYQ1P2dL
8Pojd8LrzgPxDxPVqol7i+wNaGJvBr4TVyhDmV2qL7uAha2RrDmmZO2atjMf4ej5
E537IKissSzGCbS1dwTuTEORXAXCTQx9YTWQ3LysviATHlabHt7noinOetnNfLgX
UQqjQnIaBofPQzlDMwoEJDZVQqhTDMJ2bi7oFtNsowhLWfbMU/tqdDBkQMnfts1e
dRIN7orMv/8vL3yMZMa0o8sp2QOTHL9g8NRMFF6f/2M7PoLyBBdJgolQMvfLqbIC
VPYepu2S7t8SlGp7eKjCRHtywcjWmUIrKeDC0vKtQPZRcHVTXKMlZ1CmM/ohCXEg
GetR2laUpOokAVHB/82vQWDqCN9gmL3nJXiyg43duoAdOip0No8rxkej6cvcsS2S
o9GwhzM8TPONkA3POlqkchXzSgqsSCwB4MTc51TN9VixXnNwerZZdpczpiutvd8B
Cb0U9/efekJD39AmW6ZSyXhURN9Kq3STklE1atf06UpvgjzHVqjV0ul5yqp9Ukyd
YGa25zyALyUE01p7wmFOQsPtPyfyxvnhRmRdK/jLT2pFYUm9CWzF7BFyUDVovk4o
ZXi6DI2SJaVelTxQl0D7IBm6grOguX7GVXxpzps1vispRPfjphDo2lL7F8Q8OyBR
ZEK+8iDBQRC4x+lJl5rUjCKqIeMimDdV9TJzgdsJH7w+zXCUkP01A94h/cZT0GgO
BPUhhaQSHt0W5HC7lFG80jYtZY0K3DF0iTzEVjJqKaOMfDx154L6vzD9xJmB9Dne
k00MZwYuHn1au2P1ZM/PPFT/GlYUq80WBrs2Nlrn2k0M+GaKVWFbP6KEMDs2rI67
C0wSyzkyj5fR0oa5Zj4M+gnJ1m5TQY2Y0mnJ4r2cTibPCqNDcYObs3PVIHZUEsUJ
6xawfdjbTeF9qXkdOrw2ehkLYDDFJk8VxSJ0k52kY9fRi3jciEkPwkyGPXYE80/p
NiRORnVB0FhHD1d54+EbW7yw9xdxfz4ShhgRGuuhYFmEXKImFBeGF3doTeLYj3Of
7oE0Nobr2c2aOo3Tq8d1o2se4UnkardLh6+1qutRjajwfbLxM/+GTXU0Oxc97IMO
nCocXDq9ZnmC1DIw0RYiuL03nVNEvMm6h8L8DOO3Z+mhLdpIZF1n6jjT/G+ScodH
SWTzsF/3NfYgCjKX7eZE6oVcXyhiFRKHtlZF+TEbifC7I3/Mxjrf9yvQVQ3che2y
M/55Y7KpzVowLVmcdEprThimtrF4Bq8WkU1D74LDBaRrJrbXpD+KnONTt9p2Sw5S
h/XBLSixDrMlbfyDgQu8w1aG1ykFpZRjo6w/BhPv4nDZWWRiwZqDaCD0GaDky0Z0
Q+iokbBK16jm8vPHpU5ZfBKr62n0sb8zkOefYgWlxnrEmfYNbJZAeUgReLOpZgwk
WU3lstVL+8J1kHGhpd6QNfHUIsqCNy2W6Mn266KjxeiqXwV4xc1Grl0xcorUj0n5
B+3PtWJl6AFe3PEimgxH5U7jHHYYxAz5E6kpgO+i+R5eIFS5kB8IE5p/DSmQRIBB
kgEac1b3lifDr240V/4nqX9dGzYt2NVQIhdVIB7/SJzg9PSottd4FyRJfHpY5U43
KkQZ1d3jMVFDmh9oBK1nMu2CzyyIJA3AtrNYg1w+4IEGZ/7vz3zltGCOqadx+NEh
ctoDzW+qVY9wy+Hkfk7HaV0foN3P7CwzIsXdMlnW53CkDCT7AOPTdEiJwY6Z+Ses
v/iH7A6VF4KYWU93c/a76XZLIQN0GIowxu7tzd/Yj4Xwa6NmR5Dwfw8qEPb1ThY6
AY9fv2lWoJXT/Jd21dKukg/5kl1s32rjKVM1Y1VUGgR/3kmEoQvZ/fQBMkJ/n/UF
u5SH0yLP6B2be9foKpkJBsOke4BCF8ARKa7CMIhx35vJwN9UTkTka8wDCq04AO+j
bjH05MdWww87KX0Rrn6X2DEAQ96kG3im8AJLWXt3ZspPZ+OKflOfjNKWZM0bmP36
KtFhLaOD+I+ROjxtPV5+Ppyba+zE5B1daV43fH7fPQzb2c0kPW5gyC49SQU3uCEI
jz0ZPE5B3ijjp8UlSBuIry0Y28NagguMNNxZL+PNuO7cTMcEMnseQwHcTdCLm5jc
NP2gDswb7u1XDzQ0OdT5Jlf0ns+ZUxXWbVB+3Ul3Q17eVtVYBodPqVipZYucGetm
EILwrfzMqPKcU/kLzBLNmE3wKQqQIAaTvbuNI+XXcQRFMHTpjRcys6HCsKGsdB3X
tjkgYKRu8eJnVFjYM9HuXeIIVq9/KC9wP3pw4Pt4+aDIznm0UhGqHjJfmKH0Smjp
0vo7itqU5KsLKqUV/16lTrtRJolcSh2wEjnrnKy0QPO4oD3XZamMBoIPNKmtMOKg
5knthK8kMYRfPielYRVv6JmOCJI7WQUShHkQRpSYZGguRLEawQKlqQuhj0D+wyfd
eghwHNBEg35UBlzCxLSmQ2llGXFAQLkYhlChisOP1y8fl4hOE1BDKpMhi3D7Lbwf
MO2t2UPlu/VQwrh+247sHbhD8WydkBCtnHCSk86wFgxPjQik/Ow55sxv4A+irD+F
7pnhVkDFCmHcnNe5G4Ihp1S5VaAcBuplWEKDQGjK4Dyn52G1OVYjMoe/0Nj5gPr/
q1atja7vCbGiZrPR/aJpRNlfJOMQuHxeQ4NCeTkfJ07+/MldAQLDne+zuSRfaR+4
TbR0u2ZL319EmWtF1URdg/BUtzcxF5Ti9Yht8yOzRupinXrf+TuiaN/rOsl1cK5f
T9DnwMORYisZUF/4ju6D3xNkJ1dBZBytSJ4kwzLDmoILD2oZ9cWgwtOnRkLAxPT0
7KxEWvTZmU+an6weEN6WlAXwjMo022ffjnO+kM2yF/TRiICebNruW7Ai1raTTJ8D
TL4+Gee6nqwEtIe+LmQrd56O17k5RSwapJ8sN6t0/ul/8B4YQ9S8H5Dt1et/HUDu
KJ7tyreZ5UuDUetPwizi+fmwBa6f+oe/vSOuhgWgrQ1taBkHqOpMLqvNHIyfVO59
4XNHmeXXIBeXdwXzaac/a1j5AhUvehZR0oFaT5mPrW/F4AhNaEF7FFO/HXPq9rEq
DBSlOm4IwtxUU1Gl6y0FyPhS3lEuu8yVCfGATDqz5qSmkS7MeMZF8CIBTjwgIPYN
Ls/l1yCW01euVLrwIOYhusr3XMI6hdcwDevcOUOYlGCB3tKNpaS61akMA1srwxc7
VzEy37QgPxcwqCj5CBXsTckU+VkrZGT+4ka7Uetzu5uIp6p/i5uGu/IjNcAoxP6W
cXcea5AUS/W8d4rENo8DNRy4JG6xybttVEAM9pDtUeL+bIVgeQqNjmOMoE9xrCQF
Jm9d90q4MHXPVelUaI+HbuNN4698YrxoFTH57YEp6txBwMvFDG68q8J2SlaZsC6A
QnXI04pQn4t7fOkXi2VT3zGIM0koF2cu5bOrjb/ptWs9hyF7RG+gtdXpgFVNZA6/
av+xgAsf67N33W76SH0AhuQZBllr18nN2WuryIE1CApx5rjnCBdv+gZZq8gTneN8
Goi+hCddb2lu6iEA8oPsPO9L2kWrmKbhuS5WkaAUhjFs/uYLXETP72JKiAz+VdHE
PpQ9eGHFtulPeKnZ/wMtQKg5WkONW+JTKNPGT6/YIt9gHLpi54uY+UkcVjHQjdtn
40O+UP2phKJO8jtnSiSIVBL60BaclcErDgkEMHUskDntTcv8C140h6R5WwAuvlRp
3MczP9Ct6CeaKe9l/tW5+ooq9hiFXUQcyPz+fMIXq+Grlg5ehRw1idbNS1LGaWzh
J1nfFR7uyyXxB/EEoTOD+gHa5SS0hDMP8KUopYJIP271RVcRx0avfMfpE0A0+qk3
/jT+D8a5DRk3V6sfSoCHq4wEep4lMAF3NKCndV91Kt0i9Lfob0fCoL993f26dkVh
EPiCvaAJO6n45ztyuMTx8emWLlPt4JmUzZDF8ocbUHFP0sjy2m/AqgHq6gKy30/Q
Ej4h/atgiu8OChzeyRYQYV2iZ9kDBrLQGkKxjyj99m7g0gQ3SM2MfFKtag1hZb/W
nBeMOwJXHR9QyCMX7sAcCiepGVmEtM2jWoQqRFa2iNGAgrkQu2grY0F0fRPdjahm
Olnx9kiRNkHK/iuIV4GWbQifLHMFTH+v/0K2Yrdrs4fgF5iHUzhPypF005HXBUcJ
DvizCNjSebFpCqrZvNjNxofGey+B81cCLpWWHGHL6zSI2xXr+5aSvNdL8d6MthJZ
86eh4fNZet1Z+QjLmVp38VSdzixKcTx8QrHND+6zfKHlDFhDKgnOnBc7jVq4YhAW
oGpkhDJjsQ86I13jI/HongccuZf57f/E+H6ZegbokbboVCkeAIqh8/vLGnXuD+Me
a51kLBwyl50sDQozLEOHGNr+Bi24PYVQ5A01xSdyukWudUe9OWUlkuXxXI+ZALJ5
PsHAFgnH1eXpT9q6faLyHvF25TND96aQ4bsTDNtF884qmOxiD5EIcj32y4Odb9F2
iUwRsN4xfIbFCKQcLhgYvE9Rl+icXElT6QkmYoFnzoRFb72vig7eX4Ljc39Q9Re2
pRwCoI9Cuc8u/3cDrQSmHslxGACx4Ol16xBQtfD3Eu2eXeI4QkSqXGijwr1vJfMc
Dp8x2JuVbAPJOdFyD0DLfnpeeTBQZ1eyJQvstW3AaHC2KQN24qH2h6+uV22w7LBF
fRs5XJMnSIff6+YQnjD5X0lzehgTMpuCoi4VRNRCclvwaOsQxqAazMZpQW0wJkKu
x0koqwWUJeVn9AOWd4QHtDbAtcPQ8G7xHhEKN+NvRu3SS+0GqUY+YDkAxgB1yu+r
ppdCPGTMfpoIj+fO5+4hqYREA+IvKlPhKcgP7scuC4Bi3iPfH7Z4LYTNnF/w5xv4
2x61LNheqyIwfMd8ewXekAswfCV+P486EsYy2Sw0BwmZnaKLjdEn/FZYUxgu4hp4
bWNbCDVPgd27nsL9/N1A26usOVwfEDoISjGgHB9qvFmdKxuzBGLNrwc2OatvD62n
Qb7TN/qkJILKYMwnTEFoBk9i0XWnuxN9JfnpEReTS70xt/e8jeFrBDYUBPhIWlYG
136cF/QVT8wcppoBuLZAqDQets2orEmrQRZHx8ATKTI/R4gL+yS1nKTtN/Eu01QL
8cl5f3Fmd3Ys7VE6S5pHY1vejn6dEIfDwZn9WIFndvILhMr0yJx6cpLUdUeyo1hr
d4b5aEsWeUtkOyY7NR5s1sL0ifQ0HyLH193HxgGs0q7YqmMpNUA8ZxsT+GIKkYar
I39r38kDteOPZUULwP4DlHQDWtY53TYO6LWULv/HroqtOkV8KQ8XV9YMIqfYNj5d
BQUYuWQ/ttqvSa+polAUVBzAQW76lv7Le2VkBjKud/R8LSr7loOLKt0chC6o3hvi
MVtnCka80pVOrXqhHCT45pWk8OMP7W3hqPHjaPCLS78J8GhpN9U0HVQRcq4lISI1
el5EiAShfgJLOLD3cqKaObICLf+D7pI26kjVS4fi6oI2y4JX1y/XcXkDwxBBNwwn
q2FGU1vfFTdWiu3IeY90dkpIHEFbdI6bm6l2lWugavHP8s2QYIy0DBvOkptvAlI1
E9QfWVq4b8G1VWmdyd+aA7Lww+dMVgFf/obvG65+r4qslTzeinFunl2a8B9xEBpF
5gM01PM6gIlV4ct9dUmPyBDDZQFWRbQR4SSFmimHAl0vW4bxNG91wl76aLJInVnq
21jENw9TEdhHZNZfNUklrba8diQJ5wCCywnWzgVa1XI1lU0jF+gir/DUQFywF6mf
nExEUhFCGy6qo8VCCkYaG3vWNkT8Qk7jVhyJYxXzu18U0BSz6/rT2wcML9/J4oVK
6tbdWGXhCjTKulttL1L8WrdDgNT2iYsPfWLF0vGzoxeAakxOPubr6lJsUAbS1LID
tiKZx4zS1R6X5ccqtXDlNRurZt/OyV2YKVdIL/0toErxlcGiuottGLAOsBRVgORU
p1pH3PNkXwbJTGF+h0TSMyvvHDMnN/2wyojTuYBYd2jQjhA4ffjMRRfSYll13q/g
BAPnZCSkrVR2ZFTobzCTGcXRxQbgXkD+dzupXhoReCcNEyuqMyrFSHC6A1rjfXDm
tyO/AyepdP6Lx8We0K18c2b4zhzMaJvgxoWz771IQT0/ixqa1bc+HNka5V1hQy2n
EflDGJLkqg99WrZmWnepk12VDKgHrBmul7UmbgzMcYlgDuWbQSh57ZXVIk+U4/5y
OdsbbYb1YvTH0AP68IHRnEFlBRcdch+WY4FPR/VxL3hnE4uocQHk6eo41qGuRY8o
uQsB6OWz5Jzug7cvzSD7TRBvHIBuLR/pLPCBs3uK2eTN5skEXNVORahdYUZCEEkB
gTLLooSpgjaAgYfYMPx6hi2h64Oa/8JNkW4ijiwtV1jZMsjJ9WEkYt2r99mSIHmx
FJWVWuKzFYS3PW1iStrA/ffFezahAbHhmpi9dnK4jFcs93rT8OzFc8MS+WT53/eR
7+chOJl8QOCCyFSm9bevGFXJduzcI5QzH8O42ohzkBkHLeUwVH3ahQ59PtE5fg0K
Amu7e/72BWW/cuS7xFcFix7d6u3kddyyn2/HpR9UD7wtO2TbQk241tDdbNmiHl7m
S9AOxh2OFJKcMUoWYHd+h7f6KEKKpIB7eMc2BvsSTgc80yhIM/3N+KG+WwEelOCt
MPf0vNt4I+onKXNoSXbPr0AhOPdiW/cht1XlKWDtgOtvykw4Fi0Xzif/f4Ck8yqT
MIKLB3MO/5H7nwFss4pmZZBdo5fcPN5TAJCJMWdze8G8hR8b8LNRGHEiMGH5lJLG
sb5WFwb3wdGYBTNfhWfMUYEwj4O0h8OiiGf1W48HEKP2trlDizWzXFlHOlNCTTjv
BTEAPr7u4XwU2WbjpLmv7wS/Ix7BuzCc08rTY+C2Cx4Zk/1occVDWhiZbSOmgMb2
VUx9Cqawrcrxb9bRTI8lSkWGB+bWRPjUudjcz4dDWMnAhyec7i5L8/lkxsGpYBn8
QrQzdwCwBNHPJgp80Lqpkl4ncPGp1Ul9rUqZCsdH8uiDEPzjEIHA1vy0VgBd5f5b
hAOuadn2gmQhg0so4AUI80QDuPUk6YLzh4c1zd0bd8GceAgUN8YCnTlW0zqUnOUh
dCSlJ4ZPIEUMl23RXXqaQCOHhIpT2v801zmH9qAooHcQypig1uSCykf4GBEIod23
vLeseMyvNvkLv8CZ+5dXst9ImH0Jmogug+TihyZZRtRB9fBYNu1HO0X8jSbakDlR
TjGv8DFkeqX5m0ucrI+pTJcMBYTEshJNGm+LHianm86lXdQczElhj2VnTR4UXHL7
QpwRgBFxlvftNqCsigaflSI9Mnhs3Q4BmT4DAefRmHlpg4C5kNdWqTr9XEGpIfVN
JVBaYlmDh3Q2qaC+KqHe5z/u4nlwULspdJkQvn0LgDAKOht07IFAT5O19mgXwJsB
UIzNPLZqtI2nhcdoIowzYYhlxgwRnXcJVMzjW7TrdOh8Ht3Cw+drdd0OpE0s+SeE
DihRmgT6bNMWwKKEDyjyA9QfcBJfKjSZwydKui0kwEKWKdLkJyW+uIPW2EpzI4yn
0CqsJdfm8iqw6iFaAF3FpZKMoKU/OfzpvM+zYYUEvSt32JPWzSBf3qTGzzorHlz5
Y5rZkMO8laKXSTct6lK4hGm65uk5PIBfT9XulGBaUCPIDXHgPhxd5pGQtLI1fA63
iJX3fi/j83UoZcO/ZfxCdEnIz2g3Kx2oYE6YxFkBECK1Kfaw9gaRMY02PS1b3CtH
N01OeEuRMyJlRX9bVDXJ6TUq5eaObZVn27N7jaYFLWEBWv3GZ7e19IWRwkO6HrW4
6ApG7zopd52M+Ts37NiPrfK7wxcYQ1J8sMVY7e7zJeQKDR6JOoM5s1+NEPK6eZN6
YInhfXp5SYTRSF3RrMVd3h0NjCRy0vpVBIonOrbjgjTuEqhFtt6gV3NmVBjZtDYB
5t2P+1UEJAKMVDiQwiG/CNEJ2l2aIsaP1ZcmJrrsGrX/jid7cX263nC1QMs0BLEu
MLvpIE/P2ux10GVNnXl5wM+acmYOwVeQolrPe5+HbFcbhxWdxLjxe0dWY2bqJ7EX
Gh1eYP3rpWVaQ4FDNpxpw4KDuKYIakl1JAlylQf+XJpwulNGZeIQu05LU/0+Wunx
GSCeRIurmwSipOfYW3p4T4OtMjEfFTfIOFAv4ze9S/DMsehUlbBXS8Uq+J8sMC4C
tPWUI/BWzYUkoNjQ6lfFqzM75y/GBhYhwGHLaRjQDJBA6ShvyU5pZFkQtjLqZ8tB
XN7r7W/7Kdtwg90X3g9pTyuem7FGMnFqg/q64JU+J4+U95+orZEa5v7EiY+NIJ39
Z+y2XgyU2jIO4LNRNAC71ZKeC+fWOfcGo5/o3isEu7sVuLIsOqNIDwBkum28RmsE
Wp3iY4nB6HZwC0pnM/rDt8l9tWqWzVLfe+xXrFH8Zk1r+kT2VVdxzUo/Kzez+hx8
XWT7p5ORhAjE4rAaPikDR+z1eYPfekbB9iyXsqXGWWwFy2uL0JDzU6c8SH3F4+UU
UIkqxf06LCzEt6M4vXxBg9oEmDW8g60f4FJJyBLWrljzsXlWdcphs/AOc6OdkiQW
laPVsG7c49UmAX4DEuaDE9T0M4kQ1zqYL/n1FzcpGh65fqVq9q6mDmv8Cw1DUAaC
0xIYPevMNzDllEVvYaEy5HfYjHWLpsKLrG8JooJVncpC2ylHgAur96bFXlo9Ikim
Pe7DXJcVGBtVlYJoMQNNCpm5Eq32FYEdlhlRoaTw3FjwuwIvmfUaVIfsf9RFNRNW
vPkPkR4d/tuZxIXFZ27qqD1qYlmreFMiF4psNohIxeviB79OfU4fN6KhzasLW2G5
vlKJ4XAmFQJfxfYYhgu3jo3+1+cyQxT5HEUoP4XYqI6yluPKmIABZ0/fNUNf5Np9
2+u2q/iIUZwFj1E4B6zYtrmO3oQDZaEpt5VIUYWBAChuIEbO+x4ZW+Qil28gprE6
bQXsukuKNEuhyJdNRV5GTUFenqPob3SEcDsSbPSRvo65beDj9R5UTPX/psBApBbp
6ubKlAPSO0tYaMT5Q6IUyCJ0QlACMjBm9DAKtiowFcRuo0mP9Azbv79IJPol8J1N
iXQeEJf/XJWuI0KXZbhTnsbKgnspsillC6XWSRxOC4PV/iEnSuwFZdJRN7aNoItU
kvmrNnrVDZQzbck0d5WzQQph+HOE1P4MER85ZgzauFd0HDrYOayOE7CzyTh9fp5J
Awq1oeItsZVpNMK5h4xSVcqvV5MAbAYszyEFgo35j7whs/wFbZ4/n6pAg/OYOfsG
5m35ZG0/vVo4yaq7DabXkVibPEualvbXjJFAXJXtg1WRGAMTr/MI9S7hl0P43bWN
MLddGSWwxnfcxqiLiQCAMS5NgwCt9aHnc/qisR3CebTAxlNlNXtWwLy43Abn3hX0
jbp5E8LhU3CkrPOhq4RsrmYGLqdz5SjsF2scnYSt077oIKRJINI5SWL3RowhQ9Z9
Cd8Hglt13vLgHm6vvWrkTzwL5j7FWgWeFPd4JwyWme9gaZpn04EexBNW7KUPg6wK
dQtCeG/l85aRrdkxDDXYRclYZd6FsgkaHpNwEpp+trozM9U+sLct54oTFclsllpb
58rCNH7+gplK+aCRZiegu20tXCICGclNxlGL+KSpk3/yfCh11O+XJ72dJ5J0E5Fe
aZC3e/nJzlGxwzCAqAY1vesfLOL18WmQX8YBhN5zpTYGrbL8dvulRuuzen1Z6mLA
K37r2mZAObSSax7jodFXVHHR1Ve7m2KrdXFOEhEJwKkPsmPrlIehXb599PIT0TKl
zI8WotKonPVK78Jam+KCSVrcrnP3N4xsX6aq6pYZ+q8WMX9Pmy9wP1HWsodvJYtm
3vXKz7aXkcCNCGMvCP3RynPE2LQDLySM0vgkpMmpT6Z7Yw37D68gZwQ4/4GHGLxK
GPX+4PQnBV5f0DOKah8i3KLH9+AKOcTJan2Z6xlt2t8cOA8+RqEHA0jXgEahG2Sv
2wU0IZxbOkxjwdFltceSY6tBxIMVC6SEa7tjcUn5LjJvU9bgT1p4O11AIVuvWVpX
PE7IkF4/KU/NVLq9kTlEP+O+NSB0w9d6OTELcM3FQckdxG4Eu5rz7Zb+AtRkqOMC
F59mN1Lvq+nXtHTkWU1DCd/Ar2w9uvZlmefR2dQ5H+HqT9fysCMWO70EmQyFt0gb
0bvFh/Q/G+LQP4Vp8spIKGoXchqqeIPmSu64Ugb6hNI2e6bTGQkZDaa4hagDyW1Y
am3/c45nQNj17eB+jkQEfGa+W/4q9jEJ2hQGxnz6ddl0dDYLtPFrAbhbbSD2k+63
8/69LVo75oJkiVruN47+iHy20/bnEk8riJ15WWQrfUzXz8S/WWSm0Gx1bJbuVDmh
C7BgrsnvF+8CMGa3oB2HL5YjeeUWXHM7ZpRCAbkLkeZ2o/LtRUNc+o4lxu9YWc57
yasoiSRq3OW7cv+GwwY4xXPEkdARX7P69UbjWoj0h2W1akYkwxfRUBkTDTve3YER
9p5f9ZKq0L4SZvD/PBEWMkBHZzW+ACjg2msdvKlMhbUh6BEJS0WcmixJeCJdXEhO
1knS85GCYroGgLc4KNRYexUUqagqhtTXxNI7U154vVVVc3Fe2Ce8AGtNX7UYuurp
sRUsPOf7DWas345TtaN0X83VlzaeN9zansLSFDRCW7/7FEc9/0ZCSo5L2LxQ2OIp
y881nSdDF5jhVVu8cUfIXO+HMxl6FS9yKLGZVVhAeCFdWzMxl95PzWqeEhbg8lg+
qRPgY89h1x1NPyUleta4p3wuy3O48zu7th67kXyi/gLC5/bEoTi5BkMBuHACCxUq
Ge6hA0/32qEizYrokXpRuXrHIS+11tiGW6/hUKe+/KsFLtjcOOt7zPvBB2mNQI/j
FQIsJvdgAeVlknoE6gZXlejUcQUhswd81sLSdEssgXeqUIr97g3yv7zT50xmdpZS
UzQgagDJuJ9beYdhZGXX/reZ+3NtJNT4YzExVTZhJzMqU/QiNJsl//mUUYQmvn3e
r95qcgkQp1ZGtD82w+ybwxT/TdJ3vmY9nuRYIUITfSFUvquX1YaABnfOn0B0Rw2u
NPX/yuM0Ygs3A3H34QJZxRTISOFt8bLApEcj/cF0r3M9Gwe1InM8LyWVy3mb0ptt
IY7pjOLAQjVe37ePux2t76tIHQIosrMhMTxUSuctE7vpubbm7YlxSBOaEd7Qpef5
GGE2skRNwc3rmuCQ4H73QYBBsz5nJJIt0cS7/Yol2iKGNHwIsj5l48ZbV2tP7qbk
Y0j6d6egh23oeq/uwYiKY03LyW+loz6fMv+NwhYkGUQnAxG6Rnh23a9XlVnz/+Fo
IfnUXTWu/8qhU+COr8p1couXCCvDFJEKEw437of6c4iuzkmLgJ8lgQT0qWdWlqAa
/QxT+QO1jepWEgp2tlFpqIcdGPLWsC5JlAobgYqK2jdxYhQTpp8z7SSVVnKOfZTb
BW/GtRmbscpKDzfJv+hyi5XHlkLRKK6M2oQAqba3vYtF0rM3eUK5w0qdQMxNkvCb
cvME/HhKnozsboR1QgBIoq+DKFhFpNVFb+8N/hle26/VDFYsQc2c7ROHpTHeyv14
SuWBbm0aQgT3G4R6vzC2ZsMVswyK0i3StzpeKa4XcAOp7E5HSZny/Dfw86N+kHGf
VC6rQfH9CrDsv8tr5sH974DfnFRuHjdaGns3OiDuRkHLzNEd/H9kKlZCo1l3DqYM
iFLS2w5EQLYjQZp5gwhzxcOLLAlRYYFDten8DDaozBmtzxLa4rI3+XV7vEktfENa
SVhbY8U3YwsRWv/3x5ZIqZesiOdc8evY+FbSR47MM2KhQdLn7cvrqqeeo7GV/rPM
V9j+MwaWPZZN6Cjo9rWvrVoW8DCAcNJvb9eDksePcf1x7CX2kzTAAMVFrBX7f5VA
F+ybbX7BVCDAM7sCAD/y0JUJ05XvMrh4y5rHp4il2Lr1q9kGQ0CGgtxxG9YaZJgf
+e7vVVbflMXvKv6B9olhkK9E/WmrFW+yDzqJ/VS3w37iymRqVqhliCk35HcstHBO
o/ebhNEU0E93ALikgvylDiB+quDRvuSmCpuQEVAb2SRkrR4Vsgiz6JKZ72b96pNd
TuplZquYPpahb3YD/BgrC2sYMo2mH113kVPwSvJudbzPBONjYk8XrFb5cWNV6IqA
8VnqxshU5RPWnxvCRjWjHE4wwddmtsReZ//gJaoFE/vckSs8T/MyKpsXEH5brslj
4yFyWv+lJ0UOQ/pw/eK34nyvHlp+q4fvTfahJsOPEZS471XWlpaw6LLfEQilVBBo
nwZswI+EyrM6fmpG3t8GARqpiSsAxJiE2zK4KTGOGc5lltKpSAgapPnnn8WoSNA8
4ONrZZZetvng+CiKt6h+IL6pXiGOgrt2DieXNed5COlkRLb4gJ8+y75Iq+knMlEe
qiUfScSP5J/4rmAqW9uTjcDnC4ZFDHC65SyKKM329tHdVXxgIHQdXrOjUd1qvDeO
w3/Nb4koQDdloHDSA/M++bdwWDDy6Ihj0Cpa0yWi531dyJYqen+DwSWG5+rGsnyR
xEYmiQ1nG2/OQrQqC7VLIVAReTPav5dCYQ3DCD2oVpaYP8LIlW/mlBcuF3MdxCWW
HoSYKZ0qdWOELvyh/mfCfr35bYO1y9PnDgGAuIBR+RBXrbatLAIUdJR4AnZ9hikE
7tKkRkE6cOILAIYrxpgxZcU+rhv1FNiCZLmYYVu74v51nCPPH0hksQVpvpygpNvx
ccJRIsSKn5iHbdaRRt5TARJu/xCCXQ7t/O5qWG1+/7mwwkEPrCtpJsx06JXZM4tQ
NEd2onvUkbNDLF/5OX65P8/DabE6YKhuM+V/ar5SXDdzejaHh+St0G9n5Iqcqlk7
BrZ6CT24Vp9AqYGx8+8pCmcVSDDyJN+kzI8sgnd2vCw0DlM4RIJjEwCGQVmEx25M
qNxJASrGj3zdcp4sbrZ+bXXy36Wd+SIQasXDwMT0tMlXPyJLYRBdtdmXuOGiQpsI
k8KCcsdgcynfV/GDA6aZW+ucjk9tbZ5o8FaVcpIaRHGB71yo+UmMmryu+qhe50ai
rJcFYb8rkhgdI5Zf6SsnNu/cSM2TJNPvpsV5csIeBm5flDNe4ejSroiXdES7dqqG
4y/yZqIK/FipPBw/yoIQmhnEaI5h3CDT3yT2kx4kpdOfGDlIRToz7dWZRYDiMKUd
r0HRB2256nXqG+lt0ejqB2Wr3bAPo73cJkgBH45RHGoN9qTZcBN7q/L5LU+sDVp1
wXQqGAP14kLZrACvGHd0BDQqIw7Pp3j7HuF3vouMfp8o0CoVY3j1W/EOgbZwlHO4
3Fu9txDfhGa1N75JntCXHWvv3blSYMHp4gGQxHZn1UlfYhPgdBuCWpqWbtJPoxvl
N8hmsDyFlR17i9+zERIVMcqmkwoamdb/7/9otOzoOZpRCF5MB7OUfoMubIFYk4Tw
hZ2vz0aFv5FQ+/Aj3skRjWU6slKfEVaQmVgVhTNeU2gwIhnicreio9CfJwEqknaq
QDUL4GHT28TcgMLBJKePCj38Sn0wMLRuyUYD3kl3exy7dAng0YgB6ma66OzLdmiW
dZrNG3Ll3joWZIgKh37Jv4VbMVcSRobYctphf2eQY2K25v85lXiewDYT+CLaDTSe
TriAzAiptTByhTw5+UK+p/Qvs2WuVyd+K27AExh9YVBEjXza6CtIdaOpok9VftkZ
eL4AuS6oPf+998RlL6p5Oe/ioNl2Z5m3qcgLJrDx2Pj1JYCSSg/M7lJUkOBTCj1I
gpFBTeF040+M0/AAUlhk8yfKBaUOY9wfjyPj9pE2eGeja/Bt5PLaIQc+pFGl6wGk
vnZ5nDfgIFmZTg1yv35gs/H/gv7ICBz0gbqUqPWo08O5Dzrrqq0QpVfGHc1rnxbh
41gN8i2P9bQ51jYLjApGL1sqkskdVVWLUd01SDWqZbJfllXQvGQYRQDe6El28uEW
veMZYYjo3aiaBn0cq4JmYAiDC0/pr9OUQJRVxWpjjcvOLsRXQ7TKHgqFFIOL9vhj
WNDTj9V1zxu8hhN9qQohS2RoPNyk7bTAGSK/3mRDcBrQfKJAmy70E83AMokwSfOE
XzDG9NrW0w8SOKCW1jDcGsOtxOkFZQvwcsKEWevR12HRnQQcp28OfYx5B8Mz7N9y
sjhQOTM0OrcMG2N6dInY2Rh3TndHUjxktMo1i25dEbxzO28mJNtmvTzPUQXREZBt
XNddhBKHYDUchCZDStWRO8ir8eyLr2l/bBy/8n0MpzhYhSFP2ZaGuev3VjgqLyMr
SJcPx9swVeFl1/6zuSeVkjOJ82NPWE4J6wRqxL3fpzokEOwVLAXzEA36LEq24Dlq
k+VdhD+gw3i+9QmGoMDpMjA4i2OPcvmxl2nxPr0zlYs4mzlaF8uv5+WVUJBs6Vlj
WInvlo4rX4UKT8tOSM9pW5wXJQbxC0NMhly7wdj7ieN2QDkGMylGFDkqgv7pMRC4
/SSDJHQcN+supyHwVlrxhOyF6DMMi7dA05MFiOHT3TXcKgZLk3SP9MvHVUA2R7es
VSyrif0C6A2NsgmHxGFDJMLOzshMM715qcvxNuJjsIxOWUxop47+nPoMS6syE9nE
fclLnsaTl9BQSyUlZGFppjNrZv/JfbUKVHyQgrOYJmN38G1eK4wQ5cDvwKuqAe5o
xVC63qc1/f6G0osUd1VM4CiLq2klizgy6OTxqY04GdRq6bJIAkLPVNT9cihK2I9r
5QarfbpN6ZBqSOcI+WIW5sMTuPFn+d69ki6yr6pxtGrNVylNNP1QSNowxQkvi2e9
kB2wHpM+8F7eG+8IcvEK1ZDefD2kt/AABExWNYJ4MsdaUcGBP6SAVfSLXPXDw/hm
3Y6w0qdqPcvSjTIHf0LNydl3Iz8pWImxBEOjO22pWWQ1e+gO8dlK8gl8UJafbsOj
vjRdvHc2+NDdtG2Ak5zRtsijlLTN4hURZ+HopllS8I1ZSKaN6Odg+f7jRYrqPSVb
Eym3/bZHq//WwtldM1rhYwro7JVCLlkioaNxs9xDPbDj6aUpdKeU/Nd4psaJQD2Y
fSZuT9NMt1DaN8WFyjgh2y00Hu3r5YJsHxgDMSJQAHVzO69Cthoxv/agAfrENRrj
lZm8DIasDosGIA9O+kvjBRH+pAOj+sn3KKr9vX2Ep0CMRvg+FE3CFQuw7thvdPI1
itEcENgYohnX4L4bQakXE08k70P5LqyICQi1Wp3hH8fdUgLPEsmUV1nsF2IaxXoH
TY/kogblEbfnEjqRmc5PDV9AfOlWePn8+fxhKzjXrgU7JNVzFAd4diywB/Rk5wDD
AaFBC3KUa3MPLhhG7RzrVeuj5G3W0fnADCCh3Phh5seK/lAbLpC15v2LXFyXEPpQ
WnniC/lrizLpV9ClHhB3DG0/3ZrIYrplUvJSJTgFlCO7vuz3gkL180an/b2tkNqa
/gYIv9rWOgalB8e2NHPwrxev/Fpe83q2uH3OCtFVLEZfrBRsEvO/rBSSexVfqUVM
t5KI2OT4UQ9731w4ZhrZ2q1HkFgwXcyeVg1ZcZXkRezMkWYUKNuIQZmoitZ+IJa7
5nbZ4fiFn1LSylUiQKO/8BfdemcfltsTahttTD6meaLFooEpwDLLYHF1LfpfjxmH
C9cNtuzJZvDWWPeZMoRg/Xj4XqCXr5noi0G0oi2ae3nNEKxNpl0rbvkh9UHchYBh
lQAKjg91If0lPyMmy4vBwk8Av0STTDOKe4zIJn1WlrTWzBXq33rB8+8e3bw+WzVC
s1zxrutxj7Dq5TZXuXQD9Rir/i1BoSU5HowZvoGUMhEevS9l/LB1LiI+Jo2P8YTX
Af5u9q/iioJOuL74r9q/BPKTw3EBaILPOaERshabv0yJh7wXPPJ6WJFwBaP6bcPE
puXE5v/8hoqOHLJN/qeeA93aQdbR7xg/htO554J5OpbE4a8/MxSW0hbjFTTKijYn
agDjLDqsEXIRvKUOy87FiiXlLjun4vXcCsWIRbMSmHLXA000mGLZeGOkLcauqbMj
Gk6AaRZeLqjUQ8QAHDu9daVlc5T4zoWIxLq3vkZKWVYyJ6pLyePot/tnSq3ctY9d
s0QwQ3kr5J79aSIXAB/STgctZilBR04QfRBwUvtHwVr8YnL+vHlVE/eQ0ePBJp8p
gvRWedmoKZy4WT2de+hnrA8UWmlUMUqlfL73kUCsc29Ilb6OWOFoUBxugzlrLiTg
LKd3eWhrt2nZwnNFp6HC5U9uKJ2QgvjTjjxXqOcvAOPAmsrEgTJQhw3f6ruuA2VD
uDnkVUuLYIlvKi/lYslEMNS+hpKnD5m1MymviMflQeArtBKHcWS2gtXukzgytl2n
AnmVqOMpyDuYizPcXr1PZ0Q08lBIucvQDoe+HW01zjOzU2znjcrLi6ImGbZfcYtW
KziuXgAiS/vAXHcW1/JZjzC4orUQDFM4yz2rWCvsoBKCJLVfmJRjH+Gzobj0wptq
Rx9qKwSu2Y3UKExrL0MGhMkoyAVLUN4Rq2IAEAepZ+uLuJgllk2M0Vzff7bpPrjw
t4Jz8B7JV20/dSr1U7IUzgm1c8VaoJe1eIWR3+sf2n9Hu+o+Klv3FAHFJ+yuq4kn
rrUAum0tgpoBZZ+Wz/QFxSK8z1od/pkljWtSk75O3f4Y5Rk5O61sXWTsCQAsxdCw
4vaQiWEZ+aX7s/rV9CJML+9RkeYn9N9sHcmpusra7fnRxg6d9H45E6fmO3wX5/Ch
MELZ0bxxhrlMcUAyv6FkMKP8eU7gGcAf95L8M31eViPYU0LWKi2yvdelxXGb0iqn
2uy9plVmmHn51ZjoW+RgUvd843glbt1JZERPepFYD7wDyam4cM8WcH34LHOX6K3w
xcJWnJM11dGTx45NdrDE79OrTnpyKvx/SJbhaHFcvpmaZDLSiH07QRzOINE9ozms
5+RyL2WraezpHC/Q+7qrl4rPdth3M3KgeCYA083QLEUaOc27W3+3RhD35JAF+0n7
y7EnTR9k2vB7RfXvhH8zdgSgVa+uKe/MldMtmfbE7SdH3cuP4WxquupZ/w4nMwIn
NVUjxAJ+GRMpNrQmphlVn/+D6NPsCdpEOjCk7a2YUDaOeRehTF1TaggUFQWtkXJ2
tEXWKpxExxZqf+A59FIvRci65WzRpnqEOcNCRbRtPcG9f1c2+g54Hor7ITgWKPsV
xxAm09E0wmz+9U083+2p1GI7/UdHqSn7QFKp/dIrUhsZND4n7ec4QYUDntvHwa5Z
b7pt/ZV44+C1wm6UNEZFa6IZiUSf2USDGthrU5QASCSND666eLU/ItvUeh4v30En
pvBG2JSfmltMc1voc60tWnBsn6SFdl+szA5vQ6uYk5Zz2D0U6vJxuDRGMNjrGKdE
HdOh4A0PBTB4qGe6vct3QmgZiOokYxLgdifQ49bv3UO+KqTwRdKTk2Sn4tg29X0E
LFqhktw4/Vf0r5sMx1AsB9M2/lRyjHzxd2MUTjg8DRp/hxTkjkiF7ru8PzvGR9No
/zPYX8LWyVanYsz9gwCCuwdD0ZgmcFwRwXBiaT0QeIxif897J8lusdQwczR0ZfZ3
Q1NQ5KnKUYItrDjVm+MjNnXwzaqR5bi8kiUXg3jvo3R4O6xVIa6OOBZwowkurY5x
/K6OPQzRCEl47VnTdYtnK6l9OTLK9fmxoBYDe2aYvSzGHZTRGGONhU52GQCtNUSh
139HUEasx9uynA5oQOjJkH8FW2w2rpB2HmZ6u0BfcbaKbGqc0JX+6CtjIoxXyF2P
u9S2wNQmMADRQDY9E9kQPXzyh9xwJy351i6A29RlMvFogrQedfKvBLsIN0rtRPP9
J9bstWU7e0ttVIzzKD+POskDCCaC21rrV3inUuN5heBw6TpA2/d9FzWIaZS4fDwI
ifx3R10rssNHFuA6cbf1gWYnsrFhfX8xtt9OgKqEgMJWS6N8mr9TKK9m8SlRDNT0
T2en6apLD2xhNibvmR7mu9UKtOvFQSYjAURwXqxhyIIq90L+1eN/+ujo8co0EbM9
5gYhdm2I3eB99hOLkr9ZcQcjXThty1ui84MYVrv0e5kke4jv/zjg5qdF3o+NCTd5
3gD/mnnQA6V05PGI1ETLoW0/x9V7PiInz/HFb/2fd4g+U46mT4nmFqITRlcNLcjS
U5MfFSiNP2xl2fpC1a1ESOqNdxW9on+foDNwLyt9eRJhF1nnmSZ8dCtPcgdLXrB3
k/18LrcZdmENSwdjnLWidl0olaVB0bHFdjKXiUpKaS4GsMX59IretyBpx/TzuAeW
h8p3EXm4zNB/mInrV0UTRG3jvoBiuLP+kQdjT7YtqDXJKHDTrLBBFJqkcK2xsEjo
tdSBSDpvcIWuck4rCHzMSXSMjIz8KX+RoG6bCdHVPmeHQ5oEROs2UozXt7mEqgqj
vrPqxgmkWITH/1/QSg3frh0bHE09PlnsecAVLDSpk1UOsU9lvLwvLtkjP0yfg3mM
5jNCtL0yBfucwKJWQn3ksTPER+2rcEGnaHRFLr3quK7mrDZxrUg1q7ZZ40d73XhQ
M3ItE47EikEfJDMjP0Xz5mFRjhlBeE9KkouMp5cxTOTJQpMACJLvjegWW8QIFp5G
xrBviPMA+Xp93mXBYlXZIP44ChuLN3mZfv/TeaoA+t2VtSo8fPuwdqdWfo6mgcBf
T7XJOKWanzw1u0VTHZi95I8eh5h3xdhal1ZHBWAzc7Em18tjQkFuK8WhezjrDtyd
npyYNA6Tr2UA7/2aA23n/kmqTou1IM6XnUxDAHtK2tM03Oy1dEOoprEt3aML5C0G
oo0UdwlZk8rnrhzSKz8z7aIgqoMHukMFQiZ2XL6n+U+x/Mkxl+AFU2jj/ukCXczA
5uxTypHTGKBnlgl4fs684MuQSD/JkEzxI7nSSc3LR40rYw89MyLUvInkNhFAH7OF
bJCbmkcGWKhSmKveP+oaMdGaOWOSUfCtNE/9eV0pes1r/H8btrXfdz6/haGRO3fx
FMHbaYj8tDjMA5dYQTQJPqYeSrSiWkyvY4EmU5RwUPeNlAT+FO1H1A1sOJlFQ/IT
61pHbyQ/aWRG0YaCP228Tre2MoxZEPAAEIoHslieCqqLBpFPXauKzvMYHatYLhzx
FO2M32yjXFQYe0skIIIx8pRgiDCJfJV745c3/LahfA5AZ3syHl3+xTaRdCMsbGEX
S2cPx3mwqITbG9i+59AWZdJkmVAqInWNFJhlCVIBvD2kYrhPnvRGqN4BF1RTLRax
cpVnPuCLmebAjcVJjCVJMWVE9DtSdXsrEvRXeyJtOtMUKCW3V9iy2KnHqjBq3U1G
aiV6DMV++/mWmT1R2ccGalGxX4Np+iGoEfob7TfY1e1fw3c3wA37AY/h4Ink+gI4
hk2TG8dmG/5wAZSvkLVVKfKA8bMFaGN+LV5/jgoHbujuQz20r6aPOpfIA0HRkrFC
ebAaZo6mSGEyBS0jdyEJzs6GeTZ7rGMxm3AUkViElPo1l+sywhgOydD+8lcgmG0w
xMOELc9ChNrwVFEQcIf8LfzkRYnbpPDNqvUCF/yNnqcceiak5h0KvDsZn/cFrqZ0
XgFxpe9qXfovBecIWMwI5P3gEFw+v1YmCVNq408vZCGz0RzGUC5gNQy6yVCmQHRj
oqyggHQCQF06cIsbYjpa08NbDtEXgXNeTEWZCs9wkqo6hA546r/ixblcnSCnqNqX
N+4UdHb7ePlHaAjDXhg+wHEdqG/DD/FVPAw5GimYV8mZ4xxAr6ntRdNiuidwp6bU
dN/u6y9tcCsKC4kQEQgkuICh/HthgC5ZHZgVcdgBiOdXwsypl749liwZ6LEAmpgR
1M/ng9qDYyzJy1ZiKjALAYuDvLi9QzwP+eWMId6hIrGaNjdcWDhnAP3INA+saJ3U
5w1AUZ9OC4IJJTE9/MboCmi4Vq5bDXjTDrDceIvPRDaxSjVvm7Tb4EyQsjD0G62x
yHuNI8lkW8j7QG1be8T172p9TtX/TAWvBzMhiZdnUPqq6VDmz6cw4W9qp/yjpRf6
142/O+XUaX9huECmkEos1gRZqQ3Q2tZtBsjw740tDTRoKidCC0W9rb0Gph3JpmTN
JaUg1iHVtvzGU98sItCWjUcVIoLxtAxy40UKeNZIEW1b4YsM4HVjz/T/3aAaVPEz
ReE6rEOuSrqQbx+2JlSTL9olg9+l8T/ysV3I2vHw8LaSq0lOhCkIArbcSq7+C/R2
YqYrVj0eGKWmqqHp5jOuTGBJRtl2vfbG3CujuwawYCp2/DdgETHUyouu5HUsPNkp
WebO/kRYBcmsuwcENKLsykdUfGOB5WoCNTe9nHIhMKjJT25yHjE4F5srF2AmTjM5
hC2Ot6AyfPnvmoaUIS+SvVbSw+q5P/YltpTzkCKUODO1ZsgySohW+xzJ1OcimaSK
YtY1snc599hsHMXZB+vzsGau9kbEp91wDuoALZRcknlK95+ynZjlyV13PLdprjOz
H6Ca0oB72ax2jkfNL1RHegjRrn70mZ0MOpX2dRRH9T3quaXNnEhSJZkHFm4d1VUl
uyeVcNzFtirXK9MkWOwTDiFYYxKqbH6X6o7fFlCMIuCYgJyR4Np/zXGzLWhV/BsX
zlpnBEbYvyjGGGv8A34fRUYBaPHn9WtKYktXe44X0sNZwkSNVJaywzu2cFsG70N9
5EfShb/lw98RpvedibapDoOSys8idaAGly9mr/bFJrzliqfHga9ELLqXEbaWWJmA
TR/g7Xt39tKyMfP0JT8kQ4wUxP2ZQi8Txtr7eqCsIy0RqMUxGOEWBpS4UpElfnAX
qd37kU0Fve0PUzVzSlIg1cNmTDNg2rP309RLCN7OZCmYfztAEYesfzQ4LMmX9ZOu
0L30yY9xf9u8cqbg4fZI+cYYioKFH8rMUmNojwItuPQhvwHh7yiyN90vnLkBbga4
Ww25ema41deqdmWPjcyj68nP8M6HyVCYGgSHGeocBHlgh2m2uwZDNTMtkLOIcsWB
N11B3BbTWuvi8JNhlRLLx0upfPAe+K1nJlHPI6mIww8dsp69utJUWQgJ6GOCN7tQ
2rFbJpfDEGFYJSofmWeBdFKhF/244PWhcsUmvTvr3CHbpIQRtnloovtRqxU+GK66
bK9NTYu3evrLADQIxy2CDGkBAP1aCkvJEiXqs4TnUiG51jjfazE0epsBVDus1OML
E4RnXpsUO7jMegc0G8HLEaK3poXucvbnnfujfpkUrlrIeEdb3dYCnO6/te2jgtpT
yRz24GoHCMvpGyqHgfz0pAtL4jmteBLMNRKkd5rRE9wzfSxATIhaKZFECp03NJvu
VDwA3Un+w7HXt2xts5lDLKN7c2GTVgF87aRnArhSZfPBPu9RsqlV2zVdX+7b/fk1
/HMG6U2zUlHAvgESOQUGkvrnP/BwVTU0FXBHy7FrYVpFd17VL0HvQJFFvbjKP81e
Lgult9hPTiXnv9wUShbtNLkDI3E3WytNhBo2nsnA8D1kr5M/t0POWOFdCBDw1iyV
7gmRDUigWFFCI0jXm9sC2XFKObDIIXqR5amiKSzp4UyMZRdWo+1CTdiWJzkDNEwi
w3v1vaWud90lh+8ZqQqfTCcxeklUJIWLafSOe55nGNnP6lHADSJzHfkJm9Ny2uz1
WFNrt6BdOMjcqQzzFCaxcDk+f/R9PVgknezDnP58X4sjujD/ifFjEfHhVmUu/COM
eghesVJN0V0/qQjXZvKUYWiV49Df9EN6J9Id8uR16IA32aQGYzUxwJHa1Pux2Jbl
faLnlpslj9h749UH6mYS/EICkh6BbI7KN1b8M8yab815J4qBMmlUt5FrqSc3zpOj
GvrhilnLnFClQtMNaIhn0Ead9ckj+j5uIZWRZMgpNnE2OSNNHozUHt+5xmoIRUD6
5tQNVA0I2PcX42MPCmmVD7ryCcAlnDAclOjATbhx5kfOS/XL1EY4l4azwjg0JhNG
36BG6D0wEIfMHEEQAyN/JXwVIeqZperJ9C3tZ9tTFA5jGwTCr+gWpSViGv5kXrVQ
57I2yQaCF3B5h1i4AxOQFDFaq9yt7Xfh4xQAQutA9Ca++mTaKs0sTCmSxwP8iMdz
t1T1NLnlHPB7/G/qfA+8hqJMe9Fqx5sAfLc2kUMFXT8s4SWhbHDj9k4CxGAhFRE8
F8ZzSOyWgc+ih16k1yB0ede/sJ+d8AIr2/puWJ1lyvpCNRSHIjZBzJR1vBxbZxJ0
KHmdy9FvF7JAbPEYs96uPZbxPdPMtj7JNvv3WPhqeQxjX3Qw0+Ue3qghv9gT6koY
a9rasvzpwEFc8UZKdcZyYU1+r7gfVBMGlRlKn69zYfF1I1vZmprk0et6I2hFhO6D
O3ri2vqi0PF7Pyq1p8B4dDreYS6I5sDz+8e2Pr394dFbLOxC19PY2mi+FRWuyRuA
BWWkPwnQFVKMtuR0mAfOAAsoV7pNrKUHL3Djr2gYFCy3d+I1FVdaTCMBBirPsxK0
wSVXbyzg3MmIYhuW4W/NlXEVn3L/jhhGHGaS3uf82/sgYGVjYzAhgtcUApXd5FGu
b2zCsEAlbZY9SxLWGmNNcWo45hqcREWV+Fw4ss2l5KhOdASuzm3VWfMWuliSqNRO
rwK7DDKKMENAO3kEXY0sRGu8wLjS/mDDFyrZIp8VBLwuo6iUOh0wxP48alX2X43H
SQUW8pFTu3rzNUXoFHZIGf9hgxE9YpLmYWkpp+eAKf2oOurqndX57UVwdOx0hqMv
3xSukaZn4AaVVPYYTjHFDoXaukzRaO0xZ4GIebEJy7eUjDUMg9XxFD+tG7ybJSaH
2kGsHGwgKDWTnPXZbHPJRqWHD4MQEv2AZFOSned4N+vK5+bgCd3MEEHtLV924XkC
Mxz7g6bp3+BPwnYtIfUp+AFD15bjQ69lUN2V1Q0a8ddegCD8nWObBE4I9e9hDfDX
DhxsWpEfqS+YdWdjF0pOZfXdDX4w7canA49JwGXQvaC7rOB5Ni6/G1AaKyxPtt9J
QaukzAL0+0NIT8zM3/pmOm390SHgFXCbYF7Jll6oRHvHVAuhI2NyHq+2LhJZgr+X
85Y4/6w+7rJbDkeDjZoLRARLlUu/TDvYU/gMPk9+IFsOsDBOXSCDligtCutMUZ/j
ClBj/FRZQTgEVvpfPCs5LJF5QcvLIhVjqv9RE/quZhpLFkHiHqKAHqZgNSmnavxa
ft7ZRFck3QiPbY39EIxtnFEwf5MhaJJJ8v0nzAmVVYULztB3LYpuKDdLae6VM5yP
bV99CJX4NHmU9LlSwmXEUDJtgdcktIa7Jm3CMwH36Aedan3pLED/i4K2CSNNQ4aX
oF0iGM3+MBSwsCT8zn3wzagmjn7V2LseLQPNm64pkfGiZY+PnlOn7n5tForCzDrw
obeTTJGq1iPL80beFKB3vRxd7+JJzKDMjFjJmXASBF0HMSH6ew8SHrgjAIuHpM0X
zNgkbkLgDSr64fHcgO5oBB30NFiBwQxpymWTGdm8jcCdZJGeGO08hJQBZW2bsTvF
2IDM5cgFLOul4BJEDVQxyEEjpxvX0etNHI1CEdJXyMWEH8OlFT299nXP8PiOWki9
4DLvR0qTaVWXengUalQZRsrIm5hwUOKMeaP+IIpDMRjIErfplfyx0YWdFC9ig5vm
H4vM/orYqmidNP78QV9AfWQUqhCro8bMIGmXvlNP3DRlkZkFDYA90AcOBxRFOFhJ
a/DSPIUApOsDXo7WyZ3SQLrLyD4ABENlHAhMa8tSi9CprfSTlHQ6GCL2GJlhMUjA
uVWrHBLaVP1mEwMi/p7AnRbVzsnml3dpqjbZ1ytOqnmNdWJJxqDhdlvg1oecySNN
SohXCeWoQljRsytCJYtmqWR3Hd92i+tha7Y/0hqTkj/ks11/yj+8oYQBSo1n0wHh
LoW/H4ugt73RP/gtxJtPnppHFbJZzxIlRFx/UczS49casJ2VwZDE5nn/aeq/N1js
HvxM4oi9ZMlhNn5fBi/wv8nRHaM3guj3NNFhBoeJyQo8gyNvo/R2cD6bntAeXkM8
WfjQVjgAr7yTPsKcH7x0Cgs5Ar3qDWtUN956cmKTXYyoEtCrjAAd5cjwqpYgtnI5
tdTZotLeJ5Kl19NJDiwVR+glKaBmoWL72Y+G38PBp+squztN1phdTkNm/u8sFVSd
y/cdIVi7HveNTO8wjZA5CPQaJbM98sVg7jI3FMfll2DzQpwwNq7dx5YdbjS2R/+m
1ZVjqoNmOV9+a7Z/uEFxg0pIPFiw5FUencMuSDvEQA59abIUiizyC4k2Qml+e/Yg
2RZ9SGPBIJFCzHsjyN2uYyundd6Eo+svKyN3QdBIIVqXTFbeKuENmpAB/+y7Oc/u
AwLKz7dI3+mRHwSW8EEAmrNU2l11GOgaRaYeqTqGTWrPbA86vqJoIXn/GMEATPUW
M55bUgCrU5qrX25HdFvbK5NdTftPtogUA+wPxaQ3VooEGpWLQp9nFi2QX5kFM3De
WJhniBDFOcOyRe5WYCZ5/+Wwq8prM8H6gQVPBy/N+XVnKN/4p5Y0GWRVTZSFRarD
FPX/0QHJTMRO5Ie+cKk0MH+b1elEa1DRPn86tpQoE066vZGGaDiid8zwO0kKvL7/
dJV2edbftS5tscAoXxQ5SU6/FbGD5KYKfmVQ33QB2+1JhpwlAbGFP0xjtFQXBdVH
hak28y3RoZwz6Ljv/YpNK23lzFrpEjKRgmfhfzJflYl+/zyyTWwTbOuQvc+LHvwX
Ssr9/twOhT7+opZMJ0JIJFarDOZpzRiAcEHlUeigbQ8ZQWHMr/Od0r4te/ZAj/Vf
2SwPp9fwTH6yXYVW2vG/19cyA7qq0hFs5QHpMXBXbewN4qOhQvE+/JUmVr2tdpTN
phaAZmnO5Jgpdwj7IN+XMchZp3lDX2W8vx/NWV7yJ84S0bhEH3urCO5vapALfz6V
quWFY39jvExDmadqJeQr6dVcCsXDKyTFvnPY8wLDuFp6KRuDMSRUfmvlqcK9cWgF
c9Gy95S38Mgt1DrDzQIavw1w6MsgU64aQt5N5nV/whwkrQO8roF/bbetCzCEWqlU
I5xThu18wJxuXG9wJJTZzbH/jyJ6lJUnYfFnJDpNbDVVGZ1v2LTaSnQgxD5MJFtG
uYyIdQ/f19Y0g+ZR0vhXh2RXku5/1jg5dxrJ20hs2YRJPIShKxdzAJVITxDvMwTe
udCqSqxhYgd+0Ik3KXyM6EuUAQOd+0DBlZR7D/++anLgjyGI6H+laK3SCSCa1Fhn
+MASe2zgCFuaZhd5s7XA3KiD0WeAwV0myVlHtXcmACHYISrDGN0sZb3+w2KI22Qm
lzHklRrtJAOE21AjnEj1EfaJ37hnIk+Ue1GO6UvivabONqs8ywY3p2OezFYC5pFZ
H8az9or/v/xbnuQDGOJNu8LisCXfe8B0FFTgr0kAJQbnSBZaPrAOkHPW+woFgvEN
g78hWlkJTmZ6yhGfl9vf67y0f+WJzu+QVdXJebTV377I28Wnn/pd3u9AwnUIobCe
RXWqqoltuQz5wYQVjXR9CEgI7yhCFwgmYI0gI033kHalSlS+gaW61RS8+kLHqxdL
ApR7r03nsqcQkoaR1U0mN2cX24+WQVP4BiN+YXvV9E3cq2w7sljw5iYJUOnzMtmu
ukSoBUkQpPaYWPGNQE3HHPJMecYUQZ+tSVPT6Jbhe4wQhTvKngM/LIsaHfxS2JIS
fs9chI70k25v30RX07ZZZ75IeuAnkYDdNkYA/BgDwtmdpbasqH0Mn9PVhecLJgMd
q99NCnNDg0bC+wvw21sbnH/yGvqLa7+r/AyYKKNmUCsbfXhPD6YWDhwJoD3oK3r8
JdqFb4UyrZVlGGXg7XmgqSJEGuMGrh2kLkm/5os9KZxmVpY4X1SsMTbZifjs9BQW
1Rdnea60oE4ooa0vczXS3CSiJvFudmPx9wDYD3CrxXiZxz3PH81k/k31ERXX9vdK
/m750pyPxdAN2PybjmjjXh+RBDcPxXTq5j7ELC5z9EK0wLSx4EMx2BrH1bcu2Z9M
jo9MzHhYXWtqW6bN/LQbPgScEuvDTMS7ooGj0O078WZh/5JYSPeo8SghZF5WgNDW
q19aJAcYd+aAKZEHcLTso2ghyczeU+3qgKPgkP3GyImVu+syAZUmZgis5ncAb4un
/6r+BP/vIyWgrmHXVD4yt/V8691HEMiBFf4oAnXhVFBd1Ss83+NirwGNXaHxBzbc
GFgqPmDxY3Q0HH614FfgCBlz/ERxiS2XmNFogdEiPEbxLRkdu+oDnWm9YVaUd555
dMrazEZb8C97qC4NN4e7KboIzCd/cd8cmykndP1hUDDxj9hptm6LOE2tia5Igv1m
i9C9+OagUgBEnjH4LVjqxn8PYHVN5OlvoRKMGL+4iEHzAGdXWioe8oVByMs7bdC2
gL2tUzOoR3PVwjNlGVi31Ak709E4Vu2GC5njLiNix/rCeLGbO/Ma0JQn7UEVZ7rZ
yjwE7fVpuBXpxjimo159M2JaGTwcrX2ytaLGnfME5rBVN4PrA+OfCrg5j0Jn1nL3
aBPmvlN/E5Lz7NiOBiN5fg9s1HVXcWiiG1hV4oSHeeEJ10jNyCtxNJijrDGfU5QL
vyddZMcnp45wx6jfxIFn/lleFxBgrdUqQO9SCr+hgAF1pdLOCTb5f5Hy0Wgs4BiS
2KDWAOl6HI/BRAbaQHJEt9SnDM55W4XaKoHPz6E5ymNAjHXtw7z7lRVo1rrYnmnM
v585Klq1bsPDW0aGsvGqHSPoX5lCX1NY6LNURdqUN2GaCqlmsZxRvd9guvg6SxPS
St86WDF+L6XZ9Z0WZ5bE+bVqvHnpiyH9rCnzitEu9en35nHHBm9Eq4CL1KQGiQaq
Fkfh1a3KVG2PWiHZncDq2sLxWFfDMJj6cv65ClDg6CGfn3uxg01zX9mgPN1zbZCz
9xXV5mmeyyHpNmF2Ou0VSWjeoxI6IlO9qfgFhlVJWsp9NntgKvEYU2EG+yxhHWod
NxgILEMnP5rW9czf6l4jovF0Bqtc9mn3tevhawQ+lEQEsevJGCKXgObrVYhOTh1D
1UAxgWsJgs3w4ELU/Vg+k05XpRAZJjPZVsn4P4POPWo5W9Qul9xx79/N4730lYfH
OoRAJZRN0Vs6O31ySUCWA60tlddecSbAQph7jN2UoxfJuYuosufKSmCfJQVKVPls
TQSltCrSlSqU0mKJi0o1UTrMjU5moVaZHxInKI+M+ASzHxO21sOJme7ZssMgfYEw
KZI71sgbndQAbGzY7rGcy5mEqnOhc+cQc06k8eXvGd75UxMP6pUFLsJ0vDLFluES
BCdilq1dmqrsGbF1uqmmed3prTs8mpC8T6jKkPk3HKaoHSfEiAD+RLf79r1LaG8B
4111iQMzHo+f9lr+sPD7aeqMansVYvMVMvQqbti3tM+JPr95I1wyKT87UdkQSInf
zOPKvfREU+hRybPPq9JPtHxA4enEjWmN3EFeZfhX5OgHe6Zcqght7ngckCWhTT6/
AD+zmWHE67M9k/0YP+uRWciG+o2vw+Du07oDsFBa6JVnGgC1Px5fpss8Bu1glacF
8aV+cdauoidRu5zkASieIa+nYKyvH4PMwbUKwLq0OMpAo2EU79Uk17RNoF0W+MfW
lS9lMcDlXu4nvItillRdiIWxwu3BD+NhFgmiCgN7uCbIssnLhrcHvU84rm2zSsyN
vIFTIum4KhpuhiMz0T0ZHziSc3UKuLGVLY8Baa8t5G2WQpuGlF+1e7SyTQ6Mb8yX
idtu4hjnNUA7A1LFoaYauXVhkcwaYwuieHj2CtQzUhr618ehnoQjumBxBqh9aJAs
hVneg+pGnicGFoGrY5FE1xMPgU+bId8jRTxjIb+mgYu5uJqVZ6/B+Z5xuVblv6zq
R9eo4QI7rnP3n7/g5M6EJ9DvJZl/l3oOwqGItPCITOcLKAVdDXaJ+wRPDOoPq2W6
WzQ5RC1CmkbhpdXf9XvK3Dl7who2lUjOAHa+z2VkdXo8ux0hJKe6akAwW1fSqiuw
aqMYAmQMgdzZ+NQaQed+bGjiMhFgSXIVDNDaIrx5tz4YCl2+PA8pq1cEIuw7xGSH
wsqMlgCkDm47+FEJJHZ/Utd87uiwd/8twWeZ0l+GqH53TdZO9KMk2vMJyIV6thbk
frXkD+R+Fv6xmgPlaYUnWSGgODlpGXYDcgxF8AbLue1vi33Y8E99sQ+8Lks1do2l
BVp2fbisalnw2YGl9R3IFBaMAWgFeUv2sDabHYnDlIzN9bx43O6OHMLF6I8P/O7W
qK9xB1njQKaHw2Pe0Vd4DsqlqtR8HQA9z3VSFvzONhGouAxrcdB9v4/AQdAXh5/M
wXWKnKCp0jUfRZo2xScvr8H2fFewgqVTPXmITykBXEPszSCMxzKpmnOvQNIA+JYv
cLZocikcBOCwmYIj4ks37pXbft/TkbBRxKcny5i1hd8oAam6d2WbeJJp+H3ILRvP
tGllvJMdqi5hpd0zGvGQOE9hRIN0ZT3l5aRGQTKMFTvlxWds7CuHIu6PzJ2Pl9yX
cbQIoc/ay5gV6EyYlz48JDiwFV4xbMYWkznVAXNI6EbnLNK/3Qj61Os7yX7PRN8M
TpCyr2BsvSQWt/GjcMoHsZk2E+FRCptya4zgzTFrVkz6CfFXbeFoy3Kg0EdFxbAy
pBupnJ7f6tt6yoxB5q6A6sc9jqaEcXDM8GD+IsUVwpIgsbCyj+h1XVoDal6lkLhn
9847su4Hr4ZuWIdV3QLmslLV+bT5zMNiC1fRSEPkaYuxsXEXRxB37F5PpzMNIcCy
+jRpzuN9ls3B9uB+GOen+jocx29+kgfj74NtQETW5yhtCekdljHlJXhS41BhEn5V
WBPaDbTwKmSAeHCMHY2xv3uvyBehJa54psUJrXjLQsbJztwwVMPu15SkWIfdbgEP
2pw7IJ5IU6FZF5AfsQ4GJ45ww/MptldfQTJkzQmviTITEddwdHy2H60kqrvjp288
LyQkNOQR6tlppaPUcUfscIKsPTBTee75JahBNJhIV1YMihrNUSEuJzP2ft1E79YN
in/KSFDo0rv/Wuj/cnlHK/Xt5NofDEn+T+dp9oVbDwqaxRzk3Dg3udpakTCX/Zrt
SjJtKBupwrtT0ySOxPsydo92fW3yB/3qCxuh6HdFBUfS8XGD/92VspoOYIR3PuLU
md+ku44Jv/GOw8grHVlQvOgH3pdTAuWOcxBT2nqeMy5qGOFwPMUQkZttW1PSmyjn
JfwOmJfd0i2YAJ/0cdWLBPnjuz+SLEnQKE5biwXg3UV2CI2h1HCnqQ1WVNpdiGdp
hd+Ze0OWwuTjP6eEkoG1c3AqW1KQGIkF0DnX8UeEPtnA3znv0+HoZP9K6ktUaiVH
j+L52in4X3JfD5mjQs6QTiy9qVuNJc0pcqtxxxTzoRFdXQih4xkt/cp2loXc7rjZ
1dCmaQVMKPav+s5HeNNSgy3H/d94XU+ku4lo4N6u9is1nohJUk0R7sbf7vjmfCox
fnQkOXzkhzBxEBw20h51xnyUbPDj+rzCA2sATwqQie7bEBxBfnK789cPMr7oYTgC
ljWZxpiT0uq5ImxRVFlsDmLvUox6vjB4LVurNqAV5NFUNbw5t2AC55xVzlfIOv00
ePP8Ps8Bo14cJTcP1VMkv+TEwWhz3GfkGJ+Rq6a38b0wBjkzbsk6fRoMJ6oGWT3w
dBG4d+h3GbeYr5XnBNgb4RgHmw6RfGktG8t4eIhb9O6mebV1hmtfa0qzKVsgqNZK
oIjWthlEp3eGexDrnCQAKfyfSOZReg5ChhexIz1WYEtA2f0IF8icQxTRbxWq63Vb
JasdKnqzUYNL2aZuwIsH/K7RxBkOd0PR/pd+/52+RaVSaJctY4h11lDRvlLFDYxe
nwXNRVTDt9bgPxT34EkV1OpECLx//IvvkLiVoVaBIPsJpyspj+MPmdFdJzdY11Ya
PfaazBKRDFdQB0Vb9ZQiIY7Peq8674Vc94l1q+OtDZfGu+l7c2lEyFH+wtXbE4Zu
m3gvmCiwbchoSzSh/0uEM5Sw7xbHnbSW8ftX45UJgkVtvO11zuZS6m9uWixg0n1k
RQuWDwuQBD+bhD6u6jU6uOclEoGFEngtEiDQJnko6l96xVHskOGRb94TVRRHrovH
0i7W0KXMdLfN5jHlo0BVoWaRkZ3LwGOcLjmzahzvBk9GLyeU/7Ocv08jY85YgiWS
TjvEQvtEGi8WeVqNYlVJ5ELyGZ91615vbpWrX2/x2+JEkoulZAioX7RNy7LbF/JC
FksX2YFl/uMQZJJDgpr6nQu4nCVl3k0Rfxffw78KsgMVLT3p2aWC612CyqS92Bhl
ttXXKuLnf40iJ0PQlK3kgDfobWpCQsJmbMII+ijWf7UISCusK09o31hL8EJFdQOh
8J8efxjvqkM+iKbuXMjKZjfUf9QwPx8hiiPGFwS8sJ0iWD6BjKAR2Gj7cd8c7eyC
CSeMWaUISisXi4JIpVo0O9gNyNXgKH9fF/xtQ+RAQAbWPrEihHbsJsBzAbYg+8Gz
U0ad/Yw7y/BuLcKjXofQbSttfk9cjDJAOHbHkrvRPMCX1EiHgU3nxJbAQmclNpms
mpJ42IvJu5lvsGlIot6aMGPE506vM/uREJCJaDGd5gQifbGgyY1NkS3KcObEMrP9
ySA3AvbtBd9hG9Z+8MQbgGKPNw/l78vIa/cZW2iAjluBqXGHZlTLLGs4cwV0ZfOy
jLHQx4ieR/X0FnJ/lKtalspvX7zFrIRdAtW9dAccuhF/IBYa2gL+vBDfR7iqUa6D
4Ts8XbLn0IEtWZ/1fy/5zveI65AKusgtK+vHCq8wCJnVrGMxnC+1mBXm+nmfa4PK
OioliGD9o78WsJ7h6V/43t9fnd4XNqyPjmhRh30qjfa6UH8FNUXYNhf+chjIux2o
9o29/aMxCc3KYAutPANZi4SYLaz5gaA3ommT5LBovWmx0lKxBkcwvtdOk/7JB8Q9
+ECYvUC4huXoG7lAxdjbGl8bEiLUzurGKjA1L7gfSB10sOBvCewRL9YPRnZfNgJy
kioErI5jSmcQI4qdg0t9jcvcC4LrtJSMKVRMsBay9DzF+bFPtinqwr2VgQpIZL6q
D8kctjDN4jqlQ7fEp3/hqWahQbYMXGJUN13nBDnTpEdhxBrnkoEx2JLN9+WekuNk
1KGymvROe7+L0mi5FCxwp3pSxwXLYHNuxL1Wqd4CYLXsGJOM+SX+yv20ED/ut7cl
tv5V6Yvo0/gD4/xydQnweu4WMSSINyqOhlwVkYWDGcnbfz66Hr9V5vpjuTUFGel9
EhrVpAPAsV1hWqOgbITOt/1BIJ8HvQQgtJtzMJ7F6a9WXSFPoB8I64HMcTgu8t6Q
v2TP724ZLUDR6YnfYe83FLw1BdRGBg+qFB1230VKZztCRKvGZpxGj2DxYbuvrU1W
EakRNeZH8Dr7iknbY9AkaW8yv1RJyqfWTxSPCfWdVlj9+2RIwnGH7eWl6+yZPWSY
G2chIPKJDJDBGRsZyqELk3GQff3XYN+WKAgwyC1UYrsUdsmNmi66B5WKPsUuVxWL
YUocTf9MUPsYg2Xwxyu8XSN+NQxwordXFRDkzteUpKG08NAmggI1wQfh+pWFgx50
UP5Zzzaj33vFJarnvhdgOnVygLhxYvFXYWze6XmwM7lFvzyrRw7K5bOGmiPnokFL
iGMAgXYDgzzQkkcGrOVUAetUlEIrE5b+kKKIavxEGzcItdcrPBB4ZCrsvcUmCDqo
USb7QU8RVWCMmai6WZzb57OgLXiGBiGcexCa50bnoyocJRcZ457JkOK8x/y4nAQC
VWBdUyMunUQM9sQRs4HqT6CLwcz4Bwl/GhrKJOaEFwqOxzWHBG41SNNOn2LYySkR
ZrOHNv0kpuMsjKqjThaSa4xdj9eD4tkbZmhJJIQq7Wqworsu9+AEGcsnamA/+84X
8gs9mA4SB/d66L2RN/fyNaGu4Y5pn2HwSnOmAW1g8aBdCbAI/+q+KAaT8lEs2vA5
IMp/WJZKrlEYmjrDqCNT8eoaGFs/BhN/pSzAR8qCDmrGM8udkffZNDzuP5vZSO/f
cqTryqk3v+eUnUtj+S31WYGP0ahlxgKSQS/DrCqRQRPdJY5QtAF0RF69IejwBCMa
kd0vXPUXFLDSLOdlIAf8imIFeKaClu61E4SMB419tT2FBY/qiRU1udu/msjSyy+w
aUxm6cM8ztcrT0/S+w4+esdsoL9dHOxleHw6oGlJKqlw08J4hCxUulvHjsj1bS97
z+qMRn4ltly6tev+9cOF6AuzWES+HT+QuS/Y3Q7GGc3YZHvDAM/IODPmdmjOjyaS
UQ7cMMD1r8Vki5j8/SM8Kh+2SJrVYnwc0wDig74tvRqWbNBLh7eFXpmhCx9n/mkR
Lg8lOp4/ywxZ5p/GvwgYVKg7QNal3QS3VRE+YlX65jBDzwRZWExrTwPgwssEaw7p
dzNLreEWv6Qx9PBF6I+mWD8nzGOvpzfXy96YH0MvECylRiRiB9BpXu/bOI4CNuJj
2MG6oHtWinuD9XwGA4FspvMRkARLVHUq0Psoekmhcumdp0H1EDyVER7A0g1HZV+N
ZtL1pwD8LjZt+AYitLL5crd7zAbFypVczcYE4y5Jrj+NEtCInC4JSPAVeBe9iJOk
rW7Yb6bk3ip+7YvkbuiNUT/r3fMLgmsZYMrixhya0yNRRvp+gnxLaqRHtNr2HEY8
MBzUK8YxRcWkQdj/ubkbGZaE6qM/n6s/rMU+/2hGBX7UUGVLDzuNkS6f9Rhvm1g0
fdJtzFsqY4ViVIGqXaAHO5WV21pa+b04o+SlezxgsJrgRsD+bDmQh1R1wFouT/EN
SWSgcg6V1UbXX4a8BLwhD6tqr2v5qhD027ZN2XTJvGKm5grkwzvDPw5iY/31ZZUU
ixfXFYT849ugxupijsR0F1Gri1aVku3fz00RLrrhLlq2ff3/w7aTlqfSjz8e0OKl
s6WoTiDJthr6yu2rHQ2gmNGr0ThzeqvwZSqDH4AA04UD6XDYRgJhouZ/XjA40yz1
b/89NdU0gRb6CD4SQIWHHM/w45j3uy3coPTIhrJOm74Vkak/HM5C+5Jjtpx77sK+
w3fIhKk0RgEZxRZDjPLTnOMbBzZP8mbvmiqe20J7vcp5BJ3/g6Zl+JIWqpWHAxR6
3Gof01QgF64DM1mygW8ZgTx1IotBzpaNsS92SdDsPn20+fIk1XYpy3mSjPUPvUgs
aRC+hIIIxQDXRa9ZppSNbM5i7GREb9a55lwLl4gEnYkwt5UEs4RyoMqbtFnRv5kh
I/0aUUNr67Or+5ND8bFK//geeL+VNVupjkn4TTcQ2Q5IfhoMFmKYWgZcfGxugcro
cn0Zqke8S5GlLIrir+X99CHRN+mzYOqBs4QdWOZfVNHQDIvpeyV69kz5s0dltcsG
eC0l4Jvht/kh/PkRvM08apjymn8aUrsg0JVzWfRRLQiirXFlv9j+S0R+lNlT+UrV
vBat79qA8E0/+de8djkQPLhgGY8kXjG5NRl4ZG/QnY8KHAiVZCW1RgO4MpkBbdxj
gLUdaQ/TbLUSRHZJUdFZBiPXzbWn6yPnCw5mfY6138sWhNbO+OU16n6Q0nzAX81E
pn0MQYizK24g3QTIAzykhroRk1/o2LAOr4ZcKkPs8FcJNzNrMeHmMAeVgrSGkYw/
h5vS5wCdqA9P7PFWn5uwyR8onAFtF4UM2gnocwc2LuiyPoXrS3b5ing0QkWGOz5x
PQkOljdZIiFXWx6qqgfKuGBMQ4XWrEfJf0SCQLZEZD7YU336gdGpueHzw0KLyby5
CMZNOn9LliGDqFjlqsVSICFXMVQAdczHLVkEce8wHQTKmpMfs0v5HUcO1lrgspu/
+C0uvSTpK7ov7KjlGYNsZyRmEPvSq/DC3zAvFgBbYj1U8IJsl+nNFWnA6v9R0sMI
28MrEMVcjjw872lTilQcFy4U+BwjHpBU5ZZ12MXl7iTHZmF0cX+qDvMG/Aj2fEEx
8DJYBLp2X7fAslug54KA3KqUTZVdpH8+mX1JrkYEDICyIlKuE3b/YcapH7d6T/SY
HgfOG2qPq0nyl/QIieBZEZMYkCsbQu3O1ymRIHnuK/o9/vvd5hGWWP3/Rx5rMGqQ
pNjvCZY507L4gcrPfXPqAq73tWtqVOEJG/F1tcB0LlT8Sf317SShVwx+4+VP47z0
ofacJBpY9EiiraZs95Fm9W7ZF4zqlhC9tjBbARLn5mII6lBoGPDLiWgpPCQUDJ1g
Z+6qowgDrlm6bXsEbmMrEa2opxxdej0CjdQmkASHbLR6/JO6S8LKS66VxuNeB3P1
CPRXiS2j+Ixtg+kcztMGS/pDRtdWmo7z/WhxIOwm9OfCGNNM76lIeV0+ulTtygMD
R2pPZMapgNeRJ3D19LIDiy/AQZ97pyQ4OC7Kt/u74gaEvI+3pbHVMc+xRd0CRgfH
8PiIvnW4rb6uQeDtJScHN0CmaH9/dfru6kDbP6v4wzIbWMVy7RlG1DVWryxwtmY7
GFbnqqmAS20MhhV5YA8a3D3WbvDNRcdVjycn3tInFs7jqjnCp0jU4MHBTP9vZItN
tdcsx3oppPTqWVtSiTjN8KM3f8iwrfvREbj217ZK3Kc01sslASCKpwymfwKuXAFy
Jl6wPTM6C6WSA0D1aRp95u8zJYMh2daWTc12FAJUtDjxldGqH8SWO6YL0/H6uCg4
EocnKsflou/1LY8TAkEZve6bXW0lBe4Qo8Lha5mULoHGc4IsMaDykM/DQa62Et7L
qzeVG4jzEs78AeEFlgyKuAiW/HV8GB8FVI9h+dXVxXO/TDSdmDJvb1j4AGF61jOE
d4vuwJXUNSiMQUOmnP3XScMs9goufaV9VxIykZi1+wu0XgeUgRv8kB+kPf9EuvtY
SLArdQNmOOI2WfxU4Z3FJS1ZB7lk6xJZds/cNKO1qauL5jeIcA8H2WaBJNuMCiLR
/yvYJ8feW2EPM5sdJC/gDQE0QmrSIPf87VnenlsHgiLC9T+Zd6bCZJrVDUrfeMTB
ZTzwIdDQy7e1+1hVtFv88GhPC1jstRFXQf7r5QnFDwXuuNh4owGU/Ge91wLT0+Em
HMYSTAWFLslT/q/YvlsHClDfhjf7bVt38nsQjUQZ9s2rKhUOZQ3N9QzZUn8uZFZl
aq77XY5VZQyHsSGQOSWB0Gmi6K6bkK99W4je1JXRfqglSo12OQZLNJbmbJwUL59o
A+A57dh5Dd5z0xBl1nOgsi1hLccXmf0qAWyb5XaIZQthP4TGG44dHZEgLLvqG+br
IGiZXAxEPXBYg6hLVTqWOq58ExQZYg/aCLLyWtCUu/e4Lr6v7mRz0d7ZeVDhs9na
twVS/uji1TupJrlKsrzhlPZdUiU+eFKyfnff/po3EDMRTN1elZeAus58DEgULAgd
mxC4K3L1/T0Fw+pOO24URnk0SJlV69WNAuSzNqZBexs+nHJY8Tb0k2+1oq7pMhX2
c3fprr1aYNP/7e3TKOwgB2Lgz2U9IckMC87T6Ep6gmFp4YZfgxTuk0WWXHB7u/0Z
pWk8o2WRPQSyDBE04Wu4WfD21rA4HN69mwxibOsobFlbryNiAth9wQNJrSxkRczG
s6uuVSqnQ80puXeRzuILuBPmKQSAV3mYxpKg7beSH8gEj39gHEh1PICQzKT2Ys88
Aa9C1PPHIGYRNi4D/pLmE4E3QOXFqkrYrFWoJtSrf80uRrV/FjME9izq5IHQP/0W
NSshjMLaTMFnfSZe8eos4WtgVhGmnSHxxfvrQ9cnODSeqSUJqumlX8LmMBbmKh5f
vF+J+HkvQuZxnSd6goINhfoLjnoAHVgoRn+hCrlYAMJon8P/Osjkycwua+FGUUIE
xncW8CVDSu66JnPic+XK99NrhQxomk2Jde0GTeu0obQND0In9E+FknrA5BQFtOAE
RVQ0FMh6YIN7wj+AnOyyofz1xg48LaHLVD9CuuA5RG+AJOD4X0HHC12C3UfuSDzb
N1SVOZ3YvOdWFovwmpYAZEFi9SAo/tlImRVeLc8XqsasreWY0Rq6gXi5C9w1hcd1
3zXcWN99NKVrSWn0Jw8f+CzULl7BYdN9qD5nNGZotuMBkwi1DfdQ+/UTuJR9tQlV
XAGEYZEPwNW5V1sFDzb835ttWQe+lPszsSAnA4raZV57OQ1BiDWioi2UfApKot3j
ZxC1RTPOpY/P9napZwdzMXNq9A4qKrfNEm4o270xBC8SJM/tF2mmGZMZ4YRcWRta
LdbFFsPiK+jeikGz3SQsZkIRrtGSX54wZnidia4wKIVb+YfgkoKdTsDedce0ULTk
08Gu3cHcKVkXq6A4qpAAGDGBaEQQaYu+REq6Bhe5zlBsUxsGObEeq+tRtM7y2SqI
KWddQoc8qt1bupCTOR1jL/sgFfe0eOgS1oUhTFFNpy2U7j+TNlDrPnrYIbcDsDLy
u2gQDRTRmwYPRgHe3neFmRP7gZVRlo9w7dnOeRB1nt9faFFa5MxOjze6tZ5QMoqn
+ogaKNMfJ4+8kMT8FPIES+DMa8Si++82zZ+D5pE3JjH3afnkRL66/oTnkIXbAadU
di9F/orVc/GhMqRYEmmycDk3YwbUBNJGIwSHn70QQ0LPpziboZxnt4cGp27Tgz0c
PiZxpl9LTC+mC+uJ+4Gkwc0aE0ZUyPNmeNggAjt9wQRyhH+xQajUXel1px0c6tpD
67tKjhS6+QAcVTIkMdJ1mFiBBNW1pMAUIrq52OZ4h7OCjV/PZUirs2X7jTI8sUC7
8TJFfzW61yAYbhKGwgpldXvu/E1oOI77TA2gPf8qaJarF3dikw5wU9xNQc2ddnB0
9Hoolun3AIFzpi2QlnYduteiZKWwyXUnunES8vx+ON9/0shYGAWrkcK1WL4nN/3d
LF8ok9vyLUq+NbY7P3kS4pCy0EyPalHrhA8ZnUybhlXGolFYHVr/ramhBSknrF3W
fwuaq/UA5ajRYVuJmiaZwj5UFkwGv6/VBVM9BTqJZMKtUJDE1AZhJ+lSvclYi36l
OK7BP4aEGGYV9FDK57hDqsDMwWGn1oUY1R3Z25t79Rri+BHZ40s1rFBYx0y8y0Gl
5lHt3+lPER/VhaNzlk9raBU/96n8VLrkjRrU5ej9JFpINnJpr+isGL2k+H6svEpg
xBTCtGngnDImYQmqOMH9TMkChVfLlYPRIlyNUxnWLmt4xY2GHU0uOFKSQaAUmieu
CgBBEUwiCiG6laK2txg6yFTH72vhJzjpP8VSIyYu4EiI9MbWz0Q9/cig3q3lj4sp
0em3R72kg+ms28TPz2DA3kMDHY3IWJNG+8N07mIOo7npfHUGX6H+xeRGSoc1Ybn6
BXUjFXpFXAWPmKfQILc7+3txfM+5qkfCOvqScCsPQpAG/o25nlNWm2u/FbX5jUnY
uC+q8UIWjrFUwK3UgxdSau0DaiZpj6Azbp+89oAwzS7JIaL+ALS3bQXzJZDE3Sg+
qH6aQz/8xCd0hdthiux/uLKdVaJ8CMdHsRyjuY/uYpjeDVW9iQc0xrWF1jeH4f1l
brb5+xRPsAteHeYMHqTQDX4m5GM1eNKJT0aV3b3NxQ2usqYfKVtz8ERygpkYVzkH
PkrwALbCJ/qYsIkC2ABHT3Bl88q0cNIGFA7fMeZPAdXAXZTpHZGbGrsxHASLSyCG
vGsnFEpcnSNkqotoBEyKPOmKMpInJskFfG8FjQzurWJgwjp/P7/33Yl6zQXqCVgO
nitcLfXsP6nUj+GY3hEzgQSedvn1OWTAXQkbIXN3NmWgNbh4bYbSDGXe8ODNzUQc
IiCqu3LWw3CuJ++gnQXz7ktrz5hvJzq1MmMF1eB97ELQaTYhfZYbHemeJlw0oZ6d
UgDo8Kd3WDrbS8ufUvwPszDYeib+pdtHuvCK6D7/7MT0Ze7XlBjW16hleg7iHraP
XHZQhV6d6j2cVBkeUN2hsGfk1SeiNraEy/kMEelUiAzF14EEeOml+CuJXIwpJiqN
1+koQ4cibMssqYtwr44nkVNrPetu1Y+YzuPV/6KfNTAGM6DjnJOQJq+IlxIff9Hp
XUXx8ZNZeIZE0jMkRpIRHoMVM3ZxXkFg1ZmlQaSs+mwEnvzA8LSOcJeoKYwXbsTw
9RbdUSXUNss9dj4TlG9yPsUCR7CiiEyLD+osjUqMHsMAIEDJ0Bk1zQ10s3azG5j8
i75awFuHM8R6bfDxYVU9MkSCKx7PJWdPx/9/L/Xc8am35tM543HdtMEdg66ZXvM4
Yud1vgzP3VYCkxZkOPAxhla2Lpnz5Vhj32szkIGo/wSRTsVqrqkwFo2xSd/XXcEi
40pELavxf5D2u3i9I2ixt1NwPwGmmHmn+HNQoMlBPt2fIw8USxBvan1iKgg+ishl
VSY2kFvbxa7Fpyam+9n8SqVz8AQFByGo1DcdelTQLPHKtPLATRYiBxPRtjmxzCr0
SyzQ/EYlJZGoEyEfvsRHiu+qyhOl2gJWGpcp9uGLG5jngU7G326jN3UMwljmnPDy
UbWdUoACrpy1dny0Q+FM1VaqejEv5V/PShOd6+o5HLthahKu9c8iMy/7OfsQUPjv
N9RgZjkYA6ohomN/sq4y40H+DQxh1BhTIvHtF+sDVppa42J5cefYj18TwUOULCQ3
oeZ58XVJ5bFJPSXujwLw2EusVtFCW5Gf5jwQSA29Ft0UIFEJMsQfUmYzEoMZReki
Pescjab0LL41yF3ULDVIxOEGk8Jm6gQOIJlYtBOxFZ9udTqDTMOf57IFMteqc6LB
QNrXECGb213OsXNMg8RoBJEK94aoaz+wqRRplrNG3Z3bxDHD389Rp9/+fUDgE9SR
LUPj2jC2x10dfMxTB9Cuk/Bee9d7nlgOvIowV6K8LHYPlmPKG2EyMLhbNXjFTGL5
FTIU2w5yAwJGS7oN6KakJ9qaX7t8BARWwRlW8qRz7ki3BOUOQ80N21hk3/fQy+nl
TCCsEo6Vf5348skjGmDZrnz14gagrod1qqtkTRs/2YkgK0O3sBMxFk7509hJI0XM
G/GphMFY6lyS5h2UVa50+l6YzFFwUDcMhXKCBuimg8Lk9jDeVN7M8DzUHkNE9bJW
LxiACwBbvfAov0okCq4iNXeBU1qlCJZyKGvXnhKu7Jgn/XBLtQDJ2J1tN9LNYK9x
cGLILxVyaLP32UVeZKBd4zrOmv+4Xbv+/hS1imF/tIK3rurNhEH/nkad+dAElq4m
j4UxTlczcjCpopMM9E3ZSfCRh0UvpT/YUv2X2SshOL5iDpbJc8D6aqP2Y818th7b
fSlitr9uRPymju0jG7xMzSRp73w8koDQw/H0x2gRtYRWbAQlelY6aG4oxaJ1TMjQ
IKPWQ91uf6D63Ts9GERnQxuHEro96Q6TqAU7rOY3/vtA0PmL1EGml5cRquDhP8yx
MZnITL832sS4Svv00dz/8QKvFr/gi/DiuyeGlBtIP1l8KjWelWNxTFco7ZE4MB8B
8nSgAcp+uQxiTcqXYXGQK2P4Qc0naznnEhNmV3Xj3Awg/tJK4/qxppFieaVQ4ots
2SXKuOoMwDebZf8daZeydKqZHXvJSJK66wOn//oLM5hm1+HX6Y/44QeLvztp6EgF
ab8l/h1hAWiSw5BwnRuX2iNaxwn0ff1d89fijbSAznGCUNg9cOnQkUyDKSvL0/1D
/Hamw+5cNX00qweIk7XU0NExU30sUiX3+f6dSDkhsZJ+R9QJ0qVTmTsDIyc7ylp8
J+Jo93oxeZ0R9fePtEmWDVB5G2HgTXZtwpvY8sZpr38wTloBlF2ODYblN/1fbN48
2MjXOerhDVQvOFKX7m4C3y5ngrrKuy+BzXjz3xxUMEIV35PjZOuMNzXYHNZ2fYu1
jYd+DgIVPuBexUQXmThZ4+bLTr3cEB0N47fuRYGmqInCyJKELHduYGi33j8d2884
xcetwRVlZG+ksdAI/cCMUcFPOxV1uITg15fEFH3CUUNIuliIKhz/4HQUXdcNHk3C
oCHSFbLpIKliELkh0h5i03WU2XWtRySzUHakosOjspRh9nhVkZXmfGQQjP3WGzbZ
5f2gmWNGExvDqB2pW7snoAgIDgZFIGoRf8UCqxiK/3t91DJe8K81LBxZjIqYfHsv
xPyYaKom8QLuVtjLVPhcwbnugHQ+y0uFBDkja0LxxvjbNIf2aFugoiOw3YZdu9dW
RzKs6pDyH3nugs994aa/f7QYU/rCDoi8IUZffHtr+zhrMu5KUJxbWBCVFY9ifpsD
Hah/ESmhJNZ+qxTjo/uCEDNLL89j9SlT6/epH6WD1yVrv62hYAdJcrAnytHV0BpC
a2hheMCU0cGsVbig5zMNod/GG2ylRlfeqVMHqMQnEiUCoMevSybhORiHJ4/K3Fqb
MjD9NCfWi3JTf3so9AD0B9P15Ok2q9wcohhbS7GirZnhPVvpcmm7Td4BBq05XGw3
8TWx7xGjfl8i4N6SSiYhwPdA9jubLhIScf6JfT5VW9ATIwBt0iYDg3BiPYApnafo
ff3ysujA71NXKMciJTkyoV51HtWQJRPVmS7MNSo/KxJy8ZJBjxC8bdMGv4dJRA+q
VQUH93o32FYiytYFYgTlQuvC7Sxh/p+6DGKI+f4gGwrZe3SJU4JSKGGa3nQBYKJg
QwFT131IRuPDjFf0jxqCASTCPn/Iwhw/nVOlbf7DJZeS2paLciDIbCLE4naBokv4
BXp1q8ImamNM0PT6WD6eRs8N+V5s0CDo7CMtMemER5kwXzFNDWIM03xt2x6THeXl
cN1YPoWN1ipX9bq1ZAYEQOdSdlydu/WmbV+jeKMmyBg1K1eht2YVjFEcZuG3tNH/
UpmGCi5Z++BexgSggQ426fBPqRP9j/4hnJ3KWskUKVVAR4jvZpqwI9bbPiDl8xN3
KvfsVDDbEiGxGfeLtGuJ7PinvUOEdyU1VE1FDJkk3baBTFRPXaJ9FdEY8uN+LmpQ
+tQGHJZFQGipsLz7ahL6nbS41fW38toFfqYVrQ/URbwrF/w5OvBebVPq19RlkMiD
SskHFtWu8Nbpu2atNsKITLE9mb/TG6Pzu7j4V/stFJ1L/iy4B8oW90nqVU2ZYgf2
CJcZHjvRi6dpFofaG1n8ASYMFBiAJJECi/mhuqEFFoDPLUuWRB410s5bS9w+9ESh
YIdZtVyuf12Kr96b1QL9KJ73zHJANt058LpDNqgiTvI4Dw801w3eLVsxwC0jVK68
2a9bEgIpoeruZY0E6ayvGHo9RZ38F4+6yd50uRBPhl1AXe6OGzRRleqXJHqdZXTY
Mf6+yp14k73Gnzkn9xxsT/m+zhBuZYzRZCU7GA2OdMvQixFMwUImcea6WpYfOFQB
+y77XWOz+OEhFEfKHaHj4dgAeALWiSc5KDciCsBurMFn5OvK30jPxuXudcRSoFES
FASU8jYnYbwfmUKqXg+60luyG9p7wdKYegSpcUbofOsZ4GyPK65hXVfzb6nUWzIT
AEarOVOxU1rVfU0aqC5MOk9MzxZbLhcznsSqfd79wcp7nc0JiOxiLnsEAUJ6w/hu
zEKumuKRD4i6WOISzjnuudh6XEIbvyi/waT39cUpiYfW1Uq+ApYU/TWps8A+zx77
W2O0UDgyEgmbkeGZiRGWkL6ukH7KJvEyldUL2VOvi+VziN7K5b1vj9Ez/siA839E
rub4qB4IbK/ydRoPye3bxZKV6JT4tnltEzBIcEP7CDFK4X6IOrQT6PAOgz2X73fG
LBhIiYpcmHTumowJ7JDubQVGtqbAbTYHSDYsxnkV399zcSbg9iMiFp2t1Euxqv1o
NWkF079/CpR+STcYS0EgAhpblHq/4tWeCWHXd30n8YKu73B0MJLoHcy2DDFpdTiI
2Sjo7/oE3YkPzetpSzZ4QkffMSC+CPkS0wBbJTmsSkwo6zbSCNREPDAcSSYSnp78
1ILxIiZcqQZLWMvoptL7RjCVJy9eKoPTqRSIF+pVFzWw/yVJ4sA0kIAYqDs4QAJR
EmS5E0+u0bqmyNpxw+D1BCIpGLm6LyzuENsBz3iznBVzj+F8rVcfMQdqwiGphbEC
J2kG0wr53/ByZNyZwxUcjHp72GCU6oORHKQX0c/1GUPAgYPwm4t2vZIRSm7QxS66
Jd7Qg+Gf2Z/Xk93sfJXdLB5yv7EzZfQ1taM/3jfLb42DOzMN1e5YEFSfXpAZWX4i
HSOrRRC9P1L2uqYSYnDwOQJnwKaG+12DLoNq4cJFZ2hd5gegxbr9n7vsBn8KO/DZ
RTYxaaKnNjL9NZWJuI5bQYsdrLGUNYBIPHqoMG5ntGt4Rh2veHV0U/7AWuKP5Pjs
591Cd5XY6SeYYuVneJ60SCoxuIz8JE2ZtSoxDlm1f7rdszWczWLlmfULlphNgeqK
gNAZMs6d0z6x8f9XRgkysuaMq9KL+LEb45ZuUJCIBi+8GYmP7Bq2bIuYFtDic79Y
QEZYgUs8dhRl0G9dKQnCxzaaYxAU1457wHl5sbScC1ELZzr43CDCX0dkFFQgUgLN
9F026NJ/3sX2WbyKX9H7NRDDF95RT0/+Ypl/s9Qtl4jSbVHUJT65gIj8KJEOyBWo
JiHNsDM3cvNTR9SEJuv8a8nNA+d2r/wjlKa/eGrJ1T9ADYRTphPE3xyWPAvauz+k
NUKdu9r9Sa8uZm+B5V98hHNqIihW4YH8IYPHK7wphZBWGWrpX18trWEFQCXFI1QB
LvH2Kr59nBzrOfaDeMR3vx8xOcGcPuELQcanVOs8azFAmat8mjhbmMs9MAs3Boi9
0Oaq+e/aP4XAwBSmtyd2NkvxMHxGCrEvuibH32FmZT7qimgYJ4czr+5TIN1xVRMS
sm8V/pS5qJ5qOuQx8fbU9yIuzXp7MbEp8IxgwXZz9Mlh5eieKTl0xzI2+pKy7IAS
K6GE/R5UhhFlEfodpfGOhRUdYwxAkBIgTnwr8C5Wyg4P20/arnBEWEUIrWLi6pMo
jNC3VARfALX/kDVIAsVY+wBj7ZokziLP/KGMzLxdnWL/bg1YKtV8eW4HyATBSRFd
jqVGfmKpgyu71Fiubx8J0S08a6hbieru4Po6Tz+pzsVgqOIURkmFKW2oXXyjZGYL
dBJqI7RgMmr9U1kl2PALKCOXS/lNtO62HzZf3hJ2EiYkvkUMR+2RdR1NQyl22UCR
a4tBlpArpAy+avPJVMYhLj4kbUK3r2CKbr9JpgABXg3OyRuikTDDhBCHvG5aVpb6
ZFeJ3ynwGUevfE3k+mvC5K76/V7tvZJrmwE8GNX+Y4BEPnrlrbxltrrakC/0CX5E
8m8BT//sx7V1FU0ZTk7KG/j9BwNsi25kTtV2Kq859y237v8pebH99fccLhQGmRVc
15d1V60IHdegMr9l8bvVoTtXXHNXpcF9+M83PF4TyKHlZO3EQbSDw3gXnHN+4Fa3
RXdfA9lKF2DloDu8bRnKW96heTWGm9Hf0t4q2yZU/vuuAWjXoS5PnErnIWv+WlrK
JGW0sTHiB+lK9JDWFJYx+gaLi/KfOyNRGizGlAWNzR8lVYMZsyRi0D3it44IclyT
oCM5Dy9Icwm0Ef92n90IyNL1r4FX4EZU85L5fkNj7y12LtG7kM2bytDkxX2ATcru
N+QpbQ75vuJOZaFhqVwOAT+G4IWlUl2QHekF3WilnEK1T2RnBOjlRof9+G/L+xzr
f6qxj6x0q602nrZWmN1zDxWKoGp6WC09zMqp6zYl3Y4G+FSCugzwtw1ozgf680K0
iRFoEadponEybjex2D0LKyOa983rEFx7eUZInTIrn73QDiUDXTjOu/QRrCobko0d
L2y8ZWKwIBh0PfyRpjADv01TVgcs6F2CLz/fE0n+kRipFs0E8efEu4uskbbRzIv1
MyrB+dQvBRF0WSHdKEEOEFM9Qh5O1cXJ2y5GbJ2teBqKDZ/hEvPMqUgYLE15rYuv
Uv4qYgl2Nbql4TU8d4pzrarQkeangvQUH3Th+UtB3KuuivWAHFiZtKPnOQkN/LIq
HAMvZjb8KNhPJRv5LL5XHQElCd6SM1OwrLy//o6BMXJhFRnGE8jR7x7jBP90SetP
sr4BqxrAvroh0u0rjkrT/pzvdCLMxUhrcQ3b7qFwCNKGggAJNTZ2qXcf9NwskDm+
BsEaanOqQO61uVgt25OGrPBV2PmrkC5D8sgU+yvbcrADJv4wusOgzKokJnab5o/l
4MFGkMu7Z+Gh2mYfGvLLZSvfJHCrus4EoJ9sEG/L0A2ggJShWxZH2GwdbC2ZALza
3SdO2AvihilzrwwLu58wBa/YW6YgdQzH14E05Oyr+khVUpfFMJKt3o89Ohqs1K4E
fI2B1tR1JyadupJM8WYzjNUAeBsAUwd3A3OBf4sfrjLcS8AA2Hya43PgGvOtDi66
6y7R0IO8dz+pE1aMNl7EOFIpTGlyp64R5dg3b57m0FiyjSzmLZQpU/30n9Ua6+Rh
MSgLBgb5vaNTzRQ1qcZFSyw17ZEAUayLYZMfyuar5Kh3gOfMleqzctp0vngZdbMd
Zu8wU8IZSD3CdLnhhh9truh0qW0zwTp51xOgq1GQk8WambmJFjFvRIVUS81lNFpt
X56GlG/EtUsGcoQ5DvISYs55CblSMi7ex8b7ra2Jx2iDD1akyPBlqYlUn4q6UJWv
Gh3eM0Iiv8XkidoVq9JOJ44aKNPQpbM1ymnF81HNfgZnmaM9TBlD0a/ppc67KWv9
xWMxfId4APqsxd1H5H23zVdpNp31wG2Z8Z7tAS0xhY0HvHR3gJMxrSRd1YV0XJ8O
H2Ma3SBP/l/MK0xPGpSpGyW5MDzlmMfzgk12Gelt6CY8x9uWuXjz9S/sgGFJ0EdN
kc8fkvQ9yx3YDUKg1Ahm6UaYQwI3zCPTOd4qWa2hFRWBZ91fFQoHY3AsLgL+fpXH
ClkKiISNhHqsyaOgvRAzL5eALl6+iRaAlei8axkVluhQLThlgKIwfMSUt+zTc2eI
B/N0ODClyVuA5S0x5oKmnlGBc9AoOuCq24mT21jPVhqStFuvhydk4R87rLJJKN79
itEFHz5yEZUn68aEOtKc6F9wVM91mMIBT7rRXaDK19Vmv+h3mnMw4FpKdNqZ1hiy
ys5MDsW3NUgDNodkCyzljGc2V49A7FS0BgawoJpyq9AG9WN9x8S8tG6jd7drjkb7
Or2x1AFI9HGoUJ/B9G1wIMotzyneiJMSrQLxAQlQowdIq06VB0Rx7+jtQWOQCgmv
rEkJ3kSTJ2r82nmVTxiNzRY6nfcf1O2rpC2frSp3xuwDfh1kEVYjVU3ngqJbeY4g
riFEJC7sqTOigOtZR5bMqvSGqapFN8YKNHLJb1U+UzwwZkdVG1JJNOuRdnuu3ZzX
fgT7g/SDFx7Bp6UsuQv1hPiC2N5xkSCmqhIMFLdQvnyV6nfSfK1pCjDGo0OZj0Rd
UHEk4PrF8/0HeWWt1fXysCOjSvc69TLNRO2CDdzcZHkmxc61IWbDsLQhyLzmWcl/
7D1xYNqEb2uSECWpKMc1dJ/gZn6fHRd4vR1K2KRQhMDxVFFX7Ni0TtsSQ/O447FR
EqpFf161mr6cmggImwrpZwVpRAKR8BQ67Oaelbl4yce04bY0W5U6lAKw05W3BKhJ
/4bmbQh2CE3kxrApVGg/eVf08bbSLBHZxTjv+w4OqmGd5qnGmQntpM8IMnmzwsbU
Ip3t8t7jkCJwe7U6pQCUDyrCQ+QYO0tCjO91Sf0oeIuNxwWom+DujqL+F37RoX3L
hn/FUI7FzPgiIQaTc5bjZ7veUJrlRuoh8Rihvg5kzO8ra0uj+81WToM8ZrVLB5nt
xrBnoQZQmHMZ6JsudYgcHMpna3mQEyGX9vSmp0WI+b+rPwxk7nVBpAnum38jnGUL
ncbYQLvkWrQR0H2ASpvxGXadhloFPzZuv2xXv/3lXDmiubvcPcbN7RQjs27/XzsC
6NEzSXHzW5n9BPG7OzuxROianOhpPLbTZpOn2zHUfmNpo8waHb1EvCkmsoDvMi1D
YEMJ4Ytc5qBdjsnr6azAwFL9QU0RcHj42FGt5a/1aBeVc0RtvRCDsIBH3IUxxG/I
y9vxMYd1JeF6O83oCtiutiCuknhtJNTbj+nd1Elr+M7s/oLkFp6Z9KiPGJZQFdqK
FEqX1nDu63PUDBRhkOZQ/0XeVnYSmzZhF2brvuPhDDmK9nHZTZ8CY8cy3d0mkRad
mBZ20K14FskFVaCq72Q9j2iMkgjj4jJZuQsN19KqP5+XEfsevb0zFC9YWk0Crsqs
982QF6m2M7cCfKrUVRrRMloPv1v/V6SPoOj07+iWOmwUUeDJF/APxlk6V4HoUb1J
GLG4qw7NJqe9cC5ld7kd04O/orNUQVUFGxrD2ilMoy/KoJaqp42yH9DysD5Krwpy
3yZYUFwFgJ0gYnjScZPvSYTwc4d9FWCS5TdDmsA6Er/lZTdfKWaLCMgknnwRoB4n
Eueo+MkbfGKTj7r4NEsRegpwvQ6DPdP8akDMKFBYUgkQtZ1OeKYBlX3vSauByMY3
PdFvi4mrxDD/oFiCIfrB4eIkjvqRvqdm3y0yUwUnPOoahOZDz0mC1Y76S6dH0vsZ
h/TsWLmyPk52/oZXIK5brFkriHo9p7CphDTOuPenJOy2vfOS7E0pOJTAeNvL9rOC
H5dwz4xFvKrADdylb4R1OSQqF/sa5Dm6TYpsLlO+AiAso0DOqXwKz6K7SRCKVn8F
7md0ctjxcIV1p1C0fN8XmhGLbHubL1Sylm7rcHJsIs3BucixAI45sT/DxDRVB6Ry
crjZKlK+N6Ei0jLJRQ8H47s24USNQZICMI1jQuwBDl1o4GtgllTIi5AfMy3AMTPf
MruE/s1cswQVo36SQ6u8L8AhZJUKT8JRMiowbMfU2sNtPWX8IeydDGVGzJyp8fPW
lT83j9oWtrYUo8pXbyuHxQcr+4uxTWpJT69o81dRkse9nYjY0wC/eRqyjYN84FZN
/PVQksUtl5068QTPkbeECu8dadXLE+oKmsG3abCxCHwW5hYWdiI2ResbWosBjnMN
CoMBhv+lS2C1flnGCa26qEKPOshz1R/Bcc5OjVrmieqhIgHjajAMaa2b9X6jahwj
t1Rxw0lZYvtiR1HsGC34Y+Vve2uM8gEwB5zccV05JiY88mX49ysejMiMlOc9hh1P
Tfh5s0wytpBlmUJpzDVCmWk2ckaU9A0KhIcWmodXR4E1jD4jdQGdqFa7+tMatHO+
YAJbq9Txhf/aRSyvPEg3o/KP29aqWSMdNmkJMm7UW0BHsbQmnlqKgQDp4gjJFSCj
E2db9Jruu/OGxJra7PCoOh+HwyshYxabmWG1rL+8ei9ANvXItoCR6XABYDPd+CMm
qjBr+JPsfrcJK2GKZX2iANGZS3TtbOMbpRMmj1eqE27Qt+kLn9Ie9WedB+PpMGqh
DU1mTLroTy8YEreikBi98QoEdOvfsQpcAnqSHcxgWLuYs63BccA2M4jd3MQ6YXRG
lr13iQuQJRAF/RiLKhcjUiuQLRS9mWdNH2FH38DLgiGXTWn8h/Foymw3l5bjoGgU
yuc33XphFMIJW7EFyiSeKBH837TPSPh5OBZPsOMhCjM9rbUqHwzgcq5lUz3BPbb4
gDsw/Y6sVcu2sPHxpstTUbxcmBKWEoJSLrtD0VBky86Wvs8/BjpsERJdTQp528Pp
0UwaKlewWDIGMwvIYy89S+ms0MP0cjuF6/K+Db0Wlp30TFtKsehYOuSYJrJZqwfT
7lAe8ljeBCkx8yTEu0MCYCHAkL33FcT7hPj8SitaVacYYYyBXJkD0MiJ0ht1YpnX
CvU5P20vKmahPmoEJLKLDyVmL+sGjJe4xnNEnLOwoN4Y814XkkC6RLCRpV0ANRXC
oCtYNYphSs10sEgtg+L8mGUOVQzQC5YUcsnnLeAPU6qaaW8fcHOt6TJMW3wUqKTJ
XCFqNzJSAMIQq8IfXbxIvyy4ZflmSfSeKevVJZ4ZH3EpObFkK4BGHWk92ZbX1WcN
FG8HqvPkr8QdKO+vkxSbAG5k1yIERrvXCGXeqqR5yc+G1wA+1/B2uJekXIU6EUvf
bMk61H4Jf87HFDqWosqf1TeUWE7YANCtxHxcDl25TWhehij2cvOt77KdGKkz2FVo
R+o5IRSbCySZAZIEaDs0y3G/3Hml+opFgnwN57y/yT4XeCGGa1Naeb9NuF0/t8Z2
y8J9Yr/0UMIPYtzCxtB+ADGEMTuOYU9r5pNXJFQFtHShGJMc7ewIdzYbmf59Y2bo
JFT3MrHLe1DEyYTVIN0eSzJw9SP/I0NICNdlafH6vDjoRaIBofLTLbSywq22Uwzc
s6orNkV1KO/Ycp46wNoJ3O6Q268YzQ/4k6WrjqR0KKbxJ2TQNXhhMstvBT1vuVtE
S2cE/FJvBB/4pjrhYrt120YjXNE1ak22RUicKUrkebHneY0HeQN6E7vz6uucaj1B
LxooL2zxTQjdWZqE56MZu6EZUMpyr28nugSRPTdIEy4QrsdQkSgtU2jdAwMbgI80
vLGxfiej9WNJPHeZQQceJjehg8Hq0QNIxx+IspvsB2QkRuD1jIfdQHhpYRCGOhPd
t8ifqd6PNsHbG2Xgc91FzuIjglCzJopcoWj+Wpqo6Z19nM8j+I5pEsV6VnbPi51d
5plXIe9c+PQZmv2ihgpCv/w0zcGXEVQu6AbBXjmwbuKUH6cAlPbMwQ4gJBPHS0LX
92Zwwo8X1WofsJcXQPZcmavOD2/pKYfjjOAmLHXnI/oU3M+6ZWaV5Ygu+xsnxNTZ
3mMAycGIoX78gv8lvXLeCagbMblYIYcYqzoo8JWDb3Xm7LGmIDpqsntNBRJ9tfXO
xNHpm1DJ3NMip81sR3U46Q0d7XLIu6BO3dHvZa8Kg7QUF5CZ271wguIeLd+dnxgV
1bcEOl2PR9ZCGstmPTh0loQg9zg0bBfh0PNYjUiAVzgnePaASZlJc53gLW5PqC78
wCpq6VDW2TC0dm3QM8UW37ESi84GfFXzUudNeCppwUhxcUzZVW9G7u4r0o1HkA95
0R5c5jgX7246qCVSxLGfdPzcBaOx1LjmDnlWxeouLcvBOiBDSnhWfE941OrZPzO2
QcYTmoBfdZg44en/tI9DCmxVjCV6sGYSLVmV3yyv7TgYwmslEBfxW2WOpl0uVV4e
GA+JH6SdRjYXvgDUdmGzVf56eCnt94xdUQgsv5A5wfLBRlqqjZ1iSwkJqcs0uvGn
8dLe+V8eabyKvnp6lgi6D0xFtwiHRIf9KfeT3BGhZGNmQXhX+AoV64RGcUlCAmNF
llesZ6Oz4X/7K5U11WluYRfiy/ykZIjvvdBVGIxiGmd2ePnucXEUCx5P1QBkvIfT
8Dn4DrI2iN7i6OSh2Va1nGGJGwpESL1M7JV5uts8IA4CkkjZKmfVLl7aSKVcC8io
TWuoxc7+HzSKzzRaf56Amo3YcjNLLp4qORaZyU1IrIgSZKsPFjGeVPRkroAGqFWZ
noqfYwhvEpdNk5LPtL8WAewk/87j7q6kaeWeEZ5g1BqZ5cgNR3ojWntoe1dFIZoS
FBAmK6u/fM+97mtJq7w1gUtF9uAe48pH7EoGY+3BD2mXIfCxVYH7t01jyTp/NuI6
fRZTf9ZGXC8+UUrjqEa1ET4Ol3uXa3EvliYqYNMYtvpljgRmnuU2xPNtLqnbYQk3
mzPOEm3VhU0A6k457UfQe/FaT+i6q3SGbJF1tBKF9/Mqjs7elllMkM35zqrurIeT
dsF8KalGvyBOStb9FSJ36H1IFNqG16JxStPaWPgjh8a4r/Qdaaea54J3fpZ0DTIh
liCTvkJk0HDfzUnmUDNwV494SrS852vhBmtbDSTYFCgv8ifOPkfwxrjVxBMH9jQy
ComuFJl/dhv5YbwnX6BGi42jSn28pKu2A4MdLaLy91dActh8XOYKfCwGKlLARtaH
CuSzt6OsrJX1B1KdNUfl516P6e8EWlB2qUngcmrgyqsxvmQCIgdjm0nuXpdgPaT4
wpbspVjoutPya2XhwLjB7AD+2ekKaSzaC5O46uaHtge/ZhmL1pdHxt2CIYjMHHnv
S+SMzH1l5BvRgMWRMr2oxoowfEficV7hlzddAbYDqlLshcQxDlbRTVCZMTV8rkwa
jV3WNA8VBR5B3C7qbslmei843wWUVnJ1wn5Tyh9dEzigstc3yRWUDUL4XQ9bGlqw
IgT+3APs7NiwxsRt3Yo2+Luu5JK6aADDGFfl6LFfbuIaxE0nN2ta36+4mKs5WaZT
HL3e5KlcJ9vWTkzf/xtbAMYKsxS2Q7Z7o2lxHtJIE6ZSimQi+ok1EU/jas9JpfOp
4BDLfNS91Tq+K8ETzxJL+KnBTY5BvirmO/res6kFvRN5yhequDIbxDFUgU9wmEQd
I3vlcTASsWM+s4iEmcYxftW5irwNkq1ZVHiFjSetnSO5PsQolho1gVxzPCKtFJ9N
hdgv6VS4Cw48LtXdITdZ4n5hdIJpcwaJiU9IWezxtjkevCBdH1gurxIVoq5lYgM5
bx92WIyMPTTDt9ntsiWVMgRz2751klCQlDWcENHIfOqnB3N/tLZS+WGTuPWcV2Qt
pQEWYh12JsamZNjsBnizGgJKCDLai6+0EvIE6+V0MSZM5fhj2ufkvNN6XWmQ0V+Y
FFpd4dj/tkH9rV9IAFNJPKMN33Jjj8udqFyaaAZ03YArl1fwrh+Rv4dR3LfwiEK+
iDwy2lhTugwaVB89ZW6p7GH3NAcwl+f64OqhHzD1RcwbF/dRDZkU3dMfX9dzcU3+
JuN8G2o92PrTkEpaxsdvTUkebQ58LwdPrRaG3h3hrNUB/hnZ3+Q29mI+Yxvaib1y
wEOaZZpiKbWeiz7VwbRYHXHQp8/rSCw3uPc8F5ggPCW6kzFOcUayDpJpU1t+E1CC
U3sZjmrqvE0AHfOWileoQnV89IQh5ydTk5KYXPuISv2MyQLBTEbCddgfG/MyHRRl
3+q7m3EyUDMOnD6E6duVAiSiApZljR51s1kF0URgaOCH3gX3hJqaFCrtagPJnWjv
oTD/GrdOKWHzPH8WPXFFqNU2n/eMfGneOBZ8mECUiEvg/Hrby1LugSvafnJa7VzM
ikNm/OApo6FywFBTPDPxyovgK0fu1sDl/iLfe0uQiS6tuLwx2oVdZV/ecbS/D8p1
MDmmeNmuTnz7O+m5BupKIfb7X8aRLFJNsKdMZ1r0mUu6sXifWfZ527SML3ksadUq
vaW3Gcg701tEDJyEoTwCqUGGGeEqrcPnXt5SImi6J98u7qEsCBVwyHdbmUOhXtaE
WCej7EpgLd2GsW0tdi5Becgan86udD+SuGBKdngpHJOiG/Xhnz4GgKsY3uHsfu2u
LtLwEXL6TVG269T+HJwF2hRORIoe9kb5gkKP78fnxuh70McmnhliwXnL+FFKP2s/
tm8XZbS8BwESaNj4YAhJIBnKoVF2iMqqXAS2USZk6mKUGgkbqmt+gLsU2N9APFCX
J4oRMPcC9TbVfwwQewdPnfPvwScFJeh2HGl+U0TnvWvYxMw57bnjDUjljvOytxxp
+EvxQcRsZBgNzC1/1gUp7PMmBWE/pI03up/VW8vC5hZD1S7qbRimODShYVY+z3Za
xlgEoetkRw8FXtQ5sURinkJI8z7NVwMtev+KsMiaRydUFJGDiIYKLLFgQaFga1b5
d2U4P0n/H4yy4bkYt5L6uvBHFFJQAXA8z6zcwsYfqIXJVGm5ln2DVohuVy0Xxaxv
PlcT44Qk9CW8SWJc0JiEXDX5MVxSka33XYt7FuDAPW1L+h4+xmFz1mmxZa/okmqp
B86r3mRjipcCRf1+cx8sbl9Hg4jhs7BrhxmbBlffX5H2orbPdK2H/4Gf26VSEcJr
ag/HTeqRGCe6PRKWTt+T8Ey6aW7RLwT9Yae4x3LETA+YMQfiJnoSIJllT2XRQpwC
4+zJ+imrqBiEJORO2l0dNE7ICssqFw8CeG4tHw9tQWWUezmqZ0u6GhGh/UdBV+7i
uOrZPBKNn+8rlMyJU21ePVkRsEEnTy7QFEsUyFOXO1fUCHz9dTYFNQO8oIiMmEJa
/R6vsuVKHplkCa/1fiJ6PAIAme/OQdBU0SHbr7CGvO+3ILm5YBgzbc4lBWLRkhwK
sM9N03u0VKOyj/jRnXaKGF11nyzzC9KbF39yuhMmYEcAzDKlmWFZ1Xp20SirBhoy
DLSxkpIz/h5Mzf+gSUtczZF3vSRyFogN+JvNUkgPazHUwBhH/GomqcmYyBE8gZWP
P+Ul2OvJ45Tn65C7WZYJfULP/0eI+QhOmmv5OvXzfGEAE2ARaAeLUzv8Rmg9SDko
WYQh8XUkG6bmsYxMrrY/tkNDSgWpWJ5nWqCptiXkL+pscWiyXal1v2WVc2F+Uq5o
ZwiMVY8ZLEiQ9gTvwtyFFWzGkPm8iq3kX1CSGdmj5N24RaR27psJ15R+u6ABghOb
PmLmp7XrJFcUOM+CyzWTkcWXRFqF9EDrIPDIyW+B7PGEcdGbF7Bdi41dr/IACltT
vZ6ZHI1ocQOeP4wpBMiP2aNI0AjCfnU+ZEccGcF2a6+VsAtPmXiIHEv0wx39b0Jo
SjV26i4RT/CrNLYCQ89JRmrfZwZvMzNQX475KXTlOl5+Lr9aJiuMrQiyi5SBggyq
fzjjd/NxH9HCgLDzPwP6IG/sJhKQHdbCcYOLwCweMufqpSi5Vv37PdodLVZm8ZH/
qrnUZNhHt1USecfAPW/v+HCOvg0FW0IO+iYpPqVLfxekC8vvw+ysR6yibQAqvwgF
t8l2GilqpJ7mdi/gT8V8Sx8t1kmTMwbRBzR1ju+mRagtFJzIHOOW/DVqcIhYP0gc
eMszXbxgw+EJgyXmzRHSsocWFzCbVYp2jVjod27Oh1c/hW6Ev//4ai7znsPqyry3
+uF19GCbXBa8vH3n/UYaT/FG5CX5ySH+ndCWhUMTTKWyy9Cezl6cSQJHxKl2jzdr
3IHRnrKmVdX0wNWujxUvdsle62Z1SoaZG65nSUDD+dCba0WTM8hqLVmG7ocVoSvn
Ahva0hm8Iy5Bnzvyu80vUqEeVHK18uKmZI+1eupsbGs3KK5NxgiIGSMJJ38Gh7hk
uijPNiC1X4qfyCA3jRIyDYzktavZ5sR8XAD6Wjj8DOUncUu/ZBKmFozzV3ClxbfC
aalPZN4JkEeuS7X2r5m96SblXe2OsMeB1tLxSx8YD3p8D7VODEDnSZRuOuE16kPi
BCDoTXYJPVRrSoe+NCQdkQqEQ0oDopI8K1Lz39f8xtCvAByFHDWpxR8c52pYQ+ZI
sH8B98eV5S9cIWEst52QHzqoULRjzEYSTZsYQcOXTbDb92AWGlgHp75o3Xi3jUCh
uos4RleyPxLxLPd/KTp6v1ixq5X7X35MkSafF7mYPsEbgoPpBXtW8QAi1SJ6zm9O
keZa9j93lfrioUFyKGuB8xQk0oGzddHKeloWhVPzUugvmQfppiYMYHI4sv3zVcKD
nlscgIH3iMA0j60fkRFZ9dD3cDvwa+4gvZRAZ6wkMefnHsqkWmWq7EH0cs67PTD5
slMZuWkXgNidSdHTSREZJH31fJkH0G4UeeKuPLfNgOAFoRT3lJk3fpdwmrYG46Ma
XkH4XBcyfXygjQe0QtblkMG1vnuTcHqO8fGtR+vBcRNqxIObevQbn87LmR2Z0b8c
IHFKxhnCaGy29mKdIeArWDg6IzT/h1TYJa/O15i2b2i5Z/Mj9/s5Wd9JxcQh+Qi6
osOSXVK9emzGSwOwohdghLxkVeSjGPsWaLAAMMT0DTNEE880E79NNv14jM9ouvHn
28METdJnsa6mRC5RgYMmuRys2wwWWJ0II2jwI2oh2DwsXcRgbnpGuRQ1Fkrzo8b5
BmbXJaW8T0xDCKuoivd2l98nfisEzDLZRpBHZljpdU+TdkLifFzg+51W3S/IHic2
m0ZqeIX2BFxJWXDmPlROOIDChIcIXFsvI5lAWOsYrfmFZqGHi9tIDQndOn+ws0LP
LoO/sEEekg7ja6CCFouTwMFOH69Ydj9EuugATir/08zOCHG/g+JdgevqRFcV/Z0w
fsr/IPfiF9ZEJoZoFK6F/8PgCQLNCucFbYWwevQOthY7+lN3trOOzuACqIC9Zlac
3eAJlVtHAagMnC4XuWhvaESZ9TredUpPiyWlT24jyFlPG3Pgcnab3xh748g/gExx
flU4mBDooIhB7Clv6iJh2xsYAQiNgVdk803NSS0OHSjsFAbRcMcgx4hC4/2GxWAG
dKE4lmJeZ+79qy+aUFH166ctArcTIUW1CIP69O5TiQg1HvKEHuRsEwJ7u2RcQW5z
r6z6npCawJDy68SheFXMQyFGyQ8C+ysHLBBV2fHP4bUy3Y5OMqUu+u3mc3I4p5+m
IjmtNejGBxp5dW0d9qss8e8qFfXHgCG9uwzM2h6h/GZoWROeDvveSFXVrnUc1D7d
Kago1aPEmDPOdQLUcTdBfg//Ju5jcLM6tdUKmzAgOCAWEKwctm4scYkgkCVRNQiN
B50e4J7e3zgQA4L1jbQEoG2PkFqfXIfmmVBbC9xgRppC5u1pV5H1fSbXKkESsKPB
KOJElyWLTRGM0AXjrXVhdsDzzntiYDJqj+SsFsyqmSDwp+6l4HZUGZJ/Pexg1g2P
I5A/6AYxV+XYxjJHJMNNvimf3tUfdciJfluCyDzRI1Y0aJJ0M9Q9Qy5G8fQYGPr6
9LM3QxQvRsj3609u7VsZhhwQqyTpcwt52637/gfJHahFvibErV2y98Z7t0FLfGnA
gqE9SvBixKm4lmrANqy8tyzt9PxnmahDM5J9AC6OzwPVczyIfDOsSpHC4+ROdsVw
dFjQULtGz8WXEUZ4mn2RZ1cjlV8Pab25HZdO7Rnwx5T0r5dMg1uqdrVf1AY53gnW
E1p0rANnnRRfJITDhSeRvLJLobEghXT5MDcrcvsrogCjdjF3D+iMgB3EnggvGlqA
4dTVR60VtDGxo/qwwjMH35S5091VyUeHAKW+dCe0EQVHamUrpareV2r730JlTZ14
lec2aloR4IqcHUv8XgAHKwUDslOTokQ0IhBYDVyHpGGbKCl4HBo4aSO4SKzioCqV
PqYLhNnGIU/W9tQ9Kn2sr//fCxw/unXSOxbYAJPqn4zIpWac+x9ZwvZOr5kc/caf
vQdzGlqB0aRQSjDcwDDx6rclpR8wFktd39zQJNQcHSR4zjtqL4DYQxargwmF10lE
hnJX98/65ugzF+kAPsZxWAnxeM5eU9yaUBC9CSfnIeYz7lWrix3jj3EwNAsjFMiT
1NyhDviLE4ddBgyeHikRcWVfslFsdiw2aPPyUP5Zxf7pa4szXgqKJrPFuycjnKCT
pcP2mreqtOylr3YqPlXwdgR//JyXcp2iaOu1J3HcdLkoPVVE8wkFVAnLklti2xJh
J8BREYG3/o6dH+I76zRuPeXji6QdX8cyj1L0+aLUn23pOLdAxwWzMEqEYfteePA0
r6/APyA4Ceix7McvNmCITocdDA9TeW4ZyCDDgaMRBxzfONx6qK6Izu1wE5xWPPLf
t+xQbbCzcatVo6iK5JXyGYqdFElRltQ6+PmFVZvoVgGLz1BAbCfgAXQZF1zBGnEo
TqAk/V19cj/Y88OlSnsZWJfprOPWKO3L61obHHvgjezm9pinbjGUKjb1FcqSvbQF
fyaXhOKKItp9hejxdie9iXKWiufKzI/Bg+mbh4qn/tRFeKqswcCnnPvoY1LqqKux
HaCcOFrfbVIOs7GWvfzIagu9DTdi20RauT9deLNlAXMGfdAN06tjAPpjgf+kJOjp
Go9lCiBA8fpPAF47mUee4v77jcUgl++7xq/SD9oSxikBGFSPEjhSkQpgUqQ/qFpC
OAKplgbiPMysZgHOubWNaVFEm2pTzDyDhawJN544l1zK1emfkrs5yIYUaueMpiQf
RDCAthrLiUWx+UKcdFGxPymuuNumGVqdBS8BvObVDmGCMeReX85pQAqZDJUVxcoP
VgrlsZcRJSCKsAZVzYZL7HvyQYMWCJpauXFAzDmhSL+a6bYi5x58kOI/j+J9xhLV
XGFXRosaCdPM5I+jCJRENVcZ6L2a9TKYpV/mHJjXKhal1xkgQgq2qlhKxURMHhzf
bJOicUagCbSyUyyit/yPXh0TvyWVZvev68dQhA+R70KQvcVOXae8jHU4pdC+52+F
RzTCd/0NJRNhIkbtBd23UmA9UYFx3B5+Spna4qoddc5JNjhzs0odGCI0pHHigUuf
ePQ2ilDVOh0xr1OeO5dN7/02RepgxVb8LTlwVUYrgSFMA3uh3T2ZizltlrCzrXbF
5tjmYjUgW2Z9Lo1qiJYPI0KmMl6IqIA7IbZDMxXRkVrWSJKhk92zS3+/Mupmus+J
onCFBPnnacYuCiz6TmooJdq++HL3OoHa9f9BRvM+7vNMbMz+D8XEBIVnBUKkPu5J
ksQOJjscI5PSCUE6xbQjR44rpCc6Lsszh0wOdCt+fPoxJQ09yNdS6rUEenOV24kF
ki8Oko2nEYaYi7sVECn6fLgBtwsusAmJteU6u7gGYOjGdPBwb9tQ217pP0wUReTS
RFX6xON4okfZq4aIadDC1VmJFAZ2J6ntANeEzD8pOM+8aW4KwfVbMkEu/zwgSLVQ
vanQpT8vxb4NexhPwppivgN8Nxd1B2dql6nhTSTWLMqfmsXRUEvT2eH61KC2eKcx
3mimuUHxyUIo2XagLvfQQeLlRXIoHKSzNhLnsvpqO8YpU01iMI5tK5cGzBjm7Mre
nLLhykQMLmmA7WFDjX8udl1UFZyYCHbgRWc6e3UMdMAMEhQf/iyyapnyh2sfLZTB
ycCTD6/ijwbAS9bEUyWP3Mxmf3hXrZKlRe2//IMKq8RpkYEEUHEEp04ETLqMgLXs
1Zf+sYaNtDLLotwZyPtxhYWcGu0y6suDgSnY/mdKaQHoI1x7akhwVGpV6jeD8AsL
9rjxoW5YGIGG7FHAlkjnptVVVwxsyd1pf6kazfB26tlNsDyyLh4z0qH1kr0AQ7tG
dGTnD07EkebYxkS2DWGw7zq9emDfWQe2GAKV13ed6aa0/FCic3piQ3WFhofOOHa9
owr39wN+VBamBf7/43Lqo4yM7F5891eJRBBf0jPddoMSNm2fDw3dN+lRUMVLwZVH
Zkij0kDul45dKATV6gtwWMsyKKZAc9R2Fn1taNba8denvmeCaGzoBbS7kEtJlP3Z
x10UIe5hBGED/f9EygRarq5Fe42nOFR4A6kNAeG9hJBT034OmO/MUeUQm9b2f/GW
tLucN0Qwq3LzUXsK5+4v9vah5mTIs7WRN67IQEmcoNHoLT4n5RTWTv1OcpVIUAyS
q66OyJH9Yy+hR8PJqq9W/CCK74C1iGOfb3PTRSWIKNwVDSfGDP23zJGGo4kGSgLj
6w36VBD56Adit3PDwsoJImjYEQBYKg5gaC7t1u5ZWfTimeX1hIBVa2swgMu16bvH
UYRlnF8jiwSDLj9C1M+UCF+XnJSIgv/fJFgWM3yiGc0Ei8FtVz5yuuVpuDubkXC9
Q2WJ5R1qzAq/3g7xLnXL7Oj3Fh4eSdRi3GoKpI4r3cop2ACW2e9ewLlewfadHfMd
7qBACvWejBNl2wynhdNuZK/fnKEnIvzorVdmt5GvCXrX2GQFctRk7SQiFzXNRavV
zox8rC+VglaKA/qigKuElSk97UND2CbEtHMJC/hUOHCo0jsM6AiIwmsnMDfSjNKh
Cgf16uy0OkQ69DTtD+isoPZwzwtmRpjBo8kozqs3JDiPNSI1AqPmQLKJFsfMBquI
zi5m8hjiEfpGXRQZWj2m/ImpbfzQF6wWP95xUBQ3PEkTK8VPte6XZhMN2vKGBiOU
kqjNDEJptjrRc1CdDRxGJtk54AERy08Sx5vehPwoIXI+H7q7GaPRgLU/BFjFZtvj
cAYuto6Xrf4lMQLakJlpsHSefOzkHvd1qB1glFEZBvQCt/Bu8zr82mU7w5Cs/5nn
9SFFyHP76aockP/BzS0IgXZ8OyrfwVtSmCSJkReB8ixBYX2I9Y3EKnLx/OaO3sBs
AIFDIpJTfAHPMqtHWsRZfdNM0dKLxx7ROQ6hyQc4TWdywO2owF8WveXOScTr7+rw
0OFVoZAP5voniyEaqB5T6ZFgZTdHAZP8/dcgAVZ+rd6t42ObUtOg7U9Fmopma1iV
d7NAzx9fT2yF+1F4EK4xKDLBwtKlKThCM6zoziZhV8PcFN/HhZsbjBYCiu54nmCo
/QE5ImOFecDGvGQiu4I8eipL+KHZ8RfznkRzVlOO1ckkhG05o5riWzKBdF+n/3qP
+SkXU728bb6kAPykL08BASAzXlnUKRfiJt4Lq6Jtdtu0mc9P7BBTBj61BEhwwjsd
SdI3yBnm8+xYAjWK5exHpGAqOfzoJthQLuRYRrVqv5nbSyXvCsqV/FLK/Y5IvBlL
UCDLhNCLEfU0GusxySDNuS1ze8iadu2hekPUS26YWrxl+Me6HT/NdKP8+vym4dW1
KMANy6ctct9BsoDWcSa1L4vm3Htb0JwNQzqF1+aXInu/Zf0EpmdCNJejekVrlJWt
MZ3HB3ij6kCYuCiG3o1XMA+6imx+jYVM3A/ZcLNB0M2ybREG1iUVvtasLvBxpxzk
NnsjgSZCDP9m3VIracQuWuPXGiCyICD+KLEPNwdb8xrwW0caFrQqui7AtcY+o5GX
Ywt+fhtsfEdhTi+4XuVEkfWFfCjvqhIAFK8jZz2S+VCz6I8U4IK44H1hXHAFOqDR
gZpw0gAiw3Bt3b08acB29jdVeed+6PnBjvlsm4bY65t4oNuct0CRDyqwmnXZvn4/
079BfRy+wF4G6bmFHOzPq8mtXML+HoOPFTZyGMNKpQwALl6NFwEkO66sSMbPSLHM
m+0Kx4MZbbstEv18W8MS11jGxsDpVNi49K1l7FBJdeQ21dNOUXp68ysSVDAGfBCJ
KUYpBfeGr7a+YY6l8mygWFOMBMsiO22/7uaAjDN736Gq4Cc3g0KzW77deL5DDHWP
1JSIKnOcIJvLEeKQID5YwZLjr1cGGm+6v2sfvfz/t9+qFpFraLxf5uDSWiShWYEz
oXWrOdMgfX5aTo0XoYKxmERUj4WwzwPqVcr6xG93kldiJ2UAA+R/yEhnrS3E5A9n
XKWgt2GTFaPxcTT+cF0iqkLNqYImZnOKnBEVpXyfcPlkfML0sk321Ts2s7Iyi1Tn
Ls/NqJIyjuZS3zelmWvZQ8UblMDELPU1ary8mYpz8oLu8gdFkTVWYioPFttZylbK
003gIlBd69lFlW5Y1KCGLC66NwytC/DQ78eDiITi/KUZCIJix118zhayRc3gQMX7
iRrQnVc7L5ZBxvPlHRWaM/RFZE4vpjsj+3jEdBZEu5Fq4SLx06mX3xqdO6/W0Jh5
2blXOdAO92q5QGFNU9LY1tkITPBjBmE21jR7fay48+oS0savKHtWSlzkuavU4GPC
P2AF6WAVWKsUXQVZgrMamGK5nfAyAbUFxmn3JB2BN4wuJGvptCUeC69/YHPD1s7d
+b4SgiPgkZhx/iOMDUWX2QVAngdgfVvZoudhpUFU8cceGxfgwwPN4QwSB0+g8rQQ
DnxOYSSQS+Ym85rRJocVX9+0X+TAKGi7E3k/vzaFQYq40//1ucBphZLJVRQdwZC3
NdMvnd3KRzE4oTl8gBeeFrwfb6zYGUmPKxU93fLNdhVKqIm+Y813/7o5ZeVWF4Pn
CWXW/xVkT64wHsRz929jHVRH/WYVgSLSfpXRgEVtCtiDp7VyKXr32R2crcn55LYT
wDK4eF1tLE0XC+nVsfbBw4O0KotUQIXQthxVzRBqujvt1YYhL3lj9r1SiE1xzy0s
4wxuU5OK/+IJDqiSWS5FLvoXR7Mwaaga54a+ASAAA3xBnnWmmiKg8g/IEHKLzUvh
t8/60ofeeT3pDFGtFtP1Rx4sZVltYcxlWpLwqYWIR+M49RVv8PJd40Af9hmAHxmV
kwPTEOtIPQl1n+XsAm/7mR0g1WFe/fjXx6qCDS0LVocB3yOEP+238cozBoZd0ReQ
2Ao9DR5JSD1uObf4jlALyT3X8wco+np7PAw14MKSQzb4iq1TfROQiki3Qg6wrSHt
4rFInP5DyPezh8zseaaeXuhl56jY83XJa2rgf7Y/GsLwCJHrwA4sQFtgPElarHQH
LJv9PaMt6IaGOAbiXDzPzPmVMppIJOWHOkVNX0wY1gIRa4WrguubBEqAWsd5VUDT
SvxvbA2NdcNtfZWLgsGsKNR0H1Aj8RMov6e1xMACryZ6UycA8nJpT/fXZF+8aREv
SROSpE+MScfJCRJHmgYTSrEi9/o7uQ+p82cAxue3H8C3yCz2gKEVU++VGwLpkiVs
ZKOqLd1G2hplFfzZabr7BA/J3BAnZNDV0ejgbHdnACEBhxUyIKe7zD3K4sWkYfe4
ymN9sIMk0HDpe1LY3nA+frH3Fk+LC1DkamYQJc9blSa29ScKipsAE1B+eAbU2TZz
btqLXA3fL8X/iSOjqkW+IW/ppqYhQrKd+nxgFjK2xZZAljAq8TuwN/Deg9wn8sZR
hymKGefOsen3Ktg7DNeKwr6yE8ZlCmATgk5VbxnYk/AcAzNDidOKRf/dmmKrKXB6
6hmYVofkIlHePF0tJEzK1mVu6JgwrIlrrYkbH9V1uImGtyHlrwJ2xokzjlptl/4W
ka6PVFixNZLFFPHtuHVEU7P981xvrZwjNClKlt6Kw4C93snXvc4KazciNH3mRlpS
kiLXr6TLHIQAfghGf+cpzo3VSv24WNH4pvk6dFXzA1XK3TohQbA5AQU8d/40FZiS
qO5WvdRlgES7+mBZjoBri2lbNCPYkdsPRWpF0sXfbSyVdHMzd3S1LhqhXvBb7dzR
/cEAM5YmclU6ERw2TjWQkavnxuDm5aR/ZkT0+7HMlHwSlOrNIxjgZoIQC4DVbs9/
J/PqJ0HwuK9F1wNeuDuUovHDJJmSoRTtFd9x+XLrFZ65hFnjP4oan2g+tORPaMR8
ikIqLeREPgkddXesSbfs/nbbdl3+Ibn6+sr7Sl9ZYB/vTYLntQYfTGSgezMhciT0
hT48rzZuyZ7EvHAJTUDrBLmeFZsYKhwMb648vlFksTm+TKEQDzH2CbygCQXy+gOw
x2ZAO8pX54cHRlW8UHoSYPf9fAmPFfzK65IzHi8iZ3tQm5jHw0bgkNAhpDa981On
2ffUdswz5eoJQCICQcxX8LfKAxGSkkx3SxCa1mUxZD6B/T+2sNTbiFmDw9sgsLwo
QELq2neeVmJS32HbFHUaqYY5aQm4huf8v72yvo2TPfcN/b+jOcs/B/K3yFbxqtWp
SoSNSW6qRBne0EbRa8Jzc5NItJfxjdph76LdqYkVFf/GiBEFR1t9njs/x+pH+h9B
fJF5fHQw9SYgu5ge8RBPgVhRD/RN66/FmWmxUJ1y5bMXYDPgJ04bBHBWwrfMBMAi
Ba2Ie+X8sDCbHgj/dyGiHjdRs9v6O7PRZQIqgHov6i266x08WPEWCbZ7z2FkQ2Jv
7KUK32yqprjQIT5qr/zG0kzcorbnSJYLzn28CMIucQ67s2SOgeq5j3UdohOzXyMv
J2dUH7eFEHHE75qwOBIryo62xV4RXqM9tYm304y5dqdUWPKxeN8bhYXiCZjsSOOm
yDAiGlhFTRSkawQqnJ8Lq0IiQsPVyzLfrnlQKCQECUihp/W1ldaQz/poOk7d3i8b
WRo+915GHtHd9RXY94x5fJGVdWZiB3Q2iFMgi/u/5FzDTBu4OlrzPTNq/6bGUZQD
+nyAFIhUfZQ5auhNr7ycZbD32gD6RvIn4mPSWUXGQP7zxB1hdANFZ1vL4ZeOiEbt
dmKrFjm/f1QKsZ7YNP/k7IbM7rUEQP+70x7OHsZqCRCYEbGV7w8VqJdeWm+GXuYS
BsKDIm13rKZ9vC7sF6pcRhoNTKTXSqXhtZWUmGm0UwF8e/dh2LZsHYZzP0Hd9CM/
9UratdHKeeMCDix+reawBCl1j6Au5HAC8npBtiVnKkSTUvVOIx5p/IA5vrzeNv7J
jZdDwttLGNFmeJpT3j8nIJxLPSSZwlVcEoes7WdJ1mGQ42kiB0Wyyo3fXYkrxBnu
9LkZEupOzr6oQQVHUzjyB75dcn9vabUP9bJuDZ0PEA2z4LuTb1CvKuohxsPp7RBk
xksdu0OUXrMBcly4okQzWMvuBF0fNwOjukWmir1HoaSmRtbPTBRW/WhSgxoy+8Iu
Q5dKUYui6FxfdEcwXGoT8T51lq6FJQWiUKrbejvMUCHtzcMqAipYLSC+cgvsDmLp
kjxu+9PaaqF7DNwIf7m+D9zZR+vekPdRnVviw578bDZJadrW8Veb+85y6yyiRuGz
ZGE7TzNHhCK5WQnzzz+cRFGIM7fE4BUoT5Cyi4546IOz0fwJFZI1mJxgSYBiSWbR
Bqiap/jExGqZTedBJglyj+ql0bgWyh+Wvo3fe0vfRwRMD47Jp3yIi+WkKC93Qt6I
vZAD6JjD3VRoI0yXtSR5gxC3YdnXL9a9RT1Gb3igLD6OWWncksWAVmO4Iavb/6sh
w76LZ2136Xn6Osm/1VftQ0Ki+DHi95rnKFgX+ZslXJ1C55nXjRhR+fhS7KZfIMTK
2Q48N5dGsIdKEsZQZR2K5poUFeAJ9ofzu5kstkxU2PEgfk7xUMdl5rYdv/c+1DGi
83eHCfF4rdy4g8/fSC2+QbZ/+GDmGJopY2CSJykOIE7Wel37MtYYhGmWxyLAx3Qo
wFs1fl5rWOBm9zV0hJqR4ISj4P54v+yhXD7C7SBPWWcYQX9dEPXTZQw7UNonvYPb
QsLuOilOTob8j1Hh7kWPEk8joeckfeuj55Oqn5fAcVXyVfXacoOU49oDUCMcj+tz
G3N1Rbjrx8HSEStAebtY7WPXk1xV0a3EOnf8CL/FPRgRGN/2YAs5ta55GvawhFsS
jZ6F7akglSd0iW2hY3CU0E2QhtkAmZ1UiubTE3tKmWpQO1o6yDAkqgciOvWs3Mcf
BDrJiJyhcACvejcQHkjKXJ/6xpDwmhDGLo6OqcqbhLMtsbLxpyv19hluMspwNUyW
x6PdTuekTcoQ99rvckHM+hsdqYzQh3LjVKF3Obg9vc4wh6+9n6CCZmnKSUI/K8V8
QYlN2wvdtc7t7MubbVSgaOnMYSiuBpAyFC4m+VWHutANpZqnTqiPZfmfWffKrLrS
CvpdPL/LBeLhyHna8WByLSQeMBDWlrPw1d33wZqXSFmyDTe/QhOQ8rjHZEOBqPRI
5KbDJ3M3z6McyxOcDFSE3OO0PMEbqWMirvK6urxyQGFjQCJJNiupGVCtLrhHLui5
D/XEh783Kb0TDn8+OqsZixKUk4lU/1uTE0uGtFryT5BTe+nTK6f3hld0vvmCAd4w
auP9N8vEUlx8nhvTB2kUPc/YgjpkCdbT2M7Mc38KV0FVQLbIOiICS14VF90cu4Z4
jCKDsgXEtX9gSBR4lSkZvNI+3H/g7nmyd1oXT2xSDbNjSNsjS2r+JRkuj2JLdixd
xGMSnuwZTalel0bpirWEKWxyPdgvzwBwgheA2iK8uOYDqWoOCWs25QpeRM+Anm7f
DYAUlX3RJ1/DIthjYEP0cKeUGUMWgNXrY/1lCrPD0iU19atplqnL6fOjBrMxLg7r
T00oBBstKpBzJ0N2ohlEq0mTPKbP6Gs7gJTgyw0nBTpMBqLUdU+bI/2vd55+noWg
Kp3wYAozQrKWdOy+mHO4Kid/5qV9vkQb+NWhlQtwRcXWsT28ozt3BsnpkLhwfxMh
tVQXcsCOeuVMOLWhTGH9XoM7P/OBTTrSPt1EGm9b6VM6wszopADSUQXf0bAgk7TI
tgtjqV3+0bXIFkuzku7c/HGyS2W67UA4LGWciyIp4mmfF6qfnRjWXOzzJoyFwbzr
gO7QZ8+/NliiwO5hM5PzOI907dMhZmOU0dBXS950vDvcz/z833NztZhitnrIuxYP
gt4v6mdE3rnZEJHsesxLYCNgcMMPSHsCAobeoVG9ordpRjLXLZyR7vDjAp4SzwFl
6hWCW0CkyqW7iNaj9Jof+gqsw3n7oB2ExFRqUJ+/qRHp85XqGRV7OsuPMR6VMTRl
jTCU3phsjJmjS76EJgNCPO8JlcSqTXkxtbVcqrJBr1BRHgM6XdFJK2TtLM9ffuvp
123PvULRuiA8Nh4UKSjBtMWDH61UlBD/0VKie8lz1oVJ9iCiRPCEZR7v8kaEC0Dj
V91eUiAwblb+lYh37rkLXLI0UQwxNbBnTTHmDwFhi3TARc+SKKbND/2MFM3TdcRz
Py9nYmxY/ezD4WOVwPN+9BWx6XpkiVb3HW5DCgK+j0VpzIyNGNoTvtN2UT5oe9/Q
+Z5+MHfa4jNhIIDRcJrfacatS/hzv+KtvFc2fRPY8PUIKw/+dy4zRG4uZOHxsMQy
qhU4U1TsFxVVXHXz3f2DBtdM/LMlzlBFkcmAvWK264vb5eEgaOfFkgQhxMv2lJ0I
IrF4h58gYFMSefmYZ+dyCpDwQB3N+Q3Yu0yCHSuRpjYIMROi/eE7WhwJY88vzCOL
1nJEN2NFys34gvE39earfzTpS+LmM1vILCXkqT2xHI+M+oDSsTQVi4vuyfK8CXSC
2k0LSY8T0/JX8/LXNu/OH0CwvXw8VRjkvDAu8n4HIuqv6sPOdGYXjy9wpTplM7MF
b1wDGF/0q2d5TBR6lNUWi2x/Ln7Zhzblh+RDP9Op+DntKP317/I3oYhVtTAqKAJp
KyALbzYJlJqQjxvF3r0OFDkFpp6+wCH4RjaxOLeKB77Ew5qNOIqEKR1vcBGfw/zn
xd8996x5xT7l6bnj+zn2Lxq61peVdFVdVMjXEucignu727KeR66iyLq67mLmzzEb
fJZsY3D8n+0XbWa5KGAE9uMPF4i5VXO9pGZeNXp9Ck1fcJaJMeKFbqQ3mRQDZV6e
x2SOtRiLe8Q7+ygveLhDid9VgRBNODPcmv9VjD/4F10hMKWQjJfzqY9ENDXdihAf
O1TSw4Y/1WIWqGVUqLIFky9ycjkZn36m/1qbDb7LSIxBEbbhnfYkI6u0Oo65lI4y
kfDCFWl/43XM3EhKn6kv8LPOmN6sQUebmixNoMY/GRSBr9fSvteDK8oXF6WbhDIp
mMwwFu9B3zMVkBWyA/9Aouv31Ly2McT/Bna7XNywvhzdkxpoTJQHU/Dr6GMmQGIH
DI22+eg5LlL138I5BWa9yy9v6LtQvfjQC5nwhq7xV8mkt4r6SJX+oSB/qtJmIhYl
HPvIlebm9TbuVdNARFbauQamM4fDg0lPZxZdncNR7EiAEzlibx9y3YSxb1E0TmZC
Rw6GZRL6b505jXonvtLoUeBHbpNhlxTiduYsOe5un34XLtrWAAvJLlqLFrUbl3Rb
l/c3lb8LBpWzdEU/FivfhrvQaO6h1GsA9fkMQE1sG5mC2OvTcAL3BAk671QT/2B9
4GoAgd0tVqtTi31BV8a0kSGM2oqBD6ZhDo5d6hGeqaBhtKPG1E7CSymtz9Vk/iia
IawArAoVZrzNEbd4/mLLLGp1NpiNecwmeJAKIOLqUNqVMSjSAX00NZYI+y3uxUEa
O877SObuD/uRhqcCcGd92UCVVbmYadm9DPvX3iPvMxjMG3JlVe2Kis7HJ47cyv+S
NEdNBCHjrFllR1T66nmH0kATO0WBLSbaYP4hEovrcMb9YLbAKtdfXZuF9bD7B/rT
k3E12AXEd15rrAnUVi1IcZdkdbjOjZtPVdtGCBzfg4zanbZqcPFNQJBcyyFvuvPK
010moa5EXn3ATYACSPrU0Gkrl63b8StzjmiM49CEet2Iq9gIs9yVqZsapl59ZO+U
kgeu0LitducF/26PuHz0fvJmyqo3fWPoo31KFuexUGaEI0/IviS0vdPIhVvHAdfP
y2wQ1OAhODFJWhWs105XE52haFCDiwiFO1dd2s3olXbKKO/IQy0o9awL+CvBkZAV
CPbXpk3j7xEzhRD4aE3VfnmF2K5+QmKeMPBWYJ7IxGIp8J/G1O0F/Cz7NzYNWHTD
BeHYchxEMsygj5jMVWv5NF33rg3mBC1M2iX2zi61Nh2p5FJfMN7D8I3Cf2uepT/E
oPYwgr/cZsLu5dPdwSIV8J7OqbiOWCg9HriUhzstwZ6s6wEKq8a0TlpD67OfMfzs
ey54Honx11zyBPEnRaKO3kDVVBsMaok5gUEqkwzHdkQushSm0DuO8LFN/EPs/Vo2
rvnKe7YHhjiXNMhd03NcBux4OeZ7D+v7L7J8PdvtJqPAuT6N9CaouASxoe4SMiUb
itLd55nrMMPhMcbFBUtfxMSxtSxFjvJOtt8luIFWVDB1oDveu08Q5IZeRKfS5dOU
EVswOa0L6hn0SU25bAjvtc1kYghSATY5BzE704MODPwBw4XKsGTUdtcm1iBQaPq5
j43DPcXtWGvUrzFA/XxzIfhhWbFpRg5OGzbBLbACbSxCJhpvHwWmW2053iX88ZGa
jGiixCg0Q31f74fiSHc2gty/zvo7lc7SsMwZmg99uVXYC6bzhBu87C2qH1m4qcbJ
Q0qTchswISdfWvHx5ul/Gwez9tBS6d1+J2e5Hrz7oLU2D/cOEMJ84Je+46Um/XcJ
huZe8/2QWfhaHlqGgLNv4ONnfQcjH/8XhXDaqGiLj/jXpNBA04jo0cUf1eRJ4V/K
RnNVu5vLnLeKFnvf43g14ehlTXdPBIiiQlKqWjufC9Q5nKkKnk606uRQDcNlLfTW
A3EyVwZ8hzrlkGhXOpQ9UXbzXXuRQVVK2q9jTZmRrCALgPN/gL/CSKesca/H9QDn
ILmA+Nz015iqtrgvt7MMzaaFi0Jq4K1krdIdCzlbF02MEs2Sm78yViKeI35isVEz
D7Jx37bS9LLfQlT9qs6NwwuHg9EQZ7/+MavMQAX5rxetKoubw15a/S0+1jIWEV9f
fRD9Mv/mXF1SH9986WpQ4e4cSmXxa5ZF7iWmOhxBm72OJ3EY4rhfGYjt8aiqa7Sc
yOkGgqCAKSKzSOT6wuvUIYgvp/6Hy7He3JqdaK3WpIE7lrbksmq6KQi+UXFChlac
IrhiJrfIMxGW5fteKGlut+yyhmyyA4lD3Ka9lPcSIx7buEH26HrxWGnDxLeAc6zZ
ybpi9JqnTAAqGxRB0wkqgT4B6O3qSObhCNLbXfXG5lPFGxMSI7iNf3dfm1xRIE44
rAB0cltj8ZQssiXK8lWx5WISomQf5x9mZOb9zNENngS/6sUeP0ZOHW7xHIsM+qGF
N0vSPzUSSPIZwCXKr+x+Q3aBMe41Mq2EpFapr0NGHdMS6hbjTMeXBq4eHbMvFfz5
8xuZ+XLyZVZP+zcEXaQx4mF2cE45GwJ97NYMc5ABpQp5X8sw3ZOLRiMBoMHSuIuK
tcyFBLW5O5oFn7VbRGY9tQTO6vftwK/5LcDLwPSTjf36r4zkexyIjIKwqRzB0Hg/
yWRO9cmSWIv+qYE7st8pZSK4NbJkXoG7gUB4DJHEfS0GnVmVNtVuRwNDae8rSzk/
3Yn0secBHpwwHYZ3tZgsI4wZgabs0asMU5fsycNkSdjISgzpE6il4F0n/fjm85fb
fpsHyYG1PxMJs0ld/6Obp8dtY2QT5IeWTREGNMekNhLR68Cp0Drc61uMo0nsMsnN
NWc81Lj94bo5dwZy3dbG20ShcJ0riE4sHzm7oYSEebvsaHa7OQa29BegpbGbF7oe
+7QoiBmGpT6a7tDkkIZrEwE11kq/FhnZ2COXx0adDMVIQdiYjtSrSPG42PsjIbBm
72ZqZdAP67cPdy9keK1j1DWcNUA6J+1gK2brWSlLdgPbcJmkiG/wI1vJtLCYGFWb
phLi4tB72XgMXWBdGkVtEHTABBTyvBk1I2rUlvVOqquE3v2Hf/Hvn6OTQZrZUAaG
SDhl3yE6RsToSvn4lFbr9bPMpGY6aYnOpbiwWqzt7d6BHGU3vLJ4w9P7OTz/2GYV
WpEXZwf5mOhRPnMiy9wM9g43rkv2NbQZfXuGcsQRtGNwVfupSzj5ZzqHkWHJs5MQ
POJL9ScH3nWoBnsnWN//pka1aZp8T5HVMGCyOlCofgDCT+P/w9TtvtKOTfYmuqu0
52c+rtQatpJ+Qud0fVqsX21z55V2bIPqoA4Pc/FuubRAoFsyIb0/ewcsV9iBCjTh
FnS5D6h8wz5ehKXKj/M4oQ6CYbjd+SJ6PDbzsmuH6zWzjySp5vTfoCjXDHriXoMn
7bhb9IU2I9mC8hU8yPwhebN2eofyWH5vND7Bwl2CRIxrIElHvR6kW5qPj1PshM0E
7Z16S4HNG830x+CrVht89ZBiGKNvato5Cys7D4eNSoWWYJbJAxE7lDDNnNia3UDx
vNMoDmjS7xnby+UR5YMfiQLxoaBnrk1wXbnjqbjkSNA8j6Vx2TuzmVb0GfzPU4yr
AnUjlK9jG+rSZQZveRHmJexD2DIaBKeaUEsqFyWHKmMgZrydE926ZpwqBQhMidxm
3nHUtDVUqflfp0KwDKK+Bg94+eZsTjII2pxR72e5ew2T9x4oa9uRydJWZxMdnXOa
LBAhiozMklK1TSIWRHnJr7GvXsAspJGy7Gf/FRW8P88kS4/EX4Yxex3UJ+ZUo372
Yc8pDFQGPHM4a0mpwg6zmtS+QZwCmdW4fiJ0o3woqy6flmaClXxZ+C2gLaC5q9Wh
3Sqolykt9GXHQBtfMm6dhRXG7oOXVT9GM8/+NpHNCyr9mpfrEkXWsqhDZODXCtpW
LmrIGRf4OR+rVfrCRkjC/25jPTGqCJe8xWgVXhxxwtiFi/NVCDvlJjyVYCuLM0UI
9bSmEbPiIzYEiZca2dku5lVDbR4EPHa1WlcytAoFPwvIch18c/KwxU6kzR/eyS56
trbkgjUhncoKLjRUoyvKXPa2GdCeaQ49Ed0DZ8YlBSy3wpPXluDURmESgR3+kIZ3
GGEHv+g47D1DwnHod11eD7D12phsvCJWI6snyskXWFdG6Kw/9HxJGXFgzVs1/QJw
o7DLDlCDC3LEQ08en7gap0slYC1MrVHB67ifsVVrpmtbgzC1dgtoOpREWbsZbg59
n6Tk4+ygkT+NKPjOFJWtYmV37C1q0Cd32P7uY0VAMnScL9rp1icz15AEQsacvLmQ
jBj/2QO8i1qtbi3uLRqzKW74M5EpzLhWI/5CABVRDIzO5lnIBMIlqT7n0ei9QlBb
FEpQnIvmXc5LVmzfVigb1ALaGBqM3d0udPEilJpGXic7Ju9OOhz2u2YrAl3ItWbI
PCAg6aeRXdahUAdjWKKQQJZTaXby+qSUjvt8LBc70uqHWov1UWfEp2NjCHIGNstM
0KQXS6cJWMMuwdLWPmtwvKrUEWe/CKJeC1dV7E//IEaZvX3W/WN/WhYfSWFT5nVe
nybBrrtfCTI5GE60mbrqX1BTDOdbSeAsB/Jtpe36H1tnDtz0XqUxkz59IiClDBgC
9+tWImglnmw/Lll9RqId90y5jfSNwXScaZfCn1ukSdJwxaOAMe5Ubr2M0LtBT2Z/
4RVcMaZsEUO3x1ywZQe+vybJxDhZQt8BuRb1xmtxOdpdQI0sVKUochdmn598JwoI
0ir97aQsNoFGFc+tqNaLRP4IJjdf3ghHNVKiG0+NaGwR35HVhNidZSZO9AKEreHk
qR/ojprebRboyeFFBoL+e0AcuZNpOY1vlBshyWLbzd4Q1UZgtO5/XsDk5gxlGt8l
4eANneozr9StdFsA0XDXBJ/RZL1SGjoqRqGUWdD/acvYbApADR4mdRc+jOmg2ELH
2UkfVJooLw1hMmPiVh1tS3Hlv8w0fJz4o7C+u2fFz/DL7xOYlkGvelu+YczEFKcK
rW9EDKKjCRzrvbbh22zK9ENVJmBX4bfN8JLp5Ctq8touOoK0GP7xoRjkbVWtUS4f
AA0tler3ikpHQLBRKi1Oi0DsMhAF0k2w6Jknigs1lPZYADmrayp9vLkd64WT7Aq/
rhg1/lX5gK3X0kzUaFDZIB0wKE9IRoo1fW3u9IzZozpYhIOZPeoDWEoG1v6p0tHk
N2p+/lP/RObl/AysXHHZPx7qNP4ElanWGc0x2XyHurduOmg14FGB/WSkUSoPe09/
YzNxnlQ/pNXH51GJgRyGs0W6+lL4/RIf96ryrfwIJlNySKBqPuj6APr4Stb0KABG
V2UdvS/xcLPxWS9A/6etWx38Dk5Ac8NZ+jtf2jh1NxM/JzY7GQbTOhe6p7IUYHLY
Xk8tjsrEQPZUhODimhRj+0QWF8Cp/zJd03MXFJ69TCTT0gCxIUdqxPoEwUmy2crB
WtzlitwF0L/0SwXbxOEsct7cklIKOX4+ciXEG++r/uh8UfVs+rtGvCG2Sq6cmytZ
4agrikEmTwcx0qy0AFFgU/K+EAH/rrV+eE5KfwUYIbqh87FWNVlviK0GQ0qtvwie
XR4geJeyf8X+fN8UHitoQJV5Ds8Y6wpK6teYN3lZiVapjXKk8rGLXcMfgcL5qMfQ
B8VAHUE6V08xutvKlncranOcX5UubP8Tq7vs+7RXcDtWODnvSDMAK2Jgl+sZiq6C
j9zupHiovQAnjLXvc2B+zMoPzRBd8VeWmr8oui92Ke+zSyTX/2Q9EX1ksCO/BdMI
qL7hc7A2/1QDkxCVNZeHKRMvSGQONHavPU5MHZsAw2Mjs1zNlS/UQMT1SWwJ4KrD
LkTPlbRzKGMHoA87fz8JGGvSMnqvfSH/6miYS4fRhMeJqqv7uSEtsaf21Hg4Bw20
HbojOfgsZ5S6ZaVdQVRkdadAre9AXbMu1+Tiny8Ru9RrtZodkMU46hT8hFUyJAVw
eovLFV+vnIq8yCfZjFiPpwsH8HJDpdgqTYxLq82nf+uBxZa0ju9V/7s8cOS/+sNC
c5dfZviS96jE8kfYeVhWVUYK2sIdTqy+/0uuWk7RqnJnxpfre1z7S5Ihc8d4/B+N
8iULnIWVWeTPyzuYg5nYsdSQBDeneIEkF0Qj5c4KfxE2zNaJsNEmH6ZcOkk0YPBd
GMZxbZgxQNu/8ZQuYAMNb4qgAMOKVHP13kWtG4JXEOHrNuByOpvpLz7gdGxxw0D8
ToqqTVfCsmHLuyJOBVYlL/zveZDQB7RSSQt6oxm984pAgnMMoy6ST77o4dWlP6zb
q5KTpUBW62YB8wiqAhP6zFeNUXjDxMCGOFgiA/izDfmdibos6zrQG6XNm9nRuLYD
DMzbixiMu7UVfGNPsml4O5/pLsMf4KVwKzpFObM/obFwJA+4sIiDr4SjHWgyp2H/
el2wqWKfbtmp35T2bAGk1eh+5OLxrrSS2Tym8YIEECLTL7S2e+fRq970mEqEbMpa
lRbGIG6d4RdPAWvaFJABd6L9yg4BNsCK8NqaRnwny7TCBRwZW9nb7Xz8J34Ul7F3
KYj5gQkVVseJXTakaoIJcar54AjgRFix6fRxYWAyfyou/EWk+nsY9wgISNYxtII3
iweIbV6+4WfvsrHI+F2p1jcjFG6S4tSJaJA8LXZxWR18QduCoTZ+MKVZk7+g2Rnq
vR/tSWiX97xpjVgvBdydg2nnTnBuk9KlLzxnZeq7Ok6mfNDsLFu5BccVAw0EJuTv
KpcrH5MGKe1mNeek0ARUdaA47khambB9ayMju1u98gYalTg9u6vG0H51c09wE8fz
el7TIITnpjpNnxDOg2IIKzhlgWpO4hy1OuVHyZ02nZ1gJc9P00TPVFgO0j6dZY1J
RGgG0/XCIS8SvGUJZlXokahCdw4qMtx7tOR5lX6AbKEmcLc6qfA8SoKwqDZ4UKir
N6oDXP3cN3XHuNg+VdsXzwPtDSeyH0Nfl+ONVSQKorrYWorlcAfF2kRnUxTKCuWK
pOewJukHOKOsf17UmLoUSThHs60mzfN56nhnU9TsjU3LS1e5X5twf7xfLhCWBCun
OMUPX4feOE5Ck2sDjtBT0DmCaJhicavC+98sUWv3CPwlGdU9iAKdqXEu0QKjls0k
Q+3OWUZNTFbgotpoSocun4TuLC2Hgf09W8iRRzXmf8Ar4v55XYXsGMSWJKKo8dGa
9IwHh3AFWVtFuqQF7RIs7O+MWjWTTBnJ0T9GzVqo8taoVnrFOpP5WMh/GGPUVeu7
uqrbn/DtrPF6P35nZ36T+bnLZ3tsNT+kZhD4WyvMEI+obeFzBblHGvGrclIcFPZ0
mGShOggDjH2coD2nAYLScVx/rjka3eNM+g7avxVmZsyxkud9J4eNcOtn4KLxTY3w
HkOGBfzrNkAOHBSYdi1ERx4/s0mc0CtDH4tjSG6fzjtrJgRkXdxA9HbkD4qaTEzD
Idhbz/Er/f8I/LjT+UkK0AeYgsZ27Hc2MhTyfHw0cK52dkVodIp2jAC4769fVX4X
WGZ6ukZXEV73f1P6JIlEqBp4YKtDVq3fQM69z4kzywob0AzkzaA5JhJxATxM6uNM
Y4zD3Tww8G/8+W1vgF62JFIBGs4qdrg0rqv/esIETk1YsTqkq30SFP2zTDfr+VCG
3UNmHr0Mb1phzEr20DQAblTPvWsIjOdZnazLnaRmks61kSm3Tnw6fhq+JXNISqCC
Oi2oIwuDRXC3/5Pn4JaYFYkKU+Gf2UPEc8Q9XLBok70OdCcxIjCYnv9sKtxRVdlx
avNn+C1rDw30Ya3fDtxpCi5dgKRHrsMAWzUNGtZP/6i0ZKg/6nX2yS1+uwfMHBKV
dI/GjpkXADLFLGe+xOCYEiM0Qluf/JQ5cCK7lKng+yocBoLdbPdswqbreHQd19cq
GM1TKeq2NKO3XqCtL1MyoUJFxeoc0gs761yxOH0jxPzyorM/2oTAH7cXZqMc4oxj
xMDTbUrsi2DyC8dRPYnG1+5gX0A29bbMF4qO8J6v/4hjahs319bQz6pUQOEPpHjf
5Wa+fqSqBCEVbD1+z6MgorkeOtF04i+K6pdGmYk7T4Cp6ITBhhgUXTUATx6aA/Y+
ZNX6c1DWsxA5/kj6hW94Rx7G9lnptD+tNp7v9EIIdPyGEY+Tfl9Tlx0G6lMlfdBy
cPoQn7IqoXl0h8xY+F0uTBWMi0L7XbVl1DuxjCfiJdCn1lDXNo6FaZlTadMonc1W
R81TAHvrrc1rgiRYLQ5H4h8lvXMYMnyQjG2dJ8+AJFM48T9ydEd7e8F200zHZ3Ev
Nf3gsy/KYJo80G8Od3w45bfXL+3or2GrluN9/5Ru/ddPRVGFN7gA6qsM2LgM3IY4
Vqiv2p4fnLMLxCaQhWB/iYx6evMW1HetOwxYXtjpsT9TwgQA3ToX0AP46vm1jvMd
kdeygX3/YqVXzbv+Dn5H2R0qBRtTratXtUTUzkAhe5YUdU2xY8ccVRaixRANjCcA
ph0hYI9oD2l6bni9zsxDD4PcFdZAAVtWKCAnM4WzOxDgullRMYU2+7vctgIkURg8
tyOC9Fbe1ruIiDd1aTMZAJnWdVaCkgHZ18ZvMnzeEE+YBxmlmtKMeKIE+aDZZ3G6
EuX6L7tZZM4YsjvokQmSNomyjWr/gEO32wANoAyZdJujCNJ6PHt/0dEyVY3g/JeA
UsyvqEn1w8KfIac/zxCsOK45RdGUAIXLhNbbsBdhuwwn9CRbyWxIr5iX0kI+9+ZC
tDXR/k22iMosHfGz5Tn/0+LWe1zWyViM1URdbV+XxIipeVSx1YQHonHfGKkB2CGB
63po9bUeEf6L+OBICkgtKbn6C9vbc2gDzw5Ul4atRF+HPvDbzxA6IRUDlCIEu/37
t2bgQ7PlRNFTsKP2bSevBQRVGOwaeVIhlQo6i3YQhPY6HWYYbCwFkTuZwkIIVt9j
nignr80JSlF3uou3/CcATRKSB1c/NRYciv4Er/XWOoyJnM+OpU19Z5mFYAi0tkW0
Az/xOouS2Fb9T0NdQZ+gWcH41f5U22iekA4AoCXnZwdORd/eHKEVpwDoIR3wyxhf
MrI9SgY24erMgaRWrW/rgrySGa/Tt2CY4yxUMrZrifvl4gqQEIW2KKZdmMRbpKso
sYXlfU3tOBQGrr9pFnipgHHPl0slpTV6dmvQYssS0HCEpGNUixMTnA7F+PJkl5t8
1cDotNXZfBmTdTa3Ka0mVXn6/WYJqgqQFkSHuAiqzC0xCvdy0obzGsaRz2Ul9+S3
tZyM4hGAjvIQ7utBvjqEJISyHUhzjoXKt4BgXVfgjg0ery41WJQEVo0LHHaDq43V
6TBxEE17i1Uz83bVXudNjEuW/uR3F5jBa8XJZMy/ehaYrUGWmOEpSzodpYiBdq8q
na5S3FsDrEJFXBEvcyuqSc/cG2mjrCBwxTe/NZDVIbxmfAUls3u41s4o9Dp17C6/
pqCYOtXM5nZ7exY/+nM8mE8oTsjNFQ6nUbNkhtiLh1qmUJ8bUVjyhImvbWI4I6fP
0EaeizPXmoa1r+bgyTHUQjbYxFsGoL+BtToTru0k1cB5CVAWaEx68Qjny9nGo8u4
8sCul1gj9I8BWJPPl9mWcBy1Q73M/UbQ4JozoGT5LLdHmH3NxOArABUv60g3UHjP
YWI9O/IqKfoxCtGEuWwCgcY5KqFpT268TxONLciSmL5v+HLI7mJIA3f7+97pk41Y
QsOtlUU/GzLze2+t6mULCI2+Enrt/a9vy1JXjFsKy4wvOXzNLgfYAPkk3xOLWlkK
/4mx5llqUGHk/9qncxXpil7BP5+5pFktB/zwyd+J8fPcbH90Dc4Y8H5AK6J0Lssw
TtEYdmp5hoLhTgovm6UOxbTzt4rZXTXxWySGM1NItDT61OnC1Rk7gJPEPzUfH2NQ
hgw/yDdOGN4WVXEJiU4iiPZ08aLZ7jhrpJ9JwZkUXVyR0OVIeINer5oBbqZbVFQF
6WS4n3CY+oQg4uXWBL+U5KSN91ir9Z697LSjj5pW7haIs3j5VUD98aT8ObsjMz9a
n8HUKi7Y6VFxS/5llBv+CIu5yE0FU9eeFiqQcjQxZ4jz3aQgjr5JyAEv0hEOe3ku
CFuEYeQnN6c704FzDalbKVKioaDfjU7X/06BtidVq17+Qv6W/Erqbw4u5MLfqhbD
Nf3hZ9HKv4/26SBu/aVlfLX4yUcQhBlJaJpdEMd2/o5HIN2Ie0jxJedAnnuvRQPj
EjQoZpKDl6Vq421iZY2Ie0GfBHgYNcfUYMoS4b53sp3zUtFsffOlXwASaWM2b6tY
DvWi4PN65j/COfJnMOGWCE71uCXJc/TWMriNC4myIRcagvzFZI/RmzZ4nYjKt/kg
Dsd4AYGt6OAi256cCKL3+zpnDAEfctFn8tU7070KdkBuU0H18o9D7CHRRU1Cn4zK
+t9NNK/9ct8If1lRiTEKVIGOCwYTj6ayb/PCco/g/zv04zZEYjfKsec5H4oESEQl
VkE6tW/oaAcqjbbN9/1h89j/s00WM5cMzxBf3TIeBBZgKwRU9H+7gwBB8skAi/aq
9pPcow12dUPkJswm6TQE2Cn4aEeuFZtnvQu4lc3ZQcaOigP+rRsvNWFK8LrdVhtm
vtdXc9iPj903BvLYMk5TTGJPlKqNpSqMzZ7iC235pMm2ptxYubkCvqMELk9YuFMV
ah9ed6LVjG/5lqR9FLI/A5KS9z80a8HCUKnDVsy2KcpRpPhS2EQCio/C2UBitPlG
NF9FioUofv0DoLV6eVq+oXzR7ABhCtP0xWXag38gt+Hj8cGZhTbeeYO1AfAHGXm5
RQgRW2QRPTp5egK+EZpdF27GJnSDzOWDY6JMmyZygWFc2J80Y4N6hZaAbD/vcuIE
CDEDPb4xPz4Tb9uWukzWtkUwIfAN2COipMEP9Q3bxnuf4cu9r7gwhbZD4YIuWuB2
Ua0jnFK4Qh5N4+cc5PENh74WDqc5IR+wpNJmcC9C+AiBzwF9PHU0uaBEIA/MBhRT
8pHvx2cQ0KxBG26hP4wNlFoa0iJrgealJZaoUr552evjg9Owj4Nqc8XWIH2KQBWL
iZMT47i3YuIgaC8JlCzCbJCoZZa1Eg0MeUmXOsWUZ7kTrnedhQJCklmj4LyhZNHN
fTXIY88n7ywAOPAR2PqV5A4DlQ/lqimN6N6WFuXakaAxL7KViANaBUemo/T0lPF3
DGw8GR75u4avVfc55yzkKkfy/rQhN9IMe3CN0bUX5LMDFZVqFc2jagJ30QbgJhLl
5XWKMdKo+5ej9sxM2yRhlEIthDwMXBa7M2IG7Kz7YkUgCHdghqxYat9RJivA18MG
aYjTFoKcSEcYp6EDdG2s2KCfV3aRr4eYd0msesQ7XylGyvCzA3HL/gFTNyqHItZ7
QwJpELlpmAleqJitoeWHNA6sTWZWDb6dFSrAjVpvJJ/0CFrAR0bu8R03GdnIm5KR
8DCRbrRZb3MHvj9YySP2/iILf3goG1bi6FsVQPzo7DoLKj0H6SzbfwQLT9CcaMGF
UqCabSzFYNdD118Op9pjGCVlFPxtm/8sONbChsUa7szgoSiuGAWv8UMuk7Ch2IGx
IhFEU2SdzbySJ1Z63byZRRuA16RiHP8Tk07gLNfqwDw8GCjAPNp8qM9FycVRrO9C
EDoyB8X+0Hh8lUn6F9x9sV5zFC1ylfn/6P97NyZ9y1zY8VVS0xzvZlbWjSct6xhe
ELYtE79wo9s57aiBERPio0nXyfDOgP/loItV5EmcaB648fxd1s6LVP6A4AuRVXGy
lyTjHvWf4/P4sAW8qIuygP7ojGajlQXLCfS0Y32U9W7/UUKRyjfwyrT8LwvMN9U2
Yws3IF+2HmF2Q7pRBv85rCMdFk6M+0KNmogpPLdsGEyKp+fgfLAdRHo20t4aMrgT
KozqK59HoKQi8AVmVU+tx8hfQk2PNFFyDMksh7VBrX9YyY9mNVV8i7tV21ybf2Rg
n5pBUYBqc6sZsDybNjgwmdONF1+wP/ABDp2PBexEakk+oHEa5+k1AyZIRztBS17J
D4oYgoGlnBpm5jVOJEPa/6QR9JISs2imRooBbzr5OPxbLiEPRY+a7zyhQiTFHHe1
zRSMumjGiT83TmvvMkSZzhF94qlvgUUmFO4ssiCcKrj8EJw33RaGA9JbUspuct69
9+W58rrBPsQ59fRAMqg8K5s7LA1UszRHpP2zPly3b7jmwOiUs3StdsEBl1fy7+pn
j+FcxSvjxP57cSXfBXyYr28/Vm6d8+k5z6lLetpG2IUC9MIf0/DeuCL2rSaw2l8G
VKIYYY8zqL51Kb8TvFbjL8tAkNNSoWzwDQZZRH7ZNtgBDvQzblpLTOK4XLvuxcQ8
571kQ4ZrCr/aDNyZHtDP2dT5cCP52Jt+6NlxpUtan5Y5cxkwZ9vDrH5vMAha+M0X
YXanN84V1MTAZJUIvCXHyURaYRyS1nPLfM60alUmD7012eJvqK6mlxLngs+rNLFV
FxyBSNSgg465dEXot8dDF+ZkBhESXmn/nthm28yD9lZ9xG/niy0VsQGvtY5rEqhR
k9kj384tVUJ2TOMZdVhckjtsLoMI+A+RmT3Dh7lkCkooSAWknfjWBD6XyGgoLUT/
N7fo459BtdVMRr4eHZUc+yCdtcKHlXr2c9bnmYT8RQsjVHkRiTTQ9LAI0pwVVsUl
7ymKIYnh3KGcU4nG0l0SU8hzaX+8JSq8gPFyvwfmeD7aYpF/aOTgWBMYOmShBgHT
RCYVFysAq6GoniyUAgPw96jpG1z90PrljD+mshdQm4LjP56G0BVZej6nnjTyT0D3
Ska5vNwuaju2iqWTWvJitm1IfxXiDbjuom/hM/hJ6UMC3A2088syLnu3YH1m1V6V
Fy23flavrdh6+tUlxDhKQVcxRmv17DgVcyHqZjG8PH1+7XL/dU2VM3P+0NOgftJ6
/GIVCJDrKo3jh/pGuupVKgtvfmKmP11dE99DX9NKHiPNlvjuqf2gVUXS5E4ASUVn
GkRQGztrKhFmRM+yDBteZDjoD/tZUUpOCQ4V0ziBCjWWCUJnXkMfWS/GFOnyA+sn
wSshC2XtYD+0u23cwfSGj/PT4JHix+vKBY6gSjV95juKIbKJIDD8+Ncswqa2D30j
JnyS4VpaIw2E5k7e5s78UsY9PQRN+dSUJt/eb1RX+LMxNvI36S/syL646MURegNr
Xpwd/DaIOcBfaDIN5dYSAye/rCjvr8B4CLPr1BMeUcU/vFhDZDyGtRwIeHQTJFkz
Z/k03pfz5KQlPk3FauKcDfPdgyy2LPlVjxD2XSSxryCeotLuUm0Z0j2TCkVWVgcZ
8EpTsCTyKgyI382zRQn3+VCcK9ePovtygpuP1KGp13aNHmI2e5t3SP1qUFqvyIKE
M6fSabNTCarVn5lH29qsR22LDyRu5eaEYsSfGy1Um3LMTNqJQuTSnBKxLc4xJyHC
nBBmmaYbR8es2wjmzHqNOB/uuh8TYA6OBhgpVAIkWr7LMTo3I/bGzBGlomR0b6QM
BWnTgEpo1VauaoW/2URFY9+qlmBPxhMrzeejasHXxUDjL7YzOqHFHRnoij2Cy6Og
iZgq8tydFC94pNcyX899IBiBndwHQhEPcp+J901DS/rtLpKyaNmXTpKtn7U7M3iU
Fi7GiZaDuFd9lrjWb+5XR7IBu6E6IM3SuqzAvTLDGhOuE+Y6POEpsxcLvBTd2EEQ
Ttomvno4aPiHxZ56PMQ6oAdU8sB92UEUcGmyiadiyuHNheSAg2swWB+OCjIwItXD
J05J6iS2LcRPXpJGWh/XTJXR+70rA0zTBFE2a9I6q99ESSke25DRp11nUOPQFaBd
7riJpfkmklPBoSN9RBFlqqVP9NXPQTeW97Krrs4JsqcsPuPGN2j8rfFDmbbHKbH7
tQHe5FU/O9ExuqEX4z1pq1VKZ/h0+Zo9l2A31DkRL36cMfX07xyydOlh7vak1UJM
j2VEfAakfbINLXia7qd1FhE+dm2FeAGi87r0HNTdCxu+u4sEoy+gvAJ37qYgmMDF
GnIH9RoEr/Ow8QuxiLYfs2R8q2zh0Do5ADOjpp38pkHd/ZN7rNDGB/ptnjxI9ykK
xV1JzcPa/bfdwoWY1oQHI8fdwAs7e3zmALX+jcYkhhiGtuUbPru0jQsdfnq64DEc
os/SsS71JhU1EmKRWWjFmLyhzhWPhg9mhXfLl5PSvWR+78xjDpQtiGjfRFc3J3qj
0L/n9I7RVYq+uD+FF2u3Z/RLerZCtwNYanTPWaSEmZMGUbaExyohrcq0sSU3yOoE
Z6RdsCqPd20d5puX99zpO35QYFItuZCRhzadH0p/7HSAfv47SvMS+Seyhlp63XwX
cRzoZxMEynvesDa7iXHTgrg9tY+r6Os9XjOkYBl9UyLx8pI4nRlOM46z+rZkNVdN
oxs2Qf9BknN0kfHT1fr072t+YtMOkHKS1DDuap85q4zIgbBKwFrFkb8Z2IWAoohv
LDW5CTNkNiBHzlMcwlwOkKTuVlTeFypM4qSJXC7XrR9y0qFwf9mFsURIgfTokqpB
bhOMNH3SKAWg1jkk0DAmZCTxQv0AJUBdW0eSUVGVkb36XtDnQSHNdHK4PpMG+mfu
z98RBJh3Sn59bZTJQRN9PhFJGM6l0rl908h3oJKxoPeN6wlA+JLD8zlDQyGaOPOy
qDtBUsqMV3b5JXF7CXAy/d9+IBsWeSXv+X7fqViW8SrfbDFesW3E/SCx1LWY51Sj
sHgwefDs6xVsvwHIo/1mWEVS2hiCWZfVoZrXsT9VKcGgWs9cxlpzfXnoJiSgOfdz
FMnk1eDDSYWQy4+hp/AEX63kJRzdTt4Gxfc2apy4OOvzvtzpNzYIna+yED75DezS
HgbUbN7QS3EHJBF9uHYHn1KYywXzZZHFxvZC23azqOXEKT/W6um7HCHw8Q/Iblaq
Uz9Wl5l7wVH91OTUQN6kkgumsBBfq8vLowxBBKVCgPYaqqrH3qnS1Ew7mxAI+VoZ
3q3XSddLxCvE/1FiARyggqs/099/pkZYnCtQqEbA2NZR7BY+bd2ky3wqDzTcS2NH
iHyrSiHg82zbWzr8/ZoJtI3gnrDgOj1YXC+EnwB9J2c/8jTwfftkC9ecqoeON98x
26CNrH3+7q534H6bLrnX0TFLuD/bFtywQ95M1OgvF1DSGWW/twi8c/uPl+4JtiLh
DfOaJdI9RGuxxzQd+B/S+1V5I5vYQt+/1PTtveBmmCjZBaDDkkg9vkjFyn6mucHv
BEz0gKCElFLUpmJa5E4Oc+Kf9KhaNoA16Cc7wcCG64nLiVbow02j9FhWzEw8D2T6
9vTMY9Kiqgp3dj/ozjkvyGwtR/zwxv54L7Hri1iOmL3CVtplbmaRupYdxjQnd4yo
29ZYcj5kXZNLU3epLajGD8g3mGRabSzN1s9HprZSs+QblGtHcg0gmkzTbFZCcGEK
xnaZfFJVLdVjj3CNBzoIrw4k+u+HB2cOTAIHkBzYfPEAssPb87sTV3SSnJuJsjd8
Yeb/tTBwXzg74uYdAoDD4jSXmDK0Sld/7TeMw2IYaXZ6eohHlMbcHgyuXb2HUUC4
A8TEpyO6ZUgxE3DUbCoIJIWheDQYpSVUezd6bdgEtLpe1dQOppgfcWqOV02T2ycl
8HzcEFbgsTQXEfM3Sn0830PjDmUP0EDZX1X6j62sUUTR4JXCcHZ2rUjF2wZ+nP+T
oF05W9f7kiSve5g8KF3Ik8fCFkN545VmcBlYYoJsDm3aX/Iozc3Ly35zVriKe56O
iOQfktD034TRlRccuY86lZM7V0+veWvyGasi+ZVIA6IE3eR96rc/4s08PPjCw5Tu
EwEqc8n17pdSllEr6dlQgA1mWLYvM2qcglgBf7oAMisSn2QNf+oTHO7BKFkbk9P1
q5XCAtD88P7KRwM54JKXwXzCINhsi+NrLo622vkdneOItSnnE42xxI+vTIYtuKo3
tgIFq20mlpX4S4Bg8D4O7Jx5OFfhHYKuX2hDHDNiOkrbtOfjLCGM/ww8pxZylYai
zIrVSrqxSuqlZMtIrDmMgjH+2gnGEv8LpcwbWRSIp6DCU0FQw8OZIxDB6XllDokq
MrJyD8YkM4A2zTCuuO6bvHVj8rg1Bq1gJ0GzIdu16O4BH6MXaz7Mh78KD3y12Coc
G7CdcMxJY5aBvlWRwgMYI53tcuv/V74RAW0hhZr5MtwuPgHANGL151iKiphyaVWg
KcWu6lzMRGbB89HH+ZimvevXaWgKKouL7NugVp+S9xvtfdYfiCealtU7nXly+hk7
s/r9VChte91gEfUT1arusiyW0uDhys86yCvPdVr0IUaWy97bUir6iyIEKSG+sqie
TA3+3KKr0vkhCYJl+uqPQFxuGBGHCCy6cU5Yy/49zBSTOnfikKpLcxVlQF8ujgmP
K3+lSbmEUSZ0NdJ3q7FdYYw+/gu7FHmWbPg/kpGiojEOebyFJCP65Cg1pq8Ob2UY
47pL4o0WuUJGJrEMhaO4Xm2yCq0rOLb/jrvlmhnDXRutyh4l7rM/T5MGRN9K4Jwy
OWxYR30gjTvpmWaysdg++XQ//oojYAc0hoIvDoj8An3+WX9DosjLYzFJEjP510Yc
l+GhCx4azeTfsaEFB1OigwsTTLP2bxWhw/Ezb6k/ccK2sTk+S0l2aYdwZt8Ax8fG
xrj52wVtLXbF3NkHgRgvJHww/cUxMUXsZWX296XpYtNNrSOQP5I0o5Gmmaco24L9
K5YI4vbFAuzPtDHNiaC0YKBe8WP8VEeF66h6s0T46y7owO7lcLJuL3lItlFgGpY6
ZH1WFS/fl9F8GeunF29bKE15siFuvoAc2C2G0wNd6kkPGZZ2ReTZVKtJBG1cXoSz
t0QKQ+mD5AMBSDgd7hQrzoNdu+96GLT1eyxCMRbLTov4q5E5b/jlB5PV/jWy/o5c
MiPOz7m7/mU2ZzuCxgq0Nn1WmA/zhnCzA6MdkEU1HOogOL2N4Sl/8N9Ne7cRxFcV
qEh/4k4HKileQpnhUFDrgFaCUDUywiu7ut2gbKq6hOH3hZJuUu7XB2X55UfvWzjU
pHSlV2Irh9Lx2RoSehCkb78w8q2Nzom6t7H17pjRZpKnCAVqb8T54zLt1wKJQXL0
tJeDzS8JOvhtALbEf9e4bS7YgwUJyTJ0V6dU/mLCvB22n5DxTR44WJf6MXeGPXKM
8FIdX9TTLYG4Gf0/NFmeMFgkg+Wgq64VuD7rbUIOYR4KbisrKEt24abnNkXRIEqE
0CUK6hlDlxvqLlJ8hsGUGhpKhKJHkAExX24b4WCHJREQ1XqHEWx4tpMGq+1gJeWZ
PnaEX/JTumxRMsKMl1Sn397kGvyE8S+M9MusCHmQ2aSNQRloV7pm3P4wHuH+xkJW
p/NeWcHJhJP06kSuTxc2ppTKDyq3X1QxqcO4TXnZV0XGUIwSkBZp5+Ig9CeRGpWB
D1yhZZFXNuVlvs3gemiYO46TfNrhOAoO9vhcA66DXgMps1qm5Q9ZNuNeES3Eokqc
wqGJsu0nnXGxkiH6lwrIRzeNUL4f4p97LpdmoPClEuhx/BnnB+mqN0+F8BPdIHRs
6H440K3D6tQ3z/WgJh1P1fVp3dL2DhfjhY2K5wIXnw0zXhnXuBF9mNZ+FZmPD1Sq
1zLXwoiS0XDYeyXCpKSFZtY4RMNdizehJk+jkmDo71oMKtWu7dtXc8RyRjlWoi+7
S5BXs3uUmAEu8+il/NfMpM/9CFTyibXX7XPEACK7aTtM/jQ0q3OTlUdPkYjnjVhM
LM5fdtsYo6LymqaSLtCVOcx7iVP3R0Juwp1WihQft8zkAHaYU60arTrZiaeoTLWa
wudA4I1S8Nvecw0iXrW9pTHAj+5XYaRUgOLYZYc6R5mmrWmwFr+nKqM33GCi0o6H
9r92N12JrR7rY27KLlbeci4E/Di9TkzB4M/9Pos/gFvzRujzn5UT+F/l9qtTtdzK
FaQHjKeql6iyIqT13medf/1AacKWGOYjCr1ZPPmVc9GKQqFLRxedQ75fQ0xgJdGK
QC0TT93EB6I5trweFiZUsu//tJ0KPj/uGyEtNfw/sUx3I+mTc287p+aPv6i9nU0i
yR3UOQkXFKHUXo8dVmF3Mjpkzr1KjBnyoT+teU6ri9EjCTPm8ZOoSHVyv3sOINY2
Qj69IGSGZUyPA9ZzZs+8Ug/a1mO+KS7vjld0Q4ILLrAvvEAojXVfe+H/kNpmUzVf
OYlc+O4swogHNVLXCcOof0j+r4Nm7JqAzx5CiOwBpP40vWcFwnHXXskwARH7pgu9
Sy41xzQmANM7XB5Runnd4bKphoLd4Lp24RJ9j/u9Lto8/LNYB0jAr447gJY+fYpJ
83E9T/9VKsQnbIT6AcbImr7DJurWNJeZVk7g2SKPCQBZdXiyrMZj7/JLvyP+8bew
z/HQEM8OUINUEp4XJXt/pjhJ9hA6shmE+cWzY+M3+1Fgm44xWECyQcso/vkZ7FOs
o3Z4cCoeW3Kekzhb00nN8AViDnt6b+y0uZ7xhrQ1jYmpLUmLPv8luiJNU1e/d0Oi
R/WevCItHmv4gzkWGpy6AVzb00J2uuws+p4sV4VfbBslUh2NgdFdd3zDxVzyfo9A
Nkcwtq1N+uc/yfA/0J9gN1Sx2Tk/bFIzZr/2zGdQvGo6pcJaK0Wm/Yy2jiZAk26T
1CDkLehX6B0YX9UebVXb/znTicRQNGG3IxaA3SqR/XJkZw5piiNl0AUC2ut5qSeA
YlU8Y7aqhcRmDoUizXVCOs8VwaaS84Uw1iEsHAXSnnvveq9Lyrdlf/NkXifDDDVI
/3vrE0sv0Nw3ewnwDQHu9Zq6erIb//oTK9gMyWvBbC9q5AYPohdL0ZaRhsHzLy+i
1fc0ehQffm+OsVkxMiKPa+ESbLWV+grsMuz0Qs9BW+m+nSHhTFIL9rRzZ+1HFmTx
7EKW+WoOh87HSE5C62WkTVXWkGE+WeexE8kgB1Tsb2Q+mZ7ZT18/4otPv4DFnW5A
tHrlGD/3F57A+7O1n7xUcrAkOOTUwr7M8O3Z+x0WG8qqp4ASYi5HMIgF8AaBCngx
T/M3qamCV08RE46hUTEPGlKlbdE/Ad55ppfaSye7aNNc92A2+c9E5UBwohiHXW7c
UgWWyFI4T3WiU5V7swDxM4Knr3gO4uyl0MDcaezY+0TvylIefSJ1n6bHzs3hKIzk
SM92g+iwdEqBt7AAMORTDLHByAxH0rvrb0co/QAaQXS+0YDi2EcWVBmuuM8aMgsS
pBVPreVTamR4GPoWiIWXVruRUrmUI96JE2VMflOP3szo31Utwl7bkLLdrp6hOJSw
xxU8nyuCnTvwlEVrBQApxy0LM641F/BOuERAnSSz7yl9S+MPplro4BogSw2Hz1+A
n8Vg031wXRuxS9WHZy2cqDtvNqf11XagjqyQ2yndIQXwlI0nadZ3FLUckjaxQNZB
ZIWqhMXWVUSHGlT1EKfDO5VktGE+XMq7xK5L7bhWnWfe8kL3C3dqx05SKRQT5hXO
6LzFotcPFHtzQJ0EvsPLp44xVIX0ByP+XvV5Ia6a9KIKc7Mwc1y9kRJEq/Ds/tI3
icMkCCO9W18/6YKUZ7rlzmszDG/pVSs94VFWMFt8PUpBPk8bCbRs/6bTZAf/+CTH
GoH+RziJyPee7n2q7d+xKqlgKQ3L7XajlETgQoxHZmKxtQIWz74/FLAV/lMcUoeZ
76Gk4IsL5wluLY1csymgakEEL5m/O7JJIyoC6Fy9vpZjLe7bawpubCQ1+6hOe89p
3DHOfgbinxg6ssYutxT0U78LeD+2tWLxUAdUlF9ftc/K/h3UrrINuKRivguxuFUu
Gi3P0jwg3SxPaLpq+EBgXnpddpz7NjXfhXpn8NliKmXP6pYDdRJcIN4S+ltZpIUn
rSEQXWU8y9TvY6zoxw/dmw16SjLvOzQbtCZLMaIMhhrlXksxVzQNiFRUeFHiZyUR
9BejSVLlZ3oFKlJcNaNRfJ+QLhdaW5in67pThxYpRT3b1q+Id8qNnNXfwbK79ON/
J9rL3mQJYddJ5tkstDT6FGipAgybsHuirCFK5dQci/SEERdwnruNfJPAfX0fVsAT
sMYE52vtvaOBp6wtDLZOi9Th/9hM9OnmdHGOPHOA++PE/8yn/5FM2P42og9xze48
jd9t/stHsYx0TRyD2LAUhsxcshTKayKZWUqXVKM8V6zKHzMTAHMCfdV/d7hYD4VF
5q65cLOaUynafySRTueSENQtWwp0qKCiV8gmWiM2Im4AsqBXa0MJNGrH6WN2jN+/
9HPVwpvHEFLryVY3S8WOyqLKNs7VEa/MlNBRCDwfCfUPRY7gKB6E/6T0Ix3+NUag
f5Pd1Ag/Nr8qZA+KwMbGI4tbZgK1lfx/KxAzYdSRzbmkQqXZCV4xYAgFeAQng4Kd
Iq+L8zbUiUXEFzDh9M6Yz7gyaMVlCadLm4VBej8RDRb5GsVlhxk4dZ+Oun9zSt1Z
t1gjrU1nmt+Ov67JOgSdZhzzjvx8XDIygciMHQYgghEP1v4ReS4XeAjOBxuLnG9g
ecXntkddRebQ5qZQaM+Gm+ZVPhG6+S5Oh6ftwjOClgQ0/egYdm0OUeA5HQ7QkzBS
ZmhBxhI+BCaLtz3b+rTKyNnusjTU8p7anA0wVHPeB+C3/w3ybB7IuCWx0RZME4Qf
DtP0nlnmcg6crrCNaQ6gAflFzVd3HsGzykmlgGGTALoaMZNc6atxwWv+570FEVN0
wvOIXe0r8EReOouZcKhsjgq7a7kTeOwwminI0iAovv9mOLg9Pjb+yZCtMm8ey/WG
VTkPR+G/QEUS4cOgJXXz26tDOXjQ6ndhtTCxV2CC9f0rLjDFZHvil0db97K5Gmsm
8a7myvcslhzIeZBnozQziA4d8ry9Ozmf0vKMVDZVzRwSJqPgTnPj0Ig8yJfWK0GU
BCsL2boDf3dbZAYP16ygRUES1e5bxy8ZmpntKKJqDAmVqg72C1Fi38NqiKchCHiQ
Y7GRnSP14YfhugG/LaOklm1IyV77grRw92Q0aByoO6feDb0z2tEzfdCBHSWdvPH0
QD8oHWwfjQOLpFfHneP0CJ/uBlo1s8hdu97nVWRcyL8RkoLHM6TkuIHvxeC8hYyw
P+qoWjXCNm/Ho9NeygeiAEsoLd8Q7Nk3AwvSENrelFOPplCJX4FQ8POSjOxEMjVS
b043XEwaVofmiEZTTT3G8scni2lQwJwMqlG+oi/KOoNhczxSpPPREOkaJYfycrns
HmPkRo+j9OBzgAOTKLTZ9L0UxeBODSRRhArJpg2SMPHQ1DnpdAVnVLZnNJCHkswL
gHY4z24OrlL8krPDxJve96Pmb+jSKqmPveYIeUR6cTVNxJ2XgOwYuy4j7QQFMom/
GdNJNG4pPUe7hMyS4prS/mnEk7BVzGi5U+IDQP4mb/gt0snScnIDGv7KWk7McvBe
NikMDrjJrAxNuQQdQOP2NQShURTAf0wxEKWcGO9SznSyW1eEOCzQNKp4/TtY5/fN
IS8YOUQ93COxBZ9kb+2Gl5Owq/Ysk1ZorJEYWoSltUX2fYOam7WKibYN9b7ZfK1L
AI457l+172KV67AGFkBgQSF/riG1JCOYYyZd8wAEH9P+abLetjHgLRQEKa84HbxW
E/+wybWmMlwdT8mxbuhxcKxuscZndn9mJbz6Q/R0ZouJjQoYEHOumtG/s+4Xe5mP
rTDQqGf/zbfm/CT6BM0Hux387p0kHaCYtoFp1xFDr7yOlBOpTnh9nDpkp1x2z77X
CtfJ8edOX5/6Pk+1WSZPha8XC9+/WYiSoPgDpAY0fo8SLm05wF0o1bwOcoXDd5ZV
JxZrOjtNhKBObtBLk7A/WPDd8wMf1WnGgZWo/vj2Hv51pwa4thyKAoZX1/XMBDNQ
eLcTc1txfCA1dI09WICbUca7kkvtcAxk04TZl4EygR0g/gGgPpEzqoGozcfxcVv1
LWg3St2Pyw9eSlvzxpGm0nPJy4FUBAIZq9aAktkLmTOdDkb0Etbg5tncD0qTUA/V
ezc/HRzffYXJ4doSjE43WGkC6vyoEY2o37JR/W7SqgzzQGE5+tdqYaMPXstxUba6
yO2gfIg5O61xjxCypCEOLmTTDgLUjk11KPnVxOwwZX+FdZrGDNu7P3ov6QjRFQGo
BdVd1/PsyLi+Ew+/1njJ2UAMZICkrxKaHu+x3hOkBUBRADdpdRQoQL8uLz7si+i4
M8UXzTTU/5/9WUqalIXW4LRpiUNUn8BZRl43MyaKDNZOXo3lBRMJT+mKpq9OlzR3
GlnLS9k6mztUt4uOmVt/8AUFRjR5BKE3IcJe3ot8c8OzOsvzYnuBxU4+cTJVS+fJ
LvgUwbA/kQTKmTsSUSIrTupCIU1GMZqSAayoudODBKwSN86/jtTzsMjaJQgnU02m
U99Wi0pP5InnhsX405jyRyK6QuTq0a4c2sosycgrzN3tbIip+y/b+bqJ6wGgxJCR
glpMeCklnShLUbuMi2/zV5KS0rKq7abB2iv1zSf1HL0wdk3qTNgo1VOnM8FRwOlE
z8arvd7C/9KO/EeudgfrWme1RpCEM/PAIK13myURlnUDivv7Dc+Mnx4L8N/DjjPs
G8sgfzAbzLOMT9BQwEknmHSCi+4Q0h+vrxRGQuUhQd+7cJz3xFpYzg2FN0u7INZV
amskY5DCaNArgPVd7POqqgpGPOpGUbsBsIRk7jaiVIBAn1OjVVza0l5F+zdC1zbG
aTiATGJwQdC5K3NOs6DFdUQ2am6tXQsMrnrSH7L+MVaBqJ6ytaGfi+XymCsDCLZ1
um//ZKAQfIDjUAMhqjXSugAmY1UPUtNbW2OfmSHlAtHhxIYRl3LnmKa036E81Asc
5HVn3Ltusdw3lcoxF0QyfzjRZw+xIdXu7Plk66D/Bb2CTkQoIHyltyG4swOr/rCV
9sAhWLn55fn5atRqZptDv7snbIvHTsZvgwCMLi4HiePfPDNLm5EfjQ2Bq41n+NgU
fvWCBytXeBQN5oRgeS/oVtgs3/oysCMItbgmDzq0z0LRzU4P+DZ1PJi7WyMHYTsF
jps7O2F9U2PU3Xj3awv5hxy+KqjTkbEpl8iHTrO3c1U9TDTeuo1HQ0tdDiB9RwZH
HRUitGRxW51he4fa4CLtAIEzEfqOcH8nPh2fvL1RwP5VdtyqCp/DG90QmeXYgTyJ
uI3O/B98FvGKA2VCCKX3tsScINBn4AP4kwF7dRA4Cm1g1Jdv8bIIJDCjEQVVYT90
L2/GLwFwFv3wLyNEVWrGbhb1T6vRwVI/yEOiOHzNv3uN6uYIk3Du+5gcnAVEd+mZ
u9jmSE4xo/thdqE2EQFoHe6/gvxGo2yam+XtUd5+QOLBDk9qruRsG997Y5/VqP2j
CnRc0ZL9qoo4AeltvvaHJMH1GkhGi+3d4fb6CrI28oNHyNiDNPLDtYWo6FAF51pV
GhkU9MxsBFsY1q3ekevinBFMK7PtuPlcdQJWmfFZmLVbShGhG59EBkt7/iPPUPga
hvBnKaSnrvKiLZOeq1dHXNFi+2QQBB68y+gry5MhcCcUiS3LmguqZoFIe282HPJi
HiKUHkwr4jzKf3qSaQzUFvb1ZMLZ7T59V54jCpHwq8h/mzSOvcTWe8OqTvRudh+a
9uLu5YhUXxda1y/Qao/6rRTmP9icTUH0KnHZE0Z7rAUSi67Z19/UTiYJlZgICU2Q
GwzIaG/J21x5IAlWzhX3sHrObAo7DuVB+Qo5+ZHumg7X741xbvAkcxGjY1jChBft
M8tv9tB8HS2xA8xAekCdiqperhW0v83kGVFImt6SnUMnH2zY5PwPrCx0Le8KNyG9
RA8WLwQV+a+Sx5+lqw9ca33ZL9mpT3XwwXpx6NI3aPOyVS9hWC61JVAPOUzENZ4S
NTsOaPfOhHTcbStThVjCHJbkNtNA5uTvJ8AmKreNqL8889TAHxtJ+ULTHCN4suoY
gWOJRtQ7J8OMhaErcvetS1YT3az9PWBChxJWDfUhtGdCUexUeH/Ad/gBn+OqIdF7
5LW9loowGqYDqZgyZ2Vt7+2p4FlyoGb4EXSjsylLYps90RTtRq4KOeNNxvLkFkjO
w6BXBfNs0PAao2vk93rRzZYJvzkyVgByJXY6kqTiR5b5AUaQtgYWh1tMPiCspKft
EilLPtwaxCQ+PMq6f8P0u9LZsmsddCZPgCmy9XRMbKJsewQv0C4hhBRoDowryBw3
UhluTXYqdUF6TbM+P9jeba9/usC9EidivgxZx/sSOKzFc+OnVMTp8bTteUTZHrOY
ynRgouOrPcd74ewx7zGooQzaGBHl4WnHFpad23YpvvsxtYBHEZaIgYoe/aw13Njw
3bGfGtqEeow8sLy9puas7sjStcVxqtL7mgHErin7G5TBW4Lc6XO8GVE1Nr8h10mP
B7sw2CqMUbEYE9W8oxxMbh7NF5SKDLY/3UplbMyHmTtwOO0FI/Ex+rCMzGgY3hUX
PkjIbIV+SHSMd33FkG50LAaHRGMIdpqtrUXYNiorCifrsBzmMwLE8/GTFmkJV1eA
IL7tFudXxhv+FDkz5ABXHPIuw2WmrY/9yN/QM5SqKWVpIYbAiz5yTXDRMBsrnSrl
L6DenvkYU6Dfz+IBKA+sDP7jNJPHr5rslxOeBDCpyBTpjQ+5iKaVgstCQhJGet8/
y0fvQF5N3lJviskMzy8vRbSjZZo4MKU1YQIsYfES6mKDbzl/tA6YEfrc9d1TC/r/
L7l/9DNsUgs8VTdoV/4vf8LDxuY+pn6HUntUoDQT/7udaQHvuqbsw6NBxEXU4vEL
g5PzRqlyYmm+xLgL7UT0l1UnfABrCTfzsZbQL3lmIbYsel6GCTwC+KeHPfz7sum4
jpa/cEQihFS6YsXmhrZJm0A1RwFQrAUuwgG6IX7GIjhQ2WB4LHpGocEv4NMntSOA
gUIQG5UWjtHuVekAHQggsTYlUqXryk1X8/Zc6QAkj7F5KdAAw2l8vx300RwBExUR
LQjxXL7U2YEK67A7yU70jOVKV+I5Rk1KCxyL2VOvqeVDUlTF0x1iEGen3gzIcWDc
g3PVP22Tn5s1EVlDlbE2eCsgICj1UFW077MjIpX5F215ygpoNcRyswKESvYQcVsB
odFBhD+tB1Z90aCR1Cb+6CczcGP4vWdKTBViDfP3UItYSG44Qe/OepIOV5A+5tCx
u7K0U7McTT3JP9pQnkJF4Ih+k9fhMMXAKzRKAk2FslYopy+2/GkiqoZFxTkmT17A
+BIxXtmBCyOv821u/bjwJEI9t0hGXblG79rOc1IE8h0zxEQuCYjxBtauspeDV5DG
5d5CjsLoEc+fo8DODiDRze3OIzWa5Dwqvhenwfd17bcXd4PvpbLhlAUzoCiAXBRp
riNZcrmAShkAPCj0t9w8aVsJLp7J1lGiJLC+St4V2VSJYvauxyf6C5TvDEcGYJW9
pcdKDElpRBsJ35ZqXbCFENcpigH85SWILdI332IbpBaRwHyZz5Q+YEnzcpyoJMt3
89s0OQrNbP70UUPwj02AeT0L7n7WK78gXNWSOR4WhOhkKTS4CYbaq0P/P9hJdXGm
ZOVPfg8G1qcHfKVfvqzoATEd5BFqokTpsBvW78Zqghrqf6oE8dmy3QIyrB2BsbAc
cJGDkbWOsDFio+4MGKlnaemLiipxhE3LuNYChkj5pdJm4zEQ4edA8fusFyUKdN5e
oh0bJtDmpgSGzwS3X4B/bvUMu/JawhrbIDKfaW7ybzMO1UGowY97yts50BgRXh9a
ahH2xo9X8uYfTvENQwogXdSm564AvWrq2fWbUkZkHcNT9eGd+YJfKD2Rx+qwSUYV
Oi/JwAnhoGlmywsDEgdb3atAEVnrxr0QjZlbjLGIP5kuA7RIC6JtXqN5hiVSqRsN
3sewzR6+77CbrCn7zpvBZCTh4uvI/WJRKInzinLO80caE/k4JnsRal1LYLxIukoo
PtS8CLREGeQYxvN5HNI3HCw+9QV5/v1jjozlPMwzB1LV5201LJtttduA9SM/1crS
tG/rtA+qICCUG5+RePaTFwnZJwfYT1lLg65IIDtJYdif2ECiC4EjZSM1p5zYlf8Z
UhvRkJaoI77pzLRcsAV5t+j2mr7T5BgkECexxQHnkCugGIlBmxaRb/yndg4ygBjK
zsZSZfevJb3ql9uqWSgz/8RDMyxM+djWF+AQy1Ow4jfgTJJT99EvP9Vaf/mJPqJu
OD+LvO01t4RqOQabsKj2D0t0Cc9amByzKqw0UQb01+4/CSZkWakgz3h6N10g0SWf
ROwP4SJ1Pjj0E6iCFmk0KSCwhm8ZmY8v0dJVHfFBjIEaNqDD6/BI0OaSVfhMW1jB
APOevAkt1s9u8QxOvr9E6uW8Xv6Ov/HdJ2s/P2V4GrwlWfwuwnhdsz3uxdBTQT5z
f2/SH+CL7g922uRJxUM3T5T1hASzrWSy2kLUe+68yOWP/QywYBuCa6WfF7XiX7+a
WDaZLzBORSCFx+7wDFhuJkn1ydA0sLXbz+5YQY1eRx8xBOkSPPVWc9swysTnJgMO
C2YrFuWzi8lnce5coxGCfGKUS5nC5z6VKSyAyYKSsUQuPXrWVM6Kc2yOXZU883dh
baM6Q9Lt1VENMW7+kK5t4qq5sn0Kg+H+MRNQnhv3BujLP2Ph5aFB4kggKY7q57om
CiUGQ0b7rahNma+eX0dZ76SPV+4v3wpleiGKrvzUWvEENKBhRIlc6lSISi+Lpoch
Pb2EHk1Og+UTZDO2bWF/RoTGW6QEOoSlQtSrBCuezIA9SgNphUU2fZ/yDbM6noq0
xg5vT0mxApkrpSyGH2cDsAqfBsI6aT79XWD6oeQQU0GWwpIIBKiWFbYgWPsK2D+/
1MSTH8ZnmGrQgT9XsGVvEpAnROwpCIXjT8OXPyfjZYtXyZQxqZUxZLGXpItQg4az
Q/+302b6TCV2xREbEhv14AivSROA6O7lneW2hI4lQq0Z8mWd8UgiQm9lKV/duVNQ
81ZT02K7v2rWCuxW01WpKOPMncJU7GpeU4errypYgmfyoNKbsYf5B0jGyZ/Eo577
JuDsf5jibJYJx5nuBBg1XTUZYlJdKwIyd7oLDgE97G1REm62zwXAuOu7/j7AiSn1
OOd4HW6W8/pnlgw0PRFh15uVl4whtWdXfB2a+IXF3w5iKtu9JzRB0Sj46edfCM4P
wl0UD3+SlbmKAkzAXxkr+GTRtDGoGTNLfhxmdsaOKphVrMBRp6fWpY5YX/HlGImY
7sdK0MonXq3v6kWTO/TCrwxB9qmyfK+sBesh3pr5reB5bpGqF14WmgSnXJ6jydA8
3bBfrH6bUkWoRmbZ5aRrhNQ64evL+jPV7z7UaI7sGZQIULJ12FnUrxCx4LQvRVLs
ZxjqrVcw8FPVtaWSuyzVbrZKRIzUI0iCYEwJOYzohYioDS1f9YDupuonGuIAMVNO
7Eanx7P7kYuRZ+a0OXJt5w5Yb+BDIer6Nsyb+PC/ghDx6amVhxEdpyi67nSI0EzI
KRemSjHjJAPrFz8aFoZd6S7LAwcobyvCEDxnf0fPF2SFaUWY9fkZAc3QgKbflKOD
vgsAk7rwG9NSmVLYdag9tXY2YivdJu0JaVNseFeZTlU/u0X0XnaB1whq4i12tzYn
OCRJC2sVII8YFGCXCHFBoIcGuHLwNoiUC7j3V6CsPc4dypw+nA4BZmEezU+9aLP2
rbv0oCO6psGaZ8y+3UbT8h0GRTKsySTF1S5PNqyPRW46Wtg+fIR4KRtSB6R3QkgN
XFjZbn8/cLRFu7yW9Piswgqhx7l7po/pQFDyp/DlK0EmUV0yO1cKJid8R7ESoEd7
Iz72VCgaZ96oaroeeRADfsXMccBylId6b0mZTdGY/qpzZn9/GYSlWdBLYrgMnfkh
jONiOSomQVLA+CtfOYd0xqbKkzxndnDmtiBttGokhkgVv2ofFlAYLiI7bcBfK026
PHDAqt8+Du8+SUh2K34Ck+xUC+SPurEAf7XvYq+N6UWuRpbW+TTn+i5rns5AH1BF
dmIMBNwJ7uyiqfylaqvkf3V/XDLf2OmRVYQe2OMk1QLv1Vgco5rm1M4djcW2pXge
Ihol+Bg5YFgMZp/ZP1a1AEJqBJYaCrzoryOg/ZH6KnSZpQ1kbPlFowVLxZwZM4SB
lB+mbu1JCqzkfY9iNr5dN/tQjpdFHd38uZeHxAhfZg1aEWVuvwWHq0ov0gUCVvpP
4OUGERjRL8ocvGiDfd8Z7ljnha7odtv6qnNNMIX8XqGbVEIRUGzJwECcSAuUVxYa
Hq6mCK6JCtme5aJrq80qQEaJbKqrJyEi/l+j0ruQw8Q7ZJ5eVBONJNmTxXxLuU15
v995X5xi/xY3/bWgARTJfWoeUPG5Xdnhw6DW5Lb/7wUSXAsTlgaaVgjmm5jUqrvm
3ol5CAnsV9rBf9+WNZ1ePUK3bl3BZM3fRVNcODErpnOvf6V82rqyx8IzDjL1Kq6m
ahX08knYO4oBi87Z1+GLdCARdQa2avdLJiiFIMmkwEILE2dELxh/Ly1c8qShdVLF
/pJWz4RaBxsMpRAH5M6bUUWbv2RxiJh2EkFa3of0u5+2M49d2dpWaHLP18VsBTzt
HnzSanklZvb4cWzNlBGnOniD/7CpHMcO7eZeI4Leqh2Q33ugWrw/i05qCJvpKn01
hMPKfXYjloULsANiikJW05PE6V7fUNl7Y2+YRfkvGU/V/AGP9EtIba8sPEXyBlJ8
i0LrgxK6d7J7Vq/ajvla0GIdSIqBHSEN+p32/2WtYuD42GDFXwn4IU5Uyl1hgEEe
CNtMcKeiD5RS+is/Lhqelip/d6SLrRRppDBKWDBu8m7i2Sq6GLE2H7CjS63YqbIM
ShuZhDLqt13R+L6+0+YdUpm1Ne9DcM/6zG6ugUSmbLzLD+/RxMxIwms+gDe0D7vy
sTf2HRDg12QmedarGLbk7n1tmBPBrwT8w9oZMr1GFew6lwiYmoCbNXDz7WtzX0Pv
+2lKqUkw1a6KYqyspSyY8HwmW3zKdB96T6GuXCvAslzV2TjZbG6JfY2hNIHKBkZ6
AFTuEwJZjPjn0Tyg+bSjgrmWA/WIhz/gKVL/EQJ4sUHwGA2opY62MVIYvDS1KJRu
8acHVQkO0vUgxCLmsPBJLehqe54Yk4qza3f95Djv8lKEUaqbnX9JWJsrW9wzcLNY
lPykQn0pIQmzw2DFySgHz1aQUTMxlqNTPlRZSd8fjcpzVY4ZpmUdMNHX7MA236mT
FhxQVvSQrWKdzLnIIa7IW0ZWSsjAo3JSAyOC/RPE+3qKEAti87wpa9osyfG+H/jR
EvZDqfBZ6d1YC1itAwe+rSD1pf0nSpS+mKD6gdFIBhG7sWha+YWY8GhlEQsP4qO1
Zjc5MpY7vYy8U+abGrmQQftQwedqAsWfaC1ejQqkyAVsomxtzYb9mbwiznrTLaV0
ASGQ8BZaZEWe2bm3EQM7JXrno8gMWqWvnvQ/aAIqG950bA0Rv+gjRPXdJFuJYsQc
T/SHDdFltr3VO26r2DxGzeFcHZ6kWCbQuzJffQLoCky8vprLOT0Q9JeXuqVoPKu1
+oInRUyXl1Mi+zDWhzltZVfcS9SdzBZ/tkFUiF8vJXv6tk+bfAcgiqj1dLJ76IKt
8Rabo1p73Ko32KzafymXiMlKdODdKh2rFQ/KBCKFAD4J9Nw6rmi+Tr2jawYGiVLu
Wvv3UDZN7oqX+Wda5GRd8lIdIWGmsg+gwZ0hbh1OEFlPyWJfde0Nlr4HEZZc0+xe
5J+PpAeTAjFFguOr8cCantMekzSmAE1MgRD3B3eIAMvE0lX9DUx/sn/fDVmrxoBc
g37OkwwXo6akAOes7YR4Fk/a0ZtdttP8kLOcOYyl2t6pGtYkShtKHi44LD7RmQ+c
JmB2NfJp+Ez0zWmvfigzsyt9D9T5Dqod/yotcKPcNn68xXFO1v0rh0eUfLcGCGGd
cfqQrPqmMl7Zoq+8eP/3cetJRAJfwjn8SRFKkmvCF1mW4eKStQjUVhD55BDf45EG
Ib+XLqrrYv25wfoaGGA5yJKWW2cl9gtyIgwfWahATn/dR4/K7lKWd5Pgfotc9Ai1
pGSQMBSDGZZbFyfR1+3diGnIwyLoieTKDYaDnIOMS8T63Pwz4H/DyVvl1echGR8S
IEy1r0lDtvm9g/MkxDMogvijr8mA5/qnfrx4VOAkln3x5KTVlQ4yijQOz+WXBxso
OvKLyTeahQw7zAj0/mBHVzBAJFiEf0k6TxND3kwj1qIUAGg6IHiEQXx4bsNne4l/
4Bp1DnHGvrYsOG69oGTXjIL4iPjHosPv0C3mbkh9G743UTWXMAplYvV3D1xRj1N7
zSGZ8fHGDzMPfm0f/Q2L+/GfXBSu3jVgTYSaYq58ggB3VwnIAiiemHjFTQ6M6rFr
i58OGJLEsn2ztkvf+5arD04s2Gq9M/0UVkBy3/gh9ch6jSR4Cd+Qc0+Vw/6eRq2V
MRFMNyahCL1HoWZOQMo/dM3/n2n5Hza8eZTZmwtPQwFMiWlsE+8ONowdUckHZ9MO
krdOKdpUBwm/7gPTcrkDNSj4XZqX7LUr5Nj84dTWaLZc8ZCr3aQ7b51llBeUWUfH
Wzkg1CGueniYq4bKRb1yWfzBRTRvMP+PUC/cXJ2X7HiAUU7cNloPf/1v5YNLR7vh
yJI2C5Ak8ECm44O7itcCaIbVnL+O+C+gIbVe0z6hg4r8rKpILgFN6hv4nQpUkNvn
ovKKekR9pZE6Pj87QxUPWBpVyZkya1de9Q8+A8z5PGJUzYjm0lTZEBFeBB9aCyOQ
gV5EFJ4Xg4pR7BS/BbzXnO2WjJGYnTfulaM5JP8i7Jn4bMWuELc6QQHSLjkaBJUJ
Xct83GZN9PrcOoqjGpKLQQkUQioTalDj9X7DNPAhIxpSwLQQv7uRhs3DvZw741Su
cFcS6UFKMyNKzQu3anjjKgcsxpqsnUCfPgGqdfP8hOrlJduietaCz63ouXQOaoxe
bP825tBXFCSyN7rsLroAMjvbBIJ9Azg8QkG8UCd4fnrC+ZFzDrOqUYiufOJ9v3ky
pCgble+4rZ5V45cSFg2Hx+40gv0Pl2GlfKRfh6QJv7yfdgNU57xlgjc87jdQloGN
baA9+XEpIcZU0+HvN1CMkUrhv1XhRPvYGeZd21hhtpJ7wEF/TTP90OVjk9OSdL9Z
T49oRLNgAL2om8Tt59AAt92Ry2P2IIhx7Vqur8p4lYBA1SELGyv3jGQnuMbOm2ys
f+/82ykdKoKKL6UgQMtpYfyNIuJYRckFuOS/Z+AoKNHscl9H1AYkRsHE3hV5eSNM
RnIIVz/CK1b2YwmTNbXbZOOfZr+VRrvhfS2WfWUHx7RDfwRjWU/mD4sRdsd7aDud
vMgYq9Am5c3AK+pmGYvJDWN0ZzI+9y/zjRzanB9cMTJEgxqyadurUYoD1mKSUkJE
3al5+rc/dzEcgkHNklf2/Cs+VCEk/q1PWyxkDQUqu5Ku3Qmwp9SxjcM2zW+ZDtB2
1+Gm2FOhQjxnVLJMMwwPpQCGiWx60qbDu95bmByuq0yrxFXJvI+aFj3NH6Lh4rfw
BsgudlsYNiixCfL6qxkVxqKNMlPbIqlviUCd2I1AcHPLz65Oo4eymwp2aGpCTdUW
LkHAfxYbVZhVVqbxCCcwzy0+4wrFsxZpwmeqpNqzCt9bztvvStr9ALBkODtHlM3C
2gLoEGrVUxohT/RQti1DI8ziG7XhJJkb5bqO9ogLIetHnTouw48sB5sdHnf3+mU6
MJ7/bXei4UKkyFCjTf6cYNNKTmqTPxE3qYIjQyB+IGeMGez392wVLW1DWZAxmLNs
hyly0QNsG5iWZLpVyzh+veLRj6Jrgtf7ImSOw6rd3h3i/bd5MmwIX0YCTYozUTig
7okHXPjoZDeEFyjIzZV3i9mieTEwGmoylBQDZhVK2ssqtmukq4Z6hqfxk7S7g6YY
sBZQcgu/lYUoeG4vzty3fYqr0u0Xy2Dhfu7YmlduDNbTbbM16gHKaYpgJRlnakCn
KSowNsGf+If5171FdduTtU2jDEQwpdSE5U3UTs+obAnGyOuAEXZCqrChE5IJYVdQ
WWUy9PePqMJWMjSpvWafoKbHU6yL0rZw2EOSPaSKElyT4LzYbXf+ohFIWmEny7Nl
JQax4Deu/vjvhFxo1PuD6ImLRi0jDJwJGrIh+PbjSYgFriZiQlJU99nta06ucnsC
dmKyjHbdAtLnBNY6aRKe0a8KjAS3tFqErfbx9TO7S3woKoKpawbIgrMuEclwmfII
NdjmQ9hYLRxB6O66lLO9qCVh3YmCDyvDMh9KhotRzB0x3M2gtlp2D/HVrr054kZ8
kvC3234Q4V2CakmkATeCplZ5t26eyK6D9RSG3vzepSuxYeBVz7GrVXl+fF1CXxRp
e48NveZiRtVp/D4Sgxc3KtMWchfI1uc7c5EITYSWEnoA0lnYH9an0VVCKANFN+0S
KeFjhEZeVZynLT2aEddNULvWpu9JFPQYBmF9OPmh06sS/cl6cTihoVpsLInB9lRD
TK+4Ew13cwvFoGtYryNpiv51HjoYA/laM0Bikq112qXZdQJW3mhnmWiM5vlFm/oz
v7qJz7ThtUnsGuFZ4441X3iqXpuJHOg1tzw2eW/ybiOYV6KZLvoZx3capvqURpGF
h6Za20YhBhUl79rtrOL7ZIb9odcj/2j//Jt/wxlu3BJp51HfJw5ambr1hLyDIAgf
hskqpZRsBVWzDgKkZ1MRJLYXUSVO+zDa6f8DkH0fTuLYOW5KK7ZbmVv0TJDo9rvO
kNiNQV0D29V15W0SfJCYk5uxKfOia1yiv6XfgQybX3XWwN6oqjgEpNqJCXVFK6ur
Ldj8oFYxmvty9sGIIUgzGjYXY+KwFh+UbxHzhKvvQ42Wvz7XkJndtunbt3p+eTta
pWl9sde/lNPiTro3jNXOr4k49AKKU/WU1XBn4v6GDJuUHi0pJUZoIdHZTAoP3Pru
d3ulAHDB5lbBvQZHXvO6j8xNxiHEPbRheGuBpesRMsx56PieWjLB1p2UElK7pPsi
7W41ouS8YHdLkoy0qKx2Micb2VOPJ3sszq0VRspYQZUC9rzy3MCgxvET5PodGWEi
n0MNMV+FdNfKECOC/Q7Ltyr8e57obDONCqhIFDI6n+5/5Y83h/Bce+oOkoHOHk3F
ax5WUe+Ap7u8+RA82uW20VcD8y2rMpsLFJne3xPol+GuKHtlK6Mc0vhJMoCDs3OS
SLDeJqn4AqppslbVtE54DV1k+S2xmjKjDAY6VtSRQiemZdePBUrMNoVjBLvtf47l
U5eDGsrZl0VvQdXchlOV41YZtai0yk4C+aQYoxJ28syC530IAggtdDaubY5w3yJn
ibzH3PuTe+4UxfbSrgk9fbuAL1Lfp1n6wrfjKMHN28CtRYYMJxJkGXfRkHCirf14
mDXyHmMqOIXK6NYHlMijR10kxxULfUuRfSNPTCB7oAmCLb/GLI1F5L2dz0yVNdkP
e0GHE/AQtA6iY4LDfaUJlyVyK8VgipbjfHTrADZiWoTzWkm9uHTnLjFiUiK+9YV7
Vt4BOA1DBVDMI13qZ/qqOThw0Xql5YPPmLgIf1S542HdAAr4NAEF2wuNolMCk7M8
3Loc6IZJN8lJ2OaouvnlQi+eb0C8tXYPmD6iLqS44BhqpDLQg/JKsjlFM9/UA+Lm
3WaS7in0BK2phsRLVOlD4TEFwhjoujrMiw46LgnQz4CY0sBWbxO4KFqwWkI+V7Da
WGFkbpXrl4n/NrJslXbcZtx9cL4EEfmJkgdsX92njggMOq1ClRebQudjxi1y7u+n
QeGtyuKQPeeWwN5zEGHv0Efntsdpwru5MMLkBv3sS7da7XU3o+8iP+5mxIyPs8EK
a/f7MXUiXLA9VF/FB9ezm80kllyr027Fb7TF4t1+qBNdGBlRAV/7R+8U4mBhxme/
mFsa7LSgp3uIo551iKY3fRImp0IjmKHNFO/iTnZa2UYVY2sJikHr+7c+qoSgZvjT
D30M9lkREERM/7gJcOSDaDdzG9Ra1CuHqr0iIgSWeaHnThxXsRJQzRKpu5Sj5f3i
yb0Wkk11MDu3Mbrc570uYppJAtBiuvv88QEp+BKS1nys5JkVH40ttbAoBw91PpP0
gtdbYnAGA5toukWdtVv9IUe7HkPyBH6HVtaxvM9N/67183smeOsP8tFAnzozrh82
oJyOCMEjrz2TCDPruTZtKpYUrG9U81l7mE0uEC6vJg9UNjU5nY4kjAkvIi6stcKI
+24WHJI9wYzTQOr2AJH30ssD610ASS9sLT75fXP0/YWWzJgHo2/CqF/r+gwCZY8b
XGQQ/G0+YoHtRKl/7z5lvAdCsgT5TC3iu9CjPIEqs7LIL9dJH3yAwPIWxdDYpmfM
BnkTTx3GL7LVWllwU2kOZZqLhp1+l2L86/31eOJ7nj+F+j4Nh9sfbauaINC65YSu
My73+bxGjfPZ/Q6xBAPJWrn9hQRCuAnYxB2pPTZ/+mmQ0vup9S8PAJ5L4wBpfqTi
KdXoVYn+lDQR6hy9r5GDeGOvziVTS/7ZFTgGj9iVl+C7Hz8Tmt954gONihl5bAnx
HDabu4Qq12tXmiC+J++fJJj6OkducJtpWTv4cP4xbuI+7nps/d84JB9Qf3uMxzSk
FWUVMU5SPQ0P1e9Zaq33QQJwdXG3Nux/7WqkVTgkr75oI7ueEgDGbMSbODoe2vlk
d/lnXFc8a1f0sG5aUs/JBtUNo1TkEO98CT+bxEB78+5ggooGPIhQ6j9yVC6dZwvu
8K60Wj8eJDvGmB7RiByVrFfBN3dOUKTt+XYZzK4PzY7VvpgqMPFGL8B0hCCRCAkL
n3WtE4YLKdZ9clXvwO3rf5YHZakTPGTT2nZEAmpDkgxmij0Z4xdoWZHniDTVxYjv
8oKjlOdzq3yVuduaoLBptjOCRSWrRggvppFz65thAin9Ctkwvc7gVe/AxhAJjfMl
3zGBiEDx57xzD52KKI1xjQ+Bv9bN0kIZxyU+HVVWqwylh5KeZnZzSCWtb2xWJpKY
wVl1lmZOl95yClaf7j7dZzu63Tr19iG6wBzrfNs+TwzrxfKoqbHbJ8tPWNTwUsSF
Pg+Dq514GyN9fK2qlOECJ21td0Io2KIFvu2GOoDEKLQ4eFdNXzLDmBwFmaIR4h+m
AGurFOH/FeirD4Cqjs+x8SAZtp0mRCYL55AQkR+tkPp5IIbA5Ghq0o3FByjfU1Gb
QnYJPVDp/tMs2raEDh9ENn3He7aOQvO5WA5PugB61oQs/DezdGaxT29CsLg9hGZP
70tOC0J2Ewok1mrLllA6Z0dIQFURV2yEmryjCFHCBYEwo4sz45wbAcdcVHSZ+pQJ
s1TbHCmezMiTh03ncff0TKM4R8tey95nXglx4KuRh3NIDl2/IcltCebhY1iR09M/
SCxnifpETaNnpAySpUy0ZCJ3p/hQYN2bjGDGCanA3Zm8LJkSE9UKWgnETro8W0Ez
Rr1gnC0WSuJl4hRkemrhU3NfEMcL/hLizR0LmR8IiaR1xC4uGDiDv5kwFBq1OSNN
1KUePpgg+sxXLR5w2ArrX49eOBlSJwY4rMw96BY32vHJQHu47k9HF/gkvwocBG/A
81Ll6kiLeTwj7DP95jvLV9kMIo9r0i7n4pyn8wQxOTn+3Y+IGrAYsDzW6ON1cKS6
OccGKC1y2TqsRaHqmgNXkoxTz/VFmTXOl0NCB5UuEWiR8akmtLum1lDlCZsSeq/s
hxZxfewNAGym/M4bgMnJh7qX61CH71zL2yjhUy7xJtzPsCUK13htS5EBn1qMpyO9
UGirbdq75Ty5PK7a+jm4brxwTX2iqoyZh3LcGq32v5nC5zNns1FEgpwILdITyZkM
bT9Q/hp6og78zUVR6qvE8w6DQbnlqbJkneJ71flCwUW/VDv7v7la9I7Ft/iknKpl
k7OuERBVGBvsDQY5fhX98A2nYOgdEXTLZ3+oXpDzfWY48lE6rKdfvWvId6Q4rX/3
J97qDoDTeGYfazEu2YE+gyVa6/pGV02Lqpzzpud+Z8CUndZyl4OHbEAXoN/nEOn7
8I5ajrNDYsHr1W6zqfiveE/Q/I5PfOaUDhtfPF0vVOsd5OYIyimZRPlD3RxxldWC
sIdXQws3WD/+RWtbANplO63m6sNt1Gz/7fnT9kZvXqBs9dGwYtkmk2pSRMqWLOXM
vQREGxRpftFxGqKvS+IniUdh+Im+gyL+AAQOixpXku2jP5ry4lVp1EXvX/wqohvq
/5Wk9RfTC/szCKmU1IG2SFksUhJ0cJQq9Vl39kiOrSftKtQsJbxvTfw4BOumg8hL
jxqZ3ihsFX3ftY8lZcOq197bCqEWY3OSHOW7vK6bU3pB0Is/xAwvtFtUhgt59ALX
UKVmuLH4PDSaBl4UZ+j6Z7tcNnOD310JQYmApMkv3gY1ye1GiwNwCyIoATBIwR0Y
27KQbnoFQRyLg47WCZUN4ncUllurTCiIAgqjwDZPmRMnCs+Ju1OktC4xke3aJrI7
/SSxwszB0bVJhtP6w9ht2c+LEWu7s4vkk2rhqrU7JnR1xUKhSPt8ZfnIGKKaqpQH
Er3SAvnwsZwPWFIeJbkQ8VMQdYc2J6dy6aRWqwyPK73k/Q8RcP5/JMl3zwktx8+R
PrML0p33LN/Ii9GWHUYMqV/dAkRgHCXfCMibWHat4YffaP9ow6Ki7YmFT+1hdxL2
LNRvDNfHBZeG5oq+dpDEsJBbH8U9IP9YxP+jpeco5E40zbNB46md1Bng3EhbkzNM
0vXwZl1bBkbiBeQPfV/GVmL3OZxLPlTvlqByIQRMctl7byjbFjUR/eGd3cj7KvHL
DkQVdjqQ0JYEoCH7inW8/1BD++wtmCLsjya8bC44iyK6nHGmRDvROznKXceAT7MA
yfKnOZgkv3t/nBJ3C+6Ky2hYzeRzfDatm8guWGk6SdhKhzR5Otga/0aKU3ceudMe
L0sdwlClyfvr9/OUuHdcc+dHiWbvstLIcsO+nuX1CJgS6gmkRFpIOoyN1oTcicoE
qFaACzJaVCPAuGWOF//LFPeg05SkSs5evtV1wZG7kgMuP0IOokmobIEZGigK9EeP
/wF9ubhEuoxUCmpNm/dgzIclatZqCtHRq6QvrDRi7R8h+8s2p8/jxMYQuNjXESOC
rk/6eWmKosNfOnhMzjkjkCiRvJicRSIMGjuC6b3N5qiawaPoDtIp9fYkhIpSMGuB
PdWxgQSfjJVrmO3aF7fYEb2gAOxJGNHGT6cCymNz08iJJeUuneduFkjJoInkRCC7
2iUW6KdNpOspVGNHiYaitaaBdvPareTHWLCXmaQRsLrRiRG+iAq+3Wqn0sor5Opu
9S8D10n9EQK7lywKad0P8r8zAGbsZTjjS5b14x8uxKMy700f5m0MeVUq1ClFt0+4
BoxSu0CC1vXqVOoPQB9POBrPIjsV0W6klqe3NISUWcS2bu/TsQgmZ515FmINJEMI
MxxZN+Y6aE6sF2D87fukDQRUGmi62Bx90PX+qXNHq5XiCWSu/+QYAB6cikL017BR
ip4hfKqOyAz58eAKoq1SjY5Cw4WApIkq3Gd2aAfP0jKRy+imXN6SzzqisaEEcIKi
1JrGTNqZYRqSq5Mv9tN6bTbw1UTnYcwAjQ1hEdszVbXxoF6ssYRVFgDPE6p/L44g
nuyXDm+h2hBcSjdwWcnnu+HrHBY2CY9c9XSTG9XMy37M18qqSzLLfDIJvo+htxMh
gYXLgqD1Sox37IlE3ytroWbnaLoWhzhaWRaPkaUV3mBwozyhwJVPPGxCKATpaGgd
5f5fkUku9nagZ0hmW3oikcI4dQhc49I4nBdQz9ZL7KlaAeMP7L72r1QzR8GcjaBY
k+Pl0HriixRYn9uJwDgykdSF0gRBuHjALHXPr+zkOoHr0oL2J35T3DjY7DpgRX5w
zXznCo/kWkb+3OBWtcrHoFlp48juq970HQOZJiLPw9qZBUO6jx0Xqb8NmMHLUUjc
PugZy/R4Dh5uf8OaCgH8+fJoNNAZO1Omw+gLpyKx5tNqU7JBOwaMyBAMaTXwCC/n
NiQ7elxvG044eU6wwvHIUXDg5CwnLM91b8GGgfAlF6+vYUsOjbAG1fuBaC8GkpXj
r8+omblNpJmj8p6Pa5tiSFFVo8uODGsvGJ8wNddSVHOKZTIQNHThS3bhrr7BhZTl
VH8IcTeekj9ZNVJCzjYK60Xf7GhIbmvY8ygKnte2gJ74+fWN67XRovqAHf0rWgm8
tmOY1poHL6RQTvSB3Kz2H1ot9pz9CuoF5dp6URwLtyti49GHFS5AeoJuVqghBk2k
cVz85cmOW2v1tfNK0fIXcd+Opa4Y9VnEcPUK2aY0mDNOdENEXYLIa+ZD1kB6sJHY
ItLs8gWfOTXidYB/PbAJodPpdQD6xuIEnP9MFVCazdYoa3E5mQj1c+5e9+LHN8Ak
Wiu1aFg/lYHQJfHKdLcMS9V0OJ5f3S63Y71R1C5XtTgLv63celNx0BU5SJbkwUwN
rOhmpEQaQHF5QF37zR3zEAW/ege8WKhfQzJw9W+rPKvEP3n3Q40qVoMboSBIGLSv
kvZUI8VEAssQ5k0LPGKOTE5dCOfe/kMrLIT5a2VKUb29LT3jpRfbPH77PqFgTl00
9Z8CN56iBrX+2l5Wq/PNZtw55MQbsRIM7/Fih99TTz0ZoN+28I1ZTrRfz2rm0iUP
JV2SZ73WrLsjm6XIgi2SQhTUgw/6jKAMipKsYWSYb/JJOjVLJlqLLt1sgI2ecZkp
79sAGg8z1xStlMVYToiMEXDKOIBvCV8b/cVY7N4nX6ois/gQ/oFQilHmvljeBXtd
QTBA15NDqns70Qd4Fuek1pFOhftPZxtwCNRaTZsQ2B8+StJNv8xBLZ+2JXFqFXnO
DafshQXia+pl+LXoNK9xSWVtwmVwUykCcN1Cz/GuvPNScg+rsAGoJJQKXONpwn2f
IUE5I4Op5uJcmlwyjM+vRBquFc+9lvnG75Hk0j3CebUP6x+Qtl+u1ZxzXjrGzbcd
X36ccgBVgk5yUaqlMokUE6yfz/e3edm/nOMychBhy/vY9WQO9q2sdGqk2BQIxvU8
hz7Dn9dJ/bWWek4VHGKWJmdOLPjQuflGfwaLYSPiRJbEWpQC+YIiqE9tXtec9/7y
Khz3fU4Fu+shWECzC/Xb8uCPtn0jk5ci5SuF7mgNt17AWtOH0V9JlD/WMyedeBSX
sTbpqGx46z+8psxXWKehgbFhyYzLsRMepRUlNbkgu2zerUX60JuEMSdCWP3Q6ofh
b+MbY6hz4JPhU9oT1NlPe0EMPF6MIp2z45vGeqhzc+P2ggxpdpcblpOPPqA1J0DE
JQLa/jdAsSIqqDs8Q8HI0X5PoWkwQVPGKes1go1Xlypk3wyesm/IY/5TiC6vynPo
YuEw34gbEImCOGyL1iaWo53AqyeAaFlf3KHmrziQ4MS88pqz1o/zon0nPu9myiSJ
/HumIyBQZjV/Sw+8vl4Kfoz6BNLRYU3AeYmsOku7bTUqo8SjsQqKFVHz5fLXvNHL
O0ImDyZXtGfzIlCOd1FSKrBGa2E2vfrAnfB2GMjPkhryjOnp80sEhvhr89yUCDC4
pR7hRYcLiZMQa90VkqTSGdpOM2jctAQgHuHF3ogYs/c+RlMgQJbi946tfAuIoX0S
f8ceDfHs3SBXJCLhKrpdO64YtStGIGiZpBIgRcq4ZooWK9HBk8sBPjZnBnW8oO9v
r7C/t8MoIuQCryJQ3rAmcdk/ZggU1oIdNcFkTu5sSREXldsgHFcAsvKGcDUEfL2b
s5BalSzydNf1181Nz2f9bu2kzU9Xqn/C3X4zQh7n8M8lmI0TnQWyaWUaOWkjbaeP
R1h4XwsS1qnOt3FKrrZe02uGEiBUmTW+71k/ViIzl5RdICXKpAowwO9xHz/l+oKJ
mJknbeTLxorzwg76C9O1AFhahbOSN6I9pntR3e8a9ighQMhKIAACy3sknB7PTr2v
m42XMOJk7aUeuBYk4eOkHB0uuZUKb9k3LfJ8Z4GxPJK21Ka2EkTASjV9841BdB0u
h7rTBrDLX2xlya9uQExhUuaRBLn6OJNZS5kNckeThiSUJU3+SsfP8BJGcJqt524L
Y+T6nt2ZcJR0tvZr12k2MDioDqkzHdf5h6+kPLhpT6AyZCFVc22nnV5BfBXJb08b
MAKXy5pXyabjceI7WLg2Lqhpgi6c+d5c5LYatuDQAp9Q3HlBnWsu1itkxgK8Ofbj
DCBnD2f+nhP+zPyzQ+5JOOWJ+GIwbAIccSLXgXgMbWLpzZnWKOmeUA75ccM5LTH4
yVRdXLLhXaeIXUoIV32tiTLLum1xpRk7tqBpO7+ILuxpgyF7sZU4x+sNdWEmXRXo
OVZfTGOKyj4Pko/DhMhONoL4nEo0E+jQop9gVbpgqCtdN4kZ2QzvlfH1QC0/yBub
FmK0tYiSwfyAZqpgGV5zTDiYJeSytUPKMihpwWEqUDt4TgJpfdAHcm9NCIpd6L/U
wk6ZIuukZ3xZUlNN7IAljpFolk8HVqmggKNdsB6o3/5nHSKsrqxI2xHdddpduUYG
VqGhuflIRJ71IQ7SBEhy0KucczsxM+QpYsrJHghvni06MoNug9Pc6GL3LrWiPF08
iGbynuOF5STohzPErLsjPRHdLJdKo/yiQEmRg6BlLbhJfHMawVF+4rAiwHmvcOyI
JB11mIydyTsSFpnsl9+IBmk0QfJumb0HlIGn784vX/gfssZFqBDZS1jrzdW8E1wZ
ZjM/KRluIswvJCmMUKmhpN3OB7X3NxGXOuM8/rXPM4y36GShOleSEmvE8KHrXdKG
6M4eiF5C9aAAKiQ8VQy/e8dp/T14wgesnhkvdd1InBOKJy1LMqLgi3ujvjSCVzQx
H8ShW9DgBrRwqVlHg1uvF2S6lgxuGGZCtvAQiCPPxwzbGRno1EMCRBKZdKUJTD8P
EFoLgOXsc7fxPSfmqkDl3v23GJOxOjWH2d/QTatboRCRtB1czQm8fu7DMhEqQ8tn
/jnAvtkxRZbiQeKVflsCBWelO02ORx5T0x8Yj5yXG05b1j3CpbhKg8zoL/MG1rqG
0Vc13CafU5skWLs741edcKxWoSDoinQ5YLPL6U38T8+p922YSmG4rSxYQA9vqg1P
f3tLSnVCNVtqr5XlXOmMcndrsAJIZEkdi+XmoSjiZ2WhZOpNg3E70+0DtxZ5FEp5
t29XVVziOtso6DMkmNqLr47RZUhQAwhz/qfKs6UGo29eOMP8/zKO0TXuo0euICgl
n/6Adqd+QP8BPPLlaqQ+MNdjPN3Uox9sGPBAlo7eT1c5feCYmFWYqiGs3QnD/8Q0
5EtD6jrP4cqP/vSsUN6HL3i6xeENKIwLeKOhrUAhEciMKWXbY03XQyVf/RqTUp8V
CfI97vY5iZ1+1goXrvg/2+RRC1rPhUzTBC64F+f/AtudONQFlIv1DrYG8zJk/j16
QHIeGpYCTi0UJ24Tu8+wvSNptNzd+Gm7fFjHS+hG4bEmo/70lFzc18k3d4XT29PG
/uKBcwew9f20dHI2cEb8YEliAu2OHQNcKi79c0B0NCa90iWA/FHrCW1126RBCuKU
UcLYy/ZkTWU5980Uvu/RI3UhlMQmTm5ErMJajWcllnc2XG/9zObjBeVB2CLSnu+H
RxGD9F73IA0YqB+hGLF3Rg7kmdQi3JHC+LvaSY8InyanhQtW1nOc+YW6ExD/T+oT
2BPw3dX5iUx9TemX2P2rwIxYQpYSyCBxjab9z/Xbes5liv25MRRALrz/jAdAObGI
PW4MT54banLr6nn4kQMeeDl5bb328yz6/F+YKko1/92DpMHrXZA3XiHkEBqY7Qu3
+HuIQ3XNH6w+jyPbCjUzvoVDX+MUF0508MHSLb42UraAdgEZwInBbvOPNoujBcGh
PXof98PraUGZ3H0d2JB1cDtLTVMAVPY751aSte4IoDKICWXse5p+CqQdSKZ8DHKj
vPiTPlHR91sCso/QNiecAh6uqjo0EOamAOoLTsoZ4QEUJg3yd/MDXrPpVC/G3j73
ze4XIbVt5J8QGNexE27QoMkt1O4IBf+rn14VFOm0HrmMZ4WhAFyHrX+p+Z+Tgkcr
lf4+rW+j0j7YF+7ime7Aymfyj/BUJqNKtUS0p9RAhm4Fb3ytZVVwtgnBGQm3qX1Q
yrP6pTxRRjCy9/Xmdm68pQEiWS99L6t9qeRUSFWSDs/ibjMBHDwCRTvENdAxnoq+
RVYcqi9D37e1v8hey+q3Vd7VjIMvKGAhDKD43xuRPHkrRaO34kklXmnt/2RqtJu0
FMOdoN4CP7q3NyuY6LiTzSbfvfl9Q4kA3wxfT68Dudhr7mX8LAt0yGfsmh/LquNi
dgBwGwtRpwGfJIlxRbkNWNrmiW35Gs3ME9TemxS7pFPahU5LL3aZVeiG7BN96rkH
TFLXOutZpkW3lpanKef88yshXdrimuUgN070dUJkhfBzzvPoxQn4Hpd9DuCIiwk4
hHFcG+7I/M9nSDLCb45ZOQBUdio2crtx1K/55lh3/SDHP16eaD6oFb2VTOFDOvgb
hckJe64PRWFPh7+eAiQP+oOrjn943RgxpsxRFfBr3liT08zwxdDn0GjqaWgJDreq
r8Yq8hdgOoWXA6jgObFw+qwGqzlAeMHDvtqDMl7wVxPr9F+R3ikr0odKAlhj0lLj
I7DTBvatgUF49VdmgjxwqRbafGGlu/Ov23kTLYuUf+WiI9tqxJ/JmmsWxlcN/Kg9
ba5eSteP/ExTPrhJxqizdudCj6tBitETOi3Ai+vP0Db0ahSW1NrVniARzhzlivQy
3MR04SgXsFzy9QoSDHZGwCK/prz2nTe2QA0aPCRqP29TB9XJBvmovFG/Se1QPZy9
nliprRBi1wGmDL4kod4zDM71yc98Dd8R7MDfgt1Eqoh3VetuzIYIM+he3uPVc9Bv
/WjyfUJ7qasW6YpG1mJ9CGh+kojCU9jhLFfScwl6qkYWbx6v23r+fV92tTj2GsJh
BUKF+AhCsGo6RK7HLZQqNSOkUkm4xgHuRRVNFhkLtw2FtZwL+4gB6Ri8cvxeUZUI
3KIbIV/cYVU6arr9OH6G1JEA9qPXNtIxFdsilC0n/R+jVdbBcfVJVcXxx7gk4tgF
Qybx0dh0Ekfo1lsvsQ0Y1DgBzVYSRtPBJ/2b95k76ZJP0kaAorqeP86hHKiFZkp8
7wC3dkL23DH6EdJGx5u4gjPQJ4m9l2G68SYCDL69aJR0HRa1eU/oz6SBpaTNuqyR
B/vzPCLVDWk7z2ALPah+l4hZ9vEolxM2YLlkbYL6gA0slS+s1nm0uiH2cC6Pxh5F
aNLBaKmVErNLsniYeNLVXo10ptNA7Mz7yRE0HKlQXT9d5bIfRaEcRafgFiiyIrMv
ioe9Bpvbymxmk1gvPVqXvYwcwaGFECP6J+/RdgpAwI3YUWvZJYV2DWx3UzckaHUc
fTEctBUGtXEd5mbWslqFhLgVUmdt7wDCx6h+Y09A82zYxGEHs9mJBRCLJJX6dHO8
2McwTa7KjELFcRVfVDnxs4g+1b5MGJ7BMNcnblBIHTvFjMejnBO2OWHGUqIp786e
lcDlJA0fQO82Wo20Cf2toLLQCUBFOhqGhkxR4qTZCyKOUvjzqsRcQLnz77T04MWQ
pqg6IJHpPsWGiN//uNl4zIoOv53k4+FLMgnF4IAXHrqWtse9+GKKAoZVK4wQKfGr
QjlETZe1VIuAsv4S/MtEbPgOxvEbuURp4o0hTT2vTSKDRJi6tvSgoWTX7J5bRxYz
/vjrb536bF+f1/dSvltBYV3+E+asN6D6t9VSCmu4BY7nPc8Cj5BGEyqRQeSB79Q8
EIbtNL+SfaU/ef4oRonbMJSKO7a3nBZhH1Jqgd1ilevY7CVejvLPJMhKk9NadU6z
LCwD8iDGFvSX8VkBp5OjcR2IpRmwyAk0urYuT6HzfSsvJbXO7fpLfusgWdjw2RRB
RqXrMUaRA/VnRQmmX3zE27NkUI7fafD9Twcc/Hwtm8lGhP40VGm0SL3CpM05wO6R
QmHDEF6Ol5k+NhLZnzKMEPX3ilbIZOSWNECyK+v5d3Q89Gibf4qS/oKhBI191x6S
KtzXn1vgkmhBsWZZoLTM/cWoL++x3qsusq8JAJk0KB+8iimfv7KHW30w4Y78txCR
/Vkhf1NAbN6ocFjHUBeVFkpiKmZ9XAt1yH97RqoutumBX2I7vHkyBbrBkXWUtJ2D
d3hlHHFjoGjuSDj3SrZ6HQkds9Nptue56Pfr+UacMMNNSGt1MRa7lQiJWWlF9uRi
Zp6sZzhBd+IimGT0yIoSBRSdJZ7NuuSc3UeeeV0Irkju/qRR7wcyNwc+FpsTKSwD
JlLL1d4vjuEAUiCQX+qwr1jB8ns7nknl9GlbiASlnFZk78bH/Nyd1AY4FgA2GrQb
Pdrnk1JStOkI7Kkh9U9UWtAReKcvhmzJWprHmGecK5SBpSx2NalnKXRrS1OyRYX8
lPhcxQTdsPG0mDoGpsw1+zXvPhYjq7/RHqOnNIIQpxAFtgNNLd7TuFQ5og3Q1PMM
mVMwW4bWryq2vxGkRFfPpHhZ44bvVdYKKwoZVVdgZCa0B6B6dq5LPQmd9fMaeGNC
M/8s59EUa1vsH0jRR71cSVb57oI6lE9r+/Jh+sMwoZhO2vCnlUdRVV9pjhS+JZkC
cls+fXd/rLwyEUX9O4Z5FiMuA/tHuujt2Y8pGpBKHSNzuptKI37sFtNe5CT7ltG7
DUIJoHyZenO6AETHLP3Krsxr5/IREfWtlbgmcAczdMVMnSJleFcKA2gyP3dd0zqt
UA+eip2oix3w7tHE9easEhvRmo2FIflyTvFAb02VnfZBw3baXmD6vbcgs72ntF9T
p1HvJcwbLm008C/a48hBcxQap1xRMvUC0piT6kwzN5dW+tVXYPU3CrNn7wcxZ8+j
HhxaMhMlkW90GGDp5HJnXcRakolmKngzl553WOv+W5RF5EbZu+a79ST7TIriZgC4
RyUL5muTh7GR0kZTeW7NZsjdCpwMSIUUgcC49bZzWb3gy1vGhy031kp4dltFtYJm
wmltVcfh2usV9w+IvEI2KCevuRPjIsIyNwETWapMmDCjbc3xI82SFyR6JaNAqVLr
oH1VSvtIqce7g2kiZsoki+CKMtEpeZ2ymFvsKua09L8eAzsaAo8U89wENelCLUKS
AU4jZR9QwcB0VBcoJztfD6zr5s/b0/rb5VF1cmjJ9ZaDb61ERC8OcAyrrJNCHz2d
Do4Gf47jdkPt9Qy2IIGounODO+2W49Te1DNopwN/zN9YmhLqlpknNh7y9tQ4hcx7
Gxvdsunm80DuYzl/Akqj9VQqPEjKPbu03cCnJki+r4r+deGWmnGF5pFO8nLgS/V1
1NxWVTc50ObIsX+Q2svNdak9IbG3c3WHfhaAf8P27o1Tjh8QAHqYkIRKvcmCL4MF
H6Uwe3DIQYA8HvnjzVyw4x9vVjnp85PpEJDksroUz9ChCxdQ4kJCd/UUR/1j7iRS
H7ph4ONTcK4IUPdhcn+4LVFKYeF15rT3jyfmqQpCxEedKdWQFqZXkzFA8obtbdjJ
RMFIJoB48T+6fsbfKRGhiPRJlwv1hYax6sNlx9auszb5190v9W5aO5BakjPRB2Kr
L5IIJpttGTcYnCUbDaJPJU4q2p92gYj+zozAjEBfBxDNz/MPN9uxop03VO6vT6n6
74xw/3Dy4CDANXgvJzXoATBYBlVxmeq4EKwqAdDZ2cFG0JVpuVC5tXS4lEXBrPG1
w4azws63yS/BfyZAzHWTiUnlKqjAoqya6euR+iKHPWiYgpKli44+PptqC/DPgDT5
2yFsW5Oo+ZUxiCjURC3gyZPwnLqjObHoTFcR9C8/AEUsub2Vc2KtzWzJknn5fNYv
+MyK0Xws53m4gic+Elnp92C/nTJgJjW0dIE9d3/jIY3PAcSbrKzQ8WGtckegbwsd
sozjcGhTpDEXBpPMhaybj1JMXNocxC5VSgeQKSazXBztcNCEKeXcP/n8/FjF6u5M
KdC7eRh4ApE8mL44zbWnOaIwPmcWyiDzRICI1ChjkOd4L5+3eTFuThQGEeJR5zXb
aWx/keg7zMTmy6GnL07Yn6Eu1A3k1fXEmq0lZCUB6/8JO8kx83wagtKHmLNa2hoc
DLMQCTpTj4eh80NcrJCLCucBVFQc37VLUr7V67YM3TJI4/NgWnln3i33heiMtvHN
PORzI3G+eL4vg9uF8+q6ExhRW2vYjqDYROp2v5hhDn+L75ksQBPg7skLd8COAmKw
2xda5Oxvdo9+sGJu7h70mT8e2xUOY/M04TtEls22zq2lsbRkHzsyOet6bLhYndBY
BP06sk6ViaMumF8iDQdEYPXvZ/EBT0A4v/+xSds67fAZf39kNZNTuO8e0XuIzhSv
EKpgVT8TbWRpWSN3B2ZwwgyyAOs5bOn/KuNSyofs90RTqKkRAt/3pZpwTKH8LeUB
ppAdOQm61GvhFnpLr9xxcNcyHL5W0EnzCuff2IrisnjAzl7xj03BLZLtTKMjDXSC
uYheMmmEBUZSat3OhL+xbHAvO5E4jbILRmfE2N5BLrf3hD69wzV3XKsG9DihXVet
SfychhpIkhoQw2EeV7YjXkhU/mBg1Ku5jFwvhDYSnHA2zZSYlGo/+ta6K4PuCx3E
aNisEK2TLZImpb2LXPYgChMQQko+5AAFiwXpIru9JFIguaxkGMW9vYTklZSMqT7r
Hb3+Lr1cWAwsVNBusKFmWyXLBaxhSbokAwSDx/5jEMR+i4OjkukBXysPGX6Je2oI
Woi9MeGmOsq6J09YR+TaN3da4zoef2kG9oJhZ/xnUZHGDp46X6w6d5HTm6BvBkcb
l6gTInMR3k3ljUi++5SxDS6HMw/yLtuV5HVo7BMsTdiIrZVI+1GfJawgkJhcs0IL
GXoyt+rfdADEfDoHmH61aIVwVFqeMtIMM6MXh9bdUxnJip0CVsDZjnsD74g7voRp
8htoBdyABBB5rM+zQW+Ip6yi4QStAHHdTEoqCVl7aaky6sVZhG35MriOderMqy1N
FotyQ1ZmNGFTia/pKejdlqhbYEO71bYhKQBGWPR7wBbm8h6tI382nxC23BB1hsQm
wRvVs0S4btNQwvMpkQqW12TcGdAHp4442Z8aO4raP8/VhbwWSbHOfqoDkXWzCvfi
jOJJfLbqsndyC6pALz/sey2I2Xm1VaunH14+wnHsXc/U/HTnxikbNXrF5dU1s3eS
Tl8nRnV5nbHcs5v8B4ynP8vBwAkbfmeq+cGA+YAoRzFCHIoWqVH040U4CDH23mPr
JA1dyCJdq/fYiThSYWUl7F85v1JalqwXk5rZCHt06IF4KpobH5eCGkJtc/v6w33p
3QoZvEqYM0oxdalxFMpWid7zlpUQuih01bX4NVgYyuWkuY/xSit1tHbychN4iAF6
+Tzv21hi25rB0NQIn+IMmHS1NMeKv+B63PDrdnlNBgPNMIehfOnPvPQNQpuhgck6
37HJIM47BfCFYwEU5emCICuu85R7gSkJYU/mKRwZGszoT9isB23hl2VvLORDsL6d
NPriTO/G7luSdTHErazrxN3C2dSfKypdqmW9Yunu3z2GxzTHqiWYx1pFEVZHzm69
KkVcSTz47GeirJfr6QbyRtqPx9PKlBD6Ies05XQszg7WMtixS6cs7l3tk8x2GpnE
XwMtZiBh7CX2AwrphAwjckOWwVzWhuXvvgLDaoEsLog0i1/OAJpdC9hxtOnpMgrj
+mWqlu+S4+rFb9I9hTvP7IvusNjjwEkf6sHB+rI+we8AhiiHTFD6dJ2RoYg2OdRo
sV2CtsOwWYvx5dRCnnD6nOap6vEYe4Y879s+nEv/YIalz+z63Bx5fFUZ89medsKn
qoSvfws0mN6MQrwMr6aFcfzwYD3xnb2P1Bl1rs8faeUgSZepKGrn7MbC5GAAbEjW
ZKi5poUeqz0giPMsHzdlnuDDtJQacg+aAT217r6c5U/C2BC08uYO7e8Yup0jENmy
MGdfi5TY4KhTO0TBcFinwbvZc4cx7xNQjAfZtasfeEp6IHmyadWmb5uzxMzyf4ED
NdpD3RMgBpv1F4rz3zxWADCzmlyrAsUBbx2lLVxwPts5Kru9ptmzQyCZ7BWKzRbc
6Rv5OEDylpawTtlIJCQKieIST37lTfVSKdvblUxn6CKuTcgO81Wa2sL+IOMUp646
6pQwmwd5DtoMQdfrC7PLkJePU/1R2XTxVTQAprEspmRw3XsJYx0mgCffgrBP67ba
ydNvE97Czufz4wbCRfa/fcR1WDV7E6waoJu0+SPeobESEDHUfhqsOk8XbX24pZ+r
l169xF60O688ytdBN9BsxbltvR6vduw2L0qrJ8EAq02LQx7a747nvp47BeT/30em
OBNtjB2l0toQtonCvRnm8zpgkWUw5H68yMbYigzA9APqDXcm4tusahRGB/lEKqIQ
qOxD6X745kASr7zaw2sFA7jWW83kV/vJuMaq3gXQiSO61V5Vtg/1VlKeikHvuDFo
7PUQyHWgrCC6uDKWJg1ffrCr4jZA3dLlH6K5YOhRy4W4sA7x3j6Rmvkkcj+16vir
8J1TQf9uzepA0tC4z8th1o/zH/MlV957JiVkA+eAYKssZv97pD5rJtJi90qKdFuW
mQ67K7fR1+JHjcNX2o5bWxNLufwx5nnqkBAqlA7l8DSupCrdBBga6f8v/twzR4Hq
5yXGt61n7NQ1M9SVA7+gIo4AkoW++LlFLU5pZ1cwJcgPI/ciesGt+rFem/d0PbbZ
uGTePVcnqIDdXAeJREwd58x2RmJWWnkVoE6o9p2kseKwT5Cpd+NBzDIK93Vj7MkF
KoU3JJkrsJ7Qg1iq8khM6u5ZQw+TGqcukljMCq/CwAJyCp7KytjsxNt1sN7/2/k/
E32FC8s0R34EqDrLuGduBUviqTBwgsRU3i5FS2DvFg6pqgIlGXl+0LtaxohsukG4
dQZxdXm8lPKfuLZBrG8YX7Z3r4WkhLjUYQSqLfZihWN6aU8AiWaxvRu71C9O30/1
fckdR8bPpEMXw5Q6bCTwNKa9bfawdrqpzU20uXiphW6HE2xpk2RyXZj9pZSXrSN4
5CKTwsyT7aIdEoRJ8JTLCj8Sm0bITjbqaxQCr/7TVgcWJinikKn5qtiSeCsziYI5
1ONkDWjW7X8VJsEjJ16ot0Y/tkXex+GKHZGVYzdjE9alcuzsct0Ezb1NRm3NB0oD
LPGKP2TCSV0S40Jg1F8oTmNlZs6tpYiTIlkDDl3y0MeIogWFsTiUJkBIK5tltr14
J9ud7GP+YNkP0BYhT+J8CyJ2PiUDUxDOVSIFEFjP95K/6Sa8TQxxTqDq7ansq0eO
sk8imBtZ3Nfw8lLAXOmSn1PmxbggjZRKSeBZP7C2wTwzvyO3nRrISfJrGRVpwDg0
/sMWXVLADF39umWMN1vjBo6YlqD2w0i9Tfp2fYDIG/XneYERWsvq9Kpaunuo3m6C
H+ptf+2xjcW9JxQN4Sg1T/5/saTCMLBsUxKIuDXnRP6XI/69dk0elg3oAeM3DDcg
hko8iSKCWcYxCKNmaJtgIkHawRC0lo3ZToP7oLkNH/XspU7DBlH8hq62LgqKqm3D
l3QAKB17YmXWSPtlM8wAFAFFi2KBR1imhppyJCaWWEtty45cpyJIbAmIyKJSO+K6
OKK8Mx9Pp/oshRZ72dFTHhv2XPNBPIFXwGAD2TUsJdZ5SLlTrm5GazAUj9QbpGdN
wW8x8X59LjLMXnWf6cBpCYarPmOTt3Rml3t+mdGpxCGmKHkRr3MLavtS7pmili7J
vjuCSmJC9K8NDXOHpj1ICl3MM9hi3L65NdFSkx5Xe1NGbGlPMGki2DkZMo3lseGM
WqDfrhwnvQC0d0zAuAv6M0DTQ2u0Byc6fP9/cVhtmamXP6uArYxaamnYUBhvjTCy
lVmTZ2CBOVwhpVJjfou5S3L9Sir+mNgvDe0JfTD4GuMntVqdcLikrKi7e4TVfFH7
z7CL/tBYbjTbcun2wN2J7KkNxKCDYuelaa51kHlilYCQ/fc6JKm0nSJWm5a2XtPE
2xGoAk1/IihZLiVH6dWhgngl05z+pqyyqrOWP4f3cpen2NMkpP/lKsyBVK7ik0Ty
TgO5z+Ly/ZdnEi91mBuURdJdyHkWeUmF8kEEPBZrHji1Vw6u2f8g1SxV/Pg+DMYq
2W5ZYsOo2dYW6+3YfTeY/COt2QE2MLxvjrVikEZ3JykbsrIzI6YlZXi3IlkBck+S
O1TCYaqfEFn8m91UAjwhcN0O1u0/zbJRDl0KPqVwr9WjR4bEHJU/T5/PAzgs0cVx
bq2rZMDXdONL/emsUiehzanxTojlyfe0YgJYfcNo8MQIgrWEDTy4r0w6c4glcdI9
BWak/AHmNl6HmtMpFci10J5iKyrzrFpw3e9GHv3mfIW9re/bnBYkkgsOWPh+k7C8
owbhA/q1O/RvPFVKQYxP4/LmSPuX/rv3UK75o29ovLYmtIhC7kLYCuOntV23D/Dn
1TNbBuJgxKhuvGjfgank3WCBvF/V5+ru2qipvRVb5jaUrqDtj5yT5qauFd2j5EJB
GUzUJPxOxG4xfabAJWI0ZN0k/A2oR6GTx3hBBeVqZsuj/zlsBNA832FPjA/rPx7B
rIyp55Ay7sd0PeMYEjoTspO6lvZdWY/meaHOdDk6eH8i6DPyk6xvY7JndFIF+RlE
c03hXGDod6GfwIlXPNpqRtEgjV6y1niBVIjIt95KHr4Vt7TrBY8vKoFNFbXu17Ir
feh3IyHTDSw3rGUU9/xwIbnP1aWhQnzwJ7+mCqeyHaMIu2hL2swCT7pC9xe/XesD
w43Llb+MFH0nywraFHhSMsZtvq6iC9rDWuo5p6QIVLXp1HcjDDpHzLuILTxNOe8l
x6hzm/pyJ03eVmvG6OvUDt736HL0qyb8vJNRu75woPI4XnThVytUDa0h33Tz/UcS
/6VNewYqdNzXYE3rjLBygyHZDQXH9XcIqLisLVjMYQikwt6fkEOvPGPsk++47wFv
ac5S5Giu2Og5E2Q/a2ZAsfZmcB0IbrZrKRB3BA0XzM0IWYZvuYWrKZsDAvB+O1/u
1xyHZo72/zmT/FKOdfS4bhklcSct+4sbFAWOKTfXXugqHYczYQJhJDb633CisMQl
YDZRITRAz5Y6/Cft5eDE0jDjRuDGd4/4+HKRPTpmJ5p/anrk1pkBmragJ1b0YlEz
gmVm3n2x/2gWm3Ik233S7GYsMvEpJhYhc6gI3dkpweTfYXgg0a7MYlRm7qPN9M0t
whfrjZJ56T8RAjo93WNLMr5D2RcoYHq762D4w06ISjA4xbPyPP4/4bpgQkd4aIr+
slLEkeSxsdRFrPncugsagRzzBLMKx4zQTQyPu+2fHOqQFbRnzD4aimy9/i8Ey+5B
+PPndc3z+iQs2BOaPWKBe49IN+lBD0YV47CLAG5KU6UJaBKEMJa9S2z3EfrJHdi3
XXG3ZUZRKU3GGaHHA0EcipoRsDBrwXgA4ZzpkNsZG51CrF9DUYAuvUMIRmAR4sCC
8dmzwl+9NtnFfKNcr3MMR4LARiX5itoJjTdRFBUKRYp61JhS5sfPdOkbSgQWSXHF
QGDo6VEYU5o9Wt84xuRev2Vrh5WdNe2skhDuerDaUJ8+pkUA6TPC2WRIX3uL3fDD
caeHhEMl8F3fV6k0rMjNnF+toa+DcVNTTe2HQbp9lh/xwh7pwy/5ZqxX+Nch9UXD
r1r+/3huRJgLlgOG3L1vrtn8lZ5g/cZYhR9gAkqcTttMXzUgv5qX041sUDvQQAoe
KqdLPW44D4ueaf/4z92yRHGKReoryyBreRFYk+Szb1jsj7VzA9+Usvi0/AI9RQFQ
fH7kIJu91dvTEND0dKz/6yRTlxAuimtbuiryRon2HVFEEMXuT21bH5nOo14PvR9d
OBBpdbqatq2dHCvxebak3GS92XUK/X5D9uwMYNm9DwJaCd2yLjF5KXAbZAAAmWwX
9z6YG7ZiPvcelHOnFe3OiR+ld1ffS5XXe81xWJ8n5BTrXLYM6LuRXxvon6H1UZIr
9gAwwaGx+si0XwuL9XZybJyWiE6iQcWqpc29EtE4GlJrVu3dFG2pPOhg52anD35+
R+a8armxq/YVYTatigMciHRf3Ew1PZv1cWj95pfvFfX3JDBA+Sb1qW1Ia2BsSVuP
JBR72tccXeIo5wOwfn7pU2AdywL4k1C/cRbL3GOTQx0YdkbJUaVsPpwciFsxGRYp
iQtrYt18hkhmRSEITISw3s7tUmFpAy/2mwNVRQ5noFaxxdn5mN8Sn3+B7pHJm+HJ
A/m82ZnjtMJxr3MQBN1Yt0/BdSjpI7dbRKOtNgQRKrgYfotnFi9kTgZxsO5iiENs
jHboHim00BZFHu//ctls73VLhwFQvvWzowi2ITVyzWwehOYSdlg2e0EK2yNsUOOQ
CUneUbm/ZrRGGQoD9mrbHPWXvcraYzw2m0SsNODk0ZG1MhNOmubzNfCtzlxbo//A
9mv36RED4A2Vh+c+9W3e1nj/6kbjOSv8Zg6UvIOtrpMthGS3xgLRCDEgLGl5Q7Zr
9vXBH563FUgdSAbhxmK0YQhPTqkNtWQ6YtsAw7Ac0Bq7yCUn25gYMdatcvRSUN6x
rFHs7yafprLbXapKUPxUuviagR+xUnzLya0MG6r0jtK+Rh7rGFfx2QbZSwxaQvwP
LY78vi0aguGYZuKEL9hxUfzKV3OzSmS7ATTmb+v0XA2oeRH3Bq8ojGshwp+Ze/RZ
UfrF7co6ZEnHpq5pM5o+z7ixAQ0LNd7VnXNGHSNMvWvtKyXLo5Jgx/IMDl0OXc+S
dbeGXiT+9suGip+CR3PDADppHa35i8HiyRvKKneEBxjh/ByUuq5zw3OVnm7DQuxO
EuWF7tmkjJ44oTpOlAmvGUJEtkM8Li0Mlid44Yyf94L/leUD07g58VpTOZmz4HGk
idmvs4jfrg8r20swtlQ969RJz+tYgNAk6/jeqNU5fBZAXdLfMBZZA4pi62CXMTxE
XUUQTg0cwzo5KVeZo5IM3PnlckQ6kjiFGuZk8RT6ViaFRbwvSdrQmY5QEpqqOY3n
2Ul0KTPv3msBm59DW3DZfoxIq5lKuZGZ1Ih2k1R+SWmdvyFR7bG1Cfido1wKWV/s
BfNDCn6hVGwXAFZDkZXk8pdHksVfGeZtphAj5ntaHMm1Jq+yzg0otlAkLFF0ye4r
MkntXUJjMMRY+PXdflHVBTjUkTRiComexUxMdoYpaeOr81+syPsp9TEknoDr4PcQ
mEqFDpbrYr/KR4Kr6XLjfEI0SY9SRrBVbBqe4aqrYp7kOa8Iqq1pSWuKxeEl9lRC
v/f/xDe+p05BXhHrgQr9gsxd9pWSCx8O8P9MnjJ5Nzad7uogNCNHe8gLU1M5lYYP
JK+xqYCIsCHZtcfvuWACJIrCEgxKljQGLsvs7Cg4jrNfhF67nAH7+bPDqDf70Gw6
3UT+KGuZOcLFuRAKQ9SFd75uuUFYhRdIWhOpAeAMeme58WEVeRhxjf/434rVFJEH
vb6a4+QxubyRXViqUsyudl/5bql3infYZDO+a/3p59O7QWmXGQg3k+97oOqTIXD3
mZI4P1ekoR430dLu4DlqnTaNZBHwE37YQSpvnvBXhLWm8Ukbvyu4Q1Pu5DyNFNFD
4cK5kiBNSFF5Vs8zhWTwzalwximgLkFTsnONxCQI/wvjWBaYf6O//kbKDOpW1KbS
RZw1EBEkYIEtMoprsalcrn2Y/cJRNkZJQY3QuAg3ZT51yfV5W7l60Nn7Rp2CQrmw
b+5ajOtLV5meX9qR3BVirwWl5aLk49V3E31ALtHSsxWO0TLMmb3Gg1KQyvqw9mGG
7KhTqe5Hq/eWaLBpNJZOlZbzjJWWegAGNiUZiSEbgNIjEnf8/2tk5d0D319Hxktk
/2R/jJBi/vWqwd5Bafb81qsuhnKpFaZU8biRKJX4/WLOX/MRuI5J4moylF+e7Hym
MLLcCDbbQD7MZkUun0HMJnpwpauPoaeNvqcu0wjUBX6ZB9SOfg9ja5IXuYFZuyKr
sMguKNfA7IiIMFm0uHBzOFTafkajzCCtXFlEQaxwUx8IwrXKIZnJQg6q+W9Rnvlg
CErNomHJYqUiOXr5qFAhOBFs2+nA/vJ1AiNdss8rRnSa56o/FrL9J+99WpZypjIX
JJWFyH6FInz6nIVnZOQt7SUTULQE0BlJGX6dmr3/AeAbO9Sj08Ty2FfGDXVJRMua
a4jwSCpq5AQs/vMBCBTrFmvNq7pq0M9ir5d2Gd72+6Zzf5AjbwxUIyV/RbVtZJgu
5DLuEkz/Ec6yXXzY6PegcWoLt9Z96DVEkvKmfWX0cjpmd52dpAjiFB9xosYfjnCi
jblQbKpFIwjftzo40uqm8ywMtOBW78/T9H/1Lq4OChuXlOOoFDSi7dag1z7MdWEH
sTGOLU9RMDLXsNFUoU4ZNDE6UGG4jYTnYKntdG08HgDNiOx+ROQnJVC+67oJjV9e
fyzrlDX42GUSpVad/3sMNOXNVKBcI+KEMYFHKKElTi6hCU0tDit+/N7q3aoa9zes
eF71WEg+xvbB6iGfanJNz5ewqQMTMg1HnlROatirTCOSSPNQEoHhEYmF5Wsml+mL
2rztNt/aVs68J8VDTGx6mxKTMCG6hiePtR6OQpchi8tp3qcxI8oC1Kz51dEu99n7
wrNtrU0DMCppXhEDLaduUKLJ5vY5tH+P7a6qS6PfJDwj6qr2v0rDK9tH35XZL+98
/Uxa/vJBPrr95GDt1Bwx/2zHMEPzUhK5xxPW8mEbolmp3iUv7m1360v/g9lz5d3P
eenSJ3zBG8ec5dXmEJ7HJYz5hjnlwbVdbyWxFtjglGGugxtnUKO7uar5EUIdbo8e
cL2tdCAz2PEduYqIey7l/543wfm5SjaPlyY7Ycaweei3ooY5f3VhZMDlWv6jAbeL
qtI9Vm0hP/ts7xRK4ni14dxId4/NoDc8PIIUuf6w02DpxrNWbm5zHN+J6fLeSCtD
qb6I+iOoptr3JRaE0qarkFDT3P8Y+zsMQ05JVj+MLM9DOzzTQZ/BG83P7LjAKaaq
TroEGkqSmpbThVtUbKLl6nmIPSkBBX1RBTMaBBHFoSovxuO5PWhmYCyS8qtUpE/l
ejtuDWbVYEKLtShpt3Vq94Gk4JjkROFU2G3s3c5/KE6dGUgKCvvlY9U/BlWtXOO+
L55EpDti1WhGdxHE53jWrOMMNdxjW2B5qO6uQx8zT2zZlhRtF+HN5+lFONgZ18oV
3exu2eASOkFsfOXHXcyyIw3HILG8TBeKQ4t2erEh1e7HRCBN+32xijjFDCMAIbH5
+VldgMMOOzOAYlaCecYO0FRjPLDH66my/AY4KsZsP+fWqEdjaMDOkyBpFb1P5JXP
qJ1vQw7c32pL/FzWcnfeyav2t2zWWRH2CLBQdRlzg7xCKyrDgMKWVgGOnglh+2sf
Pvqtl/UHh5gczHYRSMhgE7Jw7/VoHXTBbDrJUKYWBY0UnmwT6trJXWFniApTpC14
q3pnymZNTH0HavbkcZPxma6RRDZsTiLuObjTdVcqNxhwybUV1nAIy0tUi5ZwX8TR
tYSUoXI1GtTq/qtCopH0qyFj9j0q3Tb429u9BJhn0x0r9anjLz/n5Qq6ncRpwXLp
PrmeAXf/EXdwJa8P7KgUjMQn+u2GrrXFOwxDpWfaSAeMyqgqK09D8P3rc7atExp1
qG5XoqeEXVjKvIX5D28RPEmev1PnYYaziW52gaQq6PrQA4me8M6o7KeTkHoWipYa
8d/WivpNFrc64aY24IY/Sx2mS6n6IrC9uEyCmZ+PLErSu5upS+ACZWrsJKzO7c+Z
W8gUINIAaimZDSEkMuXo+gelg7nlTCJ/tUKyu+LNrVvs7Fy6MSu2Xrc4Dy1qI1HA
YBc1Ek1iGIX4XhKFIE8NfIVPpZIRgmU+yqYA9lcFgBgCB73kO1THJk/85ofOpPia
+aO4t7A34yRD6cyPBf0SEBesYMbzkdN0b5ZK7Ayapu1Bt5ljawDLxuOiW0WmQtTv
xI5iVgI7kRIfubF3eb3Wv5O9Zkt9VqQqUA/VvzjAslOePy4k+CMefpYq3sYB1E8/
oNoanHfb8bB0D7CQ5HWLdvFaIX+2E1v94oVsgRAUxumZQdrLM80MxcZYqUKd6b20
qQn29qwvnhrMNqJ5Aakyhe5No9IU+x1qJOlA8BWpLJ3poxzU/ty+7LgNhh1sEWwV
NtySYPQe+xLrMHJnMAKok3uy2/unUsSvwELX2ZrO5SNRlToFjywkzwQbHXHqJSU1
kS68QpBQZmGEK9tDGGkpgqWZOzGs2ZDjzX+Dqz4ZLyJwSPuLFxHJPDstB47JtC9F
bI6fJERun33C2XMA68J9xdt7Qwj4PAJh+18sQg0NHiKNlzMZJgFeMsJLwU5Ah32e
91SykYzjki7Br2UQ7GL5QpLjgVzhGkQPOVwkM/N1JRZaYXdTyQ66+f1ywC/w3znJ
J5/xU/0X1G9TILQsmgNR9Lz6U30oxQoDrqIz8m3ssoDHaIno9YIwa3PLd0hxyUY0
r4rhEEtN1sK1SVHdSiG4SID4zQkH9VoYlOfe5ZYHw+xGxh1g5Ite6pAuWgO+ugZT
LxRlnrNEqXh2Dyz0bfqvC64jIw/Vj52XWHk2BiHRuGFHoE4ZQ/uN33V2qVEg4NJg
X7Tp2kR4VNmmKW+2YAXW2jkR5dQga7ayo64Zx7Oib3MhbpcMfQWSSwmYS3uw1f3N
Yf760NbA1UCkFMBdz39jAURR4jARQtv11Sta2GszcqFYmSjbFTUzCGupiDFqg6oI
1nT94TKVWGtsXNbLI44ReUy/llMzgqJTJfRdDh5qgN2T4T1Kxq+jVQO35CFHxKaX
usCEaQd+CYztodmU7MnN4vxpjTeiEeD5aNdp3w8NYEGbZ6whCQ67pMo0DnYak5+n
h9ClQ4j8fTswWn6iqcbXkx1y0/mfK3b48/wEXy9jKvFpdHPVxLPockTsNssXGKZZ
vO1SsdFkDTOaRhWSs5h/ebU43Df21a+7FaQCJ8KRTlEo5LLcrpNskijH7TYoPSul
DseEiAcbV+FOMr4477rpaQ+FoT+W2yz8iFHVl9Tuf0GQrzjkvi5jmupKwQv+lnW4
hLlq7E/CU4V/t5dgoPmohFn/4llFL17kOdPoWkvaxxSyFsHosA85WP67BrSWaFmi
mnSUVp/5Jx7Iv8xRXjoQQa7yfzI04fDhe1IIAGIFXz0XMqYQWPfnjSXHVmlWJ3u5
wsdbLftnp6+ra4Xs/YocePL42cFAjp0S6Q51f0LVS3t7xLM6TfkU1LlS7T+rphWh
t/jxlFIxY90Ys6VvhJA/K+tl+g7KYqOpklRKLQarq6Fdb1nAjz4fUZwFk6fErsDF
EfJ1gEnoB6OvOgy8YCOMUbxWYLiJi743ms0XYQV4HM1KTFprebH+1EGNkWOe9qZx
Ppd5Fjx2sE7WfODf9ImfGyULHZs1cKDnS8jHL7lP+zsZ3itsNOhMHKZjlR9EEByY
bgME/T29fh2oBNaiqhQVW9zgdVFQFRqIDnomj4GNmAUPSrsdF/I4MUSaNYLxit8c
TtqQeUlJzDbYS3VKKyxusUniMvJ1/GGGMXgmahaOiPhYFfXRY55UJiTidcW0z35d
kip3f5dQ5sBeAZitvKOL3KgI2PiAu3Ii36Ohzxtu37TJ+BBi9TS3CowSqf5bjjjk
6TP41SYqAFRsDuvXmJNaD3jM3es5nV6qCAZ8mhiDGffgufcBM0Nt451BMHZ1spGo
iDg0OCuHmUcZysavmz3tihrdEqjix6iaYLZgIr37zpWeE1mK7/VFP5p3rMdSv+0Y
ohT63XPV6sKOwvfpYNjWg9FWkzWkfzPq/UscJJM8WxXULXx6WO5Tma0HcBKs3LgV
mH9GSA7FlQR8gZxKNAxZhWWFUfybYnVO1BTTJgU6HnMgL63TJyEL97nB+9DsR64F
LcrM6tm7dSkTL+ShsycNd1VQ4gGuNwYID5ctPfd8qtWlUwOgrBv9zho2ZI4iVH4R
wl5MXen13XPVH1Jt46r4HGnHt7URsmu37k2MFIdG9/e8XwfMH0svjazSr02aRD43
zScYh+arKnfBDhlOqoafQ912McvSPI0J3f3t7ifrBWptXPYLiVnQka4gnB4FU9vK
9PgUkNF3ccw6DqxeAqC3lSAB7yMJljgDZ35ynknuQ6fVfFOe4fvj8CDXRA4nRt54
cBLaMAu8pB/Rv5kXSdTiIw1vDgSbsZ9DEFMyz8UnQHULKD7vqhFzj3qXWsUQA0hi
pfh8vhIm/lM4mqDdtEXq4Tm+4+ndEButZbLjOdTF2nf7Ct0ifAeEQJOK96E6tqN0
Q9CNvfDh/oC4suy/GdHTKZfrRq5jskHE5AymURN0wvYQlCPnNMhqc0T+nSW3Nyfh
ZNIylcD1W2OOVoqtXHIk7QM8Ox7FNpNMZYwX9cPBjwHY4IAhM5XgYQhYFB1SOmOl
O8nJPtt7UnMsv9L49h3lES0Bv8/4kFOGMUrR2KrQQ2aqw81i5WEKSy9khXv1Giml
uKISG8h09ZP6/VnpDKddcZ4qssSbF65sw8Efu3ra24ZyX00FhY4hEHo2fqJjSR3D
rgmgxhnN7P2bNClgGlH3oRMTmmXGiw42M6PCKJ3FCTZuxm44ZepBhvfFg+hXTpqb
kCL2Lyn9h2U2POSxPdxqxNJFZTNfWgG7pbcZl1gsB+5lI+YaNeLxsuVOjWz5QCPP
6730aIl3MWJG0jHAx3jvGvN9+oC5KcPcIbxYUqD7M+oMBImHlkIj+C36U/fBZuy+
Gj776D8durAoq6NIc4IUd5gCIuKXJOurdJygmGcualbRfIqCPzc+3MuiMZeNyIfr
SlGWiLQHp6ut+pMYQB1hrjPk357mu5qU2w1MZPbaA4MYMiwB5L5hMkBhgcfaO/Eq
7NTcZz4ff5/+T2FhEV/wwEmtaXtKNHxJM+yJ3DuUooqRmkxhYCYgQADa+fsJuiTC
SdeSnnmPnxWmhlwhgFtOBw9vR25ZyRBwU0G5x5Bjf2ez7fb7lWMelbhFrWV3DlMV
V2i7TI0C8ErBFj9Rnk9nOoKqEn6xyhzWy8wz9HiQXw7pGzPXkupLa/yU06unbzaM
jYgnIX0I246kXipQcBin3tr2/viMROMgiWjpkDLubX4QA7sOnecySV4hxObmhPAm
nmOk5QOqrpOtKEb8zcKHXd2/YtvBN/tCuaVl1VFQyRiULyUFqaN7SIymN9zKvt6G
qsODg+enpbjrrsCDbYQWdMb+OA4nGM6jAIIGT1s04vO/GgHY2Z1NqnO+Nm9OUK2I
Ut2CYdUp6CuR8ljn8SIdEgDWMN81CBhpnQsOBHqODxVQvvK3qzUMCKPjChNy6e7Z
KVaZ3dm6B0ijKW1aCDeGgZbs/ip6kR0oQ8fiNHT46szvKo029Y6Fapc5BweOPdd1
C9JcY0K71fkawXXdMKJSULPtdx/OjQDx/g9qzn/8aD0C3OBJjqwZ71JhLKwpeNs9
fs87uG/VrxF8pF4Aitt186XgZ+sPS8oShsymlN3xAd6OG3vHApqjzNSWzCX3uEv8
RbG0hZkO7/40x4PhCVInScTKKAksZrcqQ4vCoKNn6nd2t165duBNoDpaLA7DzSnK
H9mYBn0OT6tJvYhoIINKWnqW0+klqKCM5l0ySyjPMvo6ntgN+uMJhdO26tpRbwiW
lxTbdxbsqvAbu4e/9YdpoqGLbhQXoHI2MfAAlGTklh8rx+Wv/flXuf2Ze2aKZ+1U
H9HcThlCA0qMxEMY/7afa8jl0YChtfWSGm4Q6K/S5Ar0YgsYaoTSmeen4YbSvzTE
BNLPxlEt+koKhvmcLOQmjAO/sKWc+dfnMPtNC6MFycf6IsBf4AeVmOBoUWBDr4DM
ZPnVwUZBBXZuHx0349yrvo1q5mZv79UX6REx1UA4Nd9uAiakuPPmluZNhIttJ2hc
dSXF4kALf7sD4tVecDBIQ9MOCpKHdmCyp8Y6qXeDELdU/BC/Qs7JoxOt2HK+jUtT
gMV80H5ROGzeNFjhAQhxeuLNMmeD4X2kR1OteTzduODa+6o0SfHHGUcthKwX0W9x
iDFeSYjWjgZU2P2oEndO0Suh1m6aliVKW7hkoYmVTkTLWbxhr4sIUUMHwDQfiv4y
HFf/BtDPH/IeXp7Bd7WaZfSIC0OouGGB1hXUlI6l4cAHAyEyHa/j9IsnAd5TceIp
AwVbDOvFBZk1i4RBVqmbkN4Zx5LriZkvKsxlDbrl5Y4St81bsFL2ehcogBp2tICx
4NQnJRUQT3TOFscueqNRcuFoicOP/szeLSb3S90qwKJvLw+kMOyhb2SQz4Y+1adD
FGdT/l4yBz86Yz4vfENS/B+lGaKkOFDhoZ4AR6sYhuMluFhK/r7y8wOotUY2rj4c
lEmR39KiFYHGWe9EY2NmS4Fm7s+RuG4InOis8CaWK8P0HrFbFzGQ9JaXoCrz0nuZ
cxNVTf3hDUPDk2L9WP9IhG0YWDvMYBG7wQ4qj4Lk76eahaORoE3ustC60qUJTFA5
7KVX5BMcUBIKqiqqrhjB8ZVpCawMFj5zJ1Co0af2w5VcxeHcUNxMyjmm3rvYK4N8
Pow4sPVr/P6gJJliR/6n2UKc4CNgDyradXitq8afOrZhjVMh93O/W56jD7wsbARG
2i3nK/PpzncnsFohMhECzCuHm2dEnQoj7vuQnRUvq7mFztxxpPKDBGjAbn/BgjIc
B/LZEW2bkUTXV5DK6pYc+4WWbF73OwtEkkmwtzsIM3EqB+qKM6qQEkiFXdMCcoyD
VyfrXlqSddnhKNKxazKBCHlvoRl4Ip0MD6aFJnvRBodd4/H66Ph0fuU14iuCudrp
j8hrjxbwAsQqaJ6fn+U2TH7W3KcFZDNXEwRDlccMrSpk74o0AGZHVov+Vy5P0JSz
vxKiYcy9O3vTe2QnJaIJV/aMKoeqEF5+10fFc4tq1ZKQaTyltYCYNtHGNT8B9ShQ
Ir98lAzki3LmS4ApWXDSKgGupGgdIMmqoRXaXBI+7D9ebDAXUKLZShm4SB8NBvQX
V+iLyX+KQImB4ho5xtJzUqJLCtQ/7O+9Vl/DPgDePS1kOPx9J8WXR1BRIA+lGrzg
b4xVa9ms0xNBgfXzAGvNCAl19FJw0NjIP/qT5HSq5MY8FUzc4xnCKc/aeWRVjgww
oAxhaA48Ml25NoHYza0fu15EOIu8qaI3Qb1HbZt+g8JZGZjZqN/2R0324nBwilPh
acCCKvKmiukLlLTfaqONuoGHyTONNfVQOQdIt6aAPgSF8Fdz8TOrrZOi240KZPCR
kz1w8n/GuYobTeSX1q1OK+i9n0QJFOq0NWWaqASpbOkeVh7CHoNUx83g3UBCuZf5
5Hv4sERPsfL+TNLY0O66teGDpFBO8h6gV7rzntx2LV+1s0tWIjITOCFHsTwa1EZp
/QH3VNXBkAsYmVpyHyk/ySy++A+hf5KVd6CGKCW8vRFeh1Y/4VTIMatnMzitQt50
w6Jd0B75js8nfwWtuj2cVbCCfxnJnBjM92b0Mf2y3xcpH+G2nWVLrc0KnnF6BtXI
SNC5LiyinZ8RzcHw9Df1xAxtCfmLhE5OO51zBUuu0R5gsIUerzd48i+5dwwEKzIV
qQVfi/zneJZSCSV0P2XwiSKkzj3WIfYalxakHlauBTV8CLW4tx/XjX+HrEVYOmrO
RQiG18hOVV2TiupJRpJVw/Hv4e0GtuoA1xkMcQkhuXCNbE6GfTTssT5pyBWHdF+c
+7kCr3KQhBiUIgzGxxqGKZeQ5Ed9OQtlRAjqOQFFBTrZGS3HlJrp14gSR2szzDFT
2uaL9VrMKZnr64OlbJIWCLpAtoElN/h/5c6w1LEozS8zE8OCcbPcfJAnSPSqHOn1
E7RenSfXGWwwRKyIsyGbOugkmmr1SVhtU0+oWUL8E13R7NIJMuhfYlj4I0xDO4R6
88F2v3lMkWJ0Kd6xYSBAWtzNLWnsz1y7n7/DSag3aMStt7ED8kmwC3S2RfiplJ8Z
N9DZ2mntoi9JIHOUNWPrpImWzuQGa3M7zvw4L2zTcJgKV4g7fmR8rEic7DgrjNBC
T037Jx1hNW6sHh0mG/dVJ6Z2uaCoqLb4lLLP2yHQ9JBrV6NxWEmPknFIv2E3Cehg
gpy5hHcUT6bsdxSgczSnk0zzdG+tueNQ9zGG0xal4F8OwrNZfEFh6ABRHEUZfq3a
jpSoyVfDVR9bRcoVGqENAXl1T0t9HNGoFdoHDNxICHo4aOwWK0v+tIH3wTcqT65X
rD7XSM7FxZJIUnjo4jmYcyjxYGYzV3zDgJMS1pwUIvtB6K9ZHRjj1iNwbkqTJTB6
+yntWfXjVAveCCF6zAk/Taz2XbOKw4TD5ykRmWLPlXH8/CAYDOedj4nKw3PlA00j
tBdWEl4Ffc6l98srzmkMQf7HQQO7GbOjOCkGUMH2CHBBYnNi7Gtv8tWeNnqHw9RS
JdhAWMF3wEofqvTQRacZ3oWmlrNV8XDrUGcpI7xE2fAIoBh5Nh3YJ23/RWiANmr/
NiOSsiO19qqS1OsNp4NgTSPuAFbL5chPLgQf75myGvWLZFjxnn31NH6VnJ8Z+Yuv
Kbhr2/ZmotTb0Afb+5t9Py5MzScyVXJOgtAsa//0ueKsqip2yy1WGdx8MWQwTVQ0
ncG/WqTT1pVp/LHKeDo6hD6z1QW8+41W9woPbPljL4k6FfZdiDLridMqUcWKKmeG
hvRIBOj6OZmRDMGQp2KP7us/KxxAC2j0FwOap4NpGfspQOTqaudQqUFLZ6VkOAuW
XaXxqNzTnDrribJeQ5ffp1jv//LRlJJHuMqS//Gp/3Z/XM5Jp0d2QweGHXyciVFp
R8HAtjYAk9UcLKfV/dZ0e0T5Btl49aQZP2AVWyvZx7Cl7CplGjHMjckgTYAD9iBd
ndhQ2kqZN+wjn/4liSDczLw2Dl3GhyFLKSrwYOXuIoVoSRmgpp+PAt+dTdxOcD+l
Cd079SWRfE/+V3gAJ8+W/mZRCrijZ6/Ssa9CYyuuIi1sipbpudsEabPvvUXVf8dK
o3eVYjFhfm5+kePLJlCPxWkHGqrfQeYtZzMhhCKB0eTRBVCvu2hI448WdxRSR1um
zlnMZ8uRUfPHRcOQP9o4nUdLW8rtcT+1QW8pdU4rq8QBwpOXvpbZqmS4aRyTmhc2
lw2VpI61spGR4AgDGDOgZk6Wj9OG40uzte+fu6zkNs6VNd3k0qjavgkClU5efLPU
fGSi+TtTLYh7FLxYOgSfcAW0FLmSebPvqDXPcoFShnbk9VRlSmez+tZSiJEsVRFR
UgNqOLhstlT5B1egz471GOhjb4r4B8gxsdWzm4RG/9zhgNeczshm5A4Us+AOlsnw
FjSMGLCZ1umcJBO3JjWFWDpq31hO16U3tvMbVM0Hq9CyTQBhvtMVIcv2+pO//VLF
tTXvCQ3PUePemFZDdrif4TM44mOtGSoVubKCio6/kXoVqPa/M3U8Gh4rSYKVTN/m
WCk7QKfjF3wjjb+Ahvh4aoNuKuzHfhGrq8uoEtwzJn7NPLLekZdz7kLdv+XpVlol
njYHyvnthgt/Z8kATt0SS1DX5hCCefvV9KPHOyJ0T/QLc7DP6rtLAZmVWwKc7lmz
bcKKiaztDA6CGvDRbzRs5QUVHoojO5t0YV88MvBjHeeQT6LJS74/kK++o8TskQ/T
JSz/ecwo2/qwyqVeF17HeePUlQwHYZHq9/KnSjep4hcB2Lfw25D3bhOnlQYvV7i8
z9CJ3ohim/Yq09vYYIxfUvyLIrf8X1m26kmB5df3ClidgdliW2utQLq0Ev36PkCF
jF1Zo7p9Gly1KB0n16KJRJBDn6skVwySGN/fXZfduazCXcTg9N9+duM3aDCWxeS4
eH2tACQ4SsQWtfWTsZQmG4JjjglBqE9iuhBwXf7PZC1DmqPDFFlgSap2jwEGUXwp
z5hN4lqwQHuIs0P5OPoCYEJlLnV/mLVzjdjAsnS1jgwpINKjOBzOzjIB87gMMciw
Do1PuhbiP6PM4XPaj8N+mBZ7+6/TW9lOgHcL87Z9WGPnSZp5RgbulaXtGM03uDGn
EXwuSNCVaeJVPuSqq9S83z4eWIMRgBmcdMsftyPFQxQr6zgiasQuxvMgfLOgAShf
lF5yssAQdYa2Cl2DL55DZxppLtoNdG+4RTzlGeHqFy0HbDDUFr3b3toegEooHpB8
jyySwWlO5oU+ItXi+HKPMLIk27XoQbH69TWEVIg/vZnoYjjoYqzofFlN5xSqOA6K
8yxALz+5ZBs6L/tlgZm1CJ5Wze3bPoleUSSm4zAVLvcY7E4CNpZ6Oj9DVFJCmLpR
2cFeNQMNRnJ5zpZTUR/FJTR5i6VCtDOuixfmTtueXUtxo1BPb8YNrTLwmQBBlgeP
5llYtPYiQjpn2C76okPGPC94PcyNg0S5tjnM+Hk4Gv2uZql64mpeLRMG9pIZqjvx
hAZLloJ3nCy7sLcQaM7y1zNkeWcS0x3RlwgGEw/twSFWx1cWx5UCHvYHd838cMzq
IMMu5BL+1TkePugHSCfiv6S9c46AGUNqooCOuOIHgvZAgEl5jjDzN2v9klKkDXt1
Yxv5vpijnKnjEx0VfshKdkchJ5HmKAQxqOp6vVeoYhvH/T2OXIg4kObVuJgSAOb2
6UqR9jmzDgRmeeXrO3rw1US7ZsNz7PJnSvamw/lr5XPtZ3ixmLhbsuxMU167mrpX
+6A/BhiWUJFCMiZxeV6QQm/vkxMjhYwlTqcP2qCu1RO7m3b1eMT4seTZC8D4Wvxp
7v8cPEEDYWHH90paR/MYr1Vsphw7U+vDknO5mDkTddhW/h7exS5MebKr5Eq/piVw
Ohk1SvoUyKOEE7E/Qywl7eyV4OfaVkTR7Y1fRA7g5/mIajui8pbQuAXifyW3xU2j
zCfF2t8+9JPQRislBolRFzXsc6oQFwCSUnoc5/oKzGpIYTmARorbYtn9bOKltADJ
Cp+ReDf78UKWbPIb58ZuWybz3/aCYJZUZ7TFe4meiSyDu9sf7QKY+g9RhdnlxcJS
vqAJeo0K0jZdR6Ap6rlfnYlquk9eKsROY5xuR/LIDldo/LtQxB7330pn7uOXGhtK
A0Uaa5IpTi698qOEScksEcGhP0ktwxTXyzoaUHMvMPgVWs6aIYDPVQfYeKczvmpH
CIaLGG6QYRd18Jval59A/OtEYPBjdjImYxJiC7WCua2aYUc8vrLIoNgfdCT1n62N
YndlIcPXvwHB1YxZy29fEZHIi4kwbK92A9n16a3rIQgrjFH12AbdAFoTzPoAVzpa
FpuP+3Fec6YFfK8XUAatk0JBN6PCL1B6G0uYcXnBbkZYjojy+D+CyS+c7nI1LoEo
a1tclttLtd2cqi0wfTlYlb8OwOcELg7F0X5GDsv6aXFMszrlxtvF5fzzCTAk21oD
eko1UoblWFcVpdes0wWZkEc7kJ5PYxsf4YDQTsV2K/gPDMLegxb6YOCA4IfUs+eo
F19GWzidjWLl1wDBVgpngVNpbKG3MhD/NTa8ccVglEqMS00+1oS/yuIDkVLo4VzR
FeNYD9thxkSUCCRVP+YOo2+Ro6OkVAXM+GKgjgw8tz2ngRRHvldOtLmou40roSQC
GRNutDaVAK8PS9Qjysf3A6cahye89D/pQWb8bxgXXNEjM+DvoiJDXoblJ68obr7X
6ds1ABnJ/pUtDZfY8NMsaOb1Iy1uYHB+jQ01gud4QMtcU3I6CEnRVVBC/1zJ24Np
me8rVPgP7l/+JwTc1ilSvHo0Of5dY5xUaDPzkwGtl7UdgR2mT63CCImHEvsVXc0D
ubdyI5G3c3TsdEQOH4LhaI1gOl3jPQF/nx3xVv9RRDlJgwh7dFbBkS15ntz2rAtU
J4HKQiNsZKSsb+wt7TE05b/PoMlj6/J39NoNdtMNsVuvMOQs0ip4vzxqliFvkS60
8DuqayUu4/9jxnDME40YRIyAOr/WZ7h2u86nmO7xgxhDLSPAzmDUe6UJ6/eeNzp5
UZX2+C2e3573HHP241FzL7t89dYWI49nPZ4xfKC/qF0wpmeq8F+50axN3+skCIQ2
SikZHKzzUcpJhgdzWPNRRnJ12vs4zLKVYR1fvY/wQDgdda+1EIhDyw+wNnOflNZH
8h9MoZkbgFAynAk+SPMkzwc5XEDHQTh0RHEYSB+7dxseBKg9FMTM84Tp6tiuSBMs
BZgira4IFzSgld6Q/6vnv9hArlSMwiTBtdVAbCuQ7RsolONVE/3DMmhTNSlfeCdK
5DeJqGFZXENexgXSSBXpTV9DAyZak/WL81Z3z9esMbNDjfphUFkd53SC7FiZUMzq
8dFBPwKfwMliTuwFeKw5HCyQ8KPKEfxiLYsz4Jxcq6VqAFj+vmEiFYwDqfrpAqLS
qP96t2dQSwI9G2obmZH7oWMVi1l0BJRCvS5xCeQrYZXkhQ5WmLr5D6yjyQ4Y6F6n
n+/WhMPNMosctUawRxV4bzK7u/GOtm9Bxy6REshSODsAGFkyo/iwtwgo1xzNV+Nc
zD09bK/DMLt7TtnSxifPHKEuXu0g5u/i6M2YQafOJ7EL+ejv17cfn0ZbCS+goAWe
RqjPtfoQcly+1cfB9K4N045pc9mrE20NfstTPbXqL33wT16hsdctQIAN3l5VoslS
FqTxrWIsCETrnKaeD2P3q4lWw+5GYkUrT+j5wMiaKM3+9zECvw6NJeeUh2OGEnjO
mP4fQA3++P98EaPKsfZTRV76+BYspz1TgK1i84iqn50EKp99AXcB39+ImZHbPuS9
riWRkobojJJX7HVEViiw2ek7g4dwdIX/kVbNPBP7Uy6fdoYi92TzvbZ0JTt2dHJy
Ntj2tf4Ii8ULiPtCtacZQ7QkMZbeJ4YWCLHTZqieReO5R4Zpan0KY6k5+O3gmAgH
foyRuXDANVFsOYxTBZmDhBsQmGZ0h56/MXOX97XkBYI+tu+8VN7Ld/2+80Qgsfnc
1CxeJT+0QLyv1WSupPgZjiqzOSuFGKAvpphvg5iEmaKGkREfdK1MCjb59P+SWuh1
XWA725OzGAihU+sfkUztOt77Pi7CLujMpxnXcEF/Hd8j7tMkU1glMHEDScdyP7Vk
irYWskHqMa26QRlvWRdUqmY3JRT7ubLUksY+H5FaAZK24vI1qpX0W6vrPiDDatHl
M9a/XFIuUdFzxao/lheG5BoLMpUfgBGylCpuVRgOU+fHOHcbEfau4gWcOzJsz5Cq
OYseUBSJ/31XPaLbt7rbEg4sYcRx/8G6ZsPXvg235o5zSMsyoDWmBGVaElPvA08X
K/fGAF8HiyFeZa2/MNJh57JqdSiRDPeWqm18oTd5HVAwiG4eMD95mFPvrhSzsZoj
vGDk283la+g0XFd6vByedmx5XtU/eCwNYgGljrCdel6X3yfi9PVreMvELOIeSYaQ
MtZn2Nvgs9wlMHB+0hkd3s6Sf+dGh4DPKkfMtmlod77+kCdtuZKluNShyoXIFBee
RJnlo0vBIODzA++zXNCGe23N1P9TnflPG1LUpWS7i6Qf0ojh3IZfY/2NrnkMEha5
Y2s1L//HB/FqWXSrfGTi2xPujxysDMUAvJyI+iexdkz4yxIKJIkq45P/c6VCS/Mm
DalXj2N4GexnrB+stl2yfwu9Girk+BQjTorzzc8wDlck+FzO18pSvoJCp/BivWUu
skdA9tUneVGcdxXofeBVoZNF6g4vl1LKSP+mwuqyJDSsoNCC/9POvw1cD+5zDUz8
W9ySDyWUld9WFnd6ICvGarV/qPhJeo6ZgbTJsOh6La3yrR4K4KgC+5sv4TQwAKDx
/wbDgvnGwjOkmR26gMdR+j6xY0j3TxHJqxHqZJ+oY+GoE/5AL8jaoPHW8ayR0wTm
J7dXRq+rsoYqTdUGjvqN7yVW7Ekbi2/hPC/x0dA/PNNbefJZLAf7p4P+fnXPzSPT
7P0Vq1SkzaeFZXe8oCRw2nubyEXL3dWLeU9scHuCZv7eMSGdmLlXDFKwHX5kmRAQ
YrZajfnBSeLZHeC/sl+zZapPew9XhCvu1H73XTAgpNJKBXCdrAIvAlOjOnhpjIzC
jOIywlslJNusCQDZMnUxEWWJuTMcyy+biaNn1g6PDj2nr7Z3rF3gptfBQhe7abU4
+6qfzvvGXKwblz1Uv3kX4497/UFy3O6JFq9KAuNM77i6eCuX13BFqB1pGfDnVcJs
nIz8ZTRgOlhEjgTUFol7z2RI/YuarvYcwGXbeFP0eGHT/x9s6nh+2UCNUKPxTXD7
plulyBvD1z/nKVLc2V26toYU6S3EnjXxrM9B0ElofySpU7I85pQa36vrpSUahRjD
5+WkXcP0zcscX+AJ/npt4Lk6encnNSlzwG4TpWa/3ZC+nju9vTtGlulMCQxNvXmm
Pd2292rbkvXtrx5Z3C2IK4S//76cvdD96ZGVy44uNNUjbIyNwhg9NahhXae2T/0V
0ybk4plu9KF5MCgokc6C/yGM21+FqNdLK6spXpelRMM4ztv4+NFX6BSJBU35ieDO
JXUaMjXwirLanczEt4/vyFbOB3ELU2b70OAyfXZ+S60//z7b9b4rCel0m+/NEEoF
tVj/Du4+n3JsAKRBnR3FagGQ8cGnt324yxW7kmWymMtANiHRiszFtvUlYEavloX+
FbVgSZMfJJV07WcfGkx90oSKSPSm5L5AOfwPuUM79EJ+5vHj/44SvY+Xytke5Gvo
YeOCUaBfzqVQdrHs/gRJgeesQ1fD2ksaOAob/e6mCvGFyZwQ1UXLEY67Gtqogpso
d43NiUJ/VW7p88DYbmIrky6VQctA0W5MejZuj7b/ZRBCsXomNikRan7NlaCVrO0F
EbM6Mhveg6pk+LQiMAsGTzApdAyexxNzxXaNVSYwVijKMQYigeVMHEsxzVBaRDd1
Pxy2Zc616MAOWHBQl8hh+hk+IjJ6VVwXcJTsWcM3QNeedLakZQZm8u+vAb/LMzCv
37b6KJHOZxd+w1f7pyGvFGC7+n7c/SfYgJIuatx35kSiGyWV+uhfLOh9NmFfledH
/TYUcuHpdnQZpDrxm8+O2ygqBNLOAzX/JfoyN4tloQ7PdX8bDNuXJAMxFf7iyS9k
vllRNQrkEtuKb/8l1zANDZwMWAcYZ2p0EojUfZpWrUsVx5bm1LMxNyHacD9zXaVX
imCcgEtyk8hP/27kIkYV8E9BCrDQSbFmwrmoPthJiKdvLVVyeyMVapJ4eBQqt89p
r6hUTrK+1K8kYuy2PL6co1cOg5VfuJppXjo7LwPbsHjxoLM47okeRRS3h6b8M4cD
Rc/6Q1Hcj+BWZGWRWKjM023OdhWB9LY9X1D0erIFYJyFH71owpBdnqNm3Otkbpmd
WAj63ivKwQFYqa4dsqL5hk3wHnbdSexucW7/133XsUDS6wzmI43OIRczP2W85GA3
WG1wDNusefNAuwNY8SrPlUzsuwmav/ZUmmq+pP/ND/6XYSoI9UtUuvb3lUhlEZ6f
ScdijKTTvcF2tyLfvn9Zd9h7QDh+IGk/JJ+OvzKIh4wr7bzpRue09KC4AMgmroJ/
yEndIRXE0wrsRIsdaHmkDWmLADSjOfGWdnb3ICkkheSiz5pp/kAyG1Xbu6BDA/6A
EzW5Lzg7Bgd1PLrZ954FbvzYIptXiLeEoBC7Udg8w7lLgQI/QDYNjDRGyvvVS+Lv
Ob4BaSyzpWxxkx3qRH5fADKLBSAPc32TMHOvomquloTYG67D/K5pXKjrt60kUvsz
HG8+G4a6P3An4AnaDxF/mZY8RaHimGUBnZqoF7NAy7Yc16GFaXVVDOOE3xL2ugFF
ODabkom5b3qLQ4A7e6HlgHDm6agOJ8nwgAUc5ryLfCNlwf5k+1ODzE4+r7ckQGJa
VQ/kz8oBMg32Ig6Qvf363TNrNhFs4WqGrQanZVx+MMVPw5Nago4lvRLi4MXWWqE7
JNoUJIdv6RPFw5y6P7K8FPEW5IaXmFYQwfihll4kTXnZLRPE88nF13rjL0yKfywz
gBURw5yxwegzobOxhSVdXp3DpNYl7A24bo/gVjcCIrodQqMcut53J73yH7MuSFSw
/NKYkqm7Tb0WVqIQrqnezPBi/QVdAUrf7UgbzoDpj7oDYpJaZl+Qi0GYcQEnuY6G
jPU7A8Uc9iwkwOBTtHK8oJNYeVj/REC817v1an9TY9Uksd4wDUyETnPgWZINgQbK
J0hliOuRfApt9vP8q4XD4lELvotlgiICV8Iux8DbPndRiPL7hZfIh9nqsKZfxVfv
hcNcI4l31D5/p8tmDNkEiCBIjfxgE83aNaFwTHefJKT9rxN9D0X1oTSK0dfcnPAJ
3oBuU4M57eSD5wLLTbmk/EF3hEcevidVcgnmkP/iq4oHa8HomGn/mRQ8sjEkuurf
6bOYvKf1/Y3+3nX3gY1P+tTAhVz3nlHSMqf6cqAlpOZyN30qZWqZIMGsDWRCiRpH
uceNlfjncJeGKaOAk4z6C5OkPLO4abe2+xtz+mbnjabhEfWDnlJc30yAyp8RMD5w
If296wrIzGvsoejUeXNOgO2yU13pCYE8TikYvAy5JzPTuq0t3tbq0y2EBXb2v6Pp
HbygnXiP2cRgiS1rAbeM84tiGESdmd+wPCvvZfBQmbrFuVeIxCHutiMqVY+Qgn+Y
seXM1c+vxXHNj47fH7xbWgjv34YdH3KoHzmfGiNb/r2SX+0UKBXIggxZzQK7aZbK
zXVxvfoHaNgMLhaiu8KE9waP71AufTFHwEn6WqVQwMWz3QoNlYc5GxKHFMsXv3Xb
37DWhr/tCG9WTXE+xYPr7x+PTQWqtWSpvjpe3SQ6mzU+rJcjh4vBptckmO+I0uqH
pABG9yaL4WCgaef8cKHmiaKUpD8ydxXIDVOQQTEOobJ+tTPfa9fAiZA5MVYcUPJq
8ABIUxWanW7VlmpTUJq3ixltYg72O0HnE7uPFJ2nVNxFZ2wQ6MNgpnqc2g05aoMY
Ef+iO8Aj+KtgjYyKOkLH/GFXWIHdL8FsBvED4fwLK6i6mXoH5SRXUNxEdsn87TyT
2UWl2hkmLkjNMi9ciUNwKrAMscGG1flu48MfXwmoEgJE/C/Oxu5f++uaEnTum2yH
RoJsdA0nO8XwnApKbMkSdR16XfCY/7vbfPiu63AyJiDNg3mw6pohlhRGC71wPI4O
H8ZNr7ks8VmENd30/ihHclMsb2DOKfUvyeV2cPCXjuUUSG+0NTk9EdoHnFhnRY3m
O32eSSUHbR79AQICwuCpuOHXduR4mJj+sKyiOlaNvlVN4kM5I74Z72ldnXiROKTs
FenV2I/dzPh06HYohXxM7CigG6UOsj1PA5tlia7eUnEG9GlwJwtAXYN5JFk5vhPt
eXlIrp626XvaPBW5dmj5qEQdaP4bkBj8ugxL/N7OBnTaD++dzciWpJAs9BoTBnKN
JoKkGGFipKS0oVAGvcYtgVkFQF0WZcYYnuJYTeL04bJCYPTTiB2X956+VoSMyYwH
iDCK5zcuXAxVJqKd19XZjzEun221QE7Jo6gxZiEx1U6NuGPB8Gs4cfp14RJDwfS6
w6bIoL9NgP9RjaIPh1Lv/3pF+PYJEyw9XPYLcOj8KUm2czPCL9GlrgFD7trcXGkb
aTEIxYru1LoFBFN5G3YyJtW55vCGKKWKg8MAjQH7Bfd8alB0UTrE12iAbc4GzMwZ
W8yR3xp8TJrT6VjylTRFs6WyGYaXwMdf4FBbJ2Pu801lasLZTP70tar72NzEDabA
gjWg4TeE7UQNzW7defzROdM+rre/PsGj55gEfNLGbagsYKlMvrc8lLwf4oAkTSyg
yaVxnAi+70AIUCrOvQP70EGZbzwrwKVfPSUy3VS3E5z7PdMXGpAUIrQ/UYuhnXnC
S1rvEQLr6f5FA/z3HbnwAFiF9suhfAcJ/OcBijr9Mu5o+Rb1Iy2lmFjaCppFFxfs
bHmO4GWxRJnk6BCkIMM/Lpm/3obaZtiNSoQEy8GW92QdNV86ld8G1JQlKn3STPql
+FdKG429mqScj33TESz2m7p/F5zsz9jT0UEzt3jZtbHxu08tnkqF8EzMkmm5CONt
GGyMFH6hZn+qghx9thtc1qMjRtGxJfJq323/cw8Rfcg/8Q83zJ8vgvE07RYXc+yV
76bZygfGToTswJEKwi3lfQR9yoWVMKQzM8UZl4RoSbjUSfaXb1j2yd81Ol8Lyvv7
c4TieED+sSxeLQ8/6dd5xnacLR/zr74ro+nQ9GXxjguQyodg8gT3uUsbz4bbT6dv
oUw6LTNNMtpJlvrMoDFycaA8hQLR+l7DLKomosrKcnSyvaMPceti9c0OzcySBjUh
a59T0Vshl7Asdj2/XXQpSbto4gOFYpdtCTIUbw+4iDNt6DrH+QT9EqUYzFxppmrY
nNC7uAxNLJtUdhdpgWUoGUmf80OlJSq30n7TlS3982XojhYxnuSCxOJe9cTre3Y9
DSJlgeFAlOp90z19pgahuFGMWc6avlW9/NwxgxGdPqW4SmmgXZpRmr7mZT5Hdb1Q
8mynaPdShs7/n6z3mETT9kk5dudEfaZ+4mErQjyk1iQJcOP8ntRGAXYLlD0BdP60
cUJ53TjDwA4MbcKf9+quklrOGiPvIfvXosovSlig1gSEtFD765PJzA+plHxtuS4t
qy73pTJeVXZ9r9ImdD10lA1K/YVKCC8uKdr9QUliv+v9UDnnPA6g3ehr+P0t7OQ2
pqkn0IfrKdq07i629GXjfnhCQEtNSFNxBomquJlNzxsiTZ7QRPg9dMhsD4weCJhr
WIdmaxE4ipnEZhaHBycsmxxnWHnt79rhRlhkUDT2RgR/cG0MhNv93UwXa78UuqDN
XLL2joggwgyXbPTQYAS/PUBorYbssswFOCnPbhZhlaqe1CZxuyjIugvKraAHitcj
yKA0UeuCKL+/jfZ/+TkeTNRlQNg9OaOwcmQDbNaakHGl44e7zswiRkSjpIvhJtZ0
ZYXGPswprsGDxAggQPjwCqP8vqwARaORkSC9TwO92XF4lUkmn2msWYStvgvdzgl0
BQyvrQvQe7Wty/GcOF4ZaAuwJ9bxNsaQJxZDWhVg2RPMrSUXOrnnjZFxOoQHrv5v
Ebsg6RfRdj8GU+1SMWSxig9aooAm0AC/0fFAJBhQffzKZi9JcZqfYlbHvs7xMVA8
bM69zBAtF7Xu0Yfi3V+O4kyiVE8V7aVaFPNvsHe1VEMKEWHKugBlyD+mHPbp5Pqy
ab4sp+EYRIEJDt4ltYXcpZeR69pWFHg5a8Y3K3Q7nU3NlPPgy7qYik645g2Mt3Az
PnzmTL3GolStRwjMFoZvcpZqUbyU5MO4j5ovEFx6t5uvCQaoj40GMhuhcu14nAqt
FAlA6VbVsL9GyrHxZd9XQkqQYZsgaexdRm3Q+RtgjCTX5rAcLLP8R9/L1i5rSck/
IhbSgnWw2iGsdOooAtLiOuMEj5/KhbVM8XVhpf1sBqio8By9n9pt16Au+Mi/FGAw
Sq4pi4pXK3JXOyk6PjdyANKt2muiK39LAey52KepthfRInOFTLcU2ZwiGtbLZ0Np
pTb2n6aXhwP21HUg4a19OpHREA8vaGpdVLc+BT9Fs6FSHLn6w4qqpUNZh0hT0uQq
1kScjkMaeZMTRNb5tMwJkpmndwCwxRuKb2C7ev2FwTsQdQDX9GkDu6bF5vfVg3bU
XcftOLiv+LBnDVO77nI+LVRFCGOTB6o4Zi59bzBc+4Z5SzSAq+OUmvd+DceYTyNQ
umLFqZb5LeDyjPln2W+bWzcwInhqfcDfTNPB28AgCjluoZaT+aDKNeQ4ulQNlyBI
Vm9mDuRMaz94I/7VCadpy78ll/rlcqzEqDXX/zdgDvROfGkLGWr1rdldPpsNs5Mo
k9pDU8vQqQeEJilqzs9/JZMZn2GclKzia0tEA/CQqCxM1S8keziPItfJ/kk7oDxK
mo/7EfuvLuQQ43wLxnyJrEbkj6DV4mzlAHaAnMcaV9Ht3DDxbhh4YeA19JU62lZW
/QBoFtaztf8cMrsRGuV8AKG6bhOSfuTRUeAIaoRQTWZK2AQNX6vHb22oM7wFX0cg
LgZiJyw3d3Ih3TsihhcuiZLJXrOrY1I/JwbrrhedajO5bENSWW153P61K0oHPBXD
S92Y0pFliJpi/mDttXfQ0I2Vhj8JQ1652Eb3uXV8ch8xfccW9JRjjLHdtzVJatfc
mqbDl1Vf/4YUo1lkq0ZW5LTAOpdIv/6KPv0pmcMfzUWuO6Nk5WYYfD3SwjtvwP5D
1r+j6t2hHvCqX5yt57UsEvIfX4NqGNPWal3daVdBnCUStlPTqh/rDUcCJKoPLDhF
4aq0iEyEzvGYgIpp6qtUWddSYSHLmVzhJdqhU2I4pQp9koiC0tef3P3v4hlZU5uk
a2Tuj/2f9FMUamOIp4sxywN+7UyD/UAKUnYIP7GOtQ/51RDY5Hc0AVFMaBuBY2mW
KS4Z72jVcyUJCEk4E9BR51VN1NZ8Yex3J5kQElrXuCSCf7Vb0k2BpI0zxYlm6je1
y7BIf12hLoTvaMob3t7W3QnEGNBBBFwaH+PZ/pYYJwyIV4sKq+Hwrtnn+ShUyd9I
Sk4WyazB6f376oS0Qu9yS37IZrF8ovl0yyd/qLkKUXXcRGzx6c4Wml0cy2is2SHQ
iKJffUjkg7XtknOyOW3hRvoBr4IWo4tpPDvitTHfF0oe60gJI0PJ2NkBP4AuDJPJ
yxg7d2lKaTD3txvqjK5OhVVsoOaqs0MJiIJLVfa93Jkvnw0b/XYkJDlAux4auFHj
2hDDa50waQyKnobKRf7RKTkhBwMDDJNRhJaatlaIvqyoBSS9a4BeMIaiihp6pEIK
ER8XJSVbkcRTe85gnrY0YgZWQm2ijw1gV9JiADxy9+VwSwbA7rStvuay1cel0a8L
KifwUH32O2FJD3oQ40/WzQ7naTOEW/PCDVffEiGUw4W8ejr+PA3nb6DU9mB8ztVx
mQI6fPv9apFbgpjI4lKi7zaic5kPdmiDI8fqbEQ64UceCS1s/HJPycEgImUQvdda
zuVNdJ+ssMp8XtSBZjD3j3lUpyNTvChx8+UZFTk5hGkt1iF5hjCYLfV/1Ws3B7zZ
YrTX/H04Mm/WPEqFlmgRFB38REP/HhFME4w3gDuM4IYGTVWeACTG1v/+yvnxTt/w
UOACweNtz8qjSkBkjyvK3z5CdwLMZbB+hKXN+JmWuN9cJBEvkhffHz1ep+jUsUD4
KJot6q/++ATX9qaiCwLbbM4YBO5xxOxKZi7fm/Po1Ysg7+AaulfM/Mpobv4J99aY
b1SB3DphTmFUztQklmYm++HUtKkrIOTZHAzkpsfWStntc6aUUkIQNDu+mP6WEyZk
k9SZ/n4EL2zDzII66HX7waMcF7QAugNAVrIuQOnSavZh33B0JvzBiGxMFgfGdECU
NFUZgci77dBCcz8T5nZY28axxqIxxXNi75SGxejAzKG1W+1I4imM4KEAxfbA2iMG
XN9OsWKfhjMmMYk9xYiMvtNdDtvbiRYuPQe5Tc5vAqKCHCgF1kWEc09TNPvA5xYe
Kaa8cl9NGWOkCjTHpTZdIOvWoIRQqGfTwg4rkBJ/Ju+POljoxN3m3i4kkSSZaAL8
vA1n9N+Soo7NwkRAIr3rRPnF1zH5OGPC4gnMfynyKuR4ezDcHcGbui+AXXyeHfiK
xV5ldc24AgIF3wdpAplCLjeE3Qzfm0MKO/VZ0jZ3yctuMB6iyJhpp7rEcmwjWV9G
XN82t99GxBYtHzpFpLfJ9/WspV06DKnPYsn3ktnJta1mmR4gxHieYr7C5QcYoUlo
GLBS0elpm0SK+ZZCqQ29tpnAGPTeYvBH3oY/qJcSBwesG6nY20EkhxSvE8KIqRE8
lehZwIwfEc1gkSZf6g+XwsWHPZMKUdSQlOuc5jloh7eLatnU+leCaOKK5xsFHxkY
u+vt3y6BaX4fEi7gMrrISMe/sn2Chi+zpltofVM+CLuaYTY9/z7pv1fr2xjgocGV
M5VvcRNrSO3iJnOyVdf1YFhjbAGc7kQCFcvJrrIK45gC8IdCmVrg20Lz5M0HF3vD
Je1xNhfIOOfRT/LfSYClyw9X+RggZcq5iUNIJAqJgqKB2NI2/nD+xSCDUND/4Zky
QAXCceuegQVInC0LcBt8jqSaG1EU5MR2TrHM9irC/dbcP+gvsrCOylr5yc99uWEN
Ilhha4q0MaFKG+Nx/Zb6fFb2MsJiAuNHzdAetqJgbG58/NMvoRP4rIwJrmnh5ax1
TPkhU0X2l0/KcL4b3WouoUNu/hVQBh67k6oFqQc6rmwIpokMd7eatwYtcMekjUgn
GaoGRY0ecH3+uwr5f4B7iFBJQs7Cjv3SsfniOko8NxFSZIY3UC7foRXP6JuiAZhG
UsO+ZKMl0zglOy0KsUr2g6+6NuX2S8dRCnpfo8OjjQ7UK8AsI9KyiqZELFQDqiPH
lm30XMJeQnvF5DS3lM2QjJwzSAjeTeBMM2qS5a5W/v7Z1t8R7KsjzviVWerqU6+4
a8Kymwqroy55gGFYpAd7fhNH1yABIrtzC1lMS5aBgdSXxS1N7WW2wAYGSDYfSoTu
3N/gmDvwfuGfefxj8dqL4AXTvJ0C6gqqa1D/0eMQmH35L2CRXUvK2/WBO99legoU
pxM3kfyCtB7IVu9kNhxAls3T4UNJIkly3bwp/IW9bxM2KdstG7GhHHYKVCx5X56h
jUXFZKBk8j6YCQIfpLbKj83Y8XxY7TRbNKmqdeAX8vV6KJfgbFDPO9y9NvVGGtL9
2P0IfakclQJAd/n/Ok7mWYOFac+YD7lq1hzyUax3KQT91CN5pic8jt/axfy9SmvK
7AJFPI7HWhbFiBieFsdXpBlehUGS5QXI4O9N7/OazLHqbs0hMBR5+2ZOxXRfN6XO
QpZ++IQ4n9BFo+yHLA7JI+/RqT1F/Zc+8fyZG4gOgBkwmai/c+Y+Ig2BqrixchvS
R1WH7aG8uTQoeurSp6NxqpT9X1KQiQCaO89oekyQQeB28eSVzD69j+u828qoo90b
l9OgMlafsgeBHsN0oVGfN1arSOXLFxxuphfSpuuTuPn4/zCATqKQ2iyES4nFE0EL
Nu/FSKiDPMzUDd06PIcuFgkf/TnnNrdPzeQ6lKX7TGUzTVhHw30i6ls7y7XrABl2
zG2gkDY6pz1c0XiWGoy1gMrXmUwLW9Bx77yzXtZKJ6H2e0eRxR3YUF6Deh3xm5l6
byd06oxifYb1HcleO1QgRGTGK5ry+mfbEazE2qUBKxM+F0pooXgiGfulw8W68UTO
kZqmxM+AIZZGu5qF01VajuJCdsvwl86W4lVRJk/IVjpZW5cViEpJyOpFvYcag/B1
gHw/+J0p+PCwG7Vb21/U0jEHQCQQvhBSR1+YTzyVOT+bZ3+iKR0vKWpgqImQvPl1
e5+dsws+Xtz4dTgHBkyzMHkaCIl4kj7y97/yf4BiLAziMin8YxWty2U15i7ipk/f
qcAc2iplv33HJm48pUE7BtTUzzJV4Fz33le5azV2RPaZmrPtnTZcuCIlvshmGep7
VI/TD9Lei5d/qz0zOhSlVqK6R61vqVA+9AIBbeBZGtyNqByT3UoIvhejNFLjr9Ck
jZTlVeY1raNQ8Nhpn/8n2tECi039uoTAir5xJUVPUA9wVwMIe0cA86ZJPMGmosjz
Texy7L8+lNGOSj/rA/sgFXn64kvoQVJXPiVXcmVA5QNrBoetcZH3d5EMVHyxWJei
lKBvPPhpGV3Od12TNok3qhpUiX7sze0p/Zy9bSnokdm72TVmqbuEMOk+zlDUX8LI
NN2b7OpPT1lj0Z3Lfw+EW6ByHfC1tEiwgz5T/n+BXbWjOed/u195EkckseF+HTph
JGf0nXJ9zs9ByNU0UXeq4c0TbI27lZvxbN13wOL+YGpYBbF7Oh7FSgVs3L+JrmKQ
jsa3gXewX3NwrAE9f1QnKBXti6V4dFwpr8Soer1pTYLllPZcA+w0RPeNuiLwkqB4
rqMj/P6RzHmOkx19BinnQRR6KrPm7lQNIjRW8PI+zhiwrx0fQnYu2bcYjqG0+RJM
nVrVKrMMHIXNZsrPEosJ5qIoBtKmyDmqDVEKUzaXWxinpkf0ZO7UYoqAuevucPwN
vmIBl69ZURaTWAAibUmSVw/OmF0Z7iMmWiOmWuuKQX7XHVV+KJ2sQW7+sT0a0iDY
VtLNrsBdf7VM8pr1fC3euotsEERlsVANDIqeinEuHjNSvN27dE25wAS4chMY90Ze
xjsBdazUio3/7TlBo2gKhta598gu9CY8zF1lfpHOnyFOSoUsTbTTvs/avHLeygP+
uO6I+nf33r4uDfuLrqd/IB5XHkyC5xdnAJ85vsNA4yzANOUhF/zeV0QeK1H/7u98
xxvRi5fXTlxHJWsDsFRxyEv0fASX1DCygqq/pBBvnuQ4sC8n2GzcU+EWEHa713AD
i7yI6JFJz8DfNcel0F/7CCWyJWvGNfE0kPcilT6VFLejDFNzxDbUZnjyZEtYnGLT
0+w4Yfzz0IcahT2IX42QbQL93ct/bDCcF2bG9sVmYxUsVuMjvpadVRQthDeBsCYL
bSKwt8WFDBLpPgByg4mp+iGaiekhmXcq8eaokMpraZ8NlFPpUi0WCCIfaNV86qfQ
sp0ze4AzWTFQE2GFJZKw4qVNxy48J4fwxYbldevP5VL3QXA6FLBhfgzdydIUwe7i
2n4yTM5leY4hFyN65qwAiTM/lFdq/62xsq6aa8x9g7Cu2XPiP84WGCFi/ATb6IUm
za0pxgWSNeNnrX1AtLpS7tBwk5lNADOC/W3KmENCGo6QxwaZuTBZRC2RbHOeVJ0o
sI8Izv6WRCDlf2DbxMXiFYHuJWwrF1DKUoTuV5KArwTUW2vY06xPCnnU66APIQWu
s3i78CVAOPyCfFJ8gKFV3BWHpNN3+l3Jx1KWS53loNCG8caaBgXIzu+ulUEI5TwH
ddGgmq+2tV3uFzL8txoC1fwnqcvalrlF/5l7ZJ1ry/9zsKBmKPJ8rSQujfZZZ86d
27E5j3G/kLKsbvZoFv8jIaOHrv7W87mFQJ6mvxQdTn4dTpJHra/EbIXdSEeTZOa2
UEh/d5NU9yJ/KBU930R/NHfttSuN2MGKBHjobnFa3ttbx0Mys1jTLGQDgZMAgk+B
oiMgjJXS6iF1+QdJBmtrfIm5bIA/H4kZxGwpBUwtnrrHQ5/LMYbHlP5+13q10951
c/JbcUzSJig9TkeI1/RCnQPXMwAp6lIzMH6afQxphNnjzQhAkj1VGa0lLRRnsTKo
NYj4uZH8FiboiapP/ifroGJnKPJEHkycbH4DhWZ9sf/sqsuGeo9hLBI2R5EvAo83
iZ0xWUO8bLjjQhgC4bvBHN/hq0QGxdUjKFawFHUqlLIh+d452Np9fmfsxlL+2G51
wgT+l47vWNFTy1HUf/IfIklDypxFqjTPnsEccCq7ttuMIkxsFk5D0bRDECTAgAoS
muYAvi09lD+xi2GbDJNp8MqAUL7Rl6gJxWdJ0aMl86NGtao1i8C9xg3qv8lMyK8e
t4VOKEgP0hKdTPA2D+Jq0z6W2pruuDEmFk8m7bm+dwYrtwdQQkQXQsGf7kRQtCx6
1JJC/HBcZqaZhjUCRXZmnFXTvRZwTlKS4VMypD/JIxjildxCbjukzUicIN4Kc7TW
mQDCq+O47IPvWzJc3Do4ywhrCHRPG4cdznB/VY2HEPISbEzVg6zaxRxhyDMjrl+B
7wDIZ1jvtUEafYPY/GbPMxqnSbNzGPSFQGZwIp70xXPn0j/phLPeiI1d3DzUZOHT
TSPSQ3b1G99IAfuxSJcoItENNazpb1sYT/cDJxsAq7xbdfft5t3gmmk+cde28pmf
Sl68VAtM+d6AB6GjrOB85UyNikaeFsqd2NzTg899VqJAGKq7O0pXMmhHS8L4r7pW
HJIEaN5YP5CmBzyGAkiVxFF+p782Ol9Ss6sJtW3g3x2QL1/Ufgto6UYWAslWcwLq
jbGfEi+5EQ8SWIfKrcvOWy58MKsaKm4x+KcAGArgQYv4P319EH8e+uA6dWr9CdUE
B/1XIgml6JqSHWb0WGImBibZ3Hc5vwE2ki1ts4MTDzCRHXkL7iGDw22ZrgWBVt5n
rTKWWsYgXVUeNJwnEsPdOH+teRCRTZjvIp/jV4q3aDIqtfaXk0mMbk8bLcSu4g5g
1YnYXQnJi4bqzVnC0nNT81WdubTewRK+Q3uxV3j6L8YQdVVNZquVwk619iz5Xq6Z
JGociPbbgw7j5ZW+8NytW5cdoQKEkag9FXQzMvQqRoOtgzt3KFJf9kzqPYqyV7UN
hWdImiUAPbz7ExFGmxGan7xZzolJbw/QmG+qgP4aeYr0EdA4K/UgX/lLmjCc2rCX
FAnaS2wKZ5TCQjBS7z0MEPOG4oBz/wmusp/tjlJsr+Lg+axxAzjtBRmJS/1Nvnmw
jo87NZ/DbXQhVWQvum30hQnXr2f+p/e9HH4oeuMiuD+dfVOPn3qOc7Ph7Rtf3EmV
lGfF/M1c6TJXNxbZyegIJ8FPg/hW6pYJB7Rp8+hzW3AmWLRYn0+ckWB8htyrxXbo
PQ7uLDLrO6ldomrzKuwaX0SXtG8N3qf854KuTu3laIndNgN1e/r/V8HsshsIs070
WcmOd3RvxMZmGxxqztawJemLw1V+gBO/8G29IBLgwbridCqJggqB2W15UStdT9fB
EuyDYqdySknPk0hadNnOGYiCk33rXyJ5vr74zt+eYNmoNUQMaZpQ6HKQDUExu6+N
JSyRGJz+Ep84HwwOkYF02YdwOD/aBhmdM9aJkLCAQvZaPURVdH7SpBw+JBCBY6ZA
gFRcb2xJE89kNgWtVnJo2DhX4wSMy+TWR3vHFur9CAJ83FsZTjDJr5BF62c8WNmP
QboI7RewpwPzQiqow5/4ykyv7xEyR0myn44UXJlZ+bEWbXB4bzSJFfRyxu01po0u
9NPlVydO7PfBCMF+iwheMCho2nsBtbUlbYM6GrRcVxUYDbWaZoFl24HwmKKE4FDr
YaD1PwyG+XwQ2v28wOOB7ROKRo11e5gkXM4NFTiq+3BIqb/6kYoexVoZ89r/O8e9
vFfXlrLbMOLClq8fGNYPayyhNAEwPratW9qttTZm0D4CgUhRz1zPbhV+v6INKBiN
Nla6i8ZpZgNPNnyDhEF8o6weRSOzAatYtXdmsl3hW54N7a4Sg2P3mhUf6F3XMeK7
rBvuvalNzvaWP4uthdHkMbQ7/+t+s+DIEtwxZP/aFjLp88qhNFCb4yS/sfQ9LcDG
/ZMzeYp8k++SzgOxstZUt2G9/XytNFHO6RCEADqmMdxzgVInbW+5HwRHkkZjEJjf
ASZ4P6yUq39A2iKBIdQqzA0V2eRpPeStclgRMz8+7pixa/qbw69CLzkZThFWlqdv
E0AwCjQOr4KJDHqcYvQ+oUZPJpLdIz61IZRIh7sy3rkXo5lrUqdKbi5+9/ngZGC9
E0vRi5ptnOWrCfkTA7X5T4RuJmhJLzXLgOkJyXYixlKNIn5tHqXT7xLhjkZB5ww0
lt+h5kytkPKs5LxI3XO2Elnozr6aISkXk8pSyCNMz1cAr+n6lmSX5BMjvsST9qr2
ThDM2n1uZ8Zf6jcY1bPnGDLtw8YANGLwBIgrhAI9MhBUqhUTd8FBJdtA+2FmfNdk
142AA1ux8upWPLDvjYpmxv4GmYoayvFqMqb1J5hYx/Ehno7fSpI+GkJmq78iZnX1
CKm/eRn8pAD2plMjSvMUlkjoIeEXxhofV6OcFOCz00TwiHBQ+lemVQifOj2Lp4nL
idaHH0+b7f+rZ/qoH4vm/haM63lV1BSfJmITv94LPYl6XjANLmmSWzz1qrq4bMOW
baHQwt8dNe03ZxfsMZ4huNvbg96k4BOXD2s0k6vYdoeD94qjbAeE3NFA4/1heS42
XWqk+bginlKB6VmXLLevfuiqyIxRqO+vGCabouZduU7vO9EbUis1UMVGX/le8TkV
QJeRxBwECayEQmtaWgxjrFHtUGQg6lKqGsxxEBOLAEC5AAXyKribU39MUFZhDAtT
QyCEFw1BZbexvHzZgAJrXQofJGGX2BE61CZ6xqX/yWgoTnzrhMQTV5qoHI2KWniQ
j+guhwiRKYlJ/QP5A4Jy3xxUPtGthkJHLD/oELp233liODXvnr+EpStsju7DQRr0
4aSQig/DoOPFkDNI4i8kjXFcRKqK2jqwkr02f4ncVJk8RzF45vwEU2i3N/2k7qER
w+3KWPkFLT4cbt5Og5bYLGr1c8MXX6vtc2ecZ5+QEVxiCkcWAzSs2cNh56XGEmFJ
IaYkFsYoLx0qkWirwVYjeRTq7y2WBrxxZ6Mi+AriLbppIrOeamgwCcsdKZmPpObT
4YPCu4gifaTNW2vIadFtCz4r9UlClqYnXqED16tIoIzWqJ8iD/H3WWZdv3B1E6UX
l1N9g5EKOythvD8ijHJwYzEPj2wNpvb3/AMwKz3/AdfsO6jWYyxEpJ+A2cflEGuH
JCH8LJ2kG2m5QcYFhFs661ydqX66E/2NFy+srQq2lnTacCO8oLRz9JvfbeQdgbEP
iJRTJ2e65cn0h8HuuINcy2usihvN5Dg5IiE1sKQJIx53KCVnpB/aotnLDGoSqpQi
Fr8rOLzCrrlpsDL4RqRn5rg5mg6zejYlHgNwdpiqJPUZr6IbTUFdnG6y3LgwsFKW
j3RbqeuBtQ6lMDsI3kU5fWvwyAJF7EGlccl4UUSM4VO6tSwO/emgCPSNH91I+ycL
SNpu7Fi/DoIsQHmaB2V/49EXBZ28nVHaOcetbcISNBBCgy9oVThxh2U5m22wwmDk
KDs6HYK9byN56MNBXtgP18q9s3vJAW96PHtnWdPz5I2sz+C25qy4o3UrNmS7s91G
JAEgrttqadn6xIUN2lNA2uDdN6E2OhlrgSJEqzbLTPx0ratP+sNfeBkGx5GHwxee
ppb0pNxdw5rZxScSkCrc/YAQkkhVNUGxo0le5Y7rlBbPyDgra+OrS4ToVy/aini/
g4ulX8A+e11R3mQq9atpJvBK6/T+Qz4olkuIpFhqgtDnxbDaBfn3AQXtAw62PrPn
uLCVtwOLuiFUDhzUvq3Vw1yc1V0YOrcJA17A6tPZbf5rSwc0KGN5kjgu1Mj5Ewlk
cTdKAwA+VbyFq9cgAwvstgzj56+vRsImMJnzPFZW9Cu7Zjd9rSYUIyBBerUi162M
kk4hFENk0fU+dYWJ0I31WWXCkFcjg4VZxc3iO6fX9o5U8OYiZW6DLLESKJHoUqHZ
76A4ZCyuIxFxShFkvOGqKS7YDL77oiqx+K/laNWk7P17tfZaMR5Rmd5NAczB4ITT
I3fAcg5Nat2omvjsn3Hw8SJTuhnNItLFmI794fntnOwvMFU4/+GzohU1oSveY/sK
ccxpWBzmlt74E3BnupUZt3PSSbVkoPV+YL7i1aWbJPs5+XSl3OTM2SGJ8ViU8aBF
0qSt50118xOxOc6kYJl4aNtEEcID4eu9UKnVQkcwvgnqby1B5o3H8OMxNKTaJQY9
2h/pmOs/Hb0REGFiZAa4+c/TvKMP+IDeXTtWMoJHDKUjxFevgzxH1W60ZzlJiiZE
0ybP64/mcNkZqN+OyaLRhyBM9SWnA1qvG/wybo40LpRgBk+c7j6ScOzRn+/snWS0
p9BLBN4Z9/x/pIC1Nl1V3IS7kvLgW8iiOwPhXpYTvPcUelYV0TFH2wfORgxAE2ux
H0qstblY67eW7q00GtBHnptdPpu+RelB4MC08kC51dC/O71vVTG/jwehXLG2m8Kj
g/GocZjdbZSkshpDyyLc8rn7FScCjHmGZHL7Ss3L3MGJqFJZnd76W8TNS02RvMKP
pGvbOq6Xf6P9NuTdwU/c64r1cDvrSxP3JZVEkeRpChf/nxy2qNEL11hNMvP/WEMm
UKCCuPqnL0ttFlatsEJzwFX60Jg1TgpHXZev9BUyqFrmBiWpvG9xIzbbaccgVMb7
32dvOvBgDHgIkbXr1gqwJnLv76Sm5pR32o0rmlSUPtTjmM6CZNfKpmx4kHxzyIEV
hUjv5yQRsp6drma+wi/Aropvx4Xz4ZTt+XMTklLW5idwYG3R0dIHneJTUJNk85s5
zja7m1yhFSGOTSgBGyK0+U1VbCp5QoYTXoXUc42Z2KrXaBW413g0eJGeKbcu5qF9
H0QKPiVkqbxNu/t2GHvMOKd0QIgni0g2K0fFnmM0mBP8rb3oSox3PRQ+x//LU3zm
al6VwpmZ8qC6OTLV8LayULBs6tE5pP5qehxXMuqvm+GTl61NiNbDNXLBXfwQhEOj
r36+4+QWIcqN78vJfSaLvruKyCM8Fjm+HsTwy9C6O5cOYMBuJ6OtgT5H+DNfr/zF
e0AvEEdaScAqXY5cow7f0ZoYIYGqpfi+O89wxhTej26bfimLZAmLaHOHF++k8L56
oagNX9qzpPnWeFKvQO3+IY1wfxgx2P32u8AbZiA+7+rWW4jNMa0GNANaQ25xxuZq
aly+BhmcidQOw2qPa8wR6zopWcokxIav7aSMDyJHRiAhgit8SkcdJbjVj3s0QZq3
3urlX6O5AvNBd+44Na35Iu9nJXwyQpQJppHvGGs1sYTa3Wj97fFtwRNYtse00s4S
MAWSxwMA9J4F29slR6hPdKvGsy2VYR8H6fQ6yQvkkC5M63GZJ+pfBkV1aehdimq0
ECi5OQmNJezdOkvMy8ROo7wITtP6to0ybkeUDcbM5WsoJ5+xAVz7p3kyunW2qyBR
znOC33au1z3PeRA2Vug8KLxV4epWtaGEYQ+0GmRRfETgUb9N9g76xOGjFIwYVFyH
d9IZthMa4+EAUDAIrRJEsm46RtK3MpI42fEGAmVxtoLaKm/g8stX45F+ePn+liXJ
zKZyAUj3qrxRbfmEBaG1TRaapaVqFiszjCJtIpmY8wpFX/lwKJBtAz+/wti2RUdL
AQydtpbWQ3xiJz0LyPn0LUKEBjr/qJECdhTGwRMM0jPlEZOrQqSJXyaIGG/zEFK3
ELvNDvpcdGDBrKkZ4Spuk41+bHMyUuBpIY67Bs2odJvLdQzS7IEKg+SZpaAt/un6
Ffl/4EKgGI44at0rveSK1eq9FtFj4qM+qB5QPn9tWXf5HFaEv30ChVAF5Ih9zozq
6C6pfJIskdlTpqb8gbz2qlDcZE8oLT5VGo6pORPtNJ+tdFjhjyg88YRTCLTjfaRQ
GR+b+uVpwz4C+75/uOq5UN1ckFExR7y4SB/5vyJMJR71OKdtOTPqG8dbwODJ06vU
AQMW1szY1sirqKXRPi/C+5NAAPCsJv309fIVw9x9pb7oaoiEuohmCjJWfLSduU+x
AJyRzf/in3GMN5JJtsi+FLbnrs7YGkrEII3+Bi/3jHfrZYmJp4+hK1cHjTLNBfG4
hD6ADh1NcS0Uk2i9wBU/GDFUShd1gEjnMaiO51n9I5Sv4feiRL5IWbeow8l7Nc3K
2tU2+AEyzYu0pZ4S3UhSPsan7JSNQPMFWSkrR1x7TzbOg3JdRYkcbUcds4ZFKA8E
ykGyNq5miYOsfZEh9k3j+hnuyh+T7BjF3dHVqicgdDG/46YNTSKm7n57Irdauqlw
hk4r6CzrP7LZj2NmmF/IV3Cdxb4lBzFKjKYSoYcdDNrdmXRxgvsapPR6/pvLaG76
gyevmL8SpRPD56wnd15qqEBFYIw/R7ykCMpj1MnuqCoSsfUdDWVQNNPxpEsyBMiw
ytc9XpdQVlF9z7DQFob9jX9SUjhWbJxG23twwsolvNh32D8jIBUexnCC1y2O8Py4
6qsZs7aRoA0z4BBfT4y/ylPncRIcIygVoZHWx/Y1am6XMnAPVsm6Uu7NGGteDzqG
xr70kvGLUKkoTjgP6nHYLnvx2JIYxo7S2O/3PBcE2p8e9qwGESlyaUslucCrcnEK
px+XEFrGjob5yULgZXG4eX0LBiNxzCRHJhArm3JaxZ8RrDbHfyc3rD7GdeG+aGdz
tF+cEsyJ1niq3WsbACu5IvYnKAZtjWDXWnccXdAwlmHZkKhcM78fKBT7DEW8zJI1
HT6LEpJXJIu9CFuym0GYm5PIPwi6YQHbsN7UoPrSuPeoqJ9XiUs/rHGuEXsFWU1A
DMMQaj0y3ec0pJ+h4az1SAS77q5W+ePQKf4+sXyfFEaxoZhY7UtSdSSL0ow4R69X
9Bm0zneoSukfJNYsj5qMYnY6AUkZVbwOCGWOQnnFs/ZJMB6M9dnrg4XJzg2fiq8u
3cmZW5iaDKgEz7qVv0Ewnh9WOXQCF2vh9Vb9bwhXFSipx0Ry3SgV2S02mFNpcavf
Dsr0RixecI+jnIfS3EpXOuXgFSpMC8jrP7bL40K08vP72v31PZCxTOHxIRanp71r
24pc+yp1LIq/Uwfgr3haMTWB7CY2xOZvwuv7YS2KUW0goEfYzoqqfRhfrw3EsONJ
QqKnmqc3KVwxjBqeT0Y0zhMwQvskHa032zrNpYUZIJGh4F+/s5nSpVa+mJiAC8wh
adRn6lGjdHIb1WBz0VTR1VeM/mLa4hOaGIAC3SqTqJbHpS2b58VTNipV7CdyMBhH
wMn+YvUpVOz+ZOodnzMJo5CtBaoGFXDr5bS5WPTwVSRMm/l1YhW5KMH4JYFa11Dl
ND0iLggne4kqZ9HozuI3s9WqwuXVxqCq6lGEy/DyNrlm1XyvFuMLcrBx2zh0ALoP
J//si5r8s0Qd0Z0jCvUCO9Ed/cgcMpeqdaT+4fJbCgboADmWqzn5wdkpFy8i3Ggv
M3OoKI1ag0Ls/lzqGK8NT32K60UbWDrKtTSOuJ7cTHfb3UxU/lG7p2ehDAUpwwoH
yRm5jAVtOZOjUWdEatDogeEdDf1mjdC7v6zWFby1ad0qQjcoEiW1TdbuoIhrth8P
RY7QZzsATo8AC4DE4z/DnJUD7rmVwZ4KzDEg94OTfNk1FA+g6I4RgWQkGLth23tx
1VVN0o/p4abSVezJbbS/fZcub96VzOdgucMc6+tllZo/uWCbQEwvVnmp3T7bl07H
1CP86fmtm+g1ke4CI0ZcLaC7I6Hz92O2TdTmCLVojS4+0+tompaO9EQgj4Ir9rl2
MlBhpsxUDeJOdDIbblNGRI6T8v4ky/VquN/KUN7zv4J/9hPlb3/M6csP2k1Izirz
hhMWbBxF5OcIzdMaO+ksnTQbRZodFuruYjsI9qJCod1ddeU8XGKjgwCxE7f4RAT/
Rc1DMoWi2XiHz1SBLQIs6G7Lyr1tpt4msSr/5SOXz/gXmkrXWRi+dHNo/x6VQwWb
NHx0r3lXe+Tu6P+X1/qw79k1nlpiXMQ6yy9jMx74PUPFBW7sDe3aA0LciCkv0c0H
zpfY5Wh3x+P84hx5Ik6cR+v9V6WqXP6KYee1FQCQjUhPaEgQEa749U/eOB/vVWN6
ykFcMW8OePev3VF6cdwRBInfR7Uyo6VcmxXSdwMRQugUzooQt4aBLT1tT7AheVwW
oE2v1rRsHSWbmD8pjKixrhVOAo3CmX37v7Js83C2shPzhDWXXQBeqW/bwknFM9pi
2JnZ3nE3mNvb3qBmb8qgcuIuFVXRmk1uTI430nPkAUaxBz0MxIQeXmeBJDcsgMuC
SoCI0gafTpvzRSn6Fa/jnD/IqWOEOln0t1uAbraBu0Tu4pNqlZfDbqXg9EEwm/fA
iDbjrOIlpi39ozXeDWzfXhzxGV6pDdBi8/XRu20HAR6ahePgFgx0lIeVIQSN2Lh0
BI09hqediPUQg8fnwYxD67dEbIVHaS+nT65K4RavGmeC22HP0awJ+jU66zpLAo37
vWninxB2GlOxk1MmgFUNEecRgp7N8KgTrYPTNePK4LIKnre9jIp3LKLJK0R2e2dR
DcMGlJoUXLM32vVAswZdnThvyNKAZX7R0JHnXhs89iU4rK6UgLaxwS16u1ghQxQN
zjjIRGr4hT5zizjuAV6tXcg0uLznP4hAx4oHZaW6Fe2Hkx0daAjy+F8nhM5Y2cRF
T9GDwm83GR8ZEya5ogb1NEmy2qilivQDHxeR84jSSvHkBHRsOEmlvOsSdqfkJmnQ
bYrpIQ0qiPQzismInmWaSIMQhbinOB3b40ugYUtm+leiF1/FICLe+MO7LIqky+Bb
iiWos25FK9JwryFTQi3NAqVZdT6Zwgysagwv6WbvxB/VsotQaIdazTEilgFAaWSR
IS0ZumJs1KF8faDIE0/3WKEqrlWZAtRvHFb/YkSYvlP66GJ25EmbM0UEBAqgCEjs
Y9nu9XDJg4rkH3D8ahwE8WIVrUjCskVY0uWTihPWnS7zJeBYONBuTyfctgRATH+O
Pu23jU1TmFVnYMVJia+f87ln+BMpIrY7HE/K7sd0ONaxMY7DFU5JUOgYg7aONn4u
mmYyyvObGPxWo4O200x4LKv2SRA02649SDRjZthvHSjTZ+ZaGZJp3In9jJqDnPwA
Fv+z072By6DLwwQxjX4IPSrI00xeBJhzsL5lL7egJfDrBM/QP62iNd+ZiCzxMjnc
RQBU11+VjB2f8K28VPwqUxPc8F9gxtT6AXwhOG+kAJens05FSBcHGHTgv77z8wzm
3KyBIYsIpJacKPU9HHdgmTuU2zLB8xfF6KjN3dwO1xEzJeFAIaU9ZJaR+JEx/JW3
NPRaHfasdAbDTIDnyk57sq6MfCdh42o6YO6r5SHdkkLRHHbFXaL/ClfK3tVa376t
zWom4DxanF1oRlKWwnIL6xd+X3+fN5w7ojw+P1/n2pNHPQH1cEn1LYk8C12E05cy
Jk+7EwTg5rxggkRpDyg09bY24UOaQ9SdVBoqa3fCE9lj4QDg0AY6X1W+pBOvFFdU
xhGTfHOrl2mFyQujHe4AoC95+6syx13XfvfAaEccnDd+PZhxA+RAtmzCZd23fiaZ
6QHO3K9Q5aGog1Uvhyfph08BpaGgy/1dvjp2CT05H0nle2jQGVrjZGhpA+uM8vdb
SAJ44G2mC7m7VxPXHW+B7jkN+BMMNg0Yz7wFs8M5Qez7rv9BMsH9OrhkGU8lu5w0
RZJfAET5DOVBYTb96LBRH0yBvz5j0inu+za0dhTGODzew8sWaGNk0U2hhx46HC5f
gI6xKTOnQOumHF+/0J/lrIy1yw4ad2qNioXOIv+sOqr4V/CAPdjWoIRQn5YbzZc+
Tp5WdWVIYZgSNtYqXsc7Qso1SBb336r9n3JfIjjj6MOIzWvY1OSWxcHGh3I+wcLk
rz2vbKT0xIVmCT6mh5ITvbopsLaBporjyOuIicLxyfcrXXDWvh1xbxP6jHsIwfxU
yW3Sbbrrc2WBJijDWoCIgeaCPwktnVyNMoXS5be+l2IgdL3W3IiR3Id1896PzSEE
HLgdGMEsSpHODdyY1uJo4WZH0YNnTlNmQNOEmrxcc7KwAG1ZNVGyImrtg3mctrYa
s+vNhDD7PEwUzBLk0stPZvI8exNwm+TGWus2EZYMnDxX7l2gOj9wwRfO31R6Z2Zw
6wv/F2ysFgK6rMFm77Y1BK5/Ea/Ay8IENmWNKvhM3iKp/mPL/XeIq5u6AhvrkKat
Itm3qaLfJGOB/cE0/BdEA4LdrLZZmmFeGM3YuWDVjaQkrwvYqVe9DdWt6fD++Q2k
/Xa2A9bTejo4DVrM1btUDtwrwZVBakgVuTIR8tB/8ORXJsbjyj62j5UUKY9AlA2i
RH3wOWDvQCQeXib4bdt6UIVkW9b1MrIDeMDj5XWwaYN/HSWN10zOWMgge0l3+xWH
mtxPSGypsgc7bCp7aKKZrUL5O4DPt1ADsr3NPQ51JpAZ6NZnZKXG91mK2Hnx6yjS
5tElaXX3HRUOzsiKcUVNmeVOLnr2yahYulkSzBtuqdp8B3GO2xi5s25Hed+BMsSq
f8+nszJCBS0yInDY6ZUUkq24pGdipq8+LZu27gdbUj/KabD+OoIjWe/Z83iPgdMR
PMj2GneRZ3X0WeJ8p1nce7KuGFsD3WIf0FdaUz0lwkDVxOZunVcg55swROjwfe7q
Hm1AfYHJ39M41vPRW9Fk2Cc2+swQ4ul+fcgw8e4Uvxn24MLBe9pEgnST7PKT4ep4
mXdIhOcB/fTQFpQfTU708DvBAeypi1aB484o63Nxv/cfF6P7FNPVkzYLeURjNURW
5TRFPIhllhCOJ7rxzMtG2NX/U99wBj/AD3qEkKX9s3wg3nF/QH/A/ddtx5aUhtwA
fkaP16MLwGH6z73ubkGDrGyxcaxn/iS5N+9gae72fEKiWiXC3l+jjWtQb2ono46J
WOx44iAFtZ5xHaWe77/Cqiu682Zhj6QIGQAfGTqij/yBaqpy8XiUruuVJ68ZFQl/
YNzTUutlZqt72m/csESHfwP6VAoMuH+jn/E+HqJvGwfmqK2nNmkOHlM3+i2tyK0X
wPiDPg1Xk5YTD9Gke0sCwTPXEQOy4JhuZ6bR6bXjtJsd5a/JuB+YPOyY/BxWdfXF
XxaURucgVEdRJ/ZkFaLk7nsnxhZEXKaew+ki5P35Rtgbd15Sx1sKVvbHsLgB5HNM
nQKIkGMTA7QIYYD0MXz0P5DVC5Xf0QZl14aad5q8bFyvihHIn5pNzFgDN1n5pb7j
jNalK1XXk1rDu07mhuQhks1zLbHdMAWh9HUVVndzNQSfPQLOPDve9rLp1CsNcPDt
RRq71reG2tNpTd/6ivG2QYYhIIsHnAHltVHTjANAd+kOlG3qDnBOzxuP+RTyfDqy
oPmMVxouTX0YN5XC7aMgijTQsZbk9UfZ7Wg9Sn4bKqqW5kF9N5esqw7tTxGNQSNx
B4eyui476TbM41FHgrGM/q8X5tZX7fJyM37qXp2VpFxQZdelwB2yVUeA1EQxkCMA
OvQ4KEigtqnsWZH/WqOIC/DVLNHe0ntIvKef4G2auzAAyN91hUG50tNiZP6xNiPw
7ZTPQBudYJoJSilPIEqOrhF8YqYyBKwREWElGzSW//0IceKCUuFH7KTozO9S5fFo
J3GBwKciCouYAzyKmGG3bVaCwa42vxUGpidfgdR8/0TBHClzeI5XhAQNP+dhHnW7
qmllR2SndPKYeBo9mh1Ayo28swFhisxuIAN6P4bnn5iEOolA05Pdr1bGKZCa0wpw
alrTYTT1U7XeYQe5LJ27DqWnTgluIcYdAewphRtjf+F0izyDW+gst1Sh+A+YS//0
RVdGbQer2Idt6HSQcixR+8cUmpBqgXZ+FwchlRJD6e7/2ipEGwYBAhF+4pFgeX/U
rbbhken+5QPjEN/IRQe+6v2mqx623aSS8X29ENipyYU3kYoorQMNJDWf7VZVZkCi
8j6lYWAXjbnPqPiZA8ShhV+kNKY7tX/igHBL64q9caqO7PBWl71sVVaIR2uxGaH0
rcuuXVzR8LDLTQznBY1L9snKwjOkkF01E9pc0em2KDkye/tedbt2Vw3OIoz7q6tL
dFyZk7YKKyJL3GsDGg95aw9lg848sGLc+HQUXYg7WddpzeFRPI4/m/hpg/YV6801
TFLSX/BPM/mEYjJR7Pk6E4TnZeQn0G1vqe7eiw04iTT0/Nq1McykzgxjhDcew1Ii
l5sMUyt7l7Nfk5pTK3A7F//O940KDuRXR43Zw7jWheovsZnpTKp8fGv6owc7hXjN
tLj05attlUK8NbpfTTbtXsKJy3Sr/uSmKQLQm1UGyR3+yk0I64DtTrPlU9rYpl27
JHoQvRJOW4JgzCelLVx4XxqELICdm5/1TMx8cxImmrcT2VKqdpWu8epzzjgwWFwd
6ZCilOMgBFUNKJpqKA9AsvTXclAu25N7NXOtwcVE3dINMBrH3VsuMHR59H2JjNcI
3aLM1IQ0jjQS7B+F/1PXy7vpacKyySOudZ2byRwD2G1XxJwSxUkLvV6Caxby1Kjg
cme9dCPo/N1oV7x2NpFRu1F4E4bBAVPqbyBQbzEa4xEkay771/SMk++nbs2dzZF2
vYNdMvaq2bq1LmSYDwhi8mld2+t9oav+4TBRoUN/tNSFgfnrdmGkphuyl2hevtgl
2HgkLFnNJDiYo5+cbMyy1nAxKQ1/bcWbFDUgIrldKQFcRDPD8Xp0JfYpQhdZYVgy
BGQwJ1zri18cQsIj8kAo8U7dpbHIvqZa2kuf44/SLA4yB0Ir90Oz2efbhj35fpIk
GH542lAeDYEo0vCsyIZitjTGV6FZGbZaAvrUrP19lf0VVmuMR1fuoflfQ8toAjvI
DUlijXQWdYY5Pj686zmmSvb18fgnLVuOvhXYMMMYsoeCk0bIFtbJodwjwn226pLL
3rDLrDaDlDgyrzNzOkioA5bntPBosoWInV6StKTMdv9ix79aFubDau67Gc/QeAU3
c1Iji0NTzyGxmRo83Iqwr7kn0jz9I0OYQ7Ra2yGcHbal4xYMe5UUgw/XC+PVed4q
O42zqlCcwJxp7I3ZfXCgZevWdayc663+zfqVzkdkfWq8KHPw+yAkuAaytBQn2QBE
vmOHHaah9Ke+iZb4DstSfSDtLJKOujLtTzpudMDTg/EfGDfhstQIwIhvBYJ2E0PB
HdlUK89hMw8828KJryzFzQthm+Cd+cnWwX80eB2q+y7GLmBX4ubBLMpXcFn4Q3sU
+K9aGMyTz1ZGPXq3MOpga63xkJa3YFn88uEAngzKbdmWPigdsaGu+pQf6vLOT6jR
lZvrPnR2O+i3w6XoB5Dre7yTSh4Dm78b/Z7QQdbFp/B1WLynE2jgziEhToZcW5/Y
92BLp7FnHRg/oZuBdCo59x/qvvqz1ZCXesCdFYW8AnCHe63MQ2e4CnucsyrLpKDT
eBnklpSbK8UDWk7GzqrxKhk7Lrt8Tp9MkHyfQQ2Jxfd3RJOpkkFq13Pa7ol+1ABd
1/+BlGfVzgrhIMfk7GhDS9knjOs8gct9Kyg3iH1c9RdWoapoC8sDHmXzNJiHhatp
8sHqvsSC/CUq+HJS/qNhEPSIOHuBsqLoZgz2ImQqiW37GnVRfrRnQkvJFhsmtgB3
pczS1umelL/vXVNMpkHveYHH0oYrtiLcA1tlnMZ08HOjVfeGyO/dr5zA0JoHDMpf
j9O+WaaA3lEDitiIPiJ6qjJb8i4LR0ZRLUSn7OSNW+g6TwFstv/hwZf7Z3d9HGmG
jldjFYbOjmYfOe6aEqALUlkjTYVOfO2/nibqu+8kmvRv5vy9M23KV94mAlk2v3vK
rX42gFnU9GwVVtFuXT9ByL3t34ATpALbAcsbOyxcTY4TSc5EqHHCEgdBTQUyRd/f
xJMfFrlgkHxK/EAKAonZw9NILeCIGEXWxTrBgZuJIlOTY8IrtAOTbYfGNGIW4oen
rODGSoBZiWsychN1JgtaxIMhHdnh4aWiIbm3B//dxJv4PVU4feQNyfFxrM2zAjP+
UPsEnq97vPZI5byccjvcxGS3HnWXhOC+arfyVmEtx0mJKz4qw1iT0veYT9e5wBu8
q6U60TiDZ8TNDz7Rr21WvHOFV/NLYHh47dEeP9ihpzgi0TnKTz6QwKWhsrpxegdx
gyIjdKr/L7TeeD0U+XPkhZruRJQkTB9t4HI/KKRuT4DieCR1xKJ4fTrMzieZiNjA
kTxClF9I9V1oz3RNVsXjGgJzP1F3H81PRploWA21KdSaOzYGqiHFE5uOFR+ByEld
4iIPzbKpMeqlUw36TFhfxNEBPPkPLdL3TKuymfJLFmTWdpDkkSLv+7/QWyYPTxok
I3YXkA4Fs7iKajHu+40RBFBFfDFHHjeXftq4T5uHeMoH5JJOaRz/1jQ9n9hbNq64
LdORqsWyMPY5e7sWQCibcmIVF5KhDxsftbADyOocDtIkMZ7NqWc2oMcWu+fAiRzS
PHv2WBzTRD9WGyf7quSyNHz39lDofCPetPA+y0BtzIky12mlLafyoq0YO1808rH9
ppasncBoF07zx9LtBmnA5Ld/Vt3qGRHOrR/6YuopfLFLvoZOWcB0XjQWjZXt+vyM
pKPRuZ7PUw4QyrXm5KxiDNWT9PnHd+pqi62GFAoTdJnvMt7H1KqOp8H16rOiVhHj
rYOyVOWtNzhAgJPfiRLnPTSwGrp1IepKMKkCKjo9XNpVdi2Dzn1j6IeE0uSBlTU7
i6rtmsqLvIhqu/WMyQMjjOpkQJ03goaCY7Yodhe3vNHiRPAOCwwdcASiYLdutExu
4GBXOKUKRiwn0WZ18cHKwdJn8LsG5GrqNVosMSkpHCF1HI3d7qRl1b+lGoJQKAuI
Aix4HqcjxjEYaKCfRxWFRIWJW/m23B5RyPhX3iHvi4ahHXKkFqY3ovUa5UDijtAZ
1rVi4kSwvdAofitySRnsxrWf0LigICvsGoifsjTcp55PG+PiH6p/8CmtcWUiUhv6
8okO5YYFdsIGhrBMBJeZYf02iaymWB1nV3u7iy/9mOA/imleUUzW2DhPHbaPbGcw
m241N32aSUsWcfwPtSh9Jrt/UL3E2vMx3cXZ61CYeB+8/q+RTN+OvJTiX35YzZAo
qMxA4kOJ8iktwo8kEl+I0IFJO3v8i7gvBoHaSYTHp4uL+A1nzEpjlQuyv/Ma3vAS
KHnZIqx5gf61X8ggCFJOC9HLSqxU9vSe1VNCSCprW1v9yYQwwTxD2UKpf6eU549y
ejblqG+V1dpFRw5PO5cU8Qm2tYwe3rFUREc2D+G3ZzGiLsIsBs5Mdu4f7XiD+H45
lYcsKO++E1Fr3TMcds+7ZB2qgqqelSSaa45fWD2hoed9bGoEmIHNc+47DlbaYB7T
StmPI5Fqmu2fBmffEGtZ6p853/zs7FMgcfQuMRESHg3T1e6uzhkgiQSvm15tsT+1
D+2p+meCykD3xJsMNigvxsQasuJVHzDI32SrFdDb4e6Ao0gmCIb25cHH6U6lr7ME
vLD07PmrjcKnW2UjcNTPE19sYju1916XIEjOkEIN4I+gBYZRO2lsXkVdGAGQjUjx
mvr5rMJVTccrkaqHT4XRTwN0IF2vVW/R19E9L26VWIrdBTHP8aSuheqY3YHp/4hc
iGH7vbOhDcpXqE2cNmCQndQoj40I+ZCkySu5IvOP0R2VPNrkwtygwj9Yd/NMeI24
QKd22alQDoaLSZ6zkW107FVob+lst+fBGzZdkPXzaA8+lUT0KJCLgp+eNw3TrBok
fRWTMAdrQnOEX58eEW0/wTYnC9vTZRJeW/GjhuYE/U3a0VyTSNKVjhMBsdDdr23V
87GPeHuRhfP4JWkA4B+VQTlIvuA3WQ2kCGep4MujcFOBmWkiEPRMX3M+0MXufork
FleRNcfrvOkZ9EdzSPlRNJEmRau1kfKQKbzNDyZOExNchIxB9RVqRmY8vzAD2Qfv
bDZulSp4kFRtJZ8r01HFcf0Kwhr9L/2HrLxMyx2EbVqHhaEnkTxbiVOc/4RsIqR/
BZktU3g4hLNyTfJPbLHJd54NKh2sYpsX3JZQhe9pgqO7ZLo5Y71gSCRh9ZoWV5oQ
as8VH4vltcAraOtTh3OyXZgQgWGxo9djGxcG3CMO81vPAp8Ke80VscIihEr5KQJJ
Q7mI8kuGbgmXfPOIy84AxPELisJQ1HSbFXHgHiXltmQeFn/l+QPeulSeh4YQ7If3
fQQCYpEX1rJv/d8q//1Qz8guJG/orlN4amlU30gRdh9ra22/hyG++oGVMq7LOF+Y
XmIgyoKVmBwTfoUDPK151WkH9ohO7LSdRHc51s+FQRxrD93ET7jXnxeHYSragN86
Kem6cPUFgI/ZYJNBPefE996sXF9VfASaQOxd/RWEDNNoOxctQSlIFliB2oWt5p7/
aRvb69JeUh04GH3trxdNJ266Lp2Aiv2peYWzwTpvwyDzbh0A0/4Xxkx0Hbexz04Z
amKf3x/lD8RLNyksJ1CiqBDkD+Ro1Ue22tXGB+MvURyHgo36ry6zT5wumjDsi8Xk
0piAK/6mAfk/BErTAjf0agv/MWVokyOyo71QleakDgcRK2Qkul9M986CZDnPKmib
SPOJ9cJFRymKJfhfuan2kNs0T2jzepf8Vfi3iDbCdsBkb7JvaeCOXEjJlR2rfr/P
LZd98LH+wIcI51+Zy11pefPKuniCx0c1QjgsZl1S8JPiCFWGWYjQgJJqzdfOMaMP
PvCwqsS3xokhClcXEdI17lK9ahsY9phrsnwxFOgqe4oqor3njgJFNoJnfJeKRb/b
cHZvfWmXQstLPN3qGrKT3ljnJnLyXQgGVlP/c0oK4Plk7u/M4u3Ac6Ol0zeZ44zi
B1v7fSKtXkcYuloJCeCpIjdMGiUnhMQtiyBn2m7HDmbL8uJ2vXmdXuHEIBJXWcXU
yEtEE338AWokOYApz1+mBl9vtVpOW9L8ybPmpkI1DZgGFCHalyiQcnXqLdOR9OQT
r9wDx43ygjUfGIolXU4ctxfIDcOpZfAwt+p/GPsTCDAJ0wSAskUzIeH2mxiIeGFT
tImJKyKmr8fml+MbVcQ6LlvIoTprpMOsnJPE8sJd6EfQGcVNwWlLRAoSLikdrj32
sOV/jwgMA8NeKmH750g6CNzJyrff2dBi17u9QH2RxnyXE2Eq4iUa++eLKhOqqK2b
k+MHCGrqf4qmIaeHs8pFyD3OGp4E2sZcop4r3p42LCLCb5VDZel3poTPZcJeqrNz
I2esx/iDxZY+qvyL5sGP6xdv7YVHKz/4hNKCZr8mT3PAYWxDZA+EFVHgsAmNLz5d
umuUxv5hGwjVgJVvYfzH5irsfKLE83qmL/uAVVUeT0Ub4uybZe8e3Tsj2wMyjNoC
W5C7+nFXpTI/dUBgMFksCKcdOx84UkHSwjsdQhmuuEw5Z9kwiTlFHmTlpO59Bac5
6/Rg88i2S9u3F1EjVaf1flaVn+2Bql/s0gJBVQTjIdmJCEQEEIfuDLQZYLo6hCbM
UmNF4e6PbJmfIBU5LqsperAr0/BuCK+6/cD9+wiM4SnIt0U4/OZFbM6mbDc2vtBP
WVr0ePCdjkDu97oJSYP6Qkq3MXSOrC1A1C9cAsmDuiXhgXajMM6JGrdrspZkpZ5G
60RFZIzpPWExo0+EbyLHEX3uS49QQB0RMABnv8njKF3Vu/ek43e6FwjcmUTRwmJL
Ne8xw9yxxUZQ50KzYt64OxQLRJSe6psDh9zQ3YFqN2Cwu2eNrJYWZh76TDLmNiMy
xy0qz/dYlLlS6NZPqtgW74+L/qgZjmnxR2mDbPN+Tqpw2W8JtAoTuPSK2wXnMLhj
IDoafYgoyYITC11DedV40KkgO+wRLk6+gLA4RpKJrur3I61OmDHXVjkPNAeMmb79
g/MGOJA7IbC7dTUuKSfFP8blpdNEiF6KIyOYYa9bQynVEUEMf8/mTOY7qOfkKVJv
ccpkIwlIQD863iU8gU7e6ZrtHWzRRhumqEF469LiDGPWwqLuWsQVXcvBBGdqV6ha
mXYkrl1vgzEHPfgd/iiLbdxtEOu46ZN1AX/4nkC8QY3gPhJppfu5bbMlewNCOUgS
3Ae93Fuu6TpI0b8nAFQsmcuDhRwfiO6azSGcNoesl/dZXL3WqBzIfMOfM1lk8dft
LL+yKGLQbAl58b1qhMCstctSXUsRl6xFEDdacSRWETIAlt0WhMzGj7fuyKPdOgfa
YphcewYgrWzx2iPw0UYQpujdS0Gkbn2amf3OjXvGlbtIsga1wNeiD38PfVxbr3f6
YarvnSNBrRdXQL+k2dWN/lzA6T5d76ifU6H+9UXPYemZwlf87Yxz/SKAvnfhbr9p
wOFJHEjdnxfXl959zMFgEKsf6zM//A+ZTW9NwKZgXYFQZMKXcj9PTcj7WYdKCa5q
YXymm/6FctWSbkScxhQNaj8EiWa4veuBFAVbeotBhS7d9Ni7uYUSqNdPLQyNDrju
KKWM/+v8fjfoJNPYnPW6PNKe407OVVH+RVa9FKpQNJsjbxzZSWM+SE+ThgJ9LDnC
FMcsyxgeVuaZTydlpk86c04FbgaZ9L60jondfiuq1Dh5TUSRe2D3EnUB+UKia78l
trIuUWci8MM2zDC++Z0Y0NoBdLSWj4Tou37ZvGFrh0pqM/BN/wOy5bLd9vG4o2rb
XHXQnge5L6s1C4dL3DrOwvFBA3l/VLWeESS5M8iIojWEHjaF/8bh0C02bbY6f0UC
Mzv1GHLI9pnAeP0BlvSag1LePcgnSsSJb87txOntHEaLUIaGvLdmKzYVITbIvU8C
sPOx2MHGSRxIpXfUrwqGDw95kBx6234vceZ2i7mzW1gAhyeBVzidbSXh60AYFwrJ
Q1Y70AJlCZHz3zH+bd5MziX5vMdub5jcKvWsiuhDsnfb4b9B3grkaa8+u9RUklRv
/0L9E3eMWubXKqqEK95IyD75BxUyvT19FJd9NwM5VsQm4Kuh3KnMCGbRBhOeNk7F
voE5+PumrpzaOHKZv8geuOLOZhNnyZI2hgLbwEVFHSNn0p4wP9o0xvtNGAqnF0Cz
vUg+U88+uEOcKv/+CsemWt0Q5bbj2MVT+lk+d0YasPIm7ViO4UOSvzv7+Bs+02IE
H1v+lGHE/hJcyqwlJaoYGu7vMvcjcbmiEH8ws8HwOfmQP8Jea0Dz2XA0xr9ATuVV
J/nZ+bg7cYtwPZY8pMaJ/xf5n16F9vUK0PpMHZOUpF6C3KlUBW5rSf7rC3zsNk/5
GtyaMBV1AKqCImV3tVL6tDbdf00JgYHwq6y/A3k0/V2iI9WSmgHeGCIK/r7UiwDb
3vrvyK725/lbLzLAMA1dXD3DlhTA+7iOCX4QvsgmGCmSECNFscuQGtZiM4cFfU5l
piB2jQxiYNhzHwIxLBxU8UVJJGw1UTmHuwiIi1hLZngBoOr+kAKFB3hC5+9ISuGY
TAmXQz1pD+WANmLVuO8f9k2nDHgwLoUjoq+9KMp4vvLHisrZJqrBKSLa8t0shIOo
RIN18gAC4wbEd6pHOPEJxMF7Ml5li38YffAyqwVS7V4gcv6h2yW+/st4PViungJw
1s2Axun362X6g00oKFGosBdIAOyKEZDY+AHQG/g2Rp4ZQfsjj1F58WgdkaiywyxH
cvwDAFpuif4wXDgWz+EIm/GAjwkvZmmEuE1rSMk0jzR+rjF2LVu+Ux/tv3S5Ei/V
53/ARLDNFWC2xSXvhq8TbIjqL18XvgqwCiGpvZnF5F2ni9BQdb26x216j3J2hQnU
/b1eU3PV0w19Q5LVoM25OxTJ9ISO/6NGl2dgT6Eio7Bu9sTK3DgKwifnwgHr2XyA
1iQAqgLRtNmoHeibZ4n+re3QWOEOfoVam/MJtRZI02Pnl0Op3Mqnw1FzLJYwqiNG
dVCOCPnBwRzTTNuQrO0ol4F8MEyno40tX4vx6OSVtJuPusdLv5WkQutHTm/0EJ2N
Rchhyhv4mB7p9Q+Ozf6iDsTbDsY9vGI6fMrwWQ51YN3UlW4TRo8dZcJYWMi3YJ7u
OA5EPUf0N/JG2QzcBkcYuECPWIEs5NjjPPE3NdJXlrgstEi/HF83XiRk0g5NN6lh
JCInpUzE4M2d3bDaK3MNYqik4T1VYcAM2eekH11BUULd1gk4b3s3aJqflDiUmezn
1wQn7qnO1AD7qJ1mkNK/9CQCg/zDKSx/cgzst7I4NJ3P2JU5hLBKAhqrbU/Y4yEL
I/yMeIOpofPSyjNoozgtgkNTEb1PBe8sq0Y2iyC5e245/3/PznQio2kP5weyr9cd
/35xAgIGS1Yj1FV4wosmFPtdOH5fR89w04YUO9YHmxS3JNfYVZt8pvIU75cT9gtP
BrKeEDPC50gMHh2QZe9SThbGUKk4KkrZ6GpYTjhXQESeXiQ9y6jw4UE5lq8vF3pM
sMPSMFRN0RJJsEitV7lt0ULDn5rluuWyIreh5Giu9AwpGc86Wap2HkCrvKaQFYsB
YuGtM8ZWl5afzz3mU7Aj4+AZtSeu/ykfSPH6ZXoPT5G5/uUAfmQ4INA7K8luxevr
4c2bPDCGE5Du2HIwFjjTAVIrDRxUjgVUdBRjbCR1GGrlXNkTSHWGkoKymdTNnwJ2
4rcDG1I9e06c+Sd9zy1VDZYYKEAq50GMIEtpC84XxByw1aJlE+6RdFSQAQWU5x7R
fhLi5MMIkewHWgE7XdFvmstffayITM3aZeD5TZCjBoDYLzHez3y22FP96DTmluc7
LTJN9nntBmlqJiOlgOjEzQa3UNpUI3frfwcieq5tZGVmOR3RzrJHIrnAC5fnDqtW
WQQx+AOLXb3tRPCNUUAOKlq3wZRwVcLnuIR33sYRD0PQno2QHk0DZSmfLN0UCrFk
qkjtpxx4YDyb7VkmsWqC23M2hScz8xRu1NZSHM4pnAjWJhdq7G4LFdnhB2V9tFBh
0bUvJZe7PboLZVfvnETaA/+fYLI78QAiP2Vqo6P1/ItT++YaWRI+2il5XK3iHh0o
WSf2pjDx5n+POhflOQ2NKAe8ZXbeqKMbxCr5+FS2C8LjYlbM6h4h4KZecg9MiunN
MROK2MdQBC8dA6m8r2/Gz0rUYkc+ac3DyfoReIzBuktuHSy+0DP2TEMEBQjPTR5i
OrXGpK1ZlPzh0T8hV/fRqeqLmZv5CZdFl9Sqb8SJ4UIAXceU2viBmN4Hbw6DTGkT
hmvHdBdX59qPKZE4HPw/0G5JugZ5HR9ZVzSbtlRhGBWn5mZhM9XLmrJuyuAZDnEj
mPwUAUBqKSRFggnVEKa76thtcNChqQNFIicHuc/Vi3b5614BjBVhC+KksqTm047K
gB9bW+hRYyBJA1NnnFbrry1QKyPwOSHDBzgyOlPzO7Wip3jNjcvIFItECsBU4C0v
PVwJODnjbCgN0Ke912iIYqJF9nc0hugkJFbYXvAeOmk+kr4gwgmN3/Q+fzkUwHtq
EI5tZcUPNmN5+TjGOEhsNr6wlQnELkIr3dpxgeaW47XJ5cIyAZ130V2uD5htAJCQ
HTpZh5IO91s9kBzZeLdudPh0DN5VV2cYi0RZePHdX7HEeISX+xWDy6eFUtXFcGdm
ea4nOqpbgxeo3T9AbZ6ykdTay4T3hf+pLMVHQwy4KkQZ3qDuHDrFC/exLhgTmnmu
cU7ulFs89XeNFuVHGlQbZ2xvjMZcVTeoTSm97BsmcI40bEYtX8Np5LVj3ZZGzzgA
3J8DcA+50uc0P1RTa6KAFEAPlQ/rYMKR7Y5xHUxdzzb7WB8J+5E7S3Cgh162g6lh
YX/JVYb9f7iN54/cu9h0+Dy7pqEXaDd61y7sfWxINi6tbR3Q8zjWXgtjqlnB5zCC
oJNEgPFHYEsE5UoBh7c8+SpPqOlfP23hdAY+ZEzCJHYzlUdnLAgPpZdVULxJHI9z
5yKAXjZKSxh2/E15UyF15bFMPYw/9IVku9BGdzQfMFBQsQNE0d9GlQUooiLMtkaG
s27ZbYv4wqLqVB2lhcA36xa8yuUXJVs5Mr/ovfdcb8VztDQycvE2sKIpJ0pv5zND
nxGDWKujRkt67eSnv3cpcu68m0wF/ytVomB9BjSKzRl7QovQFC+2BWNRFfixg9CK
jCBuLrMxD2qDVgnaTnImoKuj6RIQDsgSkyKc6eMqysc1Vwzgec8pt/CgLAW785Fw
jIxsKK/EwAbLm8Frzm3dGQc/S3RYsk5NA6s1GMLkJaWtDA90/v1NHwyWc0poFehZ
arIMPWdtYqITL9Kh9/JfK3UfdCE7zfHsRirNbADDB+og8I6S2azWNJjhE+8JZGna
wLme+fYBtE5PZVcZra+b+vBkC/P/ixvwExlBnpDLXzh8Q/ldhIIOC3/8Ybnys3fH
a3KF7mRdA7j/EsyNiJozbymFECjUyz1czAknqWUoNlA8qrCQCiCMMgjdcoESGvw4
r5p6Sq5TQ53c7EEAflcHSFvx9h3/zmJLzcsLcC40ukCdQV/ehBxHcCRJ8REUk5R9
G9GQPAlptWybccHNdAq0A/dt3tf21uFJAU+yY3AZplJuklM1gHcxQF5jbjS780Yl
bFFcZlxiVibzFLmmEZVWOexAwHrgNlYDPyD9qEwO1WTh5Tq2uNbI+aZb1j7fUjDx
gN3kRuJfONMxKsv8UKawHJY9pZnzhxjfAGrrz5g7xwxX631UyDK53Tppimw9rcTl
RzeLfuQ5AcZDzXrKeW8Hxkemv5aSINVCAg0MtTn1wUmdRBRMJZ9e/i5Cy0q24hlN
Z7+V97ECNC8bDQy3IUuQbNOowYFEgDJEeMTDybuK4vpxqXdOCVtjKP0Q7TpdPTbH
2kAvt2jLANxNvrG4sqWUO3hYuC06Ihk9N53DT1RJL2lAlhFFI0qqEcHrxrb8Xnq3
0AOrU3+nntJ1W2xyblLe5Y3u5LM8lJW+9IShN9FJs+k9jdL4qve84CqhDG3NS5w2
QwKKXutr071aJJR8neJDYFPo/LFooxdaqQ16PK7FrKdyb91UGxrgfRbF8Tz5/1NC
VkCmm3KuMz0pEJyPzmUKkN6muLhd6/KV8lBpE0j/ZMiQKrueEtofgu43TQZZdmqE
oKB/mbOi7piFjDsZTg7+0C3bGyZV2+xyR7/xwrZQ41P5NdRLHRK65oFDjqdp0ZiS
sl1IjMwKxQKS9RZ8cz7s2OUf3umLLVCByJ/fbWVBXs/0bBEAR5Ovhj1jgHlVQq4t
WFBrMUQsGjk1VwyMD6MGJXrlpKCM/z7HqF+V9B2I8+AADOuY7+JbR+mc1cQVVnor
Ry0SsINIFxavGW8juZRAiA2IfM9Jia6AKIwiLCiAU6rH3VyuryOehpm4z1GnN/vd
C23wxLiucy2IpPEXt/Qm5wqASY7AmyZmCduDbQLj+1XLiYW/zQLGk2ObvxGoWQdV
Eiiuri3ydJK4rGKHempfhEdIEvyN118Occ6CJ3QeSiXNk2xoV4oKTVhEjqg67X91
CePQfUiHldDIBaBp6oRYjo8go4npUBkWbeUo+qdkLwuEF0N4n73zhy7wrz4pOsjt
oMrJEjR/3dZfBmxovk2yA3aSNFGNhsN8myIbcl+IWk1KORlywNkcjHDGEv0Mfs1I
gTvQo/ZZKFmcxccqYEPkaNDORYxrWzEoKkRD1lveMXooBTdoNhDSbuy15qfuJFKZ
+S6MmkJJOLC8luZ0yzLyWHabjN9wOq4DNJg3v4zZkRKmndAOVKohdMUtq+Kt7t2X
xr+EJ6hqb9rZ+vxjui6H6IlbfpAuTRJrHb1h0i/8XANr9cUw/xfAe5T3EwmEp2Fv
+Fczu/pskG3h3xh2GOlkN6zGZh/gB4m4mn1CAlcnbeDFmiz3XJbW6t4hnS4hw5hb
xqau24pxHcGhtNqdBKndXDCAhT/xqOa+AQYeDW47f0AbAm3JHT7CEjuTHC9ZUvEW
606pRLsxL2d6OXez1rzfcZyp4pYLsm7eQg3VUWZINuLpDvCmp4YN2upoATpfmvDb
qxvf1xurCifsWZDmUvhcEHd3B9Ph/lMmFsS1aFvkAws2/LiKCKmCNhK3HMN6FCkh
3BhDi03w97ZUiaDsXWV9olNwzzLAzJeaXOFUP2zdNgcbXmurGMfk0Y//xUKQD3su
5jqVNHmYoJdePdmGn2rk6hkgX9kW+j/E1feSrdhKYwBrrXmXq82jJwR41aChjk2z
4u6Qqm4RM2wmJFkkWHFwvl2Ctf8LnQ/uyDSPWcvAoYZxTOL6R9wjzikGKSKNAmXG
QkdV/me8zmV/vUd04LB6JKx3anjZmba0z/nqOptkdGL9ccM6JQ+qv0lAp76iFY9+
PP+EUuYIHNeOiSAoQfJhw9UzxFs+Bodnz3HTHiklJRr+9mre2IILsqEdWOo5peDC
C+DJVG4wAtj5II7NjHUtfarsnoBEK5/fiFk5y2MBUujD0shUP/B5ngCix0PwvNqb
hkSk8pqlXTJYkQ6EfILHLFUH+tJmWl07pxAE5rFI2SiC8c1iOcH5QsWUccf1Knar
zHucnzHzrghpt7QTacm7HyV2BlT56zbR1gIv7pOeamMIo5A6JIwJxXMr781vmV28
jqQRl+lJ3vzQ7Z+XVmGg7GTT26kl4pErXMj+tIoCFs9rmK9LK1vx+nbJaLAGg+tB
sbVCn7mMzYsnFwa8vBvnt9jGhEf8o6hp0TEl61zI+tA6vwwE2njy2IXTWu234wK6
96u134dDhGReuGhxsYAt2og9kfFqdtPCsSChwgDnJUqN2ylQCc1dGqI1aSR1i0La
fNcAYdd+0THUFC9ppbwMs/qno/7DKeSAjalrzPayg3akAXg6aULkBA52mV2zqKP0
n/XTqCF5Vy7YTalC6ndsXeDe3QYSG48OiktP7Jj3cx5kxpoS+jA4MZp/8MxZgQOG
O0Abtfjmnh9nyIXI1ETvUHD7ykXtcnOiMvh887rjGGerDtf5GHbCfxKF7on2eigy
zdx4JH1Vr6fHEqkEX1JYBOySq1E/EgPqMH8fuKBULEbeMbz9aR3vJV3kuJM3uVrw
UWLhgqeBNZh5Sa91mdmSR5OAloHZUY0R+Rfp7QIJu26fe2aXS0Xv4vCOnOfA1iRn
hejMEU6aUnqVEq5lyeUeYMPD1vIFNSUOQydgszCtaV5JGtiHi10Kb3YZSmLvp6De
riVlB4QO+zRCmsLQpDdYsR6gvZ8snWghcIDkBd4Z/k7EHx+5WjXv0T2RT2oV972c
TMnL4CYkdqOXO3nRyd3XeA0VMyab1Am+CImv5pRavtqAb3YIq1E+/QKCCBUaD8/Y
wgv4wFx//Z+4LpBnArIJJPTk+xoC5Nq86GcwkiIYC+L9PKCm0A16NNaLEhgJ4ZsA
2//b9M9IlS4uOwPDjnxmgxcLh8cjdgyN2cBR0zQUPVDiSJXto7x4FFmkQn7W4dx2
O3XpzFWZts/F1S5zMnDiyr/B2N5uj8atFvpMclKaY9a2wDhUD7fVZ5QrAzVgrizW
KUSF7CAQwLKk3TKpLGKSvFK+M1kQhDufRRYugjQEJsA1y7uj16QkKII1KuzPxJBN
tC1OCx52MkD9GLHO2USAMTKaYx+f3SG8bxD7lwsUe2Odq+mRLJLTdHD0Y2kPBVgV
drTfDHhfIjNIiHfiekxOKvw3zFE6+guTfKuC/SBlzXNuV7/efVcxy294YbfHMMfx
YH0wYNdt1xJI+Gsiylz/oC3lKQFpHZTDHsA+TqSM+yarpgN22/ObGp5PMzNlhu6O
zvec6KwAM5wbNam5UdCSA/2CYlqWrH7lbRIzr3Vpbfmm8O89Dk/YNhmRNzTBezHZ
TCKAtSyeWP0l0VG26RegfPKot4gUkeDqBfxua/h603rgU/CjM3jgKq46W2f4fVkJ
FCwan1G83Cj9LRTQwdvGd/5AtfIUjb+qUqjaZSJ7JxHTwy6fpo5BabmvYmliqSOE
JM5Wt043GSR0I+KevRBqs7ieqQ3aTYqzOrODTpyfk9mRrB/0UaYb5W7WPvZu4Nfy
HVyvy+uMd+OJIIBRtrI5D780cEEIi1njcGm8aQM894jB0rnbyrA1w352vVFUfVXQ
VdtCM+6T9ts7WKqtGwdhbNvKx6IRUG8ZkljfYDBqwtzWLJzX0t0pruOsAmbTi4tE
UAWTmm/91+o3fPuXC8pJHYg2Tg3xGxvgrkpfeEL496GYd/klz2ACIrB1l0SAbDrs
Syxp4tYwoOeZqbHYsb7xqvIa24eFUrwd66KV+kfFdWlRBw/IJqGI/lzf8FA4iBzc
g4oFXskg4vhbbKyR9ezAbtUGQGB9qRBKmSrlc0tmzonDCoST6+uJj30iy4TQ3+gr
Yxt+11Oak82xk9BajHFAWAsVoWRAHAiOzAdFjXTuc73MbFrV8pUEdfDfvNj+r4MC
zrwDihHsf4mjJhNkZI+59x1mGDqbmToUQX7JgdtSpeFqievBYuweEm//C4vZqmGz
eJ6CYGrYzrucg/mX5yTyBAg0aYlGU5+vb+MZnZ7HpJCC3/bAQJlLd4kyi+By2+VA
TsCCwdBdnGUbiGd+gudAcqRttalWh5/d6N/nFNTZgaxfjD+4SP7eCg+O5NlUEYPl
LmJidWgUELhbGmPAV5mSShSbOgohSHvmwpisDd+jqMCCTpdq257M462unGuZRwYB
ihwLFYwBst3lFNFsjTH6X7KRioKIbPPCEFWoN2tRqlUsPYD0JIB58Glaa8tL7IE8
RIZN09p9dxdyp77eIZab6f9rbRJykcid4haJ7D6/zigzmwrwQKVIyN4uy7pb/AR2
OrgoBjwZ9BXTocnyed4dK78PWS5Xg+1ZVmo+2eXIFt4sZcFqKRLCBzAyLr/QB4Ea
5yjFaMpYPFaU0Cne1EJIgd0AN7vJx/3Z3W12oHiLDFmoxs00G/UCIXN3A08z52in
CQFZy/zU1YO8uHdBEZ9ys3o5t5d2609hwiiLILONv+zeCBNkxcGy8Rl1vxMt+7oW
QOwrGI9Uul9tdgNGx3IOpviCiTr9szWeekgBaqS+TWSJEKysnh/J8QpJFbb0HmgI
0Ul4XcVSvwAZGeic+qdAZdF5LVQMp+/VQNyFKPOs30Y8GLNOms5T2/v+u8MOy7bK
P8sQrMP/P8CoE+xGjDa1FNzcxK3Uhr15N3diNlLXqfLwusFnGD9dgW6QJHxN4Td5
3W9LRngIlUmochbDSzRmff+3t8dD4FkPaTtTquoWF6mTbpIyLmWpxh88/c5hJSMB
b8wQAUjj7B27d2gIGYKnN19wyiKSDcFiRwnCsOjWsLiL6Tfa8LcyMmrXt1cwbe8S
CqIxKLuOoFMgbUOofV7wWLxcyH/Zsdkwm2IY9wr03MgWq0R2b6blbdWSqgyaLYCe
XRFmnHONNb8wWY2fDGeLT4AYfBhRzuw1IThMw4nsrhUtOhCVvwy/NC71nJMbgf+P
sqQgI/DcmOVxybCQ4Apj70PevkpB4Hz3e50jiQGuEXJ9i/WM4SsIkhtpu11dvUTI
hG/c8J8u0MWii+NCdKZtCOQbT2iJegL6Ukb4YR3IcLn7kASHzX94DqwjN1f7rrLz
4AsjqVTRuYeaaUMgF3+TOF9OWtWsAnQc0XTwC2N6w1a+yjo3LwU+IuyKIRdYdW5Q
5nRlntFesb317DSvK/pv5I7xjzeSAUUvGe9IuzJdcsxYP11HsgOE1Kn9ZjqxxBbq
6mNDAlPmkMqp0cR0oKGoUOy1/ns8yyhID7UXXUNy2FQlbovXs95FFj/Se6I+0wI2
K0Iv/Ucgl+sF+NN2L2jHf5h/WoZf7TDFCsmcgTTT7I42N3R/GIpXJT8wQv29+CNF
cMZgAHJLoqlGA14QnRK0vbCrYrShHbQHNUo0uFGuz0/HbHDfhpBd6+OWa0px1CO3
MaYTc16jhhTn6JzbynjFcBz69crR/oyEa3vKrQ2OpaOehIG/7vkcu0XCROWvDfEj
5VZGutb+yamFT/XIVxVD2ppSeMwQypMYGm0Fix0Sh31PxNyVZ04ypXaWM/o3XjOB
3/fudcmkkBBON/WgObEPGri+xCmewDCpwNWsLmoE1Hhd5DrosvzkABoFJCor3Xgj
L2LEaw/H6BCCEHWNTleknVaGTnvybUV+lVX69aq9t/yi31BzYbYOG+383FBHVrbK
zrD9vRyW3tHXYZh+y89UF5uKJgxPgp/NLnDbUpr7lyvsp664fFHRxp2ETTTyyBdg
d20lEkBHJDVAGbov5Ufcuv7nSYAF3Bw0T4EDyLjmB8GywAKyRF0Os+dHtQfBg1Fm
HdjpObMSE0k/7DfVtDW/d8T7FEiAniFCeHUrvkSSG8UZS6sNQ2X3fEhToyhaNSbI
/4+EPxnLLOqethhK2i0/yCEtm+a9Aau0amvh160XwWVvq5QvxHinmup6HoruQWZe
Wl3pxX6+W/IkVWd4ONmMyiA44YKkD4c+SmFZA1kWMHRU2RU9qedpSRgfKD01lfa/
FFy0hTy8ARC1Md42wvVYBe26mtCRYOHubeNqbNrjiUZwGHmQilm/b4ITGgzm+TCf
swOb1w0sbCFTkI/BZPaeV6C2ULWFj0MGOMq9T/+Tn3jFrqWnRFVVS+f8vb4auPLu
dYavK7b7zXDMApggZkykR00Jvhu17Vi6wS37FKw5oUCEBh/FhCb5Sk0a9pgEjsOx
6qW36K5KzAETJcp1pkEIzl2b7WKxyHXBLOQqsrJToUFyFtC5EvUooc9K6m+mihY0
H+hKNOWmPW8hsD6ULLF+IbXgEvar2SHa4mtwaNgraezZo9ZM56lMJ1pyqjTm/FT/
l2bysxFJBcAybeXS9zP9HcRgaTMIKGShICibMfh0ieB6T7sxm8JxFTuaua0KRdCq
CTyEh4HEdqIE6sGaAQoUKYos0FTenNaZ8jJzJkv9EVFhdDtwwrpqmOJXAtmATB5c
/pTJOywZv3dc4dLjmvzyaSOxOFDPRsPg3qig8z6jY3wqoUPeoqyyi1OXhTE2Jqdz
b3q4fYEzM65P3jQT0oLMAhLUgNG9HNQmuz6Zo6KwJgA8n2QGEkZN3UUcBUzvCWZd
tllGDYdarGbQpihFfw5IWOTNjKd4N1LX4FVBYdUR1SX1MUsjPbJMOenjII/dnug4
62NMSvD/5QxU2fKhR7KquwQq+Iafevn2mRS+lZUlngW3wKULItBOarb8x7x6n//h
esU09DPi/ovF6hx6hbqygBQ3/GCYO93XRi+asbjcTN5J4vXasuS2DkPFD7gpYi+3
1bbDK0uROJf27rYK+MLPCK+0TNPMiuBPKllFyfyTFYsXQPJPJ9bM6nJlhyQg/c9z
ddLya6muuuj5Vpy/4600MQxNUdff6wkhKWrNQLGUw/uLpFogHeKJAx+fnQKdGvZ3
i333iCOodeN9YVzM+4q5il/C+RtKH7qbz62V5Fs8CnoOuXe7NiHzDHX/Rf2xExhT
MA6gJwZYD0h2wau+XBfBF7n7P07uWMzOh+8AdlBcQQ5feBrKT2W4CtkYqBarsVxL
Y+v0dQreNxTULtrctnVNd6C20MqnE6mRBVvRyAnNiZAzDxem6HKFPPSz34zX7wR9
UK3Kl+kgP9mMnktBz2gSekh0XibT/sJrymmD55xVBqtoaiXjZGVXura+TLIg80EA
69ei73clRlPnJJkjxHVv3Smu3watBanQsHvo/7CELrk5X+pmlaylBd5SRUHTWs6Z
Gs13sptkedIk1su9ZOJENsEOAnErrfTd+zYp31gZafp65wWVaVxFX3YmByHEaWLX
Ns5Y4dfdEYrFcuYxcjUbIQcqJYJzJL4wiEiIi0lzPz4MD0Of1Ygkr/AX1QWa6IU1
kpq89wLEmcowCHBQYooNXELbjxrA/DX4gh/7bhtCmEMH6XTIwslYRL9ilJLnSOuu
wdB4+LdUmBQb1h8OSGVGpQL6fEcNJGrh7IBKhRQ63gV4GmemYnV2+fmhNXwh+8uX
79YUwGB0mNez7VPS89v0OUQb9PIv+Jva6LCkPyHRe3g1jMMAZvFSch2bBCuhbXQE
Dn84xyjwzgVQxAgk5H5dL4WbjDYXM338cxc6Bv8P7idjRRNH4+kTsEr/zWtreQ6g
PSv76dh48dL79ZNqT4TWjN97fQMkmimz4Xl9aHHso3IOcdSxgrUSvJ4CQYC5ggJv
yYJataG6iJ9I8qNe3Z5lfv9xN0FYEHXYfBQOj9njWSlO7nqe9ghAnfcXLABYlhHY
7Zx6YzmJh5SAXVpWhNTvrj4vFnJzsAgUCtU5piVRLZSjemws8I+InRd04w9MxJO0
atE1aaGynIS+Gn/Qa16FqI+xfn06nWQ2atCMjzAs1Lj3t97PLobx6NH63eScdUx2
z+DJUs5WegBfkxIMMNcEj/u8A3cLwFvQ/jrunATEd9ICqIX999/68fYiMDS7+jm1
ilVpBgLkw36dFPQHWPWHM4wOaJmM8Q0dHeQ3p+9W5GR/ijhn+U5OMqC+UMTpsqtS
qQ644czBC7IkS+AAkzEwrUKGWJbg54aZ5BMvcKkUKYWvPlNEa8R49QgP32xM/Bwx
28i9qJiuIghcOL2UYBxcg3aOpD3obR7pTNbVPF6KY/oOhVOkTBNv8riM2FUIfyXE
hgBY12A5vtF6OY3t+7JbkmiuJnccNmqbsDwSoVGTcZxoZBz5pEVZ9k1TYm69QJeb
4UXCQNeSQVcOiAHQ8SRpeDi/+fArkPu4kn/gugydb0OB1H+2Q44icKOIFHLq0UJ5
sd3C51xCO7+gN2/+o3Waahpham9CTJZU1Kucm1iJGd9z9Jh5ZDHJ3MBt+L7w7UcN
5N+Yz7WZ6sWWCdw/kjqp9pWbJzFrwVgvYJXgrFQUY3UXwsGRHwcTzBFvbYjgjADe
yavV+7Yeyersd/wWoJpvUw+QIH0fQI7ChdIJRUZp5mpXMHUBC5RbC1QM3tMsOhMJ
VNquQEBiWcZ7Pfbbz5lXcyVipgez7jAdOJZ6hNDm8sPWn7lSBhZ9X7YpQopnR9jW
YM8W8NP+8GQjreT/JNLbT83zvToeRJSNWMc1ATzcIQTB++jcSP+6mCxEzUY39dvO
bm9tzXsjXEGGhdjNrJm6Vd0FofTygAYSIfWWGY+hvo/43tQZu50CTYlvScfuERG1
EHsCOYeXYC/FV5EBXPftZ5uA8bNUmIA66VI9W66oYQiHBp83BLyeKHqQXtwpjJ50
uxq7642iIWzfq9cNA4b2a2xNtEZWZfh3OqTphlidRVdOV3ZLpqcVUysYRYwi9FyM
NQn5QZjktx+jZnR7SISRn8IgFRp/ylH/FGOCQiZ3Kj/1pbPPdjQmEetiQKKlrnnT
8MJbiiXYJcb9JDdN0dgsUcg5KmnXbGVY3v5S7M4B0z6eLtLkCasV1LDVuLQ0U/nD
MdypUbBFQV7sQS2eZ0eXfAUk2CoKbUR0hreg0VqAXZDqOhBioAifN05LpoNHTbPk
DPZMhbfexw5W60CbQ9HGPX5934JW1XR2NY20RDKrqQscbNjOS7a81F869Ap11AyF
IAZXlTWGwKlNkswo96wnpJnG86jG/CURYRWAxoGWelrFtzwHU5wxcaUPRErrF/h5
l/AaWQiEeDRzaodCOz7/JVHrm2alhQ7yAQ5TjOG26haJXhHt1rRmsiy6qbRNS8sn
rz2RgRKcK8PYQbxG/koIsvvvdF7Lw0bC+QAuPfJYlG+zF/hsn/HdEMhSCJ7qFLuu
KriG+bONlGJlNUQijC7111HjU8povB4w2belFTCXPs0xcKFKi+bZH2gL1ZrCCNCO
+wj2VcIVeVyz72d2V6jStOj6IZGDWOgJJ63F4AquPnqT45U3ROCSIKJl2Kt0yxGM
rTFL0L8D3Y+wpqMEy/MkjaGhxUR0+Ftjou3GMMrlyEOpyXghwlxB32HxKsInX6+a
5cJbqcnq/7r1WnYW5SSpIrDsdA5zkKYVWkee4WZBOqrzqJ127rJvgtQmD8rtoE5S
yZ+GAKpyyORD+iGpAi52qGwIVTSqwdPp+Xz2A06zqFAejZepWo0Amxj3J9S/Dk5w
Dtas0VHSKrJsfq617h0A/XwRt5HyRqdigyO5EF5ptW471V3nR5notAChJUgrZA8e
hYRtTE73NvqM1vRijkth2+321TB0TSy39vgFZ/Gb4kBifw0kKYRnViteroynM7+N
Y/QTmTv0jkCQeb7Fv/dXypeZYXHDrFSafGF9qBVkwoKD1qW7sNKy53g0dFCMG/nF
jdh/sHHjfWgWQXz4q60ANaXdUl2w81ua+CtyIehXFLlNRlb9+hsHWASP/gftWDBl
+7INUSdjBUxeSVtXmismP4XCgjnkt6xRWCC5nhW8kRYvLSRWfRJptQ2HqH+72ddJ
Brhnm6yLIoGxzOIxHssEfGsCVB0+9QO1auTUdEsIRT381UVHBHQaAEKmdDkhpoSi
Lwe7cQxudWaRJYIfbgblsO2vQnHwcOIFVItIP486OE5g4yGgst6bsdptS/Cgy3dP
HJiIyQV/grLgyoM9skNBjyADYHOzdgHQILvr9nRiRZkVNu5NA6osV+rX4GfjtZ3N
bxcAcsQNusKYOi7oLpwbFcxMny7tZBA4fKkeRGYSyr/Z+0skqVEYMOMWO3wlPj3R
ect5Ska62Tc2SxLyV4K8zPQNg7fuAxrOfM5T/B375C9+EtEt92NzH1yvv46Q+BA2
7HVR8xCR5DOrasjdf9imdm+ArgF5lyq2ZMEoypg6zKHhBdJ/jgw88dyVAwiombFw
4p2l5Suhpns3KcJLcG1vajM+k76s5wtyuJGehshYU417/JzCnVUqK4GLwCK0H/HB
SmtftXtb8qXuOMNjq3XiM37q5LNWskbl62SbwlOKHbmBlbxa5EgBPO6XS28qfU5D
h3mFoMYs9/6DakMxMVAiU76QyUgqWLpNS+wLmvf93NxjhjJnxatzkV/BnZIuYQA9
nvoi/R2+Wo7mK3vnz1gZXYO+IQhhjjo/5y37NQjcWJZUCJAIn7SmdD1PN+TOwHtl
/dXTELeaCtyfCvYjXDGPEbAbrlPu3XUB1h+Uvcq4cFViCLu5iHNa90g1YNbNT40n
2pYxombNQ5FtBLtAmAoJBDgP3pZRPyIKRGx/lg+rbZ3eIiXFs2GJSOxxzJ5RIuLD
V6YFauO/t3ysOBPZZs4MvvasCV7xr76ExMk448G/YCnUPzvPXDMiDbuM8uCrcvyL
9jBn1xjP3cuUxWI652s6SmStdG6urqaWHXNpLSqChBWzMT1TvBgC0lLFHff97X24
loGoAcyL0RCvezIIwIo82iadUL+8n+orp3UNRa5kHYnCdrkLwvY8TAiFWkhg/Y4F
T6c+rYIjqspRTNvNEjHLZ/L+RR8Wey+A9R/GvrMAxfdlpz6OvTcxuT8Ox1y6sCSL
WVQnC2KC/lzH+LnOe46NjhNF1LRSoM04/gS+EThjItRgbZ0qjTLolNWmiqvCdPrY
QG0YeO/toimLKrnpaf4leizi995PudpiHSGqn9NcRu+bnDt0PexGe2fCyLE4s875
hlLIdGXgaXi420O8lPJ7gYIOhHK1evRUjJqVqahKdisAh0Wwb8KOgQw+VPcEOIJk
9IthsftXRk7nbm6oUwCUIVz92vmIcojJoyCSXZ1QrV+D37ONhPB99RIIh+X7PKPR
sx6gADofeD2PLLVXb1CdBDcWvKmvz++PE6aSJhFEYGk1TSElCAB/HCRzjT20zAKh
JE+hfGcG6Q9i7TQhY5qVF99sgu8rw8JfMMUSdEUo60+NuhvyWOzWkFjwK3psngme
kCFIq7riSfICM6jDgn7i6bAMzDlSPA9/IF/ILO0gMDuVoFnMjejn4VlvjEo2dKQg
dXAGOUvB8djFjY7Tl9uKZspehs2p1t/d90wxH1TMPV521Xs+ypSZFmWSL3NcB3Z6
bNDWGU8rvVbUvQZ3pzNgdJm/tttoCBe3GyKrVBnQqbyphcE3pw/WZuIQJ/9wapCl
FBeWAvwDzz3ATb8BLTkHSjimlVCRibH/gjCLrIHz2mXrb5EgZUcTDeLU4TlqIAcw
PeF2vAXQL47pO5B8a6Q2HbExd7CnMrEO8eomgniIAtdHSUDw+Wl3uOKG6ysIE30e
UE6+aCY3rnOQNGUKFPtocj13l9qgjp8pYgRf1sXJYM8lL1GfvU4i8WozFu06JN61
StFeg6AzDLb73IH3QY+YwGvX/3Uy5hjmHVc+GsFAzXsmu87nmDefUz4OIx93IBGp
P9Kc44OOH1Ej8oJrkij2UzZFQD68fOsHQ0ocgYFwKDUDabBE7JbuupzXmq53v2H7
/fEh7MevxV41//Z6zHsXyMhISe/EOx2Urpl096wifN3+0X7Y5T2J4UtzCRzr1Tge
LLqtvOALmXS/qz9eofSnBYbOcr/DaE18gHoPhhVJlbXY9lA8jO1M95vTdv8KgJLM
WwL0XqoX7PyLP7uri2ukicj1sksuG2tp0iLPXfV9NcWz2paC9MKIDsqBCp3A9TdZ
B+bPFPjHDL88UK0EX/+ygrC4rvzszLVzN/XzquFtr3P/1/ohxJubbq4SBoJ0dMcx
F3xwO2camzATIKqpHQ5yKEDwo+3WfhYe70kqG6QdLpbPWXp9tSTQQDXlwcbUpyMG
AvGo3eo4rOpud9Ph89cKEZ2QwPESaZaOgiXiaCKilF5+hM7VEJnnizke1bklrxDZ
YMAgY1pWHY9VGfNZhem7R98iqJ/TUgc5n+l6187pEjsKIrf0euKKHdnUYg1NU6IO
IljTQvWq9UZa/lJjgfkrKsU2+y7Sok0cs55QkHa37Hqfip6/5Kv1RzTkV8OukgaO
Smrl7o3JGHViGitNpFhw7hwSfLrnakNq4YSeeauOxcyKr/AzOmEFBz/d0Pmu9owO
l+SjVmdnYARQfrrul9g7WocVq4cswJ+cPfMjL8Bb9cuUyiF2bXsObtRkL/HUynuB
0PbmjI72QgmYBr2Dn+aYZKC1hCDxYP4bJnsuWQgk9oQkpdDUM4B4ah07XDCxcQKQ
Q5rTCXt1qSsZ1s/YTkOWI4V+aJyMMQ0W2oDIrJJEn1ntXdr3zeF4utVTbBBi8V0x
UTweLyVnXpCiicnc8Z9s5lThiPxY2dPdpJBGdS3pUnxdTQUkCpt2dl0qWl4XItyO
kF3my0lQtt43knRyNbeYsWIvLQ1ammtOI9AvVyA+lOSWwdQxqiZY/NF1qNbMpkwW
C7R5mkcXPaqkcoUUXZCwE1Lg3LNwWY29dXNzNG9FEMQr56Jk3hI8aI3saV13GVLR
2/WSXA/Y+wwVxvvmKHYDBXytlpl5QmiJZmEOeM1nbsClbmYjuUe9WD89cOfOu6BA
CeZ+NcEm4f3VfLeu3j/Jb3PI/44x15BrI0c+LtbI2Dih6HbUYhqqXfitMI2SRs63
P8gdS1SeQg++j+1+VhBcgyjxlsP7pWYLD1mAP56VBq5qJghGe1m4aurFUD/el4lx
eA9jE+X1oXA77x81eWQF0UaPa265K8lTg1P6Dtacb06cAK1d8Le0wydUliBRYs1V
bXcx7su7d+qn5snw6IY2eVxWJTku+v8Gobdnqd37DrBjUJGHM5rQfnf37Lm80+sh
i4zNPQCE49LtQ5jODBgew+ym6S/7/qPzK+WEF3sPrOJThuAigg499qgiB+7CzVbC
qioZ6d5T3Twi5I00aexzdnR/08UN5IqFHSwk/N2Cb5HvwbHPcFD+acCDHMyfui5K
vpjplWfIfTeyT1+Ea2B+BZCSDE71GN+rMLGhUVc19DBsvlIsoOqWiuUfpBTYb/FT
L7sQXriDoZZjZfiBkPK6KP21J0lgFTHj5EfMc2J3zs3n3XUhj8Ex39Yw5T/cG8Ed
NM+jkOl2sC0/LLr5jdBv+4u+2BZ7yXT1P2ivPwJLZGEkdBvW/yyeeqljbPyCGFBz
3FMY9MwzYLfE+iKpgJTcWvmdq+Szgyh4UyQw44B3JtKr7tZxlbHPgvRIh2QNuh35
BVVfjHM80QybgAjFDvWy109wn4x40ch2BRiD5g8sT6obZzO6mRVah2iRiMmJf+LA
Qj9WXs6Lg2ZUly5dv5p35erjUNrrN06Iw8sWOo4lihMonL+V2Qs/1uvqfadQNPhr
/KmRcb/0WUU2QH0NhHEgfBank08BCGxSmNOM9DHfuddNb/sXuVSWGbc5J79Yn+9L
jujsTzOfLmlL+D7DR/J6FeeACa3JrZ+ZEmXZ2AXmBf0TfQ5ONCg3UJabHraYQ2vj
DMZxg9YelrpiZZEkLLruqrZ7qGjGV/BTOfqQIU51SiXyy2pkA2b5D/OY+do5Y700
AucW8dz0dD8P+Qbg/BOjzyprzj+iZMEOW9zWU6SSaFClwm9SQWO0D5Z2PJf1p76g
EX/jvaKI4e75t1SJc5nNOFg5y8xQeEMUwQhXOZL5umIt55mZaF6pe/wFKDJoRmyw
2gOhjmKHkUXoBL4y2ewDbt6LjtAkeAAbTGMUv1hctPD9tvyDrjmGErlDQouh94fR
TAsh12rx0ctz7zfWvNPghIvglJv1Ow3NP0U+3gQTXxLkApmeYpO8vtBEbcQdwptm
HXyQ7LXh6Inzpv48x1Q6Kn6Fmv33uKxnRARwt32uELZYWVqhf3f3omPOBBbDik5W
NYOwcpUivPqKb3zIWh5n+7Ul6HyR1Y4v4JIbb8XNYOftdr8jJrI/Jn1R1Cii5+VP
lnwNKqMiJXbqamR5+ClRRR4DwnIg7frlnRMCV0EXamqYvT3D64e3BkB1EqjxPxBu
AGTcrQEib9yqUOkrsOiBpVqSVGwiafYI1m1a3GYCCT6osVxqHl3TR9j24PxoIbn+
w8X5oNJ7u/CnFu1WKzOM7CxB0YFkUdlCYFQEQd/PjmgPiILbfwGR+7fxXnPIZOPy
qud5uzr/loqevZNOwPNGKUeZmngDZtBni4uXhdfxFg00TiWJ79xCH+G9NMmzczyc
UQLbyLp6jYdCHNX3UMlGu1M1/25DF+OFpdtteNEyOvQa3cxR3y5UZoVuI+a+5hVM
ikE3FkbKg2DmisD1J5bORpkaaYBaE0jJUKpjLMB+c9R37iSHYji4kH/mr0UVL+Ba
vYpQ7nmYMOM7aJuhFWaKpMIrY6eYKlpWloMvA0ClHa4rKHaAvzu9yf7g8QBaxcpb
UJLFr+2tWjQGzI6eQtOJI4uS65RGOm9sYgMonUrPqvWhtYtQ2oqJ5LU3Q3om/LBq
cgj8Aexw/xYKXXyvHuyqCrR+0TO14nl67zDgAYpdT6f7DObhfszcUr2+os0R28vO
6gKZ/LNhFp8ip2QcQi0oiwTISudHs7YwVZKBX6Z5KANMUlyBMR0d7Bc9MDDLfLaA
U+P8y10jsdXw8pl3RguF2POsjMC0v2EDyAdtfyRF3dZbnH5nEFKGYUYZzEIYLk1x
/xoQjZn8+lbvAbPdkt/Fm0zHIVNKXPNjosSu+QBgsxIbk8EVZ3XAiGvaJ237nBe0
jKva/iOl8vMMy8snN+P02Oa11296WTi51A2EySki0Vm3CrtYwFk8V/US13KPYuwS
6LUoDZvmAmv5vJVIsW9HGrMwlJJtDFj0OfuM+1yTBTrBSdanysLbq30AGDvNZK5S
QpbIqJlrUqRQdkEWK74/Xz/9KgSnfzDAyixmhsAsOBKs5Byr21CdBiUsJ3n57qf8
Ms7ZpEe1iTBQRsvOkRjqD9jOFDrgimOCNzNbblHPQPpA6eChC6t5lHlEKEvM661G
gPb7Bz7LfLunZuT4YiQeBnGVd5Xycg9Tf8fCF+72DVKHpxCZ+bn9z9CVb5hhvKuT
AKJlewApBvpWp6lwniEkJ8SdSb08GA/HiwzGGqMcRtNWKHt6UOVm5SMw3700taFt
OVknPR4GewtPJEF16Z0XDNZbsXdZK7BN2NZKSNwXkG8o6fhb1dvxmTTK+heKJKzx
YSxP4uootw4lwa4pXvULikFbRYLkIN8HGrNWX0DZezsdB+kZxOG4ixFsttJWfT2T
9KRRGevB5NIdeS9sS1NQwIcY7spJxierDAHyCLHxtotAt+Qzv7OxqLzCgRMunBbP
C12PqXorNydGHWKx7aJdNmcvGejy2/Z/dnhNCXuzlaihm1pNzFUC2X0mNSzJjdyQ
cNhgX7QJ1YotZZmbUIp7facRhDc2jHn8/DChBh2Whnzak+sKNY+MOCu/gI+cnQHI
TYLuGGw27sMrD7QFpYuEbIN5E8w5TJZ58OrI+VJocMFGUGcyXLzMNVWyoovGNL58
OIwCUXHpg1zw/5I94gwmCwUmu1gckm5Z5RieMWpJN/sWA9IB/SnciE+GlwyQleJ/
aDNv2d6fKx8x+rXd2rI+zWhnnvogy4RFahM6Kwy1o5yl11QZJydhMyP+Il4ZTW/p
VtBfBZBQZpJXwAgcuA2LLQ2wAtixHxxm77uA5VFH+23wJw15SkKzPPcwUyz1lp8k
rlR3edpmyaojyvtsxajWUvDb4HAfNzN/KMK5qnAfR8RFT7JvDMg6s7KEVzkJSxYq
7kZpKpI1J0HUuvxK/gocH0BuUTon5M8F7N/zkkUjYBLHc1e8yU+1IQuAt1waURB8
4XoBfsLd4+LvYfytGDd5VQqK2TLMixANvGZyDT8T7Fb/VCTglok3DQJ1O7CtEabS
G3jiO4h4jyS3mf+QTwJe38Uy0cXn54vPZzVGI1yAZ+Bs600ufgJy7Oj18Q3rrLdB
tE3ERqRUo06cbdwRX/k9PlwjsW0fwBUdzASdWD9+1IqCtZ53MrfUl/c6slqwoPpx
CZpLTFXsI2qQnPlyPM5rQOAbGS5Kd/RKdfmVD5hzjLrxnDvogpq1OC3YaFeeU5be
UxGD0OSkT94J79AFHoQ1D3n4SdV49T9k7FlD6bSeENzRMVH9HcThJaTMsTPMUQi3
K3TnIwHYoAtzaKQkGrRzB+B8tYPIvWgcVJnUio0lHjsmaG+4M/q8VmgSxpCBVQpI
4FVtTfcAB/3taQ6+BYxoqhMovl+qB70c4MjrSGMRqrHxuAuZwXBYMk539iFm/+QS
GwlF/3w8dFpOOCNUzm4YvBSIh3KH0HEtfRdqKCguuAjmtsN2LcBqDJMJNia408na
vuU6Z1XY0nBfcwOdc7oB1H1/vffmBxVhfMohovIbZMCOwguClNJaPsmbPuYnI4xk
DnuLT43Lscq08CUgUKFEKRrKaKn4pfkRckR0Y4NW0+6xvy1zOSmUFT8STSv+rSq/
wonb1DEvJCuw9bAEvbYSe/ZkQFjmT8LpfVDof3QNK46e1f8Vn+Xde0ySfJyN6nrn
Igen9crSaPVg/uQ3n0Rw3x3LgSpb/VPP8zBrWm51RPIqqH5sCDjM3kCMsxUihLfp
V9nb6dgxwdinoGjuBbLEj01FpArsxf+X1yb0pn2d0p6QE4Y2jPAexcGxUZ8GRxxL
9bqibvqEsfeITVAkUMJ9ix3m1QBHrEnfVv5hZGyfdK5eN+3ghL164UE6Yihp7cjJ
lfIklnsUDKLjlGZQT2ssKxoRqrRrJXIOWbZx+g5Ci0LLNDfMg8arg4OoI7NVCbSY
A23yU8U9KhQShOx0ILD0k4K/gmesbcDqJPTZTATj2bydDn0w777wnmQRLx6aYL+c
p/DXOkGaFyV9Yqz6eFLXkYYKaU8xP4TCc2WXoq6ELXOMHBdMz04dodLH2wi3HVqT
WoPFQcfKqoGyTaikHyf8wIZD+9Y0wnALr0YgRBq/kXvwH6NYoZzUid+20MZwtlzw
4g8666FY7eyiUwyBkPxOT6Nv0o0UYk8p9FcVYq/Q9WFLN94EW5WxBGi2NW8U4drH
pzMN7qvaEzMrZv4MpQ1uEL4yzw5EQWLS1qba8hPOh3tO7Dr6dB6jzuCXc9Qz1CcA
3R7dUCqUBserSsIR/DnU9qMBCSi6LeGufoER64Ke5j25cG72kIxWnqBE+bKn8XwP
6D1teM6kOJRNlXbXsvmk5qpOyTvYZuwtKotnnvJm6FtkxTUYESXSycbKQkcBfmUf
AMqqooMIskHg2se01+EaavF3XxcL+yG8RtHslh2+wBT8N2aSnA+7msL87KzpqG7w
oHMv/eKOm/IKTVJ7/MU/dXp3PVYqRF8iwrKmpxTB7SQeWWlck7Tlvy8kiNFPp5jQ
WEMAM2t0Mxr6HadJTzL/psLjoF8rHoPE4eTlSygSS/7m20wHoe9kZnefeHAbIpY8
bsPy0uBrCZMpxqSkLpDYkP69MGdNNXtb0smICC1HjA1QUKem1fD38OQkqsxxC9W/
0DlDcRp6yEl34GrfbxY07lb3sfc6omPs6bd50dB9xIILUZWJOP7OwAjqpkPRWb0y
SFs2PlFFXSU3Cz96C0hdjLLCiURDx76ZyaWGFOo+GK9J367TW4wLdUGqTIKeuY56
6c5YIYmiJVvfA3WZIs15QzrY9mlLhOobLpqqleqt1yU5kmLrMHCZmEbThQCQMdBK
k7d8LxrglyttF/hcnF5Q0xU62JtLI5EKr6/ISw6LQGqMAvPTezCZPkCRSoBkjkgo
GVal2QOtn5OSsCSgxY4FfKDzsaX3OQFrBPvVZaczoZOxiDDpYetp3Pn15du90bFs
HaF+6xDhqQ8xP56Nnq61TKQ/llcU9JOlwwINJBZHv3oUdSAY9rUIBfNrur8fNuOU
PYqE6i0o6BpvIbMlxNBLm8VgJMS6tc3rhpCuRKIA890va12I3mDjyGfClb5tsG8W
BoP+2NTdgb8PW0eD5l8iSZHfcL7Q0k99eTCF7rAJAMs/1TXTj9VLFui7oeEIcWJp
iK/5E3Z63k1cwKZYi2yhMuYGymVa+qJFpqSdQbZFrjRJ2pBu3Ax3gaxdSqhl9sye
nocKmGR0YQHrxGumiywsL0LViuaRsl+qidwnAvLV0Cem7nysCUTMSo5kQFcTJ3UY
VnbII2RrQ3JeInCDAD46szX1Jj7NCdJf8QE/tUwbmH7lU8hN38P43Zfhea6rHc+l
EcmsJt63S8GcAHaDMn8OFmAQvyX3Rk6hDzzuO6qTnqLjz7BTRhaRPZ84OmgTVrze
x1Tb4torLNsl47kINqb9GqsvRXSaERfMBrDFAo+m4z5955fNvZfVKYD0whxbNznZ
7wp4VKjiMG5/hCXnQwhyZY+1Mh+DiRvLPGJ+a5m1VJZwgjVVKEskCiYKLdqDVjTZ
jsvFzSP6Kxx034QHSyj/suS25LbkkxDLHP9fRpNJalXsQOnAUpdKB9Z7bxJEWjvt
2fi8+PdHi1VX7ZToYq2cGyO+hGSwLdgGjiDR2I7doFmlkZf1Do4asdxzJHw6XYDU
vZVjA8daQfUZL8aHrTZTYsyLWow28+z1uJhu0jIHNTlALauTjFwx6lZ/7R14e7qB
SRs/p4jgkxS0rf+ncxmze9cCNg5YzQKHvQmklLNCg7lhZN5vNcFiupEycEBIUaM4
e5b/lGPA417qcjXkUgk5Oz7B0FcdWo8jSpDVI0Nzxi+c/o0M/YQMtxaCyhz0fCHm
pcESe+N6NNZfwIQzkrQrSq3MK5lXOS66t+14ukBFbTrXDblsGa+Et21g/rgJvRhv
fuVOmt7JKyz3FDscxhZVZRNKKhAhNLY6lr6rHB4CuPRMdjDy6JDboRYYFSZywgWG
RGZXTM0kxpBaoAWptX5FzmQH5DXRfY0h9Tpa/OdZ2MklYau8Q18Q9/EirlG1hGjh
5R9Qtrg5em1cd369qyxcRYovP1GcXZ4iR/t1iY4oqW9SzGg1LIVGFvk0J7DFRVZX
nhggfySBV0eE0vd01ugN3e8piyhLc2If426HNs4Y0lO4hJtOo/8qRRqVmULn0eh3
N85dqAiIBoHdsH5bQQUI1WOpLToU3fzMdgVi5fixIDgJ2S6vmlG+Ssx8PhB+UmYi
atZyPaLbglPrsFmrI3InYceb+6LP/aRJM40/+6yGO888lNc8ssE8y+xd5/DuY3E0
orzfQ+G1d5jpHa8LwfT/sdwplLFZ7cCsAtU2t/7ydDE+V5OuZPtkF9ljA3qVwpnw
sENzWCOMuEvccrr74OH6EIt07FvOeVN9wJvrANFNByi13vCMRr9lPBmUQ2H01vJ7
Fp+tXiujqaUX2r/Ouqdsvdau9Hj/wC8qXx8kTdQ8Y+V+DubQMEJ+G3z2/kXJ1ZXx
UQGRcG41m7NUEqxp47wtK/J9bJkDiWI2oTjIF9UgRYAdNATphlzyk/kFrujcMZxH
yQGpWzS0WxPoiRR8RKs6EMQD1CBCiD8pBG+yKuTgnBDLkUk3Tbv7gKR8gUTzeqok
tu/n/Os3E+jrx/UitJqSgz2GR40KM9b8ZWwzNZ+qjN1JQVsacZ1GAt0wgcKeZN0e
RqE6Z+ye/9+5nOMnaX/9kPyLuRCF1wzPkHmmppYmHK582mCnNuiiC/ECd55JLsG2
1YrP8oQ7/bXiA8Av6MCzYfARx+3SlSpWRUAp6y0RKy3XbhhSp3vETA/rkwkZtScP
ehhVpIdN7UiR++9HKyt6exdTtJoCNY8RbBxt/K4WfxEGWu14cBk6W3R+6pDwnbWo
TLDSL4Cy1QZtKkVuYGYdeiSLzOYB4CJ7kD3prsZHwtg7/ot8OaHMVVIa3psLs+KS
ZXsxKNX06gK2kja+OfvQZBv7zpTvzcjnverkoKa/F19tETHe6X81GRiAnhKSytEN
c/DJzi8+lpLEuJyVO5ImtPcOVEgIhdzOFsKCXjwz8JvRgXg59KVhge2R/pxLyVvo
kSAisws/1mo18N6/nahXIIPl2sFfXRGykWaduPyhuqg2NcpqMAzESnW6lhOqGp/z
a8Ed7XjArs9EX5gQP3tJ+smNHdllTNhAJi0rfOC/CSIZ18Ci/Cjc8RHmbrpWR6jp
ssVu0D4IIKft4LfjUclSNm7ugHre5W1IKCzBy/vFzBWyd2z8luOUHCFhWa4tVKlA
NwLMcHZZ7iSXxBvYC5ufMGi8JwUhUP2pcO0WayvN3Lhk01in0piXGkbB8aNScDux
1QRJbjrjTGAp36EJDncw3PB17L3mTrkpDmfbcnONh6tCwnGB3qWSQyRO/c+FmkWj
/AVde9+7fj3G6qPAiwiCchvFDjHJdSb3DlnXMTvKVxmzq2yuWT0ShCnybsq+hu/J
m+wZa9oHK2M9SfYd9eWsPkwFegTV391ItA8KJFj/+DvafPBP8E+GK5VH3pX2dr9x
TaPtSoOoOG5ZM8Weqx6tx9Cp5l45kHgSH4NCy8ZTb9nmVVKDZExvjPhXhHOMSScD
NcwbYk8pbkqFE9HMd9RTPCEgOORtvuJA3FL6zty1UA9831t6APHW+wa9OItmJc51
U/XVltf0ZxpsZYGdI7C7MtkValRKHVpII4qTVKNLWsP6ktoVGKQP++ZkGhZgHxpq
Sb4V8btHXExQbtytXFE6aCRAxQKiQklUPMq/4r4wcqXWldk5j0TmI3ae40WC66VY
QLIqd5ftWH6CSNboPsTErv4f0IGWx5i3mySXmcc53hIZfKWtNlhUzW5HWBbnY8Mm
LlWZHVb7/PqkP578K5porWyZCMwwcL3G8bw05OBlciBPa9xLgt/WJmDol/Z/2yXp
kJoO4a1iVIQnPxPrXo9U1A+3KChrLnLLc0Zy8xWptY+jzN7IRIOmAyRvQhIhe5qE
YPqvcG7q5JwZU0dxT5t5D25zoUoLGkoQWCRqWFZKwnSSZkzIkgwY+kPcyi1fqbKi
7E+GEhuz9IVZHcwPRTNfHUR1u9Fc6SmoTcn1rw2ui+E4AbTqeRv0ZAGWInCIoq8A
b30gy1yrq1oVAcYTtmFpWtVnxX92rPde8ae5Jay6bGUTM3wqYBQ5OrQGMteKMj3q
RKY6wC6pHpR/QMjQtusf2b5UR8otiGgsx8+n9hB9j1qgTSgg8g5hQAngcPKtXyR+
8B2UTEkaMewAEPhLv5xnmmI4H8ANRASO0shB8ZVkp+yCCH60orKEBCoOW4nxjqIp
7F0Sy/hdoKdK7AksYkDM8gOu4vfhlJtoCRd4MTjtdX4//obi+inCOdE1ip714MwV
6OvhxjZzxHeoD3DRTilTUebGJztuOGT+GW5wF1c8829p7aDY3SxZkOkAdlFxmuom
k11XU/5DDyjmqgBs9cRMVhiwwN2wKQHJHf9+2CVTI3hREKdAAx6YQPA//ZaoORW2
qZoT8XaCLPGkqnfgz+dARDzPO2T5o+PjKTGC8ZKyDuTepKYWIzBMz/zRYLph5SbE
q5ml3XCfG2YIKYZtTBkMzeWObPwmi0A/tgcVuia1VYw3dPlkunOeMRj9sjBK2qlS
SEsgR01Vlsh3nNSWzAnYjawuER+lgyMfHuD2dpU2wJsMfYYFarNoQr/5GxWcRFNP
62oyYiDdUMb7+8Ry4rbdzjk+9Bqb/TttbCYSWgOLkX09/V1LOvmqtgrJwsbQnO7S
yyhYduip6F7JOVT43jGmlWrL17D3k44FRXgKVsdYWiP1DO0W+mB30oJoTVl+9BHi
DvQjT/6BzOJsbQ/zjTgwJqYkL4kDplxIE7cocjIoPENcOM1zrrHsuXKcx9kJlbHd
+TEMtDw21mTUca1Chr4dSfKdBdgSLclCOg4rYy/f8GOB73tdpUZWs2Jg4vwaCFTg
LIQxox5uFY50mUfgp3ckOwiJqgz6v4xB059157d3TDV/EhCRu/m3LScuDjvwQiZP
a2kVeg/GdlfOR80yy24BHYWjGBMPzwePmquywLx6cXRdrDtpeHSpWkJLrTjy+VIa
u3H8Ek7SY34VcPLCt2nNptM/8DMGknFch2/UViIgKYH2wQvoYOylmQPJGno7wM6j
BtGLc6fPg1tf6UZC/tL1XGA46UDQGHxHA7dp/EfVQFeVqy3Q3mvoUEiLOPd3xhgu
A8OOyWmBAiJCx2WMGq92+BD7njXw7Rslet8lAmssKp3RUkuS7sJ/ugnfd0aoSH73
0NxZCPp3h1n4Vd7dV2q+i0qvNFtZB7WJW2BHj0tJ3sfq2knvZyke6idwv64nwYWL
Lyi7jmqD3Na7dD4fJ/RaPhz3oLdd1iy0X8iVIHBk94R9RXz4x4o+4PGJLE275V4K
OTIMgLKto82vp6dw5c/EYVLNGkD8bHL3d2yEQwodRK1Vwlx8k5VcVt26YBtlHBdc
mIXLY7Ggh48SuDlEVYSwGTvUsSUvz6A9yQ6hA0xv2ax36xLiuLN1iszQicPQGxSQ
OC5czITDTxhaKLaCWKofYZRtqK8eQmXZ30SwgNoGlvgxBjQ3PRJlNICt9qBYBzrv
wbKnxnEYHMiK+slHZ3fbDXMda64ixWoDd4EXgOe5eDVBat5C5pwhfLMTVbBv7dTF
hGUBIT6CkXNl7JqNEI6tLxVZjk/WQNkgZDRw/LJgj4Hi/Zw92vKXYjE8XeH3Le7p
ghBTtqB+EyxwV7Jwig+2N8ct9Jui5MdHJBTKVEOTpTgqV6VYB6AOvQ/Dh35N0Iiz
AxVk9wYoTSlb9sp84tzyAD7AENVjh90DVywUAMZkY+Dm4jjzTj5X5rTauE+eb2uy
L2tV2IhCN26cl5LGXw/B+9IGEnWzaN38Ba/TZRDWOZ3hWRbAbHEYKEb7BIFrkFmH
HzcRODPPTE8w1uGueENJCJIohMQRMMrJpHxHQoPFNYWDXC2flRH2/72AjGB6jWSX
E57avf243dKzqct7ky01QUJNybTpsYrLQq/KDtOqByqE2sdmVDlMurUUKg5R/uOE
Rlb1MAezo3Ag9qKP6czBhN2tNWtd/+bX9CwboZs9BBtRaC2+kCek7rH8sJgjOxXj
XX0bVhQ2siDp2yXYKRNpLDZHAdytSA7sOoCfaCFJrWa/SWhjLRqMVgA1Itr8ePJs
YhkMyqqONtJSyMPaCkcnKavWUIo43lPqOj6V5J09Ah4keMdl1DdLTkbNNBmGTEpH
ISGWkFVsEIccgr+2TuR7UCrC1OATczwemZoiV9fLmwd8/BqAkD+W1u73k5r3KeLL
aTbXGLWszXXPX1rQUMbAY9bIOFAU8C7PGa07ApHEIRRp+ybKNAwlZit32gtIhdcp
v4YuyykKlE3559aSSpIav+2EwJfVoZ/uIgp5I2wwXGXGD/4QoUuTl4MUEyJCl5U0
RoareyTwDrFY5UNsYEtvy2XtqUuka9CD92Do90508cCWcweECJEoBUq1t1PH7cGw
GzKKMfY1X75KPREJdaPrY/qji4Dli39r49a/Uw8pq9Y5IqHqvWSDaibnzLW9jEQg
FYB8WQxLYFR3k+uFk3VnpMoa8YGKBWg0bLZapsSXQtagOri3Dg5IUx+jiOxNtPXo
JsOABODeHHfUxCVKTn96+ZsPgxIwzwdLbjWv9LIP942reFDhr2Qii1uHCFySLmjT
ygVYLorX+QOaagKIYQKS86oZy0OBT76lHBuU0bG/3TkutNus4xRuIzQFZ7s5O6Jf
j/XAJweLnIdjTJdA8Q/+GddueIz3MPbeURf9GLCtS41iYHbOuRPJpjsOM3KZ0Adp
8gGX5ov+HqFPkQ9JD4bAqEK3YVfZzkXGfcvlZEcSVPkMjqqb4aEeui6/A9tiNYpd
6P0nwvX4OB92KmBRiKpljckFZdPDdjRDcHqAyqvJwf4hFiC7K7EITnM8aGgbUU4k
2L6jdROYV77vwO8COwJIy1f4ERyVW822mQQKICDgympy20772huJb5vZxrgitWPe
ym+zKOutbjkDXJ3GGyAuqc0hC9P1y1jixcpJ0VUxrtLh3vuMS8PeCW+f1SpIlb5W
Do5LOp76Eyz5ZIN4lnemdPV5C0lnaE+orUyNDMG5QALM3Z76rb6zPm+YIgY/NIxZ
00jSXrD5zTKVMPZyTz54CO7C8EJ7pr5tSp1gSoxeFQ7ms4bdvzs+7sRI5Vk+r6iu
VKm4wT7KRjN4/7oHtN3DGTwX5AyfCOxRyqtOXLGsXMyiKrjDVMSPr+ygtpo7Hc8t
UlSZ1ttvdhtnlNRwrrSA4mSHoW115LR0UFFrHrtRA9MEZWVq694sOFSrBPoeE2MJ
k/fqSVsLyMshsnv/WaP690YTpQbWLEEr/M6C40wkMaPxeMzUJNRpottMTvlVqHhN
+VegnueYOmit3Li67PWs1z//MEWy8WDMUMNDKrRZweWogzTe/epxtUtWCqPxFrdi
V+C0gshh+GJdLDV9gyjM/hvwUepG830nHl6jiiJgHwb/q/trplh5kFZ0h9bWpOi7
QL7l5LTr2eeUt250o05KBGG+XayEM7qIeebGCxc0jdH/eCZsmsrS3KonGoRYyD+N
J0dtXnCk6N2Qd4H67YnCawwpGog2406jK6edudZ+R35f74m+rlHACFdux/QhR+uK
Fd0ZoWGIRhUlhWszqeZKK8qJk2kkkf/syJBtw21QhL2JCqyA5panhPOtvyuxPOWU
C2kgMUPipnikqJe4xlnF50Ge9CP1Z/OAous/F9eGiPheQpSZvnkhdx1cmREgXn5E
6n4VOQJaE+c1H+ztBATKvtkRtaFNy6Db4oHUOEbg+d5kB/s6lWuZIPAKJWD418dG
wMebmzC/cqgoocVgH4tOTYf1iZPeN+qaQ3VycYyfRsxpuSRU48s5cnEr3kq9KoVA
8r3YrEojxDvgeJsV2DE926kElaNpUdUNvBAGI8Bpi7SyyJdqeXWiULUn6SGEXcfb
1+Omr3t6GkIUB6pF32J6n7hv+5IIiHm+GuXIVrExDqdqDb3uX2Yw1vBvyJeJiGc0
7t8+CDQH6n1KEDT8uqvMAF16Q2afIJAyKSDq8Wem3t22N/oH5YJPt0skG5bl1G20
D2fC5ocZDAECJ6hrnbLlWXYihXrO4AIm7hTcWdCsby4A56jK9FKjIc9uNB0zt1T0
AcMYCKe4QlSSc9vYw5vjYem1+nPWr9jh32/Lxwdf8e9U9S9yfb7Ne0k4kKGyDu7i
gl+4BY+PsWLxER1uR9IPiyi9Osgrky8tXWQFehf40RUsFoFZxBZlImomVt0VEugz
l03FqvCZ9P483enXMMh8KNi46GlakSGQRAqgwAUnipPqA7SpZvY7LpE4eKfF/3kG
jc8itx3IX8OHtQ9c94CxNmliJeEYWveYM5WSmZWpSvu5n5aa0JC15y7vw+XNMpTk
FxRX+wRXiny2jsG01LSEiV/VposHI0wzFnuhgpmHRROaugF3iAE3PQpLBCKxchtc
pSL1sAEcwjnEiFu70mZScyenzDynW3n/WMMo/+4P4nfB40ZeCP0mlz7sjKBPbvVn
lqkjMtTTWpsAp8GPWru1+JIG3LD9R33qID01x15BsXNIFzUFl8DVD3eMnl8jCZal
O9p25jA62ZDIZw7Z9znBVTSINDz4N8lA0g+IsoT4SK9lF43yBXq9b5Uy4TBGkaOo
yLYpPyoqsbPB0AcC7qJeiYn6qUXVXP5RjY0Li1cdkwXBVAEwCugdasIBj4NBMwzb
92/m98KwM4GvnqxCj5F9tL4/zOObgMNSj/EreNxSV6LSBhhdwlaaCZ5iJZ77R9Wp
LxK3GdI9mv+a1Gaqp4k0CJUC+xGbUugLS9B4PmMPmyIbO7eMnSM5mq6TKTxTbt74
9YqOwyowYAH5oAVcDkISIU3AQLzHjiGVbX2G6ojCquRHejCMXAgO3Lf5n7RLO+9m
2H5iYS6SPPgbNJOmaabI+hWT832P8QoBK5fWEPZQB856sf/Upcu/BGa66L2tXDAE
wmvTrkj6rHFYg6VyNGVr68gdmGgIX5og1e1dfCJsUGazuIGvQglslQIs20mc+DBl
Y9ZctZT1u+FEbEw+11WMXc4tiKQABfubkXZz9kr8gzgHBfW77UN+1ZsbJzUV1Jco
jeBq3i1E4m6Jh5cOs67Cdp71gaJj2sl1vnBJZ+C2e8E3YI4NjM8LnEBJ3w35zAbU
4AN9iCHh7yplkepJb38nU+Ns/EYNDrFiJ2gg+/+FAxaYW+1LFIIXP2e43Z+rhZxw
vLiAlrbw4aeI4rrLXyoB9V+toGSw5x1v5L6S6bIF/XPJ8zn6eOir4n0uEBSJMRk4
7jTJvxMbnHhXNFiSlaXCRmctf4ik2ClsQOB+wHfcKhKBJ1evM19CUuqaXFEGtC8P
d3dv2FEPT+SZwIN3+SZ24EPo0ntcgh6HsWE0uWqlPkdw9bVJYFTWwLtpS0hAr3Wp
2UqqWuWlnYLsiq78NHPiB9v1xuNqPIXLYsEO7ve4Cy0IP+MVQbIsfmKmQ32N3k8z
qh5AQXR08RYf4QYRVR9RcvTfklzzoQuqCfgokE2I3kW3sj0lORZA7GOvodtbpCMC
EVW2wpeU8PSWn4yLl0TLJv0J5czmi2+aEPnd3LfMtco46ik/KN+yqlal3KaORtmc
z5srZaMMsSlGHj98EQ7iSIt8PJ/Rdb1WhvSQ1BCOPX08+iKiKh6Cycfd+kBQff+S
vur2gKSsHpp88UtwNR2E2Y/k9n0QoNU7RhSNQ0dskZdYhPUxVQXTQHa936hsdhnm
T08UAS1FGDumFhL4JbqnLVtB9Er+QOlsWuI7CcdRnrtJWAHZr68H5oij1Gf48QJB
yjrfkXJGeZoPR6BEl8wuunFsmNhLKkYwAqHz33wDLQADMHUSfGdZmhiys2epIdBP
CIGQIZUVdqPC+r89v40MGmwoirtOESg9S6VV6Oqh3X/6yLiCx1508mhlrgdUGx6Z
Ov3YMHeRWzFMxSL6IufPMknldannSycMFv7dyxTT+j6At+c5NpIXEI6JmQRqTkID
c7qsXxRCfN664qlJduhVUqU3ULgfiC4CivEB20UghIJOY28x1IWUl4MRQ+mBnBBz
0W9xT1KdFdDLktnamoQwqok1ta84ZZ0sWlD+IFFBBoVBFoUB9R1EeJ4WZyJDPI/C
977GbJmc5N0s+Kt97WkwRgO5uwaIiyRp2pw4IFHqzx8HTFyrkwimM7W3+C8Icymj
zdNWqFDKW0iEYpbH4ayAqvi+Vu9Cj9IVQ3iI1ftFIvvhKOhHZM+pEH2cAwOrICak
2zcF98D4my+yyvtFLqpFcYxd1/I1FX69SlFb31WR+UuVzPLyO4T0d0UXeUplQuQm
f9+RukmhIAUJWHbECRAMdnJch6Ur+Atoicna+pzIED9Nwceih/cJIlGFIvcKp9NO
CC3UjVLJMPS5FcWf8BjtC6My0ep1mzQDu0h+vbva0IEep/Rg4shh3vfwy+1vJDxS
ntAXc30EP+rFt6Ew4NvILeAtAbJDexXQs5db2GfK59WwYeNeKJM16PV4pAE7ZAmP
vQxAGNG8rxkAPK7K902GPcO0i1s966JzLfmpYkdhdweqiLBa4AB94IPT94uiqMu9
ondHpoaYQsu7aeK3mFWyJqhX/uZAZG09DQidIp8gcQRl901cjT7t9rV5/vsscr3C
asrp+RTly6L7uXXjjlCQZrodVzS5PbbvobcW4YbLbBDJ8OTOq8KPYDwK4pd71VYx
cl/r1XqN9DGF42sJKH5ixjZgSEuipQdQM3xUweHchbI/xb5TX7EFCEz8CvlUNnc5
AhGqnfSYJCUmlOAdtn7/fwAViK21369GXNjOH8eA8Ls9lxCRMcJ1qXdSLgmq63SD
4zFTlC5PNadSpdwC7NKnfSxIA9kVgN4jSbnLtrgLQ290mZpR4vHWCXUz+ZSoY3sd
O/ePnC58Ank/8L3hD0mF2eoRGp6ZR67myR8fZp783Td8Fe5YeXFWNwmMdreo7JBe
AbDzoc2zfvcVVN7GdXoLsSe0aPfIEi/CeIm+w1ay/xi89iXYlQsUN+7D5D68Ir9X
6hOjsqPGDdF+RBvPwTrWqd1NzYWFRM3L2ueoD2xar9pIEn/jMokfhVn/APZQVVjV
IyxXAFERM1qqAL+G0nlEbcKtXMBzkZkWmk2yBtRqTxEg3cFtJGj13UWNAkSvLWP8
wfIjfM6GQAQ3UFUp/0InDRrSk5DlZWKN0FKlH0Fw4ff5CRbtkbblQx+17goFpoky
vCD5oH7Es96nw6Q1vQiFS8wLo3IBKD/o86i2spiaPoHqNuq/T0apjnjY4Ujoyajb
jl1VT0XRcBy/P+5V9Qi9absMxFH3jyT1bIMDJmR7d/wNAf3h/toyHRrisF50ribW
GXQ2lecCehE34tenrVn0rJg/1+/c5VTfnNbqTGPBWrD2Qb86MBe8RyTvu4qSt0HK
8G6iK4OOaUPtZaL/+ChJpogoaJV+EuP2fCKUsE+NPBodgsgzoI4oXlS88g3LkygV
K1+Tl7VewpBjPX2gZBtcY8tvNi2OlLqG7yRQYigCBMbl2ggZmUvC6YDJcdLnP2d8
L9gAfygyUJ1CcrsiFg7dXF+oBxcKel+K9RjYEpRzMh6QHA5WwNUSxYEEPOWsKI9r
PcFu3jN/O09p+X6CkRqWCoYaw+jD2Asv6FipvnlbOcN/yjx3kbAtRBgwh2nzuCRk
j6BLyGy269zNhUkgJFjLZSuPr5zxN4SmvNj+bRNTL7o6sSvhsaMR0cOZBfUx3EKg
a6yXw6h57/NIbMlzXKNcH6fhW1RtfVdRj5QxVs374Rd7wlgXfti5YZ1TMwh3OBJu
J8VMeGi3y7p4vYez22sHc9EdwvVWw4GwKu8hmF0ZhcUgVhDwSvy9BzBe0BWyrj/3
xlQ4zl5GCNqgjwglBjUCTHfUJEeV+dmO03EI730x3zx/PwyocZv5EWdnteFe6+Wx
6/LHZ3cdzgg4nioJDB+jNe8V43g65TfVEGypUsMLm/RlvyA3Tc+Uhj80zX+GCnF0
/RzA4Y+tG7GOElsSZVHwzPGbuVmax/VFpRfQmCbjWyDZkt47nCV4Zk6Mg2tQ9w6V
b5z//mvorW3ZPIS+9aSRMEV4qJKhWfXbkCRQpkFhdGNFXtPnuFpdMpzHP/655GY2
ahzVoTxa3Ujuo0yhRw0qG8fMTRWwe2mcY2cegfvoVc+ej7vihf9GiDfkhQLZXjCz
2mwaZ9unRoihz60IoV3yA/c+9RQuLzLToE56MCgEZR39Q/p/UYkl6JPW6cwNxjNl
2KBe23PSsdC94S52xL7zjIKLSd6QO3bRddoTwzpozhucs7R2tBgqH7iX1u7CSJxx
6e1JIbYu1B9J6prK4203qP4cJxnfoFRq5MKGuBv5vkfVjubwc0yT2D77tZ9yrIou
4zIO01pwRMyVhTdACZIFjqpk4mnOLphM/jHkuH6gnvJZVc3aqu1eW9sBlsVRjESz
Fnxmd2RtRW9/GnGy6/kL96TUsOjPLYoGtKFZOOfyBl0etPlD2dwxsSFZTw918txy
hC/JiuXXm7nWQ6j1By0GdJPMdyX65YPYeHL90n5BvbGeSUAd2Ro9ltad+Hb/hTaw
01Z70VKcZLIIy8Yefb7OlQe1KuD7mCBi3YWW9FKexjM/vQ+M0eu3DX9zPjzmkZ8H
p7SsI71QVmQH1SwkDUc4q6npb27knHcf1KD0Jp9AmVNTIeUQfujN3y3LFv3igAw9
c0xqStqKDJlVo6CtT/4keTdQP5ZrR0M742x0wDW699DRh3PfnhrmcQiuin1GpzWj
GdENTm6rtBdnHtPZ9fykBROP9beXePjdYBzvjs161wdHpwfuqOC/iSQGLf5NI9xJ
F65CsIcCAH9EsGRy2GXb7vfJjqBGRRBio493EptI08xnJcdtLHypHqhjZbiGXI0J
LXIi5ifkdsLgsdGfqczh3shIE9SttKq77ENEN2V+1oE/XowLAYAAhsxCQ0eb1O+V
84aw6VYTIsnXNDWV3pt6NmXXMWo+aisSwjltHJyg6EwDRmvEg7W0YsJ8rFgq8BqA
GthBqw7y/nXpdyS4Fr50ByRqDvWKg43Q0Ldp3KAgHpWSz4w+LQ75I3c/DB+iI/4V
alxNna+mFqPahAy09pwW1H2t5cHe1EzJkdnkoF0IEr8apvaCKajOnhT5QIx1Am4q
UZY+l/5wzhLUM1ifmeZb1frBJ06QfN7oR1hS9d5TK/WHxYtBgKkimCzUHilt8FY9
/aN2Q69kFPxtPDJ7gJD7xvZ/EmLmJXfHvo3dsUa2EtbE52HCgrlv3tUShugSaqMv
CzDu577j79LUOU6pPrzysZ4Qe7t4+isKVJoWq8diKArsSl1Z8U9ODr420kkLoAX4
brFFgEtDajgQUriyf8oac5mwynP2A2nYVHU2RzIew8kEfShaEIWsOSFy+UYfcxY7
R7GS1E2StqouppAr6FQqpxMdTeE1JtmRY3lMIjOg4cWbzghFg5cTkWmHnbKBn/nh
tm42vGh98OoOHziOnWiKukwxqqJuIyCI/SlMLp1TPyQPkeA9q6tAXyQtgR2a8qp4
jt/iPkNRNqXVMmG/Bnfc1wIoucGl2peZZ0gmJbBHFfC9szv+rlNpGFiT+h3x2yTK
71h46X3CyHq+Zn55pGCzIpEVazGvBXhlv2aEnbsaPwzjHxdB6F5dAqYt9N3ss7Xd
L50/v0aepjnAbTpMH2h2y7CgrB8VYw9O/tl926fz02C4l0JIwZkEnJMDzjc2YZx4
OSSZYEzRmA2IzipVG+855jA+gH4Qf+ahrxCe//gHu9CWs4HRgbBMBJZEXBNrfYx5
IkKPw/yKWgaob8JrCXdgg6oGDzhr1SHt2IFYesgInZoilIly0oH4BO1Q1uirnsVV
BNrJTaEO2RxQ0f1BPx6GktOJjjcn/joTRAr77USo3qtsN6PHPyZGgueLS4SKEUt+
eBy1Z9AoJfhirtn1u5jsbMH8TZFO5Pm3JdUR7zqgY7RNyHf5f8ZhtzwmXhqNENHT
eWD3LqS8eTNvnaCc/Zs+QIwmVOVApNPJS/8GdyLwc/GWkfGogj7oGz4lbIvsn1ZZ
ZdO4J4lrWrfhjArXOtt4DWVcpDMSvol1X7kUuqgNsGAbQCiWP0KwkywA1/9Yzj4M
U5Yy4+XrLgyOE1F4dFI/r21Rqss5tmMVmCD3BD0+bLXg//38VSd0baH1hgcda8jY
89oeKQvcqlW27xBpfS3BTtMkaj6ZsODCrEnWBgiAsHdodyCoofxuq8kUIT5zgae9
2sTOlXJIN3/4Eb6M5dvW3Za4MFGeALpFG2jPVYXmh/tbUXG5Oi65Hnp9KiyGv/Uk
4ZFB/nkpOtdZfjQ1ADtzz1UKpZ91fjPlTa63dM0mMiu2JUzXSr3ldGZkbzCo74FE
rAi2MTcVjF2516XopyU44K5LAV1IxWojAkfCjU9h9Z6LuGGYbuRr5hQD0gAirESn
FttL6RvA2lgiYmmKhwPi/Ko0wjjiTwwhI0/Bydv3m9E1uHVP3yHdotN80dtQNrkA
YNyXrz+n+2+KFSQa3zMu8tQaOR97ycPD0dfkovfpTniWEhE0wEU0Wy7gUJlklwyE
FUAZCkSlIY8K+zKmjCeiLhkOx+NEaxIu2NcgOq2E9ZTh+qGdrzSyTHwocrtwRVXd
0wKPj+uPDp2cOYxFBk/OIht8mlMDfSTi+JJwRGA0ImlZs+uucm5/VWJ7S4JFG8Ff
D+FB8NFS17ufc3oDhmGgY5q9MtsShOtBLgIAGTiob+twPMuNJmsYYPaxP4741EM5
4LNM3NI+DxvpcFb2CE3gFYQRJ7ZABvnAUuTf8J0PZlWSDIElI6QtwcHm11vB5bXf
je9Umw6fmw7k7pUqmSXkXxoVVqchvWTYznsnreiMNuqousrS1q0dnAfz6sqfrJoo
nG+Phs7HsBzF5hlPzoKYChmjoiLNSdog2GU4xXCzT5MtOBYlt/Wcs2xxcAWSdRfD
+J3jv+aWfKvUNlp5PvcE0VVPfTzPo0cs+WD+tCzzvRMkZVfOIG4hGh7CBDLUpLue
4Udx6mYNP2MV8/Jd/Pa+e5mKQjk8UYpSrZO1m5DByNZtRi455NNTr8n7xWRBeAMu
NId1t8xkHU/d8/gLLSuCBfYJdxdjmD8U6gogjMAUs/sQj3bToDifZPTXVNnkdUr8
pciKoYyKkSKbT6A+4Rxa16XtffxyPqWS0AUQz9dXeFL6IZEkbHRWXYLkGFQtYcaV
B6r3Wt2BnoA4NA+eqp7tYyioGEBX3mkcn/QpbPO6QDiCt/ZAedrmq4JPbeE80crW
O5GSGRJem+6lOx7mQ6GsPcibK4oI61+oeMY+/tWQ6BHZvq5S6SVtOvF8/o0gQhAE
RVakxHhTfR+Vhet34zPl9O9Bm1mgl27l3VUHUFcXTog9YowH3OQlCZoAl5ugxnUw
4xlxw8q2cx3dBQ21G3QOLhiE06Aw8nG6cAd93R+SPZ582jZLUoDFGziLI6d6x1xk
3uvDtIFwhHY2rLN1vtAJDREtAR7Oh746euWGX/A4qmKyJVaBwLJbXsp19GqXm7kz
ZE6ABVUxAhMUgMDtVeomxzJPjwHQiPMxNH8uV4UNXTEL8Kv+lgnAi1l/Gii/HgOW
0bcyo0mGgB3jnh42hYKu/cwG6ybmyQv9RtR6Ru7uK+6BchBEvPjrTABTmzXl/1Ty
X2LJkDX1JAACtkJtC6QY5cA5bHt3jo26xOVqhIa3HBkdCqVBbA2x29/gKrw47EMI
lA1gJi7mfKjYyQyDlPFC9Ir7VMK2sty1mdvekLpdOBQ4ko78z73VQdqDCrTjuZKu
gkdrFVUsr70Mqk/40yTnbpc1P7B5QoL4AGqq9q/e0OsXB+aghhPjPGvNWF+QNXlx
A8VSIMUmqNAmlp6ZhoWbZX7Vb85BmM4d5/Tk9gZcTlm4/6pliWKL3dB9CwMloe3e
509e21EAop/ClssGIYx7nQZnTCNHrzW16F4DJtnMagURafGGH/nOqwntBIUy6IiY
FDJU3iYIRurBv/z6uV1+3iX3b1DACgn1/4e/ugbB5sogV9m4DowY4tA0viIYUe69
kkpGH2BnG71DY0Lq2/mKpvI6SWGjKMHCzVnCOzjA3dj24Y+K2gtj1XX50ahQbynh
yO5aDZRMpDMOp9Mi1Pf3YwyE0nngUU27BmYgtYSBF5hyTVqP8LXw/wimRj45yhxk
ua4KJsnuEP0846D72wvn7P+ih3f8KOLyUe025VgjTR/C0fh9U599BNXWGoTmRCQx
G6Lef0Tm/XTBK7QVeROfq21ciEbqfB05QsT22ygOkf5YrM5mzUb7gSbWq7v8fIY6
3DrPGSLuUB8F7QsZZHpy/GP2wIRTMTfXQuu1bQxofqsLCkUya65ZKA5PQP0ouGTA
zkpfDQbHh2doJwsdxm2T4Y1mfGufQpYwMZPaRSLjaidmChd1Yl0ayDWiMZr91MnS
FeGBrx2FYlC5FCYoYb3Fbtn76+YZjEIJJMKpNR17H+ilxh84FfcF+3SvVkLuWW23
SO6UGOXAauR35zyDyCUwUfRcPV41WXse0EYABgrgKZS2WKcwksTO8GZL1z7+1wLU
TV4Z4r/bZZUZ2EK87tvKLPf1VXtmfOTRpiuu5j5fmXQwvYCtiM6LpYAUoY8FWrJv
+4s8xgYjWKe9D471XbBANfNVbFi/57GMgWZFfBV6PGREkSzPKTgd8OCjvVsItzBh
fDxvaCnM5NaH560nlH0a5GAH2cQi74K29Rl3gsYS6gxjHgGfqg6xhd7pnF6YY8fZ
VzbdJ1xdg2tuRbNUCRyRwTwvEkhlPbjpuGgj9IXY6N6yhiulyUZa4ml9xd2Nxdc+
zJrBNdJWI5W+qeR6NpaFnsUp367wnAVTTx4dvPZAAIcjNdpLparOArgLWGHdHohs
WzS7sqxkV9oGcFEJN0wsKb3I5UgN/EkPTbVpwKikNHstsJHFiTlPbTKY3rGKOHqv
8nhvvvnTFWleiMh/aHhWSMZ4ZlLuPyaRWxuSoIcFjwX+Ect7uRSkq0cVbS4o4Btc
/VnLH5zzkFzRg4qtHOfjYUNFeOpgTQj7Ztl30n0ExHzUdik9WAKSYhBp902tdLss
aOFkvFBYp9vNIkgK8CKDbLAMf+el5cPxQTv9WIJseDhYcSaO6/gGD9emzHtST4Ru
z21b2ODqUXYY0sokm0rRtSqmdvChczvMZsG8aTwJ/YvQxn6t+cAAukz11cjA3s+h
4EOGpvUgDDRJeGaIooNTvqqJvd0f/GtgAttOGVKQKvG8Hza+ed+0Xca1kMZqCA5B
sjcSlOK7SWZdgk44n0UsuEDKrO+r9wHb9X+gVJYv4BHa0dPLzKlkYsZowZwGAf4C
73bDHuzrCeXrEdxbfG+MwPQrch9Hdl5lp/AkNE76EwHBokN0MTW0+PWUnAzgsblw
1pqa1pElwMI9xhgSB8uTSUMtrfxJ7V3dGSp7yAGzIoAYfJozD6U2L0FBZxmzqDLQ
HZ86tyEtriNDTDXoD5ZY7qo4rWzoB/j8fAkM+carBfWt07jb0lbwk+/aX1bBowR5
YBcSML0m0Rvq+dSQPgfmuhMy0DaKrq49eMWR3ofbnHoQkhBCmaSL3SA0cy/u1Zzk
Gy72T1NpQUrd9U/XVtZAEUyZBCG4vqmYp5+QOcHTQLFrJqILDhyjX8lRsn1jagmV
dCA1IAEhuAx6FcJH45rvF7tlq/LpFhiFwtgYWH4QkReJPAZPbnNWNTAjTLgobMQx
YHMiG2wcA5D3WVmm2rPvfT4RbsSa5OmYLF/YHnrWTBwD+p82kGxXpAIt2HZcQUST
QNJ3nYx6o3DbjOm+9rGsT99ysofvYWOpJDHnTOU3T34U+WPYaP27q6Vd4+NS8Boh
JUr3zKgJfe7so5sbSpR4qw1nSX33OurWIs2ZjAFihuzeFguWo9WTAqS0O1128qgK
NKC+IEabPbHftfAFQsz/uVTAAKJWyQ2tHz3hRTAWoUZySu3Kol/A+czz+sVMOarz
BvYkK68D04UUdDUSfYvsAOPQHUJ8AmX3tDjI2J4OOOzWkdPgDLzgrkNYN88mpZsT
kU0bxdhY+BegAijgBq/KqZ/qHZCcKawjx8ndEYJRSf3KKatjqhoqD1Wta5ryYU1z
SDUXtGgGWBUZzBZmV9fxcqQY+FbY5zpu8DPrzoytLYmGKNqhRC/guglIFjWC8n2l
CZUnpu4DCY1goKBezyLO0c9705TXaw6oJ3uFhEftHs/tX0ILwtD2QuBcs3J80j9c
1+GBGI/fEeYVhNiFJQTchZn29PPd30v8hvi60Rk6S/DQR6kz8RBnxM45EqEz+Rt4
fCxwKt4WbL/7rj47bbxXb6dzODAsI3RrfIXtSW94fYWGdGTPqpiX6OsBZzaoc+By
3BvDyG2/Q8evnOnEZ8qF7E+4ixZmgdCxJNoYUgGFAsHpj74l5IRfn5o0W5vpxr8U
MvJQkSM/8PRO6EIPuPmWoDOdQr7FRJIOemXTXnE9O6PiO6ykkbW4NgHJS+p+0wEt
Z78kmCA1j2P3Ydl/d/1hlH0KwXgCdvt5+AYc8OAkiK1pT4WmNpkWxCmPvn0Egdau
KWiefo6/XsCpT3MvJpRaeG5RbUyQyo71ZY9L4cBIt6vSI30Pzuk4P9jaY2tWI4be
pZNoY5svz3zJcTNK68hZw5TVUG38KzKQbhUKSQoRZa1Ks36pRr17AiN5SJVtinYs
1MC60s4x6NyzD1X5laYfMcC+clAICHYVCTLn2LxIbxXx+qzk6vhEhQm+pOQ7bFQU
NcIeLCzvnk94fHn1Msm+smXV9a8esBb1XIu0hB569b7ZJ992cQUA6uZme4+t+tSZ
a2VdDl20ywhycuF9g7rmdWYsVhz4yNq5XUYFrhcj1c3JVSF+uXiNEuJm6/f4lO7g
gaijd+SNLELNhkhH6s33/Puhe8vdBTrKYLlhmgSCvqs2ELRQnZ0Wpdjm6xjatP9X
zd2hboYcyX2bKqjFyZmwVIkAdd4nm1DJoCEKND2GC0wA2q0kwPtz+3m+glnLUQUv
BTabXOQ7qmgnQf/4NVBoEE0N2jG4WeHeUFEBKXs54g7Vep052HpcZy89v74FZvYw
OYCj7qgox8YPyIrep+p2KBr1QYXG3Yxs6CUTYJP/Je/Jp3woYs8x10lMNg0Qzw3o
f3JHsEcbBltvRVuYIs03YkRz3CmNAOvD8ZD8fguLgKNVIbztW2T2wbqlN4p6SRSj
iNI/f88cTIlkeukRMyRmrcOT/b+8ogCDoFsttBt2qqv7lL90r7Tcgtm2Op0z6IFk
iIDX6UgG2iRVuUHaVkP/TnZYTJAwc7jEfVsrnpv2gO4S/7P2iw4ctIsSDlhQ9SiN
kaeB0iQZw1mp68CVNKf/crXdSxXdRy96R4n3/e66+0S6NURbJ0c515qj1BWrvo4S
vxqZWkaNq1cO7j6MnrnLHwlJQqKnYKJm1tQD2HD9atsClQuJSz85CeB3ZA3P+wZw
NqXoJS0gMbT9qWMrxnaeKkao0gGgiGai/hDw8RnLOslF7ERwlFQ34x5mR4uHGlww
vdlFn467ofF2dCq/1xPKjrv9Fz3ZMDBiIM43qSBFerklxEXQwv3Uz1Sw1SBb5Y2U
lwTTKjHknGVPwhGfft0CSNYsDq9b086s6QihebtHT+LJfCQQvm+A4nRi0BLyTnld
x5s0hKXG+kiiPzTBGn66HZJq0u2Z0DNx7KUarrcL8dbX+GNIwBlfmS6KWPnq/R2v
kJJ1bzG4LELMb1/1BVItSQJpO2Mari6p3B1ekR7G5agukW49FjNehMG0/qo5m4c/
xRjTPzCh3fDTmNp9CsGrU7OiAfxkqvcvHCi/AmzS7KMVX5rGIQokHODwZYQwKbkB
bcjzWYbuHD74AVA7eDxrv5cRaqvhrnC7kXBZberlUwtt6vTv+eMnneSAhX44huhE
XPS8vN3/3HUXBQ2hcmg47hmiZFwswchSwIx+aFJkNbdueYgXC/lUkLwFhdcCXlVP
//QUGQLcE9LT3TLE/P7IxESeWGZaol6C/FqQi9PhJjZTq4oy5VvS9adDbrU3qpbg
yyGvJyrwguTl3KsTDNtADwo9Df1fdlzrJ71OS0v4VHZRp3vpwA6q5ChLCaimOGjH
GPvY8uGhXrJFh3i4RlozsWuL9tNk+4hpi6FNwEZzqF2gElxueEK8X5xR323xnCOk
2hcc12w97zYqpbOJ0L/2DCbcKAg/iyV1QKPwh2pYco+GVkzxS3GOHQHG1b7fzjPB
SqCHujBf8ha6ZXhunHCcSAJHUvDYJfhH6z+MacuOjhM6+166vxJsyvLZEeUgVyuM
f8CqKXatBz2IGhF2927Mkcg/r3VvqC3f9Xy+3r40fd3nX8KwcuWAMKAqttno1PpR
KKfeYU/nv1SsM2d4hK8OkoLqSgFYiL7vCzHqDPBeOQLtODZg8auq3CnzOd1ajNwd
xMdsGct5OpxFO7CNmHyGJ3Bhqd8dWdYOEZbOj6sbJGu9OzvERi7OSgDzNP+EmLpq
3yQ49epy88dxmrsLf4XYvWy4OpekdHQ1ZgcDPavXvqe5BCD4Kdd/fU4a/UrJY132
xr/+nobY6mFr3KZKBOB1f4vPOJiufYVX2Z3qARtGfe4SFMKWkwB11TP+xQuEsxXb
rJPKdn++beOHj26SSKzudDrAvJzqIbcEr6TEZ4YJ6A9wlidLq+vYqtKAjeHDGKHx
q+sfW5pbMK8DY01XAVWGFffSHHY/pK+H/Y/xcDz8hdW4IogNfx4eDsazN1sjmp/+
7apLhYMt+eKd8sN4f/Lc8BZxe9gRPKWAVGgK7debwxijqdrelSvdCpLAayuKGKMc
J1ZMheemn7I7S2/ywOdG3GmeyrmMG4yG/nA4s7D/MZ1ZRbLv7KkQPUtDcYbFhnCJ
tPo89Cis6ATB9MLh1yAj3XZtX81NROX87DhoO9iVHadsHxbQlMwKnIV5QQX0zNNU
3iRsN/26E8AJqrKonvVZRFMhiQX5/HCR1A7Yx3ljyr7efUY00JLSv3ddeEX187V0
qm59pftDPOix6i2i4VDNoKt4MDSkVBO9WjNd/414fXlerTMHbRmkxlMPUsaOf8h+
7/YfBlvN1Xyjc9Pqv8jzpkG0Y+XC+G3xywfvBsWol0R89yBA0gNpXxTCJjHlJ9kh
gl8q/8oU/uEJ4lVGLzHTZ0fASTNfj9KM5FU2Ww8gUFaSG68WDfhkiSDlroKW0ri8
Rdr1BCeBCP8njgleIQksM2SnNz+Ygj+qYGOIJGViSKSWH0IDxvPtnitGzMxna9Su
rjNetM/HBb+r5q6Sa1nDhWIjoe6rU2LwAnHrmygDbTDAySV1ubtsnqTHx0eKNbl0
2q4XA6za7lasl0sQoih+x1DAQpuoBjcaCSy//WbwOuIj5g52Hr00zmROEa6Ccm8d
G+UrRL4pU3cw08nvfvS9FsxRnqyA9vzrxzkYylXlC50FDsnYkil9UHP5lS7hlNHd
eqVbUGoLQzen+UxcnrKp7ReAH7Q1LXBa/XMl8UkJi01UrEySmtNGuiZb1Lf1rdBo
OgVq//a/jR7IufoIVCuo6TSBfNvbo2xkVjpC2csFb1qp/K7WSw/B9mGUIMosq6dj
sPN9qXPMRNCKKCcE37k9vR6vKH3Z9im63B6z3ffjlUGyLOn7dYxZtWLovRQ81gxe
4pOctKxYPPRlbglRpjcVWSRYu/Q7bqGbJz7/5o1OnyzAguFC3CIwnkOjb5cjBf3T
TARicmQsVpoIKoBhI4En/sTHXbr4SqdJYtZfcPICuDjpAceMrGBZYa5oWMaXom1C
NdVWFauP7vpD27EDQqr1O4oK++gievabcAmcDop9O6jmvljWjQa9cF0bJ/JGhcIP
IEFYQaZ+LrY1gVB0uSg6MMuRCSxjeI95zoHbhVAdFyPiLgV72+eoILVmDcrgsF3G
/7ETxReqG7bcw6/BBKf2QpN/uB9SMChoPyJAemjAXVJ1SzKkBFDCa/NJ9iuqB+D/
WjdpKYQ5mj8wTriYvMn1hJFreyiJ2UdLpZuPLPiSC4w+KYJRYxHE1kZca2vHF7rX
5Hd+/lq6eQpxIrVzAMlxVCy6MsZ+tsMSrsOdUCVECNw42lvFjHsAM+v1WcrQDplF
qrKr1Xrd07hYPtFY6rz0wgEU60w5B9twnH82rkpFBLbA557tzb2kgook3ckW1f/k
9vQTDSvxpOTyh3q/EkNDAack93+jBINmvj+JKDbuDBttf0E2rTVA7rb8VfNG2e+3
cK67/aiPXjjyI46iEdH7ntpb6XqmKUpG2M5WvjMvYxZnGMvXphI+wcS/iC6ZsddC
YR/TEZYvQYuM5Yq1lBKXzg8H9sfPO2HLxiDSELZx6FgRbRHcFN4jbOARDbPu8QBs
wftMO5galjIW+n07yr+KVk29uYcTjj8GfMEZHN7MR1Mvlvz/t7NccQuyTtOKhIEW
9ac0OpbP7QoEhKphTkt/8yTOzYRIkn5GEQXftgmjRj7ncuA39G26v9mwCbEnzo9y
JWDQLAMzwGbFI3wly6YCaJgpOrrfb0iZlbwu7Ow+zfKdYzfVIfIUpxQBzHyRrIHm
e3/bfJpXHiWIHvlBTl/egRO9jhznaFTEXSkGJKkkyrsSxfSk20+/OknmtWp+cX4S
ompWLH3+sgjLGLp1QidtV0PqCXiGl5w60p8z2F+YSIIEog+J2FQUKlYgbFoZQn13
hGWSx8ZWGYK1PYQYz6n/z95yYRBiVI3/zDt9uYvOCtHyCiYeqO+81kd1WstcX4A1
tTKvQ6/GWi+LaIY8Mk8iX5lZd8qUVdrlkPP5NfMb1gUv24nzr1bvLCwPbfRYtSAb
ud8/jmqAon4FuiD9JXMQiFSg/psaV3W3Q8utz5UbNnqh4OzXg+vXutnlTDRiR/VD
0UChXEZroTrF5oCpMQnif3uhGdGBCpGrHvcJp6Vvy4o+v2aayazbLADLshjp9Ld2
yAk/Ldglh5AyGHn6hQxW2dqNRUiXxYXokB0UxpK1Z220uYu9MkMCLkQIzUWG9MCK
P11yd2epI8jEC43/YKCfR1whZBpuDf6xo0j0mtNSabbXkMWPve/Z+j7WyZAmcsH4
y+K6V9tS4r+8FyQbrgnV5QZfBVRvFRq8QsS1SpbtznA4wwpcxYfMhy9khHGGYoM4
vAhul0xeleKvTouxsBl+J91xvCVrcN/F8xxB24gqf+nXQcfFhg26ppAsAQgserXk
95L8KC2j3qrsTQTf+v2MJTjeEEsjklMiNFdFI2mZPfdst4PBnJdV0hQgZ9IT04od
v/XfcR3EBIfDCtP2Gaveb0KL7H9b6jl8bXX7KklNG3OW2oO/tQwLG+H6pl7G4lrB
A3xOBGlwarrqAthJpjbv1UDrPxkfTBk0fNoQeaaRc7oEHFi3nL6SZp3fdH6pGM7A
IiJZePyfmiTp/Kic4RZJF7Sj4fyKziTVHvkHBwpPdESks+lKUiI1NSFWmvCZL1vo
o3NQudsuigqD2VE3moy5iJOtMh6gHurzTfGOpOnnqgLHUvlWE856nT4nznlz9sK+
HvBqfDt2fnMea187CG1VkU5/DFpN0sbcguh+S/Lhw+GHsJz5g9EsA0QqNVPef+Bh
GRVagzPt3vZCc3K1GrTwWfeXnzni84Q0slSAKB4x/MKSOH58UAS3jI5kaciRxP1Z
mKQA1h+8Gir/UC0PgT17NiWrQec5QMWyGqIyBnMd+zLdMnKND5VkSqTrdooZ1kMC
jS1wa8nMFks1hUwVQFOt8Aj4S5eWWGaBo/Y0qogAaGEpDMMLmvj8ue8SxdOwnVlF
0aMIZi1UWaQXZTk3mKl5eyrLa8Z7ScOP/D7UcitFtJbiZnfgUkhH8/thedGEzgTd
iOmWS+6xZaZr2BfZwHfBPXahUkGCk7gPT3rn7MxVvJCboWrshNmt1RFBxAKfw7Zh
cLgBwXz8Fyopkpi/w9Gl/GuZd1UZdXlCw84duv8SnuxdQVyqSrZxiamuaU0oxgIL
oGVneVoPqVRu3W3g3ZMG8Viu9UQYpkxzE7Yevuii97Dg5jI0CxMvD3Bfl/wSr4fV
qPZ3u0u4u+4p52AERWRVGX/4cxnknsiE5grgucUr8mCGF++YpSG3sYvwn/iHGadN
4/hWqmhmxew1+nnh+xmjfGwiJV+ejhvZwQc/Q87mJ2ItQXcBhHxh/4Us+7iYpRGL
K1kCIYADvIt0kwKuRY4jN4emwrCAlIcVTd2b9Of0w5g/fWkBZgnv717xbbe7mGPp
e1D4PYL8xbGfZjxqkMvBPs8y4FNwyqE+VGJf+oMm/VNeT9n6WVk2UHH8HPRO1iFg
DgHXPxiYNOYpQmWvPjcX6MTfxHBIZhNHBC/4+xRliOB1T6YwZ0Vl1gRBsmg61bbR
VfgjMBlCS70NGm8+oQbFDyInKPFYx2jETjxX/lSQbL1vej/X98Yn0r40vMc0Piiz
E+8ZekYh9IowzCvsKriJlUkzO1YbCIaqi/j4qNa1KWuvVB34DkEbwNzc0nVYLguf
27JXvcDQ6rD6IFD+X6glCh0tkJ75FgZ5SFp3694UYWXKC2aucd3jCoKsAqU//Hr9
UIdiLf9DSzQ0HL655uPDFkYhriRut0rkYXaYS/KY2M5KTtN13HFkthM56mRIcI1H
NVFuJAPkhFlgsTt1567N23/Y1ySLtBoqn9K2mYBENJFsfbw2o2QXEQCrkUEHcLUB
P69IfNlJrnm+CcamxYjCyR5A7JSBC4l0PXcVZamtSBdrRN5ajY1oAgjQpxVaMbfH
v1UbF9cqzZqMJfdtKCHL3OilQWYB9QRFBU2cshZO9k8XNUdkJzvYfSkuXYSvMtGP
AHm5dGPx9tfwoCCXVZ+U+fVGTmEUtc/9qRIqw5v8eo1HVmSLLRUjjMWOU1zCh0v9
TZwAer7V6gWfUoxbfy2ffwQkG4XmRvHCzt4scqJbYsOzB1nomMXBA9ZNw2J/y/Ws
LrAmIgaF9aSZf+Pb88vk5rno7Wzig4+ovx5nIujE7um21GcbPX/++2E44PH9aSua
lq7I6gKL1/AvzuoNCDO/kHaf4/X97YBrWLrGFy9zPC2hfHfMjIP+88Fcs3lGaTB2
PVGOaxwKvd1+dvLAU/TUdeYyjRH6KYIMCdWOn/7kOkluDSShr+vGa+BZUH9jCMhL
fg/muO8AfzPqxM61K83n3ctqYIaudGBAfEWqVR1nA9aYpr6CaGgLxEcfiMdsDo7H
Aoth9Rl4vj6glU3pwh2uo966NdycSl4dgziMfB4sJdPsj7fKimmhazITLZDT4Qhu
4ckgTLSmujVmAnpMdj4BdIoheSa74XtFH4oKdg7gCbujvuOVyEzOhDHURunG/MMd
tbxe8KENZjVS/ydwfTQVY+PpQP0qedU0sgPsl1Zapo0RqXuuyGxIYhQ636njpwuy
UBTLlq1srvUadaP7G1NN+yt/frdHRurMRKnchPje2jU+obkaocHqdi7cMIyViC8v
Jq6WdxH1okoBQgBw42K9T45CeQ0QNzz8UEc40jNPyZS61X8xodEGb7Xw+bKt21bd
04D/wvHSsZQW9Tjvdrp10n0QmoZfESWlo5ur0KJeFprvCqeIX2HNBqMX02tVmLC/
7QksMUw+hDVHE5uNCoEFN8JtzAKZ+wfQEyuIE1ChB3Xnr53ePItcFk9CwG8ssp5R
ziyvjzywPTZj+uQhTb/JD0sVWP0usqd70OJouyiDYp8p6QLfgI1Ir+wy6C/B1azk
U2Q9T7Hfzjdb4BAWs3YggKfIGPc1r0OfoN8GrJbOSgq0envoXwPB2ZwKYmV2Fy3w
h2CF01fWAs9f6gr1utcVNL+226KUrPuaOn+4uv4n5MCCz5RXn+0Qdxry4ItO37ds
v2NnIULiW4OlUlTJEKQcdc2Yk2xD9CwYmu0zx0s5ab9iUkqmoMMQlzOUybtsYqY8
xmhb6mW63PrLBMEPBNCWLDHElQ9IG3A26VJq1J9VrictNsdcVoEwmlVT8YtwvDl/
QVqq+OtaEbsYruYD73LxUomO3XBYnLFZV4qqLiveWZioOJVIyHr1x4BRGSvJh0dt
+wSbWkm38Qlw/0LRV8/ndaU7DXsQNZ85GrOQf/QeEqeK69lkkxQ9CoT6j8wGi7u0
nvE997INeMiLBx6oSVeD2CZAO/AHUGz6T/V/2EaN6uJjgY9Q1bd9iozVRjxVCiFX
O+P+VARmZEUQ0hicM2bdqhww3YrMywAblpY33of10HChU9Mb6JsQgwQ/0vHg4DEx
COn6RT1iYl64V7ZhLVG7YMRYUaMLJfwfxxuUJW6kxckWcJ0qiLxaKx6QIpBxXGiH
kcj3cz3pAGhNBiaQxkxrFw+snWAn+dcjxqWnfxc/mcj0eUJJpO/TqwE9dqCt3r/n
BRDt+cIHAiRffhaNcyqOJ/CuRniEjmxhEmn+k236jzgIfN5SKdSjc9fiKJKWERcA
IqoUecNcVz48P3PnwGsMbsNHyW31ezLUNUm3Va4a1yRe+CuAhY2pLaqxyxeKQvfs
vxPp9QVXMKETgJgKwHZCI3Y79ZT+n5XmbyKRRkaYKRtkC/1+Pe7O69MntTnANGgm
v6mkq3stSET4cBCwoUuozV/AMnXCKVaXnBdMNbZFC6yBwGhfaA3Md5rH6t0tSoTM
ATiShD0L6ylkDY7v33K6VWps9XpoA+NfsLaD0eM0UfvqWPLT/WYie8eTApJeaa7j
mST3MOmjtAc7aI17wItj2wrpzxwLOKGb8E31rzZmqf8sA21M1q6YleaArdfnBkPg
PdegkgN2rQ8lPnKonei4sV8ShLgxTS4e+mZMGFvhZB/ykOjzT0poj7Mb5CPJyplC
H0jf2VKtCmeZMVHMiyPUwm8QzUn/C+XIaWnvzYMnl5XRDTIOWyA79Pndbd4E+RuO
47ZbX06idA+gLSn3RDl29uIj34Gy8/3vWplnxZP+lnamGPqq5abJ1lMkpdlUH70o
bFRvn6Il9yUY2o+kBi8nhui1+CTT+QBIRPAomSNlZ7bmXPa/oVbLy9OLuTt+yIH6
b9ksq5eHwMzjk87jtMMYEcYX+SDC8GybF+T9vQDSiBjM66maoyiEKnLGHJWAcLpy
P/3DOONAvsS043e/xxaTl7hdUyBYa8PIlF5jHNmgZR9/aLNi7U2MP4IOPfO1MyUd
QcYOiwO/Ovp2QW0tqpyDo8FL7sUxe0LlThSQh3V7rx6nB2PdJZo/C9Jiqb+h0oDR
dSBSNuBVx3icOlgucWndsFDA1vW5Dim72+WoKdCgvx7sRZ1PNJIYZ39/cnO5WjMs
y1eYv2D0uya7JZO7K9ZZ0GPn+5Ap8If8N3yGO6iDyrN7vx1X/bpADbjbEMYE89Qz
NMpskXUfuo7m1YJnTLHcXrVRnoSl8cN7UsmpMi/RIpljxn1tlEZpkaqc1eMPn4rJ
k7l2ddrzV5MlMwvlne+gWYC2P56LkA/oz5kjmtXXZdJgJ1c5vXLEfqdVnMEh+4IW
NkP0t2qOzVR/vOaqyXJby6ZRrn9Rz2f+YEj7EOikhtNmm/H9E2HP7pJ5L/wra9EQ
4okuuHGYIVllxlFDE/YPXKWXwDrE+n47LiU93/ZW1V0xCCtXfjS+qCJnz59WNI4B
/Tv62F/9q4pze0GMat5FktffItzxLQ50gB0nBUbQzmlr1wbLynMV6JTFkSfKSWUy
MIbbzIbBtAIXEC6vv60Gk6hdUplAKV9MVbiyr8IxO3+wNEa5Sjb7KxXiaYjBa7ud
+1mT//LJ7rxVhp3jEYWScwSRHmGFNWTw4bYj+0LszefUC85WbYtka6k6VQTCc5R4
7yJXEloZxEEj6XMw474Jt/APCvvAvmHV58eCNC3bLuw4/CbSnw/wPKUckbbt5/4h
w3MOPfEaBtQ+f47LFRlcq/mAsz2gf0PTXWfTKuxiX0+VFIOG9X2V+dKbns0mocsB
BWSjneu+kQKEAu2X47WOlB7ZzMn6WG37122x9PMb2MwBzKqhvFY/IXoEbsdGm7hb
O4/sKQiXB+Buj6TWFz4b8IAuLU3nvgIwwC0bkSUQ2fkvPIWfc7lntA0u/NuBffBB
91PWXMq90XyRo1AqSx5BqxcLSsYgvDrJrbptZeXJmL39+lElASy5hK5DFnItbD9X
UXdgjsBuQzFFBPu0NHRqK4HI3iS+QubqQg38tusqcxKZH/JN0CLIxCP/eiQw1dUA
FiDnuoP2eftIQgQbVmsId2r7xrlS/nnHTxPrE2D5y1cXac2MDRfYOKFh9/WxW/GB
VWlebdlO1TkDcGGCGa+AeFx1RZhXZ8HhcffvpFtyFQTCx3mmxhDBHHwBILwcvqMN
pyQE5iSfCG+XgV8KQyAOHu7Kjc+0TuYdgDshzh6mH0JWDCxXHz7MgvhEn4WvuFjA
YqihnUai+d44rOO6IY6Cit2uymJ2fkWx1PFi2V8SF8NSde3ZD1CJJislWCdjYeSP
0BcqOTRLzKiy1bxrL4bHDFlSl6y6QkZoD+LSrRI/d7PaU4mmFEwj+BiQeQPJuR8W
ZPVWWZNZ/SEiS91u69qhxoGF3EmYX7V29A+C3aYiOj8XQDeOtnrdGC9L0Q1yTnjj
nB72tuCA2Z4OegqfmdGHtjITG9mxHRb4AgnYDhkkkmCckTsiRnpBWzYCr8UG4LsM
k8SvyngXZCHMfkL3Gr0vQPLoeIh5r7nw1A30mzPv27Falmc+HJ6AQErGaF8fUmrM
EcV5IYKXOutB4zcghXypgWKB5EfCB6x6Lu1nk6leBPpSUbMHhDFz5TIMnwXlh9wM
BABxpZoQB2Rd104n2f823KS+1qoirCTfXER87iu4VDZaarvR2TtGpn4KfWWS/E8D
WHFA4r8i5NBteyD++I2L2s8mIq0QTCe+9MO+zgOJSXcTcHxGNYyCBZMuJlPVZbZD
Rvw7ZyMTzjdvua19ZOaCz9vp6nhoSrmEMVmmr0wpY4kfeXQr8RDwxeIw9lTE1COM
uigVQew5uJtg0GLMvQSCRefzBfH+jH8c/pxdE1BxCxb8AT1eH6e08ur8T6oaVly2
DzG1e2RDZan/B4aJ1w22to5KFckLHDjzebZtEybxy7OQ+tsm5ija3gJJT27D+5Cf
zEQMtdM+ioSs3y/dIJ0V0aowc1zu7ufJQUrnj7NN3UZU1CGOzryC+gB8WCwWKzoq
65/yxVRuDR4zTV61kv10z0kkGV2kBVSuSWkSCTM/OzX2AIav2Wm9ZnnQ6HoPjo5P
vyyPqJZEepgw/z4n29RDgv1FMcRXw2bPVKgrKQnKwk0vuANqaS/3llLwtSApqFZV
1C4e00bQwRW0dEJKCOuE6SI0QbcHVjDVtb6L8ubhJ1hcPC8tv1tmugw+XrCIO9zb
K2UPJi3Ajy5EO252QT6cETiAlhPtIVFLh/5JX6p4nX+vMqdFbzEiFASdQzBbawhP
uedru/0Jiuj4UxEx7YZuU3T0ZPyTqmziSmBMTmMBWXjp6u0X6I9H8dt1wtDdUBgu
1hwfJ/fm74pkOYEYgdxpD3QLX9foHwFUWpFLlVg/5YoYbvTGhR9TkQJNnNjuZNXy
kaBXAojDbLjbCCCnlnFybBdKzhImLPo+QSCEqCI1vRSoe1RUYAVIwvQXztcbaJbK
yolVbGSr8SUubpSVGXMOUv7Y6QRg67BfeqnX2tuRuPkSBKa/78zJzxJiIceqn8vc
3HKQrZCSPmS42RcrvZXMawnl3pUi/hloduPYAMNvle2orNZjrqXMWkzzeCtzNVdJ
a86zGWafHEPFw5UwWaWpSeCDdWKxgjmPjUiHkzlD596h8vrEFTDj2z368rWiSeg7
BiqNpNrSK8cXf8+uvFL/wyNFuMZAm9f/E0m5dDIFJ+z20SmjkLlqoL2dwONzhmCU
ytB2vjazcE30g3gi+0GgbVgXBleIa31qEia4x0tdwmtVrcwcA2SyVsDHz/0gDd6S
RsYrrh9Kk5jE7xvUY9cuSDoXCYcFdC/p6m+jBCTduKQ6F13YuKeN4gSMWYqyP/o3
7Xz2PPxJg/IAOaG2DjwxUvcqqQxq/y9uNkWZYistsSnwcnj1bsTzGjjJDmEIoyvI
lgEyKfzmm6SuCQ8XOda3/xbnKQMfnoxE/Kc/mfYNb+8RiQt0bHp25U3fT9//G8ot
aizWQoxM/S90bSWyy99Tz4IZ43/lpyof9JQXsz3OzUVHIaeyFILYvGe6IRVeKlEo
+pLdZVW3hB7NEaE3svXW+oDrKUrJSdf2hkIWA5tP2zVEGWBxcmlU2JK8Y893Vb54
7Mk23eDC/Hgtem4KPUjsDWpXgIXwJAHhkp8uB4mOitGsuibZc/MxepeMtg9FInwg
jQCKdmMBHhmuB+0OTIpKLkQLkanHLi494yfoBKvaJzub8QY8oNrtboRfpq/lNjBg
4viF4C6hkkk/sw627u629sQOZiAC1jEbEYZlDOobd7UZzmJRVAtJkAho1lVJc51f
nCWkiK0AEUogsPBjhHfNr3j/SgtEH7iZlTFwgsOXEBlEBCEBMCsZ4mRAuQM8aFYo
GxEvUfBzuSHy5LIOI0nWS1Ubh/m111YZMq+ieCS7N3TRExLiLusxlsukzkzZldTP
Uh5dVSmxguEaBKulghvbh3M+VjhI5Z0QoCK5TIFVQorr7/nkEgOoJzLd7D+CAE+c
GUfagFoXjAaynZCZD6D5VonvGa7o2bEEWK52mzP9SYnozTeK6JKAPrQajqkanfmp
uTZGG6SHQWuBYRQeIZzwb8m1dlAUh0l+J9szMPJjC76y0AIFV45tSE4UGO+ex4gw
zrth6x09BtxKhvmAT+joDqDB0pgu+OmtWDVTvAwn4jwLxk6NrpXhfYiJ1P4ptSBO
Ys5S3oN4TMP9QFfQrzqiDZ/dRoQuG1c5F4ctLgeB0oNAjTEKwKUHDYDT2Hq05drN
RBOeH1wLCTIYd3V+YVYxNAU4B5zHCC5ZYtiTCAJe95F/drpsqnf8Q+e5ktXdTavZ
LsfFVsMQNfMq/VUBF4LRuAJyfzULprR3IBnOGNtkgOl8nefDJSSMtAyThTlaobQt
5etcWZO7pvMHHnhWbP/IYSufa/EjGr8/J140J56IAYOQ0U26rEO5Zo8CfjzSOMRR
1+pTJMFiHyz1GRBfFLpCZzuGo0IQ8d1/zWrD+mxSMOHZFuqO1eciJryOprcWBouj
VtM2gdJ3PhnHM3b5J8iStX3S8DsLGj1+S1vSJVsxGnWF370jP8egOjtLSUDzrLSd
1Dfrz3Dhvk2P1MmF1on8Zz8Iu69HNasyVuZ2I270HRTeRoZw5cm32xy+VIxKHUbW
dHtJE0+3uy22nvgxBeyUQI9vH9eCUdJ2mHxO7QJYcgVYRaI7mUrKwapkgYPujlfb
egBbmzDAppvsfHkD//wg+QZxXKrN4R1gSGlmbm9d4ZivqjmQAnfg+1+1Hoy9MMte
nvCDlG3zXAF4u1Ym2oVBtQbuaKGYIV0aXKTDTytzob7Ed8GevpFf32E9y4hi3qBZ
BkYXr/Vq+f98+6sUvs4y368tlLA+h2S6h5tYGEyfotA1ZgBr/YcgqAjZPguCRk0A
1RGTs0kiZO+An7HeOqkj/rmtOcj5dtFAk+dRpgEYXKDiv18Ur7vgcA2N8qzjEJCf
TdrDVWmhMwaLNHzMTYaIXSuatUws19aDpeMO49zZ8NEbsYDbxL39y8g88Et3c9fv
VSrnpKiHEtsifiHr+oqS7jNBgMtBejExt/Q+9TZtko/LyehKBDqDnZoArxcTYDz5
X8eFFgv3/ijU67+hO8aNtjYB/kIXJKJwODjag0mpX+zLSR1BybJLioGM1nZiazCW
JEMl26kiuFwC1ElbGHJML3JUl/D6DUedPrYqSFZY1N+8/smtca+fbBBzv86UN5E2
jEWYZIE9rUjfD1y6hxi3WwaiH//WFcIR9YW2dpjiwxHTuLs/+rxjcLLXq0DDukvm
hU9V/Nni5R47cMIe15CP+nh7+q4ebWKhIawRmZjrzDREdzKw1XIpNx3QyrEw0sEM
UEGeU3h3R5G/GkZrcY8Q/43O0gyiR0iBEt07MgwrshRz55E+ZdrP/BIW+x4/poj4
RHoh0PdAgVzNlUnrscaVLHweikNLTjyoZTl1i6gRwmKVcH7xGhZKp6cccyolTTpY
BJVZi9mlomih0+O6ZYwEMNlhKf7UVEyUV99a+o8okDe12x056+4ZD/V8ivOHtpH1
pEjy09FJ42ha1twplpSqkULVFw5W7zDETL8HyNcVpqzIlovnu8D8t6aWVVqbL8wx
n7m2fyjXausQxoBwdVRIA7tZeBk5r8LJK8QkYLJhbjIIU5n5snDH9gmxYMZDY3z3
ib/E5IiCTsqAcMn//QBaSJTPJN9XMnp8oPSnBNHiw83S6h/N3oeVEfqQOZNSRKdN
pimoJWBGeLSWzrG0nlkaTc+IJgRsNTxoWB6wav/gSPO8vLESyv9VGcDEs9y/PtpB
r1N1FbydGfF//KRO+G1mUgcEkocwDCBQAuS2fZXUf2zLDx0bkjrTmUSWXD0tUxF+
FUEEHlt0LbuFYte+VFy87/eTP+D3L1tT9Cx/xeRc2mRAG7LrKL8x4OxBiUVfQa2q
1BKMwjg3bpZELEmpYYJ1SDiUcdB48TeswjRBbo3LY8KQ85tLgUuG6NJSaCSya5Mx
l0ZkpsjPhcRYZIf3zl+YRWfg9jPgxFN91oiQWZEWThqtf0mVGv8GfPPd2bYoTPZV
NFoMottPaZIHJJtwZSi9a98MJR0FXn6+U/17Vs8r66Gi1JpyPTa0pDEd5ZUa1dP4
lVXKmm5EPp4zdc++R0FCHes+seIldL9bU0rC5+q1phk36rHnCq/2/MDBfjekqiv6
RJqamuu+cPM8Z6cCR3ZDhohTPdtJre1DOmVhOv/Pth38KqMpKgRj6ohhAsHBdFyX
XJS62xbjVxsYudjh+uagd3aG3BdRE3cbi7UEbUT71+uoLTNfnqSN2YQgNq2/MnCo
5CP1G+OGXAWR0jE70VtZralXaTjer2rb9HcaRcOD+Q4+xXIG62HtrZQbsJrNLZno
+Nf6J6W8R9ZWKaKDo37CAgUlWr9Q0QJdQdoFFOcXLOXzCfUSoIQH6fbylOozMzOw
vomAWfalv4GS/zfPtZHYtPrYn4rSfSGA5nsEzvMCl6z9MxYaT/BML88U7+7+17mV
Czti3ZRUg1iEPezeAp2k/NEpVT5XUPk9qrfNPcyr78p3cOwCrHT9qOfpuG1HLrVg
ycngliar5xBo5TkKanYJFL6ibDv0qkO29YDSxOk866JQYL4EJoRNgoR0lXSxLRmL
GZx/fYP/vY7iq3sDYFcRUpK6bUM1hQSr+0GgZO7AsAimZNgSQ1ZQUaUqAk20uEeE
cbL3TUSWE/L8cEPC7v3SMr58IZxZoaUC17a9BwUwH5d9U0UUSU3nnrpSjvfqtqt8
ThvURV0me4LjaW0uS7Kpxog3QYjDfsRumo4bocqqlHYsuZDd8BFLDcH2+UD2jZbJ
Q6sAoP2EYLvBWAv6aT3D6AWsYf9in/SQlmkwL26gU66F0lORvpYZD2mqqQBuZJ91
hOc1IQxvpahxLZgrr9K7VRry+tuFqmv/XcK1yC+/JsfD/QHwdwMm7cdGcimWGHDd
vO9Yj+YMb45yLw1qz1lauCgwYhTXvFXFFRjm/I1nfUIQKJGzvqW/fwvMb55Rz0nW
qXn/N/kRDzSRjOin5xrjeTDPkhLcRwkvFlO9ElYWAd44H/MQBpk4g4f99SZ1ZJs6
S1Lt81bIqerTtJnILerPLae0EILCuPexe45X59z1FseSC0DmDU3idZeKBmQcgrtz
HhG1w/05/xE72d3zO5JVAiMoVYHWwNmJzULUKzrt/vZY8rCR0pXw0nWo9IpQnrpi
LLKDy2BosoRsihnt7hYjlYP8eA0pysAAYj13SozWl6yd0CVuF3zO3CgY2ebprcuJ
p5aX0SCwwRh2Oi4VWruMXbpoR/xRcCg4lUKOaIxGW0uFXpYUGz3MhzjVVtzC1BKW
SBSuYjBh1F3tBNnPk/ASbupICgE7b3SnV94G38sEAHPaAUWndvguH++mhy+HXdkh
1ogl9n7DcqxHmjNspNHKiNoZ3R0xFAx8irPJVSpzOqtGW+A40ws6Pse7B3ZutwxV
Iy/IOkXpnjbbUV8AnCwKyRKOKJZ+br75aGUnzJjwf1TlEQecJOLABrylgS5FJ+HY
i5+ytDX4HqcFsnVrmnUb4qTnx8U0v6jVPHCzHBJt9E5MyhOPRHA3Z3iGv5ipRqhM
BwbCaLJKptaCh7pKcItfYdN9WsYdOmTyQia+r8LyLMZZAsIgmKeiN9SVO5R4vD72
AYu84832vBzcbv5cqN6zdD7l4rhm0JWykFzNF81P6HogBR+QAp66w9E2AdNzKmvI
ruYrghQol/LXR7WR1JwPx2S8qcw6HBCMpISruyKZRUKZRtTOec+e1zP4ck4z7jgf
kGiFUIzasx/Bl+l6Of+Yxyt9VZV1j4RX7Kv4CERWvE0Wc9pCW3WqR4b6cIp2B6jI
UiH+h4dk9M+7F4KACUf/AoKsn+wEmD3tNNCDvz1eGZ4oad+bNwQWW0hMzxeH1Ysq
Xwokiwa3a5fzcnQoJoPye894pFOcDZadwQR7TwGwZyTwyTyTC6GsljRkvxtxAfrv
MXuo/tVn++XR/vYUud57eoo28SnSlb/cWHNHN90Ktt3HCk85YH21YoV9NtSnnRv5
k76Xcu/h0K8zQ3laqwiXC5SaWX61tOdR6FpiI0oK1z2JA/P38wkaj0xTRQlkRSM7
n/9e56Mhn1I9RPSwJgWhhj48Qd4MZRds0pTW53TwHJM=
//pragma protect end_data_block
//pragma protect digest_block
TUVpYLmDclmTp6DvYVMMoKXYt98=
//pragma protect end_digest_block
//pragma protect end_protected

`endif
