
`ifndef GUARD_SVT_AMBA_PERF_BASE_SV
`define GUARD_SVT_AMBA_PERF_BASE_SV
//`include "svt_amba_defines.svi"

/**
  * Class used internally by the VIP to calculate performance. Typically an
  * instance of this class is created by the VIP for each performance metric. At
  * the end of each interval the values of this class are used for
  * checking/reporting as well as updating an instance of svt_amba_perf_rec_base
  * class which stores the performance summary for an interval
  */ 
class svt_amba_perf_calc_base extends `SVT_TRANSACTION_TYPE;

`protected
\SO(+LHU\#B.NRe329X2:\:a.U:&L0d)3.R\aA(V4Pf,HU,dV^RT/)>[ddMLL/B]
9?M,d&,4WO3fMfV+&>_0aADU\D3E_>2NC_JY6c8?OKR]-X0&MW_T<HB-Zg<100a/
g,N=V?]CFYg;Y@=8(W@7V,D.VJ:e5QOdLDggXSQAW?ae7-gDSJ.VQ#e:(:05XS4P
U&Ja8?FWPgdWI57??(5d2^OV;=J^e9d1\(UQ&2e:49?>4HfYcJDH)94L)?\V[.N@
3</&4@,a@K:5FCdgF)R8XcO/XK4RWRK,dV9eCFVUDXHSA0;//8Y_gI5c)b+/5^-S
C:Z@+L_.&U>&g2N.R1YcCb.-d]cC7ZR[TDgPP#>WVB8bQL^5LN_9,BT.\YggUfGg
Z[L9]Q-W)8CH/2dL&P]FODT#</]8F@SFcL.+UUKfN4aAHIAJ\96ef8>MFS@Y6Y9e
<[>Oc#g]cGPcR2-ELaTL,ECb-UV_]#5V+?dO,[WCI5NV#,RX7JUG0c68G=^W9A[<
WH3[g_:S#@^2:P[,S^C7,VS1g;6UcG-OOf2Q@R.E;@37Y.1d8#JH0_C:;DT;H?X?
174B8a?>]I,+3aZWdM^XR=].0\CV7W#JT.4KX/\W55;3QE+=c@_NX7CaWW4;LYM?
(,N<,<5KFU4:bCMZb5UKT:GE1^gHc_]+]/B[-7-d,/&2gBAUPRV?>PFUNN=874,Y
Y&>^,&OK(I)OQd]GVX^:/#C5V8cWS\@[/XL3cS,7gZF(Ab1R1[\[?JcNC_(OITN)
@dXfDU;aM6G0H4XGb9W-R5WJ;-CE\3NW:(d7->NOTTI0U0-79^RdQ.539A4/(&YX
D3S#?@U-NJAc.GJQB,8G/1]]37#?5=9XRLbS(/eP>1B+?]R1XV(aNJ=X6ZRa/LJK
X=9-X;<G_,4bC9,;:bSXUDF/&PODYcY\b8>U;J,3<T2FbcUEG?G1da)KL[@cH<#,
R,U7(L87F6/1E2()Q-@Za=aU3Nf[Z-UWZ6OZ4<3K1Y)+X:SR9)g_5e895NKPb&6F
^[5XE\cZ]cMePE9\;gWaG?+NP@<]T;]V2IXC(KAUg=>22(<?+_e\MH1PE\GWMGI<
cSK#P/fNf4IN/ZZ05>^_e>[=)ZO/^INE]VQ9OH8d#<SXV.7.UV9:2[:fd+ee@-XC
R)J&3B6g]TM;Wb8BKd\X?S#XC&P<a)9K-87>__=gS=<)g/2H=MH^c5VP8BZT&=US
)ZW/cNG;;)5;HMD+>gT>S9b^=f9gP]KJ<BA?C<\c)@RE0WVEP0#F@cE5<>UKfc.A
B9P8YH]TAJgFVW1b_2)g2^(+;OZBHSWA&,:_K8MI&3Z.\e(X/35GF#c^HPA1IG(3
5UC6VCfUBM606GZaW&GaU4?(7LJV;>CFV]UE,_NRK6@Q4C+R9QLX>\R=_UYS]KUf
20a(;O)7T)cO)Q:,WKI&T6U?OJ/=cQUBPKSc/TZ//G-/-^DU\\97aGY/C^VTQ7S[
afR)8YMgIEY0e:>4Ie;OFM_0I@Q67_[^_VIN/BW85,8dQ(A92f71cAF9Hg7cEf,J
PTKEFaG]^_1WadXB(H028W4d;8GZ1-OXBW@QZG0fRVH1C1HW.R8\U;YK6I#WE)K1
\4eCfa9S26baQDMcS5<^U/TNILL\4]95,IQ.QE]H#N:dSMBW<gR_WE>ZbC1>[\BU
1f_O527[.C]C01NgIR.QM\G.EIQ6cd7KSa,^1YM=a@1772(?_MJLMANd<K+[(98V
YDTOU7<R/:HID8QTfgea9E\6EGCE4a<YYY[=J01/X-<&FR(VfP[P.^Y4=baJW]#&
+KGRL^-T36+.,,aP,J1/dU_Y5cYF3=5:M,XcN@T8YS9O1SGE=Pb5.fNU5J7F5<?Q
GGO)V;f>]NH=6X,_adeQ3=LF9VL6:Q4(4N+7U<RgG8BAJ#V=UfGC2:;Nf-a63>@^
Cc[ITVB,E0fOSe8.7\8,]6&W\=^/3H&TV_Bd+4IDKLW2cA12ZIaP=ed?<2Rc3MCT
GdUDQdPUYAKWB7eg2>WM&,CJ;TI<MGIHEX1If,YIGRA,gOIY\1:.)eAOgK4.eBWG
26=XJ53BaA=Z-D>c#aDROU]c:&>M7)^(OW8\0WW0O&>ZC[Z5+8fF+af=5+f8NNeQ
LT84\^O+1=Q_b^8\)]+T7M\<K9#01F</X^,6+NRA^FW#4F\=6:A>8L#4KK3388E/
#>Ea(TV59\JC]WIHF-_?((LAcQ?B9dWJ4BO=[93NNI)Og3)TdI3-J_FdENSBGc)c
CY\/F@3(+D&8EI/40#V;0\)R/V(Yf,d]-PT\gV28YE;dBf_]FV/8b(00B>R/+FZM
-SPR.:D)2TSf-d#><R_#>64&-E;@J:\TE9J7GWI,OeF-D2^TVI4SI6Z6D;gXQ98X
\2QDL84WR))Ja#8HAL2:EGN7[K)OZORU;H93]\Q3&<#\bbKVIgRf^;M._JI.^(0G
XL\SRaLeD+/bUEL#e\Rg@\5@d,a[QO_a.(VPG8UJLXB.JQ17\VG@bJD0a0^+5B(S
?HDb/LeRKePEBMN^&Z_TFZ63+0-UW?6N_U\L>P]IB>d.G+8cYAL);+I2L\DSVKb_
LJTHb1gW1Q:A8aLEVQfQ9X@/]Ag;NK>V=$
`endprotected

endclass

`protected
d_WN.NbQJ1>SL]TSKK;K,f,Y;YXC#OIY@CE>AfLWQ[AZ[g7),aa>&)C(28e;G[c>
Z\Ie&JVI5c4:+cg38]V,+T^:VU7gAYX-A\4Td_^P@g+Y>[55)aO.>)8\+GUcE9c5
eAZ<:+E/99>2?#[&8,S3I&d/<TN6UOC[P&C9aa0g.3dQB;QGG6T?Q_;\(QgRB:c[
&G8X3(_CW6+G0bBLbNN40F_-(.g_fK(?W_d:_CT)[(\)HAZWfK<;g\5g&)B8KJ@&
6550UBE9.]1N20R;6+^IQg0@TCJ(I;20-#fR@Ha>=Y<ZJGf3=IJc1Z6B2-f^/A)@
,GA3SM8@6\d--S6W,Z_2,TG<#V)D+R(AbB)X<?.d>VG(=WKR-<eX;^4,:C0+DWU5
[EX=#K>4f4)ZG7VObdaC0DG58)b?MJ+#@<+2SZX-5W&3aDRd(6Q--R,@=]Y<e\&#
>7K8VI:.>?K&dWMP5aH#dQ<,.I/M[.-+6XO#8808JYIS:>DLC@AcS)L+Cg,<,Me/
K7NYf>;-dfe\EKIT&:_6U5c&NTdU=[dg3+^X]?4Y.B(N_WVINK3Rf+1HZLc,T0V;
9J)_dV:=(9_MPHdbM50NP,]XT.??)9<0YUa9:/TCSMb8SL@MM7d\=N]D4PD.0/F;
/aJc#D2M)\#GSQfc0?X0CZ5\Y<^\cA1fbf+#4C4af^Q3IfK^LDUW4YZJ]Ud9_#CA
@<T5.17I@6.MLN:=_MCO9Tbc=4)F@]</UegR^+NCNSZ>43J]TR@=H.L<.O6>b6^2
-+Iag&ga7\B[X&(eQJRC,T^a0E>Qa.IHDBgaI7<T,bCT\U<W7D0R/d6HW07.SZ#f
\WNG;]D;9^EAc+A4N&-J9&c:D-I/B:[Hc#T7cDQ8LU,RZ#NNH2&Y:&<N3MB;/P>>
7+a3W#^]RIJ99P_^08R+-?C^d3D?@69?XD7,(UKaPDb.-M\Deg[bX)DOMQ+(JUC@
)W#cc4?53S,,LI>a]50XV\>cKJc4N0B^g[B-GP^]Z/)N+G-H2<)-CU1UV+b8ACD_
4CV#-.I;MW2.-UVf\gC<(@4DL^XR/G>K,\W4&#5UDE,0\A6D:=7P17-V2Lg3HIGI
dVOB-cRV[[G+bPWBGPfV-LP6]8)AO[^KQ\-R8&X;<]GW8_cSC\eXU1.Fe(D/ZJ\Z
6IcDH0[<+FJ2(5IG^01=R@3c<XKa7(?D/_]aN8;91.G)gK3EgUE4D/+aL/b]^995
1,KC.e6FJ]Fd;eB1=&8SNQ2L+O];16/Y/:7G=W^LOLTQ1b9=/)G2P_+2a/8MD,BI
Pe^,ZABB][+C,V:I?N&R;<Q918?O1BeP=Y1P/5I((=#T^KQI+ZXDAX9(N90VL^\(
BSR4,IJ\\-&:Cb2AZ<KV79.7,7=C=&638;SKDIb@W[8,7GMZ@d0IE^PSHH=?JP.Y
O)c]fCQ;2P(Y/A2Q59M:gP7Fc+7fC)HB@:FDBA_6TA<cH<Dfg/;0/S_Qe\a^_Z0E
3Z0PB.dV-FaX;&S]L,4#E-8B=K(THGF04Tg[GU6YJ(OOg5D+5)fgYX?e1?1E/G=S
<Q-/(C<>J1-JN/7IC7R\/RZ_)Q1L@#Ac^/B]NZVKO]b^3/DYDK;WA,1_5;/(6ea6
O-Y^9<PbCf,Z7#E?:=77JIUQc)SZb+I00@AHOW/B5+3AC5+?EC\]7CFfL(,UM:W[
G>F.);2-dDT0SdS6@C0NR#,VSf1)XV/HZ];P#d()fdQeP,JA5G,0&Y#?-^JU)T(]
)0N4XOR1,O?:/bLUV5@Nc2>(H,>&[&L+KFXQVQ0D5N2NGNELcYC/,V3M@_=aM>]V
=e:T?SZV6WF#-^;/Wf[AEH::T4-.ZIV2cW\RIANg(-<\WC?0J#:=KE=9T71HQOM?
<g0,ECO4g:-HRT&d1I_PW-+V;1N__(\=<;e_9gF\./#,7GEcDH-#SF=?\#fJ)Tg&
O[HYO>U^[OGM(NBX50b:S0?O:&VZL:aTRG3TbA(,)d@\7bYBI5,:fc/IZ?XBNR[E
S]2VC?b,-4;X9DKe_CL@e/fGf.O-CeZfJ6_5S<a>2CY:P#TR--,9]/3dI7d&0e_W
5S_-I4#H?[P;,A(OR0#]@4V<De]ZK+S)Q8UFbaG?g>Y9eS40IDGIPgQ:W,ObEQbG
BC+,^PYA-B0W;2;[8++C#4(2JPC]/8LeM.d_M>RS+\<BRN<T(IH>&5D075g6=M==
^gWd571+@;B=?WU/P:,Q.DLH04)_]ZR;(C,4fJYTMZ)<@IVg_9@KWR[(RbS]6#a>
9;ZC75.W+f4eOC;b>F;RGbe9W5=M\>FYBL-I4a>6@dFcHfM6)[D</]-DQ]PE3:3G
INI<<YIgTWd?+4WVG)-O4^7YCE^T#SKAXOXW4K<O2XfENI1aOS\D/E?9?SU9+1]?
f4&fQVR2Te\RBBM[Ya&VaN3#GSVY#a4a6KeJHH8bIL.)6g_/+N6bC>@CA;XX7,3<
/@)Y4&PfTVNRS0H(-KR@ae96Ia2gG2U(YU>7K<Mbf,0\F6b]\4gg]G^ZLD&T4/;@
=UV=XX02UJAI?8UN5;:C).[5V;3ECZVG#@gC<ZY5_;_0_EESa6B]JNP3FI,F:)a[
CbUG4R8;Gf?bPJ8U9E/fTI=<H.0,,/eKCd9;6I1&4_:_]3N.cfDV^)5dYBSP#d+g
fVM(D=Ef==6IG59&^@KO]NO5#,^24/g[K9^<V]+?.85<LN9dGfPg#+JaT\g+KT4H
J-:[L;GcYG?7+>58<RANS>^d\ARV4ZfV(X,SGUC-^bZbQRd?/gN?Q.gb/>2<=2ES
(.1DV]GdS6KYOEDKfWL6:#I.A4H=#7E]PH>MD(^&Z9CXS_FA(K&-=b/(>W9c/0NM
59^)2X&QJ9f-bVFWR8&1ZLI.5$
`endprotected

/**
  * This class records the performance activity in a given performance interval.
  * Typcially, an instance of this class is created at the end of each
  * performance interval configured by the user and is updated with the
  * performance results for that period. This is stored by the monitor for
  * reporting
  */
class svt_amba_perf_rec_base extends `SVT_TRANSACTION_TYPE;
`protected
7/2c6eGSaF8,C.TOW\F2IQ@WMR:=)g_WVg-TX:#PLQ&W&dfc4,f,,)6f0)&EX3S\
cOUb)Je,(1aNQFF+WJ>/ZaDB.eK>EA?&)X1I[G&52.H[CBR3RJFX\A?(-?H(?H7^
gUSUOSDWIdG.e=AcI8NfSU?W6f#S93-/HWTCb6QMV<c-_e/[GV3N8M#\BL^HXSP(
d^SAG]Q:(,g;)ZF;INgS\fD]/5UXdX6U?/f7M5Q&31/LF-2cdBBKB[I]+/CI<L0<
<:,f[&3b=_XgObHF4UG6Y]D8E5A17[Q#VY\E/?HT#7+>9M;#E<VW2-A]LK5&W:[L
IX=KEX@978O/O90EE#^KSD9<OBU\_6\79^fY081JBGAaI>[>(cZ;U,=3b;I;W8D0
\R)N9d53Q?Id?1A#g[SZGdA2+(ec=3:-DKGW>f^A/6^W(>V;;L[gB.;WIBVdFBFc
_-X2]U-Hb+c,#dd\[G7JH3b7(FHX/0X04;@BMJER=#R8&UGGMX:A12D^<O/66#&A
>@Yc447+H[06B3eMK5YSg4+[>S+BJ:=N,OJ_-1XV8,B+_/KSdCKfKNgMRV6G]TZN
H-OGe_JLV9c:TEUJJ^WdN5d^/_;a2C]V\664KTPC<-aLQ2[)+Q<35P,EPL4gWNA9
93+@6^.3@/Q4fJO/d.cM2_g#GR)0HJeD/RQ#ZK?ff.]H-S2T0RKW,48aUWS9LUfc
BcYH6NM2CfA6UET98UXa@Jd4?fQTT\P_&HaH_e-J>bFVG<#SJ#?P?0MBG-V&P,FN
Q4&:A:4c]_-b)E_T31]eN/,PS[O7@5@8F<0??c[WN#5Q/.JWec(\\a2bB8#+6H+7
:+@,7C7W0>7\\Z1E(ONF<.99.71;E;^B)^IVJfYVLc/]cF&1K;0.Z6gB\+/Pc3YE
af>?1M=.:^/H=NCG3JJSEBa64b+3Y^T?ZBa^]3&dYS(=<5=_;#.]Fb?0)4>2T/b2
T/ZfZL3C>V5[HWT)E(4>6>#M4Rcb5VfROMV5P0XfcRfNW]KO/?g5X<e/ebSWb/1N
cc_6V;gbP12c8_@I34S31GMCee&fNDEC_/Pf)8BTHcN+1D6aL,cV-U3#89dVFOBT
80AB>K(F]H=I]GLa1GI>Z>-[Y7R0J52[&,OeTaYb?=LdWDe5ZA?5)WL4^e,&E0K&
;WQXHZCD#9e>B\#.d>4^\S;Y&<D87>B+Wf@XO[\7:QZMa4G]aa>XTE?c0bZ+Ec:E
>WK1G7:MXS@d/.A7=LQKeUL0bIX(3RWeD/a^.X;NY,J63DT9S@AJ]Z0.GLTa1O1<
@e3V<VVC+(@VJ.(HG,HcRTRW6;60#GHgR+)fP44MKL.>3HT55I@Q\/e/X>>Y@R(J
(;7]S#Tcg330Y0Z>@)[37MbL;A_L-(JVMY^e(c,0Kb3FJ7CI(H8DIfJ1]>gYP(0+
f#8cK>/KP+1AL,T07=F/W.c4V)[\,7D-;<TdG&0/Q#:Q8g6I(M-S15LISE9)_E(Y
>6HaI6K.gJ3a,=5FDYg+)dKQB\NfKH,c]/XJO\6FX(:^T8#8Q23VV]3ZYePb_SSE
Af>;G2Bg\DD#THOLQE:BZP+A8FF&ENVLK^CGZb,(()YST?c)&Z.R;ac;+1e7DOTD
>[Sb=eI,bX5.A3X7ASN6PL--,;9?;1O+J@JASLEABBS6VVfFM_H4P-GVGG/>PR_+
dZ6W?N+J>]^&:DQ5B@C&61M1D@IY?ABc?SASe>GBL2-U-bD(G5&GD,(G)+b:NRZ5
R>DF24J>:+:]dcW0=YA0P?5a((<)G&O,VWCD[I+=?[CXG)g,V>gd(f8cFTJI-7UW
EEDO>O2NCYTSA3(#/=-(8(Q1R<_MQ\HT9fNO1^\:2Qae5G[G:5Qa:^N2Kf+2IR4R
dI)NRNB2WeIC7ADWf2.a(YF^a0&#4]/NINDM[X[c>+@2Vde#C]5SXS_IWU1)C^W2
X.;27,)47+OaD]@.2Pd(:P9g^1V9]9cDdF/-2JdCfS;RYIZ)3L3R0ONKR8<8+dN,
cNcOTQf<3cd4(6)fX6O)97^?B_e1:,dY_c/KK-aZRZS1<]O2N<;TCA,g)LE?f3Le
dMKaFcaHT?;Ee)f?4E)EcNe@T3D1<8/5F2N74M_P:HLX9AM6bNV[JRGc=ML;Y\+Y
OMBOYH^]]dE]P3&Uaf^UQ#;[=NFT&TA4f&dc:W(_B[(fH3WeB(Mg/FNKYeggUGKK
FE3f-IKAX.,E[++>2>1c/gJ;Z-fgR@EJ/P9]E:P98aF-C8YH9b2W&5)6A)];+6:b
/B5b+/a/V/@,gGW6IJQdHXe9@>,gMK2DLRcV[QOaN2EJTJg4?Z68FKK15\F@_XSE
,Fg3XA)#c_Y1VUBe7Y/JU=J]QR/>c7X9c9Z,L;[#X5/fWaFP)b7#W6+\_/J/(<Kg
HCH/d.;cV)3_++7d>O].a/W[f-I1F6[MTY@3B?<c9e;4A#O4HbJZb;SaI=;S6D0c
W+9aZ)+=Ade-BHOR(;@]G:fYAA,GNdROM<7[ZGeT5^(]6@N/_.6.Y?58_(/1]Y,W
FZe4HOIRNFS.A_(FF+a<Y:&81HS\>a8[E1JbMg>9IOQ65&Y7J+Za7VF4d(MZHY)F
&X0T\H,d[VB2<gdV,8g6Wg9)H1+V))>HT&9Q9<Q4]IL\3KgQQBLCUNY=-)<I-8:#
Ue4)F6>6Vf9V<fB?O)>:aTDK,592GdcII#A+^E<LOMQH\_FQ/F4,98&VJ(@ZAaL9
.7.WE#48c>8W]M]40YZQ;V/?Cf:&,b01<fDR5g9eIGTA=(5LdZA6P.,]dK):@gdA
-f;dLHX[cFIGJ?O&bOCGUT=:<FaR\U3dfVc:=QE[deSQITLfcO,4YIdY1eS1-4H<
E:g,RF67+E/aX/D<JZUd]5@P)-LHBIgCJ+\ZbXDbFSbAC;2,a9D?UL=W:+48EI1A
f;M0#D7LQB6LaM)5GVTKI5^4G4#1:MM:9d<^RNg>^=20V_-CR_U]A)VD_Y2e;?>Z
ca74V+;V@5&e\[EV\7d,:29E;T70@V]c]eV1ZFL4L6V\,FK>d1?^2IfD>F1RcI/G
U0Q<_L8^S=(ETD@WLAS/UFc[^<(@QUEQ3c+#ACBJK#g3<c9OZC[9eDgD=16:fBe^
#^,8cQ8:D_UA?)O)RF=QJMR)O>c)U2UPfQ,/5H/O0.g?7fcA_+=bC982WQF6aDB,
Z08bLN8.-3F[MXT4dS:Y@d00?M5Hc;fWHg==ZZ)[XT=L=5).N^(:/aeZ^&K0LDLG
&=\c&?OOE^/^<<dU2]H.e<MD;?,\@Ig)OTc7Kcd/<PLV&>[#1T1>fF\bMV#C581:
9+&S<-XSPD4<UaJ>EP]F&JNB12\#4,a6,>ALP^N3;W&L:CXZ3##FHC1WO#V\/TJN
U\,X+B3M2R6&=<G0V>O:fC8V=G+YIY.J1[VPPL)dY\3d,VcDZOQS+1-4EUS[>LOI
KXb-#)NH)P2bKF_<bgXNF_U6(U^FA=,e1b3&LAPe,?,KH?MVKgRLc]6D<S12gIWg
/G95AQb]FBH5Q:@,U3T/&&>^JbeLgNY=K3,1Z3V>7PW](S4;PW(JDc2YNL_N?S48
a[=[T\f1ZR;&PEWaMN/d6LW39&)4d6TV.d4NHY>>WI[_1\WM_:<N28(>a5U=.(J;
dL<Je1b3-c;;/UJ1B_a_e>V)88cfM5a,QF<-T4#;5b4.+8VH:]K_D.4UYB-WTIDH
3_6J0?9AO[HHZ(8DVVXc)RODPJ>K?8VDH8a07\GR9LQZMbaV&2@6QFIX98T91&IU
O>-<S9ea.E,(_X#V[/E>+8::QB[@<Y.#-&<K/0DbLdK0>Z:eg>LM@;#&&+8;#6H8
A>1#(Z\5<MOdV<@+TS<0UM=:-JN3,1?Zd5934I\[Cd/2f3@-L<D<aT[A+)d755DJ
LR=F3UU]./04P2&[A(2U]?>[>eB2b@Ka0G?5dJ]a&C/#2E9Q@9#DXX4C0:g>2(]?
d[b7dK;8(J)UdZfa5,904T92/=NSeXb/-<a@#^NK[(JF:-IcVU7(ML(@E.&9:\e^
W^8]1ZT57HY))BQ]4-<OELYd#Sg2W2I_MDBCY#:_>7D9bD4>V6HQN\TTPTM/LKdT
R^_bc5FVf=ITbPcUPVgD;LI86O.P)ZM:f5]7=cb/CXGUA&NLZ7V5(&7c&_A4fBDg
UP(<5=JGXX&TTT4DNE.R(XN;;JW^(V(M^/R[[H>>7#<Gg=.B>b^@^g/XGQ?G63QU
M8CeX3#NB,gAFV5:K&MK<9>DHC,b+6U:;=9ZJ<Pd]EIM1\(H@Mf#Cd9,^f,aU<J1
-aYQQ;1Kc+CFTU)CQ>1(AZQ57Q)gWC6DSG34:bI@4gSLZ+9(K#R:Y;\.GCaE4:K6
1WFHb&O-.@]/:JPDWA:Z&Bc8VE;[IAdL<_(HB,aCV]+[Q2\,:Le25M)B=XLN02]5
Ya:+bFH_6,VLY#[-a@NaB<NH3RU1;,1U5K=1@-8D#4aP)6W9Q+#__MR4Q/f[B\eL
VQ=H]cKZ&QRE2#J3=.#OV?MU2B.#)fbR7USOMcgZF[#96^D-A-g2QSXA2Y6a2C<-
,ReWb=9ORJ,]C[UM#cf70:>Eb]3?R(JZ\?.D1dPcY_/00XKJ.RGLR/)b+^(RUYIU
?\PW=AEJ7-2BfO,;e,VcHM,XL(fMaY4HLBS;,1VJC0;)_XMEBC/gScLO^A@PNdZQ
\J,_U+1EOG9_RIKgY_9S#QCQ>0#]AYBBOM],U9T/1U5(f[<FGS=9:I<CcdI<I7@H
P)_dAI56dH79LF1G]+dd[=cR\CCHXa?;c>aXKaWE#aU\VDd>7BL^WTbVdH24.g2^
W9X3I1L&6TcC-JF=ABLdCW;&#H[NWNR^?^9,cN?;/\GI\9L0.V=dDS(6^bWJVD7_
:MdP0GJ_P5A3Cd-LEXMVGcW/7AM=\1]L#3@DeD]IW>:6CV)Fb5Za0WKCfCbN_4@-
g1NdcVKL_+a1#e92^F,If9F>ZP=E5&-95O-0/[]XX)L?KK_NS:I[3:(>A5-AR]18
9:#:Pcd.]D=T,&W/3bQ4LM?CIg4=PMRMJMMM^(GQ;d80,0W76KS).(Z68^=7P&\S
YM-R>6Wc8aX2H?f&9K028OM-/.BgY_a)=VcB&SWc3WAHI,9/CVIfO-<O;9HOc)1f
RBP9,4[)5dUNcd/e,FN^L/5=,07I?.1.WQ?Z9;d[1VTf0LY3\\6)ELMEdZL909&f
4>@[f3LP8HXU&c@db&\C8Df\5EdfF-cX7ORQ/7CH,S(3@6g#[5L6IP3T-[OO93)b
L?B3^-<CQ:A(83>ZIdQaUNSVO0U?bK)3HIg=YDc6[62Q^9ZS;I[RT\6RM(.FE@<H
Fd1WX=4bQC(A<4)C]PDG9(2I]-)7_e:2I,R7Kg).H-I3fE8JAX80_Z&PP943a\D1
>_UK37.V=3cMMe.8eR1;FL<D-^3^YI.\Q]GD>Z>4.L<W4R2#d]?7.#>V6+[O-I^Y
W5\[;P06#KRJHK(J@:Ye2Me:-edZCZ7T/e5FXT</F^;.:<9<43L4c&A\160&,XfB
CQRXKD,7J_HLgGbPXV<R6AHKWR[5.4C3_LBJ3EJ(W_O,bZdg8:IIf316YN?XZfHB
fLUH@E\.B^4dWZ33NR+58dZ@5G9/0ce=STPRe2MTCTN6\-E>MQL.7\TH_JB&bN&.
RN8A>2QAd]Ng+2)U4_Y-a.e>,^->Pf-]KN#e=ZSN@A,cE[R]Ye-KO8TX>[-5K4Mf
VQ@NbUgYR?9MH&[Q9\[PO66BJ9:&&IPd)O=6X778>cET\=?=Uc/;JdP]+J5-G0LD
CL</L\LEH#UgO^PP#0S0\f^)(7ZS^A3:TUN9=7>?MT+9C4)[HM_H<e5?Xb@7Yc\F
AfIJ(agBKDUa)IM464GO=-H;DDg?DU&YE4ZG(_2(Y)[:X.aFLdE5;95e_=M0.0,U
RV]Q4[N(@__&#KC.cX48E;-K@9=RWVL.?1a[&Q1fCS+NdNB]2:,\H+W(BX#+GI,a
&0R(B[MX\RdU8>O<UGO:=L^<EaN<aTAFHb0G>CUf,#8+=G7f]e(/7SN&^G=]JUaA
g0[EFBK41f6S9/81:C@3HgN6\eT<U8LeVU<3.BZJ,L(C3YJSGg^,_Z4WF0Ee0K<.
LA7H>Z,eE6]AJQ0AS(Kc0DG@1BgZcV,SB5+JNDg(?aEB1QcEW;eCABZUcfaPaPD6
DUO>Z.3K(N;7_>XJNXPb,HAS=Z4&HW=9N+0B;<74O.2JI9#&3WS=e2<gVY6gSD</
c4+1Pc3U48Q=]Z2XBH345G=bFUT>EbIF8(YMA#?,Hb3[=(E.eSW<];]H[[T)LIE_
2CNNNG7bLQTC&CC<U?#bg,c]QT\)8C6C9f)H,<]5G?IS@-N7SC#cAPOJf_-01X.F
KNc0]>HE=+RXIS3V1RP-<^C]YBW]?,M#H&MI9#(;4C,G8:Y(c)6FJL&ZgESU87IW
gR]_e?CaJ-[R.DJ7)cKU&;c7ZJZ>1eQ=[2VW&6?FT[,6JHS-DDMgQ1C=e._NODYd
dJU=/GPde(IaB<J3VIEf(OFZ@1Y3/E^KT<Ndd(?^R>#STO0<7>0PS6b^,35g]Nb\
_77/D=EPFZd23G+SdA(C?0U6WE3O[#fH/b?;>N;HPKdeK6PT;bW.\gg&UB9IL.[6
f4@=M-<;5Db^7&9a&=C3P\?eJ4Ig,/^NO;HW=U0(cJcJe\BQ;#):bZ.E9IC]B@]H
.HWd@>7NKe+1]W9E#-cM)cC[/Z:d1_I)g1SX7?CLCaK3Z[(YAM-g3]=;3GL6QN1)
0N@<D5-J6BTDK3,_S<XL@OU7+\T8;aHf9#A&c+?Q6W1^M)]a]9E?WSZ,-D^;:KI-
]aB&3afgIL_c\B7W8@Z9G00W=_2YX4dIN=QLM.dZdYLCd3UMd)O>Y<fb&UQ7UU\W
9ObNFG#>ZMW0-0N<77\LN[=8daF@-2(A<86V5^:EI[N-^FL<87J+55S@R.Y?F<RX
=GZ:Z8X+[D9Xb?gW#5;Q9CSG?dRU+L&/B-?[B#S6de(>TgbB&;0[.2E[1K#gS4HXS$
`endprotected

endclass

`protected
agHHJ)D\8c])&RN#>97;_JeTg/:\]AT+/?U-Q[#X;O@H>EDV7((83)M:fG^I<Z@F
0(6]Be@PD8T-b[53>Mf7VGDWLTA_I1),g=gEE91O@c^RU5^0cJK&;QCX-3dAgcO;
OMYSOEAN^ZWHJZgLZ4@([d]6SH4Z,8.]Dg#/bV^Y1)1JRd/6ZWP7DM.bgNB;G=49
K^/cM8dD:?G3/d>/J@\1S=GXbca]/fXR>0/W>51R+]X0)O&:PP5aVBELDdC\(bKU
(:+ZJ\HP-8DbWJ1F87_2T]C9V+SBf=MRL+K/Y(PYHJ_[9XWfF_7J2RFb?R<BG-c1
Ic;826U,HB(+]39)CKO39OR+G&RbgK+@+I/2LI^96dBCUIaaU&>#ZV\A76H9O#O,
Uc5:?g2.]a/2K\][SY6-2?I8bV<RXXd2&LQ/Tcc,51:eH_N6T]=,?1-CJ(?JKE4E
,4LMaMc,TGA[<F@.3/VMT7]TTS(9,HT>;Zg,4?>:P&5dBK>g3E/:?ff,g_&;\HZQ
5^g@\GF=-YWFYW^_I1[gX]X.>B?=SOZ@K[VQV79@c\f3.d2C<d8f3^WeY>&R.Tb0
T/<#Q;V=+^AN2_d]SG&1]IL6:+7F-H0WOdS<MD#+94(<7Nda84&,+_N:QVdZK>@3
0aN=fb5H6_^[VU&@H4;7OHg#>dYa<fD);M,7fS#8TZEKRg,1,E(Qf6YU\\)O^I1A
Be9dVX8P]dB\@df=P=CKVI+T=[^W<7AKS^AH8N[SHGS\DSZMYcF;I#3OQ-G9a9[;
A=/?R:(LZc.K7TOCE^AcW0W(R_/PVAgD1&BCb0Y8QC.YKSE_GZQN?]:B0e=?#0d-
1^Z3^@;,JU[ceUCOW1[7[@[U+b.KL;IdK,KL5IEJ&79:+EN\3HgL2YJ6C5LEXQMZ
]M0W)0WYe,&KBV(_H,NagKIIca2PU2XQ==^f#,W@MYI1DB;GR2>2X;2;2[_O&V:d
aDf^5CK)<Z1S4VB#_JgZa]@&0P&g+>Fg,(ZW:NL]#D+gGaQ0CRFO]V^6W>GKaF>F
,Y07,;<7>8I^9/THMc_3]KSS2GCMA<46+JD?XVPUL,B@d(_gg106C-__9<?F/g;<
f8;+_3M3;ad:P-Ic+3WD\NdX@Z&f6UY\=S(E_H&\\TX<eAS?\GbRK:eUe:gd].QC
+R,Y7_6Y/;U,Q=;LM[\>LJeGG^W#,3S7ae/g(cg<ITKTX-Vb#+ZVL@EEE[HWS((Y
B6+]FVY@aEf(<If58XJ0c0C3=;>GdT?0f9O7[aC+X;V/BBX33Fb6FgEfZc6WQ40(
11^-;b>(Q4V4990TT^4Z8gJ#C62^ggL&+TAcK3d):+99II[T[c,BRK2^^/fA\]Pc
?=B[Z1&(UV8F#:X[4]CQb)R1dX5D6I6;_=##+=L:.MQIOI^g=W8DBGV/AQO1GWIQ
A?a4d5067Cc4RHgCb5\;87;T[VYNJE\GW>L+CX&EM=V2:9U7CLT6M@ZGFU[[,/fa
dc?f+GPfEYGF>=7S7fIP?FAU?)R/eR?ecG>fC#K#/6Fe3#a/5@-ePTX=::I@7J00
70IEZ.C)_NY@,W?)#:IJQND/HB]0#cU.-Y<(AW.ZM90I9G:3,\5:2(WR.(6P0.8,
)1)5;=I&UE5I;EZfe:cBYPO=575D.E=\P][G#@[@=aS1e3Z.Q6=SG-[32ELP5MQ8
[[1>N(UI/aWUe=>?8eCc8</Z-JICYF0cFCWUD\g<?d->1,,g.4He0<9d8(C00_,>
DS>NZ=2U,=a;SBZ64O/NQ/IV<39J8_J?YbSZ2:S713.L/df(/Y8R?a6I)B(=d6^:
.HD4b_P=E8E8/[2,R.=./fRX3a-?IeN7U/g@MXUZS8U</eMN4A\+=CA:,,P?C]Bf
9B4)XU\]HDe0W>O3@WB6Y\5.3\1Fd>>_5SHR;eRd\FdD:RcDY0I8HJE(-5XbfRe(
.#8L5FL^ML&gG@TDTZ[VX4\H):\g+/:]X.^#GQ=8;N52HQ@#<+E1WG6+@DFN#N6;
KP_M_R^#6=\>.EY8e58#;,<=@\0;^g=5LQGA_Z?Q^LXV:.LXWJ]2AT)W8G/_U]-T
)8+..&/78=R;@Z99eL;,VDg[6@]78I6]1R)#AQZ.^F_W74VAb3a,O/#U_?N-;_MB
=UO/b&;1=;@5T<TG(9Ygb0PB\SRQ-A4HVCZ/dYKfLI5NZ^L[OD2-K]7A76d:]:?,
13<./&^XL.E?53eM]>KFY?-HED>ZW)W(@A/3YC&9c7?>3#M;?D&R&\#REV]_)fe6
B=KT=[0gFXQR:E;N5b;?KT#1:=S@fF,).>6LLIW=17((ODO_eL5X;CO_aO_6TU5Y
BRCUL;B=[-,S;IV6?)H=?TAd^^]?Jg,_f7.)V63C0X<6(^Q[g=<aae+5B_\\S4+:
A_aeT>X>M<+MZ02[=@WD+(RX;0e.K=e4cXY.R,3bR8<,2MFBGMX)2^\(E4a+B.01
INMR1X>8U7W)b9LU)GT]NB\57TYBLbN,<9-N+\61\a5d=0(&1c_Q.1=B9T(1F\Q=
3LdMNUSQUNF64;ASCdbZ-bZ3Oe>TWM3?0P^YN7N.,C]aLb[TT]N8T&9;DgY9HJg[
8X>Hb[&CRCE;XP+R,KCX?VH,M68AHW^E#XXNW;c].PW0X1/#MHW/V6@gLO?.f3,,
IYL<]24AEL>@V#3Be5F8:fIc;9IIb^bTWW=R09L-^1BKdI^d@8BL-O>?I\Eg06@R
9f)K7XV+L-O=a[8SXXB);4SgNY:,4:/HP8HMM]g4S(XE#Z(RRdSc_HBH(Y=X93^I
2eWVBW9/VK^7gM^DV;XNS))#S;\K^Kc/1bTC^ZGO9P2(,Jb0Fc^@XfHc&FT5TLYR
=:71]#TY[<TT)4fXLa-/6,3]TdNHb@=C:d.MZ)dG4[(.K:0@J=-g@6gLWN-afS&d
NL5>:2:]X40Ve,PDbZ-e4c(:288EY=4+4TD:E8&N\[()CA:^N8:CQ<S9XUCMa0=4
<M0@X^^VA@bB9,M5bBc2K<TITO;B]B)=15egJ2K@R5aS=G@A9[&CGD3SR\=0GDa5
TN2f;,8VPT3V/VUbNY][LREH)>S<5PaTNY-[LfCb)cE.c]?NF4Q@YbTSS#3)6@gc
\e=7IQ]O-E:A6P9K[&(0N?7XRO1.+d[-#QRA88<?A-O:,.R_KJUc2?=;S[c+2JfS
4bH5YDDaX,fTI=Eg?LN1.@7X6$
`endprotected

`endif

