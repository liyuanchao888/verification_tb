
`ifndef GUARD_SVT_AXI_SLAVE_CMD_ASSISTANT_OVM_SV
`define GUARD_SVT_AXI_SLAVE_CMD_ASSISTANT_OVM_SV

// =============================================================================
/**
 * Extends the base OVM command assistant to customize it for the AXI Slave
 * Driver.
 */
class svt_axi_slave_cmd_assistant extends svt_ovm_cmd_assistant;

`protected
8UTPg,VJ),Z>;9<=9g1(#3#;a(8<LeY;U=?NC1.&4E\d;.VCgF.53)8L+28U\0BN
K0NbFHD5KU/_LJICT0:.Ke-ZQOaeO+4dVTE9d(3=(_(9Qd8;PdZC)CeO654EWIE.
+)T9e2c@aA]#e-2;^c;L#?+]c/;-CgcQ:aG/,b;>XEQc28(41;fZXSZVA2_ATH)[
N=5&BIQ&5gD-R)V].GK]BGF(aW)I-5DW1)19O].:7CeSd8FgRK.g#dBNPVd[[^LK
<;)N?OUVH3cG+c(0XFB^J+@:HX3:@J14@MF_4F,DZ^0:ZX]\3,G-_65HVJWND8J,
C1(Y1IcK@U86P)c&4#2S[Q3KIF.g/Y]1c:>1,::8I:8Q-\>JL1dbT]cMI^dCK<Nf
2e67065XMR\2HQ_]0C.f[3b#^_(f@&,P4.67UWdSc_R+Q:7A-c]dGYS3Pg_00fZ8
ASQHFFf>\>5EA.KHC;94YPEDSP@b]W2ZN_V9SdeJ;N]1Sd_I=;)UI,YKT2;a^JV[
Q<Kd/4a1.6]9S1N1_W,gKAfLg\8&CbG9Q_K#L9+]#Md]Gc7:[^TY-5BScZ.8LeaN
HH[V@FYN>7]DCb#)S;<2/cP(c=SPD@S3HQPZ]cfDO<F=RMWQ#bT2?FA00;^HY8UX
JS/E?M4GJGTYHVXMN80]MDJcLH+:0QU,D</_(A)?QaQc?aDa)P)M^8H8B;UF+GX>
90F0dE0Y;D:YN(1aV+Y#&?K0NY^<3EX(4D\.WH5/.bR]-a;\G2@CL1Q>@8#<P&?,
(B_Y.e[MHfOdNQ\ZW+^Xd,<WCWg6g1fc:@-=Y\=B@&,8_f)3>;/&Z(87bU^=GaAf
&(@cOaY+6+e)@H0P<Na,T6<W8$
`endprotected


endclass

`protected
^1GaHO5G?F-dPN\&=Q9Cg<R9dB/9NTcIH9,Xff423Lf@B<1Z5=OU2)dD[bMTG=a>
N93gNRIb2]=JdR+0K64(OC.G0DU4DDR?4[4TcAT.HG88GQLFGITGT+DHNP];.^U&
S1I[K84eI10d;cc:W[B0^Me\?E-IYS9T4\g_4QeeL&a@Q8<X\;MEH7IS-XN12PF?
].Yeg6XWJK;-G&9O,W_f@QD3aa+4_KDQJ19[L-Ef7#QcXT#6UCWa#G055SE(N<PJ
<GPKO&=N(75dEH9=0[4#f&eU[Z5D/f=:<D9aH:d<_H4Eb+@F:B_#XTJJ4&=16TJ9
8eSfS::X)1_GIC,910NN/J^MfKY@_]a1&OI/KXLcEO[T22:Tcf_EJc-8-MAGQ,3C
K^XVPHJ&b?LMU>aU7>A6&@WN](VR:+d:OR:g.=:^GD:I5aQ;/)QP[,ZC/[MM]Q8P
;9U)#CCNKc(EAB-Q>4@@_/2VfMeK@_2@7+gGY_38<>dA>&1V?O_O=K1<^9e[8b.C
A48:ZI9_VC8:DDLI[K-(SG03RZ9--eE^e(Pa/I:D]X4P<J-fE&W?@VbXDX^PMOc[
_e/UXONY,55_>T2+Ga4@QbO&&J^^V(=bdC-YN^DNEM3B.N[g4a5_L.QASN8_QL=]
BQR1PVd<&362TPRR4GL\6D7?,K@ZX@fMe]PZR3b29@8F\c(eRPgA2b78.0;P+ZNL
KZg]C0f4L&;9@ERJ;6,bV)\-VVHfIK)_(U:?Yg\3R3,Z?7P=JPcFK.8(f2);Q93M
WP&<#(_2aZH>e:GIdR76EV&V3.FD-(12VJPI5U>IW)D9CA7V\38dgUWC&:U_^W6X
\E19MW(cCPCO?YfWKGM+=(R-V-?4dGE;_TK6TNPG1OaZ78Cd/Y#Ue8f&.>gF=+D3
IE1Y\RL#EfFV@&UV.E?WJ:C[@W4:2+N6CE4CdJA=c1M1GAT8=/@]SCVG4.f43F=O
7Z?FUbg^7)df09J\28;6SO6BMXE0Cd3DD7ONN^T?@+V/^10WU^4g/LSMHJC3MRAQ
5)+/g4aUMWeD+fGd:=KC71O;gFaU3,@8<Z8g(RNWA_a&X<<?L+#:(X_ed_9JIA#3
Lb4&;Ne\VVC=^1d>6/PSMF1PRMC=QX7CZ:FU><VdfCCe7EQ>/37[+R(T(9+Ta--F
a&XXB\,g<A4[)\77;>WRb<<WOO,_X9^BGS8I-Y49+F/9LUH4&T>Q2];?\XePE@R>
g_c_GK[69)c70R3Z1<4Qd72R]<J706_=/4REITJQ(,[fN-b]<_Z6fQ^EY]ZJ<<E5
;+YB>;Z9&(_.Q_&c.<W?O[BY3WRNe]VC>2N@:Y;YSIeV5:TbMc)LPW@-aMP6fDU]
H]be:>]Qe&H?M5+aGXITE9eQ8OP@fQOUGW@40d\>>Q?K/>(6I/9W]C7?[-80^2dY
5JN^GW1O_5(4GI>e8@JcL>)eC7cdU=?USALEJ2G<5X/KQ^ZOZLI5DQ&RJ:F(0T?]
L>,(:+[KWU=bU=\.@;g[3R(FT#?X76c7bQU>e750VQ84_X]]?eBUaZO)R6,O6:dH
+dX5GKDegP:VG].42:Y#[9AK1EHecDQT@gdcFg4NWN+g&#gLQL4Kf-CFX11cK_PJ
L0081R@78XSM,Z^##H[[K3/Q7>9;.TY4PW_7RP/]_OR>+g=^)&D?9HfW(Y)=Td8]
CeXA\)QeQ(?E2GE<T-5&XD,-H)S&]OOHbGM(Q<4F;=gTb>6G6O\]P15H/&3K6[.T
N6X[T9/.3c[_]XPd)cR8gJ+cTbC7SC\K+HZ\=C/;F:2V8OZNPAL<^1>TU?YTG3LJQ$
`endprotected


`endif // GUARD_SVT_AXI_SLAVE_CMD_ASSISTANT_OVM_SV
