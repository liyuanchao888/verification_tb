
`ifndef GUARD_SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_SV
`define GUARD_SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_SV
`ifndef __SVDOC__
typedef class svt_axi_snoop_transaction;
typedef class svt_axi_snoop_transaction_exception;

//----------------------------------------------------------------------------
/** Local constants. */
// ---------------------------------------------------------------------------

`ifndef SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_MAX_NUM_EXCEPTIONS
/**
 * This value is used by the svt_axi_snoop_transaction_exception_list constructor
 * to define the initial value for svt_exception_list::max_num_exceptions.
 * This field is used by the exception list to define the maximum number of
 * exceptions which can be generated for a single transaction. The user
 * testbench can override this constant value to define a different maximum
 * value for use by all svt_axi_snoop_transaction_exception_list instances or
 * can change the value of the svt_exception_list::max_num_exceptions field
 * directly to define a different maximum value for use by that
 * svt_axi_snoop_transaction_exception_list instance.
 */
`define SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_MAX_NUM_EXCEPTIONS   1
`endif

// =============================================================================
/** @cond PRIVATE */
/**
 * This class represents the exception list for a transaction.
 */
class svt_axi_snoop_transaction_exception_list extends svt_exception_list;

  // ****************************************************************************
  // Local Data
  // ****************************************************************************

  // ****************************************************************************
  // Public Data
  // ****************************************************************************

  /**
   * Array of exceptions, setup in pre_randomize to match the base class 'exceptions'.
   *
   * THIS FIELD CANNOT BE TRUSTED OUTSIDE OF RANDOMIZATION
   */
  rand svt_axi_snoop_transaction_exception typed_exceptions[];

  // ****************************************************************************
  // Constraints
  // ****************************************************************************

`ifndef SVT_HDL_CONTROL

`ifdef __SVDOC__
`define SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_ENABLE_TEST_CONSTRAINTS
`endif

`ifdef SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_ENABLE_TEST_CONSTRAINTS
  /**
   * External constraint definitions which can be used for test level constraint addition.
   * By default, VMM recommended "test_constraintsX" constraints are not enabled
   * in svt_axi_snoop_transaction_exception_list. A test can enable them by defining the following
   * before this file is compiled at compile time:
   *     SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_ENABLE_TEST_CONSTRAINTS
   */
  constraint test_constraints1;
  constraint test_constraints2;
  constraint test_constraints3;
`endif
`endif

  // ****************************************************************************
  // Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new exception list instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the instance
   */
  extern function new(string name = "svt_axi_snoop_transaction_exception_list_inst", svt_axi_snoop_transaction_exception randomized_exception = null);
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new exception list instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the instance
   */
  extern function new(string name = "svt_axi_snoop_transaction_exception_list_inst", svt_axi_snoop_transaction_exception randomized_exception = null);
`else
`ifndef __SVDOC__
  `svt_vmm_data_new(svt_axi_snoop_transaction_exception_list)
`endif
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new exception list instance, passing the appropriate
   *             argument values to the <b>svt_exception_list</b> parent class.
   *
   * @param log                   Sets the log file that is used for status output.
   *
   * @param randomized_exception  Sets the randomized exception used to generate
   *                              exceptions during randomization.
   */
  extern function new( vmm_log log = null, svt_axi_snoop_transaction_exception randomized_exception = null );
`endif

  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************
`ifndef __SVDOC__
  `svt_data_member_begin(svt_axi_snoop_transaction_exception_list)
  `svt_data_member_end(svt_axi_snoop_transaction_exception_list)
`endif

  //----------------------------------------------------------------------------
  /**
   * Populate the exceptions array to allow for the randomization.
   */
  extern function void pre_randomize();

  //----------------------------------------------------------------------------
  /**
   * Cleanup #exceptions by getting rid of no-op exceptions and sizing to match num_exceptions.
   */
  extern function void post_randomize();

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Compares the object with to. Differences are placed in diff.  The only
   * supported kind values are -1 and svt_data::COMPLETE.  Both values result
   * in a COMPLETE compare.
   */
  extern virtual function bit do_compare( `SVT_DATA_BASE_TYPE to, output string diff, input int kind = -1 );
`endif

  // ---------------------------------------------------------------------------
  /**
   * Performs basic validation of the object contents.  The only supported kind 
   * values are -1 and `SVT_DATA_TYPE::COMPLETE.  Both values result in a COMPLETE 
   * compare.
   */
  extern virtual function bit do_is_valid( bit silent = 1, int kind = -1 );

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Returns the size (in bytes) required by the byte_pack operation.  Only
   * supports a COMPLETE pack so kind must be svt_data::COMPLETE.
   */
  extern virtual function int unsigned byte_size( int kind = -1 );

  //----------------------------------------------------------------------------
  /**
   * Packs the object into the bytes buffer, beginning at offset.  Only supports
   * aCOMPLETE pack so kind must be svt_data::COMPLETE.
   */
  extern virtual function int unsigned do_byte_pack( ref logic [7:0] bytes[],
                                                     input int unsigned offset = 0,
                                                     input int kind = -1 );

  //----------------------------------------------------------------------------
  /**
   * Unpacks the object from the bytes buffer, beginning at offset.  Only supports
   * a COMPLETE unpack so kind must be svt_data::COMPLETE.
   */
  extern virtual function int unsigned do_byte_unpack( const ref logic [7:0] bytes[],
                                                       input int unsigned offset = 0,
                                                       input int len = -1,
                                                       input int kind = -1 );
`endif

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>write</i> access to public data members of this class.
   */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);

  //----------------------------------------------------------------------------
  /**
   * Gets the exception indicated by ix as a strongly typed object.
   */
  extern function svt_axi_snoop_transaction_exception get_exception( int ix );

  //----------------------------------------------------------------------------
  /**
   * Gets the randomized exception as a strongly typed object.
   */
  extern function svt_axi_snoop_transaction_exception get_randomized_exception();

  //----------------------------------------------------------------------------
  /**
   * Pushes the configuration and transaction into the randomized exception object.
   */
  extern virtual function void setup_randomized_exception( svt_axi_port_configuration cfg, svt_axi_snoop_transaction xact );

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object.
   */
  extern virtual function string get_mcd_class_name();

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Allocates a new object of type svt_axi_snoop_transaction_exception_list.
   */
  extern virtual function `SVT_DATA_BASE_TYPE do_allocate();
`endif

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: Provides <i>read</i> access to the public data members or other
   *              "derived properties" of this class.
   */
  extern virtual function bit get_prop_val( string prop_name, ref bit [1023:0] prop_val, 
                                            input int array_ix, ref `SVT_DATA_TYPE data_obj );

  // ---------------------------------------------------------------------------
  /**
   * Add a new exception with the specified content to the exception list.
   * 
   * @param xact The svt_axi_snoop_transaction that this exception is associated with.
   * @param found_error_kind This is the detected error_kind of the exception.
   */
  extern virtual function void add_new_exception(
    svt_axi_snoop_transaction xact, svt_axi_snoop_transaction_exception::error_kind_enum found_error_kind
    );

  // ---------------------------------------------------------------------------
  /**
   * Searches the exception list of the transaction (if it has one), and returns
   * a 1 if there are any exceptions of the specified type, or 0, if none were
   * found.
   * 
   * @param error_kind           The kind of exception to look for.
   * 
   * @return                     Returns 1 if the transaction's exception list  
   *                             has at least one exception of the specified type 
   *                             Returns 0 if it  does not, or if the exception list is null.
   */
  extern virtual function bit has_exception( svt_axi_snoop_transaction_exception::error_kind_enum error_kind);

  // ---------------------------------------------------------------------------
  /** 
   * Utility function which generates an string describing the currently applicable exceptions.
   *
   * @return String describing the applicable exceptions.
   */ 
  extern virtual function string get_applied_exception_kinds();

  // ---------------------------------------------------------------------------
  /** 
   * The svt_axi_snoop_transaction_exception class contains a reference, xact, to the transaction the exception
   * is for. The exception_list copy leaves xact pointing to the 'original' transaction, not the copied
   * into transaction.  This function adjusts the xact reference in any transaction exceptions present. 
   *  
   * @param new_inst The svt_axi_snoop_transaction that this exception is associated with.
   */ 
  extern virtual function void adjust_xact_reference(svt_axi_snoop_transaction new_inst);
 
  // ---------------------------------------------------------------------------
  /**
   * Searches the exception list of the transaction (if it has one), and removes
   * any exceptions of the specified type.
   * 
   * @param error_kind      The kind of exception to remove.
   * 
   * @return                Provides a handle to the updated exception list. 
   *                        This will be null if all of the exceptions have been
   *                        removed or if the exception list was null when the
   *                        function was called.
   */
  extern virtual function svt_axi_snoop_transaction_exception_list remove_exceptions(
    svt_axi_snoop_transaction_exception::error_kind_enum error_kind );

  // ---------------------------------------------------------------------------
endclass
/** @endcond */


// =============================================================================


`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
CxOLYS/sChR0zgPFYfLiRKVuMwKyV4M9DoQlepR0roEG1hR8K8ZJ0x+Uy4c5RyLR
Mh5wEHdFAaij2vRPo+k1zXVf6j0b9MIoM5CDW4T/2SLqEjriaFqpMlJUM+R6Pfki
0+vyB98b5l9ARwue88WTmAl4M2pMXGYJUCO8as3Lo5w=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 1400      )
tvkbs5T6kVC//lWj8S1P7/0k8jni/rVfxYQFisPwS0MQuy184el1iAVfmrisqpzD
yJEKr0B797mgKhNPkV/nk+jEdp8fXWBi0SSuki4htM4A/I/Er8F5cK6OvfLVxnKU
v2QwS7MRRjCNMMEPVBdv8+HqEoV/UiknfqbvN3ONFlpaNAWHJZ2AOHaXHnMbeW3A
2o8TjAMXSDt3kb6fx8a2y4tkydQYp1uKXikbAFH7cd6AY0mnBHaASBVAIXVVdH2O
nxOmFn9+/LQJAJYCfH3JO+5k1QwQLJo8WuwjvuoLEQGJauMJloab93t9dfTmntBj
W2Id1q1gRbWQPHqGX1ZhFbdqENF/RglOVHMpv29+zUfxqd4A8dt+bTorlSVakn+f
TgmZjqz/E3RmCDhaiaw4RKlCh5F2ho2JgEcP9eYaQGyFCfyqMEoWxSMuHjw0ItVh
VYmmBEUTi4z1RiqhzHYJ9s5u26eTsFyqyWwklBok6Ymdp1iTGQnkBKSCIfVYTfco
ebtu2w+CKOjxRLzyeN8G9fhwx0BgCUkues/97YwOrVRVEEdVA5QE+3YCe//pJLUZ
MIDvsjtV/M3iVCfTb0Hy2vLmaXzh8u+4bdoAb72HwmrUBcKWSdN9wZ5HugsuaTRU
lzg/4jFzuI9dMZ+JmGD62a3mMfKCkTBLMvWG4afyhgh7PLEjVOmUgJbxxIDjfY9m
G13ah6FUevbtvRUQAAkqv4fPmceWKE5OSivWj9EX0DVcyOEpxv7kKz8bj/s92DEj
nOs22J7WX2mHYs1Y0ejeV8COAxt0KAGCk04XYhmqWtnBLVstQc9+5daLgXW39704
PDFmi83f5ZyqkbHDXpAnMjG0Zb6ul31bgrBKfKjCj1WSDsyb9L30odaw/jSzGiWT
D2kDXKX8ygW0vNDB/RSB31U+Fm02M8rVevJaqh7EG/hNDzEYAYRtmUMIO6QrNrMF
rgd35BmA8w5JzpI4XqGqp+tN8eBiSZ2ksjjolTmw+8+EYzF0GNnfskHaJ/laCgIN
n0Qfl1mlKyC+MtfcZP1+Z+SeijHdCRhkpZwSUL93PKSXfnoSI2lyBQANFPwSfUXa
z+3hYUplaZccmSVaeq2C+bclhIlM9rkzhllS6zcGqM1vKU1Ubrs0agLSdoW2yTLs
tckUYa3crouXX2he9mi0FKfvFjXFrhBPEKPzwBv8ohSl0a9ulV5yt965ibEWeEq9
RKmzAyU7RRjMp1b28kD9M8YdnVmqf8QCL8Fd6lgUn9hUhrYQE2qntGcOcUCf89Pp
YEAEWTIFFXXCvzVOmuv96t5JTNtkHCN36zsXr/k1jgBHMtIGUCq4V1nSoOjD1LL+
LW32OCvfKkevW0Q25d2vO5wI6LFEOIzXAEMvpVBy/i8rrWe7LkKf0p2mViaRNJzd
lIVybz8QfoGlR9UveUaDuvFDSRaaC7IGaSFSRfXTdA7MuDMSb8LLdxus3Ecp5lnF
Y5A6nEhY85cQQl31HBM/EvRDX7nwik/rZAPl2Lk1tRcdlbY7+5eQHAqaN0h51Ulk
k/YXdECIcQtZL/lDqiZH9J4wc0vimdNUf2PIn5Ny1BF66zGK0Ffr3oJyyTfWPOXl
HAWLN/jdadYeQSMnhBN5eaGLoJMimOcS9Q5pLtDGT0CpHFzuHPizzYCPT+9Byvvr
Fu6z+a1E+cuqzstfRH7gOm+9/ow5yNmj9X9fLZne8ornOaSGd1Ev35shSunb5vJ6
UvYZnRqoabKw4iDXu7s5g7TPwZ+5OOdPEuar9//gEZ8DbDzu4ZAE9HBsFFWCKEj4
iNyGD4xidGXqXBq2vGmztV9SQTo8wecw3uodcPzYE2rDnDBCbgPqxDLoGXdwTvps
IZFXldpJCJzLgf9re7xvRg==
`pragma protect end_protected

//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
bejpIrVrIG1LB0QMYwlCZNCwGbEiLQq4h/SuHRrI0s2ByLj8OCdABo0cH72/nwKT
yR8uIo0kjT0PTAjymYPcKgt0S9VVX3rZSDxeSFelCs0yoDY6A/QdL9F91B54p/Rb
VQ5e+E5sJkBMoeuProdriYpKnOZYidX+NlP1gpm6SN0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 20057     )
41/jJw4RO5lQZFXfs+WKS3nNxqkHHZEk6rHZnaJF3cBwgXLEexk7SzaBwgvwnn2R
qt8jyRMFH06YJIKqKTQtwSTkYKuNPkp+Jy/2Pf5ssjnM286S9QGHkDJK0LSOhCuY
lQhYIKC7DwDO0tI1TU2n9Sqt0xVPEo5Nmc4nj86EWjZAaUSdd8f7tLojBf7UMUQr
jWBOweSI1aRXwsobvJbkL0BP8u8X1UTsGHk5bTQtNL+vkKA1OS3dVMd3RtgUzViP
/cdPy5X2xn+aUyhhXrXfk6+9oejuTyKt/6jJe4zWbQevuwThP/Hodr+5E2A8HFkm
tH4HL/xlBuYT4ZxzI52gKxUa+LqRxRqku359RbFiEdg/ioGw4eJ0SFJWfERaJKLm
mkmcdjiwlEKcL8Z1Ym+gEg+bY7dTd8D3VW3X0lB+/YN6kQCLh+/i0xrRwkCAhyu4
9tTUBjubgru9QwzlmqqJY62olDGRWYh+xq4FuUEZFVfHitbeYaPL0KtQ45e2zLFb
UIcAMvN27ckbPWEflZIte1HcIC2vVeY8QZ0ovIE1OqJ361jyhB3YHFuu9yFFeonq
Jj3M3eQSnvNyILb6euMvN7XqtTMjgyekscOBffrCbrwjk5jxtNleftEaeBDj/LXb
srVIzu5rG354Yx+xkNqQJNrmbTPpAuJZbI/XTbAenM+WSZYUwU8oSNCTaahRtNwU
iTuw5YvcWf6e2YAjsFP3tDsliS+2daLyyixMcM4/1Dn2SMbd4u8jyTW0jIElg44q
DLEb/VayqGh9qskI9X8khKGc7FpMD9teI6zgJUKyuZaO+amcc+3N6cZdM8vcFWHt
IQLtG+sv8Xl01X3Fm7M37V6Jira5DQ/US8qg2C+aT5J2j4fggStKaxxtRGYvDSRs
GTWa0UtDUiLTO5k5HuKElo5DsrKeguV8r68uv5bBeLsitNCrDDvWdXvslXvA0/4V
bbBkBgq9M8HhzGLGQoaFH13PHNc85QsCSWluATLAypcDnmYXA9Xfy6vH04ScpUg0
e6epz752saOT8MT/ULCU1yJkvPoFwCNfPJIn4T9mZCHqadHoK1h4tahdhXNfSK2G
bHgAqELlQEAJT9nImr11jr8zeXNdbZvTUaWrGJNcswblA8vSQX5d4Rg6RP7ngc1Z
svp8+70dNGNn0KGSs0p9UAOf7wHBAbnClaW6UtkVTwSrZyiDQtk/r/bIs/ebbqEx
mNSgm7dWW3qhawYlNupRuwsCFcjuFXHuluC2RQm+wwQxjvWdyEDWqgt26JPUCDRC
v72jvqjCCIt4eKzh3n4u8GE/Dj1NcWOmH1VAhW54Gk4jCdVgcyEEX1lKea0Yg6Pf
t93XXS9TVLP2fYVKHxS3mzCEx+PgzZploZ6KzXXu8IS9EP8ILqaXBUGVTseDGclo
dS73lalCV4ILYAd2JtEy1mFJh2mX8g2eKY4gROom8Y09aOU2vkGVkDFNGcujYUPi
/+DHTRwHPXl7DhtNGAVITKB9/OqqnAqVwzB0KH2+VYnKEIIySaG+7Ni5Cf0TzkIn
j3P6imLVNSXTXot+T3Hg5+k1heGegDbsOCy7ulrqfXUg/pbek/ES0Ik7ikyr9Z1O
UKNMbN+jiLD7WXVBD+G/1KPBmbDQdrTaDLsC2wkV30VRMtSz5EgfBZ6VROleB9v4
Ba9/4598NpR4B02w5DODzkvHmbYsarCQnLKnsnvwmW7dprfdX5dd9JDcZCMAglWO
2o+bBT2DRIWjTkV1ZBS0pHk+lOk24zo8kN9PN5DTu9Mq9bATAgOWDeoDCgs9kNwM
Ke8qngvdFg8LiArXDnh1ZbcGaLOh//fIlfaFoNLrYVKym7zxT0PJT3W460/Dia8z
gdL3rc/kdG1eCkHgZcLMvv+Ta+n9GdiZbeBIpcfLm1qK7bycx3pZ/DAnxfTkblp2
2cs347TSWTQS9ZKSC9FeHZcTd/UZmbmy/cQxEpOmUTqqWTteTzluJuymdUb0sCoq
EEdN0wvfw4XoSqW8ps9slIwRBeGFnbkIlIX45tQB+UUu8lbxfNHuiC01l/Od1Tqb
ZC7FOiBWJcfe7MvmwFkW8CuAruRXZgr1+T5n6jLTfal/hkJwhIkSTeXlilBvsdjm
Fo4UYKxmNJNguVFeOhXhoQcM/sfi7SlrlzVsNEuwvaWA/W5WiLX/pLmHrSltvRe7
5oLJuUE4Uz/50NFn9w1ah03n3EFA9Wy9sxke9TWimat6+LAk0V7B1N1bkbSDKmCD
Vm3Kr3naNpFIbXnSl2sM2tOacREbKoOY76ctMvSDDHfQcRsH4aCifX3axQw11R5G
Yw8k+tteeBRoTb9hyfM44nA6doDne1DqGGbKWErko+eRs/W7NToPnWGNs+8YS5Ek
hVtFM3lvbezR3VppKJz5RUOdKkemxijBPFKV5dwtpB3cqwLnIAK1YGWX9rKbzous
0UxE2Ov72ui8TYJp+AiOagrtB2YLFCFtaFPgtWkmSlQxSHswpBMdvAbkSyLsKUF5
IqGy/Nvv01Od+rneylaj7L8lAHTTpVG+pOXDcZUpr7ZPcHzPuY4WTBUKZ97Rnr0y
tJNjuP5xsvfQAjEbP82qEZb539HmrlsmBVVSAedp/uYiDyeMuZe5+npjDpbBb40N
XJrStA+YUZsZOjxaJIUzewsv+kojSGmRfDV7OkR/KmA8iTTXNI8dh+KnM//VIxnt
CTUcqm0VKJ+8t3TIskdUJxJ+q6CfCy4fGwA9/BI2V0SqpXsKaf7we3pK2hLAYWLa
bGflBab/IvJchFq8yazUn//cm3d5orgcCa3OJGTX4fHhuDYx/ocpZ8ujfO/bYemw
BUzvyR9ihAoZbweN4SogHcWOdXOdClPfcItaBIDdAVkgWQ6HVgJTEYSs7+bjV08t
xuMDweLsq2k9SQw0Iek8zAInM1Lh8Iid4Es5GeaapWuOpFjnzZfZiU7XO1MGL/pz
8JozUVBpCdLECUdvUGZWzOxl4YaPFXmsIOrkOYyNyLXYuKwwfsjn7+ECNcCdhrLf
oLPs2TB/5kZbE3clsBmZotMQ1krzEQUiLDWYCPN/sQ7RxZYL+DBXT9qd5Bs4oUCk
ptzb9gRJbWKyJaWCtMGvImL+DHGzhxd2XSd6Z5v4T8zNxaVsbL6y0XN9IrWV+cJW
PmEYG1KihcIg9yWjFG01GrFEr/wEKgm07A1yOsoo1wO5VHUdE6qmVcv6NY6LHGNV
bka3+hHvNGjaSFK8VqzIqq6fsdTn3B53BXznIEIP4kwtZ27YSOrXgNjl1Fn8YCUH
q8MfVQhKm9dnycyZqKhbH7WM3f30esf7XaX5D1Rs5OCz9j9b/kFyKNDHadf9Tn+Y
97PyAOw/q4NKirukEKr2yVHWvgRPphsF//dv0pebCHCosxR36gj33mf+XlRMCBMl
/0aS13eq5VthSVdlIGc4ixgU4QMKQ6h6HKDHCndYiIFqL2diaAQBO6uLE1woECbC
j56HnxtXDJyviLWc15XPdqibpPZfSsYrHHVONqFJg1z8VXFIqE8KxuwGBvPOx0Xo
bwWV6atZm0kvoZttptFU0YJQ6FabjnTcw2d6rGzfW3ieHFasLgyYwWdA9rhspF4P
n8mb0irTPmaBHHUVhjIEF3oRDgSjpMJDD7QYDe4VgV8cuZCFqZ16cnTrb0hBU47h
HYmBlChiEkMmsM27hQcyqQDnrt3HddPwjhczhLIvzB7ECEtHlPzBB92bVCZ/DYc8
kcTC8hO/ExSWB4CUDesoj7VDwDd9xCWLDNd62hIDnUPbwQ4N/XK5plaijmLMBB6C
VeU3f7PQuWKNMhl0mQmxm6C1c1l8zOIhIwHndz027FMFAGQXKV9DB6SXiykHxc+Y
//GBfdnRUPwAbAUPNtB0Ahh2nETOUDkflUX1fw2PM4b/Dqj3h1/yGsxeXo99tkQP
1VBGcDu7EjHu9U4sBFKPH8sFfiSJaQ9Ho41U/uYKbXjNUJVsFokPp7lTjzOeiaKy
uQrJATBtm3OXk2J/zbX/gnA6UYea0Jm1MVxI4cgzGoY60eeB5AkpR9sopi8UfieZ
5hTr7EPek1ujSpEFIexplRgcYlGiniSym5P01uc0ofvchNQhX8cscIwkw18Wx0Fs
u+jVXMJq9nKKdy3dmxFJMLbVL3tQ8puqJA3BQYmoAiwJaU/L6A15cBXU5xu2w8G+
CqfY9sbRbmiArfxiUiO6TgHYbJPTDbxJkAZ26KJFeur53OXfnfP0CsBAuwXQKPST
OVtD7Gii+pfgvH50vFy/YUDtbQAxyCHUDxnTZ/7QglFP9oOevFQCbfoInhblULRl
Pgp4hnKvgjF+cMyw9EGBH5BjWopIvNamfiGe0qLk85sjC3YD1vPssa+psdMYWUBm
w5cq2baSksozfNk/c7dXQfUwzMgbbDTqBdDEOrivie5UnUkiFZ+TZ33FwvY8Ald9
3ebdAoGeJnp6cbwaOuGPbil+c4mH3sE0gOpwISMfbEpplScRuRj2cWGj7LRdA1Ba
a67FI0/rgKgKivH6glecBfMWpVauXiQyKa43AMKb3373e5nwMYFroJNW1XIms3Fz
btJ1LZ2tilgaDabUt8vxq5NPElL1SjRvfoG/mOdBLjCx46adwEjS5xNuhJR1IBYu
1onFhwRUIpJsZoprHjWmIkbd1BuWzYIpShXfMt+roAC1FmB9c+sLEYpCMFdsBfOi
DLTZYpod1JctCtSKkrwJPQnnUdxP3dwszCIGyEr6Wkb4Va49wHdwBLOW3kSbuF9m
tnf0uN9u+uLJL8utQQTHMhcYriTTtmMBFM2VHw6zX9wGJML2m19kagbZ/HMR9tYD
7sNm5ZM42wC/GDZStc5Nnw8Vw1vXtbB4w4NETpfQEWUIfMs45WI8c4zJftmIrsBR
LlOFyZCTUoP27emUjUkk0Gm3GypQqd/r0lalC7lz/KiFXfwwiJANXJzdMPHNPU6n
PCZiAojYS3yzt2pxxTwJm72ldHz0pj6iOBUrZvZ7BuIwvHMPk+7G/jvIpMltAOtL
f1NyBdDWhX1TEEMTtpCBMr5wc0orLaFuILqEzYhzSsxWqLtVJWs9Mh2mcF0mk31g
HXAhykyFV9cU9Y5eEqtxjI50KvkwhtH2XEa4ietuhZe5K1bZIsjC3flQFJv7MsmM
T0wGi9UYcxsZu9gqMe4TgQPY0GT//7US23gSEaEvOjIIqkwJ+SLyv7WNMyEgvZa2
4h66GbHh4oskD/J0MqzF+aYJlbhOcAfGQ3d3VPnBW5e+bCQpSWBrqcFmmkDS77MU
pbbBankNOXPG2gaKw8WFlGHObi9lHADGitmJvJpp0ODgZQmXCZzkUKNKhBZSR9jV
SCybYZXj4u2Tm8anYYEVO5P7UhCp2XhW4wEpanOFBfmH55TExPaZ260c4BXHTLoZ
NL1m4E9GUX9h7AuVuUZuemgSc4VqzfKR5GySOH29wS94Oy6SvZ/Z9sdKReyY+8NV
JlXpmOwAWzgm9UpbP+9/F33ZCbKagcYwPPZRiJ5YT4rr/jaERUACcKdz/ROi4iro
FwlYl4GUCb6s7juOJ+g1vU3ao26vz5G6U+bNticlL+ARdSqKWVGaqHDt7oymsR70
hNWobEmI1NhutzXd06Frxa1+6glwsCpv2iOHVe1WJwENLx4p4Kd+XaFXlAeQECVI
DcIktW5/PeUr2nTE+NbkUUqjXCLJMyizMkm1qXltHUxD00TSmxbLRpDQZy930C/x
kt6exlpZG7UXjLwUXz5UAACC9SfngIoT2i4SkUU6zZzEkmtcYLj+Rcn4Gwwy7RWp
hbFvKVL16t1fBJ45QRcq45AbwUXxkqe7UABc6hW2LIfN7sXa41tl4ZSgtt6wm1Bc
UcfLI5jl4XL/G8JshWS4Pxgd+8Rf9jCPfCQSnPABUHsMU/mfQSiVPzb3fXSAwBxH
gJ0YdKxGOqnMTbxslS0G06xFq5uSlU7khW84N7D4j7QLs2gccZ1iAloxn01xol30
g+/VOt1cebKQyd/zudKN8WODqMcSXmS1TvjJw6g8OBFQ+FB4t4ZX0bSijhPAb7qq
kUDFVRfz1Uq+W8DVpl6GyT0VGNmj3cR2+/IRj8+2lUW1DIeaVOt8dEFPqh0DOh2N
sPpnVsE1Jw1ADcZeaC02X57QJOWiEaHcA4LT5spwAzOeSOm3CvYp50Mid0x0BFUc
nBbWG6cG368poVlMAavJyZe2XC9Xu5XPuAPTrl8EpqtEj1SailZ7B9ui2vJcE6FR
p8HqfXtXXk9I8+y+4v5VMUsGZxs0sAKrofCCy2FXy4a6TSDuwFU7KNzPN41DVxaP
Fiw8dJR5Fc9h0DlCZXDznDDD7t9Ze+OQloVVCLPPdTjk1ViTyw+ZIvJn+w84VVYP
ZuMRoC/7q+n/GVz/idoy/ydAqcGQxi+zQC77MVO8NQ7CGdyYbEX8CZWhfhbL7D+3
WhQLQ/71BjbtApqm3df3NIj+GsrrfwBuPi3wfWxXtHBaTRP5I9RC7we0cNC5ktrn
21KkEvRxuDdjFWMRDiTGkjed9ds69JXQgrLFSDity5Fp5mtiONeqwWScj4XUf6xh
sha2ulVmsfVVgwCddscBL3UM70w+IZLl4y6QqsZAPsZjdOiJwyJlJm8c9pZHdocQ
hZMCmiQ7oZyv+YiwYReK7k7dT1BY68a4ANNGhJW4//XY+DH35CAcEsPzy4CAzuhY
JhQQVl1cjd4A6+T+HZxNU9UQIAEzzs+r963VKsXJ34kNaEUXLRmZZM1n2VVz2IJa
zmdH/WTZVGQa/ZGkhnjS1zNdG07THK6qUmxvuIQSc2BkCN7OS0VtGJ90lC1dtjbM
C3ac1SWGkS6oB9513HVocMtyQMIeAhFzuAf08DMr8lEIX6mBmyoJ9CeJG25NMMfN
2iT1bU+6eBBHkZvgyquwsVLnKroSlId8L1rzYdKMcnTYcBqjp+qmj0y0bqhle3G6
P0wXfhYG7LmxLkKtAmaTEz5htOUFdkEZwAc/har2jyVusdqA6zEKnJs+I8ynIKsD
tDTIipCaM/ST7uMYuMnQTDa4el0HasHWuBh99B44oEARk939B/Nczgbo4w0LwFwC
uKj17KN4RgJWOdSWkmbttqSAtb54EnC62lX2nu0xbuAzd2qljAIoGOSge6vsvNh4
8e5iXLrl5MeRV2jicGxYxmnQYRp7Cs3WvUyCOqjQxyENNDuXBzsl9yDN+Ohgy+ua
TfTWxo9ZkiIWlap0WYuUPZlfUQbHLPS9ev4ta8gp6rvgJcIGCDRQ3wopLb8Luax8
uRS/x4t5GZyyCmEoZ1CFHeAm6fIkMXC4vHw3Aj4Sznyx4f738Z3ag6VUVuFfS7qi
ldiyjSinqZot+sdJIvj6IRDRfs0GF3QC6lw8QgbrS2qF7617DXQWevwrYyMADAph
3JRIe43tQF18SZxcCLGTtTvZ5dPVAsZ2143S+De9w5zTKnNjKgemXgPbY3Ss79eh
uVy9L4xSMFL5REdEI0rNhwNcPdj9NCe1SjycZrczR3olnDtJbK9N9YyXu/66S7i0
fkm1u3sk/HIJM6s8V+cmNpee7gprE0wztFULy1T57kSeoQ1ie6UUjH9Ro7aPv6ur
MFN5x158+2oBQccFCWC2F9y3cgNOMzaYbWKwU4rmqa8B3vAy2V1T9NK0zj7KQK9G
7iEeqGv5M9hVKCgUkxUQhKZUHJcH/4VEEhoR1eUb/xfBX9evbFWtMGc9XniOdaAQ
LHmRVZCw0xtBgZwknnNB2+symXiHFqFWZWXbIgBf7N+tLxuxFFOQ7ASo180PXEUq
JiPCt4y6HSDLzDZmEr9T5pqlgIRy8ixiSf6wN5s3c+JIGRzJ33T1tDjwFD8uYm6E
1mwJyIUOyHwSEOk3gBNYxHgdAPjXPkRB9tihnNUJCNvwuq+votZaXjvUA2Gp6ApW
7IcyXQ1QfiuZFIbb8zgS+lwdE6l57zy/Zm0Tb0BaYPDg3SUl41Tp/h/Mno9rEXZ6
7hJdNNZUXeg31RmScd7msRw06BWgE4jdhfaKkBcgKucNKAecjQQI73akOq3zKrwI
+r3TkD+1lqMKWnhEOnMW1+tSUxHns8aOCi68Ytf6Ve3WBYvuzsctjjnjeom9RquB
cVLxYycI8fNgymwu1UGIv89uFOcQrpu4tiy0M8LI+0wuEC0erBe+2uHQSlf7YO0+
pUPq6Qr2mVQD+BYyjEyeqF78DW+T7P2I76PQZ95tKVvR193VARF70TXD8wY3Qb/O
mAOvDTWqEZhm7myO5wX9eHDEVOuN5HxXO5aR7uk3mIaN6Q1b0xsiXW0D6x49PEub
JZug5OPark1NvxZ5HCN5+tpiZiHbT15XJ7j+S5EaWAH0XDmIv0bx3VxtwFZ5a04O
yldhfcwxNN0O4nYspMqrHfphXs3YK+siAWl0P0NFahVQH7em1vprX7iOyR2n2TMQ
O+GHKLzDA2KTvTM2niFhXRjTL539vczf6DBmnAWHF1R2Ey8ZrehIK3pLkTfNUtPS
gM1X+229rp5LcbgL7QQHDuwbsu1hZMgqU8hQwnGPFLdnWnaUPXkx7iqWHwEb+Kqw
CypxnrMiuOVwkjWYfG4ORKU9AxYTl7L6X/Bueo7ugAvTbdIVu3PzEpbv5QMYsEHY
T11/klidW/D0GzkCya+kVxvVR15c8HhAoMh9QGV1nsWJS+eT5BYpslX52Whh3NUp
XU9TLkpuwwRzoiClIYxNNH8nHXFUFftMDHipc7bkWVWaTqjpCFL0xx25lz3By1V9
er1RN8vievUK9jq8WBArOUQKeOEC6Xktq/ttyX6wQyQFflp9wvXmduMofLsBNPPs
j7VjDmCkQMADMjgHgGRUMgFEfsYsYpzBeZl4CeC3RJ3UOVGgv126XWTOVY7mMJtp
C3f4wOYE93QTeLoobXDf6N+qXnVVHAR1dOAqy8ortYKtuPdK+uS+ZLDpURw2RBBF
uEp9Glh/kXEDjo8NlO3dqnwFoaSwvVliku5fAbfaWveDPFJF4JgaU6fOwTjcSFHD
RlO2QcunI+0dJ+p1JTNcBPbLHk3z6Mhi07Of+gLiIei0Yq0mYx23bpzt8NsRpPgW
sXQaX9lE1BIH4NdwSc5TB4yOYQFHSXOZcLkXnLbG9MwNtCBR54XRUBf6qwZ8GUj+
OhQLjEu3P+i250X5lyDWzqJR4lfTrJM5KiMyyp3R2Ajgt6rchsWQi5bgTG7UktTu
5Lot8n2NJZt+mWAMT41yLumdH+rvD2+6BlNOTwtbAityOnz24VpFpgZygZiYH9og
PcWBJoe+9AkqCIAygfnnb1+GMblSDd3c+63HHm1FUE5B9SGUot/4aAWwKTy70Xvp
DuUBPuMw+WBgaVGhm/ngpWbh5Nq7nx0oVWQQ2u4x7Y4AldzJkWHErZgs9IpRLJ3e
dxk5XAkH+Ke67cS1i+nCej+mmR26avzEzqzCewv0LJ8Gdi83iQ0JRYs/z0w0y0Ke
NhT7o0EtUz1uaa2A6gibnBB1pqisBuHOOwQbuCAZJqbEfQtMtxxr+fAACA/dwoVn
Qzz5GlWQNuKKPJfwABQaCl02JrNk6R3j8wwcLwatDC0CuGAIVc/hf7qZ2E2peGTC
rH5iUQPXWyVnb4yhjuZEg+V8vMByVWjiGFnkISpui7hBUXvnXkFQ4iogBXSqKK5i
/Er2jtz4eaI37t4cZBAtN7iYM17hfHEzZMDtLRE5lcjYdMOljJH+jS+YiByeATpt
CesAyjY0tx8iezDNcFzvIuUM5F/gRQMi3Rl/u6cy/QIKSxTUEqLrYLPa6RlDkO5F
RNtmsxyu2DI2k7XMSv6ufdQ1ox56gpyBYTAmCIhPUxMnAhSAoTIrkkMbFyV4rq01
JTOdZc37D12l1flKFLGD2Hdm1UlYPkX2V0BUO+TOMY9MRcstpJJ3PwLD1geVVzzy
rSxiVebiTKzZvoFPW87+fDRt60uVbAC0qIJ+f8bIrU7RWoiWJ4tKWxP4g72CeFSh
zmGg724N2PPECKklSciARO+gnTR0QHOhpZ3Bt9MZya26lzmwtV0f2zsCc0uoAcm7
WORWNcqTHSpLAF6tkSaY1hTyjPkA8n3rLdMZyYJcmcKMOThm0IBqTWVOf8aua5rI
YNSU/ZrUibzpyw4FokstZBirLVFcEjZC0e/WqT9vwcHyJni79Tys7KSMWq6Vh9lR
TyeQuAMEeYCa0ZjR2oqiGJXN14fi6Ze+6YWVonjJ/AvpoArwRFP7+YE2aHhOwyHL
sGKS19nTtYVhSbTy3qL/dUClcmPAScYAN/k9RVyuXdCPvukV/98uZlZ/KedyUz2d
epAlNy7et9C2jyMkMWrN6sLHYxL8KAq3CAp6LwGAvq9OQZZB7vKeptiYJyaXcc6D
xllBRVTjd22zk12vHdL5maxGMkuU+h5mEcttGjs++Ujxf1ggtz4LPMPjuuZKTr21
y5EZcWZShd4kkdQowLrj9hPHCRkcSTXWruwxzjl/JnGJMXWEzs6mUwZquQT8kB+0
ODS9JwpdnxU6L+Coo6JbE2V5HI78NrPZ1mVcnpY2cdgsv1E7UAXaa8fkUtpzg1ys
YKpBcBSLzdb7MB/yfQ6iUHd2DoXZHMNp+rvh4BLBpA6T6uLjvcK82YgRt6lk+Jb+
ZEEtUTziwA2U1zCwA8du9+ts9j0pSdZDUSZ1SvCl/Gx3UQYvjcZ9kLrha6ztWbpU
mYXuQUCefpcmkKbDANGCp7L+NFOzj4rh75VJuYZyo55gPw+vo2wvgSiN5BjbXT4c
zgbAe/VqLFViz0UubXaAyQKDu7kne3mgt50Bkw4BOXI4Sih9mEN9JXYy3SSCf+ZR
33AQCZ9099plpr9ueh06uweZuhx7r614c7TSHQakSoSox9hHEY7ApOIIK5JM6Ke/
faPSjxdmvKyOgPVMeY/Ghq0Xt3uaSSkQKHeS2rzuqDn1DPLC50Qb/1RvQc4xndlZ
2TdNXf+atUuIBieWxeqFi7wn0txCGM3SsGvb0J9tFkoUSLjHuUnu7htw7e9Sw1oY
96DZnSd6NgB04N5Qy9aqiNglXhZU6o/eoSiwQeXFYI0iPJRMt0M1Il5StumE17f3
MS6oS0RrtBZ++vejYfyuVQldTndbC18A6wwHuPFIp5PnJTL58WXX6YLa7wgrmhx4
pi7uQxMp4C4QLny4mt489AtMPcAwoNjNR4R27sQXkNoDgFuMsAIOc/qxNpuQW9/E
73fmNoSVDb1tmzah3X0IOAhyEaXlvTlz1vME74mOWbpUVqueKa5JvdXPuqiCy5rV
vqJNoj24IlfJ9SnwuetYWbKyPg3efpJCjapRzmxlQie2XGVyNO8ybqOv52u1cuc/
zJFrnde/tQAprJ7QMV5jpGT3MDs/Te121Qp63/IX0BwL6CcRDLzoC9Af8jZU0Tm1
bbjvlDF2Rf8xpMf06OWdg/2swa1lbY0yhURYkH5H8zdtx/nPwFlqYdUAgMbm+JdO
jvaB9B7/dFykDJdr1EMqqvB2Hfu9QxjWJ9u1iEetew5BEd5xChiUU9lzZgMV4rx2
QrVE1Wh2h5oYe1rVcHyWacv8k08UMlVC0R4090pHiZw2IQUrY/RAID2eXue2GHfS
yWMsO6ucHVsFQF0A1BgjDexFDKhL0/Xxcr4xYaDWU5v2uNZ7BhYV/ltLmjOT75cH
XhlIIsrvrPQXOS2NKGElT0XV6/TkgMeLcVq1WsHIeEvWTW7c8oO8Fl4Pa8z5MGWK
6WYSo7WGB7KvbILh4EwrqHkwW7CbXV8C1LULAjlbHRpZ5QScYjizBomUjk4GaI2x
bT0c2RvbhCOa2q2EyNJcIPoilgliR3l/anoEeGq/gpT15Q1BL4MWAERM2g5ORiqZ
HKwpr+aXBIsXAMpchvqbjHZxX4h22N7s4VlzQ45TDtLFVm7vouGi4iisPUzJmFPM
HimDpKlLZ41TL+Bd8PCSeyBLZcB0lzU5XAaC5YqYSn2mbUBhS6s3LzUwfeGVdah8
cAZxkL+oqiAd77c21yNgk1arIwr+VeHWyjnBzKmgIJhKa5w+L5u5/xLtweXQPbAn
+H8/5qmFNF1QdYd+mNLkzR60F5xROS5ef47DDWmN53nWD5oyprqVyP5ZdsBQHrdx
Dh3qGvOx9Kt315tvtcdwFDnPJAw8alkVxAB1YaTn4bd18ihS9A+0aN4U2Q2ZA2I2
Apf9CZdbVq7p4Gg5s3aTx5iFBHAlGIS3qgzypMBFP1XFuDrgElzE8pf7xCZVs7t9
kIQOCfU/I+9lh2+dPXOBna/eUwI6TrRXJMdocUQHRUThd4q035zh0U31VVGhvOtq
x1A29/RA+BlDpLaxZ4UocxLiJPHv1jjMZXCaLkWINVWNXeSJ7RHpadDmuLFuetNw
6awv8QnlZ1UZGCy3EZqzO+n0Uz470LJuMZD3/ubqzbHu6qZ8WtbmULYhKlyMUhSU
iO1kcqzl1hyfTRFeERMbylHlIV0eLQuij0GUDqXvrH7Q6Z4FifvmNwXGyn+IpUvO
6n7UguGJiKDbWog90+/047zkGbRx+p2v4g3ORLYpy/btwKI20XZtSTiqwXNmMp7y
2IDvwgqLFlt1miy2njSkKe+oGYTSlX0fqzolsoSYty8iejcgYIgD8cJqqwShZhR9
aEzAffNSabEW5b22lCOPFRqDic8eaSaj94gaZUBWmxL2+iTwM/j9CCBqLH/AraCj
kdJ14wRU2im80n+Jms379QOd3Wpqrv2h6B7hDnxY6LGQbwEefDWhRdojiXVMQPbD
8/G2JQTI4672YWBEJ7rrzXZJ3+D3+PwE0rAyQ/KXe0rizF0TZTljgeJgXYNBLNoO
ON962nn7PRMHbJ2EUO6AlsX9lRb7r72AX2c26E3o4UQYxt9VEpa5mJ7K4Z/X1gYr
e6PAJ0NXmNz2Q73KrfxrPAckmZ2wV7ngR3pWrIqqsoUfNrIHvahSuCEqKR0UGUaS
35lFsxPH5cz+6/Obj6rZNObAhlM34f0aOdfE9pc0+AiDc0VWwVBzW0ybgddGWwjm
ijtHfini6tdhN3Z9tPteYcmmPBbIbNFJVgiObTU9eCyQ8qHadI/hVhsoJlSVjTzG
rsDyMrRPrwJ/i5zJ6ilhmLRaFk73LOz57TXB4cwe1iAco/82JujnSkMfk9dL3s/i
9OVjeZvuTbMil35Cwjs62LFwZw3qeCoTr3/HidS0L4vb1qYVaJ/0ZG0CuC2x0Gip
9eYHhjHu8QnoEc2CW3IRAnTPjHn2zz6MDssjsgUHY4Xg9yKrtw0qOgH9G1eSb2PO
6+RkfVBn5rsRxPEaCNPRFt/aO4CtGirsf5YK1j8UQ+8GJeQfXFWixDLqDw0/ETpf
1CanRdqTBFglrph/NOuh3sbwxp1ZoZV9/39E4i43F3Xa9XjgBMnZbqM7BFfbK+Wc
cIPzBbz4eUanBFauV3v5kLEpYRGEDhN2/eMVglOsZVWKrP9Oi1JZGOcJ4iZATKgX
k0RYS20hQnRQYjHCRFdCLtBCHrt+b0od2/KEmk7i3sePpVI5Ra+/cHEunlmRukvy
3Tj9VLzHMlWDbW/qdlDIDDIVtEIV5AFa4krSIlB/0UAm4dnrcGIAKogshHPZox1p
u7J4S+Nn4++mIetvdLQM2HZvpDzPq8hLJQfvh1pgmjCQ3HHgyrh/gMPAuexnSG6N
6hiYaWHtxEYgohGqdoypTCWqfwr06Ao/dSPWKAznAPUFl/gMSrOdrgEcGN3SFpa0
GVdzLL2aJp+oiEC9XPpnCCoYBoQHf70HeqbXYUslrxQcS6+iKTs+qrP0lctgDf3Y
4yTz5zS/phORnTfP3SvQYrb21UdZUpJzCbnBaRMGVR64xj3HbA2ZEcS0+JXmTjgz
+JvlhIkqjQNUEUq7P75T1tjJG7XChWLf6YqcibbcjnKFIwAZKuZJkTGyI6XKoQ07
6353GWai1vkBOFPYAFiwJ4CqZClZ/aRlR7YqfvgtyVP1IslDU+nFm78Ngs/0u7e0
akROL1wxpgW6vLsJwUw/WHSNfS/kvMPvaLnXAU+9myENIvCu8z4/aIfN40u16b5W
9jzs9ylXb6Pct1doPh3xdDUShcmGK+tJJiZD+lQlxEI5BIhO6+oJBX7QWHI1Z0hY
JhijRvtYR82IRSMAL1CS2qF9llQiUJtNG8BNl9wmXi1JDnJ+nLaOCOBs/nScHezS
A6QoHTvkYgI2dMp9MDuaC7c9//Bv0g9QpJ4LBVJ5/VoQThFZ0jsXYozX+YvEbEWU
WSksEiwLON2PUg7NB+XOzmsKNMOp0kvTQXGEiSU2ZhKvgQkVXehBMvWr4QRV3vvc
z7YewswicS2bWEvXnvMCjT/tZ49XzNGve4eynIwgAUFfo3OqhlInXWl9kdsZ++ul
8s7Z5H2Bz6bAPYp4OjuM0Pw4KHO7d8/Xw4Bb0RYYLGRpiQRv0TnGlejEFelxEjyh
1pza1M+Ckg/Fi9EUdgQIth8PI18WrvmaT3jmu1RGRVqAWpd0QKyRkyWeID89pm4s
59295MKO6tagS+DdpdQG5KNZVczkS+V/MaOCsPXIulqsTfKko9hAjsmiiUTDUXgP
aFYV76RNoOvPbYT6LLbIaDgW86x8jlkMMDqjtE5LzfIxCoJi798/Cdm6+VHJGSly
cDSzT42IM4BNIEe+SILGYd58PZpRCBHzuc+aOfkDEM7MemoRk1s9MiVYvaRFDmSS
tjckcL3sCmbfJdo9PW//uBxrwU2jrjJW4qdG3Id8sFTyIHPrvrU2WvTkkRGWK+Xz
pGc5wQsq2Si2uJtpWnwBfEM8zqj/00xfPEvlSlUY3r3cto6XNMSgSL0B6m5lyxdT
8AZAqhK6Rq+aTMbiuw4kDM6ccIN2aajuXYHFnkjqPA+9EysC+1OaZDU7TJHRF1XT
0l8TebSgR1CeN1iIavYNGwlhAdC+SNvLzTaJIaGL1IL/bQuvrQtjmJlOVookq808
BBLX6p6gId/X4Dy2YmkyF/2Tey1bl2+uYCZSYDHFtF/CMeq6kb9XnWmQ2FXE5rZ9
8LcChYdTwu9KyceHV1Mnz6IjyNS836ctZwBJJ6pN+IHco0RGx9o0flYAahhwjSOP
+OWTbe24pgCVWCBlmdiydqFelsA9maJtED/l9Nh+xiPIAj+o7rotDBzwHNRfC6lj
inxOWuUXVZdu21WStTl7PtnjzfEIWumXZkuanzQx+D5ue60DhDlW/bX6Af10S3st
y7X4z5pcrdCEtzXTocSs/MbxmcEigHDD1EqaHNUbiKJDwXcj3MP2varBTZgF7ZxM
+i/kWjq83Ls2YHjSeABj+OzFCuwdHMLqWHsnQ8iGwM9fTz1MMNtsMj7YIzVk7a8y
2sSmJ4QCdHbkl41tBf77M7/ixisurs1sWHoGNoQrxO+W0AtHiXFQJtvPfXJ7q+L7
L5mg0XRrvBGNJPou+dgXH3s8nJgbTLnBq2Xq4dkRAYUgZXXXDhu/xPSNwGCEvDMo
ntKbUm17L5Mc7B7wNwjfS/GCbCzL7/6N9bZ8WECt22VhhUO4CBRCASbb0v9g/NCA
L8nBo9TN1MgKCVdb3EK7l89qSVyGFX7Zc1duB3VXu9pqbfgT7k2tNCMKaK/qWUi+
+3j5byb9KgXgtHV759PZheADrhdQd3AOJsGjjPMdgZ7PwqC+6Gr/44ZkNd23wgDw
UOrESIKiTvyRrd63ANVoJz7S+038hSq4VNdwbG1zT6jZnj9UNYZgpBiSZO+hP4UT
5tE9c28GtsW+RLGw2N7c20H26Z3U2l20v29GMv3E7nI4v1FqWNi9bSp5Jtb5Iny/
sIbVSv6VoUqHfVbjwU+Wlk5LMrjYJL6SkTJQ9KJSabesdKTGfNI5zbHMprrEy+9c
i8vh399RRUvA+7ohYNvYStHtK4qD50D0+HvuSLdVah/tBHEeZtHmUbOr3Ay02BPN
eqDwGBoYppak1M4VoYjctWJCec003Bm0XY/AxNVFCFk9aDJ92D/H3VtGQIgqEbE4
DGcgYtUzwAqsgbfhwX8NpNRNqRNMLpw+qmCT50p9EmCx/VORhIKBXF4IQ7WhZY2F
Mb72eBJnLqguysLxy0HxLGrgw9JEbRe2w6LkujK3zU2E2DkX8nl/agfkjk161lzT
incOC5wrEl4aEmlZgz1cbw43oEcPTzEB0OmtDxGWSOMYPLFhDWlmNIQrDmAjhxx+
v2qfTK1CeurQOGo8iCUoWdeqt4qu5rosu02CZ2XaV3UVrqlgmL5qPILm/eSbxjs6
Bz1cAFvuzHqBF+Dfp/hA6LyIFifwePbZApp/QGW40dxVy6leBYNFEzPvNjkDwHDO
77xSd1TfPTzcLsnC5t/d0fsl3BVnOefCCS/ZJpiGAdgZ6Ao7XcCiV+i4Wh+0ds9i
LSC83xOxKLs4A/KEGmGY7V+m1/28jYaJhJzRJD376ILC1v6EpPfrisucDjJbYP+G
QXTi+QFxZpWtzxBhHD17xlyL+BAxP8GvtDKdPnLtGj+OfN6Mclmo+0ZimYaPIzJs
SSOW7lf4USWNTZuGoZLPje19BJHThuV/sLf4G08HMig7XjC/jC++zmc2tlLRC6eu
gIeW4Z7Xd8/abQ8vojC2cQl7/eB/p/9XyVUtTYYCLuoXYlVsaZD5RE82rSqguvUd
MRUoS/sX0VSc2Tygh6nyZ1Hl13ob+mls6NPg1dhCwNeH7lmyfGc9cHO568ovVDPg
z6mfRclN6+OzcABbmuRSNmykKpYL3kb+oPmexPe9kXLAYamoMKtEZjddk5vY46nA
f/zfv7eqoq3fEJArRHjBXPEAfsK3WZTd1jC344xkw7btJFLrNnhMadtcWo89Gy2U
miO0hgg6/5paCsoUkOCkrPVdOoCIp2V9fPNisd2JXHYS2sKjGiC4HcenjFq2UaP8
cHLMFkIavaC9EsnSD2sLIKjQyHORezm48tHzaLPxKoLKG/kCh6jTZNOcuomgBiiO
mjrLVNG7A6BWBr2t+tIuhieeze752oB0pz3sH1v+OXe2k3Hc7ZslRhbT68bHNi7m
ikK2D1MZwQb1BEtLsMBE63kzzRdESh8vxB4gDhSUxBmIWuZBl8vXb1t5RnL7TJcG
xK0mQdkYW1kiyKubJQWnvQPvQPqVcFADUeHM6nMuRvNrxl5YnGfmvVN5oS2P1vd3
FiKVJfgd+gZl96F8amB3nPATLt4GEpTLcT131VD29DTvtADCDcqEU5uqr6ZKZvNE
LfOrAYmrVdBnEc58IpTU1pIahlRKpW3ZA5smtIEoC+3mr2Bdhbb6PCeGo/R2HFgM
M23gwcnXWbi1BItq+2HjzDa1G4+dxT4Svm5G99JqXHMpbJtSuOBxqCO3QoReZfEc
EIj5gvOCPjitp4aEbEITtLya0/trIbZOqELjS7tfRYonJlCAiXhPujs8gphb/VJu
C1uJW0JI+rmazw7UorE0KN5LzSn26kZEf/tpbOfrxjKk1lhrHQ63A4Lk2CIj5UUt
PT1Z5FPeyRFSw+tHQ8EdCrSjuM7fyQsXDQQ1xVdDcl0lqkgR7qyayPbEbQmRzIMv
OicUx35eJfOGvt++qksUTolwdAkC1pORjvqh9KkwTXXUtook6VjMhSu1eyv0nG3s
uHXB+pRmJODxKzARxeTNd+UAxLCPTiUwI3WiSUMlrFEOSDDro9PLM49rtQLKLSQa
tNKtE1F6WyPcBDSHawSuNQxG5FZx5zNpCe8YqVFFdUsp7GnQvpcTOyfXwM+xexGq
RZGg/VCcq4Ek4UKyayva5euJCygCyy/vZjc8xFyVLQ1fBRGZt6TLCXYVRwyNWTYv
DGQQR7S0KDqRXite5AnvINOxtgXk+EOvkWyJpd11Fqkm8mB4Lb/eukiTmggRwEnl
8ayKTM4T8Sf8/Saj5DkM5pz1nmffATyo/tVqZACPTzEDFEsFt7YNnr74LOp85aAJ
oUZVtXD5/jlK/F/chPlZF52SmWFGiImEdJnQOYbo9QWM6WKuONLD6U7y+APzhr/m
wPhu6jKeHGCWZ4htaQ66BZzpQqdu1EsL6VcgNtmHnFbaphXO2hNqmnZ6U6uEO0pT
VXtpWbT6itjf6PswLQH20KjgcKM0qXMWUGfRE4X2d719vbVwyrVwfBEsPPcZ1zS4
JbX/Ckq+SHIIDspBQ16pBERslSQ0IsuEe5dxp6FzOrFmEZAt/P5plBaMFr5X1Pv6
54/Nj8VNi+njSEfQ0+lu0aUA6b4qqujAQZkfVL9/U5QrqI1sGKTSWjgbpsyQWXh0
FhKXXrA2RGIFkFQAYrdqxS0uHJKM3PL3fJPh14AawifrxwXu/F+YbpON45nChW1Y
Ru+1i2VsMATC6h9YScFinfHc4eHgA+cdhtgHHFZoBTzTfVglMjOZ2qQXnZuH+ZLi
8b1DdiyPfy5yovLbx+abYzgepzqySFIwiI5JVtPxYeJgfqzDVITB+6vFLY4ztoLw
vg4cHGSq58jocx6hFpYrbYR5C6H/j9Xq/KECcuU9ZJLksoGwbw93icPfXLjtJPp3
Oa/V0/qkT+KosV7FcrDfuGq24YTWq5l9d0SciowEyQS5d1SSbkJylbugq23B9Ffu
05ZM6ZoIao73/Dg1Ihdw0HtGgvlivYCEqW3xUztR/Xn68ElN7+Y4DyZWCFG2OWhr
iqtK9u8CXjXCQGvHaag1U3MQJp/CIwD9Y8jKwgEfdHrhZA2YFjlLeoZUbDSh09lI
kf79Qf9lAbsIVlbGe+HN2InfdZgdCD516atJpMFrvg1oJifau7FfXaHWS+5YPdf2
m8GR1fbf7IkiSCRLD9Wzu3vXwnjEwlrQU7NKrwFUL3zifoaAp4ercWiLGaVfJtA1
4NByx7dlLa1McxWw6eyV7iRErH6dgkvELZfTIoq86nS5a7jWtQwgiY7qYVL//nRB
987FnGkUmtsoeiZ/Rn3FqCjtXm7ThPxuybK/3o9ypWFjFggVxfQHlf6vhSYGtqyI
DgewlAPfFTviUXYjq+Axaaj246LB3fltG9YfGjhxaOO3J4J1ojCr/wRpzwT4xuz8
mZ8y10ar3W8yHbxcct+l+ZliTY6oF/Onk2ZBm8v2ivLSRsBsvHjfAvdjSo7Ye0JH
EGrm1EMSNCrWHXIXgjtrifTvC4AJAEl8hojOEwjbNZ+5+Gd30wNAltbYv51UCun4
Jnuryked1ZB3d6fRz7THEUAopQvFzRAXz1grZsgLAI2QojbTFH3tJNQw+hTUMyB/
VhxLQ0bxeW9DTDY5UBWPyBWV7RJj/z6hmsxovnV0voULcbK+p7+r68fe50A0J4p8
iMsbu34ryH5IXvbijNI+dP2egJjBnPl4iKvSRMPz4Fmt1W7/78ERyxiqZ7TpFc1c
y2cLzy+eEtClxCJWWYS6TTMpQDbaIDuFKhJnVt9yuYQjo6+ipoDcp5JYzvtBokJR
OU3BSQ43Cs1XIJmsPBY/vmCGv628n6iDLKK/m0pBBP8Mxoq7vpPKKAnnoR68ZiuV
hN3E//Q8Btqcuzb8XTCYCdpGWATGMMvCpKAdEKWfBCgp6PYwONBrKJyXxI8Maq/8
nTTVOxArwT7pAt8O/imI6xRa9nmPp/1TAdlrv6qTOKrKPqW9ZyBud7Lm0yOtN23v
lOobA1fm//L4eG3XvVaFkm5jpbn49lD6UrUSYp7Ps7GSPL9dT/KXc4AmUQXVP3bf
DExNTqqxhqZR6EA45/PsK3nJ1OhTAs9z9AAm8WM3LrvAJy/1xZVjYRXACziksbQ9
WRRO/MgGrqxoKTOEsp+eRkQdjfyR/rVKsZCR8cSAedyqUamj1bPMq8nun0DobBBL
PRZfE2bL6yRf6NTVCEq4nA5enzfmSwNSfcS6fvq26tjlVl4mEeaATRr/7nVXDGvt
LLh2V8xYmBMeQ41tQwKaIFQSl+A2R8dYBOna+XKk4QClyU2Cl6u5VCcu/xHOx5IU
wvtisP4lfDrEC5lt0Wc469N7+667K/z+mo+rtxjDbXIQ8Xpn0VnkRhg5x0cA4uzE
Q7baH95sJTiOf55ajfF/3xzPZ9aYkvPU5UPk7FObUdAN2lh4ssrcSh86LlXf//7/
w9WN0Em4QlCnNbPwDD2jxMAdNvbnQTKFYf9fk3cjdIl+tZ7JFO5EzpBFEBucmTNj
OUIRCpFM/gwbObeCZV9QG49lYYxy/0T7N7X6Zzf7z52rkVd/WSH/PEHuNuIcF0xx
sXg0zYI3OKE1A9msHfHgN//D36XJUanPSEuSnu9cEzyMdufculSVnjls5zA7CBOd
V02NLCZHH2/X+6TTlC4CdQf7fycTv31CTipWR5dxIiVs+g5KD4eZLdAvbK22o7RW
YLW1DKNyiU3Z6YcCYR2BIwuQLNYcBPipQwr/nY+6O66lTgx3D/JfCeXRCsHo3sWm
t8yacxg3ZP0QEU1gz0RD6tPZVn1+hNkTcWLJQDD8UlCEP2Bz47y6vvdhisoIp9+Z
6tk+hfuHBDMppSHE8ihDhlAxkom8orM3AKZkYt4dDFMsUWXNbGibJdvbSoCS1d87
u7K1EeL9v5mf5QxOXpqhHAW0GZOyWMyKmfUoT2MLLqFMrgSm9FJm1swtoYAAqo1d
FGnY/ZFDAXOFgEP8aHWyTyUB2MH67aeeLyxuz/ClYz1SCADCelkiirEuE6cmHqIM
5K+hNPTpIgYlyfaZYP3hLBL+2Sdt+lmdoOYctT0ZK5MuMWBowOu5yC0zirOKr1QK
OyUSUDmwFCIDws4fTNFVdhRQOUM8s2kjxX1Ol+D0cG9qRg/aKOOePK9I6vjHvgp9
JJ2bcKWhLyjZpZO+8/hKYrnWa/qD7uLvghwzQZXWESe/dub+ZwFYW2dEMMehbaOC
G3K36qSVVI+JOajiWjIl3yIpbzQ8YxOl6CXaoCrvJ3CbOLJ5oAElS+/KtYIxr5au
a+PYY5d9c1Qr9GAARuI/FeCQ5JVk89OeKueZ26lzEC9nb7Ng+nd7l/nXdV8TH0IG
koBYZGjlC8sdz9G2H0SVcFMu555lYt63fOyHf8Agk14ZRoBTUuf4+/z2qkgjFM9a
Xh5KUt+MvC3aNI/yyjPJ/auT3mJ3CzoZlVSNVqe5e7Y8Nw/L/NrxUvGpSFdd0OLd
ODjzunbzrXr6pr3++eeG5dmMtJ/mXv8Izw/YYWqAfPajFtaWKCP/EOAf7uAYHFle
O60q31pOEeuyVNfR2kBPbU29EoX8fpDupeNTmGkL5uXZqNn5iKY5eoe148ABkNpS
jW3YqeaudGAtushbW55xfGi72P3fNZs4+qXX2v7ykGFilXjl6RgaiP/rc+DUyzut
Tqup/4Jjy1Up1jspzLbguI5Cu3hv5oz/22qtyjX8HHY8OSPI2THZmwC4hStuFRWH
ZarbuqMQJ3PLkbIwYJBXWEQHJTKrLlH4rZt+bvVAg9oUWRZaVR3MFRZIz6PlnLpL
otW9brtTOPymvFfBE31mxbji1FL5eAzmTzcz2NKCVAbAhJDyiugZjBsd/VVS22uQ
P04H9J3vpIAtt7suPLY6uFXxvuFliTyiMapXClHGrc7npGYG1NnkKBNv32itX3Zb
GoZyd6RFPmwv3725JahPDrCYCOmbucGwGroKLYaXKFVw6snend7HK1e0UUiAQisY
SLOd8DTT5WM7kIgDqIZp+5vlNGCRRkHqnYZMd8ZNCjQDLDAz2NIWfrtpIBgDXVOH
/b7dbCpvWh5eiS6kKNsqmTMyhy4gDamC2Sc+wYGbKIW3JIBhFV31AeADl1eH1fKN
AZWfnpv2PX8zV6eIZHVNgh7/Pu6qfV6MZpMUnR7JddMtLySqlqyFHO0D6QlFWPTw
TkNOpz0Q/P7jvCCKnSmV7Y2Kuq3bzk8IbNZH22yL1qpTnL9VVU/6+L17Z9RvC+J/
YxOwi3NAAI3I08FM5jPexv3V0EHgpC2M2YvAL63rrKT85i1xA5cMItqJ41CniiyZ
vbYWGnmlxIKAhxwXQQGhxcg6FFtFhRKr6bCO2JibNbegkq5N/2KgiMj8kc9g4Fxj
VkwmGnGuUlHn5gm4egTai6Xc/2YBR4/P8C7wEZBb8gNNS+Y/dr6xoOAMkxrtbHlm
eST5sPAZLpg1SZPPm5BtDMGXNpgUavUn0AoJ6zWKVnccMi2ktv6aBLXdJdZlKSRA
Oz11mKBd5ZSyDtFBW7KR6NxpFwuuv6O0ATGcUfmkEqSQ7LLpkpoHK5S4RKxHsbhb
MXm4ah49x52Xavsv+KtzYcoYxOA2IbNGo5X5Q38ZUnPwxCZRjoYbM3SORDHkbAMh
C1/nz7QWXw38i7FlN08ZvcZcRALaI7RKslfAO9rJejLKVIvSmW7X4a2HpOIlcUTu
plQEVJlyw8t5WNkqndcC0zdri6/RfZM3/XM00/lqRossrjbMvh8kdXb2eusO+Qxt
jUe71NRe9wZtcS5UTdZ0tYQZfQWcwpVheHxs5WmGdOIcuCCkyfOi0lzsqRu6+BF+
1GNSSg5Y0RIgVPxwJrrwB1CKwh2YqCxSHsvFWC5kNVwf2CjvOVAC2aba5IKKJ+s8
em1OJL0KmbQlzrf9jiXGG5EdwIpWjeotQbUDsEIgcxu4DXGYOcwQlCVBoTmtZezd
7dcxremRPVARs+gFmJbMwYkAMOY2AhSfqsOrfz1OgnqYCPRPOf/R+XIZLtKxNkdA
DdeAtl4DoLwfZfM2fRiicHEDdZhTLNBkPFYKHe7cShIcYhU50Gu1FeDzbIGTBqxb
lIbxcq+lLmf7Ybbfs6ql2TXo/748c5ElQ6yA+vvyZ6rSDV0kkeh5hHNcCzDikBen
8cdE3sMllktJiJIhVRTbS3glqcriuWq8IXAI/qNFDXN4Y3I8JNuueMsl6o5XpFqZ
hKb5+t/BM6D7W9kZ4UE3MeGT/QQVL9dLpG7ExnOd9uqxKIroXdRjkcOHDqWXUUkr
JBI+6XKugrMMnndjM8tIZLUenHUS8fxnM7zYm4AsdIaBcei/WyBMSnqIKZebYp2I
ooFuG2EDrmOZu8aS50hEONPTbnZTraNnCQTW6xZJvZpHBh5bJXYLK0ldt4gn8Nud
zqycbG3FyejQSJzd0pGECqGqCd8ntESZt+r774Z0EmHq/JCW3LAeH81Zy35l1xX7
HfZ/WaRjbsurpDo8EQ4S++/kExMbIej4b/VmmG3T26eM6txUR8bTB79FNgaRgINE
q091JQNr0/aB30IHRYo8kP5pTki+DpeqOcnyeLYSpYZloYdxuulmmZO42HmDPejR
tzpKURV6VbrAPOj89442asfN3W1JZwj9gk3F9RIgYQJU0FOkTcBwOBYMa7htO/v+
s4kJcIFUDjyHfeoD+tlxfdL3M6vry+b/JbaboCqpQefjOHas0vwZj8MwLPSqDALL
BVmwO3qI7+eBonqr2LMtyGSf4niFpQ1wogeRxhrnDvvG17lDTFUJvZSCllIGlUXr
AvNdOFQ0II7VyLxwbPS45QFIGOzA3gdkqgPxxnjmqgynOGx9/mZXQ5X6Jc5wvVxS
U3FlyA4OT3wNlPmhLhz010535E1osznO29gy2gl+LpDR7c2EMYHzz02MYsBmCvQp
z63qVk46NPQuHhdvUheABsMjcPQj2T9tNw4KjwB0sVRzbZxq0LrQnkJf5jEC/642
dPo0X9NX0Adstb7wLqUZ/g5BcyKAKOKjLEid1crxpCJx1/jlNeQdT8WzG4CLM0t/
RT85Ht/6fuUsqWXejZwqnqo3CC/IpDzLs9eZp8qdej7pDCdAzDjBPXUZrnC4muSd
dcamsIXxREPmZ7Sp0PDSzH/vCP11QEiEF+Ifig3WPQoA7tEpSg8B4l59QreKd40C
V8FRqAaExti8wpjzrS4iDAfmFMwMNGZVng4ZeaREqad7KIofHnJvtf/8C23k0yKR
GMJBb+3ZlAKukO2rxXAfPhmM1QXCPynHWhqklEYsg9Gzi7y1b26Xcc6i6ieMuD8g
erXnB8yEhThdkIEf4PjWdILQDGjpuTh3eAdKZVlbmWhurBlbSbLNd/yuoRtfV9ol
rto5fWrBBKyy6t/PGUl/I5hUxO7wYuhAc9U3vVHsKTISAiLYWapNK6sE6cav4/Mz
tJbxoLOI0KnIRBSRL9dHK/pZnGhHhX2qrtH4JEkTfzguIfgLId882CgXUxNbBhDa
q48W1RpfpgugqbfMrpGE1bFhPzo/+xzZbExmC49e5DixjquvlXyEEKnVVCGP5ygK
hbHqkwHE/PulvDL4zRsb7z9nrpI9wWUezX6yvnzh7QhO05BEk9xttNvGLASzypnk
e88n4LefsVHb46hcSINUvZle6ATq9rUZ0tZENqBd1yCmMGdEl/QLBHuNMqIsurnt
ltuvwGRDOlej+gk7+U8z+jB6P0ujmcQa9ExGCwfwmNAdswC5wsncfp++4A01RbB/
HQp/0IlUddMW5VVj+KJWAPDyZSXjehC+XkIYNKcooR77cF8ZTmsqFb6P/CMQKgIq
39k/18kMlX7BmftMy1l7+sud6fHxWEl5WsY2+jGWwCWcYhPh/3IDkRoH9fLyW3Ce
bNvsUgmHLKYLieLN2J00Fxu+ehNNa5z2MfImCrqzOk9ONqbSXuzxuJlMqqeESWUt
GELQid0rjJOLXLtiMHwgpjyn+oRtD06PxpIaa5ghNwvRDWf3rxGvFPhzlghQ75R4
bQCnIHayJ6PxIU0SLKNFIbyrIlt5p30xtVJh2L7OfjuBt7TV4LNByIHQimFmkW94
8l8wx2NWNc6pDeV82d/jWabMb98YmuD+pgD+zOvX/6bKSh/HN5bGUTjsNcXUdNjY
A4N4G8OW/ncdkFBpblF8tsy59e6leOaHquTaGYuu7jLKxTECntlVH6bz57QxiPu5
ROLIiko/NToJoNMSJ5uxUsvbDJILoDeKq2uYOkl5uKdZ78KqotNO/+6seexjTE9Z
vemC1NHQi6oqbgvJSEyMR0W/vVJROENc/7qylKOATpNO1w2/P7PrKqX9uKdgELhV
P9AqU794R0UC1WK4bxxCE+y0nTM+JiGk2qZGDX457CKynX5TdKSw0BZ3a8vfDTBs
bIxW3E6k2KlDI18hdRItbkUXZ0LUqcViVSZx8uPOQ56HZNiIwXaw0I8BQvpZEJAx
`pragma protect end_protected
`endif
`endif // GUARD_SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
dELEIwFqGdx0vYr3oabhbJwFQsK5BH7JUQpS3j/a/HBIEPXmaQQVunHsCzu8VF0E
I/pxYVPEOxEuhQy4/Yhb6b8goua13t9jnwFHiHuYXrg+z7O5Dfu5wDAyR3w1pNQV
Vy8/oalPGkK2Z2ZhXjSsguhMTOoWZ/em5VvMU4n/qc0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 20140     )
SCM/M9rqyAH4iWgKKGlKPD8fFT52uoRuClGrdAEJaMOt7Hl47fovhULbrl0dfxDW
LsiqjI9cVwNvHjFmDGhtpMn+m0umxp34r+kIN0zzY0oqHiSQzG/gr4pp3pQcbDBM
`pragma protect end_protected
