
`ifndef GUARD_SVT_AXI_PORT_MONITOR_COMMON_SV
`define GUARD_SVT_AXI_PORT_MONITOR_COMMON_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi" 
`endif
`include "svt_axi_defines.svi"

//vcs_lic_vip_protect
  `protected
8.FM.c2NMHBTV55X&M81R>TM-9BU@_L.Xe]Q8338f9XY:4g,6C>=((LG\+0W=5FB
/X>0b[)c-SR7:5;P[J:UW6M4_QcY__C8+6EHeB>aVdUEO?^K=HTD;.ec.EcT<1<0
P2W2,a=30=GE2]/4S88g=RI+,]<-O<L4K-R/T?[N2OC.)V/393)-XV7a=(N.\g.@
[2S1U=&b52LB=C00XE6D636YU4FDP)YY)e6_9\[f00<\=:A^f?V\-0B@HR2+#B1M
A1MdfAM5859XcQTJ/F[3DX&_&HM[Z:58(3K)S,&.G13f48G(,;7cfeg[F1Hg#U@E
@:8]F+QWI/8a^50JRfL#,g)6.@HJNfT\GM8I;1)6^:>-];#SfYN7=QFfe2@g9[8:
SH(L@ZN&<M9?PO\)N5b(Ge+;KWFV2.V#S8A=XHKAEH1I@39+&C^^G\;_AG@RRbFO
Z;/_MXK2_0FKUWEDSN>QVcK_P@<TcV&b2@GB)HW=FW@53S_3GFegDd--Cf<F7b;P
_=YZQ=;.SINQ[f?gETc4,854F7cXR,>AADTFD]d2V.;CdB6eULfe@Rd[0]Y>eRRI
eC<GQ8-,=2&TZS/X8Ua/-[-PUYaA=JCG0cC7:9,PXJEBUHO:H4MF#(DV8@93T]?M
+g_406Z2;6aca(G,5WL#^4FcIS&[Z.A4/(F;^A^/b;1[5DS\SW50MB_FGTOD6c()
HMg]b(S:L-/b;O),e?6Z7M2J,:F4b:JdJ=9^PKF/CNd-FRV8GQ2M^4SYZ#Nff1[^
PPMa5LGG7,N2GMR2^?dMT3:8K#UOK;F]LM?7KF=EZ9J;:&aOg2X[gb:B8]eG2#)F
3^@\dZ+/6f5gKZ>S:O3FYHF)CgM[JMAR>4aC#9[@#(dZBM_A6b>C#\<BLY_dcTbL
AdGPPgP)TH8dLa)B;Pd:agAL0f\Z8X3AL4@fa15T/O/^-6aU7>B^AT@]/@R>;4=O
OXHXM/MDeb>:b,LVZ_ObL-L<KDbHXN?GP1+[0aK9>aGN@;JXc5E5?C_PPf]28W=B
ca.9NY>5FGG)beA&I;F?XUe85/FA^08XTVG_JAGbLdcS/<d#TEO6V)eOT@3Ea#AL
\F_K,/9VGg9=79K=VP8,\H/g<D_AQ<eeQ[<\3&4#(b0gTQBKU.>:AHB1bSWO8deg
1BPbG[9I;UTcB4M@bDKc,0\RR/AAf+VH(bO^-9WWI>T+>TK(Z_b.b#/O6]f-U&/E
Q-c(O9P_U=;/^:3+=]5I6])=E;EcMa9K;(=e,B0/,T-9)2:G&F=5H^Q#-GT)3-JM
6?.G]d0>XgN49=F5H?+<[M63/QgGXO6-5&(Q?S[H7CX;AYO#\?Z.L;MN[,cD#C-D
#WJ8MW6/AP>O9=<@H>;)[Ze;,A85EDLFL49JJ3:Bf:L.81<f>.067P.c72TO-@2.
-(E=1O/\bQ+PcO=0aI8M1>8NLba@dUL7<XTQK9(Q..8:<;M\-OP5_#gaLQ6L+EA0
\G1)MOVFLG>5U]E@g=M=)1DAM+QI1dT+6\.aC3VNO+ESF<e\?M0B+[?6&TW?J#ED
U:YRXOJ/WVe\Q<NAaIM0MPZ<)Y,bGJFII=DLTaZ_QZD)<Kb\R>@]eJX:UFeW8P]9
65+U):);/7Q(d;(PLWWSE:B/BLg[e&Q4<HXH@+YU.C@BN@04dfaFZ8/;dL@>7Pc2
[aYP&=B+P+U2IDH.cM:6(bO15].<I(Y6.1@X,SaaRX4J-7GS8M>W#N_=S7E2OW+g
-W4\04-Y)5KN=^=S0_gVa3J1<3_:6X(dEQ,9>2I25/)AW>Y:QB=dAN;4eL^:C:5J
GEO^&]Z;&A):.gHaG)0ebNZYeN+3]B7Jde3N@LdPd]P(]52S041#R]-dE@TP\UUM
OQ_)PUIY19gD;24/Z&>I;e[@H+1,IfdS&HT0Y4e5QfX>M\O]:4R+\=(C,gVQ,+)Y
a6_&RN6=2)IG2TKc+0=&Yf<6<AUXcZBb:e[f<5O(IC/=--NZ_VNAD/e4_Ee_I9A,
/O2=>e>4I/+TbDY;?JEd.X56ZMYQS0BTV?WV1>POZ_;+7VE=;TE?d;c889&+(K9]
ef&:/5_V(=&>c\)ASTU^L3g(3GRfC#(^db(GA6db-1@/bLG@L4J3MP[]^DHQJ]A?
fSK;J;)K#JG>0$
`endprotected
   
   

/** @cond PRIVATE */
typedef class svt_axi_checker;
typedef class svt_axi_port_monitor;
//typedef class svt_axi_cache_monitor_common;
`ifdef SVT_VMM_TECHNOLOGY
typedef class svt_axi_master_group;
`else
typedef class svt_axi_master_agent;
`endif

`ifndef SVT_AXI_DISABLE_DEBUG_PORTS
class svt_axi_port_monitor_common#(type MONITOR_MP=virtual `SVT_AXI_SLAVE_IF.svt_axi_monitor_modport,
                                   type DEBUG_MP=virtual `SVT_AXI_SLAVE_IF.svt_axi_debug_modport) extends svt_axi_common;
`else
class svt_axi_port_monitor_common#(type MONITOR_MP=virtual `SVT_AXI_SLAVE_IF.svt_axi_monitor_modport) extends svt_axi_common;
`endif

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************
  /** Custom type definition for virtual AXI interface */
  typedef virtual svt_axi_stream_if.svt_axi_stream_monitor_modport STREAM_MONITOR_MP;


  // ****************************************************************************
  //vcs_lic_vip_protect
`protected
K4cfWDEd\X15P5S?TDcBf?c^cTJ4Sf]W>Da_N3.<\LQXAKK6P/Y;)(0W);KR7TbM
Ag3398]@eKDX]P/1-,Q[O36>^[93.[@4cQBL#=)>&ZIV#D3KA\2DMXOcgJ_f8=:b
:F5G^3/7IbC1ZA-C.D4FN6aF/POM9YB&c45Ac2@.(5Td8>Jg3A:K,?M5aa8,T,P&
@_Pc\X4=P,Z4c/&I76M[A^[=>&Sd4f>K&L)H9ZN,P9<&<a5F4eQPY(WHV=NgRZ6a
YVV]P;),:HWeUO#^CU,\(V6J,5,E.LQ?1@O.Q?5fRXEfX@I@gRd5N9gU107U/?Tf
dF_Y9,P_O<#P]173_8)#)7C,?.M2KW]gb2dV1V=?U7/AZMKa_b[G/-5=Ka>f)PPW
42T#&Le[3NIe2[<B<eY(QO4V4<gY5I2d3ATHb_)]165(JKAE@\efGN=#H\eLENJS
2E1b5A^9.+(@7K7,J6bODLgNE>3+d8C4^UJgYe5W5L_;13.bHf2&fD0CX,GVJ?1e
1<>@&C68=_.;0C1-PE#SUQXb4>Ma\4EFT?g(a,K=_&HG/S3O:W=6?=/Ma2FRI;-V
F@_U&]08Q0&Q9TaH__MUY9^/gPET0SN_VMeN)ONe6R2L19>IV[]WJU0X-<+R?Q.F
FPeI/)@7Cd<E0/E?(9-9/Z?)VM40ZWAE<2D]FU.A@ZNQ>I)?M\7Q@>A=^DR)DW06
1f]1MB(G3He[=K._ZV:09&N?=3?KWbA2b#4QXDFPQ>[(E=,QR\<SH,0&U1[RN<A0
W)U@SN+g&XQfU3E5?I@0M#\HR3UDE564]&bPTRA)J3/b>PIaUSeg/8R?RW#2/]R_
;L8/5<TI#])dO;>.UNgBSO\-WAbI.J3D[Vd.D21a2=-KYQSZ-NEBO-GKVdWAR<^C
D#1&N/6EFcdA^2PV[T(0OB]INdE0d71<XSKU1E12T,=J<85&#ZfZTaJcZReV0/5N
-GbN_?EIT+D55V4&;SQZLOe/3]05F6T9JYfO[C9>g]NW-3U^<XDCeDT?UNFbdPb_
-RU4ITReN,DIO+Y=ag864&ZIOIP:6TVE7JJ]YB::7BaW;0&YRLTR3#6QE&]f,/=a
#</BT<JEa4b9H3(NdV3?-55,2fVX+dE7J&aE8XYA\9>^H)O/<ZaU-c4?2[fN0S@2
]d93P+7IaSacdae<;ME_=R\FA/.P;==.7<,M5X/CK2,CSS4R53;RVe&a_L;@fUDJ
LL)+G/ZH8?ML\RXX[:F-U?2)FZ9V_YS>7JK,fXg(LfUZK_DK&Jc631@?O47DY[ZW
TFa::=T#VDS7M_9]C2(Y6QQ7Jg^;5IKGW3K<V</=]H.g-T.LU\^;^^g#/b5YF:?4
NG<W9KX54/;&8?PMG-IR+=]^K_d@3^2MZZZ6\1-,BCgA1GIWF5-g+X._(4Z+G-<<
e2GUTL>53:(E8./C-2f)SSXeOZ&^QLEY+0:G[]-BA.D6DNR)aec;G,5#986W3ba0
+=;UX5BR7BP?OeT/9#TH,9G:Z1OJ(]PP<$
`endprotected



  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
 //svt_axi_checker axi_checker;
   svt_axi_port_monitor axi_port_monitor;

   svt_axi_cache_monitor_common passive_cache_monitor;
  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Master VIP modport */
  protected MONITOR_MP monitor_mp;
  protected STREAM_MONITOR_MP stream_monitor_mp;
`ifndef SVT_AXI_DISABLE_DEBUG_PORTS
  protected DEBUG_MP debug_mp;
`endif

  /** Factory used to create transactions. */
  svt_axi_transaction xact_factory = null;

  // ****************************************************************************
  // protected Data Properties
  // ****************************************************************************
  /** @cond PRIVATE */
   // NC gives this error for these declarations (not currently supported)
  // Associative array uses an element data type that is not currently supported [SystemVerilog]
`ifndef INCA
  /** Associative array of the receive_read_addr process indexed by
    * the transaction handle */ 
  protected process receive_read_addr_proc_q [svt_axi_transaction];

  /** Associative array of the receive_read_data process indexed by
    * the transaction handle */ 
  protected process receive_read_data_proc_q [svt_axi_transaction];

  /** Associative array of the receive_write_addr process indexed by
    * the transaction handle */ 
  protected process receive_write_addr_proc_q [svt_axi_transaction];

  /** Associative array of the receive_write_data process indexed by
    * the transaction handle */ 
  protected process receive_write_data_proc_q [svt_axi_transaction];

  /** Associative array of the receive_write_resp process indexed by
    * the transaction handle */ 
  protected process receive_write_resp_proc_q[svt_axi_transaction];

  /** Associative array of the receive_snoop_addr process indexed by
    * the transaction handle */ 
  protected process receive_snoop_addr_proc_q [svt_axi_snoop_transaction];

  /** Associative array of the receive_snoop_data process indexed by
    * the transaction handle */ 
  protected process receive_snoop_data_proc_q [svt_axi_snoop_transaction];

  /** Associative array of the receive_snoop_resp process indexed by
    * the transaction handle */ 
  protected process receive_snoop_resp_proc_q[svt_axi_snoop_transaction];

  /** Associative array of the receive_data_stream process indexed by
    * the transaction handle */ 
  protected process receive_data_stream_proc_q[svt_axi_transaction];
`endif

  /** Internal queue of active transactions */
  protected svt_axi_transaction active_xact_queue[$];
  
   /** Internal queue of active transactions */
  protected svt_axi_transaction active_memory_update_queue[$];

 /** Internal queue of active snoop transactions */
  protected svt_axi_snoop_transaction active_snoop_xact_queue[$];
  
  /** Internal queue of transactions in locked sequence */
  protected svt_axi_transaction locked_xact_queue[$];

  /** Mask for valid bytes on read data */
  bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] curr_read_data_mask;

   /** Mask for valid bytes on read poison */
  bit[`SVT_AXI_MAX_POISON_WIDTH-1:0] curr_read_poison_mask;
  
  /** Internal queue to store write transactions in the order in which address is recieved*/
  protected svt_axi_transaction  write_addr_order_xacts[$];

  /** Internal queue to store write transactions in the order in which data is received*/
  protected svt_axi_transaction  write_data_order_xacts[$];

 /** The cycle in which last arvalid was driven high*/
  //protected int last_arvalid_cycle = 0;

  /** The cycle in which last arready was sampled high*/
  //protected int last_arready_cycle = 0;

  /** The cycle in which last awvalid was driven high*/
  //protected int last_awvalid_cycle = 0;

  /** The cycle in which last awready was sampled high*/
  //protected int last_awready_cycle = 0;

  /** The cycle in which last wvalid was driven high*/
  //protected int last_wvalid_cycle = 0;

  /** The cycle in which last wready was sampled high*/
  //protected int last_wready_cycle = 0;

  /** The cycle in which last rvalid was sampled high*/
  //protected int last_rvalid_cycle = 0;

  /** The cycle in which last rready was sampled high*/
  //protected int last_rready_cycle = 0;

  /** The cycle in which last bvalid was sampled high*/
  //protected int last_bvalid_cycle = 0;

  /** The cycle in which last bready was driven high*/
  //protected int last_bready_cycle = 0;

  /** log_base_2 of data width in bytes */
  protected int log_base_2_data_width_in_bytes;

  /** data width in bytes */
  protected int data_width_in_bytes;

  /** Internal clock count from arvalid to arready.*/
  protected int arvalid_to_arready_delay;
  
  /** Internal clock count from rvalid to rready.*/
  protected int rvalid_to_rready_delay;
  
  /** Internal clock count from awvalid to awready.*/
  protected int awvalid_to_awready_delay;
  
  /** Internal clock count from wvalid to wready.*/
  protected int wvalid_to_wready_delay;
  
  /** Internal clock count from bvalid to bready.*/
  protected int bvalid_to_bready_delay;

  /** mask used for sampling data based on data_width*/
  protected bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] sample_data_mask;

  /** mask used for sampling tdata based on tdata_width*/
  protected bit[`SVT_AXI_MAX_TDATA_WIDTH-1:0] sample_tdata_mask;

   /** mask used for sampling poison based on data_width*/
  protected bit[`SVT_AXI_MAX_POISON_WIDTH-1:0] sample_poison_mask;

 /** mask used for sampling data_user based on data_user_width*/
  protected bit[`SVT_AXI_MAX_DATA_USER_WIDTH-1 :0] sample_data_user_mask;

 /** mask used for sampling tuser based on tuser_width*/
  protected bit[`SVT_AXI_MAX_TUSER_WIDTH-1 :0] sample_tuser_mask;
    
  /** mask used for sampling data based on data_width*/
  protected bit[`SVT_AXI_ACE_SNOOP_DATA_WIDTH-1:0] sample_snoopdata_mask;

 /** mask used for sampling poison based on data_width*/
  protected bit[`SVT_AXI_ACE_SNOOP_POISON_WIDTH-1:0] sample_snoop_poison_mask;

  /** mask used for sampling addr based on addr_width*/
  protected bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] sample_addr_mask;

  /** mask used for sampling addr_user based on addr_user_width*/
  protected bit[`SVT_AXI_MAX_ADDR_USER_WIDTH-1 :0] sample_addr_user_mask;
  
  /** mask used for sampling addr based on snoop_addr_width*/
  protected bit[`SVT_AXI_ACE_SNOOP_ADDR_WIDTH-1:0] sample_snoopaddr_mask;

  /** mask used for sampling ID based on id_width*/
  protected bit[`SVT_AXI_MAX_ID_WIDTH-1:0] sample_id_mask;

  /** mask used for sampling TID based on tid_width*/
  protected bit[`SVT_AXI_MAX_TID_WIDTH-1:0] sample_tid_mask;

  /** mask used for sampling ARID and RID based on read_chan_id_width*/
  protected bit[`SVT_AXI_MAX_ID_WIDTH-1:0] sample_read_id_mask;

  /** mask used for sampling AWID,WID and BID based on write_chan_id_width*/
  protected bit[`SVT_AXI_MAX_ID_WIDTH-1:0] sample_write_id_mask;

  /** mask used for sampling addr based on resp_user_width*/
  protected bit[`SVT_AXI_MAX_BRESP_USER_WIDTH-1:0] sample_resp_user_mask;
  
  /** mask used for sampling tdest based on tdest_width*/
  protected bit[`SVT_AXI_MAX_TDEST_WIDTH-1:0] sample_tdest_mask;

  /** Variable that stores the read transaction count */
  protected int read_xact_count = 0;

  /** Variable that stores the DVM complete transaction count */
  protected static int dvm_complete_count[];

  /** Variable that stores the DVM Snoop sync's count */
  protected static int dvm_sync_count[];
 
  /** Variable that stores the stream transaction count */
  protected int stream_xact_count = 0;

  /** Variable that stores the write transaction count */
  protected int write_xact_count = `SVT_AXI_WRITE_XACT_COUNT_BASE;
  
  /** Variable that stores the snoop transaction count */
  protected int snoop_xact_count = 0;

  /** this flag is set when reset is asserted synchronous or asynchronously */
  protected bit dynamic_reset_flag = 0;

  /** log_base_2 of cache_line_size */
  protected int log_base_2_cache_line_size;

  // ****************************************************************************
  // EVENTS 
  // ****************************************************************************
  /** Event that indicates that ARREADY is received */
  protected event arready_received;
  
  /** Event that indicates that ACREADY is received */
  protected event acready_received;

  /** Event that indicates that RREADY is received */
  protected event rready_received;

  /** Event that indicates that AWREADY is received */
  protected event awready_received;

  /** Event that indicates that WREADY is received */
  protected event wready_received;

  /** Event that indicates that BREADY is received */
  protected event bready_received;
  
  /** Event that indicates that CDREADY is received */
  protected event cdready_received;
  
  /** Event that indicates that CRREADY is received */
  protected event crready_received;
  
  /** Event that indicates that RACK is received */
  protected event rack_received;
  
  /** Event that indicates that WACK is received */
  protected event wack_received;

  /** Event that indicates that TREADY is received */
  protected event tready_received;

  /** Event that is triggered when the process that waits for AWVALID has started */
  protected event ev_wait_for_awvalid;

  /** Event that is triggered when the process that waits for WVALID has started */
  protected event ev_wait_for_wvalid;

  /** Event that is triggered when the process that waits for TVALID has started */
  protected event ev_wait_for_tvalid;

  /** Event that is triggered when the process receive_snoop_addr has started */
  protected event ev_snoop_addr_started;

  /** Event that is triggered when the process receive_snoop_resp has started */
  protected event ev_snoop_resp_started;

  /** Event that is triggered when the process receive_snoop_data has started */
  protected event ev_snoop_data_started;

  /** Event that is triggered when we have entered receive_read_addr task*/
  protected event ev_receive_read_addr;

  /** Event that is triggered after every sample. Other processes synchronize with
    * this event to ensure that all signals are sampled. Note that if a reset is in
    * progress, the reset_received event is triggered prior to this event. This will
    * ensure that processes that are synchronized with this event will be terminated
    * at reset.
    */
  protected event is_sampled;

`ifdef SVT_AXI_QVN_ENABLE
  /**
    * Each master needs at least one QVN Token to be available for a particular Virtual Network
    * in order to make a transfer to an Axi Channel targeted to same VN. For this purpose, each
    * master needs to keep track of each Token it has requested, granted, when it was granted,
    * tokens that remain unused and remove a token when it has been used to make a transfer.
    * It also contains semaphore for getting token statistics and requesting a token consuming time.
    *
    * Following QVN Token object queue (one for each Virtual Network) is used for Read Address Channel
    */
  protected qvn_token_pool qvn_read_addr_token_pool_of_vn[int];

  /**
    * Following QVN Token object queue (one for each Virtual Network) is used for Write Address Channel
    */
  protected qvn_token_pool qvn_write_addr_token_pool_of_vn[int];

  /**
    * Following QVN Token object queue (one for each Virtual Network) is used for Write Data Channel
    */
  protected qvn_token_pool qvn_write_data_token_pool_of_vn[int];


  protected logic previous_arvalid;
  protected logic previous_arready;
  
  protected logic previous_awvalid;
  protected logic previous_awready;

  protected logic previous_wvalid;
  protected logic previous_wready;

  /**
    * Flage to prevent call to process_qvn_reset() for every clock of reset 
    */  
  protected bit  process_qvn_reset_called;
 
`endif
   
      

   // ****************************************************************************
  // SEMAPHORES
  // ****************************************************************************
  /** Semaphore that controls access to the active xact queue. */
  protected semaphore active_xact_queue_sema;
 
  /** Semaphore that controls access to the active xact queue. */
  protected semaphore active_memory_update_queue_sema;
 
  /** Semaphore that controls access to the active snoop xact queue. */
  protected semaphore active_snoop_xact_queue_sema;
  
  /** Semaphore that controls access to the barrier xact queue. */
  protected semaphore barrier_xact_queue_sema;

  // ****************************************************************************
  // TIMERS 
  // ****************************************************************************
  /** Timer that monitors arready assertion */
  svt_timer arvalid_arready_timer;

  /** Timer that monitors rready assertion */
  svt_timer rvalid_rready_timer;

  /** Timer that monitors awready assertion */
  svt_timer awvalid_awready_timer;

  /** Timer that monitors wready assertion */
  svt_timer wvalid_wready_timer;

  /** Timer that monitors bready assertion */
  svt_timer bvalid_bready_timer;
  
  /** Timer that monitors acready assertion */
  svt_timer acvalid_acready_timer;
  
  /** Timer that monitors crready assertion */
  svt_timer crvalid_crready_timer;
  
  /** Timer that monitors cdready assertion */
  svt_timer cdvalid_cdready_timer;

  /** Timer that monitors tready assertion */
  svt_timer tvalid_tready_timer;


  local bit passive_cache_monitor_enable = 0;
  local int wr_count=0, rd_count=0, snp_count=0;
 
  local svt_axi_transaction local_xact;

  /** Master Transaction */
  svt_axi_transaction global_parity_xact;

  /** @endcond */
  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (svt_axi_port_configuration cfg, uvm_report_object reporter);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param reporter OVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (svt_axi_port_configuration cfg, ovm_report_object reporter);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_axi_port_configuration cfg, svt_xactor xactor);
`endif
 
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);
  
  /** Called in order to construct a new svt_axi_transaction object using a local
   * factory */
  extern virtual function void create_axi_xact (svt_axi_port_configuration cfg,ref svt_axi_transaction xact,ref svt_axi_transaction xact_factory);

  /**
   * If reset happens before the transaction is added to the add_to_active queue
   * the transaction is aborted and written to the analysis port.
   */
  extern virtual task process_reset_for_new_transaction(svt_axi_transaction xact);

  /** 
    * Adds the transaction to the internal queue. 
    */
  extern virtual task add_to_active(svt_axi_transaction xact);

  /** 
    * Removes transaction xact from the internal queue. 
    */
  extern virtual task remove_from_active(svt_axi_transaction xact);


  /** 
    * Removes transaction xact from the internal queue. 
    */
  extern virtual task remove_from_memory_update_queue(svt_axi_transaction xact);


  /** Receives read address */
  extern virtual task receive_read_addr(svt_axi_transaction xact);

  /** Receives read data */
  extern virtual task receive_read_data(svt_axi_transaction xact);

  /** Receives read data */
  extern virtual task receive_read_chunk_data(svt_axi_transaction xact);

  /** Receives write address */
  extern virtual task receive_write_addr(svt_axi_transaction xact);

  /** Receives write data */
  extern virtual task receive_write_data(svt_axi_transaction xact);

  /** Receives write response */
  extern virtual task receive_write_resp(svt_axi_transaction xact);

`ifdef SVT_AXI_QVN_ENABLE
  extern virtual task process_qvn_reset(bit initial_reset);
  extern virtual task process_qvn_token_handshake_signals();
  extern virtual task perform_read_addr_channel_qvn_checks(logic [3:0] arvnet_val, logic arvalid_val, logic arready_val, bit arbar_bit0, logic [`SVT_AXI_MAX_ID_WIDTH - 1:0] arid_val);
  extern virtual task perform_write_addr_channel_qvn_checks(logic [3:0] awvnet_val, logic awvalid_val, logic awready_val, bit awbar_bit0, logic [`SVT_AXI_MAX_ID_WIDTH - 1:0] awid_val);
  extern virtual task perform_write_data_channel_qvn_checks(logic [3:0] wvnet_val, logic wvalid_val, logic wready_val);
  extern virtual task check_token_availability_for_vn(logic [3:0] vnet_val, string channel_name, output bit token_available);
  extern virtual task check_slave_wr_addr_max_outstanding_token(logic [3:0] vnet_id);
  extern virtual task check_slave_wr_data_max_outstanding_token(logic [3:0] vnet_id);
  extern virtual task check_slave_rd_addr_max_outstanding_token(logic [3:0] vnet_id);
`endif

    extern virtual task process_read_addr_channel(ref int arvalid_to_arready_delay,
                                          output svt_axi_transaction curr_read_addr_xact);

    extern virtual task process_read_data_channel(ref int rvalid_to_rready_delay,
                                          output svt_axi_transaction curr_read_data_xact);

    extern virtual task process_write_addr_channel(ref int awvalid_to_awready_delay,
                                           output svt_axi_transaction curr_write_addr_xact);

    extern virtual task process_write_data_channel(ref int wvalid_to_wready_delay,
                                           output svt_axi_transaction curr_write_data_xact,
                                           input svt_axi_transaction curr_write_addr_xact);

    extern virtual task process_write_resp_channel(ref int bvalid_to_bready_delay,
                                         output svt_axi_transaction curr_write_resp_xact);

  /** Processes signals in the data stream channel */
  extern virtual task process_data_stream_signals(ref int tvalid_to_tready_delay, output svt_axi_transaction curr_data_stream_xact);
  
  /** function that compares the expected and configured RRESP for exclusive
   * read transactions */
  extern virtual function void perform_exclusive_read_resp_checks(svt_axi_transaction excl_resp_xact);
  
  /** It monitors the response for exclusive read transaction */
  extern virtual function void process_exclusive_read_response(svt_axi_transaction excl_resp_xact, input bit excl_read_error);
  
  /** function that compares the expected and configured BRESP for exclusive
   * write transactions */
  extern virtual function void perform_exclusive_write_resp_checks(svt_axi_transaction excl_resp_xact);
  
  /** Waits for exclusive write transaction after exclusive read*/
  extern virtual task wait_for_exclusive_write(svt_axi_transaction xact);

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Advances clock */
  extern virtual task advance_clock(int num_clocks);

  /** Reports end-of-simulation summary report, checks etc */
  extern virtual function void report();

  /** Samples the reset signal */
  extern virtual task sample_reset();
   /**samples initial reset async*/
   extern virtual task sample_reset_async();

   extern virtual function void detect_initial_reset();

  /**Performs checks related to reset and update variables*/
  extern virtual task process_initial_reset();

  /** Perform reset related checks*/
  extern virtual task perform_reset_checks();

  /** task to sample parity check signals and calculate respective signal parity values for parity check comparision */
  extern virtual task sample_and_check_parity_check_signal();
  
  /** Waits until rvalid corresponding to xact is received */
  extern virtual task wait_for_rvalid(svt_axi_transaction xact);
  
  /** Waits for rdata */
  extern virtual task wait_for_rdata(svt_axi_transaction xact);

  /** Waits until awvalid corresponding to xact is received */
  extern virtual task wait_for_awvalid(svt_axi_transaction xact);
  
  /** Waits for awaddr */
  extern virtual task wait_for_awaddr(svt_axi_transaction xact);

  /** Waits until wvalid corresponding to xact is received */
  extern virtual task wait_for_wvalid(svt_axi_transaction xact);

  /** Waits for wdata */
  extern virtual task wait_for_wdata(svt_axi_transaction xact);

  /** Waits until bvalid corresponding to xact is received */
  extern virtual task wait_for_bvalid(svt_axi_transaction xact);

  /** Waits until bvalid with the id of this transaction is received */
  extern virtual task wait_for_bresp(svt_axi_transaction xact);
  
  /** Sets the configuration */
  extern virtual function void set_cfg(svt_axi_port_configuration cfg);

  /** Utility task to set internal variables */
  extern virtual function void set_internal_variables(svt_axi_port_configuration cfg);

  /** Constructs the timers used */
  extern virtual function void create_timers();

  /** Waits for awready assertion. Times out based on the awvalid-awready timeout */
  extern virtual task wait_for_awready(svt_axi_transaction xact);

  /** Waits for wready assertion. Times out based on the wvalid-wready timeout */
  extern virtual task wait_for_wready(svt_axi_transaction xact);

  /** Waits for bready assertion. Times out based on the bvalid-bready timeout */
  extern virtual task wait_for_bready(svt_axi_transaction xact);
  
  /** Waits for arready assertion. Times out based on the arvalid-arready timeout */
  extern virtual task wait_for_arready(svt_axi_transaction xact);

  /** Waits for rready assertion. Times out based on the rvalid-rready timeout */
  extern virtual task wait_for_rready(svt_axi_transaction xact);
  
  /** 
    * Resizes arrays and aligns data based on the address. 
    * Used in data_before_addr scenario, where information needed for
    * size of arrays of alignment of data is received only after the data
    * is received
    */ 
  extern virtual function void resize_and_align_data(svt_axi_transaction xact);
 
  /** Writes data into a shadow memory */
  extern virtual task write_data_to_mem(svt_axi_transaction xact);

  /**
    * Creates the transaction inactivity timer
    */
  extern virtual function svt_timer create_xact_inactivity_timer();

  // ACE RELATED METHODS
  /** 
    * Adds the snoop transaction to the internal queue. 
    */
  extern virtual task add_to_snoop_active(svt_axi_snoop_transaction xact);

  /** 
    * Removes snoop transaction xact from the internal queue. 
    */
  extern virtual task remove_from_snoop_active(svt_axi_snoop_transaction xact);

  /** Receives snoop address */
  extern virtual task receive_snoop_addr(svt_axi_snoop_transaction xact);

  /** Receives snoop data */
  extern virtual task receive_snoop_data(svt_axi_snoop_transaction xact);

  /** Receives snoop response */
  extern virtual task receive_snoop_resp(svt_axi_snoop_transaction xact);

  extern virtual task process_snoop_addr_channel(ref int acvalid_to_acready_delay,
                                         output svt_axi_snoop_transaction curr_snp_addr_xact);

  extern virtual task process_snoop_resp_channel(ref int crvalid_to_crready_delay,
                                         output svt_axi_snoop_transaction curr_snp_resp_xact);

  extern virtual task process_snoop_data_channel(ref int cdvalid_to_cdready_delay,
                                         input svt_axi_snoop_transaction curr_snp_resp_xact,
                                         output svt_axi_snoop_transaction curr_snp_data_xact);

  /** Waits until cdvalid corresponding to snoop xact is received */
  extern virtual task wait_for_cdvalid(svt_axi_snoop_transaction xact);
  
  /** Waits until crvalid corresponding to snoop xact is received */
  extern virtual task wait_for_crvalid(svt_axi_snoop_transaction xact);

  /** Waits for rack assertion. Times out based on the rack timeout */
  extern virtual task wait_for_rack(svt_axi_transaction xact);
  
  /** Waits for wack assertion. Times out based on the wack timeout */
  extern virtual task wait_for_wack(svt_axi_transaction xact);

  /** Waits for acready assertion. Times out based on the acvalid-acready timeout */
  extern virtual task wait_for_acready(svt_axi_snoop_transaction xact);
  
  /** Waits for crready assertion. Times out based on the crvalid-crready timeout */
  extern virtual task wait_for_crready(svt_axi_snoop_transaction xact);
  
  /** Waits for cdready assertion. Times out based on the cdvalid-cdready timeout */
  extern virtual task wait_for_cdready(svt_axi_snoop_transaction xact);

  /** Checks if there is a snoop to the same cache line addressed by xact */
  extern virtual function svt_axi_snoop_transaction check_snoop_to_same_cache_line(svt_axi_transaction xact, output bit is_snoop_to_same_cache_line);

  /** Checks if there is a resp to the same cache line addressed by xact */
  extern virtual function svt_axi_transaction check_resp_to_same_cache_line(svt_axi_snoop_transaction xact, output bit is_resp_to_same_cache_line);

  /** Checks if this is a barrier transaction */
  extern virtual function bit is_write_barrier_or_evict(logic [`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] awsnoop, logic [`SVT_AXI_ACE_BARRIER_WIDTH-1:0]  awbar); 

`ifdef SVT_ACE5_ENABLE
/** Checks if this is a STASHONCEUNIQUE or STASHONCESHARED transaction */
  extern virtual function bit is_stashonceshared_or_stashonceunique(logic [`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] awsnoop, logic [`SVT_AXI_ACE_BARRIER_WIDTH-1:0]  awbar); 
`endif

  /** Triggers events for snoop processing based on sampled signals */
  extern virtual task trigger_snoop_events(svt_axi_snoop_transaction curr_snp_addr_xact,
                                           svt_axi_snoop_transaction curr_snp_resp_xact,
                                           svt_axi_snoop_transaction curr_snp_data_xact);

  /** Waits for active threads working on snoop transctions to terminate */
  `ifndef INCA
  extern virtual task wait_for_active_snoop_threads_to_terminate();
  `endif

  /** Processes reset for ACE related transactions */
  extern virtual task process_ace_reset();

  /** Sample ACE read address channel signals */
  extern virtual task sample_ace_read_addr_chan_signals(
                                ref logic [`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop,
                                ref logic [`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar,
                                ref logic [`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_ardomain
                      );

  /** Sample ACE write address channel signals */
  extern virtual task sample_ace_write_addr_chan_signals(
                                ref logic [`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] observed_awsnoop,
                                ref logic [`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_awbar,
                                ref logic [`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_awdomain,
`ifdef SVT_ACE5_ENABLE
                                ref logic[`SVT_AXI_STASH_NID_WIDTH-1:0]observed_stash_nid,
                                ref logic[`SVT_AXI_STASH_LPID_WIDTH-1:0]observed_stash_lpid,
                                ref logic observed_stash_nid_valid,
                                ref logic observed_stash_lpid_valid,
`endif

                                ref logic observed_awunique
                      );

  /** Samples rack */
  extern virtual task sample_rack(ref logic observed_rack);

  /** Samples wack */
  extern virtual task sample_wack(ref logic observed_wack);

  extern virtual task wait_for_tvalid(svt_axi_transaction xact);

  /** Task that controls reception of data stream signals */
  extern virtual task receive_data_stream(svt_axi_transaction xact);

  /** Waits for assertion of tready */
 extern task wait_for_tready(svt_axi_transaction xact);

 /** Performs checks on locked transactions */
 extern task check_locked_xact_sequence(svt_axi_transaction curr_locked_xacts[$]);

 /** Pushes external coherent transaction to the port monitor */
 extern virtual task push_external_coherent_xact(svt_axi_transaction xact);

 /** Pushes external snoop transaction to the port monitor */
 extern virtual task push_external_snoop_xact(svt_axi_snoop_transaction xact);
 
 /** Task for setting update_mem_in_req_order field */ 
 extern virtual task set_update_mem_in_req_order_field(svt_axi_transaction xact);

  /** 
    * Returns the number of READ transcations that have started and
    * in active queue 
    */
  extern virtual function int get_num_started_read_xacts();

  /** 
    * Returns the number of WRITE transcations that have started and
    * in active queue 
    */
  extern virtual function int get_num_started_write_xacts();

`ifdef SVT_ACE5_ENABLE
 /** 
    * Returns the number of WRITE transcations that have started  and in 
    * active queue
    */
  extern virtual function int get_num_started_atomic_xacts ();
`endif

 /**
   * Checks if the number of outstanding transactions send by the master are not more than the configured max value
   */
  extern virtual function void get_num_outstanding_xacts(output int total_outstanding_xacts, output int num_rd_outstanding_xacts, output int num_wr_outstanding_xacts,output int num_atomic_outstanding_xacts);
 
 /**
   * Gets the handle of the active transaction queue to be used by other components.
   */
 extern virtual function void get_active_transaction_queue_handle(output svt_axi_transaction active_trans_queue[]);

  /** Processes RACK */
  extern task process_rack();

  /** Processes WACK */
  extern task process_wack();

endclass
/** @endcond */
//----------------------------------------------------------------------------

`protected
F./Y5WfdR(P]9=2bdPUZcQ-/]6]&/;Y0K&,SaTWM_9_S2[5OG&Mf))W^c-?KA^(Q
APX/[&QYa==]gGA&5A@be:#&e]\,?(Z>]C[GU3c_YT/JF>./CYaGa,d8C#X=YCD[
09,7PMEPK@cEOC0@M^IcAb)VWQB]+F[b]]3U\C=PL:J<&[I9;TD<[S;P?@/aT[=.
<aE<H0,3,<W3+/Ib-YT=8=:2>a_ZB=A3UJMDbZ)XIF24FX]H1U-5(2aF>dS,C[)C
bRfX&#5K3LC[&9d]M/6)M=A]gI_>gAM&UORWF-g4=XLAL.Y1NSB+.feUL,f+@>VM
->?1U4CL5NIRQKQ?&aHQ/Nb/<fc.-VV/O?ZN4M/Tg)MMDSR\)[-LfJ>0fUE>,&]-
4SP@I3.O,P]W>e0];a6P\3ZGQEXa5a;.:.B;PZVgd4S859#;L=d=,S/5>PL:=#bZ
?2#eB<F=_W7Z<bPI3SNe:7COKg(DOXQ^9_BTE(9[C@I8=;6SX?O1La?7F@YU>U(M
gOO-VMHKYMdgTU=f=Ye9=4:9-Y)E4cRK6.Z\0EEG<HQ,];5I+>aNI+>1QV1V9LX-
a4O@AQ_)A5#92>]?Q&dfeS];GAf=ZZBYFICW:,a#bVT)FdW+eZ(VH/SfcOaC5b6.
,e9=5SOPB@TeY?Z)5PCCV@1f2);?O4/:4a@WBZ6DE11#?04QXe/fNI)Re:D0X<Sf
)AJ[5+DSCG+D3CLQ#a9UCELWEYb4V[HG@):YcES_AHc39BaI:]WCd^XGK^LE:OZ9
,_C(9?AbZE;+HPHQ5VZ=5>bg\+1<&7:\@AH#VON?c?.B3J?B()4C1ZIL998d@G1W
YY_fd^9FDgf74U_C,>>H7]Y;@gg38J(?HO[N9[V#0,C0?4T8a(=d8?K=TZ0dD259
95D,/Ra@H\A=V025R[S-,IUD_FMYF6[E+]EB5/\6R<,^<F]EN7I0=>O+2#PLZ77P
,Pd(QW6=Uf7N[?XecIe<g#51U_+XQ38<GF=],c(;:7;])>X@Hg<cZ_bM&4GdE2S@
H\8F)LgJIT6VbZX]-dEL,.80A\f&HfQ[:b5&40(>)PGEG&-2cZ)[U038#<6I_K)_
U]0,)CD-O;]#@&5bF;+^fH;X_Q0GI?XaUB///f_.<^>cWg2BO-Cc&4IO=Y84YR/C
M&4IEc+,4LVGB_OQ1GQ7-Q8/eZ1MMKd=bbCcCTLZgf(b7Q2.-/A99O7\ReUS777)
HA:<-2Y,QL2X;S:RG7b1(@WL-Y;)cH&YMQ-97X&S=4W)NEEAgW@_[U@VE8GHe9UA
fcX7GXY9_O3C?JFC-=V<1B@KRGH>QQ^8YI]cZPeS,bF,g(-[&,7E0:@2Q,R1Y7YC
43?_RP84bNd02DcK<fCd7LRdeM55N81dQX@XFJ4N^.1RR/XC_:92W/X+VTH5N3>3
0fFO&HC2=SZT&#=c0:5,]eM7)F6(6#\0B\M<++\(<C6g[ONNd>5M@AJU\dZL/#WM
5aOEAa#493LDW](^LaCI9TIA?(P+dKJ6P\)c_Ug2.-&6+H&=(W-M2_ENB\=.MOf_
P@.UII.K7.<JX12=N?F2E^^QWVB&W<NSMACR,DZ@>0F1YM8S?X3,H-2N3eVGW[8_
e=VH:KW=d&BQ[B1,ag#;9L7Q:[O)bg8-R4#K[2TE2UL8+KTHSfCQbZM@@9dAWMW&
FMLReHCM-6(<SC0N]I4??EM7eZ3@]6Z8)FEY_7=EI\?\K?WY?L0T=TXW+4XYabd9
Z8RBGMP1E#-M>aEG:2KK@Q<;DKTg#69(^:DJ.273G5:RZJ\F\8d_05d7GTOIOSBA
c.)G(O>c&N9WS9Og#5cOCF_b4ceLR>+F<OR3d.?AUF1Nc-=/?b=.K#MT+]3V3X3C
/O,QeTU=-V[<;3c>&K57=R#IZb:DL8aCVI6KWa.0=KD8B6+OASO2&70WS@Be(ML[
31\g8=U;.2+49+(00B@M;WL711@efJ[>:M=&[I1NA&VS-(:WU4[Mf6aJJ[R2+Lc1
H8a6<F6X@^(?D=RGH3bP;<R3bQ3P]U_;W.9Y1G00X>Off4Ff:YfE<a&BF[e^KPG3
e^CD<]7@F]SVX8LLc(2[=SgTe^_5N@\:dJI7\dOF]AC2I4N5;I<^f9ZUFI#][ZE1
2/O2&2\:8a6J(CeeEJ1=8\NJ3(QQ7QW&dGA;&T352:2fM0>)7D2?7V_T(dXO_2Ab
:V:3Mc+4:DcUg2.D#[MBBI5bXJf;:E?,\A?CZ8H-I:QZX_#9@-_>+\QJLRf90JZ/
<Z0K=g.@g-;f7@O2W^6TaL+cS_T8-g++\8JMH^VUY@gMU&WW8J/-/_d88C[;(-VB
G@\G#TET8&JecA6LgH5X-@\ZA+KK1OXNA6e/Y&UC^8;aHT[/3IT>9NHbc[dAgIPG
,X(ZB.:U]\+d6Z<XGY[J7\cU^?2I&;00QbA\^bZ7U3U;d1#(7KB2@NLKX6K-H<<)
LZVV-A+D>+WOY9N(eZVdMZfZ&g]<e4d3Q\,I+[E.-5f&GGO5]Y;_cEc\VG@YI16X
AK7][G45JI8BOQQBf:FV5dC(N)W1;8^C&&<1GFPM0@gZe7\_;5AcKbT&@[J>a:1Z
>_A40[JYL-#6_Vd_L0P\XLE,)OFK0937UY?)P.SFXA+.P>;52IKc;aIe+,8G^4,I
gH:QL85d0U6ZH?M=MJ>0b(;0TUZRD)1RZA,67Z0)#Y@)Q2#HS6<K/\Z5FUF\).UI
b/AD<RCHH707fK5C@+E-Qf::8.3X;2T>f@^(D]:88IFJSWAU=670?2;Y(\+1\Z#C
W8W^M+LTb\&XGEK3f+#U&)]-d.G):X[P74UMF]F4CNS&MQC_(Yg7;WC^5+HWC\fJ
E,EQW6QAXI>.>LM@;^Z?LS=[M1NGf/ZUJ;Z-f>04ZY46-.)A^3DCAb<LI<SZ1M^R
10:=YF@[B52aMTg5JHN(^8\-GVaRAG(C\/C#F7OSC2&;1aC5[0F],e[O=SWOZO#J
^PB#);;fY]6TN]L)1:84UfaAaK\1.OR+KbFZY0U]()H_C3G1DVJ,P&V6HY7Z@05Q
.<]N.\c?-W/>YdMb;^6@1I^3[@QP3XT72)D#Z>8P&@S&_R69b/Ma+UV(bIU><PX;
:C(7B72&0JJC)P)5,L2.:F[NI&?)]#\S(G8SOTYU=9X=Ea#NGB:JH>Q2cJW?<Q[0
#0g-ba,-S77=]e>ZVaQ,Z^A,D8[Y4M\N5AJ)e4W6b1Y99@R8D14;<..AMQ.Y15:L
b]dMc78KgX&P#5gTgF=ZF0V1<KfDK2dgTYOfbP&&97^;)_8&RfOdcd)-]8O(^C7e
[N,9Pc_IEcT7;;bC5=V8AKR:?-WK682QLEV;)QZ;-gH7\,>L<c&3X3b;T#<.7g46
eE=TGA]I;][(\-X]]YH4_57aV2=d6A]OO#FE]X=9>+QDHB=aCWf@8D^Hc@;\^)C:
(HR3\B5_-,@T9)gN7E4D-2DbCC5\FS&N;65KYR0^SER7EddVfb7V-@-GRPRcFAYO
9c;(09A9U+5AC5Q4U(2feUE<0@&2_::caOX1H)eA4VV?AVR5(2M+;[f=6.J>EPVe
-BZ@KG.]S(WEZSD_.2R^F?)#FJ2bVR2\F7[#Hd,R/^)_&3?9U1Kb\:3:A@-5&YCL
1c=)HMFI<4USZd;XY;G#ZG143PHc[.E8OeeWEH)EU)FA+LHCR\8?;Y3gQ/N8U]^F
Ce/KV8B7cO&0DCbS/,d/PJ&O8U&<0LKFXf-BP#<KEa3ge#DTT(,cF6^gYYG?[</C
:0,ae.:g47Rc4&f_-_=7J=Y3:[J.d\@6/@40eHG/CN&=1)&0TG]V>.W+4a&.#d3^
Bb9(.DP2>2]b;a>e2J_.>>]VJ0c-16gbXfAbb3UI/H40T55=5RJg&A+\-^VHf5VG
e_c&/e,?):0OQW6V:E7&ACCZ=)e^6?W/Je&fV8XA=cF];M&01JD5(W4?Vc38eWQW
@85O>4Ud/cKe-U_eTE.E_SeG\C^96;=Y@5aU0T43@(5X64)f6-H5RXI8-H0@X\MV
E&S^5#g?X5d)B#_Ya0MK8UCYE4eH-\0K6;[3L@4,S]99ePd;CL2/Q:DGE^UIg\:Z
>A@K4.-Y#IQM+E)=UQ?S?:IaX?G_XHd++4U;(N8JI>.@]f&<aW9+KN_#&/HbSLfB
-ddD+U(<b?8e2WCd,YJS.aK:SR6IM_ZU\Gf8:7)J#SBF.5T3D6&/?Q/YBC]:&2eO
HGdO[f&U<U7^]I>6aCD.\86g@.f#a?5EgVG)XVTCREC/[e.D)Q72,SV6)&H>&LB<
7YKaL9-[aT=^6K.Y/<<V0<=2&bc,[Dca[GQNH):?8e-]3X_J]EIZ?LI(&a0YAA,J
RVPG,G=&B.9a^0J]\GB=^BO6AZRWRQSV.S79#)DI))5<&6GXGfc7HGA<O2+a)JW>
@8DAJOE72&Rb/]KJO0M-d=be&1\^>Yf?<@P3\X_--QQ?cS5.ATe9>YXQZ/@,KJSI
Y^?O^C#)/R-^YRK)<-VVa<Z<W,Bd^R3UHI3QP@R6g?Dc+HReeSH8:AA,.NWN/J^[
gE3\#H4RFYN.KF8f=[)>;G/OKT)6UPAc:B.V^0]9.:cB7Vf[S3,7;H#F[##).[bO
RIBd@/^3;HY=((2X2L(@P:RX_--5RP;@#;f2,9>8LW3Q]M7=LMd[:]ODY,b2J0;P
733GV,=XYN]dTC+3@d/fT#4CMIAHZ<DI<caaV)(]#;C1MI[98b?PQ);)DU20(Ra8
4W[eMeF^XX5R\@BWA13-9O.S[C-L+Y:VI.[^]?c3X;.?EE0C&f^1>:JO;=+900HM
U?)+Hd^[/aO[cJB#94?_TBg5<F03Y+@\3BR)Q2O=0bYN6&8[b)I^;-TLdbHXUN2Y
5)7_BI]DJaDPZ609#3-G/RC><30FHJF[B.X100BbR19IS2#7M#X&LGe3W1+=WB9;
WJBZ=@#X7NE6E6/KMc-G+8\b)A7-]1\d;:;J/f86;..;;#\0#^0gH2-<M<<9B63C
.6O(aISbFNeX^NLfEK(7e()RA=H&<)].>CON/b2g45O]a_VQLU#6P]?F21egPQN=
C@/O@H^a&G9_)LSY\.P4]R[O@?Qd-+N-0/gX/b(#YLcQEF7#RFN1J[+S<>^_9<C]
1fU_+TfDPRN6.Y3e9E.eH1TV5EQ-B<E<,Y07O7dT5bM=3VEQ2Q7KY[H@8cEOS4R8
Tf-J<^0)G]W=5^)G&4c+,5DH58+AVBH7+N/2.=A)HRBdX&SI/eFE)>H@M$
`endprotected



// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
`protected
gS,JRb@)=/\:4Z6)&>G8gH_5@74PUc>>1ZCTK<:TdeR(5,-AT<=5/(.2]bDQ13dI
7<=9;K5F(.c;O9=cT(U#J3Yd55,D,@YDXQ_X;3I9=RJ>MZ2fb6+Z^FEG:;AG0Z^0
574.UX5]#H51CP5_c943c54WK3TH[U>_]-<2GZ.VT-8RT1E_Q=D7b3_K;HaK<3M(
cN5#fa,_VA/.,CDd-PP1KJ)FJH_\76@FdFL[@D\0e@?H3DQ9Xd@fe&NVNbIYR&QQ
[/4RL2QebM)(Q>0#a\WDQ_FGgC9:M-G]Z^6?ZT9bGa&3cU;6CN&fSQNI<7T:4#@6
GId[FgD(]4U+X\4J^>b3RP1O.05I;:OTFPXG+)d:;.WW2.e3QC67^N423C#a,>4E
P3TB=eFX3F=.-8[4F8;]JaN#(&c^f=4V@)/(e9P\(?Q<CE[V):b47;\X?(ST^],3
CCQ:@:aB&FOW7bRG2<RA3FX4]1@==W8N(Y<I;EX8QEQ?TZKK@8(M7XJW36+f39N(
fOH6GQd0</9]g?b[G1[)L[_9WZDR+d;RU>ZU8#a&\H?c+bP#BD0:6&9CDNN0MOce
GCWg7#V61Oe)P6EYH##D=PP;^?1dCX-E8ZO3Dc=<J3O]bR;SAN:=#.WQDgdTS+2#
c-H1,JN#0GOS<>@C;:d>BbS1>JQ]^7dIg:9]dbW6=FPDc:1MaC3EGUK]AMX2U7:.
eD>I&L+^=V)e_g0O)JaNRX(O5dJ/0R9#aba>376IJZB\,BWdeNTUM=J]FX/Y(Cb8
5=XdPGAVWN<4+29ObQW]Md8QI2f[-K)dNd]Ta5XG\8GIHbSTTTN<@_J6e_5=_[-Q
LA#_HQL9N4GM,3g3Kg&AV(Bfg3(N[b\Z:4HPY,_Dd0_A@<?YOcVd3,<BHW3KW600
^F^#CB-KF,WT@fWKYVeP=GQe^G+&]_W>ZT_8LDLPMFR@I+HcOWNW^de;7_R/(@+2
I:5XSJFX\)DS?f2RQ2cc^G+1^_WM]:Y-9@HHL5\;?B#[/gR]cFAd0I).V,0B:9Bd
1;HFYCI?3W.B18O?(TDG538Z\e_@F/).JAZA,=-5#VEHQ[?@+]EXeOIQP@2U50H>
8-e?eQZN>2+K?40g^6&-Z#.Zd:0#SH1I[.MA\SW^RH=CATc_4ga<@MSQK>RQHNN@
K#RN9\&6<TQ87Efc@L9F01>^\]FS\=gWFO0b2_UfN:^A,B90#D#9S]3W?4\\T),<
HX@F-7B?d8B3>aV=b#f4[E:fE\/FH:?(@EXV4NVg[6P?+=D<CX,4VN-cW2[2<:+F
)5P82a3]XF>P]\C^G[EKX>Xd3UP?I<,5UbNMI#:DdSfT+?WQ9>^Q9O,(,L]),]L4
OdQTX8/V+f<UDFC:E8^)V#-fB:H)KF7HR8bYRGSIK&Nd@&P\T]AJ;+#GVTS9GcEE
[(F2^M>EDJII\aC+=3R:f.a#3Nf_EZfZ[)FY?^L<)HU;6+[/6#3+g.PQV\d-=e#Q
<.5Ye;^>;OgXdOW=>MT1b8D@>C5(?/@a/b?LYN:<EZT^#U5E_aORZCJa;I]XQ5MZ
V#&cVYZ^U^c^6#5)U0[VG;\+Z<:Y2B2a1K[#_e2Q,X[OFO?Z\LHQEXI2+g7?b^:#
R:=D(BR=Y6[QJN8_K:[gRg@R4GK>QGM0NV\/_(RSWJK]_<;=cW>I,fIUAV?@(X=O
?ba[,GMc&ORI47VbY8AF)).+.fYK81ED>-J5.(P,APba2N<T&V@#1EFA>.e<],]@
eN;Oba85SGJ>X_,ZYM+0X_g@9_8g+&>3BLV4UZ?O5/V8M7]&)0I8O_A?Gf_&OK+8
[WVR>JH0B17#V=R_FcfPFB:gBS=g6T@>cS^Jd3&#bI+9SJOa>]SabDJdI&25AH6a
5GJTYZ&D.V(9EYgRc&@H&ZJ0.H8XZ,WUFCD.IB]V<L#-DCDbO>;AES^(W9@Q<fI/
&7&\[K0K]_S<AJea+7NGRAJb3=0PK,W4TAcK3.56eLG:E?;f@/QSc6)+YM_[cU2H
dQX:^KK=B>edY19MH5Jg^G=<J.cdMCf8ZT5YP=]KPS\AaT+/cJH_:>ZQDb;dgK,A
GK&1c_eE,Y:@U-4E\c_Q^+NZWZPa)K0[?-V<BE8eG_4agF6]&?cR(CQ@)##2eYg#
YbD2?0<HPJGa[G0YZ[;7/8f@Jc7,dOSVO-;^2fcU>W;110DB7L[L[1L??ae>^/;C
82RZ)S^X&Tff9,&<WA>534,++E/Q@7KFD(&IMG@,<9Y4D3Bb?M:6CQ^6#e=8I-@9
6HH7EH-<.\Hf<=B^LRT6BB4(Q4=M/<CXR:7[^@B<\Q-eNP--0J@c6BD0;I2&@\N:
9_bN(2f_(<OFL-g]E]J:aWccL]?5EOT#XQQ5aJ1#^-a3Taf28NPW8P^IbC71\)ON
;GW5&[=BYQ17GG.\.eCE8+FB,ET=cS#5VL-NBF3:Q8=aF7=VA.R?@=<?O._gA84J
X:J@N&D\5>WJ_,LP/DWOS4.>@^^J)W>C);WB?d+KIGSe<:JBOgOT<\MG,?d^^Y(C
?;I0Rf;VSY_d\F]4EeY<19a\:,9MJ]Ed</CQfdJ2Y_Baf9b,>Ig=-Y,96\/+\6gf
1XI;,^64C(9XGJGa;G:_-1Ta\VS:4cC-?cIR?@5\6]=^N)&W9b4L0(Ne:5Q.a4TQ
Q2@J\X(dCK&Cfe<[8=H3c+;:95A&NQ#7A4?HP1+b_W#S(5R#=_bOVBF(QPPE;dFO
@+#_HI[+MYYV5.?,7YA8226f6Y<AIFb/b@&Z8<EAYfUYEg<HG&81]9/40c>Q^+;(
G?AI?0&.3\]]KG<]_:gC,F6LRF?UbQ,,UX^TT.]=2)7EM-b,#ddJF_Z4(W:<F,;O
7UAA7TRU+H6/V65Pc@d18bc>e^)XZC?>Rb8c=X?^ee)aa(UbgJ4]YAd5Y8J]&BZ+
6Z4]ad_(g5D3:3U5-L#fG,g+_D;0I,I&50O+7N>TNIf_)R;?+PT/-Z3:JDaTI?C(
3[CMV>V&=g=65VQR;]X6772S@NC6)gbPXR[3S9Yb[.IbWgPI&QP[F^CXeL^JP,MP
NS&d#+Ua#Y-PMX-eG+_d(+C.>#&4]bdL]))@+.R]Qd8+GK#=2F5bH><Xb<W?/DP@
/4b4&[EB1=SBFQI9G_0O?0/;N63dV#dZB@2Q5fJC3(46CAB]22.J;TdQJUP\&\He
bcZd8>&(S8)IVYeLVdRJDe2^6L<c?I^F?9YGH((aBEgF89J(E:(A6-MLNBSRE5S3
_<F=d^XIJ_1^_e6V/:5L0f1gZ]eL=VAQQ?Y;(Q)_&+[2^d4b5\bV=KWG<^V_<ZN#
YP[Y>H(aLVQYP7?I5KM6PX:7<=:e)dYAK(cM,4JESgP]baR+BXCOIOHMG=E/^@0&
F:fZV,S4&M=G,U+XI/Mde@>.6T7a^1S]\W#1(#(](=17.5g>ge)Q41a4FI(FB.P#
B-aOg\V_Sb#,Z+K?YMHX(^0fVUH/#FY+MXGF6L[MI4)a=X+Ua85W:d]I(@R<Y6C=
8A/YDM:+O6B)Q:D>8KCF5U@.GQ^M)3^Ea>[UHUR(VE:Nb;<..:.X6EN9Cg3X?PFf
NXAfe6_1YPc;0b4@&e;T?[NccgHY2T.:<TdT:;bEWAc^AeMWWa9HFb\G._e#dNAS
P\VOQ??2-5=6P[@@LR3HfZ8d3)a_ER7^?8QD3N7?>MZ#W@=82Wca:gAV/C,D#7,f
Q+bG&8@Y9>cU971,\(;aD3]&ef;/0#.RRYK)e?NXTFKOcdU/fgE0U-.VQR#YPO]@
5<W76C^2-Q082GUNX(L3]5Y-,#b6V4@^>[_:d.W_7e94P/dY<Y5Sc_5=H(7eIJ,.
HGZ04[T[/,;5UA4OaaH\PS1a&e&BV\Y8JO\_Ab0VQ[?>UCFgZAN<FB:T-1:YK,YP
C8aLHI91MFEM(B9V<&H;>EfY]N;gLI1].dPb&:f>AJUYe;LLQTO]E<EQ\9;>:KZ?
7ef(,G,7e2B&4D8,6<AQI(+>\fX.4[g=VW7T9E#+UU_=4^EB(I37KB76827<@c#^
X794g,eEF-g\f4\\T0(7&R>UI_d>:e548H2->_[e--9HW44I(NA9\DXfTZ2(C6DM
X__0&VD(]&#^D&R1A)@G\Fdb4BKeG2YQQ3ABA1VR050_cLP]<U<OCB)V1=)S)/>e
?\?4PgT3;A,G#&bNg=WO^&cB6KVH\^_];g]_?)5^U?2RWM&O0#N[5b8A@d7>]FR-
V<]8R8TI]-(8P0>HQCe6:;&Rg:+U_:eJO\#5MNV8=@Q]=)>3+N^&]=;?:Y9dUfbY
-BZ084+_g8.,4gCJ/b0?gL&E8JX)I&JbXBC3W?dB=P>A1Da67QN0GCZY42)f4Xg3
F6-J?;C:^7+Hd31;RHDR0e4dT;1(J<&W?Cc?Z3M.2VK6U]IKT7ZcHOLM:.[>-E_F
@9F-=PN?NSXHf(P-(S<?5HKAL4gT33fEQ8:M8S@K;3+c/3.[R]K(.XIT@S?ReXB/
KSfX&;>(F4PQM2Y<XWe]F5gg41B1]PTIMX:VD5g&HH?f<G,0-(c1O]0/F_1c(e_/
bfX9FO6QC#QF11aHb[VPZ=TH3LaRBgJMM.SYAaW^=FGN57_Q7F[PFW,.MPE,e=AZ
(:1a:FHH2544H+fPS84MG(b@T&Y[_I#T>cHE/D_+Jde,aOg;QEP6&T(;S(M@OVK5
LQSS@+5I(B)T6KfO/JF(5V0?B]>_F93O]:&5\/\c@I/+/42Da/S?:.26C[?VPKX,
)/>bUTT0a+13+D0JKUJ/aVM7IXAI4N5X[ARXP5TZA\+DfeAO&UU4D48R[B](Pg(=
S3322#:6a[5QU-R7OeXHV2Z-?(3SZOT3ML-@;N#]PIJ7+\T/f2GgM/HR5NJ))^PW
-0J9FF0YB-Pc3@>21UB-d&X#+[S=0E@^0-gM_E0-aLIGEGF_)-GNG[eK:BBZJ[,\
6/[?PARG,D]MD#LT]N^=Zc[AT-P49Q8JdX[aT;5R/8G-&7@X91H:_5dA)H?IFa:-
8MI/^5)ZbK1D(Z.N^<P1aX6F_;ZU-URO+EJ#Ob>#[[V^4H:Te;:E?8>bJd1Y49?>
_PDaWK1<g6I)7dedf1Y).@L7>;,&>7(>aQF2+fY<_5O-7?EaO:L@JM?W84YMNWR]
BS+d;S>KFbgZ)R>^a0Ya2\e\_bc3YfDT46<A_g10NeGbP<X.\>DUMS>?WYB#A<RN
D]3K7CJ.HLDa&_5bY&:KO+?S4XUVf1_#:BYB)?BeeA3#@Mb>327(6VF-/-A/4a=S
,M=#5NTG;P(534^2dXG2INe/9J111TW3XNQ<F1BPWg34\8]K:^fAAcFE2Xb^#>IJ
fM7P@IQQXa/UM5E[[CARJ@a9BTF\ATI,MX,6^8.NLVCJA<)];a<)LAg+]<:MEPZ[
5E5FW(75dG8J@5_))A5:/WF+8,O8+4:M<DQWIM[I7=GDB-?H)4a#&/1,>76T(JLK
MA?D2CJL.VJfcRb7.#.NXQ/Z(O(]dX\bQ<8]COG1;4JAC=&NKG4:_6GgCA+T]([8
d#>F=L+JQ>.1\YSLJI^V:]N#X44=F&NJ?P&Y&@W[97:(H0GI99OPT@0/D@@Q=-=(
1T847QC6[OQcLVQ1X<V)R]TR-9(L=QAX;@JB<O(_EMW\V71b;b0\(5&WO9A-eae1
_/J)aGS./0RfdL/b_eAbV=3A>A\^3YMXA)J/WR,\JVGL?ZScNJgRTD07[\B;5g>F
]6U;gcgEP&TBN-.4+QGbKRQ8V8d)5I/;:.\a8A_C^PIbFJU[6Z15,?5DF4V^U>(.
AaV68L\2+(+.)K16WVD5:FHGJa;SaB1M:S-GgPA\+\R==&Pcd_1^JH&E>0fb.4+,
[.7T#04Bb?7N18X31Lf;d@-WH1a5S]FL>DQ+T\feGd?e;N(PDWf\-JKBD2KP85/D
(IHgcg2=2JQab1A>D:&]X>)J\/1=LZNRT)3[6]3Q(T^<<[d\G\[4.?2,fZaJe0WP
+54O5;f]W@BH?\Sc.CZZ9dbX>;[2#N4&dKEG3T5A-^^f1)R7387WHR#\](8KAPG]
\HWH>T6bFd=HQZO8JPZQeCcLdJDH?2Gc0GUE_&7])dc)d^\=/W\FU0MH;]8aN/aM
a5a@^BGP[/Z>QGY?aFe+fJZIA974gP]+;E_c..4e:-1Vc/8)T:_M9DG]T.U<fGY@
NZ5VeOJ40D1T&0-/][[8@b11\+T[^UQDbPSX;(1Df9>S,ZT(>UK;97N1V7<..EZb
a,G\9d^626O/O4M4GI9-J4LV99D6>_6+-80;R?Z0UO5)g=B.4EVCTA9P0/81(.&(
d5-SM)P,>XOJYOR(cFKO?^bJ_d(2=[@)#823?)OHDfa@FRY[:9PT)TXPc@8D9F1/
RA:+W3_IPD+-;C\U5WL5,Q4E,f7V<-G,>#Za+S8PC,FP1RTeYB[#G(7]cRR]14QH
^(a5\->LbCATI6P>V\+UbRaU[CR&,PI(b?J,)bHfbR>,:^\.(dR.TG;A3-#QgOJQ
d?)(B:.HAFZ^5X>[U#+:edM.6TKA;cMR5.7K4C;]UEdd68VGdF>O\Q/e>LYYSQ_>
_V#9((bLg1._,R.<S_M01>Q-aWaF/C2/+=F1J727LH_aWTdTXJ8PR45eJH(;3J[c
bb\IRB9&#e<[E_f1B)[G0&DVX@ZRJc?W<0/F&+7IWB_fP4g^fP9_GO-I&c0_@g?C
#1NK]NNca+P9-<M)ZPW]3Z[:G[4HC<B..=PQO95&S@?V@7=B>a2KMa_dZeWU<>)A
?6S:=a,-Bg/)[0A):KBU6J;JDLaHVB>2fCbZ#:L\Ed4F.(QKg9b>YWFfW/KXPPW1
cU_gSYH/aM?+ZH4K,-L0&_Y3KO^0^F]JOAaC(I?[RS..PIS(]UYXIS7-<c:Gc+X]
eNCSU4d9>F3)L_,O=DBK2=>;Z_fYeBG:0@a;eAUD[\(,]:[:CXPU9@=#@2XLCb-+
-EG,cW7cT5=41Og9A26)+027eD@6JT.D_;6-R:,<6^dN>QV7TDSB[7<H5-&@WTc+
KY2@(4/CJ_#FBgT;.(-MNc+Y,2&H9WO>b0bF+L8W[<P:R@N8C9ETB;1H9B#Tg,7-
4FLf27Obf2;9WX,6:A=95a1]>?)F45+_BMY[(:<Q@R5&15UD],dY@L-CNJ/2X#OJ
M_EMcW](O;J=b9d3e2N?,4:N,PL)5J8FLL(3(1-N@ZVc^Vfc5fT_LCYZgM1g-6P5
2(TEF58M(MGB0HF^fX:#DJfNY?BcPG/WTb^:C5[-&8:-7e1Of<f3L(fSK_JN;[a<
QV1Z9gC)Q+=Mb\IQcF2PS<;Ne)<EFGSQ?_[LWa7e_DRJ_]+=WUVSV40BN4/NCeW<
9P\G9J?N#=XCU3=,dZYA;Z5fSc])J.[f8;cW&<dNJDVSJcB#eK7<[&SLC]7Ic3-E
162AL8eX@Gd@.HI\U_<B_EHLc9LB<JNd(Nd:5Y\2e?W+7G)/?:ZIM<BHQ(V6dWXI
V9ARGG@c;JSCRA.+d&@YDNXYEA:OFe[4a^LU-Gc7Zg8^]@-&\Fc_2-=6]GSU+dD0
IUHA.6(cPK8JMS)RDMZKRL9.bEe:,eEP9LfRT:P^IH]N4dYFcW#/DE\M;c;54:Y2
[I\3A1+2SYV[8F9NMDg:NAHF6KQL(,Ib1.VDT(+F_9:V<;T6S^#N-Y]A1=C0K<J^
4>=;)A2L#0OUTWGB?4FSN<V5F[6SdD6=SMD)/YJO.?<<]2D;6.S#Ed3YN^dKDC^Y
)A)D17U[[:=Z8^,G&F,?dZI>O32g/M=\Ma=?I.YRNIA\XK,]#XfD3(>CW];J3\O>
Tf\3_NT@H(YK#Xa1KTR3&LaeOK]_>gfD;1RZ+.NV<+E<Qa)fa@F&B)7&b/QH#WCU
QDgZ,W1KeBMVW?F&&HKZ4-O3YP=Jb608)fd_ZHFXI7F1RN<Z_#-(=7GBOT/e7I?N
DZTZ6.Z[[\gV9c6aQQV+Q6cT_?]QaF9&JDF4O=]I5NB)fE55#5Vd=0_#2JHeJ]e/
<X4N&[ZF,5RF?NU@]>WW>5817RdO68Lc7L>NJec_f(&5SE#\8Z\+E6Hf6?,LS+b?
)^<,#5HW&=35eBX,29>9QQB)>U8W8<d;T947W7=_;]YJFDS:[QRAM?<RK,bICVIE
&\/4b=\ED::+/)_6+A&VYFU68N2WAQ++8Q,fQf:U;fPH_fJG02bfRVR53<EJ^F)8
L9/1[J^Oc#4;0&TTR=4^A>;_#(UEQC[?4:6S(U5G4<EJFa+CYOS?:^eCT(IS-X<K
LU(<XA3#NWCPQ=c[7aX^P3.&_;]d=:>L&&Z^?L,9@P7Td242?F0TRU_FM73-3O3Y
Z,S0_B/JR^E3-M0gJTU^bJG9U+R1Lb[Z,>=?c,1GJ725<&X&^#4NgX_ZS3QE[[VA
/-:bT;YD0/^I#9X\0:5\F:L8Z.U]3A6>_EVa#:5,\3T3;85XR)aGJ&@-S_a/ffMC
-5HUTT5cJ^4JX7Fcf)X2_T-O.\F<?.).;8]e?3#AFPQ6.5/XSKAcHYSI#_=8C=Zf
V[9=A9CCA@+_O>80;FS&TJET\J1.9Ddf/)[fNb1+.YQRF8@8TP4D_&5aMQ+T,f2?
WXJFNX8H/6UAOR&E41_IS0X273K_<(1#0??D\]?M9b8(fC/;ecCf[Z_\>e8C9dQ[
5WQ8QMQ:>M\AO(_4^\Q@)1C\f9F5_CcNTa+YO./WHEG+@+5eTA2H(@.18TFGZg0?
.UG^c\R)PS-8P\WMFF9VXOGL9(A9b#^\3\e8NX7c:FG2I/N2GR=_cLEZKR\=_eL[
?,CGSR+KJ/VLc#1#b#+5T))Y:_Q?.#RZgcg2-X[J+<:64cg5[&[\?KaMIa-Ga_LO
e\b#X8[3CG)^GRgTVa07^]]SI-^d/H-64WZbOcEAP2^S78&ANcf4I/2SGc4A/e]G
Y1+(#\UYIRE]dgC4.6g/EL-PB,-SdR06<X>bG0;3/)a=e.STT&[b.S+JK\36O(d,
2;Mf,(;Kd?WV6CJ[+J-C,;52IY3-HUM9/b,6gDWORB5W>XY-0Of[O_1;KQJ/+RSg
E4SdVOdaCdMGT,eXCR3([;R3fb,;4Ab^EXc4E=A#8D/HMH]D(1:5Wac5W]>Hdd1e
GB.TaD,g7B9S>YCXM(W6CQE0W@1TZ-++/g)F(1G&@dJF=W9DZQAGc&COT7\PM5E_
K]R(?&fUECP6F]KOfTIQYN3I)eaCfN,I,0a]_P</OWS?B5?[&NJ&^AE[7VGTP:JX
L76d+2XX7AU<.R)bY=?4S>=B9Sc>SNWZ(8DZ?MFgD^)d4PMMM,I]L@0;T1WPBdeY
624NYCQ;=34??T^JAKL/XVUO9H/#8J)8]3-Le4b6JgLebL+d@P6PSGUE=4]aRR^>
YWX1bEXYAFf).;eV68D.EO\_K=:P_.LIgP8>VW/:KCT>bfB)A)KL_GAGSa9>Va<_
D_1b:?HW@O(A.g]b([U2Nb3DB5F95Aa]\#>a[K,b;GBOF=0N6W[R=JGWSCI_]WKc
2Zg)5I2gK?B;.e;1FZaPb[eY_LbaUX_^O(N?IF+UE6IJO=I;Y\?ST;^FZ\Y@a)4P
A\]2Q#MgGZTH.a^O\\aUg8CT3(VdW19C;f)d@C_&HG#A7L5=eU;6Mecg;WX&)9[C
[F0?f;=8<D8EUI4cC9FGXaegW/eIP;Z75GUVW(I6,KC30DGfL8G_23HaOZ/[SN&(
>@3D&-0ZNG;a0\a?e.23B1BNL]EfW-Id)AX;gD>I01&A#C7SR6g>^,1XKb1@]b32
BX(Je75B-,XJgSQL^LT3&#@0]a\(/BV.H4M_WgFceVY@[2^P(<E]=+476;H]Ye4H
(HIaWc\g>;U@;Ld.c5U9a^<N,+RY:8BHR,J6XAKE?._JHND:@H2,(;.;SNV@=Q:#
VcQ^-W0gRK#T+g._OC[(N(?MG?UL.\C>GX0,B]KPE;\5Df\WMg?Zeg;&N@J;X#V>
cCB1BR].a<F@+YH[8gfB.6Q??AU=FH#cW##<]B),6D<DE#&0+_a)@X4#BIc7-#PN
O/F@e-_@Ic==65Y?9GR/Q;6+@5>(bb[(=6.S4_[EI<X#EfIT[\dZI)9AT\K)FMIQ
C4bB-]YRdGDJ(MI1UG@_M_PF>eD5=.]CFXJ#3=(0Z@8WID#KK^IGb;,QC&/D;QJ3
G6,_=SP]Of#WC:E_1J84=OJEKT5?2_M[Q\(6-2#Y9H^DRbTO7#^VUdHP0?IA]e]E
_fQUR3]/UQD]\(g#;/,bP]0Y2==7(^4De^IG0XFccb,gbdDK9,EJee(9-B<fX&R<
/Y9:;9><O09Gc9Tb.FCZ0gcZOR0Z@T,^3&EZ=^/(2E]R8KfSR;;YL\#aN9JfV)]0
0B><BZfZ2V;\<cC5+(5NWVa]]&7L-DaK\aAHS:I63D+K-C\C(V#-KZP&0BJcgE]+
-dgLg+S^W3#[g8Y@@P5YF396==cdM@FG@fT@+b]Z&f.K4fbVUQP^0Bg0P-WT>T/.
,PfF1gc_6OT3LK@EfT/49[#=TK5RdHeVSe7Z87c7f#V#g9Zg0Zf6+c&+VC2NYJF8
HeEKJ9;N88D9E_KBRU1+&>5c.AUBD]C&K_8aS#SPP-Y<@9_RK(V9#AXMO7f\G&XN
((S_.U<?IX#?G\M51I52)X@XG8[1WGF[P?;CW7HG(ZfYOK^=//KB.JE-DO_SM2-&
&a6EA76/Ie-]X:?d??<9,GbHT?9g?L#be6@#8UR1^Y=2/6dYOWb@a6HNK<ag=Y2-
cAL@N_5P#]]9YO/fIB(^=-O,3dVH82/NQ<#O;bDZN42c+VE]]&HF66J(gPP.O3Tc
TZ+cA6(6WAC+3-9IVEK,SJS_0Q2bWV(;Rda0=1.]ddQ]f\WTP851,<c4)3)+7\A>
g8)F9GL(\,,@I_fXg?<T]1ZK^U?)>C<cW+?<YC21=3P3L_RD0+E,C\Y.HIFg@0[?
OQ?<.ca2S8H3Hc41P54:O&[PAJ2&F?[]>Z-S[[Y]-)/I06HCO#8D8YJ/X0]H5P)g
4F2b#D#9&9\5F(c?ggH<<F++G:\252P+R@4GBbIZ<SR+dJFYX3XY(O<P(GRITA8^
Id/7I_MKKVcg_U-ZNc6,O2M\/)<Y?:a;D)-5:-1G+E31#_;(d:52A@c]GLO1LDP>
PO=M9,MX()E:4XPb=NZ+Kb_TX8NH>LRI&:gZGGEO]@)OaZZWdA\;[f900.U3L]^>
<5JND45HQZb8bgU)#RO=5EP[W>:L>?HV1B+GS+\D<cA7BSf+e+Cc\X8ET(f,YB@D
;<Pgf+ZOZYI92/BR[CB0:f,TM1@8C2fNDBD.B67ReC[3>WWcN^e>,9,&I@abg;3,
DE_N,>#SUDGH,<D-/#9Z],ZO)2\<e;VdLNO18T/g6VAad9[SHW8F2WcI<L:efS;6
SQNQK_KJ4B@&2HBW5e[.^[^MH?=58MO].ITKS=5TIE[/I\]VBIfVBW-2PU@ZI6Xe
P3JLQYY:=5MBfb:=dS50=18>YcBZD<B21\^CWA3T2)M;LX?d2ML0>afdb;Ff>BXa
?GH9L_/1D6<N3e^BdD@bLcf:Oe&.4/9Y5W4N0g\@1PK7SbFN&b-M_D6KFRNBM3QF
9@a+Y7-9PG80/USCQBX-U)R/Y7ZG<8.4ZL6GD72\=SQA-Y9O-RD:_J]:=_]@gTH)
DKSgDfaQU.@NK@,d8GTO:QDf8c(+),NEfSNKfGc0URZ[.Jc&[e#[B<-ZA@Ud(1&C
eZ-LX)bTJ#NR<Cg#)0RSaLe<^dB[F?.b)(J^d6L6>C\&<>QC/g1H.E32^?7B_LK\
:Q+]+7O3.;=>YaOVK=c+9.H=d3a?dMecE;eI6^87dbJYI\OgWL2Wb^TaVdK9LQ-6
FH9)5XbM_^eY.X1)B.=;^V\U(_R,YdLV97S<9NdCgEXHQ,IN9Z+XXVb2[:6Q<EL;
574S4#b#6e@JK&^[>0LQV#9,d#gdGEPUJ-=VDH]MONc.0MG0?7YE8N-ff@>.?W&X
2NXQ0;CLg>N(7g0=&4S.[H>MS<UaS7,I<T]N[.?LC343H-HIS:)]9;Q26GH-(=B_
M9<>-,;Eb]M78Z9Lg;f[+H]DCaZPEI?7:&75)-+]_SXa4VTH9YRVHG][BK[0A6&2
G(JO=Fc/&#Rb4dYUZJ6M5(MAe]YOG^bdTGZJ@NT.F7ee,O3M<49Lfg1(2@a:G7g]
?X/F9C4]/8W>4e8CD-ZSc(Dg1ICf(/9UKR[\BHb,b.J]@6de2E3/dG?X.9Eb^K3T
?S]3>7;+P(MECF,WfAK>dO^Z<BCPEabFGcG@Z,,PER>Q#1TB=Q=(FJL(d,PBKgKe
\,c)B/NH.fdeNNW+O-Pg&U7^#&SW)MUc301A8EL#.,PHe_#dc&DHNe;B;/g8b-=f
+Cd/\A?cL.J](ZbM5LII;.AW>(@H-;K-]9bDPB)32#eLMK8-Y^A^a\2;L?(VU++;
W&<b(3Oe9=e6E=1PDDUBB3_c?CP,GEMC9QaFLSWJ,-.ET=^b:g.=]OG;OOCJFeXD
YY,9I34E?7cQ^VcMSSRfFd:[+EX_5bA0=UZPY:B^N_\QNM<H6bF;:Xa#R8Z60BEG
+O)/YNcEe^cFdHRLdePHKE=NT#^CB5#J^I7[,<)0ZQ#&9b\M^-Q:e:GX4KT@60CY
cB#W8Q\IUXJ(:cAO2Kf_ET#_C)KU[6\R[]1;A&U5^E+QMY3OZP\AZ/[^ZEF2]2Ba
L40d<VMZ5GG#]0@REGV#J6IZO.866S^J7FecLd1[<R(a\,g.a>QF-<U>Wbb-WMD(
UK==6T@68[OIV6K2:=((:0aQ4+Q:Y;&5eKYJB=[U>fEILX=8I&f^)-=+>#.:C1NZ
R#db#>b_V<,&G(eI\@VJ^8PeU_2B=IcA8(dMLJN27gFGFU>?JY:3R&ZKYO3-3=6I
Z=-/<L4PH0>[\#AJE_I>(;-b1^[fY8KZ:E&8)F;&dFaIZ,G>Jg<+.>c),^eGJN/F
4N:<QT^>@aebSG+?O>fTSKdX<)aR4H=T-Ke-SL6c85F,3f,39KNGSc]M&,VTd:4g
1gLBN[:fWIIWLdQ[S]D#FG;eWPP(7_?_&G=G;W2e,G?\HIC(\T+E=e4IBBTCPePe
H1aTBY\VHOa1c.;)H_6KBS7(GOXb>+&:5QcI[2Sd3)QA\V=Lg52OMFa/]a9Q)AX2
aW79]KAH;3[P^QB,+9?F>K4Z8U:PG1@4]KZ/5@CD9/Q:M)^]8L?b0-d-VRV?>ZS]
U.GKN-a[QG-<K<CTE)NXKWF(TK(=FZY(DRf(F=/JT_.fH\b[XceS+)b(.Aa42fHU
J7dCfF/Ra2-@a5fE:L0[XLf(>,Nb-@\/(7d.WcV)5&cFQW>R_#-T:R2O3,Q(XD,L
0AQ@&4TO.^O/3Bd]MZ=/5;>^DS+Z_+:(>QU<DN#F,,TM?c#aL.=V6L&B=Gad-OKW
[&[+W2cb1^Ug(PDP5>X#acdT>B0201\WH__GHg\Cb>6_196b&TOfHT?7/cc3=R6:
/G(e7JBg:fc5S:2:^V=]U?=Qgc_YL<eCSabO3=<P[XE/&4)3/P(cSI:=_;C.7bW^
SbN^fNN3)fD.1B[:PgEP?LE09#4A0O[.I<TSb6QX=W.JD8<9-_S+SK<3IDgS[\\#
O@_d95\bCPWFI0-NV9U0\(IKO&,L/g8:\AT/.X;T:F0e6Z?ADL3YL(MEVU4]Z?:/
=;#J,RM0K3(XP;.,@[CgSCWX5.XQX=>0,dX7PQ)>;[687cX/TCdCc_D7]E_a\&QR
\-gbV3(<636MMDEJU:6A4\4f/X__K.FCU/ILI#TJR[4V34dDI#,ZgV?gCbMP5Je2
?U>]?EU1V@,/)-N&-YJRf/U3N\5b_Y:EV2D74T:)ARaX?R&5Y8c6,\LU/]KB,GRD
OYHX1V5MgG(J_+Ec9\<O@C8S\JLSUaWCK,=9[)dY@0L^W5e?e2Tf;4.Q\\V/=M]^
#2)NU]I5KO3G[9(-ag+7?-C^/Q(]E,2c,]?LQFZNd@Pa.XgO0+HSOEcU<9FQd)_S
Agf1-O6PFMEI_gNH+=.c(7(E)&&4]SEZT,c.be1J7ZYTY@1XZJ])J_-56/Ag:D/3
LZ2TIJZ<Uf5@&/.d5D3G\]9V_/;J\=_Y)LZI=6^LDA)G2b2a#c>4JG/LFUD>d(,.
1&3SLe+&\0KDVTNa36Y07-6[PR<\>L54N-W07.V>LZ6][))ROXRVAH^(.KbK8A25
:F<V3EB4))2/HD.ZHP,fD7C6fXRREGQ,:<Q4Ve8Mf44,DU090>QWYG3U\e^>6>.9
8W^R-0?G(,KV=Y\-Q=@4E47NP+SH^H>B2ECO,I=4^Kg/2-BdG2X&0DfGA9d/<a3J
^S2.?D;RX#QK9-[BGXXAB:3L46UEI&>eQg3B5GZ5g&JdV467a(3]Z=f<(ecE_KB\
KOLT)X_BbAB1^:-,XR>C?CX-7EEWX.(.1)8/AL>/773W0Z@-6>CDFGY.g:D9b469
<D))JCZ/HV68JL(0K56W@8[:A^.#B8]EZGP/A6T.8,?>gKgS>V8Y(Q?b38()Q-WD
>N:96O?R_eeU1<]@PaT,]W#1ZaS00b;)AMAP5bg6=LC25(UQ60>\LQ&GG1/)=59A
J+3KWTG4>S-aL[&30c;H_Q)_\FYCX]?;2@bGFU(?QV4>>0Y<1YK3EGaC@;P3NF.D
1,LM?8-=Y]@(6EV#EW=_ZQ=G9M1>#T?bCR9Pb=MM&32K?@NC>TM[6>4P-H_fYR,E
:Uc@b.26TQee_aZMD_gdQ=(;#=M[P)E#8_#;Y;VK5,E@L\G_>S=g/Z[#U^B)>@TA
fOO.Na/0e#eLQ;S_MK-&[2WIf6\ScAAU.H5=W0<>(C8H_4XFY/-++@8W[87(3+H2
E8U>:9&LU:IAY,AFURV.<L(61>.N=;>9^a\MgPNR_ae?J\@f>3>FCIQG6LPD_3(9
g:]0CL]S0:DK1W^KO-KFJXL<Y0<_WU]./J1K+CPTdg:_9=CI:>3@,HNXUe@1;L1^
JcE34ScN@KegJVMc6?VN:]LNgC/M0^B@9/HDVU/08D-:P(RaE7-(-e:3M)3SL11M
(4:\Aeeb9ASaEDWQN.B=4A@;IfYEd29-YI=-,YZ4K&&UAOd<6Taa:3/e#&G(((0\
(R07gN,ZVA^J6f8G5Ha9Cf/YS6F)O(Y2UHZ:RH]A#Y@OQBMICKU23\Z91=2_S.CV
4QK\W<2<XNQNMeZQ,::5V?+3D)8711a5Kc^c+X16fa3Z-B9.\N9\PIX(7/\8(=-K
S8=geQa0RE\c)Z#\?dI=7@H27^]U^RHIR9##QUW(K#)RVSW;C]E\#H4VPdcT0_7f
ADKFbQRDDIY9]+(NF?ODL<MWT4,2e7PF7P^ebf-]^7g@b&GRS2)eR;S9[+D2OF^=
Z3;4eXN5_4)aHGM8(c=@W]_>GfLS#L1F+5A;Q:\ZD,3350^DL_dA#WbC4.P(aV,+
bZaX+X6P54PP:4E_&1OFLbY8Q_>Y]G6&)d\_PP[4HZM^g<KG;(g1P0_1-^9CJ<W7
Bbe0W^:A?.VJ1e,)(a:4)dUa1FQGNV>ZH,35HV0#fbR_g7&Q3=:8263CDFSW1=?N
M3:(4\#G<^gOTP_=I,@HB#S]F&W63Z_^WF4OPZZFP+b,cIc7\XX2J)]JLQTHV3-8
4.f<7g>53?d[G14UQb#^CR-P&)<OZb9DS>-cLVGJJJc.OTT7V<RT=fC7ISGBAF=?
G)9QM:H8#)_?6:3e_)b#[ZY>D34^8PWSYBfdHfP+L1]cIWUC2.Ja<+0XV-3gH,C.
7_ecc9WLef/_fE?-+U7O3P1EgXY/@I>F=PWfQCG]):8OeR:<EK5Ge?VT(:)BGe)#
-=;gMN6@<DUgGgRc@#a9JQc>^JUDB\B;T7Df->>SY>-6NJ9E&?7(R/?eWFJWZP+5
/GYbb-9WYW&NH\bJ..&@RC9#^F:#eCC/ZU9FDgM[G_1J??32AIV(F;8:gF&^3+gJ
[_36[]ZJ1OCCMY3XH/aeEe>QKFC(c#OD]Q(fHf5?0CVR_JaC^(FGeRe2I2BaK[U5
F>#AKePG/<O-FR)F3L&463g=),]<Y&:;eLEKJHDJfCFHD&8>QI9/)F.>NT=7&fK:
,.LFL_7,T3O9>ZC/AVF:eN4R,&@]B_&R.FfTYS2C]Z=g[SFYC-9FgR7D,_Qe;VRN
BG</P,+<W)MQ=KV_]5E.-;/W&60;:P#A?\a>#(1X9W:G>+?TQ_3C-^_ZcFK(EKeA
DTg+\>#KU44Q[bJ&I?9OQWCY-OO9b1b8ee.KHe&KTSY/WAD&f9J=,9MD4]_UA?0H
@([)^LZ_C>_O1dE^O:efBZGG[fP\YG4X6fb9P3R9/1;E(UA4W[JLRgQ+MEO61a=_
KZX(WTbR)BWUL0a<O7]+<NKARWMN:C?-]LU;N>4160_Hb@[)@I#R)V8ASG=]6cR]
00]e0RSTT9.6M[gY@<M2^UB]?M@D4,_d,&_,-.]-c242MA?9T1,)X)56<M[2(GH6
K#b_)J=@DVIHU<HX]GX#&Ud:4_7YNf;g]HDO)]77N)2;1UaabT4\.)^?2IV)>V5f
QQ-^4]WZO4<SGd9>6_4,>5].f646H7)(WRG7I+O9b.],3G53.TAPPQ(W;1DK)+XJ
=W^R@]R5-\6TUc,4)f5SR4&f&gO)..BM8.fX1[].ag@+QI(1H]fYN1f0/GQbW/&L
:5X(JODV]Z8#-SE55G278,gJSd:^^^#A_4(dRI0#7@.)-BJc6Z\59WR3Ce<J1X>=
?bEa&cb=L.X.YT/X7D9&#I93b+NGef&D0\bE6[HIa<SONGE&#;]\QTN7gYWJb63E
J4R0-Q@.f6D-Y^c3053cYc.,Ac#O>,g6V5+aE;V)J&@#Bd-MUP\\<ZZMA2ISE8BK
X1?+8]):Q_G[g+W1YZ(g.0?6LJTV/S?I=DGcQORU?f&6S;L<c@@H3-E+AYU4L[ZP
+=RD]N[Tb\EKR,Z+>4a>BB7=/ee2317QaX.V2G&JN6bdd6)]+b<,eJ,fA8/G<MMZ
SUWMd-22[J0G,FWF@312_NVPMS-Y\TLcE;]26I68]:U:Y,)@A\#C267^MH7)0cX?
bRNU75T30KW6fL46YdVJ>.AI<X20Vf=#a<S:/d.aWOCA1;:E)YOc0UA#5/^76=HV
1dfF.5RVJ12OO5OG&8=_ODf>#Afa(B)<\Y>O3a3=O:1cDC(9O5)fR+_JQ_(6;SX\
a;,R5RJU1OD8]C=YFCD;@R8MbEFH8_^Ce&>6JA?AE8S<2M+\GBZf@0:W;W[6Y8:>
;bO/>PGW-XI^Y+g#8TCV0?f_][GL<1RT#K<YM[NU:5+D;73V_<QfUKEf/;J?dPAP
WC&E,X]AC^J#P\S/-\NG&(MIZeKedQRa>YRUQ:3CUUYW8B,8>:+>;e-M4EFfD:WI
Sb94GL>:9#]I;XBU@7KM\La+E9VIc+LbZER;HKBI5PRg_S9bOJg+F<^\.,45IaC^
+ef,aR@.+[M+IP_KV6;V+E-XUTb>?)ZQN]G^dFO14dGgG^K9eMX5K[WT;ccRTGH4
ddB_+4PB(=16NRD5K_3gW_QGCTa-fVc[86FLBdNd1a9MG7S7V6J7H&I=0>M#f?6Q
CNP>1B;+=0<e4IVU]DINe9[FQ/D#;/H(UQO+DMADN/_c=eHK/3724MZH.PHM+.3I
X/N_,T)G^D8>+_<b[14WI+F^,PWA=7\U_-:]M-SYYL<a;f#=HM[+8XfLNH&W8Xa2
&cSO^ZT^>(7g=FUZ?K1_eNF:B^fH/419,KI>8,89S7\e;a[K[L(OS-\V7PE4G2<5
fdYg9PBN+f;<;Z+N/CJ8HCR34MO#E6=^Z)Rg=(3a]H_P,U23(6?MR)aH^A1E7LX#
EHbYS@W_Q/H?E<4#KSI\K8cNb9U5Y^MO_1^D<gDMEdHT+XSIbZ@NO<I8NK;Q4Ub@
+5K1[4&CXXS5HHb42[TL<RbX>F3;K0G&4]Mb/DD4IDGWL\c5b67JDYEcKC,f?)ZH
0N]I0+UVV?(E#;.X3bW;_DKBHCEG0X#?J?/:Q;D8HV)7/L3Yc&=8^0^#[[\6VWH\
;>A1:;dgAC5NSfTY/[+N3Fgd(X_;eA8cf0PY<5bBM\]Q1BYX\;DA#HU(@>(2-NBZ
31K849.O;3fXMUFCA.?YJD/bG.,VcX,a9&K;VQ1Z(ggOO]@bbFV,g<KX3Yg\eZ;;
]_0M-(OVGYcE?C=A5Z\3RVN<dX3a+Gb0bRD(gIcMgeLJNQJJN7,QR]b@D(_FF;&[
S05AUC^&@XTRV,H.TQRX7/5c]2^.\3)<bU0\e_-9.>M:MKWS[AJ8\Xd^Ng@41FA7
S#G:/@:1]f(@d#=e;_:J2](:SE:SD-)dX/33T2R1()@^R6=9fJSZfc[CM]9X.4<^
KIO#8J)7&J+@L,@La9/KDN3DWO]/_)M[f=54/K<_F#Jde65S.>U>@MOQKT@28gH?
+2(,DB]D_&,]RK;gM_\P(bc=Z8:egW(_U\dU5T6]VS8JA@1#//EM,&I/La.d9N\T
BW\0UV5RC=28H/4-M&WP]TLabc?>aE(?8PVMSHbE&9T+bF;HL/aUI^^dcR99S?Y+
GMTI.8>(.J:U9/I+b6E+?:aGa8e4HPfO7YB;-Q_1^0?g03E&NI=MJ])aFe#5FEF1
R03;8:NTEOV_#&[M4U(2:fb<PC+CWAaJd6-Og)K+MI]e-;D8?S[GI-^c\TWM<:O7
GAfY^]e_/3T2abIGd2JWJM>KM+&F\>b0gULd9d+cC7\9Gd&QQ4UM+[F[Z.2R4JcO
L6+&;0.):<T@R/Wg.)>2aI:JFBJH3H4,CU7L_eBGZ3I+=U4b\)?LGJ@W,]E1a(5L
IacRfJLH6#JfcY5cLMI:M@><\[]M0-[3?Q/&dWY1cVPc.UG-X0(\:a1N2(J4e[+A
UQUDEb>3<,HR?1QdAH7GJK7=C_g+dI+aXD7/G.-TBGT.F\DT[JO/IYeRbE4OU3DQ
?EER#JD=T5YC)?@37VdP1T05]8J6Td];KeZKg.7DSJNc6P7+GF_:/EH;IJTDXQL(
68O:S8/;(7d0LQ<8^S9g1Ld6PSLc,,0bcDYV:S:6.74=-\GL0W(03Q[QdJPdg>B7
([+-6\=28(8P.R#M#COZ29-Z(USFWe\ee=gZBPU-L(91-2?FWR/R^4=gT1;&-[K=
D(VebeRQER0.QV^cU;&O.DDS.EL.(&&(1@<JW[.C_5-bRcG9V9;H7e\[9(c6fADd
V[gS]=Va4ATV4HdM=aHS?4e+/;N90Xa[W8VM\)-@AdO[=.fD9B2^=a[DS[\1=5:@
5WPVK4[Dd&^:Z5D#fQSf.(D4>^U([I>(<@g,RHLNK6g2e\U1Q6<C1(W?(?HW35cG
ffAH^\ON_CgcO0ea72JP7]3\V03/9d30.Z,OP]:dIc5R+O.ZDB(]d2]_0Y]>2ac1
07a+8dKHHG#\=_1;-2Df=635a._9O121AH&F^X.Z2fBS\e22\6_S^HS],ZEbQ;f@
>-L=)2/(2JNM:CTf6@0\NQJ1IHIQ<+;2cedX98GKE0RK)FE6424TYc#X=F9+<(C#
VKU-c6@eg/))WJM_5PC8HNI4OF8G8YLeYe&8TE>ZM.9+RKYS-\^M<#?,EX4MIP4L
fL/A,.X36[GG3AT6L9MgLE+>\F,4:\SSG)9]E#S7>75CU-7V6C>/+IW.BA7;02+7
I77=EWg+W[4D1gCgA;/[a+4:QGfAQT)LH8a:b/RRE^=U>M<M1\,DIQbQW3YQ<3:a
;_LQX/]9<0Q7/FC@T_\=0M1.._(UAQ[2]BD,d4Q^[?33R27;AYCCO[YdD5XeAG\>
&-I9Z^I_+#D++S7G^R9(5GL_)d0P#K(SIH5M^E5^/_4Z:&M@@N,B.gKUdI<_5<W:
Ra>I@0;S4H.Kb6P<@.S1O]B]<fXDX/\)X8=R-W-2LIV?MFaC_A)N\4@:L:I]aC55
=/W<c@0C-VeGUY(MLQ<S>(SWg,]2aH1)_UFTaL\S1E)cO9C[R-e^#Y&D2[gVU]IO
SD4SQ#&cW>/HGZ-NY/R_7ZGW9X8,g+8#E81T;I[6=78dP?68.&1C02D++?WE+#R,
Q=+X<^3O\TB26^0A?9#>VF0CJID0f-+.2<)X/ER[=BW7g7Q__2IIf\#3CWJTB#]S
-GTM+D8f@12)ddDUf@O\&JR:1Lb78Z#=cC5<9,bL3[[8264=?ZfG1CP,UA=>@ER@
47WbIBE6&P:8H:VKZRHYJF7I.<6WVUU<HR?0LE8Z7BQ@[;55cBT&f_PMFGFb\BS/
C\Q0dWTCEL5Pf<6faK+)=KD9eK7+:+(6;>gTZL8H+/W<L5UJGaM,O=L9:Ug](LO7
E1&C>R_RR=;.E.@0K>GC/FVdU5E99/LZ/Kf#+b^)Qf/O2E>Y]=IFESQLOKZMNUPK
X8#>+(>Wa+()D+\,bVLR2]MQM&DQWN[835HRI<dV5F5;]SK<5QI0ADe53)dRGOSH
/fGAeM6AEcW<-I9U2ag[^MEb<BbVBT-a,<E-/E9.5Fc1Z8&0ePXP#)R]4X/J)(+T
cV:UZLX<NIIN[-Sd>2g6F1Je9:GRE3.XS;+HTZN@[G.,EbLM<DL2aYSVV@BIL9/U
+.5T#M6I304O04S?O(8g4#.I[_K?g2C1L3F06I1&KS)\3a#L2D#-PJ+fN3/<\;MP
AF2P+^#cJ^c>&N3[YOXI,Pe\78.;X#JK)WQW>@Wa8[T;E,D/>]YK8,5W&CKVOQ;&
XA1f0TS^?>7A&;]g-3+XMb^&c2;USd^9UgeBGg;c=JPJDY(5Eg\Y]3E>SO-QHd+[
JVAZOgU)d+,#COa037I[1+2gB5R/(RTWMOD4dZ+KWHDMIWIF2^)74EBI)8d5YQLA
32a/2FHAE^dSCF,U[MBSC+89:=PLA=eO;d&OMP[CJH&dTV10NE]I-D+L\Z[(NbK#
TY^.C6Ca[L:A(gMWRa4H]Eggb(4&-f.RV.,)<eP(HA3f_FPCYGJeSXGREW-7L8(>
bP])R_LJ1Yc7ORLMUYagb3)]3<;\C3,SfJ^;2c&?e+>f5S=D@SE^ILPC;O6KcS16
T1ac:E\ZP[bKOEegdN6U>:=I[.N_#C2+DYY]^89I)[V=_[30LKI&8\ZD?FWJUM1W
(f63^RFQ6&7;AP&)LMI\D5@4gI2B/#5J,A\1977DTc3>HOHK^D\=#5)PS38RCG@;
,b3>KD(e(bB.3PP^RJJ\fT,KR(4?QLf+Fg.P4#8c3FGR2?V\c>^>a#PeD[>[+fSe
e[KWB7N<,2V^T(,E.(=9Nd?5^@/V0Ya/(1g1(^<#QQa+HEe-:#]98E-U2NEH]EL^
JV&V_aGN-PE4R==,Sg(>+33A94Y,?K>T=7;1)\S&9dSJ_-KJ<,&_J)=H0E91,29&
0+.@>^fR\Y_A5BCGX1A)?(YW)[[6D)Q.bg6:?gIg?,B=0>VD.A(SBB1.eU_[V(>X
5a/g1TB1>)Tc<cfJ+L/+Q9=RCTV&I>47>Y@SK\cMJ?Id^H?E(WZGJ?EPE@P3(.LT
-2LaBZS;U\V82@#]/fM@d1/]?_H-FTg0g#Y,P9FZ;1&1]_a7113cXX8>>2<(Wbf4
MXRZ)5859&:(,O^V45P:J8)+2Fc\9[2&BUJ409620@P6AGA#M6N86W(_J.SD9T:e
9^WSK3)N+:&U5a8f6Cd(<X#;O1IBB_88GXUYPLB#AP<VYd?\]N\K^8<1=@<#aUgK
67+5/9WBU6#O.AY)QD@U4-^X_0<@(:]O]:[RLNa6U(A)S./=-K;#+fYWbW]1//P@
(A0CfbW&g4R-W-GDNFE0G:&](WA^P8-Z^[262:IP=>)E;-GL=/EfYa>8f<C6(OPD
TJ/V8@ZWDBT6.P6HP7?6;NcPC6XRN&9I\b\0^G=c@FR@^S_-/T,O+OBPX(KB4.8[
61gf+Z6g>#dbBg+WB#G:#:TKEUC/g&?#T[D[_dX=CJD&3OOU2dZ-E<1UZD55C=7c
9Mg^91SMORb&.8QLJ,_.?Z:/?M3I@UePL0\K:??TS^\,)@U0>DGMK=436dLW6IGW
AKP;&TM.AbFKe94,_(?HNM7DfMgGV-6;E@QA0BQ3&;C46,XTTAg43O=B95O@/-+(
S1V_-g?[9(?b75SJ#F-eM)318IY#+2KO3\6NYa#2MVT2-]bTK[UU+gN0KV>0S9KG
ZD)J#Ob=)92126;(T9&.EU1TL5DHUD6FX&,#WR0NQ6.8FE))G.BW)S9&(EN1/AI/
-C^0X<H4]MP#62aUQ=e=Vaa,IdAWCKdZ>:FAD-cF748(KK:.D<:^Ogeca@@S]gb^
f4I-4SIF:.4gBO>[O6].\N]K/AL(DBeeDaW>b7B_8-#+3;/MRIMCJUE=cfM5R<FG
G:YG4RBIP<B<.7^;.GR]BRJCD<,GJQ8c\e.20&_b];S43Z\IMHc#?#d(UJ:[,L^S
S?=D-e@:?O<GX8Y;:3BZXb0YE.A^XCTbSQLXbI;DLT+/BFPU[/b2SUAY@>3O<YOV
dU7e_A_0UV8<NR9&a,=UQXZANOV]<(\Wf-<J&B[V+Ecacd-WfD#<:?DBSG@HcM>d
e)BKU3\5Z3:RdM7K6]MT@e=EPbPP/I47:RC@-SdNOB8bE>b2eU4X8a;CC<+.?=0(
KA/6c9Ee[,F]VQ=WF3X\Nc#L^@UH==f8O,c^g7e2R4WGD2K&0U=-VR.MT-bFf>8K
;;WC7@dVbbR=P:W-PXGZ3120I/-G^e/?Sgca)gb_U0(NdL1+b/DMc3(Geb6>OXe\
Cg0QH)M-N1]4<I8=-^Y,N0=;S2>3KWX0LS,<@;/1.KO2M:V)9gRQ(HAA&[Bc3XWZ
V-H4Z)P;/ET0@9&(e@2&Kf[bRY2+aBS&<].PI.fH?(0#6-PU]XPeM=5#]7DN9cAc
&HIeHT[B@LDV25>1)POP[6RQ\@1.SBO181&-WC@ZH>CeFb#_7378a^g[NfL>LONY
TGC5FcB@f_ETf]J??WQUdX1:@/G80VGMCJ01?.f/R@BI4[Mg-Q^C+#c;IMNaM1ea
2#UUBc-3_/eLc?ad.=a]BB@#O#.2MJ0?CMO_8eV)b+/\g#Z+-/_LZLGV;aAP#\#4
d/gd\O<7dPQ:GfARgO@U;dVeN5/0-:I;9HaLJe:c89--9;XKS=-L4eY0=W<6f])c
5644bE;VN#R<=DHKAU#d]1AfAFg2fV]c:4S^E::W58FCKIS:ZGZ#]98a[eg-UC_/
6H0?I<_a@82M^>J^0?ABLdY_.U(0fI]Yc:3cAe<&fT5[O[#PPg0.:T2\c-B96-.#
&S\?ARS0]AXXff+2Y;Y.K:KGIg2+R8CALB8_O#ePe7:#1ES?Ce<4P[;6W8b65#/0
gYWU2_Gf3CPfML_9.=6DJU)7^:1P\7O)H9edW1U2T\XMY:XOB&(bcTcRd5M]4_@H
b5ea1>(2feS2YcYCCS>Y(+PG4(1O/?E(Tg6b0X&F5QE3dIW[/LA:=].B2?YR#^@/
.O6Me?YddSgBE9#=)?Nf.>T\SJSUT6GTC4\2^L,fD;I7SZQ^gC;#fbJGZ(KZJ>QR
5GS_=a\]^MKJKLQ-3YS<9(.a11cPVL2DXQe<,65MQFeF_]QI&JADH+10fQ,5(1J0
-?EfXcS4ME@GGdb.OI#O,ca?KZJ;fgHFcQ0-\\]g,WL-=53gHe&1_\&PMIW?6]A6
e67B;QF]1C>#?2XaSb_H3QA=Ce2)gZKF.3:WaIQ&\d@;)MJ&FYbE;aJf&TP53Bb:
^VS1ZfE-Qed,MQS1BRgZ/NP>+^1ID0IRGd_O.IV3MMY>,ULTA9D\R]7ML1LZXg^W
1X];\Jg(>G8^T[HOS3&825DJ<UD+e4[N<=LV,P#W6g0L-4VG?gDZS?6Pa.\#cd]5
COgNc6-B7+JUASY<8D9>UHOSDgJ/.8b)X)[[B(0?YC_89N[LYERJ?GWbd_K#O09@
+K@N9SD0?3_YUd\Na2J0CFJ7^(&@@AE6<+QYOeUd<e2Na_TP2UB]6f;.;7FH0H&I
+<Q,@V@8:3Ega>EcUBH(e(RCb-RUSD,A86SH1KMc=aK8:,[3;8^\W^@WF(^@SdOc
gI5K@I6O5^61\P?e.#6KWFLBOR<T)24LBf/\^bHK9(6Be)YG)5Q9/?bd[^;U+M4/
UJfGfgJMEK6X)<ePNE3(CFKe(.Y[9P)PZ18^4+6CD+a(RbM,3/)/_c3[aU0<Z:;^
c7M^fV@dX#XUV+eP^eL=O4#a19&f4^19#(\G>PaU,fH=LbL./+)WRCeT8@gf3\^]
_?/_&AYLg,aL&PQBcCUI98Da^681(bG[6e0G&8ed@;GYMXfH?MINQ=5701)AOSTD
fZYPB??:Q4bQKA7f(5XOJe<Y#-_f#W?9[48RQ0^aI<>(6-0#W4_ZbDK,=a^+TKVK
9L5eG.SOX[>=SdHP;^NW^[K_\d=KG63a;.&1Z(.CJLNQSfJ?F2Y)X/OQD5SaffE:
bY9-?_<Wc^H+?YbP?IfF.fC\E]_/(BeMD]WP)4:bfTKWEg2(H]TND2d^1_O)&eAO
65KUgR+GeB8_G./D7bX^DL_eXJ^G:C=Tg?V04&/gCPW60)VNfWPJ45S@>\.9dBSD
LCJF&Kd]Q5XH\YAG138HUE=Y:]=&KdI6E)V9HOO+G6RXWUCa_DS(ZY@NYbX#c(^(
GGL[[d(88]_Ja7/g6P)<Zd,bEb9HD069]SP4B(@F3aXRNg0,J^LDa?=]../6#PX9
T]QWOb49Ae=T5_02M?d?;ICH(M]B<S+aWY4RE[+^bV_+D2d;Q79VMK0a6SWX(3OE
OE^g-\CYKXGYAa@@Q=bg^O08HAf-N=A8C?F)L;aDU(Sd5P;&X[T20<NPUGe[QJ-X
fM8OY9cYLK(.W^56&3T5KJ4HG+6102(-DaMSE64ZQf_a2BQ>=N@JaU;)WDCT9f(+
2aIOc9b3)d]SI#DGZM>dNU25g3MA--Y_Vf&:G+OVeH,8S<XeGPM];EdZOPe/?fDN
=V:<^CW]>f53?JW0;e^X9NRGf&CT.S2bg/YdXb9N?B&X5bGBOMWZ)>+\[DDRB-2a
BQW/9JUOX3^UN78:Me/)-E8:08fXJQOF0]U2+g.O2SQ3.X^CbD4[:D;GJ#I/9aJT
?F406A(\;7O7N@LbCJ&4+E5R>^b+=&5>?E#I1<OZ^8XCTV;B:0;:S</?a6F/a7RV
>LE<DPIXSgK6NQ\#_0O2D-^OIPW_f<=U=/L86KE6AMH^=AK:CG-\GaXc_a,[IMDa
Q]M&7@cJ_B]SH_+NgDZLL_:Y[J&I;E,XVJ>ePUZ3g_OeYG_/XQ6@<2a>H9Y[)VXQ
d/+3,?MS&N[MaUbWB?FW(Ha?K8UGBe348,Ob[]^3Z6:Q28O8H]L#_0]f\:g;U,1#
D\T+^eE6f3?2Ff\f-/90FSS(8\1?54f;B5P_7)T3bPE?;2RI+?Y0Yg+FK?aXE6?-
^^@<JC)[AVe=&1+QgZ8)&f73@:I+a#7CZ\ZZN-2U/9TMPT\R:[T=^CF^WOP#V2cA
439(/]B81E5(5=9EZe=c^Re6265GgF=c5]H(OT8#=9_bL2N:+?0RCCT4RC>#9)_)
D,SB:A1b21.<BX+ga8cb:aL+YLX)#00>X;R/#+O]6cP@AZK^DNBcb<.@0(J/@(-R
.K=?JS2VGI-#F@8F2OfN:[(J5V;9fcRgOfC3]IEgBD4.<8ARNZS15/dJAP84#:/V
)WL.3FNCEF.:dfDdJU)cZ[J:aA(:@B.LcMG]d_9DRU-LY/27.V1_EKOBMVe@cb;@
@T27=OZHYgZ?<;6)593>[FB[R7R72E_;046<(>G:D\0N@GLNODZ@g7fEOB6)X34H
@851&,N-)cQK0C4#?gN@/C3N:cKSbc3;[fWa[?SZICbFHDV[2Wg+aW==<:TZ)(+d
OPIG&Wb.<1^)c_H)d,=feYN[]-=OAQCg=Kcf(85&S4:+-3Y.=X</J=BPKLLS>9B2
LVLI=_3)=CQbLO856+W@gd(93<6b2+,C1\,OBEfQ#-f?JV,ag##f>V9&:GG8><O>
F@3\X(:>X;R0.FV8JWaM-gcC]^6=YSUGf5Z+5[@e_Y;:L.PIZ[GeZFOCdNddfBT3
XUM\?[fH^R2b0]--5O+LEY;^PSA+c:OI6J-Z(89NaJ_T2#OcU8/5@QMG;7HQHZKN
5.H0f&A#5W<66OBW[A4BV3>9XT#VYOaEESUZT\(UL,;3Z,]5?9=06HgJ>)L<c#Kg
84XMMa<[>I,Q@FJJQJfH1^7Y<f+R]cbcZ8E>R2;SA4VeD26G#Z3ZMOW3SA<#YUW;
/7-gU+9gAEQ8FLHbZ-]b(VNH&#</f-3)5ae_AMBg0D53fPMe,.Q]9+O>YEUL96;8
?8aLOH>J85_+9ScK&(@G+CdD<):)F.f6\cTKXAO>eB4/2\-&51VA;3gIAC9:fb?/
SRD]02b^2>&\0+5X:IU76:P?YF0=<MW?G=#9B<7IS;W;<bA/KJV5=a@_+EA^]Ug8
0;W^7U\bO1G:.aB@A&R=#\NP/V0Lc8^dTEdMI.@>;)W]W[KH]&&E^MdJ/)3>ZeH4
QVRSFS&9/aX@#M]85Q1/DDFD#JH8A49E_ML3:YX]HbK0-Xd;RT.AGg2H5MV\3W(9
A;0N2d)JG0[Y)#WS-\5[>ZBVFD<CGfO2Dc4dT&<#GKOMI.=8U]e=5.)/>;,FHL16
&5N,PQA4T^cOYCE:Z=+MaNROW_Gf&D@1_]<>8G+bJIK:SegcL0RQPGdH6RaL&=Zc
\e,?\B\U[19CP@e^fbLc+>W3_MQ72(7\QV7.]c-N,9R(;?cN_[P<cL/FVF(Lb,dc
;5Ta>-0e&82?f^[D746V\ZTZX>g=Bd8=:&egHOHg/]_9++;,N96fLGB682?,cX9]
a4f)?c,Y+2)RN7fJAB@Bf]K)9Se@dP=^Y>#[Y15D\&ScUR1..\f<FJG327;/KOXL
CL+@VO-T^@DUJ+FJ/4db>RD6]/a6IFc4e\4,V6;IAKG\DGdgdHK-afP0VUH--)/0
LeU6EVdX]@-7@W1.WYeN9E3PE6A^:G6Uf1A./Z9B.^>E=QUUMS1+W#L0.c-@H5>U
:D8\-=SBC^-:P=6V2IC1I:J)XF1KbW2+ID?I>98)RR9[,5J_32=9)V)0]-7d[.6?
_LPdF<#La.]9J:C4CR7]Id]VDIO_K/H20d#C/RB^(Q7^G]H9&^R^PC\P<#VF33M#
VCHa7<QVWd/?Rc;/4H3FA+g1S?e(X#,IA7+3I32RF[NF\H.dD/N)U.0HPFb4W0^Q
E?LNd:KS51#XKBOV0]b0Y=Wg4J^H>OHS3V:3P&UT)-PZ9?gXWY4,&b9Mc/,bJaA;
0(KZZU:P^3V#Q,2/+>O99V3_Y6gb[WXVCX,.(+FHOVCG\SSc_]=5_K=K8>Zd/<eN
NO;7.):4HC()bP0CR9g+3efYcG7?G488FRPHT8[fYFcQ?,;)SC3F4V++#@;?<5^;
ASZP:W]SQ1:2&TRHWLUP#6U<K_Y3a=H2@/Cb]5^cY4gf6-9S#YA5OU.#NbDB?4;[
R+#9,3-)aGNL\[4>CL9U&9VXR5SPHL^NV7S:TH1Z6Ue2HG#3PV^Gg8[CZK-SJO@O
[MCAebQH3W./][eCV-4B[J1eEG9#?G#F_#HKZ4^DU2fKXgC4J6?UBF0HR]I15KN:
A.A&=)[a5-Z[W?6]XMe6Z:\NFA+&cF.KV]WQ1/H=/H6G\ZK7[HDT?0_7f4JP->@F
S=\d;5&.1Ze(6^WSfY0A1MTMHAV3NN_-TeF_AI2H,WH?C44SDFBC;P]ULF3./VNC
\TZ?/fXScQG&(/S1Y8?BC)e@@2XI]I_^1dgI2)MBfF-W]]&JA@P73:SdDcWYBU7<
IPEL.Sg.^LEHL86D.ASUL<C234_I<.\-QRQ>e1XE2S^TO2H.cWBQVEUOL@XU+(G,
d1P+,f1/S3K4ddX\c51H-5U#bU<a549FS[b2S.7D2eMXWTB=Je[fc0/OHL13LW7B
#d<Ac>Q>[R8g#]>1+1N,O]1UZRIaZ;O?;edeBMe#>@G,cN;DeIVKINTP>\Fe\-<-
[Z.g+ZXEIeS9M3A1Ng=NIf?);H2S\/3IdZ3Q3c_1C-AD-Z7P>gV.W(6?e2^dda7E
3fAKECSEAR:YDATaL1S.UNI=LG?S;3)2A5._]AZbUNI:WJ-Z1V@<YeMUT&@F_N5_
Xa]f3OJDWN/ST,>RdNL)8KdEOBES2KZ92E3Bgc6]df7VfQg9O(T3E-&]W=^F3@gd
>\g0E?W@?PCX3EENFNF:,,0/6f<9b-TU?89\(;7SJ;>XX(04LA3=,-Y/VV05F(.&
O3.(0D?f^^@ZAcIHUF4-OVGDOT8V0MH(#,<G=S64PW)N=_/^_11E_cC:A^X>4/=c
(2FZ64Q:?GfT]8G]_C2CWBc\0fAf[HT]dH+-E&,;LQD=TE8.I,g)C=#:LC&We@4K
M85aCJ_1;9f=dOU\MLfdfP#(^fPA#H3HbI;Y9dN\6[7_GKDBDgD9?=/IDCRNMOWG
?JDa02_]@@@U=;\WIX)<PFU897R8_gVeJS:PF)22,bV^WdL9V5?7YFM.IDIRHPQZ
5dMFL)>;S&(G93X4dD(eZ7M3=V+E1BH8_#HPZ;<TKWfS^<dVT#_7H=GAZQNg]80/
BN8<KgYSB5,X^L6Ud#ZSdJ+S+OUVW1G+?KYB>YDW3ZIb7<W5ABOdcOC07I\7fK/S
e1(e&@@dN:gHaa6&fI-/31gfKN;28>I:5+VZ^&WL<75ICH+E46WG1:?+(Ib&FP0a
dGD(UA;a2E/ZE>)2H,LdV2+X_^>+<Dd,K@;aFP5dd=,#4+3eKdZ0GOJ;7Egg?(XS
91YZMGQ90e54UFV5R96(VWg1fLT;9U]M9dA[:3+W?4OK37^S&958OXV-#d+c17O1
bUY)3=Bb&453-5(NL_I3g3,4G5E#I^I1H]#C0gO]@f:4H/;T;BRN^gG&G[5^[V;9
dV-3S;(dP.M=^.7DQ2Z2;bBCCUc2R3C+6B].X7I9+XfG2\\G\8S9/JRa@0^P3IY=
4A9=VP19@7<F#YS=1)L03@a#d#fD^.SS2>\BT]c)IL+CZQ.\&?aJ_LP]N5+TFcQ7
VSf[(D,8.2/I?0VTM04?0=RN85C/LEYZTW2S+bO8A?bRd;H,+:H5&D7I5A3/YW@J
41QE/O8O]\Me8N#PM_eUCTZ_4N6\XXdO74[^CSb\C)dgca(a?ge(ce_N^R(@&dUO
][XKXFG3U4ZS/F_9;b;ggbH@bJNa:BS5,;S/CLF>fNCY-0/b4.65J7MfQFX)7\.5
OXI=^<eP(1WJfDd[8U2,CZ[BT>gZ=\)4Jf12cJ6ce]eZ=Z/^FM8;e<R]&)6FMa27
0JL/G?f6L--L>5@Y:M@\?2\KR/(.UJB#CP51R(LE6g3>5XCNIfI(/7Q7SdJK5M)Z
K#E&T5^&6WSbCL7^TccdY4)M44\5B5VIQ8Y6eMS(W@^,4LP]N9#.<44QWH+B]5:Q
QHe_4E.<d);NPa5+E[+?8#39Cg<Td[ZICagfU:636O909>LL4W4QTI2N:gO3MRVO
HT+\()V=gf>Xb-Z(QX_23#:3(N@U22Pa+/?_g4=SS]?eb^T]XKD5)B21]fK:Q_5Y
eT;gQ7?6,dYCA^Z7:U/V#8bT@5144g=]83+d-KM(g#:H#WD=]YX+[2A0@fIPU4]=
\6@KCH9[B>\Te6>Y<,I3C77Nc+MZZ<CWP2+[5(bA@V88Y[Q6T<^5,M>6?D7)eE;a
#IU79f9Nc_.[VBG_W)/7HXZGg.)cM-aH/V_bB-)+8C492d?E]9ZXON\FN4cKJ_-?
N]EUNI8Y4M(fB\9M;gO\:C-VeKI-6[:#0UL2R<b&9?IW>L.,E&7fTeNeQ:#>c[@/
3H0&Z/G\VY8=1)f\S\N3,A+E0>/)GRBP2X)#&^a<8+eSgM>a7K82\7e.L?]fAI)H
,O&\bO^GVB0eHYD4S-7&<:(.960<Dg06P[7>75UZQRDdbf_3Ka@/0DcLY\,\SED]
D598EQ[1.WN0PI[XN3J+CFg.5Q9UFC/^S_0cE#\.PYb3YAH0&\eB\WRG<f9(K)L_
LX_X,a<-^fR-_&I;[WIM>O5[^>FM0\N&f5BJ/^2:.PWS,dZNQXcOK3C,QR9V>AF^
5EEIK:B-XP;FNbR<Qbc5-Q0Zd/N,gD0F<g5KU4WP;[GYc#GY_10\]1L#D4&FM]._
/SW5#dbZ2cadPfK32cBZ0W]PV]8d+G,_D#;-EA+>+^5J?8),UN?C#3?]YESedNCS
<FH-Ng_9R]TfG&F+6>]DPQ#QcS@9(HDUScaY#8-YQL0Nd#]]FL=J?=K+[P;<A:TT
bJ7569?S(61df)IJdLV+FO473#S:)V/)64SF;AMOb8?+^[f+EXEDQfa,))KSa0ME
5N_AQATK_>c9\I<?B\A-PS,1eS&],#MdEdA.-N]IRRd2c1&=_R:@:Q?VfDZ&cL8E
3EDDZD<^HTBPS]6\CdMWPG61HFb@U]H=U5&\;V6Q9JC?J8(27Y7@f,B+,^V2>D3K
[GS/S0^HbX2&D4ed],D57&C(^B8Bee5MX/RUU,V<3PHH#BU9Bc>PNP)]b.4(W,4(
Bef0-g_4aP&0#.QB4fL[X^f(EXRGc<cV3f>e;,O@3e:=4f-;2fR9+RSRF.c:=gA,
ZLe[B,XQHNZQ+@0EbS0_7DI\1?T0HTIAXc>()P@5=2\b,eKEE?KM7>GPb2:27(/Y
BN4+AV6X8]-g@60_J#Y)F41IF8ZBGVb0HE(2EY-#fCXHbVEM;FV.NWLK@RD@E?,F
<R.WeW.D++Bc[0@ZW8Z.(L6]e:a/:E<8daU]](3W^a]?YIeE4XTV[[3>[=[LYHU=
<#-6C&KO_J\PM>TD,#8AA0\9RC6:ES.0Ne7K_Hbc2GW#<9#9g+3,(OE\OLA@^bLV
WFY[61-2A(@BaYbC0T8fOR5H([Z6dS=<Qc&JKD5W&HMG?>AfCW\UERJ9_RJ(+d\d
?);J(_\J1Tc7\K\0F>g,[5W8_K4aJMe<S)Ae3R(0LZD,GM+1M456c9(TOac7,V7P
b:D=];(-):ULB62BXI#g?aYA:FPbXgZfS&4a^2M&EZH_Xa_:Q^=,,FZWH+SLB(@+
@J5>KgR;3I73GI>N;TU+ea?O67CbbTEEGM,f46WJ@],>[,81H>AX@-#A2/ND,T>0
I#XO#CDJJf\DTgE&TTH-K=IUOK#&5gWgF4Q=&(Cc-eQ:GKN/Q=L9H3Z>5?>TKAb_
.2<c[AZ]N>(0gUG=d/(5:YM>bc+<RIPDN?6/d1@B8854c[[2E(EPY=2eYR2bE[A\
+DLJ[OK[N=YZIcdH>^ZSX&-f39H;><R/.E8C<RJM=?aX^>KcKNF[G]8R6CE=YSWb
a/9@DZ_&\dYUDR0@8^)KJ:4>fYLK+PF[0IZC&=a+697E]7=-Z5N@NE(IV_OeE0d#
2aZXFcXJR:)^[N\VJU=H5;ba947]8@7aK8DL[Pfc5^UVKG5U/L\=+#CdU2Z,;GX0
C==;50D><P)E@/(S055IdQH)2fdDXDa?:UO;,4gOC5/8T]Nb)H2,K_Z104TgdZ0_
P6Z+\(ce;4f+U(I0MPX-LAYT@S(?MPE3)9W9Q24\>,5LBSC.K8gFV-MUB@#PN[Z^
e;d==(6J+c3LE:<:+1NagV;D(O<(e;V;^f>:Vd_\+,1Y.0W+TbKd^=?GJE@^P[B+
/11E4^Y:3Ib3F+UP1Ke6#_@N9V:a?;Q[0E:G0M.Ud@>/.+:0f[e\:_14)C#5E(3#
<Z;5;53F602&14]g0)](<VBO+c)@a32K<geBW^@M:XG;1d2a_J<M-B(Ag:&9&fPW
^eS24TY^E5cZ-VE89//.R5,VFM=W.:B1bbO:U7+@9:M0TYQfI;Tb?XDJ/g?gdGfW
>4\P(dgdREgABM=7MHcTeZZ4_34K2U2JEX6eN29#4<C\M1_Z,?.=/L7NALa\+PA.
Z\:b^P8V@=(=\c0P#WT7_I4#=3RP2WLLPI&cfQ5\E5bcb48#+\X]<;Q5-bX:f^N1
b\NDB&KM&aU[P^[?RUTe2GbMB?09W=)N6#=>f#:OO=a>-c)MAQ?7=Ggf>?69-HZe
QNI?<<#,Eg#2Z;b9QXL.8Pd[N:+\M&81@T80SX@c<QS6QDJcKQT]P[&c[P\=#+I)
>AN+e6Z5eCS48?5(K::&g.>3d]6cEb8JcL&UST4E?-aRDRc>EfO_fe5d2V5gY9#E
6H)3J7B>)R-d;Zd#_N5-bINC38dDP-e6_[>JYAOGY?E_S,_9B/>UdX_OW>0RRa;J
IS>7=gJ(=cX&0HY[a@,08[B5<J2F[f,cgP7NBHVB>ZcETG?,W^AJ.2=aNBGd?(^T
C1DXH)9W,J=\e.dG^S)AOb2WS,d#?<[4C+DXC#DMZ1g4X4F)c:1g15O2/8G](^V,
Z<a4X-Q:SWQ&[BFd7K6.,c3NL(MD3fR)^^cFAY)EcMbY(<GML?L,5HQG)#3FJ7YA
g08<KMGYQI/AGYWKJS9;\>d-Rg&)b@fG_M5SZBJUU(5,;01D,,TK^UaENP:c#,d&
8TX0aOd3=3M+9]Y@>,a]6R^UaE(;c+A&B@.;1V,<U?[1Ga>cV;Y<14e.+4.];JZ+
5;ab7N27/ge)GNBT3DfQUAD08M@HCAM4S1DRb=bYe._TcI?>WE>33=G>DB;,2-_3
-R4RWR#&9:?=Q=Ygb6Z:c9,TgH97N5b8d=_TA5g?.YR65P\_;?.=1T8?.V?Ud81J
,62&0TbQ(D&M?&22YCd(HT;Ag&g,?)_g)+E&H9Y\_[W1\N6(5.WgTQNGUgb3\E.4
?<W0DY#3NGXY)<T:IAWeJ83<KLcXZ4@-QdW<8b7/-d;a>(e3/QD@27_H3^\+:eaL
7U&:(),cIf2a=Hf4Z#[eNL3/S9K\=FIfUfW8MO3RVJ-f/=8Y?-\EA4>>PWb@7N7[
@U=]=SY?46XQZ?5J5V<CN(A(AI-6ZEEBTaP[7/eF,J3BYO^4_89\W8bFXIN49:0b
=2/@Y2N@P9VX4PCSe)=+]2SQGFF5/e39D6CM:^aKU_7@&HRA<(-P-2,#4fB?J8BY
U(E1:[79^,=93AN,@(ZQ6&KO9f_e:C<PLdM.^^QYf[\fXFK3T2O:F7cP#Z0ed@I_
LJ8FdNUSX1_GJd)]b,1C,-Y&C)1^.A[&@.,J2KE+c.U#d.>\WDd@7FYe.2:PV1H?
K/ROO0S@4b]Eef<@DRa(^MXV]N:09LG>\.[DA]80Xa(QE^OG19_aMEGDb7>+=]dA
@\CV32O&(8:9\Z_>5JDO6eK5ME<dXW@?9XJ_5;+4L:M\JAe^N\;IF=Y6)YD;EGbU
1+]Y?L9JJSg&N&O,cDUOAcd63>N^KQI?9OX_c@[2e&#>UVZFU72181dFKWfY6I3M
SIOa9F4?GE\>UUZ]>4d@)->dO)_)Q2P+MD+7(N3+=;VEQ8P&X+UBe47GA]9MEIB;
a,E_Bf0I4_\Cf0F]a=M;S6F));>1<2XL4B@PGOQacLFb2,CC8.3(&Le0b4X9?5<U
cWaNTaUc4]0BY8eE[Q=O]XGK,[fcf.O^e61^+_,NC:5[A_MH+#&DTb;6Z;I_J>B+
YQIBU6\;\&)JJSID\HYgY<HR#\-8B(QB_AT:\2E]&FNWN(,<>7E96^+\@?Z2X9&:
=,.c<&#F1G7##].8KM#-E:d,>B;&b&^A9)^@b]DJ8EA[:)F459S?/df5,W160UOc
S9&g+G8DE#bdZ1/;@935);8[JC)<8S6\Y>.SVKJM33IS5/87;[=5D+\/Wd^^Lef(
5ROLHdXUATa^3C,ZKIP2S^L0Q_^@R+&EO+LO=S(,@8(P]8I>-LGAX1EYT/?BZP-W
M(O\R6EI(]Lb@YB7(3Uc)<[51Kc<c8N]HgKBP8?5G74_,S)MOB28eZVcb-;QBY=W
bN[DaSef1\>&=&LGR&W8YB[I6gZV=IWZ(b?)>[TbVSR:NT+8<ccU)g>;<O5gEO,e
\;S0>-9DC=X93=Q4W7/[4+U7I?@B.^c7U=F(fFS:Y#MdZ(5c>/+EJ6FYaNI_42R9
L(WG>8e>W;7UaL18/?POCQ3+ZKZI(=D\SAP2UFL.HP6WDf/b\Ob@0O;/U=X>WFGE
ecc9O/-#EVF6XEgNZfK0-9VQ)K@FWM0d>)VHddb?0<C7dPO<<XS25gN:Kd;^3KX?
),aL@E:#5CG3X_;\L[NG3f084>cZC5XW&),a(GM^2XW<a)],S7cF@OQ2Y_[QE<b&
bH9V8PMOA<W=6F]#10J-W.:O;YF8AYUPI[5,V\2,6Vf2FK5cNdA#:2NQ;FgOM;VD
X]0@a4\7W(V-OZcI\EEBX&4RD4Y1-<bKG8==1YdF[ecW=5T11(dSJ;(3C&EOAbgc
VK-42U^#:)_W\bb[gYP+N<cdA5REd+]W5KR>Zd8H+Q7K7BEDO#G/BHf8VC4E&#17
>+,^3SD>1LJR[,ZBB\:A.Y=(5//d3?8e_F1S)0S#8[D:5WF@YFD:XD]S<bZI>E2E
,cDdAf2d<3bZTB/7&,<UXK0)#N4(^1SM]X1g7^9E8<\HXgf0<bMJ07N>Ld#9+EUD
[/ZZTXRFHYf2\J#JAWP_,_U(EG^[V&8HaOJ.b2,4]SeT23C35dWM<]JJ:A^fdEF0
aIH=b4B@+&I7&LR9gY.3Q/O>0M[@_6)eGePUQR<N7OJ>XRE2^#.@<XSHEb1K4EIS
;HdeOB65Tba,^N933^&S-aQ+5CKWde=egKfV-M9:N<=#?8U(7)&XG#;N4g5NI^4S
+W,ZHF+Z,@X0XYU^O(H#VNLV:^H?Q^WDb7?H:A2=KgR.e_2\=a@AZ4RIa.cKL9DQ
IAGH81aH+,7D&0<]9]6Y4A^=-c9:;:Xed],CI<gZ[Tc\a7]YZK&.ISV[2R0LeC..
L6Fe&YF#fKW057Cc+AOb;<0Lg1W2&JQROdeWTa@D;VCBTVB2F.(UTO3B0^#S+HP.
R<25>0&M&F?4=FXCDcRZXS:@?Q:^O\5)I\\QNOM3a7P&ZF^DbF<;G7^d<aT3JL-;
T=WX>D\cMS\6J0gC]EcO[[<V\E+Zae22_XdSbS40f&MF5&7/CBA2E[X8NIM^H3[E
:f@GCR3HB5cRJB=[Ud>OG#IcMCJbd\cR>VQ;B<V&7_W&[I.R46I1+Q[L.d5FT0\I
6eRP=5(X+.4D3K#(?eV/4bK+4M2Qc^8US/)&_8)OE9NfQKX,Ze9,da2IP5GdVW(+
KdfIMVFG.&AQ7NHNQ+>c8\2@g\0.8<bT2:KPdS>_CfO&ETNB\J9\G?),7ME0T?GK
WLc0UT]V@=^YZ834CCg1M>gA-Hd4ZfR6JB3)^bgYH&BKK.S<1O;b;e?:VRWZD+G7
&C:?OXMUMHbPRWd=P_642Ie+UAZ/^)35DJ,/(JU.L6dGJ^NPHGP98,M.IH63D(HH
aa8ATT?e+HbB6CBQ1?EVYISdbO-:7\9g5fBQ]Z::_YBf_R+Xc5R\>.dM;5?f:P0+
OcgHKYH:XRU4U9LJfa\a\^J(8^D_WQ\QLP5^^&9F?>CT4H15Hd/A&<1CBXMGgb^X
5d#g/#a+aNbIfPG:]ZWG/NN/<F:UAM_:1f>&/P9:ON^VTC(N#R:RO1[a)<.&<-8@
_:6AP-D9g7,PQd)+DG[CDa3WW(\I)U1,]+\GgL^ZWf[EZ<Q835)NNaKPU1&AA7R)
[;@V)N),KDS1ATfKJ68>BB<D]N7-F&VJI.I/Y-]+AE,27_TLY:?KgTbI50F7,O1.
JfeW;UO89V]d[aF?5J1Z#69Z-3N#WDc[:V7F)0?;^]9f))2JO;Y.e5Ia/@.,3K9D
)0g0gN[9V8,JPHXU8^J/ddNTbT>Uaa;f7b?<5dI:17OL<(abc<-b/Da2CY2/#>e\
Ba;&L/H#b7VKLVee8R>R-:ST:VBaOZ,WL)B5QROaC&4#1JGH?EZ8<.d&AP/aE+dX
S</5@=EQe<8\eMe6QUBA,3;C&ZM6dee1F0^5T]UYM^;L<B:5ZD>-6-WcL/A:B]aI
YR#.f7JbRX7>0+2b.^9\QZQBC3?NT51a,;V:a92P,&V1((T82JHRfcYd&d/bY[R:
72cE87OQZ8#L^EQH+e6A-/.?T+#FZX=0-EQTf<]0ZgIX\;G:LPUB(e)+U,T5^[8g
3c)G)J>?W13/FQ\)BEbWT])N.J8M^4H\aV<.>\I(_:7aOZ#3c<EJ+\a+?IeT\A>K
aSX2^[RKU.>Z9MSAf=;&Jf25UQF&I^3>b(7+,ZZ)W#.HTdY]E52_AFS=b.(U7R,?
)<7@L=A_W<.]NcXI.BF.OIR/W/.^.b>N0,U5aE[M]IZ+H1WE:CG-6=[fC),)_>PX
S&.dIC[JW&SQ?KDBf?#=UU7>bVUFbT&\1>2-?fRfe?SF@OSI-^MUM.865^N96Ce8
]XP5E]?F]g?d:,BHV##F^_FJ..]@I<K<<I87ZH(Ed@G3+2#c1ag3N+a_eYN9?PfC
#5\]^[;g.FdQI;_N)=9J+]Y+:-Z#2Y^;U@18Q_-&,(UFbQ6;B3EPCJF-56WU:IQ5
^2:W/H:;O5)=JIZfBQ:O00EFC:MHNNBT;B_6KSUH(KLSJ1#?F0VQ&+#5^R9&9,@Y
>2QBMLA4/G[dREH@7ZADbPSQ=IA=]gL>G5^JaSWN1g?FX\LVZ1>GN]&#0G42V?9D
421eXU9EeSADWS.<d9ZS[:2@EgCKPP/),SB=E8M?U6aHN^OE6[/OVKBb@:I#4Z>S
P)(&@L\;#39M\G2TgKK937.<SW&:SEIQ3UIR8=?VW]X,\cV@9cdBQ:g2<T+0Y#HS
.WV1\,2-J,7gB0,c^5-DDOYCVO&F7eb,P-U_OA=/DF3^(0afRK3,abLcYK_HEQ)d
<1NQ;3-73?U6R8<U\LXM;YeDCS&>Oa7PQU](BQHO@.HE)fO58YC\JS,S-F1/QC06
b0USR3<UTeT9_ca3C\gb6HdA;Z=7742[V86HBK;AecA;O0b5I,<SfaM=J7gIOb2#
Q?5\0[PUG\18ZL71GV;EJ,eI@@7E\./CN=_X>(XMFMS><F<T3Q-9X#-fG.HGZVC2
)(0?/E4GXFH@]e(YK-=HGfT-7cc9:_fc+ZDKTIA/2B=3GR7R1F0@]]7X,2&N)gXB
1(1KL7JXEZ8UC<NLT8<N^R8J;@=E7O0Q9P^VGR<:.BX]F:/?1LTDT(0SP:)3e3T)
d6CN\aQ]YS/KJ<Ed/BdE2>2^U?KK75fRT][:[1]C)]1CESPN]H]<=8.c7^2CS,3.
7X3U95c(gJ8P6YT8^2?.Y0[598OX:6FE^+7G)=&2b0^V85]/NeI=CYRa<cIHVRG&
Q1aH4d(W2MUEQ3^:@E2>O&=^?<8c(O#&WC9K]DMAY)78]fKA4aL_2JK>Hgc4Q2Xg
I&[20C5=IF/WZV0+(F2ZZ:()9KV-8?1VN^PYI09E,\<JfeLNf>HR\WS7ZF^M=&N/
Mecc?W<R#-C30Q/+5CgfU;&AX/8Z)^RC2fcEFX9L4S-UM[P&+YA2cEN891\aZ^cC
gZe4U@JJV@Ce42cB3ga.J]V(gA>5=-BS8a<NDTB)-=L6G=ea5#0e]K/GXVa?adL;
HFT(QV;IZ\-1W-/445P,fYgb]U57+BX<Q8a\W?/a;:_YLF>MJDU@^#.H#9SS9N2/
-GC4Q7)-W2;fMVf3V:7N&G:/_KKQ)TALTT^cEK9\(?W(^YG4L\R_YbNc@KQ1]??^
U[NBb5;1H=S[+2^J&]TVLX1FCP?SP2fV<5&f[21dS8L4g:X]+UHb:#McE2PI=BOI
=S&-[)Y]CKWTMb5VLKB01G>2/e<#ZAHZVQZ7==JXV:b;LJ_V_gO97N3_8X/5,3NE
TT;Z;8ZQF/@F&R[]GN)-Q=a80EbAP>gM?Ke2[OaR,J^U4b&_#8&,ZU=)_3U0._CJ
Ta.SbD#KM85F&?bP16Je@]d(GK)\6YI8If89BF#cQWaUC\V.bdF_T(cWf@)\9Re5
I=X24MWLM1UE7SFReX\dS7)eS3PMI+1OaWWf(1e1ME9&6@CG[aX7CX9?H>6/L>?S
)#6#L;fHM+NZ/3W/L1CJ3d[eRMdee<,8cZ65UeI;?\JNcO12;,\<g(<\A@IVeV-.
=RWC)@f]88HU84Z?[UcL#X4FB/IP0I4<NASKc?INE>XNVGPPTR1UV.I.,cEH2?H-
342CXAO59P2+W^_RC>VZ+8#SW=_;2)B>/.<EE72&[L;@-bR(]_EB_(H+7(T\[_Ia
4#][9\>(CJ^+d<0>X3B>SX.TSKe#CbdGgXG)/&?GaUQUE+(2c(-_I6@6X<737aXJ
>0<\KI1TQILRIY-a]#cTV?T^63a[cN<TO7:I7L6-.)d2Zf/8(2Jc9/>,I;]M7MI]
)PKJH<Fg52LD)(H4&):GG@RC2(1#6JK/&&QcYQCCQHH^=,S30[]_.N;2TV06A6JS
-S>1#DVQ0ET^XHIB.A4@G^>5MCH&bR;Z?/+#+-+12,e>If6HZ]XZ_?D,e^bTJU)M
VM+]ST(>IaE@GV(?R@K-=3]HP[H3M5ATbc.G:C&=>c===M_GD[:c9L4BVYLCa\]E
Pc-]U0>E\-\_KfO1ISMBL13JMSFY8/Id7(6^[5GW>21,>XB,GP/F:+D8V<Y?PVgd
cBfS5[4Ae1&QX[D-S55(?\dEYZPX]=)7:6?cN<;W,CCUdfHI4O&?Vb/D(a7@V68F
8A\8;UgRSa6_Wc,5Vffb)0/cWGg\UM[DbAN5O8B>eC1CS=E&.@f--RKf=&F+7K&+
;H8Ig[>]1fNeUD2E^A:O3N5.SS<J#dJ]2@dE(\K_WX&1PGS-AfG)SFHXRI/<[5RA
J5)WUa@Ide7/L_P1>(LW2;-8])+5O@XEO?>CAeBU[5RJ]-9F1=?8OZQAcZDI7HUF
RZ_AEbWLR5]@>>.Kg8WY\KNdEDBPP#E6(5=aSf13D3:<AKFD3KSdfdYGP9[A.VQ6
>)0DfaB89@A1KX>fR&+S<GRTIO]=R=5BA54@&_E4N61F[eH-fLJDed?^/LaJ\/.=
@?)PRG<+\.aRg^)^?TKMITTX)CTAS/0c(UL;f=04PN1RJf8@O\D/<S+gQ(<9ZT#K
dQ29(1+^-ITOII>@2#eJ.4^8Pa-MTM=_9&Y03+D,<FgBCZ4\5O4>&2,PDMd?(UC0
7gH2\(^13b[N<VRH-d?KT][AG)\<L<D@(^HEGCENA._Z/E^7KVR_TY43&CGUVQ^F
(_f:1H3O[@a&92LJ6e8Z>f8B)Z6PX/<J4B7(U^PO,([ANX&4K80O2cMfcX]?WH_0
g=WMJ-2\UJ0+P8;;Q7.&7a97+G0@Z1[DU9+>V&/L];<\,E+Y9aB?G,51Z;YDWQ)<
f\A]4[56&e>XCH5S0a_W1-JSI92[H)fSZ#g_XD&4S?H7/>[:c6eT^Q\.VADY.Jf;
HD^F<)/YQ[7)S-6@_YWZfbVEX].6?a<_bZ);PDE:,-ea\9ZR:U8</HT]_-/(X=.?
+&KU>+#@CDU]VVAEHa>4<ZD3S4[_=89/Z:W8GG2eR=64:6dED@L:5>#491N]MT^O
+B],:G3I:I62[)P(6#cd]UYC?OYacCA2\cJK(,PR7SUbcf\H5.6E,LQ,G6Q-E\gR
f#+T]=cM_?3@R[HD\4NHN8P@1cK:&01UWL@MJRX5F-Q?4UBYIRK?>.XB1P:U^#0\
BT:E3RB5X^<gPYS8gGU>?-VbKCB[CT)Hf)E1(fPIE7M0bJ,Df+(_N:[0f.1/59(H
K^2]H<,(&bNZ-O@&);IA2&W1DX:,f&5[bHDb>@V6dA8GP9TREM+GO5>4;\gWBVHR
UQb]F8@=W@&CQW(ZcF.]W8,/-7J4>O)L7YFEb3cT<3cS8S:EJSS)7UIaBC_aaU5\
C7f/E6QJB_ZXPJ7Y_B>g\9)[3)Qd4+E6R\AO1PMGbaN7-KPIe&_G753UI0dD.#(a
]Y)_ZXY78?+c>A3HQ/,5I,GLR1f.=2c16b1.QN.#-:KRM^V:Qe^J.;RUV0E7N(PV
C94+eU<O3]Pa?PY,PA0D[1eHda_[\BJDS::efdRegG=H&cRBb[bTdGeVU&)59;;N
H-&+4O5,d&]eeGKUgV/X-\Ec7H?8MB)HOBgX(c<db17eV#6Mf7XXX0#RfL)eQQ[W
W]K>0II>@=9^K&g6,c>6.IY59U<]afC(,LDL)3:Bg)9)J1b@S-5_28-,38J>0VLJ
G?OS_A8UBf:D,WQ+.C?d7#SR-O4RIQF_4O2W=5.ZY5YN3>&7+E=W7]CN)T.V0/?)
7M33Y@b\&4YZ<\Y]e=89T4/Y7^AC47<GJ3ILe&F<U,NNe6=dMG\eV5Q;WTQ?5)AL
V2=a-KXgOO[GDF9@J.-V[4B>ZZDDKXLS;K20N9J\S.P@[4NBNc?VKNb[JRHC)RR>
Q^7G>Ne^Df]6NZ@NJH)AA#5@1H[9\AQ>N+P\)3<BTdE<9dE(5IS=,W\XUCDf\VLB
>ReS]A[>NbeCcI^/:3)6KLFIJ<:H1eV,1MF4(L<3)gIg_O1O4AX<W[X=Z.?GXBeF
Wb5.c^C^cWeNdL@]gN.M?eQJP1ddS=T/58KgF30BIPg^d7>L+2URNVVHJT#G3JcV
M90QEPeIXWdb.7<Md;ZNH1^e(0R?>8+FJSeW6a6.@LOS_2Y)51TB1Ja-B\4eD8,V
DJKYO;G_^63e#LU^P]@Ab+&Of[<5_XGH@,b587&CC7]-3J.HF43J,,9ZH@W>[TED
/61&;&Wf@:&aXE>^S9?YW?-b(0[#Z:/Q]L8,ZQe7=3BG7=eaR2B:cX>:44</?Ca]
1KHHZJ2_N-Y_c-ZCJ3f7-e&SAI<Y4H1Z7L]Kf5^M42-4?CeMZ_@51&^+6^MQK1?Y
d6[=-,B0HL@OLD6+\;Y]EgMRd_f0+>)<2R,LPFY7E8U59[bG1c#\P.E?XY@G)8_2
,-g9^L5dR&0]=VQ9]79#JTbAE=Q)45be#L/71b,ENE2X<OI=V]=18X2[V4IFSfB4
PM\076V3T#/[c(P3cCHUF]bW#05ee&e@GKHS=P@c5)9&7K-JQ=T[T:AJJ(?c1OU:
;27;6(NH@W4/6C01U644dO+]KaQ:;^a+WCO>/7g(@O^S/NJ73JXSHZSFf5&>I?+.
33+:B5-A/be#C@(]f1K8eE:J#7PcZBB/ZZT^F,OAS+,Z0b\B0U#+<61HOJ3GBODW
B#BN_3c7XV)@R1-=_P&9[)?R6He^F5B64M0EfJ1VG,2Q(a7TA@)_>A=72U0DX.\\
F7;>EHH]9gJCLA@NNOScZC8^f>(LHU)-=.CVF]DIB)#[\73J\<=dAFZH_<bH87QI
;\JOLf1PYRJ-V2G)d.X/(eDeSD8Jc?:dUF[1:bJ22/f#3G@PNNKN?4N7X0/UN\Hg
K>cFW[A8egHWG8Icf^GCTS9=U/6:I,P>T+U7)DeOM,<@g5#/S[,e=5?VNZ=(]U:P
J:F[_1_gSUB_P2KUT5AJJ33?<2L<V;M9-.=d7M<PM00O[704K,_E8:K93<[O?2AI
de(a7XT:dTgKFZ?(a;W7MZ7/f)IID1^,.\Q;WN/S@)8TdQV:T?W[6a=><V\#=T)e
<N,UM)d1YX.D71590_Z)BcGH&9PICXc,)D-ME;^_=TOAF\d6(-I#5C6I6KWQZW/O
_f^,W8Z[JOYVRaCW[b;?:cR-=QP2B-X@ZML5_(2:=?[AQ;FU6)0GMTL5<XJQNRZ-
b4DA..\Xd5Y+[1Jb[H,>([Z8,&_JZCI;C3M?(Wce\B&@B5YCVIT8[8ZB5GD9aNF-
Q2Ce5FO)_A\<#C6^643g(9Y6H[?^X.3<bgM^)D+X(9C[\^\5A6/>f)(FR;XE@XM,
FUK=dRf\GO3L22ceAaBfI)6O\)a;MO\g/^JPRUU<AIC+7e5ZO83IQ7O@#X\SeF-A
GOXU.TSP4Hb&/.RU:JA\\Z7,H)#5ABKK_OXO6+N;<R4D^e/:OObTSMOM_?K&-N;b
<B/cDRYAK5f:)\LegBU99:gRVGX0cAc;V]S?;R7bG4S5c]_:SAbAX2+g9]I5(4EZ
MWK5CdT[)POKVOHfT7E0#D>TbPLaP&YZK2V)TN\e9QDMU/V=J<L1=g9U/3<O5B7J
[C)d(XZN5/f1@6Y][/BDS\&Y1=Nb7RB(f&>ISV&3f\VYI7]9.;6+@+6Q_HQ?XBJI
[5,C2V7TVY[Z.=:aH^e<>BO[Dg^&]E=3eQYC979\LV3,YIG.:6\:)R?AP8DOZEOX
cf]P1,KW][Z]d<_:12B\EA/]G4Yb9SPP1NO=&_YWA/[TX,6M@gdc;T&O]PS]HaFV
.YE_5JYDMOE78K3@W[1:9Qc1D0FG(G8,cdHHG5JG0B_LAKe8D9cA??321=(/H@GY
^7Fcd(TeY\<;R@Y1[Bb?\7>GSGVUAK.JH7V69N9O?63)8LN<MNHK?T)/a7KKSAQL
2a3@;6-_aFW^S+A?F2W(77GW:3A:b=MM]+WVC1N0W@g_W6P^+@NKWX]Z.?)?VBRS
X.]a0?d1\bgQ5Eeg(\SHR?e]2XfK)X7TIYP?/ZIRc+50dT<GNJ(fM@JdV7WX@2bg
5Z=c+@I_VTQ8.MU2/GDZRGEVbd4<Y9#J/DF]VVDXd2G/f3_B8HCg0;Vb:c.I6[eQ
ZF6US?XQL=76:[+O+aU=&=e4..e@0E>&8/9-ZIGfNCJbC>c:5K&B;]&6TV4^&4b[
dTFXF;0VJ3Fa1HBaH[#W2]@;20dFf]792]7b)SA_=FBY@.EPNe[OB42/V^f/@7IL
@7O[ZC4Le\\CJ9BIfK=Z;HLJXcb)>#D\Xfcb&S)J[>K?Qc7F(#YW?5;IRcCO(L77
(NPd+S/FSJ_GgX3f3a:B[;cT_3R#-f9[VWHXFEL#3W0^_fg6cK\U@,V4e.YX/g,2
NL1.^+,RJaOE>]1,(_(@8,3X7&[B]T.VP>JFW?)HA[>gD[Faa:&MMOFcV39._A(d
bX+(+<V35++^:V@^9_G]#IJU7H]a_\2.Y?V.<RV,dW/;A9:I5=>5aMH/=2SA]I;?
9IZII.77&[2FK=R[D/Z\LKOG09VT++1#WQXJW:-W@QX0F4Y@&LDfY2^M42I\_S);
#_&I<5Gg?-)JL-9Jg]g>^(Q7?.F7DWELIOPZRGX\]23eI2E-NT9?PGMMLg.Z;gE.
VGd;5TfCK(@-K9W<EI]?=FdB>B_X>/cWP0:JB0Ee2aZZ_e-eZe#Z[@\3[c^3@+fF
_Z)BJ;I1\N0#cdNHN[-E:dMdG^HVW\aFTQMRX>91NeJJ??YK,eQ2.KV08X>gb8Re
7a>?,]#6f4<c,V)&ELG<B796(,d:Q>HW4G\4NY@6J3,IQL@5.&N#G)]H.8_[&0YJ
OdU9I>fPbTa?8>Sc1T;F0K.6BO:d=H/5WQK.+75R7]WL-;DQ)KN<_B.:=Y3O5/+b
KgBWMA+N3+_;)JbcE@/,AN&2S(NGP>=f40C6,4)-SJ@797(;OIX_eG9^e9DAQ)H8
^:dQ=VRGcf_8LaT[0:ZYGZBT[OK_1#&\84^AP2>L\ScDLcB,JR7-R[BA@#G=T9:?
O1;BeOH;^BO4M_b]O(?A\U^<2^3<];T[L<-@]93<O^(75-:9.NJ>O(\GD-WG^a@0
<JIL2b4]cKM@&TER3g,Y@e7Y=D<C1^bJ]8T1UOL?H^+[.Q-ARM77@Q^GB_Z\=7\[
72O\g0AVY\_aC_b)I2(MX@==af.?<.4G<MMgb)7.?TD)U/.bACcA\D,C\Kc/a;9J
PMcT?R+E].cWSJBSBHeb@<D4(fbgO#S6Y?cG0IOY[0dU#)Iee)2-#-SIb\gB+@3f
#_^[BU4NX[@QEd;RZ#,^2O]Y^X3eL?=&^PDW\)EQE60\5HPE)J1OId&^33AUBY7X
O;9?;PFNQ_EB(QIYDS+1bTYBbD26:2R/#gE#I).67fXI;(P&f?DA8QI#Z-3;:g:4
b(b9V2ZVb-W]Z[de,Zd>Z7?(5=-f&0YNaC;,GdGaF]Vb+J5JLC5MC#R.\21,+g:2
MY<+<3@eVgV;<A5K6e05C[5<0P+?&CW,_W4A4Ne:DPO^O<3:_Y]6=[AMZSZ6F1\g
/3,^7/J2K)U-&&&,:4<L5\eAgcXCbH3^A5CWF+95IQYgUQ9^DYE>-P0fU(I+<JSX
;KHg4,\<#XK7D=9aRI9e+8Y\D^150b23A[QKIa_NN(0-?KQ.df^M[JWQN/)VJXF#
_COH4YRUV\f)BIEdTBY5W8(Z4fcT,I]]SAD<VN@&ZOZ2aM7A^-/G776eZX31JG5b
^7PQ-FE6@HR)JX]Va0N913g/3F#]N+FfX.bF;+gdUf7&1R,K?)2PgA,3#dRNC1QY
G\-1BGQ_=eWSHZa5V5.D8-5,GR2MaV&IE.8(5c,KTEEN?5HEY6PV19J(Y-g.LZg#
8<V42<fZeC_fHZY]6X3eUEM7@a&cV9c<+(E[57[6K-UGY\@KZe-0#TCSE(NgE^(5
<VIgB^bP0Q9:437eZ2_J4:S)E41;M5Y=/O<B4950a(MK8N>NM1c;d;X\8QR.I1Q8
[WF5+b-OHS1.VE9](@]M_QKICd^cSWaLIHGLO.CfReBg/=@YSD&d>0-LW<CG0US:
L7d<H#SeV4ZN1<XSgAP\W12OBY1OPPT/(@3V_-P).fS0-)I7N<)P@XFFC[Fd)8C\
OR&8cgX)3.MT]1MYaRM246C[+7=)5\2Y00.\c\X(KPfHYY_/L[BHcNYFSa#=I,b6
=a-F-b?RK6LDcdM:DN\19D7BB]SN>gKXT;.Z+HTgG.:2e#8dD[O0-JEEdNeI;2g9
@[+JL,Y-K;97>4XaId.P&YdSF6X>5UGP4KF(/VF6ac^#-\2c6^&F2DYBBN5T0B96
eJ.KGD=(cW0@:;<PF2]0L.],3^U0dCW3)ZRRSXT?9.F9<I5f5AOL\4GDS/<ZT8<S
Qcc_Zg#^3;7+0<X+X@ed0NT=ZHbgZ/Y[5(WeX4eLag:4:?R]c@@>cYZOLg4=M]QY
UNXa089X2B>R,=dK4<EHFJg0I:9Q,F6CM:I5FUDR,#]AcZ0/D.07dWP@cVFCcZb)
_cR916e9HC_6Vbf06#E:DYUEX0b&gHINDR]XB-K;J/R/RC=LZ10^BV=PdA591ce[
FV]a_4:4VO6fA_O3.Q7aS8Qgb[eZQ&01.68R-Mf5^^D<Z@_9XI@<#^UQ\bO(+SB&
(UCT[K9c]fR8\2K\]6:?7]751ACIR3bY_QT6TN1QOC_JY-JMeb+_CBB]/09fg[V]
EAeRX[=,0DD9)AbN()JA=CA<gVTGIVcR:QO#139O@+ED:[]E,Q#f5CgLgYE;>Y]d
^2,1-,O;KEdT\Z+E7S[IO:2WVc+N6^=aI/8UOXB0VB:TWc918-N[//E-YRAX=?ee
BQ-U(\NKTa7[#3PI4bfVD-XUGDP4A#&QD&K4f86N56WEg^TfKARS-+#,V0XZO2?1
WfT37YCaBA]0M&ZI>7W\ge-IA_?8#1X4=G&68FQdN?0#:Sd-&:XS^_X<APND?3;Q
<c/WZ+?F?/PIG2@2.2ZL0SeA,+aT<DS:^M[Y&4],7H+:B,5a/2UN41(0)/MYUHcI
a]T8=5C]8;WLPDMUa;),c(/WXA@Cf]Y-d.PQ@RfR]WWb<ND)L+PHC;e3?K+Jb5\:
,\X\M80ZO?4\f7/A()&^F=AU2A-3cYO;F^HYgYf]5eAFU,.QL13:Z#T,R(S?UV(#
0E[fEP1P6RWNEI1W^O(:#ZEd;+\SXOcJ[I?V;RgH>eC].9.45\0LRDTT:L&,)JXa
)fS,?WCISYfVVg._@8aW4L&\HX82/dZ+C@,Za_\DfG?UN7a\E;RS7Z3M=.EE(Be<
W-f_1_]4M3,eS#V/9)6#9)09N[\[W2>8]U0:7TD7M^1<I6XO7TUOb[G-B759&5aR
&)e3MP;8,@ND>6f@U]96c0aM?Cf;#gg8[Z:/FAc.&/VK7QPUK,9=O[Q>9X_P3Nd@
,[N3/EMBQ5OO?R\@8QP9M&15_&BAKFHL3T09b3DV3?CYb>/,W(]]TSF(.W\D/2P)
0a=4YNTb18#O71/-)C)V-VZ4^7gBSFBc4fY6&Y4VgKM59W88/=YU-;(<AT\022YT
e:/g)XU,f:EMQ,ZYWg>#H5KcDI:59]UaSfPfK\@CgFdF:+2A?0Q(Y#EDad\MI#_>
gE:^\gJ[56C(M.2J>Ob3_.BO,FS=Ma2]gW>Oe5,9caM):RM<Sf;8G?65WIXAKO<2
V=9g8Z,J&>P-59)O]YN6_>ARX6Nge=f7NE[4:\/?bgIc,gT9[V89@<I5+GFLJ_Za
/P>VQOJQ\RdVI(B5VSX/6dOdC)PS\50[NEV@28,SSA&@S)>DF4gR^d6J&2LZ2RZg
S_JbCIa_fQ5D,/&S\>-_c3^gQ15Z^R<MQ,80RP4dCb##GJG3McQ+feCe724_50)6
K)0d4X(P=;2R/U(/O^WCMgfdN^1DVdC/XMX&#ZZ:Hb;@R@cQ9WEH9++GScbE?NKB
HGP)?QM\#^>>>c,d3O2STf5c@2UTa^I\_4R4H](9L(04b1GJ=a]8.D]3A[DVVDZV
6.53VJ;GNb56L<PMZJ7Cg/>.4X/]]?RY:@3eV#4+dAR]3=(F:(O>FX3U3?O&QKSS
BR>)_7d0NWTLL\(D,O,HB,3&)Q7Lfd?6^,Z?f4OMOUNcBI49^7AP>A&c;]Lc/LJd
9gb)Y]dQCO_]0[6f,NB1EZLFI0dfZ5VQ2OPT+g4L.WMCdGc<AKf6XF[N\]4Y+AY,
B#@PaB1#8\Hg^;4_PIR7La<=_&3.fB&[4,.+U08d9)T1P,?[6MWP>LYIAReC3^;4
-;@UC2G\QaR6_Y5<N4-2e^[,[./M=L(P5KaK)B^:T4R70cVV,@IU<ca3-E^W:aYa
Rg2_+7J(>A636^RK[e[KWegND;cGN>6F_AL+Q.bZPJPL_06>(N;:279O<6?9[8+.
1<LV[@Fb;DP].Vd.TYFd6HCU.^U(2^#Y23WVNV2MBWLb#8JD1@)g&YW:INTABFPI
HLOGc1H;X=XA\X1?BGNV4I7LU_,^Q>,HO^\KZAca@f8LQ4cNM4E?K:#\f3M@0[1,
331AR5GN]>a+@baV0YU8K=H^>2^NgMT@df^TE2M&)MPF,&2;ZV.,:E.(CISYN2Z&
JN]?Ub\71F7>ZR3Y6<6>79Rd(1L;VP8BccL:26O@GUJ8&)cW]D)<Zg_R^0^F)C6]
?APSK:PW(X9S@Z9/6^WV,^G9+KL8ZSQB-FVc?JOF#.XbKMJ=@>MBgY]W#UF47VQK
)FPfcC=K,^Z97T,K]_@&I43IWPI-I,#g/gF&;TTfVC(Aa4EIa-:)?VUHT?cFCE[8
P[F(=df\/+DJ&^,0c[;^D6>\L0NWL>cg^CT3QYAL37W;.#5)@364\#RD.?)WY)8:
SOH7JOX=4/Q9^MA2]BS;,M/g49OVWDd\^H+3K4F0_e&?&1=@?R1MS=<&L4RVb@HR
<e&VT+QEIBUHKaMQXFEMeZ+<)1e&:3EX,>8CN2;F@B:2a^PSb0POEXPMC0]WSR1a
ADALV&+JV#F)-828H(^R.:d:/)@=S^+7R\e07Y+,_TG>LgbP:Af=b7GQ6LY(<SI1
)VXK_HVeW27J0D#cc4AY/X-D/XXI8d<g1,&Ngg@@5BQ6gK13V&M18&e>O[dbU2Y8
c<JO/&Q<Y>6X_g_[#@(fRCWZadL4f]BcX-1N)&R[&&TDRbVU])6&C^A#QQ4D3-)-
:C;O4)bX(?MdI&[:,]ePJecL:/PB1b\#5BZHD9aNAB/TE+dgR[)52geU]UOaVW.#
525g1T4R:-?YfV?5HCU9<V-3?KWAVNT?64ZST<<=)?IYTXcDP052DfYBe:V07Mg=
YfY_eec3R2UZgeD&R7><P,/L^02S+2Ud+RRS]7GUB<<T1]YIJX3V&R7-QSNYbF&6
&0[^D5XDH^cIg2?I00@gcNV8-gPZKaIAS=/+&]QIZeB(+eFN:8G9fM1_5W-]WFUW
JU8E,C3\:MXMG-C7:U\L9<dXDF@>O3QU[PZN8Qd126CX<51)_?8X90,[2?g8Y\<?
f-93=JM/Xd^#fIY\S+)D@?W3]IDHfC<VK([X=;YTJS@<bW=Af.0;\O09DOXE)<E6
<e63Q&I<@;G_00A(#<b&HZ/_G[>=:F/G945<c;^GH^?ELZZXPEIT>3?B&ZK^2^H7
I>=6T:0,P?e]#SZZAd4WB=4Z&E=6(0W46fZO]KZ?NSD=6]LEa?TIUBcH-E\;g2GU
85MZ9/KFS\XT@CQ4beFQX5RPHC(;K[<VW(@9VBT(#SDT3?:EV=JWd#eeZOWa;>U-
0#S0\83_>3EG&e1S0g5V&4b^[)_:.IB-P?6fXg+G3CCeKV,[E\=XBTFD.MFO/AD.
5.\=#XS2WKB#JWQ8aXW-:VAFJ]Q3I:I&G#+O8>F=1<Ig87:8VWVS][aFX=Y5-1[0
]J/NcL)L@Y)L5>W,8c#68-T>N9OY&]V>gDCU]/gRC/#D5.ZIM)J74<LbaW,J0(2.
5+#5ac&YMX9)B5QfS/DAaF-^N=WAgAD?K>Ba;--&^,K@cEJ(bP,+fKJB?CJ:@EED
):EL28YQ+;#7IH/:3)3\=-Xc>@=gN;aF6VE-?_M6BefQeHF9)+2[L-]Na(JO[a6)
gY_/Y5)S4GdBB<4_]ZV<LbROA6RK<0G4.W83CWV2_5bF;=0,LVSe>?5cSJN]9\J=
EDEeDRcFI?+d#bZABVbYdKHAKY.R1d-/b^7+\H_[d202M[;R_6I-\cE8MgGB?eHR
,PSaU2HO+V,Kc^421X#D&d[)_Ne&GPGQ^PAF63f+6D&N.>B^ZQ^d,YDCNP>ZcKg:
+TYNXXG.S>H39&HJ&_Zg#A^E[eZLB0OV7V9N)PJB>\)/P4U/Xf6aF]cb=Yb0-Vg4
C,V4X?\N80CEVb53Q,YY:N&gVae<)a-TNe#-70]/&1A=8#@eHBF_K180b6>e;R-+
@/KgcbEf_3];fL,)#EVNe?L1DA8W06dbR\?N_9G&6b[G/d-#APGHbK;Mg-dbL[_O
g7XK5+<eG^fI;R/OD.Z9:1M]Eg)=)9/V-EQ8SG7PG#Zc&)9\I=T;ge.0[VH[@R@:
X(^Z9H+0)aGeR-DMY08[&W6UGGYf0]>4RY://1:=0GI^:.+>^8ONO:^S\+8L>/W,
3#ZR#B)Y>78c/4NN\.E=_LS110O:Ff;R;G#N,O1,>g:HJCL38>g-M4?e-)E-7Sc?
24#c\0/]5@fY(L+ON[)\&UX,>O7>(b(GI-;Sd?;DZF,Lb#04;KYS)dC@CQ32;.f8
+X^=4<9U&7+CP7efLde6R(<gH01BSBA)LcE+83Bc66W\C2.LVaT_3g/4,^]7TV>P
J22P+f?G6=47cQNRPNO=2Bcc[F.M:TD.0V+WV]#(,L38XN8M@3g:4JD_(5Q_.(=G
d?#82Q#;/Dfb^4_S)UO#_-Me^N^+TN[F_UEVKB^ZH<(Lb?J-RJ?<eIC0JE&_e=#7
:5X6UH>17e2<1G4I_7dcCG01<_^1@+]7Pdc\O^54S3J?[9@Id=c)J@C14AV.])T5
9IQD(+>BUR0LUR[&3N;NLMOgf/P7G12@&_R->abJg:86Fa.IYS;.P#J+.3-IFLX6
W7QBB-dCbc;2C)TM/<9S1&2Y+aHV6A9+d46XYW6GSR6R,SY72a[g[;0A;^4LDFM+
/BOAHD+.U2Y#^[V5A0[WEUgG:RX#QD.O<UaC^R]3b90@@I\:=F4_T0_g8:LLPO.I
Fc8OYZRN_Y?;OI=c-Bb]2aS\+@LMM6@MI7_cH1TF<8)28:c>4bC:bcLgG-IXCZPW
_B:BO0OMIZgE_\b)B5CMJg)/dC87(J5\IYEga39b3=-:?VbcMCTD-2P?WK28X_.#
Ye9=#5@-<:76V:>CHI#ND8PO_:gQIQT-I2V7UCfGBB8Ja@M-93@e\HR?S6J_YEX)
a2YL]LTeaMV;=QRZX/d.d4f[A0./d\-&aXe0.:<&>:Q@6,Y64<@&Cf<3=Mb_9ECE
H0[,2/I__H6]]N@#_:=G)&LfE?T=3-8e7L\bGLZJQBRQ;V<-V.:_#0D;.>:M3=?5
YdSbQVL>PVH>\A-F6:8VZ]#D^cDe&EA+GZG.9C,\;PAV_IXCG;(\#M[,3N;?_d6(
[?WL8A7eX?O4a5;,I8]W7Jd,,_S0-0?;,#Vf4:[^<&9c()0bO@BHY>ZL=I@8IE:c
::[Y79PU>+bD)(WbBAaXJ\9e4>g7;3<G4E9R7JIQd\-)7:NT3U8(f^4N[]9Wb=84
+5b)0S83U=]bL:H<&Ld5[LK8MOHA?@5[Z?g4^&SFHSMU<4#H[QIDXTR.Ud.YW@GF
A;H)RKN<6T^=g\>9GE]4SMGVQ.QAWAQScX+5?E^Mg2\?#^GF#8;[3:g5Hc@J1+c>
WaEQH9?:E,f69L.e@H;59E:UG7f=9:^EEJa-0b]B9UO2PL]MPFB;[FX.LeU?N_L5
_N2(41T5UKH3I0OSAdW7WA[Y]5K,#b18VF2Ne>[:N3-N0<3,^aCP0A:@-dNS7KPH
L_;Q7C=MM\c_XN.DNXL4OM0=)]V-dT.O1=IAeZ=LBU_cMc5^&BX]5;]DFC/d?CK6
-:fW[6dgedTK]QN_cCRT^CP1G4E@6b/F+Q;@R33,DE;,fGYO@JLBAeKVX0V_@6^J
W#[1I^QFdU-(>f<KEV,LNY]D7I;\aK0O#L3;L+-<BZaKV>Ob.:YWOY&ITP.38GG#
[PWNIa3;3\]RCMX[Ue(0(\,?L/6#2VC9/OJIIHGIH7)J)W@FbT1J-Y23PW1Q^.AG
bHCQgG7.Z]<:BMEU#S[7?YVQTPMSE^BZOY.\^DCF]-]ZI6K>XabCMcEC9;K6WD9^
S\1YU8WPcbQbMPJ&c2b,d>@4R.&f6OV3#UI951R^ICN+g[[2e@FGf[OGH\O=PIAI
XKAOJVNK9Rcgb?b40)EDG4@]4#-FY#H8+&+A)3gQ+7.7_eN\:\@JW](dS/+ADVA@
+c9[);,<W]ZT6&]]]0Ff94#KcI/(e2E8/5#DUB:;Ra@IB60IIg#L2b-W62Uc76R#
Q3QCEQ6#NF5L4WWd&]7.AU?\5P_I(EOJ@e/1^R3_:^(>URf?8WMJ6MV7VXc@P-R;
_+XcB+M(4U9PB3Y^O25g=TMEUU9[fH6(I2aDMN3<)#cUPW58]DSd[V8<B3(f#:WX
N54>N[D,5?X68Q08S;K(KUI]:D/[=gAA<66G&KH)e9WA.^4FF7Y6O,S;AA9G=9HI
E(1b67(cD(TPeZa)6HNd-<e>2))X>T0;5,SA-PCaZ^eaL62IEZ0S)/&+8],82/HF
4<7DIHZ(c\Y]?7FHI<T\VH3.d5@=K+NETQc3C>>L9N5I;aI?H?2GNXdUeQ.IHLX,
5a\S:RO/LC/?5/<5MXZ#]#cL+CPB39TC;CQgQ,e:V(&\e,V#ZAA\_3+,X?]cQ.,B
a)],]I/N6(NU?7W)GC7&:_EYJJ0:SC[,g(U;E)=F1.I88/Q_-2I;[H)\H-ANe&E_
)>2G7SEgeQQ3/1Y6E4295C>(YM91]XHaJfC@4UE^YNTQ=5/AUF?A=F.RQ<_d]3H&
O:;13ABgV4Q,O>STPP,+IM_3QR71P4-7Q.Pcb+4]S6F63fY6,BC&QW<,@P)d3ZP_
Tb2RZ,0OK&f6B1PPA6:&VX&T9cVa-GA.B:Q.\(.R0bVAcH?@eQ,D+4?:4,@c<?.e
C4<JVfR/dH>cJ)aP8[LU,(^>J[J55WJ-87GGeW-/g34:)D2CZRJ[9KK>e?\C25WF
?3OG]\GPa:RMC2\,(_VU@Pea^B,+M3-(CWW+JNAF,\0K7NGN/6ebSLC)KN&VOfXI
<,A.\_]=JEG=88/NBe;JC7Id\_1c:GB:8L1eH+VJJCI6aWC_++2JcK;^.N4?7+VP
ZJ>U&K1J2\P,Y>8KCReQc(/,67VNDfcA2,Da&W&(6&ANg<1^-E7YKdIP6Wf1-,\E
Z<E];KD_ED320-0D&E_^-E\)F[]eN3Z1_M(^+KK5I9cY#S0&aW#32O)@1:<>T>);
U?15L.U,R7_]SS22/KQ8SZ^1K+TKFW,6-U.XJ,H<4H/E?G@UWD9</(#Db-0Y]YS<
CYG\X^C#KL:305D5_&HFLfKC9.X<Y[N2\D?O=X&G7NQRWd8K+WSW:?8Nb#16,=10
3Sc]E\agEBK9FN])LE(edEIJ4eB/;+9RQ@51\6\&8PXSR;^(M+X(NT4CD;C]AECb
TXS^V8T2D>RPECHa8T1Z5TVSSLCg6HfgQYI<2PGD45/]:ZL6-SOFP)aC664<U>:4
;\X>=M9(/_3C\IUS5+dA;<ELDB2dHE4/CMA;35G3DBX?)3:e0Wf\YYQ2YCF1g6eK
\.A&_)9gS[TK]Ua3F0/M[b_KUMW+BUUHf_@WY0)OD[3P<0-[Z_GH3bH7;0TZ/2B2
\NM1]Z;-1><>#HP:YBeH3[J45+1//<Q#.BJ1KHR-9EF=cNCXJfRc7(?\_ZE?A6Mg
a&7e#J@=Gd:BEc;F2PdKT_0OUQ7M1M10#>KO6G?R^/WX8N,LXJ)RF<4.[E?T1PdS
(=-[,))GH&W^IKEFESL&0RX7195d12RI)_F6g>);d:5><g+[&#2<VaUC<<c[^.GR
LF&<7S#L1=+FBX)MB6bWFI[A6(\N.JEF/dS4/##1BR>MWR2R=^b^&8+4_8c+VL_e
g-MRIQAeM\a0-JEWQV;9O9H+D9BU.[Z-f063d+g,(UGSO]^^AXK[SQ,eU4&HAVLI
eU)PV/c;JJPegU;BFcI0TUW&/g<af\J\JJ;DQ)4.6e0/A3afcHV&VIUdX4WN)QE\
1CK2K(6?AdW]O3T#];Q<MN45]BaAL1:>^FWO.JKeJ=B,H4:C@>L9SVP==FZ?W5S-
g]/=L9=^f,Y0eF;]Q;4SJD4>-(75Y5+P_ABTGI7^R^U135<KUR#AN<[J+09A>]8Y
0V^[R-]bS?aCC78c-gS0=-E:fO&1;>6OX4)\=C&93YbBO[YA^3H+1JNA1^aL9EY9
#6B+fKYbb=ER.TF0Z]NZM1C7I[\,;d]>X>KM,24a7_.(W)]S:VN+]?V)QJ,;-J.T
9ESb>QT5EJd:L+.47?Z#0-\9NN+>@\&<:2dcXECKCK4=P+.Qe;g_X0Qc\g/U05@-
V==A6X5?QUeN(b^#C^5@02#T=,#(ST1-I6\LB6,PC8X@<91c7a72-a/3IKSDa0ZK
EL2NBA[YTS#C\Yf?^Dbg;2/ILKOE,Q[IG(e6;V8LQ)FL8G>?]M-@XG1&7bZ2AL<I
ZZX2ORMJ;^=_];&,9d#QTK\=W/R/K^C2WS/3#=+aJ@Q(^=++[Y]U_29Q64>V3Z@8
>US9#F8+\Z=YUgY-\YP5/:4,#SS=;de4M<f2P0IO7;SN1dHFdDD;OH<BfT8JPP?e
b.>HNceKL.fH>RO_5?NGCV9Qe?Y#1.PD3[Q6,A4:AZcU)32UWV/9U0RLWYXMQ\T8
E@;Ag@AZ5KW;JRAN3=.<)eS<;HLTKfX#FMeFUHbTJFcLTS;L75B8-VFP>YJ9&LDe
O/E;EYKNf8,eTS)0;3Y9\6T>_KV2/g)H8RSfZ6AG?;g0d3E>QHd0UXI@U=#Yf=[@
X<),f@HCC))c.)DBG5K])O49ND?A2LD^,KdPffDGW/)?f.Y?.H&O]UTfLe:=(L&>
HHd1Aa)RaG^-N:840=@/\LO12fa^dS,2YV>I_1L4/QDP1g,/TH.AS<544/aV2G6,
;R3>bgSF5?E6d>JQN+&ZaY<eB[<W-W-75,4>[2Q^BX<dL<8.)2V)dGZ95S<?Z/M>
G@aTJ@FVaLNXA/X7+A(J=A(Z-@JW0;ZU(a#@d9KL(1,L&QLW8d0;OWYGF+-UVK=G
dCW.(.X<TL#T=+&+#M,aa;B[(g5[eJ9;I-O/ZTSSM_:Z(AIXO7eWRV]0S04E5PS.
S=-@LL=D+X1Z[RJg87S88e/:YMK&&egC+XY>PGJN[CILDdMU]#=^VUXY?Z)Q]]1@
-,.+2PPXeR6=(MS>cI2gOBA(d1UTF5OM9C6=a(fY:X;/?JZF]45.Q#.0,]<^]ZC<
77F7GA70GPF8Z93H],,X61^7S7IeBVVgPfJJLgc@[N=R?TIBb1D@E2D3<+9XT_7_
DCOB/XL[R#6@YCB[=dQR1;TQ0RLbZ^=VQ1C[24E+/4_3_99\>OLYe@[&FGSVgXN/
\&d;(WaYJUF9T9=+ebR\N+@_F2O1c>CaI+V[60-+9>[b&0^T><>@eeNf\1R8,>AX
X20L05>LOXUa5IWT\W&0+;>)bdL>f,1,(gf5#(LP3\A4cRSg(OP\PITMP>5DB-YK
[>I7EZgK]4M\&daXM&J]cVKc4K62\]?7@Ld7>_(JJ,)b)C?^XZ5KYFO[1)@?H-96
B4gVRF-_6A:05Z8>eR)(W[T4SD3R@[N0=H1bU20280_.3]GdHG(3#dCWZO^42J_e
TE?[@-U9G;HIaKg/>VI7]<S.,8Y5KT+F=ZA6eCfU)N&d];]@g?fE8g=NdGE>+SY<
2+6HTeTOOI+]6BZD4MM60;(Z=CTGPP3O\_,)&=-F.7gfO4>7UCBgFQ3KYF,8)BBb
>M0=#,P[+[1QTS5B.+O,D.8#dN9E18./SJ-7LD0MU#GFZ[<D];gI-:]2L[2MfTEX
SQ>b;NZ0Mg?41F1Z/??]]Za<=;_(7XDP9-M,?5BaQD;MW([G:E6Gc]I\NPPfS<Y0
9F<R_)E(dE1\I-353UR#N#4&>@8W20II@g7N,/8;[S65Ad2^.NECF\a.P666-2dT
7?JTd7?A0N4#W8-REdQ8?8gC\@]dBIL_aC?JJU+787N2\QGQ]],=XN;U&I]G+0TA
[9PE^=3ACfaR\Z2e.&XJddAead557Q[NS9-5_<,(S)_MOFQ0(_-S61=N2G@CL\M[
a?;IK(Sa3/Y[:Vc91f5^\8:d/[()68c1Q[B^VAP.B/Pe&DP\E<X>0GCbOfQ)TNW.
F<KYHK_TWQ[IbbH<^b=JY#-FFK4+1MGNUC^,)T#87#b;OT)J3Q+.ZFU5TR_OW8-[
VdI-C57A,E4f/C:IKH-&4a&8Y[LgH@O=/PV+W@>MMcZ[_T;ML<KLC.K)DHc(<E@f
7R#J>Z_;\X=A:H](g?7[MLaQU>9,adCM]#O?Z/4RIU<Q5<I(5CG0R\0aNfHBf9RB
ZH+TU8Q<9S0A,RG+/fHe_.XC8Q,LTFV-3P;HeN&PJ]ef5^:9O)[FCfEKVJEW(ff7
J]3R//4A2<?bZSa>4=,B)0P/>Y0]8J@cACe)[,cF@FX]aRYQI9J1R.+TI+:==a.W
#&]CCN\QQPY,0&T.Ff?a3HMV>1PK87UHD360R<,INP\G)/Y@MH^IJA(Ee:\KeP;.
R67_4EMB6K?L0RIS=T?8LLC^_E+CCHQ8>K[/LEG,61.<cEK6[1&a:IT]GRMMM.U/
bG<YT&4]\f618JMQKc21K^J1#;&DbdIg/6dPS8<E0:AH#?dg]U.Wb>L[113c+N)@
Z?R/:X/?O(_#J__:D9?<#Ba)91I/=XU_I6HCB5eS]RZFa\AM,1b5P0IKO?F@YIGX
Nd^Q5]VCKQ<.?LB-Bb?(Y(^<2=3-VC?6\3G0f7;>.@ddY7;LMga[OTX=6T:)0G7/
faR#SMbYb9CZJ99@)ZX?-IVL7IHDYNW]U5]V/eY?#TbeUgWDD\=eM2,8Cg]-T;;F
L(PLW.IQTe7,1=/eP]MD918SS&EP&TL;0.+^dTP6#R2#XAa-ZAYCHMPM>BFfff:9
7/J0;Z]ZSJbO4OI)VWWe1<Rg0>_I/4JH,b/]1UV&=I&daO\#f?YJ,>Wd9QDIgC9U
B0[gX//<F)PaNfZ[b/#_]IZV,;6dOeb>.+)GWD=::c&3ZCOCSNK5K+7?cS29]a6;
\OTK8@RPY11a3[X&a16WcPBV33CE+^=2\d=@9;ZE?Xc[2cbN(\AE6]C4^Y>+-P>]
9H1D4SIIY?@g&.Ofb(HTW6.c/\E/^+T)O#Qb,.TUd5H_GB^JR;N++562d4d/OfgZ
Z@b1CT6c?.0YH=FX1IH.59#G]Y6Ed.5?<?#E@/9[,4YFgOa@_:EP2E#3Cb_fB^dZ
&X-]<O?/eGEJ.AdIF/.\@^4Q6c-J\.5a5>P\GNe\1A_Y0>M7D,JN3B\2PD/+W/LN
TU[O]&.:C_Hc&dIMAKCXG\OL;#UY98]ce/8I.IK,(f;CVbF_E03BIZ=[<((KDHE?
9eBPG_VLQ?ZaZ;^^)8@P,]TMCO/TCWYIH>>5Y?Cd?WZ2<6JD?TZ]?8Z2Z.e7\Y3E
[W-d4+7cKB0-)E8V623/cF>7P1J1_K>=d:a0-_HQFE,6gPNX;]EeT#-@HJDgADC?
\PF_D?:OP^eE5Yc#Y9^^U1R?I)9(Ob_L6/UC=&E\5bg<U3:7?.PUdW=]X5VBf.S-
g9RFVafAZYUK5O(=DJfB(Y6d\7^^OgIRWT+(I]+gXbP,ce)B;Ze2-XVK0KCM_RK)
3JI?YacdA45U8:#0WV>R<U6cSX5aBRCT4Uf3Hc;6PH1\U8>[>8FM[)^A&(fRXRY\
)X#-ac)WA96DgdLDf\FgL2NNRWCAHFOZ?2Gf?0QdJ\4V9\UJ\-MBF+YBcDE3LX@(
GD;7?W]<RXE_H<P^?GHbQO96Q^^PDRGc>gW(=TeA61cR4[Q1.G9U#ABNb0OMKO55
<TI,=CET_>bE\Q]AbLf1SCeKOK=L5DZ16G@C0)Q3;TQ,dDIBUf7=RQN0NbcB#W[7
?IaB;FIUgRKCD1Y(04F+D0fC(-,RA<UQH@,GP;VIQe(-g9/X#E6&^DZ2O6a+XUF^
WKK9BZ:95WL@fYFF.<Z8,Z]dRd5VaeE7.6H<AL13Q00+^@g?ecC)--c^@SGBS,YH
TQVPO5L^9f-FT-849^M2KCVC&7Z@1MYZS)CaY5,g_Y+&d/0e)]_/P.A(O\VK<:KI
J0f.PX8I,)+e:Y;4+&NO(?G2e\>bY/GPDKTdK5W&Z-a^&T,<6C3bL-]];].b,R6U
O2dPaR@C;Fdb:2+d\5gHWMI<,g>bDIV&?/USZ<a7e_2gUP[X[>B+?(;:U0[Ddg8=
K1d9X\TVZKAT@>0c2QJ_-\M&/^C.OaL?OAZ6dR<.g0Z&1dad7Z1T[^LTT4)H,4=X
c+5K=>B#20=OZ_>:[<:a2K64=,5FSPG+0>J04S7YW625I4=_Xd</C42UPW)C]:aR
,PP(8.B<0(6BU^#/A,Jf28[OM^IIN(1X?GH0<J2^@,M.BG7^;=.P=RUIW0g:/V.1
^+=_D6:GH+9Gf92=>OUKO8M?:MAR<=LTX_R&a(&;6JMLVFUB@:;R+[H<6C8=8FQ[
(9LL<\\LbD45CS59;C:cU6O5APCS4I2BL.7LcHWX;Ne/@<./=3@PXODFMRV3NgT_
VUGJE?\&?McbY9SC\WS4-;>M..#9Q,5R_N+-4PPa[[4RUdAY2),\IQ]433453;YS
JgG<&8&T;V-^(5g_BQ=2.COW9#g(T+B\f&][S.;>0GF=]R<#O<GM.^2<\UO@+?VQ
<L@OFRUDMUUSN[2XNM;NYC[Lf,e,cAK<Jf]NCFbHU>IS>CJ6RT_V7RU)F,WH(-d>
gNE^<DWI:/e]IFPOXR-fP/K+UW\EXcAICW0aeTUVc</:f:0;<cQ7QGK/XfPQ3KDa
5/BS?A+0?/.X=P=3/aZ<2+c&^CSI#)W\:@cG#]H6FY-9TO6BP8a.aW5#XReLfT)V
B.:,KH1-OX>]T#W5,VNfT3D9R9)g4aW4.),bAHNC.G19I-GNIAEKV3D]JAe/BBOE
7QCMWPdY).)EgGTBS#Ed>bX8(eE8?]R0YPK<Z,URNT>S97aQ)#IK(O)MT/a.(KPG
GFgML^JPJ^d=\0<YC9>SAHAL<:^>.\b\W9)OeCbT:DK5#=JGXZ^LHXLZdE)8DTf+
PB;<1OedL&(-,R/SOcOeWJ5b/OgeaLHY=^DC^5?4W;gAQ\;UP=\6+OM2Aaa&I6I:
#MSaVZAZa.YSA.bNN+]+PI[R>#;d0Ua\3[&1e_RU:)TT#C-[+__b.:Y+.Z6a<YP=
8(D=Y\Q(aGLR00)I_YA\H:G>OIV0K70<^&U4Q&.UbD\F]X;f&[e/B.d8(Y)<KD=M
AJSC4Q+LKS[FR#1^dcUVa8Mc+VRO]R^g\B(8OY9\NLO:F(]Q\9ML0gX.Ve5Z,eG#
L)CM2Z^TIG&(Y&bPQ0U1?9F6&WT6\7^^D>58K0,O[Q:H3PTL)g)0W-I.6M\DA=7A
[,.g07UN=\f).)MU<8?A>:9Lg\H5:>U?/d8J=AKGc6^5IA.J#\K=[Kc#fXZ;6b)]
UHAB?FM?;6>dDY/>7:F3&egggOBJ+.2,6#I,bSB_-6O5CfM]Y9[?f=<]KKW_^K^1
c?D?1EDI]Q@AI;-NAO7eXH0)+Q.4FXEB,10>L^GA1\B=)8XcT\>[DGIG]8UYAQA5
EYV]+<9cE71S?1dEA:FZ]8:PUb6K]3_cFBXO32OXgVN;GS_T#2GJB0GH3CgQU7R.
@@T>H;KTK?8b5LO-Q4P9.P:aNgV<PfA7eJ@>F?Hb\7RP@T(&P(g^2EZLILGAaY4/
QfeLBB1\UXO3gHgcKA?KH<?fJNR0MR[7@aUF<P45^9)SMXWbPPI0MLU:IN34XJXV
#&=BO3bdbf>cKED3J-:98e;ad;:^E(+eQd&,JD/R8GUOG9-@\-JQ<6_4dZZDHc1M
+CE?LB6SE)aAHd.1E2P]()80:CT_J&&Y+GM<b_7&2?9XbK9AT[TGQ&Z(7P_H\2&T
YH,:P7JAgB_dZTI>[[DCA.KL<QZ920,TA,ZJ9_ML]WGH@B)JE@J1MbcB&_3MJDKT
KIN:#IFURDQ9b0c<>Bd.6MO1YVP)O;GW^16HKF,;J0=[+H]<WC7+L/[34I1[S6Q1
eaaM=2_N6:5,e4[_O]0THLG2];^&BKcX\]^f614GL[0c,/:.?ON]d40E;N8=D,KQ
]YCGY3bQYf._#MeGg;#@PFQ50A3:KEBD2b?<HO_->7cV;/(dQOg[7P;4-4/).:IK
IUUS9[ZO&R/+Q_,9W0\52]0J^D\6SL,RKd8JVMIQ#]X1S&RDP]0dPFaJV@dQ=R3)
9JWWdJ2@JaTP,4@.O?:\8.0/CL@:c=gZ6K13<<Qe9NfVP67e@.e/-&3.5)-d4IcH
.eQ23+cYd((6#BZR]9[GAF@4YaPe55eWR+)#HXe4#43EC?-8-4ag::<2LL&Oc#F=
eE+L7VdN+R]#Pa4WdSca9W(JMW7-C^_cYe\F9/3\DE<c-YZPa,1Y+VVf7LgCc.J0
_<K2JVGD:c)5\0FUS?FS87_U9>)1TT;R&O?aYa0R8ORM+@\)Y3(VL/\](4S(,1Y,
XeKTCGXaS])#69(TG.LHG-V+,9ZQFcSfg6DD)IA09F#,I9UX&;]A[/6#I:[I5#?<
XNcN4(0.UIWWMRI99RNY.,_6Ie.H7b;:9B-5+=-dC5^eF85ADDa+FRDFd40]Fb:W
\b5AAb=?^OO-YJG]B:b,6N:;FJ<\E.VdL&[_XUD8LBKbf4\FB/>C#.9OL;5KY:QD
0A?a=B+?dD&Mb]2SA1(Q^-:gUSK(2B&?U#HE@>9U>&:]<6#MRY_/2=ZU+fIWbM78
;d(a2dN/TI/-RN-A5]=#:e.7TYI?QT2@K-N<?UR8WC_.:U:gg^WC0bG=T_9/Q&MF
..B^?@A[A8TaKW#-Ef2aICC46MM=RJLd7[5,/dZX4gJAg)6RRcBgM?^X@W]D4:<L
Y=KH.W7.,.0>J.\3.g^#e27:UMLLR,PZ<[;2938.QKB1+-@Z8./L@:<=V/5\NS)8
SS7cUYc2d/9I_^AYYO]BLEY>LEN46S_&B.F0TS7+;&JJ^&);S^IKfS0;T<Vf6G@0
#0dXb+Q+KTZ^N84LY(@A#1f]2WX6<ROPWIeST&E,FHA2@6&]Y5=2HE)X8Z:7S5JR
c64=6cTB2C7S)[Q98d..8F<U3&<bYdKgg^MD@E,g.Fd52PfVAIWU1)PM;1I8=8YU
K^M62e5He^fW/a7D6,I3TGcR\]]76e:A^-]0K<Q]M@)Eg66K^19H_4QEN&.)272S
eJFCGQBZZ<ESdcKB8<5S2+V4F2U0]J+[E@-(UN0fN;]?DD,^S1b()f>EI;HRV):-
[U\EA<](>5FAA^YGW]WF8/#5PgddRE@#GeM]R3&28:FK2P5?[#R2/#GG^)4S:4PT
D3Z2G@]IefB6R#\PVTIbWJH/EcS)bOIQ7]R-aIEV&Q22e.Q303Z68GLPaV6&5=]T
7(RHKSbGgZbJ3_L.+dIe4g7PF[05Xg&U+@4S6//N)V-Y^G75RO6<U,:T4W(b3>@X
CQE/7M]/4+4cW?2;?9N)946U@a1QUS53R&))[);&/a7#V&[:IAE#6DOX)<:,,9QU
J?1ZeC2>QJ)ZC/gE2VKC]U5;VD97F=_DNX7OMJfT3SF.WIHdMbFT+7O<CHg#dUXd
#?(5MU4(C)-@(>YERT06H.E<7Td]=(2-KbbW6QFJ33/;2F@7A7IX2\b\]S7_M.gT
D;(@J>H53,a(\5]Sab?O.9EI9SG8DdZYa;b<TEQ&AfIC:6dA;<ZfBU1;JMA4CbFL
;>]\CZM(41&KKcfGSb;.M3SQK;F];XZ&SW&-5HOIC+.>HP:^e=ELL#3A;2L3bR9P
.[@/SfNN^JY3]?SCY5^A:EQ)>\L9^a7T6CAXf85Q:;=3;BI.S&dDg[BN8f3^-gAc
9>UW\-]91F8)&A>H^#8?BJ9.4^WQ?J]+Q@05Mc4)K<f;eBH@bPb<J_41=\\g9D8J
K4gNUgAC+E_VdAV#R.?A@&_J1Q+7cf++PDbZ9;c1FI\<1Bbce?bVV[\e0-<B>UEA
]B(0\^+&c9BQ0IF?@,?--gCa^W=R.:RYTP_W=:K,CDS.79^I,Z8)Pa=adT/R=M\[
JH7GG^>TA>.9M0f4)A:D;a<4dHZQQaJ,/(GGO3-1C@aHX9PRB]IMd/QPfXS6W:9[
CCWP8cY<,a0E&^e0/@ZNT5P#cI>3f?ZWG>2JJ/ZFU4I4?YRIf5f_@-2A8]Va>ATS
/<NX_>[#,A)1HW(7f[Ud1fOUV<IQe[a@\9OcE0TO+W4dFIc(3LDG>5B>,]XS37R;
K:]UB<^4a4;O)WPSNR#^.8FP.SJ0S9&@;R6L0TW[bBCfCJ.+D:A&<KHL0e1X/HNP
JG+KUfY7=;;)Z5-U=JagS7aMS1YgO]M@5P9GbLYQ#0PW-YH3O/DUJAT3aP+9417=
>>6VgJ(?6@;WWg\FB9JS?\HTfED;,]EBMF@9JV&.ICE_fVE=C<[Y;0T+X53E?4\W
Pg7A]2NS&b3.5)9fTIJC)F\\&)J8B1JH,XCCT\+@0I^)c1&8LRM[b>Y#&81_6PMe
[bO^PX@eP4NYWFL)K>M43PP6bIQ6#&Dd/N>QWFJ,@4?MY.1f&DZ?B,]I,&&TUJR2
e??D.Z[>CD@/0e3:F\]Ub2F.fUK5e/(S:aHVDR.P3L:BDDP<^8R8]LCCcbg,5\e]
S1(P\VYYXY(4PXGaH0P0T_)4(S-?)(@UOZ=;Ga]J,FEdDPHJV-7)Tb;]Q6?b4>D1
><8(I&?RS7TRHL\:9K,MeB62GKba3fLCUPD&;,eF@9S/:-H>gW-#Eb\KGW:<-?-,
\O:0<\I^]Q-E?K:SSF8SLR/dRTD&Yg0D29>a=D\#T.gA.S.,aSIU&XZ-\\#J2HdW
FY/DB^S>ON+N5DYQ4f(I@03J](EDg[7NIS^M+QVK+8V\=)8))0?S#UQ(G?/e?OdW
S@W+eEa659RcDN=5P=79>D_9\gbeZJJEaEW_dL6dX<>KA##ZE4&HfVBC#N,fW=_0
4?Q=4566JaI\C8.=Y84H2HBF4&[-=)6-.(0<d[&0A+3)8C\X8PT7GC8-a/AB]dV-
ac58&/7=XCT&FKb4>V]<3M^a9PGS?SRG?A,X3+2X?Q-KP7XC7&PM3C&PENM^=Q0L
2\dBbZ?b097efg@CR1&VN/WbRGTO3fDL>QA@JR&e@)X)GU@+Q3C9FWU)60?NRS=(
FAdV?68.]Z#A.@SM+R_.L_JMRSOedBDLZNRJ)WGOZC7KZ8Q:3&\e-d&K.gX^JbL2
W_O>Lg=AQO&,e;6>HS\SbNa#W)3I.,.P(/>c7,W>3SDXO8:SDgfge)/:3.L^6T,J
C//efTX@9W=9EVC39KE&DNDFU=3bY>f?U,dY5>J.)Off1c.5KLW=1=bIY-4+Y989
HI[eO7/AZ<<PF+YEJGKe;W#:;FO7YS+S\48gQ[F@Jb,+dBJP\8()B5&:G&R.8HK.
XL=#aF[Kg]bK98667dM+T]:3B6<P6XS440=MO6M)JNVW\\.;-GdELfVFMY1g2ZJ_
@^)6K)11Nce25,NDYL1N7Nb5[MHY&IJYfUO+M[O,Q40UdO5Gbf4Lb:;6XgUJN9U;
a.TH267&T5MJEZQZP;?LB:\CWP#6;;(Q+bT(XNGH@+>#G7.O\,dKg9gRE(YC>2Fa
/2.ED^6M6c+L7W65Y_FRVRA;_YUc--cB@,Aa6A8aB^:_)FU0Vae#2UdXSO&A[IQ<
&.7[SF>=7#GB[IaQE=_:Y7,dM0S751[S9Y_\T?SCNZ+J]+_Q;G+Z035g:GS\/[aW
=K9=O,Q9IXa@:__4Df:QVEbIRV>DKfN+>PcFSdCeFM#RAG@LO3JSB-YAH63[89g@
b#9AF&/S+<L5=2:c:5a[:]65QIUH3_NHIY1)I1M4)W.M:>a9-U,[2P[,b:8964WY
8f;Ga<WW.<\9CFSQ:g]IC]F\JK,/B+)B3eK-8Qa4&R+QK^<?&8XEZ]>JI@G?dPT+
Q>KWb66[RY7R/?_DY64-N#Qd<?7ULT\]07I6f?S.R7>AFHM<D2#Y/:Z7E^L84K2Z
(KQ#)dZVIYDS9M,0>5TBAVS_c(6.LTU3I22PN9gD7XTW7C#&fdF5ca/D:,g]fMK:
ACYg,,D06@F9ce:2&GBJ8P-C50)4+,ULMcYHd#05a;J5RRA5F&8Y6X;4(NS-eW&^
AD+bO-O0Y]/G:X5.&eV4>2729d@=,K];6F_RQP3_OF(9V:M0;U;E^#Tf\-fG0aN7
gC[a3VYR((@4]S#B/)b-f3?R/eG;_aG4,07?S,9-T3Q&g5;\(]?aB3:HF]:NfM4@
(N))31L;K@_O,cZNdBC4H/IL).^[3#DGc>M(#\BcI1^^:>bACDU,;Ff<c^e)7>dS
?P4CHR^bZ/UBI:@X2\d;bG[LBOWc]c<)H^)D0]F1BX:>5g/]9UZa2[5@XfbG0>[S
^;&UX]C1]&TW==KJ:IHB/D@X+aMBd6;N=>O(63N0#]7]2Z>X>4DQc?-gHSKN8JGR
MHZ9d+?C:;)JQC?[T#Z\I7gN#G\9Y:Z=a,VOP?OPHQFB4MFc\5ZAR49eN>0_BATS
7a:>J-91H<PG91QOB^-[\XAZW&VPF4=]D^T/TD;HT:C(V6AbQF13+56^39eWc;6(
5_KZKgBMGEPSF:TC9M_FJIdC_:Y=5Hb#gYL?-HeAR&>169(M3gG1(0[Q0GcE=NNN
47&#)MEDEI?Fa@,0KB6D>(5III+8(5dIbR\ORa9=<7(d:6:IU.2LG/8PeVLQ]3:Q
HeK>AQ2d13SVGEBD[;/&913A;Yc1A&f05>ed]2&3#]B9,[e7@D;C.(f7edQ@.e\#
f9JJf+)NT9?1Q(Y::)_1R;GP+5Y;O4E+ZCb4J2,-f\7EP=Yb<P=1F-CD)4IHGB?W
#_J(dg2((?1bT2^FAKb,_E0DU,9]0[5c:]<2YPC[5U_HJ.0)&PGd\+1fMBX-.d(M
Y4FSNIJIU3SX)aXQQcFO=bUfW?0T1<O>K?M)8FbfMb5].,HKPcQfJHSPKW5GI;]Y
T;2T9@WS;)CWZ.:;_fHN)V6X4066#e=LCO5-G.=DgB1XU+,g=^C;C70Z8QPSN8\\
E5g(MEL9EPCOA>H#Q6bR@=JgF&eb>EX>:U_W5+:dZ9d+Y<K,[[f[=U\732G6BSF?
Vd^UbX(_57a;;CSXZa(a9gf<2dVLJ1>2RM4?ST46O>DT:gBPc&?\Uc&(PZDWgKFV
ZER0I:CE<NTa&=4<M=4:_)CVHbd<Z,g>MIU;38=8;-256V./g\c0[T;C&36^UW1S
Pa_MTPfc\&+;6f;<Wf;<81TSB\edf65RFL<H<<aM\U7,A-e5Q:7-UX(VVMgJfAYI
]M,[gOL)F?0@BK);9:5C/YMUQdFTS4[g9VeVQ6XSV0-#8FAPX#Wf\_e@;SK#Wg;V
#ZW/a\gU9eb/UA:VFEIUNN_M7T6afOaD=<+_K@V7b@1(W&KJV.P8@F6F@_SIg#Ke
3O\OLBg+[WW\MP9Z)aGS<cPQ9GB#8AWKITK,#;1?R4DAaCE/AK)g/+L&4aE8fJ\2
Ka+9=bb[AV6AcN/g_ODG]N56_f8aGCeM.Y^Gea^ZV/M@J=_\.HgIa&VHG31(7A8(
Lb?=ecDd/.2K?NP@IWIWUPQ/V>N@T+LM85E6-55FA,V]QCUO6:\T=Q1CdH48bb18
4GCDQWT_BOcO29[OB5=38?#+@g3:R@eKKdL]:e\ZFd=Ob_9K2W>G4A[aaYA6D[V8
@c:3>bE1+BWf\aB6^&<JQ:-UO\Y1UNf@:/+R7S8).7MScRW)_2:<gdSaQ;#19WEX
DONYLWV^Xe(\NRV23]VYTZOL;D:+<4=c]c]A4JI8TD)SLPL/@QPU0DL7@F)R5TeM
95,@/)5W6J5H;\a(BVeXEK6WK&S?1T5V.(d)YB+YaHZ+953a[P<c;BNMRHPU#U=T
TBU3(/KLEDf;>6ZL2)6AeAf4<KWJ[UfS;+VQ[AVX5>1[H9C+TNWVDbELB1(&(EJ(
;[.a[R&?5E+bg54(+6N779OI(2UXX_#PcD(J+/\V^:@CaWHHRIBD1T-NE>E#QSN@
B\7#7/2AO-M>B&R)HBD0-@Uc8S.:PQ&]PXA3=2R)bT>-bGZ8eY+-(e;N.9@4.[+0
e8^Pa&R[bb)VLSReCd+L5/0+7II.a)1(fF5@9d#=G#/82Ld2^7ZSN#)996LF=G(g
5ZKaf2LHH\8ICXU(\?=UU.UCcMEJ<XWI#<b+Y?g/<b>19b[,L#4Z\NC2I7JS8g8N
_\_g0?:P3:N,AB1J@4(ISE:_P_a?FI<DNd1?FDdRJMaf(bHC(&EIVXT?b^b4c3JC
cBM(FfD-6<3:OLcVMPPX>19<#Z?bF@e@@__T0DMM.d>+aRTEf_]QAO<()Q>XdE&M
\]/\b_W9ZJ@O)<9Id1/QRTeI<=9ZRgUH0JO;d&^<9U=AE0D@BJ[<53L]e1c)=EN^
LIa>g,@XQ<CfB;JUM-I.DJV.H+(#>b]44bVGZCLgW^c#MYZY#c3:&.+7R/\=MOYe
&V6f((AO3;aN=ZTg-;d6H52f&fO)QTfU9T#@4,?&OVYYCJ9_?;IXLRD?VdSU(Qab
HGZ#YFC:09N3OUa&6NcFbfAI::[4S[S=-F9JDJT#,>]Z?1MDOgAKa-N2_=Ob2V]N
+9#NddP-<E:&,\eIYL[]DECTPdO>9]O6KeD>fSG1b]U<,9XTLZ0fY[a;2?b.dXR8
)VcbOO.)VITDaU3C@6A8/@/1P_&c+MB>XK<ZJ[=_&VQG.ZfE_Y9NU5<4.O(fBDKB
L:eK77E;=)4XEUF[&(b)\T<g;4F[TZcM^:f,<JL<\G8FSL,WMAc^N.U7/ID22MV?
#UU5.2),R#VME/J:FXBPe\&Ueg4N-.-g4]]V8S=HH]1#E-0f2dT5:X)gAeJc;3aQ
O/RV/EP)+N;RfFQbPE_IS&LBE+VK>b;S3AZC3AT5b,40886;I+,P7@MR8GQZJB;T
=LC,_&94,b,&FLHH\aQ0)\(b+7NF#;IE<&12T)6(QK#5;])8N4fA8XIeI>4NJeC,
R57d:(&=XPPPX3DAKLV54?2@QScae:/^d3J/HWJ2EO57>A>b.^<Y.9P?ZY>QSU/H
CWGQ>B)9VYfd@S+6@\OPcd1MG(LA&MdK3?09=GZG7B]#J1RJM(R(W-?K7HX?-1,]
L#8T>HYH(VCWS=T\\J]:J[U,F9A+[V.U=H,(>KB[g@U.3[O&e#&c^9;G^,TP+++P
A+Q2G>QD^fQ>-/?I,T<:A[ZQ#45J0(VL^af=L?YEdNKQYeKPa,I;Xc6G9;5;e2-I
]@?6O8B)1_8U#=OE:X)V/bOQT_.O;>:CXH-75BISRET(/bT\=UBcI>#ZW#4:7>0V
IWb^=+^@V;FJVFZV961_TDAHSe)7HS<fXSEAC;,3ddQK&E7C@7=ILFM1BR98aG6Y
@=/8d;5.fUS],XV_D]33/DdAge_\JG&G5ZK64B46=&H1?79@\U8I?P@FHfR161bW
>&3I+8I45?e8IW7L9(P(TIN1.80]OWJ=\:.\\XIK<H?G_#R]DSBd5P,c,0@X+O<O
JOJ6b[abS7Ke5^]OEgcUfceCOZ#X]-Sg7OfHbV>U@P,P=Q85J3CKR-fDFbG5IRI.
+E;+/OU?f(>f4g2#@Z+ZT>6b/BYcZeD7eYW159XA9a3DJ?@GPOU^LUD8&c@E3/LJ
H:OJ3L>QC[6^-6GJ36=X.)9[PGVXaW<T2V_)5ege;E@D)c5X<E.?Z@@F;Y2&dB=#
XF\H&Wd>E#U_1-e&YD_f>;DbU^_9DS(77,?gZbT&R[0.EZBERb0XUdQVaK;fd[]U
OeR5gVD;/A5MFZ\f?.ITI/QfC4&2>#668COXTd+,6IgIYe,S6:K_6G&#cO3DET:C
3^b^C4V020;/1GV.7:4]]OTY=)aAFI.TI-[<N3fOY41gM(@Nbc30Z/IN.E?T;Zfg
?<-2eV0dM_KXPa?\_6gKe@KS(U0/,XbG4edWW.YS57-+FH1[,,+QQ96)?4SR;DN6
IM+L1A&/FMHGbg4b?KP4V^&=WZ<ZV:dUWf=W/?W)FZXP/H^73.@34>,W2<0(-FbN
^4U<AfO>;+B-]P_P?LJJf7I#A(Ib6K#[ZG-EYRG]BOf5Y,?-<[M,W.9\.FTD.;(b
C8\XG_U-&?/_-D2)BCM/4L@(#3:bN<Eg#\XK];XgYMY8O&MCE442@O7<W<Y;69H<
&?-]f)Hf#4RE^C;27W^9<DSJ>HICUXFO=P;/2VLXY_HGYQgK[)G3QN/4^]Q[&gI<
Y(g5_;Oc1YJAaYDN-?J]YS<?P=.2EHgFM2S:<@_=IdB]F?1S9WH7K6JKQMQgPJ.F
^M-I:dcI\I)L3PJ3f.96TAOZO^PV=5Q-OE9SJ8_91R764_O4@>+4@B+d547Z4Vb&
8PU(D4]KZ3NDFLg6)A?B<--#2U<T:IJL?PcKV7>OZ#<)649=PX<M0&GLL:&IJ-E0
?[X=(W0^(KWNE^7dJO?K@X/JIF<HR7_ceWbadUa):bG?f@B@a..b0Lc?@F&Z;P-S
LCWf\6[0+2[IFe1+BZc#c+:@F<YH;e^/<9>E23;CbA[)X,]=PS8(=^P0A\<H(HJL
@S9)AA.Ib;F?M-/:JTRGD[@9S\?=&_ad,J#0(E.BEAeVKXeAOb]C9c^GJ25;C:+)
N:5FNO_J6gQ[2Z[5S)ZB9_5,E9P5SU>O+Ia;6,JDLVSQ>WZW(PLdL/48H55MR7F>
<R#Md(_M54^8RNbF3,aHfFJd#PdHaHBC>(819;;V9)XWe2@Kg)FYaO\QQV]WNQBT
O<3001[.37\RZ/-)V>=[d(VOP:UVF8D]NZ(WPgW@0^6_Lg2We>+UEGIaNaX,(,YP
8[C\7?)XW>E<V/SM>>?@#bIC+g56cP-Jd,LLA\,7VU_R6I?GZQ)6\9I4X+.Xa7.Q
\F[Wb_]?]M-X9OW5A=WC3+QNVYKI8X)dM)WgHAB#]:8\/J\^>@>,XC6Z_bO[??;]
bW&)Z6?,#TX=Y-&KCCL:V&La5[EJFc2.LX?)T#QEG;(]Rdg:G#]@:e](cTTC@=;F
KUEY?L&#8DV2H\7[DWAIKCEY)5=b=2=QKWJ]2&;SW-H?@FX34R&XfeX0Qc]-36Nc
VPCC+6bN)<DV2KJ:,K]XYBB[C9e]ALFW\HVYc+10=&_1Wd,<d36T>.IY0M4T&?4P
,51;#8GE1D3+DY7>+)WN_U;F0RJ\<7b[WV1WH#SYET84]@^WDRda;,IQc1V[;YIZ
2:6VGaC^I0KbaaeNU4Z6G.&K/A]VVV7YXM9L/1-^A[[XYE6V#9;&dH++QK-L6\9/
J9)2JVRXV=E01S,e1BL]DC8?F/&12SN4^]0[#0TFeb/>?TfCA;=V+D/LeH^1cI?A
f]3FfIc.MO4XdK7D=\H_N8-E@bRQ-A5@#-LY<SfSZ113@,RK#@2^87<36>&?aD-X
=DeHUY)GB5c[O,70bcJIA;49aA_67Bb=KZU-Aedc8/57;g.UQWfVVDU[DC;B<&]:
QKN04:?G=Zb:D5Wb\)GdK^A:H,bBMHFQTCY<cb8KZUYM5eP>K/U_\<V[06YTdIUa
Ae-WI4ZH;.S8P1SM+[DG.Z33dQdRKA\0=aQ408K[]f@P/M(T.K&29ICF\_>dW:b@
(9J=Sc72D7NgIW?3H>?5EeNN_VY\&RH4_4]]W;MDQd,UH-F=6.@V6g,W;4=VefW;
c2[WS.f5E:7+I5V[@Af,fXe,fI.QgXC&N>1Z/PD^fXU8dK5P+PS;F\J8>bL3U:e?
V=8&^Ibc^<NOI->>WB#cKSXQ-GI>,;#4=-.:=JB\X(cHZaD.DGZJ-U+N_f:6B3>1
_OJ<^YOG<Y+La9f;H;:P^^c_AXD,5b2K(R3a^S.YZMfUT1CV.D<))\A)IgI&7/9?
Y;WR;:[4?:267/[OWc)b?/G&W(5&]@OMa\:d?DX1/Q/D5fad[+G<=a3be^D#F[f^
Hba(:?:<;aU-X?>f&#I@(dW,82)<?V/Y#d#G^62+Ze4V:Zg-)CB3MDFJNI/dRWA?
>&BcG?31GM]c/eI4?E;0:(F;2R^U-Q8)EDZ/QA7JTHdO4(O_UaAKWf?eE5L^A#YD
5K+<c=ZaB,X\GZV&]S1gBeBg55JK#7TDN+)41G#0W<Qf2[0HB5[8FcB53f@@CW2a
O5Ig?Q+\XffH>V-3?/6TW@ad#XPWHg@aRB(DZUYcR[,fNC-HGa6KN?#OU1/W>+R(
FEWK4+-:]TcdgY><.)X(?dQHKa?P:OS6B2WREG->_>90ZP@Q0Se>:3<-JH1eCS?P
]2A4OSC_S)6b#bVSYeWXP(C#>;]+D@=cI66;44;U,NAMZ_cFX-bKdaW&6JWKAd2H
C:EGXW\BbZ]HAg,a=QRYg/VJ8PG4>;>f#;[\(K)U02CA;.&d#D\C(_VMY+GYN1CW
ga45.C(S3Qc=]GX.aGc#,7OK<8+cf@SZ3KL.18H(L;fQ+e,P)f+5c,2E<<&.RF?C
4.DM2@K#;:W2H:IE/E5fOGO?)W?0PEf?8PELR<R539:8WgQ[3WIX[/.0Q+<2Q^Q[
Y,M_0GNVGE0-D,:ag3>&7.fMU(c7X-29_[aXBME8A3)V6-aeV>?_K\FYN0Pa<0_=
?LD<)H_EdH,KP>1J:,bVMJAe4G\T(=.H_&UV^Ra+8H9S4<dDM&7EMOPfO\=VL(X.
<.A?:9)S4XU28SfZd=>G3f0H068VDIF.3O-[[K^&HFAb4>-YZ^B\X3F/.gc)528;
@H3G@&1a3Ff?UPNcZG9+Ofb0.UKL[_AUA2902>5f7OB>gO-f>3--T#?Yb4-A+MYK
(ISTd(+;L_Y;7A#M.BAU&7/EOIFNO8C+T-d+ge+cKP1M6.EKaUUX]&F=?_^,BMI)
PIZ?UW)ML?g3L4?.:8cHfT^a.GET7)RRZ25<^f^S4N)NZGGBJfDPFbecYg@HC>F3
(O#U)T+B2_)f)g/)CEJPgcETbG@K6T\4.[@ffI3gN\Sc7.aV91:;g)4fRE5Gd)?F
3K?PB9gJ:(2FK8e/<7f:=1_agK_G7NXD[c7UD\[Td@#M+;<eg#)SX@d(1I9IM>[N
I?9,MODU/:939GZ(7)EQ\8dI0E]S#7^/5>(2(I)AEIbN>:OU=Y6ELTY<B+]-(5Wb
9c\ZYSQgK/MF(I+S5N#g>f^@T]\PF(dH1/Pa45;OOILa9/AI<9(8:U28BgaBXGVe
&2C(YAG>J&bLM3^E+75](>1eZOH_)cZ>W@H9LGR<fRO+5@gF(QC&J7d>^9c@-cR9
=V9OL&?DaL&1DIZW\Gg-ZYP^=#H45V#U45@P>;V8BF3.Qa9@;4Xdd6I^.&SOR>Nc
5a((e3?78f=bB=:-E0L1)R#6QO^+[XeQfUG&7D])FH:+3+OUQU8XTC&3GEaP=NW.
D(NdK:F/U(()B+=dPF.X.=AW@64^AKHP:dT0[\R_AB0aG5K#10/BeM2geL(,]af]
6RW3N-S>6G+AUKOXA0ZU.c&RN-X>7U?ZD5C=.0OQPZ(PS[&LXF&a6#/3>40dH8MF
8=V/1f1L4T+-DCE/51,+.3f7d1IV6BIbZR#e?_gTJ:1K]c@L^SQK.IJ3=_+&7E3T
a@YPRG;O;A]6eg_4+M-F(7.<6J9+RZg0<G>F2?,H]H1^;XL2Y.DM#&S,[.RDc]A+
-Z-=^#3;I/1EaXA3^<<<PVY/c))2S>Z,LO.;ae[ONZ?JV>&(fe2^)[DTX<BdC9>c
BUUc1R36I32ZLSW3+acD9[A?N@S6/8gHWfM[ag>EWIg]R+6X]//T71/><cA9]9-8
aH]83d^ZF4?DQKJTZ+.(P]OVS;d=CG3Q<:_N7EQL5<[O#U^HOdfcAd^R(-995E<V
?>C/SScVE^N>]/90+dA=(B,-IF/eA[a5Z.Q/GaJAA\UT15N1Y.-eV)N=fOS\NX_A
.:4?2_U(QWL)>X2;9.9C;M2#+aCXP4D\<9b8WBWb7.&^1d1d8N@U9.VWQf=G\[;G
DEC/=gG)[f(dRC]11-03VI.M+4\@Hf_D2Vb<c:QTe6ff1>\/(EHg3JZ;#X(S7a54
9geDRYKg+;M1=M9=0T/]HLGV0V7:VaOfWT?P-D43ANMPGOX33NBA:&<+--K-4)LK
Ue4?PI&?6_7;AW\7=OOUI3B2Ae=3(1cE[?\+-:WZ/L9UX5AcdN=NHN&^GLXb>3?3
Ma:S73D=WD;9d.^c\:@U=8f>M90A8b>78P7F(WRX[6?b:WQ,,Ie^R1Of)GJ&UV70
.L04b[C&.AP.7QGHJ<09/&0K+^<dGa@6/#1>-OU>T>gW72GfO6#f\EF^RcAfK_.G
.X5-GJF3ab\G[EfFZ]8S>GdB<F,<+#AbegAgB]2.RfWVS;bCe=_e//fMFCVb<NXZ
\e1WLX5:\D2.2(fA\C#Z-=F0cS<;Z4@VMPg)/fgJ)+=)40L^.=MFcUWI9CdK(4J<
cTGF<H9J&NQRK5cQcFcA?dK4JR\UAbS,([:KXS?22+RS9=gV@)+EDYI=,5K,+PAF
J5K<65fVHHZ/+Gb)0YP,@63;f3<T\B-b)2_#ZY/g)&c7&^C/ZK0TT/5#XM)K:&^N
.LdK89)cV<#b0^V/7aSbG9<OaULU)5:&K>S7FI6HS6.<#e?X)J,;2ER\Z;&KW/GG
AAC&&:8D3Mec\SaT>LQ<N(B?X;Ha;^f6?cdgCd[\deQH+^Me<[PLIe&f1ba_Q)HV
,:V??AFFTU(^A#+M./01IGZJK<7fcFW1SMVQ#I_7[K]dELXLH.VV4DU?=<=6Oag8
O\_,6_J\OSS5N54bI:2aZ?J535TL4J;&P_&3U2X#5NI_PZ0G#7)IcPfDP4WX6U4B
Va#<CfPfEB7&g6ca)#E+KaG:/-3]AH=4\Y?#L3>GOd[7Y&7ABU:aKO-e465FU6]&
O.+af@PBHT8T5EV3@H-(cPD:M+>2SG;+)bO;-:\+#]/B/[_8:RG6^WS@F@9[9;[(
XgY+7>JL6,CNYeOJ2WL-,=dTfHa6K^6+ZPG)[:c:29e7+d@eT3-aXO^Db1H=R)RP
c,P&0HX_4,P3L\(:GQ>;MC\gc[-T/-\Z,A.B@>cH/\Y[.d(a-d[\9bHE&CA61;4B
.>Y:_2H:d/Qc/ROZ51Z]SM4LTE&.A[QZQ_^CE2N^EC\Qa)P4;&gZGVJN#a:^L.1N
S1G/6-&P<N5aO.KKDD?5eSEcC<Q\&=6g9YeX/(/L6,bB-CB#04?L-Dg]-KcG+828
PSX0J0;^W#]+96_f.N+3JK=ADW;(fa?SL0_KNKM/]]d2eE?cL:)_9F:\2TLYA#b8
BK0\?P,?J8I0fdd#S<@)S:HA?(FU:K>^B8d28:^Ja5DN5:\>1E#@PWAa_8S>8TTL
B=@/VI0+eTcN)GZ[E52]ff.B^]Q[DLT=Z+;7>Sb4[&AFV-27MVf\gAa1@BVWgY]F
L\TI\Ma,2>H9bZMd@BQ?D#:6H+R^OU>TNCcK-@7@,,<51_9-C]OdMXW9eDb)58bH
EMM[cc_CNKS6M>J]AE4RGR@2AIF[[G7=TVR1HX-8P4(48:V+3bNY9^+MV#5&c9PH
]S[]^DG3gX2IgN^9>]1;_bH;\F[\M^AF0(KW8<\ES>Y<=?W4BQ,RC=&A;3W3WeC(
]BagMJG\FD)>.L6@9@Xg@B)PNP>8B08T\a[^TMB-;7\0)<+-@7C/:75bR8+GQ,A[
+KQS^,8a]LPLO_:N&EZeCHRJ=AN^U-E&87afd8@O5J^e=b)6+>;+:_Gf<bbENVD_
I:Aa_.&)OdAZ-)8P/\b#XL5LNOQC(ARU#-L/3KO6ABZ05GG&^cG]&HH8d(S,\O\Z
+T.79NMTI0gRJ<^PS@IWZYYS608JDM]DZd6:LW(OSX40Sg6WYZ4FAD5G6T:EMFX]
C0,AcHbDMOfP7K/LXe^Y&:/=;SU[MOLXJaNR9N]Z;P-A(/W/=<GG?:<(SC+a0V-V
?4WP@fIV]>W(e+B)gKI/.LUa_,+1\JT3K[Y84;U?\X;ZKXFUgU-#Mea&M8-a>)Y?
g4VQQ@f\=UR109Sg6H6Lc&67P_ZZP\-3gL?B]FM#Q&J12WeL7Y^ffH].P#:BFe2B
gZ2R.10Ke-aE)C:GdNfW+:P:]LS9a-LWU>T5^:NIM^FVIBgaWMgIQ/7Z8#abKS[;
^6B2fH)2H]XRQ#LW(g(L^^YYCGBa1##F)T+[J^X8DZ^cW(@JaY,2H6JgfQE3_TIX
/fC,0d/ZAAL[&b8gADT&UYGP1-fUKB>(HC29L=<,QWINbY\>??-PWd,8G&GTg5d9
D?.fR?d,JA:2+_+[8aAII51e=gB581WN[bP9ADHS38;\F4V94d]2[d+?fG3dE\V_
b[8LObMXP42/KW3L,T0<CKPeE28dM_:>J7ZB-7eY_)L]O@/]XH^O4?M8[_aV#(2e
V1]MN96?)QIRUGd?3])W@-/I6]baZ@a2LaV6KRA]AO;(/3+.71G=Q^;D6@J=.AO2
.g<\T]TF8-BCW4_8.V)OHN#HGR_\B=J3/NQ1K5?86[:ETQ5@A:.0+6QUIHQRTQcB
W[E+BK6,d8K_Ya-cTN#e43_@:4-Q)?X[16M_Y?VW?67J\BGCe\C6901#<a2)[6[_
gAR+V/>X<U[V5/b;Jg0X5ZO0C9^?X9bCL+LPC.EN@.7/cGc)>O#IFLd&dCFLdDAB
#AC#5VgKcEF7dec4IT8RJ<(;3VT?EGbK(GTdZDH/7/@gE.2OKSI<eDd7_G-bY5QK
C1M<=f=2RTJG_+[a[(bK./HZHP\d8YFRJ47]LQKeDG_dN03J,FRH79:ST,Y3.[L]
e0+D#afB1YG)9._XLMdB#8TI1_)e#>@VBT>LP50V=a]f_H;8fbgW(>ARUK:cgTA4
FS+A9@MVV:7NQ#e2)1@UD=)-B5>N[?=MfbH:\S_P,U4>7J@IAgIK-Dc3?TW6\c__
JM^E[Ae<(Z[HeXYV#=@O^.c2RE:?5;YO1-RY,/1ce8HBZE<,=/bWO/WXLEfJ-D<T
Ra+.e=5g>IG<@O&V-:^+?U4JRC4YANI@ZCWc-83)=-23H;D&,SbL_@;UN;I=&Y]:
I#;Y5fXC6Qbc]<MTDXLS9FW_=C#:C>T3P-2E3,_1(/JAf:RH3W5R;e8X)\DdHZbH
IDRIK&U7Y^fI?Q-S+O]]1FI.:K]<fYC0<3RVeF:UD&c)&/7=O=1\c[Y-YJ);J7:?
WZ?#&9P_9B,gX0\Xc9\K))gZAOHcS=TMZb)RDYQ;BXIZOV2Cb@/R]+g<1.+,_D@)
eVC2f35f?A8:[=Lf)_W-+CGH0OCbBZ]eO--+MQ7NB(aK#Q>LO0Y3e1KN.P3XCHD(
(<&KX(YUe(M.;?#;;B9aC&)U785g5UFYPX\PU.C_Q6HH=e@Mc4#8=IK)W4.-1g/W
4PW=.ZPR-SUWgeMWdPMH6S=gW+?+2F=#KJF5(5T_dB?1Zg@7c/6f_]8GXHS3NN:M
6LQ7.d6,<.FGGLR]8_Y9IHK)[?K]#YO^I]^),NF\Cd()\<E[Z7GU+8:IX[EI,VM)
2#I62<BOSATfT(P@IZ=-aYL>1A@W0KX&4,20\dVED;1M6Q[]d[>Y2A:W?UU0,-1\
2M/D]EK&,,gSO4MR_9W/QIX,=E1L_IbGM/0Q=YS(EU=UHIGDNAL.O#&U2@^_]90(
ORf8J2Z42FLCO==ZVHOH+[+ZV9>L^D2^PcTT0&>?XeTA.>7Vgeg](A;0#DKV_[>L
=AZAL7RX+)96)XCW.&K6&9LOb#&[\1NV0c;AH.-#aSEa7WZKUBWX<LVg^F<1PDA=
GQGOg(<NeZI>6AaT8gb)a-\#]?d@DG-^6>O5:^H#C8dD)eXD6Y[?\ACH\deOUB@R
YH[4ENb?M]e=??T=ECbY#Z4?cg;H.>6cV):JV4)7]X2;2>ZV[@794DGG&eRc4>-X
@=8)WC-7Eb?W+d2IeCJg7CA<47f)\;-/575KU2DDPgB1,JNKK2EVTC@X86JSH&gX
LSXH3\cXPP#RfCa2H.A@TLgg_L4Pe+1B(_E=X\OR_8AdO10SX7UB38(@e8.4@[(1
[IXU8,_#&K=<LfF6GRfW[&AWOXS?C;3,375(Pe99dgSGBVCH#.G23G>\;7\D1VbU
\^7Z>[,6f;WH.ScMX@g1WP3@_Y^R?R&bS+Z6=LeP0/0G<[Qf0R4>X4<(,V7b;;1C
/T9OQT_R]eVQW3H=S#0,;#(KcF1W\WUaPLK>Z34Md.@a#XL^?g@Z:?;MCM(FZ#36
]?VcU7U8OVWNM@4E(04BCHX8Hfb[74Waf\R:W+==Z1>>\PM0g/R+N)&[/_.:d4D@
;c3A>E:O=JM\-Hf_RO5F##4#WPHVgS2\M0PQC>[.[_RNOTR3YK^@D-@Q+e7-VP(H
MU5H8@1dO6J]TTS/1>?AK]8ZU]^&P[Y[V7bIRH49+:\fQ4J9L,Db16.4[<3BOSZ&
;eV,eaY5(?K6RIJ+2&Y)NEW#?41Td;.G]48];U5eRN4W(8RNdSfgV^9_RT6FWVaI
/WD.0&(7KB]O^@4/?>a1>&d&.I[]G<_+^1a&?U/OR(9c=.PGIK7\R?c(e9:L[A&#
/P)Vf9.2W=bdQ[=a(E=30WBHZe:M_^/>>6Z901^4SQP+CaN?+TGPL]SeWZ\ZHMXT
?QXQ32@f]\8RQ0\VeJ8+BO.5HDF5S)A5AS:&,9=>90\3YE0TPbG.HcSJQ[::MZ8_
g??YdC>e@&O<.LX.V/[_BRCYKXeTC/aNTYVVSYU1+I8K4NO=:7f8,?<])3\F86YC
I_\Z6X81=LYg\7\7fKL+e6P&/Y=>]5)?SFX(5:(?RE96(:EU2BbX2_1c>6FAR@cd
N?Zg,POUGJMcfR42PAE9I9J>5SUc+A]V6g-[Z8HVW?:ZD[Y9.Z<2BHfI22RT7(6U
#&#SIS7T@L^&f^5L&>Ha.aPTV^c6DSP6-?DUP94<XUJOSa](ME<+aZ3/TdcCZF7\
cRa3.OZZ);08FW&dA;DO,[\/a^O>H_Ia,B:0?Lf/BZf+Pb#WT28LXWJdb1eJK]SH
[V9K>2gZ#dJXe0;gW@a43A@E=8&L65:UU&NMF-;#EY8Y(X>+TBQ+]SQY,+b4PI)c
)cdY.dJWJ&QbbcVSd;NLcK=C7=.\CM86<W+>DHFWAT&Eb70U1S2_JQUJ(]:^S>8,
P8;G3-aGA@/+\:\a6e#WTEb^6R<.4d:N,<QB]L?3AF1MaE_X)WT@XJDa9/f^RN,A
a0-VU6SVGaBHEUc]=VI^3@8H@\[)\c(KHfKZ,[8+@eVE]gBQ3)7XZ,7^XZ,NBC6E
Hf^ZOX:AbGL<_Z0GVb(2A<_C1B78MUF=OQdWN^(c<&-dMR5e^e=OOSWIUC>I=[9O
YDe\==SJ?M\?:F6JUL8GY1=.He??61+b7U9>d/PZJ,3c^A1d:f+O/;bB26eDBOYI
&@7N-X@UO,-G.IK[U@8E\.5K/;05gIA-GIAQ5E[,D4S7Q/U,WKDd>@MCG&YdcI@/
0F@0]&M4ENK(GADNJKeKMD=4[P?T6K.b&K2L^<5=H>>1c=FG9dXT+NFU]5&A_RP8
^N,f(_eRU#)HML+P#^@(N]F^GEeEOee;.2BQ/J]&e\GVfg;=R^?<G-fCQA)/NgCY
#^_E(3X7TA.,eL<VRFa=AcdA9b><:+e[+f=4]H>S6aD95M()MVR#2.J#5L6cFSca
O/e;4c6c5I^5C;_ef7U8EA>bL8E]GLE529Z/W:C2g0<S3:?QZ8-@6a9ZBdOEYGR\
LTb8+Dd_((192G<H^UNJ1^b)QB^XMK1Y&YO3RB@C#.9F<;g@/M+JQCQT\NcY1&VR
(,Z\@&?>][FAZL8HW\6JeB]?RVWa#dbT_\aTN^K<=^W)?E]g&;1)W1:G)C2]4+(U
ENN/V)()E6Z;KW8ILJ<IgHQ?Z<N.;.d:VF0H<6@^/LDLe?QR+L5=Z.VRc\0Ig&UI
<O=gQ/6+7g2BQY-AFR#[HEM+O-d(</;;PLc_<6b&2b@&PF?J07dHAa/Y.@_1Z3WJ
FQ;H;^?)/#N(W;F4E5eWe^R1OPC)Nc<:B_5G^TT<gf)<WQY-W9K](=L.BXF89W@6
2>cb@727_Q\=LdH+MM8V2=VC+e?L&.YNTP[\ZBGV/3eB)J.-GSV]/Ke2_V;Jc\3>
-Q),)Q\BOLR9S0A2JGE814:e5NI0Nb[M3E2Y&X]]P7Q:[SH7<,O2K\CX(H8V@L]#
1/7b,4EN[9g&1)_<HJLB5GOS[?4M-NI&N(O@K+WK>_,J56.H[E+ffaL/_QY9>&)P
0bV(Z8.fQFK5.,JIIU.CNG4E\3eF-eVaM5G=<d07>SU^RSNfTH[30N0e91L2VI<_
<ZC.@//A\,Zgd1bfVFG:R09b&B7YT4<7-3b\>/adOU\.WET^>]#UYVC+SUSYIDX@
_AOCY#OPD79G>-Xf;-;IELEa.#02c__FJ1FPKUg(6_//(R;(8/UG>=g,#RN5L#?>
eTdA[=/g-).])YKZTRaHb_ZK0T;2:dH];UNYWC6R,_g(71-,b35db>F#3aFd[M2,
\g7J>BS.)C083WUb83A7A6WYWC3gfa8=QA4(K7_G=+1FF=9WB_8QC)QH+42>(C=M
U2E=.(@cdXgHE#W[UP2YVIEJ88R\I>P(NOHHB((D7E#@0dUAO9]U6C>)a>bI)C(8
/g^c;N_M3X=#)ZXOe=4@P.V#F#YJ[2]7fU+,YaP<bIXM7&P6FLOJC=+@X5SPbTF[
4E#Z_U09-DX>ea.N0FgB8]9aBLU(+-B_<HONG6&,;+BEJ]P>.3cWNYV5+gd85+LW
DJA/#?C71&bM=^C^&D3=3_>Cd-B7NG,#e.\O+5fdSR\.=;(Q=,8ZWK=>.&\f3@R2
>cbc:/WOA833eSRAdCP:.O)9?gBX[@XX:C8>N1@W/\1G;9R)7EP>5Z(aKSc<VHYY
]H]6P@Dd84YT7G0UD/GC1c6;G:XBYGYX^3984Eab8R0Af&4V=IT#RLHU)_(^4Ca<
N>,>&[cf[#Q_,RK6L+/PV87eV2DBEO+6&^M52K?HQ+_fRb.dE@[M^:B+(3Yg7F^O
3@DUZ-Kc^LJ0BQQP5RT2[7Eef1PWO@/S7[,,Q=+/aIQ:2/-,dXW:T)@Wb,G7b#1J
2NV?KUF3D2O8E:dNQ??E)\TccJd,eUG<.eH6a_641CPAKWWQ+0]]Pd?e;E8a=SB,
JVg/T+QHe^e(>Z)\6]U;K@5eSW)+[eDa5_#F^18g63A>WNIPBgbd[F0N1#S/=W?e
/R)@FQcM/P2eHH#-Ng4.&(7fNgJH;[ZA3]W620F0?>8U3)EW8IdA.)7_-P]W;UdG
YAT<=fQC:#_/7^dH,YA[YeEV?RLePF1-(#[?1<X[URIH9D3eZ^9VfB2MKR[LXaZ)
^-,,S-/W[f@+Se+dJa#_Q=fY_3bb:<S;J@\Y1-@fLOQ8CM[BaEae#L/AF[V]ICVU
AgUVeeF(WcY4PS\&(Z;g>42Q4\,?eF<8Og58NNXO5\,a0N@ZX>ISGS?(Q5?,UA]=
KgI=2;6I24.OLA7.VSWd_ZTT#2dQcOGF3S@e66#=_JJNEc.[^WXG.##V/0c)F1RC
D7V1VUVG2S=gMQ-K7,aN;TI&,OUd4>M\J8YbK.A--VMD1_:1Z?23KXAN^@3^KeE?
OZ;XIX=)MG_6ZSI>WT0,[5X0ENI_AOY:B\E._XS(8dQ&aB8R(D5WP-#H3aO6,UO7
V/@c&O=\e_&U.BgfK@4:V;GK/g+TS-3;#W30>g4bHPT+\,-\Y)J_5C&J(fQ@WS7B
G?Sf>:1MB3#0VUR(,-JFXCFEW8fg-OIE1JW.(MU_MHBTE]A90J=F_W]6?;)7I4dG
JXA#(0Kf3^B(1/;A2Nag(Fa3KPFXG8,Pbg0:T<G,;WYb1-5[_KJ]:0<T5PL<?L<4
;78YETB=]02(SZXQ@1A^gN@f<K#_W&4[Z65CfLR<ET9E:14aEETbC^eKb_JNFfB^
3G0ggFT:eQM1X+MX^_f<U(>W#S-JNaLUX)0R104FKS1;?3W&aO7FbbF^CY-Y)4\N
Q6,b6LB#EVU&YbL^?7]A3Pg-<-D-a86IBaLF#a;BWQ&,SEUX91/B/gE=J.-4(U9V
DKSOJef>@gcf(6_bR+/XI67949(7d#?8CX6fe5fcF?_(B/&cbD@@&c>,+<X1_D[J
KU8U1/2RQbAVWJU+1L/FQ?Kb</:E+FeF^FPN2Y)&IP+2BP1/<dEbXN==ZB.DPb1?
5+GD--SgZOD\2)@O&K6Cce@gH.bOAG]1S;Ua=-]O\TX[5?TeKK\d+H+I@e+C.)2G
dTg5eN;CG5LS(9V5f=-c#PI>&#D\#J&U/gRK17Z44gUHBNBS.E+7JacT4^ZGNSHd
5W0P:^MVa[2T[G/[91T,c]A6H&R:)U@2F((UTU?Dg/HSCWd#?=#NUCW6Hc5]ccT@
)bN8d^^BUB)(6?M+Qf8a^>9_[JA[<7C3/&=@G>^SMPe5>fF#Z4WJ,U6TR:Rc/33N
QFOUVTN;[E++D1D;O;QTHf&8#0K0P.;F+B[PdL)@2;@NY@2a,dOaMK=J194D\d8-
)g1OL2)H^P(:.VSIK\5DE(41UFH@e<@I&T@D?4Ob[A)4QG+:/c?,7J8,,1]PJT3+
<2GZ.YD;&3G6c-[-4HL^bTOSDU].LS<LAV)>DBcI;>0F^OYYd+ZZ4<\6EY-=6?1^
;V>TP06S:&-:M(SDAF-38gNMWMfS,OVO-gW/_d#e-KD,c,[M-S^L3g5W@Z.V-?VR
XdXXX/2,T&WR3CF\X/QSdCGc.a]J\\9f8]JT^PN15dJeNJ4;AfJg&[/gU>[\(>>9
Q,9+HD>WG3X#UgJ/F5P=#^(.O;XP1+W\8Z_Yg#.OS3A4eQaQH_E@4PO^+@.Y@RZ^
:cU._EM\8<=GeNg8OZ))D1FaZ\eM_RWM-0)L9YD#9fY56.<VfY-9eB5:AMP[S(N+
I6g4ZXV2F5M<d2(P?7#IR>1\U7:9?&7cbFd:DNVP\P>I:W37DLEE,PPMJdeRF7I^
2UgS/,8AYC&/A?Ad?>c;-X+=I,NH_J5@\XJ,C\XDcZcHbb?fI99HbZ6=dPaD-IPW
S#(<D=LH(.=O(SI,=Q1B1?\;fO96d[?Nf#Z-0=I2/gM>N#X9UG)#&ZT_=d<PO#J^
(968F#6QG9Jg\POYY;V3P;E7Cb>@/aFdQKRX5]&1bFbT(>-/,XXZ>bXJAYNT<&7<
_YJI0:;)MT@.GA]@XOJ_CE>W;IOYIaPdSUXMaEd-Ja8ZS3>,9Y?d4XBf;Ia)^U#P
1BLf)Z11@MW9=AS>#0>4[SW^g0]GROC9VaGEVK4)>ZN<[\J>fO;)4F=W+N=c[PEI
RNOXSKaAFF?e,9+6.SYPaIF@gB^faZW5e<X@,EK(=WeJ8Y/J^BcJIALP.MB[OJPG
2;\[D7I)AOMR8]]^-f:LR,<[OMJ+62g.4E&AOX:Pf\+,J-a\XR8W0@9d4^Hf[IIE
(,^d?HLKQ4a75H@1ZEM9g[HG4;,4(?;?fbW2#EXY.a-=MJ;<8+>U+05)U2T6]+S+
g5VWUN.,J,K.SU+5gB12[S.]X4)JdJ<1.&N0eYaZCBD))P4Q>cA7bAZ#_9.&;S?&
K3,3:([1DeC3gV/d?)J3cd_-6H_\@G>R4TA&(CDF,<,4NSOSNS?VCDM,Y-EN&Mad
A[5T&-UZM<42V,BPfdNFRbEY76^@CSHRR5;\VJ@&Bc:KT+2d.,Sag[ICKbEVgcRW
fa63/.^Lg]_QdgBef#gg#G#5(0Q2e^9STY5MPD,2E0UU+bb)?K.&1<bF?P)-UZe\
XJ:-.=J151aN[&UAMJ1gHHSM>JdD&4I84MD]46dM;bgG5GKZ^K^eWIZ=.G^K/0I6
3R+Wg[W:&KB)a>3^bWc>4HVgURd.2>Z7NA]?FfCZ^GGTI;L9P-1cQLbcV>#0c;?S
);M=NF?3FJ1I]?L7&3B3K-CbL;b#T<EO8LM/THFZA)44L_7de&bQ0L5JAHde3T4P
@D;K#fI=]S,7YA^f^P=8+J(\]5c<7O2BMe3OD>TTKOcYM(c9K8N\;+0@O;.5SaMO
X:[R?6\_O@\U[G\d1N<T9c8<KTOQQ\X/AMLad2A^FIag66C)X79eeCDH;+#CF>2^
Z)GC3-RZc\?O4e+UAP,.bGIEX/;MXDV8H+<U)#IE?,&W=#8B6AR@]>1N39L5L@?>
]P^F^[9X:KSeHM(C)7@8+,=2GY6[RUC\.0&D2Rd=N=)cO4-gPb<T,,RB[B5-B.fA
6ZK\Y>M0:G+[/XZ91EC)UT47Z;aAECP>1c4#d:2E^@=TC,R]X1Qcc9M6S@fc-;]Y
dD9-F0H7[>]SO<bb]K:@UI/P[;5Z)g+eW+@1)4H<TAfU>55/_[(^ZNFVW4P<gWL6
+.S7V-?/X?Ke)<,6f<(KJ//]ebf7T7Y#?^XO1cCg:b-SC8CB9[21e=GQCd]A<)F8
/LW9Y?Tbf0Vc;A&-6;&VEfPbJGA:1Y,QK<X7(E-NT<+]6^Z@LB:RC>FUeX4RA2W(
5+WL^Z9>(10aC&--DMM]f44X)AAHM6/TY[76Q&@XWQ^\[34^78cI,L\A91c<RZ4+
XH+V;<;JQ2TF4WS>K:9Z5GQ;VeEV9UFf/6;N:OU6;TF&bCY4.Q7CQPD@4c\d_^J,
,>@1/(6L1SXUS?UVQPS<:a<bdPa06#0)>5QCG+<Q\<C-5\@EOHCR5@P?(/[2cc<D
@Jb]70;>2>J]CPCM70M<2DJVO26#_/[FOS-=<R6U@g-II;,?&EX#c/\N5K?H-^Z5
M1>8V=T_L]DMdN\ED:C7b&(XHedQ20?E3U/Q70)3,^ZcdY@B+HS)Xc6^A?G[?@7@
3fFN0D.#ZW9(V&/IfH.K4W)F]G,GbeDe0O\SXA2<P2(Fa+&?N@T0dV7C[ZHW/<UY
1701@(Z18=T_M24]R[QQe7/=Va0IL[O@a6Ng)A18UaZ7H6<X-_1.D?\BD(C9<A?a
B^egK(,JJg&J/D_YO>I+CM0[M+(e.>N34IU[Y1d_\F6?E\NAC:G/C.NLd/,]4?ES
6@26[e.KIKabXXHe2=\D[/++&+[54cSO1FS_54N&fU[NAO4=[X5+,[g>F5E0BJ^K
_TZ@5H5.^_DgOA>e_<+6]&2aFK88bY]7cW.=(M)29\@a252UI/-@]IeWbTAEOZ?M
,IcSdKQ:P:K-R</cdS]L,1PfX?bV1\[4Sf^WR\9A2G3[].cLc2Y=^Q<W\(Ab.?R>
Lc55STV;P8CCb2ON7bU([+2KN<,Cfa,dW:3)9P:KdU9e>2RR?Z0HA@TY38[7RJ45
,7I2<[?J8M8aJ:_W5101+fODH3dWb#_\6\YA74[P5[41+BQQJKZEPcM4JZE.W/MF
...P#,WdOO&,5V]>@_BN73+/.1;e/,)=C]]T;>3^-0FE1:^6P>-3>e\a:).F2W9#
e#S/c(=FL:&]OXTgP\)@9_f-WQYJc:A<N4\)MFPSPE2F2K]ERJc(SM-H1eE)PK+N
E1^=LPY<X5Pe]?a-_Rc7(OIM)<^QAEC^C+W64,630B/S5b/Y<)@XN(MM<NT,LUdB
bQ7XOTEONabUK#-FK;I7QA_KHLT3JNV&d@.eL8C&7&Z&YCZ&RN?&8PT53OeaWGb7
[>]R[5CXfVW_.SgHSW<a]88)IO<gPdQRD5b>T2:K+BEgMg+,_5NNYg;OD4M7g]26
P>Eef<9I=KB6S++8/?H83&@^O?U<3d6#O-YI7KH[E[@6N3ZVUa882H11Lag[ZDPT
+U=F8g,:f:FK4bR@>JW<[8Z6C\F\C6.7UW:+b1L7F&M7&G3#C;bQVZd;^edebX0W
MCVNbe66(_CM8SGJ1R>Fa6QKC&gb:14WB^Q#Ka#[Gf9?;,@\L>?R9;/,L5,?S85&
EG+U-9Tg47>>KB.(ZR:P5H3f5:31\)N0[XeY,14BdK2]@Y\5b1>ed,&R\BF+__a1
QZ-\H.>8?Y3^K[X0>aZJZ:SHcEZ4/HfJcZMVMD&Kg)KQPJ2:W8#([?g[MbG-JW./
]L&/KL>GQXSeQ@;K7_cON9&3Z;JX:=#K)Y4gcONL-Ib1@BHae0MA5F(bY(MO((_M
E(C>BDMD>fIG]ZOT=WD#GY3BKYf-M1:9#bT(HCS7O_TQ;P0S#\b3#J_LfU;&/K]&
@)@@9^;a#g\Q?PDYf1MN[Y[]=b1])1\VCRH_>&F^PB31)NQcSMD0+IU@H6FL\VQ>
L;[4#NW.7@XG^V>QTP=PIN9GL@<eERgJ\WUd=Q/fB8^@J&LN_9SZ+c[6/K^gTd>[
H@/+>TFW@8S_-b#]U^<UMC;P#U]G;\##=G#;b8B(S>Z=PaPW\XX_=<6&F/MM]6&c
=?_aa<8eB-P1c[OZe0dT?/,8MCFHF^Z\C<KcDKE57X=>IY=J=V_c<E3L/)M6@TXN
_CUX9_1H^N\a^E4TX56<_?.VC,Q\.0^)AY#[4CaW>91.VT2.UE[a[T[DITE<<=EG
8N\8S[B2I-972/&3^-P39GOa9DD4M83\e+G>K]/XXX#7R#:(HIg5_9VEdgSZ6=,W
DJ]\YYT>.BNEX>KU8:_<)00>GO,=X&7_IFU:6?@3)<HD8[99EP64>HJ9IbK/fX2/
>8.]>1T6Z6OQ(f,N+e98cXMO4X[GA@\)/1:<LQgb0:fV>9XUa9..SDNTCM7dUB@7
.Sd#M^#5V4F-3<NG[7NQ;+/VQ>V#WR-R]<UH_>Q1d&J0AfZ0M1&gUeANcA2g)G.8
8.(E40E3CRcb,U[@cF9.,QNXBPOJM3PWKfe4-D@d1+Xc:_0DKTEPa-I<JD0=WBIT
/YM6ELV3<_S[OdZ+aZD@E)LKZ-AE2RH549TK3&#>X8Re;^EXER&TgQXV[2RK^PL5
f6&3ZTJM.5IGI&JTZ=MS5A+:d2(Gc(1C)NTTB_KaFTAK@]e9U\TV=6MABBTaX98V
EMaR>,La?E3D+7[=[-#:EB:9N)DL(7SQD;cM:TW7HZ&SO^FT#>PUQ:&6XF\.VCIZ
eY8:CF>\CO05[OBgLE5M.:;aCbR-)O#(H](3BEfb]U9G^&OZOY3IZ@Z8#068>YV@
CGVd#c,^FWg)],gFZ_J##0A3#b8A:?GgeB@>UGT^X+R(245X^7dB/(B7?BPc4W&8
Q-75g&)OI@YX;6;]?B\J[K&g_-(KVc.4YdVD1A^#7L&O#N)=DcNG&^5T4:^S;aOL
X^Q=F1(YT7.)WQ)23@.R_2-A;@C&365341V7c>?f^9aW6\e-L\06&:@7?F/I9(L+
35,Ff9c@[Z>HCbNSR/TVS5]cR37,>@T?>8cKY:=N)R@_6SQB75=cJ(7;_e^P\==L
>dO<]gUddL>YdYa^T^:40XTH..4g7RS:fM5FS_ZZ2(XS?R&9/]ZAK1f.8AY-)ad;
Oec4,]@A,NTaFe7>\+(^Ve=fgJ4NP+^J1:W85GY[BEA.CfVgS3GPKI?]G6R3+&^7
;Q(QaAT<DM<R:G_Gc+QVXJ:]:K<P5c@cHN_+a#gH&OTcaDR97Q:fX&WbI7;&/8I.
<FF;g@8E,[ITG#FfeC8MH[d+dQ:Q^F7-[-d^Xd<,B4b)\NAY@PHMCbRLg\.&ND+<
Y,V.gSPQe<JVW3DYKX(dg=H_[8M2@PJ@9ZKE28#V>W<&C?)W6(a-F3a,NNW16_0Z
)0HK6>R,Z?WP9MSdY94AA6YV94Kf0]\>?Ae<,bLA]R6,3eHa7>G\OPMR636<c\b.
b8JZ[IAUVGT=#TaR;_QWZ<a-+T)1a9Z<A73_1:P(;-6a/551c[]E1abbODSQPDI2
YZYZUYR]?=E_eaf</L)CWRH:bCT]9]Q3?WWI?BOM=R1&HL@9]YaM^&EH#Icd14S>
I6GS>RcFa2KO/FIPcVYF=DgCWWLI5C]8)db<-#gI,CV65O\BPFaFWV64FS,99\LI
:/e5GC7(77Y7YA+3CAGcSC@:+GU5(c_gKK&+BaRc:CGA2g?@O.H_>4VJ-P3Lf(U@
[2VdZ4=82-cXeU9:.9H=;7AD;GaT]FX#1<3N\D/-IJ:NFBR#A(4VXcTQgM,U#A\3
Mf=FC[]_611dCIO/g6B0FP_D&I=H1H2G(3FL(SQOE?.J.REF=#UQbBU\_HUP)(RF
>WZ3I;(d.8YD\]7KPGZZUU<fEK.(5>RM4HYK4-a(bR+?_;_U,.+GgTR[(R[[QDKQ
C#g,J-LF:96.ENNaA7\77AW\IL.2/2a/J-g.fUE87IMK)bBb8\-0#T7QLd^F2PT_
c3FB(P^2Zfda_gAV@.Z,Mc#NF8J((L4MJ9K^D[UCN2,f((^d/)(+EIXZ>B(2-[U^
1@fY;d#0b.R0[8S]<JH-MAA-=0PGUL)7UgK7@-MQ]<D^6)];/gT^5]/H;J/K?36I
fP\@6-S4TF/__J3TO]N:+B\64=9MH]<]WgPPXDF3_EJ4U)d:1e:S5Y(5(f5Q40,.
)QLg=2Q<QW-=Q#OMRR?EYE<M:OHXL4JR?M9QZ5Q-W85)@/QEM.:H4O\4OGggKfLP
9CG/+O&>Df]<]GKOX;S:TO5S2.@a8dF,G^@KI\FZUBTKFb9<H3JNS:^E0[MVMTC?
@2dQ?PX-&ZgGg:[^ZC#;0(T#Oa]U#YCUYBNTP^K=.NdUcCONWI6Qeb(C-K]f[W>Q
K749<?CK--8T.JO\CcTU7OHXASZUaF/@dND&HbJ>)7b92D1&TCg/UYc?E(;Fa44A
1IDcF3c\?dD\MYS_U@g#,MM8MP?V-59VAN>XAffUd[6XO8G(Y\G].gP4E3G]bJ8K
BD:Z\Q89=@2IZ?\F=:5U)Q60P/9F2/[[;6ACHC;BF3T<1N\E@aCV;gQfXV^,ZgZ2
ZRSEF]N4c:7C024[S<9.6Z(TS(SVS8,;ALHXO12SIc\YAG3;e-^7d^C47bI/;QM_
.d385/MBgd\N7QF,J8O[=Ka@3f(FGFHGP_4DP]-b39_QDD;GIER.;QdO9X#@PHN&
<#X3LWJ_V1&eRARbWTNTIaC?>NSRg>&+J,(ECQ8DZ(^O;c5<BSERJQ9]Jd-/4E@F
AX?W_@U_U8JXXc^.dB\7B)EcKGQd3D/F+dU=9FJ_+@LU8dMTQL&ETDH.)_@DCE.O
<-:6Sa-CCP6H87VP+FQ.:H&4EF0a8R1QMdNOPMDNQKSSJ]@0G:PJEX1=0#(,<_&<
,@)16@RUSXJL3D#a=6HEe@H0DLS<Z?6Q2F42a-#<c)g8G->Z\RKd&60(P<O(UK>S
3<.EJIS^?)&SB3MEOK>G+^ZC6MU#H<1YV4HeQEVBD77&JXL@<94e1/IKH-:,+L\c
_f1:#,,aD/DHUU\^2UVVWFEG(EfSM?4-Y[(A.FKWFFT9d=_Q#>]JME_4C26bRdCL
[g>ZB,T2Z>).\)8^P(LY4]:V--8HI3D@-/b)3&&5\;ZM[]E.<d:D=Dd;g(EeI-:H
7ecLAUfJ)bPdCM9;@M[c3E^\2=0&T_5fP[\LD:BZ#fL#SESD1cE&),_FN6EKJaM^
:[#2+SUE6?=E68#R?(<HZ&9N6^S@])63K5.VAdE.\CXG270f]Lcg0fR1YN;Kf4HR
I??JC]_Y6eR-=3)[Z[GU,aI1;eP<.6;PY;FdUO7cUQD8U-(W&bDbaXV9N?)C[,\>
_0HX9]Zf3:e3NA6O,KXH\=Z]T@T(+U1-b@186W1>g109gVM59J1W&Y/0(P_>a>bG
998M\38,93Da^#bb#Q4=QaJ]6:TC0\dARF/513:+Fg6[]H#IFJ?ZZ.-Y3f>I^K^e
X96;8]_4T].b_Y;c7cALUP44=N-N=U#00S:_@1R6V@0HUDPK:L4QVfcI<<?2W-<0
2Re81NcDVa=AWX(80T;YX36-b=IMda<-:C^(&#:YcU5BLJg&/<L)1-S&#C)P^S?K
(SRPDFC5>c/e6g(DZ>L2XN-699dUV>c<JAA,ITd9eO2PRK(TS1R>)(;\ZXQ)^^92
LH<P/#bX-LQ3U9;6Lb:@6DTbBTC<&_[GBXHN);^MLH;dg=#-9VQ&e/N29g(R=/R9
/Pcg:@J7K-J(VBNb:32T4Z2_2VJPCLaI0.9469dAg;J:4@@=,TZSU(DJJ_)VX;?8
0L9;8<VQ([\EPE,:&<B>N.H2G1(4YIS9FFZK2]b77ZU;55&=NUR>#V4<U^F6GNf+
cRT_TA/.4_Q@H50Ec_K[PUP?LU##RJLK-53Q7cMYV.P:#<<S?dd:0Q1)bT?Vfc7-
\LUggdc^HTD_>K8eG5Bd<6K:;e+9Tf8eR?dB,f3)N>W[5D\;9Xa2[c+14dQ4+FUL
CDYfMS:<Z=\3e91&H^HPFe<X<YIbQVH/FbLV3^]=-fV(:),FQ7g?GFc(W?I(Q&VI
CTW6SEeMF5^4U-.,CP23c_g+PYZO]T24:BZQWL1IEODV]P13-/BHd&Y2ae[&][/.
c(8c@ga41E+Y2bH+610(Y6cFD(OLT&^Z),d6g[)UND9c@OJLW.2f5BGZ5Q5HEZ7H
7>ScX4BHKT8dR>I(6\;GV5D8b0PR2DC&K@_B@?cLJ-F31.HfMf#I=+((gWWT\c+d
2^QOWH-LBaPI,7(4.dG00(ZH@:HW=8C2WcUc(<(]/J6<ZDBITNGZeI,B(eE85MAf
\M\M]\D^FfG5_=9CLJf^&b_);#<I3P2X&d1P+I)R<U>&g,\)/-&F(1a[361F;W)0
0gJLbgB62X#VfN@;SaA.@F6X;-W<=8J<4ESO&2RX&W\aAOVL@+EN>L6FAZ&><@Z,
I]VC)SWTPL=KGBH;.&I9+NI0YFKU7/I.4TP9Z8cL^#fBZ5;WB0-&PfDA:MT);If5
-ZHe(WJ2@47\VI9\Le=Cd8ZX\AdJR]U;3a^&>@L=Z<ZSVF\f6V)=0FH0gE,L-G.4
_J:?\A,;9&-H\<7@PNP(D6XQ1?IKe>=D:HFJ2M>O((bA1g9WFN2#=:2ZVTZVIa1c
[:?;?+-1_I:@.(8;]0_5)<I9?#._[f_S^?I&[e_LabY=V9]_c2YN1>2<@YOR[?K6
^TKc5@H<Ld,1B&gPK8X@LD?87/BVcBg<JQ;P&<T7#ZT3,#A]T1gS0OLGSV/6FQU<
;9D[QY-P,^f(H5_H6)c0Z?(8=(2bQ(e><e7;\?+5>bg2MK^cV<2Ea)-:?F^<e.O[
6D^Vbd3VLHVOBO01bNQ^;@D55I)E6B9@R0a8g(=a9X<gV7g:<F<KHg9F]C-c-C<;
-WV>Dff#@eY:MSI2PB4NL.P^?X]ggOWPZOZRLbH+#4/L/6TN5/?;c+dSNU&7.JGf
AYagC=7)E)7\BaQcWM^0P3>RKKMN0/U-]?PBe_LH?T9dMNbP+UJf+_UA)fE\E1:]
-J1??D29a4fUQAJ1(U)1<ZHG?<?K.ZbY_+c-;Oc_CAZ+-U(<PBLbFAD8G))A>A^0
P?C[RM<MecVeLVK(R_J-7YX?OE^cR>4UIBe1b]/([;/2PH2=GbX;U<M#@[<X]8cX
^)(^0.UeR+e;ESL+QVgH9=23>.;dBBg-/S]];E7M2X^N^6O1=)YP3I0?_5G1Y)&#
4OYedaPd17&U>/((L>&C^1F_YJDZ@<d8B/N4S=5VZ[]6B3UJQAIBIX0CLO[=R\;8
;X2281VZ9JTL36WD3JAf(U1WGCST,1>/8O7#G>T:28.#P<;0\A3:A/ad_K<aaG/K
-E+WF;S#ED_;V5Qa5D[[@M9P\3^1&@:8fD896K+&/4gR#E-;P565\\^PFACMaCU@
^W3,)TA4[^&_NGE53b&/2]YPZMDITAFNYJc;1NVM\C^MIZUSRH6Z<g<[35PXBIc_
6\CS2aLYWfgBeR:0R<8-+TO3==T?/41eL4U)6FYg]R[<:Xd04)S_GM0A+5?44PTa
-I#8_af.4<[0BS[X&:M[g5:MXV6OEaFa3EgC-a<)Pg>?YK9]I?MT)L&.6ga0Rb_2
JS&;]F/H)GM#-O/a)_7/[N-CJA;>f/e.a#=?R^\G]ALQQ[)EfY_F#XY9Sb;BK+@2
9?I#Z8YQ;>/UX6&&\36<W@bQcPA;=TPRBDS;5BVISOH1&;SF7aA,84#gBT6V.Mf4
[R[6_UM0FH#6V_,DEG2g2L<X_AUDJ-9a_Yb3f]2MSL:@#1[KaA(YEVR#<T=Zb\MV
F9;;#H5/cc17XB-M3O63,DS+NT7<W)5b;=SE#dA<0C-.4-&PZJ&<U66U:)LO22g;
gaA\R)cX/SXc+deAAW@)7KIf(>E:/=9N@\#c35H?2@.f4#bFC9I?bKJ=DZ<30<1E
ZVaL-b8\VQ5KI1>.:6fFGg1SE+2gFQF^9#?\QZ;?4b]d\H6e9c]^BI+.,BZU\>XO
&Y-=0]47c6/L(eBEVHbg<B>/D2DM/I?0Qc.6([?W8A@P&A#9PR9RV(M@PGO40?Q4
f26A^A[)&W5J]6W[a)\c[9\L:UK=NKc@L=PSUN9;),QK8+RY7f<X^Y^KWZ5U6]C]
&#>_]TZR342XL9IKS7QE8XV;6+M=g.67T,RU:FBK7e9,=OB:De=PB7K=QB2;cAS<
Q_/@BBSE_A>E.;eU_QE[L0__KAN;f<#9SC<?CY--;,F2UAQfK2X7cVE?4+3BG1.e
OEG@X.B&W>Z&#@U/I1OJFKFF]L>-T]?BGb^74SY<6HRKaBXC[5#JC(#M:3TPG?J<
#UF/g;MR<Oe\YD^:OVT?Ue@H,-<JM,HDbZI[8]:>N04T2Q)dH[MZK91KWDH8F,X6
G#C5#3eF1S;=?dR#D.geN[Z6)8+>.Ad\#YWd9M@LMOWBB6Z9_9g>K/V=eQKd?2cS
@5V/.KU2)<A>FN4c/?Z@X38,MXAb_/-<-6+RQB[;N0bAH3L_;(8cAU,97;^;=a-K
9)@,0#L6K:4WAW=0b3b&2WM_SL1aU&NE#dfgKWg8D_7F(0+a5<JKC-4baN=]\(G;
cY@4=L0@QNdKT2U[9_DSag774_&@U^S+a]GF(#</4>+Q+V1Dbf;N\>KML/-DH4GF
X]/_Y;a/?#EG)#WfbO66&+L08IQ+^-WQ_AbJI/O<aC8F/ZG^S@84PaE3Q<2YU?59
61X#L45<)[D9Zc1gI1gbE5SVc?7?HF,BB_P3=&3^1Qf5-]N:NZ=\>TK]/MXVM+[_
[/II=0::QR0\I&FDD-<H6L:>Q(b/7&5H<2/MPWKfCYPc5\<WC(TF4f8M+OE6,50e
^+J8:WF0caMd/IL0+Od;TR.A0N36<GV4?\<S(KN36]I<d]))]RX)8B<a66QMY:W)
3#VO45g1,CBdg21XB]M#]KZ(>=K@2CdW<1fZQEAO^e+bSM#U[_b7OTdAP+,B.KI/
2>Lb8dF_;_<7FH093g-g[?+.a]-GXcFQ50g;@#C75@#936EYL2.aU5Of1Zd9LO+0
:c3M&AW0DNUT969GTJeW0C[ZbCF>,NJ#)d@Y3BMFAPU-,fW9Ib\VN)7Q;@f[e2(b
#T<M>=^W.AH&AE.1,)#-=5,V_4+,30aW?6PCXYS\C/TS9DF;2LQTfg=[FScL3,&7
C--DAY[F>_[3,P-U;QUCfU[(f4e+TWI_dH;@7?RB@ZGTf+<]6P9Ka2gK<>KFM]YY
b0CBX=:L=2O1/D>(U,JJ2JE9bD:5[GR+dP1&Z07NCJRPHVH7VNHR0OEUE??;1b+4
9aS<d4G=e9P_SK5LCVX@YV4A176#U_3V/6/_B99/PSQDW>bLIX(_Ca\HQN2a?]B5
+;3SVbF2Q\\FD@8a(O]KD+.Ke;2SA;U(K@W-OL/^80YY(:OE)Bg6b]NS1ZcVK##K
,.<KdbeHg8XF9[<X_AJ(_XW/C7[RVJ8.ac8Y2Y^N/1Y?1YS.gI3FeK7Z:(R4UV^G
c_O02P1C/CDcS>U9=1#MFMBO)4^+,Z<ObB<eRVSL]0-GeQ3a^S&EUQYc:dg7UaE[
4c\_UTY4/A&g/N:8CXc+>J#Qc^??O5)5OX?Be@POcUTXD<=FeIYZ+>Q<I,,I,+QY
UFJR3W5^:dSgUU,-G-(<V<;fb/P5O_&C^R1;Ec\CDUEJBX[5/R:(]A[N(g1,,>R^
J@4C_9KZI3:AQBJ2]M,BggJ)]&CG#JUQO3J\3_DD9fAJ;[964g?cG_/P:WF<Becf
f,WJcHI>dVf)1SQK^5c<S6UJ5;>dTI)S3-29aRg<J93F]cNQQ\fK)eQYHB@eUJV?
^\Ba)g+[2U4:K0L7XeNVX6f5Q+P<E]dcFQd.WO35>Q207dNT<D.,0J+aBF=/40?B
.Q>Y&MCK@Qe>/cbRPc/\B5?FQ(QUe-6#?[AZ-+TJ4@Y,?b[M];6&XH@?d&.g95]0
EdObAV6TT/DCe@<?-(-@=JTEXFJ4cC+H(MG,?7PSaP1A[46<:F&FR,/L08Ta#S(_
0AFI#NbF(cR0<f+:CeCe.Oe?>VcY#_CZPdeKBbUC(#M:B_I@I=,^RATO#4:;;(Pe
DbZ6>g-5X9d<J_TcV3LWO3R30RCW4>a2_f@T?\@]Q<XWe.9:10dX:SYc<>bU4W,&
1Ge3bK?IWQgd04e,U_^<56AC;)_PbHPXFPCKKQ6GKZ,6,B&0\QL@]<2c;9b(S(NR
DF3O@GL&</XT6cO.3]2KNB>B/UJT.IXNf7X>d)bC)g;ZfGRP8M/fMBE6.d#?(=(C
]@(cE39,Le)1a0V[G]9^,Vba3gA[0B[T^YVK9R(e\cU>LVJeN:UG=<LHV(43A:=R
<7NV5;4TPEdd;(,>&g2#eg6>.82Jb<bT?2#[\1+^FPgGY(U&e9(:NVWYZe#]aJ7]
J@9YEX8)03-I@2V86=1EY?e\<aBC]eG5T..W(9HCX8F.E;g0b2WHMK>b&N9Ve6OM
7-;?Z9#3TLA7<@Ef?#Fd9SWH^&V\A/D-[I/UWFB]<.X7GPR^bebaZWB,6a>);4+D
H/?3\34OBNOOX?V[TD>a#7IC0UIAO0N8;g)1cg-]9gW8O>NWgHF),Bcd>D4eF8C1
a[&-,eW1dS,@HMSd@3HU)OL-\?K_V&SQ3Y,bO,Q55fP#C+[?&_V&OI=G1E@KLH#4
WS-G3I(fI8GL>2I>3cDdHb<JVG57R#(QP8W)4Z^TVJ8Z95>@,g>H,4BS.PY90eO)
D;90cAAa03:Xa(GT:3]EcR5=91N</:N_9(dS>,E=5;#@Fb)HN]<Ue57_+1>5Y#2d
d;@AE3(@)^8<OOPK1:Pc_B<KQY-XDd3<B7B+-ZEAFB#SG,@&1e2cGA#4N38OV]_c
]KVL.&5]Y(9DD/.,02RB.34MNHBU)<[]8XQfOTVWcDM/gSE1?W?g45F63M>6Ze)4
FOa6\3;E;gO^>-20F1F;MN9/KG+2@P-fY-PadU3#;@5Q+-8b.DZ:LAKXe^SSL;.7
[>;,JX@ELS;G]44RJ1E<VC58]I>DUJS#FV8HV/cWG^Zb&LPPA[MDg_&,W#-W,::/
LIc6DgF1cQ?PH3XbYUO??Fb_dA&C6^P+C48,:0Ua80,E^UDTF4^?P6<e9HgH-H>a
+eBL<39M@gLIJ<-@daO(3cW)G8=EC0CM2>-Q,H4SB+f8(5a]Z#9bU,@]<CVKIT)Z
ZL9G@X?G&BEBVO?SVVTJ;&MFUA___/8,^bU8()=:00#R5WSUBZ)7RM47U2_CJ3M5
U=G#QeRR#;_N^UWbI\^g)X+:H@]dB)A_2;V/7Xg0Gg6\4WN64AMaE4XYRJ)f4_JS
(E,(_E[,M/7BRKcIS[1#D06<,#3Z<EE(#=QWZ4>HE)<,0>-K.gZ)D_>I9WP\TF>O
<>c&/4AG>,(6(gf?d<:;I(>);0R:00,Pdb^1/QCCU5/;RE@KC<D+>^OZ+ZAA(A^a
<+[U7d04L0MSd?G,)gV]-Of+03IFO2HFCT&[gN-QFQW+UQJ1_,6(_TXIO\31]E\M
OP]K.X\:82ZJ@VQ;3WDZ=J)?#1\2NM)BXG@^[_-.d^J)VO0)GM=5ERUJ[Eg[N(@]
[>6U#^Z1LW0&=S39,FVgNd0J[.-FEK&L0fK3gDVAe?a8\fGPc\JFU-2E7b,A?.\L
O<^4?_EHFMB-7B4@8+4<a4\gO;f@I&^BX^&.Y8c\;+4+PEH4Q(_#M5R\.2:1gb-X
T>9+C]S0<V@JA+f2_WUe,>J/)N8>W:=fNLIOO.f,T96^Lgf]6K8+K7;3V?=,Y,-Y
a0[DMBYWd6b,-3[@dORTD&LZ-ZV=?U]AfYIN#\+/CH0K_<F>8>1NZ;8aA@SPJ7f&
4B2+NM&FO0=OZdBTTM63X_2JgU+JO8ICHPeb4<9WS6HKeWDMEcSG_MfMBZC.BLd.
U-MS.dD/J#dP?<7cKLFUAL_DJBM>&/P8+Ra7.=WET3QOGc.?]+)1HF9T7O2M?=]a
0^H86,12GfGad>H:7I_.(.];JQ1KD5,SF=T_a#6XT/<0.U)b_0=.OH91:74#3edA
Y<BDYF(H\JZN9\Ga#3ZfPAXYBOB.>4;=<&BDO>2@I3A#1^C1a@)?MTT^f^PU/CAW
M@>J<7Q&KI-dE^?aF,_E.:O;#,LQV;2eT#A+=d]ON/_&R57.^,7LILB#P]CZEbZ[
,7G1:PR^&dMKG).^F652Y)S]Rc7J-7[SfOIWT]eTV_OSNMQTNF8+R]Fa^[-UI9eA
5H#5#b#L;\0M3FL&,OS(G][IPG@L[H>)R5f-M)J#9gdHUI&(V9WQ]=gJdRIYYU;)
VI\U]Oad,NcCJJLM?1OLQ>YHO7W+#<]8M7Ec0@-V[,gCQ9g1QBe_HS?9KH6?U&eJ
O-O(9#[\7R(^2cE[KNDa^-C)@85NR&-cC5<;:)Wc-9+/NDN2Td]4R/7_UC_0>^KS
BCO>..4UM,]I/E_B6P<.1/P99;2PTSE9U,(L/2FbHGDFe0AP(1[1D9))1,eEVBGc
ARG3Ff[(W/E:PbR\-X\02#8NM2YVIPYfKFFGf\EFaG5GS4B7A[b_Q<J?&3a>8O.F
H94[;+LP0bQW:)G-(E<dB(\1RfXG.M_A:<C&VD<GJTHR])M2Og?E&?=#JT^(FD#5
S>H96dRMSb.6J-7Y[(13<9Z)2Ce[e@PJa(6D8;^gNG3F&,\Y4OXA>II.NOfUC<DD
D\:Q]5Sc6FTFd32Z0)f[SfOGGJ7\7KA6eQ9.P\9LQ@_[M+VBJY&-</ed=,SW3CfT
>PaLT67]8K]J(KCD;=M7L#>(^;Adg5b,&BR9Y+7;cEfE,I(BY9V&\QQFJ?Q.8Od>
c6M(6a#dA2&<a]KOKgXOB8#FgGY.@TY,.T;7V-X_S=:QLC2.OM8gLID6,];5T1AQ
I7L7[cfAfHN)/TVB[<ZPOAf4<_eN][I.E++O.d-L.\EMKV+^Q/S>1.L&-]7FT;.B
Kgdf_I&UA/?bC=P_],EV<bOCQg<R->MP;X-eF@971WA_5=bM@](VbE7E8WX&Fg;O
4B7:#9Z,ZB;c&:U\K.:@[c[5EfeAX4a5AgO&W@QbOgQ>dPdWSc1GT=&T3_R7OdI]
7Q@a^.1X?FW-R6\T_,EJV#>IK,[B3XW/CeG9cEZ@&Dc,JHMfZ5aF6/M_>f(<P<87
)f9>2Y?(7MW>RgD?VZf<3&9L:He]JV-74MERO8S[aS/YAANYVR;F(DI,;3T=a6IH
5(&OT0.LW4E]&]/-[=7.5_JSY)1RWgG12Y;1LM^P\_(K-1G;2D,a5f:f>]05532(
Le4Ce7OE6&S\Q_,579b6FBA2XAV[Ya.K?FNEdNgTJ7TOC;Ie9Q8c4Q-gHdVb](7Y
eU[[-3N^SLX)[5MZFJaE?57JNO_[&_4BNCa+^3_H7^aK85_GIJ#^DL:9H8\A(ZEX
&WUJQ&MC1gTE5c#\ZADDNQG4RM6DD4.5(_ACg&;gb.HP:/7#PK_?P8I(_/&bL&K=
Yg7:7fKG&YRN(06))DBdaDGPAY.:K.7JW)_7K+M5(NPJH;f8?)H(-?=IXBM48V.V
RT]H/b&P1CBV+LT)8:IMLG:H,cc3Y>gN_7KFe6/6CP,J^RHWcF02T/B]KA;fY+\<
2U.Z\4#?5BdBW>O]:+aZS[KE_)Z1=T0=gcbWM):I9GH9S/cQ[MZ2EYE,)0fNJ#f4
b<#bYC4K-FY8I+HDDc90c1Q&Ha9C]W+68KY.+/d]\>ceJ^O4+9NBf&R=7^9+eCLU
=_6F.0Ib:F)cT8QgX8Fb=(39KPV+;5N-AJ7HL>@IUV0O6PfAPYERa+FYX&e8I<K#
+HAdWc2+fN(,#2Y51ZQM1X13XSWT@0]9)2[APPPeRAG,K5B?+9EI,E#ZT?)U&IJd
]eL+=CP_&4JE,#<GB80;)2+gRfM=RR3\JD6E;GB6DG/I=E.@:J8&e#U6@d3eeSB5
;g(bF][A4?:]E\eXY[,#OfT0dDX(D.GE@0E.EXQgROBPg/g6_:URgX5)(U\3KG5L
fFL@RC(B>6D:((M#7eY-^LG6R(D3-bRdg@8VGc9WXACU-XM9eNHfg>;9:LE2N\Z\
Ce.Z.@M..7cB&HMM9/+:28a;4Xf;+fF9-];2&[e8(655.7>]K;5M7,_+]_Y6)e;X
6QV.g_e7VX[X43(_^:-?;Rd^L.PLeDNUY/LHQ=DA>QXCW[O#PU#.4/(CQ@DL+X7#
+5M1?PM1LcBNgNc7agGUZ&X2&e)<#Yf2OFYQTSGLS^[LQ;-FT68YD<>AYZBE?1+)
?4^T8-#OL:PFdD4IQOM,]9?WAWOaI;<MRge8ZUXGB?51K7#.8XK[Qe++H48\PXKL
+@X\YgL9[(1e=65Bb]\N6-^_W/M_Y1G7bD>>WgN);Sc=18.=;^Q\b;=]:RI#>dK>
D@&6G1cV,PBFN^H;_^fO1KZ5OWL=fPPI5:aND4L18Ie+SO+f-OMc_5TQ7[b7X3MF
AQ/eTC;P-#\<54>(1c/BA#LIS0LL_[FR<9Nb=G8RB#b#TT0-B)K=0)-dA:.]:UXE
5?;=A7C^NVO^?Kg(<M<Be[PIJPT9ePTQV)3CTIB1#\W/::QIaP<75&W&M&>FCe=?
PO9&,X:e9ff393S:&N_@g7+I:[Y_b0?aZg,ZQTS8\1H02T^ND9GfWgT,_CQ9,M/Q
@RZc2S&VLG^OJ-a.JN.b62?0<\D>^35QW0:H/-I-\eN,0fS^T(?_N>SY5-C^J;F^
E2G?]d;g.=IJf^>AI-@7fWc-Y&IFP6dWYgRKf:#+Q2M4[=L9Ngf.M]TY]bTF)6MF
2&Zg6d)KB>WGe9_B1X4/eMOXKR-]&=\(SB-I.f40AYYG@H)P0.Eb^FKIFgR^fLfa
DbbG?O2:OB;_;^E^H-PU>b?2V:S1#U^5)B)QG^]J_X3P/&#[K,fS158RP([T=_M0
VGDF[[,B_9#\Aa/9E\N(Qd:3#[W9<TP08YfW[d9A?S]0dd\+e_\I(5BG.@=[]NJ.
e_6/RB2TfX=9\bDD[&H>C5_/g:45F&4PUSLVT278W;2Z)51;=RID1Rc&Q3g>UH>D
dE4:F0X,C5?KQ0P_W^XF@g0D]IQF5M_W0;&L-?@>/E2XY8c011)d(^SG&2EV.d@J
91TfOcSLLf0V,H#@,36@1D&TTbfYYg]__+ZOS?@FcAgA8bYOLU0N7-:O1VEUG,d6
Hd(9,K1eF8^IO+_UE;ZZT.eUbGgXgWfL2^WDK(#15[I?UNGbG^M,7U5SdTH4X1EY
4Z6F76[B/47)<(Fe58D)N9IVc4\SH-)\eV+;+B6+c+I>a.L[adWMUJNbT/7BS=.T
dOg0ReVHeN-RD?1;)Q6IECBL462e3T(UQDgJ;1Z3&WS1:.1J2PDN<.TN<XI7H_X7
4L@633ARAd3Y7=LSdK(93,)^Z8BJR#2dM0PO8H\IEX1]R2H=\e_Y:(Z)<&e5>#8f
-8;ggg/bg18R.OC:FMZE0V)cTJ@9)MZD[]T\JRO)&<&VOAH5A8Y/[75>Jgc+a@6)
MS(O&Q=ZXH-GE>94+J[_S@O/A0W\Sg/<e?X)>FQ2+X\@E.daB/5bZ_+LRT159>:D
)TCcHCMZ#P66&FU_&NR1;cYJKd_;-MVVR.Ae>+K#+PU/6(>+>M#\/E&2MJ\@/3^3
@RUebDL?Y>#\6R1H\YDOBaQM_S0OdL)>UgM15-R4bJC<QA4Z1.F4g:WINIOgGb,2
EXGB,X1HCZYNFH7QL0.^>4IP\.#U5C<K#E/?IZ2EZ[,/T.SY?G_)Q#c^&Cf5QAeV
32dE+cAU+53\f0+PJSFEAZKN-H<;&3Q03U_50XOKCQ[,C[a25Q]d;5F]g5dUO76[
)1<2=Pg_X(4gJ#Za/427IT:e:&J5?\W1R4XDUaNQU/\g2I,2BT/ISL<+g6.D.CEc
L(];3C0-[IT4a59fG=^a49a:>dd,TD1GLg6TI_6_DYAVHMQ))3TC?]>SDW=5Z;eL
b1CB[RaA6CX1\PbC[]=b2@,e,YS8HG@geefPP-/M)Vf8B#ER1[RdH-LBd_Zbb>4d
S:-I@C7cV,&/bDQ3Dbe#3,/eU605.^09(G:_6HC/RR/AL-0ECJf59C(\47.JNC<R
^1)F)C58R/-gCV#eJJ]1E([L80(;<Z9BP^b0,&KP-b0A(Og8.@F&E8#?^>DF#P#+
CQ3>N[f4(:d5TcZLZWd<5(LL:B\(2\[=fDf@;)+H08QW4F8)-(cGJfN,d76N(UFG
Dd34_UL/>(^?X4H;8_L\^@de#ec0@M;e^4]C35]<D]BDa)(,fHZHU3&eLQV0P55>
5f:JG2.Ud?@EVCFG9eU;O6<BaA)C\Vc#VC22+T5O<QY5+SgDfW9.)L+QLACcACT@
f-..0+@c7VS_^d>?21+d<[EV#1(L?C(IJ6/V+AR_&0VG4LcD1X8LT92:8X-&S<YS
_2GD+,0+>12DbP8c,79_-MJcM)7<-72E#YB=JVa?1G6+Xd#&6^YP=>WNT5,,Wd<D
eL?fCEC2SgNT=ZJ0V@Pc.a5=Xb?>eC&Yc]gEa?aIT?NRYWe6:(EX&[+f^KCcGD)L
A0@c-cS#66(;RE#/X1cK^76B=&>?Mdg#0.eI.V>T4JF8HY#Q640/_+HV3Z/TW813
(?aY=2B8:_;Z8=1D2,bd#^PZDH.0LYOVNO?H5@cRV;N[OU,KTD&C(>F2IS)8(P;S
;W=CQ?UP;9d5e@Yd9=N<^b;7RT/ET#]9HC5g++\P^&/II3eK0R\1IZ-gU&EfUY1Y
Mf=O&7Z2=DEa+6Yg(UG2Q2V#dZTb,3KVPT\\._7\cd_d+gGc;2J[XB(&RGHRDdeb
G#-f=+5e<,.I#eVKVeCZHc=CJ34-(,bVFO/,?\HS/I#0:QY@D<)3ff.RY)D82RR(
H0M_Bb2QM3BNZ_gP./2O@8b#3b4YHPIZH+,BDZZ/U9P,da::E7[JRM6MHU(c6S&K
RS.]2]a6CJ1\A_-HQ[.3cedS5]e8?9-14aUZGPe?Y6=/\)gL-^d(7@C6]9647T^a
IC&O,,DU5f80\+(TVU8E@JNZ@-W,3VD,VTG+4gN44\63)(-/0Y;B1V((#_N>:-QJ
E^142Cg-RH#fa-G]6AU(&624@P(QL?NHd,?#5Q-GY8JDgg.[&J@6\<_0DDJ),f5X
IW2d5K&H\&9/W^f=RTS/A>[Z3aba]Gb\HEF/9+3eGU<,UK+(fAK4F62N,DG0:.Tg
g[QO=1;7D2:;gU-TaWe0-;LSeU3>+(YQcMM)<dKWG>fK]1ScFCU>CGM7MRC@&@Z]
93Mc^Ze5:OETY@ZK)C&3XM2c5T2d)5b2Q.&4<^^U=B)#_&eSOd<E5@B@OYR]K,Be
d4J@a--d-<@[=S2+(aT52f[,\Ca(O_e&BfU?4DX,EZ7E\dX<TD4</?9VS7Fd-B4?
AS_S4YVD:Qf9K)&A.G]PH,c.CHG33U(QSV7]D-]FW;2RK73c3&_;K&_3/1L;/4cP
SE_@;\8d0N35F<(#R,EfSC)fe0ca.T7]<dHUWF_aMcYVC9@-AW(B:##5LJ+Qe2[#
[a85B^1<B>cN2>8MI=<NQfUaN=EAQEE-eRba(IO(0[VD0F]b3(W59:-)P_Z:/XDZ
]-2<7]BW7;--UU#A-8Q8&/[f:-U#9/KPZ2<N9=eXY::KWBSW3QJUe<BHc]+@_38J
.=)C?HE0PL:0J-OJW6SE,ccCG;g1BcdCDFIaP;DKA[a2W=@ATRVgc32TSD-Q0gKV
bHW2c/1R\PW.8abI1^RGAc9UJERU\&5][5)]IGK:<DU96XD_f_e2L)\HR;/N#Ta,
U((:,)9<ZHF)OXQRDdYe>K\=VLLD_,DMZ5b[)A\\9)]BZ+HE)@cM&8#T.^_VFYSc
;_VV^c]>+/eT#fJEA.+2:GMdZJ:VKBD5\&d1UKdO>+g;cZ8g8OK+8PM[QQS-M3,6
L^+4Qe-G1BEfU3JR3LMLU7.d.QM&QDSZ5RQ#;c#M&?f(A[Q[NL[4-:A>C=48-J-C
MI4J#+TKKC2SWE\DCe7e2gS_^,:_dN#eG[@Q^fG4U[<Fg5g&R653^2<eQ4L\O[L8
9/KSb@+C/5Bb6F[QNU8-0Zed4=f2]g-Eb-_V[6Q)7EE9ZH-aJ2:\cX=W-G8M-7[b
8.T&=IPG(MCaeF(ABX1J[Kfc>B1U+1L&NNSTYPe<Nc@7)YL:V<dKH-47D[NRfb8P
c=a):(?YE3E\4D+N^U3A.Wg09B(T/8K4I,-HgfU5Sd#WO;_6A]PQ,^#_4Dg5d)UE
E5RYM<P,Q8e_ZMP8:+_GeY22GE5>)R&;RJ=8+BX/4+f\a9=JW;VNfd126bOFRb2=
Y]]]D>MKO(c\1YVYOT6]dT-ZgTT4W#D/)FfJg1A-OI@0>?@g=E,-_c=#PQ-W-AV&
462a>/2F>8&\&/8;A&NN:a=U<-HMN/?8aZ@&R4<g<R,3E))UC(]^,?3U8TQYH_&3
=.IL0d3^fJ=2WQCZ0&ZEd25Z78;#^e+1@HY/eDRO[X:]8.dAeeKBd^/a]N+VddF(
6\7M]&>4.1Z+5;Ca4W\B@S\C-HC[E=GgY>FBaAKN=W.W-\aN<,PRQVeI-M6.J?X#
+MZ&&>2>][29aKII-U>eCHO.?,cS3AaRcY;#&NTV8=JY<a]L@4;75H))X.fK23,V
f9:_)&Be)DaZBU0)Hb2+#O<;DM##fdN0GE/4WaJ,Ld^HRQ_Xf@F<],2e+NffaV:\
;E/PZQ_YA&2ZcO@5I2_O6/C(&NGP4KW2>:^5]]RM.<Z(HH](FU\Q\X;Q,IV9JR=I
7&N#<gV4AGfW1@Y3Q+@STABe^7-#.]+XZ/T_]a^^TQ0=4WTb68(;f?KFU=_Ba0(g
d#e,XgS:=P1D0AY5[,:Y^X+C<ZS2+=1RD(H-<^<;8Z.77;?5[Y,a4&P5J]dPYN[(
6F(W1E);.5:dD+E9\JEff7AAFCcRX_=P?)N7,&M.[VVV=5adUa+@B3R;6XbZL<Se
?f5(PIBd#&KS;L=1Ud<TJ]-QIT=(&,5_F#eVIY8O#-D:,V.f2GeFH.Pb@-22gS8:
:/fISA22Q<AGdBF3F+>fMM_,NC;/AO=CYH4-M9Jd=UFaZG]9X77@YQcTY,4<4D-1
b@[-V>W]aaO?K-S4K)>H;e9.V.D(Q^<.DEJ94:KF67_=&_4.F8&:6M/7>/1QB1^U
.2O/)eK+SMadDANdHW+<YFa,0^E3cXP6OW)fY6Z.44JI&6.IA5@9LbR@Fe@g->W:
))IF_T)X@]1\RCf]I]Wf3>F28@L+I+KBS)GUA-_Ef+_^P(G/PE^Q2>.;5P9J8U[6
cO<.\#G:Y1g0e;U0O=NX82&aS(X/\HE5M\fP[=J62#\Ef3Ub.KX,9^33.,#F^Ja=
FO14f@GW@5;P+ETS=D@QT[J4+)cdc#c5+g3XRK<J)MK=QE.^Y[)9Q?QS61TW=D?[
d_JT0(6-E<NK:_>T/M<3d<f+&gbO64HCQ,\598_,Jg@I7300S36bb2HS8Q=7JB66
.Ee#<JXWX^15GT(5T(->eaaZS<A12,OUdg8+9<KL47V?F]G9@[^T8TdfSAb?3DF9
L;V0ZM:2H@+48U^cbGgGc47P,Y.?,_,Kd^\_\PXDHQQO/4bQdbVf)<L<+JWH(eA+
9d-D&5U]^Q-URVMR5gdPBP6?\5)ER3E((HR:N]_gP+VSC[NfF=eE7aXId<#0fg89
Dc8Ia]8RS0<(G4=L=(Ne74=\a2WPI>7AXc-dW/-@eL,-T&R5Q1gcf<;R?#E?#U?H
J]V4W^]S&H3XP74&fD=L>EC;ID+aRY4X0,6HO_cPYTd0&/1R<5:_e^)8S48,F]Z-
X>dXZSSaS2fT;5#C,Ng_d=GcAOKg>b>S(4M\SbSH]1CS.Wc6-47f0X^TIBR_.HWa
DXe1)2K5Q9aAEFQEP(8IIRG^?BQCY[4^1UAd,YMPLTa/]CfKRL6<GO--=Qb9?Yce
&=>W=39#IS>:)<gHHV&@74^1T(UCUZ]KO5QQGP96+B2S9]R_-1W6IY0<SNgTBfX8
fDQ>GQ6ZD=@Nc>)2\Uea\<<A5,b2E7-d.)8/K9VGB(F5L^VK;V1HT@T6W&C;8VMZ
2I.c[;(7=4e/#(DL>)]FS0gcG=)(g;HLX88C#HP,/_T,+/@S7O5I:fgA/e(D#c8[
QcA0#b&2HX>B>6<>-17Ka06_Ig&K/Gb&&P)dMg4>:SaF&E=X-A:d<K5:F>>229-V
.S_L6(#?&TW,2fedC(T<(Y;JRAa0IKO2caL/473VIQRXS.,UVVBf^V/G270dd.f.
N21J9[M]HUL@S7-.VD6&BM6f@0ACY<Ta;Hg]:\Z^?LV[?Y,[a8LF2&&SWM>2TV2)
d_MSRYX1/SZ2^>Sd5=1AM09HK&=-GYd/+9+FeLYfAJ_4=a;X:R#8S#QV<_P_0]R=
a.f:Z#KEUA;0CUC@fB-G_^K(_g<<YZ7OY,HBDA2WP/HMW.]Q2,c;LcJK4bX]Lf#I
6F0ESSM>:aG#GQ_Y:[^-G4A5b-V)K@cgKQUDAE_AA\DIeC>]JfaWa^2SPK..d&@#
<QK6-f>+20:XWBEF5E:]]X[[F)-;HI.gTa<F>6N3d?F(Oe(b.-PEO[()E4:cdBOY
GGGV:\+[_2fZe&<?R4H=67I+\F^K8X#BS6YII/VEeOF8HF>E&>NLU1.WUF]eN?ZG
fMTHGc7.HVA=0SU;Ac<A^H49.SD3M^(<[U4I?#,W9T_=-IdHfMZF[/G]W+\T5LQ1
-6ROQ=94W/+/8@d]FX,JXN>97CRAB]D9P238(dW6dM8V,fSR1<KT3-7bV=AX=?1R
0I+GIHVCA9)^E:T?YO?IY^UCeb.;9,R)c2A=2Q[XWcaK?EVaY=:0+YLH_[1&&:0G
FID105VY@XF_G2QL2dC\8^8FA)eLdDg=aB-SJC(00cDdM,-V9TF#67a&SHdO<P-F
GUc_;.FBUHNg+HM-(N7<0V]@C\D0QU;2<&C]b+T;cII;CWK3?16ANabc&]]4@3CA
(/D_N_^I?]-URa.<?FKSERaGN:Gb_?9GJJcFa_d=bXCUP-3QW[SM4DM;4Q#bCdb#
?VG4D+\MYL5).Z;efR+d=/,;MIBBa>Q9/JA,,)eE(^&R6Y,-8+:X,QCLV1=R-]Qf
Y<aEg6#F)X9ARKT6cYMd62g(3MPMQ;f\L3,aU2FF>RV[&0/&:a0&FRE-0d7ScgV,
+/Ma?,3=+C7]eD_-N@\;/eYOTWYX1:RER\:)@<:OWcA][dAYVMC4J#XB8:G2(=9d
&]Y]e=1)7\-_3<2N@/,^9+0)0/_cPca69f?DecRNa](cF+;O(<XO=7)gQ4gadNc0
bD,O:>.].40T4YE8A1_QZ,A+6DF71IO,G/V#bD7)?FP[U-/(d]>5R-MP8-2Lb:MQ
eeU3:6:?_e:/3-V>.Z.-T-AO?#@(WY+;F7d9\Q_9M>0g6.bU_T<K3.8LM.ND3]B:
6_\.=8c/\HHJLS0780_XUY8OQ9[HO/R9F?AWU?1-MTP)3Q7R0)FFWAT.Y_=T=VG?
,+C328AUG;E=5\JdfYg>284QH;-M>2AeQE7B46=BEb?2bW0#6LEBU@5MB;VJ-\1Z
<,f[PR5V0S-bV:\\A^g</P,[,?N[&7^DD6cI5&(/fY-Z7>P/&CE0aI&P_64Zb=LE
-?>-_6#P^>>.I^F]\ZV[N/MUNLW=Wc;J#aQGaMJ[8(L;d[>4#7+6_DO>0(Ob0S=L
c313105S[7.Q\4I41:g,C@->^[DJFF<.4J.T]YIV6+1dE3bFIS[-#C;JgI[2Rc/W
X1L.EVE[5B]Lc)HgL\;)XCAM@5TL)7WJI2BG;A\&(R/4^K/S.P>=J[2fPKUQ#5PE
R=YIH#dQbA)eX+1V^_3eN,1K82/0&=,^6,\?_Y_N/28EYDC2>5Z@<R)-^Eb2XP:R
7@P+-I6bWbJ8;[T@;-8.M7dd@?1#J+\1.4ATNLM/dF]A:=Z<4GN<e]30T,O:GCde
\/6()b:G>SWEDWZ;8]6Td:1#GQSUUKD/0=Z0MYX^_NWS2)U@QB3?8DZ&@.5]S@RU
PH+?8:8^cAUTG-SK@\:JU,XYB\)0FR3C-CIO[>GMT)JG]:#fO.D-_G.a95W3e3QI
@^-LDgf.@9<(OZ@+YR<\@ZKE_7XA=g>MJ9_9W-X0@1@F.]_7WQUV-BAZG2+Z,Z+\
-RW1deCSf;R)-OHb[DBO3@8MEF\B5d)4,18;4IGG/SVfdDXFB#^P)G@.=X[T\E#R
/=QDN=UK9E0fYD^UY)DXNVUH8[/]Kb)AF+G]A2fDeIJCECL#0Z=].ELXLd)HB2K>
?#&O3(3)LVd6KBa^+8@TfWU:d7?^\VCJeTf,DUgQ9\7W1HLY]VNHK_WTGA?JU2#M
AF8WJGF_=CaYb2PM2IFd96,fL9C<WcJ-?4Tg\[-KP;c^W]Eb7O/;?.U#dCLLX1[/
36(I-HJPU?Y0;#R@dA+KKV[5)UcQ(aJ;MM.EI7?c:Y@2ZJSUf&:#7J#OcfX3\Mb=
8GXP/R.#5C<0aa7_<1TS61eSJ.MEPYM9Xccf)WcEZK0IJdK&4cWaH[-e3&5:1O+P
BSC1gCef#2?DRY1aWC.?_@O6L;JX4/4CH;3(WgagN-M05>Z6?^b=_I5<BZ+LDE,(
5P_8_b4K9=VGbG6e(5O77V0^0]RH0gQeaFGQ1_,&XYYbCA#>e<X86K^ETL/Z/9UC
B;(M4=PI3TU0C1T+>L9R2>Jd.;Vf44L7Ad;\ZgOK1:;.;Y#_V4a5M4a,[2.?./9P
BdZINa5K.KVHWYME8ZCP_)b;F>0>@H.@E5/).CA(:ZFW9)4](WS_<[Y=,O>cdA;1
GN]7U6&<-ABFJ:E&HgcL1_21[^.MCAIV2PI0Mbg>7.BFWM=T0]/F)]YMI&?L]gRH
5BFSVH1F3,U252Z)JLT3I<_6X6L3]MKHb^EH.]P=@Fb&+IE>#@016Gf;XK>ERY8L
P=_S7Ff8A/aS+=8SZ^7VHBU&.<&JS[6BHZd40D;d/3_BS=ZTQPL^KW;0Y96V.e^-
e)^_K+(40N(<JY2@[f&EQP^I?WUYWe4M<,=+5=f8#I-;.DEaRIS4=JD8[^-0:XGT
g-aGL3,6AfcDK/+:bQdOQRY6COT4R?Dcg4b-U9ISfbJHFTHEDdON.6Q=9QfC/XQ7
21\EX@T0WVM>f,W?>CE5Z><C)RJeQ4:>W@-B-5g:4<b#LURQJRG_20c\4.#)3/1;
bUNc\M6[XI.BRNE4,Kg:fdA\V@KZTZ=YX<[O><>7^3A-1IV90RE#OUJX/S/F:L#V
E//_6X?;,E,<]H]AB8RC),6g)/YgZ653=WVS46L/0\#<JT^M@7?63/[@-5fC;fXU
D96#SU.TLLI\A/1CUGQAae]Qd@g;bB,^[dR@/O;Cg3XR^#,.N?,.D201bYE9<-HS
_b31Q_,+Q]UF#][+6Z&B9<<U+fa7YP<U0#R]I+eF9B>)I(^YgI)7:=Y64NBJ]F^X
6,KC1,2Z1TPQ4FD=3]V(-?4Og#\eWJ:><D[T++(P;D<8O7.0,>QO<Hc>352FeBUA
Y_77OD5-U[LOaO_-Z^I]cK#\^-#7b&_1_g9I)?PVWg,MPYP1adFT]d:bc_IO5+^A
;Y&8:ZeQ.eg=;HH#S_2/,ADX9JJ35T^=MXG?J\0aP+VBG\5P0L(+.b,V5\Gb;.gW
]QD5#E>BR/2E^KLM_Ic1C0cgR)+M-9bE6CX#d,EJc@M=@2R2>?E=PD=BA]Y)\K\V
N_6_21]<eI>0]a/@\6GAbPR3VaX]gOQA_Rf9[0T\Q0c<K49ZP(^?5R9QU7CEATcB
YS:HEaB<Yf+7_cc?;T.\KXcV>[8926)/Y,XgMH0#B<((Ag@ID28PVbfSa8:?ZW23
]GY@\EBaT0\N.X-7Fg(Qd8P]b:6Rf+9\S@OY?K6:8fY,JWVP):2(X1@_8^^>SB[/
_b9RFYc3gU&T766cD=PVc>^/J7K:^IWC./QH1V#CB>2N4D871aG2PIcLI#4U:22^
3QK0_MK3T;SDUCCQM[faG/CUg1e,M8#DQSY&L3N?e0O&7Of#AA6VU;=8N<#_-6Ia
da5R8V+NZ>;,CgZZb?=Mb+GZ1NOfI5P[J;O#PdEI3/=2Sa)]MK?-LB[ZX<A8E7a/
0-dKREcgO5GgW[gP1XL611If^(CAc&781<C6[M,)d20_?8Q3,2BUW?@[Lc?\P=T)
\^DC-J9c;70R1P(Nc1=0BJ>&6L;g7&0>7a(1Xa^06OfGQP4AdAN-5:d#NN@+g\RK
3#Ea>DdCKU<cd@EN#5f@/0OfOd5a1DN7G;N3#V,b)BZUMCaADgAaJ1,,1_V_&WeC
PUa&6O1/a?=WDKX[&T0&;DDR=;?<<3Z73?7TS-aS:UQIH4_P]b\G#RP7bE;7RL.]
?-CQb7cBE^?ZGRRc8/^?<?geZB\FXe>geNP_C&&AJL>7_]da]1_,;[?Y]XNdV=BD
NNe_YRVW#4@;1/MMPf]?_@VPAI.a8VLFRe1J#82MF;_:<,V,,_5,)d:<T]N)ISXL
4&e,[P[\HfH.,J]G>0a6K8&G/fQCY]HJQcRXaU@0?@<3N-Ce<R6U+6Ke@;KYX)EZ
R5#c2W12EAgWM2>,_#N5?^JPJ]bBPC,BI(RG(J_aA=D-]]HQP&3Tg&>D9<^U@HU]
5Rc#>Q2a88@/dORQRLA>O@.L;GZU^Oa[[QB-S@(+&#L(DG54A])^[OCFG4]M#HI_
_E8EWRgKQ1H+33D:4\#,CDP>NELf5@YeV,H+fZ\1J9_gR5a[H.U.3-e^0]SO,@]Y
V9L_+g64S,1BM/Xc6Q1,=)eSP4T>>MC1E<:+TXFAR)DeTdW3SX/57bYV.Z&&e1g&
&+1NC_/LA[[<\TOH0&Fa>]NR[9AGX2gV[5:PaTY]Y>gf2.:)4X>F.OM/YDS7GS&G
JTYO8[X5^:,c?B)YL\W6_B(^FWR+X2\Z,UA7MG=d7fM?L1bOKKUGN;P=3dQS3c#V
)HQUANNAJ@5-C>4EXb_Z27K?^IQYAI4_1#FL5>S5^??_./Oe-7#&]1IZaW)+X_eF
K(=U;L@7GJB6BUNN6U?#_-G\U7;T^X>g_K:A(^P/=32A1Z0bU1GN//b^S-Q+.DdE
DA9?./3b:PV5EZW^][EbA<#\^:.Q,>UR5CXf:--4O0OgfN.@7Gc.f_K/36S>[6(.
g+8])Q8a2ZTb#<[De#OYb^FVBT/X<RGfUc^@E2=K@RX1N0^S/.TdS^0=?RUPN,)<
B9?Q-NN+e)>LN.bBDB-SKSaUfH\3H.RLJ><ZLCT(),1X,#D]5d_R>_+3g@Q2VO]Q
N:W@;\JKBA=#G^X?f=A?KPPZW<@(ADf279YC_78g74HD(FRTdM.8IA6-\8_D4R/J
UH1U:cc:)NEgU]gb4,=6>3Ae?2??JS2U;-IGBN<_[/W0JXgM2K>&,R(A]E5_YEeD
L@KL)f;1c<86IBZ.U]H3VZ-_;K=/W@c+,aD<B6WHceE0\Gcgga4IIJ#H-gWHW0@2
VaPF^]gMfU6R801a6#c4/CM6<EMbR[df^(UJe\K2YeMLBR3Cd.K3EU,L5_=a6Q-#
ZX/b[\2\6(8+9@>:7-YQC<_?c_EHReQD:LL(?Lg;F+eZ>),>#aLE(7)C-OV9>X16
E:#N?BZ/fJ0D&O#[7S6JAF7C&bPgXLNIcJ,D]d,afA[/4EPIe=LJBRNEY0)<WL20
-]b^C/V5KC;5U&U./U?Y9RCQ_e9Uc:PcFAU5F5.5<UeZ3ZGP?281M2OFFc,d+EeZ
B;]cO]8GL[B@1b+.fJAC=S.FL]2RAR/0BALM2?1PA<3?I\<f_JP20=U4WIN>gG)d
MRQfc7@I<Hf>XTa8D&ZE/I3G]X3^>KPEeV;<c:c/5FW92M1+@?g@[YLG/e6BB60=
6fc2ZDCd.E+/9d@6@6>J>CB01N4[eX_NJ7=Vb0T3CW.TRK^0WSOQJ0YB^]C,KcQ_
82G:ENJ78S.WaW[KB-;3#&-H66)HeCXQ#>\PXB1-B))fe_BH6(d^+PWMJF<.34?7
+8Bg^Ta[B8JY3Oef]&HZ;d\Z-7-6>2.N-P1XNBO\:0JZKg0)-&4V)e6TMc_Z7@[-
:0#RXL1)MLC6=:dfeZEI(Y[R(_E=Ma.(FdH>>#+4)2#:V]?028//Z2fF&,8?IQAg
F&7X^K7WJBW3IZN/SQXd+[L7gD<-_HKP9F1/LL]ZIEdZVbPALH8K,T+G0a^V<a\K
CM/(2O0(7SMY)<2Id=H<1=QJEC.RS]@EgbY]fS7T&30:I=f>+1?<CL\42BA2aGRF
d:\OEdB8?^WQB/@b94J5d]:JPG@3X7(C^O4-G&K96>L>F#<Y)f01c=C>O]W>Zd[Q
b/N7]3COC=PJcZe(QXDaQ2<?L@TAIQg4NbZUf^0U+cK55.bP50FC5>H6:--OgN(P
L_3^KOeAab)/:5:,QGVYY51cF@P7@_cDR1W3]L;IW7g\N3(;E1-P07J>7^G_<S25
<VC^Jf@=9XMVD.L?^A(R^-b3QeY#\^gDD:Lf]/^D^QR-c[M@8V+(3f-F#Qg_S^?E
:X47U#;[/)X5ZKRG+[P=A);Jf(I(XGPR@F\@TRg_Ea5Y@6Y0X8EA_9L_T[fIV21Y
g\L/3NSJ0D7M9e]<^R2WOY4N@bDQ8NY-P)U.5#?dEDgXT:#[_@f(KTbK,NY_1bUF
4dgd2?++<JW-)MSb_V7-BcR@fVBWAG>[Z(:d^-0G46O4<)EZKNH2b])+NUPP]Ub4
YfF492JLFPW7&M>LYWCJD.6,<ID?K1SZS^>/F]Z._B^&4S?@2Z@5\5_P(U+=\^H0
:_W-T;+7bTQPHf&P1Y[MY@U?TR@,\_GU3@5eXT6.6H(?L>/?:b@8+???I(6E^];D
e-F8BO1RQ7+6fc4^HPd;g_HZ=;1COaU3C7OEWN^G8J5a&-HL?7#D)f+gU9#c9R.-
E_).bTN>Pf5)CbJJ2Ddc<9aV)Q7TG&OS.IRF1e9V.B+CD),\g1ePdYM7W?f6U#5X
+W&Cb(W\NKIee[Y#ZM+,>=g_W=/UE,1O<=eU6L1T0.>-e=WB,8@,=b/1##N&Df@&
V&W?TBbE?cWNF#,C5&(fXT(0g.((JS/]aHSNIKgF0YPSFfYbU3Egc765g<.a7S^=
G#4gbgE@(AI?faME1[=bC)W.2HKQ6EY5J6QBe#0]1eDd:DFBHH1./d;&I);OQTPQ
cRT(JNg&62QeJc8-fN/JQ4_a+CXZJd@-;9\=IAf<V6F:+>>D&Da[GUT+B8/eb3LI
C7f?KEE@[a/X+:XC^[)\98;5WIG)5/^4&F6LPSKU\CL/M5=AU+@-Z<C57#;JP8,#
@O=?cfVO.99QHG\Y6P#&-<e+85D2/\O0-EQ9TGY3efg)):<]7&7.e3W/fZTZ6^f_
bF<PbBLWVL(K^KH+;3(X62ZIRX5:TGb[6YF#=HD?\S@/UH;6Tc^NGQH)#C4b9?SZ
MBbS\4\LDE9.YT:S/]XbcXfXSA:.AbXT6MO7PMb2g>GD@Ff\5W5eU<Y:Q#&E)#R,
/)#1#G8DHOLW\:I<=KJ2OgY7eVb#J_2O<g@7fLb)Z39KEGBeIgKD-6J3EA4ZgaI+
B.DcFN;c7,@+CDbaCFJ,aMW2IeU(JES9U;<+^g_H,IH-ZbI/c95,aLBAD8/dKKBf
IE[37UQ\^ZB-aKDaXWc3e7TE]/N&FO1aVPX:aI:g+c>AY=_\YN[]AR1#5FBcggRZ
PF.OA@(7#(6JEg1g03,Ng0382^2(#_K?W?AaX@:SHZ>?BE?dA5bDBN1,>S\f<CF5
_U,6M/_E>ZO[1/661<fV:8;06C\P<-(H3R@QPI^3bM9K69.4[SKa2XcGY^&MWa47
7F+O+Ka1fL3#NJS8NgLQWZLF#DB>b)EWH1A1LeZB\)Y:HNT;D2d<d&B:D&6EG+C#
US#,Y4LF=@ebIeY+AEde@6a6ZS2)W2d6b,S8M-W](OW=KVS5-fc2gF6Pb11P=aOe
NE\#Z[>Vb\2Z0F44DA;)S1)O=CbT3.faG)[=5Y.Pc:R?IBbMNJQaH/0E:AgYE]YP
^[W0aDKG2X5P&,Nc]A^S7a/LB1:.RMd/cH97_PecbBDc<OOFO]V-Lf+@CV-[K\I-
MaMb;#VM6;)-66I:GF)->W:(XdFb_O:e)7Z\eMFKT@5>WMb(PFXM]B#W>fF.1aa&
Z#bAU?Q1O@=AIOB].08L1G9<XeSe>O4g-LBL.8\dUZCXSFW,580+&^,\6EH89^f:
Ne/[6Z5KSHVOIE\9#&dEN5F]C<6dJP:b]R[[PIWa,CGa2GI9QL&LYK[DTBX7d6IZ
KPc?.FA4LWcE?+[K-&1K.O,YA\BAM#R^<4T6Y_1,B^QZ2CU58\H5c?(HP^MEGLRI
]+-D^4U^=O7H5K6X,O&,dDc8^Y=TRIPcC;><8#+LLfbL3Z-dd?8:dH\L7T]/,JHb
OTK45LTDg;.e,N(SL[WDDPEXEZ)fa6b.U(R2#LM@=PY.XfDB>XMg/14+\XK83c4N
H^9e1WD6dbMQU=8/LK6[9\BV+2+P(1^T:J7U7/G@d?;V=:gdT5833#Z?dR]g=/43
<D@24LB49J#_9dC\U_?.ERaPIEB;X:3+(b4O=2V3C7]3#ZX9OgcXF9(@S@WC@VNb
AM/0EA12TZO[aK5<?#AGd,XW+NF\<4OYT>4C5e:@F0FY&J]S^T5\<PA((V1OeSe^
13&;UMFRDH;HR@N(.H4+&W+\239)7fS_eHD,QXgU,3((EEdeCPL,#F<Ke;Hdd;P&
&:cB8IVM]?/&.@:/27)]6]59Zfdc66XXX]KV&X@_5.I7>0G3SNN.gEHAX7ag)g_-
TbWc,19?NR4)9U2g_GT33^28F<1(OEY>4WR&+6[.c5T83;=g5,0C&C[1)WISZ=#>
S5V)\a3f^6:T\7Ba@G,R2W/O(9;7GdBX98[=NUAI/@0AOda]R;DEeeT:@?Qf),(2
g@=>,_XZW@A95LDDgM>2\<UUR[.G0W#.O-Y9]ILW(Tc3)L?c,:US&ZU.M)T#6(fB
Yc(=2\b5ZA5.IH;-AcAW_AeH99g89R/DfCG\=_B8W[/5P[0.#<>W6<E2V.HU103H
T:_WBfVC3f<W6]UAEY8NXcX:=JP._/^/eUPG9<#Sa-M90cZgNWLY_]VDQCOUVb&[
6Ga1MA:1B9B0/Z&Q.O/K)R,QUE--X2?RI])T9:M,Vdg-H;F7Z6M=E_JPG:VCVgUf
&YZID+eNgI+SQ]/\e[;N=J2G79e;2M#2[TVUQWf\59LSOc>GRHSQA6SF:EK0NF&O
(I1dP]S@YJ^;O4HW[X<.fF2aH#/D^fC^L3\:M/F^6R5S#B?0BZcB,ZCM7RNc6_NC
eQM:g+^PUV(7.;FTN8M1KTSJ#^W(Aed8HgB47/+\Ka-dEgNI:/@)#OBZIe^Oa.^6
f@\7L7>KF^9BJMNAIgGAT_aSbR2@>]PJ<??1=@cd(EO+c^AFPa:4AQFb2e3^;^<R
6>-]@H-d@c]XOYIY84(=^RA\&:dPK=D3O:a_<]86+-#X++4N7_[f7MbD.12&9RW^
6C5N\3#(bU=.b1Zg18RRF(TCM6?;249DN]B,cEP]E/-#_LZBV+6&??IgDGSXL;gF
.O><RGB8Yb[?<1FO;&(<O)ML79(O>Je-ZPdF/fSBe/T]\Q_/>4b)b7(&dW)[XLJ+
D13M8Id(P@/LQ8NBN27EH^G]3U3@>C2QTZD[J4DDI>]>NXcIObWg^S?1(^QCGS6^
)7-(F6QGJ0BX98]DE>I^=)ME-XD&+Z/(g@BKMFO?ETP.D;^:\XJ2^^,Q-]\@OC8_
c8/a<SESO28aS?/XEO0f6I6A\G[YDJ/ZWXaH]a-GRT,H,.U2FK18IA>ZI@]+)TZ\
\67gL?Pg)<3Q=7]G;^5b?UcTg(K[\c9V.>E1B9SMAKK4\0I03bQ<H-H5c7):/62H
CCN5c/2ggbfEf@&4X=9MbbO[Y=#L,\X)ND4K:A(_KD^[^P2,IGWf@@Lc7C.C>HTG
]f6OI++\4O<@,2BTgS_<_c:_d&dJ1(3816.NAg#V]T4COReScGSGP9MGG/@JH[#[
&?M5CSK;RC&OE=bQY&@;Ce)1\4?5VXdOaX+[V9NU>EVEP9HCONEfZE/[^9EN6UC0
4aCLNRdWE(Y8/7^1_6IIQ[TQZWWZc(,UGTJd.?c07I:;C;.dD-gG^@gC(];&0:)T
ecYS;)L9.I\e[9<N>OAg5,F:Y>NEP^T2H2Se,ZG+K-//-0ab5gbOeQ[[bMTJH,PB
3gX;+>R_/A9:[S-@cIPEd6>Oa.UOXAUaJ84,:PaUG65<18AN819>0&4YBdR-[4<S
RWHZ>-1=(UgO+SX9G;Z?aC.[CA_:_XGHgFeZHHF54RRE#d3SIUL3b0:>ASW/OMd;
P@=BPX,LSL718<d,MdGKX_@?EP.8@d6F=WeQb(CaQ^FK9fK)U(NE&C][C^GefOH1
XF@[+@.4>0egd1DcF@1>VQ)^)7MPC7U2.fZ&X:W@UbA;]QEUK;SeF-2Ma-@gH4MH
FXfgc\]3)dCgV?L1559H@5E&I=_f6S98/3J=#fDeWd/7&fBTF^6(7@,JgD?O]8Mg
VM.6P>&;F+,cKN&27Zg+GH>;JVgSDLHT;^f1)G4SOMAQ>a[SV4aeBcAZ]7>LC]#L
ee]>2&8@gM\Yb@aC=1K4.D]/0&)\G/W4^QcT3)S]UHT4CIS5H_<ICM1A&UdgaX_O
^<X]R#)W^.:eMYg./DQ>[/-Y>E3T1J7C(EN]d1YX5K=-4U9V;T)@<;4C0N&9La__
6Y<TEVc?;[GFg=D(=W4?;d)@<5fO?+R?=94E_SH,9+cW4W)EXL]GP>>AFX=361B^
\J-C:&T>^V9bMDG/;;KSO0+;U#O#Q3<]@2-G6CG(B9)a]SS9G#J\91PXcQK5WP=R
>HMe\^W6PJTHW_,4,<DQE^6X_=28?Hb6MbZI^X:fB7K=F59HJW_[54T+7VUF3+9=
BYVGE?]QIB(Mb6VKF0fIMMFFA5=@.)3Tb/@U1T3=W9A1V>U2;V^M/5SgEO&L52d6
)4b<ET\8X2aS_L8#CLc<@A(SOMGU.4bL3:96de^f/)4Kc+MI6(d@H<X)HN1@a^UD
2.V),6YdAJW3Yce][(,_cPNYc9_5\M+<8Q#SgYV)2)5_eG_7,4f>CW:0[(K1+I<^
YYPf[Yb8/9cH)QAE#2(T2&4BKb3V8<(EETZaDYWAW138/KCG#UBQS/G5J;3K<(4[
5@=SC]1OGV&=X8S@U:<).Yfa3Kg\\P<6CB]#;d0]DGK5^\O#QGSG4=<Xea:e?]NW
O\3aIL#=7:(fF+,2^97B0,&@S2(\9M.]+,PGP>DO.QJ[4AJ>;3#BXcUXdPKgBJ1V
U\9M,?F9Wc@[R<.N(EO+JZcZGD+gXc]a^2X6H^LUVBS,D/XL[1:O#WbV<)=1Q=5]
QBbPJZGH\-A8F)[.IMK;,U(1ZH&&EHb^I_SdK>C\2AegOIRH+ZcE?<]\H[WgPK1.
If>,F#6SV]&g/+>dQbe6TFCa^[\2W.JQ<dO\dHHY;^EE+N5KWU]&WPF>Seg1M3V[
(-626,aP7F0aL-TS23(ATJ_Zc[XO21?K(2R>&#RJP>RZ(#0c.8,B5CWGYTHC3>#0
SQVge]K5VDAa,(D429@.SXYeD?B+OJ3fPP[6&XcKZ6)-_gb6US>/0(>/)\bOV^<]
SM):32\Ca=BVE?_XQIC6X4V6[-e3-7U@,+F>:WZaced/SdFD;/RR]U#L^=-]6DI@
bM(TJMB172#&9Y:2W(>=9><e5XSO<F<-8S[0Ed0I?/0RGN(YZNQaWcBa^=[]<1?:
;UU)[46E#K0NE?LD@)1+e<OKB3#E\#EGU016ZD\TcO.cdREJb>]FfFXNg6:aHT/J
HL&#X.^G;;GKZ2FPGg;b=:]\[0eA0AEFW21<45GT#A?4(TQOHES5--[,::=<#?,]
;_9MGERAdbY/A89H2d,#G8K5>?635+7=g>6ccU=F&=[81/H?:8X/5[IZL<3a\W2H
-8EaJ.)ZWa9=GD.c.S+T(GSAZf3JBQK8SHU/(1>Te/<S\,U;A\JTdQ:W/9@\ES]L
a^E#28GPCY<A-fgF2S,M?J=bL;R.96@JDK#R&PcEMWW0<I\Z0PQ07<fP8W8f)A/a
7cV><V?dZ8W@U.Z/PF#6YCdd#QcEO5QcPV0Ub2<-X-/^YAHE\VI@b>XXfECd\b+8
5O0WE:0OM>-QL8EeT?aJ=e6e]:GTW()<Z6@cZ(ZeI&IWB)U^a4.N>Q])NP+=cb^3
Y@^KYM[PR=56L2C,8V(0bG,I2WBY=#,Ygbd=2Na6L<ZI64F06KeP&WMI2T40Td4g
R/(,,82bdRO7VB;].03]+R0.Y66f-&6aZ7][\V-Y/VeP9..^2cDHeW1@_3(ZH]./
C,4L<bL/1af-(;X2@\K&.<.7aKSR(LX,/[?c[>(9/11@2_F8AK+#A->Ce3[(;-;W
d>WB@03V-H;@FM_7cU7^;?G(/Td6H5+HD:X#](.B)(>4HB6dKf?H?g.6f?NeeTU]
_W87#eCI_QF6D]1A-5f66eT1N5e?H+O^J9#J&[UL@6Y#C8G0=,^0e\+/@B-#4&.e
-LP^\UC9@:<3LXC#:TBR)U48IMIB8XO>T7Z_BA1BeC0R@98Z,M4[^EQ_#_5eb&9<
QQTGG_9P4JDZ=Ib0>+WXMfg9\ZK1H>F64<U[_(>(:Yg;0A:]F4-R9Q,I1^]&L<NN
GG15g9).ed?VeUX]6a^1\,^2\FI68]:.\))0]FZf@O@\DOB[\>X9^.VX#EZ@Qd1<
<&N<c;JT^WR.E>=+a]72GZ#\?:Z,05RK=eWGG6C6-X]b;b5AT58#MZ8;8c(5H:,H
RN2B0E(N#D\]eF+4b<\49D&A^/^CeI0P2dM6e-f9M,e[<BBQ1G_@2>f:,[JXAaCR
JD:S?U02g2e+W.I(bc?8\68fJ6EX[3Y+I9ZE,5F/0(^8[V\Vf8J&WJ0Y(OZE&_G[
8TY\=3Xg>>UI:&J)&CDg)1#&((bOY^Le/48I?7Y(^6ZJ\\\UgL_S-@,8PW^&LGa2
-ScWc4Leed8b-_EWSWO-9:OXdH>cU]^4,0M5#@e_:Y5gV?Y4ELIWKYZ]2Y@aH]#R
5TQ/BcUV>[;Q8WDVB[bEd(4RG:EcX^MSDf9R#H>QF01]bX22g)0Q-48_7:\)LTb+
81/f5TR9gU;641[9047SeJF7YTaQZE>@@Z8/<]0_])A)LD>O5,Cef&FA&072+.\C
MNU_g-,ROS&a6\V@.@H]82]EAZCYcFMb08DS_OB:)YN6U9<-e36HQ+>M-MZ1#80Z
&Q+8a97PfWC1AA)M;Z05@8#LJ16/,@E.Bg_6F_IPMA0ZGgcNbee_g&T6RR?b4@2?
HWGOLK2TIR(<05f,P6Z/:[4DJ37G&Ag>-I:Vd]Gd?_QVH&#U/g<cE9]X?NY&2Hb;
^ACR-@/=O02/#>Kg,>/.OgAe#F0Mb\SQ<Rf4IaWPEN\K?-XYELWB(e=O/_8OLMf_
d,\+_I+32<R6AST3/4C<f83YF?0b_Oga.[3O-<<]D:MgV+R<fS-\G((CD^?_(?U@
L[P0XVgVb4UYbc+34?KX7DMLN[/6cT=RK[&g.e?J)_JO3E@,Vge:1I7+1PQWTPLN
[M#GCF6E:NX(GPdFX(d^U9_bPdZ+]5.9dJ@Tfc/V]._M.#;LQ\9R[d?]MMgC?0g=
bUY5B+:_,^H3aF1eOIWb6cJg&:V>,5\EO<cGLDFOF.g0WbZ3JXD:WNMO^=E-]PF,
HdcP2ag\>(aDC9=:?SK..g&#X1LX>L>7YTS&CR2ZG1f:bOgf^F>GL5;&&C)-_IaU
aQ4)d:fA73K<e/@7LQYHe]Z7ZY3>A.IYA#bfBJ)U<1+d/QN-aJ[R2ZF^FFO,ZRT-
/F[I\b-5,-/XH_2I&5:g7^0^@^WLcc:TV=F]NW.ZF;c9TCKCMOKXIG+3-@\N[e[L
KUe7BWSXPS7O80GV32c-L=#Nb;VVR&cO\FfGV.S+0T>ZU/6_JLJEbX;LbS2U,^C(
O#eFL<T=R=Z33DV::PY^:<>8O-H7)S+2(B7,gU>\W5<>&T^E8fTU]QIZDQOFBU&M
/f:]:R9:Ka@6+CX]/EU\V)Y1TMZJG#)\E+G106XaV@GY]-XGJN4:1g-0M?4_fOMU
3WYfbR,BdJ_=3:5<<aGbK8]6S_UGKY(Y_(^+#>Rf;a3VdR)RK.U[C&Db#/f,4V>T
BQTgF7d(XGK-J)E,OQ4C9OPU<W;X.;<(E;/6OcRL:PV:QD2,UD<9^9^d0g+Cb,,-
+:I#geXYW^3T7P3N3e+gSE0P1Mf?6]UcX?[P>IBS\TafQ(CfdbS,V8+4N>LQ)3-/
0R(N54&(94g=T8Z++URRXC0DV>B3[=0TgK)JTQ;DH23Wgc]Q0gB4Fg,>G4[AcF3Q
,CVE_[<,O64DJ,a.50BEB]1Rg6N\98KVaUG]2GWHD/0V(Le]WMD4GF\]eFa_.78>
G4AVBgd^Deac&5\\#5L5)35(fbPeNMA4Cf5R:P_?8T[M@<-AT9._[&ELV.KbRe0]
(Pf/V^/bMCJbXHCQI0Kb@c03X[CPdRY@,f^gXMHLbf&9AD_0Y6[HG^g8dQ\KaaCE
@N8C7-1G1KEBV+^(I-NE,&IG:OH_ea.#dcB6SR.\[8&I2Cg,UBQeLa<JDI-D7WPW
&PQH-.:7#J?Z7-F1D)-Y5;W^]g<+]d@U3K>F&eaA\1S:gdHDeW):4#IDEfNPISf#
W1P+U^IVNGG_4-KD&8Zg0[/MAf&166bO8Q\/NZ3I>cF@(+e@C)g0cgW3IF3E-Q5b
497B#;2<c+PV#R?+L+#E2#V91N/X^)>a@#Ue5#M:e3?J=-YUfN,KH<[@\E<<L;LT
X2NB54H9H77aBJ\][,^MA8@da+MQ3bVI_LD;Le(E>X#Q/-P\Y1;0;ON)c>?[4&.>
g5>BL0E=R7QL4cOZT)c>99I_#S?TfP=1&_SeY^463-9?Rf5MLPc9fAD_:dCMLO)4
5PAU>DV=U_eBP#cLI:f3^0J-K0SRC[T3[c1C0X[ZOV0R6;Uae\0/M0T;(cTa+;ST
a(N:I;/=D_Y)7888)VA=.MH4@#b=83]6ag+,&[(F+:GG33;fW/J&cI2GT=b^L\:2
IYCF[&6,6&(WZ-eJ\XP,RU1cG<e,N;P=YWF1Tf8Pa8b=5UPTNF(#R#-Zf[d14Fb&
<DZFB6c?TK1Q7U/R]\.&.cB9BH<1)2\6B^]03GC6R&>#3+/XGPT0R.>fB/KZEL^b
3V49/LI7E2ST-A(-e+f9>9eSc6d^^,ARXGLX(WHY:64XQe__/=+\BCL)A4.E-VY#
LY1[4;=Nf=\_X^d1DXM>8M[g+X>Y@P_^[V:WUTgOb-eWUM,96,WH_\S&IN]Y^Tg,
4dVE8@SWA?>;=E)YI;@f[K)g^46ZA_e@NSH;f;P#9E3cHT/gg5MGf4BMJ\YJTZ=]
5T)LgeL3T88,f;e/M0AeFIIf+BGSXQBa1]&1@NJR=;f(W9_1?:&^ZI#;L(4MIb5S
+LUS,RHTbgC0<E:aQGD(GSGB2TQ1A>.5?BV85Q1>=]5.cSLcV.^dEEEKc5QZ.?^G
H]1M[8<9=XG]_BT.E)PE:ILRU8=3X&-.SR-1FKLWg=ad?gNbZ=-J4gc@[4,;BR\,
_T&WHE>d)6(1W@KeAXZN)]CFJ7DaM=\S?V,gDO>]JB@\TPZJ:Ne3(;5W(\CVTd1J
#/:,E9UY4^0VS)Lb7UEWCC@F+912&/IcTZ_?,7;?R\T;\1=B/Xe9eYO+HEVX=d+X
PfKceL^ZMdHO4.59bc^AT3<MdVI965M[XEVG1H&F8=7>>HIWX#BR0eReec&3DR:O
TM@+EYf<\:9bdM[XI22cA8:8(R)/@;?&Y)f/@LTLS1O3eJ:bFb1Je?#AVHdIc]Ud
MebF/YTL2E)TE3+12E,81;Mb8GO231b69.4V#73.AX,ZAee)e.Z?c681bM+eG]5T
bJ[<^&.e=/HHDUR\SCLI53HAe5T[R1MTN<,16F+I2aHfB@=\T:3eTR6bBM6C-O\3
^OZSZL+1+@JO_&(Y<ZQA@DUa=&VZVO9()RTd20B=\7Q8>S3<@ZGgU7_@Q8MbNYK,
7S:0a[2(g@e9dU)dRVPYT0Z/J7eR7>Vge71<bG\=_d:<&IBTg+>BA.(\[P/L^+1I
7dPfTBSUdKCfggeLKd;#E\C0f;HH+A-U21_Vf@;C##e>ZIgD;7;GG]9cL1&H,/^/
GH:?K-D44,7?M^G;ZPXLaAa)9D1O+E=Gc@S>WPY?CF;[RW8UgbEH3Y-@JD@T=CSP
)A50D8W6OPTMG1/):DQ<QYOVT9=[\<E7UY8)[ZG<#@b3NB81-6L=DSA1C][HB>dR
1H_?gf0.2b<+MIJ?_F:#cdE\5#\9UX[U9&\/0+K5>-3YX3/b26[NE9e[b62PPa0>
MI&-GV6eBdB(eU_I_<Acg]Q8TDU64BJa7?NT@90<[efP78HQ^;VF#UXN]ENg<S1:
Z#HDT9HfbSM+\dedeZ5Ufg[=@eN^LNgBBf-V>HB]-2N93J1<:0H&6TBAL\R[W+[S
W[K^-3)b-,AA84Y37X-\KY4CMV5D-Q+OZ6]R,e_5WXP[HYc)f7SEB>E92#K&K.>(
Q7P5:(G=2Q^BQ\4WM-.SJRL5#5&GW,4_eWH9>=\Qb[>D-02AH2--N0>J&GTEK2<,
:1K_e_eYK0eS3b.[N=N_1+W[H]PQN=IP&9:R2RF86IEe[9dd-KPKJc-SH:0W\VAI
7DGMS-;[ITEO9+I)#Pf>b]VgSCZDF;UTY1Ef]dA5()G]c@H)Y1/5O+/+T.4SP.E^
:,J>+dHPN)2Q)Y#C&;CY+XME<6g>LUW>64GOUY:P>I6E26O1d;TW6a;cSJc0//Q[
_5?Y9+9)eGQ,(@(UXQ\AUE5SU(7(DO_40LURU-<+g.8>KD0YfBda^7MZ9&T83Ce.
.K\C[V7>>:S:\_\X;Z,H;G;(Z3FKeB>E5+><Jb=e#B;4Hg_OQ2/W-0((PF#+CRQ8
;UP(ebP^&XB^[:&<6_PU&Y4[4\HD-YfHF]#M1_\S8>2HN&aC:RM,E.d?.I9(eD]:
@B:T;MaZQSDLCUgd:6D=AcCG,S1=aA<bSK>b]G8A&]4;8=\&5_>V[@K6(I4F3MTT
9=&gb)ZNS&_E6::c0G@KYHZ)[>+EEN7W32ZI5-Ma4GfFb4\4cJRYG\cTagWC_-K,
H-gI?E-RQSTABD(T.V?_cL:]FeeYbJ:PS<MESY<b_Z+#NOa]4(C8f7J+c,e_T-Q@
IKgEMM@[V3MFDgVdBO+/A[8QX:bJX&E6cYP#O&R_EU[;>CI1Y.L@cB3d6\[2@aA&
M^J/02+0AHg87[Y&W<0P;feT7W/?4[(gT2+XcdFK4ZLI;KXcR8V50MJ\<:(&?LeX
-E5KfU0J(6U0W=e/&A4\6:+W.()86/N6PVa5^c6M(I&IfRePe:FZe4AY99:N.M/=
c,I@Oda\Y);<9de]SZ;E;<4O6C&W_70TfXH+K7PY^OQG1H3;C>^eN58W3</R=7c/
;\CVR:>3X>=MRdP&>7<KfKZFZHMVB=?F/f)A/3:@G4LP:H6-SZ@I]+4c>g/6QN;,
.ZTPaSKZe1:0S(?g)O6)R[LUGSXdgH8C6d.P:EJfW&g:_9bZD[P66f3L:&E;R#50
XG(#KYSI&[<Y2E&+1e+OC8Q7T-eOJ><e;DU34&0)fg,>6@d[^19+8#a90W-=Hc(T
/;[LLVH6#5RMV<\BYL]BB8[WBFF@9O@</30C?aA9BP5K,.AO=0Zc6fa,#/fU5H,&
:R-LXb.^KOR23,F2&]Z>dbZ^#8+P(J+OB;^>D6@W?I-[VT_IM>N^4Wc;]?M=I+QY
F>F8)Qb@B(<.?W4IeAQT2NK89O=MXUF6c1NN1:SFQ-MTVXb3GX?4YTO:[>(<Te@f
^HP<e9\gC],O.=M^C7[78ZM^e&:U@g6Y,J-aQMXA[,[3<=7\ZKVcAe&D\FOUOgHM
-^:c+3TZV9=U))ZBF?VV]430S^/I6&S(G:FQI:USeE.WX:AADcKL=c\I^2bW(JgZ
d96/T-@=[cG>[V)LQWcd2JIT8&<6f<RW:_4;X?5eVY.O5&A?_\CZQ83,,Gd?,;PQ
<^/d^(.cV>a1@UNZ?T/2JXS6f[&2-Z)D&?F\A/&.:QT::F(\/E?Vb;BBCdLf5F(W
)S.):(3Q;3)1&ISSW0DJ-)ZA629GC.RE[>+c/<aPc&>T:XN;_W.W]8<-ZKTNFW>K
Y8\0\b2I1L<9A40dG7U6BY;.D<BM17/C4Q?f5U697McP[C8]/#>:2SQ@YW>JfYR@
<5Yfa@MJdbd[<edY;)QFg1\+bSZOXT#/<L+ReY0b7]KA0T8#Y2=R/#e3P6;b=(c;
fa7&T0R]e9^Oe_.@RGYDI,0HJCHf85<?<_>baP<EfO7P)-1K;0=F3W&:5ZB:\P3^
[0]PHFJ+E_I5+,MKBH/a)@8ATPM[I_QC5>8dFUCg^-^&-YR6@41R:FH7IN]Rea;P
?28UC&8@>fGFD(d2-)fMMD^?7^U-BHFW@Q2JLNN7G\8c\Kf(BD/@Ha?2O,E;HO>8
E,7]R9M2IL)FEEIKeNW:7/>HEEGXdR6ER+7EW5KN&C<H_/RH;K\9U.K9N<-85;3W
?;&APJ=UDTS(BWAY>5:Gd^>6(fB0O;#;/6e#JV/>&]BOgYR6U7b06M]JdfZQO4D[
WaPS0YP?^L;3YB7Z61M#PHA1a]@ITEb@\59+eJ9FNH1[?9)K(YWNe/e91//0bI3@
JCM68]H<9GM_]>2P0NX)abZP1)VH56&\-^>9?)EM<b30S=>UIKX>^7^a=JU:GSE\
-93?^^f[_]Z&:I@03&S<O21eQ@Q)YBR(ZSf88@aa0Ae=#d>OegE:2M@#W1V).7P9
SK/F+7SfZ/;Ae;IAP8-=Ef/9a&O)@5G44.5J9:V]1??7B@I#Y@9;68N<9BVF->dK
LRXLDK/?;8d;Df>DQ0\HB(P1BQdZZe)?^A7X-g_25CI+f_ZP8[;/UcA#6(?C\O1=
T2^8UaK<G#_PI+4PE?6=@O4\@KNJK5N<@LH,_T]/RRSBOED)S:Bg]?B^Qe,U#]=?
A2f2A/39,d(&:K/SadS^:->-226=D9F(7GbD8^STHYA)eWY43H;G[(@J>e-J3edg
#6E:H0<>(45V2f&M[UA7(XA?L)Oc&[8L@3f]=VcI]bDV.g=\@R^KaM3+\Of.+UG?
#0VHQ+\M73ME@1>.?e?HL49_:N.9A4a>R\58[<1I7#03F\)<DPY,RL6_.W<8+K<5
V_4e=0/<H45=GG>4g0KAG49_I4];Q1Ga@Z(9<L+8BV-b)&b_PRN_G1,.O&g26V0P
I_b7[#ZJX6OcdU]>012SWVQ4[dDF6B?.Q]73USZNa[Q-NAK6Kg+e0e+@9+,M=V]g
O3>UQIJZ_[X1bMYDd?:H+D46Xc@(1CeJXOeA1?/MDbc_aY7BZ)G^6@eK>+PLge4e
-\a_Y(JdgbN5XF(FcB63B:=P;fA&@SZ0.(T/E)3PcOEGCLY]IVcRRS;I(CC^NTGc
RXNAgW4KH?9/-Sf[IW(a/\0c:OBg1L\a@6;_9GR.YJ&#e;:3)2@1R#NM8K\HK0KL
X__cg;PK2CIScCG#Of:VgeR@<]HVQL,8;9VaAGIR=;L2,@cBN-0TFe+DVc.AJW)+
R9SO]4(_0(I@>W?;5@^H_C9^E8([0c1GG#UPcD)5^DJ[54.^eUUN52MZ)&YTTYIM
g,C0A4844YKHLEe8Pc8)\/7_A^-?dCf0GP^_TR6Qe<IC]efC#MN>(O^aE>Z0I(G=
?+[5H1dgC(=U/.LT+FIRTFc,]b4+=#b4[_<F49DeI5IHE-E&VL^@CH3;D?[@&>Y7
^X+24JMcAb_9bL;S:cL7-2ADQa@VXZF7W+5f1Z#SAV+5Q<)2PM8:>#TWA&\IOC3X
16EI_P.7cQF-3\1_(>V@)7R:2gI/\<4ICbO9+Og@3Z<.=K>>,W_[3;G-H[bA#2eK
+-f+[[SA/f=9<73QdO?3fTMNd/WG_:E8F#/CKJ);6S8M\S5RBeYPWaFf]RJA;Z#8
F@Z+Q:&,H;X@_-2/GH)]LgH>=c;+#U59AQ;@VI\N<J1@80dB2BI7Sg9faeI(e;Ta
7]/XbS,SS](D@CZ>^-H)&TfX-Zg7LV]9WFffU:IZg4I2^B&cGaGKW>/KY(^T._SK
R&[LEc8;N-/Q30GfLgQ7<>F:SR8,AaeD&1]IHf+(D/D4&K_K3J/f,BEQ[&WRQ[Y]
ebeV0K:dc?,)eS)#@;ILN5,SR=C49Y-(ZSYJdMV54-#g(]&=0dS[0@O;+1]Ib[Kb
MAP-D/1baV/XSM@\ESDQIYPH#cfgJ]CJA6]3J(AKT&OJEEY.^MCgM6eMCA7WJRb7
YIZ]BR8OVW&E76-8DVJ.HE,7\(1N1F;U7\W]Y5K)1Z/eTYWQR=fTLG)2)VZ:_&M6
UXZWLLQS]1+,AA0aWF>5&9(VYL(=.=_^H+E@6YM:0<)f<U#fW+]T+P/)QeZA=AB4
)HOg(F[&K>-67g[>KH(XYH1-0<=ObaSe<Q54ObJK/HOPF7LZf?Td^@RIW9ZV7)#7
Dc1V-;N=c\W=(8#2f@e9/.BMU@f:+?T8RKAfWZ)W08X9NCTD1PYC,:]cHU2G;(,>
?1C,XK3#8R7[4.(^+Q.eW.7,=YF@_N#=G.VH3/S:S-;2+9/V>H,UVcR?3LN.0d:0
625V8Q+S41BTUK<?(1]KR+UP^J76-^3E:+_L(9TN8P3;G,/1\^MP[BH:;W1.5FE2
WC(g?@e[2NO4cU4f2ag-_(X]N07I:#^fN8::gE3#S#6adQ<-/W&Ie6C<Me4AWOUZ
N<\T/0T0-+O\8QC2<OO828(&X]Qg5^EN6V\_1=Q=V(Cc]/IZQB,]\Q.@0WYAI^9:
>MLHK\U;8B_J_E^P^::)SVd@G;P/C^-Z=8?Nf7FL?IHZH[?QPYZO?,Rb?aBcA3U;
,be(E86Jg&ND8:#Lb0=5K[@<9PT]+a-5(L>UV&LM#&?F/;IYKY34,cR1f:EY<a#f
f:,<D=DSeT3F>9FT:EMGddQ[c3UJC3U92].I#/cfLO_YD^>3I=ZdeADb@)(2?NU>
QO_W#gAWb=T:>B#KZGE?DMa7=Z5eHScSS+c09bLM\F9L3_AICYa:J3MTLU^R]S<]
48DTa,U._Q3^Z@-Q4JP)E\UUM<?IC=FALISBSEAHNRIT,]@M)T<(1e1#:YGM]M\Q
&N(4-;&#b]PUJWNZ\M])[QVS,TXYRe+1TSM6Q:KZ=?CJ.Uf;S#2P63bGHBf2S3Fg
,)@EZ+.=F+F[I<RD0d&E-K/QM(PWP]^/fV?aGaFB[?dI-/>R5(H#Fa936A=DRV12
9/?+TA5?fPVH+__2#I5=+0EFA&K#7XKP8b5g0-J,+/=IQT9FcXWAZ>-RM94TY]<E
;L@IL:B)N]5Zc8Q;f>I(QDV+K@B9Qa6)#:dOKf=EI:]G)@4a5gS(-OV,&+W(b+SW
Y:LRLf[Q)?aTBAYC@^a4R30ORURQY\c@T.TP+Z0fG/^-6c(EJ4NFPe]g[?4e1)MD
3W:/25C5U9a\bV<GSY=P75]<Q&TG3=\;YJJB]b>^/UFV@?I6F(]/:@]9I(WBaERL
d<9]_JZcR+KWI;I-/XS^65ZcPC@;DW,0)&3+:O0W)M.dMYEI,cGN;?C<E+FWQg]#
S\5P8X9F\R@&(YLM(\RZ7AL1:1C@CJJ<:5L9R_(/P<G>1-,WTb1O1Nd?8]:TgIMM
a/XP;T#.Q6EZ?Y(F(V;dN+VPF4b@8NJ(feE-6fOD\eD:F]0\M^f0\@Bg8gH+IB]D
R2Ub5MT]X9ZDPUESELVC<;cgFS;RX<DAb/g>5LDHUG<HZcg]aM8M>_A6^46+AO^D
QKeH:b?2/1^N]a.6JfJ&YN0=1&(@C@TS8C)VSCC9I]W52@2C?IG9?+H:XM:gV,20
B]A-4[_H7D/[ZTKX,7_1JK0b^46:,4]HOY->EEK_:D=U8&]3>BcGRbf7(N3BSN+F
2Z[2/CC)T609H]4Hb6O#,P;a0,TMW@GGR-;R8;WG,RMTF=Z\R:C]/]d:<\c@Y#P4
5_OaAA),4=#T)8]SG:1a[,<g8K&JaW0#RE0WbHROfD6T7@a/@[2dWE,8CELdcMgG
ZMVbA+C2YAb\\ZC/8d=g#58>UbdNO^9((#4ZRbD2FVEA)+33g5#OMRXBbf&OA+4A
Y+NLDETSETHH]@(X1J?ga6S]@YSe0GA,)b_93](#4<b4K@UbMOVeINT\0<HDIWe(
CeED0A>Q1Z4Ff+30Og<+gK7=\Nb3.M/<Z>E-dUJ63E.R#9Tb@[#ZcKM<,<<F=1O6
DAHW:F1)5(WgZBE22&C5cA?<c/K]WURKG5H;:1fSJCc,HNd+Z08W<^/[;e]_e7/;
1<E6?6GBEaT0:@/OR8RW>_E8/;AR7QTAMf6XM&=4.Ea2(=T+0?X:M__Y-I,8)D=S
54;P]OU^ga.bZU,T31>^1)QTN7+bSUUI:VOF,]0U\?_T/EQe+2=daP5W<JA.JVf.
\@b\>-JRfNL<RW7ZR]-BKW()K^_Rc/BT]4DVVVMU0-cdT?.<b/N@N@_=G)(>TC;5
=Q7g54TbRDZ2/:;6C+O6d2c.)ID@CO1\GeH&Ja(3)X^eTaPT0:BQ98B._S_KK&^F
.S;Ab=-WK)H=[FI>a5HD_fD/NYVTU(c#c/]:6e5DaUUQZXEIVV4PXU#>_aYaR/WX
eM&TT<g2A<;F,Q:40I]3MADQV#]CKU^F=?&f@<,g2H?2ZW@B5,)FGJ:5gAMUJ9Rc
==DXUXWRE@3H/D8W7&E.+d+D__1TF,gaO5=U6b[4-32J4?Ee@:1TL3O>>WU+TWb+
@EaLUaN=_PKJS8&:NJO=@X@?>dSY_;2@^0IT@?F:/S:GSN9<fRIUG>7TV_IMX^&\
cb1A\@_<[9\\IM]\5@E82.dE0M,-[e9eT(D0_J3/#<V1D>/TgT/^XXKe5<Z,]>JB
X\7JOaf3]:2Ve_3FYY&C+cH)8EVRdbLFCZGCU^ff^O1\U>QgU8dZD1LS\;^,H@fE
M&3<g^f#G1WA&9E]fE\M&0V8aLf\DOdGDEAN;W;(LYGBgb2ELb=cVL+UV/3L[<X[
AI&5;17^PA&c+S1aI+-K#FA_GBXF@Z@/W^g]MR)SY;fc5be>F/W+NS<bN?/H3[&\
U8+M9-EMfBZB3A[WEgV14@@Q]@6fAbHdDXBce1UVSG5DY=.gMM5J4_JIAU64YV90
M_I3\CTH8#\1VXA.MEZ)Q.:W0@Oa?GGMe8[V;X>_BWQ_b:UE=A(JJ=6UZdSb2C+<
5)KFJ74EY8^+Z-4F[T@)K6_RF@I4B):_0G_8B8MQ4U0XLbZJBCG5#bJ),41[6._>
b+aG2Qe-GT\bDB[VN)G2S]PC/&)S)4XS#ARF-8]S0-d;#e=c9cL9dC1QHOe9C-IQ
NP29)2CSQfeM,Y]8gV_12SQQ6,@d1_b>9Y85IYE>\dC8<T>DZeVVP.ANQ(Bg/URA
Vd=+/&bT]2S#fgD9:e]K_Mc7>9g6L[^RPUQ,0HGIRWeIdH[IaEW,<W9Bc&0H:-OH
>(O;P</<.=T<(=D@&+6S0I0C8>EH23FC]g6O+F>)fI[QLd:g<^^+5M\FA#5gg3YH
]4/\),RI>_Md9W,e@6&X.ZRdf[_3E[XI#9,bd^A1Ye1JKTA))\fe[K3FFcE&2?1?
^;7;PP[PJ:WW^:;+X\Z=]JY.eQBSFaEMZQPB]e-X[5;T)6\)H0>]4P;&),6S928.
0G=]M9H11-M@(,Ff)9##6cd5-e7MHH.\ATZ)Deb4FWMWOMIP7cWGDZ4ZX[;N9UbY
+1C/5S^FaZ=S3I2.5F]AK14TV#e_T9+W_MJ_3E(UQ=4;<@>>(V,f89AG@],N7d(D
=cQ.1&P<@);3dP_74\eO+E3FXa/#[:FP,?@1&Ne/W?:&g/9IU\+OZ7[LV+gX9_(C
J@#TU#S[=K>3edOZFZWc,ECE\UM8?Y;9&37Z5<_P+<8.Og[g,T8&=]M2]8T194cE
JQYPS\1PFY4;VD^)aDWdXR@Eg=gf&.bBgFOg5CV<;B#MJ_>fH1B/JX3@bGT6N8;Q
;9\H([/QRO7OdI>=F4Q_@[ON(,8KP/15OXfN+CGHA?UL53CC7<4LITX?;TSF<9SK
1E_39>AIgCSeF#4BgCX^^G9c:(+CG@b3KQS=)<CS.R@?N+.5J6Y.Y8X_8M:>49C9
#cXJ-,_<YDWT<CVYD(=eGZDa<#K[;A7VLJYV]/J+L1bNd&B4CA9@KOF,DSW(<MPa
b7CDM)(\#VE7CJ_/L+=F8:6G/]\@FIFWGfbg-#?MdR#A>OJ8BNa_a5cY)JdIY?+:
8KFV-#:B9>eUJ;(:X#-/P&;#E)>[D-V7,>HbD8\P161<Y0>ZfNGC0bN,LV-ADT7Z
-,IRAQOH)dfLW1g&ZFd560M[WVH?XU,YUe<V4AN5T//=4(6-SP5?T9ST1RL:3+CX
69M3+8@A+Y.(S4QdU^?)=Id4A4EZWP89Q-U.@CcW2MD6TB];>=J]DgfQ;&B2.VBG
9?3Ka+CdH+6PYLAY^^gYB-6M#&D@PF6bVV>2WN^)<IgVAaK:](T@Jc/:0,EMFT9U
ROF>/DY@feSOZ,G0&UL+BVWZCG_1+H]LX3^C,1@3R[,7,5?57^O@FZL>;7XJ4>[_
-Y=P&J8TQ#MOCXcXg/3Z<aV[F<WUJ7]IB[USIYH0]K;9PO11DKFI]7BJG@WJ6a,N
\6X?>@ROSYHBa2XZ?<W;&0(NSK;QRT[RG5[GICDec@O]@LfN,/5bfRO#8@Y7DAg@
S5WLI#AK?Y@E_)YddC#c>#0M)A3aQ_?I&,YQFb9^U6-K)^Nc(V?FEO)MX>D[OR8:
_?Te&3LC?4bG2<OGCD71^=N6D88;K\FLe\CVde:6PJJX@7<Fcg]a-Bg6gJY79<D(
8a[)Mg8dd.+,fMR7^@^\#K4AdY5eT/FHJ9>M33.HG\:@__?GK[4P0g7,4X]#7BQT
#?DN6VSZa3Q_F/QE^0aaMRNA=@Q;71/UHQ#7=IHUa+<eTDX>F2PF>_L#&NC1KGJX
TC=PMgE:7IaX8^+9#,U7C@1J[3MTREE9?d;]b)gMJ]Z=QJ?WD\]2aVY1R\-#6AE7
R<e8Z)e_#;VNDO\cD9B;@8(G<dC02e5N\APHA1JDbTQW_,,DU2cY>4^ZfR>AQc/8
P;;/092Z3XD=_b>fgKK:XIY36SAT]L@X-Y@1?;0#Z7R3\YL:\8ae?;g\a_;@)#JE
.ME@9@A)Y66_<M@?.7^-g1M23KG@g9Db[4O8>9H<Cd.\C<Q[=^)_3Pe8:<AP=?7.
8Q7d#YQT]UC_dT0FN^N/HNLMgHIKaRL8-ER6Z7<\PM8L;W-G^eR(@gX:9_D9RC43
35b2GJe8O9X3ERBbE<5?KKJR+;(MU3/YP0^>LEJ//@U0[FSTKRI[Eec@-)BKcZDG
3<;9XA)>T,E\:ON,+S^cbS&G7#]ZZ9_\J_c=YX?g3T)E7>ad0ZEYf(FCa9\YG,2A
8XW(.SK,Y=+43FSJ4;U2&_^E#]Q,/-E(Ua27EDAB2[bD]N?dB\Z/.X=/3\&g&RC/
9US;<;-WU,1DJDK4[7G?8QVR9O+6W1I^2&>7A>^/eeGJ<]AB,\E3Zafb<@M-YO6c
4P[IcJKd:(_F)7,B:CV+JP,G<_TF>#SZO.^[d1)O7/Y<SFM;=L(THUdI,J9+HWBH
PH8A0SA+KJ+4,bRQ/V>b1E+A^Fa9RL7X7RcD\L.;@;I.9U.6CKNJCA=1WKJJE@1,
(_B1:EdSST9bDSJ\Y&HM7+HbOe3G^_(29gRW_:K_I03;L[-O2?+L0J,b2NYC@-8V
:J<_[(V4C=Yb&We/._W3-V)8]E8LGQ?#f]NXU@]>0dY(7?W10Ua.>\]W_RSUOGU7
-DaDR]2#)I<VZ>9F]K9[:7\V)6KT?H&XLd1,916.M>B?0GT:2\M7+fgA;^f&5I@R
_eBfNQgK;g@5geAI]dL7Y=A+Z3A#)^)D,<deSg_O<\=P;\MRH83LWfR<ZNY?01_a
7.#(KM1EaPVC#=[US.4OBJU<6:)dTe78(XQbYcJ1G72835[R3[#[HeESNCeH=8dZ
F>[d9aHW6+JJ[#MVN>T<DDD0gWDN0.PQ;2+HRQ2U4BJ@S+_^cKaRW+,EdT->f#RE
HbYVNYbD:M70T?F2NUYd]RDfR1_LG:0>@X\RJ>8WK48fB-GgMR=LB/GQ,)3G+[;@
ICTSZVI#PL/SZ@>#O5U9a&-2,8TfO.dK>/9Z[U-PXY_&9[SdIa]J#dQY1a73BV-E
NOR7_;G10<7W0;?/T>OK,#.7(IO<:DD)I.d5A>.?/=,49bA+#=Z<@R1c(X,R7-8[
deb,bD&FU:\),YK1BcV8&&XJD9-E2)9?M<W_Z5/\Y(b&-_dVQQaU0e2Dg75D6MHI
<_I6GbM]F_>+PSY)+gF6F[=H=(SGX.b6a<6-^cTCf,aTL/=US7cNDXYM/VVLTaJ,
PCSINF&\3E0[g+f51>Y_]6^^)6ZB/X_G3,,BA@(/GF/DJCU65&HXAR[@6U#<A@Gf
aIHZH8>gR@NK5a>9+I[#/da(,#4#?.7M]/ddY_;e69R[<7FFWBS-=Y5Nf(:L2HPB
.;DXH+68a4^6f?TM=#8,XR\/,aNP>JCf]g,f6b5PR&,aQJF-GcJR@J<UH<D(CN;g
802Y3AJg:=E9f4:]CO6-Z?#1F-9VDS&Z;_C/<@C14[H_(WX7LE[d<W,FVL_7P;S?
FJ<\Sbc4FY70?F0:\V&PefLa\K@-TN\&-CUf\9;VK3(9M29g&Q[Ifa6][D+VLf.^
gMS+=._:D:RZQ)#9/<1O9D7e==WO(1Jeg\.N0JL_N:X-)IN8P#aL[WO@>2b-+13P
E<0:4QU+.GSO7X?/V.Q<8Z;\XK-);+3-ES/#O(<.X<0?=+&7B@[2DTPe8.2S4YC\
Vf(bNV1\&Lc5WT5Y^PIC+TZ2c<@7(BE4cY-3R?]-L+g3WQ8E-.V9NM]Wg,RR+2??
QFQS:P^URZ/IbTN1#5>&La:Z:>PD3<c)?HXZ(bJ;#6fXE=bZWbY9;1W?dd.I)^S-
Cf1VCgSRGK,?=\Y1[\6J/\#?;S.V?Z94+;YYLW;<R,.L1I3T&U3CVBRH/G6[V)ZL
8RS+?3)bB(9=P0[WK9S#c+QR@-)bJ537IV3B]4/07BfaFa\_@RCHgR0^_4@eMR4V
&>cBJU>+L[_PO=FaEgb\S1K[8,g)[]\85E_X[ZP31gY[LO-61B_V5GN-d78F<\bQ
fAYdT33DBL0P?J_8UfE3U+V@;8IR)LYZ+N/\S;)gI,bPX=LS]:AF33)(+N\cX07C
+UfABN#/FLA)g+I2JZ=5J]TBe>PB34&>OLfGG<F>ES1DS_CCV0+K_18gF/0.dXEF
e-X(+3N+Ue@P+Zg)3g#FXa-_OOGcB&5a=0_=?g>H3Zf,C@?2XXc)a,IWK^.)J+:9
DQ2);@L#,7JX#KZL4<HBS<GGU==GZ7U?b3C.bE)/AY7HD#N,[cBFM9CLV)V#b58+
N.[BGa\3C,APP-=)UWX(8)NMPc=R5,J\2(#^<YcW7B_6GZW</.41R@_JW;C&)(M=
5>A?0Q.g+S=1ISNKBXY;A[>B>[cJ+d3+1JOW[^U>#?7]PUK)E@\I851X4,V;(&W<
.McA&>6I,K&U;KdF(I^;3#HH/3BA-,<M6MF-\AY:IUQ&XOcD^=^22N)Xd\]c55^.
-O#U)\M;(8M=IR0M]1NA[[;G.X0X)E.A^22X]R:P8WLa#90.HVE2Y0:8WZ1]#6G]
08L4)HPWCb149J(.H&V:f[)D>=dCe?7d>HN.PUX/4g<SCDefJ@MGO4XCQbc0AW(.
,WHOVG19#c7RNUX5JdUET1NJ6>8DZ_e8XO#OfV_fFQPa=NF5bI>KOV]54.1BI6#g
G9@cb6g[a\AcIb0g9169XDVcXH<bNSZVSc3^@[S#ZZ_RANC+B^US;MUJ\DZD>#dL
Q>[/KUP;9a[A6WX[Y):d,T901&d>H\W,GaRHEe39EgO;,76&M)T@AO:)71-S[E.-
Na@+CD0U.=:VERWN9XcBgb+1+cL>9WK>Xg>E197fCUX)?)=IDS9#^BQJOVZM3<OZ
aZ(#+ARZCP9Ie6:?PH+>XGOG9/C4,TYQ#@3YNM(.R;]V\e&M6cB3..=C0M(\Sg2X
N&\F=26Vg.]XKF.Z4Ofg2^]Za:JW\Z>bM2BTKZ^A>O-4H\fb4d-M[^E/Y?R,g7<N
2\24cKIZY77V^8La39<8O<XO/ReSX7LSMO&@D-ADa/9=RV,-F/bcAH&>4JU_M6ZM
-Fa_e36YG<T?P,N5J.3S9b>V@KT#W[9&K7FGRVGRQ2EU@?(XJ6A7Pa#ZeG,f58HQ
:N]4?YSQ,@6I8@FS6G>HU-a[ND,6(\MLSa4[\UO7GIS_R[SLVg:#-<30(:.ZVBb3
H;U8<E<bRg[c\5-MR4_6F)BPf;4Y]>)NMca^R3?-)b+#^cA+b3MXX&7[B:KW[E:L
P[HX+5XC\WS>([3]gY?^;;5e9>TbSQ&>Hg0[+PT^1FS=FHYBU\P02b[_a77aEV,J
69JO3XK6?3?@?#.b//[4#]5150_MWI7=)b3I(36.:9HN\eYF(,:_011IM^VPL5XU
+.@L#a.#W)b0YCbJPYWOeFL]6e)RPf>_<[9R[dJ<9-RfYR+#ef<N4U_.6H=9Vf3a
V;JWPR=4U?FX4OUO;0-7WVU3HYL.O6K&.5A](f4V.d^W[e6=J\6-XVQZ(D,3YNZR
a+.GRI1HGZ0dVP@^dB:NTQ;;eI.QH0bB1NT:W7c(e3\)&>@<H>H3R?8;VJKSY5U>
_F8&=0G7II^MK/#+I<\fAWTJIb8CaZ[@TA=SF?I)L3T2)+=GcL-eNN>4d5M317S5
/T819_L9AB&TE/\=\ECE>,NQc-dGL1<:R4aP1S4IQ^MJTU6+985KZQOJY,S@FGRK
<LM80S-+)>LA:M:RI?bRQT,/XQ9E=aWFb;8g2WN@;RZ_437W(@3=1Ub)FW96GDEg
Ne7\BL#4cMMTM2g;0Q?0A1gb+a)<NPT\9,_7U2>S9MdIN/3;DM;bHg=F)L,VQ6@&
77e><W(3^?5eCQ\IIYMEd0ZS:<R3<53RY-MK<XbRA1e9MGT(JH(C_;<^C+:D&1&8
E-JV8I?Q5dX3#<P?I#\_@DDgI1T6cYPOWGb;O(.&5dODW<;S@9g7JTRT]2V3QK_T
T6g9GBCgZ(-.LUKJ[CR:YWOO(;[#=Kga(V,@IdE<(7.DeA#(,HX4>J#\W]#SLG.L
Z#Qd,[.^&@UGTe&I(60I:=M_O</CXY0dRTG&g;(TU;a^0RI=dfIQEeT[6SW7^\Ca
EW@I6e?MZBJE0>L.JAf)#X2#\5P_,SKeD6Fc[;GV\-=ZKI5]L__&LCAAVNf2U)\E
>H[FW:BfUL+.WDgeV^L;KI:RCb1=7FUR-\5[)&&0f<V)5#dLDARgCZ=GWcf\8?-@
QMa4FL#?<Y>8gV+..YEB+YC/bDQZS_eO76c:0]JgUN1:gRW@;B6dVKECQ43+IU-f
\Og^d,P<@f#FE[?K=fOXE<PR^CD.]AYd1AX+N,F:RF-A+^EXA>EH>-72A]b4>>V=
eEc;CC0W34M7OO]4/=1-Y;J.N+_C85V_Y@e,@7U<.=Se+]Y&fW1UbANXf15)=<^B
(3:))M-YXSBY9B;1>^-e5E.F;[)8-L2>(8^\>#cQA0KFP2HaT@aEVQWRNF#1HZ<@
=BdK7:^#e(>J:K<>P(Z?&FFNdVD3SNXRCZWc8\5g4gX3TFQIRKd.D/(MQ#g-OA-5
MZ(TSd-BT<CgUJ^QCVdS-#S]O)_;8\IMEQ8Q8a4)fd:7:M9B(4LF@@f(W.f-9H-I
+B7)2V6M1RLf)37B#+TPd(-WaZW1RTL5U;FU.&Z@VR=O[V)]bJY=]I6.F0@[+\1D
._6D\\?TLSc7Y:U;]>BJ-QX6/Y0AcCKP-;M:/&Z0g\&>&9H-\SJOK]c@:Cc\P08A
TK4=_GGIAR9IA8B]=6&:U]S/Q&Q,Y.:B:ZSOHLZ>:EPC(AYgT9ZcD@#?I2gH2P1M
MfXAMg6Te38F(gHX;C<C#^\IY5)6^2Jc&79cXX7fbBZB4[2</eKS).R-Z^IJ+CQ0
&HS-@9-JB<KB=cDRGI/-RU9VbE27&I.R?Og7d\XJ^J-T;0GFeZV\EYQ9:;K5e^\^
7-\(M-J8g;dYK(#L,=d,MA8^b3I)]6BH#ZBb+^g1:I,VA)SN)QY2)Gdc^VF+U;]\
acOQ09dAF54?NSfL?1^-@PWC.\J:HZ(dC+6NbAX6J.Z_1Y1gS9<JcGDXWS?GW^=c
/3,U_@H5]Y0K6TYJT)+,534=4e;1MN,6+dI>2H<7<>:VAYd>U8:1CNWS^TF49&g.
49<,+.Z/BBT>BWKcB6/,)Oacg,A<T?MN;&F,AS1DTN(2F)0Q@cf_BMZeR<B,&[L[
KG_g\RbgEK7DWDII[M6IL57=W_KME8OQ@4,c5gI8X+a71#EE1;d+[N.8Oa-X\U]D
&4X+G<8HXBEWG6?JPKGeVOe>AD<[^[.>CJ827Db,AR_DGJ5LB@c3.5KS1(_Ef7^Z
+VfOTYD5)6,bN?OSVLKXY_;E]=0A9c>^3A]1fG(F8&e,^Z_I@HbT?_e,3(V->b9^
6ZNVW&XbPM8Y\,.]=@d0>4FXV-/(1#/?Q;G5fTQR(JFR6KLcT(dZ7caHIUEd;W@)
[/;<9^\6R26W5^W@S,QD.Z<1E_cQe?G@A,FZe.2IYcO51G>ZG_NB@daXW1\ZM6PQ
^F5d2^bM/=SV@gKT;UQ=OEN_EG2.USfH[QH8<-0:S)eZL;)NIb4EWD;C<Qa0@0GX
LOFU3L0E:#AQDcT:-)HVQ^fHWK,=0=.C64NTW3_6FNAGg;6H]3c,^.G/Z9P1feE?
8D,21U7CDHO[D1c;&K.]_2OJSA(O]S&U8VLU)B>Q4-T-+[fIU1-<dIRA2V],Qed^
HK]#d&AXJIIC?d;gRU[U5A<#M7CL<YS.ES,X(4RJA=LaIQ1?#>a:E-\:G893-Ga7
)HdMU@DIP3OH4WfdadNWCL)4JJDUBWA23OLRY=GGWY^/;4gf;WP4+L9S:=-TB.I.
7KZZD[@>(T.V&2(JCSCFI+dadB38c5.N^]LU.g(PXQJ]\U5;F+\6OZY(Z0FCH^/O
_ABWP42]X(OA]Q?@IKO[Wf^XWc2S^;9,5<d6)ZG3KTf9/)P0E^>Q8DA4+8R(YR]U
.JPQ]+f(4:a]<MQKQ@,,3;cTHYT7]QRS@A(5f]1=Yg(]^0LP@X?L#Lb;DKaGWWZ\
)RP8F3a,Of,[RQT-eVK?:S&RgL4X@R9;C&N6f]S1Y?E@df::/\BT</JHF)+7K2L/
#2=QWBL8;@1JO9HP/W\G6F18HKF;.5NIV<>^=SQ(>-Vea2N&UcNF@/J.0>S<B3/L
.>(YUc.F\HQ^D))D,:SC,/XYH9.c/Qe9^@N#NE>8b.\T-+M[,GY=c2,BR@:AC;O7
GP5]@_]E;>gJV1JMM]@E.d,;FYNJBJJ^E:RE[\gPSgX+AOHT,9K^CQ-AI,[I(f:_
?-D>@6S:@#:=L6UJ@b?aAgG4f&P^SG[Q:IZO2,#RS[C-.ZI1SI/MY35Nd1JL/B5D
#\\VK\QB5A>8/eB86&-[W>4GOeLH)#Le?/6QTeD/^0Reg3GUVLD/IAB=#dM^RG\&
bKGXT[;^ee2EfHK7^2@b:+gEQ#ZGA.PV3Q]1;f0MeJ<FUGVfEJE;]E):_RSIQUR[
73DTHb@d7K0=V?+Na)cg+]HLH@=X37Zgg:]^L/U]c42BE#]Ka8.da<eW-BXB(,70
1KO/RAH<8f=?.;F&2;\b#I63EF6FacUEdfC4R0QO5[I1H9e8caP8e9/2>d@H.9eN
UA();+73QQ,8271711I.+bUeW&ad+8Z19)9OFJ52_AEgTeNUEH]M4^(aMP8a0@4f
I<-L0@P\^cD,KZ>]>W+H\&]Eb6>Q=YA&1_U2FD3/@8.Y0NZI,&Q^-5E=<dKU-d5_
/eWCY(.Dc@g1eCdSPd-#f7X_@BcK74;Q7-X[RgN^<_:0C8_LM0<X4/:G1>;OA[:<
IU\X?>e=ed@JfI&EDM4If1?IW2STF;b.,P&1\]R?aCfX>+P:ee4:S#WYUE()G=+O
>-80PFFOTKgQSfc:2-?&<4dK:9<ce9Ha2T>MBeF#)K&dN&e5_Z;X-g1FEU3DBZ9Y
>O<YK[[>X8#\KA,E5H0ZSbLf\2S&QQR.QZ@M#]\KR&4WFE#R08N>SV:@G\UQ3L)D
JE?ZaE<LYHDV+OABeTWQ/VDU39AS^g)/U^>8HC0&FJa<41<M82X(?WJ6J#&KR>Fa
DD4MM.BN?<Q5JF])_TgY.=LV(JdD4M-Sab^,TbY>@_B,aTDR1G^BR,CEdN)2N\Rd
WU+(_<MG84Zg380Ya;G3@Va<>7R,dLR+LTQW,:_/(9)2(fATHOQM_.K\J(a)(Dg\
Z.=f+RA9XfN7:^K/)F2UZ=.U6]d)Df^=V5)B8,^V3Y+A39d07EQ7OZCgEI79UF(V
Z#UT#KX)YJae78f8O@.X_<&<,GFR:;A#X]<,O._a-H5+gdd&Wc7E._)]66;fA(Xc
f76=J5[6ecWWX^(UecZdME#7^GVR)6AKR1B4L+=T<O8O_g_7&M<I_&4WE]8UK;;c
)#.b-^O/^?C\Z>47/e969+@D&95\&_&XI(H?J0AF9E)/g7ge3c)(QJK@O5N@XH8a
=fY>VN-[9^V+O)CYa^W[[e?G3GQMG2/:C/<HYPML;@[=\I#S)G::IY0S?9I8c6Z;
[=F6D,53?NAVcA.b<e9H&ZOJ:>_CZ).bM9YN;][M_03+2Z_DRVP<P(#<9LA&NV??
4b<@9)>)D)M#+6_,+(G&6.EIAE>>71O_;/XV=@c>G_c]dG5&LFWJW@#-YJdAbJ\D
N,Gbd0^<69WC0_I)T)(R1LUTLJ;PLfPcaLd_^DE?:2cND<4>L_O1E:[24T0SO_J2
O#@UB]TX2[3#&91-ARa&YILeBC)>2R<#Kf83K\7S?U1[7g[b4]V^V4#9XaI#bHSQ
=0BX)X<P3DO38A]BEJ6(/_Q-[Ec.adE-8H8O6R=5P8=Hc3(&6VXa)XQ3YREBTUHZ
AbgQO@Q,4]g]N-/\S6,M[8WaM:8O7+OC^8K)2cG3?:4N.b_F0W^#>TgcW-1;T842
B(d6,@eR0gFB6=.0YUSA[JX[@@+/E_7.eJN0b(W4XZ:+#Y=ON^.H,eO[0W9.;O-N
=IKH82c9J3,PDWUH>>X(#E^4)H2K?8^>.X5:J=F5(U0SXZ-0]U1V[J->TgMgdg?I
_<H4&AVd2d,TNOH&c;AbNQeb-4D]f8MHa@+FI/Fd.bZI5adNbg5d9:F_3WfN=HGI
a0+-QT+5[F?5cgE_[M8QY^,?_>1]53XYMI^D:5<eBO[NO.c5<H/)(gLV<Z0=gZ#]
Td#\H\?c8<8L[b:@L];;]67Q?]>TOQZT)\1R#0LgCP:>C;14?<-X?1;K(b+c)dUC
D>ZZG_YVAaWWC)P\gU)#LNNT7,;HMPQV?Hc,d7Y.49)YC=)1)B^AP\UD(@?0I&;3
MWb\\K^>B/d;=AXB-UZf=FZ)@[<29IIf;=8SF7Q9QcfED=Gc3Q9,QP#);1=eF@4a
7bS3^V\L0bf(R)VNDK8IZ(#a)6R((6SV.7<O,PW=C0<LXBfURN@>7UX)@eEEBBg(
7_W@MPJC:-F31S,:AM>1J)&.Ee?P-O;QLZ#F((+^08+WVG5Z,d]#&e1;MMO/]G08
QH-UP95U<-8IL\4U\SFD1L1R:e&FI>W:XE6VSYW1G8QG6G,H22)5Db[Z-J\f#_Db
.B2PP2-c.LDcY)eN\8WNg14VKRNc=:>E7M)=+EL-/6;HD9AY>+@+Q@LW[0J1[@E5
:Za23A@ff4H+UCMJ=2C@R@81P56aGXI.Q/I5gS?KA]P^T#_>(C[a/S;0]0:2;N=)
/<]M+\_c6D5JL-SE??\[P]X_OH^Y#P&V>TG44?1\VI7IZ@dg9@@8>Ie6]aAXH+B+
TCW_:d=D2)M&;ZXI28_4RVdL4F_9U4R_ecOLK&,HN_J62AY4VDEcR^3dWQ,U,QdP
8;/aJ_4OfK-.J15L/XGB>Qe<A?<PY]4P[4YX-#LZH<e>_E-ACR]Y//S]LG9HCc7Q
W&;UVdJ_Q_5^KeUa;=GbG5b).2R7>b8dT#(.DOdgT1U35H229g6b+EP4VN\(;6.c
:DbJ9=\_D>><\1ZIK.38f-\cQ04PWR:fJ/3MKUT-A,^SI3QdF&-1J>Q)eTS<85f2
U#=]2/L-<,]]?V2/XH1R#JUd/JgVWIb<:/a0,U@^OCKVL5Sa[d6_.-g@GEY<?)]8
_];I[)A]NJ?/\64OS&1J<XQ<:=M0bPaRGT&[\?d8G1bRK2TdAS9J1HC#QR@\J@V5
^/J4(LJ;3?GOeWUX-K5O/1+U0<1cQMPLI;_VJgQ)D+=:(N&O]=A^H.@Z\)442VM=
+D?Lb2a(M06J]WD(B98&:B8Tg>X#=YSLW6EEP80(TQ>M3ABN?029EUQ#AeAKF)Bd
FA/BZJ;MHDD^fD6,/fS/<@IUV]6T=WabSe7U_-M:9/?JUOJH-eaNGLVQ2KP5b2<L
01?M#N?aS/g)U;V;<GY)?-_W]>.DS+SV=/K=e,9RQ<UP]X-M+bVfeKS@-UNWXf8=
gH,XKGBHd36D+Te-=O)[QJ2\UD4]GR_S@>.7cOE7fXcDO?9&C1S@Y#.fN;EA<Z](
W[D>[=3_0XXL?3aIN8[bf0X_Hg6,LOC&2A[J0@eRM=L>bY>MUSKbWF_(LL5dN0>D
Y=AT9dGT(GeL->f_5,5GISM/3UR8BO9dL+M4?HWQRR&G]0GRfHe@X<K&(UZ.=0:J
RF(4I3d_f68-@XF=A5WE;Y>:.:@ETeNX>\2d?OeZF^T7D6UEA5_\7K@H8.d\b>9B
))2J2&S>)A>(TMg=_)XSG5L+#N(ZdZaUKV8<-[CS9XG8eY5Nc/MabF0_XAH34UOO
cZ:5#cg=N(>PL;O&]/N:EbQ82O^9535EJaMX5^^DK?UI#.IZBUF6/99GP78eHN2J
aeU,JZRS]U=+]Cb.__59?WMN#/SME)fccPU?M6-2:aXRG[G(dTfYNGYQX<=(HJPd
WR9AH;+2@1#bDP7J8AfE5(e:)M0W^b;a<-OQTcDaV:g.F(:NeeZDKNHd[f.TABd4
d8:).c2&-6gX@YVTI9U/7_CTLOHF>Ja^MEZXLOU<<O8TA<-SYJF/JO+)=D@D7eGX
V<V3US)NE^(gML)R,9\aX>,;PO9+EW]ca5^NV?eO@6RIL2]02DL;:WN0(ZL/JS(a
,.2]IZ8=,\eK_7[M0Y=-c]dQ-.30^2Z]_MTJ]78)Re8VAMf9\V^6=/>;B8Y[Q@)K
8T]WTUEV[GXSQFNeGL8D=>[Zb^OX&(D.CeCPfFS]:(gN/G777^S,QHD0.Bf1GC^M
V-cL5#+/HaCc1\EPfe@[WY/e>(LXIdA=_\TE9YC/1TZK\/;U]OBf8RI4#^Ne1;LA
.+HFFZ@daK73YCU,d4;e0b7O08/6fHD3/]+:a&6H?T5-8/bG,)AIDB9,9[^bg0dg
,XW\fW,.8\C+MF,/3<\]LQ;+_\TD510CbO&]MYFXGC@a&(B:Qf:\I.&];dWdF):b
;2aNdBT[Yg)<A92(IYVOY[W))D@6F5FIQF.9;9^_=N/RB#dP-AJS:H5:<2P[N)M0
-aME0a4]:V(A-We8b+e0^)YV.gf&0,CWeU9X]fG?a>5SY>fYW&X-Z>J.1b#X9d4&
Q_aH@.NJ=98fgcc./Z.a><V&KQK+;)<D7&9==[ZPcM<a;DS+24M/g[SH;.>RNM+5
?T1/(C_FaaFI6LI0BbfP+eTWbg-eN]/?@9-.\;[\d@#D)RJ9O<+J<,>VY><.H;5Y
U[P8[TXEF3H?_>[OI,^7>MAAYabJA9[[GMeMV3;P#\C,,7&;RQ[?@1>:&[Fg),;;
Na^g.R]Z0>>WKLV63HPCBa):2K\)+[I-e:1]?6X31(MOgd)a8D4_WB1QW+#IaZ@9
,2MOeEV@7b1-c(^)JY6A?ab:^TZaPMA2Ce:)).F6Tc,3KPW8<B@9d_T.[\A#:0XK
d>f5A0&+3>LBS/CbFW^?We[&9-MO&A78KN7<ONQTA&;AI25V@d=_)YJ9N@6(Z65R
P)6]aKSdWa]bg0Sa<W;aWAR[<>b:39=6dM^_&&3QaW[WD\R&#G#dZ6X2g>@Y@G>f
^Hb531ADgZb4D,b@6DR^+O3-^XF:T]HVeUb7_QJ(:<RfW;(S=gDKb.9deWT,4+R,
V4-?gcK[NFY=FCe7F-T&&@1/<Ia@)5@&7ZO3YYYS:JOJH9ba+)?JcMN)/Id&=K=:
O96//Fa]ega<a,1NA46d@M:bS,:YO.W0JM^VDBgP]);GGe9-[#2?,07-c3dBE2Db
,/AR#TGLc+]L7)];c7N7WXC:fZ.)Xe-?PXT7G<B>K_ULCe__]Y=\1N:,d?AWAR-+
W;>PRX&XdZ<KU;T]cJG6QTcV3L0I80+/D5a+\N&<;^&bf;g:>;PZ41/S1/e99f#f
AYP#g^W6fNFV\/Lb[.-B_Q3BD2Z1FOD^c5;1VO^M]9I?N>Na/\269LNN^2Gg>?T2
J0MX7(TZ]-(Ce48eS:daV2d2M0)094=Ug@G.b93cNF+a>/L2+DU?V_b<d8QVXKR:
X/NXBI@HNf/&Z#@)(A4FY>X9ReD2<1NM)JIZGP)O)AI7Zc_6V88Z;=^XJDYbP6J4
)3=/58f7WBf;7TBaTC10\IF]COc?15#BLT0G@a7PJdMg/4.5HbQF2&8-4OQ;R=(M
+)PP)/XA@a6)++Q?\S?g3PF:cIKO>WG?A0JNEbYX,7/<N9TOM.J7a-M(Ua(@6VEI
XO-8\]a\<bO)#+&8\[Ec>0O:R_4]G)IFW0K]D@B#+I>F\,Rf#:3b9M6gACB[9Ac_
c]06^S:P@g,+D]Xg-eDWL0:F3=(]Aa)8/HYV1=ETY8g@GeF>6FaMCDXC?Ja97ZH]
BMJ>fZPY4V7^Y\WKUUf\7Zb@WY-D^)\G_5L.b::M8/N<f=LgT\1+@V1eFWCQA(H\
^7+V;4PH[6EaSUBDLE[Re+&XTX9[7=I8LEcKH\Re])6@,PLAWXgg^]RT6Ia9?C2U
g(1QWRNbP[M5LOACK9@bfG\01>.F_1f.8BK)9PF,5EEYg>G=Ye(W6ULUK\;b.>\X
Y_\VcPSOFT_P6P.4SPMCd]F:SJ^X/&2:@QMcY19.LZUJFO707C&K8(91>,PNHZO\
BJZVb\G&>eRcM#N_S:<fE2,\FPO=HA&:CV&BO1<3JSeO-::59>U[;V3=G_QS8K2,
=f2__KUFU6BN_UMUB_,&L:/fVHf]F-[(7UZW@&?2,/O;FT,X3:eZd)5H^9TDJ43^
:J)W.0BF)BDZ9c5AY1IKL;HR8V6]H>EU//a(Cd5Y;F_T>?_[g^)8CT[=G)4UeMOG
?TD]Eg;_\fJ9M&-)HJ]@10@Z<^?Z8;D?)U+67_QF0P\)8[2Wg(f_6,OYIb?\.(KS
Tc:]D(:_(,6f^ICNC,_CY9/b<a@32RXBRd>OK05RULN0O7Ie52cK-<_PJSHS;X<3
QM>fZ>/c5^f=]A]ZWAQ]SKO<1U/?G/5+b?LT<;gLAdMU+//F&64A54eGG3(<.GG7
LeX=0Ib.=M<A/AB3YW;Nd82K=J06XJA5UOIbB[R<FDgRT88P()-2Nd]@#7,@fMZI
HZg.O@6^QI]6I1(/T3?CH^(G+XO/S+.^.(6(0RT(.)ffMEaC<d,/T:]GR\Xc/#[_
73?_P-R9B=GgU=MKPfJd7QJ0dYKW99J>AF@L>QX?7CW]OdE_ZN<W</25aA0bAKT<
1[b/IPFOZA;1D_F><6_d]<D7KDGe<W2P^?1IVRg;7ccSe[>bY3OII;>_O]a(;UNf
)d,_?c69/)_OefSc/U?&A3=a^6R=U#-b#0&GH(##^//<_D@;GS?55RTKIeUd,c3b
AdXY62dT+@Kf9N^G,(4:9IURS]=+>S=3e,E:9R3[;H(>Y4-B#&;A1?eUWMVE:V?N
1\X/N2@PYG.BcT=8SQAA&JZ/&#^Ke+VU039\U/GI-4K+0V8=?@VX(b=50UNBUXIg
I/,ZU,Y=C?/2WZ7<QP(EQUd6Rd.8S:dNEO3?]PQB)6]V]MT1_:R;D\a@^DcW6[/5
CQ-e:ZgTLZE^./5Ccb3;V@L_6&RWR=C^KP>A88?G_/SG:<\T88(@1g3G;J[LOed@
]6W^>ZCGVf0/Kf7K]#K/=&/b.WZc;2Yf-EBJHJ[I.V>WFKLEJN;<>a+[@;VW\IXP
e^48/d-B=:-)F/6=BeF;HIQ+-F]\]GT[(Q9(60BK)_9dTgdZBMA,@(:QK>19&UC=
R>Ob@<O9]A&Z4L8CTd=&0N6,CH;a08W<gCT&5.G2G&P^)3@<Xa6_gC4R05^T5V-U
=R<BI(WF@c4-0KfX/,b_<J10b.1HScd,U88R5A#g\EN[:_^@?cTc<Y=A).&9C(16
H#7PXPZOCXB5dG-bcU@_8CI;E)&89KMc_,aW^-XG4HZ)G?cACM^U=[@(7.W+Uc>@
Y2e?N1Y^<61]/GP,\PU/E02c\BN4NBJUaF0cSJc6O?AU;X?<,&><<N2X?YG(9T]W
V<^5JLLWQ\>f6>Y4;#,[2:Tb4[6e;1Z#>\bg>g.?bCU+QM8Q.Sbc6OGa5=0+cG-f
CaW+dS)a8AXDCIL-g^#(<NUN[[11]JT(F7.7d#-R]:6e>(SB8NLQ-@5Y/L])BYZX
Ha:e&&F69.A(^N,1^39?baX-;DXeX#A+O3IeT;Ed4cPb^RY^;NOVgECL3cff(ZTG
_eg2BILaWK/P=\cGU_:]\-+(-0K9;?OCE;U^?,RC8#B?0XB7,>CI<)0O<+gO82eS
(H\OX2H5N/8\Y#5_@F[SZZE25N=\;E(=@[L/,&/X/]9G>P:44b12K(<,U#3YMP8M
F=Z([fA_WPV,0-J<=SNF\B^[R@>IY347W6_GIZd^g:+V5Rb>1Z_PN:&-0,&BASAR
\LDK<(M1OZ4/g@f#&L>I5d@>:OZd@726?<OaT;4ZA62_.BLCI?B^+)5C68IJ;T)_
#1-gT^LX:g/,ZedB.aBaDUB<:?0-T9\65@6a=P6Q_QCBXM;KEN2XX?2)D3N>CM2=
J,O0+Y.SZTKM@&PKXfBL??bU)2aeHO(2=#V3)Tc;PI(-Q=>Q0eVF^&N=e?-I6GL.
B7.c^9T\J?M1>:#[^@C?=fIc)(>DDa[ZPVNRD,^A[5M;)8dW6;Ea-U4;MZY-2-^f
YMYK#RS&E9:E(X17UKE<Q[A)Y77)WQTgX_6BJ6_Ea\E^V\]#/Ec#8.SK52+)[9:g
6;Pd<XXTW(HaCM=PD.;f#g#[c-U(1(3BY&GDZZ:?F@&?^a;2,UfP[4MBZ,U-EVX7
B(dZEd&+FKF72)M+]7P6ODDP^1<U]33H9X^2-Ce;JSG3FE+I&bC=EA,A:aC>AaHK
J65F6-=1TZQE.+c_=]6KfST?MRGA?_a>;BJD7#)80Ve[Z+[eUP;8,b#=:>\&[KRS
O(_M;9DKTC-S^&&eT&WMaaea7_S;@&Ce\&8#cf]>aBc[+WMS.@L/b;GFVG7]>@PB
C6\]ZfA]JZ7fRF8@K9f7)DX(\)2KV]UaDBWd1NgA=)=,6KM8d[(Vg]LG7+L<]?J9
5;/b\T?c;c<K7006Q9[bSEgQP.eO=+L[Y1[3?cNZ(O&B:#>Z0_GAI.OF&+FM+8H\
S;_,YY9CK09N#]Kb;D9>#]^e+YL:[=73&M2+.bcWYC:Z-8?AX_8,=QXAML-=6cY]
:ONZ+)a5I,HK=;2IF<,C)0#]+Ga?6fW9B_7W&;\T]OCGb.A<&g;@FJg[ND4DJb8V
_Q0_ZTE,O)Y(E\UQ.AM3N#-L7WGGaQe]@5XO5<[JK01BL(T4;JSd.JT2+bIJ>)U2
F8)2DKUCIHQ+[VfHEDa&G5G?Q_2H?CW1HF0D81^Gg75@]5AYcA^T@+V-aB_gOSCN
=gaV=OXQXR&#:fV(a?.QEVQ<)9KFMDM->D(FJ8-NR[WZE-VQ<INTY#??]+G.,+4C
Z(JdQOPLdUb]2b?>&PIUdZD@e/)eJ87X[IRXH^?8EMGX/938P/Je6<EO.KFAS_81
M]72L);6M(>16.0UbFe?9L[#_(R,)^8E\:_);[&<gX6AX<3BB0<ML:?[@(S1=aPI
9cOK6[BW3/L/ZM70SRb)fC,BJO\TN>aX5D6+87.S4]Ub\^AP_VOg0^3V?8@6[(@P
BA)<]:1eR6<:<>/+2)Nc;P6645a6Y9NITN6VL\/3ZS>G;^f71^eGceLfa;YGD^eZ
fYcc7\16WKKbcKU,,18<_#eA_NAVXH91])HgFWXbL4HX;453gV;Fe[Z5.bRJ(IL=
/34,S#BN<JJDg3Pe,W:(fg9=OS/C]I-5V]CZd1@_FI53a<eI\ND#/-W3&NJ5JR2.
#GX^A3eJ]:6OF)c1bKK)&R(H^dJO(#JU24V_PJ(<YdY_XBbSW_ID?Z971c0?gKJ:
P\&QTES\23^L/CZ=L-O?a&YFKJHV3QL5^=5-W-gP4a9.J3U/7<_dK:E2;b]<\aJ.
IM1U<9XX1&]G+5+(B3e)MgC)&d6UG,V-\3G3U\9,7:32?#S0aZ_SWc_Z_f8=_<:.
3^a/#SHF#cYSS1,^O=:HAZ;YE<1Q,9(]bQ@7eI4Y)KR.IAWYc^X[Ib;^Ig:#4[gJ
84NY,B9BOGdI)S,J1/<K)(d1,8OKZBW_07X14ea2AUgJT4D#ZgUPN#M]YD<9TgAK
GH=\++Dd9,HES]\Y4=b:P(?YPX,(:6Z/VS2Z9FTS7RcQ/#(2dD,VJ[P?4dLLb[.-
f..Ta_V0#b/6F):/_,cPIQC>G=,#MEJ@aOLFXN8Z5B3@bfQ<@GROTFda(IbMZ4<e
\)c4JEgC<W<_)I&7RYAPP=dgRHe@<E53>c(GbA(5R]b(W^(X6]-DT)HbQ7S<35KC
#RC-RO5YO)fe:ERWS]LT33=,VMUWe/RH/@D:I+NDF0B:U3@:/Xgc.M)()FE.aNg0
dJ86]3,AAd(E;+9b@Pe[EPP&_()R.D&@EB;;DL&3?6KD?\e7OV:;HM45&DOeeFa1
9/3gX-P>bH#d[Q7OGL?MY>AV1N[:-X6:3)eGSLB=2NVc=NQ;<J,c8V@ZN(70,_5Y
0;E)#ebC\P,5L;OSIeU>bLR8F[Zga]X?aU1XEQ,R<)H?FC=0KFS)#ET,3+<_N/GV
MDOXW;[KO#9/Sa9VT=GT_FK[KB]a<A@=Z([>UFERQXO&XSHbJ/NdO<R-?Y9=-fXP
,<VaR_2M33.2#&QKLZDO75G2I3e.2Q[\>6Ja+;LTH[-#90E9&):[>F@)5YHR:+N]
E<S^@@FTIWVQ2LfHSga3&,=g65T5H(?+;JYc#1DY]^]H)>PU1d0[\#7.8-:P(CJ6
P&+^^K]EXI8QZe]WS>bPVg@M/fVaB_c22=+3TVK[&P_.0</RgK2S(f/cD>G;0b6B
fPI<7[G8U-M,((D][/?NY<S0.(.N\P0SYG58,N>7KVPdSRY7&E0g\&J[?8)T7UK,
db&cM=,#NLW&^?H=:&[BVBNJ\CC\I(1.0bF]abTH;e1A;E?U]XP(ec):,ZdXGd&6
1dY53]7=LA;1LBQR5?&L].d2C3XeB7+=+,HZ#U3fN8O7cL9dE-?>24BJ1-cYNB98
(F5DM#6O7EbGQBR35R..U/U;RgfV2FNTYdMba:fLf8U7eG8D6,HQWMJ6^G<5L=@-
d)&C&g5R^FHCMS_]8O9:.[7#/[BXKUJ;g+6cV/2<2<I7Wa-bW0^8B_B\=70RM?A<
7MSb54V6ZSB47BH68Y&-R[[?F+UC_cS/ea)>L4X[RENX7&df2ODE;O^Oe?]]6ELf
^1U2C>.>cEVRMEU\ac>gY;ZO^O4&4&e\J/+a3JQJ7;<_BSP^,@7\\RX>XFX_]A)W
f[N6Yb2MBb38K#Wd@C0gL<0L;K/d5B)E;;Q3_W3NG/[2=[F9(;O@]E\RIf;#KIX9
d.bK;Q.aW/[a\NQJAPJ-bR>G:YYJGA)@-)<B:[71XJ7ZAMaM<CYe1f.;J6eFDUY0
-3DH\MK+HQ.3B=+M1F+Pg,<2N(M_M(G7-[X1:c1C(IT:97A&V=[R;IK)6QC/2/BC
Z=KC9LNHJW=(=;;1JdHeN:Oc;_\Z[]Z]/=J#R&RgC9DVS)MEe^b&b.>)TU.J0C(@
:/Xc0#0)R)PbG#-.)ae,\(>)e42R/IDJS??>O34D/#S.F7.e/VE6Hc^#dQN:Bg6.
/HV+61E.[YESU6dSGDQ_UIf,CH2gB@<[b?D/K=Og#O3,XNe(Ugg1.MBY3VGJa5aa
&45ZPR_&&+.+C6ZD:g=ef3:eH?H0Q6)Hd;;\P[WdS;Jb.K9Z@K?/;RR(Sc]b1P&6
\4<c5&S;f/6TSQ+M].WAX087G-8eL5+BKWH4@Q:S+IbeJY5_a\4J[W>?G>:6aNLD
+GQP.Va0X6&-gc->K2>6]df2Qd89WCQ?F7_0&2YY:_QRMO:bLb[5]+AeG:1#78U6
^C0ASdF9<&,2[T<US0CF+3++SCfT<gf3P7=;Z7OP9D=9-F6PIGCWEa@HG_0A8B2M
:02e<9CbKE8a.4QHFZVIc2]U7ZSG=W,X[M]d<FeL@-)>7#fZHc<C;G?d?G.()+24
f(FUC1YZYb;HKK4=N3#Kd=6X)bTD2N(D&@;U7a<P+aNB^BNbc(<aObIY)fgMb-DR
,&01[7MMe;BBD#)1IZ:I=)_9>KQ/V]ZL+FFON?T]dd7&Q1>OE;SF/b@c_c;K(K)I
d;P>\4=5\:Q9R_)?:ZY9adHX8LN0J=\#f4,\S#:[ALTXQ?P+3QR1Od.JD>b1R];R
\1&(6_XGc:#6,T+FRC8.,VCFJC6@Q&U1[d2W1#(TIW&-c1,g[Ab\..NgI7NK_==#
a;dN4I):T+S\gMPa[WA<AFa&62<ZO2#f2R:5C991^(>T/QD5F.SQOF-9)YaYX9B^
6BE_]58/MB82)J8,YSY04E-_T\O=>fELW^3CGNV/2U)YgOR&=X<5g(,Tg#EHIUY=
e)?CC<Q#I1cJN9eDDZgRURVVffQ#[P.J#c5T(cB7316F;Pgg)dB7QUOg?[AHQ=GI
@62+D<c>C+[V(-BD=d?Vb5O3Dc1F-]/c@c8X:VJ6CTe/8979bK_Mg:eP5EJMg[DR
W=ODG<_:U\7-gY:B2<^@UY\aO9#Ic5B<5Z@3fN9^PXPM?;+2Ne.XfKJ,@,M,R&HJ
M:PT[KPBN+6W?XI;CbINbOE,,8-0A>OYZS87&WI@^+=6U28,V9WYV2?6X;7B?ACK
fF0XIB#&NRc:S(#XaGV)K),H0BD#>f\B/VI180L]Mf^TIF[.GE#/c8/YH9,?+SIW
W;Ua;\TAJa7<38AI6f1CU#HJRUXBbDQ>64+81b/&(f#540FTTXA_Q9<ZJZQ0\L.T
+bfKJ&)4@H7Y>.=?LK?)>((:4@MRK<PC=XgCg>L(&DJc(HD:Y+aQ>c/d4^45[H=3
BY<c+]VbG.CY6@^Bea07Ag]5EcW]L\5-#AKD=V?+a^QFJR[A45YS\:#_-QDa6RQ2
NWMc&8=4D;A0SR:ed;g@+71WEKc_[TB)GV?-2Me1IA6YD?f_M(?7UN1g5EY;_G,1
9VS([)4cdQ>,74X/PL_0BTR^;J#AS0=,W7JLV0]>&0,LTbc?7=If]I01IUeRHC#;
MIX]5VNcV2?ZO/P.[FfE.<dAgOQ\2e8F@^Y[2NU&(8);<FeWd0:N13.FX?a4[2GZ
68#^\;WL@.59[]++S<UCSNOfff\IeKD7G:HE]H)=c6:UP2fYTXc\+[;V1gc(U[_T
O5)6U7cY]cMBI3BVXE(TN1<QTQXU@X>9e@&?R):J=9J/\8W=]?gJ16dVF]+#?:NX
b]&b/1/L(D:(Jd)>2Peb]aS<dJ9I#eEZ38&aVVeXVfJ8_V5F,6:0/ZF5H:EP=Z49
63I@A[\1]A#MOVVLC>7d(8BD;P;3YHW5]GZ]f/\[==@[C8^6@9ae9QGNPR[Z7@Eg
:WUB2dSbP<YE\75CA&SP@0ZRU;576(#2aN_A5>\cRdA&+.?,0Ie]^JDI+)JZZ5V:
41gf]c4,d\@d1/9KGa]P&C=AgHZMc7D-#e+/4RX9#gD-SG&;^f=HHV_0R/_Kdg_2
5.@T:\OO;(,N069=T/\9[\;OaA0[]#SEJ4W<>8);TJ?[A/gCX^\;O/#[O/3_<U:P
FUN,8:_,UeHaF1/PdGDZ=@.ed8&(T3GWYe.VT<-C.X0^V0V@TM\YHK;0,KQ.UTWd
eB#XPe>)?V)>O8=&eWHW8+T0DQ[6c3J\^U&Md1_OXRd0X6U[K&546g3[NE;&SNT0
#NI>(If/SO=1>OINaY+QE2d_aGg/8HRHJOU30Q-L6(O&#I?[ff]>cFg<715C)6^P
eN7:Kc\&G9LGfKJV4>)RE?W5;1IP@311YP_G\B._KcUQ1bd0U_9U\c0+T;3O_&2W
V(<g#^RS6\?:_=XdRI^Z4O\8G5NBB8RgJ-YXBSd\?;,DR#+5UF09-D3/H3@Mg]3W
d0@Dc)O61_:5_3fAb\7CN@.CQ]<FE8E^((Ige+5?RH:&d#0HJJO^_DY]=LB7_<R:
1B2&MHISJS>.eG&U@gbR1c5J#QFDc[32),4a>a7^\^+C\[ACTPZ&1J5]XQ+I3WR,
SDVGX,gFQc6&MQ1XSRGa8X3ZH#.e,-GCJ,+M8J2YWX\:0e./IS512:OWBW917[)>
35=,fYXOL;3Z2\YId_RGRQg(_Z3EIeLfBX\ISc?S#(P]::EFV:]Z@RY@=H).&WeF
FAXL3;,=.,Lc]HD=4?1<_]C<&3:A<5WX]B4bG?>0(dO4XBU(U&I>;D&&Q5C^]^Q0
f#TL_P4MV_^P?G.)c5GZQ-3fM;PcLKdT7?2<U^EGXOX9^#,a:G0M3CGHOFOd,ab3
eM<S3:EG<-8XN+;?WHS?=7=IF-398.fFH:9RNSbY?_Kd/ZV;K47@=S?IX4gOT3_8
7M0aFG=([;9&6aP=/2XA7F(UJ3I=U/[Me(@SNS>(;(e2(Jf>,W5[UVD)aI641c#\
cVWV&5[gJ4eV5f2>JT9c)\/Bb&@AS09OcOO>TK);#6L@W(WS9dI.@KF-cCbY0dE:
Ef@M#16e&/6>@L[eJ<F?2H_D,,=WE,7<46=;;G1ADGB2L2HM5XXgOEJJ5e>JA-.>
NYc7[T^K=&T.b&gHc-DeC)DYGg-2V3fF\SEP06(+)JXe5J(=8;MZVD&P:7_J]6?d
QMG0_,8^Eb^IHF4&VOMLS&Y:5=OEE<#4P?]ENS20?5B;3Pg_NZ/XMQf:PF263ZVM
8#E9,)R^,5L.a3A&(FF)TH)(-Qb<ZDf363&CEKcGAV[94G5<cM[B8;QU=9,Q377e
g3f-c<eX<AM&81D357YU-,&QYGLE28b;e(aP.9dS0TD?F.P?F/cHWN6A\LY](2+0
I2aZAQ&8([.]505PAWVQaIHM5dT]::a#a++1-Q=GKaRA&&S@VD)(cc\L&G8M?M+b
@3X,)C1&_NNI-9_4ZZEVKe(7bg67;8[P<fN[cbbY&QZW,:dO-7BWED_QY/XDd_HB
OB1/.SaFUf-9#,-G>:a\A9_(,6)/Hf5CEN0bF]K@2g/)_JRLaVEgZ<R?gHf5R+Z8
MFUc@EMG5)4XeG_FDSPXPQCc4)f2[JF23G\Y6e?6=gCN>Z>LS/-8=27OF1=6Q/AG
\=2/F0A:V-/a.3I_#b:e#3P\/=Q+T#Y=@#D5OM=/@)fbb6A.RN9D^<G5Q5FP1>?,
GP<(_A23&RANZd6_=B,DXRgW9BJJfeIJ9JRF229(H=0I-dYC0C+?V\bC(J>FHVG(
<faR#@YBHYO_B\5F+EHQ1Pc)@S>P^?<CZKA[9];c5I7-7EBW04PG9Z7GQEC;.8MT
,dcD;?]b4/gb7U;e)MV]?V(69J=NX+GGW[;f??ZSE1.b6FA+@EA[PGdXNV:K)V;R
=IT0b&<c,<J,Q+9<I&P+Nf48S2ScKN3#6X\^O6G;[,bZ45GaQZdg>3S7e)LfQ<V:
Ed;SN2W0,;MBS)c:@MQHdKEP1>LREcDUA)8PK((KU,@9:)@aLX(U+Me.C/HT9fDF
_=SX\,@UF0d]Nf]NfQM&X5-B(T0PTY1bU_?-5D(XW[S]\@W7GCWDG.ab?[MNWH29
&D,734<LE813EIA^PKeFX:^2USEVdNL-(Vdbf>>ZPR>Y1Z73cb<)_)1E?-7+]YBI
LBCJ@?E7GUY\<DC)8OR(E?\Aa/9G^Zb<(4UA(R2>aHOgdT5A2eIa2Ie(HA5V?,^D
CIR0L/YR8U^ePL/(.cF)a/ZV^Seg\T9XS_24+.\]XM:JAZa&_?8cg47R]8:O68(g
78N_6d9NRGa<gT.a)MI,69M@D<aFW(O3)J-,+1&9Y(RdPC@[J-g[d2Rf<e8((M7K
ScIUXU-eW7N6(7gRa+QF,e@6:D6)Y/U,9F:&g5c&aD:=.QcfG-M=]PYgC,C&868H
S6]IHEc2/8SJG=M?;5BDf=Y&aETG8+(c0;(N67^)ZCCgI?/QO^f[M&_B,FNG_N@A
f_NYCgc>8EdTbf9WVYX-TG&K;.7GG0+AU:f4C,<N[]LW1;e<Z2bU0:J-[a\Ya5J_
g[9@L>AAS)Ga8O,0YVM7KCGCHDIK0^[>NZ^@<\/aRT?^5^EbYQ)/BA0Y\S<:Q8GE
<06eXb6I;3LUV6B:La]O85ODg7KR2CPW.(NAC5\HUY]g:?=_ZZCUD4F-XBJU,:J+
K;4eNZKY:2f[d<c(A^&13A-J>6EP7&L#+F9YG>DBQQM@_M9,]:adg@F&BGY+,R[1
9b)V<TOB.ZX,:9=@I_)LabHKf9-BALRROI+84>f=Q#KMJPM0O-V^(XH)DgO)@&af
4f.+^(e+J=3+b0.:46BZT[S?HTSb+5/f@D<N]Zg?.8=e,X),gXCI/7G+KS9V,/?\
>??;2(.=;SJB+?KbKHEJ+A^e1FP?FJ3O>VOM:LTcU><MT#^8GRPB]R@f(5_7H>@7
NZU9HW[>K4DD:W(UC4)#<?,>F#TU\ULB9-&GT]3T5>-IC5E2(BSb8PF/GF^KHG20
2D04:-=DG5)b;=-E8VREM&DKc015-f^0,8,F#=1G28.d#aX3eO6#=IFNGK^9T0I-
YWDD26V/MYA877<BSGP<f/RA:,;BX9RGMH75O&EPWR=VG4=T=K1+Rc;80dQDCK)5
<a-4,4@JRc@fY0G=IbRT?,-fa3QUHDL@_1S;PcgZS1]T_,HdO1#F+OS)_7@W-WMC
++E<[;Zd?[T<OA+?NSE+Yg]W4@]-:GYIgcX+JFO01:HF7f;YH0N;.:HCXbWB8(7:
VX5I6XP+D0@cSN559>;MD5@2M]@IM(125=VVS33LN[Pf3f3H9_X]F_<fOT#XbUI:
E]b,&OOOVB?NS]_&X-Wc#e0H]9bI4AC3XfJ:Y<L1YDPG,>d&C/?WPeNQNVXB?PU1
ZS9;-<E.=J.9==V(]ABFQ8C?_@BE5=\0Y#\3&8EN,K0NCE92O[05&)>e,[6E28,S
,=J+65,1VR>bE1H)=42G;ZNBH@[(5S4E==gUJ)V9SN(>.W.^6d5@^DPHR0a_g7fO
_<8.bMVRE]XX5IF_fP_a^<((N[MP&Y9#ZNMOHI5a:MZ#7Z;//OO4@6Oe=cRF9Mef
D]+IIARD4d9Q?NeXQ<-7c3?8dD&He3,H[XR2>YXVe8RQBU(gYXLL4H)MF9QP0S=(
#9E9CIAWH1[5F5fc(S0d2]Gg_dQJJKY._^MTE?GMDFeN05-b7G)Z<G47L:=KWOXb
IP(7MJ;)5Y[5897G>[,Ma_S.(&#<QAD>LQQdL3KH.R9,G67L:aT;E1/8X6+U_MOf
19g#>X5J\J,X;2/5-HZ<<@EI,K4F7#FdI&e\3[eF.41(][BI42&2;N7PZV:G<U_b
0Ob7R;/.9Z),/)Kee4GF8COQV#Y1T=6b99<P]C?VVL3G,>30:<209SCL^d6>8V9M
<.]b+We?<_>NS,69\F4)<#cKCe_(@V8/3N)gDW2I]67M&/=]ULR[QaC?J@WUJca[
BD<fgCNXTFF[Eeb)[_>1c8/O.U<0AB]e[:\NG=K<358>Hf[5E2fO<6\D0?e>1.;1
1R\\CDF5/dfOeb.YQG#(cBKST?d_CHD)OOZ/:A2<MQ[W>#8cI>D&LBYGU,dEgg5#
W\9Z_JBV;2JRHDb[<Q#D^#/D:&IXPYSY3#OY2SND]S&36XE_SGM)-E6I_cQ-?JQe
IO0?CLRE9F/>=5AKK1A3adb-Vd.;\_=G-W=dPS8YM:K<)Q,W/WZLXC6X:3XP?f@S
V0#LSZ?XOK^SP>1b,cEc/IYKBa4[^e0LY:WbI;E,Lg8c3b/>@\[@<dU_fI//eQ\[
c5c^MH.^Fd_fI-/:0GFaVCC<23c2@>YZ?Xd202O,7?1-\KJPYFK?R1P.,7/(-#.-
NbX<M_];HK)_MPQ63^g99CP7II>R#FeL@_=<U/[#8Jd21VE-5L.We&_:PPFY/F91
X<[UZM;DH:;<>DRc\?d9eB:G=GQJOf7DE>E@>CYC25P-O@47d.^8a=4H-Ee?1gKZ
?;\S38_X7VR.BU6L\>\,f(_]^F2B5CX]d\FT8;J3S#b&JL>[FJKJ@=PF:_0FIJD:
@P(XUNLXR@X/HKLN#4=UE^91.X/eLa:S,3VQCUZ,e@:_1X.N@+T85FEY/&3YV_N5
<3YTLGC</fC2\^;8F-TZ:DVAW4KSD#L:(+ZQOZ[V8CV2_LW)479:fJL.\<_\W+,f
=R7ZKEN&;>L6O,EA<Wg,T6/N&PMN.I&(H37)ZeJN9<+(QZU5GSXbLKGMQ>ZSTVP;
SE#e:QS=(C>9^\2=Z+Q?U-G8^T.Wbf<gS)A[K/HXPCJaJF+cBcc24/;3P&fV3#1A
G><).=W_4fC0AYX>Ob8RI&9^F[V6^A0Yg=Z\N/9g3T^=W_C0P)KNX&36ZTKY(.FB
QV<4GJG#bBfL1(fL>5Y=9,_bY>CBA,<M[3cU@7>/[^#[M]3_+EZ:Z1E<MPDY1ZSI
.LUX303F3MfVfLdOFKX,bG5KF9QL8=Sd>LZKaJ&K:_I?7_4JB74M:c4H1F;&&0M4
#2,VA\63QXLZLT=M.Q+)A,M>1Ydg-I1>&KOc3O(L;Wg?O2O.FQb>bVX/d:a=2M>_
J:]:7LcCf6@89PJ3M;2-_@?P5@FJ1QXCa+3,OB9_(#+bIBSPPg)5FPOGC^ANH@>G
Bd1.?.?MT5]88IHOTfA;JFE:S7[I[fc<2(@)U6aHH3&4Gde]R#.@S&@V5S;MNV-2
OF=)U&dd@6AU17DFDgXK_?HB&P#;fL\@V?D)CH=C-Ya\]@W,<:0+Z\aCPEaV0_#F
GP>eU@EQdeZ#c22/IFS0A07+U[F]Ed,<:(45>(bR9H?Bc/ccX-I.@<BMVa<1M+@O
IBVaS=+XFQ&[8IMR1(/BESDH^[BNZg4]I@?L::&Z=\?2JX\B0.SQ\E^.=E=&TJT2
V-8YRcea5A)DA634LYeF=dHZE4<]VSe/PY<Na(F;^9FNC@R-T@a&.2bTF0TR_RVH
>R4G9IX-\Yc7gM_W?OaNIf8eT7f\^P1HXDUS^D10-OL)B)a<X-:5FGTC3<<0\;8A
_.XQE&TZ54M9=W(BVAQe0Ua@,<,<S&1QUa)(]YC=-IgC_;)GWLKb:BF2=T_HJW6M
-NB\OJ5=CC+PMP(T;f+B8H(/S\.a[Y.Dbb2^3SOB_2C#@(J^3F#QE-?L^BYC7d;Q
U.W93NSRXDDaIWX[.L>faC/;V;6PF_-;4e\-@La\SYPE]]D4b2gc7EaHe,,?d[.Q
:gg0PI&W:)=OfAOMWIDCU_VV2L7g#R5AK[Y/;79c:GR:1.2b115/T,5SRL4gb/A:
S2LK[7Ga1DA)?TRF:1Z27&V2dL=C88,I#(=>YSF#)V3Y.gBLGH4E^:M)VD?;=bS8
PHVf<>b2bR/YD3g@AD@=Z7Z3MA1U:;N^;N4/>5^)4A\4+Cf^P9VVb=O+H7>T>F?1
g4B,K][O^&73+@Z#=f88KV+P1B>g-5)Z-)B(TMVK-/G?ISU6KQ+\D:67N:24[g9)
bUSW@TRL)8fURLLQKaLef.-cVfJUTe3&ZdE02._8=SJVNE[,EABFZ7E,FV,R[RY)
8.YL_S_EN1Eb5g1.V&.=MU<\L;^PcPPUL.,7F&)8AU(8+d8dJc_2445M>11M^=&8
FD.XSRRU-H,F0OJNULBY<C8Xa)A]4SLcPU-5F27]-)TbA-RSad4^U/,KgafE-->J
.&831(;.^,0OBZ(WXH,4OQ9AU_P&-ON/<07/a3,KI1#)a9ECGN.#NX;,?_.+@I<=
,Q\]^FGf5Wac(,&6K60JRA_C5-@7gF4>ZRN7#BcEK#GYP?,X?JSgYb]-RN>ef;04
cKB&H)^a,CN,#J^e+0#]^MYBW+140R/bUb]#]CJ9M7V-5Wc85HQOZHP3CX<<=S<7
.d,=HUE@QE:;HMY(,RC:G;KAD]D5>X/#>^V\=[J9BHC909I?ZXHC<U2a>..->QTI
1/J>KC5BWc@R#J@1=,gc91KJ?[5?(aS.Ug3I#g5>(d=5QPVB8]27f<\?c^U&-H6J
WJUZAE:IV_d\NXd(AV/_5K^)(#bgBQ(3:bb4L5b6>>O(_WUCZBSGC&I6a,0XPHVe
5+[D2FaKUQGTg1fZfceLW961KT@JcQ8F?C/3N4#e5L8M_ROE<=3F-6])3eHc.gTV
KFgWH11f<c\]eQ50/dR,6H(#0OM=Ec9757Y[+BYGd[1@YEA:C6\AcEMX=c)8[(OQ
_+MA>._I5&(b6ETT4&Jf0Z1>W1_C@K3)1LO;Y.QSYTM^T83C-Vce7EQAM?[>;8]9
d0K@ZOLc/LTbUCZYFV9CIRK&Q;S^V6)aDFBVSA?S/3,@9#33Q=4VM+M8VY)3AWf8
NX9Z.OW#bf5b\@TMb.B#.BI;,YN[3RQO6:EH4g8[C;TN]fg_d@AMMH&5XgNSdDMd
+KT(J+BTT;W7CELX\W3G#4ID?MUJHSI4ZDNb_eBA8.O^7f9Q1g86#,45Q<65EDfd
6XLF9P=:=KgH\U6LCbW:H9d:3NbT5:.6_QE?V0LS^gA:]J)=(3B].gY\NDS5;73C
9G].:?]a-QS:OB1/N9,)R&;HN;.f=RXdZdaeeP2RX(ZI:AS(S0QV7.>Pc3B#I3K2
6CIDgc]D2<Q=ZQ2IN/)L+IM;6+7<&/94;O^.2T(CR@BUE;LbSd4DeV:4XgCJf1LA
(_]GU(d&ePQHaa]70P8GJBQ=TR[)\6C,M-.MRPFT@I;7>@c4M-4BEY-9(\OF<@BS
1<&SVJ1_AdF3Ldc4VBG4\Qc-2MV(-Q5V87CaJU&729;ba,YS.,,_],V=,5>+BT.d
G?:FGW[D86Faf8&2^a4,#R<cAH-2UFEFGUZ&PZH]YJ6I57D;cY]&=Y6C+CFB5R8T
?c@d.^;(WRg?B<dL7c,TK8Z8Eg(4RMJW6,.LUcEcgE9GKfKQRXDb3>)44S8I/c^)
f@9[@<,^E2Gdbe(UfMK@/TBHf;PT_c=X/Q>RLW);^f&/Y?)1<WSd[[ga94O^CFC@
.BM\2[YP#gb62\4<2CcKB&7UE14K5SaKdd1#;LNP-=[/7d2A14@K9a-Re@-VZ<\-
E@I6\;.03cHZ@f+S,O3>ZRGH4W[CQ7&f6Ia)?De5g#-W]GbgU6RRZaN6[=&dY/WM
ZX@6Ab>R.(bA<9BCNI3?)9X,6B#+Kbb;gRR4GF2]N<Y#J8OT6;Z3APYC7^;c.6U)
?CM<+\FHgabc?:U^V<Y,0U9cM3[.>P\Q6PLZZG,D^/6R,\_L+Y4&bUD[+6c:;2?1
fXND0VBO/0KHF#OH:@J#\&&bVIK4JW.Xa8KHfP+J:+TI[034cK<FY0\58=ZM5..O
KE\g5T:9X<+D99?YcdEFE[bTX>YQ[-,_,DTQ1d)U]4M<=+9B_O]UO]]4CQQQDN#=
7:7_VY3@ZSea.,d;<>ZZ\@EB,>#a31Cc4P3[?P)[)eV/G4J3Y41S[<B.C9f1^>R;
H(^gc00,P-\@PYL7,(8c8I)T0CBL<8LLD-UKRUV^4/OB7^+#fWZ>dAFVIOG+WX4W
U9\,#<bU2df;8D+W4IAF.9N0\HK33cUJH;NAS/M6UFI<MH5^2@P^&D)Z9/+WZSNf
=XA>PVAM&/8?B4UBS2e1N,<,;,:KX&N-1Ue-XECL+ICWM.ZVaaf=DG3(RPZ5\Kb[
759Gc0Wd)F@RYW9=fBa32@P=9+2I)<]?1]BI]_4+&&]SR0D=A@COVQ5^YBQJc&QJ
POTYN:Q4fO[8.cU)N5[7HH?OfA_.:E,KJMBIJ,d+[9GLCPbM8c-1=)<<C&0ZYEdC
1.UIe-b74:V5aI8@2eeR6]f,05C<HSB3/Ga31I)O9Xe@4CWNO>b+0N.K5\Fa.5EJ
ZQa57DA^SXb-,dCR83X_A,W8DS0aU^F&Sfaf.FB@N/8A^gc=a5gIO[BJA:0_gJ?7
@(?N;Tg)ADaY&@EFNF5-/H.?(ddYV_ER8WOMV#X#aG64e45QQXINA(Q?RIMb##g@
8CWM8[7Vaa0+Rd[H]@C2T3H(YaObJ@(??1c:I3@FK29fF].c_6f4P2UNSVfHZXYV
;(<\bK=-+5AfG4SAa0&937)&#HD8I?P6GAV]&C2&P)7K>6e8F-LCd-@=>)d:e?<D
a8P>4^c#&^QD&B;Y?X?#=,MG5IDXbH\0YI/AdH>B_2d4S,SDPB,-);@50H(,MW,>
KZR18D+6>BadD(VQPH:A7BNGP6I\bcMA&gWW8_^J_7/7,HKRTS8.]^aK50^<XfXG
M74T4aUVd\Q;&,OVV\Vg/HLTR#6bN+_5U<bV2#Z-b94P>AB6(:Z9fg3TS-/G&CZW
<TR)g_5#408KI3IF@A&OUHCZBBgU0>SR_cP;b)P8PedJ/3e8^@Hg\FX0G/W,>B=2
WVK>0=-dBE<e]RMC#-C7=LMZffd>Ae6-5F[\9:0e4Q\45?&+]KEeAC2G.@Xa(.PG
M#(>a6G;EF4M?U9P4Xb#@H=?GBLd3VV8QB,=\9YacL?2]SIWZ36TeW\9G[IB10E+
,1-0NWT36+EP=;3-(3g.Y2?DHD?+P8S1Y;3L338^-e6NDR-MCPfX3Wd-DgQQV_IZ
(Ng9D=d\71I,TX^67dW?@()Ee>#EJgP-d4^d:e9C)]=F\][8J,JY56A/[W\d(\]K
0GRDVa-H[K++&Y<[2+cD.T?-^S[:(=?aM\IfI,1AMA6]-NU[@)c/-_?B\P7[U9X8
UOg(4TT:Na:5Ha1Q0-c.e&aOK7FQWEDf]>eX1OMQBMR=O[Pb:./Ng)1<I#c6+ZTG
cHgA]2&4VG?_+.008Je=VD3c\@]EV.W-(RGMQdcZQfbA)M\1PH)&_4PW>9QH/[E\
^@(1Jgd3-PPS@Q3=PV03WI^0?N.d?OP-18/CN8+LN<dRcIUZNV_>R&J:-OG@DV))
<46E[_N&<NAF3Y>0)E-O:1c84=4GA5<\QP.N@G1Z>N,W)KdX?cNg3Yg^L9b;AER#
F=IA-ERQ(D4\?XIX;4NLFYS=)SOR)TKH#PUZ_=L8MH-5>88P+e;]Xe#9>I>f]#f(
1R7V1?>17Wd.?Y2N<g^(OPIV\Ed)^YCZ@[?O0Y:dCbHX+)Z1S:VT,ZDMD.f[\G]e
Ie6VC),<GC[3[_6VP\QNFJBI3-g,50O?@[/B1GJe-IUQ0XS&3Z(3U?bePO^Gd2>W
+1I4#f8<g:,aCUgOK,[M6^+[2[VP?=4=Q[NB?4IOP7,5b\B8R+eY[SF9L_3J=GX#
3^KEScIB9b2=2:^\V-WFDOg#DEae<2(HYfV]Ug1LEU-dSd_7\BGa,E7HJTGN+6Kb
/Ca/K?#K:PdfGS2C/PY;G_P/EJdWP&0;+9SFgd)eO0]cUX4V=MY\[bQH27VAP4f?
E@8\9d6VJIgZ@;gFP^90&V[@IGM&SEJ9\M:X6YFAbKXX8XeC3]UPVN4c?GdaAag\
\E-C+SJG\U3aX[4?QScA#P[[EX5=Z)a92dOP[7W:JE<;K^]X5SM05=8U@+M?<af1
W54U3e3#:)7b6?KZ_RIOdWSR)7gNJ440T8.&P@/Q/&c&\PWZ7JBIM^Ffe/Ab4>M)
a;+NK5RZ_Y2If(d]RFES&FX\dCWCE[:_T_-R9I-aUVEZGbIE27S(0GH-QU_5&fN^
G&:U\eHNX;V_-YYT,?[STOC>,?X7g9JACD[BU(:aB;b)?:fM2bIFQ1C#ND<e#QKU
94=E/UXX>#C.8QSPP;;bbIL3_GZ3/7M_dE]YIG\dW1g_LG<MFR-4/?DF7##dc_P?
,Q1_f1J8N90:d_-gg:MMK-:B;O7WU5P,dZH7d,EB8b9F30YLF0<AF8c#AM4&\\95
Q/U=TG93I^6GY]KJ@^/bBEdYfW2KY=PR;;T]d+ZMY.E)&@(_Q8HAR;d5CV)0K&C/
\NZ_/-KBbe^c=@E#CJY>e_O?RZQXR7^BQFa=UJYKCJ2(d2CF6g\)+^Xe=\M8CO2E
ADJZL2//;2=04/DQCXU^<fY0Da96AWPWQQ_IdOWY:ba+09Z_Wcab\_XYa-7J0dXS
bc)I&WG<7V:_\cOE9:6EPNa/cKNET+aB\2V&E@@/XI3OOeJ.OV_4A2-/f=&8YYX-
]#TgaLE#=]E#>KWAU7&=P_#0SAVU:E1Q2c;#DR69)#;YA9dd.)OdO87W\ggJ)a.7
MF@8VV,VH411(;?\c@M4#J[.G87Y3OA/NcI40:6fLS]@fL&JS-N0#\?6OdEed:0-
dB=K)F#PS)9J(?8IG:J-T@OMFN#d;:F>HC(0^NTJeW11,_#X24DR;Ha3E>93@)F+
e(d7,<A]X9fFUG\++]FCI8.PY[UH0.0N(&\5;3T&9+56U2&d;LR@B\fJJYJHB)VX
ada7AJ>?>XRR=eI:8d9,Ig)7ETL4UcQ[HH:I#)M?8NCN],-?7KYfZ@M#Q;O[GKKC
)3U^c0C^[8C>8G80S@-4W)FH8ZTPd+]Y1Z[V,@6Mb?fC7V,5NgCT[@e4VC&L6A6U
9eU<TH=\GY@Kfg?Vec-\:UA[QggKC?4Oa41CDT:3Ec?0X&#MK^NgXXX=2e,@?7Qe
f.W6N</4_@>9>M3F9.(E\Ue9Dc;,gV4]B9<+]EE\7.7dO7SFgK2QRUI2b;=EP>4c
aW?LY&E_S^GMK.#6PUI6>74J8#(8;/)/c6DPgY39\b-/e0H7_+HE4&G#cN[MV[C&
HG>^I2WHL/17&(d_4T84.B88QKI:^IDT>Z;;NRRXSI(Pe+a,2B=EKGHNNM1T2]9g
\a9;5He_PF<-Za=03FY_gSGU>9][I0.-B-,LOXD&@.25K,3&/K3dCADY6F)XW9>.
2S]DV@ID4DDRdN&CV57eRBY9W&#05[0K+>I]bUK8F_>MG28^.061T2cB9bFKO3.8
LS:>&QQGEa;(c(@-fF3S6-bGO_C(H;BeTH#;.Y2^b&ZI.cV-&a\C.A:/U7>O3)Tf
#N5T#PFLI3PV@fA/6HDbIAZ-fb_\P?)e75\.JE/,+.0Q@g[,R^89?NI^@9B]LRJV
&HIPQZTg9cgZ0?D[9+LcRZ6PA#/6#-ALC4c09AKP1Ce+O5D2?4.7P/9X@=]9N2TD
CEUHB]-fEH8a4/6GWf1_45H;g?IeTc/a\HQ31T@;Me5g&?AW)FW;aUd)3N&c0d8;
\ERAgG/@=MY(>NRcQa.W:^^YTK9@^6b+D@3M7LTJ[RBL2GA3NLV_DgNa7-7N-,B\
IR:(J;=^_-\g9#R0HbQTTU0>92-3,^V=a9^H<6JCGQca4a7Ma;U)A.=+9+UK8VRP
Z@30?Q=bQ&OTR)d0<8@?5=eLMd/D82GOB_Y^-dA#IW;((KGX-,[2c^&HXR@VcIQe
-8cd1e;9H7)cS5,1SJ;+e)G&b3=)L0S_JEUI0,<#46RFO,#2Mc[]G\@:a)L/X<@S
7fFO#I:I?UK6G42]V;G_#7RSDXOW=NQBZ+AM@bS+HR5b8/-Y<gB.)O,Q.AU0gWMI
c5O.-8<XX+=:W5WNeV):MM5b.X.KNT-f09JX0f_?d:0[/ZG6Y&>_XW,9_;LZQXd=
/FMbXPeD1f13ee0B_)#&=8CG/A<1:#[#D/9L5SSbc=VJE5YH_R#cW.gNU#8c=FI-
eRK>9H[\3)[^ec/^E)7EeRDKRGT]/J6f5e(-Z;S7JO2Z_-K?.QQF)2:<TGSK?8]S
B>C2WVK7Q#0/&?aV_</f^MOJGY\USM[E?1E[QM7VaAf?)6GMbc71=S1^<GU)RcB[
gbWZ:d:H+J3,,a0aJ_3WAe)Dd>KLD64K]:G952_b2I:U./SJIa=&WZ6+4e40X^:0
H5B#M;8aaZEAKg3854<,QUK,_O,V2EH#W#E(^RFXSaCT0@HWf;DBeGGXW55Ag.Oa
aVB<F/T+XgXV3MMd)/S26_7.fSGMg8H><LM;]Y;EN?<e:Ta<\JBa[C]Y<X(9V:7?
ZU2Od4:WTN7aRHFKD@3#IY?C@Ed)d87^.QM2HVGXW@@_-bC._(S1IH=8d>:WXFb5
]I/;H0<^.ZcX7.DUCX:E::Ka+0OI8-Q;:NaTN3#Q0D^2KMJXDB4@RG9DX1=>\0V=
PZHDBf(]N?37.2\PE^J?2;C[KKZM+[#>e3O4]D;HF(K<^EG5gS?>UOOFTJ,\P@W9
NVQ1PT(e?bY>[__/VI[,7/4.@<F[-/GD,(9/&?9(f=VMcafWS>57JF;c5W;?LO62
2RU>U]0DfOA\a,g)3^28V+U/HNX-Z?,PSZ5W,_&F6Z3&GL^Aa2B-Y&#@5V)e&Y95
b1C9C3SDC?E3-Y>#371dF8H3\GNS:#f):(Sc8=1B,[G@YOHW4YP+B.6eC_-A2dC[
]L/F\Ge1W/;;O)31,IOICAC/3^=P\)JJ5>UdfFe>FJI=)6>fOg&Z/+@K)g[@Z=/R
\f2QPZQN:+O]D/<@+M\SYN?,/f@=#4IKA9<88BZ,?S+CFeMF@#dO=b2/eSUfc@#Y
ZA>.;7YO>+e]YM9/A6K^_CG+&9SU]_JP:S@3SKa)9\-PFK6OWWR-1gQB&TLb-81^
d5[KW_5OZJ2;--Ca_@F,78G5?=?I?+O7NGT6CL.L=P_8ad/5fR]\aIUOXY^_f1->
Oe2f\Laff]I__29<I\73M@?HR4JICc:^CSe5-IPGQ8)+[M+KY&e=Mf?5Y[d6Fgb3
XG?9.;UH;M>)AbVgMFSVE38QYg<7W5;K\b?G;7Q?/>:Q#adY[gM>A4A<KNN-_cCZ
KYWc,4\LV]J4PW;TJUBaZe3217)#O,K(X,_FgY,CM>^;:(4/#)GBW\G19<KGVc7?
G;eZM6gYHb&U5;Ha@CE(=IK]HG>U5_UQA?b__[:aR6bDEM<.GL\;&&c]2AcW:?S7
:J9^\V/@L#0>f^#66\-N?gKV2?W&fW1<S-E;;XOTF<.I9=eX5_N7EH3QSD<6OY0f
,N/\+\0XcX#]H1C1dAcaI;g4)Teg1<D:H>DIZM+5WT]GL[K8dP#dD)\c;e;R]NQ<
+7eREBe9IJaZ.D3@\2](>UW/-<2ZCC9-Q/W;1eJ/M8[M#1<NH.Q[a:HSO8gQ<c0C
#.6dSX5J.<J=7S;f.HbSb[aAW3T8:G.P>,^Ce3IW2ER262&Nd_<ED&S?6;;8.R0d
LJe0eM^OET;K;d4RP>M17<BEFGG6=H@,07LQc)K=1c3MX4(DOEcCJUCd09,Ye4U)
QPYVIN,(A)D1W[F[>b]R&5LQV2cVAAF1+&ARZc6-JS\1?ZLY^U]:cTJDEVgM53N6
H,\UeP=(RQ?A(T+Q+YYa30S]\NH^(?<>eN+H@T#I,P[:\=KO^KFa#[E)7J;(BVK1
IPKM-Y=g2CIfVeMPMUZE--XUSJ74ST6<gC25+e+N+e>S6,+(N-U)X>U1T3(DL=8G
OJ7:Z5NB[g:?]CIbABWF@GP]UdgeT.TaOU]&LISEW)]_bK)Zef,D>H>7c?/MIFE&
Q5RG/IDJd;AQG<6R]14a-J,+9c;DeKIb3#gfb+?53bS#BF67\AGF+Jc7/6#N3X@D
;W29Q]dfODXF^)+.QB?OH0QObN-:@Vb4D#fV\^@P>VAL(1M?IXO:\E4;QNYWN?D[
Q3V1XaVJKLH;E>25Vc>NJA@gf(/J:V+V=?3^S]QV_E@47<Vd)(<O+.WccZB@Z4#Y
+=^(e?UNTY1.7Q@U/b.(\D<LZ7S?^4YO9:8N.O]\N?ZKDQX<FQ\7U<Dfa+=[?b2[
G>SKSQM;[:30Jb69(&>PWZb^F[W7^0dQJ^a+1\7=D=[2BZQA>1<:F:b4?MFK1_^6
S;BcW7IgGYZ-Nf(D/]:&07QLBaeW5#FZd5-N+OD-RFKL+,;ER<6M1FE;>cEW.bB^
BV,=A>G</@)=4/@KaF,P0TTf@WYQ2U@?,K_24^Ed/H,D&eH/Y8fNO=:1ZA=0bPYX
UW>^RIQRT8f;\&e7#[:;F=@b5fd(2PU>F:8<#:KJ.OCMRWGU-f,M4L4[Y)_?4P_M
R26XICL=A+)T#N.gJ0<8QHGG1aQ0T^I[N))?WC82b2=0RLBGMN0[M8Cg(@_7N;1.
@B]CGTA1I1.>1K]_:@3,#8L?<\683?&]1<WVY;cRI)7R5+L8/^cPQ(L6\U(FT,dH
@7?0\@+IGS>fXK7eN\XNXI?C(U+9E_f>]TeF]c7c:/+_TZ/][/@VP(.27+O.>e,^
>_/J2YA=.7+TEM7I]]C_JTHB>e09DCTVMW?5f=dT>^-0;AH[TYCXI8:dWAMTV>NM
G@3ZD@(aHFfLH^1(#K8HF_?XN<#X1?93(3a\g.82X.<(-<5YYaILB<:<4TNbdZKL
YfeIABNEJS)1JSg-=4&X4e7^QDOUAC.)BbYbdRXO>#NK]B,U@#8;)8I1I.S0HC-W
bE[2;8c4P9CHa4._8[[TM<7ZCJf\].6;[TN<UX^TMZ(>I<F^^NV?GQHI,0:B^NXF
6=#O_\;d\V\(?A4R^-[T8+3.NQTJXKc#T;=cQ=F=VZ]_SR-N1P;>^PH-AZ,7NT94
-16QT6OLX,YY45JIcROE0EI2UF^-59Z,(Y^LC0VO-K+c=ZEebJ[/a2\I[<^R_,SV
Y1L3&PRL0dZbSaK+:NAR3)/P[4a):FGNcacX9&N2e\#]-UU/8H3_JHf72RB,V,7(
3GZ\.BaO,ZDYD2MQ5GL:)L+IAKWOgRSW=NY2_,(2>gI^.WV9dHB:]D##F9Cg,3R(
S7G0\85HA3ST1>+;V@S8OV<1a=_OeM<1+&D04dY3@DY+GFVKI[;0K+H,\FPUH7I#
>#8(DOBXcIVGM=YQ=SH@+4-gR?.dL:aI9FC#3\Pb-(SK8[GKPa3PE):LJ>6#X)+B
S[\I8OYIFD2C:b(C:YWC5Q3Hg>P97CULZ+Z37?6Q^<@gCbg55<NYBe&SH75(Of:.
Z0XSQ2>9Ieg9(c[QIQ(^a,X;?0[>;&N9&8>7QPGH356<7-_]+-A3We+.Z?RBB9U>
:)+B08/P6L;a36-g@gK>VN&T@E[bFSU.MBE-Ic4UOe.K6X;OaBL,UUCLJfW[e01:
RV6^cEA-(KDV#F<OH2VGL\N5\;+1NOH[MWg4@-ST,c5^#?a=3TO:bS<2MN7(_]eV
1dN#,CdDB^IBS\Y4>WIQ+6QF8=Qc>N4E9PL1?2S/_G8/JL7LHY4(GDN,A5fd7JD:
d,]CKD3PUReN8V#Y]a[+/:&2H<aPDINRW08Q;LH1^K?/@V&P&_-\@GZ+/1DG]+0&
2YG[R0(^H=UY:EX>5H73R/HfdHg:<G&V_[#+K/+]2>.Q;6&6bCRgVLg##,Q71JTE
M7e6D)1GBZ7]V&33g:@#UdMXE[U1O5&]A.FNQOK1<U]\OS3;Ia;::,-A/&?fD#\:
\7cLG2#9F0b?4I?+.?fJYb3;IKKP>&ON.#C]:>bJ.?2R;MO@=9H^&4;T0,c;(+.F
.FB/4C_88)TH<,C,Y0)C=D.RcXE9BNG=2^;T[MQL2ba3ARLG?RH2W.APM,d,:A#f
>T]+YF??d-QK1fW7bS<?=A2H_#g)2UE\af0.8f/.H;>BLC^D<Yc0E.R[-IBIa&W/
=LSNHZR1Q]GGcI#[P@:EMM4ff=;^NFYO3U02@f4Z+/gBF(f)<7gKD6@2KN1[e,f,
A2C&LdF]ggJeCa4<N:PU16,^D=S2I9JE&D(VXG9UZb>PLg@A#IN&,e1ENBU:1?>O
:[LI+#KgDc(^+LSc?c>24Y5=&C._[7-dfe-PW2A8L;XREB)FOM\;(#^5Q2.&K/1K
D>:)?56L&SHPTWCPFeMD#f.M]_M)^]C[R6D=#WCcPXA46__0?F=Ff_Y78\4@[#>E
6,)8eK&LN7c\;VNbFB+5TM4<Kd_gf,Q?5bX06039L\7#K952,U_MH?\c:G5O\9O4
Q_#(]J8D[V1P5CK306H@fC\RX;BJe_PdV_S(gE0L0;][._cETgJF-J/:?^A=BUH/
A0J4(KT@XY4g5/[abAU&0(9X\;)3\Q>dDbCNJ:,RfbEM>>6Efg[?B3\_T#<7UGP=
9)GdSZ@O6&29Gf2R;Sg8We(<T2#YfcFWNbB.?I;PDPfdaM]2AI];Y+D1GB&6e5db
ZNF7Y=W>8c4@cNW7.@YWOTHL8&E(RO-SL/XB>6V<9<Ed57f5RJ0L3=d\@DHEK(\G
//Ke?7D;7TYWBOXB)e:3\+0g=g[_CC/9\\Wb=dVMF-TU+c?c+TL[F?_Z+VH+[H(O
/\B.>Bb)NXV5AYc1e6P4;3Q,[eT_[T._=eKTUOD[B4LJ<9EBdQ0&@Y-EX<3d+0>b
4<<H[HdJ7)A3_U,f62(aNKBd,T&M[@f/McZD6=3U::JN5P+>.9N1gOV,[VT)^?50
<#3H]\cAFdW-/-(I5BH@[RSP7c(_EXP\XNB2K9D?6J<0\G,RW)]2V;Oa+PWR;EJ(
Ie+E<AAZ#dEH,_V9&Rafa8Jg^2de[;J:Y1F)]a8W;GIaH-ASBCbJ3@b[4BZH8NPM
Xc[1EG)bE=]K<3DPSC^P(SS7\V#AJ+(D5TQ&Q#cELLFY=V6d]4H-2,a?Y1dQ/G88
NeT[R/d&5U3^2:9A<LHA&8+Y?-YI;<NWb/UPQ(<g[BQHN<<R^OU5g+3bHU77>OCT
[?.Og#WLDT;5IVOD-6J,:Q])8DWA2&K5)g2ZGT0>R<==<9#O362D;X+a/:9TY\Je
ce,#[9H/bYAc&cSbgCa,Zf1J2Z1dZaCdEGYUXE1D=5K?d,3;W<PeCI5C5[P7]ZY3
LR/YTE.,H0L9Z@[:NHV2NQgd>R6D44Jb7/TRD9VH+0THZd16dT+\#Y31DWNCY7)]
8gLP^0Q+R1GA?(<;].U3/9A^37bC.90E+g_+E#-Q]EZg^6dAW8.9=J>#b7]bGZ(2
@?:\9_fAVG2S=R=WbM<ZeH1L=+VaK;1B3H+@V#LYe?JSJ5DRR@=6)I)JM<MY]3?&
2Y6e9(Bb:_]U(+[O7;@;gf]+a-CC?O<IIf4DKb4VJ0B#O.YV(GO.CcBK>PL?_eH6
6)cW2=.,\ac+.a45.[JBL1_/.EdZN2F@.-E;D:&e_cRU=E-;fMYCKYIfG6)#F(/0
+c^39#Z(c9,OR^F=EATVRR.bL,b3]VZc=P](Z&502/&R3ecVCFeD5a-eW6G2&.QD
J>B?&PCX-N\\)OSP>D]TfC<2.)Y=)5GN\eHf#QZg-eY_DF6;GTeU[-FN(:>H)83(
T26/.V3#U:=@_[ED+F;/N]Yf;FAUffFLB?O:,U:]X=9J.:4bX/IJE322LSI?4^Ed
F<KdaYHI9C37995M+=a<JU@gU/F#34bP,AA#U(66;0e=V#,.(D5KF&&;T9&We-CX
;Rd\9GC@:XCJO].8B85S>QcQ790B,U:[9,f.XXf^,Re9=b2gXXK;CNU76B5^://A
^&gNXN8;X9HDH8/U_(X:U0C.,\75@_W_7[7F,&>eeF2<I(&adK?Cd8aU[]:Z5?Mf
L[)^;)L]Fef]<W&OE3fMHV[@HdL3&N8Y/d5cTB3W8<W2cb?SE)J8dE5S)G^Jc@\I
8&g5I<0VGYZ9)Tg0GPALA_5e\KgK9c)@3S[;I@QD._\5SbEb^JJLEb6=F>a@X7#=
bKb_+:E3(_HJEb\DfY@O?.b)GA93e0/.6<J5RI)PZD)RECbAD@F95OYaW/5W-V>P
ZN@3+R6M&9I\3KAI+[Yb(=9aC70QKF4&+V.MeBbRO80\33<fcFC2IXG+P.bW6_fQ
@X5cBO4U_,eQf8KQ[?0cK90N:3XG8ZQ5eDIW0BO)146.=R=C/M+:?.ZQ;^7a.DD8
+TK_>4Sb&=g^A<VE90DX36OB_PX:K-@gCE^N/D(6B(0=aP=gI>-d&/V=_YTH>RLf
9F-Ccb_#/Dga<dWWUOB+f;>6U,,KfOHXg#P(M,Rd^YMH[DREC]A5PPRZERD5b3&.
/GLa1fN];6,32^S-.U6_PRf9T^&g;OWS6)9AJ6#Mg<7_AKKHIRUgd&0/PX.:1;SI
47TN6#FW/-OL+[@Z?YGFP1e]FHW-6D6W^2@..@:6,,OEI9KKU<Bc/50#]3JN6bQF
LD&GMQ#^5QGR?@:P3^YS+TEQQ8cXG)3:T/6fN=&I<T5+@H(PP_:FR(_TCcHE<+/E
S(&1_GC&<+1<9(3#,F;3ag3#PGE6&X]Q];?TLNC/0K<9fWLOQHTgR?KK;9?fW#3P
fWS_>edg(O-?,VBRHA9+@NF5e4eEZAPVRKd;a:7eIK^K#:X.GMX0R24R:/b\<-C[
SPJGXD8^?4^HQaC(HJL;+@/:W(6=[C]O8/QdW88R[,-f,bZfFc\2@(J.8?9gG&K5
Xg68@47&E)[],]1(GeEaG;:[8HV&&MUJO28&#IPUJ7]G.Ed7.JZ\38dEQMJBM[V\
d9U^>VH17]TXLfG<RR-Ke_\K6,?V(?_D14R?Z.e+]+]QCaQ6D^Z9bcH)K4A?D<>J
.70F[)U,[aeKf92Oc8UC4[\9fSP[B@-Q\9W(:BQ9YJ6gGBc8;8eF9G,,b-I=AaDD
G4ZF:UF]QO,:K;E^D,dO3cY0D4L-F,cX:,;;XUJ)/2_)/88,T&V/;g;50[XTE@7#
PY8TV)E]@URH=[#/(bDJATCf9ETLC:P#4.QWVa;WC[=7;4W-,c[TfE7AYY@=EDP9
?]B4G_gFTXe4eIJgRD6JYeBVT_=(U1D_RfR2=C)1I;L&PaA?)@[/g.NUIOXe^cS7
_C;S.YcA3]Ze8[>(c#9TCB>dW0]4^UWdf4_8Acc#,A^&V-C8-C)d1>a@<@fN37Y<
@I1YG4LeUT/2/.\<^(BH;V[7[5:8)AcE9b1:;S=e3@8-).;2)3_fVZc;ADK?QII<
N@:a9#7]<;=L99H^8ENUK>JV54>Q&0B,;_;+C:?CJN2a;&f0M#XI8>;5Z=->e_UW
e:H^@U>3fA\\d,N>XHFK/g/QG@[W7XQ94H@;&S<Yc6?]7PVBAHO7[CMC3fW,0O=M
KZd;EcdF9HR8#ef0T.dZ(#_:6):3LNa:_faQ8O.=2YDf043ADBb=^NcA557Q-UK]
F,YNFDZU?N+MQ1Q;^A(BHP84<G3_U^+P.HeeD9IYKB82L3N^Xd(gaT1;Ea#)dK\,
bf/T?5fD,e8N_QR8GPg1&)NX7ZJ5VO:3=J^O)B?[?U<S5XE:WECPER6V2#0>_)U4
.[\>,4W(A37HVKTB1abZJ;JLM1abK/Z36^1d&<MHcScPWd-25.e[4Y+(:8PZHQVT
Y0R5=0gEc,QXaH0)S](N5]KPCCgHaS-MOPbNEEO9)F->?<(?1]&>e>Mdf:g9>S[U
?=Q1:Kd=PLOZO,4U?.+_dWVJ(Z+<P1==HS3=CNUJG,GJU(X8+ffdU4I-e[>8M,OR
NU+LS&7LJ.?3XTC0af1T\Q^M;];J4(-2VGFgS2T_T3VbaEN)+(09Z2Ab-DB_[&:1
B5#Z_0(A02M]&ZbRU-g-;4&fT<QCB1&GX2<bYF\5_10&Igg(+fADYJ_#.dcDFL+d
-dSe8M[aZ,6&KR4M5M+gUFCRL(^T=M42FF02_8RG,L1](&8FWfC7OH?fA9]^:f/E
8<<Cf?S[YIB&JS>IC191ZN&?c^,AA;^C=,<][D^EM?TYb,e(H?5N5=_4VFc0YC,L
#\U^4W(I7c:.LIPP6NDEHP:CQd##A=\d_U35LI)UfJYG3Vf1ZdGR::Jc=#DO<P#)
MXPB=0Q=OEB(0NZ#V6Qa=5:^d/Z?D__C\GdFZ-\JK4U,GT4;4AJ8<(()JKQ&UBF?
8:WET5K;Y\8W<e556eWFP+V]66J9XE&2:WLS(Td=KY5X=IIM#=2eTH<J(a,9>dY0
A3e_-X\FV,VXDOJJ8N0N[X//;&e1EL-dW(8d)J#O\R7.B.5?JBadH+AT>>^3eR]F
AB[BECU^/=L[fVU+LXO1XbF<]AQ7T.YJ#\e2AO&K]/O1@Oe3,KSP7=DaIE.ENg^^
>)bf-XYbbLIZ^O^ab5>da5U,2^(WRg5A35YFO_VXN0W,M/L7>;dX2&FgHS6VEC1F
_F5EX.;PJVW9:_#.=cR0]B9+K:XD9(:FK)ff=g__OJ&QdZgRa;Ma_O4?K)6LaL6Y
H>GbUN(.-WCgD&G]WW;6VD(RWWSN\fb]0cf\DOHM#3V8-R&ZIZUSTg(d#+acRA_]
]]NS2]W^1a22adN+B,33JGN+9)\d14N4^.9cS,VaH2[(gGN0GO-4J1T>(-DR,;K0
(gbY@Ze[):1L=@4QA9,P79N24)23d.4E9#_LgJ#AAWY7&\77+8M#T#B-.TM;IWU2
FDfRId56.K:3IQ,ASD=)>LW(g2-]9B45T<74f2[GY3N,01#@YJMG^HGJ@2HG<R?6
a:TK(_3eINM&Xfbg0R2g6G)E,D,U]=6(BL[J10>4CeDIB(e:f=PbF)L\_NOF^=29
G]XGL8>Tb0N.6b7L+=TbNLMfSI8/RbDF7???KSUa3C#-4b8gN6I/-P]J#QJOO/b[
71a14d0/EYA/gHOZP:Q4fPPS.CB4+F77.X=cPXZXKZ=@X5DOOP;X#FSR72b2[(=Z
<=aS<?U;_2cV-^bR=R/Xd]G+URI;O(.>^P&T6]Na3+.74XS30E2X-eg02:JUC=3E
7AU1fZ_>F^dc)f7(^(7[IR.f00X=U#CE@6c;2N>XV7X31M(:#G05JCcT09D5O\CI
SKDQ^6-?&TVTXSeY@R<YAXFAV-9A79dPA1EO?Xa03ZX+M-M:8Z=/3=\2SLE44.I;
ZdB(LdM_RV&S0bNDRR@=.:,)b#29d6IQGV,_FEIdGgZFc9e[8HHP9OG=Q,T#0Q>:
T\7a2>4RVXdR65O=PDagPBJ-fLJ9b\D/(O50YE9U<e1f+:&^V//PNIFNJ)U(A<K6
71<KeN@_If4CMHY3>;B(B35UfVQ9_F8Sa6dJU1bX/[g4?gW]#HGU.?RDe<LLYJ:c
^RAR[?N)0>-V/C(34+6@WcUYCUSfL51#2#B.Ig+5#><\(a^W(69P4gHMU(?TCLYZ
(C2W9U26K18eD[H8S]f-I=;6Q3.HQ(VLYU+O?WE9_\R>/Z?T-A:1FT7QBZE:3,aX
.R8\aVAU<+IU:-CKSUP-Z2,d?Y@9g/E:;cJI8F#R9??4c=DXCb4N.g723U##9A3W
1_A,P[1#70L(2AM-#[Ca;7T&S>7bT6\(442eIcA3SYCMD1Q=Ac<>Y)VcgMM?\BWU
DCQ]W?TC[<JU#1^eVS)\I\3gHGDCV,=7RU9(1GG^83PMS\5?[4YUb+5);6OIgK6E
:0\e+6T1S<>VT_3S&[E4S&d=)VISUd6(CM91TVBCI1R\H<<1<>Z6F.K\8O+CPGc5
8+Y)FCdTMRM@/bb;45CKF4K1fL]I&Q3gQ7Y&I]/:eX6H?_2VeX(8/GQ2]W>AcF&E
1XF=.f@g92P;cbO+\.U3S?NJ:EWCUa07)IRYU6]d2PBdOcVI>5].Z570GM<=R-Zg
<K/1#2;.363QR[NXK8-gLL7Y.>OWACD=T)3]8cK&0JW#M,0.BW[XBKI-_Y)\Hc(U
[^5HSZ^TKHV^\^O@aI=SHaI_/d9K&Q;C\/WO-T4E-TE<D-AG6GUFbPDY<3^_^/L3
RL3Fd[?eaJ=Z9RI#)IRV2K&&L0]C[>#K#JLgUcZVFDI1_91LbEN/^XeQ.5F;>1-#
DdaAX6>KS>ER;a2D=<[N]-ebKeCHWU_VRFND@NA;e[A#<[&G7+7NJ8CX1YF>JLBd
6dNH_KPAE+)]0Z-a<BAW)Gef[J,G9>P3M(1F.Yf8-6()EM[Gg>S<9-378+E9J(S.
aF0RB/PY?(b0T;Yc8D1&R#O(LN#X8ScQL)3Zf4]_)WZG^=\8Z65b9LLE.J=dC3NI
&7=(W<]L<f:YdK8,TS6KR5W9;J?Y=T<7Tc58PadC\eP8f^A-)YMB4+-JKSYU?83F
_DFWZgK:D_0EeK=Wa4GgXUS4>RL2ODb.>:3Ua5KK8IQfBXBPW;b9a)2fRYDHZXH_
aA(K.KdH63WI.aae@]H9Bg&b#=PQW\T91^044:YV4C7gfU/UMW)I>;DL]UeW;GY/
1V@(7d^Y<B5JN:E4OB_CX/fQ9=1RR<HZUF.#cI^-U54&1/8C)@&,HU2B7]FZ9Kg4
c<);NZLZ4;])0^6+f(D(0fKS2QX/O6LH;JAPC)-cYO_;>TP3F2X?,eFTW0)J.7H]
J0bQa8:^9)99+0:=7W8]]K_W7?1XFW\4T6bJ8SV7EKdRZX.aG\\@;K2b_9.<f^J/
aK()>@#1+0WeU[geQ@\<3]<CVe-RZc28@b453D@P9E>U-.&7]+d[cEc(][.NKbLK
Zg&8G5LJ<1Ud<FZ&Sc4E<>7H@D]H9@2Mg:HC3P_XS=U8-.W;(8P2;4S7OQM>fCgK
9RJSUOF:M<4NbAO/WLb2YH2g0K-VA5&,)UN>gF?T+_Y>;^MROL+<Q<\9BZdf<0:-
]PgKK?ZG9)SS1WX4#bIX7W8G&_>1bKVW4(c0dTD\&S_(^,+M2c^6,BH[5O>?JHN4
6341AEa7B[:D5R-MX/87D9.2NZLM1LN?f=1c7Z\1)g)c8/[cG(9F^YKPE)A4HAP1
M_,2)?NbMO92gLcUFZbOb_:R1g58CYIfEE(ESD831WTbJ11[aBYG42T@4X<JM/??
RW^-(;IAQ;,B=[&/1XAK14)-I&L.EV-P5N7,M<TS,>-:bT+c6CDY4C7:[IGcFX?<
A0U6d[6547+9MJB=4F2M5#6Z7)-X^/]_C:[Y74/O#\VY/E??<<9/5eXE)Oc4#L<9
dOf1G@bZc:WC>JD+b+_f#ODd4f0\Sf0bM/LVFeB&/b<IEDSM[KGOUP1NYSB^+;VG
^BN0]A1ceaaQ,#cL9JX6[?XAS2T.:&\J7C#8)\eY203,_E?8V&#U,)?EfbJaIK/M
/fL#9+DHE;,F&UCUCK=^4bbKNO0=a\17VG-)QgZW<VR1;WD/F#]E7G(Q(R33HKQE
B2O0BO3B;O?7FNF/03<f-:4V?R1N8[d(P[+Q7gG>+Y0D:0KE-BXL_;D.N2e2\NNC
R>6.1e5)IVZVJMFb_+3g3J]U+VS5U)NW(D\E+\2QUM]HR;^BW?V00>LaQQ]d6@V8
U=?E<aT.X_Z5\d?/WWAZa5\@(2<(F5g5b9G>ECC@^X_5+_NP);aG0H\&eKa?3Q6X
_81N<-2T56@Z5K_L]F5&(X?H:.+SKPJbQH5CZb&79AVZ^HGMcPN&NXIKPZE>gU=S
9TEId?O[Qa5>O:PXa:_]#d2aQFK\\:ICHZf51]F<P&ZXf&f]QO[Wg,FZ8:)J.M55
1Y7A&bUdaTPZDUJX(=E-9S&dQX51>ZO/9f7WFdbLd[LR8RYWUJ3CYA;GSGE_VO;U
cN5I8O2KbBTf+N#B&5BgDDc1PN7GQ;)[4JIKEV@eMe>@^&a4I(U#cB0&6UD\6dA[
YMD2S?UXS184Dc_54fgICRMEdV6S_4L[)\GJY#:^MKK9/>+1<GP)UOFD(,De?d-(
PA77GS>R1_g8eL@]0ZT9=<fV5.R&^>;?2X^gG7PWNA,cXZE(4Q)[A6#.Wc70P-,N
,H@W]=8#@6gD-,IcCZQ+;MK[NE.be[DF892&V2&QV:[6J8E3&=W=4XKg&+G/.?-D
ORYAdTB#^IZSdYI>5U5H_;B,f/Z)R@cAf//]JEIg5ZYAB82fSF8@bX@4)57e2[:B
W>#WgMQ4DD+27X7:N9><._)5PI@)3D?T@G+/2UE@&eNGNgVM;0@D-&bX^?d45:D.
TU\/?97<I5=ff2;d5L.)=C;6<[N08SgB@L#Z7EDDNV#8aFLV(eCP[cMB\HR=#LSS
,T\=6WT<?&5:<B/HRU2J1:b]I.GS3A3Cg<&+.K?]1@>6=Q;\GPBGX_^5A1@SEE36
X]U@.[(?]IA;_EdG.1C#8?MA]FZb))CWg)CC=Zc\bN[F/7c,RM;U,bK^<;5@K_HD
+(I&PB6<1;HTNR6b7?EI_4=@[M>AX-](X3+6J9)4f:\B/+5/aAPVg;&0;N&V-Lb#
^C(/8=@=PKLB9\a&JN]+B/U]@7^)7+OVLdOgeJ65X;dFOJI11Z14=T-UG(S,X.,T
^;S)d[[Z0aX.>c:9d1Y?d^L.cUE(e?0,=8O,fQ:Y+PJ2]<L7-#eJDXaT+/HgOXZg
UfM90E5PP\,Y=bCQg_8@8K345=ZG;S1QZ#CA8ZS#BF(2H/PcU?MLXTXLcWW18-7/
7DAR3WTKaWeDaUN]ZKdd>-8S-VMfLagcH2P7Y^O)@06T+YQE[g]76f@?@+>MPCAc
^@/;5D9M1NdPb-\)T.AZ5?_R?D^6#&A59YCC9-B^C[1NP6d3SI(^]]V93XU\/YYL
=NX-UXZR.3^b]&E]\,7C-.\HCNS/TFAaD>6CYY:<WP(P7GeVV7D.0+D3BD4J&V59
,YUZ#Z66I4AV/?d9WA50:9V[d-?YOY?;KY[6c9HD@)aKFP26GfU(OCY3X4@;=C)=
,.a@2(#:AB84#3g)9<0D\6VCf=I]/RO#PSUL96-Ia\dEKF^?a>aFQ3/+fKD?(U#U
@-SO4J;/B9&[MMGP[3SfI[,ORMX)3:NF8Xg-UB0AG;b/=)EOJE\;_d4>,H=))F.O
Q&)d202:9g:DX8eS3ONQ^CG2@bCEaEaPdHW(W.g,-KEd7O#_TdR4F\eB/=0C^2DD
S5>MR2XQA7QV,/]0c-+[YZ5BE/NYZB,H<1Ee5Sf=+RI&5G/XU=)C/0N2gea5WO.1
9=EZ2>^E,\)?@B0#7E2#Y2:H\18cfEC4S6@R;,5QX6T#21)87>DWd)_C_YW5/@18
FWZ6cQK8[X/=8>;M^AY04(f^40QBMb/1BQ_<W-eZ&b(C/5Q@Q=[e,D[AcBc?GV6L
L,5\@6Df7+P2FHVKC1S9M\WNSMA7Fe_F(bQL8Nb8V;^g#:f+,T2C;A]W.B&@D(/-
[<ZZD5A]&^FX1&.O:1(8H0\U>dT#BATaMQZ.A0I)2APOX;c;YgU+2<T2T2XPM?#C
KY(>aD^BG#/_f>Og69ZT68;84<#M(^Q;<\4>=8R4MD5XEF;U.H,89c^K8WPI6>1A
\MZWX(AL:U:X;4E,1U_Y>)NdeGDU[BBb-=O44/[LOIX(WGDY[_>_82gfPULRf\c8
6C5WKd70=BQD<\.eGY1d,A53JKb47b13O[8A-dHQ3K:4bIX@BTL\YfKN9Y1&b/^\
3TUVF(fV7&N47CVU+V\<F_TL,Z(a8N>ge)0U;.WY:_P87Qbee>-82[]#T>=dMXZZ
W8NdVYJ7\Z[DQS2/#ZfSVH+5SSULRd1X;26.\R\ZeB3eBS96?f@-fJg5;8YY>9&E
3MYIQ9L[c3:6GP[YTc2BD4[CRefT&b1>(CJbecJG;1b9^D=33GSWe#K@.:38CHgS
)WbcY]Pf(&&;>.,?BI?W[7QA7+^ca(4,EBReZ<FQPI.;#1L(@RDE=5aW731Z]2<,
2VEY;3>)W\cGX\eJLA>?=RE)cFWZ>&2CRDN,_edUA^e@3^835&R:AF8gFW5BZ5Nf
K6OP<9AS=TUZVU_=H9.93YHgGNF),X27e)HAK/+&H.0O:d?=GOB_[J0&COU/6#4,
6Yg^M?>W5cNFZRYe)40F(P0L9&40D@J:466bM,TLM:(58SATA??]5IMfIE/Yb8eL
0V/KB0BOQ3fHC?6-8X>6BRTC3XGUZNZ#0&7#1[(>WZdg+O6Zf45Z7a^gW38dR,.5
?I4GSL=C6g^K4HB?_UD0[3;-P0SQQUBE8Xb5__F81?5[[@A.4IKRFA8QOF016e?A
JCG.;FNXO+F&>21RZUeQP8dW]LUR/UED=cKX<@ZZ[WZ4BWM]ZFS2/@N[DfgKNH0C
<e>[U//G^GY/&^M:gCe.T(-I,D:59HTbbQ;M(CAWeVH/P?,dLB8LPT(MeH^b]Fa@
<ML2APJB97e:R[5RLP+:WcR8e7R58WK;D\O-1A=,K93V>7\=W\X20@:=+XaSMP87
dg/3W/9Vb8+#ZNb@gdM?)<ARQ#4ZY9A9:)&KYVeD7gg4/QKZG998L0PPGf@B)-55
Mg]LO/@G)W4X?LgE_H92&X-CWU7&1WWbFQ^_I)3#:S#&W4K()@9/75CEBN]>;T^[
Q[Xe@]&F6BMY+J[?=V(g38H-J8/X5/Ob@[Z[EIA-&gU<48UZDMVF[>SVVA.QC5dV
HFbE^;dH3(]+W-fQ^@g)D\A[I?A>(#C>61CA1a5G;.5N+4:2dRK_\A>Y1+B&IUcG
+WF\gc2(b07.MLO;5XD)SZ42YG0FcI;7@--?R+NSWR+Q?(@-b:aZe)7I??@;bRLa
4P654Zgg,dI+]WT\]g_)Td:L:U=d)6ScN([T6CO#R4f._J3Y\O/da-JW@^1d2-B&
b,H9H==JQ0:\7Vg6b4ISGK2G1-S[.<Q\]<=<C;RW)^YfW?\5a/X\GXd3;;F,LY,M
DU3=SU[f&,O,,cG]BVRPM;gdbD.2\11bKOZc-@BbdJ\c#V9^,GdG8S02D[2_/H)F
UH([]<1SLa1>2)LX^Sg8=PSf^YQ>.96@_._=)(@6gC_7LR;WUBg^_Mb[;D/?:@/\
^GDX[,<D)M7<^6[3PNC=.)W4bJ##H+Q@]&(H6J3O/?UO/?@KAfaM?LYR7,VRT56L
f8dNU52;A5FX5K33YEecL#.Q8MF5Q^dZL6LMd[,HWb;]b-gW(AR27O_D<@J32#+K
YE&F+gZ28+/(MG,NOQBQ+.EP]I43J?1(/J_X64PcC0R/+@+;8RcK+Fc-bMG,ASd/
P38;a.YHebR4#9NcH5=7bgE-KA(980-MQf6NG\YLZ_5KVF>E\@(325.@bS3aQe9E
AQSF_V0XK_L1P.&L35;gKU.83e2OL_@f95B#5UFgb6&)Kd7JN_c[SS,DGQ?@9c:>
^bE:F/MFZ;)UC+a84;Oc]]?):<NKSE;TS/_Lb852PG_1-dQaU>?Sa,AR4I_:gHJW
@_>@KeYCR7G7af[]@]BP7.?NgaAPAB5=dDUObJ7b:dURO#8fa]0c?9[(-(6<e+AH
WVIAQ^A;#PRFYf+QS)X_g-/7,U,d?3_#3R)]6^0GdV09EFOaa86#U>LWQ&<AR7.]
<TV==cNOKFAP]WWN/MSOL+47?JF-J(TRG5A6LE)g8?A4MdIW5E?FF:1>C&/a+ML8
7+7FV>6Y@>eEK:I.gSfeK^9a\PP1fG(AO?;M=b.^@A.3d0R^]45]D6LG#)KR<acQ
00Q#a>A)&,&XN\Y5J#O.PL/:2a-5I?GdGKXE+D?;P?Z-__X^^_M[VS[FRLfJf@WC
e:MOT+e3CQeUJ,,AX0M+S)#SR3L<FX67=0EO2HMZ+C80-9@3fZ1EKEZ.>)F-eK\1
<4H1V,HK/g?.TQ#L=?9^X.7H@PPHLS:5G44<ca[gXcVIJQeYSVZ52>NVVLIKS)FE
@0BE?BVXZ;)\B:E4KG++]&AQSKVXYYfIg&a[;YRa:c4:O_H=c@dUAbF9cQb_XCOM
,Xe4\,\#MJ^UQaU;CRE7=Z,3YdW77W:RR<464DE[9WWP;V//P::,YbP(#QWQNTKY
HXODeaO7D&D;UbW0Ld2b2PO-Og4C/;R)695WgE@/Y?]_9K=.+=b/OG9N[ZYO?@Ng
DH=(#L@)\9;S9,7&8;(QcYH](W,#YWK+WJ>>U.PHAeO]dO+^-AD\Y5X?bTf[9D@U
R;C1Z^]7^^PI&CY6J-Y8\fQ/YWX=Q/]0H2.ARE\KYH4U=N#24=_]Ab;W&-GLZQFd
b^TS(+(CQ.afgO4b.PT\d]]]/bK#?_AfM9=\TNYPV+[E2XJ+B<6NM8<W+/B#\M7#
V(;^fSfg8Y4(7HA.5bFG#=c?;8)G#dfEG[(Nb]fbM#>;LZWdS6&YN/X:f+<3,B:?
aZN]cWe5DC@S?31@HfEdMZVaZVdP2:Edeb9gP[7M;6@AfTS6EA,[aXX8eP3XV?aa
c&X>@ZJ6,E,_>0:BD1,;S@DZ\HOaHfB@J/Nd0dV[d5>[M,_P?Ud)Z7ge>5Db97K9
T:4T,?@>F,Ba^/-#B@GXDdA?T5\ULgV:ANT;NJ;K8fc3#WIDXgZMU.NSL?_4^\fA
=DWJ?^aM3:6))445@UTDN88525Ve7.Y]N30g+,\g=dC)/+&->]-H)C(171_XZ&/2
e0L30[@?)Z?G>8:cK&4]T^T]Rg,KA6-9=TE]HCaA/JWb-F>T,He1f+F\>(NGA</D
FcdJ.Ce@A3HI[K>9UH9@@)g3?8U+]\Z-/6=S(N:?g.03R&?:Pe94AV,+,_gfJT27
:0BRV8,Ud9^,XdKZE58B@c7M=\89f6.Bc;V\)\HRE&,5J;EQ7McR,-68T/8&_e[P
[5(:J6c;W2H-_+;e=546TORa/b9.-#^Z^#.@Sa1B)WV4MHJd]6RC::@J#e[QTcJ]
3f]M)A7J(R^1]ZMFPZNA:aE?IOXEMIH<VI,V-c:;OUV306cH(\WX>[6W+5>DF+U&
>(Lg^>-A>.K8]/.T1V,_AQ6bVZ11&dC65U9Lf#SJcF/J(ILg7We.S4P+]W+#)^FH
Y9,9M5f:P-L@:^AcaVg.8.=06P&L\9W]Y^15);X6G#8@5B9e<B>AGC,S-a0+ONWI
7_)EOU\SZBYWMe:^T>aPNW;cI>8Z5b44I<[9<c:Z_=RW=POeDc><8U&AX1/TV0I2
U_M,,KA>6NT+dZOI=_ER8bX@8FT8QA3g^-;K-[>TReM:R6N6S#FKEQ890(C)52AK
XZP>G&XDDSLg5N\=f@.5A@I-d+a/b:PdfO@&H1-[,T;]C:Bf,Ib40:(>-+;IFHA&
)eKFUD]a1-J[1)bLdV@8BWY6WeS)\_=^;O6X:_2MNA1?I7RL_eM?EU=+g<EY_a^e
eXV5HU.GDHA]SD0S5J34IbdX#Xb7]I4Y=2J7Q)(+SOc^a;:[bD^41a23B[b:-D[5
LTQDGB)f]VPa3&Kb\7WM=UD(DXRAJ[Tdg5bDUgP^N.GS7HVQTg>R]R,+/BHBa<6Q
VYTa@>Y(L\E7H\I@ASYULK/THCTTB:XFD<)\.ERTd@9M)7[a)fY[O.)e?60>f_A<
[ag67-^SSQO-7J9\-RDAb^fD>AADGfCD>T^d@d4_UO)Ya^1PJ0bUNb,C]3TK]#36
\D8C0:0B@K.I@IPQ82:b/WeN1&<<;GGFHE[<ON&:TWAF_[-BFbUAH2)GBDHBK)_-
<S6Y]D6cUgQb/8beX/.@&NDDcHTQaZG.\W+0;0XQd+/F]-_&TYZLQ/=<\Q=HA#eH
&6@(?[Gf48]/b/[-NCc(bFUDd1P]FJJ,Q)/?H-EZ;8=X9++=CSZ#S<^#4:aBD,LM
=Dg+,>JX4/1#\77f2)VX\P.;N8=;#9L<33=0f)TUJS+W;VO7.V@]a:]#QeM,8d:/
_6g=R.&GI72[bFHcPb;0fZg4EUY\(C>R8]fMcY2L.(_/eGA#W>PA_ADF)_GBA6G+
+>Dd7+)5b[Z5M3C0MCObfIgbJ<L([HFGbE=<]9AK0g=U;af#ecR^OY]^f9cJaCVg
A)21JdD9IJI3T90:43F32SM]D9O8U^Tb7^;KLX.f&,0-Lb_7/bH57L_50YHXB@@M
bOc(#\P_P[\+_Z.MS0Lc@+,8>O7Sf+>.=Gg0bLUfMIRP1XALf&LHNE52-Y\JdM]6
TP>dIbAY?1e@Ma8C,eaD>aCJC8(c8;JZ((=#[b.2&5VM\f(@=WU](a&R;NK>c2Of
MI_+P/FNN-YV0FWGTa+5/DZ->c<70,d]>=@\:(a)NJ?S=>V:\a5a)&7=a69CO&+a
Ia.0@?\9->g5F:C^+\/Z0]8X]f.0JM<)9.8F<,cN,b>@E1(aL_G+IZ<08\dD=dOO
#PCVBg)F\b2N/<7K^IYJZ@-(]Q7I:B@g9UQ.#;[Q,AC;^BD_L7O/-;[/WNY4a/H/
gfI]5Gf1+B\77:+B.9d6G/<@FOMEL;fA2.I8X6cbeCbNQ@:gZ@978;MefBE)97^a
f(cg36H:?G<,<8/@9^D?H8WM;>+X/1=2?<Kc6F0@IW]7Q[UJ2]@&N[I,d==6U5RL
OL=aUQQ@X(fc>I773YCXJ7a+QWD8E21Z[c,@#/#]#Sd>\0;]+R3e.e.f)//3c4)R
/,b:CY?#ZC-g]6)^cff1(Q7DE:Y^e8G];aK0DDBM??\#]YC8fM2#AgR4-6&SUJ^Y
g+WV_EbKaY<Yd02E7b+9Ff?=F<ZeOR;a9a:fFI3b8b<S;^IK)PCY.<([bC&<&P>;
&G@\KRZ4NZ2d--U1^,2Ja)1X1@HN;P3ZBXc-@G.2LLHG\;2A6ERE^)9Z,FM:1:B)
5RYC7VE_+VX;:(.BaggH_AU5e2K1KSYag@72\bcW/IbQO1H>2\g6D#JKa&+1>d/V
1eX>>Q9(f;W[+g)6fF]:d3g[B]?<JA)Q<KTF0DEB.0M=H9gg>N[@bC7>dPJC2:/5
7bLHIX^UI,)bY5YGeGWUU<3Y?NG_]31f<;Lc:,;3IJ1OXGWTN10@gI_UeHKJ)?Z0
1.ZSI0FW9]adG,HWa#9&S<L7DadHcT56bg8,OUG5bI<G^#Q^TTef@QN:7R2I_1OI
=J]#Uc\YNX-6FIa?Jf1RIPT(9A[eCOc2?+;FgRaJ&I3EV1eLSEd#AM<PdA,73-C+
RfQ#].&F3Qb9f]>.Q/DG6V:NUMV2AGP/J=W@&_H\ac2[/4B@gd_8e_[FLCe]02GJ
<Od4]UN3:&I7TH(]0_Ra\ZAN9<IUSDf:be7I^.X:\aR>[DW\@PZd?c92=Caa\A^,
)69]A2A]KG+d&&Ae<-Q1Xaba>)#OBa,FJ_44]@VB=3M4d544G+\0M^<:BSB_8#aZ
)RbIIeJE;H)(He9,P(QJB66P\)3/5<^=&]c/EKg:4ORCO5WW,TD;(G=6g5aa2Y)d
IJV(c5(=_dD-\/f/YY_2[R6J]7E-CHa20[M.1,KXHb_d2MIV?4AJ28T2\e@](QgK
d_>6U3429C@2[6?T.D-V??&?P^Z(QJ10@/H#TM[/6D]7.M:N_./=^JW3R.>b@3]?
<gHQ(WYdR(#5:fG#9(\c0V2+X<L.NAZaM1]?6K[&F&I[CNT/9SS][PITV\B1FWLA
e-4fKG=RQ>0342V9D2Tef&f#Y_J++VJU-Q7+Z0)>RWeYPA^F4Ld7?)EPV.13MeZf
b<>-.,W1?cH8Z3@[cO<(81a.CZ;Z^@d/]]#<RR_2/P(#[f[?0TcY0J\7\II>ND0V
4@L..a+#?-Q6..,AgD4U2A\JW-cUD//5L;QfI2(I-ES-U2Fa2U[R)@Q.>L&>G027
,,KL[L?#W;69dYWLTL?6=^a;--GF^e=UbGB=f],<R^?[TAWe)@c.JHON-I4<<]7N
VS#d&R.C\N[O?S]+5fCO\:=UFN5N=]M<SH16DO<_W6H\TX_W7,8YJGV6H6T-RdTg
<6:XY7T#d8-_-J./I(N:Q[+3T+1O8&d.KV;aBH\)C0eLX>SJL>g@(?g=Y;Rb<g>_
2L3G3^-B7+MUfPXQ;=+cRYf;@g;_N5])cb9=8c]7:^=Y0e-GQ\W^TId4&[IS>807
#:A)b]G<Y:=P?\=PL-ec_546EF0;3IIH-?UOYFORT8Q)_&0)Hc;;L;^Q&#f+TCe+
U6-/@MTaKFLbY/3QDL4g25D.N/\N)d+,0bH-@)[P=DN1S)TXPKXNU72>7HP4VMCL
]TI>/PI?EdD1[<2YOb5]WT63]b26GBPJISWT;85;/\UQD?CKb3Q(VE1<+V0[M6Cf
I0V3O@5fL[A_SVS62N+d\FC23PB)GV,b/9AEBQQ[+dEO:7)8g85cTPUYCf:gG=UN
]X-Te6QdUV:g+_R[TMH\X#01&1PX&H\e4YOA^.Q3.CH[egSSO(g[>0_2:4+d>W58
[IBV_@I,K=Yf&ME7NgDN:]Lb&a#TQ(UZ0e1V[e=0Y05^TOM8.N/6g7YY6F2J?,b0
]<LPYdM]g4A/e,B>cS7=(B/_9Q9=;Ca6J#Y:#,+7O8?-W<:[4.d&AgZPM[HCf1-0
3bM^N4[1(_<e>J6XF[5,1>gCbLZN[T+Re&T39UK:Q.a^CFJ?I[GCJg^Z^O^VC77R
[C&C.0]D]KWT6H(CJ1Xe^CM<fY7PT)E>B<J#X;C;R3QWN?,9IFH2g<d@^,=BVP>]
ZQYZ/86#:N73NHW</&RJNf<G,HG9?gIgBU]UC:@W;<6?R&1(P]ZKUT35^4FV=W@9
\1)9fbTeJJ?c0=]G;V\H??^dbbCIQ]VD]LWI/L#eTN&]\#^MURd4Q+=H:@/Y4Web
K_7a==>b#XJ)6PXJfc<XO(,C]d[C5PX\(-g0Fb2YJV:P]#&YPgJ@[XKf-8=<030#
e@7I._IgcQQMJeT30BR35C8)PMe:AZ2=+5VD.c9GQ[8;bZb>Q?5P+(#V.GDaSXeb
4JB=f-eBd6P05f9K#_Z[/Rf5;.:bGg9YUX#+Q+?9(C+,75L(d65^eV?UF^@SOeM2
a>@,O-NJ;cY.;E);;JC;aI;-e4Q#I8b:>[MdV;;R^.4Z-F-?=9a3;J)MSM&VF\(4
f<CSSHMdL?3eXfH9OL@E4g4dK&5UE/1Ef^=44P6+D9>YCGVU1=dU\.4;+3UL]:;U
Y=4EM]4IH/C-J0SO#fNQ4d?B+;K]MC+EFXYULC+3=c==a[53[+<:B75Vd1g<5A+Y
CKTA9:AVTV=H^>FK9)\U78>T;3GXZVde&L30B@HW,+:[<cd&RKW^ET5UIEK;/HO]
bgd@5SFG1VQb)8Ke-ROg2/FfOC.d&[,)=WDJDBOIeC5E)#/).)=7A]<\OU+>[I@Q
^-ZNOf[W=SZ=g1_Hb[37JMaRgKHQCAH.Q:C3027^GaPT_J(KCJ(bFdN0,.U34EM[
ISY[=_[#7V)N\C2P7+7O38c+&72&C0D^[eSD\a>(&b^\?DBPS>Zd50G>7AO>GdcO
X6^YIJ6,4C9CYQY/ER^C^V8#LBD7WV(J1<=88g]56\JMT:K7B35,ZMef8U#d@6Sc
/M-SQ[4(9HPN<WJ]gRJ9caU[[PAdG=@M]G064/WZ]53;c1KR9/C[E1KD.II\?V+9
\^G@6\4GEZPYDHOT4M&LFD=.0#O)S7>eVK@SFS:LO=/#>R=0d:1eUO9gZ1T8:#6N
QP2gVC?YgbR_\^bTS\K5YI3#:SZ[E_UDWJTIDUZ+6,S=Q7[.2C2[1S)94WAP\dT#
2cZU6X\2L1\N)YWA7baGfb<T4e3ALEP8#.Y)BG-5:Sg6-OBS[(6E-9>7\GX13B3@
bRbEOOH\43CI+;0eY33BH,8=BMBM5P::WI-+g6P5cf&I3QA1Z)M,JZHY?/-K+I4&
:N.dJC#D3HQA\F)VKY:=#Q)I[8<.YBI0c^YL+Bf+KH2Q)^_bMW8Y(?LRK<@Y6]HE
2]E8P+DR&N]GV,IOH@KdC-KI>VA;K+TXb9Z#_B=RA-fVJ\TRV\c4W>f61c_adE4K
Ic11MGg0>OTM&d)Lb2aURUMZd6.f(6@.0\>-CLS/>4fEQ/+=HGcJ<(5<8CI1;ESL
a:JAR0MP-LT=B^?VdUF2;9?;[=51[XL;f5_6UUEROH[b\,gNP^TY[I/&9GT4F^e1
H5MVOTIM-#9bV&Ne?8A6JWG0_)N?SZZYWCBI57-SI:77/M\.N=0BaIZ?MIR3QB@e
d?53UQ[V3;IJ.+,S_A-FaVT8_eG@5W)#DdAWSN8@F:ba^9^P]Z>FdeK(4O@ZL@QG
O/_MZ:NQ3VD&PIOVZ0&[<@010cT.<DGLc@cR#D(25ECb&6C+1]]>SL^,YaRJ5/4M
K/_^OLROUbMPJATF7T2eN?EMg:&]SS]U^[,5;>#3+1A:>Y8BC/^c?:KRYQK6f]c&
&?B0>bY(5,S.C.9^85C:?bO:;;gY236-Z[]NYJRdO74.U<KS?AOMV364AFQ9a&AZ
EGN4FU;-/RF5U2?WBgT:3J).cM-MaE9D(X;-/L[36A.(UO5.[8T_]#G@LOY.aW+;
e;43HCH9)<gW1Xe/,a^8C(d0NRY5F7O@@^]J2gNgUHC)gcYIZ218]7I9&()B[=BY
BQIOLXYJ@e2.S2:^LDO,\^6SJ8;+B<D.(,R&FE@K_NVHR4:U>++[]=-Rg#O<7,0K
MTO6cMT^LYN6.6Q&b[77Q^S\+C^,=5Z=05YF>AObW\&W\,<-Z.gaLZ5;1AS4bW6F
dV+R5OD9G[3_C]D(FHB1/5<#^I0:M1K/F\\K>Y+V]XcQY:3bH&4Hd;5Jf4FBI>D-
gNIV>T##,dG?A(fd;B+@4S_]4CIb?<2b:I6CU(I^6fNEXC:dD+MU-RHb4@Z81WNX
#9:aGV-X0]39d.1Ya#CY&bgSRSWX/[+O;WYfW8P^=5?FLHZE<UFFPQ=L\?0]_GcO
<?=9L3BJI0T1X>Qc_-<gW/HL:b]I?b&eF77:<3OAeP]9TbaW+06-[eJfJ[dH&#(f
]EgR+6\MM9<9PD?RI(-O>;SR4O.&9f/S.(0Y6S](T<AVe]>c2HP>?dEX2.8\E1M5
//2F]Z8;O&GI^?-0X4@Q/edAU+)3Pgd)2<1Y/2MN>1aT7J]DA;,g:b\:R-\FSYTH
P67#@.)8.P^>S,P6#4(d9_UH-GDW_a:VB03Vg)e,B@J+cXV1eB5(f#b4X>H#A9Q?
2F35(\?J;(M\->;[V+@J&\/4\f4]O)0?Bb(a-&M3RaT@V]1S>OdAcUBB>>P/\([?
CZPc8^/=Y;W,59Y:6&11P691NOF#,16QTV^RII0V&:+c)T;59;FHRHReAO+PC:L#
FQZ(\KYUR=:gK_HP7a,G@D\P\9>f7>d#WQ7+L7b?cMQafHP^#@?]g[P8=X4/U)9[
UWBBT;c6AL(W,VUa)JgY?&;/)3_\M.R]b^)3<GC8QU=AR0Z#K4+3/;UPFEZ?ICA#
77S-9Qa+C[H<K0B&C9T>A6P0A8H\dAS0-d&+a#X_TR+&I&T.^1Sf5ASdAL=6&F/L
MQLJ[3/3IXf)HKSZ:P]JAa<8=[4N42Z;NZ[;4(GL1SVRH=TLCLUeBDK^1cF29JK(
.XC@47\UA3SAQFQ3(+d_EKIaIA#bd]KZ-Q\W_82?d=E/];J@_MOe07a,@e2O9\&V
VX-_>?E1CJe3;U<UG@^0g_@0QK1&81^L&_X:dM_GRMKL@=.Oc7UFE3I+(AAI/TY,
8M/<=Z\8\c_,;0H:IQ^@?1NO8L#SfSXO8HO3S?4SW.b6g([E4BgMf3C)2BIMf5FN
IXE+L>f_MSO,JK+;eeY_8L(ME[.B1],KL/SH5TMPBZZ]JQWS=)R>&W:TKAL\5]<g
ACR1bb9S4D8fRXaDf9L/^WF9&)QXLYcYV#C7HMQS1V0:JNd5^N,<G0&fQcb^:>T0
\T46#ZE\9#QF&<Bg3F\44c09f6=g;Y)1WcQOe/A2;Oa;?dFA?.<G_B?E\dKeQaa^
F^]SC4X<NF2M.72CZV&DPXJSOF1B#50A6f;T]P?AX,D:3A:.ZA7_O[Q;c,/gUO^5
&c<0?+EMA[_>:62bg5W01Y;AXcKE[Z>76#EQ=IcJZ_<N,WLQ:7#JY([LQ2Y,FeKb
H1eSDGde1RS5DZRg[(Mba\e0BNV4?cdZ6-B=-H//1FI1gBdKV7^a\.X>37f>>U:I
(S:]V.T7:\,X4_&=81G8_8V1]H.:KZ[4N0W?eJA;[_b/=Mf;;8OOX:2b?TN<XJ?)
Pd[+GQFF8D:-^cP^>5]E65d?94U665^GWAgWN(FIS8.VPATH\8DX^CX0)V2X-7UJ
gGcT<I3eLace.^2VM@[:WYJL,8@Kf?NPb7]Ud175-J9YQ?U:D^8JgL>3<(H3LTM:
\QgcbPRX(+\=\_)<Q.460@b@B<^2,IO-R2TMO1IZC9^\QQ1#6-B@O7C^6:PfQ1Y#
Qb334g<<-WHI[<eLH3gL4LIULQ>>fX.ME>g_=N(>_f\#=(]S4(SN<L2/_?/:&&\W
Q7D&EOL0O9P[5?;HD>96IcP+N;7(fT0d?HdcMe//MUA-8SG2L1&6:#D3AAfc&,\>
HH^eDVU8<fNYTL2T._(2_eaT^e<\4DVA\YeH0\[MbfbAWC\Qe(W=510a_7I2SFD>
(VPSM]4dY_?HUQ^)ENSb\1C8:DY8)P^CF_>0#VL&/3^<_F7(Og#(^LZC#>/).QJ[
:d+]-;68-ZOcO.M7K:O]/?,\&Z\1I@</7g7.+e&TL._WeS]D5ZT\8FXU//OR/a#N
eWBP=G>fGXg7V+S9C8HcFGO-cI&_EDQd>HD91B)P6f_e,d\C(@SUfa=TB-FGf7Jg
SbVLCK>PS3IA-WGfF^F_(MRZ[82G+HCXD,.^+_NFW>F/C]-5K->4,61baLT?A0?^
P<2g4^#FJ1<\44c50^aT.+8\?20\98AH0dAGL;8:-@7Mf5aM#+dUe/-:Q7UA,DGC
HRH\J&(7VaLSTWH>FR>\R7A:c=8>HRH8>ACgB80:M/TKA,EXc:)H48B;@B+35GSA
Ya)g&<BT>RIJCC\D-51BMPaH<8^UW#gGdB#H>_O\<O&gZNB&>)/3I[5DZbT)M;/P
^N2,7@e,5<2V+;[->PA1C>S2OWY7.0f;D&9=0LL]6Vd-[+<<.SObJI4Wc8/H;8AL
VBN/HR0)Z[g(M4C8Q.E+JUd+GW2/5gFJ)[d.HFL?9^4K?/4,=9+]WD[.c3fb0#T]
_YD@6R^:C2ZH8A]T_5/V5gLT)eC/[0e/QA@#fR<47ab:;P859#7?GXC9X[5:7L<^
LQ96P.&P]/;0RN^[]?Je,,@LP^?BCVY(e5L)(&)FNeP#;:5Z1\]1Wdf]]e866J?1
_]d#Ig&535HBX+FDHbg\b7e9g#ZDGf3^[:9US9]B35[NMMH#W.f8O6\PGdI7>gLA
D2[JEdF2CLcCLdcK>?ZNaa\Dc-c(_8?eA.fQe\I_LTKB&cV1GB&X;Y=SGFKHT/R@
/14cZR\#XN,>^PF?/eJaUR98_N/@Q)U6,aa^.@7V/+=]XTDV.PVF/7[6KQP/BG@0
#8cED2R,cC0]12U:E@ZMQg\Z)O1^OU&S?K9[G=#252#MIXO1Gg^BV&HFL=[SeLB6
2bJ=02Q,f&E=SH7R85Q@cOY8Q/A+D[S&8,,02]#(OS,21V8]]Cb??[\)L^>>9U@a
d9@[;/.:cDQWV)M0VUdgUN7c-_Og]4THB2bQ]bHbU)bX_-L.L;/&CSFK?09J=5WG
3222Z)S05&^S(X_SVJ2I>+?d=,W?dQYe>J>9V-W/X;P.fOZd[UBA#OKbc^?UAMCN
=LM:CaBGSRFY[Y2a1.^Z,94-ef?_Q.58WagA=80:TgIRB0,O<3Kf\YJ/gZ#);2\>
SL\;P]8#DYMG57[fCX]\E&9;PS,(e#,DAT:bKF?c]d\@>S9\EgC;>C>5X5NA?f3\
.(^fWXMRfX4?V[DM2-#N,=\G2NKX39:0_^FPDM:0KUC=_GB3N[=S+7e-5EdRO9eg
NQ/f3BO[L&,8?KI0PZ-N_@8=.\?J\6Db[A+CKZ2?_FVLT2ZOc3W9,Of?&]LTN.eA
?R9,G\V6c,&gR3Q,?MgV75T(VO/CagQ8fJ)N[6+SMgN=V4-df9#]>.G-E\\Q;ecd
^P#Ta54)@#FMD>A@T7>LJB@5c__XBf_9_[I;gaS_R1D@2H/R[-:&^&d[bV:c\:-W
O5\.:Q3=,AEIKc:,_Oa&42<:@ZfD@D\a\f7WF#;9bWLL9Ff);7f;-^2EeJ)LIMc8
gb<L6Z#<3OGEffT<TCS3W6/</c4Q6@<b6^WFIaEXX3[Z0P6@D_TOXHR8&9OdBRW7
4Z[]De:1)33;R^:NS;\#6F9FEe[&</VSKX#ABTd_P;QH>=+#f;9d+N(7CZN+P38R
XI<S^ELN8/D1Z>;2RV;>O4a4SMDSY3.f7XbVM5+WeE+6?3XI<[J;_K-2aFfCb6B-
PISdFPJ1P)6dK;-+BcGIS,b6_MO2NK2YbO?>8H2Bf0eI)FI0&6a6<D#(]BQO3U+a
THI8]>GW2.O-)Q+g])EeYJKRBcP6HCVDY>58T:GKS7N&WQT2dMV_BLVF2219N):F
[>4dI]DCZ/XH1Q#UX09+?EF@&D@6F8Ye,&>Jf)ObAIODd.DJ58-5R=BLQI,?gfC]
MGQU063F>WVL+SXO,NOR+Z2a;)=1A<@a8)>)eDQ1O(,8_GN9E?)6&77gF0U<bX:&
:;NT[HTBOe?\)^,4&ZYc=eF:SMV,gOHHB(g0WZ=&e@S8\(TIHVZ,JT>09d;:;,.=
TgL^B_9]BfFD<UV<S\&c8Y5LJ72O0f5+02E5-,cXa&TfJ>YG6K-3IC;LgZB97P?_
fa9B:\MV27GdZ?2M^EXZ[-V2YfIg#.#(XFd1[MReaB)I0Ugf^bTgQ9LB<96-M6[T
-9W_;KR[G[AdC=XJQ\g,8E^1A?37HVgIgT;X5#X6-:0K51+7W5[G5WI;c.>ebgcA
+DfC=6Ode9(^=c>J+=(5J?FeLa^0DJ#eR)RFY;Nd(2R49_^b72ScSd93W9Ia?c&7
NB]d6[cYD&a+7U9?=XJ2b+C,XK?UL?f).fT?_GW@-3.XWFM-Hd>?3:bVYFI:[=E-
M-S&<A/bE&A4;8_0L^QOX&>AZR>4UPXgO<?1cOa+DgV[Z107:O.&J9@d&BJ1UD;K
[2VLT&-@V@DDAOKcBC>c:;^Z7A>..B-D_D#1ABDcY36SX>FV/A+SCCB;DE4d#6FW
5->PHMAPe/P+C&RO&0=gCgM)@C1KHDOIF6W+3J8f8=__8M87#D7bQ#Q(?KgPX)JX
R,?-a6GLbI97Y>Q:>G-WGGe(R(@OZbP&1ge+a8^CXO<7>.-^-<fJ7#bgH0(fD?M3
&5]c+I<,JK^.@QFb^I=ZO-;eg_gaX?S>3bg.)7@F5aC+b;#JN(T,G84fS5CPe;HD
V;K5S&bNTQ[NE<AVT?,:cR-)8BMYN3&8RU;f4+1.LZCeM54VC9^Ng/A-0]f,4\>N
1B#b72g9Wcda)_A5B87BVS=D)HPR_\9;;SH18G3eUbgWLZeR=;O,W+3R6NCS8&R4
P31NAG+IT1;\SAHRHN.b0eXfFEW11;YF]\CNM_N674+149ELCSQ]M([J4<0WH.C(
b7+6LGVSE1H0@)[AG^1dNZK=VXHV(CLUGf/H//cX=0BA3;)FW^D;5Hg)C=Vd;&->
>+)K?PX<?&(2U-5?WRND0F296Scg5Wc<aR++LRA32DQSYO\-_<Z-76Q^S0OSDQ<?
e19,)JL\M.f:D2c6@f&cYCLD+UOSWE:>g:T&gYGYY8dZ^?)IJA]X[8B#<9(ZYFgA
_^b8^?(DH-7fZ58=_bRAUM:0fP_NE,AD0@BY<JCMDN9Q5/[@TJQCc9OHb@VMPJE(
()d41W/X+&QdD^BM[L#JB#JbKA-F2UTE\EFNZ9@^>GPLWSEL@->S/8[=C.7HGF:W
7GXa=T@5.66YL;Re9e;_gSZAA<G&GFR/8ZV5;.^+E1]W1;HD(6OS1^EJ7H67fL;&
F2??O-<@K?M_+<2Q\YQ700Kg)U<]2.B;9BdH.2(d[,b8LZ5K9c#RcK80[6^O;(ad
7]HGSb3/,M3#^1_gR\2F;1.@JH8AFYV>7aXHYHBfNHY=1VYaC]PfKI_80)[QF^EN
TYZOC@30MeK75F@LU>?Y7VgQE?+4NQS95B&.@Kf9Q^>.Z5,ZcWdK2_ABQY-&T<M=
HQC0XS.#4e-JaA;YZ-/#R0;Ff2?MN?1^(d:Pcc:H+/^OS6=3N;P:(YRAZ_1M#YgQ
11QT9f2.V50,g[[Z]gOM<7QLY1V;G:\\/eNSX^P8563FYcN<(?HR>LCPH_E[5Z)=
H]Q-4AHNgLACNUa.1V+-Hb1@&7117dRRH=cQ7>9+WZ;H\]XE17A&e?GK5e&L6Ab;
[?H@7CVMd>Cg<]SKFLE\Wg997YUTW9V6Q7T<+/)>.3I5>a+YNg+=]RHV#A3X:GK;
aK2W6H(-WG038(V(55=,[J[K2,^GY>I_Ze6=-AGBP?4Z\?0]XQ[c.Y^J0+e@)-4B
PIF4L1U^e7\VI?gOAA&T9Wb+,=QUU02^@?a)CEUg((6:[-,KZN^J9HEfbCIHK(Y^
&N.Je5/Zfc6Q:@>?-1VXX#,X(P.Q4/g#A/H<\S9TA.X<4QC@_\GE,PWZWLc=\-58
+[.T=c6,IEHD6(Ed\cS?PSaQ4)98E])?=H.QNQ#\?gIPRgC1fL.bK?ZVHSA,fE&4
_#=[JYL_,T]WU&-I@MaZB,?PEWc2^(c0g_=3I=D<2>A?5g]QST7Z\c^?>-GXH:;(
b=F5KeL:AR6@aMe8@8XYL<RI\Q7^OQ:ZUG\/RP\W/R3E]b>JK=f2-@A?OfI3A^8_
b0.VRX[],D,XPOV/-?>>I/4)4Ed0?;CNc+&Pb5GFXfIB>KBfC=4GT5JDW:5W=5<0
YKTd0A;aT=\DQ[/dNS#d2)SgGA\S9)_?7R,UT48VL+Q[ZVTcDOP6)4(+.bED]IW_
8_(0CK4eAL+P;W7Y3R8[-QR+9#Y]X4+-25fTCSR=_)^?\7^aW&IX)W)1V8>(-EK#
(5AZHH6g,7D<UK\f45Cd[[#D5OFT=:G9,4&W(&R=;PQ\UFb^AD(ZBA6=^#e:I=)O
ER-C_gM#B8V+CfHIQ]=MUE4#9GA<b_@c7+Y;AeDT;VJ/#LI_UCX5ec:>Df2DSNQJ
KV;MB8D#JNA<:,/Z^==<N300JA&?K&B9\VV_=(H&VF&5IY6R=(_0\f/&EYDGUI8,
HJbT+]>d4f2Bb+<NVeKfY<HB+SC\-e4W/4?:/+7(<CUYFL[=U+5+JQ.H?U:AWE&9
G.Ucbfc2.Z@WKdS[>OFN8K?eKVH()-bCJ#-JP+WH_RPd#[b)=().g:B,g\fd2L4V
@d4(Vdb]->KI:e^\fZ3@6S9b;@FfN<BfWIWe9VJ7L2VH2T8VO8J/D@gDB);S/EHO
&E>\ZL43I-03[K<I[cag<FIAVI+KP8S1CdQR2b-.=03V&\((NT:7D,c8&WdE8_O[
XOP1EHRWLd.cH8dQ]362YXg[U=N7Wg8Z.Bf)L:OUYRMaK68H1D+HNCIC.&7GB4G0
ZZ-X-V.[=+eVU5cL9A@JcgB+Z)JKO[NL/^BP-Y6B[CC/JEMS=,[Ya6=8Q^>0VV#&
FT0A:-(Ca<[19/GN8Fd.WfbK>:L7EI/^>#7;FcL5O@0f7+Z)/#,=&\]-[HedgZ+c
8P>SN?,95INOL@Q-4<(]Y2P@?[A>WDUR.S)1)0THE>fKFCU-4IKB5BcLQX&c@&JV
-Q40-?I:IR5++H2XY)bg,N)HV<7X)fGKQS?G4QK^+^&L=g\dfPDcA]4c#)C,:&3^
dA]SM]4BZL-b5DYR88F0D9-&:YT3XSWRFL=[V/U0e\-WS>HVM24OZ6=>;Ld[#Rd1
,7:#-3BR^-5Ta+08BNH@^Jeca<G\bEd)2>Ve^7g@K24<S2b))bK9b5K(=).gc27f
4-ba=6>-HCT-J(GgTA097U&J_;Q-EWQ@5T)6(H-8LgMLA/g^9KPdG1GD&e_=332-
?M,HcILN6Gg[KC5-^YdT9;X-bKDCGTGG,f7&=NdBYbTA(\0_Y<]2O=UW#G49JIM[
@gADTL;6gdf8YeeF^)&C:8#/JH\96>aV[=(Jf=QO^O5]4@JY8KRYeN-N3>[^&9#7
dG5R1Qc6]bXG<>2C[XfEI_OOP/QXW2)-YE,^bcX@PcD[+[E1Ja7]673/[[5)O@eM
a?3X,<bfK<9FJST+4E&>74LJ(_d[\<fZLG2]5C0(aUSA;DbK7_QUVXOSeVL=UP7^
M9]f[^PDC^d=9(A/EJMDT7H;_If6eX]<<X.4CceK?4>F=#[eW.<@,Va[XI,<L02W
5#8R#D29a\D:&HPVCPR^BcdVNdZH5JVM4[LBRcUd/fa_;-+X6@I:E@f^DWYJVQUb
N5W9&W<AM#/3D:P:U(,<9<\D&bJNE2bJ\AW343;H+U\[+.&f]Pf.M>I;,G_0#Bg>
Q/EJ=BIe#T&A[CaXB7+(@d6dX?5=C3RG<>@d-_9PaG-5-a?.],R?SD?SC.9e\?SF
1c_;GJeeCW(:6d>PY9LTC^EWG<]G;7K6a+0)NQ6]/X?Q<0A#.B<QXC_CAf]]]A9V
fRSG;gT3dG1>LSC#ebA]\FJC@B&6C(D0?5[I&/5IC10LODg<;RCS2L).9QOdN)=I
g.K43U>J9B24UfKa3>INVeP)cAQQ>W-8B<SG7KAE>5,RVV5YM:d(@?]?)OQO]3S:
=LKMbJf9F-^7:\&>bY.]0QB/S:5fBb.T5HcOE,B[?S#Ja:-X0CR<>?N4(34,/fTB
OA[9:TaEV:ONYFR;W3I^-)L<J5\(8?O>[F]2D=_d5X(WV/;fcO@<L:I/NYV/LMdN
A0=2USNOacBFQ&3;+(R#&W<WE?g57:<^b_=UG9L(dcRf@6-T7R=FLC=[6Fa,1#7.
V-U1&<O^A)R#I4/:H#cDb.b.CZ>IbH-,AN0CY[I+3FMNEb^U?6M\;0ZY1BMBC1+S
=;:cP#gaX?PH4U8)a4)AMc4Ydc4R<&CH4e(BAg43_L=82P/G[1b8.cP/->#ZA+(d
/==Z-:)5Q,eVD#d;;?S\0QS2Q9=e;F9V/:gZ?Cg2ec^HK5(94-fON;Ja9+MX5<bH
f?A^S0,M<FHeMIO__eYc>PD.BXC=UDXYJ6F9?SPaTgA;Mg5?#BebG?QF>1L>DEFB
>N#OBbLDaCLKQZPCE)f)SFU;=DA6A/H3S.;E9A0JG&9@)H3dc@:@5Y?;9[#<.VMI
gQW4(5e^LPf=-9CHUcCZ?,2e3I:S?J@DCP_>\Z/K6:Ie[27GJ1O,Ec]@a[N;WH#A
ebXP6HW+8UDVDY:HIMCGTO0,82gaI^MH]\CgTTF/?#Kc+_5?GKBYe\X8\gEXJcPW
3\MR]4+U7C7@8=_F1?E69g#_)B<K[gJPa--fLD,,BfI#C,\KXK--SAHU1+@<eCJK
T]YVfG>.-UK:Nag@W-gMK<>MDPc[N@Y8ge>\X+Xa_H^9+?[(,N)EZ/K#:]8ag5=H
JWN5[e46PW13X>LC649)=b)O3,X08&.e9Kc4,>OVb[g2O,T18W7)WMPAO]WSG-H1
a#;eHWVd3[S;7c(:6+Q:A-E/5eNRR-80,L;OV.);^E.E>)4ZDI0b^B(aW078F+:E
-e&D_^EO1WQH9#+Y9EF0Ea+A<+dac:ZdA]C5@TO&IQ&)]ZP6_NEH;S,c)4=(6XE3
M-dST+2M#ULf?e,AXVS.e\JK-afc_4N3?9]Ig\I7GW9==ccUV:R);H9^@53;Ag]J
MF7@L,BPaf)]_#IBDYCL<O:4#SO4+ILUKfZf:a1\MN>FD&R:D80&&7[[B36@:?:[
gJS(0K]>RED7@d]+=c5;)^1GbY6Sd_c+.057SW5Ad?G/;9M>37V-[0Y&52S,3I1.
YbOCb7\&T]]PZ@6;Y^K4(UL>ZHCE6&e;LY#1R9&Eb)99W(HHb@c@O+CW6(If6HJb
fB5[Xad+edF;7+IUUBM+CHb\#\bWfG,.(@FGN_//TC\gRTE[24Q0;dM;YQOYH.<R
I]5e]])=&bSd;8NC5=#A@\G)3aE=DV9_UfB=N^R\P+]JRc]7_NbZ]&B_7I,BTX#e
c#A5e=eMW/Hg#.:SWOG2GY6>T#^d]FP:HN&6[^eb39E:cH>V2538(L>OZg+W]9=L
c]f2AVG8B_@/eA,)1fG1]/?>>&-3BbPK5DgeeCMA0ec-=G^8:K9caIO(YC+6WG33
@6E@J/D+M=D<A^Kg\5XGE\\JcTM2Y9aZ&4H^XgRC&84fHZ<(dJP-T@+DB_g,/^UR
F@?f3aGWU.&Pa\R5d].UN2W)H??dYAY_((XXANdVcG]F.<ae1J7.,B8UN544TJ/#
aDYK]&2>gHfID3XgUK.DdQ7LDJW14HX@CN+R7Z@a0PM5#B_:YG/02T5NY/1=&g[-
P/7=2Oc\-S?(WLQNRIB6+2Z9S^;G_Rg9,IA/W984SN?DV-70YgYAQ4]Gb[b/;XM)
VMK+XXS#R?(aOYBCa9a0@-KM#AU&g6\#V9H+QC@G(]dA#aAK->33e-N?EZXJ#4FO
QW5P#g0NDY,FQG;UQOP[#_=PPDGH4#^CBdW.^,)C^Yfd@A;7f(fED[.?5/DZ.12F
G\F)W]7L)46UK+X:V/:cTW6NFGe=I7,:(VJJ.Q>6@\I-1Sg:VDObOAdN/NM0B4-,
7g2:H]:GN9Q>XI)?]#>(8dLQE+LJNX?^,)4K:MIZdV)AHO7G1]@-7X?;;/c4eMJ>
abG?V?XDR?4#&?\Y=86WEY/DbK+?E#A-VDNe&@?1)S7?ZdQ25;GZ(S[#PFRb?]b-
].(>A_5CFY,N)>G=2A/VI?=JOZ.(WD@P1f-5:c9dVeATH1CQ>bFTIYB88NA?9UNd
OBCS,@9?c:)41g[&GBO==:LGDcY,@c:He/\\5;M8_f0[59XeB5HU<If&P+M-)T4R
e@5N@VeQ[T\3#O^=)<&eCaPb1-0U_)Qb[<R0gcFV/L0,e?QXC<cRHX@I9MWD.)GX
:,+7VU\6eCHSa)e@\GD=E.SKG;GcfcBM9K16,1Z@YH9R[-WP6Daf2Jg^AQJPK@<D
JY?3[9ZUJ70)E&+Y),SI.#E@8=;7)T>OFQB&V[Yg8+dMa<=<:ROWg]5\W9_ZMc9S
&.I74U02CL9/R&Wa@)<07+SP.Vd4M(XO9H&cIA8gPN1g-=P<]H97]]]&L6R4BFWa
BE^/c#]N^75JfE@;_I,+Z03BTK;I_)SJ1R/BBKGb&8W#@>_.)BR7:\ZS3:baL[c(
TgGJd4JNLRTD4g_B7c#^_HRa-)3bHg+eV)51^;?U_EP]fLeOGTD175ME/_<8b/[&
FOXg3CDY02+bJKUL-5T\3Q>C1R90Y6dAgLSO<A>8ZPIeMKJf0VG-B]=S^V:,2]d0
,L@V-:5Ja/2d?-b=Q[N>53TW?<E+S@((]X8aF=8<FUe0SP#B8dW,P#X^bc0.-.QA
S@506_3UQIdA;9IPU761;1XgC\FV2Z[2V(Z6@^@A05#(dC_P,Ge;J743UeIJ_M/T
UP0Zfa>#4FJ]DV:b_,gJbR],1Q38AbVC8HOG>-07/WF?\^5[&1P?XL)7WEMF)]Oe
(7M]=(-d(/)]K_\E0fVJ0bSR_9KYg_b(VFEM7X5<L3Z\T^4^BPUcB?P3DHGAGDaK
(,LB?-]OM)3Qg5]_cB]Q3)2X,C9Td@->@X(+#;K4f2<d;L.Ig]OFN->fU:,61498
ZdKM2061;U0c^EP7CbQS?ef&JT7aXAGZLSV\9dFbSa1WdBc-O6=U8=\[4@,=ge--
JGScY6Q;IU=/C@0PA6c);QSb]Hc;BCQC=Wd_R^Zb2IZJ+JgbVX3,X57<[U<6M74-
a.K/H[2U@,]_1HdZd6Q[S>E#gca\]YDHc\<I#Z3X@FfLL>=VEfM4AHL^->+cObK1
9.ZRY=7PX6cLG:0f/QZ]aB+5QKGEVV4R?O&\?R9g)L^9f:4DX<W,aZJ:T6Ogg8?9
S\&4#0>T/Pg.L/fAH2\#b6M9B.Md[L\=[_8H>&_3e8XU=KTQ+T[]aCP(C#d>?<_J
/.V/H617&Ab^OW,\Dd^_\/O]Q1YDeCa##OTMO)dd?[+Y25T7R/;30gHGb\8MAJOQ
>W(-G9VOcXDCbK((Qb:g(&Xd?c[;PL15cP#@GCCa3aIFTY=KG0UbR(FcJQ_][P;g
/]</=.7O4f7CINS\0NTH#D[:43BgZ&^NYSYdSa/KB)A&U]@:AARJ@B5K,=&#I@fZ
e)6#+U/g01Z0#=HKII@.J_6b&;D@XV8g4558#Wdd9gY0XFfVXcE+1Q_c/5XS(WT\
W.XKTd_C<69R8KGW[0_&,8VHEI=(X-@8Y2f1-,b\\HN3)IVB2V@T_)G3&Z-c>3dF
A#&;)Q=62?V1N3aW,DD<5^<A6MJ.7ST.(<4c.d;MLHTUc58];e6eB)fbP2.edBY[
VTT\YY6X\YBc[LO?D.f)#SR4@?7(T_^+N_Z0AMW<_BS<d5BNE+;+1HJLYKfLXHT9
>?5C0V]AWA9DeTdY8(E7:-V9^:Z.L4:9,BM<c].aZFZ\C:=+G,1Kd<E5I<#SKc->
f[GP;[F)HBeA5;M85/,J4G3Vg-&XgQ^P,T[DF[)./\CUQf^4Mc\d.(O]0.T-14Pa
:MY6IS?\L8P]GG8VHMS^^[9>g1&N[62^J_BEKF#9Q-/G5]E?U[f:gOGD9d:/>/[H
ETDU_&O-;-VZe8://V[3BTN](,WITF.VcSYMI8VG3^1[J?<^(Ga(.:&9,E;ccAW\
2V[0,F^c(AY\Z8:KB:dJ[=5;TERN9C(?0c<O^NTbP2@1R+FGQR\g[E/9YON^@gdD
W+7>d3+<BB4;DGa=:d:GYN\6b,#X\N)4<[AL_<LB.M.<3)=-9-03/aWRSe7\W[<M
[CESLS?4S0KaO+1a<fP+74S4^A1)KRN72\bQLOZ0.eIDSPIJcb;If(RD]ERZ.U,8
O+0&(12<\8R7^/>Gf9OG#HN1DCZ@fYZ<@KP(7NJZcbVP/#5Ib>9<.CaU/BOH/M[e
_57<ge]O=4L(KZDRGQgO,6([Y<c.KRBJ24ALNILR4cO;d-EQS+7O6@(<N)->HDg[
G#g_:^WZ]&a1W6)N:Y+L_OW98T+=XW0@:W-JWE(\&E3R<2M]4cXN]+G48<f2@)B/
G:HBR&e2[faZ6c2Fa/)<W47I@_K4GV&--9X.&L6Q)F>9>d[\fL^P9Td^?S0fAZT4
V=\>0dXNO[.+Q:HQ/aGc;N,g\.^Dg?NOf-3LD-G6N<RCeI49SA[P<&NZ:RH^R+&6
E)#bOg?4&\GM8E6X,]fU8S/OJW<NS.JTP=M:EABDFO1#?U6G)8O\4[6c]f;G,aEV
XLVR/_(1c^@L#RY[M6UFD?5@^Q85>W/b:&ASE<#(E[ORJ]=1+)F4]:7G#1D.O](]
PZFaIcJ8RJBXb]eRf92<&J:?KE>UR@dOQEWQ#QV]+Z)?8gDe4ZPgQ=T@VQ1LFYXA
cX[Le9ZYWeY.APJKU?AU156gWG,1Ce9\UE^VCT?U:^_X994NW;>b]);2?(R\6?TS
-d8acUBbR:.CbYVbHK1Wg6GEbPGL+B@d>Y<&YD<gKK7:&3]QZC<)^8QQ9H=EKS3D
ICX^V;2.[,F#XMQPTQf.28TH:4dcb28LeO>X4KBTJ1\e?FE6f2A^gd#9X2D3+E7P
Ag.MIB&?42BNJ4=g]UA6.3e+I[T:]P,L1b&Bg[E^\Z/HIIREQS&^fd&dGY=EIcN/
LG]WZT_;QDX=Y[K&]E-/TB_T9e#:#[3IY-8FD[f.#O6/3-.^:a3]R\B8S\dYJQ7f
Bbb8Y)7;BP,<&+_Q1;(?<8T2TK=,#+Y/b^M)+Ag1K+cG&,61W.C_DKZ7MZE_DIfO
)4LCNYCL934O16be(,6-&DR/@T1KfX=B8-Bc^9B;Q0^P4GIg5@&Z/._7=YOd2M^]
=-/CTZ9=Y4H46K++Ld-X+;8W2Y+aY;HE7f\fVW=\(C/0J[@P\3G)KWCL(gUC_:M1
ZQ-73B2ZDdV@^M>P?AdZe36#+MT,C4?e3PS1/<3UB&?bW1Y_(,.ECBU6OX9Y75\>
1gMQUXYa)O6)T67df:G,LeF>)25+IAI]_<HB-P.Z-MDe-=[Dg2;YQ.0\JYe(/3DM
DIAKRCVLO4eE(ZC(-6]XR[Bdd8<LB@</F^L)-?e#8PBV.d7S#W^bbOYULUc.EE1(
G_dc9#?fW@f_T72QDbfY2QbMOR/I(<:^N#[HDU5MEH5Aa(Z=P_S:W_L)([c@0J-T
M7A4M)d]9LBcf1e&g\R1P?=F@\U6X&)bRJ_@,K?HK0<QJ@:/I_G_-A4dB#=&B#1A
=@8f+O]LWRQ&/Eg,9S^16-]+Z5._.[.<aQPe3HG0F:S4F=)7fTI.DJ2a_Q]+B9UP
,f@WJ,4f/a:IZ-c9SEfd;ca-V6+6W1\JDWRE/BSde@#HE#:5feJVH=eC\b5d-E[;
3&6W.:ZX+]US4I=0@1<ggBSV^DRf;T((eOf9P,1GMM9;Y)bdZF)JSXZUUUM7/W+:
E4F&/Xf^X[)4\]fP=65(0&Z_.G,1>40WcWa19MIgN&(BG6KW]M5(48#0_\dG5=,P
;4Sf1A2cX\>g(eF^F.3HMDX<A:CN/b\<@9ARHM4_BYOXJ8I4SNV]W&e&GYa35,?1
(6+_GLQ;+^fR5B6g#c[f#ZAMeKUbT(.#WA1/52:V1[4EW#W(D(6:[KN9&U3:Ua:O
.AVa]CR]2MSNY^H/d;[0f-eLS+=N=Z@?S4DcZ;V<Q7W,)(OYb&.@AO7UN)R?UcDH
,#76Q\=]Q?7:bQ6N-fJ][RDO25bc.f3I4eZ)eL.:XV042_>b?UT&@2P_^[B00#-6
65L@G?P:I.VbESD?TO?4,1.L5>WQg>N9TMD[c?K95fNF=Og?RV\,X,:SPOA/.Je_
dR;\+2</b]d)[\\39M:[VX54?6,Z#RKVD\I31VeLDQgc8IFe?.0K+;:6UL<E^SB-
)W4=L14?5c=e_Q,d?>^DAG#4JX(&aYVZf^@3S@5d]G:TK,4FR;R^a+=QdXD43V<Z
.aO0Xg96UWbID^A)(=dN1VL:bb]Ba513?Vb<gPKa]G@[a?VUFD4V)@+:K_#4F8BL
,:Q2]2?Q\T#J7_ddEM;O,)PIH6b[\9O(@,60\A6/4XF;91)O4=Q)EN/L94+[PGB(
X43L.5#96OL:7B0JB8/XB\_@_@ca:U?S_R/-bF1,Z+?2MX7UedCC6]#RbN]]a3V>
;GX#Z\HH18(+Se3C+F;Q3]5Yd;^]2E2DX@:e2EaQ=RBTLb=c1G?E-OBV1_1.TH&-
T@V2U0I)4@O/>@L(f>+IU&9J7Q2.YU+0Ma=ODS#3K3WU[L+7M^KXEIO>UbYK=O[6
6(RP3+W9^^DCW?Z0)?S7Pb1.;+,Q,BE6F65C)Cd1=ETL_^OI;]LI[>ESWLX\P.K0
.(g2R(=>]3=Q]S1g[Se:HXMK9:E#3L0O8/KU0QR<-&;_>.0a_LKH)81\-fHJ:6,W
V/C(E[e>\R2?5<_0bGM1;:CXT+P\#0/QeS]+UGB61\ZGOM)MSePJ6<,4+;9+==3N
IU[d5bM4&.K:F(,G<P^.bHJg)::CE:EU.g^^X0f4J7@A/Ma[;U4Edc:[N>\G>3Z?
XAgYc.gBU/A#60E4]VO5a[5=_OdS:0.X0Bd0-Te26545[g5f8B@XEBP39\SBC7A(
J2V((.:-[JffZ;CGA;[?Hf8YEAY5]gS.,71\g-fH&3eI@-#@\GKNVAGBN9&241eN
-1GZJU<#^./0/ee@)3L3>XHbK;I&[#X9.V^\(/EXN@5gL/7VH<<e]2TP](CH-I(9
F4FXG;0GUQ)BOf^G+AZ^G;_\58IVO-ETOF&;<1.XW?,EM1gVYXM:JG1I7Kd9;EWG
gB3=TI[>@<]ESLDaX-3H&9H?M5dJX=DERA=39fU5C7_PgSOR;:)+1_Vaa[D@OP8K
&9eOKLNCIFVZ(^dVf^Ya,Cb_NV4E4./JCXJ2U?KR@5JBTGKUA)K.DM6>L?AdTOYd
-R9W9b5803#gW^eE<WVUbJAM?@71-(H0eV=HOECC3)fV:+2(fNC\gS@PR)dA(@)7
fL9]>5#&([edPXZb6d?,>,M8+Rf>^>X^dV5g=c+aOW:0MP^OfQ>bNFQ=86BH(3YB
.0U_G>#cQ^3C<B21[6=b<b1PT(2,Ib#Oa,8)<&-0(d+cV?X8+fdd\W);ZZ5-5JcQ
-@#AUB@Ag@=bNB_6dQN>1,,SDM;?EZ=PE<Fa-DQZ;3=]a>/eWU+-KS/-fFD2G[@G
\WZGE(a)aXg-cX((V^.NCAAY,aS\9BZ6VgF2[X<,aEISO;b#eJ[<A]A6XI9XMPX:
DEJZS&8d9MW?^1O.eY@+.g\54J.afFR=:PLSNLa)dZ/f,LbceHeJdLULZ333&dG)
IAgSBg?JBP#W\D49ga[RAe#Z9[[)[K9Sa1V\W=T;CGMI(aZ3/,@ce.M@1,QV-@=X
@VNEgMV3CG4>=5Cd#8-_7H(+ZgB]N_8,E4eddfH++VQQF@1fcSd+5NS-\OCPOJ8M
31:)ae=dM,2UegXY4<4ddH9-d5Z;BS98AFK)8PG2B#IY=d]10]NGEagZ&Q(NG,>R
F]33\ffBce^f,]REBJL2dGPPeGHNfT.\P-A\=0)Pca?=A^;G-=7WgPD#WOL#Ad/Y
A(Ig@EfW>TK@?GHc;d<C?Z(#AEWH8K>\77La[U/@J_1b8R>QVc+bVf/^98&@S;N_
JWe2-f@b0-cR.BZVJMHZFL+23M5K3DZ?b<\G,D)=>dgO^-?8ZC2KU4T#UX,AB6I(
6:G)=dHP3D2f3.&Y>1@\\3a^6UI637]1E+B<R5[@4/f_.Y1gEH4>3R</RS)+J8.R
^A9[/Q.04e8&W^W>Of7[>O1Ff/V)K3L_I3TY@&Ve0;\geP?.e=OaYX=2Q[&^NV+G
d)801)+Da.(8\?HPD=,?(^Fe:c_7.CHIZHa]83O.3+=I\g)g2eKO)C2Z):,?Y&Y[
EF]e30QDebMB-QbE#.P.eNQRJ.;4[/0I,-HKYA+QEXGD)0S]UDL1RG<9>[FY#>&O
Q8HYKE9H4L[,:fP@adF>(f(_R_>ETE<RJcPE(XHg;[bNQ._XeG[TLETBPMB3APe-
J;60f/YYHHU]eN6fR?=S;Q\)\/=/I38HI,d;e2[D?4b4(c06B;/M1fD(0_?6XR>)
]CB3XRE7QSN-=Va4:SW(3MTAUda:.D@,,&CcHIW_\&40<+5)3U/OD\\WcFKfU.27
&Q2Bg7GNQAB,OdgeB<gGDJ4)WK1L-903)Q<Q6CF?7:2HAB6+@<cCcAV)_#LCc=,[
?Q:PIb_[[T,OGK0,9UWB;^C_./,4PbINAX1aE>Nb5=-d8Oa2+dVgd7,VLc5J;\<H
af&LLgIHP,]O&R-)K-9Dd>PNB2WY;E45__[?96:g753;E0L/@RX_O53d&2.WYWR5
&CI3[@EILBgU:QLa[O456HK#JNKf3@#TTT-.CF9)NS0b(D3645Y/V\.g<@KL\7C4
\V@aCJ;Q,]eOf1U0NG/VO-,46N;E2FbA:g.F;?g&YD3?8)]2X1+7O:e48Te\F9CN
5,;=@RG-T:8=<NLM?,F8^/&ZF3(9TQXZ9;)B>&,OUF_)FF&IA3c@-Z#XKMR>S;J6
Q-C1MI0U.6Kc_(&U]@9e9^(+BQ7ffU__Q:^6UCRaKQ+WIT=b<F[0^LVY3N<Xd][W
8>9GWD2@YR(_B_J&W[&[,0CLQ^IASYTXKAc_S+QZR\eM6IcdH^V5V.WWGIK58)e_
B@1@7a-e>3\f9Q:P(LECK8G2e5=fS6&(38]6M>9aYTP0^5,&8F?>YcQIHc=U5U8M
3>a9B#;F0,+bAD&->HJ)69E?g4d\FgOc:d>15&_:(.-aR,&.HP#KCU(,6;]XNV5X
H,@dE06g(f)]a0ZBOM-,R@RZKA[1=3A7Y]cBQ&A#M5,c;HA1.8P69?.WY@UgAJdT
G4]8PPKP_0U&1I;@e.QF/>FF7C6F;FfDJG?4@ZRZI8@9ZZY#eQbd2^fZ-Z18M4RW
Y57PH5Z;>GA-(XM=6?N=?<-9]7b[9CFX.eB)EP5[C>B[>9/LeMX3d^4WYGFc)<#_
bafZX_)^2N8V/TDOZWgXLXIIe\\f4G6ZVZ)[PM=C5KN-+Z2F..TOAH1/9I^7^+O9
TC6]d#XeU3aF+c3]&<OV36;V6+12d=YHe9^5<e18I4ORH>9;Wf]4T^6F@ZfAP.eF
R@;D?FB;M#I8K16WX]&JBWI;,+Bd]1@MRBKN37c<,00AQSbIP[eL13H/=7MAZX(A
F7eb?Ec.;H@R/O..U]J2MK;#<TVR7.F7=6HV0XUO#a-92.3=VgP[f]@5NE[\34(b
5CJ1L7c=4B\f?eEV1feUd@PgI6&)50QU)9KERU]=\O/0[Ib)EfSPM3/d\RAH^:FA
d]7PI^ROc+9<IAW1&)J3.IK9E6aWKVK7?3[/UF[N7(>ENcRN]IXfHgYS8?=ZSe_M
GB4Ge#AfIV+fSH3E7H(^fU9;7T8fa^<?V_aL..30V]+NY4?[T6-4XKA:Vdg,Z#O2
</adc>D(Z]-RcEA/Q/Y#H]_OaU&6Q]@D.2E4MN?;\9#6YbQ::50]cHS1(:>2bJ:1
=?Y?6=4ER5V3IO3JVX4;f<e/LCSN<aP4E_d<FB;eTO\a(Kc?8F)QN=Me0(:4^Mfd
>ddU[YY]4,]/3febXC(L[5Ze?J-X^RB)F9.ZJ;cHY=)F]D71KYFg2OR?1TC5c82B
D6@8K?1X6O6=)PcM&K&FG?c96c]BQM4AHMfHVU2cVG4<W-fJJV;:X?gCXOZDWPBG
I&?9M?,IZ#4gYO@FAGe#1?Cgg/D]^OZe+<L4HZ33</4/A^EMU&)J[Q?^.T247ML8
MW+G5&KTdbOb3N2#B+?&.9^,WC^?J2)c[UL)-YEQ_NRb5E(2_=.dec2d4_KPa?2:
?IW7Gga_KS#4WSL1F9AN[4HQc84A9Ab+J,3,Y/2/:#3RDG&FLg>UOAL5CD=6(6UI
:aGaH+cRa-,Cd@OgGR3HFf&@E:GPOc9b2JY7@La<FOG]1/>4-E2f86EDQHbEZP=0
SJUYK03_-8KS9ca&POVd0XUH6[b<V\\.AX,5.BO?<3SVX;#5E<RBTT3g4K_W&#2?
9OcDBgJ.YcLYA2YL96NF_1/0@SGILcd9??.T+I6:dA2QFCdcK5BMD_[^N)SRfWe,
T1HaZ>g>3F1.HG&D6=ID8I-^>ZAE/bS5PbL?E:X3FgX8_@1B>&D[U67g)S@NH[O>
=>a/HRG=/_>WI0DPV63[.JU=1LX1A#^#;5XZO50G9;;P1W9BYZYGe?SbV^Ed(Yc-
b@.G::U=1N(7cKNE(^R/6A6NQ<34fMW\)N)RDb@))EgQeC,/f4P8a42e_0Q0>T\c
8A[TH1Q/.TE-@B,4TY7:MV=QY;O.NDf@[=cF=e6e8EY8K1+9PIaN<S7\V3Zg75A;
XT9::XA9-,FIY,&8./0VH+,ORe;C1b7)07S2X&KE<b[<G]WW>6QLb>c]]/<I+fOa
d3a?cUX\>dJ)aRcX)aBL?]==IKL/WNU3.BXc8#_97&(QK4=]MY(JL_KU[Y1SdEYQ
G-9GYA-cR,]FK21)H-fN,0F1;928UB:c4b&/J4JcU,T+-Pf13=8GA[B#?DGL\7E;
(J>J+0a.gB.9,4a?[8g0<7D,cY2aMf8\/RebKbW]Y#aB:Z@CW#WA\LA5TQHG=\:b
K+&W)4&c[P2=/@Xg#d^MYGP&J//8Ua7adS-[26@b_Y#>eJCZ^2&UJTU0X;?\G)La
EJ=5M-IK81@a0dD(XdG7#-D)[,>6cP8TE+BAH59eTC@c/VdTG;<fJF,._;RgcMFC
cU8=;f65(9P,f><D#e_6C:434WM^5CB8FQ6,D)dP;3H##@7=\:cV(\gKAND5CS83
AX-LfYQBY94b@O2F\Q]WT>2\])9BC6PCgHF_7BeA,OBJY(XbA0#_bVV&A;?30D;,
N<QZ7?<=Hb231I(R8ZV[2YCb9g(]])1,?XMTRa=6Cf-F2f_9_\KN:W/1[=EJ\:;Z
,H,V@/eBT,:@S=L<.BINb11;7b+8ac7.-.(=TK=MI2W+D:L2:D+TVQ4<TVE@2Z:0
9W\eU?7a-dO<#<Wc;]>?Q._4\a]aJ2A7YBZdH#TJ#TPc(E@;Fe=7.Ic:#Z4e\)=;
-N4P:M37/N],7BI>/eUQ_<2e9Y:#=D+LNIV_QFUQ2XJTVAAeDcb)U1(Fb-b3XV:;
L@g<K5)U2ZU0H[a,8bKB((PW]>Kgfb6Z:U2S.G-H@SUe,G_J&5+fW1OFOMY<e6IF
gGBgVX=,(55.7D)_8/d3Da;3eb47_O#,K@#?5TJ(O:GB[T)b?D-Va,B(&6]\beR\
#1VYaDbc9&@<a-(2GT-J5J_EH.BW8#]6AAHYKO1D_#eDHRQ[S@5a0#3+3R-8D1L@
3aVO:2d_Xf8(>?cT@?UV<T\ARUa3XKO.)6-;]2#d7K&4>+KXg82=Zg>1:SXMS_<,
fOCSD8bUbd4UWCO=5+86BW([@BF@Wd^8Z]YdX_9b3M-EFdE0E0T&=7APFc8K]5?g
8GJZe\>75RNTC-MH^c647,c)H_MK/JIY,HKO\M;e-(Q\7G2Sb,O5@\ZIaYA2R?aU
F+<3:V@P>>eIJQ^cKN0TSf/K4f5AD<)QAH=Pc&__b9NR9YZ[bbNa&?,MW@b<KS5C
JY&J&?.^<3b=WGV@K(dFc,e_G2Tc)/1=a,6AHe-X_FdCdc@(d=P?(J+Q.fI3#Jb4
MAaS-,?HF,839+P)XQ?:;:LD6b1]#37>Z:c(eCE,d4bL1/6HLXN(,FGef+.8FeGU
a=O,UH]-WWM_BTDf?W3(QfN#C5AAD/R+(\HWB,9ALM)\,S@FQU@HY0POaDPgM>_+
aRSd832b3KCV+,JG;d0@2?&I96?@-QP(BA94VP<3HP^;-+#-(aLa2(Da]:M#ge\Y
\=:Y_eVM9(=0+]+@Y;L<_-e.eRFf&YD<3B67<U(FK2e(QC.BGY9V+LdL_1Sd@/42
3(OTfbHGGV5Pf(H3>ef[PfO.+LeEJB\65dH;#gG3geSVDAH1\4_\Cd0V?e8U:W)G
7eTMfPDbY519F@2+,R)Sf3YG3;=T[6_G50Q4P75;9[8ZHMZFYc+3YRd56I_YdKMZ
/aK#:1edI>dXUQ5O96>:QPC5>&[,?R((?.DPDS3GGXW1QY^5(4<Td46IFA^Z,_@K
Q<+Q0==+9FH1gfb60@4d91:c?\(82V;QUFHAH>2DO51F7=b;XH?,J7+>9AMW6N3c
=((=6SUSQCd=?FNQX2^D:dJf,agf#M/PPAF+Qf2;X8_QCfcgFDaFZ0<g^EP:-ZJ;
/cSN)cOLI#;Z;-08&gP-&>VELb\[RbSQM\cNObV<L=8WbB5GLN][1)f7BFSJZf-2
7VIEbef)=@_:.eB,I]22_S?OL;/VF\=5\-EMH?.g&ENE0J877[;-He+De7T\H.D9
KOI_J)/.0UaA6H5@Z@.KZ(+cY]BOI@b5#8d,NA<^>JA=-7S,VdH)3;)SM]g+29HU
YD-dT^Ae:F47HNM(HG[(O[_b4#UTT?^bXR90XRT##T&]9Pb#G><=+bG9/:?_d8cO
JZH46ZPg;(N25R)V:@H<E9[0+]LLDL;T^\60fM.,WZA24\UcJ)13eQ_<CaU4B7B=
S>gR2-&ZHa.RN4O:LgHFA-_)P2c@]BMS[791e&A,SU@?J&#WUFL,c;;cM5=SJ.8P
55;Ja?@4;T^d<CP6aVB5e8e5#(X^S\)R:-?Ld-5W@[5KdC)0^<,B,e5-TPC_X(U)
T/\WZ?-0,Q@f#G85d+5cY:McA(0^bM\P6^;T92Hd_1#LE8:DZ]5=7f[.\4N>Zcg\
g-I+RN112G2EWfb2S;fPXZVF?KT.R^bB5<1[3_,)]OX+ILcB:gRQM[XeBOPRT-LK
C0IX@eEDJQZVW?g8>]7E5UGE;egH2DaQV?>;ag.V_#g-fGe?D>>0<=KHV(Z&LJ>:
/RQ:#DVV#FJU?>K0HdEN;5-7[U9<dNfg^,_S0R&.f1H&M;@DRe[L>T_SaG0=SC<K
XSdSW?,-0)c:.+PX2//#I1D#;-8&HWI@4TJ[EbJ&=L6QPB=KVWBVf0;RCQT1PJQ<
a;,Nb4V_5d\DJ#&bbW]HJ4+-@8Z6Y:^)gV7/([7.Cg#9[TdW4=JQZ]DYfX]J;fT,
WMd]B0dLPb2E(WgKceN0g>9/@OUD;.)@Q+.:QWA;gVOI6_K<L<<+42cAC^-/YVUD
d1A<\OUI8(S26;4#5(M(7CUWYQ8#He\Cg0XM69LR)+.D,PeARQP2/4TV7^HABZ?<
Z3-BBW0(<\Y(6IR@.UB;d;8Z>ROd\/;QBGSBIM<a<EA/0Peg4HO-fYP<<J)V)<=;
JE@;,251LLfI:CIaN2FC#SXQ^_F4,9=/G,Z<>=P5fE7cBM0K)O-H#RUc]AMK@7(K
N=K5-\(5&_TJ+[&C/Q16O.V??#,eJAg4TN(_.8M)c^@:OWG-G?]6CB+[HXeA6&6#
T,Z[d5ad]fO_4/X20Y(/fC7Re:7XX&(1aWR3K]_8C.(<^R(]KL\0ZT@E,JUO0\Gc
M=2&CIG]_PJbRE<3/bacCT@ETMGa@gD7F7C&=HSKbI0_:5(\FXP;::U+bW?TZ^<Z
5@JCe(ZKT09H10<@4)7>/gfL:C6)OfRO1.PP5:Od1@fX]TQ1K;-,Q>&aXdS9;:b+
J#[KcD22+K[7K#Z>6K)5V_JLB37@>aG0_?@+Y@]D_>,Q2Td62LYWKUdX,).[SVJB
KQ^#g@#b=&67Q@4D>WfFJUge2C>M3J_d3(A/Wb>,OS<1^#4d\OFNNE#QT5)\6aGX
-X0S6)5>c7-9?+[9UOH38^):5OK,5d78QKb+CX2ZFH@6EDLIZZgaACb+aX@4b(U@
[5ILDJ+P)I8Uf0/+?H_++0HaBM0(?_D3V3/#J<Kf.O8Q&^.J\[1,-G_ac36KHWB5
/2g/6.gQ.J/IX8<MF+ILAH3\L]3&Vcf-(C/Db+U2B(1CR<d:gaVM=E>QfcEQ5&?R
&)64]TLbVDc+#J0H6DE)O<Q>S:eIJ;,)Y++^a7WgS,;YTdK2a].0S2a//[Ld06^P
cDY9EUf)H7=+b6P6Q\IMVF/PB/P@-EWM/DceB+8.eEOC+@30O&(fO4?B8)S;Z]2A
A(d>M:0<OJ?E9,/4b)ME(c<6?Xg\X)3RF0^-EMMZT[D<T(N3Wb7K+eaHJK4BJ5Q8
TS[=Mf;1IY]):GRB#29PU@]7SdXNX3T[L;9>Q;4\ZcAHaeSM]T;,5aVTe&a+#2XF
)97Rf<P8OYd-(Ze=[^F#YH,V#1dF1)J)5Na0,U/@N=PV\Pf+T(=Y]66AL@6THD-(
(#2KU2ME.>Qc&,AO1cA@B[f6GgR8R1B_7]0Mb3Rb4c<N5?4O^YO<]3@6WdG2;M)0
,I6gf(_.e)G9WBA)EDd/Y(5E>PTM+1e^B?.V&.IJ#FTJ+]#W=H8#T:#6/93c5LIW
\^g5;V#BM+5bKcB]P&aUX^J]X0L+]F<?+O^23M?IQ\TU+R6U=N_[^4M6F1e^0V>:
G6LF]3L?HDPN0d6<(;\\?GgQFQ;+X\/@g@IC)RXGaFP@+ZF^X:eTV,6?M<3N1>4,
#>c[\(X:,3MMEF125_M5,b-e=&_M]B7)HbC^62S/dJ=-(BdcJ0MY3VT#ZCI?-]3V
bRZ\QAC+gM9FG9.d^TbS=R+gP]=g#,G60?6BF5=UJbY4<7(=P]-6(bJW,_?UEZ^5
FY)\MS1H+e+(4\T0@egTdfacFI4dA,3[UaC,25UOPV87F/ON2/D#\9X_)[=J<\Wg
GHCXg<93aW)6TF9<D;fA[G:FVgVRbd0d+41(eN12H@I+@)U;ZY5UWd75Xe0E/&?L
IU0\9JBTTf^d2.[HGYI(?#K).D</QAgf\a70LTS:2PZ8X6E+45_M1]e.7]@ERfg5
0SPOWg9I9ZPQD<<4:dLUOdRAf3@/#Bea,;1;[7A6ZEK99c22K9E<A2Cgfge=9e5Z
/CJ5GTbJS?9=2P1).WDXg(@KL<aGVg5F;TO)T_DFc@a8(0PY9TD:B@cX.LT;?C4W
&fF-U44fT]7cWa4?,<VOLe158F^[7]3_T0eA?a]^NMW[21XIc?fMfW5K7AL0YIE-
C&.ZT4K6RC&>YH(A?eE(U=V3ZDW@C@gT25SZAB4J#3?<,:;2VAFWVO9PGSRJ(8HE
(\MeQZ@ZTTZdUY/\VaM)_WDNg5JI3V5YB:&g^^cBg@JI1BKcE25)NIdM#(^3A[g1
@g@C-CP6gg[b+[Uc\07-2=_NCET,NXLE[SQcPFU(I72e-9GNd+I//L5/M,NFD:YQ
NTL#fECg\fVVN_Y+>1BDg#?0G,e](B,#>_,>=#X_a;6;N1&>c(Q+@a&>d4<LCOEg
P<:D05W)L#g^4IJRWgP@Y41J:cEC@aR4IMBUT]L=3L.e-7A@,T,CC51MaFJ,@]:@
;fUg5,^;KM;^a3Z\Ec0C.OC]Z-0]_&ZH])C\U-(gW)Bc+:Ta)5DeWEWc6effV^^.
(8[+)[9NT&dL_0S#XLd4DdJaBCEZ-OUB</XeNTUB;c,+]_)7ZH:U9\HB(05OPc8e
OADGKP=A:FX?2Q:-,Q>(fbY_gOAgRUMdgOI>D7fO#JZ_?.f&G4:(O))2(]6I+f4C
84-ecQN]7Cg+U8&)]@4?#B0EYd>80QQIZOQg<W&6Y59)ORQ/63KX]?B+V?]^1JOI
fAKT1]S+AT,8T#[4bDLL+3/+,SAHgQZ<6@QHePeBD_5dVWD=M>8.dcH-NdM/Q]E:
@5:-[I3C)#O5.J1Q_IY(5Ge<353Ag<gf(8=7@V))8)b88.>N5K1()GWWVVOEL7A&
/EWQ/B_TB7(><2)7C9((KCRN30e+0CB8OQ/;^[)AfN&)aNG<[V/>&[_+85^@\9&N
Ded_VTZD;;BMBZ7^C?O9@/[cXc-VffeHdM=b7@Z2U5AUf>G(.CFG.UDdOETA5U9K
Ne8]B:E.55FC5H5+J/:PaJf]R\GT3+FY>ICd-9GOW-GU_9V\6b4GQ4RMSHGU5ZfP
&T_f1Rb45:-f(O/f05AA2L/gP6/XB\YPJEU,?NaY-5#a+-4Z&INcBXfK^9N0b?-2
/50+fOT9JS)(BQf84L=U(3K<Mc->#:4C2YdB<XZ]d/1<RSJ>NXG,?G=dL66T.J51
>Ld.gS>(X5F.9LIc70?)@RKO8+bXE1UY)Nd48#=--_6)2:O.X(?@0HF3^Z:D.?AF
2(LAV[YG&f(:(1#A?LVU@/=K3?a/-_<P(SL<_DU31aMHVWUX45Y)>fc)R0J_H9YK
BK<Mec6O8T1OLcC[#,6I:c4(AJO/I?cWVf?M615LOPbM<8fOgAO3(5d(W>aaKbKa
Be+aTB^28VDD/fR_^Eb-N]#b-^.;<Q^O;@9FI=PNK&H56KaP9T\5<GB23fZXJZ,#
K:1ZC1A_M_-5Y4WA^_d_G@8[_)I2b<QKg]@A]3#HePdE+K&g@W\e?HUWP;c=VQ9g
F33-ZD;@[8EeG:ZZcYAMaXZBaGG,T;?X(/(LQLLD<Z\U)OJE]=M50EP?+I7S5V/O
bPNUH)>7eZJ7&&Y[))HVO8^9+OdQ[,#K:SM;_R21dP/3WLC6,-^FWZU0-&)\9X..
BXU0a/CZVR]UABE_88\+[&:fO>aeBTN=H@C#.;DW/R-:_#<cITYBIK_F,/gZUVW8
8L[A-J:NbF5Za->(+7+[dAS;FV8AJ+F:9aG[O\F)/QDZ1[YaMbC-(OJ_E@@T2feb
2^5G\U;ZVYW#cb=MLGC1N+FU=UDdfJ(]cH?NcR.0()NTHT&5N28OX>Xcge<-cIO7
;WZ0TI@CDT#0YEfX+,XR</A-K7ZW&01dMI46OJ3:GZ\K:CC>0NRP?aRNaQ(TIPb7
)?](4^3VMR?K4&B<6->&c]M@W_7Da58W0?B8S&:3aE=>^?Z:P8H.R5g-RJNF1O3X
bG^,a<N:P,A7a-]:#0@Y_\af#EQ5]RcQ/I+cVd7Z#1a&:fc9RDRBQPd.;;TM]FP2
0+U>JM&:;F-];U92B>7#9.V95b@6(-0PeJ_QB.67#<9=PFc6PV8=aT34g/[2=[5<
]be2XCD:FY2YAe.NR3GfI<+B_aSM,MQYGZ+^gg>,XFDWQ,E@63B[CegYB7Fb3YKc
a&V/0cP7TGFa@L+;#AH_fMYCC:NZS1dbc^V5^#cI&2]:_>?4M;96,A1Z)8.KJ0R^
<0LP[Q+MI.=BGBK7f=:XJE3;5QdaM_;;.C]2)0ZH&FTJ4>Z>QQF4Ja3.]bX)#7]U
g^\XA<&gP6U_AH\ZANMSXffMX09-_N&GQ8[&YXZ&5NOVWcW&#dg#I:3:c#&<JQ&,
J)U9S7P>9U5NG@b:DVFEeX^]YHF7\/KUeY[UG9@\S0SV2<8/BQ<]fd5J\CQ_]3KH
(d:OT@P4T8.dR+c\g:\QUKJ+4O[#df\>[RX+@D57(1gdgVCA^KgE[e61G9GaeAcf
Fe42dcbf57aCO3WGZeFd:4,-:->b=PR>),9YRRV,1,EXFO2?9a+YM[63.ZeeRLYW
3DZOYdTaG1ZD;B.:V:>?;3&Z;/\^>#6(&;C4;AddDa##5F(JHH.#dO_AA:5P,8;2
@^cVe6-<B0NS4NCNA,#1LSY]OU_GdVBVY#eJ_M3E<,2M7,dO1T/>VLGP57gI)DZc
PB=>DTBXCX7&3X:QM[.O)3;\-:7aeF7a)L)\E1_=9f9V--VdZIdDcB+CR45OKg>@
32a)PJF]<NaKM\aKb.T5Z^IDW#;0GDXJ(B6_O:Z?FZ&N]9X?7J,;/2(^ZDQJfQ4H
aJd\BD3]Q&[4@#(K[WSWX&XVVBUX64H=eR&fCY^CDD.G)EX[MO\15c(@cadUE+>T
PN^7BCK+a0:<g2=TLU.3b3^<D79YMZ>X?A^Y(W_.7b&KH]fa5N)C(>Yb3SQ>eA[)
Ved&JA1fR.8^?OA(QUbB;gT=_>42M?M(JPMf@@J@:&>U/#f3:@;@1=]MR2;[1=(\
L.M92?Ke\0dBW+?d?W40P)2LYW//I3UDND7f59#4dXEZ)E4gSP-U:C2Hd&:/L3B1
_R(,Q;BES171_6GfM/6^D>UWL_P,?0<Ne.bWOH#MUZ1@#I4+?2Q>]11a1DI7P@9C
L[efA>3:aIS[)+,70I>A^<W6F&>2E\PKFHNc\NP18[06c2g6RM-f9_E[^?[A^\2A
\FdeH.(0PXP&45?85,?_;97\:3,Kg<0Db=IDIIJ^A5cKQD]UTUCF<c]98d#-?N-B
-PZ#d=-8-UXe;bL&OX(6Y@W)(S\Uf[Q;TbZ\5M10R_a&<BV8+/&5Jg7T#S=A@E00
^J96a?Q,NM71=#FRWa</9MC8Kfe\G::6I88_8Gg9S+>EY<H\N8YGYaEfH@64&VB7
N[SIPAH(VR]TdX8NdeEB3(W52MAc&&OW]c7:@Y[4S9:O\)MT==T]SPSN<.FK036Y
J];YUF_-Ldg61A^S7BeE0^4Z=]95A,=U/+60K4I,FDa&Vb&3,d2>.dTeA\[TVQe<
X;bVSL.GN?LE:4I\#^M(VbNRX/-aT_M6P&]7&Lf\:;L.@U1W\eK:^L9,&bRa/JE9
==]@^<N][+X>Oa3<+^&Q]5Tg0T8;G4V^P^^PdCCQ0:G:A)MWX]Y>K9M)=\(GK+T6
>_C1.K[)ZAgB^;gSI7^5N@,@eVd>8>:D&A:MA:\?c;gX,#+5?dTSfQ(<Rd/=>0H+
7a,8bc0688(ed]76^RSV@H^J5GT<-6DL9bKN&EO/C:bcF8_f@3X([@&\ULVG[Qg5
G8DA;@0<96Y6>Z7)fOZ)ZVa^f94FL(OJ])+G;EefRMGA-ANKeMSWH@+&Ldc[[W9@
H)a#[=g2b<5A-?Q?_D2-#Z5VN<AJ<^cZ-=(V@ccZXWdQ?]I)e[[(1&OT)f1G;U0F
:;P(;1c>1>-:aF?Q5S40]Y\3I3GI4SYDbQ\Z4)1@HMgT;84W?bfVV.EM):)?Z4A=
gZQPX+?T1>IV.8:(;dZS9_YABZX8KX&UZD<K2aJJL&?WW)#(;9g>[]TXO&5LK3S3
G2CJfN#W3YLea(.:^DaK^16BMI\,CYQQK9YY&JID0I9]S:\UFF;,TU&4C7fL<<.;
,Y/O:E51H>R=-N5D;Eb3BDA?X:7UNI&B3\D8.d6^BR_X.-8IX-R3#8>eQ>#_ABJ)
<_(Q[f-TWg]+:eNb#MT.]^DLH\g<V:LG_JaaJ0V?GXPJMOR<eM-YLFHdCSVR(JV4
[3/@4RV+E3\J6^OENcaD\<=\41/YNEE81.-Yb[M6<2N3.>-OCg(L[5G#HJV5S7OO
N60M1E74W/XFB7?;40:DXGD.>g/.,6UJ.]eaM.(@=Lb;OMOfZb#&;P(U)6A1?##=
MG3&fEI:B;W_>8YUPU9-M6O7W5VGW14_DHA<TU:8-5ZbKFM@P=2.8G711;1UfUGJ
>cL9/YY<f7WB^5?^1O#=:.)U0)E?GUPVR29W,D1N-WJ;;D+Y/<3X<\&D#]C1Ag0X
T2e\SGOTYW+D4XfONROK#WBH2E.VEXAY\9JFNV/))_CgMM>15<:RfV41SEB<L0aN
P_.\J=/9_#KV6R@f()@7EJaYfZ&efK^&G9G3E=Y]Y-_43H3d:L0J3(09>8Z2([Ld
#(8XD,bDW@#A60ASE+[9=3357;bZ#G\.,F8M7a&^>/_80HOIcILCfDIeb1A0B9E\
RZ1?>Y7&6A0A3):5JTdGOUX-Fd\#0MBASCMW;e_62)G2MHOd..4g)c1DL^+gIQ:&
0b#JCEB/:/7QfEG;M3WJ,ObKDe7@eW6@PMD35>98,gX,D,bJP0W7B75LX/:OF/23
.XK?2,/EdegH4=a_UP)+cZO+IK)+0dN)\B8P&Hef1Q0O7>G1e7H-/HU+e_Q^;G9@
O4)0&dEG[IGRD7-f?:9N(EB,DYPV13NY#B[R&T(?/F(IB.?Y9KEJ88G^Na64\<.-
e,FdaQB>&RKga:/e_C2XKcM8<KU]C<5-BYK:?J97c-9WK6b3ISPgY0J9aI-V@4,T
7d:)eGAKfOP9LO_V2]+_7d&8],\a[G8AbYc(QR3dV]P/,4T[-70+(gY2\ZaEXMcI
&I=3)+IgB[;F#0.cKAU&TMAI]0R>gE8O&=Uc7MTMND#,12cc<FNUcC?W=6SR;&J+
?f<f]27=dCUG]a)bN@4_DI6I)aYdZ-#<.SbTbVN/?aNZX0fPa/.ET+SGb)GB_>Tf
OVJMcC9M0FXA9@O,3aQ94-D+^\7WOd_FBO_?P(1VLV4369+@<Q/JL;T2NF)+(Vd0
W&JKYHT[NTDa;TJBS.-@2cb?^5Z(.JJK7<QcMW3>dI-Q_X]PIe:-\FWPLF&J+RPI
RM3Af;)a_Q50H@gEAHaLYb4/NSFdf163.,YX6Md7WCOTX;AVZ03G@/8\WgU+IUB,
.P,MWLBV,[R,;A?[1Dff@>X=/?Q9_TAT7b^/S168V^B)XcIK(.1T]E_7T58f<5a5
TEZ8<AO^AK[DVd\=7UK8cR:#e4)FJ+9T_GCA,5T]U#FN(O@cCCMPV#-;d<GM2=[P
-:E[WNc.7QZ;-J(+UQK@]IC:<9JbZ^H7Z9X.=-=C;H^46U&YP[;=Q78J,5E81B>\
HgD7HD7]QK02fLAfE@6QWUITK;Q),A89#UMRF<0&0)Q9+ZNXGA3;S.7ACbZZLALJ
bHaW/<O2TB@5^LMW&9]E2AKEFS;M1Z=;=@8MC/d:f6b/RU\L:FEDf3TP5D@Ma[>b
K/S[H7aaYS4NU?I9#6d:3:eB5Qb@_0=a)[>#K@Ie5J<9aM:FMM^]Y^LX@.])9:N(
J].A6EWdCZN(U2F>W@d+U]2F>9(77L.dZQ<^9cXL<05-L7WL5(=P_dFJO>WB4Rgb
g=6W;EUF19/[E+XRAf\YFBST(6dNR7gcc,V,G.K5g9(dE\5=VZ?&BPCV#K7LDc@G
&cTGFD/]4_/bC6HeW7Z#9F47R>XTJAHK/0=2V@1NI@5EIb4eLRF]A>^IFaEfX#@>
KD_EC^=06NQ&1IEOU[TFZP_HZg^#=/80_3aML(F]246.HSJKU-OE[)PVSd5,-B5f
GS668Ka/c4D<;]6]Z3e;fg/Cg1&d.3Y>BDOD<e\Na.7Gd8C(OL2T(dRB]VTa97)a
IS8^G(;^SR]?fV04JL4G3MfM3+(YgGLaM-R@NG6Z3S_](?fO+8#B\Q1U;/P@A5,#
WGbN-B:KU69S06F_?>X)DPJF6,E?TFgS^<=DW=9>0-T4)aV(LJ8P94\SWU2E((=b
EeF0N?Z:7/WL-#F6&]U,C^4T@I,B^:KZ,7N9/72).CWF(aR0H8M9<)Z9fE1A_ZHG
g=T<2WN8G1B,gUeg4J;@g<CaCK_V<W-S-7<e9/gXGT:@Nf8BL]E106V0IMf/>X>=
ReL(>6DO+&:F;WgLVYXS\HGYA:52He(5__#GL)6T94;&NIb+ALXAL4d9DFN6gc#e
Ie?9a-HfZ(]EE@TR,748@JWaHO+6Ief-0gSDPF(.caD&&J/[>I]=e-.E[=I,#)eP
YJCX0cccAb@LI/4gQ/BM]:?2P=>E-6c6E88;#K@/]3>3Nb:AdH=2JD/,)A/RL54C
c]:X0X&e:HG\Q(VY>L<;EIFH;U0H,D#g0f,)If<4bM@T2,8bAcB<d6[(RJ;X?Y4,
W&\_V=2K:F-\2(S[HD\F?#+c-#VcfCK\(EN;/5;Z\W/OV8I@cd1L@1KC7Md&(-@f
DaBD=>V/=Y#g4>;,.J-@b+;4J94H^P]f<CDeNbYW(Ye-eA3MeBPeLANFK#.[4IM5
EK_M@690GV\Y+AKfHS2C4e^UYIQbcEI<fY5.K0]K_I]c.33;CN>674X<54aBf-#K
L0DSJI=VW>J6KO\4)E>3AY>DVP:3>-EbH>?F,c-W-LUf(_5D?7X,g:c.g;cf(I4M
J>/LKgY<=eQYF_Db[df@N2&C3F:2dRKHR)_.I4S7\N0?:80B1:<:^-SM)=c+?fZ?
c?6Z6;Ya)#JW+P.&]\A)[IV),(g8.(MKJ<aDSJ4>)-([_-D0Td[T9Ng#U,AZPTIN
H]B93R^Hf<D[ZU5Y9]FRP[Q&W8-6&IaOK.:bYaO,+^I9;E@?+]=),/A9<\>;TPe_
+_[G@NWTY0@(YB5GcMMg_fC=E.QG:JTDCWBG:Xa2(#912=e00cP1&I=U,@gc33-Q
T;Xc2I6f)c]I6aM3^QgB[KELW;5BG=Q4?=]\^+[RAH35)OS35OM\TT_C1[E4VH^9
Lcf5I#V#f-1gT8D7;(7)Sc+X?Zb7J0P>.BFdK(0(Y5aR6K\0aCb>D06CWJ_?Wa(\
[:)2d^HWa.[1DPX==YB]]<_28=7b,4a1gf;ZLO<GEUe;#A,=4K(QQca4:c),3b<2
d)KM=4?(-M#W/ZM-P7O[NGL@F=F(<ZQ7bY1J8^6F<ON5WCZ2,W)b[-XS:6a;_=26
N]:a@ea6OMF,?4.RcI#SR3PIfFE-==1WAFQ;TFeHFRA/7D50#H/+QMB952_FMSZT
7]/LRcBXg7\MQ08L6G7gK87EGb27.^VGcQR+T6aBfLG-Fb.6\1L0L]EK;eMOSKJ)
d/PHWfNbY2\VAP\1U_H/M[eW(=Y?g0?A3fG(=YVd9JgC+(Ag:G.++N,A&R+S_,+^
5Y]Q]RI5/-^=eQC1D)]g2B]SQ5YNJL_B[]68[UTKc--fe2I9T?7ae2g83/WLeg&.
7Q,71XIRILR0NF6X:<Md9CM[7-\KF4+D1Te)GXU1;NLQ6.B#BaE2a]@L?Yc&<=a_
aJ<5EM9J\(eAIS3)][ea>YHIDA9EA:eR=3a>abJMJ><aNKJV-1K^]#2\V7Cg#IZ\
Z/a+?R,QM:YA[UG@<<RJ-B0acX)?1HAfT6CAMGg=5D,&-2X3]SU<M_Z<_8TWDJMY
K,;>6)TMW]<>N[/g]=VQZ9K,1dW]5g9PVVJD<LgPW.8Q>GT0B;@VbNCWIa/+#@:R
8c&QdL[9M4;PG293<+WT>A>:5?8[S,W#FL1.GO&:_XP7aD<]/ZKU7PYScY4(Y\dD
4UTf,TYHa@94K[5NB>)/0Q/;aM\BJ[LE:HVXaBd[<Sb)Xa@CI&4Z.Y6EeY&LK_5Z
-&-(0OXR(G7Ng)PES4OAV;/Z]W5[72K+La1\d8b+/(beB1dedc3Rd51KV6R8RWHH
?IU_+(b,8G=)E+Nde./,@N)/>X[L.?5Eg+E75(aINPb&>@_WVZJPL4JFM<DJJ\eP
+4B]DUZ._M>(>DXAKA5N.>^TJe\-XS:SM_:=6e<2FY:=ANcf9),T]/4WG41J[V7a
(e@RQINZ<.-IGTf]>9:,SSLceFC]8AC<Y<=DP[]=P.bR03IDPXg94^<^cb45+E9&
eM_=KebIAd7Z89W9GNTIG[K51_Q(UB_f:JQ3Z7_J:,8eBVDG=.=_P#(&<.Ja5)GG
3f+>5#(URW[PDAQ+Z<P&PNfQM>Vb_?5-/cWEd=Y5,bDf8213EN(<R-+DC?d[UMJN
IDTJP@N\5&[(W9>J;Vc#7Z2EV8fU@FAFbb9b(@<^,6Z[^:?49?>XL4bbeVEg8C5W
eDBUeBLD>N2FZ4+4FfIg#IeP1X?EU/<P#>+WeS,C,]g5)L.f=I#S6NDKDcL4fQPf
\8.\6dGXScP7Y7RN9@a3,J@Se7[R7L]1J?dK-3EdaBH296f0>;gKSG_AcVH6GZL3
g6Y]5@<-eL2I2VJ60#Y]5R-GLK8ObM]eAC7BU+&BS(b?5.N::C#e9(=ead3K]QUg
9L_AT<;\R]E4,>O+;:T#-?/Y?#)WVWAFf(WeJ3Ye98a:fC>.J&c)VbeD9eH_+8If
IH/?@)LaK:B&F.g)d-9N]2[(<A@#Z5Y/[(ZW?_+[P2:^.<XRe^g:M+a//&BH:M:b
UZER0[acf>&-_.J;FFa=Q=Z=4D.79dJ8<fFaR#7O<[CDWQM=N#RbK1\PI8Kd1@IF
(bZ/BO<QIGKb>P>DO[RE,@I;6@NMYg5#EcH-K4]&#VMNL]8?1WM.Pa)E?I(N-SDP
37=V-dW9:JDE4W:O[AO]gV?PAJKM69bWNP.ADWQUOBEBaE<@3N\W5M]&P)8Tfg6Z
SC@6[J>8X:#]X55A#J,9BFJg+;fc[BK5.K)cB5].OQKf-B5X1(B;<C[bB\[aHRL_
-+181^-94H]@G[:UgH_@U+3:A=E[\5DRZ.)FP\)U70@ETU5H6NW7d;@HL2PU0IP:
LL3:b8QgGDJR;=G71bL9Mb0W_L=-\fKA3;\G6@#FV\?E\d4_Ke<J=cSSM6-J,7=[
1;>W,3:)A1S91dN_,Z4@D,aY#V5V\O1BMZ3:a1X(+I<K?VXX\[aeF8B5B.Y^K;;=
QBGfQZ5GfgAMEDR/fcQU+GYZS4aHOA[9d1)2J>FVH[H,O+:@R\WT0X?J.FVb2BZQ
W?SYEFP@5WSWV:PE,S@Q?Y]&JcRe=C:]cMSg;3YZcO;#YPEI9TT&Y;VM<;gfN_T\
.FTIeY1dXQAZ+U5^AZ);:aE\gY9.5=L256f6QZ,cUaa5H@UQXJ;gZ1<ZE;Xc-F>0
&\@)8ef0AV98VNHgcVI>_19c_?(LJ>/gN40-9?(&RMTBSf[aE1(S8^)fJD]Z4]-;
F6@M?:Gd-KK<.7BF3B;2<^<0B&8+XZW6e>g:,LB1Ef5g[U(TNSHd@JfBWWeS9FG?
P@;.d>/f?6DP:^J\G1(]WcDN)03[I[^@X/@64<AO^_77&9Q@.0W:R.P?6?5I>LDB
J9]g=+=]Zc_82@g)4G_RCd\+<#.)=]aM1b(8/f3TW]X<^B:7MFYQHeJJb9bTA^N&
1RDEcABPa]f=+fd2<<bADQADgIDWQb7Te((LZY:,VbV-ZP/S0,fgFd)>K\I&A&#>
:B=05/a#?U6SE/J9+?TD9AIXTY4G4e>:]EDI4YZABOgcO(\7IE4+A?f[.4+HH-[a
&IbQUX^=DPR[;7N>A+6D-]G?HMJBG+;6KDL&Og;g\3/WBQ&VQ+U6>DJd.D:He051
f@=X3N547@Y9;AYeB/N[,Z&F?Ucdb4KD6a=OAD<L(5Z>O)fQ,<f\U4O;S8MYA<Y/
92@51YPXP_2g+L.YWA/DA>6&E4U6<D\Ba/UD(K2XgR<=\WDD6,9(e:4UJXbOGPEI
^9=C@5MgSEVT,E3-#Q=beC9B^-+=ZUeMe#(C-1KM199DC@XT3LQ];,1<J?P0dSEP
0gMSP1f4SH75E+E1fNLTg<#OF6,Z;_U7,I.3I:TBK:UP\Q@V45KJLPD_ITYBJ6Ff
+JXYX?K(/3RJD9UdfYDNCWE@7MP449OfNagA5KCNVPE)],9/IbB:J([]L+P=5>MI
P4,UV/PGY7;-EKZI9-gHC8aAP7/[KZ<AT)a#=2PUC,W/F7c(6=cC]^&A#7[\^71I
KFMBM0AP5T-0<ONV#&V#Y_@VU,N&[0/J?Uc:K=M2?gUa-ZeJ2_R1eF8;gARL+g#d
(7\SAee)FC+)#a^Sc5TS>X(-_5QR/0D.+6B7E?7NRe=8.[c);V7e5((74D^XR/;[
J\_S[Y<O#?D9aHPW3S#(DD2f^[<2J<)E)0NJ@D1)9>#^X.[T0fL126eRI3N)VZSQ
G)(:eID)F\-5P3APPcd7JRf-)A4I.[[bN)_5+Td]PT2U#<+R>C=@6?PMeRX/S(>T
c@W\gNG@F[+U&YX:E2BY+Mb=&<A9K<3XV=G-D85:?6SPSfQEeSVS,XD7/(IAR&a7
O\C]M&R:Kg/C,Z]X4328_Q:WT6,VX;;<\=fS?NUf2,1)G?JSaAVRDVW/3>V/+]V<
M8a/5U@5aBJ/-<MV\eVN([b3)B1;DW(_?)JGRQf/Z4P&^6+7H7HP]1H5K:I,,JX&
&P>VN[0D[#1#C?-)T/bK9?+R&cT,bYEf,bBHAX=d,<WUdb\d@g>VD..JPDMSPU&:
YbP)#eUA()2FScA=\LH./b;E?dfRbDB1D>00#d(66[I+0QcG<?ZH20Y\C@02=aBd
HN@B6QPeS&KcD:MCLBTW[SMeICN9D/QR+B_U=@c+VG&X/M?C=N3B#YgAH.H7Hf:@
?KgKT]MLNK9BYZ\?B:UQbMTDJZ3RM0\RCd_S@ZOVRK4^>AgNg#eRQd]LTBG-cAJY
aaQ9-FB5Q3O2]]I#c+e^NKa+^LZ9;_9.<Y&]NCFP21RZ>&X9.9?7?Ub3)cF7GDg0
4gWKDXSJ;EdbIAQ?,WAEVCfSH[b743_\CbM1.9Ad:.JC/XU:O6O2I;Z0U(8\^aKY
U@cR)O]+QOb^DPZ-::O@&1#LP[+H9N4@?O585.2Bf?/Q3OHE1./R:3cH:ag(gXb+
DMH4V/9Y+K?_LV8A3HC@\L7N)d8Y9R/+^OFW741+T=P_?OWWX#</7YNB@&/9)#/W
7Ge#^,)>Q^1W3.0gT9.^0@+?8+2+gd71+]WPQSJ3;?ef4(bUd0&/1#U5&C.Eb_<H
KQS-_./V16;DVegG2&EW)[1WRDQ:ZgH]N&eaB680&P)IYJUB\/XdL=&U2]D)I9gA
I9_LM?CWKNAaU=QAc-#MZY><R^0cZ;^C:.U]?;\5-OE+c+2&]VFVC)S)I:f30=e7
e2cYg/gGRN\5>6SQ09CHgHM&;e,G#\2U?.>79<JW/0Tb+Vg1[c+GGPO5Q2^cV8e)
D=#;F&=1CTCFS9E4#MF7#;3POWJFPQ7e@,F)MLP&06ee<8(RI\PPQF/P2->8HWZf
P?J(U:(R#?8,@=@:3a[/YKaNg[3BV>aB2=1>@^9_8:E>//aeP=:6dKXD][CfUM4A
#f5O[Qd/c+4J?1d0XRH0Ia9G+BbG8A_UXVfDcE_C-38TN](Z;T56I/0:;0L4(fDe
Z&4>K;FQ^4_^04eD5aW&+bOd3N;_+OfdQZ]N1gT:<+bFRcQ3)X5>X[P;B\ff&^NA
3e1^W)7_Dd6V[?PIK^Z;P5Z#_]/B1/M\YO2fY9XFPc0L@]92Ibe^,&_]NOHE/dda
O#19[9=6.dg_gbcZE:O;OWW)gV=Y84=RG>f55>5M3POf-F^0;J+/A#C)TA]IcO/R
TS-L[Q<a,7=#>L9D+-9PBN,W3BJeWb-^b>^V\NLQLYPDS12Ad?8ZO>THPT:B_X]H
XW-)G5Y4-ZT_YWZJS332(EXR)Ve/E23_(2\9O)]#80UKb]KJJR_e0Q(CCEHdBQJc
),_8c9Y_]#L>HL6#X@afAFKf-T7X^,Y8]\ROK4fZ&AE5U#ZgVNPO0G4[>8[AQ^Ga
GeNJC:[<gE_EK[E6Z2=MY_(-gRaD6>CZN)R3_1-7g#O.I?(;R66Me\RB+Z;?6cF;
#;R9)+)-H;1X,cM4cgR3(6PM&_W./3c4#W9a=PYLO&^=+)dE<&G4RWN>N>DZ;,1-
U7?^d=IIGBYIS#@UWGdK15V/[bU;JT]>f>XDL3Y6=D30PVHK0,2RB),BFEP5./Y-
RYV6D71GJ,SG3Gd16=G6&6&>DdH/F47D-\CYg1YI/N1Uc>;;a+XQDLT\EYc[gGX-
2\5N.C#WD6>d]3Cg;d^9LF4(]4N>><cMa+QSS1<;&/6H_N4U;aPS&Z?22/e,g=Aa
=YDR2U\=ROJeG#^,345V322<QXDMd;<XccISJ.9AZ_JaaY\4ZaAH?HWW<P[O#5N?
SMBUa2D:R&;ZS8;b4e\]SN4X6-?TAG9gGGY:.\((H#RI1DO>KKae=cP+:)?Oe?c1
J3J/[P[.HQ@GF;L(\&3DDL[gHfE9>d\0BDH70OAHeK&O]AJKLPB=34STIY[NOf_e
bZHH](&-bH97HF^3aCTM/NE#-IeIc\Y3LKS_U+[9^JY#T?,Y/S\X@]XO@c#Za:d)
2QJ>(b6<BO<fWU.93089:.@)9NQS]]_.GK\Z#MF4FVY2;9L.EX>cR6-\YOL69V.B
D_#f^LOd1[WBc2<.#OO?[U&BNR+3BVcc6UcWTSBVb951@I4DaIQ-Z1UNa;^1N_Tg
e/LN+O3_5-CFc+9Z+D(KSQL)EBHHZX8U/JUe+N84K[)&(?)&5c2Ee7_NcPZ[KSBZ
YT-3W<46;<e)U-aAQF(A_2HP9X^0dF)fNJZ^(_O:.Q:YH_fJ(D5C5+cHW\\Ob^BF
IC^+d_g2+dN.RORQ.AgQc5g8WIcA#P5++cE\/V\aPU#@G3.55A\1EQV]/F>U/gCa
XQ<X0)cX6EV,<.B8CE0dMdDbSD2;T@QE\c[E6IBBe3OFHFW+P[A2)CZI,6gTZ615
==bU-N2[-Pe_OJT<:7H58);@:_dX^9H<VDaM-+@NEW5X)0b\EeP\UO?a&34CL<J7
^&\1EgXY,D-a&RZZM>O+Lg>2\CE/7I1OG3UfV_.UCCVea.UcTCRfPeW;)OgUO=OT
b0W7PdF3_gYU1H51JQ^VJGTTI45F;^bT4NSS:N[.J2Eb&TAdaRc-1X?]4B+UF&5]
aYK0a?aag3P7?S@eOSKEdQeV(B<9K3PB7+CGF&V-IY)>V(XdW<_7?/MW#)7,+gCV
gS(;IcAZZ8Y.O?;C]-6fV7KVa0[FY^Y)_)gM15ENbRHSfEW8V/;4&RR&IfDXG?SS
,>ZM2@C_J-@614cT&8aK]1^Ydb+79eRR1Y^?,]NQ\^PW]8Q=<3AUMHfNB;<]W^V:
+e7C?J(K#bOO:9C\A8QJMad\2=7>G?C&]HV-2QEVHbW\^@EbZ.=cg_OG8B)AcdN0
I^<EPB-X)-DO?=^VR)-TND)<LSR=26>O2ZeDTQg)3edD^UN^MgW5^7f1F1H<9M4?
)LHAgfJS^//_3>0f7#]H8Y/BVgaT/;+-b],?H@?K.2M6;K@GeGH;XA.7,YNZ\b91
a+@+1W+/YF;-.YX221[aW2JS=KAf1/U_M^P:R3FF-X5;ROd[01E;<92V55UV7,=L
0O^+@LF_CUL-6..\R/T^KY@F-^7Bf0UYK5P_cM:-2,4GIEYZ-8^AD)[RNS^e&I1-
6R_SMO\90B\X0bI()E?H],N;P0aE8\^(U&[#]1)FbN&@@_5e9FS2QKHa(30)47Bf
\-SGAO7B_fgK+_#,1?:8DW+=NEPJ1aI[)b>WF\[Z@>F:eeF7IODYAA2-fX6(\aW>
Rfd16@;M+\g7O]b21a@Z\eGfd8^:3VSTO[WU@RRd+VGV?K4>CM[WRJ24X=ALg5@b
.Q82:P5P9?MFARKB:@6#;IV]X(4K6X?c2^#I_69<PF(:1FTM-ZRaM][.QMX\,5<e
gR,4LDL>),=Y.(ODK-?.]P7:&XT6UaDB1Q)BPH)UNYKIGG[.(G3@^4FQF3O=W342
Hc@U+T)>RY&JTYbW3[D_g:DQ:S9R)R+1(2(AU=Yee==)?OAG,2IYK;08G94C8@cV
eA8>0D.K9:W-WAJ4RT[U7;6S>IKe4--NS?V\9[AB3^Eag,880RN[V@#C[dTgB.L,
<\5>aB9AU3M\Q=V?I4^:U;VgCEDN>ad9]d\XE(JU-?X]45#2Q?B&b,-]3&BI5@#O
GeOK2L_[E.F[:N3=3NVgKOG)R.gRLE7@XUNG&\f2C+,&IaQJ.2(MH:+JLf?G#PQ2
Y8C>^8_Te)WZ1eJ>C;6FKc6K9\XE;X&Sa9:3()O)Gg?C<,\CQLfQ.T:]P2NCJUT_
=?&X#:3;G5B[NN>:O6AH;28IeN>&^bf:7H??P>_T3@>cKENZYWc/fcTUM,KKQAH<
T]C]5KJ?LQ#BTK3]?+#&6E,UPNdg=0Q9B4V+5\a^B2N\<F)9+ET<XCP1g.3c#_Z&
a9E^?eK7?LaBI)O<1YcF5R>O.5Z<#M_W;>]Kd8VQ/OA^7H8#ef)&g3N9&?Z+8cBc
Z;+,<-cYFJMXgIQ^<B1Bgb04JAVV=?_Ra+\?9+_@8H=C_HUKK,4PVX8fA>,-_<-)
4N17:9e/R1NaLC<(0D/HKNagf7/IMC:_&O-IID\@8cJ+.B);^T-ePF>7fWF:N]<?
<Xg3gAc1RV2JO5;Q0^-be.E-;>d;V(,5.U&d400?MS[&=W-,UY,C?S9AM.GRg28d
c5//5=VS-Lg9<RNW3cC;-?(4[b^<&8QDf?]H8-NM_GP[YRG=LV8;SC3WLL85=9)X
U(S&1RDMJ#eR;\Jfc+aN)\-NKJ#7^fSE?2e-D0c:](1Y(ER-XC@F_:-Ie=^fTe[.
VCUZ_S7XK\@-CE0F&[GN4>b&X5R.F?V].Y=>2-#[5J2#7=HE#MQ+;VbW2&=.EFbA
MUVM8DRJdSN?V(GbLW?5e;0Y]+[GMM0>g=(Y.NK#QLKCg[H\E#c3GW(H.6I&<U:Z
)e6\=V#9K-6B-N0^K?T8.>.dBdNP#WZE8A,d.POU9f.G+:C;I3bPANcLB>S?+5b^
/@G919N_FBJ:^W1IRWDg:=2Xaf:;MZ^b7:A<e<27U<KI6W/fR=(aa_,dL_a.+5#_
GP^V;fVIRXSK@YR-_C?=GGLU\.,F]XWcb_&.eM9b;NPOPa#X5TEQ5HgaBgFWDTHP
[+GT7^4)a3)ZE=XYMg=4OC4NQ5P7a4\g<eKY7)e1/ACNcg0PQAa7W:3-K[eL?/Y+
:6U:/8DG8,@/@T24c_K8+=\g)8cL\f12_B[I=U-6D<66KF90(M7gB#R=g6014PFK
KE=JEaICS?HEQS8;U4Maec5IZSE]L05&R:AR^O3VW-Rd#0@D<4>O2#4_K5M>T=eN
8MMB=b1<^B.G1=-W>S93Gd+g\&L^U2I6[W=76?W.Ua?EZ?L0#0:108c15b3gVPJc
\0W;;aecO59SfX@\(C;SDEY@F[_?Y&+VT7WNgZ8,TH.Qd=)@a..OaJ3R=WGf=/N#
<??e>Ic0(2EI-PQ&.fNEFB7KCQUE294[?E&>L;.^[Y\?@M+1Pag,KUX9.9\UMd;,
H[)8bCbCPO5N6I-T+30&=H#AJ:B3162^M_e#FC(Z5ZaeaC4eZ[X@G+^Y[bfDJOb.
D#J:XNfI92_g2GH]E:J\G/3DQD<O9.f56VV2AY+(2+3K@M-2f:[[;^]X\(b>5.:J
QR>MeBL/MO(CWeW?P@f=e9d5Q2^BW-D^We_IIZY-c=I.YOY>54<&<(bQW;Y^R^7G
Y?UC&SObH-XW&[2OGYZ_(Ae9_:KY\<@3@]ZQV7a:YHaR2N6#[GaZ<9M^7Gd\KKb)
aXOW;ZT.J-HB,7UCN1XU:g5]<4gg>\AQe]0KfRV&.M;2]&5UB/2PY/4=EPS6d#FR
46#W.#.c;H/8H?JCE:1,9W<R.#aUC=]c-[ec4YT>B[BNNI&7?RA^C?W)5+eZTDK0
fEOX>EZ.4PeGf(+S5>,QV#UD:\VL>AQ(:EgKTHN.eAbW,8)fT5>]^W.WSffg\Ic9
XcdR=R[4U[8/]eQIdV.YX&8(^Z\3.QHCY;_aD6N+M601V0]6+,I:C3eY@-)]>BE]
=VE@[,005;M^Fg4Wc[Va(P8Q,b=PW.C4WOXL_S@T?/6>d]Y,Y;<E_N]A>GKF^FJ<
6)>_]X7:/Y)Gf&:45L-H5A/(HEOaE0T1/Q64fA+(1WR0)PZcTMUIfTX1.BTWM,KP
9;#GcQH9,7fQ-XLL:SC@1Yc,Ve9c<&9#5a=TfXQX3NgL/-2Ke@fe9K[@S+>6Se7>
5e^N26E5X(O^cBN29_6_=R8)^_daZJ.f[J]&ADP[FU>IcS.(>[6UGI;&bI+P7->;
GUL[EH#JR8#XF@;A5BZ6;dd;f_I6AVFWDcZ#6C<_=Z<V5XV_BH\30V+WD@U+0TB/
]NCZM4\TbLSH5OFbfXNfB]KO9IHQ:+C#N>[-:(IGLI(+3Me-SUgNX;UcKFRV;JSX
AN/N8),L+J<@@&0@DEF9I/5\9//b5JXDM3SH(5ENc_YFT,_49^6,PH]4IT=61V?#
g/&\/1<Pd9)(NTa33=2<Y1GW7<<C._6#1,_M.O+XR)+D>@Ab6HW14d7D0IfIDD0)
;J9&&P9dCgfAZVQ/9ZPXO;D^Q\#RM_J?;PQ#?XVe&ce(C9Q-R-g:(;99Z,59[IO2
(2#AX&]HC6AHHbf\.C8ZKgR?S+,.OfQ50B01C\5L>;b=Q1^#OcJRePgRVYPQdJY4
AD5.KU5;N7#W^_W+QKR.#9\IVK[IZB+A>4<#V/)f((R0?^+R&0LW<V[+W>GA;P,I
L(6A0Af-C\GJb\Cf52N67T84X3N?5G+(BDQ8#KWL2(18Z?-ZO3R@](-aCCQ^:M^K
Z;C6Ae.#D]T\UZUP,ZEa578H]DV[\]bV\>R)Zb\UJK(#LID7WTY)D(J_/;LLI>3+
BBM2R+L]<&L@VNO#4:<\(/e7MYMQKRQ_A32ZWV9gf]42O.FVX/]H(/CY70[@J)c)
KWR[.VQdT323&]:I=-Z@L0]b:MQIU=^/2VKc?\O<WEfV?&Hc;EW?g\QcY(1/U2ZU
BA9;g]1:e[d0+AW_];5&aQH1GH/)N4+BZO?>G9PZMWMe\c2J9^O:A[^2MX;Q&]>W
.cR.dLIFca+\H3#^e(J<Ba>FK:F9C@KGb.ZKf]\N;2#f]dX6MfK9?.&U\L?1FVR5
PL]&-F^F.8GcdGY8M2>DG2)6B-2R<W/CeI)XK.)c^]^IZH]Z.-=7c0]75I3]HJcL
VgX#Gf6;3);5+\T9V\NYKbDAQ>ES]?(+60=gac7)G4ZXCOF7I,d6H:MP.EK&OG&H
C>B[(YD1:]9D[fgCJ.(\_-H,5<<>__GeI\FZGV0YXT(BD6,6/,/7^b+1D(c>b]OQ
4,-M9#(J?H1LVBLT/24:J5Q]:=,\++H=5BP::O&I45[<SU;L:048\P@aTWF/>&TF
#@Y<L^J@WKW&MZ5^AGS22J)Se8]#V+eXg(<IWL\\AYAK;NPa63@]6AW6=E[e1DW7
FR\30;;5V3A9F+6<Mf2DOFI[SJ9:^a;7]#RUb0ZA1C#5RDXJQ4R89E&0#Ag>XJX5
<Z+]-3#9P-g9>-+VC&BW@]gPZKNV:gB4W=b/SgYdJCSO75bVdT2?OY\\VTg(M6,J
@4.bN;Xd#J-UBS_c.,g,8B6Id+YH#aZS0E<RDN)Fa\RK4:Dcb9CPRPLJ,=N:IC4)
P^>M4+SUN3g#X_M23>Je_-LH=RRFKG2?b-Y,;25B79=LJ41VP>.g5G:4@E(FV=bP
f#O#77<;#=5J]7QEc,W:>V>_@SX:@[.dABQce[F)-L.T7GAbVd(Fg>SbL9(<DJOS
^XPR3cASa[1=IY:fKLGW;/.0O=f[HQCf54([8[INd-VAJR1(S+Ld#bP_:O9YN[_G
N8>-[J=,\H#)0_(8)H[P^Q0@X4TYDF]eJ<-3&\ea5GZGKOC1_34FED,CcGW5J3Q8
P\F7S9Te=-G5eJbB&ERLSa_&4XJ.B^/TCUPJZPH/&E]R);5NQ,e&:_?@V^@a+4E[
M3DGWY503#7N[:EO7&P]F=E?IKfba:?cN1@V4O@MNUVF[>a4_(#;1(7-4BU0-C\#
3>eUJDUJB(I_3OV+1L;Hf@1:@Zb_&H&3_Y^L3E>0FZAN?Ye3WC;+c<Q]K9\15R]1
+[]JC)68c4+7=QE_[g.H1<:=++ab[20Ta2_HZ@_+>cbKXMHUAIT4fEB-]0KTb8^4
ES:aQ]RUfJWSM>US^cM7HQN^UQ0M;SgN2RdD8X/LJHJfV)PAL>=\a&/ac/@)g6SN
XLA;C-RQ5HfXDP?-[Y2;U:S)g(G1U318P7])AH:4/Y\29QaeHDX9Z[+Af6^(?&P[
9UW5LC0/IZ9IF6T/US6Zd=9XNM72J([c#=RJ@:..ST)#WUcJ-;&.5J6A4<?W,S.?
-C^WF4f&2RRN9H;N15QYD^6NT[:N?T+,d^J(75/aOYd7MT8aR[RPL([702fR[BU<
_RV#678G>Be>,?Re;)RAVY4D9&2YaOZKEX9GJ@RCX8IXe(,TZ0b,YBKQb],YP.:[
-^H[,2_#(\MaIYV@1dJTWXE_bQG,3G6P.)])6CJCe/Y-ISLD=_9Cb.Rg^.e9,AP9
bc<5IM-Og52Z_[d<C+P_XZ1L4LI:f],<[\ERfSgD/8T2_\PK1PTM@e3ZR[c\dYbD
_gX7-;.,g)?446DV@Lda\&,=dbN_ggLN3&=fZP.:?2,?0P4+[e0KNGNSBCT[I)6]
G^UD]CJZN0;]),G.R-]U)LUfEaAU:?T/].XAdeQ/H&(aF?YEMeDWLDOb#JF,,1PQ
]UBGW?;D&NYP-G[fAe(L-@\g9RYZgR@@eb/GDL?0=Oa.;NI)C(Ba/9\)R#:^VQMQ
\KR_ZIZMgQ_KE(0d^PL\X.7.94(baMTEe3-c;GIDTg3M;&K<Q1Q<1W1Y<4(PI:OE
2NZDa[J38.Y36)=db>DSI<;32L.S;g@R@>A9ID8\H8e[H,Y]N@<0(<\]ORRe<2U7
G?LS\DB7&7T3gCFb_4X-WZfbE>I<a?H>:Ag0Q)(_G;RbFfOTafG3<L4-DN(Z+d@D
>-WUDH27bED:fJ_)5JCS2fdUQKX28GWQXE4Z2F<I6BWUV[@_]2BXQNV&1ID3)QRg
d9_KCe_XOJO71ebdJ62GQFZ#?EY0&C4d<UVX=@_;O;^#Sg-c/-(SgDD^9aOK.c)g
:4:3(P,/-XY21fQ_G7BQU[\.=TD]3/-3WI2dTW9/CFcTf-;Y1C3HFIgc2)cA]9?a
?96-&2J/P\4d-K:[X_18DAK83>J98K#I^.R8V[6=7Xg_b,NR<d?8P;5V(.-RN(.4
?,0PN[N==65]@=dH)a>=2dQe[.YF@Pc]gd]/>F(+Lb.@.:9-4F=240SSRHW_FV\@
4#d#,?<#_9M]X?]^&@ET.QXed2f,-3_;XC9I?7[2#A=eL>ITO/Z62?Y^;gW=)G:Q
3B;Vd.V<b(7)5Q-3<f+-ae^74;34(,GYdA#a<MXIdCVZH23Y3b-2_N]CY#C3?=;I
1A=d_+;=EERWDTURJTEfF8RZJ4>-af]#1)b<5IG6BME_M#W&/MU+TY+CMd2I[3L&
&E&_aP)dAHcWX9H_QBH1JS<9LOCIO+1WU/d8#H5-a25g;YeP]8+<<8:PC.U[AA[A
DI[90Z1@W6GSD37,8g,T-6]O-.=+V2[3<&.M/9]JTe5)<I+B-6I\1(Y/?:EZ->A>
XATdBD&U#?_]C^GP?TSZeR(S=D2R.QfE[NfX^?#MIfaQWA842JX;R,74&@WPeQPQ
Fa8d7()EO1BY&:_Qc_a:SQLXX7b+8;NSA<X.bKg<3]QKgB&JNP+&CPd::1)-W)P8
d;F5\:5HgXS\R6SW<E.eMMeQF7;b5R1G11>UQF4Pd7MV1Z/+PEMTB1A7TO0c5Za?
]gO[RbeO)OV1]OR5_WdKRDCP+C2I?)2:J2c,-Q&L[>M^MU+35c>L-^))c#cX&1I[
OXI7b.:/A&aPD\<(8fG>28<KSHZ<.Za;1#0,OY3W+,NfgCYUN&dCVXNU[<M^G-VQ
_D\;A5KCT[4QdU+Y&bZWU<cR&eZ_U_MI65N,HX1&].,E@B_Mf&1FG5((BNE^O6Xe
S-NBCH5:+D)H4FeMZ8YO;fc;@M_QKHN/GA;+HE229:6ZIAN+dIUReUN]VM/cMNBI
2=/8WYXG-a0bZ[ZW76Se-Vf153U<7//A@K#a3dB(@99P]\@VUaH,..ONC1;^a5NQ
R;][,U0_Yb)MVR8U4gR)R,CFg8gOAAJ:T8\#&T1]JTKL-<6J]T+(GFSGb[1T+F1#
)_GX8AdGgJ<)\WQLE[Q)A#H]2I.FdO4=#[Od.EKFFb&ASPU1aZ.V9X(UGF,#&d03
gO\I8NS(Vf7;AL5XWK=IDg57b7S<#V=AP#K^8&]:Ff-508#[dNB5]fBC^=35WR,9
:>AU4UYJ>a^H(@XUPZG_GDH^4RV,P.H2b<<1)LG24]X(91<5fJP)JO77JU\C@eK\
-a<L:1=5,2R^:R9#2b9&/IgBdI1;.Ja/9N.]87XV<-H;B-eA)/4SL,/e^N/[-IGK
(aZE;@69b8T44XU]-UIWQ\RPVD41AcbQJV7Q1K[OV,E_V:58:X&+IK27,ec0DDC0
&aC[A(IS6<]2+S(V4U#gd;&S,<(4.QU)@M6[9?1eDT03[AJ1.GB+2cD:VA5F-_&V
CWX1Q]6?#37&7/e8VJ1PdEE&9_+^U#fD1C:U#b<+EMNd?#)e\VQa8R\VK4)OL1L<
[3#6K\);f,f\(Jc/G?HR1]L&]]JH_/K>5FGLQSNN3DP0W+(=_9]ecc\W3Q#9>3YS
#2C_.Z&gA^DAT,UdbR@#V_J0,8,D,W7f-Q,4+dHGbW3A@aCCZe3>ABS0BEWg<<Kg
fOV;/-?(bC-<Fa:N]]aVfMSAOOZDa-D[7f4(.I,<aK-D--<O)/c38NIP+(],+LSC
4(;SZ/@V=KBFdJ@M]fJ04+?U+5dEH7gcbSZ<;\7)=SZZ/YeXR[7SQH,3[O5U]A9<
8Uc/MC9@Wg/O4W&GAOa.A7(OR,DWG/aWS<dgPa])3X:CC&dVWTA^QgWWbZVYT3L5
SRTdV,A[d/[P#)]Z&69R5JE60V9gd-6@AT(&ZQ8G(5P3[GV,)II/CHT?eB_TY\A:
I<NOF2U]&Q+RG(XCDg(#64)@3T8EF^=JdbJ2?E0aI):(>(:J68E47LNE#Q8E2CO3
];;4AFBZH)KCS20K;AX5&cX^cc+g[1T)XJ0/RbAD)D(?;E4WGZ5E_J?_I#M+,?#Z
c^=-B-[M3J_.QA(<=[6@cM=.2fI=f(=W>UB&USC0LTVfd>c]I6/V2Qf=\6,)/).I
@(47JM?Td(HNHTFFB?^a90LK<T<AY=X1aCZaA:0fT:=(X.gQaQ,J7W&fAOI0Z);)
)8Z1cQJLW6RK(S#Z6)LP)4)XO+We1B(E;dNX5\FZ+;fLZ:>PPTJ&T.UJ;IgRA609
S-&MC,<EeU3V.f6CGVfM4KN1RQ=:BV&O5&MZd-f>6f4GZI;^NAICITS2F4ZK9YO[
VRaMTA6J8e\g(BV1_&Y(GVLIa-+X)Cdc&Q&TI<Pfc;>e]dV4P6IIY2(,O&SX:cbM
a?P53&&egFCX)]e5>_3SH-d3D(DX/:?CX@6B1]L,_/gUJQd:>XU_5_#A#:5A>I4W
H\XMY^JM/]A:fCe3D^Z^EOK00M0)=)_P]TB)/?0]01PZBac<4D.AYV[\gg/Abc/f
67PLF6&Q(<D]388QY7Q9EM12D@ac-c+2/IFKTWP(T)Kb_ab]c=7-G7=?U\Hd6:E.
M-5B+/Q^I9aLbeM)ZK.OS+eN<2Z@5^S/0a8;gKG]46<<Q:[[aH+R7SdNVTY,bQZa
8feAW&bU>e>RCJL&_0=+5]bBScNaL.@<XDLDJFHCfS^=E&[Ya7TS<=WHJ3,Y_9^0
\Y:d5bf=<L\>KWB6T8_O_cfc#U7AEc\RGK=7+-0T&+adA<+-QYe\.8EG7:)SB7)d
GJ\cPA0DNW8S-eDWbFCL&31a/c-MAgRJVFWKHK,bIZ[]+W<&SA8/?IRWWZ^Af+)T
OIe\<DC<9?OFF:IXHOV:M0K&cc(=S:QL/6=XV>]?SEg>L6Sb:+U&bg^e#>(:)>PQ
CH<4ZFXI@6/Y>(cFWIOL@=AB^7@IPdg7YK2(?Re:K[D\S6^fgN)b[LfQ)Q3-4/7K
ZLH44W1XUfJ?.\XcGPFcIIN998\cNR(\ggUdeEC.-Y9L.6JX1K@?\[[e:/Kg8UI[
eGK>69E/[F<M]#\)T)+1R&/H&==6/1L1g4:aOS7)ZO(=/?OY&J7^UT24V4.T&O_H
dC(I@,aD&@g4GfeYNPBEG]Y+/4[0g/K=Wf+1ZP0D^[_\a(?N;O&#PMM/XbIT+FI&
P33OEDUe@cA.Y,.feaXVE>RT2>GZ=7.T0Y1;fd+R0bGY0?]AV.7@M&:9FWZM.Yd3
,7)C>.]J-,SV(M.#2/#@82Y,V@DbO<2ddc,QTe882_^,_Z>E32\3JbLP[IY-]W@3
Mdf:VE;>MI6A@I6;)2N=fdLSD4ED(F9DLSY.;cZDIe7G?U[BI7PRD\&N^;GaUK4K
,Z=I-\/@KJ-)/eI=HA)J5+DJ;Cf-8W=B7#PeO4cG];2<9?,BP/QaL2X83I+6\WJ<
W7-f4&cT&H/L<ce245b#<:)_R\6d(\O3_[6M\IW0OCLP.^31E\_^.eaGWd\f(bf(
@SJ.P3^A8LeLCQ:6+V7\cQA;JJU9.5A8;69R]F8[Q-G6O9H\>[H)AZRR;1dK+B^N
S(]W06FQ&25Tbc<(_4c-ZKJea;W7>b4C@:=+ZPTCDHI\^>cA]Lb2a/Tfb2#C@EZ4
0f+aPT>J/XD=Cbg1>EH\0M/b5J?@b.KDYPY)FGXFSH^D>0#0)4d04gWOSTP^P^dN
FF@G-0eL^?KIXKR0V85_-;3f)dQ07^Q9(5/DA?VR,5b&YI_F@T-(fEV6Le\Adgd8
8YL;L0-T_9Y@<[9gbOQ7GPOV=YDH2bE5R:H,L2,b88O2W9?@-YVH=(eGSO/>:]/O
fW0BUEMbDeg):,_VVS:AHD]P.J@C+::=bdcC.LB8)Y6NL,WZ#,^0[7MR]KI)I+ab
H<@02?&7W+EJX)]K7=<7-(7=VB,@N=PG_@VYCLg,WE+LNNb&SN\(15D4S2b(W:Ub
CV3]QZG4Y2OT3de.,-@2^C#a38KU5&#W3+>+1bdEE/McY/(G/EC:MK/JfY@<K6OA
cYa-Da:9g\f,)M1_X0\?IZI]fG8_?SFT+.WT1L@LZ[G[UNgTM@H-X]:K1\0Vf9QO
,]A3AB(RO>?:0(JHG\0[b.^,e@LWJG;0CGU,+H3=Z<NA,RO-0USIR;OZVX-AH4b)
)^Bd6AL:H-?=+c&M]aX<+WH]#G.F5V]RA6G#A7R/1W-dN8(IALK_4GGTW@#d#\0_
FC\2DXWaUbD7K)&f+Kd=AJ&^g3ITJQXf0#[G2W_+G82d<TA@aCaCJ#P&Y6-G.>gZ
f7(>OHAR^+K^-[(3@.?/c489WU>)&7L_RB61Y(eX/_^SN;5JFF=]TS.W_a\=fR3(
KMgX#f44ITV:2#eTER]bDTYC4gB/]&@g+Fa?_Kb1[P0VSB#fCV9Ua5H;dg_@IS9Y
,\4Z+JN\^(?GW9/2f<61V#b]3:B(Vc_Ca#[Y@\<=,aYE@fP>0NX?OR<YB)1bCVW^
Q\3/=f=>=)A+6;]5#KZf[8aW96D=^b9=/?LdUN<P92QX@=Lg79CEPKE4?UD):B=H
7RW6Y<8BB,16f<TU-;BF3<@JCag5bf#C\.)-ZZE9KTRJQ^:UL/8\H,2O0gP1OU0,
J;]/cA=.dHD6K^2NR),U9+I;XD/4A:,CJ_C37Gb#&G@][+S2+16S7fL_\2f.CD5C
Y4HRb]ALTGE-8E=_(M(QM@78M&4X+242(af.5^f<TI#>L6KOEK_7\B2L7Jda#4b)
UYZ<6J@9DS\JT8BOH&L:[f^H1(0]#E0)@O\TFIgL[aD(d6:P5A[:H(G6WOe75F7S
EEJ35?_A0=Y?1cX/)^7/-CEV=IYC7_5\2f<F\45ZYAdF]_Le]?Wa9,SK5SP;.a0,
^TR+?+6DcP].YUcVBA&1:SIF:Ce?#a]@?9a6bd\9,MCe4^(dHB]P^Q+/+FW\1/MF
@:<F=K[AbXX_^ee#3gCT^GCB?d1QT1\TXgEb[U,8F6d+O1dc]H.Nf-W3X,C=@=]9
#6dPYNX)<NJ/I?8IKJDU.O6?Cb)#aeQ)..7LDAT:H/fa9MGX_P<.X#Ed6F;7997f
X,1+)I/H(IH_[c:[[:(ZAO]P5AMX\f_4MS[&U3)HBgNb8AVHSPVD9B9]eLK6Z(]+
(R<dW+eXVRSF<U_51Q^JDJT@O/I&G3GK@A-.HE4V#15BgdLFUCe>LG]\Q;W8Q:X]
(2:OB;1e8X.cK2W+)A;AA^ce(>ge?_G:@YT2\INJI5_>G-_OSMD,HMBN1:D3IGb@
7P?b^MQ6)MV4Tg3@++12ffM^abae_L]#<cUdC._4P]e/<H^.3EdI2&[#UB_fQBMe
cS:Z[@7PTUH8.F3b<aK,-7TD2Y=;+/Y<^&dC<88.1]TY@1fLe+)d99,_NT>GZ\_C
c.\AfOQO[g:B5_A6O8E?<:\bP9fQLY>+?g^3Y5LU@eN@DT2]8Kc_D/Q\&V3//D(H
&\6CNO7W?O[OUcO9Ff1<bS[/#KQ<E/\^]T#<BaU-7ge0Y[9\KCU?U,-;2Q9-;YD6
1K9IU3Q6]SI+d,Ud;8#f@1T,/L/_;J@T[,C;#]VU=dV4N@7S,I8L<0]V[fQX#0c4
<INN>BEH3;d.?@JMLg)Hdd#M&2JHPAO5#a\Qb#A8DS<K&Gb8Qd3c+eD]TaEYHU1(
ZGD^Z3(U,?.TDH+_.JAI-@1<,2bS@8IV\B^(DDc,(1Y6XSTTC5d^+88aN:+2a105
T@;<6+N>#_W+@Qd.A5[d8[K/OP1eA-@P154:@CFK]/=d@daQ,RDPQD<eX_S4\Y(7
gAH3FcfBS,2e-W054D5]5U(,8[#,VCJOaAVbB6FB4dH[2\DKcO(aVH(C_RI7S2X/
FDK^P#6A4U.^\ad+BNaV99Xd/e0aS[/(+<X#]55ULU0@_95(<6S4fEf9;-)41V;b
A-&@@7a2D9SU>GU:9LV:N>)[f3VA0O?GbIOPDBQHTPC:c0,SCXMZe?f^Y48a3E[b
LA\6CdBC4\)L)Za]Z4^?];dN-8HYWZ8=55e^BNB>Q@aJ=#:O0@Q6bMd2QL\.):/f
E&]5@&D[+-DN)R=<UPMZ_HbcTQ)7W4DB5.72WBfZ/0TE)J>]80eZK3?G>SA1V?=2
fO=<B769<\SEd>W[#bXeE=JMKJQ^aL7@],6QO<8I4b#=ZUJ=EX.9f(209SEK@<GU
+\G_+>)-DAMX:Cf[[JX90.W_;QfcWIT.\W)U4>?>b>RHcMW#CD1+S=?<I(>EP876
MQA1DQA+Y]SRO&Ng6AM8I(7B8K=^>@HO)6+Y#Sc6?#^QF]O\S]M&BQd9cJEL+3?-
DcX@Y\\^aD(?@a8)@X4g=0,8R(NG=S5WB1WbL-QQ(L-KTXZ6J2(][HF#a9&2@S&<
aIN4C@VYV?6\?6L-[(_AX)RKNK>ETbZK(SIA:5_:b=UQ/W)REQRZ/b+\U?I?RA7\
bOdb@)[IXBa:OKQL8e(]>S<5.L]_#b01;_)8>GMYK@D6U&,ggKYPG@fFcPA3S.D&
c[^Qc07f=NIH>3NA]T#_TMbC+GYM=/I6-A,BCTQXFA^<Y\4J1LJUNd9<g;VdH>X?
CC>]c/b@:2B&-N63.&4VV7^VgLJeV)YM/9603>_IHL5cB)3aIG0)YXbR[4Ud\QK@
;cX7Q_5KGXHDN9DFLM9R+B(105T2&IMcM?D2WE30);SXO8P/Y?-2MZM@TDI,<Fb1
IBA>1HBW+CU5g;75=<.48@21f=\88UKAfKG?0g.?<<AJ?].BQ.TO8L8Ab9I0G-VJ
V(FCSGUc;fYaXG9DCcX/L4GNcJN]a<A4ALST&<82G(47CSTg:6M<+:63gS,^_2b&
cD(]K2Y&0<:-\/Bg8ZER#[KaVb<;#IM2eQMOU;.Y?0RCT\DX<U]=8U@J]Hc5Pa&b
VD2aX^XCK\gKJZ)<KHW-=]@@,C_,[#4R5KUg)?1XZ,g0Lf^ISF)e>.BZXI6X&J<<
INQE05MR;?8b>XeX:-Ybb?3(Hd3,Oe6&NX;SA#\K]cMd?EFA@#ZLbS@Ec[Rc=,\6
G(>4TgQ9&_4@PF(bg?.;Z9+WOZQ#<af,a9U6ABUA]8;LRf1/B=;C9b&;A4ZYBY+a
FG6BNb0>Z(,:U89><&RPQ4]WP&V,fJ.X.>I>b8DDU:P2O@8_O]g88W;,XDcU=&[G
_A3I94.@C=:DF]-HTJD4g)[3#9#7+P:g[F,VJS82\>D-I&(U2_+C4E[1;d7c2+44
/f\_g_Yd:Ue#&f-\MNH-Y58@)Z9EC;5Ea[&I\7+c\V-T0.;RXMd2,.9X7K0]fF+)
fb0c_dV;5#VRZ.,XQS_9+8PUA:(+,#-YQNWEfcC:O.d&LLG\B039;d3R#VRd#>U3
FQXa6Yg/2N9LaO7L<_\Cb=8I?&A@?4EgO_^N#Zg&I9,NKObe_U=\@;8\QU)]?_bJ
cfd.5ID:g<7VJAeG@0<V_MQGa8ZeDP;aWY,9:-1EG:fG/\KI)P/<,;_)eFVSVcVd
ae#caAaNVL7Z50R/SP1H\?R3.fXaWU\aK>8IP1LK@5&b(dJfQbb,Y4UN3H\((W^4
(CQ5;#8N6?eY#;]EbQc]&[V<Jf>LOK^?II80N??EUS[A)D31/gOVfG4eaIT><]((
#bCM00U,#Zc)_1QaEA]B,b:C6U\YP@);N(aG0JOBP&28[I^,FY5.dd?c-,+TH^Q6
^dC.)P1=9Aag?5e#9Ye2cIW/#TB[J3V.;FcLJ2BQGb^+65GF99VDe^2L2K7[6L<1
M-&9dfag@_gH/DV/g,L>cLZ.@^.=e9,1W.8RAT[;51H;@@2Eg5;f5N,LCZY2M0JJ
=07/1+Q+@0D/D8LWgF(QNJ,YB_9aY5b@SB#J:&bHC7:c(fT:?O]\C#VeeO=@U\SN
GPNgOge8g+a2Q\/F,H(E7LSE1Og:&R>C,SYBMSG>@RdWSYG&5(6(GD,D1Tf)bacW
6fW_+S)eE>ABV.)@&A@9EO@I,]1P]HE&RQC.6,Ob>.C3@B=gB+(:..EZWF5NGAE>
:/@0TWC:+=fJT/ZOJEeO.IHVW-d2^bHZR8YR;Ge;e7W=;aZTHQH#O1\X2TO5XdZa
FQ.7d6KY6YSJ,-.PUA&\@T;;AP7Z[X6/@/W3=)8FeO>,NJ9.--+02]QUAdHXU+&J
c#3=EQE/,&.+F7T(EJ&TX?d18S_3c#2SRQV5,-MI<Dg;XQ(#^6gJfJMgV1S]0T,?
bL2V-(<]?-aXGae-5g2EYa2[4[QHR+Le:5A(b7:,:f>3AP-RT7BNEL0GED<]DO39
Eb,?H7aHKHd/cbYS\=U<6+G3KT@IL8[K-@S_]d4S0eg6aT,fAO:MSL9U^L6X8PcA
.b@NPKa+_&B&bcFXN1FJP&Kf1cKd9M-bFS:1Y^^O4)YO+4?86ZG?gD=(A7HYLVKO
BK8F3SLfa705O-Z]9c[I2VFTd+W1VQ@gGCCXb0<(_^FGL09(3]f@g@=PAMF01L4^
9598AG71VAU?1/P)WBQL,J7eI>?0Q&SEEdKcG@(\4dL+&-Y2@E3=V.5\UG))(;IB
6YJf7=+],<>8VJAA.\6HFEMOH#^DcW,5;c@\HV\X5d3,GdC(+^MTTXKaQ;RD:?Z4
WdMaEV(86M,;],AUIQT6\Z7#-U)G[9cNVV=SQ:)78:/7A3-DI(FM=G1Lad;.ba>H
M_JMW>.<L/TWTR(1VJ=\[J])XHKeAcPSX:=8I66\c<Z&9-]7^=7U3_P#-K<V&7WP
W:SbV^1T1R-ZDDO9MV<Q;De1R6XT?(V/B(CfXa6WWDK6gbIU5Y4C5#a1C;d&B=:]
BN>2J@EALX:8M,SDE2_.4\YXFeFa109]e=VdBe8PL9RKZ)M/I0YC9+]_,X4:JK7?
N921Y8-[EG58>,0[[4YA,&8CD-K]Z<_]@TO8TG;4XRdO^6KIP&=J^2N5Qc?L.X).
L@GCAWMS.5;BMX9,:/O/R4<]Y/+S@cKTD:0S:-?eN/<V<V;?4Z_HVB&=fdgB&;X\
/\<.VHa&eAeLaWHf<&BK_Vd60f.()PQ<MfN@S4=L4L3,OWBOOFeMOPTg+K)7-490
HdD(TD[Y;35eV)B92a:J]NWUJ@/7.@c]29-C9@/7E>+W)H^#5OR@_b2_CM;O)P-(
VW2-@9_F<G:U<M9E)X1UBC,&PN=;bG<ZZR5a@gaAf:35B+LQ/Z)TEU;/8CYgKMH1
-A=_)8\6<@+C&1e(cDY@_]H9()Ub+,B^0#ST>X6TeGdBH1Z5?0G37?6Z2Pg9J;A\
A62DGCZS4/0cS1+-ca(@>.QC^RKNIRa<JT)Q[f(H:dC]J[LJ\:H3=Ngg6]X>#[:J
#CdN]N/e35<<=NMT[POOTeO-=UL.@.ER8eTd2G0]PDISgPd^K<[cC]?VP=Q=(QWS
d+WN=/H/f#Y]_4-QO,)U.)G)VZN_AAUY&0<1CBaBEU?E)DD.N+8a1QSZN#(JT;99
VD4BUe8Xga_CO(F[(aE:a0ILfg6U=BFUXa4>ad0W15PQEe49/I&f1T)M07VL3A,E
@2f.?+T.Tb2:<_[ADS3#bU:g^0&[)b2#e\)]\G^8Q#dKX24f0OV3[B+ER:-#OcR=
-95bXX@+TOCSPV;daI@&d-N[\@3VUKNI^X1^8ONg;+TK#cRD/B8bURF&2X@F-c)c
F-_@4MH:fO268UU1SG3&d+8P>(4/da1HTD@0RRB)&JJ#cBd5E[c8>e+e_:aXI/W4
3VC.N42-/>IDHacB2#/IJ+fIP9<^GF/d&]H+cH]><f>?AIVdPgNE,C-ESO9bD>&H
R.G8\RA@bWf#29TQGb6[987_I12DY<fJ(Z^PadXf0cW]M&e\e4\QWOLTD><FZe[B
-+&9ff80J9Q4,\7(M>8\M6&N4D]JE(f2/ZX26<38VP(X26.Ug)((D][DPO4g\f>F
/XX95BaZ3Q^ADCG9d#;dSU2.#4(;0V].BX)b4_5T76:+B98@RGR+CfMG[[DRf?B>
T]b?^,^;))PUd?=C_OO(RMQH<dJX216BMQ,FM#X,)U>\ZWHTa<\8#W[/FIYcP]8Q
CHAGG3,58/U;cfJ5dQQcdP.EeX)]Ce6C0[)O6G0aQN^@V:B1JF-?8MV64gY.8JJ6
.2=@2Q1bPgAY3.E9cQCI_-^Zb/;NF+?NK=@T45U1^[:1)Ndc2QXCdd:5J&PGb5BR
<-U/+9/7,UYbEJaF.NUV]BQ0FU?L;_cBQ[LPX5@daH=XB_DXf@G]]BFS(gg:db[F
;U1=JX9B)DdC#&NKec8a->/aXQ/VQU[(b;1HMgZXH__B-T+VgEO5B;If6PL[fW#<
+/Q1g^+-,15[K+O5WDBTM.2Q_=cKN64W[8P^U63DF;\W2BRf4f)AVd9XRV&4ZgAT
M#R^-[P4T^B:3+7&^>?+S>?:1MKN<UR<;ODIA<3CRJB-JWT)P[RA@gGP9aM]Zf?a
UA6bAG7IJL)+/;9f1BOaX31R5g296C/;(X<7eXf76LXBd)W(N(P4U+-6/;,3.c;c
(gKJA015QdL;(T6T@U05&K;BO#/G1L=^_)cJPA_O&)BQ>5M]Y6)__?(MVX<,@4Yb
S8/6ALOFMd8N,FQ7ZHeEGDA>>[fN7]Y<b@Y6);e^A/D4QD<Z@W6)WZ_WG9RA2gB5
&20Id/G06f>UUQS1?@HeW]3d2T4Q604:Q3dOfLN?>cEA/&C]dGCHNA/^,WZSH5ID
57MZeVIHYHa1_C]P@J#d;;OG?eDIZT))7_=7VK9L:H,c4BML;T.P_<EeQ@\LaIR\
XJFe:F[\4K<Y4C?TS@G^D;Tb[PWU]:,cd/R\>Tc.30a\2#BH)4MK<#?344O@.U81
0+ZT;R1((F7QQ,;WBd\[[]Sd=.91>5PCV-?>5,HI[<59&gGH[O8A#469(e7=;;.W
+CJM#Je2R/X,\5P9Z>T2++GISSgN#.V[1gJHaLd=RIBBce94W]+)]BY-B1ZLGK&H
14)8B-<2W2I,WYKQA?9\]/DTb/JRF7U)@)K<YUgR2+;O-VR4G8]_3dM4@HDF@[(O
:+GE7#^8Wc8#]:4N#[_<D?=@W<CQ^S/-^dF9,8e;N,F2f&#80Ef@U;(NgF07TKTD
=1M<XF\_;U)0e<(^-;]6.;PgV2Y(&<&L3fP.2\B:)#c1bQg1g)46>#QSRS[/A:B;
T5P40]=8dZSAN.BP2JTNPdId1F]08IV?^dP?F#HG3)CMd9YXAdCK85#8#R]?\f[S
W)4@5U]H7@8CV7>Y]-7JeTW9GUgaB308I74.AF,KB.CS@P=0,]3Gg2C=UM1X7H?g
:V?__2[^RYR\5J5=/1V=cVJB]\W_69?]ARX_c/,-_GL,T3NMg(17[8ZQ@..EQ:Z#
L>?4IWRd?VIHEJ&KD=<H>R+B#X[FGg?1.Ya/1A^GD9A40=<e@.(P&eSG/3>,27O[
)acMX51B05gKPK7,Web6FSWVRZ7NEE_G5RE7\/WaUEUBX(>=8?0?N4/\W.40#6Fb
ZL\D4LH]<V6=>75;5+(aYT?#g:Y.;ABEcW@L[4@gQe]Xg7@((G6XMWG/]3&9gf8Z
9[)71<_FF_&K67T\6,aFOBf[DG&_A/1R?J/WK@KT;(A)+C>e3MP#-H3XV</#C,LY
[f^VLgU6NB-RK4.#XH/Ce__#Yc<AaS5I+OX)[HEY#/[&W5Q97U-aGF,c_[gZBOON
_OP(;6gIcBI+M,DO+2R>QV>?VR1gH[gABH9+^I@JI)Z&ZFC;V0CA-:]6Od/G9=0I
3[;C)2MJUaYTXUW8c\]TKGE03dI4c^KOART];3d?BGAf(.2PDDbfAOae<]<S)GVb
P,Z^KF])4BY8Rd60XZ(/Q23@^Jc@GD59IXP]N:(J-,ASSeO-H>1<?M[QgCAN\?aN
TQ3+._gQ_(-+9d.B+QK4JL7GRH=L5WSF)ZETZ^33/ZN?(Y7U+2^:I0aNB0H)Eb<V
dDb\XdPdY_EfJQ00)F1]aZ^V6/.MFV<f<03D:Q3NAW:cBGLeU=Ef7)/Q04&L_\HD
<N3g6)f>6^a[#_GWG,F0BEC<Y371B?6XC6\#?VbbO8^HJ4.;TNJW)P.#[N/:=\4V
c9@:?]<,V.P(b2EFa4d#d,A#]^RNF9(<9aC\OS9FeBA&ADR38XN\D^8@Ba(a77C;
#>M<aT^eZ@N[2^>ZJ2J5fNgI0D@IcI[@=W=^3YObb9)R[6C;7)Gg2e[PEA[3B^/Y
Zd_X984Jg3TM9T;=FBOBQ_2&MP:=8R>Kg30C(OJJcU[)A7YB44Wf(g8\-C+X-GDM
0@?HB@f1ZABN9D&L4M:?MaVHOcWdPO8O1[+=O<<2?5M9559JCYd(gV,\fF/)H9fN
/d1Ada=GTA;.7;Q?eRV-6g9.2a,aMQ>]Bg[6/U:WC95@XCR:68BOTA7]Rc/Q6FSP
IBVRB@[0086fDKRGVe]H7f3[b_0JTJ(X.;+=4Y//M3F]B=b1XPQE#L1(J(f&()[@
SN_.7,_4[c6-<_X6T\G>geK/:-#V/NNcNFKQH=)8bF),&N,])JV[,bX0MGUU(<+K
dL9J6\:c9[;SYGOfRb?f1?7,IaY6eFMJE/Z<ICDEZHDBcCFHOX_71&#WI#+g[3QQ
WJ<0[_)YL(V&GgDRF,T-)98,8D8S)[,#EH]P?M@<3F?R.4E1AGV\Q8af,HF6;]EL
;/+d/Ja8NG>VE#SdGP4XO9)U\VXffO0(J&KFO4O/NAe54Q,J/^:K]2J\PUJ,C(9B
10WMG=]f]V7;?9c/^<J7d96ZIC12=TVV<Q1^6D)4G&N?&#]0^,Cg4:##eBJ:5QdL
4OAfeR5.U[La=cJ)JMUfgN_OZ1?,:\GK&V455DDH_R^J5;N&B6ff,Q]8AW;TLe/9
8e[=_1L:8_5NT=EgR3\)4Q[7116b:0g8OX1[N5P&1JAZ>a1F;<Jf8L1,-8=6\VaF
Q(-:&V^fg<g+BYd>Q:&.SJX:)8[2^\B\->^]UG/<A;:N^P0&(?T@)/[.E65+,f[B
:;I(=7OXaE,#2XXe#]34Vb,cX)2]UBe;4UI.f;@9ed8D?SEb+>#:Y;OO<EVY#-JE
.33DaLFQBL3SA#(8][1d:b[PUc]->Md[8^9#BI[+V4>7AZ\eCP40:XU,)2]S\J64
R+<U6^B&WM?-1RCbPRD56fS3aDU[<NYbOE],>TAW,g4#D9B-_+8940+eT+2NAa&-
7:9d^7..1F<SITEG\>eR-?VeX;R>5S3d,=;A2<?4FK5AWFT/]HE=<]L4DXGeL8(+
Q^H:TeUO[D5SO1A]=)fQPT1369afXbW4J#L0++XOf_FOQR/^PXI^_3<^N&1O6/=4
_AW=LVU/bTTdU2Q12(6W@)RI/K)=L3632NN7I\27/=\fcR69X8<CRJf<25_5TgbW
M.#E)\/Z(85=7P8RB_>[.=eaBLSOZ-IABAA4>.GKSHd<+U5;(AQG@A4O83/S>,67
0?:9[_FNAP=2Mg1^\g?^^QOTPMU1[I\PA)/N@1S6./a6^9f(CfH,H-@R^5]D#2?3
6S+4]I_V]aI.6B.UaFQ.8B.KK#4;R4c33WGa^d2M@STY+c7&T[7fX#738N2FEVFY
_D>KE#IM7.VFRe=UE#&X#NEaXOZ1d?O)MIR.8?5MWB5eE[A;K?[W?feIUX_)Bb-1
JS+/(F=-M-=<694gJ&\T??=d.7QM:I+37_R-:C[/LE7P,FP^a@H<:>gB[dV\#+=K
NR4U]>[:;ZcgP:=:>PP^GZRQ:EJ5-P@RH(Z8Y2TI8PT[KO9P#UG&:OSU#+DIfUaG
1DW(.=EV1)T@<c6+^@=L:D]P\#cUB..A?/WZJ(<XJe#fK/V+1L5.LZ-6OGP0eD?.
XUG(CG>D7ZPFb&AWf])C,JE:+4JU2g9Q)@OU(ePL(?8-RGZ[2L^G_=4<6gK0d;UI
fCB:8gIMLZ?95LeXJB.dX#&I7&K@DZ8aXg[#E8LF.YXUC\4L42V(^K_7g>IQ?G9:
S63fMc#aN4INdO[/NeL_:b8R;W4GVL8O5D=E7g0cO?.X;2)1M=AcQNAGb5E02EFE
&.)Y71HUD&C\YKV60dfIQbb8[@B/L/WDO+)XIR40?Pc[96b=cPLW5Ff?TQB#9/T0
7]1>51/0VYKND<3.,:;E^M-N5gE\X])-:PdZ7b^^&_Q,?Rf[Ife,g(5Z[Z5Q#YN1
.KP0&Fg>28D\aXM>(cTT9K^97Y?Y6e&JU]<:)aQK=,8+S;\Y,;Bd&ET.1JgOJ;S&
9^@aSG[O+@?G@Q;DQ,IDBbJYAeOLGcO@6H<VE>Y)fOI-gIZI,ED?V_)E^LadCFdV
@WF?]J(#V6DW#CS@c8QK^H)W,,SI#Ke9MEfdgUHA-/QDVE8^RC123_.)@g/^f&?f
YUT[\Q=U1DNSM0Q:G08#HY>)/N(:)1Fg/^WG/EUa:2@Ub,gCS4C>6N\N_6\b_1JH
69_@F]S4-VP]<Z2+aS)OYW6eZ]\c11P5=7#4d<=[B1UN.GS823C3A,A7?LO9)HYC
M\a8:Y.^[W1,V(dSQ]GDQ8?U0-Efe8OETVM;.<D95AI>MK?6H0Y51Z]>W5CH#O<<
<V(.?abba1fBR#]#SPIKdVCE]UHGXB[\K+3J5+1^PF:=Z;?cQ=8Tc;B51QMAT,d,
+NO,C4IW]MAPP\_+5O:_O>c=9K2RC[EDORN^NA4GadQ,@G+Mf8BXc7O\K0@5=JO\
O73(Q^P^9P1\d;7X7?W7&O,#GLRg3ATN2?NJ0SC:)a/.1Y(eQF0UEL24^-[0HYB6
WJ?a[d(Y\9cd[Ac659dI)(-&86J?_XX?[MZ[:@EHN>44f58Be++N4U<):ZaeI;7f
FS7HC3-F6O4;FaZ7]aeHX^&=QEc_&/VgIWDf[?SUK/a>A=]YT8+M7C_UIG(MU3[a
ZO85ZXgWIQD>OdBRCUF<K)MO,<32FgT</:S6X8?AW1NI;S@bcZ7S_JP_a<UN[\N-
c1);1F[;f;dM6&6?TL#+PC#HeSY,K_\/J8Y7<U[>H<<71MKXJ<\UMFNDH>D&+9AC
g[O7REA.HaDL-Mc?-?\YeKQ>[U],W48)_ANQN4XGO?IWJ+_J@)4T</)EB4<S+6)?
(IK#[+8FK2S1bPJV)8_Ae./(=4+=1]K,L4f#E:G,7>IS7S=?1HaEH9^I2E=/FE-+
,;I-0KJEHP.]#Ef)KH6NT()4WBURMI[af()_.;/^6+M=M0(a[&_BcU@geASC5,ME
Q6]74-bN9++MW;,Z:N=gAPZa.]gMNVBdac1=#)a(9D]5g-I&;KM&NYLb@P+].89M
(TT)F?DG#.-b14^RPUE=Bd>X6eSPR>;:3<\WI4&D<LID\QCEIAG4<b7S9@bF5bLB
/\@)e5I&1:RFC&GQK#CZC1)ZEUg?F^WLfTe8^8B[W45Q:PBRZRdI12M<XGbJ9)2O
CIf3YE/^DIC2(<.U\(GL:Ff0?d-XYIETWa@cB6N,BIcGK:&IHDA(CP@FB0?W91+5
LPeUY<gc&gPV(Ie(?L^Ce/5)R&LA@aMCD?(TRd(NabaK6\&D(?(__e>7P1CF1KA4
>B6E.Q5Y625H<2)_>P=RNR2=DFXK#Y()J:2^Y[>&+dQ3]VdG9<-I&36OWI.MJA[^
O>G)>fD^eDZ<0MAM=^6fR37UU;&?+.M=SXF.Q#7OGP3WQ;[61/\+^@OC]&3JZPGI
\Rb3#64<RU3E9Z6JG05((R&KLO(,67A#J4c1#5XB<ZUNCN9GPgd-+@99M36RUJLK
#HQ]NY/c;,=]2YJ>DM?H1eOfgT7<gb1f2^AAQ2#+P^677-2bHBg1]IdfZCN?WL/,
SO8Z[]fM07)[]JW9&2;QF+T=H<Q7->7/]IHFQeb^KKD@PMJR6GVY8[3OTd4DbZ>B
5/(].(e99)6XGEGBL-601fQN7&F1Pa5,3M8I91T5-2W6-\EB0;-PL93;7_Gc]\.c
A0,L(K#>]9]U;+S)8N5NJ9T(KXBI2YO\^-#LF8^7Qb:X7TB;#/@QLCN5)>31I^PX
R4&Y>8>W+cW?1SdG+LL4OGe3&c^)-LV:de/[2JAGM)N837JZ#dH^6:/2(K^_Bc[d
,#/(H#JW?M]\199cB:cM=gMKf(K7?Z8ADX91g=UO[1[YgCF2<9cWP/;Ac68Wf>;\
eW00SDDI[HTZ+E8FACTb:DYR#JWb:(3\X8&<2)DD)(PAW[(fW.D\:.X8RAcT107B
BGRVA1?=F]CSB:=<#2g/a_WV3C^DNWR^KJe)(</P(Z-M]eU=^\^9D(2TW1ZR#[F:
e1V8,-6V[@)RHU[RXR]Q=bcF_W&+GEbbQg]F#1YDI-Q>_bO:X[e;VSa.9Q<H)R#F
08\)Q)(2#EN&60YL_CMZX]Be+SX:8MX;@-V\)Q+3V(?L?84X7;[Z:b-)7[X)&>Q9
IM?IW.CaK9FTG[,]4[T2bW2SC]_21cV[L51)BW0L^fSS&[+NR?SN)PM.6#B#J#Z:
gZAHXDb.>()Zdb>]_[KY&WO#JU&_P^9_2,O;<W[3.<-eYb<DbC2Od#?cFYfFL;f9
L4gGP3BXS>c+X/5TK,=:2IF?FC42b?R(?^O3MGC,\?QM-_Gd==99:Zd6AG6;OUcf
N3WP>71C/?gF6U+5VR;[7FLY<SJeJ^0YMQ1SMc;)b,/8b?>?4Y+EeR@\?VV0SMD,
/</A,3\+7:J(T+ZcX\f<O29#/8GbKfd/DM6_d2bI6)9gV\cA=3=cJ]g[\^TPE/=L
QGCbL\NE@aWZBO^7V/F;CK#7(c?8+SGdNBL9QQIC^WfKe06J]RVX\EbOR26^[@H)
C22)@&HU4\/T<eQdfL_B\dYgKJ#VLd[\T(3M]QV@\^-0OU>TQTS8+JER1027IF##
2C@D8JRND6QA+cXR7):3KTNTNS.]<+:OJ_D<dPULgR9IRL>1UNAO\)gKU5A#U1Fb
#(MO[g)((OC@K6bG>:e=fbRD#YD>;5HT4a3c^8NddgXH7&8YDJ7bI4>^Jb=6:,2>
M=CGf+XCX6YP4+?2N65d<d:O]0KV6_1/]5K+NU_U2=^DO>=f76_A@6e4Z#1QYRC3
XFCddZ,(Z_Y(VScC#EL)0PZe-/JaHdWfXc7@)ER1J\B]X.Z&=XN9]4FB\QD,)\3&
8C/ZR4V-X4I:@<3H5NQ(7=(Ha^bGPe?F,5G],K/EULF[=\P)N7M<O.<VccDG+EJ<
gRIfBEJ5G9-Hd2eT3<Ne2U^^6E81GP.JE(g0G0D5?c4f)R0#&aaDFS-b<5,0)<)M
Z8a>;6@IONUEM#X2VSAK7^O+ANZ0=0?7ZNWfg7D;[#Mg9TLBbfKCB.3B[LeY[FYI
L^,D5SWI1YI6b[/]O.aFXc<&NF)a[RZIg&a(H;[X<DB8_J-f1ZFFSQ5aW##1=1AA
H=DJEg.b&V6aR5PcR7]#0Z(3=S6>B3T.^11#g#b&<+]eUdEaH?8MJf<.AK:AaP)(
<_IE+.N+;b#:L;#UD2#<c/(cGQ(CTFc:Aa+J^R<WGO7gf;A1H/OIYgfW;<1/E7fb
,>Ma+?0TF6f2VGCW4&H?.cJ)f--IBMP.RKD@EH(:GKfQ6FPP[U]b5X#g^?&&2P<@
g^70fZ.K<c_Y8XUG,+G1Pf>7QYfb-;&NC[\?],V)S0/UX@b<H(g_16\4[#X811b(
14g984#Zd^N.K(12JY?[d?,+&^RX1?=bGZQU9<VLNC9_9@Ke\;_\N_Y.G^_b&Af/
+YL6<2&^?Dc2Ac<.7cP]-SV=Rc7#b)NaD#N+aCAA[B\CfUAR,bWEY^&66&[4G)aB
RH-H9RbZe7H2K,4^AJH(;0JEJYBI8Jc1^OA,D&Yb+A>^),=?J;Pg:Ea7XWSOCA2T
FT6+D4d4^X6/>_@SXT0]K.21@AR9:f)=AEd,EF@?+PGE027Hf2CC.e:a@^+eJ:[/
UZ,.9UdT.eLPR]=9aV5\QEXJY/6Te]P;0_M?>QJ97&K7_-(>O;LEH;e(\LaXWFb;
>YQgS2AVW^c\VZQReSbKD-K283VUMDUWc,[CXGNI+LM5gcU0<_HSH<?He]HH;^-3
:(W&/N]_I@(7O83P^HUP9Y1<0RA?JEC<+Z>B3LXAgLUcZBW#Z<c(6T+6::d80MAI
.gE.JDR-8R7cWFW^KTE#P0TXVQYW,AS#:VH.@OdT;bgD#Q=?,/D>FJP?NB-5&H;S
@F(,H:GOIa7QXCMTZ#&Ka0cMBdV:0)bWXce@<P-R,e9_ac>:=&^7&0d0.M_PVfD/
>MC.:Ta6&HBGB)1A[RcKI^16X4\e&#_3W.^YBWTR_QK+@=29NVPL:a13?0:@..(N
P]f6I0b3KPfZEFROdK=fR9YE/+;#MNaNSM)6R>;LZSESA1^=L:]U9&]7cJf8&Q]4
TR0[d/<>SA?XT7B6[7PK3@R:M@J/DOLN^>BfZXOd5P);5RD+^[ZO46XAVCU<2K87
GJB2R(LSLUT,TO&1e4_QD(;2[=,A.]EZFX[2PPc9+P4<_\P)9AJ6cWRB-\[+g=c?
EI)-]&8bISe3eaK((295L=.7EH0NPH,Q@UFKMZZP](UQe/4\[JT#:9#5NdO(2SB3
QQG)\L18<U(^M^_5#0Yd6bT6fDJ?gJdC]LEZ(Pf)7,VFPES&Fc8._1]YQ-83([UZ
65fG3[fa@LC7E7#XYEASF,&I7C9[UW.N1SF8O_[MGXS#3-P[bOID39]60^</ENOc
MLH??aLDUIM6=7X8b(LaT?76<LTW0[:.,Q1\.2.9Eg<54\04>.VS@)62P9I@QM/G
&H@a?,Q_6TR.<Zf#_2V_59VST48VV/9,dF<@1AK.g_MfgH+>J-WcVA#)@VbA@32H
O74]KgTg#g1;TO[Jd,-D@;7S&-I5:bb8YR[]T])(H/^E:T84K02]DW^2L5DG][&B
4c41@6Le.S4Y)CB1-HQX3PW0Q=?-MLY:?RQ.CX_CBcW5,b>\#)9W,WP@+4DX1H+\
2a[2XETOcPe672XKgC=9DO:H7d:B5I[02f53[3.RdSafCDMeJC6W-Z\cP)QS(:EQ
4b<HgS^#+4Dd_-3&<e]M)RAS09H&1H.b#f6G2:G1=^VP\5D,(2==U.L4L+Jg>d(D
&H.+;:b.OGfR(CS:?[WLI^/,C@_KF/WS]XSMVP8@[@D^Pf(f-7,13CRK\OJg(5X&
HL/V(aFOOS3TQJB6V?c?-WXD)C+I@-G]a.DGaT[1GO.J/^WSOE&\KEL+V<[0AMbO
]eS7/+,1(KX6GLf.g:JO_ZMSW.d1+5d)dWfXRU^CEX+;8\f6ES930XHKOL#X&3:I
B76JBQ.F,/FWJBPWEJZd;5geLVXMXbX(EI&ZDY.B[P<OU&I2IS_9M,4&1:EM>MT)
9+5O/G7g(6)>/4W6K5E0ZJ#?VUXU0e4+IJdCCWfC/2D[R6R[4?D;:SJT#=&ARaT)
MaHfK@\.#30746<XI62X_)@JN[3Q7-M#4JIYC+T/Q;L(15,632L:R;VdBg:W?bD8
XD7>#.-L-YR&[VZILM@7TgGTc1(2YB]^8QW<XAO27Y7-I#P4+ZW(Y[HQ)MVI]BOP
c7?XL_WV;HMfcI2KGbIcGZ.UZc?Og)T:SH+K-H@aMR+&>fY^<K\8J0T;8T]Jb3/_
^A&[9MRTgEO__AR1RV2&.^3BKK;8a6<U>K-,PK]:+BNFY^0KbP:E[?TEc)]+dT\C
Z4S2aE1(_MAcQ=Ee4X4DD[FC6>4Eg[[RI#1)B/1.5A80@P8C?W#\M0S[=_5A[86T
F/aY61E_dY2#AYXV;8^TO1>UKNWZZV/):d:B/?dWXb/8@OMaf>0/&T99P\P(ILeE
=F3D.IedQPb@4;790#[5UTe6<5;-4.CMX@3DWF24B7\#[AVfaeR-@ZY-d28@JH^B
,6_U<C.aOD3e,aPaH4WY/9J(8X.[=2ELC1Q(;44S(3A:;_Q8]3R3)I<V2+@7E4a1
_#(XC_CT+COGW?P\C6S^/A#aW4IYeWNH1N?e#)QD#OEHTB3Ha>W);\\@NYObP3_D
?86X@P>.\(_MdLCA3&(.6;P[S0M3+;<Jgc-?ZT[?@S=;L-GB[([_gMHA9fIV>D1^
.E,e,0CP0PMcR40eEET:FFGL=N5Q>AAA^PHGU9RNL9=OgL;7P[:.,<<G>H-NV#Wd
<+IEN,^3H[DKS7Lb&#/.\H;-.4IPTJ5HGfWD^aZM[:4)Of]D+?NGO)^]_4J;d^8L
FZ?Q&F@NJ^@9fG,0bKB0?YSMS,<90CAFOdSMag>MB.16:eF-XeXW3F.T7=1F2T[>
4;Z+fD]9HcTEYaJEfZ=:e_8O(.Kga))NggQ+&TIO/Dd#<;OQP5<b,&LY)\aQD&Te
RcBb<[/U&a=2b[.&+AX_Ha&J=Y#;DH(b\U@YWVS-e0HIQW/&9_(GI&Z_//+7)a43
LTT&e\G75Zc\T)@(f&P?0#^c[g&+IA5W.V83(G>+0B/&Ya7,26JFFa7:fgM7?Jcf
@^NUDD>BOX_E564]L--BQ:g&[3/20Bg)W/4gN<^2T6KeaJW6456M;SKaY+6LP;3I
Pd/+US2H^B\CODM@Y(/-b.W>;=\]aG\5ER&b[HgP(ZOOQU5&,TJ;G?:MYQB.#7T4
P1&=#IFPfH1G5RRVL?\J/TcG.DP_TaOOXLM&=_X>N#V30=-QRL\R@&ea0>_44-9H
?aT8F>S\T]DF2Zc1^_#BQ+K=EU1L)IM:NKGI3]B7G&]5fF#6F64?II0:AUGL3U--
Q)Z9UNH,6Wb.,+^[e:;N&bO:-SL;SD#?:.]TUG,AEaeE4+KgY741+7E#-@VS0gIP
/GABJWT8&&FgXb-\0-><-)K&T^F]ODcJ>cZc460HM+0RNIXZ?1.<]]@A@:5YY0df
.P:?XEdFNYfAC\^0KG@M1YOGLH4eI2U7B(_V\aW#4\#U/NN;R4YOA9)CSE=4E;]E
R8ZEX;:2X&JD4.=8:56ODXG;)\#G.:WI=]dY2/\_W?B+FY-JZE)C.)b/N>\:AU]D
7HXZG5(N.:IU6]E;Z]\?(R;EW=Md=54aW&/BcBBOO,>4]G2KH6A9=3g&]NW5A,d^
^@NJRc;0V&dSB71OW4d(XA6F+R85.)6AL9\HPW8K6D8(5Hc@0Re0)[MSV(=@28@b
7I15<=5Ae<Y9.B9,4P#,O335/7(SZSE\_gRO@MVW-d4YTLc+3_b?f>9]X6EH?E]S
UO;U&M&,8>N7Hg+#)\/-;-Nf;.;]g)>58E46C]FbVMQdVK-\@#f(K.#T_@JbH6GE
-cc7K;VG@?,<-P1142AS<f9/<_/OKWX&2C5edB.B^1NCT-65S46\,ZW(:gL,eTP9
62^]LV3^_^@[b.S-2fX#+&^S4@F:N,Bf)b@Sb4/8ZE;I6TXI8?]Qc)dJCdU5.\_O
9Y5M[7N<9)L+0N<e@e\Pa_5D-UGE]2&S@4#6Z>+E>Sd#:[,PD^??d-FJ0JHUGA2a
-4La)1e=<bS8>BE&8Raf?2Y>DB[[#I2c17&@F4\K;K^Zg5^K7d1Q(N@OH(F\(L:U
,XT]b.aS2M6SVM/cPa+c<gXUaYdZYYdN]0^V?)<QJdeD?N.&=B959W?eSe-LT#8R
aG?EF0U8;)-228L.Yg6,A]3eFW:?/VPg[?]^WE-B@?:Y2JK\B@E_K@GHMO1Hg.,b
S];8ZdAB\<@bDbCCg7e,F2;R#,4&B86_/;,=^e=)AVF.54^5UCa9dNLPa4e=,)BO
3DXbD#_;AS.8]5:(9<&d@IVMK;WCG^R]5eFI8G17\0WZ-34eAPGX01TL\,Y2)DM^
P^-gTPCA0H6R>ROd]8-W_K5e3=4K,JJUU.TP>=@7:)Y5FgJ&9?1daB=?7gb>.YWc
/L98VD^-.1[RCBF&8d[;B&2<dTET/L)Ec199+WCW;ED,Q64/0Q7\GY6Z&<J5M)-^
NV2&S9>eL)ZCBU-;>GeA_cV<.bHKYBOV,9N++E7WZbAI/5)b;@V#.S(YYP(&GPD,
50VWcXgf;58^/_[7E-@U3C@;AB+3/a;/^O4Nd3##[)44X+#^BONWUQ-H?Z>TF\JT
c?0))DOYM<RB7HW@Qc#4+ZQ^&DEL(+H.X.9Z9T87=LN9WWNF#CSE)4F@P>8#;c42
cQ_(E&F0EWZ;7B)Y+[T.9#DJMY6BD:e+Vf;gb5\723M56Qc;f.3<d5H\L7_Ge:+-
I=e5&7&?^/_gfNe4Q@1QA/cgQ.S-=-^gBQ^=JI(fE:gS4IA@JBH+ZS=OT4W8H/>>
?)/+?Vb4c/YM+^ZcZ^8B6FVIBY#K/9U^G3g<a#8UEfUU0GEa^RbP^H(/CfP/9]6S
)7W[e0/DIX&][X3RDIR9aWNM0d(gVHQCCaXJXINbHbQ.ee-9fBaPKH:>I#@W)/OH
)YI@G)TRLJ17(#N)?K-]@PSK^TZFg1]4GaSaK=<VF[X]Wf@XAXH?ZKITa^A]K7F(
c#<RGSZUH1GC6gES=>/6?7+=9:Q7^OV)B=a5<#7@GQg(I01I0@3.0K-]b2G/bKd,
I\VND;D]U@:A;e?d8&aA:c+HT+OW(/f8SEK4_M6,4/[E9cIGSa_R2#TFGPN2b<HT
6eLOTEP526TI7DN[GBC2P;0);Z38060]F3G#bH/;LSKX.OZ=D#8YX?N8??A\]=Ka
FKL7Z,ObI5/CNIS6-gaVdAXIW\V-=LE#IP.5C^K1R#9?_R)_QJ:(d]FYbMQ1S/TP
)CYIU;.Q(GBCO3.&=L1727[,Qb=XSY+M.?/-Z&TdMJ26A:USM?:KY\&)]S^c:fFe
B#XWdX5WDC7CBY.15UaRb756CQ9WR[/1GH/c:NE09dd,)86L9(]g7eD+_HDLK1QN
^0WHfEB^9;Q,:\aXPZX&X&GO8<>C<7Y6Yc[/VC&53:/FTM1\Q>Be9YUR&0g6dBWG
89WT&43K=;F4CMdP8NH2;H-ES,S9.),RQ&Q)3]8dP;AEXSJe]D/1<UeO,S7:EIF/
+Gde,O)egW6)H<.::ASbN>Z0JG7)(R:d-2(g?XL0]N9dXaI4-F.<]]B6R[<+;Zba
TZR3LKK9(7GEO,[P+5ZE_E76]f0Y>T2WH:DcU1Mbc\\)fU[AZfZQ6:^Ja&AU#e3,
Q]Na==EFXW?U8=SBfdK_Uf2M8ZOXc&83f.g<fgPK,00\ZUO)DQ_=,-FPL@bLRG^(
\U2-?T&CHd-(ATa#U<P245^JP;c-]C/a;X;U(]Q_=;Q[S\R=\]Z.fb2@7=\;HQ[d
KCG^4^.(TP7,@R#Z@=:dd>MM+5Z[A<0WC/e7fST:Md76c_CRBcRT5a];\Td\6\Nd
(a-4WZH=&607@(V1AbHHW70O@4GL]G##7[+_784d?S-XTfV&.])?X)+I,:XdQc2+
gC86@Bd5g-ELE:/0C/gCX.Y(U<ET1Ta,M9OXYC581HU-LK_8f@VH)cXD:10.]35F
_+>/cG1N\C_:1YSYQRD[dbgY:aO[6K42df.4D2^[405A<cB\)0bC.TL=\AE@T^\/
]?.9TA_ec51DeD1-Y4S/XN#LU0OM:bLee7IdD2=HJBDE<cVTB.>YTOA#:HJLLVd9
,??X(B7AF;_Z<&c(;,4/IXR57E=P?+U9_4J,=.c<HS9<F>Da2)0bbX/<_=f\MDK(
9HOZ])0CJ@Rb8V1a9\;ec,b\SK#]@>TM^R.:S(H?>:W4<YPP6ML+QI^E\WT;J_Rg
0d,R:I2],+/d5f[,]EIFRXd]9NPc7X0Fd-C<eGO=#=Z+&a9)I^<J(Z9;[#a_2JN@
RP6(KL==M>2,4^b-(E)FG,_)9KNCCXV+NL-+KH900Kg_J=P7>ZW2bG+MBfRgcFa3
K2E7g5&BaGZF)?Z0^6:1d>X3PF\,TM(UR?]QF>Nc--62#IfA7I<@3M<>#ZeV&BPg
IWTMX=1FXS^)\PW?-@D0V)7.KIHJ\cLWW7P)O8;QCOXXJ5fdC@@NOQ4@bL\Lc@/&
8ZQ)EHb_S1)>eLHNN,9NZ+:D35T2(,Z0d)KAW)dIIN?E2&BMU^Ve79629,5&Z8>a
4e8P0?^J8-^AD.1aId3AP+FOKX=UGg=XB;/Pa+C04P#5=X_W^XSQZIM^WX@EEeW7
ISHW\NA5B&2WgE_>d\b0b&(<]@AWC#PggORYHZ8(G9V2fIR?1QGYVg&?+@D/MdYc
J?V]6ObYb2]<4OHD1VB<&VJ103G\]c:?Y;O,FcSPK\4H;RO)_:R;[=AXJQMZJKL]
^15<9-.eb-):EK_/S-[,#Q:[(SO_.8@/:ZFIXPBK?.H[1D+PI3YU1.Jf#5CHd^,+
XPLAG(KJR3KeOUdW.;;-D:f5BFd09P#-Q\_3GUAX/Y=#R7:Zg?)<Z9Kf<M=dOE/+
NF[3##Q^/__KQYP&gaZ>7=K:3ML?_RXZc/>W0J\eY45H-8H]6HFG.6Wg//cT#]=2
2:XO_cL2eMC;YSPA6X^VC>Oe^[CfK2(V^>6;M_Z^00)FY1#JOY;9P]e)=6YG(49G
.;(NgT]=d,&5@N(U,6FE0==G4VR^GBQ1K(GR81RI1N<,eV3VgLXdPM+M/Vd0Tc#P
MCT+9EF&UFSG85H?D_(GL-AMVBeD,g.#=2O_2Ue<dF?T;BB#3IYFWc,1L_a#HH#H
DX9[>DH8+X4>1e+562]FZ<R/fXX^B])GCP+(&G;;W+K#Z9c9>A4,B4.\^(a#W247
-[@SW:XX?JQ53M9B31Q<d?Kc0#<d]?FfeQRICF&)V5aPUa6bLR-Xe^56TYBMSJP:
L4EAJ,N.NA@&6IL2[SS-Z.5caLWFCeH8^HOeRKNf=^_^+fT0T]R&1D5TU_b(;MT@
&C\9]&X:IH1XO)6TY<0VTg,Yc7+fd?I@Ocb(1W5CZ@>>[_97UFM1cF^EJ55B:#O3
PU2e4.4K98V3Z\3HV@TU89M6O=N]#&B>f\8GD+FMf>)\d[e:L_ORFCX6Y3T&2MP>
Y[<#Y=\?RSE#N+MF>X-AaN@P/]aBBGeb^\;IIQIZ5H6-SU\/])C04#e3V0MBFge+
f.<N_QcX+0W#R(D@WF#[[FPgN>g;e>:\?8a52<S6T>YNN.dX/4,fLX8K^Wd<Ugb-
5AR.X[Ie9^XO((X5Tf^KAF-R[[4eE,aEG.]a_07?<EPA>OFPV[OM=-Za70Y6F8>e
SS<#f]g>8<&Ka4CK?a&&NM5(T^Ne&aYHK^\JT_6HAD;cFL))]8Yg..;8M[L[bJ&F
JZ7A@<N/(T0LE14+?0\FTB30KCZIC+3CM18-d-c>eJ6a8@Dc]01/EVQ6_g:+JOC,
+:Ub,(Hb^N7&W^__<]?LGK>7T]Fg9X-&[G58.R31GPXAE;?E@3_E)?QEW@K(4XQT
7;7A7C95[eb1UQQYBe[[46aGG#DQ<D#^-96+W<G8URJU9MeJD4Z.J+YF-fb2T7.C
aC3:eRK0LF>I+6S/Y8&VB=GT(Y.9[EY_E_/J1U7JL?2U?#;EP5-9]:d=ZOPD(fJ9
#XKf4B[R,:&3@YcR<-(MDR/(K,7^3]Ma[fDC@H:5=/T@[]??DD;6aL/MO>&,R?L\
BQ-T&TEdY)b:<g9ZFS(/[M-7e8FcIP<)JS_B+eF\c-a[LRaMJ+BF]W>G;+J<_QP-
/,;4f-bBdc217#+<?CU=:>SWK+bX;1c_f92X(D7=>e-aa[2)NECU5.Q3<ZE&TS@(
ZT.HEFD]6[?Ag?#UL4a8<Y-9\fCX#GAAcZ3c@JL.CYFUIOb[^B?EW=X0^6g7,;LP
<;HEHFL.<X/b[(8[5+.,)=a=56?1F>I[)3]Y]FBG1=GW(EQ04,N-Z9(V23b>F/U@
)g2DG1H/,A79I-2Rb0UV95-IQ7MP93.b^#NS,/XYG;J,dI7MVIYVSFe+G+>,J9A+
b<GAO&_/TeIXY)C/,\RS7>/?;CE0R,_:RQ@HI0Oggf)VJ\A<R9[eV74K,X]8RAM,
a=f=;;;Z2:I/#]bUIe6CFTUe@7NEYZ4b)###&UYP)[YZ(1/ROHV;8YND,8JI=:WJ
-Pa[^PUCC:FS5ZL55^gIW\[&AX_CAFO.@-bGHW7O.;_=&c-8>gX88#9);E)DgCUM
5L+10D,YQ<@CU#(>XHI8^]A>S.TXJC44L_a\8@1^SANVP>LaI0?,_OO_.Be(?Vf&
<9[;J-4O17:6=Q[fS_ZPUCMUU>Ne#Te_TAKGSG+7Z[\1Q4,eBIYU[^OROg3a2;FB
9RR@^D1F>:L=eH<TVd@O+#XW3-K=2D4.&LZGe@_#2:8G<C-bDBB^eEQ23B<L9gX7
J<1FK;K:R^C7d<&BM=5/XVDHA>>QWS8e(V9/XE7;LL5Jg?C(IaT8Md\L0\G.g@gZ
@SE@IbNgg9LL2I1:85e+a+P=R&Ta7dJAAf?eQ?(6N,+EB053(gPK<[NQX_SE.U6#
cZ;2RFO[g0FBcYL[FCfLJQZ0g,+.N?\]4>^/RC7^G:4O2CCIVAd#E)W.>S7:QO83
S:PAD,RIfF46fF]F^=+N#LgY&M<S1S@@WW\S]0TX(.^]0Cc>-b--_dBS[DeE=ZP4
IPSUQSR[SY-^52&IVV_;;?IPYdLN]g]8(1=(=?WO6f^G+A@C_2]C@fK.I6@eEB0a
EGa5NSSNL<466,W-LC=Cf\,),^TUN-BJ8_a1eGA(2I)cL00[NSfFa/RfMKSa0_IG
B(NdgAUOd&+2T@Z.9_KODdJ2P@)E52dZ+FaUQCY,=<W2O1D^fFXg1>:\dK6PT-:S
CaaLd95LFN4\UDf1g2J<&,H.>Hf+TD\?XE.(14UG)KgG<Q9&WN5_A[;54F3]Udga
2IT;J88[H0S;S=)2UP/+74BHP<D[<Tc\LQ[^MdRD5[6<d53C0LY6]fSS-X]>K)9S
Af.[c5gc+/#73O[DZ5J=d0;;86L/R?RR9aE6T;Sgb[QD?J(Sf5E2U;=J/.4P680O
UZdYW8=N4SeQG9BeAMD6]F2Y[BP5J30Wf3.8Y@(:U/4c3=S3_>7A6R]15=1P@Z:.
YQ,R(WN9#++.I0<-B)Dg47HVPGG8.489+H4@\UG770Sga[B#CSUG9@L)TgFfN)9<
ScFZI0WM4>8=H/RVR#2=U(+RJD-:1><c3Y0.RKA6AK=(FMU#,1c716]R?fU#J@I,
<&,defJIKO0H?XLW+T2TIDcOHX0:cWPcX\J].8+1g8YN,USLZ_U95]?I(YE?>dM5
AYV?(,.FgYPEVbaDSA<+^<^5IL8DZW;>K;IF8R&JJQP_UKI<b3N5&9/1==ec-dFZ
32TB=>Jf\Z6#aDQN&SN[YcS2:RGbEeb<-Q/@HZ_5+]@5[1BBS&.PXH#I<1SH&/49
AWKNNPT.M1bXKCQ&8D#U(/cMFY14:2B+bg29LV+\fTc/a\3d8d]U\Y+ASAH5<;UL
,)#[F]#d[>;N<(\NMM>dKN21+K-bY?=K^STQ-OBB2b+2O5O0U5.5Jda_&0g=FPIH
a6BG_>0_/PS:4<7\0c_(B9?F&K244ZgV3F&/+,>ZK[9VE;R(TYB0gN@a,(-XH-dI
-)5/eA][OfY(.Ccd55X,OBU[Q?:c:]6/1aWf/+Z2&+K5\,K4AdO3P^C?+/5<>4gE
<Ig:VW3JgR=)HRd)@3-eP^^QC^.Yg&B(?e,=:P>NRMcB>6\&\WLZ/@?g-a:I,FR,
L;;)X;&)P1EG+DHJFWe4B+;@KCfHTJ1.VNWd2=AfMM9cf:9@6.JYROYYEYG&&Q]7
6^f(PC-8bX;MMG#7&U.E5^-T=;WA_UZaX&2CWHB+]&+9PGL:?)]&#VKA-b<)YD7]
\?JddB@H)<[;YMF>Q::HRH_a/0^E&SSWR9f(HJ;/8OGBN2QWMZKZ0>,H1UT^>\;\
7U(4+L;NSXHM7697</F65\RZ0bBX\=K],25C2VP37cga6(\ND]Z\Oc]2NGVBJ/45
NcgJOd>[QYf_cTAXMY]2BC_aNd(g4U5):PE([#YCHWYbZV-E5UGU[JBZfX8;dY#5
#=-PXfW)QPZ.0EVGSKKFg1e=de1_aM_];8[bSaG;[K82(WN\C^ZB9EG2H9P1:KLU
fBAaY,^b0&,O8g#FfUG8K8_XB:bV8OaP;TBM=^N9LV#@AY,PR-1_DN6;9a=VZ?O+
B8P-bY\KF)@#a4^B.UW6.=2Z<ARFfGT1QHUBBW8#@2bYUFMIg>H)FTfRS8O0aQ>@
Eg7D&)A+04Yg7?]\L@Ef_2bB4@1+8Ha<IfU.6-FAX^McC<=cDHK+7D-eKG6]MJF&
O?EJc:dE:MdD/@X;[7RTI5:0;UYCH.38Z,)a_^TL^CX,#f#RaIS<>d4[<LIc-B^G
0CeFUd=TV1E^FcfA]GFF^VH+PD(LJECDNb)B9]9cS\54UdS:f\c^2ZIa]JUZUG;9
[WFGAeO@-1_QeLd]WgHb]G-LJ/&CcQg#:(af=F9@Mf+U^QFgR+7&HL8RRA,KU_R^
)KdXO.90YO9F0UWXOK4CCVO=Na0/Ca1R8TYF-d1<Y2?QLQQ53NgA^D1d^#dc^b\,
QHCM8VNY:cG@S0<>bJKaFJ-0GcDV#)I/V/5YU-5+GSZ<TeCTMdQgJXg8N][[YCX,
V?4MGT_dK?JOCTVJ.IUH51:#H,\8fHMSgCTB^fYUU>K==S4Q2R(N>-[WD27CT(K/
8+O+.SJ7LSCUfgZ=d_Q_K?]QW[\3#-LNOUf^AJ>?^fACK^BdS4eg319BPCX[c,30
GS]W.VK>R)A]<TL@L;NT:.@U<?(eSXCZ4dJ?G2]J>AB^L02@\00A>/DDW_N[WTJc
bX(E>fRRMT/M;1K:8QD/U1Z1HfT-KFK^=bb(4[B;II=N7Lda5[E4\GagZgf825@0
P^1)DY?K9ORgD]^AUf)SS+Y=@B6?;[^YL)&2RB5/P,UCfce?dK(+BLKL)#;56(SV
g\I:+#d/;/AXJRV=OZWJP+E?<Y5GTQHX=8XJ/75#BN\Y6OR_e0ZVWN6ONDUf@V:^
REA<2S?O3KHf:d.Zf59(?ZW/Wf/2,QI=(U.&P9#De-<O)1RP9IHZ9_W\e2+[Ha0#
:/=<5;2dXO+3UZ^R;A)&2@&<CTW-,X766BZg1NGQ^TTg+b<d_P7JUVNOH8]-_c.E
a5?J6S/EH8KP\Vb:Ye6ZTD:;ASf[M2eBT)f.&=\7RXU4[/QFdWH&L&0C3d[^\_FI
JLP5L3+Yb98]a#6g#@,?3R<BZ[?VLG_YU>D]&\G:&eP)N<eOSI/=(:f]f8Hd_bBR
NTfcWM65;.V-d<6D^c.E6NG)11B5G,GZ(fAMS;<+<FM9AWX.BZGX-e^T4>M_G2D8
EdT#UZBN6]-44\KQ?L[(9Y^FAOP22f<@UIX&)L\-e9M4]4M>/SY>EV/^U-]g&@<)
H/c,]]#UN]3;U8&^#?V?^<F2VTTSY8EKTHRFH<6CAPAdT13?4+a6gP++&3f:;PV?
ET@-MNWNDfN+E[@Og_=?(FC;3_68CfEG3PZC9<4b>.V4R@T18T)Xb]1d9WF(=aFA
&NVX^>DbD,Z.FX]#bX#Z#9Q?e1WR,^Ka7NLbEI.Ud7N56JR/D_2T(,QeaOfNG1#J
CZd^=QKeO:UYLZRCK-Y-Y<GJ][E2]_&+\#@M4agcL<^TM1FSbIW+IfNBI6O9D@31
7[\DDd&^4VBRAe0#==<DC@(V-_L#[BBd&HP[[a:P021-EBbZJQ>@;7QgVL[DCL?H
TCg#7&P_+3X^CN,cX)H6J;<_-0?[L2L55)fA7)fDL&P#[2IJ4G\.9E2Of&a.O\9<
=Y4,.ed:<KJc\T&>DABO.KFI>#ZATOaO7_,,+]YUJTf>_^f13.#VPR#8V=QSW6],
bGCH&&R_A,M@Ed[.=YMI_7SD>(ZOf+\]&B7E8]J&R>\\FS16M+=QeX[VF@fO(Z5=
9C\_1Hd@KJ=G9DGG;7,4ba3=A)9>);1^OM5^WH06E2[ga,HV/B,6^XRU)@I@&4)3
Pf^&KTO?A3RQg-FgaWbdeOITRe9F=XC[MWP)eb67->CH_cdZ#[B(ScZ3N:T>#L3T
G:)S#)^@7T49FFG^])J&/A9?VW2c,5ESF/;\eW^@)<a6)7,L:>8_7:6e=BR=M1^L
P_4Lf71C?_;5:RZKN]^e^7A.3.Y#3H+/7-f(8a@6CUbe5]O8V&eZOae,KAF>c++e
g6@d>L9-f)_ff9(P\:A]-6N\;aX.P\A+3.BB\1CQCTXLJ=MUd)5f_5<W:_]VKd;N
fb\[UY5I^gOEU1Bf/J2UD4U>IAJfKI-/d/RFTMI[?#@FPd4L6EIE(g1I1Y1,:B^-
<Y70-0/K;#XA#5P(_@a&g00K#G-[b/:-P/4OU^:;TV@PQ1EJO+A\2T>P#>O4[#NR
eRSLf0G&+YO/52VfT0:Q)W8:]CUVgT,S]#+,DW4S-#Q7O[1Fb##>PM/GIS5/MH?J
@Z[XS/BKdS@4P)75)OTB+_<[U61;[K,+dH=K08#-&/PW9EFcc.FB+6:&\U(SKg2)
BRZ7QR#W)R[gaB9cFe^:eKO.6Q?<d?M0CC-c8cO5I9fA8NQ)U^ROFT9[^I)gRCJ_
F109-EaeL2^[g=I]&B^beD)OfU(9&5SagFdGI(:<FB8_(\T(Y=HPQc91X#(fA950
2aL]_Y;L<(e?./==2@_]8866X>f7RPOY.32:<5QN[>S3O3L>A:3PL:2?)NO(&0K3
[3HcK6EJ8EFd:20O+b#^dA&&VS>LF<:S9.A1.AfFLOFf9aWdPZNJ\H(\+UgOIf-5
;/8:3L8Z[]KW7+Q4c5\7>GQa8>=ZeM9fU\=1=K90@9ICdfHSFFZYB8)ggd4[ULaE
WGA#U2K&BXDJV9Q0#D5bYQAX,ca,69)]Z,fO@MT#<[G.T>RL/-H4O,-IZ8@RN?bg
ffC87[;6R4F(#IRG?fXH+6_Yc5NNBKRL\ZV-KHCV+G[JG0a^(e1RC&(F\0B,UWFb
9:+(SNB.f._2LVCZ<D:51>&=(17GD8(ee+UCQ4I]b@bdT>5>7+A2:=#bFe08Vc5K
e@FTM==Iaf3]:/fVX8P>]W_eIe,dQ:@HA8K2b2XaCO^:>/5aacHd[/+DS92MDRM1
H@92QQRWPHTN_1Pa6]b-fK,IX2^XP^@SI]V[8X&S8D:8.=IG)HSXAHGY)A6T2&ac
YHSE+D?Da-1Bc&XYKb?4?EM^TE0L91G-eB:^E0\)]XWAF200>H@JQg8af/]6;X)d
S0XJY3HJ9J5+L0^[M1UQ+A\B_PZB\QQ_T-TUI31?Qf0])?@9,L:,R<76)4:MEQIc
I=UQC?982D[BRKYC9+<:/P8=d;573F7b9g)IYX#bL9CSYgF5^>(M/=M7\#\#.:eg
1c,.\K>Q^ZHK)(@M\g:O#2Yc9VPd9,25^M=g8fPA;/P:R:=2NN<bgIYB_/4WBI;B
+>Yf+J:::CKNRR3gI2SJ:a18P>[3-R)99KFe1@&_>:YdR2<^g@AE7=0g&^>VD3OG
I]6#g?S9-\0dF6?;,(Ba6),A:NM;<?8P2=He_e-;9bOX=?6YC@.,]23He3;fO4&;
/@8JV[AQ5G^d,#;a\<H9c[75b?V,J]X3?=12]F;4ITO8.Nd(WE;12(?=DU/L?.1G
[7dS/]Q\>I1+\Wg246)9g5<9?cGVN1-05Wb61?a)DLS;-ULE7=/GHR(ILdOVWGCK
#;4\5eaM5KII\9]+EDUIZf8GVVK9GF<;I3R-@4Ec20>W2_If7K;;E/Q6SABF@&3[
c99+C5aH<;CbbB7DRP1Y?+7YF=:Yf2gB=.QBgabY16HaXY36SW0@@+T.9&gF12F5
LS]WL3FDE(5)V@_@8EIY2H#a7^Df8Ob[cNDaa^QKfYE4\7)OEM+VL_LJgZD+?MLP
QZa-]=LC1)2:G8HH]AX0G2agR1dc9&_g,)=&IKF<\TP&1WMd0Gf\M2)ORcFLL#LI
Z<?^L157(bN)=[,4B(&&VNDBAHf?9-&4(E\1ODJ0?HRgI?Q]58_-[SP0XZ3?Wb==
.Ob07Db1bTG&H->3G6#FC<GRP8-0GSG6KYN9(Q^MNKcP2d&W?#FA#/A\5#Z_4Y[P
1#U)@M@E49a.eg6#.b+BG0>0)VCJ1\2(V_3H0gBDSC=.)ADcF/6eEd4gfDDd61cA
^g;:?M3U^Zb5RaDP2?a/V]3<16[PZ@:,-Q73LO8bR/#,d9=CR75CPSE=MI@Q1Ed/
f_bCH\S+8<QSI8QF4,[UbS(1[?9BJGNP0Q@LFAG,O=c^^e/9X\BS1VRLICa:;a6)
U?:+,.a10c//EF5S8(BGHNHHB^-<#gSd+=/C,Tcca._:0HGT(/GJ\=e1#:/_207:
SJGa\Z\#<5,XAaFD2VUIgbF;Q2,SX<?3A>>.4VYS8,VZAJ1=.EfI5?G=2=f6K_L+
[;77QT6QgN],TW/4B0RP5_JESG./[1f#bEF,QA9?]R(?\eMg..O[E/d-=\B=Qb09
KU5(B+E.\KTG:HLNeY]L18fVSK1TX\?U.e.K[,:YYcXGVb@?HC-]:Y8@-VCQ\RRQ
&;WRN1#JJY?gT=GDFQE_(#B6GSR5B3]O]YNUOKS1geGcR2Z0?g/S853];C1#DQd]
4WNH26e<^eQeKA6C9,O8UN_HA6g>Sb#NcfQgdBN:-#Q;0F^)#dg^)8X?IYYee)0d
Xg&&eBUKG-P(S.8\H98dc<AYD4H=^Vc#@[LK9UAVTO^NdLb4Xe][(2L#)6Lb>Bee
59>&We6fI6_>1Q7ZNDE(P3cT82QYF?E7.YS-Hd&Gb([IAWJ<1AdQQXeU0</2g/Z_
EK82.,6F_,TdG[(H3Ge8DSJK[LMa&EX^O=]#:8CW8268_deZF:<2d5G<SeB>L2TS
,eO-K;E_+Yd4Q+&,BH)e0DV,^P>8fPQ@XPF4FI1,GG5MTT0CKE32P_B=)cPa<)GN
baU7LH1Bee[VJd[b/G-fY6c:Y&D5M220<=,CSQ5M2X8/@=&FE99H+3L)O??Bc=6Y
C,P+XL;MfCcbABX&+78IgXK2_dV#g,16K@gLP/Z_?a<^IYMJ.<<4Y90H[T9AUb\8
Ae_:Mf_geX2c2#4\?XU41cdRDPWLZf/X7OJNeb_0K6Ke1PI1cJeFYULTBAcEQMX6
K5R#3P_)XdM+9QQ&U,]E6XgAcc)/\K&CER\+K2gG7<gZLXFS,4GcB+5K2OQ+f1fZ
]MTRMd.8RG^@R;c;-9_C)17:]S-H=RHT+&:ZVE/9]e0YXD(]QK;>>J7FC)gA?923
ZG,QF))E(9FdDaIQg5=XO/>aQ617)MCE>K4AU#&705]@&+OQP-E=NIBgO:P#4W98
[>?5a1/QEU?c=KS6TOMb+5O)+200aXU2UK]V@[Z[S6=#6L3YLGU1=WC<]&M\N#-@
?FbIMgCfW_AC+T+3TW+<C/d6+b-(+K>+A<6)K6W+8Ff.:C5H5Wd<6gM2TD:Z>LRF
[14SggGS3W#V1aeJ.&:[3+(#X7=4[#CNL4-0;M?T@D<IJ3UdHa@cWe8@_HXe[0)&
c1B]W=3D@]fH-\F0e<QJ=>_5+X;GM^9OUP1,HZBecS&FaOVXFTH4Rb)Tef;NMSO(
,a<KZdN,381USE:eX:+Fg?eNLBCO]V1S;JRVN(CfP&@(FaS@5F=SfECKRQeM6-Lc
g5MU[T/E[U2Qb5gZ@@6-^WT2-20U6)<Q#YSUdAI8eH@C@D?<<>&9G-gTBA7fJV,0
=gJ14=Q9QZdZWDTB)VY-/MG:+Cc;[H5I(_L/##?0fQGKEaD2VM6/HKRf\LK61UbG
dP\I_45a504T@c.<cZZ\MSa>C<VaOfR-8bXX#(:@0>2975bU7^G9=XY=L^AMWT9/
5@G&H>A3D75g)>_8=#7Zg5#SKG)H7=)d\g+6BCFZM&\=M5-2BN;:E_;#_,aF2/dY
[Xd+,_\fUe1c4QU[1T3[G(D]::N)3S)c<XAT5C,]O@PFKNFBFP,S(La\#HSE7;L[
W;[4Q6[+=X7W+B.Y>ZY/?=0)B(W+L8TeT2XV/J1HTN5J]d.\+#:Ob^F;K?7UaBCQ
=8@18BFLgXb,=@E?4JR41Wa#a_F5c6e5N+V,3HE2MM3A^/6b95(W3L()>?M:Y&Rf
<O@9Re2.QR-NO^G[8XfP)X(;X40-P)fZIa)VGZIZc>ND0\>V9W]EI\[.X6LQYNR1
;]N4#T=:JJ#3e[T-[(M5b[>0U]+(>+a]QN3,e9/A?(IH#Rf+?5e\>?QaA9Z-U5aa
L4]]b4,ZP54eg.&Z6B]3-TP^OA[\8Q5-H\44(/3O,0FK1STEfFNE+9WC)H;\(531
&GT0c?X>75HL)15J[bA&/efF6I)#)RHO2fM.N?S0V@P5M2KY]RQDNIg3XVKZM#>c
CNaRS7;0[=>^SU05H-:]1=T\:]4E;90W:5N_1=af2eIZY3(CCVgDU[6;c6c@-OCO
L7>B75gXWE@bW>:A5/\6S:VK)L?)@W],B,TTDUH]P]N>\8\P>5[,(94<-.Yf:K_Y
O:6\9GT+_)O?O41BG15e#?9Xf@2>[LH-:+;\cN5+2&RNKG1K#Y,DXV\#4HF/CO+@
@g[RWbC-#-6\R?\#G#bSS@(.)<OMaW^]N9:DN:A;DcfUR/G]g<N5P#-a0U-ON)9/
DLIZQ#;^J&J,QMR?)/]bO?5a=L?]d&(6:MV7&g6/+T0NUV+ZGT;81>VeY<YSQTT.
cMJ9H\a@1DE?G=139]T=+/[>LW,FD2C_3Z&@IVb@WKB^0:cK?ZJ:bbET8^+^78)>
+1+RfI_&7.ID@/ZIc_+Q-.D()L2<H_>c#Ue(ASP&>9O-=JcXdGcSZ7Z94f6,T)b.
B][/4#:S3a6J<G.A)463b\<O2,\dY)DO?PPSB-TTP)XZg)eG+H.=&g6>).3?S;Hc
6a2;a<Z>IB.C^IUagKMR9S;R@&c/_?M8VL,74d>=ffFE:,gZ9=05ff\)/KLA16IP
>8QP27bSf4aXQVcb+WQ@5/T^&,6F9_LXBM@?&5c_NZ^WU8NA=01A7U;Ub\AVLcJ/
MZ:E1-8X6Yf.R6e<S^Ha>WBJD@=Y)c8N4,6K,HVJJe?OFDOS?^##2fddc.-\]M+9
<SBDc(35>89NL==e7UO#,f1<<126^+\3)_VM^Qc1UG09Cgd;;8W:f/@Q#e+^5DRO
)6XU)]X9a2/SdQ[?W#0ELg@aa^A@O_#daVN(VM5_EES?/J.D&SecVFK+E40d#]&&
6L87Lc8S5,Lg,Jf;BG>UUV8e5>9KL)38VgH<H0GYPRK<RSf[YDDZ0M]b6]L.O84X
gadLNZId.ZO>]Ke6\2K4QBKBFRQPF^K72/(3,Q1R.b[QO;UDe:DFN]e+F<1)8U#Q
5,_bfJYP&+PC(:_Y@?+dQ0WR@ZIZQLa=QD2UH&((L7X??&.5>3.+KgGG=XSX=IA9
39,/?+2LI^;QZ9fLb_I@)5gAQ):d-F2<,A\][b#(@1QKP95(&F[N1a-b2#Q6WY]]
\\_c6D=I8V;Ab5WeFNE;eeG0^A_]M\&Z<A80?Z_+Bg\->@[gWV>UKR8ZUXU<52OK
7XZ+1EAV-KCGCZd9\OX&]:<GL:736+e1-8d^\L/g&G;8TSXTNKZAP#b^_W3]H?]X
5\bdb-^TQT^@7_TV?BMD:4&3-MYP/C80E&Yd#Ncd:,Z.^K02Y#N?9\.@7RL^D9\0
)IaY=?3g9,A)cA/YT3FFMf)GC#\5291cb@E48;d0Y9:5&H6#>(O\,?WbV73dN0]+
0=PP3+RZL1WC0_(_->SZFQOOAI8^^^DS6[_JEZYc8c6MS@A+dZ4c<B<\:]a+6=4J
RX8&Hc_+\cgRS17cVW[UfCgXZgB3LTL+BWKZUXWO)OS->J&C4-\eYb0^)WH4]dD?
<60\O?JY==9#3#(YGF=D^\JM6H6RT<^:4a@Q4g&7<B)3X9c4]?O\&6T_G@](3C8N
Ng,^>^Q97,E[R8([KbC][2+Hg#F:If&f=CMJE?M@KbE+CYU>/M,C>/Uc;8H[53&P
Qa9+?61K&Lc,cKe8A0)#N57;;a]VNDd_LU:\-dY0dQ04ITOd,#)71:\fE:C7[\OJ
9\\PU\[cM?D#X=G=:#??5^HF]&ON:4NX;C[@R3a]1X\fDP+T=;IF+&<28\:ZG[FR
&GU,T7<);L,@)dfSd\cHEK[^Qb&2PN+OOY=&_4(S586J:JfUD6Pded@g.3&E+[0K
ISe[)N]AB./MNcV0[cd?L8C::51CGLZ\(N?E\7?R_8Me13^TM=1#GQeZMXfg?)BJ
<DL-CNL1d=W<<Bb4\R[]DD;@6R6_H&-</EWdNdO##b7YJgE^7^YAY?_88GH2P,ID
2H9eTX=4.V2)-fD#7A9)egdV(2MI](50Z4O\U,:R_@f</6da&J0@N-O4^+g=CM>Q
9.OCIP/\YIS<0b)D#QZDW;Y:cBTA&87NHLF,&FgYeG,.Nb>5\E(cMEaN/a&F-b4I
+GF:f+DZD-P_<c(1U^C;CTPG45#f#5/Pg,&Sf+UD?eS1=bcW78\=D+9Rg)XEWFYa
[=a:9aLfQgIXB<e6[_T-PZ_U)Xb8aeQ+O1=3UH8AdRKN.UE:SRb0P\Y&ceV]7)LJ
6cF\-4BF:K@U,X]VH^RMO=6,]aLAV,Ob04WYQ1A8QF5.c.-Q.IE.0+MF8G,Y.&LP
,-bYML[QF?GMJ+&M:9)RFB;U755HP&UNbg:NEYIF=F6.7/M,EV>2+P-_1PL7L,gH
PI1Ra4,BAeYE>X4deA^<ET=1?Z<FP:.__JR\LEbTT,Z3(]I-QQbEedN.6X#4#b5T
?X9a0-93c-E)]D2:g6-A5+BZR9]Uag<CfM2H3RdU:KY/L;S5]=NY=S/#A_G+gLY]
NHR;bJcd3O/LENfb(G3U-;.9Q=Z0,9_EX?OXB,/^NXf6ddaHBII\0bK1HbAGGB7<
L8PaRTMU=[a_A+R(fXG\5F??WY1)T@f<M1]0;Q0E#]Z9d8CNAB6OR8\1+S)5J#]8
B9TD2aQSX^XP0SVTQKN-2[-bb&=6+<Z>=>9?07g?J;=5#>0)Ef,V<bBU(R#SX7F9
)c_KLVb\N1S8/f<KZaGH;<#(R<^,D1NF+,9JH6EcHS@WE1Y.R/=W:I+6fJ?]C52M
./ZVIMCB24I^ec:?&COT?1?)4HIZYKOf0BPcDOEMAR\6Xb?MaZ(MK.(P^fCYYXR7
XOgMI3^]=7HK,,M-E8G+P>0I:O5@9D_:.E=5/g2I1/ZWW4YEfF5K9^7=Q9B)_\Yc
]C#Cdc=M@4CSc,,]#:g)=G3QP()ad&=f,e)g:YI\TL(1+R:O8LaP?8>#_]DQQX?N
>bDL=bN^<b871bcE5DcO,=-V#A;c#UKCW?#^=JSdXG#GG]6])NR=,F64/Wa1\TW,
6):0]H:TJX82S_E+H=#=@CSC>OKFHR0^XP7STbbfCE0X0WGB2B8e4L>K,:\.^C,_
H7(WTP4T9NF9RX-fZ+76g0)7=BeLM1/7Gd:@O#1A4<13T0UX)=.\O0Rgd4G-MMG>
G_N_e4I=R0)]9H1bQS^cM<-Eb>#);G.IPb::Z.U#WI;1+MKBX7MZMeF),JG&).YL
f(<K:/C-IX#6CH)K^S-0QAMU5TDOg[><eBcZL?53M>^gg899\.ZLMa)?-=]C7#LK
AbX@,d5)a?&U9d@LbPO1V?;)=J?8^XKMWF]J6AT.=]]0+,IaAf3:SV6G^g[O)N<7
,[5+3/(gg97Uf;O8@0CHB79)>[:eY>RIP-RRb<4g/L3_bNfEgZ2PLge^g6a5V(_W
SS6cT-0IE9P7_RP2e]&/?Yd:cD@AE3VaY=dF0Z@G/QNV=NCDI<GXbS\2P.8M=AaL
OP=J:#GTG]N3&[Q\c5:g](6KX(\g[6@&FV7=#_KV\QA_OH-5d5EI9>PBQ=aOdFTM
2DQ,K-(T\a4X0:<6?4g,X8T0A_:b7OKJQNAbE#)XUQgd(<-:VCW?(S=fZW=([[,[
,fZ]FX<)H[_EC/\U(:I:-TMSE=YX3AV=[\,a<#YW(-/B::D(<?OL6\NRf8fZSUg7
8a->Db]P2Bg^F=&7QX-;Z-LLE\e5N]/L3J[A9A994H.-FVBEJdPIP^9O(=CMMK)1
?)1fLKHgV++<a:&QLU68P0D&R9N.0g4,X>7J^^[;]IY(PAUR[IDZcg>#fOB;a/cM
)5.d:;)U#:eQ7g;YF[aaUa\IKe;(g:&_/K3WePYb5#H\0UFV]QdJ]AfC-GWXQB,M
aE,O8T>46e6W[NHb&[<\L1?1XMgRYZL#:#5X5_Z]GOH5249^0gJg=+\+@>X7)I&+
E>8dFOXHgI[\O+-e<dVD-YWP/Caf5b=^3V<ZQ[U)L@PEO)Hg:QdBB<FeMS^OVY#,
_?O2QBA^M7<LHR>IXHFQ<[Y9(3DA,3-(-&:XGLYY5cbW,SaD2I(YDO0\8@c1PIHb
\M_&Q9>,<&Y1f(VU>5J6[Y4J147YT;0HGQ&W&YBSZGF=.Z+;_.N4B[,TQ(6eSTM\
IHHH@K,dZf7OKK.RCU&MOO-\R&?N7V?.f=Ua?79b90G:>PQ1d^=RXSGd]]\C159W
/]^1_=Ic/NCJHW)7PGfSSE,-M7AXgG7IIK#D\B;5gD=+3dLV-<2W&#5(.9NcU,WA
[?;a?3X(TEXN@dYaME6EH(2>[C0PdZ1A<\[-3T0?XD]H<@^4]]W0_B5)Jc=;-be<
?0U]?_RgCI9#GQ+L?;7V3P2G\4(HcTA6>LA7G+:R-cDY@Q//a^XUT)2X3B:,[1We
@7N\KY<OOd[Z\e&-WeQQD[)1MV>A19BAR2UVYSHGg-Hfa9f5BYR[9;^@d,?/-=ZV
^&>LVBIfbHN-7B8TC<B3@BB0FGb,]4[M)@6g-_B9IQ[bI=\]b+9KJ@3)_:KMK^Sa
Tb&&IJ\?0^@J<bfE#VXSaQDTXdJdJT^_P6@HM+Y9/02B-HWJ>5/+g1K.<CGU-I_/
OS_g]4EMbb4B-\H;XJ&7-CV6QS5ZfdgcQOfWF\&5-8dUHO,U36YV7MOBP.+]8E&C
0A.7NUBM6NNTV_?(C)SY\F0?=U)Z>7HdK>P3MfJTe5,XK7O&G,f>X,SY3G,UWJLW
[.g]8Y@0Xf]LIC/G0DXRN^cBVX1;PFR/FT&K3bV<,(^B,^(T5N9cF@gd?S1]b2T,
eV.(/O.A[:9(dHG;4B,;&H)3Y;>5B_Ya:KQC7C<:;I;9P9G4W@9HI6+7=W,&_dY_
@O;LaN_X-:O3>Ce/EG2K?f969d5MC_45R;9)A52U:aAK#Z7#d2+9M42XM/M>a=&I
-a,0FL+GGMf-1DX9g7)f+\fCW8]VU4H1B/T#@TT+M^VK==3OE93d[V]0OE.5gNJP
gfV/[OUW60^K4,L=g,&QL&^DF&->+-9O:-?Z#4]8_aUP4.A^E&^d>WZ;51;I8X[+
JE_N;RIUEF/VEF9_/Pcc:eF?TJ[<3SN7L3I-F06Za)3\OLEWD3N67S.>T9KY);#;
^68Q\&8QCb=,gH@E=3/K7W.:7G\=X5?d@]cICaC;2O@8(KUM6AE[7TT6.)De-;8F
-U4a5CK[:cZ5OZ6&ABM==;Q,Mf[@U(+(f51gA,^gIMIN2VV9@V5;?=&,-a<J7FF.
J\:2g:7ZOZ0[Ug5\D05[QE\[NCHXe)&WMaC-aDZLRe_4CCC1,+gG8##^G^<e[)b4
E\;bJMP1H&^:;#\O5_gC#L5.?Oe>A(M)C<OC?1]>?S_/bU;(f0V,E\/O(7FI_J1M
0QDA9+<4]W6.G&[ACX1DM&2U+)>Va(6P<\CQ[C@(OI4]7G0AgTQB5HJ^#2SNggAT
#gB9@::;E?A]C5-[;H@Za?Y5_^GX5fbPL3>FM#-=/N\SM\L6]^?5FOH;g4YS)]cD
\/c^>51?[TCeA9+E33J@R(2,a8dVDO[Q5-@C#1;_/d-GYNe6/fW@;PbOUZK[f(T.
V><Og=1=&DSV>Z0^[:#W?.4KVP[,(U)\7S@O24CSJdg4LWeObaXP5XLACEJD^:/8
ZE:8FODIFf2LIMTH6L,A+a]FBT@&dOgLWa.7_ZMMeU/E1C_DQcG7D>_0a\+KaXPS
Z4GUeO#([)G(1e+cV,64]3VD=R2AS)\3]^ZP;29_FTe+>H\L/3Jc#^O8gNd^-d[)
Ug_B;D+@_31<HgGA_SK#+L-8C_/N0HL3A7+Z205K]G+(\[K/e>8M[DbRBXW1@dL>
30)L8)ML\TE=+XBA>Z0TWY8a98PSgMU<d1BD[19_M6]D?bPV^2TAVPWAU4;#^84)
5g6&a=R?9[44&6;WgP\&^7.W:PH<+SJ9EG7PIR@8cS=.50J>L5V^2>M(]4>QXP]K
N\TDF:NUeT;\ReU-@8N6MP[CV7T1YS9ZD3>H\C&WROPc9A\HR=S+7:Vg6GbC;U+1
>cP-c:+67E;APO5(d(OVYDA;Q7PD55V:3B/##D9V0PYb]ZZI+aB_K)Y)7deJPB)g
[bD@=PLF_Me,#N.NR5@^95(K4bBfZX-,\M)F\a4Ag^N95:::3UD#<g=Y=fNYT..b
b\_)?EcDGaHe3H;+28a=M:O9EJGHK^bb7df7LDTT;XVX7cF6C.4?@W2K.4NJf,CI
U0K?Z5GW_NW=2T#+.DKM6&XH0=[48N8;XW@?R,NCT)3DZ_M]PN1@-N(^LTG-GHW9
,_O+JbX+]UOdZ;G6X0UbG.4(=SNI0RG=U8ccU019^OXd\EPA3#dgK@#V0<XPBR0.
7(8E+_Q)3AB=?T:Dg-+HFJY\6F)RL+@D@d0E6S;[&PUSPddN[G#EB5.)LQPELbb^
dCbBQSSg11MQ&\GC=4RRN.dA>6\@d<Mbfb,bN;XR[:T^3>0R=1N-@R0Z4TRHg/O\
Q&SATAg[-PH9W81=ZJCGXA4>f/AUcW2ZAIc>T&XQNV<P8HHF>@\<KRP(Jb<0;_^X
_4c7TM->Z/YM]U-MT_S0Y20?NX>.5=;@DE3b(_V7NJIGE47R?\[Kf>b87_MgGAX=
:&.)OAb:GGdNBF=X(b1b1TCdbbgV2K\L?[NQ_0SXaWLHaHR;Ef;c@3\TRMIecd._
>8WDA88P:P5YHLda?KFK.]1T/bOa4Rf\LJ,G+^_NPSe[N\@RO+,H[Hb\RZT.0#We
=FCSOQ+dGGbRLYZ#TJW_\309-H56](d/#Fb/Ac.e4VJK&P=YXb5#a^81N-I9UZHB
_Y,Hb9=7A,KO64F3c.O9A=CAZ@P\@13,@2L^dUO=Xf)=V@<#SBe\4^=XRWW)BeNZ
1dU;E-F<AO?8[eAS>5)-Y(?Q0P]Y985Xeb40,WGBaPKYU4K>ZXX/aRHgb@_-_fTG
,aF^NEc]M;P:P^?cBD^D\/5\3BBY3b^3FB)?^O2G0NBT8>fGRD;)=VSGFOOTfaZ@
FIV0)8W<#M@bO6PU47;)98DMT5_cg5#</I5e]TW++JVg_C\S)#)0(-aH]/X].a.Q
8ZTAbL]e)e#8VY?R9CC)K?Q#TTV>F@SKFI,MO3QNOAYE/7?2^SNU9ZGQ8f41T,2b
f;J+4-TMXPK0dBD+74+2==30A(.SZ<WA(R)<(+/E:PP6^cb8W7<F>ZgG.6cMCbGT
,\g(e(IdEP4DJIS5WRb.2H2.D\Q6@PH9A/1P0LSA2.-8[GSL7ZN7f>4d1ePF>K[V
T>G::O-/aV]R.R,]ZO#^B2C0fO=]S(LJMKBY3U-gX+[DGW-f6ACMTEG6XO4g/>8K
Q<2P#7,R\9RTg-)T9G9,C)#8Hb7MVMZEO?:@b-9fNZZ(->f&?A3.RCR(a9JM9.X\
#CG;600-S8+G)1\eX.\d89I36_4NI7:CK/gCPNd=-T:F3#V7T[UfFXI8Hf.3A+Wd
Ja<B8Bf,<(I.[5Fc_-E+S^+<:2]L3D?ceC)A4+gJB5>K6<b.\9cV[-IST3V+TaCa
+4B_PI6BNc.bB&8dHXM01@^88W1W?:WK(+)FN3D.GPNaO3N#[e2-<<(B[D):T]XL
H>bH#>E\P#NK6Z4D3R:\S[Kca[1Ba(6WG:QBBLD?FSg6[J(6_3Ub7^((dfVCK2U(
WY4f=M#U_@[^7H&c5W)^8,bUfLQW0YHeM&^be2#CDOJW+R=X\../e;UQ3fA,0;2J
ZHQbb6Xe)<^YZ>#e)R[ff5Yf;15V\[/96:E=E\Y^:(,dBZ\E2d+O?PCR(eE?I1IU
]RDBW3\Le-X(L5-54GEX:\OR5C^ed@@b\Tb>GL;7e];^@O6=bD44cGL[g,UKKPdH
SQP8dWW95Q.,+)MVggHPf^O)UQ1Ycg?BLM7_g+>[1\_&-74gDNS-XGJ3\&A2=X/A
M^>KdbNf#gNDdK_T6gS&\G46A)beD\LODO).5IV#3DHP&RI]M&e>48NVcOCZ:5O-
4;AFg^.\.3Tfbd\9gfC[RK1UYY0UB)cJ=+&9]#6BB-AQ8#8-E<[2#V=+8e)c,8DH
LO<@X55G??\a#<K1[-(LOKUc9DaCY7g&6J&I28SK1)52RE#bZR3DN@Lg-6+JX@He
59O^9UcG+H[<50B6M5dPNR04A,gb>BNU?3@XU@cGM=/>[CRc&5^;=f9&V_(>W(?7
dZF;=K1AODe/5,)A)2S:[-&1]c<JbK//U4^KB4T?\OWW,+)67&S-[C1Jgc0ZeW7(
7d95XGWMMJa;Ee\/M5H?;W4)]B_M0Z.,K8YF:S521,G@5@BJ7+Kf@:=ge#R:<6f1
RF2Q<BQX)7.+/)eg?dX&aBTgLV.XA2TB7c/FAD1_QO4__RVLMgQQVX#gIFg(CD(+
>Tb=KEPfD>e^[;g6Z,gG,c6271;X#HX?5X6;gdY\29;)W\0\02Pd,V^OM51&:P?>
FZReYF42dM/#bTdeG6)XTZ5:b>LD])DK\H?0NZ#^5b[\2F[G<E;J@2B:HCH2@LRa
dU>ME@1NU?6++@8K.g1VCbgHV/,V0gVaX6?RZ)P]88@7#(eA3]dZI]2/1d=^B,-W
/Gb@O/Gd8Vd#e]FB;2HcUYX&e>ZNG0bgWYVFG#C=S,Z8Uc91)LR[N3>fO,d]PadV
XY,QQ?31(\Hf^B5/^?aYL>&DY^62^70;ONC<2bTWPM>7;6./.H?</S][CfUR7DQb
-a5-JTE7[)cO&IO4NYD@&^,_JYMF@Z-J^JUXgXEQ@\J-O1e;VI:F+3eV+C\1LJdb
0(96F::T0J4\d]cYD_ZP4S@R6#/6dGXf3Ad0U-#5bN8<@7KSdH_B73.R/^.1d5J]
ZI<]bMB#Y?2Q\1R&[3_:1523M]5(D?T25&ad:eA-GaA>TS-&P@MKQT:[>9\EJFFL
T9+cIaWCaAOYL+9-.0Y>O0?RaNg09O#CKa6@eV-d@3aGEX1Y_1C#abe)M]CYQ&df
WOJ7D1NbR1\=\@f8^aTQ_5^ST3GN],G,>^^>RA.1;5BQdbE=^?ABgK#?/b:LgW76
@Lb7Gb.fdIZ/-b:-_:2W,4TSITERfK7HK09X9PFT6?AcCG9#a/gC7##JIORM2LA7
65N,(?L7YL#4LS7=7X]26c-X(@FB07PFDOgb,7S+AJ^A6ZN59E?S(8J^HXRUcTdA
b7F,A[g#0MaQ6:=<cU[NYdWH5c#LGJW0g2+:)20S@GJ+YQN+YKTgd&bKRfW0[G;<
B9BI\F]6YTDL\7I79XfYa7fD^O8b6<:.&(;ITLSF;7-V6SKaYfL;H5TV//WWEAJ7
?)gF+4EJ?4LMMYK7ZfcP&_YDK1]g4#]fSXY[[feO?/<8/H=)cAYANSEcXL^W;6\J
QS+IXd.#2ZPa&(RH(bY,-GVb3UgI,K&V(Gg>(&@/Rg-3=B_TeX]:UJ.51T26\eb]
:f4D5HRQMBDWCDJ,#ff6XP[T7cP);WaX?=BZg18Rf0dE\;)R?/@5HG:AJe6#GG78
#G#H8-,I6JP8J@),SMaZ[cV[ORA)8afTHa<1GW\(6#;8K\f>DF@<QJ4[@>CW4Q6U
AQJ7F7X88HM]:X?)d.HJWVZ-,1bf@0N.@@?EODX8K&_KR0\b)/g<f+=?7YO1<(4T
.3Q7Zbe1,S[LIKS2A+<<0#>f<]Xc1#P@>+OSbb#fA?Nc_WT(6+KE:aGOQKReebH6
N6bSU->Wd/:D^ff7(B:L,,XF@ZYZ.][8KUg9^Q5(HP014T\9[HM&1EC/B8_#><5(
92ESYO\^g7,=B6e4?gK0a1VOa84b8I93Z8O3a0cBa.D+9J=;AaaB-=PSN6E2&<=c
fI@1b=VTGHBZ5BW]P5QJF#fNQHR/LMA::YB,GA3=6RE7FPU\cX[cO6PTV8#(M=d?
3@Qce0BNSZ8g7=(6a(;VT,3;X/+8Ze9HA+\F@gW(=VKZ))Z^4U\1.f/(:=5)NVWD
A;DXf&PHB\?1&Ug/+1<&K7GeY?\:><^Z=6<@cV_X&#RUH-S1LG.ZU0QZA+(e;1cc
#@WIE95GVSHb\?[OY/fX&DL,SK][Gb:27#Cc&_ZcLFM4Igd1\QJUf)IBK5Y-F.FP
YZ-OfAZgcX:YP)3_N7g](6[eAG1R/N.]+;.eA??NLVW#J=31g4LGUU_C<A_,e7d#
f1D\Fcd).4RLOdM<V_ZLTDOL0a5fF0=e::#HI<1eKf^=;YS0@F6R8N4fC##91IdH
^U,BZ\A#O@)2(HWgH:>4NH]A3dJQK>P7<,[1F8Ma(>LLB:7Q-Y&@W>CAb5b88M2+
<TW@#YLYfF;DQR&@f#bLR@.Md:fV./:Q__YU9Bb=2b&PH@(H)&ETQ^Pbe-@SDA#E
-a8X6B67SM9.;cSE^LOR@]FaWTITfDSUGM&Q\2CKb)#/deL]24/.3\aJ5^QNAU#B
G\)4-4R#gW[5A8c#I3Me+d?_)T(ZI/SX]:P,ZUPM;\W3:P0J:H+Y_@>XJ8bXS(IO
2UUbB;g@&PO#KD\?O0N8+C5eR5[+V9DR6E-+=\5M0Yg;P:R]C(E8D?f,CG:dU>[_
-dP]?JU9)ZA9>\VB;?SXCA,cCZ)2fZNXWWa115e38P;:,,fHXR?&6:&/^A9Q94F7
]CGZ??GQ@D??<;)0XCZ/<9&>]EG<A178df@M_AOSL@2OaTY[Z213O/c2#W;;If]F
]&&X@QCdL(7<W&7#BL\U:W2.#9@);YQ8f+H(35e9TQC[H6P;2Q378._X7&R@b8\M
5;Db1eL6_X;b/c0#\S-SH.cf^AX7LW^3QL+bCf74fGFcTQ60#a-(/>D565X--^1>
(=BW#8a(gL-I;b:RaR6>,^Z-[6S.9C0)P;WaC0Ob6&\g^XD393(10]@7D<IQ;4QE
U<=H^YMT(a;[I8@MHa\(5?NB5U(.=6BgC.J7TK.XM7E6[EC(B13d=)ZfM9US-L>\
J([;>ZDWEV6#37]DE#V>ULb[+FVTc1(/]65;WB@MBa(A+ST66(&G+NbNOK>bRA&7
C5P-N\d#3.Q=DSICL9+M+1/Qe&:IDOIZ;DZU[#G295[SdLI4[eUA@.8)DD:_LRU5
+&H1>FMb/HHaWKGGW4VD#KW_[AM.YZNAUg(6?ELb4?[PGA7Z(bdNY,^&;ON<I1P\
BJ1+MMR+XBIeDb@QOWeXBcd:)H:bI)0V/P2.?JE2cF;2,8[gBIdC@EEA^>]VDD8>
IKMV_3PI,(^0],2f(XDOFV7aYWWYE.+ScD3OF=[J4CH:9RgfUB>M.L;SC,:>g-NT
#RNKBFTS8a:<P;741&:C\#+SJV#1CUKc<D2[f)DD?S857-a9IcPA##@#)U4XK6GF
M=CTW?=gN1NIKgDBNE>X0H6(b2N9\Je<\QO9\\dEC\YSS)S8&a_X0TbEZ[I0&DPV
V?CAT@102>UC3>HR&.E1K8MF+aNLQ4#]?CXIdXJMLAHBB,C1&f1EV#/QC\9_(;9I
YM3K9EK-3FX-#/P=H:A,\)M9g>^)SZND/6,[d<fb2/J0V.Y[8-7N3eTFfD?RVdDD
Y>YY.1,R0AXT>7-0S,^S-QK&5+BXdU.(><K6ON5(ab\X?Q-eZ>,.Z?-BGOO42JG\
([=HVcO6AS<gWVbbXA[+Z6P@J/\@/.B\V..8Y97,T)DP&f7LUMJQQ[:E3@7CY,:^
8_[\)RT43O3;d;_SXFY1-F:+=2-e18<K.YY,LLe;F8;)VZKK(74W86:7NCQ=-VKD
YcaPWNBI/N/9DWPFCFO<Rd\,XUHH)eC?9XM7YEfEc8VC8L69AZ[MLULG#PU&WHE3
VbJb@cFHMf:-#CF_#[+Zd+=E-,f\+E2]:\^]f0Eg)9E8b5BQH)TP5J\4G/J8[S<Y
\X&M\8EE.:8_0M(gbA2fcKS(ZE,PaBPYPBPJ_a92+T;(2_:X,ZX[H&fTRY@BE2:.
]HY&XIEIX=D:H)U2&E3()N.6Y1X[X;fM]Y-+5Z:/P_MLZ<[cPIR(fW1E.3e_UTGD
KFO]G9<dQ/;)OQ@I4@g(@>7BA)[g1P2R)\?,I/Q>[J/fH=:UNH.e8)&=<S)cN+8W
\/,_/_-5dg7<]b,=C8d/@^GS_VG#78BRfM,V<B<KI>,4+\R_&D9SFZ:Ze-.1Zba;
<eb?0+_TY8CC3dI1c6-M=1,-/;CXfbD7#3+3Z0AETXK&C(.R]dO6)QR]=K1IC\S(
BK_@H5(ZH:G#9<4]FUAfW@^K9H_8(,/SQP?Q9I@D]WdW(JWL<0Q\:I9\1Qd0MdA0
;QFQeJ^Ug[Uf?gI:)D>7OO[&3+A#cM=c@F)3\>\EE+4G@&-3JW(9\/#T3:9[)e2J
I]+6)ML=JI=[(NA1@f;@gO+@RE<EY\<cD11DUY(7#Qf=6GCTeNDK^E80(+VF_R9Q
Y]0-FYGPD_a+56fa&H#<f+FII,R9e):I[=0<D=2aPdCCSaSEBd.+>QCAXI+;:2<&
NVB6PDSL7c[JH8A6OT9:de>fJ09E<N>M66K_.=D_,VBOOI#f=<,I:UH1b<-5Ib@E
>H/BH^.XOU;G<\c8]gbQNcUK34<6T/TW\6:6NH0W=aLE=G/GYG[fOX-aGCF]/8e-
-,:bY+#X=NF_<>+C=U6D(eU.NfUOR:)O[SH18C4/\HW+]9;6@2FY+V]DgWQHY:2(
DaU?<GcIa8970X\Sa,=_A/PR/\If+#C;JS1<dagc03WeLQJFT7aH.b72fVM7)3XF
Y>.MB77d+?bJ^Y&@SWMcRY:9?M_BN(5cH(1=2#KO5@0eF4<_53+7CJB8DSf/,QF=
641X:e,KfH]W16.R+Q(>05Yca[,S4_f0N;Lf3P.JXU3X4(<9WUPG5EI#3OFD@cY4
KW,W#AIPZHf_LE[dKULe:2@QgTPA[H<H3Tg](E)RBH-S\N\+Kd<.=;^KYO_WTe.>
&FI@KDa?V>KUfFM<HMFR>J#:]L11E>g\)YO#2QeGCEe&Tc[VH(8WM[7[#RWQ0[Z/
+F2:/_R?J\RE/_@05K/:\()SV#eS2@SSKOeY\W5+YM+3Kc.I9_7?50F_NZd483?#
dNLBE,_A;9,?LMX=/V=c+NI]MO2Ka4.7Z@]F_3-#-K)YV@ff)[OXEe8<OA\W&3Y<
,5ERbL2SXd]UR_<XOS_G<8O=?83\JfaRMe[(c6MbH6HIS_Z]d:+J04@([D^ccQX6
:UK5I2_GEg;NGE,57LW544U93N/?RJgR70(.;;X]b[7=>SD@L>d:REGJKdO85LFO
SS7_QDINP1/:8^24#M1UD@Q::5C0)8RabYaeL\SCa83Q6NC_Q7M2PZOAO7T=Z^B>
MGHS<F]4cagLLgc>NAHVZE/FJ]Ee7/OW@&f?T+.UfgOIg;RX61T<#M[P<?XW+P_N
c8fF_4F_b=H2ZUBF>MW\NgF6^eI=eW^-N5@+AYKE_e8/MDD>FO[84^5]fca,Mcg=
G&.\0@OPYC,J5f?@J0Kb>gad)X_OSagE,=+8L;AA>fBI/UaPFA3W\D@;4R,N\Na^
cI?eH1?J5G>]F[/WUUQ6b],F&bY]46AWB>G^Q5W#YF]84=Z+=)Q4.UWM8IX8<2&8
5=D+H;W3PN:P6+0e-F7^)RM4][L8BaEE3A)IAa4D^0f\J)DdVM?_KR/L_W3PJBHB
U\Ac2J6]c4(3D(R[>d-48U8H,G,OPeDB]b34;I&1ae1:)R;6dYRO.^^L/ge#46^3
(C/AD6^OK8J2dFI#gBQOb24GT\4bFE#S48XX\=5:F6cFU=J_FHV[Y9Y1\Z[f<#.6
)5BTbDg2SbRM?7e1OT.::L(P]ZCLI><B@C<KgI@XT64T#SGg]?Q2cK9M&P6]<eKZ
#NdIQ(=.,9#QL[f1PG056EGE_dg^E#C/1bL<+F5]@B0)W3.GNU;d65H1UKDMK5\)
,HL&A]QcAE2]B5[=8c5TKJV_9L6+0cZS;Q.DB5/dfd.E80MXPEH/?@L/?I<c_:Cg
W#U^cG]^G.N389ZgK)[3_bZ4b]:O5OGNXI30A:9^6S?3Vd2G_P]dTR6>eTG\CGfM
A7cSDH\07#>=[3?[<;WZH:[TY>N_UPAI63?7,aO36\2CS;]9KX_#5^FZ\G/@KDF9
?DZcf+<5^)NQJ@T]KS<-4^&d[ad,0:@AX)aIMfB-53JZ<I0UEf)b+6ZO-aNLdW>C
R+[A_7:OKMbHb/Y_(#&XGS>DAM)_U#&,-+dUW]++]YYL9Qf7e3QPL,A.?4(D^^XZ
2G\P+?7#CVfOa2;8b3ga9E<dC<^Pa8@d6aHPN):-DK(LTBR[H)Q]Z?GK+WVb0F3S
-Z;+O3K1]9Q]ZT6#U=2<J?bdge_J]F#B>ZV3FM/4XF]EF#NFI^D&:[+Cb8ES?75V
YN6)cOd;e5I>d/Cg6eBVN>;,S?:[;L-FZ0-7KK:7JFMI^c(==7X>D7gLL)/dZfN.
4J;N1&aGaSPLDG31=5C#5&EUX:84OVW,ZfUc-UC8f:V4D?1?bP)J:ON8[Y-V?QO6
=A)VgX34X8+1ZAKQ;d^;BDa5eJ-M3B2d#Va<J,e;^\R-cf83Z12F7^J141RXHZ^&
?J4(G05F.0OCGBT&a2SZZ.,2\=]&6Yfd=>R/\G/SO6=B^)e\a==SNVge37:W<<I7
E;PDP/_9\Rc\P?NIY;XMPJM0#3ISZ3e1;9D=?^f.+Y0=QT&\#XX(/Jb9AG6(YKYN
A]VJP1-V8SB(LIX6,A?b-HeM2c:4MI.-ZZ&^6,7@@W(A83J3,S[[Mbfbc3+#DQg=
P=U.IGQbdEe0fZ.X;RT;2X4\MS#QM=IRJDaY1TW&,,B(#C;^@/2NCO8QE[2^#3AA
5KPE6QH\:)\Y?.H.U/d\f?A\+.g^]d;K]Y&]R-5T)\_3&;B;XF@R<b9#2UH.65(Z
/Z&eZ0E6O>N(KTZI]#Yd[c?V1MQZ9L3N?f/9[d._#H-:&X53G&<S)YgJ^bX@+gJ>
)OOgbHY<fS.ef/F@#V=LS(gPXKH+Rd8&[TES_<8AEK.EH=W,NS@[eaJ_Q]WA05^J
59<S9Z-&(TUf(U#f\Y@?H>_2@6Q&55,#\=BUFAcd,NK_/LKG.AeSAQR8ML#;&O@N
4RgL9/Gb3aHeFQg,0OQ6OcCZSgK/P\L1e8>2F+LF;ML\3Gg;R(Y>KC,,-NU]/)B^
d7/TM_A0Y>VKO^,3YSE#KT]+.4C/PF5?CDA/]Ya?]1;7d[RMMN,=L6\W;/<_9-)/
gOKK5?YN?-RY_;^M7,T+GAdfgN1aRf87f9)NT+f1>#MROU.W9J88X4d\808Q6[WP
X0@[SSE1^THfa?^#CC4&YcLQg_B\NY-JBaH]@316)#bFX4eHH,Z53V/,;gcb]((>
]JK2>ZJc4QeDOUg[X0b#]IgJ@fQ-SA2(ICZJT-VW,BA7EObA6VRE3IV(O?5U\5E_
^\<KCZ9@&5EA4MJVXNFNN9,-G-G)U)^C.:8AaOfQY8J+Hgg4C]_1f,9-M8e?<B+M
D8UfgO_ffObIfH7^F1-BNR&-BaaS:?c]NJ@_0L/[_e&W2SJ,SDT/,.SRNS5(KDce
,A/JUb#XgV8LGH#b9U#Xd8C>SCJ]+08WV,MA_EAK[a)T;b?]7eBeD9MaO0PEN(,+
PA&66X43W96&-\?bfC^RaK:3MJ(R//T]-O1IOY&[]DfQ0c;cZ2g.I&?-37DNW+d>
.WdOURCWT8HQXgHHAQCJ)cERK;:6/1\7E/.Z3)G3#U7E])[(YHQM,=R&7N_:N-eB
e5_926<@\78Eg\T6JT27()H9P\EICGOcY)4>6MfS\-8-VEd2NB73KgW?-@,c@Uc<
3Q;.L?1gQb_KKa(ZgX;=DgW^H[P:[X#4Sd=+;RQNaYXPQe&:0)>P=T<eWYYb045&
WURZ7,BKGFafQ/=MHAYH0c/-.^OFg\Z3Q9Z?BgB+Q@gGH6._a&dS-C/AL(I90]9I
E9X6c)>OE-1^fgbcDS,OG=T0:\9+5/R+_b29f<_TZBHO0,;FF\eb5WB)Ae6]H<02
7Hd56Ug;6?eQ;2gEH^[_#@FFU(W&(7:3H?^CcI:P@dOK<N/2DO<G+IggE&&NNV^-
1/G[eF5fC2D/9e=]M;T@CAeAf)Z<+N2Z(D]UQ&\G<R?7YW3+1[g/J)(SN)AN9MHI
]@(S<CQ=Ee[>VN0a^7GH>TW[FTdIMFbC<2XMf4_9XbFSWM1>@TT\@2E5Mc4LDN&2
6gMATgJa3I.,V=O8O,H?0Q5M5].ESc0fUMYe;A[VDPM3TW:c2E^>M-M>D;P=L_-A
.XMB)[(^\fgT#X7PB3c;+.aBIE3<D_YJYIb<^=cHPYR/Kd^.7;G9&RG.DQf(5@c,
B>G>S]U_/fUR#8:([<Ia.Le7S&7N.(16f/>;+WT7(V?UR4Yd0M[?)ANE=ef9=A>3
<bMN4QN;:ZR.7Y=<TSOND[M0[1CVZ96E&gAM8c=K=7S1HDVR(/>QgEg>G96/#N3W
0PKOXX??G(J+B\G1/M\+/<D6HNX4=(B=\61/MN>eWCee#49VJeNKV;.UP>@2c39(
(,NQd=Z(QP:-U>DL23D]_96#3OKIgQN0N2KOTUb6>BCGQ\(EGTbf0-V9a;@<_0aK
-BD:A&Se719e&Z6J/U6>BDQUHA/JHd[=P=MGI)8DLXIR<b.RgRV]S^_5SR&0AVEd
8bYFCg2aEce(0a7K+:2\T20@.T3b5Q>)>[3YH(2:g1J0WNUdO]1+TUBXO=LRF:\S
2<?gN^</Z=2D;YPbBEYW+\L7(gR3UMYQC-dHS[?E-Y^O+c6^KG#9DEg[\fD:NbS_
2.F5TUWC;)_:fCQ7(VZ0X+N19OQN6J]2-;_Y#eHV?4cTJ+-(1#:\Va;Q]FF3\T)F
\FfY?^^70[G54]2AF[/>AaNLfg<g,(W4CBDgAW^\Sd\A@0G:BN\7TcB2YI>?Q:<=
NL)_e^,^XaM]U<JeOE@5UU6g9[f,L\^c\1Qa?6U/6;]&dB(dcPOf6\Ze?&-XABF-
b5)f#8POR._WY7DB[40S:/I&9K7ZK:+S\E-945e?SP::1<,YG+=[.SRSO.V2(AO+
7_Cc51=A(dGef/VN\SAf,T:CeE>XbM[GS/VJ0_D;VC:(YI&1\V#)^.PAf02EK=:H
6SVGKH^3P[JHH>C2(#4BVF>5PDG.K2Tg?,2b>(,V\(OSH_Kccd;a<;Z0=1FcQ2NP
ABAfU=]OCe>ef->VY,OdM?^SJE.e:&0-\+gXHc75(SA3\4@=8cCBTSZD&J#N4R9D
0T&eFR#H+:JE5=2PFXN2/U?V#\)b]^FOLU47:4F+,T)QR4,W#R2\@I31S_86)=VO
=AYE_@YX.98GdKc9PP])(XS--3a\ea_UZ+QL,gF/9AccS:XEC6PfF3.Cf/ZY9gM_
\e864E7?4-^1DH(fY(OE@G29Y^7/?9WRd4\>UG&G.>1#.I]:ADf&@/^/Ne5(e6=@
Cg4WZ.SU2cV6@HK<.;TLFOOY,6>Gd6JZVS;#C9RVe#\P^Ne5[/\PD&//7(PW:,&W
H_2FaCcbUD6Y6B^SRY1HgXebJe.QE64OL9Ng2aDWe-\)^VN]H>PgN4(H#TB+6M#]
[Dg?C:K&(B@92WKD.2_H[IFDGC=47acA1KP,+)V483+KP=^:)VgVLJXQQ:0T5(TO
G3Cc6VNHL.>_BJBF6Q&,g6>QF6d\4P[=FTc1I\WZ^1PWdH/f_XHEMbF+@1=d]aNV
1WA\C^Vf2Yf8#caXI4_6N(>3E-&:]OP5>>?(:._1U((R:2.Vg:PFBVE,BX\;V@]Z
+CLA00^]E_DbHEJP_gFS/F]acbdF.C<H>/V/aIA9=G@W&3Z#=Na^/[70-,aL]Wg-
::4;(=ZXPS?+FW_(EAc?/^JBD]_<WCA]T:/L^-]_G40S5QUL=-cd4ec@TQITY(76
P6>4]6+R-4]LSWBMHcMgYJL2aBdL+HDgE72>;J?>H@G0T\L^/YRdIL),F)3_-DEa
Y<Gb+8LX^I[CN85&)QDH#U9Y53R=R(I+5)]I<N-QJ1SV^2SS;f;]bJd3/ZR8R4I&
N(&9IB9CV_\1]#)=BX]1/->e7:,QJZM^:)5VRY)b,W]#33^^CGNc7FA(;V>2Y[OI
Sed/G-&\Q<P\0PKbW2FPScWe@f1WQS;FR9IV[ITST7#+2bJRc<>a.5-9@b8CTTc9
g>YecB4F9WA]]E2,&IK6BD<=S#(N/99TCM,.K=Y@BX+C46\D&_gQRYIYI4XU[T<[
Ja3MFaBM#XK);?eMdE][A0FJK;=62S\/TM2FC\^E7EM.CVI\M]2-1e9,@]?(W-;Q
:=>3]47X<CJK(RB=I&A/D/;Y8\\R8JcZE=7fCN>T;A0D7V0aJ:fM,.MdITL1Xb:J
Td<MEEK+dOPBfG?4A_Z^aF-\CC^Va<.IaJ?^JTMfK,5>8)L/Ld]<I<9ge==[a4UJ
NC[LJBNS(=QE/e.ZL5.O.]D3=9GTbW_04cQc+6P/(5\YH#F[?gB5XOAd.J5^.@E]
C5WXK0g,Faa1./2-5&Z+Wa(Pg7],56-90N^-.0JdPB^_eKY4/G(Q>04B)\2eT@@f
[YIKWa_IVC<P.K/aC-.?RQC>;cMf7UTc(OBJ@4EOP[__N6e/g1e>,F&RN=8G0208
DSQ/Y_LZ\+OO\5eWDGH4LEUSeHV^Z<8c:#_/g1:/feKOK&RES?9&MW[TfKc##CcU
O91/<,EVNed&gU9KNaO720]MD#3^=7D6J9a/VTbH;^^Bc,:=BZ3b6a.D;KPQ?,5<
?0e>]X/L0C_g7.@LBXD6^.LH\5MCZ0QUM^a9COeP;V872c-C\NA]T>-,C/Z(Q_VW
47_23EQ\HPUEgC#YbOFa][ESZ(.4((?XgUHRCM6R49NDU)+0/[NG2(;(.^Z1Q:.Y
W?M.fGbF>6AD-#bHA;^<_#+Rb7CCPN/Q_TW+ZROVc4HdV)?YRXTQW]O]>C]W1db4
V&R_,dBT<COc)K3<LN1_NL24MH@][Q@aBA+7_I>3]c7R0XX/[>YC?ULACAf2SE#]
CA1.5C]C\0A\>L[HP[ge9THPAXY&10239TQGO[@8[a9@&T<[:5_)3UXQX0^Z7#HY
3OQ6\L7I8\<;Y,_fFR:DH,<8Q_VJ5S?<<T,:R_?=W?:7N6B6bH0&dU3g(-A9K<^X
@<f&8KV[M9##+dec^K<>Y2L[UW;HS0[Ua_C(I?@M.JEg2VPac]VX7J:be3R2D;1=
W[Q5U]fVW[2&3aAOd,f@0ZRdMcDgUKO\_M4W8d/9g:09::,eN,EbaeNG;BLW48=0
9OZ::eKW3eKMbHc-MGd(EBRE-H71RY_[V1aC>U=5A)Kb64Td_=6J\VNRU;A(e+c\
<)T\HNZ-,aH1)e0+6?SLY&Tf7#XU@d9JR5DTI&<^QOZR=3@aC>JUAP-7g^fJaTaC
RT6ag0?L[Db@,+QOYSJ&]L6<W&6>M<=WMJ:a@MfI(gK4f=37gY=g6UM1FF0:F0fW
#8,ebSd^LE7G:SbM^L.-+08MVU(C&;1LQ]g#?HeV:^Z;T9WfG.-@_Fa>;/=IV0K1
4b0[/;#@Fa\:AdRR2,.#&:9&>&<cK>:REM#(#S/[3DFQU9/>/J>:fR98=)E>c=:a
,H20ZTIF@7/(@Z=JHbD-<e_G2YI<)(QgN(ZaFegWdaDfE4#(ZRB=>bWe)I/>#XTa
QND+(<L.R_HMeYBM>[IJGIT4Y(9DC9^S6=0Vc?6e-Q1_1P,CI9I5P/QNR0(a?>1#
-Zc2JMH]_d+N.#Wc#ZY0QN,fDB\CHMV8[HCDKcK7WMag-BEKSMN4>9AKg=<\7eQB
,J6]3R2c-)U#bSMLf8(97J>>.V]Y/.Q,MNWR)^?A2N&YJB0g7[?J8gf7P;?(Ia@F
.?E6.GW_=R-,(G.65N\F#@_A_^U,:PB6Pfb-3)DEVdU-X^??\#d_?&RScH>GaE86
H?4H^JDS-[C0H=;M\_=R?+0f@/?HRZ#GW^^Yd5=Y1S(bB1=gdHI,f.Kd>TOFQ&+<
33HKG+A7R9^_De04,>?=XAV9ODMQ.X;HBA+,:RRed/TZSY.14BI]FWV]=HB)L-0W
Q@;SPb#2B#XA2:Y.Df9&,<@;bM).SVD8H-8Tb:W=V\RE[18P2D4TX?,)O:XB5ZO2
:aHY0_F<\5BD)\\IKYD>WLEPTWGgS455V_8RJ?I^CR3R9->/O/)5\:L06]Z3]-S?
IR1AG0<;/(9;d9BMdKgP1X5DF-<MZMPg20TTb@I=Rd:84P7eaTKP(IMQV:OFE1_N
NL0-N3F2\D;J,.^E>R7G4Q=JOb.AV#Sd4V[dPX&Qd7g4?/V)APJbZ]>3_WT-&=[)
=:>eZ]JLU??b.FA[@OZP^XIN<M,0Y5g4I[,C0WS_f_K2G?H9SF2[W7V5=EU,</[P
MTc=8RUH0H9WT&0#JFS+8DfKM5/+BIIf7>7Q4?B^T+)?OfA<K)TOU5CLX\+76/aN
@V3ZEI4U=Tc\Y<Qa;d4E>&(Jc.^0HC3d7A;;6FL>V7U84KL(DbNFI=QB[8g_9f_Q
H),+>01JV@#/57LQ6/,AK#:9Xb@]X+HZCVY\2(f;-JF,0[B#b5.<;/OdF+f>EdRA
.6<,.<1#5ScSXJWR<D@:AQ^e=b)NV(3D0(D\[WKbEK6OOL>Q[)/.SESCYPLD,aT]
M7E;UL<9,#)Gc[K95N.5bUCQK>?2^dZTT[-&32HU&cCE_\<e,c0(ZaAdOYP#\:.<
6C;7Z-8/Bag59NPeY50J(#cad^VPefXW&/+GUBXNOL8SV]GNKZ-AI)c3]KW/8/X=
[N.8,X+BM-eg4Y#Y=S:a]\C&1YJ<XMVW4W[Pfb6eO@d7]dS?[fI^,W3U2,];7[CL
9>ESfF^YIR1b3EM7XZP_=,OQY7Qg2A>+Cfa^@,e,,6FHQ^XY=7Td\D1J=:HMC@HM
T7QgZN/4=(eLUOUB<d&P,#dS/fS<cWS#/GH,B1L]#7Q7bcLc7#0YL@MI:GK+VF&J
PKWA?dKc[=QE\,;Tf5Y,eb_ZePU4O-W6a\-6c<6fgWK&@[11V0A9@&g),SbRPDJe
_B>JeO3RG)JGIN=7Y)7:JZ;7XMbX@Z]24TO?2AT0.:Xe@;MBLUbRV(1e?^NbWF&Y
J2fCHEKac?Da8M_96^dOCFFP5,)JZ#Ra7>2N_U\;=S2Kf&Df9]3G2d#,,#@_c#VZ
KfO3adCPY-COZ-;5Z+=0EK-MU8WN.<3K1=)]E8J5Yd4LYe++)3(5/aZ:#XO+]E]Q
M/];6BO::JfgN4V)^H2IH4J[,.\&W:S\4588cZ;bM6F/U\HH+)83P?I;E^e44WT^
\HLG[X<?9#=eK:N(&7T79HeSZa1)&:Y<d3RDJeDa(W)d^HTHQ]]DUZ[WaRC#gW>Q
O<cJ=dI(B6)ZM9g?&A:-P=(5OA87#V1<:6b@cWD[Hd-\-IKcKB/UWIUDR[F36-W\
89]K@a;EIg(b:;D0A^X>\]^M-HYC2fPfM^;D2U/J)QU@\ADcQ6EVFHT.M7C?e?#H
4cM@Mf9VJ->IJ95,(bNE.?U7.NQfB:BS/^e0KU[KF(/E?WA7+YI_cQQ&b9[;;WOP
JcIURLQZG8G,OPA&R4^=^4]&<T,.6gM2TJ,/10.QA<.f2Jd2e>H#@2]\TXOB;cP8
e(@6HIDHW1_OeWS@]9A&PO<P?5&R.be;c0\^ZCJ/B--&X=3.PBa^^3([F.,agTf<
7I]?P)-Og85aM^cOR(5CCLV\HYJc.J;<S+[1\#9]-@cIe1+AMU#AYA38cB@P3)Kc
_O[GXeKAZBG(:BCMZD=#\>9VYB]T9:)5YXN\3KJH=]1__&B;,I1:C85BEaH#B@;=
3^61IJU(.EcQ5Y=BA)93[P(#6]\LYg6#7;P[,[Y_;:\]UCJX#D0ZSU;d.NI36LA?
A5IQBCRddQ4a6?MB)7LB?F[19D5(\dSF_&,0PP09V[6T.aULbL20-39[R9.MR<_6
N0eca/b=M44+;J9.:/+LSb9<K2ZS\3\SF[(3?&(-_\#-&&I/N85&@f)[Q&(ZR&,8
bDVP#;;d/(:G9,(WP&@Ef+ZMfEcTQ[<:/)e=MPV;05G2)bF1_Hc=Za+>7BGfD,]A
\G,\=DZEBC1]P(D;[U.77:&WOC_aI\)P-X93H4GP.(5B\f2,I.-TI#X4QE(60]8A
?B0JW20?bO[M]);:N(fRZ))GS,A51DFgL>Z;.9T>NH]\g(/ZU,A;G?KeS+0Tg=&<
A\N?eA=K&QN?7@&R75>E^2(D<79R&O7JQ^Z9B][UWH\\;@OZTJ(/=XOgMdX\>3O9
,7=IbF.DPA5dXb]B8B>Be7(Rga2)=^/+3d-g\SHTQ3^[a@)WZD0^7C_?U^GZP=.Z
3D]8aY]J310)3;Z-&MUfRQe:_#/(X44AJ)7S=#7[9#\-7F./9[d?N;834E>41>-2
c?Wc>C=QJ^_QIeD79P^Y5444g0&=(S5)>HR;[=:8fUFXDXZ5)IbVGZ7HWO<3QBNX
L>^CL>0fO2>)XgZE&0d:S2f)6U.C:M/^IWZIHg_:_]6g2eM1U(9B[O5I)/E>T=Q3
gb\@Ma.M4F>,YF(8&[3#@#+cJ:2H,]^MWC@K9=ZeCF2?[#,;>92K-KY6HT,74XY@
\PW14-8gCWRDgZRa(I2\_)OHURMX:WO.I:)S3<849Pd>\ZJL9<6cW)g4#-TU<D91
_7Og5MG)#G.:3+::^#,C@gaEUa,9ISC.J2GPSVC;FIT#&4#?A337S#XQ11P9La3#
8<F+]P8M7OSNSU?ZXH82TE-QH.7/X2B.OeFT9A@Y[7aSH@ZJE&&&#8?K0L9DX#</
0TMH?#3[WdGdF5:Dc@]>a62J\Y]?1:c+VD@^Y3Y0f>H&C:8@QN:1\D2U:YAdSM6Y
W1J1#dRQ,YAZ/B1>2aLVZ.W+W1U:0810?YLU4M9GZ#.2,R1>5ONJb9)N3fQRIPaM
4;&cZS/;g1T#IT9f[HP:AQS[)EE9?aMCd^c-XTcg8II\LZ994]_X05a10C:QXdC-
?U=@,HCL>eZcRJ8K2,LO-<VBfG>3L0IPS5e?VQ/>#:6/B=_IQ3C_+-(_<2aA)<ZW
=KCHK1;M.)F1&WL/cZG]W=P6O\0@&\5#GMV7>R_G]U2aD]/EI[Z;/IOG1dDN,\^N
a&M[6Y]QBICZ,N<bO86\;&1>:4ZX;IXCf]K9ME8GK?^?,<ONT9KQV9Q>W7D?UO;/
c6Y0?b\D>#M3GJZY-K(&^?9.)MT23[3IO?SfXB&Y=(ES/,/^cFeF3\g)R5\1D)N3
&EE?DC7dG<ObZ7W_<JUH#Bbb)JP11VZ?6=Y(SO(>^3dFb^7#Y<F8HME0L@\(>,EW
?f4TSR\Z]GM#.8VU#>@/29U<\81TZU2cXBN.E)9OG&.e.#1WK;5;))[625O]NMCe
YD.(YPK\\=_?\,XC(^c^(gS0I4CH@5cW:T@):@NC=^2LBUT7OS0PDQGUY8N)FH6&
K<>\dQV(Y9>:cQf#HGA<_.W56+357/X0_N>&eO<IDE+1>H.]]?#@IBD-R<[LMFI)
#6L>>bL/dIHX_?5RD?e;Z),MgWa?g6-K^H,A-LXIZdf]WZf20-g,K#XT;T/GJHOK
F>W[[OQ&<3J=EN?53CaA8BN@8@0=B6Q0/SM:38?IS;,<fedP:OgB==GS)/P&D4F<
>3+_)gM8RC;DA)+^[+.:1BUdF\27e<@UIOg7Va6&2WSA8+2.>,;UWdHRUZM>1+6<
c_=g@.OVHVVZ7O/Oa?IEN)[bZJD)<S>b@J0,.1]<,)OJd4JM^;5K>HQNJade:OWT
;9Qe?5=Tga?H=\I?T)B[?bc<@-B1Pg@0K6^4We+7,/VI17]0EfI.K;SG/@GL\@B1
&-g/5#JB<0DMbY/bPee_8cGU<W[UCE8C=;24bW)GFTd_BO:MV&Xd5+G8R>HRS]J_
1CRIIgVQ809LFEE^E<^7,LR^gY&9C5a#E8I(O_\IWON?.N<5Ge6=#.b;+<EEEBS3
@6DU1_9KD]V>0.8P;FMC[(^,DgOD-J\&/ZKZQ>/573Le][a^7,Y>-S-K,W8Ve0:/
IQ#@BVL#A:_]bcbKe9\38GD:+19,[R(gd30:QMaRb/+<T3>2eg-bA[X;B;WMT1d-
ZM;83FTMaF.\1WFaDK>Rb/-;8>HHJQ,>#GZ@+^7_@=70@HMSCC_@aWS5Mb7202<I
HSg9Y#GUK7<S=(IYIXEd8_b(6,D1bb)-BN3a;79IP8\MJc<N4C_14aA0XQcQUANZ
N.g\D4/M>IDJ39U@Of\M]/PeWWE+0=29(?+EVbL-92_H4#H.c:F_eR[7/M#1_BGC
gT0UF8b,]8PKULJ4SR<9e@CHdWQIKg\I,<SDcTeGg2#:C-G.-Y)/SX=(1aLRT5_?
@&^Rb,\#PYe-RKQ/Y0EC0KK(\ZQf<Rb6XdT^Ta:3bI8,6X9UV3<ND>?&JQ&4_\cJ
90Z&1BSWN)O[CMbL8SJc[Tf4EQL5A#A@]_=OG7:#2\.^b9=TAc\-_64,ebV6&;dT
?+S2L66>K&I_.&H;faff:3W?;7d1X_3CZbMD0V@VgBHEIg5J3)977Y>\\/#g1<KA
bQ?f<SLN8GZe6V.-Z([-U<JIW1\H[M>+d7<8BTEfN.G=?DM^]Z;0_O@](WLQ?DBU
/XI(4OFQ^/90ZKEg=O6#6RT>R&6ZgW@b_&Cg=LeP^=Q@/A?K,cN;5Y9L87LZ6660
;7]]\?D?:[0N9(f046:GLeFIJFTa)U--.GF625TJ6K,K;cF^PgF^QVRCA.[:)e^J
9Bc>I]4e+Q[-?DaPY2=D&WQ=E<9H^SQ=)<S1L5<IMU:PHEB&TOB(,LC9@SLL)L4,
C4+Lf9Z0Tb7#P@Z<77abMY5ZMT.V0?&(GN]E3HB;OcW/If[8O\C>ZO]-<5ZTLB#g
,NMWB6d7P-d...+7L5dY^>.^>:-3Z<RS?O=aK-GbXQB3)#DEK4Ue8W\P]Q,#d<)5
9fKb6VHC&IQbEA.dM_0U[KfgH9:L+G<I#+g)D[X^O\W[[5eCP;B^N4O6;7Q,(Lb[
a;C4DY&B46DS/9&F=Y5b\7-GW7>A,^-NO\;egAO=3UQ#7e[TND)>De&.H(e)Tgbd
C<>:,_+[_MV77^g?#g,T^CdYd)\eNXYeMS:.]g,4D4Pbc/g5TOgSWC^A_;5+K3]5
(0A&=;0XQ8_I+/71E#f5gf_<)-3,E<9FfU61-JVODMSE[4@:#J99M8OFEcEe#5V@
bWOc2.9e),)dY+/=K^41g/U3\aY=eHJ<B_Qaf#bRb7La6\U_L_.XMNNALKOVHe3^
7O^_AYB(:T;a=DV6X[1&VcGTd-/+CT)BXD^0=e-/bN?:I:),Q.0?]L[e93WFccV.
,^3cK-6:Lc\Y5)+0?U]ed6T+E[7^-/X86gf.R9V.KQC[MdA?S_#N=()1H8JPO6Sd
?X:7VWJg^X-I3(>FKM(_MH,f^OOYZK23-<G]NE9/E=?c>KL?O>G57?),ZDXGXG)^
+J0A0.1>>8U4F)3+D6NTXSCUV@(/aQ-IfW_L(II)/gFD6a6?\L0dRD#c7NaY^E(P
?XIX#?HWVf]KCL9QE3XGG9TP&5J^.Q#ebZ=YT2c8aDd,+5S1U98gbK6V&1=bI53#
G#2H])=?K].]e6=ed)W?7?+fA(:,WTBT6]Ag@=0V^)NO]C])>.<_F4Kb.,TI;M2=
611g16()68P;QQ:_e(g3V.@:M3N27?WXQS^/WT7/#90;^14G@8dU^GV@&SF7;I80
a+7ceeD.X^_HM,]4a7+gHU7(F/f[QVdC1X1NdVF_H80gb)RWJ6@9VKG66J?NUb&3
@EPH;;#:;LRI<7[[>OV;<(4TA&>;a^;_7K7beX\AC:D?Ded9b4HV\DTG_MfLc\&T
,DRLZECJaNcMg(6HP\5aTXMfYPgJPQZ4=J-_&O3A^=R=]8P)(:XE0DM;TQ1e<\)O
L5G6[\U>]I8)@IYAE890;JBGAS(G089bETLX0W(NU8QebEA40.GS1M\K,3XCa>FA
aTKX&LJc.?cY+EPGV+\:(QS,WZ18L4;_/Z/UcY3Tf#e:3+[RJV40U8QCY#.0)1A#
[:+R5+J>(T>dYAa,>0eXg&>B)dSbbJ\cU>3I3RBP,65a]L;MfO)T0,,\<Ea/dT4X
BdB6F(?6+9<C>YWR1g2J](2)/+e-X?=<AZ[H?_FP>e^5L>c#c0]JcY3<T6F6IMV+
gZ77G<LEI?@7?\V[,0D18Y;6]F0gNI5RV=0,A>TAfLccNI?[RGFA[gJ;Q(B7#4&g
TZ8LIa@1aN84>H8MTK9:-YaM;U-9gH]@(g>+LB\>-HM>f],72#ZW3>Dd4U=9[2Y?
BWgSdKc0+.0eTJ?d_BA0(A<Xe<;(I.HI&?dXF6WKVBD;1F9G;&?Q8WA]A=/<HF:0
-@QWKCcKKAZIO<@BbcGQV&-=YLc<:)0fW8&FX^>>1VC\A591=0\M.N+LCX+,=6.b
_Nd8>>^.WVR17:[GOEJKI;:@4?QFJW_b2gC,D+?U\59<Y+V-/UU7\#J;.@M?T9)Z
6=+/;R]FTUY&Pa?V0F86(X9S9PKLK#S)cRE-D6_5+(A5d4ffT5]^VM/QX[/gPCBV
>:1^6_bQA;3V2=>GL8SQWS[:?.53Cef@OT2H4KP:#NG]_3+_N)D6F_C_cYbKcbI)
1UGA@N(O9;>X93.H5L?92cUgT@7@=<N3O=f.^R[e^\>0K42K++]<?\,V=1:5eS?0
<2F8HO<JJ7/UZK5H\Q5YNZ\SXOgU@g=4HZJ[/U=##TeHEdU4^:ZFM4GKFYQ\)5S4
_T^D#\^NHBd77>e+,KQZG/6[U(GB9Tcd0?eeD4-\SAS:CB22;<M)_bc@@MNM=ePN
;d6XOg(Y03FW4:8J:KL6\C+0;g?[VOa(ISROQ@<7;S34;_NF0MdKTQ5J[H.X;F1F
MC(^+ZMb<8S-ST@WVd(V6A_RA:>=8Ae5)77JD\?<ATLV(]?#KRO4/EM_,ZVSeG6_
76,9^\C.P?[8]TgVYGDQc]QR3U,5AaO#-8;Z9KRPP?:9[Gf_-EM]05:AP&V+GL+?
4.CRQ1]X@MDBF-9e>EL)Ge+)a3eJ:S18FfOLD.A_T.\PcE\65ff8gFQ3M+RTYQB1
^;(O1>eAV+.=Q1E;)4.K1bb#P;1/UH2e,3+@#,JULc/gd:+HYW=GWgL>I\+0\9@G
BPTR6<11T=((4eS/:[Y-Dc9?\T5c,Ua4/Aba157+Rd,1Id?XKUbCE=YaNO2\>9JF
X)71@9+X0T<CL_=?BCSU<FUN0XC0J)]MFdcTTR,V;EcHU\-O0.,#BD?I)U;2a?B8
J]5&dQEe@K439KQ,\HYO\EOOYK6)DfR^agMVB2SPONY;]4/]B4OFVDYL_@H:b#1)
e,:TIT/^Q/O(AU=dSM:R[/Fd_]4d=NG7_c:b.N#gZbD.TYTAZ]@H&YL2OEP5fcOd
O6IaR=@A-QUE]_T#DLc6W597(1E3A3-A?GT)T2HdR2#KJ+Tgd2SLNP0f0988>Y&4
^MM2fPU2^bNDM^_+)c:>+:MJQZN6L>K:,9d(Q79eQ/X0P4DC:>89\WIJ]W4\6O5,
5:/8WHP#]185eF8CS:[]HM9fBG]YDAd\];c:UJ]7ab-^7E^JUOZeD_B,./=.GdBE
Ab_^3^9U2Hf3:/;4XbR>V8<,=4d6P>4=ffD.M5+f:,BYb\P_=e4.;G+/:\.a=ZRS
=>.YD2HbH]<1-3J.GPC+C.H@[-bQOY--fBJ6-AWAZI0OGM<dY;.URSELbR3TOgdE
>da4f)?_4K5+--)^]AM+G.Ne:dPH;89D<[CA-HA=F=[&U[3Uf?>3F]&@-dUKUe3-
_6.VfJc2_CbBL[LTgdYA]egT2]WHN6,#^?)dT1-?&dIO)A5c,]/#a7]=3:)a:-LT
FHKcdLRQIObJ-J?Y)#7[=Te6S]9^^0OZ+f1&fOf<bSGT_e]DKW]\^Ed</bC=8NN9
5bF;MKZ=P[c.RDcCcWc#R54Cc0LDS5))__VQ#A23FM>C4C0[SbRV61g)=5(3W5H+
:ZQ2ROA-C[GdgZHD;8T3K(_SDQ;fK^g68TDeD_P)U.=6AX.Q?E\e0-2bF(6^)3e6
,^K5L9b_Z2Fba[=4P#Jf.b/[30/)@(H_UII+E@;e33G^)\)X01G.f^Ca_bO@K>fI
I=??IUT]55^1K2P\91(1AU2@AYgO2IATd5E/VWde=^Q>J(9#?^KDH-Mf)2_OZ8fN
6_QH?TNUY9I7)L)@PF^a:VadY=<9VbMI=6Z+0;8GAI.gP(7&86OeW)?bd2F]O=0Z
g./R;c[PVTON\]IOFLNJV1@<a\_;S):U-D2XW:ANXL9I(#=E8Fg>V#:#&U0K@gJ6
>cN1T^QJcFXBGbRYJM4NRL7BENI;0WNX1X9XSgGJ])7UceDe[G(g7#3D[Ae/7G?#
+EK&V=H)]7U8>CX(),JI[R9TB13:YQ;PNO:^S\T&C^:P16<5^Yc3_RA;2J3#O)FK
R)cW@cYIb8N6/I<RFX<5/&T2+//OZ4L8X[E>&cYNOP=g0U:>42:Y0+OQUK5MK;NU
S]RJ4(B-LKIg;V0CN]SIM,ZR\W\Ya69/4,T7B6#[bfNUb3#aIADZVMT17KJ]QS<A
OD9>UA8[C([\#.,HJC]6J3KQgDMFFMA(e@R-G;_7FI&=1PT2dOdI3KW:C^J[dM1b
eRR#K#5OQP(Qb+/PF68[L+bW_9XX4NO]J>^EZfCK:L.?9416>cE+AD,/2@RdUJSB
=<,Ug83V_55.2MKOT&H-D&KM7Ae+bUfL,-Qb:2Q#;?.9\/dd>IQ;)>AZF>M/IeW]
^ZO79F:2BI#.;I9W?aEc4_KMAC38P;>D/bae7=&.fB6E<Gg)ZV1ZG]<R9eNF.d,g
\4L9_=_3_KNC)a3NYO:1&HeO_9&@J)6XJ.Q\4=/<Mg=\7RIYS6_-EQAfeYA5P>:E
fXP)39ZRZNIW3Z1^=F=D@Q#+D:54dMc-Y)>B_@L@:6cc[daN_HT_9Db+[;>c8?Y0
3_5H46Uc:8KUe922.&^_Z)_P<;.O/#4V]00CE[3BSZ?7S?b6;2Ua=#GM1<@cNNMS
EZ,A17Oc?5Y#V_eMXOc>T=<ZUGeg74?R]8f&I>#0GOG5b_02,.W=SF]ZC=AgMDM3
_I+3Q_5(</gbM@A>A>>71XKeK^gT)OH7aWW[5CCbY\>O9+29RX94KMKT#b]d_eQ_
L6B(O:FR8LO(eM4+=eE38V<;,UZA8e_c1QW[@#a6D0FAc@HDW8BJ@T0^N]?:+DW&
-LEK2);(C85W))FL2V2R=-@;77J6S=Y(NSL/CQ69=5d,f6-_DZQ9X)I\gJ.C/7@d
?ZD=Z:EK55C8U>#/ObR>:#?(K4W0R#D)NeU)SDEB-<V=bE?C6YSIf+7>CNgF:b+f
1JX]Y9168R_1G[_7YWUc#AHgT<D+cd_2^QL=A47KdAbCg,4AY:?0_A_>Xe5<bVL:
LF>;Mc;O_cgVF;OTcGK4(?V5)5[&N/cfX<2LF]fYWT/31&\a;+Xc7V<N[HMY[CNU
^\BZK3]#^\&PM^aUe>3]9NH08aR.^TS#0a&4>3.,2)1eHZ(3Vd=ABNIce9_c40bT
[TbUb+\3X=,,G:(Z9/UZK2I45V.G3C##:Q[5\BU7UEKR6_]A))RS8fN9OH<L17-?
bUNZ6^Hb-S:_XCbSc?e4g>E48GZQ80#F-ObcIb-]#?@.U-=EJ3##9<_]\I8D_7J2
RXKJ7b9DYZKNcO6\4f1T@,M3fJ+:\+S]fK)&bZP>A7bJ3J4eE05@OK\&3d&be4_9
-L2@,eDJ-R06TQLKeJSY,JKDI8C-=d,^&(YP(AQ4Z(+;-e\,L1Q:O&B>FfWSH(A.
,@.M7S=<TD:N;UX8D)=D#4/K6QVZ]1NZ(-U=G.^S?P5D7/K)9B@g+VQOJ&ad^\X@
7\@CQ1UDRIb1IL17J:V(_V,Q.-d4#4C@51Q3FLUUYUNDacR)>U+>,MN?:R[14:4G
2dJ8KN:XeY-;9-=YI<Sf7M)M@dZ1=GN_IPCG/g1J)MQEFXTKSG5d>BNBT,1K1YeV
_S?W/J+LSUS\)@&>KXVd,#<7M#Z>a?ZKO^UP^(/I&T]A1^-3(Y@:H;f9RVUXHGN[
bCIaZeK]E>BQ67I^__Eb9<_PP_aT/Y+GA@1Yc;U^I(b8Nc-FaF+<R40#BKf^+&2a
\3C_Q8]8@?AROKIQI@\G.8\)[QWTB0a=R&bWR-P1(=,94R=d<1^9=fWaL[PcW6[A
<0F:(0O=09H/]GU-/FE?H+bXf7KYL>I<F,-C8[P^/^&NOE9<LUYX;#TBZXQ#F&E4
cdO.?DKd7fV5eE9R21,@&a_6U#8&Zb)WJ(Q>fL@Qg\KNLO?-L\a(ER&WU3TB&/):
O)E.99WD53W9Z)YQM3Na3_)-Y^Fg86eAe4a?_RT6\9Z<B77XX3N:#>_:bS<-^HFR
\bP86YF3M-PX_dT7Fb#M62WN=,9@MGW@YO96aA;\E=OT]#KA^K./K@Y=7TN)=5WT
CL>Ra,<G>12CLe[07,b<MLRY\-/gOe31I(2N)0,:H1:FI:IO9V:F.0E)9&M36VI.
8AS0+A=>Ib(ZSWb&MVAYD_-7/bML1K346/DPZ?M9f6UNONFF07PXR,@Y84IOP&L?
5W,N:d&3L[=4/()+1>FW#3-):30MHC&9#:Ya>c=#HNFgcHe(M(7RaeMd@_1d^5XF
]YIG6/;8F6ZJg^B4.&OEEPQM+Ze8@0#T:YeSV.+:UWWY2[&aA;BNb>cK,Q0BA2dJ
ANJWg27e6D]X4b5R;C_A?22WO8.[H53F,5a.cEf5,XBU@<2SDcVT3HUNeb6[PQ;D
EPQ0QET4>H@1?;UPB^D<IaFDA:__]^#d9]N:G05cA?Y/I9[X52.F+^LS#U=ZI>b-
(Wb&;HNa8:KWIXEA7,/,EMBdPTb7b94/@Gf#6Y?TDd58agZg8FU2?Y5Lbg-&SC=Q
Z-g#>.QK>DE#_7f?3?b/dCE=SQEKALfBFPg=3E6#BEc\_^.@Q]dWB668+@ECY@D#
fS,:2Ge<c>FRZZ9@=KMQ>AO1)A=EXH5;,/J6WDcV\371XGgc[]EYC>54/(Jd#bE@
aD>#Y=/;AW_=M#Y:;>7Pe^V,dBFY9:@.?4U<LW3TP+3eg0@ZP.M1)2ROcX#ZDN)S
dNMTP<]?NZ4=f+A<[XWQ)O2D@ecDg&]OT1>ZX)c^;/1]7;UQ\6eNC[Q>bEPf\3[;
TJd\PYZQPf0f=-EQ5g.\HT8;1VA)a,=Ka>?W:gc#JPA;L;_]CO7PUQ^8.48:d75V
]]A.bNU-dAL9P&I-Z&2)COE-+VNR9AK]<S#O>KN4CP(=I7=e-f<Q3eDB\.c0_dZU
5-V?[6]1S7JK/YJ<1S9Gc5CAEDFgWg6-a8L826::JM)8K&YSN@QQ4P<LP.^@2@NN
f/Z<Q;(=-:(3V[\6B70T;3gBc>/+M;L;Cb[B-X_T,Bb&:V6(IA(DL9<]X/7@>,Ud
9GdET<8#eB1>RD3YS;N/g-\g^J>7BW9BgP(_M<cN=[H#D.=a#6S@VC)(aCN\O.<7
@.1,=gdK>&V.?XI2+8BJL@f@T-Y6&C6-4LN=W3D)9B.4A_SI9VU]E/U=Z-BF4Q=)
bXSIX<YPKCCcRJbH<0:?d9a6W,bV--IcVI)4=K;:[#XMJT</#cfC-33^>DZ0<e:0
gC@H.L.<B-N>Lc)=I?/@E9,O+4b6H9HaNGV88baf&\V)YW8AABO?GUegL7C3,F(+
aS[QBLU:_c.<_Od8PSN\-CNgSBg@4GC?=.dZ,UZ&W#(0X;IAT4NL[9Q1>1XLWdDe
3Q;@PKXR^PbSYPL=1OY9)B(<F#TJ;,@0+HLC39S;GR//HE7_HOL>(Y889gUU_6SB
0(-N6R0VU1Mga\#4g,OJ;Q:g\.Y8G]NH^C((Q[a2U>g/KYK_;^&LUCW?Df4CFK?^
/Td2N,K<B.-B7(B7)58-V4\7SB-W@U7N<[Ygd_E)5=dc\G;BLB(cRKW4LM(./7[-
L86B--=_O7DY[S4W)UY(^UVWCC5(UUM>dAb>C0]J#KFW&7UNM\T3PBS\\_<#5U)]
LUO\;eGV,NDcY0,9U9K3P7HKDGQYV=(AKF)6K]VB/@N/F4KeC6P(5.ER;X[:(aD:
eO59:Lc3g]5fbW#]]MgGTe/WIR6FbKgEfB4C7^(^Q.47\T)1g#E@-@&K6)(G/1f<
e4FgfbSf]&@g@8K):11>eUJBC(ZY_Z;FH(_U6:/J@.]d:1)#LdM[SMg5B.Bb@;_Z
A\,[P>K[Wc@b_GWDXJI4<B2IC2[.4[KF&0VH09<6@+<e];;S8ggNE+&=37+__L5-
J;(@-(=?c7?SFS.?)B5)&L_gCQO9/B[Ge=@]OV.EI:/_BaPJ24fLP]<=QB:^bY;:
)^F_8?IE:(B7I//+;SfRbCS,HY(M0?7HI;da.\a^8?Z1;-+_g#N7B-0TA]K+.:H3
\/RZa<Sa=+,YgKCd,T60Dcg2W:U>b&;GN9@PY;9<ddW-L@)-(PcYMY<<-.T4JMaf
GOWfZQRC&M#MK)Q&FW\GO)R0XP3JN\aLWF-^R<VZ9Ng1^Y/?.M>]8G[\2W>A.6A8
L]f06H>XK+4#I\I=#+,]#7P-g^M3Z7Q;DfZK/I:f]]H8A-<WQO&5ER7VD<g8T4B@
fYV\V02H5;O8P6_7\CgR:A\aBf#/5W;/JX<]<A(DV]&g#F:Q?J:)+RGf&\K_N<UH
)3V?5:O8Z(.b\&_R3X-M5_3bN61ff_<B7;JH^X7c#SFJ#Q+\-a^@?XaZHF?aQ.=(
VO/L;L?9TND\IeJUY.Q^TScRdJRP8VG_gfaCdE^9(dF(KFY;R02E>/&G(H)MH]/4
=>KDC&M?1RS4;6,RfTSKC_/9C]TNBJeHLU0>?-9Yg)ND,LF>6T4/eIPQH96LFaDM
_@c8GMF;ZOX&6Aa+/QQ5K_;XQScbE\f]]UV+9K)I/)RTOUVB&:;d.P;)GFMM1+f/
E+ND#G:R=9baL&5fTJ_N;5OS/I<B5#>Q37SOJ-@8?6ZWUfQd=<8f]KZ,A9)0C,_9
Cfe@[aY/,_5+6V=OMF/VM+XgU_[KBPDVeOKT:S2PC;0UHa)W1;ZTK.3QYM7W_5;N
^&J&J+);1=?\N?L&eS-6We=E[E(QXK<YMJNg\cTGe[-f;L4K5eg/+R_NF[S[[5cZ
E/Db;IMF_5Bd31ETd,RA:13VBN0<DAAaA_eaU/D6(P;792Eae)36X.^RU;SL:N@F
Rb(/>X4:RBfD2=S@671:Q,OT3]VN4JQ83Q,Cg1K[7<H]QeeVPDJDI3e/=QeV3S?]
]@)UJa=gBY_D.1XOGWO>(X[PaacH=#RQ[?E6Te?6R?TA6VYEW(E4K00)R+FgKR9-
Q^KG9C^\1V[C?eaCC4Uc\(OXWEC.8]YE/XG3GFD/eW;KFBM9EI1c&C9I,>AE^U[D
4[H&,/^K(\WJ>-D_+G]-c>C^\R&<e8:4f6Je/,H7HK-]1Z0Yf2&3^N(-cI_6W8CN
HGSf25(&4RT?e1<S787FCE6aLfR.S>eGL<VJ8^1_@E]_YgQf[>),Z-_dWF\6>,3_
:.?#I+\YFA53V<SM2;e:K=.afFT06^[4fPT73g;7D3ca&agf0b@D>14O?9N(IeC+
^40aU=YIab@[WF(R,f_R2VSO[f(VG1<(7X.ebIBYdQacM(4&[2Z4/G]+TN>OTd,C
5>C_:(0R\+BSCX<^0IGAg^&#;G-A8[^d^bR<]MDY89B>F5MZa2A0,eL-2Y@^V^YW
&]9a9;1B(]6PH3de4V=HK[M;c59P;NR)E6?46-dfL20bXPWL)]5)I&F/EQ_adC.E
I((\9FaF-bGEW8J56E&>ETE(T&3#S6PQ,Ue>((=MYW;b]f;5g8WP3Y.LV0.5Df[6
K><&4a8WaU_ZI\C3&(+8C_5#+PTK2+JIb]e&PA0(O:F,\+E[\f63Y?NW5._aU#J,
ATGgA?[3Z;XX]f;]81[ZRF^LUX7(U;3K<f5[)gH+,M=(AC(T3-Ig_U=AHVKZW_IT
N;bVOBEYR@X=(RSU0@(W^U0[b#W_S-C/N&@/:K<OA;_(77S@K/O<L]7\.>)fgLJ_
OIQPWD>W[O=0ZV.g.^C7<;89geEDdIH9/0/T,G6#8Ff:62)G=WW[17MZIIe[aPf.
LPg[C6^?gR[@:,5O9N=bYW4SZ4V=)O#>A3C:]D9B1U>)R[Y:M\(()[I]c-DN>HVd
+2JcNCEMFE4/SP&F9bF\_eRF(#RFH7&Y9gd8?9-[]Gb]EJfC-B/9P0?451K6Qf2:
ASR,a;0\6bYO)/9fM<R[faG9-;4.WH&2>_D0TGR<[SWUb@]@=B+-51De1)7ZO5TE
RLQ/+R_GH+IY\_?&ZGc[Q=8eR8X6/O/K[?b@g0?M[P(Q4HFBEWPea3O-#?.T1X1O
5X6<I=/d]DI4+5Q1V5bC)8S\fN?AbN,?_J+8C6gAF:bG([+HBIdTeN=CWLV<IfSB
N\FUTDb/JR;J?,<K#&aG1G_><d9E7^Q-D8[+0^97\^VGe&IOCB0&#^XLAAF;;DG3
>I^6>,GRdf.HWYOeXO<9YT:Q?+W50[+3:.\b@C[3-L4Xc^N\&QSQOe1]7-S,BdJ,
:A6e/;2cY>[(#-HUa;-&EAdU:T[W^TNM+:+V0MX=7B5,/JG_IEf??^1@R]S,X=H0
\SaCD+D/\QZX81N#Y]F0-\6RL;#_#S@5:S3fU;6#?;A9CKUd,Y^c;PHQ3,a#5=2e
U=;8SVD?J_\)Wf?RaYS#,STWHKe_S6NQ^J64XdGLOQ:V?6eI0KAM>4S;\XX_,^=^
.SHQMR1>00-e=M_Qb._BKCc3B[ZVN/<JffS6D/IR8B,Z:0c6M6+2EB<VFB,V)EPc
#T;;1G6IURH^^>B+->V.O\?LCVV2;1_#.#Y1CWD4FFg-LW<W)]&^dVc7C<Q1Fe1c
YV0[Z51E,@/Fb78OD6];WI,FdYL(bV#E+.?aZ7[a5L_KY_YIH#J/-1L@+b@1<<@V
(N<:<GV#22(XCR67O<G7P]:_)X<DCfMS>J1B7:57N[S_<IL99eZ-+1R/Pgc57Y+I
[=;A-.I4cE[(If@PXL36-V<Q\S^)RT3/>K^IHMB75_e7GL^(=bP77+#bG0Y6U(S)
]C.063OO9d#(MHOc;MU=Q^XQZe3R#-;)f:UG[A2a9Y]T<B&^.fWJfg#e_U5)6&5M
.00K7K&;MQeQ?(@DS=bHAB\VT-&?-06eB=3d]TI@+4[e/]CT=Y#6eg5FW)7/FOAI
3aX;>5X9/;WJ&eI7d>QQ>>I5G)WNL[dMd<Z:-H&B93^cI:1Zeg+LT?8(a,(5DKMe
K/^)A>ZeTJP&\5C=AK-[>/NZFWT6J)f.K;=[e1VSR,eU5X?Pd(KC9/C3_W@^.=(\
=CC=HH+dYXa9SB\A]^Y4g9Q#AP>+ECZD#5d?W10VF3dQ-HS/<CR6=bU)N<>/PGCJ
.?&QL3HBgb-T,IF@b[Z<LXMA7U@:5D4TR&J;-4>/Y0fE/TS3X6YM\UE_ZFd?#P\(
1IYL)=Afa2F/1aU92+_g=U]UL=8R2UPW@:+:<?;B:O=d7e//bG5,HHdQ4#&G_MZX
cAWe=BVLfUY/]YMe2Y3UcH(N?=76-@;JV10R9@b2R\5H[B4aKcH92&aBc+N=7aI?
c@gS9IFWP>-QUM[8IOR3bY@8YaT/8afcfHF[@STfKE#P[(AEOf,K=3K0R.EV-eXO
8Hg)L>g28GG:J6.?5.J2CF;7,LC_N)gXA_U?9YRNP+,M2?(-?GXf(bXG,>.7d9LH
#[Ha)+M&J=+GN#5(<3e(-Gd?LKgA^gB3a_U9f[F5F)21EfaKL;8Me-1b]).f5KOW
^Cb1feV2^FYBYO)/E+63Hd6&Y0<H(6cO(RL]WO8S4\\a2baO^+aK7<J.8;_A5gT?
b]+DAX+fUGH)Y;<56^-OfDU^XR:@X/H5/V?1X;b3^08-PYM2WK,RSeVScP?Me35?
O.TK,WKU01BPD(@9>aRb]:RLBZg,<4784,5<8Qe@0QPIOFM<<UJ+(;LDd<UOUgbL
)d4&4OSM7L(V9\WHK[cNfMC&6#MV-dXYf>?#ULJ(+c/e@E+[XO.27a=+<a&[,_&3
ZacJ<&@8K68QM1ggX-#aJ?N?a2#JdTCT^eDNHJ0aBY8V-9_N(6-P@JWE^]-CKNc&
&T;6F4@;g7b<1TH(G]O3E=:#V\H&C[#98[dBY.P48Z4-Gf\3:DaF43XR-DY.=+Jb
R0>S+T)2b+@94520NF07bNI,]/+\=C7+S;A/=#@@bH;PR>NO97P43ZGg^IRL7FY=
MF4;NM5?^M\G82@186LLB]^24Uc5J5>7I@(Wd2Xc9A\33DdGXU(]RQ4NDH.eDLgZ
SG7;8g.]\3S9(/M66&6#5aJL04NV-G&AW8YAR&F8LV.JYUB+<NdFHMaL:1>WY_Id
U._4856;6#X1Ue@7XA@,WMOQY/@5C1>a25950M_[>)-_GD\\&>G_;Oe9<+eL>->@
;OADOf3GeT#CL-=PTY+(^SScSH8<d\>[@6WJX;OO<B+FJ4Q?bHO6.^.3A]8_#W:a
MK3B:ZSb-H0KdHcJR:0b)M7f5?)A=Vd_-_f@GELb(#P(+RS:;V7?565=&M5VfX99
U_XN,>IDX^.;:]H8e3,YF@Y(92#^<X_YDZ:Pg0R[fQN(#BW?VS\AZ^72;UL<=O-P
EX4FYK^D/7V2;;)Eec+\/gaGM(^<R]A?DeSM.@D7P<]-I05COdeA]DfRB#]NE=9H
d1\E[dJOS22AYa>902KMA\K[@#[dOO&S_52]KCF_P:T^#2C9A>CUOTBPEd4/+N7-
7DBMf03K:/&OMJ\_Y\CV=9@eB)KP>5I:GC:/eJO.Q@GN@6FNOQHFJ_D28gMVT@d3
/RgF]5b&T4(._ffIXH2M#(U,,[db9g,E/C.V:EH3B598)4KWI0#(/,7>LE1PBCHG
A>:/4QEPFT[B5-_Pb=D=2fG[+\)Z\79[d&78^#gWPD;N^9Q>L(6^X(.^O_>MD9)W
SO;I0<B2a#/OPePVB75&4Nd>-L[5:Z\,FL;=XFCWW92fN&J2NRMQ4D[IN+1Sb01I
XcXAX-/K;B1IfAQ4,YeY2W8H70MEMCF5#ML7PHR(J]DU:a.2#<G,?Df43b(7.AVZ
HF8eJZ]a#L>E3ATWZ35723X)<Gg[9N:B<1FC^FTDC@=9bS8cKW+YI1Qb/Z=J+:,/
?&;E#N0C8JVD#S8KA4B91A/ae+EN;E2UMgK?B]28ZAR^_79a51BF9(D\#CFDPe<I
gJ@0>eB=Z[SdQ5(-PgcMGAYO=DV\29]1cC(e1#f#IZ0#?gK(3_U\aWAQ)-O?;JS6
L):T6#O^P^fBb;DHH&E<L.dW7HU@\\UD^a[WND(@0-)L:Na8BY@Nd>T.AZ^YHV>7
A0W=F;M7@YC6gEBJ1d3A(ZTeR@&N#P8.<LWTG_;255aACV8,-;CZ,3WUS3dTcY4)
;(Ff_Xa7A27T-B-UaYHOK#-KJ_NbdZALbbDBB0M<ECJgAageR:?BE5M[[;FN+_\]
E?M,e2^9]>Pa,[DcI#S^Y)[23.JHZU<]UdWU5>cOH(c,R7(OG]F47eQW7-5+@;7Y
+BP8DL+^<^/BYaH;/C-2)OK:4;EI=N)_:2.G.Hf2QO7^#U=AJ\UCN+adBBJ?>Mg,
c[V7?+3QLaO#PI6GD>Hg8EH>B-:BgRO6AbKOHg,](d2>,Q[IXGPDe^K1X)<K[FG(
g;g#VO@?Bd^QgKc>b3[6P5a?#277^=#CL_VY8_B](.TeA9N7a-7.]0C?R0#9\&>#
+e,Q,>f?,7P9AJ:6,<8XdZ7;Na\FBV]=NT(VN#5WV[/D5&^bL)XgS&SY\)>2?V\T
XHI,)31=3aY)KbKaNQ[(7D,T8\C_aPYa8c\8JI)<FdZOag5U.9.RT[10QL/\S1:]
>3TI_[g_)1+Ifa;A#CDcU>NZS/9U?]]K9Z.PWfSdKdLW<JYO,E0]BgCd(>WC-2\P
TDRb<R,>0ZY@RCKb5#:c&0BUM1>YVDN07E#/=K8_NI]:G7L1R?4V<,6[JdL<TT.T
e6c3\79La]W5OT7DQ-XILBIT1d(\-++1IE&_@5R;P:e99B#&Ie[6,4<ND/HfX5bD
S;3ZJ:HgZ3U.,dVKA)L1<9HfWS)DYOJ;)O9EKB(6)1=63(,Uf=D3J,4(@04[X3XC
_Q72L/@FNe)#\5@0TPJgAA\:/2HLFcC]fSH&4gDCL7E+35-=:UHD\U:ELM=\7B=3
Sf_VI/=^dHDE.Z/[3\]0+bf>9<eN7ZO)/0,@I-+=(N#516-[9]?AfVT=6@.EY0)g
&.PES<LXX3KONO,G3c-CeSaF\N]Q>G=_OA/^a&W.(,T)AC-D9Q>F3]PSWPHCO?7H
c,;;TX^c2AfYK05gfY4S\?O?-.&04?R5X#F<7LD)B_1_(1@-gcfc,4KMUWV6.Eg:
(H6R.M3DRNQ(TDGO(g-7A/NO1M<EfEW&G2V)0H@,VRK>K[1;[0+Z@--WMaJ\BV,2
X>e253A72T;,EH(:<J)[A1S9)L\A9a]@bGBGb+[)dC],:0dcRgdM0=;RaCX.Q/K.
[-<1TUZNYA[fgLF44DZ4J(QI5J55G3d:B5+fH5]YR:B.(9WD._/aK\d]Q59HXBSI
f<E.dK,1@BD#?AKG=d?Z+_[)NV,5N^CGQZ08J[/M][d]1#aB(.E-:L&6KB/YOCK=
a6+b@O]f5YZ-3,_;63)#ca0M3:9cBE<&MD0#5D<e^E+-NA@@NKSTL>fY6W?C35(@
0/8SbZ8_3)fdP]BM2Y0I9<Yba).Z/CI?FDA&[]\-56PJ(K:4,69;:U+4V?\9?HSN
VHEU<dQSg6+Hb10Z=5NS=1];U97Z]c,3D&1Ug<f#Mb)5]d6A)bVPbQK7318)EEOJ
NJ;Tb\Vg@[#H-#a8#+)P#Z1&JL?L9KM4K-BDASS(EQ+?/.-3Sd-42^\4>2^HV?ZB
AT]S\Dc;R2NCTFS5J2VI7,<3g)NEZ3RA>LFT+=I717/(:M5YdfWXGOe7R&SA=K31
?-^/4VF&OCVSMV[e8GE^:He=U_P<<[:aHIYOI:4gZTCF5bGPg+Y8GgJbDKU4K&D[
Xf6X[\#WJCE7<L;ESJ@]_?^<eY;R;2^fDgF(:?28@]=@FRAf.3QIVa\IPgXETN6X
3VNW#O;7<fb,\W&HKfJb@fOXOGa6gQH(P=g7[AMd;Y#IS[B8\dOV4QEE;6(gH[2H
a&,^_4f9DO4V_6F0g[+V))N[;3M-W4\4EFcK9I>?d98=cd<TF@2BL3SBDG193#[J
_gE72Ffa(Ee-?;@9Ed,B4M0_0f4)I]:\14/#PHcX?/VKbDaPX6,8S-V@.MMDLQ;a
BKgIP?2-3<3EVUJ?7aK/\LVBEPK:=&-/P7Ua#f18#=B1&;8&/AAQ03=V4Q]N]4+E
RG#MJ2N>[98^Q(bAQ\3+_,F3dAM/Ed]cSCJQ=1,cME)=c9O9N[<ORbf4B7,cK_cI
36e49Z/JP17d8\I7WZ=Ng1O0AV)9/EH98\JG]BOO&-62@PfFg9W[41KN7gWSVPWD
/YHdEUO)g<(^cL2;)9;]cWXVDN6BO-e]5CfVP5dRbH3_:;,O1Td67DR0UO9VT543
gN#9XQ>T&@D)4R^EZ3TS-@\3[O0YL,^DBEgQ8ZYWW_3E8@.D0gNK&g0>f&;.BQON
]a2+N_OZR<:3[1&D1PT7IR+8[Q(@<D,YK\c.0.f48dgZPZK#=MFSaX/;NT<EQ#?J
5J[TGN6:Jb9[VM^;E1L/dS015-ZO?RJQ:14&gKGQXd@?GP;UN01fA4&JS&Ka0b7V
I#&P+bP5H(0Q6+(O;?MLV(8a.d,09[E&Q4Ed<RDTO1Q(JLTaR@@bUZC@OgdE/O>M
Og/;WKEH;<^g&RES+GbW\Y8]UIG=B:T>.6QO:B_K)9@@M.SC@EW;8_R8CfdX4//,
)f#>EaQ/aY2bJQRU2SSBXg:N-[R3/7-5HGMQ<YN32W//dQH#M9]XAH+ZC0Z3gRC2
XQ0^?:<E[A]b@<PD-_94J?4WO40]M@T+b2(7X@ZUWRaBR?V#TS-+3#>eDXIQ#+N(
S&4?.bKI)O89)>be+[]GJ>f?:I31L=9.&G8+.WAXP_g[Ke=O;Y\Q=6TSPW@b;G6(
:O.G>B7R\DD90==^E\(:OM,3e;EKJ\36\YX7JK:HZ\=W0+Ae>aU3//6ee5f:bNWG
ERI3[)L(-)d&7#efT]H,fV?g\,7)0\,(Ra2c^/KcYDE&EVdXX54&Q+5O-B=^a0J^
+f3T\&7GOLS8+ZYX+(=5Y>HV[+5.UEBP9?U8-#c0+/E/.LgDC<=(b_[7K5,eO16.
ZFd8WU6&QR-.E=[>I-XTT@WDbB<,1M3#YHNC[M4D>eaS_&@)S^34WI^1:67VI7JH
2S=VJB>AaU]]Pg37><2U9UdP>8Z@a\6JZ-FNY;WN_5,YX5Q[@AT/aZ0=[;1SNe>B
_/9I7<NOM2+U9L4[KWPc)[/6Vd&T2PY+1U&Q><B5I3W>+VB_[U-I^L?HW:aIQgZE
&?IPeL7eOGG;FBHSEMcUS6]WSL6b\8&ZZQXEO[1<G=.=\1gB2IfG5_EJ9@YS6aH+
J1PeXXKJQ0RJX9(-PB,3\9<G)(EZdJX,B58D[c(Cf7Xg-58CIcb+FR+D=RCWXXRO
IVXb:GIf7=QVGfW#V(J=eZVcZTd\PIbD;.[E[#^<dRO9TJe,LPQ&:P_IS:]8NQ1^
&8==T5Jg4a?-+HR/JB1==PeF(.dBZ?0,7SP=S>(R(1TL2NgPdR/3Cg/V&<fN5H=2
WN;eQG#,TK;MN:;&I)H81bV/1d(+V0KNgc8f@Od^.KI/c>^-JGMLF97#&O_HKeaL
Yd##I&\,,O;<QBCQN4R\8=KJ<aO).)bG+BQCNG\R:;D^YT?KI^LaDUQ/>e6KQ/g)
_.BaC2SbL:W2?_g1]PDTF3,BGcIgP.5,;KWb/:g>3(_.YSL02XLZ)[(70\gWXf@A
X:R4c1-3NDUa=S=3c<Yfeg]@ON=MNW:JWS?d+aB@V=cZF)UNY6^=7YB?Z+BL<+@7
J[)FK-.TA+dA<c>/(C3^3873]22J>NcGL/XHDLMRY(<T6?3,O55U,[f9fgC-8B:/
SF^:/B(,PN.PF?JK_)60OIS+BfNf^_d9P++8^R-Mb2942731+C3bNb1.BB#;cB[R
D1^,0?.;e:W^2)Lg)QF950##>a<H&8>/-7:DLea@.12K<D;@+H-_9MNP2XFXAYe@
Q3Fa-B9UCXEMMOe>&2,^X58@8+V&Q4_JfN.a_>H]+/+2[5J<>H#VO3Bb1fC/DL9&
CNc>g>]DB6&BgR]aaAb:=VW3@,J]Jc?S(>MNAIa9+eT^,;+1P];C^T_>3Z4Y805I
]8E;H9fRJ,b9V50d[Vc4a?;M5HY>Z7c,REbXT)/ZD&+6SR[J?/CH[B[_?\c><SY4
8Z)d/AY:37DONZ-[Ob77e=0aY>8QfBC=KW3TFRQ7M:,/PSY_)SXAf74_0QBNI9(>
/5K+cTJ6c.@<H,PS=T.CZ(a3Jda\_^/R0b#3]Q:X1=bP#gfW+7M7,[M:TLA3N\IQ
-DSN;DINU#&)eD>Q2NdN7<?4<QCNH&bgZF5D3I.2>LLG6.XNE3KM[7e8QC;X/=f@
?U:b0C234\6cY.TH5__/c<6)ON7HXMFXBTQH(121.U\4d8FLX<0:8^08H8@494\N
NT@-2I8.<Ga8SCZLQOR/DTN_)J]S>YOS_Kd3F\H^3Hg#DP:GObVTO:@4#LXSAO,1
(XD_XdRIV9=_F5BVSL;#gWCTDJM2\cO]Z]9_<@&,70LV(8]R,&MYF5\]D4-eC79I
A?07OfLI&b\eaN[aX;bJ_B.-OK)-cX(8W/2[TSKWZH?f1J&[C;ca<EK9JG0d^X+;
[RRM/[.^WG+9.fP]#M-AYW843M&QGXeSM-+;E(X7JG3I_VF64\&K&V12WB:J]e.F
FR\C<NRRQ;(=X\gc9)R86:>L)=c]5P<B?,Z8X^fX4#D@-CgY</W.7?b&6(I89VI&
W75A.XR/b0=Gfd-7eU1e1R_f43G\ac9HKG)L].WFRd7Z@K#bR[&H.Y_Ea5aB4_([
;_W_83.=JdGc79fK7M_Q[<AIAOC&WWW<:2Z^_Bd=1.ZIQZHe_9BZ(1fKeCHV,90K
#<]CA]C/WKc&2B[>0BO^D,C\Y^&X59EDaVUd7#80PK[-?MGQ@_0F2)(5T4LO4Ya\
)aBD?J(deHXQLgT>CPHVWZUV<=5/9L=-0G)JCLCW[C>_K:O7JY[W+@7c_aG#J@Z>
GHD?XFPe;(_3:X-)7F(9@7BO)37&=12<-8UC:Q?J[-[aC+B]@)B=aOfNaD=T[f>c
-Y:EXEE:/3UPL,30K/eQFV@.F47,<1:--^Z^J<:W6c&]M3,?DcaJHKYX#,;+fMJ\
,TG-B95bEB_#S[4C4N/bC6e\gB8/4,4e)aHZRMRda/S[b.EBa\&e2Ng6PVKIb6E7
:aRQ@J3N;\VeZ55C@e:[T)d]&HVA0FUY,,beNW;&PY?Qf2PM3[@9QU>VW3YW=FPK
7#KcL_XU2HA/aM0/R8^4JLEbac.<TTbD4<@H[eb/CPTC&(37^5=W(9.\@6R(QTRR
1;8O]9Qf^g_@f,>JGQaS\U=1.&W6.;;CgT5:YQ+TQO.BN9Y<:T,[dAAf,Z+WO_eD
=^^>PD.Df,V0=H1]RXEOB4NJ03]H8L\(6RNf4fSND@f/4U+]#)cF4VdV=QXAD7CR
?:;2W_B?01&F9ZH[->?bX06;79XFS31;[QUSNHG@JLWY1PKaO0(1eQ(_T8?6X@Sg
a+YT]aDNddA+HI.FS6O81^2dZEZ3BISP_8@.IC4/0KFe&S=#W@K^;H?00\1?VMVb
1)?U-V,84<eX89]V_6PX:@AK1JUA+>EY=?G\FLS]4d;:fEY(c8F6UaS6&ZQ)D_CP
T1D6<V6X)+5b;U]KS_N6^QBe?..Bd=JK52:+UWbfcZZ)_H8e28]K6LAA5MSW@RWV
QI/<CB?=6^dMRY6Q#C0W[NgdbO<??V3Z7@(5;gNd1Pb)\c=FHAA2)FAfI)9HX&;9
4C^W]B-DV&H.)UW2UaePGDR)bV?,MIZf@=_QD1@72&2O71VWTR6?E)C/0\5LJ#R+
=Y95#I6M?M\W=]dLPcRA#8X[7e)]EVB,3X#+F^66+_?@3EV9@&DS1(BBad>2A<g&
(0?G20\9CD0+?cPS2P=^+6.gC2F#eO_e6P2Z#=FKRW^?\G04LC+9(6PgC)8H;X[O
b:;B7:c.A[LG6#.^3R2-4/XDH?L_DDTD=)4\GX1e-YL9KVHB6Q\&H]+B3(/e5UZ7
L8UK(dbG1ROEMQ[T-]K/bcSaSW<0B@ZU#?PICL@W95E23<fT[(VdX5@\Y_8;EE@F
f]@/[X:8EEVZ3O>/CVe=[dAb5/c<(DFG[?5TT8CFF=_:G>:?.@Q2EbK/BL\/bP0F
>H0ZAC0=VfP1SC<C4TNU.\ZId[V5D+WdDRb[/#7,RF3=S:d@91<TC5Z>TM?>?]^>
+8,T4,7;1-WUH88R+4>,Z].)8=<+d>ROYQTaTT3MEe+DP]Yb=3M?:#1(]GB6bRK(
O.7MW#GB^1L17,a3\f]eW:gFYYV+_BPXX#E[2D(&HaGM_M#>OQ[Z/,<OQZ<LD6MT
dN22E>(FfK27d]ZXW?+J>8SU8V(d,-KNP?,&2cQ<fKHIO[CDJcEGQEHKM.)W_P_[
L5?67AM&.7RM)K9_Sf4Ua^Q<(OgbD58-R,c4P7B.UWVVMUV:U0AT[aL-03#c;SR2
AYDNKSUW31J,_;\?>&_ZecR(@g(3][3J(T.FE7A\c)FF:WdC;Ka=Pe=0&2gV+/A6
3],44-W=E-YD@#B_6CQ=TNRVUD:c(I4[G)ee;_^./gbB#F84Gb&#eAV7Gf^BR?Fb
@dL2TeK+OTdI74XXG0EN-_b2I>XL4;Cb_U(-[R7)0G,9g14?ZHe9[M.JIaDT/\VN
+XeRR-9]580&(]7>aF0:3<:GES.^71RgI-QKO=fD21V5]PO1(X65Z2efW3aN6\NB
36_(JH4H]#)^(4:FFKM^X:_03E\d&dUBGf;8NP&FgAJC)W;+?[1)_#E?\^RH6.6=
e4_9(c4@[e58HN5A[=T0FM9WY>,&aA]Y00Yg[JbF34:2_I/W]8bAW8VX7Z_agSD(
CD1Of+GW[Jb4JT/Y__?=)8Uce3SWQE:Q>C&(61;fTOC+d^5N/+(RIZG8(^TdU]XL
f1^YT.)KJW#ReH<cdK4fZGbg\:-^;YEL_,MOg>GBVL^=VV@g3YHCaK_/O,_M([C[
QZeGfH?OO@g8E0Ag/3Z/.(VMOMI<O[JA1MR.J11GA0XB4@VZE49.XHYLOQ0MEUSQ
O5V(,238W)TXOB(7R,+bIHTR^:QJUB5<4#VX(LN5?N,#)bCJY9R-T#J/QPe;HQE@
DT2.b@E8SXegRUA,<X5CE3/]9N#E;&9UZHDf(V5:J_J7J4QCUHUL65@J.-#2a@52
N2VaRR/5Q<>G8ZKf9_RPV^XQ\]D80^>gGQf,.HgYH1UG/=a[R8_B0bWfYI;C;3(Z
G.3L3X^\L_3:-Tc1bPTSO55c)g1K.T3I9Fb#7Y7JI/&6TgPAU7TGK/PL=>;<N=5S
+0M+AdPSA#&9fbEP>#-GVK@#Z;4<eQA(::ZQ37J3bd8TUW-9f+_4c:9GNVgOVf>P
2UG=O6a0eEI\W@NaK<>LZUf&^+(e)O.1\;40;89C+:9B,4J;0UO5\<X(9]B5B73.
6FL>;GH/g^f&7(O56VYMIE3;WdZ/LT-_@Y:a[FF0P(8OWGJbK@290#/Vf3ZG&KJL
1?gD6<be@HEM7eL2#R\Z_P3fBfUN?&&\T:BG=V3J/2P1XVQ#3ME+6(MFA\W4.UCg
:T^c4KLR#fN?#IHXD<],JUSEX\<BB@COVTM]C6]<6;DaAcWS4f761_7I,8.Se#8@
?[\_Wb)J-^WY3VG>62083)M[/d-)YbW:PGG0fL\^&R-52LWPf62@-AT[DGAG2IC9
/I6I/1a@U\):dNEVC1HE=.8NJWCDF=E5)::aO+R[QX0USRE;+]=<Gd9Kb7[=D0RU
LeN=bb&6@5?<I3_1Q(O_&cKGe(#Z(Jb>1+@0?#H=9+eY#^W7B8g@TIXF:<X2TfDM
-M9VZ[E:#U^dB<A7YJ:U)^0Df(?OMgc<,VXUYP>C7^4,\;\e?+C[g37X@Q+?T?\Q
92SW6N3J1R[NTK4V/H+P@DcFaN<b6?0?aaBc;Q^#Q6U?GYY43D]aNR+K]&-=.+:H
+e348-SF?79DKMSJfP-J/]S+7#-b;Q9<21,f_T.E=]E^YB&8L>d<<a;0gHZUU]V6
Y\eT7XTSE,JMEJOCbREFC]DD[01,H=1bMeaBF0PE<QZ;Qd;H,PXeL^bG)[aD8Ug3
7b[LQ0?g<aRf[WV)_J::(R1,gf_7CZGPb4RWV6G;f.X\L21.CO]F&KEBJM;>-@D:
,Qb_V#IUSe2/Hd=?.5V>Z6WWNS9A&>gP8RJ7-35@<N:4-LE)DG1[ME6KRG3[)1ZD
gEKH(6H9M8[/FeX@3>8eTdK&LcB<3/]H9?O\3.BI=_W5.VcPD.R,.TUg.0V(Sa)C
#7G@48FE0-Da[VKA3HPG>S43;6+99^@<5HKR^SK]J#8Ab6=MO(P^;AGG66HdG)/b
[WO-^;:::)Aa,OC5eUJ6[@:B@0W7K=BQAa#,A@E;8YdD((&fJ&=&R<JXb\SW9W>3
f@)J=EN]I:=dTZ:^R<Id,ZF,B3b\J.K#4b<d/4YA/#L?CE@?JSRBRb=GbR/Z7,bU
F0(FD+9\=+6A9E;->3T#\MZEH[E]\]5[EBc&JY6W=;VS(YVY,WHS>aG@]-GQ(TZW
(O9I^EBPE<=-RF=Ceb4MbM)=.=ETb].7f0bE,=X&bTM^:cUS++3HCWJN[gC[VUc7
=.^Q?H,e_B-<S)e;Bf<S4.MW#,8WHAO9]RXAOF?,_DOB?Sd]#D9N<5O,9K(ZT=f^
E[c<#bO@(OJQC@,)P&eS2</^:/FP\<73HN4-M?6<?Nge_cF-\ZA912C>);bK2\GG
EUdCbT,:R@NBL.5IL[]RSMYS7PbZK:fO.E_;0M2V&RCYc>eZJ@^W+-VD1^_+CD(I
R&R831MU9QJ,G)]/STD_\4_6.==d:92VNR>JLDGO#1HcGXbU4I>KFO+@MX_XB[YK
K/5XA=H6[FQ^^AXZ0aI]+adeTS.8Y5Z>NQ-+HEOL=Kf5dEV+A7YU\_Zd:^@E=K,=
?Q/__VE=S6a./F:1@R/Z=ZOBY8.1&f:bdd0OC(AVNLWQWQRN:JRD];>OD454:I/>
PNCY+P7Qce5EB\HIUE1R/_Q))30cC3EASRMQ\,:^f?P<N?,G3^+:W\gA/,FT.T(#
1O(1JFU+\XO2BG=cHE+0L_H(@JW+]4Q7eVZ3ET1#gEWZaK^2:HC#gYeKU-7dQS]I
>6,ON^VW.[RG9+)cLcVN@QH@/]TZ]DVe[9-@^[9Q8)N#97SVX<+a7M3E_9Pe97?2
\URDCGCWKEP/3>2QKI\SRS?40SFD7RQ?Oa9+X/#Zc=LUS=K>,7aR7?<#--M6K1ZC
T85657##S88+>#JIN581I#_ILbbXNJ\D)5QcG5WaEc(IP0<]3+W=@M@TYV0Pf0T7
Z43EHFLOFV^)8<g;1@&>aB5AI)/S=NV5A//4G;@2L>2?7&O^4MW3^5Y[fHLV&;R4
O,c,FGK4aD=;(=2+60M=[DTOW9Jc(,+/]JIfISYTD\SMX&JaH7,[eGF38b>90)]L
ZQ]L<4B^EgS]b]d[@8.XNQR>[MHY:WXW3_-VU:P1#2?ba7B;O5V8)Wd7(c()VIa[
=V3d6\9LRJb_<FV[9V)Hb?Zg);dUfU&2]2,EgZ>33BL7__R]EIY:7fGSY^A:O)>1
DPD_ASeb=<65>.J5d:B5@0(H0J1PI),M=E10bE_AFg0[WC66(F0;BGSBZ0ZJc+++
QPKIE.]JR9J/bQX[_+HdZU3&P(PUM]Mcfe-gD/];(?/=9aa0KYD:e.)S0E^+_>N7
@9VgFAL\?RFW+YDX&Yd<d-V?.J#)g<^df?]B#L^/O?Qf:JdC?dfb8gKXg9=>6,P?
B\T_6J)];HbDVCW][,(\CT96)JbV<F)PDZCPc:<+Z7/8,H6.UX\RA,.?>6;46g<P
HO;JKC^.X^9aOC^Cf8g4\W4eOY3aWbHb8FKBS\=:P9J^G<RX-4&7^(&>@/M,3HcV
:IAe9eX#XI28#_;\,S.TZE5-(aZ5Q]:<GH)1?S4bF>cRW52B\R[c(7[fG0fSGFeY
f->#:,Y5e^V]NOH@K/Q^UDdHHI6A7,#>VS[LW9@?(RN[TcUbEb:&2AK?ZWZI/513
d2SP6W<Ea\e#H\6,R;2^1a(e:I98[Ba#[Rb4fP(TaS7@+fT/F5(f:,2;gXU)PKO5
K+(YLHb&90Y4I&0:3,0XTA<-74Y=\2g2[Vc)C>-bRSe=>>WHFQX8B8(BB[O1T\eK
]gKd;[GG9?320KV3_<dUZ@;7UcdDX]#)X1L(4;QK?1eSN;:50fg/4GV-aaM)&2<,
7REG6<I+NCA0P+)>+T.g(IV@4Da,.,+:I;X>I+5-Q,2I&Rdg12]^fDV3We&^dJU=
2,b^,+ME#WZ&NBD\/U;^7E]):T#:#XEb<F[D5EeF&T(^TC>.4[LXBE)&S;6;2B^R
]g((DU,^V6&JH]GeMBHN2^,VBV\PO\5;B?DO47=G<S:KOKaWHJ(DEI<eF>BdR<+K
NJ&(YY:,H5V:E_Q>gXGZO6^2>QRGX<@Dg)ES6(#QBX+77Ra9I_gXX[F@L(e/&2^T
FI3^QG0I2H5da:Of2=85<g.@;HTY_F7:N;Af^KXf#L,C\)7b=f[9RL#3=WW+4#QN
AN\>eA5?4T6E4a=LL;Z]\>3/WggQBP7AH=YLY;gF+VY0IYUM&f2\=;U4^CCc.bK4
2AI/N0+,Z3gY6@<^dd,BCLgMA^6WYI-aK,I&#V.1L2eCOd20PGdO+1(@K)GP#+T;
Sg598>MfeV0/SMYgDE+;]<8ZVKf>g0c/-B8@1<aQVU>a&\8f42]->F>()B8XM.BP
IC2=;6IC[3L9N<c)=4XYO,L8Z.2:bO8HLf7C4,<I\[=_LBV2QSI6#DD.deCQ:ZF0
JbF11MQUTf4;WPYN>0f28T.^M0g>_D@<\8fNC.]MO=\B#bQPQYF-WI_#BO6^3bXg
1&Zf<ANc\Va,1,?8V6_T3S#@U8EN8F]F3QLKdPeHGVG7):PC@b-EO&Z--,NHU;].
56B(_L5#ZNH:[6^[P>EDI==,9<RC&cAOc\(&2S&B#^EgIdJ\WM=WaT@X?0J?Ja3_
+0A1H.J=#eZVXUB-Hb2W^W4F^Nd4LaW^T=LDbR0_,:)G5[[P8[YYU^;IaH-<2g@7
;MXQcbHJ92KV:6@,6(V,(a6&Qe)0-24K>-7R(^R93==.V=aMEXZaabJ[H0>gg,AO
eN\B<AZbQELd#[DV;f4b9aXe,V1C<-)Tge1J;P.ZW/6IbO?IA5FT\),VQP_fOO</
aB@]M66\HPSDJVU4.+.+<P4K<_gV,=K,TCf;_596_FHB63-S4H:H[NKJ;/2?EBg:
<TaE3c8PD38&)/Padg92W84F#RLa,P)bdeNPNd2<Z7#:/^.70YFG0>Y5e&.M,V-W
Z2M]?HK0@P])gOLe/HDREMQSZ&9Pb[,_.,_4#9FT[@[GIa[YD##@L1bZ7TW-;a_^
<E:8K[AB6B?AB25E)e3e(NC8S/gOAR&G\;@29C]MS;B685Uf-.d0g0(GR9]15Edg
[c2&M-^:2;5.32I_FPX?b8e)f:cce&K)&g7C([A<=XNL2IT]eAJS[?DNF^8bG+b]
M=>-3S-VRFYIc]&??9-d#,]Y#[&YEX&[g[+TE#-QN9Va@JWJJ\eU45/b=#X[OU^(
+G<LVVcF22\7ZCK?;S_&??#+MC(&N+B98E,\(OMOJU>&<5QIH];&O(\e5#ID\ccW
_I2(58>&P6]2U,ZD,R_TV86.dgHdW&=B3-c0@6PI=GOU_?)(1NF;26KN)-=LJ3]e
<1T&@;VF);=bCQZA9:DB2J\TL&E#DFg?3YV3J)I.NX]C-VYF+G;b.89<\BPcUSTP
.1fX;5.MH,c8;Vg9I<TX/C6)KcWEW\SfC:L=.5R1R_g)>R>WfgKcW3SXG:J)),25
[[ZI:>O(.fd^P[+[RDJCD_7)\f_)86W#/baZ3;fA?]Z:SLK1P>JF>T0F>/@-]HN&
IDMbd,SR>A&+EH5Q.+M.S;P1C22WQZ1:;HNH5563V]AJ1;0M@0K-]CbWL)\,eJ[H
)1/H@:Ab.[C.Y=K?&7gd;A8bSX7=a&0F0S753S<RDNcO#P8(RgB)[<Wa\-<4U6?V
0HDQMN5&EG^<SZR/XVIRf^b:D9IFSIK?1f7:#<.VKS/3c^&eYfIOA)/F=eOYQ7?5
YW5TbFH2YP9AIEDU/&6.cY8:]g^\P;&2/3A\3P1a:Xe.e,CEC_<=,4+b&D>@F@Sa
d+2dZO7Zb@fSWdWXO>CQ,)1GC:F,A@80:eGDcJU<J,/H?c7&a[A<(40E]6Q(22TR
CWW_-:(3aJe#Q7<^WZ(M93^@\),>+TOOENR(SZ/<^4[/06TFIgYM0C9R4<VD1[;g
#7])/_Z@Y?0d\XAL<_U-A0\5FeHff\Z3JB04OV(CN]QSDf--B?3a-C40&Z.\,3^c
gXC1)+P(a2e0&T,;TGILM=WVcZ:+/b,dOIW=EKd<GL<B^L__]:SU[^&HJIdYRY8F
X(:T?2HN+11VH@WJINeN=V5^9>=)e-ddEXFf2\1f9:fg;0<=W+X7:+P)B<,MH<7^
3BDZd4QI#R0_M+4R0GC5H>CT.dc@I,=C-5-^GPF+@ZgW80X/>]a8>O3U50dZA;1U
4f:AYe2QbJF&OQ\WVVYcA#QMX+b/SbA/D#QCM[WU6DACH&P+?LB<Z)IgYaW<>b6K
N).cALX6;b0cV3>SbL:,-64aSfY1X=Rf:.Jg?###<a6.8^U_4SEH7MC\?=+ZC9W(
BCT_XFcK973[AR60VYPfSH=+:UK@DNV=3(ILRacQNX<-<2YBGI@\+TdgNS2Q_UgK
>]NF,00NL&PH0+Bga#PH&^(1fZI[X+?YJTe/RFAN;.:WN?\,X;OR65-QXFDIU-Kb
_[)H0D3C;7\F.9OB>6cEdLQWb&I:E>L-YfQ8AS<6/&NaS8UGIC>RHc#Z(5QYEbB\
bZ0f+Ua@G<JKe9;@@e8-U077[U4\QNCOEWI0@/JKASaY)/P-W[;0CLaR1VV,U^Jb
?T,SL,/:OC9#D2&F??FS/MAbG2S>[aMO1:._HgfP#T(C61\F3aZO1,7fZcQ1.[>Z
<3XVfM.LI95XF:?M93<:FcDC<=+,BDS1BWgB#?SV?cJWGc,&;052856N;DTLOQU3
74J4&ETD_>J6QLc\,ZN:1D4bPg_+1OgN6FWX(>49,\C>LKaW]N^)BR/.<U6\WaTe
)bd#0CTT.K0ZDS9\&HAH;:f7R45JD8:eeFg4;1aVE1Y=(:]4_TI;_Q+U0@3U;ORM
V+B=<J2[=g\a.RV0L/<a>d]@0N6&)e5Qe[X3b;DW7@.g:JHN\VgKKE];W&WRd.BS
K1H)7X[Z]KP,;Y8IFf@M_EJ_H66_2a1f(WZ>/JKdCW5E^EgZJDEV<HHbY33^9Gg+
\-Mf+b[]B^31c;I7I?6FX@@3F]f(=#02gNK:S,DBfM42JFa,.&H>;Tc/@B3N?_7[
=&R?6b6XcC/+J-M)-[O;G/FGf<EP@EE=^Lb?S(;F.\&=B04/CDCQ:VWf;<00,b@e
5:;EQ3=@L_:G8EeB4EZ=B4WS\+/OM5QIfP.-fSV_P2]^F[4ObBaS,7C>?O@Z<0Q2
_g_3IAVHR;TNfa893&c<:P6(45fHUEa#_^0#]+.&=_@QGB>1^TL?+LR>VbT5@4NY
K<EgN4)-WZ93\W4PV):d:(?+.c)BALLUO4_)YIdZ4;\EgJ33C:SLfB:RFABTL^8?
c.\M#+\U/I+2,8FM@SGMfS>^2<c/Z?==;E]A^/.9QL]]Z.>R?N?@[FG0@3/]OE(9
1;@D]53H&c3Y+@SO^WK&C.)CEJ?B7+J0Na[aJgg[<FRBe9,eUdWM6JLPB/HO[Ne7
;aP+cLA]90DH#f8CMSVW)T9S]F4HAQ0..\:aTO94e&DO9(UQW[-<ES@+Z8Z6YOF5
+\WE3ZA;DOcNE+MSK?K[QWEe=A3a2.E=/1d\)#=Ug9ZG+d;-6c-5aA=^;8&7^)bI
b(Y.ZY-?F,>#5Q5MaXF;FS-]?f).Q?LAMCEYCb[:E;3;If11gab2YfL?,e&QTgA)
M1g&(]2+_#@VZXQbSX=192+,_UadS5>>NA4Q8PHNF<TJ,8aCQUc5Cd.e)_)<_3cL
T,07[?QY+fBP:Ic:^TL:5.g4Z9;5V.B,F>+K&>=A[bQ<)=P/g_R?HJfJ1[TKU&5B
;UdaRB>4GI_FFGeX-5-187:M4VI+EVYI^7@fC0IOg)Z?f\7]UMaS8Ef:-&;a(-=E
X5d(7HGdCb3A0M#Z3e/-MHM587+DgIV=58N+HGd:ATQ2T.g7U,+\Cf>P;=A>=O@4
a=3L>UDS1\,5#5>BYSKIg8FU;W_)c^N9F]<+/Lf2?S+GbX_5+/1MeC^^dAY,NDMV
X(I4\72-B2D048OE(?1G)[?RIM1GE1T8=g.<Y4V36&dEGG=\>JAR9T77K2f+/;C]
91Te#5/5Da]??eUb:4;=L=\=;R7/Z-Nf2MHHN<L,>T,1#>]::fQ/@P?14M]TN]M,
QGC:FHbFJCY\((<QI6EY-&g>>@W8..]5.#I3dg8EgXM:?Ye>KeAYR;Q46GU:BH@H
FICI]KVaTG=6B?U.XK:G5UAQ6\<D<La46MT_7CfRLS,5]W&^S,Oa\@#>OL/RKWDU
H<LEMBOb#,3;]+)NE@1JUdLU)U/FZTe)3,T(A?2fR5,);TP4Y:Q)XNLEZ8CAd546
\IKZK?;R[+TPR/(5EQ-Hac_/Eb0J^9R@P@AY57Zd:-D.B.<:GOLN#U[S#P=JV@0V
TB>RcgQNL9>eVDW.^M&76N-7I_&.&ES>OJGQ.2U>#@>6/WeP)3_6F]OZc7JDPXLf
8FGTMF09]\;=?#?PKTM)-91M+IU_bEc?QK<e[KP\@(;YCC@XXC-1]_#[0(EZK7>M
.ANPHIP1f@5IVX)7S_E9)^^QC5RUQE&G1f@JA)-f5552)X82W^;IJRH@<f1[d+dc
S]gg_-6&7d2+,=UW^g.#4[e99+CY(^GTOgE\+d=;7RgFMO\@^>f/Fc(@<1-KREeM
g4YXYfJY9ZEVW;]RY9.;A;b8C^H+0YME,;+D(EKP.(c&WBSG(5<;TGCNf)@(eU58
QKGOA#Z/V831062T1XC5(&1YT<H_\1/ed-Xb2b#?H#1ZOfDT.Bee4K5?<)OgaFCI
1c?C776P)</4Z1:60&TBBPP_GR/fGPHd3G1Q>Z:NLTQ(&#Q]baH;ZK^=PeN<8KT0
:AafRFYFZ@[1A[RG&7C]A:#/#I2V)\_2;/08#BU;)PTXTSV2]1SUd8GSR_U8_KbX
PT,8])XCDJc(G_6f9,P7CcI+C5+AN3HC[6F:^;D#Le;+Z#3.?=L)--XU08-@X)f,
g#U2E-LVVIO83ID5C]7VV<&a/QCWg+;TL@6dHR1WIB6g;C[.#\-1(1U0V(7CLb>/
2)G9JaF>QI>=QW(E&:Y/0a\0UCa:E>Q6>ZX&_.?YZ4gS+[,Z(]UGfe_DD49DaHYf
V29DK#d94/d;M^ENM=Wee:MI>H5e9&^R^^5WgYI_JR:NGDC.F9C<JbS>9U9=/TcC
1fZE+cMM9MIbB).MYON2I9V#3ML,.g=c&-_\B#75/P@QX<KJ<GIf:\Oa[\4958)D
Kd0>F+AW_M9I#H+VcH^U0KfbR]c.6856CCf3c:B\gf-(EVI9f<+<K>NS7YJ=&J::
VX(^L&^J#38gK1B9YR5:)T]M@2S9>g]5D4AR)CR-][#^[(e/b[aIKQ_X2W6)W2H(
^5b77H,MJC+=JX4H&YdQYCR]e-/BI1WMHgf0LEU&\e^gJ6=eM=7&H;7aINK/JZ+;
,#J.T91VFJ+./33S#H.6X8\(Q=N9C]35N,\[H:JQQJ&^[IaOT543-GPQDd.BZ,SG
?[BE;d)3H;B.[BE[fa/aF8e1A2BLW^,eKPQB;4H>^VQSQ5;/5FVZLGTbM/aT?/I)
(5/G[MEU?HI/.\ZaJ]Ec,N>1H/DGV>EE+1Qb(V4Z#DN9V<]];>U6(E_ZOB>B.A@]
@[UGH+d?(DdFSFH,C>51>_]g:]?+6&;<+R+UHT\GcL,]d#Qa6BZ+,_Z3C?267@;S
<-:22-3.XF>@4O_-0g::<V(;(6T0\#UGd5,,ac?QD.cLaV2=IEQS0??WOe7g^cVM
=bYb(LY(P5F>X/?YYCJA>U#F_/a7@Nbb]Kb-ggDQg>[T@-UO&.3MXM\_CIYB0W49
S\a;4<bG]+ILHVLA/?.)AR?g_3G-F>TH,@5f&^e?&77K;@8934:P_WD@XC3)DG1(
U7@c_T<GHbX1?ZE_EG<BK>Vff:J<1PZDf</:9T_3,a))[<1FL=CT.]K3=@&(,#A3
8DNB3</<96A;ME(&&+M\06IbY^@0aW(3:9R?NcBUZUKX/QaR9N1-I6W0.GVV-W0>
.3MV&_aJgf4MbC6eHP3)_CI?\W>eTV4]M;6[(AMZ;Z<;E\a#23[?[QdB\;B]G+J#
3Rd8[b#@I:WYXJ@RfYD@4gN8E;Z(G+(;2ed,DBQd<22[d2]3-CWC]:C]gWDg0EUS
;6YfSg+F>]VJ[^E8R&]TQdTgL=VM<##Fd:2+0:I.2]TXe36JcZ?YQ0BD:.82NMdU
HD(=\B6CW9#Y<baP2@_+<,@X^?_;dD))8MVIQKMLNIfU?VS\b(JEf_d>7D&2Yc\]
D8)YBd\D1d,6SWH=:)9XQ?U4;9Ga:efVdMJgcDdRc>KWb-0YY<H08daZaF8afXE>
6Y6[cgba^MX6[4DX4@W[5=8fNf+[^WK)1E5UbGB2W4S:;Z@OZ\Jb,f.1A?#62e:F
EQFC[->5bMF]1KZW6D8<S5SfCgH\PD(HSY3LReQDO@4Nf^DMG6F)5.FCHY\85)./
e,-/(:ZKcff)KN&D)?5G.<Q)818/#PgE0S](IM9MF6+(U1CREMFXX)cH?4Q&/EO;
0fT6I],N@7SC1<(aBS=CRV-INS7Oc_:bRQ7A\JOKG>364TbN\:TUE3DCKFc=([]H
41EeaG#\bb/0/DZN)fedUS#KCY#UL2]=X-64GI?16PJZg:-R.dNNTLS:DMK_-K<<
RN]-6eR^g:T?DE9dV_@5Ceg7EU)4BEJAf&H]>]Q;IUBB/3ddBNf323eAID8_:=aX
d9N&JXC[Be9Y#4WAe^IgH.WIO,XKfN<2PX508UYV5Sbd^fR@;,58+TV5P@D)4L6=
e?)D59,g(JRfO-QP-#3ZbR-?CM-6dCJ]6//a6)&Hcad5gCf[TPMIKXXDMQ#8dWcF
M(16J-NW]P<Z(9((6Z\,:\DQH[A@Z(5C@I,&DB\0&H\_#[A)dZcJN8L(4#C[<YcA
PDLZ;Fc=cRU)&WK,-?96).[0bXN[D.KB&0OCO9O@eG1\?&X>C-^<g^IALP1PL6DU
Aa;J7G_N=XK@WG6LQR/,85OX&:c#.KE1JIYbSY@R+IP;YBZ)SSQ+Q.>FK.:V1S>W
6WC5M0a#I3gP7AU,1[Wb8#Q=,]S\^.gW8VW2._BP_R?E(71LdE52-QS?cbA9<E8f
PTGUF?LAfX7LK>,7UBW6QYW27e9IAN.@5-eTa#>PaDZRQ_12.R)B=(.\S(5T5Z<2
QPeB[da;.KgIO2+B2BD5-/Pf\]6V/Bg2aL82W4I.SH#4(5#/<V:NA]K)fe-JS+A\
/a<g-K\5WG#[f.aX^\6/<=-+:f8A?Q;3X>>,>]O^IOZFU_WW9Y)E-g<cA)=Z:E;,
F,<[_2<BD45C;YGeN5FQ.X&3gV4X2ceXeUHTS<G5O<<#;fdVaT/,JBJ=Cg-LN?<^
^T)aKW;/_O9J5F_<.XL13EDXV\S9K\+V(</GD;01#T^c#@RfO/WE7&;9a&T&4Bb:
7\IR[2Tg-WQ+aQ8WF=.Reb>H(713@cL,N2;36a[7F?&5f<=[TEM4c=b@B/5egMfd
N5:_O#,]CP/E(<&I/3MU88f+3R,I)M1^R(2VOgM4S1W8#N&GZ,e4(,D71D[W/66=
L+,\)49fH.>g\7;=KQQ[Q#d-eG&Z1IU.H@Fb5EScIfRM=X/AI]X]Ycd<7XE0B,9I
Gd)<=/]d[,dORa;?UHK3B6Zf>=^PG?gf-0aWVHa,2>?--42)SHA]\G/CCU2MUQ8+
CCW(#98N+gA^LU4+UW=_.-)I(\Uc_+1NLMNEWE71-7BO#;9WcDK<H7GUQY.&K&^:
d3JabCD1@FCP)Q4Q[8c_F-2^8/aNPZB[c+L+Q&N-e_TfAf._-<X-TY#2QT<U7?QN
Q9R;ZDeK@Q[R+J>>7gK#O9Q\g&Y1V3R#[.[D9O^]<DJ::Z.<QFMH<d^WdEA[a;T5
-@NV]@I;2.NUCaT+04OVZC#Y(\fTH9VC&P/1OHc+P=D[d[@#A>4]E](_QG?TdJEN
A@<B:+4Z+H4J:5R],Y7-U@RSL;]e9@J/R,GYYP;&f1#b+fZ\NAOA@XBSb6EE@E.^
O<3Q3L1\Y/e^=(g/ZdJ>F2O);Y<N4g9NJ11^39YZI0DRLUJ_R0.dI?e.<14c9#Tb
cI6?T(R[?cd+M]VFXDYB[eR>f/QUdYP>&cN5?Q:g.\1EU,@UX&bE16_+H=_3KSb6
dWHefT/;(3a:KPYJTKc@(5,G.GE+YG>0-TFXA-AHQ4#c0fR=X,-]0JC7Z2)DD]3b
VcI2HgHf5LM[5)#P;LeFc0XT56dC@1cd=V.YDD@e28JN?RQI-=P<C8cDYg5Z:gD9
.[&5ffFb:cQVM4VWB(&e-?-6KMdAJH@/T(+PG_aV6aH^<f@aI3]^O-TRK-1UfA>\
0LGN2=\ba2af7=HaKXW6U=_Y4)9H497:J1+]YJVNgL85/K2E);Z&P(9dRL7_>(N<
4cNfV,]F+g.D1@=_(MF2VN>IE#VcCEVGA,E=B6#D^K4.#ZY[a+WYH2EJQ4R>2DId
#VP8Y[U#:KH_I6&d1;ZKGZ&Y5;O6HVP-+RTW/?Y>D5?RN@<?c.T87K-JCUMO3f_R
+K?48Q@a>CBQ.FU.Q;/;9WA^5[eIf_D9K:b7R[XM17<,D]XZ2;^E>aF3[+MLcH69
\ZY_M3A4aTNbFFQf-.g??I3^=>IPU^4I03V_#g8F.CG\/)A@P8^P9Y,[FQGUFSG_
XT1ZeI)=\XCK^8DK(6A0#(LE(^G6,=HUSF,F+dO[ZI+)8)CE(b1@U\,A:@&;:1M3
d<MO+S9/FM3KW#0VAaDRd</ScBF=L,f8,GKNZ5G(./;fHBHC],>GT#e7dad>7<W@
bESK_=Oc/QQ-FK:>,IMX]>-aTe6@\@-cL-^I-g;=.J3@V?eg^<A5X=fS884P\O^-
]M.V8-GMUG&6OUHG__;#&4&HO9Oe1Y;-G(W5[Z5\JFg4IL/EfCN0N>;#Z>@c<849
(WQOC?F-([-OaPX988I=>XdEbCFSC&A0G^16fP8A4PMW2>4;GK-CNXR4WVB[eDb=
V]e>PMQ\,EaO4<J@@:U=O?5\_9^WW,H\XW\06I:\LL/ERMZ(C>+eD,2W+bG>D,1b
=<HH]-<a+:1+/]d7T;\^)AAYaQUD,Qe&A^P_-\JX>C-g#\G#X7eB&dB2^N17)FgL
^dI(MM\>0MF+K#N@.ceDJ4I47&ZQ//OU;7@<Ra_UOPAV<X2+9Q;BR,gNS-G4QJA+
E+5@c4C#eWT+O&[&D629J;ZA+Z>R8O>a8?eQ7:A]?A=79=V#=TSc]A,.1^M:)04Z
QZ<_HXB&AJS[eW@;/1?A^WH?CWR2VNAC8g&OUKHY:eWLYEI25C4(GE5YM#W=0?T1
[O.DX0DXQIV@6Y[I?]fHCNCW=>,C??0H&C.GPLK+BLXc?3D;_>9f#:@C99/dgAE^
Rd<Jb,2a[AcJ>]F0bYX(@<_#BCO6TCS)>+W-5AMH:#0@_=AI;,P9JNeGPE^-ULRK
I^Z<bL[7CL+TZ&f^Z?]1N(-=f34QM&UX0ZVN[a05Z#:dM4,/TP-;ebK0>N]<E25P
U.18d83O?g20(f@&/Vf)KP63+MKRRG+gOMUdg97X:I;#gK0R+&NUGaB-a(g@5@Y6
Kg6[Y[QDa[7^BP+X9(HPBOFC25]@4+7ESAVQ6LW/[Fg5g/FRXa?>60Ga605I5H3#
;COPBNLZ6#_7L#(5VBM,6@4=G-eA(94G)BAYKO1LDHXL5E&df3-FFd)>/Z/K=?K1
54\9>SVJ_-A)4&ZOgF]>M7g#)XYE[K&bM?A1K[W<<O8deUTFHJ6UM<SAc(@XQIJ[
?)#PE(5Y8F>>PVFgX[JDOI6A47Z^7[JHGU#27H7dMd;E]?@OY/LaA?JC5Q714,VA
\BU+^@6f7E-[^E<,&F7&=feEgWaU13=e2=a=N(]-&8^::3B/&@IZG<eUg&K4;UT<
XE5QOb5<BVf_>41(+#^Uc[-A]^1b\bbBR?JeJc5ADCA]CE\^WW?aBQAb_^(TWVb+
?D-O8)6/+P[.&7AV0^)]WVTK\LeY5)E=cbAY3=a\CUE1F_L;<+ONe<<UU3;D8^RV
W4Z:#&T5H_SS9]Ta[]a3].2#R#VFCYc9K;dQ)U):U0I:^M8e?V@>Me7/I(PLV4I@
\H?&b@A#1\-IBAE5eIV/fO);]3<;f(ZDD9G;VAEb=CJ7Zc>^2-_-(_LFdM1fATVL
?&WD:FcT<BdX:.T?gK[_RJ]L^A>DK&Z+QE>dQ9K?fO;dU0-MUg@/P#U/+<@b^\0c
XUHCJ_b^80NGFWD_/S[KR2OfCaB,X8NcI;ZH?7K,V/a^G:-MaY:WJ=R8MV,d.B3R
]B+?<3.[TH7SDeX].S-]R>VfG9C6E849D4.3XKegW+-OO+UUc<49TO>(<==S9ED:
f5S0BY2E^D9@V=Q&Y0>,L/WD?8b=@>AQNBGMcUC3.WUJKXYR50Y(ZAT-GU]7I/8>
XWUF=c5>1PX467@Q1N)2YE&\/;5B;Ib<_V,\:-3UMQe-FLY^G1[2ET[Jf+4;/IdB
C09UX(G#S8T.C^>efCJD+ZN4X1#O\b,T)?;MSdfFIf@).3I@d7@VS51NR[_.?=b=
b6FEV_B619a9cf>M)>6bEdRASJN3<F3<3<16E9f6_3c6?^-PJ=a/13dRVe3>XA/R
/_[.C8FC+I>aX(W[dD4b]?-5Y;-?g&VD2TI@Pe&(5TGaSg.YZ[G[e9PVYcgOe>7:
)b)E9)7g\ZCRPBGR?]d+O[,UE(UD(JS04?_[/7WUb:;=X7>M-fE#-EFdgV,,RY<8
cMD[74H7a;[(KMILgf-(S7POEb>4@_F-5RB(H-\R&U:R2;0Z.[ZGFJ<M2FK9OT#T
SLegd)O:Of.&/S;EDGd_)VFOcTZK][Y4&(R-/@RZ6QF7P9,/e?/>CN7gU[?H;R8F
_TOR)MA?@a++=<BMAD4\GYaS]7dJKUIf-_[YAV3gAXd.ZD&[aHQ+Gb]ZW\57PX/0
W3Xe:I2NXIED<R-)9AJT9bN/Wd_T0R-D^9OYA1IG+7,R7HU90BVEAG=@)>/Y^/8]
4a.^9U&OZ/_>ROPaPH<f)C;G:5X:7;-]SK+G_@OO[J>[K8GQ=O\6SH1/.1Z_.X8G
5@/1@,C+2\e>E3OLEW,;/Z8gFPX>G(NX-[AVDf745J;Z1+[dU0fE-I?@_2TUQZ]1
8+Z1>,gd5VBdc\P.TLY,\=)-@/+KCPECgQEDcPE[FT+0@\PDJN-.d-7)E_WaA4K;
4KP#]Ud+6VB,52,]96F6;)QV:K);Z&,0TZ_99K+9@^LYG,2=66OO>G,@9dE??UGG
cS#1a<C_3A:JZ/V-Jd.#JN&R0a&;95)Fe##::-#0EDD)^]CP2&c?dg?YcG1Sb1[#
c_YR;gc->[E.SRTBVUFR]\I/Q-SCJD9]CCaCY3-(7LDgFYKda-=89,W@ReD0ZP#.
6&d/,6a#1(Z_U1]OTQRV73.AU^HKE=.A&_E9<aXB4@g]eSaSfDP1W9eU:;8)[PB;
V,,;TAYCKPVF&.d0gZRVQOOS:HNJMa#/.=+Y1&P1DY(+^Z&YYe:UEI8D,81A?.g[
Dg8K15:T9c0c))ZM^(^1^ME.CZdcNY?Q>S[@RL1DX>]cWJRY?>^OC^H3e8_E^HR;
R7c>ED.25DF6D&BBQae=.3)T]OGd\Y#<9W/QQGd76-d09feQ4V4LB_=K.]<\7aWR
3A]]MAB.H(S#/KK[-ZUTLA+XN=/:Z4gV)\PCV(V[/3Q8VZ29;.g>-NHXd5\+^[Z,
\SgT:+/^M<BTWZdFc9N88U;.[TKcb#H+V5<&cNJgV+[I4(b>e=:X(DEGW6a][(@P
0f:LO\D+eH[a3.[<DaD]@7c>eMLI@YLSAFKcM^X+0@?fQd044TaZa1E>N5_aHD8g
5EGK0cQaM+SUW)SI]L^+UPWZ1WWO@)LA+Xec8PYR,\ZXP/bN4(ZaH79H<^+]?398
=CMAQ2F.=]cW9UP7]C1A_XH<2[8X>INUK#E31.AVVVDB732W0M<XS9[@3@a7B1<V
/-_3LIE>g03?&LCM#G[cA&?Tg&2-?2#3dA5=#&[WXH_0,.P@660KLDO]O\b_cE<)
K/>,-C4(O(3c^PEXB;>B&(FE#/_DKZL;.N_c8P)<Hd/7I[[WKbWQTXDI;#DT8YS>
UgV+LHH#X[^0,bCJH[d&DC7?^A4NKJ6U&_7G4>=fOMc;^,b0RXYY&Nc#KOP(cCY:
6S003/F)B#XQEXN5]+APG/6Sg^)<<g[SV[,(Lac\S/&VBOg.+8:S@=6FP(_\&6S_
0(8O<666I;b/V5[g\g^I4T2bDI.H)gaYG3X1,.MO7+B[D>13+gNCa:=^6aR4bU;5
^-JPJWD./A+U\RC^\6Df.HIKK&)cOd#YdESH?-2I\9H[f&./Wc#.O[X5+cbgNFP5
[#,)G7(\Jg_COPW:(6=C9BEJ&TC7Bb=dcbEgR=8E++;&?NLdO(aSed/JTAP[3I?X
/E;EL9E-KE,_U2-E4gF#)R43U0GDK8,0dD><6)d-C]H9U_+6d&\3D&-T0bXH@AXW
.HPM_f-4:/:4C9&00YEDg753gFBa=\[,GG6LeF>[L?_8YLV<fZ?c\F8V^X0JDg0S
B(a8L=/TB_0MM]^\.]D@K#@VR0SRGA]<b=cPJ-RCTLKMSa8;X8c5]SF:SFXA^(Y#
_YFQ6QU_CaAPMMRO(d2=a:=@cM3+1/[ZW;C0B426]K_B(A[\E13B^408B#HWKZ^8
;/PF;5fFM4C2LT^(?<M0YgN[/9>^9RJg?5YWRZS8T9UeS#-87,K&:V-1+<DZO97c
4WA?cA>^:>TAJgOA37gK8;CR:28K[f,,A@7+D^?PD=\^KJBdL3Q&&PIb.L^?,TDK
#7Ud5A:f=&HP#&8C^W<bfNG]-G^KcR1^G8)F3Q82a>PSZ140C<NPVM6^1M6L/&N=
#,9^K??C8)<49bHH=5TT4DLU\TV9JUNHc&48gbS/TX1S5N<-UZgDK9K\&c#^bOeR
+=(L;Z7ga;CZWSc0RT<[L;E[OP(J(YJGTNA\+V:U:Pa[K(GMNP(F\:;8[Ka2_[WO
E\.XFcea+5]ZHMU82I1^a.AWa7>,-&a,P>\;=:RZ?fB:1+DfB_04PM&+RP&VY0R>
HBd(gd01SQT3[VHgG#F5VU.D-g55gV4.4W2D[E4+R9Y]_F&T@PKHVdTDD+[QFc<A
a^]eQJ\L-\2;D.S;LGdXUXD,HH82YX-8R.57W#76U:O96C&b]VQK85,b9X0DC6>.
N\02F6-e?A)c=<Jc+G8RcT1?G,I/f1&TTN2fTM-ab9FCF1H3f@O-:gGG#d5QefT]
N4.MAgERT/M>f01)DI_UBU3Z\a:F^Z36\cC.U#TCcS&6,S(\25PNL0JC,,5cS<P_
X0N&I@K96=^bO4a4D,gJVQVQ?FT[PF,1NJO\U?C80>e2V)3/MYU&NV_1MKNB]&1)
@F)7N\1E5R:(=LN343/4^0H0dTX0T]L[:N.CZ9KKBE#O5OcgdDF4JFa^U+8N9^7&
g(&U>.d1(F6^/]?&eN@E=/4X0>^0e)O0=&.31KYJcadc8YB[cWJ^]3QSP1^D&Zd]
CX+bHQW?92G<O>/#AV9>KW?^O(=(RIR[4B>BKe7:7Hcf@;8.S,6Of\DFEANH[#SE
7f]Za.d9=J3;(EEQT8#\Wa6Dd+4;g#5MB&e>YWI7)9/.S=4MM=M>COT4Ob)^de]<
.DgA,@efB(cZ.:>IA0+IV9>e#OHW#J5,894S4\G<G)_&<HHadOTWS^^=[_+UK)<)
VD7HM]2Q^fK<Y0Hb\R\P:>815]8TW?bYS@KN1Id]a?.eHE26G7d]HdCJBH&f32,f
K3R;8cT<?OdTY1[cK(?A,Rc+RAM21Fcd0KYG8Q\,/APXZTb^F^bO0-5)T/4W/^_F
@:b[Q+QYL@0(/.2TdN^VcE_IY4,7de_<e7R27+UbKaZYX(4+8c]d^FPPWC)Y/OG2
F3e5g9&4aR[=a6ga#285>DJbb[A#N6E(P&M>eX(U>cBT3N@RX=g9U([7=eZ(=;0X
QZaYg[cOa/SK?=Fb58egFC8=<1-D;NdHbe4XX(X_[/aR)c^(PaUX/cCTA_0_Q:DN
16#.FXIFXUR=5^T3[4@Ga^E6CL2[K,L(MF(_3?JU5ELR3R)4EZE7d<.[5XY16>/Y
LM&O3GOC#D:))\O\MJ7-P(&?4RL=MK:=f+bWf[fbYI0W;/-/b[F4J#7HAS=<UA,&
+D?.VN^+?NDSC2:6:5#XKf5&Z\RAb@#(VDbS3a)05MRR^ZLSCUB=03]_KD4J_/B5
T;X8L5<F>P0]XA;<F;D3dS7M?W>VS&I-])I^?LV\.:M,+fR,S?Q>DbQWT&+:.aSW
3XbUR<?)L__&?8H1_-C>3:MEgOUfAf)4B>,YQdBD8+\_ZZg>FVVJB,a1S3HV-L[;
J6)7YLW4::RReZTBJY=.?M]AP#,AFDDg6fbe-CJ5[,K>fG]P6Oae.732W/cCD;AC
fH&]dbWR9=87>(K9A)D/64&&\S(80X4f_=IB,K/PC1#4d:eK1I3+=2\FB]3,33D2
;T8Rd?gA=J)dV68f3-],MIFcM9.ET5PIZ5;FGa9[JJNd7b:GLe0f_a&O?Uf3;P:f
CW]34(CXeCPU8=5eB.\T<M,V)bUP;YEY\g1>7N9-S-GR+M2R)>ARf=XIH78/^TTC
e/3>(a4d/+b\@3.V@>.UKKHX9d&#.PGGIQSI\6a2@;McJgIgf4R3S;cQP==a,5/Y
eeOd(AQ?bg(WHQ)E50LC64M;B-28K-CELZ/\)TfCT[[0Q;61RB_&c@>&P^VZZUSD
3N\J3>-&f7WNA?0FAUfIac@L7a/BTXd<;eP#QI<a^_\7@[0C#VQa@IS3?O1O8,\S
>FL-I]GUYKQ^]AHWXaS1CeLC?HGP[=A9Sg_I^(6_6Ud=QOBb1=J/+XLXJa=FS\J-
X#23+a(e<5DXGV[M+/QQG>9V;(0=Q]6aQ1a#6H-Qg_-@6R.?C_-&1KHO7/@4d(>V
aHA-,VcK&/e[<JSX_>WHG&7I9[K+-ULB,_>F\SA>3&.BAc=W8Sg;)PT5J)fdFQY-
#N2Q3bMV@VH?4dHNB]c]D:G)fE<5A)IR7VXVD9cMd>@e6,J@<CM<_K8b;_fPeU)g
1g.^U8Z&BT.O>eYFbg7&W5B<T##97YeRdA?7?WGFfYR-:V+3Pe9KFZgXASA>WKW?
dD?&+2#>K&&f2K@51/]g@]./Tg33ZfB;FM:]ALD4^#8[HUJ3Ba6LKe/NXMA:QV&F
_ZT<4F;7+7,?<JB=72Eb:3#GI5TPe\_;S,B&NSYYN6DV+TZ<D:?:HYg&De4DC/be
f/S)Z0d_a>]^L-aQ2/+7HV5g=QKcEK&ODV]^#_JU599P/]Ifg,@Re;CY3R6BD_PC
MWKBA#OU_YEW)H>O7D+39[//>\Q4-^C=1A1(467J#Y<CF3eQ0VW,<#&AeAfV6N9X
5OFObWU8:64aSD\cMO4,2^64eD/=60#AUL[1K32TgGeaL.F-\(1VD35:FMC7#WDE
G10NBM4-gAKCA8RHFXZ+=))/3D(.f-0P\DZ7L>B\Q9CNK/eP7@:[@9LRD\\UZZT^
9/F\[U+G1-)e3WFIYVaeZCD:-M\)W26.fA>4/6OgEMIaE,A,R#>W2&e&-aIRaFPb
(+XX0eU,38UG#Z)2G.Z\C0BWO\^T,XcZL=f9B7JPSb>O[.YWBQBAaPVSXD2E9JaN
bD8J_(-&2Z7\g>Z+PZ5<U.UET&EQ;M^N8]\ZZAH0GUB_7Q\PU8_0bd6X?>OeOf&^
g;+=7HI,])E@:eL&f]Q6NCNU-aZJ0X9,2F,8M&;cDQ\Ef;DYINU6RG9Tg/(JWDX\
9>LMB1XE^D._ZYIaF^V@0X6BRbCDO2J2bb)g#F[5I?1#D=6;)AS_b-fNM-<&BP[W
]:[a@AH\=EeM=1[6\[>^8b+RV]HK@EC&:ZAc_bIIN5I8LFEf\a\F7efKSODULPC^
U.UfeUTCYX22QRVDTCN[WK3:/Y&Q9++bKI#\_N6HST):IF&NT4La>b<Y(_VPaLf5
c=0A:JR3FA=NOVb?X9ZNL^//1FcIJ)/5YL.\3JcF0Vc>/UGN2PP6953RT2BB)\98
_D),6ca3+/X;Q_N7HZ>B,Za@@_D2WUK^]^JOU?L[>7#;&_fSZ#/&c+59_b[5R/=^
J5J#QQ-X?#/78a_#_;NMJ;NDKF0-4=+H=##47[f1RB>2Ha,)+&I@Q<H]V)B9dQYW
g^S,-U<L:C(Pb_2TKWUc.,.D)0]](#;3#=PU2B88:2EWR.Q86]G\cG)2N@6L=cB9
IHE=D).f,=cXIe:G3EN,_NA:)KN44>e,DO#3KEd_#+A:DNUYGL2/)8D;e2MDE=gL
B8()#\a2N(3^:(D[;A;=?H9A&O=0B(W]0:<-&.+4d4[91Yg2#FX1FG1bO?@FNG#Z
b-eM+AA\#2W#(V#=?>O+[1;0S[C+]HQ<a78QX?ZKH.P_K[N.>b++MGL#^Ab[>5H>
MPQdWVTO<NX_&X1,daP_W?T:S)L_e/CSW8=_SFN]_0I.b)PCL]JN,gVYe@COgJE\
V&L<ca#+UNHO8X;f35@X/7(BFC]F/Z-(:\GH?[3aF4F=OF\<\<E9FEf7WBN=O@Ac
gNdbK@OdS4e)3Eca8\dBeMd7GKD1dTJ.cYC88.K,ONK=f/<M^HaC5JR94EPM4gIZ
_<AFJGN+S4TT+-X;_:@6^D#>9O5[PTQO.B4[MZ\Vfg.Z-gRQJ)QARM5J,1^4/EaJ
&G92DAbN99;,XK<X<a1eJ+LZa@I@-dR0L8?9PS]6aaXGA7[TP=0Uf]J].-29M<)6
aKf.-?CfETQCMTE)e=PXgg]F>E]OY&;2O)1P<9FOUd?<1Z@2fg.98H:Y84RgWPP7
E.>8SbRb&U&-Vb1I-c5:a,V(#?#B)#-#7GXFcWR2_TB2IaQ([>0^0L0Sc1GKC>\Z
9<)/TdARV)D,:4_F(RW9<-<V^ED;:,44FTLg?X2?L>7P3#\;a^;H>R0ES=#8;_b;
[-0O1)VKRZ1=62O#UK^_52>BYgAV6WQ97,cH2.B+?fg60UQbAOQTe\G&XM5LC92H
RbV.P-M4=\4N3G&NH=]NEXgX9G^-&a&/PLV1g<[>&7L]78QZ=Y=NBDHP(CR,C]Sb
gbd58PUB@6WI28G4bd5)ZNK/bA07b8U?>@[PO8)F>[Xg(=R.@5=JR<HM64^.Sa;3
+^2-K>Ga.ZX_U,(PJI/R7@EQ2#?-gOW9Cb+6(\+NO0?H@:gZVOebFA,<:-A:bfWN
RIPC\?^DGN2dT&/&MPe1eE//D+[f)5TR<+<Z0d3Pf^aKNXA^K>cK0[7B_?&5&Cb4
4F=MD;FO?SK<.aC?O68f4dVb@0cC.UH(W+#]--Vf3J6F&e11aa>XF7:.6VKFWMdP
FB84VH/(cW?cH^fQTR5gN4QA?EAe9[2T^b:P&DXc;eJ>3@V>T&MY0>VSGG(E6N>N
96+:5#ZMV-#>A_5]COB0e:=9AW:MD8BL+31N-)AA-;[>-OZTRD6N>O/<3__-ZZ6Z
D9A0.0&4c-#)//5ELJYJTdG3F0Hb;?EaY3DHEHAY:K@_&3FH2.ScQH-NI;B15IN\
4d<_?/:]>5]83SU-/Y_d[gc1\R\[MYU>+(JP2#QXeAQCF_>99<[CDPET]PU/P/:I
KYF8[ed:HgT0cf#(/HX+34:JadJIXbbId=KW6dP889#N]0E&T?a/S^Zb9\6P38e>
^DN@C9H<DBa&XFA<A[M6/3@:>GU,aE#A_,3aO=Y(KU8M&M<@d-P&0a/VJWZS3N@D
Pe5XDOB,1RV[_GE0dSXO4W/&YB_d<&;&JFJ(ZN=4a_>F@S<\Z;X,@6KfgR&S#eNI
U<-b2C&7e0@1L-&F;L9H9VbRUcDI\O)8WUdZG@K(./OCeYOYS-2dGQ9;P_ZURgU]
PfC^-FX8#ZL;PL4/8(7PR^/]-Wf7;Q)?O?INY6^_HSVG7?+;_32ZV0&QCAfH<?\g
@Sc/G1ZD]TN>3&-W.;0Wa5YSU<Y_^/@(]cPO8C\RVFO+Q9?_[daV>[2@#J/D5U=U
/_.)64f38g2>&AFa3U7.C/J(]eQL,&b5gMKTaMGe^-OWP26T[CG]+]AO)>W_]F:G
+-O@S)QU\F8UVcP@<OL/CLeKET-]Da^7UVB<?Jg)9B,=:@=bdJ:Ac4^Y)AXKJ9VE
9Ef(Ge/XH+WW@Ee[H=68:[M.dFAbDaHEdV4^f<AGF1_D)g>dDKBGU4/=LMX,eLIY
^.H(T_d&D9E=\/+fWDgV6?KcaJ&L=-(6(EJ@\R(J]]8Y]X,-.9^G65#_.9-+gf6[
?64dF^Jg&C,[/L07gc3+[.88P4c#d>+&O98O=f1.f/a)#:ddR3X_:,C0+Hg>5O>&
O&@(cK3_+]/DDFN78ULPCce<KfZP;]OXSZWLTFCDS@M1H8>PL9Y@Q<G)T94caN,N
I5Ve<N1VWf^\4ZXa75Y9f-]4K,Zb8>D6@KC^F44[6IB<ff/L_P=D5+WMO;F/4dOd
/e4[Eg]+A0AD/F^1UNZ)PXG87c3D?W2/Q99GGIC)IRQ#=IVdG?7;6.dE,bM+F@+O
ISZB&a0+\/:+?ScZM\RL4C=^YU-4VN8=(&0+_^6.)=3X?;OWTf0Z)3H+Qf[JHfSG
8A,V]HVeZ_(a-T+E81>7+/][bHa?>NHM?c_c3ZJeI\AG11<87.-E06gN7:MAPDH+
??^.QMb#CfY0;f>-5:1b-H.#&WWA36?)X&80U8BZYO)KFc24V?c#H/ZTE^KL4IL-
B=d=b5>5HC_P1(e^2G&B)<.FAggG)TYN9Z7Y>,QC[^HT&])^<Q)M/Q^QS9X>0=-^
=AOSaKV=UFf\bU]OJ-fM=>[RfL(3+RZ7W8I_\2WGd#;(RX[3RW[6@B?M14ULLa3Z
=&X8JC#?:Cac+Eg(PE)006\W&>]6J=e0<_G&I\H>>cZI,d@UeP9^-f++aMfBG-2g
VLcB34#<&4BF[I_0:>9#RJW;<]QA>(?]deKc5c19U@&beZfT-]E2a0bD<a7fG_g8
_WY>NcR2eWcVA14GV6-D7UNVTNC_,UL,DVMRGZNSBb@3)W\fBWI32H:LM62:TR<;
bY41-^<ZNZMYHH=UeaJJ++fD0fM\8)[&AgH[.:Dc9MGdTPL#b+T^LF;OM=Ud@IYK
\(_E[L_&<JCPY(gVF/[Fb0<cE,I;,AR=#4<[[SNHT8FeMY5aX]0#JBB01K,M@M5.
Z/f[dBN]^.FeUL1)LT9(<dX?J/7)76QITea\0/3OcY:-(MgD)T,3c3Ca<SVQf-B)
>+EcVVbUfgVdR=cB\O=>4,5L10I,L)D0,Gc&HT;+P5GeTJ4EI][88/4_E/BE#.>g
V&1Ie4@f)L^KVb;#(8G,af&^Q6-dKJV?RXNO1TfPD\bZ-GN-((NL,>(UW?4d/9aR
&^2B_WUfHG[gCRZK8LK_2\PgO^\&gB+>#DCS^QZ1/>Rg1N0+6\=<aF+ZK>HOZ94M
J3-A]F_TfYLM_4a.^2@P@W@8_KR5>>W8J&@W_@#:g^]>]IZE2M4_g7g4gEV;fP,a
3C+3S).<QKM@>FQbSN,I7A9FS,=:_P(+F95Pe7GZXZ]83^-URKC^;0#+F[9Mb95&
[6XRNF]/K@-V\-c5ZPc9EZ70A9QdR,.C\/C\OKV?K&RN)-dQ[MJ+OC#X58FT_aS<
S3#1G;)4DUW0.5BgZMR3d;(S6,1H:SQUJ<?T/\PTY8WADLEI#FY#Z2<bBd5OJb=d
S&gK,<>NK\2W:c:>7+=]OFMNd-A+RUSO/&9FLP0A:(:C8+\O81ONN&4QGc-^bF_O
-:\#8^?_+a^X,^JaNg5_KAcRMH;D(4VXKTW@-_4UN<d9C0],FUGX#G\/-;TS3^:F
0,1)2;AYJ&B.G8\:DdM(KEN_>AYNQLI1VJ4\cbGGFDc6DM8>?1U0aP,Se3,(:WT4
&;],KNa@?^W+NM=>ZVZ/Kea:UWLJZ8\&^01UF\Y?:W^?L:LZ_b,TWa\/S.WQJ\GX
@]SW3?=fJb.OA]&F>E>./aPA1cN#>WdXV?RV/^_8>S7DYXR+G-R](EGA9\IRaP>]
Qdb//+MZ^7II29IP=R^XHLY3#SX,1S2&>eGM/G:VBXD,QXd=[-4K9S.]G_fFYE3S
5GLV-O8RN@VAVV?bN2QGY@,5GMCU?Y;/+GIN0A4)16&6JX9M&>2[)HJ[>\#H5Fc?
g_D&fdAHeA_&O[[,[)<BHd/.H?cIVV<],&\:+_+/8be>3c.acJ+85C;PR9B7\X-V
eU@,D)F+CAAd.bHdDS1/?K#@B0b:8?4,_)Ue9W_Sa+1cS2J94,0gRbHZeMb2]d+8
R/R))0FI;J68]fGf\2-0NDe6VPZ9#]N)BC3VWGJ<K5:KGf8gCQ)FT:9[f3\=#D:.
S<-+A?\?8)HSG)4,5f4dW:R3P0PT+aSd^,1]d/C;1NE4/A\PG.YcOc(V9C@H02Od
.fbH8-_f)/:<e9cC?_3YF70U1?UMBPb9[-Z8IMA3:/UOJI-3D7UW5-M6QW_eN)PB
3JM;M-HB-KQ[459ZaIAEb&?3=b/)MZ,MW]c\4M2)JZKQJ^0U3dgP?YRP1a)P.Jc5
JL5#aX8G@YDR:J45+ZQH8SGHZ8\ga6/=J<SV,L&V6BeT\g,(feL3)Pb;>\3]gY^3
?0>]]B/R[(RD(&6>QBf66+2VCIfC88GU+RV?PM#__f5.M3R=]=V(B@fIS1K>FK3?
@c>V-US7Cc^C.2gU^Z<6\F>9e6MQ9+GF];P_3;)aD?&_O-GY^R^3WTDYc8P_/JV?
A.0])DRZFK^MOH>X)-HAMUC^=KW5fSLD4V\4+(F)OKETJH8QS?(..>D8e7e\Q3^S
51]B0c16Ug#7-]-c;f/2HX5GfeFN#CVNF-A:6V-5Vd_OH?-_@_^?+&;:YJ[2]HG0
e20]<+M^3NI@AG:U9V7(S0^O1gC^8d><H7W^=+0I9O=4fJ>(Yg\H;K/-?OCb00Y_
.T&).FB(>TdT9>)^I;8_W,:H&4AHE(T#-<M<,?O=ZGR[F,J?de6P]2(.TcO8)KG-
SL+I\N,B>4ES;f;0(HSMO-QM,0URd(S56,-7#;]V84(Y1=[02N#e-M6&YA9N&3TF
?R/62/eED=QUAI8<KSY&V4>]M(#XWTWOOETT2E2cG3K=;IfP].EVW4Y;a?.(K-CS
MFL9&CO;^]Z80bN43VC,7f-e;\^+8+)=O-7#2[-YE<Je1\].+NC=U&TAe&>\NV>D
<W)fK_7E]c/&W85T=X>Q5\L,O&L>DR./)RK[P;HD;3\?S,\SGS6V]WAT<0b9M436
aIU/QR/UNHB];)BCVO[b8;?2X.ZA5G2P\MR-_530+GXJ_>GE[R0/X<UWMRdMfcd>
TYF&[?gNPeDL:]cc4X;@K0\DY_g/^8Ya=-U#3A2W-9LSB6ebLECR^IO@69I->[g9
D(JSR8X.A3<&N/FRG8H?-5G\S2IVK8C)38^JGT_>N)W,/3F;OHA[S59RO7eC#G5U
]Ad,=-X>VV5^E^5QY)GfYRWE.L1Ogf?CV&08N_RV>P9A22/#TKI&\_bJ2)6NK7NT
9DGW7ENI\D^+O9b#/1/Fd-#G9>7Lg>Z09/8MM&T.J+G@,?a^.&9W]S):<9AU8T&4
N)03B.&ea6c<<ec:D^=\4M,D8@P4D.&d?V2IKfWJ]^(W=@\UWGDJfQ(-K1#\A]E&
5U2_).6KA[@12HaEXM.^QSPb/E((f+.E)c9>@1cC,WdZ5#9C5@eeHS569NPC-_3T
N:]b-6abc]F0,QZ8X+MI@ZNQ+1UA]8\G=A]E\L#BI-<J]0&//I:OD,AVLASZ-:5d
NJ6J5Y668V?>BL_Ra/FW9S:LFL^W(:SNKa6Y:8JWJPPD_.41001f0]0W<_d]XZE0
2K85N-KSAT+@N^G7Kb#,cO\#d@cC6Q)^_N#\&X82Vg<dTSPO6&RZ[FcF7@8d@f]_
/>:cR>6+S[TK)-G>IJ=3ecd\=GP6?-X5MUX(E&BKE5B&G<K#,D:Z@:fH3G^2;O7^
,^[P<3_P.RIEVbASBF&C6f5c@Jf35Z[OO/\M7U3?0JbLB^:NcRHY[fYK/;<Z2U<5
1ZPcZ9d]:]gOPU6eDKVgD?/#:,;?T?gC[DY.WI>(IA^DA+.g5EA1XC4A-H(Ub9-2
UK,eaQb>WK3?7=Ff[@;],.,7cD88g5BWb>S.;:fbUU/?HcG]F0N=FaGX]UHE&3_V
L>Y\EBb4/.Y(UJ49f]7b:d6e+KgS[Ug]Oa?D_g^7[/KbM9DTK;<OC4Z+-HFS-TWI
C&L-2]Ne_Ag[B#VG_OW.S2<;-#Q+8cGC.L/X,YBK5Xe<@UCR&e22GLH18=V,d9X^
gCXQa+4V\W^O2MTWD18D,OUCG<LU;RA549N>LPd+Hb.@?de7^LL3-K\8<UT@=5,T
fR2Z1D6N]]g;UMT^J@SC,3B>ea0XaeC_[HMC>EE<W)fH+-Y\ZLI5)M2KM9eC57)I
6eD,E_e&M39S#QA+[GQPVIe?XQeH<WS3@:_DG&:_@4H-Y2]S?A^JfE/g@4UBT_GY
ITO\CWgU-CaF&(JT)006;-dJMLe@#UXQ?OT^7K8/);1N<+9Q>_UJ=N254>=DUXa4
[[R1f,N7@agH^JU7e?BKcO/F[6A^PCg\<O^;R?JY49Y3S()8T4610MT=0>1T?;1<
ZWFXTCV@?F,J08>\a=Z,(d&92)FMd[O?FAf4cNWZCP8d18?M?P>M23+IDHQJ8G-Q
VL6\,B,7@.BCg1=Z_>?HSgZGY8,bWQ>3GZ(+^T.U547g1>?Xc>.^-LOT9W]:+>Af
:cEJD;4TGB;/MU.Q<K98+VX8FNQ;bMc5PM58DNYJS+=fRfcY9DN+cHXD?XIgeGAe
(E/F,/_(CeE,5B6L1#3U#VY0TEbQePUCP(V4d3]>]&:YF(J<T:WO(b025?,1Y\2A
SK_64KN.&fB522g/GEMHcaIE8W=W(\P2e-OdZ<-JEd<F;TA<-SZ8ENfER[cE(fA]
-BS+D11Y&Ab;IM&g8_gYJ<0=UFa2FX-71NOU9d2))NV5@+Ee0[FadPd<:Oa.bR.C
3OR(FSg:_N/-?/)I=\gK21;MK_5-Z1/XY#?K96,]_]2-#[=#IYgN6(C/Qg_(J]:I
_:g<B7]4(NgB_V]1/<2>&+YEPP8d32TK[E)R&?:6)OS4\M(8C7b.,BWeMAJBAX:c
c6KJ]J5/e?,L]G-@0f[X(X)GWZSa+SBeW94Lc],2JER4YC0(a)WPTY?6:I1B0cU7
4EA/_AL&@,g51aWRJI<1f^.C><MW?c^Pa<Wa8EL>KE_3IMg29[4)FRHUWJF1dVU(
;b6G\]U@[JJ6LQI1eU8Y0_Xd=dOc3S3JA4,?=20,6GRT3^e\@-M81ReKO1_22UKe
eY#dg_RgfWZ#TY?Z5[?6&2fKP=d@10@T,4RgNSd;B)1Pd4cfG[d/0bQ>K8;IgS^_
XaR:KZ4;+]M/T@OCRPO#^1TQ_VfI719P5V4T8M]GVKMfK1LOH]SGYe8:9P3)M2V/
A/Fg);2KA8ANcD<_efe#IJS#cOeU;=G+V72YFOR?:OW@/)>2f#?PbYY_1N]I1018
^/V&CE4?(2L#/BN67+X3_;J2O1CCMJf?.gG\E<7aGCWge\XSTMF,5ZPR>(E9YFg]
U3gUQP0e8@D#PWG:daa1eVg;Z9_3L@7dK]():]^aPK,)AD6Be.GQG5cRL_#UMW#V
C91@7Hg[&V@O(bM+U.0I)F]7)C:;c(NQ0T1[\Va_Y#1__BR+O?SfV/3a0fS(7-^+
42/P0RY0].HWRE?=>9FP.<=&U+_fR;0.+ef^T)1F2>WOSbg4:QW&[8&)fMRYb858
3,.,Yc]17]a)?IG[;209TDZ(@2bLF/4#/69]731HI<RQ0H;XW3fJ5B.B2\)Wc/W\
cQ:)\)=V-e\XQJ(cMXH-SP7+U9^K/1OgKTDS#c.EdNI7U-[EPfE3e>#Y8(4a[P7]
5\3L86-F^H40T&+/A^;1Y.@[c&2CG/G.7F4^H#Y,12#4fK\8@3cFd.7TRRa@PO(^
)A52=5O8,Z;3e,:_LQ@MX>22SeM/e2[XI5Ma?WGU&/=P;GGP]gIQ[R&@Q[b/88]]
+D=7X#SFaP8Ib;d9U^gJ?LBO0f^B9<Qb56/#2UTZ3PFc1VQGU_AG#UUd;1/.XU(6
]>(6fIM_#+AOP[_YX+,KWXM?1cRG[O8PME/c9@&,FR(PZ\Tgb:M.=1MS18Q59<9(
+cTR3L]+10)\J,.U96D\_HK/#8[eA=4#CB.N&OI>4LG06AU><b9b:S7?(HQ.MEgK
d1]RgG6V@-U4R9C=eL.gc-:Y=e#ETIR3d)FE/16O635R/.L+7cQ>F<^K=>BV_PcU
13-/Na>L9[CcIT84->a:IJg>[gNWSc+F0BW#KEZ6))H3e8bX\X>Gg\6TGL:9HcdF
4d//4AOO^7LFX;MMXTQ;ALc(@SZNTE.5;97A/Ib5(M?1H92a]J[V/UMJN6Q.YE3D
SA6>LIDb<1Z7LR5>JWFP/EaKZ,,Y2ga.1DSW?4I1TU=gJcRIX9)?(K>d#C(/>\Ub
,_406g0#-VPWc[_@a#GT@0#@@>LE=FSeb#9b1)&dWf^.6(Y7\5CJPL(:#M[GU2]_
eWcK;1754F\Gf9HbbTT+7(KWOXJ_c4Z,=>N,T<V/[Z_bf86-&QK@-\Y[6]7b.>f=
ED.2/5>T]^KZN2L,EMd&1d_=DLd_T24F,37<J=##B-]db,L::#Oe18TDM/d]/Z>&
_DZ>b-eT[WJaU87;M27IgFg4WD/0PFTCK=9_2<>e;O71D<OI,HZ(:+)F[^4TSQdP
O0?,20UJL:)30O\_[/[X2;4O;^;L2A_+)K&,MH0=017ZIeGGHII&F7Je?5ILf]WA
FW8][QE9dSQ&/=g/a>4gMH+5E0B?4C)J5A8U=(RZdQZ&&2XD/:DU/A#B._Z.-:C@
#^B#G4JA1W&>\g+g:I51(=\.3;F<CbgFb>4HQSf>+KaK[bE)6P6g@=36#I[cSR_9
d?ENa>QBWcB[&W6K]5M,Y^K4([?LHH/1XA\bb2R/B]_#?gMC)]#T8@4aA[>M7;HW
9()&J]P-LT]0f?.31Df1/@XD-(Z^4M2,&C5T=HQV;&FQ0BTZ,=0XFB]XW#:2S2+6
ZA3Dc=NBa.FHO2),NgH<\]6L>\QG86S<?HYM@=-P[U>MXYPPTf(&2\)1Me<Nc-Q7
):3@,2FTXE>_KHZM8;DUMAKLb[^Ce(W/AdUKFYF3CN</(R#5(DZ674e?ABU0,^(_
5bM27c8EP5V)T5.DD,dcG93Ca(3(X7S/d7(:6P.G<ZfB@8<OBPdPMba8bRfDE,/c
?721,^DWDH+MD=V?8gJ;?3QeP5Id\Xd5a6,b:8I8R)g]1_,&;)RR6?/R1:1^.PCY
F.U<f459IVc</c6_@S-?0)I?I8RJ6GW;I0(/V]>P]OC^QV;J>^;fUI]=MLN/BgYf
-._ebGN/_Y0_@cG-f\^O2)Q&VeLS3cLfN&&0N2&=Ib6KLB_:CB#?aK)5ZY8@/5;7
\[@Sebf&<,OUY1YHI=3&T1);T,.2#7(DD1/b-ee(A+.QS920/N1[1WL(,X-bZ4IB
@?AEY[D5Ma#F_0-).UQI/[:@e,cSc1[]<UeE+IFR;M^^dfJgMNcEQ,YR+L,\<=HV
[7K]4VU/5H-V(a/INNNSWBd3:f?I7@B)GbQ._#SG@<LbX.EMB[fgabbI#PE=:_a7
4)/d>9N<MX&)IdKJe:>R]WPXc..gCd=;.(_3::W=-1WSES#S9aM0Z8485dUgQLX<
_9P6CZG>)cL^?B46cS;=HcM7N#RN\:D3JYA1eLgN?c+-&>-VQ-6c./[\Kf0\I-Pa
W>Te0gN81SQ^:2[86NY8g(FEA/88J6/@&WD=./9?^RFHgVJT4eB-e_+GG2#3&M#-
6CJ-dHC+R_WEG7^XOOLU1O#2bcAJDc9K/Tg@I84@A(&BQ0&I,I,T,OVH6[/ePG)+
/W-LT/9@KEgEBe/&7(3Q&Q+-D&KgFOIO3ON728V&5;]5;>cULTGf=W&aA=UF1Y1Z
=E+8:1S)1##bL+@C[/.<LO):]fBCgCDAaL[T^L>fXcZZg]@(FJNZ9MBcG\6&T4+a
0<gRG)NZ4I3D&LPHd^H?8eb52edLH3(/#P2+BQT6g+7S7C]PgQ9A-c,/NW1,N:J\
UKa<1#.HF2K_V)C,E@:Nb)ZX,EaKH)/DGKV=MK4bB&)<@2J@V1P(cPD4]LW,bY)F
\H<eQTL.fdYR-7-<g#8g63,RL.[KLVSGZ?4=Z35T.aUeHJZ^+I(<.FXVO7g@d)GR
TV5d?=bZ.L:0_1O?d:)SN<;)6A:&@I5JFcU/g/P<4d22Q<QJ;=7[+RU3OP<V&8Q=
?EUZC&S)U(/OE5>#K;?YJ2fL4HWRA[7SQGC+SfUYY_/=YODc7+/DNHTBNG?a8JdF
8f=0RKXU0F=UG=@BPb[/4GV:F(@ED0+I7E_+MZ/+bB9_S^;5N@QGScd<]fDK7?Q@
6IG(b27\6ZV_#f6?7JLSG+>Keff6)D]DEW.VH#(dS@ZLSOe[?Q;acLcb;G#_KV5B
_7@6:[XNLA<ROJ>M\+I.)a9B0c3N6K^OO1d=EKgY4N?P,;FbH_7QP^ZD1=V5\c?-
/fL+;>X_](&B1Ua\;_QRDC2Xd_\7&2NfT(_FL]+e,5_/\NE8-FKbF7^?=OL-7;QH
JgRB.c^Gb8\9_W2A?K?+Y(TEN8:2ZbeS8P::b6VV=+2;+6H?5M,61fG<:NFReARA
K@?=M&H/ga>40[;PB.4^<\WVfVYU[7B)^97Va?B[&O2LNd27gQ[<[ZYOYHD^]a?2
^ZV[M[6KV][D4aF@EOdJWRL5Z\e_UAf_L81QfQ8QPIdc<<+9<).KQ^&F=:NE_eDP
,#L)NJe,MG;]aabJA65Eg/O@<#a2BPf8[Ed\)IAaTaIASCZ0T4GWfVf#<ZXW-=]E
.[]&4\SJBX+;e==FJb\MID3^GZ_<<V&JT4Zaa5f&9,U^WU3TSWbPfRX.bg2aVVSM
@JI,Eb6caQ(DN#/Fg@<&>/[K4e9eHQPZW])8C=P3I=5#dN4P[7YFB^Mf8@1QJFXC
_BaaF0N[2QLIG)Q(K:3F\adHZ48e1.Rb@U&VHaScIaLc71CSU3@##L#+.UMAS#0R
RH]:(2D?.)a\)U0]9]fdMXND<GGRN310S)F:ZRB_RBXgRBE;HC#e,OKHRY0&/&&:
eHU4VG@E;CJS-7AY8(]b,a<4\[bQ4S9@NJ>]Qg;_VGgbN;DGK](6gOeGARSA26Ra
0B[;;\ST>-DOKYdS@/@19L/)Y&;OI<_OdCZE@PONDOXA0gY1#Y&I:P+C>AUY]FH0
7GR41dGg/4D?,fd@O8g?@FBb\H.b.<_S+T\FDV51:1fIZ^ebH[6LYK5-8fg]JAQg
a0EbfCO:^_#(DA&_;E:0>cXADAIaRSe?X+V#+AceA1C+0N]g)?F8Q_<?H+>-F07g
ZP/a-SKS@Q49F9C0-7\,XZ47KT9C\Q#:Y6\6EOW-gb8/T(Z>#;:&&:#VJVI)d>>@
X_Y7T>)XU=9?+5V]]+@@[<c)=X(JfNB)G.Q4Y#e>^S32\,:]4=3dd_fL5#H.++2S
X]T[Q)CW6dF>WNU]W/[a)-P4Wc,@V/.SD;aQ=[>F<GS=S7Vd[4>U\_86+=<+-.a\
5HO-R06VA-]HAM\_)T:40.5EeWD=P)L_IDd^)5L:7CO<D(J@_dM8:/XK<^@K3Kc5
2\310CE5CI)\JW5B6LagNRC5[Z8FS]O_YM-9O]>cK6V1P.6<TWSUJW1Qd]TNBIX[
=/E[WOW64>He6g-@=f+VFE1JX:MTf=)EcBBCAc/&FNW^9A=2/LA.\/ZR<(=2H^?B
.ZW.R-;,MQ,#7aD6(NLf<8M8J25,N/XW0Q&FXYCffV_:^@gUb,HaB]WK7VJeLKS1
9P+aG&S#)OKY]7F;X?XYMX0Y)bY6/\3g/_Y>/:+Z2(cKBM7d+beGS;9,6H]WR;]d
7FNRQIQfT\Qc6:RG_L>0/_9Ef2CfUX=C)[6.NGS#DaO)QALBJ40F,[,9F>0H9A\X
eC>7J8+E;W=6;a/H8@N[49[P+):[+\NQAaNfHG45.M8AJW.].b^7#DN<X,PL-7P:
BY4e?CG2g.[FTGag7@>Ef:>_2e\b(\R@6:3[/2L?^TG]RROg;F/9GMZeBY[H:PaM
:dPe:T)fa2<HIEXf(=JB#[1[g#Ac:WK9IgN_[E8g63VH^WA7U-[,Y3;N&/Q,a/2_
)\O;58N8S\,^)@S,4-F6bLV)D-\WVN?:@V&E,YN=KGHa?Hgc4.]CW=+]0?Id0ZNX
M8UaO=>FV.ME[K7U6B@0R)4+J2P6a7d.SQOf_UX5\AKN?O59/cbAN<#JYUAH(ULO
VXY>6@c@X\B/OAPIJTE^/E7FUdO)J]EW+],=<EDH+c8ISN@)Gcd)+?#SDbMN?5bV
G#RD2a9=+@QTF^5a2([.&&EZI6;3D+5=TDa[#Bb#Ig+3+2K+_Za6?TcKg1(_6I&=
gbc[daC,85XW[Q>0G-\e1M;cEK8NVB9<C<<cO_//5\gg\XU@29@CX@KW7W??6M/J
-F&D+8N0N5/PL:McBAGAK,&F(C)c=?FdaE+MG6ZQ=HU_KeV#5Gd9HV\E,QL<4e6U
#YH<E)YK/MT8QN_<\:cRL.F^](NI6DGc?4JM_IEDAQBEPR8[8D92;WaU,?#+&SUH
(+f-JNa_NDVSc;)Y<f#P>f90B-PUCVH]Ed[9[]64:<eG-Ke)UU:L6;)K]+-E1a.e
>X<9-7HH_ZOLU&4=IAC45@(M:(\@[L0)cdA:4V_YIU;64&4^?Ja;&8O>,KVMS\d_
dG61;+3b-J34:IHYCIIW095BJ/_eK)S/BFI]U3TBD9^VV^3IgM<F[\L]-/M1)DgU
OW_.;\)^94/\ce,f1a1L>f3XG\10[U:?bcdZSCT;WQg<CP4V>QGE3SM@PS0d2#4W
f3:\UN,OPg9S-V;Z5?Dbad>Y,W^DXUV-X=GCPEG2>09,&,=F&gdHfb=VJ293Sd?4
9SUBMc.11R_V1CDa]92V,GG8-+DcUIPZg=087]He0)]OO990/dac<9SEQeHL<J4_
4QH&7STJTK#1^Z&OR[>BF5eK=L1Y/MYM#UN>7AL1S<U2KG#.C&)?T88GNTIOgOTB
Q12/L#WN,6UGV5^6X]J-PAaWFLQ-F(?NL=EEbUK6\P8<LAU2Se\HB.CG(8e9I[CS
,,S]JeT9XZAX[P^,[T@=,2M=L)X>Cf9ES1,7O5e1#B=HO@YK+2S@VbNMPF8b)KA+
N:&OdQ@Q(Y,N2UAKEX0\:eYO<1RK&3CeAa>X1c+7PCgW:aa8#8;6MHbZ#/8_Pf(W
3Tg.d;A-_c/f:&8IQEYJV#50@[>=G.FE<ABKMYc:-R@F[/QFEYJ:gZJZ5[[1:=4[
N0D,^MgaS]6)KJ_dZ14JEGNY-:::0#F4ZQ>/W5@/3,X<,,QgELQE8(TXW@6+fc:.
5AUC^X3C]O3.Ad?DU(ReXD=2[8R]R)Q=]5ZF_adeKE1GW3K\gFP:g32bPSNZJa=Z
dLDM&7c\\HJ@NY9-We^?>(D#0H\7N].=@243W>2TC.agIT4/HH=#KbB1#UZ-PZ:L
f[ER9+P,=>f]06]7UK63PVNH>1CV>0=\Y&(BZN..CR70Qe4KYP1/B8U+53J#6@aK
&S+ZM9YCR<^T@??);AfV\e5;^W->6&TXOM42#:]##3DM?DLabF_YEQaA4@]T-HJ<
@bR5+ecL);ge8+I-M2ULV2K3J;Kg#E=bKD>bH5,(>X>UBLe8@WLW77fQ5LG]UdCU
g56=cDV<OTg)MCEfc3QQ-4,/LcbOK03C]B+aaf1UM^DP?[.=fgDf2U8#W7gR2)NV
14L4gZ35PCUJVYXa-dbfSYZAOe&]DAI,SQ28^?E3d2<XB9@4@4&E@6+B3E>TMSbN
4b&MXGAN[Z,\c-\[\K/A.:[Neb:_I1)geU8^0f=/.BAe_I7ZA-gQ4R:JgZ^#,ceF
P]@M?aRR_2_VePL3-D;1bT&RX>K2Cc6T^BRW1FG;(g/M<K?WGK5(34L07<>F@66:
=#?TME^=IQ)G18:@N4AU[]c3b+H04Q_)3COFeg+>/Dfg5G[(\H1NCdOgDd7]cbP0
2SZ27?A<L#/P,g6:KO&#JHJ(GKVVK_LW8e@<@W3Z_WK7IXRG/f14)+8.8;S30B@[
Vdf\a&JgUd3T;NCUZf_BT,:S:4DeS6.BI1;7O0;]@\Z[fREP#bD?A65(c[MXEJB4
4-#>KOK_[-.4&7F/>TQN8f<NZTGI_CH0\bH8]>C8=-ULT9.]T\CC9LRBgA+JX/5:
N+a#UQc6Y<Qf^C;MH=F@?a2+/91d_Z>\4_LQ#]O<(gC,.OZ:C0+ZM09W#ZPcAL\Z
U?2Z#,B@CF][L#eM\^,O;&>9bEF4G0DG?XB1bCI2(4,TeR@7UFHH,gE.F7Vd:Y+6
#335H[7:d.#LFZ2ROe=1-2P&,@F/ca^UX0:BT6<&):2GI#P+d3@RBaV2,;gFd?K_
SOS38KYU36LW9_JZb7=_gECSL/60[04TMC+g_CbF5S69MdVD[M?/6<KV[@9;X)Md
fEX@b@7Z([V9@eR_BW1@+QX^e<>Qg.U3HWT:PAD<EVb9-,5@>gf-FGYaX=04ad^[
IN,.N9]b[a0.YXJeTVJd:OI;V.f==c.eNf<30L].WPb?>+_^BD-CT2]UNQFP+OD3
SDZF)YA7=73JdE2F1ZUY9YLM1b70L-3ZT=2OV5\3S^+(dc0bEQV#@)T_Q1;8?X1J
^XKg,57-c^UV^c1f;7;@1MAAZWc-??F8P]]a-:cHc6fZ#?R(_^FXaaZL?c<(7egS
aZ#D8):2,feNI=e#_T-TDC,5eY#e,GC/eAbe(@<EC&e4R-)]Q-C)JMOXEAE^g=W+
:XYKHNIA9I&[DfD]=6?bJe1XVBTZ8G&\#eE#@VLI6(Q41+6E>PW2/J36A20CE+LX
<YSO5-eZZ<eXX7\W-KV0Vg\bVI>U8]?DBF^?1(FZDbFDeNKIcH.6d,_c;HLWS-5B
,FgL6\.]63)S0N,;8cCQ>[V7bdWVH32=T..7K29Q(J4da3cY5d@VaT0LBN/72>)a
H/7S8\.R+<UJ+<2V=&Bb;\11<eeU1/5KD:a<69[0DaJ&>#Y-0)MSF&d84T.3[W7\
e(<(SXQRDb[[G?PX.Xf:I\<T[V;PW5.?X_AC6L<MGYIML3G0D5;+<&)1Ga+g]f5<
a:C9H6?P?[Z;)\c?JVSV\@e:c6cL0b/5eOd93I-2]aCB-EO]:G/,=O&b^DI5:I#:
c@;N/HZe+]2QJF^=1[/E;<GH2BcF_f:HI6^ageU&ZNGO[=@FWPZTT?)LW9-BVB+c
Q]RD4R2AW^=.&OY(A1ICdIf=,/Y8RG+b/T/@:V)QD2MVFULXY8:##X+@9=U7(B0(
NagQ9OR+S&+=5]5(FNNIF7d;FCNZ,\M<9\#H-\.7__dI_EaV-H0U<_<#gUNRR\EB
0ZFV7,?YW\^[-MT+6N2GL]O69c,\,7-E;SaYZ=e&Pf8NA:7-Ng:KgX:^OE+7\EaP
UJa#,[Qa@U,X@R.6KF]d9eDbSFZZe/ZBNX5[KDX//=T/aVBR#+FeN9a^)f)K<>#3
BFHRC\b=/c]dAd?W6IGM=1S9]2I.U8(D\[KTH43W0Q/)4:7BbI96I7be\T+:@DX3
4QX6J4F)5:3\bE)a[>+b=4D9;S=&dUHQOL\=6N&CP^;HH,RU[caabb_06C#)fg1;
JIJ@HBEI\J\L;ge+f;YAH>E^9d1J.e2;/g22R\#c4R#JX#f]D=<_5RJ6.b-Q^a]?
fRIEE76B:>X/_EP;Q?Q[]^[O4J3B/Fb#ggTW#:)576\4,R0SB/FNeOUMXPRC/Q^<
B.QFEA.Ta5&EA>JZ74JH50K09KV^<MTM1K]))WYL:Ne;_;(E6]1DE5W33.G?[<@N
.P]T,.^:B@JF>[H_BDK>2d3cdL#:8gbL.aG9eA[2_-<d]c)W&B:V4:]WDa0&2A&H
3K(738)/<bA[[L5UCO:FBBggARa0b7NYeR85V^ZeK2d[:@[T(@N)^WdV<=c]XEWX
H]@BS<0\K\SW?2FGFA#WPd/6#=.M8Z+<S;GROYQRYU^<EaP+5T=1MG(+F1>LbDHP
4)W>?6LfE^b--VVd-B6aE(Wd7G^[O<,NW&?H4A-dg^&VcdL/&-\WV&<C)+KG@S)P
CC/4L=:S;[Z?]=#=CI2GUL/S^b6/H)?dV@/,F[L:].-[N/_Gc)3J1d)FEgGCLNVG
@Y@ZSU/dB6>J8gU@89/\(2fOWV6PJ/d6WSH<dUXaU@S#Le/Z/HD/W<;+#DZA6G5T
OX4;@+8+1D^N7N22.5,af3fd==(KVCJ5-2:-:?Ia<4.R]\\4<R6[WYNLAaJ1R7\X
G<K>SaZ:+_&JJ_ME28)f>De,eLK_<=7Od,E+Qd/@LbZbPR=83]bW,.DV_Wb&Q&c1
>Z+#G?[.E,IGUgHT_S5E?:NXH[V2QS5/=dc5P/Xg8dd9UTcQ+P=@1a(,.08FM>DK
L6+QC;S/RJT/C\;?aVHBUL#J)/]Yb@&]KIFL/YKV(-XC>.6A]bVVS)UQ)c/?:dgU
LCKHA;/0L<F@)1E)N0OH&2HMg3Udba>.fUYcXb:<P3J@?MZ)0PK<Of0.(/S:gOU^
Z<g]FN-YP2;=]U8RH2KLQX1bVK\Ad>W5aM85;LY055(-D[+0R4=D9a,YCeR=ORX6
@P\WP]PNS>dDS70:O@Iba,/b17GF1XS<3Zb5Ifg_=^Q\X>F7.EZPP=32Ya^<IDVB
.S,F8)b:9EXZ-E2gLB4WHGPUdR\1W8+PGCd[\240bXI8W(4^K7H7=9:_/J,F8Cc:
#M7c]#JP__cI,5b5[916CPd8B#Y\0-eJ:ZTU:U3KG,A>?\HPUI_&)M2\D7a/>&fB
<QCRL26#AX2gb#1<4EQ-YbHC&F0f[1T,</-^c9C^(X\17_H]WQFW4)7d510Y9b.\
YMOH0C4HM>MC?>-&BCFS/<?GIS?Mef+=GdN[Q0&f?IQPJU\W\,O?&_,:6Zb3WJ+;
BUK#C4.XPNGS9.E3:e7RR97B)_2?D8@(67[^U:DX.NbdE3\,GadGA)JTOC34F.8Y
2?77:KAM/.+U0FLXH7NOg^AeM9L&;E8T_8=MQJ,;:/]8,d5FI(SROH)PQ^J5O_&/
JT-bfD&ATU1X#FD>]cJF=1OV3fQeaS(Y=,e8--V6cJgcaT+D8T##/5Sc+BXbR8WR
E4JR1-N391_L+?52O1aQWWNf&5/BB^1a:_)fBVOBg0X-^)b[IMGYAW/C\;+<f9[_
(F@6(g9,>K2;-,SMWZdb1-EBJ6-3420Z3MOBJ9d3(=NV,bQP_3]P^0UC?O:Z9K1P
\/+8E&e16gR3dS.1Z9N<0@X[B=-RJCEI6A[6^@6#30&<OVGe;,L5DSSY01[(N+TB
]De@a6W369WR>4I67bZVeHg>]M>c/Hbg]1W/F5:;_VK&C_O8@b+DafT:_[Cb+5;T
].f3(=(+?2[b0M:L7R0?JN05,IV?ED1\1-4AXa2/5Kb8[MfU56KTdbSd3Y4?LYc)
DXRAJ]O1Z(3KDD4[DeUM8&SL0e3PL#/7B@bA1SUSA+ZJJ66IcF&8)P))WZFZ#Sd4
-e-SPN;bTP8V3NMP&f<PB\44L[8_-10D89FRJP4(3e,3\b_?6P8N_84#BR0a)2<f
?&H9fFCANZNW@faLaNGSfEF:W>#=)UJ0.^#V&TW]fOBA7>X)XcHM=g-d?-Ug1QJZ
LF,QD([<MEgCIM)C?NCYEYWFfZ1@SPOOTSBHUC[g&X<?Z1L7:e1[EMO_E)OE:&>I
HLQY/QeAe^PN[EZ=O7ePD.JSI&>Z\I<BB;V+21c7P1;GZ9##0:X1:D2P?8X4b,ea
?Q_c#Td[8CRUT/4WZZcb>_beL#2EL.L(H7a1EJ.3a:8/LN[dR.D11&D?HbeS38B8
90)5(T1a+:2CFM\,8C#Va/ga@19B7Dd?[J)XSVdc^R+WB^N[ad4:>gDGL&,Y/V&c
bN4VK1;^;+\#+7\K-\70(-B=/>M&OWNGePBB,AfQI#G4;5,9Ac(Y+_RACc_TPTQ7
K4EX8[4^Y]Aa]F7e[^f)?I:NH2NX3Q>a)II]:LeHHGAEA#Bdg#2PMgSLN5OaX]8^
9J<#;OATV7;1&(ZV<NcgGYI0//M#c.FOgY\1#@U#ef+W&:UV[:X?eCE86Z5dFDad
@=08T\<dReCLd)&a@;X;RI<MAAM)W9S8V.gM7c8QEW&\GK<)63Mf4cD6JEX?V82J
U_WK4RcZ^_g2O_0P>#U_2,)afFHBSLeJ/NC;YQ:RSJ?5agTT8;86.W>-__(4M\@7
6EUPf:/<=PNW)-Z843&;_DTW#g9c[F_#0OeGZ0;4VFa#U(a[f_K0_U_GA3c?:bb<
DM.:Y4adO;37,5fVV<QN60I,P.4cCcC-[Vgc-a(>EaQ7Z:f:LD.DECYI[?g10D<:
G\Y5@Mg]0J?UeE6[ZL^?/PX7)/-]>8P?SO<4b[_</I<#Le:.W.S/)T/BLH5@//4>
]VQ>V?1&5D?=]\Q<E<a<c08P9D@.0Ce0ZKbW8Xb==BRC@GDQ4#5XBcf::B,NCe=Z
CV,bYcI(c=(f@cP7e3J+Had,C]82=-3Y(^@cf1#QN))=69))&U51P/QG]YT@LGV(
gNbOGg6SeHQ80f?S9+7?(BdL::7\d@1X_-,+>//,JcR1LTHBV65WO:2EA<C)WTCG
YG9]2Of.<bUF-O5(]>W(0L1Ub(_+[<Z@@fA+FUF]T24EICRP4b-eP+7A3?G05^Y2
[#BM?6A;U7M+)>c:eA82SZH^I\3b>A9XD-0(&:6D1QfTKV&a.VPEZQBeEJcX@PP+
8)aO?_=XMDVUfaVP+4a4#,+C^TX)TI,RgAD]1DaZPg\87,&70_#GFG.[XJ4JG5D<
DcXf67?/C?b[NgecH0+0Mf:9K]C7HT/6?:JX47F1MQb1aQ?457]ZM-eLRg@U]I92
7VYfEJfQG,+bQW?.T];QEOf05V&->K563Fa>Z+VJ:878/e&>S9]:Q65MU>4_5.H_
FGO)<OMR<H3BDWW:.FbPMJgQWB::[E3=HH>P.3NK&RAOVM5C#A;WKA\IYVQ8V+gG
@eT;+GegR=9^B(&_2\::#)+_8:EA]9ZXgc1)1ZB)1U\-Qc&D8EOL5&U5W:/-):N5
>/.a<U9<cGQ\6;PZ+,0/#G2Ae++86g@Ab8BfL^a)a]fZ&0(^&e:,[.Md]SNTM-]X
9[e/aeE8FWQ@ZT.>F3.6B0FaaR>+_E0V<+^?4PH-WD7=+2VZ8Pe(\]D3:_9VVJa2
W(U9:a8GX;]?_<94@0,N)5cc>c^\>QGK2eBSP@C9T7IEW)8F2649UHgf#WfgSOfR
fd90&f<G8UE]7LLf3c#fQ##6E\RT6&+bVS;L+]F,]@ZR&Z+f-dLOJ3U+_HF.\[B@
[egO<G;d\baL<CS2gA5=,cROKdF(G>]9RLMQ>0Ib=d)O=6]YUObU[a-/W+,IdVLc
N>P1&LMH2deQ6KGJ-F=Y_77DTWF]b=P>#aeSEAAG>B=.QO7<J7Y[32BK&=QH(Y.Y
,\=Ve+J#SO80?)C><]E67].5dVU.TR&WG84_S,,gf=(?:McD#3<[6d#]7(5UCDT2
_b]^(P.)\a]TC#N06-)59ZaX,G0]d3b3#T6W]XD+QU^JR9a6-/?Lg=dF3?H+MEB3
^0TE\Jb2905_d]ZC?A,KN9G6g:[ZS8/,BPL?Eg>WR#)#6)H?6WY&NfAV(J3EHYD.
TQN[.[UY6_D@NVQb0)EU-W@LdR<.&BIJ\CD>0c-#eGOV;0Mc@687)=K4E@:X#g&/
OSQ82<c=LIHF(]^&,6TEE=bMTKV+IBXTa#:fQ]S+_FQC5fD5g/)82fCb_UC6L&,/
a_T?9BXZdZ(dVd^NK:LIRO;VFKP4T#M2/=AdSGB([B0KXBg3AW@KL^E&V&+1T:b;
<OQ&VDZF.-@@,OL=V]YS,gXH-+fH.=GZ\a4g&JeD[6Xf.OKRDd5AIgDCGO5(D,A#
RN0LZIK=GO<=?^IXJ,TR&#fZX-J,IgPb1b(_9R<d0,#98]K5YbR(=;]c+KBgcZK0
N@Q;/(Xe8N?]L81bPO)AL^QO,KJWd(+-&E=<6<34\X^FEcI43:0^\10QG5W3SO54
1)J5N1WJJ>W@/]6HRVHe-KZS/SMRC,,AHgB:OL\S^[DOH]))@Mb0B_g&X<\UHH+H
Cg8MJ.:\EZV4S=Q2e=84,bP>,_eVFPF;GPf8>JGQ_+?S332B1KU(>++;;Q?.TX:G
LZ>0X3JA1G@S9DNSA9F:QLA7I&/E#73>Q((,65e>I0(.TXP)?&B\YeCg;:,+-L?S
&[_D5X7QWGaGRFCZ,b9O#ONDOTB3,IAL78_3SU6OU[:37JX>PVF]EBU[Y8+QR5M(
95^G2;MPE;#EQ/8MW+ZD,3.[OH?^KfDCSe5I]A+b]E.&:--2J1NXX@EY:7X(e&\L
A2RaUd8cQ\L.UEL2EH:X/EN[^eJ:;fCCH>?BgaR8CQD[5X97H_W>4=<MHBXdQe\V
b/5fDI+0K[:P^YfPE.b-1Q2g&/3;VUKcU1<X&PENP0HgGVQ6FZ]S1_@=U_-\1^5U
ZO[M###KTJFe(E4DE9@^C+Z]^Je^N#gKNcBF<+?U]HQeVNCfJXIMZ@N6.4NOJ709
?5QWBcX/OXZUO^#0c7GE373<D9P/]6W\+&LN=W@7U&K20(c440)YBS>,^f#6CU<_
NBCM(U26gC4GG^=3U9C)SQW0]I-G),dR>1-X/LJL0)@3./=WZHKV@8;OS,I5)fL]
BM7[A+7?VV<+>7>^X_=K9XNNRNDKE/L^_X:^bN?BDTF]&B\dDW\c#237<#PGSIQ+
F[Ve;&7;&1+/_^&0LG9S)MB31]EL_J0eGI;I_>&2.U=/YACe1Je[G1T.Y.JF+3)Z
2RXXAg&3D@I(f.:,c;FScKK^N]DDR#,[42gANdf5)AeOX:Bb@;RVX7U-,]S+JD-Z
.T)5@6<#_NT\H4a6LM#C#,:52OI^f=Pe?5<Y)1,8D1^.FAa@I1WH<+E)fdX9g7XG
>^2N8.1&cFRaeA?NXWL;7(L;K>9\-96C-FV)4(-X^HSe1(Xb1E/&R@dYYU]a3^\/
gd9,&Q0_Z7IFbYZBV#TRPFa_OYCIZA4]HKPVJ@\QNXERT=C0S_)=1784E:8Z4ZY<
c.=H:O.GDD44:F@YBbBQPaBe=NBd@RZ?If.+a5NKE]CNPJ5N[&TN98Fa>eaD<Pg2
;18EXY8@60HU:IU=L_L^]&gB<5AD7/S_05L=SCDd_#/?[P9[G@(-G,Y_>U-X3.JK
M.YI@C,RHId^?1JF-d-6+3,311\6H5OgYF7cG4a(/GeWW&84aP27,NIdEQ/dI:?9
PQdAO(=,cefJ#@[XW^H(?N8H?:b99<-MLIce@R-Z8J7OdMP_B>13\4-JAXgREIg>
RH&03JSJ+TY(eg8TVU.L965Z[YWFYNL1U&_74b<G3Cb2IO&;bgTQgQ6-3)PaWX--
BA+fR92:#e4&/J?H/F&^;=/I;4Y.OO?b?#:174TFOdTTZH@_]8J3ccE&RVF)4JHZ
JI:Q?g?aA:_/]M?E]T0We]C<W=2,Te)<K44eR<(0VdN2^CYUKSLe)6d9>[[0VP;3
KIWP@<:-+&(7Z_X)e6Na/.OSC=N39PJZB4>,)H6#<Gg4/;0a3:ge-\\CW#1K(c>8
^G;M-1b?CBBR+=>0cE7](DS]dV2DB^MLCbL.1X3RaYE:]^_73,?f5WAEYC=Z1fUV
=\cFN.WKGV[g0[./[g>dY[P)^[9gJE)=;QY&;FXbg/bE.c>a6&GPZaB444))/Q@,
2)3]^?\^N>,7UD=.M7._4?CZI)XY2LBb.b<8aC-be7e960deZ_A-CR15M>0G;<d:
OAM-XH,K1d\J5L:@RT/E<L1]ITDaJ(Ed^?ZIRZ>=#YKL>4D-8AD;b0\RC__f2_8L
NeTa8Z03f)P#.g37P]F4USOELR]L.@K2L+LDC\F=4-#e)MNT1e&U,9S3,[a@4Z5\
]a)#Q[7W8U.\7aFX3.(#b@/b\+2F1cR?P)(3I,DJ2/f;C;]Y[QS=MT+LWTV]8T#E
K\1;QX?SEHEcJ59QdS,76Q77a]AM3]C<>V+T-_HE8Y-;aM^#RE<7QTG[Z5[CO^Q6
)&-<W63B-PcB<DV=W&N(X98BC>]f@R.YV4<J_=F/B[aS7)T94B>[C[^WMEMUEIKg
F5RTF/0(^cHJMO+P\AROLZ)Q<)e^\BSBefMPD_:&>G7aDF:&>032@]^EIKdN#D,B
)G^4IGQY9QD^6??YI:aAJ<&+IB4P#^^:XQV(NYR0&YD?>&@OW]F&ZYf/J:33A<AD
1Oaf.a:(bEBSA,)-M8OOfUg1R_\8&:Cb>Dc@Ic1U1#9;^K0]f7T=V;9S_F[0CJQ-
;S9>;348Z<OIP(ZH0OHWRa=9a4LI^_L-BKe,VW#5NBZbD_REK?]2A(=.<U4<e(8T
PRNb[]--Z\GUR#)QDXC9\6S(@+,b,]BDfZ[VJ+R#0\Hg9NE,[Ag:gZ3K\X>,9&ba
S+cYcDgQ.5&@c.M0SY,\f3a3b1^@2d5A2T\gZB1b#4QK7T4GPf:Sb+gK;M5:gX/)
13S2aNW_1H[.)O:aWJ622[99PbE-R4S5+/I@d>GT1Oge+V/5E,4d<5+DD40(Wc\#
S6IOR+X4P6LTXeJGd@R.0=2eKMf[(gX43/IKg&/55\1D4B@=8f:6<T@?R>9Lc;1X
:&C:RICf.\>b0V12Cc7bb3dWIT:KcJ<)Q;,Fb[.92V.AeWI^fCBC,O?6#YIP.@=B
KY5Gg\PO+;//]]DP^e])\0=_&4@d(f;.:B4:H56:HE+)&6gX;)7T:-WR6P>/5.N/
R&_CgfP&W4522\;V/]VE77>J/QAC]8fML(MGRd<CX9e;C/L)6B4-6EAIFEX7OH/^
8</;7AKSAXVX?DMEQ[W&E/MZeDd(<ZfbNge4W<[7BWN76:QFc^]#0GWDP7=H)#@D
VR=?6#f5H#Ec4KD^C.S89X&M&,+U1L]eRQNEHSd:,cJ-.QUbAR4TJ9de+8#W0e])
36X]X)Q36ACQaR&BC8:#4=CH<RL2dFY8-9OcXNaJP2Zf8IPL]b6;HNRTBZcY[G\R
7EH]30XPV#<\aTa?_Ve\)g3QK&E1(B=92Y,G+C?TeD83\dXAJZ1;D]0@P,@+X[#9
&4A&I?IH?V:7H#KcL=(2Q#I.EYd476_]A[LR14T^ade.0Db\GS5W8#BdB5Y.G>)c
?fP^11#C:<G>7N47+Gd(>N1NRf?d1HHL@(4Af,NIFdK6UbKRS\>bA,E=P21&]f#+
.HOgNGCW958JcNI^^MC3-Dg/aFE.-?+D^/XD1-I_-8DaR):?/F<5&LZE-8,,];1R
D#:O<=P5K)KVNA4/6\6<42H/2QYYH5b13R9):3,XZD7.._^?[bE):-@&<A2Jb+7A
,UL9TX#L;]=@>ZdU5QaMc9cg.ed03G[:B,-S=S-O=<(gfg8.[.(X/Xd8e[W,L1e+
KYd-Dc4=@eQ-Aecb)e=G(+XL9V+9[G\d:4.#Oc:\[JcR<e[+gJ8(?X/QL=[66Jcg
c^gX@VH6>5.g_AV/UdW>K+)EO933-g^eWb8,aIV?T&LAPMa[AB=F,#@_+UBQ=f.L
KY>K1,]c:9>?SA7ZQX_U#@RXR:#X.+dK+>_Q(F@G7K+87:V&9VBZ#0E7\@+<5@EJ
;5e?,1J3aS59OJVWB55e:?=A,>ZEAI3\9U&0?_0-,5Z4\#F8Pe#U]MdD/;)#GH6R
O=aeR-8O).^]_,@]B643]?VB/gTeO53?L(XL(_eaXeP(8dc1g<&4^CBM[D/fb,ba
Q\aT]V7aJ@R&4G]A)<WW.ZRG.]8:bN17,JZ?(.]-Q=XH6/\gJVBJg.WNeFA-LQeL
8PRGL(\a18RGJNUXR51)e4F,-MTU\L/9=MOV<D-[d8UR6cfOS=UN2:7]F-Qg0I<R
4T2N:)U68:WAeN_5:)4B7X.Q,b3NHcaR92&YM.86)1N=?cd5\+Vc5bOPP^7]aY.A
;PC<L9Z(V/9?Z;=]@1C_^&N/H5SSFH#RDWA_6=I.E>;I+W8[\d4O(BJ\_eg?96g-
4g_eI_5B&e+]g^ZY_DEE;gKAM/MFEENG/7OS05&K]ObE88JPRE,8;3U+g6U7f&F.
FVS6f8X>U9e.CK[Q^O1:8ae7I78YP&OOK/;;?Z?VNO9_E^]WSP[JG<V9[81@=[DV
X(_+;I(?N\NG<XaDfO1VXL^0^+?:J4UYYLI5e]/2.a9gg7.TAQNU8LCTe]TfO]O]
I7Q&]c@)D\US&68\Fa&C879D3fM]cD<>8ZTLgSR^N8c&W^S#CfG2P:<:f<UNc#P=
c8&XMYHB)9ZR;N.Q6Ke@/)2J,\+MS54C2)03O6H9>2_0Z@N=JHNaWO<318.WGB@8
E2ABI8)H/17[O3RX4T,0)]?2PTJZTUYR(.H?ZO9;)WQ?89eb]UI:;]]R]&0\Zc12
^LFRHY1+9\H^dSSB#ZJ2,N\AC4[/45MDe4G]eQA84O+8+\9@I#WXF(M1]-#Eb0=g
P,2E(MB(T2@fUa\@)g>,87&8\#E/-fQQXKRCD<+G+ddbA^8=#RK_g?VI(XUR+ZGS
;c-N<[g#gX7^W9@(g#/3\1.V)D4ZK;C#RZScbKYR)]bd0B,4fI5Tc&F7_\8YfT>?
#T>O==(d/a<1F^9@9/3IeS>0-)ga_fd9,TdEX[X)@@^ZV@+0@W-:[^;-Ff8SHT71
1C+Vf^Y<\KV?YFbF#c,/7KRL\#@9[OQOXM2[+Q)@0d76RQ]fPI@3;<5^5)S7K_>5
3GWC+6HF.]=P(4V7SCHO3VV^6,9_KOL.GGg=JVeJFJ=--gR6X-ONaRA0=)a9<6gL
G;2]g.\\NDRW@0]+W\.FS[cV-R;cJI]fL]VJ[<6]cdK:[<E@?NfaHB?_(aXHG=,9
>F,JIQZ+e&bH]ZSPN4MW\3FMMOO1K[U]KI_a,ae?0HeVW3V8AUND&-MKR/A0JXH2
E.=,-[^FDK:0eQ,W^OX#cAR_]_McEfF3^.PF0SRcVc4a:JMNAC(R0c8:&F^;a040
YI3P7M?;IXPY5Y4FOg)F#?W=_0?VUB.cQ;/B)J(R^0aHEG<cT8_]#KJYVDgRY:.S
=2g3PNb=f;5XYD2Y[Qa.&3KC\[/^6a>5dK;)?5H@_\fff4ed3SA<d;IJ,Q)Z>-0X
#+SH^dD^aEH27=W3(7V^O#))3RV=@W&Pe?a&^MMe,8JbPKD&+.9=(_NL/8-XU2-G
(#Y<3#SL3J]?R(EHa0HJUSN^1b#1.<2X>>FS6.\I;&=US41JgG]&SY^Oe,W;N\b<
NO-KFN0FZUFSHdN877JM:1Kc,_VfcQ-T45F5F..5@UeZ7N4^T(\XD>8f4429[Oe#
\-ABNc3(R8DS3:e#/aD2<3;@]eI<38A<7F?M6M7PS)IV6HbW6<@a8JILIFg@V>9O
,bg_3H#;Pf=bNb_f02KR[>=#Y(fO<T5a4[SMCZ.#Z.>3VW[6-XD&SJ3&-E>Fa\@<
4R)MZ)a?6/W(ZN6D8+G-+531BNf3edaF\JEBf)G^PgO6G?7K8J=CWc&7=80DeDF;
Z-QRS2-+7/_Z41?f;H-UN^83>9Y[TP_5-T=b]b^&]e1g_O,P;,<bbd/Jg>0C+d+5
6@4\PL,E>:MDJ9/3?76L772<FO^;W?#B\6]QW<-IB+/?I#V-ZT2=<N8[&F2Y_37^
.9G8<+Y&1E4E6V&\.4I5&f<\:FVSCLFCGXdMX]E/b_Q@^N7HUK(a_F@aaXM#]3N\
dP@Z_LZZa1_A#d^U265Q.I:OP:aeQ8DFQe@JRB0P@4_@MEXC4Q+b0ERRYOF+?-a,
OIQE<4^9LDfPL07&V\7W=L.OT_/BI7.g+T6dX66#I6NXEbBI@]M_P#b;VG<H+]_4
?#1ERKYHe.?.f/ROOOS6VZ(@_54V/IK6>b+][(1WYRCIb=c=HVI5G<]_,WZDC2Hf
IX1eBA8fKI3CK,PU?U&Q3U5;E^TX&54gSH9K6eG&EPOIDR\-7:S^T78bF&<BV[@[
.aJ51)P#QO)5V,T_97#SbI2[eHOWb-YeQ8DK1K(a4#.:6N+9-6+P&.;6_QREE4#/
,Sb3<54Q@B@\N6LdM>^EC[g1GI#21UESHWG,7C6UGgXRT+=@QP\3XOM^@3A,YF;/
7R=EW8T-ZT@>VJ[+W>6DEM#+Kcc[Y5NVP-@Gb@5YMNC/MEB)9#IBR<[dBb6S./C1
=2SQ9Y+,J8JM+]PTdV#Y\Ue_J<-G=^+E4\AQcdY\K8B6V]GWOXUD@L6ABW24K:BT
P[GM6d7F3X_VRM6HD.&0N]+U1RcIV1=d-YH5&.^UY\C2?=8AEK/R=d^@HAG),G80
)BBZ8/OS4e/:J;^#f4]S=(0MA=2DDe-:-ONFbZO\.-OJR1fe.cL79cC<G?eQ@A&0
g8-S#gIe2a:_,D#bZB)G@bc6?H>/WE:+c2W4bf1c^Y><d5SA-?+KN5(#/>4FX\Ld
T8G18CcNT04gTa+@Y&]^SZP?0P+J_9e)\_N:f.:?dc:E3e5H37e_eTMbBf+b3?Z:
&<9fZ.OT8NM;(Vbg]f_d+,7\].HT=eM9DUBYRS4=6Y8UfFU<2?F,<:.+07>NOMVJ
gCXY#)7VY0.<4J,RW+3#;a]2H7A4Qg:TOW7c?;)-^N2-IXW@<d:0Y0B@;^>R+&dT
A/f.QfL1A;5;AXX0IORBVc?6@aHAOg6.HYJ#6aCFdNBQ4U/>Leg]bbE\#V952NAe
,Y)?23b4WgT^MBeBW5V336@[Q:E)MdU51IRMZG<>BDbO+RZeTWEJfRQd.;C]0Q^I
38V(QMT>R>.8bI0O1\(+cVN,>c@gS[Y2S4VR_cHU];]]UO<WLW\<cDaF@bN<MX;=
;E,E7)GM(>1-#&[3dXcb^/<O#/6RIAa_77-VSRKc1AABf>_2a@]W=5#,#5d\68e+
GKNLbLWd),V)>FPVVH;XFaP(:OWNAA/gfXa=X&g05R5=?QgP5f:,[3^<T#B4#1H8
,]#.3N@M5HP;M1S+BJQRYQ+WO<#dJf6XDGfZT[\>QVG\_LB:PF.D8#MH]=fAGb=6
[MJM()1FOg4T&]-.&]DM[Oa2dF&UbXPEYP:L0;<;H(VV#XPVC:b5[,[F,2<,9gMD
1f4(G4H7Zcf6dZ6&&b_>#c]BGHUb2\aX]6Ge1TeY0AeAZ,W6I_S0;/[A:LJ:<(H7
G#;b17BB<_PbQ0PaAbb\4KdER<S(YNE68PH+Y.MJ9RfJ^Qc/JRC_79H0e+TN\.D4
\9L@1d5X+>EdD>#DM7EgJdA/EFRG,1W@F(-J=X_99]I<aagG-UFR0XLOHV0Q/.[&
W(S8.d^,]JO<;62=QEFRNZ@<d52O(bBc@VQc]NR^Z</5gL1YC;=/J=Z/DL.6c[/1
#bA9g+[+dR0)KCJQ#1MY8-40a@9]I45Yb<K4EF(S+/@1AV/ARMYX_DI&(0V+P,29
DgGDF->DN[6XXf5WWZ:5]Q5bCXUZ27>T9XT8H/C)Jg)[7]&Og2I#6PM6[WZF59G(
bLa:5=MOGCbKa7)1AYOT;0V(/#ec4J:^X^(2L7K&D<RG=02#(B4@Pg@CU1+BDTOQ
T5EPQ+D+(>@C@\Y[cIP/ZVBTeaAAe3KZ?:?#]PYCK57cX&H_OaIS2EE5/<eM_(@&
FA=Q-8&#.&T\9R,gPK1CWL>2L=CCS/PNaRgf_EH<X]b;RfHQB9^e8Oa1T>d#1cAd
A)2W6acN>\c:RKYN??-B-MNU:N3=bP>#f?M45C<OFLVNLM4T+Y;N,=f+^CDVD/ge
UALEIR?3g&P[)F<#BSU?D9(#Q-g^((6N#YN(O4H8:3E^IL()=6f5]S<dJY]O7<N=
Dg,A)@:d:>-,+WeM+dS2]&34+YdcN\QB0<KB5.(]D-W?_Y8EGO]A#6df\2+3gM+]
20@[2U,0L/c7&Fe,[WB&)][LYDZe,1C80=)=.Z^G/T>dB&^Af\=c&Zd54[HC@@-?
W=JfI86Tf0(GLIX5S<Tb:Z/+LF13(<dT\COZWU&)(:eZ8U_^]EObBRY9U+cY7E(U
(NgB]<9.+PR_60K+=cHO/MFNCEX\LBFV+ObUXSb;K3+K0027V)]3UAf_Td]bUe1O
0#R#e3;^bDTR_7,Me8Y/0F7R_/YTU/U0OgH3M_;^fMc;I6_-&><DVEU7)5+Q)O^O
,:9D)=d]H(KL:T=\Y88UPf[B>DS_(5Hc<;LN\JU\B5\Va\g1W1R4CW3Z^ELA#<P?
0VdE^EA?VT&W53#.35BA_N8;A8?HL@0](;:gfOf[d#LH5#b.PfgY]JTIV2DT2<Te
J->^5.gJ\R2?Ge[):JN.M2H_])]Z<LX8MFURG-04=(Z8436[:gbb4,X]?^QVdG^X
.1F#:cX9@fWK?-DRda;P/O>^O8NMEF:^+)e<XUa<JbbDJUR1TEGcW&3FIbBJBGVX
\QYL\[>?N+)MD1417L\S2UF/KZ0cF+-;DS4N6baY+D=X0&d=ZQ7#VaYF&C6ReA>\
WeGZfVFQT#)B/@5LP12\0fICD414T?Qa7/[MTL27SE:@HER0eaGXR<aFD[[2;G3<
=F,UXg^/a7[<4EA1F]VV\4T_A0628B;@]8YJ?S2G=D:N9:DbA^:g_@@:fVI@E39d
X[bAd,X/IT0Z\U^aPd<>[fLCYNKa:JJNU3/V/[4UHbO7IXV^NJ68OdbWE^4&JFI0
3C<N:V:)\a_d.,8dA:WgdLW^Z?YEe?V)I;6?cd86W^#&<eIX_E<1U#G7;J97G<ZH
59.Z,g0STf5cFeUSOTXF2Ee=.Z/fPHA,&<]E)M9X8,EG)/YB?9#H14OUdZG[]5c,
0BfgEV0DU;L3AbeT6-0?d)?055<YN@=,26B5@HeE[&Kc./NO(&g.7ZC5L.K.)/7=
=L(;=ZJ]XH>.:4[VMTULc<X/b?^Q5d&#RP3b+=P:@&F7CBa\[aA_3P_.)32QgN/8
_e>\6:a\/HgV29?>IcaF&QP>9D^cJ/994#@QI-I-AQO514+K5Ee=f5M9EB[6[eEX
/:6,_F<f#M]-^QK_&.LMI(g>=[1fYQ.)Z=VYEQ3<,66C]JeQ[V;ab/MF4a;6fMKF
HEg)CO>I4J>e1^YE.6)[F5aQQ:V)3+VH2b)[D.<g[Xdc(#)[S=1ZC/>R^eU.3.DD
^c-OJ\Hbdc.97M-HPZ@>1E&D=S&Q_dN)62_:D:F6eCc2OVLSY:C#0#9:bPI:5=3-
H0E2N5FR(&:+OD7V2X30TU7aB[?&Cg/E8XI=Le5-9cA[W>a3Ja7#C^&(>RR3)-VD
#B,gKPWgaW3@[U&^<X,A32CG_DW,<Z--0C6;;H4S4Pg8Q.R.aX891.YA-__A-,-V
:XY5(X3?Uf_5gO(S/(_SZ?OMg>PY]C5+P9H7[P_Q1.+c:.XO_GSgQ;HU4+>1.d97
&5JeE@+PW0G2.JO^UQR(MU=J29+>UO6YX?9ba-.:a21UQ1;adJ?@L+CX<(1^:##[
/.\Z:J-TcO],<=Z047?06YB3bBD6U#RaHf8.).?01CGBeU4YJ=3BCB[U<gJ20\S(
.1.XWIZP<[9E^C3-C?:+Mf6gAJ^BUA8,L6#aK?WS<7V)#(cT//KS1[P+gFG7^(cS
Cbf2f>7UOGZHU8OM9@]Bd[^M/6/YN7<\d\6A<^M-TYA(8-(I8aK)RM5F0_(]e4C=
^B,,C6]>g0AQJ^N^VGeb8+8fB2?8Lg;QSKA?Y\JgZ]1N(#-\<g/d-U>8.S59?/A#
H#&d0&++XF@7FY+_WL-R^?_>&,5ZK8&Q3eQA^e#58.>QKMQ[<Qg06)56X+.WEHX,
F,D0:^S8U7\@RgU4)a=d0)G,1I36^XM.-@e(=Sc.N)CeUgK0X:geU]RSN>13(+-6
/f^JTGLMUULI>]<8d72c/NLB\\.3&Y\_/XR=^]X,SI6PY1Jc)b\aTBYaMD)c12;4
C=18+V,\U4<H99X9&d>9S#?\^ICV#?_NU/@(dTB<eAE]SE4f+eAA]=?EH_@X-[]2
()V1#(;YFD&@5P;bJ5RA=+H/J^4?d3O[<Z2EIGW=]XJSN>EGa@>E=,-Z6d^VB4F+
MXYL_Y\IBIX07<Q9=8P6)?aBFNCZEV5>5BQR41MJRSb,CP6,fD#KYP1If453O=A,
N)RgJ/<\YC3+gZSD>I3#DD-=]^.L[#d(/T#16+9YV=Nb,6.P&eg,)PVc,b1^S#-g
<\Z;&\_;X?aXd39Mg>R6H41MbW:0McfI^1Od&Vf\UHB+DeP;=gN_=HT6@dV^3@0?
O1/<)-0;cBTJRUE6I0cfeHg.\6f\8R,eE\J?fb21-YG:-)T#.WVSPT,f@S]Z^75R
,FWH?4>19I42CN6P0S<Z,6],9cfe1X27K>XKS^/+eLb,7Z_^7aL/OI@N/H+WIM]4
5&6:)(_#dfFWRU:QYKf&0BEa.F]e#EKIOD6P&MZGJB8[6I_RRGgNM9(6gW+KI(\J
&#:LBHQB>&CVV-<gG=J#9#/YANI:R;ICGOQN;f>a7A@CZLKG/WH_>gQDS.&&(8a;
ZE)QT>17^6ATHB>35<40]\MSSPNUXJPa,,1PdY;Q3M6O14>)5]g;LMSRC-Z<>.U=
O9F]JKKV.B=?a1Qc[&EXD6-GZP&[_2Q[5e>eC&X/P0:eP#DH5@?N(_bF@L(BcCcD
_?7?RPdC^.Gacb)8&[C>E\c[:EeM.?U>b/?XM9_6,CX:M62W>ZL=CdHK6Z813BTc
a0MUO9VWBW5+_\E_N=<gNgR?>&eW#+]@Z<)<I(b9W=KA8cQN2J@U#(XTUKJE<:;;
,\F(9F8Ee8II;f83?9>WEREa#FAVN642,+Q.e2U?VWGFVE\.B8MfD.&Y7GLP\/g_
GZ]1bM,&?)(L4(+^Pc>OeHT^+:f?X#a\C#MdO3@3,G0([RQN7:If_[&1&6-,[Ef1
7CK=Ha#K+;1b5cW&<)He<bKU\#Df2\BEdT03I_T2C-<-eDT]G-S^VN>B4].b];U<
)5WM.@HXAT#2;Vg:]LV;V[^I,<5T6=]-b9<Q\_4N27=QR,)L9QNZ8OdA8WV.;(cV
0O\D2KW#N5?K8g5S35VMON8^H>NTFTAD62/,-fKc_e=;#@HCT2EU>\bb,PBK<;8J
:7f4J8eCU8eDZ1_2fYOOUYQg1642[R6=_[&eDV[,CH<VOEacAPCT0H#.HI(7>#RV
&JfDR@NP66M]].:MOPPJ1&3T.eeEM0=))>[&^#)/&4Ng]RG-@=]]=-bWHKAW>Q+\
NgQ7/2@)XF<HN<2S=</\BWB=<YZ)I\dKCUQPR6-Q[?K9<,:M]=:X:CUO0DK6=Z76
<>,:(Z?X)DF_.R^@VWVWQ\]2T.OA9,G4T)T&3ecge1QAJ7BA^RFZaZ^&D/AMR]2+
NIdKdc7D5@1c^2N#ZZc3N(-^HQb8fOL[?-U8cZ4&64WUES,78bdNLe6W.c&L/.DQ
8eSOa/W6V.Ja&K4-R#WDTPQ#dB_P2510(B^J65F2G.23@^aWGFU7Z+bF3G1,+]D;
[(1#;[;Q=O_<CNRWB/=#eUe-b4BRHb9dZJY&+N]=X5S,b:\P-NH3XVB43PA@/XJ[
9#<@)UEI]K>C7M1e\-SZA(c][I+>-B4953gO)C1Rc[U8RSaV4>Af2&f(4Z7?O]V7
AfG(MNb4JS-aS&BD9#fTe/,M+_d90fM[&)C#U-J_c,[G7&FJ)8D8F1)1SB>I)d=W
6_Z35]@bWF2?D+LM=@743#9_@\[_+)C&bd>8.GPEUX.HRFY@IWF3-T5U0Ca&5404
,-BP-If15O#U(&\C7Le\UJ<,=SX.EQWL8fB/aVTPIIW.(J794;g=Z00f\O99UWV4
0G\KH_&F\[4IN+GGTYU<:Y,b#2UZUaZ?+T-=.6&a^E=Q2I6Qd8D7J7B17M^4:?Y/
Kc\bK_d;UBSNCFRKaZ@<YbX:dHM&F6e7=1Q=<_^2LQEFP20F/6&\2Oc3d4a3Ig0]
gH,:H)URXC\e6)=E9,Sc47NRF-e^4R_bd#2-Ag).P9NC6/N0,EeJa1@SQ)<[,EXc
aB1+GQ^;N/OR6;Q:O+-H9\-J->&S5gXRa>d247fU?8+g8N7>U)?G<EE@7e8:[HO9
R<4=d0-d</M.58=[;K0]faa2cJ-TMg4KN[WW1:1Q5P7+(+NYDe<.]:2.B<:c,AO]
#BFH.?3>CUSa[O5.YVG6&<TNY8R(gS\8/H8IBKV6LK_1WL@3RV?^4=(V0Xd50K:B
6XC79f-##I&SUb>OZL[aBTS2P5NUNa=2P;3BgOba0Kgd6^N1,M:M>6Y;><V1@#9?
Ig=#MD&fP,?M+MQ37=7E1,Jd\Dc]W0:JJ[AL0f\N3XFa[<^XB&b\K8/8+RC]J::&
E1_[A[DH-,9E?33@6XJ,a53bEEK6N7A6d]5Re3cZMa\OEMT]#bTZ1#FL8U?]);fF
ae[SU-f;fB#,4#?M#L@-gU)/0N(4.]U(8,W<71@P+=P\Vb+WV6@&ZECI5L_[LF9Y
;&9gOT4@_WY;[LE(e8.93U&>D(5.;;T3IQ[Q[]6SVY2@C_)4NF>Z)+EFcL+R/f7R
0edSa(;IJeNE4FS\(UdA5E]K:g8&)_d&O2L0C3;=S,;8dd6d;_LOS@X<EMMFW+JO
@CW/UJaR?ZGQVfIH0I<@.58e>HXY8,PIeS(4,8(AR9Nc;(d9N)=b.:(F6bOUS-C<
I:C5AFaMd>LAd5gB;QTN_c=/:NTe7MBQ67+3-Yc[\@)U8If,H]V/efBI+)_@7F1H
>PE-GJO1&H&(OfF<OE?2#EG(#4\H;_Od3YOcUeH6I<7dX?MU:6CaaL/QXNK5KKZE
=L?1ZB@8TLd)49^.Q<</E:DF8B(MbR:\)56OcZ+Qd4_S-D.+U@&NaK&f3N)[UHK^
6.-XBHJg-2DLdX/X(XS(D_;A&;?>7_c\^F;8_1]<BN&9@,a:J<+HbeW_G@BHO\.I
78@?@&Z_2#7#[C7=>Y\/GKK7feKK8<^Dcf9^AcS0DcQ++0aIK>M(C_I+HEaC=QN7
[\MBAM,)>I\18SAFC_/:F9YQ0/PL;X59;6e>__M(2Ha6&0;beU?OPI#^@A\B:IUS
#N(5G>IT5V.6M:53e03H.>cSD<C=L,-dd#\&3;YR^#cPGE_10@Q#=X727aT[&FbV
;VcG5#?dfA/[+fd(,<XZ>04RZ[1[a),C<B?__93>.&@AR)1OSN8g&<JU[-BRB393
JV<R?Vd=M-1]ZNHcPFe83QLNQR8QgZHLBK^A=W#.TF]Bfg28,b(GEMHI#T7&CU(4
;c3_a05F1E]UQL.ZM<]I/?.QKaS;9beWW1@8X:;,\WaD9^UP1TNKKUVQPb^d4B##
0;)1A+BA3[_[Vd],bITNc@bdL,fC+4ED+?N9\JM,5U+dGJ@:=GXSW.aK<9KJ/a(Q
H)d:Hbe^d>XL^2D_5#U.]=EeVRQTXfQ/,=4bS1CdA4J^/C3>F65)[dQD?OZea[cD
bVX,,7#c6f8;@3c5L/_.]B9EDS2E>^IROTO?aU01]F4LF9H(>&V,_2MJ#P+_U9(<
WW&0UZ_(\6F1BH+:F\7\gbd6]^?COU(I\I5)YQ(]S)2TgYB55+N#D9C6&^.d#_(U
6BFcSPI@QHFJR6]bM-eGB5=)cTHF3<P-)?VMWQ2B@KBKFMDQ_FXHVN4dXIP(=F&M
7O#(\?+A,c\RID70WVdI(_^2S_(J+LM+C^5AMM&f:1IC[&W\M;N-,9G_9Sf:Z3Wb
EU&#&/98PNO_YO1N:S;)Z@Z./X?&e;U511,5):2^4ga4F^##bdg?\T15O2&Q3V<g
^Rb]BMW2GXS7dM2g4UWM+fO_IIYD85;ERO\Ca9:&TKN:(b&I^aa/&#M(&/@@W/20
..^C2Gd+V@7-H;G-(B.ccFD/]A#SBc?&8.R0./)G7+F9f\YWaG[38a:>JW(_O]+;
R:D_.F8R#[-Y,U.KRNJVPOW#5/(:.2;YUceF=gYb^Q(C()R/&gg_<3037[2?_d12
.:/]MYbE;Yed4>gfKW\f+KC-bV@76=,QbEa#S=U+>=NU?UVN0KCOVH+FU#+NMLad
Ie-=?7DY^[5f+&bBEZX,ZdPeI3^;5K6AYQ/(da6T-FCDKO#fGT9e:-b2SfS+0^:c
fMZ0HR10MBY3X<NZ_]X,BfMO5ba24?;2&=&:2Y^OE7c3:3[b)X6PRNQ.Z=7O1<P,
;K:2]&CV(UcYA_=X@4?a@]=N^Y(U#4c,6G^LL_^I3-0=DOJaFG#Q<:##bW]4+[_a
@\a/V/(:.K,G>-P3GX5(K7,b7=><V[G=L3<=JY<E;EBX#VD\IK&OO6FO&Pa0QZSY
K,R1R:HZRbI4HZfR.J\VA@\KPB5]U1:YEf=5gK(b/A?NC>e#1&Uccb\LTgC7R,DP
W04<7&b^5F0eZKE_\+O=_VH2)OVIae78)>-F@MKg-<T[D>LRJT;REg?DMXVSHZb]
U4](EW7(;Eg3RW9F6LL,OFEfE)_-KbPLPdL=U2>ZOOS+=3SU0-&Lg@Q-ac(Z9A[B
1gVJU9b-gR5=bLV\cQ&ddPfc(?bV/#@QED:T8K0EB_E<eKI9eg]?aVg]#Z:?#H_+
LfI:1?GNR[QP&.O_F:JVbLZ^<O&JU]dE6>R[FA&cQGLId]TD-SA;=BeB:dE,[aId
R6fK5G-@UAe^I?G4e@M2H)39d0#Z?<2QPfZN5#\4&#(0Z\G,<-21=bDY.9Z7G0NO
LY&I\dS-6bE;[DDD<3\-+=S.2T>A](LU)e(>E^Z8:GBAXS/;L.6A,>LB+=Ib93-g
NMeKbN74:1MH3f4]A7)Q].LEKaWP8>6>Y(RWbW>,7<QVL^faPE@#DDTbb80e<eOH
HcF7Ua>f;3WNR,+JF&+_-WGF()=([K4,QGS09@=0#.b3C8H@KRJ:NdP==0;HgWfR
-D]G1=57+2L;3^)J.9818D=))SNQgDIS1@98TEbO+gUM7C5/_PJG6O)<S6U#P:e<
[NTJPO(bMY3DH3V&[BBY)R0=.J,/#_f#cL4-HUIZZaRPJ+_\bfG-P63H=P(ZYg)-
(#=B&)KI]CbgV>Hf@Z\<D&b1/fOC+3<?IY5SK[Ic1Hf<#K=MY)T94?.&HKgU(5V>
?9\N&1HY:.:+^871:Z.Qc03X5T4LVN,K,/)+11519D?Y:cY@<?6>?eKDY1S_c8YP
e6:;<1Af;T(FD3d@WI,:[=.;=/5AEK]Z,LbY#-_SA2gg([a+^We5&&0@aTceeWNT
R69LN&1N-I@5eNaFeK39B0/LX\dW/H4,K]PJH1-1b1(9G)7bf^gA5O).:Y)aO^3@
C;UGVH\/[/G2DfOaK:N/L.3_U2W/TJ?;M9b3B.E6\WMO:34J^8WH:[Nec.=P]VQK
QP2HMZ7L<6a#<P,]a_9R?9;USZA&gNPHOW5R,@Cg[eQg<J5=/938=+8d#URQB6?U
X\Ae+IWF7<8MA:\;>;9CE1)B(X^4\\KSJF/<47_T8@#Q1)FK-6\Fb@>VO_7(g?8:
^c6+M^<_?_)U+,,/;4/GU@#:]<+HI3a?/TZW2^LXYYMCX_MKB^,\f_aP5+8WA@;=
MaBM[e17,g0dPTE\,MZ0B_bBK?R.?0\Z_MAF:5E66]V3[5(^E,1]9H1gG9P5]e=^
P>Q:;7b_U,>SEfI&(aD3:-5agQ&O6WIe]M=X\agMDH2H\C:[,K(2?O@A/YORdJ&#
g\G)+;VZV?,8AWT0;;c?UX>C&?.QdYQTNYMb.RO0F5.TO>7@-.L;;,SN-(8MK]Z@
&3LDVUEPf4FCc6U+RJ4)CW_.;LF?GYa0K8]/MbY[d<^Ea6X[PVN>K)@62&6]/e&=
(#eB=<:,#Ig/#d(EFcX_7THQ(I>Z?U<EE;K4N/OZC-g0eX>)a\LH;B;>4<A^6-TY
.V\gXbG9gMMX5.D(Y/Q52^1a@UP[<QIf;a0WHT?,[eSb<./B(f0[2L4QecMYT6H5
edecIK)cb.(AS4Cc/S#d1H>?a</V9JK]J2/BI_TM6RNE[HRHa\0)@7_(?QfO7F=3
c@G.]TaB>;BVa);)2eD,^[HdE\1JD)&^a>U[IL>^M2]J5X+Q=:7TbD9]4b]=KNTW
H)3MPOOIdJ(^c0X>B_c2=:D09]b@aTDL4XNeg]XT<b:;^-[E/2_31F3>Xd1]VRO+
G@[^91aC38?3GOMJ&4YIJY+8C>#+40UQDAF2-S>\N#,eZQ\8&?Tg9=BGMYR74XDD
,67+,O-^+A[fa0XPgbQK[96)2E5;@aEP.c:Ub;EC@=07TbVB]^BPZK/d//,\,DYV
(f0e76;f,#)I3.R<K<E.aC)3E<.Y0F95L&6>U&f4J<995;SX6Y:6>cMVN^06FbDV
IEI2Q0[c71G6&(=:b;M<&+7OU.]gY=d.KZAgaTK]T,0^[:Q>fU9NAA@^AfWC;\8D
gb8gQ\AWX2;HX;;ZNZa2#QdS^<-ZV0]GaX1eFD2dXV,O4XGV;?I;6(6R1gER0?#e
_8BW=DY4S0eC<#eG7C@cYL6fdWfNOL0gFGV4#>R<Xgf1f)(LE9.HLVO=98]fM5T/
BId1??D,UY?@+VY52Ze74N=7&V\MQ^[W9246[gM^A:)[e(,Z+];Q0[^e(MKIS/f_
:^MMSP\/cD-H,:YD>6;J2;3g<M,)FaNKK=]WHA]V/VZWMU<#ad@2cWH]H7bC)H[7
?R/T<YU:V.59>;AP,g)_/:O>UJZ^JWNY72GdaJ+HYE7-Za7HJY57WH,,RULc+c.R
P4JAUE=,c=AW4\gV4:DU1VfGK<X75QH04[E)V(8=6,^MWG3Q>78840e(a6?\G(/4
U\[2GC.I@MW5>Ca99#?)01]1.>@+[fXYe[5a:=^dWC,<41>5.W>Nc:=6=(,2IRW^
]1UPYLa@^K^#(;541D?\>bWf5QD,bgaEU?-Q-d+]U,#XQa#RAdgKG<ZS#?U(H6U>
4]QaZ.0P)dVU:YFI.UeV&9/e>?_.R9N\N;/LgAFNfGSAJ/MN5(:LCK&ZS/a+AF1#
gXE>a#]H,9O6_#T\NU1^B>1\S.T=c<>Y4O(EdOdRSEXM>K088G[#aPH3TJ2+OJ(\
Nc+WP2CLP_N],PY\?NBg,MYUV/I2H38--F><:6=L&E/9_B5=WX5I4I6-b-O)0YLf
egZ@g?J&./F9eeV7AM<3OO8]F_XZ5ad^PT]gHNPOd>[_A>PVHgETP0@/Gb<W/6;;
G[Kd,K/2_<B9#_QMfGUC+#d6]U:^EGZR_M+_^+Ve^8\=MJ^?TWXF9S[CRDfbE:aY
M2d,MG]7RH@\W7)9EA18;3/9NMEE@(#&36X)RTbPW,?TUX<TG4aT_>7KASNW\HUI
;:9KR&0bS?VXBG#,bb70\\JFcEN^Db6&G5<0VJLL.D2)9Be8L2Ob@:+SH8B&[[KD
,HA?GI0aZ8)YEaV]GAVVF7<P.A;66B^E.J)UZO@+FK8ZD\1I<\=U/Sf&K&c-(aDG
cI@bL8_^WMHfTCTD.gV2NUY0E6]2F;8S+0P&.)c.e4eZDDU2;^S+53YVO^K;g=RR
M=X-M1CSJ3c6)5J+AR@YL[)g+RF7A_#=+;ZNN2bU7\JBGOeU\@EBW7P)X\_TbCG1
;?[R>)-XK>dXMDbb3&<44L#d/?S)2bY)Rg1&G)[GR6XeV):W3)I:&f=4RGW);HfO
=[H09G)MgU8R2H,e-]dcEQfJ&S_6:69g^BN)GE[^YKefG2&R=FEedE^I)aT+@9)B
AAdc8;)+dF1+SYMg[W;^I[U+eZ^1d1VS>cJ?BaF1?5dX-A=5+&L1LJUE1I]d\1TU
IeCU?>>E8.?&8XdH:200+ef)7G^QI@Y]J+4<<PeQaGT]2f\cJJMA)RN(]+K[EGHS
?II5aJ1aeNQ#(eVgI24O_G2P_<0[T:^&0FASTdSaIg.LDN29GLTSZGgfI<S6cgD=
B3Q1daeKS2UI&K33K4/Z&>^S=#+])JKB]A5JXL6.=VINY>AUT<bPb2V8eagR19Nc
TU=R4&,5YeRDa/=K_1R7_W@Z=d(\.fYZ^Ia\0I&eaK-#1ec1[^]6+BKW5)B&U4^9
RQJ./7^B@NGQDP#_8_dHdJbX2bT(5(4QbUfCTDKbdEVgL;4d_UBbBR&]>X;JE<B\
&L4dcaI:cTV2E:>,gD]UWa#J:3A.-fOV<;OReEeZ:YUI,X+/eCbHF+#]<A/SO^gd
.#_?Ae]>.@OBAW9/g;]7=R;bR7a-.;(eH,1>PXfa(c[2f]O:_d3/V<W\YST4L(5R
U,DU?c)RY4+0WN?6OOR/=Cg-FdUVe:8+JTP)E/)EV)\L3gW:fUM]9A/Dd8NTR1XK
-0U\YC)U@:X:Ma)bYN9LP_MMYNFHbLX,Ee[[f=CB-\,?b2Z3:Sa--G]N]e3&E/A>
W5C(0Y_/Ref0-Ad4K0CWP<YOGB@PA1E;+F@L]>F3LKcS#&aWZHTdI:@:G(beO\aK
7,Kbg8gC+JOE-d,&UCEU6e</T5[=&#]YPUafS<0F_FU4<ZXPYa];F#(+[7U6OU)3
9J7XUB9PF+JS?,3@LZIR-+H<(M][;LO+-SEB,^f5c<\4>ICK7^fEP\;-W[QQTOY#
LV\EA0V9LB?F6X?]bUA8aM<W1+EO0>L+;.ON[PJPRV\bFZ9Fg<_#>JK_f>\OF/LW
D3UKgT)7;,M=N?e2Q_1UZ,F?D^/K<KY:Z6YR_:5&^VF0(S=Uf&;PM@/P#dA]]69?
L:>26A^((8K^=;TRSRFD>eD-#&IMIH:A)c-R.4NZ1ST0Q-V\DJd6@:K-^eO_4b.8
3c>BT>XL3\>,ZP5)9/ACT[)6OBN0(#7KU<2-R+a-dL(QBB1L1c3cBJ5K:617eAJf
c3G0-)BU?RR.;[@D3_cSVcD@7KHAV/Ua61DBEa;+X\2]KYMZ/P,D?.YH#.OM-L_V
5R67BWOgQ_C;W.>;:Mbb&D@E/^cH_:XGHa58J?4#c8,>1?_Z)>gQ@:G.>CR:I7O3
6bZ,b373,-+\:L?WQLdgf+8a],D(?[,YV#d6SO36UR5Bb28Z#@Q)?:#:J<6_IOA\
dW0CRJd6(2;\.@<U6W_HW2+&#fT>3e5\eG[]aadD6]FH,;O@N2(JAV:U1:GdIeXK
\I+Yd^7[?3ZV(2Q-J:1fe8Z(.6+&?WJ2Yd:R>aTeLNeQbVB)RQ^_Q;7MRQ8&J5f>
BM/S_-+Kc[1Z^IK(e]7V-^?WZ9)&9Eab[^]FMR0.A2\aSOH^ddbZ-H#2cT-_JTYP
66];<O8WQcI^UJ4UcL<HV/<:)X]aH]>?O&6L;7H\2E:6U-=aMAPH=;ZRfAHX#,B9
-]ZcS.#73>BTTd(]&@-@ZWPQ9@6\A9J)4GPHGe6K,).U8W+/37]]CHR4[fONRB4,
_GP34SE52Q8K>MeF_\^7F;I>,;>Y6N=;K:c6fEHYCE/OWM:)>,8KPc2KP=WH\c4A
aAKfAE@W[SbRG]GNLIL5T,d.\)2)d;L+XDC@\+2>;H])\FaD/_022:Z]\RY7\MR5
K\+J6JDaJ[3CY9ec9?DP-3W-fORJEOT4R_4cfe#<+?Zf->/H=FY2R\1&cX:J==L2
Z[.MK?<F5dcI)WaFAF-Q,dREZZEWG9:_8<MGd)+FQ_:20ZIKe&X8d>18,UK:/N;E
eRYNB>a+[G-5@A]C8-L+4d#\+P=,c;0ZH11;E4O5DG(f&(3YDJ.TPUG8JEXTCT]I
A:G;@f@)]Q2VU+_F&e:LcD-eS0R<5-S4\)NZcJKYI:.]4Q15@OZ=Q\L,-.F5#F:#
dNFN23IOb2/J0D07J-Y[++2@VZZZ,4=>>2d(SHWAN]gK285B0@,g97E7c-RWf]3a
+/:,0<(6\T:H/8Ee;ZHCc\@W7c(8PWA0R=EENF0MDK,H554&Ua6,Jg&c;NB>^O;S
N6)ZUg(FQKQ#+MO>29CbGB8TV9:\_]2?QJLI[/I8_?fW&-_19\EX5;8<](;WR]+c
dQEdLC>Q(=.ALJd-GJ08d[IOGIS+aM<NeP)1+YTQ3Q9)+g0C]LeEESYX);.T+Se\
?E@dGKA^(cF<RbNT:-,?IUDOS8dX]&;cJJK0>1SNOO36[2160ZY;XTH2/YZ@6Q&9
B=#U_c(W2&=c?VNQ\>D1:Cc90S63IVU:46[.69_>EN2d.N\J-\YE\N1-PP>,OFKd
JH+V<,<0:FO:e=SV2++THI1GUVOP]L9^:>0N6NJK7U.Pd,3-Y(Rb)R:_2a7&P0#d
1&dY:?7b[KM>ORbVA5KH/B@c.#cNU([3gY7D,M:Fc]>f3)SU.D=?,R@GJI-1d\6S
7:_O-4T^-7MLL0>f4[5?0CXKGbS,[#B5Z5@F82]g+TaKfffKeWN,[F2f<g=FKdf6
Q@;F\^;/.?eSgMR8Y1f9MUDbHEVWF\^6YgDXT\L<Z6J^[U))FR(OP,b>gf#YOF,d
>_HP2XR2/H.OFN?J7I_JX+O+R.B9[AQ_7SVb&AMX]EUHL?:3PCV,DD?X#KO#0PH-
9Le_WONU/)A<L18DFcQ3VJ=;,E/dMQd^15f2P6W1)P^a^9U1d:E3RZdCe52B7>1X
0P+[<N>&L5Q>OC]d0,SB/g<:b^I7K>[E;3?PRP.3GfPZM8X.N]f-4OdAfS&C.L#^
W2)OJ;6e.1X?If<SKP4G3RJ@U:Jb&8V,O,@EXR^-8-fEZ)b-(=RTN39KCQY;TPH]
U_9FN_&gT8Jb^gRW+&OM)I0BeI:T)aI94BHXf7\cPZV.&U]@FM-X&B]#:A+/.MEK
gB+A[PFf@B2XfQ>JWKe6-eeI-(N?fC<Q;TcW5NUNgbFH?N1f:fT0/cNeY+7D#4C<
>R-8?DK/=SIX2S9aIB]H-_LA\1bG6Q:[K]MIZV&CV[BBd@VXZ]Z?,L,JKVG73[:H
_4ZMS],:9==68Mb?+<WBU_GP0L9D>\4=_cVYZ>\=1:YT2;@b_FGNH52[8=KC#f9?
<]fa-3,c\QR:O4XWA=60FX(-g/6f_1Q#WfL<:_VHcY8]^X]X.;79-.A,9P#,YGZP
#(\=G+?-/Je0=)KR110QX3FM:1LE;G8VME3EeJ&B#1[?.>d)#f^:_#;ZRN(bW:LI
D=?4cMc;P3UfUFc(\ID(Q3#-dbW,415g9)RFd2E<4/A];?&C:AOI?_EQX6f3#,aQ
72+B<6MY;&Z[g-=>:5c5J9L7+(\VP&F>=J>NRc\4-DP^a-;E;\2_F;]2WW..>GBJ
Ad+JR:<5G=IC1UV:RT?22[TSW,QJ\C-D-+6,S)G40R:IB?Z.XNcLXDTGVgacIbZ;
Y[(]4\8RbPDNIAV(eD8@FSe0^dWTdMXT[5:V.YLH;BdFX@B^R\/88Z]SQEIK\1:G
RMU&JWYT4]]<+=OCU+P4&7QRP?e_fY)MNFL&?CX>bf.3V/O&eJ82g+E[/27F@Zbg
#d93Gb/EC(/TNVBJVK;RUSW9=d,b5=[Nca<YILEEJCNR^+T_c0VbALdb0[V2c3:<
GA3\c6a1TYE:,)+LG?R:MSbd/4>XPT5Kcf_#\S8V.7JA<17_T;I1?CF+b+=E_<(T
(FfS\)_#D;bP0VHISG/0BLfYC1E0-I<]:,54IDW(B&9<ea2U_aeW)3.c;?H]ZQdK
bW@[/UU8-6f0,NRJCe=Jf3T,Db(T.@]HW:7G.>>.FMERQF9_b:cCLFZ5ADb/a&EI
6W^.TXLGT?IXX@/L0.IDH=0M+@D?Q^0-SOfYPcH:M-d[\g6,,TT0_a@O,GAMY1OM
1aI3O@4BS:D&T6ZKZHJ>/8a6CLNJ1aE=>UR^?170F1LARICA0F55LTKJ[[.4c&C?
g(4\;UST>CU_5HM=V.N(HEMBE6A_QTN>gZdc821^3>a#=Z_+2Afce]LA\+K@_VE0
c.]2;OS\\[FC(VG7ATYTPPX::A8T]0NLQG8II<(ga9-.Mde-P_ga].4-K59fH)4?
R8?H^AOWEPS5]-(QX4K<Ld##@]UK@A.[c8WV+2=E0GDL<B,ZTS./,7^3>71b)6(D
5BTK@8B:MV6LQ?D>d@^O/QRI06W?>JVJF;MN=I/PDD)PM[a;-BFL3SXe.eO440,^
DJ1C<BYgK&2aVUf(TAUd>6T)YD>a4\eCU080:g3-?PK>F\)U#DAT,,_4WQ)CV4CS
.+REPd#S8Q#<\B68bB42?A3DSW1ESM7U1#9-Se)3<9R-d<b.-86Q.NX1H15O][_e
VJ_+OR-f?(>>6E?GNT=AFHa+.(QBJ(/4I];483>8;/9U8RfN.MG8=Veg,3V_TBL5
]<M2#.?30#-(b>O&G\CWc4:Z1]aL/AP1/gY=\XY)9<?9=cd10]<C#N4WU;A&^a:^
SHZb1H-ZAYZKVB.REWS8]Q8J#F13T+S^>5gI@UWO1SB[1Z=,4YC7(/ZeCF?H6K,c
=IC@,XTR[\I380gBT1c_]g7]a7WU&0?+Ng;LHfJZ^LF.&UaW-N6(g/>_LbW2SIP+
W0g?GH1;&#Y/P3E/7PGL(f)\3:J@SO0Pf&e&5IN&I(M#[cD_V4@_(;8e8;7TL0:+
P5V/.:+P@QGJ/>\R?Ng/C[#K3LXdIaECeU^Kf3df.7IeaCJ?#Q[_)>X/F>SI.=Cc
#@9^\c))_HOLVcbB^MHQ_UI8BQKF;>KDKN:9Bf/<>YV1:N-,CAcBCR=2dd[LbM\:
2c]J=U;b&1_5Be3K/gP&;&5A9dO?<,\9#YNUPP[)7D&OJJXX1A<:JEFU-JEfbfWA
2,C-_RATa1G6^=eaQ:G&eGT3S&2UDP;0[=_.B1@fb;7#K#:/36X/2E&L71:[+_Yg
,M9+M:>SZA6G)Db#\Gg@>=)]T+C+^c]F^PE/>bH1X=RN\]EgTRfTbZP>3[2Q,<b[
OC=_DT-G6O+B?.#2dbR.V#VL4CO(.3FHL?aMN?RRI#5_#fc\&VJ-F37Q(K6bJY_<
8T\RQfA5aBfdV4BPS=@af0P2(I-aO?=?[<a[DHLFG9(.Ge:5g<PQ2;VO]^L\:JJ8
(=9+?UWA1U?@geV.G3V+>IdSCSHT(,egXT/#IP#eaP5N<=90WIOBAcbAPce/XgQf
fC=^#E?CS>DNgV+2/H/K\6UfBS201Zf=WOM<Cb1(AXKg>9IIS3W=@&=P>T;S&6=8
dD#fTg+/V>eA15O)FV4?G316S>E4:H=)=H-AdYK/)e5?I?J5c^>3TIg\B3a[f>C?
=cGS>,b9O?3Q>&[X238XT8GP03G2;?+^g\dW1f9?f<M0f89g(_FFT]B/a]c>+&T2
TKE@GUN]RIMe+g[?R]&^8#\>5fcEXWFN9LT@,-VXPZSI0V\&VIS9N3-/a7DAbFe<
#J&2R0cJef+dDgK]PVKcaFLaPIE1aT-:/<D<,IO&\MIUb<,>;A1b/]AW6,QKYg_H
Sf&KMH=Pd531^>R@6b35Ra64&g3deY<QD4fXE?)84W9(LgKWM+R#W+a[HAQ=HSXa
Rd)DTM&L&D?3=<I:^8VO4J;U85-=+b_Ia].FD01T5A?DNaH@7Ic[=MVEW>I<4OFH
T^\YWGd,^)EdQ:;A>Y#T\8[2gc6<2>#P.I=V?LNg;5ca3>0G:C3\VU_M[2YaD[O4
+ZV9IU<J.1I)\.?M=X2<_dc0?#;Y5b)-EB__/H4P).JN/<EIOR#4S1CK&e;ECG_5
(,FcGe-EZEM?PMSRAF80dK(KfY=He26#-D00&^^bWc?f&VJ[XEQ404b:O>Q.JfB\
M7&#===/5A2Z9Y]];:(WJG_Q>#_ZH8E^61/H9HFGU=,7c(,:F&eBg9W=P46FL,(P
2R73&5MZ9LI]GUg).BF-=[L)[3(T2e4D-GYNMGKXJdF\Y,=.HU9JZ_8cJ6J\\_#4
\XD-c/[2MKIY#]E875C\eT@Maa.E^.8/,-DbZ2IZ#Q(W-dNJ^^YEN0R65;5(dDd>
\(>)c66^?WBDZ:V:W9YR(e\_[=DMAPK>.7LYF[??Z^GC0KXg0)[,T)L^=8OMHX[e
WA]V1Fg3#D7R5WR<72\(/@.^TQUgTRdRaD/+.BCa&7N>4JYJWIX)BP=),ZFO:aJ7
\_?6B=.YF.fHN4+d^>CB3_g5<K;^E32B:Yd]W,WfHRf@bA^XeVOHGINR;7]JF3LR
:IaXY25QKFDW^D#e)/QM^YP\1RSGAb>bX9>YS4[S=d>/OV(Z4(A)[XUJ1Bg^^KgP
(-NY<>=c]cY9N=4I9Y7Ga+X#ScI>WCa?d[;.]X.N8D(ZJ([NIMIZ.g<B7()D06\-
N?De[5Qge3[ZH]eK/^@;g\51B3;TK;A=[XH[f;L+_:M,PF)\NO=(?9PF4DS^O[>6
>)6D6JBZ+<D,=#-Y1VC>M\&EY7Sf[H5ZT10@S&A>?#1X5fZVbAFSP[6SG&7M6NNT
DBFA?EMIY\UffWF@+>2L[GTO\ZI2R0Cb)5J&;UM#\/4JHT6-&\W2c=Z21H80MSIZ
G:KbGK5Dad&.<D?4.9VC@1<#OHNg=&ABZ@@LUKIQ<J:6Q/#d,NI<A_OEQH\GQQ^E
#;f7.JWS&#,UeQYO[.SC+(=JB^A]&D1K4Y]603G6-BSd&VSWR9<4W17S)U+59T:N
\7<5b7^1#MQ_2_H+F:)(-Qg3^Y[70QG>GTM):MTABCd]dePQ1H@X&1VeQYJ8Gg1e
d1Q_-E;Z<U][?E@1d6dOHb#^a[f)a/Mg@Kfb9E4f0AO+^M7F8^(G5/f72W;ADH1R
<I;K2HFOQPa)69_D2egQX5AYQ\/-YIeTb.O8cCL;51c;b9KI=__;cg6&E=gMcQ&\
#B[-I8(,;d8gS=[HK&,(.3<6PQ);D-?)<4)<0(/gGe\9V1.>#T<c\V-AHK?(#fME
PdH9E^::O5[P,HgLIg>CCe<B^W<=:3fPNYJ;d\MUbK>AWeH(MS4L[e;a41a,/^]&
/F-efYAF+ZXe)g#=Y&2(B6T?3S6[>OM=da/CgOX+:\=<?4G(@,B>7O,9K]aOJ6_]
_23:c:[M_K26)OYJ/eG6B2[=DbbY.=HRc>PBV?b)M26F(H]W]d5^dSac1\,],DId
(a7)H&<:K9cbZ):;<B]ed.\]-MB)bg/LS7Q:N6+T<>O?d3cR,f-b(XKEJ[YR;#LW
=-d2D&>f1Eg=O22H:II9.V=-RTeA;ND-_W^c)(KC@(NA](Fc1L,0CGAdPPZaE;SU
RJ,/:F@1:YgWOCANVeeB=]gJ0(QW)R(<\0]J&[QQaFBPe8bAb20_P:ATEKf6PXeG
8beg[/=6.TPX[cC[d:EQ+?:;>;B^<5Z#G5)SX4X,<2L;):eOFKRP)K^F[:JUe^gB
ZF6;X>779L8Q8Bf<OfETT57e?4BY&\9_Z\4CfB0O9N;.BP_9QG#9)e9DDXa86MEC
BJ6>7-YBZG29RHRf\YQTgL\Gg7#J0RQ4&@Z8A)]/T5@.)5\Q?e>>B:ZT?C.>=7Yg
g\YJ=NAH@YFE#T47bX0CANE8[^S-[3Y0ZR]F#cgH1U5+<[H&c:L[gQaQGP9ed+)&
=Y01P[67R9dD?[P((][OfTC>_6]O\Q&DHYOWI_5cb.<0ZE4@II:e+e/#a-5)6W(W
,V[^>VOLa245=WH5bUb?1.SfW@M<_bCce[+XQ2\(-=b?b;gO6UgWQF@8>&9MM;6_
:QZg).S.=.e;&d0CgK(?&]G,U1aY_MO47@8I^R1_gf6USEKK-YE#^T2.SUVT;::,
6X2P?FbeM_:^c,+P1?\OI#(PT^^YYTDN;@>JEVMH5H:B,>AL0<S#6USLSY/I3Z+G
eJ\8(I6K>bA#ZGNL4a3L\>H]a4W.a.&49\c2]S3J3[.8131\0)B3[W>/2ZKPKY50
=,R)#)[VJE?f0T[K-:fGAJ^HE=O?_P]YfgTA/cc7LA@U7MNcgB3<gKdPTa(,>4(e
5c@B2./NZ9/^71[aC\X_cPBN/65R_LaM=7<f8(fK95<;N+>4?94&@9Se9>^2#P1V
G&,/LdFa@0KRB86Z:DbAJa5X,L[aT#SG5K?[B7Q2(YaQ/L5XN;N05MWUC.:/Y:9,
?_V_e>/99Pg((@TZ\Be>WQ[Hc/;JY;V&VIA@K09[OT9[Q/0Z]dS#Y^OgRW.B:O.:
WeWR[\1-[PD8)/8P#c\=+0)Y4b]^E@g069Y0>7a2Xa]C&/>1c57_<33))e+J[H>-
X5&?/4:Fc/6a,CCU,V<:W^(ASef@H=;H[]?D5P6:[<]I9Q+8XV5^C-CMQ1(]O[&V
517?O>LR::Gg\HFTWZ#;;>.b-]1/EIH@(P)?Fgb@61JI#Z0c1P:HbL(+HcL.B+#W
G()Dac#Pa[OHC7OIBFGG@4R3NI#QgUFQQ3R&^W4DG68:edY6XbS+aUF2SNV1ZE:)
.PR4ZG;W_d^A\HfR^#Q9;&[bYXC.;/WMX\=b6bg60]GeA-L^7^)JDJMWdLIF)BII
G7AaP]KG6]7.U\3<C&A+?.OCDQWdDPYb#9^3?H-@#8/BN&QG/=GDg#N#+H0CPUN8
3RNFC;6JI,&\AB,)8N<T:<6N>PJS#8I.-QTP\?LU(VZ9G-@^_>&L8RKQH);5N9Sg
2NKW1NUI1NgZ80+e4J?B[PQ-QG.Z5:[M/f(-U7=)WP;-ZQH:BXf0?S,U5^7=/:G&
PD,W-.]YA,Xa0-eTO7/<IEZQSP;42HNM0ebJ\M[_VJ(ZNN[9f4_YAKa@-M/\Da<4
:(;A:NKCRO+EB.X[5T9@#)P8,Y:?65Z@MVOYY>8C5VW\4(@?@D7+SD1_2UEISS.G
2+g=N3_2P7ALJ,Q);F1.DMO4VEcCM0WWf=)cSf9D<=7_];G-1T\O>K^>/<)?IH_#
bJXEWK5=B?4KWNS9=E&(a@F?a+U7#H[ccb1J)YDR=_-_4&U5:.DJ[UP85DTcQaTT
J&&I>54Z)8SX5/3.848&NO^)JeB95&;d3JZR^@g2:e8FRGEEJTdDD3JD&_,:K0&;
T2&:GGFAHgM-3dVMV:2fP:eR=[Af=FG<M]1(E8),ZYKA_dQ:0b\)fWW>^,<R[4Yg
d@Oa..PCUM[Z4bF@^5\0(Ib=N^af7Q<1==OO;8FQ)^;AcUaU6_6KaO&QM;b.UU_7
.SAZ#2[DYVLHJ6/7QG^4&4HQMUQ;\I0M[9K3XD<>H?:e_85NAN[3bgNF)[fKF\5H
HYIa^[97L14W#]E+PY@>c^4e3FJc=GS.)I3.QeM^??CW&I+V(+MM)CUXCaER<@XB
#R&W]TTa;65TeDdcJ,:;[b]e.]YA5X9=<W9WBDMUfXd3LgZ8NJ75Qb0&1Ff^]&Qe
;G>O\C/P[>C7&NR0W7R^K;=2BVT\N9a5IPgJdJ;_SKDRJA#IA>6GU7S/[I)C?fC;
76;Z:2G;f&)-f/VCaN_e3Ya10V6W7/\I@bBU2gFA-/BgPK?7M:L(fa\,+N[SN,CV
(#QIBBP6<I)IcXC-8,D=01R8^L>Q[_:1?XK=,)(EK)=KH;_JQTe\:]37\_L+TWQ]
3]fV?\R.R9LbNLITTNG_YeKC0;b]4N6X[\ZU6aN?=e1-TPHG+VM79=D++4=,(cH/
7MVB3UF?GE-;DIe/E]5^3;^+NK6X+f/JL5AJ35+CNCD2T)&EdX4S_>@].K>O/ZYK
-c.?3@[<WRQYeQ7.U[H.S39N/OAd>UOf7[1DM=F^=R]MQZA<eJWKBM3?:K31;OPX
87FEA#:GK5efS^[=WHD7VL/9OY+U=KI?^H,90XAR.75-:9Yc_;\A1,I6+bS3DgSA
M(EG_0#6aRDRMG]55cVc4[BC+<aLPb0dg>FMg4)Sa_JfU8M#@d980/#<K#>gaHg:
aGNP1O[B5NZKRWR+V^.E;:IHO(IB;AW;38N.WaQHJ(6<BE\,BVT8[5,.4<?FcX@^
Y/HUXMM4;TLR34-5@-0WaV=1<;=Ma@NgH(7UIRVIN@I]&\OVeeLX1>K/H=O:\GbZ
1V;YIYWdUN.6e/8ddF\fC^+dI2b2C&8YFZ<IAQVX3\FN4aXVHZKJ(@(7=9./1\;_
0W\aVR20WD_06+^8],G=<a=OPIIENG?eb/\>(AD0O/OW>3&)dd>R@bY9V)O@c+GM
97S#@DPMYSFJ,d[WZ7gLLTQ^5O:GEIb5/=J]GF<;e1:1X)=53g#Tb\/YbXXVf4I7
MOA8O;_UCS0&#]=dFJf7(4&ef8JQO9Z1?HH-[D2>eVH;66DDbE6?,[?RcX[-\Y/G
LXFJIaMgVZ&05JD2,C:M#:cW/^2(T#YYQ6R@T?eKcP,g<V.>O^MgQ(e>FQ&11-/M
DR52QH4a2;:(BAP[X5]2bD,Z>3;1&aYGI4DRGd#S3L+]&NQNb&6@A>1c/TAFA3R9
D/>U5L#[\^]9,HEK^I8R,_W;@KO61//^Hd-:dHV7.)U))f/dVA/,2B_H;a0f][Q8
\5G)Z>GXSFP3B,>@-LBK&KR>J;Ha.I8GOg8.ZO487LKT)<f39HdFZJDEf89#9b1M
eP,R.0<Td=1YgKS@8U0;]V^g.@P8&KM<:#<#0.BF:c0\^Qb\M4-G/.b;6,BPO#+N
c[DH>fM&G5I2C+Q-4RDXe3/0\S[C8UB3P@OeU+A6?>Q[G?9f-Qf.)JYbXR^b392Q
D4OO;9@B\A]T:ONH_F-V5(4ggEBPE)O&3D0DOQ\UE[)+5&0649(&KSA3\R6?FQ29
KCcF03U]&;5.[=3L60W+NCZ?VUGBJG><^I=aRC)GPPM.T?g4OfacJYc6\AEgD(e:
@S3d-QE6cG=ccC(#a-Y6cW,M++N1@>^NA\Z;Ig4FAGfEG7B921R3b33)3K,&?LJ-
=W)L.O<7Ag-gKdN,d4W@Af1e[1HI2M8HR\IIg(?FD)gVF4Te=TeSD[cU3+VAZ600
EXf4#d<B?I4^Y>^#^g3,ND6TECC4W&T2Y:F^XP,:9F9YC;W=OJG/Yg8>G6<-+C1(
:/f@NZG(PUNEU.[FG\W0#b5=CGKWTC.]SMS[_[.N,PcU+7D]H/2QV[JH_Q8JKaAA
2fbf5I3bWLI?Sf0g>K^XfIAWf+E6:3._)X3Og6@\LW[S:=4]C.:7e1J?Z7^3)JQD
KKCP4LO;2)UR@S;._F3ffMB/EU_(Z918H;W;6BGfPd5]/G=+I[f3P)86_;@4Ga.@
Q1?]AS#M\/b,8Y)<7gG)K68\^D&)&Lc5IJ_#3<NX5,b-dH^=KO0VcZf4K9?73VX3
0781519Z=H-^[LZ<Eb3gN+^HUGAH?g_?ZW-.KNHfCIO@K9\#<dB<F:FZS,Nc/+IT
][S;Ve/f6&ZGgO#?TA1d3.D6[:cMSJbSM3XSc70fLSA?2cafV35[g?3JYS\cRR5;
dcf[9;-e?A<C?-E2X2^SFEf/fBRbFXE>3T,SFed&#[7(3)VEBU/H^aab1X_<[\Aa
6g&f.ZA,;6Ee],7\ea2(#(&,S\2=]bU:SLF,7T\@XR#,Eb(18&Q,@M4+-ed[>+[^
.K\9A,K?0R#>\AW@)@b,@RgT<B^-J.P6M\BCECa@f]=,3[cFa)Y]6R\D2G7G#MU7
HS]^SQST/fL682]_5d+#>8<E[J];F.Q_b[7&3?G[X0KP3^BRO>+AGN@##)Yd^T,c
]Z)[bFA5+761M@>QbSce+=_SL_LS0@NT(21R?K?WXDMK8J/9V\-J13(M=b]f+]KF
\afPYd3g/+C>]K13\XF-F^5083==46CefUQNGX]0[FC1Xa]AbSU\V)WF?Rf=V(38
+Y]Le]EE\2&4:^RC5d/UAE2:K.O9-K5GG4<5MDL(dWG.J.dM1.ba)LCaW^[S@-T4
TBKUB):/?bf-LZRP<FTJ0c#:?+gNBUW>D8T\7dFS]HJ_TL8REJEV#a^aISdBaI#Z
baZ3\85+PK#RC+@L2TE<3J]AZ5f\V@a@.G/R<L#F7\1N(?WP5(IR<\\K/#[W]_H\
968a7+:;,N#^)B554QNT4]?EFWBRY:KL\?VD\-B>\1M9A-=L^Abf3M/0](B(#Q74
]fY8FF08/C7ZVb/7BDT9/[A&C^Wb\NF&>gD&H82(7TJO][OP,FLJG(cPIY]C<O;D
(@DN;[FK85#JE\:C#GC>0)f#WeJ^cE;5Gf_B5:>UTBG5BROO[g4P761HcB-Hg&P]
,TY0eJAKTPC(cM<NV1fa@;QHXH17K@OS/8cOYN;&FW9?1J?0Zc3&9Ca/HF8C<35?
7P\Z+^?QD,AOB;ZY3YF9d7DG[H>GL-SSC9T^Z0>E@ZG(NabMC7e[<788&aCCO7CJ
0JWI-:Pe&5Z0+G0gBH+bc\TGRHZ=&1Od-5c-4c+>[.()22L-<-4\>+IgXB6.]+M)
3Z42]6X9NJ/PCK5\V>;X?V\=;]GGX&KbP:Y0b)+?(,I]T?N0-?V1-AVOOcgGPE(R
\MBab;AD2MSWVH#G[CNKXIggIS_\4(WI.V9.>=X8OQ]4\aG+c99&N1R\A\XE5MA\
;GCA4E[J+-(G2HF?WD:XS?c-S=JY4g\8BI-13V0_#G)>LYb7/\3WA;RdXYZYNe4(
GO^d?Zg2JT]X2B>[64#>8-B,X1B6P\L?R(/EcaH4+d+U/F?b<&JbK9cC65egcF)J
#cK=<SY6/1_,;BT5cb]bON,-A;,f;7=gU[&4Ha[V/)/R-D8#OC39_^(d9[dM-@]2
N?N2bDc>=cfUX6>cegDWfHdF3/+UbUU\b<f-\P:0:O<UHLa?6:4ML47MMZde-XT=
X1Le381IXdW#-2_Pfa7Z8TP66\:+HW<<7-_EM0QI#c2[^3PfN8aS=/G;GLN0dfa1
<;4J<Z^@cbQ-IP/RaPJ9@PAESf;S.AT4F9aBZf0BVG@LZU6[@c98GYAJ7WJbY2DP
]8(Z>PbHGX1Y)7+B?S6I=7(39YaM.AFgTdSV].-0YR1\^D^;(\f?BUb_d1aKB4Na
8YLXY,eVU@N??/N>1Z8#^NB])P&8_e^Q9(;8.:DC.JLF>23HVNHQ(.ESbQ=IgTZV
V.9ZZ(Kcf\d7YP.b9JM4_0e_OM2&)fE+4O:XB.9KE27_9KGW].UVYF[^;:97S#fK
e&4Z(/Q8HJR7NV-PAbCb5XNbOP2B0I+X=Y\\](I1R)<Y8G@UbO5)H)aBd&A-/Acg
NNRRNbX>5./]+b7Kb7a)-##)HR(OVcQ@,[201e(2^VI7R@E2[NXIXYI9fc]PN#&=
ZIdK.O,(5Z&9:(@>RcL7,N/eGM^TG)D;e.&RI=]GSES>..K3LE5:K48cTPM;QG-1
]\,cJMf(LE>O7fCc0bD6CD.ESR9S+6M]GQ)2SMK2LIOOZG6cH/2R/E;8]eHFKQU4
QGEA;?e(AY:3eSLdb<47.JLfR77:Ge+f6JSOYIH[ZFS?eR@-T>?MM4VPA1[e#-0&
<FJ<T3WI)[Uc(\]RA^D(@Eg89O;FH/L5FS6L@T\&[:(+W8_/GGC_GHV=F&0LX+9Y
9/(G_QQXJLW&XFRK4Ld;7+5bbQYe:E+55U^5L\)V5]2R,1AKK4M.c_&aT[>3T^fN
GBNK1cD4a5#f,dYUI[<>XL(79?BCS@>@,B]]7],&R0E@8J4:O@G>O?/e8+AO?FTg
9-C_H.)JEQgDPTH[Zd>bH_#UN_C_..37&PREDGSHfZPS@JP:PYS3=Ogd,OF7T]Bb
X,@^O-/2d8X3Od0CN_>.@&4da^_(),B&8Y01TcFd;L;CVN?EW)Fc.XI[2A\&#N6K
BI-V)(J2ag:(C&-)De2gFYXbEB9TS]&3Ia[?a23])b16JO=(fJ;,Tb_[7&=K?RIL
M,7_>43SZ[Ee>V(HZB4[X]dU33RQLc?(C/3Oc[__D_]ROV37NX\+B6MJV[f:FWV)
U#\E+E^b#:]P/GbXC.Ne6:^T7=.g]@9CVfPSSJAH3a@+1B.FJ\,D^+_I&aS/U77;
(AeATZ^dUA]EJISMCFP=_M[?)?@?:?[cP^#?0Zc;1R?cK7=PD5d@RE+3?+aBGJ\g
2ZT@1L\P9Gg#.M6Z/dNFXHS,,b?\4V5^LgSEZXN[/_XX9-gKG8#GQTU:K[N))-(Y
AI@H[ZJ3-J;O1L<1#TVD572R/Xc+-7>U2H[2L5YK^1#]LFRZA--VLD6^e#JZ8eb:
T&[-]+14YeL+F[Z?USNN8;OMVbG.MZLE-(9e,Z\EAd.Z.R2/3#KCbG&WFd0&[?\A
KRS]5XP@/1_-e?L_F\\=RQ\HKbZ=+\_fB>?)H[&a?1O1c9TLFVgU&U^9d=1KYGX=
#c[N_8V\J]cGNA8T6>6X\EU=Xe?=&+D=dRfQA+;SKQ-I36g3B+>#S:cMT5\6U_OV
0YaZ9+S\6(2[EfC;R56B.^OKcE/7J#<RYd;-[-=LC<:U?a\B&/:))>Z2f#EgDPeN
;Ig8e;cAW;UR^X[F)\;@d9<+@D._Pgd74.DEYC=fPcI(;;&N[;=8T.1T/FD@>]?J
e;f5I539d&\/@U8.aBC8Xg5?6V-0B3ZU9-:bVY08)^)Mca6[H+&dT3X)@6:.fcaZ
USL0H677?EE+dJdRFLS0@fDW-=LZ32ON(c1S6Q1E/M?>QNV072P0?)0O_dI(PR?#
=SI:CV3c2+7fF3[YZD.<Z]/;Y^K2>.<0[+YKRN:<6?fJKQaMc_5Pb[cQ[MUc;Cg+
dD1ee.IX@6T>f^0X:/a;P4PF#-^^#9QDC,O1OJ,A7KTa+Q=BfbX5MU7KYEb^a/\G
5E)PKG8/c[1?-#VVEVE5UF<&:.YZH-_g;7CeF#e,?+2Q<X4Y/GH(?Oeec=4UW.c<
Z7C/VC3=e;f^5X](P>gOB^>c2O8&NP[K4)#=@d?9,?E8138b<+(,ZL4)L>\KG[SF
b_^::b+SR2KF.VP_A4(N[DKXQ?FJR_=3NBF6VDZ8_1(>1^)Q?M]ZBZffa_]J13R3
7RS.2d)S>]DW@;4(,O[I6CUc:2^\G7:4g0.;HWgZGDWIM8CdZ\H.f4EH5I6O5&&+
PUN00R2M]O&TCGef<aM[fR5Bb0G7B?M74fA,+J[Pg[;UI/J7#V<]\T>O-?)MJ9<g
7^4\<EJ+8e=PO+6+I5V[DB(DQ9J9B\bX93YLI@XLN3R.[6<LWfR5R1&;7-15MG=N
YLF_:-Z/?@3g?4K6Fc&9DdcV4<3YA0Daa9_bHaAbERHF\=_d:>OS;CZU+F[SYXF?
(;CIb#O=WSXO:/^3f@?\+8;C32(E@c6#OE_<66cOZI>UFSfc0,6Ke.P.Z+BdIB([
6EBUA?Y17K?4UbP9X&P8<b9Y@(8C(.&CK)bJV@#0E&OJ(4@)XR.6)eJEVW_6+A.V
9(Z4WUSb;6T#LG&ZKLI34fLPVRf/U#deJ;W\YbAe_cXGDY69T/SW.\)Z3R.geMV7
17P.M;+(.8Jb&.T5(3]J9>H:],[083>=_.5C.X.eE>^gFM8W.X+9(ZAP[2]N?-V&
TM,70aE?)aZaf#WQH5MYBWQ4S:RL)<0GSB-NE+N]EW+>6SO3SEIeYMKAK/O7W,99
cGaV_WTV[LaYTP.?I&cPcN&&-=DH5Y3baXBU7(c)6;T.e8:#(cMB8E,PE;USUZa/
3,G1?=HaScHA;3/1N/_Ta>/0ESObCE+:NI+C\J]AD=eb^Pg2]9MBa_\A1V4=:]#.
]c2@\6ZH74&=cQ_EbX8+S+Z:A(bC;TT-.YFUU:6P[]34]VMK4\3.8g/YgI:3HU>S
A(QN1-D8]L^[0??(@C/]8_CB:c=>,GMEI(Yb)65WY6KC3aV1c.1F1B0:PSFbL]g-
RYPG9>Q&[UP_F;cVXG.A_XO8R9=8EAIJ3-;L2&M<G8KM/2<BU=&N.9N#FR,A^K9-
#2/T&X/c8J_RM8.^+5GKcX+\F66F<f-LCTC&EKY5gQ4\;^Tc+5eFeHA\2,H5KaNC
PP)]VcM,X[:2_f=d3U2e/BTc8:A8^fDeT1-27agNa2\URKM8eZ>XOKGVP\R?(Ba<
5K7::;aP8DG(F?b?5KK\ZG1=@S.?7A<Z[Mcdg7#QA95GDZM.TX,5P,DEK+Nb#Q+<
.B_FLL<gKO20c9&cT>f]PLb>#I\+S_XP<<],_7ES1fgXZSd/W6,@^79UNP^)/)64
=f)K[39D6E\O.V3P:affReRc8L2+@5VD03c6\LW1=:CK.D1Ef\31KaQCAQ;d>6+f
((AV9)geR)OJI#>2(8)CK>A;f)]</U]]U0CY#..CcAEc2f^HUcWW4KP?[>9fEbb_
LO3UQ&B+8K[@,U19E]?F#@UAg[.ZFE:]ceObEL28X0F(^\02^d@O/PI[U6RE;#J.
7>D9R^08e&ACF8=7BA<:ZT]NgS;+VFBR\e1OD0#F9>L[-1]VeTFfE.KKG\B3,b=H
^dW#He3=[-TQ3B&gFMLSE?1@R+P@L?=TEH2:;]0C^e4G^^FW3X0LWZ@Vb^YA)F>:
MgAM<L&NQG+0)BZc\.CI.b@]15IE&4?242K_4+NOTX4J5,R[&I&GG5RJ1[f.)4W(
X(+9_8cC(J?SX#1eP)HaNF?LS2[;/gI@6JZd25RCBJMbI;PVg,U57<R4OU;:ea0P
T4]KcFZN<Td.P<1&Dd-8Hc^EAV?7adH3UOHAUeWV93509YX<e)MKAX089MQ]XM?/
3._H1_-Y>c5V-4I>7@aS/20:]&U>KL#=JZc/HXW>PNaC(;GMLa(^MULQD0#B1]9<
H;b\E=D72de\593g8B>XaFg;V=@UD=&_[[WUIa;C(X[JCfK3\N-H^/P2?_D&<7_S
V0Z8JOV;@>;+W<E/4CAA4fDN>XI9c\/UT@O[:#P,:RI&2ME@bd4=K?8_&.F;@4(\
V.M\NL,0C2aJ6OWLSf-SF_P#]07;>SFcI@eZ,1\F0&NKdD=Q-6.BCT23^<dBS,KC
fcP_T8_dE]:(4g8^Q-&g@?8^IA+XO>M6d^Ze1N]#CJ;E;4)Kd<C#9,)L<+5/d>F=
+[(BH[EBK_XWF9aT?7JYT^Z>eA3/)X=5DQBDP19e:5JKB(/dNG-(^a@e,06Z&XYe
ZNSA2d&#cG;<0(8D-U[OU.G>NEKW+9-0O5:4R8Za5ScC/baL4\ACD-(DO_QT[SeC
gd_g(6[fO-<fB^g_FC6O?McSScO5g0YOX2@gN(45:OJGI.8#U,WW4Rf&)TN@fTaT
-HUaOH7#:C/H;#5VVEZBR42-/bTFMC3B)M]Rf.WECOf-2Tfg@AP<#?RDTgEe9&eZ
W>fG\<_],RKW\V/Zf/RGSDUC6g1=\6L(<BKEW>Ia]3J78YX#AHYJQ-_f0U<=+553
e@C_;_dO@-MNP<-1bLNdH?7T3GJ+G\=^SE<XBW+d\6eZ7LV>9V51YZVO>8Na7Q?.
),KE@#I^aSMR\=MC#Q,[Vea/FH)+H0Rb1bXO[d>Cd-V\e#<>AGg89T?HF[J+f6:Z
)#7&ZL/-4cG]D=?G9,,LBFZV7H0T;_?IJYQ0.J\<U.J?GU)e-b3/8;0eVJT>V-NI
<XVbGWc(5eNV\VV)WIR.GEM]8OV,?V7O38V9\EV3e>?b1:aF_CG04;FTV4#<)N0e
B&&_&G)5#.GaK/fWA/FASXF28J6G^F(_1YEG7B&C3SfcN[(egC+Z-4;:ZC(@L[@?
a4-U/.RZ00<>TL_G7a5A3GV-Xb5d^Aa)0#A5WS=N0=0VU-bb_.9U&AQ41G#F(IQ,
V#13:SSF>60QI/e81fbY@a^/TP>YZ7M^E(=5I]#WF\N3EKT,SZ_7c,]PP#3M^)ab
YIM5@HNbe5#;T\5D&G+?D\0WMBc:fOaDC&L1,]C,TdZ@Q0/?@=41-7Z?B>N&?a)X
Fc-(6VbJXR4[<I>Me-C49B4EAS119++(c_5[<<RKGM\<N#RL]8HeG9T9bAUbZa-#
^/5R5VK>]B=NbB=<_5D(+(gLfJQ8?9XXB@&,KC)N^7S>28dL;PRa[J6C.d[_587g
g301+&&(2-#W<Yaa4)VU/+7V/S02a.I+f<0@S>_KX@D:L@bB7;bM]6S@=8_:V>&8
4EY3/<OHUKN+1MPCB6[KD);>0=>dYSMc-3M>UVdA9TI<eT2L80WbV),#::N(,_TD
9,?^)dQ]A@/EeMCR+\U[1:Rd2JbL-0T@HL:J=f@,H_QXec\2WYM@[I#dAOdS\XCM
PTG?HgK1Gg#3FX];@^Z>_3ZGO;TP>D\;^2,BfaC5PJ&.Ja]cY=8@T;<9<J@H(XN9
F3=BW/<=LR7OY3VHOA7WMWJ(@=5b7S_HJ<&dO91__Q[Y9V<c/EP]]?77G=T:Q359
MPW;;U@I/b2HX40]Q1[RXV#0__,Hc_?fV[\)6ID,Kf@[P(R2C5a:6a-8cdVfC/LN
X.XT=.Ve4g_1R[,H@-Q:5_9@>+J&(WZ#2Pg3AMW-\]SRK5cY5JLA9^IF=bYX5(8;
9V[2.;f2Ga?2e2c#W0W2G.7RX5^FY<K3A#E07HCKB+U(A]Cd(;gK?O,VA,6gDEH^
;K7QeG)/SP#&BZ3:&=LAS729W8YPS\:]7>#Q_(,Z[2H3:bSa=VOH9b_IL4S,H)I2
1U42BC\9.JE4#,N3c\0432YS;\T39YWFL2.Q:Ka@E/C?,03bH1;4I+HPO5>K4SSR
>U&R+9J]c:VQB@]ae\9Z+=.CYWCMQSN,3?0H;S-_g)8I<3V-7S3Fe6P?#_F5US)Q
O8.[Fa8S@9?=a5[E>H?#.+=G#KVQ:?R>TB^cF:VdFNg<06Wf;TUNY:RBa;1_7_H>
(]+:M8BBGC2BH?WRDW=<J^[Q+AJ6F21N0?)gVJ(\I+c>8M779T#>VIbQfOdHELHH
XT#BMOY,GH05G0;](N:K_:R(,5JVR>6:7PaT,Xfc##PVACY]eb+N+BY^?,?KXEP?
@/#8>^BO6BMN0<:9c74J#VgP2V:(;?8DT:JN.5W;MLE&SHD[MEIa5HQL^=W=<Q@S
IS-5UUY>>-6<8M1[cY./6&&F-H,O>N(FcSTZNXA;8\AHNI#F_eA=K:afcOfNdR\(
B<6.]>X+P[^\P]_.[b[Ba\+W+PL?fB#FVEERZaB5dXZg-/P.6YH(\UHg7+36Q0#;
GHFB&ECEO^4:>>D2+BfQV[b/D(06Q?B7R<VC<\,0Ta9c^]IPRc5aN.3352AP[P<]
:aBTO3ZSUDW;:]KDE<3+9ZQQM0G=NO.]_M=#,J+Tf&f>Ra+.(&4]a/,@Q:/+H3TJ
PH9T[\O.7>fKW[I&?G:R^1+2a/S15dd)R:O&DT65eUC&<9BEd(PD&OYWH;MU#J1T
<8OQRY?(D.+TFU9WAG3IH>_acSFTJ#D>^WS(U9C>4T:2gc_-_eTC=GKDW8IM9e:A
0b2GK6_HcdcNF492YfDb/MZO2Qg8H,JZ\R(4bO_K+BPcCI=<5-?U;Z&=Kb6;_gS\
JSeVR)b^F-DB/,>W6+EERMJ7YP=gBMI.FCJ_@JcL(b08L-&6W52d,?&dC:Y0DF12
:TRP)aS_N<JJ6HH8VdW=b[4K?A(;)GTOFP6C9X380:I.,gK_O1SDae&U2[34c@QP
IB\cFZQ=CLa=CLJ9])N.:^fDe1#WFaV_[dAKOb0K3<=M6BDa/KM#D/CeHHY:#OA3
.-]KGS9JTc,BS<dXd(Y72YCN<,Zd[-L=.5L95?POKOOdIaQO<Be9&-Ba]1(+>b)4
U_;_ZD>?2;gTGU>cfDda&c/TL)BFOBEU]eS=#Ga&7@J>;Sb]:R0FIX</)f=H;G-R
&,Y;-@31/Ya=434SeQ1aU9WG/#cd\C,.N4LN1V8)7I8DMFOYML5?@]_V3[,8E=g,
+WfN-d(gVOC?HB4cLFg8eX3APL?1ME.eK7D3bK^(V0f.O/MS,CfIL)(H[d(dF-#0
<.)A(4aJ\XD_.)YY\L+d,+#B_>bGWf:4PT<Q(M).JC69dZ?McCJ&LKDP;(fSB1[O
,PT&FVG-3Be^bSgVE=]PIZD=QM;5b97:aQ&Q,Z2:Y#9N4?5B&_OW>Y3T5bP&LL_-
4MP6XBT;E1cH,X6X+g#7cXM3F<)5RV2O54V^-]7B05N1O1;-SM<4aY;e-NOJ-;[G
@H,[:<KDeZ-f;0I/@90@6WS:3XWIa\MRE<YABB7;?<]cJ?dH.@_:-T/-8]PVZg+<
_DPBN5Z+KT^+[JP2#90#5QBV[9A8L6WV.MTU5.I;3\7;(g<d\aHWL0Me>P#ACESZ
IG-R1b:FB3/)1/62f7M.DbaXKc1L:U>P<[X(_@UY5:E_g^<06bKQ[42c4]G:G,X5
]M,@8.97;:=G:6VTCeTV770&,2DK,5Y9Ka[&<6]<MTG-^YPRBMUTZeEH@]6WD/<2
2#[7@67<^HeSR<HNEPVZUK[a&T02Rdg0(@[RQ7W/5=,d+bc?d(V8B6NDE_I_76BV
I&,U[?@\^S\H:c@@Ee8X[7eO)PSSW5Q:Oc#^Bd//Z57TLb-c,>ebY-bI3AO,D/L/
/\8@R5(FfO^gS^=1abe?BIUL475=?f>:U-_=H+UG(C?c4.>S0QbFcF4R./QgJ0I;
.#X_WUM[N=7@/@QfcV^dA2Lc.X>=4_SS\Cg7LB/:I:Hf;WGTWAT;M3c6)@7P,L,M
gF\]FGV&.eUG2[.RQ7c55cHgHaYVPTb[@J;N@ZP1H#7Ne=]_H]3(Aa4/-[IVO<6Q
W37JZ.VW;a4U#EBS;F\YC[8;K2L(P^Z70BTegBSN\f.>N(7aBYROF=_d-F,22O,M
N-KGbC]=4GXSdRd=8.Ee./?70.2f5b<)L&>d<=486FgQ]2P[S)6?6YU#bMK:A6B7
5P5C#<Ia#]:.](.+M_OY[QD(+.Acfg)U6WPR-gg<RH5AF0@XO=R4;L-<7Gc8X+9S
LI2SgF[Y3CX9&f9YDLG_H>5KW1#9\[@4FAE=M[+5#TQ9.d1U6f([0#3J9U1bgKKZ
)@L.&.d/d=RYSANQccI;OB<H[Db8N<e#SJNPY6;H\dQ##;C?cL7F/(57bW4_^@Gf
I6\4;aAY?R#WUb\1#a]YC3VKGS9<eGB5g8#Me_T9ba\)+>,0J@KQ,;_FRIdN;g,\
DP/)7K)4@4V(O8X:&ZVJf#1,:#PFPeCW2R0>AW\Z142]0&EXY9SDbSK?URDP?BLP
#a7E11-#LX2W3cQR\OdSO6=IJ^@L0VHLO[LRf:ID@B0ID<EQ4Gf/RU1ZUV6UB+O_
^ZU_2MR+6eUaD6BA816+.bg[BYe]N\d>ZG179_/,KSXT67X>)UFU?K4b6T<DGbbM
TU3Q:\bR,+34N(bQ6VY3(#&82IW(\^a)4T)Mg9T7AaP@<,g-@&3A3c_1P;^E\de4
fDKW\3\Y_2&\(:&>EB;aG[9R4d):UO]bD2(MO&5GfJ@#46T1O9cU(-fJ2a+c=6/R
(aU=AQ-eAB1/gKK-3b;J07AeUa1JUU79K^Hb-U]4H7>TX)##OF(@RLA=c,G_CC4P
SM#MJa^&8PAWA^f+=[g>+F383R_&J?dY+TYMbI[[_)_JZBD@9_3/=C0D^CZWJ9>7
CbU+Ja?=:6YS\39FDB?7\-@7QSCM1=.Z@J<K=+3OM)TGLIe#DTAK6F3b[0N4:K-C
06\ED>GK@L05K.,4T@IBQNAbU/C?O2?bVdV5=e<gUZ[EaJK#e6JU[D+>)G_gUZfK
<F-REX.S#NDBA/8IX,+/.]&?5e6RA^+fbIFeZU4d-gP\?V+/(UL2<e@RSLfE^)4E
B+7@^VV9<bF+>J88K(M)A2QUCWRKB:MJ>FVAd0OH/^bJDINc5SH62FeX.SP+ZC?X
M-aHK&[a95[Q#^\EG4\3O9NPTP4U_;d-U+M+).DfdLcU-&Bbg<e>/8?LFT5+>1&R
>^70TY,J5\NcD?0A_AVEM.b-W0]=d6DWed#TL,Y]S^2L]eQQCe#Y(Le<a0Xg,(+_
:+&F@Ce70,Za?=M(_;R=2PP;99?);M_^-eUZS/a+;;MbUPfM9-P\dW:?c(1W9A[;
dJf:2L9]E5K#cTTLED=N,:80[&N#H-B;&F\Td.GR/QeQ?Ue+?;+\B_9GL@4L,AV9
JfeUZ87d62(@^/HU+A^.JQb=HYcePebP=<L5I?&#MHU>?Oa;aW2d)14b(_cHea;b
)O&S.aM;>,7-N8Zd2XfY2DC=]]g4^^^H-N/VZ5B\LESFN+RN9cI\;#0932f#)+?#
^NIOIOcOcd:@X-Z:0+5(7=55#14E0M&A[R0&=+=X;aFN_FG\bKbTIMLZ>^UID5fD
RWCZX1d=DL)MH6)(Y\&0c\,bH79<OMD.<aP1>1gAR=HTKQT#H?U9K_N1eF9?__.f
b+(#FDU\P^+)9][b.D/(eI6b;BFg;2[]e._9+>BCPT1M0RLLR-@4f-A<,890\_#7
[5\V4f4?]IO+X)gRSF6K958/>=7V\gFQa_IDG3(0Qg#,BPYLWPX.0gI^?V6A+]?f
RS1>1)DKJ[W1;a#>[_)P;7?[#2dG9FQ/d<K1D+#@2EAJ02aAXD>V\E@&7/STXTbI
gQ]f6<:^)0X8dDBQ6R.7gJNE7[OJ01=ASJ,(J=LL^J)]1/G2cOXTI@W4PT3E/VcC
Z-)Wf_F\Ib;SSEVTTdJ263Y3PIDF4_X;4L\6Ka^4:6gddNScOUI+?71GJ3aGPg2[
6@T]XTCESY,f0Wc(XV6+_]\0.N_\I;GW#J#7Q4TPF6D7dfffVBagI31B:P>fWHOG
;KO#[3T,<^@JT4I&;.R]_GZ<[<:YLWN-@KY[JXV_<-.8U32?WHVN,BGD15\YT/=L
?L7&P5BZWJW.+d=+.&,b+,&1B5M]2;F7O,V)\^f5ZH[@L(T,Oc^DObA8LZ_]B)Q8
8H<3XLd51SF1G<8@R^R)N^SI/=;L9:faBQ.\4T&RHMB;_MY/a=MZ?47(AW2L0@[N
<\)43Q]2@d[B0FRZ^,N4,,3L,<8-)1J_,ZR(91PCfHb#CLTOPegH(AAN^MMOT7P]
K-)E]PKWU<D.R/;cM5,HX[-2,DS:8(..37PD9I]+OW^d:E>?5JbWCIK2]PJ6Z7GF
-9?)GD8IKRgZE9-dPg[\QY=V-.X#G0/9JaVO:JB2fINH_fE8(K-9VE_HR+@:eN7I
E^5CL@G?4[Q)_7INUN&;X9?/Z737V^IY].RcU@V1-K./MN/(?f8+??P&044R:04G
ZJZcYaKF5JS32W;S6dS_\N[6+.>I_KN2XAfNH(\2Z2X9Ma30(M4g42E;V#A?/_,>
M3J&I(0-Oa48U+[JZJ]_/EOL_?>>QLdU#P+2X<PQI]fB1e+E)--.IW#>JB2_cR/R
QF^;,(f-<?OHU==b=6LDLIXd+K\WK@>U<UR4L_U3PK@0@Rb9H_.S#b-RV4W4TW91
b?TB9U7&F:3JB/B1WGS7cB.S,5_XfcDUR0R3M+9fcX[6I)?eNH[],CAUQ(gHQK1K
U@-6LSYE4gLMAB_9G3F<R(YD+0Rad<IIJ4H1F\SZ-+EWNaQI0434521g;S&L@&Z\
UN40e(8K>/B^(Oc9RgU(315,e/+U7XB3V9H.P>GL#^S9\SW<e)W+;TgY46\a2:YT
.9d3J^@fN=TG5eaV;5eV/+3&A:C&NNAKT-M;[fQ/D+3YLRbff64]D;XCHMV_JJU1
&C^/-.YNNX^EDO_a8fO]HP3<=#S#),;+KC#3D&BP?PTNRD:_HfOBI.,(?>?@ML;R
KXeX(P)QJV/GM<3@&ZRS@AFQB9BOIfcQ1dg)^9B^>FWaV6aaLMBPCDX(5QL3]Yd)
V.6SaTJ1<53]AWHC<<(>/E4M-2UX-;^2C(5OTb/6a-0,NXGbY.2I]@SOODP@fY9f
4-0cbUC&B;\KPNB9R05+3I9,a-AKC1>T6:MHZFZ\.g@8-5H45U_X6:0?0>R:IL5c
QROUCJ40G=R2Me-]>2Q/H=)>K_#[=9I3@DDY7P1Y;gY8XVN15@H3R1O7>-)71S_Y
P2COa0@>/3+a?W+H)EHg<0XU;Ab^_/FKe?7aH3UPbGBQ=QEHAf:,.OY<K_\CA&W2
f+9M[#eL]PW,7J]M9C-5ZaPZdaU.DEM;E>7/5P1&O<T0&;#4I,)YLV#e8dF>=d/H
D\MA516a&3U3:@0U&^O2CS+SP>B]<<IYce2;=-6D/d,<Z9A^)Td=+X;9(J<?6LAe
2<-/WQ0bcA^\56AI0?1QDN#5&/U&1&+(2dc<S]:f&CbY-=W<+C>,W45()RL#;bWC
3>.0)b/&#W?/_UFaM5UK-F0NX.<U5G_fK.3KHXa<&86VF(J;U89)dZ_M9If]&&;K
&#.\SMQaQ3afW]HTg&aJFb243[1-TK#a:O9eUJ9b+JVC>8O.4FUNJRS]9FO6K>GU
Oc10Y&^gfL]c1CC)cF0,7I);?B=Nd8A2_3>GS0d^S<1KGN@7fg9I]A)K.[:CWG-8
Yb(1NE9>TSfYe;OU(KQPHeSG:L;?_IN?cX)+PO1N4N@W>_MI5MAKQFJ4&+9EeF@&
=D_-F@Q:WSX,SF&ca[TDJV\8L4];.4^UF)M4f7B&^fH=ZS:^ZJA[1P>=2X7EV0U[
.3?.6ON0d?B=GU7LTJ9bCe,VO(T#9A(BA;@Qg;A=^(/QPT7adIMAYO0ZB4XA5.[U
H03]?dd51/+eAR,=7(fc2LYP&CD8:H_O5Af;,K\K.H]6OcTLc7#eNa\0Ad^&.7PS
J&PW];8[9S^FW@=Lc1;M#Q??1@DP16?G1K3ER:_RL^,IeL7U7HACfOGY^-d9LDNU
R]50K8?(&daV:Q@A9MM+WC>Y4)eeZ=If>@P=0,S];]R1GA4]RL[c3-<LAGMZ@C2a
JHe\KgdH)9c1&+-J47=?JAL+[IU?Nb/+L#)+@\(&\,BJRH.#DI^KbDT5,C=?^WXa
]\;g83-86EU,V[:@(J=,II-J?eI#>V7TeQbVN&7KZ9#08Yb,U2<@)OEF3C\0X4Md
C>8ZVe9&,YfQZT2d_1ZPg;a#Ed.Y]+2(/VSA4J8&X/YXXgURg2dDV\OS)&A#PR\]
,38:HZUeR&1c\)QR9#>:FN-&?#+\VA,-B-79+2U1FI(2C9YYL1K=8]BdZ\9Y7aQ7
eD2V=O1ZMD<#86W^\40eC+XPaT(M)U.6(=9>ZY;<A6O/?T=ZGbL#_[04;Q#DN\+J
(2A(_=RMeY>I)fMU-@-5S;[;)D\LXeZ@)@9>K.9GSGdU1;M_4XKQZQ3ccSW:RFD8
,-.7PA.:P1)8K#8+W\gfFRP:NZ3@=VPP1;4_-6K6(_+81_BB_RXAXcN)a.Mf]aJd
Q<+P@;GG4,F>5P.\E<.#(:@_4CcF53MEeRQNBdGL&3<-\aXa6YPNI-1<N-eB+Iaa
XW,Gf8f;Yg^f?-]cNQQRJ)RTPF+/:D+MZCF:6MF20dW4f_;dP&U<?^S-M#I0NNeM
_5ZBb/G]_<)bONa]a<N=^61b6\7KD,?5f/-06F81EQ,/b_U:IR@@9aWWg.87I97C
)O_H^Ta+0#.e^(-<OR0_?\,P.c127&dI(;<77XT[ZH=.#W@00.FDdV_K57R,D)XN
FH(g+KE/BMV#&)LWcKgaGUdX&U8fH&H5YZAee8HR[+;Fb-)3]_&@9<AU?/ENA_-[
_XII1N&T]9HJ_3/;/[<.,BJ3-EKYbA5,./cZc+.3D)0P6Y44b)/@UKU&c>8;G/PC
[2?G/H2]UNHeQ?H,f>+-Z[FLM2)1KFMPfO,8F<c]N6dPTBH<S=Jd=]RJL9Y]^L],
H.C;g8#0g@=X/c/\-&6aJe>5ZI75_G1e506A<gUN_QcJBZ/Pg,Bd^_B0.8V/R8Jc
,d,4<P()+XdZ76@U(D;2S3R5Y7d-Mc;9,ZE8Rc6J]O0DN^Ice61\E,fC^6I)T][)
ZY79YMES?G4^e,VM)X,(FQ[Z>23T,#P(NO<5(7W;bM16E3R>[FQBLT?g3-Y+;]VI
gZL>H[>C(PY_LQUZL(VWHN),0GYL0-Z4TP-X&0Fb.;__T.>Z]XY#];:6R143g;45
.VU8O7GT/>ZI]aYCD>UKeR#F\1B1<F/A#,(N30FEOK2??O1Q2QNT7.[M:FcFfTQ?
8NZK(.8QbG@0#1_#eZ@W10Zdd8=>?19#Z,Z1g,_<6Qc<a;;b9.(J-eE.WE0?<7)=
[:>LF7Q=JHRf0_KF]ZP^&A-Z9+T&f>S-](e=IN:H<&(dVgf1Od)gB-9)-Z[?gaa+
2MO<f25M6^N+:?-66E-EPU_C0KI?LGB-/.b.50)UA1BE+CScbICdVf((ESEO\+N,
e#?WP/(fDAgA\eMRR:KRXcK;:8:Q;I#=??g9,5^J=U&4I:Gb-4bOZ3>+P7eKHgcd
]XG[feHP:.6+,[Ie[_gaV&5N8-d(XPRFYQLQ0Z0Z92I3a)UMR;WZZ[>RJJ)T89N\
]E=\^=;=Ic:(-@0<EFbeY\)ObDQdD4L2)>4^<G<U90SbVZ>ML.W>;gHA(+J88Y3\
D8bcD^:2Hb]cA#J/=UAK12gTS=g\;]f6F\H5RDEJ,>WW[)KI<2.TM@8-IB.URPTg
[F>b-52Je:G6(f6_9)Ma[>4.Da^EfYg)NWB9c#ZS]7LCa()2Za^Y7agI4;g&KX06
3Y4/1?E^/+OV6#A#3N<;,DNJH8U>TWMK#;=[4RRB^6dCC>D-d1=;(KdA3MU>U##A
Vc)7)\F#+F8e[_9-PP[Q--?62\/e,aBSC2]][a1@5Y]M/<XRTX)=V)Q@e4&DPe5=
)@I>ZG#0ZMA/\>6(,#;T/XJLCCdN#]111-#,UF59F#@;V@gJEM0QFE\YY/+aJ>A#
B/I?U-)SUV;W15RPIEWVeM3O8I[WVW_;3<<G?K_>d?<QNJJL[?JY6R+><K_=YMS<
Q6/@9[^]K0R\@W7AEB4cF\d#+@X>MRQYTd?U7H0Z-U+ER?ERLQaUF1d44AS];:+:
e>>/Fg2Cc6FW6WSS0WV[&D^P1VGbAZ>MZ2?.;_\I@6;.BaZH-^3+KN8@X]J4N7_7
/WIeS4,RPeE.ZLQRZ^3EUFg:7cB>^P&^U,Z3SJ5_NF^0#LJ[\.Dd,gAQ82F44BTe
DI6a_f3AG8[DNDWX&K(4b/MFbb5\#\8Q,?U54X,W=8-W(b-0Ea&XH98O<d+f#7Og
4f.WW@[F)+0YY.=XNc#.R/B&OHbZbA0\MK^_+F_BZ-..(_IWKDW2R3A^5AC_#CJE
I6\N:ILKB^SNSeUJLG+)S6H1EBRE=7AY6P6d._O5Gg?YV0;\WgNIIQET#M>@bEJG
4UK4L7K?gNT7WM\?&P7EV]=,P29YBf(RT6<g<BTg6J8<bdG-,a^/[c&F_,)JFWSC
EAdX-:(TTddK>@Fb_9X/IE8],D.D[YffM7=+XfO1>C5Wa^_BG8IU_/e7:7AI<F,1
MVgIHMc??Z36WG\J4#??JW1LH?_aLR_Y<UDPf=LXf3D;T536/R4D/JZB]F-ZBZ_R
TWX)caB9YMLBI<;VT9\D\AV^b90eMeHKL2\e_YY8?9X-#B0YTO-)6gJcU[@0,6L]
Tcf/1IM1EOH<4Y/bCDP6)H4)F[@QXL&#.Z\Z72fXOD/FE=:G^JE;fH?]PJgCM)1\
O>SOC]&6??3O\RMUaBE4A94RR^TgY9PNTCQ:V\+X2Q:@4;F_WV4MT3L1&3F]0f],
7TFgSg>PR/A[KZZ9a;;:B8\.a#<I+[LKb3GKPQXI^bIZ0Yba7NS3<9J>=Z-:A,>@
TY5ZXO=SL6DaLZ7U#f(.TVcYXf;848Z<eIcK].?R/#bGC48NG\YKg@BY82S1YT?9
>gebRK[<WH^+:\Wd/-+AYV#_]/]XcR17)/,+\)6#-Dd9XM)T=G3F[07JO\\JXM7,
dJ^TJ#X^S8ZE@)2A;3gDKD?Hf<))&gO&IZ)0<YTY9PFB>GP&7aP=\GABa0Z&fV)9
>@&6/<[QdT5cUWK-X8,&,LVZKDSKObSRZW&K,g1_36U]2V_6-eQF#EJf;E,+Sf[V
>()I0g2B4+-R>.cZ94>/8eg;EKWFIES+I<Je,P)K_;\5<4V1,5KL]PBG//c:A=#3
c#gSLT2](CG\.IcP,?e[&Z7D:-M?8#a_I45-&.\H3+3-CMBW<=:U&F_)KS\<SP?T
\26EB61&,\6?58]WFJBf6L[)&MBb&]RTFc::(-JQ.^0&=<Lg+cSbTXOC1RNX4-?0
=6bBNPfJL]TX=bF9aDK^8.08IZ[ZbeN4S=XP.R(&.1Q[a(Bc2E==BIXSd3V?61L,
F_9CH1MY=QNVJ1[FW#AY\2\]?S?P+fgQ;[7FDaH7YYW:D8OI\?1cOC?-F0/C-IE5
=TJ0GZbNe>cZ^6(DT>J6F/\2.^:8FDd56;R/_L7XO_EgRNfEg<;X@X]>R5FO>_LM
Z=7)\S(5?]>>Va-=L^TF&?-e(H.cC&XCRL7,aJH2a/\/5U+(?J4[+94NV]4-ILfZ
G&Ag07GQ,aNKb2gIET(FGY1M8P#.+D^9^V4aJ^Y+>.=,,)&CNGM4S^.>fT?IKJ)f
<H7XL]+Y3NE;_#GLRZ7]1SB)UL^e)+=HP,/EW::#OPb_JgDE3HUG4(c\NE7/=2HX
?#d,Y0U7K+aSC/C?gUS&?DGA9TSc7R4L&7#>0Q4RKG\-[JW;S\U/T:(#(S5V2O6H
4KPI:QC=#U[@38(O+^NI-,XE&gAA)E8c8.U2YYaa(Z0bg.BI,Y^?^:d+OL\N+G1+
5-a3EXVFQSW:5Ng_K_.:2R^63/eE(CbGZ^KOX=Gc-MWJBIEY#,>#a8>.W:B_9QgN
-^N#OTF>[4?M<RfASXE(c@dIXOA/,8@-/f;\(Z<GT688G..2[L1cE+;c,Z+\(Le\
e/Y3LGa?g[OSb3C8K98KgH+5DY@Fea9-R<Td_<DU)O7<)e,D\+c<-A_A,Z@VTVMa
X_-O441+Z-,?2=Y]aV@UV^[b<OD[[=#H=PFU(46>+6;WW>?;_-.]Y:D8W3b@)]RA
S^WUVJ3PNR>@1,EQ>9BL/Q3EERfg/14&b+.8[+&6A@cJg#a5>[QC)R&a/[(1,+.K
+1-6,9ZIM=).<9ZM+GC\KIg7:CJ==KI2cR5E^PV5;RbCd?3D.@L/6@&LLG/<Q6&,
,=S-8g/&[CO.;)^0?6:EaC6+)-J@V;M.7bf@7S2EI9.;)\0feE&?_P\A+65&M8HO
\LX/NPAR,bB>a0],AU,(YdfV)LR[3I8ZO7_OS+aATU4C^+b&XUgURZG2OH5)aT:E
I;fA_c]BQ?@E+>9g/PP+UEX#GX#VDWX;Q=a^WG2cVeN])0.I7\?;g>aF\a5eY>7E
(-OW[2e0KDTP;eI>SKg&1ISGGF)]U;6L[AL\IEIdHTQe:9U^0&P8_EGgcA@UCF)?
]RX@Y\P4O>I/U6cbKZ/\T?7-+^eAgNTeVZe_\d9Xg9^7&f:>;LWLH6Z^E6]gW/6K
VS5N]2300)3a5/B1+:Y=7FW\RL/cW:D[G;f0YW(Z]0UF1g2G,MH&-??K.=U_D][Z
Y(1gJJ;&](fX8Z74_CJHA#eQ&<9FXI\UQfT&1A7-Q>WXXBA3UM-ASA#(e]ZD[@UO
Jf@U)fcSA9/15Y_4R.;UAdY[+,4)b,_4NL<?;9<,YQc9?1e,1+c#^@OVe1b>Ha5J
Ja+,XUSB:=T7]ELgVEe/OYC,BEJV]8=D.T;]COgBUUH6]&B,W(c>KF59D;&/BE[Q
4)_G=.;6KGN\OfV;H11B#^<cP1+fXGH(-2YP4KD@YP,C>b=J\4DL7-0-?CP136)&
?@LA@-#C[g\]KJf\.8U=6aK4f;3Y@R@4.3TQ-A^QM+=QL\/B>X=bg&E,X[0eCUcL
R:1[f]=071X+09M#XO?e)8TGZ7.Q=N8BH6b>15TaS-SU50CZLUg61L?U0QX1PAFd
R0WIVON:+L>SMNSDD]He7GES7eM,C:/,SbP0BV\_NG1Sf^f..2SfQTG(7Ze<SC>(
,(&R<SO/57O\Be/1MABaHI#ZD+&O4YK>GgF>LRgTY>dS86L>,+0eZF)TN0<#8(2g
;Y3USD,d5&;;<YY6D(R+^DD\K#acb_fU/&Ca4;O1ASXHaZG^If5X(^9AIFN_]5f3
eQ1O0JIOVcO@&cKc4Z.H=3\L)1A1b82##5e#M59AP5@325[8(9>Y[7)aP.M.fFLM
1,e3\S\:Z7bJ]W]4?8(<N6\HC4)X&^>Q3L&JJLELXA:W7gIVecX9&B2S<[HC>51&
WK9>E?]&Jd25_&(9T46eE:d\HK5S,U;WOXe^.+@?^8G0:.FO?YWE1T3I[=\ZAA\O
S&U1M&+552:5,2E+>P[/7(UW=fRB_,gG2b+T):<M]>XdT2V?36P&8?R-ZC-TUI,]
\#M?>VWHP;X&<)f-ZQNV5DFUBSYP2960e\8VIe1;)]392R]X.+4V-9b8dK7f_SEg
D]#gN^dJO=fRYN2fINSHH9K>a?,=);LZG_-HO6b+aU+UL5Q:M8[a1HZ@\D/6UcJ3
W]4619-f2;@L2C[85,D^01/BF@R+Z=L9]1,Y\Wf4fMdK\c66LfJW;H9-[Y&)WKeL
W[?LDE^>CV0W2K?;CS#gWc_J90H6EDA;)M104XD-,5gSCKN4IH/5.&GGQ-D1g[WK
>,QQPceS<O?TGF)JQTRf\[f:YQWWJ?f2VG?-=F)(b3Z5#/1@O6A=>6P#EX#8P+V&
d(&?D=_T8AUb4Q+GfRTOFU)6/>/;@2D5^d=R&3?.-V3BU>N#X^M]KD>VE_>a-ZG,
PY(+115]b>@AFN(C3/#8gdS+e8)GPM=G42R))-.ODFU5A<=Q#+bBX8?4:L7QIPG]
<?+HOZWbZOgS#&B/,)B1f,F].=cQUAe/Q+P=/f^)&I5^^+ED.Y?I>BT1.E-f3DZV
:NL9R_Q2a(\9e=RK?F6Ye6).;eGQT\_FLbCNN;;4gP[WS=)gfSJ6\JV;aVO-+<(M
_9Z5f/W_GTa?,6gf#H34-3<>JKFXT?H;:#>\Cc[\&SYdb>&U9-;]G)WFU1H;,gMc
Ac?4FQKB<0]5R9YU))g\./#b:Ne()fD:&[.S:d,G(1ALf0P>;(d)?^5OH(D31:W/
ag/gK/=0A6/FUd)+_\YdM<S4E3)H<PW],+-X+)3?_Gc2ce(bgW0V.77=C(>9H(PF
0?-^^JR@::X4b<>b8Id8QHNG?9BW4(YWa3e^7HZaY\>=.YgM3AAD5#&4ZY;Z\#FK
=P[;.EC\7LCaE7>Z=a:g6[HH]G33L^4+>7D+,g8.C5Hc)U6<WJ3SIJJV,Kg9_VD@
B7V:C6,)e3>ZZ>a0AeP;Se<LHLT1=Y0RJ+b_KHD(MOZ73@K6g<3_W>6:>1YM8]OE
Y1>Q,H2<3Ig&\\T(e<R#PE1Q:A@L66[e\@U4RTHFT)Y]GY7A<f(_=)QN=HW/IfN_
f4O^bJ=5N(@:V(TMH<P-OLJEAQYGQI58DfG@eI:<cccGOD&F/8[V?3<+PR-Me-/E
8[?_/^V/V>dgJ;LPCfSXE&eCYb.-cHF,;C;<G@.@?UK)&gBTCON9?.UaEZ1#PVGP
&=d_4#bf)_(a^Ic,[B5HQ2+#3>]+Y0eYS06NGX6?<5G3KW/>S1[=D4[DH07RcSB,
:7W9ZUQ:T]<I8bGY#V[VZ8SS4@GF(N+dSbWMQ#WfT;79:-Q&V(Z)8<9R1d,QdL^@
We/T#6JG>YEeXDBQ9.\Ya+(:7.g(-=)6bYV6U7M5&BSL+/=E.,WUgEb1Q<_HWeCT
fd287QJSFHSN5]V3[g9OF(ORFII=8SK?@-_9R?-J#2_b\RIbd2B\QU:DfZH<)<Z;
2[3G2NbV=TA5,.e_M9P7V@3Jg0&Jc9fBEXb?0GMZECT?+B40fe-gbIe]2XPNIS7M
RPJ.L@<,WHeUY9]7ZCANYF6)KOWaPT+V5G/QZFGH>6cGWbDaFC^;#5>F.M[a.;I&
DSgAQ-C@R4IZF@6:T&Qaa4;a2OXY.d(ZNYCd6M@IIWH1CcaD8BWFV,7?D-c,LF[8
T>9fHA;\V@72<8Ve]SaB@.MG/8H3]B)/)K(B4_U5N/]4D>4#5JX4V:^,#c_YEZC4
D#5e35TVIbcC^X5>F]VMgUUY:+F8b6DB6&.X[E[\HCJ,ZdT5J_HD(>46MVB=RZR<
D]CP:XXAXPU8I;J;CJ>U\6/&8Ca]L[-M+\Q:<,?L<WM@[,fF@Y-:Z2.&/eW-6CH5
fW8aQFO#+)HJBEID,0c+Q,HgD=>AB_DXV#_/<FS?<.<]Z6<-HR13/:[_967AAT:=
+)M8VgO;?#^b[X-P_;Ge=A5O,SFP.YMV]3&If/H:+BCU=/OE;W)Ve)P5I)U8-:#]
f+gQ29D)W.EYbeR\=)RDSCE:^O/-C4a>Y]dNIeH.)2+53M?]aIdVEW.c,)S.]GgL
([B5S.F(;?_:<K-<DQg>CFef<KD0IJJYO)fCDfIKO#TN[:/7A?31=-dB_I:/3dI+
SRD7NW8PU>JF2\A1IFF2AW,#<04KFYb/2bU:_W8O9K/YH+EeV;O&?^_HBK@.K)BP
g7:EDCP]eK>G2NR+JcdP?);&37C#-(-6#7E>H&;O9/C(3B..BbI4^BJ0QUAL6AI3
2)\PP(\6c2YMa=:OZ^Q.AZ]:13TV=+E>/6J++B-9/4UEfJQ#g7_G=EMZD3BfD)X7
<8/(ZBaJIE7K8T?OQ38Ua7OM;2@>WYI>Q>?,1fgV9@4N_Z&((>C3N35aGV>VF,)-
-f4[G/O[Y8X/5.Q>R^+=d+>GSOJ+:YM^&]=1/LS4LWH@C)/cN.@8)+[#0/S?]_MX
C]-M^b\@d9]V>Yg,P89.TL&:NFT3;VbLbBA)X?EM=fC0:4Y@]B(V<:.+_P)Yd&-2
e(L,DST.a_d]aYWScCY51VG32=<Jf#7K_D;=d#MJ5(^5IFT_=C28CU#6=MA5))VU
7;;UW)0#c28<]fc@J33Yge/5UR6e_B&Q8P:.8L6LF6\)Y]7Yeg)QUM:WV/AV@5>e
GDCZ=NW<Y&NBd=D[HKeaM1L]TU1E[UNEe3-Ad^BKe4)0N&0@X73C2KeH4;?705U=
(Ibc8&)bN9O;N>6N>)cc.Ua>a7IB;-7,HNcA+0SYJXDZ@<W1LJ0=1N]CcB\/F::\
Z.0(XT1bc.=41,#5L@L2BBQYB=.(\@JNc1(aDYAZ7#(L_[V=>4?b\\e(J:?I_8BC
?7J(QZB&<YL:XB<)233=V:.M3CgB=0VN4M9ZITW.Y2RGRQ=[V/O1_SBgg#aIfM/2
UOBaVGe=T70&VYH3VTa]&g+V?c-F92]ET]FD1cOL1MX-GbR+V>#=7)J^Z>4gF#>.
d<(_59(G8R6UM?_9N;Pgf5>=,BJFT9QcF]9YD>aSag/3CJ>=)3QOQfTa<]+=MLR7
W@]9Zf4[.RbZcCFM/+g5A8>4If2TR)HN=5g?\J>Pb4SIN2-JbV)eYDc@;7H5LNON
NG?KG&WM/+]e+P#@[HQX&DRT+\WML&+?FLMF3KL4^@.f&eIZWNH[H2DL]CaI>@K8
B\e;6\TTPTcB<f_YQ-4/N=0M-NX8O5_aX4YGNQE^CS3T\R:N[EgLL9HCJ>T@8KG+
\g:VK.+<UIL8/2Q\J=;(26]7fCb\Dbe3HXTNOc,..f904#V,8X?IVf8PbHYX1G=G
6>NUUM&I/TZJ#HA?&TESa:@Z8H6FE+B\a=1[6QF6-bI6)d#@Be8DfF:J;6&K1FVM
&LMY1T.SK8TdSJ9gdSJI.F::F]C,/TFD.53Tf1S[V/9fNQIV<+#(S[_Q/S78MB:,
&1b.[f-LE;XD[KQ=SR\]4aC&_,E;+T/_HIUOeb2-(4#OVKa2O[H9VDD8;TeBg0_e
6YQ.>0O/bAfG:H]^8\Gc^DE(5f8+Y.1b-BdB4E+.IH^T2YF.@-#d2&cSB:\?1P6C
_gK=7IA5SYT2O?T#]feE5/bUS.54:T(19BO=7^1CX7X&eGO/6BH@:TX6Z,:,U2KJ
HR&_ePbIEO4I8U)DNIU;-[=MP&4_8S:+e?9d\YSN:Cc@R=CZERNLgS11G;H9bUfB
I0,](TUMbc>BDE51<<4U\Ug<cCP@f=D[RgK>XFOc<SeL/CI0<f_Q>N<3da^JdB3T
+=ZYALGKQ@?9.;JI2\c6]K+QJaaP7bC6-JHWR^>T4B3-RVO77IZM3G:\AB/(D,&C
gb;/7.-aM-L[:c,SaOPLd7^7A;&=3\:>Y0/4LZe70b/,aOg\Qa.f<@T0)@.^G^#I
_8e,_(DJUOK-f=MABaa>CYR\>EK(_fe+,Qc#>HWOT],K3;9@]Q@7D;N1Q/DE[M8b
2T-U#AGKI?Ka&76N1WW)E_e+(QV/M:-J;>D.-a2?+LCOEN&fE\S&K-&1+J^[\R,E
]gE[BaY(#D0;.8R,\\cId-X9Ag\b?-HD3=BcHYZ+=N64&B]>Q;d9cIa=UV#,:Nc#
LWXR=@Hf_LUM(V]VRbBR6N+3R<5O[Q<<d)VDL9<&K@740O(&0?/;JeYb>K7A^?A8
RY7CVDU&(gQaM_L#H(f[WZA^:gZ;VBYa88&+;YI.)CH(Y[#fQOAK)af8O@9E(8;-
X/O@MX]I0eV.F&/K+\+2CVE&>-JHcDX165<.0^FL-&SFTR1K1gA+.H&ag.&X,;a>
B]G:/gZ=7]8.G^8JF:I7/:F)\5;C#G>EAT,5d.LU6VS#_P>/PQIIIa?fUCD2ZX,4
NeD1BT_-4XYW,ge^DU+(-OTQ0dNZ3+\(FeS8L;^BU]R>VWWT;IF9G-&BCGX2T^aM
V+g1<]942daCW6>0S.\g3ZHT=F7YJ3E?4PH\B[bX>8=GE_c2BB4Eb(M9#21Z=-dJ
.BUW.8\B\6CVgC(;?M(fN@R5JR\1?KS0\6b1;1<If6;@HBB@M_GAB0-9:g&,@V4K
&#V,b3J,9Cd#Qa>\8D99bR.Z\/P/OUW)b;,#(<1N4^;IUN;2[9d->HO1O8Z7JSe,
<#W-=TaRNW3Ag3O9O33;98<<>4aJV<W4=Y6:FI-H6M:eC55F\T1<2(DHe8cbZE6Y
1UaJ:Q0OgDcZ<Q-7)7OI;<D.cFV3(HC_I\,D@g.[?2;W@A4L)Pe:Y/>T3:7H]^0.
8-NH)JI;M:GB79f^N,J\eFg#M+<K(ZD9C5Nbd@66Bc)V,1Y24/W)5bc_F7N]X>M]
33T,25cZ4Vgb0Yb>4CHa1:9b]LNd=EEYaV,K44\^5H?ZF/S,-9Q7)eC\5.1+>)9I
,]&W&I,2Q#e=AQ^B@J@A8JUJ<;8,F3c<TB#;W7Z6GK(M+<>9DD3[a78;G.:#LO)F
Ug6>FOC=3?KgH9(&\9;)4\g>,gf/>0^.ZAZZdT/BK-SH0^c]YLdF:g?J<XU#M-a6
8d0e2@U&5Me&U&d1#5Y>Pd4])R7P?XdO.eZ&7BO.]+2[2O[,6f9/d=IUg<Sb8\>b
C+L&)^L=&((/-0(\7JT=^#]-4T5G38J69D[/[H,BeIK:?V1)23YcOJ/Zc^<)6/@_
IWOQC,cO-=)Z()fM;GY#K;C7C=<I<I-&P<EOC=9NSYEY4A3]Jf)()-DQ4Paa@N]f
?&L<VAAcHdWV>M3S??8DH;MP&/\B2_YC2Z2JL:20VFTd^Jb=Z9[,?4,DP&+N/KVc
e+b_ZGL3,3[LUWgcR\UgNAYD\-/,4.T9,bDg5>ER]KL;C0GgC51/-TU3/f7+P:-9
SeFA3>0Og8H#N9YW-@]NBB4DF-#Hf1YS&ff,@@6I(Ic4R+RC7&7Zc^?>+HN/E:P:
;CY0[dH:6+DSWH/N?\UBEc4&Q0J<F9(de+e_R<S910OA9)84J?_^_G>44WUaC](^
CQIdDX=#]bZb9HG3@=_#X@MDeRB)T1A6Z.VFeDSRT1(1NTKJ.dDLX@Eb14&<]B)9
SASV&S-;Q@U,\EBd8Y(@&-gZ8eVI]-29T]>H_:^WMaP8B+/7(?gD^/eXW2Teg:#T
WK[GA6)aMC@K8S;&FBW28f(^E/NGX^^e\;BDX]?G]g,#&E2Q+VIV<Rb.E#(dba^d
-,Ae_C:f\e(;eAHJS+T.VFbcV+76OB/0-.3\K6aR,?4N;BP^^f[=7U,8H5BQ>(#J
KT+GI<&3L\N?OA7@(J35//]K5-:2],AK&^,#,PW11:D(,(P.V.K/KQR2P\;4eZ52
A8G23S=B]T<e-(BTVdPEWJF7G&52VbL\g<A_:5^SMJ^;PD(]f3/MT(0,b/1g;Tf+
]:;@D3HW]5&c4Ng8;OfS8K^V.0(aVD6+V2>>4,]f2#\7F.,WE#\eS.b]K>9LG7;)
&13g_R=TdZA7ST,2g6J)YDM./8H@1Y3VaJJ)VY)?;N)E.WK>bL^\#5)SL#].\RIO
RLUA5K[C_W9#=&?X1QCABQV.N9\,JFJf3Y+H/HL-f4[Zae44<a2B/af[,6Ub6^)9
89&JZM/AHL62IFaZKA?<NfO]I</-QD8Z?d.6d@:/\>10#Y45[/XXYT5,e+]#\>b7
E/WF^(d(IV5_AI08H470@\<_+K/NccaULZ#,3SF:GAB=b-MW=[))]A,\U(^W1IKX
CCLPf(5YYSXeN\9FIMM/41=:HFg^[cZgCN(H-6:F<7M.BO=I8K&2D683PO_#7&YX
7#7+4TKRZQIY+P2/#3a2aWA^7>6f?Q@?KS4;=?afT-.F6e@VM^;Y^;T>E^W7DSH,
/Ga,D#<<4V6LJgEZ;G[W9EA2,&EW6L2LHb^CEa(I9])J8JLTb==Q.U[EcB_75K0^
B,>NM^aO,HTS&Y8.42eA/@AG8-9JP;^cCI6I>&<II&T-eF7I@:O,\)c1(f3XMS[U
EUg@(=:0273U3Y(8EXH310BSHLaJcIZdC+?f83YKNEa^Ta@W]CS/BU\6@+4Sc.RP
/RQfRU;2@ScWfK\X;NfY.C;dRe>,gSR95OVd+Bc_HPUZ6dfL(]_:(PQ3@>H?FgIV
DPW\Xgc8CIXJ3:9Y.],QR86M35V,6,-9\-Q4@FF#E^4B==g8g7/S6Zc6Y76H/V/<
<=F3_8-4Fc\AbYf+<-C;V>Bbd@/YU1OBc2&OVEPP-MRfS6\RF(.f[69(D\V0J;@K
KWPRdS/6_aF3F;([b)T/AU._)8/3P2E_BX&gCcJL.Ja5@.<BMXf<\=89-R7MIE;5
XJ<GAgJ(VfL#/X:D+:#YBBXZe=UGC\edAT(5RU1:#(-ZZ(>^+AK)1bNWBg5\>BVC
;LAb<C/_X-)+0LKIJ30)U9bTaB9(8/ef736?Zf2/W(b_/aJMC8)=1_Gg]9U&X(5U
1:UEeFLd_dGP-50_6][gQZ2eE/&1[5((X_I7]O_JU&[W3[&T^>&I[\:d&@Dac0aW
.YF9+BGV6EWZH-DY\/63-[e<E4S0<d]8X)ZMBa=T71#U#VX9T9AeC47\E7S:Dg_7
Y3E@)Vb;OeNH0>01N=H0_N2H/C^(6]fF73OM-?#2LU74COO9@F1K?K8af15fQ3)D
(c>,D:9K-)Yd?ZBb/e)P11VE/>8fFW=SUK]@[@f):31X;+@a/&B\<EH>\G6X]-eL
NJSA==VYL0EE>[?T>Oe=8=24D9+HY9a^\C\[a-8AI_56[Q^P+;?#955&deO=-1T:
D&T@:aMG_X5WRfFP4.BA4H;b>U:b2T&GW-&E/7083>Ta^?.1WZ)2QYNN7.WS([M]
Z_=6D;Wa0:]#eKSP1_ZH7]ScP>2G5P6;,7(-9d>fA1SKO6#=UZUJO#E(G^efHJ1A
YAJ^O5f_f=,P,:;8N&OSbCRCF=C&[BN/++]8cdgKGf_Te9+FA3W/eWY)c#Yd9PWe
&9g@<2GA)f3._0<1^6XL]eU<^GcSF^1=d--.2a]ZR<1H&MfH&4BOM9OQe8Jd#@5f
6/bE<Z9&OBF=M)D^F[SOfN<6(dWWOD=cQ_R=]==B^M<H^,Y8OR3dJYGK?M4,E580
WcJ7KP3,P/J6c42#S8UF9M2FL0U7@#d9WS#)K:g;FDC<>J.7;_>]^d4&KWfY;XLb
\HS(KCKAYIRAL5F11PF(,8cKBQ.^4H;TLWQI&S).J9=ST=+H6/PI?/NS1TdXV01Q
U+P,Z&S-78&M-:D791O(\9SJ[;6NRWHZR30O+L\DOc_)HT-2_:TC_]GC5Y>@0YRU
IP2&HGE_D=7,DQYK?ZD:_Pgf._YK9^OZTR<_TO@74eVK9:7>38dQ0;I4XA3TAEB.
;Y;5OMgJUb)C<\P]:J,)/(303Ha5=CGA0N>/]Ef<@DE-RI6DGXJ^bNU\D91RR[W:
4PcC-A9D#LcF3J&35B\)SI3T+(7CBO(/AgNR&R^PA=<8)\RA/Q6Y.X/)(/-FRC=&
3J\B7(.5WaS6Ke?URFKgU^RI&9><[b:@PJVFRPXE84_&cN7\I727&EgRR^2G,0(@
#e?CBYRfcLL/(:65CO>[4HZ/Y+gY7[OC,9&4Z\2HV^+&D+9A/FeVES=SWb=NG:XJ
3)58#34/X3AFUK]QS;@=9;5[GBe+-W:M,+Y...9V-UKAg.0c7L+Q_5df&bU(.4;M
EN2J69GDBeFUWZ8_4aSUD#16Xf].U5>eAe7K_YMRPa9FgA/Q<?acDBZ?MVG32&GA
7(f/d>K(1_W,?d<LCTdIF_YWE_0>WH([,?Ma#4b)<c/EZE</>J,NbDE]ZSd;1,:Q
fEGdFD6;YT9]K1g:6UecX?(ZBZ6D00L00KE?X6.?V<@]:LD)[0::.[^0Qf^E\2#V
bHS)>F4>Z&_e@0VE+J_&;F:^PZX(eIZ5?IXQLLSD?g#=S@3&MX(bV.GC2N5>Y<BZ
<N)(Y2dO)F?OD+3^7CYPTcCVP:ebeBXI@a59U?K7J#6D1eE6gg59-g^5>GD7g2#7
JK0a(1AFBYeO+7ba;Y\GW[BFF<)Qe8gd61MQ#/P/F=?WQ<2.=Q)5\,6HNHQC@_1,
c(D16_aN\gVO+E\2QcR:\K8a;eV(?Y]EST[IOb=b]6W@)LdER&W,\b26\\8NbbS\
83JaQb)7?UgGP+Oa<ON?F?,9^:Yc8XMJL<ecIY/g)_3?>5a-YOA0T,2Ig&.MNe)G
T2f/=B;VV9GWJLJXS(7D&g)O,5FF;aO2I7_dd?.60VQ8fNGa&]8259P:\M?XfMI0
Za&R4ITK8(G0(715SI1g?#(H=+KIAc#Vg&WH:O@8:ERB-NG_;E]8B@OU@+gRQe<g
A)WP>2H3WG^a6]V10/@N=aS_=:<gHVNO8Q5?FQ^gHG5]d(EI;:PV[7eadL6&92U0
=7OD<\:S:d2#9M1?Ob&_Se;gCF^DVF^D_-11^O=(VX3_4PWL5U2]>A&Ma_E5(P62
3MVOM/MHFHG,eXc\fRb/:9&;e]ETHLOWc,gW.I5LaVFQLI4E]QA[c)LOM#BHgUeW
4A6E^OJDG_Q7b_6D?<dDb32DR&#,a;JKE>&?b089[]=CDYJY:M/7Y^K,9R..O:Ud
d_ZL@8.5:FJ#,2,:B1)-f+DJUTH)2YOa#adT]QK/1[c0QLd4)TQSN(^2cDgU[H9_
+K)1^JJ?W&Z:&(aCRLcU))<4G/eDT7G(PbF;67XK)cC/@+_a23&_db(^ebRVCR=&
dNWNf?5G+;PdVRW,=d^XX(V+a72J\@)3g[f&-_8XS6.)=WCf6a[Y?#c_<b4UNKEd
D(N&;gO)b_H,>5;-A9TDGWXL0OJ:,P2Fe);0Ede0@+&XBbZVZf)5CM@fEN6c,W+f
DgY,I;F&fSWCA^gRD?/KF64=,FA2cNe<0R4-B9O#/K#PA@;d<VbR2>?9-?>0c-a1
(/PIRR_dX&I6VN9DXMD/S<a^]39,(HXOV[63O9<e-C]9<8We^85_0J93Z@PbL@,E
5GP+WFHP_=GR&^S&.O=/E9Rc0+L@G[-(7)9H_/)TT<:GSUI:R5.;6aF;UQZ0XC:6
=R+2[,@+fW2aI)e2X[+U@?K<7c#NEVAb#6_=a]Yc_d<Ye#A:#3/B-aBKW,WG<AVJ
dW9#P5G4#;UJ8Pg?E\VTf3L#3+Gf=G<dg@,Yad<2>M6MO)fXEX/R[2C(-&Yb>MMa
TPS)CRYf:13Ua\.=eU\@E)&H=YU6c7Qf0OY#0V7&,Hb&P@E,G+T3-b)\_\a2bID^
RUC@Xf<AJH34+23g1[fd+HYM4cQDYGg=(P9:G=d_G&K#N>2FA,F4,^<HO9\UY3E.
5)4O[gGA8K0Bf.:.cS.T&Y4CQ.J;OT&FF<:/^#<:&gJR-5+F8AA1=6Y+;Ue3Kb@5
H6UYbG8P+CMSXH32-CR(2IF:/M:;8],UU48HaLR\B7U<:0CQU:H-P;.4CXg;cB,d
E,#@-8P\dDB2=T@_/^8Ib(=/C883^LX8F<R/4+8UCI>=PH0[4=eG98Wb.g:7OEcWS$
`endprotected

`protected
#XRA9AHCI[VFc(3WRU0e<PJ3H&3Gcf,Lg1e()[1e3;f6K2^G(^O[/)\6S6H=#3/#
1AD2_1dEe+-F.$
`endprotected

//vcs_lic_vip_protect
  `protected
g^=I+_[3U+I,+A,32>=R2E<1dP<d4T[W9a)6G74=M.dU:?PgAAXf2(.b+BC7A,_K
[J\JK+3,dd2NJC/TM?1dN/0aJTVM-2g+O#S(RZF]&PLL2742F#3c5X4=TN.)#Ra:
9]@.+Pc<cc(>S>WRO[?E;)U7c+NC-Ud2R:+2g>H^,_O+:._Yg@8fW9.CHSEgNZeF
^MYK@I9U]<;E222ELEOLRaBI#TAO-;EI17(O)#BGY,dQ:GQEbLgS:Y.1)2#7)g[:
QS3_B&W\gY(9=L3E:G_a3#;>3QX=ggJ=.Qe:8U_2&TWY/11LD5>479@/AgWe#A_4
bI,3K:,6E)TdgJ&[W44Ig8<_cJ7<a0L6:^,@TcVRa)WJJPK2bMeZ9;)E&DX03J&/
:8G=,UP16OX:Lg9M.D8CfaWQ/Sd@=?cX]Z->XVG:5d^?R)E8.T>\5@2LF9d@E?&d
OA1b/HW.\VGEPaC,J;ObM93M0@Qc=IGV8SLHVSa.O,@VdB2fE:K]AAe_UA,HHJ6>
d<KB).b;?.8G[G9_gA#(dYMg,#5MLZZ9HXNAZ[W0Y2AV]R\+9-WOM:25H\H5D6HH
JIHKfL(>X)U9M)L;71O;1R>BB[EF[E?TCD3;J:a_)O<49V\2^bd6J#<0eG[ECPdM
<D&]f1>AdYCS&?9)_1KEBM&[]?_BQOE4^<58L5@Ra/Z#9.6DS+TI0/8ZEKKa,XLC
=I1J46Z+.HKRXI=W+@8^S8[@fAX59]DSa<e]cDXV\ZUbU[7?c&@:S;6SAX^0I.,Y
;O)6]3G3bfS#QFDQKSR<@V.(8J9723A[I4dKPNA]O(bLPT-FSM3Yf_NK8IKa+PEI
)-(H:X9K>+4S44U:aPX+2)IQM@@S:&=8>K#14<Y_^O^@B9Z+.N_Vg>FUW66N9_IA
RL@ZJ+;a3WQI,Q@]bU0]\\<=+S4RM&YBFDH4-L,VSP)agCI5>cF6@K.+]f)/45+-
&+a<-Y>bag<6MaQ6\=J[@OSE53>bTBJX>NfQW<^,@f#ASXZa_E2@OS#0(=:PW+g4
.6\)aW6:73;YIRC&/9d[fY5EV.#,SLUH>HR,TFZYV_N]ePM4HB+@F,d--d0E7FIR
ESS\3efB(3a7Af-N._)@IHXQ+)eW)_0M;1C+HbbaNATS:X-E0I?=.-Hb1CB_dfID
YgCDeeA&^--5QFS2D-XTS.^P#9G6WG:0K4(MN^OWBMU5/D8CBa9<^-#P2dV?JFN4
:FH4#gFa2?IUDAW/b@@T7GX^UR\OIbF&NUgI[^-PH0P+PP)H=b?2:<9T<O;L4X7g
:,+3,E8)H/P]?.1aLb;X0=MH<0,GU((7(?W3LD(R&0Jc-??Sc/IF[=8C,dFN>6eK
d64.RX]P.;RI]79@?IaMR6.[)_;(8YUM/:eCG^-a:OL-A-8C>fLJMRTFRM:<bZFS
2?MC=,R?-?M-0E3JB3Rea9>g].<U2P;4\4DgID>0,d4SW=P#?DBfMY@Z1^MbA\,&
>(W)1a6>R90MQcT(<[@bVZ58J4K;?#b(_77aMNe8ce>G26[OM+P0/Vc:IYD6)5X#
<FS7700OV1ZAdLE_JTL/^_A+9>c4F7CD0+g/][Q#LQY)WBYO)RV??2f>_;8WU_eC
0;UCZ^R4P6]\1KI7#0c9.I8-MK\T^WYIBPS50K\3B9GeF>:YHJ6aJK@[<P<875S9
;GD&5:&cPU@[M4/OGC8K._Cgc6Z1^P\f<0X#M;/F0@I#c]&DaW1H6LW\F830KLTN
Y&Lc()4;Da>\6A,;+3OSQ<,(^Q[;Ud<1P;X8edIJ7T1FZI@=VC91@G?PUSag<Vf#
A53)23)UE2)?=BQ&+@fe:UXZXXUE)O6TNcB]XPJ082@:=\:QOC&3NQ19?Bb\O>,a
D&86CY>[+G?K3.-1.=FV4&J9<4WKWXcgL#T@WO)#d93cL:R/O_U/ER)[=0LUc8b^
[I:[T;5;81W0,+@C/Q.BZegQ2+X[(JCFdQF/P]<dVF,bBd7eRe5\K)IbXVS9D#<1
b6.FH,a.(bE2B5aaLR+3(INT@PP\ECbR>4SMI2J&[[dU--9+&9S^K5(F-MGHH[W7
FNM;fLO6&-OD)W:,^d?Jd3Q\Z^_K,:-bGJfL<KX]^_&+@QC66B&D.;D7?SY#HI-_
ab_Z9[1KC]LU5_c@TT@Ja)_:#>Eb1=b;e406P37gM&L,^ceLZW81Qa^,H9;=JUY>
_[S&0)^/4:?H=]0YTeM>\5TUDNJgXE.+#VU&>1E.&1GdSZN&f[a?_W_S3Y]^X:>B
3(WGX&)[7XD.W:.(Y,1^/=aGP+=?KR9g.A^5L7TY5BAKZce),:?6#gG\^U\c/Kb>
8R(,4(\BdaJ]_CdOX0V#\?Y<]^-8329K.;NO)?f_B;_F[c^eO])c):IJ12SZ\8@U
V2WM26JSN;_H8Z1UQI94BUT\)A9\;\fL9]9/gBNSW+L4Z7.^.IWD38fMTEHL(8G9
NOH8RBBb4+.C9TWWBb6;I623?6/93Q()<>P;O;#dV?<&W9b@a.U/9eMB346AET(B
eAVB::MD3C+SR_2P1;W\8UAFHY1dRE6N<9SMd2PI6V#)2>9_.PLH=_-F\F;X,4b-
>d<//>W&\P^47Q=]UN0-[I;W=PXI<@7MN9#K&04/X:@->#d<M/JXe7XTOa[S:HQH
;Sf153_Dd@V442=C4,YL/IZFJS_9LEXKc7Dg>(3C7\^NfHI.<fBHGWP2<WA].;5b
MZIE3>YG+0P/N=ZS7#c&B1B5cb\WDgXLI+MRV9/f:<D81Fe_N<SNJ&:TZ@dTeEE[
GCO:DIH,/AC99KS@\PNaXGY<]f^DDU@WF7;J;:1dX2+6502&2YACCeFcSGYFP2_#
e@79<IVEdaW)_6f4,S2ZB(gbaT];cZ;&5#8@f?UQ>aG_P7@_N>?:cLD&f.a>:b]+
P08E?=31XS-V97f-b=>/3bO<Uc2fO;TVaDCM=IL8&cWN_SSE_F-e0A#AIWAU\PLA
NIeCP-#eg#=YYbdF=SO@+T15YaV@\<-@@a]58FRDS+NVJ7P=#.RW9,>cHgLG#JE>
\<.PFX]3TAf+0G<AB0ONIF1dSP^>b.@XK6]SZOC+^&3FY>g;b+D,7U>9Qf1,?T,&
=GNHE[ED7g,L8T[MVgS-&D.Q6?(BM6&]\MQgDcW[FcSZVM.]YHP:Te0a0[M783c^
>]+eZV2R,Q-BN_]W^1^)U;[I=2<99+.dO_HBC3R\MDHdgC?@I0)bH;ceFSORYUG9
;>cY_95U[(@^MO.DILR,ePMd[/6PP.][?Y[SR:14T\fVX0d80A_dOIU6027IC,3[
SWc.^+O=4<\=Z:#F>KVJ[>&-JcZTHNDCEVMgPFL)S)(bJ3N.F+ILPEWe&d177):P
cP1^HX;6(7OfdJ5(b<CdS5JWDK>0T.;&R.VGde([ZWK1/7L^X1Ue\3<Y\7Ig4N[c
W^AF1^0./WRgLdc0WOMdO[J:,W0^PKXEAJJ[A<aW#YV>J7Y3AV<Jf9D\c.:R183V
N#T&YXXdPYXD.FOAFE>NA2]L<&DJ1ES_L/d)CSBOEXK54DScbRKMGef.DgGa93Y5
Kb<[W\7NISS#[O6Z@(OAa563[c_F[GDI=[VC?gK\Y>J+&LNQI78PWaBF58<?)RE:
+L@1<\Z)a7M-.aWZXC&;),[UM,3)gc:<3D5RU8I->N<)@/7e_4=+>5OOXIgcO63+
7-EQ5dC0>.ffb3YIU4><MA\E_V:B7bb7H8IS)>F6K/V-EX3-H@MWcXZgP@G?2dU7
\^ZF&fg6UNDb2FZD0f<GYB@LB)^=)bVNIH8e-6PM0)fe14;13E8=B1&55.+;aI#T
0)XZEO2B/T[G8^W[]R_C=fOUC7&&eM1+O8=DF(26P;R]=H?#91AJNQ[KfSR/g6;M
<<K)0MQ95B[PZ5QWUK#G[f\0bcC7_L/W8PSCFGXPgKPMF4//(YOYY4fb/^J(LJN#
@@.^W/J2ENQ5PZVIe<a4VN1/X^7g2W+/d0#Q>1T1/FV@W?Q6J]ZD6A&?,[3L-fYN
O/M=PZ2N\B,d:Y#edL/>\RH<>72,5YG,^U+,6FH,ZGdDL1ZY\=;_?2+D&2+0d.B0
G3JYR8d/TD2FA(_9];@FK8BdbVN\H/#e6(YY8d[Y<3GKWLEN,;WDO+E=?0=PRH+\
]98=CPPGJEEEBbXZfLGC9a(LI>)\V7:b6L;-0a_>]WZU;(ORQLLRRg,Y+=5>YWWU
RN?A-e:JMWBBHPfL(ea+XLG[Lf>;Z#9b/W]W21A)/K^\\JEJ-IAU9DW7TG-e+2>f
7W^QI=[:Xg=9&&A3I+^2T/32P#=F&,#C2JK?OaI^,EWVLdI6cQ/db#VMS<PL\dM)
ME@d46Xd6SSF_WJ1ERR_LNbLJ#_--S?A)5f-Z3IJAN5^:]e4g,TQ,dR?fAfL_FGF
JSW70gVdKAgd\RgP7G?&YM;RS9+.2_M]TPHfB@)V\YR2]D90f?[,82KOV]-[G5)^
\C2Y=8OOH^aTV(<=gY03:W;C6]U(YPTS/&@[/F@KbZe>6-S34\MISG>P3W9_SO_@
JbDMbMe^T-P.?VZB5MO?<O@b?dXI1/6?-IH)Z+RWJU1H[\7XK>OVR=GP1H6-QI^6
[HD4OQS1\.e_0-\#C.-X4=9-]e#Z3QFWQASbG.?ZeC;41EW8e77S@g7EB4g)Cc<[
<6A:c-?77W7F@48ga2:&C)[Z6OP(c..A)0/7_86?<@ANL,/eP];(O-R2N2P#69b;
-CF6H84,A01FQ+N;LMga(3GGRf1+Sf5H,f.OIS=]1S[Nb&_^@E(0/eE_-ZggHZ#E
B-9B5O8TOfI@Jg7&(&Q9MaR(UTd=H?@<gIa?XBg72UQ4XNP2aIOINU(\fS8bbId9
9P2,Z:TNUaVW:N\A&08M-X9HG6>VS_&Y3>OHR=Lf5a9(5O&aZBEd^R^MTaEZR@F,
=8DB\RR0e/WaWM-:_QZF49A+\bXLf--\E7\J4:I,M&^K_aLQ>N]e>IB,2YfL)cRS
.[MHM<NP2:8LYNZGWI.>gW<2WS.&0=E0R9QCD<:Q=Q0.c0c+eQ.cF[>JT2FWdV\;
+G3O,>ES&E+\S#+3DA;\[4\>>D[#_.Egc#T=4Q.FK&Rd&47E26Ug0D[TK8bSdP;7
,)4CBG.[f#PC>5=UW>MJ3:UPe;P/.D?CNR#f+S@B=_\gJ0J0T_86DY]c]#ffF]G]
VU?WHB2&[P<U74.FFd@M>b(gP/MMV-SW-YNGDd0DVCeQJTbKHDUT#(eeYGI:]7a8
@98AJRGaeD,Id:e\BCcL75U#OKG[Y\8I^:]JE5T2@bB#>DHRRO-adP);;PgI55]8
gXQKGM_ZY&8EgX6,Y1GA&V524e,.PR=#cSg8=@K2)IE\_cUBC[[JD+bcVWCU-(a8
8]P(XI;?O^gCIabQ4M=]Y-P4XJV-43?WYfM/QNMZf,;Y>aRC5(VR-OdML(,5KKc<
;XV4=b0Hb7^NL2F5[c;,N]M9[FRUCNRAg&J6S-B0S]fa,Zeg0N0:CFHO3K3eU;d#
ObPO>SPg:\0T.SET<#+g0L;0]\HT8/g(F<VMA-5gV]N#AHOg2QSMd54+N[V(1E[>
8]3REZG=,Q=Wc<g__P<b,_FIPOXbaUc4CQ+H9QETN^T9G1,eg2.BU\;1\GZU),g+
BG5JZF-[cQNM(fQ@]OOBK)>+5(.Y(]5cXSI&NfadaW6LWX_Y@_2HAS7NGF?H4L7&
f0HF&1AD^GK>dVN)NV_/[66=;C=4Y1,T;9U[L66b8B+[RX]<Y:e0YLCgf[59I01^
)JPGc7NcGKE=I;c8XW]LdO@X3d6UaD/[^QbE]M,C(\H_NK6(]IIGW:O6]VIOKcGG
X;eVd>5B?63?W3-0O,0M;2AT)C;69@S_eJS28/Y<9PW\:bcL@QT5;)WU@gCNVL_g
bS+0KR?^=W>G6Z9fUJ1UDgaUFF6^,/gYA;cUN/fAY4R-ZRLcUYf@]-;2CGEBe3&8
/PHW=7,B.>@-7AVN2Oe4>P?5&Y&8W^:,QedH<CN7X_M.L#\ZA[HZ[E0eD>FB5f26
L7K8M9g=](U(SUNJ9fO5=AO^?cQ,Y[]\f]f+\C>)X.Qd6=A?QH#ATWAZSKG,=R/N
;TBUWaZ4#5+2\TTEGR4;OO&GQ(:.9Y[)7;\-aC;\H\eCR6f1-^Ge46QfA2QQUBa:
(N\fX1_eB6fT#)]C&SUZ.4\(UYN-\9:1_:IP>e4?ZW6)UDM[Z8GcV-1@3-E@B\QA
3H<G5>&7Q<SOe=SN=JUF]/(HDfE.D6e\EV.#15/FgOMOaD?bM])+MB<K7,#Q,JH6
(6J499/?K])KB4=\#5eKQ(B9B@6IXVaD4AD]:0-fBfRA2ZIOSe(<.eD2GY5QU=1N
#G\ET0fW_BM7YO[UdS:d.,gIPBLU?727Ma2B^5]:[A@,74)>+#e\W<V;JA4:aS]R
?/e-8\DCCA4G@YXJ:E6L]#9M,:&\0Og(KW-?89I+f[,dZ20&Q.]G(U1KE[F1GcIE
O=e/TK/bW[d)#(5JILCeSeH;&T>C347.++X+3^FJPQJ=GFCID4H(O<Lfc;QU&3]C
@M23&PYTY.AeC[+aTW@(fDa#Nf-;\)[K)a=&0OJG_.L<MC,gA\]0+]&B[+ON>LL1
U562R<396<M].H89F\MU,68cB3^)K,B@BUUMH?AbcNY27+EVZ2,WPO2;03ZZ<gH3
=[B]eSa@HYM>G,d.^,bQ@THI.H8-K.R,gGQf^&/0f/>EGS@)c0f;Ca3+2K5-J<;/
dGCHePE/ZR2IU:]Q9U;>9RG,O/+1-6+STCDNB87<a7RC6&eI1,AUA<V\ZbUbS&F/
RVCLNSBV1GaFb0S_e9?ag>W;C;#BMacG/G)TeBEF4^Bd;)JVUX)=XZCe57-aTa3Y
H>?cREc5?Z8+e]Q_WgNL:]]VQN&262J\:LFg[)g+Z(0Z7NK;?^6+[a;C/QJDQO1g
d2,C5)\?g72D1P@CW0f-LG-[9]K?5OY^5/GeG,d>QL2Xd0DX3OGc6b(fWa-&OY2;
HK&6dc2]Q[8?Q38JB6S[c+fgOfaX0/T0)F.&+M.UWM1P1H1V;\3I##f,Fc><g9Ge
+]NZEEJ[g,86E34W0RV,7>?Xc\4f/)8O^.#,HG]HK2NZ02QW]af+.QBb^3WO&YN0
)RDBc@,_WPEYQLI.1F;+=0P97(^F(6Y3L+QU7bfgRBf-/Yb,AR<UCCBL;H_42#bI
[K>YE_D.S-DX+H_A8OgPP9/NFe&0&/]G3C@3@]R+&KgOFg(M#]SLC+f>[9<dWfC5
OMRZI5[C4\68D?[81@(O?d]=XJ)g]GOPOU2XI/:[N_8:RUbb^2A#8fR62cQB080T
e-@I:>II9JBKO;TQ1Z7?>[H3J4STCc6N,f@0YU<V8UX\3?SAO6&-&_;&FHOa9X_D
\BUJ5e[>C^+L;&3N\)E-])Gc:A+)H:N[O-/FFacg?D19)XL1IR]8C5BW3[F0b#L<
V>AK103Ef:9@8(O3gf4/AF7#YELVaXOFL33abBBI1D],;;@+bdZ^)f/^B<(.R24F
H:M8JM5D?+#63M_g^3@DBGV1HKcA6<99:+<-9PX8)?ZX8+M:PJf^XZOG@DU(22QX
5e=e]bK[=IgKd1:60IJLd/a+F5Ub=IPX_PA:D(91cHR;0M/3_(L5/28CCAfVRUMD
M?Z5OYHWU[CfHN#W[eA]MX;O72_R5W@HHEZOc+OARV[TNa=d@D7Ed:L9BZ?5dgQb
O7NGV<_:SD&#IOYTOFXX2)Ne1B?gKd0e>L[gWM098?GN<=FLQ7D-;O-+a@(,N/H9
_cZY\G8\Q&0&T<f4_BK05&-daQfEQ=1W>4#>]LX-3K4]c7KX(_7BPG;7(RY[2YaJ
I,]dgBDKc)7Q?2[:gaF2c8&@LX(\&a.eHJ0A.8<<3XXgQ&b\]d:2O99?N06YH9UL
[>08dPSaSU@)Q]e</N4e#>eKNcEV+PaRQWW:^KXfFW4^?QX2)b/^3@>P5((_4WQ:
41g.?##Z[12WFfeAS4P4#R>M]_;W7:B[C77^U;g^_XX0c>ANf)OO[O]O-5KV/<Z-
=b1Ed+/Db8f_/0H_NQ6-_JbbB#MW&>KAWYf2T058P0f@1Fc4/D_/VBdOBOJ)a0&=
NTJd+T\W\>aZeR2+C0W?[#\N#])A^c5+2f77T9Y=I1\K?HG3IHC4&=Z/R7(9E=Ga
K8U206NG9(Vf8D=>3L#R_/X0)<_A1a,P47UeTP#PBc]=I</2LcV&cQ/@Q7HK8c.6
Ke=d\:4G<cSJ5BE(1dUba>B-@e?V5_A^>5TTKNVJe,/TT7+4Tb)gAR40]Pe^K3@B
-Lf>@WgE8cA8U_[Y@O4E<3c_M[-,cCXGOYLcA^1HfX/V6[fISSMZCe_Y3?Q<UX[4
)B#]GK]b^]3F6ZYC7Y(?L,5-9E\)aSWLZP=7d?P&3?JBUNW@7;4M1E>@8C\YGff2
#18KG&eZU\E1Z7gCH7?/\SWVXI=9ZE#0V@V,B#6&7Bc&E@-9ZOG(1X0M1([>#U<N
HY9H?78EGUVV^c33P11[21O6&93VBL\B]NP4I#5M+3)B,IeL+9LE=S\T>N(BOTET
,])?65V<).JBA#-.61M4Ma-bST2f#;8HRV0-/?9EK(OUX;JNE=4.cTBgYL;,@ELJ
-Q4^<f.513d?LUW;7<f/#9M[XHA8P2dNT:UL(>CbMcQf^5X@,bTDQG6.=7P5AU8)
O0(K-Z;#.9#_>JPd/X2D?_]9Z(Q=A[(>4?7ScU0UJPI31ABJ040V=cX=c4O^NJ?3
=If&03f25S@4KP/XOE?cZ48Z80_I4(\@8)9PL;7M9#[TTBP_.1BI[agKH,=]VD78
cGZ;V&_>Yg=?TO-,g;P4e404V=_YQR+:_1JF^>:)(O@-9QK:RJdc\b3?M^Z1:UJf
1Yg1B[.FG4>\OL#5/4/YA-TZYX3d+9+K)gdb@9L&S3G+=H/AWeZ&SO-)c90X6A\(
@N5QD:c.QD<XYUIgDVX\MQQ@+&QOW?@BU0URM.,JQ8?L_Yf/eG[,?YGTU40F,/8E
cGL]E^e7)B\SDCM_S^ZPJ(HVY3eTH/7&<?8LAEP40[ZI_EM2;:WF\60_0f#g:79b
UbYQFJf_<(S[Zf@)(BG16KV(95BS:_c8G69^&LR:=<B:YcT\CgTQM^d,IA9.]EHO
ERH0NV)9=W=#J)Y:(R6Ee3AJR9V@KdS6Z+GADH&Y[aRTJR^X&G7P..@?UCRJXPdb
IZH]<:E4H#R3cJ?1P10+4VD]?ZT#--TJJcH+8WNbGUV4T4+60?3P&->=V5^0O.;=
<e5d_d<0gDW11T?0NZDMORN,#51RF+3A58+YB>SLA,H),SZAcaK]Q+,&Q[/3<W.d
O>AF2,)V0WNaF\0-c?,+WRcQNOH>-&II=a\.+A4=V>WZdC^6CHQB)XU_D^W.b2Q+
4G08>L^KAYaJ<9d=:XKXaF,<C@D/2cP2EA@O-3C]YGXO^7/T4^>685-,\>b],AM[
>Z8^fSaCSSFR/&PPMa82^7ZRSb/O)]);YK?FgQS18dDe1KF:^^Y#1A(>RL7]P0Ze
c@Qd\cQE?dQN+D,<:+E>Gb5f-c_T)_NGIF=Ve(L&QU@+Q4Sbf9YFB^A=LCSC?KIM
?TZE/[XR)eW(WI/N:7YQ>#gROaGdc7/)X=b(^D:IXde>0MZS@b+PJHRRa<2\##a3
C&WNR<68<CPd:([2F[WC.3\Qd^Q5ERV.-0_KSTE[6dA@RQ\f3G6LfEOf[:ZX<C]_
0DH(E,4K&40MLE9FXe]=PG4bB6IP]&dO1H@>+9]5fc@_2@LW(P412^Ea1+]B)eLZ
8a#cYZLf>YG[7^7@P]G:(PF;OA+1_LN2?JPeP>F1A[86?.Gdd,_J23>8Wbg?e?gF
.:D]f(3\2gg;Z#4bCW1-+DO=dKa>4,=K#e9>A[S.#)3(55dTAE2^]#JdB#>P9a<#
:N:_^gSX>A_#)adYI?];EdNUIZd6MK<H[MNa11a4b:(CAB:NIL>IUMV3XR.[:^,&
LO._X:S6T4/XNed=\Y67d\K-2@10LB2?\1c#G.G7(Z-f/S;5FSH<;_=[gS;[^@Y9
Q4[REFAZP8[UO:Wgbb?7N&XK8L@SAP&:]E]HR]?;NLd.6gQ,OJ.&8650U167>_;;
bZg#YNaD.<--[E]gU=1BBZbH_?B+O40PU;>f_H:^N_cN9Q)g17BWTG@(824XQXE4
4&OKB<V3D8^30Hb.N/a?(VcG\=g52KC@2D0(V6RHfH4>F9dBX6JIF8[#5#=f7F1N
6E&-Ve,cgg^c0,GF3Sg;Nc9(ASHRc5-f.+SW0?VTTUae?>&YZ+^04+?IUc-41\,0
?gAY2+KH5Qf7(aMAM;5)[3R8.XP:@@9eE(P#JYcR6R-I@QWaT[QfS^99>;^8[B_\
Q5L@W@PcQb[P]M\DXY(BZ.M-@GYL5@aRG,a1dDe:=FHD3cY:79JeY8FX@65#E3(4
GW9>ST@N;.4:UYKN@B-FA_J>e_@-Y+/50]4]:TH,1RaRE(/(M/UX3fAVPa_3FT,J
?LeVY>d-Ed;^+0YHQ9a,cT3I3b7>g7IWXP3IUec8G;6=dXKUH8@S8GCDeJGMJZHc
eTaA@Ye(F6,70^e+=E+:cCg0?5MbgL_CRCI[BM)JIQ]2A0\/3bH;=eO?.[WgL,eA
bR2,=&66.6Q@I(E8-bDaKF45NEZZaG=VG4,._@dBP7<;:32TQaM^AX6FDG2V@H9g
27a8FQaYS2=I^ODfHO=5V:OREZ]JVECQ6FR#d^ec<#OZC86+\D+[V;JEb.#[#\E6
-C]W:19N7PPK:g@4#K_M2c540U,Y9HRW(K;,L.EHg\D[@8/=;f#6-S-TeG:&M<g;
BfQAFD;G=H9f_<,X?2M[ZUUMdR?>fG<DF)0<ag-8F0bFc@:H;]Bc#S=/Q22e>EeI
8Ld6g=FDM27e<=NP:4H(UNR8R(I6bU08)ZGaBT(JL\VAU<K58KPVDMO&/Y1<\A_8
64RQI\36[L[]]#aGPLe(gYgXP?AfMUf^67:IS4?e\2eU/f<_g8DP0PfPH#/]H;Df
^NNZ<g+A8ZKAa:eUJ)6@bWVOFe?Z4#P-Z(?>.M21-3?85d8e4Y+R<F-T]Z]OIdX3
-PS:@8&Fc]P&\??/+,0b4ScAEUI(06<YVVOJH8__7TC)#.A,/Y3Z(5YY-ZBT+\3[
,bE4F^9/A62R&IN8dC,+.L&2Obe2&b[KOdERG2O>B0D<Q712:MPO/PQBe(8R5(_@
\VFbc6@0DJVM&]/.gI5O5@W8[]C(@]Agff,OQ3YPJ(ZgS)(AR0&aN#\0dW_=[A&5
W=W^(HF1RG)2\e([XJ0344&L[;^V2KF1U]H)=MDV(LbT+;#:SV;&:fMT,M@#f4SF
.>(7;a_&3CB<HeB4T18WL51J^.QFW.ac,T0KLbG#9C^3.d;?Y[Y12FL\JZ^O27#:
BA+Ra,#0D3e+((I#:K)7LgQb/VZG6Sb08MAX-Ta[g=HYX9EMG#bI@<T5Ta0?,G4\
1bN(b^8>b-c99=V#=7H_:gaf]60e=[GV@N406HaUU5#9(<0J/@HE.XJa4+cWR.4.
DY;a@Ld?=_(^g>7GX#GG?7MRL/+4I4L-<,MYf3<ZS.f.R.&KA::1IH5RL)A?CAF2
@Rf8X<3SOBJ;3II+L:D=P-]N.,CH/WJ)_4H.?^2KA&_abDdSKCU]P<])gJ0b-FE(
ebg69Z[gJ5=2\.)_4X6+M5CD>7F8dSd>ac&58-YXLPJ]U]TXO[+Dg4g4=_abS_.^
DZ68IC<[&^9ID])E9,c0,fU9NF-F@e(H.:+&;fWg8IW3Z.T)>;LJ8f53GQbdTFX^
O2QAEO>VO=;#Y>JC.f#(;D;]:F0SPX8G7Ud9M.#XB=2fTDaN+G<RgUDR(R80#\02
TDQ^b0=E1^eT06cf\HOTa(PW7d?_(+(9HJOaeZ<M7VIbZ,&bKH&A0Eg&<\8GD2Ug
#NK4>QB@^g+(GOTBQ(=g:JI^KH@&(X)/e50f=f=OGPcBWC0@93T0=8RD@[7bOCV9
:\F^d+M4OD/B72NKIbYF5/]VW#Lde#(LL+4LA(4(:]^Bf\)fab8VC]cH967XWB,a
6N#-ZH]M,ONc=ZCQ@.4T=A\C6+NB@LIb[4<L6OQ3+@DHGLfRVb^FTZdJIK)2O3NY
9fV@I7^S)C(&2M.8=cO7NeD/g,UC.b[6HbYJ7&8\M(>E2;&Z1f1,3bTY_1GVMf9a
:V))DB1;41eT6R2;UCS?P3MR/c@.7]BRSCE@VGTJEf\4:]Yf>6ZOb:Y5:VUbWC8S
UF(+()?<V888P)T7^2YF_U[:B8)\GHL3g/H5EW&XbeCd[>H6^ZXUTAdP]XDHSPc@
-J.fI[><8EQ+#bXNLdA6]O#DZTgA_4T,G[LLN5WB0G2X_GW:10#cbA/&;&(b4P#e
1N/RQ@NY)c/7Y>92.^,@<]I&P061Z]E7C&IG>)@FdSO?XCe4gXVYJ:,I0[&XLf7?
[Ca1:?(IJC;Q5^/>6XKI@Y/@ga(8b\3QIE(_2R5]AOSZD(4(G@0DaEe+-HaVc:K3
b1Z#_:3.IU1d[a(eeJ=aNIA213:-@,f)CF3J[cT[cJMNN)NPdH0.IKOH8>+RddPX
JK4(gDTE=C7#e>E)S=N:bPGW_._ROgH9^XLYd>1DH.^aJXWgL2Z:+N:L4d6V]8?>
-ec5]EP<H394\g-6R(K+J@C(C^0G&[1@^+PO14>M9KL;0&J.FU<E]R>,aG_G=_)R
=I5Ia::b=F>fK/(1D?\<Y//<6J?L>gK2e/)ba<J0VUT2c:f0;(_2&#E&9A_B+F#B
S4U,+,]JQgK95+Z\K0P80f0FZ)U_0:b=#5FXYbVAD(SN4+TceKSL3bBcZ\+d7eU=
&Y9#?X/.>@=;cYg1#<35c\<cR)ITCT1R84<R5=dTUKA_#ebTDI5?0L2_BG125QXF
D-ca@3Q66Sd&Q(E5VBRYO@f+_^E53-/e+5fg;]#<+-1QI+=9cZVT8B8-#e+7UB=W
SQJbX;1CZ1]WYdN+K83KG-&)AT=ZJ0EF1)Sg,4@4^?B+[KfV>YK[G:M\d?:CNU4C
)T-90Y(8ZZ620I4EE1M<+]V+gU]H<X6d\GF8X;[\,-09>T.c?Y2M,Za^aeFPJP_W
;d#e[&&++_(\,R##&FJb#PB/9//40:U^N2-JU).NS(e&&^6/PR^VYF55GG.//D3E
&E\7Y-WfL1:dPd:aXL4EW&2POKS;Z7S<Ydd([M>#gH.gU1CFRE&Lb(P0L;[ZVWO,
Mf2D6C<=;Y2HNM=XbCCcL9@7CaEb8c&#>M.GSI2fc93=^V6U(0A;:J/9#3ZfH>5B
@V,B7Z6AQ;=D&GZ@)d-Z1RHURfUJMYdYJH>HC&Ua1/bW]9YMB7d2^6.U<L5M+ZD\
^TR:&>IV6Q(,=M^[F/12c?9agA7@P,0DP+AcFV/cZQ^MQ\=K2U2K-;3#W>DJ,AQF
PMG^R?Y=aPYPJQRd_dQ6?4++E>O4GY;WKaUOgRASHRU9NIC7IKZY(\a<DZ)O(^>O
G)g./YDPUDP\[+4JV2V[<8f#53ZU4MV]]a/\GM_bMH.4D<EcI@AcZCJY<:IO?TAc
(OIVKGQ3#QW#f2EZTXf,G>2=ZFcX&(<EQgVJeZLDXa,NIMLeKWZW?;5Hd+PY&Z_d
,A]R<&W.,S]I?>67cf4CZG/@75Z7M]J/G\_84]P][-5[WUGL.e@b@c+8B.Xd8BPL
INX82\#g+3])I>T)BG\6g^\;SDT+O6g;8QDO0JfBOL9.,e^N@/]0G9LJT,P(H](g
Q[MLW7XN9X-Ef7>ZHe1O9QGf-<&a8W9X)Y,MIZO+7.-/J(-0Z-9X)QATK&fN85#5
fIF+Vd@<,U+J>Y]WZ7T/W7(NC8@>D>AZC(HD6M:@-.[Q#fMLI7&JeY,#D_I:,IF@
NC7<Q\>aF_M\4ZA;/?Y9H:/3(5b>)Ye1-EDWgRJ(e,C0)UNgfUcL^G4)2/?B<aWa
HS6=gHW=EUV2V5T[(06DL[<;G0g0Y9+;35L8T_/+BICD)PMDR\=c6Zb0gHQJc_M@
3d\O>?JFQTJQZbF7NG:3K7f=2Y\;P4,NSKdJN.PeE;e;T;;eC;3NaD@<O125C[bL
O;c/65_8I/PXEHIU8Se36=@Y=\Kd=AG8V7.QB9LgH?bF,Rb^T,=9A0A9B75PZ+O>
(e(_I^gS->N]Wdf4C0dOR5PWGPO;9O7KJU(\@4abCe9>H6+5)D_DE6?VB64MR^;D
IaX(I0b4\;7@,ZI,S6IIU7&DO8C101aa<NJFITHW[331)7:8/\8QSX0KdB06);_K
1(K2,C1P[IEO7>((D#X5<DUZ,NPVR5565FG;dQW,K(K2ANc-&<U^02-&+efXeJU^
7T5D2(8+KE9BbDaCXIS_EX4-bMH&SO1-3I]Lf9]IGF+dY7DQ-ZWUT,I<:Qd(G]K6
MKJ6a;(R9OLT_)Tff;IVCW^E_<BZ>c_3NN\DDMfWW7MYaNO)&1P+]Z9@A51,]W1f
SVCe2^.,d]8_M<F7eMEJ7aPU-NYagJXK>gK0BXdA3YNg4U-BX?a?88<MPB)QDK,Z
g\:3PHa<XK0geRF[M2/O<@7<+2+#7CeD-;D3C3OK]g)daHYL0CQ4&(D>)#?e>9)8
-[g>I.@4,eW&OK6.EU9<2HVWB7E/7,XNX4dcKL(O0?<+Z6&X_YTR1B537(f[/#)9
/71f3GE&8CJ,;XFG5M[S6D=94T6^LgSK1=3^;I94B7+,GUED^V<I;3BG:4GKd1/L
]1I>3gIg53(Web7.G/DWR-2TX_/C^27b[L;&1EAQGD\QNBOcG2[g49.bQPU=N\PF
69ZU1IaL[?VKbF-]9HT:#-<VeH0XR0Ff0#S0VT^-W;,E+:Gg&@35M0NLJ?PXCJ\6
-(?VB#[@QM/B08F5a6NN)+E.FM.\@=H?C0#AGWV;[@AQY2@RDc[6eV,V-6L:OGcQ
4PED\]G09Z@WB1eX^S\f8ea+eBFT#WY902ZZT:&VHYGU;11a29D>A_=CIFdE4+V\
fEUMN6<U]6/AUd5b;+P0(62efR9EW?[L8L<e:K,/SXF-/Y3<fTcH1;1c0[)FIT85
TC/T0>D,)YNFXZc<+\[EECU^-ADXL1C(Ta@T[_XUa=F06;689&bP\_0b2U&aC0GG
\g(2f]PQS8=2ZETW,DX[ZI_HK=UcYU583/W&4f&?f)@:9S\G/P]#<\GG+cUL-&S_
cN,RLG6KKQ.Q>(+a+d<,.Bf>\5:(+aE.S#Wcc<11&WHJJBOHdFX1I-)#)>&.;A_6
BCIW.ZgOY5Z3ICdYag3NeaO?(-?LJU[DJLJ]H8^/WT:E[VL@\[X?:124#^H/JQ6F
F\8;@#S^\]B0+IB-?(QC=+>eJ8GYDccSZ@Z\KQ=\DJNMVS9W))8=O@PO+]K[O.R\
I_P.PU6ffVN+O/J8B(F:dI?+XX/R416BEF\0?D->)G&g=ND0fQ[1)OLf8LII[#[&
7gQEC7&EcX74Ob)C4BJ<f:b6I[B1_71P41L&CLYQ.F/XRG-)\N=C><M^<@Q9?(+[
58&8P_e/8:OV@U_@@X:N1c3D/Vd(9&#]-/SP4_&^#W>;SE9[22TT^+KQfF@T?#^W
=;V/b(+<@7c9^2YZ(EdCYOJGW(N?F4F/+APdF1U=M/\>#Qa\QDQUV7?R.6(Y?HUR
^cebb)X@UV[-/f3aV\HSU0&:a;-L+(#DWR+0bVBN^QOYFdC:F]3DU7NcYV6X0U34
\_U?0WSI;A]PD\6=@8=WK;3\0;d4/IJN,(SEg>c@)P8M#G3HQOHMHYV4>/>978J4
2KgE<aI9@FV<64^X/YO(D3[-GO5b7X#@IPVQcP(M&5;+_H#&d1VI/5L84>_Wde@d
GIPLEHQ7_0&4LUQBeKPb]<=fYMK=39+ePB1G9a9HV9KM,J-6:.S8=CZPZaYSRMff
KJcC86;W2Z;#PXA>.J@Cdg&-9eK=/ORNgD1+0,21OVAW8@H3Y>^X#,\1]V^\[gc^
[ZbWIHg1F@0d#Y-6DU()5>7>8MB:D;71G115^ZUE3DL\a.67IH+aCH><PKgL3?af
1a>0YBf7QS,N(PdAc>8^Z3cQ9SJ(R4TW+G(\K;QW5<_:5@=CGUf^?g2SD0@_F@Jd
7f+XC^U:G_RN]ZYEC:_S9M_B/<,K]</[Le]&aY?7K3EaLDC,F>Q0B=g7X>4eD(5W
+;Jd4NH,RZTI-^X(eD^3]6gYW,1dI@8?GW1[5]&V5a+8=+(ZAgAVI+.L&Ba)F<9Y
VBEbgZ9N]IOgF4&B2RJ:_4[OES3g=]d)4aPI^K3N+\.77ZN3Ta@2J.EUG;QDHDWO
4B(&d<^-=SCU/&>8X]QLffb8VCC+LHKW9KeW+8@X,GLM\1<SBfGe?DP]:I\8AeYY
1NET\Bc39K#R[M:cM.dY+N\@LaRfg+J7;P1VMa#9;VS:A0AOfH)Y[YWd/,9:@#d;
OSB9@bF=)bW5\;N#/[C?\+4-a^?].cF8LKA2_e)7B+.=Ib5I61>6>JJ6Q[[7e\.J
,,5YT/W4E4T?P,V),L^8=PU?g.=JPXQK@((a2?Y8_@IT0(@fFJ9,BY5L7dTSdKXT
6R#]P1.]Sb1BdIS?LAY8(Y_\6db=+[.#(e<+d?&63QgM?OB0I<B<aP7(=_KXBYRZ
.>H:R7Y>MM5R/X&1(@@PV0B-80YKcgab#KIYQ]E3e&KRJL]JQ4BObH/aT007B6EQ
dW[3UKA]N?:cK:TC#e#[?L@a(FC;cL6BBP,,]<&28J)@Y9a-=R1P[([[^AQ5J/O1
PE+32AK.HBdV.^M7).gI,.:G.UMEf#B,7B:.CYJK&-G]GAJ>A#P(DZ@L531)JVIT
da>ONBJU-g]^(#_T.&D,2-&#(G7_UMQ+5,g@#g2REFB5TAECIeSFJ:I]5e9bAeG-
C#g#UHM>-ZAILK,<CO@R;K7BU2<,Lec4-.=D_6?J6:6WdOE>4&ESJQR@V:9@0:2D
:#.16,#+IQ;77_=0]3:+FS/f?Xb4M>_UG1Y<;U+B#Z/HD<6W<<RAKC\KN(=eYB.U
YSV[Te5NXCFMI]9RAPX&AIXHSMJLePcSdR]M/D_X\c-]3RIYZ2dH.4NJD.KOE9)d
ILSU9.a:<N#7#V9QO6VR8SWf?F<3d=(LLU?Y#X/H98O,L8TV/Ma[;BWTNQe-ZeWH
UbX1I/2AWL8-E:OUeG<aXf.2D(B;0:6XIb_V:^2L#O5eM2Z)VG?@6SH^T-1-6,aM
[MV^(^I8,+QJ(;/dT7CWJRbTY-C3L[XXS0fB+[-DS6@a:Z?1b37GcN^YQ\.3Y]CE
V9+(\H]84UW<&4.f&e+S8/;&M,PSY,>bQ+[,/F+D_+M)Y3;CCX-Zg#QbUIYg/0#;
;HP4-HOLMID=;2DK-MI9J.H3_<O63MG.HEc8_,?aU#HWV?5H-Cg94W.f^]C>B]U>
Z\34;,0@K--C38^KgS9#+4fUP6bEJ?/ZBQ]0O];\;LGee[\.04f\5BK)IBZK#7DX
NCA:N-cEO>Xa>::H?c(d4++QY[)TH=bX1G??/608(ULJ[8)9LBgPgPHKT7&;3XJR
aa>;HN-]52LS2H<SSFL,_8QRBA-V<SH56c,Gc.^=6-53Jd]5H02eZVF-WLN3IX07
X33AP6.[69.5Ic,>1VM4Y@GT3Xfg?=2LZa[BSafBBFL<^7NNN):1g+4Y=GH682XV
U2/Ggb/W;/DAG+)1I#5H(#3+Pc]PT(bQ:J(a<B,\G/7:1I([6))2QI+<@VcFI(9?
?Sc0FO9FVSU:>O<,5(cJSFD[;Jf7_P2#?-e_=b._7/@a[1Vd@:9[.>]<;e7a-_?H
:V\>]@)EYB9VZR[?DLd<SeO@E^bJf?cJ5;5P]/-DW+ZR=g&<Q^)ZJQUFS7eBRNNf
X\06B6C?C+=fH+W5LX5KaJB6?HT6XQ>:2c^<;BCb</N.DJPZ0NNJ&0fZFB4gagc2
WD&+]WXC:K/c/^NNd9ga7Y+[9_[MgU24JR(\:[E(gXSJ--NKeDBEDBK:U(A&/+^T
eb^P0J0P5fHR5N_DY,\cY123Mf5&ZN/0[DX;PA#KWZ:M7M_P1LTJERCWP/<gVG)#
)Tf<O0YYVN5e-DI^O,aeH^4&78#6_ARgTW9Cbc]NJ7#g8;WC(W@g>UTg)@^]UIZ/
[BW]QMcA1Q@6G5DK[Y:YY@Z,7Of5/<f7dUJZQ+63-YC=B34WMM7,)Z2FK0DTBb5g
NL?3e].BF\T6Q8H[ga&PS/QK1?&FSY.\9aQNI1MbMQWTI<9(0edGQ4ACPP&:D?M4
DE9?UA:((<C73E62O2g)6K^BYCAWB-e)LARK,/3JUF_U#:7&U+H4JM8]0HSM#<RT
C-<>cS;EI7K[NZDef-OD=CVVaJ30(L,5[fd<_Med-Y^KA5P\b[C\]I:bbZ-N,AJb
_SA-QUd+_EO<Y7Q7(65SO=,(C.Q1-Mf>:G,]MecJH_C@6&GNRMEFVF@@\UK.IS\P
g5@RK?TCF<QIBGU4TAbF8+dQ]@#3^YOMfg\SYJ&<L/NK/-4-)8OCG6f@OCA5)PRJ
8H.gWCg5eQeeQ:?ZE0PNR_\4MD(BVO/FMUL(V#Z8+A0a=-[_=JgH;CE4?.VYV(CU
TgN_1]g+2;e2_LY=XdeM?-PNFEP20==CP]M9+DFF-UNBP_U+cYfP?7dE,(6<cV#5
F(SJFgR,OLR444I,WaUJ[O\eVK:Oe[N@a)GU0?5SFO+/b?Dd2;#6,Gf57H,=7G^X
<?=JPc__L@NVR/1?4NUH+,53;3Ud3K,0C2X4^^QF@gS<,8+5b?,758&bU,=&d0R;
.?]#XXK^e?Pb\dSI3:+694fc#P#<3DUC:eU=1<fD@XIVAYVCBg(XAe,,M0S3X+.g
AL^+KN>H]4I;e.A-Hc(Ja)\13VO)P.XU?F.PLEB4AW6d44.cNHXM#7MbfZ?^5M<g
I>gZ8YZfP+@1&gc8c/.M:)cbTC]H=J/Bf7bYe7R\@LX_Ud#6XSXA2VKRf0H>#0f0
#<84a=?c;<S?I9:C_7fEc6GKOH5KK4H<0:,1Z04G)T<O)-Ub7gZO:L)UX-fd?ff2
IRLSVT7H,g<Y3@A&S01-K7(6M/dZM\,ZWbfGOJWa<<gK5F:E5>U#aP+^/L&O=eKc
]GGaWP,?EHNZC)Z0X/-4@/8LLI>T^?;EJ.CYQGQ=1D8)Ge6J0F@cbd6J5;,5K#AC
D5fGb5WJ)H3P/cV8:FdWEG_e,]F61R5X>7f)a6A8IK[-7We7=<+f80/+-RV&7L39
R9:GQB8735B^7=^5Ub<_Q#Z?Q-.YW/B+2+9Xc3Z-SNC1ceSbI<_7@0)TFKI:7JO[
T;cUH#af4A:5Z:X2+D#22C\:Y7/K56/d=N\P.2?3\S&=K[[9Y^1MS/L\O&1;a/N<
:K+>OK[()9_<(?(YM_4Y1\X?>fN8GMB67BS6DHV#cZ;4B;+^fD?=BX1HZRb/OK?1
:I#4Ad/gd]b?&JGGZLOJ6BXa&fOM>#Yf)OS&\U1D-^3[[A1_RKX?83;NK?O-?.]R
81?KOg/@Q6YY_G8-[J5OL>@3a@/-/LVCg.6+d]V5=3ZX.B3eP9HgeTEK>d8SRZ]O
34^3H1eg07ZN/?B(Q#eMIJ6[1?YKcG[)C-_D3VJ(74e=VWbVd:?4dAC<GD[4OU]e
C,;/cY&(>+W#N72fLZ.:9/G?8Tgdg?CY.H.g12VZ\&_8XGdVUZ?VHPP0/)>8@,[a
M;/2VK+-d3\dYQVe3H-N-8a75_V=eS.(I>GgI3#@L[Xc:K<[1TE:W[U.[^\;NNH0
2T\fc-@/U\\9c/>U4TO<>gQ.GX,&Z-?2BgVJ-=.=A.b\\=.#Sb1DeQN7b>/T3IOO
PT+B+VH_a]QR11.41ed&<(AZQaRKRS=QIOL,HX/@Y1.Jd2_L@;8ATb-TW\CD>^9+
-IF@9S0\D7K1H00D6d.DbffM]7MUL](N1DCP,9BD^Z]?8.SV1W<MWOBNUf]cILR+
S:)YH>fXVX)U/@<ee-T-.1BX3I(\.=LE[Vceb:_aRD<4LGMA4L6[S^B+:A2c=WK)
VB5UfYIBLCLQEH75>eZU@dTVLIQH3K>=TU8bJ:0TQ7CKZOPJ<29EDfKVVG,NNXdG
BZJ;2I4E98N,5E9P^9#B@Tc1g4Z<C5J324TbdMAFG7.<03#]A<[0Q#g6&K9dYa(8
G,^ZS#T=OU:-/N5eFbeCBfB8N<TB+LRM^07<AOV]VaCIX?]cTPAS@[^OY942X8UF
Q4/_dVGI\5]V<_I<Hc0=LASX61ZH60KdAdbS1]>7b+.\3,.3@05@DDH9Me&C9P8a
VGPg<Pc57M)(5\H\Q[MX@M4NVe4[]PJT4\Z2Pg&\B\\&CTOaN.3,B35(6;8@,70]
.G.cQaAAYXL=/,3PDeW\dJOA,B8ZIC+aSK<Q=?Ja:g1NE^JMgVJ1O5R0e+TI@K@a
V#b7OW^9)X>;;aQYDKVKB8c]S]I/<f1,c>FQ&R:HWfZO)LR>M[ZFU[JO(Td-SIED
79JSETEM7dY7cDOKX:BX@FZ:/0\&K(b46e_RW670ca>Z0C7)RS]FT:O/6V,A2)[4
Yf/2V1-)7c,]P2H.^/[4A/cJe;5Egcc[Jed?QR9)<e:CY>/]@(<M5P;=(3?2d/Qg
.RL7RB@7=-YS[eA[#UL>07D>IR/2eg.(&C#RdOC9/KR..W:G3>_:B+&1HM32-SW3
ZY=YeC@)^P8.Afg)2[1HI^a<#b[D_DH9TUS1)EJ,3d3;QJRKJ@F17c:a?],TIB]>
MY8>T5#NBN&C^Q^\5+4ZDDP.X31Z43b?6+4L3?[4IE=c9VN-d:aTgER@@Y2/[QY.
0UBcS.T^6C1feSTM\/SgU4cNY#1F3SK^Zg@KUdO64YMNO2U)>TY\aXcgc0X1:VYU
B?+fIP#L>14DWKR/I=VABCVT2]?J8)2Ea6MEF70BY5ZQ3U@RO7I942QWB.3O_9BR
+Y:1D))QT7]UgPBIW:)gfU3=\V>K2a.?g,g5SEWd-DTb^0ZgBJ;3a2BI+aV(F&bL
\ce4]JB+Ud[PB?R1/bA3I^#S48M5_9?aPK-6[8/eZA9,gK(:5ABef<)ZBY-FK8\P
++_BQ<)g6.,SNUVZKRO@<)Ig,^A.068BGW+aHJ62\+-5RJ2?R)Q5?Jc7dN7a.#@F
;O[6U/7dbF8e1R51Wb[TOc;G_B;9KY-c.^D3<D7>49=YCP-T9L8W8cF1Z_89Z1ZF
69NIK:RPU_G.J?_8SLBIM1DcMf&5@>8?D#LHL,KFc@T7?JaX]^6^g=eUeQPf.OOT
:-8Wf(7N]ZN[46c.6+K>fQ]+KAGR=KV.10f\Z2,8-&L:/]FB+(eaO>ea^2_1#Sc&
5gS46ZY(9)_E>Y9:8Z)?J_dCgQVPPf1f<LQYZ5CX_(_eH5]>LX\g20bW1O@7(^7B
2</e@OWP2GW68_3PFY^=gV(R\L,K^W-BgM3&=2CdPUTRJ@Y/DDK(A6+-[g[>=&63
><4O#,0,E]RUSdZ0M6<=]N>N9_NAZLKS:4T^+>B#WaUWBI8MN30>WR,?)OA97JaS
P/:]3PO.g4E:N4;)@^T#@5HZT43I.#D?FC_[XXeXV#^f8+P9,BTTgb867Q+eR=7C
LQ?G(YPTHK=K:=deJg78CSSe^RP>f<BgQ\(;AGG<HMXV(,<SedC,.FbQN1+5MDd)
4/M?GJ2da&ZQfTC@VV-;b2fW5+ZQecZZ@GFUHS35VHUN)E#QP6WA0Kb0eC24Z\@b
f1GSPSLYT6K^HX&;b=,5=7-@=2=-CL87I1_[+E.g_c?e3e7X6G3IHUAd]WQRBY+[
^f)1IWSgOT+_=T,LXH8;F+E]b9.d&K;J\T)bS-UbSVBObD?4^afU.3.9+eHb+JCf
R=(\WHZU3[-VgVaCC=OSLXX32C7EIb(63QLQ(-(S#aa<<S0AWD/Eb1?A:SYO3R3?
^5)WA#3FJ=@G&<7)6VaKS;=e-BYKV@K:LTK#<;LS)SL8;8QL1<g]_T0BdRb&2]6X
I7eY26(Kg^>JPUBWJJ3QYHE+cN@\Y/_L?^<)HPP)7a/BU1SQD\ef97DTg@c:-;[<
<U#-L7RMGccL-XGT3,:d?Q=AH,<C4M=[NLKaO&^03PTFA2(9AA>XHCc@c:;REB;A
M#<b&&TAEFTK,T5,df:#/X^>g>93]@FdMJ?H)-cX9>KT5(Zd5KC>^#ONRF?3=PXC
J8^VU<H.6X)MRY,6\;F+JR&?5f14Y<,]VWEFFR8=a6a#?3LONfC4)3AM).D<B(:7
T[B;^25P<@a5EI=aQXPSEW^.cfbP.c<eGd7)8E?18V+IQ5c[1DD;?]9K1CFfaH,>
THEZP5DgNbU..a]S],>L(ec&5:>B-SX#6-)R&e.HGVIg_KW>EDY5JbPPLffdA6dM
gd;8Kf@Z]2HXQ(-ZB>J/D4&V)6BG783UXX?&BK?NK1S=3MLI],3d-ZS,4d1)I(G]
-COE:Sf@W[^E7:9b+-C:>)3ZLe.g6JGFAYHFHb76DU=QJ+9E^[IA>M)7cJ/,<YAW
[I&>+G4QA]H7GXFaf\&:a1D#d\.LAcGdb.BWP(M1/c6bLWU=X#2+[]<(Yb]OKFgJ
Q#Q5W92Y?2MZP_Tc)J7.,)/>bM-Q5a5cM?C4H2<&CD31@a;TJQR>.V?7_C()Z\Mg
#\B+L:gbOR8,4X2cP,aGPX0<-RNSVJ+.c/XA?<Ud]R@6BHW7S#<e\/J-.0cCY85P
CKdeK>(;.,>QF1E)_d49/9<<.N)<3CIH0?.>=GfH9SXa\<B2cR=YI823ZQCS1;Pc
>1=@::WH/\SVD1F@d;e3F;<R4>)&QTWEDc0JaT8FST<VIV1bQD)OX>)KcgC&^bPT
:XT3L<fJ?dgc4f0,FL&CJ-(XPS&Yc;D>gaTf149OZ::9NU=a+X=U+@ARV]Q8VaAe
O:[;Y<ZFU4^LbcZ_eg^[M:<8PV-]^a.P\(94UG^]6TV_M2HL0@=;Ma?]d<F<].#2
(AMIXWFLM?W;b5YCGX4a?E18<=N3)<4fa1#@WSUGE7S<e<7d>g=Y-T9+:gL5(5.3
:Ab-R+dUYY4/+4PQG<\J/)-=D8dY[C@f,/APWTTW4;2WA-cY1gRA:>#)^&eX-<Ie
W4eUeaPG8;BV^,e:X)N:bcL06G5KJR#:BL.HbD[6QAE4.1b^W@E6XP^2>BC=RFMM
_Q>d=+U2)g#b:LfFAGD0f]-L8\MU-<9?/;Tb\G1B.Wd;ZS]]ZI/N?D_CP/=A]8F\
AAPRZZSI00HX3ZJNFG@XEH[AfJdB?6[8:&?e5D4ZZP&dbQWD0E:gKJ#U5dX_SWQ2
)/S0GG#PJGJF6WN)/:VP>gI0,da&?&;0JHV_d7(87JM:A6/da:a4<HdZ)6X@+K3\
9A]8Sd2;Wb;F>2EJ33[[RVd<3?c^C,?#aYBY:(T4CeG(,Jg?YcY.,#MITZA>SIe(
J.)+eOHOWdf@PDS@^^45<I1(E019:UdQ_^T]O3HO-#3=@R7UO@0b81BGKb#R8XfG
MfeY?KWPef:R&_G&@_UW1GW?FXM.6AX[>;,.NMb^[,:0]/262TN@<:-4[?:,L.@U
:g]4M.e7RHDZ-e@1O^I[JLaSQ8QFQ:@N1bN9_RX+QHVS5O?_I8053d<6N#df_,#S
8ACD\T>_+ES175K<TS@M,f9))b>bD<&AL0^d5R-d5MDB\+NE+A-#)#X)(OUM8FVY
)0;a&WTe(TC0(Q_FMEXRCFS?@7YFWB-eaFNAQ-0;d2A(H+LD+7])X:R[cCU4F(IB
A]f.Yfcg/X0:G5Va.Uf@MHQCZ?LC4Z#+EX1PIcKZ#VY/N(\N)X,9INf&L1H2)gI3
e0JU4KY3@QB:MQ9_a[I0+Y[?M)2@JI31&g=;,I#W_)(L,FV\,)8YQfI@O;-Q;LLX
I,W<FKe&GZfI,)6O]]OE5HRGZ-8Hf)P[.K@@W,:]f]31N7&UAS=>HEI52G=d^58F
#1DZ7Kdf+:Q_]C0Cedd1/JW/PH:1)K2dS;5gSAJHSb-b\]&b8;CLFVB&(ORX.:@M
?bKX;/RB:]bg];Ce@,0UU/8B_<e-J:)GaHWGc:9^G(9CF7eCDXZbARFZ=0PJ08\)
bL\RWJIMQL42FcX=37^AWK,A.LB^K.2BV8?Z&>f/E0/E3PVJV1BS@U3I5@=J(GW[
6UZe9>TN/=_WeY-@@:<]\>C.KR&H7K;g7CY0SE&F#,10^F,]Ve6V09^QP7:Q<FUI
ZS0YT)Q,95-CY6.?,D_E9<O8S(]TVI8&6BbIPREOK:a?<,0/e2Y+V]FS/./-J:@3
T;b7gfQ/IF9&)F>;WO<Le/6,:P-41>&WCF<]d)54S6Z=22>LU.#F\EVALf0^AC9;
.-=NQNE(bI5KTD)gb&>8bI1LF\9UM8(W4?MS]S23K0QOFC<86\C>\Te>^XB+)baH
dT3e2#@LUPYA)21Gb^0P/SGdKC-FILLY;KDT@SD<d=aR27=-X@;AOM.f?bQ&(>):
>\5,YWBY\+:B.?gY:AH+\7_XV(B9S#VOF9:4W&PQY+5KG2fHLHQ_I:,f0HQG4bQc
VUURg(?7X;H6HBaBC:>5;Gb=fK4R_4=dC@+58,ZQeO>GXI.>)-McT=>BAE4+8-BN
LYc7->\e4]:8AB_gHGM65_IX<ZU#;e1@\;[2#[ddcOOV(L(:cNEbfT=<EES2UU/9
;E,0I&_9YC[R#/Xb:Zg-(e]K8TOE/QU]Z3LO/)c;b77:G:fE>/FbFC^4-&(5CO_)
N>D4?fR0P-)E21f^P)L_J5Y#,-KH44e+6.Ae@7HN07_929-UDZT7M2JBO&(b)HJf
B#,>PTN0EGTfG\4@IW\R&;T&N]\OT#BSVPTJVSN7M9.H.NB,T4/:;a9D[1(KWJCV
52_IZOY;+7cdO+X^F\cHB2gHO8IEdd+U/1\#M(eP5A,POB4S=UE5_5E#a<a(\_76
:H8aA#B#([&3=e.AL/N/IeW?UE:M>#9LD7;=0IFQ4a/6,XH6gMe82aC__X-3]DP]
Z8KWN9GT0?&T;EFY/.8Z<EM#A-(ILgD8dT9f<PO7EbQ7<gKZJZd#4I56?&NO.9/;
\d:Y9N[FNG,Y3Vg\[8O+\DJcSYeZP2BPFLAQ.7@P]C-#&78B961L&#FBWJ#&6165
0CYS0P3]1-MD)cP/_I:-<6gPV^-5CW<@]C])1O+c2LT+[:#SRQMFDOd3FT0XN5SX
JF?[;?EcNTQNMf9X41U<:AffSC.7U)L2FOVW-QG08Nd:+aO0g&]=G;OEIOHdB4V1
_H7M]UTM(LMVL:G=&C-N@RR_3JbGZKE1@S@@5XH8KM[8[RDfT59a4eOH]:fBLV@<
?4.6=]^[-=8<9LdC2I/AeSGb,LcS055N/?X9>=A7g0E#-1;I+[],Z3dV>US0Y>QE
JcIVPfI2)F0^DV7Z93[(0/YYNZJg,TO^4L19SA..RB=FC&V6OOa6<U(,TNd&GM9F
W1S1>-YI+XDD7?^4_,RM+<b0d)R<^L-_BQ9BJH/cK/c5](=+Y<+-E3bdL>,,LU8e
8K^.TXJ_,N#BX3g=3(@4Gc<H_,[9WP_6F:ZLI;@]K7MYdY8g#DE+@dW6/cUTa(aL
S5bF^bS2&>X,E]XJQ\2NID1f757/OGfH>._bdBGB&C]GJ=FIZ>NfGTRgN7DgV-^e
?YQLWABQ4T:afA#VAf^;2Q_Q+35gJ5(CdK:C&;Y+6+6Hg@(CegQXRSTD#Y@KG)aF
dZa_g5>6V8YO/(\4??FA^4<RHD3-ff8C[27]1Aa/D35CM#2?4f[C,8T@Tc?CN>8d
SOLV?#.YX?-PWK4RJB?W9.?28+g\VeVAaU?[YX)ObW;7g4V&0A?B^&>eFYP9XT_c
M&BB;<<^:ONJKR2K8db&bPZ.G+DN_b9YTWAQ/_Z7H@&Q0I:?OTS-96(<?.I[Hc3[
TI1fUO]=5.>^D-G-b2NR/E4IX=JK>ReGU&VJfKBI7P=X/(OBY3^^JCc^/U=G0O4V
N<JE,4g+=8AO(6E+^a\YTXB<64aLS&U]?2f9gR\8(c+RS(YJ.GdZGQVbF9H:YVT,
RMN3:#[21#1LMJ:>S>G)K+HR.Ye&3T:OHIFd1aS>,D;Db=#5g)@?fgYcKEM&#T5@
^H=?5<&=O(?7R1B]9K0.6]XOF_b@)>7C-OY?CCE426[^)MXGR>,RQ@O.LT3IPJ](
;d:Mg@OZO,K&3\a.;caMLO^&8;6[\0)TYO3F>O0@+S0]9GXOZ1GQ&#K#SU:DD,fM
?H?DP3KDd.&)7SQe::H8GTA0D#d;+1XB_-?a2J1#[0\@=b?f[<@.;0)?:M5ZD/#&
1&?2J#A;+<814ZL>SAeMUU+KC>VEf.YK:62]SF++=eJ(P5W\Y0MJ;YSZ#BI6QX0T
fFLFNc:V(]:\-=SZDQ-U4XI2+b19OH.#^]aY/WeDcQb@ZDX=_^H0gK@Q[6gE>O:(
&V6gSe&G30)^Y1.7Z<).f,^H,b.UB.:W_1(F@VP>2/.7#=BKX:?>#,a6cB8.3K\H
+G9&5C8;3Z.5eD6H3E9Y[B[8:RI__+46N>B:bB@&NT8).ge_/8DO-\DAU[CQ1UU.
fU<O&EgXGAba6NBbV&_TR-JcE[R5CeI6SB8M5+58fEK8WDB8JGSA-9=d2]_bG(X>
aIU&YFe9.,G[_a<SZVA#g//eV1Ea#/3WG?CHY<=^OZ,agZ=:e?9=^[RQ9I;4Q8aP
BCD16@EVBLEa61@YT,^.&0c5NSM-@<>3KcCB+V==b62bQ)e?PNM[A3U1GQM&g48#
5=N2aLWYe3G,.51>^EZW0M@5D#7[Q4.5VY4(A3I6&:D#)H6>#GSgX15XU,1<_S92
CG#FGf,)(E=<<HVL3HA98A-^VMO(8LfR0+97F4=T;e<aK79f)SU:LV<8DC0Hc+I<
ANTcKJU@CI2^K(S-BQ,SLG[?fVc\UM0<T&ZSYTW]Q79A0BD&JWdP#@.c6aS1&M\R
/DN,)60WU01V1I4D&2^PV#WUCZ6EOQYe^/]&5A,HU2H:B-I-/-JRCZ4EUET^-^O:
U@HeJW)\cM<_f;VN]WbXH;aI3c#VCWCY1C&-HGPVBeQ5S<N&NA?T-O]5D_@Lb;9X
_LH.e,.W=A2dC,Y75D(>6>^):W_I?[SFQM_ggAV2bFDV8U1OOA&I\0)A.AV_Pf^)
]@GIG4PbbfbdQC&L1,?<e#4&L+Y\]Tg)Pa_8ccOaM#@K&TX.=,.=^=-U:Y@X/2P7
bT7.#+_0f+C&R0E-;:TDC:8EA@1I<P5]L&&Z?O7R;ML8cR0dCeYNX<,:5:d4HECW
\cB^0-F@\a_LZbTdVMcM\5Y/5CSAe2MWQb5F@0L\g-LGcM@<a?(BKI?68F\fdf=>
4bM;a,&-]L5LBY\&2\NC&)JVHA67D@1BV\g\LJ#X,-MEB+YV,B5g/bZ-^6N\FMZ7
K?UOUfI01Q9Y2><g3)OI^e\VO_+YX5IKK2H5>=e70&6bS7VCHQ<<1+gFR>RVBC-&
>F^f-:L(SF\<WHEQTLEOYA;PZXS=ROGH>W+C)]UD\UcT\.9c8)c[W^[?1C)4X8<N
2f;9D0J)3(M/3049cbB@44/U,Z3V1K\EgJYW7dJ=0\21I4_ggO3@RF.)B#^@LFFf
6G6<+[1IH4.Q+Z9S)AF_;&/8WT9V=SfXUY1Zaf(f5\-ZfZPf_gY4+^cCK(GbBcZE
@=CNX42f@9aD++2d_,;P+LX;g+1gMgASNcb,&I@I3JK/D#42>HTa53_2-K1=f&IW
I>4T^HbYd,aY])QR4bT0D4;NCK(T91#DIdDNfKXGNeD>a#8PDH5\\W1aIMG\CCd-
VNd3g?26<ON-9T0;/-L))\M:<ZY3C,>;_H^>IJWMRUHB@[g3/eg-@D]LBOA?eGP#
S)\#WGW+?\I9\_>))RMMF=ROd:UV^g2FF<>:JS[V93.dgTHCB9AXcK;0>HP/a&Mb
L&M=L]E\8\G@UDCE0L+Z(NH^_,Ua9AdK0+;5[_gfRAX_4QWcbAGLagUJ+)NYGRaI
BWXaHBCUTVH3EI9fLMZA//AM\_:DZ@@N-WLZ?Q]R.dXC=I-deH@C?e/88;TN:GE)
40WA[&@#MA8?XJ]X5OUfX0+F=bUgIF8UFb33S+A]HG#SY?]QbNDR#B:WEdPa>K)O
<6dfg@K+e8fD=&,K(<<\GCNZe8.L.V132:UFWW7BLVTK6))-EM@7H#051XZPI@>+
8F0J92AU5VWO.0Y.BbCcd[g6@-/O&=)b;>NJO4_eZPK)KJ;F0_bB4.VEdSaM>VeX
#&,->:N^KP&cDGU5Qc:Z[K3[,WH,W((-;)VPSX#:@\SLLJL^gRVY@/.K0cIG=0H[
756/NI0DHP?O.NY7ZSXbLgAE39XSCAe[T>:b\EM4JH,@2feZORD;5;.d?NE#95IK
7H53\)d.c5+^]5d#AT<S75U/[O0&BK_?U(c8(CgM4T-]^#@;@247]O_XJb1WG<H?
AA1)J&R-#\;15^2Ce@7?)XT2P[gO(ME,<67:I#J?-b>\X?/65IOU1I,81O?YRI#4
WU]PPAM:MDB@J(#D^?Z,<=FHKdQ6L)2f^b]6A2gfa?I^^=VJK4NV=VYWYPd6@aHV
#.#97]d30#A81]DGPW#=Q&)Nf?@c2bNb/1.#7&1<3P/B-]cT1SIL[gcW6,[[+;K@
CQN:@\V/;M?HQ_9f06PM@J&ecTT_])\a?+gEGbW8>Q8;;,&5EdaX69:V=\2?0XU.
IR20M>Y7&c;@TJ7dRJ93c>MV1/5&H26V=[(D2Je2(V_7C-RbL<^::G)2c+-aef?K
#ZF=+2Q0UbU7Y;T#VRdP@?JF.FM^X_(K3Z11BgfKa7HE6V7IdXQ1&VHS-0=b5\U6
V&X;GNdDg:4ZN2N-#W;E36]]^6K^?M1fBTWH8&PQVPP@A24TU:F13cJ^=[fXBN,B
=,b=DXH4+e5\Ze.UT:<SO829L2;W@2,b5)8M89WV0-JYMI0EV-VT2_5+<Y]D.>PD
8/8&P,35BI2:AFNIV4-1/.[:G.U0&gCgV[CREAMJ.b.:<M,)+7G0d;DP5JUMSG.+
R:OI)f?W/745,4NOF-;_7;R=P2:dLgb/=d-),g:EfQ8\I<?4B8;QH]Z6,FGfPg(.
E6ETG/2d9+bbLAP5:?,&LCM;681dVL^&#fP_Ve?)QT]Tb/6b76;_,F3:A5209-;W
0E((->K&7c<29:(H.I(6G7P8/JVD;1O(N]Z(62=YXG@gU=g4I_/^FB@3eG.0/?Y7
ZG6_E#P#e)<Q=FI7#7U;5RK()9d/K[5;S1S/a,Y_3FLD)gL>;1F<-XL+Y>SB/KEV
Y9;NTAbGM>CNO-&94WT>\UC.79gRN<5N2?ZPaNN9B<9GUC@Cg6a1F_bccS@\1&42
9aLA;8\g>J3O1de3Ld7Y+ZW9]#5IRQ+]I21BR17M.CTHd>Y6VM[Q8[]YF[cC/M_U
+K>KTNW-Q2L-_+N(J\?MY=2MN#c/L&g<);aCAP\D9X>87_-^QRW1/G0I(&E5]W9/
(I8&7LFPUEYcd0:)KG+U;\b]VJC2-Og^<@QDW/#ZT/SA-P64F)1cd.2O.[cI2UN(
8gB+49KN0MUeJV?+2Eb;Pb200#2(70;E]dM7PD#5@Idc[P.]IHTS_-E\f-G0/_A2
PS>eb>LFb^K]0,cFD:7X,N;.<(0I1IbHT@IdYV=2-+SE7VH+>SccA@.;Z.2/((DZ
a&>0RVc6g+/=E7OdSIY0ID^dEF4A0X-5P5:),+>>&&NU\b]E3dDfC9W.WB=P5VSM
gacQH/B3AcE?(&G?YSOd2d-/Lfe5FRe9&+N[7#\V8\0M8YW>BGR;-@:&b.aT;E.5
67?B0F]&GB(D5He;Xd;L,dT&)MRFSIB9B10OBH^Z=IMU#^A-<^&<f9cM9@)^LC#H
2].AC/N+=J_SIM0:&@e//.D>&_f94(+U:QaYU9Y,P63(>AJ:3PgWNA/Og>7]0PFL
HG-/>9P>([5:V(f5\B0e>,\[8XFH6aD-:=Y8T:Db/#Q)4FeLNF#KB]3FaM582K-Q
P4Q]:K,LeQ//E-.PIRb]RYaOV_;Uf+C)7[SJV4H<V+V)7S_8aLK[MKPH:5R_]3e]
G6ZLH[U@K?H5D\1HQRUBCDZ500+HJI9S?JHW5eFVc#dRYE^:FX4F&6D\93WTG+Y+
OeBdbWed<:QdV#-f?H)Pg9e4+/Q:c+_=^ZgU/=B1NQT79a1-5KY0TQW?F0fY/Ba@
Rd<X47d)>;.EBZ&NJA0c:X:F0JgE9_G;[1()+:?8HEHT5=O7gdOXZcM&V\T#,ddf
N9;.1U+a5aUb2.(_/.e8LgP#78->->M3L\=d/TK_F0\IT]+EGPXg\W=I>QF/QfQZ
/;2B-2;X<9EaMZ?=gOW8(fJ3(QP:BZXE\-#)^;_GHRWKc:2d;YPO>S@,YUeNBR=U
.QFW;#W\X@G8.??_X[YL2X:d+^b7TKT=.NP9&/NK65DUOGKX+Mf_TIfQD>Q:6-?a
:SFBEGZ1X54EY]RU4_S-aG]][Sg^6c.]UBW#UgS6Gg9YYS&Va-(QVA(.@I,ReD>#
<]d7A^JN=dNdSDHA8KNK,EN#6.SUg[2CFKffHO/^XUcB;[Z2C8SD[8@?BA&^NX9B
Jfc/D0MMSC>a8V?fbG^Q,23(b(-1[QQ:4ZF+EN1WaY]R3J+E/)C;TJLfU<]G=YM+
0YO;><@=C36<;b11)4^0U>H&U^C^dJEPXV,I)cJ<F41ZfP]c^)C/ZN\6WI3VRKX,
M>G&_0H?=4.@])4/LfDOM^KOXX,]&/da#\F9+04HOQIO6&47O(U0eVc=2bdR0d:Q
?M]:VJGCNX8)NBB/+?E-)aWS0V0[^>g5>gSY5EB?#UYA?DW9<b<;40V)7cQJ\#.d
22X.VP]SMH-M;L\=gS>cMdZQWgZK6-<dA7\L)&_LR/Fa1KW_E0+C8cE<1[.V2F/V
PV5[XH2(H-AV0?FT&C[fJFVa/@#05d5^bW/=ee4/7ACB4<@.B1VYW4-AA;3V[0UN
,-T(>I8LP]3.;Y?WgM-E4VU_>HgQ:#,)]E8R:G=4Eb)N-O1RRB)^.IB.HH-eeeM@
,5Q=N3BS-P>A(E2=NA5VQPX_YfE[\C7,+g24L(_>YX]5QBSO/:?5=]&+=0af@9Ua
[142Vg]H2:d8ge>TBNO,/;R7+aEAWgU7RDC()ZH,Q,#CV>(8?=4]2,@Q(M[#Ua+P
==WMQbZ8d5-^.@BRV=(/3Kb3]=\1Oe#+g_P1/5KLcN[V<cgW189fQRXF<?dR[Gaf
g)+f>O<@)W;^g3Dd>f[ZEfQ@T@Z\I?KMc]AZCH?9>d/)@XXKW=?g1_^N0^FUF36L
31QgMS]<UPRcM1W:9)JF;<aX:/A:U_.Tc/2W)g_/6PLUa5bL8/f.M,^E/Q?aeOZS
&++N?3TM6c(dH\JJ;#X<K4RMA-E5F=#E&3RfC7;1gS9U@EY53KV5:WcU0Y=fS\JC
Y:ZII/KZCM]4C2JR,ZcZS[M-1F#5[ZF4b#Q18+&)ZUMINfFB9ROK4b3AGRMAGZ]^
K1N^^&]Y]MfEW6gR>_e&\C>52&BF;._PIgFHgB#OK_C7OZfQ5,c=G(+&49U+Y,I&
B:&IVG62:8&FORR8S_-Qb63aN+27CCc.E.EKW#;/,7Wd-\aE.I^E>FH=\B0M4&K4
_40-@3C6.RS9&D&;-V+U1XRDBUE&<24a)DXb_,NcdZ4[BCg>_#70@_B8N9<&;g15
P_/H(.B>V&LOH:C0[;[-::8796dXO4K=0VX;#4>-.I/^8B.22+JU@,3?]ZNH]/O_
\Y6T>34=f:JMA3PB@fW,W4CC]?9ML_ZCcB4=QOQ?9CABG.XR6]Ob+5\7DW1B17SP
\e@M):]5^O@Ef#B84X-./dcA^E4fCJ_CW4Yd<Ic_+KQYFI3fH5L/-R2fITT/LIW3
9c4+IV(RGNUHA)eL?/I>4EACGd<?C&<=L]4+_H6ddB0;@Ig.AFcgK8&;KO99U3R<
gf:MGUM\d2T&<360+DZ(I=,L_bGTXJM(MGe.[CR?@d9YTGD;0\W6<#P).B/860;c
S4^_7J&>BP&:@Y&42NgD#B:C8b-4Qf)U<N^gA8b8ZSd^+LJ()Vd2aXT\8#0gV-bd
U,?&W3(?g]>B,_./e9^SeK+@M6#PE1_dT:,CO&/@a\U7-K1D-T^D<Xg;(##W#ZP?
B@^:K2>Q(,[3A_)4ce8_V?HPa#gNQ<21Cb7:M\d6&F-7/=DEPdTIN#b)M6K&MHQ2
:e^b7a(G<OOTWdI0(KX9bN^PUMAB,cK[Z0E-#FVCSD&,5-=R1(E0]&XFHZS=HdWR
70L?<d?Xd>3XKJ6,A)1ZN[bQeUUPD3LbdKE]EK\SWdVQK5XLYGbN<\A\<?SA.fDE
\AcW_F==]J&b_-NeMOIaP#W^9eME._g7C\1LKA&RB(<5Pc]bQJG+ZAg+cHLe&=a:
PE>4RR&]GU--3(ffM,0WWB48[B__(CO6V+NBJ=eA1ZfCL21VLE[e>)_Y_],0Q3P5
85HB_I>/97C>,_^Y\edEEI(A?LJ.dgdJ_E&NX;FT>9FfN]JB^J/Lb/Ud<3NSKKHF
=FT)L+HGHJ(Tb6QIL1KfR[&BWTdcB9?QK_Z&V+B^:+=1&a>+X2WI3b]aVXM5f6g@
Xg_K=Q5:=-TG;DV)#T2EED<<=KE&Ge)6)WRD^>C\6PgRgN]W\,;JP^aa]6b-\BJc
Aed25T=HA9CVOUFI9R4PV.6&TU@d6\FeHHOMAFS]\P[3\9F.@#^IE#a<MM+P19RC
<Q5gP)@6E1gUM+d2]Z<?=;0KgcI_NdcE4OY12/&dO\eOLCC<gHB[.b]T[3G.]ITb
GJ6cO,U(W1/ba.9Q+J0GIQ<)1:_U[6X0=N\AU?)-E\WKAEaKTB_\Y=?c@BN09:f2
T\SR(2:G/88\,6NL?R2N[JJ53@@4&(T6RG&1KKN9:<L21E#&+F.+)a:_f4B#E;FW
T_@>P=V216-62>\Ud5BW_XQ]4]9&g>O3E>BfKO1B9286#Na91:Z7Z:5e+eJdHN=9
5_2HVIE@W<QA+H0M<M@+f?&R64,T.)?:)8I./W6DDfS_=g&,A9OGbI8B,CdY7EZB
2)0>G8.]M,H:D1ZMV.WL(eF83Q[f;=[ePaD76B=C#Q:K5BUL;O8AR9)DWVM,;^-P
@aP_&4;_0g)b:ER2\YE1AF])H/MT2\=MDK4@+8HYD)cSF3VED1P;//5W\W7GIb?N
OX=\?6CGgEC:AX:H)FIWg<aI2XF:M?6Ya(-g6.HDJIcYc\JI.W\Q>W)^Z\?R^7^H
50D(6BK=?O/PSg_G,-RT_?FG@67;YJAIead&gNZ9_NIR.1a:A1,-YgGFH<1S]=8e
)(eLU-&Y@A1V>SA?Ze6XW4FX/E:E[<,#9D2<VBBb,\ZE<]K1TGd[.I_+E58:>/VJ
GC>^:+5XeD,cE6=T9>b/U3/K\W>,9QUZa4FEKYE?[C>32O[M7X13dUTYS)_Y66Oa
L(HL]N8A7DW?(9b73=CbGY[;fY_d5V,B3^_Ce_DeY)6/P\b#SA\]A;f7_QJKAL??
4f]<_JK6>(C?\0K0PDgPF<]=&7.1A5fOG>V8MU78T\+Z1W#26c,9W)acB\NR3LXH
[NU4URI&47194>f5P\^<15Uf[?+S^2?W.Ea1A_5aS=+F0bIV]OZ9,8f52F;/^P<(
AbIQHL09237+HCQ8ND7\BK@+4TE>-eCNZ63e.N&QLTPdb@eA?PV&^5&JS@,V;U#Q
9Aa,UNK&[>]JgI[C>N8W+K&SfTMf8)egMf-[/5T]aIPNSH&Y(8]2Kg@A+<^eMNf[
5\65d=R(WfLX;fb7L-G<EL]MWZZZ;PI6(g6JfXM497]^#Y6Xg3X[=X0dW?@8RYCE
<1)-<VG-#2bU+G^?W<]EJ9<0=U,02H>LQ2^B&H1<6Rd_^?Q2\>HADdG;^d7_;_L<
CQ20Z+\X(\;XW/2)X0[XI)KP<JSWbgWYH;PPc\]1F8Md2W_AfR:Pa0T9b(@<CJP?
\0>T-/0)DZ,^77LK&:TM4PJSP7HVCMSDZNP)@E-0#OA2O\bO/)@9N#:W8_7Kf,16
+J9@-&5A>ET#^E>G+.4EI]P-a;RSA.f)e><?b-dcA2CRFV.-[7;Z<.84EX91-T#P
27ROD9),EG<7<c#D8_PBN8U]e_Z+eTV1UH[,,f?,=B2\YgG1]IR+2FR7#&-/>MG/
^4fW?1V7,@Fb8FUWdN1Y;b41+dMDQ=bZHN>^J0fIKXA:OQL8=.;bf3E0?fX3)ZA)
O7P@C?TZd0,-#QI;[Y853\&IcZ-+f,9Q83eXINF8@-FCDD;<3=1caXdH22;eL9IJ
LT>PLAb9&LCdS>08Ce3XLVZ>=&0GHAaT)5d[He,7V-;S_]1S_>(=SCC2?:7>T1I]
#a)PVSE>X0f6U<IVLN5d9+(A:73LdPYB8a&:[)fA.D?e8AT7(9RM^JV>+&N?^:W\
dFUM3a@14/#/>#a4Eg@+O)Z@L<9DH3/K5#^/(Aa#75H)D([]Y>Y#)LCIQJ<V9I<a
RK=;KKB0eLJEB3^[#/RYSE;NB&<53/60J^W1NFFU8ACW,X]EZ#cR\JfQf,(T.4aZ
#W/CB-Ec_QO3X1VM2TFIIQIJWKO:1Nb^@D1,VR(BeXK];7af:,:3):[T24BeSbH=
D_A0:Z<7F.=D5TI_UJfYUIURS#4EH-+#S:HV9HJ_FN>#6:1C4ZXe1&G,84-COe(4
@L+c&_<Z1ILBJE^^c;Z+&f=T>gE4.8ddFG13IbL=]J;g/E^:Cg9M^d)G\]&H07Ab
M9f/?7P7CN^8?KI]5@Y=O6C(M<S:FLAYU@HD22,\+C&Z:Ub_BUHZ^;VCDa+_^LO)
LN?O<ggI.(PV8GAIe\LM,cVQSL.&)Ke)9(#E[A&4:SN0\QgYf&a27JJH5_YX#M&D
aW\&5e\+>4J\9(Xf(?LU#FSdaD(?:)1:EgBe<,L&DeT6g>2)^H^=>Md0+Q(8Ie6C
-=#eBYe84P:CZ(6B?Z<cEV,VCI-\UKd-E(5T7C^fVCOdZ5:.PO:]G6CL2V0dAW6S
:?K,_YcW[bST@W,H930\RI9aE(eK&YQ#3#(I_^5,S5LTQHF77a:[9@>M5VYg2c7O
LU\[-?99;D9@T^/baY6-./TD4ffcfRCI2HH)CSN+BgN#MSBGbJXS&]VIR=PL:fIT
YVWOd1cVS-gNReI13./H)-g8E+7Sf18HF?Yb&NJZ6b<KG=2DUHJJV)=N6@EBNK:8
,[V^J/JJFMU=2:L+D#b4@33^Z#;<)9INc]G.PFCSb>-BWgaeYE@6^,6eKC26(\G8
f\U/>BF+HHIN_1?)aFBDEVgX[U+/&Q?FfE&=]ASP3[N8&NH0X[]<=4DcZ;1R#_SN
BQ0?@;K-BDd]DCK,P^-)_eObFW80O5fADO5b#IDafEJZ=R2YNM:F79AbX@eZM>]5
8/GFOa<#S\-gJP5MCJ[Y>_G5cT;Vf:a-WGM67fOLL5N.&1>KVFeCLX//XF<WOP=S
/74+AIbeW4(N,Y;Q#PbK8@a_RVX@@0BIH@(Sb6<XHX]df(+RYdd5[-+V.)P(+G]Q
4DTZe=?TRWbK##FI+0g]))/aXP8Ke@<_P[[[67#GSHNVC>X<GT_G#UA-g?8Z6<_1
^#V_d-^I7>WcZO.SDb3YOI?KaA4cC44a<T\6HUF=7E\:G;2LZb5JRYfM#O6QXW4T
)#7=(_5aLTcM24ccVB^>_(Ua(b32b<<aBR.<KH<YE2bdG.LgM@23>+U)#c,YVN+9
HL+=-67A&XQc.fgGa8NbRTBLS+@H(eP;LDR&5Pd53;.3,U9AF[FcJF31JR=ITKBE
?]IF^GNJ.2.dWVPK(C2L).MI6ZJ)6D2bCg?LOCf<@9I-@f#S4([XL#E5<7;+_^ZE
^bP2B83QMT-fV>DWI5EX@G6_>C0\W?:+K^d(J:\:7c]Z+gTJY[c@X;Z931+,7K#L
cQO\BEQ=d>,+8cd+d=XgKNT8DA575)0-Nf#&>0IY-P1X0;,MOHXd=-e_+/J2]eE>
dY0F5D_I\Zg>(D]@5TY_\NFXJc2_432S-BZV?LTVM0#9Q2U85Y_)f@CCeQM^g66]
:[a+MP5_#Y;R67\WXg3H>A?,gK3QcTU]FBJ93:T=bHYI,3bL@H1<aFf.>7F>>XR,
CA0<HL)2XVT5Ig&b9D(+QV734&9O@C=A<OIGIN]9GQ)I@?68a]UYE=QVB4FEccgN
a4HIKQT6JbUP8UWc)I<+gfB=X9(SW4>GTOe0444N>PC[W,eBDC3e6?;I>A(&=c:a
8_^.-CN>QA3CgDC51RE&LDU9Q,?\A#O]/aNa^L0@:0P?9MCM,g0JaW#1E\:?T,2_
XUVb<@PbRFcb?;T4NM.cYE6AJ7UfS,CP[A/_,2-J\MgFA/=aY3cD?=TK,FSFf(U]
^F->5KSG#57e2A6X#U.PMA6WZJQ:<IUJ5#BH8Pe?4D:(O>?^TLU6@0:.FSID5I]M
0#0(^)Ba94C8A\6DF>6JNaI_c=:7I//BD2ZCLa@a\75Me@S9-P4<VZC\^:^Y(@AN
B]U<M@V@,45c6?-98TF9#1O&MUdQFFQ4Xc:FIM_OTCZ(F[Y:PJ1Z>,dFAA>=5(YR
&V;BRBb+O:Agb3@7cC@HRcK=4DD]Gf2NP9SR1/=<JM4cC>X]AH+;;+IN?_/^eK3A
5?g:^0eT@e=1FYL.QG:3,5+K.CKO5BDXN,f&7^EXNdPD6&B89WNffX,c&[H0WBe#
M9cLRT\F50aNbb3,I+#+LC_IR#-g?gYV,C6ASOgbB#_Q1MZ+2UJZK7]M_JEcD73U
fVH+R=61JAY.bQM=7Kb(Y45[UR/K1&:27J#O3AN_?:50/8NB#--2@)V&g<P:ZgZN
5F)6f&EK#aYBJ7IdV:62M7TYFP;f(g1L8-eE)5CHFdV;TP1)2>9[CAK<2YHHc2C3
&D6-:K)BNI)0KTfG8/gJ?;ANZ6/)^c]-Lca&D__3aNYIb?\;;G2SA.)7cEGa7Q\Z
(<U]=Y&T#O_ZT>(?4<;cg@YXH5GCK4EFJLeB1#E@]N[Z?2:^=e94e.3]0M+([GYd
VN2(@7&Mf)>)a(R+B8\GX?\Uc8&TbPVS^/@/Q/bM8RB>LGd&:XE-(AH@-)9+YVB6
?f_c[&A9e.(OHT=c>=IMYDDB&RB-UDbc[d^)F7RW^+dUU.+CFCW_(>)aF/:.?dRd
Q]S:\ec]U[A69XW54L?4)S)<.UVZ/:1#B5Q[;O>0@a(:&,B6X_G52_gM1^+?]:&2
G@5Q_6V/Ee?RY&4;S\;_D3>DdT3Y(Y)AGDb?#H9D;NYK^>=VX9^SE6>[5^N,(+\Z
[JKV0,/P/0H+BQ<-AO#E\\6^4^#U801->E9C^&S[Zf\Z_IaAc(YOGJW3Fb33-W9K
4_BB(/KZ.;2G3&@#RD5I93L\L:9+7LBB+]S\9.;>;<7PNIK8I;YV+?e]YWU17]@=
,AdcW\WADQa:9-WHP:e^b>V,Yae/4OWQEA[XK;DVM^@E.aM0XCX9^ZJAPE(19c+g
V3H^S2[(\V.@@ZUBP/DGd51FVS:TQ+0E(38/=E>[R\B:8?L6=DEb[)VX0[IQNE:9
U+J#3F/N]9>D4+6Q;CI/e1@A3)=WAK>>FNT;eE84RR@\6bLA71V4?K5G9H=5EFE>
U6;ZI/4N5PO(ac(4#A>f>,X>W0JOIH]dd9Hb:8[f]YY]T1L=&U:)\e?X)ReL4CH1
e]@g@TNVL1GD=Wg:T0SWJ3fBMY5:^cLb87fM40f5L;VOA54CR?5Q8H35K(H[,CS,
88W&f=3UYC]d5]NP7>OL7^>^#YQJ:d-0.ONe8G5-gS(ASI+?16]6S48820#b/_T:
B.^5.DKBK2I7-,TFT^R3e?AQ/+9-M-;O2ZQY</<F^-^A\MeDMa/^YU5HWOV_Ug+9
8S7D:(R?a7M>):7_4c?BXVd(+VEONU?P[7Y-==gCV@MQ;GX:SVNfZ7\_AdANE6R_
+>b\a4T[;.eX@Ib-(T0GK6\WKe-b43HaES42B+Ub^W/^ALE(4KH)XQ+SPdE19P@X
UD)G\QOge#O2E],2&aUR+JaAB/ABVV2S4351?;XdJT_===bC7UAIe^73M>:(T8c9
=[NaH,OI]]:+2)9&,M6)6JD-7TO1C>aOA(?=eZWSXZ_<OL-5bDcGIQdKMKQBe<<T
?5g_T^Bb9NcU3.N+-VQ/(eD8:.?G&@cE<054OX)FR\7cZFS35Eb3eD^PScNW@JV]
>;^FNd8-WR3W&;S6V=VUC1V@R;((bA]_Eg/8GXE>Nc)&#AZ(7F[)P61-a7KNf\Ve
-#G#_\9NBRG).D?;#B^(_3SV5Q:IB?JVEX#X2HT2+O#4&bZS4eR&bWcd7Z)UC=L0
48=fdE+3-eJHYKH^>c,+&aQ&R<7\g8#<;HRG++O/OI3bV)9WPK;4a/e3QIEV[:]Y
7V#,;#F?aR#5Y6U5^O/O1UZ#.3Gb8U9CG:ISU<3A(&_/6aSL;L<bAVIO05>[:LWM
J8#OB_6,MJLM4MgPe.?.DL2P68e^T7?,PZb/OE0eb.SYB36b<:V6ASV]GHePY[^@
CX&UGe]KJ[LTfTO8KO8N-NK2T(abR/EOZMTH;KQ+6;PPAX/8:g2;O3dg01/Z4UUc
3=d@-JB_YYLSA1F>AVVcB2JG/O[0JM<780KMQB>#1b7W]Yc.W6TPdOB6;FGN-,3C
QX.b4OP#9^Ld:;?&;b(+;b/XBafK4T.c4&g&0-_@GNSH8><8@<#e-Lgb/#V03J)@
OE#[NN<Q0,g#?9[[X\^]ETB6Q@Z&^5:N3LO3)MRYSV.(CaF/0Mg9+DZ8+)B@GDOJ
/^0C[3efA_3H&.24.P/I__eUPNN1d,_)IPNPPN].AaAPJMX<>40L=afGQg.CMJd0
J[\XX891(#FgN5>W[4XNW#0EeH54EL(UV/J]_G(=80JXRYac)_/dBSQX=^VF]S-L
GGZd/#ATMf\,1D[9PD8LFG53^:A?=\PA.)g=MP6/1LL4/F(>f>=ONe+B0XC?N(^^
A;&8f4JTROcd4G;ZRIOM^Vce(DZWI^(ZNecbJ10=VWe7Q6.N]SUF^G5U7\7:g]4U
)]CE1&P9a#A5e4ZbAb+?WD_KR=e3>2_9O;.Z)bBfc47V5c3I+Y<W2,/J\W(@HDI=
ReT/[PJ^U0?c#M3&JTed(/a&:PfG3a6>I_##[;e1AR:^?B/<f]\@gT2-1eHQZ7?>
[:Q\aefB0/3]P_fQg^d.&_D\_R3\_7S^S;49a7:K.JdOA0Lb:WV2E&QP?gOMGIIH
+Ke-@DH9)Q@7Y0g782>/baSR]_c<IXR#0O/f0F;FAbS[IZ:8O]AWbD_#R0NROIOP
-_bX-5=de^0\#UP_J760,4Le7_J@\#+4c]32#Dc:e)M/@&X.FIRTVeG:MV:;FHT7
1Q6dQ,<KdZ/VI<_3TMc/BSaWWL/VFA[TN]:Ia8<S#1gR>M:<]ZaEG=4658U#[W=V
^XKQ)VF@^N6:_[b8OGff\?M3?3X(2@17<(#VP.F+)3U?AH2?8@CH]L/XRMHJ<J<I
83)[ZQ\LA_ZcKe,;P>QFW]G28\2S/E^10EHN>VMV_E5?3J6QaV[#QR,e[[e3YeGe
P9YRBgI1f9&<+0QD=<3bIYHf7M8dW82@c(/M^-bQ0c^:-E9_N-,Sc84:D<Pa?XI;
700RLQQJXJeb@DWN@49Yc:_21HdIdUJ/2S\De/VW&.CN-HDF40,^?;WGJcZ0g)EF
BDV<66,9K\ULQ<D6K\UKWWB7P[[3=UJWRX[72QA(9M2a8-cP)b^59NgHJ,1PdcS5
X_#D^0B5K^:]10UA2TA:3G\T)3+g-/O9RK)>)+^HT7=U\<IRc\<U^?VP&CUU+c8V
#aIPBNZZQBg=_<B/?[36A/g@^:Q)DeR7Je4ad(6]TOdOb[dQ8_gI8.-)X1SR-)A>
EPWeU&^W_\SQN/VRXf-?X,2QM>86/:OO.+UIY<[J^=JJAPF6#b83>,@V+^VQP(3E
)EI.9NAg_aWH.X&0I5)9)R]VR9Ke=Aa9VL>0BN+f@TY8B4U/@MC(L41Y0<Vg&]aO
B1Ne/Q4H:C8[VA<<>FQaa+M<?(<;K;QN?<S+/K&9L5c[]Kf]0<Hc0.-RJg.eN=Vd
+3Dc;Ob0VNeKf)+EH,#KY5aC,+B&Vc&MQ+EN;.I1B.&VG+X8+ZcSY8a/f,&.<[+H
cY8>F^/WT0#,gbK#L:1]V\M_RX^DQ6##=EGYI_D5e6MO2=<G-.R.;4I?_f0&V<2F
2)OHW2NNBFW+fJ1QFUaGf;gaAZ?U;@,PaDUQcR&,0X-NO>FcAG#+\B7BM45MN4X\
Hff7c#?\a:9dY_]ZeaHHM]RAWQ??6JY9I8;1Xd]E2]V0[Z8Oa=S&B]:-R[]K5&TB
USTZ7B=\DD/7e3=C=V40AOKRAO&9TZ.ZcfYZ-]4GO&/,XAXNf+2R.FFET-1:/KP<
Q3>W]VJEYXcU@,]O@<E[RNJW9URS/X]])CFMZOC\J9PE^X16^JJ?;;-I.TKFBK<4
3U/A-AD_:6Q-5;<E@YW5#Ja6]K<5eWUdgQ6/-T,Wc/F1#?^_+2-@<U^Me9/_;fWH
#_gc5gL_ST]_c^(ODFCZ:H@6e4-BYB4ARP2SUX0bI_aD=g^HQ9EC<f)ER4a0#_03
-M\C=VOR3I#F/,NGH_e.4TA3cAA#R>VW1N6F_b2>T5+JL;PIa4_A=G(+VB)F..L:
M.US/\MS^f0P9-X@1Y@B+5ee.]4E<dN<);KCOga>Y+.RA<Rd]<<YD1E=(4Cc[12[
.6CAT^=_-P<LF^Y/fZM&=B^@CI_AR3-M@)E/,VKT.g[Y^X[^B^JIVZ_OCdY^W]N.
71OR9I&09FS1TL[(/@1BP3,<=],]G2OS6W&@RE26SLf_6bR.?dGE&e]&>,3[=?OC
P<bKQSdC@6[WXRX3\J\>8[.S&-1QD(KH8[R,+X?V-F,_TcbZ(Ub.=VPWWa[^4S+2
T8XS6:eTGE7;OTB4:&b@E(42/A[7T(X]2bU^LX;8]H49YcY>SS,5YNIeQRaIZRN,
b7..f2b@;U=-R0;D2Dg3eB\MGC0TC6@K.KH86IO<Af;X(=S43e]OGY3SZ@67K\a0
&+LUe]H8.>31[?)IXW0gc8-=Q5:<#Q54KW13:9#e349cY(-d4a;&8E?3\[5+GJA1
8IG=<2V4,QJ1f.>R0YBWCce^64=R\:K2I=F;_SO[F]:FD3RVORSK-FF-MW+J/OUY
McZ-B,;N#>ALGL].Da<((YU+g</)];Wd:I+)+QB>gI9bKPCKEgQIE(M)QBL2ga;U
6OcA:M1QZ5E[+0QMX^HF8F)<M&g-437df(S/CWS>@E6L0@9WG4(dA\K8AB;:dO-J
CXV92RF,G_0UVB1KKdF,GXFG9?<?]d99W_8E7=9a?.M5W3;+c4U>g#D?#S]E5_<:
UJJI>S5c9(4I\LXgf&ffP2:-?&5\aD<)=(BfTNdf_I1^F->F00:/B@?AKc1OJTB:
#fL.I8N4RS7NWQ2?dPe@[<F3_;PQM0A?8/d^_PZ6^-FN[):(I;FC0H\,Q>606f=5
LP1(a&[BZ71@B3KW\KW8@W:fee^)bceV/(U\gI)06XF<A6g_4b/e34d\C,OQ.)7d
BJS:-W[YNNe1CP19YIb,<6:Za.f2O5/MIYfSJdY(aCS26BG>-QOP6cBP#H0M3@PA
KMM.8_F>[FZ3LIc+K\&K2cDN>T040-f#QK6E==)/UFY2ad0F##_7:4+Q),+Q]=J.
+J:)L9dc9acOS7+\Q@M6]=]U9-GSB\ZZa,8e9GPD8NW;,33,@G[K5,aFbB<?8Y<L
YAfSfXR6_<I\]>fL-Y4&D#79X.cM:27a;:aNDXeECa_aS_dPMeE66+f=D@TE1P6E
f=d6+LJB/cbG1X.(3ZJ]V07T+G#,\GeB#f5/d#bRNI[_Z?Te;(a#5_U<.>L3<dO5
aaSVVAPfObQ:S-?18J2HH^1:e^cC+bAOcIg5a/Z887CLE:3_@OO^69]U\]L^WB7W
]N9(,/&.#[fG)/:TTQ>c+9R1+bK>FXCDO541]eUA/SKWLb,9JgIIWGFIW>U:1+(S
+d\gdLO2&=[I3EFR);;&6?Y3c_,AEC#(R2I3Z=#F&O\O9=(U8bIWeJ72bTHIM.WZ
cJ>67STN^X1##Q(WfMG,6>2VIQX1fe2f><J>&V6XNI-bP&/CIfT,-JSHCRG6-6.G
U&7WZ)RZN1Eg^FU(b>([6I64JZ;D.d&PT8@-DIG2JN6IX0=Ga73IGD^V9<5_P>ZD
)QU=;A][PJ_3?,b_F<L.^<DT?6Y21N9()^/9X4^.3;\ZUfCb#F@eTRDOHD5OY6Tc
g?g?1.VW6PbHE7MG?(QF+;,g(5TI;,T^,b\I.>HYINDaf>IXH(La6IaH03?X5:c9
D_OLb;Sb,I>@-@fgFa[P;N?5I<2cI9/SbZ3R__(Vd/K=D57RD?M\ZJUM9AU>5O1G
E;-b\7\ZRfY6M:P\?@55R6eVS_MLIa&1B[11A\;XA5/WI\ab73&7_]YKP/3-Sc89
M>Sd8,1-/&#FQaE?HSQ8SW^bcJL.4QL/N2)\\9,@g/&(5PXV1564^LJH2P@?J#Xa
>]P.RM>OfQ<Z#L0S@ge3dX6C.N3X7/_RZ3[B>D<@bfSU@\VE5^VcIH&(_^\5K-]L
cQOa+&@bG?\YB6+F/.@]b5.D]Ff3YOJ?.IFJbU2c0MeC,QS_:d39C,__:.DA6O;0
[bBZXFT>fIL+GKALG>ZbAM.DbfCTS5):9HZ]-OCUVDBZfLCT,RRE.5M6W/Dc1gR6
&]&]DMI^R&=]RDDK5_]/9YT=).ZX#6M#5eUe()+aYF87&?_f\K4MA)FMFefL2=bN
MeV+4N:P#Y9b^=dK</4FX4JNOFITJ,fd1^[7Q+D#MUdeb:;gHC)0?_T#SE[9dC=g
#>HcNd96MLc8[NQ3Z,\G5&^eD@4@Zg]<G;2cR++V]e0P[YOd7+1QP^>0#YBRVUU&
^b=^XRIWSZI<SFeQ7.[8T;^3;SW>D,^QMOSBZ-2f.Vg>d,Z/D^KPaf)6=12(1g++
G;\8^3=gV[><TBSa<B-aF5O[T>4@\ecC#1a0-JgQgTN8X]Qb7=QIb&BF73T5/P#^
.]?f>bcS&7M<+a(9cPDZ,c0e#Tb.S/@#2]e:]]d#./LS9UN^A\++aTE8_BdEHEGc
(-C4W-IG9:NeK4<>@NQ=eVW]@S)]E&<YTD172>0NVR3RO^&YZ<AR.ZV508P@Jf:S
13:?QA+a-67YBc?>=CULN<T?0#e,BHVbVCV)8faQ]3/Z=IN<J7aBIQ+a_D?D^VOG
?gQ[_R,E<O^;dcb<HdGHaL]RL(^48_?:RgJ9URFgK0D5P=5@/@UUIZc:L73E?DHS
S<<2O@V(C1JHdRP3b0d9JgFga)adLgNI6@]gT:B04)O.Ff911G>M&JJCb>1MLaa?
8:O:Teg_VNZdCC.(gOIA]TJ&;aUg3QCLR#4<aTW161G@-+dV_3P9c:6:Q>C,E6R#
($
`endprotected

`protected
eFeYS:KKD#TSI,:^BA??L_FT.FSAb=aGT7;b[E@Xd(B+f/C/cVg\()MV=)f-Z@^J
>cQSMf0?I6_D]Bb)5P8cL.FT4$
`endprotected

//vcs_lic_vip_protect
  `protected
6L[ZSNKgZ8aAX\<XFM;<G\2g^5SH[Q],O?^&gC5_[eM.Le>;:]KF0(DdP?(7US\A
Tf1(KNUCXS]A5f(/RRDB7;+?,V8&VATC0DQ-WNG1:@O^^>>\?H1Q,--]LYd9Ce43
fN.J5LY&4/Q;2EH=_;+#>NDAW<.)-&QK1S5-,))bG-Y,5573X@N&]AQcWZ26UegN
<QBe<602VQ7WZ26BA#\I+3F/RCGEJYU-JVJ+0eC5B00^I=S82O\=98FU;^KBSEP(
M_(NXS(3gf<D\3Zcg:UH#d,g]=+,(\eK+)+RD73+,Z&2fVZcO\(cDb^Ne3gPfgg,
Kf@fa&6;&bRa:;IQQ56Mc<:.YMbSHZgcIISW3L6C3^A_^;L0JQNV0E?LK,[8-DLd
HP1a+_J:-+Z];=(FH=@M&e98e=E)[6)a]3-8A7cL^/dE/7QT&gU2X<YX\(K\3^3M
P;cc5L65B+OZO#&1RCWQ+BH=/R;B8Q2/6<2&B2>d?G<#A/d9?IL,HVH2/N/=X.C9
@H?+SYF92\gVc3.b95_3[Y<RU682QU#TN7EO@I\Q=HGZO[GUb[b.JZ6dab(=]PC/
B#BQ)-J;?9^C.-H])U7^IAC=ga=LcKeP[H.BgH9V-IcbC5J0^&TH([6IRJ?MaXe(
#Cb3<cGU2BFA,Tee:MaBgIH,#RKMOUO5eO\.?^A.f?M1J2DEO/I]ON4^M-+]DG],
MP\R0Cb7_cbYERIF6O8-B;08dc#beX267\e1fE4fQCa;>V5B:K9^_=BZR.XZ&Z8B
Q.3eYA-f]ba-EWDJGE2aa;&8)aOF[TRaD-3<#:A9<@7#X,TI56f97VHE_;NfBBa@
JG]I,dU?T=PD4Ag=.-&INCc4,/_=8N=RC0LG/=LVQ80I/O?fg5Ra9TNd=CFdEQKP
JWGe^g4KDDT0Q6=f^<abCXI@Xe4GI-J]A;HM&M?-Bg1HeT,W@Kg2=(CPYFW-,Gf\
cN3:T0F@2?ZPe>-LV0Ygf0:,L+<.MP2-;)=;GEN]WZ&;-_0eVW>AQA_EX3P1O0?R
,4)c9W8RIC[(O?]P9\eb,eO^GF)[):>:X_^G[1C,1IK_/6C;8<VLLA6=/-KAQ.@#
6KCW.QY]agZB]cFQ.ORK&@R=K#5A0C,\_ScUOKKf8WI?PM8,W0+I29DNS-C8_.)6
:TVKXaQ<6<_f.UbJV:_B(L9F.4b.PfCc#b/]bXHYRGR(<?)+H<.C0PVN.3:?1-,Y
JCSHK7G7L6?KPV4ITZQ.WOQT&0(YWQ<HFg)24a0=,WHFbbfFCcc&1&+[W84A&2J3
JI@8JCPN<SYIQ</->NfWc8;B5V#5B+BKS78ZH<P-.\BcdVOS]0G&IdUCQ9[#,:^0
c6U,bb=THI)/Q></8JJZ#JY6V4QW\3Y]VVf^(@L,K1HXLOOa6AZBO,NS(2994T.;
9Q[]NaY][P\#W;g.)/(PcQB87UO.3?X.;B@G>^KN<g+^RRd:<NABP;F<S@PdA#6a
R6SK:Ta;J(;?P060^A^5HPg1L)-BYOP/=V@U50a&7,+(gP>@.+0,REb7XYS.d8]C
FMLZV_N4XDI@fWOKN/Yaa.>c<>T9:Ma(FWN[_S=3=Ydg514V]LaI)LGDg&B?U6^I
^.4Z#01[1f=G/D&3KKAdBIXYLC971<D4;.1;F3HgG-P-;5EXA,;J?be+(&ME#Geg
ZJ(gS:\]E=2c&gHUHP1F;WBKVY_?\T?LF:-+0.\f:d?^SgQ]X[8_+H&LS1Hd6KE/
,#[E:;a<ZH1f_3L4^M+FFPQV&^5_Ad[M@1dM#A,9g4=P@F:c3(T.2@d(1LK&g:08
&O=MQ#QeBgSge_]LL/DfK/_CL<_91H,5?F<_XI9HA=L=PHdMCU#/g+D(I>f5g.2S
0@b4>+2<JY);WTCTON:,]HITDQSPFX0M=f^IGSZNa]Ea76PfJ@FXWdb;4[7]#adG
:G\(C_VZY/+cQSOLC6U?RD\W^.+0&[NJOdH0<:eX[d:BgPR:;.PXe2[6L)FbI8IZ
<>5>U\(\#J5I@1\/7N,;Y\?Za[a8W>_#FIEcbVA+1dZ5/=RdJ<S,2ZZ81^\1N)+D
.]V_&[,f9a50=Z/Ja^]2)=UTHQ_>XF;ca14U5(1_L8<ff18Z,G?V[JU1;-dT=e&U
^TZJ6^RK=X\PS-WBbg)@eF0W/,?b+=M]BO#I:;AN)B+4^GM2eb3\SJMUBb=B=+R7
d0M25_;=]GEH2Me=1UM>3XE/]AI(4XCU,]/+#4V_&Z-V3+]7<N[>SGaN.J7/,Fd9
Y]YAE=L6GL0WT&K>PM>[&KRNeSb?21??_IM<:H)DQZ94LE40F?C)Ig9^c9:;=\D8
/D+O&AV&DT19\d8X#MNC)5:_I,,2g,[U+QB)RA5W+-RNPPCXG=1gIQ:Bg#d05RH<
bG50Wb-7QCcbT=8/aHQ@9,b[[14,.=OSO8+fAD;E]O:703RW:-[<QPH\LI>39M5-
T8^NLZSb>+^=9)f28OK\Z?)RM);QH2e2,4ZF;#2N/a;_V(::G_Pb\g[/Q=P\TJL6
F1U<^#\T)4G>(cI?Xa7S_B,^9486(X>E7)Nc)aU7>e^\;2T]f(Af+1?PO.f0#5f>
\]GMYdX_#TUd-YfeB/#>@PUT;gJ0Hb^^Z0)M&7GUGU=??[+7b9e0+10Q->Jc@f@^
D/ULeYQSGE(POM:8Hc^P)MT)9;8#.X#VO9/N]FDH2Q_Lg=-E=8aKWD#YFd;VGgUU
ceH@1ZQ0/)MSa?YBC#M9JVL=IA1)TLEVI><-6+,E1JK@P=IFY:C,CX>eUH1S?Z:9
/Q>ee\L^aQVUM+SLbNE7_V,YT?@3LFQCE<(EX[eJ8]HN>,f7aG@Y.CZO0/9K:N7B
T=2:5:b1Tg.2EB&LQDVHWL,9KR7>c]cF8N<8SaC+?Q,QcO:,_>_.0<ZYJ[@ZdVEB
F@eQ]TVNd,6:QgdIA>(d-G7dCQAJ8bX[TNZNTXQ:37))J5+/#W>ZDL[Og[JF<Ec<
28^NXO+.d]_84S=+7P0Y7Q@:FAK#N^.53(.>,O0,LCMAA;^Q5dYB8LCM&83.8&c^
PA+C)GJ9_IFL@#5,gGNVY:NRA+d79_1D3V6&X,,T@d+16V[]VdacQPH87dG+NY&I
65LQ\bb:I>>=TQ;H^&-,N2.#A-HENM\SYYe>@a>QBJW),]2dSGdRDga]>E@_/cM_
+-^;N_/+U>Z(c&5#:SRdc27g?K+T)4aD)A&]T@_KMeeL\(6QFT_GU220?2\0^^(-
_f+D.YZ>#U[QU=9(4(+gOV>7<V\Z+/LNcOJG0XLYOQfM9D24cDg5K?K0[XF@H]U>
3I<>:H;2J.)_>H-^(4<E6ed=[=7.^6-PC]0IF1(=S&)@5PBHF16?-DaNJ-(R&U3Z
(/g]U_&2@&3-T+;g+_dR#9SUf:gZ8>Z>)Qf8@Ac#J7BW:W7bXR,TRd\T>BZ]?GR3
KH/5D[QbEa_,WdWR#JZ65@>bcYT3L4-QMZDC/>gZLXDe+2g0S9EV&UJfBG\>K5-:
[S]ADX1Z,PWYODKTZ/B86abHYLYSOWB=-OO=SeUY2=0?f#XaI@7X2WEGVUV\=2:A
BeJD5D;R=30cB=09W8gB0[_538^8YR0B55^UEF8f42B.Q9R=M((YR(.Iga(IQ0d9
Ef4ZeLDBIZ02LPZ\FCG)FMd@[FI\7.7RHSYe[SHH8?:V#+P;FV^cLQ;US4B<>931
G7Y:8F^:NCTQC(C4KS<7aV=c9R0M+H(fCe#])E8JRRbb[0/YLANOR<,,KM[R=VAG
g@6gZ.[@[\.FaXCgCaA54]K1\EUNBWG:;T,J<7[+I5Q9eDa[183A1.?D:UF[YOgW
]Sb62A4+DVY4+U;SSVJ0H(19^P]V4HA6WKYHBJ@/f@]:C1:8/\<f24a8F=8GCOOc
4e0;[F/WJOOF@Jc&#0CHCK0=.GO>+YgEG3,M)=Jfc\G&WaRYB:P-(7e;F?G3-UYe
[0;)JId_K9a/SA>8YR0+2PX9IfBR7K9;#[8GFc4>_GKBdLfH8aVD[A&Y5GC9(U\F
ZF.)0)/A_cc\?S._7GA(7D)C3L]VZ4<7#eT0dTRRZ2g&ABTeb.c77)2c,ZR<WHFJ
4QUaV+BD:@;XUHa@GD7V4=;MVAdLNS5Z[dQdK5]gVAgFK4/<6U/YF]<AYFC_E86e
N#Ng^b]9eS&]NTY=bcYATCMV\+)6P8W505b,)TDG)\F5)[H<B^QJa5XR5MBWU+O@
GC.,cS#g_[<M>>MS6RM[\1:#JG)?F/92[I[3TBX&?V;B8XU4&5A&&BUWD+NX3=T0
D(N#WW+=)@XM39\AQ-Y;KOVVX5BY@(Q7dS1+1DPJS&)B.T+fQ<Q6)7Ug&JVfRW.S
5#OcQdKf9WgMP[B3,XS=1]8g\gT08W@5EdReSdVUN:OWPC5/#>_4f<O8#a-0C55b
YZBf]59cLL34fVUA@9J<:dZ,IYRL23?:fK0,#RaK.GFBS9d_ODIE:)N#J[@d&/6G
G+L^Q_F6LC.K7\TFf3&8aI[=fAdO(8&c80\Vfd@/#4:9I^X9-bF6A8AQ?c7f_8]+
2b6REZG#?]_,[8OW?]C[2HWOX8+Ie+DTZ73aH+H7=g.cM>YO^Q??3NFIBN&GAcTN
2LD&-(b&\CcZM-ZXB:K1#[Y.NVT7/ee0_(><OCK&TNYB;ae).A3HWWYZAc?H,D_g
&MES?PWU7[#UY=7f=)7]V>KY,9STS&@6)K2LVSN:]#a.4)],2aEIG;AcZ8BI(E-6
dMYQ[cXcOR:FY>J?PL6Ge[e:-\:CbB?ZRZGYFbISZUX7#a5^@\1Y75E6N?Z8U56Z
,I,V2B6f+KR7f.g&9]-@KdG.)/R_TCIXL\+?dYE@7\2?[)(05JQLY4_3g>@R\@fd
\[:\\-1HU(V_^/_I#d51Rg.SOgeeT\Wf8=]:aK?I)TTL[dVW2)Z,T.4?@O2@,PKR
_/Y9A,@bD:-dPZ3_f?H97I#N-3H=^WfD,ESD\)4<LF]\AB;4e7@[<D(IE\b(=c^3
B63I#^Vg&QbgWRA6?F/CC[D2Oa8S8<ZOCZR+cCMAXZGR1g:0]ged\,QOK]<^AaTK
J2WLS/c-?1(FAKSfX4(a\GZW>eg4,_I@K7Jc)+:A-QAK6cHKab5BKKdI[ZC+F6.(
eUKFIOD>#&[7<S7L#A<39XA;T4.T[2\X:,XC+1Yb?NI/CTJWNTV.YVK;/bB;]62C
FNLTcd1E-CdN[39d_+@F)eU8bXUg-@/BU.e4\4Q27T9b[ebReE.FLA3[N?@Y^7<B
QW5gJb9@a_YG)-<+N0,-F_DBa(&VVEUTV\NM-YJ[bcO7\23Z@TBK&aV3cTLbK?b;
FaYO[dXdP/K_/JF,KWaZ9D,CaL1ZFYgg=,3Y^Y>UQ510[>c05I<4@KID3U?]\6+.
VFWT_V(bWc;5(:JVLeEC(&PcYd)-YU5gXVbbd&#Y0<-[VAR9d4&I@Pac5fc(#;Zg
A0RY=A9/+/fSc20:B\O+9.A18\9<XKDQ]FE+=++)-4^e8dJU@60]NHK0IX[>A7EI
6-3Ef>XWZD+a=^1=bU##^?TBJO@)2D<\a2H&:#:Q81<S1Z[dGZ5MEgdY5MJF+b5\
\E\N6:ADUIA^[D#AA=7Ua;8RPS\f\5WEB2=6?[SS;S71RC\S)M=KV^\#HV.eC-@K
H^f4>e]5L@?KG18e4W6V[K:GJeAY4&B8K56\/ELe[:f\aeNW#aO9dH:OZ>)TQdMe
XJ@7?9>>FKPa&7.WYFF2[RAS,^>eV.Tbg_N3(3,O[4&XE8<EG6-)4OUP,B3/<5/I
MBE)gVdZ4cJ9RQ#O_WT<JODfH:7.3+(5Y7g&,X)NJ_fM4R(L@;,V(CJNMC=LIDUO
MN^MRc1R2#A)RRc9E)SdI/?I24=@HgHSVCKd<>IN5#1B:OXGfM^D7J92/+)(\=L5
L_;X3f[P7+QJ6FaG14P/WFBRO.33UEQD^caW)8&->eUA7^5566=;DARS6C8fdEOH
9VNU;\NI7D._4K:(52<4c@7MHYZF2dd3RP?6eJEVY6fZ(#5=I;cC41E-L,aQJg(_
3W+IT9K\/g4>d5FK9E(10TT>9]K>S7##HaCfOZORCLDU@PA&@9SV/-8ga4P<L<Md
?^8T=gQTE(,d1805b5N^8Nf6LU&NFZUDJD^RQCCH4-XA=e0Ya,F>0M3>]4TQ\37Y
PN[+^QZMKPeHLgOKae#^bO2Wcf_)6>[ILCLb?f6(9Y\;A;;F9e<>>?E6J]:/d34K
(fY_#43LEU3:T;ZTD0_Vg\067(>#TC2NVBETZ:0DMJd#:G@#dMVGg\J;]NH@?-d2
J0.U397M<H<GNW.KFPRWP/LdU0L&K>G@+(eD?S9IG&H?GEbf[=D,eB:O@:#@0]fY
WEV.\7SS7=]>5R+[66&SYY,.RdJ&WLW_c,\DWGV8HU+c^>/GIBZ&->M@/[_ONDBS
cMRa->.M/#Q-TbgJU&65DRMS-[C&Q?cQ.Pg[#Y]+XX[2S@@AI-VE?_>?Q494Me09
<4_V+fK7\-5;(gMaYX[@MDWGIa\.1N>^Q.KdKL&1\aDF8D0K,>T.584Ed)XQLE[-
TSV^9P/6@UU,^R@KXGU-SY\ZLE][E7]AG6F[C#2;BYL6FW-1(IYX4IJ/JMN2Tg>9
7D.NIgZ,0gK-)U&5,9XG(NDYT4.844E9VcV5EFCJf@4JOCHQ7eX#&2_?45,KO=)^
^CfR[0ZQ33TZ8e1W/=ZOU]=A:HbA]659\C.J/>;]>U1B9>(5^ZR66N)SgA+0^Q7O
?Z@?73@:5G[]L;eMBRCPZ5JGQ]XT[12F_NeAJV[BV_4c)SKD<:OJF6RFX)-7>eN;
/=WMc:+/ZC-MLYXUAaEa(#0IMS0eR<O>A&I]^#YYbeP?cg(MY<O7&U)(#=S;(Z6/
D+)bS;BCgHP@_cY<Sc+GQ>Ba&S5d<^e6HLW@dA+)<X9^+_)7@TcLK]?E@Td7bA)@
-CHSZYB9@BB]I(?U[>,f9:(EPJ\Q&B]GW8d34V6(YZ9UU7d^1;)21WRR_,W=QNfD
I:V\R^d>J:g+OPRPF,\(]2I-T7a<RK6349AO.>=1+V[6X[e6@)]=FFaC?6N)LdN]
(4C[Wg2XH;[HYeQTR;g7/6,YT69IcR7>]+d8EfeI0Y-W2a_e=J(AB+]#[VL4U5/\
Z<A,K3RWB-_#\D2<Pf6D40I=(.&6gd<\6>a;\A_XF[P[:bK5X\HLX([2CHdP<45d
>f=_1W<F46Jb[:9=^Jad(246FH)W<d6K/10GKKUQ3WCLd&eV^YUZ1AH(fIf[[eM0
<e^X+bg:)CdO.@HLCU4eS?<2C9e9d4,6JCA?3P>9>-?#/JI2/)P(g0Rg3+A0\^IS
PO\[M19YGSR=6,FLAM#Q8QT#ITTL+5&HgDHb9[\<KaW7Y,K(4.F(5R/JcL\:]d4U
6_Z(>XZ+^[+OVB=4=T1;)fbb=]_ZaS<\JfHOLUc5Y);R#G\GINGBV+Aa1ZE0<:M\
9@KIT018S.@E,V9JGSG<Q(MQ,;]YI,?/_XRIZ=c97>SO(aBJ94a7:-^ICU<<K@+d
AZBT;J;8g(JS5FM\IUD8ANW@S\J;_\4LbN;W/RD=2+4[]c\<)Kc@?2d(P-,^B6;9
QP#.f.PL:dM<12^#_a:#G^U?]W)1]a9f4aa#O2Gb=2ZV8BReXH?D/_VSH?(e4.Y.
=_H?4dcJ)aQ]Bf6?3W^(>RK&)&K6+SV[XF]@NGbg[]7:FgL+NWcb<YbJaGb9^1CW
a6A_.Q#NN/TD=L,[9>95<be<^GdC24\0A60a]<YTJ=,1=>,:<R52-ZIU#IF#+.YE
.N6CEe9Y41c[7.0VE6_7YM9Pg,EgID>-<&9QA8JJ=G7?OT8;G=b+4<e57:\GB>XO
+fC;fJ_3:9e4?b&AF[1.Q-f3-\Z;d6>TJKW?7^/8QAI2#/:Ea;U[X_->ZWVK^E3b
U^7#J66GMT_A8Ma1VNLM.9562a(X5)8?0e;?5=M,B-0F3X2P4:IRLg;0?#+NBOX^
7&;a<P]P_FfC.Xf<K@-#]WF/6=a8R5e,<dXa4dN4Q:;\YPZ#-9H8,K(/33gC\KTJ
VO^40T0@25f_27.[TE1?b;6(K@@:#HLe@7a2S-.I6M5687257(N1@c58EYb6D+^,
gTY^1^:</</=8F:S&__43^D1Q4QOQM_/D[MAf&CB:3[0FB#V?;9_?5f/A)b,+PB4
dQRY>>8PE=2:./(]b^FTNOd9Z(UZ3.Fb]OIeJ/fc+gMBD<<2Ye,<VD?Q>G4SbA?I
8EP^IR5;LU;,90&2LZa5WJ,3V9fT8V]YM)[BRD1^IHc&NK\,D,/_@,=NIgB3ReCc
f-6;CR7d?D5,>K?:D1&(N\Q52J5C:?1d_agT#fJ+L/M,LJJC?4?MEQ9a6H/>[TYN
^.RS.3H2QfNP5=O&0?[XPN3+Sd?/&0QMS&GWbM>;C3/R-S98WLKd/f49YYTPP4M/
8ENZ7K]?&7fNT#=e9ACDC2O^Vc5LgD;d3\Y1\]g;d2JW_YZPD;2GWDM(L?HaBZWR
0[/B?G8Z/E#^GB\;HZR3KeF<a@U1H^=VY4M),[WPLC[B78,cM1+)2@N.Zd7EZbX^
.C.=S/dK+_R#Xf;gMIVO\#)_cQbAc-Ug]I;5)84eU4?YgF^CQ(EBKFW[9<+=]W6c
a;RWB93YGK42eWC.A?J;e[Sf0[73Xf+0BU#JTQP^+RTX>@PJJ,_=aEQ+5ZJI/gaN
)g_\67D4/6_78H\2Z&9&IZ5?cYG32dX8_Y]1OFHE^Lc^HKgbP;LVD4[EgWPK-M+>
COAbY6EgK(3fT?93/E)L4GAg5/]&=@eUBab72P?A-5+:a<Z\Q\KHE-5\SX5)V_XT
S1X[B@6(V8BZbHHRFUaEH=9QQ_,_M0E-8f)@41H[UO5C>AL>Ocg/(MPQPC#:FAFN
62G0L@-;.d>1gV9O;:Y5UPUENFTW020/NR]M6L5MZ)Ka>HfS//2Y^48BPEdFgB5N
I\^XL[Y.M6NE26?gXEG52GDQ-/IVVA,^]NAc)L\c1Y-EPV1)68P:P;G-,XM1P[#_
5M+IaP12<PQLH0CI_N=ebBRL4H2a]_PI>PSacX8;?YfP8/]0<_e2M/P:VG91&_DW
JPXgB,G1McMX8GW(6J&0c_KZHW#_LKH+@=L^)d3;YHDNQ9gQ;g8W7c<KCV-0@g\[
>Vb3>fRDUK#g<<LG@/eZ,,[,7\\+3OOC6a^_\cPV::GCQU/S[NSW4AOTTF#9_,9J
8Z;X+X0H5+RK^-F0Tc99MWFH>e6:T>ILG-b(e[>Z,3^(PDe=>W5gZ9::FF\?G-/Z
.U186B88Dc78J.;N[,OV4@C#@IDAYO#=cN/d15[GKH/,_3^-YNI->FM@C/Zg:ZID
:,J8L-7VLeNON4NS+e9CKI?b/DG@HS,UT(1<a?S1agPI7#W_Y9ZPXD69OWNg:MW>
0V1E>JeMVB\@cP8ETZ?.c=[bWIXf]B]O>JJg_S4>0G+/232]E_@IJB&R[TV22I1c
X:3O^AT#-\#fAg6NX@_5^;\U(A(f)N4:@D-5S5bH?AWB=OR&UeJ3HdQ?=#d9.-^J
1Y[/2;LJ9=13dE/@IWU=Zdf+#RX]RB#6+PE66c0&8Sfb1.4NTTM4\>5,@-B7H=@5
8_1[V0_XLJUARY)W28.FV2KJ0N7dT=+F8.=@NYeW;d@038Q,ML(3EC#;2<=d5V0N
YTZE?0EDOcO3>IfBB^Z@6?,[gAK,NgV73:/b_8AR(C;.I?1=]b0QAdLELF/8+V0+
FNOQ^E\)L^#4I[PNa-,8;d>Mg_=<5CV<5E)Q_4NN<PGLb.VWXOT.>_=aQ\HC07Ub
8M+\\CZaaJUC[cIT9RH0#gM8<KO@N4<Cea4@G?W^D(M#HaU/6cD0=+-67MA?141]
\EEQQL8LPF5>=-Ne\>3[VX0UZ_UQJ9G=,+[M/gI,JZ^b&4OH6Y\FJU^\c5Q9.(6#
.a-gbUfAJ6FJ.9d4C>GJQN3J^cX7MfMW,dFU/?/925H)HgNZD(K:[B,[1Ac6FY6a
g,NN(N1C4fZ+>9Kg@PZVbeNe.eNOUc6VJd0-R2:aXV-TI1FR@J_5G;&?WA04&SNN
eFPG-ZM0dCfR^YAf0L[.,M5>W<4.GLQOQG.NV.@KefFTe6KE^AN=MIe^5DO_MXeG
&CT2f68A:D,AE?A8dN#R]d)W<db>>gVW</Q[R9M7#GOa89b\G(93Y_@aaZ(I2,X4
^F58)/0[Vf(T2>GI^-=KL.+9(S&T-FT_PJ1^b8E+EP7BbX:#c/V,ORc1G>bAWYOQ
K2Hf[CN9Ja:c0O>+He58@fbBCQI/Ff:f:b=^PJ_=U61U;QKGS7D\IPd/1<2K5(-9
WWUK329KA]7H;GZFOcUcO7UW=ECIX.EY3e?Z?\R6J\G,_C>3Gd^@T54VeL?<OI=X
WPR8I6Aa61IS-d;4]7F:D8&+b,g>NV72/6I+73],IK&Y+L/:aJH>g=<S=dHT:VT=
M[5(f;>g+a&:,1;,129Z&5]\<TNG:.-V(EV2.LN&)^?)&UB\#,M/CH/W/dQO716N
Z<X[_A/NGF?O1QW\ZAL1+;FS5<^RI5egT2;UGa]@YEb+8bIBOb^M3/,@UbE\^T#I
CV<0=[TZJT^+=+M6Q:_2Xf]FGS>H>,-[e[Q_?O5MJZ@5(CbeU2R=+-VJ\U2ZC[()
Fb6@T#]WU.Ic1_3[#,e<WA:Z6dNWZIX9B:;SUb?.G-6c>@><A80Z#&cU7&+\eIZ6
ODMG-BB@TYb-R@=0BAR5YZ6NR>7G<=ZMF0JALPcDJGL6N72X6PW?.<#2G)FXbL<:
F&R8g/ccM&ON#=5ZI5VG4M45R_Fe9\b(.146[:@>-fBW:32PG4R--[ZbWI#(Qacg
e:83XZ1&g]JY/@PO3?A3^2H)P.)<I\XV[OC[Fg-[#1<I]IC;ZPXGfH;K)daB7&\/
2_?YCf#U0K/>bNWGCS\1YX+S&:MZAD]NNUaV[eYAcB#TV2\,9K8e+_[1U2c7\/,^
Lf(6=.[H9S_L=/ZG?R1E<]c<US)+YPJZHEKM^-UbaIdW/V2V@=.DQVD^H#7XF6]e
XgK[E(XOga5W2CQSMUf/9D,,_G7Ad#K=[G<C\(#UdeRS4O0.PH/]5;\,S1#?L-#T
;>^4ebEc8BS@DX)M?9)=c9QcdPb\YWTF8NB?<^c_/4/K\QSL8LP3>gcf.GK\QO2M
a-<dU9gO^^-/Eb2RQ)cXA4IaE2CM.<FWP@&UJT-GBC#Jc=CMU6;5#AZ25L06/a83
XdV(7ZK1_U4GJQ:b0b#AL=E,@>A)a,\\Pa(9FS6S6=?&+4E3Z_/&><#C96P[/38U
OW:bCGe.:&LINFSX^QU^#Y<8?a&B2L-IIaT)B3NCg:,9T<B\d^=8LW7NRQ3DN@W?
=>BT#ILNd(K0OK?:d(A-+7-f0UTOZ:3P)WI,aO(:5IVRESK41B4N]f#U8<KM+Xc>
d[0b[b;@bJf7C/WW&.\1W+5;6aT]\FV__PDEX6e7#.2HU]=DV,^&2U^W9);W_]_3
Yg&BSU>(28Q:2?)A7.6RT8X_2,;+(]=:VNKTcA5V\3T.NC.-A^[WVe8J9I?NQQV2
OKRAN<Ob3ZSH\Z][d\DgED4bfNPU]8##Y5SD04J41&(L1R13&6McTMDN388cd8NT
d\-F,A)<2+T(N(?W\/=3XL^V;2L]11BIT;+:]NcB5+7:BU2LTgIWJU&@GA;T<(ST
]IVT,+^>?Q2/D3d@E>:,BA22J^0cf->,65Z\B8(H0Y;.XLG[=(3)G^3-11):;Wg2
Y:QKCXY<.WH?9<S^0WW>(L_]2SD/=e:#YL?8F\.N=Y(D]<BDa=dcG01FPHK9Rd4+
\#1JNe4HG7OWZCE(1:0)KFbdaf?M8E[1SRE5-A-Wb6I=.Y5Je600#))8/#</AAbS
GC4:AY7)O>.PZ5D]N.OIU&O4CGcHd(6Y8@]44;HN\C#gS[^[>GTEVgIC=?[4ge78
EcF6)D#+F(H8J\D?0eL.PZC7J\J\/_Wd&TJ,4^F/W(^[3Q+CGEV0)^<7d?K/=D][
X02(?S=HFB7JcYXJC\MCceXc]-#4A2#-eSHTa.9MKO6IF(>MHTQBJK)R4^5ga&A+
=N7L21CR6\@46#6)?NXM0^\K[NU+a2E[J[J6<+0WE)467CW3>/c544(7-=IcKVWe
4.^QXQJ6B;HY;38PFZO@1LW\QHgX@J=DPc&XBQ1]@PIY)<L\/KLW7U^F??GgEPGY
,]Tf+5/B4N=-@3:aXBL1XZcgG4dA>(R(29g8<1gNJ1[60XGaV0>+NBcVY-_d:#<S
SCf&8X2@+@1=4N2=^8Se5S3KU^#\F2O7635B&CFg\X[VLFWGSE=gLFb4Y@RV6.@[
M8:Igg7OVZ\H4OQ1@>TZF-Q4QcYC42<B]f\f@RI5TD,@@#4Ug>3P[eBPNI?M0_c/
W6><&;#[TZNPU&081/=J_QQC-0d]f=Z=P0T04YPE4X&LIX\3/.TW(f,R@GdIZe)b
2-<O[L\R>L&YK&bRe<)/7[X]5-1bZ#1.;cLfY\ZG?DdbD,M5OUCfL9(O(D/e-/c;
X]M&ad]^7?O9Y:/OH8Wb(J56?-6#/@R[9,.<_cM?7^9.A^GGE8.W]^be<Jc7DSG_
IBAOB.4-e7^C\e+4Z.T]@4QH0<I(Z-/.A0L#8Acf8&2A?DSP3b50Nd-E&P;_\=&P
#g->1K^,+7]-US3=T<,W)5<-JS@J&2LaKN5ALI?BE1[E:>)F1]_-I[<+QXf]YRc&
M7?e.^Zc:@Yb8Y/ERP:(MEL1Bd[26.G@2^K897O,VIe<?ZMR58Pc)=@77:-G4U@(
<g:+dAOWLD.g^&d+93C&f=BT)Ge@:WY=<b=Fc3+7TO?7;CZ9&48-[@a;bM7&OLeM
?Xac0cEG/II-.\,HK.WSe5@+_/f&)F:cfaW,/F-KeC^&NB@PS\_gJ6=Ifa_aa?W0
.BOQfe_BU>Q3fYF>7+K6gP?JK;a1BBR3M;IG[HGgPb:8JY=82+6D1TIOVIZf.ZTP
5#8g9G\-1X^39ReAO_F8]Ga2E=>DHZ1-6P1CMbCa/X3R56]GYR-<-JHF_dYCHg:W
LbSfRCcZd./6)P;^^E@DV=8J97b>J(A;OPK>Pf104(LCdZEV@@909+)\BKgS7&25
]:^<[^2&-[3#:>^IBgH0(DeVOKO)(37T\ZWZ4Pf=AF/WdZ4Z>.B6OFJg-N^=K&()
1g3=<Q6C_P_70ZNO&9]HE(]@bAG&Q>@/3\Y:Pe@0a0?V=a):4BI+YSaSU8:(f:af
R&6C<DeU24AR_;cR^f8,Uc/]-8VT6?Ie><LEQbKCP3Z6eO+b=6BUZ?b)E:f<14E?
KfFF5Ef@G=S0<,X8-S37<\^BPaA_#Mb;A:gSH4K8:?M&[H06&1[.^)=-b7.K4g>-
_KB=_RV93C_HT?@H9^VW^Y-K:NIYWO6:5G3<)gNW8D;KR6\DBgK<E-Ab35H&5MHc
Kc0eQL]W,=3G=FAMA[QdQe?FIWeeD,TG+A[C(&NgX0f</XNP@:gJg]X9@KfH1GOC
)C^PPeVId2+BZ0=+C\HM)&NDAN0XH3bH^+cXe;O]H(8)?2NZ82O#.6I(W<WK,-P]
?TN&A9]ZbJ+M7L.F@7HT?(_.)=3HPNQg1dK[54g3Y9cR_N43cf4;1,AY_f2SM@5e
_5)H:(W>Ye4ET]R6f9U:MI&YIX;RPIa]_VZER4>TM?MTP-[e1]GadW##UTeb5)E2
c\/59\B7:@7MRf^FV12eZ&e1:6Q.aK:f7;Q37&O#f8<]46eTZ;@Nf5/YY/KHJ?YA
2ZORQR8&U^4[)3^4^Tbfc+W-JdUY?IRI>:dH84-V7b=AD4V\db0.VOW0^=KGaVKG
HcC3D87g02[\9fT2;8S@LRW)@K+Gg8^a4Z]Q<_9T8\EG;36Kd@9[A6eNVAHEVH4:
;+CHW(.FS.dO,IEAGLR2b_1g]7DF[6O2MfNZDgI7G&.BSPf0[,^HL,B;f/\EH3TL
:UaLc#gW6+7#-_#_LBfM(EY8@W.&W[W[^6UF3BZ9YX;:J9GD.9Vc6;fM^INcCK0:
;N#cI8T<Ua+;<TaBO.RQ]US\G+b-Ja^:K^UVEJ/Q.=B?-d;[L+P]SM2bg2;[]1C1
\[eP,S,0/DQ@e;X-LC\)(G.L32A9db?AYPWeA,\@WeB8AE&f-OD79LPaM@eBDe.-
>90\D+/WX(&.&YV^=A6TK[,e6P@0>+_82gYb&=YM/_De4]E/KA7G7#W,KYb8O>0(
@dcacPH#J36BOM5\@24ScXIdNf76T9b8W<)?_?T)7,DU_6DZg^^-UD0_g(V\eJH(
>+e&M3A-:R?[9;]/FbOZ^_+.:?(Za;E0?/95e>E,R0PXURZ5NU(72,ZB(G5fZ,A5
M5IZ^EP_dXdf<eKSLMD39aWdN<9E,@g_XHZ:?^.+ZQ0(d@4]MW7D->M#B0V+(B81
5;SS&/aZW.R.gSMbN0[[g/&FR<[D[;OdA[[cJ/LHG,ePEV=P-<I<//fDM?8QS(7P
J_J=3a+g@P4<DdNV70E0_U:VDN0J_)6.Uf;0DbJ+L&QU>M9E<P;9&c=A7-:05.M8
Iaa-]/bOVS?5GN1(WDT&8F4G5OB7]KMX4c:#]XRF+<Kece5(^T:>@XP72C_.YNSM
^GPELM(+_#Mc,@7593L8@NE32S?POd0TBcT?5/=I-d/W[C_RX9YQgTf8.\9)ec(>
51NbV72\+(BQP>[ade@X7MA8:Od(K@ZVSR-D+<]7J_,[&RKR]<6A:/g=\IIddS[O
(A-=92YbE]-Qb\>cEF6).U>9K\^K2@[E=4S8ZHSdH6=K(V5cZd:6X\c;He+>&:)4
be4JLR-R:945Y_aELC8;M?XcBOSN3K,;(JU.VI2EUI1^+bMYS;@D/&GF_Z&=I)D0
&CaHZO-BF3JY.a0dV6Z2HR,[C+?BU1BT\CZT&Kc^\@T71_4J87HbHNPcGc(UbZ\B
\<:\@gF?A_9(b,/Z75JBU1C1,VGNa>33@LA61c;eT7g67GI98XeF<f)3I8Mb32_L
3g<ReM9Q#3S?=__)^MV:8D-SDGPg,[.\0IFD2.DMM1Wb274V8/M<f56(g^,ZYC,J
D)[3g1G&dF_GV:D4N/ZMB&\N<VKeR_@O18G&-@^P]CMaL3==fSMZU/,X=)G6Q8&J
cV3R-XFLX@=KC]_TF0(LOR12O;T7SAGU\OCH/eOO=:;)0E1I:>U@(_2?KgL]OV]7
V:eI.EKe->TX)5f;F;+e8cG/0)#3YFJ=L/=F(FWdBPK6g803.295NK#RFM@a^@HP
.C5g9>I<<L[CIORf?ZEa3N^9>L(]2.R4Abeg[EfOYJ:F:NR/7HD7CJVUB<0/9HRU
<8XdZg0K;5(V_&DH>+DH-F+)@YQCLA-ZV?g)EGOAMC,X+Fa0\=8Mb0G4)EgHJ_H-
L^3?eTJ7_PC):b2(S(IZPID^3)R6.Q>-\4a.MIgDBJO8T47B;&7AQSB26G\_0K?[
&M8-A^BE635YS9.,VI_VX44ef[D8:.8aND0X#RGF+9U]BSRH?FNP)@9<N[,HIQRf
2Lc)G2R;f-7SDcD>CA3+X8KNHL+ONRIJTR0eK1HGgK/YKaCY^c,NOYS5IaaYY01A
S#^/^P=F\L_d3&N#O^E6MY.LT7A[MKaUJ(MLPT:6f43:O0Z04P0ZgQ#gYE\aPMRg
4VW5P3Y->b7-)OD_4E1;HO/Id/;#F)R[TK=E]Md&;]K((4F2fdfS&I7:^AY6F2de
2/?P[E/f5g6ceC/_L>HUZ9GO:(^-dY5R7Jb7>c<.TKZ]/&AR7+c^+eT#??,4OA5<
;)O?[=I@)G1EQ,MgM(MR;e6SFJPQD7QKeLg:UT8A=-G)SAe6)[O^>F,)EVc7HfbG
@Qb3E?F@86[.?=)DBE\_Lc,6BW5d(>1V(D?YVFUW8eX4<8AVQEIEI92eFcBGRD[N
H8AK(8d>B7.XR^D1X_6E1[X/)#8UaN@H@+K1g<I^68Z28FHa,X>W0[eeGK0.8H?D
cfS>K]30)],##LPP[NSTCLa?@gHGe/[A=d5Q97SQ&L,bFZ?&Z.eDZ7;WV4[BTOP4
=2OOAM[.[gY0VE#8f.]#K=cFd8gN\<(=D_[(T/SH80[3?UbQe5M&U#.-8G2LbA95
#25]YBP41HUXSBI6R=U(.Y6.0ODK&[B7LR]8@LJ(G.]@bA_,@&_D;Z9IeZbWbWCK
<\RNcX6Q&RDg<D(>4(>XKAO5]aHAKJ=_PVE,JK4(Y7bXe9^H<3eZYESY,CE;MV-A
U9.=?G<0(?Q[X8Z<2(-)f7@9(O3@E:FC;-;^[[_aN_/)&O_3NfX3CB8ISNYK0IeT
M08BWgE&f1F)-+c7-4Q?##1d+3[fJ/CW(Y5Bb+NA(0;TaeRMU[<7^aUOdW_L;D7[
,2E-&f,K>D>5;+X1.Z:e,V=Z4:D>EK[)AQ_R@[;=</FHI.3VS?V.MS_KQ1+1EWSX
6WNY=[UDG14S,GbC+<U5f>.F/8&+NYW@D,@Z5<JST5>Rb0_^\/PV=d3[]S]\&7@S
J2Sb2)(5Lb6HD]Jc4d:f]0R.gHc:O22X-?0V8\5NZEb)#+bHR:##L2O1R#U^N(<M
O0+-F.Id8CAg^Ff^X>+NG(4X_=V)Dd9M-Q(7fPJ2QNL^)KRA_-AZ,Y5@gV,GX@E8
2;2ZDF,R9b0^D2A\9/-785cE0:AeX^;bZ:AM&V]N)(YABR]#L]M<81f2ZR/?+eNU
T.;?=C/;1A^T-R,NA@a;e-/70/3FLT@HR4cK<c(b[@[&XU3P.>f>(ABgU3eI^FO3
L\/V1Y/0Sc+634eDPDNQ?[,>Seg)f5)aK2G(?XH^O,T&\RM2\D]79fEeEg9PN;90
eZ>E3ZMaM6N,ZNKUPYRG>K^YT;:e=VM^]1]dZY[>S=dGRFU\W+T#E?QEZ.eHC>K_
DND-P[1(MPa76?Z]E,,M:3#6+><LRA]7d&9gVN3NMIcZ^#L+9.c^gD1D;T#WE<KF
IH>0Wd;N[YUUeCQR[^UL/0T04PJCEbY=.eY<SA)Ce;PVN4GKKXbfMb1NA2MAH;OW
5N65\/-Ic.3cVF<+-9_0A0BDXYI(0B0SM,\#I/>H@.7KYYPS(Ic[TKP5J,caNf[T
@c?QRH;DZA(19]/4a/dN;866T^8Y>4@25Z.Q9-@^[P(I<&9)XM=HTg5b)X2Ob#BJ
3+BVU)gK[LZHWSTTF/RUEUDQUPLO@I,3:f^#^57b_53\#?d+L]7N9ER[^=[f0(Z7
MYINT]cYWTOI:RFYV2Bc.c+.OB39La0.T(W#HfTHEJNO?+K&SX,MX[?e3G?T@#A/
BH]/S\-UZEJTX[-P<5F79X3<)db8LD[bF4I,+C:Z1OBaCYV>/6KO:BT12;B_[Wdg
H9ALaB<RXT[=_dA5RfCYFW=:.-e\+NUU6b^>O(WL^f@2^BWg@Y0ZDP-DGd#.]Y4]
,:b?DDY-ANRg4:VPU[[0F2.Y6FX(7.a]K5G=Y\,/=bV]OR=7-[NORbR8WCLIeDCd
.Kc40_Q_X0bD9,TC7g7OITG<\.V,Q[E<B^#);X[73>P&HB(ZYPIPLV_YE1M4Y.;T
P^gFNbKQ2F8(JOT^1NEC&EKaf3WG2J(+DOHe=\MgK4[=6]eUGcefTa,P@RD7\?VO
4<SW-KLCc,c&6.&fH[Z_CFc-N08,6W+P7<-U>b,2<FH:g2C9/cJ#XTJ^_5a@g;QU
fOKe0I]LAN)X_A(5?.INZ2XfZL,IUS[f>.\7F9DK;H,TEF]2C#BMB:(VfXF.c=Id
:D?W0+I]V6GgV?6G_+HBK-NS0;JRbIPf_NW>9<A:CXeZc@6@IT:>Ofd0?,\DIN#R
NQTK3S,:SXZR(N#P-YBI1WFS=/3:GMM.J@2)a@[T>d(W[0;e#Sc3\@UBNA:D=V7+
I+LBYXNd48@=Hc3Fa[#C1f@DTU6-fRI\1:D^g9P1GI)9MA/A&79MeD0AHT5(@ggR
H0[D;J@WN6A,V)SYF:e1_FGH;7N\B>;R)gZ7B\AWWWX,EOaR>QaccB9gG3;3@gA-
adg_#\]0aZ@N)VZ8?9_I=V]?]9QUVa.]+0Z\1>:(&A1RVE9DVM@&5+>-FB_&M/L6
OU1P/HfS+2UBF;)@^J;+bA==9@;H.5BPWX+C^V63T@G_</dE>]F[)E9R26DR\:gQ
1+O/-CV78JVH5I5a/HSfV1ScegZO9^\=)UbY+&7HC=3](cB]-[A,NB+KJ<N.HP\c
KgTBBc9#(aL.>2cD&RJ+R],g\A^&RXPJeebRgL#NYA71fT@G7Y<EI?f9@F,^?(KA
GA?Y/2<TH<E5c@(,_RUVS9DM+2gGPa?_2gdSKf-,V8T(+=X/5ZR\#_4Pc]474DRc
#g(WG.FdWD]=#GL,@2]1(QY,WXgVg&34\AHRWC7(e5JE\^TaSI34/\;f?A1^V(b^
(3#P]-()bff#U8D7Gbcdg2.MMF&D9b&G4R[_PXMdB5#;U([[-e=@\EN=F4cL>E:Z
9YV,Y#\YfFV9gOU4+f_I]S4866,-BA-J-,BIW2==4HaL[GbLXf5aZ<GN\GUd=J@F
1/B?He)^7(ga8)(B7B(b^_18C7VH7O;J-N_gJQ(Zb,IXgZTL@2;OACY0b275C)]<
5V@f1T#HIJ9CPCV>>89[_)C,B\_6K8:AOYI5+D4XW.QH3bINB7(8[]BFIU[.Q)a]
g0U/23;T(_aU9B?MV&7c7b4N]8=FTV;G;PF7(_2X_M#@;TZTH6^K/c5]\/cE\@.>
P=K<C/46g+Kd6K^^e2:TfO&3S)T]W^e#\NZOVT)LU/);^H;@BEQ6PLK>fPGY#S,;
I7B\.7P&3_JK)URJHS,3)bbIAPJ\TE1bMc@>UI@6aMKPYW2OD0ULR_)=,^]M<=6U
[#+:HAF\]^V_S:9gF;I&)9^0#@=1CFMMU?+LO@M.:?/?H,SY1OP4782W\fB@3[ca
d+FJMC^Kc.M7JfR)3cD[V+FE1gX1;^L7/8Tg3N7_L)ZeX,WZ9E1,<e@-_5Kb_@R0
)>LeS7\/8CXE0.S1V<3fUNX2/TP@LHR<a4ZCgE+;e@J5-3O>ID7]TWNT_[+,XOSb
JZ+f/WGZ)K06J4#bDL].0RKL^cK)1E:A4]I?g5=CVeRB83&__QDFNH=G[KYa4bd?
\LL^cAgf1ceaO:fC<<J/9[LgP6^2T6:Je#YT6[[>+J5(V[4_URA&ZJ#5Z-C=C#YD
X\:QT62>^?;4/H:<^;:T4dYCC_JF,>NQYcZO]P+/I2.OAIb:BFY2/4?<K.3e)G5(
N+-G8fDOE3@KP96G\^Eb6(0#-Rg<H2I]e8:C2Y^]..AOWVaC_K47Mc7RfIeRf7<E
#O)T,5=BYe<Vf7[Q>WG]f,A.H7Q<g<4)MK///&R35e]URcd15<#-3cJ?gAg+a+U[
8F]DdZDPY.XL0TM]MF8V_&3c)UMY?DP0]A1NE?JW_\V/BaI+7e=6M4gJ-AYLEX[L
\7e:)Z0.8SB.E4g<EGe]9\6NcY8H+L_RFL/XeBC7<56-E^a[dP_X?AUSN\_<&I;B
;H;&:P2WUZeFOX<f6DFXHZT#></9^L1EJO=AbU+TD)?+T[\EMX;H./<QNdQN<;e)
d,5LB.2/f(RH=2NDPC:.)363,VU#PGgW,69CW46T]?L<NHAA+7D,M8GDQSMAA6;;
OB,2@P(+,9<aQ)849f0D]1;K<@?O:eUY[((+SE=UgL-bE\KX=&TEge@@^Y.,ed<X
LAD-3O#CX2\&aI]a>ag0Z@SEbaSAcU.,9YR4dIa:.(8C,d&5S,bU:e;gY;[SUD:G
+->Q\bFVd:;ZPNL:.)LT<89IAI,f23&E[HYH/P6(DW#geSJH3:=@>)7^6U=U^M=U
&RIV#Y4UfBSA#_?5b\3XB@e+\#)g)0H3IUV(=M-HN4.Gb)#KD&Bc59GYL@aNLUO]
[HLaMa=HA8_f=46VO&>-[KN_g]NB,SCQ>>7#:4NEgcUTbE4gbL(&[.7A[Reb@GSa
-)KYUf,aWd0ZZ+LLJXB[H4RD8MWUH;78Bc=].0A;F=,OF>ERH74+b&gO(TK7ZcYV
F7fU-XDJWOQ^;_4S+FEP1F</f](Y]Wd1=RUKX[:=)a<J6+41+R]0F[^>,FQ;c&K5
W<,:13gJT908ML&SR_Q]XJ.RgQL0Af>F\4TSX,B#7MT?OYK2d1M[8D)K3+Rg=(/4
AC0B0[OBVNgB94-Y1CR).E0K:6N9P[4aQ[T0L([1\\IS9e?60[>WD40Rd@)PDY0S
NNcZ9(RQYge@6BJMDe5KWNAVMLL0Rc/=gb]G@A6\R80eQbbC2[SRF9e+Xaf-M^^d
c18).b=O?KYH;BQ=8JP9W>R_H3DPbeSBb7@6LTT0?E5RT1?O<MTVHO[>L94O5QAL
]0ETUZ)L>^efEVMec/(0GNZJ&NH\>RfU,bbbJ=9Ee77E-R>(aQMe:+]:</a_-P3\
U5IEOTc7dB58IV\=@)J++<cYWW63&AR:J8e.B^IfZVHD[]F:eANH6C=(J^&X=7/<
^3184f4Q0OKLP/7,@H?e<2R#9a)g<P&J.B,:1:6,2:7(5/A;DK1]+O<L/GgDe/f]
._Na84WF7/M@R&JgKDge-WeN3ZOfdS]7YQ+EEDY3RCI/_@J[CSVD5>-RGSI4-/C8
3M,Ue48;)aX2=,@fY;4P=PRb+,VBMEH).3^L6ZWe->V?1GII^9,>]TBH/Fe[:0db
UJWXCR:GD;+X)13KNf/6B_QRUDHN>LO0,=(9/dV^H245&A8;>U0=QTWbO#5Z.bBC
5^^1DSD+A9C()gAd5J4]+4/#.^2G>T?@+SQ&#=bX8D)L&/P?6a:e[>_W@N]CGTFH
S?cP59SF>Q1:@<<Q,bPX@^9dRJ^9<+(g/[UJaU..H7:<B13fE/PO-F@19[&.^eF8
;fRXe4<_;>fS.0/\=]>aTJL=7TTJ/++XX6H[>U#I)IQ[:];/9e@AYW<LNb^e_V90
IC_KM)JTBZQC7CWNW&L8>eA#9&.5S::#7,H5B,#3bROME2S+Q^1KVA]4b)1NHb;Y
c760T0Fe4DA#8/_bYRcK02EAE?T]5XgI?9N#HBc/AD2V<0&BYf?SG+(cJPMUIBG.
bN#@Q5U+^)+Y,Y0+UG_1Ma_ff5?D+)[gT&=JVYeB+(0D9KPOB2^BKX>I0(W:Ef]P
12/YHL(6VFc2UU+F\?Me0C,C1)+GTI+7Z9>R;5J>(<-aCJC6eTX\YbGZ3RE4412F
?\?>7YeJa@FYAb491c6H;S,2L\U0f..5)<9WX7OO[LbWT/30^OE?^b^>0@f<L@(_
W)40P,]#N+TN4KMHS2&,<C]f02#)O8M\\V<?)H[FE^G>O9&&WVg9AH=&I7g2#:fG
NX#cc-c&eC6Q&KMN^.UI-YHN_ZA5WHS01YQ3:<#1BBFfD)\ECa#WRQI.).ZV6VY<
YOa5S9Ig6fcM:QZbIAQ7).L^NNU(ReUb1=R1R2T4eF)dKD[<S0TLR+OZ8aB;HcaC
:J=^;Wf(0^2RFT4)^5[X@c<g&\R3=:ADTF)AcPAI^#6adKBT45?gNB7;DQ^LCg(9
@B3HW7CP5FY[X(0gdP&Mb&S@Q8Jb,/Qd1dY4/>]+,dBIESFF\RB;@HN)>TC2GE-+
&CCL2NNH&8,,b<Yde?aBEc-6R3HbSee__=\T\(=cBGBde,HIN4Y<FPL.X4#(I-JW
#)08GB<O4gP>WAfJ15NJO-/0ZPF9HFV).=PEd\PF0.f>=f9#]4Q[?:ab_?2bI5U.
46d5=CfgYGP05&DdMD]Y.;=>X;5FTR4d/M1C^SF/\(0<E)O+cR:Qa6[6<=H#g?IY
<g391F4N6=-UF<XfY(\A?3NVEBW^O<L;=<B;dHCAJ\Q3507D-DOH[UR(Q3);=Z9I
-/V\9SC.3JV+f6:Q_0>L_PB.3f<;C&W(CTHeePWA:&?1SgEPO6T?C&QGFV6,g;DV
FWIMbK)f2b[T_bZLXLd55=<I+;XX4S8e,CLUI8X]]N51f6?(18XIG[Id:1fF?/da
FaAF3M&952W\<6?;-3?,g@MK:H/FYN<-A.Pe3,UZ6L;gN&-AgYYB+VY61M4?S_aH
&Pb?cW4fY?ON7EF9@#dO@U37.;,W[_VGd7.TfW9B<\#I?8c8A#G\e/V/3OMTP;N>
:K4=YZI+b[\.\I:HB4W-JRW-=>8KZ#2-JE0VO(=HVSB&RN58/?:Y#:G3BG#_gM2d
8_@ga/cUDR6@#@C;JQ>0M4D2/PN#TN4O#M.50M4=&U^e(cIYda_d?+7V)N?69K:0
#gX=DJ_TZbDcFR^WKUScV5PJ^^(<L]&PWEN[U<e4?bAc^_Le&\f\XIBU0DR(O5eC
U=V/KF/#Z,796#T@[Z6B8/17V(]?FMLVD;@c[PJ<6AI5LS?ACL\;2__X_1e/K98I
?@;&7PQ?7egbD:IH3b]T63@Z;W&9Y(9)UV/QP@X#V@@<U^L[8C&c11(c.4I:F/eE
]T,:N=#Fb#/KbL4(BVZ;(Z1P5/3P[9;YW)2:M4&(TV;\1-^\-@f:E\cM.AFa92fA
=C-OP:-KRJ\_;LBYG#74U,257eE^7.O/+@MM(9#OM6b20b(OR;4R2AY<d.g:\cYD
I]LTZ;^fQX7HM,aP6eCF?)EL8N;8^X>G>V9=+3-0D1RQ+f;163Peg2J:A+/g#(F9
Ra7?a7aAe-^S_NU&>&UV5]R.^bYg3Q>LK:.87]JX<cF)<,KE@GVC0ca__g5MA8cL
W-(^H,FFY1SJUQX>\HX)faIIV6JMNS8/Bb1b-EeVZ,2MD:K#1>:GH:I1eY<UdJ8@
:MTC^V_GOafL.V[JZ?DdReeG/I/Q-27J>)62TUPI?_;9=7^X80R;,+;)aAaGS>CN
3LU1A).[FM\Z53[.1IN=G1IV_5+_FTf.0=+@E)/8KbCFc=VP#(?@FKIdJ<AD/K?C
aUNKF>3.51e8H>RLJNJ_A627WA&?42B1De]-MP^RdM=1[E;ec[0/-KRU8fB1\a3.
S>XT/OP9L^dJGO>,B<+.,5D)]5dUHL\2.f@J95-NYXfc0==I,+R@([e,Q\JD26^N
RdTP<\K;(._:;(E=eOZ&KAKd61Qg-,1/&RcfN0f+4>HD_6;<54J_c.e=&f@A]7XS
5Y,9Z8KRP(WE9CY,aZP?60(b=[Va]>U;WWIc<Y:.(QVWFNGWQcG-#XJ.fH\IOUPH
g9_F(FC07[K>K,eaQ.6]Z-?X?FF=/862>bG4LX#IE/OLIRF#bQMW.4eCbOUQ:RN;
,PQN<=/SUAR=?6#M#2@ZD6d_M76E7(Mf]Hf6)6FH05cD+Ka>a3&D]-1J<_aK9Y<Q
[Vf&8Bf7#_bR6=a)W,+6H4SN@D2_[+18Z?G^(53T-ZRT+cVb8;bZA-[g.45=TAXc
dVD+>f0)EK1#IWU:.?/F(-_Y(e\DJGP6DDa/+ZaZA3B8FK.,M1?ULQT]1QTP&5Ab
7FL._EI_Oe1+(EUUNb9Q[PKeA),LM=64#L08bDd.9L4gU/+>3CYNZ]YS]>Q3)RUG
=;0XVdf;:KEgOEB+4GgfZ54F&7.2OAga0@S4DMEPL.0WNPHdCW=dbZ.F/8N]\6[6
DWWPK03,D(:+<@aAdeG)Jae[SOE.4#Qd>A2R^g;_@@BZN:_=5&>:BSSCQDUgHZH[
aKR#COU_N>JeZAD?_B4&d2\^9EQOSIH](c#0bEF#]-T):^^C4A,4dKUYKb-AY+Q5
_TB#7Z&cGZ67c0F>@c@=#>)>#GLDE1a8M)a?5]205:<ALLceN)[CXC;HcS(?=&6-
T[=4NVL\c(8J?Ab1UDBD6A(+E\ZBLaC,@/4#5/MMU_WXU\_7OT4EaWb2(N:/Q>-P
1>bR[O+5H(LBPFH_X,g0\Qb&SC+G/1^,<Tb4<]DeYF8,&1-KObG5D##-ecV0f,XZ
DV53>5C=R3faY,L>b,3H90VGMJ?./+UcZUWIcMbTf@=+OY72MAfCg=4ZKe1cL?-=
VB9[&#8RcYF^+b#a:OF:C36R5fYHV>/<+_<JfJ?X+JIfC_?2dE5:AGgQ+?_(C^D6
LX\@3=D1A:SN3a1PP7U8HcJ9WIWX@03(6JKPF9+-\G.\P2-geX/YHB3/e:52M?L&
/)=6-.F<JFgQ3-Gce0=W_D10BIOQc>)e;,FHFeWBCc(LeY/&R<I_c7X\21_[OdEJ
SBOU@fU:<<&;]7ZMOUb#7LFFMVYML<SX=<N_7]A(T@aXZS>2e;@Gd5ZY^GL.@ZaI
g11&]]Q?GNC<Kb@.B\AFGB-/\QEL+@+\aUEH3J>Z:F<=9=@e0>Ddf224=V2fZGb:
TVSg:UOV#?4O&_Ea@UZ2AceDBW5+0>^NDP7=?OgZ]JB<6gI8OS<:R2;ZCW>2O4?7
9<9]6P](/eW[B9CGX<3#]LT_G]Y)/5,?Fb[SVDM,/4[5g?4)6K@YRXBTeJRR/Z6a
Og05=O?)97fINd_6LDJAN136^(TQ&VU4&IUgFH07<CIF3XDWU.0cD@Y>-.C:7>:]
Y?#Pb4WdebOLBW^)L;cN(,NG&W\99^+\CcV\H/Ma@YS?2<U+X(^003/4T_O:\EJ#
)a9b3R)#J<2S;LUb8RHBD3aDFTEQ_SA=#7(.V&@XQ^O7<[L#@T><=@2(Bfe2),fD
XJ@Ib?K]YbH?6WEYf/??CGeWIY:V<a-3]ZNDQ2T\38P?)cR95IDAffIbXUS+8A7W
I1TBW;MV:-,a2cG+]VRL8TZ0JaeIP7M:?)I><<e>^L>#MO9ObPYcWdJE7>H41AcM
_O\=WZ73)/<6_\dF9X9)RWd+D5^&8U?-0AQHCA_?D&BLVb^e/aFXHKg-AM]bZf0;
:#N-2O))I]]-&TKIcR_[^PF3?IW4-?^d11GLDOF8Ya8>_QU6UL)/44APRAJF(S7>
UBUV0ZGA<W:SgJ.U<(<ICQU64]-5I]AFBY0>,)HgEDEX(/X3AX/V-2T/&F.WS0\]
S2g/]c>\P3>\WbK.L0fUAU?-6A@64gUHM#f3K^//NO_/ABK:Rg=;IO4<,=@RNTL#
V=;Hd..R>X<VZE]&J&T,N,T&dAZ02a.NaU8a.2<fWGaB@1:X>DT3#(B?f);A)U0K
ES0/BN8Ma&?LI<#WAYY_BaW1+LEH#.<)\4eH1=eX:=e,@b@2/-K?2#1ca/H#cgQG
g-E<Fa?YPB)1V1S7Yb=ZHH)5--Wcb96YfHeGL8]2T_/_.==dfPg(D0KVAaMgD3TK
T;S/^Z#X:PR#/_&&8JMG<@VF_FIH/;4Ca3#O&S15dY0ZO8cO]IK]+MU#^^8f_3&M
CG5L:dIf_cdLW2G./D4)800<-6Y7N(/,C_LT>9VESRe/#YC;Yf(73bNQ,)3]fB=F
23/_)<9I&=K4?18/URW&UMSP<c#GdN1gMg:8NP[G2-D-Y>QFH/5HALO=EUZ5ESdN
g&TH16G51g_YA^F^[;#5&C4T0(,)0:)Nb_7D#ZXQ]X5^#JXbSa;<3M)&6#cKN1G(
=3TW^MRKG3eD1be;4-5K6RBX)>Ud.Z5df](WB2+FE_FDE;&4WgJ#gKF[UGZ4bS@_
NIdbWSeQ8=V/:;+07124]N-8JKcDC65W:S-SQ_WJ?)[8=],/(7>>CR@3@V6(>dHT
(8=SCU:+^<IQffI9gPT_LYaRIe7bfZD8,9.VZG#R1E38@c=<-9G9+W>NU[fF]1?N
Z75[QFTOX)FS[(MTOcC#YA9AWY]MCBP[-[6_g<f[[a-R4U@?=@;bPbD0Ef2/XZF+
I[OZ#GD3WgAGEACgaa,Fgf8?F-L;>2R=BJAF/(E=5-bLS+8DaC^=?:3B85,@3#6#
FVe=Da]_CS&6/g4_IVA:=K)3JW(cWE5RH80-+:5L/I5>W4],&c\QTM/6ONFIP&D:
;Xd8SO_P&Df)U=TBCX.Q4(8dD4I.P/URb]Q.6gecd&c.UFP.R),=X,bIbIY48>UT
SbYM8g<BaF2-b)&C_?If8/g6K?LOH(Rbf0Ga]J+PG#S+)HbY-L-c[0\b_RJW3g2R
#Ac5Tc7:cKgTZT[-SU<+Vb#E#6:.Z<+?C.&K2;Q)LaS2?]WHP:Ha]MNP<JB.c&LZ
C);bZ9e>.M<O<A4G._E.TD\g)M]DE]J9(SJSQf_E\AJ3NI=1WHbSHO226L1?3gW5
-6g(B8X0-Q.M9IZG(M6XH#K;NPVWPY07_BIUcLJ3=#0Fae]N9,L^E3[,(g6c@QUN
F;=e^ME5eCfAGgcU9Y@D(YSA2g+,4[5?eGb+J2dV>4G=.[]<BdB.>a1f/)Y/KZY2
7#2CIH:5#HB-WO)F4eWWDac.T5<;C\1@^MR2C<7(FY]S<CAIL_UT7YRNW:L;X[Eg
2ID6?AO^Lc,7<;c2:R=QK?9&@@D#;8JDDfZ3WHG,)F]_#0H4W:]6EQCa6C7Mc_C=
AadKJdV#cIA34PJZFENO57L830aeRV4>G-fGIB,OR]I11-Q[3JV;/RbM+1SJ],df
SD+Y]=EH7R+]I?L.c_]C1+1[J6;QC[J]#U#0/PYG2(9b2>+S1OL^U;G@?^Hd)PWM
.#7f8Y:]+)C/.c6G?BDOFYb;D(=OJCG^F\R09QfYdaL)L:>,LH2:DY1X8)D65U[<
aP01V[B_>eggTDC3^0/7dOXCQ;9;Y6V\G=BU?2U(^.@U\=6+3ZY54Sg)>B,e\aQc
V8C5)3IeMGbSdCR1T5f-:U(YW5:2(#5g40=#VUU\31Md8c]5_W&W1.3B0^2Q?A]c
0P-OBNT9E8\XV@EAZcRN@B<^^PYF/N,U&BPJG?+b=AEBb(_R3.Q/,\ba,NZAHHRQ
L>F-GXSS4-a,GNN-39HMgXUE&SKR4Bg_Wc2C]VPD;#C]PD9S&FI?UdY;058=f[AR
)]c89^aT?2SR;&_JLIUYTV;fN9gYePZ(RFT//-DGK0I&0A<cR&S\Y<5/ALP?JXV,
G0Ed[KN>,Y156DJ,3\@Bc_aI4Rb=3g^,28ONADa=U2ZXNW)J]7>_AU8@c4R(=+9M
=@>@)KJ:-OUHJ-\1G/Ge:YJZ9E<<Z>Iag-Y+PcXg#RRY.7eGU;0Q7=/IY(:@:.e#
L(Z\CNb[7^.II#X5eOT]T#b]GO09DT6FIA69P2HNZG:^KV7c=]FM-512fHSGR(Zb
5[):5]0#UV8^)8gZT?>S;>c>TSd),[gSe^]YS:>L1>&6&RZSBd@<;X3,cS;.:4C=
J7XB,ccR9b<gGI^Y?DZ1&eO<>/7O@H2d^6)EP@LWGG^G)&2.N1E1cbAe=1EYR_0C
6R^Cf-ERe^E,0]U+9dTA#?DCbRP1b^I=4&L9BOO@N&e]ZbI>G=Q@--c9Bd<=5=dA
.Me:+(8NGg<f\=S)gFG3;[?9J;#1CSa_RH2:cS1T9_OKS)&O>IS5VX[I>Z^L/]Fc
#fQYeW[79-+YA<a4g0MZJ;,&T_&#6[/^7D3AELSWB@&g;(Ga4AK0bcKHKS^X>;b^
@GX^TKJL3U)a[L++FA1P7,HeERV7gK+@DeDB=K3AUI3cC1IF\4]2#M89K)]K40HG
g(UWAg3@:\D0EL/bGF-CSQ]07<6\?,3]e+=T4Q>GN8@2Ab=[^Rc60CdK-Td&:+8(
Of(1dMNA2b1#D#H?9DebX=-)F@<H9]5(5^W(S^4I,aL;LXLfLY8b0WC27OPD6[Sg
G,S>bA+>M,+ZEKA;N3VfE\f0XGT#OQ&)J2O9=CR^2_Cg0]TfX[S@7).GW5L&D;9#
<LPAKg-2O7JaHd]E=&f.<g#FG^Q1.ZR8/T?adY59),^5L.#7G74RVaPOBSAfO@?f
<fFCG/8=->;PcL.3#&IKI=^b9L13+C.N<#;3405b[96P>]]JH@QJN[7N3#)91(Hd
&ZFSFfYaR[UI5T<-G<;fT0EZ-aXCBU-bF;4Q<=G0KAFE-&)3\Z[WC=/\g38;:f?F
5.:c/b<2ZGY=Ub6/O6VW8@QJ0GG]e5/fg(2&I2?6(<(B7e(,GMR+GUCcRGSEGff(
HL)=EDL]HeF-SY^,?)/UA)^K:a6Nb5K(?b5L&?20I6a&,[N:Z8g[V;DEHcg67a]]
YbU.^3ZX;LJ8-+1X6+e/PX\EJ[a7&Z3b.[Ea+IG=OfSX2FG1a\CddX03/(<G#cdG
C080/3I6X,0>>:L@+U=@_96;,WQ31[XWK+E3g4[K/8=RU7;&VXP(f\g]D+^ULY@O
L=3SJD:78bN[<JLAA5&5A[,0A.P6D2NO[_e.[?Hb>N>NP0R--/Vab4a4_GUL=J,T
TbefaQc9-4?0K_Y8B;-B:Z[gQH[?PE,B^GbcbE>5M#(JLaBTCKG90<fCCG>_WB#7
\<d+2,Ya[VYgY.0#SB,b3SR^Va,YDW2C72C;\/feIXD::878cfX1@?54--S3;fX:
+1OT:]9-f>e4.&P/[MacdUHD4UU@E5dIJ012EO2&:@6S34,85_SU87g?:Lfd&>5H
ME/W(XI=Jf))_GM#RDD+WI0J8c,GK;5W^:5f^eG;G7NbT#e8?XaY:<cM&?F&0\c3
BSS4X&0]AWOK1EM63H<KEgXXa2,^R<KWUAa=_e5W\_WO83+.9R^7>9c#\Qg(8^/I
e;fGJ,1RS:);<-/Xb]Y&e\][CR_7-8KC)=d[&6XZTW(><.?(WF);;RaEc7Q;:7+@
gD,I:UN=fPF,Jf51CPY9M]L1.5JaK.e8Z^PeY4F@JXH7;?G:bGD6cTQFXZ2\G+<H
S@LeH<<7_OX^>NF/:O/>Y6d:)WcKTYFOdb+Q#?0[aY1+CQR5NbH+]&;X]_IV[e:<
9/,fdFE.Pb:SQ_S81VQG@?6eD25<TbO^_>.#Ag@[79)LL]FE1\I-:C-ME[5fADXE
(HOQO.,8aZYC1AK3c0K;-^E,QV0FbFIQ&4C+[eAW^gWLL5:([#&_(96FcfLB_\YC
Waa&Dg6=/e6\(S?,f)ZFPG_dZM2>2AgXQP2&db&]^MPY5/V6_PW=2IIIMFWOaE_X
NcEJ@LL<U)R[Q;HL0M.;SRD:WMVDZW=?S5B2SVfC^D+5[96P5ZeS6fCT[D4FR24^
\d;1<;/ZH:bKS7+-eNGHRE/JL[gM>JZI7N&e=BaXEZGF@Pa7Hb_IRQ+:7Z^O.B=.
3OC;N9:U,3\JacfAI\;(T._Wd.SQ^7+#8<:_T^19FCcAN2.42I2FAeA7((2f6C.g
75fXHY<:MSX&/aK>c,1g@P@?-^[PSYK;WGT?.WVAVeWVb=2WT:Ea072I]BRM4XLc
M)-5=^XfQX[dUeM-16J.8_NLZ1)N-1[0]PWX7]M9-dEOTDC;4S,4IL6.8Z6B,^#F
^c5F6&\<H6YA(][efP=C#(CW?2H>#:S9Q=?Jc4GA>5]QdWE5&OQbbZb917JJ>L@L
OTPP[gE,T\)d#-E7?cJ?JU?Q,_-0PER0ebJR+(/Y#NXcI1>J0]&66S=N+9[Ig8I>
2MRG;(c0VHYY0ff7PdLMdO1:cfN3];G[7MN/9/&b2E6(\RV]>IK\M-N0B<g3I@Od
Q6D6-5Ug29-4]CQR;E&.6H\Ng/V0@C]1)6,:fa=^gFUb)&^+#65LC(&NI]1f.SAb
.ebF,D;eZ[G4c(#Ucd7>>]NC9(.Z123-8ZH0Pe>IF-)E3JCSS:N]d0I+E&55[eF-
3>aZ8bCgAT>N6CH6V?.4<E4R3cIO\UFE:_[g4]E&(_J8MQcU;R9M8U,bbg[/YHCd
72]5>[W=3>CU1<-?_GEISC1Y5W0^GK:;UT#>#=CU;TT67<5JHPb57K[Ge&6MYK>\
J(&CA6DQQaY^Y0/cQ\N#=EScJ3O4_H/09F1GUd413YFK7D(K6\\[eX+_18J<g8Lb
3bU\\_/g5Z:70&V4e2W2@Z<PgfQ;PDLG;OOW=96HZNIMfMX686]NV)A4=ATZF^50
).:UP,NBGC#9]EHI_FP4^ZZ2,TBT1W+W^H+O>8ITE?-#D<^W>9MJ\9WA/d65T4/D
<M+\<IQIQdY6@A@4_fT8GSEL&-Y-aZPGY_I]BM(Ha)LbY0_KYJE&?U#&cc58BCeF
9d04,U+95&@GBW;GXE:Vg+AcVH/TA_KRbZ\F]9.54cGE;ba6bTB2Vb\?A2?=MVM8
[O&(QAXeX<c>ZL#XU_\K;CT6C+2bGHV-RK)I0a)TRV@#f#Z2a]WJe;KEOMa31MR>
J#:NB.MaPM(AKYGR2S-VVB#ZLd(DDVc0CVY,1g/;R/&_52?3ITN6A3FbKTH/CL^b
M-G4T7C30Z7AK>G^\)30\/2/J+^;JI3B9IK=L3X_Ff@H]OI&/>?a\C&+>7I?-T1?
6-fB,e12CR8gU9U5K6T]KF)[bN#ODSWY\_273FJ&cZ2Y<b?9beFZ0O0=>[&=C9(6
N])gG^\GWBQOS_>4gZ<C15M)&SQ;>?)KO(K-2EROZN>&TD=]8,KB3b&&B0;Q3TI.
G/c<+\4eE]7ODV91(W-0gbS1JD6LNRDeT18;\:1[ZLR=V;f)C/5GRE3?YaH/YZF9
CN<CdOLSSFCNeI,FgO3U)P0@GEKT3O^O[7?g=I3&3^g9G^9E\9MOUPX#8+(];3)D
LGKFQ\CTRIQ(@P279\E\A46Ya&&S6Mb\I8SF7[T]1LG6#:K>^GC.TA#C\9;X2DYL
<RFS?V(1Y.7N.J[O&#U&Z&HIQU9.W)L8Q8+>5V@@I#IV\U)MN>a-ST2,O6g:4I37
FU.@;;YDYd2?8N_UF2<K8Jc7/gCeI,CF.Y1JA,4^KB4gOZX0O3M,Z.@@a_)PAALU
7PN9AHIGU<>O8S1<7;OY/WOGTc;>S2IK[,J/QBZ&RSb\aHH)RD]QW_#)_9.?K?gM
_3D;ZNFDJE\aCfR4-[GU02(F\KbPCU#0,4cg4<<SBEBb08#Z\0CO1e0V.NKX0(3N
>O;BKQ8>b8,&f0]/Y2\ZX.OEKXPR]#WKLc=HaS:^<)gedYTV6B_,L7#,_&EZ:5-H
&PV_YJ^-UbC&PWEB)LELOA,=05Zc4=O9#=f?^-P_B3@Nd&M<GH,^8QZRWWN\R>X<
&c6cg5YLeK6>(3&c_#16T-T7H?@bLU7cRA7cK8a^&6Nc))QWV?D#+c\PdA3=f[G#
Q1RSeAN)f0[KDG+dGIF=I;]G9T[[-b(ecS:3L^PLd])g.f)Kb>Bg\AegE0A94:)7
>#a5_S7?VREbJHU\Fd;X-XcP]]D][gK8NF0F&+Bf_R2SNI^WGgD[M>YR+>]4EbdE
-+Y1TXQ4/0SId=O-QGYE)@7<Z>Q.A.LI>NNXb&_RFDX_5,O.]R8>;G3VQ+4/20UK
S-\O3<Cf,1WX6EYG_-Rd\,4?e(\I4aA?[WDcBOPJ9+==.GE[AV3;UD;W5,QaYBd\
3b@@]9T@Zg:@ZGdZ28cNGU21[W<f0L#W^FX:W6H\>>+B2,3^fI65gbKbH1d7UU+a
U83;;/0dV.;L_VC&QFg1:@5WC.((D[Z^:16M?g,J^H1d64U?Q&F\Q.^Y:7L,1Mf+
b:19O&Zgf9HUGI\O=?BFgZ9D6MeYPBgb9Q0YT.)7(Cac2B<8=e>U=4(@-3aNHOLW
&7C+)D-E\Ma=IJIVg:6W[a2fH\acKN;@=:9NS#ZX-D-[T_9O#/N;ZUcJ&RQfK36+
LURIGU+aHRGA5]D.eMX)<GG^cY44-C;_XOIJ.&CMRe>-E<7?55[PZSeCJ0#HJL]>
-DZI13^dY_L])PfKcX),U.D5WU)#)23Z,KQde5WB)aY.^=2MJe)_T(6A&Y:W@WNH
,eS]-;+..WMA:XfKd\;g^+]J&?7CS-=SP?P.PV]4_WE6_GfDZ^e5a(aaXJ=B97ec
O&IOEg9Q0CQKb0\O:-A38e?3TXPD\:N,.Ne?BA[+ebPTRU;X9Z-N=;H3N,5).[P6
9;ZNZaAeA:D(BX\&XLdb6SM7(XPZ2;;:LZ7cLeC>3Md/b&&U,6-Z&L8V&HC8)Lfg
34:PJbQS2aV=G;2D_D^P-@L-MWLS]Xda^D59EUH#dg\<X6ca02.Pc\^4@8&?5HEb
S/>X4B^cDY,YZ153(QdHa1Wd(U^1W.?<V4MNa_V@Xg&gQecM^9_S8KeKB(2<gL^I
fF>WX=//P2YHXIXOT_9<ZTD@]ScT^QV=4NY#Rc?A\)O3^U>D>^;2>M3Ib.cB4eS?
I5IQ)gTW;;]DKWV/@.0Y.;HN[#CH3ZY=MK\;1=X&>7Pb.c)?Y5bA:IX2L&E+0(d^
4aF@Pd]Q)QNW9f=5b_5:R^T^2#2e22dNV6EPd_g/9c^CVe.W1eb&3S/[3b3@(IC4
=ZJ&L&8QebTR=Q?^FWD>J#:?2?Qc^H&L,)6G9K2L(=S5_JYD/LV4&:4dg14GEa9G
7<GJ<@[VF2HT9R06NN21B^AT[;g]P1EJ;S4TT5MYR93CA_[T[>(YfX01Y2-CAHZX
B2eFH[^3]3(9BP)SN^BAGYQ5H[BS)G-<QKAF#)>?@IgPR.X=-D(LVSH1QRJ<[(&(
:2,&&65Y/)56bE)PS5COK6:[=VRM&P#24RA:^NKKYaIZ129H4;M1Wf,:_S[C@W>G
K&9A]K)1US<4I2F/-ZDOSBYI-M;]fRWBbbGLJM[8YePEOX#0\[2O0]B,4>RBH+HP
1EZ&fPdU>YLP@d7_fVXSL0;2.=>_Z7aAQVd]F>23M6LE05:;W./g4;dTNaG\+#1_
TMG]46/Bc,GVf&#KG/-L^T#aXa]L6]L:VG>#Zf5>VdKb&Lf@K?g<>I#21-DD]5-L
BeDIeRZ>b3E:511=#DVI=]WDE0,bB5QA2=[be_&N-N]F:6=c&;+;NN-bH_B/1).&
fA5#PE05g39G^9DMS<1/S_CgYVXVV2NN@2@IE<ADOOAQ84^cGE9G-O0E4fbP##D1
UScM#6T8JTeJK.K)O(L0:E)R3_:]GUdJ>XS<7:P-V/>KL>:OZ;7SMRdX7bYBBD<V
02=7gMQfdI<=@]QA/Q0I_RP^7C.C9E3aY5;F5g<Q_[7[.\Z107a?RPgZ?PE2?N2-
d:BED?4eCgBTJM:PD@,A=6AUSGMG62Z/JZ#<3-U##M0FZ9AE9DKe^^fgb_94)62V
>S\9=]XPF()YeWF(()MZ5\=dSg42,CYINBIFM5]C]#[]B^X>X:DNMFF,JX[;U.D?
:e?1E?YQ#S+GdBA2#->6BS#7^)0QQKS_R(^)E><1_)7G0D]Y;Kb-4,0#X#d-ZIc/
U==<B(=JG9Qa5#:>(1F3HXI7VX>\1>6HB7YXIEGaAR0b=BAg;TT?8b6OGFVY11Zf
_=G=M]6dMaC,bgNL8];^;IQW3;C3BefD21g>SCReR&f\]Z&H(BcC,H3^#N<(?&-?
N-G2/I\cIM<6B_OD9CH<MWIcbSG6)I-TPTL>K8/[<D2DHCeLU:_(W.B;)QJ@XPeM
;]c3ID6;4Q@C2EKUM57WQUFdMCDS\Ie>Xa\<dX)6^<c\LVW^SGWN^_)M92EPa,D\
]1>86d-Y+K6,L;e=3H]Q+BaddHK7=@&;4R;.Lg6H_gdUI5H6\[,3aY6_U1B^N&=c
XCeM:DPIEAJ.=ZbHO_7S54]+&:C^bVH5,eJY-Z#17EK,J2F<eOJ_g2<@4G3eW2G#
1_QX,V\@M&PXXKA54N;<D;T[/9bb\G;2BEPJ8KWJb.28XBAUYMac&)Z&TOLd+),L
<[dW1HaH4A;9NXQ/2LFZFE0;X4HbJ-MDC+HdT>J&DdLLb@=b+aY,NWYBKUURg0#V
+P-cN=QT0,P?;[G>3_dJY::DgS8WG9QeX<57FS#L>:6N^=Z:+?9I]SYf&\=Ke.QR
aUS1NR9OB9O9CNY44PE)X^@BMf.#Y5AVb6I+/KD.X;)5PdF?YDFKB5f2V>14H?Ub
2,Eec+[Y597GT4FX7C1=M#JVF<B\Q0+>^4=FH,g4AP2<B?V/OK6S>C-G\C&dQG5E
Y;5ZSc.3:9JdJFT9)5<PZf/OM.&aIfENQg>#:/MIB[O;RD:&dN8@)=JK&VL=#EF&
6gXQ5P6KZ#Ga,e@PfFWgU?:.KR+.\;7;IJ5E<L(VVQ;/30A#-#^G]5OfdcBECY:G
WY0/2\+EL8c0BZ>0;H3C+297<C@OJf.Q\fK)03N3@(@>28\fGMJeV\7eGd-7H=FE
[NA<A9C,R3WJOS+D#MQEG(T2N0?4I6\U^]@X&NJH[384_=G.]=ee0T3I@:f4KN_E
.(X?.D+Z;>CLYT4&c&6^JBG8?#UOG9dcJWTU&e#bP6:7>;-Q-?)F3KWT2I@VcU6E
eH70b.5b3,?VN7OB)1#,S]-H)MHQY-X-H]LR;?g68F1<X+@T+.G)8=U#Sg=,_V>B
H8dEUFY>6>NMCB90>R6A/Na3W:O;-g.a6;[P8@g)#-@Ng?eH#GD+;_K0/(DE2HJ9
/C9HePV65&9gRDC#^HU:)A8\b=^/6g>VO>P5^3\XHH-14+5Wc8ET40XcU/Nc.aS\
&c,^R.64[[+^(891VaSTH5@B^S[eKE(QM\A)f)=,=2.?1]=6E8WWd0:&NS@1G+#Y
Y/>BL+:9-@G=E_K/HX:e=DOD64e.(ECQ<dL-=D4fU2^AA7Neb9ONab[[Q;C,?Cf,
^FFJ9VX)N):PPV0U/&[UcL6GB-JZeM)32]D)HW^E_.FZJZdeO;V[+YJ;)MA-FWO(
<bV/I,&F2A_P@KUbY,OBZFT,09@O?HJO^Ec7XCRD6)C?d[;03>aXK#2PHd-6<1@D
R;\_FBL,Jfe8.XS1OIO1<(6].VGPfUL2EWZ>.c8QZJTHJ\6OBNZ@9?aObJFAD2eI
A28&IcAX]a#@-8@dW+]IgS3;[BH)cS_<0^K->/56&-a\-N0^24:Q-8DVK1-D<=\5
c8_gOHI46828E/^P@.QXdM1LZ[\HY]I5>JO.46M(VBKS:-2SCTSG75B8dYAObNEL
-6V0fN1.)_?ULY:;LP^I(WA3ZWX6,:3+?-9H38&FO0=g1]A8Z3^4aUL:AVE+O;1a
:<50?K[2&#[22bJ1/JY2a4Z#:Mc9d-&VF)B#HVTMKB,OR25VW\PF@11,U46C4DUa
983bS8c[56bEU;8\@3[cC]8US@(?:4c=BRH(_TCb27M_(@13L&5577FOMDOab.[Q
@e[4(L.U)@)f:O]Z5A.8P>A\R,Ac]BdV@S2KBK--]RO<TDM\L:^W#\;.)FI8-_7V
dcG:_=/(1+c:N68:]]AEWT+@98dPg<9ZYYPXf82H,P&FN.-I+dTVLGZHRS0,S:6]
1KJS#S6<d\4]/b)dBQ.gK&g]VKQ2aV#B)/Kc:g+WA,B>68-TY.@LPba[a-AB\V(I
Y+8V(>+N7;gag&BOH4T<RP)c7Rf+e@YW\4UN7fa<b@YB6^2_gJUZUJ(Me[9KdHVd
:IT^-E-/gYfMOCU?@FJDb8ROXRWE;K3KK0,,dCIR>eL6;I>^-fgRPY,Z<&[EN:#8
R(5<J>D+5IJF<)e(G4cQ(+WUM\S\M0L)g\fcOKR27E=(^(2U5CF./(AAR3C;TV3+
dg&T(4N+0KY-WMb#P#GQ#),/.+)/2HUFaZ^L&e[NWHf,M.#U_M6gM0I.:B?VY+]?
2bf/E&L5(T/9RRQDM?SW0YSQAZf_8B:B82L<_>O;_D1T=g:2AY:2aeE0V)(,QEc1
TL1IRBB+Z;K_/<BNOFFf.b6OEaKHPJOBN&Y\<KfZ(dJaKQ-/ebC3M7D:@P2b5DJ<
eO,,(f5gaTe&A=VZWB5JNQfJ7=)OK@05MYNaXfHQ,f.PaR><ed9XF[-g<b?/R\[Z
+[cD/?+Od+,2aADR2A3D]:J1XLHW\NSOQdT==:+^<T9efeHI_K/JXF(WT=<H@(;U
=/.F&bYIWg1Z=GG_4Z-8fX])Y03LJ##E):8JS-G2W@-HLV/Qb->-Y]])M5+7<NK5
(+8PYa\N(]7d05L:1-bbBYPc[MB)9-E42Y^]a^1)Ldd@>,RIf@8]-;-.O@d:c:;7
?XTbaX9G=eFF3BYOGDC(N<R+#WATI.UV2/7R=2C.01K>f5e^3S2_#@>P^UL(R7=g
8+Sb,5^AM10gI+OP@C]XPe)3N/[07TO#Jc1O-V-(RI/;bD1a@QZa#;U@MM,LD=R#
4P/a8/J5A<QAfd@6R>.ZOZa+]-W7[4^?0/4D+@fODL]WRgfPYO&CD:P<Q=<JJNG)
WQWeJRKQCKXQ2,[<XIZ;b\E?N94a?Ff4QN>E9]\F^_C6,+GLUHU-7CbE=X2E0d#V
:=ee.T>RV;</e/cMO[\3cLeT0.Tg7H?5D+YDV@\7I<0291FBAA8ACXZ1#[R=5<=8
9V9<W0c)P9BT3FI2>Q_0#e[6?454B>>,^dMP^H.F?(_2Od.aFIK\2\XP//1MGIb6
(d@dGGR1\W295D[EZC;GOJZOX25Y-cCWfK;-8F1fKM8;e=8dLGVK(E:M,HB&GOg_
)9NZcN2SMA^9fT_IHTO:5H@C-ZC^S2=IcFW^#\]:\L1B0)1_XSHWdNQY[]^UJTOV
GS<EB\C>VK>2P=,4_-D0bQDeHBLLD1)(9A7OgWXMb,T^&Z6PHC-g]7\Z1F0G\:3\
g^\M+ggA9==9H@9e5DcJ\^b?D_>a)P4AgG5(Vc_DdQYQ_&e:M0@ZGfFHD4NO_0/=
80B)HA)6B&f1OK\K\g7_IJdb4:4<=AN:\cPdZX2(_fBgMcO:?;cP5ReW?S1b7,?H
CWX-2,ea+X.3LJ9-&XH][G/#[-M1AO&[GXg648KM#=U5ZJ(Y@KU#e,/E8=ANE5e.
SWHe][(84b3MVQeKW[8&;YPbdEM+D=a5&d7^9U\\-(a(@Sb8CM2L)e<1A[2XQL-?
?P6KUL.XY05IQ0-cS.KQHb-;:O);IA4,?7d9\2a0Wc7<W_):B?gOb?c_U,d@8O9B
Sf6NR0B?DY_&,daGT^CBSQJ3TTLJ\X8a^,U\7+=M6c?X;?I>&)P<WZ(VYDP:QFO@
<.RSE[Zd4Y<<bV:1-V)cQ[B=1Bcb[C2ZQY=Z:G@NH(Y.4=WAHdU79T4?LB]NX@#:
3_S9XK9\8^b5VEMT3<g=;K36aV+OKLT;1/,1>39KM_c?.5#+I8=D0U0TZe=E99[+
#LS#R43>MO/]:6S[fbCI?^g?2N>Ha7PL,#NAb_MX8HY:4,#0RFFAU7:L]9+HAV9?
bLg0(O/\02B/&B6S,-\^Ve8ZCJd^[c(B.@KVZd6IMI3S&9^W.Z28&BYRL>C<><\T
EQdSVZ2?UZKd>C[H>X((^XK-c;@^MUF/;@2WB28VE8IJ,>.)GMCGfW>WP\XPD2>)
/_LBXKV^Q[66(\e^#(+LSe&UV.GJ)P3.K1I(D(Q=X=+;-GBJac[S;1]^KG2VXfeL
[VJ&_aIG?@(#P?NZ,a=H#BV2?+^\3+d.MY)RGHL+6([/(PV9?(P<]]GH]X<K,UDb
8RTU?DUJDK,GYdXJE@O:47)6,f-e5?c/C(G#)UBC?-?8R;;NCeN?B+bBNYQ-NM:=
<bb)BTX&AQI)S[ML7VF&5XGO2,Dc+I0\(;+I)FQ7W5Sd,=CU<-(NFHTL,f3S1H26
^#Q9.QA6DC-74_<:LIJJ#_5<SZC;1&@9,Yb&V;G[DaB^<ARBCAJ:N;30/6;C+BNa
:b8:(=Id4c@56I3-a@JbF>P=RZRb2@CPWW^9GZQ@J:b[<Q9O-=W>a@<..J(>a^:3
O.:0f8_5=6ZS_:_)R??^]V9+T.V[Y3NX@O9+T?YEO1\,:L)CO3(15IYfaF7S9Q5B
\\10,]T9G@:K,_?8K7fg?9-VR]gH1?f:2JfQa9ZI;?JV@)D7A,7/9;.bOOa^9W9<
0QC2?F(-(SFPBf_H>L:dgK)\49WB[M+=70B1X(/SHf@d^P)c;&?_3(([UQa_e#EP
?45=CQ.JDF]e_ZZ5L05e(FG@V7]C?FV8gOO2b&)[RHD82MLe4JI.:YHa6Rc/_2GJ
gG,&K=HS_1/fO+fS&VW0VIPJ3.K:@WLKBcTCa6#GgP0T@/I,fNH6V]_Q/[JLXAA&
E#^:+FT#P]C9T+#V_L^+7U<K(,N-#50_8@X+b/;QV/R0W)bR#4W;T_1E;GNE_((H
^)46+;D:FXXYSe-dg4)_bdM+XA3G.5S)@H;9&GYJYNPK85YSH7J\FGMR4H=CZ?VG
]H2:=ZXX.0bf(>2V@R?&W&f:#4C2O8TWC8TTfZS2FB=R>BJa3LWgEdUV=Sff2.Bc
G=VbE>EQ=\RXPd;&+L<E\,+?S@bQ8(0cO;J:U3S8D8fK.TQ;DHQWQa>bRb1(A+M7
9fS+LJE\F3b<J[HaM@,UO-C)>:?dKHQJUL+A;,,7V[8&4f&^?1[b[83HH:.SK&[4
PCdZ=U1If>(<=B1-=gW\MQ09MRF2-d8GTb?OR:D]+g.cJ(+gd<+J\<a>ad?F\[ES
cK<DG+3X9NRb5JcCbbA40S(N0Z_7H#-MHWEXHB)eFDQ,1TK^ZT+;3/6X(6=IAAM(
FH@-:-M>V8_USIP^@W/#M[\SM#ZUK>C65RPPNV4JIN9T(KKHY31D7^-Ze)4WEJ?.
H<2VN2g+EK?cb(;<NDQ.L>\XI,=Xd1.4)b:B3@C<A<+4M4)WHMKH);YJ7B2F&4Cg
KXA8MF4_JC@bPO^5&5.]#O40O#__3[-Sa;:RXc#LUK_JM6PaQ0d_1+:G.29THfA0
WO]Y<U.,b^S414H;VVNEg?[U.^],.S,d(AOW+(D<fXUaA0/b8PMEP,U[cEdIS(cP
gMD+a]=HG&@:aTK;B^bHI(G]T58G@a6=#-79UMb7B@M(U_HfEQIa=+cXO+Z+[,@[
Qg]bDEH/^>FC;;POaEM+?eI=g[4]YM]&,IX0d3[8^[5[JQe-Cd<DA#^4W@JM+R\F
9VFSdCSRJ01+6YK<WUP.2-4D\:1]F=#L#,G/eRTBN?.QP3.E,YMf#_SDBa8eDO,V
S2/#.H>LKS(<]9B:bC(1&Cgf^][M3a&[Y:=O<J-;TN.]O@aYbIWMXH-<1QGb2Z?-
JRVB.f4RPffcK+S&GL/EDEQPJ.:&T_\7:HHR8,GY-92e\+7H,KLg>W\.A<3MefFE
)G.7T56RMP.56K,R4JKY/f0R,O3A7XKc9A64A^bfA.aR(J-&]0g?Y]/=RHLLLFXI
bg>\OE&KB1\dU99CLF_4;>eE>gQ59C(E9\&Ad:4Y2KS&2.+L<Z-ED^L>]AF\VH&d
TX+;WNPaeY((XQ&SdP,7e-Leb4R-dMcG;KHUQP6=8Sa5G,]MbXLHWH48&[C#9:[Z
DGCKS@TQ(I+3)I>:KFA\K3OF3]G=_Vde#S\Sd]).=R/+[:8N63W2N.QP-PVA(O6F
,-aWR,=6#D4G9;,1\6S,KJ)?LYI/DV+<,F^7S0fC&NP>2=WL/MO+-G&_4U0>ZUcN
^f6+JX.[JO&,.OD51((NS[?EAAEBd\N/23<GDSL:1H#ZW#EK__E,K2CdZGYJE+KB
F>V3F:;;QO>MZ/U89,/A4WJ/YYd6N#.K4\C^SP[H+gL.#d+[K4>--KA)\,_U>GX@
?Wb0R+eZ\Cd]Q-#g_VP.R++6cEZ9J:,dWX>7#\6fN6S&\17^,TLM8Qf#\&dMf(c8
3P<4;b=>&6P?Ad,(EH\2^-UeD.Q(IOXYEW@[G-03>fOEN.)Kb0C4\-g.G^SddZQf
T&HXd+BR,S8d67(2+3W6>4@=Na].2N##ORHE,Bd0R^Le:V#C9_d>a[>)O&dEYD2,
/+fPRMLfONIfS#PA,BMT/]&;X.>VI8ZF)&E=FG)4Q4>cU.T;-9J[H#cJ@0J&Y\Q1
.9;1NB?PL?Q/=Q09/0?;D.,](LI^.->/Hb^&58_c1X]5D5JY=-3[S;[3J5HX0ZZ#
Q+IT?>X_I4]1fC,ZXSf/&N=I0EZ)6X1Kf)HRZZ#32a\\7PJQc46&=DJQ6]NNYY@>
Fa([_WC410dE?5]JYGG1>KT[VD\C8_4W&3bVeb>AD2S#U>F><9<]Y-Dg;@F<;Faa
XC3IBc=4AP^cc-[b[)BY-<Pa)SF]_c</<^CK\@<aD_/;1M8<V-;/E5I?XeJVNc^(
O)P13.<^-5PG)M)e[V9INF]9)Tc<+SR<)VFV]7:QZ1D/->b+BA>X/HPfV?-5_\IK
Odb]5:2(.S/U9g](:@eZG(>:#&b/P8c(K/e,f-?B4Yb0N0cgA:b?5;>+Ub(WASLe
6\(@_O&K<4cG.01.d/9HAC1d+]7MbA)NP#beK]SZABHCNg@Q04.^L6?C)/6QP0:O
ROTAHS51&aY_TI-G7D41WUf&GBd60&WIET5L3^8..(+0Q,4,YTMPS>bV]A=+N_O9
GLJ\_b#\aeaB9RDQ=T##7W#O?L9J2A#(&6HDLYbUB5XSeef^Ad)5L=f_1X0SgHBe
7B96gLRDf)GKR,);N&^9>Ka5[9F2N3ED(\&R+ggG7R0A-6170X8IEQ@dB]dH+HdJ
d:,G4+dD^CX5YJ5,_EfK6E^RA/\9F#7Sa9B#aMLgTL^1@<H.g97M:&=NX6N-7CbZ
W;A49cEObWO+CWLNa&&N3XQ8]f&Na_8(W4M4M/18E@.GZaG>;P14]X#EgI.C]=-@
G.)c5CNB@fd[TU;P]D25fG<dJP+[]G@)+NI7JWWBC[4PdJ9&T9(c>8J1W^/^GR-0
L52a9f9<9&cd,R:7@82(O3KHFI:@3C#b]Uc00d)::X27A2]=Bd.+f,,.;,;;Z/g?
K+Y08:9XK6^+gAaKDff7P_6+H,_39C<YW?#C[,[LOQ_YBf+GeI)9,=LN?,\+d=8,
]d;3:X_<D@[H@&V2X0#O9.U?ZI9eS0-?agg0S<(E1,+OT+,J(E+XVEW7OAGKKf3^
N.QW\8;/:?cZc(@Q#[c)8;AIZ]A,0=bf@&/,]HG8YUd38@0GXf5?)A7_2Xg;ZbK_
NZNVGP=HeH3Z.TKONe,5HM-+DS@:1P(d&-b)/agA_#X@2e6Vc_U/)S6NPP;W76T=
.0>8WX1Z;V<I8UN0K9gafeM:5Y?<PQ3SbBd(EM7E\AE/#ZL2U_aF.CA0=;_EYVa^
==O@W6b(b]H/aG^VIL#]#aSAa@D(]3Q3d_@#3PM.d45TeXaQ0CX3b^VFX@)a>3WI
:4dA<cS5SaAWT\-=:YQG4WLQ;<(BZT1P7\G5Y_LMX?eL?]@g_^A2N\cZW=\:-\7G
a/6a+f)d:]RNaYe0;a]I1V)OM?942<3(:$
`endprotected



`protected
@dNP/C[T7K7Vb7Dc:.B4Q8K#6&YGNPAb\KWc8ZBW<3?E@G_K/eLc5)P_JWW8JbfZ
dWcV2>Y7CeLV0$
`endprotected


//vcs_lic_vip_protect
`protected
Q?bBdZW?c,CS:.d-a\.0cL<<ceAT9A6=b7d+eG])I:Z,eF5L7TBY5(1TSIeZ8QJ/
?HaW3\12R+,GI6\;J@D_WEb_,ATQ6GaC-2LQV60d8>QK:+)_&[XSOH;bOK[OgBDd
?YT]+.geLg:F#Ab#IJ6S8SAT2;Mc2-1@H0O1U_N?+,M1R?GAfbPSH&6=>O<MAZ&2
^9.gE6<\P_7-gB77CA(7:,9Q.-/bAe[S:)&c_JGQC&?ZBFS3>,HQcGB@N8gG:OL7
<BAFP[G0^B=Da)6bQW7HJC5S3E.:OO+O&(Zb+-?#0O7^-3RA7:?-a&BI6YY3WY7[
#Wg[e;M6[4g2N9JON)#,<?J(-IUH93WP5[d9f@072=E&15VL42ZgHXcLUP9P(Ua@
[?=2D@MYB(IcT7b.>0)D=I[cdXD0TB/]b9Mb6AaS\-fS&XYQc_)Q?=&;L(DQI]([
&8DME9.<EQ>FNP#3c?3Q_O?E33+KR7H^.KTQOQK#T=;bebPE89]aBfETRJDUZd0(
VOLJfbaAK+S<QJ792;5,eD>MC6^L2Q88?KJ:/EN^1.K+:5C/6Cg==10I>;bf_7/&
Y&-X(4Vc2d6\VQWVdW52J\J84W>76X3FX3fFS-bcBB7Zf3RSD;GEW[KHa&;g<5XI
EUG?6<4:9^X=C/=/Dd>-]757Q:ccd2bXHX@Y7#(9,EJS?1\>>TbdZ)Z]C>GSLALK
64MA::VKJYSV:=_=NN.B,/?/ZScB6RU(Y_S.:)@=8D>abY;+LXY-KN&\g=7@DN>_
?1>T\=?&T9Xd>O:E5Me6@=fF3MO#A]4ca07M>a-&T7/VQ;,g\FD1>#FU#XI5B5QP
)4?5SdTCQ<O22)>1=3:Md#BC+0#gANa,eIRI@a0>UOX[6UH2]]+8&^8,OZfG=NTY
6Qa7f49[^HRE^4[/4F+3_7:6J(56IIgI)YW[@ecK)Q7EQ#\^3;aDe.M37[XTa6OU
WVe&FB;Y608IF530B./=HR&8cT\KM+b.IJEHTeETNbDW3VZ(3O;KLJEV&2#_PR]L
VNK/U@-)-=D+^9_ZcX:+]@6:O4d^^@V<FOPA,AS@WH=UNX,I/6\A6S]P_2LaccS4
_>?6\@?KgbI\4(Y\A4;gYE;:_Z4(BBG&+cfEaQ.#RfI:K6-=gYd]D_bZLZDARSBK
.(4RV>J2(GH-KRRQ[NPcb,d@)>@AG\^^^A@FUSKg8,^+(ES6@Z:MZ^5TJO8+47]b
,N->TSKSL=)@R=_:M9g8F@7_6:8)@1&3.FfcD3\7gW9+VD&NTgeO<c#HL)LY6BKJ
^(eA8ZENdMF4NOK:c2..,YK=L>M_cgcO2,3[TV=9Ig6)g.]UX&231L-dKW8U[9H?
RUQZ)=/PB[CWI1=.+W19]Q+INH#0D@(@@[,>SCD;_?#C&(:EOgdR;QN1J<RIc[CZ
d:Pgc<Aa@4K+6P;P)aGU#bBFd,][C79F>OZXd1gV91<gWJU]7aBD5L7fbg8TV>8;
^,[e?5:;Y4N(TEIU@a:U,+VY=ZPWeF2-fSB->@A@T\\GORd+HL\dNAN<#;e0WQ-9
,9HLK3(XC4O0&bHN#KaMRPJ+S;@HPE@7XB14ZD3OI>H+ED,1A05B8AXO1QKHVOEY
=ZD:fg2:f1c-8_dFVUMbf1c[a&+(g3,7,.+ICK[RgR5d#G.6<>@N9E/C_2C_^@TP
ee)RFJ;O=])g[K.Y#CI_;cf-)TAYWLN+NHUfJ/IU:CWT+5XX+T&Z@WP:X:=9T7ZR
51_6a>bT77NR#[;T6[P+)?VB+T@\H(UJ&266?HKbVV7/cM4&XZIRA.fbZe4:7QTP
IDDQO\(aaTd>[-)1eKfc6gK([ZH@0EN_;?QaDX(+O:RS_L8)8]#I/K]#>[UT.]0;
aA>.9>=Ne^FM@900,fcT>HfOI?TgC<>>6KLgZ9KF:C72gX4T:XaN>-6\RJ3)K8WI
0b(\5L[c41-f3+:5IIAY@OZ>T3;=^0@C,>FEf^Q_[8GfKf/Z1ScD>Q+/#)3QBAY9
E.?E#RXWVFZf>0V<)DVcDE(9ffGN_0#b(TQY+;eEd+,,2Y.BMcZYJ_U8FaeJC@>@
H&&>fA[cFMA6]U^a65P5IOWg#)TD9aJTCK04T:WDg/G@.RMfK2Z2\d_=/3b33a97
UEFU)(e0[ZPE=/[\I^S_X5]6-a4>M-),/@H/+@RP^8URd-O4)dQfFZg=g+-)<&NM
0ZB_R2RBfE:5+I^cY6Cf:Va59Y1K#O]c_<WIa;^Na;[aEfS[_F_+;1\gR#]Da-HI
AKJ&==f282eL:;-c>I(]-WVAWMWXQ<SUJ/&W3UN2V0eR>dI=fWA<#;e]^KdYMI2N
c#52S.+P@^0K,K(7;c//\Y-HWdDX,)?)Q#GIO7[.?&OP2<V8+#1[]CJK)<Gc42g[
TRJ+SIE-1=f>F^GDKC]G0@Ee/OLW9e44Q0&;OeQ95)857E)ff,42\>?:W.Q:Eb=d
F-)0_-BG1KUJ=KK(:(&HAOb:[NMF_JQLdbBQNV^6LK&/Gg\2,gBBEga+,)P0[I:#
;\<[F1YH,B6c=GOBJ-HVYUYUEQ@=HL@gf,(--.CgC8?3M-OGNSB09@eJ\bJ>[H=M
Ib,M4MGGP(\6/9a/<5GNB+VSDQETHH4\W#g&G1]4\I2>MSa8<>@H/:QES@6-d&W&
I;536^VJ(:&:G3.5D//(52H7M^^eccA7S)Q]EeV0@E2VFQU)?EeVbR42ZAgg318+
J24V8gMR5(faD07bO5;H/RO?<\W/G+R3M^4XD8U9X70Ga]7,@+V;I3/5#W2[1CXR
;9\ge\RgcWFMRU^c=cSE?-A9NeO>]RQSA]&DS1KSfaI;D;4(]S0\3^(JScF<dI,>
N,.QA[IMB]XOYb]>11XSM2D]]N9778IBU7IgBCA,_.3TP]X.&#cKP[E)8J&J7<WV
;\\X>c0df&R#D],C=;B9SfN_Ze/(YN2ED\bS0]fd9>g;ebCGF>4eEAZR5+29CJQM
14AT&0S\a#\#cULH#e6?W#PT51g>dA<4S^NQ).<+/E\S/WY-^69(0gdgQX8CXN0U
=BfEWD?_I2Je7Q&N88#Q<J0cYL]U#A_I]2dKK)96&;MNG/&VHMNY-YY?eE(F?(0d
A70^1.>gA(/DFJf<T>c2NLacYO@f],^LCCRLd&GEdQ=JELO1C7OK+(g)<9BVY/0Z
GN<AX2gC:@(@CU.QH8:CcI0.D2EH+XZfTL)caT+V7DSc6LZ6=JCS3R6E;Ld@<(,.
W?,G@cMQ_6R4C:edR_f;U4R?K=/8-7GDE[D@,PXgR;YX/9g/PT\<OBd/3H5UcPcb
>E2:^MO3c7TZHcAXDa[3+#LB:I_I?ONSCBJdS@Rgd_<D5>Pgc<;IM=#Nd;&KGgJV
47O;M].H8_J-IDR]J])BXP)fg3Bd<c6./I+7;f)X61FQTgH0PbY^A&++be-Q&>19
+L?bXU>\CKIUXXbCFRf/<#cVedN+=?M0L_D/[A7UT^3PbdCQ>[b)[Ze,FS^CaU4A
DLdeWJ(OP_CWSJbfOY.OA;&06,L(2a1IXW,2LPY6=cgD^9AIVe809T-XUbKUdDYc
ELAWPG.T27DPJLTP;OVZ.aN(K@+J=.@da/CJf_1<@G><M\[V7QX9Z.J9E<T8)OQ9
2NWG66L#@g(4dc(W)G3BAgg:K^@WS64BWG,PTA[V)5[)0-MW<AA34<XabN^3feC1
bF3<0J6+=AgNWUMZ<0JBfDM#gM71CV.)^g[g:=?&B.(X>TN31fE=F753\efI_g^;
8gWZ=HFH;-3eZ;b2=WR,V9074K)HY4a9e7\)9Q#.3@38XJP[&5?R56-SFY1Z6c3E
<NFC#b)/)b\ZR],1FIf;@H-Je<5UZ.;5,.YF-UV&KYGH:;H@R]f6WBYfX<].8E;Z
g,>273XTMW=NT0TG])=)>N#:641XU])^)XC,&E^FYPSZ@V&eRfY>3\/XJ-.]:B:N
XgN#HZ>KUO[=:bP=F79Z3ZP6-=L_RU@Zd/aD\cK<fI=^J7Od6ee9:^OAVCccT&>d
>8(>/a-:Sc\=+KK8<V_fJ6CJP0Y&E(dI06AY9QVN0KZ-gEb(D-VQJT7d9CAgJfP4
b8DOY\1RZ9;;bD8BZU7KF#BT>8MH1EO[^g<.Dd5[W[;D]Ef\+&e7c=O\f:cSc&U9
200^>)4eZ4b<?)Q^4VFY>,THA&R\-)WF2V3KOd:?ERTBXXH04J;][g+-QVH..]Gf
@;8.\^5Y079(59H=JJ\7B@(UK;;7/-?6B8OeG\YcVN9.bKeT/6_#BdRTP+,@IPXW
_;g,g,&Hf;V^O-IW5[Kd7AcQ7eF9C;0JA/A2G.JQ0NNc>EN#CA1HXf.aEcH(14Tb
=L+5Y:H#/0DdEUME6c7N#Y;c4>e\dLLV5+:c8U[4.QF_G9PSQ7OE@9(SSVNW4g;I
Z9>2[U91YNMHBfQU2IVJK?C8@d_gWT9c#96U:PER@:PH?]6HPZ#Z:Ef1/deAP?c5
\X:9A;Ab[/8C&FHOIcE#NKe6^L#.;Gc-61_]GO_VOUI:7::c6gd,Pc3X&^3^OT,C
(MT?@B&OMeLKP6,NMAIe=e,\7Y@IAF\@eLO:L(ILc9,ZL&.O/8QG=fI;F^8ScZ+=
6@&X+M=NUSga3KUDFWSU9d)gedZQL;HgE<?LJDadC[Y?(#<K&c\7#D0W>BbA.-#]
#+;ID\aeH,RX&?;B:88U,&@W^<OV6;aI>X7_2&/E3(BPQ[3IdK)(PX?^g.:Ue8:G
:\L0S,6W8ZZ9Gf-Td=He=+FW4>VOb</Z_Xf58]G_:gM0OD+<,c.F?CBSW36)/a_0
_:GfA(Y54B01ISEaXR3>PY7C]]Iec0&[6=0(62aR8RV@TX=#5^HJY^7bRV.6&.aW
2+[14E@Q0dfR#;OKMbUE2?9g=/)JK[NA8_Q=(9E>1E=Q00M6Y(MEP^(+E9U,0_//
VW/D)M9U\XTd86?I.Ka\Y)Qc:U6]8#?CXKgeaW=-Z/BXgK>0^b;1Gb,,GR_8G84W
1Y)[;21NP#YN\PV/LV@IcH(YB8R;:dM5U4,K=UF&WKVJ:;).P7a?UM#VH+F7GI8Q
G#64((LZB>XUC[>VE0(D&M48<9K10KTdeVeXO9.@:C7)1IOSa.U_#-^GO9C6,)>,
6B/4^K(R[@UMU&aXfS#)]HH4KPE;2.Bf(ETVM9CCTBPR,-.UD2VA]bANeB3H[XAg
.C):ZX^OG)1:=1>?:3/MaQUTSe+:Oe1JU9)D54PaDa,U_EH+;4I_.+ZZTHJ7=PVT
J&3=2Y[XM>J=e::e/HL,A#J[geL(3J]BVCTSYX(P3U8K.GOE.3VF(]WQO[(c&^.H
M6WcHI2.3I&HYdT[5Q;4#]YFD_U\_eUHQ.QM]NcYfS02?dH<>V=WXUb6WE(;3BR=
,\b__[&O)&<H,H7FQT.V/EBFPGLO9Y.\T_(E[@@&N4d:T=,ITIM1cXNddY2PMG0.
L+P0N@TSK3E9>EK(5OJ#N)-GH3MRg71@PZ2cG8fa=g9MBGA-XUF]SB@^Xd9fNQAc
d:\S]^,>Ya39[=V9\[a4A[ENc4JU/_PH5g9/\=9D+e0UN.):SRP/9B(L4RPI/6b>
<QK.QL.;FR[@XUHT<T<J.?>V5LWYAO;cfa+X2)[9A4H,KK3b5ONCU(-DZ1:#:.9/
G]D>JfPGabK1-UE1TT52WNOEAR-2X7,WO&4I?b_TJ>\=;.V9.4&XGSMFS48AEb;f
DK-GDLd=1SeQQLGccA==bfVVg>20;e]A,5=g)Pb3\_:cOZI5PgNc8X]Qg8>UC6Y;
6^4fYTAE10ecdQcN5\;:?M>I2B>6>=1U.Q+aT)Hc2<C230dg0XGK@dRZ<L@Uf&G9
77HEX@3@]LY+V]9f8;MH(9)X6FN[LS5&AQ-WHYNX,;2UGK6VH1@<17<]gUIK,X>5
4GQ_NQ6T<P5OOA.1a<)JM):F_<<<2X<WLXIZ-:4W>:Q+g#X/E68I[PWIVDES.2P4
;Q_DdfI==0:TUS-T+.d?&<JI9d.6FHQZ2A0H3,HW/-FWEX1R3<V2JZW#7ZBK@?g6
_=KG&1IPY_\f<(d/ECT,KeA1LM6DSJ6c6C)Q6BNAL\:77ZI1&_6&@EENW/gM8b;R
?CE_TFBc@;M#;-N5fEDO4)]0O;FfcE#CCcH]7;)&0]V-XOH_GMI8ZVOHF&)Z5V=8
AXaAbH)I]bcD)e_V,/eGbc(&e(-ZIIF4.W+eSMf9T+Ag[:HZB(gJE=-DS30BQECT
C:;B&O(c>MI#V:a+C..G9(QK9RT<1HHQSc3c+L]T+cM0be)UXF1&6M4dfHU0d>OS
L_PR_XL;H#=]F6WT>XB#f\IAEOeeE.\20]846gd=2A;-#98/^--QYO84R_\c4Xfb
DgR^eSWU@.I_C]U7Pe[aYb-bJVU:_.B3RTI/eF\[?80fNMZ1=EI-KQH7I58VbL9C
;=2N[8T:YWQFC4R@@DDeP?&[?_-C(4M^L?A3]7A,YgK;]2=^4<\1UU[b[V;a?A.3
YLX\TDEDC&@2J4)g1SQ:B_C;CL.M^^-@F\EPgGgaB,@/ET&4QUGU#J16=JS?HNgN
R0/JUUIGfDYL>QE#[9QFdW;JB.H^bK9@fd(b8;g-JB)DRG#eH(3C2E6d2AJRd)VW
HI:&d)=QG=#;/BDD:0=C49R^A[.5e,7#69)_D[:Y.+A:Ig>/P.AfJR5_V&P>.03F
ADIBCT68=8&P[\I;?HQgPXSd:A&H4MUb_<1b;ZV=3<]1C(\bSY[M0GL6JN/7CF(6
6d1G_-@.(=^NM:,<X.>Y#cLA9VYADI.K[0f7657ZHMYL_^CE2ZS8:>RaCMS7/YIA
6Q4bRB\R\NbD((NM:/F)OgZ4>P>76PHHZY2aI\Ca]W4Sd[E:N]_eb#eS,2?gX@)c
\7P=R3[gKGWeO#D(S?-\R\2eTgO-QF93K_6/],)#IY]8RgE449J12X;6La\20EFf
.\-g/M\H>9:(Ag[7g)X_bN#KKOLg5..:PW-BL8#7U-#/9STA+(bc)@=4N\EL[^J7
H.V&Y+IOf_/E1F2U:E^&]g/-00OZN#7N(+>VX7589:gbgBC;KfTSI4-SZ/PWI343
d2bFQ0PH;fSW#S0:WUJd/;?-Ca\K@?g_=F:g)DTKD^_)1?:K<^.MFFU59BOHQZ7H
AF,fPeWK1>37G;B9a8)#40_\IE2NMJ1BWC/XdI2DR_O;OZ@O;-0[aaMb9EQ\1b)#
D?_D3X93U;NaD99+^G_Jbcd^M]W#_Vg?ZS<69>0.F2O0+#2[=9[<D#DB_@ba\:-T
,J9B=Nf(4A/?RQU.2Q[)K)ZN1?LbC5;Fb(<PFTJT,)B3C__+V@0EL(_1R-D?Fc#L
e=?##JK0IX\MRVAe(T]6WZ],3,a4fP-\(_U@ZLWWV4BfF[F:<I,Yb=<A\YA)5[(N
1GA\#;>,&FK_SY?Vb7[@QW4/aBPJd]4aEI6[((VCX(B<UP]Rg2N:GN-d=:N,DZ>G
6?8AbfJI]-b4a1,WNAF@63LMG=8<=4&&9B(=.aN:BE2bCg/:&5W7F&@7(f&UB,[g
?2K(>-^Af=V;XN0ZLfX.[<[6ZJV<_T@VA/NF\Bce6ADDZB&:N&8DKA[X<:XU+VA>
?e,&E3EG:GASbb=+6fR_TNU@[&:TAFRTdVP3Y]NWWU<O0G[e<BgW/gD.1,?9NZbP
aDe36_D=6HULJJdAbF/U;d_Og<Sd-_3\/L-];30c](T?V]B?g[faM1954cB\EdRV
C24@&A]9L>9HD&N)[JXca#,;[7:G<RIf;Q-]>QCdV)a02G.aH;XA,\YdOWLWP+]L
8WDUV]W]7)/]cDSUfgB/4-7g]R+Jg3A.KKcN+6@C>MN?63d4Q);<(DSeYQ[ENY3f
4TG>8^,f+[BJ4W#0bFJBA&HY=+;((I;@?)ZSBM51C1S-8Le?)be?AE>\A8@@I8?e
Z_()MFJ?NUN)43S\_7gEcIBT>P?SN9^gC\NE>e1U5OXL61(Idaf=bD#.b@Z.Xcf8
CL0;UJ05L(Q5&SV^RgP2CPgU@&9V_Z^@4E0BS?P#\_<RGZZX#=T/[K;>\8=OYST+
&]/O=9[OR1GG^d?TV,(^O+)2[PLK[\HVSVPHRL^\G3G5?^)JDec@F&UFAb6_(a:a
I&^98A;+d77XO4AI)=[^;7Y3@2ScM\4^^JW#TS2RW+@^N\ESJ/fJU:T.C>XV;TD(
bSN,H9[\E^BBeDU:O;Fa1McD)2X:eU)aKXCYVJWUSE.>EG:6X=YP,D6\QSQZ/b==
5:GNaP_MI8bV?;H>9,E\9N/ZN&[O8HE0Y=GP,X?25;(9IJXU[Z+VZ:U-11X\6VIC
Y;+FW(K)#e<U<UE0<L:/UI2OD2N:PcF+C3O7WM:3)G<Jd?(D52I8K+\BLM[#d.Qb
H;J(+A)ag&B+.6d-H1gD?GF5R#(ZNH-CYPTO/E]U81fQf=N4)fdG8K=gG[V9b,B9
@NBeFW?1f,<)0_K+06S.AT,A9R+:NH8/+&I8YV_^>O,:7bbXe,Y<XHX8-Ne>46U#
]?^2LW&-G/]JfW#e\TZ1?0NYT#cL60=M^L=8TBTT#<PKVa#d1;7c0GL6)3.\dTTD
]Hg39f.,[d]f3;4I[P52bbV17)J]?gF)&\GWQ^,g(EH+??2@RL;T377W29@C&T@G
@)XS_:H^E9CZ?[fUU8@c?gX(#@X?WB=<Yf)Q[_GCY7BESM?]X<+OZ>\Pe1.:3JXX
WWb6)>^\&:M#8J+QQ<^9KcRA5XYR-c53#IcK>H)IU&B^\927#@];BE^=ga/c4#Y6
<?c9&L3O+1\/=X53=Z2V0/FSSRIFXI<+T9(fgO;X0_e:4LXXA@BcXYQ9OUWVXX6:
39CP=GFGMbd#H4ZTP^Z2(Ea-RF7[CYe-1]SRY+=O>K(ZAI8J2\fgBXO]edUG[-_V
J68W>L7PSD5&;E:#5aO5HR.U;.;f]aDZ23Ha.:HR77P+)O5@FX8VfR.cg4W13/QY
O9NHA[gLUW8(R5NJd/RC+#9>#U<0g-CN__4Jcb]3?]2a_SP#INS1BZQfEHE#6@8d
&P2LR8A:VAQZNfGT9NX]A3[9S2b4<LLDUKC+X8S@(8bE7g/:cENN>W)XUCBUVONa
?AB:CK)DS3R@0O^NH_(bXWX3BeX(;W0d<:/-?WR=#A^Jb0ZXI<5\/35_0a#RGRf&
A^Ba6&8454gc0LXCL1GDBA.9f6[/7Y]J[RQN+,0PfO6A?dT3:IfeF^DEJ[/S<T0^
W,3QKCPe-0:QFVEf9g;K<HI[X8T5XDS^1H>]W0BcH]+KWD@930CMEf<MX9ZJ4FQW
Q73H2N+(2Y.7;FVPg4Qa=c#[<b63JB/-D/_NPQ4ZX1HV\?AIE?Y\KH3Z[3+^M,<:
.>@F9C_]L36KTVU?I/,(1SN>RFdM?#8YEXPF8DeICVf./#1#c_JXNJc8Q:MVZ+O=
I5fT87S<3cC8NBO1g(,/E\5V)a>&HeJVT2O_C\1T)7)NNe\XZ?V1T2&:)#7ZIYRf
M^;CU3VK)8Y&\6HVUTfTNFQ4N5^3Y/B(.EGY(80Yd-Vf]@FA>^M+Ddb[5U^J&JBZ
CW<ZJ9-N.BgF#B^#&53&H<].6T8#MH9HbU]-3]<#I2([+\4+(68:Z+S60+#ICW\\
QR^#<^58S1A_2XbAM5bFTF1).W]Y]&Kf?-F_YQE8&ZgaMZd[TaA_+e9II<.<Ce&=
eZ>PO_>HN(7D,=6eY2JYH9C-T;c@ER?I@,V8I)(Ogc]B83A1dK^8d>YPKPYJB5ZY
0<RJE.UUV&Ee_N+_7FDc2&\2HWe<&N#+\e<99?QTHF46(LVYC<5@f\IO<.c@X#43
5Ba573JX#N#TJM3T:MW@GRQ>QM\_-89.(D^4-e2a-?_(KTGX-#K0IXD>VKf.SOO.
a]Q2BY2e.Tc)2YX9U@Leb((=_@b;O=6PY7FN_QPNK7Y_B(Y^Qf@8@],TB&D\,TSa
.]-)]>>8Q_/-;A)UI<4#&1d-g7);6MaDM^F=Mgd>43LRf8#3E#DEEC?Vb2F:5^PG
47ETIKbdDeD:0d3<^OW:.PGGQ/]YO-ICdU.7VMTUSC]9OA0XO(XNW[Xa9JT3MA0O
+MSC&]E(Af:\NK(54DKNK2NS[77>[</Y3R,HP4d=R?g?G>WeL[50J<5(,4e85<QO
)ZBOLV/_D^@+G[,)L4H,,4H\,5e8MYdcf;2015J[DO@R,PWc[Sfd.f?MHRa(UI^8
I>CA&T-[0_TE^,eg#FWFfQT/=0JM=f,8:XU_NYZFV<V8#3A7UMc^-F@I/IQY7GcM
@XM<-S:_AG\/SKU_^0^+W\/MR-7VSLT:LGI4Q32d(T73cI2OdG=IL(_]V,H#cIL+
J-RIXY#A-?eUSg#XEI;C=Y2ZUb.C0aN0C_gS(VU_+275P?WR1HPBd;/&O@DD;>Y/
:<;BTUT>EV)[Qf525XSA0I(<b6Y\eG/=bP\Y:PF]=7_BSNXQ91HSJ#0HfOb2FQ9-
^W)?gQ-24RaS#??Y9O1.>HJ9N[?-KG;)J3N-b&80-/G7X3]VBDC(^FF0>fE=c0Fd
K9@19d1Taa;-a-TE-0PN8K>F]CL7ZO+7GYD8P^dS1Y&7eab9\L4:^U@U]HSDRWf6
aAY+Q6#gRF6HgGa[_O-V:WGWT8A@LNg33S&DA.M2Vf0M080_LBaYYV)PJ(X-,&a8
UXbKS+dYb>dN666ZSLE=e=ZcRE7GD,O_(@>#CIT0M9e3GDNC;6<,ESR56I>)f05U
7@C[@T>(T0/DFY\8e8[PTI#ac5?+8K2?UV87H,/QIG(>)bd]LJ[9JKeI+5A@\[>7
@9VCXcCdGa)GOA^EEO;WOc#8W<-T:M3&OO[OWUAU,aJ].B?(+RQ:>93:6fE/\89_
YH^3]MHMSdI,5.=AN3(RACGS^Ff?X-bgYTW9=]KFJ:0[EM:9:ZIRQAT\KUWE4KP+
bCDeY\Q0ZNIR41F#OY93@cTED62.bcFT<2)V.,XXR@Q1=&,\3-+Kaa\X)ePJFO()
^ZZ96ZQD\L0;.].<RJ#+O?0F57I&78Na#U>GE^MZG6:-,b4EMC>##EEU[626X>b>
R5ReF(R_2a2;:;DIdRJ#T,HOQ/Pf(>ODAF9+Z#]KIPN3F8._J:4AIVUBN_^BN#KG
g0#?84.Xa34.&X4UdY();G2[O78SN0=Z#:O^D<[=F1@U);D<O(T\?Q;JR1,:V]FW
]8B6L(81RN4\H]2)NE:1+(S+A+=:1bFH9Ucd)N<=7+7EB09(SX=/QOTV9R&Re=DR
7&:LGM+KHG8TWQ;;gMdGOMUD\N.0HAR9=^MX7DF,3eGC_PCG)1JHOI3-Yb.#LMHC
[KTYH1J\//Y5+=bdd)72>?:FUYRa9@,_8+H:fe7WOTE1MF2M;S4[MOOA\[9L7#bA
;(H[UIVT/+Q??A(@G)-1K@,)PgP>g6./\e[XOXEP3H1=8<XD[.&cPP/+\<f&7#-9
La)1X&<b]:(QC/_W[g]Qe0FZKA0R/O-9S?]]SKeb2UbdVJLfU;&Q1=5?O67AbdF0
]CZ9N_7J@](,9fd8X^S:O/RTQeTQ^cUGT#@//eW#eLNB2SeN8]@9Ob?T,=TQ9DG<
=Q-a1dUN.FB.<2&BLc_MI;,g2+<8HLTN,UH.E;^f&,4M3)X4&V[H+OD&>7BX=Qg@
7T_>#3M]?[@=8+HO<S0QLHK=Cf0HbF<[=[_IA,5[8:>@,\VgJ=3KF2-.<D&ABf4^
AHd[9=V:2I(&7R=OM+\DG@G>N6/ba]X8N_b-e(IA2fJWUSH(-4NKF]\5TX-;&^[-
A)_a]V?+=ee#[HA_8)bKbR>&Z<>62MI?LA:JV[SFYgQSMGZga9+8IFD.\#XD5LB#
[?+TK;R-;]#,7/RMeGT+EVQ2)I9HSbRc_&GX&aO[KVBf7O<K90I4-J#bZ),DX5D@
D<8@,(QRDTWWH\U.-Q1P28F\VLSdNe?QN39NSWB/;f4#:La_Z1^Ca4/UL1./<@Z4
BLF);WD8bcZc>Eea]7F4\_SWLSV14KR81f-R(YZNFP1,<ZVF3-]:NQ\J+2fVSaTU
8PH-T@PaMKZP3f1T0REdfZeG?8(^3OBGG6XPFSS4ZVcgZR;D#eCOe8.(YU^Le<Uf
0JSAX,GFdZL:4c.U(YEb7LI38,fL80W]d;(#T+^0]MddGV<M;S9)K/+=](L8]W&4
_Q3G)bLXP&3A-V(/M4fEA.7E^DKDN#3QS^OS5?-eC#OI4ET(_OS69fN2CMPWG<4_
@F[H2+;_\/1&X\GcXOA\Y7Icg/e-A4IaH0OFf3()O=eG@Y_/UE4;6&+)G34[_F[C
/#+_1)-X,=,5AE&@f3RK5G^D.;<d.gFDS5c5D=Yd[#.Z#1NAWV]5?a.+8P0/95Q@
#X_?J6GfG]L:d2(e/J>=d.ZIWFVAd+WAP]]8O+5XGD]78#5DS8P=U8&E7B8>N6M1
UDVC4.7d=9ag?#0\+K4PQfa@O.(bIR)[EHI;=-Egc;?PWM5ge4_@]_Xc:eOd/;R5
S]6B4b=I\1S\37>ScWYJNbFAF_@UYc^-Vb3UFJ)dB)Z/[_\L,E]65-H=c9Z0L,^J
eMJgYS<;6B<#<)U4VWZQIbKG@+&:f[;e-XMGWUeHZC7#[7_ad+V\&=5fX,&\Tb05
BG[/4:7KT9\?1+gCOTYSS/+V7O@EfSS1gP&@H)6?NaWLO64M6@)4L;(.Ie2[6]+<
8G8Z0ENERfU8@T:N5?^?5^06&A\1bbScaK35Q7DCPC.W6D87(>(d4F<&XYUCCK#K
N<g:[G0;)0.RQG\LPSTWFWG=MKf8ADWFM0VF-V)W0d0EUG?)^BKJFTQ)AAB0B2,^
c4d3:_3^U56aO2@ZPO^.Z;>Z1Dc4>90]Ea<U^)9V[]U+NQU)a/Y.aS#5d7&+Z)Q.
O89SDY0NT6GaIG,a^[&7aFWQAO^H]aHb=2</KSLJEVUXK-+4H]AG.5cc&Y01KB80
ED<WF(7@TI^J>_[I@6Xf;/(U4;&e^T2CCO&&1\M:3OFP5\5F_FcIKH&E2B)Te4[1
0F:B\X-bS.DJ]d5)PW-.HJa?#-a@fE83@W^-TLeC5KVLVMRFJ24EOI1;cWLdQKb_
G[a5De774Y3FLGGM;Ea^cQb.J>:Jfg[MJ5[7XMYB4,HW2g=bK&WZ>(34)([cI(eW
&T0?#CBM8T6&eCT]UAgfg7JLDgA/U8IZDIKW&P99aZg&gT=SR-YbPD-P83ZdA9e6
cb/2D5&BD/;_-RX8FO>AV-S:<G2e\#G_@FBDI_=^TEf_b>G4S1VV4ID#dHU[fIED
CH?)?3VLJWCFg)Y^TdWZg[:6@14M.0NBFYED.,KNCG<:I_MVc^Bb>4FdE+.)bUL&
WNA<+@C.a<W1aa>Z&4AF1+7V2&CXFN^/\cX?8696-;39B=+22C(\8DH1?>]D=\U@
Xfc5e/<+8=H6_FNAUb/g9cSeE/#+U\[Q=<.W\-W^a/H9@2(GR7>V<SU@TCg,E&,I
\F-ILNL,V9][C\+B3(H\WHYE:?5]JJAC^GG^QfggNYVHf,@S.+;B:^Y5(H6/O0+M
7/a_b.e0-4gRZNd3<cLT_JKb&QX8&B;T<f+K;B==aVLT8)Q\Z,EZT)U8P[CHL^EN
b]L^[WI&6/-cOf:_F,Yb#KOW/O+?SMG#=4G@FQFAPM]W=E7GO?<]@ENb4W+5f,7,
aAJ4]&=#B50gIFbBXR8<-H)&Q5LXAaKA7LA0CV0?X))N-@e@ZeBKLRNb-#LF1I/V
_bE)0&3fROK&.:/dW4)7<-FcgPaD:S+JK;[P=7([&8a?=90PI]&cVOBb5&P[J\>L
+2XbXae[aF><^/>&K,b<&e-9J_3G>,ab:a7ScYWUWg;CZG:a+]+E0fZ<-W0+(a<C
B7ceZ-EZ4.FTKGA]3Q8=M&CS[-U]:dUgT_7[9\M+P)K4W#>WLFK_d_3X,S,?0GEF
MT=Q]C=UO,2d5D[;ZFeYSH=;QQN+df:Ue1A4_AU>5E0.JeC<[XH)[GbS&#&)@6&/
;GYDN7Ied1.=0;Kb[:.a?ETIeWUaK[bFc./KYcfS0SY,K>,.=T)+BA(R7#^S>/2c
O5E&\JbAP\aXTe@D9)4L)D#Tg;[g=MG(@<La=B[R&+HaSV?_]);CX].Z6T;Qb?[[
c6^K<=6SDC\^<\9EANLBO5bES1HGd29Jg)G6#SMDaL_79gAa](D@53G(RUS3.C7/
Ea@):R<\-,Ab1U#<0IJ6eSde[7#g(7=4Kg:A3PdD<XA9@X2bVTI^394a>BIbUEG\
YVC82CL\?-JYRSf)X&F5;Ka22NL+JF?7=cb<;^TN?8+R=&[(?OZ\)aL7O^]C-6P[
&Oc2X(;Je:&U^\bQ^bK.eGD-EIEfgFR6>=X]@-,.B],,\O;,<>VON:;9]=)TT>N9
/(:N\ed.-,UPOHN=R,\A<?_@fTY-IA;;7#UXI6].-)7<ZUC@dfM[<C;-,43G.TRW
-^PHHIG;a1K>F+52b495A\^a4>2LQ9T0+^#dWWb(-e\-3#()8=,5F;6-A+N+)5#Y
\A<-ILg8AS(??c<-07UaW4fAZ8/GQX&XJ>TJ:[+UAT7,5QL..RFL:/Q8:R<)I4#9
VQC3J&DF.5V@V;8H1&UTRIV(-Y?0Fc>D\3^3(5Dg2Zc\/=1Q];?</3PaNC4f9NV;
c^0.DZda)6X/6:O66\6LJV6BDKPY0@9(@1UNaGHD22WO;&UF+#BO7dNC&(/@W:LR
Q^fH/PB<ZPeV_H+@gN0K^6F73:-K_ZgeNX+-_4M[FCg;cWd]1@1^b#aJ+;>(1?)6
J@cW9E0^1H2GL6Q7GUde(S23L667G[,BcFI)Re3cg3..a/0aOG5P4eUQffCa++=g
,O-KIGA8CN?8TSO^fF=e7c223cP=R:=(+7OYW&d)U6(+\T1g;eOC>(31\aC<<4^g
26[N_^S&A_7JK048I/FSYHGMH:R^63cI=;B:Z-G_Xg9e#P]J&63Y0W>c19-3,PJQ
.IIHFgM3SD4Ae)FMK:L&dG\A)O3S.Q;B0PK:@HbH/CcG38:U1Be3<YC0=aJP&Z=U
Y(bP#U48\0>6NV]?;).&VG,38GFLMdVT77?)LE5FSc5]4C=;;D+UMKeS61(HcV=V
aU85Z.OPQ]=#-gLKd.#.eR#f5fgLPW@eH]M^HVQ5U&e&P.M7;F]^.:dLHeKZ;MUP
c6N>Xa+FN];+D>gfY:SGSTVL,\[:ZKd-1;9GMc0G.4)Qec;:(S3;IEU0&U5?,Fg5
Jd\EDGNUH?:YMb<[&LY&L(,g133Mc;9g]e<NIHUFBJ^,Y]FJTMb#7;F=@MWC7T=-
_-^>?S8?KF:0;7>4H^<AOM?)?ZT\&S(]8(^1<.cec3[g_J+0N@f2#:4G1QWWI]YD
Zc8WNX@Hc#Z#I5.@,>1(:Vc5(F_Yf3^BYe?#IgM_LJ@cg1M62)N@_OV@V7TC^.ZQ
8.IZYIJIK-K(#L?+>QJU:S?gSdGCRW2d_<K_S]^IJ>^QS5W(e6DWc7MRUK(d3_=g
gP]HeKI_A@gFMEf-XWSD<BVd-QF.fCC>F&caZA:263QJ8I:(3.X,,^I,ZG[AQ^Gd
5EX)=))/JE:H1?[>EeF-:g#8g2:fb1H9TWKWLZGGT]/\aR/db>@b3TcQ_\#R37E]
@QE,9M+8N.1=I3;_-B\N_/I24?MAP/Nbe(TIGP8Z)NUFDJJY>]4R@,D?Y_D#Za\G
bC,@K1X[?OHVgG)K)?L7S>CTX5A_:aKMBcGcS9T@D3BI_+UFNUD>)<&D&^Y@-_A7
W2GXAB<c5_AY?.c-PMG#K73=UG:A@W^f)dbE2?]:J8Je,EE#XLAT2V)cf7S5QMBV
gbB4A7H8Wf5XNURL@b=T7.eN_>8.#dZ:f/8_(C//ONA+/#Y-&<.-PcL9f(,/3b1>
XX[+:ZE3,IV4(b\LWW\\RCeX9dS\X6GdCL&dEZ@W0.^?9&b8LGb[BLf2_Z^[G,:Q
9?=&2+T-\S,T^7S/T^URENH9BCKM_MS6dZZ?X]Pb(G#e,?#8?aNffWaNPe)>7aRM
\,0#<MVKC>4eI.8Ab83AUA4#(JS/LJ\N)4GZ8,_8JT;T[GMc+^3^IZT(GZ]7=/ce
M9Yg?GZ]B:eV2_907)ZCd5P.H7KcGEUHH=&FC9]Yc-XVAa>:\]81;5f&Y=^g<?<Q
T8QQ4]Y\Ica([c/,_Ra4Y^DHbB#ZJ:,@7_DP\CE2b4SH05<TK>;;[,=VUV.(G5,Z
_H<V-HV\[20\Q@B:<.,5gHbQJN7\f#fZMCaV6OBAgYJ:+]Cbe(SL[6FXeW/SW?L1
#(EF-2U(;2_FgFT-FDCR=4@WY@eCZ)9?g,M<J\.38?S;Z3dPFGG+d\U&5YV>VMf8
6+-PWKM&U@dWC3K5K:A)6<36F+HeZS-J1^bRdWEPJVd3()(T@85_V\:V)B654.V+
0cF[G[V5KeVJE;eHPc.J3-aNY)@2/A0ZY9T@571L(b39]=UB?J)-\Va.&]TMRO5b
3.+]P#/K0JA:S0QLXRTV0B-.&fDccRY>O.42R0SMK^=R01CW2RX2_JD9>[J\.S1/
)&AV=<TK_[?3(8g#[807TYK)c-=SY;KB@=d9:IPDZ94X6gJ\C#YZC[C]VA8Me]2g
gb=M<AON\8S2U](]YUI0]Kc<?f:_G<g&8G6=[&8<D\6^_2ZgbJ<>2(TBR[RGbVB/
RP#fLJSW0&:dHGfY4HC10]Z6E<UZ^C=QOcMPLYS?S>X,WHU9P5\-YA\VSQHN3(/R
HI-WV_eZ<MKf>O7^@#]KIEe]F\=]K;VH-/ZO/)MA[@4?8BbQO4:IV^PGN;.K=8,L
gHG&-IQC0/+HSC7^JN5_J80U/M=KO8F_0YCbaFIB&.Xg#KLBagYd^(9fVK.H-7+B
Rg2g=MbANG@BGY?[02[+]1cNVZ/3CJPS[STSGbML8eJc8&PO7f3/b5EE(SN-cC_3
U84.RJ<6-,c\AY+SM8;EM<WW1,UKX?M_XG7e3gdc2J8B#M=R\(ddZKAJ3/f)dX4d
Y6HW^Faa=:I6OCM5\?feII2\D>c+JQ9UcIP;(&QX/4D:Y6@(:&ST+OZDa:8SA-(U
)GH^J+Pbc\\=EMA[bEAP#.O>]_H)B,=N4IA+YeN][3630:?1=7LLb/;Lbg8049b7
aY(JBK,:E.LId4J_#cX0e,)-#6;c<Q^G<)SHV.)WB1<2FVN@KK1)IIWX5b>Taa40
XOZ1d@?b/V.;;/fC[TM)L@6CQ/4-a2V9+1J(abbBD24cW+YSUHOd>c<ACVad/W>E
1&X#La&CNRAKQ)^I6cL:]D2+(WK8EEa\E+MBdNJV//cJVL<EH+S,1S2AUYP-dC:9
=7GeN>1;g;<UQ,FC7?-A73VfP-?AI:BL_1M.[>U^c#:]_J41Xa4E9.Z<F,^CK1T)
D=6&N&DDd-JT[UV/4IX:ZXa.dAD4#2RaWUX@\MRK<:?U64&(0W)J15LO=gD,X\S2
^8?TEK1A4;WPO?Eb2d:+###dUa,>,BL(Y<[C)#SH=9/]UNI,+5a/eW-e^<[W;NCW
,;<#PDXTdG+Sb1@gHTgLJ7>87K(NJ=XG&)UKP<]f[aFbLFWb4<P/2H/P)ZBF]:\<
;#6^a9EAH>Ob-.7cf,)Jb-#2bO2F21fSQXF6SB]+TdFCMS4+C(._)]60;@\R57;_
M])OBMX7BC((0/R8,&gM,E[_2<0KHU[>T3PRH=CXI,c>LfQ]18H_E/=XJgY2QOHK
@0(1aK+D;[MX^fHE--^\=WVe4cfaM)f.]Wb2Ua+0(KZ6R[(PE\+2T84&?bRH<_>e
_X],.BaNY7F;^VFe9YMHcQ\Hf&39XJ/[>fRS>C9/(JDE@MgHD@O?49^Y+EP4b_#Y
6=&K#MTI-OX:5Yb\6HU=4BLOD-\5::+RIMB?1M;5MK?GL9NPWE?O1-[PKc;7M;:g
@4O)^Wfe=Qe):_+\7eV87ZLLJ5Bc,d<O=GNJSX#FXUG5ZK=>XfSf^7HX)c,f>VfJ
,cYN?fdH=;/\@NeJ8,CHF#gG]Q0]4E)aDV-N(B(DRH^O=.fUbb\@X3>@6gJQ1a+N
Y5&#L#_MT?WGb-gEfgS+7EG,f0=-/,fPXKQ=_VfWB=3LS=5T04CPRX(Y=:04X-4<
<[X^7@K-#F2PBbbd\CSaOC5fgb>WYZSG/aCL.8V7TDH4K^5^X-L.NMHgL1BMG;Z3
?DU13e@-YFMH+dS;6_.@W[T0,+C=EGKAMWaXPXaQ@f]NKURWIG<][<NE<[,XR<J:
>):cH:?CZ3^GG6>b+MRE[D(,:4MD8(Z<[OX[f8=G@KDM4L<7I1>8H1.AXKK@_&LJ
[?;6R_d497YF\de40\;I>&T[B[./^XCRf_F8@U\(QK8YBE5C-/-TNKfF?8T,T.34
\?I59_d2b2H]D]:ZAV[P3TA;--B?DG<+V\c9,Hb_X&^&N6(Eg91W5DESdT3;4G8A
<+@(L-<RP&RF^LLK@_c)CV>F>U)?NY7KU#8#>&>bG8PYFUL=\VV#b6:=Xc75)4]S
L;=^&5Qe&](\(9^7<?/Ja&;3^Z:=ZB4W:ZT/;>X=BPOM^U7d2[d,D6S.0(E?W;=R
4.SQKfW)MCYYL_4Ug-<Ta(4FLTN>WHdOI&La6OPDUVNcL0-ZD.ITL/WE.6X)#(NA
ZPCf8WH6Y2aR9>8HBH9=DbBIEBK++Q./Qb=VY@^+3GBTNcE6PU&29/(-/SM0-;>G
8Y6a3D)O-:c,\IY/+6_)^c1<VWTVKO8bcF,@]4QE8H:Ib/KaW<DRcgGa\J:@(/<]
[-+-?5eYNXO>N26V0#.[b+F>(LO7\8UDWS;:f7C,-+FHD0c^BQ7O\\?SU(>a9R:d
0(d7@f/C/>a3/e41e;.cXbgK;Q<G_M^FO5XQL@+7G]TQWE<P9PdOEP>5?;1[UR.g
MP_SW#-ad#PNKabZ8eEO(b^f(F=QVV<#6c=D)V^3>@a_UTWK1_NK+QdbS_9W:7<@
>Y?XVA3//PDFaX.1V9J0_Q#S,ZSK@&a249S96<aY6NfOSMED+FK=TO^c9>?OfZEE
+BfY61MUH4G+<KKWCPVPg>BY31/-CbHc945\8;4;U59K6-)?W;36]-_9U(3b>L05
fGb>6ZaeBEFgLK[#E:RQ;^=Pc3\]Dcc/;7C/;U)AOF;7SZTG:(b_[UgLZdU71K7)
=02>>F5K&e065?U)AP3@HQ442<L-Md:,<ADHY\\bU.>3;;]SPAcXMTN(R^E:?e2N
;#>6^1-.T^&PVbBZ7eKI:NfLRR[0W;H@I-5B=)C:D?Yg>fT>c:>d6(4)+]Z2VZ)Y
G1:MeBWRE8Zg:YPNL/D9<NK;[FL?4I_]G?1YJJDOZ6U9;fP<4<_0S[H?_<<EHNde
N>-Cae0Q]a_C+61e2<^,gCSLM(f//9I+IP[ARd6gAIB^:T<].,YQH?8=[&OaGaHe
0g?RbZ(U.BL\@0-],WEd0+2__]/QcHg7@K&&K29#@;>E6B6R4f3U31eKWbcLH0XK
][]d+_K)<\ER+bR7U\^dTMP)12[<&\XU.0U/N#V\OTT:XAb.HYNfa_Z)7J&#UZHb
#L#]>^a5RQ6.2@5./8T=1T@2Y4Na]^cO_?g23HXb[-P-L(QD^,LGg7LP@M@##HVf
1_I6AAA.X.V,)>;1XOfQTY;A]-=g#[,^?>1,2PN0P@Ue?fK=JXG-08E277JC:;M>
B7N8J@31P+6[<FBBcXYaLECUXI/GLMCNPQ5d8Y1JBJ<0)11LeBI\4bLbP;40YCc;
=MKOWcK2U9:I6><#6+)EYVI<1=L.4.IgCV2Z-bU3=2B;FBR9L)[+KA&G6T:^OYWg
N#T066f(EDI\COgdS[K2IY3-\M0cR+GfB2V9CLCGXeQ7P8/UN]TfT2;N>X8\Cg,P
92?=>I-E31\X^-OK2,3PGdY5[VLgc@960B4d6-WWZ.L\QX&_g9e&K&gg2Z]&9b^D
a7F#1R_OR=)B^V+c?O=@E@bG<DKgL99>TbD1V[F:92EPf?.8S9QFOQ64;WA9f1X>
00+P5Q0_cISdaHfF:3\S?X8=MT_.;N(E=],M)\.gDV\c6f)LW6ZQF.S?fRd26;6:
#e4b2Td<>2>L6;;94TA,7BN6P7&SI&#A23J=9S/@d,=bIY)dPOZL>7@_)EW3J_#C
]U3XUL01Z=FdbJ8e)C#Yc/.VHU0fU[TC4XP&:CQdK?Kf2U?Ca9<Z7,HN4gV]bS6/
d/P.F6e,2MdH/J:(AF=-;LB1(ScC_FE.)<.:9ULXb,_>EGNf4U)K@8=X:aYNaC@(
P(]^L9f)-b6f946@&78FEM=BG91ccFK]&ccX&^QMP8b<&gNM@Q=e;^/B),da?.;D
V)):WXLZGRBPIW#P8K:[c(24c<.(7E575^RV.a:XRE.7aTa[d\2]=J<Pa/^HR##D
V,,L7@M=>c42[HVW&;0.gIV58RENgeCSIL<;cDZ&6T])M#[c.B@WeQC@.aC@e&[(
Z\][R+ZL:XT6-bWWAeZ6\TS+&9JW;d6APKYK^Sa;T_LZ:a5)TV\KL/HM[F#?/^K_
gZd0\_^,WFQSfb;9cebcB0;;\LgYMX1:]24-TK3a;5S,\:fT:@@.F+f,B(5[=LZa
d7GNX6)_.SfN?.[V=2PFIQXCX1P,YOBN2/E&V(He1UV-\TV3C3/<]]DUUcbSPC-e
6D;Md)g#2dJ[c:?#^,7G7)P+dZ?g_V-U>T#_<F69&#(8;M./f,Z9,K.R^bf3@cV3
OOc3#YYZGJ2R(/4OP\I>^IBZN#D#@^/ZU1<ZK7Q)]7@\[[?-4eK<+7F4WQ6-USB,
R61C45>4eeEMQXFPK6M3<MV>L\()9bP:,a2JKONF@<F?^NEa5(W_Z4PZa/F1#Y:<
D09_gVY8:^)gMaPc))>8E8XR#ZX,VDFS#:F6eUfUJ#RD7CJDf^J7>=G]U[T8gc0I
9_&g/OaJ4BH[T1B+91f6OGH&ggHBU)O9b)<@c\c9?C.+K^&eQ;P/3G^9?(TeTRW>
K)_@eKCK9+7a7d1fYgfX[,4,+^V7H-3>\K.GVCE).cYL9LYK0b@=47+KX,04\&@V
bP8NZ>g?58A#P&:]e6ZVI_8QbFKf6EbS&NLD2-9(DCF\)@8VU@Kg:3,770-.3@Ff
;^@GBVaFaRGdLQV)g,26EeAb1XBZISV6_L1^=C+4FWU&MSGXW\Bd8.@Iga3Af=6g
I@/.2bRQ+^a&_Ke32:@F2&R)NXfcEO#g.,G;aZBAMN<Tb9W8.9W<?JSOG>I:=1\G
/=H^[E&cUJIb&gH6Y#d@[6dMVMJ#M7024@(c5_V<-5WC&Q(f1K__0Gf:@<5:H=()
g<ZY;8LL=XRfg3M40,UTe;&XIMf<&@.N>B)?VGcL&Ha]6]\RX<8W4G/CJEFZ7f]:
KdJ8I;9a5d88DA2MK^d8Qc+K]IEP_eN3QL<)]Td0HR9E:Z/DY+1.F5>g@DE:?c0Z
KXZc^#6H#MOWLJ[M?45U?VF(3IfV<)[67;Z(0RUa9]>a^2U7(A<8adL69bT.5PRO
;\eg-R-UcGE[2&M@a8dAYPEHGgWgAI8.-9YOSZL5R:dD;EQ;[]:@J=Ee=RJ@[&/1
9\/,,3dIG4_<0BcD\D;d(JfV)<NcTRK4?35<X3BQ]MT5RE:a1YDAfXH,9=\85cCb
WG+YT+@d\WFT>5,,H;WOX?V&FRRd[f/P@C8A5[@dE:]+Be&g:-&0+-Pd+0cE+O)-
&DIPeW<GI(3af)Q-C+GVT-1I:cLMe=&a8DU]ee-Y0WHfg=H.7)aQSKO5\])ED<_;
3dKMMVBRWG=UE/Vg>?J@73^ADUOBb?NQG_,5#Q[@XV7c^.eEE_R//UVgEX8gNW:E
fVgA0VY-UI>dP/NS7^6bQG\d129A9;RH1&aUa94>8WP;U)=&c&1@3YE]LU/B[K.4
/GD#^Q3]Ud7?7\F,TW(VO?9cQ&@fKd7Ia6K[.36=?VS=]A,cW,M7V/,Uc#ObMLJ9
O=W55J2TU\If-F9WLQY,NRVDZ8BJ&(g#5cJXSI62+&A.33OSR:Scb=M<AY_2&WX:
FUf2(.2W;I1=9D#(FFAF3]?TgJ^EET+^+3f,L9.#>Ra\WMDP4SeQI)Y6<\DFS,\&
/b)DRf;GZWVMLO63<H31efa].P7cNHH@U&L9d@+b6R:4]VdXW)L]>VQ?Jb(63a.+
>4+D8c_>.(1/(M+c;a(K.(4W/GO9d_V,I21)0B7DTERLW1&ZG_-+0a#:M8A,)]01
+4C;5YVLRIOXMbCZOZ7dcLf1OO+QYag7G=JM2P=^A1Q?=ZWg-6N4aF]OLb<FX4F-
89=H?Z+.d^U?Q3^3->7e^b\/H4BZ4Z;R6R>c-#9OKY5/Qfd4a##AMD.,#CEd4f6W
0/;X<L])3?\LYB_O]-,24Q>KK1CN>Q3=K3Ke0:5CW9OIK,eB>=cELLB.#9J<^RT(
@RD.?PSTYaf/5[4(GZa:PPN??.+IgbQ2Q)QG^A=5,Y1]bD:2LGJ4\_1_OEG0e2d0
g]@b&6<5cGa@LN^D\dcBW+]@^4_X1A:U^\d)CFU:0>2,O4W0T:feWfP#[05=38DZ
SJEL=()-<2FT7<4\6cUAYT_5@_JH&ZA-NL)dE(PaI4?>KJ4>c3<0#W5TDMYSP6dZ
bf8LYWH^gE<)]N@J[?97gIV3MBUa0\@1NINJ1OOFL2<J,SER+BdA\D^6K4;PHP]3
,D(>,JaFN]bUG(F?7H0W6Q6;3LR&)a?7:6&HB)KFNWgA33+67&>9b0-^[HXFO_.L
T8Rc>Ed7I,&[AQ]P:=H:/-OY1V33HWY=6fb=)b5gXe,+A<A(GOTS-53\6]<0P7D6
\<NQ.^>K7+MQ)CIO(aA_H\T^Ze-:#8VZe&0&8QeffN<[T25#ECAF_U.]/7da)=MQ
AYd]g>BW(>@\GN;\Zb<C/4.NU[].V<85g5I@]c=_A\(BNf8.QA^b-D,cM>/.Ee46
S,c:gLI/P(OU42eMZd[+6G0)&F6X3UYW=,)c_69SaX-&>\OD#(4)SbZ4Q.QGN.>L
Sg6#B&.L@64CC9bYLd>?NTS:K#.3?>aY;,6d.]K/Z6MANa[;2c?4\X?>E?8V9N+S
dMX;?X#]>;8/[#FRGHWI^EKE:2eKP@Ng)O::<G)+MBWG&L:g1L\-=^Q=E^G]bSO\
f-aBH-U#cb(6+a.B<Z)=TSA]EDVP-DX26ZU;6#++R_2C=6)I-D-=1EdBf:32,CAA
OCP&-J..&PXb-DPTb5#e:;9f4dB<6HQPVGSf93eJG)W_&(e6a:;<cE<4)K<=\V)0
\\ZHUGUU-/[\VfeW>0aM@A:OIfXMN9QGU8eUT8H==9?V2dcL\b\R&bPAg#E4>I>>
&KL?RdFUTb][4CTA4^#?XO)69L]6WV6K1HBgC^Age#.?E7:E>bG13&4]bD.OPCeO
fL?3:^5cMO0^b?_84<KX?La^M^TaAaMe^I@NXcR\^X]#JYe#-)7MX?T,84G_K>AJ
VM88L1B9cY=@c6AYPB-+KQK8Y\W#Pa4-K\4.UO/00@>77L63fXT;C.Rd:-&3]#Nf
Q(^B)BOZ9[=(3797PL])Zg\N\O0FHUWVK[:K&+<fUQcK,?-&(N5GRg)E_9a^291-
X]>W@R[9QD,.b\#GRRgPEOb,XV(2A08E3D?+0GD7T3Y6<_fU^EJ5C/.1GR[8<e5O
Z6\-Z7L:U9;fJ_A9:Jb,:/?c40AbC]Hc8\.GWd1bY^Ug(g2\CeWFcC:e-8P;QT>#
bEVI&1MI@TQe==:5_/^<VfCOYB7(;V&)2Bc<[e^XU@<=2d7daT)ZJL/5OM7?9g.R
A5T[INF1K&a>[6?2Q]U@UdNaYO+F#6N-9SFBF+WfU19fUVe)+Zg\;KSfSOdBNDCQ
b\gaR23&OBS7:,^2:JW.Y5MA2I=5YSS(fG^_#.EUb4(2@PV:?=Za6-5YDD:cW\U7
aAeR<]/_T9;VB0K57W7(?>Fd+>bDFc/C-^a9<O?DfP94[#L&4[DC7L3@,^JF(..e
fTLU_,L\WM@Q@Db?Fb>3f\SZ3H8BfAL<-0E-^/6@5V\8ZHNM+->MV9EA_6+3b[J5
)E8>^1c^^7FL[TGD/0[)fB@H<Z/<(8MZ2gLT[+R].9BT4bJ?ZH^)).2Y<[a3RHfY
E.X1;Yf#-&ce:Q6\2F(_=[1VU_E0DN=2UcaDW\<V9B?[II3F(bb(VU8S[6RP?-0N
X?0^Te&?AZYeaO#e9DDE4?YY>0++eT_V>fTA.a@8U3+Q^:=Vg3O&A/E0](SSG/+Y
ga89OM<Z4cDY;/=GTK7U#>PNg?[Q?O@L_33/4<DM;]IHB<AH-9AM_9CV,_M4J2??
6U2A\J.YOeLU8\55&WN:KcKC1UH5UL5O-F-;RP4MfFfXXSW-@d3;OKK?BM#?OVH&
7Gc>N;EO22JaJ+&<WK?TJ;BWM5)P@N<ASHU^5V\#S.D(HS7eKS;.P[\aNV[I;,H6
&1M;\NK)W8/<\&beJN])S;/>ZOKg+LJ13@TTQFW78A>E4^_HUU(==)QHV)Q?>#QP
J^WVbZZVA.=G,Yg&D71edL-Ne68?30e1Df+f>a1DZIK6X@K7I3B3444T@ZDPQgO,
9L1\DTA\T_1>BY:=1_B5+BAR&19:.GZKb#:bbY3&Z\S];aYXc6N0LYd+Xe#A-22>
f_.#@M4PVf)KCZ?cI+?5cPZbeZJGY+aW8,K9-\TP2:\R8AMcQ6^P\ZYUGc;U6PQa
1S][f>Xb6fMF)_b&W:ZbgYXA6T9G_<dF0A--QM,?dVEa;OMJ5VDFV2W,@AL^9ff.
(A_F>=-0UfQ+;K6YS3C&HJ(f2;=(D@1TPB?C9<NC71Y<=DKQNZ&A/?L824gS<D7^
HRZg5eI^+c4bT]U-D-K1C\J.[6^&6/gX^dD+JgELZM,3M>4>CEE/COMK8;QGH@7f
>QD=G&Gc\^(4FNX7IKGS>YPMBCU82XJNf28(I=AUA6gUZ)R971DT9OVfDK9PK^<I
S,1;9/4L\cgV9V#5DGF#OKOS;X&-cP7@0N0[\N@1:Z/GG#b-1Q2<MU=.Hf@d6C?c
1.IFg]f[7.>RJ<JI-WC.@T3_@X<R@EZMG056Mf56a@Y7(O)\.Z>9JVDTY&.74]DQ
G76R-RZ>TG0aW^a@7,YEI(QdL-J@Z+D?eJfPR<+b&:Q>cKd(GCgDf7\f]--7>G&.
EM(E;)I2D<XF_8-[Z;N1^cIgb25S8T?G8P-=Ed\aReW<,N6GJK0/53S@C#P,9O\(
_ONgCe(3V/=EHB\ed,&9((5\]E^Ec]I4)UH9a8LCY&GWAG=K#+cW>^U4^YUb4/28
-RAdO8Y]QL7.9GHK;cQK/<AK1.I)VYY6);-HE_[TB3T@DL6_CAGgB/I_IdH45S1G
AP]^HHG.g,&GNCUKEObB2MU)3a9-<d@Y/5NEN#CRfS=e>CL5,efZ7S:^O<YJa7c/
?dQLI\S)=6?Q9Kb#Z_+W>.LLBE7F.P4XQ(M:-0GB]be(V&D6^1^&^c&IWE[(&2AF
M_<U,EHVK@cO#EY5RT8EOaN3R#Z6<R7BKV2?E-eR0bf2)@7&P:C4P;CB&S(S\.RW
(P9I?-H\O+_Z65^R0=9AJ975B<NfRDJfcG\>^E>eGD^)g?[(dSd^gDKE<Jb3ZV5M
Fd4C,W>PJfR-aFB^OP6,CF^bc3T[S)1Y=Z#YaSI1T1QW/-d+_B+cYQOTHW-=9?,5
&ZW2Z#QN,fG4=VBK\5b1<[@,UDe[&+dNY[/<.50=fUQ.:V8R4g-\1Ef47]C-Y:Z+
Ka&53#bUPJ^MRG1^6,DGD&YJVHH#T]/?VHM:O5KLUbR.[@#E6N4egFg?g93L.\[L
8)0+YGL+P?\Q<JF>fO8Jf8MI1E#@&Z1WBa9?,c8=8\]d6?YbS<9;Q5-eWOX3V)bB
Z,aL,P@.&ZL;8DAc4bDX>EGY0<=KfDL1NE_S)c.a<R+/Q@BbF[60Na9TVJ/4M]#c
GH=XMSUJC)DBCYG(f=a9VQ;T26&2?N<CC08PWT@GQ)=OG6ME(O54@7ZZd4-Q=9.,
MOEZ801Ta<cW8NZ=E3_AH?MM_]a1X&d4dHEf;49a:)^+fB:C.NgbR9>GXc?P(1HZ
&<C@#4e+fT6YD2dOF42dO]:cfd3\F?SbRG__>\]I).=cLYEKaM46\S6Ab<C/ccV6
OE]7AcLg4=?d4&O]b_9F@OB#/9+_eE,Xf^9T6<-H\4.Cd7N##ATJM1N-6CIH]NN1
&dU[W#+@gM_d6baCS.M]1/HUQ0)ffZ<OS>0X&PCZfDg/Y(VSM]BK@UJ8RHP)V;W.
,.Tg_KO)Z>E)?Q;(WB_3H-EYI/&NC]X@aNa#3J)3I2K8<[G&+.a30,a1W&_A7PL+
EV1C6/^04:g4J/\<OI??aRDV.O]-Kb0++,E:5_JMd08GbEW7/+#^OM<(4^ZeR@ZL
..B2?d#9#5Mc7>@B^N&6+?(f46<PP&3Z<@Q?TQFB?N?d2gQ8I<FBH4#\BB6)KCF#
++=GW]??_0L#/3?-D?9,,:>cN1-f(0@eTd>=P-?91IUd)(Q+(a@Lfc3fd\H77^M2
)_&-T7DRI^D:=L622_7+OOTH8@fb;1+aYYDf>JW](4TR8cC7=YH02N.c8FaeP88Q
PI\G54N9C2^49_RV#:Zc^CdUVgUafBd77K6:,NQUCAUF2DXW=^Hd3,a^TYT7[2fM
4B[E9O^?B.0;\[8[bMA&@=:@c^RV3MP[Kaca8]>/]:AZ)2N7Z2Le?]]NQA42&fOG
c6F)3;dggd[G4&4]0-Z?#eJMYIYW9+LSK,;?N3V-ZCHOL--O6d\>RGbE#ReFb/3/
c\/RZJKHC?JK5K2:.Fd-:+<=6:E5Uc5U<3,9;QD?bCS2PD>ea3&LM)0]BRJA;\C=
M&^-1Ya>U1OZ_1SM0G_<//Q[C3.8T]<S?R5[-Rc9TJ#>#W6PbFQD;8NRd8K9I8:.
99QcG#,FB[^PW]LWPA74AV#4ZTbdMN_OefHd18II-Z[d?^<&H=H?3]J=f?22=42M
H[H5)P6W=:6=-<>a#g;EWUN>4V^5OK+J+F1B@PS6+M@KBP=O1/g+0RWbGB(Jc?#V
NbA>LV\396UcbUQ3R?NISD_I5Af:):9P1KPegcF[E\:1HGEH\#UUEM#4LK9@^Mf=
H^P=agMW0_QLIKAKWX-O^gX/a)R0N/8ccNF^FT>-d@4FI7&VgGZbX6D04E:]FUb<
LKaN.:fZ8CH^Q?3>Pd#G=X#TbY#M>>&fKAY59-4@PII(SBE-:ADd7VPL/,AKHMJ8
9fb96f-<KRQ0dVGU&U5ObZ]IIY&&<W6)I(HOTcg3904)ZEd)J\]H=902HD/5J;=6
##=C\)X[T?89KE:T4f\^6Y0@+Sc08DF9^U2c:O5-T-)TN.GT<1a^^bQL6]3M#.ZA
W_J3<.^IefT?&R).dIXHIfL/W>GfCE0ZF_FfG8Ad-K#_,(0A5e&02a6B(gRBL:V>
fZE&O+-GPT9>UIEcH-d>eXMVeQN>TQKILY/^gCB8ee]a_G7\1W8?]YF,K8A<GO7P
D^I.A7ATD)33X<Z?WaV[^R\N;.PG/5-b99\>eWeO/(9PX>)baP]f547.I?I++,X5
8>VW^=Zca@+P>C):N@-I#_,2)MZUC.B3EWK3<_FJ(bDY@VUg+@bLQ;OYL:X)AF]2
^/>6LAQITg;W180EO->0GReW;IBDe+B^;=#+;daO\#<ZU6fB?=Ue\Ra:2Q]Q\cH/
,U[a)#^_UY9JTaA->7Pf/@E_b(GY:c1;V&K7AUM5gEY-M^F(7S2g<O&)^CP2C<J5
HQ(2T8[3TWF_:?<0A/BeWO]PC->&Y@a_2>cDb^6Ha=[E8RcVY)XF@<XM>:90O^J4
@6-f:f>Gbe7O59FgS&@SgI<\E&e8P./T2=Ce?^2+gF]I28IgU)>D[+NPESeBOW^C
0D=4?HEZXH>E&QW93,a5cJYCEXQ<KE?<-Sc<=H?C2[>2#D-a/P(:R:LM.bB2GR6M
F_#SVdW0&C]?_G]1\JC1&.XHfENR.=P8fIUc?@L9\P]Uf6?Ac>_SC+(C3LA)NG31
C&LH3eA=)dH,9LB>(H(eM+@GFJ&@f[]W0GI=g[K0H9D@DR&U:)OcD8#U.dS;TI;;
;[-#1ZPNG\_d&cZ(a<@g]A5AbbXEf>BW_SG,I4^;L2/B>L5VUS^>.Wa]g@#YULBL
L\f:4V1H)LUM<(05U@BC6=U2L:&[NA?IfI[ZGZ\Y.36XEdQa(@MQO;RZ^?IR7J&R
aL77-KGO(7KPC:F?WH1[@ddNgGfXE#GYX@3[M7;/-U&L1U:dWL@RDXUX:^M/>W/&
NV_?H=ILK?@4f6c[EL\^(7C/.:R/B_CObb/;Qc5J8A@ag.eeE<OIFdIU0_)P^JS^
Z8K)J,]<Ze9_6JQNc&/cBXOD?JJRMPK6<8I/M=:)eZ\&.6D2ad@+RD95Jc=?HfQ#
6e3R1McDTM(Z6[((+e@-gd]7MGFEREDG6V/R2G)QDM[]B6N4MI5O<;G70+eA[8K)
HBLG[Dg@+E?6V5fW)dOOc;S\4LPLF()G@5&B-+4:#71b_Cf=S(S4F@GQC@@QQ\A+
YCf14#2_T?YTcF.S3d(NN_8B1BXP[]ZP^-bU=9B89,-aN1g#[(X73V]ZLW/(;FJ_
OZ4dUfQ-3P_8fG:[/W_R0.b.H#7T:@D1egD?F1(f&=(b4@,\eOeARL<-d+.0\U=I
:#S9#EBAeE/\a.ZefN,XgA#486T,[HW9TBYHQ@P3d+):E4>T,9(<EOJ1:Z=UHBGS
-JK,U@#VPNLB_WJMR][,W5e@@W8@JN8X7aQ9[V6[=VX[Qe5.Q<=Zb2=](+f^L))R
?GD&\XNbaa_>X)TMWE=c94Dg&^>9@O)D?S3V@ZX_bf-fA6>>PW93dDVS;+B3/^TW
V3PG];IMKW12]0XW[TDKEGI,ND\25F\MWO<_Q1E8.+XS]<ZF0)-CGS:eSM[+P.,3
?e&MGWEDd+TV1Fde#@Cc.aRVT;3:FDSEICA28]3PN_-0,J_aZMWICSZK[R&#f/_N
O+SBD?Keff)5>ff.;?#K+^).=]Y=@;E4(9U50MD+;WFZP?)(:K^K;D683(Ma_=NK
BU;/QP);30<c_L6=8?M)<[71ZbINe@=f_(-X9(fb-G_eV_L.Ba1/68aC8LG#fSMW
(K;&NRG0JN:bWK8@(8)B;cAO7ATBNDK?9IKA8-408U60-66RWNIg#.G#12WHFVG3
GPRDgfW_0c5[/)+8_aMA(9-N]D>&Eb;<VYC7-da&,>79eID5DL]dc.NEg<>8e[(Z
E+RAcfQHK=YHGG0_fGG&LMUMbf#F6ROPbNZIBM_-66PN@5ZYBNO/_9)0AdO^RZL]
4#K917PQ)e7H)7FB9_IGK<S@)HP:A^BEb3PWB^O,H.g@6?RMc[MY<[f1<[HPM\;-
=O0D6-OK?YIJHRA9BU,@0VY^A;A-,/dPFF;]8R<-8C+?SJQ[2C,O(;?d(JU?],#S
GO63\GUY6ZcCYa>MT@eCe2#DB^#_Z@)50fU81c.a67J8KLLV-ag6G;0^BeZ^1D./
eG)T@[]M75FT#].,V:SSPTZ]2M:WBc-(DG(PX)FBa-9/V<?(,IgN,JF/[_KbNcB^
Db\Y0X;B?Z=96#MOM>e3F1Ca)N)(>c\=NE.cL#=P/P7C^X6)Y:K4LfM].78(P3bc
+#<aXDac<U=_2ROYRd9AL?YPc4#C&L@eL##cId=cQ2Y;M:bB6_68PR+^.T;UB\ZK
IGT6KQ9\V-R;Z>95O72c=DK-#0;L.;SWDbMM?FZZS\1RCg(0dcS\J26GWG2CJdaU
Ge,H)?EaJBMA^f3fdBYYT@.=0EMMfRffN@MQ,?/f/=XTCWDK0@3Sa9B<&Ra0Nbc=
bcI1.1JCDS<Wg]d)X-fW<3CB8bUZ(R4Bd8K8AM-d4/UE.+:LN4L\A#g6WEd2VPI#
+Y8/</Mc4X=TCR,#.O,3-XaA]=\)b.-dUf01#2>fE8V9,GO)d/;S3@3JG._=)Y31
e:A&)]O(PWEMB\.M.&KQbeEP7DODPST4bGDdAUbW>C6AbRT5F557IE_73MS.FNAa
YBS>/eSVGH=-CY.WRbaZe[(V:)Wc]T\KQO?8H3d@^B4=IIJeHPW]:OP>CI70bAGe
fEc60+b@WBbc;RWVCH/,+f#0#BM;@^?^&B]JU/a6=\BE:-/=\feO^)A<0.C+5&?.
c1<\<@>PZAFQa;ed9E,3bJ[WY2MAbQ)beGE5LB:&GZKCF)V3(F+OGRCXC=AA^].a
J=NO5JFBdYE66XYbR<C#Z/&>ZIV(\Q6XSSga.E6(9:G3Zd6I0]_@XDQNb>G]&A[+
H4PX0bc/f:D4eb\^4GMZB+_T;+5)\E)1)P3GKZG.K]XOG8Y5E69-74[^3Da)VB]&
E?.YVbU?+7PGDCaHAK531N8X9Zg)L^HF)fS3&a]cZPXOaW&?LXDX&fNK\d&&D,5@
\^(fG+PP;D-8)Hc+@)^J:)K[8<UIb=U+MJPX]90I0eBW:&M7#c(R#]7g.g6d-bDX
#HHH?GJ5.U[&g?UdU[W(A/\43-R5WVX:7B)dY+#YDA)g219CZMW+X&f,?8<HDC[,
8BH7.;:R7[RI+2dN1DI4IIZYIZ)PcA\<6&ag7\[E:JQU<cKFeC2W[+WXLW/-,F&B
8G4&I,2_]e4QL=^,fc>#D&eYYHI0XA&FT#;f#H:J><f.=e#=3HP)9D^6DbC?MY1-
VQ,:5IU<RR\>_;57H)]:<MLTT+XJY6\,C,V);e#?7UcW8UJ^78+OT4-dFO^&)Yd\
T(2ADe,+aT#6TfAYC7UNP//U+::;BDBOgaN(3;MB=@;f\8<5=,5=#c=28UOHdJ0)
gb44JMS93#_0_Odda7R<?fd.D/@_gK1ZQMX3Og,B@5V(C:=-@OY[S<LMW(C=g,87
X?<Q>@,EFFc+Q>_7(YI.6YgH).e)>,>bUXWe,ARH,P6fLdYe1<F]/P39W=A>U5A1
0T_CO)2^_b[e9OGJ]&,V8LF9P(K:XA4/@1:>eaQbgCD]S[IVHfcbN9&&8X90>K#^
RY)I^(E6E4<]eI03@XI.Q:;YBdMGVT--\Fb>5#0M=5T6bH2DbHG^.,C]?E[G(8b-
HC-f\OG/SFA5B&-0?[^ZY3+a])6\71:Y[_(1b[+;E@??9JG8),M\.ZgfV6bLV+FO
5ObH[H/<9AfZE)1a(MCS<JE0\79BY<7-UKQ2e.37RF-B_ZK:61.AK]U/Dad^J.7_
V_^-8^KQ.QBL)-bY:AVIf)\.CAZX9T@#FMNB4c3gD?8S89fdff-:7Z=<DA3.#93Z
D?:>>T-cKM+6-X97^L[(IAKZdV4Z##3,FGOZe^8BM+LKbW;-B>BV0;9;7]&/]^<J
R0SbJ4_?XQN1?dPSGZVf=1.J>Y==DIS620N#Ce>H+FgR0_(6cIJ#e)[4OO&g?&;S
GaA+9fM5G=M((M2I=?8IPRO)EF^:IM]S)\Z>[7J@X1OW[2F-.cK=g&#G71[/4E[0
cO(c(DE1ZVEMZe>-@UMETc4_R^>[P(6I2=a)\^/#cT_Z96c4+dgIb.dRA(#E3)f1
eJgdc[R_&JM4S=d9HPabSZTK8U;QbC#ZaB(2>]4?D)UG14MQP@0S&I(Uc_56Ca=5
d:DN_=\#.>:D=bH)):[CaJ<HWLT^UF^d[>)YJ8TFYO_5LJAg+K-[3WIL/T616/3X
-7cP5(#-(.1CRIW03_P]d?]EPHMLLEON&TgSSGcf,a6bX1X>0KNEKaD>B/;YX@U?
E)G29WBf;bF2O_.4e><,NDe=\O#G=b9]V]DV=-I8D,_HYS=]a@O&_#VMA7<@Y8K^
gg1OZ&P,>_Lb9,P-9TF#+AKFKFIHdW0;L?0SdB8L=^/UH9e508DG01OPVB8U>I/&
KCUZND#2g,A0]G3OI3]c=0,1C@0.Y_PCeEN/X@SL\?17UDB-?O?]NIE=J&<ZDR7-
?4c)3H#aR^)dd6MU+3C_>C?SFcM>W>R@MYB]@=W1D@TVeOZI4YW<FGH\E9Da>^(_
JM\IHNRb>_?0ONg=[.EI^JBGRP@?DM,/>1+OA-aG=6FROUAfQDK,(?,_T<#DaYD_
8+B&ET2]eX(?TEL0:?L#N[1-1PL.IZ=WL1_0V/X1D4A08\dZ1VAXUA+<MMWT0YIA
9X6;fWe=N-LPB]ZFX.f<DCET--)5SQ<S3:BaU(P>=]fTT5NaW81Qg=.:LPZ^/J95
/-<X(HHJHYAR@.5U;553TA+X@/^N2^aG2@CD(9/AaS;HK@+c3Hg8b7L2&)IWggc9
M)RY8^AB21.]2Y,,g>HQILF;]014FSF5=C:AQ)BeDQWD2V?IHP+T75Q;,ZUBIOA;
PXT0-//(a2KK]=]cACP#Q.^LRaI^.fRe3>><KdR#TA96bZDZ2fQ^D4&F4UfK@=3.
Q4LC@245_/S=I1I+;^XR.<3[Na^^>WW1TI7ZHV9g1-2<_6f:NU(8K_=.T64)LJR/
XOE7g6E8B]5XN/bSJgVT1-U,P(L0[H&@d2)?]2M5>PP\+S0Y7\T^@)a,;Y[NS]).
HGEZU)#/RAK61\G_b#-a,T@(b87PfM2f@[SN;6OT3)79-2.FS779E)A&C\TgAdN[
U>36O:[R]P.aL]L>OKR7f#UH^])S5.Rb_+H[NOV:SCbL->TCM>OLZf/1JZMQ+DGB
UBJ[dES5+eI:^A?<T05E0(-&a-P0-D\[-d.#X_]8AK>U9#/3L7OK5AOaKDT(dN_D
I@W]H,K6[TYCYEffT)46[P<B5D:^IMEYX80IGH;.f/C7T\;4W0F5?e1Ic>cN?DHG
g;YMW@?YC(?<XYV:F+,2dB+a/3RXeDXA/I6>OC)^CgC(f+VN1AYa_/+E?B(:c@EQ
>O<UFK+8_=R&1DGcMD0RHfOCOHG[+d@5&3H>X6F.GZJKD[M\R/\IT>NW0:.e#]9I
EE78B;8>b([Mg=9&24.2J5fC_6W^]fCcR&U7]/eVB6SO2^\(\FOPG.fUW?OR6]2?
a(Zb&Z<X>TE.=&+fe>4,d7E3A4(Wa<e#Q=L6Q7GRQ;7_4-f98e&Fd(<5MUTU\XE.
N,-XY.RN5_?2V.QPcVLcLID=34OK50Ze5VUf+POfI\<X+98<2IBb#SCK&3Xd##A+
5bYa1(SITK>P^+64T(7SMK2.71(Hd,KL^J/RZG&)Ag#-f&dM7,;GQTG6>4d^6A:;
R\]W>U&LNbNB[I6d>\3YC.;+B7<,GT-d-32]K&H:d(8-aO]LDAPb_DHLUgDI)WSG
5NB,N4/.,?[T,K._,c#\OMHLT#A@0PVQMdVF8K)Cc:A^)PO@UOO.Se5&43RCceCf
[1B9,[ReR(52eNb.O#aHg-93S5Og,GA?F75g9RbYI;aKMRD6.WA:cZ0e;cBH),4E
cSLgNf&SSbML]_X@c4@6,e3Yf>WN]e&HEM)Te-=b1EI0?Z;5a1&NTc-,I:6BeD?R
T1P?.;D\Qcf#,ccQ(:a?W\+BEK-\cY;QM3R/Mb)f-LSaO@5d33]/.CO0\GL<HK-@
#F4a37+dbY.M8T+@0.#4cQcbB\34Z-PPQ<B0/5<25B.aMUSefKDHG6RQV\[L\SX,
GX=cVdX)D.&K<;J=fR3DS,EG=4&.,_]#E(IB,<JFN:^I<]=B_-NL8(WWU=7\f7Z3
Z]F4WJ;?<]U#=X]8]^<VXFVNPU\d&;F3;FZ]/32>#Tda>DTVEBZHQJ:c>KI9:;SZ
M9R1@B>[>79_MK,K6:5M.[=a4D6HBDCf<^1CZC;5MXVF,=:)H<R11L])1[D;=3).
62BK&3/e6TRZ7X9CNJF[M/(Z^M#J,M^OWAR;Y+.]#^cYS80XCX?6),5cfd/V1;^c
6PE<T4:Z_AA=IN6J^-\39W-(NE6faF^R2B.:GVS9BY8>\\^GCc_GF-G<WFSD==RP
8-@.F]JY5K?^<?/\0#&BQdb@ZGXG)=Y62fM=SK:0+A=73,&=1,&T#/KD;U6Q>7R(
BUPIGTDAY5>BMNE0\XHVFC#AXC-FfM+MaBC/^&0\T/:8c)Xg<;,P29?/\90F6\C&
>1aCF94TW2#M:-_G.G7/1:.5@7H8M,=TBDIba963SYBV9@C<L(aY]&ZWME]M#<Rf
g6a):8N4C\G>F_)f^),=7MW,W#U2(W?a1&M6<f0V2@_@IDE)OF=,-AC\g?+V]77G
-/@5XU/S)d0ZE]-9K@c.f,342_MK(_Z4eIRST()3S\5]gN84:f].X[+\0>K<L>[>
[7^M5=7YRaSVI58Ne+:e.DGTg#-(+27X15(=Pc\aOdPKNMA5UYgFLD,dOfeQ:(1e
5d\SCWT3b.Yg<@2aH(7>(V]\2JX+):IN/<[NceIBVYeGYfA/:HC407=^H=17JUJe
X+WdXF6-49d54K8cQfcR4.:.d:TM^e3.Ha=cPY&>FZ?(BdN(H3+9EJ=W,4U66&ZG
:Z[O?_0a[.I#bB,,,]?T)+#R#:(#BT#<P:(F(59Y0(31D<-F&26XHWOd<GaMZ0QY
Xf-_E?/Y-F?^J[KDMW)JT(a-\W=38cfHO[)C]1MS=B<0FY7)\eb-\)KF&A1.B>L@
H^R-Zd@QJAWA))GM37;]V_;J9ZSUfe=&K_^8/#eKF#.g+Q:/3;Z(/OaMNIL7/;Pd
??@6g\8&McR5A,Ec&+/&7XICIRX12HPGbUbW2b40-V(0IfDL_.S4#QZHa#CH3BIf
3]VTHZcL&_;8,_e^YH;Z(?DTJ&BW.](:EBgA;Z&]MPM0D$
`endprotected

`protected
gA-d)Cc19JTPAgOFHga.MfVeJLH)Y<d2>)D/V[-PJaK<c].2\2V62)MVE3KO;8J=
I]G:35]2-FdP,$
`endprotected

//vcs_lic_vip_protect
  `protected
G2U3_>IZ0RM43F58g..9+6Ga85LGY<9+.&CN;QS0+f4c_5-J\&/M,(_81fd=771Z
a<^#b1I+g1(Bb3LBg&Zd;>TF2LP:C#AO\N-C1^88e=VC@PgIgV\I<CW3@_(d13TQ
/#f\=_O<T#f[DK_6:DHQObY(aeA;TAeWI_X_/P+Sd=5KcgUO:J:+A>\65V^S=(&5
<eAQ:JV6N;[b(^bKIM1QMGZAg2d(@63?bH:(&M0MQfERZY>(5&@gCR-6cRK_)3\@
Z;)KWEJgP21NUa[^E^[6&+?XEV0.UQCa-]OCD-eaaC4F4V=&?[,&c8B<55FAFC19
U^Xc6U=XOY20+#@bJE2:_^/)85J<0:XYKG-&V&LG-(XJ2F8@P\L/40/;TG9?g5<a
dDVKWRfYb5Bg).g3g<cb#F)JT@;<]O)e4+#\YOI#)AcY@?M\2H69JDXKc2[.;7[G
O73d??KGB8Z]I#1[Rg8^KIaH78=A+E]\:a6>TIDWR4TXNBdVS/F5)ZIJ8f3PV;@J
^P/@gV>.]>[0W(1KgSWVPW#aBX0RXgeHVaGVbg0MaR1TH1-SL;c)EcUMBS(](bM9
E6J,;35#?J+R9#R\T2c[KbC[G;dYg(@(cFAB]E+=4IV7,6:EEZGWIJ>Z)NcN)Waf
.UU3f^ROFO/47YT0GB=(]AH4OPCV)eeCVCQ/U6X>#\<7c&BUCSE=YQ5a#&K)2M)<
#<3D,?EGET,J[2Ug:0S=/ATB(+D)F_M:53\5ec&NS^Qg6Da2M)HD<W6J,W4S2-N1
W1N,Le/9CR@c0dK?6?d2.^_.gEdTf<V^#O6PGDFfTCNeKF9457I\U9aEa?DE+.Fd
]>:Q]Na_d\K08S#6TEW#8F8+_7-YRC-[0Z>Se5>P8=+/>Z)T(PDLH:>8?cU^C_AB
VG(gQIKKWc-^?R&[[f\[YD15IHRB=N9O3R=C03J9)7J(U5[>3YQS)_GS6NU,Z6.a
)XIWHfN(f3M\_T-DH3UFf(5>,:&>7?_[3,E2P(<I>HPQBTg-,Ac0]CRBPHB)6FLI
KQJGI7@=SY@?B4b;D(F3I@N_e0H8FYPWg]\WU8-_?<K4+3ZBf=K&C=PT59-6L#ZV
TYggBFV/Nb^9_+P<40LKf2+1Ic^6EaJ=Ddcg4Se,WIeI1Q;BSLUD..9_=K8U20,U
8VQ0C-HON5B.K)R/3X5Y3C](QJ>2VfXTM>gcQ=&T,64:F-U(D8/6KHHXDeaKSV@@
,=Ne>(TPZC?LaK\Q+8d2]8OJZN5#&9KHH@a?28,)a1545JeLG+&FU+PdL7&V/K<a
d-_]CPY(fDZ,WHg[;CYG198)dYg<-5ALKXf=Ba;A_W1T6;^X#:c(f)OS]@BS(22P
F8a^J@4J_3:[D:1F])W<#1ag&/;-7@W2I+2FR>D9DA#AF^URT:)>11?]^5A>?@#D
#cN,Z]6cgU:_AbK=gN4>[F\gD)BL^.5O)4WJ(L>b3HVMGW]ZN34Z,E4(DUc@#[f&
>S>O.dCM;#2>;5K74D^+Q2^ec[fI&ePP-^)DD@.BS(K];JD-3AN5^,)N)REPc6MX
c)D+3/9I_)(L5_U:-#\7RS=2T9KOBF>@^X-=Z@JfH/73)H5[NDUG5&F6+WXRA:TG
eR.1JS6T/Gc\)MT/LY>&0ZbJ;e@g]K56-]EV&+?M;U0VfBX#X+fW&BQ_.B@I:S0;
9+NY_U6Kg(+=G(H>=&(FY3bUHZ\/8S@4N2[\H@ecCdeDQIN8f+RA.=2SfUa,J0U4
<Ca=-TIQF5X=D4GNH0fa85B)>M1//c>?22L^#U8Y?K<c\eR,3KB:WA>b_RR):5;H
[W>62]Q]=Vf@39]BM5(^5JSX)/bQW.UdMG2,3BT5_#WKW@Q7R85#=KX+=TGIfI?5
=GUN9@&F[XV0A^/PBB\VI2_#dO+2Q]ZdbRgK6-O>_1838Y<aMU[94ef].YYN6L3?
M1B,LFJE-SY)a^9]V[dHA08UFJ)O9?MN:<.H?B^HSB>@U9YKe;HB+Q(4)S_Za-U(
LAa45f@D-47M1BcJ,eD4Wc\T+e0[&cM_3SKY+88X)IFQE(_=10QHR0._Y),BL2J&
3WPKb:d\GW&U99]J&U,WO^\8]7Fd9DJ_PPQS-[S6<<A4:c-6=>7QC@6(g&X.b+fe
:];U/@PE#+^FUcd(ABRW+7bZ&NA#-)T@c:_Rdc(\_Q9)1_3dSPS[U_L=D&<.QQ#)
30[?Z2ELfOC^9(/1UM7bHZ,;@B#69]KCRgcZFN;66)#[#9WER:ba0gXPSD_:3?3S
@e:67RdYRCX=7T1Gb5Jb9SDb7ZROQ>TfW)[G-f-\DD=f;T47[NaM426:/GDD><Y8
.M@SLBdEP_PfDY@D=#N,]bCET\EgaSe-&SY9Tg^1R04&ZWdSaM9H,N31U\&P=@GU
PTJ)0cA+Y+TC0SA2Q3->)B8a?=B,gSK?[O,@ZVbBZ[3V:IB8X.2\22Jc7AfCbSWA
dDLXJ=bV2?=U(>?))IQQ<(=5;7FK:gW7.^<+XF\7Y)NZCH\,<8_U>ZO0P9^9LFfV
6bE^3bZXc4S3U0DT6OD2BCUAGf)Fb8g3bU>T_&+[Dc]eX,=a@1ZfbIIVM;/c:N^X
]44S<CS5E&1QZP?L_9dAQSWS@X^G]ZLV+)BO\I.<BdEW/C(dg.U7bV.^HbHe^6W(
cGbT^2XcIQ01A,bg09_.fA3bP7D65eYS:5X^;SBNV-GR.b]<JBE181)4+-DH7L1[
9baW3e@I-TB;c8//(YZ@.B7KKR1H:/GcCQa(=+[MQ3c3G[fSUO?gL@=IU[[QX9ae
FAb8]B-5N\4TKB0M]_,([bALYP^K:0F6W,Z##[3C-f4fD,,776Q+LW3XL1H5FGFI
9-,4K5fNb5c7Q2fP^H>\C6;dbG?P=?B-13__[S[L]3.N\gd-8F]G;(2?9d08[O<M
]:P4H>C6C5NDbXO:@Q#H-8-+>5bOKb9SQHBe5H<GX,ObZI2&3]B_gSDECL4c/=D(
NJ[fVQfc?\+()cAbC/RgY9/A9+9C-B0K(Ia3[3U[fU^;F\>3R32Y&\8STEBI]+3K
dX04S<X5:P<FNIg5e[8DS\:UId#Cd5A+NfP(:fG19E8?dO<3P+F0BQ,]IUgIA>7Z
=,dT9\Je/Z-PSc>]6(7^P#?&ce>]=UR:.[-;;;4>#(fL]bX=>O8)5^fS8#4C<G98
Zg-X-(BU1OJVaRGb=d6TP;POBAR_+Q>RO>MJd)5ea-d7,8@EVQ9-&R(,-0DMg,^8
1I\B((HCdXB#;@OP@I3&Y[TGWaMZT#-5[(?<]1T.9e5KC45F0Ia)JR</@>Vf0G7/
SZELWE:].2STM2_[#XQC8B8Va<Nd/QAA.]gb;;^Q99]>G,+-?JBD9]25V-D4;)5g
aC<B)H+_X1ece7:[M<R>7LF=^f3NFG&V-^MDJgI_#W)c+DSKIBfS<;5AV<E3Dg;#
^G,e5QY]g(_WAHc.-8_E<W@6M5&>+&W/faP@>.&RCW/2e>1WfcL_+UH7=#U0<OPZ
B3MV0?-,^JD9_T).eS.OYUYSb@D6XT>^g>IVgIAd^-V^Bc(;G^Q2a4YGKY0e)?Mc
ZX&Q1K]A=)<_)-P6JI7=&9WUS4:Q71NJbHMdc9RUD[&_N@dK\;TK=:.?0R<U_+;R
><;f,RH&?HOLXcBE:=cX+OdJc?FU;2Q5bZL;)L/F>Ld4#UJG/&g+@0ZHIQ[BGK=,
Q<)7-ZM(CMY5]8JRE[SNR7@7#DBD6)/&.CI?EXQg?RcU\586[8C&]+TD,RaCZ;J=
F>B@G.?96TYb58;2&<=b-6F#;Kf/eL3Dc.#&V8S3<]daQK,2BCe&Q<38+8JcLV3J
dIF/&##41Y0R<DB\.4T5?KP#\O,bb27[>KXYDYR@/9Dg>g^.FO>^&88/ET.TJ&RR
/UEFYO.b&;]-61][/\@f4P;K:<[8Xa:K?_IQ](YPb-f(E\J)?&^(dKGKEA3BFbE+
T5:+,MWgI&e/KQLg=Nf2,5]XGEPO#7E+6J(HgFfbCg/L#^YEP9D9+8RU13P+#TZ]
@d#c[=.:X1W),La,H6V1_f=MM8WT(GFA1PCf9-J-Q^FS[(?P@JV?c68)ZGf6eWJM
/F2JR+8_1F1++e/LH(MTQdXT:AbGL:S\@[ZM0dL43d1?+O-aebYRU?J^4,[0?+M7
3LZ<+RBXc^D0YYDdFg5NN=(IO-=GRD-FELW4U,CBKX,]_C2[(A0b>g3VIW\=&+5E
O9bDcVCRB^)89;1K]71,c,Y63RYQ(X/IV_;ZPFE/BOR52\7Q\(P?W;]G2A/bU>:.
g#G//b3cBGfB=[3,]T3K:(TdF\:a,.;JR:-^,#9ZCBFN+H6J1@1.7(A:;9_+-4P[
Q:OeM9C2aa7O__K3^Wb]=E<dDPYQC5<KJ2e.7a8X8=Ee[c<A/G;)2PY]K>9738VZ
DTP3HE4W(be&+K<#:DKYFH^\=)Rb10aabZ;A\96\3G)fLT\V_9_R#g[9?T]b6DN0
JT74VOUAG5-O:.;QJ_V.B605]^Uc2g)g13KO1>L4Q+ee@W.g&O4-8-(:Xb-9S,A(
6\&5:BMQ9.A,SDNWeTLZN(/)-#,^DVJ:>=,S?UHF_+FTKZ>=M32//I\D/G1Tg[GJ
a;Sd,\F/gZ.>XVWV@Nd&dPbF[58+UY5,B651c0Q09+SQf)gQHKUb)L#:.e4VMgd4
KdGDQO7bB>+0gFaIWO5LgE]7#WB76KM369TOX^g/1IZCU:dWKaTI3]e=ZdT(IT.7
/F8-(81/\D>3\@7LL;AU7gD2O99OGYb+[BK^bCRJg@cV_==#(,8;KPJ4/2d=O-52
f+XB_@eQ\(_5_YG>dU_FC(>)eV]IGTW]_;fg/D5(NVD>gG93:c9RC-f;bMg3F^be
&W(QNDBQQU5;Q;Z4>PdeBc..7R:+#Dd0Rd[)a>GcX8,f_SU-GeH\L[Lc:e=f1E7E
-dg2YU^L@B?bceE]SDTbg6MT=I^KU38D@7X+Qb,U6C#6+5&f9M:#5E+e,X_cBF/>
>Ie-I58#_,E)F?GL&M)5#@X^db88aQe/(^C6V439^)\RQ,91>/@(AEYPI(gYCH2F
+\I5LYO(\J<GcXSO]db6Cf0T&AS:?>;(-9gVb_)ULPAW0Y=(J=LdE=T454J[=RSM
PXEg\CEVDHWg]aSe^3LJg<a#17W2;+K5d/9]77>W>[(9@)J?86L]1]PA=9UH;b?8
@&2:UgFNS?,<aEEV:W3,53GXA0WQN&;&R@0V=fZ&VQ[bMeVOec>WA(2IaNWIH2Bd
O3[\2f>]aLD4O);I._BSKU8QU9#+=4=dA?>8KVA[VF2PGSDSB,DCDY,GJQ(NeU+5
/0a.A9\(NZ.3>+)RKLB&MV<f\bL:<YML-6U&)W9X8\/EZ&@R)]341NT(F-9<[+5,
.>[3</O94(>[Qf;U0LUY-UT\,>@97cQYPBc+)A<9(9OZART5=R40A:9#I4+59JG8
QF7+(/VFbVA;-X0B=8<,BQHB1.C;^0QQXAYU7Y+EfD@(S>ABaSRK40OfI^B_Gee\
I8]SVAYIB<[Ua6_HOfb,(.\#\N-;]C:cK[JBSH/fdL^NQC9]>,1,A)>9L/C27YGD
f&fHaaT)Kg,KdGZb8a=+CE7F8PO3SU6QBW/;L;4\/0>@,WS(FB\HeDUP=#0]7@WD
X6HWaH[0)(fBY&SLWRG1g^cJ5IZDHO:VP:cKCdEM[M,#VfWFFILW29J6001;Lf/S
TV^:>.0N0?M1V0FK3fLN.R,fgJ6L)^YP5Wef)HQXX:S73e3B&V98?8):c5TV?N,D
&T\EBK981K(4LO_LO)5RX-R5OT[a0G28Zd]C63U@a/7aS3EJ3QN8<C=d^C).[L)a
g2#G80fOG;.cU#>WZ6S1aO.&e-X5T0/B=.).fH)6HPUdM0BSb+6)8O97S,:<FN/c
2:CY?f@(2IUD6b;HT,LICO1NYd@>TBfOW:8+dLUeZ6_&(/F;AB.cL1]H@T4=H>+#
\PRO][a,0NE3MSOM176D1IM+dFNHM56T2&dLI+Bf/?#[;?&K(G4Y?8@\Veg+1NF5
ZZ&6#5;[\#W+KIF7WE([0.EQd8[?<=J2]^M(#DDNJ#/Tf7^VAa?(d-d4CFOKX[VC
ZbYbHd:ZA)SfbA5@Z,EV<F&9Y;0d:d[3g^Y?ME2Occ#1G2[,dCO-#3O7V-PL4#)f
N:&I?7WTI[W_gf0U,cZ4)4G7RL,VSN1V-Qb-WWM-+:4aN[-?SZ1?<UA_,aK&GQ])
D<d[<]QWE6H-gI[ES.?ReWHcXf3R7HaK2<>7?E=)X:DU,00)=P#\Q)WI3]0H/Q\=
=M-OI59ON=5U8O1OAYQb,ZKR6117:5ca/:80(9ODTFT;:L>@GC>L/&8>OMP-OJK9
1M9bNCZ.S+Q<^N_+cKO1c6(O=[OLEO.aTZH.9WC+=JeFd@PTf9(SS-VeA^5BH6fX
=L13V]YP44D#A=<SQ;&3D2N12-:,cXWZf3PD0Cf58A;2ABT0KQ90EWDaf.PG?PZO
J0NO;FTW.+KM0d>2T(S8(NF]8g4/1&H;UE1]WKb)_5c\c.II\99C9#&RC\]_:F6;
;O1KZ1[GO(7V,c;;(+/#+fgf^KG2;QYb]M6b+^fIL-Z\ec+e_X-7ae597eU01<,?
L@KJ,6)=],QCN,6g4X4H76ZC7CYZ7];fHSF+N0D2;5Rc\+;Ng,K?^UY\(UHCQG3B
?_MR7XYS?d+_eA-?^X7E(=EQ=WY]bcdYe3bP[[^4^<)E[X7>YLKXHK:2MP.B/P75
Ib-7(5U+>=;Kc/(,+68WPWNX0OfRB^@HfAda_&+_cI?GG8U^dPIdbM:;D=(_0>H<
K5JID>^&+O#NWXDQ<)[3N?-O]I&/12P(?bX;MYVg(E&UfT[?UX&T\7AR-PGee/C=
Y7GTeQ;VS+Z1-&G]N8#/G(_ZPAC8_DCRLG1#KA;?eK9BN31RU776T:.WF96=8]GA
]RDFU3(bB8IE?E.>6;FYD&(OZ_Y&79=9&aL9(bD\B=Ge8&WTe/K&1bH8\#X8J[G9
<^YfQDHY=JP_(;/43]V6^7:?-GO\RUPCQBU=2^e@;P2B2Va8S95IWbQe[R-Z/;.^
GJI(H[=#FU6F8_WR]ICEL+G34:W09aXB61.^<ERO[L8AUBEE)7J?U(>()e;?DdVK
CR-F[e0eNKXR-P4KE1Ud<D_];\_0dQg9RNM(H1T->?_Y=PU7POU0LA2[U+?L>AOJ
(,0OOZSAa;I2VDRa+3-J93(dZ8\JXO3.Af=,.^2:7e:e3;6e_>A-\SeX:?PU,DQW
gfNPFgW;R<@-P;OLQVEL:GD;<,V?KVRR#E7VU.XTDOZOb7K_GV[XBRI.[b?gM7+1
,U9de(D7FI/[TZX65.>)PI[T+W4;VO8d;-RS?VKXTc8,,74;5V^cLNOE<?P0OL5T
[:E.(&CDTF\>BD5VBA__5+3O@.[7We)G(YI<>Td^VPI/X#?3Y3=E;_WV618/BT;;
.LYG1LD_8XK.U93[T888/+3(#.XcLac6<2[dKQc16S0?G;8;/=FXfK7M-3(J/GEV
=c4O1<S7E[@KYY3VSN)Y&R/JR+CU<A]2IXYSB=8HH/RC#3bG4eYZOL]eP].]-g[P
-__(e4NbXPF)IAV,M91)Q2SRg;2,K:00:+eY5VIfY<aaBYFe\IaN;S#>7+D,Y8f;
23eISa60NWNH/N@&BG+K<[?8VT2&YP:9d@_HLG5+2RDYN,=HV79A.0][,f[8&&70
HD;2XJ^XAFO5>C74b>+HY(Y)V]gANF&0<]K_E9E3UX)4(1R-[Zb-Z@e^V\O41X,M
[c-ZIWM(J&JWSBTg_V.?].e-=@F^>-Z>13gU1?,JL[DPBS4CEHWHC&^g66LTT4MP
,TJ/I&1SeR4LI)0PXXD@Q=5KW2ZAX\g/P7+c-3^N@La&B):[OGfZA0I/6X-Q#=^,
e\Z5-J@?Y\&^YP1+6M)XAMSOLTWA-#7)Pb\@U1eT>LI9UKUWD>ZDRUW=IG_J6[4)
#2gH@CREKHO;c;FaB35XIX]L0VBa<3OE>KNPB)b969SO-NZ,26KLI=8B89aL]-_X
^RDQS@QYM/Z5(d8_L7@SCbMD,a=ME6S(9SI\S)gH-B:J^P1U>Ba:_\6F1Y<H[^+>
OB<)HW\N-3/2_SH6:OF+B1cQ.L9A,X0OaagQE1[BH\_D6-=E):?_5F@/TF(WfbXH
+J-g/.GfEWb?DC?>-M80\XK[B-EW4M/-Z]YID<5O?Wa9eNCeIG[fFH#cc[RB6//;
S1M3.MSYXP81eg=>AK3[Y,XE]e_W]4>LfKQ.Y8GSRM3@b,4gNeaBC_)W8V.ZHY;;
6Y+\QUP.:&NFa#S]DadcOcB/:fVB#YK^:>E6J\F6A2C8W_O97GGVDNc;):G6H?KQ
KYBUgY:cJ)K\HKIDcS?c6E[ATFff()6_VD2FW&?cf?/ZGH3GNQVcI8bPFVC_?ZO#
\+3e\I8R?]6cVYbBM7F(>5Ub,]<e6B9UQTTb9HUM;@K@SQM5P1_O0Q29F-b5f+(L
DR4Id9a[\<Z=Cf2>JN=6.9_KVaLB@D<#ULf;J,0EZKTYZVNI8(+F-2@9^>MdZSRD
A7c&af<ae,Z;E=X\dIQTQ^ce4>Y-bdF6<F/X9[WW:Y+64@=a5PVY1D8e8c7W8Q2Z
e[Q#XR+X#6[50gbOFP9/)U9M\[dYOYBTA;308Qb&g@4J](J)3A+TBV^b,[PT0+2K
V_6/E1AB+;1HY6OT+:1+:K<[Q^D5.I/B9\5YY<H[K?J5F?ZN(a8BB0(g4EWBcA:/
))K+\XYP^(JA&cdZ5Z&abf37]>1d[(,3fcOM[W?_A3e#@eE8_aR8?&.D&=@7S_8D
.\K:6:+.LdD)IZ/+C\<F<;Rf@PR?:R4B?X1M#-4?A9LSfJ4PP.[QPZLUgJIZffQ]
UXN,&G_[EER_D@HO96a5<3KRbPI2,#bG03-dL2M0\LGb-C^J\e1#=W)>D>X>IF8/
91P@&3^9)b96:6(=93@g0F2MeLf+5+89[b)?IK>8J^38-13:_Kd+P4YV/AGW2;9g
PP5;5WS&X;,<>dK-WQV)UL.L->B>O==6Be^>M#aA?3_S?_@bV7KPbC(/[]D=+:50
O-[M[C_:gPOZe<:&[^DHUOg^JNO3W><\TReM3I4>NOb)PRLbd,=CXdO=W?PU=EC<
KHLW/7>WES+HF>_4b1a;f]O=,KJQO=Vf:0=18\DG[&^[agMH(^<<6<de,aG[CQf6
T=a7\4b[LMH^(#<I[EMW@UecR_?_eTM03V4[eP7HG=MG(U1gQ+.B[DFOd[H2<PN5
P]dOP,PO#g+0/-.K/Sa==>2Y=c,=<<7E583[Kd7?K[V(-W5e@7b>c#,C(4J.c#H,
P;JdE1F.I8_J.N8@GKY6a)/cOD?1Aa\\XT[XXR.FRTOPU<N@8GNL5&+>DZ8Q#LXb
F_/dSL]<B_<Y)CHg_BR:.-41La9WJ;H57dYR=aK[cZ>b5&@\<X9fICg3g:8(eOC,
W85EGX=;4_.SB1OKK:f6S\[)MYVJX9^VJ[Y5H8;NcBW+f<R2H4-PF/G^cMW&PbM;
=M//U03T+?;[F5)V6AgT_f^,_PEFaGYIHfSf@,RF68g#JbM>,D5]X^1.4JdTF)PR
,-6-<D#\dFd3D-/3XHDfOTC/?F5ZLbQ;OHOWcV4B@VS@@)Q9gc<6(^K-X5RQA15(
JP5Xb@&68N50g&R:TEDI:G3JE^SY8(A_8@N1+^F,95ZZ#4:IO[,6&+)JP^O>A#0^
I+A<^e4e&E),I-)W?3G(24I^a6:PGDR1Z^X<2?K0Gfc<^\<M6RWO?C<MRZL([3f2
Y@L/121TcI<;eLSWXa:KLKb?VHU8\B.MU[CgLP_SS<IT@^FF?_Z1)+6=Yg]U?M5<
RV?=QbQ@Z(G=b_TggT&VFV18MTcMJ+.\-KF56cUZbY8;8MX>I;1cM#V9D[/a4BQS
;cP><XP&JV&JgaMC10J:-XH0ANWeL(_+aKBe;75:YY60?R6a+XfEDC-AcO=MP=&T
fOa[K2ZN-S.5?\Jf>_FTW7V<Rd5;(a1GWAC_&[_Y6V];<6e^aL540M4US]N33bE]
D(YI1-V9?4PQ&[;#]PE&RTMU;[VH&U<H:LbV4U.RaVNT[-7^ZC\25S#_+N3JQeTd
ERI/(>?N_J3&9Fg\5<0O+\/eX)PM)C_ZDBN\YCbK+F-R+2]aP1SRb8gP>@Y+HQ:M
@^5<47Z_HbHXZ=eOT0SBAOcMd_g1>&X<f?K;PR/<5H@D]Pg\ccZW-TXS\<9(cA<6
,bc&[T?3d2-c)J0];ZW@@,)_1,46&:XG_eX,KD=RKVU;&U;QRQg.&85:,RISNAEP
UQ-c#OGKH9SF6]05f[._O]Z:G&=O)d_:Y&.\<?1T=-#eSf6)1.8T=+&fV/7,F>_:
?[-\U]/Ud-A(fJ&<\>@/TSfYM)a:dK1HXMW7]?_W?LG1GDQ0NAOE@G-JY^8:W)(.
RWK]CWZ4-I\9]LQ0NO1Q^[J>RcP872-gJ.8fQ=+DZ.S-T>QV5]-J1:=A_B(#12gT
\4LZa2@aMW5M5gNfG^N_N\H(5\<_fR=L0O47E(ADZJ&7&dJF[C_-&cU5UXa/=M6H
^_V0+H<.56C5>3_J4dN]SPb=M(H7GCg@K>Y79@4U&bYD_BTLg21Y(J.5NB:?:IQ\
:KNACc+J1G.XVS+>KaDZ8)#;eIEP(NWMM&g?:2+Ib>ZGJ=8/M6T&.K8T=Y=KfOE4
M19Q,3CV5^Q4cVa](^>98KEZ10]VA02cA5KZU\1Uf7B:<cU1NQM54[6ZW3Y][EbU
TSROIP7@\=F+36eb5;A#>V6g&=K54W@2=_I,\^c6B[2QOEYNQ?C_Y4C=I_7JDY&6
]#TD^-+a^:>4Y\b^fB0d?28UDBF<WD-#TL]]OL9R[=Xb.@C\(@=#OcA5<[4,3@Q@
I4^C[6Vf<decH\_@fIP?PDceW_g)Z606TG1>ZWB^6AVH]GK7Bce\g-_?(gP52H.W
D(,JR.[36J?F[@8;Q-@>N?,_fO].B:5bD<.3,?UTA(>VJBcRU.EC=Z5)c555/XgC
9DK;Y>\(\@-.O8MP.A-C]<MbI[M>D6/U>=,Qg4DdGT6/]F9f+_f0dc>LHZScSYUF
&Q,.T[QP6Fb_>YA5Hb5;A)5@[OeU6[RaQI5F633PRW_(E^8)AEPUS<,F(3G9&PF+
[9]^Z1<RG03GLEB&0H)YV3LMR]c_=S1&Mb9&bAYBIH>B3)IHa&731TN?UVa#_,-[
?84&=S[L9YM[,RUA]ZVT/Ib0S\1HJU>=.#eF=X)[Y/I@?[XNCc_5:,:3:0gT_YK(
,@2<e4J0O//-+cJ9\9LcZ#3e7<B,T+-X+Dg/VJ6Fc@TR/>e(:A4a)0UKBQO=3QTY
[GE_Ic=Qc0da<I+GIgKd[#..e=FCJT88O?ZBKJ.@V\M]9E(B)RfQM#55CRQ/g&Cd
P7C<,X>;-dZ7=D)b;X-;NL=3M6Ia6WG;3M6f7)S-cX6=_c.gYegJTg1BVOQAA^L7
V@VD6]W++JRLRDZP2V4cAZ:S)G\HYZH6P,)PUYE5-)P?@)#M@KA8B.e9_IP+A2c,
.CMD:N0C\Mg4\eVFH<cUHT5V+@e+b2MFd6C<KU0O6NADH^O(6OA6::L7_c5R3520
b@b\0)Jg-O.ZGc9f8_-ZQ.d#.b\:V4:H0X7Q7NHL=2U+C[V^<-]KZ>M&I(9HN((A
0B>93=X87Y[FgDgbDDB3CEVQa,Xb_c4;XU>gOBM\7]9/Z>^-g/)]cD&PYOG-B=83
Bf\S>CAd[]X?V&/G5FQ-^Y[C+:N_eH&^@VaKH7d<IL6CA/D-\cR\SDeH7((fX2[.
7\+.ZUE098GO(eIB@^^]GZ]MHCbc]OS,P+eP+ER:?0_G:gg2/#4,f(cN8/g;+eLZ
HUdH(TK[P2DQZ7>4T:M7]B<5VS0_N=<YN6a,RLV\IO8V9/3K<.AX\b@cd]NUQLbW
[O;S>)LQ,bJ1KCF3b=6QV4:KMdMXIJM0NNC1Jd^L=&2^H?CHSCC_X[[/.SV\7N_?
T4:+74N]/fGCc-He/fD]ITZ[U^(@:IH6T=:1PTQ\HSQe&:X.9P^[(Se6JF&6GB^W
R7:/GV2FIAV8e1_+A#?J9Ha,78Y:1gZ,c7+;QfZdT0WR:X3[GOJ[A3B/a8#]:9O6
>#EO=TRJ+g.d\22.dff89ML,&D7AgcTLV=RETeL,)IY]d(^;=g@6D[N&3R:d>[1f
+5[K.L-,05;e,Jf\.eLO_\?c:,/7#dD2XcN^f2[6&KN(Y#36I.BZbaKERXW[)16a
<M#>4#F^TM>NBg?M\6Sc8AZ;(SV=BQI/a^@D15TH2.NTK#CBHZdH=:JC@OK9>eDE
N[Z+/dcA/6U-M8&Kg(JW6YNLe(YEKbV0]D[71g+dU:a\.,RYQYQbWC(UB:a8RE?_
I^4O1(e,@N2_:/ZXG,?c3H9;0d#W8-\1>]O^[IK)YCS47/9G0T5G@NefC#c#fNIW
=cKY2OF=H8g6K]f+MHD51?3dW.<8X4\Z,cQA_K8Y&OL;SE9PZOUS3eJ0841GAQ^\
Zbf2XDCT_;/-Uc9M?6;08]43W6@b^Aa23<FfBf-2/))a<GOODJ/(Ie_bB?ID\^O;
Md<9;[.&dCJ_^3W9+a=gQWaF_?/O9TR[/VN@\]=ceK66HEHX/1HdV8K_[S[Y[R8K
D>f5+JgTW^06GZ_]2Z8(M27Mg(9Za&OF,=,QY8#I?cBAKR81IfKdQ2?,XF1;DIPA
\1,,6)_.1HKg5:<KWMO[I?;f:8,HS4A5UdK.Ic-JLL94Ya,gS39Y7X)>Q07H<X05
4J?&Z,CY5YO;HBgf]c-@a/26=3cTdcf+B;Q/2G8XF_,;Y^HJCaZQ.0_;_3\>ZGAO
EFXN;X=d>9^ZK[/gUH)[f[R?]E0#e+#YK8G6>eD3(,E65N:@]B13A4efb_HPP<eO
V\CROT4f&fa8W+U1YX6aK-AH41N+\/M-MS#=5b9XQMe9:AK&ZX=3QIL1PK<L^X,@
4&\JEa74MFX=;WNgA^P\R@S@BG8C;>)6UT<f(Ta8?@aZG><+:K5(B^0L#a;[AO,+
1))0(\SJ;gg5Wb^T6KQ(OTRIV>).HbSd\)J64K:K?IZfUX4b6e2V5JP5#[Ke#B6W
W5LV_aIL9_,,[N>\c+bR?dJf-N975M6YLH>63#20&a6,d7)1W4)A974L38Gbe[?6
HBFMZX5.2:),7:^EL5,17_Z8THLVY_K4(HfD<<&CYXZVD0.R9REF_a&@AfD;(bP@
HRJG+7b&Q\f>,-KQUaUCDEO\T:80E(f><Ng2=cVT9)ELD=9SeQ_BB#aYKFS--9[\
.K=ZM\YDB3SU>G8g[12794AE[a._2WCE<3fETd^N]I)H0,,1##e1fd[92DeNOW/N
AS#C-TL-3@EO7f&6(Z:5EN:6f0ZC-aX?Nf)2ZX+Y2XYW>]P;gYL_>\5>2#_-L=PC
I9LH+gZMISJ^Y#YBN#QQ3T80/<R58PT1<&J,,&SU-&F(Z5=c;_M=)<Ta6dW7US6Y
]:e+Z_U0DgS3I\<IQ_G.bWMRda]a/c6]a][8+\7A>7+^RZA4#<>eA[MN22]=eBfM
_4fBD119>O@Zd^961C+XF<)=g]K/PacU(JLN?2[0\=]e60OP=E/2A0P/=STLJI.U
Eeg-K^(_C.M)550aD8RJ<&bGMXIO(XL;d?eJ-F2W6QPJ1)cGU(\N->2J(,E;,A9+
PXaI8U8#&<?#)^\@O5d+EQA.7S<;,NQ/EZg0KI.>Z&gZ4&+2?,6HG8D+KEdUVJ#K
B-:OA>VNe;BMbDZD8dPTJ:(/T523N@.+K_EV/D8D>]gJ1,=#8XK19Mf3G,OKd^F\
aY@Eca?bE&5ZT?D[V-<CY9MAGFPKd6]bW>d_)^-e+6AEa6BY:.+605(7H#/6?GOg
NV+(b9XKI<A1>Xb7(4XQ6#D[?[1cF2Xd04B0a548MPKN+/]eb_71AC?#F86I/e[/
38aFN:E6<5N[0W^FC+(APO5:>=CDPfQSI@6#ccZRM,+Yg(9b&[>-[TA-?5U82O\C
fWI8UJ0&S2?+O5HJLQZT:Y=(;-8:f6@A2J8([O\5+ef.6-<;Q+;ebKWY]W\c2e+:
WA/;KAX80a;7VH>-D=TYA;;H5RS@1A6PO)X6&@QVWcK-]-6CJU==UPPIFS;B4ag2
49SMP/N^?-9051_0gI66ZbMB]MX3^;MUG),#VDT#,b<SBXJ+dSP50I\Ofg#U_NCW
4(+NMH7+&b4FUf?TO=Zb..?9Oa2+1=7H5PP.#DZ[D8,W.fAM^XQ((BY_N@f\eDcM
##0ZFO6VNJTKAdGRg&2HXQHX=/4GgD3I?0,(O+QR/.F(aM,X,M,3S3[9dCA9@gbQ
(,X#_C(EG7.RP_UPABZYbK(X9PC]ZH<TLgHLG6aEWA)5#1>S3+ZK/e]&S79M1dCJ
82IIacM2#V]+\>XbH+-@.8PMGdH8e_7AC,UBgSP<A^IXWM^e)C.V?UPRIg.;F_W[
3>9UFd->f#)S#,:G:J^:QK\/b2798/X]:9;M2;7[E;(PGTBWaQQ0W=U>LKOQ-H(5
DGJRb>QTRB=3C8DU3<IS+6L6IZg253EQ]dEZQ>A)6Q/22Y3PE+E9[S0C5AcR1@6&
<G\&R9(A:_JA5gL@/>aQO.KfB1@)>L4H?B0E._H\Z(9P^Yb.86ONNBH:K);A=0Y4
a)=L;BIIfM9N/?MF6M=f)1;[KFafge/=?SF3Lb5@-AeO<X\FaVOd]\[c]2G^RMbd
I8>R2<80AD4)TQ(=+:&e?_T2O8gC21A:20KgL@V-W?.7TZ=\(?\F&:bK<dSI+66@
:2aWZ=[e10IZ2d3]C?MBO\@(L8a:/7^c[a1HY-:4NS;&TH,aRAB78_[Z@Q;6UaJ,
3>HDP1?,&=4P<\Ye<:U?4d0/87ZI9C-CbAOd-+=Ca/dgb(fdHV.(d:EH4QFQNKR1
07<c0d>7;][4X5M?+7RO<db6>Xg]\@.b,?1SQ.@&I23aIC82Wg5_Y+I_Ma]?F@+[
>Y:K1<W&=;]/EI[Q=@P:81H9N_60W:0):9B,C-IRKAI[)Ya3)G#=F^e_#JA73IBS
g,aSM<1#,NM8BH<I1WFI>_c(Q<9bTRXCL]TJZBF-9HcB6PNPCK24?/,Qc0^VK[aG
1e&3UT34;+4g?J,.7[+PH.:WR_c9]Y9_Bd]1Y607^>/<,)[JK704JM37>]9c/eNb
GDaP(Jb>41:be]-\1:4cNL95LE-N2a.](M5.BO:4OG^.eDDb_C1TS7#3f4>:FS9X
OS[JaYH#>M(<B=O3YFV[a5Q2Y359abP-:/g&Y,\W0TdCD]EFA^7B,Ug\BZB?Y=Nf
UQX6,?##dSHaX]<6-B_R4.9C<^R^dbJ9JU6_IMEY3DSI+<CYA^AGJMM,?M/D]_9Y
V8Lee_H+ED&N8-d=S8Ed6Y@^CJ,U2b:WQQXG38BR@0DYXK;=E@89]VQ.bXPg1#@I
?4SBA-K)c1,=MTbcW5H:>dRX@B[#f[D/a:(QL)Q5+GN9<C]:L3&;?)7F@\0Z.P))
_aM]@[][6#;K.#fWaHAGPT+LE3:]W?,3JZ+fRb]<9S5D0#a/Ye\5S)#5cS?XP3L+
O)V+]3VZTI52:VU1R6ZT;PJG@\:9e9@,P96/C3)\RE>[f1d?#O97HFM<AP=Z.974
JI0?W;@(/aETTDfU2EFLO[/GOJO\]3(T0Q]#@g4,J1NYPM/\)0eeOQ>+J\FHO+&A
E5R:_219fHJBS=T.O?bT?G]YUAd-M@;fbYL?L?aS(5;,,>)1>F8^GaT.SX)MJL=7
8eeT=0P<5f126#STGV:B@KATA6#(W?5VG=\=d:AR_f4K(c&93KM;=-C@:E__(S(9
.>Y2\]Ib7RF-T=ec8KDQOE09-KI<KT,F:9gR@YDPQNc-WKG[T>5HagGa#g^^66gW
Wb<O.SPREfT##\>8\AU>1UD\bbR,<H9K;I.7dR1P,5S4c>1HeD4Z/8Wd6Q=.X(c?
=d@E==AQ^)FT:c0Qf1KgSDQ&(+Q:3f4__f]8?S#&SW#I6>2HYCI.UP2gH(H3CgNB
Y(bZ+1GR:TQ,NM.S;\^^DDPe(^=bL6UZ-Z_VeJ-3S#)JK<<^QcV[#)6BN0^ePO#E
9YI)6O/R_J]==_E.M4aL?.56QR_fAW&7HR)I>TI.N&U\@,C5[M5]]Ja9?F.6_##S
ES,V_I@(,[E]?Xe(ZX-LZ)TaC9#8F\]NBga#S)M[JW?X,#+\:.e.SR4gV;E_2cC<
O]A_^359NgC,L;RL>T<e3DP;7)XLC8LW?=5L7>0DMNF8&>1^M@Z&bMeIP642W1J<
R#E]GRH]8/F[@YCKL8BA;H;d>-BSX=eD@/)S>\T2-RA1IUJG+JbHAS\5(\-T&)U/
b@a@&7XD3g(ZG?<XQAaCfS1a-R\GVWRL+#-T:&=85g#8L&;L_6#O(@d_-F6O8I9+
;)GO2f9cK:O21c4BA2Z3NSS;I8^/^Q3+NHG4ILZWQ\(@=BIRgJg>bR48d8VKCfI\
fY5,gALd=KZ;aDNC+1gFfXYV&/5V6>]HM>IAA8<N__bc;0KMRZJ]?B,?/.g?/^\E
Q+?2b,_0GFDeQ(NI1]d1/HDIZ=]Q=83^]9)X/K41RV/9NH1&&edI?15TCM\3BN8A
d/eVb]TTR<F;VRTK[>+K4CMW,VS@8/5aEBUX\<.K_8)>93Bb]_L7G+bO#B&^&[\2
H&K7:GZUJ_HR@;ZZ:U2_)RE07aef377CZ1PJC8Sc5d>5f@d:-D707VR^CM:a9,WB
;_;K:18<K=T0M+XO+Z36HFa:cGAT)U.MR1F_fFHQNFGb=13N78FbfCVYWXW\f=DL
-4D(gXFSRFE-E3Z_+c[)CRR1;,]VP#Xb@&ILdVd,/.]2)J&9H^a_>Lbf(1g7\9H,
-KZ<>0#UJ[eT6c]T8g5J-OY0^IPA4/3J534fE&HZL+bC9RaRg4J/\HQ@Fa6(G3R?
\M#(?,T/=c.&\f_Y/4&]#JHAC)3gGeQNZ.-P<3SM?C;d07\QV(K8;7XXDWBS7E#b
c0R9J.Y>(1:^0)g(.+eJ80Y_:6;J,S<XU_[b<8IS5H.7&2f<HZ_RZ&@PLeAE,Q@K
_4^#;dQ8_+7UeYZ:K,LNg>M&IN,UMPZB\<FbWF@S9&4;2EYe&T^W<R@.g_[^-JS)
bgQ6.OgU[L:IR?=8:^Ecg_)R<L6P/@9f4\]-eEG0f]dMALTF)RAg>W&/aR=1aK.f
>QX9,P]@LAaa[I):NdH,Y/aAJ2NH0GW47#e8+(.4-IL0S=YPQ5S)S_-Nc[><?9eG
[5,4YG_&T3>_ca-&e1<HS&L5#dL^BT[+\5@IXLU?#[3bgQ/__gWeF<4]b?[KSfVS
Eac/0B)>KVTQUcELWDDN;aDg5Y,af-\Yf?WaF632K7YgVOP[f,<YIYOK^Se4/d(8
d,2(D&I8(V4O3:8PZA9IgJL2(LX4P4+-F>4Db>\d=,#f:fINV+g=@#ZcdK=T]QFE
S/900NCaf^?^\WE9D]S7g1[5Zg>/9e..QS-J/6(HUd(ZE^f@ITCFDEAe)ecWH+d-
ff?I),BIS^VaU1bP(94U.adQQC@KC:dBQ1]E+RWR4>>J\6Z>EY\D3556A\@0,5MA
>L&1cG8^f/dfXZ>BA=Q1/)8=U.S,2#5\>5Q>V]6L?&9>,GZZf^f&[HaQ[5/V6[8M
Q6e7T](bYX1(@65STD&6Xf+dN\T1)E#(UPbUAR?5W4e4:S;RKdQ3a&Q5aC)RJ1O;
]IH2T[O7.]6.5G[^+&dUFR_VKW3g>a2\BD9\H96AHO&S)J4@?[RTaF6c#N6SUS-d
H07&ZM_]EOY,gE+BR]B79E-RZ2<8LTJE4LgSU:Rc,fW]P8F4S],3S&6-<LSI^.^<
g#C#6fd^cVfP>3ALb,>1g0P>K_NI/NcA^U.G]_Ae4gc^KDUR8W/TI;N4.6EWd8J(
9bS-H_WDTGU1-4c];f@=9PMZ37;=+HAWN;PW5a]VON8@+6B+bIW;6ggb1I<@]60D
5?20.)GKLJ/+O6,MN&4,83QY/FK,)6>_>YagRTc(VVH)@[DQ),<94d<?D>_aA;##
C:=0)ME\TS\U,Ree2:,39^4aK#KZX:d;eUT[abM>6cM:>XF@aH8LaLPIWH,6H?Y>
W)X(dNW_B9\;90IZ+5WDW4,N^\VMWY\;EJ</&DY#bH&UAXM2QKFJa/Kf=dXgHD_U
KU<=NSILcO2YB/b=M75.8>2/b9?aQ?WX5HV02GPDA/ZC:\b@YS8_I\_.[Dg\ba.W
.+E0<-+&4+E,DL=YXPa&1HIYBMQ[TSMSC([<+MgU^@6D(Td:Y^YTR6R)Cd.c(R:e
S6b5M&NP(_,XTC#:G-d+PEGcZ]gJ4503S?A)/P#.6JP=&75Ib@.+d0Q3I3OfC_X3
b6#:K<ZgSV?98?(IO/\AD^;XI--L3<dN[)<N<25Z9fbO<<gb7;3A?=4R3;Pb=2J7
Dc7NJ=P_:BI:0;^>O:^^4PY]\3P8N[J?EDc)&fUb]2Zc7]Q6c)4Pc9a7\_=9&4]I
5,=?+KaW)2P9b\6L1Idd&6\JR3(Ld]#dQ0e-J\[=RedH8MeW:c0&f)^(R.(H\PL<
1@430a&Y8?6P^JGXa@?#@Z3OLAY9Y1H-LB</OYbSXHa2:6K/EFO[fFLGP(EAR^W>
4E/FU3(Q5G\[-KCG+C5/Y/9e6FfXdKJ:=8.I\#C=?\7^OZP2;^DK7E2&I^W@-OK0
&_@Z^SO;RQaMM6GE]7HXX-^(c5G;0MP4-<EeONZ]KBR.<Wf[;GX=V;Z)N<2MF^\f
NR0ZB8=P#4SEQ/Uc7G<>F9-14ER61aBL4@3DRB08GJ5J&&Y)[:M[?=NGA;b>^C/I
EJ21fGXU:UZBPWQ9cKGQgO^H2c3U?]N.[P3.WE/+V[=gC^KKe)G0N(&_QEXc&5W1
2O^;9#aF8K4LCPIF=2c/HFgMS?Qe=fZPZU:H@4=XA]71:8H7RbL)DDTI6b[(JSac
ML65\\2MWU@S(ab)HV(.Fc-d/Vf4[#P@7a?-b,7P;-#KFIC^<X[Q(fBF,#?UdBbY
ef2bb+4f]@])<]GEE]LA)^V,.DP36XcQ5L,L#.;#<I>/VU++Rb#?>8&H,f&d.8#c
;McFY:PLTYELRA4GXVE=0>?U[YAOb)Y><V7++3P9GUS2F5D]VK#.8352>;C_K2Jf
PMPE<RZfU0/gWN].C.T3KDTFg5_C&/1)F8875+9^]UGWd/Df+#Y/BD_D06[G@JGH
1K32D;,FQWUTE?.1/X27=U&>Q_fGaA1e.V-KddKI1-5^<[C?FM&JDZ;6L-\\TcB3
U+Xa5HE(7WW#,1T^A_0-A4);UDRaEY2_f#-10U]RL7K/DI+]U>cBMCVZNRVA?U[8
B9[Tf;OG388DMSVEEEA2db\IZIOg#N8aCTP(Z1.TYKSQF:M+V:,BaEF6,B[^L^XZ
1[AG_<E:64cF(6&YT>77BZE@9VYbKJY(Q90,GOVA6WHd7KD93I[6HP_Ig77P+)41
1OUM-R:1gR5g6OG)/2G,<_GTO>3R1HaE7-A5a(QZYg3:L&L1^+=M+=gQ>e=E?KB+
V,F45Y5EV)+Y9a>X-EdVHOTAOD&I\5-;f>b>OF:#?3cH46QgIQ:885a4eN,Q^.7I
XKEO>Ude6#BPD@?UNaFCP<L^+H);BPB(T+=8Dg/?X;cd\7\<?2V3CA[V5+_d@QXV
d(a,gfU@g.TLR9Lcd1E_1YU+VZ5DNDK6[&[V,P1WU&g0V:J>c3I+Qe;-8WIX,<>A
8<9:D=d=G\2fV4fLc^\M7;]XQf]R2I+:R7:PNU6,2Ma<7]8FX047J-cgKPHc1Ugc
3Y.B4DH<P^BS8aCZC3XCe4N.#_9HbMSEbI66U0/?5=KAH9]@bS:17?<]1/@C9bY&
RC-#\V-:8GL8@?7&_c#?UaX+\P-5PTBNWO,KV-=##CKX+5]\.c&KFT:@)@.\OLK/
XK[8Z20)cC(?V@dX4;M_/KEHGVSZ0@?C.L3_DSALH+39T[@FR(1e:eYcGc.TG#6I
5KMOEQaA\^>_.6:WMWfA/AAC@BdO6Y8TgF.a4A&I9WaM@VLYKa.#bFL49F/_bd+\
9G],;W;BAE5ZT14N:?SIHMEd-CR\:=IB/@UES<[a-GdBS-Sg0<STR\R7NGNJ2P68
Z[OF@C.ZUX/cW\?gZ+Ked1O3_e:6JD1]=SEeA.YD?CKR\1+VH#OIF,_^QHVM-JEg
5B9/N><1.XABc55[&[f3>^cQeN(2ZG0&HeHEL.PXNd[f8eEO:(.G6Y].BCQ:<U3(
Q]?b.TL;GCB(8a/gLQXQ9X?<c<O:XgaZ0V+\E;gAWU6,fXT.T&Hb;(9PO8)+0=.?
&TH=80_81^3].;CXZ.?b[OD)dJ6]T].:<TBS?Z7Z:HQ2?db.ag&O(;UMC;P&L#_,
2<(Q\>8fB61:00=L3C;=RJ83VK9QCg/45NHc>Q[E@TR\:\APOS2^>f2LCAHb0Qb@
5DKcZ)>g]D7U&be?G\ZN8H8UHJSV3bM7cefb4/=&G1XMSe/e(S=X4V#<4SK3N6Jg
HUXHVN.I9W5:]9TKE#NS8D\URdb@OR>JFIaO)C6P]G=c>B2Kc@;<fAdUKdF&9T6[
\M.MKb513Z(75?bb,2dAY&==X^b>-Y(P,JRAVa/?3@L35K]ABV)fP4GAfNRQT:MW
Od5g)<gKe:@U(^AF=@&a&UV+DU;75#,/_+1FS009)/Y8e&1+UXJ@W_?4Y0#e[]E]
/I=+=V5d@(H8a1IA2G6eQ,a4Z7NG038-CP=M4XJKBY^)37[/;.X7WG.)S=_XPK3D
EZR6Y_9gDN2>1L0C^THM3I^=-TJX2Z[d75CMd,X@54\=OfZOc+_>&\J2]VCNX-2J
JaW7.;BI9O&dLU8^KGGAZ1I9HeVN_[bAQ,,,,_1P#)_g+a6f.eZDE:gT[9&1H\PB
4;REF\@&&#Y]@]<-CgG[6X3XFXI@^K_&;D.;U@)cZ>ed]7O,<^,N3X[J#-(/aKdX
agHFaR_(.@,Ie9U]c^J6cV-eN:F7[f4eSGD/.]dDWf7+T_+JM-=V:MM,gE1\&1-/
DQ-c>_-3ZV+D-Ia2Cf:#<\4_)UHM>4G2GE1dUWTD?L\GY6/N3A1KW?AR5-SATHYB
-.=BMITTK\I0#AME/b0X5f&2DU1-Y;,0AC6@c8G-K3D4eQNH\-)21P+DG>)0@>2\
R\CMTHBJeWBG(ZT9PW17:g91KT;OT3e2&FE7g^<>AD+ZUN\=^)]@Q5)_33KZV3ae
ab&LW+4/U0fD,NNGHTK?=(M0,\65T+U2[]^18<2NQRdc2,;UU:Xc4X.WXVQI.FKT
F,ePQ<U)<4R:,-UCM--Y@[f#IGV;,58P6:TWda6Q?1;2[2Vf,;K1BU=aZM;cXS>e
U=PVPFF]\#K=87efg3?27@]48ASc^#XF=I+MY-SGeX7&aNYUE)V<1F57CEe=WNEd
>P?.O;e7JXUb1D/c\[I,UQCE+aOZ48Hg-gP\bd;;PeFX1QE1W1)0S36A/VK3W2Tc
cGPDc2N^FBK-7+>,8]dX-#7gXX02@/fE-ORPXZ;@a]d7)K2QVFPcSK2MDU,W2<)b
9WHQ8Z+cecBS,,6YCNd\V?=U-5Ca-;6NdR.^<FLUEQW78I1(N?GZ\H9gA\C-RP(9
YO#9,aL(Y0BB==.4K\:PNJW>2(c5?9Fb<1OggFUTEYFN._g/bS+S&&6@\RU#=I]2
<K^==-E5)M-7?^0SD0934G2CF2IQ]GV[7ee1U@PI\,09D>e,ZQdM?43@\+F#@d],
@HG,Q2NL89Gdd,DM<Y2>L4@@NZ.fQ2(CUX\/B,4]UK_F\CF.>2PLMP4,Cfc.5V<+
W-/EKV23C+07).268;U4RLC&JP(F5c0R4VX-L1bWA?TOCfV8[=<YF?OLI<b<I(e:
)@\]6@]:P4#W1K)Og<EIf(e@U,FaU5[S9>J6:bGW?MKFc#DIe=d_0RPI,I?d:DcA
)0;#K4QJg-PC86Y5Ha2^>c4A<?4eHO;B)IeA33SB9X(FMg0AR^e.b(LYLE.Ne#Z-
3NB]a]RPF33FTD].N)=MXAaOR7Q:7f3RMC<RI1f?@M=FC(U<[D\XU=c&5RO;#I]=
=_T[^#;32@U4f8N;3S5WI,B0#_G>NJc)+GMbM5[Wf5DX\YMAV)DG)-+3TA]I]K\8
1d-L62ef8eV4?1Q#3.LZ8J9@02MCV2LdJ<e-HK0:KQSW&)H=CFB41XES#7V>-HD<
-f2;V;8Eb;eN84#_9Q_SeU1cT#>Y7F/?d8]TU-cZ[/VT61;^KK[L[^EIe/;K&bH-
G<;+.^6VJ:91]3<fbPR([C+\<CcCA:f,AdLM88,Z.MVJD_M&E(aCb(<Sf5:&K))8
JWE>Z;1RcAY,PedQP:YU80@(HgU7NZIT)0CUH2M_c.AOWX(@D\gIU4BO5HQ0@9W6
MO<)SP]Ra4>GB6db)T2VNe>)PEEBQ-c85DL+Rc;QW:a5I0>H(#BH--DIN4PCIN>a
:H@4c3BAbe<A]I-T^\2A#)WaG8IJV53D36e5>dKT/Xc-/Y5A54bH6M>;8>L7+G;R
4cD]Ig.2?GWL=KQJQ+aHLa0OgT?A.I#SA?L??JTaF6@O\R:Q-:8KIVIQMRVGLaJ=
N:\eI4[V_JL^ea02;Nc?XP#HeFRA;HffUN-2/:FT^VL1PfSC_12d^0&JOQ5=(:fS
O^56X9D9Eb1=Z+Z5[,2_aZ@Ce7RY<?cZMSb&F#5)W@E7_398UU\DR.<FH2UcZ:);
)@UT-KR+2=?/XL+R5,IPS-f3K13JY<HaX3CcSQ\F,KC3TNa;NECf65EMS=FU.^Nc
\6eRY1IYC&\X8#<3(7@^=@3cgEcc.H^2[=B#<gW)#:GbU.Y2NbTF5BVF.,T&4D>c
+Y.\6A6[ga^BV]]fdAK)AY\>NL^^g;f7+J&U:D9W/S;+LbC2,TXG&JO4.f10gfD^
FXX#<?BfNU1+8dT)(c+&BJHIDT+1a5Nc7KaEM//F1UW/OBI3\/Vb@UQG:ab48KZB
CXG9dB#5V;H<FfH(_G+cKSU_,,&(O-9?VH?aZ,O7.9RCF590Ee/QG4S:OQGecSfG
bMH>5X2.;51R\3:MOA-/T5N,^\SRc5X>MV\&YBL.MW-c78Y4\W;\#R3<37/)Bd2@
2OF-#:>RaO)HS4)VDMO,1,gY9)4WfB0JVD]5^1AEDcU8(?TOTFYV:44?+&D#/C4^
UFPJDb]>0f87BN1Z\;=YgJ&[MWQVe(KdO71bII=@6OJ9+NXY#?L)7;)]X]S;EL>)
D5TX(HE_0)PEOAI66bD_G52Af0:VP_:G/\&HH4VK_+Q<^F@Q9FRB&ZWb#TeeQ,Tg
^M2DC7;?0(Hf/LUP(HJ1O>,gN&AX<gaA]\06O]c2F>-4[6#NJIZ4a#Y;>31KUHQZ
+/W?^L?#&[cHAeOA,E;>U><WY]We15B?TE=Y\ZB_5-WVU2WV7@-Fe)^ed:-[NH>A
:+#N5<_8f+Gg4FRTX@W[Kd;KSUWf/MT,GZ#S1b_W0KSbc\<KA(?aVKTLW\FDX[__
aE8L/-YY(@Dc;bHNP\V4PDZQQ#[A5PLRWW#9\^+04^Q&LeL\e)BH5&.fC_2SCTDe
<;3DM2IILfb2aQX)UUINLDd#4[WdQ?CMBYfedfMQ]+c0[;>Pd>R&U_I?1S3bdKd-
1QD38Y7Pf3]1Z1EGGU<9OHDM3^f[9DN[^d5;#VRb9+<d/^(O(.DR-U^8&.>/HPW?
_:0_=KD9L2IA1482U8C?)AV+e^e-bP>3_JV3XWVBVX#/R[23QWa.]X]?gfK3c_/-
J:.2#Cd::\AU:HagWVB>96C@:VDaPI&?cLH7:&GLD6X,Ka@ZX\Ka:-69<S\W=J4P
@L9H(:;L2K^#CI5^M]F;-d+]&Vg_:Tc976b]QVM))=\A45_(QcN1>KLa09F&#e]@
cZ)Y1P.9B\MfP[K_S)7_C:WZAe_Z5UY^KB]W556A]H#K3U4fe8JIXf(SU_g0e/S=
[[FIH8R@IS=N_ZL^Be4[:Mf#Zeb?7Rc1H(SRNM-b;J@_+B#4?GSELa?SB&S@DDC_
LIgBVH5/9_;8YWf3(Q&dL7Jc0P8Re/BST6R2fE^\WAHa/WQKM@=?R(MQZ-,cV7.B
E,B]+.DS:K]1WEb>T2c,\X80FD8301MKYY_ea6N,9<?<JaIKNScRb(ZOMXS=EWTb
dU[PgHd)L/CZ>5JM]15LCUZ_]PENaE@JOQdD/:I0W7B)f[ZATF&6L5V@.WY1f(?#
H6c3O8S/URAZVS5D0:BZK(TK\99+ZR1ObdW5DH5+e8c7BF=TBR,Tefa1C6+<E5+L
,?5_9:fD1;eDKGT912)g((<Ga1O^R&1:53UHGA#.IfD+6P<e5RPJIUAMbf6G//3f
UW4<&);ac7@;RdSZ,6OaCCIZ_T,MCG7D;c-;JGOgQT[4N+I,KGM_>]](g9N][I(4
_EHS#U8I+G(7.#,>M3gNI0MV##[:P=fM:<^S6VbMJ<JBFR[\fD2D28PNIOC6=GXI
89DQ#2VWN<O9)2F[?IC;);Y6:V-;(R,,(5TY=::])e(&;R7-e7=R+_>@G-eU(?V4
IN7,[bG=I7PfNCFLK6Sf5?3+fdCC5HPU>0,2Z_80RKYg<?>,RN<c-IBM0[fV)F)N
\\TI?1/^5TIQN1.HX>__WSFb>[UV9G8]3WF=^4ad6Y-,J0eY#CgFT3>7>7[V5,=6
TY([J-P]]GdO]WLZ]/@A(O.;g;YL2L>E]Zb54L,O_F(QBT_;46cb7]ZO7Od1OPT8
g]eL>L(QRK,Q95Z]f+<.]2Z/JIaR?MaD5(H=-@EUPML4#\1=FBH2,4Y#f4cW_F42
-CU+]7[G4[b)78;#3a4f5NdM6eV/O25L)H#+_E0fX@aaLcKe-5+?eHG#9aZEI(7T
E&YGX18F9;X-(ceF2S:;TM/8RCe^^T4XCU4,9ZTX+P2:.<<CMGVaE+;&:VVHgg>/
aTdDK0T?X<]4&,)5W7:P1AQKLcY?Q4103?00,W6HU>2Q=BLf&G6P/GV4#NVdg9-J
Nga><D>/E=/#d(@0;b=I#0;Z7N<M1BH8]P8>S@X6d/4HAJ?b_@0QQ+#5-4c4[<)A
YM/)45dT7)PJf#a)^=_YHT(Y-cO]1JYU^a77:LCD4AC,a1=6VF]bUC0A.d>6aD:D
&;SB]J9b&,GJ-C_C,9N5R=N9>dAb?<ZeALAa]_Y+85-;&3I-aeXD;<J4Y0cF;KTe
/N)CM\U(T+a6A,N>N^+V7K;#.J_.GM3WbMWa)X]&Y48+g=&D<-ZEKK@K<RZf6(H)
b/5Q&Qa>^43e3HN\7e>8eAHJ@D8:+3G3I+)De2^c/Q,><0(PVP.,>7dg6=Q>UPFF
1>)aGg=VF^#3g:-#>&fGO[>C=IQYb?]0S,7SCcGF;716?T,0g?=5DHBTC^KR[/T?
6=80[W_.FHDXaTF:@JU?/OOXU,4I2@[Z9<?YIbTJ3.?,;dU#QOa[L)W8XE,#Y_\Z
+#QNa[9UHbfe)LZY:>EF]a,B4J<#:JSM^#TUdI0/P[OP9(U:&F4T0L1?8S#<?YU0
Scc-GR\9Y0_d0_K(B3f+<UN,Z]Y91fDUcLCNCd/Of,V[VYaI9-FEA,D.Pc7D<Z=[
<QKFAfX]cJ#2YE:RD278G46?N;,FHd]2:498O(.K)fNVD^\OF7])0,H2@-IRWbF]
5WQ0\7,,+9/H#APU2F.X=?fJV1&\c.Yb>]@K1[7e6VD^)([BI)JgT13)<.GSR-e8
C^f&==7=5(5SV/@9F]gf38BB<SXcB9a1gW0f<&BN4Q7Ma7\18[#N.3ZDgK#SJ&CL
B;bABSV7K/F)ebR2+42SY<f1]K-K+AL23TY\b2Q/[M_#S<V#KN040;U9_QJaf[Q3
\NgEb_a9#DFe@6_TUT2fb,gK=6b@MdJ[/G)2LfGDFUc=/B:Y2^&OQ]O#VH&#,db]
[33FQ0Q&f>N1EI#VbfIC68EZc[M1.@S>#KL+4AWKcF)69[,[Y3MO[&H@>T7S\G1D
f9.8E[I[gO\Ib8-.X[JgH<FB)bCUdb\ec.Bfa?N\@)W<[)X54f=GTeTb#:KZ;)/M
HK(B+9(e69.BQZR]Y[7-ER/X99c(>ac7-@@4WM^BI1;Ogb=&Ke@@N-C3\=R44FO;
Q)[bABYI-LN+I/GW7aXZ@&C^#:SIgaP+[,_Q]GfAKGKN>VTXCX+0cC2(H4O(+[V[
DM8K.<gM6PBQ<^ZH)T2@B1^H,>L93/XY+.)YE]B5c?O0Jb\2:9H)B48D,&T3#S@=
_Q1(-^E_O&,IdLF7WAP<#/4I4JgE,CNP0@TMMW#C>XYSSL9T>\A.,c0])9O>?E]>
aP(@2,(Z:ZgOD2Mg#=</@-P0=I)]1#(f1TUg(cION3LScNQT/KFR#b7K1La76U59
0fZa,2MBbW]c-O-a6:KV467XLY)+0g2\@Z#N=&3M4PL_]A-O7c=993Xa:67^22N_
YDP^aNQ(KIcO?0,?eS5\4<K=_>C3b0fI8(g-^C+_)L9eCgD:;(e[GBW_Q2VQ(c1.
L9>-C:+<0=6=Hd544;8S;Y52EO2,:@[_d/H^fE(>=Y&/AQO9dCN3V&Z(&D?28EF+
_+24/N<HJE[2ZeKY3\2AA[7gMa\[5cC.]_/\.DP406H<)UP4e8)BI@#X[8=bLGIb
=g5DXfa;D#[SQ(V3&CBA_,X05N?c-cG3RDHC5#TZbLfbA_=059D8P[[7O2VaSUTf
240N+GVU=:R4RG-Jc@32SfN>4d[]<MI+(I[fS>:\B(9^g79b0^?f5:38dVM>U:QL
7^GMIa/\__H6/\;G(E._UGJgPL?X\#\E]/UK-AgL)R<?QPJ97ND:MCPGgY[D60)K
:Z<BX,KR/]J.JB,LNgULUWE@115];?,SXZ^/264b-^9B[V\X1B=Z./Xg4R_F=_M\
BI2QOPV].S#T<N?E=O3fW[:]O^@W#bWEW:XPU:R;20PJ2ZcMgT2/FZ?eA82A,K:6
4Jg7VO(DK=@IbH[;G2fR,P)0NPcN^e\B(9>Y>.;c[SAT)-I=;I)6d\OC6=@<_O?[
.2O#<Vg&KE^7..fgX-?/5F+3M/NXU8L=-[69IH/CAC0;JVM034&]@.A#?_<Y]+CC
)VVV)TeR/OSK1-X):0/D@?:Ucb@6NC0WcB:XU#.&N,-]S>JB/eM<g]CV\K2.@Z&.
(P.#KAUJQg:.cQ?U7g^2O)[Sb=VTIeFXC9O>DTT8W#\_V?7LP:L]E]U>E9[g?LQ_
99L6M1U[.A3Nd4+[Y:0M_+[U+a2XD@:S<X@F[+8Vf-05#E5K;.gd</]D4;SNP98A
@5WEMV#3g@BgagcH99Xd#G6&Z2P/a/AAF/UXON\/,e:TTL0Bf?TV1OZ9c5WGZTBd
R4.=Of<9-CdQFALU+GdaH#.K7>.7AIA(Y-M.Ra\,SWR)6JLI4.@)FV6++KS]Ub8>
4(UK#EL4gQ9Igc5#,1gSE0bb<f=GAH[>b8;-X9Z_.Na@ZOa,^B)a8g,ca8X>/IC8
17=M_c2,RCe.27E.,D=1>Q1Y7e3:/JNA]K](5A;gBB8L&[UT[>SU-VZTINJ(HgPR
O,W=fbP3O;SQ-JcT5J82gANdL)I?O9B0gHO7+V@[U@L3&XWUXHVD5[XJ)0bO2&QR
??X;5T<N-e+6=))cNH8Ya/bF2,2:R3O+NIA[L2S9NTA(,aVT.f]Z=Y(7<CZdF+@(
)aEc#VTO39&dOY)C;>;X=.QM,O]NbB<3E>J/[e)@8e6dY(11-I<:EY:d^<Aa>&e[
&b86Q#.@A(&g[C3+#eDT90KW+/a.bH?SMQD:F4[F=7D/?SL<B>AIV:X@;fZ0^9\H
1/KT@^ML+576-b:c9f-P/(>/=BV8@Q7VO?_3FZ\D=_IXZ9^R,9VS6.X@L$
`endprotected



`endif
