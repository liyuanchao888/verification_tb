
`ifndef GUARD_SVT_AMBA_GP_UTILS_SV
`define GUARD_SVT_AMBA_GP_UTILS_SV

 // =============================================================================
/**
 * Utility class with a collection of routines to assist with Generic Protocol
 * transaction conversions.
 */
class svt_axi_gp_utils;

  `SVT_XVM(report_object) reporter;

  svt_axi_port_configuration cfg;

  extern function new (`SVT_XVM(report_object) reporter, svt_axi_port_configuration cfg);

  extern function void expand_gp_streams(bit response_data_valid,
                                         uvm_tlm_generic_payload gp_req,
                                         output uvm_tlm_generic_payload gp_streams[$]);

  extern function void gp_to_axi_master_xacts(bit response_data_valid,
                                              uvm_tlm_generic_payload causal_gp_item,
                                              int sub_tlm_xact_counter,
                                              uvm_tlm_generic_payload tlm_gp_item,
                                              svt_amba_pv_extension pv_ext,
                                              ref bit[`SVT_AXI_MAX_ID_WIDTH-1:0] gp_xact_id,
                                              output `SVT_AXI_MASTER_TRANSACTION_TYPE master_xacts[$]);
endclass

`protected
?5)OH2HVB/eXRHK]Y<U1O+E8;RJ<6Z3)Qf)g\>E?UVYc&e,AN\Gg/)N,C3aYK<e5
X:.MZA1]@ID7T/BCOd,ZES0P8a[]..gYb_X2&_fVd0W0QI4V:::#G&02C,SI(S2B
7^QOf=FB,WW9ZQ?0=a]&fFce[JLacIT_<C5)@J-Cc,@9HTD>H\b-bL?3[(ET#3bM
+cJSUfV]<N:K:cG48_9(MAAO2^V+DNTJ@_=gOOAdJG+RF\0]]W6C3fUA6B5.Z[OY
+9S/6;8W=-f]g_d#N&I2U3^Ce>eaCIKS=$
`endprotected


//--------------------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
/,GB0)M9ZR/d,_TB[5BDW]GWV]-]<?DCSCO;25b8^AEI>H)2KWP66(,68@:O6]..
\1#2WO2<V^F2OBS2M\1@=ZINf.8[_-5W[eJ0]g1McE_PX:Qe,:bDfS.S+0^0.4>K
DJZdEMKC/Z#31<AAU.C&H;:PXH.eGCXMW9,QR(ab8UdISC/WGbCM(-Y<Q-Qb7dJe
]e&Z+Y9IUBY+5G)L:_6cKb<0QV.D+8UfWUd63-1;/a?-0>M7Of@@RX]7PDN5Z8>f
2&-6P=44PMJ<@.#eGK_1U7I[gV^LUf,-dE^Q:9+<6:J7)>\JW]X25WUI-dMVf<6E
:XM_Y=1BT46e?WYDP:TDQ@g[cb9MU;IKKH#UWE)ZUJU\M6b)R@\[-RCTXN8()6C2
a)-d-Z?d8B=J/fRA]CT9F1^cIP;0^49ea;4XJB>@Le,ARPLYb:f]5FgVe6bA3@W3
<5Nf(&+D+8,>J-;RV2<F+YC_.T4.SA1LTDTfdZ.4ZXJE^NFI6=7RKGg=#9.:?.?I
GLK\K7]gN[Ga)g7>0_H#:<5OSX<bBTb1LTDBFZHT@@2ZM[eP9D?RLLD0LZ4YR;aI
N;D^8D\Ge8:^f)L+[X^INLPQ@X)KKCL;(+Cf#fJLIAAC@>dVCX29I,;Z70OVfcFF
Od6DDU3BD4KP_7NJ6/,0+6[SQR.P,d=WGd\@b+J9GA3.c\\FP269+]C63MfUdcP<
^^DS<X7aN3Of?=;38]_W3HYg9;AN^CIEU<=I\=1Wb3LU-OZ>ZYd\FNP=\8C=[2V)
<=KBf0:[f;/QdMI/V^T;a]Z.FV]2PHNI7XF,HC&DQCZSENYB[17e,;<Y67Nb&G_9
LBa]f;@<GBHd;JO]4JGM(ZZ:USI&,^=^]H/d0cb^[EO#34R<Y[\@CHB1SG)I\ZHL
3],TM^PA^B6OY^RYM(2V/7G;<0<&KYZM&[+[_Z>JZW@97-g?>\S3:T193);BT_eB
RUV]LI[N:=0Z(#BHOd6JVM9A]YG,5F5Gf:cK8>YX+L<1-(@R#0c,5-HP4TG&63=.
:>3X/,.FSAC>L1_03CGOVBdR?2\206edVeC\;^_+5J0[Hb@M4C2D9XG=d_TcSFU@
Acb.HE3U#=>9@Bc/^@WQbAI7_YXZW@&T>CE@cfG(dYPC?E=88cSKVTW6CHR=@[9.
-@,Z)CPX(&BIFT8TW@.eW#M>IVNA4TJ/LHW<Db1\/G8&@D_Z^Z@9DSPVE7fR^PVd
]0VXV)G:3/cYAN[M:\Q\]&S?Oa14D>]HKZH[,M>#83:^.7cQ7/16^f4E9Q5DX4PI
4@59_?Y8=8FGag<F+][eM5ZE1LKF6ebf0SU.c06&<Y2eBFd,2.Tb]5Z0J8YVJ=QK
9AgIgP=N63?FH/LS3<EaYg3)2LA?6_J.Og0L[aC.D_64Nb9FQ,gb,))=eIQfD1LC
7LPA+dY7_6R=.&K6/G\@XW0HeCgPW9#-<IA^TG^&0.=KSH?Y@9C;@]4JRZV+(>X#
R=-J4EQG+KOG/aFE=2ZMY.B>>1>=Q3WQFJ7CO<K\C<:^C41g5L7<;bJ2(FEM6:=K
USBJ#GF\VSMHLY_fZB?MB8=9=F0OKM_R]g8BC9?,Vd9_C_>HZ=VM/<2>Ue]+]<bB
5=HfT.N>>[H=0L(<U.b82d@I7;9?4)6C)>BgZ5HL7-)d0,[C6JL&0b9@.L,2^^6#
&?6&H6MV16^H=)X?OW<dA11]MP=OLU4XU[0BTNTf=W;JB+GOT.eb#V),4Y)<RBBS
eX>A71]PASR&)89=gNM);PU.cD9>MTK,10NM-/K2Y@?5cSZ]K,VC;^7?aL0ZPaaG
2Z][dc-eBV&DZ#\I11.@3_3@1ZdKN]YX9I8YK&GW4@(G/PO+J@Z2.&fg<bHNU-a:
]OHNO/4Wg(.>_/,_QH5C>Q.P@PILKg-Lee(0.W)>-fR6b@@DORCK2&S@(49cK#1c
;KN15X&GPDTS2>_&;A7/Web?Mde9<]YfRP=4CJV;.+_N<M?JKN(4F-g+0,b@CTef
ID5P02<;__5_-C-P:b=IS5]?5CL#TE,5.aBP)g#28D;IP?\S<af=CZ[J#][WM<af
Rd.M@AH=N2f@R1YW4WbL_33/_NJf-DD4dFI6.B-(>/;MP?(1_]]Z?_D>.&]7Tf07
POXQLbL89RZ@TW28K1IDNOPeN,D6IG.[8cCQ2:<-,3MG^Z0a##8&JJVf(f4e?(N3
+b#eGP@[Ac4OFUA2FeD@e5>YS>fY?<R6Vd;7[F,D^#VPH=A7X0Cc__TCLf93.ILb
e1Z^dEV:\ZMM2P[_fV1O[gV;08>FLFOL=?0C5Sc,K+M&F6F59LOQH>8AFP0:c1Mc
d:>KVVcCHXGEZYCdc]GE7a^J<EF:-GZOUYgX<ZReV)QB1YUL[QW2?2Ug[FEPaQeD
;WD1J<-V_(FaSXKNKR;JDDgTIE@6Q)&C]b@E1J(Kae[+f<AV])LU>2147#=)]Ha/
20;W^4eEL^XWTH^7B0G_+Y[[3_PZZ3=4:&7)7U8BO(4SXK8ZM.?E=E8,N=Z:Vc<N
9HEFa(8N1>#-d/D4W_/Yg(1@f/,PCI7;K6bP\W+6/M@Z]_,aMECG>ad9MI-P?V@9
d/L;?CNWB0#BbA#/_^U[NJ&F5>#]D0TCfbC_R4S737SOLQ,b35f=1PbRA5[IJHP,
(Z/(?72b3g#M(R#G\FaHBecN>MRFIQE)FMK<XcLQ]FD:&A#0J>2/1.MX_?=gPMOB
+FQRQ<+XHN3]2CHETJL2BcD5V/=c#L>bNYXHH.d;=HY@@U<9CFIV@@b4J:-#/Dg:
4O(YA.O7M7,;<1-L2^M@=e+XZCJ7J^ICXe;V[D[fAP/#7.[[[7H8[4J3ZXHA8G0a
67?2&(WT[&G343A+9QMQ1X#+#S2_=<J[\[<bOb#,T9]WI2-C.68BF47LMc:1(P4f
(:BIOf6.SXPQc1<?7OeS)cf5\f_<YZaZ^\-bcT<1.M_DVOefJ3?c6JAU&-J,?CYT
=4EIN5DWa@S.+4@ZfWaACRJ,E[S+UQJJW/>-db>7\&-/;BNHG&b;C4V,3E[MME+f
?+]Of:VMW>BAMAQ-UDJBYT]?^E34S9;I93ba:.#-c?8@9E\,/5QLf\/L;^(O[9YB
/=[:=ZLH\,X_[F>V5GU63#U8CRB&=7P1W1(F+T(5D+^)[d5S6ed+0d,^;M7d:[d+
@f@K_f>ZF&?9\FOg_AVKZ4S)AS4\FP:3Haf_da3M\eUNU?08b)Z^>KIPW[U(.KIE
G9O_;2@S<Q6WQJ1GQ+YeCBS/0e8K\:L\)[UU-M7TQb-@6=e(E?aJ9a.<Q<X5E?V.
??c=.W>D3EV@fe7gb(PV7917]-S+4=\86+JcMOgV;/@=?B]M9e>?I+P4=PBd<X5J
PIa?MB2ZSBC-/YaA/U9?-Y=e;dG-PeAM;TG)&Y8K7abFDD#N&d[eW&aW<<Pee>^O
fg\/\CD][d3Q0B5;\F_,d&CCLR61#PIJDLS7?;:[@[ZR:CI]^TSZ:.3JA6D^UD3-
E]A3ENS]]d,ZB_KS8KM2@=KcS[FB&S,,^NT>V&I,+)L5HNL2W[4:GFK:0P?HF?X.
aEBS9LIB.T4R=]7E.+_^-:IP+-Y_cYNb)<CS#U_USE[/O\OVH1[A[&(@^W^FT+#@
/GJN^f?cPPg#FIKdbZ@C2ag=DK:RWRceO/?b]0?E;7;((ebF;C=R-BR&C,BdZ^#<
,=UWdP?J;N-;=><#eb56/Xf];IF&]DSG9N2(9CG:dWf)K+,EKD-(FE-FRR&Y./+g
-HZR>@<beU4(&,8\[ZbfSWGf4<)9/(1/#b1]XUK@G[P0Oa_Y?X3Me6J.3+&\Z]-]
.XKH]#XGJ,Bc]H6?b;f4gH6IP2G:@:A0F.AQ.N:__#)Q?cZa<#=-eB#9(XN=H/LN
L;Q;fbGbX)8@.-IGTANB@<R;a<a#XCC;9g;HENC(-QM=?Z=D&6.](TM;C=SCH\a(
1f_JY5/FFRH>I\9AVR5BFD5+_+Y900+)X@DOA;Z5?I\_e&7;RVC5f4_REb_19K\9
R-Q;X&MHX-MW?R93J:I+=7B.<1c-KW6d^=&:-Y<aN[[b)7I[#FLCIP9./?N_c6G9
>-6EZAZ6DVGX3f?8BP_#+?OQP0AFGTa)ZCdBW=X:AHScQec^.JGQVFb5YN4W-#R_
W8C(FC&(&YVf:ZCG\?KDBLFO\<D9RbVHJ?bCKY7=0e]3+-A_?6cHIWfHW28IggS9
P]F,1PFfbJ[[8.8]g4?(TB,7;T/\\_N(+Z+:dV>J@aUM8#O&:QL\V4F9.^(>C>e;
Q0,4VH((FGTG-H?[LA9N?8BR6aWZ.JV<_bSX#8[>;6.b3a95TcXOS=XG3VF:BX(;
dg3G8?O&]Z6a;(NJA^^SS;YecIZ5X.,1&@(A]9V[fY]CV9RbR>e5+e6BUEac(;cC
8+1GZG9U4_5KOSU1EYD6+II7;,e=&/aEP;BGgO(C,&Xf/2:\(\D4:X3&-O0>H\7N
BIH9e51AWP6:8KJ<4]3<Wd=C-__6ObLNH5Y(@1-Qc&TSf:(#4VFIKL2:G@KO_ZDC
M02[8.dE:_LK8IGG15_\e?E0273RLOS=DJXQPYOBRd9GAKcT]d-SU#P,B\K044a6
M;Tba^[NRFR3;GJDKHZ+6002G>@2:.YacE6NVD(/I5VYVfbU>GJ8FS8>Wg<?(,cK
=fB)WG3;:?/Z6D^KD-Ye5Y/OGD:9J:CFSESY4O8&b]&UG\?YRZ+g[3+&YZAP]](-
9(^:3ST>2=<=M4(5aSL4acI9CAV>@647P+MUAA<K8<-Q]KX1^NJc7B?Q<J2:#@@,
a?HJBeQZCQ3-1RL-D^L,PHgC.c7Mc674V5Y,S,SVe5HXVS<(Q4f12[]CTAA34A00
-9?7I,805R&E#N/#=CGCMd=)&I[aJ/8)LIQQc/dX8+c;+O<6]BTB<-VM?#;XbaA1
U[D3ZV\0AEHRI.#-L#T4/>>6a^E&64a_@57PL1<.E+T8c=,SZM?NFWC5\<QE0G4>
(JaVR=9KBSTU@\VZXaC>dJVMG,_aT2<21Y3bVM24SVY@c8B3]YeO6FHIDUUg\J3B
JY&:Q7MTEQOI@5RA[QdNT1RY>[F.+bFDNRPTL;5.5-/J<gRU+LS#ZY>-YgB7KTId
@fI,P/=(aSKE-:JVF8e)f1IT>@4M08;Z7+D3F+,R?BYLefGVNGZa/Y;Ofab3,#\Y
B2T78W/OMe[ZFC?&HW??J.LS#+D:d<E=OO(QOO_^VC)F[Re)G._@@(XX^\.X&V)9
GQE:A)=CGWNd0#EY75:TU],_VNG-XdB\&HHZEa8<C_3Q(N;dK1\;b-3^.Gc/]MG#
TXe/8O0KOB=M=:L7C:#V#&>\M_76A)UKE[dcU>I,W-.A_CAc/-D+A6:QTKFRcdMX
]M>Y60(P#Q]W/2ZIQ0M^/.Cg61UH013,Sa)[6[RB15af/1IE_>6^UW_&WeT<GU]c
=6e(9QLB7C(TS2FbaVKL,B=a07OS[f>0F2G><NWR@EIYM2ALE20_;[?#CbF5M1c5
;V?2EH/&KJ,)f_gNc9D:c[TC#A,#dW2?AUT#L2-V#U[C=5feI^Xc<2aMLT(=4I#6
#^fJd6B.CD[.>@UCeOB\_K64C5eK:03RPT#@Bg&/XgUS4FPQA&M4aH.2C_8?N?5?
V?V&;BB6KM;AN1TVC8E,?DSTE=MQ6D^:&43_M:PEFM\:/0H/1FAQ3K14(:S>MPEU
L_-4V(ON<#?aZ?_Ag>EUaLLcI\P]Z7[H/:c2L1:B(\-6CDP^]1F82[bH.;Te/TXF
LB,@f,\<YY,IA)DN,9&fN>6^M##YO;W>+&)6eTf+J-8=M;[^;4]:(IMJ3c-/:J^M
b5(?8P0,PFC=/OI>K<BS:@S1ecd>F\FKNEG_QQH@HO:0Q<[dV+]928JO;Ub-MER/
5[/2&93V@0[JH)H1(]7AD/eDY6U,GFDY#3(.?-Z4=AF9L7#)5A-)]^(N:?)S)(YV
9LA]K((+e3MH015Sc<2T@+,bX>?4WaXG5>a29EN;IBQWZ)JRfH6)PPTD[?DO_HZ@
7[Q)6?@C1N5@Q4_,<bC2F-R2DYUWBDgeU1<[^C?>@NaP.REKb@3H9JB<A1EJ#&5C
U/\f1JRK;#2:g&9GD2ULTOb<[7_SDdcEY0\e[]H506W5.FI5S4+JJM&7^L:\=9->
-5BU7N&g/Y3D#aT5H<]c[;22)GcfD\^a4fX48\f)E+9Fa8-T:,GdA8fMfaR<d)&b
We?=f#b?ac)9LZT/_Y#:U0DRTgd/c<0;H+3/a=/W;E]1Zg.<2cPS&ADQ5S0RGbfS
5ZGM^^>5EJd=&KaB_XQ=XPNBO-/0,)73;gBgWI#J:JQ^L(?F_a+B&EA;L78?e+E5
\-aaN_X=[_/+ZCe0K:][/1Z-[&e7fTN-(S[GKd?JD8\9_\A#ZI6L6:4[Yc?H9#WD
Jc/AVJ@JD[30gLg8-VHBIdY4.CLBY9@+SU=K?9YX91N/XE2FA3P=7f(3+I(<fRLO
&HdGS@=cJ23G)V@fe=7_^W_g<VZQJN1EO\\C(/?:[[2,Ve>9GTP6,47?/aFD[QIb
TEI+V3;3Bd2GP)6>97T_V:?(#6CV5@@K61KFSa7?=b@[eG@W1S0[NLf=#fC=:X4C
Hg.<?VLX3c-HQS(65VdO6G=?FD@)R;XA7dI[_)e:95Da:#^/IIFND[O;>;Yf[124
?Z5Lf]/J7c^5=UL>P)LCPLcEL_7BB<C:ZE]B@/Y<b55B^&CUD;X,3(IbNF3DV?3-
)5X3]6b64W5+T2\HeOUVHCZNB1=#S2ge?,X=.)=4;/LON^eSN[/B3NSJC^M6393Z
eGQ]H2_IOO@M#M]eGGK8=?47^+g@ZZSR9K8M1aOgQaY(A9.b0EAY9PgTXIWGVIf4
:J?Vg)[];I?c_&f=YYL<fZ(>BPW7U6O>FfWD8\4V,S0bH6C1B@9a&bNISa&e13_c
H,(^=8?UY&03+&P)S7+(INeYE?@MO0c+L9\FGUP?:JO&P7]I;d@>Se-+@Mc[:E7^
DVL/a#3J9(c5_(#?0UQ;0P4Q1.N^gIf1ERAE?IgR8SNP^MM<9Uc.E_O&-\fG3X44
^8)U5@dP>dc?Ma)SH6C(9VWMO(/&P0P^5\9CQ+E#RQJVgH+>Z(b4QV/C3>_E,90&
+^TMYM<^gQ6J.2d^\/X+<F;=<ZR<2@ZeF0FObSA[W==+agX+@fTb4EOVUACeV\YO
J98V6GC17F;c5K[=FA;A:MKSUGHUS0F+CL)OG(.J#(J=aDGO3:22@4KA(\-69FVI
6:88-N^(C;aQ6bO)Oc?\dTG&#F;D6aW7Y_C]16cFG\5fI(F7JJ/Uf)=VEF.XA]KT
->DBU_]X3N9Z>(0d[+?FTMBDU;P9DYcb9eK;-c:0L88FAXL1,D:dd0e\[K_W,63M
K>NCVG64I^S6K\F7b45K,BfcKI,JFBN7<](2ZX>J\09<>3L&9e7N/_]?KaC0T47.
H&(cSbeQc8^B^)(E6,W^fQ+KT@)??c[(J<BV+Xc)HXK^e]c4KPDAI6X0R5O&a)/@
H@-M\MBE16\g/U#M,6JJDJB\gfW\#3UAT+1^3IRF&ZcVd/BSH\\Ged,;0BU:(f)I
:EX:L[>G=a7T5aC_Vd1]XOaR4e4]Q]USQNGO3f&K4]&K5_7LTU4IFIX_7WG;0aA.
ffe_5HG\2a:WX^\FRgHS=QC?7AO=+-gC/A+\38FV#?6AQ(gAM7>8X77>2;d(E:7R
IZ>\<Z@BTI)).D5N+EbN<7^OFXU.;R)1Y]c#/@=@@)&(O=OO2-14\cXGf_8PS[6f
c\.?PSP1[UBC@NT9aASS&N68@5[Z;,<T5:3-P5?c]<aB(H_:/2LFB<)-ZDI(E_O7
XV&<NMXQSZ802BL6\:)L&7STEFDOAa9]I,()SHQ@<EH-c[[^gE<5X:B_W;DR^/_F
>R4a,2F,OU(1NN+Fbag&f-G3)8.^&VO(<X/&g.&P6<\D.8#ef\d)0Z73SYOX&b?V
_Pa4H.)<eb7@3\()\9d0N3@8eg1+]cC2W[U&=Q+7e:I-E[EV4QT9fgC9X5KKb:@&
ZFdeT(MHRD>dM9DS+F/2+a1S8MW(e6?T-=/5>80-bTT,<W_Z5?3/V,a)V6U6KZ+F
O9SXX4dD>W=+eS/?2ZR#Q/g93BU8-<M:W-X),9d&dab06D@\HEK2(_?L:^2;WCbJ
..g[]2EU9\1XJA/&##Ue7@&H48?BgS.]1FXI?1G-&[N7&8L2O^U4L@L7NOW/=Q-;
d\FPa>eTL0L>)#@76J;22].Y,3BWY7W)GS(W@K.CP.<H9eA,MP>A)I<Nd:P9IX:I
\Z#]N>51/48?Z_9-(FY0N:1MGQagH-Ua_IKKS.>MA^gc[:4WJg38GK=?\Y+4Yd1=
ZVF=GZRO4.J?R58FFCbbTNZ-WYEWeEKVK].,c\gdN;A#\^LO=+NV-:_aHc,SZ/O@
XNB](?,,)VZ@+a+(=B6Y/I&<0B?:]3C;(WB(\(;FCT8N8T)g[^47-a4MOQ[L3J6C
95578,;5A#fW&HcJaHC,+bI,31R:c9-SGG0MZI1EWY3B]MdCDZaI<_PPNRZAE)Za
KXEZ:G/))E2-Y?V^+/0?GPYQb3?H9?E1-ES4EWHP(c9RUaQ_#J/_/#11AW).NV@S
La+;T:-V8W>^=A7>4-^W#ZG-E&R3&ACUA+XPOR/Y74,.B+1\C8aM#9MZRK,S/43V
HY:[fSWZ1Z=N[=PNK0?/Q9g0F,B?I9G=;gdffVY<gXA9ZQdLVeMPQFDR81J\7WKM
gb@C4eV6b-OJbSb3HUW@JKF=\<QP#aXSGcgC0+1^+,Ga;RN0Uc3=WI&/P0YLMQRJ
J>eC2aC_02IKH.Y94L<7+&Y4RYZ7C5^.H.gcQ=J#R<a>bSBW=1/6XOIN<OETS:E;
()JEHNOMeg)A_B&D,IbQQeZ62RJ2(cgE1f7a6Oc+K1W[PR/9[/Z4B0UZSF;G^g@S
V?)MR[=[10WaPN+&-a;X=gecV]?QWJGIdJCGLRU69]aM8^Dc#,6(:ZE#R7D3<:BA
dSccB1[YT91XM8dCF5LDZ?.Ce+N9G\:>EP4.#.;2<WE)V@003@),^EL+^&A;eMTT
@CZQeKL,XWMQ5^d#T=Y&G<@?Y#VI]FS8Z7d2TP:_>Q;9cKM\LX#aaHf4H07U0BZP
/<@[8H?U3gf>a_EBFZecd0ZbDbEGIIUJ8>aCc#bd,J@+9M:RBBBRbfe:9a^\^1-A
A.&72K6NQU5FfJ?JTBO6/J:(B)O),1<0g7TS[A1.)>A3J0Fb8&4VTW7FS:G7(BT@
P<T)C97,?X4?8NbW(0OgILN+R\RD;<831V.C8gd0T_8a/d+QeB#CfBS.4geNBU/f
LO>#K=3F0T=],G;R.(dXB<XD.gX@^<PRS+QJHZ)_4(gX&)=U:6#a>fIA8/E>GU1U
:[-Vb(FF<];e@.W[+BELLSA&[P@7LO@[@Qb[\f#R^D]S,._8b1)&c4_0H-0GaI0^
_RG<J8J&H[+K>W#Bg-L0@3K;S5HTbg3_,^GUE=\H[WSLJZ+@R6X50Ca2W_JJQAXL
@&F_A2/:BLJ@S4UY),cEMM6^b(<3NT4JgO@-;>2f(_)aD<\?->6ZRMH6G21Q\./1
Q),ObF&,TP]XY.RH3&SX;Z2;<C(b(37cXg2g+-1#S7@R_BV?[]?I[dDPF#g>&:L;
gG)F?MIBXPVEPS1766]3B@=#WVTK3bN5,f;.Z..>8HY9A6^?YUVJQ[A<e7gUJN.B
?IR/XM8V-^@Fa,/K9,d-Wg,/3-@]-f-a,g4B(>DeF>,1STT;@(cY<@N;[.>]c75V
,9NPCdbXEW)R7Z]_YAI_bDK[d4M?_)K>K,LDWM7Y:AXICf0113RC7cDYBVg57NAA
3WbN1T/FbD.#QD/8,cJ_cWN^Cd:B7TJEQ:1P6.C.8#,ISAL=Z47-<Db@KX0/0H/f
2=c,A^&XQAO&DcGPHgdVg&479b<f^RKZ_K=I^G6?[-6XE,>3]U]T7FT^)dL)bD20
<HYOR0Ge[+5HN_V7aV#ITA(>Zg?K(5bK;?Q58TN1;P,<_c:g</[S^:>:XHWgYZ=_
@fa\CDd<H2TQb.2HZA.@P.,DI)C1Y[R,=\=_gH9-@(#:C^1/+R6#/__;OHSQY7b<
=36/gZa8/WR/Lf^/KN=UGTW8WBC[@3/\/8_Fe[GZ3e\QP.2dLb:GRRVaG&\1SQC.
^C+4a1-VM^]W\5(;)>9EXR;/A8OJ>eZ)]_G9F_O2VL@@Y;?;Yb<Rf\g8[2K(Ka/c
LP:cg.fX&(33AD,O>9^WXKO->K\Z^eJNZ)O?7>Y3M(W#4Q4(aB90?I+NU-TI4,9g
/gc@7&d^:S;)f__-Mf-E9(2#U^>)AP5(HfJH50/.eSZ+6g.14P35:)6e^BK^7<^#
[dRa\B\bEUD6177^P-C_MZ<>-\2R9DD\D2N[-dY/)X+T._KBIHd&ET5F@+d:<d9#
++R<2+]FA?:f^&a;5>bZ,-0We)V-gad_VEW?KL9d<4M[Q6=/5M(g]d/9[_WOFRW0
T5dU&e3@V\_fcfdV,./(T3C_SJYR)\8_cTS&19bKHSA),923<4Xe<NOIgF-TGQ\#
/J8-&DS<gg;2RBHgTRM<XB(BJGef+^/gOUG@=<2(07f?(C]bYS[5dIeI+EPU)Pdd
778W]LVX475E_#TAP?P>.3-P#]R4C1:[JC/EV-#7G^MQ4X]g#I\)g:(\\R4FWed&
_O:448O?JX8P)J?LXM)+=UC0D3_.WHNf&?MN;Ac5C\09_G;Ad<UHfZOW6Q<T2cKL
H;)@@].HL/#05EFESa4&5dc]&BaC[1:/@26G],_R2_S=+&Z)QMX-#Y.Aa8X6>6O7
OcHK>]I)TEZIK8_Ga]XF+d>+Id1a_WO=RY;=-f^27X)4Ng:F>Wg>1#NHG+-<>ZXV
5YgT4UeQ^AT(:&G(ZVIMIAa60.V&,1]e&1c@?8dOeDaJ7I7TQc.2gDG\2\Q??1D\
WESQ@f#XYGEAcZBE0Cd.<Z<e7>(ad<NJ?1N,bHU=f;Z2050VMaPfT[?g1TI:V_?,
#cR@LbT2_JO2d^Z^/d0E^ID]UeIJKK5bd/C-24c,4bE9N@AK9:2GgV<UT-ZaS>]B
CLXF[e8TC5Z,L#+NeA^dgR<GNIE0>?^Rg,Re<f=F7HO[)#]V2Q9U1<AP#gQAN6V3
US9b.0-23SVbM7Q#eD+,A0PVR96H:/LNI6BE^GN,(2L]eUB:KfL)(4@?VH@K.?dc
Q<WbSANY(gA2ED#..[QP:BOTeR:?X5MPC&GR_E))#PU1ZKII]RUbT-/YB_6,c0dG
#c_Z+NWK?SP.bcc-FbS3O>JMA7[VK[Se7cd^W+-(2T=\\4NE5-LA]FTCJ\\)AWS3
IW1Y)242/U:#]OPO041()2XIc^adRRZ&U,6IY?><g58KW(\Qc:63NWW>-)A4.G?M
\9(JA#@DPXI<<,\Af7W4,49U,V=5ZR+?7fcd(-gLL9#YF-aJ9L6-(IF14Nd6Z[=T
[fK#\5&Wc0Y<[],1:a[X&XK7P8M.CcM<[Z1&VFC7b;WU<_f#3[G##A#<bOY-_?G(
eW@_G4f;KF0FK,5c:_.Jf@<8<JN0gE93-[VIJ13A>a4;ZTWYg02]KC?64BNfEZ6d
e^M)F&f\d=N9=Rf9c)H8R7JLW\(,5BJ:(D;K\OgRKK>:J#bS.UL,R._NBGAWR0VQ
fK18c-K(6G+ET7KfN&:)[OSYW.0TeRg=fK&)BL8a5-J:<D?YdPYLKK@>^),9AFaU
BVO_S0VVe,2&7.fJW^WF:c9Kd3/fI4XeQFR,2IeHT5?bYNAfIR8aR0f)(D@KI2-#
UZN)EF&O60-5JgQ6BF_[&@F(G3Xe=HS71F[5^?]Lb_Ef6]J91&SbTAX51WJN9:<W
VT:WX1@T\-IS;[=;HN-HYA;>9TFg9^I:3&GMU]U4Gg[#R,<LY4M>ABH6-5?WN_A&
Z.&T3&##JgB(5Q3U0[<KHaV_3-:f45Xb]E2:M=.dTM6e.^6=RDcFH&(YSe7;ZEC?
[1cMEMKXeXeN-2[Vbd+?8a.8B]UI;:6?_VHdW8SC&gU\g0U3M=Y;g0ZFgK1&9,Rc
bV/RT3?_LXVQ]<VDc]LXDE.ZJCc\K2,a0I._5D9=)?T/6R#N&#:OgAR)0C^a.AX0
d@\I)LMT[dR2D]5d03Z:X7ONdG^-IY?,)EYJ5RYLU4060)G,33&>OWS]3>CS5aSU
)g&JggQW>Z^XWYf6U#NgW:CI[R;><JM1U-TH/);>b#F5^=+42AE6NGSU;QSeV27A
.>@#S4eO7gG[Hd.UND/[4I\18KEC1V#aXFJVF98bTgK,MQ_<Og33_f_GCea?]#U-
]HMLO7Oc,.1fX2ME7J>,\1d8QV10]dT[TD0&#Ng2IPU&g4f-.J6XKRY\YFb8_Q(7
:XEKUH]0,VUW\@_R&X25)\U>JR.[)dGXQe4FUdA4e1<<=&[SHR+EN=,+b:T^(V6-
[\B8gDDK:;PWcT6\]./7O,GG\0\3]@=41Y8NI)I-NT78INQ5BKJ9)P+9[TJ8L-E/
YAR2)aDO<Hgd;]-YbHV<#8H0AFX^MM3ZZgK8fafSC=bUM+>gD)fAEE0YB,Ib@FJ_
bZ2O?AATGU)^_6EfZ4K2>@d&XMI<FC>WI)^P(\>)WBD2VTFV5E=7M-NHRB^@efK,
F)-1Bc3\bY[Y&J(PY>/=]8??Xc&#?H<a+L\G&HRcG>:@Y()0Ha1[^bZ,37.cEUIS
Y[\e-8N]=Z,.aU7FZ+A0MP7G-fN99a:5f7C)O(Od@&(P;S5CcC2]F4:g-d[:#\f-
<6e9bG#@EM4XH4=EKeU7:0+P#V]e88bA9Ob[LJOC)XE7#J3ST_+Te^aD1fZbJ,-5
2_cIfXXZ)9H0BWMGeRLfWDDX&&>0<^;G,_,[XOcSR7>G[9U2.?4_IY9P=e]>WA,A
fT.EBQR-^-=W@L5\QCba3_<MHA,]aaT5<,3ReQd]@c,]_UCb<>^=OH(?LMB,Z@40
6Xb/#e5cY?g54W[E=K=386^4/a1MS_XWAaRaPV2:Q8[<8V8?6e78OD5bF@f7VeT\
H7d45HFD.VZ,OD;R<N;1(1<96BUfG:gFION)ZR8d-2d]?V6-/I]1)A\+54S6CXKH
F^AH]<]#Q\A&/OeOJd<M0Y<SFE8&D#@&;NSaL5dcdd.&@/_3f(M^V]ac_C7\^]b7
&MHA81<W,F@5cGJ3BO=8\Q/>IQ3>=?C8P;H_;HPRM&4((T[GGC.3YR5OC3=b)R)a
9,VI1A?@bB]E6_e)e6TEJ=N9L[EH6CW4ag_WFB+8?D6ga=9e&Q3D6CQTE#=SAfIM
4Yg,NHPG1D#LA\T0I2@eDQegc,aB#1[N@?Y5V48R].W]E-J/_>dM:JB0GN-NgLL6
A@f1I:g;EHLF]Da93./0S+:4YOE#Z5IMB]L7D0XI=Ic=N]]_Z>X.CRSS\M^gS1]d
A221QK;,Ic253]c6<Q[C3adVRXCT74Sd7=NT7G?A7EM6;L(QSO-Q_8,f#-STSCK.
H/)^FO(g/3<bO4BEI\GZa/AJd(_3a:):B8WB^cc?.VB1fB_FS>-ACR;:@86\F32O
DcPg)Sb1+:?.0^Q82\VfGBU)dd()VQGFLP17bD+c6]&PY:0BB_Ge3COP#3@bK\LC
MRF;fS<[ObD/ef0?3;e=LCK@@BPg\D-WM([7c__RX:2<1GGKIC\T?07)WKI6/+.]
^A_&83)&_B5a@T_a:NK2,)^H>=Wa+G?QS8\IEL,@GPNLgCbGU+/G(57=F?A>fLKH
[V54U;3/13#+\dV,:M\Q5&;U+GCQ_#>Db/PZ>\[,VB:JaHH=VB(YNHK]E@?8a5eX
eM&>UFU.VES.c#6LCQ)S4<+U0_0>\0L:]MOROC(W162a3DZKI+L>9?Nf6+d9Eb/b
d@>TN(4[_Me/JCFL8NS(AHFeJUa^PUN3D\fA&>MbW1\/2#W],]7/GeHQSY0B-d\)
&04cLe1Lb108S,6_@))34C4P^1^U@=B9_V?UaUI/g;E64HNLZXd:K<3QH#=/4FRT
6+MVdc,KfAcZ7JBG^J:eVg)8#G_-32g?3?+P[V#Sd)CS5PM<M,UC-SNC;d[eM^+?
M/eWI61Y-K.#S809BQ]c83Y(QcELP?3G.&NEX;H,ET(1OZ-a\N\6RWL;IP8C<#31
,W+H3MZb3IA-P6EHf./]GJF^TBI162Z2W^cCG3d;1/7J,+DL\X_K5Y6d?6gg8[IO
g-\:OF]LTc0OfL=2I,cUaA5-8_&A9HgD9YC8OGL&8>DOYfA1C5GS&\9>I50K4_DS
A1fDKPCQHUF6.\/Bg9g=dMIM/&7<Y,+N)HVO=gSVMW,V1;9<1QM,JCg]L7@NW3f[
3]6@+&>+)]\K&Sc+K86I8APG\#1P?g:#Y_EV3.6LCa7@];g9PDN2+]e/@GV_FW:g
b9S7bXB[T:eI>908K.N@K5^.eW4H#JCKSD<6ff7SUAB29bWG_YM(<+WcWN_g?b4(
P=LMW_?&&FIbS:1B\YKZfa:O;V>U0@2\:bd)7=[GM6XK/(eg+dYMG[V=02@fP:f=
RF=:^/1,>XI<=.W4_HQ(&PD(.N-ebM]9]f+KRdCW@^K50D_ZI[3H[RU2a\f,^\?<
V]]E(ERFBcGKR,5C+<=b)VQZdHR@&\,2RG-;ZXFZ_F(b+\3T7#V.P;c07LfgK\6Z
7]KbV2V#)d-@3g><DVG3TZS737UK(6Rb5fK_WLaf#9J8TO[gV=fJML?4..P\-^e:
]-C-D0+)Nc\a94>Kg0g?<A+@JJ^fN>eDR:/VUAXPaJeOUIRCHe1EV(&ZW,&]PQ]E
7HBL-;g:JRYF4TFXdPD=@gP8>:49DK^NU=77^da;)B[5BeQ]&(ITL]CTWNKcae3^
d8=K^JKDVXY]4DCC,\-/,P4(f?..KWLa<>2A=+(.]-RO(G0\;/O]8Z?P1g4dZ;>T
V90Td/0GRE&@PE&fLeKb,A:.U?&I3cada.7=-GC>?<Q2TUdP<f2]@b-@Jf_MHF[T
6b9ZQ/1_^eLG&(0;9bbOF/H]aV&eJKP>R&@<g)J\U&CcBRa#SLeF/SE<0cB(;He(
/A6H:g^/NfT,\/@N5[9P^J)0f_H#9J6/b&NW;FY\=GYX;KOG]e89_HcQ5-\JK8gN
Z447_6[=PUH-8D-LN(9#\I#&46>P6Pf0404>&?\g_KIQ\05SB3G^f1d5\K&Od67K
V^(RE-?Xa@Q_M3U=ESP^G5SHO:C/Td@MLSc7#HETT&34+>LDGg0]/2Wg5-,=YO\@
AZaA22VQAW;M#BG^V/gEdbITd>]EAc0N1Cba@PQ\\5P-]JOT7^agQ&QD4Qb(cZ+Z
Y:d=^LQgDX;V75(T[7]B9NL;Ffa7)WI1Nd;5?SL_efBe_\<GKUB]:Wg0/(XQWc<F
9/?;17QZW:8R62.5YZ&:dO^e0;=:c&3X#-FM1N(H7bbFc,KY4-\2+c<;KW/:c/&d
dP1ZeI^Z_EIf,+2^_D>f,JaFe<UF.<HPDa.M5:Y]5KLJ0@g]IUMe^-eS--AW00+G
TA)^<3f_0HRAg4b9T2AKfc])SacSI2e7V[HAYA9cfRK;B6M27TP:HF>NDI@8Jf7S
I>[H+ADX)=P-WFRFdFa0L1?(UD&,10O#-(P(5]5/+bOCLYg^Qe@[_.Cg^:6\V5b1
Z]J3AaOf)#UCDD,b[N>X#E3=>P,]1\C=TH^Y]<:IE6U?2@)3;6;#.2X0Y1Ng4be^
3KIRfY;92],W]V9)[_J>J7bT/bI8?WUB?$
`endprotected
        
      
`protected
Z2^DO;&S;@^5>/a/<>:MI3Cb0AF0UbE4Y/]E>VRKd[G&eKK-@a<N))H=Lb]O9F))
YN#I8<29H4Vd-aM]RJPe[JCNKOg_::c\Xe:NA=VC5^@/^L,YZ8VEYeH=N$
`endprotected

//vcs_lic_vip_protect
  `protected
BFY<&@1XCM/X)00B5ScPc0b5J#HNO<:.BQ4cT7Qc8813[-BNA7OL-(;0/]e&7D-d
F7K\9ZcO2IbNA../<J0=.<A]SY#2_?B9.R5&B;D6NY1O&e:X,VK:_4EaR705?N.Y
GSU_7.B?gQ=DH@LDYH:8ULJ00=AM@4]Q8,FR0::7_-1D<KD6+-aNf\Xf(GYgQMRU
@W>:Dc;cI)cLF:L=6=LNfGP0&9ZgGCKcC[)EWU4,IOA/==#TaE8M9>.S:=VWQ7)9
Xgb\cY5E(QA47F6LJX=d:PL19VfX^^dU,1)F0Vc];<V@[Da4[G5e5VG(KH4\f&<[
O\#a\4#MCHS0E=[Zb.GG\W-FbfUONL1@A8+OLX1<BN1K&C<=[:Q0[YY2JGO9R&/_
5:7;O.=Md+GPAN\@G8H;N=^Y2<GK>(F[[fXgM](AIb71XZACdc[\-8TKS<6f+K\O
YeaSZHaA/.WUR5YFY><_76V(-26e^);W-#(N.=OA=&T4?WHfg]MU9;f8_@CWccaS
+W9BONfM:8]eC7[8PT70:78P64Nd)U2Z[(X5)e3QK61XBe/TKG=<_GScMHcVQGM/
LROF=)<REK(W+RPKTXR4[@^/3gA[PO511,]gQ7&N=c[0IA)C-@e0K]SZ8gIU>f?<
cG0JG\&UT?fL<cSdX;#FMBL8DBN2,,D?5U)BA05J.,e2K?>7P-X30&&XaDF6TI>5
>a8RAA&,,/GM0/Y3=J)eL;Pe0(EVG3,;Q-/S]GK#(V5OJQHZA/N3(da]Y=@?^0.d
O.>9_A/\f7^T98)9M2_Vb8.DF_b:gV<ON_I6OV6TTVKEY,AeZYH6,W:Jg><5KVg4
>-gW=GUEAR>6=D[F&=(S(Le)KGGJQ+..-J<b;8-[T(ACPD.,[b;6dNPdVB]Y^[J1
/[+NZVMEFY(EEbb-4#;D6C@JC+0SEbPQ>^.1d.7eNT<#]R9#gMe7^4/f/IL;STUb
2:95.DNE;UBL)SJ]b>\=I&LUJLE<#TO5,3Jc9(fac\gCU#1:6GeHI<W7@4H_N@<D
2/T_4)&/\A@_:V2cN)RLNMd<OFY)7eBZeP;GdA,4RZ[E.cTNH7&VCU@OU306eWQZ
Mg24:Rf(035)JWIB4Ka6L(Cdg5>/a\TXZF#Z;c?SBX=.>Q\e3?a.W3L.G_)EZ6FC
BVN^0WFEMPLPeM9ZS6]\HFAYITN?XaMX4I>G4Fd]&F5H=,#c6I1O6=.ObS\7;70@
T+8(JN]WRL.09A)UYcAZ_(PXHZ;K7ST;SB^==Qb>#:HKVOI-/]EQTO0)>e=C+3Vg
R;gFS(6Se?^]><WM#EJ\1RI:U,U=[7Ye,+,?N.WfE\V(-P\f/YU,UMESgHJB.Nf#
Me(]JFW[)3R=C0f,G;\22H-SdbXYOY7XU#e)^//ZVU@a-OeB#Q_&S/DEAd=M0M3;
WUf#ef,[HEW5300:3J(6H[a4QWP9,V\&4VFM;CV7B]=-OA(068HKI5d8+6/2W7HE
1MY0<((bJJd\5gL\RZe3T]=3JXLgW^<RDL>1aL\TGN))\+>100;:T.JX#EYbU]SQ
;O1&/8J?W7:TL52KCO]LU<^cKZ[:PMAN:[Jf\U4W9F=-1^QE7C7efbbcfH.gHf5Q
-\E#:N07>?A+3^J(3>H3@44fW6bMbe2U6XSbE@aX@e)Ac1Z#J\.X2VYQ:7TAB=[>
.#LT.H]_5]V0_=dQ)338RIYI]O(bZ1V@E&7963XF47gZ7YIP1V2eO.(C8Z9>HC[R
RN>4@RN,RS8D<Vf5d1deC>?:Oe36eXc/HG8MQ+afA^I1aF@WMR.fdI/4_&CK\55.
T[ga,^X?GU,<FU(63IBb:]/Md2#@1Pd/,[C<&4fM55,P9EE^@R&Z,H\6Y.CI7=,\
eeZB\^#NgFe0:gJ)#;IQGA=+CUK\,WM0\A=.[9QC#E1O\PH]ZB4/8[Lf>,VBOL_^
/c(c>0g??[ZA@8^:@I[9d9JW@&DJ(E#;H#,[?]O><5QReX##]1&-\@MSCL]BY@:O
3@GR@<)]ML,&IHYV)=ME9CI&aZSc=ZLdCJVPb_)fb&(I&:g<MM8\]L&42=LQJ.8X
A0D,4=Y>T>;O:SKHT\a;P:@J(\c1Pc.EUU[R,P3<cBEdX0_>AOC2/97PM7EU)G>W
>6=JBK3LfU(-eEKe2T6GXB7aD:4b4E+@Z;NBQ10F+68J:</1[JYfV4?Q&3F4gHPO
Pb7a93<XM[[?BSQ:V6PT9e]UNOeFAH6[BSPVH_gLe20J.\8_-]X[#(QMZ/c8-M5a
JZ44ILX\TK@)RVM1WS0E6NDc?P^VI<7+]62=6[9&685R312M])ROR#DD6QMM,dL7
Pe@LZT+7Vc66JCNcL@a)S(c><B],A;d/E#<:dSNK(P@=H8I5F:e.151K#V10//(.
gR#1N;PM]6-X=6(6QJ[?>;;?2/[Y<J9[6&:=.>,&^]ZD/aT)G0-I:X3&TDN)U[_5
DPT,AI<D/DH6c(G_&]W)7_e\N_L)K9J^B]NYGYN[bQJ_H7OE\;&8U#,2332P0<d#
VeY/8-L=^f3ISVKJ<b(,;VPQb8].CbXF_TQ&A.N:dW2X]T.&H5-,?c]J,J\f]g#;
^-E<TW-YK45g8.=JP1=H]+#.+M8APD@9NK,CQO-g,aC-#XcYG0P.:V(+.1R-55#(
6ULe6/:.+7Z]e0BcMA10XRMe7^:F4?[X0@6.O=)GR7Ja[IT<a4QNF_&70?cY)aYP
#Y375X@c]W;+V?Z]B7A96fJ<I-:e3N2R:a_34#/)7^BgS9ME\.T09A:.2cGNN@=(
N5F<6(N]ZBeB>41a@U2W6X74WNXM(6L>W#0]H0g7O/JQ[TJ)A[2bY,PQRMLOS2>)
Pg@f^Xd71<P=))G-;6CaD^<GgLIEK5fW20UD0@6OA#I7P:L-&0@+Jf:LD84MW+.V
[JGT\?L^==QA([e:VP<e6;)b1NB^GG&RNL.gb+>A@92?^DBB0MaWfO22-MQBIaZF
OWd8N?.<bU2EJ@\c/E\8TGR.@TgSC2-cV=^d:JZ=5?gNObDR7Q#fdcSJT59-B8K9
]><DSKR?2JP?C97fFbTX#/-e?0U&d_,)4G)OR-]/T^b8GZPMZP@ZH5H\ZKSFPU=e
.0;OVQ;KUG?A8[Gd1VeUG@-5]d[M+_Y(cX4)/V(D.=F?\X)C_[5IO4c@eV,B<]Cg
239/P[0e@&F)GO:.=MY-QdXde+e=XZA:Q\GaWVe.Qe_@\FfXG<CI;5SXM)\b<DL&
2=L+13VM]HfJ0,/cG2MY(9.&MBIg=IR<5;ALQA&Yb6>7_b@\1:WEJNJfUR9A?Q@H
5/>>C0Y296_IV3VC<_gR)MXgEPW7/D4<EOgSb\JU:]@VR6?ScDH/O<9W+;UX:((X
D:0_>0eY(Z7.UVCS2VdCJMbTLGW)<<_B9]f2JKMbfRXfJ2:]G7X2:^XT7F+Bg2E0
U?-B8dW_^-TA8O/0#-CGcEK\)(U8I.)E2TYXcEA#Y53O&eJPOCL9CE.RfM6AMgBC
\U:4,)@L+8+b0[XY+Ic5)D911Z0KF+E0ef7a_M.1ZRP5Bc62D8V30R#Vb<3F;]>)
A#b+gMCD2Gc)6T0#XbYIH]-(E3<G6d)Z]+^C6V,#?Xe=FG<FOB[\#f.=UY.Bbf#6
SMDZ\N:(,4;)9UP,4_3ceJ<+[K:)Oa21L<8@Z9X=/\2#NM8#;^Z##8H,HKMC5?23
>;b(Gg3<PCc89F:,6JcHN>-N<dJ3NU>g25WU,9N^@Rcg#Vg_g6K3ZYV(G-@D\O;a
?H?Ege#b6Z/Ud]K\?(?SabX?G74?EHf\5[0>02D?,5-dc:0/[R[RP(^(4=(/5>G.
O?UR_C:?W.(]W]S5aCRX_29bOZe;F)[b0UHa_^#>Zed]+N9eM,K.S\S5&cIZK51.
)TVSUYXHfYV]J:beM[gHJ<IT[5HY#W./X>>MWTgWe6Y(9B&1We][>LPPBN;O+[)U
Q6P6YJTB)&3ZVXHW:<21]]Q,Z8]<Tf.8,9@PfAL7<eb4PYea[d-^QJ4]DZdT7Db&
]a?,);#0:CD<@]XPA0SNPR>(FC:N&0>0AS[fGOWa\_gLSLc_b>b/7.E=Db^>63:f
.+D:P2AXaI4YdA7f6MW]7\89+dXd5B<fCOcD@9L)?7W<dA)Y,A(?17c_YUPc/Y&]
E/&+(bER<?@^Pe[;NN3&=cT1,8@3<,VDOSQA0][T/UP)]Q&?1\4DT+@^=Gb/.ZNG
1N=M>/0#cI7DI-;Db6^A/H:0e[CQdE0X:+^X8/7)7WW(3<E)<DMV]ET2WR.F3A)Z
8\RgHC,N_dV0UUI=0P>W92G1/eAJL&2^[I;:]WL7]6FJT-7X.=<9KdE_M:1XXd[M
V-:(ZL=e2MC7=cG2P-HYV#IBb0G:5O-=6;[:V02^a,AUF:&CYO#SCCT@E@f.g^P5
dQY3RQI/F/ZX5Ze6C/Q>J;,]If7OcR9#5-[&fD(d[Lbe2MDH@Ng=V\6IF5e-b?S^
8RW^K^=D05^We_L<^N,X@HUS:CbW[K(V&&Y[W[(Seg^HT-TZN7=E(bHORE1d7gL>
VP87SNMKCK,:?SR<H#/)2/8L/?#fM)b>@9XX6X(Y;8G^VC5Lb.CS;0Hf1d=gI,<-
\>8<:U#D39)6c)/1[#6G.6)N,\7G(Nd4@.J3dP266&c?FT/Md8.0W3UB[JLB-,dI
Oc<L-6I7735EC9d<].49#4/S/,&FRMAWM3BaX9[R\9cA).T-[G;@@+YBEKTT-E\c
<@.6G1SCI8ZCJAF)RM.O#E7eTOWcMD?@EEIaVM2E=]]G(@b[#JJLY,(?&E^WX(PM
=e<>>?H\b9J5egQ6S6&Y)c:+gMUeT1;G<-&)\_T1c+<U=IS?AUVWU7D_KEA[_97b
8D<4ZBR<(39Cf-+7M7=T2#J>6FeERI3#aae]Ag?27L];WgKB7e30QD7)V;-Y?3P0
4,>]^AB?<dfZY<\QCcX[&VOQGU#?fU[S&??T6YP@^0CbUbI=Q6KW_<3\8aa8Z_(g
3,c02Oe?3A?YTQD8Q4W53#D(]QPMV].C9UZ.ILdKe+V.\ZQ,Q1\AN/e]SO;MZcRW
Q=_abNCL\G>\O7_:fUS0:EMD,PMf@LWW0WP2/a,A1,-7,_:>+940@,FY/JPF?O&B
_eSMfa4dALBgSa?Y6)M2JDY[fJ\OcG-f#G1\8XFHN,BdfI)7#M,e-FY]&X1J4&30
f^DCBFB3=N-/U7.ED3S6Z@([(gWa8M>KPMURKLIF^88GC7?K0-D@>]FRfFH^TVZ?
?K(:/]L^K]IbSJQ]7O2GBJ<OOKf5>KO>Z:U:(Agf0,6[(6[&cV?@P=,Sg7([&N5b
[+]X1H;TJ3?ENf@8SAY:W>8D/;^SOeV-KSNV(MB@9KTbNB7JK+2LI&9R.V[Z#(3B
V)3/7gX?CFG<.6OKGLNZW3KMZ>P,F7;AZf9SD-0bR]-,BAf(CN8MZD\UUXHNYN_[
R=MK[523;5,P::=.#+I:+-)WPN>LN19HISQ6#5BWWTEaRIZ=HVBGQXL=e(O.@(5J
KR7SBQNc4a,^Tdc7eV(F01;:6^HU;]W#2G?YLeWQ0POJKc,KW,dH.2C:^EDb;6X:
O^)HV32Je97(Of3@G30)Jd:^E1Kc<gBM?g@L#I70PZYSC<-O,5Y1UIVdQf<b?0gb
\0H4(26S3EG_.=I^77>BAZPd)e?/]2a[eRB[6+M](^M.b&+E09aG)P37]9(;CBMK
NeRW?B#8?A=##(-ULO.SMg,TITf/K:VGTQ#ae6[+Qge-3#=MgZ8W9d/G?<<f?,#?
;WLY=/?8fF9)8_G^aP??\]#CN4f\,SL8V\RRD0<gNeeU4@G>W3)SUT#UgSHJ),M^
ZYc9C.AX+#d-1A<+bXX;UaD(.I24C&S/+/:EK=:g)0/ddB14J<A3JO[8\8R>,9OL
_SMAR8Q/:;1&+I)CCH/VAW7B1I83_Dc;IHKf(J,YUR1U+?H=J_?V#J?^B(SV)#&a
dKB>C4:,a-fU.d)]6J3a<QFK#\4^<_Z4LHbHf#QAKV[JM7H/I:/9:b:,c9\bLA42
XI2ff:<[?]cJU48R64?T5R.D[CJ3<P(//1V=O11@-STP&,]&W</YKGa.d0#2:/Mb
A3ZG-BV&)F>1Rd3UgEJbEBV;ffa&\VC_@DXBJOJ,gPNI8MF:^/-4]CK;>Y><@,c(
/1IL;[Q5YS&)1@f2S9_X77-HgE2LJ7a?6dfWOCXMI32G+PQ-b6+e<f[#2/PJ1<U>
&0&^:=B.IUAJdJ^/9D8[e9O7J&:\+LM6AT?^MVFg_2.G>6C[0;TeSQ()ZQdLZ;X;
^74SZ0.KIY,b1-R3F>N<HMdP0e)Q-3g,NecYGcX;.&SBW)Fe/+D7NTOD+ZfA>#?a
JbaKI0U1_61aOWa^[(A-1Z6F\QV:GI;IE(,EFC)>[3&1=eP@0F3WbfM-F#fG5EU\
6LKf;E-b0g4)#EI6<PJgM@8\PP7U5_43>XZ3W<RCX;<Sgb@H5g;GdeBE;BAQP&Ye
IbIbA]e?Hc]3T>I3832S#S4A?_fY,J/JP9KFE@g,(IT+2HW3MC#5Df-JXH>P=0XM
^fQ&4]e&WRHL2AQXT;H\Sb7e<bJNc_G8-&;a@_L/6_d@VT;^b4@T[0NE6F4R;\6U
-/VTVc,PYB6IeT=b-OL0-YRY[1Q1dH7^Jg94Jd];82DbER27N/#<<TIE1/ICLf_M
^A5F+OHd]IQ?991D,2#eSF2:F:59fQg525g&B^=[R?fIX09Pb#,:)>_JDOWgNg=X
_:35&^bA6H6XMY]3DIVB5.H<P5IZ\R:CQ,Y1WZ:1<:I@TI6W^C[9K^e_\RIc82LQ
9)CPgf?UAICf286.4Q87bXNU/?+5A#be&5&.cT7>8I)ZI_dG,5,]TgN0_^?^4d>d
6Hf0Y0L2a9a#XP1dZ.OB_XX1>A393H,8g8dN#],(A7SFaU(LRLD<1;Od@BNW=d<&
fa7XDAQ2&6M\BT2Y.:fS2.\&O29N>/08#.)=gGZ?S-ec6V4=QcQ0D9IJU8e?PcK9
\BJ5V(,JU-WG_Y>A:5cXX2;fU[T7XTA4XaF6,#2)LH(++VFJ4cL2eDB0GEMO&,V5
M.+4JI=><_/-HdJ:bBe6[O=)WFQM.6O#?;3TaKE&06<OP_MLC&O>0a\+=7,0EbD<
O\QXLQN/T8:I[>8&&+87JJ]J_O(=FV[?\IGXea-L>&9+8V/RH;U^T=N30:Z)(?4P
dZJaY]74+[SLQ_SKD<&NCM,:e,#LEE-<;+W9]K[<LW[;/>B0;A8Ha@S,I4;JWBH=
VaV4PL.R3=J9b1V)NNBd_:57FcY.(]P,>D\,1Og]KC[3^.JGe(Dae2gSY,\OKYN0
M<aUN/+A3?&dAWNZ-1VadO0a16(NYR=O8dK]O-?&.H,#UYENJ:,C#A-VPC-^87_M
2#cbf(&BFRXd/D^1fIUKCI2KTKRE@([L:VBI=?TSTWZL_D=8:J^#FeCP:&?[&HP/
B5WJ=L,6X?SCYb4=7:UbNJMc_@=M\+L9-F<HZ5ceU=6,+B<YB),99b]XG2f#W)(f
#@?TTN[4(L=S@\:(>K/Z#UH_a_EZ^7;]X,FJV37K0L_NN62Xd.]KQ1D-&6VU,/QO
>XV3M_P)#@2#H)856\=-eF7Sf@++aC=g8[=44:2eOWBfTCJFd7d1E+fJ:+;#R7GS
DFIb7>#9egS&:Q.PAgXVP>0G+?BM4CgW,&ZJ?UI/>G2FZ@:J,AY)3,LB+8b5W)M3
7g)SJE)g[I#[P1HTe2g:7?^BM,?Rb)AZ+OG2.6R.Q9N0geRFV+aga0INg[Y<>Gb2
[?9FT+U?(>aV,X=N:1c4>d?d:4YcSWcT)H_R5IT1:]2@@4)X880[^R;VNS?:1+f;
=_^)RKPNY&cE\H:AF2MBIK-FC,f-:^]eELR#,f]+::VGe=\ecBb,Re\DZeKUKS#d
X,MG(Id)#LdGf8S)41)WZ=^-9e8gga?f2U09:aeIK&GBdA#GM1>_P?[HX^37.4bS
J;GLO;&&VPD5F78W-@gOQT8Q^ERU/1KZ&;=YKgC&V<MS&c&_D?cF?be?G1,dIXVA
egF.AER@:Y/=>H?(T@gd8/L0Wf2QI<QQ?G:4IQ#&NU.U-g+.,BH;a==N#BB0^S?d
(d0-6P-&+<1@)A?3861S.K2IAPeb#YN=2_;()TN25a^BNR94gAIEINDGLIZa#;Bg
YeE]T#:,KP]3[&TdSUaFY4DS\>:B./36eN,KBQ5R:.XE7O4D16^3NL^>;(49QGAU
,GOgS59(-32dLK??Z1BdWY=,ENR-0=324IHMHX=V,HA9DQ7RV(3:E\)-bT-5;gW=
Ue>WS^8.Z;<Lef80+#P81HUH<^\V#\WR->1cFg[6;TXF3L(U69f0?WL<P]PY6AYc
+K,>6]/B^L3H6OV,YfCP],5B;JYJ;/<8O4f3+HCIUL[_&()OfL278REe1[LG,dKS
(YG?:_fD9@;NASE=O7^[\\W;a?61?eN2[Z8b<9)X^6Q(TI]J6KSP7aEYS1)PO3VQ
L7Rf&P-^&-4+X@/dA;A,2&7OCIXD6[34fdQ0Pc5=]]Z0UKg3_c#CgcE4T_N<+=\)
[,SZLE+D1VDV9C,CELF=gUV>I7S<fCOV<aK:-6NG3f9;(O)4G;UIfCJ-XQT^_CVJ
.;,+Kb\SWP/TS&4&Wc>+I>2Y->:#<>IEBJ[4b\Cd(V^&HeU0IXL3SXC@aE[cNc(.
B3/;F7V>DX(O)=>(dWO232g&QG=JW1DZL[6:=YJ9+SCU1+2KT+P-XZE.C_PA3X1]
fag&X1b:JL&=J::W;JO_DPZI+CMD8/0&C;R]S6MVUG^A:>WU<:dFZ9/5fR,R34Se
P?.JB<L)BFM-:KA.OIcHYP:Q;+UEdS+b<7,@\70&:8[OKA2\@F:H/fP8@@(3G9^T
J)T[G#cUf47b3H>&&(ME;BNA&Nc#C[VT-HYO<WZSP;)=6],9P:9DD1\Lb[ZJFCOB
\9Zb,ZDK=VZR?)H;6=P+3JS[;HY\Y-^8eY,=\&&(,F#8K:a/UcEDQN_SNU+Qg<e0
]8/(=<5O/)F&94P924?JJA@7=FA_DF+a0[ga(:46P,AIIY3_^-[,:?HUJCI<4PO]
dg?Z]FB?>DGbR--b/<9PA.5fD^?9g,Z64GLGVCT^>@-UX[\G@@8\&SCIY1:Q>E@0
SV?e9#W30<#TYI>X/_LGH@QRZ(.@,^&Bd])cR^gI1dSF7N42/Z5aBTCQ;g;4#DE_
SM)7G(\02Zc6cLbDF-7J#aP)e6_Z)45acR0J]Te^TO8Db]^YD:f9@Vc\WK1^EY9+
KD4\+I+g+WML;DFK1/L_UO)9:L&g&7GM9Wb/?+)ROE:a<>-T0;e^JU,Dg+fM,1=<
\.]<Z+SM/8\fXV#J6O7/4[<R.bHO/]cZRAWMEe4OG5]e20LCDaSL7HPPVK\U=[A,
^?9#6(ZE+M(G373YK1D1MJFgJ#1CT_#1&&C(R-X2a0Z@-]&6[fegE)_V7WAG/3Ia
I,40,#KKUP4[=V1)f@@#+O^3Z4P0PW2Y^T_KBFX,HWZfa[L\GF?eaPHHc(A],cI=
)T=5@PW^TF6@MY]&ZIPFgF@.\S1[AL8NOTR;TU.))G.[P[QPFQQ#L4LB9/@+I&P3
X>#OYgZKF16@^]07K^/4-_3@1(#;[1dQfYNMCeb\(/C]Q)V3/U0Y62?&:=SYeV(M
E9EOc6A(@E27acgZ90JZK[bceNB/aR1Bab08IFBY2FYL=L;^ZRgSDD/55c^/]dI3
YX.cQ=b]QY/2S1(1#;;G>e6O4XY\a\\fDW-L,fI11=O3fZbb[G8YK19CPd4?]H]X
Oa#af)1YT3?959Id:2S7)Z,Nd]BO;)OE#QfW?fWYFEJA9;U[@e.HO8U;8FQ2&F3+
?7[>VP/@LPfa[4;dXc>+R4BI7LeXa()[3.JbS4]9ATMe3H7&bD?[d@\SKUcF,\a+
3D^QBA917@-;ZNEHSV@R>:?LVg9^58ffK99[HO&[;GG;5N>Z#^,):G\Occ2dEL4G
-&@5gI>3dEE-)eIf1M_COOe4UCaJB7@]\R6Q1<f,0DG4CKW[g@IOE73e#?.:320A
.dR&<,]C)P/#db3KH#?;7O]R>eB@Pd,Z0G3PUUYa#YO^Q)Me_8UV@g;BG0>6fS50
d]gVGKS#U/LZ:-e5)=5:UUd9)<_b/&(g<);4ZWa9OSTRJ8[SJOI2GXK\87]D=(TJ
6F7BJKGWFM&UFQ/G(17C?@_]CG?RJ4J_#^W>?PS7PHO;1[RdbS#1X83=Uc)#)A^A
XIT2MaSdW_,Q#:&W+#:KW0J&^Q#+IMaZQ)Eg&&<>cI))X4Fg+98\eBaX6^F(cK-PU$
`endprotected


`endif // GUARD_SVT_AXI_GP_UTILS_SV
