
`ifndef GUARD_SVT_AHB_MASTER_PASSIVE_COMMON_SV
`define GUARD_SVT_AHB_MASTER_PASSIVE_COMMON_SV

/** @cond PRIVATE */
class svt_ahb_master_passive_common#(type MONITOR_MP = virtual svt_ahb_master_if.svt_ahb_monitor_modport,
                                     type DEBUG_MP = virtual svt_ahb_master_if.svt_ahb_debug_modport)
  extends svt_ahb_master_common#(MONITOR_MP, DEBUG_MP);

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
  /** Tracking number for address phase transactions */
  local int addr_phase_xact_num = 0;

  /** Tracking number for data phase transactions */
  local int data_phase_xact_num = 0;

  /** Track the previous HLOCK value */
  local bit last_hlock;
  
  /** To track if the hunalign value is changed in middle of a transfer */
  local bit initial_hunalign_value;
  
  /** This flag is used to disable the EBT due to loss of grant check
   under the genuine conditions of the grant getting changed to 
   other master after the bus samples penultimate beat address. */
  local bit   bypass_ebt_check_flag;
  
  /** This flag is used to indicate that EBT occured during address phase */
  local bit   ebt_address_phase_flag;
  
  /** This flag is used to indicate that EBT occured during data phase */
  local bit   ebt_data_phase_flag;
  
  /** This flag is set once the data for the beat for which the EBT occured
   * is fetched */
  local bit   updated_data_for_ebt;
  
  /** This flag is set when complete transaction method is called for the
   * original transaction for which EBT occured */
  local bit   triggered_complete_transaction_for_ebt_xact;

  /** Track whether write data got sampled for current_data_beat_num */
  local bit is_wdata_sampled[];

  /** This member is used to track if htrans is driven to SEQ for current_data_beat_num. */
  local bit updated_htrans_to_seq[];

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new passive common instance
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param monitor transactor instance
   */
  extern function new (svt_ahb_master_configuration cfg, svt_ahb_master_monitor monitor);
`else
  /**
   * CONSTRUCTOR: Create a new passive common instance
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (svt_ahb_master_configuration cfg, `SVT_XVM(report_object) reporter);
`endif
 
  // ---------------------------------------------------------------------------
  /** Initializes signals to default values */
  extern virtual task initialize_signals();

  // ---------------------------------------------------------------------------
  /** Update flags and drive initial signal values when reset is detected */
  extern virtual task update_on_reset();

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the address phase signals */
  extern virtual task sample_passive();

  /**
   * Creates a new transaction and updates with information from the first cycle of the
   * address phase.
   */
  extern virtual function void start_addr_phase();

  /** Terminates the current address phase in preparation for a new transaction */
  extern virtual function void end_addr_phase();

  /** Moves the current address phase transaction to the data phase. */
  extern virtual function void start_data_phase();

  /**
   * Terminates the current data phase in preparation for a new transaction
   * 
   * This method is a task because is calls complete_transaction() which is a task.  The
   * implementation of complete_transaction() is a task in the svt_ahb_master_common, but
   * it doesn't consume time.
   */
  extern virtual task end_data_phase();

  /** Abort the transaction for which the ERROR response is for. */
  extern virtual task process_error_response();
  
  /** Update the trace arrays for SPLIT response. */
  extern virtual task process_split_response();
  
  /** Update the trace arrays for RETRY response. */
  extern virtual task process_retry_response();
  
  /** Update the trace arrays for EBT conditions due to loss of grant. */
  extern virtual task process_ebt_due_to_loss_of_grant();

  /** 
   * Abort any transaction currently in progress. The argument indicates whether this method 
   * should wait for reset de-assertion or not 
   */
  extern virtual task process_reset(bit wait_for_reset_deassertion = 1);

  /**
   * Utility which can be used to determine if the common file is used in a passive
   * context.
   */
  extern virtual function bit is_passive_mode();

  /** handling of rebuild_tracking_xact on active reset: called from update_on_reset() */
  extern virtual task complete_rebuild_track_xact_on_active_reset();
endclass
/** @endcond */
//----------------------------------------------------------------------------

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
EriSVMiYnn/pIQ4KRd1yPwuicrcLHX3+Oa9nFqLuHF/zxdH1EAMf4Lym269VVG+R
ogTzoPdxpv7L2+kCTNpbBe/R8BaeYlx6l4nNzyEmHvqWq+V6UREceVtAJwTiiVSg
CG1noBkBUQjCLOLUzUWou6S8Uuh7uK/q+M1ZiR8yW4s=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 435       )
icVORTFEtTnRV8nmpUDYjdke1zjTIC8ZD54B/vBs5xiktTxzXxIJF/aUCJRSHrQe
Uhttre2tI2A+33l1RXOfNZNQ3Ffe0NufcI7SdRfPQb9GTn5wgSFO48/yex8jXoNX
j33y5CV67rSgexLHJ1fT6xgVna0qRh5M0rgdaqiC2fU3oVzDOgFiVT9mQ65wn8fp
ILRpnZm1TXwdzK2cixCItPUuuGvb8V06ZEp5yLnOAcH8lRi8rVChl0sSnTv91Duw
4yBK9Z3Ps9gaCT0WZ7lWVf9raip2HRM59X0Ntzlfxp0iIkCrA9MI4xnJYl5hoo0r
xyDM4uN0Yx8rXUSz4EJEADObQnYp3wSMrrJlX/wbc1A2WbCMHNvrN1PuLiQBEVEJ
6XVheApdNNoX2SchnXRVSVEPiGMAp4RfxyP6VO3HIyj/ocyFn5AQ/HSGY2dCMnOe
ds2oKETPuJ493XJqmc2iosC0fPCJptn5bN/ZimHUT7PuajIKNRxDkwJnVMDfQp9y
z9JQhrgw8TOXAknNbb0/UzjyrGidEU4A2w0VI4SCzbophw+DILIgq8bSSprI5hdU
0W5/zFFJCtTu9k2bNphdmQ==
`pragma protect end_protected  

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
iOFyzTJlfwmYtYECf22aRPTUjlTVax+jL+0nGaAPcBFKLZgV4MjXU7fdeYUr6ksZ
61QOX/8Hf47EBlQYx/8NOfi+SODy++5pMxDEnEELk2/JbZ9k2EjDAh7DW+Xb+gU2
S2qMJiks/e9N/t3sSVcNkSDEu3DqJLL8VMXgESM+14w=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 4001      )
n3rBIvR4+PyFdEGibuft/sjxVIubXE2oBqisGlVzcZtr+41o4xoQL+QszUI/t7Y0
jfzYcK4ZsRpxynDG1Uvv/H1067bl+7rEgUPFzdyT5o+OnsDkYIuPZ+As3BG0f2Y0
Xvt4XlASPeov10Citerti5lmgFm160BXIAGtaDTn17tLXlQ1P58Lmy5RbC5wJc/8
Tw2N4j8e3Flu2k7k+NXLuJe5OC0OqMQNgUFWWOpyEEpDs4JY+O/agCyPxpk8V1OU
eYhfNohFZPifcwuoLn4ytq8TMvh8n0NsM89j82eJyuOX41BUXyf/rhtG/1JhoexA
HasLlhHrQxUtCHa4gohATyce8zduV8B+0SXo/Rnj0zvE3uOYXWgRxD8Vg92CJ+kh
dl4q5dpIlJKvsGRCvsjtMKtWUx0cMKQ3Fh9aBEUWn07XLIOL+gNTBTYURWBOZQz4
9JTriBukz8hmiFsx/poiplCminKQhpdcuGHxkPEmvjytemgStAi2RNQWeAToG6aY
/0a+E1pWQ8PktQWzYJo927oVnUsOmbbgKnCVj1FmqorWlqdaYJAV2OcKJAawXfcu
gLL+9KzdTLcybdUexbukPUxDbZXhsNt+x/vGLEWZYabGlpyMRmyxkLJ0cSXcV7k5
9RoYGuB/7hmfJE1hD6easBCfJE849ifZtVS4pFO/A2CWqMqC9DZiKxh6cflHFnoz
aeMyr4aVi7XzYnRysxscjVRsnRpTmDDt6lbwxe4e/QCDdi1DZT5W2nwBRWu8QIja
JQxPzY3SiMknfLrnrfn7aVYC2HyGHeVefBFB8mf/GI5ffMKzqiM5VOUVA3eFdqz4
Fh3OGDiPRe71ezIzFkgpIA+tMIvIfgyF9y0cO5RyLWnNeml1+/ukG/iihYcWMPkJ
rS6LGRFxTvRJ0vtBrjczwp8rjNxFFBx7T9tfs2WRpP8QRO4ouxga86vO2bu9elRK
31JCPv2ZPY1Q0GKtixdvmFg2ujuaQrq0gW4UbvcpSJWOT+E8CR8rDElUTt2l62+X
RL7nQ9Rf0RTVylhSQOQDgEmKFLd/OkMedx9kHn6hMVL0iecsmNwo6SjPi2cOo0pJ
7TZX9FFI4ugbnNwssPfvg21zY76zc1yo2e3Bn3frYfYF7U18TP1QdDwEQTZ3wycb
NTBhfgg1YC/2gmOtvVJO8jZ9uI1PkbMmrGryS0JLwj5oja4aGLYb2xYeK5/opcPG
EcWoMnBllvS426O1SNxcOKcQSlsAI7w6JY925N53GwWrJmeDJgI7ucS/RA+sn/Zs
5iTIWizM+FYpxDpdNpjjiS7x420aFXVt0NzKZABtP5HrwtmPBPtgb6hvOjrjvWMt
hMAuxgzGPi2ifGSbbutiLcsqkpW7x3eY2hKm44oIAWAB1QClefobxjSozDgcyCAc
wk36KO7v02/YBcFtr/Vpqzzp7AT8fzBSxQpNG4tpO4ou/7WpDYd0iPUOBUJdQB06
gC4XuLv5QfqTNRA+ibkvEqK23PY3Vw4kcfj58rh5vpt1vPoVK1J4OxC22SOnRK2C
HSQ5eZ8zgHxh7ASuG0HZX+6x78NUbaAQyjcmeqoYR8bh66o0f7ocmI79MAz757vk
ywLMF0JfXwZYPkXxleS7xhGrBjCdP6N1b12cY2lTpJt+jqGM3H8nv0YvNU9Nxru9
kNn4eUrNIuqlgZmYqqZ5fj/OvbWQylQ+h/CT4gss14F4N8NRW+03ZT8oSu3+kxhR
Wyl9JaVlsP10jiXXU5E/M16hOyvw6A5Rkv7GWQuL083FU2Y5qq3uzwDJDaR0pNzA
54TgYTMIiY9w9owujDJX6ot6Q4UMCSC1onFfNbNodJxRHwtNjtSHWlXK/LLjJ3ID
Hm2RKin/aXGg2z+0fu0/G0QSiLkqLECCNnAqHa0v49evbGff9gK/zG5mE3w4PlqI
K1EfzN0SSHbvwRcQUxtrWocrSAvrymT13d5ClJS6M14i6zkZOhRYK1d0eRnY4Q6o
gNDvrzzjUPN3waTpzrZt1qRX98oOFaNQWTpED17sjZBPxg6pbTGJx5JRBu+Z/Oi5
cGgQ3jpWyNQekQnywtR6h2u7eBetRcbgsJ68ri3Aqp4jCsbTbSdmm0XrqI2AIqrZ
U+P7q/l2i6HnzlLW73zL3XGdH9k86Tpj/uamMRRinzhCQRAdaafChAnhh+KdkiFR
kMJ5WvqqAsKL0SSwekgcawHClyyDQcTBWT/GzB1zqBj1Q4OP4RDp/0IVgUdDj60Y
KlXE9fS5++EfqWXOqysxgvS9ys88OVaUrtowRXF2emjOLi1QUSBk8uL+b/wWZimZ
6kPSGWMqwr3OAJiNIgHSAs35wdff7GjHxSIA22yFmsrbHQs4EV1ygUlQWm2C/j2T
3n4ps/sd3SkLTpbRHtpFF/T/o2M4ib7ap8bUgk7V5NapyixSNPfL+gf5DyDwaczv
cv84M/q/m9Fr2iyfx95clipM6/1Uz+0RNLiNfHAT3vDUATq6wXuIyb06aBDWvtQR
qiqkdoDW/WmP0yQxE5rbdfr7Cv8RSs4J8aead0Q4Zwk7mARLQfkdK5iGbY7OsafT
Yuc0h89RSXpeGs5g/f1OKHnl09K7n3KEfE3a3FOYs0pR8wJz6YDNhzwJMxdksUNX
7uFbAZkzw6XUJ7teSuV5mXsHnyE1LxhgAfz0zCD2qaQmRRtmjJCh+zcQeOzc96Sj
5bWFU+JJy43/FKXLItsWM3uDWQfu4e0oU/0mpzRCOYVnXDL2d/BPFvsGqUyc06FJ
HPZaaBznRpg11ElGgHxkj2Lkoaruoa6BlPqmiZ5uCh9EA3x2cidFmW/ENvOqu0n1
PCHhJzDmIJrosPQj2ryA1rUn0MyJAj8ntgbDkL2FF7Jt72wsuxzgulXjlj1bTeX4
2bWoatTYYQainHigsBpOJXpsfKjrLgnCbGAx+KTPUciqDBwnd+5XOx2oq+h4LemD
+I/oClUb0F53roCxOV1jA5XPliqX4gl+/3c8cJQ/0XqyNvx0bYVKDSxxc1PD5k7w
38JO92F3grld6Rgw2gxOmYvWDRHCQbUQIdu9wdqdsMhq4/9Pur/9VQsDncIowfdE
qsrnvOEuGV3s1PzVjHmAPf6DJ5JtWIJlDhSo29bsgVqM9nUk0et+F2SZXK7GqArT
Ef76a+SOM50IsD63KaYib+kgujk+YsgnhQ29UIWHTrCA8yQXGwUr00moChyc8vlO
8sRSlFLB8EusqVZVtenZ+1/iJetvQD/YENSxfbwitaiAbJoYkEBFxpWNwQn3881k
TWBat7FPtWNLlk9m/sLDeZewbfk1py02ROBDY9X7qXYudZKoyJLdq37mSOvMvLzC
9HL9S4xeMRNgfAMq59P3dJKuclmDrlSwHlRAtmZLDYJ6EGNPRdQYcL0Z78yEHc61
FKkkJZjok2dVjKmdsS9IPTge3skzeGuTA995DzZB5tibhlIqa5apa65+x17aLcGp
ChKitNZC1Mhz/Jm55RNgt2FyFzD2yTX08RzguFECgdm4bOEj9TrP+UvMuBvy0bO3
qq+KccyMKQX53B0fENBnK3jj7FNfChnXZPd7X9tEcIYEhOyCHF6Y5/yvqhsrcv6A
n4D/mfckaT4ingoGfRAJNHxQdgYlD/Fi1slgIeBYetxpou06Obvweq6Moxb9wyoY
QUCN3YVQZAo1SILRGrTqYQ3SOia6sMZP2p1Ni31HjWCuRnWWvLtpHLu1dJGKIGUT
e1bDoF11uzLiesTli/b7Y3hZzd0yV+gT/3zSbebnioDMoY+rsnxq44Z+RKQbCO3F
BDBy0CQDtq2W1+JbiFaACwdSsmbqm1d52aAvwowKgGOPos/G0bo6FQxLQZytDPiw
neBCAe+aZbEo1dDGf+ZOZnI5XvrZ+js4v1Rh5oJcMA4aaC39falxQvLAROPJKV1J
nOxSYMNheSIp/54Vg6sW+qNMEShH8Q8oQI1ALjwH1Kz2OYEevUf+q/JuU32RbXzV
nmRqyTkodT6mtuup26zUGch2Wpa7HSWCR0W0bLDDyAC8g80/5UNrj4fHQTPwAXqi
/V+rZRRrPa1suEmqIKaGSU9bOWxTUS9ryX7FHmGz810DvTMLmf5roufnq5IxK1mI
gO2lwjwSWQWjnJvC5/HMgUDWjXmiZAr8UDguINnx3T33+vM1zClllSdqVkYJu9oo
jYULkbEByi84PXO6cHYTRBjwO9tSAydFYAJMWV+rwVuVwKcCPvDJdgOzaSP8I3kL
iYYjdetUAKc7vtB1iZUSu0C+OlyCLj8vvMqaWLjYyKWcKWVhYdVwxkcUYpbiKwa0
fU2xFvuUUquJEIyr1h2wiVoh+WzPIZhrKDpNc5Xc6spYvADXp+xc+xCvJPD+iSGj
xfV/mGv5OK4VuBKDtpfR1kFtmk1XTkFcBIZxYG3+7uPBNxeLkwRdQOC3x8mBCV+P
E6TYZVb7IFw9p4RHAuubQU3naCYBUhAzUU5ML2vQ2V86hHs1Hdr+wks0rzRwM9NY
QQ55rF7fsRp3HeGKE2ZBl1I5IaW06Kl62+thrJd3zGB0v3OZiwVJ39gRIAOngJRS
dhM2/2/KtGbK1vDqeFHIU5MpVqn1qjAz0O4E9YK4ZTo6Q5T+7fOM51xJjWcUje3S
/+wiiRdfFZCHK9byMNkNNBb82QR1ZhasnZKN7M221i3d5vFqWkYmeW7+UTPLLVnO
F1Sol0iasXZ9NCnCBTWlMwf52Kz1JyfrjvxSWbpLh2BL4s21UHh/ytvEnmn+0JLz
YIWEWm/5/omuFTUGOXPODQ==
`pragma protect end_protected  

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
g5p5CwxCNwhka2NzJi7Epg2+RuivOi/ZcyyakfIq/1+nIeSFiQf7bKNd7jgMYXSz
XoOwf7QC+cgAVfzZLzExsfgZi7wUC6zYUk8LVbXG9q7dVNBoA8zm9deh9B+OhfBM
ovL6kfs+uIMO9s4QydVUdW3z9PDly6Kvp7WMM+23w0s=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 4287      )
WHH7e8XIgDEWtrf44jnX0WVbE4mcUr83jbi4DWdDhOFcwmeS8ACD8Rw3NArvnk+T
FTfRN2kUcojjUdOqGD13uoocXRfIFIt9sjgmVG8jDDzY30HJn+fs7DUa7mjKHdK4
44zm91OL27R8RsU/Wcp+s2Z/gIXagX18KKJg0dAbBZJ9RPrM3TBWs+iGMtaxJ3gr
/wG/lIj2bbvfQyRptiFfR5rCXwIZcj+uMcEoV19BWCl0RtlvIx0y62ezY/QE+V99
8gWa/+Rmk1ujI8n/yaYRGj2/f6X1ObJmokxXBimlC+f73QvJ/4/lFbkHsXUzt/Wz
yc348MXLdlWLMLby7V8PLYrz6osFheHF9oDJVr8vtiVW8VpT4c2ods44TiWT8ULR
`pragma protect end_protected    

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
bYtc/UB4TTqol1MvNHO3+dKbXcKi9PiWDE6c3qJ/XsLxwT6k0QXmTAFyT0pcIXE4
ZoRwN1a4xnKA+EAzeMwbM6lbR9Ae/ZAqoRzs44XMzqpcQaJDI8iW07p2r6Zgcgau
rQy3/hlbZ9/QDITlxU5SBUERz+YkVfWfYX/xvLo27JE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 113129    )
qhf3kvXPjKbdglxJgAmuvptMhFLnKJ14aRIHr/gb61qpAFlF4HqjdCkCTADf2dff
SccTdwNsEqwxgsu85T2Yex0MIV6mfXr3yOgZuzDtt2MS7JcizbyB/fySFKHrHx4c
ih1twZYBlRdPWya4hTAJ3YF7AnQdDm407sQAtGxrGzSV2iJTclUJ6qVkJq0/7VJK
YhHFmAzSz8T+PksfYdsikWr9z3iNLswFcqHX2cihbGRx/f8i4pIVVHHMTZkQlKyg
zeweXXQTsD+8L/aRtBSQd2srx6Ni2EDyGaC6SF2jzRopUERYG6MXJ5U5blmA7wgj
ygay3lR9mmnhAABNN6/Hd3kFUtaO62IFow8bXGea+qnKc1zkMNqB4Bb4f9vsAFY1
4x1TG3kjZ7zh5Ii7Zq6TMYk2hiVv6Kqu6rfB4XMl/QJf/RKzVoenudu3Cavw20O8
QEdJERMbs+BFHjz5nHl9WFANDkEw89pQ1/1DByBD6GenNPOkvf46pYyVloHLE7e6
+oQ9GUpzvr6kSLJ2ATAr0KMdD70IotoSaZ4R0tCG2fCJAW5EmdeGAT5QfZJd+Q7z
S/nZlhRNh9lIRfKX0RRC6kVKue/6TciB4gOifCdVcLF/NxhDt0pb1yhG3mO8+PYv
xCxboeorLL9IX6kcQsDoVTqFGbFWQiAO3NfbkJGdsSy4TOXGuyErKaaGPgwxK6Vy
r2ioZKtrCyUQqV/eFosmukEVKSqysx6Fuuo0xvhzGuBm8p4Hl8imxkbbqUxGJ7f/
UDv/Z8sSyWc1NHRUVUlLyakJKEvy3CMX+gJcLQAM4nenY0MQ2M48Jnz4jxezwpNu
9AcXeb6BoEDHlzNzBfkbhju68DxXmFQy/CWuPfd/GWPXLE97XaotDkI8X7pwFTLp
be743lHake8znBk++pFiCd4NtrQIIc9NZjMH4PLjWBXMGkfi2/S2IOWYaoLSYS7e
EfRA79C/GkeH0YYtyeLWijC4DjURofrGQ+SYJbFbe/Jih3nuKySsBgpLOqWpe6HE
fA/XJlqDPqJF1XZY1pbUCZQ00tVI6Q1xcn7+H1hyxf2g4ihusuA0yah5L95CXmBs
vteuRZU6a9unGSuwPKD2hMVBlKMMNVCTAtFb4SkQW0DkmErQUT+PV6ZRsuu9BEWj
nOGZrgfIf9D/4HxZhJjarosNOjeRoGPFnD+gPdAPWBuGOUFjdUw0DYqQHga+qrKw
mPBJabqfw9N6rYIDHUCqK9omObfaT6XVUcQf++eRY2+XO7wzQXjUwhyiXub4n7KW
3QWd696sDKlNdfNwHbPtZUaffCUTYypOG/eXB1/4yQxykqiPgab2gW1XhV5qFDlL
X2DfN8mPWOb8qwdLC4zOzsBNmOKX+lGHEHv72z8yQLFYn+D8T0KkFrTewtrDAMh/
SNV2ckF13gx072FFjVO0EJwf/3UnxKvyEbDMhzRxcTfL7kok0YHp1zGthuqjEENf
l/RHkkpUfn2LLtr8qAzkzBGjXHwLtJ0RhlIqGzpXNpbkFd/WnrMX9F+FJ8/KrxCS
mBojAQh/+pQAN9oIhf62VKKLYyeU7PGiqdbJ80tv7+YHNETnzYsRNlsWfoS6UXj7
qCbmL85W4xLfPq2g3YYPKugKjQBDpq0NpBDM9nkUj3+I6AOJvF3WKDz7yu5kI4JT
j8s0MpRuQc9SuUrX3vTtuwpLrTlWZ3C3F2yolwknvFdAuxDBW6Q0Uj9JAAn6IyyA
f/4LDyFlCM3cE28yWGxHU2wVtrQGhFsGUBT7T0uwYJ3j5o9UiJdXbrKmHMY3p/Ry
jTWOc3DlwRtdkuQonIzBiJZ23buyPVRU1aPsz9gJV1pXnM6iSTPpEgsfQZraIv3s
apIx/S6DDZtca3QieEuUMKlImkXWaY9Npl/rdHmD+5XhjxvoZhJ0QETvZwDLwPmK
31Mj99RqY5H7G8gyXJ2Hsumy3xR6nCnLeV6Am9myuEXfMkefxj2scPKM3QDk9V+f
Rnv8SJgyB5WvUspAbdHDEiNmWJdrXO2AAG9dwZU3yG57RqGxFoBYTPfr6HLX7yuG
VoD08wDpIs5+OTdCMTelUhBh00fSl5WXZ7TpBceuBsJICQ/zWSZ+eEBbOAPC7l99
YnlXzxhpYl9tFBK7TgqcEOG8Pyj0bVO3vVw7xNgB2Ehq7FKDAv0mPn80cl+tWooD
QmCSz5c+DYYAgsYcwGjKytoxx3rqk2jxFWB/Kkt1sZqZEcA082GkWGhmHqsQY9of
Vysm9wc0KE9F4xYIj9hx+6bIuPjkgkYSpdcMjYoX3CGRRKD9Qxn2g0LGUsgT1mUX
/9pX8SeFqtQD8vkQhatL/3gn+KJ5iTvNH5n2qFAB2jAJwA81x/VJnw1b6h7SdQvw
rNsOrgiJSyXxPqFbmxHNr2TZ4ajfBmYsO6/0qmxilwbDWdi2x0UMYAacZXGg9XXG
chOlsvC6zWYOEzyGM9fPHdhUskH/AAcMZwO3UJT6GkrrEcxyVvL+dupKeCh67+4J
f1LISUGwF8EBE75k2/gmST7BmOJbw0uvUZbOHMjV/Q9E+4dUsASImMg31bYk77Dw
2OC+bl5wfnhSl0GxMkbJTxrZmc6oTI4ZNdA9hRCjBFhlQEIBp52WM5m52RP6Y6fu
FmLVXwF2ztL9TwWFFg+MWDbbu/mC0L4BEGBLg7rwJrET/aCeKdTVHyOBeTOhoUV9
Qb8KPsHnP458WDm+EQHjQlg4+ovZU/x7KHXmHtulQjtBRfdz9qMEE+tRaHg3cFeJ
5OykxuFDI1+x7qTRX0R580OMywTCGw32uNIsV6oO/7QsG3kpM+ru/+e6E/Umudsf
CuDiX1iYnYqJ8NImpN2IqqqiJdUEEVcQpZtVzA0p/JVeBx6T8qSXF83Clw7F6cFG
cTJAppzLeq8UVdY+Agb1yH1HUR3u/u0pypODH6/jTFnNFLZXPpj6AA3IuAYHwP7c
rj3kISXg6Dpcps7Zd4eF9cm3n6CSaLUBGqje11ItF68xWjWAB0gOlb0WSWkk67cG
2d3jDOiRhxSbQoJPrAgFC03NVzf+Ye4BYUj9dqLMGcO81Zp+vSPSEx5RepqxI1/d
99pcXFlwh/DOzXwuos3WtjCno584f9PX9U5bDwreDIVPEFKzsB0VLfZ2uD1f6YGs
Yk63oap0ywjinZRl+qpkIvuvrNNq84K7u+Z7PRphkVvsLRpeDc7+0fNNrzU1gY1U
dVeKf6AEeqJWP21z/+MLkAulVAyy8EzUQrHdikrD1QVkQG1P/zoV7s6SkmNfzCpM
WKP52EdSCpkW3TmaMoa62WTbQhGtf74vl5e34qZKm4moMWfME3uvUFNW2TiD28UP
fUCs7Zutjv1a5K5FNvMIhvrCSWzV29HWbfeHkoDR4sXIcbseSX214+zMFRN3D1tD
32iXVCaPrDmbYvvKC5cvoDfHLRUyhMhtIxrZYXTVfPt6WmfN0DjkefMcD738qQL5
EZT7ulmYzjImadeyH6akZKr6vMCb8fhu2Bq05R4UFloKKgYo1/BxzfNfy8tlFZ1E
R/E063pMc2UkVHtAAXGvUecJAFda01ejl2pdg1OKAppwc8JcUvlDKnDAri/Dfpn9
3d8hygbdlwGqxP6kQEX0AH8DyfPhcwhVo+PDVzIP2BoAWo9u1Xz5YxpYExn0bWtt
cZAFVGW6r7CiaA8Wppwve3hG/BECjkTV4Wyxoj7HGXYEJcmwF4z8KBMNIOf6ukBb
zW9yWHacEFreN6hLoSQCiF/QBiGOFTmI7+fMbWz2xnyAOkqjhVq1HesOlxKWjKXu
GkqIdqFvPcgsbEOt3C27WgwTZG9qbDLXS88gWAxVobOEWXDrRFcAni3CEnkowrw3
w5cHmLwtq0b5Ik4CsQVk4PJCb1ljSMhWZqfDzofQNjDJaw/73XF9qVqQZfE3p58l
hIL4Y+guc3tU7ZADrRPi8wzl3sN8wolsp3EBvXkOrADWQXEEVdfJC9jYLhSUV1z5
dbeCmPweMaKhnLHlkZOj8jtjS6IarHTYsexzwHQ1oa7mc3v1KnhicqgZbMqAHyv/
O/ZClOy0Q2cWOLFBf9otZwJ8Dy6CZ3tcuYay4bWLpqF/n/Zsy0lrgFy1sNanD+mc
UXNvrYOIbTOJ/gitxPfg56xY5A/v+dYa+yeTFIAJHTi8qdV36r1lJ8YpDcy23X1D
XRak9i6hWgc02sF4C/errTQOjeIyU2MsqFj1w1RhRRMFQwe7CjZfefWNug6p5j75
p78/jPf6WUhPso/SRBU/5PRP+fl/kRWy5Vf5j6QixC4RSvUBkmhnjwTrpbmiHvir
7EWpXKQiVf0iJXwNlV+Zb4BsA5+dG0Ts7MG0uq2+Rwtt0TX47PyOI4jkCOkAtoFw
t3W1K4yGYaaRGMly9LKQQJM+rYdrHD0JTQNwphhbyBUpwQDW4ykVPjRLlXpBJPUH
JaUGpHRZ+vp7xBWAPTjCyfNyRxcociugSiTpupVdFKDUEa1etUvmQ/PYl6EPJqWf
m2XXphrN8FlbxJDhibOzQ57AeZhb3YFxYBvuzrJ82OzHDvv4mKqohHzBrnbWuPzx
RU+8bnBchQZ+8muPjA8p9wVpackZ5BmCzr3JhnbMneU8QbQtYYUAZL7ETTyjP2rt
KrNO9x4Jajp5lOah7zq3fes3vjAH4zy3bvSU6t8wary3qME1HaLQS53D4FxVnBAx
56GvnlD+eR1DEs+W1IA1ASIBI43rEGHvmDSV5DXEwmLRStdk+Q4nXV/5TxH2UriP
GnJAGhupKb6ESaTYhSEYPCo9Jx7VmEnxIdDnsmT0tYBuYwr7GNWP8lMZCWJxQkuX
ug8h0kpv/Zzi30/ilkHAJ995MnvQReL+0u46S0rvACj5MM8Zeoi37VCWs2lsESCz
0UuEgYn9UIHatXzcgnjD+A5agQU1HKe65oTtcNOaNDdbxATWNMHND4Ahr5giOlU2
qGOne60T9ZzAV3yZMlsV0jS+M00LcWCZnQlyI1vK1PkNV/ZcKHLyiSu1I86hTirK
Qtisw1Cinz+gyZBenXc3u0+HMeI2KAKlplCi9zyYM1bEL8wgcU0RpXHh9Cnmm+cE
3gLvMqClNulzuJ5F7piMqRN589yp+CNB0MO/YBD9te8ao8hhbPJvvThzRaydffMi
wg4Cpypeqx7EH03ay7CG2GdEs3JQJuB2D3gYkCc6FPYBGnGtIml9da/tku5KNt/4
8q6qYQ98slgQ16nFDthjxv9UFMXyBbNut+iXCMcJBZ5EHBP/RX1sSaUo/Nz2sbcc
tLceD/c4hwnVL4JTnhPMXmjVIBRvydqETY15DMfjV3Mxp8PmcgH+jOrqyyaqiJ+6
FisIU8yhVWZHo/zgBRQRvVX3BVVbIRj3C/oUF5pI0MwoEefnhv5dxxEpuYI1pQWa
YnVnd4qmEDOQmN8lRMz87KKlovHhMf43fxgbrJLg5xBmUOV1DBBvFRcaUMTMYriT
3hpIdRGQkBTNzOJAaUB/TaZwj0mRVSvMHaxUz2uHuY/XGddeYPk/ZcjiUOaMeKFX
QUYjI7cL/S3+J14lrQIPZLy66JVQzsFQ5ijWtl+t2aIscDogkhX5NvZSGZLJOe5R
fTZ67ItqeqibKpqIDXZeOVGkzAht04xyG0rynfPl99UHp2NCofC8wfBhGJZYaT+j
sBdkscQvhw1dx2av8jD2hFdKB1DLgd/qT0fswKneZ4cjH3PHqkTAoxrWDevi83/S
ic7pE5UrsbTD7b4+dgkZBOLctIQeySVNLL5od7/1gfrkC2CLQSNlXprAD7i8IwrJ
n/+0KIycrQ1T94d40zuwPY+mma6bOhGdssBp0e2Ab/HSgfVW/ketRDSX0DJNNxyE
xx3ClYXKXG8CICAP6aR20sgKTE8WH7AK+dAeX/iCBrInNVB3Gr+5IyMojfYJYelI
DhQvJHC0wDoUiOUONnBCzvg1b8DfKbbty90QfikjyvuG5I/VSe0scAM89vHZ+6GQ
INGRtqeiktlWpk79EOlm/WD3rAmhhDMgh1vKLbbwmno1dV/h+D4GEGr7ZDVULP7r
EJDdxb6QDSYwnvrMxek5dcuh2orEqbHig8EfMxcbDZ/O9fRtRVN1AF08UYMj0cQE
6pojfaRMXcT3G2L4CE3s0q7BX2OBTF/B9gyRkKRX0JsJ5si1hFSPXKn4VTAFCROJ
V+t/hA7EJRW4LIwOAegB+JUWZTkUFaJmNZqm0+94FfnoAhNWJ4ZIIF7uCHRlnxEc
Lmjrn1WuAsFOunomgiaga9uVJhxsCqX/ET41k2WhOu7LnbhLOPEYRj6bM4lQyL1G
gFJTGMo15JY1RT4tvcrDNnbsUK46aJggKS/gJ96lyjzNaPs/kZCljrAC0aKqTSXp
zkVtHF455VEW9YyDe/POVbGoP4rLOT0VH7zhfPjP2UBTui2d0aUgbwEGpSskgRVn
IX9/axh/RpQtac4ucKmQ6EeJ13WDP1svCu9rqB7aFBz3PEuLqF5+qwLzlx0lYcXn
R1Ty0sWdMaqwJ9/TDXC0Z//wXoCkZOgNLxkSQoZGX4pRZ4EKYESwudX2YZ+Be//g
LPh/ZG0OafeFoUhQ2fU7kB7eHHqCqg1Ghe9Y8Y8gXXTUIj6eHZquAUoOiEBjIjYt
Fiw9W5pMC8CqhIzCqlm+WKcPTfZkdVAJtEJNLsLQi9EKJYOnmQzYCWDjv6f0kZai
iUGJfWOH1jFV2Qtu9/8VfC+JDB01Sob24YHP8uG7GbQkzcSUjNSCI5QDPNSbMfiZ
WRUdQAx+W1TeALKV2nCmyhFjkiYeQ79if6h0haGsWC+HwU7LBY9Q0Gzoep1NVtF6
xSLs+ypdTiKa7oOXfWoYlgoSpEqzzw5bOet95ow6WMdcr5IS0Y8r+8qAvuwNo2I2
bHkYbMHvI/FAHKeMZ8unjbOrCmIb10yZqzKppFPIlN6UoMd4g0i11iUm96ArpBxS
aCpn7fx/+PiQ73m9RDOwKgH8HDs7Td3jtwYPbUK1P06xo96Mo0xZW//S6qxmd8N2
3+NZVEmFIcoudg6sVVNOGCbHOvFMQQZvpKiiyGDLK9MAHnU4gAfPB15B6beBnLLv
wX0Qeo8Aw4OhqVuCaZ1DT1U+iWqKv3qn5fbpORDngcohkCp7hTQhwli+O+xwC4xw
3wgmVxDuwOIyFTXQVbDe9swSZNl9eocOpUQGpNaQRy2MS5zWssyBqzDRXwP/0Ssa
pFslwZ9pznKE8V1MdEwsNyfGO6is5RQRPG+DC7punOUDEv6q3lmTHHni5nT0YzdU
oO0hwikSJuz4GUb5vDTJQaZ12det1HYW6CF3fWgqIzOQa3ctE1WHUyo9ggTD/Qs+
h8pA6RMnAjNzUsk63u8cgzFmOl89FwY34hamjRrX+hljjJwBetzH7DtcZ8SxpDPW
VYJ28hk3jcHJ2bHhM/khtVs7We5XaRz8HGWhkgvETlV1R1VLru0N184x2NPecGqI
pMz9f5oPyxJcmer0u7ojoV6MA5Ej84IZyMkK0mDviBBwDFsQdvwu1GsQb1yuHMAV
SIWJ2DtxEaEnp0Q7NGa0vp/ckBJjolfBzdiZLjeCeDlPH809IN3oM6creDjQN//a
gNQSKdP0tzHdDgyxh+3c7n72IWauuWIo5K9cXOd3KIqtyLo3BkLa0RYqh21ovYzJ
2HU3hT4Dx1pRN/HjkLet32CyFn0hyqQRIgY/Y225ZfOg7FGgY3OAtl/iS7hHpUX8
T/kxBjxVUPz3h5Umqjg6StaGS5W5ECPp6gFBE5xRs60/PS23fDGUIBsQYBRfDIW5
cVIYO/8QzsKztA3s38vxfSAFjeeCbDXE0QY7I2Te5vhKUqC9jyPvsXynKoKE1+ta
qbQRBwHWVOP8f+15953c8NZiLBflB4JJc/QjifgSdQO1bXGQpJ5tc6VSo10G3IXP
8CKLgeqHMBAU/Y6usHKhafJXDbQE7m6o2xlnFN+o5yukhXhAEst8wmskTjym/U7X
iCdxKnzZd4HvFaAEnvfJu8xTGKo6mZviO0RmhiixSwhv+8o4ECUC7gkiG3AbREBN
xLklnn+yx1N98G59jny4055BJYexJ9UVSGX3CWHK2ZSA0v9UVV7IE4MsL7JHGm36
/lqKMq2LTuLgrrPAOpNtZmmKL0bslbN6LXnTwMKUeRSAEo8jyUyZZoRulc7/qC+i
q8yODQM8wG3gHEHFGfZoAXh6qQFbwcou3wH5CYJ6BoncE7XSspIa+MJwaCq0x50w
34Y9ljOOiW7rKNPSlicQTrwisavJUle/MhS0bkiy78OQqw7r5rYyktlJdKBHDp26
XRcg7wce7qoXR6DhoJseSsVCN4IuGySXdCVhRvf0sNSIrJYoK6QtDFnWO1DGyobf
WoCMAhQO8Wc4PKq8AcY5DxxHfvZbLglVzsHZMjUCez4Zjm7YGqfB9FNyMjoywvV8
LmvwHuHxbwp28kPtRg8+BOJ8o7/BGeUM0l62CBl6rbXDfNYVojBIeC2y2cTL8DRx
PlExml1/Y/jqhK0+XVSiypzvIQrS9xsfDj8HUdv/dd7HJJEbkAINQJXTFWTWcqyP
6DDQbxovogqbRJ8Ceo2zlEtc1zPSrjMDDsfeGYMdHhFPIi/UKfCYRRUgNS1oP8rv
gguPdz4EBSqfeHxKT0Ewa/TfszYrRsOBcRpGR+kVuNwTpXkJBBt+vgSx1klD8GkA
W1k2swIptOxfrYF4sE3KMVVm3pd0l1z1PHxxThrc8y13DsMrva+H88AJXNbLPC0D
jtTyktp9Eeock+0vCGIVKtxkSfQyuRzQMP+9fsItQ7MqTKQYw4UCDju2QyTqdlJn
RLZgCqPf3/lIJozbR4k1ABfpZOZNv0tYGzv/Ei4szxFtB96y71cMceKye1r/nbV3
AyhXsHzVFxpE7xo+1gwYonJbML7KrezpmJymB+pDgrdwBcmQATvn/fQDEWZCjhud
vIvizl6Ys5I8DnP0NyOpXFNZt0CCmcNpgLsxDsBwIv7NJg0Cbbnbykfo3zzMQpun
bgPw3OjXDttEy+mO5RfTpa3g2kyEjfPOjq4C8QbRvF5uuHWVqOaoA4L/+blN5nQz
/+M/ByvRhgJWQP+zFkt48aZ4twS3pVRvaetjc0RGEtfngZG89UCz0PG0d6hh9bSN
T1yrtv8O1A+PWiiva2+biDxnRyNXXsToN5DBshSfacVW4YW2t3ZYaMph+xlXHDlX
wssdgglxkqFjFzZ+zZyYR5LjDgvyfZb1HGO0T0ePe9VErX50p2IhM/10gIMUI6yY
j0eDDUE+6Ct9T33fhvBQ+R0TS2ePAg3DAQX14IaihhPeYnP1iS2eNLnKJhYjHcNA
BwF+iDI4SY473PUi2wIqy6tsjJLDagIqaTXTRmgd6P44EYoPcgECCNPZKp0dMCpS
QHcbk5v8bG1QSOWHbuTOq6cBVGgabaNaPCnDo5mKfm8xa7KbaqgRMkntduJMcXFY
dKWMX4iMh06OBgSxuf05+oy6UbU5f8/DLsRHWj2tQUnNKq3dklNBjv+n1sndrUoy
oqYbo2iwshTLGCUDzUgug/77SGvDk/QoBIfZ0FV5PC5Y1TB3s0JQu6lta1SnuFzb
E0yiSMaL/xnjEacrOUHQ4xJgTsmXgqwLwhWVew7VpDovz3MPuMa4Vlh9ZdG4/Hlh
X5zdolXS4JWZ5Pv9xOkgsOhDpS9iDLCIcw0MdYY08JTkwvfcgb03pb4MyY04AWSK
uMo9Na30PPVh4qsOfSAJ+U549LK/xRxSWp3rGdofC9KjpXIsbWB47ln+WrIQeW75
6y2bzCmNLGOJ54NFRJDuAMqmFX8sQ/lu+PRJ/RpUOxIsZGbwNF7bSGUK2W44cvim
cnbcd/m2RuINauveJ9XuWo1t8kkL240omgwuSJjxLM+4KuzJZZNWNHyiv5ev1Cab
2FDHQ7Zw4qKxsnaN482kUFqPzRi4fubM+GK7mugabNWn0wgwYeRTS1O/oVxRYWSS
bmm4McjXojrydqSFwufNdi07KU29JfGvET/LEWDtZAl/KMdusX06C2FJtBaKS3O6
J+dcYZN/KThQMuay2E8gUghQ4v4fyisQpJmYTL9OABHatdW87nvfld0r4mUQT2U2
pwC8dHjXmuD8cSnF9JcraHtMabtLVmOg1ha81FE+DQIvltGkBlC2XKp3m0sTQJsb
WX4ftHIcNIEVPvLQ6aI3N7qNUuYsp5xt4EsJNnz8bDKaK1pAubHMnxX8P2lWZZNt
5+TgQNnN+LQeRYb3bxX3yoMqiExCosuIs5SFtf2sMbGD7ceFPl0oTWExME0BWncS
lqi9b6Ji0DYwUnM9YOPlcViHL5FEP2XZBPJG91Ib0S8VZ/YDn8RopfofXyT32YsQ
FhHdKD34pxc8oSfF7XLt0cGw5BXbnjr4/ntYIAIgQgvFwAbMwOrDP5VLva0rK3fw
nU98UuIWj0huUfawgTmyv0kK6K5Mf5DzxajqLF6STj6FtIKzUVgA9H7ne+dB45Bl
HzumWo5vVeONYJkgR02dkzxiKO30xSzmJlM70ICJtlg8MxmnuRBm7sDzmKbz4qGH
zWUEoySduyplmCHKbCBkDZY5jqWzpKWt4Ys6XTO2+E6WXP4As+tYkQGpiD+Y0yN3
AuxeS66oaJUoG7VLShK+XrSdJi5A5/VRh38rOI7i3V4ni8adRQLEPstA/0LEWsCg
QZRkkgjuxcl930rN6jzObR/r4jYEYrALCTKk3LvCgOTU4dtv5SDn6WBqtIA8PDlL
ugiupBfq4Wye4t/ivE2+/3hC50uvvPh5CLXjd1JAlKXlBDDmhKYrHmIKk47h4DM4
NvNJ1gRZ7GQ6a4S4hCvJG21FyN2ylxVGe+Qbb+WcTgXKlTtWXXOuug7NxSMMvwFX
Jhm2ItS2IsBZnuWK38p7fZhwYK+1XBQAwXSQ8cfpvne/SvZyL3KkYotYwPWL/u8u
L/H0rM/IQejIoRNF94xoZeMUUviN1hqfDtE4YZEEqFoDge7DnNvkqAQvx0cfXR9f
XGxdi4d1OYbe8PyiuA30XvsH4HmAlFrfHxFUW0V5LeJcMQ98nPCfk7/hSnPnFIds
4WMXzHlAAnYfz3Pp1FP4JSqWLwPquBEif7iIJq1wQEAb1Bt012A9J+IWz53eowPv
H0ezwhmhvBjcw1+fTpfcpiv6ix+4Gks5utUIX7Y323Hm4bED3hyBwjDF0KLxUnlZ
sPXFVSygB5giSXaHRuwi/T23Z+fmAf+DW9S9D6nVxoAvuExcIDzG3kiXSrIhLUj7
HR1h2341XECc8hnPKklAtc+ANYekgPINbx9XpJOk/zQTjR/h91htOeuZWC906rgf
YZsWuSK4ectfhFa6k1T1LmGQ9ISE0wxws6K6qZNurJ0gLYzXEz16SFY4fyP4m93a
qpBi5XNWzAgeWZIWR6KDmcA1SR32qiZQB8cG1AObe2fZw62PLWWmcxA3nKGw7MzQ
x1lHED6G8vKolLJUCsGY0Li5xHlPV2RRU45EDaRW/SMGCioML7m3q3ZDIDFDxYC9
GKnXwLHbSKXUSptWi+CVhFJ5sBFyNfAbuYQq1eCFchkYPJ346aqyKkwmhnbQEOVk
SIxuqcFAQWods9UWh4OqEcXlZeQasbyoSKELr918f4q1Zaobbs/obpC+iddyTZTJ
1DQ8IrYD8nkqLzHQ2E7uFlqzh6ME9I8rSG1kS/C9n8gTxjwhkVZsYSWd4hgznDsm
DzWwaPIHOLDsmBwclFwXNB5TjSmG0CWJLX9dIe0PSdAlyDuH4YiPv3vuhJm2DSCq
WCJs90vSV1urVQCKYXjEKhbPv6RgdsYAWa8+bG8sk9oDZOQCn39oBBgxjdHFhL+q
7YwHlHicSZp0K3P8FOjFCKbXEw+GmMENe9Z734AgxjrSmJdah0MIatHJbWLYondG
F8CQ08Jxff1+QSiexq1o9OvfyAkkHSgbT9UCJhZ23kb0kGr6BPiS9SSqzOVNvwpZ
0OUBRBDxhp42LiN6fIOcQH+WQSDeJzgNnDhehcZpsmOQYda/NRB11r0R/x8OeN1Y
fmlRNQ1VfNcqJOmEG4ZODLpn6mykDz4BTiqrMhxBOza9WeleC0BPzOw9VRPKjCii
G/B9uw0QgvxqeAiRkGSL+MK9hpbxidSTTaPdspEjhXH5h6m4W1bpEPT4HY2jumXo
gqPZoAh8ltbDJ18wDLhd8I1EL651Q4AmYONDMpcnch6m8iumtmItTRobXx1AZU5I
C1tWn3dfJ8kyBcmsBtH2GAflra5T6iIA34BY7RjDmX7DCOx83//dZ7seVUjg9T71
tPSIbwg3KOaEGvuoStGj0wV8jhAH/qpuuV49ayK4Ts4qAdfXU4ADEVGoR027MXLn
NTYRTJiPVZADp7x8VXqEaOCVMBiIQI4CdKR0QJ6sejXns/xh0zCkEkV0IoxHawmg
9g6N9AdCqIMNFmgEBJOICJkCEx++hMcjzLhoKzCpMb7mayr1pO++Tc41iVkAQTQb
uNTXPBoE+A+MGJMDpL2n84TqD9T6Pc/FiwgyHIukX6ls7/JJopbwQmQRr1PTAwca
9vU/M76MPATMyM6LDdMH9RWv2IM7K5IdPoZzrGfiIzmywoeukPM1NqFWcoA4EUVQ
0o2FzLmjf0Qp8VP/74IJgZL2y9CeyADwMZjG2L6n1mLwiXY84WcaMe2pei1602ww
FEe/vYgi9vFGvdWH5nooTMuUICkbLMQ55oqpWIGhAO8qlHb6st6OKEhT4rBwKb3r
OW08W+31GfNhyPhpbzZJJiqsWsX/aDtHnCJcniV2qqlPFBfRJEtPLHZtDagmSMTx
PZ6oochM2YIPJGyD2qmPkDX6m0vemqmk1UO49zW9WYYsT72d/8LO4NbySU58uB41
B5Jcx1eJYW1xYurlzHVDfERfgi+X1JkOgJ5MAeo9gVV7Auk9VmhmUOLV3MCO6CWd
1d1knoBI1FI0bT8VaIqsVRTmvebNuGy/G6ZOXcAzzJhqh/YhpWvMpOPXAXVhY5lD
Pw5/0s1hw0YgKsYPz3vDe9Sug12kpIeaeyvFoigzqHDybwemWZugG8RSBcfQ0iAa
Qc6LMSjy8i4DZTtXPAWwC9p92pv/dI0/E6pHrxFonfQcxJXjMg8/XzWjujHJn41e
rHuif7PWNR+YzhqGONACgM2tIXWQ/KuvG384C645X6e+fzuEjC2LdiSTv2BoixPI
jrxkmXO2KgxhHQ3Sa5JukBZ0zQE1DITQRrm6MrOrG538OczpYLu7tTf9vyz5xrMS
Kj3uEQCZYbHU8YZNpeltkgQPHWVZteVAyWqXyP/BG9rYyvpW3xBnlL1es1PhUfQE
7ONmmxWSbssQQUqLBkt7VXsGvtzv4pSXEbb6SzwUxT8IURQCo/1sXbVamEvdmMrV
CqxUiPwLmX+ayjm0Fbwgzin+i3HdvlUBVgqxybSLXyko9ZNCAa68qzwRXScFOTTi
JeAfaLW9XMcvnykj5BI761DfZbcOjqAPOB1QKHRX4bErl33us+xkZDOZOcFZBPbN
2iu9BYoavVZAXyc6xqxr1PaERTB1cLBJ5gc1036eGkqCj2XU27PzN64BwjOgrOAE
pPTjVynbLltrfEg7HwzmEIA13hm8opLKVUynOSN9T670hrq0d27wa5PKLBNqBkPa
ugrH/3sdQzpU9ArvkgMD3GFp7sU3sDAhrptB4Yt+Dhtf0rtns8FmV/OjLU1K456s
YbgQE8hFLtW1aMxk5/+LM+L6Fpuef1bGhh1n1kxfAB/3F203y16njtFODFkAnP19
SAvQFefqEJtF9dWZE7EPIioVtpGSpGuzJkZuk8wcgze8hKERg1kjEOOy3qsdXRAx
VjYrsmvGxbaJS3G3NcVK7TFEtFW7YeoFlA+9lIyvfQ5yQ1XmwJwAIC6tbi4CItF9
/H4vA4Av+b7mDuvR3I43ic1bGiHonCRpgJf2Dvhb6+PBiULlAW6huA0418q2tnBL
mbgxUkX5+3OdDDk8+HWp1GcuNAhktB7TJTwbugTY68Azwho1x7y2qyiL/Xf1tfqU
EgtuWnhaA3+RWdsUUYs0n+u0fVdaa2Vey8KQ4nHnONNgo47PCKMbswLTvn0Pq2J7
6G7JMiZ6p1q28U6scpKxJAOvmJKazsnbaEMkYA7AY785FCljuDj/3j+3NQiHXlDt
pYHPFFFY1IqaHZoF08bQhF0oc6VAn6GUTH+vYlNYYvCdEzyJmNH7b9xfHbInGZFc
IBRkLKnJ4yNmB614akvWvnhrqrc6xA/G9XosgFTmWE+mdZhfHB0dK3F70CXkMRpP
sk5+fnPpNV/l6jVAeR2z/vx1DypIOT0vcVQxMuJFXe/ekeAu/8TO8I5zTvlfGWrI
2r78Y4MYOqfhPEfJviSys4q1ujBcAFLX818rk/i35WGLDffXvqnAZ95r3UymDV3n
4cjDAc/YMR5A6CefpFPLwYbkSgoLxdccr7qEOuRHa9z5GrfjKLQ794tXMWovHs2L
HRN06YdAoskDJ4PdS9EceixV7xrLQO1Ns1qdMcAdYmr7roAWqPpOD5pz+PpXdbR9
rWM+Mv/dJ/VrSvUqa0vF2Hmo+XYcP1wm6q99xxjqcrTUc9SYOVEwWpHzrgGBF1wR
OMuTkua35wZHwYn87EpB4QtfLXT8UPGK96IzzrlFFeFS87nzNSTuaixIy0wW2OPY
HEO2kIOxLlyeN1OovcZCwlNhyrqlo8nLYVlX5UXtoSmBNCYpbrKVmGE5uHW0hhLz
KeDyey9hSfB4n7JutdP1REX47OrfCP8DCPNSY/c0XRek7F2Nfo7Io0rVGRsw0OYj
2wqonb00VRyHMazSPkBxTeaoD450uvNBAnSCtGuxc7KvH1HW0uY6rj6czZQPKuxr
h28jPPjFgRfHRfsaYaPBHlyAATd0tJaiZwTfilXyTgXc80xvpdwPCu/wrN5bDphW
nExfg6BU6G+Q6uv3z2SnrT0be8KNrLd/DrxTosLYV9ZVT941YNQPL//0Ewko2K3n
QC2Tfo2i5f85xrpH09OhHysuFWbwrE6A6PCaUMbJErkcis5Iiv57fAbiq0sG7bcX
aVAcuZrujO9O0H5lN9Gk20wtQv5fziIH+YeWDVZOfw3ymipZpXK4P3NZI2fOJ6yC
8hnATFlTal3IWN5RXu9AssdAdX4/4zKAI1E/diwSLxrwxLj9m9y8lJQ9HEgGGOEK
ruUjCiVKJZ12io2ggnieyNAv+a9fdUn8QdvLr9CqC0tq6EXIRju+uR7OpSRv+bDb
58+4qVoRgQecdR5Er2zn3a+we9vPvWM6fkTetF3QQ9ZjplD23BEW3sLGWayLk44E
ruxSvOtOd32v7pYATE7x9c71ZqhpY6kMIGKogZUDS7a+kjAffXXG0Eg7eTnWyHdo
PLGiBTTjhKI3UqV0+qP9AgTMWh6n54La4OGaxfRtyYf08Wc9cRW5q9z+56dONtRs
Pa2AJJ6qmfgbAh2d8exGabULrLIv4EPu1UqY8OAHRJH250xgZHNsDR5Rx1YD3J3J
sFz1PCaLGecAGtOjbmcHXcU+YEsFzkEi2WHYWFfCauJM6B5ztQ8SJjhgCSBgAlsU
1YAEHoDAfIpIhz/fwHPT7q1U/j8SmsoEB7FNl2utd7RrcQII5CwbvsCxf1JwdaLv
fo+kvzl8J13DTgGYlcVYAD1KMawwGvIDNnYHJWOFjQ2zE+YpSVczLWwSzh4isEMH
hfCkXMqijXVijmzqPGm9CpeBhTJcU6F11T+uKCIRPutCHYd50CaJBzP80zcTH4Tl
WJMeFwjOceFet042WZy7h+e8wu+3pZ8CNJF+pb1zoD2t8ooc0Twq9X/13Oo4yPgI
HvcC1f5DG5QixcV9rhKx1hyWmJzmDLVDVwgOaICEBrex0zvQ4Yq9rx+x9usDOViC
OhIWx2opUDXNzYZChFoKPpMiU88kkGBLglWfSI/SyAw5ABse6jF9mXcO+qAh+d8P
NT2wzRwSWCFKOG2A5w8RW8TBRXOkdjOqJppowytMnuo4jV2iFAmhLxn4biPseDwT
wQ4/7mx2It2bw+NR0Z8j+MGEZaNbHkgnxRcs8zr0Awld+X44wa+14vaUrc6vFTyJ
I0oJ6K5Bzuf9Znxv+7cPOFsH025+EP9vlSoaUKLBqSVhdNgJkad2lJBAHsO0ML4U
/axazGiKgwLBrLE9c2Tbp/BYwXkl2neBqjPs6h8xquj2QTv717/hWuWLYUFs4YGe
b410oTz9NKqMmniGj3DqAjQTps+MRFFcej2mlWyW8yjU0C8Gmqs+Jg1sSi5G+ESd
x0OTVUml/osL9pLuDD4s00TeQOFyMFmDjgo7kc3an1ks8Be4GcvfHXYmpjhBcuj4
6N6H9sKox4iEJYMgyp/fp1IQIwVh0SYVgqIzMvxDR0vxx0M2+efhfLpN84d5xn8q
x0HOjDaSCGBltyW0FZ4H5/evsuACORwjjQJzXNUR0qWO1dhBn1OM+yukpCafnql4
EJTuAja5jWwkB/HACWYFTgkFuXj/D3xtI2Y7SGoRUyiqNbOx9RcRFTW0B4FynZ81
3uh8RjfDgwPXgR3Fdu+wowujBI1jaLxx3uTYkz2y4nHtTmIGrt7jm4Cy7VBqotln
wXAmvM9O39MbQ/q5VFxWtARAghVg5DLxegdkOsPM1LttxGjxRzO+0KkSH7MDk5VZ
CIrJlo3ZZcYwDt3iWTSv2SFfE1sY2nKeQ4lVkwBGNyEOBv4fj8+kgEu61nwIhdRI
T95198FyEecWGTWsLuVQz60EPYREsqYOdDC/8w+JdBHamhDYvS8QCCJ9D2FwWOaD
4VCo22rcwbrzjsnmWCaLLaFpqvfAUkp8IO4yjq4h6P7Q3LcY0uukiOeAYiq+c65C
ovQqzPJ1J2v03hFwFZgoJYGkgkAytT1FVbVZW9Csd1AcNf2m47JcvdkF450mM1xo
GaCNv7kmNHcFDYZkR8YVexC3ZWaEgMHGDenerk3HPQy4akhxaik0yd4ElcA+dE9k
UeUIbYX8hu37cq7WitevVAIBKsgnvGfIU/PJ2MOXScz50OFxM9D3WkSH+BXsPKRI
/fPixuhgPRvA+QcxeVw45hjQedfbh8mwhGgvJm5YdMViygn3C4RnuXrYLSgLEQtA
IoaO6fpBqLaToTzyupqvXwr2hAuppQMEiDbBncurCPtsTsO8zfegucyrE/lvd8Z4
Mc5Q660PXUyd0tlWB6D6m9rhwaJgBVChrTG4DdR4QAmz3/R3ipAMnJ5Usmi0YzL1
g8BdqwhqFtq79PJyAOdtDB8spy/qzp0vHmznt5SphSVQFSYraPx6Oxl4dlelTaGv
M3aC/0c+hQIv/fWh+7XnlLfFMsvaYBmp5dPMOHOI3dy4k9nLL8VoUYCMsozVTE17
BEOyqHrLgsxQjWOA9dNPaBUb1BwE6O3guvqJlt0zILnYiTkecoU5WdTvVITMEG80
adcqK2Q0p3dYh3vC9BZPILCO9mwLkCfj0oxIf3eX+djYC5KPBNdGkA6dqTlP0D7U
nTaYcGzmIp43jpRtd5wzMncS5Zqt4TndOxjsIpo6obXhZEv2Zxteg1RV/6tlJZHT
maIr1tibOKLO0Z0uqFigD+IJZvPVAc5qhYU7YA9SB3RLQcadfZK6L6e86VLpYwVi
MyAHXxihkJo71Gogc4LIwUhi7E+7eubEG18qIpOysDdiHBApz0kTGoziFSzTT8Pl
5XaurO46I8ZFP2SvjB0U7bON/hCaj+twty6wFOA0+4z6p/2xunYJ0ieL7/834qSR
K2jRG41Qv74L7AIqgMJaATkrFFeK+9YRnF4xd2a5e1i4unMy0LRIilAsdN4N/6Ag
rfSYO8zrfXeCExxW+rj0PEOHbca6X9DTu+VvSw5sJxVJZILy4HxLugKwvS2vu/4Q
wFjv8ucdGx5Lxn3TSh5FeWkmWzK+Nx29TMedquI/EnX0DrOwdjMW7vcOiXIwSNed
NtEBilKntjB8vrz8G+r+ArZj581LXthMND26x5LzcqlljR6VNXcgi+gJrL0lHXjJ
EDPFLwgjI5UuXKyQqKI7oCPHfGYS9C3yPJRCoYsdM152PlEQ8NfuvGx0Tnx9uzz+
CFcZUKKIl5lJO8Ejk35Lq3oP1Cgywf7lpJRyMQuojoevsUa18zTpv5IuG83G5Rt7
4il1nHpqLWMIiNQiO7o8/yFtLAvsxbitLqpt43F7dll+PDjp5jaG68N2NFLGeiB9
tJ4oHm9sQK1V/C5M+HvS7mrrOBvFmpoJHHo+Lob0I+X8f39jCOIZClW50+wpku2l
Af8LNoYFRbiO9NAI1nKdcGTNdK4C0Ut4CevGElPMkWGNWndO8WVFSCMuuPd72bEY
KSBm+Hcpzu90HoRaxnxWaxpJKtDJ3QVkUiTMwN0K34NJVE0rPsp0xkOQWlrkg7tG
wyGvruAK/dLtU8vrVDFMzTn1LyUf5NVt0zkXgq00P6LSKbwUOKBj3fJ7QdvPqjul
8vWyTdZ6eXn1UoMYN9d/UklR62NcTEI/Q81xYMtMB5zQ8/RyqVH8pqd4rL/D9Jn2
rcXBmBtPfW1tcJDLodC9L8vZAXowNmPZ1a+yKydicCtPLm65FU8i2xCCRbbRqsbo
OtgSZGRlSmrcXdzu/qG00gisecTvzWt4FaqiJXHYUxiMtN4M3CYNcqkKZNH5qJPT
ydW8GnLZblwZ13lvPNeaPocwSSQruVoQq8YerCuTN2Soqk+6uXrrEktl15UmWTcA
CTosRtazPfj0bj7bf/1fw4btig+2h/k1X6JeJYseDHZi4JT2aYwxqIH8oAFV+6RB
sG1adiuL6M1f1UCkCkWf97bcP9QX5W0dfTVBvsJSdZbiwi/2j9smwwAOMKHfNyIx
7VaxJMmFtrx2lKNYBMYxQyVem8RTGRxsUpjxvPmp1kiYtf0DUEw0rriKBS+haUIo
nRzR98yPNGse6O28YvtOIvcjX4StnS+M1mwjVLk8Jj5E7kcHqOtu/xfU7zaHxViC
FRQTxJJv72jdFD4hCBu2kv9RLgxgL0NycMheD+2FyqN+JK+xTGxKk0Nv8TcvF+pK
6zx20pTHBnXwgNLBOXHvVVUwEzNiHVZyTKJ3AvCoNl6cEA8zusbiu7ICkBNkUhUa
SpF1PV9Px+k9gHFi1OrZac0IDAq/66cxw6CyD6mt0GctrBLahKKeSGCdkM4Vns/6
4Epr6MOkbc9k+8czMnTWikjdixZeEkiCIxKIp9Nh/ZuXpygTYiA3+GKDPuqqSnQ/
ONvwE+eUv/yQor/XysfaeSy7W+QKegEsc90IbtbUaE0krSIE/PDPt5CZdIKRBtIX
1gxOgrMFzAqbO0cZi2mGNHVnYAriPb3IqN+tLhmddtyAebT6T6ealbNMhES+WfRo
cvBgx1q6E8vMPjqnReJqZs6NfdNju0gUCQHayN+MwJkCox2sEywnwzI7NTVcPAmK
l3yX1S61y1SbOfsw6N8u+VHhic8+KJ9DmsNN8+P4zb4tpVIPkQj5z3+H3cqS8cy2
0O5/H1F5JDzYq+mgmdqhZIZ/lm+1aQUV/OlPzmd0g8pgYQ3Qsl2B3bPxmZpTOdCd
ROboTZZPZfBEQ2kkBBvaJ9VWzwAGHGCdzGuwENCKN7EMyQxO9vGFvgoZOuUqxTnO
gH+SBVi5yVuIqJbGevcQy5JagCaw4uKYcF2sCgVHF7nGeGxLGLDWp7rZ+K8YUtQk
cJec61E1nDL3pWopjjl49FExLtEbbB6KswzHf6NwvBWsFdwvzlxL5TITIIOR7lim
G2ztHJno+qhy/N82rT5FkJhYprRCvAbdqFxuWq2IUH67z25fuUF2gdsXohfH3s0X
+w7IEkyBh/nyWxpJTbv5h0jdm+y6ElcpFbhgiuOHwXQE04CL7zTBZbYgi2KlbCrO
m91VJiAkPW7QWrZxHQ6X86y8B6gLtrVmCy6ouoj3hhQMlvP3ZR+gCVtPdtkHiCg6
rd/iDYV9xicNGzbsRQssOk2odC4cRKepTZatTYEwOYsIe/0PgY6m/zWvSzl4SF+8
AX8eYKSGfZFdVhDAAVg5DiKa4iYYBdVWmtsrRxLwnKoW5/PyLmfMDI65Eb2pu6ew
LwS2/V93hTHtT+tlgnD2Qn4sjCb9bOyveooY8d0spCNalLnR7Npa2lxiYYpGaSXx
CvUpTOiRPxk0QoiAHytLHNJs8SwJLd6l8nHll94P7jH56BTX2bue+rfutrSlFwHu
H3ktKvJwJrNW1ikVQ/os3vAvFp/QRauNtG762CGa+NENLze0nXb2VIC8HKUQSTeb
KbPWpPkTtlsieLX7hCNPurExN/PCDNTleCkR/dxmu6RzDRjdivMTHYvMyuVUfn/i
lhvXHc1huPohUj61Uh57pj8s4UCqFaq+5IY+D1l4qa266zSkBLz/Q7NAtrIqaISt
9C+2mVw2i2QDeRgoNentmUXfCXePkA3iz0narGqe4Fm5Mn8V2FUb+p1/DZK+7FYW
m7Ibd+lUDe2uG+aq0mp3l7pa5ixeX7RUWffdYTuzpT0rLhBCUSptoDCX4FGdHTrh
I7b6+kc/+fOFXxjQDA6IDQrXmP6XiSAq4s8rtDpgvuh6TxbNYWNzWop+daIRb5a4
JuqijKdQIRJAAAPaKg+JF0ldJoJLmU05aJXl4PQPOM+3miZbbJjplNVP9NYKUVV3
ZawknNF8hPjoPn4+AsSdenMDYa68+MD+GhWVPpIUPPUDXS9Q9MMhWhg47ZnoGFKH
S6L7ZE17IfHe36SC2dGpWZBiO3kfN2QgFUPY3gAFAGwMTDbyIE409XVyyRd4hw9S
j0WyWkUBnq1xx92bM8XlH6uYEyigB6nYsyaUMt39MC95t8OdMdBFRSCPhFOMFP5f
D9pP+XnWwKt4FTZZDp3SAgupQg1c+enXmAVJNEsxf4yA8NIha7BVHq2kDQuYyFGB
Cu6D6VPvhwrp/XaOIuEHCCuS2fvGKux7GW3nPxiwr438O0FODXzyLtFNVBllbyOS
RsmQaqzGQ+J7ePie2U5h2z1wKs0pxC5r5AjJnPTMVzC+D9EnYwY6nntMGaGoDFR/
OGl9hgcZQJxmN6Ws3lO+nFsILtAz2PldjJ+Tx33MSKZYaC1wRDl+D+bc8z/3+Enf
EDn2R2jCA2WZf4gWqksFY3O4YGjb6gVYSBCVJiy7QB536RhwCHfN1gDBRWvbZA6o
Ssmn+14HfxYanYgHHJeZoYRDY576YNuhdFwFwjsJalN9BJvpkxyT5bpnd3OtMiyb
a8w1oQ/uGlRj2ZKKCHi5V2utk9UPBfR0qQSegAobNClLAxKppGEbld7Jt4zKXOEf
OBTk1h5N9FUZx8Gc/UZNUM5Y7kzSiQHPU4OFxJeMeB0alBFI4R11bBtDDUFgcVm3
ELOBs9CJC5pCm0ttGdqcCvkLAUO+5rdm7BrOZN1axo7z4WGnvEuql0F80yVg5rCN
APcdXvO2A602KJ30mSzPMcsU88KpArmzvPkUwFw9BAb21hA/Z/n9on4DvAgGov3O
mc18y9XTkWdAgGrnnX6JRlmNrMmkrCH8xbfb6KcpqpC4bZKx1O8iUj3cqx2LoCXz
gw/Mx935w8CodqgGIYHA/h+BgmbPfrnfGFt82O/vfRHeD7V4fE8DFNmqCpIKm4jA
TUXMRcqD/4TpP2hNfrPhgoPxCJZjC2Ia+W9z1uTJCCn1Ex0FaRnjh7qpG22/YtmL
yH9R9VxcGmb+d81yimbVr7WgRlZtnfltoi2LYoNnlbIRgZ9L4pThjtMDCgAbd//M
xY2w2F15aLw+BnArmxW0axY4VsmcETQ0IN21BX8CRb13plrEGy9gGvpUM8s6n3NN
aclU+Q5YmRshT8H8GTkxgQtLtlnkHPgQN33KXOa+5X3Xy9WRqBeSPG2nsq7zfXFt
25fgQHVYIEPAgBMk2Tx9gAe0kuUgaGMCYBoaFEvt8prM7VezUjEsG4SS1ydysNWS
wjFezUIYKB04Tcq+dozEY4px+2vH44TJ6qLC/3YaKM0EOG1HdLaD53RBnCHOJ9Lz
VrlH+/O2no9T7PKSFvNdaRjU8Kq++4FlyzSJWu01j31QK63lIwvHQ+BtnFKYPy74
z7wUHYBsM0Hzjxe6ZdtdCTH2f1DgeB8zp2m7eb9QVqbhOBPgM4O0X+N1WiIg/mJN
oDT0eovAFwOuuh4IIH/e8rYx/IhFBSkqTAhpNREB2rHnW+IpIVHHBvhaPs4v33Jn
w2rN/lxWCnqQfBXVsZTosYXcJqt2DPAmvRm+DGhUYCZJkvKluK745EVR8XCtRsCH
xypAdNYELBojg/bp2CRVDLq8BoSw3zng+1Sk8KJ+tYX8vLWW8tQG3qCH3OnwZuCb
zyOKkKj42n3nREXOZfn2537e5PQ4pzyA7XZoFvNHgl5Oot9K/4n6QGC6taZs1KpI
ew2kh1sybY/FQ9z83EyUZSSmFkTEvwu9hqX/2kKHL9lVakUuzJ/L31wm6MAQS0Jw
S5PdJDo40QS3BiTKGtn3gpoPu93953DfFcju3RgN7M548Ez3xZoWnXWEmZqthsCn
JawE0U2rIElBrsrF6toB2U9Ov3JBb1joP9R6cOzrYv8KFFHgBpF4RxmNxGXz4PEQ
ylpbY3eJx3YS9gWRn5gBQbzEXtskWDh1VoHa5JyE6lvSCTGIOCl5BXM8PvRAzYDj
57nVwwnrx05yobv1N2KfhxDA5R5zHG2pE5qFGIRqlsKzLHuEYowAFGl5y3kwTP7M
4H7/75VqlmMZ9Un2sn1A5L1Z07e2ku9vefqKbKLTRHVQkiYcGoU2PaOUcsXndcJ/
nQ/p45yPqmrj12NX4y8WBiKHhkJwnKGpCV5RQgrn0lB78kzgqdwZR/nt6eTTeIfg
0NBxnZt81WadE+WPG0buv3eMgcw3rVzw3kWA+iY/Jkmp2eWlnVFQuibzXTqVDdrV
ejO3Jq45fDfyiSYeXOUxBQ9To2yUZmZnyNIEgV6cmgAtYtOvGswRTAoy/84iVD42
217AOezvoTzYsn+pTCdPyVJoT7LebycEYA3mboUCuP117sCb3qjDf3pDFTrTUv6d
GaJjyWhYCFH5b3st3Xlu89cUbfsFTI475A/hZNj+Z2ZTZyflLfDdEkKWW4Znzpfs
L1C/NyCcsvAy2WItB2MNNd3B4M1kKA77V4VFxCI2U/UHMZQqlK25U+i1I/IgCVT7
tXjwpseMSdAukbBx9sF5WyEFM70kA/qKZ03Phu7JQEXLfEF/rdcp7RoaghJlNMwC
9D54nFnBcn0F+86Lknm8z/sWvXrqzvyDdc7QhdFBmMQ7T4Vze9evZ7mdDeAN0/5D
BCL2Os/cXB6rWxWGY1FAPanSRZcGcaK3zhpgFvi94F74FCLnazDtCdFvY/MdU5KZ
l/Hw2r6RcV0VESgre+Lw3s7MpJYGgU+76fy8IiuzXPcTENX6apG/rknNqQEKBQyG
+LIVqHVvCsv7E8o15gRGbtIEKiawrAnhgArn+wqPVGt4mWuT9wvuyJ32z+cxaqRG
uQCjeZunt9mfKEYFDTf4RMw6WNtrl45NZ5NnEpCK5pOPpqJ2y0H4s0zoruObsBrH
RISs2TK8atupEieHUZmqCs+unnXwqfE9efBAp7X5hPR01jyDMwsAyIx0uKk90R05
Kx6Pfg0eIG6S6alVSJE9WtLHxRgXSGvp3qfZL+CEJD7jjafJ+USIhT+shcEdMOgi
MXaQOdUchErRZdFbqOxnVCXNVw69l5NqcohlTkMKiKXvxxRvjJX6kNuqHN8e/jV9
Lf6k1QG9qKTIZWMm7YSjNNl6dZepO6oNkZQtwlgZh3ItylGOinNad9zu7sf7DLhh
qmL5YN7ue/k9dv7i4D9IUYgfiYS6enQQvAPjQ3LNQRiLumlyz69N2BYiYuYhY5WN
WkMRrNSa/mnI6rVsqUMeSNkViqmugAVrSofnHH3BkM0H0B0Q9NYs+eYjtom8vvPt
bsIxX2GaQB3ScQNzQKJ7oVXxkDfswBL2By+2IYplX64evvTxSGn0uovSR0taGADi
2p6JronRwNPv+RWvu2e0uEnwTgohR9sAikyKD9Yz/h+eyGZlregW3smuKUgi8jRY
Sb+5RxivrY1pPNrqZzVS3yu11CDsUNv3tY/tgbZdubtbT6Rp0Z+dJUF9hMyvlI3X
9w7I24nBRQDvBm7IM0bXG/NfciFGxWdaleJmONT+gP/Du25dw4mRPKzW2M8LCk5L
CPNE31bxPMaXddgi2D5iY+34t96IlVPDVbUYb1ZS++NyEjqm6IAzm0fJmINW6HvT
DpoWCbuKzKTixmCdhui6/tP1sQguMZITYfqKzKP8YAheyPFGvNMC3Q4p8tr7I7+R
nqwlI19B0cmD6XVU/PjRj7kwE3VqEJosmBzu7SB4ZeEaiV5BxlLCkFFdFEOaZkWZ
bNhJ1oZhjT5pcEwusQ90IpbAd1priuybEPKTb+2xC96pSzC2iyYelNrXhLA1Pn1m
WRRoKIvctAwYBQBiWLo0H2yvjz6mXJm+uEQ3pObBmpyDQrRsdfnLDr0S0DR/rggh
Wl8s1qfv1o1bQ+nNb37j8FZnt05eGxaxfpst6SjRClyC/JVLTJ2X9B47Dk+sl9gc
Ndg5CFH3jAeRuVsmt/yTNFJNWER4cF2/S99ReRgWtwP7dzqoSOrBxZnxwGTQLSoc
YUjFU2KYlp8s1jgv3legmoBE9/T5rLVy54PKfPT/z70r+9G1v2qI0um0Hn5JBR4H
ytM/ZI17wACPCSlCL20UK8Ia8a8HAUs7tEUMf2IMOmR5IS62mZd6fh/B/Ly8g0bx
q+sGhRBT29W2D5/Cx6QSMk7mVqNCDIZ7pgHZvAHKsgU8d1mpiRDHMbPypvjO7fGk
m1CcFHW4Z9hYRajFswyjf9Ifc41dA4T47A8zf4H3Uf1fLvHVEnJGbiaGVg0BrHLn
DEL6u3Thd+0OHcro6of+K7hfpkU20NdLga7MaZBSdf24nLLGrvkhK/v8yoURxWmN
Xso2B3kjrxdrowzwtC98zF8yE1nW5LbeO8jeEBs93spWufS9tCC+9KNkDS8a40n2
X9HBfYPIWwZxlvOWYQE0I6LIBkRwb9frbnuqLTM8zMpy2neUCSwaRFwkWKZ70CgU
QFGDIharFARTuscaFSVd9n4bgrplxoQ271ybQ/kbW/imZ4loFIZjp5yTdfObZ/zr
Xm4F6J5BQE1+Qv2MwJ0CYOCGLNkNVVVGTtfVzsFXdOaCyRoyScJpmNT7t5ElEZ4H
IDwb04YPvV9/URT9Gsx3N6luAxXn9TTcH6tabX0FSw+WXbwZPoxx5XFjoEnlwese
bhsqtxhJZYaFDmrT6Q5IfckCKEm7aRUtPoNYjirXEdOtI0R5l4EWcoEemTg3BlSf
Xq8qsuai03FPOBQv9WBoesI/717N8tNOQgguNiGJR7/lkOubo0C1h3/SDjg1q8Yf
weWnMTmeTethlS4JPi3G6evEsmDHMIVASisz9wXU08i9LcHYxRh81BUP0s+DsKHv
qK6Y+M+r/7mXnxrZWEbWgutsLd+wL1/9VD2ba34i4PvUiPYZxvQX+OlecJbX3F5E
LCcTV26wnORhlrAtgRoB7LGRzo1I4y2haUS2kQzwrK30tsrTkOCXRCh77GfpL/12
feJH7WRlUYffOBOKgyowCqJ5c0fVZioBi2Rtt/XErQZDUOfqGg16a9/2owNy/fwe
ociJ+i2DH7L0iBZrFh/oAYrePuH/V8utHJNNEUdp3KBee9dQmqbdri4bK1SKRfoW
QBrmSLoO0cyjTBqkVIDeYwelEI/i6jT8cHX87OZMFxuc+kff9CJikl00vCwWd5aq
TtzkGpfR6UEe0SxuEmPWxAP75+mf1XejqHxGHedFtXDVyqfETYjzHTX/J0Y00+n9
AFcvOk5W9feJyoi66r8FySuTov1fqNhme0+5diGA9lqHHvZYFhECcSl2IXJUOZPF
5JeL7S643XBbw7rsah86x0cnUP+sUrsx733gFXeusVDwZuKL+tLRjsNIGyBQ2tAV
lcV8Zl0Nf+TpT590Ytzc5lFf/Q+YzuRGAZVsCc2GXuZ0M4+CAZLrFlXUJDTNe3mz
xcqwEtjvTeXt+p76qIfg0P5OMxU6c8boWMf9hpvXvQkQFVq5jjXgfnJwepeyeUCz
L0rcl8Hc4oxAEankV0V8NR2zCC6rE9UWGRxXLlMKwfDI4IaqxB2BEdMI8TzJEGTx
w9mm+S9WfZEckf/ttWvxuIh1Tslnv1OkkZEEnmy6gmu1reGN7NMV8lG4X7RYekhp
jk6AtQzPMia8qRLKQW10zW486OhD7OOoVIFA2BKSU6rR19+yKCgmqWfXExm2g9G/
MMhTCj+rhTcrm2YmdhIrTZe0xkIoFiGCDLZMBlSzSZfiQyNiUgKZ9uOkCVO6Qpcf
FzjaTR/oXp/8iSO7S9MNs2VWVgV52XXMbJCATfa7IBZkUVYg/4+LKYsODHiwWQFF
DRrkD4pHZ0iJuaUlkmqVUPWDzWR1G2BbsFgQvKFIdVGxbBeU5GRBHNHS1QEBGzVP
rSHpIVczPQ1NFAJAXBMdSbbQ9f0NRS2poEfRXo4LAMo9mUwQB7YTC2bfKemqqhoa
cyXsmiAuLRIoouLFv5JHRblO6sfOB4LAVBuN3mJbbZGq1msFDx2QA/j3UrmVgfTi
kExS41WklERsbT51zr9uVRPvzp2c59NOi0y1WGbk7jvR9qjMmm3lDWVSeUMgLiOQ
XAqmMbdFSiptLSmMI7UvYk46jOws0IAL6gIZgmHDALSyp3y3L0eu1nKvV5XTtr+/
8MVzvPi8bcMW1JjortPgnI9zXsirvFkqN1FScgVl+QnovfJWG754qdExd++zPhZA
oCpm9bHCZcmYvhQ0un/V4ekMRifeoWwdlD5qTKElttvw4VCaMtkyi+i26lZwu94i
2EMEJQz21Pymp5RUwVJEsGIP/Hi+dn2W42KAxM+87WqufhHQqrE5AamQp4Pj5WvU
/Vu0Tuj5wNSjkVWD1GcWURaurbkYeaaPODcyb6UMA3oqAnnFFGNGnJKwZ/ZZH0sX
fq5HuZkJqtUA81DBj9gwc/iWFbb/XuZiJn6K8Z3gt5cJZqe37nTaDjlZczyQau3Z
sF7hXFZbn2PhhrqXyVSjuSVkxFGNzKuFdGzLL25K02/1D07it3BZepOwTJFPkQTu
RemabZV0rZTFU1tBykU0+i+svNSqkoNUDDIeQ+DLz/C3QZ38yzLg8rDN6gjAumxH
IYKlu4kFkrdgBAY/vq5DYS5wOp++kAzuiLMRgf0SUBe2lo1Elq4fsyPfDN2W0qKL
RFwpc8p1aJ5ufLtZo9qECNpYPmy5VKpSzb2sDarcx8NRNuMT/K/AWWEmYw2TLIjf
hOUI8uxDNCbRrFdiWSKHCrhYaKWNDz8W8U8Zlpdl6L/JpEyYodEqBpGQaAzblvgX
pAp4fGiPe3dH+/3Nt3kYKUgnyeSGlBc9Z2S1pzUkSZvMUh8LZB7jS9HY5ircrqOp
Pr8m0p9SLmQ1jfoHMri8b9JZJq+fi+n7zKdCfxtuhxTzJaMaYMeCVSUkirEwDk4N
MCArYqxpBcOBNk7VXDesXTCfXz7aBvrq25QVlaJhC18LIoO4ExgNlnT7NjMtpXqe
l7pjTp3DKxcXBJOnxZXEJ2eJayZoyofCYiAQjVJ6J1xMTRacd2B52Oz/NsUnuapE
s5nCgW4B1N4maaLqaOU1R427HGIJ9wJbmteCSWHQxuRcb2kGpT1n5pqJ780HmNnN
n0sFlR+80cM8NLYKT0j6GsrE9PdGC1Xaz6g+Gano21klH4f4KDhe2EV0equqMTW2
dZ+tunkj7d47NyuBL9WDhLrQhzBLktgPaUdaCFkQ9Lnp3oMS4SPJdGzlwDCHBlux
pFteu3xNcUmkj4VsIpa1tjeDqXXTkTnA69XdCCzUXV35UQMdi95didYMenDzmEU0
SjFOE69DkwsP+8e+8GDEQYimIQH4Brq9qIbArkN+eXWEvWGXViBMMLCTCfEcT+mW
DxrjrjUzVCNKXe5dZ5fgU86CckAviFiv+8Zx+vdLzvC5Nz1r9aZO6kOyuUfek81y
WoDZb6S0j2JMy8ReH6pPb0nS49GwJ3vtadTtJFxw4Vun9J7dmhv7E5z+Z83hVWOt
eHA7KIhRY0NaXsyvigkMdiHPHA5oj2CIcH6XFAdJB+5DMh1oBRnF59mQD7nszU+X
Ieg7causiAxmwGBAY6UaJI2Q5Jr1uBs/+6iwWKH89BqpSjhkZHS/K5rbPbMobCCI
SIzDXYtpNv54WJrwcZvAodSRcljKSmnDUI77KUO0ms2IwXdC7gq9WXotg0UsPzUp
L/jrQPZiswRe++WpcVRdaLzyvvNmAPJe15/E3UnOfFJ8WwJO0FtJGOOaKMci8KVl
jooKQXMzv+Amm7FpnnzzTO/6wGt+9tW71+FXb507v3FwR+yBIbfjLQfx0w3B82Of
MNEQafNc0UIGJCsU5Szqejn5Hp/zLI/j1tqt2haKDErgdYUSMgXS8NQkFReDhWl4
j+xisq8bg88sTB267KzMxTp+US4yiztZFlWGTjRAgMfrIL8J+evMerAu1jpeIqnn
WHZgcnLPx4rgOJEajDQM4jgwWhz8u826/fQqEoD60zFh/lXUapCV2yIeqFmSoIxt
v85X8mKtzDDawZIAnz+EBEGToMIkF+qVPj80NhfVRG1Lbw4cO56YDHQiMvpZ09P8
KWrL1FKG8ElClMlCnHHCDqnBfS6KkIKMIUvzBGN0JfB2imTm4l5T/R5wXKkVhLeq
4tiGJYCLHyG/oui2Pf15/UfEPxFI9+iTVKfXWHeSx4YUfkSkThLO80QAfkUVmGRj
mx2Xv7tzn1OKwlW6SlQKTJug+bGKogoBeC6xmTJRhrWgcC9uy3yGanYbjXudzeuW
+nJttzmCJySAMvoFro9tyzS5fDS2eh9fn9M88NtERAapmLyXRDsqApGjW96OwR/q
pgEmlq2ptnJSyMIWbnL6ilVaQ2a7J0c/LiPp527Y6REirJ56ZJDsDid3pNGfx5So
jUxFbik5Vj/Lqmk8OIEFagKmI54RQrCkwC3K11yDKxrl1xiAD4f4btQhJZPLO0af
LdXKX7vifTZCJlKNMl3NYAJZyTVIP2CYZucsKdTm7B4EoJ+MkbP0damOm19aLyyG
yMOs5TO3yAL/FrcuBgAP1If4HhtYUt9jNJCvOojaxM3ZtDvTv1/ZcQ4RA3X5B6wi
gxNOzhvdfvydGMGCuEU6ot816YZAndw3tT9BzUUCEu0WRhU28Zb3GD1625sSRcVN
1Ky2FoNOPolzRaksdX+ju81oOfsD87VSOlzLT9HkjSR6DhCnhCJL9POu3OOOU/wV
9EZQHR0UsqsDhHT/c372xc+Sc7RZn59zEwCB5N2qFLHYstIU2MA8S0axhdQF6ca9
Yifeu/Xyz6y2UyFlMwquYjgY3jHNjGn6+ZhFKSG29i1N7xQDu3J9nTIfHuyATLD0
by17ypQ0nMm/3s7BDPd41SQ87rVExa9HLorUiuhZYWE0D3Kn0kGQgUrPr4N5H7jD
Dz7x9APnSGH2ETuAmGN8QCQP4obEE4EbodD7eH1TSlNQ3koLngN/x4E2KdVwnZdM
atc2mG/c2/Gysap6BXHoMZkXjHr6AOxkgT+PhGd6dCr9x9VYOSPfAMy3gwxcOjwu
+eWMMQM4jk6i99Jr2n6xVXtYvTAOtcPIauj0du5/mn/NaEJ9r4lpptNOxEVRpGIJ
A2lAEkKuy+73k9yLSZ8+xaYP4cLmEHcb64g/T3IZgI6wa5oo9FvMOkBTcxGcKMIJ
/s4WE8vQQ7P2iCmjI3hczQfLA3/be7/WfQvcrL/auiU/PlCveBOjuLNuyRddXRWj
klTly7RPCTou1ZvAvp5oUASScTb6EXNTmtHceGZwU9odK+7opVr2Wvsq7uyTvhts
vXb+XcrUHzLIY8zag5iFZ5T2Jqd41dWSKPjGWJRJ6XLFaA3UYk672kyWIH8k2QFh
O740lNLm1TathD6x/HFEGZostIo6u9UF0mc/H7ZGEMRQL04nsvsSevfDO69g9Xmh
7btOcQizY+mQQlQz0MMV01lf1huAHW0aML4MeXzly49fGymALgbf0luKDFb3GP1s
ptMLVjegeEm6WN4OASUH665wO+M6j0NQNOSv4iriOFsUbFFChNyLSWTwWez7dy4J
eY8Vs5iAtOn7l+oeN10TcqKs/5d560OKrh3AdPGcQoPY0kBEwUjoRyL+B6ss8UhG
MKjvzl9ytvoiwDIvZL7TSpXaIPSHx47ccy9AoiXkuPhlzMFy9v1MvNAh+8FjKXla
r1y5YQbHfE/MDIEncSf54YwvaYj8s12PxneD/fynhk3BxJgOIi8sWM0+yyCaSBYN
oNmIpVj0YNV+jqp0EoPjhiZ8QJiYJLBVYIYp4VbKjpqjX0G95LQbmXrtXe9JQsM9
Dov79lDSu0he8HRk19n2d/zL0GLEw+JGivwCZ7bt4i/npxKTLjxZgUk5kuv+7GWH
C+DrGzSGaaD7wqo1pqx6/FOo9FJcUIpNYs15LLB3QS/tHeDvkYKyB43KWCUNUnLx
RpvTkHvEF8A8Sw8M//i8s5nYHw2XyZ8qa7W1UC+SM3Drtg75pVcqQMLy8osdK54y
iHcwDVwfq2CNu3Lb7W8BC++5Tvow77V25hk4SAtqlrgBAFb7IPnn0TzNYps5XmyD
4lWjN2KoGeDYYUe7tJf0H0oyS11aBPNz+ElDZnAw29uOfClPYhX+UbbQiix3hI1a
aawLMkrQQ14Vcggoqx/r3sJphzIq6DOFPhft+Kls8nn1sh0fAgk39HbpER1K5Atm
dGsu3+rhi/T7wscHvn9bJQ97+XcaZCye5DclvPpv3jIiKp5D2jtzrO5vvA2EhyCY
T1L+hFm5Z27X5GQNCL2wkn1sIWHI6mYBJde+yHBiyfN+2UHlo3Ah4gufSskAAUzH
U4eUDJFsFQcdeJY+DWUexCf0f0zxmykMxt2d3F+/cO7l5s5QbKJdSvaa8dQFvVGu
LH9UGWYz2QvplG3gir4Y8GhdnBnI79sQahAoOdyTT5joBJQdfv93Wl5C9TaZg5TI
8IfAwZwKGAGw2ByufyT+e4uv8pIn9r+/yA32Dg0UrKpUv3S+hccFeD/w3AkmsqnF
dgeHVPLkaO+q4sJdwqvdeKloiJXziXQlEaKjz9ooYpI9yNM9QxQ02MiR4DG1RVHl
z5/i92uqy2EPR8OQDl4HrA++Wgiu3t792Y55m/C9LBJAogHflhRz0oywLKJEAuLC
luZBr00nz/eGY0eVMFZ6RfWl0gB8FMHyuKp3uZjZoXJJXzDcRDCxeXdllcGkgZYK
64YQy8TKNR2cuVxivb3N7j3uhVlLmU2fboH3I1WR+Z+Cb0CnZyBjNc7h7T63YluH
eLXs896doVL18kSOI0f03yDdb7J83mL412xYkFCDDdrVE8HrIWboWYTcuKZa5q+h
4mV19bpsCnE1Tkm8t44AdBmY+wt4TP1W7uVHiZhO4Kv3RJcOOwHUTE0RzPExC9aI
DyYXu2L1mOzrpi/S07tZHsk58x1acTpkwVeuMwgOO/d/1Rvbe55v35IgNO88b3Id
J8GH14SpXriWp3HY9/8Htt8KRg4nfPdYs+tcBJ+nm3toNnjQCg12+LrW+TIz4hB1
sQOY3/i6LnuvIpEiRdJ2OiF2E5rZfjaBis2w42SKBwYqd0N2YOkKfuJCMnMJm6dx
tlnfbMFcjDHvEV3OlAi59SeYyB+42vOAIO0ffsl//+ykmjCemHeDNijntHa66hb2
0QFaLVAvtYfG6UfZTqMORq8s5Jge7G7EuWR0NRHwU3XURGcEPhwT31w0vjxdXR4I
t7R1TgSpOQ59RqKGCj52IEYopQJvJTkkBBPF0Fp8o7F1DwowWfkzJgMb6ND7abXo
YB9197sse9Bn/hNQY2NhklhNrq4AbsepBs3bb1SCg6XQ/071byAB5KA4ix2KaGr/
ev0gAXRpF4k0jV4eFhpEtI/krbkrYg2q3/hGb4mMJCae9hIWEJ3d+hZbRl3vUZ3/
BJLin3xVYsvuNjpQK8NWDEKzi8E3YEfurh1kQuk+LWPq79ZpbSl3yXb+vVIFGQyE
ypmw86IlKrIfurg9v/7DsyQxQKiS4J9wprWYnbGNQOLgt6ieyapJhNpRT0Z6Eju2
umSFuiIJ9ztaGzovhj0SML+6AE67LS2kGbTXdqgqZfPNCw+UciQzr8I4UisuOpke
Z6BcZb6yx12g/Xvr3akZE5ROXKziARq5fpsTXFeUfRWcv6Yls8n4h0g0QMQppcto
GIgXmCMQugWjOwwRqMh8IwCou0jfGHV5Y0qqQkF3DdUUMA7twXvHyYLH0AKQily0
qIEDiATTPMtC2nq/0vaGA9BmizIVxDAFuXolYRjkC+AH1QqT9WWAvTgZI9FRQ2Me
5J432wBzeTZ8rMJDjSrsFgGrVeq7c9bsFcTh6TfV3ya1vQSyQK9e7StdnMX8ZEQM
sdxZFsBGJSKSvhJ3dzO0m1jgJLGlic7FdJcfgJcmbgK25qziQws/q6cE5ufpXEdb
MKphQV3s5A1puuzcxMF/0im2hiLvJqgq4IluscOuZoWSQkUgD43v5hPwmM7mbYX0
1hv1ABSQSBS+EbeM8v3cr6JTHgvxvX8gMhBU1FcpvgO+DvAxQ6WkvK6gBFouee6n
BkFSlh9ZC8K4pdmC3kppfFEukxK0504piP+BQ2DSajjwx7wChPDHMh6bI/REe7EQ
U8D5bo1t3YrCVBMT9M+I+RWidd68CswoZUGjoHihrGTUJZLg01pkWG3MIORNb89G
hLWMY2hTbi5ZqAksyjrBDx0likKBFAa3oeXCfTVTcmymQe1+fBXiKiPr9UQIXcx6
HWB6BipKxb6Nr8ypKLGk1S9Rg3hGw9zBq3UV/AT75E5AaKWBLGX4aVZwLsrlBfyb
mV6mr2LFqqNbBP2gGdFFSNO+dUjbdOWmizs1eADqefhIq59SvvDdMcdpBm5Yb24d
VQEcm/4ENJFF6T6WnnqcO0p59IQXBxIjFioQPnhVxhTqo8QHhYaQvbMa64CKORQ9
zPh6BlBJ7dBJTVuYBbOT+cSKxR3lhh/he6OTs4kUypgHr6mv6pjtlPm7jisD6CUc
a2hdKq7EaJLk3cNaPSJu/KQbAaUqO5ResMLESZ8Tn7zu0OzS6eKtI7RelyNIg7wT
8wupWctt7m8JmGC41GZKTiCJFVCQjQP2HkyhmZlrg0hfsKooTqAQB10MCWSoLOAO
BVdzDFrA/UURpqgU0+3weMyxtRqybASjTmfjwJtU+zq9jcRHvrbpUe2Gjo5L4VNH
G8zzUoBWphCafW6Do21oszfRe+YhD9rpfBEHCYP/qah6igvl156Dp846GYl39v5N
00zjTo1tIvqaeqwNoi/e4Ya0qm6VIlmTgo3QiqE3IKaHDS28ZNYtjciPNqEkywji
zalm9NI1QPhYaUBRQ3pPT4AAUCazgZ0R8LcSQVB5r/um33CN9fi3Y2kJaqgRdVa7
PjMDrgoUJRpYkq79gfn4HFICEbKFjMGuV76aDSMT4TIvUKToBWGrfusGYL6HCa8H
FOfq1DgDGlCJHsVVxeb8DSz3gctb9i1XWvYuXPG+2J7VrUGJm3v4kyrs9mm/vQQ4
kKjVOXYp7OJBiR4sBE8j/baArOhBaziWfWYkvMOYjxrxR521+Kp5AsFvEuI+WLZ9
LeChd82KVFi/hISUM/LHkRYMbDHmxRQwU7XAo6F6b6tgt3hw16/SCABOCEKxfxja
HFjGOje4CWZ8A3h0iF0CjOyGZk1Gls3VRHsgBAe577TRnAQaF4LleZ9OFpXFAsEE
aeIqwGqeHXUENusvduXJvWfW4LvqAUcnisKy975FAR85xeGfyKbNc0WxeZJEV0XL
VKHUPOzOLDpfsQJRosG27vZuhvGAV24NjOs1DNbGnvggr5ktOvoZ33Zns+hUigSh
qzV/H8MGLUDq5Vmr6sIIYCZY7U8QXC/9Y3DRDl4u8X2LV1oXV1pjF8s0cboYokOu
2OI5MQTCan5bplZyNBQIxrDjOX9R2Co/FdK+tH0647hmHRrjMvE0sVFd/e4oWesx
MHeEIERnKeXpN3xKWoWiHjlfjXpEj1pLQn6SC6zrrYslpfICFEtJn1W3OYNjiIYa
rHd84xEM0xZX21VUgRbV10qSJi8uzd7u3gkzkRpRjDYBErjbCLTQxz5gEREJh4lA
i02km+kCeedOmzW4maH6WHTqruZg/98ttny71MiUp7s54nphZPfD7DquAvf6+8+P
B2aogJMLHCDfMOlm+YJeKE+3akCvN1qUnZqbvFkiWLyVoYOA6irKCEHxz4x/CnUi
i+BAGuLHfwM82MwrKTyNs0IV/Qwp+uOF6zG0KhBUE22AcBr51o3go1sadLQC0lt4
4TWEM7ysCUQOlp0nQYivNaJFJ/kCajWyzUyfttFiJRxOABdQsIEDx7X/OPeJofQ3
N2zup3+74OV3A9NjuIfbHtXxMOqQoSRS3zDGgj/6GItOdf/RZ8hPnD39tmkX+6ty
07mCEThBDTLElGehxDU4NVvcSP0e2XStu+a/uVwhsQyC8SLc8pHI+jbfnp799KWq
2jzV7r6fQru1qFD8/RjK0+P9TxhD0u6SduR+cnl5tTMstcUjd86aRc6N8CkP3Kgt
ZrUpDnW/Qdu8Z8eHN6NX34SYH0gQrTyKrIQeKewsPlQxq8D2TdENOMI6U1TuS76I
mNGviRv/FaBZR25yPFHy4weHm/MHkbOM+xiUnpa465oNxcc/w469MAlyfg2wpInU
pAClRf1zKqUt0iLHa/mG1Kzy3CSFwtbwAYQZLTz5NdDOTJvX4DONQ8wn6B/w0FPG
oYHIkmQHxjv2bCSeO3FnflrCgJs7G5OppdnfMHJwrRlU/XF3A9+xc8XozF/QjQug
KK0RAzIJ984xGAtCr9y9nIIr5QHrYXNCvajXvHvp3ilPNXKm1eMWMezHa1LrCcUL
mDn7Z1z1HVPURcohPeGZO6/PTjDc0Ih7J6tnjZgO5/14oLYvLFdM0PDf5FY8iRKn
wgzFB8HYG9LANEhHkkamAzIjgTD4WzRdTUvs9M33bSZhY5Wpj/F5yyd3Ox9NdX8T
3gMkFTaBXN1LL+P/ndbzs8X1P8xv5640iSDFhtEzUuoHkaMhPM10pptk4PFCwMzc
2tsnWKREFhERH8Sv0plolmSc+0EcQ+fIzspB8Cabr3nxG3Io5nwvnr3Mw15FlVt4
Qmf3gepv1/w6YYOzPZ1ziUmFwLwK9vmMjtAKeK44sXQNMqmxYyPBEFouLikJ1guE
CF6xDMF6plOg9B4ZjQifJRcmwcNpIGbLix0jHhxW2sa7HmJ/7TkXGSogMxKFJSTb
8F+XvWXSdYanJ7tGWwynExxmK+N27gWjJLqgSfHMhX9dmyRiuzt9RdmGmK6BMFkb
DRhYqnFMe4L/1Sd/53yaqWlLRF2Hl5PO9XTer7d0mjvoTs/6a9ej1v65Tj0juT2B
1EJffwvTibfM2HfOiMcv82GBbnG9oOiTr7JljXaknuOEagnw2Z2EXIhAD4hYXHX/
zleVpC+KUKv0B1oLbshkE/sCnkER/xOj9yYyK3XW5xvZWHsqp4/AHrUWRPtJXBAg
NsAaTXX/9sXmTkZ/vYEZJFEYqM1AaLlA9U0ZszN9/aqtwjcVTfG0ZgljwRLqEz7e
WglZx47/P/Cw2LlhuIDPCxIeshZzYuy/sKNhqRFUpok8CeZBe9DEPoVFcvV7/Xdp
12arZNFko0ICCfePcFAIJPmMprHlxibSt91I6UmNEcmXbUwNKdmCMhZUf40v7DSc
mmM5cTNvUnyssOIY5271dOGKKn7eSciv/lWbMe4shFihBssKV9/Hu2yJNPTSAk/y
C9FfNxQoX82kqa+dtvpCOVAoYXUuQvjfPJSf7ZBFiecQCFFQDITZlKaVab4m2PvE
ft5frqN64zeN30UG59kSgCg8c7rvwIhSrKkkSbUoNV0mbHJ+f+qWVQdPe31H/yBK
X5uy/5vBV/lLqNN5LGGAfSCXTOiNc2czA7I2hT2bvuNnlYIjI2r3fqXkDRJy5hNJ
RwXzmWVXGpnZbiSY6cjbIqxUz2AsANFSkyyZZEVyNslL65ccVOHaJyA6ayVayGzu
0VVlG8mX4fq15E+9vct7LWtJWgh0kOdBklSRRrzc0uHHuodUzWma6Hb9+eoG5Za6
v+svpL9ecUhSXI8oTCOwXfuwD+nT8OS+/OWP1Pnb9NTzojCR3WAadSCK5DP88TZ7
JFkIMY4qOuj2t9/HWJoTTd1MzUEDHsKSpfYQSuxLt05qrSEl/umKHQAKxEzpjA7j
SRYu1U2BXbdWSUwysgjx6ngKURnEzDS53US28TVCrTlZFhXPHWNVcP0+U89QZ1a2
cq2HMS9UPAi89vbGf0TZm0dpdKZTb23m+NOGOWfk8Dbvme+lYMRCmtTtQ5Kz5BUb
JdiQD2ipygafuS975KTKRECrCjFGRpLQUPEUz+sCvYAtCzRGw+NXX6WnkMjpLYCF
CVodg3QTsKVLtkEWZ5vgYlqoofESse2cTddQFYWxVoyPtytTWuo51qCzDxlvuNgr
c303xsrVqmeNMelWBjmFLWplhnvMf7YPpVVH08bfyjOKAPwm/1FNsD+YGe3x/qHh
TDugjn0K9jx88Zj7VIRjB0mXU0+3VmLuoxph4HYKAFe89hyHsVjvfn5AP3CM3StR
dUFoLxvbdYgQfhOKAPWFkKfQOPAojewtjJI/Jkqdih+NWaTCBDWqCTGf4hcA+4//
Bc5jEB5Eye6hVGFSEYHulWLjcHB+vBv5v4Exd1wYWLJhM/Wq5UiITJBq/8OiBELq
PfswE9kyVBPBZ7JnypdjhDykshkFp+03Lum4kKetnAvodxJ3Rv/A+mrlRtnkKm9Q
jOIh2qcGbIrxM0+0Ejbc+Oqw5c6DH/nU4mH0caNZO00jTUtJgo2O/mJhc3dYLymg
GLZJ5N8/mwhyFIJZrMFD+u0T3I2mplx87zz8YSygol4tDtiRXk5WLWsPmCNdw34g
C1uIF9cJ94NakEGJDV7nm0b2bEVO5zbUCHaQ1QcXf5xF2HO6rzXjfbdmRuyLaAn8
mh7cxeTHHKR5h5UfuCuPRdkWIjlyB9jLe8/9utvIV4b7PqtGVcRBOX0IBhI/D9br
2g9d2NqA6RlnccY1pTRiuKv/h45jAfLE0tfH3R4vkgoAgv1vT6xZEA4AGWLEwUHL
/WBFF4ShDYd8gNyxddefDtgnto2bBEOflx/A26OIXsLAynwFCl0XJNpnXUMbdj5H
zv5+q4uziL9PhfUrUqQz9gc9RX0UtDrkeLHl0UcffWPuNPk8H+sDZtSWGFwwhhpd
gdcCzHcbZN8Ml61ywV62ZwwcEvSEB+OIisviAkBekny1WAT0Nx2iP3Mm+Ne2LRfh
9R1maSiKuZt15/NjAH9FRTfYJlya7dRhZ4CpZOliAGKq7+5kWMovNkT1TXtgMhnJ
WhR/f3Tn8tsgfk0eMu59D9VZVwDuhl7/caZgLAWkKZVbQhY02rjU9ZZtTUgrSsC/
M1Z348A9K7pp9z+RcQFNT6lrBXgJqnV3on2TEAX77oP26EO1JiOlPzZTWwEpIL6P
MQ3MP91v1uizEmTjKN7Lk8YPI2JPw3BrEApBGuDgAuoZ6UFsMyIjhSdXu7KmqXqv
BjvMtiRC2nRpScIn6Bes5QigYRiZgMa2ZJPIJP0W1fN5vfmJELjbA8osuy6UtWub
OkZP5ioG5hyrqRu+MnBQvD3Xy8a/vvze/OoyTG3pxmEUT+T2Je/ac3E7ip25NG5E
eXY+hFuyS/CZtx8efNG48SVIREYo605Woh0xf/teFMaYxsjHyO8U9IK1shZkZPTQ
i+CRhCclEsDRA2LUInuEgp+5UReu5c613izvpAVU8h9f84l2saDmD/XwlZtzgM8e
Z5uGW/NdOtAM+YlmpqnLWamlCnIsEFgmagaNhfU82bji/1VVXvBmnGK31D3rBcfV
xoCDy6/S79rg78FQdDthEK6Bqsn/vaZtvpgu9fLg0G9G3HzQfSln4MG+IR3vYrGF
YE3BI4ZsCd/AbXWfwzdkcTWlHrm6Is0o+Qqo8CGcxdbtA6LWwUOn+jjQl1DN3EH8
DjU+t7jPN+r4fucJ/pJgKP/4PAzzEYCpIMQL2N9r6fcA7MeeTHV7azsMIwDLgRYw
f3y5AH+SLEWAIHrgxwE7LpD/NM+rN0rq5CInGrNijhzcl06QMJ3zLPfb9Cg5iP9j
H0Fs/OirHiGDt0qgpEGeDJAYTykeYpV3IMjYGeztnFL25ybSCJ1Msdejs8zAw3cH
LapqvVN7cKya0qXOO+CPd7XVb043NDTdNVaII1ijCAD8nt2aFA6KiPRtSRuPSlSa
PgNiD12+NqzbxhE/5YHQ4mdBN3VJ3c+D7h6tS8yMdz/3D1Zh7Qa3aXaEpkaEzxKX
xiHbWnThQwARxWdckQ7+BxqyO5k8ji56aj8mKPJ4wntgLEWYjGQXolbJmSExCGeX
qDyCo+vu8ejYlH+H7hrPHgrzfRkUTvKNZlYkQ40g+uffezNU+Nxqt/zmR5m5IV6E
cGSNHsuaa5JGv4Tlqmnns8mRuptzuA0plvSdOEkV75/AKtWeNpUu7BNN2E7akp7n
7/vJwWfp32WARDQrscXu06v9nB4Qme2B7/qz4qv670GwKs2HDV9aJChiLdY9wPP5
s8pqoYfDwaKgyQa8SYZbrw/4aeh6XkWVVq8oFHk0Cto0M6nJn1PbkKoMUypk21hf
4LtvS8ahcvBfQD/Domexnjati3nV5VqJtYsmkWVHJqerWYNhodwWHNZjiyr0bg3e
3amd/cSqY5xd2c5Bnn6/G8DynK/7wUr85t8KltNbXaNs9+CNV1dsST2YDjHas7n7
UyBC1I3Ga4iTk5vN+SuXpZjEsZ9wgCIu+dBco2dWNJZsIoVAsTZxKWqjNgj7bWwQ
MVwul/ROtJLEBxk6HuEDtPCyxart8HRUCJl5Yg/MPI3ZpY4vb5eSRKH3+qNbXdKf
S+YZRWqF+N0j90wJLsrfL85cMwfD2c/dpeN+QrTciz0JhTL6zZZOMv7wjjv4n1Nw
kSoFJ4cNAfk3vY9eykar41ufia8FbALiNt+yPxG0tTpYvfdZganeMI5JN34IngSX
bnBQU5VHftaLKYTGCaXW75PxZ2+G3pQOjHUNE5388/9rcSIhW/DkFrW4S5vpKQeO
NLjmiEpAmkhMiC/59oV5pqBDFCz8iacTpvkXH2FgpZrpHqLre9F09Ehc7OqCybmW
WR7pknXTJZl2KlmKudaFZl/ndSBHwOteG1V3SXvgZH/rcQXZtlzQhRgQoffuuhP1
uRNH5B/7p4Bq43wViwZRQ09dv4J//IcaPFH1Vv5g/dLhECquXHWIf3j/D5JPC9UL
wlAR5O+eYN4ZkPpQ9uFAxiSoJEq8eAvvz53OYO5f3u9fQ7+3tQUabvyn/Ee/2riE
1BPpsBiz6cRJkEW8/42NdG+IJi8NnMU1Y6dx3jqIXYFKXuFVM13/wn5SgLCxOdpv
jx+QqK/bSO2Qu4yd4+Rrzb7W4uIbxLIxGhBZS8z3VUMJRcfFac8+l/Znzzn3QLVT
gfR2NDwLp03qLNFDEaytgT/k+b/axVtApNLIcBPAfg+wxZ6/MY35Cf/cqElccKMI
+aHPQ9MtmzoDPmP7mQz/Fyu+0dTSBijHpDkkPiOlXUe/z5k+CkuD5I3l45nJUyj3
wigfdX9TEY6KSj/Q3o7NusPJIjVEyiRigNK9NLXeLSnE5hQ7bghkhZRaU9dq8o8m
F4l7kiJFSi+S/7lQdPDbW2bcHrDj24yIxFFDjJOyZkZUBvmoWyDSYGtgHzDRclu7
XablnohxS38bKmGr9GruFghG0WcF4bgb5nyizZqhsWbrQtGJ2NrEV6CUZsdZEdf8
mb6InZOkDeZibKWj52YT6av1QHth0+H1DdzA+3ZxEiJ1Y2sulhFUq51KuncJQT+q
lnsZYsUl8hgkKGk4ItsTsF/XeJnPEXuXWyGcw5x4d6GKyw2Hk8a89NikAtCFj/bX
sAShTaBjH/hN0OTHAT9TDHr76ySChVfaWx482cKwOUI+UThcxPzIYxuavDXc0USR
WyKAqnW6B26o/+vUvv50NDLIT5WfmY74BYSlTgPbOqfDs7bfqU1C/t/cxs59jeKv
F6NUNonF58FZQCnM6Ylrn2wxNOrs1CHtD6rFiYyXI8qBWaVW4Y8BLfgUArrke/EO
wmA8iwyHp1NHR2LuSyxf3Phj26zUPIBWd8KCiUGDS/39AaEhpXLTxnP0AaeOVqGT
3Bx/eUJrDno8ztisBy9q8VS94D4x/M/4Y9IhASq4STsaKMkGGDX+hKzaAJBJ1t3Q
KqhzuhEx5zaMl7qIZUSUtODU9C2TnkXcdoN+gF4AR8wlBvkD81r/H6TtTrTpvALP
c45hy6N4gQx8Py+huk96otHBjJMVlny+CtXi6mx1HdwnHUWnu0p+UwhNlXYRqmf4
w/muL/mIBLNHLUnL3EzTZxd66YsziTZWR1td1h6RtHzDUnvNSinFLip/GEbUNFGn
X+FASqODgZAyJyxxNER8XwwT5AYL8+o4Bt6OuyZGNHYbipLTqc0ko/NebbNcpRKM
wEZu08u0LkKbi8mgOCJnhjXlAK36o8uqbYEjc8HKVmhL2NnEN29BoHpLAiW0kMUn
nrajlDpw8my5R6QV0i/mhZTvG01vaLPqt9uy9AfLjZqCFH821LvxBDfLs6VEa1wi
oWQ2oaqldm9uQJ07r5ZY+3wMhHKhbtp5N+z36GxKPeVJhqPlLCsciAPJKTkPFfcF
zuXvYZNqYwOIqjdn1KBV8l1wS5XKeNWMygxKSWI4U9ZCguAQx9q40GQqqLIX7V4C
peCMG0AKbS7LzwKXLVP77jkaYS70Og80CNKtFn3yc731Fird/ZdgzIanb8WOaAnG
1mg+FoA8ME1MfYvuncA/pA22mSKzpljwgssvNmDi5OKm9yOPl1A5YrdiwyTi4Mvj
Cubn4KWO5KALWb3HZAVONuowLlkpBjA45QS/TENSZUKxRAjSqU7LPOPZPip2OMWy
3n06uHpXW+C/Zd7FCgF8Wx5spJmpYbLaH3q4WxvPlDuDtybnevGX0z5KHeYomkWW
GXka4QIrSB8N3q7v/ThOkKhVPfIXxESV0PUgPilqeFHhqiX5pz/AzPQtAtrkvo3e
JuQoOJdZxwtpNleUlubBV5FTOPSMLUac5lmZ5f1NJUzXOKwAjB7rAuD39jxN0mBM
Mjlyy/TdOgk74NYtUtyJzzz1MudIzJuu99B+vPo1L2Rhezl9XlfDmeZ7dcEAfbw8
PmeAbuP9LdjAoXL6Aj4fXKrij1jONdBZGVIPdsAzEXcSb+uKbMCJF3+mJQn5k1FJ
Qb4MNXvMRNNxqDS6Joo2tLmzRFKPr4qiebZ8lVFlUk0gSHN4V2+pe1Eo7EgZhG/i
k6AZcAzso59JkxDA+l8PduuSWI0FyiKv7GbFwQHna93l9biLDzqsPTlzd7I+kSJU
IJQYb7RM2WqsNUnCoKa1Pf5a8YLHV7VqT/+nxKcwxt7hFBJpN5c7uqcIOu6N69v9
9TL6MLBJQ2xLBXFRi8N4j7VH7U0rO0WVkvRmedmItnW8GegC0XIQ6ay2u1p8yqtD
z4xPYDUc4frXuFdO89uEsfB3sQNHHZ5VhhxszWPqGUVpoweQePFi/zSqBdTIfFRJ
jjGueoO44PWCPhGqvSYLZ/1D6Rq5SgNDRPGsAbquhD9i6SuR18zSUdaTEIUb6Mou
Ko0qZh9phlAJtpRpRcRWVhlMmeKtBpJUJErrNHnELxQigpBFfROk+3KpHFPePN6W
3O4dZF+xX1YefqLNy2IdGLrgdoe5R8d49Ox4vucW0gzUIQAkCjwogcj0ikPbaZMn
jrVseiEi+evuRdG86J5xnX/d52BE+Qk9HAYpr0w/nd7vR8ET2O9FV2vnDu1Og2Uo
vGW6hVYETbL+bqCb7HPRyDFZmzLbEtS0cO/VeGepAZvSw0dR7ra5OFSp06Zr8jTF
MaEIWjSxapOZ2kUDO4rRYAf5Z37ssdD0wBlK5HeB/IhqfhiS8dBGFiLj2x3h2zBK
VMYxXIYnAR9BomwTDUl/7VurinNN3neiBGDEUViQD8A9yivbOpfObWoZ5uOc6DQ8
+a9D4guDx04sdAXtpnRg1577lzmCSBmvBNS99uV+VKx6KdhrCxwXTDhW/9BEKnTW
zyRW9LY9Cc7lJKTNFi2QNrTrtCWDE+8hFdmi8LlLJLFPv+FBGkvmyrFsi2Ryk4le
5mG73xdvltUgES4SxCoZtx9kmU1i9GW4wp0LNUwanOw9snUBnoeXL0HRAF1eneLj
P0WR7hvtGXS6G9q3L/+83hGr3IeAWf454/7bDFso8K4hFwapwe8z8rgsB7TXupDo
DPKDzyuyKp90o+69ph9i06gU5l6l3U5hAN/OyS0H/vTa890knEFPQCKZ32sJeTKx
1oaliGr4CuU38uVKBqc0iEmhEg2ubRDXLcxYc16OE8gLZCrcWgt1yQzr9guA4sWu
Vc+5AvS4k1IOfnz5GQ3Vit4fLGCBEmA4lxH7IypjdAjsAz/k5SKIVpYOFU+MBaj6
HeiWkk+bwgiYUZ7kWQxB8tP8xif7LkH/AnzRJ8WTSaa9i9E2yZVXLXOgDRJneSdZ
+VGPOIwdyhWvFmyPISK0cB/fQAUHzQLLs/X0qtpjdE/y+ZyPsv3j/kS9nT7hdTnq
Xannkb86g3NWs6pHUQKcF8Ewa6nimkngyyxjOy9qM7Nv+IFyxqyx6GhU9sQeFefU
gBMKdPeQYlFZyyZYQ1qIu0sCaXXjrwkv9Dm7xzw6K5UBlvjMHddPBWl1MDRtfx6p
RqM1X2ZzCZyNZ6jv0LrWkDhK+bh4GglrjtepngBdpLsVK+fcqgv3q2SmHLLMh3fG
kwj8AJWavqK7iYOKybRvHkCsdgBnMxd8zlhmnftYj+N8NW8Kyz2U+Y48HORvuL9k
y1tMBQgQv4XJqi3/ctLJLsWuZJYJP28JFieLO2CTnyIa5dyJ/20ZKcgKHJ8GTcMu
oGIOWn+W96w5/CZ1jGRfav5BrB6Dii8OjyzLVFnLUAojD/Ue70G9+pQff371MRgT
Q6y5vkP3+ONmYeWZw5PzW5kt4Ecyo2sk9nznNiG9TjgpQhdTXlLomW9BRckvnaRl
Y1mpFDYTghyQL/a3Pk/88snAvgR+z+bbwTbMf7bLfTzkzRD0/3/MRuCflZAo1kiO
WeqwY/+RGuRnp77rcyZWJ2stQ6d7ZqZqF3Zv+TWk+lSzaMjGfy9Xz/byN+JsE2Gd
jEHGjU1W6E8Y0GbKDh9NoRz+YraHTQmsPu8Lv0EDC9qLGnppofK4adYQb4lGV6bU
DL69JFh6ehkXhbVehOo+9iCevulIjXIy8Yw9dtb2/101Ck4t+LFBb3TlQcWEaQRY
vAMtzzPP1OrcbGUDqR3BR+tJg9GC2ois52mCd26uEtmPEGiOBROp+ZvIFltX6fFx
7FV5+y9IMZJ74nyXr0H2q/HyLI5UJpOSiMi07ORsJ1GbO8m8Uo0r3YFVo+29HtZv
xaQsB9j0Nag6cANA8TmAc5RsUzzESzUmw1lYOvuC3NCuBV6mNXVOB5+WcPQvG8VB
s6D8sbkLekNLtmmTZoomYoaCYQhpqoaU+NW737Fxe4flvLimEEV9JptN/PybXlhO
rzL/Dr/seFF64mjU1t1XaATBaDi3MUUffz2jZn/2hRi+IdGDX2MAdakIP3AIgqwD
fW9CLbH9d5qPM5GNJXSrT0cWeBIxvGM02wH67dyKTM9rZyv1/51giCMnPW1Dnh2Y
zid7MozuNxy30ThfnVirFd2v2sB6qbQvxKaMDpQisxOFZgXLoTgmLLksOiENoMxd
Da+sbuT8H+vKqbKVUrSDhfxQ/O5vHrKCRMWDFjgO/Q02HhprzFlgdjwogQOQY0S4
OEF6JYg67ejK6pUchBt6nukESv7u5USN/+h1QdWdTTGSrdxugBMitAx+0rAec2B+
54jXD0LQzV9IrTrwCdf66sEa48ysoa77LFpPHNX19tQmDSeROjl3/d0bywLLcfDI
8SU3WYkV+/5SoN45gCeR9otmn6cWWh48a0Ph09k9MTVR2pHq83ZXIrnQ+mLWmx2r
cV4mDoe0C6mCLtKseD58WuAMs3OhYTATaVuBFY/LxoWLZPrqUfpNPozZldYY8/iy
njlfUK5Mz1XpyC4geplx0CVHXbkgwWnHwZ788bzt/1kmKdwQwFjVEHwp+GE9QAF+
xHVSwkvJfv9NRcbp6QIUD/8zA++Q+vmUNxJYZ0JLnLUwuzeQpWKWGZe43FV0oPa4
Cb9oJtJW3JBUzbnHog3Jgs/I150yjMPXZJiryqEgVNbYDm4c/uSDQW3j9e8h5det
P+91cuyqAG9NFekakHh3pi8K46NQPJMiz0DfPASZn8P0A6GDJhTlKg9mD82X9OEL
Njfvw2oll9HyIUucb9/B21r+ER+HGJXnqxRvhv9oNLBezzB0Y8XB2yzfNZYdzdA/
iip5szJbpMw92+EmWE4bd3uKzs8OfCE0APvwU4SyHftDIWonyXKmg+su7DTLa1BL
T79Z/eIMafvTnEe/oMxeF8uXl7cbrMBya6VZMgwctExBDXB/N29svqn1gF8gjOc5
fruYjF9AQPPVPx//qk6QJGt3q4YT0FqvHHJxLFFWAPjY9qcdzVu8RYkx1i3rqO/d
zhJjRZ5XhmP6qYWwPZ4O8dcD3tdwA9wGGkCt0sZqvJmO60wR4UwmjZ8T2IR89nGs
KLbG1Jnq0PgyOtZ6Age+SUK69LdjAYwrqzDs1qH8YC5cJH778THPvQm1OKFQva35
kb1zfycYpvmGkNDCtiFKHrMsdR+hmDq9PaprdRfx/XOP6cdbFjpKUeCNTQ1kb0w5
WLH5/FiUv0f/fJQbt//fIVLdO/7osTOvCDuLXK44fxN/sLgcNQkE4c4A4YM0VzlA
FTswok8HWzdaLUqNqQUek5ezVfkBXnUUBEGfFAsGHKJ67EOyjQ2XlC84I0ahBn9O
mnSBod+uSLurO/gJ4XOP715MqHPwpslOkTAwYu20M+M0JVfxatyfT2wGrvubFXX1
FqRkptV4vkKMtX4y4cN4+LQQ0jUG/BfbwRvzWcIj846+4AxQyIYj7/ZoCjaWffmp
/TINAJ1BV6SdGQkRSvupJtcci4/ns4F4myQde2m6BVxt+UiUIdx1p7r9N0sKoGLS
kfsqJDeOh5b/G1obC31PkeBClMBVufpvD5hx7DZjvv3ZMVYjHhOb7oZSO5KLBWdE
mq3tpiF9QNYogolyNrY6+P2yvLvbJt+TZmsmHXx14EwpJ5gIQqWVS6ETUsGIQ8fF
Ptj/i17Ud/UuuFCBI16g5oaXwhsUTlcTOlcidUov/5DZ+7VUMhbfizw0ttGq0wuG
V4WOGTFzufDWP4PUWORzgRvALSFd6aYIrdQEDG/h7Mje7hbmm8DhraX5k1zLUYHF
sfL/qxdYkpd3F1BF8bbLKYy3swA+SPRh1jNKmx7bYu0ACMErrM/jMjsvpBN41soY
vbimpA1Daq/4FxgqKmyDAayhpL31jtczrJ1pMuwMU0cSclQU9XdqU9/etupEMKjT
lcLlvLoVa+yIGY0lYSntfMhaiFpN3kv/riNX0maNcw1Lm0Ow+Z3jn5n/AdSV4WCn
2pRsUAqT7Svp5ghqjkmQzRWX9RtrmIyxrMPayPbsw6qt1h7LZvjZGvIB1LVwqUx0
WG6j4v/DVbF4BeEoBzUwWMGC1YKpAJKssPbu90PztOB+2GsTQAAKY9W4oyferk1F
xidk45yVzzJFXzrru5D/ZMILaEzKGsKmXLEa6c89G4QGtwqof4bTDVI0APtqpJ/U
mfp7W8zteR0HnadG24ngmGA+xrsEhET1QiflnLtqk1iqlAJkd0KaMyuBtn+DBBIh
Op6fDUB2MZfrggjOP7qN/iIR9tTZHNXNN5EOVBiHQSnOdMaHLJz28r6dzoAospXP
WugnTjtCZg+uwxBS/nM1DBgqnybLYbYBpUTYPjQfDbFeiJyRXYA+r+I0N4jeXOa8
/7SRS7dCcdb0sFRCFKEGqBVn6mYuYinCFkyRiCDhwzEqhl1YrBDsrnbPjjgBPYU5
GzbGvrR+6Uy2KjKmFmpbJh4EsamH33A0dqt4lj/WaPfoqP6PWBD9yHQRIxdUFh0D
CdHK1m2RAerp75pVVt6XX7mv2GxKEio1tcq3y0E8mMK13aMls7NalS20ffQUqMe3
IJGeuusoWv/81SlcKEayrkyas+hKDHLdI5+M5ma4Z6miCRsvO2Mbb2/0PjIrgU2e
2Dk7d53gnwypkmRLK/174q+J8D87JiCSfgQ6dlm268OsAmbw6p/dzkPaJuIs21lE
AhDGUbsZKXxJ2HGMf+TSrI1F4W638APfjTgUjSm1tDO+HS23sOczVk9N4XSG/Ebd
BzTDVQXLbt9re0ZptiiFfPbVkE06fJB8T/GwG1sDHNLYGIDXDhxXDCmJldivtmzN
U3dgDCm+axGWox7chhxGHg+NRaquuMBq1pmx5S1KhKmPSfRLgp1piCuckr53fdKR
yFvcW48M97BPbwADZ1byOMBtB8EVYZMs7bt1LAeuNAlzTJqyCaexFL1yhK+EbZ9k
1LgVAv7j57ziGDCMuDWz7VoNSnC/X5ObdZkPvKYU0evKwC+RNUDWTl58EtguopHU
dDXwyowxusxWlp84tJM1+sKl2vydaznLU0KrKaI6NsiTxA1WVk7DXwuWx8l2dLwM
Ia+cdm9iaPXdgaBT/ZhfE9hz+QvyLxgyqXaKDNmqQDvnjan6eCs+SwlUfRDzZU06
cCs1BJwhEehb06yoqQM8x7MyyfI+Y/rIUwvzoHIu/xJkRRctXd5VLCX7bhr6SONe
omSBCts9FQUyjLjgzs1iOaBFZYAyV6ftJFyzEopYIH76mdU5L4zRU6pcT0nJNZPm
kQt7BAU7y/iOPDPHrBwtPhnIO/346lxCnBbQ+OdqoMUIMAZaLXcwicrnq3Qlq4an
aHy9tLS/NzcCYv5yvwGyBQ0el7U8irpUiZMGuAdYQimBiD/F5oVX4yGhuR3mGKlN
wxN5+EFgpapKRaV798fOCpgnHLVmdGZPFytQpvC4/IjNA6I7xwo9roUy84Kf5nBV
2Al3Jg/UZEz00jNhAvtWTqT0mgXAbHcdNObaLnpA9Na5d1r9+WiKd8y6ljHyZ94A
8QKFyVx38+17lL6Vprz35Byvig4zL8FKNhRABAsXLm9fS99iibrT47e7Wuxkh9og
QOdAkSziC1wyYG018PSKeOMk5cmQwit/OqHuZKtNl9z6ogkt6r48cKQmS026fyD7
AGN1tAza1mPEjkLqPagCPK6SgPdSjJoybpw0R5DQjUom00e84mZC8JTcb4I2lYZO
diUhSk50JcvK1w1zGh2SRbSa+XGZWMLDuL0P/w2OyTjlfSBb6ddUMhy1D9VFpTCi
GPT17wwxcML5lPn4GS01RjqoDIv+Se0vRo8pgUYVQQTAH/IB3QprRaa++Wmj24bL
BQZbvHgRRZGLGLo0oqVu2dXT8Ku+gufXm7gBIu2QwVQdMW/SdfWnrREKoZP/jc8r
RuysSlebFttMwLBd6Rku1VyY639wtZCGkQFSIQ0242I+XdgWKLkborvD1qbdL/+Q
Urgn16uBpP9RHCowBzg9s87w/pZyss5DK13shr7OlEfP/5le7JbC5AqzT8byFraD
AD+ruzOq6Q8vJUunH4OvDz9iYkc9nUUX1d1w5WPFs7P0DUfdqJQ7bbfoSNXEwTqp
8MyhKnUWIh787gI7gwarhWk8+edd9WCCht+xQHWyAk2g+gRU1OBBVd6rJqcrfPZo
yNLJ8u64B2xXI6eGTSViXUxojAd+K/841xnk8YuztDtPoGsJf8RNtS+Y+Q2STZUf
aMa//dwUcw/EsPazZ4Npzi2av9pFH4rhp3WDg84wsK39rxuItFjjQElJFLLkm/Ox
jaJw2Mb0eQMHsLPmsJRvSu116o+JH84rY5MuDwNS8AqqLyaNnVxYA+SSuGPs5LeK
WiNd/3S+daVSUhGB3D6xJmNDZvRG88mr0zyWtRu00zgMFPvSAvxmeULWK0rIB8Ju
Nv10VK4d6iWHGC7peBi7W3v0zIXKveH5JUGxMtYeoiVsBO5B166eAqQr6H4UGJcL
9NoerqgO55dR3cpN1lYsWtkpWmQqsPXaLDl4GhJ2t83McnG3RwWirVm5EXwsG8SF
n5CcnXW9j2JUnSa8W3pXkVvtVSIPLPZSpCftWaQoWdIZEwEkEBMoF4Cdkp1MASNt
+rA/60jZ1xCdZXhlrp2bgh9akeAn7UolGO6W3Sp2TJX9VIrZXhb3C8wLIpE7A/bD
KO8jHi+2b/zkl2rByfSkV4ZPcUvIiCjNEbYBHq73MiUq+fnDYxKhvOxYPGgKWYFK
BV3JlBVy2GQIWYFHXYgs7XNZjCKFi/DdePIzROKOZC5sJYaN0ytHBU3gFkCTee/R
RuPTi67bfXli+ZEqLEmsd4TKdjsliD1BhaDi1ttrUQH+4wN18W0Wfb/RQAtq3yPv
63eXT10tei0Og7HzusXKFYPVbWUxasa3fIm5m8Y1pwuy4n11ugR2MgttX7cPXOA1
KMMN9rf3dBqekxCFJNS+h/th4ulZzUpOSZSC3PpHMXXQyKG4bP/3149YKFJbQxir
8PYu40ZMtAFIsQaw4NJ8tLNPoh/dp4VASi8VU4StdR2N9sQXdaqM0KjPxIyIRdgJ
2oR4unETwKG1n2Sw14RZQoS3IuLK5oQcF7gfEI6RpXJUQN2BOYykwTqqmaXzy9WD
vjl740dfaHszK7lXDMvUcXGwgaZ5mAedKClRxaHBYSYqR2X5YdnnT6YfB1bkprKI
cy1whBjXrUB6lpMwYuEkC4yVvJRXC0ZSM5+5e0YEMRGgw9jyKgkOEx5XENRfgzuP
phHHw/YHykTeEx04NjNGxBLjI8ioxgGapR1x+OfValYihJa69ld9h0VgefY3DZmc
557pEhmwdm07/55iyEB7ih8vbYBHZS+HcLYUS7jOys4oMnwfaA9JAWGFljTCO13x
K7blmPbtkMniWEp6wxgmZ2Dq/cR17cETkBMTmLTABsZbNGzvRfWjXJCb6NAnjMFM
AT202+abuoIklJCrEJxfuGHMm3c/2DMszyFEbg7k+Oasxx/h833ZBiFtubx7XoHx
yJQsAAxjr1XOdzbpYSBB14/umt2qXCLPpLU/mzCTTwW3Ij1Xr7AnVS7bMHRaYSJe
tENI/pPQRF01xRF+Cs+eIKnjpmOaxZzCfBfouJ1+qBYHJlXTDX/YTixlkLIpNj/D
FiVdFO7nVwSYVbJPd2oUXxDLpaufBI2qz3+kZnmPjF0IypUpv+kXsV7ux9Wb6JIC
FfXuuWTYAaU/8cDd9ctFbNNojb1F5FNs30nXpA+FmMnbCBB38YSir+jtkyXeUdrQ
jc/XRA+7uissYlbV+I2cXehC9+pBoStUFAnCRmBhdE3Sop3jv/maqaCYyZ2v2ccn
esIscol3fqinyjMqh/8LtbkzvBaZ7S0qedPSOHM/3M+sYGb3JrElC9C7IrIbabaR
hZQr0OE/c4hkaRD4cpkG/d1QRczw+0I1efYJu/fn7elX6AXpxs1oad13c42tp/Kx
X4iFWJsyt9o1ewun9tb97U0VzXbVVHAZEqfOB/FrV2D0FE2Bw30p8E0S4M85mz5w
UDg1TtoXWtVOpOmVpiwJokTMMb8DPOjwQAV92ITW/OpfiDpby2RzhABkY6mDnpie
d+wY68XJumTgwXDm2jhims5gIIhgW+t/nlPepLkiT23U9GUE7HwfFv5bZGRDJvEe
L9uc865ec2kKhuAgA8oWEr93HOAJMH5aI6zzz7pbIRG22sTrJHQfiVviEMubISug
HoiYDEVDmojfIR/7INCEo7RseEK8abMwQz1wEO+giIiYt0llmhzKfR4APOMcA2t8
rNrhRpMAgCclN35+s5vrQEk2j2P2PT4oNEV59VSPd5EPC2xaLVgX+BsXRZnNMb4O
ocURrvAUWofI5YsrZbtIZcvfC/M6K3iD4sLyNmDRGVMRNq+L/BPYi7Jswr4DG5R/
ZqmpiaAMsZ1qNvMF15LEuIz5O6Fr0O7UZvdkeD4Q/P7MtHgHqo89nIu7ZvwoOEd8
sS8sZtiaalrO65YuQ7ApAyRT7ePcbzpbdmE69ERotWMFh/QYr3ktybWmnTJbGCC6
cCI05tHnh0ZOqKcebeXXOHUOTauFatx6Yr07lWfv6+VDrSIX8xBg1C5nhr9qc6fd
boGVXadjb1efWkzElV6d2SgV79z0qquAYkpSDa9nSEMQSU8BYLRmavlrslu8MaTW
z5MkuqUodPuij2cMooRUYz9aQpMkuA1BowWB5soAUq8ZWcX4Ttw7kOKhf4s1UeHJ
MU1Q7trZBA++LVAcKZckqYcrUniK0E34U+dT5EALTNsadq4U/bEDwvypY0DTbzqW
c8hTsxzAt7i9hYQT0z9gx6EqGuShdxOQPFRlKKdQzFWIH1p+39/q0nwG8sZ9lh5p
UvJzfLXWxQZJledgdWPrG7beZRVZoU3PNWPe3Fmc/n73pJaQjViTjsnY/R4rdI0c
z6YVsMTnHZHjsjQ7PYs29efs48x75KCzjDkHzzpoUSbzrCDOUax3NYuyFDKG8MKl
eFJrs8yHfQM2c241CljQuPAIzlh/hkPgkdREOvrtVcUuyfIy4armANctVt78+b5D
0ddu9+5mbHHDsmZInLKpy430dda7/Tw1Aj5JUdjEejD9NFR19IeA2hy9PptgvwdR
zQyF54hTDLzq2mM/Y3l1zSPrToOkZq+Xlc+dK8NkmBUMx7MZsbQf90nuqxGUSW8U
0CaP2bu+AHc6nDjiMBd3vKO5kuECnOkPTY4Z+JneHvTXArwi+TmRsrikjUJtL9Gy
eqsmhiTfYD8YlaVBGY4HrQcMRYaGd3tQLtVZQsjCbYXI7AUtWlzUmeAg1gVrehiw
++ikvWTlsHj+C/4WrHNp4vETilFkux5EJuMVedyiXHH+Q0uFHVcaFh+LdZUvl9cw
WLjvu673EUA9d3P8r92sw4fZ3q4UHo5+0Zey3Id7skT8ZNVwvQIYU6505VOXZObI
WUDVhR/RjDLh3HxFdVvMC/zVTwItxkJyqIMUsE1zt3stsAmFEYPaYbYsJgszYxHC
jPm+KS0G2q/xBL6vnf5oaTi/V0KrGjEOZvSSQoEkBHvI3QWoW937WbUupvjyPWOK
OnDSx3WXlttwXogYFi7Zv3hHQI4GjCTYhaXquGR92pwBdmNvxeuh4IH2fmx9uFZw
PtC0RA9MPBg5QX4ZqLrlugm6q7TK29uVNXO2FAzqgcR79yY9eKwVCHPMliX1mecm
mcvnezXCuL3/OfGpGU0bFfN/IU/exUlhe4sfe15aYMBh4UzsxyUWt34AXyj2PV8+
Ghm+XxU0ZBQL5XX2oTsB3CS9f/dKRNgJCyCFBTC3RW5DHIdGu11GkpBPg4wThgpC
24NimsXPhQdpQna1UytY8s7LGHtbqubEBbJ7rgncJwioBc4TdYkxRId6mTMBhW7X
TYfGq+UCa8mXsx7IFB/60CYHbdezREvWSR9He8qifrnGyGBvOhzIRCdjMRh7zaD4
wdloX/AoHFDiAx5DIhgA73O/0NNsN7g3c5vnCeFmgoTbfcM5mqrIDF58oCOgnlK3
1aF10CdDjlnNqkfEcnmzfd49S4Zn5iNlPyb9lvDCv89MLWtOsgMKj0CG9ZX6pPMX
JDO28iNwkRcR+rWwpVA9v9odoZVxO68wXCyl7bJpNJ9KEvPAWhVWZrCZuwoCXJKw
/IfFDGzOLjpULAc5MkRbsWLEAAZbV9fdqpzEgzzWnrf8kpBc/O2dyuoN247UgamX
dpOb+hlXy1h54qRpPyjcFswV6axePnZ6Greg1iFAckZfiZjxgp6jNSsWRf7B0cHX
NPzbJjKloF2vrcQhwh9gmnRse5c2eawl86KDLejhJeDq8efm3xCXD1CRxLOKSDLc
H9u+fI2tj1oxhi/LY1Mo9ApXLL4VUCk6VmyGi8xDTL7+mnDGmMa88nSofSxM6Mhg
8mlPX0lckRqQfZ7VuavgqH9yqbOwIsBYi5BELwOtlTZG9TNDCMkrg4gamgQQDzu5
A1vv3axidz98gCNxSbqc2fqJhfLxpG4KpwlOVFYOhNlgqUGnCECb/QPys+XYe+WM
6M/EQoNsj7aNeroN+FCf6tTpgOX0z2wToq/eU68DuSRNMaNqMeD+SVf+UlpWdpkR
pCw4Eo7eM6hm2awAUWl2IfvB/vx8joLGGWHffiwlM9fh71QPIuyFRgnsyHxYUbpg
O09tBJZi5Xfm7uIttDpnwc6wSYXyTSn7SnCZMbnkfyJOmrSm9M04tFtDpRFv5PV3
nALHRsfol6psZ4OaFBQsrAILH374X+NNX9S02ck8TERtADEMO/uH2acPH20z99+w
06FsaeWn2rnT0SqOOIQmvhj634QhzYVHW/bBxbDlpVwdfoY3O+zhm1k2GwXZgvlZ
pqV9hqitZU4U4BxTfRVANpml8MxKdS6zTQvr20kiTKEqHugkSmYhEYylngVugebX
c619eg58fLkbC6uCALZc5J+1cPeBJJLuHcFmX7x39USRAClGxXwx+pThW4o3Zp4a
QJXyE9CouLRx/SQ+CcFqQanoKwSUWFXHNSqmMjJUNeXLNXm+3OfDIjVFew1DRG9Y
ACYHGbUeoMng8VHZzXyOZ4jNghreEzktppoAAP+bZqfFsXuQeFxWGmMvosYwMhpS
+n7NhrqemdsGGGyP5UyM5ouxWmsmFS5eCuj8oWZnn6O547aQScLx7CsdLQVF+g/X
lyB0dGwDxhiOH+4P5E/AxNfjw6zd7BoV6bu8vQqNCS/KvtnF+vzwH+/H/WueHc+T
uuMSlyH2763euTODB6mg6Gtd7fnboK7tymRqqVLppx5J8rwtiA/MTu11cCi7Da6X
21N2FuKJtUcP3sYFuGOs9XgxNV1vCgA2EPazuFwDv33f3rOtHW+drtuP/7u1+Ojx
1wkh3yczfgJUT0DoK4BlRF01gekp30gfLBJG/3GaSlxKs6m5blt8YOEe2t5c9LBY
NEdb0eX/IC10z1yPpBV1CgrDMFVaQB4FRRrwR3s8eCTkvYohYrXVeQk9bwGrfeF2
Yb2FnZjvmbAD6gjyVZXONIG2SznOEizvTx3zdySvpsGJEXsv5OJSx0Gjwq3rSndU
5zMgcxwPOEK2ux0aQBTqQr1gRiioa3Gc9RqaFKgp7dK6VY1cUq/yF6MnZhS87o4u
blaJZkhJ/BXB1pJ3D9g1RFI57AsNyoE6DOBD/9iqq5oeXwPj8hpptvFNAOU5Bvwf
nThPd9/oKx0NC19911M3ItsYK/N4twken44Pa0YZC89RdGPTOROt2htjHye7Mrg+
eUoJ6CJM5sAEUeN4yp3I5MDZxJViZAeMZMdv1EjTFsTgZ+++RPcrj6+1bTIL7JqM
CulnjR2zdD3tuoJADEIFnmkRdm+AA3rhzoIg/OvB08nP2F14ZQ8W2rkoDz/do5Hx
zO0Rq5j8cEQnlBPqwBgIV3vsxt/Pt2IB5J6LKZhj+kX9UVFelbgIAWC5v6dza2yA
slZ/2nznldMGDOubUDxKHACvAa3QpDUDVYJeGv9AlO59Vn1bAUuJRkO3g3yjg2zp
ePlqTyWoQW/pFqzogKCypqZdZteIcyXyEFz6WS6hQdunNJbvvR6AsKq7WEytKBQz
wzKP7rABiA8U28PrFMnx6XrBzlkuzIXYfaZK5ZfqNLKzbOLa41x+d53g3VRjOedi
SVRKCh4FxQsDDYlr8S9fH4dBO5CFQFCDCKmycwGYcdo0FsAyFWYpvFNlY+lbb+j9
ti8o4KKnU8/EE6lfVux7Um33rPLyBr2q4cxWwKbRL+FvltJ6qZfaQFnxqMoQYUIh
nboS53EUSyO2Dj3o/aSxKEhDyE0ELVYCrR85hej5u6U/Y1YjQTeUwslXNEXkl+J1
luL4j8DPsbuo2JUWPWa9FrsqIBwSdbMpgrzG15BZ1s5GELoh/9W1zWCBhfOlmn6h
shpSjBQYTYot8gE4JqcnRhw0SVPurqL0JTTitLkbEacaS+yIzme2WdNDezPioo5C
BNFk7bTHr5e+ygBV8HtcSqDtYsORARtFr4TMxALjklIfu72MtTW9efxy7NYeTVgl
HsDRUegCAG0ttZyhQcKy2PqoPoBqE3BUdu+dZPKgN0Tj8BxITmBWI71rb2PC+Gh4
3d+rbOq77gGCtQv+NsaQ6wdAJ+kVCH+q4FzRFReOJJeGYwrX/lOe2nlAWN1Kutl9
DEQDihIZgWzaGtzy+pizpPbJUxiCCsdpzVKs4nasX+LFhHzMEuRSXfWndCEbTX4K
9e7s9RA4ioYTNNLCm5La1H+ej+KZSSGtnSpi2sPN3GR0GQU85EH7cXRBnG2Rrv6C
NN2YMP+etU5nlSeC7nV8I5Ek6Pcp4vkXuhcxduzPfzpvtjR7YafxXR3VkFUXW9PO
x8qeDj2T01wPo9GORXk5hkyjqRFMVNBHn3IIeA4EKrzHYof6OuW23Kf7QYSejnAT
L3wNjbD3ie4sSVZi45mXnw0nPNeTq6N2P6yW3E3zVdz1+gWFXWs48TVN5L8aQnVu
tZI8EzCcGtk/5zcjUkwN3zd+qmynsoPmDf8xWWtJHVqTMYp5cDAjrvQiFGJ+Ziy8
/d81NWVeTInZDltRUoYlUPHVuhhUxaHjQiB2ix4+VDCj7JHmzEfIVC1R0BWkYfRn
NXQO0QjeiAjjXXebbDQUS21tXZPAcI0mb03dpZkbavDbenoZY7d8UKEYmCzCV3TC
U8Zeuj2cFYYgZHZVQ7TrIidzP7nws2EoBIc4Vd3IJzm2lvXlS8Er5l1g8b+hb/h+
gAPrAdZ+8wsACbmRJsFdw2tTi+ECbCqnLRLhEe/NGSsb/uHfbjyj/Pqzx+DMr9qM
5kZDWvbLoHiv5t/tQj5P5nMGUftG6ii4CdinnK6BfGpuAaQaFhTithKtjOoFq6Lo
MtMHbnHCyMErzZd1ltRhPz8uXYh0dIYqxOFjLUy0KlPK6Fv2UTAE22QzJYCeXJrK
IgzO0Qj4cOB0Get4UAtjGoG83VsquLggpDvRQn8CzIX9VBcgaKNC9/M8hCLhcyvM
zA8xJPD+fzi103LQ0s6q4VI/qRMCW1txE54Q73bOu3GIhmSPuZq1kZH1awidYCTO
dj5nGF+7H3bK3waNfShxuUBtKg1fpC7ox+ssE88xQC6x6AgaXGo+oq0xOs4wUMQA
/Vvj5Vp+1fWqIp2jQadNPEfeaw0CAJcAZCnwo6nu2wbbftw68RbjE4DjIEl8T/4i
T1U4RASS9zekVzO9KjWwebsnS3CAWUda9wGulr1VBkwqIWj+G/ksVUDvXsZ3dU4J
8yOSQuiQHMQ3/06Yn3ov53Rinn9kvcyr1M2VgmEcdVr61AjG2iUBiQpMFaYQSLOc
5M1UKibLrq/fKfQ+eeT52eCYlxZTxLkHCGLp6NS7YTk0ztM0OgeyAudevdzeOkuL
wArppGBs23L819Je1VRcY1DqIQTfFBQINUY2RLSepbRUeDw5QhZFAY0nF7FSxQgT
eMPJ+yaFRCM3ILACQwBfJ8lZmKc9OwFQ+HCjE42en/Kb28QV5MrI0nreUM6TnT9W
p/SUbqFHseONwyyAy+WKTS6cYnGZpxdwcxLCsOAblKQXG7NydLqdzMo1SJUu4wa7
Atyd0iKkaCOFPxUw0Q/kNelDJe3RdeCwRNJr93LwQmUi2va+bXF8QcpGP3PtCP+a
hXetxYCrCrCl4rYnf/+l5fOgGfmvcDcwdf6jPMnfwvG/Xs/GBqAvz1qSxY4QwtDV
57EkxUq3lWUVbkla23EqaVRIvzeFGAHgkvMHJphKRcdPS6LT396zTcnGj/0AWpOi
uG7BZXHr60Qxd6OUZXfNB4G9n4VgFq4VLNNZD1JmCHz79M4BBwwiYMGWHpLdG7Nj
RtQJsuW1LQ358JDVlU8NUllz+JMqtYxpYqdBN7+jQUGdGZLqCYw+IYcszCISXwFQ
fhGQ4Y4Q6Q40frrWzt4JQGe0Cx3m8DUblkrNG6bbI10s/0Ila+9+0KWFrBCFXLfP
5ARX5+kqpv5nZtTSVg8X+9xWFmYD0TGwq7WAxr/50jakJ+MY/1OrnIDtypp9Rsda
9ZiZ5QiGWHGDuFIxTR8LQIhPnLSH8k7nqyPrsZQuxX1QKsZnScC5HE0Jq3ftJwxB
q1z4NdaVIFZFyDFzXjzGbvp4zAeUabqFIzxYlwKbBZzPVBCMmkRvGl9EKvPUld6M
nSQLyxwHKjjdm8xbHOVQKZHVDicsNTngJa/XraHs68iZsnnnKVTYro+HMRRqWx/U
OO7W6q3NdVrbPPq+0VhrDUbPPjAcLcXv5b+L4PMsFopr29JQdNO2FWGswxPsmXTW
uv8F6LlKgzcffIIsEUJObzWnFiSpLLoAx021h/iCexRXxPorHgrhxVYacRkpTBdM
CXxSuwlaSl6Z+5uKVXCTT1lVNNtSVJc11C4qGvukOSYzhiwQOjohTPQX7TYL3nJM
9+oHPQkknNkV76wyQoPo5uJDTM8s1CcnM3PNeXiTWSjfQUCjKvlE1BSm8YqlA7I9
DlYZtIGGr0EPynVz5gXRun19BpsHh9W7wJop40XaC5c8Yt/dCMuGJCoVQVgVoMyC
N31TyCGlDD9Hd1Cv8AwbOaajZwYd1lx6Un2K0o9GBdwSivJ3d4TZ6zZYJ/f14auU
gbePX+ybsQUBi+dtVjgJUDcOoQlFS591AvIOctKgcVNvcD4IW8QVvTwTsYlJH+h6
Rpqt++nAx5Z/N2OQ5Nxzy6abKTuJAcjt2Gziq18gF6nO9rdPgagQ1Cef1hrSErKm
kV8Q5YTmDhV8mbxOoFJLgWrJPibaSdUY5/mjbV2UA8kqypfzt4CdGBAx8j/bEANL
ZlW3PcOBQS59I8pGcHMI5GJISsS35i/peDgLgfQJPQWvW/ce/je4b6sczZvDgtH3
qGKHMf1z7tiD3j+YA1Tea9b/Nan0cN3t0FE/qKE2Of6B1Aumq1XOb5v61jxNL0BC
MJgn//WvZ80F0I/S+cVmsGtssookSxYW5uyMR3Z5/1ABmayYh6qnaBonFEwK+c/H
0KZCK6AkudZ9qRyKyR/ifQyAoMyN+Ybjp5Xi/uBLcGVs6aSZqqjtJphqYltOJggn
knnGd008/r4vyoOrQoxCS5JvciGnI4nUE7jzVfmoIMVZXe2OWfYnAQE1oMkxz3PJ
aD00WIA0hqdWh61yjeD84r7uo/no3o/ksoSNaBwRueiG+G6/VauquK9efjkhDyED
DIOBuVS+JZdmqJTMv6v0l/NyfuiL0/rkao4Bp/5iC66hIT4Ly1Rx10Xm55W3b+Hq
HkwPA9HBZcouWC2tQ1LCSif5SmSZWv4TGf1LhZrsDFwlcv7kH5bnfvFNywtGkoXK
w9LcZ1dj90iFUyEi3QkyLduWnbNkKYuIdsEAY9mH1IJMigRz1qEE4wKM655lDIEJ
b+TBMKGnH/jTHMGnDAqePU5wAJL0hgpj7d/Pu+Z5fd2fx8J470BV1M8ewaQAbwKC
yQM4ROXoYtJXXugMGwd1IAyVHMXGx/YbzFDjJGVIbxcksGhHDsTuWWbPOcyoDkeV
C40RPK2NQypY94hFTArCgLh3K+xb9QuPVZ2NWLtruWNuvkLywK7FekoKkrQqgwNV
k/G2EJ82tLS2y+oSeplYVCRI05Gh/GZYva+qdu95Egml6JotuoxPUBEWyFtfzJEh
eAI7H73EX1q9sgExb5B7keslttMlHU8JF0W+N9NVcDtfVlMK7CWPxkhSlKw+KB8M
Gq8efk9fyiBXo9iIbEkbGoFBBFYmvoECILy0Ahx0cNpJL7lCT2CCbbez51aw8TWM
XszwdIj1prnH1ndwa4hrgj4kwbfzAzlMVkOthnBFNiGqHnwbuLiPCU5lYMZxriSN
yxn7yj76EdbBAXXCDj1rP8uaMC4kxRpt7pEqnk/LvQ6sNOAewNnnaiRvqEgTZOeE
S9uxO6XyLCp3SHZr7j13t1txgaa+IGIwcwuzLxgwOBTG7F2o3H+8QCBAt0veYDhU
DjRgmqrRocbCyXldZrAG0kEt5vgaF80hbXTdvKX8ICSl0iAybyBlql0eWqOpaFu2
9rFmGRKG2cFf+mGkeHbue34QxTpXY8nWh/9xFUZx9oQyJK2PMqc4bD4qc0onHof9
0obBoqekfxw9kBcyUlD1YKuZSnpW8Gms80y/nBWcTXKmLEfT2fOGARU3IaRbY6V5
WWIdOVQIUF9rXc/z2YUWQinTRRGIJoJlC72yJCySdRqw9A/rAnksDUzDob50PAjk
yAJQd8jjabpS9ep79Earx+yDMqWbM+w0ygic0zF7MvKqYGwfqlrCVTf1nsW40KcP
ZzkcAzKnVyxuT27bmjZIwCYr9Xw8swdaEHHu/8b7icDJVoediDbHkJAwBwYczOBS
Yk8gEZQzv0lx8A2/Hxd88ZHXmaukZd1KEROIqKPOyh2M3JSDPU3SKiiM3DZhwGFk
qsNdC/oXoWCEGK4nfgtW2B3qdYNpbRFifHoAoPk5H8YnKPMu2934iNGjmZOy0Q+P
Qp1VqC2PBFZMy6tEy+Kfsl6yMCinVPHAcR3F2MPiAjxQNSpTm5U+6k37wF1wK8Jf
J7A1KZZzcIDqYeRmLnE+az8oWhqRcfxwb69W+voaMgIRSiC4mi3RLQDmnGUTN7GA
v7+PfaXbO0OE30BJ0svtWqki+G8+C38mUlq/eaglfig5bWc+Vt+tg/7hHfQlhSGF
FpeTTLJlIQXVPiA7JSoJ2zrElgxfBpw4KZSGahT/kND4LJwUY+XbcNjtJ443Jskh
hNSFXEU0ktu7Vsgbj1kawLBy40qsL8EKvTcjV4C0QEuq+su7ioRuMBqG5KdZAKh4
n1lGMhnr7h8CpBmC3TsniTdilvL4wHrcKxGqgXFvG6P3auPTS8qrhUHjhxZ1uBim
WfmVdtUbrkQxbVRhlilgwAzH+O4K67ld+8TXGDdiDpuzSjsb61C5wDSPvyXQOJcF
5lZJpus2xxSaGNQw00HEWQ2ebgmm3Exb1u6ZLU+PwcJAawg59qE3MJO/mMS9IIxC
b7WfnGyXK4HIBVFpN/KfnqhWr60gaXJwbZPRHkZJehqu6WnWloXrdesjMJzMx18S
29o84oSf3ZKg9gN96CjHSxdIeP7j9GYG8YpiTbvDJmpmCziKsFktFmqHej8BeKRv
lFdryCbA1tnAaipMXerFuLiIdyqCque5hHD613CeH/NtrdVcBCxHwCOmttiYDtf8
M4+pYZDxkuhu68QL5Aa9ogHMChiX7mxHh4eUt409KcSypyDVmhnlFJB600z/fzf/
6kEVWuUw5jFA0Aej2rubcmtrRAH915YssMqqknEP0WI+T+qJUh8jDTQVutShkMFI
kRnqQyEaZVk+vEZNS7w+VZDQuCaeY2d4DXq/On2pf0rO8ovG+zJTOzUxgimPTgfA
perpFHffAPmuVbaW9JhSHhFpA6dXTCrQbwsCGl7MwevLJF7iIggTCJh5aGOssayD
urGQ9uQ9Z7f4zUkSCN5CDwc1n8ftqqSF/DyYhH23GE2PkPBJVYg7tmmqodfMpdez
2RmUuq8tyl3Y070nloXsAff+5MQbHdfkniS7H2AmJN87KusAIGdf/z7fDBgKtgsJ
WCDiy2Mgp1L5+JdJumI6babON8rWUmezBQJj5qrsRO9A6lICFaY3MnZxeTwNcqdl
+2Bdj8onopcTMSDlmrPCYhEAX8VLzP7eTxJF18t8aRaFyrTLtMCtAtmFeM1ffKfD
Cy5vmtBbtHO3Od6T8R+fPNdD8L/TB0SSqIzypn6/yts710g8MxX8JENFWR7AwgvR
WX6WxAx0THy/fJmkIJmzCHgxS9QrzU7DAMJEsTTaBvNBnC+f15YYhXGskx8n0RX7
R9Og2r2IIovMsskMmdxXh00OiHWts9TZv2yni94Glm7VvGd21y5bjqabX93Ywu9+
O6pzfNX6n4WHn7wFdyCOcUv0aSD/d1WBU03U8hS8Xo67FUrG8CEIRpGHB2ByOaZx
ix3JmSU0FhqL0E0MuIilL1meQ+z3bS/RLvgVK0mcsOnpkgM7QQf6AUmfwVpZQTEZ
/A8ydg5l6pPzlgM7vWCiqeXMEuwrbsK9fV/YhsvaG3mBKvX/14jtOB5UUeBD2D1t
XcucaBdxYvIf7HfaRYfe8y4y13sBiXHduNHfHW2YgeiJB8GaH9UU2ru6aWLnhl74
puRXtjBqMu9LD+/ljg2+b/Mug5AFaFohP9a4PBUri7pzuuP0hOSf1pXrC7TAr19Y
CxbZeSyQqtY7pnkrv9GKlsFniXLXHoNpeFURh8cSDGBNl3fug+BKO+I1FaTFVj+E
uvavo6+MW1EEtp5WNB71RSxvA36KTXk31aWCp7dvyWrXE+OzOGzV05SZvRItQqqa
4OX5leKWwN7S3DqVwa1lGNitlyXhsdD8GHKViGE4dE1OiXBDPg0FqU5+/NV3bpq2
uoyN40kp1bK86s4q75X4SJzWQVL9DOE/Sl/eQJbbO1k4z2YnGe4JdR2k3edsK/xV
kv/xQqwsemqY9DQp7yWoRck5qC6ADWxrmoSGSugcaQVkOLqJANh4u5YBJXYVJw3w
8TdXzeUJ092m7KURhSv0p+VbxKPtg1j1RNBoz/Ev+0XSNVlM5wdGI12+ELkezKAx
ZJ8YdrxqtP0++w/fXxsdRq9M7Yhd/q2CW0ccstqpZqvxRDQ8YwbIIv9z7gfz/qyY
MJJFfNz0kYeFHllSIYtgUfWvLTe50p22dvfqOjW+6n88rpKpmtWC5AU4vsskp7WA
a7ITRzIqH+XCexnpKcrJbza6lqZcBTVRDmkwptuXnAxFI5mXKISlgvyO54sa+h6E
i96YTgiJ7MjuwMI5UE8qzmmO7qreJtIoKcLLN66q6DNVneGHfud3wsAaqPtnYaOp
RXACb5Nb0IPmVWFfiwFbT344CJx53LIQHBz7Op7lXN1i0TCxGHA9Q+S+AD0fF/Ji
QnhACprg8uFx5FAobkWmRhX0KKUFKfbIDX9/t2nixzwEoioB8D0u0TDYMDKnszwZ
qZsbN3M60RWcDJLkAcFw8slxzywM5THWr3diQ561tqoS6tgMalCbFrHp6M8kgNi9
4hstCYl6LhVVSwMP3CXlyzI9/GnQ9olPeIZs6qNLjxtAwHHA4YNjzbH1OPH7ShX6
I/DfBxIeITYv0/oyLZq1QJEMSaD3GP6NMpJN28sZ9fc+6ThGA4HBb9PCT13ZeJLu
W02Wk4eOQ0roExe8eu1LZSlywxM29qrk3WuLm/5iTypIMoQfY8ktKWWWgB+vQzW/
gqrwLSU3WbLo7z70ZpSgksSggj8MjBlhZibpPEe3qbK4SXp09uhHmoUmLjCcOLfq
j37XLeMAo/SAdqvL23tBjnq9uMmnz8qPF2V4+Hs9aBkEeLkxX2ZSrlQoHErofNfe
r67EP4ca1GbMSLVV2z5uwOM04XESTCb3ijzdPwirR4n+R2O/yoUWzbxXyhZyBEfj
QPru+H/9zPegl8xTAa/xb6tFAqeKErjz/dC0acDKZg32GBPM3WJHEkOwy7sibDJH
FxN3U9aYORKeeDsgHxcDqdEu4vkGvOBO+UGUzm6JrygnLKYGu605j39cAgzYAxQ2
ZoAMwlxKDiyPyyJUpXIDUsbVU4320xe0S+OVLSmraGuwYg2XT7TiPyeExGuctC3K
286+1B9kjhVBD7f8piRPJCbIS2nFWCBP+lNXjrQyJ8ydGhBOoowlvODiDI+Fbh+x
m6FjOrydCmslFPui+3eHDZiCCfPAPD5Oo78JYPOdduEUn/sB5YxM8ecfRjW7xNKz
mvagdzaB+HvFKNYDj88pjEWNt7gTMW1Agb+rOESuq8WxSOqGbJkzFDvVF/v7O2WH
tM/YzeQlSWETk46E74b9BNggpNnehbvRLa3NX6Aljiwp2J2604gjv0PZd9ICBz+y
ri9uIQtd/oSp7eOgOrSIkq8+eNYn8CLTXPh7Ie0asVCqY486Q+cOHyUSSHA+XgA+
8FPPcZgf66b7xy0/4+iSmmrKBI6qrJhrdG1ttKL2pc8BUSPcOXowaZN7AWi9tQLb
iidtrLn6VguP5qjiFD/jn1HfWY2Pm7fGmfJ48BzxN9e1AedrLVVW2EagEkAavyUD
JoQ5jgZzdl+Boq0vgIFJhZXKyqvaR0u1g6+0pbO/XgvAna4EssNJw1NwetIGNX/s
E4X9eJ7CUHbfOCyVttmUFJDeTC2ABYzILwmfn0oGaq4qg9xJSJ2G8QfphHp2caQx
htcI1bg5EEYb0GtPYqlz9Dqr8EyJ2J3TudwMNY3zQZPtzI/f6OR/bBvanovT80bj
5G1YshyHgAAtozg6RotuGYNo8utGAs5Kyv3C7xMrnw8s4I56ueLAdtqcxsvEQeQs
MSIWHkNQs9TOV7/RjM7guPfp2LFwc0OoVM8SNK5btt4wvQmoaINx7jo8D7e4VfzN
HsETWrFQIQljDh7tfVDVx5CePbcwTFDEbg332ayAxpEzab/Dfy3e3KvjnEidR+qG
L7oO5HwKlymH62Blme5gLazBO7mDhBjd8okwMGuVKOs9QKUUWXKyy3oQymLW+iFv
Kin1soocF5JIMNjk4rZVClnPCFVQz80Q1hTviKe0yHg+ajkfdGSs+MjbbFjXyg0e
HJVqN3/jdfWdVPo5Z6RoCGrdrzY23KjytPjTQwUVBFgxaHUjhAD/tSH1K9Vu96fB
QWoOxEjTuHOuCu6tGVKWXmDPralF+ODwdRnBUVp78sRwGeX+j88zbFRfVKyr4NXu
xwzlPcrKC2Kuz8fysJOTLxTPOF2xiRGNPr42eQFqVTjyNP/x4Zh3Daiq2y4nxR7q
2bC4aj8joegLNcEYleDONpbrUKO6AO2idwswA8QnxfXwHEaBUF5S7cAoCAt15nEW
HsAdWQzY5jYrdZC6PZYnsBsQU6crAgZlSwCmc/Wn2V4z7jlvnertUBDBvMQNa8xI
Aj3dkiqTroXEfw0/SsZ4Zd8iC9i1MXnllsiFUvalMnyiV/VOUEnqmzLzx1S+VZuY
EMHOXQM0IfUEyl8MhsaAXAKSpkjlTUBT4sx3XeRA9JhFhGFwLLz+pnWuObg9CnsD
ItkYZrF/kCzdW0BjYYP70AdDC3XEC4lJku/Uw8AXjSIsLumbTntZMcjx3ZnQqned
EfpcdmkOOnbwX4o/wfxcv642R0AclaBHwNlljuAIGqKVtXDp3KCNm/ayOdKXFQg4
K0TkePirZeVphpJIl45KpcjhdvchMocTmcSIn5/YO+KZZtr+Uq6O4NiXoqubCp0P
9cfm9B1l1Ln/AklwOj1jVeR7tqk0bFdkZi68v1iWKMHSQmGJaXw0CtBqsWIzZ0YB
WyLcvaqtkaBbI+YVDZno0p7VLO5kCLcr+lB8PeZXXJJJ90EINH7wmI4jlQP5yVHZ
0s+bYJBDr5I9VvdEI6iOtWa9GULMzERLmGxmtwevfVAaODDdQp7ZB5kSe/R/rVum
6fWVbbhTj8hxZ3iKNygo1N3jDeGzgnodQxgvcUpfi377VLBtJDPHMg9A77FE7fBl
JleOjkldt3X7vS+XcdbfrqkZtiyz65+xMBQU3JS3Gi8wH29Z7M37jMe7Sl6OMp0u
bZIaIDsy954B6SBiqruh4EEphGJxRkjcKp5BGMhXBK76amuwEpogadX4PhBKBH4V
UMNjIfBz2Ri2M3maFpWrFrSouxttA/sZ584t+HwDI2co/ZBGIvDQeOFN6ac7UaLV
DqgeuZY0MC9oF5sxYd7/1+x+PTR/8SSU1gwzj4sVQJL58oH6eoWj7ryHcH28As1O
jPja9X/DttcQ76krH/zR5GRVO+xuZA5J/YXGRfGP4vICr99Ynaksjgisp2xVu1XZ
HnAXx2IBUxlAhcFM/wrqDbrT/OL6nSM3Qo2Tioo1+zOy703wFtVK0Z3djFJJG3H4
U+qxDBFTJziS2qem5RftAQe7c6LrFspCmMFpzNs4UelbdqPtWBkTti/YVtcypRqt
50Fg880Weqk0x2VgfBcr4lwdW7lqRXIj8x1SLKn5yvZLmDg1pkJLtPcTxgfxXHkd
GVoFCuewSxal2MHXNVt3IHj6y8/6uBt2p7ia3ZvEyOtKoTn8/BBcAG374bc0TJgi
p+vspqYDf4Skd7VqsGRTwswhUyo5AkErMzprSIlDMTjmOsz7lLogz/TS5VKX0dBW
rtDMsVC/w26iIy17alJ+4+Q3ZgbAwjzYTqjFN41SBhaPS1gZoMX3JDd+zzRKr5vp
Wzj/WYsN7E1Uy0aMUoBu7n4kjyUKkDBoKyyRvSCom/bHViDFtFjCeBOjrmz2Htly
Ock/zbZqU1f0QRpLhUTeZCrRn1iGz+bEAMuIaB86yNnGk5o9Gf13M+vPb0+mjh7w
PjWiKdBYW/ttj93fvTrDY13bTzIZ5S7dl8aAqOxWWkQUM3Qa++a9llGGXvl7VPks
cFPIPFknbcxquG1McqdN3epZMwfNaUq9q6Ob90OX711RbuPxQNSHVFQu2sn6b5kz
MsHXpdURxqJ/M3w/gWL5DkMqBJF+99dydvvoU2Z5Vgf3nyTD0jfp5GSnuFyS0Ll0
/rcs338xkeSRrAPcfcEJembSJqVm16658oBo8gUaf7PJt2AMvK0bgI3SyxQP4Pgl
yx3qIqdafwNjWCvpd+oScmOAXb0g09DMqwxDsp3LCXVAxh0CNr94/wLEcmSvkH+k
DqiD+57ztXKqTm3T3IHfeO8dpsBA1t0VZS5PBTH0qmoyiZc4RZDMYs4K42dLGr9/
efiTwUkYdqfwKt1toECG4XhjQQJrBv5yCzR2Ab8Lqkmh4p/CVUONYvyl/UC255uD
6edKnKMPjKxqeLgaHVKQIHiBpRNkBFjq+ZIoWStvcB64GzmP9hKUqjspM13z31fc
82bPanfGg+MhteXgb9tyeicrz88J5atV7bThR9olrJGN+JSxwOnv1No0EC4tmZLW
bc1WpAc+Tg9baz8LAeQsTF3NMF/5WrcjD+ua4EXm+lnqjPQKtBtLtHrHCpRGvemb
HQvOMffgHmyS++rhXMV9GSJaki6Bvp4QDYJrcMDVS18U2Ok0Z95n5dvTxKXk6I4B
HKWeVA1wGSA2m2GsZ3sE7ufssXQNOk0TVS6TYzaC38W0pNCpxIf6a5ECHGOpJewi
5AVjsshB09moO6DIaSNorHIebWmodOuE9fWHkOO9tHEtp13sRAbV1Il1evJAU8mx
NPN7Vf7AE1NsLH2r6aHS9t8JaT0Sy1N6whGb2ONvJH8aTI12FLMi1fomjOHn1Ejf
NOJ0dLAsZwTpBFIlv1G5o+NHWHzXoQCUe0iI3iG323HAdxCw/ATTsl3SQsmoREDn
tuSiNQwBES8/09Ht10psGq9ZbUXLo8Cuca/wjOUTWd6Hmc0BBOe51wbn5Bw9jMI6
CTJK9bPigWSqArBPfSSyNrXDB/aIBjwIp2AMdnwPXITehOMDVo+TIDAGsGNMj+8Q
1QMBF19Nd6q66sgjWb3mSsuTNGSHkPnJiBOfPBY8xtI1yNk9rJpp4Gz0Q5zmdrap
J1IYRDpBx6LV9uIUgxxRLRP794cUrdcj2k5TCflPym12t70K5jRNd+zsDKAl1cVF
uZK1Hagma3qyH66W5TfL4W7nqJFroIP0M0z/03Whp5XZf2Xu54aKDCx3nwfiEdjO
rykLN8wFXtmiYwrPEP4ZxVU34071/4oCgOHYdtP3ocNhUn0fPqyAJd2u++/CcgUO
Yu7fGaF3OzO40HYCX3GgV9c82cBUv71IIjrSqoDmdfDsQEfzBSVGogMUV379OBoS
Xv6G4EjM/sOoYqdmFOaLhRiO7oaJOuC6i1SSsI/BgMP6l6wQaNYJCwt4thu3/E7v
WmgUtmK1fJAT6x6EG5DJskUh0sU2qwWTkxbsstjO52c90V4w2pLyJTzGmM/ur1N/
0mzo/JWPA7SgKkH5uwoacGcvERy+8FKqLOCuJIiXEWi275sZevWx+DF7CxZ60fZx
2qvscSKwxFyjMZbzP0WZh7zfLaBcaDJX9d/DoGpjwqU07Ze/3pD27W84iFxlsZao
I4sb5p1sSvttQUe4MwwtBa8E448s6Ewbj4Hy+AXRQ29HBsoJC6VxaNMcltXjn9+2
Kb0jiA0mY0bAFZ1ByoT3PZO2R/cTca17wbHIdkFoVg5XS0A2y1kyOsSckTvo5TPI
Efug9r/VqjL6Rv+qdMFHOl91AAIFLzOfggbv2P+4fzClibkVZhUHtqcFmTQK6GPb
zJjCGpwGb0deBOZDdwvumbUolACcNfgUHsUUuJZns20K1EC9CUIHlj6MrYD0Ee5n
nitXGABfWC928vsqIa3buWGkSR8hk/+/ZV7MMERZoXNH4fXU2Tj3/ictXASRLsfE
Kw86OvHnOY1hhRgSgEkXmaO/zfUzzC42a1XT+Stlqe0Ah3+ZOUdj5tgsMZtDpzpK
eHs3o+CVb9X6Ajlq/9LGf7L1uWsvi54IuId18h9thcS0OMCSDckZVjPDMbvia6E3
PqyFpEGQBvdJfK+3OnzUeQzXcL2/o/wdqya4nauYBuBGjph+8Cb9xFjU0LjgaqeP
blH2Q/zjYp0gFa4Dm0eGPlnHYm+41eVsUPHPFjcsuTFsyVShGzhssy+5q2KrXPzt
MEL0M/njKDciOE4bb/7Yoahis9W6yHN0PgNEY666EY+0WWcrdReqxgIBY8vXGCsH
wNLEExUTGrrA8wWGpRd8d9kIfXQ6G5ab3XsU/YIktWTyKQBe2V6v35zR4KUO5fp0
ezE7IEkehpODXgbO6tiN9KGvy6pJxd06UlQXHPHRIW3lrsZ7mKOgBys+Fq7lM0p1
/tRCSuWjsltL+SWnlSl6erxRyFnnH7e9G2c6eILKMqqWyq5ftQ8KSThfodFGY15k
ULHCYk40phizi8lkhrEH9GylY0C1cuE4L6ULQCIQ6FQZlSMlACsL3wyzXiU4KdK2
2Px1WLIptq/8Lwm3PTmfa/ec/qzJlGrwVB1JlCOQ4jq7jC8Y//n6Rj2nZUkZ0IuA
OMJaTtPDXwyQN61PA9YqR0OQq0gYOh5kktIxaeFRgcSB4KsNdXMdMN8mtE6fe9z4
29Y6GTGEt+9O6nQ8Omv1Pa8bmGb8U5Vg6ZjuVdp2zzqBYAV8qWZI7dKywj8ZEmkH
yDpE2Ox9BbabQDGRI4K3jAvEOeSnTELIDvOP9VoDLhDcT7v1cya3y0H5gyQGALrs
7KnCf3nC6OmIe3Aasi2n5GS8HRb4lh4A4pvVaAPDJhF99/Q6jrn4oD13Fbzt2074
EjNphXoFKfiK/NeT9TA0hBrX1ZnHYhr8Yg8PeCAH1d8oyicqNx68OWfPLQP6UA4l
635OF968G4PwZ7H8U5PqFjB+8UsQ6z//EMec77MsEn2o6RSQhqHl2QPkXxjtNHYW
fPupQC9lN11cAxWPK9hR2eUs70llNGXVmxOOdQmiQS38kg47XKMnI7LwiLjtq0AC
R7iPfAPgKJrmDlKhqlgOwHmgb3QqY7+rZ5CJtIBdqj/jrFLVzT4sVUDtiw+T6bow
cbZgiVt9Eyz8zBLV44BMPRc03lLaVrPTMQbopfM2GGU//4kYBzSIxlS/T9bANdBr
3e6F34NYHh5zRDtwCN1tW3AtGjVhJpdLDep7LfmkiM6eWbUZMHMX+OON5Z98NX15
Mho1K6PBz8dZRTsyVoj7Dp6bOzEH38b3y35VaYrxtw85KyeftVWS7hKfR2MzHyoH
SmGm7T9Y/O4JVROqmyjVvXlmAdMKzALkctY0pJg+AwCqmRJw3Apc8XNoANczFn0D
KK35sOD2ryTYy7H3uIhAY469G+Nyr87Lt1ytChXYUKlJzrb8Fotp5EDuwCeROHea
+GSSerKREAtKpPHqDnjorZ2Vrru4tU6U6dV0SPSpkK/fB+wZUfQWe6EpUUiGAekp
9UhZe6XLuCUscRFYsl/FBRb2BnrNVvIGb1/+lAdQDt4FQv77RUZWu+iPDNB8Uknu
pFAnvvqxaK3X8BJWfuYzEGUPxlOsp4qtAU5+bEjlyo51HWtA+U4cC+Tzoo34hokr
5JkBa/IrAn940uZNIz3LJOS6ttYPvQXs9gaCvKVRJyAIRtYLnoHh5ZiMI88RIzWi
ZfVnRf4RuDiJcMt5Yhqs7g4nTA4N+qKgoP5Rc8/qLpDMEpZq5CpvW2bboida9dJ+
nhU2v0i3p+Msk05GkknncjqgE48o9DpUXg0m1JphUTj9CS+ncR6pcz6dy3ZO/36/
RbUJjsRQLs4z/Du7oIgDGVK08doRQaB88Oi2Ae69o6W3LbkfcVosqgDWK34nhDyg
hR0deKX5HR51FAcMw8F/id35nu+Jt1Z/S+BGTXDUx70W4EgtgPSwo5W5ILOz1+CA
WbBa3gcRq1/tK9WEAhpA1QdJps8HzzCqsUMaf/WWuHIhCyKpFcdl2KpvFlBdxbdj
oh2w+Ljbv2fpxF7T5oHf1ruEkFi0IgB5ydFlSuPC3OdtTtFoIlZAzXI6nUmGkTF5
GpGVa0GjMeCSSNa7PMMxeX+MBeTbE2MGxtkzf/30ZYVXF1LZ3FKvw/hZ0UTQtKve
WRt/z3KdSc7fpZViq8pPVUuIBBKBvR40bXWd7wWwZA4+hJRJdcre2DtsD09dTWTz
9ATPqUDDAxnvld/EPzC+xkogY3XyAwecyqbYaHfp2JQg3B1aOdrlOqZyJw24h0aq
26WGm3IuaLHBXfXLgKKlM4w8dvX/61SOQf5cojy4Rp1A0OBPOhaS0pke3AfvjZP8
ths8OIpA58y2zPLRZ3KypMLsL32nNXjq7WIwpKpKRAZwAIzIKdz7AGrot5Kd+B1T
S/OEKAAU4qZiiAR3dF/QiCTPROIQGBcpGiRHiCZG9yoQHE66ntzpJ0pMW5q4NqEi
8oaRl+/gLV6dC750JnHH5TzvFeumub4mvNv83fQg+JkNU7duekrKR4c0CaftIcyN
+TpDKFhzOIq7BDv5IvdEf+5hNn4BHheWHx4EYCmvTry4MbQcFoGmOW7qIca64GHO
6ATFH8wFxupiC4klzmC025sFEU2c9fKeNdAlAeAzwdVw4tzGeZtVuWMR2OHOOa6G
39KMfI80Q9uU8my02Dm/YiQb/7XhsEHX6fWOJ57LqCjzfh7ug0zAZZ4u9xBeY4wv
+Scx0tIEEM1cKtbXD5KPgZZpaa8nf1yHgzaPoIz2sHO48Zvq3sYIUXa7iDxozfhm
rGk7sn+MZ84KETqsM9VN2VOCQDvlSN2lxYTLgibOTz2Npt7ZiDlbqg14ZGzooWB/
+41PgHHAGPTkwcH7FjZa3AiEo9cRRDrnFDzZh4AxeUabgFpudfZWsn9rVV9hTBUd
4iARLkW9laobcoPq94XursfyYwBY/S4d/8Xg0q2lFXksqxKfBhmuxc67l1OedwFm
0+k+DuIprJjY00caVqq1UPThbHjqops+rVy3HxH7QOKYYCPcJjEjHdmVx75OYNLX
FG3J8XTcZR2A6urQETZH/C/9zpnZH/zRxou/cs1ICtSmCz6LIwGmSjhoNl9xAQ/j
T684VlSL/O/8OE8dVa3mx81PS651q8fQdUXte2khR2edxbr0KWBqZ7vRgwHFgDq+
5qWTJyGPbRduaYcvwy+AlU8ucIQbry1DgZFibvrLsVmTiInay9mCPCzjBMVxFKVE
DYpNERLMVsq/xZ6JC8aQ9lC68G9I+hMYFi+nEmy6/nwxdVYgyYQ5bmcMkOgj+qAe
Ywe3G6ZhPJeofNoOcUkIpdwDEQfaPRXeyS7b2YmZ5yKPfAa4lieUF5q6POiiJOhq
BDPrLAyaLkIblSfO3zGkHfkqg0o5n+PYjiBqHjoszpcbhpAMi/r5YbwPBvL45R8d
i5FTW0QhGkAiZd2ZowgicN+/dIZGhVwwiJJOsHPyVYDJdVZ3DiBuFeGVWGkGMir/
TQJeC5ovK7D3789/ul2JrhnP/jogLR4Q2KvVV7zN4HUMCDuHyyCzidvvmGzfX345
VpDB88qbGezTWJcYLOCuyw99pt0+DMXyVe2HvZxeRu6NCcSI2bi+C5FQi8U8lLAf
UqPf35ThEFtuDTucmoaHvQmef7hqU+PBZO2jgXcwedeuZ7Pru8ZlebcmY6Z/ql3q
MPIyDEmHecKWyl5u3u7dDTHCNoVjePoabk+vzw8ihTm1zspXXBPs0SqA/ieqNa6r
9hGyCxs+KdNsTZpaCYYc9bzPK3Dsj9YAGQrY6yLLivFL9Zd5c3sNsKHKTPA5Xb0V
1cm71pQZfDpjVthtmDoVMlvB7AbUCg+FGobdb6cruMa3Dc/OnGOag+4QwTEcbpt+
YehD3jB2DtSHO/O2Lncd4FQy0eoOZzlCqRAPRsJ43hx766QSixKrOKPhPJBTi1i5
CqAQZNtR7KQOV/Jkq/HX2rijDqvTOwaSseLVnSNualQUSycrZjlvamnQxhzIJEYp
l4qKWj6X/2z/OiH+hXdW060TODfE+Mj3+woZauLS4hsc/KZo1eD0CIXgEPD3k/1c
U7gqKS7gYdBGJWXdQFhOjzL6/Eprou3CeHUUSBBBXTIKilHXCfAixlyc3Nso9dpz
bTRldAw/JBqoGIh671ue8hv5+qU2MGPvpKScjRAnjwzYvqWtXMKbFGvtLMxKrwu9
1frtX2/OAvRUmv8owgOuBGlwK2lM5KhnBHosk8JFmFNA+UkrvnTY2Hasvlmt13+g
OJWRlfwyb83NIzZFCpBWv/JvIa+ko5id1gjQvsVRqMhrioK82EMb9J2JqBe80pDS
7cdgdL4I3d88XaPOoI7zI+EN6+14RwT5vpRGi3bGHI+y+wPow8nxnTHhGGijOIBj
tjLgdEXU2B7MNUY61PLrewS6cJDDxNlJZioBk0eamfEToY8nYgye/lEHNU3xvS+3
177xfXhmzNa8/aja0jV1EHLw37IwwAfaGxImMQ3uHdnW1fRBSvqnGvtaSOVvxCzM
xUCSWRklrM9rBbCBxUXV46Q8FFtl/FHiQmnkHinBfwH3TMFd/db8OkJZG5vKOPUQ
cK3BdAq6pS7VWxKZ3d7eLlHBMhu+N4led4OZIu6mNnKLyfrmWbuI0VVFfSKziNzY
a+6wC0RSPk4M+x06217QlTvnjD6K/lZ06ayPnFesZDkAanTxhfCmQ6Dk9pVfn1W1
mqcnk+n2k6KKYT/L+fs+RO8JNjftHwta6t4RQrGsezZt8CT/tl5wUy+e4h/hMiTc
YvOwjPUaNNxllYOOHWigUSSAgOYy6avKTZbqSuwJYCRFFf5doYgAfgZv2keG6Qoh
qkXGEqcpYQzPg1Zcy/I4cl5XiZ+udqe7HiZEkQ8MEq7OiAMfjpW7VKvTJRZgUI7i
CKG4y/NKwRCH2mEq30nnxPji8pZx+yAMJN66rUbn/I9u4/0fKYHkswVs2wlyDpjA
4O1H0ivFEMQba3QIyXM8ubYm/TQnD6vrWf/stewG3uq9V1GF+hgcgVUKl2ywo9GQ
UOCEFd9r75s5ADm1AH1X10cx9tJpl+im+I29G0mwb5suREpzdoH3FnxsVaSfSh4C
A+iXqedvziNIY1ZxMcFPoFnhAeoJWFrrTLVQISdMGwFehkU6IpkQfRHuD7apnzZf
NaSx/1Jk+pcx4qAMoClvdxK42VPR8xQdsVD+77R/LveVZhvScqo2cUcDKDMUxfF0
bR2Ll5m+JMvMbXzqqVzj3j+BZ7ng2ZFq0vdz8qqLf0Ag/+2iG8HYFQB/EBwhUNvU
ePCDkHFQifvusW8W8VAXXb6BVBAP1Is+GIGStXZyXlJU66bILl6hQsu7hjZt27be
BQRNFRp/qhUqxgqjPVtjR0rddqkDlKzYymF6tm/nLVnyvEWkJkY8kacWyrYSxS1e
CcxSRvkZFROPkSFlXVqnb+cqnMGPGBc6kM8DER59mIVFY7qNJgIXBsYuruqhE7ai
lXvHeKEmBoPTb6YU1MwtewjUfQIMlwAFNYwHFxUx/obdCC9NJEvK651QzGZrgIPT
1x6yohCaOOIdMfDtg54udSZ325wxkJFPDAZ95oZpBKVt1gahuArThgcGI24/agc1
34fe/V+o1iKV0vu5jPNQIfaz7F74/fz9BzxTNjQyfe1Ah9QwgolvsZwfI7YjieCa
zcnl7XTcPf+4Nq3rxCGQijtdhW1RNxK00Tny3luKAG89/LUnmN/kFOOrU6tVyXnJ
UZaP/ZrYkuxSpunYRFKv9xID14Osa3+BXRbKDY+BxgGE6oxZtrOZroxguEkSalDD
q1951DyhvweVXpEeV1CM7SEIxuvHx1d9nH3wmSYL8a+nZLD5goCEYLyMKtLAlB22
AcwhcTtJtx5kA7POMUsgCl/+PWiP4cvBVMmcHIwzhDPBCgj7aUMibiaYYtS6y6Or
9B+YGj7iheV7mLi8zqSLTUsRuE73vEe4NWIJC0zrNSMNNBjvtlKm7AoVHGoCmqU4
Q7Ox1XiA+uwbJhh44wBouNTyd7wgnUdh5ulEHXUmwNV9Z6CNS9fl0z7TiYqTi/8b
C99HqcrmictaS6PGBLCCJsCO7Sy16e/LF0/0aJv47YCh7HEfscla+VS+mOWS9X3A
WELfTVQjcCGoySq7A0n9Rw7A/Y8ue5S9HKui9OHYhTmLvag8gVx+YJGSZbva1P1R
TImh2UzTklbglmngC9gC1LG//Cvo0WSepMQvYIdQ3VlyL/N4ZrEwVGeFUnIc8hvC
UbkNFgIMM6iOnRu1J71bHp0ziKjntOyQl4y2KGWeOL8fRv9fnWD+KZfeY7wSBk2H
Fj98/vnlQ5MtdjEGQIMgaxKS9oHy7KjZl9jQD8r1qiEYi3vyK+bSg25+an/xVq9w
e+V4FWQg5ashpDmnL2KhrEAqYD0DaFE4Ixrz+cney0zJJG9TfTvLlsFk4vwZjQW2
KGjmYt8kj/IH/bVKzvl+8OA//3htH68jaupXYewO3TOd6oJZfY/l7xfrrOx/0VKJ
M0Xgr6wefulSiVQlocL7uO2eOmxvqDqCe2JOGLzix/BYlpzfXlhjKN/MK4CmRcjL
JoI20csUysBhBGsuFP2e6V6vp9yhEcBUxJeVfdyCue2nvXdWoD8GIfZWIrpWrXN7
NxvKT1KjrzI5Zq9vPSv6rj7n6F0sHtsm0U247gWosqSyCfdgYJvTS5pWsz0lPscb
BbT0rls7tgbXD4EYrRNwhJZUiFEXhk/X73NpEi3Ue+Eq3qLzDKlEyhuQx6PIceRb
nMvMStV/drGJPBBr19tNTRdZ2G6WrJrt7zfV9qTQLvBCGsanblMIvG23kRDJSbOv
GVFSr+JxCDG7Hq6tVTQyTHn8edvVkjoBNCl2Wtmh51Enk/4w5ELLs9FGQXPi6uio
tUxZQ9mhmasQ70k66Qb5l9ALghLT6WITZf+3rVsX7+0+gRI/h/5Cj8xil1+JQpSS
8WXmDThit7qnlSchOM24acIhn7VjKVrI2yDK1rSpGH9sH42ZLBn3At9swU6zRSO+
c38EYOogF+FRqAUWy91BM+ZR9C+xjA57ZoeMfOsq6VwlKf6yKuwD1YBmjp9KMVIJ
YXtzQEfXqr/5RN7pKWHn7qgaQkg1T3rx0lM6xAIzybcDACsyUoAzeNDRxBr2x0Iq
elRQE4Q8ncMz1J+c5xSePq8prsm8xqLsWNxmj0JSugEvb5g56Toj8/dlcTa94yiv
32WCSZXTRB9yYm/nxgmz7cPayZGXTyM3fl9zUdD1b4nRiZpY8QcrD6xJJGsGmDc5
gqDEKPanpQmryPBWVysqa3pnyLNBwyOK6NrgU/9m2npnYVpjGuxB09qcaibaKdVh
N/R2e9bgURBvmVLTwQ3CT7bkL9B7X2OhjikHcfyYs4nTCP0FR/62PFp5DWYNKHXQ
ZjsYlnRtp51TmU7KMHxYrm6dRE3Kg9ZgtsZH1w++3ejnAMd0VbzJhR3ONZicYx1M
qKeW23eihzzPCP6gQ35olShzqsvZVM+WyQq4tGvA6za9fCDnMzEoBC4EOLcXDPyb
aRoUwvCV+4Ov0NgYL3t7Rk2/NQWzVXWbN+fEgcFQuzcaw9+aahU4wjnoG5UqNUBT
fC/Ejgpv6EePBhQ71iZRPNOSC1OjiP/Y0rIlx87ccOacTjIV9mDaZdbF5OwykGEx
9oR7X1NEaBbxhwrhJjN3a6BAmXGerd+aeKFYD37lyKvgaYA0GODVVfRhCFUIjnaG
B1ZbFNYSpsI5nU5XNgWI8BfHLmxigNFsvTSyG4Cp2LLKZHXAEB7g5qh769iEhU17
WCiLEgBY2Oq+NVpXgCfTGzUNzEOTg/s/T8mJwAHNriu0eG4ktb8KV/mJJwJ7N8jq
2dxp63YrfbllQvuIkBN9MwxloiqSmGfRbIx60AglUPhbrh47bcq+I4UCFEYWNKxf
Jn/I0hpg5vjNbNmeFwpsQ3uMRN8D4ayTuRKtl46U0zu4aXkXYuZ3dcQvgGi48GjL
s0ZKpfomgfueKFvhZcfBO/QDpfucYYlt4EvXIuSeAgAVjxAgRWVe7QFinvq3f2OY
avyB0ZS4wpHypEdw2lH8CeENs496iNmtcOehBBgm+n3tBX1jy5QR8pVpbgagWyIT
I/SkFC5FhETirD+N6+5B6ermUPqBk/KRKw/R82aOWtCpnVECOfamADwstsTQrhxy
mIDS9muyGnvK7TSWdRuS91wL/huO6Xn77A0gcSYdUENg44/33TfhGjDZxqz8C5VT
V7a0G+FmqaJdqsJUzmLiTEnRpDkqqMB/nATUJ+E86n09/R9evO6gLNZ9Ws4f2lRT
QH/E6ZGmiHB2t+15FbGpWuRIGXDQQVQZIPOjfLQMj3X5VVjPL9qLJ3fzV9g7SOpE
QddC9vf0V1aukjfsGTTvTDhWXkRlYL7nGo8oE8zR4btk80YNNMaa/R17SaAFI3SQ
n5Knhlag+hAxKGoKAbB6+gYvd2ja2GYxUBZRnNIv1RPJzRWhAOj7CefzWZ+WhrDC
1Pb5pWvS1WVCbY5h7SJDPFMZaBh8NyVuhVqGBLe7WllGT4WPFaijabSILYDABsXv
BzL+c4ZgSwr/7b58Sp8D67W9omG9VFKnb4d5+L+JyPpysEap9yKLTgVlM/ra1gDo
GZAMCXF7vcbYtgFxHfiy7ELDGRGfwxZhyAorwR3YVUDPv5TdcvFEia7sC2NsOH04
I3qhzu3Ha1uVpEbDYTfYO1L/EGbIaOXlHftJz6P3RkxsM8AgisUTCWIBZ+3b/lLA
Fa1R8iZrGRfOOK0h7Y8wrGkIlCPSeRUGOVFQiUx+sG157n06Ppxyxhij/XNcz1Ur
UUFxEjTaeNv7nWzlt2CyhphDXtfO0HvXpCM5BOxPUbHlvpkQ3zdf1scdJXRmDmDS
T9pvPy85/px84Gw6gbfb2S3ASkOtC9ftM6b+Gls6i8/2kfTPtp2TAoP/l5o4eMFV
fw3xYO+xTUKmcFli0MHXrMRQHcHMSt6eGCMWqODeOCLUM8tYU5I9uY+F7av5IkAw
LcEToWZhwyh9VA1VjXKomi+SMm36vyRDpqSB93zDtwjdS4c3e1oof3UaTattrII7
vrQq/+WDhoNQ2l1ZF1el4QzzPFwXjvkzjbY8HKxrdWItCHH04sk5yGGxHpdFCyQd
RCKC4hE2Klx3tyfdVb94dATrgnQnRN9ftsXfr/4r5jpQIahwjE0cvAamKOLMJ+oh
GvlFUPio+GC8rKPSeBQjalOC7q0n4+DVRCgb96HkL3CAzgGvKNWjV8QIHFEFTc2v
KZtJXsFykeVpFWeTusZoPhTl5MNwIcvdbDEQyFse5Ijq+xhEi0IAEUi4Byo223SB
v9tzQdRD7w8WtjVh3sLCnb731vnaDi9CdNpBw0x64fqVyv8nxwj7tGKotXU3yN1b
nW7XnPmM8VVNvAtqN/5xmXFkGj9hBIXmj1+MQTSScYw11rWleNQeILD6JRFr8Jm2
A+4xiyACvNe+8DsoaLSR6v9Y0I0nmYwfR1SAoTpDTGt/Yrn4YK0dMec3Oy9Ji/m3
G51RrFPZzLgnX0SSa6vL5jObRfWblEA8+j19JB6WMaRJ9z/bBejjWpubqDE9T7Qk
09EpZ++ivUqksODrMCz6bEEjdr83zJkCZ9o8OxkRMLSpfWSJoxbKxRJGLJmE1e5O
PmGIeSlkyCt0BfsDwxIROtWF4r5hJKhOaSXiOnDvnpnUD0LJ/1RADCXa5eHUHgor
B9su4/H/mXUswYOrQ3HnTq6AgMpO1ARt6Ghj9Ny7W14kY8I8Lj9iSp8x5GpHOKzB
B50Nv5Grcg4lhBdEZ1oZdkyvQcagFoW8mqsY9YXYDMWIcF5w0+Cv4aVsmkNqgtSW
8PfGZI5Rg+3ulX6o/eLOm7L+1hb7GgztwWkbglx3m71d/z+7N4UsT8NDg6vrnZhj
AdgJhW4WkJiTbCIgNWi/nuKy8xscvGu2pc3oglIw7ARiyXB4oAecD0YLBWRFVAdY
5Ig5MQakbSsk6pfLOhFFAEL3l+4bSH4UgCO3n3XVppcl94o1HMQpPWJVA1GoQV6n
Q0UbVNU+o6gOMkFx7nfWmZ+F3uc8Ou07uqBm2FN+bzUCFVHdvLh+xhG0KsCv4Ybs
wrtC6sXA5N0sQhtwkIIFEOqpRu4wbvzo81hCSl5YZyfWKmj3/PrPDkcl+/KhP02N
KjyLQFi5Z++SQeafBdhQqWQ72DO1a4eWcVmiRjXChP3t7VgazcjvjFC1lH6pUFBf
xP0kNQWboooZsQu+Y0L6Gfwy864DjfUW2irAPK3CRtIgG5c5V+H8JGIBWzeFVlOu
yAjrWbA4VmhvOse3xDDNum7gqx2yFNZR8PS4geN8FV1yoBPbU3x4UbQeunFae2PI
kC+HdNxePGY1ndPfRN/5ksP7/e10DWJeT9ZpVnqZQSL+T0+xUA5IkkPoDryzIy6v
WIaHgwJsDoGS6g1VEcAlsGP8DztNpdH5FzpcvOd3AUJFLpzyJlNZvYp5afkdc69Q
0C8Ff4ZDtPNsPTVatcbsGsQMceDabeCQXfuyyp1FbMmKCo/KpK0+9BjJQ4f1e4kS
qbzM75l2KU+zkGeArCC186wfWP3cnI+gXp7aBZtqJ8OZwjVaVxNLXWzUSuLb3XMf
K+FGdHb3/QMk3po2omt5afldWKdLuGTps7xPzPOSaGkTFaq2MwxFpe2Vr28ZnCV6
p6tXOJT5oTuviT4HmN+fc0mDRLuMN5FFsbiZlNw9LS2HNDA0Arx34eqjXeQ5OXPS
hpti7F0mESzd1apFHJ89koualp9mys9809zpe1MDc8VrXdxCrKOIxcgTqa1uRmk/
roPEfZ9xYfP5HMvOF3xqBZsudHk+1I2TU+KDgnaD24IhbaK3XSik4XS49Ea9PQLx
hjPEshR+W65lrYgFwtcO0/G77AND+ijbCU6rQWo9wANivxpGDJkCBG/hTVkCvbDw
179qu8gWfUTw82bOb4HclRxKOGP1ODz969SNtun8vlxTmR+8vQ91Oadg+MNIoxZ6
emUOVnbGtaYdEDESNTmmNrdS6X+dqq8D9LLtgm7mQCWp+vsO9EuzwfCmtAWwFXpp
eBH3zgb4ctwcUv0Abe+kBFntetHiV9eedRbC6KeR3+h7EipNMX0HmukcmkvJTSp7
HNY8yPbtVOkLTd+cu16tQVGEsIHAoVE9voWzZKQHa9tDyvLnd4hwW7BZ7DHJl5rX
N+f4+Kdqp9Vainmqw9iIiMET8fRjOLNqcpFv+YD+TNzpgHTq58jOV93zWi8KtvKv
rG93K/3JpWtKH6xHqxn1ZqFtbsZTJoYg/aNV7ZH0xQ2Fw9Ta/6GxIwZ++pfMjQ/V
18a8YkoHQeB3dcyyNxLlsEuS96MqzYPCJjjsxf6UtfwOfiSqPBLvXr4/PyWtmmNg
Ps9m1QnFWMA7AvQsvIYw5hSP5aRJBL4WOxqsf+kqOqrTP2MR4mgTzZQr7S8rpkyE
4Vljk9ZpxpqGS8LIZHqCH5OLfy/wD0FAmcvbETp9E8g3dWOQzxl76vAhVEZvUXyD
rvcum+VrX3Rieu+HotScSXvvkQn2ioKr1nqrMj130z1WV9j03BlfQqkaxlUP87Am
NtPX32bniVE9EvkSWJAYJl3s3eEx32j+OGgySK4C/0RAC0d6zEBLQPHydTMGG8vF
t+/NaTzf6PB5z03wv8D7nCdGpd2hbjdf0xd8Jr1UZDEe3tne6k26TQJI/mM6OgVa
SE2haVFcd9Kv6DoENi08ITvQW8nyiHAPx/nIgZkMxW1PoCiE4veagdsW6WV/seZW
9Lv6Gf2ag1jCY3O4z4f3nfEUrveM0oIwk5EW42iLdRdmbymUzlmP23LDXSwz1NhI
gg1rnCZsh68C2YGLrsmdSAs7kn66D7bwhuGj07cDEOui9ZZgGnnRULxW/drgPMK/
ESWOG7b2PbSsi9Mqq+9MtykIuY59GeQp4ROuLOJgXNJ9wMLHZKMg01i/b6cIHaJA
0YiZBkGAZ1zXPKiMKJJzTyAiXc6dXR5UlpM5ornSDnxi6EVEnY/GeQk8iyYopE5x
p4jg/V9hyp0YpO35mnZMBLJM1qvn0HQ3b0llyIzJ/Iw027htrcq+YNuGz133/aZe
bxKQe4Ua6+H12uN3fSbmu+SmgarCRsk2Pn6hQSDTAQAEGqvEosck4DHjKwrB5MrF
1cAvJ1/Vn0d8HKcgyTMtHejeOHWeMV/eE/R7g8DBnRlLo4kwxYxbwKjHl1r6WQ/u
9LArQfn2I9ED3zY3Jdtcb1QWhhK4oGUhnT2ja4hsft8GmA43+fuGvasI5ReNvpC/
C6FWOTNLTWJGEardiV3M+OspGAQxssjOZapRX83qxooJYLOxOqWJ00lrmWrRV3fv
AppaSBTt8OY7FSJBnhowk6AoUmKn17QB0rsER3XG/Q1xKZ9nEtvpn8E/2WEatUvh
SKZybYA2MDjq8uLM325dN+CW5mM7i/S+jvzqu7vdSZeRorZ1f+ChnzSYPDdRfAfw
BetdvGbEWlE68IgZhLwJVNj+FiNyPbfSs4q1+BhmeHCrcee5U5/eWaqpvtV5HUZO
+c4sebtgN2dlWFLS+5061jwNzbufYynVBpyHr1nPIVDMuE0sc3D5gDht+fiHiZ2J
rs7rlSJMk+Yu4c1BWhoqRkqEtO8oGx+CRPXPK1VmqKf8W2L/5/7gfJTRYSb2DKEL
3Em6iLpD0fMEKuTrayJvKaP74hFEisBBnrxZC3aq/sYBE6B+W3o6xLrcoI2jGRSQ
t+w/MPg7oRs6u3MtcI5qakF7hBxoPaPZcZu2T8W8wlBVa3TTmO24eHscBK/H+z1E
5OCUyhW9X4qQ1Ss1d97UWgpb3xWqAl4fCxWRL7xsQ2dvnIxww77iWrS8Jewpga+G
B/+e7Kdf8NDJvlARNQnX31pv7VD7b59453fr0gUkljaP0RD5Cw7QGkE86GMjDa1v
+EYR1gtVGO9fpicl7Bas4ZwYBFmlIrZP7GBQDCXFTmuDh0w5ZvWObKB3M1o+uuE2
VtaNZc45ABUYf3mkWJuYhVePQ+nk1rygniZ/nLohUk9if1wsUHgh5HsIPRtp3dSV
hkJcAa3KNj7Has4K0RX0VhpOCnPUaGEHXFTs8c6wxcufsVWdabJYnJe+Jf2B2DOW
b7y/WcQ74lS5tVemxIW9/TdprpjCrvhJJm6rI7QgPNtk4O1Vqq/z0wfP7oYeDQk4
LartgyQWpvRnwDb/t6r+hTBtT1qSXzZdOd83dqW9vYWhqk0WR71yIYar7731ovaV
DVtP20UpM+FQ1e6PLwpUqj077OXpdktatXlYeMpQBdlWmhAEAPyJ50TojSXPO5lE
mtrwYf+33xRRV43muBRzAG9HGRlDuWX8AXYrih7OlBdQV0LttsrdTfVjqrdVS04c
QJdTB65IjGWYZWg9ATLdZKzsKoW9lYRqgptOJcfEcFP8EOr0Zwepn9w2PvBFkm/W
+HofU9rWH7xz1yjSCQ4qifp/kgvn9nVRrD2ao1oEw6U4NRrRWEWPe94M3x8PatPL
KzuYLbkSEbEf1HT9mgl8h3W+Th1v7nNG7hxApFwCGaMzGduEjKEFTrLwA0Isz6cS
KtdST2xPitl719+h+JdjGtJRSBzQrELuwoYDAwDgKYumIG79G17tBgXKPcf8jQOP
D+D3OCJR2nL/Fi59uUfrcXKC66Ld8gkIeTRTWYdFDHwAnSE3kexhiwURGKg46BTt
yi40v9zY3fdK4XksRxAL9osen7QjHv4KVKkvDPF8cIWVW7Kf9iSfYkMKRoqniN+i
tyOMqLYeqCmDuPuxc9S7pXN3KgGuq15Fzgd6/NsmIMl8yZH7DPuIR2MKki/hsKxv
9REp62KO6Jud+/cfSexXPX0Gag+vQcU5ypnIEaIo4xoN8OPHTTfwaSDvnfzImdt+
LEQ/zGCotBIacOm+8YiLvnPjAi7I1kpuMWPLgxudpz6pJJ7sDtaqEuLx374W0vXm
BlMOqrV1hhSY0nXv4VOF30Ki6aHAZbnuTLozs1x1FOjrkOHf9qcvicc91Haes3ji
C33p3g6MnvxQIR0lsRjoCy0FltGiw9eB4ckSpUyJbxuzzI9gj76Uy7e9q7EQMHO1
WeKFO3NcoWiD9yZ0MgSJ6zn7LOUKGcauBaCKzWbdGHODKRApNv3Cqnj1ilSTTMbs
tzbatORdQROfsQ33GvXByibHQWgi837RqhkGNTJZVlciimHBWrWFqX3zW7xUB//I
gfBA7vkrcS1Y08KQHrFKV3HvtFkkdD03Oa2AVhbZuHOXHLugsE5cBUzHR6LPWUMw
nkDRHAurS/CjkxKTWH6rRF0BSAIgHzLL2MvUOHq5l57FzA65KyYBXaVInW6ysvDN
AuKOqsegWiBbqY0wvCHKgaD6fU7UtmE0DAAFocuroo310/URW2f6d+2FTCsFiEDH
C7HuPQQPcM/knKsFsPRuckZIbeh4xW6CHJxK6mdsd9OO6L5+GPohXn3Low14rfwL
4F97T2vtyoyL/iRFpyM21aEk4x5Nh5jw5B2FQNG0oP0rInCR3AlnpN3BxVYEi50H
IgPXqizhrABlg2Ghdrf/D5ZdBcskMv/pynQDjrMLMP+nSY7NCPFCNAWDysSAwE3v
iLO21D4Zkym/7EUVGZng5UAXmnw5iVPcg4qDanpOyd+vL1etaXnKrVtcYgLoHbyj
FOg8fZwTU/w+ngphU/Xw7xqmOTNlwAtTehqOoZwwmZJevL5XSbzHBthLTP0cWC+I
lYeZFNkQZUTR9TQDgJ/+kBltLzMrAHj9+6OBY8Mec64LkqrK8cQTJXV7kKX8hqzJ
jj1Lt0nQwg6O70WdH4KnGHyWVq4JirfKvJcbE737uWrdfcNxjKpbKjRVH4kL79NC
mNAOX9M12HdpsHmGnKDoZmG08Ry4ZjqDSPOcIw1TDjhY64xc1+5LTf7YaobBuxQ3
hHyDWjeCc5jgiDsqr+i8zD1oD2iBuRAS8zONsf2MXbC1y6HLH1mS2vlwZkhkhTi6
H9E7LpC9N3w+Qd0fDu13NJQZsNOcPj70LJwjJWwLURrS6Oqi+Is9moVd1CPgm4b2
15rPpzB0bvyntRXwMHUl8rmgcr8TKs9XOTbkVee3f27ZeqCV1geF/+eq0aoa2HG6
QT0oIwlO8qU3UPw1VH9XswxayJy6ArcmIOVjVCw6pNnXbUb1uM8sVDOA4eWQSMLt
Ycf3HmBhO+2N77SUdZeHT17ib374zLTF6xw35FYRfKwsUf5m/YTyzkb7NMcPmtjj
tPZMLlzgviY6j4U4BqRiEuz7P+JGE8e1tMs6ot6Tv/TLttD/RF0xDmaPnUfaXJbo
c7PnwEPxuaj5m1zPzoZQI2Fx6Gc+qy2TGBBI5J9xmBp5urgY1M8nWBxu1O3sV1Hb
QEYev3DWV67MMGJjFLe5/myJFhmL9LiAKRdn6Q1jRy0Hc3jMxwKAPAYUIvVphcMb
fFNx7mqLVVLbD46BcNU/PHAO517Ei0qqeX1jyqcL6BVsEa0HsngKgStd/SGEUBrL
uRqNgYj++SfDP+VfBFatASeERNe9r7qlHW4i8yJQUQjzlFqx1IaDNfz1z8Dhx1aX
e+FnSnLmwG2rgptmVCNzv44N+SKyJAi9e9pFYJJnliiX2AoCB/ZqFjX9IsvoFD7l
khm2aG7H37EpkYYHEfS7qy1o+LPBXRUxCPoWbszGlUAhsQcHtelHL1NrJV35w1QN
KyIAxYJJAVt6ptqak8s/esbANPMmmH7FMKuMmw6yGzO+GPHwe0uu4xR2aQjI3Y9/
Z0jzX0h6xNmPYFJbC8jdrOXAOR/UrVHdJH88CAtED4vAEOFuGyzNqVNJB9NAHR51
s0AX8qZh55G/+6XcJlD9WYaKx3BGjvx+hRGKahL9kLYNBrC1OAl4SbjuQy32K6T+
0a+dQ4urhidXD64dao6R7t5wnq7Yah3lvHISSR69Jo4Mx5wF9sx2wwKV2wPwu6wB
ihrOPkS/riCqEBAJuYpOhjLA2JX09OjVUWZvxQV6BIn+mFgbs6zKvDfgk1Eo2WBL
mO6Z5k425vqTqQ7m4ibu2QmXFjpAP/+COSxmiUjdd3BaolnuoO3R4Cpaw0QLeck6
w80bK670TRla5gQSVsQtODGsow0gIsJd4vUQ2nz12K2B7+ZEIw7/6MaRCv5FnZkx
AGPmkDplKD0cHTfsxoUOEElbWG92QtsqLyVsXAfkFggpekUfISR85wrdU7Br+TQv
M05Vgw1HkDAYzyqinpuDpxE2sRiNHV18X4EL6GrHeAsXxHHba3JH3ZBpE93Vcwti
9N03/mt+az6erIS1qyMh8QEvMBrWvNk4fXqVkBApAmy4ZQIDy/QwtzONzl+n/sKe
wZOfGpeHEuiqkgWoMDZQib9BU1rheqzHfKRspbaIVBX2wHhonAsRyPVQRNXBYVGR
+ZE09E64QcfcTays+3/qMTfpHO4JS4vwKONcZraOZOGQkjw9M5Rd672gyQoXdn+o
EhADEFUZc7oCfUxDrQZWMxmJkJTD6umEqssJiuLa+Dst9vdYYEEnutdQsjo4079e
NC8kmp2hUsxP7wbAqTFToP5L7vd51Y9qaWimL5Q2qDvnr2wxCreOwbCN/ru1s8XA
WmoeB/LxY8KpLGi0ezGAjA2qAWvxe6sjBKXZMT6R9PFmUj0BpAX9vErhqNgzmG+O
J8f4Du37srM5BN9Y+vKFub3oFOo3IP6n5pd/CKUjk96WB3CHaYdvZ486SKF9TqkJ
DbNqStOodkGJXZ33SE1pdij/aiWCKa54EZ8CXP6CdrWopbrVZP05iuY3gKqj54zt
9mp+SVKm4TStzqL1O8L7NjkH8XSlD9dO49+37TDj2hCF4trjQnoWxFY8P4bfJiHf
ow4EkFAwWoHmLcmfXr4IMCJnZkVolTODb3pkalsMnv+xPYk8szF5vip5W9oTWJsv
Swi6JFaN4781U2jELg96YZyQ/5nWjBsB65lDDi92MubTEs4P+cxQ3FM+NgAskNAx
oxyTZZJm+VjYKKb8lJ2O5fhEX6WdCb7bdy7bNG3VYlYd6msajUAH+zkb+YmkNaH1
NKLBT4Xvl03OGuGuXqDZHGPUNhZC68yJkqB/cSqwyByCAiNXuBUkQFoeU6XST3sN
D2iV6wHYQrn8wo4zqRS8wXua8qLoKDHSQUFhuCGyWNMRlT6xqex6iuAaE7E8Yufn
lLMzjYQdV177Hsuu3avvteEMY39kPSzYdT1M7hSk9+AtdKm1NkiBpslfGtUkXzUI
846XXj11eiJ8RwoRunnPOxxpoW/6EuRZqZ0kZ+jxQcLWKVowHPfWUUsTshKN6FEQ
WTRHyAWJTzhWeGc5ohMD7Q6/vQH2WO7qb1h6Yr4BJFD+/WXiPxCNB1ZF2Wo/UIvH
wEZoO+QgVFxybAQmC1fXL41mgLgzYWMsAoDGkyTGgjwC9lcKZ1HX/+G+5pjummMT
NjV7duBPdsbzAMuGj/eNMVjyP6GTAhGNkpuJT6WV9DzmZpOgl9eP57V0Ir55aE0n
e33xQVwCmf/3hWQMipVtOTJxRB3Zp63GlS0RVym0Q3srjuykAm2jqwrikNP2lq7h
+HGB85wbi60gR67XlQz1ewOGMyNoq9Ks8ISPZh4/gJfj2vv5KxzepjL8m2rZ2WIF
kM3PsCXDXTlWDj+myzsF7FQgcv9QmWuAX94Vnb85fbc5ruaUEj1hav+BLPud1UOe
CCLskNgzqZCWhWlzw5TqoNPZ8qZLh2Y/MEONdXS859o5lSBi3HJB6cEHcs1w0VA+
M8a01+Ul58xoKCRUhbFme8MFLrPZ8V41DYheAMHU4YRH8djQdbzO0GaYID75ZPZ1
jY7gP+aO03Qj7L3U8rnHIGfXog+aDfceuUufqhR3+gFOf8az7A4o/pxOmPEaGBD8
DIP/cbPU4PJXN4mTTVOEZe1qKNTrsr/CTpOyiwIjB7debFRjPuty3bk8KfX6G8uX
iklqzXEe5WOtvgYls2PCUNcIuaScbNfoJtTkOTsR7dEyiwgu44OKYJaV6rIDj+yK
tI2uL+7ryyLocPjFq+IfxLnpaqh23TUoQbkXavF+QRl6U8D/UcWR5kcSGOxDZuqI
ionXwhcskBbk+lHFobAjTPKxMIJHSQJRWJ/10EgbV19924tcfmPibSePOOVaxQT3
ZeCQ9xXzGS21WTetwZh0osEGOtpXnuZWcNVplPHjKQQEW4K1T6CbsB4QAvZ3du6U
6VndinWkq9kd/oC663sU+aKmxmCCuQea0og2jhG9HeMDhOG4PUERau8Uc0CDvQJj
w8+71BSMNxFtTA4F+ZlPy5oyqAdqjtS5cKU3kGR2g9zQzMHk8boBDeMWm6+TR4NU
2SJmTBanoDF0mp3rh7en0dCynt/Jp5ODRCMPRBizUZo+ZeI2dK9nIAbFw8AL2rBF
hu7yrejqitsZTq0wr/wl2cnABxneKEU2yKsF8Ppc7gbgjuAngaGLCVNo9kKatVrT
IPMUjLKsbefHijrhCIlwvpssYrsw7/JExwmVo3J3hkdBI1YI84ZmEdiml69UeRZF
7yXQ0xw0u6svnA2VtHgmHliuW+BmO9fWHTzScV3slCZAj5yRsVM0SqGmVkzVxwHi
SIhICprJCZJpxqSnJg2ndKeK1Ocm3WwYvIdTTPrdd+164wskN5R4Tb+XQJhzNKfH
sjRpjHXwYNTJHV38WFaaZQxz0Hh5AvOhhjo4smo0kJcndke4cCMz5SdQxNg+IdSA
RLDrbUuUqxPk+S0k6kGUpqYJa+8NqLsYWGim/85WbZKrrUaTYApTFc1R3IVAs35e
0hEfjRznpTPJowKN5Cv4OzL0fb9D9JuyCWK4EpGn8RGBWS70vLgu/ScWGgQsvqtp
CNQqQuxgICCOuNl2nLh3m/ZgalP1KvTKFpJgS7Hu/nnmJYFJgOc/yh0MnJZgxlju
b5K4FXnNfwfBSbbXfO63toQpjH2K11kqejFmRw4PlGNfkhVWl5ckbdVdr74xXqpm
kAOiDxiMJRnGHhb4kDnl03AP6lvKj7wepwUom9aloGgprys3Kjycn6hN2aDXZ7mx
w0sem802hieshfWvxOx4z2D7sWb5CBZRAkdTQJPcihG/S34FJ9r9qQ9MOopOAwGl
ZLtVDWVNUSncQnPXsTslbD1F8YYyZ0CytTEltkyU9KA0h8qd6mpHrV9wJIcI/YvX
HLtXEUzIrTTkegkT0HKXuujyo1cE8wZIlS9k5NDwQLOovQXAVts/bhVab91LsKzD
uIzFnB9S+/nn9fe/rXOuHnBXgeuTuLswz8h6NGmoai2TpYZz7k2IQ1pqPY75EbU1
L2WfTZCO/Bkc5Dc0Otd0Yd+9TbY55pxPWYn6k3jRDy+6O5ed/fbruIfFktf97O3b
bwad5OKuOm1QOJYNOUBpD44l6Q163+y2q+kw6QqSgTixs/0ARzZeu63SdoEE0D4J
ABb8kJ/fgrT2juh31Tj9HD0G6Fyb6qLW6Ntj370NHuCZEvA+AucN1mxyow0Ff9Py
pRX12751nAveY+A1k5bnG5JPwqm57Ignbcq1+y1aVqx/qkuSDNlH8uK5SMhjZmjm
4LDwpeViDDozay5zltTxbMi70TpVhfOrEdKpnjYLcdwNMb9VSEnWPW/dq5iu4Bho
MJR/jM99jA2Owx3mF8vD5bPr+JtFdB92GJP3oVKs+7LcZAxOjNdLmw25E2uM6wIX
+YH4NmLqHncPBbky3P/U4zt0jiJp9J+RHoJZYxGoj26lKIia8lNiG+KQ6Iq5AfVT
iGHBo7Z0xDUtVzORllA61pp5BvKePoIyCPwL81jSd2Z7k0gWDqrvgt5J70pW86qG
nBVyjWZ/MqnJE4HD0sjKeDtb4qK/LLKuMatsjyAMY4ysGedo+UQChiV1zYXGf4qk
Zey2Ru98AXgr9FAgPKN0mUYPnTnJ8QYdsxNBgCLRp0U+3ILNh3qrUrFc6hGxBFBt
AGMM++PpRpBgr/iXipi8CmvChCZHz3yA6sQIU5NkKiutR2SivxYCzFO8s9wqbJlt
lsTGBt7cbY4ge2Iaw22fxoH1EzYpb0q6sKQ+d7x9OXYKmm5mh+VtD89KBMb27CGM
KRfMKHPWPBLj1sBKaTN209lTvX77uJqgNF84GwYNmCyI5OEdbcplfL/hoSectwUY
feyqtVlpcoVJcqNEwBmK+Loyb3lZk5Bo6SbLQ7aB5cxo69FXxom8ykZWwADEc/os
ZoOuX5b5PgGGCyvd/s8FjwudGEz9YcYnIOtLF5Aemw/xLyFmiriJ3+aouMEApjRp
LNYKOiiscGQhJjkl98M9wY2dlD+UckcGUNgfuGDBmM4s1kTXeUPQYy3jYSSsj8AU
kJIhUpHHO6NOuRUpwYnbaDkA/7U+67bZu1E/iYpXGjQ71BQJeV0pcL1x/QeoZO6+
1eyk+UT8RFosKITrLIYIJ2YQSqx4uKhv1s5iVfyzWuIpQVCdqACQzt+oVcSWFs4s
g9pasGusULmApjNrx7r2wbtgG4USpF4R9kIkQLPMgyGQLGhCi+/JTenQBYQiMtp1
m24etiQSnETB5E5uDwdZ+qGGstkp5gy/iNhhYz3Ppv/2WrqqToNm6Qgvcln7mS37
gsPkbyIF7p0On6Nn2OVdnDpluHCWRDEus2T8iDLBP1t9lKMCOodaHMSOuAEnKqJZ
88ZonL+CS+RIj6znPfRo73hbwZxHvT1LQ7fxRzAKEFc/usxghNykD/PjxBl17pWE
suUk0buwa3uDPSIIGqUKBSlD4XhXmdk5BupdajCSnMx1WGFFuM4EU1Xhc8AVyNiX
mDJIefMPDAWqVmezPbK4ZkSGeH2OyyCWksDSvBR74r/x8T9Pgf7pKtGwMTTmxXZn
89SjSJABWTb6sugMoLEVQQnAmcqeY07AgCcmE2wqHY7N63R+JbAs/ziKiRUi9ERm
iC8o/tcl519zv1nqVwcbPFndUmO1pK+d+7dFLGjRxvkZmORhPDTf3ljnQD/7fKKy
gsoBnT67XzAfEhbV1bgwD/cSH/gO4WvDFXE3VjpCBnEKN5qbkGYJDEH6oSqd+dUt
dsHNifym7vEvgSRcMbFb2JXpry54gvew/UZJNouCTb3Q7VcEl+8rpfkvg1KqnBqA
vqEFItV+Mh2yh5YBRngFKB9Pmd8Lj9IzvCdw0Rl6WBgHHkF0CxrHgg31XfDQT9Y3
iBViDStrsVym2Zale2m2enBsOgo3h02zvrPQ9zGNwyQQ8TNco04V9kubc3wPVEIt
jZMoMGUZR222f3NTLlfGbEb6NFkgbelLtUQo+HYiRZG8CoS0Cgi7Azq/9dpphFFU
uGkv3ezgrQZVlJV5Q79d509EMnxohixYmkGB1W8SECIF2yOC1vyPkXgCWLfTf8CM
qx1cUO3dFDVYNmaCe6FN7QB0h4IKFFRe7j/4a7NvvgnKrUEaNX5Odga+AlJ2+H2d
cbMJyRpnqZUziR8p99YjsKPV4xb9bd0N7hhFrt3AEONnmrjL4zve9PvtNUjOPcCq
KgMHeGNv2Bw5wffzNZcAUBlX3v2Rp0LqFjkDOZeWISFqn4RFQ3BP4ErQlELi5i8q
WYvj3CaMRDs1ao/zYrdfmxKcCVv9o3oXHO0XXyV2JvRTCCUoDQlWPPwM4uizJBOy
obmYhopajgvAKPeacTUN2Q/O/vYeJ9KSymJ4Q2udtPBCPJ5Z1unUY8L7cPFOk5KP
QQQQTeh9DChZ5bLv7+eMWtozxfqTahiVgZ3pgihrg3iL9al0s7MSsB8Jd976+WyA
etqzCT3u+bHa3dDtCQf2I1+HHVVKR/Ak9aQORjxPzr1rtQ3Dgkgy+6Qic633MQKm
YPMwVf6jccddjeuegg1LpoOITQyTVIErt8YfDbsdS17XourmUsjIujQqErJXyvZl
eNsC9OmUHmDUdmK5IPHkSf2NjiHx4ZQ8kS90UoerQxzDnJ0Q5cOaaPgCMKhI+owr
e4Ebz5HSHVs8/eAmKQEeNE+qwqqj2sLbiY+WVHZnYxNZloiVC+Un2s9np+SY3DQy
cWqhUMADmO2DTGojZPvOVd8W5008juWyoDHhaqiqsWC3F8X/kWZO3Ek7SEQ7DOb2
NpokVkUSQgs/7PCnWwHRsfcT2bqzZZRgQI0KaMa+2pFs2CSCUc9wVW0A3of9cueP
/J3CtyznhsW8nO8+jAvBo7phCXe5MfMJ6GM3nCtU3018tBPtQDxmQToLi/hSmZq1
3M4GLC52+hLqlrTHJvwbN2JJnHa1X0gAXelSsrSVxnMefWKDoflXTIWJTrEpm9oa
9Qrl6HTXtuOKTpjGQUTta4TlFRPdcuBvRCsM3LSyrUMX0yy3TCloq60egOuovtc3
30vRNWnynTqkfuVCbxQRNiz9dID7iqMAr2bwXfT45HS7NFRep2QQvOL6lrrNbDeP
+fgkYdZvN5we6d+giGqUy6WptHp7AFIRZJ/O5/ujuWOXV+jtLvCHV+SIJYEnKOga
WHJw/Dr6GqnFRLONip1RccVjp9bulH49OE7zqZKhQPLNvhUK7b0GnxrLKYhcvzyd
xlUqHvahm4Ci++oRwAuDzUAeioPTt8iwB5zkkk3/xBD1fDjfr5laOs4U5p5+KNbk
cyNRjxkp/LEfoGLRl4WdnH26VlFl36he7d27GK9zva4e8fCnTDEOJw7/X8sV27Ba
B9/9VvW5z+IQan1VGBw6DhQoDYnbY+izNCQhIWrATFhBe9MuJSyWGur/HoKBlgpd
rQmSIMOHk326lpNZ2+aBWNmDUeQHMGt00sN20ui5OiaqdUqCk4Rnt8GLzy3GRP3v
Rd+LsHxB6iGrPXYDS4VnFYvpoZQ30Cy4v09BbisRnZd2Bil6pAni22C7t5w6b8rv
NtPsTTKk3yeiFX3WchgLyWw//Uq3Zr+1FFui6oNt8GtYv+Fv5f5C+dgH03wdlVvk
wPkU7x22+Tb8KCvM/zSPRpaVOh6LWk3kIJgBAuag7kZVqzj1rA2NZI0HN89McfOa
MQ42vn71/w5+aNGDI5iPzxrSmyQXVy0oXQDHAdtU5QWiuMojBPGJQoIH0MsmUXyA
elcUa4XK1jwMLDR0pGnZb1Zcc4dZW7vYCtbUVbaFnFfAsejbLKA+3yR/RXJIJhYv
kNkQDEbM7lUerQ0RDAsd76woHaphjfjyC1t9Yxjtqqohs1hmPdZI0cTZPJoIlURx
0HDD8lakOcwqLpAoiI4pDkwSaXf4lYOuRM9ku26BbBzr5JoIEnoy/1SjjHxb8WGT
XEh8zAqdaUQumbNTtBFacFJClHmT/29AggdZ67r32z+a8cTz+w+10HNWxkiV73OV
14n1bOMVXf5G3NkfveHiiXE58tWh4y5r6rn25cIK6zcJDSbSzbUNsrZXXWcOny7P
UirD2bjQcGcbynUGqaLzzftIv+5G34hmnCgrM/YhbiEQayrZBTa7uwz0AySPoeV2
SpdrL1Kdk5a6IVKtjuIaBHfzLHKQnPniBy/zdUQm7HTT/T07nwcn4xIYtNLvL5Cj
CkuzAs6nIPjp5nC2sNM2BK7AQbNNXv3bYRCHnRUoFBZw0rPImV3qEwBYZ2kzxvnd
EV5XNW0zxQC+OoDI/wG/LqOBsypn8M3TFYuve+Ag3G2On3ItEkDGXb0WQ7ghu4oa
B6RiOpgmwTktelO+fAAx8FYrcxTMBYX2cmk8bV+tat7tNl3D/vlZLRuSxKP4MMOT
Q2aAMk4y+Uqle8ovSaRPTrGvbEq/qCR8QSDzXDPXitoNuHX01Qgy6EowJ0pXYtwA
W0w+5KfQu44YBcSEN6bPoHAPi5QzUth/JgldGKGPGJdfLVJNR42fxHEeWhBPraOr
IYwFkkkVaJjqpyJphJPF7W/FqKt7QUgPAmCUdrBzhebU9K2V3ljpXt9/GZBYb1I1
GjYD/w/xvuYYqEGm0QNg1KBD6TlankAui4rj1Nge69y/4btuzqjxra64HfVFZKPw
htlJchJxOHqZrmHNTVyKGBI472qNc3dWoAA2DYJAdovxKIf3rudl30LsgEsLrIuQ
5JR8CWxrvDOLlfdr7mU7yZdYU8FXHL4VVR9/VRnApc+e7y8pzYgfOV1HmTpWN43t
NTfKwGMTVfuXMtFwAnVk+INMyHFIp7lNsUzJgKpBcXCIjd27AK8b9Q6fA/N6tfV/
s6PUz84UFxmYUts/pV7UCidNWecDUXQWS9ZEiW3Ux1b4q98RW/fGzUV1SO+ocWkk
k3LSEQJBFDhR/cmC3sihyhnIE2G8a8go7Ni5pUmDF1Ormb3CPorryl00HIdl6Tg9
cEBEmT1VoHHAFidwuTm+0UrGyFOkAAIEcrB8U93w65fVU83BL6ZlekNUQAPrnVVC
V/I+na+aYpru8f9rLqD+cat1wYSzqYWU0ZDqqVhthVWP0Zhe/qDlqzVUXAkORD1l
1+dbtqD1733xtZm98oT+pNkKEBO7tOh3m2VJczD2fHj7ZWjlnH8eEUd73KNFnOGH
TfZ1xsp0K8cs8od1B9On/695Vo4fqEtHTt1QGzSHOjQCwLEo22U/HHbNkoS1HxlH
VosyoDVde/2VtyiOX6lfZXO4BFSDbpyMJ1Cn1zyyWn5p/NAGt2sQRDYXyeR0dqBP
ngzJgbfFcLpcv14+BndglHOEOsuNITO2NXav3j9XrBdj3Pwu4kOScVWaUajatZ0x
oOZvgMCDgkvZjebidljUgCuMG5nPz5oeA18g71dEbqxrBnfjFtZVgHZIt5uNbwfA
isFtAjrYcb21ofSida2YJSnUzGtaaTdpk/9s0/WiMdllk8ijhXW0lHzg6v2GTb9x
IuU52l5ggPe25HNlbywrYUZKzrOZeZoRRtk2kdtCDnka97hjo4JoETbc1GaBWtHr
eYIJvSWXmgHECnaSCbwZE/FTGIZWkgnQrMGAcCEAEbziX0WB0EN4v63y30N+z60e
OQEjAKlpejpcP3Nebw2z54eoUujA3uCLSEBF2lgUGVMu8/6A9/QNODtELQIYx49p
h0x2LXErdh3A93f8xUOCJ89F16iiKCXlK4ygPU42soP/Y7jtShH4hRxd5dFIxNrC
s2dzVMw7kOwMquHYH4ORaqyR4XEIm+P4LE6yGg1YX+87KZeaG103hPydJNH14RPR
zHDrQW2LeSxCsGO+gXbNzNUmoqRq1lOgRTokoq2OTmsJS3fJeIwXxlQ2cYTOL23A
Qj1u/vmY8pEplZfb0pNUGxmuTlIWY8czl84rrObqBhZldc4Yuar/2HoxaJMOoEQT
VCblPL1pA74LFqfOPm+NyA6wSpv09mHMJfKG2UIWT6GKiEARL1c5wf7KCmvPmeKQ
W84kcMCOmFlsBnGN9XRHgiZ7neRL8YMwcfuDZ7SVTrNIKifXAN5QGvJ0cyqoVtgs
nMsOGHF548ILLHmcyi3W4hgxXyFnUTVdwQnFl3casyxLZftraZMfJYk8LtOShNDn
xtr0wGsMbRwvTjnNw/v3kYZFFheNwmYARwHuzoNQHyVmoHK/BwtKYSmce7IsGqFa
NIl14gAjDWYz5wsNQbOZaBb8MTjN2xWhW4UtbUD5D2enCnl4kbVOAmajTLSaRV4m
yXOze9jCY+1vW9l/ZmO4UDyQuWCVXzJ3Xwu1i+xOtuaSHIMkS5ipOy+lXjRRlzlT
88wTsYvIwJ4og5JOorE5Fv3b5R3AJpkQvyETQ1sbfxfO2nUtkd0fGNw3uXW28Cjc
iIWHiufZk1fbKbAS2c6k4pQC3EM8OWIG50FiTjtNvndpsyUPAUUcCfuZAFM2qz2u
yzreJ2A+haFnWiA6O/pyQCahdgte7lc3Ul/SwFMnkqT+njlAsTiYRvyj2EDA4qJR
Qfg0LscTblchFngplZX/A2nW2zst38Dw0kHzyrnqZHKKSW7+iFwrHq8hZR01D98R
K1go4Oq+WJ8QrIugaWOaQj1ANIt+pBue402qUREbkxaDQZ/3yiEZvoPDqRQh6kuR
07aUBzWSXw74Um8Kp13Qa63Gw5RCWXIIM+suo/mc/akm/KgSQaR2QfiIOBjP5WVX
7MvTQ/AmtTX3hR36tB1Nmvasm+wCU9CDLsicPR11jXe9t1w9Y9XWzb0hh/a8Bxxh
r+U2l2ckxBoL5W58yKJ8lV4PVBy7hV3hKBKUR12ZT1JwkPPtmxvvwJHLLQjdVEQd
DERC25UUn1eSQRHOyEJNzkVGRjXMbY66l9pMs99D8MvBbSL/oGn+4Eit/w/BhGMg
x1hcwpnQPF3WBizgynXV8eSla4UbvN7iaTS2lnuKUpM2ffm2fp6g6AF4yADgRlcZ
wryOZdx/oG43JL3J6omtHxQDZ1xnvlvx04eTcdd3758zeGR51cxlj1mpPBzOTkHn
PJ+tyGrjcJau0seWDheSlx64z8BOgpy9mgBDYJVHEVJq+COnCV6wUho1jEq6PJnu
XqSYuOpOf4MByKiDyidNNzUJPY/UuJ7ShOlXdT7P6BxRhZ61LtcId9BjL4h0sMem
o4zvupNLwdc24eutu91sa2FDxzBIpUc6XAIbj793/MrSnF9/KaVD3MwMD8gmhgz9
WTO8aOLBW4oTA/13TBhKbSgttkkooxcCrle9J1tIBupdPFXSpaATm8oj5jMV1NFz
w+VUxUH9hCla1YHVedCpBsBWRmNgcNvA8Y3umebCOaGTWGng/vStUAWN8MbrmZJ6
Mxj8KgvVgkZ2Jz7DqJHoy+RPX0YYIgCzG6fgpR8FJN9No6rzl0JNhp6scVXV+oFN
njXwEKuoEMt1EEFooHj6NJxUho++4Olxbw+AuWfGqTyXJ0Y289p9R3CCXhadj7Ig
+pXl/fPVBbymibRFu4Tw9JiSTlDbpFL6XzWA6f1uCIaKqEB5+35Wf8t5ADcRohRq
nai7yM61F9XQ8XTnqiMGex60xC/OP64vR5z7ugQSf/4kK8OVb4w/53CvukFH8aGv
ppNbINfd0tFZzwNyuV+GnO+IwgQxrtzSqHfwI0GAG89HM22PGJFwUjfaNE0VA4K1
Zj9JPx1ef5VZ9NdXeWWT7L8hH1iaz/0NS72s5DMaBgWqn6v+eb/mF2SYBQKs86zD
FiHetWyeuriXJm+EhvYs7m+sDR6D6PCMDTqsOO4Y2vtu4yvcbxeUxacteaRVtuc0
Q9cyvObgBfWRaf19LV1RUdKQ+A8HfMiO8WvSy4b61n7Rle+VIgs8n/3scDmvB2FZ
jH3IiMsyJychAYDj9wiYoASwXgI+jbw6vhQLQMBvfciDiD3iMlfXrFM4uJCqdeSA
me+E959TOedKMit6pdzeFwaG4LDqxZm0GFt/nElHlWKuRaMN+6ip0htf6I+kG2rr
rIEuOmN+Tiz27wsXiD5HyoEERGBWs//Cvz7HYszWAnpNSDj76qvHdk9Ck4Jrz6OL
6U9Zq4W0ljhadYLsHZKAbV73vg9AV2ioUZXxFEm1LjdrN1XcOI8/2pvDXcBnoRXR
qG83eR0FYefmikydaDN5kXX0zh4UTqYF6Ka2VOmAjkAxDTf4pqGCC6P6NDdCRvXC
A3NQpUsr9sZSldQCCc/VCo2LkzvbRExPpVGccQYg+y5YBXUT/EmPiUC8JJKI1OMk
Ed5JiNx0XffSmR98XDkhrCsM+e/zxdSjGUZa82cOaK9slytqtqX5w68+vG//Bot0
ezwHPTnE8ebpYbgmwlpfZ7qtS5AhwmhPgXr/cESS8QAKCHOSiGn3ZKifk51c23bL
lq+9MU2b3tfDEG1ueIzkWIk4D44vOiV8Bvmd2BZcQkTSraIIU0kzJqKz8bHzJouO
Kn2/zQBmVUoHcmpshWQVruTvxLAg8qDoKg/RlcjJD4bjygASbiL+LjQ9cyAmrzFE
fB68nwM3mg66/5dl62L6WaS0/Bg5tKb142HWdU+bCmskw/83T+CdSic28XzV/wRz
Pp7MvsdmNwCbwf5hZLxePIPRAcjHFmnHTVAADySjAMTKiQAYhLmazQZn3vOdjLOl
XtE0SLPP1LsSePq09PpZQdVs4IhJisoqh77oRrTGACxAwJg5JH8F93oW3hUQXH2/
FGhvUoszOlRSq/tcLrrqoH1t0s6ZrAuALe9QKvo85EXdJWx+QJ681240GRqMsTOY
96vuwarvRpx16zWEzKDnf5PWL6+oP1jFFrbSgBxgRIuGbYH8Jqd5hLhi6c7MzPvV
klW0P1/Ru6ADWTHBxydElt2JlHkqnyeNhphEEDv1kRGHDkz2+8N0149rxPGCIll6
erDll3Gi07DOTVlB1G9lwzE+Fa3msU3Z8nIgzyncqQMl5r2Uk3XnZp1z7j/+yOjB
U+YmatG2lpAU0oRG4ucX+Ei77YTzPprLUX0OujBLi4vx6+OkyPE+47xD2I6U+TOS
b9gD5kMLpjfW5h3BGb71fLmS8Y6eY7AhtEswA4BvdduT+n0JlFsjCGjjdlLeg5zl
REy7vNvJst23vEQSufVnsg4mhgdU0gcyyHn6TT0BPb5QDD/Fs7p1kA7WStfFRn1J
+C+5RkEHoNsGLcSWN+j6dko16nyVMXBgBFTP+xMIeyICjvrJKFuYkaJGEMYUGmKx
eygSJeoMLMjHE1YBq7igWtZN7y61L72nB1neyD+qar9Qgy0XD0BmxAyy3l6UXTIj
ROuj6ge7qUh1a8TdFmPvInZFHczZhihSNcPwF+TkL23eJ73ofGP82ZsVI0/N8uWf
DzA2y3U/uFnmGEbWB45P9I/BMN2FbwY6JKR5PnoyP+uz7UJNl54T5JREwwA3RnW4
B1xFGtEOwvjCXpVgsGNe2vQY+aONUZX69BFGZEF0XMeRXx1K9ve5lroShxlsczCH
6E275EaTux23jXHAjZ9a0FPY3fR8CxJ5XIWot1aaEKw2B4JD1ZI4leeOSTanEW66
/vr9Jlpvp1gOyWHr7jR6LoHfZa+SL0AxqqftMoy5vt6Lc2LpJc70ixy3tjKu2K1U
0YxZBC6P6YYK0+w+o3IQqKgYWqKX8/uthWg9Ufa7MRBAO9Zr1xXfaE3kLijOb/YC
l4HEvwm4xupLszDPvJ0YD6rF53vHslPnh84vYZQ+JSZSeg5fid9ppLX7PJp7L2dK
kzRJCk6EM7kGR3c6DHCy4DpaHRGDOxggCuLvRI4/d07vNqSy2x00MwABJ1bmU/rV
mLSOJ644T69ADwkPn2Xp55B7pNOA+qIjuY/VNgGjYQnr9LnlS8I+ueDMAgBeMDvi
sGgRcgePONuv7ZVbzcJS1H0qdM03UvQDmAXPCWDLg8DOFZhj2ZXzg1rLznLszMCV
g318NFAyvC4PujnX7NPgOLXJJbQDO0Q+xcQ8gYcApooVg02qcjPim97Toaro6gna
0ahzP6LRm1REBUEFy2bC15LEDnK8wgBouxXPbxzW6hqdbk4WjfR8o9DVFznLPiS8
GCTZvZz4mod3OidhujAJ+iebORK4WTQbrChfSVSPjRgvKN7PqQA6reQu8ex8KmkA
MBpeJAw1whM7OEb+SvLGZx3tjkbVNKNfCnmtcu8iflxo8mvqkSEzhrT0zEzytkyB
46U2PsV3uJ/WV5m+fb00YQmohM8GmZerqjMjMN2K0aAYcNqXPI27SaopaHYr4llc
dETqD1Zujam3GCr+zcGKznpZqAZ8fRhR/lPYtKvK37DRvKgtcYwLh6FG17Ws13lF
svuiVulQ+JqHXrdmfGZYH+ztujzWAfKW5469RSpdBTDfRKgjTO7f3PqTdAzMYT2l
DQm4K5jjfTq26iIcpEQsJDyglStkcDkSOZgu/11y4to35AsERNIf3FDeUuUzivr/
fJauk0OU9ShPgL1iGnjft7MQFNJqGpsIL4PCwip3dwmW2Q8UVMtbHpusT9XNZU3K
I3Rv1cFtTIkpj7QOUl0SYN6TRLgcvkfNriOsP9/z1GESW52l50zHaUNpioe6GDAB
aKsMerLcN4Q7Wow4/Pn3tyvzmuqy96/QS+XM6cQmmuTs2zx51R8c+rnjwF2bYyZ2
MAQLytcJNPpDMpfuH9q/3YJGDY8WxJYC6KXG/HKt+w8xfQ4su9ECt9zxDvoLlOYi
LsNQRjoHBvuJPj9Dvy9xXjsu+c0UWva9KWN4IcLXdgSwZxkMv6w0JdcM+rJ5FTg9
b/XYYGwjUdPYnt/w0WcrZc6z7h8mJ1EzVFg1V/rzqJFRAVlznLbySBL6O1fUlfWy
vhFyS33OdpHyr7lK0PBG3HTfZ9nCiFkymtAP+93s9whKGFKzUGthDCla6IHi/7TK
dCX3675ubtI7BUolJAddW1iRQbrRHBdf/foyCz/gpP27ClxmrRevZ67aZ342IGph
paasG7iFE7c+r63aAmYvca2nAV3oCuU3GlZG+jCQTIbGKr08j1BzTOQzv1/xFJZb
O1aiBTUW+7+jgwK0d4LmkAic9Qgfgl7v1mgbDrAlGNuNWZF4T8zTuh7aunNtUJ+v
/lEkfwtPkPkv2sUqNp5n7dsVuyrLh2heVlGw/gZNnoif76IFoUoV//31PTcHi+1L
TpT2HYEfr+qfTLuob5rb9sR+3rz/JHBz9yohGQDEQhili51+/uNoIU+6xvku4y6O
iUfMNVuhAQNkzwRVfr48+VXyVT76pxIrPKItZVw9hn2A6Nst6Duf+1mG5jgf2x2N
2WuqqPjRNpFSyd7AoJ++9CRWp4NqZC7gjMZz9QtaDES8stqe4xar/HNG40eQMDPp
njQU+N44zLd5lShz7HREr+mTN+MH4DItyJ0RLa6V5TaqPkx8guv4gUIjUY4Hjyam
No8Z1Vev1R5iMe2i3EDmmOcCUpB3PLRzwBvu5WgLR33cERjYRJPZ3CbivDJDaRjc
rTsPbwGXiYw8ePivLtwCk4A1QWkdbbeTYsjPD5Q5muXuKWOaepEXLIq8jS/NfYAJ
5R6Koo7ZuKQaxRZ3DU+WpA98EvzllZZM33bZztTV8GZiXBEc+s5wq3QUBLbrltek
l0qysFPznCSu5/dG0YlJDmSz1b7iAUWtJfmss/WH1uChlGSw3mk4vDWxF0zBJsCN
m3Rd0r3dqLYa743Rk4AcCCgOAVjl7T5VbncZMB5nFjCSyZSFg7aJtDsEuqcSEvRO
qMVZ8LpGRnM04w23oDdvK1eJjbKkpWtpXGtqINM9fnzmbvdyecOsBhBFE2OTzrrk
8b2HqUAQre6UYcNeD4oO6HgJI7XO9XI5OZcIj9d1Q5PDWCSIkbU9AXlmvC4RbBWu
WPM86NiKPRclimc5rInX9gvcbPWR3kEBiLa7t97kjd1ejEnaxRq3dmnTGufs4Up8
k9IyGhsSgFSIA2inZFRjz8uy0DyaqZOmJEKvgvgyY6pH73UZsJppVcGYnAK2FDxS
oZ2X9UmXRz60qRCkooqhBOPIx5PQU5vJPO8Hqlj3zTyFjXLiXtOa81Z/rMnJtY4g
o/MWi6liNDq2xqqhLWJtJGyby+rFf/uPxCdEHd/4HxwNTl69xUhrPiHavVD4eRfB
7vU+bEzU0VeoPA0qFX61/G2yaAmiHC62wsvzHTj2iso6anGwub67AM9JMJAkqKGm
fcbBqy/4OLoqcVWobbnuBcwLf0tM6xk8zjFseScfLJROj1j7Ai247aV3SCCH47j3
4CtrvpcaXTaEd5xTWuvwY8aHoa/tvrMFtetNrJ78qnG1TwzXnXhLMAkSkJltBlvM
L2ky7IA7HHq8ZMvvL4wEDpPcdQ5ZGNQ5lF5ANwglp0ySGpKY7iN8Tk3pUX6PYKR+
24ha5UXUtbHI+t+j9OTH/gmQvTou6QRQpUBDtl2nWQAHQxno3aK8qY/8kYB+8Sef
mQJk93z1jq0MjP0SsloOx7zdfTCUapdaL/wZYazORxMaCdSSX4ifUSq44/zwWHAo
XevZDjg2IR09h7I7i64DWsRL30lQuNHTNWRYH0ZhFNXDT6zGMDYJZWvkss3Lc9g5
ML3/y3qbtsKB6sJbgk/mFnZ2fPn74iReQwBzkHFyZUdtw+u51u+pThPcbmNLzE4G
5QggErzK6rVpISyvpj1aj7YxcrrlR9+WaAV/yohfg6cf/WRCyw+f2L3Sumo/ZW/8
Dfs3k45pAfCC0CU9IGa/wXzVbuND1PfnPZcrs685D78PsSHAJGylirvrkj08yBJW
/pJxpwE3BRupTXBG0EpJ1mdLOXuDi9NNlin+hSLOJLd7VYZDgVg6AjYk6VMfX/uP
qYvAwx1g+kiix2rg6h32MQQiHQF+ZniPwbbMhEHsCEi8zXvDr/y/7r0pSwzqJAwo
F/H0ZwgH3dOSWiTR4DBfd0z163ha/xQ8Phc2K3N9FCTUMJfDsdFOzyVw2Fo2Bxq3
v1lncCAv4wNhY3QDllVUmEuqa1zGUfanNayd7y8DSMoXdxWX80IcPXYscWPjFeoT
MPe8iNc/IAvyRgxI1DIkwp2Yli1ODRUf58Whk+nm774sLq/DMpIBVyeLba8ajyES
sg72UiYF4PNFcOhPUYnKbwlUNA72bAsqEzKb0sAbFKVvU46lA2plMQVzazw8UNrG
0aCxc8wNIxXLfQsBnU2w16I9mCgXqkTFdj6ueeOArph8WtRmYwt9xxrUwhqxyS9I
unlmyft099rSis/q6aS3gtEw1tQ99cO63IsvGS7gESib/1j+HIe/jyLcJutV/ell
ghDGfrNgZBVEi6BeOV6U+0c9VgSIUT6gqPX7029LH8npEb5GKiCEEHF4KTxkkmaV
i8tv0QzTUEKgNGa3OJUHfD4pt6U4XGdEgtrnQ8ag0RAsTg7I7DNHMLIG7psTS6HK
WNZKodrQs3z7zA2UVgsgjWwfMkMWF0C/9kVcjJJy9HpLeSuyN6Fx0lwwLDInhV3V
T8k2+qzCl0DFc4m1DCKMEenPXPB+QKhmVt10QkCNRna1MWcsEhRB4kJTuSCJpYXn
+TI79kQGEuwtKiCNBoixkNpZL42SLsn/bdqhxJBJWOjOUZBLymDOEcdeyIe85ucx
fY+3W4IDnAdgCw9JYEvYtIwhszr5iRVuwsH7ni9Z+N+DfGAT2/9vMvICWqd4OWXr
OOwE6Ddn1JbyRaKUT4Ep5t+nBGro0o8AxiM8QRVtnzxJuqSoEDSzBPySCJlVdxk9
8y6LKhfjNlDhGsoLjmMhTJ+Px2Pzto+cDkv7FMq9v5XazYIj+hvjq0BK13g8klth
0uv2fc07Fl7MosfPEeKMhaLFIzuODExg4AFEZ13cCOvp/5WYVlE+lPLz7Uo48L4j
ZefSzQSiJIkdMEdZmm3KzadUbNyo25Ja2xIJSNFRQXB9Eci+e8BVDTusl3hs8mF5
my7bwHFUqL9ThfAj1mhUHWz9X1pPr2qTASgjOPjZuFVHBQ9zJTYNaTGB+DQggyRH
Ambiz65JAUhfwed8l8dZnqZJg+mIZG6DZQlC2nhp+gUy9bWdBOiVKhz+X5EFszVb
1jlpRn+yeTTDF8qcaGN84/Zof5NILxnnF46FjJQfmAYr9cV8qd9vBoUTKBmniJH0
6sjLsIbfVzpV4gq1v7HSp78T6zHIogF6u14d275j52xo7xhBtKWncBoXJ30bsMnm
RdRXhZurWumrAtg+0LjhN83yu/UEd/zH6Ot7fMukIVHL30cBN/aXb07DrrlFtZw+
BEy9rBqK3R6Zc+NfTJkhjm83/Ar8YYUF+vZvbDJZBntJN2/c81ysnDE0eb/vVC/7
gExxFLFJq5cOA82zpEwsIXAS9+pGaZkz9PiWdabq06/FoRMnr4KKz06j5xxL71Hv
xytOklmIWTVlmzpfITld/Z9uMi2HCtZU0Roxirapli3+DRALMgEtDbsK6TtPZmT/
Au31E6wC8nevxEF1VHPOYgsE7PSNEzXsShZgDiZhkfgUdlcXrY07RTSgM4Pf+0F1
CQT5Vbr82EkJOLSEbPBCWmJhWyEKIBm/9OJGwwWZzFLZij8FQC7P8Do5bZ3k5/7q
Fz+0DppEu2Yqj6PmYlnKXWiF09NYdym9hvstJw50CXg/rj5ITrkvkMRhAXP8JAN6
DyB+59JR1XAGyPxJqmZ0Ry/CfZNdkADLdjOyH1n/KURX6uunFMB4qgtLqI/Kj9aA
kIuCJKSRjk+MwNtUCoWCHKaA5q8BbkHRyft1D8NXBfDjyG4EGXAqjOFGWAgnCNN5
K0SeVuw2wXdrDC49wt8QbBAJrbNrqplFUixGFX1aVHGQ2JE+A3JQw7DOjyCq3jlm
m7eJkX899oeLEsHZAmgfegnwaRgjHbwErq1FBdglYbEfmW91vDIKd8CHW5bFDZme
wEFaa3p6qwN8DcIdXXo8Tp2ryRCV+vwrJsYhPSLzaH0ziRo2KwNvFZZ4msijk3oE
KhkE7NeP42e+PEyhJXMStUqbhIZmjvTf2fM7YHXxighOHq9K6K7BRkBBmMljAzyG
OO9dN3jtTfv968/uBz6DkNo2HAV5YpJkc2v8b2OIzBLZ0uupTcsGrikP/3roYXw2
WCLIgZhDBbLue3WtEek/UcKwKLvLSNeLw9PgKlpnu1s88MpKwKlyWkZN5SGTLz9y
SWUTYWgq0PAKwHK/9o2j6as+KrVuN2Z1lOHYwZcfot4gJD6lHKBKRlCuKNNn/3VZ
z9pJ6xz8pqELVtdp1KitCHhx7v+lK2Z7c4LQGHcilqftpMI3h7YqdaWdj+aiS0TG
XB++f4CIr6h/wM6crdNoS5kxbCttH5O7dwwcC+bmXVW/OJvneQ4QErZ3HVTAaFi2
vF9gIQE3gwgeLJhvL5B9rLqEN7CjalIfPRjmoy8WKD9tQ3EwuKYH7pLkuR/fMuEN
hz3F8k/i/8lDUEi6hbWK3Pp8aaOynnqRli5u8PVMebU80Xt/+A8qfDnw0GVt+TQk
M7hD7I/sz8vBvFNFs3AxqA80goyI54RD61lKDXDZReg0Aj8VHdbVIwz3EiQd6LDs
B7cy8A2M35+D+p3vJDcri+yFV+dupsXau+Kvz1aGoDQfrU7UL+jNcrE9SViIOO6j
MLdvYaLjja1sHZRQqMG9ML9cH4CBatoM2lTXyyeqsEmxBuHeamAMjpP3+9oxR/AJ
05ywGkJ5fan3bkW40SzPOHGf9Ig/J7nkL037zYWfz/uXHEnJZIIvDWkx3X1YDdJo
2YOgWm9lOnOH58vjw/3GOO76QHasZ2UMrBhRCMyAS9vGaUytnY0Lk/qldBr0zpXm
ipcbwYgziOEImK56G5bto9QvBEFWvZ/zIBKrOQ4OdMm3o9l6ZeAPXnfMpgq+YIPm
PQMJZQn4KRKwz6dFjo/DZUFgprATHOBQR+b04Kw61qUdh00Ydbu2Nx9DPC+T1Z0h
S6NTcomyMzjK7V5tGzure+hruicqquJ70eQJsGKp+YU2UPYEWPC0O0aKHtz70Dc/
KlDLcH93XQk/oinz/aygS3mIl5saZ66R07zoeAlqPRXxlLrGBeML0uh/DrcPbmht
pDVP2hjsyXxjaudNVsyInX9xC4yQPFx5bJm8Ccg8fySrJ3urNP4rFCcyWi4xfwBg
vrNq5VXnMj/OC6tQdln5CUig+emWKRzi2w8uoj5WFUFqWrEb5OiwRgD/2zafW+JW
6EsCw0eW5W1TbllY3SEDDyz2iUChV8Yy3YeuFtKdi4STyvnTEflL/AQHZJ+CdbOT
UnPGnzWwH7mgrhqTtYdeGwYdzAnrwaSTspMBLX+FJgVgd21BWBfw9PJVzqSBNcug
A/9mw2OpBPl/E+tQtMcYkXgFefILNmGu4gLYvvxTPrCNkDThAaF5HncdtYGvA5ck
SYLKYor+B3wjo00LXsEZLaO6HXq21i1HMg5PEdPwoSTzRJyAOa/6u57XhCgjib8b
wFRfOiNKSO/yKMHa7Drbf+VusvQdIh/Arvgft4eQwNAVkxl5ABRvKVn3jsjS5mb5
JtRuPkyR+4WYwjUEuuMSV58TOZgq2V0wYvlpvyq2MN/Xuy7C8MdoabmN/1ErY+2O
sTZhoF5omh1q4h8pe1RLQkMCeYT8vlQzp+Dfa/ftSQznfTGujzxbic4YGoB+7N5c
ZT4oRvTzE0uhqiosJkix/J4ZVLqSnQuM+qVKLiEFvhONQUPoONwL8tj+no0zfBW9
l7bUJRNmfsiMbrqG7VppbXopCy610J1vSABj4PdKsJEqt/mOIzllJHr/C/13VpKH
lrufqzXDE+MkJ5QIUwLDfmUxviJl5Bo7q0CKcD8YmkNGF/ncdK1RQDZWy5qpaTi1
Hj7dLHAUGe6A0sxv9gZKn6dgcQ7R6CbH+mP1WEgJGcbB7nCUux0dvxlHqtPrT7+V
BnvnJvyJG5VHpPqSsm7BxO11HMI/iYCHWv/2uVR9gbyTpdEX7Ms9YCJwCqMifXdW
ClDFV/23KAO5y4lmvx56sEtL7zWz4aELANzvXuhcBZ3c+LASEZqWz1Fn4rbB4mh2
Y5FwrNayHBRVjDI5f+GM7NcErGdYdxLenGW+VqIDjNuF3eerD0dVe8dgtBsb7YlQ
hiPg8mImlVArv/aAhFJP/Qi7DzCnWe0rgPb7x0fBKDSeo8PjuIsf3JbJ77R5Dzzz
AQr3/9+yaDXISn/CiWjSxtAS0Y05GAR18ojhs/hZMm6k/7dr3OrcsVBUVD6jn2GA
aX+1hPy12WOqA0JXmCyIXoFTukcVLUma+aDxq7zsuxHEmUEIQbRZj6pRjkOw4YqK
Oct0aJ/o9bkv3ski2r1xBA11pbD+B6BvY6mZtkaROsLJVr6QPUKBUQG46fpJ3Qxg
vM0tHPC5zJwQtUFQODVocAuiGb7l8Hr4sTfB4SIplPMXXZMsAJIZ5VtssyHKYd65
D4Dt9thK6DfzFd5zsQ9MjT2J2vTvMa69ngwiafw1RS2pUmO+WHp0bLt5yPO+OjQX
UkH06xNVz17XO8EP6RzM0IHy3N9tjR4QkDEolo1mvVVh3cdZRVSwmyh85Cmw0obR
CZT3cMBMlSYZmhSxJzIZ2FMlertZU5e2alGScWz2faTKobS906LlxeWOf6D8Fevs
718Qmwvq6Ht4tDTM9+iZaPhm/PoisydOhNvFWOdeGiP2BWwSc07l02NcI/Y2Awc8
FjrVbyf/DeP04uPhHnAmgubVsEvOjzpEQt2lKD9gHArxEkoqVTZ4X9pnrI6TCSVa
pBNCbAC9AhogEBmbaJRvsQJLLPoQN/GMyO+lOPULRPFX+oAwWWS86UnqmicS4MGR
+Un/fuZOJNbAcuSeWa/3JesufWxWgGx8ewjNcr5sFm5IMrHxNLLumGhOqO26MxXI
3pRM4/qw7VA2Fs2eO1evP3Wg/bnDIImftez4x/RnNDGYR2VYoMJPctndYhuwhlmb
JyYhgnkrnR82MPDerUcgtW6mpzdgKJgMe6zLQpf8t93Oq89D+pHYjs8CTrApe6g1
NdqVwXLsqibQ9UVsQGLgNzydEFQ9daYQ1xN/B0S9oIVh1rVrHsv7YqbIsCbAMq1H
nrUyzn8aK+je63FJPBRREc+hAafJS8zrMPWCOy//ts/zYe9x26VYzHxz2XsUtwpr
7NxEY+bv82GU5y0ilxo0kROtn90Th4boVK+IMWhUrGI8RWAP0DyaWrsIlDZl5MHv
iznD+u4Dmn9lzYMmFqEFSFUxEAgWvLBCThoCypyNsjXL+IhCmc/5RMNeNQb5k0KN
WkfK28YRObGFuf/NBfpT/Hycp1SsbH8G2deq7V1dO62YWxjaZB93V/Yd6X4b69x+
YksWngpL6wnzAIFYB/pHPpMqpC9EdaaIbFxub9Y6FQrpOEXmi7eOQ09uFBJeuana
HaixDmVclmFnC+aM/5hntC0o9lFaPWbDfHnSrQToS55zsgTVD+VwtDwaQ8Ni27LF
zJCjKXLjTryPKSq15R8iT0BUw9OhaOn9LZDXdBctsInH3FreGcoOFBvFdJkSIZGh
d4meaWXf1I+769U43zUW/b0EdjcdchF/CtxQtIhrRviubz1mkPaNzGveMdwIDLiK
YWqaoh++ND5BJG39Fn9lL2n2jHU1Pp657GC1Kn6Ft8gP6YUD3eaQb9D92oZ21fdN
XLWuefw81d4E8kEn1lx3Pn2VsbnnCjXcUqaKxYtfoZSMDLiaVsr/UIWuLCLyOjR2
s/5tEuzRf5QukHqPGRI/zbZjyheR4V4Du2EsYNcHvteplKBkm5BGMpPc55jf2Di9
JFLs31JpnmT3uWeQyaPbjxyhlXfYS89XiCh6uPin1ByvxsGSGHGfgA1ep+Hdikul
WbovSq7y3X18j9Y3BnRi4uqB064TAyNjYHhXFo8DaRGuC1RsKYWdeF/jb5N5aNzc
y5a1XmWjB9QzHAV0Il9FL40l3qzzUs0DhSiZRPSfleAs5mexj5r0fOAlI0J+FQUe
wN9h/IA9hDEeaiJc2/hlmC5WxnNlQJs50bPM5v247U2KlwODaX3fss72XorHv7AY
oee0tpYNfrGLKuZUAkb4Agh/5KiGktKQKOr13EPsSzhbOHgnPwrX+jNCvZqGagh2
ibn/oLR9RIL7988c+8ZFNaJ+tXrRDsiCDAr5euDg8ntw3PRGrugbsYdzAwa2m5av
VWYXllvJ5g0Ig752vFY1T9YhEb+xW3HB04rSPSR71IyOfNddLe3zosNObvh0WCR0
kN9OjJR8CDxyDTR9/e8L0UjhdEX20KLsgXyxZGj++bVYDlMgzFyKUYjB+g7h27FH
mreSFzIJEKq1VQU4HsqELRj5ZLvwCSq1QOMaMEZ/MrHb0QJh+cWxty+Qt2L88gyt
d8rgH4JsfR2YwmQ7MuuJ2mFssUxXmcsQKEkBLDyApNdND070TMGxuBBq1JFmTPKx
1iy/XWFZnycImn9bFwBp2vpl9qAE0Ns4WFMH/g9H4sUGKf+nvVI/WjYAJ05obqo9
d7703eeLOaW+3M1bQGE/C+110EETKVYctj/XOGV9hRUs85kT+tJjVC8nHhE4nmYl
SzhFiNy3sZ1VXIIeWqJQu3Z38XFt5gaerSruDedETWVG/Y1b+NlQr5baMQhqSl5/
9oiUZNXswysgPxqJveYnEp+PDoisd3D91UFbwXTV3E6v0TbfWeqUG4H66l3dH3bJ
bpmDhm/E3PplzTG6pdSbk09LZgg/Hycim1bu80CtALigMFTweLsfu1MjZndNP6xx
IsBI1KuGBhnRu+6GrGsRy5Q1yuJD1loCKTdh80ySiBRyEthMETVIqlkrcHhY3FvU
idJFomVQhtGyZx6sH9BpZayH6zHZ/4UtOKQ+EdePVZeM0jvBXTLesDBAeeLQy3gv
PNUpTeFTdtm4dC5uziLXyO/N9Anc/I6r2dYo5PZFAPITw2NtqdKdAM736WXO+f4+
QYSbsXes7rCnGQkOIkkyMzF4P0S+ybytY6A/RY3zUXeVCDR4B6KO8usH3uihs6wl
PAT6PuBR2dlU8U+RhI/OW2xbMYUMmgvxruA2tJ3eScqFuAioS9Jg58fZ9cu+0Pke
jTPlCqFTncEQSsJPiBawdsY9AFr68J41SwjDOeqLmXE466kZTCPCxVRl5k+HapIw
3qzvEBTC7eZ2iUj9PmPVh+JXHWuuh9wERKh8pIoNKCdRjNpEh42kjjzbFWovUiMH
cuOV9qX6eh4V5jlI4d20VaFVq11dE3AkUbjcwLW3BPlpDXT+D64TtCdKVg8V23jo
Ss1c/moM+MeTSHi0tY1yknUYEBN/MW6kaM20CRv1kzxac1xKuBA+jSfQW9ysghv9
W7DvOT1dze7S3Ys7imRC4ogrz1+tW5F9l8dD+t6gOfIIRUgrkNMgCNPaJo0dmPWF
3jNkBfhMeP4zNyK+NQM5hsNghQ9fIqGU+olg514KMzAYQeIHgOJj9WGFVEwzXTNN
QN5/ul2OrQQ3zMCQSjdjjtbuIJfzC1gfYE085KsnZ1UdeEI+1qV5WtDQ08Emm/5L
CQQY6ciqRmh82qwmFxJGBDyUMzttzTMOmHP/vgPYueN3MYqZ6cVnzvl5Y+M3irtA
ANA0mmP1Sy8spsz6bXIZ6hmzPB1v0cNozc1TUyoPWLpGc8AOHctlLhkBT+y+kf7m
OvlugPItb/W/TLSXJ+8HLGDnut0rUr6V92fQmnmj/KAlcpwFok4dWE339csMQpxF
9Y54NfyARtv9OeYB0pB4ZJKGd+z5WRwUUtQQB+6PVyGez/PSzvp3J2K8CGh/DS8g
wzXjpMsQuc0aqRcE8MTkambqsTWx23oh+LzdDw15Qb4L8E9aiw6U1WZmVI8DJJ9m
r+3eI0gY5KBibaFr26K+Ip2Pq2sGHv68LXgIaKnmXb0lEoTcJhi5kpdvylz+d6l7
mW77bYJLWozqENsg+6Lf/G2awD9nF3ZZ3NkLiCOjxnMrIuUdIIUImm4tbHPldMeP
AWU+xih54Ai2ODd8XCyQa46hV+LWRdyKW7oQjHOw3VHeDxl3PpyjodXJtSLwSEUM
sCUVTOJgadb8ZWRpQ7XumtO5fbfaTmGlC/yfS7JUc2LxJ45YEXf6zEsu/3++kPyD
iLZDLlPAxSmLYEAifQ0gESx2y5yrSICKwzm2Ax8FZ1xbSw8wgSc8aTdL1zriPTio
XHmWJ7bZFIn5EmUyyzSBzRYuJkEJaJJ1sYfvBkcIOmPcG4uIhyzIN47mNwEk9yui
jiM1y1Z1fSsT/FBRy3rvinogynMNmvOMdF6dyzbLpXNUu1IKGTt3vzCqbjTOHW5A
dsmF+1AZSzr+tFypJkF+mj1crz/pxibq4FZwEztxgeyLIFa70d50Sdg1EtmT/qvf
qshE9fd90QDR+mitgkx62cjlFPeuDjUErYJ9uxE4rmooCO3FIJbPv04GuD6UCxbV
SDq9+Wc7DNHlkvoWJvkQ8n98x1K9I1aDNGX1dB43mcMnE8tzQBVZI+aTvPXNeRcG
Ie+f0RZnlC8vsYcfGNAjFlZm8vQl+6F4P0Lvwy8lVem11meT2w1LsfnHWxJTso9z
7G+V0e5GUDbxyNSD/22Pno2hEkVAPHHeFHJvqrLrwdjfSqTKO5ybxTf38aTMqdFf
/kZwIUgKxrrudhON8a0QKT4FK5LRFj8ZdIERDXVrzzf7/53dCGqWZnZtZIhCY7Er
s2WZtgo90DWcqsEtrfY1/lYkqjwLJqg9kxiJfGHFdEbt6L9stN/XMK+2hZ3Ub73D
de6PjTZt7NlUAsXQfOwM28aP9iVxwEU7vWC7MM4XVxp7ae2Y1oh47O9G9iBKAnkA
kOVpHWnGD+3j2K33QHBdVvw5GyAsp7gm0BWkp2A/IcDJlBRFy6q10z76Wf147c+F
C/T+7fjW5B70Cw6AjUHk20Ub54wBDvNn5L2iChlzCDViRUmLxPRN9ei0Prekw+7y
qp2l6y3kzFcdBOjinVxQ/hKpyY5W9R18FYuUfw1/nddz9FlA/uvW7RDbRFBYB/4H
B7MBjQxkoDjjePOjJAxGLx3mzJpGXnQKLcObwCfDFHvUF5/FARxoeZ+l6U8JFoCN
BkNXGlkz0QtcaHSdO29BNMUcTHYwHUF3arSuqE5Qb4RC/nyOG3Li6gEAPzPJokKx
jyRA7LaKpBfMMVIPVTn05idK+X4jkmazfFaPTeY71/wShAaPtV9nj8SRsjDayF1f
5DnsWNKngMxpDyOu60SvQ6qAWuj+anbwdfskGjEPvVXFfTguWM8LJIgAxnpqVFti
WDGREo38aDmO4RcnN+8nrS15/QSfQXQeU2loV3QkyUsZirID9I+jD6W7rIewEem0
TwVR0H0kuENflngpJs675SrF6QE7EQ4WHuBtHADjPvQInONVdcDs2pwj8xQNFtaR
BUb1IMKEOZyQzsEzu0fuoQPST7TFWBIWQHGSU3IibOJ2DXeI2xhDHt6jVPNpST/g
bmcrNaYrkF9JMJhUbdtQ4ztDj0nJWARNsUlC2Gd8nwrJR/fTae8bNVJcj4PsovEp
Y0PvPm9n/UOYkuhLSRUWJhPjlc6RW7JghxhaIhFaqz2DnlD/1Dkcdv7vhdcrtRiF
f7t49Dp8rxAotn93yl95jnsGp+ww75nBDaMMfPGioYMJcct+47fq1rLw4suEOD4s
haD/z/ZtkkgsCld1ab21RaUTaPFwl4grBNPU6GXIXSbtpJyKekWdtEMDHtinCJJz
CBbMTStQBgesX2vqgfv668Nd2GJkbEwmmbQKbTPPg4dhqpclNevGVM2xvNcrJs1J
dulMu21voo6s0o3WALdNJJLHPYoQX+W9XDwlwN7Ndbz/j0KeexAMPCRINF64wUol
62nb+5M4aXjaDXBZMt3h9hNYHCehvGVGuzpqnUeHl1mPDWQZSAz8OxOSwJbtsDzI
gPRQCuwtJGmM7dIz+nHESDgXFNhfyrP/ntv6iziPXcEnkA3WY0+Kc2EPYVfxUUOL
5QczD2SM6L/kkTaWpHnFZqANp/1L9i+0qSWVwCuzs63m+Marm8Y/dLhJIoQy558T
kASDLoETUejIRQx/4MD2ztcFBXfLv+RsCyiXur0begLHsFcFQTZ3c3Qk1urk7PIW
7XwpC5IBUH+lb5SR5wZaTzH0GeT3dfnWoWbiwF8E6lLcYO4jDl1qdY59we0/1Hfj
vHTgYvnIT1UukxgZUrq2KPBZOM+rRrT6NYVyHPOQvBG7Rw26jbdYY9nDF6CN7+ig
+lxVTAFsrwHgA7War3A/R8hxhaDoVN3VHC+vZZlgLdu+1Wl66pFz58uZ+KRKcq2T
AIFRfx7a+66VxvaKp8KxQtR67NCrx7fXnbaHypC0QokdiCQur8RSpzkBo88yOquF
83zKpKUH2+NZCeKH/InP7fmVE0FBvLDS8471u2K7pXUuZ5Uz07p8v3AeGHIKr8Jp
KyS1bCVcQStzNg1EYocKWO8pa9BKvQdV6m0Lz6Ixrfg15PCrRISuMvtLkmcZSGyq
1Q3G7Oo6aMk9wt64oCYsNgaYBcQdfH4NPhK/5ILZzGxs9YuFuN0xeR41N57lMp8D
yiEF61O0YcxQ7eXtYsKe+mYuU/wA63uxNmsspfNvma8xHbH8DXxmmEIPP30iMImd
x4rOdhuhC2h7RMeA1RTOM/Gf0jh7lvTpF5Z7KLIvPqeYAL698qQ6wIn3C9P8pruo
zp7CYBCmqDilwtcpJI8rlpWUOKVLPf5cPQgc2H8IyrEXQBZgVAeChdjeYPGTW5lx
1wLwvMddb5VJCw3DZFxelguGaL5lZUcKj343GS55q06z3CcLsDFXUZIqy5Ou6jsy
tYi0Byn8+uYJAD7xWKMm8elrFHE725ZpwDDbgSY9TivlyPlgQ36vVuaLojwdKvTY
rKadEwwmgmJCEUql0GvhpI+V5Lpi+oNwVZHLzZ6k/93iK1yAgkLmgWLIH1axGXoU
SE3dcKt4ZuThmsXdfD+zItA5CdpKkuQo/4E1VSwrYAtF5PQRkd+wbMDTn9duxsyj
Fes0dYCWg86dx0cljq41ra14wNMJfk6oO1fCD7mKZlSrYQrUV/N+OBr2Q1bg233z
YE0djl7F1HRiLdsrMYjerpI/R/rTqN2EPl9K854curn+/bti98BSz5dPa0MhormK
1qn+AAn2Y5bnPRLMUabjYuNpDWID69lRf7vKtGCMlSPCCNaoYbk2hNlGYO+/6KUP
b0BsKj20xUpTEtO1BmXYztcCn2EIqvZAHtUdfsCrV+jd6yba2bFOL6sEkjtD/Ciq
2pnv7RmDxWpmyBXcFp+876JNoy2oHuO9PP+YSZjxzUBipdoJtRGJ15RXee4I7tYK
g+1GDw+Hdln2x7y+XXOsoOx/pRjZ3j/xOwz4JKFBI/tFGD1/LJ29wOcl2COdXg+8
frZJWe1d+8KC3BPVW8wSQb25EiXOoiin4fXsCqAQ0dmDlrJmXK4U9Q6va/TlUWLH
dP1d95AtknHGEiApeLrXbDpVeGNdELdBU80IS6+sO1i0WXwEru61tl4cn8TPxODA
GeALz9FupatVOplGAb4tWOEVKIItqz347D7owJlN7sYHRtI3DW4Daq91gMWnX7so
IpSncq/Z3TLYVk0q9zhnhRKFtdEtziTxMFKCcW6+r0mwv5PUXtfRFKy89SfwdoRv
ulKC4zzb8DWD2/+Kx9wma8R9ULUvmp63T6ZoRrXy44RcDxLAcPHmqq+Q0klqQbG0
2YEXVlPxzXn+xI4wlmWIj4n94Y07Bwheydlzgs2ms4BDG/Zc46M+PW8oNwbbyeAB
p+vUeSNekKxtsUhXQD8neC+0REH+Qzc6Y+An3XvZRqZmkumcxfqyELqUDvJp+5tw
GpS6tmlGcO+efMscloq15vH3Ir1y8GI3JDM9FOToJ11WZi6XEQe5044LgR1+6B4b
Mf5MemEkzU+FPSGKPaM+x7OrnGHyS/BsTZvRe1d9rzFDU50FXTe5fvvgszwXwp4g
vzfzVRIDvQM3CWr/QWoTtTb2v6+xh5KCKiHoL75+1HyHsH32UeU9ECJWnrZQ8npp
YLt3J7KzfvXbK9jvP01KSaF2E2zd+1MIAoGeEl01nquDcaUfH2Tie7KFeqJ3GbT+
LbidN88s4rbhqLKhor1kibzWk1tLHnOFVsfX7atS9RWC+LIyv2gPc/flc3cHGcBP
nlZsheCeRQIVNR5fywBku6EjDFRGslwGaFHCLZnU2NuZddzBl+62cEDfe/X35eY9
Xnat2NrAbo+B8FwQTRzJYl6ZrXZs/KtFSxPPr2D0jDgV55u2l6jS8y/V/Ipxp//c
DSLj97WZ2kl7/3/tquUfvGCasn9Z2h3PSZTvnsk8WudeisJpeN6cR9EkMQPo4pPZ
J3Z6oGO2Ujts32Bxzoe34IKlMfzlyx1o6fb/YZnJ6+cQO8On4lI2+O0EgaAEQ+dC
4K5t2cmshHAUqimsKObU52Z+f3nRsZQIN8OHQIcZ9A8SDPfVxo29VdbV3YHrBaoN
NNBu6D77V7I06AcQsgyOx9i1s3cgAOL8l17BmgSq2KzSLBymfTxSPhVMk1W76sgB
HyrU2oXIHbaWBjqcsgll3ceK26Hjj/A03xFNhe/bT1x7lHl5e3UsUuR63sLwBNGS
WC88N80mJjfkc30ik0EuSksAz5ut85w5amM3RiWOOk/hjVP7Q7I9OMbO+MLQqz2r
g89O2xVQayXWEphFw+ZK5hzF6nl04M5n2G/llmZd7bxruaHh4x9MtoBAio7u8BCK
7REKxY5RurI/bWL8aLxONk8UsoQCSFt2rHVuFvhUsYnqaXdfaBcNAiRdJvCLIFht
iAJ9Nf2EeLICfw7YAiI3OFLYRsQzU59OpE1caac2khReFpm95i6JeHNHPtcXl5BR
Lz40ojcsj3WVubCPTkTv88DVoa1CdEpNqYls6n1ugzUPWbqKfLiDPWl2bLwoDpeb
j5qBMTfn1xrWYDncL5Xwxbq3HRhp2EuglXMB7kgaPOCxXt7d5EtW6tlI4x7UTZTS
sc9qhSWpb0dJYtKctLg/PS7j4v1Rn21l9ipy1Z7KH3i1eGHPbwy3OMa/VRjYs1yy
WvppPiPomDICEN8h5I3TzCcgRlg90re6dT3r37TF+XGCOj1qov9e+azTA8i3r5gu
/LCUhrnPK8HAZ5+zIhsFXowRimXp0Z/oM349QGjs4DzYUQRPfhOvsWLygtk5wxY3
Yq3UpI4bO6HLP/QHTNHztfVU9734+3pNsAPtfxF6dA6FlDeu969Rq0h/VNFNrKKI
PGgRPBlYjd+iXVzIKktUCVdnuJIMjwWFaqgOm80kxls09H803591MXJl323cKjbn
rfJKVJ5Gz69peifSG8OVGleiwKhdY7TWcocartX/dzFHUQFVbKyqCU+2RPqoWCwo
k90/g2/1Ikc7I8z8ImOUSSQwt4yMnlGK31VAebZMOkoAftpQ9XGX1v2w680ExKKi
+cMccRN2r07WOgHmLbrfppz0HomhmcpNsD+ljDdwU+2jEZ1qj76foCn4jVSu9CDE
KOdK9LzZYcvKmcEOniZ9FaPxgvgD0Iztbmop3SX+IvLPRZia8wmvurrm2799lJ4d
o9kkLdceBuWvZBB0KE8mL8IMlhy3D3BM6XnGmzXFdOVKMkJDA6Jjvh7XQ/wViUYg
4vRxoi1MGqsN3J2Gm1acsPcNqdzdTCqvBH72ijAMv86IPl8aaCfs+L+qAcUxEEjy
y4R2lAZVATa+oINzh+KEIxCMSt+0xadfCYoTQcu/T2DvabMToielXGO/7dk6MCzV
v71XV9m92waKByUzJakwzdzLaM4U6jdwWuOlsX0sl9gGP+d95vjH9b23qVhAEASS
BgVmCYL4NE9Bdb9w1ATkZovnNSBlUgwbtF7ESRjcUPdnjH0Ms+CCCqHfzcHFWBtC
gdwtqGzacUaFR5aMpLVudlbO7Cmr3kX/bTOcotBPxm0TX3PEruOWfwEnItLm+9bZ
WCUV//l974VfOZ1NcgdH21lD6M3S2hF+3yq14XWTqktwPOv3rWxFgcGG1Fx/lwtP
fEWlGAO52+1Gitp/E87U2KZdpx+TGZxec5GDuVpHUZ9tVVfqaPU/sa3p9P37lxkS
vlqnSryP0LCPT0VG5UCGpL8Rnr0PqM36t/WaUX+wbHjjONpRsgiZcmI0Gpg+STjp
DTqVelWjf9tA2PLR95Di28SPy1djk9mGQ3K8+7KMSgyDB76/AybzcVSJ6g/QbcEJ
xF34LSOeCee4+ejrYWTzvalkNlg64US9ECFbT8C9LockQKOpnvvhjYPq/uVHI/II
t9yawD+jpJMePrxmUCGSxxCwpN2cpjt8LRMWWhrTGqgehD1vgwCjhwRCOrF1CXvM
m83Q7imLsNGBWHSCw+DvO2cIGIPPGuB7OpkQGL7xS9tP4Z9nkaif+yEu6aWd27uW
G6ziBhLB/4Sau8mvpWbYeZCp8KJXNHFehaGvXKyqNa6l1pdRgxZfjaEbNRD5JKWy
CvTYLaLe5njDGS/PJeZi0aP5c1IAwF5LdppEGyvCfIPJCDHtROdTF94j1EfohXLU
LHoAxXRMzbg9Y/8BkZLD/DMVpziNPeQlI2/hSAVVKYvnVYpdiFlSxvDvusIDEzbf
BEChGTRO0Qoi8yERowT8KmKn+joJu15eMpuS+A5COqzQ7vs9lCBpdpbdIhA3sxJO
vwuSwPIhr3/4wfAHuGj8ksve5+VFIOPdX5yxJRuNzF9d7P+tuLU/FvvWdYN4afDN
rER7WORIBsHl9cLt7s1StfSQ9FM2ea87QO2w3SYEIHu9dgC64cil4ee09GHF3vhR
Gxjt2KQJViRxxg/xd/HIk7ITGeYum3fuHjc3W84q5W0HznLvZtzAR2I8+L2JErms
JRj6pJ5JEaRvQSj1ZLwwLl+nbDUdIR229jpjNPzZIEox0DgYYRYrj5ZWl14YmX6O
RkcrJNDesKNguvo+VUSfbzcmc8UakxrAXDLcAkmD/aHf1HVhOv0modCpQY+2HX+U
eeP4YBOs7TS7+sph30ZFHy2YSLD4LLFa1tL9hSfofJO2G6WjMyRV/BxMl5IxtLa5
Ele/srP/BgWbIOMBtIf/11eLFkHLJkwsyCLGHs5g9+RYAvwukmrnb7eq/CYzsRjH
oRgqPj8vaY2G+0Vml+up825gBSwtMT/6IqzkLyrPSzYHvnE8q8NPZXzyFizjwlKm
U9GH6CFRdQB0Gh0mW3ztKVYOFPleeVQ5+WKoxNsuGJUGZmxYqcj+p7NqxO69Ztgf
BHSIjMu9EjP4dFJHQenRMLN+zXlpKKgZAEBJayzPfOVB6Z2uKVabP6TIi/1sOC/F
noHHklkecBjQMWzEbml2D6lQd4Xi2W70IwQuzss+8MMqAK7aCyLkPbctxTyw/8GV
M7vNXPOfUahe3byccapf1RcVO+YGSdRNYwUUg/qQdULwSU8/AnvIOslWXiTmzXNs
q10YnlDh77odt1shVdjZfbTT6zQgkalWxvP8VDqS8fmkjj2AO3cg8tSXZy6g5c+Y
qpfnDZzeRtQS3x/h0+ocgMz+xcE8EcH2aP8tRKrgIn2tRhdeSX6YRu/aiZu81asZ
erduxQDfc/4Hvws3Krcgrm+aeN3kL6iW5H8zA/bJ31SJR5m0pzlcYNmTrLCX0sDQ
b+SEKa9KRmSe12C3uBsfcWcI972RHfEOo9/WwdxJ9qe+iqeAtYZIOCFarFSaxuHl
Jw3qexlhgbGMb11TJfssczhpB/PbRnbx9upMh23wvHigt+/uIgmPjnbZj67wXudD
7msKioT8NwiQTA+j9l4rcWkkhLjRQmeiVTr20TmbbWf69nqLC8UhQXm1HVz1p29O
GoiZPd9zM2h7eDiL4sQs//5C8ZQQsECA/S2izzW8r4ev6dbhYbqdZMj4kOAzXqUi
m75YgSUYhbDfZxYZSAe33ImbU3OM7eRlPoRTqPNdOqAg+NDry23geQGzTLRbvMU0
BsghG0hPQnRdmQTZ+Px/m2zc9SeX4aFehrNJYfn0ZHaNaEweeXoMKafIZBux/Fwj
eiY8ZVG1r4t6UWDeYx2taqzv/IUf4ZBghggkkVv7ILnvpdNgP+v2doRckTxViWzK
h4QCwl42oTFSpy+6LFxOK74+L/2x4mAkCBP81zGd4SpRhMdz1qgY6/Wn9FgjQmO7
R+9pLElcHuBY6orIGj7xfCXPuZisIgq1w4Zc3cFiKUStutdrujYWTiLOJXPENA6d
jrbDrlK7Xnx0ktk78R7sX6vianZadpJMH+HSINnANgn1FhOF/NR7I5lV/zYjWDZD
mO8xO+JNxWzGlO1EJehY6jFGxwwMtfFCtyS7JIblgKa6ISgu4KJbo+yysWf30PTk
UEhGRNgM3CXhh0Y6jkSa9zcLK8bngqmRy4+agGm+AJ+de82st7xgVbBm5PLKpe14
xV9Uhu0N7FKgFjsvPDx7PZ81F1KAETTN0DWeXRu/IhtnSerhP5L7aZxQTLeptywo
3WoZOLDr7oowM0XetB55fNXU3UrbB8aQXC8MGOiHwjocPBOwNJRxkkXl3q2WO1fc
wvUL3muFU8P95VaSyuxez+1WrQE9OA2dDeZBja5zWH7f3RcUFvWr9tFHMvio4ab4
QXI92pKu4KMusZPmAJeJq4ArjhA5GWrqCL8fZGdWopoPMmtcBGnQeVtPI3xoVkU5
nxHy326KWyz5Y3Wgl19oqrqR1K5woKbgJCf9T1NaIY6s5KRLjhIFrtsX83N8Z4Iz
LjY2y9/W3SNsPuyVl3e3W1LdjhSU3ErKkyZmZp2hRwnpaHr/zP7VyW9RpP7YX/Df
AQ4qwICjMvotGWM/RHVY9tjVN0QFmMs+A0CfsfDdIZtcnjOomVMZ36iIZpvJdfqN
SFBlmRdxXhMmO8vKXn7aZfcvA8EBqi15s2OM2k4/syGpYcwDzUfHqwoQkcln4d08
0NC/dx/9QPunawRkyze2AoUQjKcVrURNDmwFME1QJYonZnEqDEaB/SSVfSe1SBQI
a9TJ11FMNpaOne/c06XFxg7nSVWIQ1JehUbFoNc/nTndpWFf3GWs/QZDYsQuZp8P
swK15GUNyKBqCwSGi7WNxVsV/1C/sVZSfgijtRTVdEIOvE/i0dzNEXqfsmPzY+KE
ZLPSmGodE8G9g27Ppdx+eXvfYrpz1lrpdxh3Akk4rdMLbodzPI6RKQtz44mXw8UV
AFnUSnfyVdb7fjAcyMrcLV2BjaYBtVtw4FnS2kBdV7l3vJ/mA60uCvTnlCLio04C
BpZen9xBMLgyO/S7+m2Wt79OudjRGe4dvZlCKQArvc4SgWhXCLU/k/J3QJr/Dest
Oq3AoMc0HQQHP9CnvsZVu1ni5Q4Msz8lD78UQiVe0fGVjP5Rlwe+4sfZtXAYM9sM
OKDm72dniVr10moqPkhDkWKApweU+5xHjs8xe3JyrzbjLa7TrauYnWd8A9xBotV3
IF3onA7+LZalRUh4tgLjR8t5ycpjDBeyy2VV9Z8ejzGBE6M7YMEOhhgbNMDpT+3/
2IKJTLIi/1eTDCDbTf2768kWaRW4KlWcmegTTMVhPshHMDA3fE52q/e9YgivQVyu
IJwvuub+T1qvQ+2szNhX/XO6/dqP/+JziOjL5CcnV4wyAGXKKtGhNHR6yDnN/ulk
KQhc6kAHYQERAR5PCpq+W2UBzQbs+vlddJ4yJLeD6DNkZSAG/rfwfBqM5TVKL2s3
GgNZ7O3dSxcslLjNWhyhOrmVkRpB88IgS625seECZLl2e8AajF/z5HzIMVqG0BYN
przfSlBJVjFqHcrAtWuvwC4ZUwsoECGTPKU8Q5dtifvaeeZVN2z20iAOS6Qa6FcE
ZJCLI2sA0SM8gE7jaBjZkzpBurj64fuadkh6sGuvgld3juhDjJ3r1wXJtytNUbh1
XVKqXIzP6BGkMXWx8IyLtEWuCwntnqc3j6Wp4r+JWmu53J75C6kkNrOKpeHF6rdh
Jbvq0Mc/tcHs14X90te3JGs94t4pASd6rUK5R7jxo+YWEVSAj0KVUcVg8CdpyZ3i
YNVXNJ6iGskcXqpk5nZD8VohFtVMUqB9h591mLX4mOssvH+0+ZrBpn38G2qh6CZ9
c/20FQ5/vfmkuEuMQfiPrqvqeCllYxsLmTdhXUGhqKraj3PDnvUzyAXitwj2KWX9
1XMS4WSiNTy/e4fgr011N7Ca9/DmEgS+LrLqy1uxt3oRZsNSka+lSEOiZiG/H0PE
kM6+6FzthJQZvfFTH/35fvBD/nV90l+9Nt3J43xw0SUzrfEV15fgzhbHrrrmgUkH
jRsK5+Ht54cHXxUjL9yDySnH1VGhcWYQ8v0fVUEWk5yewyyqdORmE2gN+0V/htnc
vMzEdofcA+p2dr3YKYXcReuJJPDUgjLgkg6RENAE2rNrpn8ObJiIMhJ+qZuYFMV9
bnoL79bQIlsrj0lF8Jj2THvE7paVEhoikmnRNw0WfXqW+uVZWqMN+KhttDlFO8Yd
rFpggy/k7zKsewuisELhjhkF4FTHVwlvW0sc1npMAmj73nMZSkTSuw5uuczsS91V
zE2k9tXoRG2QJ71XgM1Yiqzssafd7St4JXQaBnOZbS2YKlxpzzJhIMw+Hui4IebV
ZOr4Nn3Dk6mHp61HdG9JxXpQGr8fTyl0g2/9piNAoXoYLt1WtVaY30RnXB3d6Jog
A+0MPYztzNsWzD+SoDGXhjrsy22Vrd7iOGDlf4eyJMcOgFQmv628EcjEz0Mz+ijr
752sNeUJWznFWKPL2BOuN3Rgjr6iwLDtCUbpo9qzDP4HsQ6or8ETsxn5DGR4Di0f
GLw6swMOdQk0VvdSLnEbB4uC+H8ktKMPCM4NQbhPCB55a+la6cmqqUXBgwUW8mx3
8B43dmEzpOBOJvxfnrCXi24i+0dHP3uxEiPWAyKpe74DDt6IhYEn+aqezNycaiH+
EFQdlIaNdoPns52NFldsMMsFceioDRC0HZhYZ+pYij7DUTuyOdZye35i6x1hqPuP
Jzf3a95X/ObCLdW8gbdBGd/eUSOL+pA7lcCE9/AOa4nQCfYtZi15KSdnF5VEck6g
+LO+ukOpNaprhaNhufx0eK5ZTKYt3DM615CiLnhR3kTjdjMd8ghz84Ph42mr62p9
/yxUQwQ37giqrFZk6y1VzwCTTwxKqb4gHy9tT7eXxZw3LtKrwe9LlLrrxsAGGcif
gSPkuNZQi2w7C8WoU97itFfJLR4I2So9FrbqGO0DPxHCM2anXDVRxEooMkjSrDl3
h7OofROhNjk8oEfnB4SI+Wr4ATJqHpFtWBTw9lgqNQMfpz6j///ScRcid/b31yXD
fahiFS4LwQVzK0K518RH12f+PHwHhmLrIOoIV2JUJYguDkM5+EEvIDMsJnpNFu/Z
fSdVFbgx/z3wEXvANxheuWmm0/rPnVz6WV9lLHGmoETmhgxLYI9gPsMdcvXwHuQE
OuKWlkgyXMHV+m6Z58cRDYwmUUSmCMWJBHxhNVddB5mIV6ELL5q5uAeVFeZ6WfpE
pWkayREmsXfOvCVnStE3R2YMz3czFgtqMrWbrsY1V5xNilwp9ZpHT2kL3llr5ybR
xVWeilEcTb4PePBUbDPADfHpjvHJ1zVxxsx8ZcirCFDvlrh/o32GH1fT5N9WlOsQ
G2NgLzyrNFOMh9v1XV9mPe1RYcfTHb5SemulsMXCe5XHZecu65BtGM8BRALzm9qW
szkA7JUvnnwgDi+5ae4FQPzf5Iu0fWhTK7lExHtMjQAYj3OcOQMaguLn1xvxRykq
Nym6t/ntZX2G0JF01VCb0m0f+JyxJ/tbgVIrDeZVCIZfg4jj3nuDxKZw83IOr8pg
bCv/ylxdT3dgtVkfBv+Q4Ah7dwqgSladpoA5aU5R4H/55mPgZCudMRxToUgcq92C
a4SqjC67XdYJ4ezgFt+b1n55ydIg21xHh0bOAyP902tMA90e5z4ULE0gkl53PTmX
F+C+DeWbZViY8cnMf05EwW29tSybyIbwM/POnYiDw2n8CqGA3kOEZeGW3EcrFNs0
P07mhym9geoZnXyTogeGZcqActft93IQYHPHUU3WiQtgKpNtOC3eXqt1MauZ2I0v
rv3Jn+Grdkallu5KLmUvOReP6/lY4kanMSViLJONBw37785fbG+wEhXgQf/JMJPd
246Hn9Z5qXNz3u2+mPd0UF4i8VmhUwHY0KSkx9F3LnQC0YWl9ZBePZ1d3OYAyiLz
X8EdXA6FqbVrA/V7QNOCSsGNCk+OgMQxvKMUpWOM13fWQ7/1iBh+qWTn0MNs0+93
SesDJ/jTzpnzG5ftRxJfVznJDIZ1pVIersgkgyJ8Dl51xiIGIQQxZMSiDYlQFOL1
jo+On76JDKGcyLIm06iuoSUsKD8/Ck41OS7hOQRv3jsx1PLLycPC9cMtq40ZfffG
Yr1Fe1vQ+Y/JJdhIFLIhXVvxCQsln4aUgaExHXiOFXRVnTVcej7OYOgyWicMr1yW
UqKo22aud03eGAqSSyA+YUi7bi6itq0PVIxQXBXL256ODYbaAbOooHZQmfeWDMB/
TPmuOd7g72BkzTxlwtcSLyW3Y5dbqfw5wfueCcULon1DUUfAJXRw8A67WqNap5XP
2tuF9I6uTsDwxojkYFgdxQect+niN963UqfC89kq6Oz8mlCmG62O+rsNFMxXNr8J
1ef8eSQe+MR+G6bZiBUf9X+ZZCWC850N0I6ujr2e8eU5ny9FcPAaPe77mSruU/O2
B3YlmgVTnABKtzgxU/uW9Cc+bn7Bs488YiMZXX8oGAZZE88vOyNyfQSiGwG6vfdQ
y6TaZT8i9CEhb2dpivVfb4mS0qaKtlUlctstjY+GKtPXmx38h7REIZaznpe5vuC3
g2xLFnjfnv/H+gtEr9d+fZTlrA72gojP2OzbwMeDtoaCMx1RBmFqUROJW5wTV5Cz
DIWY5UEZ11Jy3fVZnJ5Vx+qUycWV+iSTS+YyHqHzxJ77J8+4TLO8uiLz0Oymikqo
agLn8b7+5PbC/jr/kVAnDlk42/CewkQ+jcPJrG07VWlhkSaZOuBPOMlJKmlHvdKT
wJ78Nn51v8CgkQ/mfoQd/rXhZ8tPDj3Spk3ILaf+iMx7ZjZhtgYOle+0ybbXTk7r
z87AW67X4uY1eeIThOiqtJfeqewz2z/dGR6mIVbbJfFk99+P3Qvn14UNZV+PHrJZ
/1MuPt3KHd1zXLryt9WqHhSZc1DvD+3D+g1rV0Hs4ktQeIF0GUIqP/qEfIsiB0ua
ZlDpT7hZhyR+pYzp3cX0QS2RSvuP0gcLdAxXbnUQvNfCx/bqovE06kTNqsL2vzAQ
3YIt/uyDLmf6ouhOeP+/sHI88XNyz7qGt9N3xhxWTHjiF4Vpk+WtDQyLAA5mqU0v
C8CHrUg21QyJ1OU0r7PdOFkqwncuzinFmp78NGZDSx0G9hyybzz/pj0SVk2PN9y9
4wfEkqvvaf7SfK84qYBoXRsrbkyeeFneC9Lvbn2oUeemoVy/T5dORN83MR/LjtHH
FICHO/iYoYEErtOTStWcjAFcOI9l9ixJvvnVdoO/PVAoR1LozofOq3XBnoPD/rZk
bhcWp05QOmLUxO8JduhVcNvYJRW6VAgc2qser6CgmsWsqkHo7xeYJHQgHaadkzi+
/HwbGwUPaB92OcGIi4RBpc63vA8Z/80RTrXwKj6vGdvsbS/BTI0kJqavSl681rzd
aP1k0NNfDtO1aI874sqiGjSy6NZH2z++TyBLXpyyqcVe4fkTAKXk3dvMmW9ff6MZ
qh/OmZPseuF+lGln4aiFWRsLozQtxL4cGIQ+4yzUJRwzHrBwLEL7UWnIUNtObO/U
xQpvv6O9fUolTAyLT1kbkk3ABa92LJndUBTsqhE1P/7/W53w0feTJLCIJDWdSduv
LDRj353F6xTuhW6OgKld6YkyAY3bdLFkgUn57WOGqDURvPNMT17WgbsXUJ7HfDli
a90z1ZdPfeULoklGsD6e89Mbmu5iQ2Tnzcz3GQ1JJ+EzT+kHA2POWmFSGEsKk2+A
r1yxISvlHjL9iQOHN9kPl80mcZbPOzH7ZmqruTLf8Ily0kVz4fr2adj/YgR2NT+l
MbxJ7aaQk+I6V5GcV5NHOLz+vlKGm+Td4GUoGVdop+VaCTEVlb47YZ3WsvxShnqL
1i1XzfhkKRG0BQFT9oAGuWg0Nhtnu7I78soUFXysXxH/Ex5/4LzqGyQ0lrmvxSUf
9tXrdmsT4+sDXpfyOp6SDKo0m8xMTJNV8XmR+J5/8OXBC/K3MiJ/RIP8js7SG1+P
JYu5yRXUo20EsQNxH44s55JMXX660Zr8/MCVOjh+E4etDjx/xrTdd/L6e8wwmZSQ
/p2JpCQPHqoYHIcA7zu/yqzQ/kSw13SxTWA5SfSYXVrqH+0PMsSKVRlcNBLimlm/
zP4g6wEFGGSLeyNv354oQWHY104Tne7PyKyuEz0Gf9Di87xUrUits+m0VZP6ke2P
ZbW5mUdW0ZaxVek76W2ExZYSeI1+e239UCD0GScRnlWCJaVaJUsfY1lsCwxUL/BC
cCn9iKKt8e/0JqN9JJ3f69BT4eE38sqvo8kb2+78niq6kHm2Gwvg0H+2evwFIApb
6+SDQ8CsQvVaTA8Z14mgzcOF83ygu5EcbSfpnauw1Or2TK+f7VDFPCDACYvxyfVV
BsMeTwGNf3YajQn+SfqHNymWif8OtyXDV0ocN69xGsV014AD4q4dRbjKDJgxtqP4
FxyZY89GpZmHsxPYo/9G9cNZ22pyIzXH0Q9gUqJfIndf1ER6WpKdgDCdtXVA3xTp
IYUlxYhEb9DO1wg4FkPrrffKArw9auNFHuk8s8RyecJMCBx3SdVC2t1yLfa+70nF
T+zIBvf6CwT/uNhD5MCYn8lFk1H7RhaFM8bDIIeyxBOrtgy3RefTJh7tindijYtA
DLxVqKcyymG2ZSAd7cQiAUwaeSTP8tZ0QKBIOXDNP0drf+KduvS/6Jv7feGDZmo+
8x58lBP4d1dhVzDkEBEkiey0Rpaxoh5n6IAqrjVYL7k3alBnYF3bwojhOXezfEna
GAS6FbatfRDC1kJYhrlLpjt/YYAYw2jphzNeRYeTLj1lWT24+eauN5ErevPTAFl2
W+6Z4+/Y9ozq1SHtu8pWQbQ3+p+/otCVxb3LVHwBRVU5zLqkYrxm+ZBN27WnSZJy
0g7mV8EhDQHe5S7TSVEYO/GLXyHK+xzJ44vV/kz8/c9EqTrRvAjBX6N96dLcxc//
TM/r1AJMKdIeiAru1rLMne0dCb+cY0vaYB9hRVS69sPahbrpAYNwo6P2nMwgGs5p
H+2fPkwxWyCEXG3DlIJlgihNS5tAzCPT+XzzkTaQdu70xUnuIB5Cq3891/ZJmuvL
9LC7wEnWzrLwubgExHbNy/jaS8W2ZO6vLYLI6wna4bNqD9sS6kIpqkM0L2Ypa33+
GiOIXtmyYKwwWuoVHV8EJwgFthPXdA+S0Ma5pcsA9mOjLlX9i97DT/vNAcMbozRd
sGeXDqrSfeR77v7VSO7IqCgvaDwMr3fWN+/0BJezQroSzAs/Ei+Csi+KNruLDS1k
Qv+RcRALBbdPesEIYAL5L0+SQ1Cbj9dDR0KTtPpPSUE5I6GtVEAMnrtRiI4+XZbL
n0Z7PX60+V0JVM05ier6c1fPLsNYI3gPWV73oQkRtpY9R+hhVOl6u+80QlumjuyV
yb2IoIDp7Q4DYkBcssgJZs4cTMMxzAQOlvE+NxLr+MTWahKaJQjWvC/0Rd7+1LAi
kZmmpovoXa47Sx3JIylrvXFhYDSCMiYU5rZAX8IvPl8u+Cy+E8C9L9dhtUoRlPkI
0hu+VJ4rEKq5MiR9wFCGGwf39zDYa4ILw+n2IvKPOmmus6iaXMfsOp75VEl/qopg
lhGSxdE96uI2pi8RRUSTBsMe28MF1yxKBqTqwZ5YNeNIYZpwkR32UnLKH8LbpCc2
Njel4aO1FfnSwwGmlzdvsGEZFKVwpS0F20g52zVRvLKdVzWJ11USg2Tp4uflSepg
J6ihNmwYd2D8AWSpLL/4GpRnrV3utgLff1WYWT8rrqipREMEOWihm/Y30Yq7G2Mm
AmHwhia2cKTWiqJzddE5eIarvYEcwzzktZSEcFFX88f93FHeRCqEuz25cWVxhXOu
yyMsGU66xYH1H9hLySZ9umEmuLYy+SAi52fZD9hbPaXHD705fOAm8o4SwwTbf67o
kFfrOSIa/2u6uMeoYusbLYpM/9wUu82TzWlnlcHa+exh8no0w71pR77eWkmx7+5P
EmgTYXI+v53QCJrZPmsnJ6zmN2sPpjLFbbJRp2DGk+OJAjRf+KtZcSTMByj5aIlQ
8zNCy2cTy9gkt+Fpo84qIaFqo5OnOsNKvmM4dcUBe75Usi4EiFbn/kfca1Gj074J
vS1oIdiw0905XmxxadEdb012gjvOpgF425s7nOgs7kgJAHpsw+lLaWIHpJzGM1Xi
NgO/nO3U2ZXe+sDtWFe4EC+FhQA5SN8+OMFKTTb8MOCjIXJ0lDEFN2t5J7b6Skz/
VCm3Pc5nYIq+lwLl51Dp4kFLaq05/W3eQlQ3Y9wSGhJ82+EaJWARTDFu8KoCKtrm
un3s3xYevGErf4xvIfhIFR7aTT3TvNcn0aJ4mVx11L+G9/tsGdVwhCh9KH7CsMtG
x1rm2IidGf40WbFogzK+ZSHSGNxunajupVcBgBKBZpjlGtAenOCwaxCvheCR16su
uUEXAfZkY0Yl9L/L0Ndx1GH54xad4tz7YetzSbQkXapUPwf6aHOM17hR7o7sfsda
33wP0B/Y1n/jZbL6POSp8axwWQKPqJMLK4XbT4wl2yPW41JQLGOpZniXLr1jlRT6
74zt7z8s+7Kru9cw1Tc54qher1klVvkAtCLrcuGuWleyRGXULm+S+D51OzDqNpZq
M4jY4X369ppO3++TqeIK3hifCl0ltsyNWx5VHSRr/mosbiGK89Kcebn/zZ/WXcCI
HBnb6KIcGpSHM+6pIicnGQ9JWP8kMWhB2OyCajkiF6tWMUmp+3BQ7ag3bWVOZCpd
rAU2xleXud/IxwG5656vrsVBAKnZIDgjyn1tGAxFwUXMeeIhrIKuy3QrX0saaMD5
4jjcWpbg2aHKcbdNblzGygRAX1e1JlBqxrhij9zxqN2KTDnmjQ7299FrcFxYIGv2
2pQGiZ0XvCWpxTSu3pJMFa13YaEBokjzzu6RXDSj84CJ4TOm2NHEmaF5fMuhW6F7
KQiNoynrQOKC9VXoytzRe+UMGozzu8kbDSGDxsltUpPPpPqcog2N51bQsy+htPqv
S5y5Wx+VqjP5W1mJ0HEwEIbCCPEniPY6PXHZAcEE4a5XTKX5jafipTHMHTxKDD8E
8GDFSLCBF1IcyN/FKdNMWjip6hliEmOtzZWjJLUqSE7lDgNyMG8dfufczUTJElKJ
OuOvJ11tUPhK8zcKJFBavDdk2de6dDaDsmyYyQs5l65DkDUk+faG19U2zbfiZhk8
3Qr0Gx7MO/piI7L+B4MzuMFVZFs88cdcTINgZEHip9XbDv4N5RkISyiDoFCIFCU1
S0apS0BCXlQm78RV8eurwmULhvat5D//y15hkkeDictjl5XZ8pJoBrJobCGuhEn8
18sUlwIpkSEGDBgLahc6GVV7tbar6RP25DbVyQbf8QQAol/0sHoz/Y7kkOKZRiZT
j8xHC65x1ecHq95nK6ZpHDbeltTdu5grxOY4C7iAmSxEIWhirjFshp8ppmfnBolb
IPtHgZYMdRkycBn0sVLFwiGTSMXQvOd6GapXwoTIlyqQwG3LCDUH7T9CXQH/BrDg
uN+slaAz6MlHsHeAtBXzuwia/GXGMFTzMgjcdcilYo9BBbPs7pnkQHNwjIhmztmN
BvLhQPRbrjsjNvHI784WTKW1fnnKTLoCTiT8sFWxG/kz7UjDcnuU8vx+iDS66wAD
NGphsF7YQBeBvoGfoXQIlqlX3kzH1D9V3qcrWUhC8ktnNovoG8vhMeUDaO0FSUX4
dEAegJfu+liYq3hJ1lwHezpyB+QXcBpVnwboDNhnNAoUXG+pAR0nC8J5xSMnI5Jr
EkLEgXbxZvX7VBJNy7jZDSH+pG4x9M3F6+lTndz07dTAI226MIx9bFf/IMiFkBvx
RrS60wpVoo23t8aiWYHbUe2U/1TJwTxBXLfbZATglsOOeUIfPJ+nOhKCc/dURzZg
nSBC5XATuf9SBuS63h3mGbkp4n+XZtSg14uYCuxlKLLGB0/TW179jmAl+UeCjzab
0Nq2Qwhf6gJTHz1Tfl/28CVzfLnIRv4xXuskjLbh3oH/F+v0XPeLkHASnAXtTZNC
oH6ho2B68/IWM3jq4kWWH3K7Ml5Y31xov2Gm4E2BgmZ+EyIynubEWKCQZxFilkMb
iCWDuYSNgHWfJpYAF2hMKOPAs/+XitSBd+c2ko2M+KQPiHCEraUrtrE4e7hOu4BW
39H7JFQAe5DK0GnHYgE6YX2oLEZP7kFTqVlO+gKczY35imssoF0Yet5HLkHIB3pE
dZwyJAY6+EAos7dQLy1eUWvRUraiBXIggW9llzQvB/800k1meMx7r4qJY81STisc
xaILBcdjBl2Kr/O98p/xMZ79wps6JDSZnQTEkOPgTXyE0GnvO2T5gkvPUZi9uW+y
JVB77c71YiAi7LLUu9PXLrKCvnJ7IxvZ4ntidXgN/UHiM84NdoQ13e5zZm9n8BNt
Yt4WQiZxzq3a8tFBmjRktfUjdti/OFfANDuJ/f1m7OWb5TM92s9cIGkVwifc5XMB
AlEpeUCGt/BS9b1aOsajOJBxNpUisdTKtVeL9u/BaOUbhEn0ekUjYUlKAQtwMQbx
KGB2ABIf7hXH9Pk5sjmtQyNGPrYW4NmxVSEkvfaaiNfgi534v+EjIvwkK/DX7o6l
v2VTujy3gJgi4Q8Q+h757+ujP95LGg8Aa+vGL2s0dWdgnp1TE394ozMnMwuZdW3Z
RGxWs/XJgRze47m6Y15LH0u5NV1yiEH5EIgdSRbul3AdQ1wx7M606/wF5EaLhAPv
2d+M9Bf9DVYGc4LbxsJqbQsA9Jyv1jIXs/bcRraXgpEhkdvH/doZHC6Fygb2mB0j
ipsl/4jGzc5yEMwQtQpiSvnLLYHVUoymqr0mpg8AAomN85A+PHuaT31eYiZdKoiL
k98oIugFDHQGWSraXka7R0xRxBdsP3iRZwT7LN6tmlD7Edu1/pdWJa6uG0XSP47n
qhlKBV87tHHVGhnTBGtbUFYj+56CNjAl0bPL5hq8ReCYJWEWo5b9Xg1vOfYbRUOR
Opy55K++G7mLXYLkLoFRmHp4ZX/q1wiZufUqBc4LIKwlzr3SKf6kwWeO5LTjB9L+
YodR+7EMpfSdrDIrXJIbJyjPxG0UWJjjNCsOTnizD8D5TUgdhcjQjQfyAd+fbPG0
hOBjAH8uHmLKoFdVUxVVyCH7c6aDBx9FprQ428k+7dsye48538z/kf2E7DV1TdII
VF21sMBoOTZZHIt8B6314/2OI33ByLpwmDNWx8JsHY744XuC2kzdxOzWYde8UrtI
XlZ+/1TtMmh2eYG/zRs4oOcPuIfHyIyBkbRqmP/kuI5kNRNRme+mCKmUkS4VjHuI
6g/mkfkdL9PC7n0KAQFdMe0fGmjX+Dc7bT16GbceT7O0TB8hdHiPTCgqzu4GB3mq
wjcW1HC+ZEJMerlcOjfwYipdjO/TorNkzThAspAy34vK2Z9y0rQ+ji5muMlNEknQ
Z/ZoTJq9smwuCJJ2s3ynyRj7WCYGOj1MVzI78KxOeqr+LTcl6mHmE9shyYVL+0cQ
UkiowTu2iJEyYrsnujVUpM8SRYmvL+GGdH7H4Sc27k/CtgWJ/NF3rVWbmCU9v4sA
Kd+o+8tKBj9CVkIMw6IpofDAer4DpMlGSgR4+yGdaQejZlgJF/WhHcTlFLnU5NJ2
L08xKDz+EFRICfzozX4OSkVh2tOAQiV0fGwIQJopNCQNe06LmHRD3VWgHeiET3GE
DRUffIPLJjHmAPFrrFnCaugJBec9SKWha3w+HIcjjMCqChY8p83Tg8FMA5KLLYjh
QoGjVpeqwaYRGDWIaqPcatp0Dd5eVouZxEbe5LSn6Wej0zS89sVpXmilSuefEwSl
0l44Hbd18YXCTI0/ziU4/Nc5mrMAJ5NOXcPbl5B4rJYZZd1oG10mT7XQ8TlMufj8
ZCM3Wbid7PTVszjAKwavhAltJLMSIM6mufeb1s5fiVM64zrTkxzwYPla9BOtfG0R
biCo5MlV6CfLeapixn80UtbU4PGACd04pX/ZiD0Z6bhKsBplxhR420GFgqF5uRAC
Q9SJW3Y0S136FNSd7mPBbN6DN5NrzHYIvhx1jWynw0V6I8PrxelgdJ2BrV+ImdDO
gkPWi5ld/0Vit1FLEXyXeOD5i1vhMivpn5lp9MGvQ9cGasIOyRtOUqIRQzBzSu5I
gakFS1kmDVLiXfFV83/wr/+uZ46ItSC1B5OywxUoBIU7eiFZQay0UIJX+gdPSLRC
BRh/Rg5iBSW3E6SlXIgUVme62Wn6ai/phF2VSNpj4WV4I7/isnymZwkk9TKunXD+
8wE77GceNfBuvFICTFpVBkCFWuZ5GMNjZCU2+IMGvOXeWF1SBlBVEr305ow1Aqqn
1LMpEQExVibm+w63E40ACvncrGB1USKzF0qTQiKfCYdqxXxLTn9r6SrGcI0CbgLQ
3TrOn9ndP1GbI1OFAndbQgKRryG7HVCY9GSCTvrN+oi4lGO5DM6WjolV23m7LaLP
k9JvJvyuX+OQe/0kMu5M4nxWuFeC26ZKUCMR2Hf3uRy5waB8dn9qI6VCSuOFsKYv
L9Ji7tCVBEV4CAHOEY7Bmk8561+FYwBc01Sr/5j8dZPRb2EgvdMcMJEIr8ZpQVV+
ZUVHRfLhhhXLTSZzbTwp9f4dGAMasSZAItca5ck5wAWlehShyrahF7ZN6pEEA37k
TVVs2Y4EJtDzLXvqrdtiY4B1M2X7cRCa4olXJdfCwt98MV0wynQS/K9CovLKkICv
/hs/Ve3dCY6ztSbM8mHRJpdIkQFmRvB5B7+v1ySFPew6059vC6uN66nWxKuMrMhq
SHK3dxGHAOjLDcJtaaRuIwwq0sqkh0w2iQLbaH9VdfJ36ampNUUwx2hjQ5xrPrHT
ujER4HUtrtGNdL9QCv0o6y1fG6Dni8LiVl6rbVyjaZFZompgpUWAPapk4IjeSB1x
d6PaWXZcq9WArwBDS0hTdFiN7Bg/WjZeS3A1tUaS0aO3NmrsrrB8XRvWGYW6H0EB
heuVqCDARpDKbEy48uwwWNzzn/3QBScXQQo4xVIc9Y8od+iRhTtPGA2jP+jgwXUm
3TlMDh/0ZFBqm7GA/ZORqacQIwYP7VxyJJ+ukUO6Okr9BWMN9lWoA9XJVqz5+4ab
e7tEBtXgaWksYkdQnU7AJYVbLdqmrSdAR0PO6PoNgneVMNlLaHeB4aPtmPkyIkC5
1e7TnOF9YL9Vr3g4gEBnaQVGlgmFBHgfPntguXf+V4/3PfgWEQfIhRdMGS6vZvEM
32nNEq3pfjz3ss9IIGASYckt4+UKa6UHpiGyDNdNgmPx1pJ2Lx3RYYniU//DOsmx
ZBsGCCwflVdWbUz5Yrxcb44eYO3WXH+lLoblU2m9zgmY9kGHTdoYyToLpIyMAvDm
XR1tZJyxzaGAOKrx6ISKvhLjafgzGsUhmhekq0E/QCSgPPo1rFk6cJuYbXTUbu0A
QZdf0auyHHxKuYhx3Wcc2lDLUs4lVdB9X3DJ78Ewx82kZeZ04FCzOnhccmjx7IZ4
xz3b5AD/Et1PohwgogxpM2rsah2gwv9QoZeC7TgPrmM4wDZplARgT0QfgTpG1FiX
pxBDj9tjcewV9I6AZLjK2BA/PLbi2L5HulRFGnRyPv/Yuv8wcIPykgXtYa79Ndky
2RP+8b2lb4+FwtbatvPIuEvZ0LgGdMIPC3ZDGAPs1iVdjY6jofzN2gm2Q5zZsCv3
ahMzItWucTYifhfK+xCbVozMKnp4bB/GLbSzO0ALe919keQKOgeLypKsrW3NpMJZ
FrJuZ/4FMKA/7F4rfCYE8b9jsGKMwxOITRnZ6/P/HrBI0QRqAqXeke43oT2zT56A
TYzwen/9LXAQHpURp8eZ81TZfBuiiE5YbcL2o23XRvhYUM7x4D2fWtlTRhHyLA/D
0tu8+lTrHXyu9UlLvq/2Tn4BYanha3NGDYwIR4TXebHaDDvRdEPFfo0dLQdBnDQm
MQHPDn9Upu3BkT4AGY90IAbdFkrbjSHv6lM+0OlMFEgAObX4pUTUNx/Sep0IEvY2
/cMpoAVdndc+b5hmigV61Bt5Ol3TEVMeDXCX2jyDXBHhkdUoQNRtrz/FPKWS8Fmh
QiiOnaKqRYQDDrRRGjR6iswDzS+h9YkK435fi/H8raoUriiiQVgdmri+p73nlTJJ
74iSRqA8KS2lWwn8++xJMOUWs+v6ARxeqbMXLTQCSA5eLNMJwaSclBRs1MFi2j2d
CLr1VXbQZUnfL2xN6w1EJSuqyiRg7bKBXTQXlTkpkdT97elG2GIxbqP8JP7vl7+2
uujxQ3r+Hpp1evmAKSvc38qgRPiytisGjKkpijmaQdkY/ExOamwLfQs2CbBoj8RA
bPyqzfIIgNA0FFMHhkpLWcsa2HHcAI/ISE3oOEmC/0jWY+rQS8Gu1xwCSpaHeU0e
0gxGK73fbxus6itgtvs407y3YVLj25Vlvf5TGt0NbnzYx7FV/HoIB0x92X5+vo8X
ZDYGDrkUIf5sdVpH5dRXnmltnzXaHM9T+bTJZL+3Gs3wBR3iYKKwCAgWSrJkIuIv
A1wFT5hA0d5H13o5L3KhEu/9DM4SW49VwzijG33W6I/1H9MXayrlFaVmVLI6QZwH
PYxBgosvH400W7/Sg7+c/Xg6GtPusWSIWsL7HLq5KBUz03CS9yRnXyEFn8ouQ6EQ
Q1EIjimpGTsoC5xrWJr8G8BpiEnCD7kM21MnhKSXhsB0IAYWNlV6mhehMxPX3jNK
UXV6RQeBFtT11U8j7BwNDoAluAG3kGFG+CloimgRVZCZtdInNQAB8iQzt1zKzvuo
jxvZRMEO31dqvpK/ay85VZP6GWscRu3/5DHB80vlKOl4vVanfBrgrCav369OLt9w
es2MJJ8u33TpulC2sY5uzGFibzzkJ7wWcQU9rrnhw9FbT8kcZ7GMttqGB3evRUtm
Ue2x0QzI+dvMbw9p94YesaVQkszAnP5pRmag1kcd16qpal9FQGPMRHwTVXSf+OwH
lNt5HXj0gMkCPHth+a+um7yNkUwwm6zaAGMcy2hENg2l0f7zpnx8NVJFlnCccX4S
EB33dE9qZZ9GIvryzJaChyyk0RnL8G3Zi8kDcWjTsHSvHhcVVyYkNf4FkxO7ExyG
eLxGFKjjxdy2DIx0Qrql6esiQUg5TtRl9zPB3OnL5LqPWGNpL5C5lHSaCeA7TBGH
C6BngOC7yA11QotUdqyBtbybRJuo6GSEMaBANsZ+FceuklvX7kAs8rWasBQoVVp/
0weKxYUTPuxGk+F/OjRA+ZstplvA1pdaZXDhVb28K2sj1VPA9acwH1hfGHgtq4rJ
rc3ai9VQT9/xJlxhRuvvkAYWuS+QEsN2ll9gV94LBjINYfb8eU/KbDy7MoygUDh2
yYf7gsTLfXZfnb2ttdyW9OFTwrCEqGZUjze4ubMfvRya76TvtxRuw6M8CYa5+g3e
jp8pFhrUWXZ1whSh/gpA8F8siLGJ9/WtJ2QAxI+PHwPDJ65hdj4kuywzj32oQ1C3
rVPO/5PcuPISoQAzyjBpvmUx9nW2zlwFz7vw3XG66iUR5rQDoCf/T+Oiaz5/zCyi
aXbHwIBQD0GELrAVxRiyHlpdq61fuw8HcMB/gMgPtYgLa3ZkqL8xYmzxeoA86XdL
z11sdIgkj3SwHrw9X2+7aobm6uoSXYpV8BcojNaKggpnH1si7TYWzuxrrJbKlYOK
YMjmjJrsfAfTVzmOf5M5uGC4najrPH8syHYYm/P9GwNAWE28+T+98GhCA7hkPMle
pU267Fh/GKRBvMSrSgWCBxeRgIHveN881b5T+LqqTnuFvIPZYY4C8jRL7RFsKKzf
WZum2GSs81MWshpkdhSd0RDBZlasCNLNZP2cL5rFgqZyxhmTeEFWWmrPil1WR04n
RV0wfgIKrTvbS0olbKgzmsCN673FxmHQ85Nt/a4FoG41T7CUTqM7Le7vl2b2yNRv
JG8DnLH//uEvkGfk2ZSh03WdNCVuYX4u0IUFcInpWKAcOs9kGoilv/Fe1tvgLJ1K
wXBf+LWNmPdDKB+3H2XHvsBFYnenpvpMaaXdD9hmOvzkK+JkAAzteSERRLGt9z0G
LbU/keN+c+DdUV86LokQd5pwAOY1+9AYIew21HtWBEJp9mrX0+Y9DPDq23zFKogB
CQ+JYFKBVM9gk52hs1FiJm5K928d8Nwb2A6PayCKHjbUq5CM2Krr3EL7NiW8oErO
tO1IsaHNBbPKMSlMfwzgsoI4YVHN/17CN3xEtAoTJK4zGY+6D6jXEW/JD6z2jYgu
SkW2xdUvsahj7MnUS597jZ4e2tIhDNHQT00ssO8Krc6RTapHIC9SupeT1ZeyUHRQ
lAZMYSImTObrhdYeekI3KerH6KPZtuK+APSJCZEiJXhy/nO+KLjWLHPgM03JwEbk
4rZMuYZzgBDqfm7qB5Ymgc7JqPrFZzEsiytNUenwo1vG+toDssG+j91m/hpGEmko
jECcKw44jCpr+26En0E2rWG96jrLNDlq0BlTzEuwz4FDXZ1e8KTFZxI3LvVNhybO
eyyVVI2M/YSLUU2YkVgQ2smd61CiNH2W4LypG6gmn1mpjTpveJnsPWeGkwh0j0A8
oUFlbut6qu7ASNTH6/w3BmI66hqHCDHzmPNX4IeDjcpqKrmNxnlPR0w6xKcPhIKU
itN+qxaZ3az+VtHXQRBUa6mNhgE9ZhCcZdIEyObYG6ylVDcp2hxa80REvdsZwITE
sYBvxX/qYBETcLqF+0nTkSREl3/J1PAMRNusupOJEz6bQH4iZT9VXyOmR07eVVqv
V2k3P0P4m+rgK1GPlhA4Adt7mXJL6mp+Emday3dMKqAXgBlqmT6+vGl1xf/v8AM7
a6dHcxcxGR1NnSl56u5nVVLMQp+hMq3n0k3UAsCIfQ0I90hAxMjpUIhHdmK1PtEz
A1BgNUrSXgfVM61kiMVytSeI4l2OfI5/8z8YlM/HJqgOb6uMBNDFKKZ8zirM9y5m
nxiRiOp6wXAPeHQ6FV186Cc2Y4qXWTQE76HhcXyQxZVpUbP28QUV3M3T75ZJNRiy
Aqp7SjoPmUObpa/JVS7qGv5n07WtuXi4SeSYkFqYiUflerAnP1ljc9uwL/TjNDge
4UXBhigofUvN53FA92Ap2T4ZsJYmRSSv3X3O3MSboGWRKsC++F6BUgQ9ivU5zU4v
H/SGjNPFHLCX1FqmrzdSWEG7OrYrRu/H3VVoTzq0xvqQZATiYhn1qN6S2CpqlAnh
5wxtOwwG8yJ6ssvq0fGqowrX3sHRX8dAkto3MblgMJ5IgMuzLt14OCbYaGjQ6T6v
anfpUfEBF8iWMOQ4ow6ADG5ClOdWFYjCfRzqR7w31vA5ArN6sl8uSvdlZJTPdRTD
DMbhUEOQteQJn7jr7cWCVoxw4i/M0X+Vk1NGT4HVXy7v5ynS98lJOFMXm9FhcMq6
LeJE7daT14upU6ELHEe7DBOecLmZq9nITzT0hZCsDfBMksuvkZObLLyxBRGS+I4m
98LJOTIpkdH34TypypNflvf97m+ChEcympz6T3D5tJxJN7lg0LrisajBobtxQ8Kx
VZMPtfPscih2/GLN3n0Q0QVhqYoEDiBo++1qNn11fco7OCgB7SIGa3VOvEJxuwHZ
jtSSzJ93fLDgoYUuoINUgykz8ceOFyFKog8K8jmdQqiFaWeprcUQ3WsFBXyhU5+L
8sho5X+JRiAdbA0DIdSPgYt2JPuSIx2dmKlCWuKku1eAhQHTUC2W3fpfFZ5qHewH
aKrBg9nVpG+ev+K5DJ0onqIwsL/9v0g9UzqYFaE/KR32cr8Al0cTCHV6bysWIioi
cUcWfKu5zxLQEwMXC2jl0gWSjKVJenyeC89OSr2Z5o9mKstbBW11fITL5Xzpxnkm
7X7gCfR85ooxtjL3QOgWY7eE0JjwJCpxf8maxRQQo5S0WXI25MpsrZKMdFbeanrm
ZNKluiVV6Pq72y4vE0vsf4NKy89Phv2eAEznxq4TCIFz0i2ljYXDvtEaz7DmMgrB
wuoI1RN+Ioi4laY/Q5feD96lq560iUTrs43ggIqduNSulCAh1bahQljU4QgtZgrL
sfEl7fd3I1oIWLOu4D0YUzb6gPaMPKFj1W8zt3w7AxVzZBIcoRxt8C85lyx+XTMQ
EtIKtYLffA9nNCChOCT50Y6juoHjkNGhIj4qh8A2HuM/Z7y20mQ3Z1xwOnbaH0tm
GxxVWqSUG2lLuvCSp6BB/WXRpnVO1KwhtCXbXvfPh23/pM3OCHk+Yf+wC4Wnw9WY
DS1bWJ7gmb3H0DHjdwG0udixsb3YpaqQR9jQEtCR4puSw2lHMBT2ra2moDL6d6QR
TCxxq/khlK0pMtLyhKr05RaDuBFqb9mu7tsBjcmggMJxf3M16X1QeX6LjjcLNmVo
dASM3/QuhdHoCBpssHbv7a4kU4AJFLkWFQ3n18GLeGQYYi0N+hM/AcoROx/rqL1x
y3gZ3oDnAKLmJNO/+KK9xlGkYKPlPqPaLRQuJdCmHKsz7rhz018Bnv4pbHlAzHLa
ntmIaLmYwtIIBwU8R03RG4LVdbdHuiTdoLeFD/ohSL9hMVxywQ1I5FiG1ieRljXM
hl6kiNsIogmcaM2CwiwZIWnoTjwdASykbE+WSuU/oE5lzbaP8gFbYniGMAErt4ol
i9ThsC00HcxYYb6F7yLx+2FvQ79SE7XPN6cPH0xjByxUSjXIhiLYLVSu4G3qjA6T
6veYb/iGvc8bGLfjJfvnKKHnP3V+pUqzDWW4+KLqfF2wGzJkhzfKQ7rXIoPlRWX5
dseTnF+tdyCJK45XzqK5SybVY82SDBjlmhhZbVCuEEcxbsCAlwjtdYtMsyKWZCni
M3Trf0B+PIvyQeevu/yk+U/Xs35hG4ZY6egR3zSwOb8hcXbUmm3wYijp+f1V/xZg
3Ps/U4R4tQmGY2TPKeOrK5qr3np9pKmZIRtW0s+HzBX+Sru7a+YK9efz1dztKbH+
3i9XMvFnviPRTVNvicZd/61W5l98PZ1qErNIIfign3uTPnnHyt9Viz2u0c6bvFiv
dmcdTXAt/Rvfulk1HEt84wZfwtTs6vI8CFOn+Tjq+MuUTh0444Qjo0lSujoJyBBV
aNEtjjSb0FPahfmIaGHWca4rj+zbYvtc8ADAoLb1elrhp/Jbv+P7FJkzULwisZel
B602kH7V4z26o4LUIMJsgxXtUHHj5P89LW36feaxVTQwSzz6q8YQN8CYUEavYFNG
b24Cu0C2nOXWyKgr/u5ULw2b3moTUc0cRePzSouVrYe6jyitIHJ2BHW5BlaUo2cS
uOsG8Efg5z7HxxlH314loTfwfi53u3XmLkmRBIesGa4eihFxoTmmbKzKToelHZ0j
57il6uyU3VFpJ73gkm2TEm87dD5Z5xa5HqvJ+HhRRHXATaynd5/1noT/tPdYab5X
nu/JuiPSDfVbB/rYNUVdwmTzqcvxwoKuhRXDP/0Y48wvBL8CwBUghSEMltlG7a82
RbpiXYj7UwvvbYtIBlrEiHa8lsswq2NQj+NRxWasz//TQeLCFo0TK67wuqMug+Cp
PqjbqiftCvNfLEkupHdZo8nswVIYITkxL8nq4leEhwsA9Ihd9et6s0QToXvdrD0i
sC5dDAhWu2CYrjKT/g5QOimT4cifJt35dmLFqP6nFwcbIzr8itUPKvoTI8YhS4Tu
PMIVV23XJNTvyxitmsvXr1JZqaY+hy4JxMMEGmt/mpClagb+z4+1mdn6ODQGLpSJ
qrB70Zq0qtPQwuaP9hcZl0EAEGzyiuFi1oRQib2Fy+5n9/KXB3xeWUtGVslU66yr
1l9PtUAaFlsp9lz0g5QwKQVSmaAlKbkW6EKN63LeCQ30WzvftQSatUJ0v5/AatSt
bQ0+1CuzuxJknePhscv/5FYfhNJTjD1wGpcJ9GDhYJDTzt1GSwCNZgkJXWNMDqln
tPAtv4FjcS4vawTENJukwO0xc8TCZXw7IQUle2mSIR/EKSphqhd4cjD2u0b8sOzN
qlj/omfTIxEsXLdm8/QBUBQVhRySkVF1mVq/9lbl4iwXe5rBsqDRcO+ezOiMthpA
Eyt3zFi6fhNQR7QDHT0RAt+oNv2OgAx5cHac6HD44HmL413w65RosWBTrR7jqRJX
N5tZuD3jrA3xuoKHWhznAcbUsFg98OkqYGJ5wB5vpqrGdj/IyP2Yi0dpYw74PnRb
LrL+GaHYZoz0DrigBcLd6F4QpN/tR80b21kjPd6KRKsFI/64Bdoo2zviyd/4MiVY
RxkG6G48mjvudwxhRk5ZZ6iSgsLvq8dZbaa5EaDJOGZO/OOeFelnXGf2++VoYrJD
YEgB6Pt57GvioPNLokScn29Ygg06tPhc3t4s9ePyxAo/At84arI7+YxHFXEj70H9
Yz//XsP0NVm1sQi8E3I16dm74JitxFvxpLF+VJGAZkgHQXVTjeVklZ6Tzu6Ms+ky
N9BMadx4FtfYcls9KdYEgJ/Kgcj7NKnP7OzIKPZjGXvXq9lkkUq2IjEOBUZgTqo8
dPYqgIRDjcVRmdfa9/g/0sQ1YGPBpbGj6kBd9Zni4/pMiC32aqD28NuefHGS9nUq
0egCSCHVv5NEn3GH2a7+VOgM7IX0dX845a7bsZizCoj+nHWN8UymU7d0rswgHEzR
AEpqxtqFKW35yAvDt5c7cv7zdAamCTaAvQbYAacEpI35xnZjAWuCdpwTnSVAWXib
GuLGMdGnXhmRYD5OZRJUDCu7uQj9QHeR7bQFNKHOISkSYJy5Q3Zylm3348CZPZl9
pRTHeg3i+G1+ewXyB/8JlmPsl14tpqZSQ3O2f0dn2tRtE6qEok16ZpLF98ZD8PO5
jk4R/VMN+rzcJidr9YDDlD6abLb206HX5InrYCKMB2BR/Ou/j5pBZXo+w0VSVFvE
mJVxU6vIvEq1qnjyhErHAhbtPyGbP3MDRG//k597n3Cr7XOrIE5JF6X6ZE1JGtH5
eoVmfaKECwlVlGmDDg/uFOGcW1vaioMsQmugqRbR/IaeuGZPxy6YLxoEvVRbg48n
atw9vsdO6BUtWNB4yB/psk+Mc0Wga+yZGZw/opWsRw/ji+FV5qdefqtbkBV3UWGB
VJEyk75ATgTzlgx9yB8LhjwJ1ONDhnBrFKbnqvDptLtS90lwOtSc/Elu1rvoBQEx
eiwOrnSsLzpe2i+ArOKmax+S+MsrdOrc4OPWUX0++QgWnnCEDjFp5vwTqek36ri2
mWQGiFK4YifG6LUsqv65i0eDnedtrXkPiJZPIrYs5Ffad8OSsPOyr9YmlgKHdN04
UxSuU1kWUumVxteP6sVWRNc0hSUHCN5u1iFjYHfaW12E8VQk0KvJk7wYpVB6q5y5
0fXtoeZDQRBh5K3T7J8mb4k0r7GPydYybFx+Jf8qvBXmEqyZtmemfoxKyUInjn73
cq1vAvmNapue5Di+tcC7lzyeW6QyduEklpR2fap+TMvi5J3p9h1CBOUMlheY33QI
A+usAui11ZttMzU3G0172MX1Bx3cn/VbBEpyTpXscqrI9B3lq9nzE9bi0YzD0e0W
jIzuWmIwvR8WUu9ZSKMomGkGV/0S57+ZfI1geMKzqzkQz5EglMEPz+ljXSrpBFZc
uf7/gpzHEE6Zb2/e7c9FYXdZc7gZCMYHHbT5HfOiXvkUx3znF8+cpB9EFKYf6Imb
PRE6K6K0qvW+yrLHMaUgj/+IMdVEfiRDufWhXTF+x0NpOuUHzAUle1q/RZBl/6eN
L/YKceitSeEA6T+LFbyONIDH5NuzP136wnnXof/7Q7pxQq+JWgfFXfgCFh3GVDnf
InyDKBK1IKCrTMcYUas1Sx2c/efOWBWhB5CwThgvqWW/95afP0AsWNyIjwJ8jE58
Mrr9+3GfbZemjJJsFGl+MO6BN5umL4g7mQDHAITekh/eCac5kXyNMYhkLW/HeWTp
HVIROul3qlC+RTzT9Hyy+kwtlzYhUbMnCPjPQGjmI70e/nSrBu+xGUJUIIHeR6aX
Td6dwlo46sbYYmm5OoT5hIudG5+1O6s0cLuUCcVeeHjZX3zRNCvsLYsz+1lD/B2y
4OtczELTt5j6fA5MMZTOP1SC75WR3ex18V8YDQ9wer5ZuIj9NS1IR7UEAT8DQYVu
xZT145oVvd/0VYyt07HmwGRp9rUH0683DQeNMf9ypvTBUR9wIV9roNI7jU80EFAs
mWPYegs0Z9JF+Y8lWw2lraZZdzWlDxNcpbNQgLLDWMd/xug5sq13uH6DvqE3eBGd
Vqo0WgY4N01yHe423rEIj5XdBZHKeGmqm/N7A0XQZc0k/yp/SaKaFwSftcR6CbCk
bBRhR26H5tMo/V5TNSPjWr76L1yP30sa3d+LEblGz3S9gBpErC+cuByuVAw55g/u
LXi3VzjnsKyrq7j7itYZ2vGaEofZM0p5mf9oktomsMvvBwYknsGg4mjT7qMms89n
6oxJMW9IFlMkIXKsTY6mHYpl402+Wd6hEKEpqyhOWe9r8TyFFd175FBKNsz+topC
7g4Mv08SX4o2Ng4CFZGdPQV/6elpUcCARRCDRI2Rp90u1AajH8bU9h90sK2BzwBP
gw9Ob3Z9kfesa+3TfAeRVwW844pRXkZYYDvXh7sA5x85/I4JqxtT4yvd/DJY1q6Z
iNpMPWnzwFZpT2Yf/E272+mNi3BU/JHkr9jyItNh2Eixvm6NxW1QagAEWw7mmeIa
XH3HlAQ62+JT/DiTO4ZLklPK/R8NOye97Zms0VoiPMqI95j3fSoPhZ05qVk4DFiF
ABC9GcvIeBfn2iFkYROjHK3Ght4Xsu0n6qaXhlZLgZUMp/UCHj33fb5Ed3vBxv41
5hOqnl6gEv2uQQpNAxeBkGq2/kPpMvzaa18JJ5YwfdA/LUSw4ba07cETJWveQtlo
iimD9yn8kQhLHUDeVkIR0moDOAsXeEPTQzV6WPEW5gi0MEAxn1QVwF5jFBQGYzpP
Kv4EYzrND/KtgmBd73pQZvLydG+zgUlCe5MkCR/3ASxfMLkb9kIyGgMYXBDxN2W6
kIGI8vVMx2yrxRzzGCC9zfesOp14PwskWvjIw4Cr1q1RS7QmvXZ+uGnlBo4rlrXO
I8DxjBUvixLjRK1BY1RurDS2slN/U0t5FC7jqLwAyzPUfd12c5uAk75fehVs7ACJ
N1RxMtosIiCIoARFPA4rjKi1Xc9ZIa8W/U/eAQJk30qvPJ/ArLKo4kcOqU52csZ2
2wbz4c5cl3/kuT3FK2uzmdZaIyiI5o/PndpteeHV1j6UrHonftH6seE2ZTDWTU4t
vPtFTPVXhX8/SPLEcY6KwbFIFUVmqhUcZL2fHy9PUs+mfVJgHpDVwZyIEy/ojnM9
08xgbnfm1shlIqdPDFvMlk+12ry4DHtpIzpbcQuTW95tGuXHag+robtmifOCIN5L
SQEf7KzfP8BsOc3L216Q32fTnS3ntZbdqQxwxenPgg3A5VkG54Nl1ie5DE1B8y+p
ZwCA3y2VV0SqqqqVNR77dns9ohbFld7piRaTdtma9wu+vMANTBXmBPy8FhokI0wd
yk2qVqdEJzZCc1GSUQPcE4WSn0ceSlybdEz89kgQ5/RttY6DrR45unG3xngWOh87
YCk8plHSr6IdmzXFgJhNZPSR6c9Si349DOKy3OpmhN+Wx+zFh9MGXXcu3hDx6QTX
w6JdSODGBDkj4n1Uxho0BnLog5LeVF5V47aMk1wx8aNr0rcLNoaHopD3vBKCVI40
IDL7qvgC93MFTVqcNKTtMkwr+bCPQEvw9vV8yqhY7kyKwMWtInbWVIUlugrhzQ1c
nIvX+64NxDBbno7ZZYE4167zZ2C0VhhdHS5iuSNpGxf6ehWkTXEvcqM4q6LbI1IK
REn8rlyNLWzXv6rUXEluilJ2RMW6XclYlQiPLTdgfV15NWdDw0qug8kvxD3jL/cH
lw2llcZw4pmxktqTEW8votat3yFRslTH3m1NNW9gEXhmSJ7KMMPcZ7Er1smXRM1+
UPPj6bffRIIfqTIMZquAjiQq2a4Ha49vmISgRvNTJXm1vHLO63dGv/mrSdFjH8fD
ClD4fhp04TrV+rxjgxXoEw1OyYXhWWxWA7KGXIyPq0ACpkzv1D+6tp5Db3h0GNCt
TE+rWl6uOUCRx0PFei5D0tMZIZqIZVY8hnzp+Djn7poyBkA0ZpVZLPZ2JgRBvpih
dmvXYYEwRyBOeR5Fdojae1zTOcNozISMEoLi5jblyXcS4mhFShTjVGDwbs1Gj1mI
0kZ/tr5nNLiHTrHKnH/SZFETVBY+Vk2e9ViTzrzhUQP01KusRWdDqTwK232SmBXJ
+RDXL1m77rgs0O7c0Zmii3QGLx2yhl5CKSMIGxPhD6CJYDLtPxdWq+iTLrsFFgk3
ojos2B64dgHFyQhI48rnvft7OJW7pvdAMRk+E1gemohbVlKFEFqsMKNmFlZMdUNa
R9BhV6sTcGYkKuzekIU6pV2o8TjAMnK/khxl4J/umVBPMS+t7YTLCSKna0QDqOpP
wFm6AYR1qQR2H0gWTBeyD4sZwjthxHLDKVyxDeF+FHl67g4VQi5dOrkyRKJjMPEb
3lvtJWm4K85jgaFqFIvJ5K/WEfYowF35XAgrhFG8O08Hxxfh8Ny8fiE1wj7kRfZS
MOHlvuS+sMiXCTDmpv7zXnAFCk0sXXuWg3mEjvbJmQovhFSVVxdWsODITOty3xjU
616zPhMZtp6TVGWWPz4NLSQdtSsWRbZWCafuL2pz3wXY/Ib2yv7vrJV4RV2pp8y4
VkhKo9rAK3WWZxe7WVtcnhBWoJgTSzNngnzXGnBpVyBi4G8aK07wpoBZZA9KVdOu
+6unDDqQ4ivyxitlxoHTPxQcHrg2tE7v9DsCYMHekEswFValwsAFX3ZSoWFyQfTE
XLT/Wp0XHd/ggRQgrcTXsZdc7bnWYE1c3i3vxwyMH0P44jk8okxeyKExzovzZINm
tJbB9YgfTSKuMtB0ugd+7beP/LMkC6vBTen6S9zCZHGkSxyaP0aKgMytJAl9Pxzt
wHC/kg5OMEqmtta0Dr1DruFl2AS1ua7L6xsi5Mnf/MJGbWKtx2mFFnX1+w3BDD7M
B+Na5j+SDs4xyJOK84hN6sjAsoW+TbUKZ6/rwOZ2x8njsdKhFlL0loh7tFoXFOi8
qANwGZBA59PV3XLvkzUYrqs6zOey5h77/w3iUnDwX2C2GtDfYJN6WPi5DuRB3cdU
MTsXmDyO5SCFVqS0RY+vsOO02cAm6h0G5Z/cTYxar7cdFF/eZfNXP1vCqGb8EHxV
v9VpXmtLxpk8BwW/Ks3lht7CA6FIDUlRtKnKNSAPwSlGLe1oNsQk2AYbZBpGhdoE
VH6UcwDP8Z5aL1isQMckbdT2Pm/fdrkVT40R4CEx2xv1bC/lAn01NxHU3AclRgy5
Nxneds77sZ69ZTGa0Ubv69nxuBHKKaX0DuU5yEvwzBqElCH2J3IdTZs9FjypAGg2
fC8c7KPRcBx3Hv8YaO0mnbuarYSRtiVPNRnr2ZQ8MV0KY06ltUkxq2RNHf2LoUbj
dUcUluo2i3Vq5Q8u4Nqc+tUnLjaASATcCbKAoTf3IGdpS/aKT6beR1GLJj9vbAtH
x6AK2vf0glirUWdfR4TtiDZhoQOc8BCtSYAyT1pvz5zkoLryDbaPINfwI1Aa609L
Z66gHwSO/w957bXGiVnnOJc0cKYDCgWixwDxVNk6K5GVZhp5V66S55pcUON05SEY
4awC5cLsgEX4diFQfvg0UOtLk1X4uKXMvqOBE9HVb5Hgh8Z9h6yFbX6o5HaBOCJI
slFYfbIjjuWliL8h6H7H2sySasK96teNvTL2Cn5EKmM89wDFNPXpKvuad+sNrnzk
jhM+w31d5UuQk0toHvlUqjOi4jbylW2AH3QV8b3TdtOf36Zl0RaBpC+rJ6w4oiBs
Ck0mMyPwUmh2sSoCrpe9y5o4J8EvgaaWoRp1AH/bQswaxMziUTJj0YUw2Rc4j8HU
MsEKYBy+uNlX+blIP/L5zuPvbLxVc/MnJVSQLuG9d2nktewrkVaVt8UGYUMChIWK
w0rqRwi0lGUKgxFx6h9ED7tMJXe6MQmSIyYt0j2HJ42Sx9S0xxdu+OXbASAhPwcB
ZHnwKrUQ8e67rJi/Of8YYDTIHAN44YV/FPAypfuxkSdgIApSSh7vMGTqB+WyAroA
3Ktb9GN4JuyX5vzcJ4lZsSQVCarksZoW8p5NSahRSzjIggJ4DGbt6I6ae5Og83Xh
fkLL1ulght4cDpRbgpsJpYOfBQm9KLuetHZkXGUt+zM5k1kk9K2qvvvh/VlU2g6i
o0qXVeF9JIP9zuzBsGI7Ca0syFwbyGRg6UXY7qZ8ay96DlF3KNvxQ/8FJtvIl2N8
Z63+0LRZ+OazT1aLpJF9b6hNvwafBs6GsXoHcRr726PQRsEsrghCgYdl//aLqXND
MiAuuCpw92PhVycgXylYXzedf9sytlO5wSMrIrCnX88QV4hZT9ERGg4jl+OXFDHb
xHI5qssuuZ1aZBRVwGhPczwH4fVXu2+RwmORsBaZN5Fhl3EpEpB1Yj8teDZFHj7Q
PEfmAfQpRwfErRSLTgZUJ6c1/+jJUEOzSbjBsMtP8MRz7JAFZHzuJQhAv+nnwcic
+UMDYFyHNL8MbenP6egRrUSdDfHgDFlesgXNQa2GdHr3rTmbhuRQX/o7SO/eOYCD
ecuhLSt1pTut/DkhC2GTE55O0f0OqgydFSB0RMZLRYFOyJ8uNe/Gu4XQwuzWQ5YJ
kxldLaOtVnCHEyhMkYAX4NOQuStVdFV00GjD75vEDrSA5EnNkewowtgZQyPo76pO
29K/+HFSa6O89/E4s3OIobiW7tCbET51xUt8YVji6300m3/3QljoAiSZg6xxmieG
cw4fH4vW+BzphrUzbUsOu5f0G5LPhBrYJy0ct89LPQAZGM769EZgEs3nvS5LvEOw
ObfXdH5CX6z0fhNYZBDB5hm+zANmUNJ7jZTT4pqncngi7hEirDTnwcO48Ezv8iL3
Q8ARPmFp1V1jmV1fBVd/RB8wM+Ar2j2GTzh/vkGS3sJOBEPe0asDUEqKyzN79/V2
jA48Kci6uUbtBuX8ekQQdggf1epNpjGuQFLEeO8GfE6rtSf1K1YTqy7cM902/XAI
8Yp5r+Xo4ToTRGFWjXp+xtl0C+QUeQ9kyRbgv0BwvZ57NvKnPWtN13lv2Ysq0Nlm
zAb+R0Hjm8sZORKiS5Vp2XhPIuOWXoR9leuzI7TcaJ3XyClxgRvmL7duY+ROIFzt
1GNnEkbHABexXxBNJb+uptmGFelhYPs2iMNfNVcX23IEOCwNnQKbfwvzms1SWDF8
7c7F5Tv2jiMTOR5daZeQKijlFgKLBfCQq+cCTCLmrP0o21lFv8NRIZvuKelelzEa
EYRk8LHwowxE5Bjkhb3DgKgKdko/JuJAWDGtletCq28zV+bqSAplUTRGyWS4NR7P
x3URWvK5gJVgXkADMNGbEsToCTvI/lswVkT/yzbzScTFmD8I1/OlMJSDNTYc/FnT
QUtKSz0r+y93gas+0FxUhJuN6jRmFb0EdBzVi2weSVj1/taXHj+ZHOnNmN21SGs2
GLbTqrXQOpODW7h/mOTunPCCik+LtKwRLZoshrePRygy/F83deCLJByxbbEzizk+
lAk8bytNnx+nE+T3bzxREt8Le2xCit1MPPhzcv75xFyPwTbywVI8pYOdZI7qsRSc
XoJTozf/c9PDhFm3Xjf+XuaPoFzZytl68+t291Mumeaa6XHojGBE225TI5Sqnycc
vZtxk9Ant1gPhRETQSuIIbhsaazdRUq80nI0AoFrA3Wq8zL/DCKE8jAooCz1ZbPU
HpZhm7wSlnmUU92sdLnd4YHEYEq2nzVsfFzMw2ZxKOukqNmKgWXJAhsbwhyo+dfH
saSAdKVSJUVBuENuTWLm+ZOt9p7kR+e1Ze6lgqWOCOOiYuoLGOciXjM/piYmp1m/
IQlh0BsYn0IK33Bo87NUcWvJEtX5I25czKnaY0GbHoXocxrGVycELaQO9fi61Pac
o3GzL7DnKLjL4IKBC2bSh0gBZs+Llfbn7BBRvoKKWeoKNVUSBIztt7VTyRHEPX2Y
+wOgq2MV6Y7x4wH4PsVRGXYTh1m1HhpZDbW3GBR4p4ZybYIfnjuocMXEGjlWbXRB
IJnXEiYF+UET0xkvMOy1Xb8QtO9DUoqFhWumnezbcGfghsUYhj94g7UYkuQdQpLs
qTl5yH7whLP+LnGU8kXt2y/HCyzb6n4IcgBAG1N2oITB3c16gbX//JtWb4sTL+nj
NOsv3Y9XYBJ0uEl8uX76r1YwuVxpEwPubTZtOz7WPxFQ8AC1oUh133MseCmVt4KO
QLTddgeiMhirgOocGPwWtheRbAnmVQ9wrD6mgMkcQNkDASy4o1Y+IHEahc8FoOPs
RA45+c5t9dOgAAVTFH9l/dms9w9ml9KABwZWsm6uBMNLc2tY/FtOFuPPXre4H2Nv
SsPlxZlIP0swYIMq0fWSTB5xbM5Lx7wdujan90FkpzBXlke9/yIZM0MNMsatQtad
/hbXGpHA3SDzZpE5DySZZlQa/JYVMzPJL8yrK9jKLPa+yT7NwdQnSxrIHfzcClX2
+JIDm2sAT+1JqaMSShwV5CHRcGMQD3bF4UbE22tuE/U/rgfj+9+z26fy5++pAJlF
dqRUAuMBGv7HK7XqWVs/EiVTYny/l0zh2owZ3BAO7U2bsfeCexx99x05Praj7PEW
YP5oJNW50gBBQm6hVBBkzbdbdCqqh0PBpa6PzhdhuwmRuUzEMkNj4QSYfRfYxU+u
91y/a1LaoVYV9+RxAEiXviP5R1ORaqB4AR7KyHineIi6qLzpj0l7q1aZKQHCc3tn
WMVi4tV2oU9TvtrJKilcsossqYwXktN+eHXe0qmOnk2JrSEWowmBRfHnjGYzP2Sc
9T1K7pXSerPzgvE/pWk+CeLR+iGXaarHZY4wIDXoFBNaVTKoI6dBnpghcAMtJHxw
1dxHEswsH+FzEOQPSphWKgxnfrJ3J/fx2WpHzsdelJXvwxTfZlGfsViNTE5M5jb+
2eULo5PycXsqGIu8dk7J92lJHnE4C0uLpuKW/Pn39gvhvfdO0/PQs/X0ROcS8lB6
btDUJ6m/hOBb0KeDZx4z4InPyClPMncCGwmMAniVf7HwpDHjUE3upo+Ek4IR/cP7
JZWvm8HJw7TlkX71wogCnM8B1KMwHPtDvT/QtNMMwPOnUfo+iZop2s747030KMRg
O/63d5YU/wo+7WkOERMRACZnB+jn9LHwOaH9Lm7mj8zBIgPBZwWZLKMUzYTY4jZQ
0pgIl+NDX6Sg26QzLt7yfkIxopPL/jOkRnNU1UR1DE08UygihR3DNSyLKsuz+Ye4
Q1e6oGu2yrBdhOSy1AkY6uRdMY/5qCObAerysnNw0x6003epUnBsJ9RINIJEBJn9
gbhq6Krb0GjSATgvK8stpCGgbJ1syHbs3pA5NjSVDJFSvRgbsum1rg9Ls2wYoY4W
54cLeMEndoLOcSY5/Bws4oAWaWAOeh2c0tjeSmPzCYTjkwbx1xZ1LBVedU1KBZUa
jhpswXSuOypljKxKTik/A8vUTJDNwquxQsYwwmPKqPlSW1LevaIqwOLPLmyPRKrx
JJ78fuNIHx9pVj7nMax1UDmWbOjQqdAQFeHwrhD3exIUaPPPAQGf8t7du0qpDmAA
Ixbbd9/nLLvMcYIs4700jY3EGFS0JYkWWUG4Uq+uN2p+2+IxgUF1QWm3HBYd8/c9
0uX/23EUiEAmasOrhpUHXfVuLBrukIVBd8H5i4haa5w6O/ouwjUQpor55F3PHNRZ
8Ih72QH7CMd+SXjtxKMjD9fRDajUdFTJ28VE+SPguEbIMU1P3j35CrGIcErPLEBP
GfyOiwGz4uyRfpLiqpSxdjx2qUf+qs6Snkq2AkpG2UiXICMEV9oJqfL20bcGqtmC
IiKeAIoJZKhVQRtSObRH0zLCBQdQXsbU2uynSYii0G1EymR+43GKFrLTO5FtNA7M
WVKPlXeuPCWhp64pFTjZiRMQMArwzrNd88EXPuUx8iOjZG8ZsmAVgk3XaG1gT6ZI
sNrHA4lcUenyJPUxEaaWAgwiyxgKEXWKvqOJ8c9T1H2jVAEiSNT6Rinx0pJKg3XV
Y4apysK2qJmmyofL60sbBSs3xrLPqfv41Q10Jt5Ps6o/3YUIp3N8hA1XKO7kSg15
KM2K77s/1nXteVjxuqvSmIQmwGRaMpdBe0eiA/LxfWo6bgdRpqB5Anu6qZM0tbg0
zxGdchCzJSeSNQ2mWSdFWC0ijMP915a50v6/HHUzsqccweBmynVrL6RYjIVZH108
lBCE0/VmqbRn0vTsQdvOKZTQ3GPO6ULxaEn/iPbzmRJkzpbW6jKZrypc+0bxo1nc
KV8MEMpJ8llDov4rVT9VP/5EpZEU8OCJUBrkqaWmEV+YnvfCelTRdbgQp1FLCW/b
cHPD7Ykov+pxiRpBgzVfSydCt9OtSfn1gyclsUDXy/hCI1wT+svqdtC9CjK0QtlY
usnF298M+wDkJsm5Bdz5qitslXyxCVDjg7nng1DaYuGWDez1yLWZx3DHjM+b1/9m
gYXMoK1ejLTRC7TilJzPRtPfE5ltgOmwVbdlK5r3iQueSirEi6VS7Wmc6nK7+Fv0
B2I71KFnTNexFB9fjqwu7j8L/ndF9xbAxOMyJlxnm7Q=
`pragma protect end_protected

`endif










`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
e1gvKs4lrBejvhuSk2pqsC7it51jGlkA1tyr6wzAWrFJa60oYOTSJfGzyi21P5rr
0lJK1GAyrRvZjVNjtkl2IpTP9dBrFopMXvwwDeUHLjC5qP+NZFz5tCi0NCK1NkED
m28Pg7OTrnK1Nd5ECCNNdxpzNLNBTCS37llv+eUvuZ8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 113212    )
EfhEZa72TFEaraenJ/0GnOQdVsSVojodlIH0vwYCLmxbG0oylyknuX3p9cXlyjxE
+cjylVZ3Ci0bdGWFvVdpSAa8VRuNRNF4+mCER0xXVE9jSA0dY1o8q+XJNMGsbRU5
`pragma protect end_protected
