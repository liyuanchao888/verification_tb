`ifndef ADDRESS_WIDTH
    `define ADDRESS_WIDTH 32
`endif
`ifndef DATA_WIDTH
    `define DATA_WIDTH 32
`endif
`ifndef NO_OF_SLAVES
    `define NO_OF_SLAVES 8
`endif
int number_of_transactions = 100;

