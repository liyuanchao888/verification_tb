
`ifndef GUARD_SVT_AHB_CHECKER_SV
`define GUARD_SVT_AHB_CHECKER_SV

/**
 * Class declaration of each of the error check stats instances using the 
 * `SVT_ERR_CHECK_STATS_COV_EXTENDED_CLASS_DECL(stats_name) MACRO.
 * 
 * Each call of the MACRO would declare an extended "svt_err_check_stats_cov.sv" class
 * named as "svt_err_check_stats_cov_<stats_name>".
 */
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
KJmxfuJA7tfo73uO6TC1e8l5b/RBnwnIhCH3SkR7VUsyGGSBjhqaRIvmjcD3w7qO
bByW7r4p1aOlVKxT2Yy27+LXC5nDG4jYpKgjmPibQiA+MzcMVldFyTuDK849k6cR
KruC+iuGSd/P0nxZemN4iJcNXcMIA6X43EIYvJIRpd8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 5847      )
6Y+4kuZ+lvYzA9Ah6trtyDAbypW5V7Z/5AhMIhsMJy/pebdXoYTEd+m/kgG4nsSs
OrKY4NcMgai5CYoGVPzPA1751nuLgD9z/1VozdQhZZC+0CP/EZhitqwmh7VOlCBJ
9m+Vxpiwa9NVDhAeMYFYNDhHqhUJu/yGcz9zPCXhR5WsdGOxoEmC1cx8V03H8B3s
Kbvazo6H4H/573I1WJ10852LHHkUdD+sSaX6Y1b1L2b8rBLWs3qd31XWRKReR6Ek
uChLqKGB7/dsVec3PZqaqSpXDgVnE6mlYDXoaed4WKYAiL4GThOGzDa0RWyp/nfD
NpSHgEEGJl7SiE9nBmDKjq0nIG+xwRG0mt/NtdiHtR4M11BAqoo8O+XcoRyfEngC
3cDyeWK2cYCxTHSLCMsc5Mb2BPmbpgnLImOHwFP8AUKIudMR3undhK22g6aS5Q0U
pPRoX3ct0BfsQKfcOIaOIZBybEtQnInt/aQb+2SNoKV66e9lIyscPK9kzpXALkn4
YsLChkz1Cq2ZPk/LXUEk/WE12oNcIyPUOPtpefpr8Ci5As7lZOVT0SfY3UDHdbnF
kiim/3SRdQ8TVRYjKIl93F5DR6rYzjdqKPW4VXvikwuZ1X1rvGWpvs5RHeFw0re/
UKCy0Fj1d6DLYS4VFxrLAf/DueG/DRyMmrIQNLk2VUSRjKO6yu8R13eMrR1t8zG4
EOFWS93XTFDvKJmIUbeLBw4hssvf6em2Q2HFCPtv4BzMVcx5zzv2hRpGVt50Zbqz
tGPT+3qKoFHHNO5hjCJGvNkpefu59SA4YMkgO0CST/5sxzTGA8eG4uTf4I+tRjT2
XjacPLTyBoZRLDjJIf6Sq6AWlM2PjyKYtUG5Ep17JhhKy36vl8eJ+15A62k5wdTD
kob8uxwZrDY0snfM/wA2HZSuCFALC00ndV3XezqfCnuzaZqka5IMsqHNOofK3OLB
9nxrsKSSIYUAgwH+ldjJpopmfeO12e47aBTlVCV85F7CC1fNMitHHK6QHa/YAfW5
AB7r8r33ReIhKqN5qbPpmc4bnhk0wJHebynuZ3mh0viLywCXdov4U5H3eA0Mqv2O
kjrApbPMaWw/ipafDgwx6f0ua0cGAv8mAHNlr+VQLX3NiCIjeKdreKA53lGV+FqU
i8nS/Kl5GG7I8NLzZK+VRZyHPT41ClBNjrb2nUejL/+HvovJRtZ43RmBrKxxBFAF
n5MVEF1jw0AoQ/honfSzaVDji3DKzrbb1CgNeF8HWuEcbLJqR3J42YVBMtNEMTdy
f5k9KfZPxHE2/YQtAqjfOGeMAUcto/4knPB/4pEtYBklVE9cdY3UQxKjJY1UACDk
gw2Jb+yVF0zuEfVKWU47fG1kYGwCS0qjF3G58Dvy+or0FejXxcWN9KAGwsCFCVF+
FF/Z5EqtwlsfBXREjiHihJlKD/XdpnFjlkUKrO+D1Ha8dd4LmuxmsZ1pJVlgwRpJ
cGW2VW5F+zgxSqNdYiQiD2w3GdG/lI4v0qr0M6NKjhpwF1y1Epm4V9cEYD9C0acb
2Uf2NFBVPm8Dy36bYP8+OEOsVDmQWYg0K+iOMN6MSfMimwBwDgqqr8jy+ediJ0XL
xeNHsXsOVrHgI+yCaKyBhEBjiAVFCMPofGRD0fZcCXupCq9lmzY4eIGCO3iTPluM
zzPg+vHmlfOzdHErGuR9OEYI3L5IZFNB7x1k0LqBoQKeeE7NmhSxwE6X1NDxYUAe
UNkhbGxRr8SpSL6EsNFgoJntE88aPWls8C7Ik+Uu7JMzVj7WRZ5jQj9caydCRpR1
zSPt/dQd9qZ0dMhHkWjWfPyZEYmxrOjXoaDtIOw7EBJVngCuu9Nk7NDBS0EjlBK3
gh4SwnsoFl6GoHVL+SrkGqr03oRNHyt6a7UU9PWGf1XPSLxAtNe+VsXWHhCMH3tC
Muca8s7kYQks/0GhBgVaHJOwFVc5iTiPNe6o5oH0oZiZEfSOvJ3vqhKCpLi8vGDQ
gVkJuixf3vLzy6OBpsR7Yg82p1B67S4prWN4QMyMTVnpIRrZBjY5Xlqds53TaYZs
VDncjgVphRah0/hybIk4RK1g1aE1xtRhhnSDl/qVym5ZAw/Wu0axXiuo0j8HAHFy
Q4D1p4KrESr3C02btpUzRZkZnsWb0ehTtHfLaYdTHlC9qsdbLXiQyRp7GXYnwp+U
oohtdRTOzEq/8OTJxWPweDgD+EWiSUfy5j+ejJk6EE0TJATPNBQJG2UUda5g5wPv
pAWXPVWAUn3ibde5YcMQPXRnidVo2Wx9hORXnHL8aZFLGj/sLPd8q6FX2hZhFwxe
dWpDbTVcks9mole42zzMXpiMC1a65CUY7vYaoqtw1Mw5isyZLsWApuAJk+/s2vpZ
36eVkRo9Bowga55JvWyQRugkIX7oRXmUY5x9qA/ZeV71Xi04Z87Z/t6H3Z0XSLoh
ajDFvPzu2DpNnGQ+r3epfJnbqWS1A2El1Cg10OK7su7gw8xCFNef3LGyHtLJemZe
wET7sCIYx9RPTO8dRqt2xSxLitEgY3fCx2KQzBaR/+s2aFgvSF4Ij9Z+KmoFg/Fb
VC/iEdY14heifmGzi8dqu0Hma3lmuy4o0b0oQyXf5SsU3FzBfc2KFg7Yxf/9gdwt
AJ0gdMh/9knXg+QwBW9PYuXgQfCJDc7W9Aj/YnCX10H+6E4T31x3xE15iYWhoZ9b
ictQ+IBQi156y5o31890pUMcWiBB0duoxlDHvVGEzWeNxczwIofjcqZWZrrsXLgQ
Zcji4E1Pt8DiZSWkms92d+BvnBDBTcCmyDnQESrB9541B1hjszBGMrMNkxIctBa6
AT/6Xr7glMjgGpf4ZeEb8b2z8VV888pK/Cj/xtzroEWCUH7adtogg72SShKRVIvH
BZrzEVHVq0VE14ktcVKUf6mylKMfnlEzY9gwNDish5a5NmqDWKjxvXi1g0J3TUNN
QtamZYrRJD3D/A088Wd5MXUTJDE2AlokuQeQty66HodRicnu/kcrz4oy1loO2OFk
unws8zXeSBazpd8esLqjuaWO8qsoSXI5PKje9EpQyi08MIWQyoq/IOcCVno9aR4w
RnIvBoVm1VAu3FmKFb3GuAxv1qFxAXRGcwIeP3VPS4Q+waW3t0HrdPIqNEhxWP60
7IHcfaD3AhHPx1cFY/ZUvFtUIRHr4ScO7/5pDlqLjwmOqjvJlNDa9Y8LuAx01wBl
OSTS6O+laUPDv0wtVSOsGj61Rv1jpNlEKc0cXlXEQ8jSPoWduH9sWc8Ty8lGQyYv
x/YkkKuJlW2WoWbZu5qKdygBQlxM4WuQSLEQomRkvbVPlKcm+RWc5ZrNBPuBoyMf
A7ZJTjBDpK0nezJkwTiQmc2DPGxtHJY7dvFDSzOYyz0+Rbmk3Dts1L6pkS1evwW8
LM7DtZ19A8tEmB/hwnaKMMTlEeTMIH2qVoMXXP0UCJTPz33Gq3FPSfQluD1xg2AC
gXDGoFAp9ovalP4RBL7p6xHobgZbrtDcwuD7NiwNP6BPyC3Julv5bwxiQIcxybFV
UW2RDrRlAWNzJfy6I2Q980mY32xTRsJmKHbVkffUeq7Qdifrf2gvUYFP0g2jhK4H
jv57Bd5zrpnk1QnS6oy0o8hQu46oLeDVDrACiSQohM/gU+wevFVmlMWTf9Bgs9pS
O2dVP67192FuLxzwlUbG2Xk6gVelEMfvxvofzY4WdFbtyQwpbwLbAV2lxnJ2hnFe
68OrdL5CKhUCdZ4SWBIP1qDcZekW383x2WuJ3JgIxZFAnB5nN6KNGoXE1zL/SUbR
AxA2HqOWaYiv55BqCEPSyLD/HABm27gyTK3+f5aN+zZQ0aRvwv6AQlftssF2p5XD
eGIhatsCtf6iShI99M0XrhAWnEMBcLmDj7ZNQ/OGM21UW9+dC8XwGllTriQUH8J/
M2ORsgqPxdDDiqro8911lMA2/AOyKMQWI3ZEI+OVhVrcJbUJPQFDBUTs+WpWyg/p
gUkWo2y/+I5dMXiqeSbEUU1wezrYWvPulz7jQOJqJoGMvOCGXOKoyGToPZJ2cfO/
MY+74rbTnOWS8jGmaG7GnNcXPIEJa3IwvMQmhyKDbbcJZyhgy3rovm3DH7ZCm+CR
cET7ocGVzaGBDTgRDhv20ya/iFc3AiCKI4p0WOJAhr9NiBoeQcSyhMnZXU4VV0aw
cjeCYaVfL7gt4FU94YTcfr98/EOFsNoxh95w7ncppFHSmkNsxQle10fi5QOxMCtc
CUTEhLvYABTI0ErF6Yjr4Hor2ANTG0J639Lm20w9QS7GkdNDVfMFsVTZHYju2V1b
Kdm9jdLYaA+f8JFhP/bXZmGMGvFY6EZ0X2iiHG50wj3nrbdADoY8qKNfAUGEzL89
uaDPob6F9UodhW3Gd75KwHXbUxDWmG+JRITKp2/XSY1anK18VLdBJOdKU5mIrRt8
Wdo/dAJrB3VWOHF684E/EqDSd0d4qaVKCEcSi5L30LmdIZhrHvHd63wUIVb3Ukwg
mjwLs8S0Eq+3A4bL12ooR2Wa49tWr+Fv4kR+6HVkYpE75/coPs62YYmMxss9qbkR
tdl+2K0samhcfKMJ1BXxDvtsh/MtvVRg3NznACcewb7vbhsIdBVm8xowzvyEP36N
BHUTksS7FTdECouLq85kA7B9sZrPqkqNJcmp1jNFnpHm0o+pjtIxuEBOt9vsUGrW
qH31tuaDqWKP7bm1+magJsUTSFt1NRroM+p2MX0JS3ELIoSHmTxEO/dPScf2C8sF
PFD9lRfwvY8wPUDudNRtF2S9aAZJmRhS7o+/cgEetjZsxxmF1F4jAZ3/sAlJ/kpF
sofZJHHggCoavr3If6GudNw9Hl8gRa8Vba4SSPyk4FyU4HjMH1g9BxHlUxLt/k+Q
51DGrwG32eZUZUj9Yp9tywi+zgQAKX77+R9U2VXvXA4rBc2XINm7YrAyIF1fo9Y5
LhaclGc5bE0EFC1iPkEr/+m7M1XGanmo7rkD8jiftYcr/e0XM8fhH3CHIFGmsQxJ
gXMD19JcfZVEltuAUDn7LdgXB7Uchbhjuuj8V8dAKuf2+KBcwnw8ixEdwBq70KMc
Jh6cT/h60kJo++cPKYvrW/9TOVr0MJKpQZ2uebtXgkggf5bp7njiT0qCwQpGtL59
vY27kgBwQhaRYDKs4yaLbwjrUp/3oN9ggluWz8FkQO5w7PkYrTmUOE16zyl4YKtb
ihhDITAsRI8LS5ORPSTT8MLA+7TaNPqwwKna7AzJ5OIHLT3WZTFh6DaQ2dEy6fI4
Jx5lxAdpZijVqe3waeFBYiw0UQS9RTHNDV5nbGlYWllKLhH9xdpKDZVEgEM7x4sM
k9sPihDNGNbsPLd3Pv/8dwaBtDd7DJfWzygWIZtlCvm1b7bcDOTB4eZXosIiqqsx
Tn+hjwKqzi+8dAPQhtam1RyRpNHqlvtnsi/LQ9UD8uvddeJipKnfesOflbZT6h8M
IU9CKWLaJh+lgwVWIrbMGlDnKyEfBdc7PNCMI/zeifNFWQJ5SUo2sx5KNfIYoutz
L2odFiO//iXbFvCFdD9HHU9pTnP+Abcuz0Qwu69IIZSbL2PvLOOJEvIMVXYXNDCR
MLlliwFE08GjGeul/5gJxGxIPv0jo36oRDNj34TciJp98f53lg9UgZXEJEktze0R
jOuwTdhR4vWyre5uIg+8VOKnGcLopiTfrjMQmvkpaeMXfO1SsdPfa+zxGEUv8QP7
aKv6Iqx4H/bXPOGcTLjEUpKMkx2jjQ3PjmSz0SJbHO8sBuHritSzjUNh10ETyllt
Y6ZZxArSGgLm5Y6Kl7IsNE2UuUG9Wluf83WVcz9SmRM9ZaXbjNEE7hlI98Dq1Go8
vU5LfvMiSuShlvKugAHImocy/mL+4gP8wvQ7sI6ZNB+5gcPWEb3EgDbZbZinpPyA
D2VPuJnDQpJSamaqrSb5d3IEYbUXJLXCmB8wcLSPFJ7xZcvjTNvn0vajv4ZYImQn
Okbrb90XCTHkZPldVzxqb8AFw1Fw/6+pKt+hFNWK7s2lOylE+O9OZfG/JAKkQ2gs
qCN9j94iQz5tRBC4angQUepYEbP3SqyRVxcHoHjXEGa9FLKkUBNT3sIE3SdGKVAY
wuRDYOb/xfEeu2098ZELx3VOmJhwoN+TJ7rK12WzKx5wopgCnGGL2AIMAclIoI3w
+6zV2p8ykHVPUPY41Zoxm+kF/tyd7SmdDdD1uklFU70QvIf3CRUltNffzgEoCNyW
JbnjuoX6x3ZcnnOWUjRQSe3lKTsP5MrZ9Ma0rjP5Yg3XblySPu8/n8OVnYJuy2XA
6n8cmrl8FG289uWxnloxK7SWtbvsn+xHmcJ6qMkcrtloSWio3hrieLGX8nVLqrjw
Z/msUXluVkTzFA5WIIMdPM8i8DEgh47HBbzQu9V3sDz2vUiMRnaqaU9DhD5fhnea
M+NJ1vAVmWCMORfwdsc/kjDPS1c4OmHMmW/islJnARlROesGw1yWe5QXPbMwKjVW
Dizvka9sTzXKeHb9EMGfUYidC5/EIIjZVYlgp4dylM7gURupfM1TMRQdPAPa7olF
0/VnkawGDEnqD2O7RfSg2f8SE4+7+Nab7NqZmYIFg/A0nCtUtM1t1Akq8ZrAWrGT
fHjhmVe3+psBw2qegpGPe/3khpjGhAWooKqhoMTuozLaY8cCtqHG2AKHZPDGzjKN
4cuymrABQSl4FImtAaNz8B4WRH4KpRFPIRbnpzLGyWXoMafmZQiKbXta0TVO/uT+
7Rw+XwvVq1TdJn/g0os2pD7oF28XWI3q4mRTHPX3MBfj+o9e++alfNbY2QdpK1N4
1ZI3V9y59pGvZbEdoFhrxkwnXC9ZkhMxnmArycAeYYWkZZHvz7Dk7Ivzqz2I1WwC
ycxkl52xJXyuFR0bDocWTqqvNs834nsXKQ26PvPMcFJqnUHfzVX/Nm5iZNBFZEZP
VIaG81mEBlazMUB28PjRSvu2bSRpkwMyC5RMYVRYNopEXQF7xL5WdmGrb7xsxtrN
3CSaKJXOVh1lZqk8y+6JqY8w70J4iAlBsR9xN/zYTeRc8h+pshXdFo9NSpiuhFmx
U83AU7oPcGr+ey9NJXGDw8Gcmn9RDrwaRaqf74boHdYABYOu5HnIa3/PvLI6pFFa
Jr4rufPQbMhMpeUjkryxUPocgMZRVO9rptwrQDShx6VhgguOURYQ4xY2lDFoQ/1e
pCqzO+ST78sy/bLzBfds2Hsy643CV/tMjwgNd6A+WIgPYg/ttMsiMxb2AuiEeR7u
9jASpio5Gcy23NSQJj9dzamkOPvTb5O+8JPB4tBCrkOHe1tGX3yhXLtmMP2uI+g5
rkpG6VCRbiETLHU5SQP3dvEghPSQXDQIFci31tXiRWCqPaBay8T2M8SWx5YSymdT
R2SUL4ZDZR86HG2JYjCw95/6HzdjjBLAHLqC4H/u9d0CSs5FqwqqK6tNtA6wBuGw
JodP+/eCEQFJpiRJnOPVdvnFwTX+nYAKH8MnfRb1CBTLFjDwQU+5Qp4crITHiOiL
C9bdjEWtY9ww0+LH02QdsS+Ook7x8QPU4amVSlAA3wpO/aVC3aOgduG8RkMlKUuV
2HX0G+M2Oh/mrZMZZlDThQFkNNq8RvdIWT75ftBXV8yA5nsO2U41nMaNm82V8hsO
gdNfH+CapQ8ot4c9HaX4nf2E6A64u5eoF+Wvaw4n9Y27BJWulFMtBZ0qofUPUDXW
zZUkoNk/ZUi7IW2kHNm2Bq8Qo1kjqGcEhcMEHIN9E0qa5uuh6JQgk+B57METtJRB
uW5iKz0XHRiGRYFztzvt+6YhtnFQhwoeejue2LntL3bO44WFTU6w0ME8ED8wlGtV
`pragma protect end_protected

  class svt_ahb_checker extends svt_err_check;

  // ****************************************************************************
  // Public Data
  // ****************************************************************************

  // Signal level Checks
  //--------------------------------------------------------------
  /** 
   * Checks that HSEL is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   */
  svt_err_check_stats signal_valid_hsel_check;

  /**  
   * Checks that HADDR is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.  
   */
  svt_err_check_stats signal_valid_haddr_check;

  /**  
   * Checks that HWRITE is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   */
  svt_err_check_stats signal_valid_hwrite_check;

  /**  
   * Checks that HBSTRB is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   * Applicable for AHB_V6 extention AHB_LITE
   */
  svt_err_check_stats signal_valid_hbstrb_check;

  /**  
   * Checks that HUNALIGN is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   * Applicable for AHB_V6 extention AHB_LITE
   */
  svt_err_check_stats signal_valid_hunalign_check;
  /**  
   * Checks that HTRANS is not X or Z  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   */
  svt_err_check_stats signal_valid_htrans_check;
 
  /**  
   * Checks that HSIZE is not X or Z  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.  
   */
  svt_err_check_stats signal_valid_hsize_check;
 
  /**  
   * Checks that HBURST is not X or Z   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   */
  svt_err_check_stats signal_valid_hburst_check;
 
  /**  
   * Checks that HBUSREQ is not X or Z  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hbusreq_check;
 
 /** Checks that HWDATA is not X or Z   */
  svt_err_check_stats signal_valid_hwdata_check;

  /** Checks that HRDATA is not X or Z   */
  svt_err_check_stats signal_valid_hrdata_check;

  /**  
   * Checks that HREADY is not X or Z   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hready_check;
  
  /**  
   * Checks that HREADY_IN is not X or Z  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hready_in_check;
  
  /** Checks that HRESP is not X or Z   */
  svt_err_check_stats signal_valid_hresp_check;
 
  /**  
   * Checks that HMASTER is not X or Z. This is performed in full-AHB mode.  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hmaster_check;
 
  /**  
   * Checks that HMASTLOCK is not X or Z on slave interface. <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hmastlock_check;
 
  /**  
   * Checks that HPROT is not X or Z   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hprot_check;

  /**  
   * Checks that Extended_Memory_Type supporting HPROT[6:2] is having valid
   * values   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hprot_ex_range_check;

  /**  
   * Checks that HNONSEC is not X or Z   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hnonsec_check;

  /**  
   * Checks that HLOCK is not X or Z on master interface.  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hlock_check;
  
  /**  
   * Checks that HGRANT is not X or Z    <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hgrant_check;

  /**  
   * Checks that HREADY output signal from bus is HIGH when reset is active. <br>
   *  This is applicable for:
   *  - Master in Active and Passive modes
   *  - Slave in active and Passive modes
   *  .
   *  This check is performed when svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1.
   */
  svt_err_check_stats hready_out_from_bus_high_during_reset;
    
  /**  
   * Checks that HREADY output signal from slave is either HIGH or LOW when reset is active. <br>
   *  This is applicable for:
   *  - Slave in Passive mode
   *  .
   *  This check is performed when svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1.
   */
  svt_err_check_stats hready_out_from_slave_not_X_or_Z_during_reset;

  /**  
   * Checks that HTRANS output signal from master/bus is IDLE when reset is active. <br>
   *  This is applicable for:
   *  - Master in Passive mode
   *  - Slave in Active and Passive modes
   *  .
   *  This check is performed when svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1.
   */
  svt_err_check_stats htrans_idle_during_reset;   

  /**  
   * Checks that HRDATA/HWDATA byte lanes are selected corresponding to
   * bits HBSTRB signal which have value 1 . <br>
   *  This is applicable for:
   *  - Master in Passive mode
   *  - Slave in Active and Passive modes
   *  .
   */
  svt_err_check_stats valid_byte_lane_for_hbstrb;

  /**  
   * Checks that HUNALIGN output signal from master dosenot changes its value
   * in middle of a transfer. <br>
   *  This is applicable for:
   *  - Master in Passive mode
   *  - Slave in Active and Passive modes
   *  .
   */
  svt_err_check_stats hunalign_changed_during_transfer; 

  // Slave Checks
  //--------------------------------------------------------------
  /** Checks that RETRY responses are not received when configured for AHB Lite */
  svt_err_check_stats ahb_lite_retry_response;

  /** Checks that SPLIT responses are not received when configured for AHB Lite */
  svt_err_check_stats ahb_lite_split_response;

  /** Checks that only OKAY responses are received during wait state */
  svt_err_check_stats non_okay_response_in_wait_state;

  /** Checks that ERROR response completes in two cycles */
  svt_err_check_stats two_cycle_error_resp;

  /** Checks that XFAIL response completes in two cycles */
  svt_err_check_stats two_cycle_xfail_resp;
  
  /**  
   * Checks that HTRANS changes to IDLE during second cycle of ERROR response. <br>
   *  This is applicable for:
   *  - Master in Passive mode
   *  - Slave in Active and Passive modes
   *  . 
   */
  svt_err_check_stats htrans_not_changed_to_idle_during_error;
  
  /** Checks that SPLIT response completes in two cycles */
  svt_err_check_stats two_cycle_split_resp;
  
  /** Checks that HTRANS changes to IDLE during second cycle of SPLIT 
   * response */
  svt_err_check_stats htrans_not_changed_to_idle_during_split;
  
  /** Checks that RETRY response completes in two cycles */
  svt_err_check_stats two_cycle_retry_resp;
  
  /** Checks that HTRANS changes to IDLE during second cycle of RETRY 
   * response */
  svt_err_check_stats htrans_not_changed_to_idle_during_retry;

  /** Checks that IDLE and BUSY transfers receive zero wait cycle OKAY response */
  svt_err_check_stats zero_wait_cycle_okay;
  
  /** Checks that if invalid HSEL is asserted for selected slave. This is applicable only in mutli_hsel_enable mode */
  svt_err_check_stats invalid_hsel_assert_check;

  /** 
   * Checks that HREADY output from slave must be either HIGH or LOW when there is no data phase
   * pending. That is, checks that the slave cannot request that the address phase
   * is extended.
   * This is applicable for:
   * - Slave in Passive mode
   * .
   * 
   */
  svt_err_check_stats hready_out_from_slave_not_X_or_Z_when_data_phase_not_pending;

  /**  
   * Checks that HSPLIT is asserted for only one clock cycle. <br>
   *  This is applicable for:
   *  - Slave in Passive mode
   *  . 
   */
  svt_err_check_stats hsplit_asserted_for_one_cycle;

  /**  
   * Checks that HSPLIT is asserted for a master that has not SPLIT earlier. <br>
   *  This is applicable for:
   *  - Slave in Passive mode
   *  . 
   */
  svt_err_check_stats hsplit_asserted_for_non_split_master;

  // Master checks
  //--------------------------------------------------------------
  /** Checks that transfer type of a SINGLE burst is NSEQ */
  svt_err_check_stats trans_during_single_is_nseq;

  /** Checks that a SEQ or BUSY trans only occur during active transaction */
  svt_err_check_stats seq_or_busy_during_active_xact;

  /** Checks that htrans does not change during wait state except when
   * htrans changes from 
   * - IDLE to NSEQ during wait state for all burst types
   * - BUSY to SEQ during wait state for all burst types
   * - BUSY to NSEQ during wait state for unspecified length burst
   * - BUSY to IDLE during wait state for unspecified length burst 
   * .
   */
  svt_err_check_stats htrans_changed_during_wait_state;

  /** Checks that contol and address does not change during wait state
   * except when htrans changes from IDLE to NSEQ */
  svt_err_check_stats ctrl_or_addr_changed_during_wait_state;

  /** Checks that write data does not change during waited writes */
  svt_err_check_stats hwdata_changed_during_wait_state;

  /** Checks that burst transaction was not terminated early: 
   *  - AHB master should never terminate a burst transfer when OKAY
   *    response is received.
   *  - In case of Full-AHB mode, the master should rebuild the burst
   *    transfer in case of EBT/SPLIT/RETRY before initiating new burst.
   *  .
   */
  svt_err_check_stats burst_terminated_early_after_okay;

  /** Checks that master attempted transfer size greater than data bus width. */
  svt_err_check_stats hsize_too_big_for_data_width;

  /** Checks that burst transfer does not cross 1 KB boundary */
  svt_err_check_stats one_k_boundry_check;

  /** Checks that burst transfer does not cross configured boundary limit */
  svt_err_check_stats boundry_crossing_check;

  /** Checks for illegal address transition during burst */
  svt_err_check_stats illegal_address_transition;

  /** Checks whether control signals (other than HTRANS) changed during burst */
  svt_err_check_stats illegal_control_transition;
  
  /** Checks whether control signals(other than HTRANS) or address changed during BUSY */
  svt_err_check_stats ctrl_or_addr_changed_during_busy;

  /** Checks for IDLE changed to SEQ during wait state */
  svt_err_check_stats idle_changed_to_seq_during_wait_state;
  
  /** Checks for IDLE changed to BUSY during wait state */
  svt_err_check_stats idle_changed_to_busy_during_wait_state;
  
  /** Checks for IDLE changed to BUSY */
  svt_err_check_stats illegal_idle2busy;
  
  /** Checks for IDLE changed to SEQ */
  svt_err_check_stats illegal_idle2seq;
  
  /** Checks number of beats in a fixed length burst */
  svt_err_check_stats burst_length_exceeded;
  
  /** Checks that a master started burst with SEQ or BUSY instead of NSEQ. */
  svt_err_check_stats seq_or_busy_before_nseq_during_xfer;

  /** 
   * Checks that for non existent memory location default slave should provide
   * ERROR response for NSEQ/SEQ transfers. 
   * This is applicable for:
   * - Master in Active and Passive mode
   * .
   */
  svt_err_check_stats illegal_default_slave_resp_to_nseq_seq;  

  /** 
   * Checks that master loses the bus once it gets the split response
   * from the slave. 
   * This is applicable for:
   * - Master in Active and Passive mode
   * .
   */  
  svt_err_check_stats illegal_hgrant_on_split_resp;  

  /** 
   * Checks that master asserted hlock in the middle of a
   * non-locked transaction. 
   * This is applicable for:
   * - Master in Passive mode
   * .
   */  
  svt_err_check_stats hlock_asserted_during_non_locked_xact;

  /** 
   * Checks that master drives HTRANS to IDLE or NSEQ when it
   * does not have access to the bus. 
   * This is applicable for:
   * - Master in Passive mode
   * .
   */  
  svt_err_check_stats htrans_not_idle_or_nseq_during_no_grant;

  //-------------------------------------------------------------
  // START OF PERFORMANCE CHECKS
  /**
    * Checks that the latency of a write transaction is not greater than the
    * configured max value
    */
  svt_err_check_stats perf_max_write_xact_latency;
  
  /**
    * Checks that the latency of a write transaction is not lesser than the
    * configured min value
    */
  svt_err_check_stats perf_min_write_xact_latency;
  
  /**
    * Checks that the average latency of write transactions in a given interval
    * is not more than the configured max value
    */
  svt_err_check_stats perf_avg_max_write_xact_latency;
  
  /**
    * Checks that the average latency of write transactions in a given interval
    * is not less than the configured min value
    */
  svt_err_check_stats perf_avg_min_write_xact_latency;
  
  /**
    * Checks that the latency of a read transaction is not greater than the
    * configured max value
    */
  svt_err_check_stats perf_max_read_xact_latency;
  
  /**
    * Checks that the latency of a read transaction is not lesser than the
    * configured min value
    */
  svt_err_check_stats perf_min_read_xact_latency;
  
  /**
    * Checks that the average latency of read transactions in a given interval
    * is not more than the configured max value
    */
  svt_err_check_stats perf_avg_max_read_xact_latency;
  
  /**
    * Checks that the average latency of read transactions in a given interval
    * is not less than the configured min value
    */
  svt_err_check_stats perf_avg_min_read_xact_latency;
  
  /**
    * Checks that the throughput of read transactions in a given interval is
    * not more that the configured max value
    */
  svt_err_check_stats perf_max_read_throughput;
  
  /**
    * Checks that the throughput of read transactions in a given interval is
    * not less that the configured min value
    */
  svt_err_check_stats perf_min_read_throughput;

  /**
  * Checks that the throughput of write transactions in a given interval is
  * not more that the configured max value
  */
  svt_err_check_stats perf_max_write_throughput;


  
  /**
    * Checks that the throughput of write transactions in a given interval is
    * not less that the configured min value
    */
  svt_err_check_stats perf_min_write_throughput;
  
  // END OF PERFORMANCE CHECKS
  //-------------------------------------------------------------

  
  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

/** @cond PRIVATE */
  /** Reference to the system configuration */
  local svt_ahb_system_configuration sys_cfg;
  
  /** Reference to the master configuration */
  local svt_ahb_master_configuration master_cfg;
  
  /** Reference to the slave configuration */
  local svt_ahb_slave_configuration slave_cfg;

  /** Identifies from agent cfg whether a master agent */
  local bit is_master = 0;
  
  /** Identifies from agent cfg whether a slave agent */
  local bit is_slave = 0;
  
  /** Instance name */
  local string inst_name;

  /** String used in macros */
  local string macro_str = "";
/** @endcond */

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param name Checker name
   * 
   * @param cfg Required argument used to set (copy data into) cfg
   * 
   * @param log VMM log instance used for messaging
   */
  extern function new (string name, svt_ahb_configuration cfg, vmm_log log = null);
`else
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param name Checker name
   * 
   * @param cfg Required argument used to set (copy data into) cfg
   * 
   * @param reporter Report object used for messaging
   */
  extern function new (string name, svt_ahb_configuration cfg, `SVT_XVM(report_object) reporter = null);
`endif

  /**
   * Execute signal level checks on the read path signals (driven by the slave)
   */
  extern function void perform_read_signal_level_checks(
    bit                                    checks_enabled,
    ref logic[`SVT_AHB_MAX_DATA_WIDTH-1:0] observed_hrdata,
    ref logic                              observed_hready,
    ref logic[(`SVT_AHB_HRESP_PORT_WIDTH-1):0]                         observed_hresp, 
    output bit is_hrdata_valid,
    output bit is_hready_valid,
    output bit is_hresp_valid
  );
     
  /**
   * Execute signal level checks on the write path signals (driven by the master)
   */
  extern function void perform_write_signal_level_checks(
    bit                                      checks_enabled,
    ref logic[`SVT_AHB_MAX_ADDR_WIDTH-1:0]   observed_haddr,
    `ifdef SVT_AHB_V6_ENABLE
    ref logic[`SVT_AHB_HBSTRB_PORT_WIDTH-1 :0] observed_hbstrb,
    ref logic                                observed_hunalign,
    `endif
    ref logic                                observed_hwrite,
    ref logic[1:0]                           observed_htrans,
    ref logic[2:0]                           observed_hsize,
    ref logic[2:0]                           observed_hburst,
    ref logic[`SVT_AHB_MAX_DATA_WIDTH-1:0]   observed_hwdata,
    ref logic[`SVT_AHB_HPROT_PORT_WIDTH-1:0] observed_hprot,
    ref logic                                observed_hnonsec,
    output bit is_haddr_valid,
    `ifdef SVT_AHB_V6_ENABLE
    output bit is_hbstrb_valid,
    output bit is_hunalign_valid,
    `endif
    output bit is_hwrite_valid,
    output bit is_htrans_valid,
    output bit is_hsize_valid,
    output bit is_hburst_valid,
    output bit is_hwdata_valid,
    output bit is_hprot_valid,
    output bit is_hprot_ex_range_valid,
    output bit is_hnonsec_valid
  );

  /**
   * Execute signal level checks on the write path signals (driven by the arbiter)
   */
  extern function void perform_slave_write_signal_level_checks(
    bit            checks_enabled,
    ref logic[(`SVT_AHB_MAX_HSEL_WIDTH-1):0]     observed_hsel,
    ref logic[(`SVT_AHB_HMASTER_PORT_WIDTH-1):0] observed_hmaster,
    ref logic[1:0]                           observed_htrans,
    ref logic      observed_hmastlock,
    ref logic      observed_hready_in,
    output bit     is_hsel_valid,
    output bit     is_hmaster_valid,
    output bit     is_hmastlock_valid,
    output bit     is_hready_in_valid 
  );

  /**
   * Execute signal level checks on the write path signals (driven by the master)
   */
  extern function void perform_master_write_signal_level_checks(
    bit        checks_enabled,
    ref logic  observed_hlock,
    ref logic  observed_hbusreq,
    output bit is_hlock_valid,
    output bit is_hbusreq_valid
  );

endclass

//----------------------------------------------------------------

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
OJJb+I3UbEgLWow4gmC9DJpIBAMG1W5MuJ478Q0B14hlsZWx9o7qa6hf9HDd7gJO
1UwKBKLdjwDKuV183dOUnB08/dsxfna85XtHtTJhlEHj9wx5qcdTs8eEiUVGh0Kb
sblDp2+ZXjVtaWIryF4Oayg9engUjFnfPO3Dj12Yfxk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 24457     )
b2/TvdXzUquOwI9RqgSLrtIn60WzjN1DW5i8PZnNAgwgwrcUnBW03lgIfrPXRq9/
xKPmO0mvbhT9OadUKZG4IV39iMj2Fk36yMPjTPxmPNvvu6XGZCHoHzNt3ls5NLKf
OpXZao54WCNkLvPElN2z57nSf7Xk2g4J7wdyQmRtAv4jNnIibntRo6wsUcXEUeHi
G4OhuPI7XvKLZWeujqu9M6zRNH+ldwxwf+FhxBza8YWSVESH2fwOtVibJw7Q6DjA
+tsOsjSvwXoRrMbVZfPaOjhA7F96m+BXyIK5l0jOyW1G3SsCMKwzoKMJJSkBeqGG
p+qIytqUIR4ADhrT/CNys4y5qxVjvKiCJctHn7Z3N9Qp+Ne49yO13ZgmAJc7JMEM
P1lBuMfaJ2J383qA9XhPIjKqBE7SQJ7L8DqX9xx3vrQ/I+BhaiFiylSA5VyPrVK5
9b3Ol0v7YcydUeSbeJHwrtKswSJ3cpXKnVKidpF1ZjaryUX56nkvRaek2qxGwRLh
pWndFzc1Drp3N+z67HCj7R3LQx4UfLmWHRd6JkHiCRoO9KiD/3MguL+oNmfc37Mq
xxRQJfHMwPT0BUH/pf82DUr90rVkFkdNCocv9X5FhWQWl62eXFI3TaNm15d9aKuR
5IW/BdX+nK1GNdlH17eBoBTiocTqf/GlnUhKPFCO2PyK8lo0duTV1u6Z6M7Nkbnr
UMkZpF5u9CgtMgUKQfQXnGxdyE4P4jrqyATNhvnnMeQ+gicJvVQ43rQnpk9B//CY
t5y1SEbeZS+PpFK1tW2RuORnHRAHcs6LQm1vB36rgO4PZl9Tto1szQjIMZi+KaRJ
1o1br1Y27cxlMF2q/GmuTrkLzUaDnFbNY+M0Qh4pNFzYfia34kcrJ6Zi4Ar5TK6z
yPN67IAyeU/+PuACz4kt4LHugslojyvvOxWWiC/slSZeLUysJ8dEt7NQtONR1+I7
0UapyJQElevpbgpU2Ag92lvlZQAXKvTQXHB8WA9dNf6h8S/A2UxYHu05J06HlyVH
6iXUrVezMzYgi/18H/VosXpxHvbGhov5xB8gWpxYoGXhkeCBEXE5SUl8MHogNPnb
JGZ9UNTIdL0ydFbSHfZbshHtsPlWshRoJBm0jQ7HPZgDgnFzIIIe0gav7vQtSLYg
Tcw3s8cte4UFKHeibCsgVrEoxtxLLnfyPEKj3R+/edZX8Cj3oI21R1N9FZ9lRgLI
baZWrLYv7/5YWfVg/jDnYXZ0wKUreO2YidKk/1sIt4IFFUg3Sko2/1K0i3leff06
Rfa+QrXI4wp2jvfpDjAGCU+7VKSfeUvgxZwdRD/I3fSjojk8zVFMHYA2e4Z3HDel
BrYkBdOT2o3NkBopMxqIeN+dMm1g8RnOUlAyPEcytTEwKpZG/f26vTEhCNplCmFg
WslLhXplDcr5nKGaL9GldT/bNsC5VL0e38Z31FMjjPU3SQXV2cK3GjC4q75Hd+Pm
YhEau0gI+O/NCQGXwOD9usE/K8y6IgcjyfRGwbGhzZgdu+8/19GOZ7qtmRtIio6t
dBGlpx1Vg3xj0v67SpO8BkINi8zkmwIoYBWRDfM0a9uJxIMSB1CDuem9r+EASpaf
GSCT3jJG5937lI2MYTCHGMkWKcg7MEueKpsdOWuv8mQAg6ZRwiGoz1DtTimdfBp2
nPXHKPhv9XHdr78k24PDuUE9PeSfybLWX4dk52imoQomc/fWL7qq3/0BKbGcFilt
zZTsqctgOxb7615vB/Ur4g6z4pt2KIg5iT/i9R4WYFyb70YLDmiPkE4jDUh1xYt9
mI/U8PPPJm9z6IuPfXmTn4jPm1X2zyGWDEoipAlhPQgM6dDyun/PjCNxIJqGTj7I
5qYwEQZkGBPL6GKP8Ew8mLla90WBt9xIV22HuQnQONH7QKjEneK8wlZ/FkfmYcn3
i4uZDc7Y224f0vQAs9qGBqRyEBqebqr/pM7NNSRhlJxBhwNbAm8gHe6GZNhmTRY5
KKDAqROQV3EUvYoykoQ7v8P1ngsdMdBToot6SBWQAnucFJOJhY9K7p5XkCU3FWxd
5t/A9hYPNkTROST7MPBqJ/DuLKlcg4oIFd19LcsoTN6vXP3C63kO9HpoAwbZMYi9
5We/Z9aLZIdmbACH9ZijOXJmfFUFl57VIjEpTpSX44u3P0dCUeIXRGeQ8ROvKupY
OQhj0o1gTxmhEKLYNHXT+4azRYI6YcSnAdPHA7V7ZYuRAdSy/VHQenKOT55/broQ
61A5OY52gP6y3MCUXiA7VPS849XMWjpiozdwPIlW/PG8aPOB9hPFvNrBfFy0A28h
uK4Zuk9n49P+TIyh/qvaHtgoGtszqUnR+PdzNk6CtINw3Q7y793h27thFD7za+gI
4Q+39pHyyOibPpYTiFX+i2ozs+1W7ZQZ3w28mP5esv6pqN5hTrxx8dACsCVWL2bZ
sQZ9LjAhipQCTiMbI1WCkUYMy6N862HzbtS+zfvp2ULkLpHj1mkl+Z1EV86PWOt/
Vu2uTdqetSEmTZ0mua55OB++L2tdV5YRFyf/j7ON8/wm5OUn1xbnddZ2EMhXfGGD
HG8MlO3ipiqXoNxnqseXiMa5zvJ5gvVrIjwrxQHv4V4AI6jegORGC8UPARNmYmSr
wF/Ob/mt8mEszLWllBIdzd3B1Sbt5gAKJM2dWf8233u80sZhEwhXBGVQ4RO++Z48
tpVf1yKtpvoIN6fgfOhMLIcNLgf37ndu2wGjiT6dfuyRsOqAoEF7avVmfjVDQi6M
8C/d63NHjnNItzExgOVFgDQbvBPpMjmKl1tYBWtzjo/vt8HFyW5FVvpvl+5BLtwd
khGMhxvu5FvLOWEAD8F0iu3RbRZj5YkcMWCw5FIsvXxqsXRCqhIuXPlvWY/7xFh6
dH8EbRS84gvyNZw2RyXRrb2dunFdyi0Y2wBsXDfgAiyP8TfnW6rqRqVOvi+Q2gTZ
Ou6UnSuB3+NOHIp9cXZDVTvskfTiscOrGlqAZ1Az4PZxKhbgNKTAxrURTXj79jwj
+onMbX8ooRCyxQaCniubZVpH8KW1Ty9GRRAtX3a8RQSCw1XdE2Xk+0jjgQJ7jl+K
PIxku71iT3bZ2Jz091jrABK4P8LvD1VSYJXDjux0/98p8SPKwk63mhjhJ0nkfLVg
nSqsG6fnAfd+MpgMO6l+1NK8ulKQxHPdvf7SlwtOlhZczFjnIbYa4xH+wtdR9e/g
wxexsAwW6yyr0TRuSacrYBYq+PjHuARMQmrhub2+IwaA0DVWYOJl6NvHfbtqLsY5
yrCHWRE8tvColOrjqWaY/QyHzIV3CqiG5s2BMjcVCIuKgxPQivVtumRJpBl4wznV
jvGnKiz3Y6t9e1GeuMFhC/Fz7QwVGZkGxRUaaOwVbciFCdYGbDio96ltJoshLtxe
DqbJBVlGHGbo8iZB4J0yp71qTcjhST1o4c7GxblAmlNeHoSm51sdqzcgxJAhvLBN
/XKH9bzAXC/mAxuAIZ4cNRPRXLnmdBrl5scS77fPOH3Wl/3ggUxG/V1lUoMLafF6
zrQyQDG3oHe6kwi16GM5/FMcAZQd39pFjaxsdo/fEv1zWfASyp3lifv2yrbF/SXA
arJOHDuZSqKEi9whT61nnQpscNCv8vj4LYQDr26K9PIAP7e/7VzC80wzZrP9xoWe
5iVWSP130Z96mS3Tggvy0TNtW+84bWOkaSLTSCtXj4kxL/2jicJqF3K04QcLPBlb
+x9dVY4GOKj0pVZrKPgREUrHWOYCgO+dY2n8MCt3ERKmokPd5xQ4vINwutN/ern2
EKmKd+uAkbyuJ4fysPGHKqy99Jlpzkg/iQd8fIt6S6z9b6wLMqyZX2jQE/lYxJeg
mnZUn8HWKONp+texaBNm6x8suWRhYMq9fS3lWsiAU5JARNeUvQ/x4oQFhXDS4zIt
9X2SAf7Jln/ustK4jl7g27FiUa5IXIUONNmDQc0x9mN1+21yEw9bGj9zZW7M5kB9
N7EiQYQAhgcRzILeQLBijaz1pnGzmYnjHlyYf57HuFasoyPukiCPdyUaHrYJm+5e
MpZ9XxYXYAzwNvEGffoJCXCdgVRbnS4YMcDQYfkNsl4L0B95nPWzLkJgqD9G/6rt
sGKMM7f831NkWtD/hqtZTE2Zy+2Iu7KmblUuWnqfCVyTA76dFemTth+aWisdiUUe
QCUyb4JkseEQGDrlJukSRhXDfzvUoViMbrn5p1nZlMPL0fl1o3aJcHSepsl3lVOW
j1dkvczSHXNkNHN1jvD1wDaovSqlkLUPjsUWGI4pUCf8CsadqGsEiiLLgHPY3wiW
4F6N7yzeYLgpZvs/aG4gqYG93R97iYa8O2gpO0n2Zf439D9d7mQayNcgf/ihzfDs
W7cshsG+CbwhDxiEvNoy4NskSMue04NbgHAusBKFVJPYDfYpNegIwUeESe042+ah
KxEOdCzuPBMGx/6oNPXkzJpYbd8aHD59JC/a2ZV9WdkR/T7yBrrNFw6EwG3uZtzE
i5Gu7eifZlTN/8sw4yDJI5SzOxmi63A4ia8IRj0td7DiB5XH3PKlYP4z0Ruxvb+G
VmgYo2S52J4BZpsxyNLQF2cjsKuY2waK5d9VskFt8lbHFq92iIsJkdA5S0r08ttr
1hjglXNb+yF0ekwouWLXuV4QPM9SWqCkGJjT2NBDKfwgV1aw+L6MEHAH0QZsHW6m
YZs1ZeVeQZoD7C6L93va10NfYEeEQZJn95hKHwkY/Pm9dmGUgR7v7fqI2QsvKIKv
oZs3aBoysIUFGKUcT5WN4riEfPDpuHJ8vrEi1ELdA64pC3FF2ki9cKaZSOZ7p+si
IdsFPdLFGsOkc7j2TYGEje8g2WldreBcU0bRiQqyAHMC8Vn80D1R0juohnDlnGpM
SH477+lg2zXtaayK4n2gEyU90wRKXYEwYzyjUPBXqZyXMdRSL42IvbMN0mlUpdc2
k/SaMzSYje0FQJ1GmB4cMbmsfYGJmRRItHaPoInnBBrmo3GLP6y1z10/GSc0E4TW
pG6IHR9nI4BCBiyOos33SD7YXEEA8L0TWHPS8ZKOWoaZ87EiOjGADLCbkS9dQI2r
0deai9KlIujgbKnsfitPP0RnGXn4ANVTba+3zDly45gnfNxZNSfI7mHf4VtPiY30
ZlM+QvANuzEfoILWy5F0+H1bLYQV1TqhAo6cFgFele1CWHjQXuQN3sLEesT1C739
s0NS8lftIi63+vz8l35T8CsVU+ij8w9PTMGH0pTZqK8LxxIe7kAnTyDtPxtdHJKj
sO7GP55Yqy8rw8seObFvbnWPvFxgI4f3RNMGiJMg5ADi8oV0dYZLtO050MOn8Pp9
9V+6YjvEbhYb25KPm/aZKiO9zUFfCANzl9L3+J7Gex9iTcBsZ2y64KwLwFUhWxft
dilBts5f4m4aA6JNpgAr+WQ8GkZ9HnC/jNEJtpMqbVYkbGpKOJyuXLuckz5tKfeW
NA/fpX+NZnucRgNHfq5NEDdcHYPg8S8ItmUNV6jrbPzEtT6dMyyG8zMMdjrNn3wC
tWP5QrVJGl1LiZtbdoOXq6ihqqcZuLj+nWwzjupPBw5T6MXtFRkiRrmQW7WDpkF+
kcN+JDWAyFlU6OQ5MGj8pJE64Rzr1YR1XF1kCAOJec/DRnp9xucWn1k/g/RGJBGP
AxnKl7YxIwZ5bS5fdP+KWposhDG9gcj7OK1duCbmo6V9Oo99rns5xkQXzzsihJTM
qnb1Vn7t3PHnWwd7xghjskTsG/rS/D8K0LtStP4iXgUwuHnqeMQ6winT1AOTwBf/
46NMBtHq3zBnyr2a3RxgLBcTUAgL+JK9eDAs54XfkJFNHzGhFUJ7cZpqZCkw/oVq
h004g9x7WguJdLDqv0v4U8xz83Ey5iHGmKPRU+86ovYJNL+cbOyhji8npBFMQCCv
OHlA2B/W7hL4DFEfObBHsZdnUUoukGp9oLgqygNzJ8xrl1YfxD3GN31ILH0C0QR9
ulGu9e8bIuJ/FBltXuONYRWby00Pol78jWZzA6rFnXgMNuUa4Q6i5SFboAFZwjqC
A86Qz9s+I1I7Ec1Jtg5TQz7qUSd5BothU4PkohAhdakeSBmT7eRnnueHSjxjDvF7
hFU3OdHB9LWK0wkj80yxSqbDiF5WFAPpR4JUbq/N1W37wK1tt8Vp1SyPk5C8Y9s+
PgstY5rfaL6wifRrVBdbmEKUcYibDCfQRl2y2LGm/sAixbVENaReo0RNTURbUayB
iiWm4+riys+RzytlXwRBWNX8LGTp6ukzaCC3uktQs0a1Li1oNTaLMRmzD2c46qCu
5Gnzx2zbNmsgPxDmIP3s8e3fWiJo2Mng8xYLn2dEEeQLTNjpqv0+Pg2JjCuLe/ex
XDkPo0AswF8D036yo5dcvDulR7/DCsbH6aLgGqXwMvk0ITZqlSFXmcbK/0ZYr5h3
ZvlVvulfgAFAEgdpgcZNXOEwZUllmO16zpmJREDyLmziVnF6mKK6CrM8XLV/P9+1
ItlnkxAG6FgxqLt26/PIgdRKuknG+JGUYd3am/9ID4AtQypj94kSKkeKt86vQf5t
T7CXzy9NifGrj3nbTsgXsQx12Vvszt7okPuhSS7FUaL3lESyflfmsYxyPzCodr7Q
8+0kTmYsZ5rScNaDfn5/S301OnKvTELWm4UAEHyN81YIehPe7/4uYPThbn2nhdgs
Vm9uVFTPAuFlRVwZddEwcO14CtFI+ky7D3dkyhriiWNJXKcvHM1xbVLl7l4saoUR
o/bBctE+dsr5+MoB61oIODHW4gGikDm6XivSYacFy30x9ExTRin2exsbeAJ7IFAc
tscszoRXfjeXVmfqyjoY0C03SJNTAzD7ytvZRx1yMjhHfKhs5UyY2eT00troIETD
PcGIadCJbtG4HBDgsb81uz21EdpvYHJH9/sEehq4vE6Rr6GB0jgGW8l05FyzMlgs
D8IBn2MLl1OX8rgCZd+x6no5BMGMRIlolgqTDVKcxKuCwNRfbhKRPh7lKpbo6FTY
5hi25fs+9bhCNopVMHgL8jaHM3buxpWpfkq7r8rZK+MTUJLZp6jLzjhheCvkrEia
rUl7koPvRRD92AU/xXuVIXj2l9dhUk1UCoGcnslsvED/r2417PvXOqgRjkcyE4ZV
VHRKDfiU/dFATnD1XPCHbpONqkB/GPVQMbMwTbU5VKgj93sRwM2D9Et2VTpbNC3j
XbhznUhFNxsoViGp4Wt7f7eNNeTwz4EzffTGVmbYynFBZyIsxIO22pkIUpmA1dh3
53/dhWXGvyelMPYNrgF6sQ5+T5yQKff/RLjh5qje3mQTp+KqfbVF1NOF8blSt0ET
92XXSUMZqgsnCnGNhMZ3XwNHp3bzP+S6wIndP5OrKe5Hb5MOuW1pNMiIk/fuE+J+
FLQCdmuAMn71OhJ0OYr+rVH35Qov66yFsOcGmnzRa8KMLtbW0WLGOdCjZdQcln6B
M1gNCBS79nwerjamTreaYDpamNhvAWasGqKRQidrWd/fC9vAjTu1JK9zuki09dto
U5Ds7aeqNKZzJ9ouNBmwypnS1nByRBpvOycrzwcY0gjYq78lIkXD8sm0onBqe6z9
2BxdbkbMXOLXgwpMB/ZWTHBWrxnIvwTjWGsUt8DHLuAbmSQgJzsS0KBIsMkZDj6w
nuc8oanjcJqamkeJJXyuVm4God89EmnOeZj7o49hgHgHW2m9YTfhGKub8TTvyTJp
Jt2amXd6WS85JBejlFJJEO65naY3VegmOYhBm5uGAkLJLuDb7C3I+V3hWOj5Esjo
tNF/1YDzoR2+8owW7PldKGAwdibgrmDJt7LBOmhA4B7BoYm/U4PDrSMLJUgP+czM
faUJj84mgXDD180WmVpdXPlm9dXppySTg8EjB8cvqew87QUoG1i47xpRgiQODzSl
eJJFJb5U0wT1VB686Nj5lW+hkxhpwqwp2Wm4zI1jXRRYejGWFQgp9EF9VEd/FAMT
oAZdLgL3QZ2OGzK0dxh1znvZbs8iwfMvA8CPkuvt1GYN2shq2y6qrdaasf9++EU6
QTaS66La2I211myn792YRoGBb7CWU154OS+Q56bWo8no11haGaZq2fdx2E4JuPe3
BuUWwFG+n0GJ0EfqMeaWs7hSYqutMkvTbfdXTEubTb2L0b/fzVx/2YryJAMGsvTr
ZmoTscwt6w9S8mHTybIW/D8/soD1xVPBRDZe/N9SXR3l9yzx+warSnksLs2UrLeh
KESZ2Josalgx32w7Auvh/UlgSjbnd7UmnbUMrQsSit8rhhNvPKCV1A0DeQ1a2iKl
4fmBaDMh7kmmoUt6VAVB/N4U5jSrNTb6YEiJSgKARNFJNpXoWPtYQxJ9c/1oYY2K
GVI7o1Vw7pAAlT3R+0i9HGYMDk2XHHXwPlq5NshxZcaIt3FAIk17r63qk2M6H4Dy
mtc1+4d9nIEQPbx43Z1AUthdAyTu9pE4WYnq2Ef2NNcBP3tgequhuPIdeFNZsJSE
J5QXQ5OxrrUtLShlcXXmd86utb4IJjwLiBsTOSMU0z6uitnRvaiCfHO39L92QwAX
1grEUBCVKjILS4lyZuuN8PM3xrPJ3SreI41RJ7dx0Po58o/uVStg8CeWBwXmeGwL
bulO14IqPSSuiDWwMbZVJtZe240+ya56tmFJBg11DUIMzgdQFt1jhvumyOrizVjI
D3kW/Hy7rgbBKNSFuMFBbj9ohiu7saJeyWGPfKZcOv2NS9+JRemeI1HPmt2QY8g0
m+c+NxyDPyuzpXcR6q5LVukogb6NE3LEFx7QI+hXjDfk4eHOfrvFdrw3myMKOZIu
IWuIL0xEW9hk57Y6CDPmd1mzYp72RZXAlS5LoBPXm10PSoBgN6FDpXt89t4qD8Vb
uCwXtGnaeuF75R+2c8KS/WeuJ+iy+lr3ylrNrVLCm7RfFiqD/g+K4sJ/P+DwDi+c
alOdZx35Jk1pQDpAxEGPkkYhXkJIy0o4IorUPMVhliPHfqucY2KvY9zRWm+5Ai2q
5lf6GO7BbYFBlm5WbK0qg2MirFG4cb7kOpYlvY9knb7hpKt5OfcZIWs0MzAhkei3
s8HcHYFOGHjK/cdMbmXbZO7hjc6WkCJ0ybt+UOKfGVHR7QP/UzO19NTDnrvlvF3N
J9yxQfGNq0zCNhPZbrXxfVWR9zQ/s/JSWfuTW9R4mLi2HXfYR0nlTH+WzpWRAGCZ
mPCb5n8zZ1sc5QcHMcM5VM36RPUOKcnj2eJ4CnYnetWvMOfvPv2qgWrM27S6bcwp
Dn+vilUDBrmhZqr0d9nC5kDwWTvxUFLjYGwCy+XUkhgSTlDDSgteAvGVI5uHeRLf
5sLY7u3y0uFCA1cnWGB4Cs4qZ/RCyS8Qw2KZXJHqRK8EXUP7cwhsLptuHiRX/aBB
Tc4P90K2ybwb46rGbYeGcsdmnb0p5GFU6evdHqstOizUmZ08XWGCO1wW8MqGeMG0
zmSwEU5DGqo9XirO1Os+SrJMX0dHsTMvyMKtRC9CZy/oqoWCTRkVsNq8g0jdw3et
4l1o9cypJ9eWdSga6yQA4LvpVyZ91E44nYMUX9Lkq1BEPOdPnx7PCglz9uK0CmtP
/Sh433DWAHLAIsIEwzbq2puP9WCxzrL0q/RZ9zwht4G4llySR8aQSVyksnkLY9H9
DhOv3iAC5KwurV+JJggir+Cq4ibDsjbf32YyzLHqhDGIy/Ap8dFCEnktC9v0MhXD
5QrPcZAPFIs0LCyoTjSey6vlmnvSOu2wQNTPIyRUUVNNnVcd8NZNQDLttMqUu1Wq
GR7xlheqehRKBZy2FIRew9AfuoT0DLraXVKonmcdPM9+29KX6XwA7y1mdcGpJseR
KuH6TN0JJ7c3dWcd6cRwl3fbNiJo+pI+dcs9JJZZEW0KH3OltCa0Mp+dHX/zAUiM
x/2n+SYCp2rubb/2wFIdcGs+9xbpFeVoPXI9gu8OcqnOwv6aWIwarEtNjXGRzusR
fPQSO6Ef/7OaAeiVIqiXVDLbluwC9DjZTeKSrhlumh7xBXaCrqIhSqtShzbBIY9b
DsSg8kDXuexZHyP+v5PEOlfcX3Wi5ZLRwx76ldo0p1zlwLhCKI6WDp69L7+e5yQD
r4OTdQelWA69MySuMntHz4/rT7xGIxRD8yS2/Ko29sfbzQRiKXtyHNV2ykiUZ1dv
R6hmN/Ncm8KwlS4xnGrIlBUBk3iQI0wnYIZOJvQnEvr/NscXH7jnnTHJOQjBQld0
kg4GJioDclx8N1q8xsq6f4rV6tRSeRp/IMjMZijkva1lllI0sTTwb72R7cgebzN+
rGsRMCXuesppD/Q0lRvjkMTpwH8FzHCmb2Z6CH5JfXZl+cp3SnUwVxYv+o98ejvb
/sDSlYa94BeNcVGSZkMjHmjDgrus7csakPEbhmuSdYktyHMf++aZoBCfSr7B4dkH
yVqZMSADuzpGnqY2+KUuuFuOxMx5b4sXF/EIQ9BaTgGGXsfEVz7KQIwdoP22OdTy
sOdklV36dVP0zYx/8eikqhbhJpMpqGKfMq743tBgVABeIt8I1/9HKDYhPF4ev+Nk
xPu+hxXdS9a8vPw2a0mzUvYGCGIv6Oj+fqY4CJDRgi+P+ArakxqCKLjz34+FtJ+g
wZZppbTc5pUM4eskJ/qjjqz0l+iLGfdCt84VMhUZW6vme75biAahQap39c0oPMVC
FRZbsBhTkdVA2FbKCrgNqgoq1ye9aaBe2nK/SpK0/ZrkYOq+EFNyHC6XGSpl+k6S
JbPoPTibnrtI4sOb9UoKdqViiE0yGNhHQcmV/TnlXciH9bwraRqDjOodAe1WT1wt
A9+OOyaRuLG0B5bczC/PAHXAoG6DP2c/R9gTixgJ2AjekmZE7qRKttGq7JtvwLxR
P88KoPnfQc5Pr+BuGOoQUljpG30Wu7EdcJHgK+54+hX6zzA2oY6ftYLMFJVrC7kv
oR/2R2p17n5jJdN0oR0l+kS+2WeCexP4dAfJ0t4Xgu0XpSb8En0fGZp2btquLj4U
r57mXv7xhHS94Wo5BG4hDEuWGhhQq7eWcH0AIvr3Hg9hpn2ULvaTbxvHaQ8RHS8F
tdvS9MlhnAYVj1SV2y2/VvhimrGd16urj736/vX33Qzx7cJ3vc66Po3cx+l4+DEM
0pqnqyEOv7HbqZYgOJ+Kjw88ufMU8mrFXtzDfAW3fs3t4cO0EOfGmEmJtATTjORf
g8sygl1c2jHNtfIVYALXi+RML49IigbswadEpVyzSLS/T4WhVIC22fs1DidZHHWZ
D3+EcEQEpf8n/X5rOEMLssUS+65DZRABsG3H4IWLpmhdnDr6O5nLw+1jJmNnIkIi
xK5emHsX+W2So14atMGA8CplooQ9BjKwlfXR4t+iC/eDHnObWLbYaOnrSShtADwf
dzt1wM1jFjYOG+8jHz2kdOC/M38k0eV3SMn+UKuNDy7EwZ2W+18wH5UnSQX6LKOu
ESUMMZ/lSuoaRN65y+CHGa16rJu5UGKy3zncKtEdaNBUzgf+xx1AupRSCziQ+Lce
/8gEs0kkgLgRAMIjXxN6IPSNM4UyaWbntLgwwua5BrsxpEJNlRJvjY1mGKLnwXk9
QI6QrwXjBzv5b3LxHqj0+YB3owLr+HYOy7F5v1QjNT2fp7tEJGOgay297b3viulX
gAXyvN3BmmaAk1vcICzt0CC8Yiw9iVPd0k5KzlVjhthOGI0IzCXrr2i60P3BO6tG
ykhUkXUrF8myYh2CbplCApnq7mvbIPvjodE8isoiMAeYuDH/gMPh8XfFFSe9lZ3H
byqN7sVW4AUoLiInuZTrTdt/nuqwteBS5JYDsReOtgucPWk0eiLYJcjKy4ZnxYZG
BBzy829qY8qq/HekDtF0xxPYsx0YmM+Yed5igDDdPDTrvZpX6XcXa+2qzPfq0W2v
THpHHl7+yLro+cG6pFqFYLihghexlKTbIx1g8jUB2xJ0xJtwbruF1FYelHpI3TCJ
9Xb+svHYHX4qAQsSZ6pR2I9Wstk2gFB8IUF4Ow5njfFu+2yc3KbNLubmu7duT3sm
HeqKWHYxvaNsYdQegGLuSD9tyJnzrb0XbSUzvQ6Ir2hQzwortfzR/ZNM8PyUB1u3
GNAwI2ggTjzylR0evugchTtNt0ZxI+sqWj84BEu5d53HjbCZ/G/2FgPkq98AtTVu
/RJWClhVDEiwjY8YCPfTIWzq32DeUf6O3QXwS+tdhCQarP073WXsHjvUb1YTEWGo
q1NBAf9ptFbZVbu13ipcT7DxnQ2bjUWU8IOxO3a2mOdwg+O4AF6oavbiqtj1SA0e
0SZ7EVK/ZPXNMfVrdlfiCYv2oWd0ZQ4z+GUMONkFU6E/nAZARQkerM1oBMmpDj06
blEdhuKc4Wen3syV0gjQSabZLCxc7nVnPAeI+xYTz+xpUUavhCCJj73vZy7phglU
9H0zCh49Xgl75x9rkq0jZddvtqsqTcCFpYufvAwhgmRd+7zG/ssjW2JcdM1kGMCI
43HCKwnWohZRX5XuXGG0vFnLi/vPuWyS9FTgDVTOxrMIFs3jWbyPJbfKSEG3tmE5
IvjmrRmBG/kMXB/9o7N7TduhuBAmoTQVcT3QFBspkrkNSEsrJ/0fd/eNRCM2W4XA
n2RHoSU9NU60+Wrbgn26OB8+/NiW+5IYc0pb2LpIe2fV8vIfJMTCuYCSrTVIf2ru
7glRsIjBFxXVi82eRnenpYvM1Ig59WOyv8OJikA6gwGsfbsD3ksaWF5upfuJbTNJ
Z2rpYObWiMaoDvELxmyNUtpvNnfeuN4IYMpIrx8adKMYrJmlht844fh0cH3tsTYV
4wxZ27Rtxwe08e/cUC3OJutPl+yA+9pnpeWD0nIZulcfKqFNbj2DanoxNgqOMmjR
chdeVVKYC6saRwLXtQbhlNwP3pBAIW6AkuuQxMuSm5VPhiLE/Is1NkW51AyWj2ef
tCYCeEp2iYz7WQWeW15+4g1CCwBzKVrvmf6oayudDoOF7NQ5x79eR3CHm11C8+5z
gWn4KA9GXxE8/6c3xCFtfAKprEzS8BMB9ci6cRzUzoVLkDRIyJirNyRJuNzYn3At
Deu4axBOa1rVJ1+WXwYzcfqmfY3PsaIfb+IsbXk2VuDWtYjFhmws7GwwWfqk54pU
cM7yBc3aei33XB80Jaly7n3avsgWIB5Bzsqcc/CYQjr6ZdPv45YaCNRW3ti12Nqr
yVXVxB3gTEkT5Stqe17WgoeRvBLsNN6FBLz2V3EyR3mruU8GSjcChDyKVOsxjVB2
sACOlAv4ooYEdJWRSXisHbeyL/pzMd6MaAJ5VbNJ0Z8Aj4+YuRBdtQKn7qr/8yPp
QMfxGbUXiVopfIn9Nv1aMrbweJSZccoNEWPh8StOgSHNW8J7qMFAVIHCoPDa5hCv
olW1z0xm77/CjtJt66ShC0XxO2e2oyErmL5HXOl9Owpe8/mJzwC3mmUIWEMDPYqZ
oJhuJpwG9k1rt9RvLo88iLMl2keAHsqtx6OAfW+3y86TbG9jPLX8mwO6iFWgumHM
NcixlPlhAB11cD+dJvviDHBwlpCjAAUHBEkDfJO4qzYsnyJ29s4C8RB9cscaKnyq
Y5CIfCihEZLTl8U+74c9D8MijmrAWwRhePpr67f7qxZ6a7UodSODUgloqUQTlfnY
7lRvcG8I+ftYueRfMEZxx0XW57hHciH7AKXOkJSUknvbtIcYQR3bpcpFSGNmcJi/
DypowSZpiBEoFme6AszW67gnKd26sooUYnfWcwDLNykUsCF7hlsz9H3Tl4A962re
7ALZSzglzroh54FVezsPNKFLB3wpbmLaS+K7Nru1sAnzArXOmX6r+ANG8VZ0B+P8
ncizD8GDPnVWKFh1bTFPtdyHW+60vqMVGV5a+m5DjtKUWrbHv/+ZL5Yly2jb4fED
Q/1goyMw8xahUyqVqcoEtnDRwhzT3xtUfL3DoHtzVdLJE0Hs0LVnxBcUdc/Af+vp
uNpAEi0N7+Bkup927fL57pHRc1urHNRU9C4pArYpsp4dl0d7Kbc0buzLt/rOJGMU
ieMnd8NMw2U6JZnhlEir/0dsx2VGjwRnQZ6lq0ZiONiEVCkMrOTLwsZho/MqgoF+
t572RwZstuHzmDTeRpCHklO0j8JwPg0l56qDKDvru6ohDFA8LOiazIL2zPsHMvU8
wUgqjJ6RjwvsUibAb5Csq+mNTTcyKhqP74MHAIUi5UrHEmKKj9fqKjjfHQ0FEDXK
g8eQ09Xuw/4RkE/foj6VOWK2RrhIlj10cHufaHRL+dh8jy8mWIv/J/qPHfg2VyxJ
c1KYeRz2YHX57qUctS+4YWjBxWRXAGL/zUZiNLXtTeyyWsFQ5e3ExU9nH1aSw4on
2qXJain8YGFxPJgrLqEOALnbWCXeviXw4mnlsi09sdvtvTjgfo6zWNADQwzZtRiI
eMPKurGglcLA3ugdkckWyfvuIGX/5m4oBw7h+ckywfWkDXi0i5keA71fCv0v3JCg
wO4B3SG9rFzVsEmqMsrgF3xQtAlKKFKW2vIsvQgiXypepNfLrJXAyXYcB6ukAeVd
BXVtuYnnrinUMbz61I1gzP+OjgupU81y4NRberXEHRPo0IVJDLfa3QgiiJNBG3tt
iHkuBG2PGI2cs0mXAukGUwDk00qwFLWmqFjtofbcil+tdt5V+0twnVlurzmOMY57
YNndkhzMy3QKGDKulZnuBTvGX8HEmLHyH4Ti77MiYoDQg24OmrXJnHtaFGrJ+6Ro
XSactcvoNUHefNNBeePbbBYamJuO4F7KhCYLLbIr79XdLIJsNE05LUKC0LKesyNS
okkmiD5IfcVROemBm5yqgYbX0o0vUPIaAkWMx+utuk2KcEf77sTy7tkHIoM4N8er
rfMnG+knMFmSIdtLOhX4RPon2uNS9+cNQ4lt8gFcFuHxG8ymwZD0ecb6/04ABFIw
IlGVmaHbzzDh5xlJ9UUDDREw2bq88TAkZx+LT0GYWJSK1Jym50Q36gz8xP39aGWs
iuq+shOSc+5F7PgJOgbZh8bD7fOFC/r5K0nSbahrjTEuK3Bwcm947qg8QAkIXV7p
lBQXUHJ/iRQvVJLdSOts+vt5HTPuL3iL9AA8CMZG8IGWnYMrqDUrAqsd5WBifewi
TVMwsjAB8kUYJe/9fJZpYVAFhJ8sd+UjsC8A0chxQhWmCXENC+WeNE0WoerlYSXg
5ozstThwalS5XDAuQN5io8mS4Hi4+gC53ed3POmL40dnfoAzbYqte+FLTpftRDze
nfJFWqwXKKz0arEm+VsbIVv9uBALEehLEpQhvM2t26U/80UXWCeLsmT+8BCtEvwn
x9dvFQDouYyWGciBhYFMoBaMKhgkbe3Nf7g0xV5SbLNyKcds/2gGGAUae6yMkjRc
TaTHxNBekm2e9NLP0J6vnawVnbwJcXa7dkN+dACiRyBni9dP9/x+a7Y+tJS5VFXs
QV7cfxC8RcQxTcJtcbxS1pbaVYrZVnlC3XdzyRPG0LzKKbCcXMoIwq0zmTSjWFU4
VUo8GqKd62JsVsLCVbzqvDJ5KfxztLjk6s58jcHwzTQ39H0rCT2kntCUIN2LAOtu
JnsMMl9W1VuVKwb2makfVX9sgKdVL5hun/iKr+ckeh2C4O6OQZR0wPnekE3mEhaX
etsIJQUxOwz4aDu3Sjby1QUPDEOdmNe0isHRPcdmt3jM81We6h036SPZzVcGhBaE
k9EMbLspyuwhY7or1+f4rGhp1hfKiGWQ/2DgbGAklKV0eOaIUVFWiMsu/Cm+modR
eIThpnXBc8xu1ctFiFUGHifU72TntJij4b6wlRYq6J0ou/dinLAdiZA1PpYGmNX6
KMHksA0RpR6BKnfnOD7QtoXQ12KWhtv5ulC6jZPvEJobj9SVunNV1QRf5i9bDn6h
wP6CwsHjgrQNGnvB6paSMYCOMJV5QNuQnDbR6VERYmW3zywzem+ZME87bkzRZK+z
zvG4gyby8jmvjaXnNwD/1xhgajh+XHh//JaecqLnUVfrQ5Vvo8YQO088T5wEOjOd
HGtOnWYrQl0WPXLBsK/WTmSBY614joEHO7VBrC923qvw6+ubAEKKPvs4AjbBE2nA
Kz5tsnEFZIrSD4vLxwhYTiKiBvMheap3zwabPG54W0+8T1Omy7ynnNl5pXb1LNjn
9PMkeDxsWqTVohUfmbVF6hHZtlUCoE9OkpuQEe+uD6/gUcluP6v/k4fGaEPFEeUc
ZchMNN/qXZGaeuplAxEHvUkybc/Kljg+eZKcoyPeu0kjJWXtoeMgXZrkYlIbmczC
LvwFaVKmgT4Sl/40h/+6A1+6vMPDHk9751L/bEqvTI2bA2Wjj+071HLSTxmQlsrT
LrkZQUE67pYg4QW/yLfVZYzFymksS4eaEQuF7yj0hxYNQ10BmLBPdISwjaCED10N
BhhBrBWi/cibmu6SlDvnFimEIz3vDOK1MuazvDmisBzdHU57Lr9yHHMVQdh+Y5bt
crGemRtilQ+A2rR4xQuyW92CNLvhxfs+INGNiUY6NYMDZwvPU1rSocIusGzl3EXc
9sJvgvtCq5JIfU+yh41E4Vbc1zwXkZsCKarXFLxL1QaKxazt8xOVvzZ0TkpufBBt
FTqYKvER4zsE4dYty0H8XjuGqf4ph56DCeniIV+Qs7SHTP5LRB2MQq9soM4EH8rp
mVtuKJSUwONdZM+xWfVSXnOzI1p9W0EXzo9mHQDLH6dkeuQxVpFaibxzZ5yG/i6F
rc1o/oOOdrnR74R2LLnHQExa0G1qjnbV6Oe9+NnezA8VKAHkvRkZL5+FpmVfmAcb
5aOQ2Nlo/PQb7A8DhxBXVFQpyUmX/+St1n+3PWHLPvDR9H0BMrcvCPtUXuYmVE1s
XJ0HYw5YU4VKWMrZK9XJTmisErxVaH2Rja5slVyuRxn+wSvEF0En3uRqjlygpmlA
qrEJqItVQoOBePalrWGySNoq07zYHXX5DmoEfJrubpkQ4oBoj5ra+KMA6bClLujL
9tLCdDk6JnXAMHO6ZfUK1lhn6Hok/gqMSw6pKh15I+XutdOTdUZVEdY2m3oW8IKL
2qrRDSInjhWlqjLkkzSnnp+WdDQ+tTHyTBqablYDwADGDMCXfO2xkJA+1utUuUtI
OXj5ioWCGEino9R+aGvAof+extPQVgPGpA6fBUkAT4bDKTezAOxNnp54BOiN8SMj
451wnP4EVvYz+n9PCZJ1WxdIu8cffS++Qhv2qwVCVDgmG0/fcfo7tQf8yFxsMGGD
nQXih3/g/7dI3UTkH3ZHbGKF2DhF9QPDoGngaQTC8fRHjQfUs6s/na6YhUab1VAe
d0uboKXqnh8NTsRdiiI2XMoBDZh/nH3UClS8HV7lEdVNevtiXTQ13hq7HvkyvEUh
9/WjJYQdG6v6uVrRzMHY0YsGfqpeM6KkEZWN6mCTRhvSyhhamMJmeqko70TkyXWm
pQ4DE4pFU54nBDyb+/fKAp4z62djdUHf/po+O5dXRgAQePsR0aWAFCJS5GOt/UFD
KIxZbflazQYA1cEj+j2mb5W43OD2+tAabRtdCLywEnEFe75Cy2eRxTMRa4L4OK/s
tZpAmzZRPmrtYW413/efyQ/0njLGuPjDAdaancPaT8gddtjErAxZOIE+1UZSuCt6
iZtyF2HOwtDhzVfbBzn3qW58CVX4rznyV0Gqjpxg9KM175SPoiBsDoAl4LGzLsZ8
1bMBh3bFUqOaOp8jCJwS7R7u0WqfN3Axfqrl95uTjnP8tqxFrrobYgpmiNsjVEBz
Ksd2k5CYJO7uS1KA6E06xqi+I5E3eX8CSsaT/EMtBQAqpxTKBAh7ZZS+cMYC41ny
k1+94xNxDcZBf7Sv5bjhgA9Wev/tk2VHxkYfkes1pTGy3TKU3mwpiETNweFSUN64
MpibO1Laqi903CMRoBeaue3pdGXQ17r0bBzG9On3q/J6lDAaj/YvexyDwg+6EqNM
Op7coYkiWs/0xUZq3JfTbt0X7dXQA97l9fZR3X2CKkSW820OO6DlujhWIjj0f1zQ
JXWpMenlbMy7wqmY8Pt3lVQDJ0qJBudpHe2HQASQynCsJDeIV3FLJ7wKB5G89/TB
4e8om1PMOzWCB9KJt+eJHtKQvuyP95+d3P7EE3Avp/21/cVpV+5sJdVpcKDSE5gB
bb2KOU9oQAakbJ5jjg71eg0xYFRElhonejyXp24PtGRGW2aEfJ5+7NUFbVJkW1F5
wn1+U4aP4Qr55dPUYX3m7r/pzuORn1/v90ckBsz7YgsvjvZrDQzJ7tojoMrL+VmX
xl4t6t9D7qAAN483pNubbFWJIGvEalTvDAITOn9iK4DT4M9uufMwT1/ddQ/ImGDp
SH5gCsF/PPcAWLcc4uv9CLSXmCgPTKqTEkOf1ski314epT3biUOym8TPwEy1vYm/
mqG9LZxvYskVy5wL69kXVepKFwfSGw76Bsph+ai3u6L+fz4HYY49To3FXZLyyg2S
Vf/ohuWhPS/39Kzbl9G35btIVckm7paK5K7MfHhS9cOT53ePCqUFocZ+d0jNLwum
Abp1XPhwnZBdjVdEBjIQQ5FhtXAxy4IoDpR+AR0XqrBmEXR920at+1WvOp6MlLfq
PFUvo8h9hW05seahyQTclVGYxiCPNeF3/vlxkS8OjlX4m7M8q/qPAWCke9eUKR4Q
kDPj4IQeqUTKRG3HSEzOw4j2jidj//2cdBdNZ81yJYIxzW65U34rzUkQn/07QhT4
sS9Bc6ZOr5XjrMrXepl+CnUtAanruQQ8yt7R+GoH98NPJXRP1Qpm8bxfXcT7HdhW
nov/oc7PwL/26zS2bFxyW2zZJdMojSUGF0ghTl4b3i52lp9F5ttP2b6XJHPBgm7u
5IjRYss3mg52VIi8xXGQR+naeNgjlHIkTGBuwlDnJVzIGtHax+J2C8RYcHwmnUrc
QCQj5kGkCKh48ZMAG0AEO64rjHByox9EItfKnf0/P62oRiFDFbQeC6pfESfDEo6M
1BGaR9beMyW54Qd2+wBe056QM+7T2FmEr5H5o5cTIyG2dcRfcrmt4o4OjzFFuPbk
EGXfo576cfSMBLb3sKM2BGtBCb2diGsfRzCcnQcDhsMKehd6FTUo2bdYcJ26GqlP
ftBYxy6DxrokpGo9o/dtZ8PtFBNKV/gZs2R2p/teYoNMXp0Ch4gwATqUpBxvX7jl
ZzLelczA/kNOxhV0Zjki2LuEfee37IlNHi9NLUhilygFEhw/QDlRpYRLdK+PZ955
4INiZNr68qhsJIU08bWwGu5XUcTLAOmJRl02IV24SYQGUOMZs+6+4UNEved1XEwe
PTRzppDnoNS/FJxay5ezEheUqlHFqenWzD4zUnVz+xbg4PHZUI11Oo/2M2ThyFdb
iZR8sEoPwgvvQHJJFayYFUIYw8nztuRK6os7kOncPnbntB3C7gYH8xo1iLV+r3uu
2qqOEJktzzxugQ1CwyGiSi0cJapmSy1VNi9H1+FtH17oLHNsEcZEqMvX/ePMjOp0
xe/3OxmreaaIl9n9xrZwLhZinbCLBcEg/WbcRllTg4Snytqr5M8fdMsoliEARi1K
16HJBZRBTajjpxNXFm126tYhTXYkElncRClJts4Xeo6TyOBVS4PgG9U8K5bVX4K5
hI4yOqXGyU5QJrcJkneZaptxflXxjurZYb0mztEzxLvz6YP7/YVm/OiRQiGkjN7t
V67vVNA3itkB4DFknFUV5XSOdGE0gIUe6w2mJP5YCt9080FwWCBPkAlvd0ONi8bC
K6nrk1BGSBCuDpgpXp6EJ6FSGaccrigTTtJcNS5vF33XGkEnr5twikmOQs7oVAbZ
eGZIc364L1vrkPzDWQMP3bhtFbSbem0R5Yr2zwx+8kwySK1M+ezmCwkqd/2TB06v
JP4HFpvfAo0dYJZ5Sro/X7MwSCAI8b76u+XD9c/sEj3Pzky6QtbU50y8htaXbOyc
1MwdUfE/MP2Xs1ARm8/mLMuJUCvilOWbV+JH/SXdLKDOpKPu3GGSU6LjF4OLvTPp
KnBKrvWwBa7+8jZm5y4YCxipDvYhPImD3IfkWnqonKUBpQuxmowPAKD7FkEWFjxP
fSPGAuSOxN9pPiFtSiap2D58To/YYvPIZbfaj0HEHPEtA80/3FemyXp5WH/XwmiS
464wUQuO3vMXlTBQu3q7IX+uHM71ARRwmEErWhxAD05puCb63cNl2cQrbiNlFq3K
qOQjBsP9ZfbGEWLO/HVMJOcLi0nmCx6OOYAQBPof+vVf6eOMqD5xWOHSRDXZuAyR
bPt1A2eJoj8dce26nzg4cNU9FeAKW1+5t47pwvUgDZyHx2fatCSNz7jZTzbWBwkF
QpQpy6iDw775Cg5ilUIIiy3nDe3wjAvrYM+hC2VFKrkaHK7RlorRWR8p3/d9R1vT
nYPb5LR9GDtPDvO6ySOlzr42QU6SDIL7XOO0e0cPsHFVDAWwcDeJIq2E8H+oJt9M
iIp1m3H5mKyz1SNa+gSUXdnHGLf4clp5kq0L68OLM7p3B6NyYhHtIClyTYWGjUin
yLii8CsR40o1btZP4jYQsRK7hOwjiasCX5MXI5G6FQ9xCBkGgBlDLmkH3MT8c00I
8WsbmedikgU4Gyn6WaHWHNZvHzBWgfcDdTVYX9AZQg8vbQlXYT3uMhuT+68rBE6C
ty59nNmJ6oNRCtxrLyvcIJixhiUAsVuUHlqqeW1sklRcK3VGWyTtBsU+7EQ7ctWm
H7fgQH8YfU1I2emR7Sgd+jR3QKbEywGk1sfLajEy0j6mXDGQEd9x3D/R52bhykr8
EWLOxyZnHFz0unS+TSogOdl9YYjScyuPGCwdpdAGj3CuBaie3uL6fQbsKQ4rfAtQ
pRfupPCxeyYCMuYxVLQP4RxJCCpy1Hvj1MqoPnPoY5P1ofLKnI7fc5lBGYW3OC8/
2EJeMoC3Ceb8jMRkLYoxTWnPedE19LUd3HlPLs8/fCCENZa8eiwNRrY1EDeR9hXM
lSC7buDAwqeTjwx83BXAyubxXLxSQ8timkEnKnlOpj5HtlqppZK3tR/sN/WIepYC
MZMLy0tFU3mhjE2yATDKAXBHy6TtsSeViY5Ou+IMC1VD8MsQviDeGFVt/0XHVBzy
uEO1LAYGRa44auHaVSBJNVH2Y5+vD9LfCrr1cgVOO325fFyQb10Og5xnpCLtwquQ
pQO9Oo8vv2kaoyqTmuoWW1HjwSOzuClTBpuNYw3JheduHraYkTX1tKN05QSj7zwp
wqeIcUD7j9fWUflzM5/+V+mcO34VcqfCiNInp21R5qvtX70pQqL8DkV2qZwx3TFJ
mqvneyqfIyEg+NFmgHgj+5v4A1ey8YeUGmpnqd97JPEyxkP9PynxlJt8M50zUvY3
oZ3OpYCMGMnVY1bs5gYfm2CQfn66cTnCwMH/FsrGSlNDG+0k7JIuvHhZEuKD+DsY
S4kBG2HEQfE2sLN305Ak716XRJMCjkycuR9ALe7DitRukO8tZTs+sYAQYOBPcwIl
b/4bC6LVo02M9dRSxupkJARAJWF+EUtYlFweYzY8MAvMvCXNHxsZ6Qepk2IdVM0p
hi8u99yxVWJi7KYAsvTx5HSPwqrj63DoYT5N3RjkSZWykwLC+lhaMQCxNRswHU/k
hUgfBp7viBwiYmMoCNhUZHcgOBQNqiWZt0yYR83ijvjCaKMH4rvKyl3QVprPpu+x
bXLhTnz+S7R/ZqB1oGXCDGxhv9i0aFmG2ygcuC+zWxU5wwrJdRhmejwFUy4VDyVA
snJ8SsaFGVJlHye3qbtSKE4J7bNe6CYrvVShmUS9/yflJVgZvyxJGWIm+yfIK8zp
xQwpQa+DwCkoa8CtPf8afgYaCV0lCGrjLt/PW6POwDd0Dj4DrP1No/J+VvMkHsI8
IPq3gsUNzgN/aarHYgf82sFxKlJuZdjdHSuNx67zHyHoyTiEZ7J+If+8Dkkv70kz
bcTm1imGX9rvajCgiI8AYLMFY2392hfH67MyobvcfRBx2fFFAoe2oLYSjoOY7f1t
p4SC1WBj7yFBIxaw0T55nIb2OsVP2b80R1BO9nnyk6Jx68hyzZEh1/2FebBrYlsG
WlCbE8YA+sbggynNLARkQxTgsiahRhiKR+anckopHvXtliidUgb7+xbSGZ5kd3Tq
R9iRO1/ZnXJUZC2JofhySwcncXzQc0k6I3BAPvud0UGd0QbTJBSsknzNqN3X63SO
Ck3gbkzfSYi0k6Qr6fvaN4LlIwB9NTHhCB3aDcxDNmyIXLe0RbWQGqnhSbQEF4xH
A8eJ95QjS3HwEqdpMvecYfDgQLi9kYKbvue1Iei9Rdeo0K6VMPf2fQQSu8mY1NZi
PhGebbYOBsIM14gLpUJgxeyTIhNqlDEf41yOeZbRr7jZo3qqcO6g0Fezwe1Vu14t
rV6TeIGsmJln0clxRvSNns53U695Q7HSXuDNnpgJCpG691WIY3nKPWBvRtfEpyhj
JKMWV+CoZEVR0l7LnDn8D1erhWzNUZ18UzylcaxG/sqIDGwVoMIy4b5c8o+0Wi4k
KJHsH3L9wglw4MJRLodLybeLvXSVWw76bOIl73j/mrqLHspFHSaoc8z0kKi5CyQo
ZFPk1vDtu11IsOJYKW2ax5keIoq8FObJ3M1cWzSLIobWCtgBLQrObOFi4urlbNkL
E5yEtNnjAzuWdcaiuFbU3IMdECGN63tWXrZHhebcyWhyrxfm8ADMyJVxjIWMYlk0
88N1S7F36ZjoBir0ecfw+T8a0WLL/RhAloj+mlgJVZx1FTrimqh6Q91kwDojPcd7
0zckScnNfR1gVtA5IpXvMjn4NqQr1tEXAYKUJsHNo+Z8gXDeV88nSxYEL2tWhI73
BcT4IC/yzFHyCOkxsUubz24+BCmoRbnPeNeyOxWSWVVIzdhh9oAi0N+1eks+suAz
OOI36MHvkap94Dvhvgu1jIPWVa+Jkzdbpy4bdNbqhvC5TLTcPmH7VpShJZv+nftS
kCB/jIBkrtgsNnG50YsZ07tMfWPVtOpV6vXjLLTed6n9qSV7kHg2Q/n1egowlcf2
uMq3ua0KT+ZRyUblFz+7U22v+8tZo+/mzIVjB39y6YHkyKnE+R/HY0CAZN9+bZva
FHHRHFYD67gdTRkeRIVgMDtI/+tc8bVi8ofBb5DtXdqRU6s4OCxWV6Bz3B2KjoAK
wN7KY6S38J5XaJqusEXTKF/JkBZ/lxygQzY89rBd62UZsPY2TP4kYHIHVP7N4/6J
nZHxpkPJxcRD3qG3wlRwCjzXtJRN6dVJFZtohsZJGodJWr6tnslwND8M3sWwfk5v
v0A2XVufpS9w/HwbjQTnkVcjlq+busIVwVkwoDJtGZHmXtlI5sk4NQ8a2ygFUOc5
6HbKn8RUdyRihIT2jbAdrJQwUllnVHk7wgPACXx7WHiRL0vAuhObdQVckz3pjNwf
uTahcoB3Qp28nxgEU9FZQ1cw+H8x5WpEzViqNF/QuDkS2ipcQkyuBnCPQdER9Euw
l4KZnH3LmpS9D3D4UIte6tHO89aeR6Oik6RZ/8p7LaXLaP4daDLYBCe6PviQMJVv
njJJbfb7Gd+Ey2UtyU8PjDs8I7wQPOjXqGuUSOT0g4JSe6OxQQqi5gsVaf+BbsXu
oSL+jxuA5+h7qFiHuMaL+0XRnC8qhpOhAKfFTEgwlDF51RWMoON/gJXOZbOdF0qa
YttXu25Vag0ePcz7r2VwmJEJ+46dhs7fTCRFdu7c4H6zggxlVXpKUrl7WOfeglgw
Pd2YvztEFsoiFVecYAhJQFbnzWYQSJSzyO4PLGfcPxwPfqiswie6wdmZSHSc87PG
gi82jNAdfWVNbrImBYNjrk2HyxKPZSv+3UFViCVOb7Bysz1grICJ+yAbX/4Yqiah
DKg7WI15C3ccxmxsNbDbFTmuRTLrWLUPRKfOO9aMhUZB3y6uPOebMT0JXuNRStQR
LJsOd2pJRyE/Sy2UmR2xKfu0/urTOFYbDV7mPceFZU98T4jLmcKqB1+iX+fAKUD2
/jXmEHRV4cbz1MCn6qyLzG8131Z1XPXEhauek3znz3ijHWXZbGnD6LD52UbkQHnd
pw63FD6RlG74v0nU4bpY9u9HGj6jDAv1UV8OI7rQkuzsiX4Rg+8tT/fdaCC0QaJV
VWD5JpvL5JlC0TkuLVP/cajQjGY8dygvabmXI3BExUv7Iuhse7TajBgtaoWJVZui
ciNnrxCLnMbi2oCpE9eIl0qogI4f1q+xxbSbEQwaNokdKTXc/QIbsl3UMcGrAdqC
5OLD6CY2p7oIi3VlyCV45szstKEMqFNvJblJJW3rscHFz5x9Zaq36q+Ii8Q/JNx6
v78uWupf/kCZgLNxg/UTD3Nmv2SLOrcaY7qS0Qhn6/uYPrgRhIWvQQF4xGs6jMPr
Zy/XL5otq7Yj4Hlks7m+S8kCd5N9nzq76SxyBcJtaLLLWBuCMogrmEZB8yf0UoyC
uO8XkyDK2Qjx5uGoxMg8twiNYR+Twc7HZHvIGqJTtNpjyODJkWlAIgH9VX0MsEPR
p5XOJQZV+OV6KSUi5jnv8PlvuCfina0u54vhKy9S1P4cFGJfWwgFuAiVI6CA9m9x
Jv1hTY15h5PaxpsO1NHQClXcbhqehtu8op8q2AAQ07VUPGxEpkJztbEqoqdzqV6S
AKuNN98Xjlu7lRkY6EMllqD6nqaHFqPpdr+4zkNmcDOzJlPGed34gNMg8GXiDkTN
jVAeP7VG1yROov8YdB5oS7YLWVqDurMQ4YUBu8/NdHI6lwuvohUbpXPqqwhgeFim
J7TxmYC7oI4ybO6r+S8+BEtrfvRLfjccAdrPCXuJvfnSUNC311X48QpAdj2WIOwL
CloH5GfY2Wn/Kel0oL9/uAXt2IhdpNNayHHQXb7b1yJwOxGmDWI0X7j2C3SNzybt
Z9G2FYma7OPjsx63xJQLNksTnZ3073lz/Fh7L09eN8X/2BVKQiZADx/kQloQORI9
`pragma protect end_protected

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
A3RRcvNuGied7WEYAhw9Pljg81cslr7Gk0iS9yL8q0qO1ItibXlfI7sOsJi8M6WP
uDLQy8G8pkNEtaIM79sEFvDZNcNUB8I8NOBg/BZj4k/fDS0WxTQGeadyP6Fkj2x8
LLfV7je0zMiE7QAJ9fQldMdwtn+2MdlNyw5F2g4rXO4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 33787     )
XnuZ9KaYsjhK6E7TOcNVUVDg0SjogZIwHnSw4iRxQHelYUmf7cpXo2l4zvYHFEtv
CQW2BxstBTUbXA/IPl+2W/QnVnc9ccrDhjB88eooYLpIGaIXOnT1BCgEq2gBIVV3
BMGAsBZ4s+kkfjhiqUkZqFYMoSbaYU1JLWajZAG+uumLvJmdj4DUv6cI4Rut2SY+
32JemuXd3258Ilr7iQm9l2+MuZR8QsUtxqzICsJM0BSDeTL5t/knzXSvTSq/lNGq
2V2wzzC5KjZ20pEb0YyDiEgR5e6ly+nkj1enlYIehU2yn/WK9ktzG6IsjM5l7IgY
XA550fshIpIbR/CAMmr2uTwy11XHLyeWfvZ7Ax0hn7TJt/31mXMycp83cVqugy4E
aGhyPSrCO1W5cnIz+mbrKuLoJdw+ioeUs9wgyg7hyan3F/4qz5uvndHaNj8L+KV7
qm2EwNn5dH+xIPZwt4IQIJj0ojUgJzPjNI0JG4oW6OVwPij8NkAO40MG2JVRMmnY
C7uV9aNkmELEPVYYBnUZStoc6ZRAduk9N9Y3LRJcsZpkjdOrTExr+c+pCTXgwSRF
bCpZKOCBf1Qjg5R+MGIeU0j6NL6nL8La1vJGoq1GyIZzyt6xlOzaWK4219+JxAwv
BTSWUxHBSCF4zVr2enhqcCl+8e61uqZtahkIW3tkS5OYYNBJnMroscQiFYBs8JuR
4UNSrt6IpC61MyqcQrbpk65r0m3knXYjds49PsCX+RX218Srm/3NxL+YgSZoPjcl
WXYp944tG04xjuI6Scjle5r26scse1SswfqRmNLSDb5MqERYYN0MvOosskPJcvts
RZ6voFT+mLXAkRwblGcUayJln71OdiB2zJFLEfu4WlaKqUY520lpsh4jpOyW6iEz
o7WSagW9/gkV7+KeWQ2gcWMORc+kvldm1ips1oZ1QcJ+UDvH4eHrpfxrxdXajZoI
Lqx4nM9mqmdrtEh2m0MiuSDPe0eWkQzUHxqqJUcDDQ8ZrNQ1MGBFkPjbcxGn0qyy
7mzNnzMaAbNSSJuGAmH86oOaTKtvmGkWT8goUU4fpVxazMTG5OBWEtNa4RzFSv0C
BoAtYkFeH6bXmYjPYmEdl3kzC9D0N0m15fSwjXfN1nnQkr8o3Imwd3ApkUx0N1Lr
bs8Iab2apQWqWG5ZXM9huGx3PJ1H3Hs/MQzZgBbIHE++93CVqulQJavqXA6BBMA+
pCFFFZ78xqpHOwGRcOz0nWCqG9HcGFkgrxQox6HZwSgBLytX4KylIwjAkzI/7ZFZ
06nWjASWhr+eTJzcK9fhV4W5eSyL5IFr0ixwN/aP6NdE1nFM0pd36ZaL5KlrAAUx
9DlM7Hpy5ydkqvUgC75bY+eO7Ccr8YgOHlTk7k1YujOIVAx92+zq3TJ6/LibUf8E
Qxv3pqkjLTTMuq0q2mfUFYViNk4HUtwrCtsO1eOPeq9u5BMOrp4bMBlEgBbGwvO1
p1n0IksHu7FC/WbC7XS/1jCFQSc2GE+/PEHWRgXww31fKKCefwP65Rf8mCqVsXex
vYqmN4TeZnJzUpVFPApf9ze0ULcxd/h0XQkqXSimIhVLjpNi0X6RorXTjY9qWykA
fxyrfHR/gcJGcQOo6Js5X6+4umk+CaGiKkjnQtDW5l7oUPq9vCxFSElzvk0BIb+I
C+ImIWj/Cfg3QfuFSRJABAHl0WefRVvvAIBTSsEnKsN0wlbqZBhGGQfY/exfBvUQ
q5n70qWwPfInbbH3irYzp99yPBukoNBBETNPYeNLjsJNUfkKUQYZGLIfomJG/5/P
LmONrVKuqZ/GdX6c+FbGLz6kGRHrKsreR1V8ULVbIcinV6A8OpfVNyom1GugUh++
IR4aBx749bVQ6+meYWq+ZgbgBKBTuVbvJt07ibxvACGzgLG9xspnBlPnmFlFJnev
ImG1pZ7edhMBRIzh8PE+YALHXX1k+imX4H0NRn81LOPrP3qb74awNkSU35+Qrjzf
514Xf5JAiG37fEsH1PFKyBxSKCWR0Xo2H1FwuREvsEuAcVAV+mTYCBJNWnkHovMY
bJYDoZrZg8bxTt2WTrroj87O64ngAPEwdU+O/uU9oJyk5+T0NYIBhyd9fnDkCUgS
pSOwsWo0OFHI65jI/S74U+Jm2IWaaaOzM2eL5vjqZqwzEAZY7FqvEvXwU6/Tlf3L
HkJiqR8GdbCUfa4dxttA6uzhOES+5N1TFvjfWv0DTYU+TTUjDWlW6rUOC9E1QHlX
JSUDkwLPMYSO5YpNHrskMNgKoOzkZJSNCro3BZsYgFI/7s4V+DFw4lsGTBBZmAU8
u6L0XZ+TmianbZOLWp9JPx/1QwMPr9bHNIlgzPzy/SA9f1hWLB5OoHVbfFPJQA3b
t4d4r+X93SLsMiC724roI0xyNY0Td4OZ7wLBtjdr2ok+j1vWlHNwoaSKDO4Y6F/a
jpV0bfVJ6GwR+HA+3dWfHabWpGeCcMI8xP/fGNx/hJlLWY+1ovBDM62TAjE0Aydr
2rlLGHbYYNHrwCt4sIxRUeQRSu+Z2iTpezExToZ1iTyA1AWHps3ZMAkgcIhvCZm9
eZGIUxaanM5AA4b5FK7ATTmUnEtx91cuqzvmT2aDIPMKTrrNmwerWq50adC6aLWE
hpwflIzmoCPjx4HDrs5TeTaPDEvvqZaPUDBAWr5XCjTkd82vMb4NHMsg3CeP9GsY
rI4t7t73iqO64i+tnGN9vZ9cquDe5QDHPjPjxR5TBS9BwiphWI/DH2IgF0VazlwX
pGwDvCbVOPEJnYzZrvLZA/WGquE/6HCsZS7CkXakPqZud+p5mxivj87SwhqeYdRE
/x2Q7dJn5vt/6wLwkAF4KYqQRLsZ0R0bnYQpl/unVGEQrmcKcay9/jWM46IwAaqs
U6WwZsuo0q/NcwlOSmcK+z/SA3bHBNUlbvcoxmtFOSDR74MIMsdZTx4cq7PwOVdu
hfK6TEIssz5q13AJg+8YNTehSSfi5ssF+MB+xKV4K06lEDyl73hnWKXP5JwZCqOT
hXBGK9DJ0IfuT/Fg9Djg/CISWAfRfcVMFOQj5fjuf8P3iB8/eRTzndXRzBgKwkfd
+NCNjZnwC/DMdvgtVzTum86QWcetdarUhjENMIoElaXAoN/vMgG8IT2t4L2aR/ww
VtS16R2wcHyYKtHowEuhfrAP+Jxpl/n5NiupN6f8oP1/ybDVhXubh/IsfEnVKSxD
pDagWhRV+dkR5UC/cypkYdlPUN5Kbkc9Vao/fefKmDyaKAiJBD5dznVkVeLayDue
TNO0qW9Q8jxSwPr64+cBiCVUsHe6Ft59AiTMPWjOurBqERJrxJuUsU4LYSpWfwvL
SzkrUFwANOv2SpIbR5OcY1k0rEM4UpTWu+rSUx7Pdn+fXQALh1RbX3jKt0o296wK
QhDcYrSJFpNJuyCeqHwDr2s0v8GfR30k85G1/dTLcXZe5Etjb1QZK2euL/wGR+Oh
iPi3qN4ip8VC38bsoR+lFqKzmmADlqn23kX4dn57bETVpCVTviqqQxcHW95BG7dZ
E0GxaM7cqBniVri8DZSp4Jf/laLMsnBlhbkzOTtfXCXPhdk6Phg0XOAkBpeulfEd
thq32N+JLtODIRdcN0qYNwOH1GpRzq6PhdTvIE5PQVCtR00dZVLI2bIfPAVLqis5
D7oBTipSMPMtSg2zAdl3n9337Ehm6y+erQXTVqWYB6d+LVW0SNtAlKj19WumzDtP
XUZVUb44G56p5HoIVE8X9HsWn5N3f9azfUQbNrutWLUtePGjzHphXE8bLbKbXFTN
X9pjsl1P1cKDudJW1evSNW2ExNI0bCLjp/XxUqZlmXnXvhkcLTwfPosYoCf4juGT
ktU535KJvVmUJY9ky7ZutXZBYZxrmVZ8T1b5uBVwzLxeMJlqgsmGuipWrurc0C7j
po/4TakUpUe/qoEYfG5REUfiMczAlERuY8F5NRFW0qp9oPxtWmuNNVWLPegHVM9K
+VWAhLO79ci5EcSbp9wxFW1JJPUVLA/+Go6MsTeTBQeWdH2s4ZYhmAOUCDn84VCo
2CKLCzBrdUne+RjcBIzkzuEaI3/hCLE0Qg27IWz7aSpEHx218ic5nzLg7TUAM4CP
daBiNI39Fc0LG8kasRIiRv+qPaom0cs4Y4TAC3wE5dUqDkvl59JSeNmEEoQlRkaQ
5ApB6OlVcQs6XC4qGu8hCNBlY2TtrP2nkfothfeDXGGRYxtRnhEd4RmbzWzX2Pg0
Q8/Ao11OjnGLQPhdVZnvygSDZcX4wcXNEN3RPeJ6lgbAGh7NeTIbsnKbE35qGhGQ
/1fLjhT7cxObplijold8w4im/Ut0ArYILxZP4legLbl/nu3NZFvcQ6J25trgnBDA
xrM7uiYtrGp0FwwJFM0/ePntRiL3T5ZEkb2B8ZCYjl+w2USukuIxhuolpzE/zopM
znWPXM9VSO2SaaPiSky71JoJZnE1RzptL0KyRXL6kTWMayo6/9+BFWrnBxAtlTRZ
sr1eCiymZO25VXVOAU8T2uF0hZ+CgOof33U0uiuLwKv7MT2FiBmSb0qiNEAXzuQh
XBT3xKS6HgDqsrF8EbhdBquLRl7AqmDoC8RDyX86+JPPOFr4NSf5mkBGR18p4Wbc
mBi11dsiE0hZWjPVmv37kgPEfZObBYSg8EYXed1BufwySs22P4G/1VRaP53Jxdip
ImOM1Sl/23Y2x/7lb5fjckik5NFVnSDswaZDEsTXnAJwymGABcW3g7kP20dmDwpr
6womnSa2Afw2X0Yrul7st8GNBBL88oixujKDuAykKdSswRpugrhEeYAI06CgWeD1
ehsoQj8yL+AT9nNR66SyV77iS4Q5BYtmHwBxnhWmal4+JU0eQBt8tLmKuXSxO1cz
fxnlKJNfzuyWxmrSxV/IaeuLnMWCoqFZkQaHfM23/SCliSblAqgzFZ4YTxQw5wFu
4EXWrKUzjrJZtL3UgB8nouG9x2eZN5bdTJ2lytwT8e8KJLqV4F1rxdishQZYPzxf
pEmz5IxFKrzWxS6qELfiyQFQyDd661DqZV+RUErRMyomIhT+BaeJXj1peIVMijSv
frQrAixubieauUkdCpy45pO6quxtn9FeNBml8h0jPsb3o+7sqzp9MbjMgw8W4mdP
uBJD1anLlQ6CK0Zs38+hOY4ToQr2tvh5ISkJzFmDNoIr74+pWT8IBfddIcCG2ShS
UGwJdETrmqGJe3lbkTti7jg5Ogz+Kg9k8NZS5DomSh7C1ODZYN5eugvZIKcU5KmA
8DK+j4jtvwJswEdLP1B6wb7zvgG4i2kYpcj1efu10fC672PhH1pYEwk/NCC9WpNo
5kcmd722IneRhhmLtfOArc+CMBRN4zGwupkcMQ4wlefXfjSQyio9SO3IKWWdFcF5
dgC2IbwZ6GMfrJMRyrtOMkbM9qennwZkfI9LKwM7VXC2SIiPwms//DWe/NoGDMuq
zzMN5GaRig6hEGYPRH7qeapmT/aAPqf+hgbGNCJdJ3ExEjjDcsIhB3T7jvE/qzVR
a0ek7umlAV3xSRLtvJSoxFDIEmaChUAMJWpp/FVItAzYDaduAWC0mg7nyrnX72Qm
o+xu1Z/e3WigpUy7118AEC63wXJTXJ4tXcq+Tu+ocoJq2JQoj3covCYJVb2gCa3Q
Ujlax3dt+7yzGwNX+Kc6VX8GPu/LRK1ikWIENYgXHMWb7ORXXmasYel0cICvCTEZ
im8erwfMmvoYP0BVSOvAEM44o+EXlefy8D0rf5Sn1izmgA0Kjv2fzZWpHUnRJDxT
c6aT4h4zTWycVT5Qd3MG4tjXYAxHrSezydpnY5sx+EqwlHjW5fqs7Oyf6l1AAFCH
WuT7ex+IbPt0OCuxRUlghD7Q0wBwMsOfsUiQ2IDil2myMfiCkdVxIYnIadh90OZ0
AS+d42CjQBy0wMroqdAQgH1PBkPEHulG9vXy56kbqPLh5upiCr0ai+zKXTKnpoYL
qNZd/vgQSQqcIBt58purFiNnG3cQr5xA7L+0IVfCOD5dZftXUPlYarrA5DcyUlD0
QfVtEeZIzQRgp/Ah+afu+VP/CoY8aE1scU+p0Um2uJ/qfRI0FVvX3yWMDtPXouz7
m4t2RWtZjm5S/d+ONjR4N2cNlGJSnYBYn3W9xCsIN/nPs2A9/xK/VIK+Woh8P36p
yLX5rcwb5rTcIalaclL2+vyN7XisqCGamjTO/t3tPuh7DekOWYZDGcO2PglJRPkk
Jqgq/mHBUzH/sAu0EXW04M6ltdjTQfymF6UEcuxsQgc1Ft+tQC1Gb4l53/EORBNc
FpQAuf/k8jms0LV/NpJsnt/9ArWR5s0Aej1BljgfBGuEoUE/9k4s9OFcgvs+J4sn
GzR4E24A9A9KUvrYkYNEBZH3qQJl6b6brkLWr3E4gJYNBLFgMiCAfFomVDqRh4f3
MhrbObrW2q4q/JgQAcFzgP20tvrhZG6bZkD5FaR8GeQLngq8JXHdeOCea92L5C//
abq3NvcoLfgBLG24iUzBowTD7uTfTFIgL31y24Aug2yGgfXIkIH3fnHGp+p2i1Hi
fBzA9QOzF79ZQJbLS89rg8Dqpqaoj+8/AhC2/mMxAkfK+hmPQI8gEoNmjqM9qB3L
rzOxQHZUY7r7K66fE5KMkOqJFfuNxxPlxKdy/bFQim4VH13Mkr2qr5ltGM9Vb508
+nraOrMVcIdqwNkl65xKf9JC/xCcx7rCyKcL8jBBsm2fqWJttLk7MlDxlbl+p2oH
CKn5XgxviVLr5bn15iXrBiGrcRQZxxZxXH1eAh6EeYBLHNAuFYDpn4PyOvPTwzvg
rF+L0sGyLvrgF+0u4n1ANoa+T8oUCOgBQmeUFbVkka/2oCH12PP8SMwr5kLOe7wm
n2N9vi/equBYSfINVgDw/y0f83fyD1QINJgcJtbUuGEhwkRN+JVaW5M2tqN8HJd+
22ZcS5D16+2BklDN69LbIdwNPAC52rOboXS+MP036q4CPI4fy6mhfQ246DvvWdNG
QKU0zyAtG7T0eiGYaPfC4vWJSHhlySlXjre57EWBBqOPf1CStHnzxTIWIX2QjfLW
Is2f519Ce47k429V0DoPqIm7bV/w2Umg2mYhlpEtH/S+yxcbKbIp3I7zf50HzKVx
5mAP5exc5Dd/PxKo1bQmm36BWsUmnDT0wT9OpJxcCn1bTyPp2ufgSwXOqyRet/lL
QYtboYCLizwEdLfXFA7YQxJGrt6IQkGmWw+wcX7C+hV0kcAneYPPi40v+3K+aKRF
zzricQLJjsZzC0j9g4CjSXAgcyM/x9DYqJwM8FOToT0KhvAu0qiKNULOULX0KNJ2
VLcuAuZOMBysLgtEN31dDSjrhDL06bSIDAVMHZhBBnSTB/6zl+8Hf+pf0pqcMFCQ
21PxKidR4Dv3DgD/p5qLmYx5ZIE8TF2gS1XEI5llRG0mzCES5GW+JU8GOlnHrmsP
PMUIT9r0dIRx2bcxeyPl4bkZdmhEaTcyq71l8CYg6qHNHNrFPpskr14IaW8hkkwl
gqmDqocVVvdYibT5oYUDu2KDuHnjLm2SgdLeuX+alEPdV60nwfbkbOUO2lsazI8w
ZsxepmztKpiXprF9Zuoc+oh0h3o88Dlk/NrV6I5LJ4NX3t1tukiMBRzewX5fP8Na
ucOOHvxWdHeNCulaQJB5njhOPJgUUrNXoYEmSYUzhFdZLvgQ3s4QvN5MfXlv/65o
vdauhHaGmFCPXbpbZrtcCfjC3cZJOMtDOU2TXmyUb+jxLH/X/aMc0z7f9YdLdWvk
lgvB3S6FTXnwjCJDZei7Lw2N+YYFkMPugjuFV9uAPnZcPS4jVF3NWlRU+pIPjaYT
pJxkm403/3ClwGvZI06AJIdHYd6CKLIXfY83xfFIH3TPJRdbsgAfGqfm6d68XDFQ
YRvxYgvQvFdnuO22KOXIQVCwzF80Ltg3uUtJMTVu+l5nGBTa8878ZnhuiBCzxU36
zlmEjlY1FBglnxzSnCFTWtG3wsKu8FLWNWDTpqliahRnN7tlO4vm+gSYjJXnjELU
bJFcnRww/LHb91laNF8v5bETbCK1zPGqx+MhoANugiZoUqj6i/jRynjvq2sRvOPo
bGlRYRs+GvW/Y5iMYMTvyuAeE8w4Q4d6tp9VoWiGevI9tbxoWSQysfo1IondZdmh
zy9HzXpsNiEfr6bLr8Y/W+dPUfJe8FMF6D/n490f3QeWM2Yx19My39XaJLgQOKBs
1hHpZ4D88zrdQn5AKmJqj85KUBW46m5ZX7dQH4SpVB8aIOk4fQ+65zNgoTz7iSvy
UpEvrgyC3f9p2uX3ZmbSq2fmjxU6/P2ufibfjLs/gr+QXP+IlpHKokCsmxPh2YKm
LDkjvK2F8LRAw5fd+b/NOVLa231SxwY3LMlOeXMXeFg+s7Q7dGHvjmVGd5hkBNIT
pps67G5KzByqt/w1argbF9ZvBjGM1zjH09f+TiWIuQ4ulTzv6L4e9TxVdq3T+799
YvPXchhdZ4FUs7Mb2qHXXCb15OUrSV6uLQ/RZ9LFNorIYc1PlLjsYMITGe6QW2+Q
ZDJLkVzBQWWb9VollaKrxonYAfzU4q845H6KVuE0TaymDXOrDiK+N+LSG/WodB1+
cUxHjOrVYhEf5agS6Jljw2tAG8CwPIc3OGSDp3+bX1fEavRKjE+E1I0/YK9p+Ck9
rtlxfchKZBl9SzR11GJ4pzc1lv7LUaum7FSLmtxErgOmdD9rcfxgvG2v8I+dsJWN
yZ1ZhIa5eKOTv2NqQZCYFtw/bp/JTyaUvakNAVJWhTQRNYY0dLPeXiskNi2x0rwO
EsI0o0MCfVv/8PoTsUndR5V50WeQLFpQt1Gzy5EcAtBunHQkfvYN1VPNHb9BfPGn
1mW02yaDq/SFG1/Sbb4trW4b8Rp7gRGMl40Ue5sgCJRsRNcAPFRKZgamosj6Av4U
bbxcHMQXuGwQJX37eHMu79LwUW62y/GqXDLlL6Szlf5AIANqi/9sStQ/LAm2q8/F
8jpiA0NRLey0wtH4w/vSS8Z6ZcXAq4ALIVWD1+c54G2Kg3lp0hc7tTBuOPVAGhSd
Bh/kgcd7GU6TfY7VxFzCsrrUVoHFg0d0TQZAWnd2lWQ+h8fKL2azFM5KFmV3/GDs
DDeDYulKATn8CzlHrkukhvGsewvc4EK2cRVV/13Xd/gsN0OhUQFH6jxrWj03DHZJ
NdPS6wiGUN/HdcOJ05No9Oc0FVsIDH1sTaON0n57RJZFWnw1bF/BnDEUlYcS4/FB
kbkd96tBKJFnIyqpLS7iCLvbtQGgnOJ3xtQyTJ4XuUkNcyb4+cKyBwopJAs84Fd/
zAM1A2WbHPF7vBd1sij6QqeHs0lI11dMgZdsEKSIupjIcOyiMmMCzvzpv7M0uoBq
lu/2Ebtz0sb6Vdk3emy+hA596swW3zvEe2Fyl1Y5AOzEYZ6CC0ujbP4qI//Ml+z9
W0qhYy6895UbBU7QPK1Digz2gQW6clioC7bfYvjpaznT8SaUF3Fsy9nerwM5VlM9
5Eu4u6AjWWWLvL3px/GbbwQPT/obAk5pPVSZEmMzEFmRYqMgY5X04Tfly86Z2zDV
xeuKvm6LEJ7CXrcY1SLm21JmxlqO1bdt7OGD94N47IPUGTz5ZZuopOriI7Yk4q5K
CsULfeBxW/nnfTFAFPyXEdsWTaHrsCR59bnkl2/3Dy0t5OJGdZFWRXx7fvTcXT10
xvvSaf9Q99Y8Hz3ADXWU9mjGyUHBbqlllMbCZRy5Q7gMT0cmK/3ZqvZkYbw2b5pY
rcD3p8PTbeK2N3tEIcFwC2lmgao9yPBZ7tCVXiBZ1awSmmeK5MhoWDeTtHXQpgrg
Z+aTAa9jyiL56QmbYUih4u9rAA3h6L2xfREXIP1dL/YDlLWxIYA2ovGMVt15hKXu
S49yxvL3Y2Pq/9gMt2E7aeUyNr7vD337b1MQIMi8fSKD8pVy6cGCrzDsGmFKJ9au
I6ut1MUWE1GNI1d0kLNJIlrO7WJpIemHPyFlmbtoSQsNNW1sSSnT78shCfkZzSRd
nsQeQZqGLGOJuo1Ew1s3ugmjl2zU6omZN5qhcE6vVuSGYglhucg1AhYs7hQXXEpk
LZS68FC/8NT5l8cu+obfNGm2bL4vCBPm3jnTpcZn+hKzKrVK1cQr3+poO4Hdbz3G
G1aUEFBLC4zni4iBXFl1zo4ffcw61WUPBez0fcu/BYOX/TVPahPBnS5yEY2t2gFH
Vonhy098eCp+I0BWLlb2G1n4PIcYlwgYWEfsHf4/YApiual9CKehTd1JTW5mRjrg
SbGjuTzkjW/VgZXYSV2x0hXlHiik8upHctYOLJ7IjWjw+y1plwp3ZD9uP4JnsTnu
jSX6t5NaKy1d/aUDKef71b9tl2cVmH3g7UCNL//T3TSqQ6cCo0G3vfkMCOF6brGP
CeS0mdp2s4sNavpztjp4auzl86KdZw04UqXuxp2PZOvb0cy2MRBdSkl3Nqiy33Ky
IH42SJ/Js7H2kLDPX3o/ClXZ+fcL3Kga7ceH5ZO+CxXuOWL0XQt8kxowITPhB+hM
3QKsoaG6Fs06T4e+RTnhiUc82/XzgK0gdVq9QNIyUBJPBbL1NQIFwNzNWq6a0+NF
6UhXhvfYvyn/YbeMXH/Tx8zRJWHtyKG1f5MiCbUsn9NY9/RozhIKOL9iulWqc4AW
0hzfglp5Bdp8uOJB3Agw8uj+63jgoSjZhCn7VC599mC27iP2BZyDU73ASQNOkXgD
uhov2yjIqkuPVKp2EcWJ8+R9wsp2g6XJXctddOgLr0qp9BuwK4j8BtWv5krxlLqq
pJ6XJqVc9jTybPemYcuwvDL4zY60eq2FaYIRGVk8lLQ0gsjRci/2xMJeS2wfy+lH
MUaVPc9j++BzuMgMKrLTXRttwb1tpePMIMKhI40zfMaOqqx1EJ+o3FTEhKkxgw4m
jKlbf75rGbGCZOxWiwS54S0UrpaJ/Z4CPrqD+HoRGfxexOvR0Kv84HJX+lWu+roZ
LI/TrPbQoBIBjd6OoxPby4/DC2hbPOgBNNbn3OIdA5JOPyqZBZnZlkbVIfi5XuTN
Q7lrgYXIeYtzowOPNthz7rgEeUn534SNkEVNYoEDi34hejZMbXHzHaZ+kSvrp1mY
285YrJKwbZZ9ybY4odvJdDCMIr/DIKPmqJWbIn9Biqc9b3Ytgzo1er8F10owzvSl
MMih4/IekODuhyt9nmTVJYkZFdDNf1j+GA/XXE6CbiC1VbypohjKJHbW6imf/vxd
5fkNvKo/MeeSdEwYWOrPvFdi95fDUafWc4yw8cASXGsdHfK+tqsvXEw24RJXG7mS
Unnrr9Tpn4JZH3ydTal2KNkL225DdN6xVbEsPBCsGWidvJjqiKMjpBovf3PmdE3i
SDEU0netuz1b5hTPUzmO0SYropVa2fGImwMzCHp4c1QUJQfl69CwfsmoQZbmEJjF
t4XDY1sbLxm/AI/O4Jq7M8Cg3u/9TlFAOon3KkwNnuG+kfvzx0GHXRychDknHiRj
ATeScTzamleZPQN8S3DDzKWi0L5scKTg5+DULwcx5ruUeIAC+mXhZXgw9wN6U8rS
mfHaBWBOue8KEat7hVSeBVoiXIfxoZGcP2CIgvs3b1aqVpMSD9gaQRBX5i3VDvnR
ThfKlUohdLkCqMcnxPK2p5ak9khrcWBlkI5NFe4WzTxGYX4XkF5majtcXufMjBGP
Xkt2oKDwLHpI50iwog4bU5wJh5PNiqlVIIQGbX3rmMod5Sa/2jFjXeyYA1XzaA86
NqMEGz+oHtJIwyV8hvHJ8Bw8dafvm0FYLta99PPfUmr/KVAt5uVbq9me4i9EIG5i
CgeSlF4uf27Q56eD8a/yF3Kx68mEGz0I3VsP6NWezTaEoZYfXO6qkstM1HIbSEWH
9a0y5g21zIBcBYXoN8E/wEp+go7vGMcq0YjODLoamLFYqA+Inq8vqv9AFu6JJ5Us
xHPQf7E3tvZ4k8T+bWGubSeMz2dc3tH/6jDPELyyTAKFMJHKe0oquh6t1jy95L2I
VCITSbzdzExqqLUYjKw/45rk/EWTTuIWbpduKxNPmSpi3PJWE6lUfnCezbyhebb6
MDKtVESOPf2pW8aYVIOKsPC/jnHZt8uKRs5y8bbHsaEU+wQb7ZbGHNh6zXvapHRX
hiJdbUwWXS4VNQWXF0k5sf+xOB7L9T1N5eOVQ23WU9BT67dY0CrggUpVSi7N8175
UMaKyl7EVBhGYIaLplEecHTK9or8jPtyDLwuFrJ1dLy5cwqg8wmXmNDnLSE539dW
Eq6cfeaQhZu1WaeWDmC5k6Q4b9MKHZ2f4oVk8jas3uQ6Ds5eUTsX8NJJsPUQN1yC
gDmTMsDC0p5aISuXA8JXly54pWIuhshdXdl3yQyYlqwZ+L79tjTJHZIDJO71eCMP
vS1lhd0GX6y4ZAnDS84X2FXmtz5BsUqdf5g9BZjrI0Tph8gUqQgItv2EYMous99k
I2Af8c8Jwwm3QKEYw08QNcJOfNZoLUZQKX3nFoL3gts=
`pragma protect end_protected

`endif // GUARD_SVT_AHB_CHECKER_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
HKKWf3RZ3eNVfCGoPBLdZPmh2oy4MGQj98rPO7BIQ99hxSaz5kuzfF/x1fFjRi35
nnVGPNsf7T8e4lJrWUK6Ax9A9pWUk18NBmcuR2VNqWSKyf9ndMn0DMNl+bEV1XpZ
mhfzoFIAC4y/6y3bh7xGXIIN3NpDejoo0rQZFJq9TBc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 33870     )
N7YbNlfLst60p5qqHtnvQni8x+SUNqGuYOmxt75SbHee1ICEUVFlERZgRjXYzlih
R2tzVDbG1hHm8fQ/NHLhAmuvyyZzdEzt4ysWNIAaYeGn8agk4OZxMwPTVfByCuQK
`pragma protect end_protected
