`ifndef GUARD_SVT_AXI_SYSTEM_MONITOR_COMMON_SV
`define GUARD_SVT_AXI_SYSTEM_MONITOR_COMMON_SV

`protected
V()EFd=IdZ_KdQRBR-T0972B82FKbPT#TD&?aa@cceI(YC3@FS[,-)>Q6<B<&CQF
U-VNQY2]+H+MC5W3^)6f)2I1#^B-NN=8[Mdg>)P)_4V(E$
`endprotected
`include "svt_event_util.svi"
`protected
EFLV_WI/,H=P=MX(DHTNW(?2#?W_B>Q4+fdM^:>6=X9R-eI4UVM:))<(FaZTVGY,
RLO[Ae+KdWaP0$
`endprotected
`include "svt_axi_defines.svi"
`protected
)CT@D3/EbfV?S7VU0EF#VD0@e^A0A/:CK.35&[Rg1_&)a.W1WD4:4)OZC0+7BgG?
DSX4VEZ61M&@6d&/^Y?P-.c<+PGeS#5=4.,]8=5?F-C&ORgR]-A/dS^&WVO<;G\2
??=\WAT1FD5c<2Q==ZWP0-S/<#A7W/D#XW(a/dE@&)UaX#D2c#N<-QVc4Ce68BE;
0Xe+acE.bX0[R6I\TE,+>@PV=(8bGXe)J-\,@B7;(gF;UN;FTgWPfWHDX(9-#9.<
M@=Ef<TAc#c,R-Y\.gT/E&SDX(=2\]#Q;@M+D>N\:b)FLMT@1>HAb(WQ9BE=Z9YT
e7V85G:WEDDC/Q^/G>Xc>BgUJ2ZFGJe3b_A\ZCO>-;KZB+D?>[R5U(),DW[^)fQ+
8@,-?T^V;3L;6T6-aQMQZ]NdQ045g16O]ZbP.8QLN1V1V_E<a8X,/8>,,:X.1XAf
Z9ZT7+Mac9RK-_>ADd:P.&&ffN08^/AGAX1&BXSY&<QgM/N<aQ=V\,,@R0O2P.F\
fJ&fCBOO&aZ#GeaV.02.,@]cJYZ]d_:<W0GFLE;GPd2BWgb&_6D?[Od?8VV][JD>
,F,X^2g>JIc-XF9^,P7<:_S<PJ=+I(^Q9>Xa5VN72\Z(D07X=M;5;cA6J&fWBX1f
>MC>HcZSY4D/;LQ//(=@>@G1M@#C>1]JYE1VK4D?@K-?aW)YPe/Z39;[+,2UYPXI
He5]ZeRPJ&TCJc(RfRIaQc73L\aGWfAY_L^2+/NVHP5bO#7APg>X;HQ=aO](^THK
cVD>DY.]DD3DJE7YVDcPLY,B^.MSUcLP8)R?6S],@A8b\<45=(OJ(a>(GQMED,:7
FD\@3EJ#@<f:aXW4>5E7W#e:J/;Q(6I?S8>5KIaT,BXNT_RU4bL3?3f/+LF.JdPc
[-Z<dA;PSVI<?APfL_.>N2:)C@\V\?O3\==caPW;Cg4b/<Z#_0HJ>\9(M#TNUK:a
<eV_R>/31Q[9[+RHbU(dF8G;=5.\6]NY1WM@L3d0ADW3#(\E,M<U(@+OfD1K=^G[
T:)7+(94B>H8_3LWd9NPXRFG<e@;;&E65cN?0_b[.4L\bQM=A^ffa+H#B9?DUX66
SB@)L;M,VP(C])/)Ye[9,J^35R+)>N+Z;L+03A;cf@O8U1])JE9RBBM>VcKAF>KQ
(YT:63d2?2(@Ged_W>a]?Q6&B\2E^C\9BTc1^e[2cfPeOP9==BQ<N?eP^&P_3+#.
RY-HLCLc]cBD@,c;3-KPdBT9=?TCU3&,S@#.aPY]Y]RDCO@\P15(CI43RaCbM;JL
:Da_NLS:M1C=6:-I7REOI(58c5<MJ>Y)FT5Mg/WLPRaC7RUHBY#^:e7)MWd1<C]0
IEH7YABTeHO[ZNC)+TD#+LM?LMKO9CaDV<>3,7^:X]9/SXe1S,B&N7)=P.45?9a^
#6I&_d5#^9EQ3:PHY@I70G3(9O=PNX-&RZ>d/<4<-A/P[B+J;(EN><[_BcLT_INI
B4IJ5S?PgR4=:N:VdU85#^@S;^]A.48M.fK9W=4O<8.L\58c#TL9RRGbMK<Od\YK
5NZ73\XAEJT:Mf[#KfgQ[LeAUSQKfKKG\SHHSJUc.DB^f57JS7I.+gMDR/75-A3<
TN4KV?U+YI&6)[)&/D_9^F-cI6dS(.b1<(aKbg)ON5KA4cQ,CM8)-N;+)@;^cTGZ
;U@2b]L59HH#X-gV[UTc.5U-=L@0NRE()2WQ8c+L&C/MPV=H&W&V/,Y]8)NUCX#a
f\6>_,+V?,c_bg&+dZ-^0>JD0EF61)DL_\T=&aDPg\>NbfMfX8GGNSd:X7ZBA7>V
2Qd#HdN)):1X=IO\/N^,7=<1dgUYBf=(FC>H;a3#G@dba+M,V^8K7G53cR\85T).
(c^c=[>)BVa#3,2cVb25:Q;PB0]^J2]ZbKR;ce3JbR_QW\_0]1XTKW1b@_DKKDZ=
]EF)(VS1NYD/GTT65U..@,X^L0MaSG)#:<I_IRPIJ[-GdUEEH,/6G+&YRJRP1+KF
+:.:UVP2N>dEZ,0D/\OR,G>AO>T;2GIAE?a7G<gY>2(M7TLP:-KM)WH9d[+Q>:I6
00U8H_N_V(aP1M-6^F)7.0??OSEccB_>3PU-,M/VR,&b@,4RBd7Ba+FE)AY):+WX
+=071]Mg=c+-b5B7=N+FRV3a_f(RfTR>=8OLLC:RcAeCRBF55TOVD:7D7<BT<eQ7
BW>S?<LJ\QEd65LKf\=S>SSd&XKDP>X@&<D[IY,EQ4:>,C1?adE4FETJ&#^W/GdZ
:Dg&O<;F^d;\L:==[Q)RZJ9;(Je.3]F)(;=@N4[7X(gR(Ke3-DZS+A,3/H[-Vb45
6J9)FWdb#=[Q7\?XC><V)a#S:OWCc<BZ/S1\:N]2YfAK&YB\(c_O1_2JeX..M55A
=#[;DB2bJUZ@bgFfGWefFMR?T[==?:Z.3cCPFJOdd/f-S>.CY&fB.JE-D&S^KfTX
65TP;3\-d?P\F9C6:[F\VCa[XDe2J#P]T#ZaP\#IB24OI:&=Sed16BXFY/M\Uc8A
-61=5c;?PM;2baIb,ZeKIVJY>]5]@\RVg]2<@_T@U.IHOaB?E05=f;@&U4b0:I\?
2VQL9]TA.2]N(#(R)_&NdA^M78H=.?_Pdc.7IdPT.8PRISG\].TLa7V:/07Q+@Q&
FAe)[3<ES[&690g@R<]RdPc>#,ES50gF<=+HIYNHBM2AS#UB7INF;MB@W\;5&UPJ
[GBaY>Fdg;R#1;_N(GeeAK\J)5I@W>Q)6RNFH&YL-90II?aZV)RM=3E7Ug&FZXd;
+<GdSCOPV+&PVP-JRd)Rb_0/Y@b^a^[A/C^QME)e])f8MDKaYH:3GYa7cJ8ITH,?
2S)3_T],K+b3<=Q?/fG-R@0/3$
`endprotected


typedef class svt_axi_system_checker;
typedef class svt_axi_system_monitor;
typedef class svt_axi_system_common;
`ifdef SVT_UVM_TECHNOLOGY
typedef class svt_axi_system_env;
`elsif SVT_OVM_TECHNOLOGY
typedef class svt_axi_system_env;
`else
typedef class svt_axi_system_group;
`endif

 /** @cond PRIVATE */
class svt_axi_system_monitor_common extends svt_axi_system_common;
`protected
d_O?DLb2B<54P/<^].2.;7Z]]]^7f#8](RAa9a@@O87KH3QV&]R=.)5dX&;.41I#
4B@.67_dU[1OW0&UV0]UIX9E=>,_(a4^;>S]=Nc0MV2JJ=fQ4AS6V6OE&;Fe;cP]
S42WU3-LOcO/&ZC76ad9^VIKLU&@-BIGBX]/B:gc>F@XK5;YLGWZD\G<O[^2T#HH
C6@T]UN9Y6(L,Q5.CJd-f4[Y:[T3]g5eO;^bIN8Bcg7NK[Ib.T1SWUcb_a1Z8/,E
aW8UG<K]Z=QN2XMfM-H8Xg=TUKKS?JX@?E/f:\WXfg-YV+a]X3@+gWQ&RfBZ+3(K
LREVC3B]AW#URTE8L;=gV5@+OKbTC,9La]7RPL^JTZ-=])(aP:O9;:6.UDc<EAOF
Tf(B89ZEK@RGMTg0HbK5S=_U\aCTX2@f5:5M@eT>:@+FEbBQ]@e/&d[<SUc(8E+;
C2BQU2^R1+^NcFC=1=_S1Kb?/?WU^,EV9b1dV_)IYe^O=U1-:#+7bcb-R-<cCeML
6I5T7VKe5MV(^1,cMgJ5PL.K//>2]#6VAH\6aP5GCCZ7TW=N\Qe&@T)>#Yc0AH3a
>_B;?YdZG//02&P3(32L)C3Z,/#=;/[]ObV9(YSAY#8_WR:Q)L=9&MM&,BZXX10V
/1YDT?O;\ZYQf;^:E.6&b:[;3)fH.(MN+KZDc5<SV2f_?WgZ,Z(&W,M@IRVI9WN;
(ME0SV(<9NBb]Ge,^Kg_;;dg?+7M)Gcf1QgUF[#5TaO[95T[4#8f&:_N8DV(:e_:
\<bTD.1O(PWMP,W/&<9,O>S52<g9+FSHW3S3a1.aJeOB@FNMC?7@BM6_c<S@(1<_
e7&BU).J/779Z_#WK_&#+K+CB678H9BZX@cg8/4WTE:_aA;0;;;=U38)1c2OQdDc
_1:5W29K#FNFZ)0b36f4VHRdUWd4X3?_MV5=,e7JfRBIZ.8fd5X#<F0.:W,HGAG>
3]B0X8J,NE\PXf.fD8.?^[SB0a#JV2XKZaNJ&Z(4fbJV\348\#fJ)^DaD(9ME\Kf
NK1KUf^\2RWKS#Q3I;Q)S,G^BZAH&.QHD\#[T>A9[>GeO\:Q)dSW9H/Z_[bLL>:&
MG>D)/F&5\.:;80H3&20O3cL19[TBgZ1V3HAP#dT+X-f8W1YC[[dB7.[HK#F:XFg
H1Xc+0T5:SE8E/V&=8Oe-eM&0.fOW9>I34B+(P?A>N#<@E&eG4><YR5G<?SX;K86
Y:VCLI;;>CCO_MHEH0?6H/?&g)1d\YW_B#U9#U3-ASZ&(0TddKW9f^I)+c.#.EK>
L>7WbOgUK-+=SdDTgNE2>54b?>TE#GOOcW+K@6f39]gG)WUWZgIJ.8&)aXb4V5/X
Y>W5_@a14Y=b&\a1SfWV6VLf9,PHIR\^bG,Z.)g\=@C9Z+A\1RFX,-]@BNNXLFRC
e<_C&+KfP1+4QJ3g7(3)VYU;77SZRN6(9acUeHO\1fXT=d)7/daF<O3I\3,H@QY&
FA=fa\OPOT^a,/DXG<ZYSFK+^XfX@LO\<LJJ5a3GXFQBPG\4?.P=O&f:5J&Y>VGa
4eSXa?NV,_]PTV.,M/?]O-Y+41D.717Kf+acDR/2FU@111(1.[@/9:U4B(\.X[N;
3>?0KBB-JN]U>cce&#JgGEYLVDg9HI&IO+&b4LFA.4[ZKR,OdSBHEPO+GbKV#N0X
[S/+>OPKDPI1YAf#O:,R&3;23#Q9<QA]bBg<)H/K8aV-F9\N0+CM:45gY]-<&eTY
8a+-d,YF<Y.(a[-7>1V8d#U.(<Z,:Ng)f#N?9:6Y.CW,>@P,0NQe3LI5E4Ed+R=e
2?3TC^G6c1O\HWe7(-U+61;RdI)c82If2\P9740PSENI1dSXI65/=0@cUc_Sb_Y\
FXQV._?UB&3@PEJbQOTC&PdB,8B-Dc(4ONG^JK[2POTUL<JEEIQTeJZRTW/Rb>?b
13d>=W9\JYbEG]b9,R,e.L-@P:FFIQBc+EJMe,_3]A]K>4YNDPgAYM+@@^A(46+G
GX@a<2>BX:?YL_5C4A2:6O:7N(L648HF2:S;3>Y&L60G)Q2bPUKK<HOaEN_^I^>W
8:&DN+&7YJLb]D)Q>b7V5O8CFaJf3.LC<_,:.^^C&GeJa+IVCXd-XB-9F)U;97SA
653RT2.<5I;]_9VQ5bcII0#J7=,T^&#<RM9g[>.5K7H.VP@+G,SRdE#YcgQBOB1(
NL9S,L\JP&GUM=#AR2Qa-.L(611\RRfbG,JZ7:f;Te7_EQ7e9#FZ@+X004M.+KU9
XS^0]_]:d@0b=(X_a,O=^U)UTdMP\O&7=f)Ca;6b^6UR]T\KUZ3U7EZGM@S[9DRD
2RLZ7?/=\bKAZ\:S.S)>R;dM\&WQ=+927O#LfA//ODAK+e]O@M?H3Rf)YJS_DD6T
a-]L^K2V_dTOFAXG[9NZ9N(8C7K=XJ7,;TNZ@g[IX[a8<+V>O7)_L#R>]UXLZAP3
J/@)[^95M<4_GdBb4GF6PNT]TE1)_]D1F2J>_)<J2N7UGR(ROFA_NY_F@fU2EM7)
(@C0R6gWYIX;N3gd=2NPV.<f+R\<F85)>^_R<.bY.SG9BKD]0#N,5XQ#ZLR.4g&&
>+&HHTZgc2BeK9b0dc3)8dHeJ)e6G=^=AEITJ9d_;NWAGB3X)-DN;F@deX2_MSS#
&NO<H)2,LOMLUKSPIZAFL[72fO@?f7G9G.O:(<CBQL[>Y[<6dRfTd]2_)TW\+YLd
8a+6U5><fN5;F+PgPE9J4&4>XF.O#VFFF9T8YBZH+Wb:/fCH-O>_d+-HRGaBf_@7
L=A#WE1bTP&5WT1_54I\]]eWC(RP15Ac[[U_I3JgI&@Dd717(A^O^/XU0-\PX.CL
HB<XR,#BUMg@IA>c_GUBA]<_7)0=;QC9[@>Xc#M#^bF87W4L=DV;8E#g.7O>+\D4
g@a+g/f:8gEX=G/@P<CJ^^8P?gUBgf[a:F/\5CZV28O?AGP2/42/K9.KJQ65?Y2Q
+a>J+#(WG@c/67L>GOgBbZ@2:ACK=A:#^fJ:ge(Gc[4=M>(Y3_);3Z(_GU^Rbe&a
KE:Q[+#Wb/@g.^B(-e(1EJVGWXa^K,]W9<;\>Ad5GF<KP:8-4;gU-d6_I72,V+=e
(aSD3e>Pe^PPAIfRY:&,F6U]Kb6C)5,XQCA97NaadF@eFT\J/27c\2M<P#0Q\ZO-
Qb/6H8=2c?6QZ_RJU4/]^0&aB>>L,7HS]9.,OAFVYMIDTQddXH@Y:OJZG+;L1E(7
<Ne?[(a9ER/;UO@e12\C-^?aP:;Gfb5b7@MK,C/E(^f^^#\9>,&>;&RHMe6OYU>G
P>KYK6#g#^3f>(YLG:Kd:32A?U]=/2.EVKGG0R-RE)\(D>a8Vebb(0cW8\-[.K)U
f_[-;>g?03D)eA25^DT?><05\A]UW;WG)N2M:d?g^CKY]K#2O5>\cF;MggCd1XNZ
=DN+B5dT#C.+8b/+G25N3WNU&2+a]78X\2FO_IB7(Y9@8f_5&dOQa-,^LVY:;\>Q
76NB3[?<W8(ae7?2][ZJ..W<_\L\V9<HL&2__?YMg/WBA@\1AL=]/\c=T=;[5.WG
S5&EETSZMb4W)/DR(RNd9#?&MSE[[?-LR#9S@C/)805JI0G>Y#\g^9W35IL/b[+_
\R<Oe=E)7FW)BVHJWSI1+-8UP>aTM05#47#;T1S+V?XWSX5Y7.7&UAL2[bCJ)ATJ
3S.==LL90?X7,7?aOg;(_IBN8^QP.ZM#3be<bW=.\9XTJCGU492LSFa&#CQNZ_d/
FJG1a\?fU5^&?=>3KMa7U&5P,]aeSZ_==QM,8:LdNJf#T[#B3Z8&\]/RIT\Vb-+,
-1J2ZGeZaWT,X#CXGO3<9VOgC>R43I6)_/V>3Xe]?6?@eV@OT?POGOG>N([ZS75Q
O8#-+78aM^ERA5.FVAY5bEO5,4RM9J\+]Ig<)Z3IDFVO/1--43/K?cf\@AY0AG<Q
@50ZW,(g0gQ^I097QS)=3C@<S4+#d-0IFDP&g,\(.2AF9CCRbR,B:^?3dT[49)0[
dbC27MC4Ug3N-._VVaV/Nge6&A;7K=RL=^7S?A>HI8Y[SV/,2BX-<K&aAG1&(NU&
G3F?]QC=]N^^-M71GKI=A,UVU]5ZYF]/:^LYPT;\KFL?=JX.\?YM)9G=F,6FQJd.
>Q-RPCc#-B.?C98aV?5JZS86N@+BZ/W/6-+ca&=b=PI?.\JJUBaa?V<-W.=CgA;6
;A=@FfS1LS+D9]e/b1e\C(c8LH#FB(bU>)PJBZ^IP<53cJb&)fg80S65d)TQ9[ZS
8aa5.C=bTd#>@:)1<@e27Y2+dJ=[<&-b#e3PJeP24dbGe.FBgVFH&9Z3g4E:KA)P
L]401HcP3(=NUQSGTHYJ9596/:XP,U@[RKG@6GA;H&0ISJ1QHZHFFS=8P0bPX(f#
-aG67Y4+9R>>?<CdC;Y@/SLTcEYH;fDN50&,OdGI_XcSLW)4RQ&c]_WMUR>KO\K<
ICeM)&8UGSDbZ-_KCY7FBcTfGO=U8/PURg-S(10e,bE8^ZS&?42=a@d<U:I<1_<f
\U[TZ@L4A0O;4=8HUYHVIAI=HNKD4S=If8FIDM(@K0\7f2;QBOF=77Aa2(._)c#+
?_:Q<7(^<G__aFEVE?c\;T;G>J#b?AQO)5-4K3cef,@;-B2E#W4:Sg+ccFFLL)/A
54/+#-bWE5;A<;0d8)7aSXHFP^N-L.G].,0B2L9;HgX5W42M4bD]Oa&81U/HOH[B
5Gg8NLeeQJUaa#4O=3L#C_MGIKB-U<)WY-<U&#8B^GW+958Z.I:Z<;J99UY4fA:6
VI65<(\N1_Oa0$
`endprotected


  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

  //--------------------------------------------------------------------------------

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   *
   * @param reporter UVM report object used for messaging
   * 
   * 
   */
  extern function new (svt_axi_system_configuration cfg, uvm_report_object reporter, svt_axi_system_monitor system_monitor);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   *
   * @param reporter OVM report object used for messaging
   * 
   * 
   */
  extern function new (svt_axi_system_configuration cfg, ovm_report_object reporter, svt_axi_system_monitor system_monitor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param system_monitor A handle to the monitor class of type svt_axi_system_monitor 
   */
  extern function new (svt_axi_system_configuration cfg,svt_axi_system_monitor system_monitor);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Sets up exclusive access monitors */
  extern virtual function void set_exclusive_access_monitors();

  /** Sets the configuration */
  extern function void set_cfg(svt_axi_system_configuration cfg);

  /** Sets internal variables */
  extern function void set_internal_variables();

  /** Adds transaction from master to IC to internal queue */
  extern task add_to_master_xact_active(svt_axi_transaction xact); 

  /** Processes master transactions which must be split for system monitor use due to DUT requirements */
  extern task process_split_master_xacts(svt_axi_transaction xact, svt_axi_transaction split_xacts[$]);

  /** Processes received master transaction */
  extern task process_master_xact(svt_axi_transaction xact);

  /** Adds transactions to the queue. These are from the IC scheduler */
  extern task add_to_master_xact_active_from_ic_scheduler(svt_axi_transaction xact);

  /** Adds transaction from IC to slave to internal queue */
  extern task add_to_slave_xact_active(svt_axi_transaction xact); 

  /** Adds snoop transactions from IC to master to internal queue */
  extern task add_to_snoop_xact_active(svt_axi_snoop_transaction xact); 

  /** Add a barrier transaction to internal queue */
  extern task add_to_barrier_xact_active(svt_axi_transaction xact);

  extern task get_sys_xact(svt_axi_transaction xact,
                           bit delete_post_get,
                           output svt_axi_system_transaction sys_xact);

  // Checks correctness of data for transactions that access multiple cache lines
  extern function void check_cross_cache_line_data_consistency(svt_axi_transaction xact,svt_axi_system_transaction sys_xact,bit[7:0] mem_data[]);

  /**Checks the byte count of writes across masters and slaves */
  extern function void check_master_slave_write_byte_count();

  /** Gets list of system transactions where master xact is not fully mapped to a slave transaction */
  extern function void get_unmapped_system_transactions(output svt_axi_system_transaction unmapped_xacts[$]);

  /** Prints summary of transactions that have not been fully mapped to slave transactions */
  extern function void print_unmapped_xact_summary();

  /** Gets the fully summary report  based on entries in xacts_summary array */
  extern function string get_full_summary_report();
  extern function string get_full_summary_report1();

  /** Reports end-of-simulation summary report, checks etc */
  extern function void report();


`ifndef SVT_AXI_SNOOP_FROM_SLAVE_ENABLE_1
  /** Checks if the snoop transaction's address matches an outstanding coherent transaction */
  extern function bit check_snoop_addr_match(svt_axi_snoop_transaction xact);

  /** Process this transaction and execute relevant checks */
  extern task process_coherent_xact(svt_axi_transaction xact,svt_axi_system_transaction sys_xact);

  // Checks if there were read or write transactions which were started prior to or after xact
  // was started to an overlapping address.
  extern function void check_rd_or_wr_xacts_during_curr_xact(
                                                   svt_axi_system_transaction sys_xact, 
                                                   svt_axi_transaction xact, 
                                                   bit[4:0] overlap_xact_type_check_mode, 
                                                   output bit is_rd_or_wr_xact_before_curr_xact, 
                                                   output bit is_rd_or_wr_xact_after_curr_xact);
 
  // Checks if there were write transactions which were started prior to or after xact
  // was started to an overlapping address.
  extern function void check_write_store_cmo_xacts_during_curr_xact(svt_axi_system_transaction sys_xact, svt_axi_transaction xact, 
                       bit check_store, bit check_cmo,
                       output bit is_write_store_cmo_xact_before_curr_xact, output bit is_write_store_cmo_xact_after_curr_xact);

  // Checks if there was any transaction that overlapped current transaction and completed in different
  // order than it started
  extern function void check_overlapped_xacts_during_curr_xact(svt_axi_system_transaction sys_xact, svt_axi_transaction xact, 
                       output bit is_overlapped_xact_before_curr_xact, output bit is_overlapped_xact_after_curr_xact);

  /** Process barrier transaction and execute relevant checks */
  extern task process_barrier_xact(svt_axi_transaction barrier_pair[$]);

  /** Returns the snoop transactions associated with this coherent transaction */
  extern task associate_snoop_to_coherent(svt_axi_transaction xact, svt_axi_system_transaction sys_xact,
                                          output svt_axi_snoop_transaction associated_snoop_xacts[$]);

  /** Gets the snoop data as a string */
  extern function string get_snoop_data_string(svt_axi_snoop_transaction snoop_xact);

  /** Performs checks on associated snoop transactions */
  extern task perform_associated_snoop_checks(svt_axi_transaction xact,svt_axi_snoop_transaction snoop_xact,svt_axi_system_transaction sys_xact);

  /** Removes a coherent transaction from queue */
  extern task remove_from_master_active(svt_axi_transaction xact,svt_axi_system_transaction sys_xact);

  /** Removes a snoop transaction from queue */
  extern task remove_from_snoop_active(svt_axi_snoop_transaction xact);

  /** Removes a slave transaction from queue */
  //extern task remove_from_slave_queue(svt_axi_transaction xact,svt_axi_system_transaction sys_xact);

  /** Remove a barrier transaction from queue */
  //extern task remove_from_slave_barrier_queue(svt_axi_transaction xact);

  /** Tracks allocations of cache based on snoop transactions */
  extern task update_snoop_filter_after_snoop_xact(svt_axi_snoop_transaction xact);

  /** Indicates if a given transaction generates a snoop or not */
  extern virtual function bit has_snoop(svt_axi_transaction xact, svt_axi_system_transaction sys_xact=null);

  // Check if the snoop generated is one of the valid types for the given coherent transaction
  // Refer Table C6-1 of the AMBA4-beta specification
  extern task check_coherent_and_snoop_type_match(svt_axi_transaction xact, svt_axi_snoop_transaction snoop_xact,svt_axi_system_transaction sys_xact);

  /** Checks if the port on which snoop is received is in the domain indicated by the corresponding coherent transaction */
  extern function void check_coherent_and_snoop_domain_match(svt_axi_transaction xact, svt_axi_snoop_transaction snoop_xact);

  /** Checks that a secure coherent access results in a corresponding secure
   * access in the snoop. Similarly a non secure access results in a
   * corresponding non secure access in the snoop 
   */
  extern function void check_coherent_and_snoop_prot_match(svt_axi_transaction xact, svt_axi_snoop_transaction snoop_xact);

  /* Checks if all conditions are met before starting response to a coherent transaction */
  extern task check_snoop_transaction_issue(svt_axi_system_transaction sys_xact,svt_axi_snoop_transaction assoc_snoop_xacts[$],
                                                     bit was_unique, bit data_transfer,bit pass_dirty,int snooped_ports[$]);

  /* Checks if the is_shared response to a coherent transactions is correct */
  extern function void check_is_shared_response(svt_axi_transaction xact,bit was_unique,bit is_shared,bit is_shared_of_unique_xact,bit data_transfer);

  /* Checks if the pass_dirty response to a coherent transaction is correct */
  extern function void check_pass_dirty_response(svt_axi_transaction xact,bit pass_dirty,output bit is_pass_dirty_error);

  /* Checks if all the caches which have an allocation in the given domain are snooped. */
  extern function void check_all_caches_are_snooped(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, svt_axi_transaction xact, int snooped_ports[$], 
                                                    output bit is_snooped, output int snoop_port_with_cache_line);

  /** Checks for coherency of all cachelines which are clean with memory */
  extern function void check_all_cache_mem_coherency();
  /*
   * Updates snoop filter of a master based on the coherent transaction.
   * Refer Section C10: Optional External Snoop Filtering
   */
  extern function void update_snoop_filter_after_coherent_xact(svt_axi_system_transaction sys_xact);

  /** Data-Integrity:: Checks for coherency of cachelines which are clean for this addr */
  extern function void check_cache_consistency(svt_axi_transaction xact, svt_axi_system_transaction sys_xact);

  /** Returns 1 if all cachelines are clean for this addr, otherwise returns 0 */
  extern function bit get_clean_status_of_all_caches(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);

  /** Data-Integrity:: Checks consistency of cacheline and memory for a particular address */
  extern function void check_mem_cache_consistency_by_addr(int cache_line_size, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, bit[7:0] data[], int master_num, bit is_error, bit is_warning = 1'b1, svt_axi_transaction xact=null);

  /** Data-Integrity:: Checks consistency of snoop data with coherent data */
  extern function void check_coherent_and_snoop_data(svt_axi_transaction xact,svt_axi_system_transaction sys_xact,svt_axi_snoop_transaction associated_snoop_xacts[$]);

  /** Data-Integrity:: Checks if there was a previous writeback/writeclean transaction while a read was initiated. If so the data in the WRITEBACK/WRITECLEAN is expected */
  extern function void check_data_integrity_with_last_coherent_write(svt_axi_system_transaction sys_xact,svt_axi_transaction xact,bit[7:0] coh_resp_data[]);

  /** Gets the system env/system group */
  extern function void get_system_env();


  /** Checks read transaction timing relative to the last posted write transaction */
  extern virtual task check_read_timing_wrt_last_posted_write(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  /** Deletes transactions from sys_xact_assoc_queue */
  extern virtual task delete_from_sys_xact_assoc_queue(svt_axi_system_transaction sys_xact_map_queue[$]);

  /** Checks protocol restrictions for non modifiable transactions */
  extern virtual task check_non_modifiable_transaction_properties(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  /** Prints coherent and associated snoop information */
  extern function string print_coherent_and_snoop_xact(svt_axi_transaction xact,svt_axi_system_transaction sys_xact,svt_axi_snoop_transaction associated_snoop_xacts[$],bit do_not_display=0);

  /** Gets cache contents of address in xact for all masters */
  extern function string get_cache_line_content_string(svt_axi_transaction xact,svt_axi_system_transaction sys_xact);

  /** Adds summary report of transaction to an associative array indexed by the start time */
  extern function void add_xact_summary_report(int start_time, string xact_summary);
 extern function void add_xact_summary_report1(int start_time, string xact_summary1);

  /** Gets memory contents for address in xact */
  //extern function string get_mem_contents_string(svt_axi_transaction xact);
  extern function void get_mem_contents_string(svt_axi_transaction xact,output string mem_contents_string);
  //extern task get_mem_contents_string(svt_axi_transaction xact,output string mem_contents_string);
  // Data-Integrity:: Checks consistency of transaction data with memory data
  extern function bit check_xact_data_consistency_with_mem_data(svt_axi_transaction xact, svt_axi_system_transaction sys_xact);

  /** Gets the associated snoop transactions' data as a byte stream */
  extern virtual function void get_associated_snoop_data_as_byte_stream(svt_axi_transaction xact, svt_axi_system_transaction sys_xact, bit use_dirty_data_only, 
                                             output bit[7:0] snoop_data_as_byte_stream[], output bit is_snoop_has_data[]);

  /** Checks snoop data contents with corresonding bytes of coherent xact. Returns 1 if it matches */
  extern function bit check_snoop_xact_data_with_coherent_xact(svt_axi_snoop_transaction snoop_xact, svt_axi_system_transaction sys_xact, svt_axi_snoop_transaction assoc_snoop_xacts[$]);

  // Gets the memory contents as a byte stream
  extern function bit get_mem_contents_as_byte_stream(svt_axi_transaction xact, output bit[7:0] mem_data[], output int slave_port_id);

  // Processes DVM Operation and DVM Sync
  extern task process_dvm_message(svt_axi_transaction xact,svt_axi_system_transaction sys_xact);

  // Process DVM complete transactions
  extern function void process_dvm_complete(svt_axi_snoop_transaction snoop_xact,output svt_axi_system_transaction dvm_sync_sys_xact);

  // Associated snoop transaction to DVM Operation and DVM Sync transactions
  extern function void associate_snoop_to_dvm(svt_axi_transaction xact, 
                                     svt_axi_system_transaction sys_xact,
                                     bit skip_snoop_association_check, 
                                     output svt_axi_snoop_transaction associated_snoop_xacts[$]);

  // Gets ports that need to be snooped 
  extern function void get_snoop_route_ports(string mode="dvm", svt_axi_transaction xact, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr=0, ref int snoop_route_ports[$]);

  // Prints DVM Complete transaction
  extern task print_dvm_complete_xact(svt_axi_system_transaction sys_xact);

  // Prints DVM Message and corresponding snoop transactions
  extern task print_dvm_message_and_snoop_xact(svt_axi_transaction xact,svt_axi_snoop_transaction associated_snoop_xacts[$]);

  extern function void check_xact_decerr_response(svt_axi_transaction xact);

  /** Checks if there is an ACE-lite transaction to the address given by snoop transaction */
  extern task check_xact_from_ace_lite_to_addr(svt_axi_transaction xact, svt_axi_snoop_transaction snoop_xact, svt_axi_system_transaction input_sys_xact,output svt_axi_system_transaction sys_xact, output bit found_ace_lite_xact_to_same_addr);

  /** 
    * Registers information about association of snoop_xact to xact with the given system transaction 
    */
  extern function void register_snoop_from_ace_lite_info(
                                             svt_axi_transaction xact, 
                                             svt_axi_snoop_transaction snoop_xact, 
                                             svt_axi_system_transaction sys_xact
                       );

  /** Tracks byte count of write transactions from upstream components */
  extern task track_upstream_write_xacts_byte_count(svt_axi_system_transaction sys_xact);

  /** Tracks byte count of write transactions from downstream components */
  extern task track_downstream_write_xacts_byte_count(svt_axi_transaction xact);

  /** Track slave error response */
  extern task track_slave_error_response(svt_axi_transaction slave_xact);

  /** Checks if an error response was received at the slave for any of the addresses
    * corresponding to xact */
  extern task check_slave_error_resp(svt_axi_transaction xact, output bit is_slave_err_resp);

  /** Indicates if this transaction can be correlated to a slave transaction */
  extern function bit is_xact_correlated(svt_axi_transaction xact);

  /** Indicates if there are any full AXI_ACE master ports */
  extern virtual function bit has_ace_ports();

  // Gets a combined read response from all the individual read responses. 
`ifndef __SVDOC__
  extern function void check_read_response_status(svt_axi_transaction xact,output svt_axi_transaction::resp_type_enum rresp);
`endif
`endif

  /** task to start timer to track timeout between coherent transaction and corresponding snoop transaction */
  extern virtual task coherent_xact_to_snoop_timer_start(svt_axi_transaction xact);

  /** task to end timer to track timeout between coherent transaction and corresponding snoop transaction */
  extern virtual task coherent_xact_to_snoop_timer_end(svt_axi_snoop_transaction snoop_xact);

  /** returns 1 if a cacheline is allocated in any of the peer master's cache, if mode is set as "peer"
    * returns 1 if a cacheline is allocated in the master specified in curr_port_id, if mode is set as "self"
    * returns 1 if a cacheline is allocated in any master's cache including initiating master, if mode is set as "all"
    * if current transaction handle is provided "null" then the explicit cacheline address and port id are used instead
    * of transaction address and port id
    */
  extern virtual function bit is_cacheline_in_snoop_filter(svt_axi_transaction curr_xact, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr=0, int curr_port_id=0, string mode="peer"); 

  /** returns 1 if system transaction corresponds to master transaction that attempts to allocate a cacheline and
    *           has at least one overlapped transaction that attempts to de-allocate the same cacheline at the same time.
    *           This check is needed for system monitor to determine whether snoop filter corresponding to the port of current
    *           system transaction should be allocated or not when master sends allocating and de-allocating transactions
    *           at the same time. Please refer AXI-ACE specification IHI0022E C10.2 for further details related to this requirement.
    */
  extern virtual function bit has_overlapped_dealloc_xact(svt_axi_system_transaction sys_xact);

  /** Waits for transaction to be accepted */
  extern virtual task wait_for_transaction_accept(`SVT_TRANSACTION_TYPE xact);

  /** Waits until snoop association can start */
  extern task wait_for_snoop_association_trigger(svt_axi_transaction xact, svt_axi_system_transaction sys_xact);

  /** Executes the master_slave_xact_data_integrity_check */
  extern virtual task execute_master_slave_xact_data_integrity_check(svt_axi_transaction xact, bit is_pass = 1,string desc);

  /** Executes the interconnect_generated_write_xact_to_update_main_memory_check */
  extern virtual function void execute_interconnect_generated_write_xact_to_update_main_memory_check(svt_axi_transaction xact, bit is_pass = 1,string desc);

  /** Checks if CMOs were forwarded to the correct slaves */ 
  extern virtual function void check_cmo_forwarding_to_slaves(svt_axi_system_transaction sys_xact);

  /** Executes the interconnect_generated_dirty_data_write_detected callback */
  extern virtual task interconnect_generated_dirty_data_write_detected_cb_exec(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

  /** Executes the master_xact_fully_associated_to_slave_xacts callback */
  extern virtual task master_xact_fully_associated_to_slave_xacts_cb_exec(svt_axi_system_transaction sys_xact);

  /**
   * Returns the requester name for the supplied master transaction
   * 
   * @param xact Transaction for which to return the requester ID
   * @return The component name that generated the request
   */
  extern virtual function string get_master_xact_requester_name(svt_axi_transaction xact);

  /** Sets the expected snooped ports based on the status of snoop filter and overlapping allocating transactions */
  extern function void set_expected_snoop_ports(svt_axi_transaction xact,svt_axi_system_transaction sys_xact,bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] tagged_addr);

  /**
   * If complex address mapping is enabled, this method translates the supplied master
   * address in the transaction to a global address, and then uses that global address to
   * determine the slave address and active slave port ids.
   * 
   * If complex address mapping is not enabled then the address is converted to a slave
   * address and then the port ids are obtained using the legacy methods.
   * 
   * @param master_addr Master address to be converted (can be tagged or non-tagged)
   * @param system_id AXI System ID
   * @param is_ic_port Determines if the address originated from a port on the interconnect
   * @param xact_type Transaction type (read or write)
   * @param is_tagged_addr Determines if address tags are present within the address
   * @param is_register_addr_space Returns 1 if this address targets the register address
   *   space of a component
   * @param slave_addr Local slave address
   * @param slave_port_ids The slave port to which the given global address is destined
   *   to. In some cases, there can be multiple such slaves. If so, all such slaves must
   *   be present in the queue.
   * @return Returns 1 if a matching slave address was found, otherwise returns 0
   */
  extern virtual function bit get_slave_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] master_addr,
                                             int system_id,
                                             bit is_ic_port,
                                             bit master_port_id,
                                             svt_axi_transaction::xact_type_enum xact_type,
                                             bit is_tagged_addr,
                                             output bit is_register_addr_space,
                                             output bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr,
                                             output int slave_port_ids[$],
                                             input svt_axi_transaction xact);

  extern virtual task check_slave_routing(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact=null);

  /**
    * Checks if there are
    */
  extern task check_overlap_address_secure_and_non_secure_access(svt_axi_system_transaction sys_xact, output bit is_untagged_secure_nonsecure_overlap, output svt_axi_system_transaction overlap_xact);

  extern task update_access_type_info(svt_axi_system_transaction sys_xact);

  extern virtual function void check_mismatched_access_types(svt_axi_system_transaction sys_xact, output bit is_mismatched_access_type);

  /** updates snoop filter size by modifying total_snoop_filter_size variable based on the
    * argument number of modified entries i.e. num_entries
    *
    * @param num_entries indicates how many entries need to be increased or decreased. If
    *                    size needs to be decreased then <->ve number should be provided i.e. if
    * size needs to be decremented then -1 needs to be passed.
    */
  extern virtual function void update_snoop_filter_size(int num_entries);

  /** returns number of entries for the specified address across snoop filter of all the masters.
    * @param addr address for which number of entries in the snoop filter must be searched.
    * @return Returns number of entries 
    */
  extern virtual function int get_num_addr_entry_in_snoop_filter(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);
      
  /** This methos allocates a cacheline into L3 cache inside system monitor and returns '1' if successful else '0' */
  extern virtual function bit l3_allocate(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,
                                          bit [7:0] data[],
                                          bit byteen[],
                                          int is_unique = -1,
                                          int is_clean = -1
                                         );

  /** process current transaction to determine L3 cache allocation or deallocation and perform relevant checks */
  extern virtual task process_l3_cache(svt_axi_transaction xact, svt_axi_system_transaction sys_xact, svt_axi_snoop_transaction associated_snoop_xacts[$]);

  /** Checks restriction that WU/WLU transactions must not be sent when WB/WC/WE transactions are in progress
    * on an interleaved port */
  extern virtual task check_wu_wlu_restrictions_on_interleaved_ports(svt_axi_transaction master_xact);

  /** Invalidates snoop filter for given address */
  extern virtual task invalidate_snoop_filter(bit flush_all, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] tagged_addr=0, svt_axi_snoop_transaction::snoop_xact_type_enum snoop_type=svt_axi_snoop_transaction::CLEANINVALID);

  /** Prints outstanding snoop transaction information */
  extern function void print_outstanding_snoop_debug_info(svt_axi_system_transaction sys_xact);

  /** Checks if outstanding coherent transactions have a snoop or slave transaction associated to it */
  extern function void check_snoop_and_slave_xact_for_outstanding_xacts(svt_axi_system_transaction sys_xact, bit use_error_addr=0, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] error_addr=0);

  /** Checks if the sum of snoops and slave xacts for a set of overlapping transactions is as expected */
  extern function void do_snoop_and_slave_xact_group_check_for_outstanding_xacts(svt_axi_system_transaction sys_xact);

  /** Checks transaction data match with outstanding snoop queue */
  extern function bit check_xact_match_in_outstanding_snoop_queue(svt_axi_system_transaction sys_xact, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] expected_snoop_addr, output svt_axi_snoop_transaction snoop_xact);

  /** Checks transaction data match with slave transactions that overlap in time and address with it */
  extern function bit check_xact_match_in_overlap_slave_xact_queue(svt_axi_system_transaction sys_xact, svt_axi_system_transaction sys_concur_xact, svt_axi_transaction concur_potential_assoc_slave_xacts[$], bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] snoop_addr, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr, output svt_axi_transaction potential_assoc_slave_xacts[$], ref int potential_assoc_slave_xact_count);

  /** Process address and updates relevant fields in system transaction */
  extern task process_and_update_addr_info(svt_axi_transaction xact, svt_axi_system_transaction sys_xact);

  /** Samples Reset signal via axi_if.interconnect_resetn and detects Reset assertion and deassertion */
  extern virtual task sample_reset();
  
  /** Checks if CMOs were forwarded to the correct slaves */ 
  extern virtual function void check_data_integrity_with_outstanding_coherent_write_at_eos();

endclass
/** @endcond */

// -----------------------------------------------------------------------------

// System monitor cannot be supported in the INTERNAL ACE TESTING at port level
// This is done in the tb_ace_vmm_implicit_1m_1s testbench directory and
// the tb_ace_lite_vmm_implicit_1m_1s testbench directory where we mimick the
// behaviour of an interconnect port. However, these task need to be defined
// so that things will compile.
// -----------------------------------------------------------------------------
`protected
3e[^S,\c.P&>NaXU59gC=egP#,)VYU6cVQ855V@V;N1KQ?@-b..]7)C#_<T#5WP#
#UEAUca3Ob#Of&;EeGVF7>FP2]OSEXaa=#YaJ__S:0f8+V5d(64>:.H\#RX(2>,@
]@4I?\d[C@M?a)E>Y\-TD^SN0g:7.9E6JgHdI9Y7ZdV2fX4(G2[dH[,[_0]EB.9C
N.&G)Fe)f;_U0]eGSc9[=<+^6RW)9^BQC[d\g).0BH;Va4B/da448.NgE9B)REH@
6)11K[QC4I(UQ,DeI1JLg<[C=g[SXX53f)DH5DKHdYIeC\O8Mf:G=QTg@(]]I1,,
S36#ES2<;L/V@#?N\UdYK-;AC8KT\INHbbdTgb4TP32[52d[e0F&c.f:4B=P&1bF
aEFTBa15XS.9(H5g\KOQ;P:^.<N/4@+,F8-UcGbg\ERPL?.(J10AZeeSTc#7,5bW
0C03CadDF]96#^c#I>E7J2d69+.(VJ^_3\O<5X;@8J@5QcDZ;BN?bHW>1e1TE&OY
<BWf70#&9@^,E<4[:T(I-9970&5[;#7/_03UeX9;PcD@QbeS+NST5-B:BSMdW]V;
fI0JTf^7^62#+>8-XEH2Td&&VM^c#K_R/8)E@UDFTJbW5:RN6e&L-0UYEU1WNSG9
>JK+L>TER;dLT7YBR]JZU/OVP4R<(ge9-JJJ53:R\@=MP18fNdLe70V:c][Y4XVT
fe,]Acbfg?&&>VDN@Ue:_\0-M9RK4Q(cefd;?=S+S#YDJA5\:;d7bXe_0(2.P8X3
+98U[F&+:+ZH[ebW9/5FWAI87CX5FbP8.:OO8JGc6c[Y)C]A3f39d.WW5TBF@1_B
192@#Ya)DXS3/K@;;6R6.:>XOLF3e[g7VScY2<PH-@\4Ge2\RKZ3UeL]d^JM-5)9
Y)7GA[4cCUb6G/bcH3/dVBg@U+TN>a3]WE>S#DcTUXZ]OVLE1[KNK)BRGGMK+W(H
c;>GM;#f^@a3I?4=4.b1_59He0KVKLI^d,f57T0XIHRET1]1EW?_Q1V9PJ;15CJO
/:E>[RA9A(d_FbZ_^Sf)JJJ?@dV1SWgfL#]]<-:RP=56DOGI0<b1O+K?&[1Sb,7#
E)5O,FU0AT,06KO]-PE29/]IC^7>&fD9HX7(0a5:A:aO2#(?A4bTf_fG,g?fE&::
f,)#8gZO32G1?&#R4aPFQc@OT)(XE;=\a0#3YSCOgfGa)]\WMZcYaJ6V;_-(1/R=
62\a.FI.cEdL.MQ8Y^P-U1S4)VeKV33E0P-f,eXELOD\:eLJd/885Z^^\T)eX1D3
S#27YReYCgP=,/G^H]T:;g^7:I(gWELc6L:<V;d-=5>7-(GGA7aecN/K6P^)_1EP
9Z>2#g\9>T/-HO=K;TJ.M-^e64ID7DG>JC-\<D^28I_K#[.&(/F;2A7F&T#2Q#VW
Q^#CW#Ga9U(;Ebb(,X)aY#+8PA[/<4HYM\BZU^_V&+@\L/[8OOTW3+Z:5e3U1KAP
8[DN/KXJJ=9^_dNd&<H7NNGZ9RI_#XMb5C.BQbE)/697:gP:S\NfgXdA,GWWFV\Z
Ra,AeAZ_766#+5=+?GVQ]O1O,_0G[[+G]US_V)4D:@0/[&7OeM(LG<]W,W3XKR]=
f/01_0=(-Q9T1I5gW0XXD9[:O8\K=D^3PaHa,aR2d\F^9]9KN&]I5_?^NCM_BS;^
H.,[)Fc=-I64G-M(+_I3eL#G7TR7/35P(YK/7FeO&FK05Z]2K93Cfe\BKMfA1N).
B8_1V.Y?gd5U>=UW;L#QUDJTb&H0MJeH6P([B^<]+1?BcSPHd_]BH5?[PY>WaPLW
[Z][EQVX0I05RY<+L-R=3(O\[LK\GU&B<XIbOMd:Y/UC>:4=/EeIN[_]A&N+_W#Q
bTCPPV+c9DQ40?>7V8b=_+K/eK(KA<-If2VY(^;NDc(YK7MZZ#cICGR\-bc0e;.X
X[R9eZ,a2/N7EKR<?^5E>F82E?S8.EY#<I&;6\B&9C04U93X=.<A81L:T5\+H9J(
VGD6NdB]&Ad2Wg-=+LGTB.6M_F?>5e\g14bQ37HA<dHeReQ@7c+-4DeD^Ab>GPG0
<g&32fT-ZFIV;=.Aa=QZEJ&XYd39a#a/:=PHc9dN4-#Z9??8U])afce07--J]RFa
]JfN96I?8=SIFS3bc(96d272-1RIZAb6c0_11/M-WgJY?6,bGQ_eT2.Bfg?3W=[@
A1#^@eYD2<=C;FDgV[a+bdFY/>,-8b[H;_PJEA7[FB]&@1R+T46N9G5C-eLcgE?c
7N9PLB^(a4BNM07;9^?T())1<L9aH=BYA-a:4SA#?7TGQD1&:T?,K^COSL^D<Q_5
@<<:Q.7\Q[8E<dUb[4K()IF,/;)I,Q:VTHPP^)@LU#G?;B@6c<3.?M][OJ]cH\BG
10Hf43.Wc-#DeE;1N/8N:-R[Z3W3-:MeR-]2a\(H>?G]/X-77#AQ0b4>g7VIeC9-
9S(CEcN(T?_FE&LB5YF8YS2EDY,B@BVMZ6YNC-N)I8b\2?9BbN\LcPR/BfRU?b\#
F)&MLgbEV^H:]Zdf2M]=.#X,+WJ:Fa?/+N84I_7d38c-5=WKCH?@TbE9Z2QG=Gb;
8,Ze[+:?ECg^6:TLIUfP\eEGI5.2>#MZ<@&\06/43OBLaSQWe]U]4J75fSg=NZF&
g=29WeU/2&:_=;.YK.(Q2?M;.^;(gVe\GCD)MNVefLOV-aIaPGNO,IgZR?&Tf[M[
g;H/QfGGcf]GfSF@eKDY=@6A^K7d^TIB7NDS.J3U2#\_g9OeKA<+&OUD9MPV4<:O
NJ^Q(<?LXBMWERaZB)VS;,d>T1?5+LUbZ4,f)7TMM_FD&GR5NTCAc&3dZPX+F7#@
<E+;<IKD3TY.QIH]7Rb5)VJ:Y?Q?CFMcUc#9WI\D73F6J89RgI.;^e.cIOV#T5dV
&Y3[OL:D3IU4H[__S8J2#e4O0?0EYgCA).H.V1)QB,JVad)e=.(YQe+WDK?ABW=&
)NeAHT_NgWVTUZ(&8Q/K0F)6G5D\&8Z]8PPId0Hd\Z=@/V\_8?aa5FZ0<5C2B9N,
]UbHbeaTPZ=M5dGP4Ta-8a16V.L(:AM6C4=aYUW:cD7RgO]:5E9J^WS#D2B(.\A.
a?fg/NK\\7H#NGOcMR>RV1:6I;8#P)3K@6dR>]-geB#:c?(X3?Qe;EVEOaKeU6MI
dddVM/19T9HEfHC?R\&+HK1aZgW9TZFEG9QA32?0,D/W8)1d#TJ<0^K6ZRgPZ/Kg
&&.cMRZIE,/9^C5YQ&#-^]5a+@8XQ#=#DD07>@>I:B0a#-+g,Z(MZYDS5KgP^e+f
3=#1]?]3.52?c&[60DTD-?DDQ)B_3De[OB)b&U&7-(e1>FHaeJ=@4>c9gc\#gJ\>
/T,1S@NK=-B]LIH66JIR+47[)@9OEFFMN/V3M_HdBF4:XT@T5#(PE/0bKQTFW@0<
f6g)afT;DR[YD(=_+W:A<Y&Z\<WIbaRdQ7^861^cAMc+02VggBM@RF<IU?H;E#(H
TV&&^L?-RCO57+SF[MeL#UE;0XCc879LPOZKK2&HU]C\DW\cg)Yg&30U_Q/+Z(BO
657N]I+7ATFS?EW8L;;+gVB2IQMMYCB.fH@U]OD<S3=L\D(\@XN:IL53)RT2TQQW
FLB5b\fY49][,)7BUQC>>8,AR<)=Z0g0C,>,?5)PERSEB8<La_1dLA9,NN]&\E65
VD()O3,J?WVIa]S0N->=8=Y?cG?(^C5TS3I@S/WIAF9:;]-;Wd2U[R_b=cb;9P9J
O=6M@9PBP:,62ffB2G(3F,OH#Q.L]aXcJ63ZE@bX0gIFJ[EFJ.V3;+.<<WRO9;ML
dgeW\[&[T-DXe<20e3+8MI<bXQZ,S#UO.QP@6PdU=PbGEgaW92N\L&EGYgR]#(K@
STZ?A?O(4^VeY^6FfI#RR8H0f4WSa]J^D:&\+\6I-C2^HgR_B7^QU4F#UIaHS>.V
(2ELb-D:d]BB6b\-6<39R-+G8]aUBWVO??CY3_bEHA/+8:8S&AK:U:3b6.ZSZ\3K
RAI]^cWP)67e6GR(cPK&VC,gb>KUa/D26fa.1^01>W1EWVB:G:E[B_^P=2#Z(@&;
?Y:DFT\Z5^cB2_?T&b8K44YU@L_-Y9a3LN,+YVYgb&JWEZ4Z,YG3ITREY\d<WYQf
HdU:::GA)c\<&3DN]F^_>_#\A(_4_7EK2CCB>PJ]K)EHR-Y&N>24]SW@7\AVcQ==
H_Q2PTRS@?]R6b54<eM<Sb2>1#4SJI>BQ4EZBJb@@=>e<OQ_MFaf]0WVa4>Gc>,b
2C3?ZS8_VMgNADS/@\8:08]58DIOX8W&Q)F?2#Nb&8SZfAR:@&ILZZ&<[K.B_X+K
MbCg4,(FB=@SV.#W#GXPMT9\_7/\F&NY?[R]7]Q0]TVd/HZ.bN4CCZ32H/ED1H58
JS151Q?P:F]2Y8^66>FAPT29T\b+<>daA?=2;dJb/3&6>_>T^1#.NPHTR[ML[M48
dcB#-6^fD6@S7^-15>+OO17(YCOIJE@P:9FS42J5W>C;:8G;4dE=;R]f=\b@/JTB
\(dRT)RbI3@?gcE:eC_:O]UGI1=RA+<#GZF:dF7..N4:_/\DQE?NRPZeUBT8K8BN
(1Qa-E-^=gI]6-&UaP(L2YCVW:R4XYc]V]d=N?K:XC.S:\TMAbKJ)IMcC#9W.T07
L.3(YDK::b7MDM7UKXC0]_B?1T1dL]]H=VaVN_EL3dAI]XUHdAJ/SD;BeT(=7J&3
]COJ=366Gg6^.N=,+PL/</ED3eI0+=Q714A^KPP.@MeMc^/SFZO/OA)L1;S-_CbE
#0LX7/=EH6cU9QEUd/BbeG8(Q:=E_<_:\FdBESc;;/SU8_L:<JcC5P+C?2bbS5<I
A3X&LMNW\/F1:GZ?-2YW&</BW\>\^Z[[Z^]3B0@/\>(A]beZPUC0M@CU8ecY\P&.
H@3&7NUAL=/A,-AfMbdFbOO7XJ)SLbSRJ@N>B?U7&P]])P:<6<3[f7BQE:(/:&0<
.=A6C9>A.C@aBKS89+S/\E8b),8K^f0_>:c5/4cY;8>0MZ;[.UX.6db7W:9#IN=Q
NNXBFW6IDRF29dVF=XEO(bg8;CS5-JOfU=XV+[1E(XW9^@\>Vd=d.QT[c]6RdaEd
<U&_::d1&J89_ETIT()P?_c+ERV<TJa_1B:XK7EBGA<J\,FG7dINR_d,2<^JJ@.Z
VATdG]UP8766\_OZXEV^K8JTC[RcXK_QUU2O[P(9^_^F)dXR(@0E(AK#WMcT0:YY
3dLN.;61T-Sf6P<A?]M<D410.&N6-\N[6JgcWddNK\,7,71F1Q?CM8I]P,25G_?Q
<_:\c5QJCLa&KFefQ)Q#D,aQP<I/Z<Y>ZS:g6&+B5+&aT#I&g@+K(EE)0D3<XFL-
eRaHIFUG\g3#52LV6^M>SCVa_G[A=;Vd<Y28geL1>^5VYMMU7]UUeP^>aC?DfOSJ
MJ0WX-7(0_X([bc(?O&VYCK3HH5F=[8aVgYWWONeT,Y\OfX-0E\fS[e4LHdQ?I#f
\Ta-,QAG.G8VD&(;UH_HW9#JYR5JfWJfJM<S,/^T3ULgH/)Cfd9[>fI5Z7O_0O8I
Ga+Q(fbP32=QeE:^07Q_Hc#PKX]^J).>P1/&6JG^&7N&=@T&8H8W?04R@1>FC,aL
F2bg4#A-^TQJZ9WZH^;:3ID^?6\3Z,=G=eV5(De.YOJ:bIQP3dU,f(M[/DNCBVfg
cKBI?Lg5N3A@9A?][,dN7[&==O)?NVaJ-+=bT^\?QBAWC;7YZ5B1:CB[;>)>OP1,
V;HN@TKPF.f=-#IDJ^SS=a#32T,:Mb?6)@(8:AYcNdgRQb)dgDT^;#QWADgZQP2V
1W9K21CbKEV_O0P-40N,9]a>[\\fe#Acd8c5\O(]X4\gE/^&2-aO-[eOZff36YF^
fG8;YH]=FT4=:18a]bI/_S^8?Y?9]AF?J@2OLOS3&2KMDD/#J)&04>GSP[Y)V4AI
M?WE?aG<1I^aRG5P(=RS9Ja++YFI^6E]g^)DNZC&ZZ>8/Dc57g]+fW/R@GI<XV^=
S-SYDDBMJM^;\IM4G2ZFC@=-\Q[aEUI22G@M?AJN2);)H-L2]5>86S3XP6?SgDS0
.?IP;?ae>.P;-BI:6dH_c9=H\V(\W\T=2F?:>DUW.8IdaDS6_Kc0?HK>RC&WH0>[
85DM#;<CZa_WE/cd+:U;(<,D)A^H3-EAR/MXKBgTLAZ@eH^0B,<_9WQF&cR,cK8=
&T7#D92JNO38G^A/;2CBMeXP-(Cc?&9(S^6>.YS,FcaU^:<28][9aJdF&aEScTP#
1@(Sg7=3bPEgLIAJG0Y<BVcT1,\1CRZ;+0e/HNFB+cJY]8Q<aE0P,c6JL3#PKRI5
DZC;_P/L0^^YC8362aHHa]0cg1:98+#0^4Z^1:WYNeA=P=4Jb.4WK=\HP5>F9BME
]b+6/&WaI.FI^\3IXOg+;QJCQS^eL@,3_2[&K-Rf4?RgeCb^c-](R2bf#4;SKQd+
?9:bg;6OSDP8J\.F=B:(/4ggA8#KHUJccE:4RQ=L-OMLGVD6>7&Z=Ye5aGCD8V:9
MI(-72:B,61EZRg2[-3/OK(GEVC?:TVVMGI@LcaG;3Xd?B&<9df[CP;L52_gWVCH
a9R^]/CgM@5Zb1&@Fe^L#?.YIc3:-/MYWC.dUC_]//Z7&X23SE3P@[5D&FFf:5Gf
VH(F@\dDS@A<0=1fRB[1ZBB;=MWJb53N79FGRc1O6<c>XI7g3HIcL8<1e_A\U<7+
+@f\V,?)L@0I4(ZPM4H[c@?.Wc82Xf)H9aM4+N>VB,8Tg;cYCVKU.BK8JRGCO6V(
e.1bXI)[[W=K3N9QM8P@0/(.FE)aU2ZND_3B&?:E2b_Z4PKMXfD222@,PZX+W(,+
#Y@]cJ_[=;;0efK6(0f]HgKEN1Q^/J@X7<X8ZU8>D067-U;I.2Rge,;TFZ&X8HXB
XS#f&<SURAL55V[M#e9<T]cN.8d]9V(<A]dJZP.1KTI8C9e?U(A8c\gYGKJ<X]G4
5Sb5[0,#8<(WZ3)):,;O\28>gU/fQ_K9FbAX#>8]CQ7(^09g0d)]IC^77E=HOSWU
]W25ZAF6Oe<;edMP=#T:O]8.OgB;[-N\3W@VK^IIM5AO?GMVgGd)3d?[DZ:^GVc/
-@G9N8g<S7:b8/(REK8PNZ>Q_=NAO19J=L:^9g282+6/D>.Y2WcM>[ecYN@Q7-d)
0F1+9bS>[CA30/D;+:b+GTP44VKR@#F)cCBGb/XLWY)1JOP3e@,;X;P+[HY5G<P=
aEJ=:68I+SgR0(7PY01+K]+1WagW5;4)XASA1F>d36D395;GH2XEH)JV3C9UTb?;
4]fAN4C2(-]cJ=V^1c1_g-#]JDRBVALD2d&_0fN[aP4aO_-4:E-cXHW_UKOF^-##
<OQOWFX9#,P=9I@b/<NB_&41JZC=f@0YQS49PdIKJCNAY;:5(Z;&QIb3JNKF>LY>
3UKdaT=b8;DgNL..8+FQS17_@4;fZ7>3&EA;Kdg&UU;OB(2>\TZ4PBS-0L^=--4#
QJd_3]LMZS0/?cJ>.,6R7?K>JQ=F^[Ld2XP-V_VW/\&P?5bfOe(Z(d)IfF\9]^<U
PbUT]RFAKdO99/f8;fG?QLZ9aLQ@MPXJ3HX.K]LP7bVCED3L14F\DSGN^-^g(/V+
Z1F[0,E=b__,fJ\X,;LNb#<]@9Zb6<c][acaF:M,g>=3Q4S_9N6LJ\=QPOVNFB8J
2a;N0GNF(^U/L/7FagPfWdSM5#1,Rdd3?MKNG:>OE5fIc\G>PGFgPT3g4e4fP>a,
M5g]K-<-MZ;eGCAJ;aBNTdW]7LdgX[6ULN>K)d=C7[b^)TU4_8IOc\=JN>:A0,N#
(VgTPbLAR<.SK[K:H?aSO3^_T\U2V_MWU8gX2M6QGNIOA2cDWSKY)=27DP7J&fFd
5M^,ICa]LAL:6F9<X>]7W//N6,B4O9_HV1Q?3G<A_[\&G&-<]VR+^cXE:/D-4.:D
f<A0D_=@(M46E@N[.P/b&+ZR,La;YW,7EIFP^RX<=>IV@P4BfC8.F.dW/#&L5XF@
87G23K[UAaSJ<\@WC-EcF1.ZJXBNOB?)g<DMHfG45b0Ba998[0##<Y5A_5-FYaE#
Ubd9aTW:H>G=JW/<4eVJY=R4OQDg3^@QOHD&TfNRI2L6/W4Cd:/V2K;@;I)fN5=?
7MDH_GeT\ggD,gUWY&faNLMP^-]<eGb<S>gZgV/QV7^,FM<X4(ef0J3\]E1D1:>?
ZZD8DFK9dPS/TA3#R]TC>0V+#^TXUF<ZB0+<81E^4.RA-K4N1+F;dgVK4F-C_5M1
FV-9d)^R6JA7D^+A;,@<VLDS2G51+2>UeO])f-)ZV/H9_<Kd@5bW81QXH1:8Sd^_
8Q\<0(P7[MZac&^d#8P<W6[K;8-_S[U7dG[WLg.M&4EWga[9g[\^-H)8cD8EgdRc
L3cW\C+.-@WHVDVX-X-Z#Re?a?WI+beQ0/A.GXe:Q)TX,6_8(79^bK9C3^EP(CLd
f2^\7Y276@F-6=,;0V#dgHB-(@Bc22ga8F/U:7:JKHW>U31&7+..SSP&SQ5]A7cK
RZF]cIPaU=Xb3R3L62M+d[7Be0Nc.IFDC.dGP:1.^6d&QZ(0/BKVX85Z8RBR4PSG
UO^Qf;ZOP6)Q,3egA=B?E@4O_X@C.\+F?c7E9Ddc>e4HVO]FIQSKCf/(eHa1I:1a
LadW1cZRP[,J/E/VZ)TaO#\Y^?GW8]82F60PcM+F[K\ZbD4d;64PQa)?@EJe\;b>
.V[_b+fCY2A0&@U#,3HV_@e12FA?9)f_eTefJ<O9FSQdU371gd1IJY\52]6S454@
A5,daMc8\),(NU=0=89>:V(CZMQ;?R^&G9MW<9c<2_,4ULWY#6YN^BSaM=G)><=;
RPZN6/+g[M]OX@38]P^.2[6LJ83B\QI[GeU,SEM=[O_N--X:X8XNPH^cU\2VOXCH
H9_2/gASGfc&PF\W>?cLa2YFO1=P&+A@L3UE[cST,&[.RZCb6@-F?@c,)@YCS39g
BB]\^cNG3g#cEO/3bTeeZ(UAP#@6gSOB0J+U1FP88_dV&7J&eGUg9_>#1JX>1HS.
X0W=ZKP,3;67UGU#gA#@M8XUa)81&=>f0ZK+]NRdQ#XHVOG6aZA)+^dQC4AKdLD_
Q[?HT&E=KH>gSVLRX;KO+)52[@K./F#B5X>b5=A\/.LU&U[-XMCPSMAO7,X2UcKg
]TN^:]-g@351]C9_TE0D=-SZ-&NY;;MPY35RDU]&>Kg32,&HfbXf>[M7K9T6+PDV
S9@+]0d(R,0>+HQEKP_;+27T?#0cJ>c2O1a(bPP^T?M3@E/)QbLC(eFPTQPY]/.b
D1_HcO3eH#PYEFQP.;EF^]08e965&S9Z\UH,:(-\J&JM0UN@[,_TSBQ:A-/A1.PP
L_0JXdJH9288<g_)H:D2NQ[?9&]103V5=K/&FOZ3-J^N,T2]NT[E:7JIJ,.fJ#Xc
+<edE)6UIR[@1WI-Sd:<c]RZE&aS_Z8^Y(^+(cO_>&:84?dU,<55LMB,=I1FWS4]
&;JYAR0D.==NVJ#(2G3^A@3B\;d0(6_d=L99&gO;E[B3Pa;.HbdR7O&,8gF;KRC9
Ga/QU/;]_bB/;dS6cBE.MgF,CMOg6#7L1c_,XA=F17R,XKbf<[YYW4=##IGM6F6Y
O[Q29RX8&L,871A#GI^;@?>MTQ3S8O#-76fR[2P;,C?06Hca<4X#P\5bB4JD>0YT
I<aYFD#M@@G0QC+C)SgbA:L8G4I;&cf9=g_S,]Z[?[1cH0P8B?PBP+>VCgb7,.:<
OGgf8eJUdDB3X@^==N[EPBS6^Q[LN-O2T@92:[3U>)TUX-/7g@2377Ma&^3P&-W4
RNN#LXeR@Y_c2?@24ZS2P=bg8V](X1-CNDa2X1&.P(7GE6,V3Z<Z^aX^85G1>_RF
3OARJ,.6cgO.=d<g\^ZXZ]ae_5b(?(IeTeUd.65APXB<0E+Z[EY;DMU1N5L9H4?M
g2M0;Lgg#^M/,NRdRaK3;#[A5DG-7]8YLFRALFbCN?Y<[c5@9)/0XYFP;Qa^cRFN
L6U3&6d_E,bfJDT0d>g;25cE9?>M80TFXY3#I032V60CRSY.[24\O5A;.W/3HO21
5PIRe^c/)>E)J1OgJN)=UW1DL.XVDT.B=I#&<_S:&@a;#8LR_TM6.DS@X+OO_8S8
_1e]bLAR\-eUM8,4f>:?YI;QW9,+RDfAKJTf<4/YU1d+eDG4WGUPLJZ\GbISQN4>
^&;A@c-,F^eDOb?bB,RRLee2FCGUKO@.HNY[(4OA,\BDCEbR?^c4XeHF(NK\-HE4
3SZ3Hb,f01SHaKK\3[-9S]V?1/Gf9-.INMN)?WgdCJ873(IL+AFY_P[>WF;fB?DI
4W4ESG6W>5?<)=Q=7;M^J,VUJ46e]]f(+[U8I6e9BFY9a:FMJ?7OS(DK=c\gI3/O
F]@L\5RZ&/N3;JQgWMM(K+g1;5&BbG[N>]6A.B@MXgR(WI)FMRP8\P?a66C[:)3d
(#@?d+d&bSF?dLPXMJ7H195-@Q#T3&?O4/XA5B7,CaW)b8eB.I#Z<,XBaV56e]9)
9bM80^L)MMIYMQM@1G[>WB<@TT]RRH2ZVEXOTb;,Mg(7W,a.C6#B=WO?8d5_0:F5
UM?XFHXE12Z1_dU/LFI<KSB<E6(V^>[S^JH?L:@5;G<XIg]VZ5>+M937G3(ZYa^Y
=PF9<@(K,-1V_SJ)/^0R@A6-dCVI=fb&1MP]O;N8^e6aXK8E]aI)/[0B6d^PM5+G
UQH^VgL^V@I<;M/KX2gAA@(1Lf6Z5TI,ff,,II2_8U6LF8F@a3gO&@^EXV+O6=0.
^cDU4P;[R.VC:L.:5\F=8W=7\4Fd>H)HY^)_FQF:B+VBe2R>57DcX:Eb>&\b=Y?,
bVaU,1X32&^?(EWZ\ES&L8G4@8DCgY95MedC/,+5KLLNAUUe[,A#433Qd\5+U[7#
gN-La4bJ6gX4[XS@]^dPB;NM_S;Z?=4BVHG@P=M[140VZ6@>3/UeQ_0X7-3BU/NB
Mg>U(=\P;g&#S<\Ze5#L[X?VL[,6fD:KX5^dG5D3;N90ATHIJOMg9?eU#aXR@2C)
PEB&@0#W4PBNK;>M2]8XQKf.0[\+EQ<5=RN5IX:UR-?Q2=b=3V#C2D3,L)O5KOP3
Rc#]b2OdDGdLfO0Yg4a<MdaCVGSBe8L<IU&Qab+2UMaMJKV;-JL#5D)g[@aRW+]J
_W=gC:D+N0KFc\JC<-,=-8>1?SeL+:#@eg^\3T)>AHXe4M&:&^L=KXXIH91C8:Wf
Z?TRMB>ZRF<E>:;5-D;_5M56bg\UWK7YYI8ZW=;E9B#;-dX.6U2-bWC71]&:b+YN
F#O/VM6G>VcgSOQAE,+C/_WZTB81J-4;O7YK\=#3beM^GHg-R[PYFPJfW^g,4@b^
1]&Q3]EJ-f^6V..SPTT,NXN2]2#L#Z+<L1G;70XV=2&L6PE]cRa\CETRJ5Z7Q#[(
3/QUM.C50aR9<7JNBDQKZBM>(?]d389FAP4FMO-K?;6W2f8>2=EAI/b:R34AT;b.
Mb:T9D#3cgTE1fOFHD@?@AXS]:U2NKQ&ZMP>@W^]B-VT\D+TB6+6bR0-N;>\F2F[
GW8AB&/K1.D:B0X8[.MIC-SY@45J^ETg97RKcLYLYS:I?dc<.YG><=>D0RI&@N5B
(##UL.8a<;(X#-cS&R+fJMg]&MOZWD@UROHGL[;XV_aDa@(J3SNH41d63=#H,U(7
DU\20V<Pa83B/aJV6N.29DZ#\=+AWb-,H5cgR2_J0T-+K]T((Yf]GI/U-d>/GdDZ
^IBS]fe=K#1ZL_OAOJD(?1Y&3@^0EVde<,T<XVaeGI&@];QK3WMS6aS140b&Xac2
7]Ac(0CK./Yg6LPLT=+^H9+cMANM7Ka(eR5:].TA:R2;3VbOKaOZOZYALaW:,8#U
>0IG7T_T+>51Z8;B6EgC&I0/+S@ag^2>JbPL+KATaN,,9fPEQ2-F4V^(aL=a7ZOQ
cQ1DKLN_8VO/?a@+KZ\PXZ5?8CWV[D;Z,FNgbXIJ-01E@059^ZC3(>OaG<^I=]L^
:b:RF:3-CTP2[M2\fDJO)8O@L5DEVE;R7._T2?4Q9XfGeVZf1GRAK,^g,eVZNJHb
1T-N?gSc6cURJORPK7\_^.S_CWd/eG8U7I\N,4OD5_/=@X-/JW]3BXC^>5OG).W2
UW@43L:?4eK/+F:JaN(bc[?JKM-eDZ&@V+N0@/4fT/C(DTBXHGKT?0WG;Kd/[MY)
.G\?UZM=\=9+89fJ>e=eV([AD>;R+B<4c=,FS8SJH4Y7;4:<Nb#J#Y)@E<?CHJ,K
29:g=g43YeJb\QcIA&VOY86H9FGIJFK=>S8+5XY-=+,e1F/&#.)+?TTS/[\aS+2Z
5[62.Oa.#3,&Z14/.f,AQWgHVF3Bd>V3^WK\/gJ1f):6+Y6]Sd]5;aDB3.+42#-H
#Q_].78RU5#P._WSHW0ae2=.H(]e15?2Odf1[57GIW=a7f0=e&O4&5/a^ec(A/6-
=F68E<g4IL&=@DGVBBJSJ3.O4fO]X<Z+V-BB=e)8MW>R1.>>AdR=QV(E0eST8J,f
F0Ob[]0O.f#&6<,A\3#>O:Jf_Y3@7GNU4L5E84DFI;?;2\66YTVNf55[7^7D0ZR2
&NH.1dD[CRH0W<f?D+.IN;^Gg6:HC;IfGFFF#M^5J:__>eFPX&3/G)D;P=JdD\EB
S)LP#L>]b6XgbN44?@LXg0Q_Rf0\d3+=7O#+O)[0Tce[WN:CFePd(a?-A-GgX6A3
&7JPB:_,b9:[)7;Q1D9>D-F4W/^S(Qb<XfT\fc55<NH?S[0HDHZV?,6b_A3OdW#&
fXRV<++fKOTKDZ&e]R05/06J5ABTU8e2Qda6BSQ09]\3S8UJ=7ZE.[eX<E(EKV1W
4R;E;\>RS]PK?.5&\16,BMgF(gG#O&&a+ME1F(Y^B6BQ=7+FD.;@KGQW)[QD280E
(DZdLJ4C/?D,5W6A@(gbdZT3a\)>&82\L.63/G>\4HJGb=@Xb2aId[O?E;)IZdO6
TT,CM^-c?QJgA8@0&D2fDZC7fg#QO/]d^_6Vg0MR@8M5?-;6^<DN73/5GPW&cU/=
R&R8;;DD?Ya7R^=;-C4[a&VC>(-X590<\V9-^Of:_9-6-A<.\cJ?,NWUGe3;J1G>
RP6-dWZ9D?gHXbQEgQ10^])(D3b4RP?KVI7Ca+BDU3.Fa_BC]Qa(8^>B6eWc0dH:
c[6I;R9T6HM+E.;3e1EX]H<bQC89DZFLE#PVD4Pg7_dg/L,E-H[J66;AgRS]VBYc
MT1VC[GX<X7Y:MAKN?)181\_\=dSfNQ0(,0AZ:93QE@[bV0D/A^/(#KcYAcT4aCg
Q5>g0[eU)LaGM)1#(=,-a5S),NY]F143XB#egLF@4.FP&aD-,\9L40V]MU_\CCH&
FffcL[L4SeL.bgA1d@LC6I5H2YYf?^X/<9]@L^I<Wf#BZDd,&EHHC)C_N+X/EOE<
])PH0KN,QNF@X43]A<bO^;X<-DYZEJ&\(><P@YQJ^b3,6^?AG@5?U;IKDSQgH)eb
,5D0Fc>K4WNA-91:1=2DD2D.M>]+9_(0Za@IO[=>[VZR=Jf2NM-?MN&L<A9S?BXJ
ME1GE&4:Tc4>^Rg1N]62=Z:,>O>b^TT@2>\a\YFaQ#S?gE56)TGaXJ,[HfL]aeYB
FbDQ80Y^:G-GTSZG)Dg<Z^B8T#WbYS?YOG;F#WG2Af\D0>+I?IL].>6?@YEIVJMT
g,2EE>?J>)89@]WZLd^)PL<>#H/O9Q<:9/[]=_3(,bb652.R27K=ZSCO1\M\Eec.
PL>RQcc<1#(UcP7FVS+/@\d?D,GH3/?KE>5);;CAXPgceaQMF7E/K[+\gT=5]=JL
I?M<V\?TTZ:/]IS=O)VfU#3:+LVQ&RTZ<HX9,&LZf[@fRVCBIcRI[b6\R^RC[Z#A
8J.2Q>K\UE\=I_3JBFP3<EY>TQOGHY8&LfbNQS^90TOTYE59Gd5VI3A73Tb8VRTX
UeCY]BF<eU7K:4SV&<:JWP00DNbf;JG/a;XKAT/5W-#W)=gY@0:<#C@93RQAFGbS
/^CK?edE>TT0^W1<c?1Hb;WMBd=HGScV]@DQR,-\CVZOQYQ+^<<&VOP:PQY;#gZ(
#&,Zd&+[1Ae4E.[X#cZ,Y1CB@^&E,D>BP1X0D7(O,TN?7(T_3I=N;GKU\,0\784C
(;RbO[45e^0DgLH.DgZ:XT_TbEJg5&4G06W0&9f(4gE<B[/G^L/DJ583+:\XWd39
f7(O3N6^.)QW&YG]CA^T_VRKgeJJM9.eYXIKS56S^6b9a?+>&9@XB-AW(X<L[e.6
[M^6S_=D.ba1b_fVQ@+)G7A2OX@Cgg^W,Oe&QZ^WED@VfV(:/(2cFHN,WJSFAT1<
5cg8#(?HI\Y@>IRW6.G)N:ZgI0WGKI=;+eD80RK4(bD;Y4>EK==K_J\V@SY04/+V
A#1W+4?B_[)HbQ&OQa1R^4CN:8.FG+=_,<+?K6XQH?X_B[<eAH:f(CMO?+V&O,=N
\F4cU<K&B&/L#;1EW#(2M+L0LP<.J^5M#bQ?gC0JXc1=ge/?E6>0+?SgS3@+IFOf
Ja>K;6BX7A<Z+>fgBBI,Vg+@1ebf#UWQ?_U,D:Qg_+C78#^##Z&Rf,Fa8]G9(<b&
^465,F>gbZa,U/KVP,cM\JWP7??/^.SEMe?R(:U-6+B(T1GTNE#.]Ge6H7)WCE1N
T/4T@8;Y0R#^+FGfXQ,A6dF4D_0UHRgMO4DRWJUEfa1HSSIMJX=BN<HF^K/c,6XT
JK<5;1W=V.XN.SC#-19F&cd:_+ZP8JOY,25g)BB#-L/N>IWL-;J^S)FJVH>bK)cb
@E0?YGRg)B,K6T8;18]#9Q@;SL8^(S;K8Q1,(LM7QI4(-(GL#J=))P.^J@HAA5QB
P,^]0GJPXDU565SG8c:TNCAF?;C^D4U_ZJZ)HF5Ee0fNHWOOSe;Jf6Na)(,d/PW[
Z@>1P8JMa[&NOZ&+NNO\@I6-Ed-VWV9#PP&]7V=@.N-1]FUYV91Z6//CFCFBF7TC
+#A.bY3>+.F,(,a\TIQEQM,1KY^+AbOQZ0<2@>3[8^LQe[C:(QcgT68Y@5f0R]W-
K,G)-<dQZ@?YI(<BXMU+GaE8.=;,UdfbUTK]VgIde?_CHPZG[F:97Z>=ZTT,<<Mg
fRB\<=D]U][^7U>NMK\[AdLW7H&5X:26\X\R(^5)WU4QM9#:7IFLJWYadVCU8Qc@
d8aM68Z_a4[A^=C10e.d1daVSB.W3&;1T2bDgAH0Q2(9f,E>+Y^04N:;6ALa(S,I
J2/P&.(O)X6M8cLDE5[+U77_B^&P8aQN@._>gCLRRCg+;&1+2/;Hg-FJ?5db>dC6
Q6fA_Se/[E0LeP6^B7FCM5&a:cM.6T9)9\#f_>aH9K-01D_ggDdFF^U53TU-\/:N
N1W,Y(V\WX4gSK6W)]^^1(2G9#D_HD]L+eJ_?R4[7Q950dJAec\&UW?f&T=E=85D
?c(W3Y=F#f_9T:,(Paedd67cOL4><9dfMS,;\eecPKG;7)/)NKCP2SZ2S.1/^WG&
O^b,).9fAGgFSP?9D^<aS-OBa46UgRFMDVC=g3H;TLH4JU#?M-)+=a\HY/]:dG<0
7?Y/F/R[>?<MGEQ=\=SBYOBQe=ab3c-+fO9LR-RcM9cITXY3g\H)/61L;f>4]CVH
^A.8LNdEK,?3L,/-8RGGNWU&A49S5R</eBCQ@W51AdS40G47IGV^+J/]G-P/KX>S
GCQ4>)IGc_D8153b(8#WU-B\&M<,\7[HP_WD8d;=_G.PD#4c;He:.6IKZP5=DYDZ
aa#]gVPN\T3SX(<.^Fa=,BK?\SAABRB&7+Q\9C8SI>+3WMdN3F)><1\OHf3OK@\X
H,.IT.a8EdQ^<DRX;RM@&,<>R:NT8<SAGCEe=-)g(A\LYA>,82IU;MF4W]GL@;5>
Ge#ZTdT5C+<\a<gI6(6<YMGG<\D2FV/G:H0H:,.]H66\]L6V/-:_EGVCf5KRfAK(
X&-\?Z(1.V0GY+E^;d[RWQ0<cDRJd.@:P(;8_PZ;\YV?YZE8O>[Z]8dHgJ-?29.C
cULL+UF?B2,MFJRE=0N]If@STFO4\E#Q7<_0gGcV@gQA>Te]P@X.gfcSV69,=Z=4
(Z#aN(1-QQ\;\NW-V#dT<WJ+R&FNWS-QM>)TS1BRPV0_<+)C?Le,5)UVD:87AE7J
/WE[ZQN27@dB<.DP1+9=FETO2KPU-L799b3&J-OLAeZC25:BJ)[ZDf-^5&E1#2O;
dN5Q<A@FJZ7M.1#TX_68Z@X9/B\F[fZ]ZA>E49MCOM)&CI>:PF;=I;:g_c@X#VFg
dFAVA8bZ@)a;,GEL(fH9(#]XWB5-^cReN<@EbbC?KBK,=EOdF&RVTBe]5F4RJW6-
NZY>E;[KHgA1.cRL@ZN-]Z<.S#(8C+W,3-PGQQ91O[Z=b5Yeb&8)H8&)-L7(Y>cc
CF03@K2,#3RO=6LPXf4,eH5.&RUc)(OK;[RFI).SWV]4U0Y^_dK^\b90W>7D4U4\
94RZ,U,Z0OL,E+&,>2?ZNRX>f(c:M&eVYGORH&RIgFIeUIS+6e/;HXF6PLAB17K=
I,/6MJ7_<O8U&P;(Y?4e<LbfPY0WNcXO76V])fUHD^<AdL9g_W\-b.=<UJ:&CE/I
MEX(P<C93Z(4P.;]B-.[<b:8,\A;+1Yc3IF,>Aaf3;SW4NKP9fH[5cQ_91-753c>
5a5E-Jc>RL>Z5HQV70:.#YC5=E/e?Fb,@S;?^<T,V5FO^6B5]\46JWQ&\\IdJAX#
ca.+=H0^+YTb>C3aZ/M(YBN:R.]a9SJFNZ)<C);791OLYBMdG#,8gdKQ^8GXQS\7
Cd>/c,9<[d4(>YDMXQ?3N0:&,7KI&,A]H)2/<X8H6Y0X-Z5>3a+V=-.;YS@RHY33
UUG>.;1XCX)0E>8)L]8#[1<15^4KC>P/(2#A[@a^M.R^C#_=e@_:]gP.G>Fb@OU1
T8f\H^Y+^dB4=+VNIA]V5<GU+RRV9I_UIK6HEL4^_SGCW#Pe[ZQCTKL3M9LVFWTU
+#@5Q7?4@2+._0;?Oa&SL8fRXBP+X5a\O<#?O>,GQ_4g((,;I)Lg,/81Q5b>cBD?
c)41_E\4\fB=c:8TS>f:AfPBCZKb0BaT=\eE@C8)I:>#(7-&e]-IdPe.e\[a?a7d
HAK,3;Hf<)]c:YTR673SW4Nb7I,3H1C=Y-@bFZ3;F&(PJ6UeW=VI>Hc&?G<K<++D
OOVC.YK/<#GOa<(_beASAZeUIJNA]M(QGNe2@)[XD6LC1)AW3J9=2b^7ZR0\5.0,
1E38TTBP.M?DY0)>EC2&I@M]MLb-CJ?KCJM(XbJ)I=_MHJP/_YJb5M;=5@.:g,b@
gP8N6QLY4:b30.dB0a=8)02gZH^^Y<O88IO#1:CabR6O<5Pb0?07bUIbM5::.,VO
&PO7IHAF/fN22CH+)U8)2?J]E\U21fU^\X_2>U@TDc,&#/7M++eZ5-_dd00G2FZT
,bJS(KS8N^TCM:X=.3@;ISc22&BTPfKQFe(ZVg;OAH=CXD7OY6\52CW;Z2QccZE0
:X18VERXHf246aB?/#4K&6^-N6ES19F\O(HXHEL@RKb+-c-U_:9BCf#gNK@\P_<+
:/)PLL6^GK/):;YRA-_PdJM_>1Jg\._eKSW-IMf3_Q^)a.#ZJ7)H?4HO_=9#3aVU
?5T,])4eR]VOKGX6@Xc_PO=(U8^^(/8^Ie<T_U@5+YK?SfS(K,VZ6TBdH3(,[V:g
I9:B@2[.053.f-NKMA9A5,??)F3;c7I^ICZ+<&/&2A&Q<&ZMCfC1dU:E4,\&]fX5
CR\+HF1Q0S1^,ND(\gTP5a8E6gUOMN@af1_gU:S)9_M1AD6=AKI>-QFe=2KOX8XK
LGd(NWDW2GZ5)W@INHf;IMWR04\9F<413+TUPA;HK0)\EF)+POQ/fJP@XEWCR4:=
,2@Z,g0P+T.3\LS(Pd3eI@:)f,]H<6\CP+#30<5?U=PK-8+H)4?#T8<:M<0W7GXN
=S>--DWEJ>YW2V<c)F]&6dL&(/bgeFa7C22ZfJT0MA;&38GdHIOa&eMO5<CN#IbM
4L[J8L?1^3GRHUF>+03.30Wa/R-7H3(C.G4G_>N0XEW?9;EG1X64+N(8JIESb@Z;
/N1FNG2L?[U4eeE0R5#AA:@gUO@5LWb7]:A4.ZCg9L2<Wd]=64@VEC7cKV[bO/,[
cSI-#^;\EO?\C.78(HQ2:?YH7cefUZ8GaQ.P<Lda:R^OCX3?#fRcc-;48:Bd3/)L
#9)64IYMNH@F4Z/PT8/^.@C;+EQ6bVX#0]DP:I>3^VB?,PF3eW?N2].@U?FU,_Q?
EFZWY^RP1_U#Z-1FJC-8bEA,UJQ\_3@EK]-3g/PZD0N._\W-)_bMIbO5OLO[&DT<
W32F6K,Y9b@WCWU<7.>Wd/TWRBbR#ED++&A^AgZbAeB+dN<(^#1g<<4C?WSc)([e
F\7_Y(FUP-F5F7G\V^e1;XL3=T=6d8ON5(3A0+P[L=<9?K#[6=4d1^<5W<O-QT7=
6d.5,W-&AJHX[LJUag6d(?-dgbgP4\EJ_H[VK=b5L+a5BGK9\[I(,M+IT^&GBB1I
?)3E)3>P/[<H##T59>:Ib3>QDg=_Y6IN?a&BQe+8]NZK1748:/_O50(NU\8+W;c\
R91.P1<(6]+?)eJ8H],0->aeKJ1RDA@Ddg>YXK_Bbd<T-0(1X4WaS@_>=37\IKg>
.[3HP9D?G^O@4>WRMB@]I8-/3:)a#@]6^g2f13QE3J[5SR[=eNB)5eKKE_b-D@HW
#]P-AGCPVf8&?5H5N;).LeM2[KFC.]C;NHg,#Z)PE.7??,NE&aMa.<9+HgCQD7<Y
D5M0RR5I_#gEZFV#Qc6@7?cSYE=4;;=9=]7;U#?UCAXXP)B/a>+(;FJg&&WQ@D+,
RaC6f)/7(L8S;RFKVHfeO4BdA-PVaE+#_S#.U#1-1LC?=QV;MC20Lc@Y,>1gP+8>
7(SC/AR.^6;c3Bg-P/R/ND5V-_#f?e)fb,5)FJF=E,/H.68TFT6SI;aEFe.&f2d?
O-d3I\Hc,cAPG6_Ae@aY123G20HBX>G4ZWaGF;&V@gF,;[e#(VTD84[QUBU6PVS)
F?,?.Td9FR#eT;[[:CS:<SbBZ_EM?]4]Y:Le3VE&;_)K4T?3e),Q_=^-<JA]Q<+B
X)bB6eBV5BD8-/Aa2<^(O_-]/DEDcYBX5VB-?+?\OUHCD,Z\e+>R=HT;H5#27c9Q
A2I7/Of1PM.:Nd[4H@P#E?VF3MD2,_4bD#X&TTU-W7(8)C7V#&Z6KCCaW=HD>EeT
R2NYggJ5LV=U9D(D)U:W\3VCOBNVX/]WB[OHY62UfN&N83AQ)8bM+g&V7d=?=A,2
_]Z-5aY@aR6Kc?;R\&Jc)K_.a)))fNGC(VDQ6>:-7R=]7dW]=R2S6QZAIcfP+6W3
d-S>R#Kf6XEcN2&GAB)Y;2P0[:&e(IQN:KQa5;b<E?EfC;>[d]W,X#7NRIZf,F2&
dZ68D;@A6MZDMTL]DbFAX@8eQ&NPJ2N_8PQ9DS)1#+H+C.N3)VVU?Y>R]K4H/7<]
/C\\X@0MCLLUMYLfA\bK8</^/JH-@^P])K5;]O]=YZVbRWOJ#[#P5LaOK@]dKCY@
4(cK,TY+I6/GLI?)24/5GI5EKM=_:<c=g,6DA01H];e^:b>,UE(1V(>?#9Ag2>cZ
SMAd]Y6^]^e;aW3aC1PINA8@5/:BH->0BBKK#bE0GE7YJ,1LaH-SFKZJO<SB<cK0
.JAM2;&QC:?fgIbUPgOAP(Z)/_LD:3JJQV39T+2HG_7#U?aDPG6)N7B]b^[PV=SL
=:=ec@D#L45\bRXMH<?+UJeIRc#17&Fg&?)=L6H40SFcUUd[2L:6&dBg)TeUM1PX
b+L+ad\##C.,T&K@f=^a=f>BP_A)-Cg#>T5ZN16)M5&WEX2gVMC(PY8c^J]Ff>H6
F2a\2+L1[U5WX:R-9/&ZF+[S.H_[:9T2S5/F+DaUHE\_??ZT?Ca+IBe^fN0aZIHf
3,[/_C/DV2:>\e2XJ(EK#9T0GBXV=KIWA7[=,UEUZ?9?Mb5#:(N-.ZUdgTd^?\RE
7>W3;-aMCCMaR0Bg=;:=LMa8e/g@T5(^J3AH#JO^#90H8E+P:V^)+9[\[(_\@:TP
KFL@TOPgVPU-/FBPO8?3=K3D7=;0U.TfHg:>VA@[MDeG3@)TIX3BK+Za;3[A)BIW
(_0@@b-BN>c?<U&8-LE752GFLI_2R#JOYP;DaKQg<0H26Z;d1EAW-)1FH/7T-97^
.@F8@/25YQ^)HEMFK.)dKI([]c:NJd#<;)#29A1CN33QUcE/&Kg9,1BAC.1&@];A
d1f;A,FES1g5-Df<W]==5XQ>S.E8L,^@VNTAK;H71<[Z0KWI:W3J3545S[U^+=FS
E&Ig@E,;JNa,;AHN)7e:P@/N]@8#HQ&50]-24W8YN4]/8546&6-cV]HaBG7/44++
e5WL^)Z+[X3ScRV\=[@-V@CB1:PWLBKD?WF=74UE6V-b>ccadaA0GZ+VQF=cV<9V
fBIVIJcCfOJOJWVBgD6Qa]795Dc>a<WY[/GUQ@:XGSOAg3EFN8EaDAT7L;/Ncb((
EP+OW6+T46J3fe93eS;+-Mf=KV&@6\?@a2R]X?abI[>Y8PfHg5P,EbZP+6B:1CZ&
E7eQFe>8QP#a_a]Ed_QQE[#WcJHTO(bU3)NfU-]O0QdPPC)2>S811.-Pd<[8/P9e
(N64\dZUf?G22H.)?6D[fT&(g/bb)XUCMV1ARAF:[9YNSE2bMf?3e5BM7K5Pg_CJ
W0:ZT)UM(4LC7WFNg;9b?\FeB5+#0\dV=^ggg51JZ]+VN_:b;S2ZQ9;1JJ65-T1)
F[KV+,ZgMJST::7VM^P?_aF48P#[+&^A<-9W6BTJC.d6?B5D,IK8KTd_&Gb5P\L9
K<:_5UL++WF/,9&VN;6,[4UHS,d4G\cDfHEaf9[a5g[#6<cO3#E)Q&THPG.8H&;)
.4V0IUaEF\,=eH#eb.CUUIDYU0,/R<3VSb<S5S5f50&_=@7]B(ZD4SdQ\\f#6ZPK
&>E4MFBUO))CR76>_+.F<&a):bOQ:KS60\N9d0JdO(W=K+M^<f.b#0gYTWTFKRJ(
)fN>Q[X@K_PN37)GEZ9c^.O0B6FeT?c;TE^Va39b,@0Q,#d]).EANR+e^(3&&_F^
CIN^JbeaNX75AE0C=(.UEQ02_TDbHS,H2\FGX5O9cHZSb#[IO\c]e1I^M,N75RZF
SBLLN?b+A(QFR0?EU#NbeXH/Z=S>[]:K-UHVOKOO<PL31,II#Oc/7cc<[>C-#&cJ
6RB+d-Cd;I@6#7@0+@4<7H#275UAeZ(cU^)4LBI#cNTZa8_YRe)EdI7LQPM\,4@d
/Ga?TMQ\K2+Y6/X2FS;F13GU#)<SgdHZB7R_T^=8^TG12./b744MU+#PWJa-_H5<
(+8E4D^4a0E?;::g-420I1M2QY]a9a\\BPE-1VBEJ8,&_a1NbeYO44)UI9-:,:F8
)A<fXU8&J,R\X-Q8E<4@\GKY(=:E5Z\ZH^H[.J@MYL#[J_8MfW[[aH@2X>\XBY<Q
_<41D,Z(@d#>OAeEZM,1(O7:<e]?g#L60<afFFXFXCCB,^DF+Zb=)^\E&DLPD]&D
XT4:H^BFe/-O2VL\f1fL^Bb/g+>>7K.-^b:.(I\Q1O&_+S-BA1,2J0M/M;7PO8HN
;T7fL=6(]O\O0aF/Q+2:6fD-T2COf-JfSUIHe27A<<NHXZA>#9A05E6B(4DE(PIL
7;IZ\[H[C926;6&#]Aa\XH>C7@9E45JZ9?Z/a;R08Q4a@E4ba7>;Y@<92&WUJ5&4
S=>([PR;3+\U:29CSc=BR_Yd4OUa8WW(RP7QP1<:&NB/9aH)T/U#O/COH+fg#)5>
:&AJ)0PH_L5]<@?W+HO/^8b0TS3aAX)WXQEaP>P#f79;>M==N5R^26XeODLTXg23
SL(:-eeR03gg+PGe,EFFO#XMOE:TdO59@4M[O)Ib/(I0aSB6]WC<5/a):Y:44Z,8
BR0b7>B8e1BLDECIK,g?H2JAf:])T8ce#<3].V5T[E/=;c)F<KMb(/.>27UeJ(I7
\QOJH96adL_@@CQAZTEI1:edcKZ;)DMWD-E[OIU<Rc./-G4Ncc#a^BNO5g\H.c[g
DF21a&(H4Y5CRB9?3VLfe+K/,WAL_Lg]DAM50[K4U24I0=fE&N:;a<Q#H_ESR^UW
GNdVg0?)c^Z&)FKgXHJ/CXK/c/N1CF5J8,a?B?VRUHPf<5AK]b_fP5M[+QX?P]ea
cPO(#&99=TL\3?GM&[Z@B^2F7T3,Z;#,N47<8&;6.)\:TOV1a_=2Va,Y_2#b,3@D
R\[OCDea_HIWD?W?>2+?\?56Rd^K/MXf\eS5V[ZdGL8HZ:BC^?#UTY=A]N^I//N:
U:cQ@&bHT=\DO4H9K:bBSPSXe2QNDH\1)^e:f6+\IS?YF>DYCTNgbfOKR0L-1I):
:6)[c.=XLRHH:-B^1Y+I#;@5D+dJdJL,&<d3<N:L1RQFL#R7>_#NLfC/#=?280Va
M+)E^HF^Q25GKRSHP#&[ZV^Vc_\;W#KIQ1#O.-[WD-W_a):[@LHOge,9UN7.b=f1
OV#g[[A#2DfY\L,H@.Yg0UXUZDCc/N:/GB#VY#HJD&LM=-H9gG_C0KJeG6:c&UIP
;BJ9R2W14QMHfK?B>&6FDZ,7U?V13Oe((c1=KLYa-H@ZC_K0cGZ^P?4YH#Eb8L&@
J-IWP#;dO2[aKO>AT+U,S0L;Y7W4a,MQJR?_>PNdNOMG)/9WWJeL0\B.F1QQ6T5>
cIM1eHNJEJ^,;cS&91##9))a0V/,gf;abAVZ0GLf]/-M\_JbDg9E??IZ:a;Q#M6H
9e71<7fZXS]V_Zf6XKg\Vd-6]cGQU]#)OcA(3e]gHOe:VN,fgcNc^^MW8A6Z)#;#
/9=eNKL@@(@.\c6^0f(R+KPFH_39.f@c)7Y.,]@a_WS_-6a[RF_:)AB-..P>H.-G
N99A+G\Z\8#6b=BFGRd5U090.8-#A0Ue&O-0#GYTY]fdKXd#C#)&eXSL>a0.=X9K
0PRW9cTT.=8EG^E-4IbZ,bUR>)PDT+3I;TDSP1R?X4ZA27_6:L0HI^dOcWZS&LW\
@aI1TUgLZF9=Y#XeUZ@8BbYB<[WN[3-W-,E91<L[[>eXEYdW(aTb98X<eB:+c51-
F^Z3f[-(>\&Kc-RL]C,U<LRe>B>Gf4(eW(@c8V)2WH]DcOB?J>&CS>;NdYS9f>S;
D=1H,AGH,1c:WebAU7a[6]WFK>0HAY99DJNeEEIcO7NC4;?9NWN9d:15]EM(ScB1
53/[:\6e?8D+(\;CBA;bS)??F-X\4[.F[_O@?L66M;F)UBObQbgH4:B<.gb4ALGB
PU.3F,Q=DBK9K(/Q+N4W5AO3F>4S)XbbIg=@F<:FFSfV(e6AH,C/=.JBJ3CR-M:>
..-/?3AF(EGDHQ.&,-QS?VKPI&E,2fRJ4cc[,9B2_E\Sc1fR+O0Jg+MHKLEA:Q/:
L1.&4YOU;N^CO,H-.3.(U&1^.A8dV<68\JQS>\Z3<F=2d5\J1g=>4EFO,[1<9+2O
L+WC.8R2^1,B8H@Pd&_,N8(H9OAb_[V@,)_?VDY^W57?ER_,=ORMN84]Z>G[OJ=#
/<a@]RH?E^2Z](a];d>[4GUN:??PM,/OcNY,-V;3Y7O-f3NWWA&H&F<P4(Gg[TXX
-[JfE@<>_QD)a;AIKKAEXF;]\QU8M>\/_Q-2@;R1?C/(+4fQO6fgIII^#EZT77L5
RVbMg+&G]Z0]&^HcKKUS.J])1VT4V2(SQ#gGe^8V-Jc30^5)a^1WU2gFT303:_MX
J>3(LO.0/@RV?2ZbR2[AVT\;_a<CdC+N2YBIRIH:GH[8\IK8c<\DZ49Qf3XC<1-4
^.WK.f#27GV75\cRQBIebV7bYHM@YTNE?4BJNU[/D#[26X&5<86M0g89&23+dNQX
B+J;.O95e\gK0M_IG,;<L<;S.<9214Kg>4^,]QA)3MQ@85QVKH39XY#MAB\#H/)>
a;bEQ@6#TN@g<O._Ea^11BT;eE+fAKM&PD@NXe542E+I0=df[/)3eG-+K4b,bgG1
ABF0./>a#b=TMA<R-I::-KcBAa6b4B5Q-b\WU+TdH#M>1c2C^G>R[YM6;b#V[?De
EAFagZ)853]fK(Re^T-I?+MI)<FQ,@,Q>F71#a7-;NMM6-W0W;9LH-Wc@KCF?(9V
_\N>#0?dC(GUQMNH?<3NN\7Z+bL\W[P_TE6V9/<^3f2D,7-9JbGH.2AGcN&KR6gB
W=.LC3A\B,bc(XU]#fIb0A+7<BP6:BcE3[GGKCDLW6Q;7WZFe<2C5P]D&._M#8]3
gV:2A5XJ<gC>QfVPgd9?)F/ZV];QR3N:P6Zg0UB&/E9T^2gd9K<G(15TZ]?N+QH1
ICH?3^cb+FfN;W,4HCWKKP9J69T?A.>g\0^.Q9e6ZMP#0]PJ[2;R?O6FM?AE:,(c
BJE68a&^K1aUaDe@2A[@)7-HW9:aC1+(RXV>H]>BS>Y[6NA&&5CR)&c@)B>](X(?
G7(/D3IZ)0J40?Q5PI0#<9IVB.-bCLIdF\&^SB+Z]fK7Q/<S+VTcIdRW@W?;3agL
:cLeZ/J<dR\/bdX_bBJ,PO]YfYe3EN-,X>B@9AQ-O.A5Q@NYPKg+Ag]RDWM<6_a:
A]8=0L;UK+#a(eSO_&(17YH,Gd3SPdXfQ@VSV@F8Ue/4<>Xa)>cF@XP7@X;@5)=]
HcENE9@_[^AQgYfT]54/d_<WTRe>D-&MNCdMfP<\E4?#KV[@>#<gF?G0=HRWQ+7;
TTg87FHGZ;>:#<c&]J6WC_SF(e,gGC>F^J4YMdRH\J)ZLKBE5#Xc.HgET4e1g5a/
I-SM7OTRG:A5eDES>7&[b84N81(FZRd&#Sfc_UHD]dC6Edc(C:-bB,UPQ3BW1)A=
b#DgJb.fUd)d@/K3C[bVgCZa+I&I)4[fCT5]V3I9+V#?:b=JPcP,C^fUg#4;N_)3
M72KGf_>QgC3,M#4R@X[KWY[gCcY-d4W\CMF:DJa+4S-JFaDW]cR/Z+ON74:a_E+
<TKD(O&H14VI/HXXX[I8(c:\bb(##b6fU<LZYQG.e+>16OS+<ZL=?J+Y=\7C6f/_
MLfLYgC/C==0XT718.[TT1G\EK^(6U;2(]75Ba:G\IWLFQ8XJ\:=KFJG,CIA:8<1
WV1/LCLd<H)KE>Q&C=DX#.PIfg2KZW_AJNFKKZ[@H>1/\ZCDN8X2J>MGO92A4&^E
:.ZWN#YW075G&D];b38JG&<f;[QeMZP0DI8NWS@ENf=T3-cNQ95[E1ga0.[d?WU)
(+-((FD&ACQ9ObEWBJ&X:#fbc-&fGX5Z^#+9:0Od31):NWHO+B57\IY3:NE2d/)H
OHF-B3S(KCcO[+FV7T)BX=FdUHI:D.5(_UI)>8^_c/W=,.#GKTd&NXSYbEII\dQ>
Z-?:;VB^)86]5eGA_gYaN3LFFfOgB2g/O\FT]Q6PLO.+.BW3S]WW+.R1#+b#?Q5=
G9X\);)]Me5+&:[CfH=fPPScCEd1VY\VP().::V5)\1-B\Q<:]/)F3Z6YWK(TV?_
&_E<=^ccQTc51[57:D\GFTC^Y9WKUWCg56/4I716,JZP^UNT)1?77#0L4+MbC_df
WS]UWgKB);Z1VL04,?;8:TST_c]?9I#14ec(V.baIX;&H)UX#Gc3OIa,UKV;cG0(
E>d.,W>.EY\V3+JZ1PXJSggGXFQ<:0,EI.V;H8dBP#2BOO(G6AS972/bC_2gdT&T
B41#ga;3a;[367Y.YcWbL<Id5McX1-a=[(Jb)L<,@+S4Se1D>6&KZ^HId<AQb=:,
g6SdJEH05D=<Z>7C<<S<F/YfKb/gP9R,DFDKEB8eRK56(KE4B>ZYS2)AJJg:,H?<
4U&2dY1)6;,WIJL,TJ2@e,K(+8]a0P/F80#?OCAOP3]A8E8eYa3#8D)Xgd+<64[(
\7Q_]EY=Z4R9<XeL8?;TL1V2()MNKR\;S0IU4YF#6a0+(OCKBZDH<>>-]dGSD4N3
-:?40>0MH>D;9C\C=I6)Sd\T2,#RDMQAM+;SV6\H226Y4fL^\/4H(YCT5.;MLPR#
BLW9B2CA(TU]S9WeP.&]0VT8[/eM_@:+BB47WFeU-@V;#?b=GBN_Z;VLdJ2H0J17
8+QGgQ\,@.2<e__;@+QUBfA@6>F7^M5S>/>acJ,0#?JH4@T(V>U_BEIb<8^8HJMb
gbQ7-O]0Ybg#_9P^+>.IB#UK:O3/&L3Y&O4W/&JN(=)6;B_\)JBRP2G/]J@G&ZWN
&Zg2^UJ(UP&Le2T\SSWFf(9K4IWcHf1:Y/e\92#H+\?0BT6Q5ZE?;]#fLZaJ#L,8
_d?-H-;d(GKJMYY:TBUZ&,J]&b@O@C(5g\]UCJ](M:<@Ud+WV(Y@dgS_#)7-,Fg1
d?NT[DbeH-_&8Y7IU[RUVPc0><&#DbT-b#300-<=PS)#XAdYM,UOTX^9L7=7;X(Z
BRfS6NU&3^CW>N/(DK;6U9E+<^_VMK^HI;?6^JDVNW+<MMME/@bM1C,PbcCM;F+(
_C-D5?e(UA9]LFE((ND#GE)g5.@fL.+;JPfc]K#,//G=5BO2B)dJAY6R]AM79?#/
T7C7e3eg;^,84S3V:6T.#1&Ef-8ZZ=;;=(]9a4=;D-\:2\fg8DNQN,.Hd2H7<3N#
)@Ab-IgM-@M)YM59I8Jd<A-H&D,(DX&O=2,6G9HHJBPF.KFRGW60T,-,1MQ-97<>
bO>\WPCFYb,BQ<EH&g4QQHN)5SKbL8UXGGg^JP1L\Hd(Gb5\FTQ5+KCF:,Z\O,TH
Y0,g_,]I;VU)JOHIR(bD6AYT;/=(4S5gT^LQ;NBU10JPdL,-TI_)9#C@PeY<M8_/
dFaHf,4T/[Y;;-#\V0(&]4fFJ&L54-[f@#PSc:KFX0??SP,MV7f&B(0+9I64L?^f
A@3fJ.Y::e&?N/#UfQ.+E;R;Z)][&CM0:TI8=>=2Na7;;#]Y2eMQ,Kg.:68#5I=_
6<.HfVWYPF&&?,1S=_&\c,L+2?#eDO1XX2T]:.5e)03)1ccLgKJOK08?]K9>7C?9
&bX.gMbX?#^,cb1a<&T5a^4_Vca0&=DGSEZT7@U<;R7/]e,EceTQQCE2R^XJ?Z(\
V08,M3#e^?1LW/PD0aQU9DKT>Z\9UZf.?M4Y8(B@.=0e/?^.J,SNaJ4>W8LO3\TL
BVaaOP4L\,S]QTf>.af+&K92;;;Q&QUC-[4((=ODO@P9MDF@#6Se470GT,+f#)f2
ISZHX>T&+b:/_4W<56(0KRGI-^I_:S4KN4L;K(][\c2aDcI4IS^<KRGf<Z-f?NeW
)#@19BM>ffS,AFFGYAe9G_ZFR^#;9@M7/-PO0/cgEffZbWZ8(7].S6[:g?H:J/K\
eIgXLG(?>=9&F-dZAS@Db#_c6PL/KW0YTHCDeF:?_9]YIV90+HTRP,0&C)1-?PL;
4))QgJ3)48ac\,1c4Ee;>A&,V[XXN0/X<g=^^1&(<5^88cfH3dJgARVRDD3g916^
Y4K<_X1T:Qf<J-DK]eP)KQTDbV7-aWf8RHYDK(VQ(>&+aeHE]:g=GQLYP&F^_)[E
N.Y]?\^^bcP=_<+Of6TMCV#J,O.O_J;>_,KB&e<.Q1J#]7QJ2:-+S_gQE]Q0([7_
7)4F9^01X6&H-)M(ffKIS&4f[/>RU<Ha/YUa2H-.eNS-C6eU]D1?,J6K\WgLU@.;
5.G\LWHgXN>L1U?/Ie[BS/RPgWUK<c#WZf\HJ?F6E6:X\UUW1]XS4TV<U/JB5NU@
\W-.MbcIeg^/W-D5_e,:6LBT(]B1M3WQ76bgNVO>,a?3=cRfJ8U#bTU3D67^;-82
/QW81?Za/YP>T9.=.+0/;U2>AbHG1GSHMVNfd<[8SY-D:55K=3)/Q?N0&DL1eQBD
Q3H[8dc[6F.Q[/R6GL,>H2S4W<4IF2ZPLHUGR,)Ef-)UZ2I>75&)IL5QTN66CZ&5
7_2^B]]-Z)XFa)C1E-<3e.dWQePOM(KM/.?:Hc9C+K+E#,T]-Ie8M)CSY(8b:]NK
A4g9?\b5OK\2JMC.fRRc.M_d=<N0ZK15NNdE(Zd:UB8AN9<\961B/W2d5TU1#bF.
C/d2X9[P[<J7L6d)c4(b(AD#-1^V\d1ZT39,ISQdGC#1_fE8e+Bd+IE,fd)QDI(G
;P,cKOc_GZVY7Y8QgKC5+d]a\(-;NMAX5c>AR^WBg\QK\\]\68Jf>VZb0cE7-eQ+
EBS;fA@_2FVH.dA=Dd8b3-5\@;WF.P?39T/K9]\KZ-1>HPXP8[UJ;<SS+5f7SWO&
O<Y5WKD:BY<^L,F,?.M/PPB2AJ,G/TLZ:V-:9G?97b(cQb57L5cE9/:cC)XW?TM1
4NK35=L/YaJRXSI1W8AbIIQY-?[<0_;K&&gIJE-9R,3IQa2d=]A86NKcF:CdZ,GJ
/g>R/Ef1,GW1+46:,eTcAEHAZ+C?CEX3[D)(9_ac)QP6G\KBGC3OW+8[],Sc+LU-
,@NNB.EV2XW5JW6#8Z,><J@^g_MgH8_f(S^W\79HI-A<@JNB[]]-AA:ST=]JB#_&
G5EU[NRG:=@X/IIH4,PO_H=Cf,:De@X_+9M^;+5>N)6:^b?G:-11H&UU=c_PQee#
F;[ZJ9N[f+JF9FgfX)a<XK1V^5J_U_G_/d]R3+2e<C..2>/K>[e^=MM5:f9?7GgT
+TBd.-#_)=1\(F#)3[Y64U[>VB:SfO^EJL@6^)^.9>1PH\IP2\]3MSF==PCBX\c7
HRA988LQ5/(9aF0b,-]PV3E5Z+CHa5@]Z0<F_6gMc.(H&c,e8\2KU[AWgPWbOH.Z
;aK,DF^0-SZQ2_Y+ROMcD&7A4<?bI:.=dbJfeeL(6^>=IBNKgNa[NfWRFM1HG^/;
A^>5g3_gX_<.NADWbN+QPXD@CN.I+P.L:Z^@CSM,=1bEE.0EF:8R/gAUgHF38bIR
g?O_=5U5TWI,?b(HER?/RO2gD<VVd(?WS<Xc2YdC-6#3MW;/:YWEL9e.T0JA/NfS
XOA-c2EUNP\(RGO@IB^D6aOAQ39NQ,(WH?;R@,/:]60\7#;1,fZ>M5cb8Y7CRSQ(
g(;X)c>WZ(P<5@PBJ2,>\^V2OVU0Z#.^.aaG55(XfNP<^NSc\P@?C1DD:BF,XSA[
&g<7Y6]b9A]-UI.=f&L+YQC0()7DP_-8#[V1;Sg#GAOS3T-\BSX+Oe-_[^Y(cEfL
f7-EL<[C?/a]RVA->f<HRKS_K0Vd?8@M+G;W]-_<8;Z3,J.9b<&X]WGaL]Q-R=F;
8?0[B2fAc+/#V[R(LY4DN8If++F(1UfTPZ8)L)27/Kf-6&8@XaL&LW1V4-PBa#(H
E<]Q?/2A>E-IB^A)[21_-fWLXN[,._S\ZcT.-Yd]O-WPdDD\\0X/e/DRI:6V#A51
d^N_WM#E2>]b4R,-^GUA:c,\YH67Ud>,6U1C357UIW:SURcIB57gNdC&d[1,8,#c
TL[#^A_.CVY#1,ON@_YJY8NeWPUO<#WBOH@MbTOMHMHVKYSHKTgfZHdYD7A7cAcT
GMPU/dX)UVOZP[e,J<dR]U=f2JI49/5X.c3VCbMS@K.[\8cLP^S/0KHJIb2A[:/6
3BP)&P)J#@D]0V+@><RP@LUA0&dZaR54@4dKLBQ<K04/:eHf_7R<A2/QKdcc:^Xc
Q1G^@B+/]G9H1>P1FQKY<M2.(U-Ib8/fZ>>BQ+(g<BJ_&JgV)-[XA/eD5Q=#=3J0
eDHd@JH+AO==TCF)TX)TOUXAYRSc-TMXD,:1.+f<XLdP<@>DKCK?=Eg3SCBN.\3>
GAfd8_BPNM[CR(-13MTC(1-8JOV-3TW\IX0NGY?M-cIBK>S_D)^aZ1V?NEG6:R#G
A#gaXWS.IZd\_dO_X=e7A+0T8(2^JfgL??\dZ?^Ub(SOY.SW0CY8dL<gTE=@eY)X
&bGSI9VBA@1Me?I?F8a=CDJ(8?LQb/@A/;#EHDXHc\I@ES6,EJ.eZOVHdDGJf/BS
I)2(e<9YQ,Y&Ef_gP^>1D5]MTR_ENYZ8YMcCW<aPV,gJb8DKQGGeW]8]&Lg9Pd2<
c@N#>Q3=3MPQM^X2TB<d-DUSA<UNC7T>V[R82RB&MPADb],GNW?X91/4\^0fN29\
[C>.&bE1\DDb_7NKDY+4PKVKFA0]Be\_2\[RM84d3?-cR69#6VV(2F\IZb#VV4SQ
@-4J)NO3G8]_^)T5@2fD3/Y,PcL,Efc?eY4<ZfF]Wb6aHOW5SDe^H6SH]M>UN^SM
^;/P=P<+;<PUVcPM12:JS[;3a2Q8C_58-5QMZM1HCefN)93=<3a^9e=V#2B\Sb?O
fBAT?Z.2D1M_->2+-e&GFL;Y4IeLOgZAP=5]SAA0CK[]/eZ_3f:RZ,6KbX0O4-2/
^UfNOO(Z8H0Z-d2];-VNg-14R[,8a3c41d2aI83J@H+P13E5&,J&7AH+eJceYBEK
>7RZ1[3Ve@5O(R>#-DL>b3,UM#04G[b&_T3,QdC=1K)c+B4<<=,FbXPc(XS:>9bY
C<86_C(FSb3>#:7(CU_S^/EKKFK&6D[;GcZ7(6bQ)YBKRa]cdOLQ4feYOI(SBNB;
G:4\0JScWKZ]X)VMDW=7=>2X8WF6Q@DOFQ)\FIR7GaITN>C\AO9Z-XTKeW:9^7O+
)YaFG6c#cQP6.2fOS#4XA_O:L8;G+8&X&0-]?4d[@b:@8)S/:/:)_4]eU]&gY_51
V-:F]N5NfC1FUcNF>U:E5Y1R[.D&U=;57X;R8X#\c598J:(/gUc2Pc02I&5Z15LR
O\ZIBM59T2d(aLdTF)Z;.9BWDRMJcbBE1)M#:H;0P_Y>G>&Q#D:Z8G35Rgg1M_D2
,><I4\++M\=MJ[cd2T;3^B7/1S1K8:G]a/MgaT?(PNC6GfBQ)L55CGIW+E.A--:W
-7RTWB:ab0->M]dY)-F.)4]d=8Y):M7>CJBZI.T]&43McML4F?FVfM0/,&W_<d7A
b#1KITgdA8W#AD;1/>9;#dRS8d/Y,H6]I1Z/N_7g.(&/Rfd[-/R8OL/QE^#EFe0F
dHOO4;,HZ@]T2DFR]AV_+J6]@VPZ/23Lb(4(^cM5e;TT@VP2gfD,U)J-X6,.]+dU
YdF,OJ=])CWW_/4g5G\(41bE\4L=N5-C,UR/,K=\<>fH:E>P/FLZZ5:7=YFH14f\
/5NFUH,OfKIBYXa(UEPG5KOcVG(Qg-R/\R3EO-d&>HFdU:B9A8(D+eYHL.FLLP:Z
->ZWHTO4Kf?R&2[=Q/:[[?[1V_I+c<IY^>Z-bW@/;,/8fR+G336bC+C9g>N?.,cI
SSE,2FAW^[b_IXZbDZ\@?B1[G9^40V0#fEE(R[A/&fOL/D_c_@1&7d3f6&^E1+>_
+0O2eRS8SW_b/7?:ba(U7:g:]ed=J\UJCTD?RKH1WcZDV^;Lg?G8JT9(E2L/:2)&
-<^@1@NBI@4JUgB]]SONW]ZI?5OM_4-(W)UBSXbG[^2SIO[7QPF2-:-01HA0g,L_
R7^+<Q)D.&?T(Sfa4+.NPP6XM^ba\TP<=9P,^;e9-8@R8Q-(A.;-A;(B;+BGA\Mg
0;816V\/&[=&CY7Z_CLf7@fEL7N22L^f@E+dT^>;KR&]&9,01eM>9CVM1UV>?Q:^
/X9EX#f7VO[5L&A\L;UU=&Oc+40a#c+AV5SH@\S==UW;ccc:AO[RZ_,U[VFN=WVN
M/3DbDgL=)XgI-J_7GFJ8=@3V\@2C]2@=VYK;G^[\faP#E&=)FKK1>SQ9VdDaSF&
Q1bC1@eT<4P,KX@2QfF8IZ^Ce.-\^);6^3/4):]1IA:e2J>5gO[ZNE?0O2(+L<LD
a-)Z[TbT:U5GBMBHR#G9@IV;7T+[E&:-2GLA(ZHT/Bf&aJaCL#=#NB7UO&AD?NYE
7W4R+Od7X3aK3@JD\)(^GLAXZ@,3&VNF2.&U:=A>-(2AK59WSdZ>/?X:;(KOP)67
OZ_Wae?EfgD1.B)G7_3M@TaRA^HSQf7J<)dC6NY_8N#1-/9dH6=3]\Y#7&a;6WK^
1Z2:0NMg(c[72O==&TL,HUX8YNZ_\8X1d6FU[07,;+592Hg)>-SQN3bbN_3I6I1.
g)+#Ra)NW?D2+\M6eaR]IKgS>MPKL)./42>+>dA](1R7C>Y1fb-7a]@ZcQ6QYW8b
MVfR8)VCVX?58YO=P_e/+OR:(R8,6./73@\(YNFM[4-b5(4?g@974TZ:;HgUZfI_
cZ1THB[FB0&QF9R0\CZRaPL9H^(IMNUMZ)a\&\.\:XQgPgbETR]6D5?ETH44K3fX
\+Ua\FV>6KI7;9eD@&VgfNB4ZB395@J/&NX^f=gK(LYdZ#7\OgO?IQJNK)E)Ka5Q
Q]:bH#;eGWdBSg-I?X;HD;FZ=2+g(GTE6,2W=WZ400^FP/_#98Q4fKZCQ=Ib[JC]
f<8C)7XB5b.Zf)WgC?N_Z[O\][FU7/(91AQ-B38K&B6gSOFZZ0\L6C#-A\=MUPe1
KX[90Z0,_,XMN5=EL,@ILF.-TM:A1=f69_5(S3AEUNX40U0XCXN0#1^HC1-L9Q+4
K\&(E\bWEKBH_E-JcJ5dZ&8Q_&B_]/.+0\IM->1JPZ<)-Yd?>@NA2HY&cR>Dg3>a
Wbb)1]V/KWA)G[dRR^Q_Q(Jf.L.[)PBF\?<[fFUbKIeQ#c?B,g]3TU?W/@)><U3E
gWFIbP.^C2]^g08NZP>^9CXS&XMRa<#(<b#(<2:0dT1/Tc-F\K_cfTWa_a:.ERcI
MX+PM2&faO:?3NK^ObWVbQ&5TX:8+FgCW&XC_27@XWV&36WP.CDA9SXc,#a[@&3]
_4[c>GAEZ>ADPfM=/\L[CGdGOb^^^[E8=ecF^;BRG&4DMBL9GC9[##F,K?R52?8O
GOS+3R.GXL/D48#^M3X)W=IFH67^_BCO8f:.JIW(]87XNS;b1=X;)>0+eEHXe<S1
_;PIH)M4925Xc9;V48KY@:C2a[NcGT-)[3(7IFUc\]MS_[>49b_.Z(I1.TI94V7>
P=V=M=SMH]^9b+#b#XfU&Obe2;B/V_^a8BT[U]EA1]:28G,:(A@9aV(O6J2]U)5)
G=LSf+33#dJf&Y@Yb:7>G)0HH;+bcN^BM]Kc@0)GUHSO?\2PUT<MEJ)b8#F]GJ8Z
XNL8]_ICP8-2OcHSCGVT:5HRfedNaU0H/R5E8QY\UeIM<08;GM@@<P0D^g2VT(:L
c@5B@XF-DZcJNWbLUS6W[F4R0\OJQ/^7bB@((-24:g\dO#JW7=?8ZD^Y]XMEX\89
UT=//5A-@-8NYUZU_\R<F>VWfW0@VUcMaG/E[W5dOSXQ3]I5Q2If449>4?TL)W,+
E^L^#[Q;Yg4CN]^JMQ2Jb,@P@2K:+]EM0GX4(VP9JV??F1g1>U0&cWSQeA<YWBBZ
7([@>NHPK@1.EYU?Hc(JeZJW4YaFUWNfOHZ2V)cE7D6EReEI<N5/d=L^D(DPGKKa
QQbXMD,9aI=G&f7E5YPH38d-WN;?,7T<dX<>7PbOa2N?>/)bZbcS3Uc=8e&FE@8-
/8-;[4/4G,&=/]Q<&8e7E0<MbRT,8>?KOJ&;=<@(-e;C:Q5C;.b@1Q;;3<ZFMg@<
24.0MbZA4>4\Yc#[@P57cR1c.K#0Kf03(9&T<59M2e\E81?W\O0UEA[/7Uc[;6SG
Ab24S0)ZfY[<F,9N-dZ9A5^dR/<VFWeNKU+2W?fd.:?PA^5#d0VgPbe+M4A2]IA(
]c?Y]7ZCL2Jd4CaRFKL<[[gNBH^E1d\R]g9f15g+VLTZRVE0KB0EF5C]EG7FEITS
J@+bXFQcT^b6X)+:cD,:G@EbC:ELQ9E?=@TCaYGJ^9I[g-9L>D7XV7Rb2854_#@_
>^ZfCH85#D#5KT&(A9(ZaK.e=g-#GPee:]cWH-(XUQZML&B[<?)_/BMX^aWW-:&5
8/@(]39aNGe2]-B58,0#;MA;J44>@4F3]\FDQ>:K0Lg>])R].&[/f/\^.5.M.9E6
8A_[RI3IYK9A)0]D31bIGg#RNY=YYOMaBN,E?]UZC#2f;-8RfYQ(Ta(DP84=&]Bd
_@IB35H1BU<a8):)?ZGAaO4F=f[/1ZWaDC+4(H=eXE\<_NZ(>]V:&3I#K.KH_Ue7
68=6;FSIVX_GG1T7e/\B4ZE8#=g)JH43b#3&Cgg,Z;CGFSW<be99PV/Y@M@[GO<1
9a/-<K&WN80;>RX[#>g7bdJ-P.aYMg(\7L7SGIdUa7cGOP7<=QVIL;Q1&WN>^93g
C@bEI,9SaR+38^+<4&(&ZA@S8+G3;-P),0CTBN2AM5W&.NJ(/Pf8:^.c=-+W,(6F
9F>-XgfCMKLR5EN66RKJKCbAB-d6Y]bB;=d_Q_=8\5Qc_GY__+eeU[=F-O);\UH6
Yb/SJ7K&aM&GgJGc-FD[V.K,#E6LH9;ad=TD?6-43e>D8Ab[T3IQd@L?=fe^:6)M
a_+3Q+KaX\;=\3D9>g,1?-;Yd,U]W2Vc?2T^V-W.NO5RE:cK_X[F8G(C:^4CXW1d
^_#Z1_55,0Y.DGSQb\M7G^CIH1Dfd&ReR,f,3GCG#RbA39X_^\_S5->HSdXT9?HU
aQMB;<ABS>U70QN+5a\ec&&&YZY]79OL]<,f.]-d4?;^8MFZ.CN:\d-M4R&78;eZ
a]a_dCTOX+Te[&IeeY43WCB/E<O[cCZ_\#bKLa:^=Q>G#+OGL6SO?UE=8BbcPTBH
@dMYM(IMMU>XAP.>N#0:/YC+BO5^<)>U04Te4<<S_W/O?g]@54FHAIZ==8TY1FO;
.V=W07(8J@+=PI=c4c[MI@/UdQef=+AM&,E<I:8A<-+1J<TfcC(=:T#Z1.[[:A/@
Bb+C2,-,bWNdVU3,:M/Z06=;NL=)\0=HNC6La+c(#Q7=NJ5CU.J=Z[-MK6P.32+[
]1YKWSd;X3/.,PeYOZ^cbfAD.f]COa:^,8K9OYM=EL5eR?Q532FALHSH_9?_T\O/
J:625QeA(N(Sf\+5gOUA_McGA0SA=0S_OF)7))L[)FXdV85YS;=01\7LM:I7N0?+
HAfa71D,[^3Y?TS<.V@Qf#]JUZZ+JO;30;K@99V6NB4/+S]<I+9:;??+GU+[>?8X
@D,^)L^N3(1S)NZQ@,S.LDJ7N#C7=4FLI-=7PJ6[ZS:A\,]89S12a6,V5cUVZLVN
UBC]6OA^/e=-X5ZOS5(XGQG-_ETH5_1:&g,OV0Lb:/#DM?W\c+51d,RUUAfVMPUU
G2F8d2f/L6(SCdR,XKG:-SdZADS0g+FLKe4E^PZ3,#\)@GY-(T5N>>1EDg^g37<N
LcZEf#CB&aAD_3=?I2W?Sc2QcCML:N0N6\f,NB#Q<.@W+EAP^[-Y>[?f9MJPB8Z^
Ca;/G@QQ]Uba<37VP2>Z3e9;+I/C-eZ\)&^:;<^A0OTFF?CC6VEHBN-cGEWI]Z:g
T?eEGTfQdK<5c6([A3gGF;D6=XAU_@7I[2YPa-]JcEPCLLN\VS-Eg/=L;5fI9_:V
?X3:^5K7ec2EY<,)eX7W+;1G1H/EI_9[Z>;S7KKE<^>L/>a3d)8KQ6ZLRN7<A@BP
>>GU^Q1E00e/g_&UFI/V.L([^42B<OUgEI:50HKb>GHS&O04Z?E8=BGH>M543G30
G=#<95cW0ANbEdb^d4.A2f>H#JSAdRRL_64;_>:7_.Z0)\-H=;c98>_e5EBT\I;^
I;[Z9Bb^<3C>DV.7@4XS)\PXU20f#9dF\@)c[gdD_BH>ETX0=X:0OD\/GIQ[_]80
MFO-^5WY.R(&<fCMf9,/);&\<H+]-JI]?GA6\g^:;:#C]U6K>MHNHg/_#;-eGG=9
Jg7Idg]O4/,cBfHCYEN.A3)<^I#4::cW?RUPF@:MW1aGUV;2_WT=77)cfA1#1#U>
g+cgNTYWd\9(_/AR>g;&fQ5K2N2U>#J^IP^]O,42,O/S46KA?]Ra?W/gS;V?8d0[
U<-eK:)0?RZP,?+f3^-aFeJb.[B-fE.X&&FFR8H@V4]Y]/HYWX)0a#P78#5:cP_4
M_5\Rff.OXQfXS3c78-/S1_7,G0U.KM5\beW;FMfI-XU7<DBb^+VX\5]f_#V>(Ab
LAOZKBBFcXb#BV#7NbV;B/T/e_Y>#D^gVb]0gS;<Z?V4/;GJSKEB1YM&.R^Wc8#U
FNg0);_dTGdcVI/(5;BUX?3Z9E>VNM#U,]I?YNaB)@>23>W6g+T?(;Y#&3N^ZT1^
4[0\2V<?[?J5K9?_Z48Q/UefS5Y@Ie/Q4[4e8C:=cN<W8IV/d<.<MA#O5:Ige&IN
5HW1=)>4X>[_#PAF1e;9CbU81adE];?Ib5Z]UH6-0<L;e=IM&AZd5]@&NL+D,KEY
:&8X(VY]>ffa<]de9e^4L@LU_S0@g:_9==:5>:G:KHP>U[)4D.HO>[6/\H>F<[K,
6MQd)S=YaW4b.2NK@Y#@e8+H4X\H_RR6-TdCGf1B@5OANfH5,LV@CbcKX,=Z4I47
J);G8ITef,2;DEMLVbIbPG^+SX#6U)a@<2>?Zg2/Le<f<.2bdT^HU64F4Ga4@bUI
(N5\-JZ()SdL\,FTZF#I4B8^3?SVdbZX]K8bRJ?<a[TU0SMJ-\VHQb(+&.SSUB9f
B>F\V)]V+..M)-<[ea>^g^<SXNIfVb4)H;:Fg/=2-O?[=2.b;TgJ^IFGYUSXC1<O
#PK9a?Z\d<GR/+3V6cF.V4UbD]+S/E)eQG(JWJCfORQR@TRT=f@6;01^cN=RM5(S
NXH)?784YFF[6_aXJZQ:=QOa[C<3\P#TLJY/9H9<KQ\+A3ZeC9#1#Z+M\^HI#8R_
PF.Z26]Q&NIP/&30PcB8Adag@P#^LD;//_\1aKIgRcRce,::Q1cE6Dad5_09K9HI
a,ZKN+0/c2P_@D?-5HVW9[a(Q<R,N;2:G1BK0[fga;OBOEA<,AH]6,1-eQ#]SHY\
@-\cIKGceG@B#K33AT8C=(_f+VXfH5OL(Y,J:WWa&1;9-_a>#(PN09c6/VdTQQ6U
PW_fSVPKMIK4LR5O3>U+Tc+5S^_K_#Uf<M(<5aZcW?F,A&e;:L+=71+PU]WKE2Q+
._+VSYTKdJ[EC&()F\^MA4_GMeVd&XY2R5;UFK4R&O[W,Mc+[/b4]WaC=&9JO+d<
(W2V_<?8\OOO4bI/+1:U6Ye<W=K5cXT.SPY&OgR7=X.424&c=(P]bOO&D7&0T66#
5D8\@XWDH(R4KCg4?-7^6O>#SHU,7OY6\\YG4,(B[-<6.5CD]dW+,S-?3YJg@?10
44Waf(=3XL(b6V,LJM[7O+DKKLIS-3S6D9E];@UUY[</bYQ^a#bN.;70DR_D=0EH
f5?Fb,;W8D6X.JLG;;(_,Z@)afe\aN/3T[U\K72Ge9^O7E>5:J]Q;bT)6+G5)a_X
U5ObP4/F3UC21Wa#_=8:X9IO-UaAS/gXafOdZB2H\08L6FT#?f-Ze#JFF.0DPg<f
K6^IX-Og=&NV^Ja]J4DAE;gH0IH@HY\aV97FG=R?ZfQQ^A&+ZB&SQ]M(IP,\S/)/
Le\,@QEfB:FW_Kf9@Q.,+?;Lb8@5CN\:\F0ZX;5:4CD9<>g5R?<::M@X-K1UVLTH
Y#Nf6?J+02G1WD(2>;T4TZS+bR&7TQSf=VLY3&LC)88Fe_]PW1_;S4DQB@#9bGO2
4=-3:UPHT1)LaeJ+dQ4]Ed7-^:C[;&8cT.GM-VMWSXBZ9d5Y\ZeYFOSX&N]M\;>I
4B6<:Y7#621W@IIP;g?;K5Z.;C40H@R/KV_Id9.a8XgE#:D(C#TZ>:FRF8KfB?5G
^Y>:g&D9@Mbg:\>#)2N6UF=)g&1Rb_>cKbFa;F7Ja=AZ_<RNG_fRa2Rfb3e_3(EH
U5^f_3S7&.f4MS)NbD)a;KQU?[@CUK5HKa2WdH2HG^4gQg9^<R:PGL>0N>gdW6CP
&\6NK@/?M>]S@W3Z=PAMS9]>I=XY_c?Z]gCIcg1+,D18<5HFCd4K,1e9A?,:4;U>
+MIX[[_^0aZ?#<c?]C:.-SL/SQcG1@C@GYGOPCECEYS;4E0B[Q5SV+U8)Ce?19b7
dB9gI589#MK>X,29AYcQG>dYG>41ePg;//VH&5A[MAIEfY3?>?&g>:O2SFK6F7V>
KN,:g9FL]H0#PO()52eSJOJNf1RJ[8I?T<a+^:BAAg<5#gMdc.KFL4W_JTT@\T3#
2E->/1d@#H?6[e7IbIB0ea.I(2S<B/4;D..(?BGgf8e7PQ:QD]/F>PY]UfE\fYX5
OE\eH&3U8F,KWXH0U^TOF1,^VCa.JBaHL^,[A1A?O/EB+U,#aYGfF,g+S^JK6,),
:.#g3)-_<[T1S87/dAg/928-_9A<R=GHG;KANS>:Yfg)Ke\GaGR2&0#F,Hc-NCRX
YTS);7:S#JS8NYJOd0V9->)S[W77(Q+6(-.A#44)RY39@P3DTFB#3?Q63fWf<,(@
VO59+g9BDQR6\;7N&7ASe2OA_.J>0Yf49MA9F2>ASJQJX52,<E@N<HBZA^M=:RQ6
DAEVYA:#^II>M5C(#AE::HC?#d.:NZ,G;5eGH+QEaf4dD@B1QdPSLL,UaQW7,VKb
24.#d/BY#a8NaL@MC6fUS2)4).BF)L:-K\@;eY9TU3T_d,cY@Y=JWc\c,([[22fV
Cd=EB#:VLNY8C5R.E(T8.I]UIe)(;1MUDRIU7]N@&NEXM)AI]24G>&AfTQ\H\]@[
^K>__;f@RED3KH:ZIeK1\d(9O,g&Sd(OcHNC,Ue?4VZ1aJ_ONS/O\,+<,aS)1M5c
L16/ZC2edf.^13VMC)[PY//N+K\Cc(D?X54V(LAX/X,2B[FEfd&[-G3CY2F/?M,g
VZFeVfD\=b.S>T5=XLC(?S5>+[BJBfD6-?^Y+^_N=Td.O/6\3A.J?1.af\QV@]:.
2W.O]KQQ-,KXLdfg=^80f>13U5&Q,)J[7\A[BVQLXR05-)KHYY/[19X_5X@2;S+1
@Vc;FF+#b\=f]BL@.<e-ZQQRL3WT3R]L1PIc7P1RRF-_1(]U4S\(G=NHB27#U/Y3
c]f@=1J<+.K/L90Z?Q//=T.b.QZGIOHU>J,,NO0JY;SW3N,\4OO^#4WW.R70>Q?#
5ZZC>Y/^;_LT+;<YR42N;RTcY@VGX0_7PCO/Y-11a(5T9JR2U9fXG9(YH;I&:QE,
#162A)2^<GEJK(=;cNb/MS_380],?a:BKL#C?YRYAXebTc\5^:0Ig8JMd[\IJL&R
1[2[(/NIK_TI5DHed6@(,3_?>1&(YF7(8]/O[<afRQFSff<=O9=JgL1RV>E_0(RZ
2^-Ua3ICg8C]-1[98]9U8_&6f)F#YZQbG:Ue.@R>gW#O@8:+[4[F9&J\D^3I]<PL
d[Y3X^>I&<7?=0G^]CURcJ2=cUJ6T]DfI9L]:GT+&)Z,ZF]a6:B6?H3PSWCa?UC)
7\S4,,PQfAg_d1bS-a7,W7ffedX;I#Kf>Vg8BKZb_4]1MD/f;R-\SVMAK_-]H?3@
QJgDd>)+?dQ:RQM^/##fe3R[5TRO./bVeg>#LG6[P+?d<-\;Fa][Z&5cPG]PB4()
=CE;cN?eMWGCPQ(#/.,4R,+ZeJD9R:,?:c3K,Kg\S[d+,eaDJO@?2cW#,4Y;&,(:
][58/LPa9^c+5D[B5I;\+80e:1P-E0=L0e-1IZJ92=:2Q)^_04&ALW>WG5He&KEX
SbHf?1ITeQcBSB7#=e66^-D0_^[L=&KZe&Wc-X7Rb9_/<:O>52_&DJ4?&D)WZ(Gg
e<JgbX>2JUL9/TD,5afdd<MV9Z)]XT69PN,BF4g:PQA<]VT2<&9/_#_8>G)X]9[=
UAL&2#Z86P:8X0CN_R9XCB/SL+M:)>eFg/7fP\YD?1YDH_-9&<I++^1P7EWGWDXT
g,5\E@G@&YJ#I]162-./b=BYX-U@2NBJ^f9ID>@^7eM\c:F6_?XY(;Qff4MQb[cd
ef=1ZY3[N@ZMQ192YQbBNcVW27]]8b^;9BV4_G60FAO<cM<-3.K>c5OP/DPGQ_95
Y9;Be-JY?/WI&TJT=fDC1dGJNWORbF,M,/b?Da;JS8IFeYDF28e>9-GN?<P&Z1fA
d4]L1d2Lf#a8@-0NR/N,)M)+CLN,@gO=Fd-MST_c^3QadHI7^<A_A-dYG@Tb72O6
PadV65574F3cIR)>6aPNa:V9DFf0=2-e/<e@]_C+NC]18FWLZG1,BUQfYLRHV-_G
N_RZ&5<I[:KBb28E/;F:;Z(R0P6]V>bH@<#eR#B(/Taf_(g7N5M<#:5]\PCR6Aec
I0TUY&^5GJ)e,,7SY>VS>4fO?P3VCLW9]T>+d8=8@a3/I_BH:6?85?AM[,#Gf)])
(S3>T?P,6QDR5P[7=@3fe/T_X\C0,fGB4PL/L2dB@:0Ib11&E.6EfV5=/&#aU_&U
NR1WA;W2@Z0==eWH_UT=.R[bHE(/B@fL&[2JRJ4YG+L#]#1?FV9VDXK;&B/NH:G8
#]JE</6>]?G#H??\CQVg_Z8=GJE)[/-ceM#CeR5U,PK;U=OIDGIQPH8/fWg>f\I6
aC[^W#V<O]PXQ68/UKa>^g13BF5]=_YS4+SbG0.12[bQ;C\H@SUU:K7I5=^8NB21
&00J7/4RSC&aF_Mg7#5_Z5Q7V@\-+I<@TI-]JEQ8D5[&P(6/N_g9TV:/BdC9E6[C
WgI.d;QE11?Fa_XOE:F\fV0.ePIK/=Z52_B8=I1G>#4RQ)31P&5OI31ab2d0,a8(
1a<1_G;IQG91LJ&K;(/gDBC0&QBVE]_A\@I3>ZW,BFMRVKLC>8WEc0]I>T18facd
AZ[U10.Yf>49>QO5F_ZVQ7QWM[#PUYEfZ<]#gJPY[-^1T9FMH1BH)^K<^9__^X;S
O9V#BLKPU)dOb?R)5F3ggZ;.AHb?7XEP=UOfUGPI_DdS6WGA4DFSV_e7UVQK4fU:
;W&6LJ[E,9;?LCRAgO<?+LC2L,-CEA[\IZ_A7C#KfB#WU-742[Oa_.Q73-b;?Vfb
\ZL2&O^HLYb_[SLH5NN_RQ(SBU=[X_T8bX?>E:&-TbdK\>J.[<9D=L2(R1:<8?_6
P51]BR+]P(b\?,C,#8Z5E#;J8CZZN0_(N\TXOb#IV5Q5bT228A9:PXG=9D[4U)/R
5\b#ceM\dfe\24V][BU6EYZ]^N(N-NT3?<ZG,a>]^])@Q0EdA/(#M@A>D@);F70=
LT_))TB<7&)fa39#8<c3\.W^CW]Ib]c:PZ6fGWT<4J^9R:-B/[9//<^(>dV:<0)c
Ug/5#gX;KL5\?Vd&>5P5??V,JE&07_2bC)cM:YX&40US#1W4KTS_+3d<D8:5B5\3
8LfS:b/X6@F-59(SAFg_.K5A:[aKMQK[Ugf&A9]XSL&UXPf99@aJe>FMEeP&&fY@
^5f(:R(aJ,NCUQg[IS;0Z#B0AdLFQeDMcF7=X]-S=e]MA(WGGB70:_L(D;fEP/41
4a,0@VDG-6UdJO_PW:<1.-N^/ed&T&?Vb:0IEcZI7E(=CNg.[8VMb)[E(;6QIAW/
3S?cHDK+F]7,RF/FJX.Z^YO&c2[=82XH;_X+O-\4]Ab&;M-XcHFcMAd[e7R#9<-L
Vf-9J0FT8]?_YHW64BIH-;Q,fdDd=QbDg;]_;@aZ_eG/AN\W_+Q2.,gH1;53\4_b
&WD[YfVP/UdYEPBTU<f+YZ/JPE0b3\&):]9FG_DTdSRdHVOX;-E,&:e:bNR?+Y[=
FQ]:;]McLeFFC+PBOJc-D\P.Cb,@FaT?b:2K-OPNQV2(gIaI@V[OY.fV_>\/CG\L
c<[5\.=E;gS-W+4,N80=M2P\L_RMc7-37^[5=4C7M6/U(^5:_JG21R=C77#^cX<]
GLL+ETCT<=0]]2@()BJf:ec[^2.[;aH=IgZ]ggHG/3P^E9NDKZDQL)1.IFZ-5N(D
@T=2cWG:5#I[,H<fV)]>/SKA&()DFbcF#_TGOK?/?&X7?S[@2>CNTP7U]GO>=7Fg
SV6Kda9Y)\D\F6e=1Y:V)#_I#.<cC.B(8Qe[F;U^(?GJM>LE=P7/)>RA.<(X\O]L
9U^8JgR-aPMI+)_b35?G??Xf-d/O)8\fcgd,7R\feZ;FRKSN#=8]QVHVaU-B1/2+
]P7b<()JPI,RHQO-Ff/1+S4a:>[(b9?MVKa))-Mfa[+;cXAXPT,7O_9KLI11H);O
XI6b&N\?2LT:M0AF\2A&K4b5\=?DR,0a:^OAS;PJg(1N?F3MLCE#W;3gF&,QP8bO
;O<@bF&HCJ7a.>4e_3,[4JY(ND_/]6B.VH/F?3IT]SY1(X\(_BH:S-F:)U+[3U@+
)/ZeW+[2<XT7I&<c\<faefZP,0K7^cXISHI,^+4:KDQ^F=EK7.C2e1U-)5<BVVc2
IT#?F6@EHM(d^E+3IMNH@NaQBIK\QDU@7Gb,)dDVIcBS\GWMR\Z_Y9B7cZ?5@6VL
c1-Ee)>=Q]0DF9]D-#\R38124N,5#B;AM_[@43]V0;&.L&??A6M1eI5Ud1_QdW&F
O?/Uc8.D:1O@.eV6af@PBg^]aB763C;?A3+D3a8T[R,?#?5Sb5\UVXRa@->],g8T
GU^#Hb8aPAg4K9;29P(2STRf:?5]3R_;@eHUD36-EP6^A&1Q<=VFGMF0[HQ^?;8(
X:+f;W=aH(9&;4M(UCV3@CN##G?K7/=5^AR8TbH6:5,ZA18@?:C.&EU45^Z=gEF=
UO+J9-)H&3d;g<D_E)R_=SD2G&T]SC)=SAW)=O+b2\d_=L:J?1^+V[YZL/bS4fAF
))?35SWA(J&#Q,aVKYI3E1)&&4BW=UNAXdJL9V)1C;FE?1HX>.e&/\,A6@c5)(H&
CgZ)d+T0EgD#6[J[d^U+;Z-IeW1+8#&c562:S?J,40>e0XJR]gI&[1:E]G^NOH]W
ADd;>48E8bDT;XbW,e,ZN@CLITXW);ZVX&Ge._P]d.ba4L5)>]g1&=0Ya_;2I<f5
g;U>KGW9e]df1(44T57?7MVLd863Y^?-H>4Z[P:4_UfQ_I?5_I14;<4::#X@Gebg
gM]Y-2#SUPcJOfDOTR52B\ITf]#=4N+C[.-4gSO4Z=cMN.C84-4_-G+Lf].DMdVe
e:WNZTJHCT>Pd3d2e;<QB8>Y-?CAEUf6C928@,_RR61+>XX]?g]S[af[(X[>[.QY
^Fdg_gQ5cKJG(1.GCO[ecI1BS_:UB)E=YR_>f/T?RF0@@0#e91LK5@?3,NLOPff4
_M07TSEYC/7-Y(4\\aNeATQ5WO(8AVga(H)SNG4D2Nd)HFCec52NGMTMQ1<;c.=?
^C.>[FU7LOA=BAed@c@-GX:)<LRFL5g?5:dBU:(D>KY?O=V^SCHG.SF+&ec,d,T2
G^Ee=,LbB^9D[9._V(DQ)NaDaLW[4>D?Y5EEP=9H;H2XILBVYX[C75DOMIW=<SE?
=c35[-_XVf_dM6D:4dcKdDMC5:T865XeX^V&:8,@d+&c?\3QZH^a7Jc0Zf.T[_H+
?QP.)>XY0#eH4\6<Fe?e1HCHW@8G@[]X)LXY/9g7GA_/+.N(g?.;-BL@,Z<CLYUN
bOCNM>TFc#V3:F?b.)]/DB<gfa]1ELbFW#e^DaV>3bAH6@;@FcO]KD1K@FQV7N58
+&E=edEXD1#B,(\2DA8>I/a>;+DJ@&gDJZTDTQBA?C)K8@TKe4EK:BaaEB[^#Cb(
&(M\PIXE#Q-][F>]):^RQGJDLW?T99LDIPDV]c>#XKOcQ/::6Xg3)&^1e2MdVfeS
,D7OdZf)FJ;2K-)2dSNVO:W&(^1=V8=01ETIZW\D@^4,31P5O()Sg=[=6/N6E&1X
4#1[ZXGfE^<^2Y/<6AAY]PcCFTgE@Ab>T=2YQ:^47Z<J+VC>f=Q\DH)R[,5[_5;T
D8>1c8P,?\_0B&#0g3;_2IO.0gdK[Od1TTSa\QL420P+46Q+\;K_Z>eO3\X;U2G?
(&IWN)N,VI;)Kfb9?B:E8/L6NWBdd,6YL>JX3USb,,e]7aU2KFTBQK+g;&cG._&>
72]LBGY=58dYSV8UI_Z@@4D[VY:-X\0^F#^Q;6.g]5M<#ID/M+W)3O2M9[T>RPF.
468HR\?O#)IQT>:>+.P>C7=-I0R+@4QPTDVGVZVca##GM#^L]XO.3,ZEUF2ff(NQ
&<<3c124@d\bQ-?2Y\]+\RU^2TC_G0E:_V1KQ/-21Ef2>X83bfGGG(-g>AfP]TYP
20Y+S;41#JggW8]@[_J3_#&D(3@AeS_+4&=:XfeY4gEYe1:N>W0;S:P>fN2RcCLQ
3Kf7U/YVF4_F6,;-:#UR?bSAKBAbPTXcC4.6C)_cdW_5[c+_&@THA[WIWX,g9W\(
DW87X5PF5YZX8?PCZHDNU(Z7LI^A.XXaag#KU4)g?,9^Z69S?/&X1HU=.fEa2X:P
#/1D@7X>NI0NW\KP?+g\=da+W(@O00b?E)MAH4B2HdFBS)]2-@R?];1_41Z9(:\I
HP9+R(;<Q)PW^]S0Uc8WRGZ=+G9NY9KdEOBA0L<T=gD+]AG#O;QMafIa@&\1g>07
B3:=X6A.1-gW#XcQ=SMa5O=]bO_94<4g,J_0=4W.[-\:0<1dPWefX#f,DPHQ2EFF
Q^SY#&,AObI,F?)C@&IfdEVcE_B:;AWGBCP-?,Pf20JW(UcX,NE/&g-P)+^cHLTe
c:IAZE7a?ac2T]1MOEQ8,dA^\J9g<FGD)GVO1<5+PBf&O^eMAP^e_-.Qa5=Hb4)E
cI5eVF;9=@5\S2bVbAe-8<76ER&HWaC4#ZDYD_]\<@[HLcJQ;H1Y8B6R0))(GZ>V
Z/N>I4NAWT#SL[e[b1f0,VVge0W=0c1IXAA1)2,3]?.09M=0aKWRG#>U<e)FYcVM
\O4=P<O>/Q>;Z;&W<2#3-HS@Q156P=_D@-)_3E-1eOQE?a,4dZB5+,G.F=?0=MFB
-Sg=CUB)3QB5a&I;@\F22cC/bE2b>](C@;I\2WX?6;I]gHd/Z]TY3KUNI6gZd2D<
OKUNb@b6RaF#C.G?LUU?[)d^VD>.DAYSI^5B;YEac4GT^..W4=)^<2)dbV:E,D;Q
S]K;7B^DDLaOPP&0&SC)[=#QYUWLETKGU1J@193g1ZR3NgeWG<?d)N1#LBL=Wb(+
=+_VH+EY0\B.FVe[JKG]^NCO,;F-_R0DH7f_UXe8-\fYg_/?3Ac;T6AI>ZXeA]04
N;Q6PM-ggIG;\c;K+M]^?/dTHN,8JSZg558Ea(aD+Xc\c)C6I>cR[,F+,:=PZ630
;JFK_d>3K7e_:JZQ,-DZ=ETKTH-^.d1E6c^49\A6C13<5e]fTaQeRB-(2(&J-@&C
93TT11;^,TVRKUEGN:d6eKWb6NZ[0a)/UHN:Pb<2Z5^)=+7eIE6a=/7;8?(,IQW9
@CTUg-4A8-eMP1;X@.-[75^BgX-BXY?6fa0TVCCb5R0Q-@g\,7CU8#?IW=>6#J\a
M1P#ZY3[YX\:-)#/6(IQHV7IK=3eKT1(4Z,T?=/PW6=U/aHbP.7QSb4@1bL6^H)&
V6<MgMTL^DY1#U;/92aK;,?I]<<+fYT.a(gd5ML6f<RQ<2=b(I+(9^2\>ZD/aV[B
]eERdI=6cZ#dX<JdIN6,JNI?d9-:g41D33]ACOT4_((_E.SL(,O.d7dTWf6H7<G6
E[#aRT^3V,\7NFdHPHZ;&Ob]+]SX3RXXLScB2&R_Z2-c/Fe>^[f^eK1dIM?76g[7
CL,U2Z(6WAKJYf&FA?6HgG7,S_/e_10gMS?Fc-,SQNFX60/8\d_BJH0()4[O90#e
QNLdf[9V.1Z2eDT>,/?70\(PV[4.dA.[e2KELIB2)9<aI:PX;3\IZ5HH)L6VEU(O
@IUM?1dB?/[c[#>IDCYZ\N[GL4@X&Y#&]T>XNQSc=GZ7bS-9MIBRNGZWIfQ1#M+H
)YI.>Sf\KR+)PeKU[9@gf#?YUG=\YfMND_@GN<d2.gAL_:OW8aR)D[ADG)3V?3P]
Vb&;c;?00>3UG_8^=-YCe+N.\D<?6O[/fT0A;Fg,3&NdYDPRUB)([Y8)L[9=<=2A
8Eda:>#=E(Q:(19bDVMeX21]GYX&N7/9K+,P9Ee24FB6-dHIW>F/;G79N[E_YO=C
Y=9<6\g,QR/1VK?eRLa>e8R]UHH./)M\\=d);-=LGEMCC.E#2gU-_DP.NB?WJ-@N
=YdB7NU[OEJ/1ZQ)AHb1#6IT&HW6N82=ALCK&AW]Ie+#>5SAbN:XX1a[5QRagVX6
AA&04af&6D&MbM^<.=DfESREZ-42XH=##O+6b1VUa?V,D]5[@@QGVB_IK3;Qg7]]
O/?S:J89B#aDDSSa<3U]<>bW>Nd-6&e+@PT_=V7,Wf1/VG+P&R&f\:>)4,M)f3,0
T-T\JZ;e1@UM&P?PI^.X3UJAL:U-ZAZb7+a6=M&RB8cEGeSK;^Hg0L(JVb;TW,:\
_,2Aa7gE+37E\=1g2Z-.TTI0+JR,/1.T5PGFYc<5XS2c@c_D^B4ACA3B-QPZZ/&6
eF+WPW)DO\-?>@<]R3/,;P0N5#d?5TRG]Q44]1;5X)1/I7]cL5_-F8;:X]HD>;[;
..([L.PE>.UfR>>>CO#FQcO3]XNICBd\N,If?Vb&\fK2aR0+HTKJVYH)CI-]U#]-
c&Ae5^8R\g3I=2RPcSK2W;^MQ9ZS[2(2]HO/B3^e=g@GFX:>_Ua(bX]&N]^Sd0E7
ZQ;^KgE0DTE9V31N\=RfcSMSgM?(\MXgKPGGY07f<44]OA/N6B/M_@\>N:O,3^FT
?@1,V?MY5bBdX=NRHSN]da3RN-QL_e=C3V2.;BH03[6-]SADdUU#YLGY(_)PXMFD
^OQ0dXgQX4D^#e3d:,X,FK&T,SdHcb:A)UCBd>dKFE/H09&:W&UEQ0d6ENXP]0Y@
M3RQTK(5Rd,aY//FRb,D\IQO5=TU6:TJ&b6#cP=X(I+23+G0,D65=/VPTWV3IUKE
2(@FDdB.A(V\GB]_/\Y:K2^(b22ZIFbZd+&:4egJTbO;gG1E-K(LKea+R2@1M)S)
T0&WQ^SH]JP5YJ78DP-fNH..6:<EBV\Q9X781JEa#eb^[G@eN<V-e=:-]D2XXW18
a0W5P<,e(0LaFGLg>CF,CGWf>&RC(d?DFZIcd]c(?RLXFMLHY#YLc7(2;6-NZ9(A
--1:03]0[gaTBe<PAb#CLf_W.SXFEf9eR9d+]3[LDVM51e#RRdXZ1Q]Lf/>NXQD<
94AQ\E;:V5+U?FGZZ<VKGX=<9[eG9bg?\baIdEV>/[a&b(B2f)<E5bddN2H,SZd[
U?@bJC&@@VSMcO.?HA,JT<-Z4U)XDG&a.Dbg#3=_8;21(0c@6^)a.(&#;EOS<2.E
]3cO+KQ:CSJXF/)EU4CgD(6Kf405aF9R];R/X02W@&^fGcS8#1&EZcB>P;3gOWTb
X3H,RU:L),,&0U)./d1_6ISHD.KNgO3?=2\a_-\-6<Ha,cHfVTNXR9<UX<a2aC0V
.UPR@V>fFXVED(7d0O9D2#2ae2?cF\I3#MX\>0c4CA_=;d#4RJ1G@L.H#UU711Q;
FZQ]Jg_eZa3,V8QNI/&WK@+1<EF,S#::KXGC24(+1G?G:-2^#AMFHV3gA,eA0][T
0>/H-C1VU;96F90;^R7YS/QXC8);e\0QI&dPf>g.ea8)^L]<)3/\WE6^4[VC>F6/
>8cG/X4(<JYP3L(DX0PdUd[:He3Y+NDT>]Z@d5W?d9eIN/PbO=>ZM[YgM_AMAf,6
eV_@L-4-VGT5.;#FD)O1U0^I2G7>L<?_YW9;&b_]Y/Xafd1#R97VTZ/5MZfNBS:H
:]Ie1F<:e)RbCZOQVQ(+a<)G1>0COdS&;C2<2\MXcL[1D)e?_[-[XRK<)/5]3\bT
V4R:WVfK0>L@9TLWfFZR:PF9H:E^1CRZaTH,OY>f8]Bc]-Z4Uf1XQX7\6Ne;M97c
U_7\]WNA#:--_ALBb<IU54CUFQE_BC(>WRP+ACGUAg0_Xc3P]>VBU0J.I_#JZM_;
W:945K0J+>5AT61=+GSfN[]Cdb;RM#TS;@E8\CK5RQ@cBAH;Y3-MBLS?e#G_._WP
(Q:&QLc32@-:>F1:U?(YX9(>D0PSA;^-TCHBF;F#BTLWfHW31WN.CG7-V-?O7[H=
X/D9aD0@[F@N=I-M,UN#Y,<<,-JfC2LVF<T[XH6W1)/O2B?<+cC=cAegI]A6,(QN
UQTOg:1<GHSCgd7Za3H2.=Vf6[-gC]HNS0f]>5\X--fYU3XE[CR8ZB>]UDOM5Kg>
JGM,,b]C4(D-FK0T-D_:SYFJ6/CPYPZcgUHQe3V,T:JD[5TJ^81e0?@e4A^M<;?-
-f,J(.J;KA8.Z4eVcAa,^0N7_WP2fYKN94O1<TYgWf^UGeVaA&I;.7U7=>[FaZQ^
274SJF(/[;@I4RT&U?B5KP,Zf-O[N6[>2;C27KgQ5Y)gKf)14-8<1@f@P[dDa#03
7e9J[0DMYNc.f5O_+D2U6G>23U,[CTQO0fCOHIdfWeIFDWQQ26/a?dWR]gNQc1I\
?BCLBWZ7cJ&-5@NII94TMWYeD4>e@7b@968)eH)8YRR>I#8L>F3\-(c=M5RVDb9N
2LK\+KW.,L,)_6)c+a.aASV&Y&&WbE9Ug5]De@;ZDRM.0_<Y(6b4fe=gS<EA4[4G
1Y>L9?<b?V5?+a]f-DZEJ,8HAR9?LEa].H/C>9HgTUN3PA#K=RS?@X:L#?;JY(?1
6(:^^\=Y&O/b_OF(B7\B0W@AECN70eM(W4K&S763V#B(53_V4dacWGA=++MM\U/Z
7Fd5c)Z<bD_YePKF,7-LSH=[g5a.JgLaM7]d2e<->Q/GB.T#W9[L4N\HJKC@]>QY
#PVN4M1eLE0dVX(8;NOeC7#bI#5(.]K,3=DVL(0fCQ1SfV&U#UQf7H/+;#K4:-R_
9FJDKG)M;-F:e[#]_/&<M#a?1ZXa.L#JcB+aWF7E+fI0WM4d<2b3Y&7RV:SL&SHH
\.+N,;LE\,8NJ5aWB]@d_[+NDNNEMQ7>?.8aO0G#4G1E:&S)G-c/d9e-AH?65+LO
[.E#e4DSOHcPXd1J67.M@U0?O-++,A)[^YaFXfd;V2&?\\<Xb<[H;]Paf85OV#;,
Z8&3Z[^O4ZeI&A.12gWRCSR^8,M.f70(NZKF=WQ4/=Y^_TOL.X)Oe/cSKRNZ,2WW
WH&Vg+NOGZ24EJe@?B0:]=I;&M.aBFI/Bb9c2WG8fX).JdWD.AC<aCOFK(A2bM)b
EH7Q.VbXC:2NQ+<3\\I_R,)=W4cRBNTbb+@14C,L<8/Q-NYFO&5:OOZ_9Q,(WOW]
a>1FRI;G[#]TGMOO0Y;I=]\VG./XACbO>7;(de+5WgOFJREaMA3ADF;?cNTIAc:R
,7#G/#IY-gI;d8P,3(3XWRI.A2Y9fTF1.DEP9Td6-_)FR_P#P-TJG4&I8Wg,W?X;
M4FA8A8FXRM]@D^CafHZ_[.:DQJ0+=)E&L<)TK@W,SJLaf+]>H]/(N2QEgN.W783
]b0(#KR3,E3,d--3>V8:17gU-/A4Y/_AN8F/PUeP0((0.E:6UN1B#Hc8YA.DGCgg
)E,AT/;RN8(6[3eIEa[-)#F3SGBe^)AZE7G8]8bZ.g;W&ZgQaf3Kf<L8LZZY/^Xc
[8<dVNW,aE19)eZ23J885X_@1P]XK\?DQGJGaUT&#BDdf6E\P6=?;UV:Y3:Y9C;E
&C9AJAGfSIM[c68E0e(?7,0AX)?<=0d(eaa&I.=S#2-Y3R#?2S=]5CAQ\(fc@JY#
2J:4^TNF6fFG(F^#D:AM;fbW3PTNB9+7GY84<UVIZ&6>L@R+eeK;.+JXZa\3:@DF
8([C27a7IK[J/E0,f[/7=_Y\gH2AF3]W-QCEa\X0LB9Z1SI+-JGI+M<H;0P?[f,7
O_S^3:\XKWPC8_GE@9c3aU/M>+:4Ng\;=F(gQ(C:RA]:FGdOMIc<(Ob0a&P^/E9g
VG+T2##R#?OJb2-6)0b;CSINXN_FC7cc+JG@Z_XL/[OPH66MRK.ZP(SZcgY@@8bE
SN,OA6d]GK_1V.\O3_2P>T(ZFSD2/8d8DLI_f?6A]/3:AF@B33TUF(\Ha4Q(BGBH
:PY0UQg6.&RKfBB-7D+e]64@F2PD.ZD9V\=1,OaAZaIP+V(U25cQ7fY-PJ5BD6L7
6NPO<8JU((bQ74\585?@\OBb<3Y>CRM:-=^=a\7QRD2XP#F7?b]UDLe/M=M>-W73
=4bKcJJa-#L7C,7\X,#R2e7RX.M0Lg3GR/1^M?T<ID74>>f&.W3\NR[gb[gb9BcA
&gR(dE,#N,/>.L)SJA\U3R^,ad##U6UML[@QWHL(,/U12>A_eUFA2&@gVbUecV<+
5@KCQ7#?C\B#Q=Y1CO@WHaa4H7-6=P9+VP_#B.H?FSQW0D/IA82f]-4:7PT-MaA4
\;3ANSa\I8A7<g>Fc_6_M1#NLTaD0M>U6C:?cg?QfQ#M3d1?JFLa5(<dd)VF.I98
9gP/SF>\?dKW+L?f\L1ZZ&/NFO/42+=HNQ;5&+V8B<N=^R6:6d(CGJUK?&K<B,g.
eD[56B=[.g[.+DgdULWNd/TL[c(M4R(]83&5Q_6\S<\3QDg_H=&-.8DfebF-5-.L
GJ,Q7MVEBg+F5D5YSWAcKC;AG=.7QW6-H02FU>6U9E)SGY94Lde#LKC7LD1gDX/)
MbV9/FCC^F&F<?]LBZ47.U,[dX9-I^b9.gYG2/egVG@M6C78W9VTC]F9RF#Qf[N.
1bMJc5DYYBX?>/7(E-U+:8+Bb1@XWEHF#e1\<3.L(e/f:7GEK##c==ET@TC8]IV<
IG0@G8d0.##?@Ag\:1>@1?WCRcZQ/dU03Nd,g3ge?^Ta604(-6K(4fD_E;ASCY8C
a:fEbgS85&H#cH\6R54(@UFb[;RXfVJ2YfbX),Q>>.cFPb[bePBdfc5.O)=FRa4#
BO=J2f=WLKb\Lb.FH&1420HV8XL:3f@H<=fb<^DKD1D[+R2D0Eb6U\,L6&2O;B(7
Xf;FSdPG:W&<4S>/+:IE7b3^;^OH@Z@G)(HQ^>Y_a6\_?LI]\,PQM#><\E@I2b6T
QBD76,#0J+N4ZXS^,9JM#a-Hc1XA>Ac46Kc_EJeW6;gV1MK+E@f#WUWLM454[-:+
K)HZ(3TE_06\=QP(@M1<OPLb=H_H)/;=TUPe.]IKKAf&AM9=9]N451YU0D4[]XYX
eBY62,L)]C=U9\8=f,-KY9RK2@-,Y=RI1McU(28(_Kc[dX-D>EW#FX^b\)M>.=Ug
S+^:?T+1FZ?8fI?5G3HY=+2ZKK:TLbfWHFHIVBE9MQM@eX\/E@,J0SeGW)KWB5L+
gd9bEI6:&:B0-R-EK/V+[GVKK]bM\/NU99(>B@AIL8,#-KJMK9b/D/\-H_?6KbgA
UZK?JZ37^de&O:B)W\Z^f5?TFf/0SUU7bGN;F1g/BgXS:]K49P^7J[I:c0-U2?3E
XAGD?<(4FM-G?g4U)E&Td32H9(fIW3#d678FQ(HbHO@[0W/@,N.RL]-8ff@,:CYE
0RK#K+S2>+B&MTW61A2?5+0>PR,GEM9TXC-3E0OG[B^2,a7WX//gUbVG[)XE5E.)
J2J/Y>aXVBH(,)<>NaG;T:e94?G0GGVbJSN;N=[&gb2]6a.MJ0ZQ7c)OMZcXe6WL
.S+S&#N<[S:#:RS]0b],T(UW,4<(XQ_&+8.G8/83d/G[dVXVRE&9a.>^Xa4ZSR):
C?0=c]6W7Q]I;O9^4G(Y?WH7PZG1)NYTAL(_1\1ef]KCV/Mg-@dG7>1DdaDg]4P<
J\^9\.?FDd1[;>NW/JNZC?[ZNNgVKPe+U]Z&@6_.G1<KOLVZ\?3NH0U\=fNENc6@
\)K.MF+S5e,PT@?g3LZLE<(==2H,08C_:K#XNY-O_MB]N@eFOb+K2PV60Ue;H\K-
/f</1M><BW1Ag(:(9/_X7ST\IEZUJdeSKOS_RQNQ75B6G[&//e34ZO0CGO-IFc;A
>fC3De;[ff/;M7FX(O@DBGD.9edJ2:+H;Y(:Vg\&^a^UDULPFZP;,&XT8^J55IN_
@XA8Q,\/@?QSf7Q\@#O\aG#RVT+E6c6MP6Q0e\gH]1)5HG;P:GZ60KVBSDNU29TQ
b2=BQ;H7^V=<a7#c;RUg7aI20-K7+.)?TT=FE9O<88Qd6JH,dM^3]&b9-Y,RVZ.C
WQg:2I\#&[,dT@.,M>@XO[A(/OGUKe0FELe0g;=>4bN;Z4X-gT^M>[E2;QAIF=gf
:I=K#A-\C?Led_JAAQb6/7+Je^Z867Pc>/Zd1YFdcK/WYTa#BNJLK;<Vb@:93:D4
0\=e)N5)CdL5Q9?\Cd1:VX>_@0G>6\-#MV\PTe-D/)]FP6X\\&GR3ZgNaL9U@UP:
GXa.QX,MgfbLe]@g3X,0Y,\A-W,b?^KP4^;,3@??g[EgUK<BA8DF;)N939J]-OJ[
M2/<GHUW+LQ5>N5XPRS1YV.gb-XUN-4ADFF2U,I8:[373R^TE\-[c=IU2d+JU^V6
S11X1<dUM>cJ)XB0CKM[PX]dG@PW:&fR.g)7VcBE^]SFI;S:40@f3Q<F\2Wb)4Z7
[3.SGR1,)HQ\>DQ;f5SF2IbD(?>T.4)NO_G).?;K<#7Z[J_MDUZAY1OZe1W4\D&B
X868#V(MBcQ?[0bTYb@^^;54BYLRGPY1;6HgAB?;EN.>O6HUQG,3.875TdYKD#>H
<YM\d(R_\96Y8ZQW4<P;-^CXRH[cgHCR:W]N@g1MDb_C]4\CSg-^)6CDIJb:4Y:/
PgQFZd]Y<K+[0C0Cf4XZWBgf+Y^&IVg7f3KR<bWR?E&_c@#?S3HDSMS_.^e;[SKe
b#+^.4JGG)#9)dZ/9:dL\D.#:5+9X..5RO)V41I^e&3eT(=#EV@eG^fR.4V1f1DZ
W=.+9B-2W(W\KMb5;093?#=T0_0[&g<<V2Vf1CNEa#T_5HV(.<[:_?NHNIX^bDVN
-OLdPb+0GHFWL<ObcN:1(D0D<:>RRF\F2g]GOdJc8)=>OJ@VE\0A\7J.V.^+A&.Y
0;M&N+.MZ432R54P9Z@;@U,QF&,,\c3gL&6[=LNaZ2_>bfWH8E+9)aAKI>8b-&DQ
A+S+Lc&Q)SOCJKOe@8f#::a##>ID+GOI2;c[.UL69_&.:A65@W^AG0C(:J.K@cCG
g3D__N][LTYbU+Y@6??O)bKW7>9Xe[D@7.Sc?5ZJ464<IX8.M,H#3L^g5WJLJQG\
c(W/HE87BQT(-GI6#?I2Ue8\]A@BK[JH\98(OL:2cXP?708TD<SDXMDCVbLM:BI5
T2OUGg-e732U?R?@)J8fbcK.]+A8[][-HFgTJM)_c><]+2YAFR-WX8ceE(KNZL\)
@]1)g/[7EDD][NGTKYJ+?-]7CSg1PYSO\6e[:a=S8BPa>OKg9+N[PTZB6b<17FUG
D9bb[2aeWg^ba/1&-=S<DTELG^XUb8KHFZH;[Yd,8[Ig#<G@0RLdC0S<0+7&L?4R
\C#@6+BgaE=-@#X=>&((NZ;4b3N-PY?DJ7AVfD^-13J3VE777/+Ag7Nd_?R#,MR\
O6L]/eHJ;Vb_&@G2ESa<67I&d:J?23.,^7])X/4-gZ^Te&EF[R)DQO3cNH2DGPD&
,;M@PS)aX8PW7eO)#c=6V^3I7:=e>ZD3XgIA=5&;;=Ua:W=D_+7TL&NY5Z+L(T/Y
#OH:9>=WVaFcNKM.VWH#VDA::B__X0>O4G=].DDH#;#:A/g0X;K?5-P^Q6GAXRG]
(NT@1GK;C68b3G^?NUa5;Y9DW0.;dXRHXBGUMSDQB3e+,.8=<<+c/Fa1<W1+PVVL
eZ&O\Q_M6?@aY:Y#I@bfVa+e1b=4bBK<f:?XaQFMJ^,#.)gU&,,MeKA/eVKVZeIJ
+&?2SVL@;8R0EO&RAaEM=P<g@L-0g;?Q-Y&]_^Fb1AdfccCR_YS]9(;XbV0f1>N=
,b03:O;[VaRe=XcG8]JT&=O/5;]J>&]fId^BG]76S642&R8efC=8U/ggFI6(Z6\X
?_L<[8O(ZA9<#]BFK)cA<<2?GGV6JJLDUR2cJ6K.U3YB[TgRd<P@K=dd@ZCQd&+/
@N.FGX<@&MDW<VV[76QTdHdAF1&@NUA5[5FY\@RV6)]R-<VK<T]D>7X=YVK,&C0f
S-<HAW,Q?5P35)+]2M^cCL>(24QE<]aP4cXL/7-WA,Ka(]J;<).<6b.3S28cdGG#
(&(De3^?)QJ\B#(<BbbX9c<aI8:)F+?JNV9M<af_F0CV>N5K=7f&DJ_VL09&1dae
],)BOHR41@@#[0fIHNJ3;ae8)1A5&WI5g2GV&+\)B]OP,YM)ac^O8,JTg&/;0EHO
Ce9M0E3d=WFMFB.,e)ReZ7E2&6_7T2&1d:c2U/&=<E>0Q2Qb>E?\JX2MPN/]b=X1
Rf?6EB5VM&44&]P.S=?O,@X^-<BEgT9a+ObYWTEb#<O7PdY<e>a1#/DM/\_1cFdF
JEbOBGbSVYL,^dE:@]+QF1[-N_Pc>71\H9/O<F9R[1J^29IJ0&gOcENJ.9WWSM,?
APZ(<=70gd+ZA76X/Gb3[JALQN(KJA.>C+dO>DPO+aF72,>]Q2OI]6W8<QCg:6?c
8BEXR).AFD8TNOWS)WPS>;][NW..JH>?3fLRLG.[g30U_Vd?]0I#+N]g9_1Fg=#\
:BXXZM5N+8NSB=:DHbU0?,_QdY?6-L?I5M<3f6H:W=]a8Tb_\>.[<G)3R4eJa(RZ
B8?.?-)Xd(QQ-B&ZUKFZ,=\^R,_7)C(UQ=(B#@FA(Y^(0cO4[1QA<a]:g:NZ&O4&
[b,bEYP:4Qf6Lf=Y-7.19J&8KBCFKKTPe<b=WPP)<G2&Ae+S1Y6VOM+9J:1H3F[)
MH97a890g6,^f_HeY\c=g0Z<9D,3gWg^(N/,.T>D[_):X)03V):c/R+S1UB&c.6N
cQ860]79U1WH2eHNFTB+g7]T==RR7b1J^X?,QMI20^/I1>_EG-(b[G?2^,GJJ\;g
:A/EV41U9bLMCU-e<Y1gT&N<FKILM)XaU^+)8RLO5e7++=PZd7KR@.EYAWYg/90T
S^?9-0;/7F@NY:d/e#GLK4-7TMZ3]ETM#X>.>V8VWb[[Te?TMW.ER4,6KJ0BB#83
dYO7V+O_T@OfC9SYa/-E2fJ@PW\V]Rg0=V/fT#31H](_[K&0BJ=FB+-RG)c8Y+Ng
:+1UQg9@X0=c)?T.2U)@BB0@ZE5eI)cBQ@7/[H0:#88_GfacPf-2e3B)gecPC?L]
)a9^c+USGA@K:H=ORA--XH(2S;W(>S5.@BC]ZgF?5f>#-]bOMV/G_SWd_3b,[gON
1aOeCD7@fBO[W_.g1[Z--5.O[6TOWGO?H4B<;LV@B=WJ5;.&gCT[B3Vcc:9a@HP^
P:Hf[8#:@6Q).V&T)Q9B:1<fdI=FC]d)O4?N90BS>USZBE0bIQ?<f1^HgSfe-@a5
cO<:AXT+<+66_S^EI2A<_-HYCMg6#bU/c2beM:I.e\@5JOdT4N)>RV.VRg1+CKb^
2H<)9:\1CT6Qc-2>R61UQE(4HS@LAU>40&U+=4-1Ud9J[WE4KX7G>cUMZY@9S4-G
F>Q5_DQZB2YGg_GDaS__K\IL?2:GfNDb/dL(A&JCW&4+#\K(=EPT<L:#/XA1>OEJ
G.YcTB_&PCR:;/3d8b=)42gY8^\_WAMH[WD]YO]^N7R>]C1WaOD-e([A6\.B^D4e
8YEI]NcO:@&0P[DK;-cR>eS?@Q>b)bASK@[/[-KI\gAYKcgU6W^QSaB,[FNH=-UI
&c)]I6R2UNPIK=HT<U6666-R7R[U?NH&dg4ga(QRT>dBY?12eccaNGDRB0LH?)?)
D&EOXLQJePf+QH>[.?<4AZ54HQM,6D8;c]#O3&R;:4A?PL&+eaDYa+;7U0P_1T<U
fU4-Z[RZYBD84?-XZ\XLA/J>YJWATCb<WQ4;&TH[S&BNbSL3[VG<,V[9)B3Q_aT0
44[:-D5Ad[dQ-P4[>^Y@SERb7#/0;7Q<6C9);9Wc[Q8X1(V\[KILH)AI1OX&A)W.
D13C[)OQ-GB]R+IAJHC:BY]J)2-/3aSB;CH0[0HR9,G;(?a1#B-=)#@TS619CV.#
CWAGf?V6A[4I26KaN4S#9-XN[>fBU9\5;56#/S(D5Me_NFa\H3SPd=?SBTbbE1KP
S;@9RbPCc.4fQTZST]J+A-0[H:E\7MR5a66>1Y]:E8;]9F&UQcCQKC_(G-)48BA/
/(&P)>-6b:0Y:KDY5D?3Y6/,7M;D]+G>_VW(DgMT_C,HKE_=,SIZ_S.2Lc#NGCS0
X@CSM5b3ST&R&MMcQ<PGRf[EKIG7AbeFYL309YG8aF_XHZ^G;^>/WRS,Vd>,APXN
+_ZUK&GC:VHYc<OJ:,WWK-;Q&[O&C1KB\8Yf[7K@-PL1d3D?:\SBEGRfNWFXLK_2
O>NY4&=-aE3/L5g[]B^[M\XB<PWaZfVZKd6?f:eM@HD#CXVO/KfERM]a11Af;<YP
QG,L5>HNY5A+L?bK#bYX7HWF=M,3TbYKJX,3@ZcU:EgU:f:EH_C0cK=IU8a/.>A\
(GT+,<US_V:ZKPeD-_3C=PR>HQT^#TN0<;C3fHQPf6aReGd2@YPZ7NG/ZH3],1^d
,@D=+F3NdQBUQ7SbK=2Z;\EVE^)(,fX?]66Y,Eb0cQV)BK,]9#S<C;O8<If7K9EI
L<JZZd516>\\2g)-\7;90QM>c@20B>E)OC6gV&3;)V1KTH15T]^)Ge80&0K(@LEK
VGH@QTdHO,@_P,a\CFHG^ZDW8;-<N.2D=^@NcHIU0F#g3:^aN(9\cF0\+7Ng0R.+
</A;Ge3HR(P0EP9:PC>GHZN@?>6A,f/W^19dE2ROXS>4_\Y2G5EZ:GERV+S.NDJ^
[Q4=.Te:=&R^@&4+JcNTDgO?:1+>_T\R+2=QfHb2K;J)FK>0Qe_N]QGG(HX>)ML>
=g\J:^0FB>dDQJTYF&P>15@UcU7b+@&:TGGd1OG^F&]HP@9/cD+8H6AT+K2,8g8:
9K.e(0U(T0-8?W.KfEdcNOBR_<8gZ&\B_2feIg_O/aJ&Pa74M:-5F:K_g8O,1#Z=
BK:Y1T[16:b3[OPd[b5B7N.,-K+6gdgPe:<6Vg+0TBAB&(g)2@5J?gKB/0f84XeT
HCF;.cP(++_1-MGR[VM(JCaRN0[.E><:[S0]]KJ)f&SfP>WFgG2]\#-E-]NWdcHC
GSZ\c8=RX#DMMS=SW?RYDf4XGFN@8X38W8\>JK4.:F4>OV[AcY]+Cf:9aB9FOfdZ
?EZMRZ3_RHC&7PH.f3[B4[c#\V9R8cQ95)U/3K3,I-f6f6e8/849Q])8LC:P3-Ef
XPOSFf,&cP(V8G;+PJ<.4JcRPH7fA^Q_V@=bLVKQ):X\3LfV_ASCB;??9BDVHXRR
-.eTd)75+TMZIgTf4?=4R6F,&cXY7W[,aX5DXCcf_Q7/Id(be;\SHIScR:?M&?#J
W6\P,C;ZQ<+\07>U\eDK=#-3T/2L@Y[;g>fE.]@R3b2QEG/0-f<7U]+5U\MY&YQ2
1ER?ZETMX/X5\)-O[N,^><7Zg@G&9M=WLM?.+:0LB5fPc>&:WEe;6,4>5XT^_>WH
b0\QZ,R0][>E[Q#B-#NM6X,RFg\03K7)SeMQV2?fEY-+M3AcgN=e.YJ>@LRXMI\F
[,MJbL)[-6RW7?d#CAbWD_dA0]]OWWS9XFEJKYBFfHIF[-J,@/Z\N0Q5A)^JW9gL
J]Ke)NBKf:FE5H)556ZKSSGTgT&4RM#WM8G_+5eSQEG5OVRgM_08gCO14[^U(UHd
:Q]a]>8.bIWHSZ69IO5Re,XHEEG<5XE6RaMFD-,DC[_>(76?G>@0EU(PVS+O?8f1
+O&^F,2)a-aVH76LRQ]4fE)#O^I[eMSV2@RSF.-RU9R=fHVP.N)PeGN0W&J[]+N,
U@AN7B+O-E(N-7GNHY2PQ@Q@fEe],d(X2:bT=d=f3gZ?=(FN;\:585QfU4DHD[,G
I_[&R&H+RU1ZEaPG(#+_7EYK+S3aGGHLZGEa)N;?f4)=?c7@M18/PS5UXdEYeW>:
eTJJ\bZ@PLH4=QP8a^^#VJ9N3LOaTbc6J#?&S>JJ8(S1GW,Q.aRU5]HUD5LVG[Y:
TN-f?O\,CK1U7\T=]G@PB](a0>3^)_XdW8f1;g43,=YJ?DKKIZ;ZBWc9NPUW_W@I
[7LYEY@5(3R_:.+];7&RY2B?0SL_USg)#E>2J<R&O=d=I#P6a[OP/L+JA_AI^_#@
XM(8.=VAcWXeXA)+>?QRgK3LCgH&U;T12PB&W2?][e.U_?IPcH7M-_MGFQ/AfU0@
(6B9?#)ea31BY?b=Q#)I875S)#f:d>[#UA#Z]3X>8<<,21XOe0FVLH8:.JCSe?G[
CB+\U&DP:RLHAK<+R#C[]>Kb-f]E@cK#(LIcTaNT#9e9)g?LaUM\M7aQ4W:AcR_C
2]Va&8-GT?&X>c@5b-4LNbA?&<LE^g8)C8,GeY4.5Re;/\g;Fa76A(U0)<5.(0=]
,V[3I-F>[C+8c.=+):7)2G\I?7<@5LA\&]#\]G>X1QV4</WEINUcG/GEW@H(]HM>
DA6G/FNZD8T0?>CTYR2>>K)XAPQad5-##-Ob=A+0KfL&#?@1/2FB,ZTLHR9b1\Pa
V5_/D[b&cU8L(MQU4IX?Q&=E^NeGR(;?eNR)+;a:f]1YS^>gMUP2OCZ;TO](K66\
+?;^b]d1>B57,]R.KPS/VXK5f\UCWKH,e]g(D&O58Ub=6&b-MfO@AE.OUd[J&KV^
:N#&bSPX-[\I]MgR,BS6fK+\&&\/D9^K_)Bd:6Od<WPd(+9X\L<@0+S<O:LKg6./
I+EQ,BT5^:>,M?eMT;S0:)PNR2GGUd4eX_K.8-[48b0,DJMU(5&?D.KCC1MRSOFf
gc83:U-#<K42_1NT9gKWeTH_U=/Y@?87JZHAU._?ffFbf;+@YD@/7fFOS6V;?7d,
\dQ6;7KB8de_L#T&aeWab)>SPR9\)L09&d9[f9#ZT>_Z3L<N-Ga3gO+L13XG14(0
U;)-<33]?_a,[@3GYD=QG?_DeE@:OaI)U<8569D?/g^)^K<5geZ1443[\[WXYRK:
<L^bHB8f[WHZ^UH?F(Ye>\,[)0dc2<6S?5d,V8O6OECb^c#,d87eN@KPH1&cL<I7
b7a&?OPASI&\RIU(O&NY<4>.)Q,)KLf+#J0D.Q.M,\TcSLL1^)d,9?=C^W+ZB@_I
T&:Y@5]fZ0RMS]WDN.c3VSB,LaRR7G==<Gd?WO/?.?BT;3-G#(2@J<_4BMJ1@_6^
UL+aSeQcJ5TGSK4Ga\+AA439[O&KRKL7gcCeABE@)[=[/RfcCDOJK<MHR6N<-#5I
I-Y[&=\/0@gIg#\J\<)D(),YbI3gMH)Re5N5N6E2fOReb(d2?OHM\D:?[6RLL-2f
WO+bJ4B9A>=,IBM>ET@^M&[?8-Ta.,[@gWf>@?-F,f[V^eM&]C&Ga):/8HD=NBXM
,;gY&7BS.Yc4GT-PAEdNI?Ve^(Tc&9MPCXNe42)AN;6Z-X64<RV1XC.(1S2=1&R<
]E5Oc:5]c3[N5?-9K0.ad2-Z+H:PPY(ZGUU3d?gW9a6+S@(bTMPG5.C4F>+XgXWD
eGDKC>&<#dO505G2QQ#_ZL^L1<><CC<_bf/N;LF7K0S00[M_>G/8<V8(C4_e1gCe
NJKaF6cVKV1XUUTd\=EF?,?XM_3JJ?BY-D_>Y;@a#\U1g8V:NO#?^#8Y/,KUMT=a
e.c^E96V0M,\^&<6ZQYf7f_77fG+<<<4NW?P<U]N+DaC\L]<)3.Hf+6\:GfC-+c=
^TdRd5UEV0(abRC(7-;g9^B8ZQ0/0JWZf;8^1VQDG=JQ5J7JE5J.;:1G/MT--)_=
RBV9.V-K9.<3_0Q5TM9,)cAbdZ=K49@/16_H+#NX44;=:QOYCNUeG9X0)Jg\a^&D
F58S/<TgWLC(VZ9fg.^V[MEE]X)O=b-HR6<DPS[,V_<M\O=J>;7Wc=0I0A0,KD_6
OY.FaILTOU?F[E3PL84==]B)7E_<DgD6-<SNa/.7Z7fgE>,-FF(#2I79XGH0)T,E
KX,D]A8?(>WGbOL-ZWB7X0.\+(;YgK:KW^H9)+GY#MS[95F+D,-YWTLJVe=TL?U(
?Cc4g(:5TP^dI:RO95.=C+U_/Md5))eg:(5B],^JYeRQGN_&b,88+8#ZLKRW&eGc
H(-5D^c+Af&FaORa2UOB82G/gL&+PMXNc+K?#DM8PCZa#=<.,/W7.6O]+dSEc_Qb
;5J>):c9=>9.B&K#F\[L)^c\,?2?d0ZTbP+;QV7,LFZD:bX86=8ca\RK7IAPQ60_
]^LF7.1LCcEIc+>P7A#[LS#&,caR-F10#TF(YGVP9QKE\;OOW4f?7d.JAAKTQgVV
F?>IA-(AY^7\AD9M)BZPN+HY.Te>?f8d.;Lf3ZI-8+J]J8ZN9:77NTTeAJ:K:Q;<
QJL#TE+/Gd-I3PcQdQ^(NGF7VJ4<DXgOEKAIIU:?F?Z3.34[.3K(.H<>L>^dE8,H
7ZdgK=[d]8:23._bMa?8GY#,IA56[S9KaY4Y9H@7GIF&]IT:_?D:C\>2GHIZF1I2
:D)GDD]\&^B[J@NH2@Q7QOY2&>0U;WLf3#dLB^)>6=MaI4F2LLU(AD=IYH-S6eXN
c==M,>IVWHXY(NRBD,VZ35K0E&W>IW;d;B]]Q@dZWARSU3@CG8YNJU&>:U^WE3Gb
db_C>2GcIdGMUaM<e)>a;SPb[_>VE8<\?)03Z2IO.)Y+[/V=]JQTQVCQ^T/:.(\J
QAD,);IF)^K<N.N]O9HFWCcL):>.XDg3-FLU7;#5+O)H[bXJfK(<Rb>[\I(8@fMU
>UEB(1K)LQ9[eX2gU[GFR,)Y6[F7IX1WO.#c4/Y.-AOS3WY+2O?L^5b&FIgX&QML
QKF7/#:a6BBRA]J>7\.Q\>?fCQQF.GJ9aF006H8/L+[K^T#;.(/Z==/=gQ5_E:D?
ASY;?;2^^]ZPQ.,DBK?Z3LS0;KD#=WA]BH74@G_G#:@;QadURFg#/K(GM_N)X@S-
OI]95E5_a<R6F^e3&#cTKAA)TZTO#]#84MWNV\S4JI8Y_GRgV,_LgGU6/LTC@BK1
V+\B@JI-=));GEA?b3^TB)]#,X#]e2(8R&d^YQ/S@;R5Q.B2XC86=S[YGG?1Y3ZP
bc\:LD7EOF>O_J6//AD9aML56:fEaPX6ccQ.Pg?e6X;GObN@7c=.:H#>#KNY<2:4
#@,4CH[U>PgP;]8g/cJ9(ZT6B&,MadS_IQU5+HQ.O?Z+/]g2?Y_K>fP/ScC5b(B&
F7&^YRU]GU[IE5R0YBSK1A](E(KOBYeM.:Y#4M<\=\b:;1aV)_P,)>(cedIY0KNX
P045Q;7AEcP)f9BN+&9H5caSc\HT@A2ZPL#J66VAXZebT\JBV;ffgC\[#IEabVf+
gLf\3\09YYZOZ^TB,W;d@?Xg9E\GV5GUUPV)fO3-QNKM-8H/XT5BHVRN4R(f^?(X
,Y@4.=Q-A;R.>J)a;UI,.:(A(IJU/3=PAd=_38LX,CcCg9];b^dLV2\]M.]Jc/A:
MPVI#Q@7\<7E_(1Xd&03L]E^U8SZ;B\,9N5,f60O>Z6P<);f49];#gX:B+A-KB,?
9gV-A1E[2.2NJG-3J<KRD8f8(U+@E(D0&VSXYWGE;7KK7eV.MgTB>O=LfgJ12dI[
=E0&8615)\/JS2OJ\ZB1+AZ;\GK)ZK/AM/V9\aW7S0b,</fN4dO#g8X3D:CYC<7b
==Ad#1F\J8O(bTIfI5OD2DT(cC[=:RC0^N._\:#BZGG>ALL.[@EMGO)>4EYbXJFO
4BU4-(V\CR,.][2#K<#0=)Lc;618:LK\L7;1XCU71LZ84JP.2&(eOY>>aJg;MYXG
Zg8YYB[S\c>WXf9T5&f5&C1DE19A9eNP67^I)AM\\?]Cf]NJ6];S^[;W=78+8V+E
]d:=U[C2,5<M/V9c@-fMe18S02bXe\=0W#.1NIP^f7BEJR41?+=Oc+dBP^>Sd6F_
\9+9D++OQ5C-_L#IB:(P:QW?,1b-d4KP)5g_.B6.bE<30;<3a3N1F]B(10Tc;],I
TV#B:QQ?#8U#0>WeSKGY8E3Kd7FR=USa.gQFKNP/88+UCQ)^6P6_@HL]Z#Sc9TK-
U5<0aF0NPa/SPfWX0C-9gM9JVPPE#(M</^e0D2:AW-CRHa^DY-Z[/bEGO9c96IE(
S/de08]9];b..40K3&:DIK24NPLa2>^\D-</1&6I>7..^?,AHLD8a^K)ZG55(?O.
,Ef,&YAS,XR15WR)X\dSZ3d^TU6;Q7(4/66:I?#[I-d]I?=U>=00]:@DV-6[L]cM
\F(M9f9V<JEK0e3X6+\Y_#NE:N.1]+bWO6<><]XG]E)82XgfO[)&UK&+CU9-N)N(
<0:=_6&-6)TW>WPK.5B@SIB[UK<CHZR/8>?Wbf/(aB0.0FHQ&^:F^IUB2P+Ac,b2
F0HG5960P9^W;L0R8-@]@T93(=0Y6^;<-P,#U5\\8a[T0;/ZKIQ.bA2NaOA2>^?P
#J,/c_SNf;NUBC[NV\IW6/C,^g8b):97Ja1DW+#PMZQ487:VLS_?KD5F-baNV<WK
G]Mbe3R+2YD9,<b-UEE>0=Rb5((A7?>AB9(ON9S\c-c>bOHf?1.d(JYe<S^)eOQb
e5<[E==5<Pde3?O[BKY2HY0-Obg\+e)90BDf[EVK.KB&&J=IZMLg->f(:GX#V);)
GKO5EG&>K5/cM/&Z[:42+E/OQWN(N+<f9c1R6;3B73-/:)1Mcb4XWaGE,a:Q)YP>
?AUK#JJ=5aeB=-X39c,a_F;@aEU[YD7Y2O-]K3XOAERVY2SNG6f=[M6DHO=Z=GRB
91bNY2JLOc(=9e-18AS\eAa[T=^PTF+,5DEO-7f.O\LT)Ab\MQgaaVT6^@RIJ<&6
f1EIIRU>/<1-9Dga-LK4P>SL4Fe:Wc@W/N,]aFD+J72GTSWd7=V>,5-N^ZCYQ^b,
]?T0<L+&72Lg)13f/9aSZ/TA2&/>dCZ<#9_eId2,+QRDYN<;(bBDD75KQfN4<](]
?OE9P<YG7;^,g6_IW#=6MCXHLVXdNQQIaQ)a/P2Z&4@3/[bU_0C8Z9eX_5P31_De
38ge/07aJe.1?AgD)DCMW>:+__\KW4.&eXg<.1A(P;Z\OQO.Q:X+gXA(>d\;NWSR
eY^1eD1eB@C3LEJ#JXO=eQGbZE;T)P@E>O8+6>Ada.fd?(FUW0^G7I48+g&D;BN?
P?eV,ZHVLc=b79c<9_46C9D^AR78@3f0,;T,Q_+#1IEUaS9#LIg)9ceDL_1Y-cV)
cDgAeWS6:JDE:E/)Z>T5@a8&9?Q/4db/aUcD>=_c7<4+HU1555e0Nd?7/,6M&6,\
?&@,1Q,_EY/c->V#F1:@\G(\Y\;F<R5HRX)M\M-<4BH+SUb07^S@@2QB>P^H[>3.
d0a_O\^PP_Q.2/bGY\;_#3cXRU+3e\JU,#c8]LAcQ3NN9/ddQZTQZ=e,5/b]T[\@
5>a8^PcASQL@c]fc^Zc7.40FFPa(A[IdH^N<PW8.Q\9dXa7VX.O0V0:8/X&]gP.E
M8JZRK0(240+:K9P;B9HbBDX1]UHVg]^YZ,.a>E8C,O-FMe>^NNX)&=:fZ,=;EX0
fQ-^QN_I1>VKOT@SHa^](gITJ2FFAMQ9RdV.=L#b#LNgUgSFWJ-DZg8[EB?8#X45
F/(@<51cE16EBYPK>&aH(YV3SE)IIT,?\KLTD9>&DT8RB5]-8f-Y+]>PUK6/9JCc
eCL34E0:O<GHCJ?<HAB#F5@T9b&X,>8,G1><8bECYH0#\=93NI)bdEXTeF]VV#=G
gb3U,UgL51UJTb-)L1@cDXQL(]g:0J6\KF(=T@d(-2TPf:J9Se0U]aB+&9Yc(U<T
)?7@SHe4AF_\TAI?^J#PR<\O^]UPgYMKX<fL7SYWDfA=>W/S/L5QR.;UYTH,3-=L
N=cTP[J/6XHg#dSW1-M.0PE:G)?M3b6?@>A=<YOa8W<^U)O@?YD,/1fO?1;26[cB
DBXL?8)MO6Od-0D1ebKH?;5Z/^fZgA7X-.AF6f5=3:WKI#11QZ8PY>9&:):+U/aW
N)G030fA[?bL=_Z-:?;11I3?]\F4VTX7B)(fcP?M3ef):B#\?S1DB@3=KBZ_Z1R3
A[\N4ZgMTI[ND6V^V_Z-a/]<PQbR8-NDY-Vb0<L7Hf[1Z/>Z)BPX&RR05^?Q6^-K
eS6_6IIf0J>69GHc=W[Q3&B4HW<_/M<31D9)K56K=SZdY?CP(+eZLGTJSc>KZ87@
U1(SA:9#NB4Z6J82U?+934D<]QbQQ0;JK]0+N&:\D4169#2=IT=/BSOD^aWDRF2#
K^=cgCDP&:TUGD_OOV+\C/?9,/ELJ01U/\L?TH;+?:<DZ<=;X)+BX2Sc1Sg<OgPR
9>JCd1@e4/O-\L+5&\.(HCD(YLgYCCg2PMAgN#8FY/g4U746VPPVBb+Z4OTU\9F=
e4#M]a,-:GE6<#aN/GgeI0HB(&3OO/.)LZM;9PJc]\6^g_6E<_>g?H,9()N51ZTM
K[bZKTa<Z;,Td@/OZ9#Ne1&KIYZRDP&Z7<C_#A@dO)RN5BP[fS.VHa\CQd2XU6aN
;IgD^66T<I?9.eC8GCe>=X\>XE4C(4Of2/4bd:@fdKg.ZTGM(F#6SK+10H)OG.Hc
L1RUR8WTE6L4ACSSI\^<0)P=FM,8V-gX[3Y>I&KLJAX^C&e9)IFNgX@+U,:</47^
M(8DWgg]ZNB^dVS/F5Xf,?cQV4,&X<3]KQ2&RfIFTOT;6C4^c0_X#>JNQcF?52AH
a5[_^#(<S4/#.8<N.GW+R@c=&U0:.DG165[?]gSW]+AAZ9]OOJJQ>@:POg\FSbBV
@ORe=A7<#HXG\AdPSg<PHfLZ7=5+1R.cS>280G-F1J@_U4ADUWROV\MEK=G8#KUB
?^\#L;9f&):R3O3O.^A;(b4?4=X<ZW;TQ&#9EEMe9OeGR)K-UZSJgUA][ERVM#=3
9:eIgfYE11WBTBf9FK^PAELF_O]1e?0Z_U>aIX]PZG@K8E\^T5M3@_PZ[@\.K3b_
8DAWW92/>II-LR7NK7ELZ/N<Ufg^C8\/_#<>+>O@gUb4]b[7SIV3\3^7>NKK0:CF
^N\?2D8R]0HGHEO#U8Q,6T6K(a.7TJ62J(+,SbK?).(9d8.]-]&JPX2@6eL^4D;M
BHMDfY6])2-)1GbcH7/?BHX:&SJWUD<@U)UD<SY^2f:Y6[SQ7RJd5Y@+.@&IHF5U
V;Mf);;4C5.]TK=9+EP_JGB/T/5W8:SaW=9/D8E0a\7[;6<R8+-J;]7Y:>U5Jce1
-)LW964)a44fe<IHM.SS?REf5<TJFKBT9Xf>STJL#?JVe[(Bf=dW:B]X6^YF?Q=L
)aCD?U6>SSA:J/4b\8WGcW-e(8._1<GHT9YY<6+,6b?([D/.C\;,.MgZ>#A.XgS9
U7NTL6CM2f^05:)W=S;5<0>J04Hg>c([0XBX-UFKY/eO;,U:01=WLM-SD]C0HeQU
/\DB+9F#M^P1A#=J<Ze_^a.NLPd@(J::]XH@AGdN)FYYdF_;RAF,a43?]JXef[-C
I-];(,/@>eAHCA@+^Lb[IEK=L.]T+RZ:G4dMM)CcW5HB;1:B]C^:Y]b?;8T_WPBP
8JeB,HY>VL+d+_,I1PAG0aKVeB?dYJdfM&S+V(<V#b.&-R:[6e<6P@fKUWb/[bCP
gSa&Gce:^&e,AUACXF4/b3>Q2<4DQ9B<g)GFYYK_SCQ5?,B#G4J;)2@+LZE,#B2a
dUacY0\C_H4gfP?_0+gHe?4FcD94+\P3^H3/,SS?.NQf9JYG9fCQO5&2dW=>ad;N
2HB3WW_dMcRTdANTSG40+9?F>R7=fDL[c:3@;QJSfS\a=3(ZZV_LU^Rcf\(K1SE1
48U:BB1H>QB[RM>1g2#N][_>fDcE.]CPM#:7JFV=]B_+Gc\A>3aPVY\KR,OLIHT@
[D;XcFVU8S:a<A&Wd@+DJ?\f2O>QX@JQRM8#SB]_9>1gb/X^;XN(c]QL6YR8@^eT
[aHDQS+=:?6FSEBRc?A;LdS#YGcLK7]be&1A>VU@/=ND4G+g7b9QUNGd<Ac/f][T
7P7GWBF,Sa0K2NgR#Za\R)@YWf;&[9?aY=9IBD+26Q-7ReJ]8_G9DNL3V&OS1.=E
H/^1WDZ1Q753[7FJL97H?7+>cJCAW?1-F1>[7168S(f7^_c&KR_HF/5AX@,ONCD-
HB-aV=2[2#SR0XI>)E.[GO]K\A8]Ggb8&3..Y/YdFf_/E@bRG/IOdLAdM#:.CN.J
b_fL?9Zb(&S2b?GC>LRSTC,OH5bMQ4&EUSc;MZNa9B<b116BX3gZDQVZ?(:Yb9^a
_H9c<5N_L:A8,NC)]XS(4B87J(_2UC2=^E^[1,FA+e+_F,dXU4G7,FDC;)MMA^30
>b/0U+bI\Eed]R7dEM?HW4N4g8<J];N)UCeWKg(8TO:SNQ0&:HELIDJ(3A-B2A\@
V_LNA71U06-MbOI,LaX0d[H-Ya5?1KZPOJRL2D9;1RR\M,B\d^>4aAU[K=NCNN+e
/L:B5,>+<Q;;Ge;D?-VCZ>72D;Z:ffLB;<HL#2PE<)&L/U1<2Z#PbC?)CZ//>X&]
EU?=JM)<e?He,ECMaa59.\d?)KdC+@7J^,HPG:0HaFI4B=5#RN<g.L.K@4X#NNJ+
KeP9>>.[1OZT7dL4T(MZ(aSNX>Ec=b+6N--ZW/Da@P8T01MA=J/A7#;[^I4#JQCX
XC1=E^8=)>6Md0SNNP\-Gb+(XEbHCKaBAM\UKb&\FV;DfAe,aJ^PG[)#b/5\RRcV
e//\0I@1c7.]\NbP;_@be2Q]LM^HSgJKeP;X:U&IUbWTZ\CKf)LON^91c5d;SRAD
L3G]&Q09S[8#7U<&?,V]-Hf?K\ZbH^]Jd3J?g;aZR3AKgB&V,T2(]NV]D&-DREG_
O?38<9gTMb\BOQ_9TQ/+gc_IF9C_B#[b8d?,INcK\X#f,[g3KM2^CfCV^7[&4=7+
^8P[^(I)a:cd]NbNMK+6><77=+b&8KA94-+Lb^?=AV&TN>?X&);_F+>6K>Df6E]_
#\W7:/b#_KJ4Q3S=UbS]0&UA&.I?Y?Ha:4cfT,Z51bC8_RQ?>=J^CV6<5MgUBL.N
Q)]&^D(3846J=d+HKc60(HQ(G]Y-0V)<)9-&]=ZWNJ>,;L1&-M<5JR>^Y6/WKJN<
5M?bBe<E<R>f-I<>.5gL1:0=:P\F/d1_-7/7<&4ecVFMT<TG;#[BN7I6NIG.UU6:
b6F>IaJb-;F/A@e.\YV6\B;TIX)WVNP:2N/JRf<a6_gVdQHV=IB#X6eXVK+(DN.=
9A5[TX5(S21S&?>K5VdFcYNe4dY@b4c1dcf7W((ZBJ9Y8X#W<Xd7-aRNCV&,-c(^
.=;EYcQ#eX2f7a[-I/-B<E-1Q\>7V(2?&JfW[We?8IP3;(8(,<O1U.?W^N:=.3Ng
U2e</7J=35?[Jf56\McX9E7JZ=HOQ@(?S83f/DfI6=aQ#4EGF]R,?VVV^gT]FSE.
>VGQ3(cO_]H4Y[E\YJM22SdVDb^ZX-3:0\_FO)>[1QFMe]\Z105CdM97e1<AMA=4
5E/:3B(L(4Bb.V<K-U.82NDY:aCdD0-I880#.;?7Y9_V)K2JF10cTC)Y,1SNZVZ?
;6=dZN6c5OV44?eVO-)(/@II6BgL+G(e3Nag[1UP3\Tg\SgI)a(E(F7@;S.]Q4E3
1;5\1\gcKRHDF5J#X2]]#f\R))AL(FSV/NBVGFH:MLGWc)Xe^DOBKK;P8#Y(+C:]
U(WZ>(f\;H<#7]gLY9f4eS#W/NNH8Bd9:aB#E\EcL0AQg.4Z<9)2<I1&-aG^[JT[
6;QF-I;.#8\>_:M9dQ_?<N:&3G^=(U#/g@NCMSLcB[+,AIJ8KEDaa#K0Y-VJB.1[
E];>J.X@ag)1B,K7N[VVVW@g355bbY(PZ=HZ.H7U>P[>>IP6#10&W9?He\[>>fHY
W50=G^I6^<<+:F;2>]T2)LO)V#?OU)I_6_Z/00VPAUJ/bBb<@<5d3ZM+9LG2,(2C
3C=WK)a:]e_50DB?8Bb4N#M&+ag;ZeV14V2HPQLd[64=R_A^:L^+-9IOL<4NeO@(
#O,ZOG<fQ^TPUV&Q_A76_DY0&c:aXO1#[H<DLQ_.RMFG,49c4>PYUfB+7Fg)2G:B
5bUF,Ue28ARR+b_(@g9L]KeI-E3K0W[83QN)3[5K\6cfBP37?FQJ/cTJ4Df)/68/
-R>IK:;AQ,;X0a6_&./4.TbL,;Z>X:A9d=9,9UVdT8O:9]?dU4:&HTOHa67H\g<^
46&OI1c,?0TI,bHW@gXOJN&M:_>Q>IK(Pa?aX267Q3)XWA2LHLg&gT8O[MR&<Q;9
Y)C2O;[ZU/g,eKKJc_#7,LTU-\e2,GAa&8D=PR&a>Jc3@:BSF(0+]O;U6M/)B=9d
13=>bTZIUONI:T-ga7fGEPE1fPV-EF/-eQ2^#I;5acO[JC/gZD-QJ5geP35\U&c\
25#[-g#AFC_=U6[?PI#]@_E]E3?WR,V\6eO8c7PVGFN74URGBEHG1ZKK2UDR8A^_
P#e7K9#H4aRd7aO]@7<J8^af4LaISDDVEC71U:CMNOR^fN->Af.:VYO<G1,\T)Y;
GLL@e)H=):];Y>^[_^TO8](gfVZ8\./,AWG[QGUF,(WG[33M0AM6YQC5LQR2Nd3W
BJEN6BV6PJE#N:c9BOa449>NIbAge-S5P[/CH1Ma(Ug,_.b33=f#/ZcK^3)7[#G?
Q3><-WN6LD<EdH_O;W8?dJEVC3GR6=QLZCA5beO;AcMAL>:4U<X(O4N)E+N)+,UI
Y.--QO)G[XaCg[U]+X9a#B]AN,R5gS\A6_W;b&gR2gQ\XCf9+)<R>BEPZ#^_FYA,
8D^Ed+W4<P>B9Q6):HdQ6=USeAJJ4C-K&IZ0URT=G7D:99,Eb<P2BQ1D1DY0\9_g
ATP?4#@?M><)SE-P,5a+Lf(WVD2^Xb7g\EgOOQ_CceDPKBVU<>+LW:TQ\1POVQS(
51c6(-(cWbb40A]T1WS,N9We&EN7Db8]2ST>4Z4>OdJ/)1._2&ILKfZDb6b#ZOTC
DBS7CULR8&4I/)9P7LQc6_.R^#/9Z<L8c,C<VONWISH@P@>+BZfKQK;30A(>B4T[
3Q=eBUJT+.d_MM&C9N8B7/E)aY+^?S8<3.gdVA3[],,5=KffMEK&e:9EVDAQ;8C<
D#_=RG#+;bge++E6d1J,2:RPMZg,GaN-+<B<aHX4ZM=>\:D3\IFaYfC]^]gAb\SY
(\dAXa,QMPMDSbMCEKAXJ8I=feM7W8/BPY]4&J6P^#STA#QOW7eEBE<XAX=P:+=B
)#Q@G0LUB=/TPN^O>9A4?9T-f?+9_=bY7RfP+>D:(c>DAfWW)-[O9G6Q[f@V0Ee/
9&5:N0\G#SM(Y-Zc3]O63#YHMUI3++X:6Y?&fObW=IT^O,PP?6b;IVeP?+ZGX,.4
Q&^QRaS]5G#M<Q+_]J6PPB&Zb7\bEA1O6T#QA8\:Lb@T>YO0DN5KWWUea2+7MgI6
?gPD<-+5aG@-NAAeY56^49?WH@Y.:VA.POEgL)g^6,^K.&9f=_>E2H1c]2+2RW=f
BAFUT>E+dMgI604DM?5VVd5HNE49EX>(/(RR\/+BdYRaZ0,ENT:=;+,4Y^CLU</F
HH,6H.QGR4cVU]-IKfU,d1##O3<eDTA5d[SV)6K=E6XD)E:>H5L(+\R7-=b<)=gV
)ZBf/>]L6NVCOSEN;J+__80e+FUBB9>RLXF7SYL/VM<HKF+L[<2,N=P[941C.b9&
G/&I4#5QeVM0DJY7eX#@4.<>VO^^&]>dd@:g8gA\4,:_NS1\P-[XG7-CTW5a.@VE
XY^3;<)I==38?:;Z/DDY])DgQ1(@?T+Q)<G)QHecb-.#P3EdbRC[:?U_R?G7N^Y5
[d_fg;GJ&2a2W6E3B-W:>6b/]#6T5=^G/L(YJUNdDce&,/NCAAFAMCW/-73DCLWI
;ET6[==+\Q<J#+S7O/gU&>f<Ad+6Y;#S9PVC6FXb-Z9c9=&+L0-Pc\^0LTAW3,de
\C[3Y]4CNOY+1.<^M05KX5G7P24M-cZ]3=&4<Z53dH0M=5aA]E84G1Oc>]Q:1C>Q
SYA/B;]<C8L66VHceP5&Fg:9IP];N5,0g)B?XZ&U@Fdb5:25/(]<,88FO&>]ZIZS
>?NVF_M6A-Z[d=eD4:14L>F@W)E(g1-X.LI;6):0GI@a5UU7?01He_8_.4cIf6L]
::@ZZF&9]WSM-\Jg_6][EYRd8YDJb4W.FCB=Z;9f)&^=&G16)2HI3#ZM3fR@[@[/
(HV,Y7MX8+X4QfL:7:FZS>I&G1\1N[X2RCPIB3)QMg16_;T?CIQB7J_f<BfdZ&Eb
C5((3H;=J2X,VU>O7X(4?1/Q)MIVZ=NX.4:1X5[?4:N&XE<.5/4TA1^0TU[0JVaa
G62FH;?-R<bA;(I8eX72APYUONXA03P:77)#XNOQO.:U_>dE0O2@5SDM2ZULXg;&
=DY2OWV.\Y6?\FZERO;4:YI)<SF;K^L^U?-Re(((dUI3CZ=XI5Kf,2I60ES,&JNM
A0ZRY>7aP?IJI=6dSU=6Kf8K[,./@HN&,\QVXGd0aAP02\LJ:2Fd)]978+<&Z(e1
Da/ceb:C_G4QM9N1c\-JdQJ9S1#O^1U[(QPU<Jd>VU^\@_J]AM0f>U3S_IIL)HR1
<1-[GF6\6954a5LaXA4,bEMd7c_D+;A#-H+(Md9f6DbE(&T2\5:^bGX=&V460BgS
VbBXQK5N&^3[;+S^47SWQXM.>&&>c3P(ScP_^Z\NUEcG:Q6D6HJBXd.F2EP+:<E5
S_<=WAeRPR1MCAXB2d]QV1J1dE(W;VOUeJb=f3:-1X4.bI:U(C/A.)DI>H^.VJ>\
=g?X(#g0Eb,GI,RD[4PY(7d3c(?c#R2)afQ7VZ,eFGgV2TDNc;GcP0RAC9?eKR/f
AgL)610=&J9aYOG5LbX//(dPaa+E2USf53_<W=SE[/<,+I_f/L7+AU;gBX[#-abD
6VJ<Z^MX.a2)S/O.;QG5>7,,0b1+IHHC(YXDILBP.L0Q;+Hb@Iac+L0cC_Q2g1Q^
=,H^E/T3#OGF]fD==C\I?N],(IC1UKdVT-+NgVPdB1[)3M(@Q]OK:QP:]@H&\YA=
TGY.2UB]49=gc>)J^C;H,9f,ER?1d:ZKeFW2^WIYd0<@>M)4PN+^cY&6#RT2FZdf
T65dU<-H#86QT[U-]_FW4Xc@R+6BZC^JD8YI7)O/YPS0+6,8JR6DIQ8cQ(JCZ;+)
[&?V/BS0GYGIeX>AN8YNaF.L74DDCb\<QA.CBF;SfP][<K?96e7FN[M3Y+B0C(e^
X#\4e,1VHA(b(5Ec=Z?T-KH9E9KDA<H7a]QL;1]9<<SS2YCE>T&&7>fW\DF^2<(;
NIBJg@:IOJJ2,I;D8Q_E^SJLXWCMfUbWRXSRb.S,d)dT(F//C[LEX&<L7Pd>6;0/
5eCUB.3dPATM(fUK=L4/IU1-EVKcg7ZM5Qe39DZYPSQ::dR1O\28D=1_RM+=LCGX
LIbH.b@E@65O=Sg,<,[c:6<9)XVF6=ZG;C(D_UT3g6/+IL#(dOJ-SM55/&=X@@T]
&NfW96cfN>(E#e:X+dK[cOS-J5O6?1,[&.dZ+f:&NNQ(eZ&6#4_BUfTK(7dFYDX8
Z6HR629[AUV,^dJFW?HSB-_Mf-,M0JJE\@&P/[1?)DPI[dd[b:?D,J;KYgLcO]W)
BfFb10)^=)\3a&e,7Y\QH5HT2:HJ=Y\#c>((5f#QFK<[d4?-R@=W_cWe_;ZJ=-&9
4VQd]O2-38F2F(W&M2WF:([fRSQQ4P_:@PGaL=A3Dg,(NOU(C<6318eP_S/8b(4d
VJ@7dGd+XIMNRBK6,P_)U>CU@A+N5KXXNZB;)/dZBgI20Hb_<U1;fS-]^-@JE#XU
)<WHd2NcIJ4&Xb/D0ObTVOEaTB\c]b,02^7@YYd:;_TE4I;JKW)6/4+D#&&=-UcJ
K9PcP5+OL&602#/L:O-Y@38DV()6adXEJE=EOV\K^-39N7:)S&NQJV\eA,Ia=72(
(0S@ZLSK_>#IMbMTa?fMR+@UXa4[BZ#?W5Zf[J^U0.-JHEMVN27SS-XZ5LG41bMV
(I(7X[Q4RSU00f3)gGaGLDe6>=3HK_]M4gVAJBP)g?-A=??0UF5J]KPJaG)RJ5E,
=Sb(MK^P2bfFC?]MU1-Kf10^<^JTQ+ZdHa581GfK4H2HPKg[FAB4/(>4D1U[T-[g
LTR>-+X8[J:ZMS@MH3caLV3aWPET&.16L&/)?N2eWUaH55fS^C6W]=])/7TAQ,Y@
,67E;aBF)^X),,AUZO@^\&#_Y+2/5\g:fALdV,-I(P?#BXH0UB?aQ-X1+LI9,_D0
9?(3D-Wa,e)>EY0KIa+6Bb9ag(Ye4^1H\#VDC2_]XU>V\BVb_BWJL2\[Of26)a1[
R]C[)eR)AVX_Oa,F\g6C/?5,N+JQ^+E1-#5#6OCE8\#f]@)D&7<cIg-:5U&/UCF-
QaIgGEa7;b4B=B.T5C,3QdGaWXYbZL@O<Y-X#1<c)[IJY?.:[8F3A=T)US\3Z#^6
8V0)K0@2&e(.@UUeJVZZQUR1]?@d=A&P\/:fX]QVSe?HaP?E5[H:LOJcfA)gCI1f
F].Qcb_e1N?O1+T^^(M-AM#>EHL[&3,Y4ZFCACMC,S&bE1a^\/[QbMV?a<RA1;a:
0OIUc[4^B9?W-d5.K073HdJTHGX&KRIb2FOLI\16Z1(H[+DOdPG7X3)>^c&)B5T+
PNX0O-6:&]I_[K,P)+P2UA1]g;ZQRDI[ebTW;<-I,9JORX29H5)YTf,-HH6OeC.#
bEB7.P.)&:dNVV5D4>Hc8.M<_?+\8:=KH/VW63Yd7E9MS^+=))dY^F-@\EFYg\03
X\d2d_YTK/d(S/RDOZfNgUNMRLANgVC12^01P^Ze\63\ZS=+8J+,L?7BZ4G)LH1M
6DSW37>?8YG\d/UQ.CNFa?D\4J>H(9Ad?>#M><W.-9EF/<G2JIKM9DP3:f#17@C3
//?QCd(9&X<0@^5T#a@g:3B0O5/bJa-RVQXV0-9BY:MaUI+.@2[6:VMIS2ZAR?17
0S?V)dMFMfgUeSCb4ZXaFJQQ<3dBd,YAWBH;826(7..KYVLe+,8WJ:QG)GN,b:Z?
@E,(GIBfJAI[+DaKBXR>ZONZ5A90?dfREf->H0,e]_+b7gUH]f,Qbb+2CD)\;PJD
d#6&M=E<MOaLDE/.DTTQ70O@)-L1f;RG1bV]13aWT8XGL1b7-YUE<&^N<0/92bIg
d4ATQX;M]cf=?R(c3RKRf-DGJfH0HR3fYM&?0e^H=H&.A@:dPCdJ:.f:RI-G44U9
1;NcCO/#b:.[0IW\#;(]D781^&O=aXKO^,SVcW4_.2#RdK+]IPaNZU,0(K?@g21;
@Sg#J+8f+XJ^Z>47I3&O6S-A8<^795a0J4P,0c]&IdH2\-D#VZ:S+<-0OdCV<<?_
dTd7CBfRKO9D79J4N?)LYeEYP:)Q6C#,3NXd-Q4,JDcD],;,).I6ENK7HW]DSXU2
0&1J;DdDH42#)7\5VgZ3=_ReIc;Q)1>=C[-g^cG2R3^NaTWf,][E^,;5,g8[.U?8
F[3,7+0&41<UU9b>Cc,]FgRZO>cX3)B8@[IG>f0\:[cG/c=<VDNKY1X#?JS@.Q6U
?YH\VDJ,7(/RFUODT8@IG][\C=T,QR-;HG]&,:9>7L.V+_1gO)I)CC1?/aQgW;FZ
2RZ\J6//2Z@UT\T\J(605f+-\cg3A>eF7D9f-PF/=U;V9L\aE?@<3DPQD.(c2V@+
Y_+,06_7-;[g&1(&Dd<YB4dNcXQB[]1f(EXCRZW;=;^D?&-c._5J\48^:_)eFL5G
FcTbX;5d+bD@H^Z?KYOBJZY&A8SBXAN\&@1fN=g88<I\9A)Za1:4)R3PMNNbJZG3
bG59[;H/7[TY^>I;\02-Z<:#GYQ:\L57_Y&#:dKGO0P;WL>#ef9ge._Q5KT\<\bG
,+^#^=OWL8&+0J_A[V;[a@W8O872N#YG871R@#gS[>54X2,gEEG1aI[+Ee7:7g9:
D]5IXF(gHE[#&][O@2@CZP/AabR5\aNHOG-Ve[DcB]XAOPe)2>g9M9#3L)U:#6[N
7f;6K.ZO@@=F.DU?\<RY_KD?0g[4N/M@:bPZ;(>JZ2;;-b/AU>#.d-_L&UU[X.gR
I:5)S4[cgeA?H42/;K.0)EI;V-SR.H/@XLNE:?=D/c)Ef,gb/A=.A6Y&ALH8-N\N
d_3W=b;4ZR^e]EQ_a9Ng3L9GV2cB:NfCa58DEUI.5eNBG@/_#PRD1#fFdMM-.;+I
WgF.+e4[H6&?&ED_X&V#)6[NXe1RLHGBM#KH1ZOW3>H-7^X=[[5RR/YPLM]-5IX\
WHRE6FW>(7R>?VXJ4_d+bU#Pe&P\ZQJ>@b.@^/)A1;H.^5bY6NbRB#9A7X[S6JQO
F)SU</O[6cW3+W+D\.7KHd@T0dFdO4GC>5/5TSU;gE#+)RZ@bW-+_RV.)-NON10=
#WIU7Y^4DdS8O\^FaHQHW&_EYOKE8NE=c&8bDO=4^20b#7)a,FaLa399_A90.B?f
Vb/fOYgc)1ME74X;,-9]AQ6BPA+#8_4T-RU.\#NC(ZH/7=8I1?IJ_.,GB-gc/B2O
/\_:OG+DUHg.L;,b9=AIbTV)-;EZWb(=WI36AA\UDVOaIT&W84O49V8??&-N>\Y.
ZLNSSS0D#TSDX-^N]U5IL-XHR==#UPCH[3MNNZBD>Z4.#G)&;7e+L+XaB]Ie)C=B
gg(Pd=DJ_6J,(4:Y\6257_J,>7@+Wg7RTOVMUA885S[c,Bb2[cLX>6UY9XVVMG3+
AFfOW7F8.,(@=3d:c5f5&I25[RgD5_#H44GRgL&TNR-=9@fR=U[fF4590F@#B#,<
A)KC5\32ZScJ9,Nb3O3/2_ARB=OVBF/9E(Y/QC?12MI]5#3-)^RYH#6RFY?Q2&fR
VZa9.4=g(&VZ@YVHH8VJ<QAYag=]=,O.8#bKE22\G13A:O=E9,R=K5<+C6&/+)gI
cc>c&Q3>T.-,Oc]N6DL.&3<TNf72d/E&d0Yd;6K0bEC>bPdBQ7<_fUY>,[8f<MFQ
7L;==5.0/WB-dV0(AH=Z.3JPfB,a/,(V#T\N5X?_0Sb2O#3dC@K43G-bMEA=LU^d
H>5RI1GT&f-cYcI8Ie/fJMI47C#V7M-d6YVCWQ>2eL3B4GC\L)/_S,-1G+PSX,+=
0FA]137U3(bRH5^&4E7-VCBPK,X6(c;RWR1<MW;\fdbH66Cb4.CNRFPgdP?-7[We
fH00UW:PQZ6G17PF,f0Q(9Z7I?FT&P(4YdQ>X=d3eY^&BP\#IG^G6VGP&5ca/^KN
:9\@UK#DE>\dKdK&<-_<Z:0OdgMS2(Z9-FcQJ3-bfaP0;1:GT-)KadUgQN1e33/0
\WC,46\.9=XBMOcRV)G?+HbWSaVX?WK>T<SJKeUZU<I+6<HL(IV(&_g[6U#.I]b9
?8fXMF0ebGQV,Ne5HH#@),\LXDYC6Ja+e4NY8UZ+e+7V(NURHXUG:d156C#:MCJK
1eFJf1R4ZRS+Z.9d+QPO;+=H(NR8ED=>B2M#W=GE?9)W=Yab1<L-C@JP9fdOMIG(
B3[5(&,,-1+#Z?466FLF2UQV=/7DI&RU=7=fd>ABE]KDIH-aQUUGK].L<R))AF]T
UKe@M4gR@0DfDWK8W9De0W7CM9BR:;#]T2\RYEN=,&,[7&CVDN=<Z,>0-F>MITe7
_L0NV8[5cU54^9.C_TN))bR[05]a^9.]54F89=PU/L8BS2-)f-_/I3deGF7MfQ;>
<W9@]WXS73IXdHBF;,?W1ge5>]\JM0:GXFcP\V03BMAeEKeQgVA/QNJ?&3FNN[6I
cI&>I<27F+1M<Z.dH^:&7(/:7_cX<I;DI2:a&Y).CR/AJf@;=-;Za?YWTNZF;DHF
5PRbf+=HB9T<&B?^.F:[0Uf5deD#a.DM&+MEcd8cB@a^5-,,W6+F]77[/f3>.gSG
2ZWO74Y>)CR<a:SZJ]?O7IA=a==a/#I(92])1)EH-D<4Db5GP>#3He@2aaI)Mb6]
D#H;F6X3g[77=;-@+CZO]&ALOD[H6=K7[OOF,BJ8Ug^2O(GJ:TO::7(F^QdUM,?@
M3\RD^UCF2RZ,U^95dg5+_(@.?]@B>IUcD\dY;XO_3c5cMSM&aTM^1IK634SWDQB
Q;gEdM3ZM:L=VXGQM^HDM)6NA[+NGdJg+e5D-c[TW(L+McXbMaP0.H^U^RRTaWRg
e0TdB8F1^TFRZ\af[#V?5.c0WM(Wb^&HFHf;-2a;GeKH:[fd=L]2Xe+/Z8+8@_O=
^#H03REa7Tb-KRA/=AW>e\BP@L)(IU>V#3QAP.?ZK=_bX;5C(L0::956X3I8G)eS
?LfeI?S;g1F@4.(FDfA<>>^g.6CLWMf\Uf]#?Qa=gJaE9<QMT))7.;R;/AZ:S=CM
>RKQ?I,-C(Wc3Se;/aWZ6RIW9+?HRS/+HN5C#g-WS0V7J+(P[QZ?df#F<dWQ(aZ/
J@XF&U;b;]I+ab8DD6&=Z0daHbDd32B,8CR#Y#,^9MB;^ZE[57?dV2LPIaU:TY&e
S(<M5(SC2?E\R8:9,NN1\YZ2,HLI5KfY(fBA8b[(EV@6[_=1O3AG\2OM&R..7?H9
I4AGYQGD><OZ.=PAEHDIPfDc]a<3K>0Q92V8V@[GBg9AR[B.0B.D9Z1GZO(1S6XI
6T0Ca&:)6V#e9aO89(JA4][4@-Cg+TXbaReK7bH]ZbFVDRYKC)@e-5T(8A?.dO1P
)(FM4[@Y3(7d8?0(:9M)RR]E1E4[XK:0H19DWg461HY.,R#NV9ASXa#=0>:GTN[H
:gJI9@U:bE=]]+IE\JC>5d&MEO71X[L\#KQNBANNN5+J-O(]fIRb1H8SJ<Y(YaaH
K.,5KZNB/5]@5L00A5P7DY;Z\@f9NS3.3Q<)44JOI=7LFe+bg)?,;-+&^.GWNYXQ
C)FI(TPMCA/9DXIEJ<7VO::2aDP0A2N5ZdVc(?&KfG]H#aa\@(?DYK+J94=+T\1/
E>V_R@T-:W96-G@BR/33P#U5GC?UHeg-YQ#S4JC(bU71.d2K7+O;dEOXYZ98B5@N
JAHM.4,VH1(79X,&\bJ.X:WZ9)\8.LI38]B]#8bVKHQ1B[[Y@SQf_?#;PG7b>UZa
F5B]=5=3<&:8<PS;A#D(48S2B=??TdYS,?VF]A1S=LXEVI&DCOK&^AZ;3;9[_d_\
\IIRX_]+OXNRO8Y631WU8<LJ2Ue#[20YbTbcY@<R+NOBgMA6X9]JcBF4PQP-cMBM
4e1eJVBKfd]Z(V;/KBV<,5Q5N#50M^a.+dYVU@^T/@=FQg[.QNXS,G68.Q<AQFN^
f&;\PVQR&W#NJE=<gO8ISfZ&68eZY8P,W8]aK-/3A>O(1@[CXCSbOQ8NBDFHVVYS
A:;+SS5aUZNWbC^F>=O^2XT4J7PeFg&0YZ&RJ>V/R(OTB\9K;2?(K/XMF>:2^b[A
,\+:LK3CdB6eG[@B2W7a,NXbKR(F<RN_T4J^+T;63]NJ8Sc6QFE7HT_-/2:()ZC3
DB_WB1?(57LJd^9Z4?KG-6=G\-9YU_OYELC0,\?1.3+;V^d8N5g6Kdb?WAV2XM53
E&Q=F?#d^-6.\I?/7dX76V5b(48G3^;V/C,g)@(\[ESMfF,P??,_/X>CS:eb[aFD
V4-.Ka(:Kd+S7eM,1W@B8>D\)BK<gX4:8\EBBaf)^#-P572O=g^]fZ)e0DEVPaPL
UHf>GZSg>4c=+6VU8=2c=/8cSbXg<L[T;]KN(/^O?ZWYd5BPGHaMK._/K49V]T.A
U&LbE/-S?d)f/VUf816\agI2L;fWc:Bf.aCD>281^9-\.IFN_)P;A;>1.Lga6fGN
RLX\U/L4;bF3AO:R9#)HX&K0ZM/DMf=(Q3KWX8=OU<f\bAFW=&9@UM)^#)BeT;IE
cZN/Z_9_>8(5[R\(_&WOgU[2YgO,,,A<5ZOU,e0fXLCMCecf,cM(_DeVeIV\<Cb&
2cZA:(ZH],7Q#72++:TR\I/AK^/@fO6:_e&/e;(C@O9a<dL/cL]L<?/W<J=\YbS,
ND40?@<S3dU>1-.E)L#TgbEI\4X/WWP50R@4Y3C<cC)K]0_XeUNB=7+GSb:.9(cX
[^Q_2;aQ<3^#)]?7Xe:Mc_aBYcS//:[AW,2ZDg,b5G[K>]1F/DFL=D:A74+Z&-_b
LA(gAQ+G8DAVNJ.@ceX)T>;I:23gd4^3/+/eJM)]?K3LIP/FVaV+?K^EGeg-P_A/
89BBZfg+5HN]NM8LRUf?O+2N4915U,-V-?M9/WeF^P,H7TfOa6/.T5.+P\P\_?<V
V^)J;ZRY/-]+eAb_L/J0aFZM12&UQfE[\@Vc>?L,e)V5X3YW.g)^,?&cXHJ]cUOI
?B8Kb0:GR-;ZE;+T92C6;d_IVb/IZ:-O2WA@MMJE6O12H.IP36gCcSVD[aXZ90\]
[6Z5H6gPN.QEX<8:cH)COI)O-;N5&#Y(Wd;bR=f&3&QD&X6bH_]<aISfOI@LWAIK
#5O5#0QYMC.;4Kcga4\\AAXDP;;-O7FH_YZ7&#&HY+V9QI\HXdd3T7(FJC75?5O8
XRIM=&?-Z:GC9@)8e+XFW.a@We\ONUHM]F>?9\BW=64ZV(XX5HB[8T\e(6\4X[\S
L-J0EN;M4[3#B6NS(a?f9?)H,0MT9W?VeIH3QZJ58HU+_SY+fQU[X.5YP,fR0H&I
/-,9F_COA]a>Og,L.:<^6RK,UP=AHTfSMd^95O-,bfeY]#KJ<W(Q^3K?&f75,ZcN
Z#J14O<bG7]RU18IX0,F.Ae?aU@JM@<ZK_PNTPRS?>7c>-5O=I9A_eZJeZJL65A)
7f;]99fbTH2X[;<B79A(DDU7SK48EM&\)+AIWXdGeO_ZCF4)5[)/2^38\J^IF#38
PZ_#H:LcO/fPD.c5;UDQP.?-9W#beAVW:&Ee3#-&I]I1bRObe45[\LDBf/O4J9RX
EVWHO:X_N81BIBAe-5;A\[99e/ce0DVRCOcN<#BRWF:0@:,bVHZNRcPFI96aHMTZ
\+45U8<5bZ9V]06Q.3UVUA5.5dc0/c46RDc@SSNg[[./3F.1&0@=>NeF[)GZ6)D?
/c7&EA9Bf<>_B-6X84\MIWCAL#DD#X^D3K:Wf>])A5?NbJ]:SGYP2C[T=._Z+_6I
dZ58-;DU@#&UT0+6\aI_S?aQT;9>ec_e>.__37@=CIR3A0^ANMWXa(;5P@>bW#:]
7)[PIRDW+9,Y]U8)(/U,@L(AB.d@.CX;7KM9=,ZJ1D7=5?5(ERCXQ90c-9f&2QN3
&,E<NZ]4=^+@f/JEHRX(?dY35S.0@;4=X<:W@X_KPAC]bSKX,D.UIcDVB-N&[<;E
FeG<D_7E^UZ&F2GW>J)CV:DR\XO@4)Z0M-0D?G(^c:Ca;NAZYc0EXd(L.E.YA#+[
FU3ETE:.6g]7aL&fE+JNA=\Cb1f#JGE01g2W[@=dB)HXY/?TQ2dOIH1[OPX1V-O&
d.5E=Q0K&a;+0MP[6(V)1UY9A@[(I#3RWQG;/W=O4Y]4-N5f?(2a6;9/WN<>.],2
D+GC(:1/[TE8:VJ?HPP_CQ][N#:&^#+O2:+Z>6K^PNK-:cI/Rf56JUHH):TO^(II
WL:VR\+0d?R#:V>#\NO011ZgCVG2fSX&\>d+1N]&bbHDO4E8VOVe>\@\/[bBaM:2
XNGP,-GO7f\BK_)MGKfX;Od6YKDGE-FbA3Of2a2\,BW(.&XD_COX#\ZO3eR<SY+=
_/R:c&SfbEeV#OJTC&fB91bO3</R+,6E.e/J.W_9?bfcU=U76?#TA>.?]=@IF7+]
;.+J71YU6?0PgEO@Wb:])L(FTB5/fg=eGB\F-@MVRX#<T@=8D#SUYfCb)50[-XX4
CM3-X=7G1DA[OX0b-QU1MX72XED5S>0+b>1KH?UNVH&YZX-8WXZ8I:I;E=,6E6b(
Pd/^=&X;a-(Jf8=#JVK)5/;GfA.CFTZX.f6GGX6GeCIL=L87WSbP4a(2K&gTNY=Z
5;[f9IF7OJ,&d<>.2Rf6.N<d.GLPN4MI\-,S9?7+/d2V;M+;/J)?-;e#>B)1;1/K
9JK(/RSJ5KfFb_S5f<>ZCVCZ_0eDM3XUdOV\UHdMa<@:Hf&++S;/1S)TG)G7b4Ua
F&H,1e1c0aI:OY,X3BJ3K<6gH#fC+5C(\+U_Q?Of@,>0[c5Cb?@5+81C?Z06.8(g
1^P7XfS2bY?,LEV8TGWBYbX.)O(]M0N5D,5[.@>dO161R]&466De,]0-Cf70O?fW
aZ6G7W6L+87=7X>g#e3Zfa>QX?_\&+8b8OZ:+9&D;R1bB;AP4]I@F-1S+DLVbU<1
DT>^F[,BG6D7f3WF_N2:G(2=VI(9Y3^R=8#D<?MF,FSD_L9e41SF7R&>&)9<P0H:
09418TaJfD=aYUNZ;R?A7BGDL].cTYA#e_O=Y:,eVG,.6d@UQ.NKgd+O5f+WgF\f
a8IXVA[,4CKFc[L>DK9\>ZX-\B+;d6ZLgLB=C([\]NZ3,Jae1DVJJAdaL;Z68aQS
+JUWa4D5\K[+EM?HF1[C_3dgC2fTDAD>g<+_NFA#8VNRLQ8.90BZccSC)b.]V@=d
+Z2-.aWT^@21_V5@]@V5Fg?]#MH5O<OQ5?T8B+<_OD66D\Ng?Yed-:B#DDY:Y9<8
<Ae=(A9)BgDeYS(XSF;?E8^1D<<=@=^2OZ1PZeY]Y2(Z5VNM]G.Y41gg+TR=PF4T
#NO^eZGSETZ43JP24MUBU]<BOW/&:d.K[Gf^V0g_F5D/?8Qe+#F(UaeT[PJ_Z8>@
/+FcfOHP<cP+@0[LP;&)FYVa.R4\KN#,NHEK?bIIXP@P-/@Z##R[V4DP\XK=FZUX
dLB]4<GX.U9DJXN:P(6X#5bD3Je+-55Y7^T+/+LDP(JP53JEa3\a80UHVL,.H2/a
RJHMNaRPM.&e.Ya:D.)L+&5&&JLG3+gN_=>IMcKK,[+d(@36HV(8?&bfNK\2,2Kc
4Z,F1QD6/SI7NR.).Zf]Zf&D3C0Y2f4\L=0aG,Z8f&X#;M]/X/RF_=5H9@-+6=E@
YAPAN+YDXd4YA;29+K2[e1Hd-(,T47ZO.,W[-Sc77FWXHD-P^H#]G&bEJDf0SUNG
Y26I_..N:Fd7^f?3[L5@EB0(D7,]d>V?:?:JKcc.V/8&Y#VWCL=OXY3b?7Cf3.<c
?&[<@<Q/Z]S0(XV.V4Na.XS/OOWd&0([a0L3Z54]d[QQ<)e:_0]JCX6Yb8]Yf)]S
:F;<P904-W-A(#F25BJIZ8AG.89FEQ^]KY1@3JU11<Gd;<)V0R?:D@;?L&V7>Z&I
]LCT#Y-R;9C,BfTHRe(9EZCG6EXFT[)>2Df(&J)]?.+K,L]e(^PYUg;5PgKOKB-b
/P=_4_f25f@R5<74NCVdAaQQQEQQN7^@bAS])FL_:@F1]+d48?K-Ug,deJI8-&8M
c@1NT[7VcP[a=W?<P5=A4QXMg7]P3)e;FeO;ND#XgKeSQS4?V,EF_T\E.^bNF^VP
aYe<=+2>X#>C6#7@bCV,T75N2=18eaZUcC@7&X5e:O=B,N\4+K(AIQVF\E@\E:J_
)U;D.DbU&Q396fPRN4VOGT/d3)#)CV6Uc?/EK1P_6-GQ1S(DJA?)LI2UP@#+a6d:
3.7bbNMJCRJYL:67^1W/578IPH2I+>^;JIDda;8,FTWI3e_F-,L\MdZU3>F2_2JP
K(eSC]cVEeNDPRP8W#+]eI:WG#(7#]1,#>Y#UPJHT\/8:I6LffTG>2KUC9GM=Y+c
DZP,M:F#e3)UW>]^e(^4dW4HgC,+8HcDgKe+:AZ_WBU\cAU<b0(B2<[[GRaIW>e#
PSHP+A^\U,ZE((MM?^V?d=H6[O/:\YTG<S=aY;I+3.:+:#II1^eQ<WJeeVHQS#=7
)-PG]5e4I7.S.\Q[=gaXER>GTC<f[N1[E0Y?,U16L94e>75UFdbV#G<Kf#G=N>-#
Sc.)Xa<+WC@3Q^R+UE28A1AI3M_-8/7:QT?Ye]GN0#/Tf(XEYY2e005R]@=FfOG,
?5,Y4g=cQ2f4=Y5ZLbH]Q(3ZW[_FIE9feDDM?9U.(2-S?MW[];28c#;:Df0Qcba?
:7)9g4=@a6QG9=bE,VCV??WX>XL/1<+Nb9@XC=(D=Z+LZJ<YXM]>:R.KOB4g(71/
R[6X8-=P+=>)e1Q(,W,7XMc2YFL3S;/-M3C2PY#CNV3^-e6LRT<6[3H\M]:@ZYUU
D0\\457e/:KdPTS>aE.A=B]1#<7]\T8+<K5aYMF1]KWgYH_G)9J&\@A;@8eJZdY>
HB0cRW]R_U2M(1\_<7D2.R9Z(NCBfEU&VQ3+JUW,AP#c>/JGC_8Q/GW=IO2Q6>TH
e2#7?1VfA\?Qa,DcL.D(/Faf/4:4@M.<X8(Hf.Ug7.FRQII?b809\bIaJfR8)43b
]&bQ<d@9EGI+J:]QH;I&Q?,CeS3be3G)9\K7\HgPC+=VUcMdF4JBd)[K^-;.58Of
:EA.R&L=@HCcEOBN-:W,-\P74NaV-/8I29FOE6-TDXCM_<MZ,a=0K0W>3M\,^fEE
\BU2XA2\?O&S/:7:Ja<aX]@#</7=U^f6.:/DK/96=T))HfMGTH5Pa2fI;/T>g,US
^R9bV8948#YV>7ZG+4J_6J)FGYIOP\^<V@C(0#MI[35S&Q.TV8B0dM9WXgfK4BS<
#)_eJ^#UW<He@]&4W;3@Ne4@C+g6.(d4<1D^Cc#0G5@\U]G)/1R28]M^8=231fdE
M6Q^cdA42,@./(>H>#B3/H1==LBd]d]<,O-J12(ARf3YaW)RJ:8=ZZ?HN^0.\73I
=>1SD)5ZA203d6IL-W<&L/Od#=_7b6Q;&F+bA7G-Td#dE495.R=S1ES3(WQ]26#Q
RPLV6VCVO@g=Qd=a+f,Q-&L#:bfDdOT60G40_a;I,3c-W]]XAcJDIR=MJ+_WRBJD
\P;U=Ffd_-Q@C^-_CQ8\>T1_RN7O^(G;Lb,f>JKDcBOf?IK92@A_@D\&EQGVTN,0
FBfQG-^aQQLCO>f##BGM5<+C-INT\CRMIB1,CgbHMg+@]^V,LY/+X+>#LWLK4V<+
I>3Lg3EVF.EdG#U3QR+f?fEF+ZeZ2L95A/K9GE)/N@)-ZIF[&8eBN5g=(ZJdO-gd
,DH(ZWI=7agd+9R+0N_\,0g_e^AgYW6>N00Cc6C7S<:@fI@U+DI9g3?1ZcR#LK^#
f[P#,HH,@+#8D-(Zg1[H>ON:P(;dX:STV@+9S2YL0AAfL:4=/[)0Ug?+FP:=\ZRC
4YHJ>NCL>-D;KB4MW:D8C<e5\)D<6=C>#AVCcf-cLL4RR.4.5_&NS2b&X/88-CLE
,D\Q1\T3e>ROGRKN3)_L-OB/D-4c<9BV4Ee:8?FKJAZ[_AbPQ3GTYLXIfGH/064=
30b[3N-RIf>>eSYSfSE#G4B@>ER;Y7QLDW^.aB,c\;,MP(Gcdc=PHC/U-5[ZgaBB
#>G,64QbYEaGD-U9Y)Ed0AA4+?8QLUH-T_Y&0ZKK]9K(2U-2f1-9,K33LHVIBaVU
aWSP61MXaR+L5[@VH9&NTN&2e#Og4b\DEEG))a0JMa<^M/:#2P7c554=.S&0)U#K
Ke,LX0F+Y.a>NCJ&gcOJM-Y9IF#L.LRQW)+b1TV2>+6aLGf&A7LI#H8?aUH2IN,8
CS6_DXaY[NB69]b/-)<P8#F9R(/,TUJU]Q]_UOBWDPL09:TN&:(N;Sf/eU^2?M53
J3fd5>]Oa58V,be;U96M)^+==8-CG5N3H<SXR2A;UbKFA@GgRBfE=9K-8d=NJg72
(ILY::\:<UE-7;S0dfCZOMV#_=V6cUF<??PAE4d=K\>G,JL8P+[9.92:H0dJPJA1
B_g^#VX^BZ(f^L[,5G\1g12B1,7.b):CL30fJ]I3(4HO>aK<=.e),[-E1L#MF=d_
a?P-A>ePB=#[S_cK&/23YT78H?bLN=)BG_c0B[3<U-8;9fCWE[Z5G]4F:)cX=6N,
S[<:2&_=J-?[I18)>#JEXD==g8M3+/:)WZP=g1ZOT_6._V5gPBC.O(ER[dR?NNX<
N<H&Q4dPP<P44FaGP]23.(beJgEOF-LVHeCRZJJ8RD-I9>(+VKZ;L8&X>H;2&f7Q
8M9O>62S7@ZGd0?5[QEI4e9-^FA9L]c3/Q+1f<OV)b=0);=PTAXUYfZ\T6(+H[5F
3;:36RDT3MD/?74#Gb:e()e4d,7><QEeKLA.U;2JcgEP5V-]&VD<<CKZ];?UFC&e
N_a:WV202U][bG<(DAg_:[4\bSS7&ZT&-eG3AQe8/g6fGTgO#AbK1BH94ZSIafK/
+C_C_S93A]@cSXJNY\dF19R]9(^DI]Zc<ZPBN3P_a-/A&=g9YJ+G).?bHFQESH=&
^f4B?WeTIU@IVDV#H+\-.g;MHW&20=_=NL@NFHAPUc;E&;S]e5&&XR60NIg>O))a
Kc955;2^?L0e[ZAM(#4LBWTVT/CaE;Hg+T/Y>U(^P^Ma37Y)3>BcM)ebgg_X@CI<
[Igd>]L/XYW?A2AZ#WJ461P7U1I73Za.[_0&:9;8,Xb2A2EYKd3aCCN3Fd#Y_MX5
ZD,.;b4>UUbG-J:fX^OaXgDM<8OdEJ1KU5ZH:H9#^]G0g_B65C]@CBa)]I<RMADG
S\T3Z##Z&.OTJ#L=[Q_)QVCe[1=fQZ##IF517aBA)f]X2=+&^>IJ93.A7^2:I&V7
]^P^\[963Ud,bd)QU;a\]Cd;V(BVbST<e5.FQe0UPC6^@]K0-[LI_4RR:_PIa+Y#
7d)@.9==[NM[&U\,>b>3C+.4O]2I#,5D\@)Ddd-c@]V;PJ]9OR31KcfOPISVTaND
F<1?7^X-GcOF]MPLaKV+:KBaJA^8](^RQFQBB\aZ_X5:0H_V\J>abb)9?ABDbbB_
c4a.GKL7EZUf)C,02DQ-=RV<ZM>8?QVNRB;SJbLR8/b[GDNS&R[@I\D4GWFaZA31
M6B;TQYT4e33ZWBFb:[\YOM1J3Y;<-@;76>:0bUfQ<4/f3017R)EaH^g/=<C+OU>
:A>6B9^GE-;34WQ+0IAMb/gN=34VDLcIcMeG_,c4Y811=&Z_-P(MN=9Sb]bNOOLL
U;<=\#;e)dZX0B+YT^UW?43FDSd>J9&2dP+A@=.+-aUI;G,\=.D.\,fa]1[_IffR
<bcQ/YY9a9GLW(/X:9Bf&IDg>)9S\CN711/,4bb8:CK?:gODdT]1Bf>?B&IX)_5a
b_.SAd;W<VYdR<2T>&IR05BcH\GC70S/3/#?#ZP;L1H@LeCfg)+d:[#Kc)7,=UgU
@ddCO;/e@GD0a/,b_4FAeGI))EHI+,O=)JP6][UEaI(Qe612:YS\@FIHRgV=d+P(
3RSdO>CTJP5<<Y?7gQLDRYL.>DNg92@^-2SC:594@TXd9FJ,g?/6\DFC#7R&97#0
MaBD>:XPFEO.#Y]J7-WPO2=8QU:3:#),H_RH8GKJE83]dEBM2&eNW)C.U3c?G@5M
eN:M)H&5@&MH>f#1@+#8YVdHd33G<OFYf=5BEY+ZK2GL-BaQ9f46[&egeG1554c#
M/e:8;JCZW,7K&b,I9Y1+bH#1A3YZ#KF__VGQ9d./F-L@Zb\e(#6<WQeWfYSdFMG
N-5f0Z#ag67_feY^DDPK:)VS8BPVa&/CSK:c5B9BR@Q5JG]c;W66N?)+e:U?>(&G
c(+&4dQ&2@NdC65/@N>a#)0KS/PbC(HS^V:O[;JZc62P-,ag@6[N&J]GTNc,K6OS
N-eb9.(3d)DbTV>R=FZ_)[0\2RIEI\FLE11MYZFA:3CY-#53cVWS(1CDP[]2aVW\
?U9EXaDS&PbS<#5:V\[;95bK6?N,&^+AZH2#3MB4>#32YW;?Nf#Y6J\3eR>NP?5Q
dO>?^&M>eH>Q23@Rf=^-/S?C0IKK\@Y<]P=_._,>D4M7Y7[9.7Bb33(XV:);^,<U
6^GF(Z45Z9NE7YLS]E.E9SIQQ/L@9\FJ@AeI<]RH@-@GWL>6@2G:\A0.daRYR#^H
&a;I_bX\faVSX&/5fZ//-6-#CUH;=bHHSWV^EOE](2B8bBd3]<J#ZfN&AB(5CG#5
(NT5eEDM=&,@,f8b3NE<bf@9UI.H8aC+(&eea[UH(1J1c+&S3.3f]).7:@TS15W0
P<QgT4]912T2eHN+V?<GZ:&+IN\5[\UWSQ#g>&?(=<fCU^0gV<<(RH+A/2PZ:3Xg
@Lg0CX#d\1HEX[KFUN)5g9:]cZ\Y<2=[]U&H-N_)7O31_X)F69eFP-)/&N5[K\Yf
J&#&.&XP>8OM7(:J2INZB9Oa9MTJ+c^SUBZ5/-BY&3dX+<c:-e0=g1@+0fI#fH\Y
/;MR=/7Ud#>IgH[6DF;C82#bMA0]#f8;HGMdVb,;^D1LI>.G9O[&2+OFYMQ+(@[f
LO#E[_abWd\QI,WfX=T))&gTTa6--9<5:c?=FaUR._\8TWaQ)>0_&e,RP=I1[8UI
I#H8AQ[C9Ld9F&O2C7]gI45^5A:SVT4G.F1B&]B=RbBf;AS;f1c/K(LXB>Q_4&1O
Y9&R7#5^S_B3aJ]^5V:f1FgQN;^^H8[5Rb64KR:(Scd)@NQ6f>b97Rf/?LCVB+^3
4eAQP.\#eVD#DNdAUdO=c0Wc]cEM1\K00&N+S:\KLMcQ\,_#3)B1P,@Q0O<[X[OZ
3(d]XCBDLe0(O6eTE\G.XB06>bINg-U>\ZEB4]HN1:&=e5G+af&[g87BDf6/>1=#
9B23gRT+)3]48[Nc[^gHUZd6cXN4>+08H3>ZEFQLgB_6<#&PgE,--PUaH4aX>BAc
C:\a4BX?geTSF[UeMSIL\&(f0;;W[^bN04&2[7M?3#]=7&[cF&9S:.ISQe.9N<-D
/0\H5\N5WeGFQ=JD45SGa<AOd&e<6\EM+>DD59Y-eR/28_QO<5R2JdYb>KgYX[8I
5)HffNbfb>2VS]OQg++@b@.,U]:C\LAI:PZS3DH[e3AB[@/\-T5O\3=e8D+UeF22
:+J?f]e]0dJH+Z)LD4eVeK@\2:0G@.MH68:NLLVe:WYNLX2QSYX&A@b(S\QgZNKY
HUJBX:^EG+C@/:G0\UGA,R#<:E#@(4WG<97G37OW:@R&X/PAJ+<TU+U&7,4(2Ga_
S[/_8Oa0UTaS;ZKCS#D],5,eEJF)SYbLS=[M^Z4H]=5/B\R/aIZY<RPI9FK&Ve0=
3=F^&S;_B:FSRLIf=]GP.EJS[41Y@IE#A+S#V2WQWGBEddQSfe[@6:Z(QdZ0N<?e
[e27VUEbEU2169]MN^&RUE^0]#W8Sg]7MQ1VfB(H(A2/I48)GRPGV-cE)\:07JL_
8:.S:)8B7A6=C4,.7@&\-EZ2):46F:bLXN@=6U7CL.H#)8@K82TXJJPR[@[G-8ES
0YV[C0d_>O.K2@XO6&#K(=90N7&43R@ZY,&f]0-;N^6G8.QH87F[]e1E7D&BN3B7
.+SG(d[QeEW@.T;(;6Q?Xd79d+4.23M(e2.E@,6F3N0(J,7[/EfaB9\?HF34D(g@
/,6e/;EQ5e_M7)>MZL2@3)^/4I[RF5_XX)+S4(]8]EK-Z-C#>MO1HdKPa8SH7ZYN
<..8XBMd9DZE@XMT]GQ\7UI7U6F;G#TL6&:\A+Q>43g+#/5V8MESI>^/1gPP-3.4
7>#5#H#8HJHSP7F/)c=K3.VA?.AR)RdN)JYWNP>B4;1X2L569A8dfYZ<0E2S;;/X
JIQYKL:dK7H2@fH@dHgHCg]74fW0TS0]0,E&R>>X>c3^eSWcTUdV7Y\VMg<65Yd.
#f+f,G&bW4&e)^<2MKUeKc^;9&A97YH;;=2N(+,O29GdKQ^2>;-Q[0DY=9LgDJ<[
a>.\9ZWG3O;K/K[:P\J7[UU#aNB=3X\;A+,\\\1Uc14YR6A\[8\^S><00N3D.ZfU
?a5bC,Ief?D3.L=;Q24<e/?V^92LZ<YeT^bYM4QUf[K^DV8Z79?A0bA=O1HHZ?T1
?TO3M\\1ddR[R;GQZd@W]RQae/Ra-eFDR[XfAK/KUgN]#(c[@XJ1g7(81BIUMZJQ
+9UFS?eDJ64C#a48c6J5?(TGgPX73Z+^08bG84JWZ1>-@]?1+(eN6ae+917IXQWS
>WDUE&]\^[YP],e-Nb/Q>RJM2Md;dEGP(FR9X+.,;O_BYd&<US5,8+NK1WXCcbf[
-V.[,I&+cPQa:>@LSABBKB\V:WTSZC6(7aX6fCdNNfH_L=;GT]FUX_0&0#Z[_F2(
6MPDTNa9LEVc^-V\+/?:HG\XUUOGVA&]DGZ+^7M>KWB<g,\[BN8<ESZ@HIN)&OW\
BdY4gNM/Fc-d8?dE1&X+YM,TFY\7+@F=H7\1?A59SA]-;16?#IZA5eH\8<DUE7<C
A@(8f@GBTK6d^MHG6#;H/9:-W^g.c+,2&2[=H[ReH=H)(MF,89E)e31KfB+XTNW[
7(M]AU30/b^HKQ-a8[?e@;b&K(@L9EOK<\<R\ZH0Q&6?@?g8MX<K7T&I<9.eA1OW
7_?5aUKa+^W6<?]-g\BAO4,S,Zb/P0&EH[-GW>dZDcX2FK:U#H02OGQBgJ:dH+IC
#51=885+PKLOVLHGF[RK]aRHX.8B57I5@LRGa^89X(6:+(RDPK]EQ6Y,\(LN9Bb4
QEe-;aFN2M(eUOM4Ub>C=>O8_=FfJG:8YRIBK&.QT?JPZ5_cbQA,,#gS-/(Y>Df&
MS,W?#[<A,?OPLII^)=3]R#+dg+R5X1D7ZN=W\V2?VS9Z/;E<K6C&>30U5I2;P6f
OE+2S0XCQ:T43&;_VZ3MC()_Qa:)S-^KfQ1487G.6(R,<[-#-;(@bRELZ;/R7@gT
2#K3I,TISfG/SG0VGc@/7Cc=L.1/fH1[PO>4[T8A4)O.++,aM565-9KRS0OLRaF>
5C3GT+F0@G#7@JTDN;+=Cb__C^LB0K8N_6]77YX(W4+ZL+IdKX[^C@R,^ZF/QE?d
D.P[9V>-BJ+(T9FCA=J2V(QbM6f^X]A1a3E^HG<>d[8XK7+?@/2>4C-,@Z0MX_2X
6OB2M59@W_@WU#bOB#,M.;H>FW>RPS),0gS\fIZX)WT#Q]H=KB-gQ93I-:<bAN1b
M4=WA69,HW4Eg<441:PZ1/X[,52VB_]6Z;=PZ@[/R+@GKPbX/ZAN^@4N#UcS>XKG
>1.,a-D1g+7Q278fYH.N:O\Z16dJC^S=>?WK?(N7(^RXB_E,./9XU0_JKAb\YbGM
LSUb\Fd]F;\WLR_>O?7K(+IcO\\R^=^M5[)X+e6QASF@5[HVaFS<X)0<A(QE_+O?
K>BM1AW@V74&O_KXN299H/UB@U=d4IP=cWFNYND9E@[?BPZS.4;\U^F2g,Gg/#9Z
G+\_?<)EQW^45Ld0@B8fL)N]>(V6D,/JZ\IQ\B^YN]c4J\S9]WaXDG+Rf;DP(CF0
A<e&Caaaa+2Fce#[EHGC/UPNTBCbTJO&M56ZE/@CPa?d&X&--TT1\a/@f]/Q,G,_
X4/0UBWd2)QZ&)Dde?E^P:\\D+H2DK63YCPFL1H+@/\FZ&JWf.:2Q(42HJ3)CI\-
7,+?TY0@]M>eRUeU-]MH]L4bJCJQ0cA?804M#:_=@_]@Ge2;C0^_KZ1GAQS17&H:
LA9?g#9&Lc7+M5dXeRL/g[]1G]^FNKSa@:aF_XF6+0D(0F@Q@g4;#&.EW?EM7e;[
LbSD]f&OS?L;[[UB:,8GA[KI1;3,:7V9AVV5+QcLWdbgM7)]7(RL@YV>=<#aT7\2
;<OJ:g3J(:62Z\MbV3IUNK,J#P0UUdUeX.9KW]c[?(BQGgWPgPDDefQEH+IJA8R.
-\Ff1J2:]8^,?aaX-Be/XF\-OKZ7K(59252LZ^d?(#@(2dgN4&Wda0L985(DAeRg
V^F9@Qb@.787PcA+7MbBMQdVPT=NC6<Sd0T+eXQ/5d-BXR4Z-2TX#/XDDgK.5(P,
Y>26#J))Z:S-ZUFGeO[>8R3FaaL/HS5d3JEa)Off6@c(BQ&&RV5H[U/gT\364g;6
M;9e2Td__S]46:SEBIHWNO[ZU2RHQ-#>US^W5g&f\N[+@2)S?;03<34+_(-S,<;;
f)QEI4ZFWE(1W\KF2T3KC;?_XBPc]Q[OOCWgcOaMV+_Y86d2MfZK)OE)-.=SU2Hb
YA]VT_;@3OFS1LOCN;T63O.Od>QWaA3/ROKHIS8KYK?M\BN=[3E84EW(,MF]9KcE
eKM2A4?36O8[G5/g(YX#^@a3YLY,f]1<+T)C339P<a(Q?#;eN^T2^\;gOC;>>5NQ
).&IY1IOTUWVZ=8.L7O5:K2R(XNR=3+/ZRDCI<<G4cKYD\_CD+-V&LdX=P7&]Fd]
^d\-JAWd->-T(=\,O?QUD]P3[Ab00?F60S2f_>JeY:Y@N--#APRW=ART+9=DV&29
gP7L#-eJ88@7KYC#(+fL2<3\8K,NZI-S.H,g;@UR9(?BgQNX_fQbO@\53RgDeQbC
4N?;@,)Y4Y)LF]_\eREbbU-E_[P1AbQ10V:SL8.#]MTTQ/dTR=3XV\9^FX]KT?OR
Z:gGVQJD+_g#X9PC;NQ?S3dJcUG>TJN+>3OR;V/9?DUZF-eZI5cC;##4XT,B^;O&
JCd_IJe\]0496.7RDFQ38F_#d\+7?a/=U]&YCC4[<H\W__aFaCLSg)-ZM?2e\W?8
P4GL3F5Ca]#_Y_5IU=a?(.CW-Z&U^:&Z+<@_Y;(;:M_RP=a1[]gY;D7=.7.]F0Z8
6eF#/L^F+I:6)]N>3#D(Z9T:DJf0[Uc?f:A2fE0L-7Z/Q#DH(a(7UF4eKX3L0X,2
Z=.<I0CP;aYf+:5&R6HdeYKAa93#[5@Mb6QIQRgK4f15GJBDTK7Wf>+#]eF^[BEX
KX8RTJS>bO0[I8&#@(7d:AB6YS/8gO8712@N7\Z>Y8<&eFIGCG2?(ZB,d\Z]P4P]
b&F_T,f(MY6b)GM(MC\Ice1N>Be>dES?IF9@7f7H?/YAFdK#^?]dUG[NF87XGS7,
Va<\II/BP3]f_DJV>GTK+=_+W^D6F(S:WIa6^]JZYY=[DGWA_@CGFYeY48^VJY5H
a6:b=d],_1WSeU#<X=dOKNKe7P10=J<DN5_G>X3IU1&Z3FBL3Z1E-;PMUBB#>FRC
ZLH46DX4K+e#+SP(6<>=B67PWF2])-C#.=FdXR2Yff;74?Qa9\8DK1>daZ)gN407
U8G2];CP=0U:C^^=TcM7RF]a5<Dcg(W@g-\-(9KP7T_F9f7-_YD)3U3ND_]R?d/P
bR_8;S3-E5U>1Q&7TM/,/C2dQ&XI&\=K)@AG3fPMS0IE<J=GUV41_;5QI]C&NUe#
F&Q<-UNUNM<Q>MU/?+F2DSbZVPZ91e[?bT,V<J)_^C:d+.00H=WJ4[f1fDR;Vc\7
AOd:]@,DLERBU6/6EgdfWX4@-(2Q,),(MN.BN)T[Z/-a]&+.BJ6QAZ9703#cM;P_
93Lg&;\b&-DB2#Q[GNM=56\[07AQXGLSaNRG2KYJdg-ce&1=LfOIOHLHL>XC:Qdd
c^SL8)a5CP(KR6WS1Q)(^](55Wa#,4^<J7)cT;@97<FA+2GPa_CD==JJEgU+&9CX
TPf7,398YN]A0/AALFD[0;I6/>@S=,d6KJ[RKc(,e8eaHJ4J[OASXeZ+D(I5X=aH
a\f0:=HGOD.:>c1BY(>S_&gTE<G:XK+78(?LfMd,7R4TH@,KQ#(\a[T\QY0L-A##
Fa)ACM2;LC4+dT+KVN2]-eQf7:(beCIVE>?D;):S]:N+ERKQZ\=OYa-D4CWL5[S?
ZM&R:0EBI[QAe@PbAT@3P?><=TBO0aZZf?H),aDN_L@,Jge_PI+e&gN(@<7G12Zf
5R@KK?^NA-IUG24^5+;8Z:OTC8855Ka9LTb08f]eA@+CDUTc9KRgE->RWAK(^<gF
)Hd&<YYH^E,AUTB._AVFP@XdS1K2;\9UeXZ.dSN)GDH8.5PA3]29\E?QQfWeI=_Z
E(YAR)IC@YWKNgQ07]5,5VY300MWB5^UY/C4YHB[+4_/G8FW#-b9#.2P2;>ebL4S
4WOWG8/Ta[<eK.([.b>T18IC];_\dQ@A0?5?E=eS&#-_OR?OgC[bPa]99YG&D0e3
I\^7c-L[_f5bV7-HN__ZB=dPHc2HAELT&D83b(^H:9E+=:7&81:Q/L38M)I?ReWf
4Pce3@e;XOTI:EF\_OeHgAH9GRZS^Q0e1#1M9Na9P-V;g]&X&Ze+M6a0&@3;SQQ\
I2F[]F4W#MWCd5^>V;6[gI1[GGg[8=\:EYLAH_Y2Dg3:LPd5Hc/dU:1C=I@DTV8Y
ZYeCJPXFJ9W[g^:&Tc)BL9E&S7][aRH[K?&U<]X+)ddDOMZ2[8H?;6^Dc>O&&#)O
@;eO8cI/fC)2027(UL,JaC;0b6&P7MKF\-,KaKQ3SYTa0]&A=:P>(;AHeW](W<b\
V5A5b5_AQ8g@\&SW0[([KW/J50JF7KdC#IN_&NF8YF,gI;R)GV5a@&N2^YU;8JW9
TM6.XWR_/YC]Ad7(T=aR6aQMS6/7]V_F7,LEW-QW=Vc++X&DYaDb\1g-@&g<7ZO^
A-1#HL/aeQX#]F\Ld/7+GI0\+UAK6VE7fFS@5E8@G0\g:8Q.C6GWXcUbd:f#AaU<
f34fCYJfc\Ae&g03..40,FCA)//BeHbHWbK18XXg[S64FB3]2J<PSW_:E,X6X>Ge
GXgU[Wa^DdT98I-ZJG&1;XceD?(5SbZ#ZR\E-AJ5]I^Z2FX8?Z#cL-65N\3Bb&G5
IUHF[2?Z<bB.(0H6ZB#P5g;>RUZ5M#I(/CgWQX-G9[8FHeT9&R:UI9b7<DH_OC.-
d#d88a]HAPI:#XB\1RB\?SIZAfZa/\AC4DY84dAL+&X;[[U[efZ22c#_Z^N=L6a4
/]T3^<26g8<DU33,aHV=bOQ+U>@->(6AXQ,(LfNYS7cV2eM\1db^M5:QCW30?N79
bJYH?U-IdW,=5A9NEY2HKJI[+Jda+][IR9Ldd&9(WX&#gd-gIO67?5W>baOQY3RQ
;e8BP<<#O/6A>dXV2R<c]VC:?:Q)S^)Zc?a+LgEUS)-ZM?EW66.B@XdMdN6/4Q_H
ZJQe1:/gbN.YKJQ/gW.:H/)2c^:;ZG=R1gG(,;D#PR-J[O>Ge9.6N5NZ:)aB0O?>
DDe,-0:IFZW/PA#\e72g_c):LC3&S5.&TVS?FLR;;WM>\D9EOG+/AWa:UEZI2.9D
-?5)44X)(aNXH--8_-dD3^03#+J,X(\f:G=cK60:EGK]WH04RP+)X-Zd.KR^>Xb2
RM\3G6c:#c4C<M0KLKI:=e6(1>XJAL<3<\d3T69-/:?\WdZ?Sg?QYb2bC&,)TEIH
gH-c/DE.\T\7<FKR=.QFB.RENe6EI&9#2,IAPFHHZCg+D]&[;0P@UaV0\]V5X8[B
Y;M);O#K;F7516EM7K\15b,db+1c+]<=V4>#X(F[g]#8,J2S/]G6.6V4dfLb;L4#
fUGeF+MBV:BB=-==X:M@ab+UL+d4<J6g@/0a#;X#SID:f]-/II-8)B4g34<O(RaG
2M/b.0V,ON[^7_H4F<1=W66C+6O?OBL:.[[G@Y=VU1:f0/8BVa3&BH5R6ANg_>]@
g3EU.TO09^#SaASM4AR&4DIWKIDSZU4-6<]I?[R9>=5B5&1>]72Wd[R_#e#T=A_Q
^AB?PCG11e8a4:]I7&XF[Q5TNG0MN0fE>XI7O28/3#E<LcdgIUYca(?a_I7&>P4?
.\.GM_4^M?ND#2?C?7b&NU-^U(6[I;^SLT693,S4Gb+X/4,77.]4>;6W_T.-0f9X
HZ&6A2LU(W2NZO@P^7?^g^U.<[3/DL^0H;aL#>efNf#:cb<S:VM^B7?d]CK=J#FC
XGC6PHPM[V00ec=<e7,a?R4CJaJXO9eP=\>_UaR9A^A6SZHbK>WTLZ^<1(XHMEC+
gJK(2BcRR,E<f#^f(0(A7Oe#g8-OHe\-,02f?,LHe^AB,[];=b]6/BT/bRE+V+NQ
C.F^=\7LB^M]E.A/;V_K3a4@+a[0:_J&)[WA@?EaZ3P->_gEB0D[+5;20[MDOL@G
[fO8/ZJ5O0K;K,@3P9<7e]/a_b-^Y\fSY-9?_Ge^+QR4I>@Ee<d]c8SD5,(&[Fb:
G?(0VYd,C22g<_VJBED78#[@EW9VCN.6W=[gIIdb,1,0-fXebK,QAJF2L,/(Gc</
M5RF&15ET7ZY<0Dd>JfEMP5L6_-@FX(?TNT&\S=;Qb)]cQ5#?6O5<TLG[[-DAQ9N
#=,2>MdH2H:Y35<HIgN(\YK#:aAGbVR;>3])P@fZ<7E7#5cA_,ZA(;]TB2Q9T+7=
9)LTAE9DXNQ_>21&?[7_(5Ee6Y7VFW-06+_7BPd:b=WB0[ZLCd<R0Y0;fU=JNI#L
F><cG7/g<3VC&GbJZg4g9V.CdP)FSOOG>I)0I#-Yc?X7K7^S(W8J)\f(6=NY5DQb
=R;<G=c3;GQLOFO7:@^;GaS\D(4+@VC(PDOD54_&9Y<:RA?S0>1JO->PD0d&O<DB
-UU^gIQ+-/HFUc9TfLcd@=\S>6:ca3@2&^CYI>9bb5gGaNVc=7+F(]NfQI,.S=^L
R1OgG<MPaS[_4RT,C9JIU48W\2@HCc.?D^5D1Z\\JYcS?_KSNb>@<TV)_5,]7Kf(
5,bPP.M@W]PW@f3TE^KS;314>5;FX-YgL\L]X,A96F[KQbY[-PQ64fL]1HMU4;gb
M;2#e7/Gc#+-OGAEF8:7@?d[K_?CDTDR.BD;;Ec-OcN[-Y67Z<I7JcGL(b;Ue7/O
YB(:gX>]GWN=(e-P:9MD-I1WM+DZYY[4,?@A7d,Y73&OPUNHZP^MP7#YaL=JJ9(<
^_a;SE8aHQS:^Y0ERP9[^aI..Z\0E(PF?F^C7S\+RJ)O;,aJ4Z\H&,]O>/:93Q+L
0ZV5BPF0)SCE8d13AHS)5aGg/I+[U.-3[dgWg6/I>T]4fRQa905&A.ABX+DU/bV:
8MMN2g.T17O7?-DJ-PRLf<a\D=HMXD-;bHN=PId[BN^]8,HO)2_;/W/=IT_<VZ.g
I0P#7433d7#B:9R>dLHaDG#7bB,Y.gEB<>aRLe4U(aKb2J8HP393@CQ[8RCc7[KW
[c8KVA,_DM@NN+8HHS5H)Y^&-)>K>-U;b77&_IY?<R7CJ6\3-:04A0gY_C&7&8df
eI8WXQK=1&DF\bO4b\Q.]1=B)ceA@N4^V9fNM]SJ3O7=gMd>4VJg/5[Y@8^E.>;c
07VF.S?[&N_T-E&Q/B#+5P]0g.AE7K]?7Y:2Jg=PV1B/1YMNR:QF>,8NCc27&PaO
Vf))#A\&>@f&&740P]XMF-&@;-10C((^SYX(6K.U#P,MB@H@[Q,SPfcUD1#H8#OC
Y]N=4UVGFDf1e,TbJ)Y8<14^9C<Wc8S)XfTgCK(>J_FgL9W>4TIK_8I:RZ2<6D#P
9^#O;g-3K>-[@RHdQU>dX;@-+&Y?^.CH+\OfgbJ^Y:8f-K/?DE0S&.a&C[gUV<5^
S]&Y2]KM-A[:5gfNFKLHS2eFW@7Kc),(KE4T2^^ddJcIX=8K5SCEFU/5ff(eD.;\
,T&@gb>9-g6)]IZSM>+N4#bB<LB<,?SY<4EU+(9a\eIPGQEKe6Id.R[^GF4f(+3.
=;^-0>>&NeRD1Q4_=EaY?W&A>BC-9b68ND_5H3ZDD]Pa,>\^<IH4N.@;FY<G);#,
?RdYC)=1B[Wf)(Y>@g)6UN6M[92@eG:I?FO,TBSfG-H<A]-=@WMc@G@ac.8Q]H\K
WUeY067B6ZZ[4U(D1OE(5W5(VSU#>CgABPCUK#+WAbgFTTF&/6IP^=eJVa\K-/?R
28f4f>]P6=ZY?[Pdfd3GKM4Tf))+G>V>&06_XFKI>)V1YKQ0J85XX==:b7Ea+g?&
@E2?#/;30BK3&U/\0DY2TBba<48RDgSF7V?C];#8FU+1.N0b\&P5N^=.<\Bc.G>W
3<=0PTEA(;N9)=5DE1-9?bN?0AG<,I#TGf703?0SRU1._T&XCP&4)9RC+\7G6[XV
O3(@>c\.I81J48Gb1H6AHW+\1RW,8XG:L?8+R<-I1G/FNVQ:fSSW-Lb1cE0&C.Y?
IGKAbM<[YBbgG#=MWKb16+(Z@LMF@?5^W6P/b[N=#,]_12aED]A\BVU27gNKIG\@
M]2.XdWe@\^YT(fJASWdQ1OM2@4g>J=M0?B,\C4a)5+a+2_,TH;2b+b7JdOV?6V7
/dVg7ccFa9BQY,+4_cY(E]1X9B]S4BL7]0E6@P4IV]<f)Y5;a9L^I^GDK8CB9dDW
&/=-3D5/-[([GG<(1K9F7OG3N4LaCf;eO\[GMTdW(<>/)a?4d)KH8Ne<VGb#8ZbK
^cM93SZWKURMcK]XNe^G#a,\4Y1X5C_/H6eHEA>\Uf7CUM&d\SXFW1gY,_L/.@N<
#<e6U3d?9TXC@W2BF/[/V^JP)_SDML+AEZ/S6g)QS(&<DH7^HG7/:>H7]1MY(e39
2L#^+/7d#.5Bc8&(N387Wg_EgJC\fBAGE0a2B92P3W\#@Z,_3]@LX-fZH72WLbg0
V;FNUX?32K2LbWVJMZEZ]@,Lb6EUX(UQ(T35bE61&WRN7O::A,5>L5B&0e.K:EW6
)A_&2;e:GaOH>#I3;9SN7LbOHZcYeEJ[TRQ#Uf--3a\g\??5K@0ZWK?@JWbb3A1/
_MXNbSb(6MS#:XVU;BY;-UeT-AS0XdcGW>N8:BFBH+cGE8HLb2dR[11DDJd&6G?b
f32W<3^b<@NdNC37\VB1\_4)]Z[#VF1V.7[+SY0dQOHT9S_(O;>BBE-)d0@N;&OP
4<GF=Pc[5Oe;\R#G0O_N>(R4aL;]7:Q&#74)gE:+<e/&9\?(XKb_YM#7E4;I2c@c
BU@.5P1;_fA<>Oc8N-K?;@)9\_ES1C68B]\1eYZ;.P8=Q#LA2d6Jg>BDXD]#V4G3
V9@LL6,b./ZMCSV^5f/4KEVa?<10LBeX3Kd^YWE.]e2(=F->SEcIS)3X-c5YZDPE
37dVQVY:AeZ&fBSS:CEdQLbc=4<6;;BJ>@VN&16A,F--\IGT/PMGA45VG[eC-XLQ
c1cO8Q9,H)_I8R\/1-DWZRbE.YU@8WZ3PSJZ2@KJ0XbD]RX\I5OgQ88HPWUa#80M
SQ3J-+4>2-0SHg@9;OG_T6UFG6ce;\c5_=>b<b8N/T]5DbbQ;:c:.KA4UV9&#@0Z
,E(6.Z<)<^eQ.)-2WK.@6Xd<#8?]fHf_;?#]1X=/WS<;W=N(T5_1B19Jg=^V5PR[
L?T?-2F7TBbVFP-UaF,AE\(A&H&>KgR59.AN0G&e_)/D;3JQ@?BB-&YJGc<+MOCM
b>L;840WHA?I>SE1,><e9;&YIP;+>F@:N/QKDFI56)6@-Z\F_R?EE3--MgdfZA(P
EV+VeDb7]-1W7DQF),SedaQW:H_)C=AZJbQ1(..[>PUP]>dK9VUY0H4?RT?=1EeB
?&D-:BRZ>+I=Ff#F&9AE3+:FYZ,Q778ZG&I<TMg=.HD[Q5N6gRb5]f.91[E6d6Z6
LLY?.5JN&dP1((VcDJ_^MDY=(](,I2K\ZQXPH2/bQHg=B:M^J3]VH\>F\+AUUF=b
9BF?,g4P\E-TO>-;_FM10[(,4gWafT?X8]/cZ;e53C/T:T/QHg:NIO:dMGaE^(BT
D>&3F.2DRW)K1OWSL;BSVC.R5dP98,U:M70,:75^=^K/PYB<agV6=/#4b7G-cQ?C
6WO@X/XO7>ZI.9@Lb12+#H>>[Lb1LUUCd+H@3;#R<(UG6DaW>&03ffG.WC6)WfQV
N?B<B1D##e]FY)Ga+I[bHO<aQeY:36^cZfN#(B4@O>\>R1bf7IXbU<(aQ4Facd:&
1),XUIBf72X>K-#;/(Q^AM^#bBP-U_Z8L;Z6SHD-EUKbZVS=JF7aMP^D2RZbD^JU
0,/V):J:5.ZJQ#,Ae\6:>B-F5aU/U[RU\6C(Xb320IF3D/>IXU/_b;C(P/X,O:-X
>7>>30Rd6&PYOOS)eK)@0AeJ2]GW/M,3K@-&6O4QX]NKJf&(BQaQUQ>YVU)-</0)
g:e2#AeCXeQ?V@H&/Ja5_6D5]^@6<CS6]]J(-TM2\OfcFe+MY#gEa[SJJL-754bU
e:/4dfFJ>S1(<9dFC8G;/=7LI-PT=:N_7D4Zc5,S/\>&Vg(ZT::^=(3[@93+:TPL
>dC55=DP(YR[IFS8YVJSO-JBYH7]?.;+8Z=JLc^g9Ya2TBGd@EMY-T/7e8L[M@.-
WIZ9X(0?S\ge?Reg]Xa=>CUYU]N<=;^_7,dAR0S-=)BY)](_]R(DH:DEW/4(O#Ce
8VYBGCG>1B1-LFSLTLO285GW@3W=PH><LCSMA#_VeS^3A9/@Y3GW_N>gBG-3_WX\
DT31I:afN/2U1)E-&/Z#Q==[#6;=.H5CI-@U#5NH\:I=H:NddEU#0_DFOfL@K9?6
VL2e;9WG@J3F6]a,,X&+C5#(dO,CMa7>+afV9AA+V(R=R8JN=b3&IR<5CY(TD4Q#
C2cTSP;bRFY=aOWIZG_D4^[7e-#Yd7M\T+=aE:2(XcdMR^W54]g+RXVZCcM)dYWT
Be-?8.4MK_2Y_>>R5cd)&3Nc/A\2&7aU<1DQQS=.PCIE5P6GgYI&V)?IcALZD/9Y
e]/T2QcT1XMX9:a:U+./3F0d+G0G0SW9AdKPII\c@[EORM5cL>4E5bE>].#QYO;&
3WBVTPHFZZ<7\3cPQEO9+H(f91Xa)9YPOU>Zb?KE36>g5PLHcb79P.AVX;CfQYee
DVW;.2LcKM79<U^>Z;SgYddEAUD,d)^feBV2d;/XGg#V;#CPZEH6FgRCFEY@<C;E
\H0I)RWBcKK>XG]d4XLK\,HSZ?bT7F]O3dYAL5g,33\RR-:N=7RSZP-<N]aWS+3>
AY<gJS.,CG=N?M=M,@]g0KR[(6ed^7SUOTR7S[2T0Q:]7&#5ae0/FRA<Ic[=CHRe
^.KAdJ8?LLS(_^gS?IYeTKfZL5&Mb;)XW\=#I^]FLbd;a#F5OZF;\<>f]HT_8[2J
.9WcAA.:#TZ>G=b(eG8Q2SIdHVB=#ZB3YaHZP\@gH)Ob(3Y;\d@1C.]U:_ca7P>F
D@85[W<+a&S)BW1[6/ZV0LbR)JPV/.S^L\15E2=JHfI1RH7_93\IFUH26WE9CO]X
dYMCL5H)[PcD)fHPW4F;^,F+bc^;PH2feA)0CB4?d;)+EO#V)]>7\-_92\DPH94(
[RL_gX-/OIP^\T7JT)9U[Z?;E;6RaRe6b)Z@0;U6:2C6B0WS/I(B)6(KB:JK@\g#
Q8,5T\8DfNDMU&-cY.-7a5e>H=-\N66]TU\aOO92I2b7dJT03?@FU)>UP3@A08b;
3-b9W(d+2F:TRbE>MOgZI[UTOe)9eBd]9acY996#;DH\5J<HPBg0?Q?d8=^MC;d[
[DRSB\/\WNZ+=L0gL]AS\3dP.(3MN?5/)(\F-MW2B8+eJXGGUB1FO_\U1Z\/\:5?
8LW^G[->@gK7SEG-c9_Z@b7D(:U4-8@G4:VY(A\6bKN&f_F\OOU-(bI;8He]9^e1
GW[1UCU/GK4Z^NQ^WIXXASRNL7IL\(5?(GF\G\ISVM.S;Pbd)BRTf#g<..\aC):S
O9/UVQf:DSQ0)P<+<.\#UD3bLVaM^3N@4G1^EO.FbLMH1a351(4a@I><1WE:;/&d
a(^f7gcb;bNC)@GVTQ_TIDE;CIc-\->KB864P1ZHgIQ^L?&\2S:=L]HCRfPJ6:J:
]FAe+1NXD]Z,(>]F-87;08PIfG@J<C.c#aU@U.[DUYDR;eX5a;^J_:YHGa)XA5<=
AU?c<XN?7PN5Q--_I(61_0^?-<6cP1^=^DW4ZKU@&H:P=G1b9_#1+b[XPEb;70LF
-R=bQ0dZWL+IEKV8;McP/X[[U:dT3>WC7#[+G/QYV\E]14:BT23eT<HHRggA45MY
&6?.IV;7aQUe<c\T1baRFK,]g.F=>?#LeZF@^F&7X99<:NaUa\,J@4S>c^VX7B8F
<fPdcNbGH\bKa1<cN1&>_3)-LZ)8L@6R5OZ=[>2bSMBC6&DPY<7MZ7K)7TC>W>Qe
6#.ba8aO&/;^XQBc61N&=0[JQeE3YMd^CS()\<dIL:Q)>U003S,Wf+.dI+1.Jg\B
gUKX/OV=cf]5C=LSWC@VX=PINB(/3AI5dY8;?Xc1U5<I&]9gQ;7Oe.d?RW-9EPUA
=\Q();B?Ia#[4=_(a6@>,7PCC?HPIC@^fNRN6G<GFC[1A_64Nb#He5Tg&-6,1E1E
R6.U>Wa7U.93MPbV>A#G7a8=bb9ZdRcSb5(LP^&KWg2)BI@/:>F8>:)Nd>X2NE^F
1aEVPYS2eITY/;U;7[M.DBa@6&a_Z92KZD?bc<S.SE::JcbTcH1^6/ENW0^d-UQ(
24/3P87JPU6)\(SC5W11U,cBbK?GFD]Q]1S^_<(JIXNNUd[;Z)PBb^>6KCZcbG=R
KV(6V5fW?56DSWWe&fW,CcC^RZ7#F-f,J-+.,d.D,a\<\JH@\5.G:Hbb1+/2K_^,
>HZB3,D2>5..Bb[2A78.P@GB=GEQ(GJTTAO1dSfZRTg:>bQ(X+)EBQNa]8cXFaMF
(;\=b,C3DFWHIb3V7e=^]A,5J+<(fC4fB_AY0],1XL;>_cg3&SQPG14=]?,LVK8,
[<TG_fNbC_\]gOR#K\_XdT.MRC5bS5+:?)K:-;>8?R/4f3325N;&KOF\(XP:#^68
?+bR_T],e<+B=&,P3S^65A]B.@Dab;T+N3WZ<V<=P78B&ZPTbgH1[P&H0Ha()fD0
@cQ6:[=E:F7dX:gb_/dSAT7efOU99GFFP:Mc40;6EaT6=IJ80P@):@@5dD@H#3,\
AF^>+/C)LW=,-LBHbAX>FMdGO@8^E^JPAP>QeBA6;?OcA-\Q_1ON[,^e\C,R=U?/
TA_]H=12AGXS[&F1GJDg.).+QTHbM_8(::;EZVAL3eEQLNBN?G?Kb+2H?f:^W89e
]@[:1B.]OfR6<R<F])6>--Z4?W[7J/^PWRWcN.@;Q:0T7(=5+&QOaeQb,/>/\,CO
L\2H.9/(B@5[YFVJ-7#?Y-)+2&3e>(F\3<(Af+PaSD^,76P:P-6e^]8B[I,TTDb^
+a3Qd&gc?fN]55^K_(c]0V4@H+c?\@JP60X8#;/^X@B3\LLIR8XBT13g5/>YN9[d
eBI2]9.?c2I@_M[]0Kb:bC\a;:Z)67f<U_-bD6cK,UQRA:L]NL[2:Z8a,X4\&?L&
GdPFR92]IHUT4;+4S2JN;3BGgYb_25+@&1<I#?B]cHJOGK,_X[<Kf<Of3FBfcH\J
^cOI[0ea2Ga9W07FD;[g&L?I8D:X,I6;[]4QF5U2f=><V03TQaL::AJ<@SWN+6(g
dLPW[-abe?<8N^7?e=4#-;bZ4OIEcd#9_NaHgJ[7GBQ+CMOa]]K.+>?:d<#?:+DU
&BB6e239#BTTTTSdUF,;[IV;;K/_>?K:S1H?8F.3E@Q@Qc)E2YC.F<VN[]>I0=c/
R+0ZUMQd?A:EPY8[P6(Y+B41K/be:\-b?7LMFK5A/7g?&bZ@AUV]@X4d@A&=-a\W
1:QJ=b>F(IQ2VEVZV.T#^#]I<O+[^REQIJ22@aOPS;0C,N6/V?YTAET7NG)S(QZ+
bdd(0M]N?FDbRLf_]Z8N87M07Y3Za<+BQ)I_&1\<g)b5c_e8.(&J>2O,@Ic>HCD+
4gd;-M8gD>c[4A(:YDD-<TI/+We5[]4OOPI0)L3Q8(Z5^MQ<.[.,1Z7;,/@eC=5[
412g#NW?F+/D(_5B7KLB2T4P=A0F=0HLF4[==cF\WR0XO7QTW6=/DJ0U]::9\=Hb
W\A2Ra#DZ,Y9(UcGXFUFN\?33<GHCYBaZ55^;70?b-/0cQ>LXFY0^8UW:K<DJ_IE
P^#U?;_Zgd7QAMXg5KG0^H-[=.)Ce^=8G,U>32c8:TJfeLO[dH\DAOC0J&^JH;^V
3/7,g[]P5>93g>M>B+_FB/DTOKP;D+@GND?DS#ZAJNe?II@+Z5O5bO/(,]Lb:E9P
B-23+(+ON=:b8QNY/&5@XHG-U[NN(ESX.c_I)3D=X,D4,?8;ZUH5N/H;7<6RB&ZJ
\AJ=8D?USQ,1(Ib^T88[cS7ST._4[JB++aR^DY_cBc6#ROKO)[c<N-+V-fdTLK@W
@M5RL6eV9c+R8L6XB,MD68,M6?;,MUB.\>=D_3^988P7,KZ#.K2CPRT#(=-?BIS]
ZVAY_3Pe7_eH@XX_FG>Y98LJQE?#NOAX+Wb0U<IXIJA;<.)Q8C\4UGC;N6?XN[dS
^-cG(#C<W;,,aC^PO#g^2-[VbcX-Ma\C2W_cAT8R:::OYKT=TPY1,aeO^VN7;D8?
aA2K847KL_YE^7:I>(=HJfT(#(2ZX7,=(T(B4ZBQRDAZZJ\VJX]D3MBS;/0A6HW>
-bZP8Z?=O02.J7/H?3B4#b,fCBQN&5Q[YJWEBED+=gaI,<&4MEZTRgCI&?X++;##
F<F1CfcAcHL?f([>O3TM)O=#A^8FYS@V@#]=J30PWIW.4JJCWO2T_5BX[/g9cbaC
:WN)/1LLBZ8LB\WW@NOW)9N_^:Z]_US7B4AG3+>XM&^<?GdQ8L6JdaJbgV^J:ESa
>J3ZJ6c#EO9\8(;B\:L\AeY9&Eda1>0GB:0f<Y)W?AL?dCM,HeAWXH\X42eS<S-V
U=>@]FNL(^fL<gOQf\2?]_-U+,QEZCe-b#EcV@eH_Y#.VKHaAPQ9H5cXYL-5Q?Z@
#78AgZ#;9D<U#ZYTE=Z(@^E63;#D)bUY^VY:cVFA5Q@EL1QI0R?M@d+d&#f;5OfH
-FA;7I>,-/5OUF>6D;IH\.Jf4dOPg<ZBOU#_YM]];a(YX7AT/2=F?QS7=7RB<C7L
]I-P[9cc6C#^O,U@>+W7a6=B5\d_P1O6/YP6)>2Y0G[(bB5/^b+Y-PS0U-B)aGUf
QEA)P:?/ce0M7a]0KE6I[R>79)F?F\02UI0Tce2.^#YRA=?+CcC&=R,P,;M73Z^>
3\Y)NIO&H(.+35L&eK\[K(K5A-;MK4A;B94V#0[<,9]./IW[0WL]b;1:gT=^O<-]
U.N3^^@VT>IQTDB@\I8V8A7[S8Ub(f+UAL,E5LPP3e:>BTbSVA<2.eY/1A#Te2Yc
HDGDRQT,P#gB[S<F./.JJ28U=)SU&ISd3#PN52/)6GDUZS,,NN\03C\S>X6+Z5H(
/Xg4\H<(K94J>eNef@[XTB:_<:RW9NP?VdP;[VS+:a15]MRaAADGfVA6X,3V.R0C
gYZg_,&PMI(HLE=@19)Y-E4I>55QO6\JSSR/4^.O40-3UT.E0@-G@0\SaI[=#=C?
3&@a;6BU-P+;NG>J74Q=X^:C3A/f0-e.,bLfFM.d=,JGdKAK7H0+/)J,GbLE3]WU
#4BPQ?DAO>+d]I]4>?_a44A#2?JXAALdUSW,cX3EVO#7]a9;b\=Oc4K6/+SDO93Z
@FEc,KX]Xa^,a,W<CfggEK_R)SJ:;+(1S=TMg,Ff?4S<^G2(&+Ie6Xe]5T2,,(]0
C/;#T:IJZc6<2.Vd-d,[<>e>(5[<)LaGA5YQ/U(MgI8PC;gWF//S,e>+C0GXKZEK
b>^V=.I4.=c#+4S?)e#<<cDG7B9acdZQ8A?HUFV8_eJSU[e^I/.HZ<@e0(=e,LIT
bRVaPH=X0L])NRMQ&OQ,VV#U(3^,+6HK3;G<[8@YTW;6>fI)c9O,:\M9O3&+B\fU
AdJ)+<QVAHSf/+(_<V>PPR-X?:5,TT.#?1Vf?V.8OVM(.)UP0MG1F,_Z^,6#<4#V
?IWV-f312cK5B2S&G1L0>EOaOHP/.VPLYgEB(fI7C=V6<,F?\XD#ND.gSa]g:JV^
+CUaL00H]RA3R.DD7<>Q+[XVZO=cEa[7<VBRN\RcG&.X6<J+]2a1[bg>GILK@FIZ
N(WD5,LB7<a;_?4@b+#dZFdMV8X6)CB3N43d+EL;/RE9L_d+Ra[&FF_^.A2Lb_Y4
2Lc=W<H)O&);[Ud3]b/RHSEBX3VO&95^)?G^bWJJ3P9a@_bA:f&(U9/R=V]^?#cJ
F-R:(ef9cTB^]c;CS(VE-X&BB\NMJ1Y(bM=F\&U,96^E^X.b>?:f4FL_J(->I\E#
<Z3L,#JJ7L<TA9>^GZ+I4^6HGD@RBFN5c:=<aO7dUQ8C4TWU&G81[.=5g;SB0/)g
79a-TKZAZF8AL1HY\(JBIKLLM^DVOY[J[Ba)#7YUZ]KN4LE=27a&VG[K2+5_b0H#
P;cH:F;_Q&G5)-gCRM;HgVa<+CFL/]FTI&(e1G)WV(+]793;f[,AR<KbC:JIFYV?
e>7O<JCB2__0L7dQ@1LHbBZ;@,=.?/QKK92D?_H3X#^\/?]]/1K>eN#_]M3XNXg[
]>AZ+JSB;f;L@?&Ue./eLAX24?::^IcU&5VUO59C77DPbC>b1O<-R[/BCWK+&6]A
fd9LYC<bcY+G0Zb15Xc2&2KM(dg6X?4MC9B\37d)9DLMAW6HPEZJJe[TBE#LYC,B
R8N63\;\FOARFc::IG2G/f3UK]FGI0SV\\/[7+^659ULM0AM(NPagBX,7U+6N[]S
S&.gTAg0&KNI=D?geMO>MaSdVY#;;0&-T@&XbUHG@bQ(7K<a64F6+L5G(ag6aK++
^O[/@P41A4Ud)B&UgQ(##039OJ;0AO8ea5G^?]BQN2XFePR)V_e8Mg0,DNT[8Z7J
57AU:9Z>IC^9b[d@3Y416#8eNMWf)(=L.[b)I(;;9a+<a9+LgL06^0]#WX;^86EV
W6Q2;cVK:]G<EEU)V/b(JB](FI+R60=#[(fg0+)_ARd\Z^Id8c88U]GfNBP[:Z>>
E(&R0-F(V(AXDYFYATWZBb<,B8BEKR0/O]69P\PdFH6C_DE;\.<JV&BXTN?9daN,
JE)+M,@]+3A:XD7O>-Ue4>[^&#69J\b\DML]KNVL9PL>Z^0=17#]EVQF>_?e>+/0
3O=6=^aK/AMJ,:\]=JL8gO5E0.HY)d8;D435JeJ#@4E4O<6)N&1AZV>&;=\&?cTA
da6-(1CB1cK1>ab^=()&JYNP7Y4Y.gL)e^]89[<D:NXLZ9@=]8dbRZ7\<.1X49W4
8>;OWDe+7PLQ73\Z^Y+Ud1#XRWWK=Tb/@e:=V7P\N<)g[QHb[CVI[GLJ_(6B>?67
(DF:DD;4>:UcXC9c@3X^^3AIEL_M1<SA\Bb)GA4g9O9:DK0&d8L=JI74@7Yc4f1D
7gV&96(NLeV9e@UIg=4f0g--=#d2ZBB2cF:<Q(^,//75MBIPFAL)Dd/:P=OJ8DTT
g\,(f3QM3V7Y-3J:71f/Pg+/3G3MO5(7/(?,1ZU4=.[?+X,CT;1dDJTCXJfNF+/1
-91BD.@R.@XHdU56(I320]1E[?,WZO:AeI<N^H:76A?/L2977_/(0+Gb0cIKBS+g
FbJZg@fJa#IG[PC=897-DC#O\)D[Y<(TIPe8B<?+fALX&Y#@@:I1FUZP4B2+64R[
7O;O4X[B-5EN.-5@IfU:U<Za?(.U]G)#J\@5J-=E-<1N/,W3:?bKISVMQO&4:RWC
-RP[I+[8XV_R2U,Z&_RB/<QZKKT&Y1@J2cNQMMILT2EbW3OIN_9VS1L+:W_&4,eI
_-eE1E58b#(ZMX]B,bQXK14eX6_=B<g;N<QY2YXI6Z+U;VQ00e)Z^EXUCZX+Q/=U
M6@d/T/?3U2d&FfM:>]1QdY^6GaLE28CdIDFOVSZ9<6bT)aP]c@TW<+NCe,C3+NZ
UY?d5#V&bC?1NI\/;dCY)c4^K5BH]-?T.B1?-O)0FA&)VM)2H^dH5)/FI&f5/_XU
8RDK3DD>@W@H_/[I=8WT-#c&M<?OgW9<.:Z0PSRBMHA4CMDb9+>/[42=42D(AIb)
XI:T2IF/VKEAMdBPCGKP1?]5Tb>4)HD(3_(34GSB;;>@VUP7>C,9fBDNO;Z\a+_S
TH2S;-F]/S=@<)DW>IefWe5@ZbcXFE5@1/Y<57YSAD(Z/>0O]A591ZF6cT7=?>(W
)Oe6@7d^X]M^3U7GMRU5gIO<#KZK5(B](:/ff[&78>\E)/8P-,NUJeR>+NIA#QRa
5c+47Ra(<d=BfM.YXR68g&&C6[]#ZLO#JdG\OCaBeE&[Jd-7:8OXHP1H6+7cQ<(?
;5U,LL+gS1)7V]?e=++]HK3K<Q/?;E7)XVLCgY,AeZ=fOfdC_.WXRbM<\W,ZGVFd
ggU&Kf=7NCF=(\6PN7>#ZK&9g]aTEYTF[Y=G/E:Xgcd_.,Ld>@)MJI\dgZa#DRb1
?E;OF]AdGf7a7([GCV+-6_WEYST_H)/Wc5E3ZKSBU_<@DL7C35Fd#9a2;YJN[F--
YPb3+M.;&f8AP11E?b0#bWfZQ/707)[8I(JGC^:a+=A\A;+U]DU#88fJUc7]@8&F
9CT@QMg;c,(1a,0(UF+55?>_)TgTPBEU/EL487EQ5B9&8\fT&Yd;d_+a]1gX;AbT
_f9W&\Q5E/9.J?N+;0C=^b\f7c-B?\[_);/OM)d7<YD(+2Z3A#3F<?^EE/J&d2+Q
X0baV9)dZO);?H8KdC&M;OMaAY]=1>=82Gb7VcR=2\DB#fAL?1fN@R-T;T9/F6WO
<D65<[[D\<-\>]8X&M&6^P05dG4??MCM[.Va<.GN47L<FT6\_/V<\LN^=aYT>)He
P?7TL<Q:YOQ-/P2-M]_B7)2)R?EMBYeD_Q\L?3JM:IL,-/O2b3^J([gG7QYW3f27
g_^ZgS]Ce9N_OfX?1A=)-DN##aGJe7CO.VMK,;4T@+KcIfXJ]D@M;D_80&0B9U33
W24WDVU(\Y.MBQR_[2,8[)fZHP)[>ZCb2?V5/#>@#08d>&/EMD+6WL9@,f;9BW61
@&Q^]M\/aIdD+_3Y1VREeVDaaNN<P&ZO^UUC4O1cQ8.7_fW)XdG=?4ZTFP^a/1KL
=_3,S/D3\FA4Va;-6FAX0@JBJcXKT8/9\[](BNAF2E#7gP=N)/=_88eKQ6\ccg@Z
[:7FR986+d)\0KffY:Wc;UA\RAeQZD4-KD=a=W=0IXg2++:a5eNB_GX=DQH4aaW_
WY?8E(YALB\(3<@SZ.8fFL^A?JG+PGUG/2bR5NX]&>JEdTc1VG>C&(GBfK#,5<[I
;>fXVCf34<d=\-(6N)R?@C(;e;\gLP,0Z,5WaaI2:;c7,CY>@2(DIg](:L81a0QP
-7<,,4gB,L:[(2:;5R0:Re:gb4IVLbF#H[=CUVLMT&>UK911M26,83?@3?V58g1B
P=^WVJYQ[H,)[.^CN1X:e#XH\_QJ<MMd4=cP.98F6\4@#T8O2eV>Q2#aJB[>N@\I
B/=9gVWbLaACVU:#K(7De,V@+Z+<6/FSS>&_WH&T8RF975\4+YZZ29bQe2<2>ZgZ
/c/YK<;B3LUK;@;O?&=-^^8f9W,g<<f(e9CO5@@UZ5^;#b=7GI&_Q21#N@+IV;44
L03eF\UaSRV.X<<?(O[A4KIZ)-Ye2e+LecX@B+\?XIK^J4^WL7+Z/@\0G7B?0[_>
LOPM]E)(A[[=^#H1d03a-a..A4a6>,P:\9J)Ae0WMH^D,9@G19UPN4JN96)Pg91#
TP\L.#9L#I5->\5d,\e8/]:G-5ET)CgY\#OXN(:57Ga.@^NO+T[9R>+eN+(SJ)aX
eCDLJSZga:@D1WdE09_P5d?I(a5D/[Wgg-d^IW>ZK?E,+N;/cd9#=^47fS+?SNGC
4)eATB(X7[UTd(IQ0?7Zc4e+/b)&-0.M=5K++AK><0VPge+LHeK](9)V?6X80WQ^
dF[UO8Baf3I-C)<C4f]/\:X\9>bW(SNAH\^ERNY(2^K,;83(dP=KgeBL\2<F<EUH
=b(fAOJGTJG_OSOAE(bZ)E7A2<NJ>>/)>@)J/7;g#JI2J<=35e=NUREYef_Z4b&T
XMEVF^Z:I(Rf8?M[T.VV.W=AJBW64B(_;WZC&9R[P2[JL[=A6Af&J.e=O;g4>cIM
:]U>CCDEC.6(beRc5Uc-DSc:UOB&BNL\1;G4.6J5NK&V93=E/<RTE4C@d/gc0[O#
[3^EgA5R:fEa[c3dGY@:QJ4G9KS/6S_9@SJ\00f5\P]&W>(9H#FE+X\e0gN5<Vf[
5g002a6-d>5P\[T<\3V-O?gGL_+UUAH_O45#-U,XFfXT\\8XdCU,EeI;;=_HEc)K
@b9S2NGW_OJXZ=FB7UP_H.PVYc^64PRIXW)5/HB_5]R??_Qb.;VNATBc4Z..=HDc
9,[=^:_g=gMHK3c[[GRL6-9((AB]+F=XJ63GE3681TNGTRe/8@9dZB+Q.-HFe;]^
+IUGe3XgPX8[MeQZ&V=V9#K;5,VOfO]6aZH6c>F\+XW[=()1W\WI(-1<WNB>;HN.
6VH<&.0ESe@_2TBf[f]VLbU).CeFEC+0>[_Z_N#DL)H9d9S1GGV,]b^&eTG/AUD^
J1\DOW\&0:=g;=^eXN6ZVXWbQY?SUbX,G8QG62L4g<UAeW008M)9EBA1_-7)NVCD
O^G_U.+ERYe^PU5^/Ff#Igf#J>>UFbCPEG3IQ+4?Y]K6TbC]@?]:Oe9)8ZS[7(R9
+cKcS<GEW48(HZK-]G2VL290@Y-Hb9?(O<eb.741c]3NX=YY=f>K55CW7MgIXWK;
(/ZM6e6G^^fPMb\]MTQWV7IT9QKN77cT[:W&9[_-C9VX6.RI:dY?=+IM#C1;<4+\
UNPUL9de=/SLNRSQ+^dY2PA5;.D&Gf26ZRAT0H1LQ?+Z14aA[)[65P&ID^@K[P]7
&,F]7+#-Zb:_F-;-N[bAVb2M&C\@2E,;N1gTCJBJ4#VCP)_^?6^H2@>BbaIN=5>4
L1(DZB<K_a9)64EH]S?JS/)VX6L@&)a]NV@B?7YW71K^:3&J5Qc966T\35YQ1;+U
bZ/8KM<4MMX/0fbf2])_UKJ=]1M+;Yc;3TI]=5@#F42&GPQ:ZfPI1>N(FWKFOL80
W/X-&T41&.)(+HS>fAG1IK-)N.=@&LI39e9AZc?3WX,VEgG(UHHC[Z3b55fA>97C
&I2P:1TT@=7LHV0W=Qf#dgV)6+K,E/5#6Be)3QF0EO+L6dV^)K#c^K6?Se>.MYFL
+56PW29[#Z/1E^e<\___@2Vg=8^[CbKaVL98CLZ3QHMaRW47T3&B8e^XE/dg)@))
2GYX4S),ab_aHJZ(3facGf(N&XXKO#c9X890XF-XUS1fRJM)MaREAF&aXGKYAZ#?
4ZE]dg^CAC);4;AMZJGI4VL]+9?,K6A#@?@>OBB-Z=R.]f)&AM[=\4+C1+8C];a:
Q8Y^65J-fP@L/=]Y5RQ3=^Qa0;-_>H^]PUY2&J5SJV8T_LEQKM(K\@g=cS).B0/3
)1Ba8)L:RE>OSHT\@:3NK-/N[eJSd01O.Z0/O_ScLBdOS+\4c77>(_@AA[LS0RV#
HA#4<KUd;YDJe=;U>57E?.<:M3fI9>E4@B8DMK:LP#SDHT7[^#(BC.TU8RUZJ2BS
bP/13G[4MB[cg-ONG:VcNLd];Hf\UGL[:eKQ(B32U\+Q+\=0?GfB.3:7?;:G0-\I
c1#OJR=HDeb3L;cT<V,KIEY+MW-]LBb3)-P\B=>Q>@P..b4T6N[>=H8YYCSaOSSA
IICGYB;g6@\.-Y4a-[C23Y_A-+ELc31G;X^Y55T(fV>18:;^>)L^\;@>>^_1gY[U
cEeC@g1UCd;/]RTEdVd]CS)5eL;D3#1LCD&]KVdR]7JdUU,)#7He_#=0f]66Oe:M
cM3&-:#[9=E5L@[_I?HN?W6+TJ/H++>HG06_5V5G4.Z^+&20K7,II(5WWN9f6/MS
J,7]c/d?MTF>R2W8YZfU_T_:^gQ5SI]XS85,;;Yg&W4:<GVBM:ZMSPX1K#G=.E\V
IKL6?1X0-1]c8M8Z#IAZZ[S,NL^CYLN#EeY9XC^XXUF?\?/&;?8Scf(2UcG:[R#.
g/@F3R;fDS_(8CIMc[/:g=2E]]f6dEY<aI0T5D\@d=2Q;Ndaac__CTI7SLHXZ0<0
#&4ZB=3^F]D4)P9M4AdSeI7A1^AC]=e73[;+&/6P1F9b>SB#PWV.ZgbV,.DE;e_6
<4&<)UHdX/?,3_JKeT7c]NJA/=S-?#2FM#P^()_/.dZL8,\Z2+Vg1>MF)SQU<P]J
f4F5d-C>C&1CXYGU06-J\9LcXG^_7#K33@O=J.8^IQ_DT1LVb2>G9WN.7=2A90c2
DV(PRSH/@HD@K;<b913(@KgTYRL,#^<3B_a3O8.<.P58QQHR=521KN<&#)eS6;3B
Q#[+aY2+Q4VMMfc=+\,CG#c0-JIET79^A==S55.65b(UX(\2d<>8O6X]L[\F_@DT
9A76C?4F3X[CTC<)<Nb^da@[7+<3D.P2b8]K^=a+00aYJA-1Q0f(MEF&/AYWcMOL
gR43+X(.fgV+@OJQ@Y@>S&\d&L=)^?&M:_.N-6^cD\V]IRSW+AT\X1/?0TY,&XO2
DbK/>\?L>GV64Va=cB;;JKR7eMIH5F5H/cP9>>e+M9,ZO-aK+(ZX2a+W,NR>Z5//
DIO+;KGF=#0dZ,;Cg/\PXHL]3U,R\Z.DcYVTDW+L+5@938a#;Dgf8Y5H722E[8F8
)&DcA.cHGI)T9VCW8AafC@<;fL02SCMgT:>fe4U[B9;#D(6#KUMPSH,3IVgXP731
-32<a(7eM7+?O0d6V6PgH?F3@e)9SKWBHJ4a69/UP)J-3fR]C+VV[83D43@XM3H;
Te1BNK3H9_URO\-LT;[>Z9;QW1MCV;9ZG;RF?6_gU&?3@N9AE<@IM[9da=I+115P
eF8@HNe):,ZXNRR_[e0Z1S8]UQLH^#;VQ&3ENQ12T?8HYd)P=3b8)>aJO?PT79gX
J_gd@C#d([E,[f5]V-PE&/;<]5/8.XB9VKd)a?beD+/H(ARNIPTUF0FWgXTB,Aac
\[3LA5_)f#R92=W<K9J9K<cIa42+@X?)M=#>@YGCd.GPTY.aEeQ+da22?)GA:I6A
#B+DZQ:7#@Z/5A7S0KbdB9cO;H:+d&/^OBRIdPC>:)++(]?:1RUR&:b_\]FeSPY,
d]&.JO9)&?/MD(Wd@LJUSUWI,S[@NQ+HDY;A55MB1DR^UgG(_(B_N_(TS]:7PZ[U
;)@cWOVK+g&dbf8B5[I)9<]4M_+^Q54P-(1df.TYEda)aQe@]?&:;>/)N]OY<DZ/
U1KTX]TCJHN#3@B/&AN113J>&/_A]3Z[;5-T9A5d:D:,BEPX??E>\BTZO;M3L\V<
+]N8RVfeVMSM=78\&Y/]@H6EXYbfOOLJRR<3J=L)O.CCU7HZP];gNeY,Z4>7L;87
10[K+ICY]B5]G+/WF8]V(eQ@2-+(@,,1S<4<6:e0UA=UcAeNFgEMX=-;^P38)=R_
VZ[&)2;N@P/OBBNbP]JXP=K9@;S5d\J=;b,\;O+.TSW&8DA;7Z+K.#aQ/?FS,QO\
9?U(5.#e09@M8IF1DO1^2HF<[EgN7R:cZS\E2DXH()K\KI8,afI:DPfQ&]63PYT&
@E7YU0]OZ1F0<LIHM?GXDXNC2[EEO72^FYYT6TTQ@94?a5eX+3YS^0TMU&&T3])3
M.-A[4,CN+P?c@@9<NYC4-F0;^U\8@P[bb71GK^60dO6^JX.Q_.LX[MYP0ULKW1:
e)>-_g#Yc+@N0Gg3,;,Rb-(,<Cg=KE,?>>7=LLP66#+1,CS979b60GXR/a.G/;L\
7KQBdEZ-)11a3B:Ba6U;JDK?9NRd-JZ]K<WC6#bN_9)Z\QB]T&c@4d=AVFf3M@O6
[Z5F.@g8F)IST=P7EUfKJ<-KCKU_PMe4&/baD\7fEe9:=_f=O9YQ?OfYdJ@O+M]4
O^TIaB#U#7VDIA5I\R+cd6D>S37J6/MLA6\#U(Ne3a8(25NSIF9IJW9Y/]DO0d6/
geS4+(JTcf7>06C+[5S0M:C;J#Y_E+\VYb2F944RG)WXADe[HfO1,X2bI_>N-4fG
3+<cBO=@VA\)A]ECI:R]_Z(OOKS6V<3TH3f6L;7P+-KSS623>H.\5,HPIgJMKY@\
;FX41)5I#?Hb6@7S.ODKZX5FI9Tf-[W3.^8=>3TNE)4=N5^MM:)42=d@a5@=@4cU
gKJD=+B9Y)_0&XS#HE9g4,^_\B1U=a&?ZB:@3_&ZB@F0L.;fR?0C_MZ[8:1[WXe<
]\.&1#87\AB3/\)=C]Hg#fCP@ed\\YY0+gO]U=dJ3^F#bQDVO[_d=geF1RAWM>c?
+eS]K^A-CcFYb0f#NFRVeY&QE60(98\J+a-(.D+2K.Q+WH1Z>KP;79W1fV.[Q1e&
b[;DGH=#W2D_NbT^M_8I.^&[78Zc1fK.VUcg<eM4VK2]T5(gfd(_-0\8FFH8[V9P
ZY;7e;[[+0G;6,d^?<3EO8;@^(G:JMF\S/S+CPBdb@429Vd4bUNS;+aJd+9BCP:W
feP,H?f(OD@gU?@JM4,1O7?WRC[1D109-\W2H)?6Ge\TRa+5J=I8>E#],=I^_L(d
cVSS>0J@c@3=&9>JfB\b>(WZV4&cX,.ZM,[a]e#YgbaJAB=gTQQEe8UI5L6W^I42
Y(A8gg/\CbEc&H=G/3R+fc.6YB\+]?_1NN8dAD?^?2=H4Rc.A3e9+LWSVV\c1E_I
aP.>9Q)3_VRXJd628#5@)e6a1.a9<GQgZgGA2e5D2VNfC2UHCM>#AY3OUZMHXb]]
,#D-QR1bOW:7_S4VU9MQRfF<Eg\<5OHKGZ<MYESWN>=45Ef/@bGQ/=GB>)cKbcQ8
gI@8,B;c@ZeZDa;T-E_/V-4:46[4VC##g18^^Ce^Z/8+3W)TJ.RcZ__9A5:]4_]R
UH.W;_M9c?_c>=26g=V]\@4)I-Le\9dfI1KM3R)G[#4R?1MN)5VAO.)Y47Y(3N\g
U-/SaJ_d5UZZM2N>KgRFT0A3(Gg5BBW\WH5bG/TEQ-C+G;-0\b[3cdSH)XO7e_a-
9?b[KS_+008<9A]#^fWX6G?F>-V-[EdAQcP;;TS1J:LJ3T7A>5Ed:@?(NA10QFF@
:_Q9EPWWKeb?HLJKeGOeE8AcN=P@PJ#2@eQ@)PfMFG:IFN3?<-Fe9QObd_dW_D\d
CMX23;P-;YPQgV?:77GdW-HVeWa:96N-F4Mga5L^Z+T/G@e21d2G0bSDbHCd#\OI
=1Y#]Y77V1-8W>\XL0(PK-;F6<D?4Q</_&OI)?1b5<H4IYY@1)5C#dX,)#e^>F)3
M@2K1^2S(dZ]9S2M8fV^[]?[:H=fWf<=B;Bb:HTG0V/d]>QNc@Z.CK-5U:PKMJZ4
HJBb9&79#)[_(SZC>7RFDR&B;d(W>8FDGTUQ-.PT-bPRI]54_0HS&Q:;XR<+X8,)
74OMV=&VJZ7b+#\+fZ>Tc.4H8DQ-&d>/OeFTT0e@4>TRWed[LR(\,099B]RcF:5O
[=fSM_/dKH5W<Ye>0Ig15ZG&/U7][)ECfI;GV#(+J8]=Vbb?:AdbKg5@C?fBE8a0
#)Q?[K0.([=\g;9ER0ADRC/VeA]11I<TBb;;G^P,3NFZ:9OPKM)-5gE]>+1UE_R4
+X2P1?\@B#S)BS-a(ZNcR,5FaZ.D#:.?,AE>(=[FQd@+d]^9UF-LBD+cAUfg3B^D
<4E5D4I#0PCH5.S:d24>_4D@-cMRa.<34RGXgJ^-)0?@F?1T\\9GX,O,fQBJ/H</
J1b9:&&0gbSOF_4&77_]a>Q>F73+1XQCZ6XZWM3REF&Q3M24-&[US<?c\D4.96OO
Z;_:@O:H7VMHC9;KR1dPR5^G4N4J=26#fS2_;>8_DRBIF?Qe=0Z#NZJa.(WHF4MT
704,4Jc9]eW)B#=E08g7.U=I@W:L3\,G>O_)fLBHR^1U=YPWP6O?CGKOH&d@]=6_
]CLeMRQO#-beb)O=F[8c6Ab[PV;,SW_;2ERCZH-HTb]6M(OYaZP-T^4gWH4XCKgN
JO@N):0WFHa>g1LB0><UU:S9A=UNNQ<S]J(f:FN\H;Bb-U7ARU(??=.W/MeKdG0V
9g30De320D/8Zf^&aZTf_YHaFLMa6#(8;[KB0&Z91LJa#aNXcK;\-1fd])W+\,UC
P\J6^UW-d1Ja)^,UeRdIS[^e2aHKQ++U0gVD0_3)gAKOD0H)GW3I:V[E<22YNd)9
g;f5-YQP.NN6R^F;2e2.=+_)6#MZ\I0P-,]2ZD@7GMLNLg)7c\5BKNYM[?WOZe\H
d(CAHA6g-46]JF=Ga-SdN_R&D59g/-6,60gcb85K659F48a5[7bZ8UTeMCMFR1[1
K;QLEUU.A]>a+;8>L=XeJROgK:gJ=4Y.7-;,[WKf(ZBN8@@\L5+P7D;UVET+JFTA
=5[Ng]HW9Jc:,R.cXMN46P2)&_\J>FJIL5NV0XDMLX.fKg3+.^W4,^6J>3C5(cK3
9E9<L5E(&WXHgZVXQ),ZLSRBQ41Q[-=.gM+3B0&;OV8;J\_0e2f6OFQV^IC\L460
SUA5QJBG)>\U2]_e8#F\OUO_R6f?gEL-NabV/R+;HSSZ;HbX)Y5:K\I.51G.4I9^
I6B?V4>J:>8;cQ[dJ@J^XE#\e&@CfHTIe/LKNGd./ad.\4RW=KL>g^cAT09Rcc6Q
UW:Z]O56V#R>[g)-aY\T7PFE^+\9L6+Z8IY5T;OFJ@;TIOB(0G\NJR2gfFPH)6XP
IFIVZILYR)ZJ[#;>[=2F@QE3XK6I[J;2[<#,3dA>P^Zc+S+e1U.:^.[-SZY@a,\V
,>5</Ud[<#&:[.?ZHRW1fZYLgBN+gU+A>WS#DDI;S5PL+Fb,c,9c(YW_-PV1#&(3
:3TM)fVGTaV^^f7]0^b5fWWbGeW;Y[(9FSUF/a#XC9?&<ZBM1HaSU&OI>M)b+L)D
TT[:+HS&1^OGV8,LU4M5/TOP)G,1[,FMC.BO>/g7a_EU8H&JDY&8A@a9fV5P(b^Y
>Ig1+XWDCUg.YV)IWMSgJIcW(M<@6_8DbKe^0NKM4g0gbPQcFOW9g^Y57aaE_G[b
Kc63UQBEfJGDZ^+&.Q?]]g=FZYL=A?>0]2/:I)<JKI.0DcE94GY@UCP-:6=6.SL7
3M9=G05H0FWH&8K5</MR;,+7^Q@(aL3F+TGDO(b]&>c?A<4MAga[dIfYBLd:eX(F
(0@0[O),bZfX([^NMN;0gdfZ?H]QXHAZH<).@TeV^7/VFN6Q1CTHc02I69D>JDC&
MO);@3+182>(I-e+VF,HD[9gb\0eQP21-#KRAO2VN6+UI2QaMA9BCD?.b2.eU;0[
U@E^=5TBg-P].\e<^=I=/R?SK=eDa7f7#5,8+06&O:3=(LWbKXTIXHIX3&a9NW,d
5.]9C0Wf[Q<0#5GcSYFGW=5)G_<PRC6+XIX9#Q.^S3T([UKH=_2;T@L[@eYBUD-J
f^MIEQ[&LNLbGdZ(8@3K1Og,WY;dFe2/9>]WDURV)D@;Qg:MdGUV\>T03Za^5<NQ
ILbJXK:83U#^SD_&:F]]RJ1DI(64Y@g#?ET=+eH.>@:K/@2b1\;I?&HTJ5?\4fRa
e2.;1I\,K1W5)S+4M2HQ;OS\5fT:L;Oc0^?f&9_N,_;\99XC//]#WXFJE[<N<G^&
?4064EW.+#HR&,)d)>@Y_1+G.W[9Fd1U=(LM^S6[?543&FBSK7U@]6(AV11_(X]2
)#f5Z73)[5<BJNJ7V.a^f.E7<+/FIH[;dS?=SGb-bUVU>]]3cbdZ.UcKJP.@-&^>
bRVF\B&G==\_L179(T(QKXfSZ<&&8dG=S]/bDD@b21]=E.DC>EfGM]<X/3-^O^01
)I_9QFK@)P+-\F)>0<-ZJ7g0)X&&=B=E=U.Ud@/=W](]&LE/d@c:ID&()=M_+dG#
2Q3<a++3(^I-bFe(S7;e)Z\L0+0[7@UC.G.JeZ/K4<]D1KK<?2HHY(/3F)14C0)H
(b)T0YK4?Y[a#;EZVJ??B&-7<GBV]<L9Oc21-#5;+Xfg&V.=dU_Be5VS.]CO-<4Z
g(RJ(cbXNJ.E9ILbO=B_[;:+M/S)1.a@Ce/^K0)-[Y@c1-/7JO1HNCR(_K/7PMFg
.[FFO)^X^W2ObKI62d2=eUdT>3&)8dW+^G4/-Ke8X[aX@[BQ#0;OU70VW4F=X<3d
[M0+b_H@^=b&S27FaUOF2?(O3E#E.&BD_ZJ<]SAMLc>]7PFJEU[^,Decg>\e[DEH
WGJd2f[C:bIJQ&A:46e&397D_L,aO25TdAVAdCMS[8-,R7^L4C1N+fKC68SZ.GI@
56JX@XC6,WHD_5,RZ4@f,BS/S2;OQEaBU<ZA(_cH66N+:5HBbA4?G.J.:<A@KM1<
\Sge;#03;K&4fG@(Y:-H,5=FD(>C\K.TX]baW6YHCO?/FKPM<Q(^[X(7NdIVG<AU
>Y07KCbE[K.BIQBPTTE>GGg3EH8R9>AXKIg8(3:Fd>KJ8eJ]L/<^.I9V0([WO3F7
L?9RaDWSKaV1WE?L?R2^ZT6M6_WG1BW^fLTX0ZPdB4/=4#;?dO@N\__#BEAWPYNg
&#E>A5XIL1B_6.G5b8_>c(O>3bV-BP=/\NY+T>.&cK)25C[/ZIRC1H(IRTeKg@QM
^aXD7TRBZA9CDK@48U(G.CT]e1Ka;/,88YY,R<c/(b9OJ&6-9P8eN,L3W>09V_WR
bM0e9137&f-EJHZCL@@J:dFI/.<]&X(HH_XMM38BgXDRR2=I=_41XCBFY4ZU;+JJ
/c_4DOMg4)#<Tc3ZO=:,IcRH^/K.JS?QPP=9d6PgY+=egOKdM3+1CaTO<5]@4c)0
55)@eY1aU8+G/d55c3REUTdK+,.2J;7dKCf?T8ZYW<c]0LL@E.C=V@S<<JSBacO2
)O[RYUbN55\>Q0NG0NX-PT_9&MYdNA_&GdfND6dINA-RHKDH34fP?8D5PI;bEML1
@4>[E5-R]-G18<K#E4C1)PMJC76),0WQ4HTU#PB78TfIZ^H^D^\BgU0D69(RI<Dg
)=U@Zf]>E-99gEX@aZ;6N=_XXUdIK[UabX#e@=#>ACJ?dH=C^G<F/JB5G0gcff(,
Q<6:f5N:T(S[X7&;DVGWM.KVFSCC&Df.e<;B/fJ;H>23(I-37L::Q5:WIg-bbP(:
(LV>&;J)E9;0\=)XMHWOf6D@[J:C\,86?<R&Q4gL8MI-F:\2?:38]8^V#W=2?+Y&
A]<X>0X..M>K9>d@2)H(X&HI_cZBI][:?&6fQT(;Fbb^4aAU[5V.J<A/g&bK19FX
2@1HV/g/?KRb0.=29GH&2-\Y5PBE=N71=ZfP^F7RL1]g&3+WScCb=ZAcM)=[9/1]
\W;9;_/L&7CLg8RUe9H/9SFF=0YfeY1O?AM01GH^?,(Y\)5f\^A#V]E+-TfN7Zef
\3CL\TJbJIH3)L_3cN_;Cd6[&_a(9EH#d=.ZW1IL=O8bSH,]/A(,GNIe73UT4g[f
1^L(:gcZ6Z,7LfDO;&f(.)P?#+(<daIX=S;252:e:DeJJ[dPd^=f4)[7RRTOT8SY
U-,,NACW3:6BQ//6I3YV\ggZR)c=PdHB(D,__G)ARF-Jb776,F;>]-=0P_:>6Q:4
Y8O.dE+BLU+D#VJ2gG_SS.5&WX1(=2_c&N.Gee6E;8<OH9bVGf(EDWaX.:[X^D^+
)I1_.(gQ#-0+B+4Yf=Y#6?8g91TP[7c,KGY8UCFd0YeQ2K&U8_EcdM@cM:[4Q)-U
Z956@2H3K_?7[8T:OUC1H5-;APA,A(1FPA:H]JJ6a_g/(BEAa=9T5/aP-A@20.2:
f/_@Z)OE2MAeYK7ORVOAXb&U10/=Y/PNbWLX(Rg4@O<Y<MQUY)UKSbNVee&5eOAV
Tg;6He)@cY/[YI(0.9a1O&g5UFK7cDJ;2XUSNG?.e3;4=(J;bH1SHAY]).GW_aR1
aB4bN.KYI&K.5@_5U_@9B49V;-=(,,?J,RL&b;K_e:ea10;d>b\@PZDf>P[RHU]+
F^LgG/.[93c;U&,g1LHPAL,LX^J.eW2L#RR+c1Ic8g.NHN0#SU4e;WU^1P.>F-C+
)8gUf]?[V29-UG0,d,)QeDT((#]J#:9,\Tcd4NZ.<;\KN6>4Q,,61NAI95[3J3H+
D7ePN-7SPF=>24caV5@JG)dWI/4FW3\6M69>:?=+84G1c=]Sba_8K\:NW#YPeKC(
LW,)60?FT@3^-2L=#)PV?Bc_<;4])AMS#KU:U2;e_6?,JW;OR\PF14\A5)AeEZ5f
Nc[N0YHAEEJ;\,H[c(cfZN7X-AAeF&:T\CQO),YFe:2Jbc))=:K]OL?>6Xa0e@LL
8?4R&afK+6-@ES8;PQ=dPMLaf]Z7<4dA6FG[?EB\G+M<&6&=DZLCc)JVWV,>FafF
3:6Y3<+LCVVF8(A#H]3H\MXVMGY55?PU&bU74-c-D(W5;Z=ZRA;WNO+QS_dFNLM>
X^G<1GcS7B.G4QI2O=Z6[]0-C]FY+FAdS5-G9Lc7UAT_/AOSBRO/;G(UY^X/Y7aS
\6Lf19AT]7c>;U)4P(H&eC5\<[_b,78RM<EFMe/;f.(IF72I9a3U7L_&/UAR=I&E
e0O5Zf^<=MYb_+D[E94&J\)bSRd7,^Og]M-GbWU11aNA/f5Z6@T?7)d0SVDEfJ0N
W:]QXE-^7bY2?LRKf6ZGENH4R_R.fE[2LbJR^XLX4)_.e:Da#SQN.MZ49Ee\V3F&
ecI@cW>O/#;K:A@a-35dHQ<O[T#Vc(aQd,Q^VB6H(I8Pe6#+b9NGDNMSQ=U6&E;.
Z5@T^UgcWg,I^]ZZ4CSZNGfaS=YTNBST6R-JaGI4FLT_&K/C+VZcXPDQVa(.Zde>
+<Q4\TXf-PNC^^gAOA8eQ1]4Z]NDSb8HW][R8a#0H<L:&g70bf<7,#,UJ3#X<SV9
B^;ASGODH;B(1N<Kg^Y+VX5=VW]9(>DH9Oe)MO\Y#JNK43bDHA-[HJ1O6G<-S?FH
^E)350XPdOafgSDCX:HYD.7IRI].LHaQU3Q:3-UP4:DdQH(9W,(>,)H1TDI;FVRP
).9H-IV&I&]T6)\,</S8:XH;FcFO[561,cTa7aKM5\HL7;ZL]_,K5fVaJY]?+.;?
be#R,S(Y+]3O/Z2]JU7C>3WGIKa:cOAbfDg,TH05Tg>TJ(Q5e8S88FfLIfB>2&DC
5J^?e<2>U:<X4&6Y;2H-_S>M]]Y0TU2e9,HXD5C:,^72HRRIND&eDFEH/f4>.[-5
L7SL1Q6VgDEc^TP9d]M+=#6I:CRDI?-)@4d0KEeVcG0)D6-O><P[g;ZS-1f)9Z[Y
_D^9cD-4UXWN#52?>.)@.#TEbQOZ^Fd(4M&TVH(3.VH[V+(G1907V75_GP\CgV/(
eTB0EDg_GHG.PZ\S=90J@U7EbLK4gd\fgK>[FE\7MYZUX\c;GPWEPQ\HYVEY6/4U
-+GaVDP/b+b5OQfH.55LggcdUYI?O/Q7^\#g6g?+NAD0(\(8Lf4^g/e^,[dfF>^d
+Ca83/))=G_-2c:=/Ug<)2C>[_N:JGUbeB:1g71?C9\4gM88)G(,&=DBe6G&^?/@
LXQ9?<O7>UE65:#GP4dKRG;=;^6B[9D=HEb=N-S4><[A_@<KCgebcE[VK&CKGO@L
<V.L>d5^3P9fGU4J?^Z#5>7._Q5&9F#93EZd=YWM,FVb_Z(#Od::f:38^_U&Fd=?
B2QAb^OS>#eS/.9SA8eN_[b,:&SEF8^d\@I?M?XQN3XL.>:V6__LcG_eVZGG+]MX
JcAfA8SZ^EE)CUf\MXBUcK2:>GJF90[[95[XQU/X5\;[R)fL88I[gfP5,_@gA^BF
[CfUT5]E3eLR6TM59baC\.T<UQNV6F?0Ga0D4+W3,B7K;<NfI9<IJ>U0dP]0XA;X
<+A,.650KZ?@G^BBA8Z1ONK3_P;<KX/_C7<#?_+G232W(U6/L9;1:PBP_=;MRN24
_@adeA6H7bB<fbY\<2d^+TH^[LfS#T1+:^(A?dJSf28>?0FYUeFA[5M#DC8MC_>f
cX&_aR:B^KXI#7/TQdB?.Z.CBTW:Aa(=RAIE\JTXQMJ6^FbN&UHeOSRf4N)bQU,/
+2.(<3ZZN.Q=5OS-7A?.OWTBeX^FfSTW;8AT:HbIX2]]/Z-dXSYR]da2]V4Aec4e
I)B-;K]Q8I1cGZf_1SZ8YJFSf<L2AJ^H)]7Za,E?Zb>-/^^KWIc&7cH;1ENC8Uaa
>CA#I]d:0,/+Z??OSK.))#)TX(8P\B-QdY]&TGLJ6AT3R8g?8;\<U1SZ&@+)HFHK
7@S_C:(gacXW105@-QE7(C.VUD]-N8bKWZ:=FD>97-6-FGS6,E57HATVJAfS5L,5
=[;MIYc>)W_BYUI5?X,BO/S.0J\13LN^1RN/4HVA4>+=Q>(RI)=aW\f2O\O9J65^
6-FfY-B[_f/[-KJ)N7caeRa-;R]<KJ(5U](JLeDTSb6M51)7\X,=Xc/#?LP;-S^?
=KS/.DH=b1KgEY7W+3Y=.;c]<V8K5/>YD\RW2/?4NDAT+dRP-P,YaC30G<-Q];2S
_:K?&)GXd5J@B/R;2-.+1XafTJZH]#AN[f?-_c\/A&F[V^>Rc(CR3,Q==;,\[DbP
8V1GV;98IfX/&PK7CM0=^OZgJYY0_6QX>aT&<WLPGPZPBb[d&O=,LET:V5GY/>40
[0^E)g(=6;R)K9GA:gS_a7T3U4Q.E:31R1@9f=LPb[Vda-Rg5Q8U&>J1+YWa[(J?
-)CgOK-5\=\WE/e/Y@IMH+6dQ9#bM);Ofe]J4CLSL3\3dPX9Zd>QWR#^>_602_3>
Q]@:G-NXB#6+O_Q7c=T)A(Yea6a#[TN5+YO.(<@=N+)L+4K&dQ?&X7U[:>P5Mf9E
gFDJ)0;M9[Y;a;6L9@O:9fXM(81@\^OPCE5cL&#A<[U.06I6_S.NILFP^\EK#>\?
70]R8daL+]T3JDP4.C;(VZ-7P5J<&@:egBZIPZcE3@8]Oc0I9P?d)T[)cDID0X&e
)#T^2W0>786.?46+9=9:KZ^R#>CM^F0P&LQ,#b/;gAbVE_U.[ZPG+8/,Cb]<9-fg
QE/@4GTe5Qb4f]LXcGc:T[56I9VC(;[2_1^-Y_0\50Ld2;8(COYE,f_?IR7_V-6F
]@#E6:gd8K5ROCbEUGa=Ca>K\e76aKDKH1M_S3/UaZ@<RV3+/E766;F?\Db/@X24
gJ=+[;/-CVb<46(<H,TOU+#b-aa4CCcSb9D;c\OXR-#>H\IK8Z,CNYgB[0(.1BWG
Q^?E9T:-S\2GG<V6#9JW^:g++XbVc/cR(Z5Y?-SUU#Fe0JYMX-0[HdPUL[Y#&GM^
?LaYBNHS9GdF1G6OR9eadM=-5;3\I^088bS/VbP(c&(/J:4c]_cM(RNEBJ88(=-V
aB5/W+GU,_M<S#FA_HOa;dRcCA)^R8(/g]6>^4L#fdLd:aL<DYf5M9_W:K3U7-bV
OWSEVK3F/S#E\G7]Ed]3K3[=b\W@a>bQAJ=_P[d]VK1ZL\((+-gQG&[H1cccMZ<9
VOE1NVPa[W2<Z,(1Aa13eF3KPCE_T97K.d+/ZKIY>92FXU^A:0R_b1_36U=R520)
H]@HI>HdF;2Gb:g+.g1DEbG)+@PeHQQ+)dc50[\d/9.f972be8P,BS13f8^?V;(Y
WRA8T]MPL\NY34g3fY20gW8Rd@c^afa1],&bW<]O+dXP[I9SeDdJ:7IRdD2SXD@B
bHfF>e_1Ac_PGD\4U^KZOT8-YaD7@Zc0#c-J837_F^EGA?N[2+dZ^3]&7]3g5O(G
QE]RP6H@QE;06EJE.#<OK^fDIcK=GT?-a:SZ/>?L371A0d<1g)VA9dRc;XZNQ1NA
Y31eg-Ke(XQQd\&,^<f2UHA]F6aeZT2H+[5Y;(:RZ9.2a4H+K\b+5f=I@@^WF.<6
W2Ib?&&5e\]GMC<B(K/KMLNB7Q;OMP;;gN-=F8a=5,^6X\]E=:gc-6B[[>bAT?DV
DC[9fTY[^WT0QC=8B/&8BM07:1KgGA6_\[0E&a\JWPK,:V#_#7<T,X;;,W-XGd+:
&@V/4Q\8QC:J@-S1AbOMf_.S+Pc.=CC1>QdGO2N,UL:#0,+Ve6Q[H^Ob;.:R9(_G
\G1@gTG+C+3@G2&9VGN+-Cac7=7]#Ye3AGGg,E,\^45<gW+;6,R\_Q^UND?f)HGQ
P=W-Jb24;HF:SMWR6/Z#(U+17ReAJX^e^>F2WQ6F7;KSQ0<\GNRXT8)7T4T>dW\D
c[B&L;c@MCb(@]CTFf.6OIaY-Kb@^XHMKXL[U^EF2NOO<VBZZ2D9c][H^JNJ?:86
+IK:Z:=G1.#J^AQZ7^0BS0NN)85PY>gf^F_ELaaF\RAg^QbMd_3Yf7)7NC2FN_A/
AY<OTNU5?+MNK[E[V7W?gD>fc&aQ5-Z^(&2Z:-W<dV+/A\:](b^TW1RcaF_=BSC[
T\QE]Q3<<FUU#(G[6::P&CNT(D30OMSR1:-1<d3)AYcK,_I-<0a]g;MVC=X?\HEE
<=1WNG_c?97PC2[5/W#@A\fO\OgVM7::Q3.+4AF^EOd\KO,#a4-GM@FJ]Y:US&P7
3+bS7WCegN^>FgNDMULO6@W+>RCC?ae?D57_3W@CBNQbFPY^@Za=G=-S3,0Y^)HY
4g?RY8AOZZDcR\-]Kg-dD++=37S3FX:RJ0Rf-IdZfK4\H<8J66Ld89>gS3([+SW3
bG/V]Y)U,TU6>Md3WI=+?#4N1LMP#>L2JV>J1Z=.XA+F(g67D0^CG6571,.&/F76
LU801B?HdGK;#U@E6G364OUTL;VdTHfFLcW]gSO6A&-N/8+Q^U;RO7-[\(A@S@2+
UPO:+KD6Z3EYJ58I\CaJYaA9d0T=dZ[Z&9FDQcFXZ9K?4?8?b3MG/4Xe,5geS&La
R^,=cXBH>AGR@X\7Q_a+35\PDL^;6VT\T1J8F)VJ3JL&+PF9dTFe@_@Q#J[U3/74
8+^O?BNVe23&PG@R<C476(M&15acMUY&X1<5dOS]Md)(\)3/^FU.VVDX[#S3=>Ud
6TVYR[K./QWfYXJNIAaVII5VXaHH1#5bG9I91AG:IB,fOOI8fOEZ9-?UHbb)93Q9
UQU)H&O<7AB,D:BHC^8<Ma)7W@FIYU6=8_E/bOICQ\UE&H>7F[Q6Z9-Zb(g]c3E&
[C\Z+/fSV/9DWI:cGV6@Dc1/6Y,S-/^ZK]D5P_eZ0L(55UMDZ<9HL@6Y/K\b.=IZ
S+_;+f.TS)LQX:+R&B??6/4CNSN1FQF^V(-RV6bNRMUcRTZcZ+^<L?=>Q)[TV1Y#
I\#:;Q[[@_EWa&29L#eOg632(@BKfRJ_>cR=F38e,fV#6CI[CIe+CJ7;ZcCNW2D(
,;]N<IY@;If(L<__#]=B)RVYQFPgeQ:a/a?M<0=#G>6QQT0b(R&D8\6?9_gZ0;@=
3a+FK^>6RId6GSNbG#RZd?6;C8-;g;:;BMZ4^0;CO@01(FNM#S4Ae?H;E5a+d1=W
@>gK[LVT_A.<I].3:QCIe5R(.>2>SfYF?Z?VX?Re]T4<@]8R4&X?3G40>DBRD@[R
2T)[Ib0S^J_b4,?XI1AGV_;L_-;7?KKaZWE\5#WC#dIYKJYG6P?gPPE\GN7YQ2_D
M1H5@IL#Y^]/:#1)6Gf1X].?5>b8C_A3SES:_VL?UFR;MG@C,/2H+eE?A.)cY]4T
dNdDF<N=O;b;F_DYGQ5O+Ff_V6^;VAE(aE3C5C3YSRaYc);&EF<-X?DTV\UV7ec#
(&&?P0D<Y[+MN2fB#SJ<6N2C-6RfUVg6(1+GH]]XD1T:CS^@4YKdae14DN#91L4C
TQBgJ1B?\^(@:YaEGM\e=6g2:V)9[8Hc+F;7Pf1Zaf&T@g(\Z>9-,411\_&HKKG5
?a3H]RCNJ&DK+aP_M]g^E_MZB>de[#ZKGd8V2YEP:5F]=S=Gbf1?<.<(KNNH/OVe
N_Y)dW0]gVHVGA[eX?a)Id6eQ72d,YaCcWJS@3SDILW\@cU^O5/H1O4[9<bDDeQ7
aaY&,+<0_??Z1ZLc=O,WI(R1#6-5HWJ.TE0O#K@6;K>fdA>ZLgC[WH<(b]44=DJ;
H@D>KK?S)bbC8B4KT775dT[>+=7\bS=R=Zd61A.LY.f\WLVX4K\K:H:L4K&6YTX\
3[IS&G[9VA-OT;U.W:0O<Qa_5BW=WcbTGf12.8?[_TSV,XI:UOT0(?[/,WVM2?E=
);-A3=2\;BF&IG1>A[L/g&\=CP:MAN:9#WbWZc;HD8W+88.aD-fgJcHN\_R8]K2[
X,26.W6?U1?F0SIf/#7T1RUTR)aM^XeW&cR7<6;J(PZD_>/a<H(O54[EJWFJB0C_
9&fYF,O5dXWL1([3Ge48V1;.D[6c@aX3YD-]^CL/K_#59GT7/GUJAS-R/^35K(fI
U7Y.RHd.@+FPAKLdbO-fWR9F,N5ALKD8T\caA4F_MGR2H(/3.0;Zb[4+[L=He4U:
I(MJN8(34F=ACEG49]S5H@>><QeZ@Ie=SSJbc>1O+63EcgOOP?02^?IH3WA_gDbL
G.gf7DV]=+8)b(e.U5BWSbQ0FI[25C)EUH/G#<2#gFg8]_0U58[<7EUDKFG6cQ-f
)d<3W4Q[HJGbOU/1LKeX9G^-T>VT(gc&<f@;=1F25:KNJ;D40=W7J/;?K>5[.7C(
ObD/FSN9Z=dI]bU6gN&L4W.&K8TO91H@SPN]UWG<([g@aR2f-QAc(@Z]YM2Ed)Ma
SeT&4X=T6>&Q\LR(]JYSecISX-::;S:23=W&;N#UA7IX1:?PGW2U#-SZ=MY[Eg^e
_686\L-;fb-_R5#IL2a1<d@aD4:Hg80#J,A,TG.GbbfE8K<6Q]78@ZHULfHIF&AZ
bf[MY5D#\f@(#fUMV>(;\#J]^@]JY@2g35,7<8(SIeF0HPD&MJ?=P5d(N?f<\.P]
NNMD5D\#MaDK_SH)c&V9U:_2g3E_XN7.+RI@VagaFQgN,NBZe+U,2+[IegWb2X>W
34FL;TacOMOI@A;.>PGB5d[3783bTI],<G0&._W83f>I6]B:,RF.&YUM-R;X+SO/
.AA.XSf&cD\ePBb8AfAQ12R2;DA)(-2Q5^=3,]<Q/9R-NR>.#ec[dP48f46K>VPQ
IN<)CR0O],RU\eIP^)Z<?3CVQ:XUdZ?(+TN4.Vf#_fL:OQIbP3CUI1>:39YBAKUe
^V]]JMccXZ+UB9B@e?IUg<c@caH6RD5,_1J7[T2c^W)cH_L2E])/O0cHRgbT9[H]
4Zf(cM-^;0Td,.T=cB(;;dQH24OE5F<=9?\9=D-N6?G?C8J3:b@</SI7a>6-<K7M
OMKZ.NT/[7f<E2@2@@/Z?>gSUYW3^:]RP#B;H?9f1[HNJc3T<_P\()84JbYQ?.(4
20cR#3<4E_S^R0_PAI3f.9V5\b1#T1YKRZT??\:.2US&;e.HJ[6H#Dea9\OZO]95
AXV5PR5L@M.MeNQ0Zab/<=9BJND#KNea4d5NaL2@Y3TA5dF4:E<V6Q2NZU^FD)\H
><T;#eDH/6]@=Q07d7G=UWa&W[UG-XA+&06.Y1JbIN9CB/T78V9Ac9GK^\89[^;/
N4c951V810#_gIEQ@1#V5#1M>UTK?RF)[G2V.0SUH:=.N&AMTDX2;USbQUWG5YJc
HO:7_W@c[@L?agP)SJ5bJXCL5edFSM#J_#@YVC?LKb0aJV1N:&eT=fWW9<?.XQG[
OQ<KJ4#KbH5)7?<6]gX6d,[5#dV35_NU)bQKE6;@K5>C0716U39]BYR3(08TgN_I
cKXR^Y19-d0CX>3Y_.4J27@D@BS:SFCGX;/-;:P0C)C:fF[6^<&3g@Tf;GRQR_17
32<OEZ@U^dIg>WWBT:7e1a>HCJG9G&HO2E<g.A]B>bd2ZUgAG:dINGES/@=Y@f&]
/_+aWB#UXIC\]B33,/d39U+IPD#^d/UM@2A=)HJO<<J]fLRT[:38c(,]A#^_Ja:S
NgISg>a&]:fMF4&GR^K4E2PRNPZS^-[I;[d6b,Pdc/:AeaZ-\S+cH&K=->LaJ6M-
:GgbH6BV?@2A^?2-eT\)a.4g+3FEM]H\>[#C^#gBDFOGSQ.VO1.AY<ZgGJGH[db?
,O@aJba&MRNQ:[gFWHXCLgOSOPC;X#H5cbJEca1;]<BN,;1eTXHGF&=?KE6HDg6W
:bU]9/P6M_U+T,e(1cZ(T@?aSP0)eF1dP\g/V?)&<_(Z7[[(RXRTc=/=K5:]<:^M
;:^bHeBHU28\<YCgMbRW7d>&gKAcM]ReG<GHa8@M^2I#HWUT=fe\2[_T39R8R;,[
0N8WVR/&RG5X[SO>F73U1R]98eVVO>Y5fZgGCG.(ZUDb[X=,.S&[L3-fc37<Ve+d
+2Ed]fXK:g85Ce7HGU]LGH?5[J6=5e.::/&(VVH7E7[;P?PW[]DV4cXMf0FSgW_K
EUIGVXdF@7S_cJ1G&(Y>e])R5KE0G3L.:DKf<IE#?:?3G[a9.O8^L.[[C14X])Y[
(cA^^.fR#Y]Ua)U.ZX?.T>^E8#5_C#R5AJ?<bd8HXVa:_]W6ZU-UTFJISL:1..@C
A+IWY:eOFVM.BHUeV4+]OQW:ELd=HM4:?.-\)6+V^R8be@.\gGVb1U.RXECKOg0B
#T?0/:X65MCgbd5GZ,70Ag8b_Y-J;cF>;[N-.2=9Hf,6:V6Tf-KV^=;#Ng4V)+.@
8ecIUM#D6V_Q]_?8TaQPF-Q.KWZg@2DR(VdD6[N^]#bD\0fVc=96,O4P]S[>6B(-
PXTU;]#7b]0LB@&7I<E[fH[_#M5<Z^NW#[c929::cT+:d,<@^Q)B7N5QF2,J?#-\
K#WeT_3UTcC02,L?A(8aOg;:_69=+Z20cdNe);ROC2F/OR_N2V,aLdR>b<GC.L-L
g8F._;/@FD^HD(d<C/O(d2e-Rab]3L(OMYO[aHYRg(),g]#8TbU<a&.bNWDUK:>5
URV@F#e.Pdd=a(R.0\1(G\#?AY@YR1TDN/&I;?Oa75J)0\CX13/Q]4_#<,D:XIVR
[d#aKQfW<f21baW[^ce6ddfU:8WM-SPPU_R?4:+3?PGJQ5e]YdeY]a02MNPa?R5T
5W^+=dD3WDH+NMEJ-eNOBQ4OM?b&?OS53fgBJ]Z.&d-fS85^+UD,K:6W8,LW@G\+
PG\G4BL#cU,GaPBC6/ECg-\;JZNORU[<9#dVd)(&CW[-d0HA):L@KfI]aO0=Cg9H
)/W\Yc-:9BCO4O<KLU^/2<^fT8A4-Cc59]X<P(Ca4LRb-TTK;gR<bHSA\M\ZB61(
L[07)S3CJEQE90#aA>DP[Mb_;fYI;@W2ZD]>9/0EK1=Z?f>I/eAF8cVEN9TOIQWH
Z=P>^(Je&2\:(,7A.:cFRUcV=TNSHTTDgK:H/,5/W.[JP)0OK;U)#Z,F;bADI9J#
A=B\0Q[TO@=^IW,]3aRWT^P?VB0aY:WWD;X\e?4GcVeASZ17TK-Na_H1I::S+eS.
=?GG_c[]<;10V-TE#A(HE#_P1dbg-F_Fb,CD]b/9\&CEbNY]]-IddMZ[TU)bBG?^
WBNK<QJ0Hd^,8M3N>:W]JcPV)>CFQK2-#4=UA#\4X/\fJ48E,JN\EM8=(_9GeeKd
;[L3P-VZg<0-JF.=D2@Y=90_?I[JRW6T2.VR&<UMQ1_39E4_<RC6T9c<JgTS02EF
,D[_X/=?2R^G<DP;Gf_\[6dDce@K0B#<f0Z&H,/X&K[LDBW3WQE9OFI@)Tdd(G@=
K?]VaNT0,S15f]\5aAT\N5?7d4M1SN8\b@Q4UgVZ-Q<KOHAG@0GB8ZT>S-Y=[#aA
THBI)?TWC4SbCdF,BDBCP23S++[/gFYY9S:;;QORe4_HJc[c>#,W.I)SF,ZZdLO1
[C(0=4W2P&OV;g;8(]MP+I5SGP^(GM>F/4,]\S7WC7P8NXS\N(E3ZR5/E;+-9D39
5aJ1EC^LcFHSU-b+RB45.\E?Y83aMdW>7;F&PN72UBa@,8BYc=LbF2e<P[PaQ[KR
-4&;6U6TEF<0UWT7RW>DO2?dUS-_..8,CIZZ0>Ld^@Oec1bT;YUg\[83G-=+YNO6
^_D==?6RY^#5cZ8/bQ@DTKM):;(:>@f)0I02R&L-#0=1Q/M->c0>BUfd<:]169M1
[>JRd4HA\gg6=^C><R,-83WU_YW@DV3-RY7.+\<Y0L^&N)2cB]GfMBR\(d[bS/DU
YS/IG^)Y-TVX^/4?6D^g@+XPX]d)ZLKQSI9E(+4>JOBH(bS0gSXY(a]I#(BEC)U?
U0.F+;2[(NF^;-NbMP)_2L57S\0JT3b_4CJX_EFbR+bWP?6E+#I_&,4egMZBQJI:
W9gMa\YUS)bAVf]2_:N60-+)WL>(bUBa9NI,<D_<.N-)[<1eUOd].R;N>#M,HG8T
.M?dX_>cRSRg3F..eK_X:UT(M9c30-B#[7Z7VfbBB:f+?<=E@)2MgEPN_e:BG92@
MY]W;KQXN&\)CGNa\Y?X2X5?FABJ_18D^4+Re(QQR2M_+(#5ALOE0#Y3WESa5;3F
bC3g.&TW2KHf5VY:c<#DdGaaJ+Z+0N4JI(4):,9XQL./8[c2VAKGD@\.28BJGXUW
7?D3I]-NCUgVC@UAZ,UVI5f[eP]Z+J9U+8L,:J84R>Y@Z#E<)W8),JL(3^P]FD,L
572K134Bf7HRaHG/>JQe^AB.QN<4CIF)RJX_ZJL8:6W)97@WT:gIL\:=L?+=d08B
[N:CDC6UI&L(91I6B6a;_?XA+@I/UMA?36ZA\aZ#0QWb.d]^XPLN5dO&RNcdeD0K
CIM_O#\_D))Z:[.5R9[X5B<4.+\2)5C^d4@U48g?;9(f+b.DOZOdPg6WYUHHA;0;
)Q69>e.aCLeS(H-O#Lg4B2,UWg(7^R,/aNd\ZZVWB6FEe3J\H59c+c^@b98_RW;4
_30PFVd>VWc(gU:[48;.?c\[M:KPQ#ED&&)J=]fQcNWQT2>91L^a_5YA(aBP<56:
[+#7\PQJV,+a?9-8f3#4<b@U?HW.(JXgO+:=>9>GUXCA2^C[L0\/YSUAFG##:0EG
52BFJ?B1G;E_FXL6TRSJ[,2b=KXFK#VQ3NGMAac:&=Xf6DC(Ec91N)F7.<.>KF+[
Q([a<77NReRG44U<D]GX#B6/acd.B+[U)e9.\_/f[Tbae6X5I-9?GQ7LT\5/E0W5
RRCJg][WA-(4?Z+LZ/]gd;6]7QdGK6)eW,]CYOVLOJCGST@OP9e-];[-:;I2J&XA
MI9VT+26ZJa.P+c,,.JRbc#a1V8bL383>EF-KN/+D=M3DZ78D&]1L[_KGZ/K(EW;
f0b:XX9VQ64\Ua5]/4_g/#WR8?9b@e3KUW7U)ND0Z1\5.^ZFe2=e,]L@U#V.=7b5
Y9ELL/f=JVZUC?:9Z+b5HYP+&]?1c#_@BSb2+<SYRU]U)I5,9I8gC]g/84ZJ37OU
8K--&OC(Na?41g^02&].g9L[3Maf#;)W5W7GGU4Z/EP.V6V43Ofe-H9Dc?C5-g,&
,Q^43F\25]<L)=5L_V>&M@Z\10FD<R#QaRHHM]SFO:a76[f3<4?_O,&Rc^8D5\Xd
F;+RRIU8dEZ)J.HXG8B+3D;Z[10>&I<Y+,_C/d2e0d1Ab/,K&MGH0/Z6WX_@URL<
#D1A-G_Z\E\aI(>4DPNQd]5S3a+NX_+,,PPDM#ZGZM?X[7DB\dW(9GN./7)ED[7^
2:CJUfDgML17M;=.\@2_>GS16101^-NMI5O0X>>ZT=LOH<[HAWX0LaBENYGNRGI<
3FE#M\MD;4D+R^^S1N2AGSA\JZ()GOGWaPH&._]R:S1]_-:N[C<V94E@)?-YQ7[@
&,UU]CgUEF=[)I^UU9^e2Vc9U&\@3gT2OQPM<UI2a(V20G+T8g(5Ia:3G_-f1@_-
^&XZFPZ,b5OL+>\]Pe];HMN:LY+QVY)^+M\OOa3Qd+@Y)V,N#aRW/R[25+.ME]@0
ANTN=8?)C>ETQRO)/R&(Z5[efZ\;4+@YeNae5>MX9/RMa_Oa6Ga1<5-Q+JFfJ,3G
bXMV8WRgd/@X>N]L:+d(VXKP6Mb0cGH-e3B2GTZ<WW@/4SDH[>D48P/&bDc#fa_1
TI6)HL-X]#=26MR1LX7bff9:LcEWY#Z3>_R]c+gZe>^VT623#J_/a3,R8\/Y[T>D
L)[JN63@C:DaT&],4;/M^;M5Id1UfTa]UDG2]L(eB.LJQQ=B-J+X4cfX020LBd_\
.TgLYPW8Z87&[O0\6I\[:.Agad(;VSE:<fJ^gg1)G)S;P4W4)=9:165:6IgVa2>E
4X,/3@WXP4XRW]=5MR>S(4?W0R5Tf[VXfX9[d_<Jd<KOa=H84Ra462K2[93+FI)b
eTU3Rf3G<X-]=BK-6fH6F8RN_A/7VZ+=B?OK<D)Y^(H_.YQY@LGTcWE2Igd=,d+L
88\NYPfAd/PN;aI;3L]8abL:(_C93MH+H\WTI+gT]\6F5d\>JE_cF9DTI^.;aIBU
b,([BN#@<N?;<56&.M:#Z.5?<\?.QH->J/4dN84?RQ;=IP_C7M?7=.Ubc;@aG8XZ
NP4EdCG=8Z17TeCK,Ia(D(?7(@SA,2GWWeTgM6@A+B6G5Z?N49>_42-[Z0Y(A]X)
cdIJM+/UcN-_JDKD\2OWIB,4e+_D+NfX<XN6T_[DABQK9DbW:PJ5^YRg:]J4+6Q&
eUD10^Wa[MR;A\4dFCIe#/AQ.8U8YN0/=8a-Q04A.ZdD+^=]M1CTd#XKCB,.M&d0
NcKH,WH>JMAa(,^#WF0+=Q=VeP81A5>U;VRGCAGVH7\;L5JBZ0?6U8AHJP6<5SL8
8IGZ,0d<F_6Kc3M(<A]^PXXZN6_T8Md6]AfJY\CL6F@;LcJH;;2PW/K&?0B/).,g
Sg^=b4-cR+-HHV??8?6<DY2.?RG+ZcJ9K>@c]Uf@E_3Q]FQ#[4;9fd&dC<Y1G0^G
Ge0RS^<34b#97F&,d9\PG91?(5;K/\5d;FbKO#3>U#=T33Y2cXMX@Kg^,\U^cD5/
E,RVHJM=63E,FMEA_3GLYX/:T^b;#&M[ACH,XaV_Yf&77Y,R[_5[15cT.K9(b&g,
M4=DUfWDKQMO7+&g=<S3W\ZOXX70@<P@5&0^WPg[NYIUM.b6[CK#H5<VQG\(2(g?
3S63[.&+MYI2IY[E,B@dde2(YJc/6e\Ke8IF7X==2PKA55dW]BCA>C^TFH<D88GQ
5.JS?(fD3?ZFbGbgVS&gHTZ5<M&6_=Y<-7&=?4>ME0D;_;#e7HF0;9^[36K^8DGB
)@H-g_&8TO/AZ1^ZaUG)EH#F8^cd:]_VHJG/-5&/G0N\gVUQS\YbXY]4Bb8.aDb7
2YW#TAf>gBKP_^O)NZP0BGC7E.g75@e8T#OJ/1NL>7P)8MdV6BEba;cE;]MNH]Bd
@+LN(Te/<^9=#__[WV>VM&<gTU:H]N1-C2?0&EV+B3E]ec9]:U0Y@g;5[d.N3SI9
OL.K5[g.03g5Y@[Eg/BUbRC2U?2^)BO9XfUBZYGR@)/)6-/U;>C:T?e/&+ff\L6G
dQJ>?]J3##-.JPSB85EX(RK-S29A^0=7fY0?\LbcgY7eUE]7EC>eU0V(/&LIF7gK
^0M2=UK-(,PTF>J<#YMaZ1B/VB^SFSBZ\@E5X>7T\^AN/01C:\[Ba35?,K,JgV_Q
-Z_+U0Y>JZ3Uc;3@gXH=X91ZMfINGTAZS0IYX(_I]dMWUG<fSH?[<T[L3^UKVJ7X
=K&&3T=f:fB^@3[.9g3YK.L\_(R5I^+XJ-7A?Hg6?_6T3:I1OPRc68.@<=6Wb.BC
8Gb=YNDWcM#E\DcL+3<Dd8fVZ1>C787G_+NYS:A?]+KPSUU[RTO[-T20B]F58R:a
D.:B2OO/JeD?02=TBZ#bbKM76E#5J5VaZ5<W>7.DeA/9=)-NGRKVQ5DS,:?[cGLN
+8N+P[Med#1IGQO/\J&]]F#+gE[3-KIPe>JYSC&FGM9HRaA7A5e(dR@8Oee#cDUJ
EM#cfFLXBf/Z^Z\Y]+HYF]7f2SD(5/]^_KJ).4>VR4<GbQX7Rd8fT2LT7E@OQe-P
#d=DJ&51:D+>b(U:-LYO+F8S]2\9>:S0(Kd&+E&[OCI(7cUb59#0ad6PIaRJY]2D
PU5V4AOJd,d[NKGR.aF-X7:3\_9>d[??9U)5U&^I:Mg]f&..Tc/1U^SS28L?==@I
L9>UKC(Z@L3M<[S;?aZLEYJLS?&6T[/#;K<.17PZ;=6E0IMI;-G#:+QcdP8]:T9+
1aXPB/QTTQJD6D\VF[R3J-;393=)M@F2GNT#AN+]1[F6VJe-Wf#:;]OQ714R4cFJ
E;>C=MG.WcW9A\X8^35AS^:1^>XUe,O]7;]NZb)=V5/(F3.:9.FF__D)9)\d\1cd
G[-&/Y)M1HLdEH:OWN]1XDS2-8d]W/I\DR+Gf[=>B,,IU,-Ag_K)f]I:b(^E[d49
f4P?cW7FUT3-V)_@R?8EKMB@_<FSIXQ,S?2EC\1cOC8LLf+H@c(CbeQ-W2WU.#4_
<dNa,(D1JfF]2b,E6DVSYgN-_J(7GVDRK3#Kf;Wd/4A[0<fYACF>BdcSfe]+AD#X
<g9.^g:>(^2?&G^RP0RP&)HMeIOT/d4X&dA?FUOBN>W7:[gUTF\fABdcBKdLbCc\
^Y<W&,HJJZb8aOTJGg,JJf>5G;EY5;c7?SV61_M_.97.M<I\#4#IQ?RLE[Zdb?Gd
FE<ea_;@47&,b2&5cFG(g7#H[0LTP:Td8^c7W64QP<;CgI@._BHVB>XZOHS/2T:7
?WT;NPCPc7;;5,P&7@F:4\E(T(SGC\X&_J;-;KNOb][3eeg=WI.eJYHYQ1(T2_\K
aX_BV;W0O=BNA_ZgUd<_g6O??9,DSCHTI#;26KGI-A/J^D:4fN/XGV1/H0T,U+VC
SECW(cNH9V(/T76P2bQZ77d2PbFfPO<a5I)QI(,Y0HZ[?&FN:K,X00dEIb288b9;
&+bg1,B/L.KTeM)J#3f\U<;UL.3;Ic,(F\XL,XHT\dgXfP+g/4RO-+[<#(?;XMeM
&YdC1R6f1Y7;XdNB:/D0fP(.?g_)N>a0eD\W3(;;F8<#0@#/bAL6<^ZUBQ_UDR)<
F;f:eU6<^G(B4B=3;A9SIT&2:D2.:g7T./<M-=491(54XW&EZ^76]BD,E@+-Z.Rf
44HZY9V,JSW\9T7<4Lg)KQ1/7=Eg,N57>\/IKff7Sb=#7Ze3Z&I7ZG6CHV@1157(
?HaBE4VS7;-?U7JWc8/H@NI4VE;4.>A0<..[.C>9ag1RR\M^?W6RCSI<0GS]KIWf
9/HTI^P^7\#@/YJ0aKLB<#cCIHg^##?#G)(F4:ddEG9Kd3MP^CDW@JR[5LTUg\Tc
DKO+D_)^1NOD)]1QB\;HBIVbJSI2R(3\b_S^Je\69_OI&^@fYEY#?X6N3-,)@ST^
/U2U88ZB@]1C)2R6dD.MC4/1HFBg<\IW4.]XRH0]/Na75]):T):#4KW;E)LMI^FZ
_=W,-_KX#=QFX]/GURQ/CJDA<6:ZU4);&8H=C&A19M\9=I>+?VHc_?E[?FT:db.Y
D1c0A;U-Hc&D738/\@,B&/^87)aGFbg9X^V9J?398;&dC\MW/]A3?9#E02^Af(a2
/a\7M_#XR\C2KV6J)g\e6U0XB&D#dIeb^UeR,G>]U.Q5K17YGA^&dTMea3/U.a[@
(#IC_4e5,IWR1S@E);X[-UT2C.P>A=Z)J&]K1]PW[WQ#2:^QKD?[X(:M1.40)E:3
RQL:MgW7\f@b)FS;fB&-FeI7+g)366##2M5#8d?EYVJ>_4:\_@>aUGL80CCQIY&)
f8@ORbT9_N;[R[_D(PYPJ\c8&Pg^JB5d.71)N<D-9=)NQM^@B16DPW2B\B<NW;.Z
^:gX4cTU3ZFH/G#fQIa3H63]^7#<=c6IKcDY5WK\H,c3+&Z\HVWGP3dK5K/)KVa8
&60.]F:LP1dI:>_WQ?\:9XW?NJ5g^U&SN0E2A<)5RW-(EB&,C8C,3F<Y64&aabL?
;ZF0HS^^g#6EHWP5J^eT;NOgJ/924fJ<=(?\@HI[@XWVJ8E4M8W?_C_H+QQ58<Qb
;-KNO=aeY1/Y5AS]:5CAHfAFXe^S?P3B=K=O-.TWd_9UYPc;H4Q4SML[dD26>bQa
79)R^XR/eCAC]5/IU-f(/>(7=[_5WGU-XQF7c^=c^c>G.89:D\L@U</-A85?&8P7
QXg#9FQPFgS@K6R]3AdCD+Zc^LbEB-,J0Y2,KWH5HCJ,c_Y(P_\THC83ZI4YWdaY
KL[c0,01e@HcC?a#KR3Z7.T;D?Q>UIT,G\2IAa(66)XK:F/KR,9Jf+)3M#E@.7I^
gZY\4#[DCZAbLSY-We7]EK02d-c&]6F)EZ^g8=c.YXH+A/_50@<[-6K)+&TL6<4Q
-.8D#0(^UW0:PD2L=YC(DS1PP>=Fb.aG^Wa_^<#T6[cM0;-2>-;Y_.SJ.#\CMe+\
3EIQNNF1I+8BM;;bcV)]3S?XW/]8E/VH-G-68Ib#5(EHIUDKddg5PVO:]/^=W)7[
\FI3L3BR_\dA05dD(XY9c/7@2HHY+e7M0TcW7\BgD7Xa=-W29fX],)=YEH54&8.)
4a]GGd.ab:8M\<JS[;IB8<,^RV/IUI^T.^Qb6@-E7g2<EB;I&#]dSVJJ.>aTba)H
I5A^?X(Z5aM?CS57\R)7[<G]^T[G;JR>R?<[#8b6.Gc&P71b[(K.8F;b&DFcH;[_
Z?_RVfA0DVE\;1@8a^G#0Q+\V>V\J2],_EJD&)@T1F/(EG>C:CP52S?[>?KO@L]S
TPH_R8Z>YC)f<3P,e81dB^^_f#+A@bUgS4))DQ[U6D.<6JAC[g3QUK>3UCNTUI4J
^1K5d0>QS3Z1c#BAAV;D]gB8IfHKU6c)CeUR?MJF>8OU2,YW=&GaC2-.R@PO0U62
cNG7CC:2KS<Eea540X2KWdU.F=bA-Q^K8?>;7)bddHd;E@]4VDa&+5O)C76b6TG/
[af[SXPT)3Jc^@+[5#GMgU(\@YeEb7B5UK2[Ydd;+0A&/NJK56)K/.gg>MSLc7\0
Qb?=:I?+AGD=TT#(3):[/FaW+@IM:0<3A<^gGJ+FB=O(V329>)?5-,P]5W.,)<5<
BOR(FI<a@C&(f7b,3U90J,#,]/J0@\TP4-=>R[?6IZESF4H;<R#:N:0QSGe_B[c>
/.)D?.ATfC7c[)3I)/P2V_UEB?f2)4(.0)dA8V)fYd.3-1@;</8_8b17HaL3F9eY
BcEVX.gRLLU12:^U8+.NELgT/4:VX@/7Yb>J;Z(b)dg.dRD&ZfXH3(UQ-TWW,8N]
-__^eH^ENX3b()K(LZQ)MLIBaZ__J2]UC(UJUJ<@:d_@14+Ug&S0?/7&7eQS0Ze+
U+^6F<GgF1adf?R)JIWRO&K1@769NRMJ?6b5e1U9)2[Oe.&<8/+\Zd>?4I_#U]_U
,0Q]ZZ8,6RZ97N3-7VP(OL/99BJ@1+IWbgA6\]3R&cU);1dd6&6-8F??F5&LQP;\
5g2H<R<bD]L3/W@RH;73Z#fCd#)O1<65^WGR+-Dc,g);NE[Ad<;fe>YRO>XPF515
M?9Y(\6_8NcbBGO?S6:[K-<1WSR<87P7NB0Tg:d4e1(J;R4.DV8BM_LE+F#&7gLK
S#-8T8P\N@5Re\L^fO-aW4.MR3I<=HaAR-AJV\5(6^BJ^8/B78@X1Q&<(/JMDc^_
CJ=:0f/(U>@OJESEc4T?E2C1,<]FW&ac?[]D3cd1<Jg+_YHNB85^TB?#126(-\3C
.#E5H?(RRSEfWX\f4=bI>a5f+3U;2Q=a4>9/dF;OMA[M;J=)TQHXHa/-B)Z@-@)d
I_Q[9L,@-SGDCAH)D3JO<9D<,2\<#DCEaY+GO1&e2cN[;B<]H:0>D-G=0VH\0G.G
V-9>MN:?3d=>Q.SZefaQ([0[0MbUJK=VHbZb.&;A3#28=GDeNA?c(bJEOb(21?ge
KC2_G6c+eU_\MIc2[(9;TgXJ#d\(<O)c>MRgdJ^/-9AN23YCMdP>.B.e(A8^A=5F
]6+^b.OgG:#SI2S;5UGU,\QcELA^?:#67fD?<Ed3.D5-VRQZJJV)GG0dCHcFCNag
OW@(dLC,]&gHYSPI4M@\^U/4LdA^UKL[XL(-DL92fCUeb<QF>Keg#a/K#C,G=TQ2
II5FTTPN#SJC9aWF:;/\N.@9.I3f;OO8FFZ^DW8Mg7^^IX@0<CLQcbKWFW74H_:3
+^ZIg6(FIbgeF[;;aFP3O]T,:>=WNSc=;c>bgM.dg]R&V_CKOY_QSFIX8bDE^XWA
BD3+A8d>e4;2/#d=K1\]D<fa(GWL=1><dJ9f[T2C&F545N#0YMKTH;Z^=R]FEP&M
B5.JAc^@J)>f+90D<4,7AAU9YPTI:b8TJ;8Fb2cJS8^[:(QV9F?8@U(NN#a,<d,K
cfSSUBg0JgY8_[cW>bB4F<[J?gZ<&gDE&7eP)G7b4dgBH;M.1XZX@A;,BeQK\W,?
1-YQO).->=H_L^4WOFG_;,GRXB6Nga/>MAO/aE.1gc6)J8XeC5^7/R&B1:C@gHIJ
B;J2/900AVBc^=f&7D.?0RR0ADCS6ea?D=_1E;g/>P]EI?S[-JMD]Ea]Q[JL.KY]
MIF;V1BBA-@JcfPUEISET]=14M&_MAX[-RO;V.-I>SeI-RA&^8,HR5);ZVEZNSYA
-(f#]f[:d-#8@5>.O/S\G6=,FFV_MLS2\U581b_+M,9ED#T4QWNdXMNV^7N#g6=7
IM8?--<5^N-&TgY>\(UU(Zg0FP)0SDF=]/-C5:fEO9,Q#E:(D>3Gc(e\cfTcRfU6
g#1,_?7Q/0V35_4;G9@=Ka=ZUU^]SL#=UMQKFRTB<(V;F3O;b@gc?/^c68C\8@OS
60Y<e-A)<ggCX/;NT9/O(Y^]B<TCH9U,F;:fM-IU0[I]Z9L1M/FV#5(eQ8?TZ-O^
Nf5L;5>-.Wd6IR.>[6[;@aEf<cW<OBfC0?SfLf0+fJ?L8<2@+5G]:N(-ZNZCF?O3
F=F]YV(aL()2OP#)Q,KbRA.SO\G24fP=9>^(FR@.0_gP<_6LO_egNL=;.bHRc=-?
0NWb;5gHKLW61)K^H#@e(>QFU(G_]>,L(;=3Mc#@Z1:2+5IZ[>V&:/43gaKSLKR=
GWY,3FB5,^=9)BG>,8O8fb/[P(M[4LW]RPcLW;;cN2dQfT2#B:3#&bJ8ROM3+30Z
E.d&.bG>a#W?d&8VO==.dg=(N4EIgbLE70X^)6CSTM6NOL8T>:?^Ub,D6UOQ/efA
^.aE#Q)OZ+F>E7D^BfIU^f=d6[OLO?/]J26W.fNe5b1;PZ5eX:ccEE?@4G8J0>b/
?&6]MRW(L7N^#YM7)J?U??Q[A;LbILD4Y07f7C9;:JDJeL\@M;60[#1f[g.E?/D7
1ML^?C<bG-R85WKNA?PM#FXeVRE(J__#LKOC8gVG8Lb:MRg)NLMJ\A(R:_LN.=<<
<K4N;^G+,76AMHe0BEW/#d>.ZB@;C2;6+IUXPR)gWg<D6PaO8&OYT5?0aaDc:H9\
aQH04A(0#,OM4.\RJK(+eOU_9@S\@4GR1,<E</c1](TPT6,0WeC5If]UeXd7F:5L
EEC66E6]MCV2]#JL;Y;?f>e@N6BX<e80J2C#B;:U=U9L=+H-,EN:;][IfOaZa7<?
HN>5K?0;R\@A<N+/V3_N>9<YYVB2#D>Ug09?9/bIKCRP.#bGL2=RX/de\485U0#,
;A\6.P5c4T:d<ePT8WO9Hc>ETUM^;>]2[M#+UX_X;#e-6fR9IKN]c2HI<d(@>-/^
9+JNR_CQ0@FVMg)5ce^<bBW3dcA8-A[a82:a]EWD(G:Ue<W2#G_?cW=RHg:D>eZ[
1,^a)e)MS,MHT&&0Z/0eaFZE\>XEXI.\GY^Z93MHH)3WLXK[:[^.#4>>)cV)C2fc
^RF+&JL0cc<>-e9<eTa?O9(W--:+<F6WV;+->V@15d;L:HW&/,<c_03a.bA5K?_4
NY)^W>]QD#UD?DO=\aO<^5c>J-TZI=ZP+/CgYU0fe<I^c)9U&P@:2TN/),^FIOML
G/91f?T#.S@R91BKH;(]TO_IPd2V6]feKJb_@_6+>W_C<TW@3RM@D88IX\LSD#[g
XU7==PG;;b?@Q1>A8:TS\5D@P2M6J#89AQcb<d86@2>NgL>SeP#X/EbD^L([I-;-
YeILE?[WcdY_GJUAKNE2D9F<e@,UBYT7DR\:S#,fONgf(_?cF<PP-8MMS1)eSVRY
>/_.SB/bA;cP.Q11#fWC_-H3S=<Q3NH0e#Nf[D.K;Mce5\]N1S]8>X\cFX6_VZ55
bIM+Gb-6LVFaC#CIJLZIEWTTAJ5;K22JM\6H,:-J]#A/fGbfd+a&O5RbCIYaOI43
>^M0Kg#dV[XAT+2A7XRIU^1:]557g/d5?d/V.B-eP7Z7dWK;S.199cFH7Y9<MP]>
-9Y+&90PHcW6#YG_O_BQgCA3>cT=@,cU>L_.08M&,GD<gZOIeU)RQWU&VTQF2=8U
1_C871)C\+21@0M8RZccAPZ.FQdL[,BZ[<FO7GTZ(5-@D<S+&]?HYgNMf5V49P5F
H=GP4ZMJTY8/C0@#GKa6=.^8A<-1bSOB2M>W_R6:2:T]1YWJb+#@T7M6VYX6U+/7
)8JDLX3Te3W#L>__S0/\8VX=J(<ZB1[dc);[4_FAPM11,>SMaJZ0E)gcGI,_5N<g
Fe<b[WHT[&R[bM6Iedc5BKaVd@(7YaTIN\)C],&(\3He+U;^418@Sc7F[AeKSbD4
bE@)6bJPYB-2S0J\Ie/ER65,;E=^d>PIEYU<_TR\]E1JEXI3UEGF_X+P_d=eaD@I
J5[1#3F>ISJ>6\6K1F4)6IP,SV2N^&6\Y+(IeFNGGb8K^I^@(,7[LB479J5Qb<YD
FSZO?H\+Ye1V8^e?RI-X@]Xfd&\S<GVOgKVM8(-:Rb[@7fP1DCJ^A4]T/J+FIT_8
[_-#c;/K58<&ab4U]47bFZd3N@fH/gAPe.?.&9:Q,2Q0^>ARdLO1R7.2FH1G9aHa
_-#e=YJ+1-d_M7D>RHCR9K=BYA6c/CN^;f##(GN4E8e4:?G=]/3T<,BY]PcT-K,S
\^P(7M@1Wb4T2)Q#6a@e8-QY^&-]2LS@fQ-f1/8&c7T)WSY_77-X(a)]Nb\44g.^
3=G6DLX+>.@@D>3\F\eP@.[_NKA&bM8&R8CHe&0PR2_WS;961)O3L_AQVLD6/I4-
C28=40^7c\^<[N#:2gb2JU>TZdS6(W)aWRfL[&8-AN?R^+&#APOL<T296H7Uf85_
#g&L-1[D41a<F#XUfMI#>cO>]CM]..T]@8<>>(+[_<SU<T]QG2Y8MC0Zd=P,\)<9
)C]7_Ta[L9K3?:D?a7B\0=egUJD+0T^?K<IU49#/^+71K[RbL78O5E[-1UU=W>BN
)YLP0KFZeae3MYP<W#f<aMS&(M;f\M7ML8/dW)aE^Z\54d]V&fE1C6.&N>Z//_J[
??H:?Fc_<X>g2.1MC\UPbHE1/\T5\4IS@VSg[3KaTD2gF\25^]LXO1WUFc&0BYf)
I<PXNRQT:dYc+-M_F]SIX3Pa#A6O5CVLJGOee.2.dHN./S/==:;)^>5M2@5E\YRY
Ke0ae9S6EB^P]b&M@96F2>CAUJTI0^(\G\P+SM1)GO&T.Z=/@(\HSa=71fSg_#0g
&.\90IY?]cQ:g,NE>V9E[Jc=f,Z3PJ7B\XDW+@Ya0EgdZgHPE3ef_+_VWYT2(-d7
]IW]1S0L>Z<_e<Q=ZC,(9YCVa]<dE#e-M;+Y:O9.)T6dZ5CWU=.C?dc2LMQ:1_EJ
/@WDL&3JCGVPC[G81RNe8<6Qf&Y6B@<9(>d]0I&<ecf7Td\7E&#/Qc4F\@g;?)1/
)JB=IG2;M@JD:ARYJd;Lg<(P(#aaFMW=#RVMMX62\7?XFJZ9T.T;32HT(Bb5A60E
V3@^9b@K-AXQb(@=5I-,-4,QAHH-(V)VFP&/R7)<G_C(.^9Id/ZXD-K7Z.7UMaaX
7J2?Z,\B3^UGWE#;9VH;HKT;#H&\W336JH1gBBbL\B[<ZIGTG2;@_HXUD4^bIAZJ
)#9[?I]=LR:8WT),/_)VZ9K1Nf?T-HRW3eC0cPHN&9JPAf=1@1+cW3U63-B,L_d=
7+48f+cKG(]49e15EQ]f6JN3RFEgEE4(<4Q-/f/.#fS9bK:H@-1D9.^XQ=TLM^MS
5+BXPcHDAGLK84D(,96D?H4OO2O\XfNe5JV,.BQD<WL(=TUJ[/.eZD\^3;G^;cMA
(&c/G)EEX1Fdb:&a)NA#N(]XfV8ZgH4JMQ/JcR9GcW7)RW+X1,Z+abZ;29U9)F3H
,OHNG776E6eO[9QV)Y/e6_E+Oa(Z)F>Hg<I=d5CZ=^.8_1X_@aNX62fY_&g@gJ#6
-A(I6S9OYNQd-\3TG=Ub(MdYe[#e]JZGcT(BZJ+=F=Q.Ec>0#F1I;N8M(09V3OUR
/2Y&;KJ+:5L/IJ8RN[ebW2;AVN>V4UcGZ3>,gS,6L;ANO1J9H=ZCc@aQW7_VN/WO
)/_41LYKRWQbIN_JR5I&Vf>#<13J0C6(CORF717Y)VDU><@5JUB#M[SNEU6.&\;F
]VV;agaA)0#C2S9?7QF#Z;P>gcRb4U=MZ4:4a<;F=<-,TEe.>?8?L#=D1MJLg\5?
)K;>5-)cKdB?AOJ]8IV>HS;.a#_V(+2C8Q7e2K)QA+2(;Xb3QD[KI3b882L@6Q1)
6LO6X&>2UL>2+.HOH)d12A:=.-VJ8R2:OIT9[.K^.>U5fMBY<N==JAGCPZ_\RF&W
e/RGHU2eCVec5<V?(6MOX2cI=A96^6M6;dE(=Rea8bbY/O<46A+\+C5H(+E6/Db4
7;c(,a_>54,bc,Z1DAXL:X2;d4.dF-)=S<_MRP\]J06eS;L<Bd3OD#SIII)QA=1H
,M4V=#TVbT]V):_O0^Df4I1;P\O8/I@(^HON.I.]I5OJ33_R5Pf^Y=&a=\bSSTf_
I^//523:H8B58?e7F_6LfHUY_fI7Qg=_&J0)M(.U:f]bSQ,]6E-.86&+33(g_Xba
)52/25ZgM2Gg8B^NOcC>a:04eAN55EcK8K,-P8]a1M7&1ePQ6>A&19?6/?66Y88N
OXMWbI>>DG4S0?S_SI3/&e/:FeP+W+A.<?H_2W3ZZ&4aXKW:KHQXSb]Q#9[Z_)5O
>)IG#NW?>>bXg?>5T1Sc)=La>YLG/0FM>aO[HVDce#cN>^]F=2c[6Q)fQ=\;d@(;
48J(M1^Me9.@M5g]L.:^?8S:E\]Y>02P13@[O.(L18B6O&>0,1W2\C^cIe\ND:,J
[e&ECGVL7/S_/_+&FE:S0]JJXPY8fNDXD((TB9R2VG@UOBXL6<f(FcR]EWI7ZEI<
W)_P)Y=R5I_He0)dP1GEZd;_b@6?H.7OZOI2A@^a?8/<bB&</gF7YggPC1^[L_,E
B=^CA\QbGF;AI7G&.3M#]MdWEUTb;^)&47UG?I:EB\bTUMKK:dIM&0GTK^0^9/4=
ACS/RCACc1.U31-2SI8[,3_OMe\.@2W;4F]IaSTGUQ-eZ.9;VNNJbG2?Xf/I;\L_
L722#RU0&[54eZ-9&QL7AE9Q+/P1CIYFMO9B(C_\K<cZR0KgdO1WWDbc/+a6WULG
1/0Y1T@a8fTa)5ZK.)R&9CT&G=4&CBZO:5FBe]D<U&)5(PTg89dIJNH^Le^)RXA.
@2?C3(aKe.,0XS_Iff>I-:Ag1-#TdZUFgCG\W?P+I^#-O6>&O&W,XMd+01X,2ASW
Eab&:R+(N--E-YgUP+=J3V#>&DN4c5I#bLY=D6@_H1Yd\\&-J&J.>(dE@25M&g9-
2bdB?]-BY\e^9c.:67B4bDWZ9;KF_>[XecL?VN&(AVWO)GJdLc75]==M,[)<C,HH
AM.AS23,RF,FHSG0GaY?O#-B^DE&8cB)=2<0T#e(&)46aC,:Nc::GZ\MgGg;KcWV
L9VWGa<R9-P/6)3BZ&a.\3d)Z0/K>72]@1=QOQcd^IY.\9RW:)+(bZVA=f<gK</_
d:F<Y>UZVKd6f\)(5gd(EDMQgUME-B<f6;,8+#V]G><5e11bN_9gQ-XgR=[EOS.L
L/Gf#W,,]6#;XH>/5188E)A\XNG6]7B=2(N4H1DH8;#_(EH@Q&G_f_-<73FXLTZK
#S=H85S]Ig&()QaLEC\Ha050Y1;Ba[U>M8@]^X\44g,<.T5V1c8N]::g(YX>M?&#
eb)@CLY#X4e^0Rf^EOd9SV[B(89,cI]RZTTLY>.-Y7eXZ)aD&&W=fV.,<;DG19N6
_+#8;-=(VN=:9,Y,)2T&7LKH_\=[Q&9Q#F3^_:L+Z:e-3+<Z[GI\+TJe)/UF@E5N
_##Z\a;.>])0bS+A)59R\5+50ZCCOcceSE]4\P[bJ]6=VU/_CO7Q^@9]Z(AUN,,E
6G)7O)HY=dOW#R+9dAD3(]Hc8T?J@-)XUZc?R/HIS27_;VcLYaM^/ACWD?O:\D?L
<d/(DDS6]U#0U.+2>U42[[(6c7WV#R<#X7(60_eZ]8/QI^9.=8\X[5E[-_Kg7\B>
?V(VX]8Mg[OSS4+#=-1gE@2SQ47-6<70@=R_b9X)^YL@1S+Y-D:d0N8:PZ@.;WR-
=[C:dJZ(J=(2&_UQ<VMSe;U1:WLSHd,VDJ?5L;1AIb#H6O->@aXLU\.g\R@Z=N<b
U;QVb7D,b,HD#SNM3SKJCa&>XBBO.,KJ.&[,<?aVF+JY_2KVBCH(D0YD]C3F;&U&
[:+\[S80Z,YT(&8AMZ9D05c=9@[SY:J?N0/g]WgUD92?40F8N-9[fA9JbTd_QY#B
F-d+-2=A<<LY^eS8K:X9_0V/PD>JbJI^Z1_>:ge_\BCaNGY;.US>N0&5-Wb-NERS
@&?SH8C[I/#[FF)9\.e)&IHAdeKL\FW5fcOCBP<KD>e;+-e>a&0F>Uf1d0.0ZPb)
[4(BN+S#gceH?V9XaH+A8(dC6^g1[ZD47f.F6P/Q_@SF=MDF8JOC;ZHb3H>AU4D>
/QCVGBc2X2.SCR#-A[R1fWK_\/HRS0O3?)eV_X@NGH;>P(]LH)Z)VD[X#S&eAX\K
8\Z?g+2_K#dFG[DP#J,@W.fV^5BC+/agHZ:\70#:Cf@L<3]DI9eP,2;_8a>e5GB(
EAWD^80HNgHfA0bT([64Pb&[RLQ9eCeDL#HK]&.-g85[GY&\#+KfP80X,bC3XNd4
&Y.8>9Nbe902J^bXSOJ52\MTZ)Og+#5[aFf=b(50S&1dMEI@?22SB]^5UdJ#a4OJ
7-70O?g:GQ(5\B[.DSH87g-Jb/>9YG^2ZP610[MdefYb^1^GK<aZ2a7ccL)5f,2D
U))OZ;2W,Ld:,#KCMAa4TJ<=cWdZJ5L__H_f6a(@2dVD2CO=dL5&]6+2LYDJI9G.
DIF_1Z^fZ1:&e763W#,X>#V4)PC,aFEN4QI/[?HGLVc2IU47W?7\=S2.270+&9@,
PATJC#_W\_2X?g2GGG0ID3&TY?fWN5;9IS?I+^Wbc1@fEaSNf&,3ONegYKPKRD#S
gI)&7^C&_>H@/_[UJ?bg/b&J&I92,T1VK4];d=0^1KEMLP?>eafE9UU#97T2UD+<
YIS/Gc(IUg.M/<PdRJ#8b3[2;2d0K5U:LHZ5L_2JX7WR<75_^>O=6CNb-=YBb@;?
cD<U?2d<Ae)<ASRVX-\^JTLTOHF)43B@Oe:?a=91[G,QH81Jd]<=dB-=gY5PaBU3
I5f&^<S@cUe2XJEL?X^#WQ13Dd;bYS?^=,Q2Pb&_&Y9\8aL[<cg.=@#a5X>U<4b#
4UIeO-QCDb^<TNS].LN>B>?]\HJT,8c;bI@ADOEB^aIUFIF4e^,EVC[<D=\^5ZI\
P9TY7]QU]9>d];J=aI1@g^7+R^(JfKf6ebG,4@47M6SK=eFT5E^AP;W\U;HA4U&.
]D\,bNeQR4ZXF6NV_0RbM=O)eEF)Eg1T._ab3eXA(_^Q==F&FY-4>)3Z&/#<PE;A
;0+4MU[U:2C;fY0?.S.e_N)cZ>2_PBa\<X5)_I1dL@8[V=.^R[R7afFd]&-dGR[-
9AT4ZG1\F6,H1WNM;N/8#::N=:71A9LMEMa7P&1?gU_c\K]V(Ef7\_@[d7T?@&)G
UV&F1(UI6JO9OSU@:L9\-/13HA7[5A3ZULJSP/H1R,P)L@04)R\eG3;L&?AN_MTd
>FBF22IgSW;B0dfQH,E)eG>);693#>7HI\3[JO:4PaMEV80;PRd],Wb):UgSF1O6
);WL#5+=1WdZU_gVZ]eE0g][?C8be8Y2Q8W+@QXbV_S@PgfTLZ9e)1YV]b,EIbC_
Q[5U7@]#Ra]UDC&GS/M,Z5&4=8cfJW4BC;J1)b&VHg/6-66AC:P@LdJN#N&[-#6T
<IXYY#[ZPDaXfS^a\D1](2Gf52(LHUfS_>:cYQFJC_M3.#e?TgSC7RZ&NL_03<[a
P&YaW(<2T:0Eg)K,BJU3V?=_N^Z2JA.Z(29)N@V\[THA;fY9\IT7=Q.3M(E7P52J
GUA&W<^/]O&-BNP9[XA^H@B(GXIJ4,7gcIZ[N?^M#,.L)e/I:EA?a&WCD[8We8OP
#C34W]):Cb=B(#51e^[7;]7H2/K/3?[>G>-:O^.PNe#[/^LAI+VM[GWaYbDMR9H5
UdDL5XT1ecbdHQWWE)DR<fg97>G8RZFbO0W\&cgC+G5.59_[1QZSOXD7fE\(.R@#
Bg@BK:\,,K.Oe/>V8],4>0-B:WOf?IUYcgIFYD#L#]Y@a>T8&bF>BE3=+U04c)5[
+9fUQ<#SD&-;K74LLI2C_H8cF[/;QA<L?5b<_>C6dO/1OZW6]/fU_RHH7,S(#:@I
#->;/51fZ[(S#P3NUP&.YVZLTLL@74AGV6\#ID2a_Md>+&e\)P>9.[82GEcQ1N3Y
^1RZ2a-?,g7;bC\=<3-ANF@3H/V3&B0PbQD^ME6UO=C///<_IEPN:YJMZ;2;&-AO
6c#;<@WPWdYY.dZ37#>WW4J+_92-c;3U[&/3+0VB:Yb?ZA<_DI;6T+AMJXX?HZZU
EY6-Q],&gKGSC8+QXP>GV8U._cA0\HO-7:/80^9[&c=JJZJ_#4g\C]\VFACEFW+K
RgD,GVXaE)D7SR=Jddb&fWI995[06YEG\4PE8HEU.&gS6O]@L0gXWF9L>)_fJ@(B
//N;/4,)UEC;S(97VJ)S.I.11>4=DFW(/C&)#C,Q6@@LQ,P2KWUH?;(Dc+^U:Y=7
Dd[)9ESaTUB8GSSfdN:H4I4TS7N6>^Y]>-8N[RTGJ]2F/Mg<NQ,]4Z/6>8&MLI1K
-0RXPgW3H>RJ#PcZQQ/=c43A<=9F;+He:?[Jf7&b,M3&_1BFTKgHOD91FeK@)Z4G
D[<3?d_CXL2F/JV2_,>@1fPA<FQZWdDa22.F6^JM5fMYS-#Y\L?aY@W/?2(X+IA3
B+c[R=6V\^@a1:2bd5YaS/RTJC7GAY>9PWcPJCf/3E1;96>Y=+FB]SKVE:>L9cDJ
5[ZV.U>C5CW(Pd(8)>X26P+#2eJ4D]eD.Z<4b<,>KJ?:A/eA5c^_]>YQ?#2?&><Q
FAV8F>B[34gVHO,QB.,E&dG6[_MI<QHY/0S-#(J]256)K&D;7//KN\/MC.IA/(1;
1&eW7]I(J?_/8/WF,4>GC+JSW\VZag@A)-MF1_MJ@,)X6U)>4J;3fFgNc1>YB\2O
eR9^_8fdd8LU7e)R^.1V4AeN5SHC/6JT._#P1</D21b/a@OG9QLY;O6HRGgaagY?
[]JM(<M/V@17??>=)WQeW)XaLM0O@&D4O\XT.;,&]2cJ0&^RLZ:AJ?\UAP))1.5;
+7@;e9(^G418C=V\#=GK2dRE43FCA7&5S_8<=A3Z)^SGT,Nd;NJdCWdBUQQS5=7>
U\@9O58f?7PC=B.LV=(>R2H(]GRIMB#H0J-ZITRgU;UI0+(05c+Gc+>aV[0\K6YG
;@=Y7FJP8fE,=d8PMgI>_(2M8PXg:32RT,QX:Wc.HO&-MT\7CT@a5ZV?:aO1c=KI
C]2+I8(:)/HK_2KN0/9V061E:T/WF.ff#F70d8eOXbaX^+eE3e#^IWT0b-IS)/W-
2SY&X4T5dEDJa>[+Cd5RaXE1MINSE-Q5S;eW?9F:ED#>eTc1_+dF3N^VMZ-@\gL.
HC_D+da1&g(T\Yd#U@-Y-I[F,QR3LB#85/06G0RCe5G._2A0T7Qd9=S+V:,_KWSD
#B(=)SJO/6R.C#ZdH#M7dKJH9KY?&,cEJ+fSXL@d&.Ea\ER@2\:G/DWTYND/GBXY
cQH6XPXaV^QF1:H07J]^XN=655CV;L)=Y:9UaQNNZg-KeYfU#&dcNX3;]QW73M>G
80K1EDW#\>G<).Tc3VP<:P\))?U)8=5-[R==:RS9?P8<BMI[6C\Z;1P+-9I@=?D>
e09//JfW=4d+6)FRQgD>SefJJKRU53NI]f[3fe163H_OX[b,/QIOPO71eQbX[,;1
9:ONJ#_3^EU0S,O-FeP<:6HL<Z3-9?JE&9Y::EeF>PWf44:MJ+H/c#+D<Bd2bb;5
ZN2-HfU=(;9S.c4PN@GJ-ZB3V0^]bF]a13+Afd83aEV,AgA&=gYd6Yg7.QJO1>^d
f8[_ccB9_)MNRH2eAY9C2;[S_&c)#;OMg1ZCU0(6-Q90LQ9=0Nb]EW4a9TcN8V1/
=\(R+H#Pa)A?,4VB=V>cNXf(+?CS:UcOZV7(4+<Z#)IaE_9.]f6R5g\7ZBPM=1^?
2H<?;eF]LYMNA<#3dGd03dfO_NAOfgP<OV,J0@(98W)J)?f-29BNGN;gGCR_dDIS
K@L?>?O^/8A/CSFSO8,/IT>LG<_aB#>TOgSG1=c27E8dD^79Q]-_6987;fY076=;
3?dJWJ,g165F)GY^A;HSgdK#9,1=5MHT0/>J<;6PH.-H/)3KQ=-9M2\QFOc4?4^e
R<^Z3?#><=#b?AK4.S^#4):)d?S<gH42:1IG)-c&6^L.K<A\&:4@(?Gd1V0]bN25
8W=[eP-LRg4dF2(HYL@:1a(3..WHBT7J=Mf#32caSP8OgN[RYPMHC9]@c_UGfJRe
#.P[(_I^@.?4IIQ,A^G&7F\HeUAWP<9#23#[.&.52GIH5KU+63FFLD69E(-4d_NJ
9?4GQ63Q9R1&AUH;,OAU8V9c/\F=+;C:FeO\McM4ZAVSHA6d^CFGQ=_9R\DaZ<P2
(K&Z?E:[Jg^HFa^Z@&MBG25;2VON6fB39d)S:^Z4O/H0A8X(A>E1HO7JG[C;>c2a
MT,8-Fd(F_5PR));HCXZ;IdXD[e[g:N(0aR@_dV)aS<UO]?A:6PN7:)RcPe80D^D
?;8;,\Wd1TCEeH)TL80\3+\A]@#W35O0(bCU8]I<O-)T]SZ_;BD/7MQ0P]?17e>@
M-0F5GHS4],PJMT9=2276aEXO.e.ES>2@DE5P,7e_-Ve-FX;B9F0<A7HbGf;VE=Y
U;Z=H726883,(f4eN0+=AV7EPWd=+3?I5P=#G^>2]]M_NfgGcN][UG2_CE:c(e:;
cb4XIH]\O;.33,>6fGeQE>3XTX56cYPB6#8QC[&K8dW4SaJcW7[@D&^UF[4\ca>_
6HP&ZGGg[:,8cI_5d.^:YJ]K9,LBa-N#DPGKIaKUI(3=<&:[YAHPJdR?cDXWL7#6
Q[#NLBLT&TDY&=I9&a-8-DLc)>dCT@[B^a7M67M3X5&VV_VWg(d67<PVHO(:dYIT
]&F3+\bKgLYgPI.D2F+O=LR9?RMUZF7ZdQK[X(/LZ/?.G=:g,D,ca:.:-3R=\.X-
E?SgNSTV:++-T]cF#N7?1<G(044M]+[I:,?0YX^F<+DdI);#.:2df^bP1,b1GQ74
Se:ca.(VHE4+QMP4:gS&\E3ALSY7;9K@A+&W.41&QDFKeA[+Vgg;UNSE;R6_^,L[
),_9,W5dRTb9TRET4-\S.(dBF6IaRbB90)_=TJ@)Ag\U8L2e/5A7;FM_LQcMNYT]
)HRL#[<aFV?WN.#&)GRL;A88]E\WMY;;ML:aX9_&)Ye#c[KcJC_>PFV,D,UVdeHb
fLIBE5b7N660^(HZJ,-[e#R]#fA]S7EZL&H85;[X]+#+XF2b2^]:)32HfSN([SN3
H.<(U&0=[96#9gV#K_0/d#3A02-6Q35Acg#DgDgAeb4M#Ra3LTHH@gE/&LZIeLUX
=FE13_RgS7.?fL\^3G3#MNNQK/e[LgMTFAC)IP]YG,G+UP#TG:H+,/I4TFa9;JK[
Oc8BPSJR=]JWSL.7OEFg57-B]OCcIJO^?0-0L?V(SA4Xg>b@3fFf?<\Z1gVO9Q3?
eY\&?5)5[1YI,e#^OCg/cWQ.EYXe6RgUD]VN+]@YXH:^=P>Ne>]W6:B=+V\GG>8T
Y2\AePbRM_W[.JWdQfNccc+FJ_U\CHEP2ddf:dd?/PQ>&US:5)f-T3^K@[gBJcWY
>JPQ@TNOU/E3A<P=W5+aX.1RI44\IWS@:^6JNe\dX@0)\XY6-&TSAB+F4:f-;Y:b
PINB#]7DCY+B9/b2CFB:HG,HddF[E.@fRTSC1)RYgF1c;4f^XA(-TAS)C)Q@=7>_
Z43B7)J&K8R?EW45Q7SN6M(D;BJ\W,3MI,I99.QZ6NJ-5X9\3F5.35\0UDX+a5H.
VUCC,W=>>3#9B,0QaEfLdV/VB/;CNZO933&NgR^L3=LeJN26NN^b,70I87T);WJB
Kf-<5^V4\R;-KG]:)D#+/V59gQ->gVR]F6Xd6KETKe.?LERV29[S-2T^g2\If&55
VY\C_6g;,B/TU3F\XNY1Y2^M&D)aO^5<f<Y)FeQ<H;6\cM[&,EVMA]JVJ0:.KLg[
3R5/K//?V_=U/96K(F1H#eDK_Dg=U42<2#P.5b)f4A6GZU-&bgEF-5gB#&,]a<Oc
,DJYLS/0)a;d-5eX67=5:-?SOCXA]C7AE+e(Y@fb<<[[V+J(W6.P.XWA&QRcMTHO
K)+U_(Z3dY_&PMZ8B&/:;B9^BNJLK9FbB]8aG^BeB#5<f8?3P<Q]((Q=E)[-I>6F
[69Id8.WVMM)@f65K[aUP\a3?/9Z+KY=&NV0TR:-8Z:ZN<b3>+4P,@VB&Od3E^fe
8@R-K7SH@43^T&7:HOg?\0C#L1Q;A<KfbDNEA>R]Z+EWG#CbgJG:,/9=d.(5KR[a
&&fSUgYH37aZC(3;+gb10ZRebbYbXb@c(7V<DZY:SC\f^F:F+T7B\YCQO#J_G:Z;
&HNXbZA\?1JN;@<(:IJc;>gZ.<NV\^KZOP^+4.ALBC6W08^f3^TDXDa=H[TZc@1g
N4EXeeK[U[9OV466EW?B5Tf9KZ6^P5[a;Jb9\=A9D5V>(Df_J1Sa+_,^CMAO[g&M
F_LO(@Bf]E5f:I>[[]H]^)&;CP\dcg^Ng77WeZY_b3f2YfTFLgT5TX)6P?/O@K??
NH6caB/:^]:FL.TTKb&U:>\QI=ACMBH.,:3C&?c8QC=XRf>_4dFCC^D^Z3FR91\A
7X[/d5e@@c3]J+fd9+M<bgVT[_6@PPf-gDI6WJg,C[,\I3#,(Z;0I3gHKDRGK2b2
B_g?G5-6D=;TfB]d:7X1SfBG0^&H);TR4OBQa>6DIE@+=[16Zf=/EO??\7\b@,c0
2&H63VdUg4[>UG]DA@G?2_RKgTbA85:Tg,@OJZcD1D5B5K-]P?]SQH:[))EYB9&C
bGNC;14L@F#X3XcdQ,^6G0GZ)^^C\/@IXGB4N6CXZH[FAZC;:-PCgB+C(#5AJGH)
@\0E?=RUV+2U3^U@@eEe)12Tc_C@-FU]0--NG)O.G[<1#AQL9_2T)J&K&42Z+K?F
5Ba2<Zfe)X_>eKdWZ0MW/[KZ(?,V6,?K\M4O<c,(F4#ACW[GFE+3XA7UDCOg9K?=
0ZAa<5RJ[(D@O,>;eSg[?/_4P=-dH4CRQDE_:U\e#_(BEVVO?;_Qe4DR#H^5Z)@+
29)KR=[3Cb#ZbTD1+4>A)H2(CVGgUSJBL#BfP0?efdVJ^=dE/IRd2FILL@EJf37R
9WOBDX:b_K^IB-+@4L.F42-P9&QX;f5&gG0fMdgRaTM,@#3cE2CP3&]XP7>,5b[&
SMA>:?BX8(^fUK@D#=49dbA7>b_C81^fec+L64VTLVb,J\63P&]Z28?4G]Uf[f6&
.0Q0IS]/[:#6HfR-G0,H<ZMA=JDaUa4RYg.fP6.:SDd-\]Y:E&Z,#V])Q0ROBSOB
.(a-SH-?NeLcZ-c/42K#8D(eB(]HSaUfZ[XO_d#a86PM.4\^NKN=QD>;D>H#/U\\
PGd9Mf)c)Z6RVd[[EK9\FFBQ?BV1edS9Mb_+_&7.AYJU8GYKfEKPI3BR8Ne[M3gf
48MS@C?-FKg,#ZUGPC+10Y0[KZeZTC;#3-D<\3b(Z-QH&6PJ=3Ef9Zgfa>>#bBJP
28K:_a#XH\^ff2[Ib,.0;:N(c3&-K,eC]8M4]\=;3fOVK&^K@SU/M_8]A6d0c_aP
;YKZJ;5,KCLQ_6U4gQ,J(JV\Oc;#+R/[G+fPSg:H?6_?N[:Z,)Y5/f5<\):Q\XZ0
8;Q76FK6,LM=gd7G&F)8[FegVMaI7AcY+:d>V=\8=:MP&RMfPN>;eT0L#U66a:F2
cFa\DCFMD;d^-EE1d5g,<;[-CS<;T^d=MQ,T2-=Z#9I(KO+V+6=f)CPY-35KW0c(
UC.<+4TD9]&O>6WTZG:<X=XgSFS::E#L+ZJ0S?&L?[HV#\^KQT6-(YF52[@[(aII
E8dK25[(H&;4I-WcQOWH,<:RE&e\[MTY9Oegd;Q,1A(II9dBbOeJ3JA0HNA<[gF4
X+Y;T>^5[WS<]]LA]d5.E0LbHEUR-UYC;FL@9,\eF5MXE340J82<RZN7dI-T@aP5
?(Ab:\ZDc\H3SW2Q0O[E7VJ^NLFYB:Z(\8^W?G7Kb&XB(YP[O-C;cKgED(a[I]NZ
FB>RaZPVJBYXE9QA^X#X:]#K<\3[Q1?&XTANIFdC9d&I9:J/)Ya,GLYTV]^NSQ3T
Z1::Q0TLRc7M#a::W4KE3QUWRTL\5\_\D=U;_@J\Q)3X_c9e&4Ve^KH&EX3g:@F,
9\0R?FP1LRM,=JPbae))4RaG4f#M.F_-<F850&;8_3W:C1RF-R5g-\\;N\aGg:Y;
:@ES.Z7QJ6T,b[#@XOFT=cf]3/F^[JAU#W<BWNE4NL.()R#@UGYT;YH23&_M6&:(
;.A]1#JM.^;.JM:C:Bg1++>_eWB\8.[,^bH)5IPc<^T\AEJ)EWQAZ\Z7E6+A\La<
a>7fTC[.dIBH]50ffV29fNA0UMP;2<0(:I(#5IN\&^SL6[9\QI@9IbU2J9.8R02U
6RF#3INcVYDPN?6[^5AN\gUb.81e\O?OS<QG6DEeEXPL6Q[;9[Y6#R[@dXY=dUW@
>/[D[O.fXG]+?FZP=dWQ[/^>)2D36Q7IT010^f1SaO.87KLVVT?^_6GZQCE?#d+f
U?#GEJG@_bK<fU>C8WFe#[()WQ+Y@2&=?a#5.BLT/9T,=2ZNSL>dGC95684fG@,;
RIcWE6?/RHF=>(UVZUN&AT=FcAePNUZ0[TNIg\\JA8GNMH<#]9a=@K8Qb;#UE@<]
</&d7RTSB<[D-&fcA_MP4c:EIY]MQ,ES6XZU9U\-RY;A_))U>\dSQ\V7YI@.9a4F
XL;R?\)_5[b;X#)/<_Pg0_\74g##TJa7,CfFa9];W#<KXI-Dc0ZZ7b,0SfIO?Z./
fR@ALLX;X(UF\MCT3&VT2MT5(gTQKIXb=P_XB;W7EJQJ;STLb4c5Y,:aH\IZM2@K
&[27Ace7F]SB0[->>>a,20=AG.4^4/<^FFYc::_QV@8V1H7LU6DeFM#N6\M&\R4I
4PA9W-KJaX9/OIF-WMW&(cGb?g-3#JY5.04-Ga1c#5FJ@K/YR,67G1S>=/g#a2;V
;X^=0W)Be]G@9/<A[-:gZaB3-(Y71]TbC-[D-E#QN>?eB9VD@K&geX(g/S./c7&X
4.PC?,SbFCYKS0/E<5M:W20:0\7YIR^XMKLO\Ld:]U::;b#8(eXe,GLFe?&A;4L5
e=3:;#+>\EGQ@X.AVN,C+,IdY=)]?2=8&)6=D#E#O;2b<VO_0^[#QN;>D7BP02.=
dTHM<616#HH]gKc,dA>)J\G.Z2^IH:I1WRU0)N),B:JWM1\</F^\VBSb?&[?I#8+
E@T5^I+)3f(e9Ug1^SJ0Pb@\:0;f/@C#2U+NW2=3Z\3gW#,9M,6/#UQHfU.L=ag5
->V=6/3+b6#eNfb<10X5A^BLgg18dZ(;)1S5F)aDD]&1B:TS]]-gCcK=J5H4;OMa
I8BA&eO55>_1KFbFY7a95EBPfWRS.(OMTB,UUf<,;HcC)Y2DdV62/;dD=fM<=d[E
&NKC7P)XBELWC6PTHbR-8+FHZPD6)2B>1^_X&E9GEb3-S4H-<]GVA8)fEc=<:M[3
QR.X=fAKI@G6,e\2U(KN5)\EOX/H675.:O#F5(gUeAaL@]a0-BcDP4]+G&/)LMdJ
D.8eD^^_:MGAG<NCY#_1_RcQ4L?2&aMe8N.a7Y@#&#+b=<^><#89gH2RFNQFC:E1
C(U<T#T,9C_b3)RSBK#H7TP,F>[=^6>YM5<WRPLeTTD2WDeJ[JI1D[D06R\84^b3
H&?(KfcSQHWX&&.cb:>fDe>WC&<[L6,U>?Z6SK@J:8_ZM1a^ZIdLQgHC:C<7)BGE
5deg.3@a)DTMC6?H=&;[eJ/U>,7CHTLdKg6PFd,LK\++2-9B[3TK5Cg#=)C:gOXZ
.\A&825@)D&L8&QTWUa[gCc]2KQ)4[\S/@Z0)fSfZC]XE@c[-_VAQKC/R=aRT(c=
7@<&3?a5J@LZ+>QfTWO[58B6?7b9b0K4;0Gf5gA);OUYHL1642^f+1f\0&]bBaX_
H#ecV^I,d<R(c2HH<a1L4W7AHPK.7],+RcJ9PXH1d1&.0WWVS4)N<abbC+YG>9_W
8I?+WX)0Tf]Fa6WgR28@L^B_<1ZGeAgc@DI0&DN7G8W?Y?d72b0M&b2^,F\>V,(]
/BR4XQPVN^S9>NS</Dc;T50,>d<P4>XS-7+HW@8[eC5-GJ5E/IE?^L#WZ4)/:SE?
9^BDXU2RCI79+-C\5))[]-41eK1(;Z\+U5XGO\PM-L5\G6Q1-NRHJ4#XZLO.<SI[
JS<_#D[,A:0;FWf^<J;5BLV:Sc-819)HKb65TNQ9:B1@460g33eefS)G-54BX=f>
-#[GXF=RIWK^+Yg[3CSD3OVf5#MCLX1^2;A:(;UHBJ/-R8H53>/0JIeEB]YW.=c?
\;V;aad4O4;W)C,eKcSB89[CCT_]V-La_THDUQJ8VL6&\-W5X^X=3@,K05fZV=>,
7d+R#EAKX>P#b4/UZ>J[A]MQIWZ:/dK[^QK0_.(^TS9JD-<OK.B0IWC;F#9<O&8O
8HJbQI_abTOPO:P:1D+ad.:1[=H1]OdGD6V99SXU>[P[^/NS5X75Y=(L=Vdg^;X6
eQcaO_]6[ILNaG8@/bK2=W[K<-592<GfDQ4DNXe<-#UY4e--]1>3a7ID#CaM:A:P
d?-++HLe:ECRDC;a1HB^H>]Qc5Hb;_RU)6@?/cCT64;?&:_dFH])^8Qb(1OXP(Sg
K-NfTdeLK+_c84?AYWg>/Q93d&UHD)IOPZg>KXb)A,U0@O#\B&(>9OB^<DCYdCMF
aR,6d#/L_>RW2A72;_4/cTRZ1F=VRQMJLP&Ob(G6C;6.,=W4+H6F6Z\/#c<)X0;0
^=;=d?fD/->(EP/WD/VY+Z-=6[\(FQG(3F#K>^2DOX_6)3J(AS97\_P=d5b#)b[1
g7EA[9c[#0&^I<(Xbc5YUeZa4g3;5B28>I.B]2,LBIXD;fag,JTHg.ag,<8O0B.O
=Y+:GV5Td]#]N):&CQ<1?1FD5NS@(.2A[2ZZ.WWPL.V4])#)3d9EC@L25LXM@WU6
L+fUJO2HSDM[a1e[GF.@YY)+UGA7X;_VZ0]+gaG49?6QL>D><+f.,PM(AJa.[1]?
N8(a+a\Z&9-W@5/bCK]?9-A>.(+XYf;.YA&#=T]H67(+1>G80;K3.]87f=/YZeA>
KYWUF_5E\[YD[eQ@@g-5^H#g=E;+PN81f0BQSffQV[gWJf&TX[]V^/SXcI29;c3C
\d43@G#>HC())Gbde0FPJ2a1N)6af^)ISZ./[UL@Z)a><FLb]TSEgGC;JS;GfcBA
65\3)<f6He6SN;F7QQBVD+eEdH6TVR-9KDd]dZ<FB@M;Z]F79-Q466G8)MKQXH2X
,U]A(Y\&aMX3e-MKa,f.JVN>?XOFBT)5BO@NI^H]O]]CTJNJ9Ca+-Z:-&E-TT>,>
+]9]?M.[Y-W[9_IK3SE?YE:-3DI80S>0V@EdDA)#S?:ISO]0IQ.WGPf+KVG:U1Q]
:6SHBNb&KQE,,@>EKS7LTaKC3ZRdUf).Q8RQHNf)XM)_G^;-_fLS1HT3EL(L8AG#
0AB+6]KL,A6HPQ8QG?9_b^\)LF=gZ.[#Y-TP5=9\?FUO5f:B_17bXBd,97c(L-Zf
3-Rc:^:@VI+790DA=d7./L_WE+:QBa5SX9c,/3d0L<ON2.7-/4NAYc\B^6,B.g(9
,4Rf7bE-6;UIKRS@O:gb78?F=<eQX3gb<;AZTKNI1>0_TeI-J10cDeZQ_4=@0;Y?
VG=/-<.PN-EceL]b2dIWDf,H\ZdbCG5:9LK_<DW8JE\:b3;bZ^K3V+IOWU<+,R^I
EVTdZE)1/cX52SXg=2I7J&O;C)HGWgW;TNUT:X)#T-.2A&_S;,QV,NZR@,Y<@#C<
19PDW6/:S6[7.#Q?+abUe2U)cA(<.ePTAY0FCXeN=ZP0Na&-TYQ^GS)I.;X8=J>c
WR70Fg;VGHLLMPgO&F@dJG,C9\1K1g<M_bFc[T9@-7]eg(SZPS0eaP?,(,KOWXNM
#Sb?cD7YcY5OP6;>G1L.1HVRbQ^4&O)<d44<:.RI7<BO2_5/[AB<+K;(]dN./TF3
=6A4U[G31P@P2B01]SGab=gIYWdb-;H^?RXZ,+)WR-W.MOHQKS+9R-8VXEXgS\F4
CUCV6X]CbX[P2R3.dWc7,e^UGPafTcQ1ge/-)=9Y9S&(9Rd?D=-@PP8-)5gYObCD
G#gX;fg;L)4.?eOM>.K8;Q_O1bN.9VIAVKA(<RLRTC4[V1/CKge=I:e<(Ec3e<.a
.)7-SJ2HFI2QQ4^4<N&\2c2CDdUfZ9aS/S0?d([J(<gaX.5NUI^(G\B[;&BBQB(a
)41L4egL[L.HW0bPX?Y4ZRJ,7+f_]]J=<I<4/#64fXge^LUTQIPM8=)-168]V;gD
O-6H?fH6Q0/E_KI32;@5(])QU.Kg&]I+:B^U6,O\2R;_ZNCBC3W:,5NAc[XM,/-=
+HO[\\^B9Fa/<I\Bg__XW,=eUe8?L?4JPfNf^P8M:SJA8XO;LeG..),TBK./P8WI
/dI>+BFYU\J#NbFT3-)5?(\@)>U)gS\CT./X_BP(IgN^FS#d8b;V.#ACY9-O/+TM
OT5Q5HSG4P184>M@WSYKAZ=decA]E+086>e5Y)GcZ1^@ff0Y9X,\Fg@)/8/e-gMB
-6)_]CSe#^&<)#VDcLQd\F&ea96SX1]9OX,H=5MT_:S]#P3K8;I_JFBgX2a\#S18
49M:b^]Y495<\Cc#@3d8<.&9Y+B1&(LUc_?#<HF>cCT,0KM)K]AP)>=5WHO/#CAT
HO)[-HJ_d49I\fKXJ\D;>80LUXA8F?@(XBV04SX0a+@Y@;8Q^YA24d-agW1FPTL;
G/:+/R]6O9@EV\+J^c#FJUXP6;L9^^D.TW\9O,cLW:^VbC3U._)5cV/ZHSCQ+X-S
T&4?)L0MH+&a05\FgRBC1fb.T[I:,#XU1?8Y9;4,SB^aYPH:;Q_)<5g9Wb\=1,Ng
+fg)N>M\5Lg2(K;#+\UH&]Y6FV2C_[H)c)T^e\KU4EOc&GF;M0,J-IY&A<YRHKbC
BW_[R(3&^^&.9X)aDT;:@8HF#SM8NHK]:T.?8fA,GHLO<2,1/WEK\C&4+\FNE,eQ
L584G_Mb;#9cU9X[Q&20H7K7MS41-1?<c7.=Kde_DfC_I<E#>GZA5=N=KY)3b0F[
X;g[(>N>/V.BENZdXO),JTTfG9IYc:;V6a_B92UID96KUV^8K#^P;C1^YMA-,.@B
J/:B9YMJN1B6ULb8+?1,_/dWH0]#a&<?b?Z48eTN0e4WJaPM^+,/^Z[d2H,RQ(&3
)2g[7dX9/C5E+.T(.#E2G63TXeC]d@XU,6ICTZI-Cbf<#C0L?/T90bAM+])GO^KF
P455YfPE]WCW:,_<_I;&2QC/d+a[;E@RFcR@NAUA@5)IU3J.[GJ2-=8c\G.,70KQ
LLBcP=IV/D4G8/W[KAZPR<1NV8Z:IZ<&;8T+7VW@2WRI5Ie_N21]4cHZ;e4S\ZJX
40)U@\WKMIg_[g2XP&=PV_N;C\K]+W5beE1;MAFR=>D(C-K4EA\UH#TRcOGAFdPb
>V/0gS&<)8KO<6?XR93fb@LS7^g4/#&gSBgI;U@;TPH,00DGRDT[GdX=R9)_@HA7
&P4:aG=;T&#/T];\KfUcS7=+X6==Z7f->VDRKG^2BD(<[5U(7e\YZ</CO2,[ce?/
P<JKec]T-C+,62J=Y>S-Z&\b<<UdVc?<FQ#-+J8^:4AGR\&KUfZ(LK5S4VA[R)3.
Z,WR7@f@?B<^>\g\a+O0(AYI6)a5Bb\Q-E^V1?^b3YIeF,ZC6C<(b^#6Eg:4f06g
/-c4E\:J-RH1WZ[f7XT5>?@I]2,0855P9UN1F):[c@MeXS/ed;I_((RDCec=#OUd
5d8E4WX]14XUaUd@75R>X])QNS7&dO:ZN8BW:D)gK]N\TUdf,D2+6_33)/7]g<S;
&b;1J2TX1&X/]+Q+SX4N>NYM)d-/B]<PcAB_:MNZ_R=AJZG3ZW+02?<#I_TcbKKE
^J)PP/&Vc9WWS2LX&;:dCfLL9^+ge1:5VN-]>d_SEd_M0,c_G<T<91_b3-.?QM6e
J6BgG^J6N,[O7,b36S&R.GUO.&M2<(NGRU2T:[[FYIQ+K&LXX0IW7LZd6:-)<>4\
_f]:PKUZ=.L+J;,T)R3DAYeF-.3RPJ<f.b>RT97Y)YKM.._4QNZ3_b43ggaZPDEQ
9WF-#R)LE=E:9H-);@?R:W(eLI9b\4,KV\@/Sf7<SJ0&cVR-eaEJ)1g81:I4b8SU
2:3>?6/,(MW@a4Y.#fb+40I@RZ)O56R[[(g^.bU[]8,0(+aU3Jfb.79W1.P@.4I/
?EJ7dZZ>2]XQ&7<>5+#eM>,I.6#S?G+XZ)-_TZe+(L@@Q(.U>AA2MYF7RcS:NB@J
0V^:6)L&RWL>W[71BKSS</QDIV5-.@Z/O;N@CU#5&/B4.:MT+LO6]fDPcb+V@daD
=EJ>;2HLL(O4cI77?[<LfE8X,<;?)-[@81c_4e/86?/K;8)FL>DE+&M)GNba=FF>
DXf02.,QDDW1^JKN5MRZ>BRdM)CeW4EE=L(AJSGM0D[>P,3O4K[5@eBAR1R./8VP
7d:NBA.53I_bK.c5P[_FHYW4D^0e6E>\I.D5AJ+>@WZ&F4:)K/>YbMS7f0Nf3+O/
SMdJ<8NE<-=0e=bY5QTKc)]fe[YdaK#IJ)=X1:];VOV^T_.H4+U3[_+EdJOIE:e,
?5]@CUCWaGF.a7MS_eC#1;&+H&^QSWd7.H4.CQTX.S?N^Eag1[IgEd9JcS2Y,Z93
:.(VI&\cI+?NWeA?&6NU@7(6#:Y3_RY]+@5[&B+E2>MbCeCM\VaSTM9>-<P[fMNc
]ScaM[B7@QJ?A^;FIP^eY<8f7<FIA/g=<eR#A(K,BM]N:YBP8O<;^@53,L#C6:H^
1YJg\ETZUZL&]]#HN]U1G;<8E<:^7@V9#](66H;+#MMA#1<A&6DZH8=c+IL0(eLS
32gH?+7_/1PbfYFH6fU88;JGU0AG=<II]:SS#Cf2?QW+O@F6B5HWL)N<YMd0GWd=
.DH_2K1;F0b]W14Y\K2A)I94P)<:EB8C^cc]9=;9L9BaF>g1X?g]\eHQAO#G;4+0
eX=Cf:\UcY@aXVJfKF?7>bHU7GOX;&cQRXg;bZ+T1AT=VBIG&+VZ+Oa]B/O(>9bL
AVY57J;AA\AO\;aD[\T10V7a,W&M^EN8Z]SV#@2(.dIfSTa0(&.N^=_R0FCMXgX=
ES40eHB:\]J6M4SWFdd8Hb8AFbJ_?YbeG7cX/-)7eTSW:5+@_Y@8_9IVG7S#</P/
L9V:7K)\(ID70V)T:_9&WKb^OdF\a++F1^=S^+bIUY66/d)@bUK+W[I&;.O:-dO1
Z&RDPZ)=aD@ad=MBM]UaS0N-J#E,=:(NTeO@=YfB+;4B&WM<UNHKL>e(1d34.)Cc
W)9N=,2RF7O5^PR9P_HVU?SS5E&&c?EF/:G:3>M,/@E5-Lbd._D[bWXUO[c4>UQU
@P4e^E\d3d7Bc[NAG?6B2J>M:f>Qb8K\0eDLa6Bc:U/)RFM7B.S\K8PZaOAB,gfM
+>/J4gPKN0Y.(G?=2EOf:H]D86-KH7AbP5g6ZB>;DcN^O,5]A-N;8e@c^1c62Z@:
?;_4e4;QLTZ8#&aV1f2Q0[_)H01RN67c=-cFZ.L0)fCQ;HSHS=C;OJSN8:@>XIcB
H3M,.WGP^HL]dY-b(E3U?4WSabTKM<EZ=&3UV3)A9.4R\ST[YeT[@Ug0b;CYT6)I
.J=1#/9\1_bJD2W<9JEY+M.@W16:Hb@c=3&E]:VXI5:G92MJ/JF_=Hc?/HUE91R)
^,IS7H/+PfdAag=7;+0KJT.1X0J>;,0_:I@-3K,Gf+ZJHRa/@-^03L9Q3H+CLcV,
E@^/+N^IC7Zd](K4g:-be3>2:-P&0g6L.8RYJ9BVfTXb/4cW/U8E90>=,/8PUZ8U
eT7Z3ffEHR>/BPc\[gR1CTLR84Y/8e;GW1/9b?/V:#[PUWO@3MEB)#CaQVZCV?]S
CG<a^GTDg7EgVdGMU\d4M-B)3;e@KdS1AW,Cc,4Wa?OeB)XMHY&[gC4PHD5MM\/5
OP_2^(3Z26deCCc]A[H1@EXdAdNL<D,9,#gLBfN-+]OYe@Q3\(gA@W@4Ne)[-YC8
RKYAbS&dNHPbcZHE0<VT?BCH9,#08f@<R<414E[XX>7LFM<Wc\K@H+>0^S_L)Z0]
fgHMW3RME5O34M.3/\ZJ9LbT&P5Qe<Y5]:#,<[1.Ufg\]37:OT3O,#CI1g#RHD_)
f0[4_=-ScbIR210L(457BV_W=RA5]fYCW<=X&TRYdZK4M;D9N/??dcc7\?L=&:YX
#ec7J9[#5ZgN:<KWDf^bZUD:_a/eEMK[A8A&_:<YW?<0[BdOY79a_2A)JG=\SF&d
\;6V(:aBQ)b#9feH1+#[La.HX8NRFc(bRUZW\LD>cZ?;PdN\X[=c@ZOeILgbKU98
)RR2@a;JLAFbG#<+0H3bM#PS9:_Q9fScENJKG=Q6:0cg>;a6fUGSV?D+0&KZ7I6L
N393K/g<>SfK50[/0\QT-a(g+ATR(BfY@/cYO53P57132aT)a_;+[bIV<N=NFKc6
LCSa6.X,58H_]bZ.NLX=_g^=5cBV9e:GAO9B;&1a_VG<_.Nfe:F36b:fACZ6#43(
c+&.>X2DMC7O2MD3NN;H1)UU:F\Eb@)38/=Mc,U@9],a;,<GA0b-eO3KTg3Kg+&b
TK\.[\2Y42JD+&/KZb:2^W[HOO95+AM+?MV+MIJ+P)R7g#e(74Lb7=7f@,]4GcF-
?5VS]HOY^_/BXCFCSN3gR,XA@TR20_,e,WdKLg&a1^GYYdSSB/U_=UZ#SR1D#XK+
aY<]GT/c]318Hff5X/).&XT_R[<f,P88(&CM[5PLfJVQ[J4Q:eG(=]OcC#)IK1^,
I-E9<^9d--?C:DcVZRC7A+RG45G\SZ,<g0[6(1PY]O;/g>-)+bLLSB9e9dN#Tec[
BZXT4g>83ADM?#Y9;C=6GSV<ZX/3T4T8g+U69bYQ#E4#YX/&Z)OTc6O4WHQa9a<f
+.3TZ4P.&:6LfQIcB[K^gVQ[&#gPK(C^@TBdJ,70&G_?5SRT>f9K0A0]O>BaT>g.
dR7Y1GYg\N<J?]?_f3N_.E/CI9,caBa+B2N@baCZ+[EXE13edE]GI89.+eA&09?Y
,.]a/3Dcb\N?HOW?L]3Y5_T]a5SgD^GRD]M#6?KMMTLS>P,RH70VE;Q1XCT@\K9+
aW#842dJ[,T69+)GK\N=#=#BF3CA_IYQR=V@,6NM/B@AA^@KJ/aWVIeW3Cf)06,P
6:87NT2TE=,#AP>T-NH(K.K]gb]PL7_A85IR(SaQg++W[^M#SPf)::G6Dg9,HV^V
g1@:?+;1?ace;:M>5@;7HR5CLQ/JCb3?RAa85g5:4:/WC7/0cEM_B&.6V_P>,9,\
@G,6X?GT3,D^YdeAZ#2KPUc<LU:?_<b7:N[O8F#D+-bOJbg;c\RRR#c:&+Z/KVC:
Q3WJK2F-f7\INW_MLaN9YQCJ@e.FVB)CF)P/?PS@d:+I.RJ:PBUV^P3EL;c&/@2M
F0KX.>P\?>@g5TC\ESZG)CQIb5Ne-ZY\A_CfBN.2Q<36c(eWWfa@F03NO(RMB<I6
EIX[+X<fM0M>74Jg;K-]7DL-IBW<=SQW6DDc0-R\990I_TA:38d^^,JK]fQUOUSZ
]E</UTU30)?N\(&]0235Abb=P0)V&=P?(4=cGJV^.URLY;_AfIFU8T;Q5&3M;KHb
GTb##R-CN+U4e<TcGOPJXKI?V.CD0\X]ASEf5cS;4dg2XQTC>2H./a:OGeF;<\LK
:Z&bT5[#41,#V3&EaO_f,Z0NC0AfDT9>8MQVDH]2UUD]4,40f6NE#KY#GJ77Y3d1
1)<;HeH,PK8YDMR^cgZH\/T:d,CZDNY6I?XRa&dc#YGUD\Y6eNB36BSI67^:E9EA
W-fb](c8SI./?cD3A]abAFa]U8>#R7EZc)K30Ve5e^=;>LcG8\N+bdf/<8Gb^g/Y
Y9+:;f^6:Q49cN>bLFS\BFLWXR@f7\PU^A@4g(V(XK)-Q&Y+(KKE89d>.>I59Yd+
1V(_C+WKM3GZVK<a6)\U@L)df]E6ME@/=HG6J^#I9VYC0GHTS_7;\)24Qe_&e3,7
I?PB@c&NB5c6ed_b(O)c_.)80PA?QW4eBQ4d7E>1Y+gR/:<S_b[\BEO+^0FVQTBX
Xd\c^Bg1EQ?#&d:?Y1/9(9_^SK=_06bVRR7aKKNb>1.1VT\FFY.Lc@>SdE44BGT-
d.@8bGCH;NXJ,.)(a<&+RXW3:/A.B^\f?N]3_\(BZ0?(0f)BK1A?f^K(Q]_]5Y.E
K_G-OWK5C.^:D0UXBKO\Z]dY8cX95Y;WTAa??<&E[dgHB:gPLX?J>)&@aJ_d1X+2
Q6b5/6cR<PGP72A0ZX#B-589K3]J(,&@L[e:]4g)I4I\CRFV+LCY&1G\7D_,?IJ)
S/aS8O&TO>.BMXO@5]-K0N7;eWb@SM)_7Y2O?b/DN=29e\N?c48,3_=)6PJY,Tf\
B;^6[:6?JHJDG_-d+-&NMLA/2O#(]-<4)0?SLGa5L\@+KN]38gOfPOMYa[NY6)FE
Vf^Hf>QU@H6cKd)B\HSQ62aM1aVad-5_P\VOIJ+6W,5OcFT3/2b#f:O;#&8)+Z//
dLEU_E,g(e]@C,?T[D:K#PL_LK2<fSAOf:F.,;672ED51_:=I_)9XAd6V2-f=_MJ
c;A?@(.JY7\3\12)WNTdRQ9;6#L=6]DH^ef\5U[_&OR^=)SgbQ/2&HERFTJG2&#7
dO#E#O7D/F]H>eEb2H0=N7aL^<L4e>QQI38:5feXR,[;..b=QVN&6<S<3HC\7P(5
eSAE+&+I/gdGe=gPMeGB3c,2=g7KNZT1bHQ:9XGMf(C-=>Rd3;I.()30c]U+]MR^
^0RVWddQGTWM;DB^/(@JZ+M>^/fHRF8DX;]NI7S.AY&</Q<LR07/ATc(:Q]YR;G^
.BbT\0&#7DY3_W5e1ZJ<V\R=\@VIR35VY)\S@Of7C1S:0KW=BL67Ve1:P+DZ0e3B
/AK5c5<RMT/-a6abag)WE7P2?H<Z[7#SeNQT(1bE6?\,NAF>:3Q^.UL8GLP]BT?P
,2GIW#1bB/dK8Jf4(JRO;FFe?A1H>\c-,0B7AH8geWXZX3@?4X@J[1Q.Pa)4:EdR
V^[--bA>G_;DIgJ-N.FR\Y6E9^)^T=GL<8OFTFTWfTd?+d0=\N^,S^Ub(<Z:@4d:
cb)6f/W>AABCD2YUPCHH@CW1eG6I[-M0(@F(LL,2[BZSX\Hg<=)-NeMdb>8+0B-G
b<Qdb[[dFIFZQQ)58RC;6SdEAc/]S41L\BG&AZ1?&/Zc=.Z4+EcM]67F-M;d.#X(
=G0GJ[WG<3&U@CbXD>GPNIa6U.1HW0WXT+L+Aa6\baF3F3CB5U?KeL(/c+a5gUgQ
0ELR9JF3W.^N]eS9G<IOIAeg5)fF)ga=:&^Y7[6\UOORB&R>53&UY5=V02_)cbQ0
+X_E<KJ#OF&,^@AUH<cS<,;MJK/8)_DZSE_ccQPL=4RKgMH+@NabB4a7P9TFKQ0C
CZF4YJ^ZC&NI44G.05I3ge>;VMRHZ@Rg:a06Ue9Q8>_aVE&dTO]ZW2=Y@Y:3Y26d
OgaKFO[6e^Q1L#&f&aZ418E4@5AP<c&VBD7SO(&c:4T&U3+S1&PB?X?;bZC?c[O&
7?XK6g0,M/&L.B^C^.@E>GJOA97&QKR+N&faL8/@)P8ef=KLd3>+<G90RTO4]3f\
#_/1T]UH3@Jd=DDI&37:JR2QW:R.2^_TdS4;c<U_(FLW7WWN-GD7QIKO-P3:=GXB
Bg@A(U[O5(5=.LHLb#3DHNC:eF@,XOO6/b<Z.E/V[GR^>O)ggVHO#9NAedW9>C6I
S]X5_7H^c[[)_ZD(F<S/:Gb+XF5[:5g;,SD\W3&OV)KF#9;M=)gM(Ib\c3A?URYV
Ud_:BLQ>O#/B3Y91DgL.4PGbaP769=J&fG8^3;d\#-S02OQ8LNM6dUN@8S@50OQ=
A0-L.>R4eVR,B/MS&N:;O4P?3#,/:GL0Zd@PRQNT30R+::c?]?DF,.SY:]a9P-?8
HBFUK_a0_,4KaSQB)7POSb_CJ-d1WDOQ2G0c052&=^?W0FN;P8d4FKeWXaNKDPPM
-8+d]QaYUfe,dgVgE5H76UEBId=2JJGc7,3^=,d4,J#)2;>7O#(L->8Y@.e=:0DI
^<?2)e+E5+VJ/LX?WX7<>fX?R6[ZBP3.LBa09(eS19gLJZRga:TA/[^JS9LU\1\/
b;1YSGW7Bf#Z,IS+:.6\FD:+NVA6TAH4O0]g[DD_ReE)e7ZDTDTSbH\>ZL?&RF#N
1-Y]:M0M>YBH#8^[bT6F?8/ea,gZe?A+#:S@3NeCFTFgeQ-OA5PZ_-2&-&ADCKEL
.>4LXSN186T#Dd6XbG2YL-AW9c\IV-:WBX8V/03&:3bOHZLNGDKSM;f^J6=RX_V&
B7+\8GZ_U(QUN,.TUQ2ZK44()4;6YW^eT^1:@UEL50ME;>I))U>G5^/V<LNZHIcQ
QC2OU((W4X>U<_MV<e/b.W6_S4BAe<G:+ZB;@Q[.e8;ZN&;caYe;E36VCe5;bGRY
X-:CXCIP:FOF/,7@NP=FZWOb(cWeDV.J#>80d69X-,bgbG/PLg1@RV/8LdG5WbY&
ME<^;[.H10D?c7ff@MQ59A408P/82)fD9NJ5P3@4&ACJdSFfI(:VS<@R[ZaS)&_D
J-FgeM#:bQ>T8.cU&8HH[8F.0N4D1.^,eFP>eS+Naa4,&((&/[0,&OAU9E8:D=ca
HKJb.4>#a4J@6g#O^H[^;H><X-I=[0,)XRPb5KaT-Q)dbBg#4f4JX):\I:a7b7.Y
XRM^fE_2,B29.9bb?GN[XL-H-LD+(a1I=IBP5:.3E5W^TJC#3LG1+4_(5MF;5NOL
G93ZHb6K2.@VRe47gCZ=gc#2C8a#c@><d-ZY\eWUD.=YQg<CFEC^_.Waa/5RYG-G
4D0?F7GIT+?aS3aedW[7fHWH^57#H8M;-bR:2V-5/:/.e(ab/Qa4:<ULdF+eR>Lf
I2\1(9PAFce;_eLC)0B,O,d-SWgH6:4:ZVBZ.O6cDGYX.H-EEQ(U]DKOb3c\YG9]
VQ\RZ[&BF;[PS=HfWDXAMc+<9D5J0:=BR<OD?Z#R^5.FT7Oga?8_(-=.LeK)3O=;
@P:-LF?S(^N)C08/YV-VEAKD9#AJ8NJ)I[B[USO@4TWg;55]e&#/L@Z@&2YPV4KL
A0f(#30bf@I8K,6#0e8(6J7-QI@CRY-_7\(#b<N](J7J_4fa=3H:OMfHcg3N4#LD
aa6d2V8+PV+cFR5?Y5X0C504TU(&C,6VDeAN#I<\)QZg8[+D83e6->K([4[-a0D\
=@Z:2dfe<9U3M+DCP&P#Lf,HSZaFe9?-fYb5?ec^J5A3BG3AX>)a;X2N749(=WAb
;7^=HWENLM7d<4aUb_?3DWBZ5ML&8)4ZL+bIU8dS6-9]4Q@5?+,eV=XQ=9-PPa0\
HgZD?2/69P-/YUG@O1=:/RF384/Q<L4KS&QRRC,>K=X)WOX&>HV[a2Mf+REaG7SQ
RVI[OWE_e<eAe=D_Z244[=RF)bV^6M/R#L?[C(<ebM1Ac1.O/F<aM8,UJIgWJG.2
LWPA-BK2DSID#X10L&Vc3VIA#aJM5(ZP_90OCN3Zd1SQ)e:H(BRd^dYdP:?.^]Q5
ZGVea+QgJU5ZL3V?B<YC:657SO=6\A:PA\b8LI>ZQEf@:KU(f(d/,SJQ1,f\[4\9
S\_\OFR1Z,/-:_OBdOV7GFg_6.37V/B0AbKT4N/;,ebREfWd7)G(\f60fbLTB7.X
E7=T1WXAf&48,=CAf/2^L9@&:(:T8U4&KA2RZ^Q4PgJe=(aI420Q7_M^+7#7GYO-
-A?.5&2a8OYG],QfMc#a\>^0<VIENZf3I,ReTJ&/&0f1M@3+,6&1\+=8VR5Aa-L3
M]UfJH8@(FMNHI_]9[f0>d8Zc+PD_ZPIJTH5E+/gLbS__B1/(;75/FFcALIaTZQG
\<Q.PZ;[Z&G?&+V)G:X_TNE1.X)@fKP5TX=I6RN<c3CJ>7IWdZ[@e=\]gW[fK#=g
?ga?,8HVQJd3_MF&)Z;(@ec3?4Y4FIIaF_>/EN-d;6KS1dQ77L@g8&-VI()MXDYN
32YR/-MCbd[f&9\.[dV?BG3X8c)MHc#],f:;&a_\WJ0Ic9c+T6c&<)^_d(\CQ.]C
/^(L12?SMdU0g1Z[Z2BfDE91[L?VZe=Rf@Q/WT94WOK+WC<^V(<DRY.e;]NA]_\g
#Yea-CNG\VKQ-SGe6,RT94(1Zf1]/S7WV3_2&?=L(7Mc<UFc<3]GC;02R/5<bA7C
(,H6)\C+aV&I5TL_E;UCI&\G6Z)KXK[L10O6dI20LO?U&3ePc;eY<d6SYSY7\D03
.<\4cAWaN_VFE/^d5(>,XY.c>[><?N-&4b;.W>6]3?GeS&:gE=TDVXWF8V7I10T1
DR&;Ef,^^H0=0(OV9V0?:LY_g/]G0KdV\JeLAa1dL261]GZ^?0TPe1MPOf,ffIV;
cRR3V[,W21:4fK2FQEac(-(?YE+S-[e_.?&X7aH^Z9caWA=@;GHM-N\BW50PK^F4
P#&5H9PJ2P]eS/D+7ZgH84ZVI)U]@:MH,E9T?.M:3CX\0VL=dag0AV2_a6:7Dc\R
ea0.\GTI<KLNVL63]^UOLYAW5gaQG,R65\V6/X<#66adGIf@)M&aX#P3_SJ<[>HO
9-Za645JWN21BbMYUV-M8P;dHV&K106fP]cS<g8c_;(\C&F#76<QGPX#E<EKFL>B
,K4]aS+]J3ZYXXH(P:&1+T58)5S7=EFODJN>1Z4cWFEK,MGdB^.ZQ8)5gM1bfQ??
L2Q2S2U;F2<2I#;V,[I;P&^4T&XKV1a;004be26g=T13:M#9Y[d<Hb:8K+&?Dag;
>#6BL)>M3EU@UF<gU:\NZ)+=CUc\VUb4X?3gK+^gA9O@aEOc(-;BU[4[1:;eU/\)
E.C@?SBf9WI1C.dG(/BQ8B_QRCFE4D<@b<&#;CF-(UaY4:E_^ZJU<?B;D+J;3>-B
=K_HNT.TRc6NM^SHVQUB@<c\bI8cR5OadfSL\;)EQ>]?4\&af<@g_f6a-UT<9;:O
KQ((.EL3=A:\_C2N_1=9+6A^;eMJ#SSa)JRBHXYM>^4-L[H_dP;=g12ffX6SXDEf
-LV?.Q/V,M:ZKI4Tg6JLVE4/L&46IQJ:.H(<AJ1eUbg,+7DB?/B@8HLC.\UWHa[[
,EV)T\G#BFb?J_QS83e3\^A2\d#OeR^J&/[Y5fSQ3ZI:H6V7J0UCFZ99_fK_Q2/:
GcFCg6=+1.1d&EfcX4/BSbU>\@J;41D2R]#K<9>:D--2gW5BC3G)C\/L3gb+SLU9
B9@6_N2)aP_BRWdC9A_aMP9<^[]SVP/A3\^TcZ+EDQ=XaI5>YMeXfWMLG6]2A9KB
,0.,7/7g1I,KD]@P<>RB:Rda?PBc1WLbFb&796dC/BZE+f:FXeJf:(O(9NGIP]EE
Rc]U0=@@F,H<R(-1MBbZH-a(=Y7g>GY3FV.X)2>#(LS)Se0cY&]FCGO1?D-]_V0)
/:6^=1bQ[,K@VOY4QD?eLX=I//&Y,V)2IdeFV/;ScK?3&Sg.[@[,:V_e^HRA0b,>
FOT_R\/0D(GMMS@\F[M\7,H,EVN_2e?,T)c&&<07++#47N:7G-E=:#KF65b?92,M
caW(C14\GTP.]/7#OE1RZU5F_3J9G7ZHJ01_<6NT=5#-f1gZLAS_3B?+dIQ;Jb/P
94SRX5<MXEB8gXR<\E-<:AXQ&=8+.>S]@G3<.RC2badfE7AO(D048-84IU-8bF&D
T_=cc2ZQR08f4JLU,;I1003Gee@b=C,(O+ZO(36/0e4/,B^L+&@c>[b/9?>4egVU
;..+BFdU4=BL@=RGKfL_&.W+f_=?I?0e#H23R598\.0_3.]B6dZ>]@<ZFbSWXU2d
#-E+5Vc+1U==HLDg2\\_V,8(]c2QE/5P^:]d+43RRKCP\?4OK??T;fSBe&c7[+;d
\V;8O\-0HE58@Ke5BTH6?/;QaW04bc9A7a8N\)>c+N_d\CbaX5G&X-bcdE<==WBg
<7LSC.G\0(NC75d_M+A+N7KP59f.?9V\;BBU.W#[H2Uf7L[J;_6Q+LeUfC6WdL8.
XedI1F3f8.V1RYb[79:G8<&bI)S7O7><VX<\G^Kf5OfQa(K1O<:&dc4E]8&#X&WN
&D(LPV;(V2H(T/@E>_7JP7\J;X:#/P[@Lc8P3Ef1/GUNbZ12YK/+T/\K6PI0]\EZ
##b<V^)I&49,.9.GH3,3G18<TK(b/9K\e&aP=9QH5];[2EIXLMOAf;V_U@\-e,a@
B[H6f\C(AF2-WH76,dfPC&a9Cg;MG(R:A+^53N2GEOccLI,c^(VNaMa7W21@->CA
C-F+8c\aWUXfe\KS/@\6U]]_0@<OCH9_P5=Bc/#D9=MgX(WF:#<MNWH(7QOV8IRX
B9(6]GOL])WdSUH4MC-8R>92D\.NHdD9)1.YN^)?=F/FM&V2C&6=gRZEE@eLgB\B
L3YGbSe^B^MO/6L5=.cYDd]R=8ec=dA,[:GT-8LX@18XJ?V2?/5T\)FNGg3_4TQO
84I7@1RCGcB2&f#HU@R,0N>LJM(XTTc1QZggY8G2c?46c,50YR1=\RR=c#YA#A4J
E07_g=B=d2PX\1J^&5V#Fg50ZPa7FLC[0RTBTL\(M.MLc+R3Y1;6:gDd31=J>2NO
aSH2AV_[_(NUPSS#1YFOW\>LH[OE]B,gMW0+_ab/X[UB#R#IK5Y\gaTNBgS9-:+c
/#>X1J<gYF?fR@P)(MJCJ.c^GU57@347/OL[.<U6V)N139VGIRN2SED_bXH#\MAS
VU;Z0NN8__K<^TJ4PF,2Ufc((@2Y@7.6Q:C>;,O#e3W5@VF:)[@5cK)9Ff(YaWgK
4,I-Z??3L?.7414D/J?.,TL./.EU38K+:d3fKc,\J?6R4g2PD9gK3HS83c0KZGTg
Ta)ES?NG=R9J=cNXG3RL;d7V8fdO[ZZG5cAd.e(>L0:)ME-Y>-JPXR]^+6H0R#/f
QBZ-<P=OVF1LD_bK8[)F+7X?=--&fXeRI.A;__6\d8G#DR0e7,W&F@Qaf5I=]4)#
1P^_-?4L))-1c&c5JNd58;CI:RP#5;]G3^Ra9&26#9O_JG2f?WO-9BLH/[1)C>2:
PJAfFZAFHfb6=SL.LZa\/^(aNMAR[TaOKE.XRYbcbd9>>c2RH&#Nabbd)KUXFX01
Q\f#L/Z)IDBDDJd?)U71+6A<5DG<\3g9I+YN)I,.VTS;Ee71XA0b[d:BGUYZK.DJ
=?6Q^C32#aT[>PEcJ83)eVE7\dJJ>+_.P=\MK-</&P[,.^+fab&V39M1)-,&ALLa
4MXHVS\6g0++-Cg^4A#e68I5MV<K5ND74/_ZdIVRa3VDTF4eYHcfX]ae8b,GOWd,
X:_R0&gS>G3/<e#TS8<3@g.0GE5fY,XgY,UE><R#g<_63fdC[=)7cB_QJ\HHZSWS
[c:>78K\SN2IK5c4C(IV.f-^>08J&&@X^a>6;4[:P^)NO@CL_FeP5).N@TSWggC#
=P:e_cPSEd,J)Q1YM/5962gE3WGd+Ze#IQOTYB>?3Z)HVaf[=CVCCT48N(T95I3.
<J;3a+gR68.X)e335(19UEc?(99+FID+3T#/(ISB1ZZdY[Ja0+P7/F)5INZ5,)#+
NC<8-2\H?E9^7.@KM@XL4;2)7:/_&JIW;?AG6=8c#XJN;dbHZCP0a9\_/S1TI2(d
dP?+PSQGB&JSNg:Ba60V/LJ@4CMJ4/<O;SL76K3Le7Z451D+FYc[17HQ-O.\F8;N
.FI.#LR/:bH]WGY4NR]76HVaV.Wf+VIe5b;[X4cMI94=IN/6+L[F/+.1ZFU#>><E
G3_/ZE,0=:/4dXe;AA&RND_Y.6R8\UC[d6]9S:Y+HP:bG=A@1eLeN80[Of9;GC5X
3DVS85(EBABCH<ae1Fgg#D1\dNGS18CZX<L5.c5O+7C>=DbZI]8JKQ\=agI37F0^
MI[[MSDP94B2EIR62.Dc6).@^U8GE1]GQR(,)eXD71aS@L?2.CC5eV@#LZ\V&GC.
Yd&.,.]E&?H83KXaK0NUUZCY).W5,AB=;6_b7g,@6dZI4_I;Q=4-EdZC?Q,>FIf5
\_O^cR2=2^,eDa6/Of/f5RJD9a[=EEBd+dI64Qc1g>NPKG24(63OGH^;C?#:e?Qa
GfeFO&ZZ_&OQ-+d^_Cb0E3\03.2\R#(Qcg-2:<7^AaKA\\:Q.D+R&23#7?O@I\P^
f&eLeAD@,/8[.4YD_d.+8UZAZNe3Te2#4)-b.>HHbC6(QJ\_cVI7A6(YVOMBS:5,
WOHH[T9ZJ\@b80);B?3U1MZRAA>[f(=EV4X4f8YDSd5GB-B#4G?fS;:A=0>A^W9B
Acd,YPUa_F/1B([7KQBZ2H<MS[\&IO8^9E?TZS1A[KKMJDV#1ADJEAZg==V,-/@H
Oc#(6ULA\1+>/PC)OZRN\Mb)\^3@QTSJ+464WA0I))OA^X(?00+E_BeALWBFL,,K
D+@8ZUVK<e_(4]M6S(6V;P]+98M7[(c?0;Y--&O2H6->05=6IL25?(W)Z#YZX.).
ZP>.bX2SgM62JJL&XOXe7;EM_Oc4+]d,HXV)X#9+RL)Ic)958DC>AWFBK/a86b5P
0^/,NT/Pc/V0P,DXS7XYZc:R+X+;6eCb8IXBRX<[6Qa/F5JC+,4:TM_;5c[XM7^Q
ga&T9?0^;e-#FLfJHNIFgBOTb^=;X[E,6WM<?[a>F^(+AFTc2KM/WL5_UK(-&Q/>
3=bV-@D6_[N;&Z[>J<TPE+=RZ>IC2J8XRA_f88J#:b^g=87@PdPZFAI4QWD9GeU:
PM1AIRf/X5D?+H+<g5O5>44f(<<C39IU/[HVc_dAT^[W9&0/:9&//?=955R4JG^<
F49#]6I3F)EAZ,M,MV:((Fec;URW5TD)Qf+P=&>=bT\>[;He5Y-b.I&?JK+154X_
?\4c[5L12WB5SNTL#CP?c]LZY8Mb=Z9S1]3LICgH(SH:6KENZ,D:SRKGQ,_b2?@1
E53LX25HTg,H)WaW[5fbU?bfE7I4]JLD@\P4.<[8D>cHbeWHVC0>32BY0]=bNC\>
gd1^L#S#EcB3?YWSTVbF.&>E90T)6H.a2DQ1WGHVY7<@^J7\D#9[?.)Y1/6<V+-S
>3Xg,G3g8LeT7c6-B+5QF6I;LV0c)06MU,-5eL8Nf(XE0ISCXB#JLeYZB.)cOfLH
>f(c1d&CEMdXIAW.cdY\YPE:5)<=&M,:8Hg=3Ngf90c]UVU?G1+R-BELU()344J2
BT0RMb:=)XGcFBG+@;e]3+RC)XLIA@J<Jc50+<\><U#L@BaOQ,Z5)a4MRC<+>JSd
f3KR(5884,HYV8P>@]8W:FGV30c,+Z/=@)[(9M.[aVV^HcLE0XgB3GG\)F_\)U&L
=55RaBAYR3/PbR?:(Y/CU4aH4aCRcQ4,aUK=PRQU/Q-f#,B]7TC2@,-,]+C_<E?J
8b&F5LU70?4@X[<T]LBO.5[E?aAc[WUO=>79O2,.8Vf=dVIZU:&.G7R\HgU7fBO>
;<9Q?8:C\g,bMc]-)_6QYAAED+CaM07Ea./33)8XE9(:Q=gPB1](YZW7a9PA.6>(
H:-19G<2<3U,:a@6UdDEc]]BAK_P;P5YaW;X[?YeU0e1d-/=EX5)S=:e6WFV.#dM
3f<)L=>0=1^UX0d)>DcT(\([2CW&P7P/B]TZ__FC#Z>,3cQD1JB;e_L_&>&]WW.9
)DQK3^&\cP:e^\8HVH/6<+Fd_M]Wb>#J0(<D#_;ccNOP+&=d<ZCZGU9NeNE)F=IP
6S=W@Sb7KN+BV>K\ZNVUSM/V7fK&TZ]7Z>b+^42bLd1:7P<DM5=)/_):V#7VH0O@
I@SL(9P5beVMM,J\-PaTY?18:6XVS:WJ2,@#gaOPDCa=0cVAfg(Ig0[A##XM7V+C
0a([79e<T<E2.F=Qf;5.[ARC4JE(#8(Z=+0_JYASG,.Q=9VS0,bX-E5@E3HBbFR>
-];S](;5#;0I+Pc4PJX+S)_)fI545bNa(Sb8UU<[OVTR.^UU_g\\E)^K9CKM0d-,
)2_bH9]^B[(aUL?&/(Q\LD=1:1(23f8;TAN+99-G^4;@3MQR>?(aN?2Ua=:GJ_^S
8ZM>NO(U9RVCZc4Vgf4fY]F(c1LZHe37?G)WV\5Y5F1LODAOP41U6Q_..,e(J>-d
7R,5#cQ+M9ATK_Q7cU,(bA5)Y^4_Je+.W4BbWd+,fL\a<O@a@@U&KfY@Z]G(f;<g
Wc2\H<\T(/?fIM84_F<<9DU3?<:?<+UeHeYGEU0c\S6N\HVGI-KZ4V:;;&]VRdT,
UU8_8RJDX@4LSUL9+99D-&??JJB]011KfGa39SPE^OHVeY]:KZ(??<W<7B1UU3Z?
>/-LCI+gQW\VV^@NdU6CC6:(H7a\B/IW@6@@:OT]/a7B(KA6c],@W1=2H#P]V].P
F887H>99Ud>dcWa7+V5)7-I<)0EVg>QJ)Ga34-X4[TKTXD^S7Y;5DD<G^(f2=1PG
aCN,W::Q)G5I_U0Cf[DfNU,,HE-B4UIW;5:LR\5,^9WNRSGF[]U.N&9U_]]Z/IYX
69,e4N<?FLAJ=D.G5#KSIW)N)IZRL]#.Z7]ZIG<CR)3#YCb)WNKaMKDWFS0gF]d_
TW(.9TA0c##<6ZA8CG])3_7X9eZKGU)98ZTB[ON>&fR8.?FdK4)cG+NCVXH)W&dN
;?FDa.7G.Yf2e<E7)J+R+S)TCREc)K9)-#Z&Q@)>Ug?TbNO<a.\aecE=LafF:cY&
O6#BgA(Mb@f[YIH#:&^GcXXN0?J(9F4ce:/3?b0I)8:DILbL^:_V<V[FD8#+=)-2
<a:B5dK:0YW>d^FG_Z&>^Q[Sa-.abTNA&b&3b<<9Od=TLAZHWcNNM.4?O>MaP,2Y
\f=)&<a/_8AZ&,a3I=(eK0)&NYEb(KUFA7.Y-e#_M?#3G4-6:9bDB[B@<TfA7+GA
-aPcMQbSKFONITDWbE[RP0<3:.ZT[]AZVL(_N7d@9\+]g5Yb)C4e@@LL^ZLZ#42Q
-NW+.ZLCL2eJ0#_JFc(RW70I2>V88\\c0f3VIcKU.X]7dd.cW2Qb2(6GGce;Ke.e
^5S/^TL0(#IO[,1K(H6>;C&\_IQ71+J#?CG/O)#/+(F<[eV]/g7ZJWGeJK:M.B.1
,XT:MN9\YK(MLBFXeY3O?^QSIEfYOA1E>0&GYe2()/VG69JKW)0IbUCbFI8:<#g[
g[8)L72&.]7BZ\cOI/=QG4U4T-G[BQ9Jb;SPSV9FB>OEWe-V>OR).YE.K)HC8cNC
P-#NQ]\\Y#LDN8?(,<Gg4X<#YTBHNbG,MG9,8AWLa6ZY83.^_a\bVHAI+\(ZA.^/
RJB+^UUZBNKRF43RREL;V>2+YY6K;M7183BBc;IVcL2b?+)3g<CHRf&AfY/C9MEC
7<B.H<&6(HY<?0JK]MTJ4Z.A;9PL-34US0E]I8.P8Se1Dg\PaR)ITDM9_]VHBQ6b
5a4fdX#;0\\2VNf]#&GMLLeb?ObdN#b5g;HEZ<MU56?TP2ccgTG^4/73UNe))IRT
7a5+>GF<[>J><\)MWfPaIdg0b6DAf;V43IFWBLdBJg/XWaEJ:@4Aa/g<^Y^#VJ8&
/c:A+]L9bGa;>aE-027T.4-XCQ=VeXNfWE,X\E)-;(/(A+9CFRd_U1Eg<F_d3,3J
].ID=+3ANI1JBIb2C/-9_\0:\STO_B7]Jg^H?J3I5O\-9-)U@CbJ,3=&9&P(dG.?
Q4Mg3=)52TG6MCEHI3O>Ze=Q?7=I3QH6,S=eB8\K2GRGT&KVa8MSB0R6>IAZ)@-/
-_\f/b:Z/BTO&349S5bc5E-E7SD88L8J(NeT,2RScgWcA<AHg#ZO(1+SbDQ<V^L@
K/HM:BgAIS+e4N2^P8NZH-T>1G,D>7H#>SZ6,<^0(I\(0>M-OEXR6YbQ6\@^(.a8
a(HbbWQ,M[[A4W]?.<dE@+8,R.4J(b3=+]]a&ZF:V+3O>T,)&3NH5)EUY[5;C)9P
K^(T??+ZGM8;3[UaW+?a3G^<<YBZ408d>I7NE)HHDE,FUg^S;27\TC@O)0?083Qa
1Q\[&EG_c/U^A#=+<=PP4NP3UHe=-b[>6V4bAA;20Pf-&FdN]SF4)A9W:79HI1DD
Tc;MN+YU+4XUDA9:ec]A]+<,[_LBVIB_X)SN]J[cN8R7\TI@02Y(c@]T1Kd\[)U6
5ZWZ(O;F8BDM8/(d@@[gFRb/HMP7)901gY\^WL6K8[4ce[;BI\b5D#@Y\E;d:?)d
:OG-a><77&9MK;M#_VF@V;WN)9d&K3A+)]R,A<g,g-=;5BceV4(2PYWb_72O(R@f
IUgcOX(,aJNP1^DT<.F1]aQQND_])5?3PH+TJ(VWT93dLg\:bTPZYW+3c.BA9T^e
IRfV^X#:9@NMbE7)@[3Vf#?ZJAQ>;HI+HeG-GcXA:ODbYRE0&7IT//VTBKBYdLaQ
#LYgZa>^-G\JZKMeBeB4UHg+/(@(ZQY+CND[],EZWCXAPTZV^J_9O3?fEb+\[WP6
5>=OMPcU)#QaJ#6J<_[<,e5-V\===@f#.JNYBaW;M0O1,JV.JAd+V#f<A3<:AF=a
fZ]a]#W?;ZB@#U1BX323c:)8I20fK[,,MaBeAS(57@KJPc(]OU+R:+Z[9/(C4.H3
IG@;3FHb=Q.8GDAHeF^NNR#N/2(<X5KFM&/C0fL8WEB\Dg?Cf\J7G-^6K2TIA>)?
@[=A0;>5>#_Z=^H.E_E_:L-bX+)U/W0bRe)EIfG3Y#0;<D@eYPQ.@Y^3UEOG.99-
ZO-R92Z\6_cG=7.+a0@J@RJ:LZ:eZQF]f5HIGR^^&g2L8E.dF,=fD-\3^dO15>UN
RE<ZZ-Y^,&FW+Q?#Qb,_XQ;QJ<#DV5Cg#)Q:]0EBVRK+\^&>NYRdKQ7]c;c;]18H
#^)Qeag+0ecP)]BE:4eR3A6dJ;0c-,R<5(NX?_,F;0XSDR^VWB1D:d=\N8;O?S6(
^I4J=Y]Vc=4CSQXeHMF.#J)a?Baf@M;MZSc(57HT^\g2M#WX\?<YJc[IWfda+LPO
PH&DKe^RNUe1GR&&Z8.3))WCHSOZ3CYP&I3YW_f6U?:7JZBA1e1.(QYM(9XNXXdQ
22-<E?(LfCHJE,4W(A8SZ2>L40TEG,/V)O;VU^efP3^MF68U1YXYTZ-DVfS0G/-^
_gI)eHG?G;]/OKcBVbQ\#8-M3d31F:8OVb@-WRZ41,/NQMUJ-bR+caK1Od4RGF=?
Pb=9UE=Cb9\R=283IR[XdM2cV<,QKL;=_>T4ba_T@5K>4=_bU-eHQZ/O6?PGd\IF
-N#CPFg39WKS<HW2&OS2Z1.\AW@KA@9CRZ/8(c(3Y8G?RX4EaF4QZ)d\gaf3/0JV
M0;PPg2AA1aZF:Cgg6#?2\-KM2.e373eMZ5WSD:Dfd4X4RNO>^]++D1Vb3aX\,:S
^\:5RJP2+Z5_)<=DF(d[0\3dE#??<5eJ.[QXEB-/M:L->5#(#+I\)NYGN+AE.&S?
]-2/baW+,?.0=PDD=4AYSV\KVQG1@/8--dd2QV5F3IfGNHc3],HBYBgQ5f-c6.cA
)/:beN8&Q(P45A=cF89AHNR2IN](8IO5SMNf1e+5[3eFM6Q&M528.P107G8K-eX)
b3b+XOY0D@)X01E7LJ3P=YXIQH,8f\I,a?B<^UH&;<T_R.E=G1]8\3a&W:J^(5;G
4L86U=1&RF0CEVf-c=cT/4KH1GXJBf4:9d,Ad+<_OX-7B;?@2[D8#b@\3+?dN1@Y
X5@ELZ1PTK)NGH>4>TDdL0e<?>[MILTWT<bD>4Y)AU88[S<N^EQBZPK7f=3bX#Md
C&D(5-3g6XW8AGK0N&Z35M<]0S5eE0@,04dKAbfgLd\^8(Q[]4?LS2/?]Lab@+cG
44?F=/KD@H=QW@b(X3]-D0Y,[0YR(B84Ib>FT[Va#b@]Y)&87=2WAK9d1V1NP018
(,5IDYB1-B4O<>>9(7ZBLHdP^JY(RM9OY]]:#@(IL>8+\cI.fbULIU?</fD)fe#)
KHOVHKJ&dRY+2Y)+]A&FXc>@99T]Z7+c7B@gC;4/6&TB:g&F//6@6\6[]G0aW[V[
H9^\d52<ed^,PH4170d/>Z4S1Vc^Z7K?DE&C&db+FcK(V,K[(_7<S].a7:GM;#J3
(?JFSUL31/Ce78]5\d+Q3>>K083;?VFgPg+6CNegbTIW4cER,3<_a@)J.O9LX\b#
MDI8W#6Ca2V/1F(f=>:N=8(;[0.R1^5d6a>N,_Z?OVQ1@9>(MR:3<R8fU2:A29/.
d/bJN485ZYO0HCg5H\EVJ31MA7>(c?ZIC(/R1[0U55MUeE[&J4Q7)\[,[NPH+9I+
eY[[E)-RS1ZP@Q,PAHMMBg<,,2U]a^B_.aNYN=#R4>^VS]K_+.943O;g),7f>><Y
X,eQB]R;GIS-PH?^eO)PHC^\6F1,E-:+M#^6S1;_c,;/_<[Ygcc&VR2]RR\[L:RV
(239.L3K(50&^-gF,_;.)QQ:G2SD:7=^EH_=e,c@FWgP3-2c#>aG\2aa+XVAV^(S
8VZ2T6/YZLIE/:H:I/cY_+&8Y5a1WeGefT\E36cc;VW;X^?>V=++=dKD\V[F6,?[
#]\5L0OMML_\H124)A&G@_V^G7,_G6[MNG7KUR[LYfcS6_4K,3F+5&4VGY0aVOIN
b^T7=(V==#K8KbXa4C-2=R[VV6F.?R[3B:IH,1]=6M?PZJfL=:=^KW03@4XD)RHA
#<MI[J]<X8[FWQ:4<5M(Z0bY[HK8SbZ?](]61+#US>ff2X?7E#BR>X8E-)Jb/NT)
CQ#AOA?1MS@+Ne3/)S1DU&H,AH[f]aM^W6>B.^Sg(.,Z;U/Z@Db#_3@/7cELAN_S
cHC.d[b;)a-]A;<]W0;eHGI0^^,LO89FD8>6GC[5\d4B(V]6;Q8IVEJGgM@[F@,T
M?3aPXT0]ZAW0)gUQNF4=EC:WLG6DR_SZ/]=LA@M8_c(H=S-M=cF1V:@/SNP>>RD
[-FR<M&;cYP^XcH&A6QAZ#B\3R?+#G&.]XHT-X<>9Y7(1H@1LNe#O,g3N=OGQSD&
E-GSA(7^A5\GA7aP)T\VA#9VMXSQ83RP@@C0JHP10dSL/;.V#6Bf>;Q9#=YEXSW_
06X(NNa_Te:U+Q;?]E1^9,WFSN:46d,=VC;\V4\H>Fe<)g:+V9Q_a=\;L02O_d2A
#g<QS)N]BIO708Y?S[5UCWQBAC=[dAI(Y4A=#QF/5LX7]OA5\aZ&eQB5#M=W3_RS
:Y6@Xa)3W)HUKM=d9/a>g7c@.,,3F2[B;G9,:QY_#d.OFXCQPNf(DP=5JT]9=41\
DQe7(DJWY4CaQPDW^F9\)<0;7Wab[9+]A]98PW(698635<e@e_Hga)XSR&VaE8+:
8^#H+>9c>@7]I/Y-IN_Y40DIQ+WPV\T1.]C?R<WFVN.DYL-9U?db#&M[UBZQdFUd
eH-3?EL4/SZ2QG9fD(FCL<[K:^<<g8a&JB\bIKM01_U/cN8D(2<DP.8#3>VXB][6
)fCXa_>X8(;Y<)I)75BM6VD-bT@\5.:9G/TV<,):C:NIXVXCdCWX89/ecaLJ>XUS
ZbHZ=3M-1=2aYc<f\N,(E,W(WBb;#^FE@RBe@7Ng;B#SMG@eD(627B<\P=FTFV_[
UO.TE6\+G47>^FHMNSOX-2(K<&;Z;HJF4;30SY7EF?6\Sd\Oe\1X?,C<^SY2eNF+
[034(PfcV-_4:V7LI,e>_6&L?3^,.+V@]6gLK>W(P7TJ1@#L+CP1Ac0R+JIRJMgW
:IK80-bY)e#,Baa6][.=[8K__]F#G:2PFR=85AdeC(KcQTRP51X,aX5gX21HGIIQ
AWD_\207\I+BZA)(E/[AfG@4BKgOX:2eFPCDZ9SXN?>&-@+1O:R5fN-;<7#>QGYT
41Lb9PPJ9_(HZPXI?aL)RCJ05MW6eTI;&:,AQd_YcW?V.9/UTbZTK8+Y[3,gWRAc
4V9GB^#P-E(fJG12b-KZSDU(.24RQEG60H.3G20X7N,fGZ8,]27][>N_09UbIS[S
dbb9J&@&7E[P@Q(TaPAS;JQdYV50?_ZG3TOR@e4gPfP[3W+Cfd)LVUM)JOXDGG]/
)KBTTQb7D0V(#S<3WY?S6RLJ3NM,1D?/f+EV^@8K>]=V3GVSUCXA5URXN:JQY3d0
F3OP647CRK7A?f>-^@Y@;>gLJQYS&[\MCITFFD^1<;2c<X:dec=_0,\^NR^59R+;
TYSP>X9ZSZFg4eD;2QS-&H[f2F#1@=.H+()EeWbL#5WT5O9.CPeB1Y:F](-WVJUE
<Mb+0PRCKNL\@MB_BVYb4A7aA(f+X(AZ;25@W/^J;C90A@2N2_>Ef7U<A;L_&_5.
OP3=H2UR6EH/Sffd[BcB07(,AgLS,OLA>3gdV]#@[:Vf[11P>R)1U?=Wc6K,d^(3
b7HeRgUU46d0TW<;]5XdK,R\g^AHEgc;PR:<B8>M9LcHf&ONMD.[-)0Mb36+>7((
2ZbM<:,YMX8XR?ANHQ2N(OdfUf)[X>5D)^IH1G9bBE:YHE1(<X8^B@d88+S,&IL9
dE.7S)e=T+W-+GI=B2FS)K8ZWL8ENa:#>T68MK?Kgg+ZZ(B_7g<I[Ya2[#ZL^]OM
cc0?aBVU3PWM^COAIZ86SS4;-/+CJ&eEK-R9QK]^>.L]5>0W.0,.bLY_]KIa4IW[
7P8A]CD3LRL7GeXEEU^Eb,&T;S?)OWU>[]C(,N4Qc&bM+F>38]_NOFRVA;gL/b?(
Na?5Fc[8c:)<8B[;<AOBGOPa\.T92F&HEFC5dVg(L@UV@=]QJ0[H@cbDI,33F4f;
NgEJ(3YU;;[KGV5E(]Db20(7Y@\J?HDag_&/;L:S).&VF0X#ITK@=Y7V:AWX#:2-
V0E-G5D8gd<(/aV?Ne]<-BY#4bWHX:58^[EHE;4CZ^R,fb=Lf69X9.LEJ>7C1=CG
(=SdCP:#edeM#@CeWBT4P84gLGX>/,T<&.Z&I\Y<-PL&80TNY-[&YS^?_?f\^ZW9
Nb63/X8>;JEO3:T(dYCVFZ_W>YHa5GO5)J_8XGS5G]A,f9=?KV.acB>]MaO4eUe>
@W#D>cZOG9/P]N1U>eaZ+\4aaZQP@3>9U:F;@dHJIH@_2<5RO.JR44YXQ(^-8e]7
,bIXT8<^8aC2]@E7?S9@WT)(_)[OZP7V&Q1NX0cd7.a=Sb(;GX(M;g_e>RYJSCeS
9;Y21+:^K^g?7QE>]8@82g\a_7I7NNL/;N_dbS:#]X#9D3]XU=>#[?F=?4SQ[K;;
#3@0\ZgAL@1E:,F_^5:ZPb#KL^>^R)M0ETLV>U;#E]&G)Fc-+a534KcP;+eRg,e2
G:RE_9=QGeDbdB]58d.Y/FDN^),=1&G+Nb+;d7C;\(;JcKPCaPTR=[P[VZ?XEGQL
60_2U7\EdaLJ)f_HgJ180b7\_Z4d)PG3D9e^3VMNYEV3>K?A)L(=DY.TN=4<3XPS
RT]\Y3/cPG.U:,YXLGC+:7E=7XLUD/Q;^?^;#VcAV9VI:;;R1)gBg[@U64CdI7T.
c7cRM;V/1)9c8:fIb9MY7f.g1b)BPHJ;KY:#<CReaONWOeY=2[+B.Z[A93d1f/LE
e_>)=5ZW&-a#V^?g\L]]Y4U/PF/47cL,68?0,8Qg7(][;JVFF8;/2Rg)J&HecK1^
cK9>13f>E:#)bO:AUAfb[d1:#)C4<cI#U^]]4eea42&#,Q&[Q1;Kd.E32/dTe]>\
N/>LP7IMFG>_=2-5M)M.d?FE9B)^a>MM;TTWM1?/N:9T\(/RIe@YR7Ca+SZ,W8I,
8_L]fd/?e^IA;T@=;-D](@T8C=Ld:5X:/JW@)c=J2+K;;O9g.R271Cb1QZa?KB\S
LR1.Ud\bK/f?=4e>-<YUd5.<fC(cd2g5X=[JY7O1e)4D-(;,/^>Ie80d>(T8cB[D
NS#cT;DZc.d-<+8b&c[TMIVJ0Y)T6e#L_TJ#]NW_BXXWBSIdCP./-.cXG=7eH._g
.?8BN(B4IOU#Q(OHY0[?\72#1CT]N-g4E0&K0XRXKKGa\3;\PJNAEM?OEc1CZPB\
.]f,\@JcVJMEI=K)8ID8cJ&+]QA<9I6F^fR[(CMOeBT65]E\RBX?a^8CgI2\1A&A
0^>8Hg\#ME00G[N)X.61D4M&gM7Z@c.[@9S:d0/OU1,HM-:Nca^A@Q1/7=-b5GHQ
<?9#\.+?4AC)K>,\?)bOD+_=,E71X&:2D[#[/131&4G:CdMEO8UfCU6,@1W@X28/
fPf3GSG@::MR,96]?E1W7:g^2P4C>I@BN\EaGWE)S5a1@SQ)/^)T4O6^#eRM1J)6
P:JA)Hb4BRKc4YS++O(J]Nd5E35N=_VJT\A;>dE:W^[(a,[0dL5)8>fCFA[c65B/
@BE^Y<J-<#O,KA/IVSG#2]VV2AgV/Q19Vd3_#3SE\?YS+L\:=5EEcOED5Q9I]^J&
EP=X9?9=3X_EZXEg#Tb<+3AIM62U141)&9c;944G/f+A1LOB:3+.WW9KK[GFT<7\
Lg;PZ>9d,GWL[RAa<E/)USY>M^>d4A(75+2K5^&5VB/KK&#D^&g:)&Yg:ZZUZPGO
Y8VKa>-B]@S,Lad]5+-12=WIa9U#ZN<3Y-&4,_8Q-g)b6:ADb[#RRNaBI^\R6+IH
_V2a;IbAQO5QMa=IXWIg[[FV.4_)E\;DN9_@g+Nf&3g-HdCT1_XGZ/AE&W]137;K
\J^b9=WHdeP487IU+bKA_d?<0TdbRDcMV>U#Z_K(/IW)1H.5=IWGN[IWR]0#/+@A
bP=92-K3X.4RUWPD)8@bA,+LDeQHV5AcaH5d@>4J+.2H)SIUQ\c-f-DYQ?RIF.f@
)PZ28Wc4+R\XJVI];Y-K7Y:=Ec8TL/4Md=-7gg92^1+:&\c>=5<<IE1UDcZQ/W^b
M+Sd_8]./+,4E73:eY]-54OdTaQMAb+#I16B122)d@b)[;,cG.?BC76MO2LN+IE+
eAgGR,]^dM(>dM<T>(EXbBJP[5.;d)Ja@6T]CFGLdAV/O4c^#RfIUB<\;T4)Q9V1
T_,\GEH5DbZY0+VQ2BH,_H?ERgRYT\26V85?1C:ZRg;D;d2b?G),O>\Rd?QRd=fL
EY)d>;c(873bb(be-&e;3:.dH[\<_Y647d5X?QI5a&g;c.Q>50e-e0gE-)T)\.TR
g4?OFZ]NJ\P.8:2b4:83_RXdJ?D:W<IA4#]8988HgFJ@F),GO,?M/a3;42gcZ447
><[V,=GaC&6?BI61\Hb3MIN[?L^V(N\d9)c5(S;DaDf/BX^M_fc->;EMIIJ?A6fb
#F;.6FS4@VAH2UD@@]1^)&4I5Y-TPV:W;EN:M1[AC<b\7\+7IaKXELN:T.H.HU&W
3PBZZ[=Z^G>:6?2B)bJe&Gag?Qd)SgFIR[F?2MJ)Z3V]NS.@\)7>=GG9^5:dS#dH
Gf1MN):\MLO3+=)E1T2O5,9CPRWBKMXB[0))6[FM:KD2K)?,(/VCD4BM#==9&QD2
N]CR]If3#II32#:bXYK5M;5&XM^/^LW@b4N6:M-K:+)R-J3.)bU-G,3(>P@LH)]M
WZWbX5f=LZV;X^2&EV-faHg&G,R&1@1P&JR.R^W0WQ/eZ8WeGADdSA+fd,M&+H2G
eUR+D<,J>55E1Eg/^R;_YfN;&T^eI97^<D^AY3aU5Q_BgKd>[Q9CE]^MP-YHG,0.
f;-/4a=_K[DUEgX\<a7SE)6NS^/f(0USGY4\[&FD._XFb^=G9:gDg=^MP.d1:/We
-RN:HAdbO@1-5?)RfJ;WeVVELd>2\_9_cYFL=7#QY>X@?Qc_H]2&ZPW^.>LBabNe
7G),=(=@N1KQ<4A=JVL^M\H)&2.]O(00+aS-58DIC2E8MgfS83ESd)G@;D?e(\F6
07Mg<fGb=W825Z#42J9R+K0dI6->YfY6WTVMQG--Q/-.#K?dRBLA@2FGOeD]J;U]
#g5QUD33gY:9-4C\#LQOK5HQ5LZN#.<SOQS6A>[:Na3IA?dK8G=Y[O^:<9>8-T32
E6<dF.@ARIIWH],)1R)\:aDd]FaACKeZ-2/&bW:=CS)Kb><[__&OaD)&.G<F2C_.
\F1TGLb6<M_948;;;b(eL,cJW5_>)P)UH29GGOQ4;1Q2WQWc?UZPF67LGXPe^a,R
Z<V:J]dLU/WGK+7:#[>2f^F35Sfaf\1I9>aUcJIB_H^(^bI>@:Pd?6DO_=C&JQBN
aCD.>2ZD[2\NEDAU\7Y3[+C)<?T3ZX/@#OR4&/[UDgCJQcKG?+Gc:]L5D/R/-NA_
^Hg_9FNV6OL@eDEE1AGWHA5Y_/I+@=Ub1[<).c&JeZ2+f=b-T+6D7R8b.#80cc+B
ZNW8UN[@?5+fMGeP#LP&gP?a[G]Bf=GdPc[Ud;=3R^_@c\^4-(N?9[-=Z5#Rb34C
C)-eD[SBB,(3KYS=QL@FUN\CNAM1R;aa\g8SLRTHeZ.c9>/)5(O\=0<HDNfHM:M_
H\X1fDbBVK\6X[g;TI.VL3gD-@L]AZb2EPe;7af7>d2+[=MQ:Pg&_?R/-E<7=S^#
]#8@\+D8F5=Z/a=)8V7b+_5DX2/X.6FE@>>J9CB.L?Wf257ECX<(e_Q3eKTN,W#D
UK.OQFPa4Z)=HbANc#67eO6JB<@N\>SD9E=-NY)MYdeT97g_3f+8cC5XQ<BY8D_;
e>=,UJW3F?/5L][H5;GD6I^O+(f@\\2PVbI9@D,M90L;#a.6Bb5fRN-W1/\@^_a-
O=5SV)\,[=fM^,2OB#P1L#T,B:FNg#C(TRV/a7^>@@LF=Y&K52:g;-aF7Hb6VRGH
<E7OUceCU5R4\^E2Y6ATZ929d9&8C&/==(4F/G=VgA=RL]RT</D7bXF[,5FPN?O2
@0^(7B:-Bb(BO+LI6^eRd)a/<>]3N;7_5\0)56g4f-?gaEA]2ea/4V/Y9Dg<@@7&
abEOD&Y9C::L=RN+_IQ9O(74MJ@Ee#7T\EQO&Y\O[_?(>JLUa)>?Y?DR8L4#dD)-
EO4WAG6VVH5e[E9A.VRZ_g\5KWMa2<REc0SEXGV0>@DHEd[:)K?]&9dD<Gf_\WHT
g;.AD/8b.OcOH_8&95gcf-;@C-96V+HNQDLc;7_T<R=NH8O+HeR.2/Kg:cR&c5S^
fIY=@-?D=afaf4:QD<eBN48[[U080^CG=GffEVQ2#Q_Id;CL?F(&?_SF\DO>96:0
POD1\cRI,aC/)8.:W:_]2&[M.fA9>=7H5M?<GI0=^_d[OUE<RW0V0D@0(NMNU=]I
f.;+8JfRXW87T6=QeNb>gWU&>2[3Q8;)dM2d)MDIOTBfcJc=L2:@U@EUUdG6GF6g
5[;T:?Od8P;L+g_#(PT+I^B,(EC\c9bBNEEe16fFV]]OY=TS@;&_LA#QeQURP:^B
X_TWW:(GTgD6B5#E:]cB.Y(3;CX)BI\[I/7F?F>.51IWSf8RaCGAa,;&O2A(f4OX
7aUPTG0<+O958Y^Pa3Z8LU+cfH.US_e:R=/[\?(eOY:FH#EQ?P(GO:CXZ-D\V&8T
fK(:OY+f5.X0P#aO\@2MT:\S5]1O>:V7],-J493H?B>Q5:J,[F/&L002_E.BOIg/
0F&T9f0f[64T44HOe/Re)Z8&#D3AB16D^24+SH,DV3Vd.22QH#0<e(FH7>#O:<Ka
,B0f4#/M)NW[M.DF5gZ-^)8dO5I9;IF=867QLT#47/&G9CKU_Ea]fR/;K-@\>9,L
F/^Kb^-U6Y^2KcH(FZ\PP=A^D8&?(T<S]&WXDDE8>NcL2R07E1R81VOW)AgERJKV
fR-MQJL_93R,CD\UN5aIf^G5Ib6XI&[-Y5M&:1WE<(N;_@eIdM+cK,H^PVIW0R8\
08NU)EF89OY;M>4R#KIY[6&#WDbCf/A]G4#gCS<=G=O?#0KUZ&H/29+,Y7aQ.1?[
_fVIAK;Y/#R[01dI>.8a@[630bd37bbCe]CUVROBI4N:M]b(c7F7+[]^YL=QOZ5H
P]B4O\]8#02K_KUDg-Td-NKQ-/+HRSWCbHO/+_W+G]9C/9Z9TD/K37cPIVfI-.0/
]&=YNc)cQ=d,G>-;=?/>4:>UYEQ4PcTIO]Ra4MgbaM0>A1-F?P[,C<8K[,/E]7a^
VF\#c7EUc?4&^YF-JHMB4e4;\\\SI(:U;F.M;dbOBeA=<dU:Z/VFeUO&=I-AdY&2
\dgagLKH=cV;_/V[-ATf,05/8@7+PHDW(M7:T&\4DQ_N=4(P=N8BZb_[fYc?=AZI
RS9SMdC&9gEX5>Le&@7cIED4X;Z8:U[8f2<DXRI9O@P\HAZGc,JVU6O_4-/Q=L66
+.a[fQf^_eF+(ZY<S?BS^[?c;@1UgLa+^UU#Dd2?D9)=NZ9@@#f=5SM]N1gc3-6^
+I[IIFAJ(X_#^93>Uf16,.F[A;Lf<5aXFR]:=H0e<8\#2C2QIF8CQfBc@YCeZ@:4
(L=f=6)dLMd7?gb+VN+S/UM?TJ3#5]E9eC=?2X2#Ic@S#W8=1BWR2VR/?@gaEG,(
/<4c:NRQMC;4:M.]Ba.\)\V-Wa.gCP-L57Q/2K@KZK<K[Q[+1E5CDIRcOKN5B;(H
0][/PLS.IS]9=>g7R_c.?E&Y?O[OBUND.Sb+CPcJ4@a#P&+KN>6R30=35gD8>XfY
5MLFZF?cScNNaW_.)C8_40+L&2bU>]\;6>IMM,@NUIUX9MDWP;U<EA],.IOM(66^
5Ic_Q;Z^(00EdA^ddWf2eeRVQ\/@91L>-GX#A#.W@\17N3KZXW,8]<HPKPJV2L&^
4&D]e/4E0V_JX4=g+=\XeN:8+8(EA&>^6c=3g&Q2Z[AS=6FDg&/8/,fZZJf=EAeb
;MOc]OAU/UTY>cO@;T#)M;T]4\^LVU\GTV@M.4H@VT2[I,:\<9)THTEBVA0I.\T>
Xc<FWD=f;a40.-WDE&TA6ZL4&6Kb694K0KP+4a\F2>[\(:8KfLJ76PE##T7WDK]e
&7L1TU[#,E38AEbO[8eg<798WII>d[D:dB<Z:,fF2>X6C4B6/NGKa)U.Z1O[^]^U
:dcc6b_FbG@G@J+T\<LXO8M2ca,&I.dP3B)-,9BPL:GZ3<\MEHWUTg8N)3d0E912
=H]PXMb_7V<?4;#@-+N.D<Qa#>U,e:>FfbD<_cb.8#bTT8/.\)>]#CW^PHL417TX
>g68INSNfBd.GR3KX(H&)fJ8^d,+)NFbTT.[XL/M&6L>N;#?UfU2>gfCF9C=>f\7
F\1,e4O+D#N9WU#e[;a0Tf9U)1]d,N]2&);Scd(Yb<MJ=#Wb:9]C;FO[B4HB7T5?
SfJAQfRO+:T01K877R9K(AK[1<6:-e<Q+:01X4:5ZXV<5gR]W1O?Vbeg\?O2&DQ_
B6g[WE3D2&>4Sb]8GgJSL+[_71;..G=38^6b?(T.Pd0AY7@,gYDDP(-#W_)]1g#Q
,NY#TNB9<+P5]5f&.EMfGR\f1=Q>:)3#RJ/WH3Z5d4,HHIGD?f,Ne(O5[ZA,K^QZ
RCBG,H(WQ[E;8];CL=dUSb+EKO(1-706.c9DaVTW.7J0E][CAbU+:cUKCWKOL76Z
f>Y=cV679HF;)4(#L#E+<TP#DF84<KO\[,CI-3\=[b;.;#+>LXHZ^RRXGQ5U\7e;
A9P_+4Kc+.>GBgb+1R>T<P=;bXAK-aU#=&QVL5K,BLG(,4>DS(V-R4L(I/P]<OBN
F<cTCJeV>(]<@^eQc99VG&a99)Y(bA;fWQBUSK.5Fb,_H)aP2gTC8@9^fX_:;&Wf
=&L9NdY#4.[^9ZO?c\^G9+^<F\>BY=)>f+_?>,G/+.9E<JXPF0V/;+1g=;+JPc&-
\PZJ(-WG/=+D=fRgGHUO>K;++TF]M50T9I5S).2dWH4B6,+YIXH6aZ2IVdT1@/&&
6>\VX[QTMLLJ91JUF:R:,V\fU;@Y7fYY7G[c_CY&]SF7&E#;Pg.UKJ6D?F_46E8P
Z<SeUN(af##9APL2H@O=Q2HPQ136AbV>-KMT4#NU=TaSJ[a9F-G,Gc_UgMfN25>)
eT;RgWJ9Q8+VA-Y?OMNT@_#aT307&=R-gYf3WQ[W9D7UaS((KH211N#H7E88)><d
X@@53a&#R(eK5#-_C3O6U@YG>5ed[T[R[S[7WPK03H_#869K;7MPQAa\=I.TNB6a
L2.YYIg)L--^bX8@H/;-)D<7)C/&cOg0MP+;H9(J>CXYDfa3\GN0P(2)&_1A9#J3
#AH8#&b_->1,UJ7.M<##O)a]BJ[SRK_C4#40d[9K0+W,OMTK[1IB66gT\OCB6]:D
\JY_0P?S.:>HTFI[&eD3[0>S;&[^ea376]6A]4W.6D^LXWF\;TN6(f8;TOW-c\Eg
bW06N9+6:LTg_G+>(ObX;.8,ccTI+((D\4FQfHb;9QSU5C5KeTER1HMBf</WW1-M
E-/bEa>A_@eLTS?NOA+eM0BKW2F/EAU^XeC:1Sa64fVb<.[BRbbL^8]eTY.+HFdN
RPQ^JBf]aZP17B3JDQY,8(aJ1dgKCAfXNAMH+6U+]OK8DS2[R,@0^G?G9&,IW1SQ
Rb.)QGD>dWK([AG9Q;EP64e#(6C02E9A(gIDb]AS-.@D8[^FUc6#,cA[K6I?[O7P
MBV9J4E>,?L#cg0?=0G-:NFdQF1[(&2HA33f<1d?K2XfcML=SWQ2-+f67aS#cOWf
.41D3Habc5:TPH6(S8MU?>->5D.WeNF_HN?3f<]LD9_+LIKdg(9b[8Y.@U^P2P_a
,gI64(=Q:PU+K05;e5\Y32MbgZbC1f6)]MMaH?^NW>aABOe.5T830&@AOAV29Eeg
2[7ZH0[Q[G<5,a@c=A2G=-HJ9\D(5eH-_Q0^&SNDWS>UE-/cFI^OQ7]B9M<bD#[;
@PA&HV]).4.8&^D::;JG(EKQ_R3#08\J6?b9KJCM1V3XW)C8+Lf)H\J5UX1\D(Tb
UJYN9C8gSab9,OOM<4Y?_gR,ZZ)QOaIWI0V3JYE+c?;G27IM+:\>A7-H1c]MIEQ7
.S5gZ1Fb][WH,HTIE+DbSg>,^U;U^9GAD0ETe2LWeN4AdW8HI:32R5XFMT35dV7Q
B2#Od:_W)Fa-Z>45CaR/0_:ID,=40\]#F<)gCBHU__DgARb98_.=gXL]&eg(_ffN
G9=_F;C3_a7ND]<[J440AD\2W<YZ-2>A,c[87<Kea=<NNN8CXg;8@Z-b,RO^#+M_
59S&W8gIOdcF^EB;]Db\B:O^(-6#T.9/Ja[X9NXX-Ze>/5(V[TL\W2OC\/0fG,G&
RV##DLRH3+ZBCW?-PAT>X_,SA,4&_Yf&J/G#>SK/Vbg247J]bFVA;B-GGXL\b(-R
/<KQ&A#):=O#]KXgCFOANRN96(EXEdCT,NRLf:ISe6^aW1bdDPG(7-P.gI=c:JMR
<42\]9/]:>E,?/cR:G\[D^@<gSP8e4#O0AY@[=&=7OK[Rb9P05#9UPdNANQcLA^)
W3)Y6[+A#.\EMR/XBe,LP2@afS\BbGd)[aHD[c,WIY/LC9Y1YNY]^KEHF+SD.M/I
KIYbG1#^YQ(d#1_XY&/Q[ULV(HP=J8C2XKA&SENcg+3II-KL;(-UF,(#-c+6JH@U
):7+C&U>^O;==<cFe&0V4eg2GUL;?LLKgA#K+X>URaWPCVO@PW7E=::G:NTgOaO8
d4UT==6?B,Z[JfOZ(a./[d6IVf:1@:/7@#dLEIYR)-^fcZW,>K<:0K=43@X2L)G,
^^X+ad=:-W/_TOX9DE?[<K.DeE9G^ga>W&<1DVc<>DWL#0(#UF;/H1(_P-]]<Ff7
TF8<@J248gQ=^FJ#e\V.2TCQ[O?Q_E_L70@0dGBbXBAeE?HX6SC_&e+S&X+LKPY:
CZ5WOPJT1PW)>\?(08RQI[IOb_P.NENRVTF.cLE:JGD?)DAA9?XP=QUCKMf9L=[Y
4/2b1OGTZS\_JJ1TMbX>&F3[&U9?.gE6[A4U_MC#7B6e&86H3:8E;+Z5NGP0IfUW
Ua2>d3WGJDcTTgWRXXQUQ9=V]Rc71T.35],d_#a&;(JG-?0]fd)H@+KLM2?d4&;3
I6GI\ZRPN6c<37-]ddYg;R.S1=H6,42Pd;g_PW4_83-\\Rg];6?RcJcHJf9Yad1.
_Df[WCFg?1&b@dDF2:?(]=;32Bf0W:5BIaYJVOf8#7:TYB\Z??bfAFWcZ9?KW911
TE57F6U5Qd?,[0QD2,@(>2CF29ARB0.2NAa6MX3[20DfGgg4S)A(fLK,@Y,ZL7MZ
LH1&H+[acS)OcS:8D[[?.0TF(N2TJ?g;<F[HMC4S_\gLERZ#NZSOf6_,ISQ0IHML
5Vca9K0L6VDR.<e+;:B^,KGc6]Y3;U6C:#8&,e5):=e.ZB6APgI+g(FbJb506Xb+
+]bH+<=7(0XJ(2Be@JX>H\_)QRZ?]GP6^F#AdGee^CMCB_\C^:9)-g@B:1g6V[53
;g#5\]AX68L9.O#CVOdK#K9S20D,Ta+ePSG6N<G(R=C4f==69J0D0M_-C>4#a>[]
@16SP7I)NO^]&+d>PgN5A<J-]/BH/.aYK<=H.F-+9Deb@aQ3S64F@D[Kd[3K]=L[
^JfY_L2\\fNQTR1f((2-=Zc(6U^GSQ>QLCA,GGU4]a#a7U1V=V4VT/[Y+[f270BK
UaBQ/,]+GWE9EWT0fQ3>RC-XU5X--W]DK3?N=(Oc7TV_)ZC5-4Lf9L,-R47RWd3Y
Wg6\B,F;8I(1gMKK2V0.B_a=#KLHQ)@A#MG7R4LR0_/EPFSQUF6+C[),,HMX9&Y0
fTa?+3C0>2/H3YL?T8#4+DeW<V4V+.bJc,V[A.b/1@>JD,V&F@:,gQ3T;U]?N8.Y
ASW(ggYLI@13:&VFA/^S:ODSZON7LJUGC2?ScTBDX6H8^[.>_>?5ZQ_(f6e(HMfG
#3<XQ-5Fed2_>-=b(ED=.G6MER>V9QfDd34V?;_(?P,O;b5c[1Vb12._ga_G:GW7
6Na>BFU6e.^)(5+gd.WO^]/5TC_2B7KYR_NTedTLd,gIH08Fb-G]7-LY)/&LTYF_
QX]:=QQ8@-;bG+2HEe)9]T)1>I:QG)-5[2P+dKMb?1>+KAX3F-gO+]>H:L)[7U,1
GII]&f,2(CRc0>9IH4LSW#H^RPgUeC.g+V(ebOC:Q7#?f1(_C;G44QZ?b^O)1g.0
>VFHJ948g]E:E\Gg4YL3:]gUJJLeO8T]RC_P7O6/Z,B-IFWd2YPS/[RF+IDCN3JB
>[87-5dVPg@3;MT3Z;5a0-cEVQ6N1QP<1ARaAB@<e\eCaf+aEX[@]L>0JJFE2/<I
5<>\U2.0+c&B\;0X,:F<4.O#-K6fg:+=Rae?,&(+gbW5G2Dcf-0V-)XGI?<SGO^.
_:?AX2>,&)Lg?\2_6AK/4-?\)S-78-N0GY097BQURQGLPSe/]C>)2J47IHcSGecG
X(_a&W/#4E:;<9NU]>\e8c,d430ENN1.E\1)88bg(X94\Wf,>-2aIJgYbU2I])UK
HR-_[F>77R1CJ:P<FeY-+>gd002b>IJ216A>dI0(5)W<[FX,\HAJQ\e>PJTH(\V/
A>)E8a&+^JD2E]2BN=A4BKUSHQ8PH;e3Ac3)#J0^1K9^.T2.L&e1Q^QQ#>YR8M0\
&.W]EL\/@54D6J@)@J98B^.CXJNP=Ce2P\gUC0,ZD2W:&-6dZMEVBQ5#dPfM.\5D
-C9M1\Z;6f8b4YSL6f1GCZ3[R3/)5<.NL6ON]Vg48dY:&AJ:88Z6[:GBVPb[2T^K
SZOeR(M4GDX.9Y\ENF#XcQ-/ee-73O[1EA,fB/KP?c1Y46R7MSfQM;[]@Q2B&Q.+
Q?ZGA#V&b+>>K+FeZJ#Z4)HX-<<?>a)\RbGXYXD#ag8:[c_IRH6^LTR#Z@b)W2#H
.L:CTGHY3PeT^d/\.,#J-2.b?>BVNTe>1AWV^a?UA9X@gY<F#U5gOVe_c<7LKVKf
-H70&;3]cLSf-002fWN,9_3^EPSg[dYI<,?:D1<B#<1C=O]355@1SRd[73@M=)I\
,b+[3F0&<&>\_(#UF93#_GV^()@]-WTQ.+QV/<?-(Pf;X.K#ZPP10Pf@aKbZSPX,
Gf>EX-1N#4X#FYAV(f:MJL2J#B>LXT+^::V(Nf+E+L0Z[1#3/HFLF/,MK=2E<+K<
T,I-0;<5A8XLM\W_VH9eaKO1K,\Q]^N5e4,F53d-KF?_0T;PUP+>S,3V3Y/;ZfNY
c&=_M@]@MLHXTZ1<bfN7D8V=-<TYD3gR0>CO6+DPUCMDH3IR?#(+aaLfX^fK=J-,
1aHCAMUJ\F0#X_7135P:fEPW>4>EAbE:N;:4G1FVdYXM_;?9e/H2-9[;RfN8;V@]
E\R&RG5D#<U1L6ZbX?\1<@UBU#<0WAdg2RQJgDe//eQdZWB)04M7CK@S24DMK<X-
9#FbQB1b@A5=]1FgI+<7b<\QI^Qd(+-9e4bL=g2ed?;9O<,Q0YcQAcT=c+7D:12c
I,]YP_#O,698_eEMgg5P5H@98+B4Z.ICLVJHDGL@MS(ADBc#HbO0&MfRH>64:E?G
JRg?D,g8-]2&AKbHSfY^9+6H8cdIBN7-gV^VG.6e?g11)&W,YHeN&Hf75NJQg83^
6S=:fQ4;;e@_5/;W@MAN,7[NT5Ncb17a7=d+\JN0Y&1dMg9E\#G1f.>KU\OJ,:R3
e8T8gWGM;:K/RY2W/9g7Ec9<eb=2\2E]Xg[\QPcL(;g5A2ND6]7#WZ43:^HGeG=?
a:6A?OF&fB9e4)I5e4Kb+-?3OPYeNOcP-O/a4>M-&G7.+3:+S>S60G:Q]LaQ#<VR
5/2W7Z=e08M5YSf,T8IYBZS-KD,,\&I+J(4;A.+cgUA&M0JBV9JG5E7JZX\3(e[#
/c7-?ZSP#3:,R21I>gd072(b12D+(?7(_U?-=eU]7SJ3+[=QE8RLJYP\9PeYOb(F
5:?,;(KD/8G@I0<dSINXcGPK=2UF>_g-K;A=)]0ddVRRT;1=<PV1;:55-JM>IGFB
=-]Z,X]-OSe>6DK^U<g(HaD/\Z=,a,:[(#-(V@9dN,8a?L7&ZKRB7);2I,N7>L.^
Q>,1KfaY4d0T_\We9#V6/8^A8]Ld#U35EZ#U&L0cSOa,8e#E@M\c;M8.7BFPaEg6
OR)[[3]U15GfEBW/HX<VM9=91E4L[eWaf/P_L4+QXYD\6H2XVf9H5CPL3;PU=X1E
g>2_5.,G1I:31Q50V]3.S_<5J4<ab[L2fC1LJS8YHN)#:]YJ\A<ZN69<]807FOO0
gC=()bX.?J@#dVDB5.P>?25C[CWPA<MG##.6?IXW+65XZ:<ZXg4b#aYb,:ZGb^Z)
:HDW16,9K5OL)cY=\T;dRNg#P:,J][-geH;OH];J3;I5021/8V?4HE3E.7=7(bX2
.@0#/8R#7IZE+bbFaCb[Bf59&\CZ6cW5WW2=4\7O5:EYA3:()C4D9?H1GYd&CNR/
4SJ+KLYS.[?D7+c3^8IH73\SQT6.6:BGF)9C,YP8:PdPZaVLNT,Gf#>G/C]AEO1d
;DM46J74/dCbBJ/TIE+X@<VA63f0Z.5257bG0a+VP4?7S:G<RB,<<<J=RM1g8;LD
<Yg#<(#ONJZZ5cXc)LMeWc3QF01G:bW6eeP]>/fRWdb5LV+KMfFP2K+Dd(Z6/\8B
?D5N(6-Z=Z7YZ9S+ZcZD1N_E6^aL_<G1\E-Fg.Na;_@YXA=.246YZYD0c7=@SZ>H
K.XGVX9<Cf5;;C<dfPS@X0(03Hg>9T^1fVPXTFY@fLN+8B/NH1EG>.6WJ:YPE5/U
M1CV0>>]+3egeLgdVY4]B6O:I698L=YK)d[W#VIGDMA?HXQQB9:,#gc1@?(?KIDP
7/g^^^)KJ(:,5&J86Aa.e9#;Q[\>X7\Y.@J<Y5c[HD2G>.5]WT(1DTD41a)De4Hg
c++MgcU&/?V.aUDR&=gBF&L(P/EY4/2gba^Q8/[bHLU0;:IL.<G6BS4Be_5TK-HH
?;\cTPUZfQ_&GCJF3&6.?dZ:eV&V4[4XIJ:7-VdG)]?bMZ2BQJ?F@3<E#TgND]?N
L)7?0VL+MQ2PI1FcZg4O=5.bKebdK+92H_85&K13Q,9cd=b^R(#(6UY.A)?:5T@D
LI^N^A3[5CI\[C<LXN,NP\897X(gMAH]K.D2FF+(LC7X?(R[cSZ0VSbIe0)IUXP0
;@@)C+UWG)7d;<)ZJTM?OD5GQG()[/7g0V1\D+(eG>A]#GH7&Z.fA.TI7US4E-X#
\)C@M;bed(#UCbG(3Y9FT4;;8]9UQR\7^1?7cT65P=:T>>61b(OJ\cfF+1F1]S;1
_(fOGH/a?SUG=^KPL,&F]5Y.<CNU@NNM2R@HPCH?[[eGaQBOF]NLX09b#+F_VBXc
?TSbI>6P,T=WVWg,S^4&EMUO#?b]D>#d,1,(4+Q4M=]a)A^B(EM3:_)N71N>/0KK
@;ceJT9,BO\H:5.KdH?ORRU1CJbDW.EG.KZg-+\1SOX:4F&e>Wgf_5#3DM1F,7\.
&b[Qe+2&VL#UN[++Q5;GQ;E4ON6>fR?\>R9f+]37e]K_KQWR03O3ZMTabg4Nd;DH
N1bCdWg/bLM<9\&D1\Q@B@g<WNN)dZD?BZ:_/)J,DSGJS+I7)aCI;X71LT[eD<IL
&E5<g/TUA;0>Q2M_54IAD()1]H2JL:fJ&f8;[1Q-?669O4S?N3_)?C3I^05@PP)Y
[U:_R[bX<>]B-f(3aQ]-K4QCYOR/^/H49(,K5d3[K1b1J@EFF734L[:ZT#4=.ZYF
N0]0E@/1[cSDNKSJ&^a):D/a]/ID-L+#G]<c:T_R,c46C5<;IX4]a@aN^-7g8?O-
)4]<L,a,bOTMO)5E]4c4e:0A-PZZH]#LX0PLLc0DcBc,0W1+Ha10cC-_:Q;Z4/Vg
5DHA@OTX(9AS8&MR=/&0X,M@ebN03AbcTZI:O3W;.+0D7Eeb]2e8(T/A5D<(gXIc
78-E7CgF3d-3RQ=_F\L@AI/ALS:C&gYf/X?E2+M@LM@CbA,@6g;NGX=F[LY-RYI/
[Ke79gM&&6O6#GbdV=U32MAgd-?KNVE]HeaZZ29gca:,3,bLOIGVH7cd59Re&94#
]Yc81De=Qg7D4F?&UYd9+aHe?TRd&[XE1./2:_]?>H\X:\^[:UKY]]EfSXROU.Oa
Ja8L=7E?]X0N-eJb)YR=S-.9X=f-40?gJMbeO4d;A&]BeIe9.38HUZcJ.J1H[KXR
aN;+(>01\JN;09RR3>>;8Z#(dL3/Te?]>:)/ND8dVY9O6fXN6\W?E#&4S/?)2XJC
dNZ&E;=e8baV/+g2DKJUYZ9\YH#ME+^VbJVQ456ee1)SfHR_.\T)aH2S7LE\MgHe
A;CO]A;Y<HcfeR9CRf22f@B>-0fHZQ01E+7@:=>;A&#5gUNT/fB_--(SO1=^?:KI
DX2^,-[7c178^/FBXb;8QaMQV(UWPV701Z>bRgd@S-bLH;AN8b]-)@51c;DN2=>K
#SLd.6/+X2\B@0Q2A_K]7P7ISg9IJ[][EWQNRF#a?Q(0aSB\QdA44)?ZX6&W=C-E
b\@a7E.)0S[-Q<<Q5+9&.X,.R-N68,?eadJ:>5E;^d<;,3T=-TAd7_(PN7[8#X2Z
<,O,?:WaH)_2fL\=L0:5WMLfZK,:FCKO0Y;;FNWPOZ@bg&M&=b5EH#T#=_I(AECU
[HH<BR^)RQ.B0>e)bZL#940G\<J\>PB@0;<+OLf8+fFX]a:<d<>E]a&OLa1-^.16
_&RD2RdK_e^&4OQYL@J,QM>^\.QcdJ0:@1#&78_f:^\1ce\R]MCQ&CID=f#S#\0/
0N)9Pe/W5.eCe-&+-_Y_S@VeKN5X-9>#_G9UG[gR7W(AD;I8X@PZ:8P._\bE;HQ\
b3WGH;0MC_bTPMf^\-M..ZD[F4/8@KS24EHXJABEY^a5D:P5;W59CL02.B5GN[YX
OTfK;d]WG(^SV5YLf2/33gUeGS/IHbS)(V@Mg6a(&,e/8KbYBRKdK\-WcRf4E<49
[c6+WT+#?FM]TS?DLG\WB>f<U=cc,N1Z<W#8Dd0V<^+R#D3#&P0JdH+<IX)ES//K
=(6QfQKT_L7B/e5DDSB;[1.2dW(fPD0-QWVA:,G&a?<\g^IUUW67NW-6-GB&E)]0
X<b[7Oe#NRW,b_BK4_/]Z/GKEB=D^,4_+H9^>]3VOLAC#8FXg;T+D0c:1C#MCII=
S5P7.TV0,FRD8cc_]TX=M96;=0@0T(<,G?S;9]TPGRA#9S0f=@_T,YRU+?^-F7S;
/AO+9-J-AEQR4H1FT_D_1aZG6RKR:]IAQe4Z(6-4/?@Cd(.7^T]F.bN^2QJO:(e_
Q;6(]dDYeXD&1VbJ51e)df@bLN1/\XL])7TcKBf?OLUUgR3_H^TO-EUTe#4TW3AZ
3.8[PXE8a=Yb4@-VZPa/f-c4\=XZCP)U?OYMUYM/@.@VaVOL>F1&7_IZSd=PbW[S
VCe.7C>&-57&G;.SD8?X=Q]YOM<)]7VVdH\]7BN?R6A6Q@BBH=Z:?@D[/@)MLAPK
PC+INKPN(V_T.3dTE++ML_IXEBLg=.3CN<2R<fU>-C)P_c.H7;UDP.2ND(\0SEaK
1-DWa;78K82V@SRN/0&K/gZ3L[K<S8S,63Q508W4bJ12dFBZ_R:9\3A7X:+LHW1^
9DL^RUIQ@bO^Zc5EeaBZ_C>bZOgM9#Hf\H<STSgYM+#MSDDY>e,=>ME/9_3(03J=
UC\MO1d(JM(J4gIE6[XB(94Z5Vg_ERGB9eK23Q6R\3V,#Z_2701Z_7FN@Pb/)66W
?M;RW6RdN)/+#<??VMSJAT:XU01&MO[X4.F9@/L5U?2TcF&g&M[QP\UY[H)[.QZW
6:.E(@@:bQ8Q>Lc83HO@/CXNVR:1QON&9:KDBTZ4FV:)=g0<DcZZ8^U0D@TTc)B&
0J3F&95,1OH:aJ1#4KJ&36,_b>b61E(W)aD2UYK^61P:BdQ(HRI,VKN2U>BB[&4-
+Uc1(ECK;VI86(5-5e+#9[E8DL]+MSY^(-2^N-9#;A;JdZFQaBY^MSSILB0:T>=2
[bZ&4=4)e8YLSPC?g1:.HJR:R0(G)N/I]fPV2W/C5<>eDfQ;6U/QfN5^2]E+8Kf7
VZ=[&E&7P6FQ^O:8dV?9ZGa^IF^@HBQ&88:2,5WXCGXd_bAG7#K2cPC,N=-R2G/F
8KJMJ,@D?c?+;]M/3S/P6)_7&?3_;P+]9\7).-(B709bI0?^Y:9NaXATJ-WbBgJL
GU4AEd@N/Z7)Te@094f,22A#+2/<3EcSLb692N\OP,E>60gQRUQ;K8[,>=<-JQM_
SJVW:JB&?^eL;LO9;K,.d?a?QR#890bf-W5RS>;eIOJDQ21XASbN?7XT>+A:gF)2
7+-HA--2.P\\[_WO+=ZQ+#&dLSA,R7Rd9]HeFKV0ZG/248/]+YQ3G6])5+:/aD#)
e0[,@_-d@>]Rd,2:S774X67WO8@aI6.;FV1BG_?&,QW\\HL[O#B^c.9[A:\dG0R]
M;<8&g170IZb+GF@^3dV47\2UFJSeJ0:B.MYK<1E:<HF7OT_HJ6^MeH]>^Z:>:MH
W;1N3.4S;eZ,Z+2QP][)a-a=:(6K<[V9&VdUe30R0<8OL@9K?cUXTKaS9TT&1N/d
^f[&UeZEPJY->?8/a^R>\TSN<ES-(DQ(DcOe4F1JfGZ(:&9Idc<98NZG/gC56HEE
a/1+?H>&&NNN.EK>W0NIE+<@9fT\dH#b&A5AG-:,M0^[C0]BEf6Z<b^[2^L60.(#
PA==8LZ^a<CAGcCO2@6=J4.Pc>L=9W6(a;J<4CO<VZAU,1RLL:VMQg=S>K^X.FeZ
&7,-],3M:A:?W]F+H??.?S&^PZDWce.>[dWA)?AKL&MeL4]\<<NEfHR#&TLMTRT1
F9aF.8#-COB@L\bPCV^GWJIW+TB5KTA\?)K1TCFf0GYLTCgJ;&B7&.BC=.\IF0^5
;]:Nd/0VRbHdMEQQ71TR8@FKOB]N-84FWD0]W;XDb=Z5.ZSG)>V=LT]2TMFYg01;
+<]XO.;YYbVbR,2_aGT]5E#&290,Qf9@,3J)&2b58#B(c@>CC<P0\[<S2#D^1QgQ
NBcEFA0Hb#W<@T8BgTYYPdB&A]&aKd@Hg8[UCQ^#(#?@?dOCLeG8:F7JM]7L[=:,
VggJWCR9>aU1S6\24(@VdZMAP<5F-N)7(dUM+V>&L3ebA.c3?/f;VO#@6,K\,?_D
>&-b1>^WL#eRK5S2OUeR)c=JS+&FIF0^fbC,-VE(;194&CL]JE9aP;RXADO>cFa5
ZKRN<g\8#5?:AK)(2\:WP^6gCJWT)D8Z8S[DJ24b.1<4>bg5LS;f1d\)3YF(]C[7
>TGRIK@g]P^e7g>ME4Ab&[?K:VT3.(H&(U#2(1^,NT0V8)eIFW7Y&+^Q3556Y/19
Y&Q#P-M.M9SBJ>@MP-)SXg#4?.UZ<fWUL>6Y8e/^X_PW;S@R4QAZP1M6O<)[bHbI
JJ.LPAfH=gf9ZII)a(&3]//B_^5GI::OBD>;),LPd]H?N-VQU-Qb0ENH[<,]RGW7
O[?M_V+J1K/._\7.Z<YA>7L9J[dd,F-/;<@L,8KeQR)+C>5Ec)\+a?LG]QaZ7QK1
LY?\/N]&^<HcS&A-Z]O4XBb+g2=0gD36,20C7=:1>99aGG:&@g8GFHR#I+U#_C7N
Y[f\(K^DGQ^UgPCB8_VQR(3]?EV6TAD3HBg_(CgcOWWM_<+<.gZ-\8=@1L/TK/d^
DBR?OU<UMWG+-CSa>3S1IT/@(/^=EU-:,SG:\9J1_);?_2.LH)WC?:CE55a([POJ
:HQ_X==Zb;V?91e@#eLU2UWUMF8=H>H6G=@@K6GU[:TJFH=X..G[>UWVWB7VTRKD
PCW2B<DO(@KV20KD^L:5=1+WP1-Q:^5IeFQQIZOJ(>4ZDfMKa>cMC_L:dBQF2a5U
\O;\S/2L(R\a^<;B;\F9.:JBg?P;^E&RKQ7?6DLQ(K#_X^92+.)f(W<ZcSb[aZ=f
NFRD7b+[Ea=eS:<bdZKP2UH7L69@GKCW9fV]?R+G;#-+-:Xaf]6C)b_dU4bDg?d/
D0c(bCeA(]1L)Ze5@(46cN2]YDc@#I<B>;)G//TCSA3f)7Wc5E7+X+aeGG<C@>]1
(0DW65&^,eSTV\6.ML,\>2bSL?[E:+b91T-06QT<]8F]P_1M9S5^g6HQL)I](X?0
Q/2)<e.&L93^P;HY<dCGa=.^/IM5#Bc20CB2N0\5=+5DOaM7R=+GC39EbSS]H^BA
D]0)\K7gg^S)6UaSD=FR:=9?MdLag3?g4aBY.P\)\ZYKe(BY&eUP,3Ob?g]C.9_d
P2=_RKA5Df)+6P7A3MQ7V<=D+[[:T7&K<XF[(Me1_9041X/UPW>[]3WX8V66(C\_
H-FRDL5]cd<S=IaVX+ID.,=Pf]PMD?4-bSaP6#T:\<>Z^&-^TAT0JIbc:B1^Y]CH
VS3c?3d8C[MSP[H&V3:Y\OATNa;gC>1T)=+eE;G_XZ@7+VFTI\Q=bP<9[@REFYa3
8^JfY^MJ#-+YC@)+2.T8\38d7F2_d(1/f8cRObET5I50[/c^C0>@=WeBO[)g0DE/
#GWU2/V1&0W-VS,Mf^(P,),]PbB#fLbIaeE(GOc.BQ\F?K7]BT\ddB(-S^ACR#BI
#KY@,G.7VA3++0OI7G5Da]I>.9N7G6,B-dV]8&g<NBB^IT.J1Q8e;V\X#;JMQA)F
O<PM@G=PcB.R1b0SR7=@HG^03_>a&Z;7>g^HSQ-)^5FU.8X1PM0IabM5]\.aO+4T
:7b0MIHNg6dK):2/IcTMe]cQaGe6X6;\IUP/dZGbB0JMBU,45RH;.1g1GaDLI3G-
TFO^<R)\1NRL(>IC_F-/W1O^X44?D@,^_G7B=@N.8d=8P<A(LXcO=:(=#?-&^KWJ
0HN=<g;7E@;E8V3KJ;;e_W[(=UCCB/9==fUMX@g<[fIE)gdA#-LDXR>KDOP/Y.,D
@K@Y(f;(bRT3]Fe4>7LdKg#KfPXM?(M;6BRB-52&A@/-[b+/M6])=.>&HH::=eUQ
:C@6FYY>7?IMJQ\._FS4>#O?@+bQWe4ZeK(UY/13.RO=T:LG::DR+]..L.O74YdQ
[L=PB;/,7DB6(K(3P,,X=-HUCJPBd3;DMBa9VF&5&&U<5[+0AH0C+1Df(?:;30be
J#/L2K;,OB;C7FG5Z+&+6(V^.X]?TSXNX5cf#Igg_]FH.2C6XJW[L/b0#R&2?(3U
_OWb\PFTE#[Dgf(-aL2T0J&L,P\FA?HPC[1R[2=VbD/@92,0-<6Q8d-:&ZEKIAL^
JU+fN_J@(&/=@VYf[6P7,L:9KKHB[6=JfP;VJAcV.4c0RO9H4X5Geb),#.&WY+R8
f\-+,Q\[aY\M[[/TA0W^=KK=^AY-FaZ<P@D[OW<^:C3V,M370f;X=(C>54Lc@W1V
:X+<MbD1;JL1/ZDAJ?V,OL;IYd-<_,d4_KVAERX_b/ED;=1)>e21R24LZY8X.KXU
2c.Y2-];XW_,>&dT^Z,/)M7[L?YR6gB>;O(JE9+B@J[W_)Q5)1^HTW(ZRTbHee88
F[5/c(f^?]g1_EbC(SRd2W42-[7QF\^\^[KM1T5HN<<;1<f;^e+FS&c=.^B,NX3B
G92TH?JE+@(VL_95:WNe0&<cK:fK4-FJ>5Sb+4T1RUH3.KH2]21G>_Cf5;OMdRR1
A,GJRNGO-M9GCLPaa;0A.,1V3af3@VR5a7R<[E))4/YX&&[YMFc88>OWJ?<Gb3T6
+=^aY/<K]cO)K96LA(=db+ZdfCbNaJ+DQ)/H]B)-R39?e-A1TH?EN&c0OIWUH[22
+P26gP:3T;(-<ADDP0+7G3R(a&DST+#@L>&UZdS8;,eQ5<E<KZ([^VFOH+.ASU)W
.O2KKKTOWMXX,DP4KbY^\3FbH+III9,D/^77;0XATA,5]g5=P_U4N?=[D,#EBGT/
GB(@YCB_+/(9P\GP6G@5.Ea+E@JUXg146^)6\a994a[2c+T;_Y4cS2.P=g.HW_dI
E76KR&G_.RFZ@HU^21fZVJFI7;X::)B+7K@>IS2)2MNY?BB1=g,a[f+1Z&[I?Fg:
L2;>U]f0I[7?7:&g)c;EKce;K2(BdV@\V_M;O1C>A:P^?AV.R/Tc,_SV?Db9.+Y@
<WJg=ZRD8f[,SRbO4^F62GN<<LcH6;@UXUU/7<W/?Neg=GeQDX6W96ITEL@Nd]-g
;Leg5/->@(<dHa/CeSV.]D-B1cCEZCYZO)I+W566WRcXaN9UfdX9,dP9/5@Jf\#H
M,<S>^RQ),dT9eR#SZb[Y\HaK&HS?f5J4VC5DPAP@,0O12V>)F-:#+^0G#3)587W
4<HS+cf<[AZKW6&\J@WWU^4OSB(:)LZ4QW&:cQg1_FF_<0C--dg9DR)L11<.(W@^
FBJ(e?N(&71XQ_9TLEVRV&I7J#\/b]@cD/L,D8Z<e_^N+&-]/fHELOON<36dV<MK
CQS0+BeYEc=4?@DJYFN?RLJ\KY\B-SEY,D1RBC1]\H8]TM7O/.9_)ECH3MVL)W]e
5W\&3.PF#@VQ]P>?YS=LfZVP;X7HI8<Q>?c9JA(FbW:5)ME=EV6IT&PQK]ZJ?55/
aN+gO.CJ6#0Jc]]?^?<Y/8X0AM:e^1d/FQCI-R6fDAfFI&SfAMM+G>I-;.3<LOS\
[^31GbYX+fL531dM0WV7dEBN>d;>^1<e5e5-dG87V=/T>PP;>R)g5[M];GBSY\@U
<#9H1SYWM^BMI3WO^feCZR\0&VRL][-0.b>(]-11J8-I\LGa4K5\QZ.f0:H=.AK2
[>\.^8T.Y&F63Yf?)(7<,<Bf.aQ,Sf9AB\dIfUUCa&VOb\D[3RfDVP9_>L3&Pf>^
R)Fd,=4D&5^;Ud.U;cB]Hb#V#YQ.YPN.O05Q4FF+9L<]TGQRTB\/:^O#M=2E/3b]
Tfe&BJ4<VWP.OG=XV>;J+8&61\]8-PWIN&WK,YQH)+81?&gAM7A1]H0^D>FW5>Qa
eH@A#Q_0DeCH(SA3[/T(eX4YT?#XcA+?:J43V0W7?<Pg2MBAFR4L0PF.L>HbL3,<
K>OJ;2efJ#a@VF=K-&VC3GYSg)&8]dI]6CN4)8c68J/cYVV84T1&JCV].:TK@[Z&
WBJY)3Y#D7.-)?L+BfPAW=Dc2>)UU\B)Ld]?M9^3&Z]_:fXaMD;HSU>bNXe<U7PS
Y?NF,cF;?K&Q0:;6N2F-^Q,U-Ig\-O->(PF#I3TU6^:?,dTeX,5HH_HMEE?..QbQ
fFF:H;[f>I>)UTLFg4\8ZP-8d&&E?,,(NYJ3=PMDKfVE-02NQfWf8@;b]H@Z&)VY
=I;gaA<5dbAHIU_=-U_II(>P9QQ18UB72ESfNGSaOR7RR-U]A4B)Ma<F#&=dDP^\
EUP:4I2S_C3E[^(<#CGfBRKX<).)1K?-dWNG149^_XU7EFZ\T;;2.P?g_O0B0QG?
E&X5PR[bC;C(]_^)fg+R.4eDAB<)^O7+2)<+>SL=T;/6GE^LSe?CRaRdV;[-;_X0
W+W)3=2@,H.I(<2FEDX29KQO;BfE7RVfcKWAU?1H=\RV0DV2CJE5gI>TA,\Y0+(G
6X\2K@5JBXOB3JB<2--@J+R\(:2GE9?ND80]O]C.3329?5\>7RT>#M131#671XT?
(4_VJL42E9>(ZC6MVb6U<DUL>-9C\c8..J49W(WE^GW]4V]P@F]XURM,;4UCMagZ
:3\^BRW1gd50?Fba#9,F#T-+&#H94\=F2Yfa2eL(e5aIF^^29[BeT)5CV&G3F=LE
NA(K+KB&(0VSB>5d9^Jd/57W/6_fJXCZ7QVY,BBNgN6V]0)79G838d6ZXG@Y_gCN
[9b_3,^MDC.RFNG>VXO36?L-<FMN+7Lb,NH+gLeNM\<M[Kb/#a<?8Tbb5[Z/cBdf
Y_;[b+OfZ+ZQ:;K[_M=6):JQWE5NAOAK.S.SY^63U-FE@;I;D)PAeV,((/.&BgBG
K_V#AK&;)PK.U,NdVUT\Y;X4\<?[G^/fSR.E8=?d;WT)@.G,J)[2NPO<;F0.\b=c
]08L;#@W731-[VZ8MJ5A44PF\@9fSP/.8,>M:(Dg8d=FB/THHF=]G:^db^#@McSX
egb(V@T:Ha3NY0V-LcdQ7a]JSg693gFT:+:#6fKHX()XDZ_-2<M)E^-<(:PLeA43
8)S0d_-fRO<B]dAG54Y^+M3WE#Jf=/?0NY(Mc[BN[>4d&@Y.3)V\(#<V.OWOBROA
>[@CdX^EJQ[,3.7R/[(9/#g666,?AK<9S6fUF6L&=NS7KF&FBCDc16&S>[JSWKO-
V.,F]^>5c6;HKIVJA\=^^WL0[EE&[48>\NO(EbKA(03ZYM\E5+JM,Ne##VG+,_F=
YQ3YR@>25C?+FOW)?\-@+F+FP7-E#++W<(YK/f\:PC?J^ID1XPT4G\T\OREBAUg#
;@2QU;3:-]:^=9B5RCEdR#L8bUVc;GYZ?0G-G:KMZ[QMgb;UeS()C+[68O.Z+>OB
M:VCE12NfA@97\3c&X<Y>O3,UKN1[@Y[TdXF)FdICIK:Wg@X#M:<4?Tb4\4F-+J[
\GYBGcW+=UdS8fPOI5cZdeQ@E&6;@DK.\K)\@[OJ;.aS3?,;XIf=N&-;0JL18.8Z
FZJ./,cdJ7KSFT54cbd6+>NWR0A\=##gOEN26aI2E8EYXP)JdY49)fBH&0B]RSTS
CH3492_>?O#gdW#E+.g,+Y#d.?0J^=8?QD8HD)^B\d1H54C\=+f9;]-FT\8E9D_=
\V:^=CP@Wf1:WaHJ-G6#L+dCNNK0MYIZYCI(BF&.bKVScYdM:7;UFM#HbA_ZRX0#
bbg[#&Eg&dKSOJROPW;Gc_4Pge:F9)M6);g9aEeVMS@AQKc(HJAL3\S7A4/XcQV8
A<8=dPT9.#9BA&,V2=Y;QH^A=Lc3+?/]SJ;QWZ9Yde0\30MP\B[U7fAMF5\:/cQ+
#MaAX_?4\-?>eBFO847_@DWR&<MI:DabLd45T.^QNSA-6]+90c60Q2]+]EXQ+D7N
/dIJN]Fc9(X]?\E)6E_R5#YgH0cGObgZV/Z5Y6<#)Z[@Je+=]Z35a@bH-b1FTD@:
cT0DAHIXJXBLFBUQ(^2Y=;0.N)fGLbAII:I#Bbd)2^=>BOO/=[W>W)cE25&[Te;R
[E/JfP^@T5a5YT/-7:(?\aU(K6HX4bL0e&.B4UEUaSA1VDJ9D)6(^=W]Ig2>:NKL
Xc@N=2T:/?FI_cC/c;RF4@T,;Tbe:H_U@I,g.R;JFV^V:e&LXReZWC7)W_)CO<e-
O^R=(,7,&W?V&<FD+2:fFbJORE5K;D6:,[0\VJA?g4->+>f@f)^)dGT)]:MScgR2
X5/7;U>&Q4ZfGg1,=3GE@HMcDEIP^W<\fAA1V5_+&VNTa.J+64VBBbJLdAV^;8C.
,Q--G7&-.\OT2<ZV-E]I?fd1?8G[?B#0bC-?PWIV)_:RKTU/,fLKXIVTI95KK>44
+d[2_;>]9A?eA2]3L6,KH2R/)IZZ]L)I<b3E?;ZV6QKTT@.]T.^M_/ZW/1Y12OKF
>JYd3L^]8YT(T^S6V=F[:JI^gVJX6.R6S)X2];Z8V[cGaFIQU9aU;@5W0cR:B@1e
d.>#?8CF8:L=36Lf<RFJW3eY\_6aT4^.d=TMLS5ZV>D:H]c;GTMYZW]g<&MJJ()6
V#b>Y&DX7WVg_cOV^E3ZF&Y@Yg@2KZ]W0.dVB.<X495<_CB0F/&\GI<[\X7]9fQV
7,KQ?<I)RSMQW?QecHUe5g[O_8B-BMLRAc\AQ(.cd9g6.AFSIaYbbH=S6S.bYg4H
c54,3NURT&c_)1=Z;0\S59@<XV;JP.LD/.0^N^WLL\,c6&abFR<OU.0A&5)^[8(b
649&]Y9e7435cF=#:c>P0^a@ZAT<B2=#WQ]MB@56M/+8MB=eP:&IHA>P:+12JI<O
a)3-c4>L:1.aYdN&YdWb5U\cVOHW)M<L)Ag;dF+UQ1U0bA303/O4L\PIZ-4Y]?gW
/8<N7aX99OPFc>aS5-<7;XT;[J?#b[LSE^g[I_Z7STF/I^N(?Y(1\SDQ^,6OXYQY
J:YAWY3<cQ><[Yb0Kf/Sf729T(I+a7/>Pd9T6JOg>6LP:\=bBb_g.P5S96AYT,:S
U6eB@R,D8+;.AE7Yf3BMg&77>2?N1S9;a.1?,?,V@)8.T)L@Z)dM]^/YXD0SCBf>
cL?;52&XBg7<_PLB&O&Le.=:L0+6^4BA^ADVaLOE_++c6VLa00-:/?,H0]2)_(cM
B8,_PSVPN.<)VaVFJ-RQd(FUE3CDQQaGF4V<GX2#3@RK(:+,eS+fFU38a:&+_BcF
U1S9?GN:UV[CYNfL<3+6c]GR)^<E?N[<?ROdP3U-#RbK>A=<Ke1e7X[X>2:].O;S
;UI_59\bPAb.3-5b_\V/F>.AV+0VPP,(Yb)BTHQFfE^NEZ<&_CCUH&B&c6(ATRHd
:&2?QHA6G+V#7Y8c2LYT(\KN4_1(M&(db;Xf82M\XLc7VQB5.(Y7X\+EYH-(S9@E
G0Ca@&dL3A7EM]Dc1bb]MQG,EMLebS);)][/EY(,]IC_e1=H#+aF0]_C6)<&CP<e
N#;7(HDc_CW15GfK#;(;CA,gI4aYS\CGM@-BGW7AHHDFH[761T]<I2eb=aLPRe,]
;F9EaBSM)1906G=P8<3QU2<W]8@cVMF_PeV(>L-BLM48]c?PFAA#I^H?.>b2FT2>
)SLfd>3W,]_V;VSQ\@]=/U;+]SBc<IcXaP<K<H/&_B2V+8c7^_FTYPMVDR9P6W:P
PJ+Q&.UH(YdVPb+L<JYWGJ9+JZL+bXa/V&SH,)T[^DPe@XG5bUF^@/+S0W4MaaPd
G.d7\CW0dCY69,COfb-=H>LO_-Z^F@aH83_NgO-I>R4&&DDN-5,d49(Re[@7[Y(^
BJbEd-d29NYEXFC/aac0\\,:<9D=a+08F@eO&E:^I.6#R#@;d?b=Z(dLQbLNe\J8
(T,D6K3IYL31#5>bc\C2DFA(:?Be-Y3PJ9@)R3>=e6ZgBVG1J:D2+eUgNX<-Ucgc
=27PJ=RSO8__b1d7Wa_)=cF:QRgX<Ld[NTe7g8eb^Z5W8/K+[U\UV;5CV4#^>MG-
WG2eMR9O.T#ALNKWAKbNSZI@g=c:@]AGL0=;?MIG0]Cf&)VAGD07C?dEPe(,DP<T
T1KZ.^^KMg+R/H/8T@MR2<gZ5D]\&)D,)N^?4Xag+^+a_@E[_V,2R?c7[A1(\^Ja
-_DeAJ2(5]3M.7N2c6/0;daJa_>DCUO-fE0&HOBcb)4.;IU;KdPA0TR6d])VaGC,
\TcSaZW2+,JN?0aP&@ON?:2V5YEE.K):AJK]90?&c742Ge)NW:W2:K6W0F\L9eR8
UMfVHZT^J5XfD2a#=3;:(+\eBY+);\7U[\^HY)PCCgXANKdV?I5UFNI7V6;MPa#D
)U3HM0[ML6F;SEfL7<.L-(bITF\R94Y)1Oeag/Da9EC45XNdK5cGSd\USFY=&aMR
0SK#ET0H184-:>7>AY1D[[T2d>\[K\b:=dQ46;[9[S(8[e2UQ47K2eZMIBIMcg1O
7aC1ae^ccg_N]7;)\g6_YK)/F]7U?aY6bK2X6db?d)TQR2dSKTOIE8#@>1);S88=
[Y^U0[DP959#JE2;FSO^7?Z;;2N_,M5D&1>c<S7P[U>>)+@UdcU[H#fZJC_Y_99H
7.E(E@KI4GS:ONCRW]O8RZNZIa04gaA_8J3RGgFU[W(7L\-9O5M34C_e,4Ec>;+_
81F:XZ]Q0RgcJ.6cV(U/&aB9Fc<0^0K7@f:c4JT6Lg_FGUL;I3ZH.DEJb\Ca/:IY
@EY<6M]/9BF_1c>BAKMN::5G@,2?^G&+?/<gEaIFeB[(BD/QP)>\MYU>5,IQC5IT
@Q,VOV>Q3.K=+Oe7H\[6G</F4c>(/g>1MTN\e[DZB[B4=X9I\4:BUf;6@N:gOVXO
^)(ZU3-E(=[#eb-Re0H18).7d?Ec^[NXS,/D8JYQX4ad..?:VKX,5e>1PF5=M7@>
H/c>ZgYZeEL]/Lf+HBbE?a&f8f\3Y5:f\>&2L7;N=c-9?eWGV2Cd5dCWHJT+H8X]
FZ@93g2(HC?cKW5R7Oa?CWX),\(T-(7Fb.VO[bL,2Q7Y/2]V/F:P9:Xa(8Nc<0,M
V^&@H2f3Z5NZRK1dN4-^L@QP.S3X?Q4b?KaO_<[)g/BfdK.CBY^?#)?76Q5-fg8L
@BF2_Rd)RU_WHX7IUA=0/C?]H_F.=T_.Aa5DLRR]cG5)C29CEg3_A?b8+<2Uc=dP
JOE6(BK((>RH-)/9>S)<AV^60G)_+>E@GZb,:B.SM>BVU;d+#>6(4Y6G4ES9MI;D
G=4NcMG_e\,e#?dFH=YY07eGFC#.4a0c80(VaVGMKe#:#&R)-@b@C,5NCX(TY1]Y
H&1e5-D4_7_BHL>B0RH6,b+R0d;+f_E>869ET[><;0_L-NY?,O(FPX9fbZ15#g_Y
gQT.BbXR2+4<B_(6Q;7HZK]0>XCeNQIPP6&@J<VD3?Q^WP79aR]JFf0fEQP+A33;
f9]44,A8=?(RV?5]FBB)O-#0\gRA7Bd3b?SOP45M>)gcb:-;W220_H:\d+L9H62:
H#_)A&]V@A<:\#]MRJJ2]fU=58:dO>P^U_+-a0@S16+5^E:bKQ_ING#4e]F]5Cb-
D+7I@?^/#Z>8N&LYBF<H)5?.@=@OXebL7Q_HSZTY_I_EP/4eE-]S2=,S8^-)68&=
>BSDMDf5QZSGI(+beK@;,29J0e47(W5GP48\P?aEa71#bQFc/ED<FBI8H.6f>T\D
(:WZ:9N)7FZ?<92^QQND<&[0/g++M_RFE<@#TUZ)#6VecNV)^W;&08/4NI-2:YN5
#[@g4<)1M4\@[;;6IR]FHMY^fUL+.(OIDc+5M<;A1=1B?>]g)S0Y__Z[YSIONY>]
HX/#FSBFQNVA_0=aTTAaBP^^e?-=T)\=g^D0>(8Bc2PHMDCJ-YIW/WX9S28]cOXc
#e^QdYgaS3TR1@4L4?/\UG>UR#f9DUQ;4N>4gcD4^<AC5+DAQCB>fa7:C++<^>U=
VHIc@U:ZY3LU@EK3:;c37J5X-GcRING3,]SI/K#TTEg_FAM-a,L_Ng0@4?YC/e8A
FJT1a5/NdQ=d4=)9M,,7A(33^#QX/4Ac[BVC[[=IU68BV_U#YE_.XIPB5MQL4D<Q
H-eeOR7&ET;E9<ABL<6JCMJ[@35:.7D[.Qb8U3LY2.O?De0NA\d&;8ZcHG0)eT2[
NK;:PUAEfUZ&W()RO6E)-H81;(D\95eW#LN3UfSceIb@:EZZPeVQ[_THPcDSC,^>
FN9QLQSC+:\((ZdXb;a2L-?7,58-6V04)?f#6T58b77QE/TAg[7>UKF>9=U8cVY/
g=Z_,#NJ=KRB]3.??0_cb8&-(c)EH4NE90a73E0B)/-4XP@Z^,6eEU3;^P/?GZ3P
BcGbM#0Da6O)6CXH7V]M6@)bH^F]#bE:A.KVM,H[&_Z^N0?\O/&U7V8EI(578,:R
c:Pf07SMOe00/9R[L2F_cS@T]Ta8Q3RHG8W&(.)+\_Z24ecX\/6c.P(WbKg<0+BY
UWO8[>6C)D:)C(3&(MT;;>(I@dI\,Q8GRL2ISPVaBCF;S)BK4=f?1.K0AAFe?Ca:
FW,O7=8PbQSS8L##\]<R4a+G<;7<>a>3(/6&aVf)^LXfaX7T:HVJCWA^=aJA7160
5DQ-WY3A+>1ZC[D:-NN\4,;3SID,+(,=4LFKac5\)Y53f5:[Lg->(4SWc;A/E]]B
V+eQNQUR)/5Y:T0I-aK(Q38cJTcD4.cQ>A\gEgP#f#_f7aF3X#]Z=E52YS,:4R.D
R-1L;2\^V<WL/Vb+dZBN-0O-1^J:-G,8T+(6O0&6?/4\/LFSbXLKXJ=(^#bL]_59
f.CR?OE-c=XFQ2KO^VB_U>Z::.?OJG]0(84-aX7W6<P:GMC,X;P.<YK(9(4N(g;#
M+MCF]L8=>)+LU=#e2NbHF:8STdREg6MZBLGY#:cC1C.N19@W-OFDN[^G3/8]0b5
<E0:@74BG@JRNIJ9<#B0T-H4Fa7Qg0=dNNIY<U?EVWTLdc;Fb1M,eO.^Pe0W7dFA
/Qa)eR[7YCAcM+([DI&MJ.cA=8_dU\-^B4EUI?NM<](E4fTO9Y#YVIC9;<UEU\?K
NNbCC6XI)P@/9K-XWPf-A&GKJ?bV@2_AQ-a.8g,G@5d3Xf0MXJ7abVaL3CH/)Mab
-+9Q6]PLbVEWS71egaL#]f;DD8&VR#[O(=2^d^\;=eBORb?ERaY&5VMVQH<9JXcK
D&:7c29H7D@faUDX1\2([--\;7H7WT&,ac_Xf:ZZKP>.0(c0J,=F@e[CW4P51PZE
E@Z1G;2=3:f40+6VY&=)<+4[31A&O;ZFd:A\BI4#KIAEL3W0:AKC(M2F)Of7F7J:
:-_Z^J\5\,)K]aYK)LE5C7[7=<]-3OS@S/EfAZD<^I0(Vg?:g\aYCH3P?c//+^(G
[>cMTLLCFK+E+QfY1^W&=6@<^7B16G+BV</JQ+MZ4W(=>1X5PCU)/V:9Ud>DK(98
E0:BdJ:fS1WR<K:,HE#;W5LZE/,IGUPG&dEMK8dR,(RJ\RBOVaZ@&6?UKJAJPQXe
F\V206/4YWJ)UOO]K=CE=G4b=T[LOO<;3)]L;NX.01]L?UKN?E2),BN(XF>eIYG?
)_&G.HWf[2d&OabL>Z@GZ_EKN[f+DccGB3#L\L_?>e1QL0I6_GYW-@3A7L;#MW#8
5M5X=JeWH]V[c-Z9PM(ZI&SA]Wab9>[\TY9JJX_)B.Lb9]5Z#1K6ZDGY88[]AKBW
J-<.S#\P<L?0:dMWOG8].a(.(_gBMUd>1QU9/.McWEO&.,<g&K(Xef&#?[^O;:5W
dPMVF)/)YZ56.[OH6cA5Z^JG[\7HgW^5Cc5c<e-U;+@W[aL8:S7RK:2074:EC(B&
IJ/2)d31cdQ+>(]cdO2ZYUW+VCFc3W3Yb2:39P-^@e,/GVaafXJA#U;C@-T[YK0P
428S(;Rf3;@T0QEO(;[O6D;2P3dX6+gWW@\FE0Z#c&TfRb6a;:0OV3.C(H-=Q&@Z
\(C(RJK?[.R_VYCd9;,29LbW&cfE/6T#]X.,T\/2NBVa>^2S.Zb6:K1,Z4S?41IV
.SAWXUB=.(G7I)P3D>[cL8&DO2\IF(Y)+NaeG;.;MeL[5J-\5bOY=b=OA9;:N7;4
=MH.(W9[V(X&YU36N),I)XUFUU7)PE1]F80MXf-J55SC#GVR,<=A?WgLdGeT9.AL
2\0G;UYa1TbYEG66I:<#V[T7?20^9#LYdHP?KO)D#<1Z=.G4^CLfd#\[Y8DaPX_1
>2DI8#>,+<K<A7UbMcIA<WgP-=5I<@@/B9#BF9#cYb6cBB,]^&E3(>MfJ)c9F6W,
+J>77_dGSb5_+F0HM^4=/d8-NX4eO)b.g>OM\[:P,=^C]W_W=,GdeK_T3#ZeZ=3[
V:+F8K?OWfI&AD>VMC>Lg,;C51>K5G\5[8>]+<O[N1B6b@B\KQQ;-Md:;f,(WN(>
[AD.63WFd2D-R#IC6R58.@6>HcPc@6>&J-4F]IeD@ZX[QYZ^LaV67gM]g((6EIGY
SW:MaV1-C/VeCfBXBP,;[2<_R-S=@<4]UQ-<a^f)OOG2da,^B0#(X[AVWH9YA6SE
45\UHJb,d_1C^5A>Ob(/BP+)Jc,>TL)4)/C6<XO6^ZNL[)Le)MFV,[E+N[?YD^>\
6^9GZH0FeTbF+_DEJPNgD/#,=gKSGXa/^-1Mba].&10eK/GAUg1A0]G&N^Z]<NIW
<GdG:)TY5Z-1CYd0Hf.-KHVcEe-H&-Z.G\b=WZ:TKZSUHXg2XXI/0JI.R0G+^=MH
f>D;(9,&e[3F]a=)9:IQ996\^5E/_e<C-=A_8WAgR,0)IfCYGJ<+2)SbP#aP7baV
/0/+5IR)3K..g,.AQSO@W\H8[+@GOXPdb&dX&BDTN^W]7VacW;J?HN9#HVD,g.cG
O11BL+-BNLM56E=bY]O)G7BF+7G<W4HH<:Y\]T5C\K1.F3[_UBOU5PQAJ>LAM6OH
aN7S230[H&@_E.eedgQ2V/TEgUQ(:Lae8:,,&3=/M]#W2cR6C49SOS\^SFQ.<<@f
6M/BA@7N;HA<G0<^/HIf#HR:d6F\cU@\YST,OW\@fcEMFefM,_7e2RR^MFZR>T<H
+;Y4L[<A0Z6Y_DV_1&VUBSCA^TeB-Z-H@_74X7bJ_O=,M#[6(LD1D-=#bU0LNWfD
a.TfAf:ZdPMfdVFE)@WB>)@<Y2PA72d1f^bT@0<<X>G]9SR-.)J.5aN&D8S+ad4A
Ag8f;0K@6a;X\IgW5^=G9\5DSd_@L[>aG,@,b7JW6W<6TZ[I3YB(3D_0[e?@c5cV
4E2g[U\cR6Cd1#V;\CZ\:W8NM5CQ\V&RSE]H^/932c3?@E3[>:YB<gI>8=:QZ#_@
gAa\0)Z3\bg)Pf6-=7@\aN0]=9]B=&/fg0ZbaSNVfYCDgF^M[cKbOG#A2X<bC)ge
+PQ>-00;HAL]S,cHSNO).23H+69@/aC9FXRUE3f/,daRE]K8[#e65RZ(R&>cWW;?
bI=Q7dU//V9]9IZd8K4Z6D:eYG53]EDNI]52cb_W&M&R5e8YcbL=_/bCAZR&G1[.
Xb^A<bO/U?cMY;QA;QCONI\NYZP&S.>cBK\@^K3C-@F?79/&SU9g:NHNEZ@/EV(^
N1CFa27e7LS/EBYFDg6:1]NPNW[V9@fa=W0IE^W5Pb=S9FD)P1^XXG@PCD;4#g:<
0;FGU5+#:RZ8.c_6E53&&)NaOcB>J_+TLC#>9_I-(J2bPOZAH<7EL-60+Y<WCF0(
OA9c:JY#^&.#56VX8NCaDaa41]SF6@@1U_.1=QGW\:P=Uc7JC[(WafU7XF@/(K]X
^MUL2bFOFO-^.NS@3&;I4IX-f:(NF;NWACP\=DZKLbUABHDEgJ,XK2[+72LXL7T9
]3]H^OJFD14)H@9MG+4?,CV#7Ne;>C]8@ODG.E43&\;NIC-e^??TSbJ7JPaYRL11
#YPL8EY2ZOb;V1G2;AQTU_gF&H6UH3(X/J]E>L5(5+9<V=cPE>:.?aZAM;N4]e3H
Y&IMcBX#4[P.F(;32&7M/IK762C]&K>?+HD@/a1^.0;ZgL-1[fb59R.DQ;V+1fU0
1P=Q[UeFW0O8#Y4(.5)LF^E4X8_<R>JeMK)R].4Y-bY/X3L>(?7^P)@A1W=J,664
V]#A_2Q6cOQ8eH(TWI72c=ZI)4\2>FHeC6Z^I5-bd4GSP)2E.KK-ebeME4W?CAL,
L#edCOT??5J;I:2\USd7>@DR/@0dF0ZS2UH/:\.TKJLb.3?]^2d6U&J\DHDdL:83
_R2?-2754aA1BPBP3J+\.\a35)7([O9eF_8;U->PgFXPVG=662b)#F&P.8IBfNQa
0A-BFW]R\SN\:AfG2R(C^>U<,&<M;JC=@5,IRQC&AS3b5HFa-O<28.[]fS3]FCZ\
#3.b7@Z4\^Y0T?e^X^QW/-DSa>a#C9OO#5\@EGAD^eQ(^7e[#RR+913,:MP3c>Vg
:TZ/55<A/XR^U-9Ha_V@?K,1LHC6aP0R1b?B9U7]Y[WAO5^KN[[A4,([GN?5].PA
#+22MU<,U9gLa-Y1-N_=1YGOHSN@QH]F_\WA:E()E3GZSaNEbPa#bVb(acD<.SRR
&9RfZ[ILCcHFXDEAK6+I3-BM=FO91@81@H&TAJ[XdH_8R3(DMCO:H&09-N0-b^5Y
TfcdMLN7M<BAY&Rge(Sb&C0P5-0\(?)CPE&]-[Z&W6TBQR>8OK:P>;>.GB<Zc9N-
]^g5+:L-@NS=aA.DNP?e.\C-.MX6@..W402@U5[+QfI/e(+PDV[;X9^J7e3Pe7YO
IBSWU3C&3a@bb6#2#9&B;)GbP&&S@R=NPU.)=J^Nf<:=CZ5Z[QPbHN9V9#O/JQLH
<8IC/@g?#c06R0Ee0ZX,QZL)Ye>X9-V]K+-]+_5G2<7AFNb;-9\S6#8(b31fMJNJ
9F86Z+W(92X4MVD_?\aN<VM0<HX.d7K+U9b&Z^ZU3/<EQXM+];31^(P1/U#K8]f4
LE#6E:bDC5,7H<#Xc3>3?1B^7b>RHCI;@LYSRFTdTKLI;0BQd4e3?.agL1)JP:DS
8#.;-OU,.+>FN5e:C):/&W+fEGLA,ccG(CS#aMXTf&6.H1BEU.0/WdTH1?QL:Rf3
VUZZS>.d-S+;2E&0Qb/C+BW35.A-;#)UX-dgYbdQI?+;OF.:<_;D?@^CB5@O+/R5
g0&GfTJ5C48(-N6N(2[0:1\W/U>bd\?>+X-]>4E9M?P:Y0NLUJ<-VTge7>YR+#=5
K)bH(0eE.E(ZE7SY3HJQN<e/CJQ@?+,>)PTOL-IS_>G&CE5,#IgM1aQ/Mc8.QFYb
E3dL<+?(fS=d)8bL_J>G@#;TJ?Q+>J@dB7bgZ-AJ@Tb4BW@E__A6[?_G4?P@JLG#
OA=MH(PNb-e/8G/MC&PQW&36,HaLJZ?8N@AXMOPfC(HLK6,^A5^._>\E[7SH5TR^
c_d.<@dO5MEaS-T.3NAI/Y;d-(JDBP[E:<:ALT1b:K6Pae<;5QW(Y-9GF=:FK7;M
HQPO+Mc_FeGc]N\3(\<PK&2W_RB2:GO0G\b9BLW6AA<GEaeSM7:=E\8#)3+1Q>dG
4.CAPR#5;-?4-2UAcI0I<bZ3&(T(UM1()^1K>?O..2B5JMX;CJARcK)5+B:1)F89
([\=^VQg\0;@5R=?Z\-6]e+ZXRKg?#Gd5]Y,6Z8)U\[HJS6Lb/0E,eI]&Q-g)C@M
<2\4D77B\?F#4D6CMHX6<Y?1CR@?TH5Lc;b4>V2IG(I(;aD6?THC;1)OLK[]d_>I
,[O\P.gb_7?(/d+_.A#V,9/CI60&+cf;^X?O>@])SCX>OfT0A;:g3&RZdgU4=fT?
Z3,R7,-cI0<d)#&f3HPQ^5W?G-9394<]3&L8R95MbJ3OG/B3,gR.;A/>ET2GeM;-
YND6Wc;O0:K1T>B/P[9d[;4dc8#0G9LcKQ2RJ1<[g<\GIc?.\7PH5?:+^TB#<]c3
V)VU^M9Rb8>g@W\>)#MRBN9eg:0:KXA?P@3WPAbcNTIPZg7G\&,MDGaUa#EKIeGf
+89+0Z1TEU(1Q4^(#X&/&;)N=0VLBD;HW<\((B]?<NHe#ASQ[##\8@eUe[NQg)(G
V?<EN/9):OQ8C/8(3Z/R2YV]B,D<gTU>0CNa^XVBWC,X4#;2J&UgY0V61O66=Pd_
A/b>Q,P]O)DgTX_MO1)fHM#=[CNE,+A,eG7<D2Z#P(K/,Df,9/[#O@;D7+,>B1K(
[&TIE:gXM[UH9Z>NII?#=Qa<2;PJ)YGQ]]/#R;L=CV?05(ETSNPB1C/4&Hg2b-IS
Z>N1C&,V^.MH/FT+NLA,/125CQO&@g]A>KV.34FKaVY?]_F:<)/8\EJfU?a\FBE;
HU3XS#RaB?E&)&[;F)W4Z/#:+fT#;1H>4)aL)GB7K_dW>Ag10H\QMG_&<d,eO0HG
ER0\fJS/A2#1/-^AfKd^gQ>)(7K3QBOC7?5MgO3\60W:<70=>M,6__YR2]&8Y#P:
aC^6NY+fRc,_,IfEcbQ/g9a9@VT2L])-OQe0+/.dHDB-7>g)43a7-9gDH8Rb8,>b
348<0-6&9HcYRWAfSVX5[Q,8)-9JW<gM;O7R^Z/5;P)@E[?ETM7\?]\7:d3/ATS#
QDfMG_]N:4gac1eD?>F=M6eLKVC41(caZ,=+X<&X^D;QLJ]UHB85F@[Wff\+_=.1
9g+BDHK5=?FH9IR36eCB2D#1f56Z#dX7)M2fD[4>5]=Xg)DRT,EV8?TUcfPX6M2@
>G7V5dJ\Y];41HC?5_bI;7g,/F>G_2d;-5IcS#(F><A^_,H6bO;R_D9KL<7^(R)G
7PXUX]?[W@:,1DC/KRL?5DC>/Q?8#(g#Y;ad+(3cB;X-&MCbMZ]CBMDYS#8<;AC5
EFcQcXA.4&=fR,a]6KTYORS[#a;W66I4:5>+&f1^,W.MCQZ-DN1:.SXdI(DIFW(K
54HbRJfW:2>aF>M1>&M=>-+7P72NH9c;F=gYT5.^@.0_/59bNA[]:Pb:/_FD?Y#R
1b]MC)RE#L8LL5Q=5@2]TL&XaF0^eF@9Y=[/L/4DG@I#70=_PdK\3dR<W>5@3.A;
4c>)Cg@2-;M<0W)&RTA/6=b(&4>3FFa5KJ4C<?-A((9.[H>301:EC3N]JKCYY5UH
D4NK8d7CN=XKQOF:PF;8M=_QHY@FZXO#5eFI;&WO89=?]UF>;H#GgB&MA8=9Wa_.
D@F/eI10QQ[57ZcF[MJA,D3-9Y51&\W<dN_d;e)O@Z1>R163ggEFKD/Q^KIe9eUK
JN_cg90eW?:bEF;L)_CcT/-_OA7AIN^S>^9ZdKE;=NJ54Z2F.>2.0=P>EU0FK(g<
8,J&JX@=PX;(5aa1M7W<CR9++47(17DcE<)Y:Df2U&X,W7dB;Y26IG-F+3/AfQ9>
P/7&Z-R@:SE^C02^X&bIYL]IAJ-^Z910g<(KH0##J&4dM5AU&M>2H=(f0V5(Ud8[
)9P1&5(fVbg.E27GUBS[TM(VH+f2#/ZP_DIL.8)NV0\?:1?9F)H[\V=6_f[AXQ:O
e>?#fU#V2NLC;=PTH\WCIHg+RW3AQQ)BLL3Sd-V1E?X^+:&]E>H8Z0K#?c5;aWU&
3PP&^g#?PSN5TSRV08]LARW1c:7HTdCEFV73Fb;-dfJ_f:;ZD+2=V:1,J;_XcVE5
MbX0EeGHOT.aKHOgN+Q?4RSYNeIM]I6&WF8;J45QA?_O&7(Pg0)-[3g)5F^ZKQD>
ZK(/5V]?4_<bI?0Y;efFY#A:MI8)X,YJe[U=MQ9_;8R8P911KF-+QaaJ))3Tcgcg
T9M;EdYO(T_?5,A>bH7]CNSMFQ)fJVRSY)J4T(O]4K8fZI#6Y8,BK-fJ0MC[3AMR
?.)ZH#a5b:GYgRIe1.]F:@#+>gS[=cQ@E&O1E8?C4HDPN#NT)#HX.g1TW^N/I4PB
8W3^5@>L7H,#]&^UR#H_:A@_/H&2Q(C7]-0_-+-\c)3[[:,M^K/X\:?E8#E4\\>#
JQG6Q)W)D#U4W(QPDY:BWXdV:YdS#;3/&L3&gW_(C8d-;=#LKH8>4O##Leg\:c#4
cd1R(77]YEb6CC&d_.(1RX5g_0JEePI<[7R^Gbe49ZdTY91&Y98JN1^<?Hd9eY\K
,<LFAY<#Z#cgP+9TeO^8O<[f,E]&LgB0NKR/P)QIfUg<QI>5&4IS\N/fAV_MTC<Z
bT]-[V&QP0a6M0]^?0GN[C_(?@FGWQSR@bVQ/GDI,<)K@#DSP=M:Oe,85>Dd4O]/
9?.(dZA./]&WX_EFT=9:\MI/MAA6dUD2&4<Q^ZDC:c=0@CC0+R75Q^RaU5E9R#[;
TQb22a7XDR<8G#>8d^aba=aM@U;&7.\#Q(([5>V.OEf=?@DBEP170R643A3E1<N>
O6)E(HG[d:WF3.BREHX[V&;;;;R]PdT^a]3fg&@JVTEA7B.KN_g0@WK/2#+,MbAL
gQM6)4bBfN-3[g@d;.@6O@e\ULC;98fN-ZeZRP2eT;5gIU33,^aEK6Y=-@eAIM+0
4Q[L(Zc;O1Yce(.B\4\X6A1eB/:2W(@&ZO3HGC/\+O<\T-E;HP/4>[W[1-f=@\@N
9#8bIM,c=bFB4daCEPIP,7B<H8Xb]+[[fg)RGK@cX?_AXM<HS4#8N.0P1W==VCT\
f^ea<aZ;M^b()@D4XZMM2[T#(;D@ADQ0RCHIS_POT6_1U>VU3EaAJ0DOf?McYE:>
:&[;VIFK>C7-2K^T]I8H;dF,PE#WaIN7[^gWNAUXZI23X+(D:&+d1J;-LI5>;^ZA
SWZPRVX0CNf7/(_Q8dSPg0U9<3YU9Z0>78E)F5aaC(@DdBDR&UZ59DN[_\NU)^>e
A7aU@Y=OCcZWUZ[f,<bdM#fAMKWWB_ECQ^927M5XWXaCQ=QD)ZN9F?gXNN=HHV^W
3E)GRS<41OW=Z2PfZBR1-^Cc&EDDKeN3S:aW3M,,L)CQ;D3d,,/1,>WYa;(a2K?<
]F6T5&E+W+/VKZ<FgEd[&&0Z]VPcMES.]4Q39#g,[>A4N(L)+>_5:eGPggBV^b;6
M;A+8\eEI2<(O&8d2Z?/IWZ\N=R.>NY+F/D@UTJgbRGPaTdJJ=G4[>c9W8X16M,(
&IG\L[C_OI-Y69<5Jd8<D0FF0M\cCQ@3A:daId6PC@=+SOgSPgX2I[If6L&eDMQE
EdWM(1+Yc?D02cLR4:WW(:W4@\QK+8P?UTa-&aEg1#]B;Tg:P_VKUE:;;LAXI#SC
/dSN3VL#[3#;.Y/?:_eL=9WZNN3=4D::ccAEPTcPN@?gP7\P@TQ8gEH#50YU=T1E
5PVSd0L,S^.AE+811FW,aUPUR9(0\:9CON[?&1YXVHP40MXd3>_GN&]d#dA/<^<+
1TX8.CdO_S0C:YdP\RW=/4.4;GDN6EId+1I<8KAaaFQER:K3&;6HTN#2d;PA7;aK
[]KDZHQ]OZDA]U2]fI[<C)&&1O-H;J>GA=@:cX>M6A9e:&7\3:;KXJJ5H<(@\QXg
;U-@-(c[HD)dT@VH/cG5-K^(#Z/V]W6#f&[SFO+GSF3YM##_8ZK&K=>7?13(Ne)6
_;a\3.=b0O@S/V;44.KZ#_9L7IE3A?]\D@4DR^a0(2KL&K;df5(-)E2QT1]^S/VO
_CFU<<1geOVa9BK2NUDR--DU\RHc(06O,BPV7,59g+,bX)L@,f@UY5EWY1,4BQG_
B))R;(^=,=\:]VX9P)=8ZAQVD_8d8V_\B).;>Rf@9[P#UR5E6:UEXW84Ua\S3C9A
H(3>>V72^bQ;bHPWd(S?]E7I2f:b9OA6SSMHKGJ/d#-eZ\O,A?RaGKN,>IV;INCc
dSZS@X4c[^NV86(SBZN@^ONOW_cY\-&KZ63G@/3SUacTYD@LJ)3TMYW[4b/#6;5C
YGVI;2XY)dacP,G7FPW4P5WMIWME\+e4_5MN0GJQ9NQRPECF1,D-9U&:G)&3S40&
&cVBS?W8,&HWG>#.);8P6g&20T6V.WQ)[8_.+UTVL=LOe?7DI<18BAc^5&\CT)P=
TRXdLE.gH^Q=/0-fQe?Kc;0H18KN0e,#J;Z]GHV;_MJTRS(]G<T?&9++:D?I>5:f
gKa+:?HeE20OXe,:<B8/=e?AO@/-IH.T)D785TKWXL_-+P/\T[cCGT;R5QdM4U+d
E?MXS;Ne0fL]]:+Ve/M,4&E\^-D3=7</^=;B(OI)FAF6BJ-Kf][)ecDXY1eJ55\9
g/FDO;E>[@FTBfE49eaB4@(cOe?[E[,>-K,T)MXIV7#2Qa/G_+@JP80DgMc-gS=M
=D/\-,M6[]B9/+[ZI(6#9ZJ,NTd2^X:6M-.L8&IUB3VA442+L5@_&X&a_52dgLEV
9K&I9?a?;(C8R.JQ6C,/RF>6.CHe\fI;_6UM[NYX6^\XWB(H[#)/7R/7G(#c@NWG
&ZGI^&ccG1Z6[Q(YPKaS.(bZG-.T>YIXd=PHVND-^;gFNV1:^IY-Ga&F@RXVW):/
b\KVRQOLO2BE\8bJTB;cW+dJd?B,_XMWQN8._&1S<\Qga9J29Y/G79CP#JSG,W3K
MDef<[,agJUG>3CeA^=_/eKONRf88=D;/TXMAgf13cBVJM+).3_9Y3XN]/c&M&+]
c,#+AYV=/-Xc<X5E#>e3+8DM=Z,?BBVWbBYYI9[<Z]X+G7-N1G];aaaMH(XK93Z2
G>e>XACS;.GeVOU9/#YEa<Wa&,4.2#>db1^>(=4V<CF(@1,^(c#GMY2S8)C44VY,
eACX2[YcAH_V6?fO]IS6CbKV:2>2I7Q)-A18P?790XaK>PSID?96?TbU,^[7BLGO
H#85beV>TNSecbc)PDf8>d3@@6>S;f+L9Fcfe7Q-<^-6\.,,=U<C>OLc-ZH)?UZY
(D63?L7[0_B,)\2;(0;dBV-:=HgS>D+\eLN^[d3RB[;_/+afAaUF28cT)DRS+9H#
.+D#<MTS=9g+/O>4<IH0:M<SN](IF]8,XI-4YPe6)0I@f+#Mg0g^I)3:^TQ.7Bg7
T/^adOFg+6H<=U(@c=[8\]\E.Y75)bAX;;gSQ3.0,VYc6[9d;3;EZZ[Ac4ENJG2Y
#XFCeT1+PYH4MJ&cA>gS[RIFU+:.dEO/;YTYC#ZU8BaKY2R#O8<1L;(QS9FUTJFY
T2@GD9bQP4M]C>2:Y^?@5Ocgf?Lc5:5bU(AM+]QN7XM0@XC;#S2dCdLKYPceP]7N
5AM],N028(MC3fgdXB7<3&8]T>8F[AXdP9QZ=ZP_^7Dg[dNHE/2B<f7O\>E\5:.:
868:LLK<UP\[@?8-d8KO..[6\QNb:UH<>F\4<6O4)3K+a#M_2BYKYLNC#+4E@\Gc
ARdSb74fg+QT\MLE3NDNcA2R,eRF>=J/BB_<NJ3+&4NCaOQF]-gS2X>(\FKU>;WN
BQT;f+4D.4:[Y8XC(.G6]#f67>Q?,GgVTbJ_^;RbIQG2R#3ZFU2,A@\JSI0[d=de
=JOff)C(QeKSMYb1#;1CWA)9@-@N\E(,M+?a[#2RSDT\G]GfKN-5gOD9f9Z/+6>W
OMVbEO>[\;(WPdRfUC_],QIIWc83D?[G>&:4&:A8<[fD8MU2\9/3A>\<)d-N,.eQ
<B)F8f)C6(N>NQ;6)B(-1A0\[1?V@A^L8K0We^#VO]=a6@4b)ZS@e/C1((9?)QNR
K4\+Wg1dS:DfG/e+D\Z;O8T\E3Dda(ON7P77(b.D3Kf/>O=dQJ-LNfIU;-=GRaPF
VEXN4]\>-[P/Ia[?HE^:D:9(@&BL.9^-H_G@I-=;)1#NN^L:2(#KdE]gdU33dFB)
[IIBNVT,7DY;3JO<+RH[FX^B.UN\TSON(U^egIaN:2FRG/-:Q6,?UK)B75MKT,KP
^&Ae(>^YfTZ#<9F8M.RWR,-1(QPg_&<Q_GK;dAH=&]TV@W+U#7.FR\CJ0=@]a=1:
0d:-_JNWV3..<M(-KNF@g8c)W_/M42_/\:74Veb&VT6&Rg#.:GbgU?CcG)LfaI]8
(3G[-6_GLT64;.BFSgLZ.\NNDgG=62DS+OMJF^4MOfWT#KcL)HNHIHg9S4L/BRZ_
N:@cD8(X27#fA]c9K)-<@,0_]2MA,^_X,1[Sg0c:A>_>^fgFA?YXQ]8JLd1_Z[YX
WfW9(&8IY9_,FZHJ69(cYN(d4?1Q6fa6HP&>04OLb(E.Z]RZ\68EaUR(f0^dQY@2
Z:g@6]SGEN)e:UAP?-;A@8@)_M5H#\,&6(]115SM^WfS;GH.cdfbFdTGA\&9:7UB
9IH<FG-#_fYYX=DF@d2?P5gA74F,LgF]L)1<;7((T5I&#Y)H3/d<Wf0XD+)9O5--
8>2+O]g-+Tfa<VCEOLA_=:D59L=ceSE(aVFV<?ZGg/5O/ec12@-C(NG1(Ic4G;:@
>Bf#.D6>K?09EFfQ&1ZT+RSfC)d;KJ+9T]_<.2f,A&2P(D;fAdX[[T@\&@O0#8O2
\)?V\DbGTQ_\.EL?7]J6#DT?4f?JQbbEH&PQ64fN<Z,#INV#4-<]/(KA#^AL-2BK
7?KJ9GD.aTURT+X^]#S7CA:9]4M_T@HZH_]ASM=2_[:.#BK]:;/\Z.=O6340(XM:
F6KVL8QYS3@N0_^;GX6)[B&bYINI=5B+_<MG93=URT,^J13Nb)9)AS3J]#;9f]eE
B=&[=GX3,H.Y=-PgX&PB0;;,P[-LMR>[=RQSVHJdeUQ/,<9OcW9d/9g5:90-QSf[
JI6B:O_)UHI1g(NL=U0:ZTWCLWQB:;/5gX+KZL7?CMfX\U]#2J;Z?9E<e,1<?cD6
@YgGA9KgT38N]M:R25CWA=#=IW[:g5UBYZ22&e6#LQ:A&YdeVOOR@E@[^9MV4aGE
C0[KdLWA)/=/M&_2eK58&DcFY8QI.MX711O]93/80,W/^W+gcIEde\[]1cG^+EEX
Mc>DLYL_,F_9FZT85cKbG94<<(/V4SL8fe]:.)eI,K,3gNQ4Eb(e?2&,S?IFdG/b
_2S7^,OFg\[;HO.=d=&I(F9G&-;V^bdKC;^_Pa(5U\F;41,T(@R+-_J]E/=&<(;C
IAB82H9W],bdc\ZY?Z4aX:O_R6E[(5XFOZNK_aS<+abMYVK(]H-1.P,dJb@H<R5A
(eX.[0^HG:O;SE>8?Nb#,bVAaCTUJY.Oc;e^5[QO+.V_R6MQQ>K#W[4R4WXgfVW5
0?JEd.9)1YE/I;2^.998Tfa+194&e0Z^3M#7Cb<DQJ5AG7C01WdD/c-@V[A=D_V#
[P55H@(<&&MQg0TM<AaA)1&YCATd-fS-9PP?<3d/<4#Pa)Y+X-b(J9REd&06cdRd
\E++S[fJLS8ES28)Ze85XU4RH-VV1+&3dIa24Bf(eAE19a]1_=T+M)ZAZN2>N;LX
-QYUJ8<5dT:6PE4I,W0cB<70GX@K3X1Q7#W+GIU#g1&WA4&DAXYIf6Hefb_\c->g
\<()(W;,LHJ1Q7.Q8T<SGba97Xc^4:(^cV-PK7,8gI0>^b>gVR(VXC,FBMZNS79M
U6Z?gZK3F<+Hbg(aB&:NI6[G.fVB3</>4afdFJQV>K)fRLO]HP\02=G7U/cV,VY_
1:bW/<)#Q^HXBVGT.E5DQDUSPH-ZN>GIONSgZZ@M>W>YJ.QZTb]OMf0#aR7aO];+
UO2Ic8Y7XQ<&FcV3=d\0+2OT-aa+&+Z#;P_^-<fKB83CaI]NS?J0C9\1T-E:Y_0O
HBOP/5]O8A;E4[T8UE1ba/(<.U/gfI]:3D[NA-<-M:70YF0>WE[E9QK,+ZN&gIN=
K_#[a+IDMJ#W60B<D8\4V>AMKK<J@_bN6;1]&^YUZ,#EdeQ;?bDZc8)2@\>f60YP
W36F1aD4)&EZVY,(AN+RLc]Vb-TRTcY]^EZ>:KTa#K#RH&+-eSRL<X7/Sd>]LCIG
a:T0TRKP93_XfG)JY<#a_X<2QNM/0]\_I0a(HQS)BZF6_IO[[b:Yd;DGcYZY>9,S
2-:Y>L3O2/;a@=&MfSFEA-2RTSg=@5A7_WECg7/J<Bg;JAI_AN]Zc5aYNaLFTgXd
]dO9[WU-M>Y_>]BHe+^/C65W_L&A;K,6.A>^-[Md;BfTEL.M1J6dSRW8If<H?1N@
:Ea=PC=5b5A4V7B4C>]=T)/d&3T6PK;NLV(c0+MZKZ^>(&1/6I5a-]4WC9Da6ZP#
Ia19c#;Q1SY.#@3IJ.d\.13b9K)fGP3GC^/U<D0H<#4M+I00WED7RgX>GYgSW^MK
F:2T+W8PECQ8cD[UbO-ARAOXYPP>gO-QP6=TeNNQX2,QE.^QF=)N2W2#5N@KVJAC
L#Ca-1;W2#Qb&9OOa,H(e^Kf#S5eL7XWbAEDMFZ_8D^V?0?)WPW)^cQeDS-K0ZS_
bG1&^_;PBa2-A03EdYM[(<6VRFKC8H9,FB-)>E[)OUNU+A(9a/]J/SSE>.7?8^TO
:R?-g&gI,1b&7G##S+S85,.Vg-:R/8Tff&K4P(0g\VUQ5A07BNb5_=9CU9(cQ.AA
Z.\7=HPTT1f6Q-./29_SV+b\)=)BQ0/aV3:I[,K76B<F/e>HQaX5Fb0_]U11U4a6
N.:[A8T_.@)Q/6(Fg3^beeD?-Q2QI(14[T_B-]:7e7Q;J>5Y,A3O0TV,<J(O-<:J
.PRK_G0D^>WEK(ZMd13e]4J.gS,]_@XI#AU+\H84>JL+,X9KCM@YKVF8cCHLH8F;
?f+Fg6G?ZG@5bX.EJEe:C/G@>QNEL[QZ,4\:UWO[7,D[#2CD))1&b9#UG+.H6eUF
O5PBBN4W9g90Md0Z+GQVP+G1SQ-P8eVJ7B_IT)LBaQg9LB-+7=0>J=dRbUCJ&0OZ
2T7W0J?(&JeC>=8+YdQfQ(4E?9934ZfP(SJ3&@PX]VFHZ;1Q&d6D.OL?H]G6TD1+
5E\R2EDRgC>V/>3&Y@N2=P=<A>:7G6&Ra<SMPE25WKLU,K;/7?+1HF>25XS39P^T
(WO1c&ES^fS^5G7g4IIS+dLOa5NS>N;d0JO-:)11T/fX.ee.987EKL,Y8K61334N
]_2-/QRfd1^ZaOG9XS4JEcV,Q8L?f:g>A)D1OW?b^RDgP-=Ng\>W2O.7G4,X:e4<
6NFJ2UV<Q>2<&BGS-2D&.7e.U.fVRf?-:,>711NL^W1R)?4XaG:WN5.GGO3X34P=
[WI+/.C+LNNa.L:H&)H((QF.b<\8H)/[PGR/P)],f:.e+4)DfJ/FU:,)DP@X4&H.
BB?HKYdJ.E/ICI-;XCcFQ=VZ.1>\G.\.+UcK^cU6.M@)MY(F8OfQ0HZ-6L&C3+O_
3@0aB<FgK<^@dJHFKcJ]@NWdDd&;.EeOD9YY[:T:Y<Q.?(.VD66(AM[BWSR#@&#_
[5QOR?c7)&8Y&,Q9^#PN1TP]_ScL?BKE(N2=J:PS3BVB/731+[F,=V=gD>8@)8OE
@Dg6Na0YC?^4Pfd\)9bTB(@3];c3>;R=fU5_KdMM+dKO<<8:.8#@K.(W?@/[d+Xd
.[][.5HL/QK+SSGCRg:K1U#QU[F@:5?/UHH7_\))));@01@1OHN>>T<5gD(SZR;N
H>_g->4.QGaFgY+ESCW3>I3EL@57EZY#0;OAF:_C@<HEB(7cT<&N)?G(,3dJYYYA
4]GgS)+>,=gIT(&C,aa_e13Ib[G++,\_+c(2QCDK)FB]X5WP?4^]UY\1MaN:^eCU
>53W8PHMUQ]#(Q9DCJ[^X?A0VUgFVgg9+J<eG3aWN;WfdN7@:Bb>LSa42#cLS1-Z
4(Ygg4>&,0)=a7dcUVWMeTF6;O]e[0?ND^QL;;TeFB?Sc4<LeAa@W=#8f8@?^GJG
d0P7ZCbV97-<[D0RD:GPf_8QQ&TZ;Fg9GXd&1<ARHX0LJEY?V.VZ?R:W?b<GGT^H
+XMc6LBC?XZY_U?=bIR4Z&(b5NeI&/\G22&Z9LV<gbDIS5Ea0:;,?/DA&LY,O5=>
L._E.:OQ=^baE-T(UWaHP]Xg0@PAXcTU:4G+e&)WZ2gBVfdDLMQR.^;&d1POOdZV
=Q-[_1=QPA]=U8?>BB2JF;NK_L3e:PZBF1]F^>)#/ZL5;OF1#RWX-;(cD2:,ND21
5GE-ZDE)B8KZaDXS3_]]H(/6FO]KZFLMb9Od5+@fDd?)Q1H](_9/B&^)Rd#H-f0<
T\)G2;UVLf-:OZd+C<1-+@.IG@E:FOIegD2\Me7AZT^,TFcI#K)3:I#RZ>)TTdE;
9ZgFKU/>BUZ7fB7Xg[Y&T_fH9<f3(\/69C_aYA,,55TU3<3FC3(ScY(eK[.g]DNK
?C90gd6J-[e8QV=\#ODa\5]Z+c@)7BB,#9NBAE:MXZ<\CaC&25S)6\]<YYg1T0=I
eR&ZO47C)K_G+W+43_B1P1INUEE6X+-7J;,EHS,W8\aY.H\+aGI>)ag-Z\?EW@HL
9.QSMQZf?(GaQON^Q[XT@a\_AYB^RLU:>B,^:9AB&=HREeJ>(g[KJ:&8A.>YQRe[
Y8FP6#X1MEG.TD?#+F3c):]I=#Ige\a/24W1#(EePES/APTWZ-g0@]:11;;Q0D1a
=Q[26;MJ[/<==Y?I]\,H^201(S,-b(WNTZ\V7g,CTP=XfaU-HY>D_;cG<cK6Q@ZE
Y88J90]d]V:\IZ^3=4_MeK@O;#)S]9:Q^A)/?.gZ<)_8d3WKPER@B\L53])5Q2ML
IQ^&U/=OAM;#VH08<^5U5N@IC-C.+W<Pa1D7M;BI+N=AcKEMNZbKZ_>_PB)0d>>\
(Xb5C9).R.:g:N]D+8e>M)TYdHD8.FAE22HVO;fZ-6Lg9<-BLU,CIa,9ebZ2KG#5
#YQga/E]X?@P)U\=)+PdGBO=NSC2OH,F^1?Mbe^B@HC\NTJD;Dg/^\?LL9/&Ef_U
+gFB7#CX(TG3VK8?ACe]-2-;5;AZY;I;Wf8WB2@TP88G)gH=B;7THZaG<Na.f3dI
HRcDD0[@aaJQ:C9,?X3J6H4H&E;LV/)U3a5ZSa20DI7Z_&@GU(_dNSAKE[Nc5F6U
D\X(TggBagcX)811\(Z]>058GCCGC?46AVMJ?e>\aJJ@,&RFX9a4@GTWAI6GL[Lg
=2(3+5&L4C+?b;<F/[5eLC5I?Q#L,G#)]U#VF0J.>][6LSUGE=M3@E75U?V]<8[:
g(dQg7P;d.1]Ld:?Q5bdCIQ[.G0<AD=;X]8P,;?90bSGd-[^3Y#B0VM_>0He<.?b
KNO/ce_<NE-d[54LC&DLcAC)97-eZ7VE/EZMU^YB,B,/c?VFK<2:6_[cP(X\]MZ0
V#E,5&V]>WZBS4H^9g6f4Zb1[Pe=&7)f52:\[>e#XG_gd<T=DRJ?]\4Sf-=>A&GT
&O4K+].(M>^#M/]=.GM?V;/Z-@K(_d.U_->1SQfAg,.T7/5(dZ/8Y?-SYR)RO0A@
/>H_#AO7)6=D[g+B,.ggS09CD8[b00e<P+>eCM/5(2:C2T6YSPEM\F0@E\_3Re=E
6GUCed7&_<W&K=;gXZBfeQBa+8d9R71;GQe@?1J^>F-0]&=eH4-EecY,=YM.XKD[
:#5<R2+bQWIcE?-bcWR=-g_:<WB[Mc][Q)ZGF;Wa[^A:Q<YLO4;W(a8fe^0@f3K3
V85ZFXB8:73F7H^^0ACWM85#-1cLT6X-2Q9&?U@/GI2)#E]#)R4bfTCX;1DF?d/4
^UaOPI7L\Z,EI82#ZS2cg\12Q?ED/I=[NO;TP[2&?7aVd&McQP/CKeC\gE:GBIWH
5DK:((;C)_1R)_#K=Se,6SS2>XdU6cU\OEV=#LP.,e;8fdBH@6S686+MT156&O^Z
ac]GV=2d8/WSW>C&aNAV2@6RR7/-2YX=[B;fS2WdM+:/8X8LS-U)@ABBBT&e76bc
g.(,3C-I[2g^X;)]Z1D:I=2ZB5TIT\/#+8ZS;#4Z0a3[8\\Z8#&0#R.d[^#c=ObH
JWXb>8NVU-a27I3O\Ge2fQgD(SDa/RTC14+L&/[eg:RS5.J#:FUICGa&J=CX6eB1
>IN)NZ^BB37KGUCe&O5LLE.(#&VeeeXT@1=CW\4dfDVVVIRd97ScKNT@d\?K1SC<
7GXDX6F-c:I[M:Q-KZE<;Ze0ZYWZN,B?R]2c<L^N,:4<eRN3+-30GDLC?MZeQ5bM
cCVSgG2SRgD\Wa/L2O:?a6bU+;_C#JL25:?CCA);;YOFCV4C<dW<^,eN1@+2WQb:
(9KbeG74=>Ng</0g&N7MU>\/?@S8B/](#JU;P5-^4K[=+Kc?Xcc=ZBgMSFQR:123
/b?f^8:L.I(8;LEMJ6\-DeE^VUOga[\S.0@cLd5U31dI,8D]bd^:#--C+U<^U/+/
7Pb3bMODgWOP2S#f<8)/S^JJTZL=EB.X2@PdWXf/N_T-F52^0&^=6).\ZJ;Z2Z8_
A<POX2#,,[eC@)IW_W(JR/H:F+7(Ace6Z&=BA6ARF+EMXMZLG55[NDUH#ZZ>V3#0
c&R^ZV(P?4.QG?I:_[=OVNU8@0=#<W)b>gI:>-@bGZ5?--L2GYAPTB:8Y,5D2aI>
60810-3>P30G3VYPLL]R<ZRcX:MWKSS4.7BMN9E35O4A>6=,[>#</@&I#W+/?VB#
]4aeJMV9R(QYBdK.>BF3?HB,,U)6CXZQGb;dJ#[dV\BI;^B=>)+e)PST/;?eSJP4
@f@(T<P1IJf^KN=C/XQ@H4I=#4DO9^/Ze7B6=?M89+S3+F]MSX+.[)\VYBY^6fI5
W&@bWY@Fg0&\R+)79+G]P93c9/S3L:fZ>5aZO?agdRZ@aBdXTgI79@;Q?:@@1H<-
UB7LLc\K^bV1\F22JZVT>Mbc+:<\TggP@K)RGI7E\e@WX;PN\J^,c@H4BfKG#::C
(Kf,I^4PUgSTc17FRSAOU<7V;CP1F?E;L:g4Ld_cG.fgR.f2AV:=egT:5Q1[-5:R
C77((be:T0KXF>+&>bc/,:=6\YSK4>QUBHBfC>;-^7<MBZ7:<Sd:/Y\_9bSfd&8&
cX2N3-K5>)@aL-RSIa)T?PX,+:]D6U])C.G^Nd<SH8BWN19X)8-EY(>&6Y/E/2^_
?<6T@J5XGTDQ93SK218E4SA12==>DT@BQ+K/CfH,6X<DFXb;+1O(QUSZ.3-c9>FL
a@BE0NF-eVfR:8WPe;:FSd0YB<NV)<+Q>\8/-e5J#0GDQN3_:UIc#dX4G#R&.K+b
>Y4LfXQ,Ee[ZCCY>\9<:(EHN]LR<B6A72)c4W>N-4/6PCWD?I>.)gFAZ)EM4U\U:
,SVDSgF7JMa#G-;^.4eKb9bPCI^+UN2R6M;MU_b,6[_+JZJYgT>NF(+9<f6T)Q?.
VP0M/E/G15X>7REf+c][XYZ=2T#.FeT5:KWF8f.a_N0H8S5&08_?cFaVK0K/I>Me
8\a=ece3@\PN5/NIS+(Jf>6J#HgcVT&PIBI<a3+GP[&H&aC&^Z^(13SYC+E&:-d[
/9<]/8SR@1TVEXS0P8PdMb^10XAPI2b3U=aE2]SGc[+1?86KJTbC3OQYPLK826eV
?A,TZ?@^=X^HM:QdF4U/Xb#(P^<[;J5UH/R5/N(@E:6XYZa(9WL?f:3+5[Ig2<A<
AAb;<VRG2b(0CF##F(Fb8ff[M-GaX@G:1N\BHVDNC/DT,f#]X[f\9g23B&[+e?.<
dLaY0?QeA0MV92AK.Q<@ETK[\LISOf,L,?XB[OPbg,?JIOXR=14V^B/=gC,QWGf[
+I#8HL:/.;ZO^TS[8eI313U;39B?#\>?TAAK-O@PCC7NS11JfH0^JY9K(#@=;C#c
1MX9DRJb[<FG=R3],c(AdY/CDc;6c.Z>PJ^#1])eL86.@/S.U)063&7OUVa[I/e^
&C\_GC([O[E3XBbG957-)OKd>96IX\MOM9J6:S3J/];b(3VEQCVF3<Z69F#BP7TA
8d#6bDE(0X]2@]?,Nc=/c;/U;^HJQaO&\?34/D0\<]:9]GT1O&PT-a#)L1HE:B)U
/>23I5;BBH0Yc,F/N94LdT)c)XD(E6ICPCS_?CZ6H.^)WcIYA(0Z&d[J.=;;7a4a
;VG1+F&E[69f-GJ(RNQdYfH[9G2@\1)D\Q5g;)ARBS2?&](=A6L<1\I;^[B,8X#e
Oc4IEaeR5A?FY1:94,PPB^?9NZCWd2AQ[::24G[SEPgWcFDYO\aJ(L\4EbLWU=UR
2@2GM_1+,GHD_UMe01K0^DTQ93\HF=-RZ-8.(K0:cVd2XQ1)C,8Re)D;5=O0B4BZ
FR(5T<9Y_>ZCQQR5RJUTL#&J0R^[.;G<##.OMNTGQ]d7eOC<_?>J7>M,&T)NaT6Z
2<McQG.4ab>LU6Ubc;+.&0EBM#J?F20=<C@(ZU/<1RU2Y.@f,95S_KD&ABT1EgC)
c(]A/OCgBHDCO&AKU#)<(5LU[1QWe7,NHAL2Ya;Ld88UO0P<5_cV1GXMVDC\DK@e
U+1O::32UAaC9>SQ4,#e,fMS008+VcW1V6]4HYQSW/a;Y/;BTS6,HOc>X8J_@6Y<
S=..P/db<+1UJ\[@<)P/R5\3JfFHQ7UG]BKGZMg9<+a=>,9cLUd2gId&A:BJfg<3
Ad;JRDCGWPVb3IMC2.^K6O?[N^gVU(fW&C?C2bNX_PBF5)=3LGC&UX2619MS2YUa
S:?=<#H+Y.dE,\\09>376G/;W2c7>>E^f(3W?g7f&/@+S3.TI^/PEb[ULJV3ECAf
W/0aGc]JbeQIHX)A#819J-NZWABbNdIc;7E3;HQ@dXWLW26O[[,A2?MF;;&P[IY9
B8H[W)XF.6A?+d#9YD5/U[@c+/Df&,91V(XJcc,_U>,)>?X#J&.He:&C^6I7>d]L
@JF9WY<GgKH2LbV<4^3ZD?RW[,b,d3UHQ8,CR_G&U:D)_@(b:eG)J1ceKZ\O_e3V
RSSA:JOcW_]X+7/U81(L?]eb]:KXQBWQX[d@SGE<G:?L^Kb#+R2>a&bC<1:=5W#,
TU&.fLS?<QBVJ0/M8+eK<F@(H>XV)b3_7AD9beWDC(cW1=Cg<0SdCB0CIR?cKSeg
?:#HO15cQS=,_M]EH,Pc7a<H&2C4,O=9J?PX1cSRRfL/AfcTaaH,3,MBa__R9Q]d
[/T_R,+.GYJ=1RQ2J6WZ.5X7EL]C#-HIaH@#M&W;8?EQ1QHGAT+W0CC+244&1DN,
/R&PERYESVJ(Y7T>Y8#6UDfX>T=GbB421OK_@AQM(]ZO2QI41TU^MWX9g5/>1/>P
CKV(.+0Z-#OK[2\2=#f<1V,,/]IP5Q5YO[SWWE5MZ8]H0YP46gT:OT;&]LfTMd6O
aeFM?B5E=G=O6@N+,_B9KHQ2C0PcI:R74&Tb\)^C@9[e6L3#eOWX__XGE_Z.d5+K
K?[PaLGNJ6e8V-&_;:Y]@2E.KS(-?,CW:#9=P4T>G5@M]34=eWH.Bc?E^0NJWE/]
6Z=89dCXGVUAE0VJA?Y6&JE(EB2ZP)f-+G,3O6-(EIJQ,R9W(_F]]fXRO0G+&(,;
+-,F(7AD==MIgZ=:-HZf8>;=ECQgR5>4g,UK^Scf00WfZ<4L,+UIFdGO&M[@IAbU
474?@[T6F3)P81E2^(7MDP9]Q,V@1e?G_.Q3=]9ff\M[cf1Wa46405Ecac-3X,bM
KA&:gMA:UIEUS5P?S=T0DWU?EY@&6RC6\#Z^H>#3TXcG+2.(RI=FdW1?\-&XX2bb
FKMPKE0J9E^<E\EIM@I30g83SfLPdU,dW4PGI2?=U9,cV+FGc&K9.0;-ND\0FQ/A
ZNZ5_I7-N#=[(,4[-2MfHI;].ZM=DHVS]b?e3^WRJ:dZe6PTO>/9fRZI2,,4]fWW
V.\V(ffR8U0Sb;(7W/dHbIJLN;HF(D,LCN57O;-9f\/:L+ZK,TM0AOEWa#G)#+(d
3fg[F(;a?=)Y3RVfHWP_TP=\D:D18,6OC1YYVM-^+>Mf9L?dM8eE=>b_BTQ/f:,^
<::J[&,A/@FX<?X(g6+3[1Za]E2Pd._S^_P(DWLHRY1I]fPLU-VcaYXHN<#@S1GG
c65PdVa@R\K_a01WAS6B57>F5)=^7aVH\.#c]55_0+-BA_3_3,7NJE8&/ML^b^I3
G<cZKb8X3ZZ?aF_VNO57J@f=4)c2LbN#-TTK\4)W;W(:7=#Y&[4JOR<E6aS&,F@b
7@C<-9,>&^fTU0H(Y>&TGcP2gM\6.]42=C.BW#B1Z\EaR8BL-Z[TSI0:].F(/IUc
YfR,PT7S4ce=,F-?[bV9X4Ke)2E43)4J(b2O;;)+eIG?e<.NKF_S\86QM(YK61V.
2FgDO,YP5N3VKCW]\f1Y;Y@R<]M1[]+.B&SRM?)=3;-I4KWYVR8QZWS3,:9R>X?I
-H\6TL1JI,Y[UX:)4Sg(g3S4R@R5<E7D_TQJL8D3+b(g?DC-I0FcM6Y0Lg./:6X:
?>>6F03:1)UP>6=<O8G?4HfGA=X#;@4MNTPCP&81G&6\ebd.c=[Td[CQ/U,^Lb?7
2B(<K(5;_H,2[1EK[W<;9?6E]+0JK8[>^LIP(X(FM.eP=@8,:JVD_dO)O>SS\CK+
,3^=QJ]8E8UPS3JA99W6+gd15#eMWABWRU:HHVc?@#WQBJJRZca#eFHL_670\/_?
,+<R[A8H?XM1A?4(][WK)7I<>f#[P]4.c4HPNg7e;YLIKRgMbXUN4aS=/.J:.C@A
Y=gE@(6aPSK6cQGagMC9&F#P:a4b5bBgYUSaN@Kbd:N;B<,Fd[9]Ng-DBF]O-H)W
.4K(8ZA42BYUP24E9;)G9b<V#SHgHX4T@9bHYCVZMZ;I>[0NK2_\]\bG4_OEQFP6
Y@LBXOc<&X\c?D--M;7O(X]Tb_1Xe#38.&KggIL:LZZ#XHVP]XQCaNf>QB,=Z<0M
V2Qa\WBVZEATEQ+TF?>G]K&@B4d][c0,C37KVaXHZ05W3dW#DbRaWP0TB4^>2@(\
N-8_^bGf:]RCZCW4T,T5Uc_LcY&N7SBcM7)5TAf)NS(5G1^J4KRQ@9_V\1HWZ8SP
\3E8;gGe\THU)JcJK?d<LTS0^^gARFd[dD,#4=WG0GNQ+U+@PM&WK.T,)E?R+GN:
HA?QP.3(9@dQ-0:IRES8Db6NLI/AV?D.&);2KA6SWJ?\/J.,OK9UX=4R8R_GS9#a
L(ge8^KA,Vde0B?dAaZW&[PS?^fPO_bU-McG1C:&B&b^J>IO_<dKI=5TVQ0RZ/)L
H7D^]ZgdA(X(2>#W/_T\ZD[)E5DXMX>_2R=]U^OA\ad:NFe#8cCZ,,P[e#>d+[?S
a9RET0S/&J0G:Ic72gRb]HePc[:e)fWM\]0PKEJA._a0Q,bJ.6>WRb);U<Afe)G;
e0[ggK^+A>22XMKFWd?VO]EC[)T^ZcL-E^I:GUH1O:F?[IOKZ,,VG_f=>5_gD^H+
eWfVc(B(=],=OJK#+4_MUEZ#0R2_JE^VI#@2>>:QLHHdd:<DPb(K;N-I2eLDF,Q.
]6B87fVMMZcQA2e0M^F24K&GQM1-]RMU5W35(6CN,8:Q0Pb#(RgRX-_Z4]?GGM,^
6WXRDe/>81<>GND]0UERL,WY@61DPD9D1=K4<S&G\aM,&-SaP42LMb@Q-be@.,RB
3[3UMT.>T4SfY?Z2FL/?-M/AB\a=dX_)Oaa(K.)4G-0\WMWW<Ke-d8T\CV9]AJde
&VOT+b7:fZNW7XaJ284&2->]^@ScfF212SK.322FP/;eCJV/f6NQ\HVV7_cf6&BY
O-9c6,)+E1]I\>.EC1DT9fg[b.;]d90.8IB9/&Ye==0;=]1+/0cCbU\fJK^4+L4N
beZbca_#\E0D/N4g-RBe0EGT;N\:\)=Q6VR@Ug0&S#KbQLd\4F7I^(Z4H:#I/A7:
0MLYBMWg5c[&:eF;,7gCfO,=TbA^WBXBQ?+K8H_VRE0g3;MJW<ba(bVH8+QdZ:#U
JJHa0B8[bM,Jg(B,a#\AWA;d]7,A=D3>/,[MPT/f@U_:Y5SL7UcXN7Tf3]+PROMK
N=&Na_K[_?3d.R-60IZP+F3YObYYLOMf\X>[7P>Pg\C;bDG<+<Y_7BGX,VC_I+-1
MDS@.(J=EI]Y?RVZ8+Zf4MadNY,?,,)bd8FM/O69\PLT@&YWDZP?>5K/M605;HD0
^LVK20&CQWg6,>ARHZ73:AC?^M>=T1,KX+<5;MJL1O69b](9H\LBdOeRG&S=Xg>G
5@:8TcNNDCb];abZ.\K=A=_9@=1#Dg)I[@5WA_T(8SCRE8D&<0NgH(CT]#A?gBB=
7#VG&>(N2R;6OD1aBJ/(R^6N#Q+E1c#TZ:TH:[cXa3Z1A6XV;J>2]GTL1IA-)-gM
X[0+9JXOOd&5(OfV^@,bB+H-)K0P[&AX51(@<Vgd//@I2A_I3,#)a1>Z)(@/I\/d
PRVH/+B0fSH,]<T#UQRc:TG=11^Mg/0F^AUH6Mfa#=W[Q6+\Ve+c\.EJdP5G<b?8
E.SX;K1PES_.-^>;b:(XL+FHR15-^;-0MQ_@I)009g,NS#[A##G(H3S=NK)\TMC.
^D,8JU(/Ff3ND/>^M03.5#&c6e]eVH;1?;I8RBP6GAPJT4AWKd(^,=_8;IW4f,/9
?&g6/eb;A2,Z)M0JZGe\44bXI5M\(_d,PLaN((<MDCc;CTB?FAc.C;Z>)N05G^X4
&>1;=I?eH>ALL_;8??cQd4G9aIJKZA-)0EIUIe//O;W\<;<?1\F5.DBUJ>d6@&HG
&fOfD-=Le];7>eQ_-C9)(ZG5G_Z)ZW39LRJN6YA(FP4K0#X9H_,.Z<7SIH4UKT5>
C0).#>YOW=UXeJNbXDLc3]3&34QSTdES,GR]N<OGadJ[-_9D8Z]22R#:.Q(3S;Q^
(f\QMW&)8=?QG,T_<J7cfL4KaBgSMP632IFK<3L5E<+,2JSTK.F[^4L5-C^>QdW2
.=3R?O>8^N0,3Tg#S>^LPWENFc1fR]KCd_IIf:8S8_F/@@#\\S?348ON<N+BAMfa
TXM+XbgaN_C@e]GW94YL3,P(R_XdCPEYN<)XgRfNMP<VI\M=)SeG#(M)A(_]Y<[.
e3H>[/b\T8-24;AO?;_-BGbW,6O>0@&Y+eN/XCb]9HP-QO?cE7+SLOI9ZZ,ZM,+E
BWS8GPOG7#+&f>@9=V-A<U-SSDHK2&dXSJ6OgNV:.La&=#+;_K<Q[^-]N/eTAR&9
<K+7OV\(<;O;#E[MB,_T8=bSP[Y^V^0M84/P@Y#AVX^XK6[AQ;KdZaWD9FDA?.P6
7>37R\g9T4>FAGbgaL_a/4UFPc+8RQ]cH:6QV2],Q,SYB]:S8=X^e)dLBg6fGQ6c
-274aEdR.N;5(_b(,;:S(FCWWb<;6DfI=9D?0Y1:QRFgU2Yb^K=JKCQ,R@]-O/I1
/Pef=.3NTc8f4PEeE5>,?\,=SGP<Z^>ZGHQB]XEc/#af7Ua&E4aBT,W)-fH1#ML;
7]b9A#DHLTE0\EGMN2E8B48CM(./c0eGL[+7b5<\#5+L#9KbARK3KAX1TT-NF^QX
EDCH@W+<e5<#[48?&+M6fCDa218:gcA+R/?0:_GdgTUR4Pe=A9>W2O>(gR-:(Mf@
[b7#PXDR7AeDJCa7:C)b^cA/S0e-I47SbW8?5,#)#_TC@KF>CO4OHQ9F<Ce1F=3d
U_.N4>U1A8\,Hg>+3#^3]@[3+GbEJ6[g/cO_O(0=L_6>S1BWK2f6GW4c7-PG<G@K
cV;;6CNc-)8Qd?UE/e9S5<6Rc::=WGOd;.B6A01)E2^dGPZaW/CCE,Cf-]GHFbK0
K[#eY>]OQ?\JdB2:OO>04(,2UO6W8=FGCMXA=]BbGJ:H(,-7a:a+>,_/#H^(fQ0_
B6JA1=7(#-USYEWeTS,M^W+S-6L6=LH_XI,P/8P:A\E1a/J;[cH_afXOYR/4.=]0
/=4]M/BHJM6AK<@_.<R-]Jg8Nc^T]].@aVU6W=)O3aKC0.9,R6:1AcQ-,8gI@=W1
EVS<[)gXO_#g62g2\981L]?E2cM]f(K4O[=5\g,U:C4bcRQFW5Ld0C-UK9./Oc?1
5W6U<[;.dTFLfOeN,BT0(6+/&EeU]L-;gP67/3&SK8Xd90.&cZZg[9BbPT#]RdW+
O#D-aJGVWKW4O7[TAE\b9HG]==g6NC2^CCb;Y;/&8+I)G>[>e8H;&gW8T_#;c;+b
SC:a?KEa,PGS,c=dd>+J>1X4gT1_gVSE[MYD(RHO74D2g@H>G=a&6bW[[c_(20Z>
Q;O)YReTORPX@L&/N]DGPe._HRK(b-[K>R4Y=.O-VM3d<>WEcVD<NRQM?XO=&LD]
3TR2-NA:(+?K.cSfCN@a5.+(X9ROB_ZdE1EbLa-N2EN>Y:Y-LPgI]JUQP+W1/MWY
b\KXW7XI2gF>IOeY1XORN]c5J91\?6\d5\N_e_ac8>24F;,UU[?9EY]&\GH5Bd+Z
S4>D9-b)#B-S:=5_(4FQ3]H6>99.K8^?g8LZb.48,<:-J5@5be?AE[J#/UOe49e/
52HN]bHO@.e:e.X[VQd+:E91N\:7\>X3L3B2/:.[L^IK^Tc+,SFF29^>GW<=YWPQ
d7C&=NUYb+LUTZA<RXgQ(+ff0S.(/7BAG0aSgZCdYV@E((P9U^N>ebA=PNFX6)6_
WH-@2V\3aAdd+UI5<J)Ob>&BH=gBMW@Vc-P38MU_S9fO>+?@<(8Hfe8:2J5QU31e
[4W2)6>?VE1,:^@UaK1\(_Sd_<8K-H2K[/#X:5Xg/Ac(@TUgb(W-^&5-dJ\[#XX)
7eJEcN@C[]f0[9gd83;F#6@M#Qg4W8ZQI1<YSHHDNE8>@?f&[.G,b_^RMEbNK-J(
UD-@1)13\S4@L-L.?<@).QCHLV-EQfc-]>CV46f,&PL:VD]KZa@+WPdXFQ_(][E@
#3#3RQ&JZUO7gVUWBb0..IO1H^Og3_WL[RQ]>GAOT4#-.7JXbG85@T18^#BL_&\+
RZMSc?<3WAf)=4U/H1;M>Y9B78Wg&dJ6V0@8HB[G&2?9+O_A--A5RR>g0413KT4G
67d3<XW>AE)(C];JeLSX\gSOY^BH4T9>DbZ;R<MO/V1953IUKc_RY=&[/XERU?,Q
:bK&+][6gM=[ZEEC?c-f1A,:F71(P<\aNUAF534Hb&::CKC2DAK73==c/9R=[MB=
X8IF<Of(N-1AP:ZM,5M?&,37c6PSI7VE[0ccPG2_1<_2S^EFcEF<Q+A6VA[d?Q<T
B03I/=&QRWP_Oe&?BD#(V^:X?8d7HRN5?N0P<gVE;UHX@DX/XG7S&&2B411D&)F;
?Lgg/cQZ:cWd@2NR9[.0C71?]cC8P0-cGX.GE#T)EQb,2b?2EO&F:;\MKEOO6Ia]
>f;aI.fHG4_f3(_KL)c<LOP100DX)O+>Tf)8?dK9SU?/0#R1JbKKe?Uf;Ab<bJZ;
bEa4+]:O+8N\:[[#5SXXB^e<daR5[TT<=M=P.O/6g4:XTCKL,3]:Wb[NTe+/LLc2
596HDa\XeCggB_X<2?]KH5J>VGE7/f0<B\?H,.2C\NM>;5-J+P,<VYPAaY#7<gTB
2-XI0dYafK-3RXNX&EM3R#I?7b?P#:JU313YCBa+/PU,5E>D8=2?4A__VNHc:Oc>
#=EY3MEV0+2&PGTf[gTN^#DXIVL0XC8VB(Z?cK297e+b34DE?F>W)/b[;:33bFMO
TD:/Zbg(@;FDU?UYD&@1W5^(83[;#JR,]g\4HfO7CZfFZIGRZ#G8e_LRU::7cWgW
B\4M7Z_->GFX5GHbG#7;2J389^L@-Nf::E.2,85^7=GX<(gIKT0eRV,D.M&E/FT-
IFUBA#V];PV]5C60B?PGA-.2gNF(bL1ZLU;&BR&[SQ\MJU9Z_V(^Z+[Se:5@K:(3
aC/86_>7N)Be)3ZL\27Z/8FP4?[+(NY9/_M3Sf(R;_IEc0,.&.)GISGaZ(0_QZ29
-AfB6YEG=QSMTC.G-3XTbdHW>e.E.bc?]2[>0BMSU/#CL5[g#,<1BP8XZ=^YXBLE
^>QTO49ce0WG?;9db-S@YaXX]08JCD0D@SQe3LQ6W?9&WK2XQPQ8E2LeVJYIN-/F
M;4LX0[;5c#3H:Mb\f48-:O0CDX1^=7aUJ+fQ.D6@.-^LFeX@KMVe@<[G_9NUDIQ
(Z1<:ac^S4Jee?36N,MNU^#Ne_>]D#7S/<bD19;M&58HBN:JZC(>fP7FfDD3XegA
DW-7?bVEZ3c3KN7I/.ORa/2<XR8c.PdUcTd_<g,QCY,A#+7@YSM11cb2#A_2c&b1
H.eQ(b@[(dUKfN>8>):<&#VWMEB:/#cI5J^BB?H7]7)7?a\8WU@beQ\H4[.cPIFd
1AKaZ3C@\d/dG0QEHc#dOBL/C>;+@\@IA(0),Q:.FT[CT?a(M#,GNDYU_W-1#S9L
EQg#&G>5WT]ZY-f[?DLc>-L7[5P_XGe=CdQ5TXbI1Q[@1g#3(&CcGNRC?1eE=V0R
46>c58X?W_2K3?M9K9VA(AY<X<BY(O;e:X&4&Ic/OLFBKXNf.5^?N8(F2;\F+0L-
?3SMHIaf5_]@C3\c8_gg@QHbb@<Y\?:QDEU#&<4WK\V:-ec[KX/?8Q,A/O;8\89?
Z564eLP1SBBeP_[OP;+][-J=??HWTbY7\26<MG:g<3ST_S4,Zc/f5ORd\7X^F.=?
-@RH=A15/6QeG00A9C3;-7\4ZQD4UH7(R36SU(;[e]=_#+5S,b.J47@,T1L5GF.,
X/SB^QU6Qb4d^B]H[2S;?#R1/RcWSW?6gRbZ:gD7cD;L14@C8^P#QTg0QA2NQ\IA
JF<;<fIVC1gU_([Yg.-/F&T-):9eAT&-W#e/aR6_J2#N#9(JFWNY.KY)59C/DWQ0
eg\^A><1+.2dRDAN,8^T[D/I\3,[7C4,g:V,fWQ1Pf8U[c#cB6GSg2?dP/Q.HA=Q
f?E48XN4H;A/K-R4;^N=DS?.=)(PReb0/CZ+Fd;)09aGJ-H=c,;A:b<Z+FLcR08V
:>AL:Zdc#VD4Y=]gMNddIF&70561H]6TW/dUR\]<IcR5ZOd?_K)/26N3<G=F-L_a
MfW<R.H#7?N_[cHJBV,UW73#EQGc/1L18+Sfb1+:B9&@\SdSM(Ya(1?/UA)OF+D]
/ESW,^F>ad200C9D#8V_POf-F.gJXe1QZT,#8R.PbGUJ4T.22Za/)=5Z\KAeK4AM
/P=a8)BSIIfB^170cCTS8cZLGeOUB3+^9+3/H6IR0LaIM/YcBG5E<NQaV388BH.\
D(W#AbaUD=3+cLM>FBgF<f,3;Q)=Xg&e>:ND7P7aVcE(9aAA\?ZO9;Q.R7F.5O41
@g5Gc6+RXcUc.6Ve5MVWB_2&8VEaRGc2FE+5f?^.:C)-VWFB:fIE7I25,O+:UNPQ
HOcP;f8YQ_#b=A0B>1V@?&4C0LL;YcME+SV6WAOVfHF#,^U)PGI0]?W3Bf+>TO[U
gTD^[+@S66C8@-(@Ne<OSCF+UA3,Ld-_VM.0&d9@S@Gf@UZdYE5c+c@&<gR-8(LT
9;aF++g?AIKB;FI@>([Ce>)RgPC2_N)eFM7J1M>cTgOEZGI?&\V#JcNbU/C+\2RW
:d]=WbNW];)LR]&/2d9FE4>NXUT2E1&:^A20X<MF63F#C2+]+e,?28a8>TX2..JR
b,,=F7C^M?aDZ/1&BGHB7D.VFY8,S5USf+b@4cc1Le/;d/Q_/BE^AW__-/MSgQAB
KTZ4g<UE@_O?N<=>B5]L9EQH;IC+aB##AgE75;I#0fW[?)Z\Y<Eff=ZL,ZA.+gab
5[Z-D_I5]Y8:@LD9ZB&VT3Y+2F_c16gE11LGD0XJ)Rg5.Z5TX83R@DbV\,?TT/=G
<GDO=0eef#V5Q&Ob1/5+[gH119Qd,]e=Q.Y=22JS,,.0;\U@.BeR8HGD1EIgd:W9
O(JW>\=_UcM0a\Rcc\f3F:<J6WWc09.MWUOeP3XcPV3=@;+Qd1?Fe<:c-8NW=/68
0[]^YZ3BO\::[I5748Q_dD,F^K=V_/K_NRVgM.F2Dg)M]af_QS>g@9^8V-=f(_Q5
AMI-@KafKU&<dB(TCdEC^8]DV2d&b/aSF19.F,=Z^<Ye=EHY-b;aO1]^=X/:IG3a
Ff\TFWa0J2NC4=GSRKQ?eN<4-=\#+K+T-J6V@cPcQJDD-K/.SN_.D&ZS7FA&8>)9
_OMQ21XZR\0WgV_89Ic(Ja:MPO()LNJ#@Z,5>U9bSb+QdV;2X0663,[XTb=29JDW
M;a1>U9gB4T]V4]GaA\&TH^[gRF]UP+Qg8TNf>]&fI<=5KKIN0M3M.6R+8+bT&fP
D@64,9V^[O++UBL0W,6>JFbE0@-1YTMb2KJd7+1-3Od1VY?:B.N+S_afS_;7_)6b
>6+-(c))/OHT@J5R1<;^P0bRF_H#ed43(E8;F&TOWFLFfc)IaC[/,_5S\d4f1&dY
aMB@US5aIQ1ZS5(gI+eab#=L0d8W#S/#7\Ze2GfKXWM.[Dg:RZ?,O.8Ig3<M)F8)
C)1ZZ#bSZ8R+cT5+a@,HGLLOGYdOD=RNc45RX66V<>2DF>_4]QXQV4Y03;VfC]-f
G/e4WMM.9>FcW;]g<Z6U@8]+CG,H1C@gaIUO7Ac>S^Q:V1#<G<+#KAN_XC3C2N</
@;]bbW3cQQ_H:,Ca9PMQU,=bG&?^X<S?PIS2(08L<Ng4@M#5O+ddP#6.6\fbaO=<
0cg,[5KKCBg)dY((>50V3(-9)b1eQ>C=XS_/P,D.P5/GDAP+MJ)a9?[NU7(d5Yg\
cXS.E/#MaSc4S(0NB30&I]WH(Cce[cI26,M7Sg.4RI3,S<d3?K(UJ?0]+I+_DFTc
AdB7ZeK&5>A5D.P_SU+.dbQ8(QM9<ZN122&Y^SK1+#c0c2W9DV4TH7NXQFDOFZZ)
gQU3TF/34KNQ5O/KJ;FTO4-@69B<?022;RA0a(1BcH66/Qd(<[G^<_SaTF[<>TYM
XXK[H9gRQA=#.):B/Q5J@eCL2P7D\8-[;YG(TC)I@P3]<NT:b<[^a93^^a12#;_@
Q4Q2L?^80bX,g@+,fX.]>R/PK^Vg0R9YCVUgE2KCYV1R(:S8O9P1/^4O_.a91AL8
;d)+4<X1TC#^).EQN0\.I)2P6eP/JK]L#ZAN0fDE/;@(RH9..NXJQQ#2&(L,IXgU
:&YAa5?^0Z=5_RcDe+LeESC,:>@9W5LDWIJ3c5=KcYQG4c#H,_SX^3>1?fKd(?^(
gQ7Y<b\.NH,7g&gaXGTS8GSB)Zc^b&C^CH5-&X4VNPJ_eMU^)S^N_=64A,FDgMT9
28#0f/X7>6=3<:=W&WdT98F@HRT46L[f=D5gN7RDPBg,O6;>f9Cd1H+5.Mg_VO1+
&DcOX@d8CUY??HHOYG<XX3UR-5,[Rg3[5H^Ee8[ccc3T/_,g?P,#R]7C(U#^(aW2
0V+ed=1X3FJ5]<@A#=^?cLD?:QRW=c#WFQb)d^^>6CK@CHAZBU;?2g]=A2CF;^]8
S#[K@KH.:.DZ5aPFDKK@5)Tc]cS8&7UUDBB0#N@cgY@)V:+?Y3C/Z.U4/S2#(?HO
8G4)0:Jd<2Sc;Y3RIM6bGI0V>^/g-eg:#@NQNC-L:5fe4QNJ@449=PUe(<1<VDWZ
(2KUVeNASNCT55d:_F^CT6XRN9B+E<H<F465NK\SZ=X#:/@F>(::D(NO_:0/V49@
03V55>SZ)\9,YYA&7bW0L#-SNK/FV#A9Ed#aQ_P5E(3-5J?TdVgfcZ33g#<d#C/N
46\F@cK+5?f/QUQA/g04(ASF\Z:XKQaHICS9#:FN-+DIYa0[C^cUV[QRA\O=Ob@L
#[:[;;8M^P;=_cKV&e.g7;f:gI]Xb(,F<7&Y=(bC]=]EVM;FGI:66.BNXOYe,WTJ
/+J[S62Se?CS3197M];SW#?,Z9DQ\-67W@:\8../+Cd\^@@UZ678G-+X<>KBP:a?
cE#J4M0P6\P?=GL?RQ(.;6bB;(Ic_=c\X?,T6bLg9;KfFJSB_.R]L\e\MK4P3F:-
BH@0\Y/E((V=\SdNA?=XC)FReP\L@^d:UZJeV;4CDg;dA/,,)TBI-5(ff@GAfISE
+Y4WEJeb3LTYa]6W6IYK0,HPa7=X)7_K,K1B]f0Ga[2)b(]Ia?;F3_ee\J1c?B:f
;Kfb3aQEM8?:-44E\4XAbO7Qba&BN[CU@M_b_H=[0a_P=2#3^S@NRLL.FgT)YE;K
HdgWfRU[A_]39GVe:Y7JK8.:e;L_a,L9N2K2[eQX.TIe:M#/=R5Z9?NLb)7UacA5
U)1)(aeQ\O6UH1OBXg4a<51L4J#eO7DC#O(eZUI-T>KN;&c)B1eAYcSYe@(#M[>A
EGTYR((U&HTXW-[.]YEdROMAGYa4b56[:<T:4)bCF]Z=NQ1g8cM>0_Ufe4E2O-0:
>Y@3?QEaUfLCf>J\ZPWW[/3#@,PMR=@,[TZQH77D+R<F_;V[3@(4(bWHS[#DBT/N
\&c;SC7,\([L5EV15N^H<2N(Mc<W>eK)Z6QK1BXJeVKTY+-TUf?_/>KI_AA#cEcC
&7:/^3<-e7L7G,-&T-R2N:21g6YULB4O,PK&AV#43K;gdGKZVDOTLQBRQ3+0R&XB
OFQ^]@K8/I(5(>1dRe=JH2\FBYgI]gMYIZDRP(2LTH3&/[:GF/f\fg1<3P)_:a=L
>AS()T-N/,1XZ)UI1aG;34H46I)RgN]X&KY#8U70OG55:H6ggX;bD8_Wa(GScE0H
eOW+Q9-&]S\/J@96R?=I(GM@,?A_:>]QeLeOI2MUGY[,JYRWS)W^]+)MKZ2aDH[9
->fGDV+A7D@c+[3B<8.3Z3PZR85P1.X6b\gDERaL?695#@^MbP9b&Be/N=MY&&_c
SM&e=0>3M[L_B@,Q[,O^2Qb&H7]Y:efa06EQBYAZ_L8.CB\N]5)ZP<O<;cN=1Q)Z
],,c[JTOP^#(NMNX4D3ePK\a<7.PJZ9+<YJ?XHUSSY9b>#[:34)S,4OeF.R8K.<7
8[&aTI>+DHe_.RF]CL+M:=&8KI<\V1Xg/_DVL-:A=^[dNAY;ZE3/6._NQKE(&CUT
\=I@<6FVV9W[SB2&(bMV/PbA[KGWU^P;K,?[DK?]FXeBEdCbO_fY##b<T/ZH1d;[
c?.I_KDg607T&T,WK4Fbe22?3>Xa)<>BRS08M8,6X3C2?_(7KdGc&X9K9C1KaE-&
1?OH&^CNKY[Lc+3TOS\KDDCXW7KU[e3W)?>95/#aD\IgK<@ZP/TH1XBY0?0<&IB1
F(ZA>^4[AJV0CK7A_g31#Z=R5=&XcbEd4P9K;_VLR/E:g</F([KZZ4M#cKG<fDD7
HU0L+e8c@9aRVWJ@bSN#IEJg;]6]+B8aL[\:1,D79_PN27MVSS8M84L>P2SKX=H>
[^OA?Nb)P]TG.-HZEbVS+.L2-J[GEEb_K_0AL@3@gc6\3@4L-3<#ZU,:Q3J;0I(/
_8eJJ:<TMge:K47OI;JE)U>Z6dRI)O:ad66D[VST<eGaJ(55GG@-?VWbbN#,0)M3
.e&BM?Jf[#6LC^/b?>f@CM7/MVT3P:[:E5VFE4UF^R:YR+KF@)NCGTOcb3eabcW.
C9CM(YfdR9F)R1[a:Z9cg<b&_Ga5aUFY=^U45(Z5KTW]-fI4O+5egd7P]bO[CeO?
4_<ILDX//EK\>^ebJaCN&@3^dUdQL7/PYS8PaD-dF#&\@B&^S5?RgB,#[/cXGZ]:
Ba7bD2eZKAEIbM]7A/e_7df&12KM1gO\(//V<c(5\2(&0S:8MO_\,[D\bMO9,bJ:
?V)><RZ<cZ(AR-,Y0/^SLTd^JcP_#:EQ0>f[5H6f3aMAaD4)-\?:9P+\0FD8_aeT
:F#9MBO7>::2_XJ0AI)8OEJE4_0>3PFd9-)6,<8fa00;/G</e)3[8IW(/L1\JNVU
Sd)]DT3dVNF4c><FWUg+(P:,gH,GOIZfEYf_554MGf^]fD&@^HZS>-I9614:9S..
:dPKWEaB;8W[.H(.b#U(7^FgLBaYY0c/>GXWc&d)dBX:e>.#(=fcfIBX^L\?g8a=
);6&DC)[CL0a6/_@7#^9JO5KT)0)0-eHU3,[Td9aUI&5O<.-08K5XFLa,cBJ5?._
.GFE-P>17XX;DM7d8dS-^Q6d#/I@Ef=3bLKfZdYO#&5LJQS38I4PH1^Q\WM]X8;_
gKM#IPD>@PFF1fDT.+g9I[+?.S8>49F2F=F:;VSGZ5&bdY++Ua=<aQ/9fG,RI+,D
N&TbGK]_&L3aGB/B++E1Ie^)[MM#8Z#7#^g_>27g#^9b/<N_)0:a?:KOWU0\5S2K
2cJfa#LK.@,E2<8g3R?BNaH??+5^B@/Z8H5A5QXdJMFfG58S+08.OK5gON&Q9U8E
8dU&HgW,0A.N,9X0F8MNe15Y-T7^Rgef^YUMC=7R7ZD3GT_RD1O\<C[Jac(4HQFY
>[XJb:9GHQ.#?HUa97L<Z^O&HN@_a6>[M^gF8D8-fL+YI<V@/8;aH8-AWS2<1:a8
L&;3)V4IG&WZIWNT;d07M1[IZ#UI&fP)#6FWGB>LJM\F3UKC=a)E2cZ:E^A8G>/+
&\3:.]:JE5=:=MK+SYd.,Zd@HR-/S^C#-9F:9V[^&&Pb9f1Q+(a9KI@IE<9L-ZER
7PU_SQUS)Jg<a#;PHMYW.\=5##F8=WVL?(CCcDfF6&f,UQSf6#U_0D0/@CP<4HfW
26V#-B.bN,XZbR7ALd2<:BK:RY1d88gM1_7-&C_L:L+NHYR(J,FPQg+X[;=E<-87
YQZ4M>&EF:eX469XcR:(SN.I+_#DUDP\c(O:.DY5a5HHO=[8-b(5^SL?I9RJ8#GC
]=QY7(UIRBK\G8)G@d3)O?]\\:43Z_fE1I#<E6^-\EEadR.2X^CBfP==8[dQF@5Z
:G[eHA3)gfFaL1=L=8.Ug.X-J_#DHG15Og(:S^-=9g=]L@eBWg70Wbe<UXAB1N2V
fNN#gQPg)V4.Y83):2.BcM7>0g(VF6EGX&P\<gNN;WaP,DO<8W57)I0;G1.WLI_3
.4_E)ZMc_cXP/&51a#Vc+@FFgZK5UM]]B\8:1OQF,T7(^(KM5]=fEf8GNb/A/BGd
eOA\8BF534X^YLDMB,1N,]SAG5S42:E-8C]AC,V[KRU#\MG1GD5H\,TbD8[K2VRb
/VR8DJIGAgAc4X:d5<<Z0E01IO7PA+I:PFYLZ(de<;8=d:&)^<U6V0=I[0^:,Kb?
4Kaf01aLEG[f7EMA^DH<1A>RZ\4=9S0&9CN=&SCBE\GHT;fK3]2(19^V\A;)EEdG
+<<J//ZZ9EMH7[9O1CU9@IZ/L9J,b2f5a6S,Be>P));3[TF^TI\2+Q\];VcT.1c?
,EL+>]/^#04P5D5BH9LQIbL[6GcY812@MOPSCScPddcQ#V=BEYK\[Vc1cEM(0_-X
EdI9B#3KUfCBK_B@Qe>)V)M9-SD9=f8.[R<CDgD[HY9@KRHUFWfTfaa^:M+\N;Fg
Q7+WZK>HJ(Be<-P,N7)M1^]?b]P\&Q2KEU9Ve6&P[57cIDLeRX0AB:]f\?McK@DC
Fc,>=VSSGOZ;#a-GK2+9VC^H/Z]d-]b&T_/AXeLGT9U+R9KMPOVg9(LJTQ7-(A(R
NMNEgTN&1]I-5;0Oa?A::6gdW:Wc@.:&I/CPI/L))(@K8A-G,M-2V5]05Z=?ZV:I
VI3Y-BSB0[>9Z/0XUZ6L^DSF26B_cZD&<GBMV/Ag7NT?4c2/\ae?R3@dCVG>,0N>
V1V4:e3T#N./I.2JH\[=KQSOR@8fGY59AH]eS1;6&J)<M_O58.QHA<:)#1EQ9-K9
16.5](3f6CLYg=:RQ^-HPM^E3I_/UI^_E:#T,56O6OE3I=SDM8:J#._CYP&47[4X
-g2/g(,XNZaQLP+,PeL@U4g,-<S3\UbCe<@)>>fN-0,2\de)fd8I4gc/a8;a@>ST
[8L1@1PH3(<ZK>(1aPcNQA7=CcV8UEV-Q1;OagK7VHTS.=f:3V>HYTPW)+7N60+7
3e[JaK8Q^-I)V1<J[83bfZHWQce7.H@cc:GG](Z>&.Q8ECV?-748b)A+<=:5VHf&
7D\P1(98e;d&ALZE,(;F7=KXBXX1>b[DI8#T)M,dV94eUAV]X/Vfg3R=N2:4_L#P
Y(7:OZ<^bO@F6Jg2C[g.G@Q-5IO@[Q:ZL6J^61c;Q?ScUD#N,b+NC5HAM6\S:_A]
\L=XKXTcIM?7@JU5,F?LJ\2@Q7#8b1IgC^VG7--L0L1^bKO7g,/C(6)ccZD/JN>(
,(Nf7I?WB0DX3:^QSTLI6K;UVEc<\\c=7X?VX2J]e.4B.,:1fP>4YF]H^0RIT\)Q
.H<((E3Z2f<E,(fS)-EX8eDNUB6],Q\8dRAb:@)O9EN+F_C,VF+FZ-f+dF2Z9,6U
<]E_282?1&7SM)A\KJ01&d(Q)27G.?f4UdN4Q-5NS59<aPM^SN3S0SL4+=>T>RM/
.4+cb3Wc_4VYd/6H^9WG-[5cb;ES88<1SK[N-R8O9YKRM6/Aa?N@.&L5I20&=4B;
)J\K/;#:IY0<Hg4aNeI.V=+=B;U&5G)[>^cfD)[S:1bB3:0>O9LXD^<Uf2<PP6DX
a=#c=@?7M8>J<^6fTeeeB(gK+2(;T^?/e.^]@f=g4P.b.;6S3&CXJ.<8W/NUHd;3
Z8:DZ93V:B&Q=,&V9H@?)EAT(;YRD]PVNCF-@_@D,EO#HXc7AY\/MWg_.,Z^AUV]
PX]-,#N8PaF[L1A8Oe:fCB7F11Z4YQK]VH8ggYD\V>NWX/0??<1ObJ2cX./9BB-J
WR4YJZ=[QN0cKMLQ/B40QEB?2]EL=49BGTI.7d>30f)P;2+9TaJfQgL&NJ84Y-C/
3DeYP[WTHV1@b_CQH),;YS-B0I9K80@Dgf1@#<:)VXN]GIdPffdb.dC=JKf5[G;f
=SGT+bd])=8=c1&&-/c_a-2&)dF^]:[)BT#2IK)g<gNcE5#SS-U0:KUTY;YFDK-B
@4N-E<QUKFg;&eYQFQ6#g91N^ITFI#T9[X=dfD8>dG:_&X8(HF^aO5#DdAUV,]:J
\-Q?OZT&>>+#cG)6D#+DCK,,]1S<8.[L.-6?>1#gK7JF#J2Y33Z/J6_SOUb/9.HV
(UGJR(<\I96^08R6RR1;T>;eHB8J^+=:^ZN<_e1#4a/aJE\^^E[PZRWeDTdO34KP
?3Ge<,;)6H&WLWe:,-K8BU@1.dNM6A-aR1X/=@,VL=d>A@:J]Sg5LRGPKXE0A^F6
^HX+T&PIQ.7G?b+<dC-KQTS#e]HS1M;3=aXM9/3gXH[O0R;c,O3:28bN@WX[A2f-
9f#6;gZAODO6JW]<<(N7#1HHZ2^W.3EL)cf8:b^S?=Y]VK<_eOC@WX6g^X4OH(TW
c\<JP:M_#]ca@U.VZ[;?5F0aQZPW2Ga>cZ_C^9PEI.134#L;9O1L4PAYBN5Ld3J/
ddPJ]T?E?<L#T<IMBW#d=6S,)0a7b_YWgH9EMT&MAOPSVUKU6F(#?6cJRe.5?O#^
FTZG)H1@d&9VOcZf,:ga2LA7(^GG0STeO:=G(4=]N_GD;Q)Cc9?(T>L<eb2>CDEC
1E\,<E[MQ5/G6gWR;dEb.>0/SEF.(^Y^R5H;LA&]6S-]c-G8DC;9W^JQZ4]ES-G2
E6>GbIgVNa+QDN_O)9<QNb+6LBL8G]1]JJg3B=beH\eeZWW]&C#YO,NFAcX3.f65
(,fCZ6Q^+LZM:3P]:/J>N1-^7W5Pee:I;]B@MCWgcNF-MDFUK?V]KPBaS<fCKY@.
=>BJ@bQ3R^(GE-6>d)ZIBA[;@&fQ\WMM)T;MQ^0,SP89C6ZE+(d[WZM)XKg]@e7b
9_T,3#?O@AX=(Rf0(YQdf=,LM^2GeAF[<c8UGGK/P-GH8EESfVF76-J:&Yd^eNW0
/N2=@96Ea<ZC-Td(JHX1]/VeVC;EeU12^e&<eDI4TgXCWc<NZ&FIbG4XV4K<CTOg
fGgBD(X4<[<g.=B6?GA6[B?3Qf/29]#_<-NMN)8RF>gHN_\<5&\F#E,H7(TY^#=:
#>;@N,)=Mfe--QVM2E/W_@1NbG;;_If_<FHSPS,>?fC4^[J2R\:F);+8[-D>W,<D
f_S#H2D]T_S,cHbMSDE4A?;CII3JH7Qf5X:ffY2B,]a^d<)-P;:2IeG.9;-=P^Oe
E[e>N-838KZbD@LN;<]cf^IAMAfKAZV.5,ZeAe:d1PI/.LZ1:^WbPa.N?U3G4@fW
cW@Qd8O_J=Dc/4cC0eGFZgB;BJ:#/AG3Z2_CBB5dBHW&[_474/d:dAJ5UT9@_IV=
P_ZU5We.J4K?M@gE:LRMN+[g@6f6^4RYT;CMTKa<X2OaEg]0M3#BAIIO@RP,.8)c
fIT(WLZ5I1GUDbL^;AN8CPXPU9<[MQ\T;.1F7W3LZ<006O@M6@.593aEe3DFQE&=
+WT0BbVc9f_;N70(32/V@?.,WCT:cA2]P,5Y@J4UaE?g8X)c9.F0USWdbbY_N9OZ
YbP&9O/<53ZeY4_+L+f2g1T4ANTDT3dFA4(UHGR./:UYU^R0)C0M:;e(a7V:-XWe
X_1(=(4&=P\fV-\-YR?6/CML;0deE<g2f2SR[c,^Sd#[c:_-:SUJEA-[YT4^D(R^
Cb\K_^e[@fY^_O-Tb_&.529]R9BEN=M1/H)#0.X5Wc@DR4)OBQbCK8:532>aTZ.D
:c]GHd]I<IPeEB>df+RJb->;UOEaVD2a<3)[SJCd^,4d:&d#;7.P\@7>_cE-7O>R
@P4cDB;VW)HGTP,/,1<X/f-];CYc)a]EgW;,J3<^5HDO?d#05aa]bRDX-)8._-9F
RC;Xc?58a>E@38Q75^Eb@>Q,B6QJWL)(-_LN7QSV?W)KNO&g[3+RfbDP)<K:1E>H
+?BeTZ2-@)[+CUJDZC\<P,8QB05Fd^+\L2?M<@6\S=P?bL?bMc[\&\[f-OafQaIS
JO.bK2dR0_=:();4)XSQ)2(,7>X-WVGa).ZB(F#+cM8<)aA>A),:JNH\VUgI_4R]
HE1X4YN>=H0LLOcY/A[J#=?b>JP=8\B]A\V8.?H@8gIC(@e@KXaaI8P,N])ZR?2>
Ja4&6QN/ZLf>d(b#._ZB7PPCE7TD,<,4FL_&YF][\VTdVCdA35Lff^^@dUD3=\5>
2NGGdc_\=)1TL39=S\Hdg6,UPaBG8(I#6/@FO.F02Bd7V=(f==C8)][7<3K^JR;c
1O)WE+ZZ[+B6;LDEB88aL5f,ZTNL&S#F8\?Z.7;(K3Zc)8QYd:^196-N1,ef^QAJ
c9Y=^bbGa5I&2FBPK?+5FFBY^J9b@.f[eSSaXTDacR)1J,?gSeJQ<A:a_;1Q,5aQ
KDUS8R3Dc.BZ(.6\T2#Z_\CdJeTeccF_/VeG1V?HL11Z,f7ID\F28-]aL/a7eKXL
;+YdgLOfM0;23Of6W#);eVSLBUHVI4YSE;O0;@^E6Kc(4M:)Rd2#B?[NAI<8Tba3
TGc/0a7g([].(#?G1.JZE3HGJ@1\51Q(#L\BB9Y[<Y]N>eJ4bVWP_2K9FGH]&,#-
72)gX1a6WcC5KK3?f=IbTH8^),5H;@Sf;,;(&?QB9AK@+7;U_RBTB_c-)8JYWR1^
),A<FJ,^[]V5Sa_EAM59^Ub>GfLF\A[XKcX;a:0G<N.W9\BBF1YB(b-=<58#2K)1
3^Y6,U:5Q1PT>J8KA-;^]_FL-RXfOLF<]JA0:>RVHIACS52<F5.MFbU)FHbP/=#J
]FO>X)<9LDK/]X?f-+Y1E7TD\7^H/8aJMM/W&TG)U(7_Pbe/;CR^?#a0P-9/3@XU
JB1e(2O<gL\gVgQSAF52T6>(8AF3V#[dQ]M8V#aOJD=+#&,_4+ZUS6fgF^Q-:X@+
[MAHSCbYd,Q:fb.U89A>:T-KWf&Z.XT.BGCb6Xe&TCOa&D&R>B)@<[#5IR>LH##g
L6E:EdUc1be[ZJ<U>3.E?N@-149b45I=-T.8[_0E7aE?)T:_GB4Xb31S1:UK=?-&
SFQ7VBW_.,]Ga?A24NNe(QLYc07,4@2TLa?5:-7ScI&;31U[U?@L#C:7(#M:<c(Q
<V1gXbP):d(F[+FefTbC<;+R2#ZUA:H4RHd^gAf=61B2K:2/dWC>C2C\?MVO>9.:
=F_NZfVeUUCc2#e.,4;?UT+?8K#25T.KY60g6W7[f7<4fUN:P?DdRN^:&WF=D)@W
D1Wg.7^:G\P./JD5S#&4<093)[34GeJY#7)@[WY/N=(UY.L[:=L/.dKf)FUBI.9<
\:J4Zb_L</UR(4U58XP?cNdLJ;2J)/g/E5D4V(<@&,2S#cEL_9OfU(d2IaJ<UGQ]
YcFUdSR.915A^MbDWZDSeI<GdaRYDP]V,>UJX8SX1XRI(\HT2d4&O#TJ(/)X1;C4
/)3]T#;BWfI@:Z:FDEf3(K;4f:^@N(TI@&Pf8KZQ59L<V:P5QZAU[[(BD+OB;Be]
RI7]SNLA>-:S,_NX7dH4488&+T/fPgcHcX]L0@gU3gFHEI<E\;>,^KL<NNF(ZB3C
RNZNS?g-Bc+\V^b];__M8EWeZfMO8cE&/d-\RUde<;MTIOXCX95VGE+S+gQ&(B6a
MJ2+T<8<gDK;/aT@(PfWK1H0J?V,EV;+LUg3SUEJ//8>M?(V-,d4fS(]O]6+Xa=X
d;WU=GQdX@&2-#&TF7)@/a_+T3b8fFUXc/X[Ia.75K8<2ObBde+&Y;R.3g_GB;H2
(9aVO178b];@1ISR\&PWO&eF6EOXCNc8aBBQLZ>;JMX;1JI<]FR7eZ3XAN2?#1J6
D\fcJ2Zd@d1+]RIC9[9S&@fPK[&RDJ3K0CK>Rf2Q0K6O7F[#FW??099I8/a/YL-7
S)d0P:P/5J[fJ8I)&Z,JU@,US>[MXeV6VUW7C\\3a-0a+bJ0C\-B@MIZ;]ZOO--S
2:>G4F<H#5WK,9g2+dGfd[6X1ZY?6U/::I,0[XA=2U/\B<E:5CAI5-0>aY:f4D,Q
\c0CD[WJ+\aK96=^OdYS2@Wc4^1b/C(;;2;e-C5bESYK(>aJ134Q=+7SD32BT8F,
VZ5E9/9NS@33@2-a+4L>_=I=UQ9E=4^:A#KXF^fIaAaHD5(B^+90]30LFDL5ZR?@
=E\K.Vg:CY^Z]6cJ.Se+,b[@Z&?,\f//]V1TaYaK9U+]8C7ANNM9Q6BZ97WLS/Ac
O.\fbOP400=cE^bCFV/(/(#)CfZHg#?QPQG\O6/W1CMV3C\_A5KL4&]9&IV>O0Fd
<75?9,9dK_dg;NR7GTSP;P\FZVJZC=?e,U4Z,1+[B&2]D>LGFM79?=CWO[D;(2,H
PV[,E0Jb+?:(c-#D6))@_-HRD)bYO8J72SV&&0=F/Q4V-VU&E)6SVIS8-?_WDEe]
FcW]A=aJI67?)MMXBF[VRXP;D4PeP[J;e@<B_7KU>_MI8I?GRdH7SG;:HLSC:Kb5
376b^DAC6,6Db^4]=g)(#^:Q.I:ISBP0K1UG]ER=_(8@bReV^08YK&bce@G,P)gN
\P23EQO[0+&_&fLV1LY8:8?M_G6#d7@c]O3UdXMW\b_V61-;_+3^J.G8PH(eG/1J
DUMXI(BWQcd2d0_D;;T3+[=E#?aP_]JV6&94d;SOH\X[#Q<IbEdS/K6GHd/&->,d
bJFT&1TJ#3)^0/GXc3TgSc>]TJAURd=XcGN975U&GMKBd<;_-Pde7:RgR2I)4a<[
P^MEC>..-Q9Fa?O-[LJg3[:5>KS>-9Z:cCZDSJ^U^-DX#6,_G6TH)1(bTW)WH2L2
HM_E)5(F;U(_;1Oc08#ZK5O>;#^>c.VE9FFG8S[A=2\:dO)5.Nb9G;>\JFEESgW-
<I^/4G4V2&T)=TKQ0];QH6KW[G/^.VO9H^5YbR@J(C2@YJA.(EbYLH-.0f;I(a3.
W+I/Hb(G9L+6dP=5H@4I66ZeaG(3D16W#0&Y/63d#133@[0@V#[,32=BLaeAEGL/
S8f(&@O,UJ>U]3P+T\S>(1E-@X.4?+Xd()?6E8ZTQ.I(e1e(f^ANc]<^LaZXX/]5
#Wfb;bQ[NE)-ge&R,@=5G[ET7P4.,aT#Z+9L6,#+cDJE)K_:Va]9ZB4Q:?,&#R67
LY406-)N<\H_B35X[.CGNQO[0=:AVA-N-.FRH(<aX]@A7/=eI/^MOHgL+4<K6gPH
G<_8,B65G8&PYJbce2FSe2<>8K?7Ub7?Z9MW.d[R:cCaT.Y=++0:Z)_@aCdSeKNd
OJ+PMd]^GH:XY;8N]^FDY0#;SeL?.=(RcP78MV2LO.\KaRAQ&_fEBX[,d_.CW4c3
?:3Y9PCY:Q@0BWd-;cD@_9.(^=2T#^/MaY(?IX:],gEJ>8YcE8-g;TL0A=CQb\N#
_5Qb=DaHZ9I\V-&A-2LaEaSf#FH7eZFRLgZcOQ\]A@\Z5;].B:PbAE[7;YNG.VS<
LBP+Ha_0[UNKU&?5Hge]JR1Ga@6?gRJRK2#:E==c(B2aYQb:+ba=P80(,-V.X_YK
aS,OP\A-&Hf.7I:9eX]T>\T:fP<CR_=8[T:XN4+XUAGfD:De,\LGbX2NM\L:,>F7
P0HeO/-.UaEAaU)S,a>)(ZZHb.77b@J^#MKJ&9M<G[N12L^ReD;PAae&?D>D,4fb
d/HBJIRH]:&\>>RfJH<^RR/-JF9dJ[#;(2TH]6fgcL8fdG0Wg]R?<(F9HHJG#.NB
,J@,gUY2^\@J17=^I27FNa5O=^;,M(ea:I<NI_0,FM,CaUeNM1[bV<+/(W?(5Y4L
7L/0P4A2Y,/BH+b]CA:9(B1/.XXLfcZb+J:OM-7^5U>N()#UC5FP<ZgNSNV13I8F
/,0#24.A?A?<NeLS\f?cU,=2JWZ/f>9&]TaP@+bgIN0R[,/]bAcP@Q:2PEU#,[K^
D,;X&+dT0,dN_H\P;/\=#HP.R@.O+;<a:0#Wcb)IAe&^@8_^G:DCYSDe<GZ6P1(P
EaA4W@QDJW)9PfM^0W@)Z)O>>1b,S#IGT?,dc)OL]&G^5MTdVTSaY9FG.=7O.A?^
TEeHH0)(g]LeD3.M8]a@1@TKcWCM>H&?M1UC4F.9Xe^/^KC:R69@WQ;E@44Dbe;E
fdWAOa99T^DA,>0_#Z3^R#6-R>c0=5MAXX[c7W;N_+\_?U2H)&;9eCFA3-d80;RY
;dO^&L6LF.O[aSK,TZ45G@>&N\)-dS085f;Q>b>E:D=8I#&?&/<4g0<^6<?Aa=PJ
O@f(0Tb30Zdg]NW4QAU(Aa>bH^=SXfPI[c09I\F6fBMUHE(:3fLS^f#@R=Ra8=^@
CfccMN8Q5A<:(9/_?2E]d@0G]X7XK5b4?;83K63S6FDA[?&<UAZ-F.S5Ga\]4\7J
3,_TG=:Ub=8J>;.@<O:g:W)0aDDB8(CG+GF>bLK:V751G6KOSCFN0]<Db9;\fH\X
2/FQD3ASW?e?K/VUF@e:0]IEZLG@&8N)\U5eXQdJ;Bc?3Q1cK02XWYUN5Yc3&GX7
SFI^NIMVU@:>X9SD>OMY=3GW&#8FSM#Z8,e.LGY)Q?ea+Z<#[X1G(BR])DZaYSd+
11b#=#\fcA>Z1<J6g\9ET.0aPb7^1UNS+ORU-,@-PdJ5\V2DdDT>..+CQ3(/Q?A\
L5Gg(9b(.5\<\.?B8IOAZ<2)O^-.g@J0NePVAgZ.PCgT1=@2+BM4P]1E2<S>QaQJ
D8O?_=g)E-U5JZb8@SdS.K:O3?@&g69FXDF[J+d),1c3D87<C/WLQ.9/,d(g=P4e
UNdPC+B/N)eSgDHfC:=M\gZ0aU2@g]/M8a^OPOZ_/,S93bIOW6[=bJ6d,4cgOZ3[
>8GFg@ZF8QQS\5&GZ?,]0X[OF0O;J0?CS9_SZLUg@FI2b7&_Q7BY#JZ,Z.H8+U78
JKZJ73A8TOK)=6#63S4]H2aEUH^FLEg0:8(81]B7(Q?G39D,0gAbMa>IU[=SB8CM
BPf_+>N;)KO6O_P?,.H(B,eeGc+JJaACL<)T0eIeE9R>(FB3a-X_0FTCcdWb0Z@(
VQ1:5+A@4A(eZVbS7<C[?-eDOP,#b].SKUdCC+U.-GF_+B,:[+J7dU(F<Z\VeSGe
S3-(f?W^Z^N;f<=:_U1VeBP3ZIeU_2^@[U2,+E0)d-d,9B>(<K.-.(eHZ9LTFHSJ
+eZ^Ag_Z(?Y.PXCLSKdPNgXM9dWd0@^+2>@8YD6#?MEGd-E.a>F-W/+AD\C;cJ//
Z#(VWK]DZ_3B6;eN)-):QdEC6JWQ?5_734I2:4U.QK4?D5#A[K)Z#aP3g2:9ETX0
A3LK&,g=-\F\>EV^,Z1/SVBW=?+GX&K3Z<.[R:P=2]H_-fBVdDb8,5e?9gVY6E@d
DO;)\_<.bX[<.R&g-EVcKbNGQ?E\=K+f9M,E]+?<_&Y+(/7<e-?73BJKQ0U;+@OC
PRT><L^MXB,)OKce[3.83M\>IBQA)J2-TfM=PY==[/FAQL[.W(&K@5gKY(6U^E&8
LYOd:^/TLE1L2B/^RYHUKfPAZDK:Qd=e,U.+&C#1ON)?)&,ME^RP^P9AXNdMVM&8
O=^GR@LaRDa?_)c@Y1D>M\V,egG/FSR&O6UGGK1/,]R8a+fQZ1bRWXZ10\-6Q?W_
@42;3=DQTJG/[DGN;9YP&PRLGQ/+I?&9XC[bK6deM8FQUFXPaFVRZO].I+6(<5UQ
)7a=O\+de<OPZ13@Ob9O&SYP[L0.OaS2de3(@=c>FCC[JFY)T/4>Q.7aVW-8]>>.
/44XAYOJBff:0]e:;&[WM\<T+E,&6f7PB7IS[MYX6SP,e6IK/R=HfF3+EE-L65Tg
(?GA(f(:U+O5XT#Q;CYS@XZ90]72I-V+dVg_KL:M=1;:7IdET4P7_H3eB.bH5_Mb
<-5;5d/3H5?55#CD>Y3bSEe1gZdWXg#NO1=a-D[g0>dX5:G<H,0YJc1)G./D[Hc+
6.R9^Gde\[D.NZ(BJ(/cfN6]TbUD-1L<I6W#U^E]^NC&DI0JJ<bKRVP,,#2P?;1;
JB0QJY-LT))TE4IXc##VB<ZN\LOKA0N/)c[,Y)4bPJ24cc023YRPVQ,E8FFA\E1H
:L_P9GZ7VUAUef23P]d.RY\57PVNIb.J6LcEaacKg.[=QTKO7gWf56gR/N66<J#D
b9L7>0=N]XSMN7S+9[2)QYF:8N@APY&W+-8D<NX.?0H3?W>OBC3V9VH9U/(;.=_J
G[R732HIZ[:NW_@N86\eTgU@G?QcM>XDc?#+ZV0I0^Aa+M6:1g7..SGKLNQN5)T\
617bGG6H]0<Sac@Y7AEV<V4ZD=F)2#/(X6PGC^M>9>4T5>6E8Z8?JMf(a:)Tc[;4
)9gUb^T<.c4AH9MC_YPZL]-<D;A)afX=T9-#))M5^2HbAK>_2JS/^dHeD_,cSOf1
(-C::=1aNAe<5@/>9IUG&4MUR]+g:2<4Ma\B9<Fc@6d1NbH_]D0,0-EPY.cO07gX
.D09TIDZaf+9;J=C;c[JN4eQ,RR)P9<834f-M8RD?U3N)fO)7RWaAF@,]PcM0dON
e7L)WWAUQQ0R8_LK[=T^aYc7eMaRLOG7ZHa.4L1J\CfN,9b9FOA8.IG7>3A0SBd5
S_QWN>S3b.;/2dBHK<=>eK7bD(Xc27ff[0D-RHcT]_X_3YD-Ga.UaP?D-b562)EG
.R1@UVRUdP4_a\787PT[]FUH-6,cK2fcUH]6Ga<B05@#^dKMF31?1,9);GGV=6Y3
5N^WY5EQ#NEKOWdM]8d7adILG^NQQ68-K5]8BUHMaGOW)S(,AGO6GbZIVP09:;>f
X+/TdadU=ZRB-_G+-+[WbRN2/(XS-:W>KSGH/bP90f>D,T:1=D\W(b.&79)7\\)5
#5)OB0PWU<f5O,#?+5+/Z8<NCQeK(,MLVWYTQ\1V>>Sg9B<>Sc0d2@T0)Eb^>d_^
?0K&@:_TfBUU/:[aff=e4YS=bO/RHD^U@5]8#2S<12d?=Me\=O.]<;FW]<<8]B\,
Pgc#WDO?JGH:R\aI@)E35S8KP-2dIZX63.D#[(AB=cF_@#PG1KD4H<[TQEP/&PF[
4T5BJ9X3?+,6Z;FMJZ4eb[JX29O9R/aYCaO.;eBAG[\.=#>cY:UA8M/7D]<\.Fc2
V9gM8LZ52TaQ1E.U2K4B^K_4(8253WVB;KZVf0-)TUfVQbWU[f1e>6AXJ1)V1\cG
&6EeOXaD]>f;IPLSfG7X&8J;E[Kf#8C>\L&447&01PV]#PP1X>9TRebBXg&/g:;R
Q^g0\R6/PFcLYVebGg)3)BKY3TVYO6-Q4/&F-=@^][K^(5E_SDM@&TFM#+,H#M)f
2VYc<C3>)FET?#LZ5E,<XBPWZK[TM9)G<?CU2^FQ(S[<9.#(W:+TACT(D0NFLG;\
)O6Y<8UEE>QZbWBMM<+^XXfJUU9CBe&&9^_P,1eA-MW<5WY)JFN^O>W]TA3K,^g,
.7F1]&,K98e:U\S^dL6RU.F^bL.,6X=O9-JD.,)R[DV:7bPHbgNU7J#9B8-GNKDM
J9H+V@FQR6Q2A/4;_8+C:fQ+Z\J([N4:K41^=;0P3]I&#&]7c\+-T.fIU]^JQK60
9,d1&,0S+Z.DfF-EJ<FY&2F6DFe>RH-7d4^Y((3R94QA\#]U/-_RSNc17\Z&R@BC
5W5>L^65=D90dF=A\-0(HDY]9X2G@/eMFV1[R)0bZd+>4^C=\1T5EdY^;RCU_b83
,@]QZ)2WZ:P[L_#P;:(Q4?B[/eK;W8R>][9#VB>NB?ecGF6P?N.Y?SVJF7C(2\C9
e:0NVZ1B:QU+GPX@2H;aT#a>Y3,bMACg9Mgb^,#2NL9WLYUfbJ1J197R85G/8&\L
=K@Mc/?HRM6;4@.6>,]M\d]J1=:9#HST#X=RdR)14#0467STICWg845R,P7?YU+W
T\:ZG#F([WNWOML/AA5c65Uc#V#>]QD?;M#.PgWA>V-L4JQ-O^<S,>_UP#O^3?^M
cc\bK6W9P.4GP59CfR+/OdW2VGI2;Kbb[60DcJ?1aa5-C0c=eI0g<>]K\:2(HJ.Z
.#9d&D5J5=(cU#A,HPP^c9FbU+/WW72e_<AD^B2PM2M01>2Y9JQ?>dF9c^86D(QO
CD>SRY0(_M#5)g^dQHCAVN2W&ELe#>WG<Y^&5,X#V:^I@+AE(SE;R68E4-Eggc1X
+6:47O:6-?;ND#DP44R#E--SG#QJ[]S?LdJM)LFdQ>0b@23GXP(1L+FeN;Pf(Q8D
/>2AZ\I-C[g6@XS=L\c_g<MLPSRVR[=>#a_H<FALF]X+ccbSVIU4U#06;7QUF6+S
eS?TR7J]N<UdFf.DE0\8;KYe6#@-dQ>CO[E,>]P8?&D.TOUaZEU(<=BZPVJ0ZO<L
FH>Q<K5:fa^e(Ee055F&>,3BdGM<T86e2.N^<ON72V^<ND93ED2)27dGLD7<9aD5
7@M_212JP&gJ9Y7@[I=]R;@TP/)Z9&4\EU<I)M5TT4cWFG8,S/)R<MV:^a+<d;Y^
b@6SABS7:/+G]_R+7D(R-0H8c8V<XU^5;G)_^:T/YUC./&Y.:K9g:NfcMJbHDIPO
.ERW.0;c5T#SfZG<La/YgKf88QZ>>@g<H3DG3f3/##EL4#@_)6V0AdQMMK19VI95
c3?Z9OU=e\Od)N/PYTK#)J+Qg5S94VYE2&143+_D5J6F5?f)>beS1+=YCAK]f69c
_MYRT.fcW6<K)bFL?I0Y)gg.a]6][O/-c_837Z-]\D+8P).&b(7YE4?OELcEW>@6
0?&HHD;V+96AQJ&(8a0_<Ic,TB:f&_;69MTO=<ae\US#/(c_G0KD:X5G)5f7=-ID
LC4JX/5X:[/IWS6U^R2HU#FB9AR2e7EH7EW8EFF:NaKRKK+?#,KYG;3(I9Z544Fd
XbB3+&3KVaD^4_2]H[J\LA1]2-a[@N^RdTd[+S,(J]Y^3>Z56[g[dcW\7+R0fC\(
c&54Uf+HWG\:08EP?CZ>7ZS<>.+ag@1G+TWQMC_?_-7\@<dPB5F9eKP-2J]IdJ3C
)0FT(S8(QDZ6ID#5N\g-932a8XXNRZ.;4,6RBEAI8&IWRF_e:(1Y<-G(^eA:8]\M
S,AA3deC7c:Pf9=X.Q(74(M()gUU#ART]=CJ6VYGJF04FM(,-X,I(8FG.UdN5@#:
B/LYY-GBP7DEXZOXdPB<<aJNJU>^I+S[fc@P3?Hcd4gg[3IE@2T\28@9<]A2=g8/
bT#VKX\^R0ZBEIN6#Y2#a0g\55YKG&W3GC<ID(&LXR?Z68QSW11H\C]M\&gX/0Q@
6U[_4L2F6[1c2Uf>eM-]g(C900@T=<1Wd)&aC&.,BP5V^1\UW+\A26Q]@I(6TMH^
U[AT,IS<,;NP)<2Z)?+gF\T)4H>f?NCO87Kd@\V@O<fGa-O-1d_IfOSM/5d;9QdC
eI7W,(g_\g<^fdW+g&T2E(3UNMeG=-8WWUQc+U<]a,9cd(0Z?_G@6\3C:8fM+9Dd
5E#/G=Oc1J?f\W_W;:-NLC7=-Fc176#_:3&DAc5c-X.4.P<0&^RS9J\KT4#OZZ>1
ZX]V)FYD/):@1fb2730cRE^J_P<?GL_DQJLS,70;39QS.<:_:db#K,BgJE_=>0bS
Ge-Zg[bL+ba(Bc\d1f:4MERe[,D;IOKWaYY1NE#_3;T[E#caAUQYHFG,I[_eLX12
;59MZW0RZ_Ze,;-.@\HC#ULPU9P@QCX0HOLIB3&D>V[MAA>_Y=AW\L.P<Y)I9+[]
3C:4OeRAYe+JX)-XF__9?+VRM6O;#0gV86BYLb-L7e?+Kg\8E.FQE_=D7#Sfd^UW
/6<?6cJHDAQf_Q(c19PX+C4.EG33B\6QFF-MO,XW7,;4I]Ug#/Z0<Xf-T4]LN;fY
3:RO<5UB-?L6<1]86(,108>d;B)(HW2NBTE&g+L.gO+CF?Z4f3HeHc;RAJ:d;\X]
I.HOJ&YF8&b8ZC8QQ.HMB4MF=X#,+S=eC;d;_M@Z:@O2,S]1[,gX63ON?LNO4<WF
=>?[U^6/dDf77J&,DD&>&7LP6))(RGFFJg0:TNR^E,ZALJ/ZHbKX9RMU-;Z<FGdE
6+I5GV?^S[5H(gL9fT[TP=?4A8->_Rd]M,Hf8Pf+RY6\Q8fYP/8[EBHa\gT./W#C
.B65SBNI\J/=BU;XD0VI&IW7P.//:)<UG<HB54:2Jda_:5)23gBEc,W@-R&R(:?)
IT24Ze9;7gC,P;a?dF(1=O_3,SLRZED]>&e:(HPO5fO9?ISM@XIO1>#aMSEg,JYQ
JI@1-OCR<@[+aS&-IL&=G#\]3314aGX[I,##P6Da6WPEPa&5P?X\ZcLGL,?84gY#
+6X6/_a6)R7fA@-UZ.-<64=OFP91Q(c?@(f4@W?>:KVO5C#RKE2,0.2R,/P^Z46N
c?+@=90#--K[RK?C;_&HM2#d\QJT0A>,[Cf7Q19A2B_g[R;<9eE+EYb[XB.bVLDZ
Z(:SA.ME9N<e893,J,Q-/f(/)QHO6aBS<1NRNg8PgQKaM7^+_LGL/21R<MG?/L8#
S]\VfP48M@HK<Z5JA.\d:;K,aF#.M^4JE;FKRbSIcX3JG>,.4XXX)_bBLJDf2Pb[
V4<NcWH\?.23]151+_KP2W3R=F5#;E8@#.1^6U^Q+RMbAEW0]eEP?(#Q2OO:FCJN
N3Y77A;^E:N<\bJ?=dAc7bKML+fPHf,1,CPU@XC6QDd>8ANZI<C_<O+G3W323DU+
8Q[KC(0E1-Z^W(69[K9_O3H67g91LP3GH[HX:5#[;5V<A-d==9<1872cd//EagSH
U@eTDD;LA_MPIQP-.)-5R:Oa9N9W1bUJ3ZS-BQO3bQJHWPGC2d;?<O/D0GSXD0:P
Zg14G,Dg,9&J&_U4a6[F?-\CL54&.O0e(_Z/a=KQ8N+RFXXR2H49..0]N:aeC.ON
LG2GJ8:0fZ@@_9.9U\86@^M1N-XBZ80eK^<CW#1^K,1JLW3bf)Z;D>2QOVLO34?W
AKPSJKI,a(?BZ=:Y&FE4e5F:N&aUOfAF7=:NbB[&Y)J2H])N-GcQMS.I?ZC<VE]B
J@Ag#5H5S.;&@Z4J]?4)a1Cd6X5D3:628.T7X-<JKYQ+32Z\?]b1^JT)RF96=J.T
(XG3@Q7H_4U-2[2#]ELY9a_O5FGQS+f&d;cbN[I8aK/6/228SZR/gc0V8&VVd^V.
IR41SAVL2>Qg:&ZYa:<^C6@\WQM)3H+6R-)6#>\F?)F84RKG29OPF5],O(/ASH/A
CR:6:b/Fb,DJA&9/HVdL/-QL]0fXB1JcLa2EG\&-/Y?@^6ceadSY2C3La&S.aKZK
&AUI:<+7C1c(M<c?QGHNV6/^<L51CeV0NCa^e--.-F6E/U>M>8bf)O<6M7J84C]a
a@NaW][4#XHYN1fQX<5IV/[M<@EC]f7bFA/f/cN9[I/C1B5L74<E097T;6=X#?-@
&fA4CY31cf+8<F@WG@DM-9JO)HEc5;gB#SWG@5OV5S5Fb&<@J\d?+g_B1d5L\-eO
U?_MI#J+\Ve6W2EYX[MJb9a,;D5@K=JKAF9&,CU]7d1\U)I<cE=@B=D?P(&12N0S
TWHd[J,QVN+c]KV:\L)#bbNU)]a#28)NPG\RKN=&P?L]WZ\OA1Pf7R+dS;eG<BHR
[<a6IBTOBaSHe51Bf:]=I>?=,QOPg[_We9PIFAVa7S^0?U.3?9S.AWFQN.TXS#DY
g^/@EaFd3,(4Y#JV4YE@#L\IQgR-f04]NQ-81Oef+D1W/.]O0MH@Ff5V.PT?,:c/
eA;75f=+][b9.&f9X&KGU6@MZ?2@eb91+:gb2c832b<Od6RL/@86(KBNC(CLF+/P
V90cgE<7M=QOQI=_dWfXRMB1UE.=/52U+HNI<<-Q4F@9gE48dO&XAMX6OYZ4F)1Q
C:28DEVHfN,K03d3]+HFfRRHA<WgaYPba1aT+8I=cT1:LG/51QATLCULP\UVQ9d(
.X/:_(-BCRe@]//Od(6EdgBNX\Nfb56V2FL\ASfI]L=EK\P1W+4_(3^.8\0DL:.9
H1.\RQZ?SdZa0bPd.9,&.TIeQ<&PSL95aHURZ<f&U]egVH3U-[\E6VG@^gWI,+OO
<Q;Y7?DCVfcbgb-.G3GVdJGKYa>K91L&JR60J;?A=E(SE69;VREZ_3Ig^RY.XFc+
3FZ@2:4g/O[Sf>3FIAPRLE@1CA)DZNE-G;cYD18TAZ2QPDfKbRV@TA22[J8QL0gX
1R736B_B9U,6cB^0/KCM3#_&YG-Jf9:CJeeTFNW>_&(gQaKQaeFCS;J;)Z#?fTS3
7(Eb+<WD0A3/&DQ(Jf:6UUFegMb/LOg4eY.aDSZE#RTT+S(4[C1&aLCM39/M#8/0
L@8;ME)RWZNMG9E=HC<D=.6U-F[T]1KX2[f),Ad)C,W9+U^IS&eTP]2gV8Cc=6gg
8HU/T/LXSfJ_,3RRK3,ebB:PIaPNE2YRNbcZM6?6U+Sc4bJR,a<;<W,9OZJ[K4)D
?V6W-=9>8D]#<PXBdFV1O:ZS<2+:S9][a_//ZP1?2#.b+970bGRL<IX#bWO.W0>E
D6QR[ARaC>DU4Y<bg-dJ.7;F1FA4_Ae-7e5Sa-e3QPD5W4aKU9P>3HE6[+2aW?5Z
UUe10\F^F8&:K>Acb.:cD<,,\f9__BIf#]QGGDf9?Q+d5)K#7f0K)^X<&g<SUD9_
CF_>-XK1Wb])f_9)P^M2:U&,&-K;a#<cKOL[SM5Nd^V1P]8>J/:&N3Ke;J,:FMeb
VJVU3-X:&3?/PN<8?5dKQK#[UP4SN5[,fG\<d.+<bNCK?>L#L(OQ\^&JdVJ@LM(f
=.[ReV]NAR64=8aPYId,F).8CX@U61)RPE?3+D;bcfZTUX&JJ1Y4dVHJ?a<:+S3c
JC#3V;(3F<:1Ea.BNYUO]N.E;a,\S6_^,A./\R7YV5A0?[UGBM9#a;2;9PV;#8PV
[&UQ=+SBI5D]?K[,edB;5BEWPKD&-IEaVX,\0+Tf7KDgPIFK9T2SYY6_B7/&cH2Z
&eJ5e8LSI0GUJgF5TgGWWHVP?/>)bO4,)^H(RI2Ce=9.fd\8#\,G6J)\AY79T_)b
1O?06>FI#ICfNAH6:@87M140;ccF1.e3FJeaS+SZ.L]96[SAbVOY9]N,^+XOc#W9
:QC\27DPZT<)D5<J50cf42.d48B8Q_D^8:fNE&/.5PfJEe_(Y;WTW<ZV,,d5H4T#
-Y,;(4f4[]7Uc)1I<b1b0#5^__<HXW<\5WJOX;.:.\&5Ka3Vg3e;@3<TP+Y[PNRC
1.(=-)[CHL4<969<1+J5L05b,^Wb1bI/I\A_=([XQScD8RIB:.(02FF6A>C[O3CF
f)-8_KH#>WPU9SQK-b#&e?cEFH;#QU6;DYZX3DDD+0/PH?1C#,)Y16]aR-EUNWA6
PM\1FYLBd;]a;K)T.;VL3#2(SLQC?d(:J^)bQe7A+d>bV#d11T0B36-MO>E2D,5;
H/8KX+49U?AfJ8-WUWSE/#&K:)_H[f?HI98M_,<UA8KWM8;)XB<Z7ZX^6,?NfU20
22D#1bEK1PV+CBYK,IXBCX<(E)@0/[M5b0TRNWLV3[8+9\b]:?D6_BH-Mf2,fO-&
KFPF)4_V0O-N.L<fY>#23];(T_:fE4?,EP[<9<P6<U]2[G6JeF_L92bMFEWH[:0<
9#/-)=?Z@JD=?XQ-a2ICGf_<QJ0CCD6G9=4^(a]83]c<f^D_YY#f#eYa(B^1^4ZW
;2d^0Y9LX\c(=NF5(I^&8LK\LEQSYR4-N,41\?JUfDf//M.I><.3IUPX6WJ.N3\K
f2DdZ0CcN()-[:(4e/+\V/]3/KNK)]<)AMI_/DW4W;Rb@AXdN@Uc5+/R1@N-BNJ,
\bf=dPSgE9NOgI(@(?OdQC77MaN690ReE)D_1f24fedTEA4+.^c6/S4L5B[fJ\-#
7\Ta)G2F526F/_\LY.)Q1Q>B=[dLTRag[fF_UJJg[E,d:RK<d?[d9P)X^F&f__0#
Y/b.L=PUP#_<2E5g4TQg6?K2:7:390S^a_:VU&JJ;^.)_0[R4dGTaO]VJegPW[13
]ADd6:VWcYWNX2?0bf1GI(88?PCL?;HCY3,PGd07E<O3d2aOgL(c/6Z(bIEE?[MC
Ng.5B7F<L9HDC@FLXf2I92d(9cD::N-JHBBP5FDKUG](;S2B6.VbZN6YJ<OP(a40
6eXNY11eaS9d_1EN5_J08F],,0Y81)Gg\H+(A;V>B;;Z=P;:F1.3GIJ4_/(:f@Ug
]8+NNac3?M#LE90454gU\83W^@E)G>&/@:WX&P+f-@ZS:MT/LIE=Y-H<6OC,==MO
UEV_XGIe\(^:(Oa=I\OVfbF?9?&QK:..f(,)#;DEV0ea/631;#VLHW@.U8\;?5K7
Q5[E),R\3X[RC1aAPPNY+L#SOY(8XD;:LYZBTV9WKP-2a9ed1<\[/RJfC)2M#Q<F
0=5_O-bLH38(QUg<]A[S2HZD,XG#K4aV;5^W0;QEQ,&ZK);.?&4N6N).I4<TaK3_
R[FJ?f0bC&M7U=XbZ55_WAbcWF?F,B6N/\:E6YQ^PQB9P[X7(e\&B>+>FQ&:>/U9
WcX6M][92;(5ME-QG#[QA)e0RDV9UZ3A&TdS(L=3:B6A)[YL)98I66+^+--^2==]
LEKYg>C(6ZU[:9V=T+@]I5)3fAO9V6KP_deQ>O8b/I=NT])+E?cS\>=^TAe,.0LC
LO][>FD&.C<7eA#<>:)[=7(bU+08#3=gg_LFG6c=>LGd>dWT+-(_f)FR?FX?XQYH
)F8aF.OgQEA9/H=/9EX+-eL5T05N#[^2B1LX[5f=Z,AYDF\E?H&8+Pc6c5EE@Y(E
F44<g&UZI=7-L(@E8VXW.)^&HfK+Z(g:bYB8GR.[6;cWI7Q0GcL>SX.8+?PEF2bN
W&/_P\676G4Z^.Ka&NW-S41;68_62N0I9Z0.2Q=e\1O#G7eccJPWa:6?CAY/JENf
5[Gf,X+-S&6(UFFL+[L]NSJ=U3K92eYVFJF>Z2cLT@@T&T&?,MMT@4K5g72,GEWI
>aRRe]Y957O2.XC0R,8b\4]\V]cSEQ;&8]E34gYB8)LU4OXO^\cEg/fHP=-[TI8K
;g>(ZIXEV&S>-4YLa=P<GB1.)/0<;.4>^YHYc9I-TDbP_VLM3?WBYI1K8^]+aG?-
d+J]@8d0CQQJ;^E/W/NF&?&2ELe(:F0X[4QXZ0N8>#]G=2dJcX;9^JD/6bVb+MDR
6+2D3P;Kb[XS@7L18@3U/,AP5EWL6D[\XADV&B8f,B48U1Q?R3X\5;S,G^T40GC3
FgU6/-K:/fDN^,;HaP[Hb@/#Z_WK3aT:ZBC1F]WcE],K7eI6JLdf4?e2:A<f7HGX
4c+2\WaO,;E-fPO.D8J5Nc;)dT[9M]@;F6#@GPXc31[]ODY\4E_3S5:OdX0N?=,2
Rf94FYLG0(/FT?3++fM+@=0^]&c1I7/\I0R84Ud#(IVHRSe&Q(D?0^Gfccgg^FEM
&aXd?(P_/SC&]1\QJ+=^ZHC_CK\]FXQP=@,e9C5f(5b=^_C?W)7-]9Q21b1eb7T/
M?S9L_ZcB><X8N(<PSF\ZI6KZ@c@7aXZDIN]>(Ue4,T>=P_=ZOO/a/=A)[FX@UOV
g12B_&aS/<KdQ<P,Q0a_1L;<_b;a1+Cf-WV-Q^QN(XT)7,CUMIO-FX2?E-YXM<R#
4E)UU3FZg?#NA[P(C,#DFW>1=03LMM#B<eF1d]UC:(S>0@@c=4&R)Y=<+ZX<c+U&
V3R-\aIP6B+7b+TS]-#d8Qa/B=(8LcL\PTEJ&&?O?c/(>X.UOUV2ZRfD9cJ(9eH@
+\1PE7b=C5Wa;?X4(Ua<I5<M,_H<IM#-16]XGNf;-Y9c/N9-.-J/dBCdI?-5&#&\
N29\RD?:#1P(L?MJ7FB#Ke7H#<^@)/?CERPdf7E3S9O#3D>8<?>JT].A[I:d9E;H
\>Y&<=[?N(Se>FO>?A&bPeWZU@GbZ3Yg0(dV4-7D[?V;:.9cb;U:<FBdQ0A)bPQO
N3daS7[5g6H^\2Hc.b/S5=5f]M,VG1IVJ1RZ\@RAcHAFfQeU7UAG)#[#YUa9#cgR
6QRG6BUd#+XS_F8RHE,8;_^/WFD&^A.)<(5;\aMX=N5f?+FLF8J\3NOV8_68<8;W
B\;G[96J3GMV0d-0]+aV)I5e5J-+&[W1_>\MJGS/&8&BY=(VBgfCJ+HIBM)J18>7
A6#[>0&:d+5:2FFaST--9&JT+^B4G)=\W-JbGTJddCKH/)VR=5cI_dGM^4OSO8?>
f&7Nb.Q0;PgEXZT^VePP(70V=UBWT[JN^T74/Z/>^OE9BXQ+1da5g=<Q2geXJ]R#
H?Sf-TCf1TJ:RDA-JUOV90HA4.BAYOKZa\>YO/B)S)F>M90f[-GIISNJK<^daXc,
eOAcDFWM>DYZZd>6X(9V-PY_IdCHQWDGI=:H;/2GdO:(9cfD37d45L9P_.0:B>5(
C?>-A,IcE+e5f?-D9<2#H>4+3g\EV&+aO4YU,^==/HE(P,Y->WZF/8W:XTe--f\\
R>;I(#Y9T@,,^22T.H>dHa;U/-M?f&R1c@Vg7UJGLc+NXQT.8B)_7MZ.^d7BFXX+
RGSW4+db#&YZ4[&5K-VgIga9ZcB(KX-:@3>&[fFJ)Z</4-<MFZM>NG&8,4K;/P4?
EY[K@g;;&+Ja?_W5O^40.RQ[fY9H,Le9QGAaY2APcAU6D^QbDR7NCU7Y)U37G9Q,
V<,<b5@3NT=.C40S<&e>1Z+F;_0f=J&2;cA<:]dVR].=M0a0L7/+C#B,X+GBRN#=
^:4)N@3<<eb._#B\-6E:#+B2N(dQ?HcJ2@5C42<+g]/3[K_WfggX22-S=-UX<4^<
>VaF,TVe9^93ZN9+)G\CD7^.]9HB<3LPB>IX?/EHF;MK)d_GS/FA/Qc9+dCV>OUN
Be==3Y9_eM+DM-8(UA[ef/Vg3IVX#c>&XdBWAc@T/c[50[-V6OBH[XIFC@)Q\NIg
VA>HF^R1?5e?L[=^B,b>\Va<N/XTF9a>>7RWfVP=E,.MaT4:4VYfaLGD44X5ODD/
DO^H-dJ695(CT;^5V._=HIG&W3Z_77(ECaKLb#K=UTY+)O,];:&fU4:McQ^][/C\
S(J(L3[ZA9ZFd;Bc3?;3F&S^U/6bVDe18<dQ:T>d58:.97#J4]J\,DfBfS9>\_Kd
7XW]S1I>4L+KL0V2-]2J>FfgWEI)d_8gS7F&R02.&AW&+LS):>c+#F?QJc\1QK+5
cDI42g9AH\4:T0f-RB_GY;W[fM8_MBZ9M5aP(\c^/)E@?B0/?>CU5ac3Ne?5?gXb
TC^U>fL;We\@#]6;,5G^IN(4^H9E4\;6K)CG>7A&&ZAF_R])<]7ONVAWG+1K::0H
?e[eSD]1gN)X)1;;^_,VUPgF7;e;#Vb<995W03>&__a>V613:T6:7cLQcb-TKGb[
\Bb4J).B-1addA6DN.>c>/#(?I0HQa1Y:KQ:&FA:>1;Vf+ZH64^,A]UP-21CT.KQ
;-+cC_DK3IS6_B4PK:(H02eEDgSEM-aONg9K/,J(WJJQd4B:29SJ?EZL(JCV/3,f
#0]9aYZXY(XVEKX50-S(XIQ,NH6&9/V:MPUMT,)5Rf3GN6OWeRWF>QNZ2P57@F79
e:JZ^]N:O)Oe,@0Z>K;H0?0:AAC=eB8AMB1bQ<G.ad6^W@c?FR7>EQ2)V:3FFWKP
\DaWE:f+VFLd\cC-VJPW<1PQdMQBI,24B1ZXB=9>TZET/TZdgPcY605B2f-W\#P4
B;H&>F:1&+(Hb+CXTURf&gc#)M-W?)55XK\a5)DXfbc3)S,O5XT3ZV#TGf0@7dK8
b0L(\_c-+6]K-TGRH12L5:)KNB@V7LK[[(NK2edRgB:Ia&_ZNU:MBGMT;SeQWDWd
P&/f.]=L/8b/_]SD,W9(0PEAb?58U8d.I&JFY3,gWaIF&(gFBDYV;2-_CTYbdGJO
E&5><N]0PcV?Q?,II6OM?WUP(A:3OO@O@3C-d4CT=E.3OV8PUHPBeVMQb[17BR\L
g95WHQ>@-Qa@B2^7=WY&I)EIIH0LX<5E?&3_;?1caX[Z::ZQ9R38Ybg9[Gf/&b5F
52/Le6bb108_fXHR2]F^?06dGY\[fMa:UI@8DZe>;0LdX7@ReA:-0LH6V>4H=VO:
LP591<Y,F+E;F^)RKN;23FIKKf<^C+W=_2BCD+K^d-d3gXgBFeDX\,F4YASIJ]X=
:e,+>#K1^I6IbWTFg><Yb#\,U9IT.Bg9N7g[X/3<b;-MSZN0@CK_L2Yd7[ZXND--
\6?-CNKQ_X-7._S/OKcAIZ-CFfEJFZX@H6OE^TFb4,J5-;,aW:GC0fGQ^8@2]R@=
]ES/WGAR,SA-e);^)K<851)?SVIQK;7?1UQJ@A[dP=:6:E6^ZCOMUc>^\c1L56fA
F5L1)GOLaN)F-@f6@[CO=,Xf0;59Ia>gF)@-XCUgaP\Y<^&g9#b@T?E?Wb@+ED=#
OSgQEKFVbJHQ(bgA>gT.M]M3(0GCKZY77I4cUEOc7X^d]TA4J1662\>P<M<RPg2H
/+-d>NOMMbeOKQ4WA/.J@?V?3SbY&#M&OF;7SYCO@S#9-FT+_Cc[4RXA@C_8NCR1
bIHTdgaM,.:1g4580G\0;R?3Z;GEZFHd&BUR](P;X@+LQV<Pf;R9f3]V#)W@V3-@
0#0K_N5)L+ZDJEFM1A^ZNZ2(ZF#IL;9HRY;^S.#;H?a[#<M-KBY98OM,>H&3BeV/
fTZP8R2:;81-Sb?6]@1X-^.::R4?dAM\AIG,cB8VZg8;ZN9d[3F.a.U&#11NJ0,\
E@)K\;(D=2MAT8908#@2_WRGU7AOd4#)c5B12&H)+C^Y]Y2>IDb6;Ma8YXMLR^Ff
:V\:.MY:/Z=7Y\MU8MOP+PH.LS6R1H>OK<g?K?Pdf6UW3G-2ZM&=UN,e+SCaOd:5
cN<NIJ4X9gL0LaX-U>Wd_;;_8..7Rg[#\^9:6?8(@XVIVU[B[SQ7^53X\HFE?e+[
U(5E[^3-(3T-c-@B:,H#98&(C_N>UPgg2PL^;TGGdH1BeR:B#]8]\=\ag@P)R)7S
c1(J8EA^NQcd2[BKC\^L@,d(7.C8:HP0&TZT9I)?4@<Y,94P(FJ>=D0LN;YBL9K+
??24&:>KI/V;HJTMN6CWCI>/B3LVT^gZf4/WU-(eOe:E].1Q+bd6LPTAC1Y\dS=;
0f18VeRG=^S2326,D02+LH8ALb2:@:\I7OS<5;cUJ34ebbOVD[SeMV])L7E>:A#)
+JbFH(L>;764ST(I/A1?_)K29\I+1N,&9?HR6?:]9RAL0@ffJ:[Bd+Hf,MI0dD>c
F;F[GABFS/PQCAFP5;S8PFC97\f#a2Z9fM;@&S0W-LOCN[>P9UUeJ3@D)M^YIP7/
aJ2XD.D>QM\M:Y=9+.(5T.O/E3]8DQP0&0V4G&;B;/X9+UY-5adM20BG1aN/V.;Q
#;Mb?H5K[Z.NW^0H_^.N1A+d0\)D;TGJ^.II/>A8BBICdD?L&.C4&g.P/E6;T_(P
0RH]BB^8=7UK/(OQUL&WKZ65]/Dfa3NKF2ANGc[R44D]A-LY2<PF6:;7V_R_+\OT
=C,#KX/M_&.7J+2)U=PH_TYPG>Q+c(X_fCX/3G1GWH_4;7OJcH2Z^\CE\A:&NSRR
M#00P@/Q.3X1CPePL2WWWGcY9gQHOT3P.2A3,P:H;4=G.#YI92E<<g<a(d.V#=)Z
1a1P21&9J-=XX;Z)1:]dV)UTTNXfeAQ5X?W6QgQYT@]ZYH86I\2c.gM3KS:K4)_+
TR18SLG?a;]T=1QDLAB@aM1M_;LM#YF:Q@bG0(B8)[A_A)7C+BN[+F+M/aEW91JP
J]14SMP6FfM#1-C_7B:V)NDTW40B29J+3[bTQ:@_(fI>^1RUA3YL0ZNg0C1=-.;f
N]IZ.?Yd\T5,O,b&^@HXTW/A#ECKFaJ^bD?W@UQ45U9#@^gM3SKX.2MKFfcGI?b+
),]CDfeFMNPe]IQg5CGJ>6L]@OI6KBEER\B<I+M0;9?WA#ZH1(NKX4\/@4W8>a@H
>-/RN,&JWQ7OSW7IWW.=?>dY-27eARNK7^[(@@(W5aE0:?O22?_V9>[G.]]C&OZM
]AES1;]VbIWC<6-8VdS<T<cP#6Dg:QbD7MD_3^CAZX14M57aUO#RZL4_?IKA>eFP
f:O(dd3?V?+-d07Q5DBMXCXaW&H_T6,4aMMAAPN1&N&6GGRGF+O]HSJ+LecN.EQ2
MJAJ9A#?4E]2A3O(&;]D1=(b[I73_Zd-RY@&4>&6f>EbP>gR#8N14Z=CB)ENCN&:
0c.1;K&d(U[1YRW.(BKBeeJ?]Z^a:;aBa2ZMb@dRf-:IZH+ZYB9DKEWZU42N>FeY
N#DB4M:KLAGR(Y6^M?UAG2<_c0HY\VTd/=5O)O&#f&F9N>dAfU3Da;&ILC+0EHG(
IaQ[SBd9X@#Y9VVRLfg#UUObKU_eI<M@eI_-d-(bHF:JPYT9-DC8CSZJJF4#g3]O
S=@fK-Dd;5&>YH2E>53_[[+(@fHd=G3RK1RUR?3^STNJYW?V4FK/LZ.A^c3_AQC-
3FORcL-])/R6b/OY\O29^)BXfEI(Y<Q&[LdX,2.Y)gHFP5(_4FH1CLIM:E.O,PR9
5@E95>^==IKeI;VK97.G;4E)7-U2/W9dcfaX;VUT:.5g,(J=e9OQ6A8#^?VB:cGY
>+L2C2@8S.5S;FK#cLD)O\@;)NZJgE3O2(W[Ia;)]6AHGd+&Me2XBKSI^4WSI@9V
LW<47W)+GZ68](eP\faP-gCB7=WI\;RYB^?a00F&5PSVJ&-MH:Zg=-7ZOQ-F(,?a
[-_NRHOXJ7U#7&Vde),V1Y\OTY<3\AJ&g99eT^-AaY;&BFNMJ]20SLG[Z91^#LMW
0Tf/4@7)&HACb9CdD^JL;/R0+d5+.QIJ54G7fG4QWN.E:(R#DJD42/XN3VC#=7VV
2ZA620<J.O?MKQ25I:AQO_:22XP-N[dXL.fbRK+>4[R8b8C_M((J99eKZVMG+aL?
WgL8;PO]gf2DU@Pa-_):4d:8b([BMLHWC3dS1G#NX,<:^Y.XQS,S)8M4(O[>P2>_
T7KVH/=+AcF.,3PSf&5;\^BbRI\4A6FME-TFK)QNKP(&7&a9Sc2TcFb_M=XXCWO<
U./Q1EPdA>0&@DOQ5SE_VK&EK30D;^0OIZ0G6=V:J#;&4T\1+U[>YXa/)ZKb0?J.
=41gcR5;W\D7[:#eL+H3cP)Oa^>UR5=6G?7+[;JddCZ1(cJ1Y00H^BbB79MVN.N#
-3Z(M17/NNI4cHILYIO7]]O_U\A0EF>Bb7f)1FIdS8T=>E5fZS]PXPg7U1-H=bYM
+]E1_ZIbW+HIG8.V6N&V6BH-db,JPYG.KHFcNf=V.1#EPV2+0]#23X,#5?RJ0WKX
4f]g9E()d983?9&N-e7VTX53A:b35gU^Fd<-^Q/ceV)bSXM;_>gDDSe(9Ga^;G5g
9.YOYNMC:J#>aEW73GE+cgM]UE:T>US4O0YFR?e@_Iff\Jc)1^&B8/2I-9ZK_&\B
bIK59)@cU^X#\X:&QMZFR9R?LZ@e\K(QQCCI4F=McVI@;M1;&;a:^RQ[/2L/VeI]
4VKfRMN>\53@,PBY3[/DDd&NV3KI&YQ0LfHNA.c_\f5\Y&CdDe1Q[:-B1:.D2]JQ
:49[ZN1L+:,95Z#)AUZ#Mgc[R)1)Ha,_GA&_U7gIZ1cLT3243d^.N8G0S9S]4OA_
e]S8)4)MA5VPB&EZ@H8WCB4NdOK40X)VBSQ68bRB-DOgHG#=[+ASK-gcLXf?\T[G
)_C]gdJGLDM+adJcA;QTfcU0\K\@JYKLKE;MAL0]KXeg/4CKUEc3JS5HeSKX0OKE
(-?20EcZD-XcJCG8E-@Q984]aR&>V(#]_f7WPb&R//O^\+(CL/+[A2QT+-(D2+#g
+QY3f5bZe?.?eDS/dAH0J5\GJF,ZZ-^@#;aK&\YfB]2Q@^L,?-gZ36Q9TAKdAB+:
NP^=dT;KA[?2X(=7<SIGET[,FVY(2<4BCg4WPB,VRY4X??C:--U^@abOS4S:AHCa
B-UW1a2F:TLDT_M,7FD;QCOW/Z5BP/M3N2;V8(&&>M_9<de&f)4_21YecWQd7Hf.
SHZ+?Qb([TJH8J9GOD1b#_SI4:a67)8Tf:Z2#3Oe.KE5C0cKHeVW/\YY+24+A#He
YYCMNKGUeaNZ,8W]/=WVEVWgQLAaBX,=,:(3^7\/:OQ__M>/e-A&#;1ef^2]YX5<
L/:6aWGd<J)[00U:?Fc0)\_U=5@JZa:C.C>JNgL:YDN8\2A,,<ZQ<D)&42G2@#FL
E=:O@Q?R3gSBHF7(-M^AS^CGT0e4]^BMWPKI82EcARR#L^M0L&<5C@La37+OXYK)
&-;-RJ3B0CWdS0@;5S[X=O]bB?OOCMbaNR@8D=:?YN(2-fJE(^Q^[&9_UWZS-[Mf
RB]-;f02DMb(RYP5F7&S+M&.HR&8>YEN<0BT-X1VaAPXA)7<#cEY^72A43T:b@@.
]V<6Z@B,7[3[?Yd7M&GLAfW76,M5?6H6+2=ceMOdH93+Eb6[N7-]IbO@MT&5=M[6
?HQK&-OcTPC_MLCC8+_FBF3B3&/OI_X1SSRcQgY7ZQSEIVLDRBXWX:,V-?<b0;NJ
eZDIFS_c2RcO6A(>;B9CcY6b]V^(8QY__-W;414=6UYK]\\<2<<0R5_)7/X89=cW
&JM_]9?M1cAc-4KU(F[8Y41;f82\bXG[5V)H)#>QZQA1V8PD?d=dHK]4,+_,JC4H
;TQA7fS_K/X(AG?&4P^UFRF]6RU37Ia9F#a1[\;gfX2EfV]>PGLI29NcR)\2F,PZ
1#H67&84S5_Ma?2(:D#W\E#S0e?\+4]GP^]W0JfAU?g^\:SJ-U>?M),D[7Ff>ZAH
CN2Hc6c=N]W56H&P@5G]XDGJdNIQ@AJ9SNY7b.Wef#C+(;2a0LdG7P=RE05:A40E
#8];]VZ<;d4I,,b>=2E36c0QR1#d:cX@WYcf;[]dIT8SE@.f6+JOO-fAXLT5bB<H
3@GZ\(-<0(D2:X<,,[U6SAB,4A:6Z_I+eXET,;e8c5>KI^5a9/Y45Vd()bS=YPI/
:MR;4#=fDeS0>WTHW)^L)6g#7F\cYQP9_UaY_DS_cB(B)ZTdN7&X^/^f[1/R<NYg
2BY,KBV^SZVbL30,KgLaa1Y\+?CeL=-:Af_Ec+RHO:4.-3AbWEEB.S(=YK;T[CB:
7&@S/+ZVaW5FfLf_#\K)E=[19a9a0[-&GCYK:F2L70MJPRG;Ca[c;0)_g5&]KFU0
BZaIQ:7CNeAR:Z.ET]A).L92+?<JdY76GYN,74IQc&7QAVAB,]TeJ\XOO)V[KZWM
dCfP,Q92OF\S)_I4^G4/10PA<UOE6Zad-JE-@GPV,\\X#fUQ,L>5[7.LX/WO\EWL
32C7e[.Bb[a+?XfYOI2gH8=O#Cbe23\g)=?(2;US#[UDc\/4+]aAND22Z7XUQO=9
g[[e8W.&#V_2OJa_6^6TN/8_O&VEg?0?gfMJQ]UbGVF]0C48W(TB?U?daWDL.6&G
:R3cM-F21F0;)Z1&3TMP-PAJKB+.G>-51CRRHdZ=6,:2c&15Z]_GOR^WRPBgIW+,
O#HEaBGK-/Sg>X_0VJ6TSPYO9VK#S[K)gQJ5_CaHIG]E5+4JZ3fO2g;HbH>RT@F.
=0QfF0:dQ@Q:K.CR<4bLJ(J0QS)K8+94(/Z[A<8b:+2-H73;>)&\T;OJ96#7;3F9
U<H6D&VFC#-AANE:JA4E57ceV)ZR4Z8@(+LYBAD<#ZU:R-+6e110WT[L^/&(0BW7
AJ9FVOLM<Q+ZFR?FL7>K.IL]C7FZ_YPL-72G81R#C<bb#Mf_V^#,c)(])CT2c(0W
4MP5:MMTN0X)FbH_OW[M5;TF?TZ@,TK<OUf)R;]VcU+F@6Z,H>#0D.XFARR/>\]Z
)]O85IPT7DNRIR&6Q?DW1(N?;PWQcg/P)8)F_]eg<G.URH\;cG1?dQBQ:E:Y(T4b
LMUa?T?Y6/aX6fV8:/<T-21[A-X\0/MHYHNLAb^I/B5S.I@5(#6/20OFU4.gXY1&
TL7\a3+\3AL9_HD)fG@L>Z>Sff4;)&:/#L?X>F3U>RK=?9XF2MOUPV4bT]5(QaK;
PWQK;-OW>-MQN.4=D8eJ+H=Q\9?daRM,)]&8Eg-:15WPU-Vae(.<,LJTPb(BN2^(
YZ-Ae2bP1=SGA-Z/W]_C\M]9eR@Ob9V?QQCTR/1GdVa_]]Z&PK9d>V3=N_G-)5PH
O=9a7W9F2/KA<DI<H#7\]2U.[DJY6:#FS&W_Rc)I<GOIH+?\fgFV^Qg7T^K@O1&(
WC=O;Bf,<P[V1adN=BTfMBY539:5&IbfM=&#FA4>?Z9;+WJcgJ&IK]]:5f?3>LK[
75Xb?#fMZbID[fA]/I654,#;\@c&M-9\G_/c)B5?&BHbA)JP\WUD01^0PbZA>fc^
HgU=K_fE\Y7B(357_J?^(WM[<0#Ed___]QYc26F/7:]J6:<<Xf_)/M;IWJ)U,?83
+J@N=#:P-T7Q1dXK8,#&3;/YFM1[24/ccZeJ)=a1IEcOB&^T_:XI9b[.L9,T>XY/
F@^=(0]Ef<LKR^g[SC^a,/(0SKCF07TbCLKS/L3-TaP:HL?]bG@YGH9V3T0GM^gM
X>]0(NCH9LD6e?=Sg9KZa:)gWN??#@NF\FNQcFS#X?@MFeA#5OcM>5.2f5HRY;c-
ZHdUNWQMV[M3@HD?gA=fc=D8?aUC:NFDD?-OX<1M#&_/)Ja-(DU_62Q4,U<a1d6(
;ONd^X)(G-LUdWg>cA6S_1?&I/-42+U(5BfUJ(c0P]BP(XAR:)[/eBJ3Ad^1<)0H
b/-50,;TQ?K2>OXR(?4/cKd[;P97BXWSB,Hc6a#ZKFDZgTJ[+I92QHN=+.d(SMLO
&S=6H)MQ6J+A^?_@G,)&T>_FI6;<//04>D])+ND30J8)9^M)[(/D2fRd2Y1.AbI^
^c>60WTMZb,6WefW]97e&2c0#<c_Z83)P.P>I&ARa&X+W4&@9/c7,WdW,6_5L2(&
6.3/ec1ON>;9\48#XV3UUP>:I0d/0-+/3-YId0<Bb0LY+,6K#^FP9b0V3SCDITBZ
TGIEW+F9LD\RK[M6HL^a8ETYENQR9RQB+#P+\aXLa0aL];QHcUKU^0g:d2^6LFE^
JF-5M0JF9cS45:SXNMg@6GRJV#31.VTMe1TT_0NR:^Rg4U[-IebV<,BEO:M[P(IN
VHA9H3NQ0MWd+A><+7X;e1?)6X&/D9#Z\G.fcPDUXO(=B:&2XOHR[IIHfDSA]OY[
Q+>?/S;3VHBO_,M,b79X+&W]F?AZXHQ;A6QZfR79<0Y@N<XS_05D.U,29=+\B#7>
;=.6/E3F4G##X7aPV#7^dd4=eNG4[RU9c/,eM+#&(\H[L+#P1,O+OZWMQQQ<B/MN
S1\)IK5d(64gLc8]B^YE,]_?HE:4.7^,+gP0cEa<A38YNNegEP^d-b[=Y+:SQ5^.
7K1/^^0U[9gBP9LTKAHM;ACLga;F30.df_K6E0^6FF&DeF>KAYEW-J)LMA/H#f?=
ce<.:a9N.\R.S.cU,-)?O(@K5\03TJg.6++]-#GT#S.Y)6NQU_Y;=c&<MTNL<>Cf
\@Y6.JI6_.<R>9#VCQSFB0e4@:JSQ8/)5Y:gGY69NAY.TLPA2KEO+[Z?JWa3C3g7
A13CQc>J7;CLJ2=YYaL.<0.:8//,:(8(U[7Dab^[cR;AG_H[P1QCFIX(8NSOX\G1
MYD/\=CQc-bNEEV&>=FF#?.)<:0fE)GJdZ&89X@-W>GAXe)W:Q;47.FRO8\44_6)
LOCU-;:F8:fC,L@#1GF5Y_M8>#Y>VM8X?[dL9#B6#04(F=Ydd0_IX\@^0/(?BXB,
BE8=A=(NeCE7U:D9N9=1DON1CQN^(0SDEeX(J^?0/DQ2DSDXf8]E^bB07ERQ8f7b
b(e3VZQ/5<=].gD:M,3TA\:/WO\DOO>c9>=&?1(/C(ECH0Wd-OJ5CF:^c2<Se<PH
3bPCHc#P&IIF2&EL;;PN1K=+\Z+c[74VQ:ZVE)e4cH+<X:4A#=95HTVK5Z_PLMHe
QSNJ9@6f2N1\CT=KIYLPV8aM]&[KJ>I\?K,C^+2FY3+9U.^:c=ME_f1ZgJG^cC])
G0)3:G19_KPcUZYMY^E,bQL9&LCKE2,#[?L(E1RJI_5Z2&&T]RO:=B\=;14S)H+9
g_:<D20c9F+4-?7Md2_ZdR-O?Y3]W=0,NLJ(,,9STC7YK[a^<a]Z/R#dI)ab\AK]
9GDP9/^=LbG32_dVa&8)GZ,-/fd>/F:K/U@WFg&Y_H@[M[:8(=0aX[Fa\QI-=cCT
F>@?Ne&V9c)-L6dNR&,,_c.Z7PP8&b[Ad=E2_>I3;F61&UWDc#+T2U;[a1]^d:WT
_5c\@gfda-HXQK.^URRU<TF)d^8H>-S13B2O(Q_;B9IR0(VV<dZ]W_2[Z.)04cK9
P24C&W[E,b>KU0UV@5B,<XQ9)6-Sb-#-#AEI?>6J4cRY-&+a3^Jd2BN7,V;IB/FI
-gZb@JOOU+0^][FW_>/#4L04D^M:bb3QU/>YcD\UYMa_.9g#7IWSe&K=?f>U#EdK
J6IT:RJ.+R]YBKB.EP9>W-PS4QC]g#c[eUEUR/PM^]K?JT:60+Y.a^X=)[(=;ZC@
[.VgMd29VFIZb(9?<P92.WEM;FPR5F.=M\EfO3:U1]/GE72>NfOH]IVY5ccG;^)(
39]K,YgWJI1)UATXVEbE([K+EUMYWdA]2cJS.57^HPccf?U&)@0gBF,+6DDF/SJ7
Q\McOG43GCGVMQH1WBJX^(Xc6-=5Q,1P:#H/.<5BfP9-PAWC1>T[(I9WgL24=PHI
HV4PXH818.fVSdKc./G-.J6=1g+O,d^U<C2,PM>F=;E)\O]>4KM;g7+DcMJg&L[d
A:CI?Kc[&F+M/e8dRY9XIQ3#(K/P(NN.=GTE\(96GA^MF&E_c7U3/#>ZaPB(](IS
C0@5Gd<1/f#MVUZD?eYE#>AZ<_-dBWUR.b>@1/QQ/_3(]eH)gZ4KPDGFLQ_)T_I.
1P[\1FN[fDP=agcg8D:FI;CN#547;1O<3AcEFf8+>27PA.H=ZZMXA>&d:)(?V.d5
E/E#=_UfZaZ_:)+M]^E\QJ^=/WH&LQ(#ceZJ@dWS^XA558Z0aDGY.@X((2N.cY;4
b&G(]5R_aP_f2KF_=N>KI8(R:&#3?[KZ670-EMT1W6A8A(XL497b(_X:f-A7cNYK
0T,>#^:f-ALSVbSaJgEQZXU=+^@>2U8]]=[[5VY03T)8bF,M/IbbKSRHH56OZ]Ie
=RCZ/O-bG8VN];ANXLfcc+2ZdCH0X/N)L,-1-[D/MdCaJa?81[G2LE3HLE8U5ZFT
SaF=5\47dTZ9D-dV1?A17@2a1BN#edE,-N5ecGfF5)X1KR.HP+;0SN^8)dYY)_#7
K;I+a16[+C&cK,>ZFH,MBb(X#MPF2[L07TcLQ=CTS7D.J8O^-0+,M62Q4RD;S8dG
#5,DO<T4QT:1g)#^b/YUXY:8E;DDPD/.IRX9/cU:IT2<-X6D&+723=)KE4(EM21d
W^_ZPOIbeA,=V;Q1B[&-W;4)-08Y#-SgFP9;]O8+>K^Z833[a6#\<FA5-XJ/,E7G
@9^X<NSW[<5MT+30+DOeb[LWI,=.-8]\(O+#:Ba9(=F/GJSbL#<HU8+HZ#<0M5+/
f_e56Q/[gP_9W+^;;.NI[Ga?-dMaAc\Qf8WeE(EX;HKPY.]6Mc1f,L^Wb086dQ+>
S]@L[]AT9eC85e#29LI=53CHK):#(R(8K[1)O^+C:V.^B0TD,R:T):gO:d[GRKIB
^QgNYK)a<,f_YQ.W@JcDg^aQFU(dH+&4RB_LeL0PM(JBO2aO87/=(VNWb^-ECQIU
a8.AGg)\_BXZX-[I,NH&S>D-O4HO2H8a7#2VA#\>)OZFSTDS8/SWb;J0V>8X=DI>
?8A20]66V88f1?RY=CgNaT[GH,cXW<0A,:?6[;T7GXTR70g,77W970e=#.U/ZP#_
]]=H9.72C/L-3^;_:1V&+4A\73<(6\:f1adE?O.3A@0@3;G1FIbIb7,Ia@Gd>@2)
4f.61/\WGYa^D)9f>F+G7NPNIeR[6Y:Pb0C(.=F5@M(DY0Z#II]Cc520(_C1Z+dL
,[Q[c5_:a0>WBW::=bUW\F(U4b@2db+<_<[1^>_a;1D=:g?@)+],_8^58(eZCGVR
5&HY(2#J[6#7]_N4a-&&(75R]gCQ4e1GW>[FW\\OgX3ST-Ye]ESF&1QMUF\aAf)Y
a;:N]WW/B\@&fS0&8MGDG@#Wa>AH8[aQ<S[8AW<_QDYL3BT&dLe&0M,XLTIY.^K#
6&AWH2LMWCS4Jb+G1R<+2(dFC8^5OX/EY7Q89??0U0JeQ/X>^#G3@WM1MI534I:c
fC,;,Z05D;GHbB]G+f_88AYR?9L_/1VF\K\e&@e;D40XA0cA_I;Z9)F8K\IH50O<
OXJ(WdWH;?/VC^\^b:NWd<2f\:;5(.W6=H;K=W1Aa)-@=TZ&JcO^Gg^19SKL8Z0T
&g]/DeK<a^-,W/HH93Jd1(.cK@c_G2X?VS-88#A-<a\^F(3P27P2aZTTZ25)M9@G
M97+TZWMNUgG-ZQc0RG((:>OP-dLV>Q+,-2:+.X&d^a8B1^H9AJ=,8TY,e-g-@^5
R4+edT@/?HHe,3fgXb>Q;UW^SG)YGDOW?;dcWU.1&NWU[0.0A4MXC1H@M&W)a:F9
E#<HbEHDO;JX>124E(HNT1VZR7f41[a0_DQLSCIT<dbYO?C;9_U;1-SN):-3D5.S
J\ECfIS&:.:Z0;&#GYW7<BCK-#cD7^UI2SUDIHUE<U>bON-R+Qf7N+7,=c?PBE5>
LgU;NN2F0W(;Z5P>4ALP>4OFZE@YS^Y/>-<](..U,0FcLRRP+TXO2SZNC,,_0R2(
WQZ;4D\<>P+5dNC)9.ScDS,-A&Y^GK7]4BJ2),IH@F=dH0G-0U7X#7^AM42;5R22
UM_c_<G3@<-Lf[:J,]RC[3^cXeAADH=G;IX<SfBTAS</<@4&eXJK-)0<Y^aUHQ6)
VaV-8R(fH<K/>X:A?J;>1X:&K6V8W]SCOf57H>bPGUK95W><)f^@gdP@-Pg#]AC4
aDNI6..]CS)+]@W^.;/=:H+RM9X59CVUS==bCM(bK7ZbW0FG-_OIGGcA[IL4[Qc^
Z)@,Jdfa-AB0U--2PGK6CfM>[W+V?-]6S=T6)_.@B<=M8WPUg9FBSVXU(0R=;M</
2O)5f4Z(]2L\/JVKF9c>KP^&D9=[U=.IX>]=g/-Z@=Vf/AD:e]?;PdT>A>MEL14,
Q:Z)LH#JQ3eZ=5P7fI&98[)\Q32ODRN=I&KIGZ5&fVEN)]EDMW&8Ff6=JURf4GP[
H:>&38E55;U[b.B280cHAT>Ic;-UH0U#_FO(6d2gI<9/(6>D6PZU&;COT9;2NYN3
O5T3_+bIedFGOL_.VN=C0T=RWG8#eEGKE3LTP&I@D9>f2RU]X5HU?g.HEYBgSELO
TMPcA:CE+d1\YZ;2X6K/2@?<#3]W9(fZ0^:FRY:gRRI8+FJRcK[9XgJbSCA\1/N:
34>e,HA=@1AJ[Md<]NCb=fPG]#MN)PX>XLHT+&D+R#LM9@F1C:ZFRN4-]K026ABD
GXRIJ9^3)ER<GRa1U()]RcEHE;?NMe<d47ZSdagd<,0D9-K;UKS_=?3^cZF>)P20
RT@HMTIG/?.22GBa=+4d1gDO3N-\f-Nb#JG70LM7@ODc4D5O.&9QN<KEaI;W4HfC
+Pc3TB:M6WL1Pb\7\V]Qd\K@2>00]Z9U4>WJM2JI@0;,<T1ad;4Q\W_;cg8G<;?C
X6PA+Ae:U]gN-d668+O<J]ULg+.,LMB8NA?08:FTA>^7LgN1Q)Ed>Ya-f:bY;(^6
d(-8;D=g#@X6/fS3KBHNJ@(ZYTNH?2C,Pg8+3452OG\:-(3TC<3C@g/):0K,5@(J
U@<YISESDJ0,1\R><c.&+V]f#/B:<2IX:H#U5A:^D<>P=O-A<eKMg6^CY;[36>@G
8@.P))/?+VR8&+<7PF2I/X9PI_O52R[<KHd1&RR:TXH@cDO2H)Og63JeUCP+Pe-2
UQO^-P@C+I]2IMFPZ8WE0K44U:Jde\>af#[96\3^<3U1U&)>5>UEIgBO2^-a-N=2
WQN@N5&=REEa[1-)UKZ(47F=N,>KVeV?B(VYEF[MdH.[I?RKeX5:T1eFVGZOcOQ-
;6dT2SZZ7IX1Y5;_LZ5ACKf+[_W6NbgV[.H+^R)H/W(_,a>CXG^=e>=aVB=RaPC>
)HIPPDZ6?0AGgT[WKU#)7>953QIO9_ON+@Z7gYS^.cR]&C?R]4b;U)R5FR/X,>@F
;-B0A96aOL4d+b[RINNEe2-Z<5(LeX7TCbE8g\9?Od_+<:^STCJLIP@_ABO:GZ7O
\#Z(5_cB:b6>?DN4L_71;7ZKP?+VI?b[W>.g16&+=Fc>[91W?P_)a#(9O8E6-XX/
/2e=X5g5797[PC;:RG(0c><WDO.SA7YdE;dRW=a\LFKX,NJc,DMJ56:<79#&+-?.
HN->?22F=(27W\CL<f<Qa\>4>:@MKU@\>MNaURdd+^;SX<a\X1U+:dRb4gR0GZ>.
=0E@Z_W=,.O:fd\5O\SfGBF<S:U<I&4]G(N.f.)8\J9&7?X3X8L4_W(AR:2Y@L#g
GQcSICTU-_,GVV+<@Gab8cbF;WG-Wa6)GV5C0<fJ.)(4[A\^RET\BGdF+P>F/9O[
U[K^gOENCb;4)K.O1eA3.FP28+A3?CNY_4d<\H#f\[57T-gNdLg0?=I8FO9=a0BX
CP5DK8OLWZF=GRM?[6fReUR@L?<9W8UMc\_N2^JQM>/?)(Z2W,8Q::2Q>(LCP^Q_
_]0d;<FB88YNWKVM-R7PXF&-A(6+)2c1/BbV:5P&7VNA[gI-N.S<P=]VEP8-WC4D
T)N-V&#VOUS#@X7BQecJI.E((AEb)aSJ9RK2#gcB86K6^JL8V5A-MZVNbE-<IYZU
BDP4e0BOHB&Q0_<Y<;2g[F:L^^KcBP6[\GJgY.]<_f^IA4C+I-P@O=E0Z4788E\5
b6JK1I>B3YU9NCgf;f\8W/R+d.^:,Bb,)J-7U9e9=&/9JDR?8a7Y6X_cY(>PXN:L
XT3H_ESI\^0F[1U(?e&+,;:((F/)NSI+L1YG=TK036/^0QP>]1ZH#GOL+H#DE<8K
80,O3SVY\4JQM@E22d(:YDXaHbP@JB>V0M_6OC-YTW_3:XZR?NCOJ@28aAQ[aeP1
9R6545cR&&,5DL6YK@?e&FcC0GS:O0<+:5^+[<3C2dSLMYQ9FP+#@7W1WQQfdW])
7L8.1.YLI0e6/&//@S&@HMB^G089Y-#4ggE(Q=4KV8\-\-&L>T457^.SY?WY?N3f
\##0Z?P@B1[ZLeL>2+eTG:HOHX9S1G5SF&g_U[Y8K]>:@gg(6^bO]Hc]I^GWGMXY
O&MGT5:0SP[+V14cIQ<0c&GAIH@^NJMJ5:;I7O_gfIFZ_R2HH3ALN062K#;2dW9/
72fX1=:-MCI[(P=Y4AIG.KHC#=PIC:.X^>C>NHH^fQ:7DG6#cU/OJ@Xf6dYJR3CH
f+<U#La-\/F3SYVX[]X1^G5_UAdV<a^/@M8QJZ+)S/85<#L4Q=d.;P1Rd]#U4@Ye
gFY[N>Y[.[cAgce)(_L<FV75^b>A@>N.1d\@2c@2:7QST1Z)a;F=1^^eF>VG#_6T
-]@A>c(=)48DX<D)=(2]Mc-93]VP2)c_QdGIJ@15,@2AC:K2@<G/V:J6<8>9RKTA
/;B>Q.I9SMS<g1V,Y][[1@6ACX4WJ+gZ8)CY)K<e1-SaXY2R+1L__S147d27Z#4P
gNcRY-H3bTMPJP+\WPR:[##X&W4#):40D(PBHP)6@>F,Vg^_I9LfH\08&R]&95\9
F=JP[]df_d[]W^^#=@T(H:GSWPHNYEXf3GTK+bY5H;R03/GgM0VU&]RBa?dZ<>I5
BHZRM0ZeTI)g]G4C,5>-?\KAaV9VCfQXF?I:J0.XRA7#T]ZVW+1(H7M.V;3@JeFI
dZUR&;gGb?gG9A7R776.L(QHPQZ[dY97(&:#3;B.^+GX,P:_/;#<?H6TT7@a>U=,
8?]^YEST\4XXQg)2L])1[;bVXc=WeE92#;OEb<928XNW^/NA/dA#KQR7J<d)9/Jf
[O6H\TAC=1f7/eCDH5]NUY?<NQeK@:fc;.PfYT4\bPOP4:)>;WGZcK]?1CS:Z(6I
UNK8.4[5D^.F2_bE_:G?UEa-ES.J\S;P9RNUNIBA;2;NbJX,Be??QT[;)FXbG;(g
-SCQ[fTFU2[;LK34OGWH-2^AK-&O&2SL0U[4W=#C(:d(-@TS0?0(3E^#KK?&aY#+
_JWg1EKBG+:V.=KW9]BSMbW]d)X<f]-fR?)@=XR1fJ8(M<9eT9),99<PU6df0#HR
D+>;C83AO#d6gYQRW0THN8b:^.A3Jg_A0bB,[4/UUUGS6FS^]QI+58bG38GPLCDW
0]^b\AfS-WbH;.aKR3-W(BNQHR0UZEKJ4UdXIF^?NWP(@=BB?V>UMdF[^#&b/-)7
cCBW83-:9/#4J#O(4:#@T[.IET7>[3:+2d)a7P:2FXWYXVgS?SSg)3eec;d-H<CD
2X[1HA])3MSb,EeWF&d3E7WfUIfG+G&V1cD@A1ZR8e38GVMc0(8>(H,1FIWP9D02
e>@CXT01_HAATeTRZU-\^0edCI.d2NPATAU^S,AQfVf.05?CGRALC^-/R)eA25>T
UTc(UBN7O6dD,RT=g4QaIg@BO/d]MH0aDG\[5EGX6(ZC54LH7gDWT[g004gUfNW5
)K0ZeB;9(?a&9FfXd9+ZeRKR90X85,]9fTQd3.UT#63(L@2>TWg=4&PF<PfL[MAS
)-RM-Z)2C8@TZ3R2).?c^cG@S@Q>MWB01,ff#-I8d6E1I5G.Qc\0gUQ7Ze6\Jd\8
(N7YQO6.0f+9dI)0J_CDNKZ(Fg80LD.99RaYZ.eG1#?U\^.WNK45)E(W:5,XWKYL
?N&d/HEKG3I?7&dKW(#IXeR/U7HY,TfgORAF>23f^#RW/]0f7Le.0@J49M\X7L6Y
OHa>&P;b7K,gXV.GEP&aANL;Qb8R/S^NbOI++d)P))TgCWKH63Q1d0d)\Dd]^fW1
RL(-S,GMHO.04KQ+O)C9_F6I+GFQ,P>TJQZS_-Ka5S^ddT.GSbS:Ae4:<.JWfK_8
_246S>3FcQ,O02[F/TY5#/YaL0.5g?8Cde^092W>MF6&2YcDHH:<>(gBK;+I(N:>
OeN7SXI^QgAJPH(2N.dX]\7@S2Vb)0#5/6&f@\N,f4Eed361#J-:g_D)Q5CN+Xc3
?Qa,=]QT)1b[gH9_XF:DU?LK.QPc>XD1=M6MIK<TeOK-]T_TKMXUTA61AL9HMI:f
c1?J_D3]QfT7Za;:MYe@b9OB/6S26_3J;V?-OF)_\35A43NdDP+IDM[V/,8=\VX+
>;P2=Cc]NQ&3^VG[<W52,88B09O=).T4[K+:CWD7?-=cQG_:b?3/X]VF13?/0D]U
d<GT.9I5OHRMLLI\Vc8US_&510[IPN5gW]_<O^4SWSFf&6\-,cKY((G4P_HZ,)NF
D.R1PL13J\/U9=AY(D;8]/<6CDUA/.:2>LPJSP]>FN2AM](e8OI_7ZQcG;Z0>?ab
_9c#F:=ZUdU7ggCQ/?b91SY0K#<A&R[+ZE;9]7)HB\BS#daR6gZ6S,)E.\NXM@e?
-KcP8KYC-YXf@(M<4gbC-.#R1\)81_IaYfW)YJaYMQ_O-&96PEePN@N7>;C/W,7W
&K:1;,89[K]CMWY/Gg.7XV7PZfA(c9P9O5a.HH#YGd;CY-Q6WJ/WT>1HYc^3(92X
>X=.c^.BSNXD_WB>M8[#S(PRa,0^c8GbCC@QR72=;RZVU63SFc9+c3M#:+e24X2B
V:5UM4Pa>8Y,\LL)e409cJ3;)-L;7O;e:-Z:<(5I95b>[TE9;EEc<FCCII,5(=;@
8_a-F+,XJW\(:a8D3=81UZ.UZfC<<(81U:aW3]H<V(ZKJI6.1A^,3)\cb&Ie3\S)
LCW#NYY)=6Z4bSQ96/ASU?JTI3TV)#@2FB4@]SOH?P0)(]3ad2fM,dOQMU5E802#
>:8=FT6FUEZe8B:E(_P>e;#CGAJVcdS)1J33<YC:3^Q#aAd^Z;WYCI^EBORBIP[[
=e?/,g5>c+8@?TX)2N+g5(E.,K[M6&F51J.\fSS@(L^/AW(8b@HVa/JGZOD#19TX
cRD@4@]HUU>Da;5V&Y>0I2K;P1X#H.4C7cY1THKbWH_88c9)a9+>^/_@)HKS6Q.2
)M=;[V(G(W6a]SA<abT?>4&N\7g3B@P5.fCOEQZ\RB45T[CH;Q.^?=DFZ&Ge@GbL
GP#Xb[X<N_#g]P3Pd-O3;WBQgB[J&d/56UP0)a3T@THGYfde^Dc0?-9U_:E3ZAV[
)D5]#ee/C=;,?cbP\<S60ga9A3ZQ/X[VAKI45)OXG^)#\6LbGG)b=C&dHA1E6.e,
2,S(DLFb+3e9&DgL53+]W)W4RBRUY>Ia7?4BJ1K:?=JVZ),?\>_5\?gOKgRc51X=
,M3V)UJ^?]6/M(6,c>B83D[DHL&_Y@_aSJ2feWL8R::IF[d26=Q;=S^F@YZgSTcJ
CY3O\X+Z]c2_eZEU0_4R@L1eXJ)Y1T:VH4Y#G/L#7G1g/cD[_@]U]>a,CPQD1T&&
G,fF<6\)7BW,TAL_]G\HB5^K,,e0Ce7L\W()cD3Xd_UFR7W<ZXH>5/VdD9Q_5eab
C]X8&PD06Xg2cQc;gEH4,UGaOP.JBTdHMcB<\bE:HN,-_\](D]K,e54,df)H4S-g
CXJ8PL)>=5gZW55IRXP&Cc==_1#F8#[fYX:-TL4.,U,J5e0#aFGMI;EP:X[4N2E2
W(V9>520RX@-.6UO\D=bMdgdE,=e8?S[8V+9.TbMIH8D8LGGMK7(G+73DJ^,J7+&
:J#f>A=56F)[F(@[>[a6[<IeZ4+#<Y51e2X]6EXNNITcGXb0:WD,3F0AU5(^D3C0
[Y17P4B>P+>]f,a^cS(0VG7TWD0.&6bQXeJP=@_5F>(Y:K>4^#N&U]T<b)FgA,=K
E8.Q##:5c2UZ:I-4)](ME1D:W55:^Gb:+[Y+7\:RXGV-2dNG#-:2\2ZfL/?.5K8M
e=fV5RL;9X^@5P?YDbY)d/<Wc@-L)X4:d)@M^Q0T&7_W1O<13Y,+NGQLQQ4:eJb4
B,3c#+.TXd7AM-;;/0O40dP:b:2NP7KTH83eCU]0J=LaP8,a]#?YB[-87<-@.Ua_
@LcTcLf7dEcCDYT@4OM?E.:/2<9,>2cH:X@]^=6#fQ.d)31^)&#0IA0@G.BaZ@T:
=5b(;&J1bL-E4Y#]8>(bY#HOF.KLeB/a]+_d\2NEg:^17F/4FX:1I=TfJB;)(3IR
eF5fVV+^BC8b@ZfOc1=]5D^BMLg-4=8[33Q5ZS\OW[B\3P+Z^+9W]9>C^@Z,da6P
OVYK0IbA)3[Z,58>3;^H9?f58/K.EWJZU_&RCTB5]a>g3QP3:<aQJIgX76Eb^Vf?
FQ,g3+28LeF#N,V5a,Q(Obc1HU6dY+6(H?GfaNcZ]O&D[=MX_=1.RIQEMJ@L50>+
CT2<6N1HP)D\]K\?/I,^ddUADD]GGXcY)7U;;\cDJJ7F1ca#)a42]eX#<SU@F>?&
R+45O5-@RV,Cf0ETf<@>,HF45bTJJ-Ff.<-0OXCE;(EIZ8-,R&Aa7IDH;CO9)3Ad
8^8&R=8CF<RA2^bb4PcZ[>Bc?fd/9fFgbf[6eDS[E&YdF1YSRA1OX2KSc/QS)50T
M&[ZAT4C]\gFcI9+^MF8VAR2:&faXMQD?R47>S>GZ_=[E^ef:F?a&.M,+#=&#T(\
F=_?LJQdP8B8LVW+=MXIb-<Y>cF6B0)<?+7ceEVY+6RP,0/eAg)DfPIGM98\T?RB
.J+Qa-6U5#=[G[f8,QF8BO#IdDD.]JLZ.@6gbQUIJTJ0SM/g]cN],7K84?1&.=YS
T&K-S?[MK:1,cTXL(+a=_[6/M_AXd#;3?/&_F97V7=N#dY4c5,O,HF[.EaP>\;B&
8MJMO7FI+H^fVX1g8\Q<0-S4KD;J>.\]3K?I)XY3Y2UCY;CJ#LSAFOP^8CV).FDg
]:N&+0f#Q=;dA+AdAWP>PX(&+>FE@L36J]]_RTEG?cDU)_gf-(M0eX?_Va^&)Q4I
GK^F8HW1;g@S(Vc/9C>fUSVYCfeL3bcDC5Z^SJNT/1580^4LS\^1U(<Lcf=G:a;E
fI.ZLE.3H;aQ68Lf0KM<+MBZBg.K:Y1WWQNETf^EJGDA=BFY7824RB<YF)=3bH-Y
7IF^3QV993TW-_Mc80?gTEQ]g7)cRWGaH0).J8\@]SIZ>9-1=J/53;3_II.?baPb
.6LG:QSe36C->Vd0L9_[W6Z8)AY@HXegON[1FL8&O:#J]V^Z/9d8GVV1)&)]7DP&
YggIQ4[G_a[MJZE\TBgR<X:f<g<(+458b5_g30PKHH#YR+=G257WI6\eZOAO6aW=
.bP5@NUP1K.\5(G8=-Be&ZAG(@d:-:#Z<N:Z]J[T_1:7ebZg:bf\7=O7V>X3QFQL
a;8K2?>_4_<eeKFAHT+aOE6IP[]27-(VYIDN3]_ID,Og[#bDBYD95bfeT9=/=G:[
CaSYUb:13]A0/<R,WWM;FYeVZ0CP(+S^9?KP+_8B4,GA&A.O,g1J&)FfLI:7V@Q]
./\NI.H<E#);U-6Q50<ea)IR\Z(RLT=6F#g@,(f+^Rc,)0;13=VKCIK?db#Y7Z3:
HAL]gGTc@)TgM2g\V.\c(1AR2&)L,#,DBJ8\f<D\H2;5SNC.&>Z9QaHb+(c4V/[&
1/A?X.IA.cDHGBQ5=R60NeCE2RPXd^,Dg[eG<E9beCbL+QR1^NK+6GP;(aVf,K#;
U9JX:(L0aQ:_BKW6\Tg3F0@[_E.X;)/7dX2R2fG@He;O@FMY#JS@CX8Y\b(:Jac,
1^SU7IU3IG/6_<P?_IL\BB84e3^&1-(eAc#+8S3\Fa7FETZ^^0B&ZIH3W>M1ZU]A
-0869JHL@YNN_>@1G.?_e5dR[5<2=H0#LgR_[>f2[.&e8OU:6IIOU3@HcNeWH:[a
\ac-<,Kg\5V/g+8c],.2K:=3_]=?SYLJg7:.B.LMJQbZ_MF#(;bg,^dVaS(&2&Z?
5CIY[AUV)Z0-GQ]DcC)BIB^4H3B)VQ:0Q#O^fWdDg1S\CO>X_O6(_A?U.Mc2=\a3
<FO,+UQC,JOT-5/PdJFL94HX1HBJZLTSZcW/8@ZA-3YU@\(f;<O+\cW[9We2>-49
674IUPWZZ/TCC87KgCW?&ZaY]Z:T;05S1OO=D)8\fS>Zc#c9]gBJgLV+PM/OT/T?
9g0QY77YR)GG[BF_ZFLYX=6b]_a)e.^b#YI=12@2dQR4X5=fT_9?PO,3;bZ^Q,d3
^U<g]N4L/(>.X/9F=CMI#V=1)FIQ&#?-K2M=D>I-P,)X4?g1aD&_&1;_W>OKJ-W6
W7(fX6NT.^?fP0a#T/:-N))M:3Oa149#f)gTG5Z54^+G&H7-CC.B>A/+KEV85CXA
COg:Fd4\8;//;+XF8<DBZGeJ;2dO?LYF?5-]]]b<8.FC?a5K5L(F3,PP8-1NfDAH
,]2ZX/[58U9f\_)Q,/D:W[&4G(T&_S/Te,DJHZ1L^e1QY4^ObCZ:QXJG&R+6BV<^
DO)RXgB?2b34,-HXg87HVV<^],c3(BgEXTWK3V;&+MQ6AB)cN1.Pc8gW@eK7#LJb
8DDG0adea5[EGL]Mg7[LG#DH^9@&AQRSRJ^,+=@Z1?g[&8EBZ\D1H685F^9E;:40
L;OZBCCGb.7[GX)K<7dSCaR2IZ2CC86ga5bN.(L=bM[5H,6R)/YC?.7@d1R956Z<
KdE+[@#6-0+24MUcHXUA;T<QE0X,WgD-)J05cfEc^fF+f]>Sg?>>?O?5EB0#6]a&
M?G9?Ug\HMa2YBP480eZ<CP[;,8_8;[+^0#NO&bDfd^51B3;#E#N/dQEH2-aX1\1
1KT<5B];:HC3aa8+eL,22L##eC7aER4V,P8bHc2P/CKKP/b1NYJ?\>YXU]bG_g6<
BUdU;bA_Z)+:?/,RR?^SY023:T\LS#,#eM6[gbb0.DDd811I[I]Y7TU5g\+Z)W8A
2\83K<fBRTE4JIJK/cRL-ca,WTc_N^98SR_X?>184=XJ#?a.e#&4IJ^YXD_ORd<O
N6=bQDOYf4U:g0?<gSQV<cQDO8a0(L)fE;Z<^1Z[g1Mbb\822&74[)M/,OI6-cH,
_aD8J+ZbWYARd,fN2_)PN\+M??cA](8EZW[eZ9J;#XUgI/D4CYdZCPST[dVa(^6_
dWbL8DDA5,g<g,NE.,I4b,36H?A+^#J]C[(7+#Z1DM0O5S(D;=M\N]Mc82O)dUSQ
4B1M50M[+aBYAHEa;ea)+H5[8^H(/fAO\gXRW[-I:\SCZ^BJ(cbI\42A,ES)dOH8
GUE5843<ZQVYS1#fHRYIPR4:>61@fH]^;IJY5KN&@@(278,I=<QeU[I)D20AcP4O
?HEBTcGaLJOfJg;PeC^QJZCb_[UO,R([\@GG7(TDM=4)YVK=IFE_1.=96gX4#)4=
4Gf68)KMEJS.>PEE_Q3F8VLS0UbO7KRW<7C55228B<Xg-E5<R1W>aVYI8Q:U#R,W
OCYXZY;R5?d[XDO3&T>QYg_/&J?VSNbV#6<L@dUB0MX^Y[a1.ce0&d2d=1Z4=E2b
N]SX7PdQE>3X67Y4]M(SYe7<3b94SR\0R0WBA29L<d.=eY8f01VA7D[XTU4g6/0@
SJfW5:b:?0bH.XcS0M#@W>_cIMN?VeWPE.:+fM^fYQ-2.gCXW^V]=)7)O1]?,OW8
G[Fe,N=C-#FM&I#>;9J0DL0fO_5HTC(KTY,AF\IY+D;#AMbU3KQHG)VVgbeeD(+7
LMYNZ\>g:cGO==ZE_I.@V@2gA520([C#[.B0Mcd4K-9QUfND,3TGPe.ZgRWHGBg2
I/-E_egHVB=Xf+0@TUTO+e))UY[1ZLE_L<V/>FHW)/+G>DH]3Z,J0N2=gFe[Z;CX
^V&Sf3()@06@\+BQ;;:f=1TOg2Cb<f&[La:&3<-4V=&3bMSI0&T5.e8<S<-fN&dW
;CcD.Y&=S=1[;)Y>1Y>_,,_CLZN9B2NO5eT6:EXYALbbN/daS9+G-JX63--30Pff
:I5,7/7B1F&?IbCUY?cPC[];D0CKGGA+0A\J?2A))dCL=OG\b3K-V,FKG[OCYDRW
QWL1TTN8:-Z//<I3g<HAbC25KeY0;,8>]ZNY(JRNLQ1]6^<f(QG(0bFQ7bD-=QM(
EC];BJf9+-OS[#K\G>W.QM>6<0N@Q<&]\XEU;R4&I^M&Beg&LM\[E#;K8@H6ACOC
Y,SS\dNTUYAgVN[6,EPTa10H2+#?=<_^GcZA26QG))&6FS9UKEMEZL269,A>79Ee
GA0=0\;7d)4JQK)aG+ZT[O)T>+C@>V_,QT5[X#DW-?0R3V=V43_JQ3f4-?(9I0T[
ObU7TIMW((4A_.9/Q:-fa5FQS.0&b18R2=PVG,/GFNS<.aM/N_7YO6H@/02_;ZDe
TD5f<_YW:Nd\8-X9g_d7)?IGYFca&KG/^;L\;:FUMXU;CVM&FI+BMYALBg#OSZ@b
<FT(W[P7^D9SXN#Qa-J=)/dXe_+?L93L>SP(V<Wg#0?5UOegU]gEN?>4T<JJHg1X
B:fLCfX?GXf510CH2HV-\9OR4Yea>A&V=M<JVG1I_E30F,(CRZ38U1_J=H/>#Y0c
H6A?84365FZD]aTTZgG4\L7=_MT^c2YKS4.(cW#BZ_46/e69+(XVFN^\L7^LE.;/
94=?gTET&2SV(AM5Z@I1=2Ag[:acYG&VFASaY_aJ9K1fU3=RW=^,[CK28Z^L],P;
/M6T\3N8.fY[,&&(]KD)Q<O.QF0C/.2D8WH5_M.GI^HcQ5FJNLGMB,CYWTeJG;PH
K)3A2N:(cCJJVD8SHB5S#8Y9<VJ/>;I.X:N59;8DEQRQP.[JC9R33b1UbL>a87QL
dcDF;KAI5-c9^^-P5L1YPOa=^MY52EE5,:.1#]c^ZR7A.DEMNT)QJH\P.SBY7AW-
(WHF-3?QX.Ub@bJ/I0&X(&ER@=b2,-eNVR\N_1bP9d\IG#15KB@fW,=&6DBB=M@U
b.1&#M.GX(LPfUBY1S#Z8_Z,gZL#=+T[XRH[BT@K:L4P3:S4b:eaEI9ARcRcU\\Y
.W4[aTbV843&CP^5XH>V_cGTZZ[X@@>NC.Paa9\C>4,YG1;JUOOa[\2FaATU?P&H
IBMZK4V=_X8ZOB9LAD=</06dgL8M&;4^2?J?,ZQQ8Z@#8YcX)/=eZKH]DAC\?L@I
X\9^6)]#O:X27V9(VbAce;B=&?\ge;O<E?]R_9eR09#6+C]@e-XUM_9bK/b6Vg#6
ZXP,_M5I\e)1O\0g;\&S:)(I2SU0VfW2#(>O)d+NL]-Kfef]ZBX<TXad^2-O&Eb)
:V+cGeVdJ59[VSY<b+=94;#RfL],X-7?<>/fSfJJ0XTMX;K]WJX_cOF#7?3CY;?^
]E@M:KQCLRG^EY+F0d1)WCY#W8^S2,>8ddNffVAQJP=TNQ6EHF7fA9N_LBW:E>ZG
?#V#_))VU<B<3)cN)\W5TP]L-UfLMA[,MCH5@(feD@==\\O/TW7-LLK?eEAB3,Y>
Ce;+[A:A#TVYG<708Xc#0P]#ZA?2-W3XefN?T[Lc:01YT7aH05YZ;-gK?09a^ZX+
=A?)=.[,>EcXgW-EWM[fS5D1-Ybd(MDO[AO\FX&9@B8HONS947/>^:32=6]ZVK1W
(7]H(;GL-5U@TS9898Bf[P3++H-CG-E03Q[T(.R<Z@]6Zdc(33)F7^PLK36?/IO8
1,;2O]-:V^\V2TaQ(]50O^_0>9X::e;=FV@SbeBW>PfPTBVK&GB.5=I=DYZ.F,#7
/7PY0MC9WMX03aT_UZ^ID958I-FBDSKYV4Q/H)BQeD]\cYD5aIdHOK?K+O#b@78K
N^S2L315)e,b=V#3&WAc8I@R#DD@^AI;W[+7fK>JGK[1<FVgX9/V_g;SH<+[a<Xc
SP:45ecE>)_<9=.9[b-a\P2,E]XD668agA?I)Zd6K:IVV5V^Tf1\fd9,MfbN5N?2
P0K]J.Ie_4-U2DH\ff2@GZ3L0]UcBbU4JV\6LPZM#_79;@P@_WLeNK^^/[4B:__M
FCKfaWL6CW\W9,Ae5I.KK#K2\ea@IQJ(]L\-D6T72dT/f5HW(d1E49f:O_-BaB3[
T(W2TB..fVQ(:dM5+(8B[R_3.-2@ZVS#a]@COd9F6M&0Rge5I[F&O5P\GTPdEK/D
<I)XBEOMW?33;2Z)#aDMU<;gV.8LFb)/(V=]e8_LKee#))/2M].311/[.HJO+A\;
RPb2b<e5C9gR9:GGH)/c4CKY&,M:L0Y=POS(XFN/UPAcSBeVeV76)Y@VKG6&f\LG
:3@2WU))=^L^<@W=8UPUISgJEPEOY.?>;[?4/QE2<5dKFRM/Q1&66D^a\HU[@+WG
--acHE^bd;&>T9<9DRLPW?:_)\589\D18YR;+Sg:(fA&D6)eZ^D;+QWW-_L[D3Z@
X:,L/0.?X:A?OLCA_4L4>RENS<XaJfYA3[V?Ca?3_N<[])UIDED,P29L&fPc]]-a
JAYG11,W#Q>K59U6-47DIS)<H?De<7D7P65SEO,,;/Z-3X</^K[F&T\N/IJLO-dR
VAdQ8J6;6b;=[E>9(8cFA]2[IB=56g[\,T.LHZ5DaQE#L4VAg7dJ(0,_Of#X7-E6
<G\g;)QC/W@M-H5G)R8J1.RWSLTFT^U@Z]X,C=S.G&@:3@K70&cLPC9^_O0T#/XY
@=_^=GRWBY]#6G]0VXg#V.[#V-@9+Q5<R_b8Y0M#K/_JRPD9dTQNbUc;M5+3)RF6
bTKQS.#Fc^)\g0QGLUQLLO&.EE5YS0Y4ZaISD)6&caW5ge[/#Ia4KHD00>A6:#gC
ER;&2YX--J_?f1PI3UW;\2=+)F5(X5KP@M]Wd^R?3b1HQ97ALCJ]O/,-A8)VE?Dc
_[[U(5NQ/.>d8.eBcXgLYD<E/.GZagZQE0G@BQLGBWd1@=O[D8L/Za_7/XJL];&K
]MGdV@V67a-Qc5cg;O5E\:e+F(1Sgg&df.H3+K/Q0e_]8;JNJ+8(12MALEHHE,G\
SRJ8HG^DNX7fQ-d5P(3N#ePE.,R(5/\:JT[?O\]_Ad\WdNTR.YUEQ>X[6Nc3@]+\
[YI8PMZ1?4TbZO@XWG]K-ND^>GK_(103S:SS-_Y17,/XVP.UX0SNLY(0?6]Q-e_?
6-92),K57VTY3ONfX;bL:.bc?8J\8W8c(D.L\?_]P[:,fC-J:H(>aVCdL/=813PW
dN9b>37X@AMGT,5,#d(b?PJ:7X4[@]7)@b+T78&3g^&2YF9;V/K?P:+AYQSP+a>9
V1O#G_U3Pe[7KRJ#SOXNCa>GDO4H.>3>dZ76gC+\2N[Q7/28K.b+A2+W\.3Y=6,L
H:C6fV[Y@OM>N^6I?[/6UR^15+CEO5]RO5DeSDCE8Y3:5S5S]\U8HZ&#Rbb&b9.I
;0L,EP(;R@fDQJ)O6YOUNS@/YW7?D)dO>J[U]<@-\+Z+2:M=d,ZGgO8@d=F=HFGX
0<F-B9cPJY&_^])\a;XP_<P(8(/I-]]+P[&/c08B;L]]5?XK1(8^MLU+/S)-]8g(
Z\)]SWeD[/S_SaST2H/JRE.c8HVV12=FZ)SR<E.WPO[3#/\FZ^,7fK>J(IQa/P2=
PKHd0ODX:-PQ0e<)3\,XW;-C4@OS.N>Ff+E_5:>aMcB,5.VbG2OaDA_=<&g.AfA/
dA<&1#J=a7,P+SfUH5dcFf6+V=L>[e/.-GZ8SDRU80/[H2Z(>7WfVE+>@WB@?\>_
SdDS]eX?Z9N_3bX;A7YaV#86C-/X:gMb=IODL@=G[5Cc=0AWJ[@+_+G=Xe+3)\26
5ELI7[8d30GY()YE#gWL#PGBR^OOCa]I0cN92eN6IET<=cUN?-X)[0#L)[JXW?dQ
VPLQN0^=,M\T)=@.+Z(BcZ2HYNV.a,PC+RW/,10)(1GIY8H-P<I>[\gVDNfaQ1A?
VLY@g,V^JIG(B)>XJJa+@d<,^20CSd52_/#P?>d<_JT)Q+0Z?Z;WeL]M^;34U+O=
(._ZWXfQTELZ2aLQ,,[OR92491]cET+PH3dTH3RW@f>69Y>ZV-^c5dK/2.FIS4b6
NX-G1PH,FY#K^d<ZaJMLE^.8047S@Y(;(gP0e_.=WV+7F?Q<PDP?aFS5W+dSX8E0
,Z=bQGOZ[\\I<NDXOYQG\ERO2+c<E)e,>^TGM3O0GQ8T_f7\d,5MR.DfUeC\^3e&
QHH04L55J5HF32O:5]Q6;-XISNLDa7_b-,SXXEDR)SCDL1FgH(UT6N].TUH;D+IG
1d)7DaLKd^GZGC9bQQbTePLL):CX2G^)@_L0YPP:7IW^J#H(EK?)MbQMO[_D^FIQ
\23P9e?7SG2b;C43P?]Q)(TaWCK4(QWT<9E258EM9KdXC,9[eJLd5AV-R32XZ<P\
;XaBU^[<B,I^-R?(Pb^,/[PJWG+9K(:-JDQ9aVNE4(fdb)@3H^9#/X5J,_TC>TNG
DM5N>@5Lc3_O54S<V>S[QJ?X<LG<,KUSUHF48R4QfFG<O]3<6-,?@^9SL5@N2BT)
Q4S<+.94ML_-Ffg9d7;\14U5)0eg6Y4ccZX7;G2aB>Je^B94Z>HLf)IY;4Z@B]V&
4_#g3W.9285&aI&W+[U_.=^6MEV7O?T0R+)<>b<=_])N5;1>\R+?1O\Q[O<7:OMV
PM=I&51QG@J:N=C\KYTHGXdJ;EHfU?#[ND\b_^3IFCc]8DLPY./A:e3)E5R_)LZg
b+/1O688361GM<P-c]:PAKUB>1UH9USB&[:b3R(NCHIW1MdF-24&.VUSO=-27#<N
\I3?e+M#^HcW)PbBY:53\,[U&_S<6NffD2+g(Uf)-g/]?PBcK=D4b7g,0eJLM6Ed
I+CT:8(KPa@b:gd^9_gL[?Aee\W;JWNP#e==KOU=70a=S3cR+?d6Ye1b5^Z1fYA,
70IJOc<)G0Q=CBH+Q;-eA@+NZe?[:X)\e]>S8dQTNSHXO\R79GIKHID_2G[#P(Y;
((Z)dMH/@(ZMc@>A+5GZ++JNdXGD;3?c]Q>b1D+HFF+UXNA\-YLC7_^=+SE&B]Xa
BQ.f0\2fRJ=9VO.D.H?&LUFSU:R9:WL,M-CS#C,=:R9cGSI5PEaAbNFdQ[?,,(IH
KP_ad_1-V:^L^CQ/ZfA4>ML8.]J\M?C#9(e5M\.b8XT))KAX9;A10L6U_:<=0<\S
[WX2<9SWRfLP^U2T66.KLQZ>::1ZGf5J;Rf?=G_UFZ)CX2E,[V.#1^;4K48EU;1^
\TeL_2-.B#C\#EN&(0H0:L+(Ne,QETb7>M7GEJ4?O5dS1+/#>W.eXF8FRf@QD#LH
,+>8&Z\I(-#QE#&NRZ^VF0RWP)2fe7Z\1?CNT+[.ODAfE79V],-3K-@T-P)CZ8T3
7/2?<-.R[;=-f=>G06IKP_98;CSLBY1-9<d-),K-dF:FEPAYZ9>c6G77=04[;8KJ
R0WW^Y;HY<Ae+ce5G7:\/;1d@BA9P#8N0f./)IF+/7R0Z[J1/5TKPVT4-R[>4c8a
4c.S>^N2UfY(aN,A)?g15WL[?I[R@A>CB(eXc,CdB=#IFD:K^5O5L3-e9/_2+b@d
.&[H9:VTYMLK_0Qf#S,d91,U\Pg=:KPeAX\aUg\V_V,YJ12MV3=GB,^Kb:JT&0<]
@5MZ93G,ReKPQ_FOKZ3^8>&\gO]JTASS2^PY-4^[fdgB+RZT(X[Uf.H###^3\Z9H
A//TR;1K>#DEe(89WKf_WVb2?0=D_MG6(Sc+VbVJfO_#aV(GUc5YN.PJO]L[N:D;
Yc8;K,]BY6>3=b8>UXO?fD8C(?dL3LSY?5YH,D=ccQ1UEZ+F=JVTfb&ACfgf<)5Z
f.,P?(@QP20Nc]M6<@H[M^59(#_8+a@)(0KS2Y(XCS;XC\Heg0)@d;=d&(IFQX:+
Ebd7]&Z-><(aAeIbe59XE#K)+03G398g/C_4?J0LH72K6OE&Xd;-Y/I.UY/IbaP7
b(R8,N:)<a;)L-^a0S>=gXKOBV4]CADBa=ede9<gYc[_L?Z@8J+8UHR2M9;1[DOV
[g:M\+81dY(-0OHD.HAR<AS#/+_OPd,P&Qc#_9dIf]3dT+)7?BD)=Z)J>@4Y6QI_
Cf6JPSJ=PMWUg55d\D&JV>a2PQ.R-BDMe(>D-cMC;Y54\.=\>c-75X)Od]?YIM5C
B,,V922[P;5K?fIY[WRP3,&O;FGM->IR=,=4+PFIe([/9ZKAEBK?a5(?#eZ?_e6?
5B=0gd?,5a=E#-#;3CNb20/:c>8PDRI362aAddBW(N@9T7EU3UX7:SGO:ZeXdU(,
8bL[A</Z?IPNM,.7N6)V\Cd-EA&>Fa&52F(caJNb)d((1ZPg).-A.ECU-\39/cRY
U>POWaJ)CZ?]cVcXVOISRe9Q]I4:3]?XZc20VWR-+G,(gTAU_LS/Oe2_?_+:3c;C
7Vg)e?+W?[LP[QQGe7SX?&^[CFELQ^K/a]f)>(ET\FNA/+#fPc8\:/JWBXC/)0Q>
URL,@Z;L,Ua/EE:[31H=ELK2:D,KV.WD;NMQa>P0f4Q5OE66@?:d;bM]NR@6KKWB
^:PV-<:GJF(YE[C-KBJgR+HNaVC3]2B9bPYGB?@,.&&3D?1bL2ZKU]8eGIeMPV;O
cM,X?77BSUa3@PO^4&YE[MM2U47gSH+?Q<RL9;NS97WPQ,:KeHN4RK<J;JI++bU4
f^&<=>P-g_6+H&F3MU.<f]E-?;3_^g2)<QKa5,MR3bORB;:1__L][GU,UJ9[\/Xg
2TUV^>.V7e4AD;OHLf-dA<JW37B#C/AEfJ7O<H+.YC.WQLWNSdOL_=0OC(KBA7L-
[4G82J/E;[S&f9#C./VNA5_)@-Y=Q2C6HPYH(_CLI&^JcUCY+<-V[WG(bB>VJ,-Z
NcfaB#=Q^X1cg7,H2A;.2U+KV:)R?fYDN#c5.Y9+/IeT:9&)314CWV_=(f_>:D8O
,aL2.NFYAbCUPE&YMOc4V:LU6b,>C@ad=[DfS7c2(ON7H&LF(BEJ;MfD4,9\^N1O
#J5HF=SG(+^/JWgASRM33,gNXVg?4b,0GBg-e5Y.65XK[]4+5#NfATISP[<6Q63\
_?VQ[/T>Y4Z_4eNKTHHBJf0>\GYd?JY/MBgEF>C)^[=Y7>3cR)NDE)JOD../cC5?
T27:bJQfG.;O6F./g\^>;H3)_aB@1]KX&PD;A&M+7Q,U(\LV9bN7DR3W8?@Qd,\Q
4+OR#TV>L>(9W^21d,L8g7>e\.ZN=A9Ta_F.?g7+2L^P/\V>WfC4Sg2C_U@_d?B)
Rg&Wb@@)N_/fX4@A1K#1H5.[G/Y&-WN_7[IGYgKOVK@JU.]/C\/#XXNGL;[^IVK4
A.][)<A[?HcSK<DW0?.XVMW7R+Z:)dab._Y^JGe/.?b73DCK76P)gaI-#c]72c3_
&&W]FFH(:g>30B0ZU]-1Z5<BJ/C()\E9\E.G19QBD>+C9+XX;#(e7<XX4M6C&.PC
M&W)R[SQ1O3<O>F?C7)IB.N5<b=_^P>URe(+-+WP9XAJ=DSFK9@PbQ[<M87]UP@[
5e^H8TZU7YRVB#U@IJJ0g8PYX,];=_5AW+2<.FK2LV0K_G[,BK1/0/R.Z=W@?WE?
A[-aJ1)<-ZGY,>I\^JU.Y2UF,,BU&+cGD\:U2A9@RF6?DeBK6;.6e[-Cc10a5f?T
#S&H_+D^PcabHU&=8a1aBB.Q]HO^cV4M_Ge#:V;fMFH\SY90?/4,\Y_gLYe[(MX=
2#R5[-C-a_V<H3H2)^K)dRQ+=^RI?SA>[-7cffOA?e[eT,[SG#[DR_Y^c]\>WFLC
gY0M=.8,??a7STIZ_VX9Z41c.+_H@/\KU66,8)ZM:<O_32<=@FL^ZQT#K4))gD7R
NRcO9FX#L&?F]_GK>CJD6/,bYZN9:VgeRa\;7D6P>\ZK>gg=27bdG?RA)G@WOY><
\(3\A[/\-c+EY<=+#37/>?cQ6eP<@&K<\0XEFdI,EEPA95(VIa>>QM6R&.=F_P4C
1M6]OR?X-Q5c]==H-ZPf9&]S&W<A(2KXJGIJ.Y_gJA]+@-)\^@FV6&JMFTY##;L#
VUQUH-<1HaQ51K[@T=T7g_&BdPMK8AW2N\ET)f=R8)ZeZU6&Kd#V>YJ6a)5I_6IL
14K@955cWEd8].@E<-DQ,<#3\A+dX@MV85,.R13K?0.W:^c<[6PQ9)R,&X./5A.e
NdcPMS.\Z;N@ET(A,E)32Q0WeV=H79D03?<6C6eC.8#NJI?2Db.6ceF8SYeG&ePF
478_7IW?+1[QOgY&RBD7,a)O+J#Q)RdI^>d4Z08S]#f]aCZ=R#P=^EZY4)G0&(2L
Z.#)D7-gG;?\d#NK=+6Yd;5JMdNQF6EPFYVXUTY?,RYS^.DgE\9]9F,7^b.(+SF=
I-/8J^WIfLI_>;cW<d2;Q(QfOW/9,-G[GdP[Q]Z,)d#\<=gg3HMDSL<.Va+dK?:9
XOF.IGc,PEUO\/CU\6SZ-)858>2VNg7I6^4#T0RaL9A4R?ObATV-VMd@4CXeH.d4
I0<^X6?PAF1(;R+BHWUX#b<(3aDa?9OD87J](Y4PE3.;6ODf0..@fDSY=@JGAWUT
\+K6^\U=??05?,/W#OFV7^0NCT@Sbc?/g7E3FP\dOJJWM/cg+9CYOEKQ;O;28?cI
;N[FVBD\/G?H0R7IfAG(3/@b,W=JADdQQ=.A?.),EaQZ\./7@<>1\Z&_S)Lff/B<
Pe)gb&UH0)H=-CQIOc(2:\0>6N99^?/DJLE]?c3]Mg0J8HOWdgVKa=QVD6E-eLS9
;SVRN2Q:(S6D(4;Lg3L:Kb)];K.UI2^OUK6d3RaR]C)(BIKR<A3X3VFVg@IO(ZC@
eD:QENI\gP6/7P;P\Z=K?6(/#=0g5Yb/TS&R^U2\\Kf^(g36dP0^DGY^#BB\MNMC
Q7cH52BABa(MRc\Q:<EN0A,^ac.DHdPcfFLQ]FO0RH8LVC3:=<@3V/ZM+.:43B+[
CA)DM5fWBPS=7/-U6b_D+2[<=93b=;[]JRbgZ)]8VVd6e;[W45^-eFQ4+7I&OZa>
Q^bJ(CLDa0Wd0KFD@#b6?^UN5SJ]Y.Y9aZ3[a\TTPX:/;-IO(Q#e)?);.S=dc+B-
ag3f#AQX4CF5D(BPA#A)8R5LQZK-VZaF=eN^U@NZX>]OBeV(Nf++^_c&N>33UQ&g
B/>@a.IZLWG?C[;BMY]5d^WHP&b6d^JVG<DN<0e7DDP:GRNLW]3<fFgUK.dSBLR_
?MU(+Ja8[Z2Da(6-/bPPDaBW^Y<Lc)_YF?QC75:cDUgT:(7ca?8HN^;PJ@J7;V3H
@:V<M3f[0.gHggF(,J:5?[XX_(JE1:da_6#JOZ()?+Bg:@SG-FfS_R:)>+BWKP63
\c\OG_Q+9OIKL[MX[=b)R+U[)C]</_;C;gQHbF,QL50KF<L#T?>)Q[LJ(]D1_-b+
@e2K3VK_D>Z@[ROZ=\M8J?Q4&-0,f24(dX,8E\S^).:&\IFe<PT+Y\c3G.72d0BI
cC)^<B2bB-EeW>2M-&\H8\)KFKMV^XYaV5/H)L:6e&b1OQH,EKU+,1GXc_Vb9]M;
61K+[,9Ud)D7QaB2?WA?J,FLc?FfF:3AgaUX_HVGQO=^[d)<1QcH3=edNf:BZ&8/
3BW658(0^X&1/K_(,E#_:Nca.H&T.U2g^\.2D<B>IBJ<04#[/HSDdAY5KYFZJ,_L
5<J/8RW;XJ;YbO.5B;&0#f1c&1@_W7)K7+J20db>U^T^WED.(S/eBN:<V7<1eb8X
W/_9gc@S_J.:/ML,AT+71e]Lefc]>fGe._WE^YLF1ZeAe/I5NP-FIe(A,SG9J0UV
3[a9.aVMaH5RB<EeXfUfL#-OBbA\fQ_B=EZNP>&,GeH=4N=]31]>AL@]DYQ]CGDP
Y.7bJ4P><)Rf+A=5X13T9[7OEf#667]UBLaaZ0V3[EF=2cBSeH&cP-SA(P[R5S99
N<:/8Q&)+ISfdQ6+]&U?BSORC_#Q]X=>b;-HFTFC54BFS#a#EN5&B&_JEF[=\2W1
Eg5DZJ1L)<+C>a:M28._dQaST_;.UaQQ^b#WJ17;@#)EEH78+GYcAgg5S2fZb5c;
[N=I9>7Y-\+\BW+HPE6ACG]@dM=HRITJ5?S/VUc@RLN+X2R#c>/7C_R:LF(?BLC@
CbM78C[A>c=_@EfYQ)6)#eCOGg@b9GV/6;b^/Y@FfeA^_]SIHg[QK&>I1<8JVH3P
-Q;.1[LcJ2PXIU/\ORHODI<e\ZTWMJ;:dVW6ULSGVZEJVGNTG.e_XH\V,+e,4</S
OLICAA182O3<;c?JRDOVa/]+MKTW[PGOb@@T_92U&YQ[Z^=TaZ^@dC[+V,,5#g?U
&N9(CO:\dZAM,9c#fF:^_+.<BbB3>BL&]+8d<RU&/c.6\R2_8X(5aP7d&]DNGTM<
@K)#g_W,__BOYY]46Wd6M=6+R@ZH:)9=MVCP@G:(>ZA8b>9\c&?<C?JYD\<HW;[L
d,2b/28bY.,YM4G:)[8Za3X.IFGNEd-DPQ0#X;)Z\gFSgFY_V)4Ca@fT]?J7V;Jg
6V2N_g1,D0f6^5<9+/Y.#aRDf.SC,+-d[08bMMX[T>_XX(1_21&QH:BfG77gbNZX
R/\UU1XJG<OUdaHZca4#6Q039Qd?+S]7T7Fa4J,E;[6Y/A#_Rf(bU,@(W]]-?J7R
]>7g(VHI5g3JB8&W[DP5)Z<+GG348?b:I5QgX<^,SD;,FP&];@0GeKA&7M?X8ff-
WXc)UV^RL9VFM]],EM(:K/GOI#4NSVVV\fJ;S)[K?MUQIce)<1^PeREOd5f3P8d8
a0&Z,g5T(_C5,IYXRWNKS=N7K]76A>&;R-Mg76N&Y_KIT.PO,+Z2<M7Z)Ub.&_Y&
T.L_e.R_9QJ4M?M^e<G:2/X=Z);-Wd1:#NcG(c+Y>60/FQeg>T_/IJbT48H:e(;M
dW/>H#]?K0M:<J1:c0/_/<B5H\g.@>+CH2Od#XVbYQ\VVNc\eO/:L^@_WSX4/3R=
F#<,UT;-W\XZ8S0Og7c#]cAgPc5NYRBU4NF@A\.?G65;_Z=),;a21AU?Y(-]-7ZZ
:Z.Q_\+X4gaKaR5OeAg]>VD6bW-Kb/YU\C^NB152JKefM[R1P<^@IB247:I7T2S.
<dca(PK)S@N50HXOCP8O-MAEJ6UT0F80;7,_^BVJ\ed/FMbBXZaYTI00_2/=&b6W
WLP?O00J;_GEb29gbE_W?&-]M>(DJBJU&Og#[d#QILW7XA\<.N3)AE#.C\3\E-/Q
>AVIedU.P4Jef3Da\d]QdF9(WZ[K8SYW#.gH;.\J[]>.QF;6BB1g6/M1]L_ICTg-
L(7Pd2R.>MT3R-<3@f2+RL&&,OFGZK<D(RI)eP>V4-TD:d92SRe[FVU:?-PAK:I4
:@XX[LCV;Sa0(DSHYc5+]&Sb+CgV^8ZY>829>=:[+L1O;HP3O]N:2-PBDE:1f?LG
9dD.N^_>#Q,V^WVUAB)^APT143eUaJEB<N?c.4?G6(NcB?;c,QR]YDQ&@@#KgTF=
,C_<EMX/<-a5ZF3H11+]V;503S,HFe#13g(PY=V&=b)^f:<@M.:DHT-MM3QC_4;0
eB_=.;XDaMc#X8_DND&P6R,BOb894;H-?^#P,T@PbL09WXGK8UON6d.eZ/JbQ,B@
.BV6E.Q/3Of\/]LFB.?F7PA)HKD?9>7[Q0Z=,IH2?/]=H)YB4ECgBZ-VX^-aEZWY
0@3W>=+=UX+61IDY5O4_=C<@]/g&a:<gV_Nb4_ONR:_+#^ZW]1KC^SaJJIA[ZgOg
E:+0^7(L&1A0QCM,/B)eGV?@\IL?SgL3PBLBJ/ddG,N0f/_N].KbY-&_ET&HK_B_
Eg=Ac7L.#F^Wg)MHJ)V+1.>6MGa@<.geNe3(]H?@M\W8KBY[NV7550fb(+L(]_)g
O>F\SbDd@K#_S308BSY81+7L3.>.L6I(La2.D(SdY0DJ+@f:c3/.O8ND-\g.E81b
eCE&)86)A4EJ7NeCT,Q7=J>E7<]:Y:?.+I/-W^;4U3.C]Scc3@D_V(_RG4-O6g8C
9_UX2108>+-FSeZeg\Xe(WADe&gV-5UdG(+1GLN+WA38TGEf;J]VQcXG.g+RC/[P
<gaW\GN#?WZL)V6=Q<B,,gS/RMH(T&JU4=,0[YB\;+C0O/D7<;\f]f,S5Zd2?gE>
Y,LI/V[_(f\2I[L1QA:QUCX>ODC\05Rd]dZ/)BHXeKI9fIBA+TDOa.3AIQCf75)-
.e;EKb:D[g:f)V,BD>OB/K,_b[]9=Ec@d0d;f;d;0#5#<&9/^U]DD7gdBWCL+1KE
CRJG=f\)F]PgNHZRdRAVR90MN8FU:+O8.BY6I-UI5b29O5U3WS9FSO@9)9>]=a@;
f68Sa^aRf>&Geb[CDf:_c\>NY#PIUMMgNP+dZNAf,RfJeb\ZQcfOZ:ec/;DJ0QT#
b\_aW-V-FfGY4dT25aE2X\[;9&J^V-VW>K<,b<=dfVZf,6AFFA30a5]RSWKG#GXB
G@XH[c>Y/X(THN]:A9]EP,>(ID5H=K8JQR=H+L)1DR(\8DfTAdN8)d?L&AO2ZQW3
MbHPA&LP0<[VfMEE#F/J96TU0Ge6gVe0<.Z=ZR3T]cc\d+9DZ9<g+T,dA\NbDPf>
7g406>QOFHFdF?>H\-^1L6NXN(^,b&C?Dg02(UbaX@1WMGVbdeJUeEWQC?+YJMU/
=H=[0^N#&R2K)G7<8NR?PHQ_g_E-@cY9/,)<96XLe(d7bR-4?<?+Q0QDH1,?5))4
-2=TWB/eb78)?26cb-[YObM-NLDE^aB;gJ61#.H+edcJ?ac[&II4.S^Y_7PF8;40
6cBCV@=a&O?6]<TW6MC)Q?a<RgY<^7ddAg9K_>BD7/]SL_8PHZ6RHX55cPN21M+Y
;Da,8GAU99\1;2C6Z;4T4(cU7^>bb&1Q)AMOcM>867)U\Zb\L)@UcZ+3_bP[5a=.
g=Z28C\V+8e9,gc==BBe(^Lb-&K:g&;97();FA[DWOcF9XE8&9eC;V6V(K)I@M:R
dU9^QC7?;X/LG74GN<6A8,Q)\K7OF;HM:K(]?A]1OH-Vg531e?V5MdM]YP^4GPI:
^MLf4HVQ<R0CEK(.7IL9F]T/+[.?+D8L[/G.+P-,X^de2U0LQ-^85720LI[[gAaf
ec\DQ)bfY+2F[G0D#(FC62L&;PBEMd.;Hf,IQD.LC95+6<69^[afe)1H)&L\?V7Q
EJ<7@024.-g,_-:&a+H,Y1KA)DZY-/<VMV2?9b;,^0eD84;@53=.V]2@W+P=0/#J
7#b>]G^@b4>g@>B-#^\[D.PZJcD@BB#=GC/SRZ,F_Dfa;?;[G0(YK=a5(0?MU@]K
6\;\9R54/./[=(R+TF5@<CSJC6;<6Y18Z?N9HLO^D-Y=Y?<&XF8BI#]c\<T5M5^?
+gZ_)\#LKC9^QcW+_:(VLDe5c_e<AAaA>;AeD76=-)HLNf9a[5Y@G4><_dD3)?MG
:9\d[VCb(,DTUNO>>.eUg9V[d8<X/[.I#[I-gN?<D&VV7cUQWDc3b?bK@e@,fZG&
/1\<<?]<_#/-ER\[&PK:8:2301f-VRC\:.&^F;4gP92X83FCHRW?6CH6M_TKJL2Z
<)&GgAW@VR51[--.>[-+O@#2IJQ<,GM#W&5+Ug?KeW.7I>4M(L),&-^[#GV05NPD
7(._X@PALM.ffIIJKJW>[aYW[g\Oa)[-LDcH8^VU/8.3^9?O]N\[L1=3E,9aE#d1
<-Uf#\NYD&b7-INZ7;P\[g^aUDA8FEU;Y^M]2<C1()KgH=7be5RW8W,?56f?\([W
0Mb;.fY<d.8g=:@+U)&CPeSB/dTW(S-Pc+(5d]U\;FE^a75A^]U0bZUJ/M(a(#_b
:52+e)VI(BT=8(,>A;ZbH2AAFF#0R9N#[fAf)dIN><U[):KcLSaeG[\(3NZRV;P>
>^Dc6U.D7:L3^c=O7B(FW[=a8SV7V#bdcJ>]V;5>S+Y&WYCYAR8RfO+^F]JdG2+Y
QB7?QE^#ZL+cBc>OH=K^C0_H.5CD]P2Nb)G>VW^3bIbgWUC[GR9YVMB_d-dGT236
SAMU/CR<7JLEgFFZg_H_#+HAWXR^,4;4T9.9YJI+U=>,]KAEW-JdE<1L_YG6PF]R
d>)fU;K7Dg#<^T,L#Z@+Q63Yb=FIKX,JZKE@Pg=LW6_c;GA;]HeT6:Y,dW:eTgZ-
2]=S4[+JV1B0CK,=H=]<4N)U>JHYR3\B5EG\Le/W>2&0=b\A=IN>@&SbJT/B#a0]
;J=K&?)KMAD^TLD];?1Z9e6_eag)()NSM2]D^e08)CB8=L[1;d<bR#F-A8L#GbJZ
&8X/;:79F<^:(E+Y0I^OJ6JDR#,+bge4(4D75&(LL^U.FIHeP__OL0.W?0e>6=WN
6adOHR_R8K&3,&:/YZ[O<#LG0S@;Yf+\effT+3,+g1:G>I>Ua),#2U8FUZbG<>#)
4[ER5aIX]g<a(B#0?fI(=J\c@K@2R#Z3dY_b(0[P\Z@f)=^KY7G[:CTZ>e7dROPM
&@22+F2+93=GNFTH6<W9dJe4Z4B6N+/01TRO@D&ICY@K@3;?:(SCPEWE&JV<[]=f
9]CU/_#;M/RA<63+OTKW.T/7g^<SOK6cT.>RRL1ag.U_P?=FK:-//?=/8f@Z<D\=
_B[\>4_N)SG9S@e-B48dcZA<D+O]NMDG)@C:.<9J)S:W#S4He]d_e+F[,_MK]FZ_
H7.Y11.0M,_VE#@^fETO#f./OIE(4Qa-DNQ>&b6B916I:J1d?3^Y6B9WWf@8P+?2
P6)?1AAI>I6V\HGg4OF<RALcB_#RAX)A)K<+^:faI2;\T,XH9d\,&gYdRAV:1IeS
>71L<4F\g8fBe/R,4B:aIP+PE/gMZ<&7MCU;gE4I9[YXD(6/6A(1(SGB(H8^8dD5
,-V8>;MR&?6&>/d+UB\LJdHTA5ac>)bAN:G\&TBH7fG@LM76F_KK_H&^#^_da;B>
C+ZG63><QNbDXgfgL0RCa,FH+#&e3BEN_B0N?5d+OX4K-eG)^:AF;.7LP_]Q4>@D
AV#bC&\g5bb9DaH&1PLBNC)QA>e^A;4Q/D3N^CC&3VNAccZXG3E?-PgL]-f\(.AY
@NZ#8O^TDE#D[db(S/M:^4^bSQCCK:H\@3BGQG@83D/U+aX_U3>(2\6+V0(VG4\:
N]?4;K92dD>(HW(DKd7eP+&&<f]\Ag60:e&GE2^dDQ9a+G@.-RQDG<2=VTF?>V_b
JHOJO=?2W+AG.H5aD^&UI1LcLMG7G3-:7\[D\GU[fU?F2R0/O>4-B?7AZ?\#SFd>
&Nb</,XI;G4F4R@9/?<IdG=d62YYcW+OfC_Hb6T/B=L:?LSJP;@I8895,2gKU\8[
A)/4eY6=<]K>0;9,VZKCdE25LXG]_PX1BM5fSYHQE5?3beJ)ffSDeU/Y2e6159Vc
,P#B+Q-f>+86<Z4,E#+\M_aR<1&:Vd,7-6:aQUg3#O?dU=<M>cb7Nf;MRNUP?2GR
?.XP72g0@Y)bY?e(GPUJQ6CGZ5+]Q@)2JV5]5U^4(f=#?Y-\XL;_g8K&J>RgL^;#
P4R:200_PPC,P6H9?aLEYB0@Y5E:60A)A90NSVDTXQ0J1X\a=N01^bVQ\/;9KOYM
U;c&S4<>G^WTFN>FP7N8+aB8=1C_d?(9f(Q5<OaBZPYQ(9&W5IYWUOQ:B(_,\9a1
2741H-C5G;[SUT=d7V:HW[5(M/c^(21dD#S,&JA^aK45gIAFG[X-FJ\fY1T&6SXd
Q6aGL\>D2O=SOWf/&e;NQaWZG927eX;5@R.R=aOf>/JDb=bd;[=-U]Kc&7#4Ra8_
.SJEO&(DeIK2_BZHC,4266?A^;,)e+&[.db>(K.3M(\494@b<OZWIcc5UMb6?;O5
DXWTJ5(]ZOaDF,K^RF6OJQ_EL?F;R8=2-W80)4De4c7PP/OGCYCQ-P2NV:FQ6JY;
JO?V\OAf9[A^KI,B^BVf[R0);8;O2_E\O0CAGf2&[T)V7dWJ8O1a4OP0=2>E,d?K
5eD5-O=4HFcW#)g4@#RB-N979M)]L(5ZERZNP-DYPf2>57;HIMKdCPWW;=1.2(H-
)9^#a31IV:7:4KdAc\BYXOO^gI4JJB\]FPW.G]B_3^Cb]9-;K&NMDH_915a84bM.
C5]LX/IH<NIKV/\C-)#eM?J?(U.Lg42+J9eU,AWZg+A=:&603ISf>Z:6V5Y@_,Fa
J[,E\-+03\G1E?>#<Y=6gMRf)(V+AK>GF-@>\I0F#PZaO42EFS:<ZFY-R<OI;-+Z
F])1J;S/L7/&)LQ;/M+ZLS#(9IE0@QQCH7WcF^0U2R5<aW9D1;1Y)YF/WI:bU::U
ZG)VEGfIF=_e]N>]#W]Z:.HHg=YZ+Q,gGW.dF6G),7:99gV>>/:7+<7RGf7fKTJ/
?[:5FV[YLY)Q4Y=a.X97ZB05Xg5.N,64<cda5^-eMM)XB#E##H[BPZC:)M(eL5(]
2@+K?-eQ35#>3b-J6g3M=N,Z>LNN,]SPPFKA78Z4KJ[F47I#XOcM\TAf7GU#6D^B
SR2F21.(,^M((L):/8(-JW^BW3P2Ha/DCg>,VV\4;?8_NJa\KPcLMAN0/MHHD8K#
&RWbD3WK/:?^@3O+0Y^MTFQbf5eT9[ATSa+>#SVL>/9Sc;=M6NI89Y3,CM9K(HIY
6ZBUL;B]1Pa=/1TN)\BQ)(a:DGA.\eM7W@PH#@5cGX7e1VM=-YKZ0:I5SU==0]B)
G[CWDS#gWWJILXD4W;J;R#4[fD]N9g=I?R#1b2GGAR+5_<J:Q7adf6W],HX>W@FW
_DO+Z[WQ]2Ae=,JFJY?@a6TdL)L&FdQ#,A+W\Q9I5)aKdJ6R//(#J&P_FTWAZS5/
U3F5<_U\W.b)Pd=E&J\Ac<7ELDELQ.PZBVRDN(JD\e7(JL#V@KZ+UFI,TKXOB.3E
:c7AECe,aF)KLFE\UVAH:[a_<T0Ib2V@dK>.RE@RUG8VDO32Y7R-2IcDfeeM+3f4
DFVS4Sd[D4V\N-O)5=E.aY-?HfT/UfeR\5aR0Q<\09^U>(CG+[5CDSd6J=)=S?D]
DVVQE:.GEZHg/\S>c+]AgZL]Td,[&+:SB;\?aeb/NOLg2=0aNSRU.@c6CCAMJ^U;
BZYIYN@3?/GI-,J@=Q)_=f/@b/;VD&M8-#KOX?=4CDAT&>a)cN.+K]A5gK1P8FG_
CgdYTSIG[-+XXI_^9/0[HC/9-gC>JZQCFPCVL.^)]A/1CgO,C_I=1]c_1P1G&57L
NZ)ZC0UV=.-L5ReeR+>.AZWRDe:cf]cC-S62<4?60O#@eU(.cG25=Z6dPH79Mb7]
<4),@NB14fb+g-E4(T.#@<OIAGdIYHK29QWD#X^)PPXGbKV2VfX.Y&V^Dd1g6=L0
1dcVA7\D1?9?:[QMfZI>bF>H?1Y7-[-757_EMNN&.KW<IX4DHTXe</fO7:D2AVc]
YdD<A(^I].&ae0RY-2>EdKGGgN:IA?JV[e57V.Mf#gCB1_3:J)Cg@+G55^J=bS/E
L9?XIJA^[[Q&]L#(N1Y5A;9,:N(TIZ-W+C383N1c6HB2<HeUgG2fLM[RbN@[W)?>
#(DO8BWDW2(08D?U):@9GgAMLQC/X\P9Vf).1Jg>#8/09BI)U?]7,C3Nc9.HHX)&
>F37R)e>/Q2[Od2H=.?4KH6FN@TKK>G2(_96bB,#3cH5>+8->Oc1ERU4.B7]]TCN
M^B2M4)#N:]bNBTW^-4;=c;@U39\.FIL1<>g9gEF2e8=+X1U07;Zd@:LD+SFV54P
X_\f-=ME(@1IJ-2[c4^bg:0452[&\O&4;_]&0E<Q)d4?IL;5O#VcD7_\P431#S_V
YE3DG]\_RYDS+ECb7IK07DbETUb0FFX)XC@^5^KYFdMeV)(99D/E>,H+D#R=BN.Q
6SCQSW@(4K11G6LK&A?.OF6FB.6KaI@5/)/7b[EY94Rg^8OEM>4b?^ZIC#J;07?8
PJW_Y<aQV?OV]((e>XNE&d;2R0A+?]PSfc=A#FXZf5<?0PF(1c.1W&69+AER369d
WeB<P-U:eA)a,N>fUBZ/6\H6U:##\T]A7E(&[9;_QBR?J0[CV-fd&5E>M5Q]T=cO
GD:C&-)S:\DPBACXVN3+A8cdLa[VfOIA>,H/ZgJTe[8-QM,+de#2f@6N>D2&[PaX
(32C]5,RbN0^N;/H(S]53H1^LbV#(?Qc;=#6IY+Yc,/EY3a<_L,@KTb?M6PWR.9_
0T9Uc52B]=N<<G1-YL4P;7,?BaZDERO.N?@SLOKE(N#W;K::23-+PI&\c_g=7.3d
?Ra0a(7bH[XBGU?\:@102,C5gcL=IDf?5S[BcNZ)DJaGJZ;+&V:N0&4EE2aE-,QT
7gTV?N;<LFJA#/N](QB0R>28BXRHZXN[12JESc^P1+C+,8EQQb9R\RQ.1<e-XE4F
XcF.N1NS1Q1[97;<dC0P)IJ01WCM>2JP7K8Q4:\6O8Ob94O&E8?G6[;R>9Z^>>fT
S=/OAR>FFDKVPS_DdKI;18NK6Q</PXFLGV9CS7g.BVSXP5b;52=.\Ad10;(TJ:_=
e:c0(?/V.ANV2^,I29[.-WMd?eG1N:;>eIaI>e&US[:7A?e0#PN:EI6K\KD:OReD
4K(9-YV<[+JNRY@F4N#^.@7V^N0Ya.S\PS0N1O_O9cVO(Tg\0[GRc84?b?bN3K/I
J>JL.9KD_D;N0(W>69&EB;=6X##.;OB39RD@:F>bddB^[Fc9&g#[dZGea^Z(?a5A
M=2e2#4Z1L8WYLMKMI3;>?Z<Nc0cP4>4ZY6e_:QQ4M=IU2?&[.eNJ6)NEC=^YOJM
3G=5;L><WE]G1fZ,ZT;7O]\[;?@;^,:CRB;D3^PLL@>LQ;+^@19fS1+GA[<QDUIJ
K4&[fKX]Jee0dXfI<H>\c:OHNXc=2bPX+3_V(O3&\[?9_)^bZfR(1b@\64H)3>YU
[8M[=XgZd\F0A@5H+(YN-DZ9;IO2^OfC=(d(aG;4+2Y3HOV,CY5aVQ?#1gON72B0
Wd1:2/Ae?.bQEPZQOe1I4A,(Zg_)8A/XK+Z0&00\I?L:XZWKJ+[V]c>5S:^#3EBL
aCD-UA4S666#Wc,dT_S0;+_Wd:eDe?1V9J-&;R1R=Y6[]\1L=M_6gNTV^EV^)E9b
MHI@YPWP_)CR>S2^fQL+YC#-8eTb1/-KKf&4C&a)^OEXD0aY)&J^JRCe>C=3NVOf
cY6=S86e<)Hc=6BRZ1\:O?RLHW+.>9&OY^Q_T1)\4ZQF/D1eUB6+>=(OcN(cfTN7
c.O3;-gE46U#4E&UY8M6-HfFK(:@UX\J@/7X>;6Z,1PNX)T(./3g/-P,K9/;/W-A
)0G>P1]egTPS/N1>V]Ygd@AQ6#Yd3SE9MYTB2[JPMM5UGW;fSF#HOZM[M/UNNV-9
;eDZ>G7YE(:4K]RM>WG5^ZD_B]BU8F1d[SK[]Ab>LFaA@:OJM=40VR-Ta2>>TT,/
dLfaXCeH4L7-L>d=D>H>J8&G^cPR=g=AN=WSbYeYLS1@cDG]ONcEgNHX.]P&8(&C
S[QG,O2]G@bg#K-0J2A)c.F-+^D1L^F1P1HYD@_-]9b4D0^_Z9W);K0fP]LEM;XV
LQ(ZLL&2Z\#._H4Ld38;E4CVR:W6Le1-8,UAF^:a:c=;cH<8M(g;7AeB4PQCLIgI
fgA4BGg;4\Nec&[H)4KIUJ^Nag?]J)C&(Ta9V(gSU&B<Be5880\;DVM[;dS,ccBR
=91Fe/e7^H4=<4TU<+Qg+YbW3GVCWC/CID(J2#g<GQ(2b;K&7]E321W[e6XDHL0N
TSa,&65dMcD8g-#EaIVY1+,ZIgIRV=2AeaV-0Q>]A:U34:]ceQHJU3fTBc\4-Y6g
B#c7\b4-I>+4a0Tb.T6,JR)SdLG,F&fFeP;,>V(2Ad3(;TA]GR[bX05[MGY?##gR
6TSAG5@X4WAAe>O3?fVZ(OHaHM/(4XcZ1FAD?HSe>(6LWO]Uc-fTWXC,;O(E:OV+
7B2.]MPZAc5=>[T4/7gC@54eE9++N265U))4S7F4>G8J[@LUM4]b0f[C,Rg/b;E+
[3f+5KI(^F#J.T(_(XD3TGDe3+Z^YFTJVR-c4URIGV<B#XLCSLC,fHECd4I3O6dO
4.A.E.ccbQR13P9JSg3TfFXMB\-M[4K(Z-XZ[,,2(RTd226R@/NTP?#3B7fZ+H]:
-XF\LH.LZG9[7/(;?B?cH;O_(5G0e;XgY;T+a>Ja)/2@XRbaEO-N\aD9_65CL[]G
DbP@[0d6L2G-1,JE.;#(/I&U.G^KgJB&_]LBaD[<GLP=>ZdED8?5@QDCb68WC4)\
.3Q0e5D/HJ9A7M_#.I4O07DA04NA=F\/;Cd.QG.MVK4-([#CLC\3NI<YXBK>HZ)2
^^KP2P6\6O)W/2I98H.-OR;I5RP_AH/WJdg.U;dU+a1NNa3b4H)5_K8GFQQH9W-G
U2YESYY1O33,G#eB;\aB(.cT9.USXSDG_Oa\Yf]4]GD@)87-1YR\-N/Nd?#ZP81E
Z&@>I3&7cI()0R]f:<-<J(3(bSP4ZcOb(N,()IZE32YTH5)13A@c0=fdOQYQ]8F^
#Q,D,:Kd&YF_eTdTOb6NBaY(=4AbAVBF\,CUA+K&7)&4;SRH0TJ[7V9I#0][(##9
8=dU,[@]P=U+H\/IOTBH>g&HI4+gR^,.AV@Q]HMQ^_V.L6&F^eK\<SOfV?PG>7c^
#d):?\G2K9ZKa]?TD]<CJRLF\1Ye]5HDG]G25(LJ[3,6DcWM=cGZ1#Q6_R)RUO@V
@6FUM@e4+E1UaHf3L^UOYCf-K?;f/7&MLNJRX551I-:9HT8bX4VdHFIF7RKDgA0F
\F0UWN+<a+=ZdY?3I(\G7?IB]aAcJgXH0.AV,^3+BgPIb1N4/]7a70SFJSWfBeMQ
&;GWH7_OC+#d&6K)B-5J?^@aJ@OP,J^P>?9g\SC>9gM,L0/RL2^LeG8+KO>N1DU1
J:KWFI4A)32O5E:JH]#KP<NcP9V,43a4f_BdKSHOE(Y9gDbPA;^[cF;Q9d[2ZOVM
]8bI:]g+\2Xbe6-FY4>1@RHW]ZTP.<Beg)3eM_S4<W/06A0NZ>\JKEFWTWb=b@;K
c5A7?]AU5K^>1O4(IX.1eAH:@^=0[D0MQfeUS;S0]_Y(R:&).D>;IZfN^:2G]g;D
Y,7E=EJN,Dc-,E<3#cNK_=U>H?TWGOMAVFWUb0G[,bW8&(8\6(<G/?SF5S/B9/4P
21a>]3a^MadBa2<Z<EB/&3eD9#J85IW[O9HL?OCG0KGAf@AADO<<7fHYE9cZcfCP
6QGVVUaO?S2^YM;>_YAE/CN\_?+3HKQRZ\W[C<W\)EX07cQ[GC;NQ&\5EC4eE?9-
B9R_5H3>,-_L?&>55C\[b&;@H:KS+\@40e3D-:9A[@5b@6=623AT5I((^X>0L]6(
bNF<J#eYWgW@eAOF<_g(GJ#]MZF1+MO+O=-9)B(:^QbS1ZW.=9-S[aC_Eeg6Z\L_
\WeSJSTVPZMH\\,]JMK#3=(VXW7).FLG^NcXZ?UYPOKZZ#FVg]E/</A28TgRX?5<
TO&a1<<+M=T/RK&JSKBR_CH&&[JI:<G0aRPfKQBER.aD]G:^Dc)_]I<H]0;\>^3N
?98/;::Q;3^,:Rc_A+K^3YNNBR0;>F4JJ1dMbUcLX>51PdMJeV@4A,e>aZK[3>8,
(?]^f8eP90d@U]KC;#Nb+HX#.de4^9ZSPD/W)7=FEZ:Q2?B1U=:[a5Q2O+VbHQ+A
C1G8C-d53@+8XOL/1GS1^J7;O=K]&#REM79]Z/,VHNNF92<=4ECa/W+Z<:gE:?2f
.FbDE^DA:f0C&Q9La8f7g3ZGcC>G>5-54\0ESA7ecdgU4?<5T_f2FF5]^S4P(&KM
Q&?-FU\E)A(gN]JBaOABN:b)(.-)B#1=KgdL6.(7>&XF>(e5b@;/,WL7]4T-a:#e
5@K<?QXR@P)KObF3+VBfJRTGg^_IUR:D(_fT9UMbQADT8^F@?Mb2&3HB?2KA3=fZ
IZP]:gD_C73/B2ALX[V0ZRNU@\V:>D>&Y52E41-5-@.JCA;D)YAG@AO)7^C:6OLK
E3=dU20gNFMECRS44=EeYX>,@I3;.^DY_a_7M?3Wg#(6,N7U2MN5>&W39fbVY\@b
]fJZ#ZZM\aWC.cB:g>.WO8DL73ce<ATI9Ya12?IW-HK/RN.17_15J#I,>>(GOZ@d
UD<6C]<50/F6X3+.IddafA9#d;-P<,J1[+cXd^SFCWeK]V&,ZT4#=M^cfV=Y_fKP
Q0X23#COfa0#[ZGSWQ+9,5]W]NS/N=TFWBHdF7Og9C#1D6J:O.1FHa0@W;gTUS9&
2OJeC6212&eg=KXGM4.PSb^2?C5R@D@BDEXJ4HK^FZgY:b-:eC,A/HU>7:2Z3?Sc
/4J(_2_M^>aUYK-Df(#X:27T)WG5K?cd\4TV.Eg6?KBG[Wg20Sa6W<^B,M_N2NNf
MS3QA&6C_G6BNLb8V-/JfWNaf?=H/WT3]L1;^I]B4aJUFB/=d]7,9&5P7UT?Pb/g
?,SCTGT_,6ZPAC5F2\1BB-82d&b:X:D>(HfXIQfM,@[0J/,_@RcSQ@?3\fAb=J6_
Xece@,V7fe^0\@a2W<+0cSDbQg=BK:;Fb;[M4g6J;+aTQTg/1N:/&d>2:RG7Z/S#
cUddM6HHZ5C_E^#-9bLSaWg/W1K4F3VE+GF1V5Z53Q<PB0ZgJ1I<KGKQBU7@g69e
WSK+)\9(deD1@E:&,T-+?>_KQeL[>DX-f</Q1:F1Y55(Kc;HOD/F:^Y-6G?[Z62W
UdC9LYT58I]0@-(;P@1HV7W;\D.ZJOaY/[-9/A&CEK3eW-G1N6?8@K<#D1aEMRbK
LWO@0APK,EVN_&b&M3f0M^._KdW3R/f<_H-K1F>Kb?6[3JO]OWR\LXdZCV2DP-CC
gH<A7HeVZUC)3>KY;N.-KNF(ZC/#VUFd.7+EV:O(2I_fb=+e>R_N7Z6_C,_10a=M
^<1K<6ZR0^Y=R&.6(8_MSg3:#5;&8XMD\PdcDK(:99EJ@CEO+,]1N7E>51SDV8[J
eJ[HGI&.PR)\IY,e\Cc.12ER5QbY=f.HY#>_[)f=G\7UW(JYH4+ZENZZ4FgfB_ZL
F(7<^B/Z4,&SA3@,OEe>)+a0DN)D+Kg-M4MS.B&>De1/L1[P7W\,JE,[W>6<6^,?
>.6/VE9I]7<6]==+#^M(&IbEX[7./a5P6OD8,eSWJUE.PO_;O58<3138H_+T]I6&
UE8NU4>(=/51^G[;N^:&JO&_.H#c]a6?790=K[<04A[e3K_0YgTCP((JG#T]-d2T
R9/cA0;<I_QAfcJ-FTE0dVXR[1f6>5&:;]IFa(Zc^8a5:L>@\](;SQ?N[LYPB_I)
VHUJG9N_RMCH\HNeFQRG0@Y-gHR-6XC=4Q#Z;X3Ye\GIHXF[cX/D+W?W]P5?O@SS
+1JDZDfcK;gAUF^<L=QX3>AJE[AU5P;YTJbHP]>(IV:?J6fYVL.R0JW^Pg<ORPb3
@148-QHQ.V&IU.-Ie>5I05GE-)d7fNJ02>gY.T?=gJLg@=g@:4]eG2A#)\-fS+/(
#P88C:JDR.MF\FEJ&I)MT^LU]XVG]91.V&C^FIRNO5E]Ia]NU1A[TO]:]Eg>/9]g
TF[gP>65UT(?^HCWf8Vd72aL/4[.ga\G20/HX#f/,J@L6eC(fC(b)I?8[L9JCYZU
5dWMTd<Rdf/,:2Sc5FM__H98)U0e,Cbd8U/OKVD/#B89P-gVFg><F07R8=T4BT4J
N5\g:.WIA]:K;?GJO2c8,B?2C1)M]:M999A=;GQG/WMd</THJI]e#)b#CTH1^TeP
fE@9=Rf#V4S^?02H?F>c.Qg70W_.@7+Z)+AYC4f^E6Ee^<Of5:Y-)G09GfeUBeXW
[W4#_V\4bNK3#P+>UIY;?a.OXMb:-PYCP>-f>LPDeF1R?F/TMCTNB#N+.g##<I]4
[=F?AdR08c,26Qe3B_HT4\0WLM<ED.2[\V&Re(K9eB;?OEM-#E/4cH8gBOPA[\6<
-^S)&gV#HXP\;fL17_-:HTfC>4B-WA#\OD/3ND:(V6XX0C0;@Vd?];6P=Z#3BBG,
eEaX#[NHI)I.[D(.>G4aaBKdS7.#X#P>+=O/H26#E<:&.=598eaa4R;FFBTI\:8S
;cS0CL);Y@);[R\cdS];9L/W-Wb5I#<Ng:EIN<Q:F\H,=eARUS2/))b;>#J1E,MQ
40eM68dfZOQ<)^&X?XL9O&09QY6FN>)d.0\EWM(E[&0;<A(9I(Y?RYAF:ITJ=&a\
^6R9\MQ3<Y;B7VD9^KA_e3ATC@d(A>P:4EI-I^)BG96HX-MD@W6Y3bfd.d+?f@5B
bS83#[T>T1ZH?]Rb]_6U5A&gT5f<IUUG9ZN45XJ+G8A1WO_+XC8TE6cK2?/A_0Oc
#4L=-+00e>H7S;X[LOQW/5-M]<T)F>_[=HOL-@]IMbVafg[Df+/&4LIgA&Xe?;\<
:TEc+5Z(H>d2XWc)g7(++0_a9,FZXTM&]ECT7]g4[2=AA;-:HH3(K7KaNd/&@(MR
R:T+D,3S<5(9Q\U5-2LL_SFV8/P6I#))0&<X3LdW\6>X#->0=@1X2A(MLXWFBMR)
21WHOa4>5GL7+>,dD_ZB\O51QLK\=0Y;3Iga(<BC:&D:=0R?700^A5E:E\/4)Q[U
)@,@9;HVCEJUJG<\_:B?:A#b:QJKC=T,T9XM/-Z2MY,6,2d+\Y1-eW,X-2aZXUb)
EeP_Te8RAT/HBZ6&R?TV_f/fcCFP#Ze[:5U2=LgJ6435]#<0cH2K6VHF;IgJc,AS
->F^I-410Q,Z]LM(F^:DN1P2=R)/Q-KTTMCJN=I)N[RWPE_+(adKJ,8/_4U4=_HR
fLQ0(S3,B-J.6@WCNe00O6d3IfMgZ[f,g)VW[d5>3BMR[QUfL)@))6Q>3g7bJWXb
\TNAM5g&X^?3>Wd-XdJcUda-=Y;f)6_5A&?S]c)MP3Dg9\324\9e:@A?PG3a//Q-
8K#/S9)?,.]32_@cX,L84L8.FH,+J32\RHYNGc2cO\ZZ1E&::fE1Fff(c2Q[M?a]
Z>Q7013B51GDbPG;P@CQSOZ16H.1+DQPAE;A;a.)aCd)>.S>[3cYI:fcCE&YV#+-
X1MIFd.\2VTC_\fRO:N1H3(]/H,4I]Z4B/P[[2EIUK@bP/,d_01FH(/?&KCBI_(.
&X8OGeb\ScPP&0E0UJ:LKO?K2YTM/X&dE>\_Z9b#53D/O.G7V214I>b@P6T;2_:V
:eYR\C_D=SNWNOd0:Q4\Y5_?Uc+FOR)>4-46;fB:U86VD0=;D8NNa65;b0=:[D7>
_CQHNT2;R-D:8JVL4J<U.fR)?E?)<A9K/@2CFUQc)XF2I,;K<eZ/5]:3R<:c/AOP
-d>,^_91BC0G;Y-6SWddbK,C<X2>/^0G2=?H2WF7+f_U.,RL[:-[=f&.bc0RL4(0
b,3O,T;:G8:K=-Y>1(72[_cd\5(3:IUdO;g(3IQd:be-WD\\K--&F<0CPWAXMeEG
[T,L9WAf4/P_:;S/,_3b\@P9^/]3\LZ]JP;I?CL1CRfD_cEHKTQgg_^O</JSa)9T
e_KF5XGaKT6YTLBd8-CD5a@M>[Z4__ODQ:F#7e_R>)O,[7IUX&4+Ub/a8C@Na.8Q
(NA<&e:e\4B4\ZKT]RW3J<8eMP8@g<&J:8AW(N.0P@>DcTW_=U>1GWe;0[3[\TeN
YBY5:d#S/F_bSd.f_5U7=Q.F&cS(JN/-L<?QD,X(K[7CQ3PL)K:aa)PP46QaC65c
0&O1?#MBI#J7^c)5K^^K84MC[g6dZY:2_TU?-RB4)?>F]+^Y28)@RF@-E?/BDd<e
f1HNB3QNXbMbYeHMO]VJYX\aZAag<GT^F<RAM7J9B]/O77AWNB5cSQB\4?VE3JQ?
;J5B^ae+LFMI5_<DBL/RUYUV^5;:V5)K1L.]LbIWHAK<Jd:(#B?2a23VE2261O6E
GY^F[J+N9BKNAcI0SdIPSgOO5^^T7eN3NFYHN,=+0UXG:U/5:dN#\LO&_5VbI5N.
f#@/X?Z&UIOVD0C-.BK4dMHUQOdQ7F^UP6\&[ag6.]L^JJbO7;ZYV@HQYaHG1_Y^
QT^3[7Z;U/J2D^Fe[,\?+BKE@P#VG2H#a9\KLSQ^RN/IdG3/6LGUI8XfJF.2X,?G
D1eEP#Nf:(d6ZGJ#Y3]aAfCFL;+-Eg4)de+/U=J09_R+T.geIE7AM:M01a:bSFEb
d(d?eg?UQ^(NO7+TfA0617EbUM506=D3TAG]g7-]J.aXJgHa+T43D>c,@>]OOS+F
ICagW&I9d/>4)N^T+^NY;Y?GcXUYg=\&-VOYBD>TH@(#,_1BYEDef[c(:_-Ya-=<
5^^E=1/4Ja@6K)K.d)U+G.><@AKXWZ,/eW;T+UVe]Ga4C+7B.>OC(Q\164?,AU\2
Ib:4\\f9V>]QZFQePJ6\9dE],[AF9@.AF^N?:1N6B_dN^3DSHHZL[(Z,I0[G6/#(
db^4d6NNA9f6RW40<:Z_015_OGD??,_+FZ@(c<ee]N#)D?d&@aB?R&8O.D:;JE+<
7c6JM.d6fHTHL.[LX,KT7SDbW-MS[;fR/dbS3d@L#9PZ,H1.6b.I;,#fd+_&?NVG
B@JcD3A&aE6>>8e<d9>)c@7K7MO_bQ7@LO+e9QMKdg;&-6P)WEVN?+^0<L)_JO?[
2NS2BBfJ1U&1SD6C.f8DTK<Le.DNJ5]CA\aPB^dF;3X7#.JfM/358aEUSYFA8J68
:9.P#8NE&cZ=A+1S.BVaM]-f07d_](3G>F;b;S=1:QCO7(CU2[4L6IHFf#R;(2F=
3a@7A4EF2LW.V4\c,Ie31+:Q.<?6=UcIJ6\8?M>@7M)T9PcMEVb#c8fT#U,U,S@D
cS?TQg9+DdWf>N>U0R,Xe\Z0.XC,Bd>1Ae^7NBI>F^^b(U?K69BLL@(G@I&QANYJ
LLVa-F:E+4TH:()YAT1XM\FXEV+27E^g8/P/eMQ[\R^=QJ_(CYad>fZQ:N4#NKOU
#?CWV1/bEZC#QTd-Nga]A\T\a&dO1(Q2Y/b47Se60CB,\DBV7218cb]cg:_4Fd/E
Hb_EQ7d\3b7@0.(VT:P>Z:/#]ABNEOOeS-WNdbH]G8(5#U8652?b5&4RPAC6Q+;#
,>H._FRFgc=CY7I(@+f.<?T]A-[8g\BO9()4B4)<]VXLFQd^&+gSf0BeSbV7B1F0
8f?UG)Yaa4Vf&>eSRf8R@3cK903=45WRU@/#):9=aY7[4Y<8LX>V:VOgSdCGQ[QA
gRW8C[3AH;(UY\7M._K>RS?()\WcU]L\]AZLcBA+/REFXHBBTPTN)95O9+K]=dCI
COKAWe&>@I6]2EWFQPGe3F;9@\N&HT>EGMJU@7d>Q_G?HR;1Q;NJC1d]IU,BX9f-
<>A[8c(Mg^6T.F5S8RNfPQ4QA]W0I]b,[V3bRWa+RX[VLM2_f\)a94#S.=b-?[Q>
+/VefZGEZa-AbUL188Q573d)?]1M8LA@&R-G,8F_cbZ.>&K8Ec2b6],IG?0=2>dH
0?MWGIT\=#X?d5X+SA47,(0AM8I7C(2F_;4>&@G=+5>fWE&E@UP@;W0Ig^EfD&YF
QOO[:135NLT<gY]5&TSA0KL_AFA=d<D>g&edIA+[\N_NVK@5:Pf)(RWIJ[+MR86C
K9@S2>:CE)LM+A5J@/;;BT=TQOD(M\AgUK#?UE+4;]#J=7bOT;?4&E9N^/?[N?ZZ
Y2V-613Ce5@W;H^+aV8CVQ)&I\Q[KB4JB2g_GbY@OgMDaA][[-DQ@4e0(GE?3;_Y
F-1URP;5e_P7L;\.61e8:Jg<O&e5>WG&IB&9880)+fDYXLZ@K5;J>JT:a>X8-fa]
E:e^>H<^f[NJ0/N;>96CHc:^&7]4cZMLX-VBO/.f5W]UV<8-KV??+#Q-:&>c+Eb9
:>-3G_eK87\VaH>X8,F)IY+;TZ26N/7J)^;K_>S-.-N)gf1g5Ab56ADUc(ecc6#-
Ogef+^CY\fP1c&>I3@PG)E^S@E3587N=Z)O[SgMf#>@WXS<\cAe.f?W?0=,]ZOJ5
)<HMF,#Mg3eRbI6_b:X.Zg=NX-^FA3)(IDB9[]&-Z:PM?LE^RA_@8?^ZfNc-P#a@
_])].Eb(=#83GR^-X+0:C\O4?&9C)J_RBH?:e^0P]W.cZQZeI&b6_Og,7dM^JUVE
N(+V#VU1ZV8&:HO==TJ-[e.7MJVMLJN)+8[9]fa3>^50;B+BgXf))=Y72IML_DC:
/P/bT[-aC\Ic&Q/7S-K=7D71D[WA,/fCTG-4VGM1U)gH/3[/@V.](d#_CQBdKQ6-
XDH-&3Xf+H@dd+C)O1E^)WXFfG1P=3#Z^W^bLV3QS+LKb-AJQ[R]8+e,7b5?7ab\
#+QeD#[O^[IB.+g;5?1f;G;b_<4B[R)@dIBUg<K6HL-PFR/Sc,K>;_RFEU&\eO2b
Zc+EYfN[dEO+(AV4:g&&gD7b9[BHG&Z(B_#e1VVbX0UUe5#W>?#aOcS0#OU5)#NE
aNNX-^?IPIDY)B9#1\I5FO71=/CL03)M5#@dT&4F<^R4L/,Tc-WObLR]06QJbB5;
a:UH#?:IJ4W+0[P=4GPL(.)6<?D[UB-_YS&(F]_1:DN965)gfQ\dRC9HOCeZ80V-
NbQ1gH[)\]1-+QGdM#O&P,7_[(BDS.a3NMJZLT#>\@E80aF-C91)GCV_.X(fR>8:
a[>e&+<fIQVJT&L8?+@6F@([[TY?.ae0g2L=#(PJ.FeXFQ?]DXS,K&aQLMa7f_](
&?FdQ7@a2c5NLQ+6J1;)^?B6NO\[6O8Z+f^DU0>BVYcbLX[=ZH(:L(JPKOKb0BeN
?dIX/T=@_E5;&=,<)J3>=WeW+4)Ta.M^=3DE<LC&1VgVU-O00@aTgRMHT5@3\,NJ
:M0KD43dPMXZZ9XggcG/FHO<+99J#8?YWW7QK=7\/a(#c0dWB)<91M:=R4e>d\/Z
Hd3U9/0UC()c>@?3@bY+LCcJVPcDONe4(JJ=6.?ZgY+E.683EAFT/=A5WfUU8B&I
YS/<QM;05(I3,F)>ZO[(PCM^.C:9@5;5&^b<.d^]>[XSW1GAXCfI&6TX;/JR#^X+
7+@P-?&,bS1/-1d(eW#YagEg=_#XJ#)?P1[0>D04Z6F^+\9(K6OC)2A9FJ.=.3Lf
?8A7:3QCMb;QXKVbX/VENB9#dD]FE52gO/E#])V=3gg;@WQB&6F/0\[@.)H\XWKf
SCVSNPF^]@MGTP(Y-.+[;a.V/:,)152D^M8-V9_gO_aSVF:eVYb839DH0C)-&e92
\KKG&WYIeERe#IHFg#NE\V>\3-[ZKGLS.-MX<ee:-=J9UU&V\TcK#SRF4)ED;Qf6
2+>B=2KQ(0C14Q\1^&#fa(7>:F=FTWIMeZ>:1>@ab)X;D&R=NK4[/+[BJM=.V8/)
e9B=Mb767AMO]/I=KL6?bCU90OeeG,\VJHFF)2&WTC;LM:QYQL^)#)_K7f7(>XHJ
a_e[DCbGU:(UCd(_JZg>>\HJ=49VIc7QT6N[bWXE.HO<UUNcY2fJ79A,1Uc4g,aL
&VZLN8YO;TbP9\M[YC()TfJ9&;-Y1[EFOdF\FZF/2RSaAD8M6?MN2Xf^=29XCWbU
:Z177Nb#DF(cC-&aB+,RFAQ4J&Z1@b8OP3-&F2&>OY)U)O=<Gd_f-YCGY:Ac(Q,1
M;HH5O(60I+&#ZZL/6X:,7DU.0DZ]CJ9I]P<9Be&4C,&R?&2cc^5:3QD2B@-/<&_
E6N9J;C/)0O@/)/I:6b7I)T=1P]4U[8HM0aM/CUJ5c=6N2:,Z/CJa]75OFPA\[99
bAC+/1XV,Wd<Z,bFV19a<[#gO;2Tb&9Q)8XE3XI1\BG(LD.ff6-U1b/=8,H<4X.=
fHKaKP2&TQ#1]&RQ4TA1de6[BK(U>+T1Z#?H/IS\Z0c>fN?G-9KY/>#\O/7.cCV[
VD=_\^V)TTXFgV]0PI^2DfHc++G9U_DObb+dAVdK>ZN=.D?:eXIKc4)N5Ka;5eJ@
[e1]<ZBe0dRMEB@L(53=S0>a5/L=22)ab]&01<fY&G(\=&6PN3E0#B?I;eN&&,BO
-JC2][2MWKBWOH(bCKbJeb/4Kd&A2,7-(;T8]gY-f..E.5.L.2HO9a/7cE\2DP8E
0FVIW>CSQ3&GCf^G_+/O_7:fbPU>H3T=H\5f@Re_\a#1gIFe1,e-N[_@P]69cN82
U/eVQCMO=?c\:B]A/O4UIgN0ZeSI;,3J2FFHZ[NdEfCEO<EL:P]f/2M1H[C37c#=
]+MF9F\5MW.=G_)_6#]d&+UQNY#/3XHg,dfJ/8;,,gD7IVJP#<YXBBB0c[_D>GA[
@1bBcD4=]ZbUU](ULC)KT@0DUe;?4LM1c5&V<)0e_C@YX)THPL?ZK5+gfHY-YdW=
,89:PN+M3H),0(J7aSXUdL,2^[M@->Q(:RYDI/:XX\5QKS^LIc>R=eB[2Q7#_RBK
6])E<Aa7KgXS1P0/O2S)Fa\(?QON=A.?e+L&:GX^#B5)RK=83SE/;]N7NM0WRf>c
f(G(,eOAWW)&CPD5ERM\;/KAS^/;X@]9H+()9=6+<OC8=-<0[+/:CP=NI19PV+[N
7ID->#Vf?)\M6R4.ORB+&ZHI\c#0Wfg6;IVJe[c<A:KCgAKIcC0]=B+GUL1:R]90
0N9(Aed1CZ#I(V+N8XYEU;Y8BL,FOXK(YFQ>:A@C^&/R#X;N_;Z.8HaH?YJ,@C;d
U?J@OT?ARY#62aRM1-,4OO3[&LL:96=7N,MKR0V)(N4eT^)d7R@C_gFV)PR:W5I2
S\=9W\(^);+2@XUUH(O(/OP>fKU(b.EJ)H)D:\A@GO5/Z_LgX^YP4@J#=Ga\cL>U
1g<f]ESJXJ6+9.2M\<I\G+eYAD?\cHVHIGD&E:aIUO#HSc8Z0X(@HDM(_;@=76e^
7aBGCec_Xf+6CZaK-PK4-P#?1QVNEf@HUCQ=GLWBa&+#3Z@YK#<D=;4B.2&-fWg(
DZ.-3@;K5<38GHRHJ^W10JENDM,FXVTU[@[G1#Pb,7B#_9>D[T@@;>/PB-Y@HZeJ
fddb^bY+,]OL672VY58d=e8V>/>e_:YZMTY(6Ma_E1S#L&6G-Xg\[0WJ.X1DK7ad
PJ9HX\50=)6=YZ9A;J(HaZTc3c(FbD=CPFQSSDd2QX2?>O]dUbcBNZ_V?/I#=:D+
cN0c/(AG1g&PE^\<_-&=S\Gb9HTD2:^>8J0T4^d^\Cdd=NL@0O3e3N2-Q@QYO4B]
dU6GPd6d]7@e).5(<P>V,K&3WDPgFc[2/O+=M@6[^F5-S&GI,8UW]HC\.S_NSa2M
ZJ@\H:d,f#gdA=&DQHQ]e-B5_?@0eA/<(a[VgH>D\JKPW@9>&2#@gEIWc5_a1(Z&
CE^&eZ_K2LB@RX[E)([-H3BJ9^3&X@ff4H,.TB=E#gRDF(9Jg6[ca6:1aafD8YeX
7M/)/9RgeZdIO6_&?SK(A_;@QDb&5gf33?2aMF=?-YW>CbU0=KQ>?-YC6QNEO[)5
@\?PQ3Vf)Oca2@J]1Q[D@X.&fX/F@UXQ&B;3-@[@4JcSF7DX199TH0KcIb,=c[U<
)=E::I)\2f@aeDEHfF(7/M:?4^V5+G6.CE3T^IOf=e8XaE?=(L<MO8HbNOV0+T+K
&F#M(aXPd=4CbFU2<.[5MS/\U6;e>(F6I>&f2J541Ka)/1KS;e)NUO@F\XRMA=()
XR)+:J6=KPGeX#A:?I5DgdC[GSW<5B:ZHX/RaEgRT6D05[_D^BbQYZ+4ZG7KYV0B
9;:CZaITZTc39>8-fU.?#3/JC)F6+)9S@gQf+,]NT,L^bZ=PRT]F\a2W4IS#SW?;
3V30J(R-_@L])U@a6,78=a>cS<LaWbb8M#WW=WXdgQ9)VJMOcgY]UYKEf.,KU3bX
V)<C_5cPY#==(<SUg]59#2+@[5ACU6.6e220A?)/=XV#>#0d3F=]/b<I<R()D.0P
2Fgc?M=-.XS\350MO\g^gF4ZO[@UbTd,([(=<E51E_\Qf#]I^g7K6D.E,4f[Rc.+
KbEUO41&B6O[6GI=ca:CCFP/-;=<N1@Z^aSeS?)/@MGL4<\O1YLSL0S/Xf/b(3f]
ba&0V.VM0[c/YGUM/805O/8\OO8C1gP\?_]PQ;UdSA;OLF\8U0gf:#9,AB<=].AG
0GFN0S\e3MD>R)8PE>)GDWZ#VC]/(@2^(@ZB.c8cd^=?#YLaQOddc^+6)bG1GC-E
e6-KOHb4[,6DA[WE;=XS<X<UF^^5A0[,#9CR;4,g#SJ_1Qf-GA0(@0\=<&LaM,:1
67Zg^;c&NcPf)NGe?2+IA#Q2HLM5-O\#CaJ=8]Q&S?PW8PK:.3UbVWX1GbKSSW+,
?V90b;7Zd>H][d9S7.HW=4):g/g&V@?b&ULb#d9XSDOIKdIX/O92[aWMEQ:N&=AO
8KWP6f:9eb1<HSP)9[:cWS#_e52aS:T&[W9A18VZPN>F-_[+[-3f]HbD13A.;HZ:
-FMgZA[-F\VBBT6.(/WT<^E]I?eE).&2-0Ff+I@V4S4E+EXXPN>_(CL0OC;>GP>&
_2PF<ETC+PKSJ,K,9BBB\_\@SBR:23V<8)Gb]7GdHWVO5BRbFJ#-@7:OP(-EMHNc
V6\N((?U^UCF1a\I@U)2FMd&M4M]4=0-#45c3-OB9;/=TE3@Q<B#0XfH2e6E@X\/
XZb7S)L/2K#\6FKO\,CDD;5KU(5b_V\5&](FAN62,#0995DPU1&X05]^J-_G)8#Y
+6)T[4M_=H&P.HW,QD/Pe#]:[4NDO371^9e2dJ?+KA&45S-aG)LZK;_,DIaIIB<e
UV4b^Pa0@0D]L;5BY:fVMN^[^?_1GXFEYM#KI[J><#WF5H^HEA_;R9A,@IbcIN=J
>,WE1CD5,WINY,1dd-_M7#aX0O9_]9VG3;?-WXMQLNS0&g4cZFCE19)[c/MK;_0:
g.d\9X9=8I:6+R]\RNb5<5ZNL31\Ac21U4C;[TW(2EDU1e6D?PBg8B.99.@>\1QR
V/ccY#?=B]EY+OKERN1EMPKMJ2@ccXJVP,X4PA=TB5(5:27+cRN0@adD7>^W;7.J
?01;[?5f(<J&S:\Zd2)?c_2gS4,CXFIL>WL28#-(6__K&E9-RKJ95/a:/A0e1:a(
fHQHS,ZZ=)_)O=G5ZdV^.W]]/O@^?W3cYU7F,)A-M3R+2T6c9+_C(a3)3X,=5I;N
#)aUT;(0d]EL_FCbPU0QKEM=5DQ)cIK=g4?4<3YFQM#>bLb_S1M7XU6&gX_K(ge@
J#6D99K6eYSfMg_F:#/.NMK5Z.5G9(#AVa[OS@Bc)3&b5fTEc=[;J-5,1JI_(GLQ
##aI2&G1PUQ-/#J6PXf6(SBbgZ8A]Y(/AJDNJD7/-GAB]_dG2^\-XA0+Lg2\Tb&:
65O+<@Z9<8dF_a,M#b(I72J?LF(^cNAT3/1=&GZ:)&c;0&9?FJ>U_0GCP9]77Sf;
U?9NS&XZVLI,eMdE^\N]HF5NFTa,;eFOVW6>^YD5U2KPTSLW7)/UWY(PQNME=.9c
3.M]SG=:W[087@-TS@dI8LbRWX_MUf=TTZ6:KRcMZGH+B:,4X>MQAYCOL((I\ecO
U<)VMf[2&fGU,TG86])9=TW=TZOSf:&[EJ^>fSXJ7eT.+FDMM.5dRPEW2;QXQ>4H
LdU>K76Z:U]Z#/J1OfM\4NR^0+M/.P<&Z98<9;2FE10G;/)^M0X#L:DeH;,E,S1/
(eK;>7eK0f<KHTOWUNPL@2F7T8N?;-WRN4]&IY36=f-G<d.R&49IO5JeHIgL^A.9
[;UPMH4gc4f&Z8Q9T1DbH[6EE,VZB[X)fZO7>eT(26WZK,NPdDHKG_d-4=1?W[ee
:U3JP;96H5@,X2CWbJ928^^cL5:R93Sd.@F;A\ZC/fPY2_4ET8UJ5)\>WFQT&O/#
Xd(VXNN4Y1[Bed2)W]_a@&F3ZGI,]ZBJ60B<4FK;CSRbN\ZVIQ?cc&LT&JR:f6Q]
SX(^FO<V+\V.>9Q7DPPb]=_=NBR)6f8M,^[W(QK?H5_>:QX7B\((RZNC61\+S##N
:9BEHgG<A0W5[,@W4gcWN(>\EgeFG_^9WTR+#2RE&#;?15@JR/#UU,fGKZPX&:X:
;6[3-0GUTHK5#5:KAZSbaA2U2]92HXD9^M-^9^L34;Md>KeQGW9I;HY_Q1FL_3-M
B7g5>3B_YKaeE@D>5ZS;D@S/PcCCKDM;#8LGS65g7X^D7D&]+H]N7#O5d=<)G;_?
N2IB3L;NI\[;:H71,JA&U:(b_N>5AdfNQ+;<?F]+)N2<AO8gd^eQ-^DAKVVgDaY)
9;?#BMAeEaK>Q)f0KO?[(H4Y@]2AV7ZTM+\MCXe1Q4YUNJJ<c/g=-T9]@,6b=Y9I
0dH&8A_I^-D;KGGdH?WN5ZT/eLLEHS^WJA7Ud--cUN>a_>):V2JY8MS7RO^6:CDO
eWEUM>O@1?INX8#Z#(#QKH[5>IZD0BcPXEZ5,/I9g<<8CYBS>;f]JMFJ1(Vfb-Z<
J&4LFAeZa[f/L4Ub(?D@e/ESF&E>RQ&8BMbJ:3SHe7L?KQ_;5(aUN.NH?_C=ILKe
B47W;WCA=5Q_#6UBS?G._;I]7f2,P.-fV#4d+HXE=4eP5_GKge()UDY)JcXRNgdT
f8S>\Nd?aY=H/V?LCRe7[E-,&db^21EI\HJAK@J;c3Z5b-5+g-dZ&]eeS8T7ZQJ5
C_U?]/=/&0N4fF1&M[LHDIb7,e3d?ZJAIX_\3847fP>-Ff?Ed^eX^Qa4836(RCcB
E24.9UT8eOMWeDe;FeO<^KH=E/2d-D=/5:g<T3]Ye7[<)FV:?PcGE8f@Q/UDQF#G
/_TTEe>I)+4Q2>M8<P,c]3;QKZH8DWH0bfYC0/Y#9Q9(gbT/C-G/AQ)(+-HT4?3:
ID.]7\&7aIF4\Tab[FXB/&5HZQ#6\>8@?c^LeKV)LK@,@ZULMaf^gcfJVYW_3_fM
Kc[58>Q\M-BE\&6G,fbQ549d:.7A6fU0g83E21TPb?YTX30=?U)P<?a4B)>A[S>0
8D.GN?_DKaMSAVP@eO,Gb/FbXUS]F1B>c,Rf5Y?eZO:e,;V03a1a\H#DD4.4L\g/
MPQ8VV[0W[gdP,0ZUG?8B&F,D@WI(?:&bg+0(&S=(WcAQHQ<U?Z3QDf7BUNY<<ac
?U91QZ+3Qd>c1eE8)>[]aC].A-+PIM3R0A-dVMAB8FI8V2&cc?@.Se],1_&Q,La@
g;J^_S8?N]N=X6gN#930V1?Z@6;NG,4:&RT[0O<:PSdf^;/f_F(/J83CPYU<1T/N
6^Bg30aL6.#W=.1Hb91F0_9ZF1E6_W7N.XDP+F_1WTXLC1Xf.SA:,2>UHgH<f:6[
Lc\P7afDP&[&WTS[\&cHC@JgCE]5?@]:_VG^D71DAQS1CXP)OOY\RfB=O+MHVZAU
AXJK\]Q=#ZEZU-0PBND@,[.=52YD+DO4249D)4P->W3I3C6@22gCL-.3166eb03\
V\G((^<SLG8Tf150;OdS9b0ggVW4\Y&#0[/;&_>aGg.:L/b_:f[7ZQ7/N6GM#FAY
:+_2M29&H9=[ZJC2SFASF&\TJLMW;EZcc>TD/D_M>#Q=Og6FMN;7+1gYOM+NTa#U
B?ZFKe^VN<94J@)V1EBGE@]EVc\8MdDDZQR9F.^H?g-)?7P5Z1CGAKLV9O2W@HYY
FJ.Z3<H?\F>/TM&-4?2^GaO15]2129M/?:X8NW58);:g,IOa#?B-4BOMD+)6:,;a
^VcPb:^KB]W+7?Qeg)S>.L45DDadQ[GZKfY^cIZ2f+&K2\),)dJTRD44LG9BN]0H
?29Y.[L?:<c:>cdA3G_4JY8ZAHVCWaM4M#GJ.7^#Z6>Z0>e<0cLNL9CC=]fJMaHA
BTbE]:4Q@,S94W:Af\g#ZbA-V>Z>3.:BG^I\O2:YSG]X+/_X1dC)=_<;2a2/3=.P
8L>bGI+3M;UB),1cSKH]>[<JRQ-<_C42a>H)&?T+I2C-7SO,2,PLX6J_AbJ;a)[V
-)A+b:@#.IQ]e(aTUe-U](&L</9:eS@S@+6bY##+.<I,L:.bH(:\:dR(fLXII23M
8UTB[5&1^A+,C:P<97]Y;?+Acd:&8-eEAZU+AV[dfa^+/WV#@15+aX5U8,FA=d;B
XdE.&aU(C9S)]U/CE<?<EC;(^V^)W\322)aQYPJZ0;0-MJ:.NK7DUU>S((H(b=SP
)0S.a:L<+];Yd54@#eO7PcN&\>:P:P7Q1;U(C=E[KcB_bB4?>bdL5c0X8]3<FP+W
=S=G_8H;.T2f&4\\gG4;E;T+=X>Y+5T;+C1,WWKNMA6a.Xc;)B+c&c3:PMVd8[1:
N+Y5C85MTXYP9JQDQL;-PLIB6V/gAW?UbD&5UHa0G?/^.S?H&+T1Cc.]9fHR-;7I
GaGO^=(OX@PgI)^WL@_,F_f>EbJcF\dDO99OBR,Zaa+]9BO4GXNS\Ga16N8#ZFC9
D:&8._Ec>V-;(+G7TZ2GZNQEUe>JTI._KQCP.U8[.X](+b0\358<L8Z662>KQY&+
c7_D9T7b_a<.e?Q>XO7T#6:-:F>Ye3c>E?e+0)=9aA>K\R2D_ZK)OCPML58O,FD<
e5-7TEY^F_eI,0(8JU[#QK[YVQT,P\S(^DU4D3YMPbTbLHSX2D(d]/):O6C094NJ
=NWKcT,eKg,NP\BX((L;XGCf^Ec8A33^/1dR]C0@#aN_>29XaGOU_7gJZaV6I:19
f)5=1V&6cD-EgUVe/eQT5()_Z@9:g4N+J,H\cXG+U8GA=dY,\@1F;@DB]TS9,W#b
XRC)VJ=,MW#dL58VKJ)-Ab@HHYYYA[A-FKcNL^IYJ1KNQ9>DS;:<)#?MD[7^.g-Y
,Ke1JR.ee>fPM[D7Z.FM;<8SN\f)CUIN[\8687[7>+B:-KKX_E6#Q=.E5;eZKa?1
+\LF&^=FB+595_<Q#(<CVO4(C95aD&3ZRJLg>ZXM=(DP0\b]8R)=4=;M,BfK;f3N
R==CQ,NbbXg2bG2,H)CKTdSD5HT##ZVg4Be49[-d,f;35<c^8a<FBdAFE1N?L&3X
e>YM<ZONQ]LGRWa=E9@QROO<)>=ZGFfU#HV+U4W72+DGS57<OJEGc1#F+#[.UJ75
CdRZ83(@B?#Q[_KXA3KbFJC9e6+G-HeQaP:#E_UW-2H(+d_Y([/?cTgcJQcX.;FY
AZ@D(WOg,A:^S:TSGP#f0c,-H4<Y.]E9ga84_Va<I]C6OFL63)N^YIC?\9d8>Gc&
+(IeX),@S7/PQfP[(8MG7/.,AFDU)SE2JdZaA<R3f7)-Y?W9:VBU8VZf853#\-?-
J+=LAP#14?2X6YX&96U>]M+>SVX>&DFTM)151UYE>R,?1,79C]4IPYGNF3R/9_AY
18L3gH-6+J9R1UbMedKQX=G?/F/#DJKK+-:))C]28&4N32c1RYg)c;a-M.<P<M,6
.eZ;E\c.BB-[TeVI[IIg]a]T>d@H^DHZPL_M1EPG).3J@D=.RSeZCJLASJdL4@Mc
2T?]SB+<W#3(a<OJAK]MGX804C]>T7aO>9)[&AEE9&055Ege5J@#-UHFQc]/Pg?c
ZWKd>]Hc.TL9ZDcQ(=YX8f9)OJ1-:=/2Z25JGT79TKc7X6WEPS-_R97?fV0\Z0_H
D?fJNBHG8Q8([51]B:YW.U87d3PV0_=Qe>KMBJUIed2QWN9A&g2J5:+IfSfU.GSU
U^e,:B=?eP:#fAgeTBeS_BTKB,UA>26PYU4#C9P,_BCNYF4IFRKUOb:QTc0@Y?gE
W(_40RgH15/=,Cd?G;SFH0MS>G\eVE?BEM6@[G#=2KJVTV\4Z<C>?S0-:bbYUN=b
H+72.XR67Be.Y2@fR?2)7<(XKGRHU([EQ)37=WN,&).]QN4:T0+(c]DL)RF@_cV#
2J5Db;3XVd+D-;9TJXH4GL:1bW1Ugg+/8G2VQ8UVea>A9-0C=+UHRW9OPH#)?@FG
3Q0\M>-1Z1>T6,M?J(W)21IV;K5EQT?EC#)J7\LFTP<3R6LFaF1.d;I)X:9N;8D3
<.U>X\.PGLETWT\C;(B.]JM_.e0B8gA3;/cP0BH,3g0-5D2e3XD4?Z.SO_C5E_7[
NV9]BcYHHC8,0b/[:ZC@IJPDXX6<VEK(M+Vb;GS<W9WG^ca=IZ,YK0B/E;:?M5TS
fB1d/XF;[F^dC77FG_:@IZK?OKfg//@7M&8&ca.K#RV),J--;SQ;3GHA<H[^[cfb
QUV)22d/e3,>\0B.edPR5D5YFRO43Q15f^,VgMdJ:PaMV:b,T7F+U>JS9_S/1>;O
\K4OaZ^M0XK7,-M(RP,_P5_PS6YeW.F+KEWQKR+24_2JCY0a^-2cKSZBKZ\SaD+,
Ef[4?A5[RPYCL#JPE\LL4E3<N>235bFR)4BbN4S(S<fZS10+S-X7\0[H:.V=[:AD
(=X:V>]129QGF)B@E_Eg^AQ2cE/9WVKH+4X/DQ[,=YO&X:XF60&HPWC\;8b2JYH8
@1AcGZBO.PTLH>M/g)BW8d\bKZGG0Yd+&7)GV<B20KTK9SU^HRG\KXIBg,bVR08a
BU;Z;f_-Q&-W<]T>fNW2BaS0VSZeEb)#SC(>&IHfJMZS@8YU:7L=EZ_X1^0CS62b
a?M;VV;[S)^K2O,f5Y)M-7XQgETRS0^X+#S+DW=8JP<bWI:T5FN_+Q5(M0HAA(:?
<;ALecH:(aA&/Qb+;]@0#(1+aHCe<9I&>5dHI@\RR4RFgY:#O7bA:M1.2?[f#I;6
10WS2^:H.KM[4U>DeMK;T7[)RNQ#fdZEY+.[J2UI)::Q75YK>WBDD5H[K&760-/F
bM:;@KgRR96N[)M-I2+Y&3^V4HI(b.J?gC6]=0T4McQ-/M#cdGHSC8cI8NZX^,:6
G#gQ08,=.SK_BGS(Ig>A.E<E^U?g-c?<RV38&GEb;\\;4RMDYH4^N?c69KP5JM?f
S=>7+TTMTA[_^-^@S@,-\Pa1K#R+YCP]OIZ8G^GU<#1]bQ^Ad&@)6TK\D)CF17N+
I44#e2)#ZX86dQ^V/W)P?^AM3b#VF/&5G9O7]6I-;:>Ib>H=(#gX?&Ta+V1T_X-A
@3Uab<KB\I6cVJU]PfG=dM#FIU1Z9eQI;7L4,/;Y.;;P<@gP100J[NI^=(]S[bDa
=V]-JObYa.WPNFUU[acJK+;D4fd;QY>#gGI,<[OaE8O57:[0R_SU<(b>XE7^6.)-
:>8HG]8eS(I>(>(_61NP1Jgc-]N/EF;b4O@E5LWUaK0_H??N>L)X;\c]a(a;RJ/P
<<V4.WSgU+E<[5C_F5LJO[UFIM-6YHJ\MIB^4dX_)e=PDaf-@1+GJ,EG-d+?R79b
(FI;<>U6>#bWE+T\N6:BaZ#_+8CA8ZWAJWG3Z9M[6;8&WGX;GBYJ)LafG-ab9AZ-
XLMQ>?gR]1H#4f,5Taa)cVa1ccc&bg@RC@>1L+RW8g,VRIg5O]>XP+Z/USC4Ve&O
\U<E(O<^F]HNMIC>.@6B>F:F9\JA[b^7I#@(Qd0a?A\=<5^KMc9B-DZYKED.TGK=
e?TT&LMGQ:0=J4:H7Z;L9.;ATL2I+CS^Q1H(_C^g.E8Md)L1fd9BG=&A^,E@XX(@
?4C;@VA;FA+^?_@-dE_4&F#g?2DIQO5X)4P2b8N4;^,N3gPNW3c^Xb[.B[5L<(\A
&JKbB63U41e?6/)VRQI&#Pc&PU\\+:+M+#J#=50<1eWW-XU55NI<2Jb&+>(/C#8b
S81]<I4@9TD&@/LRQ5g>-g_DLYN[@YWQ_8S43ddB1.36GW#NQVg8YXc,&6Nf,.6.
T3^-0DM_V9VP6-1ST198VaPF0>#J#K0dUGX:.\aNY5^dXU23f]T/,)gL@?H\KR(C
5+=CU=Fb>;(&V3\IH39Z@cBB#5eD.F]16fCO9Z+1W;\&.J_@?XVN/dDR:,44YBR(
g_4.PPT3KT55>SXgT;6b).R8J\RaWKQa,RZQ,a\Xed(H)2)eJGe4Z@AAKf43&8N4
CCXGMB<)O9,W@+W.PD-B1ZffCM\<>UObc[5_?D)V@M14aZ#E-B);eC7,d?).)A,b
HE2;SNZG_b@Nb=H2_2&VG,BM+<^6BUSIXJ[-5,+9;0RAB8\+YR^WDT67,5+75VGI
QX(5Ud&LD?/F-]4aBCB#-9HA.(T.\ffPH52EL^eKFTB;-33bXWW(82J,QW4>#4WK
:KPY[d)e_(JPMFU=6PDLJ]g.,J>+TA;6W4W4?S,E_QG;Y)BEXcLNGdL9B0Z6J-W0
XSTV6Zc@<U26,6[6g-ZD=7X+A<@R2H>;b;_<[6L6b2+eI1?c/:B@0)BdSXEHQWO@
I1\cEB<M.(SC=(U.gG7#D:efS>.=_deM8-)4bDFgY;#_6)KI]SM/)b:H2d0V6F)6
=NOeK-YNg+6?WMR.OU/;C9a<6]WD0W<BS9BN-WJGRIV1[YHEee95NSDRBD7^]R6H
C2Y^(]7YHQOQe@ZT&Jf^^WGT5#7cNE_d)XQUO7f:\f+DDTa^#Z2eSET&@_MQ0F4f
^.:dB4_\Bd2TeHKd/R@E,=O&+-U8O1:WNa4[XVg>4#1Q1O+9C00cJR>>EV8ePO;E
O+&=A53ZAJbBN=IMbHcXF082HM+Y-6ZA/]Mg&]]-BZHG]ZBBG2>QVLc<e777&@)N
W3QNKKWQ97B6O]Y#8AV2dKc46G7O_/LGKFT_H]7JR(^,CZ+/]_d-GHTPf[c[>RBf
8PPO6^=/ZC4L/D3.N,Y=E]M,+FdQ^#DcGb/c2>J7@fJOZSPWN+XW)_cd,IbgcH5A
<<edCMTUCR,FX5/^D3,\LTb(<7W2.UN-[[\7GX4[?4X[(fI6M@gfQGcD_Ob-bQ=2
FfS7X7W:gg1K8880BXfAZGgOBW5#8-g#9JWV4#,1XGbC8^35(eILYCHN-K8IQR#&
>&ZDaTV)B?c\ge=g>gb;(<dA/,/&TJc7&C6g]eFE64ed>\gffA&WK?YWV:\<SV,W
?_A+-/7#ON=8g.MC=\).TXb;X8D^_)C59HQ[CI7c[P1FI(YAU>:FP>I88L(R\@62
(RPNEY7#2A)JIK\H\Y+]#K94cA+KR\8)S;HT,:BZ7IWMJ,.E-M+/+5e6P1b:64YR
\NeH&ZZB.O#Y)H@_5fC:E>@;\[?g>+[>M=B/a71Q5@c#];0<<_)-S9S>^DB^XT@?
C8Z&D2a1LT.g9?-[UQZ,-@@\DV/3PT8eR22aV]<G?Ba,_LVZa2VN+\R.>K^UHAT9
^Ca=IfJ&PH7fGf=fAU1=UF?N8K6MI;]G7YQ/X/-8<98f^bN8@^UDe+8T=J)K:d4\
-#8?(bF[IcV]DW;Id+[]Wc&,.WZDH]HJ1M:2^DTAPJfX__@BC1OVg-^C2=]1/Y[F
J=3Je9PJ#>(R0K-PMe#,_WYON8;cJVUY@[&Q(S>D691DXDcNaJKRHW6=CI[[)P3V
,,@Zd]:(>\DC]GB;0?>S#^R4fL/N(_a_QeLP,(P\.;=:SZ]O.FQ,<Tc^fZHM3:LG
)AF6WQKA&QQ1g.)^]5Mb2\fQ>M9d4A-S-e_dLM[<(V8.G@.FD[Q8R0cEAGcR[?U[
U:G8F5d4JM4Z[EXRG5dEEZ2BY@Y4@+H27O[UZYOTcW#HGP/EN-6f:DC>b+FMBGK2
B:HB=#C(ZFC))g=>:1eM1LBa6X^(_@BH#g(/5,/._CDfGM((3Zb4-.^A(;bEYd^Z
G&#S(=M?IQ/-DLAQO,ZME#CKaFSQ--K\KI@F(^R-eW1e0/H9DLXMKg=WOI^3(FHU
\BO:N8eYV=II7(N@.f;_#e=gHB1.eZbORA#-G)c&7CZYfVYA.&4<f4F+?HbZaeK;
b2gRO+DJ8@#5TYL(8DF;>5]]6CXKgF+R]-^P15VHXdJf6g+N7&B(eeP2?]U;CDX)
1.Ng/BcD/DVS.XEV.ZU>N)LLR->\.]4YYM[@O3a;S)^YW#a2D\R&X<Jd@e:?2eLA
Mb,4;ffbVXNM2;:Qg:eKK>:DES3X(b[HX\Y#_;fb5XW+USF/H:O6KeXW_;A2\9=1
dg19EQ]736=<(Q@;]R[WEBMWV[dGS&(g;F@7#)c360048ac3#FMCc_DVc/Z]2]BT
-DQ4a?].3W23(b.[LI>Db?FD7<#:A:[,5QA5Kg-K/W#C:=0<_292?CD\^GMZBgOU
6]5_8,9EfC;DfITH@3K<bU/I&J5eT][\WMe=MWS4G,K2V#BPZ[;OJ<e5C;K:V=_<
[;RU9G<O=.7>5&3?:E@Y[<Fc]HLTA>:3&VQMW&@#9,K-27Ra.[-3YcCQfc#<FMBG
IKH@6_1O)\5D_dIM@[-(W(X)5fU18e6X:_@=L\?D>Kge/g7SZWS+RgT^S:[@eHRC
@)g/H_\AQ,NKE@0?aI&JM09d;#Y+]PXU7:J_73G3>@A+#04J+GgN8(@B.F+@a4P^
.\KFX5efQD,C2c5Zc6>:TB@&eBa/7UC0X+W3&KJ<86ZL<GE=7]_CIc_4Z7a;[#fc
dOM)U-J;Db64.&,25+OC(U(^9MD^Ded,&QBVO>I?0)WaP,WC\LQdLRQeOg-WC;Tg
[RD0K-B32#@@4;CCWQL,gTKN;:]La,0=M(SF6@,0Q]T#cZW2>>S&>]a]ZObF6d>[
+:SM+cd11^Q6MfJA3^?g8ddDZdU8OV?/=OK)P6F/ef+TbC5?Y3b;M,Qd.9Kd[LP<
/0RD+QIXeAPH\fFKg2GUN4]+#=I[&0Tf,;K_H:LPDPg<1AC>CL,+S28KHR3]PFLO
[>((=(5-3QO8c:f/<0Nd<B145Q7DD#gD@DMb#SP\,#]:V\g(-Y3=OO]?Z7>RD3c<
1I^J1KK9E7X(AQ67JGPILU4=-g=L=6N0dG:9LQ<g0F8FN6E6,D-^T[5J-1P+fI-Z
]:g&KZK9)N8]P_=MO(d1>VWE[PUWRZ@+A96fT.?ZK()=F>)P9=C2F7@d(gedI9:P
8X.Q6@=Ca]3QW]^a25_O2aa2B?f]c&Jd@XNK+5L@)BQ7]X+e&.V-6YDYX_Zfg17I
ZMg1N8L2C\P1dV/D2.&I8MFP51D[8e;a[DX8HRR6fWOKHR]8M).>ZGG6c3GEB#3c
MWIgXa9J\08ZHLZfJ7&UK5F6&RS08,LA(;,P(W4Oc0(QPD^J6F)=1P<QeJ5CJCD5
UDTR:G.;G35?@151f/JM>NM8[[;A-QW.MPR-c9JS=b^H[^d@0G2ZOa-<D8Jb2g77
8TZcbHH1P0T@b(O+5V__1_=2HDQe3JL=_;GK8[Z=7)Ve:+eHTT55^9e+D;ceB&Sf
&)DD[KX^.K@WfZCOZ-WUN#KBL81GeVVDYM+5fKa&+H^c^cK<[>:M;Hb1gbd=;PY-
^b:(eOB^ZIa+HOfR.\03B.MfYaZe8d1Wg,Q7Ve1Z,D@^SB?EV+<_D)W8I-6A)M#F
W.Y8,[23I9Ze0\PF_Q004;1KQ;+eJA5#IGJLVA-J5XddV6BI)_9LV2(5+1>5@\/N
<G&c5=,BK6fNKYPP5b9H3:B=FF1J3@g&;D/+V.HTXAQf(.)34eB9_X3c_HQ^_O07
Dg<XM<Rb?<>e;D:M^RX_S\3#QHK-FL3)_0aLg9:cU>-R_UCeI2U]f@gSAQ9=[O:]
MD^AGAc4T,4Ne@e^BJ)UOIOU5AL\C(H0Z<X^fWdW]eYCLY+KIPL-3f?C1IXAf.OV
W4gR@b<^[_/^_M](eT@/<J7H(L4c;I7FAgX_Z:O(UJ>+bJJX:8G(\63A8>.5KQ5N
DW5R_a8K[cZc^CX4?IfG5Y-\K:I)f)B3]4D[OKAFTPZA1Ac3L,Z3Y)(?]A3&\)<B
P5/79)S6>\ZQVV?75;OMg&<LFS7.:d>>6G@-+8[UZS\6[WRIKKY^5_L_OWN/&Xb,
^,5M.9QQf31f1M:I>:B3S3TO=K:Z\&eTd,9/0]#/fXK3#.)A1X(L16;\]B\-UJ7_
,aCM+06f3+NIBM:c](3,:)_3XC]>_g],KESbICNH,2OQ)LF&fL1/IO+_7XK&^?>c
9#KH4_9EAU2XHCZS55_82b<8&3U6]g\VSf8@6\JE0(T&VFgV.RK>L/VT8I)-@XCR
2P[[>cH8R?4(g1Le(8N2<WaOcJG,IS6#f^ESaV_@J^?(Le6f64)TJ62JA?-NG9?7
B5B[1]20LSDTDff<K7AUP&LdBLXcAO08A.,JBU>+#TdLOe=Kcf+g(O.HeVa:_-DG
:8M7TDS#K^:?NVF.>T1SUb/#^:\;]<S./HCQ+SS1)?TE22Bf+Af9E:T]A0bDD]+=
@=L>g<HH>?22VJ^:C?W(1KPI4G,PMg?dbI8/0IU[:,95R[8;Ld2CB8bT-2;6?FV8
H=d9O87=YY7&TL?XL7P&<XYHV?X&(O;9IK(_;L.(T@+0NR[Je:Q7JT2JX7Wf_Z3)
#961QXJ8Q4Ue,91SVS3Y72<(JJ>0L\S:MW]fAJWOOYTd3[O<HV(9,^K/J:8g\;LG
-_SCZU-5e/eM9>=NDf\b3KXVNfga+SI3YP@?476Q,M2/RS^O6V=)FUf7GBb.<E,D
Q)NU::.5)d:QOKP3Y<)9ZZ0L@(P<[0O@b0V(5Z-F:fL4A82H&baM#ge[QZ5X<3^/
J0/J/TOHIH&_5NNH0Y1D&H#Cf@HL80fBNA0W7?M73QbM?V:)-2UEKdC@D.9K0Da?
9RK7-AUC[CfD.cQICC.+-f,@7W1+eGL#0IH2>b6dM30=FH8B;B^FUIDZKe+J2@+a
-KT=A]7&[GaY]HM>WH7Q^-dR7f+d=ED_-,f-S=?eY=YBL;6c[PS26EX5L&AH)]4^
P&d]N^QV+C9.]6RAPWAgB(?8B8IdW:QaEX=N&_gM\BeK>#6?&&GC3Q-/GO1dL/>5
9>(>JIIP56KMR(V9=EIC/^_TbLMC7:eUX-]SdD_6;F34ZNGU5XB>F&S\PfG.XJ>>
V4c_c&29P516ac=M41)GH]T?-_UCXJOY/AUaM@-.MaZ2ER20O[e0#1SaVT_>)N11
+E..ZQV<e/<Q0OBe;47B;P.GWC5J[7CP[UR84GF2?S&)-3?CLYe\\RTfY=V0aI.G
W7O?6S(;EfbH\#G;;TA;G[/D6(^NJgPUVX7X>Z3^N3Uc+ED-WA<g(LBNCVgR.=1&
2CRQc-ZAV9,/@YA+RPCFeP4SR;3VUDLc:XHX>6V4MFZG,++6](FTBJ0+bX6CDb2c
MM1gV,(GBF;a8IN_D#^L,;=?+0]E6X59M1+f@_/ZS)FeHeS9YK,J(E/?@_NY#@;B
;_UV-?Uf0]f>,d<TEEC+M5\XN2R[]\A[WCHCCA/4fW1XgHEET+>9aD:8;:+C4R;Q
U#cg.7+=\>VS@?<3((R&CXDIX#)OJBUR\]+Z:cDdAB#F[@Q89#P7dP\g,X_BV;T1
.<MNPTdA(9VI1K.J\aIFETG6/O,/S,KG7XLcQ)>U3@KN?eBfL+KBY5F6^IdQY977
J9^U,VARGdbMY&<P(3I^,)eFa=R##JC2#5+Pa&VX7GcTY;2B/PJNLg4fC<fDB>fc
CEG/>ZN)QV2\\8)Z(c>?6c0T9Z7<cPHA;H5Q:DM8>-?2#YGPI\^\5WCc98Sd4IeH
#KI?W_=<cB#\1+GcA.dT^S=KO,(9OfdXCX5bK?&A@#,gg1K#Kd#/BgK[d@XRd):,
f(@Q9FbIDDZLD&[g.5@3I..XU:,+_e4?-9P-C-dJK0N2YJ2)#-0)[9C,0d34b\Wg
5d2HR[bgX)RWRD+?+J_YA;:48E?++XC<6-@5O3).]^Q+C_T2P5X)?WMEM3&IG\)_
DR:\6:TX1K[E?Wg?gOc-2eN8F2E6J6,P/aZA^WefCK0-:/V0/X6eaZ<ca;\ef962
b00TVa(5DKPY9W(fFXWT.?@Q&fDO+DAJL>Y#9>EY(F<V7@_7.6)#P]PI>Pd94ON2
/6c5KbZ9&7<<2FF/\Dg8UF:Q\[LJ(EZ@I+e5(-AP:,;@0.\<b1fJNA4HFg-15+Hg
AN#U?dJRgER])D(_c5ZQZ=N[c?U:X7&cR263;E1_A[(OXeH<JY/Q0E5F49F0_,O)
/KM]?-&93[JK[.G8,IUF(2-g;W=f0^A@cbRL[Qg.U)]-0;268F^b<8(H=ec#VBe7
WH:I8,Gf9NFK_&+dY(P.O-g;]K_1Z.[C7W3UR7)#?g]>1J325,-b:8)adEe.=+&d
DQF+b=eAT1f0>+cQ_@=UQ9\^dc?FH[BY-8H+(4Z(a,&9G(_4cO,cP@36gHdf2=^:
(VT]RO.4K<Se(K&GC^TY4/Tb\[:TG@GK],G+=&IDZWbe48NUUeFU^@77FQ/,FG);
dVB^@(>M@/?+#]ec^<+]LB=eg-7:+:H=)[H?/>deOHYZ#2XSF[(+KGHS5abIRB3.
M^;Y3J7g#,KVUO#I4L07R1@LbaQe(&7.D10DUSC6([D1NA0;Y.._UB:L\N[PW8F7
L\?0#fJfUB=V9FU.>?IS\8Jd4-9X+=N9C;P_\8f/Jd0@GUZS1Ic=5>(c/B?7ZgX/
2P_ZE7V2STYDVdV:X8YcI^A.4DAH&1UIN:;>5JS[HQ7CX/3J#G_0YBDK[CRHb+\a
<USa#?2cJNed=,DH;>NgZA5<KH=^;Y^9DGf&WCP8Y#MU+SUIZ]_]8=Q:YUbdCLKZ
)XEFfFRQ+dP4U6=fW=)PS:8W=Qc9XgWWMMYXN/=\2Wd]F?:#@,N^=2EebZXe><46
,TC7PM4X+V-LYVW1C>T.[@&=K<3>VSTV)ecS)T,>,PaU9:DQ4S?5Z-:5+)\OU[I3
209RRMNSPN_d(?]/D>#J6)U42[7EUcd;&NT@@##IKVg<WT5W]3KNYg=?WMV&0/YS
3KQM/Zcb>UY(WYVW@9e-[/T+F.?A6J,FVVUZ()IbcbIFcdTT9FeK0dG0MB-:K7Y:
.QX6ZELe8OZBW&C>2NPJO8ZO5J:,N7(72.d_bB_>7HaB\OD:Q\<Y,Z(?FV@M)W?G
gZWQ-=#;PED<4dSLY/1P,Y(J^OYSKM#>TG;5TYdISLY/+55;eJDaK;a6GRbgZ?fL
@CcN&Q3H?-W46>MdL&+?/TX]IYK\0eQ[bV#?fRK?]M+2TQ;b2-?73=dEM?9GLfg(
SCEaFC&\8N@D[,<_GN,\_SA_55fJ4\]e-P0cAJ2K845O#bG)6=FHYH]=);XFTMcc
8G7e0[-L2eE_U+V.c\7=^.)+84V#EH+e4DLB-,g=Q/>P^gN-b5[63P#M97G>_];c
eBNB]R>-0&8>@MC7H@[RWdJf<T/?5&3>dEb/@:#@e,T2EM7+aUV=IKE@fe/_0FQb
LAa3X=&8JI[,:cTVS(NN40>E@+K-2\F):Ga?B4:f4PP4<0cIU;[NU.6BMZN5Md8G
g5-,E=O=)V_QYOO]^-3_d_Z,[X:JIP;PERbLbF8A-8NC:,Q+U^:#L_Pd8)GGH]f#
O;JW.J-]WM<5.Ke^JaNgNLV]M-HaAUEK=GJ[FgTDYd@?VD)aFbBZ^MQKVX4NHXN;
7S&PG(+YBZX>FQG#@cW/(<5eGIRcX?>QY4#5Y,g04I.Yc@KO09-\0TA[e,/=24;#
F>]F_[LC02g?1>O5[e=DH5KG=5.J3AI&=?X.L5c)1C[2&EW_gFa]c_:9D-9K+g;6
C]]BF#&bIA6:2[c\OW#)d8>dFBA]d5:47PQ4J</aaeDYM6_)PIRY[3^O\4@AF_4a
@ec,)=53b:8-6TKaKJO0\J1HK+;\T5bfdVBI8f/Y/:fIFHYR+:@DF1d^V>&2:HT8
23=3MfKa4f[WJH02/1,5,gbW=OS<PPDc7cV?]gF77:1([<ZR:\F<6+HE/L[IU(XC
(A3XYe8_KEK-,^Z3D+;deV#\R9OP9bN?D5?W_Ga;\OE@M0>C]CWMZYa/-QS^TM0b
U3.H;-e1@.#=6S>ZG2B8#@2UN>HPPbI@;/>VD:#[0=g26RFK<UO&B\<gLc=K,]1,
cY[UT-c/Ye[=Qd)7NLK):FVQ-ZPTG(JM.SQ/YIZV5YGR,OA;+LJgP5DgU)^L7U&M
aaH42P?>-E71gD@\GN#O8(MUC::C>RA94gU;?LZ(78RI/SW+X0ZbX>C3@)^,>g5;
+4JbK4:6EAMLNR_e]LY<)2X+=IfBQ)c@,deA&KUGG#9fC(7eYQYg<RR#IRW^OS#K
&F8=KLK1EGUG2S/Y[D(PTg8T43Y5X7bLY=e193HA&Og/P?>?aV[aN[+>EIgEPaH8
0MWe42aKH[[<)4LfX78J?^IH9;^P:19C2D&M9//I)IgBd<4GSI2VADQRZ@XLa2GT
&LA&/.&@cQ:(?g:fV=U2#3:[D+#[BC3@f=PRIda7:O9JD?PQ,CR3GKYY8QI+XBSB
J\=>DSJ?&27KU/c2N=.6:0UX;BTQL9,=dV[\aa6NcfBPa6L7VI1Jc;32+eDe[ITI
Vb\J#)c3=)P^_Z+=F4gIY.=(5:>We@WGOL97]:>K8([>7<+:RYNJWX:MWVAZCM.d
I76BQU(9=)OaZP_JYbH:IWDOGK]J@a+HK<H(W,)C7,:XOGRYMCUEJ9ZDF?F;B-9.
RLZ\A@2C#^D_Q>V;)cBgD3+dKX^O:@#&YXfRZS56T7+D0HA:03L)BEN#5P^<c5<R
N4JdP2?[O@@=J1<&86WK#gN)IT(H8>D5K#:X2]DZ77&SS_?FHFCJ=/3WD1/?27;c
ABEX\IK9-@MHdJ(:d0K_8eZ-6S-9J<^e&;ET/MAR#IfJRJ#[;fB)bXX=,N5PQVIW
Td=X;(/21g0IB+NL^0YUITadXQd,:0fMWRHLS4)#,^^6HP2T,7?,:B=G24XCUcQ>
3DRgA;+:M@\_A+5Z#0I)>\g:5<Lc6251E\=2=1=)/X@E@036COgSP5LSg(_=^Zf:
7.dL]&5.Q=MW^6G7&K:;U5ObL)6ReNI\&DKbf8Y6N:FCPc=^Q(<76/994C4=WCaW
-/SDMTe#B]3U:&QA<fY.0[@\e(?f9YB93WXe2WTVQbVH-E/92:4T\OdK31NX.?Ag
5TO2W;^_fERPYeR^(OFJQ=-K>g)OW9[c5<O6<)05PdaKI.B+6#9MZT&+]]CPP4Og
X2<;]W5bHg,Q=J]5^L9S=bL;(Ob<N]@@CeKd6+[^&+BeD;L1aAH]=]Wb>?YLbWW]
A62:UCRY=a/C+17SY2(VO[-)T^aPX\9#_KdOFK]VE<Q3(JLU7+>LS=L/d(a;&03L
@K9fYA&MdeI[c^g4/:a1@;c(W(L45a3@\)SS9YZL5a4e+OTgFULU;T-.VbCX@g<c
/f\.JPS3(?0ecU@J<_/9HTHX2UQcYXWRV>L2L)EPF6MU?=Rf+M.#/[](+cBa(RHE
A]@KPVcXTQIN.+\78(#M.(ggE2G;VSQg<N@7+VdJg+5FGCCO9LVAZWe8CV<9X,++
IcCMbQ&6IY^(ND8:B?_e=W7gc.e:-7HATf\2,D8+@g]/#W=9=@Q/\g;L88=+U,a0
Qde)O6f^^91@a>X]#(5?EE\QfPT^;E3TUP,#8JC\GF@S.db,;4Z9QLaLfI7c::Nc
TZN/K/9GRP7c2e,18_bKcbE+3[<eM;5N/#/LOO]68T&WS:Z?B60CC#MSV&c@59ef
O<;6CDB[SF0]]U?#2),/+a3^;KK5NI#H9XSPP&#]/a-OSCagHO,QHE#2?.K9T&@\
IZI\OHK-V4XRe)dQ)&[S?P#9R]@UGIX9YXO7Pd3/JcRg&@]JMBXN)8X>)]gVYZKG
N7FBZ&UcCVBLHSOFGKNBXE?F:MKg+cG/TS]AeR4aN-5Z+1V]/a=IJ[\-[gAL.0aN
fF-b0JYC6_JU[CGT@B-N8^LU,+E_G]cVeJ7)+/.aHP#K0]&SbWN,)^E:dOZ3/(<#
Xd+4BW7AV42<L3BQ8JE#?F&Q7aTG]J7)O7AeQ?;I:@X&RaH7c#E148?N^Y0AX[P>
CGLMFK:@13-,b4f+/cVVH:eV#)<^-4>R5f(RG3[P^DFBY4U:@(/CJ-S9dES6Zg]8
6&13=1=a@X(3),&aK(5H&P5PV5@_1L-U[+.W(ZD]3:A9aW7-,a@\U_[VP:&ZD;d=
SE)Oe)32+c]J68cg]12_EWA2TDc<(B[[d@/FFF.ee[NX)SQD<AA;1;4#LBL9a^TX
B4/\Y#E?fB2X7eY4^<Y,Fc7@EWQR]eXX5^<[]4@31;.#1T18Y71H<CLG/JVZCD;9
04IV-^:W6N5e9@\M^HKW1_,J)b8H+7.>SJ:6@c8+=9IPISTN4U.H._8W),S:0a1,
EBSRb>1<A3\(9G_V4]J@MX+JK?;5[4d:&g>3R&ETfJ,R,LR:_feV<d-b[\]3H6gg
ZZV42TM3gZLZXS#\>UV(ONXg\=>22Wf_+[D&B4[W0:]0+<NW5P:1,HF;)-XB(WPK
d7>,)b-QI6^.@4N9Pa95Z58(Y<c_F9)&RHdZEe,WGLJAb/=S;5DX?#d(>[/QOIGL
gPdV-8<9[<(ZR@RD-G<I5B,508)Sf8cS9WeK1XfOR7N]YWe_eP>0R@W:5Lga33;L
H@I53W@ZD@SO,WFSBTJ)KK<c:2Z/;4aNF?ZgZ_Q0[FQ2a?6S]E^cPdWG6/(cc&7(
^M\3OB;4??W0/_@6.0M]0=56B]ZB;-J2AB3JDJO(]Ag/_/GeRc\[#Zga,DacV-F.
_2SfR?e74)R78bF/QL2KWEJ<>31&L0U;-F-#C?0W]V6c37(BbL<FT^Cb-VXd]a0D
XX04Vc??(6&P&MZ]#O^\T8M]YK(X-<6^KcTeTERO=GV&PAZ4)dc^9&I[1MT:/=<@
X=POeU(_cG#D_)Ac4B1,IY;FfReF612A89(Z&FSZT<+,QdZ2VI]dES>Ga/ZR:Kdc
@@^778JbaQHVDHK;KCNYaK&/<3_d3fI,c2Pbc@cGHB0^)c&D44]]B>&3c3\75^<a
GFdf][XX-d56IUA\;K03gODO^/NJV]cd?^LT_1]V5d0,^;W_@(RERX++X-BeTU6Q
_OYI]C7\Bc6HJZ?)9)W];&e9:?9534A_W4Zb+;c;e96ZE@BI7VOS9^B3K5+6CU[\
N\?TO:W[_A05>:>RgZK&&3BcM43_GV7bEKP2[N9=G]H)1M#329Y7acUgYE0NJ;cb
@,e]Bd>bUWI#0QLbfcI1X]3IY]CT=/;DKf^DL__;&5(^22\G>Ua=aTZX.f2M^I1I
GVe\&KC&WN2-LT9d+?^P/J?12@7:bQV+[.&TA[VS?EAeZQ4ZK1D-9gL8\c.UR1d>
5;#c7eNbANf?3SRHYf01/b@??7ZR(4KP6U]WV\8]UC:,2;8XN-Z:>K[?G6YGKeMW
1U=JEYC_fCGLQ]2f06dF8.I_T#81gUZB])GV<@.(C8J4[W?_7.HT>c@-RU.K)#DG
Q_;aM2/Y-+_a?>1)?M#+2HPQU=R7/C3dJCF,8A1=-\F1INJ]:-A=PFcMbg<34(Va
f(XW@>8+aZE8\FA#GJG^+&PK=fKST@9L]G1;ZadC_\89DVc>9[DQ6PW\Y9JO_=Ga
LDOJ-O=d4S-_aCV+RM&_Y-JV;X1SaQOKC[bZIXU\WX[:F;FIAdMdJ1)VgSF+V;U3
^]@[>2&BbCY6ADT453]X8D;61)S<B_EPF>IXZaWgXPf_9JO]gQ1G.]L].-8X7UNY
9--;LBED9HMb8BG089Q7#_J8)_\V8_ZBcVJbf=;8aCEaO>NWBYZA#,JeeUAW?KFG
2RELMGX(AX5,)57^&OGagfBTI,bIL+6C?#aRG<1)Rf^ZRS.:ZP5;1g;5#+9e[;cM
eU80.WQ==XaNbdJQ<Y8(7(gZg4dW-cE:UPeWR\FIVZ-V=;V;;O)8+P2F6HRa;HJG
JRcN[f&08?VOQP.<3TI,#6D\G]K>WLcb-B5[WRO-YC6B\GA^C\Q[;bB^VP>(83X#
fH?RI:V(A-,&,Q6bT,Df3YJ?6FTCb5aJ,JV[N+0.)C3J:YUY.+CgE@WL,59B>,RD
+P,F7IU=F_M71adC[3B/+1K36PbGLIJ5gM@;MD\7X_K-^UcZ2)32VR7d6c[TF__J
>8,LC2aN23UXV_YT=BSZ@L_Zg(D<E]J8,e&#1X&9F;BAA1UOZR@QJL#9>N8c1T<2
S-c=W55VTYH8>A3E5e>IV^7J#DA2BNg(5Q+45MeS(</^-6,8c=[I.0WKWBdOV]Y=
aE?+L^+L3GB\BU1J3:b32.GT-9W0?3],L(),F#(Ub<[J@8+B1@[dV29a9e,L>IJE
=P#=Q]5>;3_^e&M@:FT^8LaD643gd)QH:C+gFFF=<B#_#ALRAPcZ-O,HWH;@NK7K
5]\DJQ(;#eYC(6UX?VOfJc9Ce5c6K,+FXOIT)ZY;NA_d6ddH;_D5G58G/FSH-[@F
<5]IPB,U0-?YMUK_)BV6/[aX[Ed8\].VD]63H[Q<FO2R?bL&R@dLUfVP^7MFVLEe
[B7I/#4,4_/];-B9c^A[.-;.S(DV5O.HTJ--JL(HZD+]@..#Kc6OCH521<Y@P_.S
DY+HH.=(a/c+@J]W^F>^97+;]cbXD(UJ;eCTSe-0FX\@XLdNJ))V9e]]K135e&W.
8C]_-O;<WPXbU84eVP9]+<+M@f[BW?ac5+d4\TM[FVZR72+0SL.Ne9\BJK\_,g0e
(Q>AE=Sb@:9<G,Q,3_U&.1;eWaZ)O;e@ge]B@9+c-=FPdNX&b5R,XJ51]g_<-<FJ
cR&cC@.#I4QdA?aTg25gdP&WQ@UXNYF6797HD6:M1LQMXMJJ32&4]e./fIKWD#H?
22L;IOWe#Ia]#e>)@e#Za5d@@QDE9bK;&GQ1<;ZI7M0Ze:YB0[cIWOK/K)U/^9TF
E<?#a/_WbHX/HT/8K4Z5:b,Fdg+#aC@cWZ:d<Z.(Ad7eAc(2X,II0;7DC0.EE]I\
?\P0Q2FNCSXZNRBD(d@JPCfN=g7LU0G3SPK5?83ZWe#0VY[GLVg+7Hb69XPccI)\
;f5AYc&=_JYLL@LKG.N;g65+;P#S=LO@=U6=Q+?J?)a3V@AP.V6UQU/5gMN;-K2K
deFe5<.4&ROR9CF.(@8OD[]];>b4X,JZYe.L@R^Zb;aH45aXG(eFXd,C&^W\S-45
@:6.(\\EC>OK99V2@/RT9\@_8G4R)a&PcgUKK=JX4L&aE6X-&@c9c;=gJfSgEGB9
-Aa9P-26d6dVgCbg.7752aLB;04CMW4cC,13ONHJV89A9,e#fCGU1Mf+aU:=+8cU
dLBA@N3<N6\YW;M34(D-YUKdD2PW^NP7S6.MJ/VL3FPG58e/-fZ&NY7A5fIR,3AQ
)3LY,Zdc:H&VT5:__99Q+bW?4QQ-8+(aB2He16-1VX1\JV&9V@>2H&(S;)-BZSEP
B58(d(Z:LV4[(@cR3-P+-g1Y;?>AfQJK(7c\>H.P3_X;Q?,8f;6IZ[6gW_?/,ggP
USTLOaX6]:4I.bKQ#g,7J@1C[]9.;7@f#(a=V0<8)?(-Ca/(2,ISP6Q-Q/W.)=Ne
HB7.^?He?Tc8A,VOb5OT?4WHDC^EdD1,abI(IA?G&1@QU<V9QJ9(gT5c6E(N++SC
^V5_G[]Qea+FSPV/#F^E.ZS=BIeXW;V[IXNPa&W=E.=.W4\[cS:,YbQd?E[gK<<T
MQb1S0>/;D-ZZ<GLFU;Md,GNBX1,^>KZgGM(\c9]6G4P[c)W=_X/:RRJZ^/Ve<QC
f7?FgS\XE)8H+\Td2QV8()7OEV^&&J=4M7ZW-b_N/KcV:\,@N/Y2FHd4TS;b.=Ug
4ML7LKJYb<X8M+3cEZ<+QIDTE-?(68DW/LKgJg\>>DA5@P,?.TFe4>#?8_MIXLL8
C_CH75S7?(ED2AKAf[)C#<VA1+><&Z([(SS^e&&11e190]3=FagN8d<#8-L,>X(R
+)6AZ?X51VH6PI25[>1c<6M3JKA-a-e]eSE#)K+,bTY&0F7b;[W)+23GU5V>0:0J
WF#-=NVc7Z15;@?EF\R97NVbY]3S7WRS(^Y[1-+.O]E/b/b.Z&NER](L?Y?8:Lf5
eTYE8C&fQWM^^129^Gg[TD=EC)0&S6f&PAB+TP-dG2,9XbbAM=<8U6B<,g_.3K5;
b:?#^QM1@I,g>71WF.?@Xa+_PO.=dDdHUDDRd8QcO0PH43g9gNTf=3Rf3DI8c@4.
6LVc:PL#3DPCP(dd(AX,[,B:UHU5XVT]?f_Xffg36G+>L9&IYW#Sb&+MM9GYQ:&V
0ScE,O?FRX0(-QM-ZPPN]6c2XG2YN&;9,8:L/ERL^VEY.c??;a?aG/6E</.SAW)>
.6PYS[K;+],2+])IV71JO.117dT0)^Y^g)A9_GX>e1HYJeYKBGL6.]>XUc3;U,g4
WZP_[&:)&XE+f=[C8JRL:Z2KZ83[XfCRegK8Y\5f++b)FXUVF3g)O1<P:#fQc[HA
377&HBg/+0&_)VD-YF6Xb7V@Q]BQ1+3>]4@T;2)3aL=G[FMFZNeHa7(f>e]\57QS
<MZ))RacOE2A94CbQOb=M3\040=_,S\/--R5XT#E18LGJ1^(#7TL^,B(>QSBc=-[
Fg?B]KNZb>&DJFBSXO(<(0NA4QD>+D@)]ENWNBJD2ZKa2O/J85cbL4cDFA:B=4YN
:OR6D.XKP.FU121O>@[XW1CI0-BT>_Q^a]=Y>SKd\+VDNG)_5g0F]WZZ4O>_0@KY
[<6ddD+.ZL17Sf<H;238+HZ9VECX,DbVJ8,)ZBXV^+,7HY]3T>G<WH3)d-;39Z;[
B6Wb1Z_C&;VI+?a_L:M9#X-EOZ;[9[eBgbd4+#-BE:/&2@6>VCgb.H7-S6F,MZ?/
PQ0V36ON&^HcS_5RC(fRG+&0[T18(ELf)dW\a#0L:>M6A+HOO=B<Z@E6&49XF?E6
#DQ9@L42TVf?.aOPY#BW[a#L0?c8+,a+8=X5?N^>X=c(K=)Lc^ZG>-0d<NZ(/Lg/
FJg>_R>BMVEMa;4]OP8^O25_<YH-b.E\B.C@RDVY4M29e3Z]EA7\Q_K9_gHRES2c
+?7[K-G65EZ.C941\;Mg?aI+9?&9CU3<DT?]TZ638M?.7P/VN^cd4+8N3RH\E:-O
/SPX5f>f#LF_4I7,>3AP^)cKZ#82</8HYK<ZA4gFcaPO>_&f[?_fP+g=..b:eL^4
P57=YYg3c5(2dMc/9&E;4E>#c\C;dHUb+JaS@LVX,JgW#Z;g39^M2\OZF]RM\=^e
69D-1PKM,:24b,eACgJ??8Q@aNb6PTd^1Cb))NSB3Z8)=][5[_.O5_5UEQ4)VTe^
(E9;TVgO+6P1gRZA2eWTIB7a(e.DB]<I[=3#</_aY[aK4K&;V8PN3UE8+15Ua.Y0
I],N[4_F3W3-,@=bXHS)-IQSILb_\S&&FF)/cEMS+a[f@O3Y,(BRf6.U(fUQ3:c_
@,9[^,W(6,4M9_E.gJ?BG,)H:0WG<L7=^BANeGSIf8\Ka(P=If7_U4]Q,:3N-ZFb
-IL7J1_@-1;1Zg&b(ON6@]d_+WS[\&;>@T-/H>@2,RD)@bLf7I(W2JcU91X]+aLa
9V]F\\>W.16e@eF+_,<#L\C?L6J2VA.6D),@W\A+1/D)+\-G4be)<=MS[YY^NIYO
ZgaBFOEA+R+1:VW1Z9>0&SNB=U6@STc2@[b?MSHYPK_LMee(-aLDBHEE&.H/=V-+
9\8D4LO/WW7XP,/._GOKR-A5S]_<^R&NI8f-@=^FQ0(4OUfKYNMZG<G#^KK-9H/N
1;,R1F9c7+10-7-+Sg.=X@5:L:g-Jc29,+M#;F5O[X(U\Y8c(T+.=]HQ&9LYBZXK
e);9dI2,5)\?FO#A5F7g5:KJ/[).7K^>Z>Y5LMU9:E0+D<_W^#C^@c]\Vg1WN+OU
#<1CSR)J<>K]d0ILbWHK.6SL2U?);8ZRK0/K-2_HQ+S4?O)._JbK:+a0TODRN,HP
(TW90)-8d[U9&_VEH9PJCIg782b)483@QS/\gMf&N1<OH2J8)5@D1DZ]bNM3]NCH
Lef[X\HSSO-_4UQ8a,e\@E7J+@86g_e6bG]G_]QXLaa(X>55Q@ISeC,TZb0#6:f+
2Yf2&?feJg1WAG=1MV40E+cIR5\cOaN20S5N2LY&>=e+b4G4W2\//>7R?d2eAGCe
:4?W7-WG:U[W<><17eGI-N8OId<0Oe7]c8+]RIXe4CbF3cZ-#UAXR)e\FVS#Sdb;
[FfF@4@A]F-<?7](X@YA>VGX[5#&0Y<K46CWJ1dA5NGdga.DZ]-X5OZ_RT#3.3QM
01Ac@F^gA=SY-+,0d=_Zdb5)@IF;,db22F]55)>]f9J82III/RF=A9VPQ/,A#7RU
3=(QL1O25G>RM/_=O^(Xf-4<8#c75J8M?L<LH.YA8/YJIg<K[G^&/\P&Qf=4)HCG
N=VI)ZdQOL-_Td45L_fHMXYHLc6E3L#.,XG)8+f14J:RcTZ:Y-(Ie>eOFZR0+8>:
3L2Q=(/078J>T<GU+=>E(D+NNYP;b9Ye?3<8/(C\T:bS:F-TN3L+eWQ&P@9^W:Af
L58(3VAN[f8+D+GCH6d5/OI<QA(09X=8BH(UEWSRIHM(>N8OY\U5O1.WAI6_:eK.
e>=552]IVEE^.L9<cCJ7.(^;##RNP=O+W;f1#ZB+8bZ+;46Nc@[;JFRXL8H(SD(\
3HHgH=>3-4)1&PJ);P<a-fT[EE(LMefKGWcV=0O;[_-/R463V[@?[I/g)A/,E,cS
bV#7\:L;4YJ.[9c15=I-2a>1<RE6Y2EY6;b;\8Q;]4/b>cK;2fVRQ7cRP1eAI6SC
P9RHH1T4b29M,5P43,7SJE(g>60Y6fNS)T3(e?U1JMK6GPX.5fH^.RDHVaBX;SM+
Ze=AQH-dP_SZa\D9fU31L;>0YVN3B=JR5<C,O6Sc(e./a?)4N>>c]LaHP(JdD3)/
Z-L3g2gVS9,4R7d2&b9/Ddb0deQf8b67e:<:^]d]>)GC1::D0-ec=E:8^MU[]b:O
]UKCRP:_)B)@^/08@Beg3V#QK&P/0:;-9U8G2M-DYNHdZ\K8C8^UcI)cgH;.1GSB
Zb^KbUdCX3F??5_eQDC8dKFV6,H(K9]ac6&)5.+<IY8X6Jg\IU&baDMA?R<agd[(
>SVE4Q9#4W&-gGXZa?dfeQWJT:SPPb35^C11)^#/becEd_@-^R^V(DJON@?XZHJQ
_BV8]9YF@DZ,f[#3D<INg]c<eH,:X6@.M6(-L,Y2WJ8;/g:]Dc+_CP)73>SJ@D8Q
33LA:Z/X,QNY-_0Y:CK\gJ2bI=e.#J(\\21(e,KE\5&RPVO+VJ#23?5WM&3X]e?C
<\K0E-bUWQg?DGQ(0:N>@#Of.,J3VR_0e:cRQ8O-9);10M7YQM[GHA)KJ)+M-_:K
_UP(R1A_He>?fYUO,Kd&0FCXc\UK;eefR8>=),2SNLIT,2.FCaNH(N:W\TBKKYT?
DdGNZcYe:fe63&QZUTaF=aUMdPK+F\]9B2.:Pb;2Yb,cf:Ga+UN]aS]]_J2d63ZE
Yd0Q-[IGIfOEA&VK+X5UO9cgc6F8]=TH?VRFP,@J#X)W\IHf[(P&:X6dbL^R93Hf
3K1&2De]K1>O0:c/D&=,K\;a.Qb:RMR?L1P\Pb;Q6P#,#CSPMD@)_#T@H<2RX2)^
(X>BN5[8S3K=AS[N)@Oc9Q[<=[L1?42U#;VT:GaVAGI2:,_QgL^HS^M,H.Z:(\DQ
dYO-U:Y>6_;c&@O38O51DP8+W8?eYQdL9Ub#T&dD)D1Sg8N/AH/JV-8;3[bW#Zb@
X#AJMb1+KNWd1AYfeb/ND&VNfOc6+RY_AWFCZ;YefUW,LRH_BG7N,g25FdVYY5PV
g#US)X:\A&VC9FAAYQ\AMSFa_Va.FSAN-?-KZS\T2.U0_]FX)N;X&?.c5CPGV@2B
YQ&BH250V_3Da5J8:eC3;Z(->J:d(UVI\U3P;N2RT:R@fQ3[Q^V.@,O;@PC\g7CU
Y4[)fC7Vd+3Vcb,]VT-70O_HP?E\AAD4<;g-6LH?8:ZBIg;)C</TSC?a?1DO0F&1
[35J#9_Z,@BMg>6-,W]QAZVG):A[fQC8d)gfIDZd2.B5d1E7MN,[HEH<]7E+\WZG
PIIIFF5=-5/H0HZ9KaeH:UL_7ONS5b)+5X2fX7(a0(Mb+c70_@<a71I2#KfQ32fN
^Gb7?#Eb:E1OWD<WHC,U\;AIC@T9.WPC+gb]PPWC]M;L0=^28]Z,7\MDV3a0Y+9L
^?Re\&J1BWRa-NQTPVJE+AMZ<[M3@PT9d[Xeb9eIPIBb#XUKN8,,J:.XB.N#XT?@
>-&7HY:F&\TUTPAdS6]1N(Z(AKKaFNG5D[c#Vf37RPO#J(/K&P<:F=?PC9?IY<AC
W3I\\gc]2b:].O#R=EY9)c.ZS,f].2F(N^,[@OV)#W3MUcR.1[2@5NTEL,8<Q9>2
=JG.e<aJV[QJ:^]df=4-PHYP/UYOK0g2KB_O7Zd>@HJW5N\R6(fL78I:<I)dSaI1
W8U3FZA0\aC5\&OH;1,0QH97\S\-K>QY1V1ZXU]A)(L9fSYP.Z^.0^@8M4Y8=0G4
eWG4O:\6S6Z^H9B(FX:7\SJZBLWb>L><7Cab<5B;8;RP#A\WZFOceI:@(0fDSU6\
VN.1)88:E]W8Nd][J_&4#_,gD-B^PVUA:2BC\g[IE=P\;K=bY9Oge1@SITYfba_L
(Z&?\=H_/]TA[=MS<HVc02&-/FMbT_f3Y1<I#]>0RFYRQ5]S,=8,@PL6+;1:b-85
Ac9cLG#eS05^81.6JLWPd[OV](JML)@,.Xe#?H4d\Y.DgYRPS>=UDDA14GQBVe20
[KaMU^>AI>2TDXVV14V&57R#3;G]LTN[fJN?+C4TBQWQ;-.3/=,V@eC@/X)-(e(X
Y>&+W9^H16,Y2L3XH<(e.4+/^JPKX\G_/(==H#Q>YXZ/9\&#81<M)\TJFc<+;]2<
2N)Z&>ZL0\@,)2V+Ng<bA.][1<4D_,<;C8>WH342cED/@4,I?T?JZ(/EI0H>#GGc
.cMQ4=4UFWbc.)->;IfI&3EC93Z;bg8aDNHY\M,V1b>Rc@A,?AK&HYfZ,3>7IUFc
353a+OUUPO(8KP)TeATGb]@aMKIeW6_]]Ea[fTcZZeaWD[_P8Nb5W1X\M)D:c75Y
FX-NN^TQ6RJ\FO#]8-[+)[53F.Z]&P/(H08[5f^gg&(A;Y)OL@(b6\CI6J+&QCd)
8R=-2beKg,5Be&W;7KeWD<MK>^H?N0ge#b&,F+-G6cJ7OQI1]AFcfC^-QF3#P.;e
DdY5a8.WV=5?H^SF-83(NMS(\bXS.]DVe)SXS(V8-(6^_9g5=SAe8OQBSO-71YLX
8.CWPgRDW=-3Cg<KHPOdWCU^R5g5S^-,bIJB:T[cCTB+6UG_10>f31Pe4Y:W[(I+
;HHDd5U>Q^a_Z]bJ,4a0eL9GTK4^X.f.1U(T,aO1ZL#G5UFN9@(XH^6PZ87b43e7
@F?U4S=eE<-b4g?G@7\CVCREfQ=;JB=Y]cdAWR82@6O,J=La>c]fSb?8(J6NO3:C
_3OU/Z?(0g>0Zb@O7GE3U8_OPU<E2BPDDY.A.WOBUU-.V0LdB];AVTBK/?OID@E,
C-]GDIS&L.RKLXe=7U0?TT,Z+#6\e&[3)B0gMI0STMQdENJFY0P9ZB@(E0+9.(/a
27ED>\ZJ4C+Z-<A#2.:LGbPZV(g0Z@c(,=GC3E51e[5&[S>eGM-5OO54:c:]8X5_
]UCb4I;\P^KZbK:O61X3gE90bP^0W.ARfgQ+9PWNc.3bbD2Z=9T[Yfgd&@1PO\@6
&Sg<]d]J1>Y2WXGb?O.V\f:CF>@1LYGBT=1>Tad<GaCQ3Bb:JJe0.I&eY_B]20:2
Rfg=C[BAKJ=YJZU,[gZ::aUW/MRa;WR&3Lb3++;BK>f4-?,)0c&fGS6XLeJCaO8:
Q(36a5Kb7<]:[Q2.O4\AE33Q.DA_\+EFdX8gHGQd=+D]&^/cX]A>3-=a8eF1QM?/
B:-L-FEABX7Y<>FV]#LZAcKMB/ZC=XE?ZIY&<ZUJMcO.R,9)+@NK^XeA7;_[<E;=
>Q&-Z(7,OL86?B5]4Ub6AM8,#3X>H[(BCb6<_\=V)\^YNf1@;M@SZd60eSg?1V1.
@U^:#4/.Yd7K[.3]f-P,KOD:eJGSZ+[C6_912AA<W?L#TfT-7[BTNH4S]\b<T0=J
6;C-DD;eGDBU?T,fG38?@C.TH@XGOODaJ,d]bcA@&=f?#b+/PcH6\>0GZ(1#^H6\
]eBgf7-HFLXP\9)bR-cWUI]#Pe#.5FGFe&eGT6bMK5aHgb0[6;^Mb6OFg<_&06M,
)M2Gd3AEaLEQT&B+HS6(LS06<,>(3Gb>ZFJ1S:T:fF/MVD9;^MNX,:WdT<F^dJEO
6LLL\cc79dD?6/gBfN.?NRa.NSX(>YTP=61SWTFTPS@b.P#_d[M^FI]>RFJN8d8Y
9Fc+?a9:,OVMTZNP3^d5+HS](f2Q,X7X>N5]O#HK0O8+Hg_(=H)aHR@1+MOY1B5/
S6_?:-II=]3UI6dI&_>DdYcZT:W?=0X<bf(XIeA7=Tc8>f\,PXeWU.Q]C].4?;YQ
N0#QSdZ-Ba0]dEc8,&)K\E)^<6,Y<106g:XX.4g&>AJY?5?VDPI5SQJ,>@\\bZP9
1-I7bgecKaeY7?d\]fQW4CI5UM)BA(;-=^^4Z@13/(-Ia]gQ6(NKfK+1c#a,afN5
ZI5B5LL9RLW6d#YN0=/I5&^\+LHA#dFH[3ACPR)<\W(]PX/,3eEH6T@/Y3?F,@DW
M2@E]8F@+CY9HDL-F+cc<.d&#,S)_G^KV#QV[/U-/?>WL=5T/N:LY4T]eG.+f.HQ
3a?_5XXTffU+TK)R)c[]I/f&eYK50IH&=PK/V#R^6/H8=AZ)X:8,ZegQg#3/2V6=
aSXX<eY4AX8[YXW<H52?-RaJHPM6E9+KcSfX=A0QZcf/fGJT^aO=^Pa7C(@eJe3F
V.3E:P63XEPJW]S67U1C9-D?=-^+ACPKa<aF;_9cA>6NOZ<X]IVg4_71,0bNDFcD
(>f;SbL+]?[E,X1=dQ4OLN3H-WS1EMge;TNWYJE^3@UQ,(J.>/f_G8J,8LO/QMIZ
-=9@K265aUPJJH4KR0e<]Y(].NO<4G#6&]&2V-FgAOa&3TUBW<+KO?/ZMQ4F6GB[
S+V-aV?9YKLE.MW2(WX8U:?I#ONeVSa9K7+).YAVf.8T#I)TPKUIH+<;B#_6470?
+Be&V?_JJM3QSWZ7>FL#g=Y/1dP^4a/+MFb7VcLRTbHJBQ?g4T_CE&gdg(#NMXd<
,=VJeb#:JO5Bb0?Hg];I.I6d8J9WL;g&DbJG?G(+@I97[Y30M:BGSbRD)Q;^VG=-
M4[?+a#-Ted))4--H/B;=,CT-EHFV\U^4>N;5+XH8d7&^0V5;8N3U0B5#T/[c9ZQ
E2c5Y.)^,ZM&I\Hc8>dR]^Z:CdCHTgLV:c&:=6=W7\6>;E.c&KBdU95:5],7)T/Z
7H+/U/cFXNJaEWT06Zf6@8.eT1fagJ7[J/5#NLd6?_W<a1R/\RBN&1J\=1M<()X.
G,IVWcL-ZWLPU&FFZY<@;]^96(R1cCVbE-)INZCS,@\40&P4STRAJTfWdLE9f3aC
A@AC>,.WKTZHb&g6)a0;(0TEL>Z@5@[>I4;W.;IC,(G4Q[X+#WLXVR,08#-+\d5a
9beO0SUO:(1Y[B)0Uf+5F_,T0#b[,0e8:;<UcMaT)fEN9Wc-^<g[T.CI&J9GSZ>T
UC(Q95)\&30#QHJDR_O2-Z)ZQB&2Rf11JG=;-eaa-gVN?A/HG0]dQCQ1J#<BfZ5G
H2&CB8VI#Kb)eDFJ0?+>=(d+(E6CELO@/9\_:,+7f@&BPD0b4>G0<:V.ID5+J9fC
X4JMS7,VDZBgN?&)FfOP,+g.<-U<b[N4g8+@bFE4W;&e90I8.G^.+D>>gKV^EGg=
<M^XU(?-a>I.&CG:UK.FEf[53HLSZ20=WWL@+_XWaL;E?]VV_b)VE01@1,A]JJZT
MAg]5]J=8dI^/bR>d/H24JReTI7#+97HK8JNGI;?_DDc>8[@I)6EVH>R[FIQ/;89
3,5LNQf&aH7+1BK>FdB76^DUX[,Og+H#3ZfC::G.6VS,Y1[)?(1JOEc6#aMKD6]Q
-)J+dFNC^&JP14:I4JL-]JW4:4>dg(IL\].N22BZ8D7.1e)\E)Wc<0RfC?e@G6S5
CM513Z389Q18/J6ICH8\J5QMf79LJ@T??Sgd,,SXW2?1;_/.O_dIZLcUNbGGC1^b
9g;Rc\K]&,FQ_+[7=SAUP_@V,<8N4fYaUI)3fJ=G_LR5c<]WRgd(^8>XbI\H3IDB
:_50D1G-bDNO/GJ>O8B].N\QdL3?<X>S3&caY_J46L5YR--G,-_GR=\/L\f\C=W>
BaYZS#R\__Zg74@e,LQ2]Z5FHZ+<Y:\;=C:SUGO#d.fUN(gMW1,d#4UgUBGYND<f
gNG?b.3aRQ)UZd3S2^YOSacX,.?U[11541d(U+T^_N.SK-/e#]?6SZ0;_J#..K0H
cgG>VFX2VG];5Nb2UL4P]2\68N(AQ5O^WI\ZG6_d_8J19RUbD(fCS9b,OZ5,bO]\
=/RB(1BZ@7>NbNf:AJ;H_7CWR7V@77Ea[A]GaW(-IPRBE591BH4O;Pc?03;(S=,7
Pa+CWO^0W#;BVK=_e0+615MQAO[.-Q(0=@#?9&aMC4]SG?JKaA=+2Ed4-TV0]@4/
dNZ;7a<0IY(X,.2aN4[2gSC0))Nc(=J@]A7<f3SU\b=4Nf\?X+0>K[>10=).8&O@
7?Y#_W=8\R#PgE\BJ]baU_E)AJ4Pa_-4/JUIT+_\1LfT:I.X.d)?VUc&EQW/?HYa
a]>5/J,7?f^\CG4A-1?2gDg:5FF91WO+4^/C;1^;=3T-0R;K81dMGWb/GK/?]gF0
Q)693&YWgHGO&<+P]-=T[9]+/#6-M2A52BSF:HeafM>=CO_@H/g9X<Y[VaYC5TYP
:[,4g6)H359OHVJ=UCWWX^;c-3#&R7Pea:217M,^#^TQP-;_5]?_<DKT8S[g=.ZV
869_K9F[);;YP85P_dI37F,^S]EF=B-;5Vd9K-BdTW0<=?C\<I&Z-PcL]>WM=SP2
Q=fObXA?2:OLB2KUSFb7L.S\/A7S\Y\E<DB#(+HHfcEH9/^fT@6aW,A^@(N3BOF(
SS/=e;\V^6A<F#Vf>a3Ag9^U@WDJGK(7OUV7PWNR(=07M)_:YRXX5H2/)=UC4NS[
^.7.VOH6NZF[Q[YbeYLZ2EA@HeH1L?4]RaI(@BbW]2S<OH82(CAK]fDG&OJ&e\I-
dK^=FTSBTEQ@@97>;FO]+.JJ0AUfN>5YZ_KXP13__HEHAHH(C=L2+JGO\Qc7R5a0
9d2g:LG#;L)+DbP;>cA@2[U(CRPdaV.Q9;L2NNXe_G>GNIcVbgZ;#^(aLYU?H+,B
c;I&CQg2WdI^U@L.PWe8\FH;B)B)\O_Qbc+<53(a?J1,#R,KM:b0Pc1R8]1O=PKG
d214[UWW/LX8J=]&;?<b8f7Ec##Q3.=,8DDbdWcS[0^.2>JR2C&#VIBb0=b570T9
]aRA7LJLeb-49I_>CEZM@a-Ue39P4B79H.0FL\^OIEAdHBDEQ9[Y<g3JH=)C#f=#
dNIZG)QPIObdcR5F]QOXe3KC^<</F&ZbR)558cLFfADY\J4F]Jc<@V-C&M7-<2<:
:SP?POU?IC_-U(H9T,7PZ9^DLSUORH-=7:We#A\GfK^==KIU\#F1ENM60UO/T)+M
)85FMGdaS60O,#DA38cF:]FG2f&3<H60Md)I&dG>)0eJ81DJ(//-\(GU0c7-a5(@
-\8=#?;Q=Q\SD)QJ9[XD_bd,+WH6K#B[K,7?^.&ec.gKA=d:Y;04?eeL06YL\c6b
QA3Tgg=+gOKAR=:A&(dCE/)]H.a+:<&gG;8E<Q/dY:2)2LN0EQ)e0&L:;:ZN/;#F
\&SX8K,L6L=ec/&W8fZ439M-(,+4cN?.0FOB7KY<:<LW@MSE9JG]]Q)]?@;P2VK@
6H)Fc@0OcJ_ST#)JL0MYUV,N7Xb\cCeYSFPK^&Jc4ZB7_6QHW1Fc-?=9^fW,#L],
OA-P=YWW&Y,&CO,B/(\\cg5OTEMcK,3:UKCQ7KaTYge+9XB,I0VFg-A)SdL4EbC]
1VaM0:[5?0GXd7]2WJ:XecM=4U\[;-d\H?)PU>^,eC<;B7VQ9<E^<dR@\5D+aA)L
1O]:Edd>?#Sf7EcA;QZQ7@X>PYW29JgM8:5^MK^W74VG=9HU&JU6PAP_.^eV(:]I
)@^Ed<cE^Ub]GVJg92-J:F:G;PU^J^;AN.FD#PMb6.g^YU=1E9+UgOJ1B6_DSf&G
BbNacgB3=Qfe,?]EI+\#YZW:ba^\FBTXQ3:FTU-;6_/UBX2,XIFg&W=.dcL9.K#^
V>OI2b_F5]U:e[-+aU_.WZSYb(g(82G&9C9487S5WVHe(]IJ77&A0ZUM+]MXeFfI
+C1#;gAT=\.)fD99X4))F<;aW_MNbe61EA[aM^M.[V35dR6\#K@/\MC;)FR4R_DC
:2:X@JGc.aV2<PEDg@Q2gM#&2&]81GdEIg6MZC_^K;^5cS?4&LETL]MQddUGIN1Y
O.M]H;EJe;DI@J3P9TU=H:++RLeb=C1\&c3cb/0+_=@WA3),0XE[SJ&49(+W8:]\
>4_KZ+#+G41#G3(#W@_@8P<<1^@]<^5]g&[gK5U88\G>g3551A1<&HH>D_\OTS[K
,]B9EKRU]NXO:cA4P_Y&Z,fL]<d64UMd9G24]--UKUWdIOdZf-DHM2QV.>Pd1URA
+NEgH8AAR\7]W6aB?C1^Q\:[6CJ>60QaBU.XM=8Y4/KXI8^D.R5\cR^IA<ZbQX0(
^fP;)6HIgI&&3>E;,4,[gZc]BU+&aUITUD31<DG]L&Vg@_#S+-,J2e8TgcdOc[_L
=+D.TCBWFWJ^R,9Uf?:ZeG(M7&3J[CY1_M&Lc35PSN0#:GbWgX;VIfC:<YgA<_C7
2HT<H>=KBR8AR1^6?CD@\EL6ggQ43Ya8),4^3a91A\2<U?aKSQIK:cgYU:(EATCX
X@>VU3ac6@46JK=5HFWZ35@9;:bZ>A\MFL2G4;<f1M<.YVOB2M2>\,\2)B\Eg.U5
.@dP>3&]Geg1;_IJ,RaE\JQWI+fXB8#N6F:fg,ad\=QS.ZOU,8=)NIL)Ud4+8(2B
CQdBPeDUPaM\LN92)>&T_.L3g+M4QY:-(;U)=L4>HVR=?/A[G+EQVVea&?H2#SAI
#-9[).N7+aC4gZ<.EZ^IgO]E9@NL_J.R28<^?;-[9.<eGC^9=P-;AZ[:NRJ5[@F1
2b[P403X6A&FW<J8#)g@56EYd+[Tb\QK)75f&M^X)DRBSc+f#Ve:/e_YFO#e[&\6
G7-&2[TDD7M2/&a;G=[SGA3?IQK9#RG-K=_bGNJ3;df/7c68[YZ2)9_I0RJbM65=
M]>g1PaL=B35dg6Z,/YWANE[,K.OGS2ZZP+;4FKGAD3G^KaaC;I-1-#@LeM(W052
T[V/VgAML&)=Z8IU6PSR;U7LaXK>c7;G-0QR5P38bQI-<9W8.))(8E(<RF4EZHI_
4C_>Z&aM-4TAL4B<f)HCWUH+K<]dB[#gWN\WgaI^fHcNE_H.S2Y9PT6\E7U^Z&<#
UOSe_N/&cL8H0)f;DfM]NOT:?VMR^^_W4D^WP@dbU93MMF<4+]]H4(<F#CAEc,C[
d&S1PJ0I&OfKeUQEDU_]2H8\V7);5TcJ23_72:4@;Y&\0]^9(F1]bfE<>0-ge);0
b_LD\]87?fNC817/21MO,QJcO51OEJE6bP;#JZ^/ZCPN@\BL=O#=([Q\S8Jd;T]d
?VAf9-91-]9M/cKI^+GB;BdC1/4M6J3_UJ(19C<<RW_,^[X01.V]<Kf0C>^-U]00
?We=GM;<[?eZGAD;P2)W@LJE^>62)G_-IbYWJBKXQZ?,_=5D4[KBGcbAI4EZVPA#
^:9D4G9-GQ0UDg>1IA\0PbALg6)JC/R8\A8?#/OPR@/,MQZgJ//^I)f9DROW7T<\
TI_Y9Z]^e2LN?LgF.GPJR]Gbe5\&.?2;c0cG3gZL(OPG,KM^LOad\1TX2F<[<]Nf
7=FLWJgg>@/@R/^2FK?ebR(?)OcV_9f_ED_4HT3Q(f]+4a&cMI?g_F6a456]^bIL
8;8JIL=^5.LJ<=]GDL;Y2M)F].H5QWX\S3CVK?Pf6RK-^FaEF4W&^@4D?=ZBB4:,
GaS8U[30P1d>^(9=8^A#f?b3ESd8f:XTUNVQ/H.,_<d,1MP9gYePfI;EFI#98)?>
c+0?G&MA?T<W+-QG4C3W2f0009dQa\]U)0=BP)^NS?_6U(52?Z5+ZXeeYE#TX2A0
,ALggJ)eHDbM\<6X[U8Cc8fQY>-D2SS89EH<CU].E=58HF\1T=4T\RFA:2?.A<Cd
U(DH-e=4^DAY53E-=Je?@5CLacQG#YEV^NcXcEKDcB.f/\FE&YC4SFb>)->\;@R9
Q?daR#A2DJZD7\O]+dDBI@GK]<]DUM&#+Hc6c[&3><Be?-Ege1R)WS0Def(;9fJY
a80>2P-AASMBJ>1ETJ+SWOWVLHe&#E@XG;.HIQGTQ<<DDUIVSHWE5NH7c^A,54+:
O,2e3G]Ye?U.f_QPA.)DXJTFPQgdEWR>[^8HG&&XN,G?a:LU7\N9Z//T[Xd-da?A
ZNRFYb^:V&\=0b6#9B1,U\M^C\2NAC7B[VT5#Ta/:CR#;;M(B2c6<.PKSO@]W4<4
L8P+4gC96EaAI63U8\>F+-gY^B3=W?92#HEaKbbD?Z>?T(#MP@>TcDLDg;5d1P4L
W9C]B:8.0\PYS?4[#--=S=M66^S1=T9g<1APAMcGg8O(:/\92<^J=Q?g^&+_HV2R
>\&53=Wf.fKM)J6TFXg.Pg5-c5Rb-E56d^S_0JF0@EB?<\/8&1:8aZXb&77aJ(/c
0V^\KD:T,AJVZ^Y=M2IX#9BD#PV,7BX)1D-deQ@)^&I=Z#-7S-b:MY9dNZPB+I[T
FA(deT;.e(L2+_E/5&Za+@_[2,Kb=HPSJLROD2+F-([/4,Z=eTX/Q[(^][D=UBZ#
E-KPYU-U(2HMB7;2N+gee:+#LI;L,TLE<6X+/&,&F+6&ZZ^N9ae>gY(:6@Ed_,D)
I+>I8CQ4(1W^Y0MCLH2D4;&@7&VcK#fH5VA/fJSR-2@B<461bcVX\<>Q35&7:b>Q
g<4fM9OV^#C68_c9UVNGXg>VEAO?bfV6^&6e/D]A^>c)2/W(4M_>VBA,9].GWQc/
M8\ObIf(D@[4-J[C2++0K>\/5XKf2@^C<:1\S.fHKG4K=U[A;81[NS:/26KD[T)-
+V;?YCW06>8#.2T:N_\\<4EU&7=aFa1BeS13KH3,,KO3V=RY,f4a)NfJYB,)5?J?
L:2<#aDY+g3dU7Va;_F-FX2YR2RQ=C6<XSefdL/b1@eWI)/K4I9:D[8NNFK7e>I1
5I]ZNHQ?:1T^XE?Fd>5L6(&-+b>/FF)9dOVOZ+a4;H5cC4I(:F9[d6[aL7fIa?&f
aO4.S-RQT28.Z\V[-HQHVJXBNS)DQ/7-.5UVae^H8+>[0SI6>Y9SK9CCg(T+9&UN
Ue7)KNUeRWTW4S??D2]0NXdSXU3HZ;EF+Y(7_Pc?-Z;._bdQSFND5N&RVW;FM^1Y
8++W?CgC^Q)6,[??IP[b35=&\.BEL>XL(F:[YdQ.-cbb3U:d-g\POg[>.DfP\7Db
[AQ4X\(T2c/&aCBA;C:>5,N;Q7,W-@AeIGTQ/SfLf0ZfV0DYEgR[,b83;TL+9A>P
1\Ac#Z/MZ@)]fS5?(87L;S5=fbOA?GX55L3_RVKbUVC8LAR:9NMZL\S4SG:PPH?,
28>3M#7SNNFeXG?UG-Qa=)X5DP[SegC<CX4XN9^N7KU3TBLS+5R3;a6Ae1_JbX71
T?:W/\-;498]:GCWN9L&=8PY;_W5<B1fORD3a>WC&=39.WD>aNf?DERa(BF&<V#1
JR,6[2@F\(^+3d\9:-;a]5R)g79<6&)(1fB]<WOIFDP]QBL9U=_LeK-KT\gRY;@B
Xc74567/4_,22B^[AbgWL_(d+>f:SJ-.A4Ge[XJ@JMfe_YcRS4^J+N9caH)-=4(<
)79\UKFJ.YZL+JPOQ>W30;(8L\^f?G6F?D=T0J4+_1PYCZOEWQ;,XHIcY)eU:<V9
<]TNEK-]@=cKC1Cg@1/9N_-9[N#5]PA(Q4ePN1B6PTKKcUAa1)GNZ7P__H0dFS4Z
L#Y(B_1^Y)QL^EL2H]0b0W?1#,6b.a6WS]WeM;8e;A6]\Ka0=1.YS])3@4d(AE-/
e;IC/#(OcBf4fR[D#7F\c.MZaPQY^240))aVSO[ALIXEB4UEYM;-R,:4]O0aaL>-
,^f9,.IL-B0]7FNZRBbef.9O3>JFcae)##R-2.b(J]8B-M1KI^dE(F#1/JTbf6QD
G^&7C-ZgZ2P66+T1)SH^5IN<C0/aOZWVG^D>B>ZFG5]#,+9E=[]-D/81=?UAT4X7
&5>#LLEf2>Vc7Q4:0]+SBN):-W;_[L3/1SF:530BIU7_\<60]/-3&4X5<EZCG](T
X.&5@DM(IYMHV=J7@0A1TE:]SX=MY\TV#\1dL^?^g6BN9)@R;&f0Q#&@VN9]F4[]
,_OcTSAC#JP7)B6U;&KN0D-Ua:^XC[d3)7>RFc0J<-Z_Mb6^_K8-(-/8E3@S\+U)
;OM(,P02:I#-g5e^(5eg[WKB=J5aLLN>3;VLM/=+Xd-bX_U8dQAf(RTUJf@;dI1:
dJ75??8Ee-H\ARR\4M&OW.<\30RTA\B>@d;fAb/C/_@FMaW>)a^4(,SVEc:BQEW2
bXT)Z(N,\Y?2Of_,9MfU0V\A+/>AQ.a1F5?RfWf511-#,FE-,8^^O(JXID+DZU]e
Hc]ec]+:d#++S?4\,H5JZd6SP_[F638;.;1b1cF;P2D=QS50cRO#A0@WT+(-WQbf
bd_M?I49I_gX=;BVQE0NUTUK6-B/fgVLEX@QGI#3\\JZ.E>Ne@-=8K5G\6>AV^SI
.CBE7;P+UI7JFDg7Sg^3:g_)T^[IL@f#[Dd#+\GI<(MU/8SeAc)8<OO7f(\Q,2)9
P4GCSU?I^3IeKZ\b#>AEJ>UADD;AWTPEFDO>N1<I;g973G1&dC@@dBa@3M-TaOd-
>HHI+N?>fYdBD;Z/Z)2V.,<Tc0,CUD6=O;GE72gUEOHPNU\cN)N#EH0(B]8WTJ@c
,+7G2;_=dZ\O[1;&1A3CaC3NfT+8\1E.&@g5Dg4U^?d6#?:d]f<HG269>6<?9f/3
-L2cX__VB?HD\=_7EG8+FGM]DF035P?a>^6N-\F5CA/RMdI,c8CB#Fe:45W6/[Pa
ZL>A46I]OQ16e21AF=4LC=_\Y+b<baTP>aGVM^S7dP;.Z^IK+<fQWIL<S:UNQ:GJ
@^G6B0D(QZ\?K#@BG(S\=BOH8^HJGD)-NbeN-P\F?4,,ADQ#cU^bg#7g,:2D&##<
P2/2U9\<@ZO)MC<aea>KG5aVH-NS]DZ@&SP2I0+IY]+\(8ACT+eH?<3_<0A,=T5Y
5L^^:240^NE=W#.,XO?<PH0W>dAT#3gRI;.9)8WFX.LA<<F6e1:(1/c6+#F:8K>c
dEK9IdgXN2f]P;6EZ+KX[cIT,8/NT[5\QVEW)gHF?U#Cdg#ZgN0?8d;FM:FRgW&>
-\CGe#VO]EB?e(/-<N.M49=dL[LL,.XWZb[K63(3>3O7Z7+1D->WED,8^TS+ZCCC
RcAd<293S#Bf/[ZDQ2,.KM#0:dS0-?D\9W?.gOY8QG6bN7cRS7V2)-NU_+S6^B&4
4)P-:SLW-?]HdT6aH@CL\),eYG0QPE-Cb=/:A[9@HbLabS8YHf[Dg-W/4]RYB/Y#
(If]f(M=2/]#g\CS2=Y]<27E;5YeG:B_PM]AaX)&4\NYQTEUd;HE,Y&bB2CNd[;:
5AF]3;c.PLYUfRW,H]E(a#9Q0S[OMC&IKISO[gL&1K^OM]HLN0DgV8I/E<&#O@7X
?Mf^8,LH\220TP:8EH?3e1f.34@@E(._-b&P^Z-XBU;9,(+M7D2Y5VFCb-Q0I1E?
XFVYG>XV.R+(7JGJUCZ#@PN?;=)P.+6fD/1c:Z91GP]-gZ/RLFJHJ)2eSFJ7NHPP
BbJEeLYHVV61Tc/NWEa=?b4Y+55WM0(2A#fC4_(_&,5XG)U/3Oc1XGF/4a&BdKT\
3SQ-\9Q.1P23G6RINb[L.#/)a/<B-_cQ=H\>9]P5>G=@E6I.G_C&bDV=WH1W\[_S
Z1J&QBAA\E=&^Q0V;cVg\a+I6OYW.L19H#FI3D#_:92OF@DWUJBRb&?2ZXEbJb-Y
^gNR7A8H?-_YP=<dH_3DA>Q)g+OS+\DaQBf9<LZ?9AGK>XaQNGR=&aA\I,YD78ZQ
LT4G:fIL-/d7Ca]?@MH+@Hg<:O^/LX/KVV(PUG<U5DcbKZ#f.JJgGf?5PILH\7@I
PI.b1:]8Iacf;1AKDK(N+g-=g^+8SfZF)S17P,ZC]>S6ORU]a=BESI[A)G(O=aeK
1Ld5[8#51L+(R3[:P<N92PD@d(c/NbI=/QUWO?\0@KN0)C&1JBQZCBL&[Sf+W(U8
T::4(Y5XVS(Bd16##fFNXT_[<&6=1GLWD1&6R>^)HR_J25DHE=R&:A5>PECd?KTJ
H70H=,[a(SQAF-0,FQgJPSAF+<9gg\P]?)U.2dc58d[A[&d=6\ed]a]/.^IVQL;>
-&[,eU@U4I2B@-W-d;[4X3(3PAXCAe-VTTHc5<YF/Kg8+-dR?3_&6R4W/3?O6F5Z
gVFY74.TRYJ5OO@C24IUM;?\W(Q_KU,1EX&UX7+5,gc7NLGJbR\^.<N<+73&;(,J
<FCO;UD;RSbC<?MBWY&.?WDJ;D&O&96&NX(A[E=H-eFSd9+f0=]?bU>K9\?V/.Ug
Mb@ZRF\.P<-#2@G^H:]&.O+65OaEf1Z,FN(gEK3GQ=>,.72NYXT_FB&?WgKI?<C:
LN?_40H<58Q;WS^QK3&E\bV.g&W^/GB_E]@WJF(]NggD1O&1QfJ-A4g3XSUcBV5d
L>\e:KI;U6P#=5A66BRD=S>2ga8)HRK?2g:(bLG=OOLNRA9eF(&;Bb)-WUN\&dOK
.CK,8,gK5MF3_Ae[L^L..6#Gg+BO0gIc]+AGRe4N2Za#5DPO4#Qe,<.1A];?H,0_
d9[@;V1\5/eB;TdB?PWccPP6c)WABaU7e]WZCTA3gHH._1X\bR\-\98.EQ,1ZObD
Y=XWf3Y>a^9C.E?Y_cA,AH6-RF]BA@K<GAKb:=4]TL:3]d,EZ?MR-H8]Ea^+XB@5
[#3JL?b5+&ab&:Md;D3S=;HAgJ<?W,YEd.D0THaS3?1?RRG;2.36G\UMcKM/3,CN
/_O#&J=)9>:[+QEcF(gE-3WB1[C5=;:EK/BDMc[f7dJd>][GD6K.c4>-^)FR)N42
T/?5a5=b\U+2X22:Od5:=L1)Vf#9MV1WF3-UT8G-\NFgVe>Q0db/CCNeE@)G&RO1
GUL/T^>K@cd&AS9^GJMT<47QAB_1d?8:O7KL>R@f#5W=ZAXX>/YN3#?Ta>6aC^+O
3cY_/MI_#MIA&V[cdLWJP4/O6J@;)AGP/OUUC<K=G8A;=/HgZJKL+Ld(aBg)#^4^
6?Qc8>9,6M0\M<\7Y)W76>a<T_A7R;Kf?)]86Y).Qg+HGT=MRMV_NDZe.Sd;Q^@<
=J6O&e2=5LOM)=^@:7JL0Mc:40.,LT(VgTE>GT29d@I@/NEB1EeKJ0g.44dLVB/J
/PHD5<#TU[W20_dag19;;>+7AWUU5UHc7\Kd\8M&2ZY]\E]\1FU#<A9&ZK>g[F36
[CP1c^C>c,C4a2/Z<92QSEf^,1_A2U,5(+LLYF:MELfaN-Z^+b;#=[=033.G-?P\
a@gJ=G_XA<L1a#U43,)8SU;^8-W&cP^+Q8IFO]Pf+S;86.WS9T&;3&LZ]4NfH(A1
/X5D>=L]C&YG+Y5G;)_Xd_7Cd@<B\2KL0_Y)U,IZ<=ERV?Z2=^,KfcO6WJNJ[?:C
_.;ATF?:2FJ/QQgF.SBZ6Z7I,5-;U6U>KIKOSQJ?K,VPVX]O1RS&AK#^A#5(_[OH
&d)-16G:a73;-&;,=NWM8XEE/@^ET4+eTR,,Scf=7ee[3DfS(CL3+A>NRZ(+90Q.
N?(2O5K7.;gLbT\O2eN6-53=@MGaSHD5._^6GZ[ONDdAYZ+ZU?(e),D(9d?+Hb3D
5H<M:D:MCIgD6SQUG]>U9H,OUP3=\0g]]/FTYHR&MCYL:9LE<\(2\F27/(cURBX,
&5TOV-eXf28=<_?G1,,,&;->,VaA<4Y7=;LNT3>^T/PX6F=:QH@I5d_JL8PQBe@A
DCcf&B.)([^KYFH6Z_0&CWcd#VSIa+1+Jb4d&<dMV[VA&;6@gVWM8?c_S409_HPH
><BCIKY;7c085+T^f9V9HT5TUDR7&+CdP[33N1J;2=MGDLPW?>)KH+YbZJ[R.eDG
IQZW<7<B=1<-F)dZ&G>3E:3KBADS@eU0\?91fd^4KKg.>4WM)JV;1_J,<=/.NG<W
@M\L<=KF655JG^]UWb5>;<BO<.86G?FB./)7F<ebHKK#5PY..DAV+/fU@ECeJ+XQ
WDLYQ18-W(.]G;VR1FEc&F>_-SO3IcD=HZ_QD5G9PU(a.?J:M29RI8R\G_9#,gLB
g>4EC^GMK,_cdeX_?F<8P6^-T&6:-92W>de:17/?V)8-H3KJ=\?,[/7XXUU>.?.L
V,V)Ca#U#_9I-MC1TK_P0^_N/.1#F>Fb#PI;Q]dDS1_D#H+a@KVFVF#I<5##IGLI
./9]ea[8]+?_O6D?#]G,ZS:8G9\9VaEK=gABe](cD(T#A;-WOEHaT9.G;A_Z?:7.
MWXd&#LQCE;4THT<S,N_P_dZdY1bITDf<X?BBK6CA?Q/cBSZT,bNIc/Nf5_/aYgY
Z?N9#;Z^></a?c^<2&5<@SQIB]L59F,];/-:gDSF#C+YRPYC<6UI5fd;K2J&G_&2
]-AX6J;cfRSaOOI\M-95cBDaG^\Re)69IHEUe6)Bc;<6d5L)&7WgdS)0>)=-DADH
AF;=NIcW2\9/eYa7]CK/QS_)KHI(bAEU,1[A0a/=.gPUF+a+P02D55:fQ)^Gc+@[
[FM3QP_MEN-6UJaa4J/#.&aA8TU@c66VF,\ZTZ(O57?<.&OXR>7;,Z6<=TI&1DI,
/92T>4S5YgIV6D6fE1Yd)V>1LVa(Fa(.)]Ae/F@]U4P<S8,ZVXd60H^fb;(WA,/.
-g)F^(a&g#cHQbFZRS;Y\e_J0]W4J9BMX)T4:#?V/4UP.&FO)R]3U[.=<a(SO^W0
+a\?+XZKYDZDaRTd(8O1)Y9QZ@TNXW@8d?6H6&)J_YLX1W4VEWg\>-C0IG:.\BD2
XGY_4LJJX<4f1Ff1EJI@-#L&KGUML/#&GfbM>F8QA_/a#AdASVQZ+_6F5_:YZ2[Z
;cU9<I@G=Q.\EGfA08Y4?aU1f6=9,OOM6WHZF[W,5BSDF/bd+=A=K.L(==4V@:@a
;g(\Cgeb>d?QKS^UL/#DE7//JKT&<c:PS(S6J43Pg/OBLTB57.09E^=;K1eN2<;;
L(:_/[,d?3_)g>7.eUF>;W/XZ[LSDF2b8N_V3/1Q=-JL3eeI5F^CI#GLBGYeBaAN
+XX-F/;g^\1<4D<UUFb.)13cM?S)B0DP:WBD]=@JL46F\\AeU++:BfH1S9/2V49S
4)5.6fUa_E([L^<+;GBa(G?>L/C&9UO\=R<5Q]9^VgOe)[>;#P2TF1dBGYV54<B/
PE2EE4+ZB+ba/09FNGEK1EQ/OQ5g[J=T<E)0]I(WT0G8H[3(K2bCL-6@gGbR@\D)
1JJ/a<S85>12<ef0JSB^ZAG29c,E&SU-QUD1e)TET9RB8SZYCU+A)5(b5(@W1:X4
&MUfM&;9F)FHRLK])L0#QVU)7^0(+VY<9Z](a1^>&dV7MX-@L7T?+,YQ/.6TQc>f
4dJ7g2ZXUG_1Qd>:MG/WG)g<Ccb;E]bC6RF0(0W#@(:W_EX.b/fb]##g:<CKJgRZ
118PdGe5bYM9Y1#RB]YdHHZDZK<XB#FD+X[FX]\,B+<.Z=[C-++JG0<Y(H5Re/2G
(>^.ZS4#=d6SFM;V4T<\DbR-&)b[RQC?N<^^NA[,8V.P^ZfLX8>c>SR)K1Y]a?fJ
\J+KUXO<1)E;3Ge.-EY@/<5=Q-d5]/Z&c)-=Z4F394K-?\.M&d)4WDHRQLB9W<#-
fI7&MZD8)FZ?+?D^4J(@^MIG+;.RDdY&Kc532NC@T<,6Hf_(:[AbKD[YDD,K)4\6
\]f<V^?][TBW1ODA\K?][;d#_g8I8Gdd?6)09X]=37B1?-):X_Y;Z?,A#)L0)LRL
e.S@)fCCY6>A&DFFb[_aK<LLZ_gN#G\U(FL)RC(O#QT\#6Y@b;5(><1+.Q\^QNS,
[4A4ZV9<ebWb.V#;/#+&ef(eX)g^L8W9J8Z-#Af@?eD+QgD9<GG7;FNEEK1[D=]S
HFQ318X4ecXbXbWY&/f7:P5UG(HTD9eJ^M?4]DdM[ALF4XgfO.[4T0F.P4(QS62Q
QQ;&SM,R;VMY0/ReEFe)7DBUU(@^9fN;>??dS3Q_2f@,E,P8eRU931AN,g5=-+AJ
6+RL7K=-EW6_[P#KSfX?9@]EI@GL:@9@13B)>0-UdP+L&aMf,M(,)>M.VPHRKC_f
F)^MYb\FKP?4S@2V^aV[4JcV#He29EDHP/&6XR9FQ2#dD7VR<+L)g)IZ_S,:0;JX
BDSJ20Lc>RGW6CFZ37YHP\WF_2F-4D-^U<3WcJLPHa?e58@.EB2eC<cedR9LXK,8
OTN^e<Z2W(:3G5K>ZM=0KfFW#J\@BfCR.4BGg5\Y-GCZA\FMYR\\I5SX:88\1/<c
ce>8F,?46\Z@DTE64+20,Sc@RM]>4]_T@(HBA#dKW2<5U4AUe,K<LV8af-:A5JQJ
b@<:^C&C@.X&((589IBO>Z;K\J/+EDM<P7?JZ@DRV&eSc^Qf^?BE#K60#-U<f:QH
5=K?@a,2H-=^X7XcV[f#M[/#X04=TV5^Z75W>+N;RCU:2EW-(Y[?9]-U/Z2KPIg(
Ed?A?Afe87c<-e7[OV[[]3.V(\1O+V?6Ng)aLX4U@PZXR?COE,6QPMW9,@d10@S;
=,Df9W.<R8]^>XT7.OY:?46):?.4Qg9?d6I)KcD;R)62Qe(VW-df4J/(?.3A2J31
R@PR?,[^K#=4&2ZU2_)S:RT+Se1;Wg#P\@K\KfY0-MYP6X:b?\G6:_,8_#Z\ZBe@
3\g>C7K+J,8UIcg0(bL2X6SfWZ5;HNQPV72Z#9CHY@]0bBcRVAc@0C<E=F>T.?X:
@,:_@edPe#2eaH?9IV\2Zb:[NF#?.c<OXXRC(@.854.TNNNY5V.X^R+GaS/3??aa
&4>:)>3R?8WJ;^M.fIH@&T7?1/I/ZJ/08c9X7(4M?8,Xc<@cM].OV.:aHPXV9I=Q
KX,b9O)/6BdQ[H=>P^TP2TEHbIN)\6gRHcI.gXc8]4EJS](G\U#6:f8bBfH]6JOM
T0d;f=Q8CI]:RPgG6NfZb^KYBK4E/V:G-c;C<1<gc65eAbJ+=Z.\8eQG5#fLf<Z_
0NISM1@=\X&RTSH?8:BJL[UWI:JTH[0(bY<1#D0Be&+?X[AH=AQNS)IT,EK>b\3O
QRcBf^\Z07BfdHc>Q0HET0/5F8C0WN]8QVH4dI1TP;><WI,dc07d0@b_A-/:&+S0
DP3I++I6IIXT]LE/MH6(3gISYX9)4S15G+]+dVB3c<FUA@dDFO=[N-_a1)@d?e2-
>a,2c0C;(b(a9RB4KcLTfD[/LQ8^9[\9;0<]\?15;.8DW^&Gdb6<D]#3=VdXE@97
VZO-7^7CS4LF8GT&df?^+KQD;+87gKe:Fb+_/#WJ&]?JYL2>+W),#QXbdc<L<I@Z
B/&^,B\+SQ]O4&b9a/UE+XZOK>BCMZ?W;?e@B2:Qe9LPF[^C-^C<L[\JE3,VgC8<
0>@4BJ<Sb923XC[[:[C2TWH^K08:X-+f:]K<2YAScZ@dENf,ZK@?gO0GOd_2F5YR
:F_3H7R/7<4PG5-LJ6RZ6L8-<FFLG.[->M9aaPD:(;P,A:6,\#.3,7gBZO@6B3PE
fd7?KE9<\</LB_3&@f94e4H[@,d\29]D+Gc&/Hf4#&E@V^Q7I_d5(cbHD8E?UI\C
gBMC?E:6?@3SSC^H8,LY.X&e8UeR-dTNfWf=U3>Fg-d2W,-@EY]RN/MU#SX8N429
1O8S7Y^QSKfVcT6WGeb(6CZJZ#SC/OLU8M4PRZIgFI^H\Q0##cRedfVb[W.bFAKZ
\=[4K7JE6a^d7L#R@Db95L.eUf@gWX5FJ&W#cS2JO_>gVgX#[_)TVH_@DP[YQgVb
+2G:(L#B&.D([deggT)6b7T.J./2,2<@[[/GJ7EFc;OC?[;08<?OG=X2T]N8U3B=
dEI48E&=aN-/8d5O)Q_Z)D4<[(5]+M>,0KI2NA&[7_]E^=fYe9[(00JG/Z(8EV6/
gGDRGG)4((KZL.XEFgRDUV+X\BJ-WH4EKIf/[:P]OFfLdKb^QS]c&K/H9W_P\?4Q
;G#@.VJ9_aNZ#e&SF;Q:O[Qb1=UeP:aTbY[NA<cZ@F_4<I\1@W?V\Z&eJ94K/MYO
/)>Sg-XYUVb6#DIAeYfa.g8R^0/&H27I]#[=d3QA+fFJM.OBIXP_;7IMSDMRG>WU
QJ85_LJS,=Jf5LPD/)3EJZc[NZL@3ILL(5B0HVJc^U.#Hgb<(^dI6P+)9ESHB[><
f^bVQ3RISW1Ke3=C0V^>UKF&HK1IQgV#eNEYCS+3AKS.NOe29((.7aEa:#e#<c[f
9&1JD3Q3_WF3>[YRc7J_9K^4A4D^+VNKK?:Y40[-+X<=3&1#0276e;H6M1O3@BQ>
8Y@0f^9Nc&9cbJ2\LE3W@)N4J@JMaU,G;dgCWRY;X6E+9I:7NFJQCa@fIH\)WMTS
dScYZ:QVOc4N^\aPO70DYeaAN^UBa7O+FBQfRfCd1(IIH#U.;7VFR_0KGX)OLd:&
^bU,7b-+IP/acF8^H7gT>,D(Z)eVZ\HJ3E046OS6gZJINBW+YT;de]?ad0#5D.N1
K#-AX=-G0aNN8JM+=I,YR6B5M-BB.^WUY^KVCJDH2?@J2US61[gM#Hg-]T\JcW+2
G.Y^>5ZVA=#&40:V3V5F/&WQ#5gT8)7@]XB(K]=b#@Ke2MTG;A_ONUQ2\WJB#JIB
;Ca51=6E505gY5D+]fV+WE+F(^@J2[@d7?L>g<[</TS82O\&6&2C\HbKO&>)/D,(
A(@=1LDT5\IAeF9.Q<KXJWHD^193)>e:;N8&T4CTZO6):cS]cX,-?TIBNXfE?c^K
AMP>#LG)Lb-]J0T_<M8@7(&,fD6<Ye2fC]ZfA(gc/4dR([73-H-DQ3GK]/A?Xd?O
EJUH9.D55JIX-7e@EC0=f>PZR->JS_0[OUV.)1?fYF7O9d-FD8[#@daZH)AU?]gY
?PgacB((5L7B&30MKF:,&(_Z>Nb9FA5U]44A82^VN=#]dQ:9Z6)X<g>LO10^X]g_
9Hd6TQ];a\agT]_Z)d]S]FM\MgYdbX,CS2]K]:CQS->DR)_QYZM-(2\+;3eaL)+E
JGV]N4e6J5eAUQJfGDG0>BTd9b;9?/d>08AK(A?DE1OfS_E.VLDP2JS.GH14cDgK
AO)gHCI0g_\KaC;L#<9N,/_c(3#B0cMN/19\4DZC?S#ZV686(CQTE9eAZWM,SdBe
1bGD;0ZaEDCK2P(<AZTMcRVWL]6W7>EN62\f0g49YSgb.3W_H9J&.5[NE62D66E.
(aTbX2HJY6;/@GFM_NV:64H54aH+1E:TeQE/FeGWHH9R:0DFI@/a8:=dbdZNROT_
<04AM?-d00d2@K@_B?:TGc_0+](29V[19Bg06-MbFEBbdQdB7]?.4&?\3@CCab?g
f=af0]gG<6FW?93COEX.J2H@,^\.GU+5#=-4#A-_4YKM?#.M-NeJN)]JPT2-P40V
=^?ANJL<PSGI_FZfIB_0dTL?I4H3[)K-KNALSa#DYE,(Q>ga39fCeP9gD#MPWSD]
+E/MF^BfHU0HS9\2e##-eGB)d(1aEH-SFZ+?-)Rc&JA3J>5RKE^<g3#;L/FWD#GW
?OcEbZQ,2@6PHFNRMW4ZG7RF;,H[AL6?<(@f/?f@c6N^aUE:\H\GdPJ&Z^Bf3<CX
#dP-aBbY,,ZS/DV:LOJTZd]RM,:,+dG>@MOd0Td4AXL]KNQAEgW/R7.F_6WCTAP0
/K(C8+&=VNX]GY:>\b67K]R,fUG:PHG(6UcI.][O(QR.E,2B8Q)@WU3YM3[A)4Ff
,D8>CXZQebd6DV=PS>&TBS_?I?a]ePGYOGI&<KA]d26g,/.:Ea3MGBaOP#B^1>(5
dbd:<LeHf]C4(ReFX76G3#3S;V5R7=VYf?)9G9R)f7XH9.8Uec9fQ1GC;GX8EU(#
fg^J[RT?3,[7_=Sd-#C@W3Z6.f2YEV#gP+bY]c<Sg0>da4XJg9F>OF(MVgR=?F<)
=;@C2R,4GQ4K:@e?&5<5bg2=Pgf(a&O-&+SGX@MRC+PVBO&=]9I<LOI;e?<^g1e+
MP#RF:,_gVE,WaF[Xf1BH27>NR/cGMeac_],1-+J</0X.6<MQC1.8,];cY)\8R1K
6;\Kf.BHDX/PYY<C&58^.AfE50#(aF1880ST(V+0FKE[,+_75L=\6R#-1.cUR\R>
H;LMMI_IQT2bTX\IaaOFPXQM,X_LeG(G@=,_-Ge<f7QA>/[]),J^d/aI4gHgDGPD
#^<R3_K&L[0I]F/+3NM0NP:#HaHA.[0f,Wa&P2f6N<>+U7TF;+M62<W,\L]_NDWS
E8I.&@MLD[d-H9L98/>ICM&GbZb4TT^a:YTH&Q^Y,B-J.KY?U1M&X.b5&C59TbTY
#d?#I<TQg:H0A=ONL-8N\Y^J<V2e4\1Y3>:B;&<?:VTRbMH2@EU20>[RQE+JW+Z)
LZ+JV4FgKACFHHM#TVE9@0)H^cG5ggBa.A)8@#C4RCIP?_AO#,4daYbXC(<;A7RL
\MKS,Z9,_e,5RC\@=@aa&Ffb4?b]=H3QJ41-MLf=35VJ7HB@4M)eQB7gU]STfU>)
J4=L/Q\8L1;#IYXgO)L9aK>43\NLN]\a8&_Y9(0I=_d>Q>A&J=+WQ;KD(?5,?E\B
NafCF:?-bY&UXK0-cR:53cD\NL+NbP)Y.>AM702>&.H\Z,I3>HY7cW\PPUcC<4.]
7.GAMBB]Ya<e+</g+8W&g2Xb_2;FGfLP@IJ;WQ;@Y=10T@Tb,)..N\<W7^)U?H0)
OYTRI[Q>HM1(3:@dYFD<.=CMHJA.,0[fdOeW36dMGPBa=MN-#&7V#9f^A71eI?I4
11Q6+9I\<YUVIFS:-]/A=gBa>1\KY=Z)/A5>NO#>T9NE2#0?K3L[/JK53^8G5HJ<
N-Ab&N9>gbN-(W.G(P4=;4QbHg6H#daTR50W:(FbFU<AgB86WCX:T_g8Q>0L=[PO
JI\LTN<=HD-3X>^g=fPGN7dU;+J+b-.[[&F<F4K(R>Q,R/9\KFDg5L,:#,7B7?;Q
JMfVE&W3.&^^:WE8:H,DF=;3IG7E3DOO\K5OQf[NdZb#FB_\O2-dZ\,#1NC2W?GO
NS&/N6[VWV/8cI8DG-<Q45Z+ObQX]SdPI>L\A>T#6K<[->G+#C0AY2P6A?/UJ3aX
;H+B=EGF&9LZW6+cV<:1_&gJf8GEML7X695VbRDS=J\Le48YUK,K::EA/=1A/09>
&(A,&U5#+L\>SRB7;7c7[5+FA</]bL5,28TW+_I<8V7WI].&:d\(=W(E@DcbI2S]
VST&>9>_\)I9[SY;WK@#+\c?UMR>KE@5IF+OTY6SBS64]33^+>aA_dIS<f7bb=#b
8]^1F=CV/2e60ME&Pe_GR=::0&F7RAG[f#(Y^[(AL/3RBV84LF7cg&SW,baB[&R6
?.U(IZDc&]:)CZL@B;82e.(0:9,e-E6;./[e.T@MG_AF8E^_=K.^&O5e7/^9+/XH
C=,7Qg=VOP.1#Zd&g6da=)BTEF^f9(N3_;M,<-H5S0<:eYW?_][/V4,BZIGW;J9L
WX3@-N8)]aa[&I([BeK_RB#IZ7>@-;f;^\P./\0@4LF)-CP9M^JfVSA&6[/_Z<ZR
7.&I,#+@=E<5^&-OeNMc.ST>^HFe)\<(8W-02TQJOWa)ePaeIHT5M(]^L?Y?VHUT
gM2+bdAgE[FCL2G=F3fY)+4f:MZ@eXc8Bd2REF]MHa>>BeQR-\Yc5/P)b@^)3#c7
?>f@4M8=V2:CG5=O6R/DWIU3d?LBQPB;,453F=<\H3>I3R94=-@JWQ(M_8@YTE^:
(#+TS/#2Ec+=Yfc+599YZH\/>HM=f5Pc_=YD46TN]>U/V4J5CB/00D>^a:T_V=e)
A<;CW#[HDKg=+c[2D/Se^NCU:]Dg+GA08gF)US0OS2(CG&5AB\BgBA>#;1J#>^Ef
I:MUS5fY5GYAUD\(L#[,fW:dJ&4g#6=V\[=M=&cB\ZEY.0ZQ=\\&be-3:[\(ANUQ
6NQCU3@+?=,&b#g&?fI_L6J\>6?UY07EY0=Wf/Qd,SR1e:+c38^.I+2aEJE[[c7e
f?3.?Y>HASc<Tc8^&@0-M8_e1E7?D<60R/]1&33Aa#88R:FJFd60g&fSA+3Cf^<:
496Sef)C??]FAU75=e<d^YY5DD66^J1E42+LKfN,gdBaDFL74L+H01Cd<8H1>L/<
,#&dW]@6<BNZUDT5IXX__Z^>2;Y=<+Se)dVa=4gS]YDCCGd)JD)F(@P&S0&[S^4L
OJ.]7H=#J[e.=;4Y6c1QB,RP0GYS#/7L;TOS&c1T)74V8)0PMQT#a_G[XHA.37I/
NN,FC]-Q;ZTN/<_aDg5;IZ68[d[S@3)[1T&5&]@I=Ig#DNB#b?@>?_NV)B+\Bff7
LNYf8L:+35P8DZI&d[1/K,:DDXE8b+(M5>,G.;Q>(QF:Ma1##A]3,;GL6eG=HeUO
]:-J&-Y0T2Y)@DF:?baZ<H/L54:9[NAM#Y^_AC6].bK]10Y]M6FKDJgOd1=U9K\B
ZC9J<NGLOdEdX5T3VNG^J&LL2F96aKTaIR>15=L\2O4K+EUAH;+3ONA66e_^M:]7
GT?=9]XTVY<Rd(cW2Ig/4gF<[GeIB<V&(7@f]aaK[3B\4Ta?)+6e2NJ^?dPQ@HO-
4gGVcC2XTKR,bGa_@DGH<:9Y1&E(T+HO6E&]b0@7dI9FLAICO9:K-PTRPG8UDN3,
]1<7BEHJ@F7TL7a705GCbNLd61:_)YEQ(E,#L;JL,M)8[b(+Gf:CcaFW&dU0K0CP
BeX\\C.>a/^]YRTZ8H3)G&_ITVQKW_FY9e#YWRCSg0[A+gH5SUfgC;0.<A5-+<<J
)5?:FQ28ZSbUKH[\PgY6O2>HgOVQZSR.^F0_W#b<PVFa<BA.Z(V4:_PM[KE=Y9^,
F>XMZEG)3?PIQf4I_/PbAeWd?,_8/P[c+#>U,@QE)X=MKN9HQ0,,/QFNS?3A<>b5
-2IVF@[DS7.-9b)&94^CHQ=Ue27O;P&X96Z<fUT2ZbdNc@]JA4bYeXdT-)--=0@S
4/G74<?,4]56e+S<[#W5?F5X;9#KYFA4?<Z/(c#FPAb(:_B[g3W[bVO1XY^FaCPW
Z5;^FP8b+:S?PE:g^NE:ATg8T,I[J,gV[KU:MXEMXJ&FRY<S[+2b:Y(IMfT&>6fA
1)bF,YVBb4@.&-Ef2L\IEJD:[9LE@Y0XbSad06?SM4<J3A0gdC&3UR[<=Y=79NJ+
B\Hg^>95<C[0U1Ke-:M0&H46Zd=6CX#Y]_/]>XNX/(6-1R\Y81Y6Q7O1]D^6C<SL
@4f8J:=7C]4;BCfMLE+-YL/YOU\6IDDc?\R#HfNQ.C\-+ZIG4=J,CBW3;HC6IOF,
-2_;]E^cgg#_eV@<O.69BCWE=1S4M9[@O5<U<.4D<EgUA=6<G,P@@94^>3Ib>^3K
:8Y5Z=X?aGXQEA2cW(#eB4,(ac#F/fMHSO?4#0>e_aV+Z0(&]eL(NF[5baag&-3^
^2(ceF[1T@;^5FX786=b1Ga\>EN6EbFG=1WI^9<:Z+G<YDSYDfKY:ILB><.E::+R
5M/aS/fW&X1>04W(;T4:SY3#ggaMSECaZgJg:W8S;GcH=,Ab,7g(5V4QQFCV/B_/
Fd7dc2gS-?,0XB>>68b0<MTYR3)9W<.M/,&FgRB)ae,dc(Z,.;2HISR/S4H=;M_D
_Z0Dc/YP?.B6&NTFT\;JS&V8GZ(f?3X52BF8^CHAV:H9MS:Z^7XQB<<=1C4W(/fZ
0LC,O2.OH6gBM04ebF6BgDP&WV?H63F]gR0P+<(,\a?fM]eS894Q=<G(,81E>M>6
a/4[P_#,0RNV0bSRKcH]C&Y5d1/P).:KXS\/=KGV^Nee92)GaTd/0@X?acOI,@?f
+S\gB&9S=,;HZXUTJ@CH)?RC#YL++eRe&)QN;5&05CY,CaD,M+Td3\2CI3LIJBCY
KT>5;Jb[5.d2?\I<1:FEALL_>cOc\T\^V/4OeUGM9+Rc4.9B>D,.(6EWfI8:f[fW
7IYA&+#XO_e\:e[8dB:LX8I,VY7GF&O<C31R4Z>/fMf/4=c4a6Y[YC(Ab_[91eHQ
1.5QPa[eS7Ad.:M6M;8?X3fb4:AO(#@:]GED>U;5^87H_J#cdI-&]H9OC3@U[Bf+
],fF?WbL]5K:R39L_,c>]+PYC+YJfHV?7MZ]8PVW23^P(KQ&LO4b-XE:VIMW,UDD
@_CP:JKL)YY=a5Ia)/d5()1a(RQb(bSe<LHI1K];R=\;23fcHNK#4cV=&EAfD6WU
RL2]:;#fT^3;ZZGK0eB(dJ74KHURD,g\Kg:GMK5)4M8?&93JR8&@.c5A=(1J=\_f
(.-).KVOc<T&Re2>cfW&OQ2[Id<<.Wb5JF2ST^;_JV)U9-GZ]89e,^2>+bHaO1AN
Id[,bbZ(gU@KKH>T.I122[/NTYa&IIKH48aRcZB?/FOee>IUMJ,.a@OE1<6gdGFf
4ITO>+?-+YDN7R1^c;N?S^b^&NI#RK.EQH@;K_V6PG_e6>@5Sc:+6a\T83_)YDMb
.W8)Z-d^9;]R+17O.:FE-f?J(_4C<X,_[g3?.&(66A\&6YO-?V)E>(:NEAH]:;YA
Q._f9(:Zd8L>Z6cC:X\^]-M/HENH.U,5DK)_/AYdB?3F0UQ0cb/0\Ic@62?>BO(Y
]D9/UVd9_UHER\6@-8#^OEOQ11SH\VIZ\e077X>3C=)U2.8P/^FTZ-7@F=V-^V7E
(C]L3+Gf?g48AYfK7V8:>@7[>NGBXW@72^3J\]97:FL]&-&L76]KSR)g:H@E>-.F
5gQ,BcOI7D(Y1YMT]W<5<dT[X?_E>,L)?L58#R_+-HAc:bW3a)\:+.1H9e&Fe2P<
eSYC9)d[(5\XZFO8;WK):;\OL>/Q22fF0M2\]H2E38TR\><Z9VG7C_L1\3#1=:37
=df2>QRg8GBOdG0:E\DbFJeG?g348c_@1;FE9BXa6\eb\C4#.=,]?P8UTb(W3.S2
F=C.:7Nef1]5B?J/L4YfP]LO0RB:4OYML2@^ONAaM>_QXLVR@/1CcV58dC4f36H_
(KB5J=\9HA+E12\KE\g-=d,)FN1WK.We_;ZGeHE9^^_Te&D&&B>]\ZJBUWLf]egE
1P_6+U666+?a8)I>CGY[?SX&gg(=.D\;NBcgYa#<g(f+FYXA&])b4M4IfZEUb0-8
KA(9,[CCd=CV&beMUB)_QgfV\\QBTTWa<[)W=f&MY73A]U:gM+e?8?Q__,FZ;VZ>
;0,:E@1QN]\L189<-HCI,TRAZ.>Y?WZ@L\c7SHMeV[H#e14Y>NOM=]eI0X=ZSa0_
PS#&4Xaf9]gBD/Vg:MT;+F26?eD6+@>USZPRG8^XFL;JRd(J+S.DC+OHT1aVP-2E
&3\-gK>8K=;6-]V\O3/;b<7&#,9]W(^aZB#SWQ<)8>WZ-2./92YD]Y(1R:@L\R9P
G5-d9H8UMR)S>3R./fZ;RTLJ[7TC)S[7=N.;a\,A-KSc102dN&F;H1LJ5X8[b3fg
JBR40\cN?;]NJZ_3-?e+:L4M-CK<\)6Q:._&3E7Y72g@dYbZX@U;\gM)O(2<0=Ge
_KG(5^-MK9/],IFcfcRN7TV7W4d^dHR[-W@#XW8/c:;4LM:c(_@B\MN;PLWJW(Pc
-U6d<,U5H.XU;60-X3#,SA=\,3HIfBVPM441c7LVW>4^3_LOb,e1g7bW^J3Mb<Uc
AWW#RU^.EY9]cRNC->/68LDBe^HG=GgMF--<f=S.f-:/]T9YHA()CQ62eCV:XUC)
,#&;;4b5^>DZ-C7<Q;84LYNfa=P[/C,_:+EAV:;,44T[_R3C,YT#M:bS\7UEU[_d
CON>f1\Re-0E]0S=C@^0)TeQTO?/8;Y&gY;D>c:QEOWT_4F)J?Q3RWRaUfI[W8J+
@?16V9LP36J<B7b,1>PO79b&HcVHe0;18BIeJ]2,3VIDHWf&F9M<7T/R:c02W+.1
1(bGGRGBI@44QJ)M0B?:=]>2A\XZE1LHF>W]9SJ(Jec8T64@Dc#S;gO5=#@IJ1:C
dSFY_1MVGf+eR5)6gU&fMP<S^cSdH^3P(1fN=E^KD.A5O?@+7NVeFJSF,.fdc@T?
0G14/Y8Y(cN+OfC>L>=PD?Pc#[7dc[f5L-IY0<CfJ[(3A+?GCS#f#4&:P.F<3>8.
2V+;8c75PD4,b\C2+c2Re38[3)X&B@?f7R<]KYcU1_=I:[LQfI\3<aZH83:>DIKG
[e+c2(4Q8,<YcJ39+MHCV:\dGV\9N?FYEY(MdF\>0\E6PXQ3e1@af,<TVG\<U\RQ
[E__TAP]15<W[&@=Z.?g)66AD]^?^--(Kf\(3G@)YfKLAJDW3_:N2:2ag;F5;F-.
Z#SXL=5U8HH>_T+28d=e#;/CgPC5G\?F9VO]#@d@<We5LQU>=APMULHIFTNLSMaF
Qa2@STW9g1+PRAAIQ,@5MWUYgLb9Tcf8M&YKSg=R<[FJA@=ZdI?:CTCHT<^K=O&<
36CK7;MAcX&OB75J+_I?T.a9TJ:2F(_K52I>77CI(XQ-8I;#I&8.K.0VAdUc/NU8
3\;K5F\A.dT:+QVL0HF>Y4aNe:AF5C-#BW=#>X:PIM_B@)WXV/81G9[bZ)S8+3c1
23L2a>3VK9S;:K4@RXN&Xe&SI-6f(5Ce-3I]2JH,.:T5>3G>L0;25[[[6Y@-,IRb
B/&+HfU6d_A3NWLBF,H78>dR?0Z\-d/f#:^QgM#=QO(Y8VV=&@2FOY<1U/g:M/:1
=&V,bOLYLJ>?G^c,52,f;OfPQebBCWK8^(97MCE=P4a9WYOZ2:=H.7T/RM)-\CAd
[)DGNX_6(THd>\#\a1(8]XU/dCUEK0eGF@Df?=cgVPJ[&&=(R0XODP7e/c=5)2^7
fa_FbST@bO=.NCXP?3;M:g,\=ZS,?Vb+g,c\)G;I9Mg04UU/MOMe:#d[20L1d44]
HV_7:(CFBI8a@:e<>dcOb:9FWd[@OY/J3#GCZegd,72+HcQO\3>-QP,=Y=I0E:S8
-:93K6f<(S+Cd83ggW7HZB4:DcIJDG6YCWELGcfBF5Y/<C_(80&2S@-L_,<bK]=@
Z3,;ZHKH0+GCXI1g&HQbbVCZTeZV3Q68R2SW>3)64J0GIcY@.ACRW[O]<.f3?E^.
>:NU93^Wfbd[40Xc85)0XDI&,E6c#d]+3VeS7G>BEM3:g3XTG;:#WVf^4/8M;<da
E;@^WQCVeYF_0WG;fV>23.QSJUe+:1E4(PA6cMN2f(SSH8^7OBENQ6N#8+6]Gag+
6>&Uef]:b#gIY<P4Z0DHaKS6D(:5Nb2&NR^gE1dU^Y@1VU>30f9.X\dg=4+QC6PH
2Q?cXPOH-&V7FUIAESF84\c?MK:S,V#:_&YLeIT483#B:FDDXVJO8;W7/@24f,_E
;=RS<I[5b)g#5GTYB)8]53R3A)J@X4Q5=d&TGaVR0(gab9-]76:N5Rb1JQZ].7P#
[\A>>U[3E#N/J-W-@#\S#)^-56gKTJK?7(U4Z#U\Q\A;?&/U8\g9_J1fPA<)WGS4
B7,[\bP0]\-J]a(&_:__Pf,5/?(>daR?7Q4F\ANRXa2?d,/IOL[5d#D,^+@XX0[;
>+1cfcE_a5cY,F-/TNJ]cL4=452&#<BB?:AP\7FB81HbCN6FXV^W8#LX3P?E.CC,
?/C/X(EdG\&6=XCCR&4_;0D?[)HFg==@).dV^(F[UH\D<JT6Yf-f_F1;#.Ba]^fY
RN7=P_.3V[]LWVTG(I3D;\Y>aR.G4#S8K#U;gC4NPQU_V>XZ1gV8;MW3CW98A//J
f73FWBZX7=0^?6?1<@5,<=07b^[:A2J;_SAM:R@N?3bd<aM,9F]fgQ3BIB[/<ZM/
gDD-.Sf/R?-C1&EM5+S>>&(gI]<^9&;,<4&MI;J5^R32O891dID)M>CUYU/d\Cb8
6be9.e_[/gBUH4T4_\]EZ6&+5-UG,DPEX?J[cIc:ed[OgT>ag6<WgA(W4[D[+L]A
6EFIfBR^/a\()^LA#gg+g7(W1bTC-HeQ)&=[4UKT94=6:gZ9-[;))C-]F/d<_WPK
R?(SB+3Q/[PO_TG1]O+J4A6JPg&76cZ6HL2SD>VcaWRB11T>&]?CP2_2^386#VBd
([B/>&7?&VBD#;fI)U)RgKNMDeLH0F/d72+BAGWSO]GWJ9K3;OQ=114)Z0W>:c38
;8/.:]A]SNY7-LZNcB,)#<,Z=#X/@0/.L7IJO?bX8C5,4fe06OFXBWWL)XCUH/1\
YK49WFdEL#[V&^V(=d[M#VRRd;WOg.T-fRJIg54B.c1KXNAXI&VL72gMQVL,U,QZ
d<8[IH:K+7+JOFKIf/&Q&#K#D)f6-QF3388G+ZE.5IM.4,gS:aE\J+VJRIOc\AXg
YHA9#\4MHXG.I<R7]5QR]/_78.P]P5C2Y#]@ZS7Me@Y78fZ]=#)[/UX-AD3;Q(:3
fTf-S)16/P,3g1>^c.\8(03KT\&\N9-gC\707WN/XI_#R<][M,6[IA^7?&aX8<B7
;c9eMZ;MCZ\P3@FO7@f9?Ha7E27<f8;Z3QG@/>I-XV?0<]VC@,gFCY.b099=(==b
G<]V@[fK0BOHf;FM0S0JT6MeZJ9-=UO/eH[#:T5AgU4#7f6[J,,c2Y#U?4O-E+Hf
W;>>6(Dc8,;=X\(G9Sc?1F(eD?5fd1^>fB;aLGFXP0CUcQOFb^e]C??2M9AfQMPO
.Uc&O-28(J/A[Yc_Ve5^1P?CJf;SB?b1A&W2R9b(1.aMbgPbIL8R_^VAWA;182)C
22>?Jc_P,f9Yd\V=(\>R0KB2AST?\1T(VDO77^LMDM8bL.Bb3VRE?PR<eMK=c#B@
;<Tc+&WM5<N#eL39ZY4(AEJ,C>_?CPC77-M--Y][.K]AT:e0CI1J:69(e5,+F:ZX
Q>3f0E/Z=8TPE&70LeM,AW[(0<:AASdB38\-E5?81=XW\\(P5Z29HbG7Hd]9CUHG
JJA?TCPP&Y:RK0M?ZW?B<I,I7K4/&/U&->?5]Q^EJg6V-0&&L2OPdNH6-G-<&>.F
UT)\&fP[cADOPd1DMd3Q4HN4IeVAJeH+3<J(?VD8^)>SV:VeM88e6f9J;\ISg/1Z
\;;=LBI9>/SDX&YIB3^98K1b\]aQTNFVId@.S-)(Tg@(7M60N5.SY:f(L[L^A6OE
^H;g5()7M].9?Na(>W29b77S9KBA?(&c8aB>544Cg;/:3:-7@FFM+X^?ZXU__86:
BYLF(bO?F2960=1WF5U8762WP8V-0N76[@Udf]T.L1N(R9_6PUa&HX+3#[KHQL\M
[gUgDB^;,3#+W?D:&4gAdAgZ&/\@N[,ZJ?aV7b<4#TQHLF6PY]+BJ9COAYAKd)_9
C>KbP3M,)O&V^)c7Y:H\K5=N\)(8P>RTSG)35#P^#2EVga>.N6+/bRQN?EZO<d_C
CF:@V)aSH?F5T)P[9&(_gNe5LEJ4N@#E;EGH8DMCbF8H&4K(BGDfG6JQQOM8&B2C
,KXGZ]U-J9B/^OGQ[=LC9LcF4\FXKH?)1fH1L,c/5_\gEA)P.4HS#CM-(/<?HI[R
UV?U,-e(J7G:Z-=G_5D1KDM7/[NJ20Zf-PUF0/W.Tc_aJB,EabTHUS86[O(FX(J2
&f:]@9)BBSN)+9RJS?F/K@3bHE_R=)f_K7IX8A3WQ:_7VN])/[U?S)L&:&7b33^H
cVY8RECXAJ1Ba\VP77eLB^20TK.LS+FVUf)+C6(\<:>^[#I(TJK>\DLW2?BIEcL>
]Z?b-(@dNG@Z,+?BY&@1I2<2(V2-NM5E@T.0(bC=b(L=?D(IP?,Z0P78CYd]0b3T
HDB)4MVP<&:E2K7Od>^>R)L+De,c.a.RPK=F1=J.Y.N7(c.Ma18E:K@HZg(Z]N\M
KQ6]4&/d@(_EIU>#+SPH]Q6-)4S7LXT1@3#N=GJB5.&Y647E5I@ARAB+0(P0A:_D
Bf@&+;7S7\_OE]bJ?Qc^H+]E#3A<-#G:f>Y)NC228AY@Q8J^(eQQa#RF8],CVDMX
BGTfd7OF:=bOD2BdS/f2;W7Og92f9/@A?[f8LaC]TDK4L-8L;aRQ3VSIY/2=2RZ-
+Cb:R1TgFZ+&:LCKJ)RTN:5DCbC/cFL6?_H-=X/SUPXK9);b>Hg[:KJ8I??<\eUS
4FP]1N7gZLEMIa0+d\>]gF_>7Ia]E\(U_VQ;8,g&XT_T.XULUS4gTeBP5\CM^_,e
O(AI0_2U1^0f?@1V?/)>^d[52)a))>XH:S]g6O<9,[0eEP^faXBTO-=>\;gP.20,
NM[(WXKS/G_I:K>(b]?+N+]&TbG:EYcQD@=],SOGB/\/Z_NEO=.WYY+2:<<\U;f-
F0S4R=(-7[7CIaR0J7UPfB^NWN;a-M9XM^P&40H/YT@b[^:@REVTR<Yd(HAMS&?K
KI1Q?0AU=&4N>+U7R0H:#e66N(,YV^g6[S=,c;g&8ZL5d/I,bR[]?e+G/gETM,LI
XH)GB&HU/TB1f<:H8[b5VASB>99&E8AId)VVY875<,5+^K?cM2HKT0-3(YRDC,<I
^f0]1dGcH;ec2cBL;+:eO)(5f=b=BU1&090&:?[H,5d]HEA?a,Z^PUZV4gP?ebYG
FY+I,B-47a\JV/7P61KGHB7?ETNVe_;?V;db@GdMK_GaZ_fTH-(U@d2.:19F?8=]
APJ,Hcg]YTYbdP0^C^?X3N]E)LTP)3-1?3E\;,7E_eFBF[4F&e,5d9F>3S_,:+e#
a3Oec5?c9CO[2D#/GO>YDC=CEG:fde/O&XX<+QK>bEHUb2cG?9APJ6.85WARc0JZ
.]YC_GGYZYF5CdcED_N&ZPVV?DW>6(O;2;COOe1G099<NGd@U<JZ]V,Q-LTA+]^f
J]JYFGBFb+HFeIYg?AV5/.6d/68gMHNB,=XX4^fgH0#XKC88Yg4EJ[^K=2P69(+.
/X.&RO8P2\HeX>\43^VNF.;QaTd3:=WZ3&VHAQH;@2^[JEDKeMNQg,JQHAcDaHD9
cAS/,FTO:9@];5V)(Jb56Z\8S?,X-JRZ>Y9Odeg[5>,M,ggLC#D73V+XE=\4=P]8
1Q9dfOAO6MIGd^2OQ5.c2<@X3<#(8+c=e;C5=B1c3H1#N&]B2H>>.KV^9O<OL[)?
J,8Z=G)O1J<9KJ<Y)GD>M(/a?IZ@FdbY2P]N+Y7N9PE7U)T5H=K=Q1c;_\I\31Ve
<Ce_+5[YCA+1Q(cY:aU40.NAK>=_a>W9R\U&1]4Q3R)U^a,cV--0I8M=[\QKE&D3
;.9LeRGQ>+#=91FP8MC:Ob8T^bIb1@?#LWJV7UOVF8X[U2\Q8ECYM&Uc-=^ERROW
S17V/g:1XdV(]P=MPU8Uc2100_W>9_\f/fS3KXcE>4#3K)T,FVM&OLDY>1Ea,XeQ
e?_0[-.ZS^Ugd&VFVN3JcZ-TA5MBN(-@1MET4\S[EeYXUI5<1V^;1ZWOOKHYHXSI
595EB\I]2R8W+ZNeYbT3C.##LRgA4-/7NAQ1AbQEgM?-2aBeGBVY9MZ.3\6I,V7T
\:[Gb:_2GX^B]=^-b]da]K7#S&7.>Bab]#-7/:CcA]F<K&MFIWUO89d)6/6FMW98
-?-A^J181(<GO>&5OWadA+dIHGY,@a#dddGI)A_b)9MDfb4]XHLEZ=Gc/:<8JWeH
R:B_B>bgK@bAU/33H5NUE^:4V&0+,O=(GKUZX^89JCge)N2<[2:M;dQc#HQgF4aO
SGf=g;Sa0?ePGN-f0N@c\@\T9>>W]e:@B_XRNKa4G/)eZVAeR0&+<LF-DQFXG>SW
L/17<IEVJdFN\&X&Ff-Of3)0CBHRb.,PKMB(4@KM4<?70&DDKVK,OD@Y>G6ATYf3
C#<Ve2ga[F0&=@7P4N7+S_HWF#?5PB9CV>18R1b,21.:7G0US0#0gd^[XK<W>c5d
@CXR3N)(BMGg)^bUSE#>CJW)FJZX/A,YN>H[,cYU0TDa-5PNFQM^W-F,2Td9=B83
>59I\OS0#TIA[8)U5UM3A<02OCU8/&=_e(2(8T1.#c;<IX12eB,;4?QEZ:)9JaC7
(-+2SIIB_IA+T&;ab^Mbd)T)6)#AO<-P?&,0MgW3D:1_VcNNFL=5-ARC;Xb#fTN;
/fcONGQ3)]<adGdV[MBD9ZEE;+.bM1[64&8@G<)<eJ63#6:6\)a4TcLfX?@L8BVF
Q0RB5eWX&X7^NX,>4@>R\Ca^-](N./-3fEGD3_?VSb,++;FBG5[S/VN<g+9TTYG<
>Q3\W@eWJ5W0dcd?>YKHP6YOFTO^b<=+bUMRZJ^K,RP[.(gJ&B^#;>gGSJ>eHG&X
4eHLGR1_=F^7fBE(ebRLK9RT:6L<gd;3\eCN+f)),R>aI)]U6bg;gLC8^1>F;Ac\
RfHc&]#8c^fB(L-5ec,:INH?S^@AN7(&[DB^/US^;FEVB&.+MdLM\CBG+J+K8(bR
)-DHP8,_ON19\RKQI=(R?_f]\R=@B/KR@aN;H]c)>4UAGL;\81,c7B]=[D;#:;>X
/cPT1X2gfA8[J<-f:/d+fV>>1;.&.EZQUC@+>W0d41L.)T6L#GCDDfHge)aY:F=(
)<-W7MWBKZ_<cLM&]HVNDcCgc?LKU+gCU2FJY-+Z&S=)DNFZ[HCPIW3(0:7<K<D+
(Z-MQ&;O.cE>d^2a&#>U<:Gg1CL\Y(S5MSH_[/Sb(<MaZL_,eKS5G9HHMLD>B?7(
WP\_F;ZW[B.+cd/<_2H#7<^@4XF&_@R9=4+,9gSMMM]N+<;^76]6#.&aaMJ7CQVg
E^:RI:2IU5?e5JV6MN7dZPM?Q>?10+XR0S(LND&Ib\[)/O)ec_;83VRaSc9E_VgQ
+Cc-dMR\17dHJcN;a9R6\Z9+HDV31B<W19A+:T<HXQ_YW]Q).R.612GBWP9LOA-g
7UNIHZZ,_3Ya&1S.>72OcBc9:#?C:P>\YN)c9d5L0M36YC2c#dT[03O?DAaJ&^cg
E^F1@]5>U.FUJP21Q=IQPQE8J.KGP:AH-Z67^&^IXe14H\U,+D7PA>Eb6-<17QMS
eGR+9APc(<FWC__]+9\3XG_,9ZI4.ZMUeEJCPZ].6/-#6;_9bITgf/f&6G\-d2L_
,83VC?S/=MQJY6f\J/.[P2KC_HQQc.762F>(Q+WA#H86K;@5(69YNF#AD>bCC/,;
E6>;MaUMb@Wa2d+WR9KEcJIQ0WQP\NJRc^b7b/Q11Vb9\TJ5>[\FFKb@2(6-bRMd
+U;4+^^-g0cXgB55\PFg34VE,Q7=<E-A<YMe&(VZ9R#=X(K_,-/g1RH6cK[gTW[O
;GRM+(1(<0>E7/K@4CR82C8FYZc\f@\XfSR;FWQVB[7-OO\XVB4HZ.-7U1_5B\GT
6L67\M=-MP-OQ73F(ed[S3,V)1,O3H.)B,3,Oa/<G:K;4EK/[01/c21U8E1=5W36
?T]-b+18#DW<+8+1&^MA=>QX\[:fQ>cS@T5\_(5fA2#f4CWK43)+86DKMX9/gT+G
L?8CG6R()gcY4Y,A>a=4Z>RbVd-?G3>H=/aJ)]#ZD,Oa=[Kf3P,]+I-,1,O6[bL.
6(EUCQ@CQTcb8Ed55?\3aN]WI7ZPbA:0B_;I#WNadJ)G,S[.S8-PZORC.1DY[#3Z
;/&cDH,cFP\<cQVK=Q2=C?<5]JH.QG3I3-.@a]>/a:X(JfIf_.CV>8M0U(T@&YQ[
;/]&X-CNV0M[=GM53Lag&2?K+^@AK)cJJe/5Q,B(?2V/4ERd@<.2[<a&(CT966U\
7N58dCJ5J7R[fXL:a\RHZ-6?OE-Hbf@EAd,BXZ)(ASB,WdN:ZCAIL32^DI=c.bS6
)HN-c_9N/8,)VQZ&)3O&UWJ<2)3?+X5g#D@,gAG+9d4A?MYG;X_#AO4_5/W/N\&9
b2-..APG28Y)JBS76>,c;Sc0\aESMdIQ4UaZ_CQ-c2UB7V3+LC1Wf\4e>C>GXK[D
DC+89RSNd5GC>9gRK?,C\YYZace[I+_Z.>^Td_@.UAE9M5KU.@3US&7c>_g_@^3f
,\?>)7+e55Kd38].X0BTWX]aU=AHLD#>SNaI5.<M4525<W4JI;P^OAaY^(TQ;W04
a5E#1^WHe4>72X9KHGU.J2/(\SBLQJ3>0Ja,dgG:ULRZ.Y,9795L-fU^I9D=A?8R
3:QKB\g.+Le-dOVcF74R;aVE2_=;Og:^=DW83e=3K\e12QV;P-YHAPeFHD1]2\8,
LFMVW[Fc<65SWV=B-J>-[NdC<)X\?)I^V<ZYb&,cV-0S7UAOSZ5:e6]g.H&)Qf^9
<@N&Og]3Q+eK=8N\K;]CZHMBJW,NgQ+<^0+T5RMaaCI80(:LaX\)@5Ed0U/;b=\J
Ke.-bY8KQ0..]1<6L6]-e8\Q)UZIJ>=_.L<aTP5V7-R_MRRN.[._VK6_2WFQF7A:
)c0:8XJ=25H&&M)IH5/WM;/[/.cYT&1]\e@7OA&GE#UL;DeY6M<;cC\B->:b6[28
1,NK5##aK]E9RCTH=;&C(,7.KC3]H<O>-OgS5]FW@GK[.OI@T7b)^bKgMA>DT(fK
J\>KXJ0ID4=P)DZLX+WD24bbBTa52C#/H]A6ZSX93cWHeY++5V:J6;E>,L6H-e&E
GWF0NGUfUTRXR7./3Y^.:OcfV,Z<TYeMLT[_LZc+YT>GSbdB?064/Z>=c)fGdIP^
I.E=]P(e9,Dc\7GB=eD93TQ(_>>B8,G@0#3,))9W1LU1Za3NReZ1=VDSd2-C3&0?
^PI5B1g7)<4OgF.P/=a<U@8P>I>&.\/<P<;?F\2R<;X;PGV>BG\]Zb]RX],+^41F
0:HBWc6?fJW\E?A>UG?<K^>_d9_&3_P@FaagRTUYA8/S@)G?7^WBd.LT5.G)TU9R
c5ZHF-&F9KM(4DI+dWT>_QD(U8_0;J@NQ4bD;:+R]I;2)?[f.5UVd/8@Pg^OE#VP
dg?eO/HX.5/2VL1@BRF^<(^WDRBEQ^87V0BTO.A]]W[</@TfYO?MXc#/SC6S1_^1
7e9LAX+>\)?&^_\A?Z,3[c51@_)J\:J<+]Z7.,(XKc&PR\//QJc6T&1F(Q:9Y^7]
.b,;L[?PBRADW#[);1UFEg@Y#/+&/;>e:HUW?d<X7YIRMeL),PIN/2J]fTDRdfX;
3V?L@FJ7X,,(D?GbHZ27?D1XV2DGNeT64\TWb_3,,,O<f#HWLdLRH\(UbV0;9;fQ
AeK/4<-798g9Ia&Nb=fRaXKM^(C?3TRAU-H5(d+-7O_I(J5PF[S_77D5MI)7<(X[
JDZ:;/L)QHJ]FdUNM/4L:,/C^TR3bIMUIUZO2?YB+^=&EP#CRA)e._&A:W?LHgIK
Q532&8#F-3NC9@JfdZ75[C\0@1&IUJINg[R[OI4#Y?6JdLP1N_4EL^)L)4+8WL3.
ZAEMbOYL6F>.Z43TN/2Q6Y4+,TMP@C6.+O1f^:0AKZ5/Q#C5P&@B]5<-D0M41.Zd
E-+0PTE_-g,WP;@U53N-&+e1=/X-.N[E^Z=BB2]2M.>Ta<YCM^;)_U8=B@/KJ)TB
^^0=_-ZW^SS>=FcDTZ9786g9LCI&#D3L,9c5-U4DY&R-d;O3b3bPdJ2^2dRRHQ@6
B(4.R_#HB);Ib]\BA[YC30W?7]#8[B_@fd<K=W.]Z34Pf7H\QPN#fB>YCJ0A=-Fg
gS<2>(L/VMO/UN@V0N3IF9;D)M11AgLL(P<F[3Nf2d-PG5VU&VHDfN):(Ld.Nf-M
US9M\#Kg]f7&NE;#bCL<VHaUS/HT+-SaK&<F8./aV360,EDV5TIf+?845;XH713Q
C05&PW24eJ?=Td1[5A3TB<J\:OG=W9IT0LV(6XVQEaG.RFb]W:L/&\0C+^[L9B[-
V)aG4696]=QN)CXPT3TfB^JNb7=I&d[UG_;-aNCGSDX^CBA33P.:TAQ(Ieg2G3K3
c1,VdCIKggFdgeF9f]^DCVKC.8G/3R(&E-<?.+#d0=Y4QME:>a3P^D:?VTO1CU6K
;T)R<&]2AS/6N69=aDPfE-7=S>6^9B@G7,;4,AT.<#geCWg]SSJZ&=(OUMO4#gIJ
T(TJ5O>MDJ;)]M/[JBFd(^3([AN05(3cZYHRWG3DUSH,UJ@eU9cXBEbJ>Vg]0B#:
V<3U3C0W-&+N?d+>^DJEF-,\C1R\K@cNFfc.J3-dPJ_=OXXG0=-689OV&^,.aV>U
D:<d5+[\gN5E.DN:F\MBP.5&#DSc:bGf+)B#<eX_7C,.0@04[684O@D</LD[1Oa/
[4?6gV;;e)RgQTCPKQ]Y=GW)_0J]<c6]I6VXB8:fV21IE3(.F(&R;2D<#fC=;@]C
0\-6(c5(^W4Y<+);X>L>8=M&d4\/+/I=4&^?+1Q?7_3,SCVXS2K)?66P&=YJ(KgD
)OBK&&EbTcH/02PeBeN@+9PE2eB8/g1XEbR8b^^&)b:T7=JQZ1_XM]9^FXAUKJ+Q
Qf#UaCGWXQ6XfaN<\A;I(EdG@_@FSX\cUB9EPI;2>B3./3X_ANEX1FJ.NG?[?e+(
NYVaE7P5DBcA?B8;L>G+W@2a0e1\C,I;6^[AV=8]N.]-b9Xc/D</e6&MR6KXC^TJ
b6E6PIB+1=B++gQR\bN)^1NPReY4[I+KXSLMKO7#-H<F1)O&-DNI61-4M@J+48;3
f4=e[a_a_@#87MFL:7FSGOHR8W?ZM11K]?aD,48[==.G<K==E\K>T&CAUYN44fR4
fA1<K]Pa9fQcIX=_#R@;N^)KP32FY]#aPa5f>+_A&3&_SHaIL])#S=^;^Wg)aLUZ
TWJgW#]2e[&e8@S/\38E4_@<FDDV\<1I41FCS(e39J2?/>]@\dXM8926@IFGG=15
QC7?d>=FEC4U)XA/@Ze773GB<_ab>K@(K#O,AcNYEAd?#U[_>aBf6g8;1#I[VUR[
X8P\@4T=JGfAFU2S.N&\T_7V0/J#GQ,efa1IZJ\Y/X/:)-<T@7)E64SV7d8;N/eZ
:ERB14I#a>3N3UG?@b6GC\&T.,4TZd79;)OKME]BG&>8C<+F0Ya,-8)>g[Dgd^5Y
:D9ESBLK,PcD>_QXQReb,I(YT4:g;V.,_CWE(,.ZIgFS&KB/TQ]2IbD:=?@DREgM
(5MP0I2XgE^0R[Y5,<>I(N_PbTFL4PXA<OfE\\IFXE;I1,QG7U.7D+TbW;[G7FEJ
N(&?R2OND(&-/T33PGPAd1Ge=WW=T]9UcRc?DGIM=/(eBS?A9I&<PT)L9[C_)XTg
GG@,42WQ]>Aa#&aNKJfQKgE?&+P:T/D;P-5Q_623]b;Mf79DSXKEKb>_-OVc;J.=
J7O#G;9CBB9N>;QH/QHH_QdRQD.+P\3-_)-84FOAb5G3eQZ6O&I^UePF2bVc=@K]
LNF#fV30f/CV]=1a1cJ9;g.:T2[)c2>U0C5J?TQZ\4-a7Q,C&M-VaBL7eZ@Cg3HJ
_5=T-CHY6;:bJf6d,/&S_g28Z>@)5@+fa@Z,CI:d?I3S0CVA7&;D(.:.D+I-JIQ7
N9KHdbBV]ZRIaJ:)+3VA:1-AN,aWF_Gd__fNC=;KD^.Y?3GQdYC_;[F;M>ebZM@@
9#])PSGUYC^<TQ<gZM^gaf^VX)1V>0)GX8S?,5=ZD,+=12beT[gH2PD5:GT>4AB5
WP71AS\+;bZL##TN?-T[:f_XYRW^0(K7_A?1RK5E.AYA4Q:[[?7a/E^6aF/@R/.4
)C&OgEefO?=(f#KZ]5/8CI=39e^19J;M\?G^bY)H:Y74NR0,Q@Bf\V7e)30>YND5
3</WYL=R,6A@]K^7C/+RR4-?PQYOX+.PQa:c7RN^BKOTAf?O1./8)cW9ED5;P&;4
UYY1&/XcNfdb^F-=6aF#R>^P>K.<?;PG<V?K(Y+/@2]7(JBJ.?6./g;S?\^RS<2S
\GO,fU+cLH&I=c?=/#Re]4LB\K7=8/+,Y^-BA6RcZaa66cOEDTU;a8WMeB,8DR&Y
5Eg^]gUa.PF+59YdJ8:&g,1BR)DRC&[TbKF2ZEAfLY0ecfKUA6_OaJ^3X,G3FG18
5ab>H^&2TO6=O6&a?SH7I3Z1G6X#F3QLL[4c5^I?@<A#b^6[YBa^#(a#/Ue;#-7^
fW_CANA_V@LcC[9]_DN;Ia1ONXX3JXWB6,;La)32<0()?6g8Ma-&bS<XIfD9H/,0
,V)d#[[A/bZg\FL_>B&bV_\X7VFA5(\#IEZSAGd@AMEAT9bT/&ZC6A:?7O3>U(&<
6\d(4S:O<B<_.<EEZ1^Hd;[McacA3EdXQ&&E?\-Y1WBe/^WJWc][_+1_Fc?dGH^P
/[P^3WIZHB95A?Ra]]ecY1_LL6eE,_>=]U>@#Rfa.F+@@^D7D68>=VVPGP00:@,R
B0/1FJAUK5>[Z?3Q4EIM9^D>d5C)Q6L3KUbTT^)M5>23#+=_;T+[A+.cE0YS(;#)
B]76[-<<UY_AF<LD_1;&S5_K=-6HD_B1P488Ve(N,BbIYM\b-TGaJ_BKW.C>>.:>
WIJ\O<5?47CQ>-f#G^7KXA+/5XX,g+Yf\>G7Rg>VeQYXY/C[#9\S4f)^H-,fHI,9
TF_DOT4WG:a+<LdH]<5928=W/LcJ2&)?6WPf/b^V_7\+3WEYgWC?g[e,FH9&8G_7
JP4?KaK<28SdOFN3ADe>bR9X;J?9:KJWE;UH,KG]ReK>XcU#SOLM+BHY\[L8]L&/
\b;DO5P1E[?bV858CNNH=CF5\,8^&&9M,eS/ENcXLQ-Z/I^N#=S^/f3E:L50WA:=
c]bObge<7I8DaQ^?/f(6_8>3IDYIHU+]caOA_]3>L4+.EF6/MKQF4LbK7WK(5X-P
/6+L9f1<b7O@G(ER[A[M9^<YS+&ORYF(bLFg&6/#>O9Nd>Y66=3D<Ed2D8]e.PeT
8D)-=gV\KKa>BM7M<8[G:>^?WHCEfF5f63M^1_2OVF]Re2?W-a>/g+Eg2#_;@IIG
J[44fCPQ7#2(0C(#>@6\NS#;&#bKHK5F8@XN=g]?b;/H\)QMUB:6,7)J7A7]B\Y1
a:,XW^a=D9Q2BMNa_H]CS&^Je)Fa3KJ-X>;Z7c9_IQY]+#WK50Y2&?CZQF472G6B
]@18gJHF;(&81aP6L9H-[LL=c^g1S<1/6EK-W>9\V^AJ1WbbZI7aQ4<6.LF#4aI8
K5=.-VKBX6I9+PaW?WUW\8IeIPCH^XF/UIO5HfJePA\HdbSJ[K,2+(V?,F]/C#[Q
TE8\#5dOPICL92B.M)eJQS(c7CL#SDeX@.?JQKe^22GU@R;fI;^XJ)>fR7H>.@XR
f-.VV-bX_;CI(4f1:TR.^3dLaI0;)>c^,WcA>9TeY.EdC&f;bAeKO1WVQbRS&S+[
O_SPOY</=F4+F<<H.EWfUDI&5YXP9/=)0JH6Q.Dg9/d/a;ZA2YBC?)3OME1+c&^d
_A<F:<H;?UeRQEA=gTJ,bMFTg-8JJRg]e6/99+dNMH,^NC8[94G<9047cD&KYXGS
W:RGaIe/;^<A7U9FK6&c8O85[L,.;/@Q_F6;VZHV_[UW@FH>Q&AE<=BCK6b=K78^
BV5<&Q?(]DAL7_?U9g\Y0_=7375\FS_B_X7/D>?U9I61J/a(M:dXH5T)C)?ZC=.Q
7Q,DZa#E/W(dO[^_:1]ddNN5RS1S7\_M[6P9[:0YG]W(^KOPFB8G?VE;0LQBK9P)
R(=MW+?6:CUL&dSfVHH8B#B-HC/&?eYV=bB<G+87;\0OMJK.O3RcS@J/9V-L+;0I
0EM[9(]J7Bb)V4IA&F7[:cY7f<T3KRSIZ_E++TM#A#0Z0K;&M[;I0,_aJUN2=TXK
_Z0TC&[GV<K2BY>PNf2(01K@a0dR8OJIe<\]3-.+d5JX/C5#5?K;A9L\FGC;/>1-
M,_QTP1U:Cf],9<1JYK\V^V:W[DW)_4eAc\_E?O5V#I)1.^J98>PH@(\-NOO_8f;
I8&)9:=WZ13#8=R=G9IN:aQMM]Le6Ac.?4PH3_\#:&#I--SZ=>aQFZ10/L;5U9)2
HR2F6&GILCJ\9,f[J4\JD)RXHQWbMQ8/&]g@f\KCRFE?0I3,D6J(d)eVROe57g68
_(C&2-Qg.W0KX\WWTB#(e\O\&E[>@A.K(93ML+=C6.-S=\FCLZP,(#,V8;6T?QB=
X<@cI&?QZPHe&V&Tc)0K+TdC(Rd\5f/<+)4J?8YC-PE\1g,f1\AEO0^J_M?]+ZAE
c/a+Z(g7R<9CAaCJS7,Q_Q]>E>&+e-:4PR<88>AUS7,4B/;ZB[MP.KXNCD_S0Te2
P>#@DZ>J^f09S@C:H1#4@]L4e]F)[Ac1@N+aM+3:e)[e+[WI6a^T-?G(6+9K862^
8]?[,/Y/[LJL88YCEN3+H3dZ4(H84N8fHce,84(]6.,D;N>Z5EFI0K03e2>IdCWG
bCCO^M-2I)XTJQ#/E90JG+E^F-.L;b;e02=+PV93F?-/DT;4.SZSPZF=7A(f#fVF
4B\,MFU\M2I=2OTBLYQH\5Q64<1gQ&9#5;BbU23.-(CJ6J\JB+V:<P8MC.=>UYe-
8cG2bb/=7Zc,53\Eb^Zf]OO7K:O0/CVAd0b(&G/7V.bK]1#_5N]Bf\SZc-P>4]YT
+f/,M;/-1RSA91K?&,Yg.OGc(I^0I.F]55EPL.L^T@AQFRE<^@(3_UgJ@DNY;>@(
gdeNYI/8120&CFRcb2<OVU>DLQ0RU+N/>B,K_W1YS;(57B#L[7(Y2SM^W;9W@04,
#>c>+01BGY=D\V@_3RDDUgc?aLEI6d4b_c1UIYO5)A6=Y_)c?=<aOY6/(R7>O@7]
^32LEFWK-&DIMY46:V9F1OOHEfI<SeC9S-HT1?^TE#V/,&VQT.1VGZg_>HT,;:L]
\LWgCG=_&[6CEZ3#VQ-b?b9#5#K+[2d[5,^ebX2Z0.;/?F3;VH/5=/6J<.NGW3HE
/>Jb86a->f^N@CYc=NF0[7Jc/UR(WT:e)7Q2\,9,Nc)SDPCc2dJ34@NYcP[HN8&4
RTJd//EC\N-V.J+b1>C,X:f.S?^1;CR0B#D#RS2;9-@-_[a@4RII8d^2(eg<Yc?4
O<f266OKU@-#0_S(=]]@L-M;fL4BI=fK^e8dC8+GZEc2--A?AL=TfUD#GIH[PW03
<CP.CS6\5?>>H4LR8K\:=/+fSDG]^6e1Q&O7P5M,91TZ021O7NVYSGIWeMEgO&0,
,,>HdH^7M^1baMOI]bb3?QM4X)M8@ZCA4JG0G[NZX207Oe\7IONK<PP.FTRb]OL,
3KW_:E<KL9X,EG2U;Ga\36(:E;1)+<WLKg[Q39SKU25=CcMU0QU?TZ\.(=1EVW>+
;BEX8(b)[AZ.;[#XL42e75AKBCcWX403\-(>0b26/+\Q^&Md\5>a6]?I^[P0<=6M
2\cZc\N8KgI9K_UYF#NDC>)bH/b-(cCB1_;+,JeB[M:cR>:3:W.8(+d\.+7LW0K-
BC<J//2M/?^_+&#ff+ZHPeFIc=eRF&7O\_fYTF)8=.bWe\.0+WIW-AXQ@_[YP&JJ
)12@.fe]0b:15?W3]0#P\.#1F&JRbE7GGX5PH76FW&Z-II5g_+DFLSFGY9W#d?\@
^2PZ5>JG]C)2]Y/PI6Y^X/\HW>]I&bCF\RVR<))a_3&C2_?9Pd3K9SGT94E_F^(_
0>O3Kd@(^P05P_P?JOMFJ5gJ=^PNE]RVXIY+fP4dW]E=;eSMQe?E&KNFM6UNV=Hb
,FUSR=O_T2U1+U179OfIYV#K4+a(@HT6c-aK3_DR(b9\T=0P4/bD,[@eHWJHF6[Z
()f]9VS-T1+?eVW-Z+CWD;Mf6FX,HHH\3TP^]2+BL]#8+W:+_3[6?DFPCAa6L?/3
7?W)K&7R:F9fMTSK_L9LZ]DOF0e>XX>&KE];D)W_Z]DCSWP7/SS3+#L_^W&fB&AS
SQ_^cgHL=)eE_MLO6++a396P3U_P6VN6a]-FZ@)9R2HYDIdfCSMNIbCdEU6#9TD3
(X,9S19FSA@SWHEF\c60HM8RO9;@?7F5MW=Y//8VKHfPL50(PONd?^=b[=gZdC(C
XJRAGX-g(F2#d^[?5VEd231D1K.NK^6IUFY1(EM97afE;NC]DE_3d;ZOTXMae[^g
]GS]M2ZBK,3@g6B9g.A;KQ<7KXe[bR1O^XRQ-e>NYcZd#+9f[7e.;,JVUG]AH4>3
aagPSb6(O+9MPH7H4QW&:dBR[>T4B52;8BRAS.QK/#OGN;1;a7[FBB)4QIWY/C\Y
,;PV6SJF4ST&?&(d+QB4Kgd]M][[P3H.\F]HDS70H[OA,O7H)1b)>P)Wb/W(5N@7
UC^R<,YAP&P?LDN3+W^0TS:+US13S(cF(1WEaS@BV/GX+R9/MN&_W:EU.)5YF]1:
\<<<Z_E8TF\U?4S3NZdO26:_RNRPY22RE0<)R+4DCTTY?[M:D_N26_NL=WD.O?[/
c2+,Z@H#::X@<Hb:a3>S=GF7-4cULF7E7^EO)&ANPa.Y3H,?d6TaXSdGEZK9@&8f
_f6>8SCO5;HfV\NY&5;1K_OGfP]>5D@:WCP/U81C=ZEY+[]81D^JY^CG3>C[SJ.I
e&V\=D/A\)TZDUXCbW-1/@+RcM7Q@AK>?)H/f#I.\#MB]R3DZa/X>B]f-ad99&L>
Hd?8fQU?^V+;BYW>HA5d9f^NWHXX)V1#^Vec@a-3F8eH69g,b<Y\MAcR^E\K.Ba,
OB?9XaY<fJYe^+U39&_D)AOBE;[eHLJALMJ&gbRZ=6F4>XbGfPXB8U3K<DV>JLSL
D;Wf3f_/B14+_J]ERF6^Gb<9JMO#DY@NEWJ2VJ],cQ;@0#K@<:<ZJ0_ZKE<Y-e>?
VB@8V]Sd4f^UYe9-:(CXDBR]+3]f(#7=A0BXER][+FRMK0-RcNMKaK/ZATF2G7)H
;3;W^4JNgMW5V98B]bWU:L_8VM+UAc\/W@VUcA33GH4Z_HJdP9LeL[O7L^B2R2=>
0e(B]gP;4#(P?OcW4SF+V+>gN09B\5O.613Q,4b_ZD-LC([_)#RYfG8AZ,>AZV9D
>@dP^3c1fC>cPfJ(>QGO1?;Z8O4E>Zf@O-5WM=#bAUg>_HA6,:2DROcf,;RY+NA]
0V]>d>Cg;bMP[6=8UTZOTT?/bZ5/.>3?V;FCVa8A.=?B]S5+;]R(]A4@PI1dMAU7
-=RV,)<E#[cJGcg[RP&XL:L05QIR:ZQYT>a_#K:=aI;P&3Bf>,4/RU38O5BPW0Ed
_\D@NRc3M.3YDIQbXE\N.Y44fa9]ZJd1V/1U4#.Sb><ebPSg11:M+?Ibf5.MfXH2
QFbY623H;8G(=M@KUaK+Z/fZg^T7OCQ<RTS(N7\BFT[21.,2+K:W#6Y2KP]ALP3)
H],-gNR^8MLU\gH4T7FD9H5IT?[^A\KcFYXe:YFACA]M0#=AGX>C]^BZ\CX74X:G
:]Gbd>ED=&HaV&/=DO\LO(^M/>]>1Ec4EdB[XEJeX+:5H@Y-D>MW)b7Z3=:@_:A\
8R-BdQ56479V3c9E7+#/K9,;AR+CD?QDVDGCFC<-.6(Y_LRI[2#_J2SAFc)-PZg:
b2RP0,GH0X730@S^E>UKT]KH;3K]MXaKIBR-U7=A3M[B0IM68\SLCc(Q/TH7RK=-
HKO,A#DJB-c(EC/<?8]IH/c,]CGT1G:T-6G=H>Pc\Y>/@)<:&=8Y.#ZTTSLL7-aA
-]NeE->8RF8f]I<<30YDJ4f&eg_IT-8O(Xe=^,,0<Rg(:(].AE(6:+=19GX?O0AI
V1_5SF<M;(E4+V[CZEX+RBQgdN]]].FA,:+HGK^=>Y1D2PR5L;9R#=c:&e=3\I]U
RHU=Q#=<;9##(GeU3-bPUgE8SJ6[]_ea1+Z^7F@@XPA)-G)KBQ-)KR_H[4YZI>J<
>g&XOeE5P-cB,Z[\H^gf)O.<.B3^GA2@gRdK6<((6fT(/[]WE1gF&Z_:7?4);R8]
fgb^LD+)>L^5RA8RS1_WX:&?)+J.KCI]&bSU8081DG,KbZ._F9WGbM^D/,.RbF=F
IePcJRYW7SR7fB)I<9^+fdRV,f=3;Kc[03KCP;@QTgL1PH-,-[FS];.E&FAEgQ[J
J3WLeLe6G,K,dM<<g&DWf5bEWZf)7DW;b6D[H^&a6J=EJ20>BLbS2f4J0U^g@FE1
\=9(\+(THI+D/0^c)JO0^_H=,eAP2gCK>cDYV2XFJB4;fe,^f/ZIF&V\^4/(]X0)
&b&LZO0W9VR6\ZP89AZI8>05c1e#MWg;NTT_9:<K-f(G2&f<\dOH/>5C-);SfJTF
D6::^Y;dZg/T_X.7_RaC):KALaZ.;?ME-1DR37O1J^J.-4Y7BMMD5fJJV:g,0ab1
<f_\GR1cHXe\<?__GZDVU+d3aH.e;dFf[_7W8YCH+K:9^>1CZ0\981#/6/19Y.EC
KL>PC-R1\&S@HNdD+MTAg:6OGDe4P3\]1QNGF@S@e_3]47G.G8=#A+-H=N/U^&WT
.HQ3J/R_9XPd]UA..a18\-).HMdF)R+L\fT>#I;I:E.S6@7T^<.\cY^8C+(EJJDQ
Kd(,1X(fT(JP#XJF5KZE@EFV&1D4\E9TJcK.?//KO.R4:2<ZB,:3[)JgU)N;VQN_
gT/fd^^Tg[Xa,?2gG)Y1,:;:]RE<NQHaSE]#<>.^WfF;:I>,,d4VQ0dWJ7<.8K7C
(?OJO?H0BUNbI+R=IX1X,5DCadEF=I@e8\KO:6SK30^NB.JQ/1f#]GF6IMCYW;5.
RDGCZJ[W=CdL?D&EQB:6ZRI-bMT&_)HMRAWEfO47e7XGQ+Fce2c]ODD+^]7:^@KE
CL90b2A(E0DdLEDG8a]QNb1EK53&XXR_Y:XB=>VV,^7ZbOE-66(TKI-+aCL\E(8@
ANfI[#;UD(2O)C-/X9Z,a8&UVCdZF#]6@gK8LeA:J4YZ(g@;=3MH/0gb/W8GdY40
a:X:+V6)ET6.D??70B#7?CFXRTcMWd<>7^-Ef0,@6aQW3RGQ,Z?991TOd]G]aKZ#
K-RD&40Pe4-EYM8gKQ]aPgDf-);,eDU(B,gA)R;KK1aea4f)A33&58X<8PG=Z/.e
O)@b#=9;_bQA=?a@DX&Ud5Xa]]PK;[fJT]Z;=QgbIZ\03a]:@fBTM\:dcOfQC1_9
C@+I#89CK.S)(U;NXe;V0:2X36R(G7,F>Zf+-;8I6G-e\(UE,RP@0aQ:1^RS63)8
K2d;A7F9V8C/--Z\,]/(BS0TU&A<f25._P8VQHI5UD\G@7MML0.M1T([)<OQMNd/
^d5X./?PdH,X>C:V042VO:/(VO/OFd_^Q1OK]^4fBLd)#>aaYgX3.7.OF5E1)Q,\
f3fT#6-R#,B.D]FKf730?DEBe8,0\fe^&#4+>UBM>6/IIbVW&-3Z_A=+)H/[K/DU
;1VGKg(7&10A4RJ-O7,HE=bJ1KBL(f?c1-Q,13F;49)2EN#eXQ^V9)M)-T;c\)<G
1AGFRF7-LHQH_MF.I#X[_OHD<XB(fRc>HDU4<]@6UJDYgTd-?&W>DWC8[-BYNL.O
-bQe-d&W8@HM:]\Pf0I1e>gW9M_f9]#?8EE_)\6g.#&_PY_]_XYEDWG;3eaJ(HKa
G/XYS<&ZB#ZZSf\B?X3XZ;>/eC(VQWa]VS&\ZC^^b(ffg;T/(T9=<+U37M(@AdM9
g7c><7+&Q2+fF,?K=H\Z&bD&D8fM>Od2M^2:,K](g,e<<e)=^TTUf_2aWLYBAIGa
H;MNd3b=W<X5(JOd6K(4+9M-KAO^g/]MZ7(&X+>d#031>a(]E0bA9@dIZ[W&MTbW
,gWcgH-:0#6AA1[)g)<^2c8TIH2WZ(<[#V6^P]LeK0_I.F\2@(6S3N:N(Vc/VBLb
M9dT1cJ@\Ce0.Q9V502C<3?A(?.ARDYcDP0C5?YKVV(H?ef)<I2;HNbMH@P+eY#c
eA-Z\-@N&2A1X:]P6a2W#O6S])/Y5GQ[J:B)f,9FSACA5dVVD(DCJ77YXZ=OBSQc
.?aKLg#I26)+D+W#IGc+<U9,\C\/)J>Y_1O[C.7JQ3^&H:aV8(@e^Y_=V>OHBKM/
@97fdgC#)ETS&c8f>R.\UV)ENGJg5;3APJBQG5V8)SUBYD_SRAfJEL[VIHXUN6cO
c4^T38bR7-0WCG/b<DK7S/@LPZY;I[5ONGGY&YC(0GG74K\Zd\__D._.bG6A,KM-
cPSfKE_dG8(:LScQc9b,#B7g_=5(CU0EME2dV@Y-D_86?P>[GIEd;Q5[3H#94<1-
]dXU2/_a64QD_LbIZb\7PCZGb1\:F+Q@U4Z#HVe>I2=2Y-Fc>&6Uf<<)PAKO?g52
cP&&9>:M/^\;]39<(V>DM;@>dJ&RQOSQLWQI2&_db<5=E#MgZOEeU^OgKW\5]\3X
ULU6F@VfF901a<5Bdb0:fbF^QEFV.65EY-:3H:_(cRLf[Fc=XX+VE#JJ)A+7RM]S
E95Cf<\1aBBQ\^@Z;A8))X\H3K1DW88gDKVF\3T<.a8;)P53TWZGc>I;5;@g.]cA
5GB@>a<bHD,<RB7Z\U3V7#fDP9,:&1)-G.CdUdG>#B9<H+9b4H6,S,V)e,X6PX/H
Y/RJAZF[,I#CGRaA0U4]#,R@7Pf=7R9_72FE6\D9cVI:d&#TfGUUQ]NMY-U)-XUC
GYaM-+^d_8RO?A+RX)[4Y/LA@.POD/GdO1cSZQGaB:J9C<2AS(Xg;aZZTDY<&XB[
Dc^Te9Yc>(f\\^R7MPH>^JN:.LDP\bU6+4Ie8OE6O34?Z9V&L:=\+S7VM6aV4)FT
[6_OM7gbb-BdHN4LU[GJ1a>H8QD6<UC;3LO0#]PV17(4XWY+e/?I7;8NMb8EQ^8f
-_SD,C?LbZ/E3P6&d03(PR3Pc:dDce[7adMe3&#/e=MHbMTAV\_gZ\;[H1;VVQQU
2E,B01b@6c[^&YF&:PEIdX+IXPZccR]&gTCGKg7C(,;.=3^AXVP2,e\g859E6Q3b
2VTNPMBF@3c-OcY[^H+1gRF41S>PCTgdTB&8)FS=J6PLMf]CTaQKJM4BQAN7<)[,
I-GAfL5BUP4X.+3/ZR+75FeHI/Y3+760>)[V(6Wb8VN\MVDL@EEM+YY^X#L[,K:G
dH3AeXU<[QDJb4^W[BPG>S#V?TM,\fX,EW?[:+M5^>B+3?SP+bPV_??fG.(,OE3<
dC9KMR&>)=@_dL1aG#)-=>(MV)]@6NEg>>9+JF]Ae]PAQNXJ=\;8TPLeQUPRQDdH
+2e7W84X\@aZBTe:C^(fI\(eSK#Va^FfA5V7=\ac+A;Z_.]F.L\(2DEWN/F96c&C
5IY@R.);9N>K<gSBNGCW8LNQ9>OZZ&[1Y_.=5TW(V7#HJ+(gQ.6FY0)BX=bHBcLG
R@=/4/VKM3L)1[T6(=MS(V<6?[+MIIBPP71_K[b)EOf5V]7#:AOQ)CH&35De^-(B
b;B\&,1_ZZ@f_13N@<ON(+dA0&3Lb0[C&da5T0K7g]I-eFdTf)Kgcb@Ea1Cb6K>E
9D##75C)TE,PQLT6T8dbDdH1W;BcZHQF;KS==PJQ@a1H18+0:_RUOS<763a(1<MW
[O9?]:G9>(IJBA&cZNXTfDdV[IM>IE/5&\1O7M1.J[3[VZ&S6K^U.E0Hc#Y1O)5H
GUa#S8:3Y5Sb4^?8V+HN:..d:\GcH\b>ZC_L>=JCIfS8(+JK5>>f^eAA8f)_EKUc
-GR6c3TUcED49:Q>]7\Q=5LJU&d,2WS@_21^<W6,=3AeF?EJ^2Q=bKe>YAS0?MN.
_]?1EYbR[I&5^)+-7LLMN:(C\4Ud_5)P6Nf_<XSL>Vc?]VfQ4]_b/KP0ZT2WRcY&
RG1dD@W/OU&bX#PAeDS/17,4IJG;Gg4],R/^Z.ROP09WK0;=B=:(3&\5Q[G<^;N#
>;#+&#a/IY-U]Sc5_e#YE6g+?f^V=K#,,c(:X[BeF6?09^3a9,4E4WHNJ>SM,F=F
aW5Ed)<@>7Y6M/8OA59\>N>N;ZUJY)Dc^>&ZWRA0?\=C0.D:-)@S&:MW5O^/;-gF
O51\)QZO/?Z1SQ&A?I?MRbH,)?YGQ_[7eTg(M8>P_44LDgC@\)Xd?/RR=QGd9_RZ
GVV?0Ob#FJ,-TC4WfD?.6ME3,gRJc#\]K/(LVGA3Z.]\.\K^PI_11)VS8L+V:,7N
g<>4Vf?.#FbQL><FG+c?@@VOR4V-T>cF-S0#a<3A]b:\eb589.+a]d:&WJ5=cNQ:
YB7+H1\]N8#SHbFgQX1J.^-GO6ME#1JY4c@YG_M:2X]2X:S_YeFBTW^A4(E8=-#,
(2VDFg<Z_<011eD.(g;O/C,+V@K6,/BJ[R@A68DF5O_9<.;&BeNfD<V>1UcIdNV^
LI.ZIP=2aXE)X]M<YaMM)>\Qe,#0Ac^H=/R9a>c@L9L78&2Y[5dB[4X#N0(H;bd=
)<37POK8&R<bR25Z,\<#aGK>BgeOBB;?HXDVZDaW>HU+W:K2=VT0Dg-^aIV\N@&^
?V\.Z/.H8T[P?G12N]&?RQE#3M_CMPe+^S6T)3&#E8b#RX0b/-\X1gZ(Y72W9EN#
T^15KCZa=#75]3NACWE.R<fR]PZW51I-(E:)C6(9&P_6M))fB.J;bb4f=JfgQ.,b
]&6@7BYE9Q6aN1,FG,-<C4RD4LGC#WL</LN&H:)3<SL-QT1\M\bSa7NT5fXIMaZ)
?_gM,M8#JfCQ(>#U&U/R:6Q&F_B3Med&c>Q/+@>ABBc@\a_#I]6c:5ZXJ9B(6F30
_3IR39bW9Oce[QG)2I6,U&P:@L6Ua=I</:W9@A/<WY1BcS7CdWHZ2G^L^2),T)LY
96X#=1SZEN].UE^PDK_D[YR9F^QSA9Z/CB-T\Df_Z3.YO;F79RH.d^<WGOX#M,c\
7:SU5c]M3@:49/9WRd498K,8c@fT(Rc=NCFQ>[1ZC.+//bQgUPX)E=XefFW=.HKM
a[D,M?H;#gTH[BF)D?IHeNG^?4#b69BXg(6<Yc?WXIUHM3@88X_UDM?6V?I7OVT5
R^F^]&:7fW.-:+,AKFXOIINMD>N@Fc]KEagTI25>?A-:&U+VF1OC>=d:aV#5#]S(
8TfKd?>g?<GRRV)_]E=aJe_0fa^:7]<+eNC=^DZ?P6\cFVc-Yc+]4FQCV8LM-KI&
3?J?[(6K#d-BO^cAC]3/Fe:?/G\\<5&Da=ca/_;E45JG_J7K9G6]MbT1GP.+g6/_
8db,+/4d)b;QD/=d@P4)VG-1F)JPOdOJ(H@2ed-P\WW7dFP+)F>#8:8f7,-L<VJ<
9PC<FfFBMFSWQZ41,1DE(UdD]9]efeELUN(3#gU2bJgUWbEACR[2BKIDe/DV+[7b
dK64RC\STG[H+A^XD0b]Ja1(?O+;XJ^E6CO+&fIC@LeO^)+,]R:<+IH0UN7/TUJ9
?DV21KNb;#97]E4YPFI3D[3<.2R/C7,7GH88)N>N9/[D9S1^KE,)WOaD])]U)Fgf
-_]^6Ac56[aEd0/&H2\?7875O]F(eYMR.a@cZ>X,SVXg(CZ^OO;&OI-@[2AZ.CU^
gU/CXXDF;-6PReU#+:07L1dG^QWT3&&N3ZSX/SI--a4[])C,B;EaVEX<I_OMEZQ6
(7J3>F6,?2WQV9Z]&9,_^Ug?CL6QPU/-(5D;27fa1[J-2gg(65D]U5^)Q2ZcPGd_
VY+;0-9](2UU6f+ccV>SfL[e_LSOQ)&;b#.56/cXJ,6STW\:DJNN#b_X^_aMY>((
-&_AV,@]VZ8PYgg?)TX/\-+XbFFCdL/FGI2IU]&Nf_+IBWGT=?Cfg=2MK3K.&E:3
#?gWXM/Ue/DSf\VY9<2(+P,@W-Y13YBH8JST\#fMVe5DIYI.\#V,P>&Kd;/c8Y#Z
7?T]2X(-G;U+5LA<a>TGQ2N+8@8bU/.d^0-fcT>>0+==aaKF#1+7fOAg>Td,D2DZ
GD?bIO+8#F7^a4-CF8=3V3SVFQKW)KVXA-cQG>?ePRg9LJ[31Eb])P1aOT97C=5.
PeSBZTV[PGG9[F;:7:,]@=7UWCd0YN/9H5BAT9N-8+eUf_U@)O#g;?ZFOQ3d7>g9
cgSH//NNX/f_PO]^YI/O;3OEb,6_9ORbf&<-gJ=0\<(164QA8^^IU_ZH5e0X)BK8
28ZCBF4ZUT2_-0XUEbEE86RW.JJL539b&e#,(\K&N@QTfIKHVXO&c8JXb7Zd,g4H
cIF#9]<DWbS^AMHLeJAG28X(V5DcV<8,];V,-TTF&7.?,J-eWZ:3(1-CeCH?]]MY
F;THI,&+F0P>5gO)L<DB)7cOJ&9VVc-ZY79C(E,W.O650WGOY>FR;M)IJ#3H?MZP
Pf=e-)Nb?)+\?f2,gg2ORTRMeRE?1CR&AfKd7-]?#&4R)<26+90XKLBJ,\07,TdQ
FH1Vfc?BM6A_K?&&L(3aC=).434=We^FIXdR>8Mf68W-G=E5K44A<85)d8D]MC\_
ISfLAcL):C8P40IB:\470f:Z&O,M&G7]B8N((DWAdADdE6CU_AgbMfFA8Z\E@N/-
O61\1&;c:g(Hg&1IBNR7<H3\>AHSBN5>YWHH@ba#\4=48J1SLPd)_V844D[e2O(J
HdH9LC]\0FEO6ZA/4O3SYQFG[O=.cd1H/XCDE=+1gfYB]OQN0K(/ZU@M0:>P^)-T
-Pg(93^^_:,.Wbc:UGOPOCC,eC3/Mf#A5)^WYT-&ZOXL]Q>eFCMg2=.R4<O>&&L6
-&L8cPG8579T@WXY]bXJG4D1<[EWJ&FY]f>LCYgZ/CZ\=3eUO/A[Jg,c8#RS49(9
?O\O;S^3F#_FGIgT_1?+UF16E)P#c&ZPALg]#H35SV-HMJ[,KQOQd\I+SNMQ4KZF
5,HY.9H2#S?\Vf7#d5I]CUF/.J<B/+BN5Q/QV)Vb1=?NE;bbH2Ib)Y3S)BC#A[NW
EHc3c<@M8E;Tg=#HSL>0:JUHDGM-)Z2/Nb)4?1U>/?4c.TRTWZX9\QW3eLO5I.[G
;K,R5fH#XMcT3V&,\HU6g9W=d:a[4_<8/^VKIO3C5X0VVaQL0P]UK4f4-_MZ3X.Q
fK?_/X2G9>OF\B5KHTD7O#B.OGZC@.+YA40IIQ/?0<=EI8M)&=O#F9a?6B\DgUTa
&XH#0?WORCec3VD\HKEa^YD3C-+Na;aea\-=GPARL>.V^\?@HXRaM@K3O^(e+L.a
JQY/a>#N/B1O91)(=R4]&MQS,#25X;d0P5Q+4,/7_UC\fBIKF+UO_;)26(_V]):8
/6B\[9@KC5N&5-;ROc<bGc4U0G0Ge2&P[-HP+b_PN]]2@-VNWOb(83:[4I3fA=bW
Y2KV#9C1&DUcD,,CLTg4VW@37UF.+YYfLDK5R_VI2]dLdg#;H9;]L-efK@[,D#V4
>2OMOLXH/eQP<?=YL/dB6K?ecR).9Q<<[\S#-O0a3QUOE)9,g1OZD[(8Z]1cg&QY
JX4EKNX;-P0_?0R,-XdG83Nd7,eN&R1__bgVdS0CR<G/>]1V)gcRC-R4YC=-6IGB
-V[ba2/\[\4fV<M:&/3+.I4D5J:CFc2MF&:GbWO/WHb4f;JWCM0T2J0PVFM3b_1]
HCGgaIP8AeMD;\IX5K6c]CC(2#J977ND22KaI6T#&06EBS[2OfFI@^#ZAbI\@[_J
<]6PK0C\\6c.DMb=GT:_C8-H\6C-HeIVUD]:/dLZXED-c^IOG0]B4<+g7G8^dW^#
e8J:)K77<JOQN<_C43LGEO_^M#J.T_(]g9)b-aZA1H38U15OVWF?X,9L^[b[()FJ
4DNV>6;Z@#):dE;BcMB<S+#g[6](YBNYXHV_GeE&,,N2/V^JNYgK(VM8?T77H^_d
KW]bXA1aU^<D6S@\Z-P?fC?UM&>V7gU8>;\;Q,c@Z4WSMKB[,;FT6AH3P_ac=gdH
?SO[<1(_HXDU];;=a>U6Z[C1P\V5LP(8eL=AVHQ6I]=_L/])8#1(&?WP+bgA(5LX
[U3;XT_X9GdA/4?-EEC+1JP/Pf#33VSF<CIObWd?:Nc.O9<=FZ)E9-4;8U&CgSKC
(GJ:X[;U)M&D7b0gW889I.:S</[0cV[#.V7X(.,&X1GBS>1Y23g8c0486^0QC_:f
OZ03?,V&>Ccf)D]5JVPTcfZ##S/+<T-2,]:g3;B,,,[V:a?DH),EgLXW+1XTI[MX
W0(HUW)@HOH,/&Eb1&;C#f>5:0)G+X-SHP+1V<+e7[WMQ1c&[17_CX7>[3,0.aYP
<Q8Rg6F)07,&=:-2J\;]Og1?DEMB6^KEG3P6Ra2(cDAdB,M]TE,E9)KHa9J>G1L^
,_JV\]I3ZZG7MHC?^)67[#g)<VN,.)#Sg17<.8DP];R3d9^97c?552bW&6<NY/A7
Lc.aIS8(2IEHFb+<B@HdRf)O1UKD(W;PZXE6@U[P+a&C/V+O_[)NRa:[]EBO@]K\
Z@LXV0[[,J9-cNICBZ@3Se\A\5U6=L\OH1I<MHabH+AZ_fPGDbR[3+3D+?:gffIA
fS7&D:a,J,ZJ.:_Zfd49A<BQ0B6E#N#C9M]4cQ\a/TCVM.R8ZC[Ib&9c1O@?eP-G
QgH4?0F(+]8<#W-/O,EM143D3^P,Z\H93g8H/)>Z.M7PG?4VLO(HPIC>T648#K_[
22g5746\KF#E_@;NTHcY[D)Wf)_@VfNQ_;6P,CEaH/MJ.LSPEb+>b;:EbG2Kf)Z1
@Z(#(5F78EOPU8d<GOOLKBY<43Bb,ZWFAcNTRAbOPa:KS6&K?JI[S)W/_FGT.b^8
4W^W.:\<3#DD3@RS2W7\TT8<Q:CP3e[>&\#J9WP\/1Pe&?VZ04#LdJ(CaZTK@]fG
I2ATFD?aX^BgQRCbJU5)bVNA]fX@OA_KAa+/R()DFG:-\d6P[B+][\K/&:5Q,?[1
O4FR8Y:8(7dg:WJ6d=a>.9>L2?IAEDJK-0@+H6bGCT3FL?bSYEAMf^EZ4<4;Yg+I
gXdb4__VQa[bGe+5342&d7\64aDSQS+_76?@L-V&3S&U3CLPP5Y@(fN39D?@)^K\
M.XJ8IWI>#e&K6WYMP&42T\42a70R=+1>2Z,_9BCFN]TJHQ]R@Ae7CFbZJV+_16K
7O)8]b4JWOCP1A^ZUC9:/XRV;3;gaVRN?U9);fN7N45d4Y0Ca3C#TORSABB;S=D.
[gDG,RgYd]fSZ9bPGXU5RPX]VQ9#^b<>d4LV6N&:g,Rg^=<Y0Y.B1DR)8:+55E:^
MCC^^cGIfN<J&Ia(N\UE2R]7T)d&CRV0W@M/PXN:&d,[f,8=>7Rd;LG4FKLSaO]5
g\P/U&AFcNPPe;P/cPQ0]=a?f_O,R8133.5:_RHBJ?9K9fYHFL+A.__KYQG-&?<:
?fF([d3W#BY@V&KLX.(JfUF:()Fd@DIZPMJU<0^2+MA.V15&g[Ug(X,H0c2CaU>@
O@XWGO?W68D&LQIHaK@A^H4RKKf2?]C9ARd/=^<:HX,G2,&31Xe6?N8Uca?_9b[&
<_:M0FFC+M4[N_YPXdT>4G:7N[AC0d;8UY6K;A:=-c,<--#BEY7>5dd:X6[;O7#3
g[HffI&,/1AP-2MDXKZCKP^BMQVO[g4<fd&Q.ZH5A1f-OT&e-<cDK;N-<]T@X>e&
OW9UI7TJAY4G?&b\7SX4(1M[3KH6IY#I\-;]1CcEL]A]8=AbQVU7SXR7KAD3Pcb[
-dK)#A2Z<XWRKT&(C&_IB\ZGX?37Da)N/QVR#c6WN?87YeWa9WXDaQ0OS\:^OK^I
H4fBB>L.Z-<,=;?/f_7e]dF.H>CWa^#dLJ/)PS,5+87G6L-U[>Y5<A[Fc2T1X+8b
46//>#29[9][)YQ2K&Y49F5O0V59^;6e#,dXKN?J<@Q3F0N_d6MXaFKM=.[GUGHd
H7>R/eK>f?X91TP8@Q?]S+@_OQ:3U@7SOIbYH\5LHe\<2fFYI1<Q_E(BQX_FWa6)
(;4\FE3.,bc#[eU7\WP@90g^<GE8DH+(]cQ#1=X6?3?3bGH=a9O&\bc/Pa6&c]RN
gG__I-]LIe>\&g3YMfA33=FcST(&I9CWS]T;9WET2RGJ#1=/R&V(/<D#=,J1VZIT
I>V]-.3K/&OJ[]0;FeR4WBK.>9cZ<;b8H(8_0_GWRDPA\P).egV,@67B1>N^>Z5>
?UMSR=^H9VE4fOX.5,1H5(87K0O1R<3\[-[,+Q2?TIA5.?&1?2H/@K8CL98g]M@8
P6eS^g6P>a-G)-OX/97eLfJId4HHZ&J&4P]>=@KD0[7U^U#FH,CRID1FNT9SI#1[
P_JN0W?[N?6@NgcV5,74gK]47T/Of6SEX;1#WPQ6a4#;WL24<VS2AUaIH@_9:/b8
Ra##,c61J><,GQS9WG:?Y&5eJ;Q3#dFN(MYJ&S[+E/WMG=H0<\-N7QM=eHTdC5#R
aQ6I)QV04E-=4:d7,ZE<V#1>/C2dV6>0+UU[-E<2ZW</E#U,1]IGGVW8DX>QJY@[
0c=U+0<J[)]9[.F,U<=S02;GbZZZ:^bcYgA<f-=:fJ;]WW@W^7ba@Xa-Y\)4CfY7
5fZ#=Z9@fIf,^2bML8WLT_4KG[IecHEfGA;>ICDPR[7ZXHcM,5V4QP2ND,X16:Ke
[7EW2.Y<ZEO1M^V9c4).666bB=JcE,58DLZQ0_dVM2JRbK+/H?CN-&fQ?9C->fRS
GH/]YBNI+^4V;[HD]?&9I09DW9Y^5SH-_V@>JcbcO+.cR)bXe);^[?I@]IPa;c+-
\II&Nc1;X]FN\d4C80CSca(&8?C@W_E2W?5ATVE(R;,-_I;d+ge@SH1BUMBJX]:E
SBJ2<FP8FT^X/6e2GdJ/g.7XBeMQ1-:4LX/LDMM.g:>2^(@([ASL,VX@&TKSVPDd
Q7XfAF>#M.gH^fa\-8K(-<U8LT#K@)+7Q9=d.V.PXNC_\#g?T-YdTLVRYDL(,4A(
V0IaCVfN-d+9_FJ)3[,f_+\[WG;7Tfc<+32f[,daFFCTd0XEHYgU\dI[KDbR&;=T
A>-?M6I(+&BAV(K6eN[?Y5&0AG.R+VZF[4PAVeb_R?UBCH6/-T5cL7#HSS6P=WR?
A2H#aY.EZIVVI[6Qb@O^>4Q@#gI;DHb;_]c+643eAXdW?(1&@?&7&GcSdP\PbIW&
7aAC<OS5@;,2_H-4UHU@.\Nc>df/WL+Dc/5IF-S)0ME<4A<O9>J;6G8I:LQc8<P<
E;1c&?acfR(T9E<#_/\/eVK719B.?+TW+(9>>\[J^+F.0:H&WGM_=9BI?KF8@]M[
dGD1G:_3<A@1X8\F6@K2#JW]De/=^ZT7R+-VZ)OY3LNA_3@NE-^D\UF/AC0RJUSN
-V/?5OD5,#>E2)aH-b(/8ZEEPXcW[7ZfTfc5F9]eC>PVe[\5IaabJ_GT)gTWM?:A
9gF(YQMKO.<;EVSgCD6)YOY6D?eg4/H^-Y<IaV5?1=/&GU11;J;c?+:-64K,,C)e
#,L6C;B2>V@VOg,G)2;d@B4J_QV^EZ88=++RSCc:\]KI]5=BgI48UYfJ?aMFC50-
:.O;7#4gRO7(,WB\Q(1C+@c)WeU.Q^f8fbKJBGJ=4DOB+A&-fW<982B/S8RTMF6I
Q3F0ZP93b7.B0I7#W#]b7R^V_-Y5XaNR&U5/\I&NbX>.4Q@P[@#7a32Z+c(7-R^?
6W););_D5/c1D\#a]R:F(2-D1;E?3bZ?A2/(e\R-OCLf&^VT.Ub&P6-:\/_ZP&7d
P)I?E(=G)6b6M@.,L2g9=_B1c3BdO_Cg>]:ZI-EC2QN6GRQ3gQTafD8QU6:G.FE1
RU^)#4?=D6OQPO#:a#</@gS_3/Ng=g4[dB;YR(53bD^_I<^GKdKe_1#O.<58/6eL
7O[fH-XQ]JR_UH?RW@NRW3Ta8FR<BIY+,/&]U.9Q1D\=+6b8D093&2>C>+EZQ/4S
S2c\+N7H8-5?/\0R=L90OT+#)GU+SIRaRGS-(a;WPVT8+[:e[G:[ESR[d-2N@e_X
G^eLJ^^^KBNADAJg51Qf4P1cV4TEVQ<0MZ7O?&@[bea8690,-5=TPc]6-8^/<a2X
CS4D?DJ2g4:7/0^EPCIV0TQ1\eM.U?2X.^0E\Ma>dG[7fR&QUaJI8=;>.-f#MbQ[
3M4V)[IKYFUQNF8/K2.T,[V]_#<R4_OY92(c@^>WRJQ4Bc2T69&E7aD@QA^_IT](
_cVcb<&H39dO6-:3)?\2(6^<d-d#,EU@=)K2._;dVg3[(5T[CC<,:/)d..AW;?:c
cE[O89GP-N2M15ZZ/<N^c[0\:S[,=#KT]1Ae^-LO]EL_d2FK[21=T0W0,RfZJBb<
/9?\>[:;LZX0,Q:>cQa+OY5F<A2FO\M:a?>d+E4^YE1bHT,:geAS8.N&-VVA9W#F
7ME[_6cSEJR[#(9c,7K]J6_OgFW92UeX9D/Jb:2F]@P^2?>QLDJ<O,D)S9F+FPU;
<KZ3#V4g6X0(6fH-0ITVJfS1GI(DP22(8YJ7a/##KLW^@+2a)b)J2-B.6TS^MP+(
SY>]cWSNdHMMQX-gJC&@EE3TMW8=0(@,MI@QLf8@VC?.+/+;AQ^FEL>L.O2Y)H8e
41GJG#9NRPJ(804bMSTce/>7IUKM9A4N-BE#L@eAM9fC:2NE#T/0Ma(_P6@,PK^B
@3KARX,M#cZJ>GW#>_YbQYUEG.TH[FJQ>8?XKF:=/49U0.Pe-5W:+G@:<BR:\EQV
><9/5HVQ-,+OIYf1-BDJ?c@9\7=6&OLOD3NReVG+BZ[F[<:#K7f7R3,;gbOBY7cM
bAC3:&f^ES>a_]bQ#ab(f&178;aCS+\[3YEIg;R1ZR:.YL2+2;?(])JgA(ec(=T:
(8f<.MG0#LJ(]O+QK30N(N]#J8[+2H7)a<=&F4<0T8N2/>M(-SR0Z]c&f]cgG[Xd
ODJdg]J]E971\,_,R:0^=2F5AO-AW3AW5V@OQ=6[>(H[YW27c]cGJbS&G<5W-.,a
8UQZ+EMSF6Ae_^G_&fZEe#=ALHD^ETSV2d=@K#7A^WFDF:Y.P5[(J(:P17cQMH+D
cJfeF[N)16(:<OXPAW#I:ac7UM(bL6fgHVTYBM>b+H?.:J7AK\ROCBdI8d6=PEf\
YTfJ]UF0JE7PBHYIT\_0/Bfcc8]Ub]O24[2]XXI79M2^^:Z[_DS;c.f3/^U<5_a4
?[2.PaG/H2ASX(^Y5JcAS40bO24g^6G1KKH-#ES4QdST71F:+FTefVA(1.e;^_cg
=Q>bZ<ZL<a@V0N-?#\_((#,L3<G-c.E7@g.UQ-c7<)HN?&JG8IS5UU&GM876/\+U
c-:7Fb2QB#&W=F<&#&[NKO?0c?GO)<9OL#<E.B=\?D&83_;Ua_3bgeEPOSNO/fWG
\:K^8@[LGX58YGQEI;?MP+:\:6T3,cM[]CJ0QaFBf-C;OUdZMdT(L4B0:G,R[V60
:T4O^IM1@IT,3&???=FMFbZF1D^M-_)a:Y8_5QOVQ@3](\-+Q/RY6>e=2I@U1C,/
(QJP<6M]2MP^UYAVaJKS&1Sc]d-?FBe@N-GfZR=dJV(;M9g2P;:6-ZQ]SfY_8/Y>
E03XNIV7@]_g[(gJ;?),VH<A(HOH(E]UUQE,JK&A>NTA49e,W[BZ664:B,;P]O<L
fYQHH\:ULf@VcKAG3f.bdg)&K[d,D4E1Y2E[OW.SXSKC</MIaBTPRfV8EX&7eA(A
B?dc3QLBNI6=/d[KT^/+,3)]E/A4\+Y2-@dTJ=;RF7G0W&Z8VX-cT,]g&]gJB##d
I@JbB_.Q6e<c2\AG[c-b4:4bUP(JaI.T]M8BO:452E(BS/-7A@a;LgWXN?+L8IXW
[;_U>^#2>5cY9OI\4RGIOgb(=VZ6GAT7+SZ1L;6IC2B>A00?QNVX<Y;S2RbN.ZAd
:/dL.eZ?HE:eQ))L,53^.:H@S;eP=H[DVX98M[K.<;?@^aTUW3R#;8X50:L5I^)=
P[=/K[1Hd0(Nc9J5>@(R7?J<0=N9HX[dHFg=Ka:d]X@\_4A@N)K8eD0N+BIUcW[d
f(#E5/Za#>)Ig,Y8VgY<FPC]Ea1<V9L1U8#;5_3Lb43C4I0CH7NOA/;H0Ic:7Q<E
TL/_NXD5O0CTJ^fALb]:;3_14XHcJ)?Q#Mbc&2bNW&BdK)Q-0gE;X65f,Q#5Y_Y0
dR?5ebGP8&_6d3-QH[Y64c1\AMc[9aKR?=egNdP[g0;(Ra>0^#d([Z<P[.R4f..8
H8bd=)Q68\E@IRX&5,8)FV2(7NG<LIeG6KJ)#eJRV>Q7B,e3(N2eIZ>6C)/9Z(HG
J/E<S9L1](2J7V7;+^a6S8OP6S0JK.Mc7D(afd/K6B8=(cB=HA\_W+fD]LQ5+Rb[
192VFJc7LgHPX,\e1.<6?)0&Ob\HU[8G#FL=9PA)PdX:T-LONXD5<@NeOEbTIN31
)=8;]RO@/NX0][16_1g;cN.g99VLTQZ2C(8GS^)>@W5)U\=(;N8NHaU_CeP^V7fH
LNZDM1MP(K[1L[XeM+-H)eb,B]JB6YB1)#N+D^T6W\e<C8QJE0GE46&A]BPa7MPF
=S<4<)>&C[&?@FHO5<J1_^K@#D0JH/CV+gM2b+g[AI2P;06Cc@PEQ:=Q:WLg2;=1
Jf;a:<,071D/P5[L/R@V-2:?(:a]:fUD2MR\,.O>@=b5RE43d955e&OUJ5UBR)A9
YcLB<L3aIVA.e7S3P,-eZB&&.1LR=D_ASV-9N8/(V/g4g.Yg9FC)3_?^)R3.c.K>
E^W\LQ6U\Qg@_9P[0.@8?ER_2aX=-,:1JT[-BM9PSLc[fPL,WS,@LM0EA@VZ7cWe
_^E#JKa>W?gYKR[4dLZAHM_OQY?1Pc7aDJ.YR.LFe;)0<O47YD&U@0Je?(VZCA8G
e)4BZ/]a3)5CF-?)<3[\CK5TT4P9_+0WJRcMII#K(cYV55b;FN3Z&5L/;7&)B\3^
;)9<LY(=>[;QJ2EVe=b5^N@6JH(ZV9KXY7KZIP>bG#&Zc\]g0Q/S-cB<WDY:E?b(
99/?-#EOLM5-&KfSDK4Y<<T0,T8I[X47M3Y?+(EJL+8He@;PF&Pa7K\K5=0=6=W,
M/PI4dO9S_.Md=A1LQ,5QfP;X9Jb=@ZFf(aLY5ePCd]aXE\ATKXF.\M]WOO;]aST
O_JH2dP[Od]@&O];@YeB+N72F9HI.4He>KQR7a3FUPULADJ,AKHV/FHEd?@D/S2M
<NZ>e.-0?YbI&Y)X9F<e#\LVZK2UQ6Q>LBT=2X-O283903OBf>1<QLJ6G#_OL9c7
V^XQQ7f6:\QN-P#dLc#.[M02=,JFNCQEU\+[-)QQ+U+#L8fCXRY)-8cQ#fea<00R
R3U06#YX^7H[UT0?VT7@6LZ0&ga@LPH6948J@4^>R1\I4<8QUE0dL<UQA-;VQ3-d
f(9@FJ7?W3.#(aXeMY<^AZbCXV:gVO/4M\=Z3\C1]L5-:f0e7_6;dF3^a7?_5Z;V
>_KT=f0/Z-=8GYgP9J/V.&dM0I>>+\P_;<9[Gc&A,aFS1CG[Y5S[g(0&-^;bHe<R
:O-[ZTQe<=-4@T=:B5AVALQAM.D]LLM5U]&RITYdV3D^d)3F_+]UU\&9a8d?QSRG
+YPR<O\DN\_X(L/(ccBE#FfK47JJ<XJ:Lg/)KGdP+MY5-JWRcZ2bXKNCW&K,_O?g
]17@-R52OXeOZ_L=J&NZgQ>,La1B)E0UZW#<_;Z:dG0+9CNWCN2PJYHP[g5>?Hb7
9#bQKP17DB^.:[aX67QKX/BL57OOV/O?7HH)fRfR,&(<N).(3?=+f:<;)f=I\_DV
>K]=MQH@RbN9GE#Ied=:dGH/I?b9@N8NffYJ:b?ZH5Y+-7)N3:4-R]_3=c+O)d(d
T63-(g8ULX9C,=Q\;Z]((Md5ZE,+Y/I^QD[+V:+.4SP=:2B&_T[83GG,XY3)@_OR
@U9-V\E-:Rd8.gB^SY&A.bB+?BW\g2e[e3;5P]]\K);gT1SMYQFe/Q5e37@&E@3<
FD)7_eC<)_XA(fEXP,d15._b+0TJeEUeH/e\BVE0N<LgK>V9ef82Y:[VRKf@U+Pc
TDLU<F=)\9&GJ_<SKKA>OeP,J2)@Y5?^5/^TD[0&(N:Y;BP]3J5B];C8dYBZ9Sg#
1#M0U.9IMSG0ANG6bQ@RfXHJQ?;]eT/eX._,56Z5;X@)GEG]TU:REN_W+T#4^(gR
LOeLZe1VWEY7L5J\0UgYfT:4I.Ab^.XC?K.4A6(1ZP4(6PF[JQOX\5/Y0bY1C?JK
:&.-EJ?8Se[7W^=deP.2&QeSR&CL,[(>U\84Y?H4O-(XH9BNYMa>@4H#6C2AVVVd
H^0a;GU6NG^#=cQ0E0D>QB^APfBK,dC/84<KK?2J<0&-;(UNTJPUacNKgA&5cZFQ
Rc610IYW^)L3VSK;bFSa5L,Z:D_).);#9EX-+\g&,1-SR->I8=Z5d05HX5E?/C]f
)g.5NU>AP&KLASII><>CEW)2F5<fW(TL39ZRfc^)+gGY1B^EYY5,X8(P;[UN5<[.
UBafUGWU&fV;4G)V)7]-6X:FRR/Id#/B/N44C^78#_UcW/.[KfCV9MPb,dEcW&PB
,A]D^e#DPa>,8BEL9.##X>WFec^DI<S8[[9Z>[OP-S^3VC9G+UaNF+G2M.[VYAE.
AG[>:e6.(=)A)9\[)TffTO8[4OQ#K<(XG+OWc?/gWY#>^W_c2@JdQPg1g4-H5@]g
gd+R5d=@_/T8Q;BJCgC+e@GF<[+gQCIFO0C3CD&N/Rca&E9[G38:#JAZ6DHG(Y]D
2Q5[6.8WHK41a=dJXI0?Wd)/C[5a9TI_8B#ULNHI-VOac0&:;S?<HK<c3N3?[+DY
gEXGfZ(QW4F1=_I7;-L2B0S6>-3C/()/OIC\eH[3^)=@ccGV<G2FI5<Aa.UQ0<5g
TeZOY,7_eEd6Ae-1#L]NE:ML29-b)cM07(EgNaW-ZNQf<7f01+#D#Jb>=G;I:\bg
9:f,#MW[9VDO>\2J?X;<d-3:T,_SgZVSBX/4/Ma=RYQ^cZZ?/bAg_bCSAUMQB5#:
R.^,O;/#>?C>\\4O:JSH^_LdDa6ATMF0FM^>576@MMdS=MU@V.?.ROB+C7(3f8/B
[L8YVA#[OY:cYa;#O[aY>O0:O,&656F^aD\e?.9ZI?SHN-\D[Y(I>=5BWbg;L@A_
>NVY3KCVFC(<5IW&)DQRT50/J2&SL22?(A4,9Z)[]UA3EPAI.F.M4IRS/MFCVHC_
MJaNMOH9UK0V1@V1P07N^cc=?DZW6A>ON.e^6.)7#?]]<:H[&DZB0fZc1bfJP1],
fR3f8?ca1,73RW5/2UD,&HXF(N<3DR4PCe2IDJ@,_Y=PM_&W/Nb?N\4R[F[=X2B5
.-D=aKfA:]96>MBRD:LN191#];Z5E7]SXa6Z7(HgWIZ<;4W._LX;^NW)=LY302>e
9S:9J2;4dDLDX8.B\ANfJWXT0#aJ8/4]<^Hc?=](#22@&.>V@4Jf6GUf@?8J_TC8
+X8<6@]eS1P#DFMW)35&eQ_?H_eM<cVW<:(XLM&5E?4Q@5N<[;]Y+2=.Y+#TdB2V
-I>-eA7d1/?WF_N7GbCgYJADZH\E/)8>&O#.,)B^Y1,[)JLK-0U+1.X4cI4(;\?9
B8R?P;/HOR=#/>.cZ;K035f9E<8+7?+)9gT,d1ZF/]N3#0P&X-AfXT+V0&&J9<RH
8Z[2CG&P3]?eLHM95Kg),Z4#W/@6F]-FT@@KK#6#gPE3+HMLaX+9GfDM=[Zb98UO
5>Gb5c@.]aAX1fFNR262T:[:86<>>e_AbEWY[Y0RH^D69D\Q>Z0,R.;gQdeeg-8;
5Cb_C7f[(@X&2V=7IAVg2HKBG72JYd6(DTT,dO>fWOMOJbHbEe-DYL[LOO975>J\
4O#0^4PFW]#R1-@FC4XfaggB;&;da87_^J0T/+d#d@Q([1KTc>5GV<R<<E7IJC2:
BF_SR9f<Pb\Z@6=O/:G#a4VUdTC[FL@+\G-W<ZXX(>^S,MfFaMJHVZXG)_6QZ>\[
^4?f(]AL_=f\QOVQY<-c]fF13&Q^\1OCS>24a^QF(P/W.[BU17E5F5MSE1bJRC6J
T4Rg5S8V-eTS+XMaHD/;TfB-9S1;g(7Te+UFFDVBgN81g?\W:a]>1RD]VHMV_&&2
L4=]ML=RHBIVfR()&1T68(-49fZ\]F[fS5-BP)gAH-PO+2YZcgaO?@W?D)^.P>#f
KFFK?#)JH=?HcXV/6U>)4/X-g9^/0ZTPfLPMfP8;8ETV.eeC8e^<9f<ZINU6MfbX
:a-R^YU\LP^\.L^8RVE/FKV^4d?47)J\a)J58@AM^fJ9.;<0dEV-UPK.Sf39/MOC
/aM[-;X[d12L4>Z(1-R-1b9Re&MQU^R8@.=G5TE+:X1FIG/[9>48P6Z??^(4&9RI
e5?4UZB3LJ]+KLXc>/g3<4O>^7UgKT&?g=SeI26;Q6N2?Q;MEAdMe=dASN)9B3VH
/CN-4=QcEc<,<5Ja[>/.EC8H]3@&ZV7ZD6GSCZ>?3<,5K90UR2S)EI7,g?L&1669
N4&f@g)c?9aO=O(P/8(b0V/b5Z3^KJdKdTL,KaRW&6=)=cF/]#;6JD>LM\3&Y2#(
F-CLgMJC?+AL0Z</#51-e>MJ[;LE(a+RT]7UgG#^M&Xd.T>I9_EAM_/0YQLdgW+A
[QO3+4]U/a]IVYHN;+d.I>>3c<a6&\6;^@e14B2;G1XfJ(8/e2V[;:L?dRLK]M/M
IZ:+GU3^)^GZLYeEdHCSb7<(+80(]P&P#]R5c0.QAM\Db[R.;+@4V(fCYbJ0FT?V
28e5A[MDHP\aG].7(\6/TT#Q:=59-JMO;@4?-\B.]S2@RM)3@#RA1]]GZ3X]^cIg
<DQG\UeM,9eN?S_WU2L5[0;;5cYDN:TbCe(#a44W9EdY1V_(a2?__CO)7=2,&Y,:
G2PQ2ccNP0>R<ZHg/#N3&@_bB8W7/gWK]<G??.-gAZ.HRVGIGJ[QOgF\E(M_f+K.
LCT:@@P20E0Yb7HO1#cS<PB3f5DXZK7+Nf3[(S<9WBW/_C+:C3-b.1[g)L38B(K?
8L#7VC^>PNQA>HKYO7<@bD9-/77CH2IW0AQBf7Wa]?_]/[48+_)?3M)Qa\5bA><:
_)I>a02GdPN5Pdf5g7B35Ad]e(1DVTbfd\/8=Q;[gYc4R5#Of-=\B[H0O+?:XCS?
\NG7?3QSX50bX.U,TC+IG98>\c^H.<DET?TNQ[3EgULJHBL[[@N9AdQE=+Hd>6CP
ZEa,1fZ3:&I4cddf(,4>^\M-0^ENL3K-c225f3I]N0]TZ>^be0(<X8b21MdKL-)+
<]P7+PbL9-(dgQC?2QMJ\Y\M.,Jf1MB]5NFNMOg4FTG;[T]??U/19a)5]N_V0Qe>
1aMDJ6+>gU)CMa.D[Y^1O+NYJX(E]9P8,/_29FB^E?VKS;?6/.e8?H8WFUee.XTV
Vf82UUF+1QTDYO00-:/,V4,2Zd]Ud.T()UO5,)PZaDC6)FK#fIG[<D1<65<+aZbe
([CN5V6>9@:<^gW(K;+&E)(2UTC#Q@;Q)\G5:HA5Zb)GgTXYJMDG2&50T.2OPTgS
^X+.Pe\-\d8f08C1#\^E35(eTLN\[M++cQI<E0dBbSKPFadX24U3a1J.HAD7W@-;
-HNf92/W=N/>3U]S?B,=--ONI(gOca;]>.f-ER@4E84DL662gJC@a#E#9Hd2SH>8
2Q(dJ6d/4Bd=&9(fb>a7?IJF_BUB#?,Pb@O(aaIG,Z]KJQO/eS-O9/,X7c5AH3,7
4T:LDa+g/V0;:PI<EX(LX7TD#4FOe)ZD#/P_1gVW5CWdG3[4eMN>f6;34[gbLL99
HV_)YZB-S59BLHCQRBc:)[#XJ7^3C^&2WA^F@]#M?fX7/.gNM/d,bMX4#(S)JJ+1
MZ\eeMO>3)W[eM(O&;A6afF?5fZVYLNMa?:@^@P<SVZa0X[a;M5W74PJL7M?64@T
1.I)FJQ<RY.dBR&(6#G/GJN13-@EQ+Da+=0R=Bda<dg=;Y,)AF39RE\TN0HBIFGB
3RK#N-Va)]<P_f67+PKW<8(EZ?gG#W2/S=H9^_;FG[]]SE/e4A1H-Q^]:RdFQ3aT
<<D.QFbX103LYC@IUS)82a:3J&,>I-VfGE[X=UEM?TWb\H2NWO/AHI4=D#/E1;;F
(I_Z-VA&gc0bVcG4K6LAUW\O9<g\CgJ-,P\JIS9.SfbS>FWX;FaFPc#5__Qc><gI
J7^AYd(g([a=FgbGNU@,5E:XA?3X&(5K.GC>VUN:6)FTWD.N[&T+dI_[2.=D89;=
Rd##\.C4C+D-a-QB-2=ZY.,K#DH<g9gdTI),>JRX+DgcJc^[=6:,e>Y]S,\.F7ZP
Z+Z_EVY?<2WVX-3\.F]PHN>45-MIfKdY8G)5?BI\7]<fU2]/604H)@(RY]>A4S@a
B3RD_M6aM<Eb&6dL1G@4#\H7Y]2Z&RSMTC91R,_;&2RF4P[0IP,CZMKf-F/M4#:3
.S/5PP//EV>VegbY[g?X0YI\(3O=dd+_A,/&6N=,e,H-MKVf_g?<)IL#9D]YH?cd
0>Q7E5eI7gP53f;F&g6?Hbc&Q_+?e\B54@P\-6@:OGe(,=3)H&5?9-+U#7Ya8&_2
g>R2g=VG8K\-.V&b_W8M9PHA)GIXSa^X0e-L71.QL/B)VJP]fG<,SD18N+[VLZTF
^2U=?EJ8I71GRC32f:eNKgbd6;=EOXAe5&=/3)dE(82CUbA<5_b],4F))[@WIN<)
B6Y^G)74N(OMAe<M@J17LK9&Q[K3UKEI0-;[Z[I\\SC9ZR37.8>@0Wd@;Q)]7[:B
-e=40ZZ(:bY_93g1CHFb9-4VO5KK=+O1S6Sb3e@X2N3:^LLg)9>.UTB5G4.IR=(V
MT+>73bO>7E?TN#HO(?Vf86B[g_92bf;REID+ULV5,UHR9]Q_-/R\+aYXL(-dZ+P
Igb@[#3+LMaV=7g,?YKVMdCG:0UgZX2@P(@&CKT)L&Jb;Y/U8(UM;g/7^@_B/CQL
Fg29b[^OC_bY7OC)9QeHFM+gQ&>Q50)(6a9V_OcYXc/XUR_fJT^&NQS(AbA>6_XZ
K-b]-UG5&eTN;^K>K^gNB[&bO5>0#UKJe5T^;-><Z^;f+@,QB08M)U[8OgbI=AMc
^O7KeI0+1V#dCdDF]##?=IC^N;7-^0:[]+.30ff9RD:/._G&gP;^1P#BQR=IUd]e
cAB<J++<bb[6:SKT:)RHbEKZ@6D09415#MPPbP4<4c)c:_7#cf6PEOd1WZVT>-]K
H3KOEea\VeM&\,8U.bb>^6[Y,2@[W,AG[ZL0@R2S\:;\R+&]NVCA25X-E?8bR\20
@SS;#UMfe+9[GOKP^>0C#G+>/-/@UGTOH:34aeF>B>a4M<,(GV40<Xa@<C3Z[e8+
:\d^3Cd+^P5\PINf#ZYLQ#;9b-?6]bHS?,#(Pg+IeXZ(>f60gI\2-,g,I)3QeYCD
<2^d1[8Xc+6A8PAEN,TP2.bZP[O</X.MGPL_H36[Y[a9\T/?NA95KBCe.=f#GS[P
ZX8P+A[08<@fWcXf@=H0&:P?OWa[MV9EAg)#)BQ+)#:]K>O41_RT>[(3H7YZ5).S
gS/dGOVU5O8V\IV7=gM,X6@A&C<(5M_\_W,g4O5R3Y(@A)HBLLSHQcBg\68cL3R@
HHaHE\,6Ab,(8(RF7I0\J8\P_gd&+]d0aWfd966A?5?4C51V:g/G9)\,57g=XE8.
QOa+3]2f:NUL/4d>N?CFO,daY[><BdddW#,O)6&LPX9EC:RY@3cS6=C13>?#2>&U
JA-9#?fD_S4YYC_,-RK/VX/V&R=L=D#;IG4D2I)3TZgFI)e9Xb[5]HV7cg2I7&V4
5JaP/Pf#6MO\2/TTGJO]SbPQW8=]#TDU;e:,IcA4@)D=I<KKT;dTCHAJ1/,SeGHM
IEI1Ce:1:dQMd8Z07JTK&;]LX#?RSNLBMAd4B&HbF?YJ1B?Vce?LOA4AXg-O[eEG
R++W=?L-HM,Q_C^1?_X3\#0UZO/-F1UG-g,2@-;QZS:)IU#^gYX,6(6QS;QO5]e:
\BMe+9=PGO#;68SN^_+.1.Og/.PbdBca/+TTMU3GZPRdO)?F11T)30\&&D3PZ8+Q
eG6API-Z.8QFS)J/NYCDMZ7D@/G03^@^6D63fRT].#EMcND4\H\gWeMDW5<a8>H@
6FI#Ya[d#&5-VC2.JV9_^c&B:5(cdf&YC[(./Ga5NIXc77abSGETU]TFM_g21M7U
/0/29JI@5d1FGB]?WBI<EY<a,(3.8)6FSP1TJ0?IbRgL?B/P_MKR]>SIQf[eJ:]e
5cRE-FLgWNBN@W[d0V0>12R\_9M9(M,33DB2LdFe;YKG3HOV&\dHL?aC^Y\\?EdW
P0M2QAc.^fcEd6/MTd&Oa_\0AVJ5#\3^4<F<2I]5)9UL]9O&\YI10@Kb;\3E0CE3
F_\HY#8/LDW=B9JY1:=M#U,8X(gFSL]dd_MI-CP&9FF/Y#I_KL[d6&3fH,KG7>bB
C?\DMJG>PM0;?0QB&aGZ#AS+e0E&?aRWEf;89e+H-[PYe(#e@&(/VK(KG@]&#-gX
T08e->H>IGK9T916;2aBgUJ]T@3cA9J[f&V6(@_-?.UBJX(cd,ILQ&M[?De8EDF^
Ig5a2&GML84_=#6^RGc5:M@LU42Q;F<a[C2E&,M/U7GX86]EKMNggc3D-HW^LG@R
@SR2I,gZC<gN2Qf&-N6M12@^B>L&cE).(OU-XTB#^]@<O>K5#<2,V2@I9MHU>/03
H\-ZN#]301O[:VX,<=d<1@S87850#1b54-6PSMXa)WL>NRP+6BA=?,SJ@QFY?a,B
860FD>RE5;Q&8.MEZ<S;]8]4#BN@OPDOd[.9R),?6^NIg(YQI]DN[T+QB-.T3XX>
ODVSDF6f72;80H<K.@S?XVI_7>;J4H4)N<1-Pa_/Z)addB?2EZ97g4K6TT<.c#e#
N64&[IfEDSHEOBcQ](ZCTB@4XWGVJTa>VXY_D;0=K&I;CZD;A8KXO^.f_>)(,(U:
0Ue+>=3ARC>3Q/+J-10K?&dP7afIK#F?\D3DCa5[P/Y]<K(RbF<DB/SfeDZ?+Kc:
;dfIO8++JbX<;L@SSM:NRRLcM/_OK5I&?_Q-;F()#cN6a/,N&AQLZJH1@[[8HD4Y
17RNSIIfe2Z#&=OJGPE<7_eY6<d#(T<70PV7_Z):9;OLc/SK6e-JU2URT0Z6M1.3
DB3SH:K?9BdLad\C/Tb8+[GIQ=P]FSJ<SGYRA[_]D]MH4&I&Ofd4F^[X&4bVe@+5
90-&2B?JM1U5;7&-3@M3\NT=fZDJ:B/X1GW32>c#=+JX9_Hg&+Zf,UJgSZ10DJ^.
D(3=&-3-\-T#;.B:X;SHN.dE]G[HGI=+-C3HO5V,1:LI9QLNf[CM<fU4:[Y-C#NG
4SS)E3I;W6+)W:TMbN=@IG/=D;IG_LJIf,S@&#37b&e=e9#OKMM(93\]QZ>.S,cG
@Z/QN?207IFA[ZV9cV#CJc>:>Q8&6;C:2(TQ9)61N;89Nb;O(A(R-A+aWIV-@,<+
=?&AB\N>\^4=3NF(gV7]cF17Z2@>PR812^D96QH7NI]NU.ZFYW9]1/8XfNBAL2,8
W\NZ&M-\8=9:5M,=_RHN1FS8ZEX,cW:,TB]\5e8=N:bAX7AB:bM:/?.E;WVQ9E8)
gYE8\FDA_Qdb-<F2AQ400#2e,eE8UL\8;OXcY4QF#[Qb,TM6d=SMP1cW>;,2(@G,
77.)_c/He^7E[C(C;eF6^F5e)W0g+@G?#GcA+IU[PV4US.fA>Nae8DE,R,4U,D(O
L]-Cf;[@^_SQ/:<^]ZB^UJF)Q\V1:@MJ?7/NL8O370cFLMN0&/f[cCYD1,feWJ(f
CE1&.L_-.:7-68GQ28fc(F)Xf(5Uc[+YQ7=4/[d.L#SQd]RTB6+Kgfd:P7M6I(R5
+\(5>D4/&TELU,d/c4.Y5>Ff[,DOb;V:SPK4:#g(3H9E-MA1HN&(+[3D8C2QFTA_
ZP?SU<+4[9>a;&/]B]U1W[Pc7]<^ZFe04J;g[]b;M&@E4Y+[#ZP]eM)TTPZ\-FCZ
?KCe-MIfCa[TQKC]a]Pd9gc2EU8O1R@MX1bAHS@MS]E=8HKVOEZ4.R5MHEeH-Rb(
M.fcC\_#8&6N8AN/?Y_EJ3#b.0V&fe.dE(D#7?DC?F-_:2/>AeA6I=C>1e]_A:-D
IRAJg?#K+464XMJOQDV6QeBU)/<<[C-85b,5?XbC2Ng.CW?cJ0Pa-XQM+/C\e)ce
[NF(A?b_1[WBD#.(E<?)P8#30RT&FX4<_U9gefERPP_A/eNaDY;&V/-FC\a[[CJ.
W84;[f983D\5EPdAB8F^S5WC<:f8Td-SgI+4a_Vb;JX.bO0W#^2^+AI&6fG[[S1Y
CW[]CZA75f_4)//,Q/8:1OegMLg[^W<YeRaa=>Va_>aX#Q_N(97NeJV:+aF8C1JD
:7,Bb,SWf?<AE__@[\P^eHOUL^,S9)V1d:WT<Ya>V&I_408aO.?g?[8ZSIfQVLOe
1&2:]817/2AK5<_&)#;ZJ4P0F74XcCbMA:CBG<d2[Hb1\#L6S2/]:Q9N<5C:B4X+
:T/PU>W;/?fUdAbO2FC0YUZ-YSHK@O+6D#E][(^bF]\E=_W:9TIb2)CXF1P_YMT5
MJ0.FR/^H]KZT#Y;_d]/S/TG>U(d0;],;:A;a4VJ#==]_,F(5VX//E\.\Fc=G/9B
HNNgNb]DM^0&00XK:UL>R9Z;)15#UZRO^c_3FU/NKOF>H+(,_5YPPN73Y>JK1Y>H
P>OP(R7/W]KI2V^0/BQPY<ED-I3WZb&b4\\OKKS@C#b/)XM)1EACSKHJ<@ESKPXc
5H+J5Kg]H>GT5,3J)1;>DT3TP(+P&a8/8P:PK6CTZBLf;0]Ue@d/K7O<O+Y55=Y/
_#cD_@3Ncf]VL>A1XUeGFNd#L&8dH&MEG]TO<1(;6]1T;MVZH-P9R:54gg7#d_JL
XVBZ2VN;^])Ggc<f)+NYR2@<1CQ\YH[c-d)-S-DECYb\]BCXTbO@->d;1G\J5&MN
6:(V;>RFaFZ-85=QR@-^32S(JN?-,^5U03U5MG4eKSb+E>)<8a&/L2<_]^02V.gD
OG&5]eFUXVJ9)7FWdF;^[Y##dVfAc1+/ePB8@<B\B:\E)EXER4e9EF79V:[I0DK0
H,:e?QFQ=2WN+f5C-ZS1f@[d>CC,L=4MR=J&N[L#V=MUIcY60767^+@866<OQWTM
WdG@,<S18)6PU=dS_^0A>VM:0SBMCX#2RS2T#INR[A=Q\BUKL(Z-V;2D+#J(;H=0
E,Kba@R+FGg79AA,_9E))(g9]Rfd[T<Y+dIWgZ5#)ga2af@LO6B:TIE_EANIY=g,
gBBe6K;=O=A.8Q-[;LAXD5XO:UaE?g<H&[<2@eaSU&Ke.e=&/QRf(T7)G;d&bd79
0aZGM0]3,WSDH3GW7#fOS4J@G8BX#++gHId,I5S+Q?4=:Me98g4K>(gMHL=6cUZN
b9[<1a2VJ\_6.TUP=d_WM75>)KG].+ffWBgWb4@YXI^b?M9B?J+HBT\,7AR,6N4W
VW-4PAReF^,TZ1J;))C[b,EfXWSQP:8M]gIg/8--+cG5-CD@GO3CbEdPQK#=-N64
dY^BOSbYOOJg0cVXcI/a\=)UQVBcLGG6(73N#f\TeO7<a177EG;5f^aE8Q<]fD46
[F?&-)9g[^GFS>dXcV3HHSB6(@Cd:]_CUN;4J]#OF8fZ;?L73HW\0<)487\=ee=+
&X+>.3f056aDDH:BcLJXaR_4=JAAaRZKg1<B_e9fQW@:&N2NdPa9=4U7PL40_BVW
[<EZc>QBMU6;#(FV^VfCHb?5VDZ;5/]9>MV5F^5L4;,cXX_^cMD@:>OZ>RCNM?Ne
7Jgd@\XG^ZEcLM-/R6H)?:JJL-bM@@^W(&)XO-gH]e-EVeE&D<.,O_bA6M1UcbfP
TYQCC,gSK>H2>=OE9bAES(1c2NL[F^c)+Y/VA1;:2W0TQ/=We.HV9=a@\3OK7RV.
7Z11+;fOC6YC#(<HA/=?^SCLfAORffSEJDH:7O2Rg.c,0<Eb[/WPP\H?=4AdAE)U
+8R505Q76U((EDB2/a9?-Y(&L>;_P&SN2+2OKE3\[J0EcZFX8f1L;?A:/@F=f9]g
#G,6bE&]Y+Mg7LW9)9=b(\<,ZLL8ZS]A7.^18J#?eO-YJac0E1,)US5Jcf.Md</1
.6E7@=/Ag43-U0^T)E]g27-LF[2(_LDeWC<ge]H0VLHW50K<W.HDB#K(^7T2+5RQ
JK^P1gFLL>7YZS</_FFQ+Pa/FD3PMB\a6PJ&^]<7QL+)HLD4(LM,YI9EH[;,NEO+
7LE/5)XJ,I5&f#aa)aLVC0d8.RUWE07]YRPBT>b8cbg;WSNeS65[<TK)&PYW6d]Z
D\deW\H4L-=]TD-RBXBd:8dT-C&]:\#.G^-]g\f<UE8R^Se(\:baMJZH;U/=7>^Z
9^I6>d8CTLQB-OA:@Ec)d=9GD#+Z>X39X140P(J(33WZPZ/6;W)90AT\d7_cWg4>
P6D+JKQ]-Mfa3[8Y]_X>-V[AJRg-Ke?_.#+P,:bGaVG0Z[QKKf)WK]9a+^D6b()_
5=FXc:LHa^8S,8#F7#Fbd@.2c,SONJWO6]PgU@/>XZb,EWAcI3M86MaXQPgFL<+4
,..IEKF+Ee_VH73d,+e29Y1MHP2RWACaHTgUeb8](Z&YO,W@U;I34-T(+G0:UIb:
:@.b1,>N;8fLC@[N/f5^3QED&F\2Y,WbV9V809O-e31X0WJG6a:@2d2GFYO+97PZ
3gM?B1OQ\@=NY9D:ZCPUT-UO]NSQDYD#GJOI&Y;?^#F\g4.[PO:1/GEN6]DL1/WK
e9Ka&AY8)0V5>Ja(NbE_DgJABQLF1@CMIb?:RIZeWOOcE5A802<e2)1N0>QAE[87
B)ZV6S)>/]Z^:ED8eVfU(1(QW5QG9eU7NPa?C;^E&N=b:d,A,.YY^+J_03;(=HW=
\.JgD5<[@=d2E[[ZYg&TL+2TIDa9CS1N/)NT@&AP\7@A([d_bVc_NLP2:26^+XH>
;DPI,FLL,94.XS[ANC;Y-/?<FH;#Hf-J;2&#(/-=KaU[6db;^-T8<,HOfL3S+M?M
2X#Jcd_/1Ef[)4ZF78DUQ(.Y]@(Q&-EZBeSM389O6ce&]W@T/^?^<0O(EL&-1Mac
=-.L.A)M@g5SA9G?-NP0cc69V[9.06D1a;bAeQ=BW0,<Yg+YDJ:?(S=RU+GX^UW,
AWB]ebXdP<:WMYU1<T@L#//I_A^OO,>\_U<SB-J-ZdW]_XSE>61B_7FAMAe^NUM+
[S<@3HXa[/YOK20EZY55E@[Y[J[^\O8ObL4:J#^fOB@M[;._Z,G.6:?1b8_Zf_3M
@\;G=3(/FP7.&=+?O@.YS7X1LITYEg=bB];aG#1:V@2c&\?A;Y4KK5+KABL7E++H
@YN291:J@[[8X;QSCd:5XfNgYQ(U?,&/AHQJ><f#A+a2HPL]<T6X,XG-b@H.S(NE
C<B#R+MP<+J<:C@e1W5N#Nd]dY?AE+YG?9c(E;#Tf8W2BZ?_G6N_+VTY&Y5FAJe2
Kg7Y^7^G+GOP1<HT@7_]]bB_(><0^f904a9-LQ?d\\-+,BdH-K1#3-ONR/1K61gG
RU6C?&ZSPb][=P1=K,P.O,H(\&\E[bLP15C[R&bG+Og;V8:P,H58EUSg0XM-=,2N
J@@c/G1#G9[(bR\-KULIA?4X0O/@<)@^,<<F8-UFF\<b;6G\FR,+U4D1GC>Tb#.A
I@\D^YK&Ha,.&IcE9QI;]USAZQVV/E1([19B=)>@Yg<&ceSB.8,>[N^+5:7eXD#\
eK^,C3ZFUX:#1:Fg3><c>/E.WTM0<(.1ZXNE:(g^-[;,>:IJN/?@EWT.U>HfL15;
QVa>[T6+<0;LO=4)cC<dY\<>Y@D>d.4/Xa<-0@PJ20Z./YP-;^EHW+BMWdGG1EFL
4^g_,ET#,^E</gd<AEFL)e\;R?bS&gQ.\.L&#-Ue&;EH0)Q2YL;B[6e.&Y]FRVD@
KHEQ\d&HF+#<#RNI\GABF<L_KN1N4fdFW.^)EX)3?dM6)IdT,F#MBBHY5-/QFVIY
,KeHc:I?Tc\LDa46S_[&1;T,<W7I[a?cWHGP2I7EZAJ;P^)QA53>L4dcB&.O#CJF
J;G&YT(FfM3YEH^A^Uc^I0V#[M,Y;_0Y=C7=IbcZ\UG<9cEH@gbR(^KeF1]B_(BX
38+e[<gYMCVg6bDMKaDG4PI55MJWOP(RbfDf&(C1V.,1G;5YD#L7g_LGTR,L-?2)
7a070R\?(;CE>@V2f=I^Ca<+P=1S#2K?1GG4A:?F,d8L[S-e^-c^0:Y]d4Q5D-g#
2FSQ\0K#_QK(+.M2J,,9Gg\7+G5FU^E?#?]A;CX-XR9HNEG<IF/VLIfg0#+&F0__
^f]\]7U.#/Y\ATPc0UIF@Rd(Z#RSM1/6:1ZM,9/8X7S3IDQE<FM)C?d[.N2H>&]-
1N+G@+W9aDW.:_4GR8N)Ie@]/2a[3O65MaNW5Z85W9L_#H^^5?TG_5PAW,]ZSQO+
8V23C@CDaD[/NdOWI(D->RS,?+BC3<D]=:O_B1270bGF((OD3\NNUYY-06@AHMSe
@9<(P<NPLF<,EB.?c@ec1^BOdB^-1,W=^X@1S@)WNZ@9X]ELg[J9c7A<;Ke&P,V]
BDWB0&0KT;P=8Ng..^_ATZ;b?ODH=DPG@;I.@Z9AH2R?D^@]&HUV?2\)\A^HcMT0
DR#H+[?RUE>e^+F:2JYA98<O-d(ZT<]:NE2FgGaMA,N5eESg<.;J/7NNTK0KGV#J
>8R[,_MO:YbNfNM<P_IQ?@\.5Z#LD1XYEG(1H#RE6-3/;)P;GGffM\P=G<9d1))-
_9&,.(ACP/9B)KK;6(-]DD\aJca4]]P[ID@0a_A,@>T=@R0.gD9&fa>/4[\88P)2
.^ZWLYPN7R5e(5XVZ:)[H\XX:dJ3=_a9fg0YIN=<R<E/4&OYcag?37VD.>+g3aXS
KP[BOTFZD0;KG+fD]>E#\Q<G^]Z0E>RYJL\O@4(,.#dd-b?5P7YHW;J0N_dC.WRM
TJ+\GK;5\=6\&D3VAE3REeW&+74<&92BJ9>CD].]0ABURBPH]F?/gKSK]UWE(aK.
0A0]eR1R.,_>A_[K.)caQSB-==KCJ2Tc[LXG\L8]S6;7Ab8IY;W\g7;2?LCGN7S3
f.81K0R(,E<3e;7@^DTU7.H@W+64,B3@;K+.EY\g74fRgO>+cF4IJJ3JA@_UP;[0
/FRQM)O_=PK33AHDDNV>(SN.;WZ/-\G-EU5.Ma,EJ^,8XOBWB5b4=.3XUA-D5d)Z
82H+WB]]^YSXRSE6P3?R:KOQZ3Y4X8+U&OE<Q]+HJfRc1(>8F#;CcAB]Y67B]K9@
_MdIBUV_O.2:--(Y,GP#?FU+-CG/(D;QRI:><+?:MgQ9U4<1-QH&JB#IQY,N&K1=
0(>K?.-V\UDK]V]&9gM:M8gA23NX^8/Q-VfMYHEVB/A/HBZ,49J@f:>N7SGD8LP.
26QD_Og@VYgG;-7OL:[TM;XO68;(1fX.g=(Nf)8S&]?JaS3X9=U_@_P,be1G_+4g
ZH8/\0\eZXB9Y(K7E?2cXOO7(DDT=2UUe,QFBOd:M\)==3Q3/V\<H_+Y.9#U?]69
FL3-eNb1PL8]b_5=@WG4FW_KFe9?GUVBfABQW)P1)N]bC1Ic>KbY\_^(+(\#g6f=
U;G&FbC2.BDY:BWYZT=FRQD,[9fQI9K6Y=P?[BII56L1:#g\SF2UbJ9<E@fL88C9
?Pa<L:BN;8>&H1@3BE3DagX19AaYBG=?U?J^XHg[-4O]^H2SM:.Y&\,-G_NJcQOI
T8Q?AR]=S8:UL7ZbZ\&aI9\F9X&Ub_eTf\D].?HBR]X\b9Xg^(T>NgQ-10U[5OF&
Gb]7B)M\^gR+UQ3;Z.9e2\Z)JKd=g@VQW)-2\Wg81O2:6(YMOZI[,aJ@](R-M7,/
VZdWG>B_#a:?3L)R8>5R(HLHVB=H(-0M__QE>>Dd^d\NU7[ED93S/KA6[RA+BB+X
Dg4A.3HIdaUAB##&HB#]0M/1H/:2M_0_VIXO[7ZP47J(RZOg5\Q#[+STHgY3(E6d
MJ:G5+9M,U,fO&LR[/dPXIIH#ARWCJa?:TVY5TdIMK@:E.;P1M\US/V]E1JD_7//
DM]fR.:]Pg(3=V<aeg)\4ID/f,U-aF[af_I;<2gb?CE4.YdLfND>P=&4g]01^<f_
Te,QHZa.\c#763;O<LA[N]K[BPecXBEO(+EaG3MD5A#1N3+]E@J#0_&GQR\SaC;X
;-CW>aW2--HQK_d&ZE5.<.2C0IKd^H3f+e)bc(^,3)fLLJT_E?a?^ddR7\LJbeB\
U1b<]+J@\cZ^KUF.b#NTD+93bLI+7V\G2Q8YVDO;C>\-X.,H/8f.)=[B.cf&Q__A
Pb6,#+PgKZ]a:&?CD1B;?GR40f#.dLK\E+]Qf#DGX)>O(W&X\+[P:aOPGg=M1H,c
CI:,3YGA@c5EDLCeY3X;2c+?]OfgOKN=,1H]US_N4P(c++1C2[6HHL<;6/0<-@ZT
ES]0[1=XP2UN#/KE89Z\R^PN5,H1M7LEf-)M^9Y@#5-=JP/1Ib:eQKKKK^7<-fN2
9TU47/J?T_L]N<eIIX,4=cJQ8aO4P()?(;<6NYAKR]a^-J\N,.GUebU9MIN[6R[f
[#E+2-.QJQE]Y3QY0c,9<.eaY(6M;P>#UK@1X\g]DV1V4N3U5L4V0\.O74\8VAK,
=\P,74/cEQ;-SgK#c>a#Jf7JC,2^@?gNAD+62BZGDX<f7=eg#_&MP@--3ab(_9BD
COd8\_Bb&UNc=:AcWXF)6&(HX=OXC.A)K(Q?:X-U<[GE7?-<dM./:F4I6)BYT&N7
FYCK3.gM@??Q2g._&KN9F1->Fe=X<MO41<]GI56-];(H;cI&)P,5U1K+Ag6RYHfK
YB-<,9&V0QYR:^3b3/Xb](b^dGVY3RZ:T5AdWP00_@<Y1b)?YId3.X\+E1;Y;^-e
>4)L4XGA+2@Q6;D(M^F.8303R?#g38LZ-_(E,?JX8C<R?54dfe4-8.DAgQ81T7T2
H0gcC[X9=aED[M5.CTdc-]:NB1G;RNN@,OQ/)?)7=c7VXR#[=4M??F28]B=9/\I)
<H^cf-C7R&BV9afG)<YA8ZC95Te:8-@SH)J\.8OV2U^aT;cZ5A+PRR(8gJU6,/W@
V=17HWa2VV]@8HN__D46Y8GQ&1a9:]G\H[gV29QWQ<8Y.I+Z#<c)eS(Z(-Z>&IN:
65]d,+fOe]3,ZI^Q2XI1^.3A)LJC^+G#UdSa#D/_HT72981NR8Z&LC-a):FHQCaC
eA#_7MaY]-\QJBeQ7GKRGUO,#73eC^JGB:X;/>HMI(1,4e4;E6e1^6UX&(:CPMgA
[&.&J;b5SSZbHAd#d2R_9EJ.a?L=88^7,):0\XF&FZ/4N0]B2#LUaOJN^^M\E7f0
@#b@1+4G[/K+)\Z>8?L\5([c1&;KA#(KGR9/,WMJ1.H^Q+NI&BKC)SDY/2FCZ#<,
gXD81L>J^Lg:0@b3@1>^cSF_Y1U&RS^QP=\AWSO\W=J0Re:e8L9DDM_&Y.(D&82U
OQ6<FP&(L;+^XK)F8RMFFTcUXd)BVWbcD@.;Ug\TVLd4O#/\.ZbD=7R_g?:c[.SW
E\>\2,N0,e9K>3aXNVFAS7L&.dAPfaQNbMd[g&;YO8@D19fJ,FgC9Q4?PNB-Y^9V
W8H#,gQ0^7\.6B4SN@3+@c,K0V:5d@a6X?1(dgYE,(?:[61(K/Y4S&574B<K0Yf)
B5@2H\D(R7-b?RSZN=@S8G2FS)SRa4XZRJ,0e#9:F^<^&<^Q13K)L2]#P#Q0EF6f
Egc]ed<H4+U6#H6?[EPOF=H#Y8f<2/+Ha]HAZD.BY/+UN6B?beM0Q.>@K[NZ?3_L
ebdUf0VKR71LI:,5\e.B/(YU.<BVXMS@bJ#8/-2(EM[U/-PHY\d(6>g^5>Z<3Qgf
_)0IE/OB1\6?Uf=JAaeS.DSX7Y0;[V[Eg7#21P1bE:0O+M+eGTLS]=/[\T8CG<JG
Hd\0]_PNcC<<(4:\2PM<Y1W3CX+?MZ7UK\T@)YKOH7e1g7d\b-Z8PZ_fB/W6ZfB2
f_6Ud21DIOIXF:^=_#:2FHBK5A.4eWNK2.4+<&TMc:g+QaU)K)>1KaC4C5D;CPA)
S+Sd,3CND^(UCa4/V/07BgQ[B5f58YBec:.YB]X0\LENGT-6,/3J=V9Z;:E&6U;[
H08^-RK>2:.ZeSSK(-.UcJ0Yf<7GS2DBC9QWa?0?eI43YIT;N@6M3+eF.C\]fL/I
;F?^?R\(S5C#:M9@C\;M^3MP=V#B,LIEZ7K?a;N9[7/Xg5C:SBU6c,3__C3QD(?@
cG@)e47X4B^050=V3B[fKKM&f8;a0bGR?R^f]=EL()V7/1cK3<6VN@K=YBI<3<S4
)YO#,dfWeW-C4>EMa4WZ@Sf1)Od]XMDX[+,<(NE:A?aB-)QUG-5gI?fJ;@LGF9:S
G[2HLJ_?f/4?[(U^bZ9O>4+18E4<[g5fH4I<;0OCf@ZX/_Dfg+Y(F<)?K^a]B/eI
9>P3H#2[0FWYL;>J\E+O/JM7T^;Q<?+@.T)f9V49Sa7]gAK3OUfC=&bW#8]D+:R5
.PR)(@22D)0^=DY<ERU.OB>M&@Qd4f3CfU,HHIYC)[G]BQB?/]OZWae+]J-(1)>7
IRTD5/>Ad@<JCTD1;1KDBQbXe;QXL(VfRXC[X?6P6E&NZS>D4Z#URA:O-B[7c\Q_
-2T=X2#cQ;H0:@SWJD.@g7;YVWA<EaQNFWFHV@Z4L]PSS2RfSQPXKNEdL[LL(b^Y
c6gG4\aUe/R,S3-ZF&:Z?7L\cX^5A8#Y\SLK?7<JI44TfBQ5dOD[0<g4>Vg3Qg)Z
+Sb#SQFPL<1[HT@.3?.B,,gUTTHFa+ReDL.VXaVT(Y?Q&Hc\bPT\\W@;dE)0?1e?
9A<3RQ+_F>P(7=U;F\?E]4=U+&e5g#Q3:<=W&6a8-AG&-2.bTTQHa:9>=_a63=SM
)beQ1VQ.c,@)ATG,0JC>Lg_E7D-U[gR:_U.Xc;@K6dQ&>aa=NYXY55EUGf(HMXQ6
J\;I.5IX1+Q2-M7^Z9a7AEI]KX](7GOeacIXZWA?C0-(7/4;]_:&PLIYZSEAZ\RO
&O^?VA4<@a])D)YO^T6YX#WcObE,=T)#2ILe4AB7J<O+dc/?J0##&gSM)]=e@J2G
S-?.]-X+.)G@=6^gGU</UTJHOOZ9JN(D^]9:XLT9-N(82D@MNH;B(0RX]+LAPaC-
>De1WUWCI_KG9McaZ+:)B_cTLJK7;X)3e>Y,e2#3Md1_G4O?K#BYDEB/+>e9]W_b
EWaEZ/-/A:.#=9c9.B[DECK]c@-N@?7IK;=EH<X-BfS5S,W0^Ba?RN=RgJTN=>;G
6e2_W5OV?\35]Aee?ePeG^O:8E7ZIN-B&Wc(CbQZ1+AH)\bd57EVP)^;JY8?FL:-
0C]>GNYHgZ0Z<FR@8+S#,#C)aYPPTaLSgF]c5C/F#V-O]-N44/#XT8,eK#]:#&Q]
7eS@0@>dR1CNKE9,968Va9P=B4MHD?=0JRVSPB=M_PE&5]B46>34H2eYgCDZZ68\
bP?cZd[cd4Pfg?g7cQN+)f#eJOV09Wegg2;bF=)SQPaBLaPY.ddg>d]C&VCQCO&c
E8GY#Ef7X@X:QS<T7e&\)BF(4[-Z(M6&(AV^0_dQW36M,E4)1RKTcSH\17cPT]N5
f-9gKKIM[>)9W0IS7gAHHeIJ<6_]K[7Z/C?TRb\2+HAg48K,OD,eOE8[@^f]\\Zb
A&)?BFb=EUU<O+RcO^>U(<RR85(EROO4]8Kga0EfFBA3Hc<,8[^-2bdA]F4DPY\U
V<^1LV,O)@Jb6:G9cKbZd/Dc<E&#JXOd.SeW(-1K59CJ?g\I)fXL@aL-3.-GO..W
?AOeL2T]D7dTWdcVSTe__L85=N@fLB@EMfc3-EWE2?1#Jb,RV&0Z5=][8V6/M1bC
6]cAa5)(7Zd@)N+IS[MQgB2#=(QY6+Zce?+/GMc0]X(3cCVWbE4C_CaS.T_NWfAe
@7+aOFO4e8UUP;47IUANX^4afCO,AWQ.I+AV:UZ01A?-I2G_5.B.Eg_5)94+V7<W
_8(4/]P+=/RRZ93a)-6JLTc4WND7F4W>EE:OSMA/C3O+W.P,T+I:CNO&53Y;::eT
8O0P]S-8A([R4#N+101_\L.#Mc\2C#?fMJRYb>f6Q4[)EPfNC(W8-f_?4Q=f1\KT
:?Mg@<?Dc>JLI0eVaNeMRXZ@fO)PUIa[G<MUZ>-Y_J9QV^2A4:cXTI:/K5HNd5BV
J64N4-<L-24dX5dOAB3?8NB3R46=V@cfF]>gADH3\/G93KKaJF4e_OCbM^gQ?)Q@
5ObR44Z2McEM9#P&A]]C\dK5PYg]5\;(ODC=>T7KD.f?3-X-Te[;XIHeC^=2>C#g
_2;\,X3L+UUXdgSVYK6^=@N6.,10dX0O4:Z9g(BF\<?>d8cPCa,,(\L:J12BQYKD
9N_K@CA#I](LHQEQ;e.<>8Jg.6?Z<6&5f6)&NLA\KbW>g\R&YEP)YOIFb5E?-]?B
S5P/&ZRcOE5?M&J:EH_Ua.DA25,NNRbJ\(?c0<B?53:H42Q=^b55MF^HDa4eWEE&
?=/,RSI1QC@)>@.^24b8#/[P6[b=U50,MceA]5b;GL\W#Edf9E9\;O7K\-1?C:I]
#aQD/VZBIN>9L512:M<B:.HD19JHO>=VD=SQ?.f3[,T,4_[ZeIBXUQAEZ&.Md<M(
N_(b>8eS2Fd&DI0C-@a9MMNIdZO\QAK0cXDA/\\N^Q#C2?N\4>#Z1[\=]+/a=cI]
=X;:c;/Q_ff(C5K-1T>FJ037V0M5E-;IeB6&1dH6R6KJYR/8HH0-c3@,&92NYb-J
gFb6]F@_+S<Sd7D5(cPJ58I>R2NPM<:+eVK46@fbF19@-T2&b\AY;U-)HcgIWU5+
eW(C,M>aC;?WNZOIEQ/)\G,&@Nc(V\83I[T7=_Z5,-<:]C[LDPFY/FKeZ3AOAeMF
#.TVSe.b):9(WC/4<K1PUOPaQdHa1VLEMW)&X2_=RdS8eb@2?WA.2/bVg]DaAS_?
@g1@F7/5?Pe0_a_]R<NR@]a_R2B_(f0<SdI](AO&fND-/\,++ZS.ADX2Id:]J;/6
CG[9<;(OIec.;RJFd7#K]5[E7BPAC<L_EX&0?]Q7+DV,e_C0<L2RZa_RgH--]4ES
>2HKefWH-9WILecFA:eO>5fD<dE?,3OPZVM\5-._6W3UC552\c)496R_J213J[V9
AY;O^R9HLWG[+W.^f3O_6OagNJ&(R9Z2P2G;S#:B.-Q_c?D-)FVPI@gJ]QUXUKH(
^GI.,0^Z7#Q8.G+93K6#1R]J#0<f6KZ[W0YI9(c#_U0:P@XV^M_(Ae@##M?WC]-8
:cGc?d821D\Y^QXD-X=@bCV?T,?OWO&=)RdVPU7^K1WOe6[P<de.O+.L7<&d9Z>H
RL-PH68+_J8.f+T4aNDK.R@_R(<\A^gF,-,7+<0K/G9V9-]KIYXb>?<2#DR+7=0E
aVJ;,N=+SVX:3[L6a>AZ(MZ>XN&[K2CN4@g;U9#W:3\g&eR]#?XaHIV>AZf6.F:X
)D.8B-[C,PYNL.6375+,_]FVM[-D&G3G&fDEY]QL>L92.RXY5[&:DJ=R4,T3c[U\
YDVM.S&C_NfF:aUZCBNIK^[MG<<1KD0IBM=6E]V-^Q?64PB+,MKT_d5[?;KRG?;=
_HIOB@7K&EfS/e/Z#c)7;32+e,JYTa&V1cU9:AW5CcDc<F7K,,[0XGd_(-]03\D(
V-#(ZA:1@\Q;\dO+:Q;D)P>bQ5\c-I2D<:]Wf?BaMDSD0GSK[]DWd-gEeAI&_W#]
fgCHKdbDaVMJ:AW-3:@UYQfZT.3U)^SFgH084FM4L[a=/_1fI<)F8.G4\6N.d>Ea
)4IeL+_B8MF@A.AISL=?C,[DNT&WfIgA(YUaf<MgBBbFH65g)F(&KdG0]L,]P+8P
f:g=NM;P7b[=bQ82CbAHWC8Be9,/<JX6f/67:EN_B/][#\_PV7OUIcH6&<.dSSCI
cO>K^JPMVDA)b25LSD\:<[#T03OD:4:Pf^DAU6)(Ba=IH=YUb,YU@[dK8)M??&)d
f:(L@(TZ1OTD-[8PVNJ1/=M7^Tb?a)YB+65[]K&d_:\W-JO>_K_aFAN5\TY2eGbI
M(VZ<4ZEH7-RG5YT3g-06@2)RZB;U0/9TVS_^KPCKe:J8ZE>ag-b9bA+DFMJ3e8(
/IDGIVdA^N<Rd:[bFN5Q^-79I/U+1g+TXX/@THZ/TX<8/;ZY+>YfR&-\1RL^ZdD.
6<e<7T/?N\KS-C1T@T.3BRK5><Y4\3=E]TWB&8af(I(=X\5daOF=?+Y7AV)PU>4O
?.BZ487?&Q^.fR=SR1LY1T:&);3P4U1Mb.(+A(dbY]6b--E38,C8f>VB(4AWfOP4
P[C4\e/&;g2RD.,6M2eQV2V1e#g8M,?YE?BK=#<fe7C[?ED?S+?K\2GV<2MbeZ2S
gHRI2#a7Y57SSZ=Y/I_-NGKgeR8:eZ[+:XdQJGBaPWB^,SDZZ>ZRI>a&?\WdY@d5
3>:I,d=g--dNFIQdH-BCS1K,D9_FS<&6dIZY<^/:R.QC@+Q](Z[e9^/6TAd=Q#e]
f2dYW__QO7&^N@/G6]9T0>1L[@[eK(BY;>CG<bI-,//\\gMecYL6_+)[)eR?@S<I
O>#cCHU83\^HLf&E5]TD]KABY(&]@;:L_]gcIE<793SP:^HeXA9E)O0?a(N)DJ]2
4+W>Y4RUQL^b@>?@DR)++<7We+^N;57F1e<=TZLV/C=SA]>VGa(d[0.1TDX-W.:/
31EJ7>Z&8DTGHa\,;a(&7f=+#C9^\ERfFM@:E>G?-L4IT,093;D648#b(5fJ-8\[
6C,Fc.J0Xd9FGbQWY-@#28;R62\d0H7HS..g6>eO+8(-D/E2K=fMBOWU5S.WE@C5
[4BP.D^@=_bC0W87(.+<.XAGS6.bBL2fVAPEDS:)A6Va20OTOQP?C2N3OY1eA?Ld
fHHH;.7ZZ8MDA,BfY8<Wb31G0?_.D=23JJfVJZ3Ke,HMC4FN1[K0N>bZd(U55A[_
eRf+=7BKWE0ec-[)d;O9f5<5GdXS@U4F1RWTa#JHcJLA1.,):2-U9:SO#)__KX<W
McYEM?R(_U\S9YYXTB#SMPFg63f>E:,g;B3NLWQ^U#/(;]1>5]^>6Y2ce#f<d;CD
#2A)?REbMeE7T//3<&cWa\_IP=UPS<0+@P9F=PQ2SR>1Q?M6;,>6S4dV0@QY.Y44
N?W&M9b5gCX)]#a2NH5\gcS:2ZU+TER4RL8IW3\TM,Hb,O)@U13M+@I]E)?c#OAG
@a:^.;5/\7^5We/PNE@e\=?G/f?5R1H];0;#&M,GEC_fTJ=I)fA+-0;_;#=gT3d/
dV?8G)>25W-d(-I_[U^\,7:79?a[PMO?9N/B7b2B2YI)=QJAb[2D80(@:PW3efR9
WG]\5I?A(LZ+Lc1:g:fNTUBGg>OHS#<_Vd<e7L)&&@b[OXc0BD+=>_a&+RT23&RC
d3Ng;ZR3A.-0U?JVcY\g3f5@(NCVd,SN]0Se?\-F+Qb07O6CE,e#/cR:aLSG/7#C
b?=B/R2cZSgdK4HK[-C9Y;/_8-dT5NfbVQ8I)D0g5-)[EV;87H=7#PZ)N-_NXBJ0
d1BS@b4N;gK.:D(+Y&#fWLdR1PZ^f7,R&C=P-@QBCR&H]X//QG#YYfD]K(UdJ6&W
W+fW95&+MD,VYNb2^eD?@:&eOMDTO?9_=ddO?)J_47@:S-Vd;MA]W\M8fY@ZOBeW
@1.1D>XAX(:6\G@=.4V?.OJcQG)6QDY:1<&VU4>#6&;f6dU)J(f^Mc)D&HFWH+<f
4f@TKgJL2RXe4;>2^&=,2R#M,&1Ke]RXSEB7=RG+C#NIM^g7TefcPS=5T=&.4>2Y
KJ))TS]BcL9A\&3QD+S.CJJRI9U,gQCALgW5#7D_-GgV\_\J]M8/WbgZ355Ydf^7
;cd6QfIP=,=fec_N#S6U@bB<FJ>TXMd;NZ?1(R=Y@LgKM4JOaaRRO.UOge84TEb<
M0Q3\Q/<>YWE:#a0._<[SWT5EATI;;J;F]8(^S(,F6.\CbSgaQb>3:_IP8/Y+c6=
+@c^_EdcdOfCA2f)9(Tfe1#I[XUKBQ#<_[d\0T5:6LAX^8(@&-6[+d9Q&L\aO7[e
72826KJRIN?G)I+Y<+7SVQVLPJfC9FI22#bF>M88ZLVB2/>Ac.ESZZ_ETf7TUDW6
]NEA)]/Rg34Y51;X;G<Ze5Z>[0^V2>(RFTS=T8(bVVIb\X0>=DBUBXXI[6OQe?5W
N/fVEB1YUOT@D-;=/@]:Y]-&^9NKC)>;eNJD3;FS)X4?AHe2/KFBE5V3W_,91^:=
_@d.Hc51aVEO5G]>4=+2&U,W:^g&,Qc^=3g[,dVf&=4;fPAXY58N8(1a[IFE8CDg
S4]aC8P7>Z,\g42RHZ=I@E/+f:8ZS_]K1V7\\BU[.Y##HDad8eA[\A1<@TS6JgR&
8PQ=QA25GbEb<O^N>6b.=,+;#>FPO=@S<f3J6OU?)C_+?Y4]ODBF=#FVHXB0)-KH
]HBO+4@9O1_-0+>H-?C?g6SeWb9_-;->75B03G<\N@&7,(O:Yg?:J[V/Y;bWb,Q=
TS_7HAMA^.?RWMc+^VKJ9([>YA:WT7EL2aFCS((7SYaJN3;5UB1]^]e+bO79aM#Z
B@)7[c&eg[&U9/R?)CO<E+BV7OFW/c#)RSKOTKDL?[K,A-B]/D8_E>^?-_:gZM2(
32<g8.@3&BH><N\bgOaWP@@P6,2cJ8JQ5TRYE)F9gC=6J&=315S@+Rf,aTBOY-M1
X_&f4e]5MG:D^QN+]T)^3[gQS_P?4MNV)@F]-KFQ(C#DPf:978&BfNDMOIU4e6P>
6XP.6+-dNcGNQ8OM)ZOMd/F5eXY2SV]N/=OF0gALJYP)L,[OA^<K,E-\1(VUMG\0
FLWc,S#g+Z(D8/UU,d^?Z3P6G&J9H\)F\@C7L4ZKQ_E&[OaNE\f+4e;SY^ICLBeC
eK;J/JCK.ERD&?Ed4L>+N>-S-,K:Ca&4JLe&\=1aPUccV2P2RCI9D.2;=eg6(&f0
FZ0Ebf-49bccHJ>50c3Q9A3)RX)MMX.YQ33d6PC(cXCUa8_Meg0Q.YF-fT[UMZ<b
gM_:7>F#[cNSH+SWNDMF+80##95<BKX14Z=_W9F=-XgcZ<CR6]Q#Q7Z9J4bXPE-W
3PYK-ENUHQ3&RPD=F9IL2+Dg2=6/;ba8fEV56S#SF>1<fE(TCXQ4YTNP7HFNFb9P
+-JdRSe).UKaON[AB6B?;C,NR.f_9a)1=U&ggA+P2+IC#I#1XGO@5UTR+.K[aH>\
JFWNTGgE]a46BAN[H,7dHA/Pg95(J#J:ZB<3O5Q@73WTOW>9WU2f.<AIeXV-/8>M
(?c)+J[bTg<d,Z;T3/T6R_[^]QH5+_?IdJ5KW[gdXYGU-dJ[4/@;SNQBU3DEQP(6
0:-JNOfDXa2/VD>[QHTaE#fYcGS\;YZ#d,WM;[X(CB7&R5\?#J=LL\S)8_YI\OTV
bJ1S_R#8cL32(CNgH#2H].2bM6K-dDZG=;1bX/+cZBBcb?gce[X/XN)FJ/>bGbF+
WZ&KBVRJYgR-=MS;^62T#@8^QTWC,Na/CZQDI_6C(::e;)DMA+XU<(>K5(SAUg4W
:/-g0VJ5R=<,\7]C^?S7\)b?CX,SS2NYW&-6Bb;d5=(B9Y3UIX7Yfg,3>=A7ND=V
:-Be8:S==b5NgY(T6#<N+OH9=^:eZf^^)Z:?J-;,TB4X.,Ode]-a4D\=KZTIF,XM
IW7LI?5Lab<F6YYgHW0?)WUGM#6d[c(M&BWYMD3>cfAPV[JH:WYYJ(&5]ZCANA^(
9ECA]a5&>.&_#]4QMAOU2Q8+OYeQ1g8f+ZLEE;.Te=8g;@cJ,;g.a>]8^DIQdTB/
5[07+6^B.PX@EJMA0@IeC-U]D&5#WRPIGSK3KL/P2I:FZAMYXe^6Ogde&O/LO.eT
<>BbgIP;69>M=Q/ZFa1_UfC;V9S7AI8GI;/9?AfC#aO0HG/c,.GMf)Y017JPFJ1V
3K6+LSdVE#?SB\bQcH,5?+e?f_01Xa.Z6(cIcP0PX0,SEEUgP&?<C#Rae3dD>5(S
Y5//8c<6CgB6ES(O#XMWKY_:UZ_bX2I=5O]W:Lg-Vf)43e09QI:6]--Y:FP=@DLV
=.KNF53IgG69P6g.8J5KE4^U_C[9K90B<J-3K&+?,edW?c>2TK&DgU<2P<MEG?dX
X4O?Tf3D0/f&I_8<5CX&T1ZbVZSZJT24-B^X)GQX]+Q[8/TOUMXG7#(RXd2VZa,.
+IY9SMQG4K6]b=d;5-J+cY/],VBR]U(.@]6BRSQSNc[)de;aDCZ]5-C30+F=\H7J
#WeE93aTJZ33b^.N\(TQ-M=g_]P0/E86-S]6=3ZJOGRR/D+FVM3bFFQPPa1^[(79
ZY#&I.\?^7RK#)@#?dSdC>1P@EeT[V<#QGe@FMRHK]#cWG?68=C(MEb,FL.P(5)>
S<g@CaJKOIU:+F?N\S].4_FS2W&:a/RR(37<+>B[QBc6@OUBC)H)Z?XAd=gaA4_;
RYMI1YEgR806ZIR,/c(2K-KYHC;QVC)_b;?DbXCQT<EDD@O4L7I5F#]>:]-de<cN
HBg[G-1BN4;D+L.Ha@-N;IaPE#T-ZgO/Q1X&S8T^(J@]e&Na=_-,::(WZc?6(,+b
Db3^bGU95B</2>I54HDFKR-:C.L3<G#F<TFf5O;EM7=fO&P?:+ac)P#gZaZRQ1VS
MOU.=A9^RFeC9ZKJ]/GD+A=BX=7P/KQ2M0f-WQ?9\gfZ28;^>?PQ71>-89fY_\,1
UM2LJ?aLf;&J3?g7d>UL0LN?P/[^OBC3SJRJ@CJg;:-b1<R1-A-V5XSXPRO691\\
3.e)]#Lde.+>A/Oe3<7G>C+&cc;8CKF@.a?BF[)7XD>)[bMWd-D]a]GYI0e<P12L
b)A3WfA_RO^IRgAJC#Y]c>4_B8XKfbDA2B2\EVd#4C/<H=UIC)Q5&gM8J2@,5^b:
H+\JT#79Dce<;]BKKcSCQQa6F7O^?,.&Bg1c\OK-1QAH]74ZD6W=HWeF+(0:N^+,
4,).b1I?SH1_2bNX2O&f-_.IRAgPIe0aST#eWaACDK=_R-db[,Mb[JKQCT,1JID^
?85I@LDPS>H#CDKN9@01c=\EM?W/Oca@K7[CB15EX#EM>4;:T<J-5UYH3HEFVD+8
EbKN31PR_D(S:gYW@e9Bea-^GPE4-L+MH:eC]De[3DdYY(K&0/0W;IB,0JM@eC,&
Q8C:SdB0=eX8U,D;BI6I@57+cFe(,VWbPE;T/0W@61B1Bb)V=[D=L0/BKE[E&;IJ
9S3JG35W+K3BS@KK@8\e<E5/d9]3/TUF6/:9223d1X?g<KXESR2\/Ha7F+TTReg<
XV3#HMVU57KLW<HD.6^,:I]T[TAd7?&09O\]4IMbYF8LJUY2TQR5H51F^H_^RK55
(;C);?HR^>H&;GONagUHd05K09_?3_4ML(7M83d.TXF9&@AK7S/fK)Z]e)]3J9N<
FV-<>A=:W#-<BE/UY-,:FKU;,=RU0J[f3PI#(/8IB@eVSX?=E#I\YfF\.UWB?(@F
2g0#c/=e[,J7AG2P:6+8b)^<;/:bX0O+S[cRDIdfEK?a?V2@/6CCARL:R<a]J_aG
GR<_)S.AR<S1NVH76,?]E_CI.aeA6)W?6_]d@PgXH#GW(07))8+P^PdCEgL#fD/W
dWDK9H#M&3JH>A,<M,:G,^0f7:a:>=P+XeXHZYB@AcS2bb),4/ef@N;3M5)9A)a+
6Z5X/7S)a;NPeKGS@T8&,=6?L(3+F1=3Z5<U6OK>[4A#;QUg0_X_7:-?G/.&-5=E
0=gJ4,R3f#?LW&ZP.7]^=:SbNUVP0/D(IX^M]RA?D9D;V>6WaHO>SGdY9U=8^5XS
;=g_8,JU4egf/(SN:Z/2F11-][^+:a&g+bZ7O?](4b&/1d^5dGY5a\>?@@>GL4+J
#c1)EL_/3)1]eGH/9R7?^Y-UD,4+b.:98<YNeb=_K#I5/FI7CD74[fA@K>gXX#2T
J<KT-#NXY=a\]3VcYKA8F6G&3FR7/Q3&UNOI\O7HUT@2UEfCV03)L5T>D&?FZ1+F
CX0XD-]U@TfA2M>gOOR=/3N<f1;V&;BO/9FLd;CX4Z=U)Pb,1CcbVIAacKB?J2bY
YM6X&:SOVJVDQeGUC(Sa@OG)Sb?b^FKC]1AB=XMFgBc:KaYJZ5C)dG=N@KVFR&;E
Q?_I?d)0_JN.B<Ig9[agabK5+I>(P05E/G6P3XZ3-:XDDVT0];;+VX[:3FZE_8G8
)P37FMfW#Z72N4[Z0FfV3<e&_d/763ZLdMZ]J7bM_fEJ@-d=cVLFReP>HH,)41=-
a8WM<dAY6EXCb.F.#Bc/(Da)Q^-A1?S/C,4S:--<f(^,-9SL6/P=LH)^_\VXJQ1b
B/^b^V[J\fR&6\OJFJ,gU^.eN;@X4IXa6,d^JG4:?BYON&SQA1)a2,E>;M1E3CdO
H><fg^K0GMBCMJB&F^eMV0&]6--=:RYR1?(M+PW?X5VHbcK3)gG8L#5TaUfEUZVR
2&MOIY6/I2>]DG&V+J48JRL0RR7d,a[E)=^<F[5@d6)agYc)A_Fe<:6ZRHA01b1,
6fJC,X[EUK30HP+W5)=.BD];182/_?QI7d8K:^8H&:DJ;D_<6XLT:,d-[RRVca&(
.a/+L).eUf>Z:R5+&<YVGET)/(7X8F9/V7?(+g1\\/A:WA10U]gc?MJe51V.X\fF
2aeS.EJC/)S)N-(S6TOM5584XcA7RbWKa,f9KE-d0Y?YMXS-9K\/=7/]FX.YC^^Y
PJ8RfJ;R(RA7=9(DE&31,dR[2]=bFTW\XfJ11MJ@Q_EX.0O2JFCEVE<&gYCH3X,5
/.KO7bCacd@BR_NaCL^6f7].13V^HGX3fD;__[IGe)LN0JHe3>&RAI>/[]85Va&7
BGVIXQ5\+,d@e-0daUJAX,E6YDP/.b[aC((O,a](<.)HY@BJ-a_gHET85MeJg,/I
RSMUWR;TL/eX)97EO=7-6<)HTE8(8\+-Z_F&NC2EO/ad/P3KE<W.K[:6c-QB;-88
Z\4<6GFJ_L^Y8)KP0M/eUN2,3M8BW?^7<AZ]/)^\ARS]<g]e4CbCIRWEVWA<X(A[
VQSJ4a[-_V(8.]Y^5IRTEJafHU_@T44?)+3CZ;2C,-fJNRO6J/3#C76K\A]UZ-);
YN6VC/OM7SX&->B8[QN&RKLS9]IQIMa3V9YMZE/@UL&\5UJA8R?aB#c+WK0A3)>:
^&[<+0^6A&UIVe(-Bbg(eB=NeRHWAaI4;]c8@SAF=7UV&:BVYg6-1;.d4L]e@RO=
X:7=ALN&=)KEHR5Q0ZS>@_cCPLa&ba^.X_Z:J\?_:;g(=4O;W^-IZ17Ge7eeF]BD
?eRV_98W3K_)9e8+Pg,B.U<-fS\d3TU<4T=24A_J+SDYP3=J=_PSAdK3K68F.KZ.
f4QP?FCR8E4AgUb=.E7Hb33E+\7OSVAaYd-WZLZ5,KPZR3+R30cW.de@e+/79=.(
VcXG=>-dJQ(<2ae;Y,a+V1,>,7_(7;PZ+(afA,+4O3AM/eA&KeGSJ0GJ],W/U,#6
D(:Q<&85c+0H=8MXP:a5L\S,_5ac]YeJ2PII[HW=bY]23I9+OLeRP)U)^>:b.EQB
#YO+9&WXV]V\TF@eSU6X#Y);=O=^VUXNZ,N]MRE.c=>XVH]7<gWcH/J7B5:7HU&V
HGVb3#AgK5CFAdb2-5-d[3eD5W4FYWHHOJc?c,U7=@H7A_-c)8:#8P9eE_MVgC)S
J/8#(Sg8HUHEG_<3gL#^6OG8:RP4Pe4V_\+2-</R/:56]I\Y@EdWb3/(@]U4cZF#
@441R1J.d4fNOEJ:?H1_eU?Z1S;Kb<+WCZ1:G>CU(MX.R(XZ=I5g^>LA[(_<JKgb
,I#[9-Xdg;PcDO0:ZOI02Y.F6b67=M/[BF?@R@NT?M,\I-c[]LOHW:EP1CFJ\QZB
NNHJ5WT-^W@;/]NH,MJUC0ULG]=GaXN7>R\QfgA(#]S-&Ge^Q/UO,XX>[aIgN>R2
)@IQA]_2GcG-\>]baDYeTa61@4#_)=<_HCP5fM,-8U@Sgf@TdJP)W8EbCO(T>.,+
)0,@WN@<O2^FJY_)Y_8\^YU.;8BeUO2f7]N/3/ADV>SgXW7Ze@/Vd,U6IKdEWJV#
^&\B:.A^9U9JORg003:GY3A:OA#T1eaUVS0@0dE\K)g#46EbNJ6E9B_:AaIL^S?a
BW2;eBJ[B0]\O,C_NU#P@bc\\X1V-C^6\&VG?OBc;-]Y9d=@9g9A)-C<7=YagF.^
ZGO>,U_+V_=eSeTBFceJLf;6<1=d+>?GYB2&CFK(6bdYC<NP1K@;^N^;4..V/S#C
,-].)Y4VZfIBL<(Q<dS?LAO1^M0c>FLC#e6?=.-\#.J\46M&^UX/9[dQ:=]8QH07
c:/S7?M8Y=^ZP+E@WF0@<G7#2]0W3X77G9T3-MPX;aY-e6K#E4SRC)7W,5)B:()#
6_daRd&+d5HC9Q@=XcHd)QWCNPP:1Ze[e]8#b)[4\e.>,:EJ_+PeR8OEHD>WG9O]
09J@c,6X<V<:S96A3?V9&F#+.7\8d&<>3#UET[Rf[#M(P,V8P@-OaUd]dE5;e\8a
1YeF/N,61OQ^819ag<5:QBgE/ad/Y<)C1_Z1PD.3XF4F;5FFR(Tb0W9f_O_/1,<?
3MY3@d1F;8[Dd.EWWK]IKEZ/,dTZgZY#0RBW<(D=)X.&d^cg;NGGA6IUa#b^/\O?
c)N,89LWG1>0<([&G=VRW4;P];DL_aD)LcB]W@L1:21:2SR^-7+>K?J1aMAIJ8JF
c\CV[D)6@:.=M+NaUA]:D/MFJ/VSL3S#<1g#+E8XK8CH@c)E=?7OBPL@Sg=953BT
B0Qeb3@397aFS.;WEQT+.PA(TH-](G8Z1RK?P1>fQ:A75ca;Ug(V9Q5NU(X,^WMU
-^3YgDJQZ,]X:)N@YMI3WK^Cf5==>;3EHS[>8\?WDf?P5&/Y.2G7H(>dJG86C[@X
-=P&US#M5T6/S+cLgH,]edf>?a^49\H#)4ENE<(VM3+QOKVM#AGd2E/.DIL+B?)A
Y8+Wfg\3A@>R),D\Y7O,5X7RA<##+/&]N-eYS&S:E54ME1E^f=)EHT=@[[bTE6Fb
8;6a/R).?QN?PFPF+,c#:)#FMY9@7N[??4R=?RORK-HJR](]8gEbE6?#K<3072:X
CZS;>F>&d:e&62cKW>8#A@L.6Wa3^S-E;-cG^V/#3ab\ePW9<Gd7;S/_CGf96:\X
GJa95-Q2Z:NZ(^S@I;6=eKe.DQ_T6AgD4?BG(P<^C#=fg=0+SgEK64UPdC(VSN9?
g=d<IQ]Xe[L>TNYSOLD6ZU#cR[Y7B[\B9(>gEAV:PNaKec5S=>Z\<#&,/&GS5IfL
[7Fb#A^CDUB7Tb:ZbKA=P>dA963,Hc?(:P[,b-QdM9a1ZJ)L-2f]XLgd7W9-dZ#O
eY,E;)c7AT2_eOA:g4LTf@Y_14787UEb4:RQ\@LS@Xc)_,.H2d,R[[4]G9c\P)YW
I]:Y[@0b=9RAC6@;KaO.b[J>F0EQI:(c;Z6E7C#1Ig^eRR,/]YH@O])QN8<(+6X1
6KbPW<BB[0]X6d4@dZ4X/\QY^8MbN3O8]Vec49I3Z/C^]5UVD_BVODHK)<OLKSPP
Z?+U)88cbAbYH>3S>AIS1O6>#Y:(DH7c\QNP;eDF6R[;FAS@Y:-/5.YT4JVJ^VTV
[J-&1]5H(KUc4C4a)e@=WVa&;;;U&@e+]0S6MRY5g./OM(WXZ&;FR(_Vd(8PVQ2R
d9^57d.AeI5Ba9_21^8F/#5W.#>[DQdW1fZ-OD?B+KO,A=#9X03/W1WC_#QVdB0E
X-F8C#>@6I3A:JV5-SB2)fYUFSPPf.Hb>OGJ5\g^4;D>I^[0S0c\&G;9_KS\)J]T
\Q2_;R7^1YH_P6c,?0:.EWa:87ODEMGg/@1=\;bP<+MP.JC?X(I8VMKU5IcVEe@@
gd]FHVc/?@b8LTW]g=NDJOSO<\+Lb._fTc)B3aR#5YV_I=34B[dDc]/7c=@N?Q6R
8J^A(XgTKfY]43Le@QLVI&_UL_IK#:Z_J+JY8,>0-#.4,HR\+/;H(.61K#g_C@-;
TFBN4bUfH2fFe[RGPP2]6@.\M,8C@5,e:3,WZL#O^^CgKAKD_C>QbIf#],SQTJ5N
Y<#=S/V^/,\Q2R]JTW3+^D+V6[c&VEbM#Q2bKYKU-,W:629>U9Le1V/75BA_.E;b
J<g<P=Gd.MCY<VF_<1a/\RcgZSKcXD>fS8\=<)<<RT5&,M>X^(@cVEbaG&5G,GT9
8>#(,fg+?-A6ZFId.1dZc(bZKIB_cV;aGY_0U+gec;gZCEVc;c0S+JGCN[dIQW3P
U;R^,L5XG-XX\]R:a>CP:WY,GCJ,3g&NH34DW@-eB\733X83=TA94WS;\=/eP(DQ
[E@HQ<R,:>BHJR\FQY8]^6aT[Kc2LVDWJ70?>#>]MdXCI5^P)MAG)#e]=,fg9Ice
]VB&&R=ZH9^>L57V.?,.^;YO0)CMG&>/V[.6+9\[R^5DgT[5&5#9SQcg_Q,UT(dX
<?ecK7M^)]6BHFc5[49@R8VWFDP-&8O??c?A3Ef-+-KR+7MYZ=bU&H=O+Z<GSgc#
?NSFdgQc365]MdAeARcVGF18=&IHS6VGf[PF?U/@]WFe[+;@b>BM/<K4F1A/EH2b
;O[C1J3S\3Q[>5?O2dZRg\g-#QA06f<F8aKAd3L(6C84HU;PZQ.1FJR6F\4>1X7R
F@PgL3+#?X.T6]@OVAJN#M6AX&.dPQa<HC=ONbcD-Qe&H+8UbCM3)\6Dbcdf(SXR
,\&c;EcK1&\O\2bF23MO:VF](.K42[A).UE?3AXc9#&9<KIK8c>;TeCMJ+XCD73;
XZ-F<>a4&[D==9&g#B&,9f/6;C;Lc;9U@gW/:0[e^EZ/bSCHX3I.&;fK6\,)H-_9
/#];/(E\2F^/)d9QB\9I-JO4CDC(T(0fSVUO=_W7B7,26+I/YDgYXEPWW)Xa((fR
-^(N0W-6106LP;ABT;a@>W:Qb<Cf6bcLP>OXEE-5^2H/e(;(QfQ;c;Ig:-UU<80H
SD<Ne\&R,bQ]cg-YVg-+f&7aX_b870)V]5?[1J1:&M.[E2Z_SSDV.-BXT20GKfCN
(+IY.R<I#4<KB_,I]98de&8@a^0RH_DfGUZ4EZ=LM&eLg-:3)f\51,VL7IU4A?A7
^6-#+F<6+\HDN(]JJTRB;E_#&^ICg[Qce=:O\:\>_J&?BGFNVU7Z7c3<\8=7V)D^
Te/?]g-b30O3?eZ,c)Qc:.C.+dOQM7R+YZ#D@?#dMY7P4N[/4P40OZ1IS@P)8;C-
[Z;NN98;g@R0V7WCf1]G-3bXacY[HDe591Y)>J9@(Q-)]GP\g6@IeJ-;g3e8Y,&O
+:dXT-fU[d@DcQ\[]dWd\:c2LPe/L^,4PVS;9/aeAOK&=4A=5\0#NRNE9FYdE7]F
31\<C2RDIQM#d2f+EEUbG8BX<4:f?Q?W0N@)S0/>UEG&fZ@C4)Ge]08+-.HVOP-A
R]Kf&^Y\:8V>./-JDF.7aR[(^214C@cf-DI7\RSD7+(2B34Z2TW/E]BQHMGISFa[
^>6(gR)9_a+Ef?Q#X0JM]59;+MT,S.ZQgMGeD0TJ:OV228-GI?^##dEfB6P6S6Se
@R:+WX?AV0POQQY],f@f6@M2U:6V/8J-NGK\d8]Bd+RDfD,B&^@D7#R(9CcJ/VNK
[\E7Ke.=(_aH-7c@JBcI2-e9VUMRG8:I#I5PE&N+X].YOL-TR0_7_[S>X&#>.ZN9
=)=ZaOP<L)HdB00X(?_\;A__[;eU_SQF+.MG^GFS)SPQF7,aC:42QLOfb8Z#2-[A
-XF2D(W]dc=276RW&N)VE)-=HOf0CZg=gCCI^>4A#9O.CdDNW]c,5OAZ3RC[)I0W
.OK)CSgMG7K3bS(AJR-X?<T>A5OR@f(>U-OL#_g,J,(bMAH[@&8Cg:/B0+a/:0eL
-,X6S.IO:\(]Dd:PPR:<#0I?Vb[[a_IO?W^=;a=40&]CD0+E(faIT.cISQWFM70L
a1D5Q@Q7-fH5aCKWIY(B]HMJ3]51<K^FFW1U;bX6^G^=8b_QX@-f9,[d-LB&P@/^
CXe324?c(I:d<7F957?[=H(W)X+7;7M9Gf?G8[;I8&ED_42bS\5L,VK?dbbAd/B_
Y[QK@?CN@M>U.<)O/O^M&?cc?79XR-A?S.0,4S)^aT<MFR[bdRIBa>:B1\=R5U8c
^(D-3&(g7O-fcSV:b=,9/DAC3X<b^CY&RF_cONQCB9U\[b\/<98G/_0-gYfUc>Vb
)^:?cCEa/aMLDQQTA6dX.4GDML=7/UgV(RS9N_R<eg44HT2BHL7OLSdVC9RJS]T4
+C\IJ)AKE(,JI<+E8S>S2?1:/K^TN:Q3BFVPa<:UgJ]@_]0#=\2^5ZF]3:f880F<
\O_2=c(Kf_\3FBY_QPb>489eILgD2K)TOf_1d7Z0)JKYa<B0O3AN,.C.L?a3B+>;
GScYcWc-R,RMQ:2,ddf[?.)D4BgfQZ8C:,T6Qg4DMHBS(XOLb<e7PEU9X)IJFVKV
R>(dXg2]\d3.^dE8J)T1fA+TI_77)DJ7#_&e[W,OZ@(f]^T:4T2cd[EIab1fTZc5
;KEea4?/S)72Va^(<Ybc0Lcgd<dW>3F?[g6eJI6]AYb/(_N,VL77M293;&_85C>W
R#VPeZ@N\(f\&9E4A985:_Mab#9P)D,24637NW)bWS9=EXf(<<Zeg]W7/C_@\4EG
Sf4DRD4Z\P45=a:bGR(BD.-L?G.<--T2A?>4CGNQE7]PY9.@0fM4N]O9FY<DGCV9
\A24e<NNa0A[S^A>=NFFD4FUg0ca[V(KBZXYQ=1WdC=QJH/R[Q7IE:?54(1KJ[<B
>C#,5.DVE9eB#U1P+1[fMag3;].@EbcZgB;?QOJD/]De&?G1SD3cB/a\1FLY1/RH
^>_A2D?g\4Fc@a+&C;6T,F9IE>U96LW.V\H<SUO0)@K53REGDIV58#]W.b>dS,IQ
>63JDUO_WC6gE24=9TR^\U0H^Y=dQY_1NDd][=#=E57X=J+4)eW&Z.,A&S52H+ZO
fMZH=_>WMgYYTE0U<+DR9UI#W[O^ALe9Z=<a&WRW[O.T<]MCGQK?Ig6Y3[<XNQ=)
D54M2B^3+IaX=a-P[M^K01P[9:e]2[SCcJgBHT;Td3RKV]YfVd(\/@8g>(&3Xc/2
/\V/a@)0V<4-Y1=<W_UUXZM,8(+aAVX=Bcg.8]Z-^Z:-F\,2/Qf/B01aSY92W;d0
(#+2@d]GFTRg&)4gUYf,I^H27?X6U6OZ.)Ja#H>[T(4fUG:K0_0U9M=O#_fA07&[
:LWT-XW>SO->G,NFW\@SAW/L>O#WMb@96gB,QZ./35&9=]78.Od&8)d,X^N#O5:A
Rg[@cXY,U^R9@TE@T4D-6@bX)S(@],Ne8TH(QUT;f]_VcSg[27c^/de]?S0b;8[B
,<,1?4g7;6XW0VAA>I5^L@//]EDFO.+G9+cc/eQ\&,W3J+>Ua9M@+_?P(>c6ZYRM
,gc^VJ#_(,,230&R@E@_)-#dU8.1fUE@MKa(G-@^5W,H]bC\P_LV^=?7g<=H&C4/
T7eP1ZedI3?,@Ebe-_S>>=Ga#Ka[NcHf466F&@Xb;TcVIbK7C=0,a.4CBXK;(C)d
B(SLCb66\/J49f\T[)C09-LBR)cM)7R>W,Qd^:K4JScC:a#QKRUTD<J8&NcC+BI;
\0fLG,dXU44/d[[9>VL,1?;NW88IB)M.9e:P;REJ/DK,g7AeA#b<aZK/L#A_&CVY
6IL?1+5\UY7HVPTe?@Q]HXI^d;4NF+@LG(JCf1S1B&WW/6>64D(/E=E8J#WY253T
C<0JU-7?2J\9IERX[PN,Ug#bST4X?cY;E_UB8Jf-;)@ST2CWd0CJWB+J]7+R(S6G
:6YXU86:YTI/c<Te/EC1W3\&N.>C;8?/X,A]f@+?0-MY@M+PK)EdIEC<[OW4XHQQ
,XRU4>g+e]SKEHdAb^S0c_+X2;^E168/2afI-&>4S&OAa&d6LL:JHE#B\LHF,9)[
IL<2Y\@fXR1NFO,610M\FAIf-BD7V4ePCD#&78c:0P(C3C2(EK9AN@0<^EDKC>SL
2/@)Y)<+DTE0N=TC<H;V6HfJ@I^3HZ&f9V_fLBYI;BFYRP.@Y>/d7-</-M5g)fg0
8R,@.,YeT-RGF/[fVPT#K18;7Yg.I<L;ZMQ;QCOVK4K26Ic0&2gR[cF-,[6[6A;J
BfYI?437gHI5S3S.+Db>2L^9,LQE7Z-OQIHXZHY]d]GO;FIN.9<R<5S@M.8AEUg0
I]BCY8],Te/eH=c/-J)BPA6J-SV-3-6=P_(.H[#;K]P1Q:]a_1F8<;(GAB)(Z\:d
&GS+82?1X&^[b/FY(W)JJB<3F-X<CBG8de]d6=_FW8#OUP:)9A+B,[Fe]R5EMCc@
A@ONY1DC5Y&V]U/P1A=3/[79L]>,Nb5_?gL_N.KWQSEfCbARcF?b.T3:+J]GYKC\
ON&1T.CKQb<gZ2H6;^>O7HC&_b+=@Z]gc/+XL\9=D8]<([16M,MGELd@C_NB7[eU
(A:LED]-a;?f9W\+fa_1C545,)OTbXBDf_IZDe[3EP]D#Q0[YX^fK?J[CY2eS99e
:S:42E<+cMZB9=;b4)RAe(U#;<4^5cd\E_=Z(J/RW^418\33MSE/6-RW):Ee,>VI
EK=REYGKBX.IcW01<b2XJ,>WfLe7WBDL&S5,)2dIJSJ4[c[]gC3X)J^A;L81e#N4
6e#CQJ-8HQUMQ^@-:6a87[5bC[NVBH)P@X8A612P.^]UNPLCUBK/5)d_K,RWOO]/
fIE,IQWD^>I5e@;REaAXQJ]6GI&F.5US9VH4g0GWYd2OC#BU)9,c)Qf,0\^ZJe03
VQYc=:;5A7g2BO#]5[[=XB=DZNaD[,YLa>,-D@-IbZ6ARGTJ61Ke#7^14d;GE=2A
&.]9aM[V#]c8:KF3>W1Z4N=K05>@Z\g.K=P<TB6X)DdN_6]+;W<\7FZZ)R67Sc2S
cT(2Y0I-TUL^U6+(_F<7EOZ[&TR+-b_0MP5Zb&JR=U[:&=3d5.4/=;]KMf92a;TF
Xa8R/SB&YF,OF<MP)]L2&Zb-/MX+Wb/>d[gGEU8(SBI(FQ;HBOg?:C)6[EMCJ999
UQ77QXSLM+=4a;G@;IY0W>XZ._^-bTgPUWIL\+?>?_0b,EgP[J,WMdg5Qe/fVafP
=]W3+JO1C/VJ2D9G/S#bf?4Q[6P=FdFgLN6KggVA:7Y9M1\/NA_U7[CC6>M(cG0/
^Z2#dFVRa;S&UQNDB98@=DBKA/I70A;6FC>)H4/bZ@]GAcb)UDGBe)969D76MBLM
9gV=@)I3X9[N4Kc+[TXW,E5[/b,UIE_>g_IDW^_\FF&Qg84W37Bd9GTY^1/;XUEb
=VWBIbBBS3,IC3^BcHAb+ZW1#9)/&N&SL4PWI@,-RN]-V>eB5+X=)X_PNWUPQZ^.
05V2FbO>:LFe@T)IUKI/\D?S<f_D2.Z-ZaYJ4T]P?G6_2)KF2[]3A;87Ed.4d(XP
,0<PU<&NGdOFH20:B>eK2QfeVg3A<&./.=VV=XeZ#DXc9H5TT>](RZ.ATPcH_a).
EggY=6_&^AI><(C0(80=8]c^2JFSJGA3c>5@Xf]Q]Of[3N([a9IZ:CX1=W+4XT\<
+1SE<U8Mf]=30-QD4]FM/88ZQ<g-cK5fQ.E^9Q4D_&R(-?E]]c;9]a204:_5S9bD
U?_U1bLN(T2FQUQec\+(.A.)d.2VZeHBE:USgBGG5:\)U?_=J3@a+<Fb-TB/M&@U
47;Lad;R_[@4[)f^d,W(?>8D:=QZ,3)M;<<+];U]D[U0>B4@EMO2G#L#X8V1:fJ>
5?&FcPE],D+d,<@7)Mc1UK[G;;2B(.dA-3XE)@:a6;E2B@B&KIC<B[U(e9Cg;cSB
VR_d@^aHA\N5#;QgU)f;VG<47TTEV;\QQ^TH_6S#V:EfPfZ>O?f<O#W,\Q)-cdM9
F2>1TPC,AfV+_VI4Lc(QCEd(Z28E+/K)LVR,d]^f&N&T#L8K#8YUL+9&gf&6]bJf
2K6A=,&/CI6L)a0O?UQfAZ?(BMTg.(/.XM_D:6.=2;(WFe&\/Gd9P#c:PR5QW)1O
D4,B2;J;_FaE/;DCf,;gGB]U+ZL+d:YI#?#PYXO7dNg9:GZIF<7IAP;),Ye#7Q6B
86+bYFK3T8;b@<H<I(Ff&N@\^bNdb[4Z@JabcAQ(IIGTKEDM:Q9(<2ePM1NC#+9W
T/XKH;4?ZKVJR@?<)5-=fHAb]=d7[,YAL-)a-&0VJe/Dc]dY-Ke:)a&VPA3T;7/4
gA?N1Y]ENeZ9QU6g)E=@Pd\>NF(@.]1:FaY,d[EaUN\\,VCHYc@,&[CDSZQJPE@[
FKN.K7W0OWb3CVcOc-H9I3VX?753LQ:?OcJK8?H]SOBd&9&=Xf&d?RKDOg;6&&1=
gc[#2J]dCGKa\HW[4a1UF7DS70.PE;-M&[QR0V:GfP7)SK3dU[0GM\f3B--TA\I^
.K6bT(VT88)4/5<:A5J0Q8W=Ma87+6CWY\2;]1<M2F[P81=UOY\+Q/&PCY&TKQ=Z
Ld5X]IIea12(]:FbYUH&c<6a.NJF16J)5NCX?UH#Z+_&RfJ(.W&>B^A(K?+0B5G_
KOcbI:YO[a/;b97O#Na-XQY)[M^7_0RO)]LM)>edCVGL.,F#1Qc@N[E-#[&L<a4O
7@;.18;Y-NX)fFII.X/a^C&Y8(Xc<;/?F0SD&V>>B61&X:4AP6Z0DG0g:>bAK7-(
U1[]FgK6Mc,Jg1[Z)>\_deBK@e[:K#gJU0D<OZ<XU[<daJ.;2HDfAO5c7N?QdC?5
Wg]T.]eGe6MeD++f4&cP,cT#&^A4)Q#4PO+++RfGfcZ]YfPVe>D7H6Q>A@(c7\^\
Y=W6B#Td<O6F.]WeOgg,(TUQAG):X2>X(a6Fe-AU,QI_FWZ>Q>AB_I3CMLQ>,V0T
7IXP,O,d+XV;RS((HH@gQ(I(74S=c[+W9F]/LHXFINON/6RICIJM^/eQf6PVPI^f
&8&+VE+2ZdV^.Eg2;_#)bNb)ILaX^_d[.?)\S11.1fG?aQT\0K:U,Z;NRP^N#V6U
BF.4C-H/ZW4L-]9K@3&1[T@fJN?DcD\:]f/5Hc\IC53I_K1)8H:+0Q4L3d(#ONL.
MB<=^g:+O9eIU:X5=SP-:Oc@])cL4XKV\0I>1,-a:J86T31@8:eR,SX3:E38ZN+,
,\LT5;0MMAg8]>T3?=4^f.KV61Y>_#^4eg?)+K+bOF/bPGW#7BYD)4?QM@JW<R:-
NNLReB)UfS^eW_cgS33A6TD<c]C-8BHaV#AQ#e8eNP:6TSY_9J8fbZZMg_^C]U#G
@XMa<2C_1a0cG]_:ZTT+?gTXH]=4MH[E7O6=E2OH?)cLK@YSA#+>=\F9\@Qg0UU.
#QCN__317eAa_adB1]9QUaLLOO]LE73Ic?/3Zgd+6aG6@0fN@M)J/OeC#/?T,?,V
/Q\#Ic29::b8f49-B3JM])J;),_;1^;Tae.+0<1E:g_9cZ<0PE#1[-gK1+X6)<SX
51^IE.VQc[ab@3c8e/-,ccQ:ETW6QR^aGQQ\9_I1NM;,GQFTYL=A]4Hf<)@W)^N9
_):,@W3^Ae&7>FEAPabAO1G60@N0,;W791Z6U6]c9J05Af7.,I<EZ;8;.6dH,X(U
H)6b&;09bT#b?1&AAPO/V+\9d1f#GUM]gDEAYeEE(#2F,U>6:Ifg:9@20gA]6;gK
UeW7(=O#2;a53#TbS?LK-,FAE&Q#0I>?<a3R\B/4^6NJ=]YRaf#T?.Y=CJB,-.F^
WL;U5:6fKGNEH#f61c/@E^A=?R-N7-8_gPTAWOY?aEXOT\bB,He>-eR8VK]V(g-T
e^CM&<&cW2B0eEOAB+3OI+G927e/#a<L+fG#I-9B6R_M/ac9PSM?d5&EJIId,]+,
S?CCD?H&CCeJ14(0&.LV:FG?c);MXcW]eP;WMNf[^6gEIZTb71+XDL=LYS5,(727
G/5/>Tg5;9g:.7bJWB#2\5g:G-a8e0;=>0,W?)f5C_aJ&W7R3(-RL^CN-CZPXS-;
\8Bf:cFG:THe)Z(Of,?HbX_BJ7NgZHbDPM77:ZTT&Ha&#a[+R]H@UNX<FO0?,b8Z
H3b&CMA4PA[Pag([Y9P>Q3W7e4B^YR.R^[ST0[H8cX\^/5J0\;<@W1<bMbSUKf(f
(+OV@aCX?\1BS5N-HF;2Q.gB^g_4Te>5THD;GdPI3?N(YPKY::>ZdI]1@MK3D++;
303SO<LZb>+[89F328cI1bX^Z8.aKQUL,6)FQO@>8T_a@a+QC\XW#B;TUG_bRI#6
&e2=/dR:P,51:YGc7KR>&9V@3&^MST=W2eV1X4I5c6OW>=c50Z6ZGY6/=1Wc3X,Z
9^CK]3b-(&CDc,8NY_]L&F36Z9g#_[4bP3adLLe?KcFdV(>F&R0?(LC0c.XF:0?e
=LKO+@(\Q2YCZe#KK[2fT(e0#8F(T?0NS>JNI7+V-H\SNW&LR3IVgPON^c1QdH[6
@_dfPF>\3PSO+SggGCAPBEM:4B&E:S&fS9&=RcPCR,0K5W]\I(XK]MACg/f;X@gD
WZfJ+cJ6S>e1=:gMW5[<<E&>ORP\J5<Y_IG6O(QDXGJdRHM+3Y>(JS@V[YX4DG_(
NE_F&@R3W+Ic1.6P-<VBdK1\<\FZ0Ug7TDE&]MDM7U,H70>5PS#L8+3[GI]-F_FJ
Ba=1&OK/-2^W=6(ROO@?;+=G9#La:=ARWG^H6.SL43SP3HcHb2\=Q.5XB&JgC:[d
]aA>Ng3PV+O6:EL/2I+D>dM=-[W#9[OO+E/fc?N&bP[8[^UW_S94SeX3:[aN\]&W
-I^^]93&E._K&H(YP;FJ@&AC0WIK-[IU0CN1?)KY;XRLOXW]A0UVLN90b<ZP&Rf(
Ie=e#fbeN<;-7c,bfeVa9/G3.05:D56gfZG;Gd^6E7\__UB(f.R1.&M+LN;QLc2/
8_]^dK,2F+-egT?MJ5W/MA=52M[a^d+Q-9Y+@EL?C;b_\7\a24FRP-M;bX/WC--0
XQeaN9+,55Ca7BgbeCQR6ZIBd;WDf5VG+CFQ^fS,_L>\USgLEdC_DER&U<9ZZ]C\
_3TGbWg3F6QUFPIXa31)OE(.4g[:O[aXF]fQY98Z5L^H8O[:?dGJ1T]d0O;1D>Sf
Rd9#VX1=[1@;a+cD]8ae0A^MJVM.&.(ga;Pc,V_[]?V7J7(1NA6>\,GZ6/]H1Y3-
f1@C9V@=8/&B,_2D<CW7C./<]fB@@<P.2Zf\#>=MKf5#4-5S@ITd_L38]9J>YY_E
76#R\6XS[Mb4Z2T[)a_Q53L(8^G91WV<G-4L2ECdB9_dO1_b#8CV3MRQQQ@<V(SX
U[0AFIJ(VF5?FcgG@b=aaI<37NP5=>.=D+If1QV:QR+QE;<TeNS)IfNaMXCHbeCI
EX\5&E-,D/H8:abNEf]8gBB/@X.YQ/;+2Z>WJ)OS)Ogd;?RF8_dVDH\gLbQc9Yca
LI0.#PF@\86+S2M#=cCdR-W#Fg,,D(=d>.(IK\9edLTE^;Y7[<-LF20C.2P?NFTB
8(:IR.^F+EQ<Z/QIU<U703I??M7,YQdK-6_0#XQHeW@;_R\O<;aT;3=DI6LLa(BZ
ffg8Z,9O>LR:7MPM#M][P>Y#N-O[^2#+X9\(fIFecg+<_c9?QKYVS9]^)Ff8ZL9S
1I552eC1VdbKI(;_1H5WCcL<YS53f<JVU#QEWI#PIADe5QM5H3#1L\;:8d>/J(e4
:K?(Ug;Wa1\a;/+^LM<^aY>4LJCH=1VSU]g<C(?IVSB6C\K^]T5N^TMOa=32[S#:
1^151aASOBgGPC<ZD>De-D]aI&_7g<TI-OUV)fN[Q\X^c1:ZXWgGD21TJUc<(aY6
bP6MegV,2)B=ZB2F02I[@AcB:=^OSf\cJ<,;>O13gd,:^LE^W9>D(3Y6Q9]9EUd]
&J.@F),SU>:&N+&(Z)]+MQ.6_abMRW;[+-=IdBL7G7F\(9B#=?_E/bP>@(]\J6EC
fCIHJC.]Q>3:_:_a[+KMHI\G2KdAZ(9SQFYI.8.6PR><b3YKg\BIYFH\#G(DRc?g
<G\&.,B>(N1823\H)A/R53OP(:2G..dAAO7=AE><4^(QcO6Q:UJUQbZWC;T=OPIc
5JG,[H>O&<B=4ER.J>bW?:64+,9e&Hg,e-&dN;ZIgJC4B)@DSHXE<(EQ^HR)4U(I
.91gP</CD/U2C[EEe9;HCY7V5^>7(Wc3MgV@,aG9+B03]RW2:5V<XP55b0#]5Pg;
>>TLOM3\cB?F_KC(]aYcQ((AA=COOSJZ7b]5JD^A4dP<fUg>7M&\gf?P+TOeDQ)(
@91\BcONIIHLF\6a@M5]MD3OHI6_8[+0aF@b[66,2NM\VWI4IC6=@;I-#I]g;]6+
>DKd\@g7^Q6EbaRbQKPX&#LKDgIOD[c6^4M[I<5L.=T)1/\MDE6HK8IYQ6_;>Z[-
eDD[J7<Q-Y@IL_SX)(JZ7a;77,1+7_N1X9=Z[;TI:8).YMRg\U-&Lg)R#YggT12P
-0,-YZHaVYX.=JFPGb+07>4f;1Og0Yd3QKd99SbZ?XeNW>;N4J\+;;M:U(7T^-Rg
3d?CgcH:FNaLK0G[K>[B:UC(1]V12/);[2IKW6B.F5<W#\:VW8]GVc,/Y(@TKQCf
N&a6c#X+cOSeIU5CdIFdeQ=33^CU&4GP+.f/FGU;LT:\XdNF7Fb\MF(AGJGc:[\8
BDI&+]-cC7C9dO././fT3K&D#^-UQ,X3_G=<BMGKdcA=K?,dUD38a[GUHGV>HIfH
P:L1QW&>,N[/NH\cX.9DZNd233NCcDJE#2,C)X5gbF]E8,B\dQ[]Y\FVW0U;QG8b
DL//AO4PSJTS/1<N2gH<I5S7.?89P9Ke3<DRH:4LR]c7H<(gb&7]6D>HDZg7DT(5
,J4O?d7XO;C.HC0D<BfP7B(@>3QQTJF..\200J;5CfeNbeXc@7SK3>B7H)0=LT(M
:;]^_WVAI_gd_N5X&15aa]6[\baQS5+WU(6,f^YOd5H]+1UbV4Tb[7?@QK(;ZV,O
^S]@FF1bXCeF_&?>X+OeH48#e&e1GWf1Mg<aJL9b^b\<P^KZ^d/BPD7&,INXgK+O
aNNf4T_VU5H2H2^^UfX-3#I\11_c#(_5/g22+[Q38dWI?EC7F#VC=\-8UDO@UUd1
1J_aCA8U9E(0-<gE&OSU1dT5[TUCd@;6.A_F?2AT<8,E#4]/f\TSD^WW)D@NeOfP
O&_A?Q2I4UYS.V0-1+J7M2=0M/g;YN8c@?FY3(C>?Y0e6IN;UKCMd_1\UQUWEIAD
@&(Rc67-g^79C6ZW[Z=@XP[&Y99KH,QXGYCSeD)\M;WL[a?Bg1>7-0XCJgN5cCe^
<UbM4^+O9>/O_(M.f:-F?2HJbLf)4;FQ]KKVY[T>P,L3MR7XJ_UfX.<E-G,Ae_fT
G6BN]&X-g8a=?:@LND7=9d&N^g/H1@_EQN#3W5ZbCZLV^UL@LY4aJWfcUUgD1SeF
;Se1.b87Z5I&7N@=VU+4>^GVEEF9eGcU6\L(H@T2\aKgKK(=5F0S;3CCAF8#\^X]
9LR<c)#<?BR)J_ggOA;N77\ZOZ1a_?<W+f1ABUANNAgU0#U/W35D?d(_,@P0>K_?
EV+0I<Q>+&>+]>HI&Y?X/d47I[YMfIJ3/UF=2GP(UD;#@=J4P3c[4R341VWT7Y0B
>QJ0N+GJ4TR0NX(S(>\-AgU+7[R<VHVF>A3,N>3@2R-/b5/@WbfAM^b+6ebKLT>R
?c8D44eJ1-U)=d5@&^:<_f^GJI--/AY2R[/E:3+.6#SG=8H@D@2g7@K35NTWa5&Y
:P(G/PAcZ(G7TL096KFT5ZGISTa.3[.AGM9MC<gXH0V,&Vf_(<15NbY-F6d;Ge[R
<8Q_]\>,g-e#bV2;7R+75F]X;M\+-Y&f\9O16(<<HDC0WA5f28JBMJ5)OXNH<WeX
_cg2?QUR&59(7(WO>a>.=[gJ8:gHP.Of?,EENCPQVM-SU9d;V(&-0/=&A:&6D.8Y
?O\-T-AJ(dYPH,g)_(R-<PZCJ9ZDJ#XRI9[UW95SUL\8BMW6Q:/b/.G6V50TARA&
ceG(d&8aFZRK?[U[>GaM^(-(@177bQLITYZ)4NeF,UELG4;,XL.0H(?Q=MdOFC]1
9Z3L@&2L=(6Ka_D_\Z+dPNJe8:H2gWH^1<E<CLb4SI7L5d43ZD>8Q9&,Z@J?GE\5
EBG0faR?QN<#=I96)^UL(;<)+0;5:@bUU1\@9;K?_T5UEI]fa>-;Y#b95&S1K4Q4
D:_(,U8CM(caTgeR54:d)E9cUGdKL+F3T05B#Q&?7NVU#V_U_Y7(WQSd@Tf1W[aC
C3UTF6.OP)4;L<F/K@cF()3TP/D13_.I7[6QfU.KW3+/T+5bC=C^9&Ob8,NP_(P_
Q&Jg,I7.-+CG<7IfPLAAU;@+FOZQgR0P_19+5I+)(_a\+47LRV>8g3)f[5UT@S+&
E(Ae#bL6:_>7R;;(1aU27>Q6aWYd^agBfP44Tg&.PG)&M5S#7MMI_gdR7cN<G5AC
[5(K^G9eWK4Dbd>cCC3@MCO.-25eXJ1/PFW:g+b_d]R4RW\#c8G@@2;O^IH=BS#Y
WLPgIf[OEUXC7N,SYbP8J^&1E@0S7AKX1O^)cVX]BN71FQEDNd7S(+K^=bba@&0[
dAgL[P.1<e&aA).gf=\3@D@H^^1-A+a+9CfKD-4JL<O9&:CK.b;WTJ^]_;Y#R,#c
X8>P)D6V\>&92)20aE02Y;6U\c3E>T/fOZ.R?bHGd2/8E6E<HLId??BQ;D_I4FV4
-D3[Rb8GQ</XT8f[O-/BH44AG>]HQK)RHS4SFQg,O3PS/[S.JIK;B7G/gN-ef9>/
cP-L)V7bZ25)KJEQD;4(T+5CRaJ0ZW?H9TdNe#MP._^K-CN2.9e/?X(K<XGB9eGb
]d^bI0MY9:(.6U@C],,T2]TgQG/RT,\TWD9Tbea+-C:X_TJa>:I;_3(AW#MM;Q1V
?WPU+9PQDO[:P=OJG8[WLZ0+9;[(_5&3D-aOM^C)O_?9L>&B6WJSN24L8<.HfWI:
YeW-Z5;/f?Y6TU?R^&3,S/2d1_c=(Q45^U0b3-TS&EfHW7-K1g2aJ8P_3=-L]?Cc
/P=UM0&&b>:FE\U.OS-3eDVc/\eB=U;X[[71+GDQ^gNd#RgH@ZQ/_f?M,;W_>@8-
.)CPEb0MQT</cJ;4d<d3-O<<1?4D.NLMN-QYaJE+H1I^8K<1NV8?D?6Y@Oa9IRaQ
5?<SHf(F((OC(Re_=0W[\2,34YTC@MH--K2#NHEeJJ7f/Be488/B@eQ646eFHB[[
J+cLB&TB;[;J@NA5FH(b4BDf,?C?^K9/3?20.FL0_Vb6T=J4YRGMG&-GK-6<L_&A
Y\+J-c&72DfN5c6.e+?WS41,V7V2U,[f60<193#DL85<\WZG2G<B&f;-e[DE?[[.
dD&)KFTX-24dYJ[O9/I1P4\H\?=..#NEX5P8ST^>O)0[Ug2e88-EMYd<1].[3=fB
ZF#_.IP+7d]f1Yb9Z.fJ,.3M:X(,7DS?A6JFQ//CKeJ6-c-(W6bHBT2F5W)IbA&;
UDXQN;[/2X/@-I\UfY,RC1g5TWd_,&eg5<B]YT\+b6K2a3_4@+HLTN+MWPfZKJ#H
;HP#EbCCP@=+&0H)VA+H_ULfMX+c:C6TN?H/DbG[/I2+5CJ\f?JBD.GP4YH)..KZ
9LEAF;ZKJJ+-8ZUP+a=+643U:3BNaQI,3GMd)05]a>XILZ)W(C75CY25V_ECNS(H
Q^^^1fPY+A26,JAAF]R_V[.RGa:@VWBDYdH,X?QLX4S2a\IQ0G_G6//:E@T_I<R5
6f(LZ4E?#7=&XR6X8Ja8fB?50FH6YdOY@66+POLX2(V6;WfH-N8M]J>-0(ZH4.)d
B\KZ[\ZN8Z?SD)2[-Sb,7[cbS(8,PBCZO@:KN=c[DZfCS=dGE39]NW9NBaf[\H&B
E2g^e2S)_L:;Q3^(GV/M(\6C7EHA@V(JD0U=RKK9H]E0OS+7+([(R>COQ,.EX)CG
Y)@cMJbf=TL.7WS]aX]OM?X+Rc5^JR;VS^]PX(eIU^,e[=3\Xe]M-NEO4O_OR.)5
H#9P&,T&ZH-OC_T#@)F>c0e2I=e)Y@\dE+M?H0Sa(SO-?ZT^CaNaf-+Z;a[f0cL6
1^UJB+/.XdS+dCX_\EP70K:,71<^\dcW^;L7(QPb3OD,<]Z)N;W530fFg23XC(--
>PfOM4&#6<Wga71CP#N7VU<OSc98bN,JYH2]O2L58T<:g0YX,F10fg);ZT8V:)Cd
OWX+&J.5-R^B.RQW(Ue.<<V8A_RQdBcB?0SN:/]NF#\#-3(>aDOV-:ILZ;EXM4:U
Wf9M_<>.;+(,A/XYQ@Pa7A(@7g-0ZYS3=4gTL)dg<+]d;XWQ<EQK-6TKMAXe(?US
--:;Vef8MT:W-aN:KfK0VMVJ#]=/8Q&/D#0&[TRR<&.QFNV[?Yf:S^/4FdB#KW?\
c=#P>EO0EbAC&5_C^a&<&>]B_O4?VF0Pf&ZX;(Gf4GJdL.02XCe(S;VDbC&U.4-N
IU)c>=8-F2H19.?de(8UI-NY_SUf9/F@\a:HW<P>0bg:L3]>4AaId>M-Rd2c)G?V
)/UC)YD<B0IcH\Nb,OGQ/S/-CB7e5Z-3a^P330C0<<dJcG#f^=MfO0#?]_dYPa(I
EA?VJP_a_;MOMWI:#A7Lb(TNVX\Z]4DL/4Db:)c=9Y1G\<F#-dI9&H93(4(3=3;Q
@7;6R?B./R?F3)[abZA9aR\?M;S\1>@9XSE2Vf]NeBb#&-=eZ-E#J9X]Ae<35c3+
.M&3Lc/7U[A2@SL;V\9+(<MUBS[+4=A9gJ_c&^17V&88#5,6OIea^e;19HFB+DFU
54O(7XI##?d-&R?-dWL5J([aXR66XJ=AVdLcTATR_ZT?eM1YZ#b]:X>f&S28AKB&
TA)2EW&_>4HGRRc<S?VUIEL[=)eQ-WH[><3ZUG,A_?GXC2aL7SB(fJJQU@9CIfW9
(#>V>0MUd;4S:gS:\MV5T,<A85^f=1:Oa&K],OQ>F#+E42,\CI;X-9SAMYS0_^G[
7?BQ9P[fO-0E2IY>UBE292XM3Qf7Xe?UXQfR.5#=&+4IN7U[HbQN#HQ+5UZF^N/@
ZIcg]M/^]S<.gJ9.DJ;S0VC==;CHLC5e_=^P=.dM80.URIdRN33@YB4[T125+<ZL
KTE:P231LFH#CZD,W1bQ(LTZ)CJ/ETMBSKT?Gb667/75b=A-G(/#;a734&SA<NFE
58JAgUT@Tf/F#P2)b#ZBBU[-J)P^>VDERA#;O]+c]d:4)E1cZL./e34YJ0S<8@eB
[)_fAYaQ@@+Vf&+EF-Y7aC57MHH\H)?&1g^9G88WM>W8Ca6d3_.D\0QVXTBR5&,;
,+P1g5Yf80H^47Z#dN5Feg;)3?<[Q>aeF8PW.f]e086e[U2UTQ-,GeD]@82+BY><
gU@W,3H6)c,-Y4:[KXbIC5N.3CdCF)I#X/WY<KSX?,>^I.[A:-52c:EXa1Z\5Y[)
0:\(IHJ7,c2.I1a<,/:\U-S\Q^C\6U#[_C=^W.;40K[<2EG=\@GCd3CBb1XK3\D4
104&5_.4XTGU/<)TR)8@+A,W9cFfW-UT;fT&P0WDZ@:>U/2?(adU<FSB,O1RH.bE
ZQFIKC91Uf2<g[BWg59W5f#g,RM[+VQ)bG1d<WK<@RE&488:JQHP:>I)0O6\NSV=
b8Q<6UC.CX2R2^Tg2[M/bC4>dYVSb60+/>0d8Yc+7RAV;L:&K;,U]AF.<87S&=:P
ZFaUc7GTeZPCEI=W6aBTLXc86(I@,QW39U7aC[<4(fZ8L32b8?K+.<GV9afK2:F?
a,6B-BZb?4;UCd52/.>IG_6G(27K.W+YO@8d&H0_KPZ^9Q]_S-adWI@C7QaCR6:O
56(3@PV@;3@2a+VB]-&8GaQKaJT_-E1Y]36^c258TLV#?D(K]3L]=N.#\6VPe.4:
0Wg28[4&d_<<K@XR7W,1M1](7\EgXaT0)-&H/8.-BX.OHa<M?@\<B(=Z7\=;YT_I
//[cJV0G>Q(dB)]@D/2Q(PK5)Rbg5L[;AGC:GWG-3_^Da\?H]WRV_-H-I<P,<,<4
L-K^O2D#=,AcRDD^J-68]a^[:E/c_@=PcN,M;&+(9.F@K?_L0a22f\0(?[g2?ba?
dG,Hb.:P\VfKH]&GV#\J:H>_XU_J<dUZ9I)V741/=(@Ge>/R;Z3OYJ2A+P+V(&9:
)83JR5BGP=T4E?.AR<9?ZUNd.KK?c.g)A&E,<F[S=\?:aP:D1G.O0a3<+bS=WO6R
S=O,7_bKBMaO:(?B(D(gKQ1(#IX@MPbNG0QdF_,f)eH49BK0&U176BF2YN,?=AHE
O]@cV_MFI:58aG@?7Oe@a0V]^?f17@Y_1)L6DXT[;B^9/gK>9gHI]eeXZ1[?GWSB
-^M3NaS._dI(]IF=/dBcY^&;d_c#TOd;KJ^S]XG:JR64b4]c/X5K,R.UO^Oe4RAH
:._AY3]PB\)_F#e@eN[\MH,3e#_Ve=1M3N.[a+/Pf5OD:OWaXMWZV1>;2U[4QU[)
89M\A9>RM+^7&X0?<I5gGgR(#(66J8/.d(2P1a-D,(LBa]6@b6KZf6ebP>8Z>V;6
3AVIW,I>9+?UYNeUf_,LSSaW)(D=Te-d2cEP7=e1,LR:\JZQLbF>GJF:<#5aK99K
IW&A,=eaI3BT0><>W<-(VT0e-WZ7M7-JBAOA<IX)I.^:2caSZO\+EQH0;#KGf5\-
>:YJ?#c32JbB4[cdRNU(58M2aOMA;KV=;M/@Y&:4-3(U)VNY8(6N;#6LILdWdfBZ
6Kf@;f-)+fOE1+BV[La12LGHQF_]G@K2B+@JY\:Gd.GR(cDE.38^;(bfK\@_FD/f
aE5d.fa@=5e#cF[NebeCR)4f6;CaLcO8/g6=,CVPV<+?J0>^.V?L7<R/8B#:?MRM
PS1LM.X?D+CSD4_XV4T_A?5&#3feG<1a256ONE6]N96@+6K/)/&CLHA3\W30QH4+
TT4e@DB6b<\=dH1-4c?:>4]J4A4\O^1.11A.@:QH:dV?GLR66UCfc?d108Ic3=SA
H/KOFaB]#9gIPW(AN011X5TG_99K0@dgJ1R)[5(VL,?;eW>-Id@dP<?cXEFVC;-^
WLTO#>,X>2P48>ZW5PZ_V]R0(:LB<D?U<)M3::UgCfM9[D5(\8/6^]E\UZMP^8Q,
1#-[U/1c.:F:KWXCFXH-Xd28KHaYZ2e(b\a\U8H4e-\f44BF^B7^44]d0U^R[TS8
O6636cC@F;IIa4;dR]9#66LXQ?2KB#:c(2bU2C1H5d56a97N0?55+)I+WWY45\[X
9=_47LcHDN(]XKN&?KUL-()>;>W@4X&)MZ,4b[aAHUb416,-RaG=Y6XX<\@=b9/[
a204]6/?J1M+.N(C;GW.@-\/1(8cDL]=dD@TQe]7O:ULa7S[_#K]7]FKM/O6&&IP
d/^b.N4DGG;d[\><bG0eS91N#CSP=B,0)4#)X85SB)>[=Me8<+M7XV+K79DPR8R6
V6/C1H^8ZTI\T2I=ccGgFK0LS]&T;]]G(G46)?X4c;f7X#0/Q8a;Y7>U:6WXX(d,
9HX\fH=bHgG5,)?R+NKeX\CTX8_gRa;88FC>XLf&AAVc]afFd;YgHZUEE)ZV-<YW
U(K)0eZAcB:1g:9)?eD-0OADJ&1^A#WA4&8Nc[,W@\VVROIYA+NgDdL3;U,7?#^;
W01TY&IWP)8O/IV,H5A<(H?(32D8&&9E&W9e<ba<]6]XTNc[(ZDS8PVHaM=fYX(O
MN[@)[,#X,&DCL-^.593N?:N/=K3M)WF]A_.;_V&\D2&?DSXfc9YX>d+)F4VE6XG
PF+2d((0:-eG,[^15.>^@dM[]+ZNf]RDb\2>6d,J\?/e&P[)eD;^?]5_TJY,70,B
fR=a:IMIa4>X#^;6J@NL;=aDLTFI6a+PfYVc62G_=LR/)&=(_^U510bVL6QZ_YPZ
bNOFX:<I_Z#dbG(Z+dO_P5/]X35(@+8C^L>@T_YD,JH/(BXQ3WT(DbPNK]^=<#@_
Z,SA>@.VZ/1-#f.]XN40JR9)4BPB+2]SSQ0:3;EMJU3f-[YMF2(Y6^FGcMBG;?FM
:^^^6&=_,f/He5cH3T:EHd)1HP/HT01<[F,L<T&Oe(+>3fP+G-C>+0U1Z6E<5ZfF
R6UV-&,J?2+1IUZTbFPaKeCP[eU0P4+(DMA^Mc6eNKFE]Wc6@Ef8G6\2^)0(<C#&
\F6\D77EdNYRLV2WA)dR6ED:US(^85KGgBYZGE,_GG#bW3K3S9IS.JD4[c=.gEH9
>J5^WE<@IdUf5NR).KfO&^AK.@Fe9(LEKZO]cJDY-[TU,-<2@<L26Wf#D9MXFVc^
H;OT&G0_5GE1>[=_JGRe8O1d\P;G#].E)-OXgU&96VF1#fJV)QW]PP@eDg)[0H[S
fM3V8a4.J;JX/1GfK^:R^b-1Le\F;d&H]9)bfF):@]O5UaN[F8d.:e46W,3WSF:e
)0]B_^S5C7(((O7E][H1NULBT)&8F)PTG6[@:G@dGa&&6>J&)OF^O\V8cD.cG;66
]g9H<O3(FJF,>6-LA;]\/_#cgU7JLLF/ANQDIUQ=#J<:+8JTU6^R^Q(Nb+aLQ]OI
).H1N5a=DYa2#MYML&]99#C:K?&O.&N,+R1XdWRbCKa&W/456PWABJ/Pb^YJ+P0#
4QVPW:G^5=(f8KF>.JV<CWTGaIC6[1B#:E=1(##b_L_9O.dQ@RPMP(<c?cO#8IA,
7,>K,5;LH@#ZSOVb0QE^HOLHGg)EfMD-&?/Eb0aQW;)CCXgQ\gLA#dX32/?aeB4O
g/M\[[/EM/=Z13UaV\Fa@6cUX_2(V,XVBS7?9W3S1^Le4,1E-+Qg9TLC[>9gJ0V=
b(///;]IT(XdM1R=+Ed2^aR;Z_NWD=\Y(;JIfd-U[YU_=dJV+1U+_b6CXJ?-/3B=
=P&ER>0GTSM87=SX>9T:2<I:_+=[eeTDAL)-ALdI\.PJ,EY4V2GS=4bB4fEeEHO1
(D[B.W8a]3:AZ1\ZeZ)edTZUbMQ93-H_AE9UYQD@Se?Y4X4I)>^W(Qa=<#g92XSI
e-0c0_-Fg\T^R.-RD@25?LMd9;b]G?00ZPV:[6GD8O+X.5?LX^P<>M147+.SBDca
+eF\QV(Jf2&XT23G^e1WBKC/-U4gCS.QIBUGK7.H8Ab>O.-=9R]S)@M>30_3(4&/
42@PT#JSQB-[Sa&0^.Q3)?3A,US1#G\?Z,dLGLL-/<d)E<cbGT(B(1P+T-VH8C9N
d;^cc,VUaaQD;E#]5KIME4^X/+T-B2Mgb=a(NRfd<YP<-(;OKD&D#6,f3b48HeV/
LY95(>KCKIUP(.#Kgfb,(MV2:1&<M1fBKfSAg,U8a9+Qa1ERaYU)[Se/WPT@P_?7
+VKQefaO(?GV\@S(U(#+&cgGf_8#B>B7U8:IT9[C-N:YJGUASCZXM/<S1S(+J>1V
7_a[(#g7C)0?KN<HDe(8f=.OgBZ)TOfb:Pf]2GV\>IV1?I4BR\U#/2L3Pg,C.#Y\
8;I[(baQdB>JHW]60Z08QAB8E:4O;dD/4^?DA2OJD+?1Jb,8=.11#N/3[66&Z,1I
>eS4YB\6DCa.&YA2TJM5Kg;KOO\49fLC_,46RL[K>I4PCeS/9,>2ZO9L<<Q_PMS,
Tc7P-TX6LU92:f_&6aS8cIfITdG6>OddCT6b\d\<I<=7IX+1f,aFA&T^).X:204N
<Vfc],J0KCP\H:+SaF\=7/UAG8IW&9&S<E55C(PSL30TG(AWQY+8CL0104UI@K&\
7CNC4/eZ&0gI<#C4249AFD/aX(LJ_[#@9@J/^TRa[H)T[J7?P11[Xc-g8->:D.T>
6H_LBD4FN@4GEG]S;XLY,e9;.]@gCD7\1.N=V:B.+>HPISQNF7bM97]G[\,gT.\^
f(D_SQ[51=gWWM:IKW_bX(NdC6gX[I;fDWJd8>0##\JdRfAYI(M?+?]bDD&];bP,
]9[8^?@I:JBG>\K).Y<>0,8N]CL7(#,<<:_fBZ31+agMDUY@>^L0HN4I1eD/5gg^
WI4>?,KX(:g;_-3.KCO)-8fff2VNc0BC=ETcAJcM^3]Da#A=Qg<&W-gS./(^ELW-
\/Z67#f_/4/<BXJG-_,WfJWM2IPeOUGbaPaAUA^1UBZ/14;FM^_<2d\Lg9c^g2:]
KF4F=g/8]g1=^]\)O,EE)?Z=?PDTec:<.&+<Z_T5[#EPI==76A49EM826@gK,9R5
H7VAF],-Vg0Bd(URJE80D.NM(/-\)9NZc=ab,V&76\:13S2a>EC)eYN3&0U-=]cM
C6S;.KHaLDUbUV135X.D6Q0HfZ;]:/,@A0-EO6f.0SIAPf+N8X@+0<IOI<AZ.c&2
RMI/+eE7ZGM]VI,BOF9fK7[HHd36@^g0G8<DW8M@J=8VG,ab6#@:e07cGR3]JU6?
_d35-O.RM3,9ccYa?NAG[(?@,Q/a\D=3:LVDcZ2F7A?+/M7?Q9P&?)AbDg+W=I,N
a[-87+?HTVHHS=Q(T2YM9CLY8Y39]<(NP0+KN)f1[A/C&.d/-VQB5W=-d#QH:Ge\
CYCU7_g.fHV=S/b#TFYGYO&G@M5MK(=dDN?YY21CMQZDLM+_[0SHR7dLF-_7>7RD
[1a#P\9d@f>^Me348bH#X3eTBV_KNZP;J]9;J6?59(A^I+\M&PI]ceHY3=@6_M0b
98A9eH=eVA-PM;F\#b#Z564-G+O&Q4L,I]8eGR8a(.L/f)J,#SVC[;56bU)fX-J7
.U;XY7Wad6.2F>L))91W>O(V\P1d/+Rc568LH[4K3^FREZ<T[9WRLA2?818,B]FS
_T0L5d2GZ(S/VDM4@-fN8gK5/7V>S(V&Me]Uf^[[B5;2/[&>^VX5S?a2S28>0cF>
4&8c&3aBOPg-dgab\<J&6\6CU1YP<GPN:TICWJMGQKTe?\P[AaZ5.\9MMSB;fE;+
ZXJ(.)f&HLF_-Q0c6597+WFa0f/Z)RJZ-2_e]eX4DC+PR4B#+B<U@YQSC?0EM1Z-
-eYM0+cP?7RV2,9U-;Z<K@QI)O83)QSAA=[48:&/,E(751:U8]WT?KD>6[d+S_Q-
.NK<M5b]LN4[9<dFCO8g;_A7/U6)/gNLD0SUAGVb(+C/KPQVU>(/-_F\E7\,ESJ]
C-TR&4\OLb:EeG_C7,0;J6U+N.5;E/-2W2&8\SX=VTHgCC:&4^4=W19#a>0:>7FP
Y7Z-CW;/WQ1#^_((H\DM4R&?:P(Pb/+Q2SE.QC&Mb8a/0)We@91M6T-?]e67e^XN
1T;;/GR-C)?Y(VW65CF=(#0:#\K4dG[/,[SZI3Q2(/\eI,B\CERd<<fcPWWd_Bb_
L>D4E-aO5DW./^?+b9_YVZP2@GMe8SK;OBS(D7VfU=.&SGF(I+1EGGa[@7E?KIS<
LO.S#1)-LUZ8A4_)XJ.4\C6&&Gd^>R[eGIT=0#X@gEDO<_]JV.#-QCR#R\N/-V(#
I7DfVY7c2cU2Sg0K[@cSFKE>M\V6JZB>47+)-,I:d1:B(\W0KgK^9W>[=.c_J?Z4
:_WZ0&b2FE=6L@XgP4B)_HM.1f&[HWLcUb3NW77;QC?fd.4\729<W[d(CgB<6d2B
ZCDDfW9M/SM8^bCO_)E;O/G+K[ag>FcK;)662@cO5bP_5R/=FeOR_(VP@C+0VD&>
._0)-U=b9WSdN3Y>g;]K<9=G>;]8F8;DN0F49O+>W@>c8Y4f1PG:=2])LPC>7(5d
E8H@E=GRLW8f0122Q4bGJG2^^c1Z,\6BP?C>5R_fI,53>#M4RP3X#P^EM8E>B\4Y
;;;1<Kg4=BYS,Efd50<NJ<BgCCEL#B+Z(P4MdaG?/VC?\D]84a&^MdR0cO5Qa)GD
?\S,VZ9].H#///V;]71]OH=C]a?P8@9&#7)#>K8UP&gK,MB:GXZ>H/gdAM>M_>[2
S/ANFW2a]dAeZ:Vf276W)N,@/HWUE75Rf>N^<U(b0+D6C-2?G9ZV#@cU3&#Mb]^P
&M/#c)@fC4@\<(:LW3>//=GQJP_Ma+OdXOgHO6H.b7V15)7KS1#)^,_I]86aXKE<
S>[e6=:>#a8?JO-@]P0E+I12^)<g(OUb?)a?<>PE#f--L&ZTRa,8,MF,=;K>19M#
Oc7P2V;D^JVgGAI5..eM;VUB>,YCbI_5\/I(6Mg9#&(&De\BWCE)^fOV6@Sd8R./
J87EQ7eRED0&850g]+Sb7JTWAc/L]EJPE]3@X/_/_:.gR3#J5a,PMRWbC=7X&/02
cOeTE4YF+WHfWQ.>\_E@bZULQf3;CY9b@S+A6b]T3<WK+^+8eNL9(.@=,[OUREQ_
0TfeSXZ\>OY4,=+A)<9MF@K;ee=cV25B)aNggbZfW+BW\LZYSW)I/,JM678=NT5c
YX4(\-Tdg(H_?dLJ=d@<bXeC7AW\gR2Y1TS-aZTdYb9WOd[V^)/W3UF[BD[2_V,4
]2,3fHH8TCHRSaPG:bVM0fF_K-9:EVXe&LgJ@gbVg25.=(P+LNU>O1,/)78MXUUG
;89XEfe)af2P^-bAM+_OTLfGSa;f5aK2A=D^@b)K0O#W>(a9?X^0(FAM^AE]eF)]
H:=V0R[]@HS#VF_<01I_Z;O:)<=Q@Ma<50G4\2^ZA&E-B>74^K3)YTabb\[6]JS1
-_e?7bF[#=5FAX&S@BbcQSB2bJ_DX;036bHD+cf+/Y&3M?JO&G0[6<db4=(NI8J_
CBK/cae79]KX]CC7R9.Z.gE;@>Hf_TY1OdG25;Z3G,,JZU7D=gD/&WUf@0?I3O)M
)RbIQZ;;_YWe)_EJW>E3\Q=4=T7T:?]GJ,A]=>\SD@8)C=,UXeSF6YH[5];gGfKP
F^=^?#^bS/5]VMWWIF=)#AWRP3=#3U=[^EE?&fG@@H?G;6NKAM=;A.(4B;BPM)-@
#EMd2fTX4Ge]_a:5E5R9]RQW,A.N<?O;30<3@9#)WbOO_DWNPLFED?F[[aHT1)/S
bCJ@&KZG0=VeDe5>98II3XZ-/C-QT#@A>#I0MMUUP##9->+BU(S#H#NTJ0dU^Pe:
+8aUM/(+V-=QC416MU>9YU.UP0[V0D;AR11O/a+;ZIFP.:]OV?8H5.T(2]AU;3FR
DBB;NH+06:QZ>c2^a1?cD#GAQ]?<K_RJ=a:C.Se9\-2EdF>(^>)HT)e)?:F]B(42
@(WHY2K,^=[6:HW&#PcLHT]WT8Uc.gHLXLaUPNg2ZJXPd>\a_JVaEDQ5T66G&F0?
Z5,&V(_XB]fRL@A^TVP0K[<gI+N5AG>TDO/PBH@HQ,Bd1NIQaBGSIFS)Z0eF0X+W
\aN+fbT3//QIV#Y=9a6=(5XX8bRQ6(]V#EDCde;:@9??\dHRE>SNH()P/aQ=#b\[
1aN2BF_J04MG]&)6^:,cN^g[K)[0JXM+Bf3c]b/bOLVJ9c836DW\&(+F#L;F7a1-
65:,&gULaL6[g[+efJ4U.L>g(G(JD<7@OcBK>C?(R;5V6)O:IG#@W(UWPgS4?S0H
>R+F68X_2fB\;V;7XZVS413Z;6)G+&BW:I.QOH;W>VFUa@STCG;,_OJ<KS;8#Y73
J\=MgK3RSWX275gffecC4TXNG<].D0:FO\1Le@_5fGV0f7A4_)89>EF?#8DK>NP<
J;61?A)7;IBW-BcbLNbW(,,e,Z]UQQfX7+[7^ZQC<^XHDGJ2\9)7IY@AAT-aE-4\
T9N0VP&/6cE?2g)NAXJdFSPfCOSSX8,Ze>.2ZSb\9Z#26>43JO[T;6(G6._)T;_3
?L>DW22MA0+&AXa17_5PG&TDc;;0NE7O37d7?X@&bKfU7D;?c4N>L6ae=5&M,(;M
2G<Lgf)8P7G2ZLWH;)4KES6ZU#@6XR]1Wf7J7ET>g_8II]]ZJJ;@:(Qe8=UB;4&L
D#?(Q<GQ\-d:Q[2]_&HfgZ6R#R\>3\6Y2I[MZb08fV50_;GL;NeN[I(bedVQ-beJ
_#=W>GJc.96_L-Oa37@ecaFR,@b=d99Y:,(Q;<e]46>BUAYHLEa/=+E^Z(;JU;^d
4IgdN:HNea#E6,5Af#DgT:d-,g<Wd&W6ED-eA;c+PYNVDU],LT,.5-;6JESM,HK5
>-^EMD0R_5.4U?.^dE<=2aNYdd9\/[FUJd@f4O&C0LCM=N[?Q[-0RbAN/H1)<52P
+G\4ac=QbMae3#R(XPC<T@1a2P4[?7Re[.OE/:Z?RVAM(>-b-(d+#7L1RM^V/QfW
K1e(PT4W-J61;[Q3#d&d,ZMK[^FNXB@[7>BAV<f3YWK>\I;C4g1eI/M/-MEAKPbg
J>JIg1QDPd7O&SVWAZ[a25X/NeUg&#a@Y=S#K>J9#YUE_b:1:P?10SK\U7)X5Ha)
&)I([eRS<FQ8A,8)Na=@-5^O^N7R&>F.;-5J1g5af&81MLGVU288-b=M/g-/&1;O
3B#Lf(<AOfHNF#/cE2^O23XQe^ZV^GN5M(]V=b;@=\e.^]J\H_bF1F5IFBEZaEDN
&;e@_0RH8?[Y/=7D/\aRR.[OM)G>W,R8&XBf9aWe)02:IGD+.FA]Rc63Q)MT1B8@
C]8CA/AeTefVa;Qd[9EPf^gf8&GV9LTb^fc(5#1;/C57X1B,OD^GCcR#63Q5-b]]
K3KI]4D[Q\H)-VY[1N3YfegR?9?/GX#Cg1W+Z8I@fAF\QEB7?<cN]c/-3I7,(M03
#716QP_7/-FW_@dE/UKA/g5U,#e&HD>F942aPDcLP8,A1g7aGdUaSBe)aJ_BI11)
e9IT-KaE;\9/=/@,21=A6MD1,L[[RD]X/cWE75/C(f=8\_A_P@2T,Lc,7,T)P>1T
&\553bW9(EGeXbZg=7a<X4@0f\3U&Q1@3^(1]2@CY69g3RJCOODYTK/a-D93BE7_
7f7bJ&bG:D6&+C+?5-_d:PWC0eNOZN5T</A<O89^UL#L\.Q5CR9@C988>XJJUQbf
b^DQI,ZWd_-3LW<-ZDZPYTGVTK;7_+,GI/ON-&:HEbS-FgH8[?LfCcf5OAB\Cg8A
LP_SE#15U,Z\&?cb/MgKDa+B:2UN?VHKWG.aO)3g9Kg2=19X59#-F?G-C3OM&,(U
X#/I.4JH8[\>_Z&17#XZB8:f3G9FQ<IBXTb^KX]b\cYL\#\:83(?I\:;1?JZ0.?3
VRC?af.H.QZAX8;AeK1/WXDC:9fF(7Z5L:&?2?)N_W.#7gJML9XUCL30\M,dHRfA
AEc&HECAXfCEbJe_.S7&dR5PT;5PZbVeH=@#LYeJA_5A_9f8XFIN=>>CTcC;F3D;
.VG1FfD^QSfIL=A\A89?KBR+Hb[73RGOFHYF?##80XBVJV?^?0S0[>&4G;--(#K[
0:cgEKfYF66,[=84QH9,/A=d7K3^Te.OdDLD^f5NA@(I<g_R62FT0)4FPUL;FfIO
bE+0VV(STC,;R1^.8GY0H_?7NG:^S]P)1@__gZ&Gb6gX&\T)/P>KdN4@US<J\@4-
Z:X24IQ#,VAcX#ASK>)N-g&>D8-.7@H=aV_6]37#69XI0@.c_\EH[A()7YA>_0^b
WFEI&2gF6f:-<8QKA>d@+.HQ=b#S#cP,/7/4\d4\+;L#LP3&/L(TUI4fK-O8TT&^
VSE0G=e&AZ1V;a.)P0[5)aAZ/].\/&6[8V18N..&V?][>IdO[,@3Y#e,CTJJ@I>O
R3K8gL^)20M++dH#LTa5eN;._+D4<BEMMY6=#Z@f/&1;.;EMOACDG,S^.CGVD@df
O)\#=I4d:1F;:+1>US1=cY4NQA3WC6dG,I6BC)<aQDM@g_M,?-,J&+-gdK>Z>\D4
JT]:gUZ&23:.F36VVaD3X<FYYBJa#(#F[-DPN?;6(Z1>38<@K5Y/H/c]CEH&Z,49
A\)G#5OZ0ZK?(CKE]-W3W)J-,70c[Z9VOOE]b]C3>(#XP\H;_3=e/A0?1M?a56<]
6HJ[_TPX>SZOgUHFV#Y#\ZX]\2TQ1<04T<WG\0bb@GRQ-Z<Y@cUN=-UI=QB2bE\b
:RZUcR1\2O[WO..5-(ERBW#aANZb[5#SX/7M\HC8)V-49URJ#A@I[U]W:MP;g]B^
&K3,Re1URc#d?WY)^Ef9DgDLJJWOBdf)S.DV@<)#I=f>.OD?[]E[>LFON>(,PHDf
JS+I[G+G]Fg^8HKG(FcS<[;\_-UT(;51(JM/Yb3d)+EUa2bc.BA]ATQLX177,DU^
_A=dO&6+SBADKd1LU2FAUX:;TZ1>]\HINWGX?Z=7)KS5SMPWff5K=#&S;]W+eJBJ
MN5VZc,D[,-g#GR_,4X08XQ=8RLA[.a0D+L=7&RafOf+YaReOUX.MFHc=B9_DeR.
-;G(B6[dIQW,9^F::e5OMX4T2P5#;a_g(G^MHVKM+C@LWCYKFF;HT(K0cN=7^.:]
TD1IN+E(HH]:]EJD,H)Z9e3HPC&/KRP.=)eE]_QO\6f3CM3Q0GE=\D32FF:e4;bc
D8251^dJDPGK\T0N?LVe1@&DZH<7g[D1#W3=0\&a&efIg#_]7=>,Y8:_9_fA[c;f
6T)CN6Ue#7G5T@3:YWRD4YgTGE4d^dRG;GD\7>ZP;V^Y&VUO0FYTT1daUe-O66^3
7#D:D9,]<@WIX2?aIGB,&)-@-Z0.L+8H@#EMO^:86^F8NZ?HBJ\<(dWL<OG4A48-
W4)J4VOL44(gORTN8PU0_ITRC0B9L4=M^X1UU:]g#SN&g]\&)I>V]PCVW+JgYAIb
[I,;6W4X9+,-UES0-X+=K2Q>_,P/7UW.+4#&:NUH^QZe,:Yf#Z/O9<+JZH=@]GQ]
bPCP2=MJLdCSOeMN13bF-<\^M>OW@aG8X?_,aYe>-:+dc;cY<1P89A-GeX8Pf#H3
03I@Rg34T#VcI8/g=B+Q+)S/39.Z=XE6L#Dg72_ZD\DWU(=#YF<OSD(2AbecO8BY
cO+_4Q.-KAYc71fXVQWdC+L@IR/#Nf_QR(4dR9(V+0?P)S8#4J;FDH1:d3TJ6?+X
C-._>JO0,(XRDZab6KU.@^J=dSeT:,T4Ec;PH;_VVdLUSZX7/U(d\3.-C/_V-+U9
2bI[b,5IA>bSfWVcM(@XF-9d>R^<+g_=S,ACHOHT\:[e/7&P:bLYRd?(LfgaG>85
NBd1ENcdK0SO,5_eW_36bGGG4U0\F)?6L7Y].e)MATSNf<^;RGa,Ic8+>VMEg<8C
e]aVUQ41@(AM_SE2(Te<SDe.UH5eMX#)WDZ>5dcQZ(YJY>PC]#G4&>A[=T;8bA#Q
\aNEccc6F_9LREE-2,,a4G3^cM.P#/+&ZI0@&):Q8/ULf8VW_<(8OSTFX&,b=2f-
3@aB#6X^11U=OTaXIDJGe0I>Z&>P2_MVO4=dU9>PVFUJfgO/K33YM[[NfeJJ^)22
S.MQ]M=U168/gIAa]I8BWMK:C@A:eK[2b,&85;6P;GLR,7W@b^ZdaUSOEbc;XU3C
N+R..&VX089UFDG8\,Tb70()9+\;^6[b^DZ<7^7<#,=:\1f&&dWNc7I4RI]Q7@N)
\D751][7,O-MG-c:]GeK:\5JCHSQeXF@>[^=SB<&])G[^g,.bY_)2;[T[P,.<f5f
4:<4C9aRgLX[RT;0MTT->P]]/Ua\XV[G/@H/X(Y57g0Uf67#Lb5@?Gb<S0aS@b[4
;D>T@UNK=cV=5]8K2;d2N>AO@Z:e\G_0.5fCH-^CXTaTJ[7WfT(N8&ObE9WA9WOf
(HQ(S[[/g7[d)X1.->XAI1<1(X:E9,:;FY=TPQN2cX-a()3(3GV#JF0SHW]_JFUJ
/HdB6R-GEWU2NbC.2agA>ZAO2PMBR8Z<H35gQ].Pggg,1Z1/Z^5C6R6eINb;LHVV
E])d;.d6P@F@+;Z9C]&,_]P+;(WE(eX(Z8E1]^JY6JB>Rg^-IQJ>LK7F8&[N0XVK
\A,>f@XH7-Oc-;Y-3c7]T+8,2/83>CbP\#L3J6Be0F-TCFMg<Sf?C+7RCR#eK1M5
b3[D9_e<:;,A4GDIaDZ7?;A=YK.:Cd4/Z8;65#YcLdK8CNP[g_YcO3aNRfI)3E^/
)G^#Q38^=;\F^R\IJPC5@9WMY.84JWe?[##R2,Eb;7-ZCR@6>U_:Ed?V.d8dY7VK
^gS,XB0a)&=R3R-F&@\-9g)25]\,PJ.c:U\Ea&XQ8O@V[\1-IU_3_]AR9BWfP75F
Z)^Y2^15D?,>]^6YgZ]J^B&JLM/&[_C:I??YK<N)DONT<WY00>g.?X[9ecCVd;NE
^))5/.MD3M4T^ZPKNH..bJ]6:BFH17H?V)M@(M<.WX8P::S:(eJe965,B([O>7BV
7AV(bTG8I^Q)c12[_g(2X^2&SD87-E:&HIK6N,X6+5dVbb,&fE,1I3&JdDN#WOWM
J-Y7b<4bO6O8G@ScLCfJ8D0\F&YKJAW5X+\36I(\J.LJBC#,\5QS:=Ua;I+LgUE.
^/SY]/6K\c,DU?0a]&,4LLEHFYSX5+8/-a[F;.]g7E;)S3)g+7/d@T<O&;F-bS@/
[;,MSMW/D,O&4VIP;7];d@=7+XZ@WXfD<:4(>6e=G];&(;L350]ZgR=e4:TGA(I8
PUV/M8WYSJ3Ic,E.d6,fYUC],U#_C##<^6K_CY;[,X9Q8b5W8P3Y2YOeQ;_(\.4f
Y]=W\7M;:#U_V]TQ8>AZ_ce&.K=UR?__],&9M>30?KT^[?0-?L28NXdU[ObJ,H=B
TReP-=<>#HH[,28UfM[+7N4H8058eM=EMOD9+_J(ZGL4bGR?[7VKfOU.Y[X[G9T/
)#QMLb9d>]TfA&\DK.BK1c:X9a/NDRC39QLgA+Y5c^8/-GS^><;+G1O>]3gWP+Q>
43)K6\Y0GJe^&KEdMKI+3SGMG.5;1HTJNf8MH6-R,d:<X/-[[gMNO_RAW[^K9MJe
aWZM0@O7TXF4f>_^<=(De99CY1+M^J96b.&]JGT>0UQU>bdFLBg<dI&&F8.J0JYe
d5Vc7UM409-P]+&X0c8VW([PDSLCD5T#MOaXOc5T=&fXeQ9[;DPS&,Y(VR8,QS?@
/\?[H,@GX,cO89,ac@PA3]e3/,?A77VUA=IBL<?P[<OLTK6([R97M]LGaR;B;KJQ
DT2bVCMJcc2\Ua+/DF9@d]Q3929WD/GR#Q87]1JVO/FJ]WQ#:7)C5?H.5JBCP[#g
D1L1Y4Z0;T=V6EM2[ba-PGf63d<#[gQUF):^FB.I\cE0d^<C8T_@cf;+;Pc3(^=>
O?gNO=U=KD-JII+LSOdP&X<TZG,bE-gCaISJ>T+^PW<ga^].f.0Kb/K;@e(:[eLL
K/@O?Lg=aADge.;#15T\_b0TO0eODMR?E&fEF#C6)75_Z02Z+4)6TB1#.WgN2J.0
)5gb_KZZPN=cgE#E+_0,ZJ.2YC6F6/.@a.-9ffKJT^)f5TP?bYY1E[P?GTEbfWD:
=Z^RY0SQ]B(-JA+00=gaHQ/DfVJ22W0:f\b_-3R[_&HPNAeW2U9g[8d+X7])5B,&
8K5(1S23/6aA@:Y)HGdEHHgc@5/,)-0VC-<&dEaG?-Q2O@/O<:D,V\2fQ8UACK\\
Wd7KY04=WC\KH^7^g)LOK</H\b(B15.=Sg=Qcc[TdbCI<L60J5>3:>7^/KaJf_gK
7V<MY4ET1ce_#7a2-YF#,5LNSdYOJ-_.bbM-@Sed99ZNRb(+XJ#Y]7M6)f[J4N8(
^]I;K728bI#N<#&0ANI9?KYd;:ORZ&:TWZI>^NBYB^+LcA1A55aD4,LG/g^V:HI2
3fP6gcbSUIBQ@#N:GD5?eJeISO-4;UJ0:);:[a3+c6H^eVPN:\YAHI,K5Nd2]=;O
Z9F,dP+NK<QUKb810Cf^]T7>1#\:Q&:F>/S9\)EZ#M:b>^NSDUW#E3D:?d[[((?P
)>e&/;a9FbYEF#D6LE?86=OV-58>Cbf]aF_>2#I(U(5T7EJ[04QA4:PVQ-97K_I6
V<+;CN]1Y<=,>C>LI]:c.-[.5N6Wf5Y4K>aQQ50A?RaV@@@D+(>,;Ce,0(@_b0IS
fXSbdHb6FQLW@52<7WEI5WM0XbFXAPW_<])eV(>8,_XVA;6\7=RAcCGQb+4Mf9)\
)3e8@R:/B5?ZCV:C8V-R0a)0J#E)#>CLVe9ceK91VAdL^)RI]7#<W-/;#aeD.0eV
@OU[8&AANLA]b&D&5GM-d@+T)-/SM18OJg5>;7a(O;KI8c=0S.>\W#EPd=<KN9Yg
W9NO>HR3LL<,UZbTc^(FFE-0(S/\:SRWc)-_0@2@OK7T[07)76/I7>CDEYY<aLZ(
Z5@a+QeI991a#LAE]JbW=:F1TD\Nd/I2:&:\4L63dRQY<4VVDgY4EWOXQ=HM;.=[
6@RY/Jdb1FW9N\U\R3)?Q4P?)JHM6=,/0eT3\XNF4O<CFg8_743^2e[bW_]NHWE]
<bY1;I+C?A@L&fZ/B(A:4</Z2a&9+XdTF\2B_0+eS7cZDUI(_O6;LP6[ab=>L#C5
R3XF4.2LMYLNS^(AZZ?&D\V:?_X&U0:7?gP\b:X+g\gJ5N15>7<;O<0]?Q)?B@F^
3PM6TGBG^[?B&J83N,M.>N_PDMZ7Q/W)WB9D?YWg_f>Y[fQCL2IYQ=4TW60?VZ;1
3OEgC5W3Z=Q142U-?:S7aZTab)U8ecGLW=0JD\e3T(6_^U5g&:2CeTFI:9PKARNC
OEN7eIIFC_(V0HW:CL(TM4N=ag+_#;G(=<D7=Z(-e6F6gKYd\RTE7^PB5d(S,D:;
eT)W[HS6Q+:J]<3&Q?LBMKVD5&Xdb,D(:YJQ[QZ@SeG05d;d:OI&QPJ]Zf,=GCd1
>)ZC0J,/.T7[JgfSb\=I^@LM/7]V6):,W1LDG^)Xe=75.6dMOVZK^-L4M0.EM[2Y
&I]8X;H@#19FRf7R-@d.FP+2>fQ8CDQ3^,::?KRN?WF<9]Ab32X;712#=WH4,V&>
c<@T0?;P<Z6-XX5@@O95=SBe61[U]90M++I\/3ZV8(Y-@N1/G<>V4aYH&6B(@)P=
G#dd&RD;,#;T9^--?FcSg/L+^AB5,>4fO+MOa.#G[_L<8EQQ]@-dJCY^2#^FfE\D
XZ6WAA3bBC/?J(ZW??3(]b@Jg8LLf1<V;72Z&aI53YNd(6(5V^4ee.([[dQN0(5Z
Xf^+?)-^N/afZ?TT7#c__U5[XPX0f@VSgPK3ZI92gGSHPOC>:P;Hdb7\GD44L?=K
;>]SZ62&>3LBY=C__6P/X7]XZ0/8.QXUO_7=VG^7]]g_bX_H6FYKeK(?J,&)A0[N
e:b#&KH+47Da3C]bf<3(SgQBP^FNK9A^TD^K._,Dg7HZ+>@<<^+08Z+2:fb&gc8:
MTSF?^MJFYC7+@ZbMa:X)F\6#eKReZ5SU)CZHb0JeXOSaI+;P/(eQ;Be#/gL1VSH
BV.GFZ1X9R0U_PMMgIJ1W:BaU;U00,g^0,+1WBPb-S-?ZSR,HI+bD/RUaK^a==?P
EWQ6:W2b[e+HZ3<L1T&171E;A>\T0YN@S)N-/PE2#&<A?<4Rc#EKM8Q@+=<6Z4gb
?MK+PY2?e?G4&@e(CHf_3ORU.EEV&Ed<<Cd@;]9J2C50SJ1CC.f,c&2B>7C;3UB>
?b;XAEQ-We3<-/CO30.UO&,dI2JbA5+L59J5AHQW217-V3,0e2cgd3HQECf_EaOF
>WIH&14:eY)TSD#1gPK[gU(IfZ56H[9/DaB=01LPUHJ@=T+]<TcJ3JGQT]fcZO^5
F]c9^WA+7U=8?.Z_OIcKH,NLEX);aRZ\4eOEML?fV.&HgWXFBQH?VDY,3fX5=&dT
1D5Z#\:F/^_:YIZ)_N5CLWbQ(V(C:g:LeXQ^CQC4=\KB&E-M]/Z7R<E6HD3\=b(;
K?QE=F>-[,(-c9+W_cXH,@V>XK&+a\A>dMJa4YP9^,\@[FB3MfH7P7(XM/?/ggXe
fAI(ee<gAKXO/87/F]G:U;aF5He&_HS;VT6C._J[9@<J1P0G:(&X,Q1fecb6<NH0
U:X_c94Z3#cC,KFZ7JK[g@d[Bf[/_/8KY+ZKAM<d-?EI2Y;@9eLNRPbN+MDKI/gb
_QcMbFOK#>eUV&K0:_\UFR+1[@LfE[B?bB_\f1=;B&A5K^P@7FZ-g0SL,6IgEW95
a3)[#<)>de-_CHfd]S25g#U?2&<JNcWV\Tgb-7e9fQef8D?V.6CH.aXC(5]ga_EA
(X:A.d^+cJU7L5P)FOT^I+K^B.OQdM&:/[.XbL.b4W\-@1bJ[MXKB=H[Q^S]O8VC
8H<)KQQ1\5MUB:Zd-EFE;A^R#]RLIe+6FS&A=[<IO&>2]7(AKL.?Q(]6<2eLdac,
#09^eaMR743a^S&.R[5ec.LXDY=F#+CB>8KAIfN1&E_d0-bf-FK]gEF>[>Ge<C8_
EAFVfLeb4:ZM>5C=I:-.69g>O=31^<Y?_]eH3LG?Kde26MN=b::e[&91bA_,?VXc
7/4W^4\(8=NDYX,.)83X<LSe-J=JRb,>BOHANH:AdWG3,X95d4@[E0C80:&Vf6;A
>LLP^FYcIS0N\#Kga6T+?[f21<bN?ZNg<N5>\+C.XdQ&EYg,/@RS=N_B_QH7_A0<
:8b<J(J/O3E+6><0>NbYO=FVgfZMX1G:4Z]Vb4,X=MRA)0e3OA52B7#eVaV_d[\W
8;RZ_T=\2aUG3PQ4K0BWdB0TOJ3+\3D@0F[N1/.Ma[1\I/;A>Q[d<(+4VE-<&29P
_]KH>930eF1)ULU@.,gQ\2=VYOT81=9BYf[/OQEE/PT6R)JKV5B#P2&\d7^_TS,6
f,6PH5]7E,/RIC3I(83g@;(=IU#<;-FcQ&ML/<-X0G/C-Ng>0)#<XCH4b@?(L^5<
>?Z=5J^C]@:0^VPeELZR+T)L09)73[2+VL0,^d#?Z:Kd6XC6C]AXGb#ZE?\K3SO7
VD>\fI8TTH^X/fd268:4bN6X&cF9&A/CH>#\-B,WMW@5N5D5DY?COMMIFK4/PIVU
We:QeS&>Y_7W[2IJ[E]c>I3+DDW0:/5#CI[=6@/DCD)WH94S^6:0.,O@SA^RdP,<
d@ZKe,L];CE(aE2?N+g7_]ZcfM;OOdSCSO]H>P_2,DX>^-B;N/3X7SD^[VF5:R#f
A6^6bd(Kgb&E8=E7XO=@V_>fD0D(_MN6f_HX4@NAR8g\YeC9O\UdXL=cVN#fPO?R
-UC3=HM41_1[b)PASI21+]0?@9P=(;>9ER;DaZA(>)6^HP_HHg7Sc.)^:>:G<[&V
]O+1#.P(IYV=RLOaR&)16-UNJ-E1L)-9\g:7U/9,gJY0A8OJ=<#[U28e>_-:_H57
B2PB)Cd<?\7<g/e19dY>^P07PMd)YVN-=\H7S5eJ7B]/4GWdI,e(6c<b[UO6.Hf2
;6Me,U1(eBbG6ZM<cF1UTESPHR+e4Wb;Q?2F@3LV=16OM:f17[a><I.Q=_EB9<6A
CT&G49_C@G>RK-F/F/A87)7R9^1UO)=:DdYfPg?;DIDHf/+abaBVAb(18f4Y>gZ<
UPF#3B.RIW,#7G&EU.ccB,;I;2FKQ<f9#-M\d76cD>JKGFN+KYaT=c^GN3<]<\K7
VJ2V6;Ld2GcVG&<;?T[8DAH^HdIGdK6:GAG44[TYa&KUGX-;Z?V3fJBS54@cD.<S
ILL9PWY6_X6:H=U@,QYL:0+P4,YF4SN_I&J)GY9AI_g350+g)<[^;9SWNX0/Ub(/
Hf.[YX8QfFF1c7Q\^KF;Y>Id_+KX7DA:.^W7-K(gT>b)^Ud2MKBMaMfXa#3.4@ca
P>-[-a/c]Q(=#QR[&6/J0(7gb6C&U[]2[VW/bDf=23_S9;5.>EW#U@NCUR^YeIL-
RO\Mdb2bEaa.M7XPF-(KS#&2G7+d>6PVgPf,0,ANZ.b06V7G?_,(Q:0,V<50U\+8
02NHL1E;_KE>7Pb]@Y6SBU0^a/M3-OI(>^]9#20e&0IQI/Z=.X#0NH&#_=9DPM,D
a=>=]Y/f,R_H.)_7?aE++bS1ZdW>FNBdND)6Y&IP<\d;Ua:QTZY6AS?7F\7ML,<L
c5YgR>>fJ7a/P)I/P7P)RW4-?KAY<#ALa<)9IPJbY0cL-AWY[GUB./H<K;DA--7C
EMK0e2b/3?;;PU&Qa]T3HQ&ZO(HCAZfC:1H.&fbJG_.A48d<;>=10;MG(U4f#)@O
E\YZ:R5O_6N(L?PePVfM5&2D6&L[(]EA,6>A&EK-^V:,F&XI<Y>=^\\eH^JcB\9@
P=1g+EM6+4ZS83M>9S5CDFSX0B8_@]cg51[b-c(J0WONY#M(N&D[[?,D>3#f,g:=
5F;b^2_YW_=Kca@Y5f3AeZ,U._L00C58IMaU6W-:^HB.=T#Z=Nd(,]=8.5Z92.KV
6\C9\d7,_)66O/+2DSRR4V=cAS1:^>DRY5_^:E49X+-8+1U^=;KMLUNcATD?I^<X
\9V&F.SEc?P\I@QcQeMALUd\XM9Z30@dbANO5R?dA&Hd34d&<()aaHTC3gE^B7P6
YEeO&d.7^#[J8>Ff)LKA,4VRUV;@M1FPR,#>aB0XAGL;XL4feG61Z.8,.S@(D@)1
5b5&XZM2^)KB2I6-XBF<])YVV\LD\COddg/dAIa3K)<-4T\.1aR]Z2BTKA\1AX:@
,:6H,[b_5;6#gISBd2&O34<We][.S??-EY+W2YZ<@^[RU,[O^Xd.B&;,CQXb;d1=
d48YOD/04CNCE8b?S?Y(TXK&)TESaV6LD7QV.=:NTARZ5fBgLeC&0&=3D7U&C.,L
;VIO61)JP;8R93<7NMAcN=0aC5L/L<e\HUQeFQCYgUO8C]?.^44I=#+JQ;HQ7YP@
Y_SNgK9JccdR7J5.XBUE,)48EUL(Y\-db&.1dX__46ON44<YWPQ::c674Y/9>9g+
_[eE&g1O9Sb.V#\G2;c6QS7+==+b<^:EXJ:H:GQ<#gd^[:GAY0IZU#[&6J[a,-BS
gW;S&4J/g-LX)]Y+e875(RHe\^.I>:Cd<^:;6+?#5C7K^_OW19==]e+IYJ?2N=4#
bL3@8a2b/]7)0LQZHeJFfMC8IVG4G1dT0P6-@QMMP@f97-;#^_(YRR?=,A.9R>]Y
=cdP>3<:,Yag,;P@GZOg[)@VO[D7)?YLM:ZKM4^?:?__..Wc\99Ff\Dd3].<P#<3
/4aJcBbGAU+R1L^&I--T+dJJdC33>W_\eQ-D5&KEIR5NJ.M#egfZG)Pg_;gH1Q<=
P\P0++/5DNZCNP[N+>Sd6H23[NE0XfV>cS#cbONIS@=ZbfdNXM__C?O]W[VU_V1f
74IDKW.>3/21NIEX>Q3DB-CRXP=O&#,<<C4TS<59[X+@0Ke)Y,M;#;]F0DWbW63K
SM+gWG+2@OEN8Z3X[>E9KL3KHQ[_2:]R,F]Wd>,cUD:DV<eb^-(2)/IaVQ_1edb7
^GHF^K39:\8Fe#RdK)e.QC_[MB>M>LTU.J?M3M_63>6AJLaJ5[=@6-6XR&X-aA=5
GOSJ\Mg..+<OO:bC9BR@P3WKMKJ&=J[JK)Q7[f#:QT?ZE88?B4U4)@;Bg5SLX0(A
X@RA^4f#KIR\,e\F?/Ee@T9_2WE[]<R#Uc/7TWCT1,[HM0T;ccV]R4ae;d<&e1RM
82WJc5f[.LP=G,U:.1FYRdNS@(VK#Ya&E-ELS7)^--DYb?eYWD>LU4K+-a,06gZc
E+?7?.UYAXbI1]RO/)0[1T)a>]9^AXE6+_KE:WSJK-ORg2=?#Xa7K5)/NeF;8B)8
ZMPfa0U+8g77]-N[;?ZDL9T7g,W.47F+cabA0PgAG<=7,X:NaYYFD+^V4;U/],.@
^ed]9+b@:Ma_K;fLa[W9_>W#QcH/>0;HHIdQb_BBdU1:^f&\]V\I+(Q&)T1@0=eU
g#g&HRT)3daaF30FUGRGg.+O,b;G.dKWYRH(M>&[Db?/0P9WTK/AELN\D4F[J&=4
HHZaJ@1-YgFfc9)g,WMb0AYd-W6+TA..F?TTKMD0+a5+&/306Xcb;=57OGgJY?FC
(BQI]V/RdXBSF)R&@6]MZ4eC(e/3<P3WHKFI(:L4L4JU#^d:acTVXNgD5^JXOA<&
:HYYSR.NBDMKT?J8M#0Y+_e/N=5<A/cQ.c_=WB2P?HDZfE\+5899@#@W;CK:=J]b
4TLKb<4=+B-e;5UY#YP3>15]N-N^4-M]3J:>LK]T3\+B;N95<5BVNC#J?(06UA44
?:RQL(GI]&eR+#00D#0,&^EGF^41NL^_6&C13Ea^#f]:797-L>MbLI+[4+N4)b[a
gK4JH)1L#_O[QW]ZRE6_P>[^5]GNcPAd&16E(>aX>ZNc@dLfU/Y+(N0_=[0P-0Y.
K/W89F4a/_O\Ie-AA6^58;FMJDL])44A_,WH::SQ21Z?CBd4QLELWXA#KH5^;f81
9Ce7>TC1U#,ULOc<#),=_dgfU\8/V[4-]c0,Eb1CI?>[XJ(gF.8XTeMYBN3f&e0X
Y@ARC-dK5R;\GGTH6gb(>KY970?<H-P>84K,1K5+cD/T?4HKTI.ZcSJWcS+]#FJ/
A=(Pc;SSSY[BGQ;1830SaSQ3^(J3.I9?O^.;4Y81#6)R[(K]BONFUO\Jc>f(+N/E
Y_f?7//cQL/2_T\-R6ZUW;?U;M78b]L+1WN,gHYZ._R/.=Eb(6;a3974YX:Qa:K;
@2KIWZa@90&8V4P4\/FHE^b_1\b^e>fd^0BZX)A7]fV#c+g)[DcU2067O7B0=YHB
d;f34FD204E/Q<ca8_);4eee9(@VBYE_L<4Ic0>,3CJ3<HH7B4W(3E5NcHe0P?V#
O8U5a6VIK>&dEW5R4HY<FXKc18K\Y[IOI7.D]?94,W(CC2P<]J\aNHW.UXE]J:]F
HEgJVU9I(2&CC]X7T794NA-]eA<FUfQc6I2g/\QLc3^)5;dM=I+7e^fMdb2a(^JZ
P0W_8.4)7[GR<2:\D9afFOATeO6>H61=<6N:+7WHd6O^OL/3(UAagR=(:g71^MHE
X#0&&]@T7QU)TRL\gF5aSBAf6K2EG\e#,&6?(+JWP6[dBQ=WG9ETK&gT:(:9WGcH
BZaSU7(a9Q54<>>LNg7E9_PN\aFOgVO74e3f3C^S_J?PD=G9?@T9,8ZHM==3=)>,
AEWI]>S_SW:<gg9GA[bGU;U(@CRMCRA/LGI09bb,5Z0)D-:Y.(X\W3Ae06.[cGJ(
V4O:YWWg7=bFa\CTK&3@aY<g]93.UdPBg=>,E27Z(=E>8F5^GG2#\-T9c3gKbdJP
TFJ,OYeCFYU6;.48-Y2HO/CSge&&0Z[H72D;.KdE5DT;O1KBJQ-KFRR1DfAbC\/3
,>F[XQQA4QGL24((ge^BSK72G++gCK(HE+5IM&gH<)/(a,gEY&dIVF@H5+K@?0B@
d1gQIUVZSZK@Q<Sc?UQ3S.D9b3,SDJ:-D&B+K>A?<O+d?0EaNMf^WSF??VEXKK8P
/@4cNaG:@M&gV@97\c6NBT=T-c.OF&YaEQGPN7&/47^G,\NAGT-aWPT>MHUG;?IN
bB=98N)A_2=B>=4IRH-f-ea7V6B?7?F>K:Q#UTN.gTPH/>bIZUb2F/T-B-D_?VIb
<.\K6:Ed5VN(cDO:#<9?^G:2G7\SQBXG/]@_ACS?[X>ccANQG#.(=6Xe<4Wee4PV
9;F54NZ&<96g<76aZ=[X>2DDdWFFP>MX1A\0eMg4fQDMS,O\]fO&?:UV9W]Z&BE-
H,.3VRAbd3Gga]fPZ[^Bf\L:W7>B[YQ9CDe;?0e==ETTSSI2(LddD]+7XDMBJ[^S
/c5KTU9NWd=PQ<>BSab4d3#9Cce<(8WE-_63^1IMU/e/+QHIM,N\):)YJS1DZ1eG
R3cVeWb8I8+C8>>3@.a(08<b.Fb>(WaNKLW2V.74;AZ+EVb)XE@)CMVXDPA(T]E<
ZOe<JcTA7#426adUeJ&AC0QLPR>+1R0c^YM1CSETf1LO;3.Ud]ZW_edgJGcC(_[N
:;11^.If)\22VB193A;-]e6e2#b,9P-:H>=@I\5N+X]e6:3f:Cg6:-G]+E+Y6e?5
=2U5+0AZd^S353UC_a^@D9>bS-,H.E#O>_gPAJSZ1=Le3L1d=D?_K?T;eBa_WSa^
TaNJTK96A)6WCDb?\f:3U?(^[E6+-T]+O8>5OGTSeATWX?NBX760@S-HU&eGE)Uf
bL>/7==C64X^B:a+e2FW^5,FRL?9DI9(UXG9[XPZC[fOE?W=2=/EH/YT?K\2ZGGL
d]fX)3=HG3WS=5c2.)5&EI?7dSM>ZBISNgg>M8H>74]OB].Qg+,:,,U+SU<dX<+H
3SC)&5d_5S87BR4G-G_\&;gH_@9F.?BFGQJPd-M0\,A4EPO[&G]2]B,2L;SeTJJ5
DN=U2Wf/d]:X=MC.3cbaZ>gX>Wd_b;=Kd2&gK?88<52<VJGV-=3X>M.&+E>be/_=
<E7>J3/7J;0MbFP_<)2O6TW044gRV&.K4)2;_[LX+S1@Yf#IVG;L6e=G4d@b:0dG
]JMS0:.I6gB]6DGSLe,_/e+1(9;:&0JJOM,+#<,N#7@J&;6I>GC(4d#N#2L(>;]g
6D6XU)U;M8M@T=ATY?K4gXE(=7)K7;LGcLX/8Q-4>C#@K(Vc:?A:]WC0KdSfU_D3
]da02JE-7=[@8[W[cgD.(LAEecD(_V3LC\_(?TTRJJ<W##+D=JS/0)K#c.9YWD:0
]e+BTE3;Gb@+?ecWK8A6e&WRDaGeUgVK2S:[Z-ZXf^=@8:4YX/D]\W?_@Lf-N8a-
[5(OdcV/1g2M)a:KW4+bIc-HC@QZA4=T(b7Z04-=-04BZ7\WX3AeDROKGB-TKY@-
=e0(DfIcW[daHDY79U8]SZg9f_c:De?-454/,++CU=:AW0Xdd+B#I#8e4Y^LD?U.
?E9JM+g7FDeXM?aI?05+]OY_FeFVV1a^_?:13,)M1AP\^+8Jc#TGCOJC6[QIIfH7
=>X6CCf69XS&)714SZ#V[dJUg&gd[.[=LQ]U_c0OSL5N:eG[MV:[0(5#RQ0d1e?.
5B&M\\DTe4X-#\<=#HFa:bc(;EV1d2=JG7,5a>TM;,_]K(8C=;T^()KO.S2Caa1I
9B44L?#cUX&,\XT@bX6RKaUZO6B#WX]5,Cca6D[\>ZUBQ@8RV\@/=bUEIgU.S<;=
0bc;1IC#U^J&429]D<Q_93KR39?V2NM=;6T[Yd?P34_bG2I3;8K4VS-)Lb9Ta[(S
Wa3KU<H3A.\7bY-6ED1149W+1f#BVGN\MJc^EEG0T<0c8H/#6gX[#T;.5gGB9g#M
.T[1=W2^/D,C95KUbWMBZa;O,S>VQ=>:B#BIA=;=bF4(X?5J#P7,aMM,?A902>^_
/fF[5Y?#K<Ab5&,H1>D0P+3b)53K+/;#67?@G,9.Q2;[RS8P1]5+BJ.8BCM<#33K
-3ZG+T:GTH\g/8D^<[Ha?C?MG7:3;]M9BWQbfYD.XC?>gW#H_c.@EQf3;fC3Vb4\
5[NYVXR_9T]WP3#[KT+P+1U1-K^X?M<N2GW+O\X9eSS0W1G8O6<ReX+\9GfX+P/:
VN&(1e1HgRc;-OgYTJ1<S3Ja615H,ZKV\AT^5YdIP4Y\N4+g:7JY@b,1=\a?6gWZ
g>cYXAU#P^@70^R>W6.JYK^\(/OT7N9?fcLZ4]cX5YBeD]1.#+L(;J9CT5d?>YgK
]]R<]2IVMM)PgTOI[0dZ[>M)eca(IR>AJJ)\edCf2)dHFfK9Fgd>B]UZ#K\CLY#1
c68V\JB;;@a@[TB9,8QY;^>#.=HM5+G#V#VUHS0S?EZd\AP=>71>0GC]fgEaCdRc
-5fM/FG<BA986+:N=NO\T&.KI#NQ,#U1.MY5<GaRZ7LK._eQ4,++^R&:gSQJab3B
U(GY?+(VA#eJDcf)(ecMWS\Q/2IMRHJ:\7M(640IK9>,HH\E4cV:[25>NT/&LNG[
@fH7L]DLcLL=fZfG0>1<[.NQI1Ld(FbE?/EfZAgOQU;RET?.dQ=-TQ.^>>JG0YDZ
30OCYN++AOZ8:,QW-K)(g,)QdMHMcX>XcB/4<+3g2YXM3Yc0=KFV2GGS3NKKEG,\
aL.T@ba0M.b4)Kg,d31I,gNHASRF:5;^<KI]VY;5IbP@5Q1&QCg0DF6Z4F^B.1@:
X5Za=1aXG>&2fX1@Y#JMN#f>;6,aSf0)#V@FFb/1_AbEGN5DO1@3(LM37^NEW2<8
NYHTNZG+3>cX+f@2Sb][A#gLNK1;5A-Z^Gd7?Vc56_H5[,R<-/g4G\:_UdZE.XC+
J9)]_<2]-HCG@a@Xbb?QXX@LDK\)\Sb@T3Q4GHJ+NH8\A(5YfWR;BC_ZVGI&S]XF
2VH-A0\P&93d1E2:Qa2M;.#)LQOX);Q21ea7)RL0532FTP_#0V@40NI^gXA/gKZ>
VIP8E6T2RK[CGeKRNM,5UBG;7FY&]K13:dO^#N(8^&--MV@Yc+4S<]0DR)MIJ<PP
_cV_Hge\Q1MIP7ZH1J@\.ac],b7A<L6[0Y3a]JFK4V5M/&N;e#eXc)Y]\H_VC4B^
Z;1^Id4SgG4M[_bg:L,]<8=>XD,8R\1GU_SbZ\KQ.8:]U,)_YL.&TQYGI:a]dJIR
8MJ9F]YUUO<cR:+d5dLd@4B^c+-97)?9cdgT;K\_BeT/LRMdY)R97(M&[,EUXK(a
OZ1ZO>C-)?QYZ-&^CQa<A-7H;KdT9b@_H]d(bH4Xe>@af,EAI74#>K_+/[IRWJ)[
PAW/FAF,N#ge+_#6a(TS&f^<ZJ=Z&1Q(([(KZM-#54(6/02BQagc5V-M=I7e1@;2
W3]DBA?@/MU1[,?2dSbD]ODH5aL,c9gIE1J=>T&#BB81G3a@>R@gV7^ULg?Y#YT^
0\28.PgeQ[\2E_,Ige3gI]TT\-GgMEF.B@)g<XbbJ^3>(6d3/<)N(0S.ACRC3)\3
\aQDVU@g?IN6/)_0b>gH^bE&0U2G/(SIM-^@4&e6ebB=3_,d]5>^#3&a5Ga&S)3=
\6gIN5;NT8e6d<9Sg:?+S_8+<b+\d[\Ga5MXL4O)<QL2]IX@^a0^YI#8fC>4X6b<
F+7d=B<VL1TG\]=+dDN1RX&)+b2_@5I[e82-QJF7><>TKD[UHO5XJ1G[X7_aYfZT
I//B6c^:8T>NE]HNO>D4N6b<B_MK_XL_R(//.JECC4OA,)YPO#2MDKW/O<IeW0,)
I6Z:^U]Te]Rc,c2Fg/Z5&eJ-2e5)@d-]=e9gL_01cICIa??.I/L+a)X72OEJL,4Y
[_5A#a/2B,#V@06H:eAA8F,TUM?C]GWMOe=\4W.cMNK6__</O;09.=;3fQ1V.[=e
?fOg/ZAFf[W@?Oa2O:LL,SSK-1-L_&FH1[ZL/Tf&^63&5fUd1aVLWc,3;I9B)P6_
DDE-4T5]4W4d6=1:.(X,F(OC\:@LN_>#a]5B#CA@_d_f+,IX:,>/d<??L?Ae@59U
Y5@>FP>b#[3MN>/H6(_?SEKc\FD\FAD@(()BV9JE/A99geNY;\W-(HXUNC(D_c?L
DV0H)L#^c@X^GR5E8;TQ[Z,7-P);9GBO41>1K<O[\A[J^:XcR,1>93XgQSM^13Vd
=)(^>T:_e_F27UJR^)AJL-RN7P7JRT/-<.Z/-?R?[gGSCRSI=01c73cPO;1df5YT
<8:BO.<FR)QMA>1IY+5,\/8#XFK\DgF>fB4_3+Q40H2+L,.7P7_06^R[1WS?,=Vg
E]UJOP3aP04#;9RM=PUO0F^,5[[T\\-.\W_f0N.>\^^gZR1B);U1HdU.H]B4;efW
ULIXZfQ95Hf=FHDNN3MBCDA:Y_d?39Cf^+992M73N6BC?)Ha)+X23<fB(OEQ?Fda
QYa3.KYaDPCU/4@=0(g(5@EHM4P?(K6Y^c9GE+G@VJ.JLXSD2INRc-PM3/#Sb\)U
87^.T5]=,LZFYbg;7g9.;)&P>@P1NG/.ZH->TMO2UC=KE^QNGeRJ(VGFR@f]b<5B
.:]]B#(VeE]2=F/5cH&M\(d4_:/5d&+I6H1.G&D5FL[12X5?GeUN[DAGM<=?BSGN
4FSOW/2EJ@K/(+GAc,RKV#a2Qe:0_JUA&FLO)E0c[bLM?@K&Z3/O#fA2->,<P]9C
=U\L](1(<;a7AE0H-4-OQ7,V@2+P=ZZbJf)8gTIVCY,J.^YZDY-2YXU8CeggB5+#
KX&#gLaX56gQWM@UY9Hc\@?ALOKJK<>QIIN7bNaeId+4,U[6D.K6>S,36FYUe[K;
FX]54X\+>N>dL:@R<2QTJ&K^Gb/fFU-U@PNS6c(:>(^BU8\P</E<,HHV?M]<Qb4Q
U)Nd[;0W4QRNFPE1+6[=>g+(/&CaPXd@O-.GA7P@03DK@2_d=Z8TVNeASR/H8]<g
bY-f]^fGObEc=/8HPR6MQ:_89If?]+)NKK4e5<c4^dG#JZ6V_F2M#dDD,U\RS@+=
Ic(UcA5@(?BTT,1PL.U,^fcb/B9?+[WY=8F998=IC^PF\]KVED.,EY#&4.0X^&O@
b;e40N_S(TK/dd_,g-.:.IHb7:[B2a&[A>STLEHeUL#[fBF>#aW66;Ta0#DD;R)P
O9\^b1[XM([cQ/6F#<S1J:M?-/1^:)GN4C:3D9JHM?f4U8XR<Qc>RJc]d2CVVVcU
ANHgK;gG=10)<#1[G)UeU=LMN@WG7\GS9E7J^)XdJTGT,GX+HX_@6;]8^6T2O(3f
-[E+7^-VR-BGJDE;+.R/7Uge3^3CW\5JgFOId=]LH22K;SDMQJ03S.Q\fW4[QO3I
7Hc\ZVWJZPXC#?F1bOWX6\A4b/Zd=eM_NJg/0P=GbR5EH,;.dY2Ub-@32BQ9IVbD
HaYV#WA-0)X>.]>;H-eKG.YQOaN@?WOgZ]g[=MPL9O0;5UbJ9f>52I<J1^dIGJ=<
C^A0((98&WC?VL14I-^NFJ,c0][X4\G0P5P,3.RO.&8TS_)7]I05--[M_J[aP6bP
JE;00+CH^fOHU(L\GVB-7.XMUd>d&3ZC-/Z/FbU(&&^e)M\fLJ5g[V_3TN-#N9F/
;.>e1T]F(:3,f-:Y.F(G6(CXYcL8)^VfT5(0FP@^+\/@MS)R,<]A6C[CdF\X+YLQ
>A.bBM\/G#=NJNC[Te&-ee_CX&@P^II>_M^HIK#R8BS2=dQWP7H:;G0-RN@2EEQW
/2b?&.eO9P7^9S-3+dG?WIc6<,G2NRQ^c^5IIPgHN?K#AVUb&AB(,]-GAR5b&\&D
QOL7LgRJQCP>a.d1,)RT:95[SCP;Y/_NS>f-e4E@cS:\^IN;=D\[/\bY+Y+@)Q9W
[]@>K_JW^I=01]AWD-CND&6X6PKD2ZIRPccGTI5dGLJ84L^c#;e\59Y0>SJ\,=OW
>b4LSE+92O15JJH#De[W4feW1;ed53-/>cL^K8GJ,OSUK0b&8_d0QKf,Q\d3R0KM
S4PcZ]<?]OU_d1>C]CE(\]c;W##K#1b(W>T-J:_Q)E)>9]7T2VBHc=6&I4CH1a4>
B2df#\dK:O-:ce#^O[)ESUe1V)gf<Y\21PR7\CGHFZ^@.\>;6LO;V=/BG36M&L-T
5I60HL^E8-C(=>\caMHTPG,QRPRE<.>,LH6R5>S=K,&ITA#&SU.,<H(FQADS2.U-
)@DI&2PQAC_WTIHP86#2Ya&X2IL4b404ZIPOP@_Q1KNL4<@HKXQBAS&V_\YDJcbD
?E#>VQM6EUR5EBE./,c5&U,gVUgN/H/1ZY,D@P85+CN/E;dP0[6P[cD0X726AUI^
8bJ)-O.,W&OgABdK4f<S_42LE)C8<b+<Dc=2&[CR2(I>Igc&.N?+WAT@T^c9Eb#5
,@KEJg]S;8gc+SUTMQ&7b_,R]:NK44XZ^7X&^L&Za&47=HL8[0ULD]c3.J]CW^f5
Z(]_e_feZHS#V0c):YZS6HLA\,OSI9f7Q,B6J#X;EM>eZRM=+B\8cOV/Bc2:FK=K
1,_^FP;eL&.Y<_27T1fXW4TI&d8T2FP[Y-(N#3VWM;2FL9W1;H_=Z2@YOTc0-_K1
4d4;-_G1N)^<),4:HBWVL;WecX0KTZ1cRcb04)<67=>#VXVJ4)fePe5O<OP>_IC:
6Wb<c==^[>.G-DR21VH[0GeddEC6Xb34?7F/bW^7Y^Gc0e)UZ7[(MIK=SUWcUbIJ
\3RFMWN##:d\A)d<@_&E_CDBIRTAZb9MGN2\<^TTXO@6C8/Oc6[+Z@SWG0aII-6)
1.K3E+JF+HN:1#)d4I3<gfFeC_FVH=)[_@0HYM0;=a?#LdbSFC[[^Oee.WgT+I@/
<SS)=SC)(c0[TeJDL7/2/Cd#A<g=;[S2?NK+1)0]Ad#Z>eee9JQ<?Q(MHI^5J\8W
^Pfeg#G=S+ggG2V^3A;Yd/=&85R8\,fGRYYe2<];C[D[D.[NdI-(.14Kgf=6XJ-4
?#_TL[GAGWS,6]5#FB/=6>2U>B2=6X[\E8SBG4#e8Y0AR&I5d>??g?=Cb@US,=P&
39&:e0.?eKgb,5WU#U_P:7ZeaEH.H@S)>6KCQL&??e,eP4G07gJ[/I@/>[?3(X:5
T]6F6<Lf/6GLD(bL[.#=DI[J\S3X9EIfc?.KF-FOPOS2</I##XMP_XFg_GJRM70X
EC,T?:_ZH7F^(7B9[A_g_<\LZYCI^]]I\IZ3^].IWR@Ma))CK3S&dWCJ,gY-VGYX
3E?_T:QVBa0EN)_J-cJY;Na]DS[@Wa12#TMBZEYZGgeW,4RHW4C701cGH],I4f<2
)=LN&41[>+/)[a.9[1+@[=ZY=GIbV)E3?83JXV05WJ=BK@KQ8\-;S+7eL-,Rc<GB
J>6D/;U\917XR#aaM0-D0CG?)<=X1gEF3/#dH>]><QXG)Le95Y;G>GPcbJb7GUb/
XEN2F-68([/PY5IV[9geU7[dKXU^I1+dg)VY+KEL2#TH7d.#V_eAPAR8K1dKW-MI
E<00J)2+5B2+>bC>#=0_;#J-XTV5JVY]@O]Q/-Ge?.6<S@4E;@#IfH?\[3>QZ?=_
I4>M#&6]LVS_12Kb/Z6@]f:])c>-AX3;6c(3,7ZT)69;82&E=HTT^a#75.CT+_48
0CF)W,g-#5W>1F+0<-aPNV<_BJZMY#6K</W:OE<V,d.0IJ,?/C@c.]\7YJBP+8b9
bKZX^:a=(bMFZaKLe??d&\]]IKTV.O.dB1a0@CaBa-==>POA:TMMTf+dbdZg:-7g
P/AdFO/JO6J=K_O:e<VI=VQ>V^?#4A=a^?6Fd@FG]5F4?F9FAPVMV-bX<D\<6-Y)
^@_=gdT5?6T^2/K+_H4\X/d@Z/Ad?BATX?PM]M<K^#Y+CDeRT(KI8S_VUFT\XL:-
N?6I,LB-I7VBL#d0[?fJb5Fa,S&NUbFT1,dHW_g/_,0<BOegV6f[M@0&?SQKQ3JC
DN>9fM1VRW.[:=J^AAH-c+)/P\bR_:-2O:WVf7TObGC@5A7.Cd>f,>ZgGRWBWYQ-
)=O;C2gZbcN=XAJ3:gI]Uc)BC3dN1bD0=JK@B(>9_UI\F39R0F/-gWPJ,=GKd[,?
<O3J?Cf4ZIYQa]C:/4fZ9D0R]<IUO>.S@VH/TSKcSP8W1?e;1=#A?+ebg^R1[Q7F
:F2)&?YWDRES+YB?AEXDQ7XCF^e>/)P4TB8?<E.:>0B2+]U74SYS1Y=#R&F=/5>R
-O[OXKQQ62^H)26fe]Y7)>+U?6#HM[a<eR0eSN2Wfg#AGcJC>YLAO]QKO:beEDYT
G_T:=LF#X+1FD;YeSgBJ.LU9X^MJ#EIf?FKcECP>MGHXNI&GZgEb(fVc;1Le\O+Q
.e(Kg(2dHDU/Ua>;\S=J+L<Qe?;D.B)JTY&+8I0)R8YdS9C#NgBZFJH[6TDgEIWR
-5K#Y70F+@;c\0);UgI-EZWdSZOYNDF8B=]b0>dWBD[EDN-9gQ0;38P<\2N[QD]:
HN9]V_]?I]AWWLO/W5DC4)&&TQ#G(+S,Se=4=aP>=39AF9aT5SA2_;JO4VO=CSOZ
=AV>+PW<6X]Q[1O1+#XdFTB57<(c\Xf,c_,#)8[g=R:G<B94#f^-S1^D(,>-B1#9
3T)>C_H.\gF3WNY(Z>a^1Gf9g8PQ3WF[;C(XUQBQ.bWGc\ISXNd2EG681K9:]E)Y
e^EY0KI8^gUZ=^6_F_]A5eXMZ-DE)g269_P^g[#7DfUf3[Y&7];W/]2;@C4X/99=
Z2(:_&HgRd+TKc1_TPSdPQ8ME@>b9O8BdH0_Hg._MC<RR[/FYOab6[aR72[UaIQ4
H-7S10>1Xa>b)B?)UN6864cJf,N[LP^f>.(;I-.\[_Z2>fT_S:F.[>O;[UOQb=Jd
NA36.\+=IA.UK5D@=eO8).IVWB<)c[>VY&-6e)+7IBEW4:\8FSa)GI?AUZP2U8Cg
Na=GgEJ37RSMAe0JSR;+fbNBN=ZeH6ATKaYM4Y_b+.\J.\[g#_+GL7g5FAeRZ]Bc
U.DJO@Y><#P&2aLTIJCHOMW)Id\Z,0b[@@e:(gE_P?f5AT])_ERDb9)0O4A)X]K:
a:gc[Y,=MEIb]M&e^M]A,aH2eHN\U3>,Y4D_BgPd+,Lc<?YFFU.f?80L4TC5+TH\
.9@c3=2g.?HQM+>&4(:d.TP[L9]CP==e=,,[2gD1W?Yg<_d[fM(ZD853R36T.3@f
[[_OYcfCdV_B?H@2\UIQ7&VY1a;WYVPD=gX/S>XTd8B?AR1Q^2-:-Jg1N)cB&0UE
&HEC=RB9d6[XU5;<d<?S372?D[D=X7_5egNMP9Y>405=1\HR4ZBVgSVC=(4WYK5>
eP>,(;/H8MV4APQ.W9<C0P/9468;=4aT_59&DD.c2^&W@TE\S:&4I<S]BNe&ggb?
-J(]_K2_a>3>#F77+#K(aS1C?_0cUA<0S8RDJJTa68d225A;GHLg2Q]7[:D:QQS\
bZ8U6<Q]ZS3)2UI&V4A9cNgD#ZT:YEf/WE0eeOdB\9.gFI;/2Z,f@R#CEI<@;Ca-
)9D/:OEQ>a9d<R7aP@dW;P^=b.[AKeeB5beI<cTOIWN)STKO?AO;KI^8DTSg<5U-
3^:?:R4,d4Y+;-]=\K93ROT+2WGI:dR>SM7^cfc4JQ/6Ea>fd_,8VU)])S,UM0CM
A^Q5UDCM+S>0V(576]+/&48II?@6F9O<UaS,166:<V[Y\EA&6+YQ&@cQ:XcSNFOI
UU\+,<[W:?/3SW18[.,4+8B?3?;]<UW3K/P:a;8L6^<(5g)efR05aMARI>=_M83f
e))TI)+C\D4CbIda\DHJbOJ^-ZLLg6\AN/I_B?.CXTQ:e04F,I6;]4d0V6U]D:J^
<F;[(g.VM_;SOJFZOdX+6WY;eF9#R&N]WP22<cQU]8f?eG6;C,1=X?;EWBP)(-D3
gY]76fTe0_0EVF_L)@OOAD\<0=\GWgf:T-C5Q7=f-O;3=5]\QI<b-])06_?[R42+
8ZE;@N/WV^MR/La-E14/77IU?NW6AEQU=HF)E(-7MYTc-:VXINg(IV#@B);Z7cQ7
#=_>>UX[U.4HFH=[?dfR4A4J63#DHX:MX\-Q8\f;Zc/Z>=N^Gcg#Ga,Q?\(bZ2a/
a9WQ8fZ>O@eN3A97,C)\:>1Jda@;<CT3FfO+]e/_\0_8<=>=]R;OTc\Q5dT]HEWN
;?4C8R0,,\C8NP=5W)3#e<gaCc4()cV=LSFaggeV15#TU^SQ9.Z95eC6+_BF5DB#
U979)bQQc,/e]FXS(]WP6/aUQLg\Q@>a&<W]?IgC#-GSE[]\N.V0C)6KO?[3ZZKG
a]NKL=,/Zdeb<-C[23F_JCC4ZDYGHI00(:CT+5)45DS9;dJLR0+a]]K8EC?H&P0#
TQ[D.S=-Hf#c41CbQORe7SNA)bC7.<?Pc4@NI;BHZ\4VRJC1/I:EgDI\WU:79_3>
\YSaC6Df,__BX\H7V//_7]#]faO:f;]]JL_dJ02IP]K6<a2MADdZ^,;U[5G.XG<F
>2[VRP-1VG[@SWg5\M,fQ=8dFgD1Y.2.bBTRAg=LSE^]:FG#&DH6,5UJJ[bC-\MT
=#R(N6-.ZWc&D7geST>9G;;XHbNf.MX0>P9Af??=_\W(a&/4PXF@#U9d5BCB.[CR
\&53[2Yg_.[f.XMeV?-e>/UL5T>SNeUJG#6R.3A\d&b.d4Hg#,_D9L4YE-caTCL7
N3)=,Y=XN-/N?XRUF[CM\a&,9AO/<);IXRB5W[E#4LPbCZ]9-Qe&\[:(0Z_:CZg[
f#L;4aG5^I<VPXRGAY9P26bP0C?,NOfJAPF#0&LT:9KbH:])/UY+>1)MQ#P.[b_3
??C1c@&T7N_XZVEZU>+7@G55.WZ5W=]M4b4@bY)1V((^]\\70PbEY.W.D1)/?QIW
8fF6&>[;DZXd,(J6Y^U]f6O)?U0JTR=J^8>gTQUa7TH7^G^A+b@16SVW_\7HF/G7
)7.>EK<#<-?.,212UCWY.HN<4gVHIP[YB5dLQ.5_0BE=WAVS_(2?]N^P;61Ie_S@
.c[1MK5Z1_)/a)K7-1N,?d?+^\<SR005O.F8?AE_>D\27a>MEEM^N0J^K97W5D:<
BGDfM335SeZ^a6T7SaJ[]HfYfd31O,+YW+SOWg?N^_Dg(S/>GdH0;G3cMecB(8Bf
548O_)gdQfgLZQ;+\M_e)B4L)Y<)H7Y0PKT1<J[#WW.>Gb01AG^a#/]6SaUNR</b
8K]ScH-3=E58ZVJ@+K>3I8a8F8@-81]7JO_?XB8bGT7=8J\-/RNWJARCT<G1N-7/
O^XS5cH>c14HRIc&M1E4HYa3R/Y37,A@07de.f)G4>S+5GLIP=5=6@d04SVBd<HQ
@dOVYAb0#+;1C5&O8a6MfTT(S2(LgP@]-I:@CFLE6@RagZO^^3JR,A:KB4gP=-PE
S4A40\X-U_2UC1<fFcdN.;/CX>(c62P#)E?df5B?7bJ.52W+?8-_?#P7(YdK,N2c
VOI1X>c7X6D7=AF]2L@(]ZTPRS&YJV>=@NHKO3<0MP\?PUQSYO,:8\DJg+e4O(3[
]21BeLfE.SLc-2gAE7--(L&gcR/_5e7Q9-MY=a?&VUYf2Y1&(J)@);OY12/<:&T.
?TT,\<b@H6VQ3G>25PU(ZD_d4MD:7W+03@LB8(IFOaYEbfE23U,>A#YMQ26=1/P_
GK)55+[g7RKdQ7eT-21&(7AN#MT^H&J/#;B]\(/b,#>d,2#-J(7?9TR-\,?46]4b
RV(>e\PD45a@QG\b_2[AT__SdAL/IL[\&EG^4YUbB85DPbY6d4#F;+d:84EY;<-[
OPZ4DKJ_E\8UKf3-b;BT2=6d34Ua:fETdHg@cNL9f]-S:7aY]J-0\2I2D8DC.PEa
<?cHGVUf8ZW<&K:)8++M<e0CW&LJS3FV.=/U38g6&+SPBS^8PG+MHD]<UKc?S:DO
eRPCfFZ_/H&@#Z8^gLU]fLg\41XE8?\Ug?S8\PHSUd>Q)Z:5GBfb;fBc>BZ3WYTF
X@(S0;;PU&/WXZI_=)C9AT;[4;UGIMC/7<]bG[]OQe7<6KOO_PZ0-J[5A>Gd)++X
+IeYHf?588:0;92/?&(RFX(fg6<SE]G-1,[?E0+SX+.>@]HeeJ<A+\TY=M-dA&0]
TR7?\2]8=)d)0L3\))^HJU#a4)#B.#DN=;Y2+VA1J#U#>0c^bOD+@G#aMDS]@b[f
1TZTOQ1;5W;R(O4[cN=C(W+b(H85fCNX>Z>Eb\Y>#3[V6_HL]4_EUV[G(dVgS=gX
cTYFS5e=1DS)-S;NA>5J.8<(0;CYa_JE,H,^]N)(.\.&UFFH?7?/2^\+.I#NN,@a
^CfZ9\/Q8M4dPZ@GNEed^CLV\SX&/eH2CH0(3#1/a.NMH=>@9S-S;9^6<67DU,A1
^cBVQ5[8SDJ,aL1B,I^=NF@MA5&Z52NP:a5R8JcF=Pg+^_[,D1RQP0aT?M3-A)/#
Qd1N41@+/#1V#F.4SQ2-OWCFN/)4\EODLU][BPBZ;d4,M?[W[U6P_G#IDL576T]7
E2bgL)Q8c&ASV)&HA+(RTX,6&7K9J_9UN\fb<R[>>8\f(=9B:4Ye9geIHWGdAWH6
3M0^E:MWV&HXfNCU6W@WI5ZLg&9\V]<TJb:ZUR^4Rec[S0]2K,:7:K8C&P?]K]HA
0DV>G37FAGFF<O&UL#=gW#@Q9c<RR^+?6c5L7+@cA\XBUL-8G3X9\&ADG64#Y\e:
<GF59/8Z[8Z/bfR4b@#U@Bd5]?XGZ<7;D::5S9FB_G5CY47CbT1J-V.ZQ#B;]TJ)
+K+@Z5FS-@cW)TNf04M)#U[VFH<^B+C&f6b(?)&O4_3aE>FK/PRS3BaT:E\EJ,eM
M36U2a&P^9W3WM_0[J@/Z<Eg\4V]8R&:@4c<B]U=FW#)AW/89YHbX[C\,_&HOX>(
]+[EKCCHU@9-;H3_T<3+N(?X+&NZMR;NLa3Y_.050eMTB7/R471ce7Hdg&]YZ7(F
B=AJJC3gcQe,.:J3)-W0/S[QB-MZ75Z.=-0-e8eDUeKBR)[Z0>b0AZTdAcWGGMCG
A1aWA5HI^BR\,c<bRMd+.YHc?<4?@4Ab,+(K<Ng#8e)g:O=[NFOFT\U\F==SOKRM
M)Z:g3Ba;I]7_68TPKX/2W;?-BTU(5f]/\36cg00E&+WV59B7+00=?C=,U?NL#@Z
[S)BcLYTV@c/3>C?141@9LN^83UU,eVP+05^N<aN.d[97#]:^^#?a3CZP#d]4d@@
JQ9F_Qe+bQ+KR;CA/1\&g15b.42^ET9O_W=>B7:bK-:#ObMQGQJJA1+7[BSAf2LX
4cg#7DKVGbD3F]5AWcZ?^PX2C?a(0_a=IS5,IO4]@,5+QM;P@N2g=/\FD#_@4cP=
+aOS3I5Rf5(A+bc#H7UV:e=/X8_77?OfD?;a59-LaFecS9[649V)#4BeJ)YL1Y05
Bfbf+P53e<G\J;U9JCfGTf[#]P#5U7.I=B8#35+AYeeGSGG7I2H4.8d?<U4BO,J#
5;8T0EZ1f8W&e2J\[.=bLYCR0LZdEHD;;Pb9M>X_J]8A?GgTBUZLP;H\9ZV2(/PP
+^,XV2HNW[aTd7#K2f^0f2VKW@-+8PM#&2+Re4=>>e=M-6B#B-N-.]]#?C73FC/^
(P=:bI<+<0MT5^&a_=+78S@[&;[YBC=b(>&.<Z_cg9T@b).LZ^_>PSD,4Je^JBF_
O0Td#+4df7,,0BH8H79V5F\gcE,_?+J4=bKC9)Vd[\>C0aAbcH=a=\I&Ad(-4fD=
LbdN>(2XVNLT>[f5,2g(9TIV;K6a,?7OggdKQJ=J3;f@[H9^QI.f\_[2FEDD(+.g
Q)Y-EZ]L4ZWbceBG>ZPLWaJW6F>:?YU(_D0\8.6++,\C;HMYLY\9:+/;=&ea#2>7
C:0//&KGa5e?08/BMV(OOYO30@C2_;:U=Q<cZ>+&)@6FA86=&Z3ZJNdLE5ENA0M@
F8:[#7KA=SC18+58gK10;2#W]T,=@BR[bJ+-P5ZP4-+?,X#?aLd_LAaYR9/)?TTL
3E8;?[Ma8<@g2RCC,<6de\SG)M=OX+A3N<03F5/A9QAc#5R>J++D_-9QC/_e6&?1
gKOC0RM+V+?4Lf/O>/(M#U&(<3ZO.D?P1RTGYJ\0JEV3,.bF5aQ@1HENUM]JMJf&
[[<J0#A;_O]#]I#QL0cM/BPJ\#27eBa7AXQeI@b4+XT8JK086+FNW:bCf1BHN_&Y
[&:_-,NWdJaAI+4BUSFMQI7((.\^]VC8]?,&FZAREI8?FCX2<_@4G\c+LC9@<^[\
UJ;)H.N:H=a[=]SR-@\Y:J)22WS0G(a?<BT#:,4_PU&SQP=EL0/7B-(TQW-YI&+O
TE8Q8g8dW7EWRfO3/aXRaT__-+HTSR;I+=3N^@KQfI2RT9G],T;?+:6T3?7HgMX[
TfUVVcAOdgO.Q^0bXWK8_CA;4Vg,Y)>V=eQ.g?-^84MbZW:/O)U^F;E2]LBGcD1/
_44&0O-<WFM5aX#a]fK>=]&NKgOObcVEI@W:C/Ka4/<90G_Z^,:B@Tac@GY#POYI
7+E-W40HOG0YaR\K==4HLJ3NOIB]CQ053R7BR>[6^?-W4QfU&/<]1VgaQWQM?ZOG
5.TAI6PNQTCUOYQ0+B3)J9fg>?[,D?dHW0dc-e>:6#+C[bO>ZCZ+D-L7FFHPT=A9
F?H-:;DZEG^JM7GB@G?cgNd6T?];.dET@A\4DW>Ib=#8[gGG\Gf;T(4EDR4FV+Y=
I/)^bABCR5@Y7N/Sg2gXYWDZ5\3H_D?J4-Q\RfN<C;5GKAa]53EJ#CJLSZPJ:FgL
KGILG)7U_R.&#\@U1WY/XVEa_]@Zfa9OEC#9&@_CM.BKSUc/dcR@:gQ6;BN?#\:6
?A_C#I)_FA-A4(@K5V7&\AGc_F5]YS15c&eecLJb#_F;6#UF,^B]bHD_YOWH;:-Z
8LY7^9&>2K_.5)Kd/O#P]\A./W@HF2@6DOQ8=cH?:J\,PBTWO^SUa1/@a?9-O7MY
0=-P:T4RcJ03eR]3#9N4_46J\e\/.KSe3fVIM7Qd\W[@RU([g(Z#()41CEJ5C)]M
Xfa)K@/W)fPR97;&/F.W,]&LNH<ZX;P6;?^E1@#NRY(<--L;F#2DX8RT<Z_2[9a6
EfZA(5\2+P\E4EcF,+[L-XNW&#E@5[d/_eNM,:LL@)4-@5D87A/fWUGU,><1RgeY
Ub5gIW2+]V?V?VcBLJ5>N+B[+6g1><_4?@KV\>D8T:8J#IU3N:8&A>V7+IA57,?+
9+Jc>4BV-JUa:FTO)A:M^Z_18G9/+><CDBS79/[;46OA-Id4=@0ZLDM=.R<ZfA>G
5eb=A@U?AQI4I^SKf>?B0ZY2,BR\G=75F.Wd^_+.0.87;EL[WZKCJc[P4/W+IL@f
Uc^((.B.TH2Oe9?aBKJRCe2:=0IS?D_(:3SIKV2H-2K<]H5A#T7(g6C<93cD;DS#
g(1=d4^(6_GX=,cYR(/6aW/6N7K27D.QCB0OMb#7J5#5@(5@f_0Z;?\[Z>L&^Da<
IKBJZ/MdG:b5de^Z\b09Z&-E,=fH@=KUb=[K3E[1@:ZX)CfU=A).R7B#OISZe8(P
:_Q28Q<:MMM_#FP_d]9L=+T;K2W/97d6[,N#a6/HU),7S=T7+5W84HOM==F)KNA_
_9L@CFX/CPQ5Y_Pg,eJHD;Y>GYO(U\W1bJ0642(HJXeW_5AKCIg>I^CZfP1&:6YG
_aM8b<P,G(c<[Uf\=)DNEQD./[_-XbJY]0Zd02HEB-[XH)6;E6>D04N[0R/O^Ce3
=]9e5/NHWLe)fY9V/NC/FQ?NVNB,_IF85F97M.,6E(<G+(8fb,f-SE=?X^X,Ve@D
XZ5W;,@:]d,c84VI_XDJSeI:2Wc-<=;Fff:L(/QSW&-cIN6-WGW4FWEMNDNGd]=3
(VYJBA1Lce??Y17(0.JI[b9=gB9;VEY-:M8\e4E6DI-RcBX;269E75CBEMY?H7G[
7&4:I9Qd6EDST,2AT_?e#0cEQ-U#LX:3QPT<28@7-RN9_^9=4VH1\QY)C19HB2-I
RCbL2D_VEJUZCSaB],U;f/F_GMB9_T9?::ZW@AdgNdg&f(XN@\dL4^()N_>NNT#7
&cT38[?LP&(J1\9R_(?U:3c/gKbS(N1.f(^Y0XF>[?/BX2[?FO6AF0DFbQ>+cg_X
SM\_HgK=B4JP/+KYHf/1_VPKETQ46\F[geA/Ubg48_WG?UF9fZJQ^N9GR)d7N@CR
F/;.c->MD+].dE;ReJO<@3@-\bbR].,1>c2<0D2/.KUB598OR3EH@(UDgc+OeZg,
aaMJ\B&/A8gOKIHD+[S#0VDa#a@<JGF1gVD0Q1e/#RB?1)Z9,1X<&U+8PecPcOG(
YSeTF>E,..OZTE7E=6EB/WO_Jcf1KG[Pc=V;JAL5cbP)DKJ[.;#J6RS<07G0[E37
A^_egb;g-AA?^OU9BJU.JE(7P5)8;:GFFE,)H(HV.51b_^-[(;d3G#GDQ9XITf0V
fF-SS&GCROD[G=66,:]?0DDHRQ9N5gNdM^ZMGO3VN;M?O&0TK\J^Y+M6C68YE3F^
C0+G_IP@DFg.DSPUTTc<_Q5CBd.J=&b;_U\W2&@.IL.UK00=_cS+gPG)>;8C8Od<
>P:B8O>6^bc<MVY7A#CD;K(&5>YS?A.E68PG:IH.a\@,8:Cg&gOSO9P&7LBZI3=>
7Z+)M)Y3&5]UNHdMX3EOJDG6))T@=aCR84\PM/RcJ>J6;C[O&=Bc/f(<fa+6)fN)
;NRf(3N>b3BR-8aQOa/CA^[\.@EMEGBdcUbS=CL<H+_QV<g;cEU7eK?:4]:O.BF7
9M__8/JB3/E2^;NGTdL)NVccL@6A\N9=g1W1Uf,g?eN5&(63#M=4B;]1(>eWS(c]
C@HSM^3a6S<:YE]JXeTE#Y75W@Y5<,B5;SR2ZZOeKgW#PJUe>Y5M6g6ZQUdZVf[g
5TINZ6]CVEcJW9WDVL@J(7,[4G+NZ,YWbe0c_I6eE5OI5=ZPScYW-;EfG+D5IJY4
NAVTO1)C9\)E50#WZ<e6)\NQ,GN1bW6_]DXM=bLBe@7MCOMdN5&QU__+T-3e-9AS
UVcbeDQNJ[AgS##c9eB@QId6\T?<c&/^&_bWdf+5CX<H+M3[&FE,DOd//QRM&bRP
DI]E(3[(\/0E]eS[^Q8_d\AJ7(Q.7][L+Y0M8\99H9;Z>^AU1a8;+EYW3]gNT.A+
>/@a82<&@cE2e\<II>I@WFg>],GV)+4C0_P?P66B07WFK1<&?151)+=S^;2L7-5J
Q-KLcRY53FcR>5I]=M)RfafQ<\27WW,1XPM>7VWR[&7<eMK/3X<>eOI@W;X6+>VD
;?>E)WVZB(-:McIG#DXgU+M?9FbfW=8U8O&&&VR[S7A#9^3JYbe([+E+J[M@J;.S
d=a-T9]-^UWG41+;-M_]#:g;HMa2-&FP;\LRdQ(;W3&gd7P.B)(P&H4&,.\QbK=.
gPO(d8P.,fS#e1W:&CeRd1C1WdVMSD75D9?[05#M1B.^d<-4K@+YD\FcCbBdL-4)
.\<RBL>6NJeIW@8<Z^(;X>a4d\W^3BW>0fe(J_.#070124aa,f>SYYH?90]MgWPG
53da^FZ@&G6+JH7:RKR&KZ)]]CO#M?A&=@[:;8,1ZSdP?+,,Oc:\B_bd/QICI?f)
C:;4LFHc+7J]^;b3B<\)3SEU4H<89;f/@Fg_d0d-C<[6QKLLeRaZ#GYWJcbMY[W1
>;E2fbdYb/Te#X/4WfU/9-?8::FT1CNaYVb6Va@Ha0;WB,+AO6[N8B;?e8.d:5(8
XN0KWNH.J7,a6A,7H51C(H5&LSY917-C0;.Z+P+O.\4&,3C,WagBQ8WB4>BaZd+U
BJO-(^UD(3_cB;fZ<QU21ADK4+663?-VF;5d+7Wg<0&bb2f5YN8ET?f;)4W44485
c@DM(0OeBR&@H0-_1<LUZI;_@OOb(e).GaK,g&2B(6c#Vc>ZdPDG0PTLTTWE@>KQ
29_dN,Z(/ZJL)5<?_aXK9fGDB75d\R^dD^DI4=KQ\gPQC-3=@HL;)^LJS0cC0^He
@@Tc<@S,TEfVIC:&a:8g;3.b/X.:EAa>3\7.-0(62,[7dI0LQIS@6K)ged^T-H,-
AJ+38,WQfW<@RWcRg7O8c4+SD[M6]HPN,CX3/>3@A<2PVA]_)+?E/1Q[\5DEg;Q&
)E]^cP[PU7_\BA=;V\I36?J-GA8:4X)a?e<fW8T_cSaCgO<.8GMK/&NI+S#8K>J)
Z5G:F39.LX9E0DQ?2fO84[,9)>F^3\/DDH@0EE>Y56QKd8L)YR5F2:,[Y4.1=NR7
C68:S(X?2g^]22>:c&A1U#W/1KKc9@TbERDXX2AW?;[Y/OGPZL1(C/_W^SUD?Cb]
\S(HO#cD^OD]-[E)-7=P+2-RMY>?O5-N>5>P7,GZ/ORLP2Y-bFf?))a<\OP0gda,
N30[D4)>3N.:cPIB)HfNc>]UF6aaIRB?EYQ4P2W]O#U_3S(]AM.^&OfCM2YST<W)
=D5R3+VRM?C^\)TG4WX+G]OV&>^F\<(EM39&I2\O6[YB&MS(H3fH.-Q0_WFUf^>X
E#Z=BVIW@V5,fAb96OKSf7VIK24<X3DVac,^L&RD\ZN?E=)AOd72dU=GX8b1dJ-d
4)7>@3f>&9cfeae=<EMeGY)IM-G4CWT6#T;Z)@)E4FG\;^L&K\a]1\)TN<:I4W\]
cI&FHY66eCXBRQXU[W+Q:L9A/(U,SN5#.@1:JTfA3?:^2QdO@@g50O(2T@0702e\
K)RZeaVU3BFgeK^&B5NUDeE]_;RI-D_Z0a\HSF,V&YR7K3S?:)M=_Ye;W..R:=MC
Y@;60L]T58gH@I+R8R0#dZ:E@Ra;.\F,JUacVeD@T@1D4QWLW_@-9DE85L_T3Q[Y
&5VFS,#gC849Q4dXfR;J&4,U[LA+&Ac@T_Z<?SZ<#4=Wfe2SH?;5C(NL:7V6<]0E
d<+]AS-J[S)Z8f1fT>#H2J6c-I,Nb._KTR#6@,3A1+PDT+0S[\YX:+b-aN[\W.V.
XX3+D+ANHUc@7J8AB3aJ#.U^eV\F/HD<BH5]9H;[\fARA6261?Y11SR\O,;)=CY9
Ad5f&R.?+V3KcT.])?cD.2BBGLJ#<NWf6+R#C5\@B+,&0)+=gaT).T?ISE+(D=5&
c0P40HLM^60d8NRcSIb9Y^-Z\KWJd/Q,=aL;P[Q6;#3_d5S&2FM^V5ON:S<X9&[O
ed\E03/IRg_<M88@1(ceeM5F)B>[5Ce5-JETS)MY,N0f,OXZ-JA^fP?A476#FU]=
_g]OU]@D[T?^)F/F.PgaWHH+eICTEeUR9TUY1/>-\Q_IBX(c;aCXOORDdc1bJY.d
MW/LTLU8eFF6GH(F],@<eQV8/YN#..Bb:0EfVaPaa4_5>QRF:X\C):X8U2[=_b@9
Tf5VG)Kd:<-L8g.E^K=F0\R75L8D?gIdOU:SRV?=9_RAPG,,M<&]J^L4UN5@Y>>8
]fLe2&2+1VP@#/(SH&Z94Pb.cRcBC?GA#].RFZ83W04@/<BA+L.g5Ra8RF9RU8e:
65M=.A8[L3;LJ;,@\)/IL8P]@,XJ[>d2R0=B7Z^E^dN;_G.g?ZaC3\@M==T&g)/_
N?GO7KK8AN[=?@^Q\J)G6-EGCSJD?Mc+C_@?f(aDR&Kf6;I;C,@,&=,34MOAB^gU
O9@IVZMe3@<D:@2L3/5:EgO?Fb(3@S=UX6d#JL?Rd/-SO?+^/B<DBN3-C>c;4_O;
Q(.HLHD&);LU/:R5-gLL^@2a^#4MJ(WTC-)3_)LTb/EBF6TVfXRC#+aCNDZDBOA=
VZFD.=aLRS@;CHVX6Bg]b.A_dKYQ_5_F,I02aRR+eGSf]8e3A+])aKR[T3]4B?98
edKc_JP_ZJ)KO0?,OX6#/fUJ6YL5\7dV)5V^Db7W-R^aC]MH]@83E5N@FTAeDG,c
RD2L,8:Ncbg2g/OH:M?87+Z772efTN&4P37I?WUK_d6#T9.&BT39TXX@DRAH?GHM
bUP;&D?+e8).GKf??4[;@455]K9E#:J\RgQ21b2X(?UF\DL=^,GCHQC=H/Q>Z]^2
2DPaQ_Y)R5(I84QcFL#/+ZH-L]<&#?9B,d<#(P7MRd.(eGFW\XRJ&RL0.H2_9)f;
)e+e30J]6&IK#dR-0JB^&;A1QM3TV85IWd=N)PEOF1aS6;68@?)d?-4d8+<OLgZ3
+(?)MK[G:#BU=:R3AW^f[SZS,3^KC23W(5\-Q(OMWSY8_M<OR?\AXNDdecaT_(8e
C/HKCHUQ\7/J_QHP3=PAWT:2\D9\c;ZRd?F^S[Pef^FdS;ETe4X)W)NY[D??PGT]
3A-(J;QQW+MBg#[(L+H5AU-\B:Y94=1G(..1:X_HddI[.QHDP;XT_gaRBISQEBWF
L0^/#WNUKB+,PQ@0.6gfYM@5JVQbf=XLH(CHgWXS@IeFba<g5^XFaE/]U6&^WAAG
?DLTC5WcBaF.B0a-;b<6D@&V],8_S?\TJ/GBK(I#<79/@[BcAVJ;)A85FR>aJ<?d
9^7Gab+@9.8gHE)(N9&U5\00/YWB?g+F>BD?5PIcA(KDgJ3dY.VcI-e3dR19-96G
7T1)D+VHW=MDVL>1=8GX&3TH?5Y.ZYeY#f\B=CIa4&AO>T_B2ag=MJe38^N1O]0-
W0#<1.<cDXGWa:I-e[;cbgX+J=L2F7(YQK9=]5P,Yg+9-1O+2<)aU[9&aRV_P>N=
RV,UF[&&-.12O88.WWR<7)+RI?;#?72G2L2WCG03DS?QRZ7\YGVSa\cOP#&IWUTB
2W?S:^9M(2S4H:3A#(G&M:GC5>7HI)1a^^QL@E[RcCF2@#K\CSg<J[C.+F=T^(0T
U,6ZHSdFgME009(ED@,QSH\_J]45:O_bS<A4VF.PD@X(@HH8YcKEf,X8VOAQa+=R
^-.9:8I5(P.ZLXbEagJ9XH#C7A8NIaO(D,D/_(T4UX;B=HRAV+L0I6=[GXD>Ic_M
e5T@C>(K8F1WPQDBVV#^@EbbePK,O58-.G<+AP:@T^7#^K3^#cM:-b>_2d9B/H(+
V\f65^O_&b(R]VH[320fA7C<F7(?2[JbB1LR)ZV++;a):#5a][J6OZW+:;75@0SB
FJEL6-;K[^R.g0&AeO0c6?-D)<[IX+_dB<\5@c/[DM+gE8I_ZKSF^?:TF,<cN^QQ
LEaPHGC6ef9I0_T-<,)#P+#<_J#8fR/S:QaXJ5dHTC022@;L=8J=5GQH0&,F[0H2
OLE06MMcTUQKC9MZYAM,c2)<<V]9T8Z@.@#=I/]IK:FbE?1#^&UD3FO1M@796f2@
RSYE@-0+A;6E?ZV9\_DOWN:?]Kf?L?;:?6.7FM/O/8]dPC0aR9.cS^D,-L)cYIHD
7/;SK5X49c(UD6+@4U59/[He35BSE\:<(_5H^<1b&;<L#?M3RS\Ldg&&WXBPeFH\
\.,98GWAaHF8VKOQA0A[K7.81SJ<]I>.CUXQF]1X2>d309&=]BTD7f9;:\19,L)U
?>L7-08#D-]FDfZ0&6FNF/[fAGB[,+WM)SQRFEWYgdL1Ka);#0S#VJ#D5d/B,]PE
6B3(J/R1Pbb2E]_R5UKM7\O:]H3;)2Q\E7D31[(_5AKRA_D(52@UW01POBOIL&6[
L2I&(g==7O)e1^-:I01>K+/7W43f=@d<a_R&JI_UYRF(1-&8-XMUg^bYU@(P]fRR
J46N\AS8OT5GU0TVCg&;bYH7a4K55=Cb+-#P/@5ag<RcT=dCHIcO6VI&HceZ9H[c
0B48XYSP]]<J?UG+L83E8-TR+J6GD8[:__D@_O]aJ,cIY7GR:b>S^Y\2@V]<N&f9
L-Leb+\TKWO?-8#=Sd5;-E14UQG2)NHRS<U/6V4>9O[gdf(;0^7P,bDa2WMbWME_
[K@II^Ybe+[J\/3-Z]4W99c&2XQK0:]H?0C3g>:/P4-#g3-[V_TRISKAQ7HX1B,F
[>388U3,(\,D,c77[:92.4/?@35[&UJJ08cH__B&c6Kg-)V2-;+=/OR#+K9<Kb9^
,aCLO1RSK_+S6?ZKb6Z6SFXHc0+8<bd_<KEP4]&EfOeLaF/=,NI)Y]-.EJ/(XQ3N
<)5K4aOV^Y65T?]W=P04fKe=a@7<0DTUNCK]Y\RYY?).ZBJV9gE/5BO&a2_N&YGO
CU))-\?g-M:7T_O[ZTY;TE(edDdFY.dcLMa&f3#V^1G3gV>=619TKW,-4Y=5:I3U
H=@3WZ-VA6]RNOEB2NPDQZ64LK.QQAEIQb0YCTYbe:FO/5^1IT4XG@D5V;RI>Q,c
YHGEW;))f9?+-d/7[F7-<0SF]>O8;6IZLLT?Z]E<acf>,b;RBXKW:GMa.5>&9S^<
f6LRL@-AS#OS[\+eb=JT7??E5>+<-?H9F>d4@ePeE9U_Y][&@_:X6>OWg-_V#B[Z
7Ae1R&cSf>+F)V1(6)e<1dBQN.^5SXGaC^#T>HV6S+]d--Ye(J+JSAXd#2BCSF=I
FdT86P5L340IZ7f=5PHBLP9U-9a\#EL5/P5+A^4)<NB2H^8D-1_H:W(b0V-U#_J)
A3N^D4YeWCAgWPJV3d]]Q3C9P5LVY-dTZ9C1>V\21;M5Y=SU5,R[N7DeLB/Ga)D?
EO^+f.+\J-+4DPVMD]2SdY-_<Q?P,0:_((^9g_2#(O)J#@^5IPN@H/<]MM33VKgd
)f2=AMc]6dNL,N^H&/\a5,fO7AGDDcff,F4=gcCL2T+KEaT/^2;cf-(f;S@;\?F1
VT4XWeJF<<aXSJ;6+A&e921XEB5UKQXP86Z/5H/ce&01NN]gW#[:FggZ\Q&8PL<7
,Af5WM:G2@6F5<ba&[/\bI.beCK3a5(&M7,AfR/2(1=F6=g-M8..OIDXT:e\gIaT
V;,8f.>FNP=XW=P5f;S:41P#g_U1F\RZXT7;[;#H.-O_fd30YfK5c1bJ<XYK<c7;
3GaN_P^4WA/ZP.U<7/>ScR(M6TbBI44OKfMZ,6@<<8,HF/bV4^ORG9)6+YXI9],f
YQV)L(43B.:Y4+(M<d/PKc#^5<\7dgA)HO2@OHYEcQ/7ZLRE(FZ&I.<.cGD;gP37
7=6>@d<?<&IN/F;Y_f_:4OE:+VI=]JU^Je5MdMR:Y:9C3\<6&1:YKTLM4Jb#]:?d
Xd^:F8QNc6K4AT]3<#f.9N#g<,b]b>+-g#GfH9RBY5^T0,HGPS#/=WV,gPV\,J,J
]4URD4PP]M4Rd\5UbJ)=_JPFe1SB6&3+\6,[gS&XDNUfDeRZBb:7HB1@,:UbX]11
I#/_VX_;)\)T?9\-IX;DX&5)3H8+[5dVfUS&=b9Ge=(;K_?7dfF@@]^8cYe+Xf(#
RG>\(7[5&K&D\2,_8G<YSP<TQ[MUVdK>\634M(a1S2[WL==gJVH2+SQV&=TJgIa^
)[WK_^e:.Z30W6P3Q-gU88]#L07bDE:b30[B5N,CNDMfXXM?E=W&5(41L&?XZQM@
LN9AFaI[0S=JN0DRZe];S<#M5C2)?@E_-JD&)?1e.E6#K7P(Y)Q73#,BU<PFH-XD
]7FGURa<H1UJP[?L2f2<Qd-c^.6D:BX-0E4gL?DP&#b5B,ANK<-1_YT)PR6A0/XC
8IT[89f5F;\Y:-/HB7d9VH_/K1&B/N6M(&30=]E4B^076<.,09a2;EX#HIdDBT#A
XR6NT&K\)T=L4=bAC&6eGXH(=BaU:^LO7E@]S/FMg\50#DA?+4.F75fcV+P7:T+O
;^)?9M7OW68EUea#;8C5O+/88b>aZ;-F5cYL9+f>0G&B>(&^CY-K9C:a9I3ZF2U^
e-,[SB#d;a1=2d5ZF1T16:H<-9@L0E[+#8E+,C@&Le:/E1WN6YI/a4DS-X,]APZ,
S@KL-6W>I_\LRTP]WK22TL4<b_D50K9PE:5QB#-PD,4EN(H9IU+C0d2=a=LEVB66
L6G8<PST>bJG?()=>QAU4ObD=TNf9Sa5CZ_4G?c>DV(g/IPO1.L4^6ZLKA)cU.I;
GVgKWgTC.H4=42XM9&XXPfU(C;3#IgC1V?9.-9+PA+EO=K&1J@_62/V6G_645,-+
_P5U?1>I9[a7>=VE4:Kg]UI+f,eV\;WV/L<R<NU=J@/D;3\:=K_V-a.Gc0Ng/Ma@
,;8;4N0#^1\[B/I4c1eC.a+B](_CLI7W2\Sec#-AMIKa7O?,VcPf_[E<5g8MFE&F
4M>W.7D,Y_HW]aPG\)\g3A562K1>C-7,AG=K@^/f42XD5G]),67QPecXDO@?UJL(
L^_813EgZO3(.LBG?c=XT^AWe1V>+IgC\34O:)\AHYC4Sg8N)>-e2@R<M]e6RbB0
ScL[K@VRH6[1ca,CESgf7UW>&7YU820)KHd)50:<DbD/<]9&\]Y;8&g[dRI,K>K,
@+LSe;.L)::WdfPa5W[Fc4_S>UU.X:<d6=9=7^ZYL(O3c44ebOGN::b]FH^0=23S
60O.M#c,+?c>[Obe8GITFA&>L4_:g1=\\02RDfE19GU6;.FSZJ21e77b0,W^PdVA
a/_,gI]MB]1Pf[FF[\PG7=[SN.C>WS>W<[][3[9ABCg?g45=K5P_P<YDP@?-OI]]
4;_XMSY&/-\ceZV].d2gQga1(]ab3^(5@d0geMCJPe9S;S>+.cX&7QH:-HOa#LI6
RKPCICe6YV@gC&U2J?/ADZ_5K3e.Xc8;dMab+8X5=Yb;<H?TI+Pf,S>DU@^(HWeG
(7YV+2MM11&(@G(g;Q(Z/HDQOdPK.;-WG/cLG5Q+Jaa=U=HcR8K<e9@[Y5X2VcOV
QB]^@+.>EIe76fPVa;e=[&9YCZVa?2];b=3E)K,+)_NO,S5Q>U-YX2Hbc19S<;g,
QZKGN]Kg=>N:#8ZRF8a6B70O[O5J\U9D16)7IK(GB;QF8MBE6M(OWWZU/^0=+?]d
fBS1b+&_fB-aaFHPd.5@93c-8Uc>PIG:e,96W^FE@e6/K[OR#?S/M)NRQ8,-HKD,
9H9?BDSeW;>aKV\8g>5[GRISS/Be\YWYV7XN)_fZ^\T#f.SeM7,a4H-(G(),LO21
fAVbK#QM@7]2WY6H-<9T1\+\Z:P3b<[G.YBabb91V&M^N-Ob4?I[^#=-CS[gd4Hb
U3Q4[8X+\>IM\\)(Tg#9\\bK_G(/cZ^_+T/RUd8\dEa=d<T1:AR,fG_EEV_7YK.H
1;>+M6JRG(c(W@E0QG:ZE]S<^^]E6-NXEPIX&2f4.11@I7=FK?4<064[U<CbDLO\
5bVSD>BQd;SeWZYL\1ETV(-c.#OX-V^]Qf^7)6bCG:5eK+IbXQ\C57Ra2@_eUaQ7
]#8F_BLAVJaBD-Dc=-,]ZWcM2R__Tb24AWf.0XEZ,#-VCK-)ZE,ECU6#WUA[fY(_
a^=[2P18BK(_.N5LTBV9)^gb;\Paf^d_:QQ,W2<Z&QU_08]HT7b=K3EQg1?ZYT\-
>gJ\VF==V;B2\TWWI,;EJZNH/?E;BSAI37?VdfGT2V2a8JSGNOUaXBF_?[R=:U>M
R?->cDCSc]-PW)R1gD.7NaO@?7ATeI(G_AI3];f:6TFV\<4A.G&@=X.</b8(E+T0
FTBVON@bA&CX:.<Y?\Oe+(_IaMPYO.L<,)]K-S?5QL1,&;:8cWBMOG(:YRE1T6SJ
AW&f)^-MSN=-31J,+X^==&DE;-Kaf,eScQ06]IUg/DE9ed<&QQ4MZ<ZAZF5@&9-\
>PNc36R^f,e+cNNT9P/XRE@8+1[6dF>Ig([PB/?@9W(TQTcUc<FS<53W<A9_#8#W
5)V.4#FJ_[gX;1QG5Z@H(Tca@YF1_@@WWg+?Z[e7H_?0E0M4FJ#@YFC>M<Zd6#QI
QUb,-^<G1?_-5=GUag1XUJQTD<#T(D15Y@UA4JNQ-<TPN;4O3QQ(Q#&?fP)^MUZb
.<()a^0Y<C=-GVJV</F^[3=U44AFg7Pa:RTG8F+aADYVd,F7ZHGE-:L(606FS?C/
TQB7c.+U=M/]6>61WBcA&:8Nc/<2<^KY9<IU3ZT)\;DPNL?A,XK\D.AH8:#3),aM
+0FLg85Q>;KWO^ZYO-bVSK:=TNX:ZY:#BN?S?2Z;PbUG4Z)L-;3)D0NbFc6Ca(^N
G:F/?E<;4Y]1V@cG:A/[LOV5gFR2ET34)W^a;<21YQ-<UOLV)QcN;g_Xa/]Z&<eK
>&2T3UUU-Z=WJB?fcN8/Q^Q?[U8?B=1&FV_OX(+\6eLGbXKKb@&C.3M0<66+\YU\
MJ7Y[5P(TbfX/5VgC)(.b=UHg]AU/S.M30d#W)D(f&LZ2JWB?73H0EZKV&0F;<cJ
c:>YMSV9bCc&_QB?cbL=1GU@H:dW9g4NO_,&4PP-/>e#.b=G/WJZZ)aF_a(HgRRb
<HEN=,C/V1YE6(&)I<9Y7[T\HP40-BHNQ+.AYQW=Y9c/ZbYPTaX3QGZXTC_:X:.+
?7;c5(a;;]DAZXAF#\Kb1[5P9<f@L^\8-.X6@Nc=R?EJ9O:T68?EaEa1,ZF6XGIR
PUK+^^QK7WF2GZP[H5U6X&<WQ]If(&c1[JgGM^7V,T4#(ZLF>A4U\];(V<gNgF&L
fg?^<JZRU\IbdCe9@=F+dea>adTC4VX77?JgTM[[ATQVN7R7^)BRCYRUHJ.OW=aQ
bGMBDZUHea,9V7.Uad;2AU[]ZAD#<AV^I--&^L04/TO#-DBB6=2-?>@MgUC/:EEI
fN&4IUT0:QW2g&I88eE=a..1.KZ_>E[Q,C?/4L/1d2P(a[\0N?>?:PJSNGg.\>&\
1&NF;CK5Y7;eC/A(JCe_IZ31CQ<&J++aI()BL1IE12/f=@V+==e7O+E8/KW38Z<F
V\fGO[?PO2[CdZg>K__/FX)^N_bF2I8]&@^Mag@&;I+f=a#2d?><]?MQ>5_=2AFZ
Y,TUM<D3&JfR8;IGD@3JfaSB#gbCTe7_f[/V5X>ef:1>;M8F8KY.+.g?)1AF[-M3
@FD,O;UY+.]:=#L=Q/KcH<,4<RHQNN:V]Vf9K&UKI6JAe2P(B_6YAMcTDO>E(Dg#
Fc+CIFWW40;&D^WEB_&?J?QM8bYI-?:TO@H=8aaDP#g@4gA:B.-3ML7HN:<K@g3[
e89,JGM@bYSZ_CPbf(KT/V;d=C(#DU3R]__N-\;D;PcXNbF+f8If)EO,cJ&HJa(I
J-IX^FRN&(b/e.61R9b=AFRaV[A4+IBIFc6R2MeJI(@^]QIQZ\^Q-H9BfG9LVZUF
1I_Q;JVX^>WT,9cC3C5PWcIXXVEb/)5gI-SAJJWS]Q\Fe0:LJ>_dFMG?VABQ,/6O
fb+8F]\040&09Y>Z?AgI(B^(/.+^56EMI_geAF0-X:SNf:=<N&+?6AGOHEb\UXF&
W&53gd2\;GbUCc^5cHgZd3&.E+ZU;b<B7C(\]UNcLXH6ROVRR.;TaF>VGe_8ScL6
UMB[0VH&I/:)NY188(PQEJFX)HR4gA)-I3KU]]BIZBE+Z28BDf-d7]4F,QH?+gSU
V\=TKOMW=5XZT?b:60AV>UBb;DX&Q5AJ\2(gTLVg?d]G.D4](1-\JaZdENXO=c^2
^g38<9VUL,L]Y4])3:B^:a/;_=P(gP:\)>_Z849[bX2N)EDTOKc[K@2aQUCK(bC.
LKUMSXS=:2>(T_5^Z3aA=eECBVG/f7a<+4d4[]HSC^KOD\_JC(2.XLK[-W]8/,GG
P;<@ZW2cPX)8dUO1\Y9&THW3f/]09[Z6J\QB23>=c+#fAa6].B?B7@LM/1];K[3c
L3eHKH?RCHd[f&[Z#I&QTGFJ3(f2bPF<_Xa(R=]dYMgNeM#-8GbJ\,&ER^ZI&F.]
V)IF=P&c0@OZ1S6C.K&a]a3.;a;.<bJ;9U,KN=_0^DM68fE5KV(+J^??=B<F,72V
E9CD\QGR(4fZTYU:X1U8AS:0ESCL)T[c1Q_>_g>6)L4EF,@)CI>PQBS^\b?MBF<A
X1&ST;<>Y(R6YC+.V[]c:H4Da35&.BDe(f_7g<).+fc4()SCJFc.K[Ofb2G5>bg^
)AA53AF?E[/3-bJK=:BWO=7,2?2d@+7[-gD(]_]3.)V3Y?6SB<G1(BL]d\)7:_&&
RCfTSa6=O0B;2@4&Y)?F7Dga_dAe7Zg6N<dK&U2NaN)9GA^D(AF8S[##F91X@([f
)]47IBZQ+FdZ8#<g5QAO\[#]D>17^0;c<M2I=^,2gI:A.(]]U0+f@6H&;Tbb6/+-
/P;J:P6HY;0Q<ge)F[05GM[IRKU8O@>2VBYeM9BF,HQ<7bY>c4=Ia(M2KQ)UT@LF
#NeJCD7_-,eSYI.2N9B7)AHMWFDe37NPAIZU;@PIP1PS.<CR4ZYa3SbBRI+L<H@_
0b>7GRVB5]dFJH9ONbV+NQ;QUAZDUPZ\8PAIe15_R@/IZ)G)b>ZDb5[TcIF2SX7d
T[-GVJ^@;f6g6=]e4D6F9H7W_K5[..-6J-P0(>f-R/Ha?S-,?TAR,EcLZ]9_Td47
33TT9.\88;FR]BF>+e]\AUAb[[N^WIT^)F,K#6P]8<G(1e^(KNI2\H0]4a#G3baM
>WM1M;)G,QbgM)FKAO^S^&9?RK#ZBHV1+X.TR[NXUTGH\e<>15T9;0J0XSOdC8a0
eggR4C-FC^@?]Y&,GAYOD__)/=GCYa]\cME>,gd[bXVTTJ);B6DU^Pb(]D/230U5
RX7>1ZO#T/6L8\^EP]\.5\3C#bd2:?/E\+.J\]b4G_NB;A@Hd5]W/CeXb67CB9,0
JQ^Lf[dU:FO4/.PgI/XIfM[?R\VJ&Ud6ITBJ-1S9KXF0ADJW9UB(8:cQ;Acc&Ye&
B&B,WVC,G+S[VGZH.SQX:a/EJ&a@->B#<T763+G,0A3CZDS&]+(,O::+6GSWEeeU
\6A/QD/.>88(.Ib/@+7;87EV8QT2[SDE+?\S.>_\SP<U7#JT[T)g93U-V)f/,?]^
d\L@G^Y98A@#Y7;Xaf/V3]L=aF)3fKV<+@,K7)?2Eb7#?BSH#c#ES]P]4UIMB@g[
T4_UC?7K>N3E[#T^MI>2++UT>KVXXd5(6P^7I[&ON<^fE#Y;S;T1GB8ZD,Oc96/?
]\Rb;FdQ@9TK=VTe@Fee/.&_;FB4;:9C/ME.JF1O9PT(XZb(K=+180F\Q;TI[>Bd
0H:E0FW9C?KA1J67QV>RD\cRZge5PT=K4,ZK?\T/&U6>4K@.-(E2XT3_F&)1CCT&
?QBK.:&_F(7[#ACPCV5D@eQ#\1f_D0BNfb8OEZ/f)#M@#S,eB]09\:--)Zf)Zb&G
<RMg4KIKGR\=.fCb8b^.CEI1W6.[+1+5>NcNZTW&cD-:+#Fc&dB]PaR1f9OKHJ6T
&?,ZX1R\A,ZJ21R&bIM5b2L,8=Nad3X;7C15J>WGL>K7](>^1JM#7A]_fR:6Y0/_
DQ)-f4_2J3CJ6T/K<,J&[b]9^B_S4_Afgdf?Jb@_9&FH31[VI5\\G&^5LQ9HEGf1
<effCO33>>eWc7YCVAEbe=[7K^1U;bUf]S-:#COd&CNbNMF\7#/PeZ&5PbLAF=bT
F=e(CA0.)IMMV>(U)@\DdX.[a2/YL4W2L#eZG]5R6B.W]<@Q73S;ET&gM]AKB6+:
=T@CFf<9I9;.(_&)/:K:3;A5f_:9M&\M#/-T;/NdKGZYUN^KJ2Zd#KEC5P_HI60;
5(\4bH1:#U1).=2e2V5^edM)/\X#6/A-=G7A6&L^,[<\[+E#?MNQg7MVC6_QWf[U
2?A65.K9;?&Bcf,TD/CEH<X/>1g.7>],N(V<<,b9C=61b,=/T6=59AfYZ5ReLKA;
=OZJS2ae=Bae<RfQ&40_4TS/Y5&\>JeGfdOK?f/d39Md-f320<KVBf[K9D5U#Y8B
aU;)V#=b;gE7/QHS@_V9,B6d03.?L-g1c<RGU+/J(FR&]IK5M&EN+6dLQZYD=C5@
W-30/JO-e=U7F)RP59d0?ZM]3Y^C8[WH[M(1\A[]22fU=Hd0=YL:@aDDba);JeK?
UHUH17&I]<][a&S4Q@f)\MZ:;/<a)0RC0&GW[P8/)&W=b#/Y_DE,WAO[NU/5H9d&
/7f\a6\,+\(&H0MMg#f_MY-JBT;/TPW&M?N)LSC&Paf3MF#@gH?7[HT=6RM_4e@@
5Z.eRQ1_;WLOXT=[?6R(^FWVd3N#e1Tc(W#R/P0LBgO#eecP1G2YK+-(HVJ1A(&7
SQ8Z[Z)BeQM4a[5gG=1R+c;>fgG\HO=BBG&7fa#.Z[<#>9844-M]JTU(UW.L++=T
05RcO5T+(BJ+Ga.Q(]=VA0+DObfPR=CAc).I<=3d[d^3<8T+c++)4;1O4MN.O^@=
aAFU1Ne<:3WC1W#(5c3.T5K2YEf:G[I#8Tgd+WgII/PP);A?[f8,QAOS1A[HW8H(
@^=]_#7#XK5E,a1eZ0<83WV&OHL,4MI.P=MAQ##MU>TTHG(cQ6XYCIJDT2cD>KC)
]#I@2\D]2VHSd?4QTM.(<K],eR[>CGb,1d;U&JL??LN,SF5T6TL;K(fA8C[)O\<<
FH4EQ_6bHJ^@.^<HCNf>Rd^@g:[-]_[G=HD=FeTOaC:C+P?^0\JXD_BA:cfEcE)>
SOPN+,QV-I[(J:I#HD?DQ^@?)9<fX=1(A?51D/+?]5KGE,-]T4:@C)^#SEeCUB?a
e3]T&a@YZA&3\R:#AB>=:eSG_QaR4,/Eef\EdHGgS_JZ>MB>M.D_bT]C#eadCQeZ
d7DUZU(YXP045-2Ac=:VQ)F<974[OY0O@fa?V[^(Z=?/(J5<Be?f=I1]QO_S-&<D
EN<YPHdVQ;\=:M:>KP[AJAB7C[29A2L9=Ye6c-4d?.>L>@;)R[2SdL)N=O(;)S8D
M[45/QF?Y:EA307_HI_X[P8?[SW7.PZUQREK<88RKQ/N93[P+?FI7:DSTHG\[Wg>
J(d.G,\P#1#)<41J2WE(7-U#ZEgZ;MdQI=N3=V__C9B5\94DB63-\Z6XN;_5WGFM
UV:KO;ZfKJ/G4:]Cff6>cR4E6)9I#-74UUQ7WEVU6BB/)LE+d\R6;c?7VEJ996G+
F3W(K:GT(LSMO9aAfK+MBB63O]EF/2[_5^3>S\<^d^CII0(7@)[g2<(f>2BG89-W
BBb)W<)(T(<Yc=Z@e]7B7Qe<<ZVE;Ja@/3;OcaH0_.@6SDK7?N4.:5/YRfKK0Q=_
64Uf,[6HAg)3QCTaU2IJ_c@N7A.9fD<:F20gGKAG[#9QPWge@=;R1I:Jc58e7?1H
>\1L#Vc5O?_Ce\,^caD-B.g7FIA8@:cV@JT?eZ9@+#&34d7Sf>J(<&XYPc8[.N.J
SGf;F^&dDS>W2Y/K2D&:gQ2(c+La=QK?f##CY&DV]][W)?@5b.A7+0ZZb_:BQSJB
.S67gX@X3;O&Y:6P=S1=H,LU@,R/cK.4V3Kg,FRe2_>VE_T;^^If+08)<cB[dOTN
XCQE]VGa^@XJX[61KFN_c9CE7>UK)#\<NY.2YA:9=_88d6a9J>GB+61.^8G>BX8P
7@W<VZAXVL4W8/=[DW2:QCg#B#H-6Z\T2=,?;K#9PdB/JI_A7-cV+118=_,/VfQX
)8#3VPVFJ35)[9##A_&?9c:0c7ZB.AD[#Y0I-V9BHWb4PFVA-NY&8g[?LN8PIZg^
gGR))._T3<dVcXQ=>2BQ6HF[Id3cg1AE3=MQ3;7;TU8Eb,#CSHKW+/G,@I7\b:Md
Y(A9@1):dc_a#a+)2O2^3e#A#J4L772E4Gf)P9F:AR?X@KA+<WI+V7_&9b>1UY<U
Z:[>HfL[Le10gd46)d?3&C=J-DL_KL:9GbfH#@CKZf6?8XX<NKBM(Q1gM5NSDN1?
NRJQ^I1cE7[U/Q=.dWGB7[[4]>C:(P04G?9R^eBA[9KW4Va05S9]3BD<cBULEDU&
D63T>W;);R-GD,aT^_5^/0T.fC([93:DVBea0(WU+<[79]M@0HRJd1.3d+X&gJ:A
3SODg2cII\_5<-#5><fZR-YPV)dYJ0G0ZTd&GS5^Q0W]L=TG5+PQLH]?G[ANZg6L
CR#1U8TN:bg9J^A3L^9<@93^R:OT,_H/5&3E?[+RC#KS:5_a9J56G6SBbgJOf+SW
D>\WTT]:_9XB4BJ>=IKD^4e.5Mg)<.P4[@JJ=YI).ed)aO=5C=\)(:I<AYCdPc?N
#02K+&EU<NG@@3]96]@QG6N4<&+\0=3A<#9g9VX]2,UBQG#(0]<&OeJ@)BBe<GT>
=8/e7#(H)<^LB=Cd1+BOZ&5YNO1?:0MU&I0-Yb0-FU^?aETa<K6HDRZ^G:X9LQfR
ZS0_-3dMOKcde<--YU7RT^UKPB;B(I5C@,^)RC_ZKRcE/TaEQ1DM>[BQcZ_b1&9R
DMRN)+HY/WJ<8=45UTZ32K]d3^ZEXJ)/X3b2V3dG1JX=04RHY:D:]V+\(O><d0HQ
<(AHa6MGLYVc>4@eO7f+EYZeKM\fW]8:eJI7[-)74T&:_g9Xf@Q]8(:140eI\S,Y
HP6_C9O9_[B@X0=O6QG0B/2Z)&gBKMWODaX5#>IWCC.TJb@Z2GU[<;)GSL?B^A_=
Y2X-e#EZ?B#OKg12c1>L\1f5NLL-+_g.<E;-3NeOWWCdVX9<)M[FEMX;_<C2(+8D
FbT8<<D.=AGRTS>Q.BV4RBVNb?_42;:<,QD_,H7&.,?df[W,M[=231DA.8K:>:(&
.ZRJ31?C/O?48/R@5]0fLOH=1cV_AbTX.4XfFcM;19EHR?+eCWPd7M.L77YOcA/G
K/,TI5#][P1TU;W=AU(T?=,7,:=>SHTI04V/UH@0QQQEQdH,9\NZcCa/_13M,,<^
g,ZLZQ<QEFBK_7C]ScOFI.[B:_da3/)LZDbAXF,A_6.[gR[0EgFaA01D-NJ;(?<?
fK-d1.-@c2U7fd=2g/AZQG\VCVSTK^c2UJdg0B[=GL;OD=7T&_PF049g_DV^([IJ
Z78Q_M5QNVJ9YM4A8VW^LgE#V1g&bD;]>@DWb7dL/Y(&QO@/_XFH;Z[cYb:Pg)?R
bOE.]_VZ.-F2@:-gcU0<V4]W(/Z1?[I?24QOBe:?NZ<aU^6^\81]=/W1;cUQTC1;
P_LM/792&;G+4d6<P)J8Z4)6I>@f9]>K7&]Ice+^4N3LZ81J^_J[6:JESJC[F2\6
W01#+LYKI^J@Jf3[E03W_TG8,A?22?]7aU0Jb\R-PU>e\][YPQ[b(;QPWJ.F0,fB
TdHV[fJ.e6.4[7cgBOa:52)=cE5C4NQU_YS)aZP&SVa@F,71^<JA3-Tf\1GR&H;g
963+@]/^[eHgF5M;52B^&14b4bY&57cSA38D,.7g5LLdAF_8aE9ReHaUWbRCfJE^
A;CPR4dLUZ4cBc7\RA)X@ZCQHb5C4YJWYOA7+2ND+FN-R8gBdJGN5-K=QCET@0@#
+=]^J&8-^A^c/Z59KR;H>H4/W0O7R9WQG((^O=a];B.6D-^H6OD)N>GQS:(2b#8/
>1c<6B(YD,4L[X,Ug488HA?DD.NU6/ADHK0@RQ)Ld\1T=3)Rc<WPU&G_1L4PTgT.
.Eb)<dfJ?B_4I4K0U0P-DZL\B_efF^cTH]Wg)@&_bOE5LJ_1CQO\N42@ZHSRO?/3
c9:SGO\(eTQaaCE]ddHPdeADc7QcN5SGK:,EC_S(G5F^:S4F[_R@UOZ7X6<U@A&a
-_EO4J3gHQLSdX#=fM[eTR5aXe_/5#7AEA^_+7=aQDEa8OL=_bEb01:dc:IXB5fe
XT^P]874O[1K7aP-.M(&(Kd&gMd#B.f_&2^#b/?d\=e)?TJY,f#(L,]O-F)(1+F@
/49?2ca&E#H_/KZY+GO/0&5MQ.?XJ>(\,JQa/8OHa&56918P0MQ(CR3>aD/)H5ae
>)S[UIe<Ca]:7K;BL4f3-eHMJKPNKABP/D/c,Wc:+&))R9=@&D=I3@Y)bc@Ug.F+
D/H,H&@2VLH1&DQVNPCYQLE3I.-?TC..9.4g6.Y]])PB9[c:V=:a46Y?:&QYEDTg
=1W^4]U9>U4D#QCF<M?QIeW]efcNGd^@JFRAc3]+HD4E(BY>b:O5,++d#2R<G<N7
#-gMR=Aa81_6EXO/O?1);4U8daC9bbEJ-//=,Rd@/B9gJC+XI4.Vd6#^9T.Z9eK_
I/5J8/I@eYKT.Z]-Mf]cFOM\NJ4M0OYe6A)aOL9@f]^gHN-.TUb#&&4=2SXN_Y+(
[1L=TM/8TdYYbXR:0AVN-L3J^e(00A(V5aY4NeZ3Y0E\^9,;A,F26+F0?Q)D9Pa2
AIZa>J<]R2PJ_>95ZN7QPac:80)fW7X,bbeO,:5<I&8NG0,>WcXN;2U^d31_6_.e
D60K>4;CE0V_(2(JR4M/_feQcO=X<A-7NM_F(=Z_gG^<b?GL-aJ^XYd9(=7[>E.4
;\[bY4;/=3CSPE:(;1]A[95B.UX-.X)SS/_S4L/N?WNG=(@H[,(H81RaV1@.9ea7
2(MaSWa2NEf/0:CVKf7cN.O0M:U2eI90T(6R3XUa&L\-d&#]\aX,W/P>5bM)?Pf8
D8Oe?3F7,DX5EU+WG2BH<c>b38L\bJdLd+R0BIfX>cP-.M:+@6ERN#He3VH=3SgT
)<Q0]7aaM36Yd9ML<1ZN-Y-9Z.B3X--0:+=0cL8S[2_JO2IW?g_1+HZI_&PU()57
^b?,N3)MW14E&8791B6;V7EUfQO(>7OBFWI@Ebb&Xa1F3[MG7AC/7Je#IC?96)/)
a0(-7F@f6T?J6YZ&F:@55^(D_b;;+FD0eH4;Sb8ca5)BNWbY4ASG6N2La]WbaLH_
]_+<EadGPH.OE@EE\_g[<;YPG4_E\AK2?LAD_I]-[.aPHX;M+B9EL.Lc0dVG/FF]
E:d1&?G8EZc/CMaY,2<Q)d4-Z,GN,&Zc62KTF2,N?Z#0S:b#[2>#ML8V+b[#/AcI
#LEQD9d^(CX^C/0<21L)(@PM5PH-&<3_beb<-05P<3UC@6L:-JL/:Xe,P==6a3\]
(e&WHE1Wd6g<-,\AQ=dLK>;Z\J5DbL;<-4IVBC[I+=J(bZ^bPNK@gP-b6(HO[(Sg
b_=C[cKT)?4456BU0&1?F>.gT@FN#1OE6:[=UAe;IbPgR;)#:0TPO9)KD)88-948
;T<1?[7&AK--+26G3E0.c6:CJRLFN+c+UgKUE60gcdE-(f^C?EH2Ha\g^?X;+g/R
0,1_/ACC?A:0Q&R5aE=D(Sf0DeYf2f+UFf_KNNcVQ3>RD?H#>9a,Q\#F9O)@W>;(
NIC</7J0(YGeW_Eb,AO,P4)bGH&(c]HIBK4U\F]VSVM3g2;c=-:WMWXIN53V,;_a
6GXe+_G\cJ#6^<,.f.W60#-><3L7;3&\&8c&]<d=/@KW:eE42<<N@E4CdeK,E3E6
@\4N]AFTVb>G5f-&&18(b<CRKP.1a\O4TWGec63CIGHD<Z<FQYPP>^X3J>]>7CT:
JS\5,XAPfbLeY8S;.LVgP[e#_(ObY07.:PQ-JYYWSRRUE)LfC/6W3K35C3.&9?<U
b/eT:[WH@KPY)MIQ;7GcgZRa?.6gXN]1RUH0JSC5TDcP(:E@e#:7dD)C-&0GA3/,
OD6A8XD-=6Z\++F-D5bL,&,=,K4Y#0E)E[dT@WJ3LK==Ddd1D:DI.C)B/^+PC.g[
I;.B4b)OB5/^c@NBR2=O&=UbecP6V=C0_3@6S&;231=S)L=QKCJLRL7E/c=XQca0
DK>>[02R+CKJAc+)#T[)&1Sb&=CL-Wb(2)EZ/0(GY7^I.BJ9>.OQcKa<+A03L1^N
IdZ(,ZW.C/3,aLI]DD0c#,\P&JFS)RTNEWZC3GbBH_FMRa9OF9\N^gg?M0XO,>E?
<ZX.=@/.CBa1.M5Q=&W?#HcRbV5+I@T4UE\N=YPJ6-[X8;a71a)/<QY]H-M+06TL
8aaK=S\)Qcg_Ha<5c_5_3PXXe+/eLV=9Aa_\8N1[>R^.aWW1O#]=;@G^dC+KMLW5
fI<gR5E>9[3AJc>De06I+5,,Bc&2A:,BbWXdOSO^2:f>4_Y5I/dd5ERXS.U=R]dZ
U/R>]gBS)DH8dE[>NLQ(Q5JG0cWK2gQg0JE/:)<;+dLbVD+9X^F80JUJBDLa2V?A
_J?T\I(]bd=?cVKS77G7\Xab#@&]Y[/=)#BCE^<GQ=0fe8G+?Oe;<;VKA_H:]Fd\
3+g>2J0WFVXE@8E_0MH.F@bV.+R?.\5+])SWLd&E>ID+38K?663CQ0ZR_]47aMBc
3?JgJPWN>FeGL;>eTF5;bH],Md#8-6#I=M<?F\S)8f\G[S(eFGN&@VO)+B>W\)dT
.#0G)J4SPPFdT[F:+Ce3[?)0WK&a2fa3AVI;^<A/TeeODBZKcK@<DM=N5&OT.d0\
b[&#-DIB+T\E=WF,O]0aSJY^D2W,a26MUV[W@VXXHfAJc;[Qc^L&)R#]S)4AK@R=
>V7cQZPGdJ+X32([35T(\(GX0XW#J50fEUD@VY?RJX5^G4RDfUZ@A_5HQQX1HN9D
??,1]EP);U7GF1(XY25YGg0OFfHBEVH<^-V1G7,=QW>N36?K;/#LE^#PGX:4(RTX
9)+H7H6,)aE37KeaQJ6_fH5Db+g_W/?TDT#8EP>Y6eSG=LV#;V-/IVY.CKV7TgJ9
LM?cbe\6Z1-,Eb;VA+RPc\b6#T1_5Z=PQLeL-NVSUc]f574g)[=ZF+HeY\=+.73c
,5Y_d-5HJ80C0e,&Q/^RXd2+HT/Nb9,\Mf.^K4R_L1(a5J.Q<GU&[382]\RHZ_^a
V3d)N_P9?_KM](PfC@?:[-GE,e/)6+;1LZ]AS\,+6Q,HA:O]BQ>OI9?\?UaL;d?2
?/6K&1?W=dFZTNbH36Q=5A>4@_&.YafN:Oa1_,e7NYFZ=@b1N_fH6bV=1f3O9B:C
e:412@:3G/3B^O/E6RN[1@#&(_4=RWg6eTL&)gXO#0_@^bZW:>2J)WDSV\]Y16CY
:,Z9&(-U>YX<fNPP\O5f&SL78cZeDYCOE6E,PLB?E?]3=Q&>D\<Zdb,&#aC@/WU8
\XP?BM);5E1BX<:aPc;]BHGI=_I.J0Y6RG)X&^@\McSK=fWbK=.&_P(Z4M7A[JgO
\D2[7YdIY6-XW?OHLb@&:L/eQgLaTN],I2N^/IF,3_aWFgTMHf?NHQ:2G=,Z,aP(
KEeN:\f.S-DL:.IC1>M=a7?-#\D3(KMUNE#=D:5,AaDggKX:7?G,#c.MJdY_43/a
=<B^TCKXW_M:6)TFACReKd+4(T+^5DTWX)X(4XKL1L=ZFD5[O+FVCZB8eQPeY,&#
4cTOP)UXJ_->-SL7BZQ633X4D^^,1Wc;,XX[058FDVD:3IZN=E)FITOaW[:6LPFK
R2M1^XeG@.,a9@+^JT\9#GeST&<CZZB/aPgf5e-C]3Ae?VcX6fDMbG_P>Z#4e)MP
><],5d;5K6a0>FHL?e.;a#Y>fEQAdQV^DI@/N.^dDd?YO#&8/7;baC=(ccC08e_H
JO#[R@+IIN5@Q0fLC6Qe>\F170NQ(Tg>QWd#YU^eM8L/&/g8(RQCJc).LAOS9CIB
-/+W5PP2()DgG]fAEfY>f1V60Z)W,,Z0/#O786F:JW?L\c/SgXf?SO4A/TK8R#0M
PRYWg2g<8M7H\Q?R<g&9b+I5QIY)7NYI_eU66J[B7PYBH1bW;aIbCA:/.@F4_BSV
+.2HL23GH#?4(6V0Y&N^6)6YO:Z>fTH)7DFXL]Y]6Pg/9W&?-TQ4O2,=8NAD]1-8
9L7a-#eFP]f.ZaNN7>6RD)V2DXgMA3a+(Z0UE1P.]GOIOD<aN.+/#ZTg2IU-VW=]
9:RX>,f&P+(7QGU\4,&9aR:;.bY66,K19TdabG(LH6QF&3=bT^.68_eQ@fTac[&D
g(6U0K7HWV=/6(D7/W&9+ffNV1AbCU@<9<d@Y>Hf@8A8O<ZQa/f+LL0WgC43&8=F
?N33;P[=T1ea2#0MQ8f0)20UVS<Jd+)DdWOb,d3LP5M)3,GLM(4&+gL>)(,0d[\1
<:4))?37B3]I1SfU6@>:;RT+WN2([=9IcVT@6_eKR9T@>+&Z1\Q?^TIM[3E=?YK3
-cRKV>6B+7+[<IN6VG8[e>,UXJ;NRg:0d>f+Z#9,3S(5]+GBI8=&M^Z^9e\7X[0:
,/NA0Q.&/aI<2TF1)#A6:[G5>f,N:GWM\^><MEE?J&L)FZc4QHUMZ^c<M]BPQSH@
3CKLf?&&CZHF)MeS71:>Q^)DP#[T_I]c?J?_^J<0FOH#^&f@_(L,\@R52FAeM>2O
DMbdV=CbSZfZ):C<KI>5N?R=J/?E96^QI\e_K<Z)AE\cG&/bG[,7VMc&ZBF&>c7J
(:7d^GT+5Y,cVg=[[D[dL76:JHX=I?6X,K7U1SQUD0@]1G.)CB_)<BM;0-1[8MSc
>VcG6<(;S1Bb9,^1V8=(56F2R&PYRH.S-R2Cd0(Q+4RO)Y-T/=Y=LK&deJ@)=726
U8B((H51N53@MBMc=g>TKJ.(Gd&LJ:CeVbDeCY;>:/E:O]FFC^6F^<cH4WUL\K37
GKEZ7)8?#fBRA@ZK9KO1.B:#IDUd:6NY&Oe2S^c;#80QBF?Ta<)UaF-69[+SeAM[
BR1L8RUUc6..4Eeg?9/_V?PdD;f=S3<#K/[.e6QY/N,-??GKRa7:[G<-UOdL3-^1
B0S6\K8?GCX-cV.[dV-^=@/H+_c&M/BHb:X]_CD67-/HQ=c<=;JFY/N+3NfM[Y4/
Z<YNM8D&CZ],D0O+@F-c?M:GaUe()HVL3edB,?WUPIOP(0W11=2M&YA:7_CKIQ5F
H,=?(gZ6&EgW6.LZ[LT>NA2O]C,BN\#DX=c,]K],4:7[=UF:Y1_cbW#B^8TUO:Q5
-HI^O-3Gbd0L^D\cC=(IbeB0RR>Qe12;Y2L=W/Y?70#e,Q[C5TGe<Y-_L(KU(3O/
b8gZ2c&]5e_293OYXV>aYM7_,2eB7d@f+BTd<-K3].N#JMH3[FZ=9TB,+Q4/F0E5
+44YMc(..I.PDEN=XU=7.0-5FYQ]8PQUdUZ7W?W;fgXFA_BO_bU)PBaI.a-;LJ/5
]?V/KC)-=eJ@fJWODJW4Q0aG[FA^\18@VgHLH_K,YeYd0Z)dL+:a7:c#[BXC+R[S
@fK[UDZXTHQCJ&BE+aX0Mf;dV:Bg&H8WN+dE&8Paf#&O,1(R6<QJ43V\fM;PD&KM
&0^J+dBd,8T,QQUE@U&]<,6<bL>(T2KFa=IRdIAOO#JN,[AOX(1cab64.WZHQ-AE
9cHJ.7VW#>[TK^],ZX[5ccAGOUa/d1CgK&HM_^PWfV@1ISO/B?RGBZD12a.X4I9=
U3D3K(W9BdIS^X6g-bfD#53]afW.J1OLTeAgZHbSXU0fOMc_4GZOO8MZF/<f=BA^
UBB=Q-D_(WA\)g>F>T5H#9.MBdUIC\a18+XaV^Jg9C,EGM^F4\dcCOI6=:SDbEDe
U>CY(F>e8;=F-E:d\^8a?-Y:^-g^2AS4cAKG/.Cb-P-L7S+4XH;D]P<bH@=JeENL
/6+H&XF,6P&_YPSLZIGM\M2JSOW6Ga[g6Q_?I,,fUST9XdAQW;7Ob0>(^#GFHN62
WfHM+DG=DB&:./]@fSbYBga<1QXMN2\\g[]:#8fJ)eQY_)8^FXdXJH?IA8Xc[@__
RWVfE(b1V5C)Pa/H>E&<)eed;S46+G1.NWLKc^EWYY-0[0gK9L/Z@JY47?&E?-^.
VRg4U0F,RZ9B:_Xec9?.=-g@^&bUdWV-9E5J0R4Dgf9g)=<H;LD8_-2P==+A?0eH
7;]F7c]cS5:F45Q)F_M3d)T78aYK8.0L=4I<X\2P0d63-5SHLL0\NPN<H-Q8O:,M
JJa&eN,fTd]GOGA?<HdF>OWRXXD;F2JO5I:UdWa1Q2NH=@/8Z_A^/OWB/#,ZUg8I
4PI9T9G]^^[T.-=QM=4;:V&P0AR[G>&AH@c7E7&f#GbL+Z#8>A=ZY5M>_V57a+BB
3V+7=Qf[>/]2U?Ic1Le.H]3W(d(OQG&B=3fdAdL_^#<^@,E=76Ve-e<-/5NR?Qf#
&?gE<O>&B.3D:MCLQ@@<Z,83M_K=d&OAXS4fcL9UJ#ZTJ,HF<A@PN2YLX=^Age^W
AbJ5R(,\McM8aJ<B,4(/KXAe&44<1M?@S60dU?CZgU&BO5CcHR?1eAdJ]_E<Z>Fd
UDOe.a55VK\;=3/c_2bg=E(ER5@3FJdeMbL4]^T:1J22V7,>D4M1S:Ya/GEQA_B8
2W98AegR9OCe<^H)0VaZQa7=&O7)cP.&=>C8:<UM#WEaKRM<O=LZ;0gM?ZdZW[fN
5716SaOZ@+#Y(7M98G],(OFb&&bF:C&(.ffCYIIMVH@-H@(:/Y0LZ,=X9aG^;3DR
WL-e^fBMVfSOPYH0B9Ve_^b.0XDNH;>g8]a_6Uc<HY&B6eaN;R;c[[b?NMUOMCc.
UY;PJ6S0b&X[K\\NJ[TULTV95]+,7+IMa/Id:J0,AdL8R1OaE#33LF2Y^2XAGE97
DJ#IY<=@[<>VOCZNGU=F5+UdVG+B4N_YWX]V/SZU8V:LIOC8B<0JINZZ]bDb]:.+
>COIY3c];J[4U9]Z.QGcGDD:^9;U&d+,/Y4RUG.9M+]Ff&5NTdS=IHDMWY_S7TG@
PaP@(c;e8A<+<<^dR\=A@IaY=SZ@-+RCJ5DA+C/UCJBSf&9f^R]E<AW=d<MWNQd3
QPZBCa>0-L)8dI3(bDCUUR>[&SB@dB\bVI/a<OAgc=PSUP1#O/:6eU5YQGJ5]e;g
IW8W0I2G5=Q3V\U,F0HS=]c/M#/;eA2DD:UM9-E@gBBY?RF59ZO^a_d[B0]]fdYR
\93^fW28EdAd=N&0b[VFM)IZ/@#NSV/4>@EO=C:<LV(8^Y5eW,M8)-&T^I\ASLNK
)Nbg0O:#Z)Z&^K5fS#87(^Nf1>LMRX<9ZI^C(.G>@SebN[R#Ucdd8[cJ</52Y)#Q
5Z.EF5+[:UX@SN[IL&@Y^F/6U79dEW8&BL/bdWBT)#1LH[CB&O89+_&1-?E9Kd=M
X(Fd<7S<faEffOV+]O56]+.T2ORVR\dSS_Ma0E^6O^_T&9,5cV(=#EA@ZKcR71GL
_DE2ZE,U3PXB[aR-dQDe),GY09O0(ZRb-W5O:^CPKPeEJ?[5g;S??(c;84>cBV39
P(.::O@/Y,?H-bE.WVB0H(GMeDE[c\d,WPQBMC(NCXb2H5E>Z139g__18J212L_Q
7#6(O;R#EFI@:Z44B;LHQG&/,VFa0a4G[d:Z7gFO08(V@M0>9XJZ@MR]MaB<<bDg
.5?,Gg_(J+P)/BTE+R0cDKJ?MSIQ\g,?UW@<>OTRa5.=R-2:a66F4.=.Q,7NfZ4;
4KUG)>=P7J3M02H6ZZ<X\?Zg)84-VBa7bY&FU:TPKN7Y==WIO&58:7E2.]BLFcEg
I5cWICO5b+T\OS92P[]KWd>e47(C93Fc3UGE_YIXE]5GQYf0bP=X8SCg#=AIYDU2
f:\0=,_WbIc6F(CKdRLb)<bJ^e2LWR=V^7=L/.VU@V77W4&#dJZ,HSA]KRCVERQ^
N/GOMDQd<0FJ\TZ@&T0I[8@NDOg.CW-Mcg2(]NRP72-I)JLD-3K9M[Y&]\)H=Y+5
;d8gaK/M-AFMO1XN(<_W(gX^8?V)?JB1>D,SfSWeT?+_E<+;g>U3L=&=_J9B8cXB
ZWa];8OA8+.Ge=7KJB<HE?gNKRD94VM5HP5KGOeDWHPA+826PKeRJ&HFQG^KE-T:
F558?I_@<3[8SYB)@MOR3>8TVDO6Tb6GgQQef>C^P0)8I32&[CPdM)_VV#D-g<df
C>e>[9N8HPBZD[<4]_9E?b0Ng66@X1)c=G]2ObW+GS;]G>X)JO-)[N@^F2ZNT^aJ
.(,.cORV2CO#PN3Y#XbFCJB4158B>[O.JPA_GE32c[22POI@,7UQ@[V#\&9/2#6[
-J8VCgNZTKV<=)U7c8WdQ0LFScMCSRT512]P)8H&c0f?WZGIAKR>?F4<R,;6X88\
UVLIXE])g-E@NDYb@/0PU\6D-)M+X-IFML.A:Hb+e?fE=dTRZH?+Vc2AYT)7.KCc
9S/&Z_CT.,:../39[._MRab-C&Q>E(6/7N-Wf[>dZ+[Q64Z+_QZ\H(^3a[52F6a/
;0>F8[8IJFA==]Y8,Q\dWI(TM-[V+^=^S10VJF94<WaGP^\GZUN?e,EeHGKK&-OQ
<C?0BOb7@8X>JIPA<3O6.H-=aS9?=TbQO?L:(AQ\JPK[MO<ICJ]3gCIYMD:UYXD?
0X,gY#()GG-VIb^.[f3NK7\)aLOMfcQgJ,>WRC==Lf>YSW7HY>@.QLeHA4d;VY]-
-7D2/1@8Z@+S8(&N3.D)A=2=<)JfB;Q.LF0\F(S#dcdH5TdNOTgN<aC30E@-3N,4
XJ3K,;9+D?c/4W;IKWQdedCR2GMGUW6?DD0ZCA<[8I+[IKYbS7[S.^37^R6S5\<J
UgPg,^Jb3ZADJgPD]Xd?8J[c9Zd\MF_dc[YEg@ZUOIU@9dBEQ,WB8@J#>=RgAb^M
WZM/J4WZfXAb71JTF>73Xg.e>WU8+c7bW?^F;_K<)9CS?IOScSCe^Vg0FIXST^NC
d1O0I]3K-E-8.BW0LZ(HdDS7UP/Jd?ZbV;\8IMS8QV?eJ8]&\5a&a)Q>2f&40,\X
;Y6:FHfd8O)>,C=R]E)PN^JaIDOf>(QDaSQWYRHb.M1VeI?QYc/B\HUS&bG\[Z)0
UaX18T=/F_&CeSTG&B2W+fF^KTW)f2-Q3ONC(Xg9UC?U_?W_[5)O.]3_Xcb(MHF(
X[QE8dH=KL;R+6KQf;T>5,I2]M#fZ9@SUFLTcH1774]9YdO0a2.aL[ab7O-UZKd#
LC(af,M48;\;IOO7#(A>OU^/e+O=\a)8=<Qb5>e@CO6@^W]#SJ1TCN^P:1RWMC)0
f/\QJ>IT6Z72e8LL1geb/f>Y-Z2Y8.EdW=/4J=HMM/[_;43.Q^/Z#BI09dQ^,LM\
b;-J0UE1T:U;LM;/F7,0UP,(R<;G&,_E)VM..2JL1[eaA;UcE(TC:@1gUF84ECIF
1WBKRMPcfbCIQ9C#]WD21VC(,Y0GP)?GA8;^.OLVgc#DEYR:/+7H,U(&5+2RFg=Z
g;)IBWJPJNGW94D7I7V,YEDcE[;=,@:+]-aC\FA^DEC1[&\aKT((Z1Z@Z2N+YbCY
.UQG+?c/dSKLZ+/b+5)eI?>TYfQT1;XP&F-<MN:]TM@XARcH)7SW5Gb<P?Ab0^4C
LU)E??a##7WQ]@=K\A_K9+7=P;82JQ_ILb1OF+Q?;OOW[9UP@+,U8(aQPH>?O+#7
TS:I8bI/Y@V?(VCP,HD<F=CLTGJAR:#GD)6B949)]QB<V2[]<YF[KH(E-cNLf3F+
ZWNECD]CK><bYVN\9dQ@/40]H=)85/@Q)<Y,1/C7L]gO4/\NU8/eS]]b,F;3I5BF
JZ#1Fd:]?52c=9S#g/2H7^A3CGKI(:Q3;8;X\A.7<7a>e-aOQaF+(-fCFOZR.=NT
X<6>^P^)VP;>@=DVe_VQ0N[&d7bY>Y&/I<(1QObeT7\S=0B:]S_KNaVR9LU&B06f
?R?FTD)cA[,#HK6KPSMKXB0a2F\.X-0P#9W@^LBL74^DE;c@2C^VC8Zf2a:@\Rg,
P<ZI_W6#F2@&14=N=,3?;7J199ddHPJ7Mg6<beUB960[Sg4E9]aL7XGeVSX5Rf?@
20X;LEe)B0ZT<>cB92UAC->HcJ7)e-<@AeCZ\/\L6GNN#.XW8_[NG#4C-:6K:=.^
;\+COM-PN@\S(#e-gOB#A#J=[eH@)J3e_T>b)NHM6XHLMM)W9[=TOIUZ#R=W4D@9
XSS+7fFL_a__2L9AV:T;/9PXBBf:_Y@\H0FB.,U21gFDI,D=Q>?g,]81HbJX<^L[
<A<caYSYI7P-@&IEZ7eY91CLdBP+61UB_3?7afd#FJ]6&>-1TQOEXMN)\U,6R;5@
K_\U+>L1<O7g\(EPK+#<2fF3e3T_A9&TRG8FAc5WTX^4?&/BfSB?U:8]N]>[#OP6
d3;=\:9]I=FK:FdaM2<#UI:HP+X\;VMe;O\RQ&<@+EFG@8(bA4F]U;AIPGI<Y@-]
1P17-S(4T8?\M6a]M#8Cebc+0,R.&_fO/&ESO_L&<<Wa,+Bc&a->3/3#:5[&_UK;
2?=5W4bBaMGVBQ<.;fZbNR;GS5UaIQDVCJ)Id9:U^YN,?UDaXX7Jg8G]B_1g@WBU
O0?FY/?J8::@[Z02=BO2:>JF^(===4/(A\O1S1T#=+&SB9_1DJ]:)[;-:F?DD^VT
5Ya4NI>VPaaBPf;@RX-9ZYfRHD1]d7_fRX.G=6D,.g7IKYHJM^]UP3Q21P9]2.#G
LA+&eeSbc[OJSNaA<XRYPNM[@)gAQ=fE[12\.WKU[0T2O1A[Y&]VcIX5b>R]1B22
#:L9Ic;]Le5DQ.F-PVI0\RbdHC_CRR>GU=376V)f+TNVQL)@2>CSRfB\KC9B7QP0
ENKc0LXb0HVCf^\_T=IQ]ORS1(1?L(A+KI>dCSK[=#9U-E0?;4aB7(4\B0e)OP3a
G.KP]e,2&K87=V.4BR8P223c8Mc(&4_@/^g>L2IIJ5/5AZ,:X>PPfYUf.U+P@7?O
7=];V/]LZN79DZH[cd&?Z<_3NG@)Y[>##@\Pa3cFaAQaAJNQ;,+N.6a=Q;_A)I[A
W)XaIcJU//2)CASCO_XTagSdK;WcTB<S>_+?#=P3gTdd8gKd5YBP@1S1?8J-;gE]
\^(aGQF<fE4fLc^O:5JI7V@C/\a05Q1eM,a=_WZ(-5f=_cM,Z,e.Gb9@SG+E)?OL
GTAY_1;ZR#K-Cf1_VL_5#ZM@C#gP1^4-#1+.eZP_A([]VNGU5H<#8-:fcO0F&K?=
#35dFG5WA)M\VZG:)<@Ua6WKLa3cC#8EW-)(\()ES32(::,(M1WS_g8DMCd1X2Hc
OER3MPULX-8Q95S\5CW>2HB.L=QJ]_9E.9M9(DUA@0TI_8gf8T^LcMF/Xb,;U-@<
WE??6/#R:g9]Df_[b/KD>4:)ABXJ2:-C0.F;L?.](F;NF5W<Tc4\MP#G.3WUB.(T
Z6+Md=4@g.<JbdW,/W2-ED:+8X1X&Ufd=ZU;c9/;?E9M4QMf<9b:)\T;?>NPce:W
R]bD31>PB5c7^F.(Z_QZB.M0OY_dMXN@]G8WT2C)@6PS3),(fQaH+\:<W1^5O6eN
1A\SH32;8K9=W)ZP?^cFTgN_\0/gbDA<]VX9Y1O8EQP(W=>N[JZb37LSFM2c-P>[
A_G2e[7(0EgaLgJ-dP,eVfW6dVL/NAI@GL,2V[PPMcU&6gAJ-VX@a7IZ4\;UfNVH
#Q2T@Uc;=MSID):Qa<+N0BPIA[)S#I>H9PRb^cI[U4+WKM0O)(?AMRU+cGR81AG:
6;;=M4<7gYQAG(c8e&RM^c[9>YJ^[],(V&)PV.2QXK8KNTb<ecD.7RUJJ:BIJ)3-
e])NcWD/?Q;#gA3?]_,;WXBGYY(e@gaM&\RH?X7-,CZ8g/GY>,GdE<=^5&0e(V^g
_NCaXM.0^68[39&6FR&DJ;gRI=3-H@D-TZ3cN#:3:&/_>+,LdZVZ^Q-]X[TX&,\L
>a].>A(/-cH/T]2,<0=BUYe>6Oe]REc>6(B-;^]\TUX32gZ@BgG-PRF,>aQN[YKS
]T,#^4X#5NPX-=1ZV:[bGTWBV.c0)+UC4)FJ5_U\1>4UNB,Tg^<<PW7J@2&SBD@Q
<4<BCA_45U;UJI(.;-(7,D6G?LNDB>a_0\A9@[;I,JQ0eded29:8]bHbZR?9#[MZ
bQLA<B(RRdS=^N:;.a0C@=RP2K5bE7_)6]@K?91ffLgP0AOV;6,F2LW^(_,9/^>H
c-4gL8Qf+2H685IO&;2ML]=K;S)<f1eSF?;R.IK8@IX#IZb+cT&O\XeUE6.-NDdM
a<T.fd8AF4NJD>Ig+9[4R2BUPgW[4CM=H+#6+QB>1:4Q[bP];0dQ<J76[7O6L#Pf
3Oa/&Ta@#HQUN^REN@C(11cND/J#1O_[BGI0aL@A93O=;6?,AMPS;&D\CcJ-fa=_
&4>G?()N0,;gB?d06(C9/+U,a#c-?Ja?(Z8_4L.LEdU^c2Ze9gJMYTU3B/FQQONF
Kf#<&/XJ^e9d],&4NO#eD>5b4Rec7M9K>O&0b-#ZWB[c)I+POV6R=&M?F6_bAFV[
]b/0BIe)^5,PXHU(2Y9+JaH:9QYYH&QSY\F:7JK6=,HHX(Y@8E/9g\T_VI#(36^Z
^48B&&9#a3>\HY+B?ZWTLZAgF&R2^LZd?eSB3CY-VD0VHE)Y1@eYC=UMBF@<\A:I
05-c:6F.C70Id2/H?&0\^7MEJ]F,BU:6N\@-f/9E?M_DH-@U4\^F7B)MGg7:8/W(
MH0C3cI3g&RR4,&?>a9TFMD[=;a^f&KOW-)@I]+B+WV3V>Y=b_,C_:)QcdRM3ZV-
Q\JKI3>@I/+X^2M/Q3^\)N6F.+S[A-ZGP9^eS@PN;+-JM?,[EMR&_e4SCYELLWX[
bK<Q;3aFAc]S4OL[Sa@MM37]3V:=HYM3=@H0_-]W2)9MdZC>6Y0-K.Q[cC7<F<_@
L-,Wb)HaANPCR#dZYgeD^=:fE\[G+_aAbANO@PX38ATXX2JP0>5XECQ_;dAD030N
@\Jd,ZYQ.GMgQ>5(>,I4[YE/_edd6/6;VE^bH<MV?2)84f:#,ggNEU&G\Xe7<AaC
Bg(DHK>6##NL:OLDf3.<f\.?ea)A]+E+7g7)1bNBNbE?3<ZRc<D25FFACFP)D(T&
P5HOCC>@e<e\6Q+^JU>3887Q0H8NJC<2f)9C_QfSD[/GgPdZBID(;BfU>6OQD>(?
)PW,@/-FIA]J:W7AQX=@@)W1E8M9A0T5GU#)HKN;A/d^dE;RIWUGF;]4_UFQM<9F
H8&SgJYa3B.HIA-LX@f[L;\//_K^3I(;f@+/+8=6V9c3[?,Y]#=R;>]OJ@BO3e+F
[10UbId+_17@LBcQ-8=JST\@C>TV4^>.R1bM14VXR]B<7QESTB[=I[+]<.=7?YGM
/-[f&1SS5Q<Q(adO:EUX782W-/[_OF9Z0e8F/W3PI6A;0DP2MON8M((BRdOGQSPd
e+UDZ#Z/,G08:YgDRQP\2cAWXc9;Z/U=6\XX(W<6NL.g4B+#V39]UA8+f.f0KLCU
&DB[HP=B4=-U.KXE/-XGYgV.CQ9FWPB6g9JB-LOS7\DZ[&YN&9Pa2M9R4[9XeUPf
-4/TR69^.2dg?XG)/@;Zb0/G:X7^UOeeQB&=39&c->1B4e,WNQUbd):VTK@IN_O@
>#@)X6DLacba3W0SB66Z<S#.D#.\Qcf+48A4=1OeO>>K2b(.S@Q+7XJCRYY]00J/
(9ZKS>\MO\C]V1f:-D:+A1?^RVKS3?UPYOY6,[2Vb5]3P49_@#.O8@cN1V)(+:0?
)Xc+I5:6:&5;:BaZXT+B1cZfHLeE^3\JeJWI\bgH<NUR>+cPDbB_RKT.GCa=5Ze2
=XX;[@D2d.&aJ2RYONJ7[HCTYdE_53@E/&83Sf<OaOKf3Y^:5D.3PPSD5FCO-B^[
3F-@7a0d#KA>K8PDGaLbM4JaJJZ?C:;7P1UTa&6Q2NFLbHNKcS&f0Ka5[H8[;A3&
4T@Md?f8Fa#A\./9E+T#&(S-@gd<bECFDM(:KP1]FQ-8Z,=VW@3>FEe@X+]=P1<)
YRCZdYTf5W:CLZf/8AePHQgU1+R#=)Q)]Kf)&P=]C8-MPc8BG1-.FfRPCQ2W@?=X
K#cORP@4RZ+c,<ZGGU0CG;2)M.?(8Q2)1#D17FA]O.]H;DIUW-0_f_7IWHFM[f4P
4I;RTY?C,-<DU4ZW^6B&fbMSeJ2d=&C#Z@0DHU?C,f4I(,ZJAGEMJ]&cXU5S?[X-
F\O.,ZIPVc[UN=V=3;2PG6V:RZ&cQT(6.Y3aQ,FE@.0.aVQJcPD>=(3:[FF9PfNO
fIRS;I1:[N:AA0XL;S7SZ?UUJO(DS:N?Te._87>4L\B0e9R(T.+;_DAA17&)N/f3
>IJW9dI5Q+gZa4AgD7B6COT4I2RS-Zb>?+46Y#5F]-)-_cB,NBL^NXa)e9:)GDMc
;+Ef0:MP9IXU;(/HH+\_TAIUB92F87THP1dK:3LeMYSf#IHY+D2T9LO7&&c5Oa^S
QFc?f9U:RF=\g>@1L7_5Xe=#K@W8ENEZ,B>Oa_c>)T5^]7A=@C3?5U;dR&P)YaFI
<gBKU741F0^IIWK(g0^0CggAA(7IDc(L(HXN@\PF@HK8a]L6gHf&Ke?2BR19/JJF
6ZP)?:,E8W)6g#GDRR#6RM/(PHU1gON;]K5F2-,KR7@1THQ3OPgV(9>F973/(HWd
4DX@P2#W-EW0-6DTU1C&eLeGVD@S^;IOFOfa1+9VFf,TRPSa6U,7g,/gB6[;cHU[
T1^(HZ0B:ST[YVAS4@&4;O[\@,?1ga>0/&U7Z6+MJBQ^1g&ZJa^fWIBL:9A=W9GP
g@aY;F-bZ0F.6f@&Z;C]4L=a-H@7QM[58(Mc1:[).(=+P//4]W0GQ>_M((S-/?41
Cf.IDgA5)N](QY>]SH2D5K094US=-OZbgP@5<6A(,8d2U/[g2ZKH:,Y9>aHe<gRB
Q,[/A#,>Nf:9RK\0/bWTJY@C^L9/RBUe6Hc\-2\ARZT..0C3c32FM81bDaJcaG=0
V2.L?GM2I.7HXd@&-@F_5\815\BAHd<[L[Q>S#V:W@_#3#B#>[M1^:J+dL63\8F>
TEd5T4+,daLa0RCc.X,ZD3L.=/;+]](P-@:H/XYDNDYdP,]HOb#F5_)2^/Q-UW2W
CBXXO21f1F0Y[TT,+X]J(ZSd,CZDDW3e,12.2JTPdR<Nd/.4FK\f(g7caK?FVD0]
TNT:6_4\TP&=LAES;\f1PgbE[Ba1a&VD^\-3R<]HRV](a6HV3<83>.8JCWJe0YD=
Z]gf:FMP;@[?MGfHca^LSPNDZ&]FT2T=(;gB9LTg5Z_-a(5A);EdK;1\c2L8\.Ab
Z:E-FfZ_6f^.P&d8ZGG4&126Q-8[_&>S@@2X^G=Gg)>J:Qb>8c(]UbDff=O5SN\@
;]ES,T-W,E3;LT>Q.Z_PEg&RgSI7[C?7c4I1)ZP+E_8-O9AQE.,:)K&WODEY:5?J
E:RY>=@\gL?^B7F^3MKW_VHbU]A.6_V4a?3:3V7Z>E)>().I>gM1XfI:?#O:=@3F
aP(^Q^<]?#cD[[G\We-F/H68(]eCa7(XW);EJ?,>ObV-E4>S[W,OaNY+cYC.EH0Z
-1U^;>E5WF2-bIEe^OGCUJF[CR\[?GbKJcEW(>W77J0LK?N>CX&O1PdZ4?NQ@>H/
(H4N&4g&@1a]5VBC0R>2G3YPXgO7[gK1.?_WHA,\Le91N=&,E=,@)(K^eVa]766#
_YT.#c6eVf8:4HG;]6Gda>]:(/G.R,RU9-5]<Ec)7N-b,f\CBLG.S1WP#:J0GVeL
NL(.O?W=)IGeE3OUf@RTTM[fJKOJ041#WbV5]V1](E_/J?1DA0\4^7U-K5Tf73ce
@)cJ5TPC-2Y)//#_a0RJ04gf]L+,)-@6B@,Y6B8Od6f_SW4.)8-]7^VgW^ffb0MV
L.J[F?&-G/6fK]+IHL7fAAJPT,MK@=7#^J)I=;9g:6Ha^c#NU#8\<Pa8\6X>L]gW
@gYLG85Q;(>D7/;A#N?dLP[+3O@YLP[2B&&3]gM.5.>&E^D-&[#3^1LI:#_(WRUg
edH>T4MJ4Q-T3\fT8?(OLN5+E<WaT<<CM+_)R^G_XFYf4PFC75c-XAd>>DQ2ON[(
T#8gO3<GW39^?@W:V7]?e+2-\L(8b&9=]I\EH3A[&1>6Y);(^KO0Cc<#T<\0>Naf
X>=GFb0^ZT^04-=0MLLcf--[4>_b62?N4.<bU&W/Fb8>&.;Ae^_C#H#E)E&2G?1W
G3O_6JZ+2>VU8P06W>7@S-;^Pe4fA[GMK]9=.OLF5N(G9HN5)=:a<4\SMbeS2>Ca
Jc;KZ]X96&4C8OSKF+Y^=6.POc5[1X3UI\2g(?_;(AZJ-?3:AT5-[]g&c3DOMD\+
7#)Q95H_;GYSY7844<F(+(b.HJ1L1bZ.?gQ^^5g6N-VL/fg5\ODcX8,;C[YFI^+c
9)0Gb=KXO6W3]Kf>Ig6fI2+KPI2UK?+]a8WM@K+PNXT>KMA.6Z5_@ZV?b_T12W]N
K/P&G<KC;_U<H(EgR.+JUbf,)ZW>KF/Q\Ka&/L\EZ4]3DE#/?AbLc5>3SC,O)D<I
8fLL;VM^:g0#JQ55=3Y;1B?\f1@CU68I1>K\W4&XKP<\KgE8L(2bO[4X[J)_4Q>C
@Ve#()&]2B<4,/&7M#1SOG[#T?6^3LDfA0:B4J_84171Wa;Y^^32&@XR/YG;3HEN
OM:WHVFPA#&.6J(5e-<WU<HE-M89TJHZCL[aPJD,a1O3S0L1@\.b/-YJZ_SIJ,/[
N7/:=_LI0N,8Wb;BH\@E>^59@0RQI#)F]Pa7+.Z/C2bYAZ[S+a]/&[7e-]K]W,?=
]M>=gX>BC84X1RF3)U)@Se9FZ2@\-=J/dS/B.L,#JY(5^_;[;(_R68f+@5(9L/OR
gOQT?O0K>e23ZLKZT=dD(cAGY\KBU>[4@3RaP)Q#I+O7d?O.E7[OT-UGa+bAb3/e
e(4F;\F-4LYZX=2\AWKWEQ)\>eRGTPM/Ye/Mc2NcL;>T]ge9H[c[)/EcgQ4D:(@c
NbX&cP?a7G0:-PQB:YY7=EAN#X705IUA_B[N<Q/RBa)Sfg0EI?LMJPS7EO)&5d;,
V:O.eCFPJS:XZ=1;DF-&0A<XMI#CZ5Z+:?WDJUES>+e@WFNS0/MVN+L50f^N^D#E
W-FGLU32Oge0)5-5bZ=MA-K+IY1c[#UU_c#4G&-]T_WD;(@/Ge=2+#(eROf[VMA5
\?bAG-]F#Qd0#YR/VDGT/&?@A6_eNHD,MRWeR-XbUWZERI;,;/0MN,TNQ;3&a)>^
^Y.B[_WQE4,TL9JD@<RMUYWSJ)&Xc@WaOQL9D8HS3<0Rf53OS5<+._Ef5+R18FG=
W=bB<2/7DZFR^SdMR^SW6S0D0>-HHOYVD&]6?LfPc-V^+.(@]^=78&c=K/=;F.]/
F8<)4G9^;.974[ICARZUA_]KVX1N_2/\U[?.NDQ:(A/<?UTT?U-]L&T6Jd-HV.AL
5_ST,4<7EU;?@69g]^J(e,Mb\P2<0)a#TgCLR<Z#e,2WS<&HB<12P;]fP]L/]3]Q
<W+4DaBg6M^_T)VI56>BF>(aX,#,e1\5(5->.7PI5)AgC(Eb^YMD30Q+4X@1Z^6F
KZ?F;)^;&&0S-]PK-9@,?^O)gLfYY?Kg/gb^XgdMGEQ:R357/HG3TSF6TMJ6K61E
>H=I2AL2IXW\8aM^6&<b#^+.U/&2E+V)=Z+;H=+8B;SDEP.O/e:>XK=a2FLOZ>?;
/fIfeBQOaYP1:45F#PXKF@T@F<@\44OENXJ46aMG)E:UTHZ<M[+1,0[)0dME,6N&
.^8#X^ZO>E5;f7gFL8>L2<5R5KQOFWfN=(#eWR=f7J@XO)VQ=C:.Hc^OSPD)aLBU
R0XYW9MeV)LHAA8aB)2?,8#8\9AI1:H_0X+U/=D@#:M>78D&[RR;B\GeA@G[XaYA
I+6Vf,f:R:18MRWKSA\Nb1B>\/Ug2,aZg&?HS+eLM1_V>0>C@]A76_\+7^Q38=CY
T]^LX.\cM(fD0HWK#AC&+6KJ4MNEN29&gUW;RIa+DYNGPdGLSe][YaU;1/G,H=21
)FEVH49@91F];Ja03P((0T(@7K=DXg[,+G\OER=Y:O>YbXM]537I+T9X\2+OUUC2
Z2&_c7E#?\[&b=LK]5f<X?9\/9^_<XbYHPG-AfOC4NMMW-DER5.8SZEd7RUJ/63G
bIcX0g49S7S[EJ38NNK)\fa&b;;E;1UVfP1=c[Z#FY_4HZZ;.31->RaE&))(H&W[
]W2>/W-&XKdHT.6GD;fWGT^<G:gO3T2.5b)5gBeVH>W,GWb7)#REOX:4ReAFcD^X
6T[LYVg,,@f1_6(QJE]<KB=WE,B,ZB>bCdaFY2LQNFEC1S4RZ/A0=AIdH0B9a_I.
aZ(_EAc:eACHTOLVJ:Dg-gXRQ1>NH[T.IX547CMd/SXE<_QBB01cdb(,D.\Y)^_Z
_+R]F=DXIG#OJFI25-\I)@T9c6YPYDU2YS3+5-[/cKKY]<g,A6;-7eYP;a-M(_a-
AD@<E1bUd?IIQeYBJ1.XLW7fQW0DC/4/>SMCWD#/Qb.W#X687CV676C:c^<1/AF)
MDU3dPS;;\fOH#HWV]YJ75O)],YSgGA,B9Y9K(8:>&8bUL<9;_HJ=]+aVTO5W,FL
aa6UYf3TTK>U;Yb57?YXP+Hbd+J2;KMI?gD41R&]^d/7aU0cbBTDW/E&K@\GFY-\
Yf.7C:E&]0IV4R.2I2T17/ABH_MY>NU89^[f?M&\OMEF]5/fggMB8)=C^V[DOBcD
G(F\>4Nfb#5L9RTfY5M=0B38F#^a7HF18BeT?aJdV<<^066H_2.:6FbQTcP2e5+P
B/IP+45RH7?>O/MIW&\(E,(:1;aMK3KHag;bOfC6IM6<LSb]]7AY]G@KD+U-\?7d
BfCR<R9L?\HA]_M;&]B7CA?Z8/EYc?L?OC:@#)OT?(#]N>7a#66=ZIT#a&=UE14=
_4>eFO&][+[R+>dIW,GO+9K2;[:1:5FB8?Y=.caSH1>dMDcGY/XW9fCOXdZ/X\<-
>H@^]Y<.<=YN(VYJ8(OdHXY?ae#78^[CTV.^f2/Q6S.W+S\=P;ZB__4R&DA\5U]1
UQGLA6A)^&C;C70e4<B:.YJ186^5#0E00C(ERAc1fUKVe=/&Y-FcBK=_,@8S1N#B
ETT?FfV&bS8_,dMM2_UWS/T4bF<:D;,.E.T=/;f-bD0CA7H.4(bE<g@>e-8bW=^<
JOJ>IeY:__AVW]B#&IQ+&P97QS=GWEcN[6&A(A@;;+Y19b=S+W9+Xf)JT?;,Q).c
\#KYd#Y8INQb>BMN[F&Qg2aaYA67SQ@##R_JeXR8HM^HK/4<;FcWb8J;-?.N3/:S
Y=DM3)@Kc3:+JV8[K>S=AQH\C4a;75P[7Pe4_QL=1\a2B,8E#&>?\H647/\PLg0K
PCb;^45CBe1>B1L,bKbE\IIe.<7(Fa+4A#KT_0Af(?7G(83?S4RE#@6E8LG5Kgd^
-K-D\SYZK4>a?(f=/J,R^A_.Tgb&7baW0AEDG5W+H=/RVLQ1gaZUSCf5?6\dbA,O
6gV(0dR\^WJbL?f2KfaHNIS^a?LOSg(](MUU-5FZ+YI>_)WW:LP\fUNO[RCW@bNX
80Ec>=b;c/:@X9X95R05eA?/]bMaAGA2,3T_R4a:4<PM35(L-:_e)KE+B5.@TPQ3
3@#+@a]V>ZaQX3DL\/^E;SYZ]S)KaFWW]\&e2+:)Yc(2C:VM[S;\Z\/-T=GQ4@8E
Z9+BGeX/@3f_fJ(f@YG[=K9f[@-<g127&\S]PNP&111J3R/X?Z]5_>_NQ4Z[]>:Y
[YUS99f]HLcB9cM(_f@Q>a8_eDX<N^D.a,cI\Ab]Z;]e#)W;./g\//DcB5#8VM4B
aIMD1T&fAa0]&baQJ@:;O2]5-#D6.b@K_]O=gW.HV7A(]=LfM:.55JB_DgXTMf<d
7>gY@.-U/ZKe.f6-]c5QK?XFTeV9AdCM6]F\OJ,[U3L2-H<;VS#H]_;1[UPS1WEg
f=7^FV]^cMK@_\ed-fQMG;69<6@Xb&VC1A.IHT0KVHbNe\2618Y\RbISY5>7K4fH
VPKY?;>7-1394Y^\M0T?).KR3?VP@+bIPUJL4X=F)\K9@TR#CbA:A?_20Fe.YfbF
.ga#5-d[.QL.Ie\(HNc<1d7g<\\b=S7b7e#8DL(RYYEP[=?6Of:T)Sc6.+6O=?-[
3X:BUKW70B>FbfaW5/=8O3_-7@gG+8];B(8?dN7INJK&QEIc3WJ7VaJIe:Y<g13X
F)KTB^<gQX\\JU)_3<CY<E5Ia#ffcZHP8P]JG9/FQ8bTPE.ST=2,b;):(J72G2=E
5DKLTZGJN#:ea[^aW.aG<O^1RUa7Y-].Bc\H/5:f:GLD^9E,GD943OKf8)UPZ(&K
5O434D]M-X0QQ7TIb1N@WL5KX.MOOJ)d#=a[25KP&&_L1JV9OM6H;c.EKFI7CegN
>R>,;KZGRT8IK-IZH<#GYI;69)UR;2-[8YY284>5A[?Kc[\f(PWR?=fY39#AD@7G
0Z^adT-2CTS:N8;>J/9@DYeT/1Sfc#edJ[aPH/4AA0[Lf.C\,26@>-:Vc-@S5,/#
WTWH[SGa9/U(F-.JG8I;9+P1M:##0R;)YIQ[L]&?0g/)-E[U;ce5A,B>J@\^Ja@K
(9,M,D96HLaB+N0P?EDJLIZa]9OO\N4>-dabL;TO1U1O&fPT0,=W)W5TF<&X102M
\8S[FB-27ACe61G17+A1>gaSM]c11)SfIL1S)<#VSDT@gfM)2/DGSdRP39QDdCb&
Be#H]9#O^@BX)gdV14+P>LJ3>4FDF_f;NLcQ2W?[[b:0UHLUN;XJSL9XNGY?WRdg
Wa3PYJ88C31DDNVB5Z2:5F2#W9I;/@Z&E:,YIBe,\G)FbO6e_HVaa:8Ug3^MBZS1
AY9_KSXYDcS?D).]+Y#Qa#bCY,9WZ\?/RJF<3aH^F:dQWO?,b6RY^FSBeIVS>67=
(M(JLPJQN3<VTD--LEdP()&[U-7D]5]V6>93THVbVb8,>B/0Z;1<Ic<,(^E^+G1Y
CWGVH39X8NCT8WMTO^.^_HCYZRS&GY>>\>;+I/T=Q>,T7NZYMJVG\-ZCZc.Ig@^<
fF6B5D#N&dVVH^df/9G)e50ea@b;&^1@Fd#4VJ0]T;UGc)88C]W<\#9Pa:QO.=41
[E3Na6[(fag130Q#6f5_+54>/0Z>PQd;[KG/e[L.RCg-<1KT7/3HG5F;FdD]IMZ5
T#LPJ0g4?N,T0,JX+>AP6?,+<2/1)Zc;C@H=bg./L:]@dMbSMW[^#2bM\[OX><GJ
=bQd\TV0=8IRGZ6[U^D_M/eOHCZ-ZIOBOa^Ye55/7QKUI(>]7SGXWg:>50HG3QSe
;_e;.@=W]e]BKd3U\C-DfdOb&+8RPffaK5H[JDD/V7Qd(c6c.3g#84[];FPT#Df4
c\&6&,,NcU45A]3D_0?/74#:D_#gC>1O+5T5bL01bMgAZZD2eOGe[Z=]P]8>^7/N
LLW)S06[K@QTfLK_&a\a89<6:XUe32H.T:Y4M^^YDRJc(g8efJCBgaI&7NA]c35>
DJf.-f#AFE):F1(fb;J+f1(IAPag6cE;.O+PAB4MUfX#DQHY;bDQe#GfQ8S@e.T(
GFEQ8>0U_(V<f[[9VF7SF6f0NfOJZ#CcQLJE1EI-_FHK//Gf?A6^\+MHaI[bK]Zb
HA7a]eLY)]GQH&G)FK?FI2ZW5LX;9_IOH(WDP_Z,\-MAWC;=g_:df?H9&]M1f99<
60U2-K?X?IaAS9SWR^XLC.O14H[J2abQ6E2aCRBI3(,MMTA8486@F0?W;(Zf?;&D
\>BSS.()A+3D\+J824gL+W]I1/c.V&cDNA\=Z=Q?^8XDT:XH[CANgW:@]46A>U#a
Yg9\@CGd#B)W6RUK:Lc@0)Y6Ld_U4EMT-c6fYPIf\,HM00bIbS/BE=?Wfa&<>a?d
b:)[.9AG(Q<X_6:Tg]4J+:G3T>?69-GLbOeY8SEBGIY3NJG(-)FC^=<0DeG3DB;U
SYR1Rb?6-DNHY\;(g\^T:IaB8R1<4/=Jg?V^>?2S)X5g7M\bOVNg9\YbTZ#f_1Q<
\SDeWL>6,;8K#VAb]EG)<D/eDV@3g\-O4P8E;b(X=DP[B/?Y<c;f(VBRN78DE8AS
fb?O(<M[M#)FM.P#&BP_3)#TgNfXa0=dI?Z\1WWSe^[JWWGcW3@EH>P:FGfe]Y)#
#53HK595O,0IF?>TT\V]Rb6F7@\0U-Of],<>:D:J>PfO<F?Ja9;JA6:gV+5P)):f
[O:XdeRX;3^0H]Z1d]&a4aBTAG4-8OZCg]+gb=)=(OVg97/WBAT[,I>&bWM2D:K1
d8-f5H--K5aD-NM^C=Qd4b1Hb50fV8RUdgI<-X_-I_RY4AEb^G#aNY=@gf3,RLNb
0>]MRTAIV6E=5.5:;7B[@GFe0UaT[KLe2bIJY(_a]#L4^D4XW1)LSO.84+@EL#=)
:DTN[JcA(bV0O:\KX@CZMJg<6S1^\af#9^YcF56\ER1?U4\1@@[f?=?8FZ:4Igf&
87##+[=A=MEb/.S.^^a4H57?c0B\,-)QX[cX6)3A6Q@HgPX((Oe58=<C#E#>BTZ4
0?VX[e&/Kd47^(>>9;I2LA</@@3SVAbHI1C;AD0<=D039P2CH,O_/29,^K)7d7V.
#ZTX@JbPgf5EDKM(WURc)/&1/ceYg4[EfHEB(S/@HK]/-ga)87,796B4CGO;V36?
/cN1_J#U^[Cc)=]0[]6+0Z23VXYXF\&2GC--CR,9NQ.d5CcF#X514T_<X2;bM1(\
USQ;GgQ7]RK1ZOM;@UDSY7A?AYA;BE^@:+Y8^,_&TL4/<(3[Z<TXVb.U)A^a-Za^
4O_^.7dB-^3dXK&Y)b3HP9L.K6A>I9?^eXP@]5))Q&7@2/cbTZ2068XH.P[ERF=0
H-VED[.K;+#JM#ZX&R\(d^6IBSZHV##[+;5\T)-gE#O1C7G)_S(b<9I7HHcH+F,4
ZE0^20&)LJ?f>P?)f^4@-+&7P\PeXI-5WFAdVE715ASg4?;N:ee@CE&Ff]2N:@>)
CNK#RY/MDZHDG.21/YH>B?32(Ig^A5fGIfAeAL.+OUC:W-AF#IDX9c<VL>EE_d2L
=.AaZ;,TXc>cI6HSNCNTDBB.=MTS)(62JI#CS-;0EAW]:,FZdSgNL=a#Q2?Z1<S@
X>L8UI?]VN=3Ec99,.(#20P2L=>cB>F[.bL=9U&6:GOe&UG&9.g(G;c_Z2>Oc<.;
ZGaIRQ&<L)e.;=F-a6R[.U@]CR&+/))//TSL<82OOT:.dYVT^=5T,LO^fREV>J_^
S?XTQ4H;Me\2QCT=/Uf&YM:12C@R0E#]>Z(aM/C^..<VR?#+5?D5+XF;J7150@#7
efICdO4+eJ7J3?SKF9:W0SG&-#\]VKa:.I4,I,TMZCSa,>9-2V#b:V[4HOaW=BdE
RGBJQ;#]9Fa3@ae?2+@P8^4/8dcA_7,11;9Q22?ea2d7//7(/^a)FGJO.^da:[eC
X)gMSAcJOR/;>XS?]L89bP)L:(:[d&:PMaW/LE0UedI^KcXNZ8.YKB^_@JU<g91_
NcK9WI@>#TgVg:G8N2X7+;&^8<\1Y2=LZX_VB[O;[#1IR,WCbF>)d^FaFB\]L9ZM
S71<=aaQ.5YAgOC+1S,DV>0Q4+\bgES:cVWUf:<=ZSFA@,ZXW/;ZMF#Q-bFMedKG
522gT9MT<J06LC2C&V+;,GMDWHG4SHCYNG][81/,Z-e7g21dB0MBL91a#WZ#Ha+G
SbFR.:K)Z]Ig2^]IcDX]QU^X5Bc5_<J]?)56D1cc?f7.DOTe@V#WX>2ZG(V0NW[6
+?Y2cG)(0ESaO3,>KW4W+9C:ad2PgEbT9(fJ&d;L9R#G+]RWFWERDI.Ub\<YcM).
8YCE;6WP3&2;BO2(O.:9SVg-7<=.GZ1>)\?.BM<dKH(Ua\?H3BP4S)7CKIRDQ@QM
\2XE1,Q_LJ,BCXaSVM6;4MC([QU>e010A.&A@g,_\TMP2FfGG@88;(aH&(LI=.W#
XD710XNcVQOROO9(-Ce(-#R)FQQT0NL,=[@9?HHV<V<<(18]CEg-CA,@?Vf2Ld3=
3bDYf&]UIOH>Y(fP243SV^Cc7g)&a34P-=&PcPe-/9[FAgdbJYQ-_?/Sb(IUT:gK
90PFUb,g6&eI=9HcZS^cFSS3G]VPa8a.G_V#,d>0c#P4HMACRUa9TNUH9D.R_BIC
(+\(PWfV=N4MKZ#dT;0,MFXEcI2:AUY,EcP]0X/Y)Ea3FUMeE1Zaa?8I>)I<[(RM
Q7_8dfA^^UZ^@^\+@9G+V1RI55b;>YZ_Uf_G5?E-P=)-@R>SYI)?YU1^^U<C?&?-
6/MJ\:/H,NZ8b=3NX/V4+WcHK>/Q)]^T7ZXUNNgIJ>H/W:bCTJGEWP2SW/d/K;Le
F5Bfb0JdNT0T4(^Pe]aC_#^#WL;SA/=5GWZ.IGY#?d04fF8?#2/eEAPdNWNH3JL@
-EW6,?](+[eH&aW9=]W]fKG0HZFQ53.bA::b>19=4]I);>&g9-LUcX@_(QXN@?<:
L25@8<DbV2-\a#:#,(.3ANWV1/;<(E__1dM,,]226:^a3MM7BI>-JLMDF[T?DIgb
fH7>PPM=e9_>cS-;c10G9@Q6f>\7=7;5[:&4A#7De=#B#PK(LOBgW)+9@Dc0[0##
V+dS^++a1.<+Y.c?#ab>HUgVD.dMKF;LIK([X&92JE0M5URBTBAg0T3N3=b<>2X[
RD3,553M\ULP-X4DP92O@P0\G_;FGF&6M&&EEB/C;29J?bI_\\]g<LM,WDQ0<BXS
N9XOb8@+U<7dKde@2UU-+dGfdDB/)^#9eg:AbP/QeEJbCN.dQD6faeN]8I<_#,Yf
)XK^.7NXI<4)^BS(-T.89c\KFMQc/8M^&XCfZ\+&TGe.J=QS&..;O1[f.7-DHBJ[
gZ6VM;JOaR=e\F]NX+JHgA<.0XSXTOQc=OE++1e9_BLZ29Y[Y@J:R?^fd-_VDVPE
]edGcg)W[392HZO#_)I12WBBZUFKU=5#8#+YB<R,;b[LU<-b:,XFQEXOS,(X-A[?
.AR&[Ff(?&VSG6X4]^HVW3VaBR,()>e)C-DL1DHE?^+98OKb_2)UV)^+bFP4?^dW
NRKKdaBFUO<ZX[9<08g/8e\:I&@<CC(]YW<bTG&AFS&/IWL^XI)K:\03;^<4/2cD
NK8L<=]ZN<BAD-F9[5>3.dcf;:FXWeLGcI&#Ea[-LdG3HRK]63:ga/AeLg),M/cN
_,:3^EK8./?19(&-9=Q-BIe\M]7Mg>@5F^f_Tc=ag_D?HL2TR#BKMbO-c]:#[f>[
DXK&_E6TSQYLFT_)ZBF,e-Ia;LLMW<<^Fga6[-K96>Ee;S4@9?&?bLCdFV_cF)2.
KbQ+,Ea\,/^+4f?0B;M.KgH0,W0Fa-+?IO+<c<L9SR#^-UP,=8d<>LNa+F[B^O58
W&GH7U)_0d_-?@TQIFd#90G/Be=)^4.;FY0BW4Bf?9ZZ:2Cd/[bg5+2<U#GA9aV0
,/NZ^9B;ZP#[bA&dX3cD\KSf5(:S7#gd/)Kf3OdU9\SWA>gJ8,-(?;#Aa(LE+E]^
RP?6:ad]ICbB)WJ:8LXU)bCR4.&B9.^F@WAWFJF3[R6]8\<Z_D;AX(2C4>M8K4K/
LP+P[=3Nd?CJSM9P[5RMSTG2?5F<O^N-H1=b<9R4D.^@@4=#Ib4ORE+4aL2JR848
Y);9IPc,8JQJFfd2f>fYc50,NQWfXKC04/39<>L<6IIaM9))C.K.I\6?TP9L1J3Z
S#>e6[e^02PX@PN.L8S-#^[WK<D8/(6TWR3WcHN+N<JBIK=a#3g#>EIWY#ZCWcHL
9/\VUL<MP#+L?&cbMA6W6=8K:4A8<W:LRAK9<B,H/R&I;GN/U;A4gI>VRcPQ><+4
.3\#XR&+ADKV[C^@@CV>/5L6:d\cON-QR.A/gU#+c3HLQ,d^I6Y82O@SC\O]gJK#
>D]AO.,<YTFfgX<,BI1<b#+BYd),QM_6B:0V[.N\(VVV^Q12]<O3ed_ZKDaI4(J9
eO1_>HXLY^(ZH&:<BMd1BeWYf#P/J>+OWDF\?JUDJaf.8\=>-NC\-I.G>EJ3HJ5?
4e:T6ZJR-9O^D-,TXB[1ZQKfFC69#0FFeH[-WU3OOUB.SVFedT_#->3d(DOJ7@:0
\#0O&JMR0ZeWPQN]^#C^^KF&(^GDWY(\gVeZOS>?3.Pc.[J>c88S5B\M1IS=(HW2
@:?#5-([F@_#.<0U/NV[@]d<C(f)XCb;Xg/.a(CT,=0YSS1bCVY_J7bG,@QZ-T0e
N@ZDf689/T4ZRS#7:9CRM#6ILc:H_e@BXg<.(/8]4)gE^d/,:59X9&8FI.MM1,^H
aIc<8^=H.2?.&0[FGYX8/#W4VLASHVfA7NS8VNV@B.3Vag3dBI1eg=f5QbcIgW:S
/HF>EO3YT;Mge]gML-U4/^+A,Z9+0Oe6gc5S8&,/+Z.=;BD-I6[g?ZD&6-]a0^45
DR/=8B6-.OE,b42]E/UTNN,dbVTYQ<f31_K=LX;?#-f0gZ,#SB1X0?JJ:\:@;OM\
,.&GF>g]ZY4A\S>f;+]^01FL0:@Xbc3VA0_JUUKHN@98T1c5Ia&-R?539BaY?_^\
([7QC46ed)FN1@OPWUCTgS6[\^N&A^4CXWC&-&3@=^B(AcB:<&b#bMfcNeZ<[f-P
L7&-3K_QCXK4F8FYDTdF#F-d1<A_[B6<_AKPLKIFCL:1)4=QEg6Of2NaABFI8&C3
U/EPH31W4.b[gf0R?@F6\?:882_+-,)07.OHE55Y=;(/cBZCI8Z[GT0LC>R?e9(V
3LdB;L&F2@_;=6Q3G6(RVWL4NcU=DE^>+P?A7,d4ebJO4S<_<1ERcZR95cZ\O[XW
YXX#a+([<F2+a[E[M>G2LCS+/5N2@FHI\G6M(>S_88>#>eWc#;G^ZD:#Lg=+NF5R
d189.@a1;QQ6cfRgbU8Q:_9S4^JRA,X8cg4ccf/Fe[QR,I/aPeV8+4O-<23Fa]Ie
17.NI#MT,M/LKJ_4KEN^ff,Y<,:2g:RSR^NS_3VTC.M4L+F9K9>W;;]b=+934M8T
9+,J+]OCKF.fgU_#a[6U2Hf02S.L\3P[WBX&A1GW^-ece4Y7.=H8IbRP;L3T8O\>
2SS=4[=R(aR_&#6@N=f0cP),K#T#E:d;;4TZS8:M^=S1RLR_U<1-N\S.TPPA87Qc
KC#MeM[[L/J6IG^5<M(6QeRP179YRIH/_9U2R0U[BcW9?C<(@FZ6R]a3S@:/R#bI
JL/[.GDJ;<9^_b)e7^/5N1O&@SJ\JYaa8;(?b0:_+^P9UCVEF<).4QZ]/S^:>F<c
aU##SK\NDWFP#5?GK8G:+3^&R(Z49gF6-@EP[7/AQ+.V\#Q+_EV=PO_a_ae#d#UR
ZK_EF^8<_^/^D-0SXbOTF1>K9T8c^RR5g)2C1J31?&E<aX1(Def0U,beARBQTL20
9@JJ.be:&V9.Q::=QMD>f[Bb\N;M^?6;CgFMdW2UBF[I5IYcA1eb#@e)MYTWca03
Q?/=:OEb?QXd(Na+Le3e2g:FX_IBKSa:DO@AR=Hf<+d?3AI?\W[?-Sd]&EE&0CRU
H)4.3-H@6#:=L[b_S62GReXdVCZN+7C0J8)QfNJL^#262f&\]T2#@\01=@F=KBf1
b7g^A9;-IeVF#1b9C>=3@b,)0_YA7<VH,ZVBeR#)KaH)Z0N5J4QW#6-=4TcQ<UK>
&IJ\SCNH0;7=5gQ[)L9B?N_cN_fQYBd0.71J;8U[+Z8.4CRJY;[,TCT&-FTcNCNT
7H_,3I@5&V-^JU&CLO;T?45-O[NU.)5d=aDfH=^Q:G?MT\\JMf/Se_EAbI<47HAC
34XX?_+<G@)T1YYYQE^G1cC<;9&9&5dd,14f4]RR@,LSJ+].8G)T)>X^1N:XS8U+
]A(OCQ20>[H/;I]]FK#Pd0B0-OFJbe0)cGWdICI[/[V]6?<V)P8f9b?=<?KKf1f_
J_@[M,@8]KV]7L-&RM=Bf1S5c(]>V(WgFK4cEEg]f6P-dMJKcd0J:+6d@a<LF&8\
=F]7#V^K5Ld#-8c(LeQdBJ]8YK[g6e<_.9b7V(.[AFf(BBIUIgUI@ET.[P,441R-
a)cf10W+46ZZ[:P[/cH_:UD^+0ea@&3(FG[+B7#Z(dbT/U,cEW\ND0[f7-R-1TWT
)TP-f#UMa+<VA67UVM/V&V_Kd0XYHZdL1XVAagP&HYLf@9E_9P>UH+&WHBaRZe@B
O32_3f@VM3WSE3FS>H@2TLBL?J0c1dH._[A)DW#G^dd=\42.[^Qa7V)3<_LI3T26
;#&1(Y./gL\<7@,/-WaOb1GE;Y1C9cfV],Y;QKG/g-\LG?SR1_Vd^WOTP4G/IAUd
DFb7(O3D5^F?NF>Ne(-eC;eSL9UEX9_VDW\8N0B._8OZCNa_[8DQT)5&@)=>RBSe
gBW?]I&a&eg>R(Q(3R\=ACF[YIbA>gB^K^VfGg.gI.NHXALDgP7=>9YG4BWYA^?K
]0W_NQ>4RO@@<A#(VG=GQ]3\MZP<a&&[7+b\GQaAG,Ea;PA9_][A]1D1X1/GT4K>
I\AgYTGS1KDG]>A1UegDE3(=?TVfW(3aU\8G._UAe&FL3;RD),DY1O>B@dO9BUa^
Vc7Y>1aHL(bH89<23]<f\0T^(D;ERQOMIX]4BA)2JeTYP^)Ha>)HUKBV_c-/&:B=
P:Oc/bRg;1&4O#;,F6;#b525M^)PATT@gd>Cb2(A0Y00IR>9X214TYJRGeP#Ig7K
;SWLU1Q@U/W?&SN00U]eB0g#;0\L7C-cS>4I-FX<&^<VC1\8d0,@GSL.#8N/9#3V
PNB78XN]TXUg]2&P\)E/6N6C]57g,gHf#^CBVT6Z/]c0/&TF_(JQ&>5::.?Fa,aJ
9UAKI;g]IW(5O7bXZA<dFIceaEfD7V9<8EGYUM+F+C47+L-DU+\?NBgVSg,gLg8W
[;M1R\2_GA71^Mf/,_&G:H(\FO,4<b5<54VUR&JD62c<E4Y30G=K_93#<a:]OF3?
f;?+^UDIgb3A9MW7c6TP]dF/OD>cM0S?1_RO+@1^dF/e^]fJbge2g1\/DRH=g5Q-
.3L.2@cfT1TYQK(a&^&5JeT&/McIRH,:(>V&Jc,2M=M84C+R+Y<?d7F1.17OAX,4
(,BM0F#YA2Xa^g^KVCSNK5R+7)\\M5@4DRY0f0Q/2I,#@BX7_60g#55&\/W0[+,[
(H&aS+SF2CLD1)P-8._SaL0Z#ffN:;B@<gC5.GOOT3a4g9_^?MR=;8R2#AH.<^JJ
2NWJ_eLBNU?,]X[JU.KX6/)T7A+R/ZX/&=(S2S4J#W3C8Cg/AIFTBH]XC>E3V.bB
T.OcS??ePQ@;16<cUD\g;/(g)>S/X5cagPU=1_XS><B)IC/733V0)]E0^9Z,abZ;
UffUF_36Sa5c70]QY6a/RFNG6XcB+WHM=0F2BY^(<F47,e^f_LeU^N/6dAD5R9R.
7,C#5(B3@PafZ-Ig3J/ZVHCXIcSXG9fcCNe9,80NUGGB0P]6A5^^ECRG?L+(VOH,
\bK/G);_JgbI\P)QfSXTJ-_bNb<ME#e^.6TE5UP)W.-<0>Xc)g8>=_F751/\dc<@
\Sa>F&3b=cf=_>R^Zg7e&]Db(+0(.7^OPQTI(Z+6dV(Z_\]1D23=<IQP)OQA).+[
5CYa>AX]^/=SH#)HZ^DQ8DKTWF#+N.RG3)U>#HC+1<dZ2f,ZBI1)CC>Jc(H4OAXS
EYeR[=dTC2Lf=[E)^bSVRAYY0Q[8U2(.6-=KCY;\B#=J\SC#R3XO-)V/Z+Eb]2V0
8+e.0#_Sb?d#@0/(+VWF@&Y?FQRDI:C)3=@AQfBaX3-?YQ.6.\/MV7e=\)R+PA::
>bS595)?0M=-^7=-f:7f]4Z;Gg47Qa=VLeSS00fBT0Rg.(TY\E-1fa/_>cFe:.Q8
5eYI/@(@a9cV6UF[;Q0WZ[d8TU=c8N-NHOb&g&#-O>D^fDb+P-OFXX7.KC8Cg,)^
W1.;I6,,7D\FRHL;H0N(85HAfS1K+V8M7AI_2Vd9>50(CKC&?5OB/B4c+d[94X#N
eBPcA,g-CZ)8P<&0#\[^W9e6-U^b+/;W<a+Z@OH,PH3aQK9c2TFJ58SK])&FCCVa
I1+B2f^.K[>0@I6JD)Q-5U]3XLKW\-.Ha6P:8I/2@GbZR.X_RMAMGF>L?/B7M&>[
C+4==Gb?5&Rb_7S&4AccCP?d3Q6FBHW-Q\FaYI-37C(F]X_McN<(gDf;_QH1LBMT
>\N63J8WVK@T-VT#a4B+W(2.g30fbOGgfW&)&A-b-g]@+5-10M,E805Q_1Cc:5gg
CQ&4N:&8#I3b;EUIU1NfgKdX@@8eb1P^b0;b3;(cQ6/7g^6bW?T+L=D7=1Q#YMU_
56(XE./c#caIH;N]f,C7#8+3bH=Z6XLBKFI3()#:^dU7;Z.5G\#g,T^J_A?)@Y&Y
]S;VeC]<?(OI9aeZ2Fac82+;1>O;Ra:00HU<N>61Q>JRFb-IW7-#NL<.KeN_+_W6
O/4P#010YJa]#0.X[V)K+;+)N,-TN+ENS#59b-b/2D[241E1)T/7aa)?c_b,K8]>
Ied6e/,#<:PQRVfI_#DcV2Z5>:90^;6D:_G&dX)+aQ:BH2(PgFZe)5c>DgL(B7a(
G+:<@XCZ5\bQ2.?<U5+5Vd:OK/V#A7cPQ;IAUL7)f7=PcFSY\75V<I25?P=)YYT:
bW[VK1=P=bPCL>cUUFXO8=H&#NVgK;EZ/g;BS/LI(A&F_9,0I83RMO@C,4;A_eW,
)AZR5Y.Q4K6UY(1GGeW)4/5B1K>:O^DM;QM7f+\,1>6V/U^d72H9@eZTE3T]WYL)
dA0/2gT?KZT.KbLFP[Jd[D?6[(8LCEEdW;8#^&7\fALQ#J7a,/.=/5B17]G6a,4/
I4SSQ8^_f,K1G3CL=.QH([,?>,;K]V(QN3+ScIaC^H2[&=WN=:W^fd2\9CI=d18@
UC&WZRe1?#Re];5e+Q)K0#0#<7K+9<.[QE3R>=ac5YT=BZV;g-4)#BXSQFUMNH^(
FP93(-c.:-=<[(QN30QC6UFbHKV4)Y_:000P+LH@##25^+W,HgYN[X+6()0)F?XB
_WDF3;8C52,VgC0P2Y21X1@Q]PSB:IL[X=N.CEdEB]3M:Z4c5:LQ;&QQ^_LIge6I
LH2=_)YY@;#?8V6]f-/)cU>UF?0A<M2;D#<L):H&]3,W6#(6HN[6.KPL;IA47#3X
D<_T0YGMB5&X76+J:=IK6]&U:?O]NNee&?3,AJa-b\]JdW1H2cY9F=Rd2^.ee+Xf
g2De[acDK@372B2KM?eN[P8:S+RAa2C5a&;bd)T5;:XB)188S^C<T(Eg05#\P3SZ
.+[8TVIBZ8)@ZH^#8DK29>#SY9YSA>]SU6VB:P9PJ]8LeHVecB2HeA1LU2cY;6G]
Q2dW8+WW#CEJV2c9ODcd1PC)<<C,aG#^;B5-M[+W;]+L[STO[gHO9N<TZTG]7.IO
IP)d]Z(:39HDLT1.2PHC.>L#,af.X6&f_F&+/f2E(J,/A<)6KC#gGBY>.^5H:DfU
J^4?/?,adQYDBLGDaS7]+;2bc=5#8DTA;,Te_:9_6Wce=a+8)55C5@Y6b7b/8&Z,
cGK]MDD1KCNFPe<.;.DE4RSIVL&,HaF7GQ\=H(;^(UB:DDMC(HIcfeaGWQc&KBNS
3;U6MH9.[TZ+:aG-92+4EX/L2HEEBE&1Kc.6g7#<IU8OCKTA)GOYWKIDe].daFS1
;IYU:Oe@:-(U14(#]=4-K[ccSUf>XO)1[ZR5K\.3;#WLJS]]?0,:3>O59]fC3.9b
@)OdT,CR@Q8bY6Q0J0Rc[(_CO#c.dPD;LC.VI+L=<X83&KCgdKa_YLC_CXQ:eCB\
/3Ddb7@7RbAXXX@,GSagZ/_dGA6R?C9L2J.Oa&c7M0\B76]MHV[/J12ZY[?RR&>5
P.g[W7B6A78XOBcD\Q7_H1#XIB&0NAZXC[PPY>.G7.d^cKI./ENI:V]GO8+\+D/4
<He.K3DbeBdZNcL47W4<4(JRLaT[c^1P>;>V7B_f-5UGZ813KTF40SJ_c6A;VaGK
H\YVBUZ,+c6XO:#4A#>?U(<0_27)@UU8eC:(9?(0Ne6-IO,ggD>Id<V/U(#TZUF3
9MLfC6(U>]R^LAZC?QA:HO@5dE^0^A8TYNf9Tc6MD3-AHD;Rf^[7EXZ,cK[aaTAI
2TFZIf3;Q^Y)b7NS.#R]\RfWeeT3L/gILZM0bFe903)@B,8X]Yg;.ZRE<L#OS6GS
PgcAPIc8Q:\N]<4L>+X<a#&XW-1GP)LXB<.-:WI0/2D[Vf,;O:W0<QF-CB3M3<N.
/^Kc^.g[G[5f?S7UOC<G,BFC,N^ER1KYB#R0:-^K(?eX?1>>[3VI-(DcXC-@<MP+
M;7/,OI+,N;EMg9U4+SOd1TR+&U<V4LU-)^YcEca>_Wc\E/1Y1(bYeZ<P@\cV2.W
9P/L/(.D.>J;2a)N<^a12@F+8M_6.@1eNY8-b31&a0GU@\6E.V:Q5/b]KfP5)-)E
JJ_6f0.Qgb3-F\,)d_@+BL/@CNRg](dA:4#=1a4O&MLd9U^@8)B)K4G1HPXA0baW
cg=b+6R;+5SKaWb=Y+9?B7-&7ZV6FEJQWAB2,>#(_5]DH@+E[Q\/.;>>R&E\/d-^
W-_L<6ZHf#A#><GaC(g2+3f2FfdLPH&#3DPBTE\.-:])7W0D/>@Q@4B)Je11FBKD
J/&L3JP\9K/d/Y:5U[9A[Z+XCb]9_[FO6^QZ.Cd.C<C.D)]2C9f_,J<W-\>EN;.^
<5;PKB+Cf>D(g^KM#-D.85,T:eFA6TdD:@4@]5=g&_N:NS>IddVJ>Q0AA=&\)-_=
EQQ,3<L_HTN@\L@#=ZH1YXcINdFTA(6M1e<.dX.PJ+#K5XZ9.4?J06KCPMd;+W\g
KTQQ,/5GXZY:/9a<#BTdg7G\C+FQDPLN9Y=b_NM44d(Q90X+N35Tf]F:W.7d?]dg
OI6UHF/bWdeeaT,3DN>>U5\f/N&B2+fHSO[d:@)3Z@\5OS9[336X/CTR8MPCN^UG
NOVO4OKIV1MXdcd0SZQ)<gDD)B.5)(L4UN)5M:W-@RaeHN7ZP?>^_TNfY],EA3c_
4#9^aH_MN2bQaM7S\]+@,F)[8BAX_]PL[[eWg2[E)+I@H<M/fG[7LJ9bT_<98&8Q
+BU[F5R@7Y9#N?[;A79(cZeAS7g>U<&f/HQZLaM[c^^&cVNR.0P_OL3Ff6T0.VT]
/&QRH[a#]H5Vd>UC>T9T\XBM:?bM_T0J^JPF0fL=A22Z->FEBe0a?LDQgJP(>5)?
,H3&^.>^gAD6^5^:-c_E?Z[F-+S^+B,g:\1V\XD:)LX6-bIJdS2.NF#aBGN6>1.e
D+_G:6aYB=CKO[&JI,,U4XZ]eK[Ia8I_,6Y=eU.DIMMCCK7g]<[^Q/R066a_#CgE
_6/B#EUH]:#Tg=_c>dMBK=@OB[[ED:BdK/e)9[LZBTRVS4AD\31O<9f#a([RBXSG
4<NRUJ=M,=6;<HW,:5fd5U,W(H1NFD[6MG^2Dg4H\:W<VQOd5>b]\DdX5&?IMPX7
dgab=1;L68UO:D;_;))(C(]=35I^e74Z,YH&/cCZ.G;Oc#dLT\:b6Xa4N-R=D&E7
=]dTM9;<LXIagGRJK?/2&#HB4[T.O&BA4><AcE#G5MO-<,Lc(:,D&>(WPI^c.GgI
;.96-55bfeQ^N/c[H^[_O2ID<5+)]=a_+&#U?UNF8O[Y6b>c+_=2RF.(Y2LUA>Y5
PTQVgVMF_73+,9=F-e_?7[g,M5<]PEZ&#?92VA<[^/5P992Gg?9I)VE>0YaT@?HG
2NG7dd-QHZg/.Z2<O3W63@J[&dU>&K@0aTE&CN1aF<H/MD=X37T+W:74E[P3_f#]
4QMV3MMSa4Y@^?=e9OI+_#fQ)LBOca<CY<R8GZ<NU0/@f^C-:O6HBdS?O(VaHY3S
e3c/Y?I=0]E]#K4RV:@N9<+ZZf?W\2Z/bL]\Dg5_J,EXZZT3:?2A#:/7>LPN>cDW
8G[_?Sa5BRc1a[K0,3a>:RORX3X8d<7CL+#G8Q+d,D(WY)9AW0#+4BQd?@<[AH=f
GE_,><\L:[;:d?9G:18:J=ZUAOM0JOa?/RSg[4=/WRGTD;dOWZ97M>0DURBPIg(>
+,4CYR<&Ug9(9^Q_ObSF-WHI;_0AbfOT^(1&#YG^_g1K1?,PAEJ/X9JUe^CS12]2
)-H\]Tg=]<KM>3f3[(bX,^W>EX<Ie@13VG2Q7<IgUeW=FFK;A#QK(Se>Ba[]P=3C
cgH(1Da6C?>=>4R]<P48W\(YL7YR8bK=2J_X/)MT-gS4V^B.4eL6I&WGYc=WI6Ug
K8K^W6-QRacY3gPJDC]ZdJPTW67)3(FW:[S#,6c)YPD.PbTeB=]C?@)]((K]OLQ3
K3C2F4\ag;];3Fe@RL:b;Y5b5R-Y=FYP>##&cX+2Id9e<a.F;@YbC8:9,9TU2WI(
&WefeGFSTdHBgWK5_C]X/R][2=SD#0[]QD&a1XA77]\WTD8Sc&Bd0]OWZ.3NLL.3
0+EQFX=O^Gd)BRKM?^VSB@6PUEG?GZ]=-PR\14@UNZ57Ve#?K80G/8ZKYR1F^b78
1<8GVdKF/GP+2@]Ib--_&)5+\2bWaUYPKEbK\X#V;:[0W>B-E;:^U=Y8.0eg:?Vc
NULWgSW3@T^gA)=&,2S<FJF->E+g165IWLQO5C[/</O0KEA&(53T3=-5SRBbI:5@
,-H8aIHI9)DMH=7(]J)?>DG8[\I<C6Z#X?#\6-bW.&>GVWSK/#F4a\>9<0AYdM=c
(cM,B=CB39=c003M2DKO:X8>4FbNCcd0V:IWEB:d+c]-A9<\Z&XcN474FSRNRgca
;DOdW82P8aIV@V<N5^bMDWDfX.g;&8>(cOMf.7JD1G0XU-)\/[Y&eIU@(6Gc6ONA
c/]Kg8)@NX=^gZ\<e<eSaOdeZSW)H2:/K6M]d(.U.,.F>FXN);0-e.3FW/deCIDT
3dcfG01:W]&<H&ID6IW^I.J.GY;?eP;E#5MR6=DCHV#]\>ODBOY03G.AI0_DYF0)
[-I.87:@,Oe9YIB(KNM?bG9)-NC=01cNG_b?CFdPDWfK/(#CQ2IQaMcE4YT2e2]8
#V)D9\cM+c(X08LYgOgEU3bW,?<6\@48S/3^786N-1a2<HLDaZUUeb?.GV<QGGTf
M#UX4)(HDWT8GIIgC:BG:#K+CP)d[/JDfKB_==g7G)(8]DL/CUU6K=;ZIbK8+NX=
<NH&(/QUZ4-Zb>X:59=(_+CP)D<EWfZg.3WO@a>E<>6SZQMK;cR-IH-a\0=G>4&6
?Z;K(#H7Lf67f(X[#29PLF[>2NL&QW;[cCFIG[BLcJ.@<PV:dE;ILg8.?YX;_ZEL
Q:0N;)aF_9c)ZVeB\;^I(-4./XFTY/.975]&A9]KN\_bbT403BK]XI)[V=3CKaOJ
/-BN?,AHN:=Y.1f^;M@.EgLM8AGJ^\GWCFSURMEgWVbPQ?ceae?K64e<FL[:<T-T
.B2fOS\B=;UXT4Nc/9d>?0fN<0>Z6W>eQPK2R9cJH7CC_-6JM<DJ)C3X]8BXd3F,
YJTVT=Z=\5bSCY(]:2HN].R3\1U8=9(?.+FQ[@8X1SCN,@-P+Lf1:PL>0UeJNLf+
6=-S/Q6N#JfD+C070CCV6#Ef1-4>O=P)6P:?\A>V/P[YFRJPf5/Q;]E=JU_7CfS#
1DdPW\:A?,,:>)HY[^==0DWU<cXR#gYKec2[];;X.WG)We:SP3HHH<?P5D4),T1c
P3gZ6<eABe9+EFJV7?2C6N+I_V^QYA0MKGK[8Ucc>=EH/H\J>b)+:XU9_\4OGSYb
7?B4aN\R\;>3\RIc9_&^\#37e-WMb+=QUf[ZH.)?/MD?b8OgP@V(FQ9PCM@T.a+1
;-(b]-;@=_YPcCCKC+GZgbECd7YRV_0CMOMY+OW?e,[VKZ\f47AQcA43f(D&#LXV
B+f4[/^^[I.f4^Qa/RXM\0FWSa__7QLA^#-,FP7Q=-;#A;&5LL))8G6daF>>8Mf8
P9GFZ:AFFaNEH&Ta)85/W3_BAC7FKTJBCU,UFTO2[^\\EBS2NAc)f].??/3D=b>+
;1CQ=[e:b@>]2;3=J9KD70_].)4<KK211Q@8-_N>_&>Y:[K:(=&AfI_P3P0VY/1I
Lg0=PG3?8@W27gJ-d>d?R=5+10dB7.>N#-1/G[9Z4QYJfOZSAK</6aZZE_8FJ)6A
7JNP_g6WVIbKT+Ha/4,T]2ZPAUR=3Sg37##C#d\24N/5AUdMf@Q>RVAT?Ge=ad[=
.OIM/L-^.Pg.e_VaZ#K0>,;+K8OaB&S<\b@aDV.C92@8D,8:#VLG._(4E_EXEcLF
T5X>2aP<DV-2/ADQOcb+g5.?^]#@TZVQ_BO#PUY;e/S+eEc\,b[J<&N)<4Y,^2XX
9X@7J\I8EgfKS:]:@I1AL#/4SS5-ZX)KVN[2?gb6PFg-LJ8H4D@(,+Y:PSd#:,eF
e_H+=L0CVBcbNX4HTF>5PU9Z2a3>VUA-(10#[cfd/[GGdS7=SVC:,;\dBR4<feRJ
9>9E[:9@D)Cg3eC\<@09^V#RaH]Q6@f+/SYWP)^/Q#d(/a(U5],:WTc:;KP6+5=.
@PfDO[da>2gYG/f[\@OKIV->,=0ZV+X@@ZRRF>?]W/FNgMf&Y;3Kc):N;@=b\[L[
X6Og4HD/^Zc_a<.,F(L^SVc;fga;>)_U97N@_Cg^ZOYU2b;PU,fR,KIM02)/J>SH
QD5Lb-TK5bMS&>2<O[2[/U+Y\]FXX481L[WS7c#XGP?e1.R@\gY>FQF5Bb+@DX3;
+f4P8PdPgd6<f8O<[S@Ne[+2FUK27H<C969D^E@U?<[V^#LJ1=HI9O+e0CVVHUSU
>)aY-JP73I1=8.MdGEIU4gCTRc.[VP5?8[WFN+fC[;P[Z+>;]SNUJ1&;;G>+WfWC
&cA\G1\Bd6>PWB_@0VBR.7]7OYQ<APf:_.S7OC6S[K/U[2D6@90<IX3^F=1D-J;S
,@D>F)YI6T2?PKa.TN(.<>:9TR^>&S3I^K0e.TE&=GP2DbV.0K.JaARI._2bS_+N
d-T8[8G;&N#?W<@T;3\4OK/MOJ2QN@e0LCQ0.II;f[c1d62FE+S09g+gN9Q-]1CV
X[B/1>B2Z-?NW+_aaOL@JNE.ebT6>UZAN4[_NaPM.e><Z5+[IRK8D;_;^d;/ZSXH
8_63P(F^IFKU&&X01)6K-Y[G@Qf-H]B86NRC>PJ^PYf_5@fbG&[#D&Bag1Be??A2
IN-X0FVTFZI[DM0]=4V5>/KXO4_MWK)0=c&)0PUf56)076[^#3A@&.B4b_B&4]]6
H@/[KVe]T+_1&S+[Ad7,E^?8M+]64gX0L+/F<UK-XEc\dC#X+f_c&eb<a>X+9;3e
aO^]MB=4YaPQP,[.7R>5=Mc?#BTeN>#bB274Le7[e1;^8;?-HT-=Df688@^^(SYC
)<:3De-bX#4C#Q6OT\[A<?W?Y0L[B@B\G#&b0E]97Y>B;[;T8BT9&3:P1.Pf&B_&
E>gG[b-gJdD?E_+(aB7[.NQ.]595?QNF;(P1QSY;:3T<Q8J@4^Ne-9YS1P)?7?6V
P]3M+JEY,&F0Y&WaIafMG5Od.1LSXX@:.QI&f;:3SQ^@^Q6c=g6DC>3=/N7B=(9I
3bD7CI=N]f.(g7\K@Q2SY2..S3QPA?,O;Lg=;-_Z1P7SL#C#]N\EAFD5B07E3Mc@
D7<G-+4K\^aD;PO-AKD6&EHFJS\7Q2?A2BYX::^L(&&/O&(<&ZW-M1b>cg9G(^c#
]X0N-YW9T,RZ/.f=1<0^)Db/IJ;DcUY2G=UZ(:@c/G;[XX[eDOO)e,GO;C/&gF;c
MQcG,(+_48T;0+Y-TT3IJM?<P]4/\\+)U5=-LJbW1a88YX7WCV8G#4VaP\ATb5JH
G<)dYZQbPf)?a?Wg;dbA/UGA^Z#gOc[0FMYP.YP37WDYG12d^D>Y9.:H@(K?.Gg3
-S)YK#ScA&ITUP<7^,D&,9e]L,H/>L7eGc41(ZD;fQBSEL25>VLG74#AKd>8eDIW
(?gSf01e5@^7c:1\@6-cM\EI5K+e_8cHYU2[J=2,/18^4=BfO.4aD#9be02#7I#;
)I/?A]\/d?7b0@R/JD^\T+gg(AO]T\_@O)_PgALO?E+HR#fQ-GaWS]dT,<?F-g<=
e>[7:V\^R2^62]e;JDM<gNH-4=37P)L4cO=;L<Y4[5d>8;.E]PE^CR_O:Nb#-,Ya
6U0Va51:0L?-WE/^F^YY.154RZQ[+M,aF0GU6/ZML=0d7d29ZF&/CU2()Je<aHVP
7&P&8(,a@\?F5O7LLGZE;+_C3NVZOA^JK^08)fCQP]O&B&FbHZaf)E:f>8MN89ZB
PdI@<QI=1If>&]?=_[?C;TF7NBY1P<,/B]X],BbUbSAF_\?&&=T_W1)JA2<^51O>
ZCbN)XH&f+VD@=cS)^d,J@]4TGb?QAa;_732;3CcRUXX,d/,YaI>4O:-AAdZCKPD
FA90<S:+Q@,JX#L,KF25>B)1W,.A9?93;g5YX+9YIZaJ#:B(@R^L_#+5V7A3)=(7
\S\;;Fe.=Nf/-#+)L[5A=Rd-EgQHVW&1@F>3cKK4@1[cbbQ\cEgQ=DRRP]>QKGgQ
/VJ?Z3_;XFLE[0-EN4Z7]fbda:#J3QM_gf=0CABaXO?c=-;,]bJ/Jg5(c=:aINZc
Fa6?;?R],LGDR5?@O8d[RYVT_e_@dEII^@V8NRB3@]b4CK>[Me2Q1g?QTZC,#C6S
2Oe(a4EC656-=RA)deJX/-.^V9+D=6IeR^V=3fB.(WB,Y-6XG]4e8^:^ITXf]CB(
#2K92=OCVFG8AgX(e78G[UP)LTF7e++V1c^82S0789X:Z4(gQ=F2W8ROQ.UUE,3e
JP]+P:5K+M1WTOECS2K4b8fd5c<:<_]O/4gM>;&,@=GX.1b0WZ?7?S4(NTdf/JcY
gG)+a_SE4;5(e21+Z1.TV6&^fe1P#V7U8J@8VCW-DU(17(-PZ=NX-3=G]a.8b8\T
W.281J:S;RKb/O?Z_,B@0?FY>;B2GU(\TXQMc+b#0[Z^-@#V\=>/V#SDf]59a[[)
V984a?4AA\eF@CDP:<&c(S9E5e19,T:fWd=I?0<CbcW>E9U979H7^Na?\)-6>D-d
C&-9@#6P@=]8dV1S3VgT&?fGFM86>:5AM^bg//2CDDa3SN7Y]YIC9H__8=P(L\]7
7QaK.0F_6<_Y8CEU?/0I@AVeF.5]UA:5_<C8FC+H<)WU=dcb06;=J<AB-1He\bDP
Y:BI3/Y&@PWVU_+[ba#N0WG[1T9U4>A8_>JCN4A5Q?1+)f;?I#.3bM_Y(:47M35P
\2N7C_^d.2WA[=)=b&5W<G@FRR=XVM^-:aX++\)&Nb6?OYM^@RE5d@/_;?/R7)[9
2TA?#K5\G-(JAM^&ACJ9ERbL<+(2bKW,3T+HPJeE@=&cKV>0M/<DRGR3:GOQGOPf
(NHbV2a=Q-[d19V&<S[_?T9R2]S8VTTW4_W0NP<1NJASZJC<gA)QAI#6c@a\\(9)
ZL>3,]GC<9/ZIb7[PXREH)NfCKf.@eKW[HES+[fQ@9NV9#\3gc4S7BG?[TEa/<:J
JV(Nd2#PdW6J&b74O,0(\fAH1#NEW[[D4WG+G]a8Y/ab#f/_B#JY[1DW0dS/-Pae
UZG03,4QE]V_6F5>5;2GX#=6C=/1GO:2T@F3eUgbf@fES)L8;-G?KE-NBA<I))f6
@6LX0MaG3.VR+b1#GB=V-TA4L0b0_E1#cW(K7[Uc2^cHAFY>9PEOLO;BYf=#^)a[
_IRg>7K=BK-9Xc7d.5TCAbK5g+399fa/2.BM&?<]2>U]LYVP7g/QeB_ME3M5.NB+
BTWOeM:d9fg]NbaDUQOPAO?/NZ<CSegc>#LQD[9#+DLa;e(W3D>U@,C(5IOA998;
,),10HO1G2e45Yd9f#^f@BS<:[QbTFP?(77:6O]B<5_K^6NPY1.,(M>=fQ+=d=-N
cXHT@>0T(I[-A^2=c=:+M&g8^R_/ZH3\X9.U^K[L)QZ5[6^OFI0AIYP1KZDX5M<G
USa2G@FM.J4aAN14^]Y+a)V[<aORFg;&ADeT<RMZN+f4Fb88-9H]eHIGOG],HCN(
6B66N@5c^Ya^Na4]eH+\eR-DUTRHg:&a(fba2^Aa@&R#AgcELMe=MU1J27N\UW0?
Cd>cJJ=Y8\0P:WL)SGZFc5I&T@U\fg0-Q(^ITDS2:/GZ5/VDRMM8Ybb3#P@Qc_LW
;/GG#<]E)@R<6W7+#_9TE4_[GH#OLC(g1KW_JUHIC]0=T#Y-dC[RY&6;R(a83f(^
Pfe><a7X]]U,C(@<R\7RAF125)aM+F<HXHXTMJW4..f:,\FSHLbfS)_FSX\/G7LB
.9/_Rd4)be[60&(+OeY)aN#UP-PF;2W(5N5;59M2d5_NB<2eRP:OU@1C&bM],332
BA1Cg;V7;MA1GUaf6<TG)QRGZXG>1I?J4<bY7A_fBe9R<(d5de3IXQ;^B&?+D;AZ
X6&eI=>eSJY4P_?.TB1M3=9XI2RPEQR?#RgNG>VJJ?W;F+2>WcSYfKIed:B9^KJ<
]);a?CfZ[4AS#,&VTO0./D@bbR)eVMSD.(.-NWT=7M4(>+Y>IHJ5MXS-5#VVB6\)
+N>4J3,L(,CfO21@ETDB8fT0,AD^A3I6^)dXH>O:\2147aCg\<1f0XC6cL9g.4=M
(=@>?#\b@V-0QATEKE=:egIN(0&P8C92-Y6E@H3TX90HF\/;^:c6]JD&G8a&G1g[
>#0@._24H?D)(+bI-ZT5+@WY#HL1NcRR9@;RS1>bH[^1>[]Q,OIReCSV(Q59Y9JT
@;679/]aFHKW6+B920-M&J6ZF@(.>@LC(AQ;4I7&\-&9&)68_LUNC&gLd\/N&ESP
DGfZFC+R62(:>LC(-eaVMCe5[UZJec/:.KCe#ECR8]>=CHa\J4a]L.T816Q\SHXR
]>S:I2G0b?FJ3d6f]DA^ZXL1O@c_c=ebDJ-YCF&5FVX^W<<9<Ied50f@V_QG,FCI
L-,>?A5Ba93<+A@@S20II211c?OfaO?T1[c.^LES[N=Yge>Z7d677[.Q@&A/2(gT
\Q;1c(Z7Ha/&V^Q[d3<;LZ1]Q14C6489/KG(3T:I-<Q4)&HW#AKP#aN=;Q&-\fC^
?B]Y;V3\aIa1gd.D#Y#&LLEMBgI^^WTN(USF^_5Q4=TEg2@cX6cXg:DgH0(8I7W^
cYdACfIG1<NUc=-M(aW,T#/(&YQb2IKW,.UXMSIHYd@I(<V1)L6:>:RF>,=LKfa5
0Yb:;Jg.Q]4D::12^4eBO=de..@VLb55Sc5Q1=Z-M>e(^CM,RMMP>0gB_KeB\Z5c
Q5a5a6B<-be9#M)F<R.U[WGI21&<+H)E_4DSZ)BcK:bc24D1/c<8L&_C[4MCccLc
[MP5/0e,V#d6E_U:9^)>;M^-NQDM+]NeSc(28TF3WdBAI^S^c],B,YPU8GSgN8Fd
ZB])Wg0+[I+Y,&DH9Q[,6\9]#CD7;.6T>f)fHd??T)d&A1B]b?5RGHUB6e2eM-P=
VC#a0Sb[@cK>BISDVC2]OJ^2D6,b4+Nb=BC7dZ_Oe=P?8(<8:^)X(MaMbGdTXC1W
f>W+,4?#/J/Xe5YY6>3(>49M72B7@TeBM9J7D4PJPF2XU-B:7e;2;I;OIQ0\L3f@
ZS8<g?\gWa#[+.gK0&K=c[HJAJ=R;KZ];\KKJcJ6]C:cJ/WS)SgUMKPDUc8KIFKT
e=ca]HU5e0D]J8]\aY;1>,U8M3eRTBS:+S]Kf^XHJ@Gd@>>U;7SUeLRNaH7]3.M^
ZED2_JVdbc9[^Dca?F)],:(T&b:Y1V^V#E,1g3IKaaDg/c6O2a7cS6:A18IeK9M)
aQLDL)0/\?DU7]J9CWKJV.&:[aAWPT1c0C+cX0VI>7PW,+,N@a9VHQ5XeC9fB:X,
9=3Q::-Jf]g2cR>9-g9SAHHR1baJ;(XTX1\F)beaY]^fVG4cY^<KBSP52;[Z;c0,
L&OIL)aZ+^ZdRc55;(NGgeI+=PRWQaJ5,C-XS4[M.@CfLN<DF\.dWV_:BN7/2+E=
C:3^]4bK(B-1J4?,^NZ]U6e=X];:6YW;7S+)Vg962RBF(0fC8J(LADA.52=5.cQC
V9^2FUAFKg15YSHbgV>H^D-T75Y;,B7ZZ&\,0+L;#T;ATbS4EU<R6\UdHV/fP^G\
1cTI4S@=+/-(CXN8#fNHAH\EDMNWe1<?OcY3)a/,HB[.3.>X-2Ta1bU(TE-+#NSL
)ZT)@NXVA\.WLATI2KLQ.;68.N]^Sd>U?+J[7]WcI@\@DAbOA^_IgLK8VJY)J0&(
OE9WS;#KHVH47;_<FEGPNdSaYH>AP4-+RW,^>MXP.Db[IX^cK-HXc@>>02U5H<U=
-J;4A=S-07MH//N5QePP#JHDa48&PZ--<N)^8EZ&JLEb>M&,2^)WbK23)[.AB,M8
\@[A>60-=<?XI[U-+XZX-S61]eQaTbMZKM08,D3F#DK2BIX7M,8:G;.I[gY]\LUc
b7]AS)7V#UV\3(WS]([dWEB:V_@&G2Oa94C)@F,2LFID[V-^=;WUYL#_(W#AKU8.
,C<\,OB]GCS&]7Q3&2]aHEK&<6&E^FGN/\-__HFLG<OI/fPCPT(_XcNNa)d@)PYR
483e)AgDT),4]&bPU>9d_:2W#&@SS#XTDXZKNGM6C<1WDU&L@P9[&41Qf72Hf2b2
^g6,Q85A4ZdRQ.RBeb]LIH<#:?cSO)fY39YJeRPaKB8_W_(TG8a/TKX[dGe1(&;U
+AaO8IK18;AVXXVF#cf<bIS-GI04RbN>H9R+F.>WX+FeE?d=.N&K[f]IR8)I(YEV
Ag;BAOZ]N^V.\=3@+a(5\ReGCEEA5<FAg?^N^O(DG4RC=9)3:[5)&.ZGcP6g3I>K
7HHW>6]J=Y&FVC6:W.EY9_5@XGLBU;<6AQY0d7[JTJVeUS+XELOI167SS&>@<^5:
+0VDQ,=g]<^-.c9ICg;I(-:)#Q3<+^<YbM4:ZI\7^)dK8<X#JMe^J4aX_5RNOMHc
KDXZd+c[bE6(5:NX(7,[A,5LF4MRE/_:cQ]4O\1-Vg:CZf9CB)K/+g[#,U(b4ZOQ
MK&?,U\D2S1GdG0-<NKO4-H9);BYWL4=TSINK7aG#_(GMS0e>)8X0&RH#23cae6@
a4V^V/1J#ZBU\H]W:F&_R<[/NXG2C5D#KCG#01f-6e)>+;aD3(E#P:&f]IC,DM>A
M3ML&1<IdLA&gMbOU)BP7f;daCU8Zfg_bL9>HZZ.P-@fFg_#]CW0:]P_(XD3<2(D
818MHU93EZ4S4/#](B&KZ=DPM\bP,-1&K-/]/9E3WD.KB<X#FWb@WZ\\J3TdFbQM
X)MT,:&aBBS[4A:IJFf_4HW^TV[2?Gc<8b&]5G67:QcB/57N2^;da6605)4LPR33
SI:3KHT16M)WVbPXJcTc)Vae>DGF]^\f.,Jc-dK-&&&#Q@&Yg7XCKPJHVCD2DHGJ
K3:^X&CZ8EQ,eQITZSRD-RZD0&(Nb=K;OLHT?ZLECG7[T;K(0e__gSL0H\AQVe0b
H#0Ab2E\X4fJE<>OS<^91AgVXYB?e=ODGYc29g/IIWA[OdX-81Q=Oab&/9a?=],?
^(^3c573>)U:BE2O?5,8(g#HT^1H5Y=V\F>_>eJe.R?]3b.;U]<;RgaB\LJSW>J8
1Y-\9I8]L??R;S=X@4bL(04f_>e>VS0]dEY5dL(QI;[f;UEc,T+IMCFgC:[D.Ya&
2DC>?SV2c^HC?e7.NcU+:=;7\6Z)B;_RFd4ac[N8[K&/@=GY/)4XBZN21b&c@@b+
I>S.eG\^;I<CWUCXc>IXNSCWHD,=O,^J)Vf\Y5&:@DTXY=>FB.PK^4:Nc-IS<SV8
E;C4MH:HL#H/]cXI[W?A]#]8KZ.18bXBXaP<E5O=X?)+1JJV0DHO;W8&;f_>7A/J
7,E(XAXCFeIO(R=b:Fba&CVM_MRM#9g86_3KD]8Q01O3(U2[)21]=&,eE&0@JN\/
a1(F<KQ2LZTY7Xd<]9QMKDE]Y3CXYOR&V9+?eXK@49:-W8UK+L92.=#5#AUT)6#A
Z\:#7@[JdXI48()EXA&B3;A(/?&g,T;&<;.Xf20E&,>750D4(NS@4>W=JQ,V]^B]
KUF^08b\a+#)/19+(Z]MM&2MH[bSf7cbgHY\W8fIfY1[HKe9@,3Je?&g4XJ@(@Oa
W](@W15P/(/?NU3fb=dV-9CUR&@;W1Q&4QGg&1OT.:d+[EABYMe8(88D63(?&SC<
5\/QASfI]dHc8eC>&#A2-T.7[ZG:^3M(]XLR=bK1g?RO=9A_Yg]YbAA89ZZ,(>gP
M3=:.#,C(NRZU=[CMRK1GCUgPDSX51)eBaIE[:@3H>.+EYcg7CRL_W9VBa^C+,E(
0C>I>5QT<3WC/RB,f.cg55a)\>=KU>9SZ/0E,Pb^E72-L>f7H.T9[bRbOHUMT9@b
;8<@Y2&@Q/H2_BN==/L2)0dP5dIbH[RH@bgZBJIC(Z7P2E,N<XSfWe+5/<N-@d?5
.b?)R^G<>/-/ceHTd.N.+d6d8\:)VD;UY,Oa9F&4R-(LgMK+9Z1D5#AHCBAfN5WG
_04SQQb/;EVNfSbcT#,6HHCI.T)DUQ@KDJ4HeggQZM5[\SAE5Pd(7;:SR]\f-e(M
)P/]aL9W&U@OJSWK</BG<3J&I9<XSW;45X#GCW;X:67E+K89dKKRb5N:4<(eAJ+F
)?ESUP5#OJ]<4A)f4Y1QA@34g6+S@8ge^_bP--JN)R(SGgb=b6.IRcgbI-_]e4\E
GL6MIfA7,eZJ]=IOaY>\WCZIP7IR071?]X:Y7IE7/Ec6bJ@I/X/ERV5d?@Xa#;-Y
\-8M=4H8+b>_T;[XM.V-@LV9f08E?+2N,35#(_JE++b[MO(LWNJ;U^X##NeO#85F
:U2TIUg>_N4Z=W53GEWWUROBO8Z(Zb->&f?e6V^TE?J(7XZ#;)7-523^)\QIEV_d
8]M6>EgU<:#1Ic0[@0)SKdG(#4/CXbCS+0e_LC[-XfPXG,b?cP7,CaW+5,\@K7K)
dI:.K[KUP[b_G_\F#F[b4gMZFe9A6)CR86#]JQRP:41TdD#cC_-a);RA-+77/+=e
cf>4)()_XR-/bP3&R&7HZVSge.ZbaFK8Kb93K4O15\MVJWV@LV_69=B>+CP]MNaP
VO):D1#X4#K(W&CeM7-ZDff@d09F;M8N2A)7Yd/RXT>?MGW24<;BWg\d9bL]#JgQ
c(1#6S[^g[fH-8,7\IX<79\4_3G0)^.@1/cbZC8=e@IXI_\e=-68H89[V/GIN8/^
WQMM5T:\7COWR^JZ^:J31+>(17V20U0_)XMg\UUBeD30QU9X;R?::GdR1<OLJK),
B]B)QU:^7GMOUWULSPSGc8R2Q0V;Y9U,=dQC]gQ:LAA>:[.>_gbC?6<RGFW&O5(T
]4Q5@]69Lf/;->(Q6.F1U18;Y-;:?&W<_a7?A,]NMAF[dM40G#((+HJSW.,.4&62
AMF3=&=8XcTH.b7cPGF\+HLFE:gPb7d&CRD:O+A#(BQ\O;0Dcg(M\&;UQSC.E^KF
Da\<X:gIA_+:/EC:RMJ.)U&I_1AXS;#@F]F2D-ILH6_M2W5(B<Hff:WI-XS)V^JB
P?X>APM-KR<bTaK1,3DV8.Z+O:-TK5MV=GAfH942(H0#?:L/C]42<,2\8C]#_[US
5K[b=Ja[@>91bTU/gDPN-6]KS9(bf.X2B.;_GY9MK8/@QOT0L6:3]IYK07VS+ZL_
bbg&gV#cI507S6f^7+.-<FXf(Wc8db4M)SRE&4>7/);FY<P6REI)VNQ&gb9#X,ZA
_GMf4G__\cT)I&4ff(MIgG30&4G9O]g7C&TW?L?(WE,NZ-/d_[?1eFb:I\W^#bMW
gZ;/NUAC2^\:[7MR?]=P:T>&]2c13I0J.:,OfLUC&e-HD5)JA.(Q\S@T^^RL509e
1I\+^2ffX:#81EWP0GfL]A)X^Z-Z17EF1>(/807M)[H</3UYL@@>R=KP,B/^XLUZ
\gH-g(d4^QB]KB8Ub)R:c6H=[b7=8?IO.f5#[C)Ad=?-PLKNO_>,4YTHOgAC.;B+
<H\Va,7HQ3=gG(OgC+_c(X/Rd3AGQ:81VA]G([aCH#9dDQa-&EfgR8G&^HW;CXH.
8;;7W.c[-\Z-ZO;A\dR[^;B;2AeC-&1GdKgGF_)YZ<a^C;/>:aPU)e-Q834-MdV[
CWc?f)ee,&7;aA^U0KW?^Z?TXNG>WEg(\;;RZLOB(_NRQH.=TdIg:Be7YE.Z<S/0
8e.WAL78-B(,bL5\8OaOVA_W(1>#g6_-)ZV#N^34e)(C&0GHgGX3=47:DDXJ-W)=
SV=2V5-QWNJ(bN/DA;X@BN;MfMN86N-E2PHMWE<<1@Nc2:=><gU7D:UG^C\fFDPD
K-Q=dAE7^gA37ZUa&)\6X_K[]f7^-._dR_1VD5&:\+C1O[#/Faa>67<bEf+E]P@&
@AAP^0b&aSN;OH>+=_SA<KV\/^fPGQ_7(HKW@Q2<NW+CQ,XRB8],.,TbcWcU3[KT
c@Mg?G1[@6]eFLe1.b0JacO,fP=7&c1f;=R2CN6?g9ce728[?I&CF_KDGJ^@M#g@
)PaLd2:<ZFB@D[g,/KWWaVZ7[bB0\)IdW3JBLCWK?#)?10?\-1E6ZY#4g=)@T]_Y
PEOeDf=E=]G/JT1]Q4PH24+<P=_?;?G0H@[5@5@7M?OK8a#)(T[TLFb]BVf2ZV\(
O+OF<L]RC1Z&.eK/1X0cAIa<P[.b+P&,@d]2:.K9Z3G0W7PC)(]Q\1]L:1GCgP-e
BR.fIVg>d;YI:D.0M::>EV1])g(7=.\/3W;RYKT_,;#UfK.d+:#WC(&BS#78AEB?
L/0D.L/EScaHg-HRY#Y\;KYL#2D>ZPgS0L.C./0?_/9]N<)NgO5e:-Pd3SV1@34Y
8MW6YU8CaFD3K6LcaMWWA[F>]U<>[#\SDUNddGT..>3;fBRS>>b_:Mc-WZ#ZG\2W
BMfZ@NHe@+.e)W@9cfCW,g?HDD:YOZ(c.cJ^ET6,9._A4RN(W-4-bRMUQ5-cJVS\
PT4EZGS0R/CG8a,/U(&O^(HW(1<f\M^X)@-I9;8;H[P14Q#L7Gg(d;GIaFgR&>B>
[+<4-N0f8]K&@63Q\>R)O7(C7>7KF^FDVD42XLF0cR^<9=NNfZ](XMN@R<<82SGY
g&CJVD@T;.8_YN0FH-WTbb=E3c6PgP\F97W4LI(M]Ba7#N&&),c=^fLWWg2YP1]0
T\6)7/Ka2Z-UeW]BB,9KHN3-H;>eY8;,c(RHC<HH1IQ(eDcJQ]W0I=]163,KQDHG
FDR\S9Z<XUQ&F#1Wa;I;=/@)8AI/FRGL8.c1G3:R2UDF<:Zf7^0N741AWU[;BU7b
HH(#5RVRC@)6Z#DM7?4^UTIIN>IQ,[W+NEOf-CeJS;^;GBf=3+S:FQ>^;KfUT7A]
CR85ObWg/Y.S^/=A&\gO,QUC[SGA(.@d1:cdg<3>GccDIKSI)aTU5_MJS8WOQA]?
3+bKZJT/e5K;7E4d/c;:<]WT-1e.c1D:H=YP-81fKG5.gWY/EWM-(0ecW(<.O+9D
=RcbM@)Ia/H<KPF[[WgTUMg4^C7BYeEcNYLZPD<aMF:46P,/I5-G=E+f5(5Gf5DM
W7A=eZLBF)\c4T(dZLKF(b^+d,_c4K)_A:/<836Z9VNSGJPQ1W4S#Q)PM:2D.E]@
DcW\@+G7>Q?,7\TX3]X0g8GY]K+(WVUca03)ZY.-I+UCNB-+QGFW7:/C-TK[(gAM
37+A,IdD#cTQL_L<gdff_+b<FY&_/5?L8X4\c0E9OP>8VG_G_XAcZ&GI3G4-;L(I
]FeU7J;?U^D9;6a1R8R(ND;C1N2TOfKRPYIHZJ7d,c9ZY[V\c,_Ke(I5J2a\ZY8^
Y8CTC>Jc=YH@V[,0-_PYO@PDKQQTf)N+:2A(/9B>KX4+0&]Na?4F/0C7<08CAZH3
U9.AG4d.048GF8P[3-aJHE:[?S?H#&U(:YH#03H02(YAOM)>N\dG\UL#Eg<4XB@\
L_3N=GD0KR1>-];e\28GA4Q@J7V><UNV8FIB,H2&W:U+5)U49O6ZJfP8cX<J/JbJ
1<Rd0#ZA\C@^F/aB,8c7GNHS^#70<+dP6W4@2SH=.cUA#V4X+cDa=QeS_\XfWA7I
@J_f/QcVF1.6)@0FeSZVPCD#K<U-<4;0I/Gb0MAH0_6??8gb+RQW?ZdNMe+[WJ>/
P\;6=e5/?eP03ZC1LY=89<^1O=dIC5Wc5/7:Jdb=P//Wg-LgYaHc]+925&4Wb4.f
.5C0caSG^3f.&;(HU7R?,WP,f-R8XUBJS>V6aX:5-(e&\RTHF(c]eVRa=\Xa3:NV
^b4.D0&P3W_XU8G^QKO5\CdgW3HY?g>gT_McCd];&R(GZ+/JM)9fd4eL?HNRU:=g
KNOcHc<7K^K-:\E^@O/GVF7XP-bJNI@,QI.+\XMX>\Q7US>e]Q_NR^L)82aBGeWC
a0b5@.)d#]]3S=-ZOM-VSE35S??&-g#>:P;&:EVK9Ae)MbVP[7B,W+5cV/>;PY>5
IGa1THD[6Y]<V)?QV)DdZU@KaZ>Fd0,VUQgTCT5)7UBDdQb:E0L-A8JECWPb)3HH
eb<[F-;5XbI>+gU2KC#I_YXc>Z#U;;QYLK]GT.\<J3QD;cL1G#FD#)HI-c=Q7WS4
E4T\ZXB>FQ3aS88&/R:_>DAQfTZ?\QW1Of)V3];W7PP)Q6;_\BLYKZ/Q-6>?C#HR
^<Cd=T=0\ODb=?\e8Y>1:<eIAcZ95WXaQLY<0)eb@X9[QagINe@5#.WN.HD7cI-Y
^ZH1_?ZB094U653#DC+&CRe_EEQaf.?+S1KW:=0-bN-)H_O.HN=M/+^OZUQM0]_@
MYfYI+@Z^<IQV2J3[J0@0)ED;&:LS4N9f>8f^E?_]9#L?#\)+Y:0JRcFegN@eP;2
,[aFCZDX^LML)0O/Mg8QH^g@^8CL:&Z^0W)6[J)[EUZZTA.=0I6IM#E-MP)^L,XW
,A4c^^25cZLQ4#MW#4IcK+-.,3E6Q>:T2T81KgWg&[:/bK\HbB3b=L:,Y(-f.H[C
MJbMOO@OgZ4QBBg>:EPOd>aP_N).IHKBSB_=2H8bBDZaV8_^X,BABc^\ASL@LGEg
:<Sb]F1D\P]FKF/bf<Bf;>N?],>OK3#&a&WWf2fZaK#Y/6T[V]_,(E,PO5IO\eU&
228>G>71NC&?ZPbJL/^eX2PX11F\#R>Wb^;@/Z=3@dH\@3IfQS8+C4Xe94YYC\@B
bYPYf#,I_1YFacN=GJDO@&&Y#bZ;FRQ+.[WOcWUARbD3VEcQ?OE[U6S@7X,CYPgb
/\]cC4faJb7^R^,_R(3T[V[0V2_:[:]7J[84fKKJg7FT891S>aMM.@_aHBOV96NP
_;2.4Zd>YJ+]@T7IA6M(A?4]S-FeT^E0#@,-g8.Y=33+/&E2,;;\MF2Z13T_+GOB
M0@;cfWK+0?M/^7]G>SC768Aec1b,\CGP(]<9N\L\L9+]T<AY:eSaJ>S(FBB?cM:
Eb8M9@PU8c.DUV)cQ>dBKXVfD&KX.McCR,P7]YJFUJ)B0=D#2YB,c;HBJ>?:S6g^
N)?65\3a0)Bdag2+[VgC=]_4YBZY&0dY-0]<a<WN1,VY^+KMg:Tg+05&+CK62Q1e
JL2JXOUG=f[bUBM+8;@e-(&+M.,[aHR[(WJ),?L>?5g,aMQ_a9G?KB,6R8TIe;>L
fP(N0cNY<-L4KDT:&Vd[T_SYY7E8:WfJ>C^S\e>4a\X.=PUb6-^TX,GWQ/=#FIaD
-(7?9_PY?WdEK9P,G=HFWS-1:(/9U0;3a[40fH,6bB39dEA14N5?J?K,_KX:U-B=
9,J4_I5Bbb8.YQDH>aC_5_2HC);M2(#2/BDM2cPDc5c5>K[VL\0#C>6/8?2=2JSb
g6OIc.]dE^d0Z0]dVV\S=38d:-0JA>>gK1F.#f^<.1&WK0b;<5HV@69:2BRF+H(I
8+B][[(ZOdBe&)=f>=>gJfHX3<(DM:KZg?B:,94JQ>_ARXG06BNdf-V(?@Dc-EHB
N487bCRYHgR&6d@/889>3\?0/^H,:KC5cI9fNfB30#UEI#S9KG/dY<?-8-ZQLZ>:
&/VcSC(e#cVM5PLac1bL3R\KgSY.9a1W.#1&e_B[/cDGcAL+D)[BK1O=&;938\V&
?FIHM_47VH,L64GJ(4fS6Ia>c9P)C0f]@4]A>KW3GMRI)3RUVU+H1:B,O-UJZ:V-
]?&5Qd@LT]=51(FSQQ^e#E,]6A;,668>WA8WNRLDQZ0S9dF]7dHfG^WMgF@98C5W
=I]gbg@\8F2>0fSM.1\AK_>;_d]@Ae[W1K:7,D2J\MR-@a&(E9K<T[>:W48U(>(.
NBAX+1KRY1e#R^(6MYf4H2A958>YIUP:_Y.U60W>25JC/KE2+bg[=657EQ:I9JE6
O=AaH?C#::c23fg#D)B8VcL\B.1)?;(US<e9&61Lf1.,&_R]MI]MFP282AJFB[Ed
XJM]]\_5;_:LH5QO#6(BEICX,^]T3QV6:c6bXX5I.Ce?_8M+RS(+]#F9.G81;J9M
LfYYFV,IXMY4ZbIZV@05&,O6L4fgcB..b>QP)g1ELVQ[Fe8@<.<8#gAE?dbeJ=OO
e#Ud42_C[#Ae5NGUA8aP]MEg+^J5@H:W+>JN+=K^UM>+BY,&XIH:-&NF_:O(dT8D
e,d(egTL]JPSd8<<L747=7Z=&UX4:OgS0:<KAZNV:d-KG_.=gM6dVC\26-H;[56(
VUS259]dLP>+#693B=Q:E1<T/aX?KBT)4VgFN]WU6Lf(T@9IOZ-bf,Hc-JNc=1C6
TXU?.@R&A3I&?:(E.U19KO+>g&H2YM)W:HT7BHLJ3)D6^1<3W.;EL=8FIg2;_K]@
085C@b=R\,BFb5c=CF-(\eb->O.REJ]a2;H&._e(KQ-;[+P#+<.CI(77LF)=[,]A
D;RV.;N06\FE;AJGMCU46bKLXLC4,\),@-UVQMO,B_^WWB8,@7cQA#f3D:ZAF?==
\HE&gINIL6,]>,94L.gK,&Efe5a(XL/@6W3g,?P31_fB-YXVCcN\dM2<TabbB#)Z
ADD?.;,1/Y_W3,+B4SY.5[f^>F0LU]D@?K5+Z=<FE<:WS<C0AF0X,[[bDYeD_2E>
^)e&<&G<_.SFOZ\S.EJ8):793OXRV18><M=b805fEb@&S4R[:;_YeSK39UVCM)4\
E.P&UF?:(:WR7(I/=:c/,0SBIN<#ZI(;Rce_Vb_CJK2#Ce.bA4e+LdG1D?8K]7b?
?QLfSYM<Y70;3[ZZK0P7;J==F4fT6L3]+aX8SDC5C=aQG(;Gb#<E16)C.g&WaeG>
]06#U-[+N?T4+KU2T)]J]CX3VN[3CgMb3ZZFbD&:/KCN9;)T:c8H65(LRF/D6,CH
</IW\;0E[N@Va]KYG3@&\VS]1+GaP2d0\P>LQTMb;+[EVa+8@:Wf(5:\d.>G:<<7
Mb02ea4SO6A,F-)NQG1=X_)-WY1;(-4:BSA--TL2&V:PL#Q(+<M@b5Af:Sg])9Q]
7U59CgNQQHI66aW-?Db_Y<g3P9DILGc&XJVJJPJ1K7PgXD1We(EEY6a&+=c;BXK1
I@2>);T51F<)0A&H:b4bPfSCIWWG7^c4eEYLCb[JC[2JV[9Z\=0.:81YgB5eRXOV
8=6]>0K>IQK,\0g0PK)6=GZ7(Yf:+bB\>.D#CXM)\WZ]J(d-+H=,d-YMD<:F]1bb
C.K=c_46Bc#.O6U:bQKa52#[Y#]U#@/H83](Y9]Le,\28<A]bHEYcYLd>.QE2<WC
]e.b:\L0C\Af8FE@<=+YB(ePZ,8&R5\<[J)A2/</UW&>GHWDdd@+F=PLNJ.//7Eb
SMO?CYH](N]Q_^/J6#R(bLI753ZPF^Y>MZ@Q_H:1/(VDHZ<>;X3)&/b:]+=cb-N9
RQ>2a12:_JG@075(:Eb^2BHF\1FPF0(QZM[Z7JbYa-O(e_YOfX[@gF6INE?3K0)7
<]Pa8TUE9b)CWN\;PSQ>Za.P1,g:A8PGJc@^#D@DdHHW^VfJU6#g2?ZSU0+Nf+Y;
D65#U8fX6-.C&J28([6ZEAGTgeOc=1AU78,=IL)]>JcB^QV>@TNWBW<WBE2GNXBZ
??:->W2+[3C\D0(SIAI;6\.,JSOfDf@09G)_[CD7V?9ZPAY+A)J<=)\RR<\a.#[>
8.0DA@bJH2:X_-<^G-EVWQOP>-9K0]G@GW_I@F#-;8aH?dIBNG^)GS,_&8e,gb;8
9)QXPHL0a;5&13.=95#.+JfKD9d(=_,LF)3N\0.KR#.G:[#:YGGLJX=9N&I4,3F1
4T-\_J^/9V3U+]>R5eN2(UcU&-_[A3L&]gJD)/>^Q>6gZcH2RF3L\JP\?8IO>1:-
:;5c3(62L.R:+^7DBQ-U6a#JZ1/=T6=XdFGPg-C^5H&6_3]d@][X<X8B&(afZSG:
,(]eG6K@U?PHG>+F&2L91GB;1IU9YKRO(eO/;DI,8\,J:30X&7cVb\dB2ZPMF>YX
T^>2T:8eMM)]1f06&I?XfQg]1&@-V#5RPECaWeK]-fDg.OXJI[VPGH1\b0NGMH&P
=OU^g7[a9bdD^QWg]6WSV#Ea.7-&KcBgNOcdI25,f;aY,AfAI<1Y;3VW&Lbg)(8D
b-MD1b93L12IF-e<X-MP6QCM^=P9?.H]\=31bW,e#MAVVa5C/H6D^637K7T&aB1Q
M)\Z]TES&P&^KK:IDg2Me2IJZ[7MTW@P72.U42#:EVQA3Bcg(R(:HAb[]>G,UgfE
eN-<HG5OLdgTR\4)YAD@X:FDSE62LH\-T8K9e+&:DDa4YU3)SF0^MG2dUJ_H\V?#
,)68]XMbQZE&bA?[c-J=1)Q/cN9V1K/1U6IY=6R#e]>bVP)WLVf#]#c@VGc<X>_Q
Na?BRGBD6-L9]UaefO_\D5N?c_;@]NJ:c1;Gd>KOT5=X:0\]fG_:?C655.b5Z[6,
8)\cQ0eU[XbP6DOOL0b#9,O=46FcPS2fSW4Qg1TEND5GW2K?0<MKZ60]6g-KGG-4
WE1+LU;F,KUUb,aO?VKQ5Q:7>C7bELJV/:fKP[.L3TX.,6T2)-_<IO/d:,S2T-T:
96B3#X)EUAd-TH+>N)H_4Y]\W(Fd0eQd2K0@H@\1bQ=RIZAYC67_a(C2^^&P,d:]
5a3J230B\2)VEJZcPgJSHL4Q[WKQf^+fV1EDA>>8YFGM^AV2SG1JUN.CUR^B-B,Z
T2c5Q#/Y7[N+A1<RA:(AXGF+[Q[HaDJ1adLJ;=1d_39Y3bO8/<4CB>7@;(fV/a.)
Q(+G6&aAO>98D3BTY,B>9Y,6WgN>-aAE-D0HCVcOV>M@.N_C7[/f4HU[3@gXU57(
ZX:NO6fJf38W+XUTQQYL#B8c1(6=ZA9[]+:QRGJK&-IeSe,>^Qe@71N3]dPO/fC-
[9](?-NZK+b<:Y4fZe;8d]OA0?/5,[=eGd2/:GR?85FSU[JOG1f-PcaVe@]E^>^V
B;-R]2K.@-a3>F8W5=5<T\]R;83H5U;)dHB]a(.BD:T4XE#eD9d&9;XBAL50A[?e
4/@7[R/5fa27;+=J:.FF[/d<S&L&Z^COS(4NgH-5O/QH-,J7J7EUARD3GC?&G]\2
3cI,ZV\WcKS7DJVY9VU9>PG&?GE.RedeN9::WXRAeIGM3R1:X8\YX9GPFM[A.P_;
:5_c/E]JA:UQ&\Q7OY[J:OTHO+_H4<f4#f;5CDV=NEK)\>)7KVS@DagAbF0I(G0S
7#-.c09b)8X_CQ9R)d=dVO))#\I)IV8.3MJ4-QVK#NcX6gHZTEATD9+EUf\+Eb&0
(9N+825X.3@MHRK_^a;b89M6.WaB&/eU[ZWW;AHBDQ8<EG+59Z2^HaaHUC=04MXO
\Ke]91N;8I(\IW2VHWKdY[\G=XCIC[P?E=9g<-C/9FdOd-,Uf6]7e0&28]/@__(@
MXZ+==&0.<+:1dFHX>7gGSM17^QZcFN4W5TQ8#]\>Jc?NM173?^:+Ee^5\BJTFPA
?Y0+)0077:[=Od/04M7#YF[bQ.Gg3dDc-:)]X17MWbP8\./W]bP0S\P)T;L/Be/^
/Ie:2<(H<&<f>3\8Z5aH-:dg[K4N;_dY5;Q#_@PF^ZbELfAQC(9e8)_P_1Sea<^/
-496]QF(QW0PLIeNa7@S9NE>5Gd[I;)RY,3F^9E?,,QW9M&^eC]PNQ+eN0(V[)/G
YeabN&K+H8CEPF:9W.^1ZJC2O3#TS_VU/eY&8CbDUU_^\,MG:-VaGSA>bMJ4=bd1
f\3VM)?@.4;PaD<V]8]aWO4+K)\>N?Yc,M#Q5_^XQ).7;V;L2/GLI58\G/1QJ@MG
Qe+8N.#<0P1;/^/B5AFRNM\P:L)>Jf9[4<dDYF_YcfP4c\PJ&4^\aCbPMV(T0W[K
<@2;gNFbR#a^Zcd0G_R:KHM6Vg1H1\8^)<#BEeE-ED;<.f1W/W=O,DAWbaZ+67E:
>X6M[23XSd:Jc4_EZd//a.G;.LWA?J;c<TT6AH.4W&A-@>>I3_cBZ.C&F5Z3QM>)
#48K@1JC5_]ea6Z>WM?3KK@cM))a(9bgY57\JVD>SR_Sc4C9BVCL>LOUadK69RM(
A5T5(Q>D?KU^79M+QV#=)1P+RY8eB3CXc(^:+T6)[cdJCH34)4;.2FK8TUEPUN,g
MPHN4LX95E/L7>=5IcN,fZ#-Ld+4\ZfN+7XZFWNM:R3\.UO(X<\3FWd7=Lg)+@44
/SB3-gN]=#I94A0(4-^LS5@#XP<ZNDC.33R;QM\]@Bb2YaFZ7M(cUb#)\b&ARMX8
4_Q80aZDOU.IIO?W.cRGYXTU1KZM>S^1,;G0CT)J=,R3/g;LL_E:[0<cCR[1)aX^
PQ(&_2]WY#J,b>^XXdJa^FEYLQ5<P,XY6G\_e\[+VN>0KO==Q<<H.;J,2+3,G&6B
GJbfYE(P\+HOP-?:WcQ]H2?X7@Ze(4R8^-(XJX\@V&ABL5:-H:W;a(05aG5Z5X&[
I\VcIB2:^4S:-N5+4eGd6)J;.4-67f^3F8D(H>4c=_7\]]]F7\:,-GcMLI(EIK+I
SI#P-Eg=(3GO9REXefR9f,_+,)PHS;d?^44.+^?@M6UQW0M+N74^_cHH4L)[/;++
+]D^ECYa^aa^J4T@##c^#AL#5[D3S6O:bQWW2ER:^dKRZ8EaTW9bE/@,YUP=>a7-
PN[OgB^W-f.Q>RGI44)f_QQQ/>U]E4C@>FD;ZK+1e?d-L#-LGJaS\f:V6/M>:K^H
Z\f\J\7ALc8^KccI)(:Y)geMSWISD8L:-&(JT(+=[IO:Ja(&\5DIdUJ[^eCWD3CM
gV1f#fQ4<a2&KJYdRRCK09)bIJR(G1S(dB;B#05]C<OG.L6eMP[ed^3^eXWP\]fN
]b;Q^dd2USV_Df=#65AORWCG8M4f\]e/EdT@d#A?VZVOICT^07VgI/H08,_8#86U
g#QV(Xb:T6I\Z521C@ZAJIbYNI-DB7DeQ0fP4gG=#[gE;Z/QBN,.Qf8Ng_-.Y#g?
XQ3(OW1?SAU7cWRHG=&W>K4E(BfcDJa#\,cbGZB-LX.F,;[7;WNg_edG(1>CE-WW
4790SVXC-8D=#5G17[PP;;(aAM]7Y81dbZ;55T#D8]cd,c13UQ+=A4?@Z)_14<4G
3U]c)(&^5+M[_6_/ADe^DC\a1Mec__JRdOX0KfA457C&6\9J+>/:]X.Dd6ZBTU)f
b<PI+7AFC/S3H:c&UEJN3710>\L=1NaG7deXdTZE4TX99/A,Sb4&57FXIg=J1FK0
<G(SAW7T[^JH/2#M)47/7M7_:_KE:&BcOB=R<IB0(N,RV[ObGJ5NB2Y&T/9PYE6.
>&V#c1+#?Va/0^[Y>@Vd0H?aR\G(OC,aR9H#Y00GF>B]e]BLQ#/9T(3DVIVJHP\&
,7FK>fK:KRE]S]^[R?15/GP3e_ZE#1SEQ#@&CB:^7#C5e9gTIdJ=:.2OY2[g0,TF
U?_?D8CDE2fAg/_7G40@;8@@R5bLD)VUWbRUD3/IaERfM#PTT.5f+7M@PbSLS+aR
:Q3bG9e06@ST#FaOW3JD?]JBQY4?V0)=N>&3e_B,8E;dH5fD(,5bEJ[\GMNQOFeP
eF,D=gd16L3G)FG4L^E[?<TXYg8b=9Va7\O#RDU#MgIWVK(eJH_A@b9[fZ+YG607
+M4c0ZP-LcL3SX-B9LLZIQDW/1XYcETT3<S@M\2Qd#3:9LfSGMTgP>B4M4S?WGBS
H?d1D_)GJ+_.0M^H-_EQ?Wd,b=a<4>>ZK<ZM]>=gKU_1Xc7N&^BM7U?/GA^HgJP(
+<2@^4Ye2O;e38?ZZFQD4/bSOV.#G>WgG@,H5AN??(3;ZK(GF4.61V\c]2S8@,:<
\?ARgZNFJCEc.d-H<P&Q[L^JW>9TKZ?8LP?C)#E<@O\G@6JI:CEPS/VSA0C?fd0c
#]@f72K;E792<UT6K>\@8\O_2Q&OTB9[Z08T02(bRB\\AOYaUS0Y7BU5>O#JW01?
.=2=6)63R\T+LH4QZS/f1,M>J@gV9Z^PKSM[WSc3>Od4@1,]dd;F@Lb97^E26+Z-
X#H(FcC.B&<_MHR93K2>FC>)>D/LGQT,]2U]HZO[[D2))TTKSAD>&,(1JLf?W,>W
;;YS,D]8\<EE0,BR-BO/5+@E3\e.M&AEN@XV<#[Z8Ca7a(CR1?3DH8E?]N?^Gcg+
G=<-BA+4>ad&-?^5WH1gFR?5RAYCR4V]ZbH/+e_W<6@K-Z<;^A6FX[Ug:3PP<8P7
ESE.5(C5K/@^FHf@>>.AO_eb8W018-gM<=Be)MBM/@76.-6L7R.>/J+N2/S03QK&
A+/QZ/SUUaJAI&G9]c=e_-=@#H@6G&^-3eeW#/(S/OT2JZXI^)=B)-a@[WfMS6.P
A@#8SE#R80S>0.1\TZD4HX)X,1(_,O\NOY:f8VVBV;CK\K>5UMVg)W7[cQb;[eW]
_7Hd\X<c3\XXRfg?I?;JA1^egMA^R.YeKEW>SVOHL(Rgg,^F>/(/Of+<@/+AWM.b
Y=@S/H):XTD>/QI<I]2cdDdZTLQg)CRb=E8A4EaK)]DF2H;O)_UBf@?=eJG&2U1G
]^/J&?[A7[JI<ZH-0aR\@^bH-dD<Z#aK6FVODO2:SP?>MX5#KGYGbbeG7(T_9P\F
K<V[8NT<#T[2PU:NME_fSJM0JI1C?]>+V[caAOQQIVE;4YFJ,\WU#T3Y^<?)EL^g
V\_f@e^MYTN4aC[D8fg=^#4\H]1E.XRf\e=K;@S@MbEU+O^+:X^&,4C=.QAEC0&6
-AEJ)UC[,CG[aFK]LRfB+SF2_@18g\UV8V)]L-.bTJZ,1)DVJ4Z=:(b_C7,I(b\5
X;?.ag,+)1&fNfVZYU3@3eH((B.6)<X=>f=@X=&c;/aO6FWJ^Q9<L2UMRPGUD_c,
,+aV(HF/^#aUYde#d/?T.f,@UTDR@.Q\)3;CYW)Bd)f\&b6T<@23BHNG_>L.2]^X
RI&3g>dL6,1&CZ]ZM?DE,U=&9\_6SgTRb\2Y,f3TKHB1X9<.G[O]T]dVP[O8T8)P
E3d<_I-S4CDWNR\\AA6]01-^63C:2_SC.W=aHHI<>dX8E[H/ILg,&@=_(+?:Tec&
\DV5OQ5=\^MaYK_(1>4>1Yf-HD51).]K6,d2^2XRRY]S8/-,^X-G45KWK5)-)YW_
c;0I#(-b@>U.<ZK@a:8Ye(d:1\+N._25@_(0+4EC5LYf.(_3]V&M?E^X@/LSJ1=^
MRb?Zg\IO7>)K#=@=T.AZ(@,ITb@4W]?5AXTZY9I.BgF0Aa5@20UIK/gYA&R<(+)
Z[@Q@91f64^RX#4<E_G#4^0G889_RW@,])9_LDUU16J6BK=K,F>OM(Q)J74LTQ]M
35cgII3SeE;#,dB(D5GZFX?E/[SVZ+6X-(BHA(INKe98+OK1/ZJ;21Ee/6PIKEdd
\,AP?4+3fNU?F<79GCXOX<UPU.#>>LY28KcfA^5e<MMKf(.Q&2A<T.H7;<E8GA.&
GA;P\7adP0U/Gb8#>eVI8712gL7.L++1QbM_IH[b4&4b3Bf-N7e@VGU\[4a17Zc-
1e\#O>Mgg;+,^O0/JFU?b]&A[,9;10NF9WN^&;),bCES/YD.d_-=CGC]ZXW(KE4E
)6;<&B1&\DF?3/3=X>K<;:DH\aL.1=gVB9URa+Z0eF7DZ@#<70M>5.PgRWZ,U:ZA
<06KR,J8M_<CG2cAMdb]C1Nc?0.dR&SfPJQ.#e-ZZG\]_D&E2VW8d,W]<GdE0Y+O
7^9,JHG@WA)JdNJ&XfI<fXI1]XR_-AGG@V@J@cU4>8X(Z4ZHcHTF+C6M,6EBL,^J
2?I(U+ZPb:R?#&3dXUDJ)dAX=L83/Fg^-/].f67STNeSa@[B&7^f5VI+O29=]MY1
2b(+#&SYeFK@)4G)CQSVeLddI<4XYQ)O\GU2H,LQEX\]W^)^9cJf,D..I=2aT<8O
EY&5:#]576N]7DW@@0RII.^BH7P1QVA0dV1TATT[[]TXVQ^O<NM=0HJba<fD_AW+
GcDE0a(8Z0>1,4@.1&HIW:]aVO[O4@X]QF3\<CY6_2[);CE];2YgU5ND#89C,+6[
25I?^IK_A;];@d?HgL809A?IQc(W(0J1A+D?=(FRH/R][PI=0DM?Q9R7(076KZYE
@FcR(E;ge[c4(R0IPY10M>4WTS:E:++0]EXXW>a88S38QK^<=PAZ5BEP>Z3(;QT&
CR.L>3cVb_^RQVIf96>]\CKY-&^\[c6V1DGM9cSPK;#;>ed2W&#&bbZHQ]7+GJ(,
LKd_1V.U?cH)?;e\0>&8K^cFRXV)X^W6J:Nc>ORX=L+QUIcRfYT2Ng9VPBMSK[9U
g8;\5W3Q64EKVOK,R[0#T+c;8N+g-g9X2C\\@5acgdO7A<V-/EB6Cf(U:bI\GT@5
5fX@Y=1Of+1JgMJ+>C#39a(PKV[>@H[MdBXg]?I/S-/)W6e0G7AXg5PfQQ]f=P]I
Ba]FHUeYI0g7e3Y./b@bJGL+,S]dE/^]O,6_9OUSJVOgGd^)I_?c#91F41JS\Y6N
cWU1O<.10+)dd.AcDL>]-:\WJ;,Q/I8?AT1=HF\TeM81:QcT/dV&BCFLL?K/Ld/7
d0/<49;D_H?FBN/T]#9)3\)?89,^_AZd#DL\3fa]W=H&^(RYN]4ZL#]1;61fZV4-
2JgT12FU+YS[_R)]DH,4&;WTZ[?42\YXTX0BP=GgfgfE0.FN(QV6M9^+[2>e?;R>
GW5g#?13Mc8X[b?AR,f9[J23YOFTZe;fbe_<b5;1[SEVY^BU@WRabW&:0T@^aH\6
V3K]MWCFM8,M9G3/[J,^eE5C.f/J#VV_J@441^bW7C7S\<c8gN@OXLff2R[/MR]N
#KdM.B@NX[D&(?JYIR6.b2LSc9J794Df<.4<,fb^DAH;fXV17I9P=V-6TDJ];d5&
AgWV=T;PK\ZTI=MJ1YNSB#]YUg=8\4g/c4ce_ga/([MZOY7g3Z,8A/_(c89.>)L#
1K[0aW3;C9)<ZC]McQAW0?^4e>=S-=_NdFa=9DeCfB7Pb^NBWQ0JJ.g7RPRR>bEO
/W]@_(8MB4U1QYU54(=TK9JVbXJe?cO77B\O7O):\G8,RC_,1P-@V&E:=FJI[)[E
^8(HU,c)-V#36MMG.T=R.[V7291>,3-#Y42BC]-a)@):Vb1>-:.\G:9#/[/<1fWR
]<XOL)WDYg6+f4X/UPPC^9g0U9\;8bD;E#2,=:7.@,V0H&e@L_JQbHe9Z.f>QPF0
KTB]B:Hf^7>a+aS^G^1B>XNK;(,.4H8:g+BDNA5B>NW_IU?C(_&A<B\1_6^LASIH
2=XB7^0IcVOY2(C<J#C<YN1AXbJF?DO]/dEX)]9U/dLDUKe/_P^Ub:@bT2e4HYb;
-<7:)9/[DIAH[C2V_4&A(L-G;Kc&-_Q3Z9H49\R<9G7>,?Z9^25(G?g&4GbRe84\
.O2B&dJ4CC6CI#cQVR=N(fb+K.+dFA>)c#^Jb.3[@>/Z5^a.dUZ\dbPcI;g]YX]3
8V1IRI1P(#AIQG<C>9&gX7faWg/B(YZD+f3eYJeAd@<J;D_)M2T,@C?)WE3YHTQ/
]X=6^JJE&FNX,.IW-0..bRX.Xa16P:a4aC2[5]B<c7PV9&7SdI@F^49[A<3U&L;#
=Z[(F@G5[1JTFU._+-eM(8c[b3R@I\gWRVKT/g8J7be>@@UH1?-F:WLKREc]>#&(
-YD_^SHZ8U+/WROQA+^3e&:Md,d9X@3-J>X6LDH8D5cA.V+.#]3B7M^D6MUW4,/2
BU-K\>\f\5])--eRV3c<LSL[;QG^Ec.@bQ.\(X:,1NFF]:CGPF\E3bM5]-RYBHAF
<I.f+eJfCU2HPT)UQ@VNaC(8gc:P-+KWFZ(PQ(LXHbDf]VEcW?7aDa<DWY@(fU+I
>(fC37eF96##)=VG4&Kg>\49IZXT6)2BPgg91&7SJURUbA_XUIKa:KSCBP^?Y.f1
Q,28E+@<O\=KL:IY2(>7\4RPQBW]Td2ZDaGWeZ;-N;,DcT2V1N1ddO4:aW,Ma9(]
+]#d,5<07cc4TQ&FOXYYPI0=S4\4_-/QKgS&7d+3A7Sc&Dc/]-8EXV51^IM9H1#=
;>[S+I1&BC4_0^+9(&(N?\_QdBDP_56:=+)G)&U2gBG3EdZWY#X=AON5G<C6Yf&e
/EL<cf+VGVc56.FMB7\,_/EL(UaGV4=FC_8TC9D6J;/.?f.Q>\]J&>g)>QG)>9JK
e>L?DNO17U;,Qbe&^UQ&3L3T[?;41A=8cTO7Y?dVFg1;3Q:]I^D9IE-KC\F1M#M3
U&g)9#Fa_]gMA&F1((C)=Q/FC\A0>&_;G(M^SUggU(UbD:X0QU_0QD3XT=+.efK9
S(F&?0H4N(^;@_K&]8#C>cV8WT9WTH\b\U_9>HWI2^SN15/af22;D:&b<4-D4[BV
I)3]JLX-L=XHJN,?Q&#<C>3AdJJ#+g,IZ2TYJHB+d0@NZY_fX,-X(=X5ZO3<8+-&
faF;9E3WUSOEZ[>X.)Z#J13K^);#,2OEgV64fF1VaUU5@[</E2CZ,e;Cd-QWPIXL
B8NYd;fUQ+22BXUaIY,F\-U2N;DV)OC#V.L.YYLMVY?,V34OV./O<JR\3QC12X?G
]HNP=N:2g#6-&./]7T9<g3IbC;YL:@0GL=T6K,3MRXM^[0)c;>OM1.]96#05N/P0
JDQ-X\U=GCD\L,M_;YBb1?=I##TP>\Mf5[6_+=Q;,S8gF6Y:EPOYT-0cO<0gZ;SS
-a02gEOO/VTZg_HdLLF3@B6fV:GMfe.,ESHTLZ^0bMJ[5K;]Wb]L_#gVW0@DG,]a
RE&[6cY3/+-GdaIO94f\NX(0[+;G515P8MZDH]Y#@^OaSEa?V\7U?4;I=MN1I(;(
e4QCKRf;1QEXgc?d=,AUdFC4U7<=FgM8.Bd6L>cD&g;T.[8PBXaQ,E<RU;98(CPc
(_2/_M^F;F<;I>eZaQU?@8D^F8R_K(;\]eL1Ff&/9R]d8Fe1W8(&,]e0-=(Z/8&D
:\&(SR\UFP-L3B,6&YaO_BRd^@U56^SD?fK&(JEeD?BFbb,19@1)8E-B-K4f1YQ-
TZI&Z&IBQAL9F1?cQ2L&e_?c:UQ5HIYW3YLME8G4C.LR6]].,NTgUe#^d=b2521E
O?9(_RAQb7X])#II6H3Ded>B(_561dd02aQFR)b4JBRKVR;.]V,ae;+-PVSY?[JD
J&b2J^764A1d&8?D2]7DO)ZEHMZ7/Y\F464T7WV)63_,2[7A+@59A<(=.?G_DF7J
/W-/>V_TG(ARWAEADM?gI)/XY=Wa#e8edTcg,=4RZ>SMS5?g,8ODaOBK7,.X#FFJ
25O(d[\O8?d/NFc.]);+:]bDZ@C4DO38dI]V>]8HVBIQ4bPJH:.VFK&+JX,@N=E0
:+D-\90S]/ReTRC25<]<Q3GKRO_JQ0T1d^f-_K_G-J?BY/B,3K#E7K]CAYIMJ8P5
Z_7RCSeH[(C;;B1OX.DPb\@?MJ27CfP+>2NUdTV/MI[YMJ;]YU7^53\fT9Q0W]Le
gG6=OC:[a^NB]Ed@Dd]#+8gDHA.gX.V=7g:CZ0\;X[X/1KC0U5f>?VK[0Q/V&:9d
+D=LRTXXVd(WBO9Dd+(&1a20]UZ1>D8,EL=&QC.(NMR4#65f3]BURAK5eF9dCadX
+8YdgD.Zg4aMZA7gF-P+8QO+FNe;fTXV7NH)9-Xc&4;^N:E7W7b1N+21E>SB7dDE
SRH/D&+M/&2d]eM^#80?fW_IXO2YZVO]V-XSK+8K/ZIM?9?>]0YgAbK6M+,7K\.#
PH?2Q(ZOf<9Va?7&D2:UZVe5)SSCa?CeH;UZZNg@Tf3Y^P593/[T7KW@Dd(L,:Z?
_Q<G(Y=MI(ZIa=H7)#UF>-F]0?WgfgT+J#+Y.J0^SV1UDQ0I&@,[QOXN/4eZBX+[
QDS9^UB^L099UZeX<?Y8Fc@XSQ0Y\X&O:Y6U6614e_IVQa,@6(Ue+EP][KCe\TBQ
@<I^9YgWW,1PVNCG5C_M/O(WIM4X9Y;L7Xc1b./Q-g+S(UY:e2NTV)NdX0I)H,ff
f;].@Z_cSBTNELfHB4D8J(5/VP8NAST,#e<\G&1Ig5(?.:FSK>;F/?#gTJbXK>Pc
U?9EHQ[daLbF_bPKfY>B[Fc949^I7R8F4_2bX@QQM_(V1NABV_V&dgIV#S-]fKT>
3]T1DbG),1\V<8HYe6VC,M^1H@]C)NXE(@FQ4(a>OXf>B.+DR6W,.P@[^44I+<aR
6P=+];=LBNaOI:O24;.6AeV10THZG(:)AEBc[J,A\J3dLWEVI-HBI@8K^RJV6\78
e2&ZL#<U:X=Yb,#=&);X;b,8-Q-[883&7[ccF&1+adV)J?MU9a^RfKXW_2V9E:Pg
aG>153ae9<J]YecLMgQAd<2(QCBcfV(fJ]4&-BBB2@).7OCTKMO#(/L+YB2F&@8f
I_WEAK:g[ILZC>a0]>B&f6X9XdS63F9]:?RJ90C[?e#MbASf,f6WK&8;NRA5fN5&
[d,1K?&)TQ<-<5,[&NGMRecW:b_M0#bg1J\G4I&CdP[X9\9LbC/=-P/2fbSN\YLW
_[?f3?;.MOBU^17&_IE_e8b=AP19P5+.1-]ggL4W7UbNRQK.We&A=>&(d^;+=1;X
dW\8CHCMeN-LIGHU[5+69NGBB9+e:290X.83&^:<&c]_-AZR>NKUaKVV;1=]CYU7
>:[S9+BI3#L5V^/SS9^5>eB8&O[Y_YP;cQ@92A+O]6V(^d9&4Z_;YS5d/UP1:XJ,
YG75Y(0a:MFF=Ec61f^O@OC5EVB8V^N,E/G\@C:Oe;Jd\NFe/e3MfKZ\WEGg87e-
@2PGL7dLLV+PXJEIWNGZG/;(P08+)Td)92W8:&3CRH/>2Yf&LIg^FFd5_]23\dEG
90VbXM:\I=8[=)(\I:(Q/O&\VQdYEW-?_]7Q4>I<4.7fV/R_:ZaM]KCA4D=8B4Fg
W;ca#e1)AL7<eORaY)9Rg3SePVb7<8I1c&0[#TJE\Ba#-1T=fRYE\[R.fQ?XVP[0
SS.FCEgfLU1XOZ(5:O1^CCN23IbX=@5EM[CSM]VT,(-Ab(OB532+:)Ff]48>FL@a
9XIg>1=/S+@-1d1d<+/GLgW;fcf-ZN26(0HJ9_,SGMM4^)9G5</9HYVTf&^,f<GY
D@V\G-[DT[-J#bFeW+.Gc\dL,VN^4eZY:V;H8-]YB[_4S(3WOS9LWMD#(VS,OVa[
Wf3I=b,gVG=;.#TOKC7U6F/^\R@1S-^QEIEC1AK^6WI.KM>LAAZ6Hd5\I@;4[19X
WF=e##Y2ZSMG+=fFHb(6bZ7XV0LXPDbFH\eV-;?FWC/^V-Wf[S5U9Ya6A9I@fJ&J
Xg6C)R45U2Z5V[G?8bC@TFf_@C#OJH5O;&/TR5,1X@S/92/OM070-O.bX[W-f:46
DdHRSbL/.:=OR/EF<&Me.5:2O0YK[#ag+=?UUO>1NJ;:K#)XdFO3EI+<;XW>g?H:
+T/[Bgd)J-YA4fJ??K?AbW1T<D))I1=JI+\3;If2_L9;G]W+.bCOVX0;\#F2P#UV
,BC&^;0;W58N=0=bd>JQHeVI)P2B1VZe=],_/)HK@BL=0_QKW]d#DX,+^/-V:Ma5
eQI;@[G\6NXS.:XQ)WQ+PKS2(]4Bb(K7X1T=JV-BJGR;@D6e[E?A47CRIN;-B07_
AD_J<S8a0&9fHDV_D@5T[M/]35C[_H57E4<20H^SaPf0PB?@.[,NO.()fWfXSPXg
,9>T+g\6\BLEg=1GJQJ;beMO=N6CM1B>:]f@c,M]IcZY&[;2@-K1JR#a:1OO[EMD
,7VT0>XH;L0d?8(b;,(<?1WLCQYGHHc^04;0>2,6XE5@(6W-:GD=B@b5DbWJ4_FC
\O#P0ebeJK+O;66Yg4QW-0Cfa9CKb<#_261_:?IN79c<W;-HHfgQE>N=7X4BRKcd
2dLP?F]T=P:O&QNH)W(?JP-T674&=GFY4JDKR)aPI?=7D>YX#@aTW\DCEVKg8cdY
<AT^<R))BDM6dd,b#O&/@_H.S[@]B9R/fHYgd8L,.)dI\LFAe0,&,8-:=5+VW7Fe
Zbb9I8=;R7:f37,1J9&S[10f@[XTY1,;5Y/U+g.-G44_&b-?:S[]Oa]]Bf0f0&HF
F9G7@M)eYERW2W6DT7JK;Q#967fd7#g&dO;OXR\Q9>TPcd22=7MReG@(&E.>2+TB
:/9&1=P7-a>a><EROMd\_MS58Wbd8\B1cTe8^@cKVbHNc2[IQgYTGWZ<#B>d?5,:
YZ)WbZ7IG2OAMCJ8K5bGZf#)g\gG5gP?G;PJNW-LEa)B(SGT07c?-1#/74TJD71g
dD=EB;b&:5Q=2H8Gg(@R_]5YGJaJU,0ZBM,Rb>Gf#a[C9:NFcaX\KY3IW#_a;DD,
[,H,3YgEA/E&B=TeTe.L9.W5,LNNZ>TCJB<_FdPVSeZ?,:C88bO5Q3V7(A_2TTA3
S80MC\b&@:_aZ[B1\^SSRZM?gceE1Q+./)[NFQ&P3-2c#6eMIWE_V(]+QU),PB7J
M=Rfe-\V/;0IN+39e>#YR-cRLSXI.E;)2&AI>]0@\#J,D[4V<(AJ9Y-?PbDe)^?1
,S?X?PB<-@/ZJ^Yd#43(0=\E4Q@<F_/[.8_Z8WS=RY2#?_(=HUK138C=[3.M,7(3
V0_,7>[F<W32PAdRP?P;A+)FN@F?@_JY@RIF+b=e@R1OI51>cT?QHP>]ZT8:5FH5
QFI0=WID;IcFBPU/^VW.O_5:#9CFd&:@N.6</\5ENfbfF:A9KZAEd7S8AD^D-\RJ
eK/+1AH<SF(<G4DF,&+TF^V):J4c[KIg#_M]V[IT/XWV\?>T9U[+(B)^,0X]fae&
QbV_fMP25Y5RFUb:<SXSRMZW9.3ZFOc3e5Jg7]OC#bU-M/+e/&K6QLa\A=@dWLHe
g>=33ZObTRGS)O7/5:_^O/L<@.N3F?,7M)b[?e/7YQaN@gY>PP,-4^CfcI>PNS\B
<4/48^^.&a#NOP/+fMW[4e\B((;e>Bf336J3LcV,0B79d3NU=[]8ILKXF+]?PYQ)
3MZ(3a7e@?[de6E2)9JC,A]S?6EMMYZ0L3NC/e:_BR2-)BAE23(.])D1#Wb=X+#G
V47N0dF]O2@>G>8PcS9dc]gNOCUVZ)Rf.\Q^^Y:2YaJQE&XKff4d]SR<X&PJ\Fa(
\D8Q-W7N,e,Q8RGLKXBVARdXDJ8Z0OPDMF2E/--(:bS1SBdI,-YfZS+;&BR1>g[/
XT=<RW8cge14?=&\)V1BGcI8UU32A-RELf7<KZP):#_\]aK3L0DPbN[<(XZd);\f
3U=?Q:6KO/S60@F_7b<8=@R@M)558AK,>W+6[VZ#,A9S5FFBT>3X-6\V6E)HM<RS
Veecc8CPTOF:;K([2e1CE/BXTegD#66S,F[XWM,1EVHWBWd)@67:>0;cUa3&LgNV
=W[J^0O,1OT6^-G\c&7Qdd#@V]-32V[:[+[<&DVF2,TJQ+;^2DI5>F(8>#\CRV+V
G]^G4H9LDU-82bU<c6_(-1QC,M_1Z\=\M(,BJ=YcJ)&I5>;/N/29YGf8gVR:2d?F
_4ePBE\I\\Vb<2&38.[K&Y]BO3QF+;(3M3NM<&\C[C:Qe=0CD2Ka)8E7Z:DOdT,A
BUQd@9Lg#g1XKJZGVMd3>)&4TO1GXQ=>XR&fWK9eQAT/O5-XLFJ&8)9aIN\YBAgQ
<2RJ2LXPCH]EZ#;L0_MP5@EGE6W\3+5?Y0I1(#RI2BU/S_aPS5e6:0KeOU&4,66T
?P[UAU11G[a=2P;FRA3aTFJU(3M:53(4((XH.g1f#KUA-;1J<f8D>](GW^9VP6a8
0>&OSO[W&Q7Q#X?;ARb=a^U,cCDO&&QUJ1M++gTbN?1K\I1e;gUAT_@(\/I_5^4V
ed.L^[/gZ1-J-S;AOE:e^Z+H6X_UTD#XR0a[@05<\f/=/J+FGF7bc(36YLRN/[WU
4Q0VBTGT]Q3D/KNSZQAWT6d(OL1Re@?M@T,]=a_ALH?77ALD7DT&PRN=ReRYg[WC
T3@G0;P:d(f1];f.EKS?]IdC-]McXFX<,^,.3c4[5Oa>?6e(NBKUC,Y0Q=f7/(U/
,=INIeaM]^UBe;4XbWH\/Hb1FUbN.:4+e6fF(M;59I0;(a6?08KN/;XVGdD49KFT
Bbg@(1\8+f8?LTB/[(]PK,fM3CT]M0J\?6#LOP4KQN9R90?7]#WHb4=N)2TXcY4/
@16&,8Jg3M>?4^?Vc]QL.VGGY;(G_22X?YCBC[W,04B]Z^)S?UeGSZ-[4HIK@PY0
1Z7C?SZ(Y;]LJdLg_8a4SM2SJdaS2\AcI_\OS[K07:.763_RVFGSE0UZIP2SbB05
Uf&eUf;e_JBV4SNP_;ZGAF902HZJYAS)aa3OB(8P2RW+TaYCEab]=F+-[7GBb5T1
HXVDLH;@dO;W5E7GC>g\W76]]9(.0a5XZ.>+32=a&2CNM&YdSA(XO#-.;)Z4HPKC
AJT(G[+]2@[aEC/a2A5,->5;K0)Zd7Wc:V(ZLP2O2F1Y=7:O>ZeWWdV+XKI_c1TN
TGL=[=G58ENJDR_-#_c+15:2M4;]^,&[#Tgc3Ra]9G-A>[93)GITVK_<DV9IPRN7
b>)WRJ2)&CO?FNFE]<G@VZP\6C3b)K(+b8X\HJQCfS@^1TAB/@D7D3\<I.gTTg[_
)77B<2Xd-#J5Q>U&?M1/&J?U_e,ddD3Y;UHcY.A6=b@ZQW=c;]e8)<R_,,3W;Fg\
&@^#.JR>+.BB;&fO(AOY8=UP>CNT7QZ)^T^ML81ff,(;PIRc)+E7;-^JQZ(T.DUP
>>e9Q?-a>&7Rb;2Q8d#GXRY:EQFI++XWX6aVTO-=P-SGe_S?C,W(]\RY4?eM4M1R
N,NaeeWH=P<VMB]6e4;(O_XYZSJA>47)H8#XbaZ=0F5e#E0LH6d<]g5C.S.S..0V
,O#cSG@9fWT3VLbT,)HXACF7XadD\ON0gOcD^UYa^(\/]cF:-gLa]fe_-@-_94EU
0.@.8[O\VaA:YB1:N^O/2PQLL7:-?dP<+X6ESTK.&JS\GN\Hg_e<R9?5P6EQI&B6
])D-GB@++V[M#@@H2U&McF_Wbc^W8DN;L6d9S<HGWd&C\IR=Ic)FfBR6]NJD15d=
MEcQ[H,63#A@f1cHY0HY,7O/Z\CO09HW/8_,Df.5fD,VBcW6V0A13+SB7+?XXCY.
bR:#=5UNK7-_^@OI0(B.RLfS(ZC5R.(/Q\PDaXMZ&dYVO>&W^03A=(8DR#>?PP+Y
0H?IE2-<>PPEL2-JcH8e?[GSaNX35RRNW17f;6Y\MU)Pf[+<QN<=+aXg=ZQMMQa4
Ke]PQ>9g;ZJW#72:MAVC:[NTcBOK1bW(-;HERYVcK[-Z:C5G+C-)RaE(6H+J@C+F
SWGeac,,W\@NC6,5UB>]6F.Z9/4Z<fBgd:PAB2(N^:^M8IT573WCIL0K;_2A]X^N
7L6Q(_&\4:XG#C.TJX2BKCPD.,6MH)9?Z^NCcgIO(DRS]A2d>2E?4-JLFL^H6a)H
?US^f:DWd07E3-IG7HA\:</Q&Lg=.)JfN93TQLSIU/R[<B/)0O4]]:38gP[,4bb+
,L^D50.(&YJT9H_@b-87Y]3Z(0Ld(Z5TUH&<Ig&Q:dQTJ#KI+NKNgf8PgQ2YGXPG
]+N3?b)We2?LC?7e),>PO92I;]L/ed_PFYC<9)a923_RV>12b3W_=8-Qd)Z+IWWK
MGH9(&ADDSAUD)95MK5&XK\EI2c<^CB#RJCT4>/<DA5R<N;/Z_W>d-.dg5=OeQFO
fbc;C)I^bI2_K,,O.^&M3Q,FMF<Q(46S<VZ^JBBXfT4FBN-0@>C^-_I,?@VC(WOL
]c5ZePK5;</D5.L4YI2K&Ya6-]VU]dQ<L#gCVQgI6^8NDVgN\.@QM7IS;\7?.][f
Vg3JBZfS8.g/H89OU1RL+C>KP1PQ_>W-))83H2W5W]T[4Z0KVbKOLLc4#@e@Lc5/
_Vb-b)J.B3_/.^g.L:A,_[TLZf>J.F=9&;QA50KbOB24H1c3W5)G2?8U<NP^d5W:
fR63/++:++C?IZCE.:;;+@(L(4\_)2I5NJ47J@,BMRDS7#BfdeNKH55Hb\Aee][/
cLZ]DX6/-R-R-LRMYb4RF_e8VX>D3+_AGTU7;45QCU9EeF6BcM:<LS,5+/4OM5^P
=N:L[2A-C/?Q3e(_gcOK54;K^bNOX;cUQB+6([PC_bb/JH_D,;MIXS72eeWeY4ZR
^O05cIc/4[1HAe1N>Q,,>2R:H[A__.g[g>>?GZM2VO)b)U)a+O12KCX9]2fP1[gW
GOZKV;-1R6F-:[DUgZ18G5F;W+I8UM:^?3KA,80=<.dXQ.FHe.gP+N3>+<NS,D:Z
eF>HJGG:eA4N@CY8-HRc6^PX(@f6^D^7YL[E<^5d>ROWDdOC[&V=B(E37b&E=MMf
8)E:bNIT&UAYL8;?0eU]@F:LT<572?Tg_)EW>6?C#;+bWW&_8FBd7SK)?RcMUFAb
XVd]DU.#S?/Dd;5?>D22cEbeL/N^XR4#+,503S\+>8bQ3e8+[eIP<:),O><PY>Ue
6FbN4^\g)#4ERd#-f:Zd)7b--ZVC\6^9gD(W))8PM9=Z4\egf-;QBOTbdecfL2bN
eD=IX>DHfa@[+WW9F_64U;-.a^Id2VZHdO/UF&CO7MZfVR0IZ5U(6FSBg+be:KW3
/6IWGW?HBMH?SRd</cZ4YWFYAg<8X1]D?=;KOd(4?RR3T=?_[F8B^8DC9d#5W9fb
KbL/e?Y-+QB,XXCae@6RDa.W@Va95ZWZCYUCT<(Wd@gJ/KWWY1&\)XV,R:[4Q=&I
@)<?BV]KYVNKHIJEPN4+ZA:W&[A5U,BF:VPHE-2>(@QKO4)LfgbTINSFH>fT4OK/
MdJdbVR@2I]d1cSI-&<UaGI898XACd&(;I,SY1^W#_(\ST93J>^VT-ZBA5UN84[U
DS3S.1MQPMRE/e#);[.ga1:++.O8IE]DEF1;O4<S@=]XCcA34B5WcD<g8eC&_A53
H6VO&3<Jd[8L/HG@D@)V/g=+Z>SCcBZS&1J1O^=&:4PGD\IZLbe28f0XWe-SREge
D/Y9fU7E(\SBdVPbM+34>/X^2@>d=KaPRN<0@.O<#DgD#e8P7+4WOJ)&D0HM\5)C
:dML[]X^0Z0VU_[-1/S8,-4BM=(.5&>=^DIbQ,5VX^QLAcT4T)F([[=^MM=:WfKQ
F9<?>XG,FYJIA99.+C/VUCPC4,fY[>D+MLD9[bP,TGO&AI=ge]\Vb^UAPLWUc=>B
NaYWZR/a)/5\,#;^?JfX/@+e_MKJC/8IbPYX/6?J+5.BgZL&Y.f)<EDH)UC#4I]^
a9QCD:T+R80M[:;T2A_LC<2N[/.Q+AB5L3B#GC]DgJ>]eLG(BM&8VPY6SS1:+0;C
6XD+dRKOG73R/=UL3Z;8<GfI60H5dN9,=a156aGe=Xb>bZSO&X^M+eC^JL/,_7:/
G\X3/NDZ3Sa@@X04,]fFI+F-XC#;92,Re#AH>T;;#&8;0E1#<Me0O0d1YFHE(U.A
I)Zg7#4;@-G8C&0+WWVVA7(+c/@1@WUfb_54aW;20E>;Z))YDW4+SGDT7\I0R-?/
B\daE/K[C,>(,>O/,bCXM]VO#9-.YZ\R28^2@&9/XWgE5e_A@>XSJTe:U&FDELP]
eUCC0V1eO+@2=E2[7HIgJP3R85<F&M:Z6:#)2JPO;<(X-9-TG>2]#QXWddWT[Fb@
E#1.-g#CDXgVM[Vac:A+PECHXBbEg3CF=&:E9/I-c-Z3cF#XR45P_7\<N<EbT.RI
5#9G:/2U[.=?@Sd3#[YS\Kg44Z)L)S]^)])aQ58VOL\JG4JHQV,&;E[?P3)C6N&M
S,fWHUb_9bT3M=]=2U;<6)Zg:D0BLKU>;B@QHVL0=VG//=\YH<,/UPB:c)fZXR5#
4beLE]1b9CDRJ-Y;D1M)g,]H;4,YM;16LV[gWTX#T44A6YFJM-;/DQ/)J:GD_8)6
S7,TH8IF0,UL&B/L[e5VR;^dQDU7OF/#HWYX)V_(4B=L_^_@M]5JL1JJB9YDZ[a;
;3.^O#MCLcO#\e:9cAD2>eM#T+K[8(^Zf2\ee+?@,Y/a]7\X=U^@O&KE;P7.bR1R
0DYW:Jg&]]<g1b6>VgKaO-1QS@P[Z1OHCT/.2AV.U2YI^+C6NMK/..+-cK2fcdbM
0VESfSCR@(I[Z@(5-2+@^Tg680/I0#NgRD-f&4FE\P;JLb7:@gR&W349Rf6ETD;V
[GZORea@R#,&B>gD-SI32fLR++49U;-N#KeVGgCZDI1Mc:CeaDX1[^CD^@Sf,\><
K7d5VG>gD@c7X7-^IHC5cXB(.B/eL(&4OX+NQ99YJT0^_b>X_Z:OF<C^O@];N95a
,P;JA?N#N?KW?K9Z\_0\Z&[Tgb5FgQQbA(I,KEH[2_B&UG0T+dg?0.+YOS9IDg1_
bYYdDFGWC]Z<C\M1_X+#FbIW<^\&OKe=-e@9FE<CaT,B+J#Pcc(XOL_b>STdAQI)
WJa6+OVdSWdAQcPEd:-/V/NO51dgb]PE:Q+gRZ&MX_d<VgL8\X&-V19PK<X+bS:)
4d8051&A@0#A4IGO@)Se/1EY@(,F)D0R/Qa2K^/7.GdOXA.1<.D#KRb&WAU<5cBM
c^DaNYNAWT/H5#gD>7,6L?&c:.],F>OcG3Z(Dd(P92/Hd.,)N(Z6-dfVO@EdcAe_
Y1&R9Mf1Kb^,Vc;f>79\gM_T3XID9#7P;X,28H)1AY?1M>CCDOV;&BO27(\,DT=5
2#/Z^OGB_/.Y0FZ8ZTf)cB3S-L+WN&+FME6<@cZYPCM8d0bBJ0Q_Q\D<?H3(:5[B
;E)J;9OST]+=397b3V,7^K>b7dSLRPOc_(V<Re;U@2>7@?g&dMEV>d93cV,5dW?>
X-BFGL.SW29JD9#>)>QS=@MV87M\:dKDUJ;5B=0fEB]IL>X?][UQEVVS3&G=L1BF
BCDa1UX>?9LfJ;R<8#U\d@,8J<M5.,JWSb)U&CHBb:cZ.FB.AOD;LfcET4CJ7U2^
B]/&J=AGDW@RPKf;:B(N3IDcCX[FCMII.,=#faR>6-4E+]FP7(E.9DbDB+e=BYE>
V:ad4U-Dc\H&aGf_XX95)D)87KK&81[3&UR>A8JG6<O@\12G.R-.e:P[IO&\YHRS
?K6CR/^^(P2#e=]8>@M(-KOZO::H)#aE;#b=EKNd[,<;bcc<9NULf.U+-GcT,aHb
\V/_,O8Z_e-94D)6G2D/U(WII-bJ]\:OS1)#ZH@\/@CNZ>TMGHe(7I8=<LJALJbf
Q2e>&?\NCFeRACS2&->4RSRA-[;.>V3a,d0:PVbMG@LWaLX-5D,dMSO.C6)6cKB]
@bR]8#g[/N=f8cFGR6AFW]e<0<R/^eR7(I1#G[BJX>.1>U(Db6:GZ@#8N>O7QS5I
^2.5[_Mb/WLX&5H[Cd(1F.0B.TN^:HS.L\9/WE3TGM6V^g^N<KCRXQI75(M?1@)9
B:WcVe:YEI_Y13T5SKQ&()RRKc#P\>IF77/MF#G\bPMY.E&\+RKWVbb8H/C[07?=
+28>g+8b[QS1K;H</5)ZC<9,e_W70A3_SQ:9U)68[2K-DX#;X0BMGTF5UC(f^:03
BGR@/D@,NEg\TM^aR&^O@-+@((8PBEPeWR\@^)X&d/d1]^=MgH>HAd&SC&U3gd#[
aY>]A/B9HYg(-N)HbH=d(UdR:_8+/Ge=[.\B(8TGUU:EC\=+[/?(V+__]XAdH6VK
ZO-RYb(^=_LG]]Q+,+M@?VZ\\J.#G9FP>_f;F4eC2TU.@6]ZEM^W/CJI@3<;Ie^:
R-g7,De(#]YK3gZdC7a6.M#S[G:/9b0:[E27Z0]TJd.4CWY0M/2>YDR_aLA0TQ4W
JH9:#;VA>\B^L,[EC(;;#0GJ@T,#1E<+8aL:K5fM,5g<U]b=cO6dPHKQS;N4M[OU
SD=&J3-H4:.8)dCYTN^>4gAH]bJ[VP9UV,IAEE8L1^KT5>VX+OdIRg=>?D\1X9aL
He>K0ZW#N3><b(<->F/0,&B[B-+L:e@P2Q5A_?#[d85f1CG7Q+.e[\P&V?7PV1B#
RM;1=a]1VR7CNBIL]\UK,G,03gRS8g4>/1;adSa/RR9M(VdU)P.LeNMaf\cBAcF<
O>egQ5:E5J?^TYd1,YAN6Mg-Aa/XXeK0AGU7e29HCY?=P@CB^B,31fV8aQLROU=J
_A-eM,=)#G&5IBG[f#=EcA<Xe;7D8/X=7I+HFa[c22DR[9;.?XbCD5eb]3,T<-cL
O;M=HRY:.:LAgT8VZ))YV)J/QMf4XOJNX8Df0_.9:&&CK2P,a)NRR?0CJ._EK27J
@9YX(D7XGcc=I-V7b=ca?]-PK]3IY\Y(4F?\9fEY\=A:,PHgCQK+;J8D#/g.0a86
HGNQU[Gf,BJAN2VU2UBUH5P+gQ5@8f2W=>CQV0^.&Cf_9L:;JY4=(OKZERK6(0?D
3K:F(]WRMKA&3(V2T(81W<.](MX@;P/6VYU#@<Tc1EK_EQF6;>=TQBY2Aa<C\=,1
(@1\Gc=66S-WM<R,bY_QHO?aL0Z11A4N0,R95O_:-a52I&1c/5g_Xd@\aC,V@@KX
\4/[[(][^#74AE_J09OQ2=RUI--UK&Hd6V+TER9EF9d5]PI-+.;LLJB0A>>RC#<\
:TP;LF1]&7YC]V+S>@aU\R0d[(<e=IA>b(8Z,B8)B#)@H^VZ/GAS/2(Ie8;g>Y9C
86b#g>[dgF0LZ]IN_[f/6#)I+Sc1E(8W8Z]<5M>,VRbgM)C+YQ]:3^&FPdObQQ.D
=A4aQ[0.FTC+),MO<2O9&JL@.B>=.d9LE3eRgC=#Q.a?^O?a9K=.=:E[Yb+W/b1c
2[)BFH^?1/c6(.(@[,DGDcSG3?Fgd>O^9_fNJA6BVe_IFDET8_@0T9b@Y3NKUIH1
WDCB=?&2S3a\^5#LK:a/G03-V_Q22a\/5bJ;VE;.0Y)=B)58(\6]WZM238MML8X]
8<;-bAEGaZ>[J)cGD;Y<KU[R#2(HSTf@e8X+a./],[(_JYFGN[>RUc>I5MRGB)NC
.+?DH6&O^K3L8^]BdQ]-IRLG:._A_1S)b;_WP3R.R8Y[GXRW9\a#W[^5XP<C1#BR
@D3O)MZPU387?FV@:0AdXRcc;b^Md1W>_g58,-^.;b_He>>0Z..O_9\b.:[VI)<B
BXY/LG4GN#A7XAFGN:/P70(SEBGZfeDX1P]@]#G)BTbd052ZR^9YEWaFK@5]aUUZ
aK_F:7TfdS/1c0:])QgOf>M1#(<-398/WB8gHGG<,X<;9>-X/R.Ge+=F3+X<aR:C
XSfPE<(O^,TL3A@Y2XNL1-8Ac1;8X_DKUd\0RMMM=7:Gf00<PJ<-(_=WJ9C#gg7d
_a>Q,<YTPB=_-dFQ&&[bMgI_GE>TDD50;3/d3f?W0-X-B@1[UOY7?\ed3(Qab]N;
Bf)JN1Pd3LS-&B1:dQY]]7g;S4,\42gA0OE,J19B)HC2=&OSdWPK.PE2g63(L<3^
)ZXOP^L69)D[eNM&\L&TAK5U1WP8b,-6NUeOV;UDa9W;,K=<A(_<NbE@0;O]4)ER
CRNYIa/V_J2Ef?OOE3))X#7O4G+R52bQRNU>G6GEG_ZI@,\G]bKV\bH?-NO36dKP
DaPJ[c3>302:b5Z2).=O?4R7\GcHe3M+W49Jf&-P72)aUE,dD/cLQa5[G4XW85\e
>>eHAA4V-aG4[MKdXZ2RTAJOc[^AFGB-K<QN5(OaHUa\F.J2-I\#R&F+W8)Z/\)2
Z8UCe9V0VH=A)-ZW=]Ac@8>@7QK6)Qad.Gb&/JB@gK5IRJEKF<T9HC))d9KK^&L6
b#&a&Lb/H-KO1.9d3,&#77H#LSGVR1#KRE?+)2,GK9/ZC)dRgeKa6@,<BWeZaI:Q
gR(EYeZIA1>#@MY>@W[IXdFLVOL3KKH6;>G^)U5QcIVJRJD>FZ.9.4A7YSdg=21F
0A@6_HDZbAU#a7M1OAQK+Q+56)8<FE1N1DcY2[agM^)JT:+B]4gSZCFQ_(,9VV1J
F=T8I6dcePTN,O8T^#P4_SCCWULF[f,R&O+_.,(>Y^>^=+eSK?g<>0,SM3^GTe0=
QW)[#b>:EJEUVRLfLEe<@UX/CbXHN>XH7+a@[+=J7<8ZE_&.cRU@MREA1.fEE;b\
)LM?O/DM-<-Y=RFHL//G6&8=I5c/FS<gH>g<-0,8T7&1^A^3@e=7cYgX:KK3Y//G
16QG+<,BVe\b2==(d7,DE?6:+U+:_)KJX)@^)cEaD0B/=V_R&#VLGC6SW<Y-<&P4
J8L6YA]_2RW94Q1Y^#QA[:?d8YH@ef4MU(]M\=cFTNg?\:a7(54U@QGOK;7ccc8&
>E5Z7/SQ>(8BQ@5\PWOPA7fB?JL,bTg1C#?PWO[D?4f4IF4+ZV-+P&Dbc18F^8K7
C<^(L<bB><2cF[@SBKO61T<K<V@(+VJ9HbD1F]Hg<,+f<R@/7&L9\g)B/FU>b;gL
WXF,g1HTHcUXU<Y,cULH11@#e?=9-XaYX[5FR2BcUJZS&SQfJ/HPTPP]-2f,a7Hb
\a,.0\?W@W@NV]&G6RTc2(1S-R_-01=]Pf0Q=V,6a2S3]1AbPYUIV09d[X#egO9L
Ef12SI>+BSdD\;X,7)fW;CH\+GGWLgcCC/10\DT@f8QPe@a.+2?82WUF7WI/:A,,
@/.d>JGNY>AZ=+&#0_4^HC\+HMZVVKIN86,aK0V+#<]+V)=c>I-,M;L]@aEc8[R<
([[d7O\-+/JDUK#AAK[@M2L[K(#CJ2)cIe]C(\_ZA>YI/4gM7PD@T]b6I01B/2S_
WdQbA.=]C80aBZf0ZIK>X5N#O\g3ECZb.g2544XcE9R8LQF\SN8V>4QE().8gO<4
cYRW^=b1Rc>WO,FYOA98JX&0+WP:>Cac5/GYZF0I+G()N9YLMC=U.?6<T-],;N[=
T9)T7O<(;_(R(.eHTC,;P5_CT>ZQKEOYCX74bTX@X^WIP8:Mg5dHAN5(J:EJ32PO
FPIeE<W=?8B=d6;4fW75VfPJQ:YH23EV;FD8gN3X;3N<P2@C/;AfDbe+;3UgcH]K
AH1(VJc1[;JGBfZd6.fY4P<cAU[c3e@7]Z4fR9\_+9@:Wf35,]#ULE[0^AIL,O72
;P^2LO9A7OPGbR@+>UQMGT_-eg&+5c1E^E?ZP2^_dUgTRc?K?JX:H,82S@R=])0F
H4a7MUc[X[1/XDS&N>CBNcLE#eA^d=G&#S440(68<dYA?c5(eL.CN^<(Dg>G+N-N
#]9LH4a1@-8HdR&EU:W]9+8@L3<<c_VV8YS_7D[;8L(#J_SOdV/9.ZK29e)K_[\c
WF<+NAAI2:(6R<U#5=?MER-S(EbXb7HVB)-JX[LE#&#<9ZXHKY@0a2cf>,]QSg,]
YV]2OP7;+FB_G22.AY^W6cYSC^^Q,?.U&9^X(3Af]EIb0PA1?R2)61LE>9?ZEf+>
.>JWA&Q?Ke1b(/-3<>-NXR,RZAfC\WGb?0N(7gJ<7]N6CSEeQC:&Ab)HQ]Hd-H-?
>Q4#F-[F<^@a@_6Q?E8H23=)f_N46)eTBRaO?9/Q\Pf\,)Y0gUV@N]51@1H^Qf1#
dd0OcdD\78-+:]e1.:Egg^)(4(?AQLUU^.4&2/&9-=<M6McPM>f9Ec4,Lg;c&\K:
b:1H@.aQS;&>&;#3G=^CCObJDG841+C>VCPD9@GFQ.NN^eBG5D[-S3A9]\:-:)8^
\KQ-YFV>?+2LLdN/RT;g:>AHb_E1-&<>]PX2.?+O]Fcb3=PD8<T2TO#W/YU@XS_Z
aN+_L^<(a(_^EgV,Wc[35>IHZJG[GZ3HZMPTTVCSRMKOO\b8&[>)WZ81AJ&M29W?
06]LZ1-5cK[&Sc3QL)f1cS&B.5B-I:0SMDN+aIR<#FNFS](IT)B3XeA[YFTP4R]E
c1[bc##DB_(E71dK&f8@c,]NTV4eCFT62^:Y2Bd[V/XRM:_Z0X;4JA6=e?Jc1DCM
Qb5CFGdL4=\FN]^PT11D<+<HF-74f.MU@GRJ+<#_<LMW4cKKQ:(_:C?U=3cTbFAg
;7?IFaW9b8UHEfN9PeH6J_LC,7R/XRZX),:TcU/JS453+/=,V#L@]/PC)fKBH#>4
D/bF>:QO0;.UA8=Q-c=&<_2>\DTV_=[&2C;EPLX+eGD4cc+\PeZ#MbX/43\fe-)3
1IP)]d8Kag=4QRa?98,FK+BMI8XW6gNN5^K=8OV6FFHA,WN=X-1YN;RG<(gGU;C4
cE:^-/S5Oe1DgCdHNC\P1QcS[;)EI\Ia;CXQ5ETOGbR.]:N27?V4+0A.6;0=3O(2
c_acBKJd,ULI:7#O?MJKBK>N/c=D#OQZOO<SPCf<<bU0a;T6fCB]QHK.>E.@Z.Z^
;X^B_LCFZO7;\@>^]\AEcF4L&\XC(b28_YH/c6X)--#_/0?0:D?HH?RFHWb8dD5B
@>_[6IK-S:=2[SQAX;S:I5V_A9NUQ0#Td2@]L)5H<A^D#;XO^VN(2F7SQ_>8RI7(
4Q]X7Y^Mgg41_)-e4G^0N2;#7@T<3M(LL-<?UX7_RJ_)]#]GA>NWc-?)D#OVIG;_
QfWXac]31[cVI+CWIH&3Td+PYS,B).523-I.HOE(5OM/4@,3Je55)2Q(IRa7CO6b
d^?XD?Y;U_C^b8=GV.)?@IG:fV:3a(M<Y1Z.T_[CI=:5TXN(JJO=&SfaRR#=_>=S
0<db4d=L<(c&_M2?R>ZU&^(@B(/.-E2&=[><3H)IJ9,NFYO20.#ZQbCbD2_:BIPI
K&YR7Ye572WdEPG>5b;ad9S\]7:aFM&S_Q77S)X;JX8ZX3?bCLARM-)^=JbHOf:S
63/;T0a=HN&+Q2da(R=bMAM<E_0\BbaALXWE7UNNA^Z3Te=;+<.0d9C>UFg1.-eP
X7T[G_b__,g39@DO((K+J-AS3[Gd2CPJ5@GHR7O@S8YH;[Y:AeEcaEH6>J#4SGV+
Q>>F0P/27]:=Ad0_MM6=_MY.Q(_gdTd=24c<<O/Od7,LX/A:1[8?F8J0RO<(G544
KG4S]+#&,f:9(F5,a1gG:?OM1E:E0U8fU_fYgOO?V1DC5+4X;V7ZKR\VZ<P^g/GS
@2JK4[_aXd0DcaL/FVI(7PLZd1f(RXN3:TVH@^DX_0;LIXT_5:)IJ-^M,[,\#34]
SA?.5UD73a35;UMTL7OYag.;/-B2W-M>Y#04>2&0@5&@:dTC#]\6Vf0NNa>5N?<,
Q4=PC305D<56_MZIU.]d6YMLZcdKf)YO9MM[O9OUDE+ACE948\^;U4C5C5E,X=>Q
^2QE>e=g<SZT@]T;B&>a2N)2:@]]X7>aWHI&.ZQL\R5;>&X[15&V-^Ka.<:-(S9e
EUK28ME2+25HU.H0cfR?E/>2d-Q[4M5])>)EgSK2HFcY7K3aRB#+GU>@3ebb;_T.
\/,IITGP2d=OP\N^g(8=/R=)2UWX4>6:93E3H6<RVL@<9/#WZPU6Z:agY=eWS76C
SRK3=f)_M?7g)T8a0:TGS(aM=I];6:2_HGT]2,XcN3/<R\ecBQJGIf#<Pe1NE+VK
^bY83&?JTTJ.L#3O^^+6?9&0HLXAb+4&F?QH+H/3c@eYT?[]R[XLTFFR89YbCZQ3
K2M@FcJ,9\QA/b&]Ga_5E\/?([Q3=6S&<0T+<?1?-?Xe.>T]ZIN#eXKe^GI>_7[<
,6XZJO=.Me#Z(H]ESB-U.R_Y]=OLWOA;[VA@>N7ggX42dQP01V6H)BQ,X0X>_0P+
Pf\.I&PZ4g3C3O?,][NbdM3;3>;3(Hb[gR9EH3W,D2YSKQ(TVHT/#ZZW>9/FbYV9
W6B\TT@#fG@D)&A)+K,]5=996F_RR&O[<?b/Z4/_KCfMKU)Fg,AGGdRJfSGYf2d@
U@TL\&e(T]M0FSfg;OO8=]&,&b>]#B(<9W0QRb.SJ^+1N\#<]Ma+R7,82^6;7c.R
;F>.@79-TDV>X(4Rc:;O982W5FS@M53\aT3RD-F4#79\7_UI,R,.8/4DfQ6Z&];-
U<5+W(3HDWa2M_+^f8>+U(7ZY7T?7K_4]aF)M5E40B2ZKdW60T69DGKFATVCTQQ<
XBdJ]F[B;=(0aNOZ:?g5Rg7XD-D;Z&70XF^\E:Of8O-43dKN<=?g;E:K)@5U)GI7
TB19V#4?d4LbEBP=385SLb)8T+OB6Tf9#:91f8A9[5M<05Ef9,92T(XV[C,E9ELA
[-gE@Uc6F6+.]3P,#R[T(1K3B6];-_a=[BRD<\aP9YE;(L)V@<=9;^]&/Af=DXQL
HK5[VDfR#FDI=e2SYS,e,3+(:>N6(:0M]Q#cP_;Z7UPY5-b/(bA:\YFNA\4ffB5>
.[U(^@E]O8V.IbZ;g3aWGcK\S4LQ,(7<GEb<;1Q9LZ@fMZ6deQ1-fA60S;GW6U8(
;JQ__a-fXX@+.<aAf:5QQf-@\@Y5/Ee:4(SOG#/[eaW.^^O7ALVM5.YeTSf;7EPb
fd;8)M5Sd>O94U)-(3=@Q@XPa+L_\./VF6=T\aSJUY<M1EAWgNa1#<bOWa3cO(O9
Te585A39_aBC/P/EU45.C0Mc#HcV#fDDT&U+MK-Hd)+cGB\>PK89HIf.\5/P/M?3
gI_#d<54.SUD+4^\<]S&ZgNFX9WR+4?26g.>H3gN_-V@OX.K+7X^&CD080J;TL:a
4XI/IQ0eFA0af7A.Y[J./K[A:5b0>EI6D0UfH]2&MVf\cAaA1CGb1(WXJW34c(f9
gJAR=</Z+JW-Q.?D2M-aC29_ETfM9-GZMA=8(Ve7aB>.&f&UbRJagK3N=SF_/5NC
I/>YN#XR:&\/C::G3[4/WKTC<Q\GHYLB]M0]&8MNE[c\AgIeV6L1.\<BWcG/Y4.g
f#5&H6CM[5BDV6(:NG:HCGgJg=[_+MZG&58,#08a&Q@gdW)-fZ0B\+Zf+8C3H[W#
5LMZ[77M7fdF+.E=G#Y0,LX+^M.7O>^K99\][M3fQD&P>#/=+\H\f+00.[BM@<>3
Y.ZT+b#G[8&4_8S)WAD=SXcNAZ:^.H\6]>HCOU-OPIXZZ1bg/>C63UFB3C@ZISV4
.MR=]#8>9QLQ_E)V6<RA9.V=HMVTLW=_&Z0aL4ETI8VEc5/@@=5FN_0)]P?ZfaUD
5HB,9L?M;F[<#QF65V==7<Bg,KZICaG3&&<.FCa-DRbVR0V9g3:,5S2?/F6OY3,F
(9LBG4+cX<X[1;R36U1Y37]3=Ng0+9RT&Z(O,+&^4.4/L7FDb1#VaI-F\fe2\YLF
4)K-ZDT/XC.\[:[fdRK)RF&R[^(6EPa_GU8a+5D@-D>Q6)a?O87X@7=W8##E0T.G
8aTG=c\CBdfbP(8<BK\-8Ba3gId]V#CX:O7VZf6-g?DA&FQ^&LLfFRW>=GBb1_P9
g,D990TV3?^4-_G7XYDYLCNSWHF(N)UHM4fQEV<FcINK20DK6/0KRKEO\G>Q2Zf8
^Vf[4N>cHT/NS)NDG>^dMY+egB?ZQ;95[_)=MGEcE#)16L-5B1JWX/;Q99a^;_dd
;MZWLgV3PN(\A,V#c6RLeB],+GZ1<AM(2M:67\,)_K(T6:+gW+NUMXW)6)M_S(??
Vb(Ze6MI?O2\?6=M=c3fP6T[XAA1bN9cXF7O1CO+7^=B=H>2e>8GLcS\^-3^c[C1
?cHG4#TM^])+D,E.]YM<4,E.b\7B^[@VI;/PW(YO-G3:=/@Dg]>PLec=?P(a(M],
3d1G\G+6,T)1Q?G[0E?@V?^E2Y(ag]:<39d>1R;.9e5c1\e+45bbZbUTb7H7LG#J
cNMGV(HacfO?<=L_48dE=aJOSag.J[?e@gAZQ5A;4b:8dHA,:b,LE2P1[,eL0RM:
DK(#>9I<a4V2IgXL@[.,X.g,N)RVYg?2b-4-DT5c^:T37a<MVFVJXE1f50U62b8E
NH(Z9JfP>JKY\;0>;C)>(30:^GE,5c5V49a8f3I=:;,#_(-4Y&VF5?>_1_+E<P7Y
dOEX6>KV(]_bF-)GOY4\\+YA\A4#SSP8/,9G-g=DL(U/dT,@H3(B#K(29^D9-UT(
6H?D<bDe=M2-VN;.=g4+3B;fL4SD:OK[\:&BFC&XW3]N3_6Vc&]eMV:\O1/^,ae2
[N[XbAHIgf#I]@dU#^>[Q1Eb;\:M,36&6LIE6d=Ic+J6c-VX9Q?W:9Y)6ZY+7Lef
2D38FC9WS(X+6]VR@A;1eA?IE+S<Hf#D3H29AbLPJg:(DM#C]B@)5C)QZH2cXe_^
3dXRPN-gH-O>MCf04RDA@T\@6O::5SR\<f,S32Y@(dX#/aH0bQT?0>?CBZ#aa8Ta
,E-X+BdN,I1KPB>eT(NQUg;G2@\4P^[,K5G:/Y8+0N>MR/_M\J>9RLKCMZO/U3,d
(M\&S82N>^7Z+V8>Y03;<g[F7Rd7afc4A&]P[-G2P?.<6fJQgSOS8:A/gBFOaU#@
?-?C+)bS1;5Y?6f.:=1;XGL>dM;Z^17fB(<IaV0-K>:FPR^^+#^4,MfePBD@XIeQ
<&ZaU>51TFF;+dJLa_[7W[IGd[X[I442f@Q8O(?-<I46ECad<^c:HR-BbX&EH#=B
D&;b@;RV,]6b=8_E1E1OW\)W:-##,\Ve=7b.0UESS50I0:N4aHCKHM++d2[#W[Q[
>gFg8Oa^8;>03=KK,c625L@cebNcG76R3C.;\S.8dJ#)V=YSL#LIbA0DE5E;cG6O
0AH>>-PXc@D+Xd-^]Jc81+FVfA>0UPEP3S-F<D75\ZR]^H3)/2Bd@/)5UK:@OUFa
cC?+Ic9-WI[dT(^/>@-?-_=XV]:TGT;^BBS3VLMIL<K40^]8Zb^AB9B;D5A\K]PC
9@;C,Q(]U#B(JN^_2_IX;3f5_XS:?4D[=5g@F2F(D:6Xe<_[6\YUfgIDE#T.XU+^
Re?gEY,fI=OUf(2<D(e#K]ZCcddY^YG[PRG4#:]/5[eg;\8B:fd+BI[d>>\,bHRB
-,-OL>N<)6f\LM=LSJX6TS]U5]+[]S#T&4-a\J<Aa8J9O+;_SN],_C6?D<.PXMMa
6J.=KAa?D@MU0&^Z(]<1cHZA(&8>aMEF5.GS),UMMJ1(0087G(gC)E:c5YSfC.^E
//T]8&ZCJG0K?e+(9#,:Z]V(L.>E@bE^\KU05f-^EG#EJO;,eTc[+\8,&[W(<b1H
P&&TO@0S-bC3J#bDO,ILHBK-V_]G;G:(S[W28L7=(aa\VM:V8RN[b==\]2)g[5SP
05+OTK\CgL.-gR+./6eCKP09V_;A(E&]<LA@@QZd]QQ[0WG&Xc(TReB-RVJQJ=P)
0a[b9DBY-7.?6:N:)E>-E&PMJ]Y3:aeL80):#gPdLA\Gb^A[B12Y-&7BNX>\bAc\
&f<GW>W\Nf.Qa#@#SV,:+f#SEa_H]I#P71L5#JA=VA)d_A4<MYd&g-1W(9<YJ_\P
cF.c)UD(<5H[/3Y_.6KFT)->OBA>.eAe]4H_;4=KLSTcC1CO4[(.>2QSH<=\?)gf
EO;B5?J7c<_\6F8Y.W7+JI>3<>If(W&3HAJB]WQU?fH5b_MA@MK6BC^e+9OA:?X3
\P6ZCEGAM.fS/PV/F@AOGX\f83./<27Q;2@Tf>D3W&@^\1RCT?gVL<<9_P<23YV<
/,F_U?(59T?YC/LDZ=]=5EG-TOFJ.(;4E4>ZIV.4EWKd[7TD(/f7X/03Z&(e,[@E
Z/4dUCS)6>1B.;\XTHRf)5fG-g#9A_dFD=\8#CGWe.YG,eeCG8-54.JGRRG[L0W\
U10O\+JH/]cBa32dT31EO326G_CGC+V7B4GUN,7?KH4-Ld;397fVQLJM>7=50:\H
G[A9N7_,897&;(cT27>A7W93bg;aJ,N]RB0KT+;9+#=:UgN.d#dc:A:&0B#^;1]>
SM^Y2^UYV=XcZdNG[R=EL+:T(,FF(=D\0L^b.HE[X>0ZgI0eg71O@+b#O[LR(5E)
7Ic^G:E?\L;]^:c;M<-L5=M:7^59DRW]V3GO)fRGPbV5YSC65+:_VNYT-T-7&B(,
HM(.NU)VX-T5#]ZMZPHa>&ZMG-\N.E-d@.fOB+O+gD-Z;eF0KEN&eBJZ[6F;77QH
&.Qf>(J4^<cAXL4VQg@\T/C4:E_UPI:Q3Q9I<#B(2,dgDE8@OL+J?\1MR=ADHWCf
III@H+=-eVRK-(QOJ<2e(1&BWMa3+=dM:0?c_e9,5fYa)^cYCMH9)T?@,GJJ+A[4
D:;9UK7L=?H[CZ:GT6V8V=Ee:B_TB/fR/(8e9Z?bPV1_;6C@4R4#ZdfRESY9b+&0
XM(97CN)[A@d\RM9CY0)+]52MBdg4J@2QBcJ?b[gIc=P,W4JCIB],/Z3_C7B#_GK
>GRgc=[2-);.ZZ3#=K76.?[PY_<2.TIA4IYdJB6g4@,]V:Y^J;XYE);LeFH69WPK
0(##3<a9fES8,Z:@R^X79YAH3cNE/A-7T^_cZM0[Z(<X/&]1\YOU@\M:8C6<#DaO
0g\.:5T^OJ)&[3\Eb;CS,T?:eYZX:9^^g.gb\TB&8=EJcP2L(\=Ff)(RFVIOe_.;
=;RY4LaPV-46[d?3LWI\fMRV,4A2QF_WdLaTN#@,7)fQ#5]-98U+2d9I-T1a#\=M
SNf4NFS8B03N-Vc&4^PO,5^_KCQ)4:g^.?YRGU&TK0SGNR0_IL]LTN[d5AKA2>NL
(07EFJ[>?YL<3a5e1&@S#1((cJQN?BKA0T)ZY-#FM>_Id94/N-1SVQ3P2YQXW1FY
BabFE\M1^80RTZ:KP:AX74[[,YA+0O(0.[]a8NMbSXdKAbF8.OAEf)U.bC>&&J+U
@TAeOWPZMJ(.BSGGRC:7ccT:A#ME4Ha_UFUGg>c@C_V]6dX<M_[=;/QTLSU4RC]Y
2dS::V<X78JBe^=+A=Q81PD&e)YM.0Z2<##YeE-&ZIN+ZV03)D>PW]SSffOf(4VU
2JG0]T+0>T,[]d0a\N2CD,<9/KL#YVM?4T3;S<Yg]8X>^cG\;e[#SQBLMQ&GWONV
@86\/?fD#DWYQ[8,XW695ae.YfVIKS0-D;=D_G0+G:\2&dMUAeQ\CT,A09;TM4:B
ZE)<SKV=b[Pe[XFAbbT39UF7fH=LB5#.UeZA).bBc;3Q.]<a1>XAVg7@P[4DDXX;
QgOACIb,cZgIC+C?GJ<L0(QRC3APPAJ/GF772V(144Q2B2[F0#Q9]Z@Q+?B/:G]=
OW^(-;:RM,^6+TY0RAg4NOQ1<+F8\MagIJCT<822_f579GYBT+=5<J9ZI>I4,8^U
aW&[<NG0Q1I_O+HALa9-D]JTFAEEU+9MY;@<CTJ@e5OR1_acTQM:RZEBF=(gFSY]
>4FM+DM@-N:aH;F@2.dW)fXB+1TW7cM.(^<ZNHCPR,;2_f4)OPK/V\eFcH,W]Z_5
WX\D<P7@2O=_HAC\M.XM4<3CY&O8D[J(YW9A0,@-?bR-dUK[YPP8[\;//0H4_2V2
804=XCD+N=U4eX2^DfMaT5[FK]6XH-8P-R&LCg5N+)_3<>G1RSB93dF)/b;NOI:+
D_[(5Nf5Q\#0(fLHb&/1d=LX8R2,[6Q+T2KO=6?<GWPX/@A1Z9(:MI;H3fU@eOOS
8?R0P3HP_349I@c_GNa?P&a.Z<AC,Z?GJ&V4GJfC)3BY0KE0R,Q(:T@V2cc9Ff@M
Rd?aVV,KMB:@(C+\O4#N^?Z+,P?Y@#]TU1/G0I^\/(P_cRI+K:_M9U??FR2A?=C?
(6CYN0N?<G<&c(/T)N?7V,ATK@Gg+2=YDcS.8DK=AQ@M3597IgN7TUPRR.VW27EW
A+MF]Wd8[/RRS;JZU:aV[C&@<=Y.Ng:_ga.3fB.9OUN<.ROO.<5J\(N#^XD/CA<Y
?O.f<6]<cWJ5-U/])AD=NaX&eWQ5M&b,^Te)2d_22>U@\(4R8-0&D9G2YfY<3b&9
Hb.0BNZY[M3fC.C3^QbCW<2@RZ)_O&eb2Q\72@@CL()VagS[>Ua0Y./U?eH66f8C
TECB;^OGKG@-XXdQSV7(U<,W/f/65YL+YC[E2,&O^C3e<<BeV5SG6M^gdPK.>6f?
2cc#QZ-&7\7S-]A[;CAVcFXRM&8/OL==5)((ScW-#<6aC.H3F/XGZ42^/=\e6YJW
/Pba.I&5Y97e9Z9ID^NGOVO_\@<8<O5[@7S23=-f/(V.=V0;&S5RB3>(PL67:Re.
KP<SbPFU1&bF9X,1LPfNE\^#5/[0#?JT<]AD<aYMTX9\AR-(F1D<^=@4#FO7d,&3
C#cFC,KXK;8C)0_.0<5CQDG>g)<7LF&T_0V8ae<6JLFd<M.6RAWW,F::05g2A^d/
,V+A&B7b\U6Z9\K1e[L>aMe?VY3&.e0D,ea)8A-RN3WOg9Q];c2_PCRN.XDe578(
.H<3g6YX+;2A08g>)C_Uf\,S56HJgXPG6W721ND/7D>UD-d,/BG+g3P79B_REWC:
)&G4Z(ZB_X^P[d6EV20Ba#RF><6M&@HeggfY#O@W.bSG?MWTdG:cU]3^YZYb.S#W
9Ra..=B?E4XCe)dFI00YG;@CH1cBIa+8VA.R^XY?:R@MY^E>CO_7a8YI+K[0_:Ub
3FY(J^5P<AV8F8,BZAJ3>dYKU[JM(-A1Ka8H@Ndce3S_=#&T8Da4F-^e)\c:J+eJ
9:AW?@+TCYJI&Ef+:<S4<C,M=R^/#+A[G6:#/G4a)UR<K>SJ#YJ6R&Ze>8(JJ=(K
<-QH]76CcLR09C@J(:8VJQ6U-)&)<S>@fX;)R/1<aMg@<(I>_g7Bdc)]aHLG=TWS
a5HW=+e[P-)?2PeHeTWB2KXLG[#_M->)?Aa(M0eY57E>_6KBa9^)SP/<\7K>TMA[
d.A43:QTI=f17I_)3=ZKYG,6JV?OX[OLTO75]F&#V]b&K,b+4g0gKC9BLc786QeD
Jb_=aMDbObI-)DF:;a9MQ<Mg>=#-)bMM;M#Y5^dM>B>X,Pd.DM/B/VCC1XN^K)RR
MP_][I/T?fR?c<UD<>Q,:b3;MGa66g,M>0\/6PX2;F\#-)A^d3PPLaJ\+7I8?.B7
Y=\1-bPUaGR:#dG:U.BS7)OGA+cYC.?#22(V+0R->@2\\VBACgZW:/1X(FVE0U#>
ACU(J^=bF-;-A(.H#1E1e4MCAH/GU(Z1g<BcGg=Q-Yb^F^((U:\GG&d#f&:BWCUf
).ZbZ;#-YWJgI<J8&F(QXR:3[b93BU4G8]E:UCNcd41AQd(W&ZXZ)#24?RTS:g-3
L]@>9CII6>@\a/];\RcKW[2X[-8?cKGd<;VL)HdFI9HGFdHU@N\WDd5APK]W0FH4
W)?:-(f[c.-c7L>\VP=-A8J[g#aW1b+3TA]dK5#/JDW=@B?Z;cM]?4)4[.Y#+Lce
5?4M&Z:-Ue]TTa9N<EI9/(SXCb&0T7MIABDEXVH/+.)LM35AU8^1\SCe?7B7dWa?
6)?8D[BRCd/OO_DZ3R-^0KSE#PD?,\Edd(\_:DA\/KCHZ_&?,15(J;#gG89TCV+(
:(1F+36L\1X(>6+1Of:bV@)2ZMMf^UK,)0f0ID9GC:C51V#EEDc9<R&&L-U&[VDO
JF/QT=,@J7g56-YW_,CM.aRJL1&??>>aLTI(+GOY+I>C;BCW5.7:1:f-EbQ551^:
TH2@)5U-_YVX,/B0eD]]+0#6fIE3MU6:6_fG=:UG;82eV9;eS[VfI3VP?&]2?K68
eP(GXTbP7:c&8<bFQG^Xd?62aY1,H1QaN7RG1<J)dUd?^\.^)e+TY>H>E&g6,1._
;C^<cZ5c3=XM0X=b5@E707,>Ub->feDd(cJC6>R.:@JF=L]_53R[:0IIGHF8FEfD
WXf@Q7;-VT0LV_g/\AcOV/Z5QM^VR3[\0SM#L>6;[SU?5X^)FB,EAOAJW>eC_Y&I
.V:)\L<T7g<e5&9G_D\[.WSe=ebb516#PA3Y9X533&/&SCHSIcE\J-8?9M\aPS94
,=IJ>JGE,FU:5_\XWfQCBT1IVeGg^9.5.@@>1E]bE:)dJaO&OM&71HQ,Ze)QNdZL
5X)@TTYJF=Z11C(eV&8MO1_\S.B8@WOD<]@2Sg^_fBPZ)?U@21_=f-0F:Q9@@NXd
JWMgHNeDC&^OW);eFLG9\X3\AgWe7<,b9(e]R[)cd@+P/A,GJZfV8&g9X&-IPgD0
#)WK4cb<RL#46OXX3O&AMOPJT?FgP1D>SO]a@PKF&;Rd)4-ASIdH=?J5:V(AV.4.
O=RHG/SM/&_F4@SY_E#Z?f<4g0BD&8MZ?bb_KX^\V7J]L&GD5A,77_fUQQ?.0FVD
RL5:A5Bg:1aHQID=41XIMA7A-[]UCK>MXBNJ+##A/SHaI]B?S.CD,V=W^_c-aTJL
\b&K4<W]O9MK9T^V#KY3ZU_39eV=VF:TNY=9FJ#]A?@X_Y0=JRcQ^0-JNY-EAgV>
ZQBZO07&KTH4^d27Cc6U^4-6D?3d4b58FRZSAHS[#/AR9>1cWLIebKU/ZNLXF9YD
;R1(6XZc9cNAIEP:]=0Ef?e2E(+B7=6C?Q2GI86#e4TeeANH9C##Y8151@>JEcK\
G03[R]Y))CS3>#?^1OV?3)[LdRg0dc^32^da]=K/SV:Uca5<+^(=SHR\Q@WgU\N-
(Y(JL608BG&A2TV#NYGI;c,I8)GQK_b1358<K>BSA(a3&5(RSRHRE5,Y,9/LEIfd
[D\&Od11::HNED11&8:e-LC2NCX.GaVbM;/QJ;a;a&<)4JYTa&dS:6:aAP;2RF&5
/-Kf6:Bc3]D3:RYF;,LQ,aFc22EXX?d<I,KFMP>O+64d:I9RUW44b;&=:36\^/K_
#IY^6Q#D?R9a11P&P>?aC2]4eL]6NO4;)&6RCISTI/3B@,^UE4,&e?L(d7RZ8FF7
LOe;\LUWSU6:#?AOg?@bGW3:P.@F_VO>,b]38ae\LMJ]d6+;68d,e6geKA8-.<(Z
Tc+F+VbQL=^bS:;MIfOF\BVeB[FD(9e43b+M\X90;_cB/>ODBY5HMO\#4)>cR/X(
]aJ6(8C?H]:9GD;W=^\)bO0JB8@+87R-\1g&5#KTGgHH1F3^>BVd=e8B7aP<@_?L
>++3dcJ5;7;9GF@gOI?,ZISF]M>CN5[RD^)TdAFUHcN,B0AXeJbB&>GVDZ]P:]B)
_d;JMeIEP1C^:@BTEgX>1;+0Q(>]0+Y8,-S&A5?)TTE,S[J/V-\9.;d1cb3KC)VW
/]AeQDHG;P^/&OadcGJV-XcD;A84@\3GB.YB63<DQR1]QV_LGTU\K^@QY#6^;Yff
_JGE7HaFb>8Id[(8?Kd5926N;U1TY4.B3],dE)f#PN2RHL0XY002SRQ=f2^&<5-J
WC-B5(O&]fW1KW)a=f?^HFa,=#4V2g>\F\/WeH;-<,]8G=70I,&DJF,_)(8I)2cZ
DHKBBdLd7JAP#6A=RcW&G^()FO?BIW<AHTa0(HQY[+Vc;a:;A(XE6__O^LC[X]G=
7]LbY#TH6a\\C[F-fI;cRZb)0FPVC^1WRVL5+_75?N^WX8L3+D>&aBM99=CV;+ZD
-=NE)29L@_:eB_d=c?I+)gR9<#)PN]O-9.>E2ZD=1I^]6(C-_Q(@&B05Y4NSIY<c
JLX73Y..R4H4bTdV?(Ic0_T0(,cH,gIK+WgGa3L-YZ>7QJCP66OXG_RGJYWZS4dV
dICI3JfDI39b0U1dZ6DFW#\;]e\M-^VFR,fXb9D95Y#QPgaB_8+>+VW43HTRYC_,
-D3OI#]/V8V;/8MOgKcA)QDGaWe>W:W/:?7Q:,B0\0c:2(GS^XBeATWefW40][J,
5=R4aDKKP7#f;e<aI(Gd5JY7GZ67,(Y7CB8&@G@-38OU5LK32aS&3a:-\eKNX@8M
1/8c5VI>72:[a,Z5OL^]2\#J-9M(KC_EVd0/Y(@[-9#9RGR2\P0H5e=D(Z4LK,LI
X\D_\<da-NF/WH=]-X+ENdDc3)),OZ&R,=&Z?4WPGU]V.AQgFMCeHJ3VC8^P^7f5
D1b3bETC=LH;Z?=PX.1AO,I>^HYHBH^E<JM:/0,YKR2X--HH+1L?3QgN/I4g[V\4
KD0)HP&&2[?U?/aAKa?FgTU76-N6F+\=2?b:DR([?2-^U9W+\>fd:U2c1(UI(?#d
/FZ9[2NEdf^2W8.J28_D6;@A6@&QYccCbHO6Nb>G[.5;4TIdX2U7JE2-,e:OB+<^
cc?VT?V)W;KZQW9;[8V1JO&::]b)9>c>6HN[3/\.5(^U8#LT0FH=;LMBR-(&=^MY
C?009+Uf>B)bBLG\?4&OM/dT8(Z,7YEWHA0Y7V85,-)a90TZ66P,;gDX9=F.=TG9
R\+7^aR7=,Oe<[^T_)>eD\AaY\8ZN,E+)31QRH,R-<_C=cb_d4[GJ&ON5U9PQe^_
H?9\O-L^B3LEe8C]CJ?R\C[K73Q#LGJ=Z06(cSNf+1_B;b1>RRDZ>92O^/fCNAD]
GRKg:Ec:dCAPCg)+cIH/C,UJe:7_e:+C6Eb>a-_SL:TUTG2NbANS8?bdD3d-W@]B
>^(a7JJLNb<O#+//.90]Ag-UD7\]BceP-U@d++BW,gS^(C/0F#e9R19b8=CG&BCM
L3AeJWfX\6d;dBI5:T6_4&NY7.PCHA[F4(_Oa4eOe43XY\;@.f_Wc2]O^/NA:A/e
63U&Q7=4Jd5S3=4&8BQ=ZW\Jc(75KgVH6=5PW3MN(O5-#7_=a/PXTXFeJ2dB:&#8
6fbf(#^FRYOL,(P6O_L[_8O67MX-F4LT_=6SR;(=NHEC+;f<PGMeb4=V\bU;]&ST
BEH,+LZ/4(HQ)NROJ(E,B7=6fJZDc#1EI(7RG:=OA8B,a5VZ&&KdMP5D5Y2FY+14
;,NTPL8(7#JI7R_7H9R7L6]?]?Z?.RH4E.GL_Rb>EZUNc.Ie6]cZYfd3a2K,RRRX
g/#(egK&f?(E]KY8[]&fcPS]N2F@FO8>AF174IWeTZe9^dV=&7RdIA=5g[6TCA)b
OSGY&D5dW7B^7^VeZ/7KD7YbfVM_0S&E@/HFBWB1P,?]ROVd(/W&Pg>c;?#Z[09,
03B/<JE:&bB/BBB?[da5I7E&JA;Z(?>6EPe\N^.\U>IKW.[\C?@g5(Y;)EFeV/[;
(L:a@N>L60[8-D6@OVH1SDH6:K#H8]/1YLC#GGC;W=ga].4d6>/_313AF^.C89=G
P;aRN6ag15Se?_9.^9;gQ75WY6RW03.AH8L67G.aEg=MS.G,,MOE22Y_/(CMJ@[/
T_2/PeGPH+9g0RX+_06N686BKM3b5c0e?[AU=(^.2;Kg>A_?M>eccO-QYRPbR,Rb
?N:A4D?1FdfQ_d19ad/,A<AD=&^4?0g5P@DWZI-5)MAH3/gcYdSXb.EGLANW0ZZf
.II[M?89-0<4,AAW@QK=5B:I/7\N:df(CRdHE0e-(D+fJ;E[W]7e,B^PH#_6\L)a
]1cARV4;gec2WQ+&-N@.:RYR^PTVL^L?-X8FAbd/^[WS\1EBWBD&dBLZWXZaXDAA
NHP++W&Y#e.+H8#=B;\@]6@>]U((LBCQPRNb37HDE+]+M_GZ8W5eZGEO#Cg+/B#I
Ga_U>S^)X??U)FKK8).YT[C>Ff5GgUKaeAH,C.^KQBgA^bDK3JLD5\PU8b_]#TIe
56D(7\QKgf6U2ddP<0A=W4OaZ8LfCJ84Z/NE7A]/d)N8/=O\2P,#QgCKe_GbBI64
4/2^NG_EUA?UX&3a>a/5gcG^d>6PR_PFDH2W\R:)COIVLJN@fdR/YM_[1.<17ADE
_WX>Tf0I>)S7WT1cg<+6_Q[-KZ8?ZdJH]Q+D#[GRO@)#bfcH_M@-.Pd)Oe46.>V)
O<&<M]MPc8IWbZ3I+I]G#c.-&9@]=WKX-Rf-OGY99d1&Z)^WI1eC6\[H\1BeeSU,
[Z7WVYf-ZTW4>@/?ee.XQBL)+8dS?JE^g(4YADGRS<@6Ag:L#ZV?.>P46U3)&+.A
U3M+QJ/G)G3F#V55[)@[f[0de7fb?KE6EfbR[52fU4@@,F7AZB-MBOKeLEJ[X.R]
L9PPRW6N/>D/UeU(-bO=@dCWDWI;T8P5c/W)8dJb_Dc>Jf[XL:X(\6:aC[&.QGFW
fHKNc[[1M0dA;ULR^3]AKMHdPHF.9[G-+^A.Y@<SBMFc@Z0VZbc3KN&MTcW/7:RC
7M/.aLQH-E_XUb<S-;e.VP?=4K&W_^T0).&JMR/X30V4OY>;GAf_Q5JO?V:1O&)A
6+=T3OaCe4bL<>5[>ODQM[><5/_9.3SUT-b?eP:17@=M]YMY>bWXF],e?b/U@36A
YB>L^)Tfe=U\9][]T>\TJc=CWaXeB/b4TJ1/\7WbKX8R7a_&,1,&9=4RS8BdE9XX
#O8JWWTJ&-B9(e51(5I(&>[<;-&/eY<>be4;d1H[0,0YD1C@3.P,>Uc?PA+/gaMU
PbY81c>T].c,Y&[?aQCZ0IDQN\2&T_?SZST6:<J]>&e1@Z/5<CJ82;EK94-QgDW0
c_^B<V<J8X<Be+).RCLd=.K0R.V(BIYbN2M#=\=b(OJV)IAT<NE@=I5&TC7D.MLM
J^&]gKdMO,6YJP)c&G+V87JJSX8GMb3@Y\S;OE_J\W-LQO9&>g8H8a,8JOTC<>JH
e9[S:DL6#(JF5,a&WCK>88FS,D8Ld=HU2&Og)U4OOAceMDWR1EWUJ1W6gV7#)>aV
NVB/[N]7<?58P9[TC3.9E=-,6[^Qb-VgC>Z<7Qd]6GW(aG0;Y/#;A)1a2.JFYY)X
Z^SIQO)J:2L])fZ]MQH;dCVA\0f<<48V^I<fZL[&GIFYHYPT@IQfUa,[-dUbD>(X
6+@+V0gb])U1S@FIQ(Wf:Z]E>H8;G]W).If85FHJX&2?[)D,;Z[WJ)e;OIH6BM<8
]+6LK)J\23IK-a3E,f7:a5)9OZ^#=+R?TFgQ=c-Z5DT04+Z;6bW:)0-<aEIQH<[Y
eN<cI-a^AIe&P@<1gU/Mc)FH@&aN,CK1^gY0)/UX>&#E=gcR6>+8C_P8[A[g]WVf
a6?D3FWHaI@DWWKD2,[f^I)>UXYG@f,eW+K31TYVcZ7<e9gX;W5^K2FB@/@)3>\.
N.MBX&XaJ,_I[:f=c@WaN^cg7-R:HF(-D_(=\3)/GH1H?E\4,SOX=&MRKaQW96TX
bO?4Uf^J&@80(SZ;?&&7)Yc-8;[D#N5fE#NKCHTdWV]aGJ-DAFeMN&Qg;MYP5_^R
,HK3/?BJd-WJ9(=FbN,Cf:3Ze+0#NYBZeB1d>7CYdHY+)LN)_F<YW_c85BSZ0]UM
^&:;ScHE@g_9RN^ZX8V][J641bgE(ILEH&01A)OGQ2d4DZOb\@>.?B#0-0I\M_-:
ZL+eIQ@DF-PWgC,I)A2^].H4@;1=[GR+[/.F]FE?RRS-(4\QYA1\8:f<?N982Z6N
W4[LHJF1Q7Da\bcRV(Vf(7BFbU2f3Nf8gS;/1^AbL:\(OOL4I]N,BR2+?4Z<RM1Z
8[:d02d&(E4cW/_YE6PQd&H4-V1A4.),1H&8C5JfTY5cYKDL&J@Eg\,gC9;INW>K
LU.(.7#_Y-;H<S?-+2.5)AB1eG6VV\4?gINRC.B+R.f=d931))b(_7Q0)9Nd^eZ0
R+P\e>X.>7.+d.=[+>\(1,+9&VLcQ[PD#BaXA;f@134fDV1g1+1X@N9O&A4ZEVZ2
9VA&PU_Y+,<15OF254-AHK@W1ZJbXP18:M7[&;fZ=62Te]UaP:PMTf6aO5#X\Q)-
[aUMaE#V\F)/cVMb.MDdO5M77ReR9ZDA-a[A52DRG/(9C&:G3dePWVJ&WP=bWag_
g+P>MbEQ3bEPc6XK>.KK+B74.;9SG?:UC<I>#/4L+FET>1N0EH1O4LP34/&OLSX1
Q88YTIPB[_;@^QQ3U;#M[Re&=#+b=<U+QHB9_&1bf>0g64POTKM0UCM?N\&AT8M(
0QS9^Dc-W+ULd1)W78T[4aPA?ZJdUT9+5I(;8Nc->I+ab(=KcD(UDUASOg==WeA>
R(NdW5HY_UBBR(PH1;SX,^0gJ8D;E,OU3@HW8MA4<f>.=MZWDIQ<Y[^_=00O,AP:
=N08#144BQ6Hcg,_0aUBY54F5GUe(A8WNGV2QGZVW/_L31/:;)G2Jf<7=5Oe__TJ
?WJ)2=HCVT\+-T\K9Z]ERbT^Qc#3J@_WZ92L-GS-N4Y_X-OCOG\EF98/C@V1D:<e
MFcH-0Gg+1+KE;c#Z#(^QBSUV^-EP5FC&C0AQ48@dC93+)GAT=Vf,>HZ?_)1PU&/
eAI_,J2I/P<B8f+WO.P?7LJ3-]2^dK/5W?8aD8YSEd/QHQgMP^eYWWUNO4F=/=2c
JZM<16P)UULUI6DVD?D@_LRNRNUSGFKEZb+b@c_I8/K&&D:3?B/,D(M&#.9JU:7K
Y,b0:7fG=f2(DE4_+gW:(81X?3EE]f@bf<eD>Ug#B=.AD\7H/c/Ub=YVK;0aTa8)
K^33;d-<(eM:S#)PH236X4,0ZVOFEHDF^d#@SQ#F>\/?0ARg2MFQfcW[YEN3;f5O
e82H_)WYB4,T-B(O/.&#J&]bE>VDF+=LC^V[=Ube#Ie^ZU65g,.]<(+C)9K#@X-@
[&P20=DO4I=)Z:(<)Ce?g-O/AO;G&?SJKP;BM>H<;B]1])9eI\_<H,7:DKYCg,JG
X_F<NV.G^=H\&]>-._8gc6A7@De9Y.@E?e:BI>=J?bL_8Na?,?Bb,eCc;J^SH?gQ
EP,7<9?Ia.Y6[OG<)(X?cZ3P.b48ZEQcg@FZKfAC_M/DT_4+L;Eg)(U9J<#;9_-&
X+d#JV93)(<b.C5]T#2Q1^Z5VUNd5?RS:20JQF)_>09@[Ng56WBaYF)SKLO=Ng#N
VJJ5VcZ[=19(c(L<N]K3DG)N;^LCK7PP,b6BRQREa[TXOUg4^B,3bD+P)g00O^e7
d;/Q555BdD)ZXY1P);L_GGUWMPJ:2\cH8L=0#L3;O-<.XEK>/7_OE&5+bLQ7YPVS
aS>BFW2>_63[3@Q#AHXZ-c7I-?M@JQH6MJO(55^XXK3VA#S^Kf0C7]#9L:dVN^P^
1I]T77=TZ]d<b6bJJ_^a^=O<4K0_/(_;RL\\=BfPC]:H.2E0cZfN)?D<OU4Vc6__
(U>)#bPIM:4JeW<>cE->&TWX6g+2<<I@@O[a3d.34^8XKZ)g6>WT4@[9Y8d2F]Kg
\0=X)PG(A[&OGSee?fd92TMM&1)F(R4D[bFc4#Y<7&[0eW#RS,EESH-USH-^&LO=
?=bW)a[2RONCCJ;bM@28O44DVGTCa,3dZ,,]M)A\.M8^d2N=d(KdcB2>SXRfA]cR
/Mba&b5QOT4V@g;TGT+>E=e#]eU4#PBGT63\02=T0,R0bS2G61XbYNgHIXeOU\.9
cQ<-f-N+_e@.bJK-MM6)cUM;5e[D<[BZ=+B6\4MUW5c(079@/[g;M&3N<:(SS636
gL#2?X;),bD/D/bRBfVHUZES52_]/+M^_R>P0\LV3aEdSPfG\V?GWZ2&>=FAU^,J
FE80#?fQ2(Bd)L:V^CHbQBHBZ,1.6^<?d\(3V<10:Zb-[;RNLNQ8Q/.]_8R,@U:=
OHgIQSMDN_].#M=I,UYcEMX,&A5W/f6/T;D_LA00cK<N+ZKHQPLLN<@OC<Aa&<<>
U\<aDWR?KW[IN49QFD7=d;],TO:14&DY.79:>2;_4&&fb0eX#4UB7d--GZOLTaON
NZgA2d3+@<&G4;2EAR\_IRgC\T]R8,;29R+eaF\c,<7eW;^_N6LI6B[S1,,.J+0F
4<[G9V&FYB0M&N_5Y_H,KY4b^f2EEHI:JNdWUR(1=#a(J_4fZ(^fBV^S2A?a:^E^
+90MA6^G);Q]<(4;SIRf+OI6G_g=+B3TTcA_E6dKB]2P(c&S=]24PRE56e3>^-.0
97Yd^=)WQ/WgH:3,0WR[1L@=Ze;Ha,,V0BfeBeH40V3dJG#-/>.?RgHQHQ5-bU>:
H7AT0bFOW>fc9/^JYLU#A[,?6cN)5\..=4=Y0fB01.2WJgAHCE>B+CbCddK&U.Re
+(JA5/\8/IB.8cALN^C39JgP:J2L@1<gNc/[0gV__EP=#AMEQaP(3=EeH_N=3B2M
2L(c>]2[5RM,Z5LBCI-5&Jb5f-6FCI7937?UFFFfD/.g9g;3N\)Jf2UC((c@YW3;
dF<_eaIVI6RHEH(E?22_bgJQ,QWMe.2KGHECa;5<<f6NJ6&8Z)K]I1B5MYSU?MP7
OLLa6c.M[)W64e1PZ/T.UAU1V;T3gNZ+@_4a;PA6dF&?#(cU=TG/E<G)S7K0:QM<
MYF5_?\g=fd;c06XWI44T,TRa2N,->6)bS:L7\Y#Nca=dSfQ;E(<f/:OLQR;CV;T
B/]3B6g-:DW+6Y3G[f#1>5CC/28]MdN>OT02deRYT/gRWQ:Y/8ZMeaSb0R)_b,[K
>1-0QAXf)SWB,(aB.a.;S<G<WBFQFJDT5H,ed2;3Pb?ME7[]&=3e5HOg[MRRWT=5
82.58Yg8a.BBWX4bJ]Ea2WY5:-8Z(V(Zd838S3]f/DC>/dNG?L8UGT(B;NJ7<W<C
R<(,=Bg/5P:YVf41)[T_(B?0X<HZ@fc@T45H50C1(:V=<F2G+\E^.1@?c4G>=)=9
;7,F_74RZ;:>>SaEf4/2;UJ/:K,S<TS\\g:]@]e#8Se;_I?JI7ed:-E3fZ(,TW)Q
O,\^=Ng]\N8&J-]dC(10Fb9RCR]EGWGG9_ZNVL#b/G^,fR44M+_KIF@#8Hf,ZgE8
&9S4WA2#;dRNNQNIVF2NF:GJHa)RId;0gQ8K,d-b.gbS@OA#]G^M+5]:R38+N,>X
3>c.H;=6EId(=Uf3IS?F[#(-Y-)V+Rc19\TB]HcN8PM;CafAb<=356K?ge2:;VQ8
N:D1]bWO^C5IeAeA4;,5@TcdT)4P5].WPQW^#\L2aP,;DJ/SC.UVIMHB77@>?U7[
-dS;FT@FQ127<8DPeEC28P+g?V<2DCTH^g5A;&RQ<>/A2E.J),;V#4N09DD?RL:+
d@bJQPfUb7B<f2R?S0.&()SSGOd(9WVKAG]#L#0L)3G#R)+YN97+#1(CV.F:+8&2
M:OWBI&5BSgD8R+>K;2W0.Ke>[eCBA@UK\fJ?_37-T2MZa6CS0F<SQG\/aXfPX:O
><J.VAX\,.&L1<g\b0Od>P,5;K7J_U/9O@Y<@QC9A46I3f]VGY)T^AR/(F)>[=Kf
\PQKUO#MI8I>K1-YFR-c?aPNM<Y:N3F:VeOJ</-aa^HH:#N#W:/W/[3JB]5dJcAI
>\g^VgX:BWC7bU^RaR^86&..XPb/TGT+WJ[(MYK.K)HD)Ze(_HV[,ZQX,A1]+U[a
f->b6XG5f,H##/2O_8?EL4@c<4<63ZWOb7/e5c@KUTXE,UU<SC=98Gd/GbdQP/7K
YQ3Y^&0c+>OE&+9=_]GN#GISPR-?gJ0]G&A\GMEVY<(c2fG7D4SKeM8P+SE0WMY7
9bVZMJQ.]Ze<egSX6a]A>(JD+3e:9Za?\)BbgVC+X0^00)9f8dgC(7U7-c?^26NW
FBa^B)6QcaG;W:^;PcPHC=.Hg]TW(VQH=8e64JXLEcE;QQ=T79PU_JDK7C878]/[
3J@\>XYEKeTXS2:J<?\A9=R)OJc3)UF[dKB)GYbYec+)KL^ZQS90\TN>#8+HgUQ^
e7QAQ115DMbIE[9+J)7T+<gIFP##?Z<J:KIJ)\f]R_TegF^QeLH-S>MK1IVEfF\E
_T#=Ca-)VNHNZV=]3b]51=;7_I-]^[Z_a1P:MQUR:;4JY-BEX8eLE((]L16MfOO-
RV.VL#8ID>KUS\CTac,aN4ObAH9?6.K\Q@IN1/=;[0,19KJV#4g:]c;DFHZ,Q2Y>
I\+R[QF?fY&G_d:>SOZ+5M4,M=VH/=Q=N#f59c]B>ENgSQ.3aUA_+b<9cG,Mg;@P
&GC3>eaMd96DEe(3.GFZA-)0#K^_EJW_MFBa/E(AR#//f/T2:KJWffUC@M(VVC#G
:M,DE\KBgJT4g3^K@d[<X8+SYR7P\H,Ig-Q(:dY-)A^>/,][2UaD>#c=]N,YdT:a
<;Q7\2<9)Q]\LP^6#^3[[-8]e\/,D;8=W2:LgQI2/OdT61B.T3C]/#FUXc^M<X4Q
cgRcD8)AO&,0=(/L/IOW[a:JWReLLN2=>+c)Zd>]VBcBF:Z(eC86aD_>(\e(SNZP
cW[MdW)DRDWSUTeP&T@#.78DgBMMLSXa?UQK^,MD#MT-/c^MYd[DfYJc<Q@E_Q>T
,O29_51C>)TK?Q?e7cO@A\BTD@6Q[8\,/CbZEPS:,60?VI<SRFgOWD^-7WCA^-US
)82V2T<LIFC__903E9ES^H4C4MMg7,GG91/.8Ygb+AC^OFMc5gQaW-;\V8LYKa9g
S-fX?8]#P4&3^3?JIeZ1N62:<P[XG;Ff9;>KPO9=3PC>4Ad1,^03\0K.1SNb(TT:
e/AgeE_VPQ4_O,K,KHTD,Y(OcKc\Y<EZ<@5Lc#5B^N:A#?53C](EIX[.#F_I@dSV
L[ccZb-<))(_.UOOe0g+5#0B,aG=8[g^1(:E33&+8]2@gT6G=<44P5d<?N3bHa[^
)EPZdbb?2=\)NHBa#)30O&0a@PEIV9[dA1@JV)f89Nb_<<L91KH7f(JG_DLSRNXa
;Q)WN?&5RccZL4WBGU+EHcX(M3DWA7BK\&P5A5-0XO68G]DSBP>(U&W)@d)-N_YF
V045A>^/B=?O]L+F<f_,UY.7WEN2K5N(Y>b^II[XI;@Z.=;=eAT__)@:KTOBU-,S
WQHeaW[MeY;H]E08TdZE7X/@ES2\dBeY;8?Ke;KF5_#=4H7E[gg;E42@N@GKQCS[
I>78b8TPV[[@6:I-_TO5LV]3YcF.Ue+ag5HBL[V@]WG=/^S.806R#((5YdM6dD75
QaO8;MI)e7P050VH),&-1&I<fB_a^/9/faK:gMEI(69E(Q(B(<\gHQ0SQ04,dTG0
?6g1W7:4@YTS?Ja)1FP#R;B/U3&;<I(3+@dMdTUG&1F+FQMG]F\AMKgS9DDYeT2G
RKL+1;48T_0eT]B=bR+R=K+RZO@9G(5FDV,P)D&<PQ3T#CY8e:EVM/X,KUL\^a<9
IPdVAS/J0A+,bDaIWF)7U^KLD>R(O\c^6:]HZ8FHf2ERg&&0=OC6D/d#e<BC]/2)
LP?bgZ?#6dM)a:WC)(8X:NeDDU@[C@UF#N6&.B.LVF&=aLD:R1.>^ZFO6R-98g](
E<edd+f/\37,Cdd<QNMCHG:ZXXY,aBI9OfNMQ3@:Q;NOcG?bWRCIV&d=ME.NLJZZ
I\f_0@S>/#ESPO1OR;E7^M3N8^,NT=GU&VP03]SAHRO#:QNLb>#8H#O)UG;O,U_0
-E=@5T+=)Y5Y-)0b),/@R_]JWJU<gCd#[deJ..^g^D]7\OD=X1a6B0J:]WZLfC_#
5,;6&G5MJPB>6&Qa(/#DZCI&Nab4-.B1EI.Lg0L.4-8ODcAXHa8b)R:8Ue>SN1W?
=\AUX,4g24BGJc0T8VBdWD-<(d(?,E4G+Mf--A19,Z>,DYf9MNG.FDB9HIX]6]6=
;J[8&V@PSH06MB:-&_)LDQ3PP;YZC9?5eff;V]dLBAT+:eeX&6M2=MP+BaL0feUG
P.4D?AgF;Xf6_(;@-BL5T7_9Mf3d?WNJXBIOc8T2@eIYQdARAX,73cR/T,:gLLf#
)JfIP4.T,Cc]Sc/>J&Q-eaIO>&H0XT,\>FWEE+MOT1#D;24/g(gYU+a0SA4DQ,F5
Y>VQY#>T9QC)./)IGY3[&=a-4HK&ObL=54Xf<SV>36bS6#:@)VW=M3ag/Y^]BMM&
(4#T[JVV7M6K+&7fN@I\->(16MQ0.\-M<L&[S)#f-=L:\IC>(-fFK,[W/TQU.CbM
XXUCZI(b.+a[@=(_A6L9+_GC(+519Z-XO5gfg/+f(=4IY3g,I7@164ebJaB29V>2
d6X=XBXM?3&g1^<_KZN9Q@68L7>B.+0B9N4:=;SV8>,SPNa\]OQPObfa^_7H5_H,
[W(KP_41R()70\@VKW<H4;g/1/5IX^MO_2WL[OJ(LS4,7C=QZ/WLA>.J\4AOIXD1
/=L&1)^R^.T5gE#7GZ=3&I)7@^[ALUG-(764\+O+0GU?gW8Ka4[)+PVHB#a-@K&L
c;_M(]L(cd1R8?N9719B\1]JRad@.<2R<Uc9AK37/L]K?f:M;5_c9R=8cVD3>a;X
aK68+=(198+^4\O^3S=eE[6gX97^^Y:F@1QCb@^;.?CD]U9^BRK=U:Z7)cO?AXTA
/SI[\60#Td/b7e?FCU^ZVHbJXf,_HF]a9>)XDXTe+WU5?cA7W\GZJ#KJQ<?]_4.8
PYe5R.YN>A?cF8E/R.9(Y+6/(aDN#ENTaZCKXS_];-Q?Qb-Jb(SFIH0E=SWe7)55
dT_Y>JEK3@.U0(<B5T6fc/HF.(0WL>3+_a)2]FFSW-7bOK[g_[Z5\0<6-KB()E#7
2.IU1V0,WNUS>fY1e96=dAdVM6@+U-5-Ze52bKQC3C9#^=X+KHA8BV=XV8W4/8<&
HRaM\a5V#E)5g5GB-b0;O/]@J9;9K32\#1692fgcPMA/_]:SX-8/fD]X^LFNC6<(
L&]7#Q1D,&F4a0YD7DfTYGefB[6gB+1&aHKR)c,O5A.P7Od)\_A#=&FX#WTDP9g-
2SIMaY<UA0@8SVLa6?YC^1#7@<gZg6&-7WD?[U0/E2AFIDNSF4XM52IM[+_RWb#c
C_^b9EW?g<]NgFPf9CTL]23b<2KH@db(BMM?ZW>H6S(PGF3dSR)K<g46WI,\;.cU
/I=&7c]EH45\S2V&?<CU.TB/X9^[IHbSZ,cbR/P:MD740(E/XXCPZ@LJT27>P3I/
fR)ZNPB6\gGKb6VdBR+4DDBRS?NGSB:ZKF81UFV^eAA79&AK.#J);VVQ5/T2e08:
QX2TM#R]@L2^28-204<+V@^^/e\[N#@#RQ8d5D7)dL;U7W)8CYC8<c2O2O#CI^gA
R+Se.V:S+_P1?G7+;7K94?+bcUJAS&@YDQ^8E5LNeQDUD26;&12Hb^QV@\L>1E^(
C:FEAG:=_B_I+Y^ZM)g(:U(E>3O>HS-(H3\YD&EUVM588f,Qe;FC2R-OcF2NT)]a
1I6\IQ=[=7fT+>b84VdI@2_##QM&=K1WX63O.PO91GH2f+LC?/\H;5ON\JY>+a=-
[A/<PXJZgZYXQefdVGM@>F.1?>NSf.5Q-=(G1.G[#4,D:M2JU8G.1KOIS^>R5/OD
[Ma/94<MTG@^YKcY=gH?7Q7<);JH8O;?aQQeJ[YZ8\0,CKPF<RUa4>7Z3bERHg4#
XS.?JE]1Z8/<QDV(8PH+;_7-N,dHF#T-dcXaMO<F+(0#\Dg51T7=2c[C[Sf4&^[#
:X1@=;;74NCHKRBG/@>?8M,CAda&F#FKZ(L31ZH/0aDBI_WZ36N)YCCb;dM5-8^I
(J/AUD_#2:H-V4-F4O3BC(a>//=,51GH40R2^g(be?fYO14\G<=MHP;gDU7>Y&fX
NN,)gEE,9a?BdDCCQa)U)._P2&[b-&NWd#E@^f)7VLTaWC5#2JKZX:;VU8FDS439
ZCCV,T[P;KcdLUCfGf?&@.aABAQZ)L41d-?DddeSET=a&M_&5&EWP/gB2X0<I@fS
RQ9A;IC+;8dCGRXHG,OQ)FTS/JA]O+7_/?dCaaKIU0R6R4JKZP>)=KI<+;#4L<.I
O+ZW21Za[=28S+/]<O@Z]8H1]=g]a6]:c1]T86HeT1_,[T>210O,0;851UcYNX[_
#L_Q1/D+];&&cdY+IFCeZ+8?a:Z.<<&E[_KT-/IZ7B)D,6AQ1aZ-B:[-EQI&BdWe
<7@D5HRb(A&D1<>_=<F;1&J[GKVR(GS1<S^1.;8c8D\7)MA2\4H,9:\+45)G@cDC
(H8,=X/=9TP:LXeQH?V[Y\S0KaP1g5U+J076a8THA\P[ZH#?LL0=B(Pa^8dHOgaT
;)]1&5).B^MILf#J/;2#]QV<QY.:F1deFSJJTM34QAHZC/Tf^37\7DfAX6M[:F/]
]?QW)8cb^KWR\;.>/X.@3]SR&fC8XN9H@?P;QJ\#[^2:+5OK5^]+XU/1]N9#9N8g
F;/G7b:PI0Lcc&H:\@,NBf865P1>_d,Qa34OOc@M_Y2Q2,=&6Q;@bg&KK55(#Y.3
Q6:?\f=1WIBT475=P0BM_:;3(0KIT=gBXMJKBgfV-_33.5U^[M8IZda<56_\3Wd<
498.a\U)GWSI,1GBL2fJ.F?RB7gRVGJRZW#:&P]b4K79E1Lb@#FXL:PL-)QR26,[
(/5A[_]81A_#\RF,;gPF[DP&N\O#:=JEOI/b&e2AI5G2d&cY9UD-bPe>BVS#&ZV5
YGI6V]R4X&+\b=@](OPJC]f5FWTVaG(&5+?(e:dRU2IS55V[KAB5AN&.WTJVY:EW
I9A,YSbT67DG9G4O)&PSBb/aSVKJ#0N.4.RfKE9=E4C?-;Td^gaSYZ0Y15Ag6C\[
HIPbVfJN)M#e:cBfABa,Bd01Y7GO/X8b(??7L38DAZ[BQ;Id_fLZYf<YfffbT#)P
?V5Pd0dEZKOM:=J<=U3<DYIBD]7C95Z<d)Z+3&cS,25bUH6V3R@?SVL/D&(gKA#O
BI[^8L3H4NN7B)bRR=Ld#05>Nf1RPG__3g\DSP?N5L7PDZW7^O+1=BS@JfA4dEg6
#EIIa\fbH@e1(^8(WF>@9G];d:9]<<Me3X6KI\=@JW4+I-GGe7VL22,f=e<AdQaN
BM+(\4P(c/^>0Y:_AZY&)58g3GT#@fWF[.DfdQaLQ^4X7b(I,7TXe]:A,T<QC@UW
ZDWc>38IKQGH6YD+J9c&[9YdTE__R9D&]cZ<1;#32:,=ARH]/C(&N/7A3H93<;2;
-.<DO07<S:321[QL)3EcCHPc=aAWJdb=[5Y[H]L3^A2J^TQ]fH:A?L+>;MW:#LC4
#T@F_@:=3\6P-4?aca?\gK6CBbe5SD_.\NB76F/-d#UC_+cETc:VIg4W/88##JOF
HfP?,O@MOBY.fYY7=QdX5QgTIQYL0.-F4LPYa>+H\KXKKN;Y93a___cSD9E&IaI2
CHf35dHLF,G?QS@@ULU<Ffb6&=8L@[eNWE#QgaL/117@L.7Of)5M:fd.[)S&)_TG
GWKGX&B(MUaaM>V7a+__S17SXUY?A/Y7>bYR.;BYfV>gJ]96Y=G0eC1DOUeEOQ3]
O3)GJY@93B#LP6Ne+ZI<DLV1K8[GX5Ta=>F3c8VdW52]X0]Z?)b\?_URgV:;#]OE
FTGVDN@V&&W21V4V?eE=GEGAUa&#:6-(A6TB\0TdVH2^EMgfC@W:LDL5d/&;>ZdA
22S;c:GRR6L1JLFEbJ-b,[IE/#4GFYUZMWBS3f(d1adF(7dL?E.D#c+/=^R^=C-[
C=^3H9?.TD@:@4V(0::=^c0PWO;5K,RY((ZXT<,E>@8Y[M_](V(/CR\B_MD00Y]F
>&Xd8N:<&b@)-b=B:>bZDZf,b.U/)AMT(>d5CLG?60J/MH[#Q_Q-EL6=J?ccH@27
XJ39PL^P0RR:Pc_41aM.&Iee<R=fQKa/L5LHLBdHV-&#<5E<RE:LNR^Ee@aU5dSC
aW:8A0bZ)K=P:AFOWX#B4FL\TN&U8QPfCJY8,Lf(d6ePHFGWB^S+S3/d\Vd)Y13)
4)D)B,)7d8^+K2:.b0LRK&8GfE8GK3W1aM,:-E>,\0K],6N41XPQ8]Mf+Z/L@T=L
]X(?AFe0]ER&?HcFb7-9b@OM4MadIFXN:A2gOT6,8#[QA;d,&_X4:fA)J]E@@+(P
J8CBPC1@&WL;1W</T1F>M#JG/I,Q::=JMXP]\W^2]TA46cSCLH0FM8K5JELd9PY.
RA&HRM.G:D5NVC3^cOG<:0HY(;\c4O[K80P_62,b^LA=(5W>W:+X50YC\F&ZGU2_
;YE6FQd(C[]D(#_M6HP.Z;9U1D252+QcG9HXd?B#Sf00d]Q5:\#:gWC3gNK-CMaV
BJ.6S6[O5:dd&+M#^+Yf@NC14<:<#A>3S5])Q+\C._dd7QW^.?2?GgbT[a_XT;U&
^d4M,E5=JEb=8DVY32V]G<S[T-aH432:W[?Db^X5=F+Z=HNH^gVRIU&Fg7&[>e<V
SQf.14b4MZV3YG9dUNA):f/7BZ1-ASS4f>:ROLWbR:T_1OcS-INQc=c61B30#1?A
VNQ:P-JM<=^C(Y<Jb1>Y1^Q1cf&0#?bN]<H+L[MZWY0V;;_E<D<-DP?,BHP8ZY@5
+?Z)&=0R]T3/J]T>40CPW)-06?J[X&?[:@ZNY0=^WKV)_U=FMVILBN>326AV=Ud[
?&M+XNK9OYWF&T\#^c>Bb1_0f0W7S[3,Pb#Ye]NO_,N07_B@([\CX49,G.?YK4Af
)?KbJfGC;&eWY0(+<9.-\/NXB)2cR4g]W_=TUC@>&P\O=C@4H&14F?4<+>,#ZAP6
CB+PEL.\G?bD=_.GO41]R)GMPZM;gQ91#N2\/;N[/Q@+c?]QD^FS3^\+c9\58gdL
F[G?KE;86^E<ba.PM6WR6L5=Td,\O0G)c-8NB8DaM?TKVWUdMEaYFBU+^=>OdLd]
SESQaKWa.T2[>BdN(2ZE3QQ=J9W8BRSQ\5dG(HPUYGfI)\(U11EVBF^Db.De?X<>
I42^<]OCCd\?+?[]^V]fTG)TLAYZ0bMT0Z7O@BLU=18<@TN\VL,HF.EZU#2+e<:4
F_^ZCK68O8e^6EM0OV3_+H8,ZY^M9]2R.M:f78;2T0=M2>6D-HN^&;XRWBTHLM,-
d18,;f?<D_9QHff/e[OINd))U1ZWP>4_a=a]-@TT;=&I16DB+c8>81D-A[E<fP77
Gd5Q:IF;KP;>g2f>TWO\X.e@>OM1DHUP<JC:.AY+K_VcM;@fd,=D.1X/?IKKf2&1
d,D?VBT=[<N@Ve<Dg<eTaW0?MC(/(e1^V2-,_7fa^d9bE.@#2WIH?XDaMI,W>0)0
STAS\<VVF24BMS]WG]^CZbG0TAcTd\-REM4UO#;Y](CK@,&EYVG63cX[G2_KV)?+
He\;9(@ZE]M3)eUYZO[)J.+>@PI:a#_eVa:28Q=AWR-;,@OV_Z_eH1RE7RJ0]c@G
e0>5IM279@;VYHaI3/XO9B<7VeY]D,\Jg[\K7T[#d)IH3.fVU;O2\,:RE=b/A5gN
(E(W:N9)ZQ.79>QX:T.]I/KMTQN>,e/JYPTM@e[<F2@<S;.F\PaY<8QP[\Y&(^=,
]5P2^E6,b4e2@Q933V_Oe&DX1U/>6]PMad7R<F4G]9f^@#BV6[ZB&UfRJG(>PA04
[F>d[ZecHE\2WOSPb+JF\\@.4VbBKeOBcdHCXYFD?50.1eGZWH[K^EJ2I.^aNU.:
ZM8dH-Ng[eJJMATf(d1)YD?(D#O+JS/Ua==RK?5(O(&g,EA&->fQWO/T7U8E=S::
X1bgS,2S#K83,I]JRF?BAPE+IF&RM79KKMeHX=WB&fPDc[+?b2=T#XWTG8H6KU0Z
:SBaU#H(W8ZNX54cJZIB-<0XZ-\UF-,\V1A=@8J:;S-UCT3>Y^W)3EYXDG+N@Z:W
/e5SNMa[b0BJIC,V9[FRE\Q.>RYX9[#6dGU6<=ARe+V9SgK\G2Nf9^P1c^+J_ccg
TA[4Hc&/fF05ORf&HF@NF=WV;FN)d^_D@7>DB,KO?1B@a::-D2/&eDa>N-12MJFd
Lg:PBbX[8XO99E,G]ad&NO.(093gW/P>?TWa56K12^:,U9D_]EfU3R)A[\Wc[TM/
[3Ag13P1;eN@aYc+5cTZ(^8_CZ@3()TO=OMJeX4#baMG4F;=ZHM)#10_Gc2b4baH
EW?/#?SAd^\:,TSXgR\c00UP8d/WA9DCg?6B1V49,HP@G@QFU[U61^.+5PWZ?2\X
-Q1BQ^gI(K?C]P1ea#KFgHLFRI)\YOgJ2U\3fO0N:d0KR0ASXV_=Z^M:Tf>MH[H)
EZf[,\?/AR.7G>B=]+]JJSId,^KWP?1?23^eQ\ZC&cN(QGDEHG0LUbDKM.F^<=SW
WY05=PCFHB84H/C41L^CU\UR&85JDI+.3P;49;K&aQQ>&W#-]SeRX-a(a3<Z(bNO
bY64MCTE1^W1RgeJCDaBO4[L:\f?_PK7F.&Q+U>76<eaDX8-Ua@b-8PaeOEfVSKP
H/#.T713LFe-2bEdS;^Fbb.3VGR:Q^62f5>]<d+76,Gf.+KK5?B&O^I59JDGG]bG
)?U@Q(Fa#W>J[U&7O)+Cb4T[:Ha+HVUd2Je\@6A=eFbG)VW[7FK[4E:6O_Wb\f(>
4B77AbF:R05W5HSZ#cfTQ0+WN3)U&=JZ2GX+1]N8-[3e<EbL3]PO6[Y5S23Fc&TY
MC=]8fg>@<0JRHJ7RWdT9^5F71>aAY+E:@<PCF3HBBX8.Qg,&LV[fb75J,[L9I_Y
29?gV[-J8Y<dNbe)d8;@^McU1ZbNc.EaZ@9LQ@G.<TKa_@/2G6_bX.PLA\b8[#AJ
<DESWW/E(&1,4gc6gV^&706V_-?2:Q7XDJN/PWH#OeGCYAc=<<O6,+\0IJH17d6S
[E#.d.+N3;?&EA:</,K6cUGD97BVQ?Q]:YTP?>I))c;7dS+A46SY&WCXaATXNJAG
MLf2,fOX5H-]aWAaEO\SZ#8Q?\b/N,1@P6S3?BH,FbLa_-4WdF@S.IBd^^36<1:W
.b/dBdD;D0?-^R<fcDH+VaTM]ME3H&GAd(e),#>UHBA(JEQ4J10,(+Kb4/C5ObfF
AG>0<^.KM\10Vab@[fDdb^1OYF51a8I4T<H=/+5P2MS2#\LQ3IDVeM8(81^@P8Ke
G)B/@A;^W.#R&a03=4I)TID:V]?8T+FgBfVSAB>G=C^]EEM23cd0+8^GY\DfAfXR
6VL\=1H5I<,)1IPG5;B^948F8=7I9/I,e-QAf<c>X^=NGOJ&5][da.+>8N(:HS7b
.6Mf]LObW=baY/81B0UJd<P3VDeC\&e6GL,FNaNKb9N8ZEe.F<5W_8\a5Sf#=1FQ
=R?=FH=bCC,XHH/=I+^8(Q_MA\7-^AN[RbW\:L/+S7AI1f.TF--RG(0^]0[E_F4E
26E^16F@OFQ&O#>a+45<1G=E?:^ZbZgaOAPO319I4DOEg<08f?N>S=]4/[&+Z5(9
_#1=EH;3->3=OPJET<ZfCY8??#_>GbU.)F?1/H-\CF:NR/BIIDX5U;;:H-K=T8HA
ZHJV<6B8WDe-Y&9C(Z:3CF_\4^05U+(E3dS&?)2\S]:0\(fN:g7&(TEIe_R,b1NT
L+gKRO39b<VV.3IE02]I8@UJ,>N#b<<,ZGDeDK-^H>T.-M@I8T;-VC8/acREELZ^
(6R?O-QUP4?Eb]0PF\^66=Q;?GX=]N-RG3PU5UbL2N9eI)=DScS7(?f]8KSYZI/W
G?@0Q#.0fKaJJ/6&>Y5=@I?C\SE]ML7dKDDZ4OgFe#=9/[[dE:9,N8.=E0?Y_#aH
N3bAD#3AWW+I#L7HTWGDZ[A9PAEU78<G<(G3HC]:2SK:+VQ<&Rff#>[AU.UGaNH[
5?&(R;fQ</^3BU9#+c).Zb8,#:,8Ba5ABBP);HGZE&gZFG4gF4L^99IFddH8,dMc
AC:AG(+]\dBX-O0#W0PKIf_YMH2d7?[NRS75RI7Dd4LCDaJNU8YF(2=SR=6)d,\R
JJ8.&f<3X[6bFV\e.g^e5CJ0b.CdODG_TXeK58;DR]825-Yc)37?g/2WVIg;D>Q(
2OfGPV2A/NPH,>#\&.50>0.[1CS.#0^Ig(^^-^>F&A&->D0DYU,XC;#.Rb8X3K57
-^QN8I,FTYYMSc:NWbHM^@<Ag8Q3[N)1J:\X@+)+gfBWd6K,KKTH)UTJMGbV(OJ-
):30->7d@CWM2+WfJ;PJGfQf#Q>S4J:DaUQF1O)OP?=UZfbDgB5R)Z\Bb@YS<+bW
a6<-=OCa:O3NeS]CP?]gWfHCI?C_18DQ(B(E(8>U\U<_3;?:a1cf3W_2DeSf>;A-
2A/VSL-+JL+;8K#c6BRNMEF2>FN74?eN[a4N5fRY5@B8;L(7?CUb03F2BH]<(6IA
BPg[92&?:UOY\(f;<0G^3/f7]SD6FE-@cG)9UPRR0E)(Y[0S[f&5B\PWg0OQ21BZ
#;@+A8V5S[9ZF3&UI(Ig5XANf@7a+]b,0#BC2Xe3370OQVX\7?X@d8+M+E)>[NcP
8?V448-<ZIag,)?X4-C3]ED#4\=L8S02S6b/PbD=e[M[,=0;A8-FL/4,G=8(c>Y[
K][75Gg]1)dT:+H//N7SE#H8&P4UT4X-8YWZ+VC+MFce4Zg;ELIAeKHE,><I+(Yg
Fb5X.6QU<X<A9SX==\_gVSW-I8)7&FS7PT=a.?f3]d^99O06D[(#8fD]47WOI]4?
P@e7e[\We;H6cc;4J\0U+;S7&\8V>6>FE6(Y??0.9+7B(cU6#C4,&SRdSB>[H=19
_B(D5AB_UZaF-T2Q#(a4LQUfPXN/T1a<fC;\WAZ2(BW#V9I7G+7;1M?C\D=G?0g#
JAGEbZ@H_g79T[dL/F+a7T;J7C>cB9U(R@+B7;:F-X&Sf.SN:SIP.TG(4?fB:1TG
c>+.;].MML=&9JAG<<AN15]=gPT+I/=[B;T#OKJ&<7)GWQ?P[22#LSVG<P[X#c#J
@a<&745LW6XC8(6fO94dOSGR6THFWcM7dBC?>SQ.QA@0:;?,VYU76,&\@\+[L<V4
.EWI4Hd&EL,fKRE\BOW8PcD(F\L;1a5+E2VD7^0/7G;@:JTf=>KTb8<A\Q8gQLOD
>C1DG?S&NOE7gU5&-<];WF^La[;dU0CVH3?_c?K)LMS[L_&IYb0df64WLFb&LPR9
XM,,@ZfM(\+\#T@OL317L)R@-B2d&3a2?e^K71fg=.-YU3.\>N72;97L[FNRB16c
f9(d7=K@GI[<F1599FTELAcQX3YDf(4,=H>)TT)6)8gEKd:a)2:E=O4=5=Ma-RZe
?(-6>Af]RY+d(,bZ>aJWNNaBZ>?6B5T?P9g/RFC\^^6HE<+;57>>ULR0LYKWM37J
Q5]Va>KT)Mc3M?eI6a@V5F63ZV)V8a9>g-(>dW+dg83eF1CeL;2/9[L-ZEUKA8O^
D#4+fPK@YD6FUd#?0_XZ2RKAEP\Ie3>PX8<L#R/5(;4Kc7U/1J7J0TJV#U8A8\?J
C\@]D=>#[US#R5S+.<DJ_DFNS#Y\>Sa.W;cJ.Df[[_7X-I1.Na7a8(UAB.g#N#dI
Y5WfPQDI34]5Z)C?3@ffVME<2=7IR-2-\5<&\9gV?P]BeYT&DI6fSJEK\d/5Kg&.
X5)&TgW_5=ROCf0?6<.)]&Ge#IF\FB3B5N7RCg]38VG7@Y,X,#<TBcTc\:L@\gfH
g;gbL2&PRT>UPfQT0\4MEX,(_P-J#1eCIJ+0;=cMc>UM=2>ARb,,Paa)#DGe4_9\
\#9M6>2\X?/;54gAH/O@bfM3e^:R:&T)A2X3Cf#)8C^ZL,WLLF45L8/[N#?<D)1e
)e5ECQLRg&8M2EV&f0I8D-CZ+G7>M:IgA7Ng&SKC2-L-.)f<3G#&R0Z=eRFg]AFd
SbE+CQdKQ.1V_NeT.3cY^[E14C1)ADK-_T(.9IK;6CII;)\?#CdL5^(29R[OaY+(
P&0d95M5>NOdEHG9N#@3]_)G3+=BbeK4L(IQJN>HUB,Y[b?D-[YDBFDZQZ\b&,[/
O?I7P<#/5B2dSeTQK=JE7\Se(Wf8>HIeRGfK<K>H:[g&Y3.-N>d;>d=VD/.E7@D=
3V;S36)L18L@12U7I_&O&/,VUY5@JIeg_b+QE?HT_\>T8+.9XTH0GV\UIO(BLM4&
VYSRM:/=3R3C:4(_>K[XRf0(:EX6CM;PcA;D-X?FbUL/8f/WEe?VX-4d<Q>?_5G3
:aff-8,8574UK2DaJ-4KR1WS^W-UC/fNOC+7:KTF(f?gN\e6W(J]G31&3.Y;^4dB
,H6\8C:U.BM(U,IL2][TKaeN=/O94S;\,7=^SRQ_=AgF6^;N,N:K>\M9bMgAP9-3
G>@VM+)E/G86B6MX+)bUeHZ[KGaTf^W^^Ea7[7JfY<?^^.:V;?>(]0C3_AW=PG2f
a\(.BVHI@K]E[\:GP0KPcgPUcXAMT,2D1G(\;g)ENf2/3aV4)e]MH;[d^[0:3]@[
?0-.(6_7DMeQYT=8<?NgYXJ>HN9W>GXg95,5G<gJEfcICUQ[0a2#OYB+FN7>=K4B
WM6^RR/:K14\(WGN6G2Z28;PU1aOPY3M#WWJfG8>42Sf8<.KO2;-J7b>_7I>6e30
cV2/aNVX42ICfNU\&_g;:1^_Z#1JEd07_N9^LJ,R0S=56/J,096-8A1K2]A))L9X
da-TC,EU(/BQCRF&Z-9D))2IUV7]f\A2.2N<7/e>P>YCb<bd(-Ee:DY<@0EGCK\T
XUYA>&Q_E5&F[f=(LZF2\G.Z(fA]2ZKL7^#eG6YY_/C0=dLeO]UER1]&#HDcX#J+
B,C,3^&R8b4UOGb9RUE#UgYG6<YG2d?Bc]B(IG+>ggHC3?D;@L&)ScDA8;C=W2_3
AO;=9dOHMT4+cGN5eY<WC&U[V75HROFJ9.?)/H_&L2NcFW\9K(#YGR?^Y;AYZT>N
7VIcIZ@GP0T>CUJB6MO1.)8=-Bg)a^0I6ZS:GV19P4LC2S#b3_XQ]dWEFa?NKL\5
@<&+M)UUNc</5cZb4;1[0fH5)3UeaZF?:FDc6X+9&X]W7:PY<]S^2M=DMOU:-9(Y
C..[[&3&CM/]^,aGCM[7^_4B?&8;^_)E92]:Da\CMIQ4Z^?4Q9UD3@Jb#6aC^T\E
cB]^<-(aF-1BgF34;^G#\d;<;VN7FbFC976gT4OMO(?fTVX<6W@D<gE##<.Sg#L9
\9<X./bBJZBgF])W,W9)7@5X)H0086>5S2O/UB.(RL6ZR@R[&fO?UD;>5;DW2Wf3
0KA12E^>3&g(_05Qfe]K,Q1\(FV.]:&35.a+/E4F=ENLB)H4DNT>).91cK:B(9Ud
SUZeUZ-NI=G.I,O33E>4U2P^WOMVR)ESD&HBZK5+]K#F>TT+)5OVZ>b,ZaH1fJQM
^225]&XSZNcBWINZ&NLcOU,3S1)5G]R0@.]=#C:gc=0-d]?<dR=R5eU)2P(2^df3
8TUR?;9aK#&2M<aT@C[aV^.N38,QUO<QI6N65/NT;S3-YAFfAbDT@IQPggW;2IHS
XV?)L+PdI6NAF8P3_WdW_c+H^37\b=;,C2J)?)g]IMd&bc#_-8D)OBDcALUQ8a<#
5_<6S_YZZ;T6;RLJCU;4IL8fdLE:MQ_G?K/6X=-.9]D8,65d9TT93L[34b:.U::?
?G/b=M)[FR>bb?]aNN7\M8:<^5XT<EPVT#QE?X#(8]Qc>4]+<#LO:;T)@7Pg>?#-
[,LG,UH)JE-OaK&YP/E\>E^#IeJ.?PI+,EM^CY((1749a,.,9ICOEN>0]ZXf^E1<
<ZKfG3;E69XU,]FgfJ-=/,c)?6<VA::Ugbc_aM5b(,PB@;NG2W<^NVM];PG>/HaQ
g\BFD[A#BA;^&<QKbBXA,7_OfX6gRACK.A7V=OAW\+#SPU4\836]5\/TUb&\6D#,
Xd?#G-T[?gD8B,2P74g-P):bEEPBF_2&R15C^(Ag#SCa/3>[1S+gD?Y[Q;VQ0D>\
T9]C#]R48A:#J]X[N(YaN54^T1MAS9aI1G)JOb95C7I4?/-e8H6g1-#G2YR=\V>g
:9_6G>N_/^W,FVBP<CZ)BM^J]MX>R9e>)[HTedB[.cdKI<.PSJ=[gg45PXcT@C._
[H##OF\/(2(=+TdNfQPQYS@IcW[J0[E.@QDa)>E03:Uf8E;:HBV8,?:18#E[=H@J
XMB1IXQgZe(T\DHW6BY^.8eN&2eM@?28eEH.YW;R;#=-NB>&7^^A8^,8]\c]1OH\
.AH,)ZX=L0FVNN=YT51BQ&3@D8-[4?-2(2E[:YZ?>N/\g7,YXa?8#c=8M-1Je7L3
V^Gf_A2W3V@JF8,8fddMHEQFOEH270C6HG.#3C&-LddbG2>#TDe98L&(SB-JY+1D
GFKOLPdK[&692;DO(d&]b@SAE/fbKI#.>;-aPYZ@PabbXIg\CZeZYF1g>a&>g4-S
P6^JXc-.U/9O=M@\S5X@29BG3;;>,f&T,864EOCD#O9_.A?aX_7A9BZ[(LBXQIC[
-U6Hf(-V695J.Q,WPP7\c)#MM+UE3HG83HX2_Ee>A]>gVN[;fe:KW=Qg+NQPQ+WU
Q-O0VDDI?:TP&++b8)OZ)D,3;G9Z9Y#VHLFJ29OF;8OFSI\F4+P06aB@g+3cN:6.
Z)@?MLD+QLAG24_.]IVL[YV75]#/]bJL#?SC?FfK<9PY&=J9Ya^66LI=V5N]++dW
==+U)(O-H:I\Q6AXeMQSVANPR49I;C9-OW3L?47EMJ7<N^W)A/LWDA(0>+/<]cc3
HP?OfZAD^Y#F.8C?[_Lge?SBP;[^4JV#GQAd=^PNS?aOYJ]G)/X=VA4dV2]>G=I-
4:c5ICDf;W;)H[PN\CW0d6FR:eX]1.83eC;\WK6TN?6]7?;K#->W]Q8XHN]ea@8d
4QPI\.&bPPV;E/<#S_81aN?]QO;VEXF0cMe_]JQEV]8d8W8M#X2JVD@.9N+&g#@+
T@)>_?^2#FSffdR6BIU@<##5LBg/;13?Ud.\C,;[IJ36K.HCY-.AS2B(a@X/S:&Y
6AB>=S9T>_D8\=-bP^6S^M^>E(eN?[Y[I/>C?,QM:&9g#387T81JSRUWOB9fY(+.
VO0a-E_B(_B2,3PY4D@5eLKU:U9\>9@ABLfV)VYZ>aa.M1+eb(&&X0R5GS&E/Pf-
K4L?/cP7\:FEUW@1E9S8gcB9Q8ZdL5IVY97He>X0(U,;a2^O6-:aV,\MB@-E^#+_
],-?Ca[^4.70>;@E<<L?M/(3[6Z-HLHR+K1d3A30U4cE-VB8@JIVTP=IQ>0<Sd11
UUA[0Q5.:?28cA?4CHbAFe+cS7AFV]A,)KV1AbDHIGeb_7LCE.fE)dSbYUd0f][S
.=)KZ??fF,&WTO(L_0MROYPbGMYERc@E9,4P0?Q@[>E-@CcGPGW8@6^5&]QJI<bD
0\Cg@ad9QY/CRKP2J70\&PPa0dHCe;?=[e_.<:a#C?S_X:T2N90d;DY7@2VRFLLG
f#OBfObaG=P02RZ,J+=^#SDIP:I^e^@;]QA/+?b8V9QfC8+Ga]9aN2HRYf>c_FT(
6gXZaI8>70>Z#IQ^E?_&19-af1>@d=39WO;VcRg6KgcS_L3)0W+Re,<c^=D6@&[f
HY&5K3>/D>X9G+^E>eO@+OLRa_9[0-6/],bdW_#A:2>,#W/LNBTYYJ]G&^V8.,PM
RA,IFF;J^9.\-^W37cK8UfWK)D?()=g)],aXc)XUJ]Hfc0Nb/=&UP\TT&&\91WOP
ZD.X2KJe@.3_b6bJc-[BPdbAO(/+QF]V8<=)&(5PE[FUK&=]Eb]NaW07W?+)-9)A
ZgM_J2_<Tf?RH\V)U?AP5?A6/aU;CV9M--O(?W5K\[+\@O4-0cX:NeSHgb<C.R^6
JKK&()K17-dWdJDVO4:f2]HF8.;-4--ZWRfEZVWH)(]T[8XP+fY49B63f?ge(YUM
@X-=]\5cCG]/0g+PYEAb-0UWNF2V9UgI:^J3)MI1&;5,H_4gg<1d1e<NUDM\<3\<
U&1\#/g35I3N:E8a<3fM55C[JT9YMG.EZ1Q\ER0BT5ILc)MDK.XaY=Y^+)EE_+d#
6I]/9BRUWLZ/RE>LVcf426<KgAHbX,X1PIPUKd4RWGDaCd7ZOC_YN_Ka0aKYdT@g
E.(GM9#MF2^-_S_:-6:=,4B:7HdWe5KC04XH.IKYBcS<DZT=ZO]1Y)[K.,b\g3OL
9,gWT7M:?<=<;?9gUWe>0BB:Lg4DS]9Z1c@U=bVZ736\NTN,8-#W4=c=W2QdeNRa
U2NF77G9UN34(RV30(JGagA#C[H:N-/(\RA[9S]e2F>bfV)bId0d#PK9QF[Ca1)<
-d)^[eE=VY6.?WBfHaPQ9eL]NLKAa32.c9Q=DXRBHQdH>(P-(3=(bWYW[e6N9TVI
E_P9,eW/agGR(N,>aJ3::aN=\CQ84X-K;Dd_2L=FNDfY)d\?d1bAS/Y=MY]P1/]&
4.;;0V87_S,W8UH/.XL.F++,:[Y4WLd_.\f>9^,01PTcS>^3Xg)]OER7]F9?=dMB
eT8Q,@CQ@D7c3^DQ=/DgCbPSRL6>WA2_G]d8adFa-Xdf]O?9aHMc5c#<M(g936g=
5DS9U7_ST\HVW(ESTI;;6K<a;37+H#M&HN7-D[TN.:TBYgTc?<1K],[UAW/3_FO+
DGVC55&,4<[QH#KfRW)GH>T=P<V]Z-A8?WE+GdTV(2f@\8T;/d(cT].[[@?Vf>:M
F,JLP-Y6.a]gL;O)B],-SHWZF?2f_AS]KA;DA)?8P[)]e@D_IaGTJ_R<XOJQP(_W
\5:SG,eKZNgKANHZ6-Z,M<8.XTO,:+GNH)5dH.VS-2[)d[L1TH2CJ_7BbTUZA.05
YIgM:;TRYF5O8AcK3:3H^HfeM#M:MIX8532X#.+_;g]QfZ<DcUZEYU(R8E#T\3/4
JBD5Q;#?/@fbY58FAdBW3KDQ95^,?YB:5?1\\UHM^+g:[[=++\(,fR2C-(B3).7a
V9?[B]:@UeO[GV+U?af:Q^=J<X=:/5Z8I82.c#S9?cLe14,JUSeIYaZ/Q6J#_0CC
]d8)A<?7D@8IR;8_@3b6TUM2OJ\D6LCVR&fUf5DUKF7(VIDPU,L805N9L+:)?W79
GP(>GIV,>?RNUefV/(>,,.R1^<V\OA7CA/=&;TF20]aS0>Z&Gc&T)/P;RQL>BW-D
+\#JOEG#;52JDc<0CU\,?#KCSHHMN=+\C3g:ZCF5(^R?.g4&7.1Y5TF]R#\,4a,5
K7&[]de6K[RQ2:dL5_91LX6Q1[HW?P<?1U2Ia2Rd10MF=f2)3aTD5]H/M28M]Qb:
TW?]OBGU&df#QYD/)NQN(6AGe7cI:REM>KL@L.f3cQW7gZ0_>&eCPZ-52]+FM>8G
g<VS07B,]f5=U_WES_Vf0VR2&-]fJBa2CF]\7T5>R/aR0f^N<f1?9P5&_g-WNMRN
Fa9_.\fA1NPTaT_HS,g#[_#K7==F:7PI^P@fRGfU]_2H-PVNJ;[Yd<2-GgK/2XDC
,b:M,Vb/AL8Qa,ObdC.Ye.6/Q4GbA]AIU+VAfVW@^;-=CS.[CR>Z&Lc^\cB^=P.d
P12;[JB_5Y-P2;a6IaJ1@N/(Sd^D\QGV_8#Y8)UZIX#&1UgE[J=^(A:f+07?[68/
@8[QI\e[QM=EeG780:YW/[_#Z,BVE;Q7Y^GA74?15#+[cMQeH#CXLW89VPR5;.&)
A[9\YZ0[-bW^P6Be@K)dB6SNb=KT3dZVXF,.1OKN-b[5U[If#SQ#SO(TDLMf-I6<
2CU-8?R1Fc(BGb@,DO1^GfH-1I1fFSF/R<Uc0YC:\.+:Ac>;:DQ9MC<aM1(48]e:
bGW5AY.D;#QMH[;O\fcdQO]+Sc.1-E.?95N2&(d\;dg@0M12a]0;aVR<G]Da[WR4
D)M5]OIW@JCQeCbS</EdBV5gfD?T,))cN5ZdR,e.+P?JA(Q=H_OXaCX-)RP)6&H]
98EI2)UN]5ed/((QWOVVgQZ:LTL/Ng@gd+4f=d83E-A2#O-A2+B#SgQI@g8BIP.=
2eYgK;EP8PbJ)6CW,([+B,cDKHA4IMe_QcGQ3TP/OaK/(,9IFKeV;.?-BKg-)LCI
?GQaV3F7Pf6)(CP,J5?JeTWVPB.cRa\c<-N361M&/CcSfb&W1IZKCFQS&HD5K47C
Q7]MP6&Q(<RB0#bFJ,8bTU/->^UP#b43CG^+f/Od5AUHWYZ@HI?[2E@Z]VKUMB5\
-V(@KgJa5c.4B?-OS/c^G3R73X^PUP6Pb_0[#?cR&PcGG<HFV+JfGM_f<g<D4<E8
5YF#Ng-PL+cX_93<8=-(e-a;^9ZP<1/A?OFOgL=<OPL^:B:f&[MH\MZF(R0gP_F@
Q=CaE5F>afBK6WX30&VL@A[0(gSdP:RbW9Te?1&Tf]:TfAX,A2]><G8:EJG9/=B&
a&LM,MA936:ZGAc2M\Q9L1K;U([55d=@QH&^1:_P:(@<_BDW-,CYHQ<M^Hd1e+7W
I764L+]<(FfB]R1T6.9]QJ,SdW<S/B8Pb]eW3B3Qf=<+LV>\_Y.T(gM&eJ34V,bK
7^/SH@a8@:Gda#SHXcd#0,I?CB1BE&M-[UA=\<6TR4HW3&1KUJD0XD;JM)X55EAa
T;R&51g=_V/.//a88W2KWU\TOCKZN4B+Q\>dS<#&B2FC7W)3GH8>BQgP8^VDT[R_
/PY?G]X>MJSeP\.[)4bcbQO/Lf)B;A[?4f(W(\V#c^Y[cDC&S\@]b1QRH,O8R[AX
(HB^=+,/SP=^Ca>@]]+VM,?+@&4.VG#bSYaZ_@V<P;A3g]7PPD(],G(,XK(OF.#b
(]1B[P:4\(/NG3<KX&Mdc:]([4;6;[R>((N#68EdB^59)g+LO6.1/-cf/L)SCC[1
@b80B-d;(9&d@/QcFO[U&J/[XO:F+Z&ZH75Zfe\c-V,+-2@5dU/AOTE#Q2UbPPV]
8C08dRSg^E<WM36JcU]71e#,Y^]O.OBebO3+17__H1/U2>WMB/7+&g2^MMW749IY
U:=g[81b@CT@8C[M\C--7ePd51[dB3e^:Q9/EKXWT2a&BWWCE\3Q7K)DZbIWQI)<
8OFE/C39X,JeG4+EYA5HM\.KKWD&SR(VJI<#Wa@RG4O=7Y/&;Zac\c&MNSBPRGPK
@BI&X2eCP=)e/7QPc[9=c]WOR2>Z^HbZ#+NLWVbbbF)/;-H7N/C#9-49&eeBM20,
M:D-fIaWUg/R11fH8@Mc_954A5+YOd_F/R2A\AO@&X,W?[OMf=\;4WWQZ?^:be8A
dS6d<2G_9NMVb4c5\(?#:A5[^E3X.Hg4^094\(6a./4\SGN2[WTPP5,K3\I,LCO8
SZ)^C=_eNVLLEF51#QVW>P/6?NE93F/aZP<\.B&C,-#dYMO.?2XSH6OAJ5/6[f3C
YP)BM3H:^#P.KMZ.K:STL@V=7M#+]L&D3__@P24)-:-SB8E[/3Y87e&Ve2L[_VK4
WEB8g.:FeHHDIUXeUe)BbAQYd>Pf1>\I+@TG(JHFgaA(-FA)M=M5a;]D=Kf,,c\4
aBT)-\d#+S]JQ8>LP)(TX[cS=AgQ4\0&DCBSf0cMNFRK>&J&-La)g;#e2Zc;F\T_
3H#<F85=g\VF&)/53faXX4^Z=+C?g>W73Vb0_JJ1Z+U275PN<<XH:;+_LLL?6<7S
YNJ)OQ+H);4K8gTHJJ8H,L;GXLIR&XK)RcGFWI:;Ca21I[)d(PV2)WN\2U^QA?XQ
<#-@D;+W)Z3#O2<SG>BJ^-1Oc9^P>NOD)-#?A1+0fVIe]e^5c0gbK[K><\GUVIGU
&KG2SA1.-,5F8NDS\Hb[;]gDa/=9GgJC49<4gfAcSR#)9;^[@ZIbQISR#C/+E;J=
>;Q[[eDSZ?+[CT.+-d-V#<[/bAf2S[XK4(I,7geYR,IKTGTc)=(:\Og#4#83S7GW
;C^3P?Wg^ZB4Uf2ZNI#6<+6WL1N@A7:2K1C4#ZW=QO7d>YScG/Z9(,QJgR(920V5
gA,6#\BeU.V>XCZ#O916Z6eU0.[g]@0BWW_H:#A.BP^8D^ETX?FSUA6^;4ZOO6)Y
B>Eb@d+,gOA(M[Gcf&a46Q5>5BOT.&_g69Sd/BXKV1Yg:X(3Vc9CJ89J0I)N/0cQ
efg._HgF^b-7U(&KQ[9:cF7TV&2PgL#-:.-1?aZT]g/Yc[)>dMMR#]I]J\DNZ#RR
/b9_36?S4]:JN<WbZ,Z_43WM)CdFGA2GW_.Pfd]ST>?e,JXKE)CYCAHAYEZ2dPCD
P=5Q&?3_5/9[a=3W?Z[AaY@A;0^J]SIg3Z[/D)M1/ReZ5ZH7(8<H95<ceZ5][7^=
,@,F_BU1PVZVA;;/3_NB/BY#C@FHQ.&)W6d?aYIID_a+^7V&C:0&;4eg_(AAN.0[
A-SFL\=0CbV4<.Q,NVLU;HX190N[IA=4&OCLOOQD,KAK60V>dX#bNZf@B0B0H;U&
+:#7<,Z&:b(d3\EKddP,bDAcRS_#IZ]C>]eW,73Kg;,OQA/8Y]D?0I2YB.N^Q5d^
+\Rc00Z:bMJN)2R655M6>.@FHHW1,^3(U/[L52+_AU@J2BP+_HVNa1fC.Gb);:6L
[S?Wf<PP3GNU\_K/ZX0dOC;+C@7&Y-YgYDC[XUbI?BgTF]Y(=G-;;H?I8R/G@[c)
K=I:Gb#GKOH6?;-;CT78d.75EbH.e>>X\6eVXbXFX6fZ#RS+N,b-:#K]88Z8REa0
7d)H92+EFLONKO8YE-8+_<^8EXF\L28GKX&cg==5U,]=14ENMBFPVPZ0bJU9V8U^
.]C1)c_VY^5IXP5]Fe<T2RKfa.1@5UHN=3be3PYVeT/ZAT4/5FNCYN8;=X97H3Y4
\Z+=bRTRZWe@YQ-;0OOBUP4BfR<:8bbbg8fHM6_3FI,Od3a.g=R+VE]YC>_[)Z^D
K6Q[I,2LR53Kg:[RWIgY0f0:4F+/dGQ=)8&E3[C>1[bP^P<JUBV7^)PFZ(C32Q?X
&HH?TXN>U-Yf0AH13HU,=4U?B)\IVDM_]HgK><(COPZ6VGV.;)(S&BFH08U#g3UP
KMg)<J[+cSF(W^D7(XEfbE<T@]4:3]>O=_,Za-C\5Y82@L<2<7;BO2gWSKg@&)^H
9UXS[A>?)TafSH&Z/0//3)@fQO2W#Q_M^=U0PO;[^cX]]c>#e\3<V\T1UGZKg9W9
HKb8)).#,FQd<.gLdV#IRJ8X?I9?8T)-4.W;>47UYEX(0L9_bFf4gWJ_YC+dS^/,
2H?TfI@g]9?4[S^23SV@db-(Y/I[gd4.@B,P42M-g0PV:a&Q05,f,bL,R^ZcL?X4
SA1F;:,MbJO+W@X9FR/-6dJUNI[T\7RIXeF-F>6a5ZHZ^]JTX6/6B0bI95JA8&YD
G3^Q_[_:<:LW-0U[XWSf;<H][SPTQcSNG]N1gQ(ZN:@A</5\EW+Q&2S,dS7T\Aab
,PSK1NBCOcN1Rf(NePDP9KfX=E>+QVX[(M)R:P]RbbcINgWHUG-\3UPaGIUVZ)M>
31<62(R=^WZ-RVO6U=V0Z<,FYTQ.e45EKbD;]BDUGdF(a8UaZI24..=?F?VHI+(g
2JA-IG:@1a3XdQ[W1=O/GZD1L.D9TC3NAZOO_Ha(71^OI=T2G-e=R[V4UD<0cG5Q
7eU6=B4/?_<^-_G(Q,ceG;M]=a6eE=Y@e^SDBFDXMUQYa;,1P&>7\eIA?)4]#CB[
<Z=8]AFHeTP&g-bS9@?()P]GZ>4@gg&Y3I)3;LEeF\_+[L2K#;@G?9BR@2R6KIga
]+VcL)B:;4/H+S]1(3e-3.Mc^\RPTD22N-11E;0BagM(.8+N@(6?f7b.W(TM-^8L
A:KNaYTP(&IHb?T<C_gRQOgD^UB:9U18W,U4eZ-ZT#X=<ICKIJ>5Ob2<W5,Q[#WH
O8A3U,_L+A5&N]UC3BSF4S[BB.D.6IdYDBcd<2@03A\V^<cKGLe=/aG[:YIB@(9B
ST.[HY+E6JEb3R9M/ZTAKI2:.gP,)ZWd60C6P(TYZUZY#-[R@g3O8PSKOBZFN9FP
EWR3K+J<&2F#^d(1X?]\3IC.7^4acY:L=<1:4-c?ad[2a0MU4\C(^L^.099;=QW4
LLeNC&5>aa#(8VCG0NdY/3\D,]:edMEf[6-3)>\?^14X5J0HI^dXB4>)c:H47]P7
21cbGF;FX);V4GXPJITOG?a_=g(,OWYL&=?..7d^R6+20;e)P(&]RI/3b2SQKL8b
CgSDTCEJXbINC9C:PGSEgbO1De@Y^H\6+H@MK.HF<495R\VUg>R:D^1SL>P;B&07
A&32D1.1#.K7a)P@M&dE,FMQ#AcOT84NS])fB:8Q+K-KZ;RQM-OKJW83a;L_9\EG
ZX&g(MPI^A5OT<<&>FLXMRT-O7F6I=cdAEeAF8(QG)QB?#G./#PYF,Y4]PcaVadM
@[KE+46]MUCH)EE_eUf1LdQSUKPO6Y]H5YC8JP=DLafI+?c(Hc.fKU6P2^bJTIP-
-O3ZU-aLeMcEZOW&bIDaWN3<,#+0,D/<WTa.f_YAC]B8@AgEVC:gaeKW^?9P8PD#
0J8,eMCCKO7JUPAE-b?&QagKKK];AZZ18ILVS&ZO#8#E_a4K7[M(X#Ld]KV-P714
0]Aa&?/9bV<e6L-)\2FM=g9OHH5,LPX)UI.LBPWGWAa8B3-7W.D=#S)AD5NKR7CX
dZ2a^3@B(#^?AH,J]P,e7e0+W2EA1SS>@=@HQFAMG#gRK#S(=aKU+g7?0;@G48<J
B3V+f_UfU2BbNMf&JM\&3N:POYR_9L.H<[1^6I.Y)N)4DM/+M^UF&_JJ<KR^<9,8
TYUG,F9BR+;QE5^_a5<DS^&:5Z(>W)dd,QUL&G6f[2G,P>Pe\CYS/0S:;Q]cP4.F
5\[WX[85FB6VF&8LT=X5E\IKEC9U;76):(TL.,8-KW[dI5GJBF;+@e5;Z7AY35^[
/,=_A#=G33WeC[I8BK9Y>_e0;<1A+Y_KbIEUNgCb)f0\Oa66GX#R1ZGLE=8ID3&,
Ia-8W0U/(4ZDdDGd]XYNe=RKQI=H,,:5<c]60g.D-<,F\IC60)0I29cd[9;J/E3;
)+QH674M8Y90Z<5@Lf24B#5aDE\C\-C(VD1g@.cTKIZK:?T@bMEA>fKL8FW?=a\F
>5b==N3c;9;0^c(&4X_?dQ#/,+YII2)X_3S#e8;9KMX4LRHa.VY;]CACXF]0]B0c
Wb[#.WTeO0E<58[QWW79FX[(MSB:+9O^4RaJCANVT3TLB_IfR#A,XQ/VdNa0VQGG
#ISaS#M:#.1=aELVYHOeJLOM_R\CO+XB3H<d;1#:XVSQT=Oda=/=C@5A/\8K&d8C
AfLHPSJ0I=[HVRN3RP^WWd2XNJdI?NgI]=>ca)HB=#XYRW337a9[1gb<[):R?,-R
\;IJ5:#H2V+Z,@KQ_Xf3^I</U_0@T<)]:JZHdA+@g)D@_;#MVB]ba4S5TAX/]YK/
Z+,:I.KD7bbg-.\L;RYOUVS9MKU1CXPF>[;FYa/I0/AT_;)+I0LNR\,)U;+&G\H(
L\QfBGD1\&1\(P#N3bd&+C0=a-C3Y5C7bd--#THZAVU9daR=0K8=;3b8GQ?QD>aE
IaK_3,,KA:?5[M;)A^:92X.,bAYAdOa=0E.2+@fS6;#(dK\(0YeIC+15[5eG272.
Tg1#U.b-VFEO6dYE[X5;0B=,5,ZZE#D(Yg+RZ7a^L5;LZSE93SOFN9J=(_8CL8+\
[YG52C_-G/.V#BU^C0,MZB(9V>,d#0W&U6Z_Z7_bU>Z3X_Y_0WJGe>LFNEW:-&],
.7Ae8;RA>\JPeV\gg4GU4IS=E,<85<5V?9<aC3Y4.=aG6L]D[Z?;E(GWLL_U8)BQ
SD2ZOGG<7(^&g94\H],P;X8,V;4<OC&+P0Zd@6gDJ&JN[8B1\HEJIT-7[_7=PQ8D
dG-g+aIga131ON97&Oc,8:KaL_d8=Eeg^O.XQbGY:SG]5/25=[Q:eSQHWQ16cJ5^
)#3:C-G#6OGd,TaD[c<EL@48Q>9,N3VN<IVCPUMKLA(N\-_fGK#9H()M[9(\2&G6
K1N^adW@KR/PR=R\7c5QE<P[[X9]60^ZBY[X-C2,P>R/EVAHF_<fMJ:>#H@a8b-C
gW<_0HZ9Zg7eO,/K0WQ5P,BdWVebN7c4a\8PI/b\-R-;@S5N8[c\aM[\HYORP(V0
K8B/?6<6JX9E&H)_5-;PSb?@64aa0+^O?F+c_NTB?VPP5E/O]Y1ZZ7@RP4/(C:C2
?:,IQLW+>DPP02,1](&G04[FF6b\3W912-TabMcga4W3f)[cRQ)U#R<gM]]0GEK8
J+B6I/KQX4UO[b4Zdd6gMZ[c\3;^RLLP^ZS2^_#9:SeZ<U@=>=YRS)A]N93;#R/=
+/33a03WTWCH+\?-f.JD867U:5+D8VW2F4S#4W4eNOI\;2BB=B3524gV#6[[.cfR
V0J?EGH=Q/I[.0L&UPF=Y4daB<MF^J9]J;5EF:Z^M@XAGfZT\6_E4SAR.)9I0;f0
G^ORH]D;0R1c4(4[0>,O-,_SD(\B4-f?)L6#SY(a>U#Na0HeffVE?/.)[OO[R1Ob
Q8?Ja3TKH8QH670(U?0B)0&[VILXU<+gR7#V<Ye3PAKW0G-Q-8/1H;]#,(FNdYg1
PQ/^I^ABKNS<GM@,Df^LQ-eMWU9,g1GT)BTARI:EA;E;Pf_6aZ6&Y+SEZW@;RCZH
,:EBC2H4LC8(@g\-V638&_=X60JMUf3J<:K#I(//3YcbAUaN\WbegSQTX-g#8U0&
ING&QTCX)\=<49gIANOZ0TgT;X_XEGdD>8M-cOF[55cb&,JX^V.M/52BWOA9)GcQ
V8Y=OPJ3=61c7</2[MD&>Pb\0IM<IL94)8G#(g_99:c_L3f-gB_<^-ANXB+Q(LI\
E7d;g1F/I;I8R]g/]Oc<b]NH[8#Fb(Yb]>f7@/D)d_Pc02;40I&2FWCAG]6fg?JZ
F/AR>4;bHPb33H;EY4)W@1]?:CgJ_JVdK=C3RF@.Ad6ge/Q/3G.P6e8&F&WZ5+FF
K:,=^-D?]82c]Ee0GFfdG_DJ6VN]gQJcS:UN9U.RfSX==#>Y76C)\,\fR>-DYTf^
,KY2HR[=HX[gDR[:.CD-)QH_Q;bbbYU\9<8-,_4@HO(JIWSg:R7U>F+XE17\(:FN
U,f)#Le4_5@,DF_F;]E3QNEFb#)P<;I;YbD4T&A1JKUdN0D?J6W_G+X+Hc,FH?.T
@VCXPg>T+e?,ZC]<D1FOGVQGJ2\10T0fNLUL[D@;0NA7(D/HOT<[(Q_NG]=/7R(/
US5LZ222(^YgH-&;NZ=c?TIe>C1@4S2B-B4A[IXW(:c+#UQZD&34NBL+P\K,F55e
BX3d0IH-L#KI.0-[gXA:&FG<fKgTAL4ZM(&>,b)aaIYUJ20Y[0aH-)DcKGda<_PM
QDW789K0G:E1,72D#aSB3PD,QC#A/4TFIW;BLfSTD@\W6C@#Y@/2(d(.LH98D5P)
KEW507PB1[+L/3:0bJ3c@:J>\5(IPOLR_48KR.eY:g,_P+86+OHagIP\=TH1,1<O
4:RV8\#W?Y#;^\9<(L/)LHZA.+Tb-SIgZFT,9D+=@H7bd6@Z?4e<D5C0Id94gSO.
DDO<05S(TLWW&T@F57<=bX<Y<1OIRN11/4XV+^c2LFARWd];R7Mg:@^Zb-],CE&U
fbb32@Q4PaR_1^2(LBA;;WRIc[15eICK,g0RTVM_#K]cBB2^.E[?38<JB[O-VCf2
XW^]U_?H:-&Z:?#AFH7X3].g>+EYIKa>-D)(^ND?T4?,de+I>f-8c-7_;93J.30O
LCV?d@&#-(PdLD>E<73IAZG0Xe7]0D>d7W-[Y>G.^E.aR-?--2+Rf-?b[76=THCP
[4<GLFYaIVQ4[PB#@<<6ZL<X]M3_Y3]_+W(VF-L)AW+6[S\&/D63IW28S@9#1:FI
bJ]c]=?S(D@9+,[N,FZDIL,2[]>6ZJ7G,fCWG^:9^C7-@;YBC8@/SB/5e<,f,?R0
1/5P]Aa2\JA/<cLf+?BKN#XN;0;396JHV_.;_1\OF19e+N7K?9@c<1J)8g9+McEA
aDFE=bM:ag1^cVM[cWW6ge:JHd7CA8A9ZHFTE-]8@QR;W>5GZ9K)UP1(_<,:Qf#U
&4]Ag<\[HZW&(Z5Y[a+;V>F0B=Oacd7W@D4ZD\d@aDQR;MH4Q[K3?V4J^eV_1d_d
.=+cIc00G#:[T,LTPOcceT#:0T[N2g4^0&JM7KEDVPQ(\[4#:^]C=T:^.:L8VJGV
2\b4bb<Z7>;;9RZOM8I\e=<0S:.RA=bRA[D;CJe]@fSFf#;N4TbMeY-_P4<H\OH<
83;/f:FC1GeJD)?CT^/c_g9LKZ?C\IR4M)]=gBN4&de]d@26@SKEBNa2c,:/,UE=
da,a/gaODJ8#541IRfUM]2@[g0\<#-P@M[f-W1CZ6c03_7OFB:V#3X?a<eTKe[I>
ScIC)85eaI>]U8S[<KKTD+^)_<MUW3KS>5V/0E@cCOZ6.,#-f0:Te:RIg;+MO>@.
9.<b1ASOVG/b(d4#2(8GXZ-EW#FDT5M<I#DBf6:&XA8\=K2PNBf,Z<KN65YY>bAJ
73+CggB,X04AI37DFL;SMP;>;T1#@@BCa,QG-O7fZH-@8b[P297&>@EK^UWOb64b
KJ,B8_9fO#R7[,\J7A&YC@/-,,/5B+:;,BJ?CD]U.fd8B<&/LKI]>&<eG7Ye-C(_
b[T#G(>VWXd<6QH=\(PT32/L//O.@<FI-G.8,EMfVP]VHUKWC0<)NX7[XJ/cfHM+
DL5188>T\Bf<M+E0b<K4K0CeM:=g=Ug3d.LW/4P::a^,JdH-Ha;3JYHfGV<b@YW;
5WXg(2Kg9Xb@2T8U<4,W2C3,cO,bVJ41W[aHXUDa2]^/R\bD85H:gC6&BS-\Z^A\
d8I+6.U_LW/L1\fU=cR39?2X>KB9D7=&\fX(C,XF7UY6+c]&0V0dfB?4cM\>2OI&
^A8FDNM6BCc6B=7_QIDZOD3I?P+#UM[L19f,c>3,J>eKO@SFFDQFfBDWR;)&7ECG
8QZ9)3=2LS@T?,f^K0BW.8W-Qb25=T;BEKg3Fd/7/<1_O4CUJBe--ZC+M@\SgWP-
D7H+L/ZLP5L.+@[+OMURY@9&D@,c?[<:b6CfG]88Y6fE2&QaR/IJ,Z4VF^GZ?S1D
a2LL8gO.#3DVW=:Q]5\Y]@PKIOL/^]+QI>CS5/VVc\PE;P>WPdDUY3I\J]NLa1:T
2E<9A.W+Tg^R@7&K?5f]7Pa:QAQ6SADcOe9^fS+B\HC:PYc#SP_:A_RI]NbZL4KU
&IY3>gL5I=Zf>4&aM>]bV.#0S:WRe4Ob=5dbRcZVLENYc&8E<@OED.FdBIaN.Ka.
KMMW@R]B97<b&>]CD[M1_S]df\X^@>bb5K6SSXMERIFM3W,-?OWGXf&+c>?H?>C(
fLcL(3.aXWS[[#A4a)C@&TfNQW31H/&W9K>faZ-a3a^#F:/a8G@#8@EId;=?fF3(
<)N#;XE0/E.FP=c@d]/cC]_W\?f)30?ZK&\PRA]NU1Df/Ce(2-=0X@B_8&.CQIWO
M.c69Q>L<9_6]@5JUXQ(,1:CRX<T_c0KaLKJ7_FYE35S2S\^JFg7@KUD1LH7^OGb
_>MJ#/,/dBY3T]Lc^WUVAZALNGIX3C#YR,V]E][g_UVTdVYdc?Ng-c<@IKA&W8BV
H5ZG&VN,dDR4#O\H<M,T)NaE)7[98^c@?[dEH;.?YNaf2//6GG9<===Z5?4c-0&?
1&PKMIB.36#@=K4]_ZFZ.Z&M0c1WBg@DR&[Y0,B=K;UOR@<0VEW#Ta-LUTF:?L1I
;NNH=EE5IgLEN72==#CE)VU81@/\UZ,28LM9eJWG<L(6<Xd\#C=C873)-=:eXcD&
;<eI9?AcHGdF^3(>@I06KLEEeYe)]Kde6TPc+R[N]QSa<?0Z_G3a^d1:2#3\ZI_J
A?,))ccFZ05cbVICXH&5Vb<#[+9>LYaU@/IAADXLVb7GP#b(&UX)ebTG.F9B#Sg2
/EZQaH\==G/,aI@c3YdNF/IG[STO9#\(J4I^8R&cNEG4NI/>Pf4&CI^POV-bO;Q6
d0GB[17H)]P5PVKRgZJB7/HZ@G\W,a4EW5TD4]QO;G5^D[>^bC)0\5cHE@gO-]fB
c2].(HNY#J0RO-=f0J5V:DV00_I\<eN3E0B+:K7PP\TQ5NQ?I<EK6+^K,5eY>\E3
,[cZLK&OD7G0.WX?P/b8eWCDR>=H6M6N2DDZ/,Rd)/^^SAAdVW<>FcE7ZLZ7aC<f
c[=T:ZW7\<J#[bZU778FMe5Mc]2ZALg0V.U0a/gR+;BLYHe8O3/ZB^C>N(adDZ++
bOV)-aXCZLM1B]T.dVQI6Z<T^XK-b,a/7,A5[W\^>PBW2T@[ER=f^-@;_+R@06QJ
4:gc[E^=_Y<\AP>\#O#:#aH\<0A;<R=.9;0<bc.#)9I3g,gY=^[&0/./1DYVW6bC
EF;Sa+;Q9;:/6R&Zb69)\TaDe:3Y6gVEWOPI_?L5P<:,R4N#QacA>+R^Aa/8cA]f
_V-(+<Mb@cUKO]T_]e3UCART)D&FQJ,P5aP<dB<)0J2(U:W5PP8N5-Z/f@,/P<g5
[GZ8D.:aA08UEE)WY03<:dM=U#\XTZ@#;^9KU]@T+GDf6]CEDEAef2Cb9gHZdTBG
?_1]:2S[^dC]\FeTZ@dXR05>1=5:Oe=3RH3XO?Le49c7,7KZV&Db#?DWK+>DI\bE
cOFdM\fbTQP/B\K@d]<W&bRF<R/ETcG.]<,2_9Pc1[6NMd(_-&#UPXIJ)fRaI0F6
MTX\EA3R5f+4>YgL&eB@dS?d5BDY[HOFWDa:6b8GW4PcIe2CVY_V@f_bFU+7I.-b
4.KO((1,YA+@)Yf1MeMR7#A8RF1=:=U_g+I]242Y3]6ZRA44_34+P9Ufb_T@[,,C
gNQXHEEA4-1JG5Y22[2E)1\QZ_@K=)_eR=g6;@]DFXIHLA^aN4@E4(_:CfS333-H
]d=ZP@@)e2IX67dabELbT5Q4V]GP6d/JD:WW-[.eU3YY##KdEa)ga#5G0YBB2;f3
aM-,<C_dJ(dYP<U^>2bKZ((WAa:@V))658>_##BM,NICPKF(9MMF20+8c/P04-EW
G=RX@G-?6Y>cK6#g4,7]):I?3<]c16;(Y(.c)b&LcAV#c&d0>N^HDdBX)7IV/5:1
_FC2/<0O<=GM<3eC@6;)\d:e[/6O\M^,^^2,:Y60=3]EO><I[2b8^Dg029a1Y5G9
HHJc)0P<@#3b:UOb\;P_EE4@Z.b)X>EX]J<1VEL8d/aaAaOfHGOULU.D.1Y<Q;90
CZJXLHNZ9P.2&>:KL2K,:W5H7#Q/ID6O9(;-<R&1ZD;cR-AZXaUCCJRaNZS:A<fY
>:X2]#Z]Kb:<4(/A7H6?H[f7Y^[gE#+7RZCMIdV)E1gMYaFP?&YGYV#8=\PfB9(Z
F](T4EAR448_^)V=ZJ-3OZ:\O=>]gf-Ba]O79T0)b@APNIZaaMdWMD?W09Ie/Z#U
9OBPO8a\.,W-,CHBCa/UK0D?ED2a(58K1]5/T2\^cR)LI<7eg.E0V42CVFb<^-#]
^bT@6?#(IN/<JDS4V>EA9?ZY#P\\IeM@XC,K#,93NY)TP\X&]H-@MI6&#3NTbOJ8
<<?W;JA7(A#T)a3IQ6Z+4DMFRUORa2a6b]=H+e+E:(CBf6aeFdcG^-1K+P,&0b^>
UQ(f4SPG8:+-0I-2:RKVbM,[^M^B+3/3[<^Z-3ILJ^cgNN5<6-M:;(ZAd&CQg?@T
9D42;cfY,JD_].)7e(ERRE/:5.SX2(;>b@LR[(GYV=4QYCQ_d.JA)M-b:=/L8V\B
6.-cT,O?UU38.\/4OEdIH^YX\TE?d:HOZ=G]8aDI6.d5_6_5#Mf5<L1W;.:(]=R^
Q>>^72,Ke[PBgeQ#7ITOF9Q-;6^+?].eb^_&R6-dGTQ7#S;TYZdEZP]NbE^L0H,7
TCLec:.^7_f\-(6=e:\.OE-#)4C=G1J+8,dSW[WfUH#0S4A:aN)@CT00bZG)/De;
BC3]Ua-E9f:5+g8Da:96d<+V^J3[29ALP8B]&P<TDaQR(=#/SE6=9O0baV879P#@
DDbe;Hb\G/ZX>@)?A6@gc5VH^F@Q(_-H8E,efFE64V(X+_0\<df2&CO-GZ@.eO+X
aW=NO6B)W]>GI_.3GSB7/2??4b<7FWWU#aE\A9M)>:2>f-4[5AS.A8GQQP\ffTeR
;)X&:<L:ZYUWF73+3RdECP053)&A(B+OAc-B4,NBAZ[L9-EYd:Sf/L+T?ad7OLKA
K].UeW2N#g7?\#FOZQX/UMLbe;NS80Se:(V_@6,-#]PCZ;IP@9SCMC3:_+IQI+Uc
55>.F=eMFc7O&O^IdMWgdaJ]3+d61B5OfZVdDW7fYDF,^AYHLK\<6A&b[_ZCIe)H
9@T1>/d-IGS6I9Y4\b#1d/MB^OJ(;E+\DBUQObfWW@_:)RBLT7-KK[C/])NBG\Nc
6<1P4^OSNVOa&TXbCNH74GG-U^OB3,Y.PV14:c>9T?>CNE#;,KLL&W5ML3a^AKTb
fT<ZA)WEc;7X>OHg8NY\:V^PG0^MdA<^G^9M35Z]ID\f\S&S=0?N>A;:A<-J3D0U
N31<g=]R+AK)K\6QZ3A03Yf3He)7fII?H82AEN_dEPAXIag@RB+a]LN3PXNE#&T[
[eO@(:1Y23>X.23-YQa2[WY\DYX[T-1?[:X/5e,@]8LWN6L;UG_1-/<Pe=6W1[KY
XNV_X<EbPCI7<,Wa#gE;IRV4@S5e:C+FDA0V(+(WGB?KGFK[?I&e:P+4\[PeB6<f
G-AV9XC_7@>M6SGA]DI(_ERc\.\3g8bT]7>Y5FWC\=G_&GHNR?E47T;9FU/;>,P>
&_/19=fd/=XMD@D(+Bbg=TK+V8&X@12U:Z.4\J^3Y)b96K@G1[@T6BQd=NKXJb,G
\e@CVE1Q:/42CHcR&g2##TG(LVEZR1?C#@,N9Q=(NT\@ZaR+1CZ&)c(M)WLJ9XJ\
#CR(5abM96TDGbBYM_Hc#VQ>:[2?1d_^+Od<,A9feVJC4&bfUJ=UZUc\NaZd7WJG
dBT1?<M0^728?)0>/]fLQ)0SD)bf9,KH70Sa[-d9.VN4c(_eGLd6=>,<^74>3.2V
Ke6&_)BD9MAS9[HN)+/8&0-1&&,CS^,>#IC2?B@S3D++-9c2@LDODAAE<AQfZDJG
?@?CN)=4LZ_eKT::12ZJ,ZW@^/>K)NWN0d#MefGB+>M91Q(+W,g9@XH(NUD<HQ/W
:[/gg0O(39M<?]03f)7N1:a6+28([S=9(06XX.KQ#Kea\O>MSbHd,EO6?3FFJc5O
Uc.DggPBMUfE^&1c=7Q^+g<O4](0>]HdFX2.NfT\F:bYH.cgD:BI:1+37CK:K4^Y
#M/LH,5>R,\FS-#e;F@_/_MRg3:I<R-b>=Fb5RY7Q3cB[>Z<S7Z@d@+7#2XEN[UJ
ceV/BAVf:\&WGcba@B\bFZGa[<EIdAV<QS8FD16?V2If@23bQ4OJ>;,>fD2MKZ_2
NCe/L[a:\]ZH^d\MGKV+FLWX>T6)?>#NN:&V2a<8#2TQ]OF:QdR.8H&.-V.K_4>,
;Vc<>CbSBSVV;,P02dO;DSC95E^KX@,2A>)_.S)A6B4?ZaU:SZEV,,MKP,Z5A>aL
UdJ<D7]D9B8I9:6&[ZE/_@O_2aYEY(VJ__+BGN,3)T_ZG[Hf5W/P/K&cccgKJ1BF
cIZJ\_X8TPe>23,bUI43NG?ZH-8Xa-T2E3M9Z(&>Q7C<cOf+ffKY:.Z_gP,^48K\
YQb7d42f5G1JO\P<SII)7dU8gZUe<S+U=bB&K1:&.-)FO\8^dYf_(1VB<J):b9\)
b>B=37d[WZ2Z)A[#]dTKY2A,4e)IG_M3D80]X30Hg05SK?;<UU0>6U2>T4^T;643
220.-cXYdB?R),6gG])B7If)Td0.U#;4@Y2?4>0bF1PV6B&>,5PKY.D_H#0B[U)K
@NR_5>Y6J_:](>C)FOI621P/M#2>3.M4VNWTaL1LQaUcC\N_SLFZbPOD;<68f0=4
3;Kf//<?E6bHaXZDSH4/6Q/4;B:8^2G7U?((K:^.B0I6eQ5fP+>Z(Z>b<3?],?L?
4\<+B;^.2Pb)\8CVF:[/e9Z?b^^0(=GG:8)g=^(b\cDFXf^^FTS5CR:PU#O.ENLW
7_9THa<5gE=,A@;+5HR?N4IG2F9g8F]6&5Y[QNJ_N63d]&,76b/Q&OT_H<#](;BS
MSO8H9@IA?G[A<fW\8WM1>](3c+?;&.TCG(6cBUeJ=d.?5C7Hec8DQdSQ]V2GOfI
8YJ\/43bZ];?E.VF[/DTVZYT._)I?c2CCOM&JXLHL=ZE=BOE,LfX>=(JHgP^8JHF
6)FgaKOd]:3ad9(>cFQgANcOW_cUWPbVP5fEL1&0W&(HGKOQY][dVeL&JWAeQd5K
71@:f^D\M^R[1^+2_8^1ZXY3_LD9YTF:BfNAH_?Z[g6Rg\5eX:/KBEY4eOdEQZSP
DJ,?HFVD[LF1e_WI_9_bVOe(=LDB;W)S,NS\82Sb2JUWT;/Z5YRPC2Z_[eOB;_,:
ZdI1Sb5GVFg41#E4L4FaQ_/@SHgb+fCH8;D1dRgQWWb_H0)M05JXgU4F/+QBX\NY
bQH#TCF+6I#T5,KNFF6D+:?A&?+VL=KM3C:c[G73e_C_+/0RL10K,=4R6YED5gTA
,(A#=R3J[4)BHG+/Q+_STcOKG#)[4=QG16YCAW\<17c1X3^Oa.A6]W;20W)fa9dZ
\F1/U0RfTLW_0Sg\eJ+3I,dUadA)@YNeBaN#L^3,R7_^Pb^(dd_^<R7TX2cPa_00
^R8CQW=1.;7GcTa@2(;1Zc3I4.Z7#UcH3Q=OACQ3PbM;L&AOLD^UL3M>2/;]C)<E
g-A)Q-4DCT;3]gM^\>DBR<;QfeLO:>1:S81.EIRaSW4\MdH@WgEYQ:Gc>6d60_Z<
IQ4MPE=SR7Z+FCcdF;:LOL1YR@3LSHNYV;&eNU6,TbWJ)&g#ZD:IGP\IbV8E&7SX
=b2<)P/MY?^/Z.,^?2)OJDSQ]]KS/M.43f6NWT:EA3MUVNL,[/cU#EUD]S0^E=b6
WJ6_eYAIG@8^]6d+2\X?J2T-8FTV\VbTC@\]>WRVEC4&e@J=Q0#._PWAPR#ef<Hb
SU?fOgU\6X;\6ScFP\M31D=f?/4@@RMU[(-K])T[D))RW137/eac-^(+Q;cZ&A]N
KBBVg^d]D]&Rd-I-Z=1@CS<-R?Eag]9:d(1dB2:G^>AS7dP]3=WMSb75\,&G.=SS
264dI+JM^V^O;3\R&>7\-O#>AY[03f1[5bLZOXG5-;J_=40EM0^g8HK@-HVURVXQ
0@\@\fGCUgX+c+F])Q7JH?46Y9H&[YN>O,>,Q_5b0QI\#6Ie.TMDLbXK^ZR4S<L#
QO=(=X74W=7cWJ^3K+a-Oe-[A(WI:QT;3fY:Xc;]J)#6:T1^Y&L@ZFEW[@/TdH7K
O],C(9>C\0<a<I_,(12bV5841=0;K<aCMfG^UF]1eb9X>QE1CQ]b3YOCc#;:_,Zg
HWYU?cAc+-0?e&_Hc=DI4NSWMNKcZ^O(KA88I5aQ/cEa6RR+G]\@VbYJA2AR72\J
X>d[50+[)G_8&H^QG//I2Ba@-H47+ZP(W]g=e<@=8423bc:#W6gF1?AL@_>FOAd5
@,S1?H/>8g]-ZN,^Q-YKOTXNe\=OY[:^-;Z(=JO?Ta=?@dd&7/-A14E64=Q;I1-]
.[.0#aH)B_6SE&NOQZ1)PbG2B>K)R&gE84]-,Y?W&3]fKW?\D1TgdH#_5=-D4GRW
VEb.-5=8DD39DOPUL&K67)IM6e5Le57YLTA.(4a#;gEgg8@USe43)JDc2PB#9QF@
_;X.1@S^GH2[)UWQEBU5I+[)<FXNVbZNHGM9bY#O-SA?)B05#3^=UM(Kf;G;7/4K
G#O_E0L:43e:W4f@C/-(^K9<:X9,VD0^Z2.@8EN&ES)@&F_g<EaTGTdSO+K,7:N#
d)c\/.VXePY3dc_;a+-Z^WY()=92gbfGdTTaHX\gYa&<<.WSZgB/-?PHNE_ZJAGR
>f#9_(cTSbRZ;,:I<AFa1)A-]IM0fP-2>JJ\X?3BX/Yg.0=5=OPQ)]&E,aKW.G(+
adC&ggQOC.I25&-F3BLB2@LJLgJI]+gge62g:C^JN#6a_[<CA.\;6KXa#H/0FN3.
g^RVRM)R5[XOMMaDK;7IKO[)-@Z)T.F:OPUaYEUeBH8YPC2:&/,OgZdW,^&H+L[;
H7436b4/TS9<E+T7UWJOfO(9RNDbDLbZ[1I]@HX@H\A\HMW8#YK.8C6<H&MbYAMH
M))HE]+<>ae+EPJe?/^F3a?D/#aUPL6N>TZ;O9+PMQc1gf?NAVS7RK@\bQEB#?Xd
F3<=YY<LW:Nc=_F[Ib.84dSPgBb<J;TCJK\(KfXT]I,3c/;U[S+A,C5GNBX3b;(b
<_W:\]M?bB07+7ATIJ,,2==IeSbdf@-=_UaS=\?_A:3G^K0RSE&Z]5.86G9.ePDD
;PL/JTUZU&3SINXfQ<fB&e&,EP:d3>]SJ+g=HQR@)X>C=QU/N<I#5(],1>O]X[T.
I&8-K0IF>4YP#:FN)Ba<+)SJ@:[#>7<3@cXg><H=-aZBP>K=X6#Rf+F[Y&/MLD0P
&aD)D-?aZ,87+4#Z8?eMF>(2U7\9a]6+gD<e/U68J)K\XB>eSHC;O3:&bbU]+O)M
4CYc>WZDJ02a(KUH:gT#--CTfV:cfM/7-7eaB]X6=2+#c=FIXY)TX;e;+O1&5:W@
XV4G.+6DI[0e?Q>OCNL5J<XcH)Nb7cc\KS@KbG)I?F<=UD8fF;5)8@S0R-SN/VX9
@@?TQ/1)cVEBUJ)bbU=]EZgPR<)bEge-FT,+:FHKa/g[8UcY41WfALbB](]e4+5<
Z+WAb<Q/gOS7Y9I]EZc?#a<+#)Re.[bfKR4d7EfLM<.9.Q@_^_HO#FX&;^)7>@dg
M9P3dSdc]/-CX=&L<PQ[G]+@Bf-3#;.2Sddg:76+37Vd<P7_B>F42gL2Re(Ub29Z
fNC.cL&I,^+,&PH+1_\HXNaB+\0ISLXJ&AL,UFAZ<36KWS4M.P&Ge^3N5fa2S^EL
G,F3=46\\YeL2B#g;.^U22U7BCWT&R.We^Y7&VC0f+#>F>@H<<A&B^B#3B=NGe/<
8]O^7LD(:WHG[d722G-V;IKf7QN[]]db;a/QBa;eU]g)9bg@3&AV#L<N(-K#<(E_
L<2)-UI#Bd1X3b\OH;72+FQ[S6^9^efKcJADML_)47C_IGYX6_]F_GXF:@(RTU0_
:G>Q]=4><B/]DR<:86Q<&?B=[KHYJX=>FA,7H1_RXS0[CT[]\G<<+P-<WQZ-1bH&
]KI,D]N98;O\c5(;D=E/V^B@e@#YSI6X^1c1TE3e-gZ+.LYF6^gGeW<TR^2Ie8,L
N@Vg-AE-(M2K\>W6]dNTfSTGBfVN/EB;<AUN=C=.],M2VM)PS(JU64d/e.G,W@_L
MJ;=0>=A-HM@;M,W_Y+RdTEQN0F?ZPIc4;;EF-V@X7ZdJCKJ+IL<(IHMcaF6[Vd:
-QKNRYeWbBbQF+R.S[LHS+1gACTN_HgRLcR:(UZO.-?)aOCW3GR:fEY_d4P=P@Oa
b4N1dY[:IO^B[SZ^QHf8-0a+d8-L?F][>L.T.Z(bL@Q@DP(4,,AQgG6C=?5T)DI9
7.X_^:D7b6=.d[Ae\QY+[^=4bW@I7-H33=ccg)e6Ve\RK8Y@HJ]MAY,-?MGKSeWP
\+7@I5KVaPX@OVXdcQ?9-b.fEa2BR3^YbUYIO19dAN5Pd716YOIFVAUKYeFC]RO2
^bSHaQ-0X;)PO^4EW24F:O/9VAXPS[+?^H7;;EJ;YYU=&N-H#8>Ic;N=-O.01=SN
[1WUL;8([DMHad]PPH-X@@6a=P?5c#/@=YBT6d&NP/f>NC61?>&d.X(S;NA(dH0O
J(,5WG;UOWU@8Q[IfURH,I-dV52A3?45O_&\-1fMH1(-,]]5a<GeDVHbEG=ARb[-
B0d(/S2abJPf_Z;(EO;RGg8H9(\V:Je+bbC.N&SgC4cc^+&=0::R]3c@_1fB8d2F
WbY8K.30>MQUX:9BZ69&MOW:S4bf4QC;G1)M-8V:Da05#6R1Rc;W5D/-;^GIBLWD
g9.>4Q2OJ(^#K.C;:7G)KBL3UaC\[M&KSb8aEOCD&:aHdJZOX\=/Hd)Y+DRgL-@#
gb-[O+F=LbT_BHR8B@dYfEDG68H+\<.+.6/J;[(W8-WDWMa_83I4FX?^BSASTU?(
[RY@)-9a2LR_,6?,dceZ-_>b4WA/5FWeFYM;Q:-6d^;4e8+>LD5b\a:LC>JDRdI:
gLU.?TdV>YR#T;OS-#0=/V-SV3&AYf8Ge4@+]W(R/ca]W88g[11T3[K(1XFRfP>C
G1ES#^IQNK[e]:gY6P5CJ^g;&PP:[QHWGJ1=c404\EPba4,TYIB^616WW:K^N^-/
O],FO+Ac.:SQR(WU>fD5f05DV.P\_UR5[WB+48^>>75aGa9E:V&RXLdN1E?JT_O(
be0S3K(Gc_b60;?^Hb/<\XdIIG?CeZUYd63,31Dg6Y;KOM,X^E23=?KMO_\,;5N9
:^?<^H;dIR15O[=?6]DaH3b-NcU^\E8:YU?_.Hg,^3NWNNLUUMJbXS.a;\V4MIH>
21D<d,LQPd-S9&.d&W>Q=81-a\R(6HWKY_YSB<5U@3>Vd184)d+01e40H//1;5.<
G;0Gb>1D806+=E&JeF,]^dLF?bQH](FOBcN/LM/X\EZe#_e]IJWeTQ\TL0V,7M,E
DZEHB]VdV\)f83W^cD(b/K,Y@3Q:IaI+860_bWH-3d\Eb06<.)5fX9[,5e#5fU/c
K,W@ggFT>((6E+bg+J1V6KQ8?f\UcaR,,GF?gfA\b9:&3gQSFb?P&]:P:;>0QS8O
+-RWJZ>cJ8Oc/7.5Q4EIaOJNU0b(&7e]3O]cM&0.IO4AEC_K2D11aN.a[++J2W9@
BDSOVW,Td-38),WgT9d/E^GAfF2-?/=A#d#5M2=/6,7Z0e@#O\d\]dMa?,Q:8U1Z
&]Na4]f[91P3NE/PK>]P#W(SH+;=A,HT]W-b?3A?dG3IY2QD?J,fMSeEA)g(LD]9
/2aSIA1gagZ>;4O:a?2I38bW+4(b7P.931X(>]JIDU3b>&8[aGDI6;E#_@4G&Rgc
8KHDV4#K-R@S91TB[\/>a0^,(S:8IRGW=UOH+2V,=68QIK]#-XJ4XES3geH=CY?(
ME^T65P/D3L<&N69Y^+),DQ<0>/Ye(]7MVIAIBAK_&cFO^dFQ[<Wg-PEZgZ>&f;8
M+=eS,-ET1Y7^T(L\a&F/b3-R>V_VW3[6fD\QO=+#8\7=(PbZ]W8T0H_ddS^IgYN
=#WN@+MNTfJd=57Aff\^3+d6TN<8bN.9VUc&Q@?P:LOQd.fg2e#Z8f6O,1eb)gAC
>[9RM&G?J:9[d:S2BP\\J3ccV?d\db7=,bF@98P(UD2]g<I/8g7I9ST&/Sa0=1,T
);K:\;_&VI:IfNS@X:\7(G@_E4,JbW7DGFHE2)eN<M-O4R:_+6O?_:4JTQJ#WQdO
.VHM+cC81gOgDf&_@\2GN,61,e^3A_=JWY7NN^0R7UW<)LCW[PD;(YW-U2N]GO4+
0,MUc8?P]B-+C6PedC>f9X@-BD1gaca=Q)^b8JUe.&T[+[.d&A\:5-#1J4A0#+A>
CUT45\#db4Nd?W4J9,S?3?AgL)Z:NJM2YT2>M&8X(J^JTDI]4JI3GR6(dPZ;Y2AX
fb(ef9E#8UbRYBcA</CJ44#&F+&AK[;<<MOc,4b;8;IBa]Z2d87<DFK#9F);(RCg
AZ.?DREH:b9=f;EMZY3fcWGg.._/X3K&)WXTXTb.1(.LM+@Z)NQH4?N3\_ZZ^7Uc
J<d(MS2K?c.G4Z\Ma1C4&_bSD?(.HSb[^^dZ]0d)[10DI3PV4K_AK(@G8.6HC^fD
H2+4g]TK_MDQ0<T1D=5>aNGE5EcN[6:?b]KVK,G/#XASGfG3FIaEa(@IY8I#]dDb
T]+3N+5/[O26(>bc?Z+PUa9[TM4T442/Q)IEUQb+41IWW^\MYSL+J[B?LXO\9(+e
)=>VML_USbE4b[d[5c>>gU^c[#8eN<3J)QOAd2A5X-9KJBK5e#G62Y?ceBJE_dL=
^&_3J(KfB_+F]gG#.PT4add_YeXedbfa+#AEC0dFZbT43;dHI(+;5_8=@P4BOg/H
A,I_NIed^]QGH]Gb:fR0LegFJ[VA_]f=:;LHXY)@-11<YKeaeE>57KgaXCe0P7KE
G\VVX2[NdZ9-gY3:]F-E/B]/VV7+1c5D3+6A(5T<4SH(e3J=DCc7X7EI#H=.c65f
>a9N8-)<@H/Se)W>C.bGI;X:VIZ=5&dV/7bV)+OKgRd?C&1aFQ,1;.0@dO:>M=)9
Z>2La>ZRI9g1FHXb3__8BE(b^-Y>=A1Gd3MNVe>?2P#LUCMdIcY3PXKTCb.?#&<)
@W^_bM.KP0eG?&[OZ?&NYJD;^6X&UZ2H]e5TV^6@\X>8I[X#/7KQ,eW4S8cV^ZRC
CTU]JF^-&?\)]/&QI)+5gaC6/K@(SC-:ZDFA2CaX-gX#+3>V1\,F5P6PZ?Z^VX+X
03G9.I4e5WY3RS(YTO?PII;G1E)MU]H(9LTLUN\WR6L:6#Y4L&O,^c0H;/I_\<[G
3a/cT6=^^+OZG49-g9=;C3,@dBgI8&KM?ZKO>TQ:,(U>53cB)Yf5\1Feef8]KfRF
+N[cYY>cdNea]+@O.5_+GBOVa1WOLOBKND3K,>>R.abR21]?B44K/d4K4NgN-ZBV
E8<F&P/HCE\c83X[6WI5)XS-daFM?6]HYfP(C^fMZdPD=WcBbbSbFbagLLQ^A8>g
I\F,/aNf:cGd,Kg&IMO9>Tda5ML>?f?0C(=;V;],-Lg3?]2O3>E/bZ5g5aX2A+YJ
JgI7?\[GD.B7]RP4JfTdS+J>SN#aZ#;MNDFD]^4K4N9MgR]a25#FeX)?-Y-RAdd)
_)f].He&)P0Y-.AMP#\[7Y]RFG=L:d;QQHbUa8CP780a&Fe)dREZX<L?^B,a1B2b
7,2cc6gA8gaF1_+JG1ce93S5=[:bcWK>6g:NZa8Kd[15ORK:,M/FcI-:J(_LT.?9
D;fSJ;L)910?#95.fK2LMUb;.J]<BW3C8UGRUgNZT@LJdc;5/0c[ZfL(>Y(/cN\S
G_Bb_[V3ZYC>5ABBI2fEPU@I0S@YB,LbXP@AEPCbRObDb^<[g&.2.QRL>R4cKbg\
RZXE6_1D59KUFbL?+(H^#1CK(+MH4PJb]f(Bf1+KT:GVGK491COaTDEXFLG77cDY
_1bD06A5[EWEBX,&\dTQKOLcE>1c[6gW:A0?8/eR?K?G#/?-?CJW#/UW]TeF:X>8
(.cA:PdK0MbK>GL9TbRV:5=K4P>\/fXN1][M=A.]-@SK6,3949CG1\@[:g]SSX5G
RfF]C,1EMF@)C=QL(3V^IB0Q2[CD[4DPO=@R#eg1(GADG=;-.cbF&-]gXWbK?FSV
:2H]Ha.D7#DQK_0XK>DD8U)\]_R^+Sb<OYQZ7/VVc>UeY0L/1CL)?SGY:FTXTMAb
Ld+6[J_L<;HVXO@>^)V8>]MS(X1Q-Tb6:Xfg#^J<BI?]2OL:)H(f;8DDD8LKe090
f@6/R4THKJE9N4/R?R#-)FSGTKLDX]&M#5KGaSV/6.df,+[1PL?a;I:UgVfR2F^@
K]?0#N4,Q-M:0+9&EI98^U:dNILM5Tf=Q7.UKNMNDH(/.5YTL&a@M+5[W-,\-1@L
V(>XPcT>1P2eU1>P8)/g:RaZGQ9<JI3=,G@.&Q,II7Jg+Y:Q3;e6/(]#B)5A_M[N
[)C=fc?QV<gMZ3b>)_:5Kd1b00GeD/9XP/R^W\VP=;G.&[a_505.>X2^O^Y<BB05
#@gNU]4VCH;Y1O#+/@\G4=<ET0G26PfFV)?NUf=SeILJ\M\c5HB@F45133USI[d6
+K4Of<N12DM^7(e@U0cWSS?C<2#S=Y4VT1;5HEH2b>9\<#E8UFCXf;XADZ9#(f.(
1VVV\]4O[?,60E7@Y.9->@+5VcEQc^T-+YMD&Bf&[C(RHe^,,SSfB4F^#-6[V4YA
6H73Z^G;\WN\gQJa&=^MV5ZMBX9EC\)\eIR6PL5b>ccMB7G<2K]7S?d[[dD7M_94
(:97A/O+d2K8)G0-bXNe>[JK_.6dd9^K=aW^#;P+RY-T>9?V:WVGF1DZEE7ZJ29[
AAH1^0BA1&40-M,Z^BC.>&Y]GDg-VQgOW?KB;\6GT-2c3B?^G(&.0bd04Q?U#:8+
Z5?ZKe5X^c:??a8BL^=5^f8&Y=0^K1Z_.WT2fI-M@)&WU]\<R-ZP9-(<:=B(3];/
#Me=Y8e6:a>3c:;<A#4H-86d4aCA:+,9<(M_e6Xc#JRgSSP9M.U>bC4VVYLG+WRY
281_M1L9]<PZ>277b(#KCX])<Y<;OXFDCMQKYU<+W<4\b(7B:<FX2.4VL$
`endprotected

`endif // GUARD_SVT_AXI_SYSTEM_MONITOR_COMMON_SV
