
`ifndef GUARD_SVT_AHB_SYSTEM_CONFIGURATION_SV
`define GUARD_SVT_AHB_SYSTEM_CONFIGURATION_SV

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
FgkzcMHRFzAdi6fI+wAOKLd9+r6BlK5LS9VoP1k/skE82nMsdyeYHb3lKzNfBqLf
zXjfgQjSP7uWL9mAYdFxmamZIGHSIiEEZYN0SooI1oO+Ct/AK1ZuMcjcPoO+OV2M
y1X768fLINCxwJ/l+VGFqO4Q0pgQiaNLy2iAWShC1+o=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 1054      )
Opt8wklFVc3gruFuEjTY06wPQOmNlX92fWbJT61ec/fYEZkoZUZ0Hu4tVbhCC2a4
72eyzygIjzeWydmkwtSjgGKAjbDrbCeGmz8mhDu6LqWXbTT+tdekkFpSrpxk2q6+
6ATcMbmMg5IwQmlxviJpt4GvdbcI5JIwy9f0Nerb6XD6UxvNX98kFgBbbGSuPRme
ccO8UTzHglsHYg5wW9A6oGbpeLKWScLipveO3dDAHWbN88uq62bAXu9pYV+QXSa4
Acz/JDZqsooziKg/hT46sOE4ex0DHx1H6040k/cBCv85G+FukIpleroF7ezdook0
dowG5QWMpfFqJQV8aebCSCjdFayXu3zV4DIG2w/FZo2iYIgSozKMX4I9xlUDOtnZ
j3k194IlrlKSSL5l2jFFPXNuEWqnht44x8H4bXs30KcHfnf/bMQeJYMCmIMKiUCc
UQzQZPMBkmEkNXMKN9F2IolbR/Uv7dsqSvGvkmw0vV5DGdyRdIlYF4B2oqQRo3cu
d32xYQuTZQXYV2cz0jlEB2JBE9xRRQmZeXhEkCxoUEY409NO2hx+qsp5cYAq02Cf
jwI36HVpDSBrxHTCeEA5FEEv+RypJeQuUtavLszHi8S+pxO7oFGaVgCUWgXPi05r
wJo1UHlYRlXPGOL+4gtz0z4T9YfG+Um4wbMKFac9huiGA3TstS+tWNtXrxI/8aR/
GpZtQL9P3MOo/EjGmBPFFJarqe/B7MQwOZ0FmEgUhldbXiidGgcXkQfzwIkE4HQK
Z4svHbUlAsLIw421uBH7msZ6iVPGJvRPkogOvbhXX1PQRpOjUe9/manIeXVcSYHW
+qyW9mKudSVtb8amg0hDleCsmMiJIXoK6QK9SMOY5qbOPH/DiUyweTR6H5vxSUtl
74Mpt7aW2qP0nQ9z2SJJT5xj01gFxAGQlxNGbug05fncDt3pQy1E680CUouwwBKc
/6GJFRAKidPZLnK6kGYW1ZGksTflwkyDNCaJGWPQAl9LMR9w8Dob7vsyxJausA/u
gT0EWDILgz409s/1j8wHPkjr9Pb8KVIyOgIYlOjPkpyTvm6QSAii1y3KaQx7gslk
dvIRCsZSY1A+zzFfZsYX2IR38gp864ummsrBbMJSx0xizx3TwNOju79PBhAr5FZy
JNBdBL3wRJphw5NZTTDBgyFWR2wSWlxfRTZCuoz3xlWt+ncCP/GohEBNR5lVMADq
eSemIV7dyifw58O8ytzJjw6HANUJbwmwC5oUce7M6gbCdfoCW9wVMDD90IrPdJJG
R2geeFnkLr5Ap6WyxqPWJDnkKshuzli9zsHR8WVydqWZmBoMySmTYleKb7/cyR0A
4cI0lOJjz6mJUueVLO/L0rzUJyDCFDZgTj03Zq1+PHhP+tFKhvqTxAYXqYUIHPb5
`pragma protect end_protected

/**
 * System configuration class contains configuration information about the entire AHB
 * system
*/
class svt_ahb_system_configuration extends svt_configuration;

  // ****************************************************************************
  // Type Definitions
  // ****************************************************************************

  /** Custom type definition for virtual AHB interface */
`ifndef __SVDOC__
  typedef virtual svt_ahb_if AHB_IF;
`endif // __SVDOC__

  // ****************************************************************************
`ifndef __SVDOC__
  typedef virtual svt_ahb_master_if AHB_MASTER_IF;
`endif // __SVDOC__

  // ****************************************************************************
  // Public Data
  // ****************************************************************************

`ifndef __SVDOC__
  /** Port interface */
  AHB_MASTER_IF master_if;
`endif

  /**
    @grouphdr ahb_generic_sys_config Generic configuration parameters
    This group contains generic attributes
    */

  /**
    @grouphdr ahb_master_slave_config Master and slave configuration
    This group contains attributes which are used to configure masters and slaves within the system
    */

  /**
    @grouphdr ahb_addr_map Address map
    This group contains attributes and methods which are used to configure address map
    */
   
   /**
   * Enumerated types that tells ERROR response handling policy for AHB Master.
   */
  typedef enum {
     CONTINUE_ON_ERROR = `SVT_AHB_CONFIGURATION_CONTINUE_ON_ERROR, /**< Master continues with the remaining transfers in a burst after receiving an ERROR response. This mode will not insert an IDLE during the second cycle of an ERROR response */
     CONTINUE_ON_ERROR_WITH_IDLE= `SVT_AHB_CONFIGURATION_CONTINUE_ON_ERROR_WITH_IDLE, /**< Master continues with the remaining transfers in a burst after receiving an ERROR response. This mode will insert an IDLE during the second cycle of an ERROR response.This mode is not yet supported */
     ABORT_ON_ERROR = `SVT_AHB_CONFIGURATION_ABORT_ON_ERROR, /**< Master will abort the burst after receiving an ERROR response. Master will not rebuild the transaction*/ 
     ABORT_ON_ERROR_WITH_REBUILD= `SVT_AHB_CONFIGURATION_ABORT_ON_ERROR_WITH_REBUILD /**< Master will abort the burst after receiving an ERROR response. Master will rebuild the transaction again from the beat which got an ERROR response.This mode is not yet supported*/
  } error_response_policy_enum;

  /** @cond PRIVATE */ 
  // This is made private due to known limitations. It should be made public once the STAR 9000993130 is fixed
  /** 
  *  Enumerated types that defines maximum address boundary limit for a given burst transfer.
  */
  typedef enum {
    ONE_KB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_1KB,
    TWO_KB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_2KB,
    FOUR_KB =            `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_4KB,
    EIGHT_KB =           `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_8KB,
    SIXTEEN_KB=          `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_16KB,
    THIRTY_TWO_KB=       `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_32KB,
    SIXTY_FOUR_KB=       `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_64KB,
    ONE_TWENTY_EIGHT_KB= `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_128KB,
    TWO_FIFTY_SIX_KB =   `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_256KB,
    FIVE_TWELVE_KB =     `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_512KB,
    
    ONE_MB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_1MB,
    TWO_MB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_2MB,
    FOUR_MB =            `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_4MB,
    EIGHT_MB =           `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_8MB,
    SIXTEEN_MB=          `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_16MB,
    THIRTY_TWO_MB=       `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_32MB,
    SIXTY_FOUR_MB=       `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_64MB,
    ONE_TWENTY_EIGHT_MB= `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_128MB,
    TWO_FIFTY_SIX_MB =   `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_256MB,
    FIVE_TWELVE_MB =     `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_512MB, 

    ONE_GB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_1GB,
    TWO_GB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_2GB,
    FOUR_GB =            `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_4GB
  } max_addr_boundary_limit_enum;

  /** @endcond */

`ifdef SVT_VMM_TECHNOLOGY  
   /**
    @grouphdr ahb_bus_sys_config Bus configuration
    This is not yet supported. <br>
    This group contains attributes which are used to configure bus within the system
    */
`else  
   /**
    @grouphdr ahb_bus_sys_config Bus configuration
    This group contains attributes which are used to configure bus within the system
    */
`endif  
  // ****************************************************************************
  // Public Data
  // ****************************************************************************

`ifndef __SVDOC__
  /** Modport providing the system view of the bus */
  AHB_IF ahb_if;
`endif

  /**
    * @groupname ahb_generic_sys_config
    * An id that is automatically assigned to this configuration based on the
    * instance number in the svt_ahb_system_configuration array in
    * svt_amba_system_configuration class.  Applicable when a system is created
    * using svt_amba_system_configuration and there are multiple ahb systems
    * This property is automaically set by VIP and must not be assigned by the
    * user.
    */ 
  int system_id = 0;

  /** 
    * @groupname ahb_clock
    * This parameter indicates whether a common clock should be used
    * for all the components in the system or not.
    * When set, a common clock supplied to the top level interface 
    * is used for all the masters, slaves and interconnect in 
    * the system. This mode is to be used if all components are
    * expected to run at the same frequency.
    * When not set, the user needs to supply a clock for each of the
    * port level interfaces. This mode is useful when some components
    * need to run at a different clock frequency from other
    * components in the system.
    */
  bit common_clock_mode = 1;

  /** 
    * @groupname reset
    * This parameter indicates whether a common reset should be used
    * for all the components in the system or not.
    * When set, a common reset supplied to the top level interface 
    * is used for all the masters, slaves and interconnect in 
    * the system. This mode is to be used if all components are
    * expected to use the same reset signal.
    * When not set, the user needs to supply a reset for each of the
    * port level interfaces. This mode is useful when some components
    * need to be reset at a different time from other
    * components in the system.
    */
  bit common_reset_mode = 1;
  
`ifdef SVT_VMM_TECHNOLOGY
  /**
   * Enables the Multi-Stream Scenario Generator
   * Configuration type: Static
   */
  bit ms_scenario_gen_enable = 0;

  /** 
   * The number of scenarios that the multi-stream generator should create.
   * Configuration type: Static
   */
  int stop_after_n_scenarios = -1;

  /** 
   * The number of instances that the multi-stream generators should create
   * Configuration type: Static
   */
  int stop_after_n_insts = -1;

  /** 
   * @groupname ahb_bus_sys_config
   * This is not yet supported. <br>
   * Determines if a VIP bus should be instantiated
   */
`else
  /** 
   * @groupname ahb_bus_sys_config
   * Determines if a VIP bus should be instantiated
   */
`endif
  bit use_bus = 0;


  /** @cond PRIVATE */ 
  // This is made private due to known limitations. It should be made public once the STAR 9000993130 is fixed
  /**
    * @groupname ahb_generic_sys_config 
    * Defines maximum address boundary limit for a given burst transfer in terms of 2's power.
    * Default value is ONE_KB=10 (here 10 indicates the 2's power ie 2^10=1024=1KB).User can define maximum value upto 4GB.
    * This feature is applicable to Active/Passive AHB Master and Slave Components 
    */
  max_addr_boundary_limit_enum max_addr_boundary_limit = ONE_KB;
  /** @endcond */

  /**
   * @groupname ahb_generic_sys_config
   * Enables system monitor
   */
  bit system_monitor_enable = 0;

  /**
    * @groupname ahb_generic_sys_config 
    * When set to '1', enables system level coverage.All covergroups enabled
    * by system_ahb_*_enable are created only if this bit is set.
    * Applicable if #system_monitor_enable=1
    * <b>type:</b> Static 
    */
  bit system_coverage_enable = 1;  

  /**
    * @groupname ahb_coverage_protocol_checks_system
    * Enables system level protocol checks coverage. 
    * <b>type:</b> Dynamic 
    */
  bit protocol_checks_coverage_enable= 0;

  /**
    * @groupname ahb_coverage_protocol_checks
    * When set to '1', enables coverage for system level positive protocol checks
    * When set to '1', enables positive protocol checks coverage.
    * When set to '0', enables negative protocol checks coverage.
    * <b>type:</b> Static 
    */
  bit pass_check_cov = 1;

  `ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to UVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to UVM_HIGH or below.
    */
  bit display_summary_report = 0;
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to OVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to OVM_HIGH or below.
    */
  bit display_summary_report = 0;
`else
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to NOTE or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to DEBUG or below. 
    */
  bit display_summary_report = 0;
`endif

`ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of performance summary report of transactions by the system env
    *
    * When set, performance summary report of transactions are printed by the system env
    * when verbosity is set to UVM_MEDIUM or below.
    *
    * When unset, performance summary report of transactions are printed by the system
    * env when verbosity is set to UVM_HIGH or above.
    */
  bit display_perf_summary_report= 0;
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of performance summary report of transactions by the system env
    *
    * When set, performance summary report of transactions are printed by the system env
    * when verbosity is set to OVM_MEDIUM or below.
    *
    * When unset, performance summary report of transactions are printed by the system
    * env when verbosity is set to OVM_HIGH or above.
    */
  bit display_perf_summary_report= 0;
`else
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of performance summary report of transactions by the system env 
    *
    * When set, performance summary report of transactions are printed by the system env 
    * when verbosity is set to NOTE or below.
    *
    * When unset, performance summary report of transactions are printed by the system
    * env when verbosity is set to DEBUG or above. 
    */
  bit display_perf_summary_report= 0;
`endif
    
  /**
   * @groupname ahb_master_slave_config
   * Used by the AHB monitor, master, and slave interfaces. When true, turns on the 
   * AHB Lite mode 
   * for AMBA AHB models. Lite mode has only one AHB Master and one or more AHB Slaves. 
   * It does not support SPLIT and RETRY.
  */
  bit ahb_lite = 0 ;

  /**
   * @groupname ahb_master_slave_config
   * When set to 1, enables AHB-3.0 features as per ARM IHI 0033A.
   * Applicable to Active and Passive Master and Slave
   * Configuration type: Static
  */
  bit ahb3 = 0 ;

  /**
   * @groupname ahb_master_slave_config
   * Used by the AHB monitor, master, and slave interfaces. 
   * AHB Lite MultiLayer Mode for AMBA AHB models. 
   * AHB Lite Multilayer mode has multiple AHB Lite Master and one or more AHB Slaves.
   * When set to '1', will enable connection of more than one AHB Lite Master in a Single System Env.
  */
  bit ahb_lite_multilayer = 0 ;
  
  /**
   * @groupname ahb_master_slave_config
   * Used by the AHB monitor, master, and slave interfaces. 
   * When set to '1', will enable AMBA 5 AHB protocol features as per ARM IHI ID102715
   * Applicable to Active and Passive Master and Slave
   * Configuration type: Static
  */
  bit ahb5 = 0 ;

  /**
   * @groupname ahb_master_slave_config
   * Used by the AHB monitor, master, and slave interfaces. 
   * When set to '1', will consider / drive the BUSY cycle only with HREADY
   * being HIGH for AHB3 / AHB5 mode
   * Applicable to Active and Passive Master and Slave
   * Configuration type: Static
  */
  bit count_busy_only_during_hready_high = 0 ;

  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------

  /** 
    * @groupname ahb_master_slave_config
    * Number of masters in the system 
    * - Min value: 1
    * - Max value: \`SVT_AHB_MAX_NUM_MASTERS
    * - Configuration type: Static 
    * .
    */
  rand int num_masters;

  /** 
    * @groupname ahb_master_slave_config
    * Number of slaves in the system 
    * - Min value: 1
    * - Max value: \`SVT_AHB_MAX_NUM_SLAVES
    * - Configuration type: Static
    * .
    */
  rand int num_slaves;

  /** 
    * @groupname ahb_master_slave_config
    * Array holding the configuration of all the masters in the system.
    * Size of the array is equal to svt_ahb_system_configuration::num_masters.
   */
  rand svt_ahb_master_configuration master_cfg[];

  /** 
    * @groupname ahb_master_slave_config
    * Array holding the configuration of all the slaves in the system.
    * Size of the array is equal to svt_ahb_system_configuration::num_slaves.
    */
  rand svt_ahb_slave_configuration slave_cfg[];

`ifdef SVT_VMM_TECHNOLOGY
   /** 
    * @groupname ahb_bus_sys_config
    * This is not yet supported. <br>
    * Holds configuration of the bus group in the system.
    */
`else
   /** 
    * @groupname ahb_bus_sys_config
    * Holds configuration of the bus ENV in the system.
    */
`endif  
  rand svt_ahb_bus_configuration bus_cfg;
 
  /**
    * @groupname ahb_addr_map
    * Address map for the slave components. This is used by system monitor for
    * performing system checks. This member is initialized through method
    * #set_addr_range.
    */
  svt_ahb_slave_addr_range slave_addr_ranges[];

   /**
    * @groupname ahb_addr_map
    * Enables mapping of two or more slaves to the same address range.  If two or more
    * slaves are mapped to the same address range through the set_addr_range
    * method and this bit is set, no warning is issued. Also, routing checks in
    * system monitor take into account the fact that a transaction initiated at
    * a master could be routed to any of these slaves.  A given address range
    * can be shared between multiple slaves, but the entire address range must
    * be shared. Note that this doesn't necessarily mean that the entire
    * address map of a slave needs to be shared with another slave. It only
    * means that an address range which lies within the address map of a slave
    * and which is shared with another slave, must be shared in its entirety
    * and not partially. This is possible because the set_addr_range method
    * allows the user to set multiple address ranges for the same slave. 
    * For example, consider two slaves S0 and S1, where S0's address map is
    * from 0-8K and S1's address map is from 4K-12K. The 4K-8K address range
    * overlaps between the two slaves.  The address map can be configured as
    * follows: <br>
    * set_addr_range(0,'h0,'h1000); //0-4K configured for slave 0 <br>
    * set_addr_range(0, 'h1001, 'h2000); //4K-8K configured for slave 0 <br>
    * set_addr_range(1, 'h1001, 'h2000); //4K-8K configured for slave 1 overlaps with slave 0 <br>
    * set_addr_range(1,'h20001, 'h3000); //8K-12K configured for slave 1. <br>
    *
    * Note that the VIP does not manage shared memory of slaves that have
    * overlapping addresses.  This needs to be managed by the testbench to
    * ensure that data integrity checks in the system monitor work correctly.
    * This can be done by passing the same instance of svt_mem from the
    * testbench to the slave agents that share memory. Refer to
    * tb_amba_svt_uvm_basic_sys example for usage. <br>
    *
    * If this bit is unset, a warning is issued when setting slaves with
    * overlapping addresses. In such a case, routing checks do not take into
    * account the fact that a transaction could be routed to any of these slaves
    * which may result in routing check failure. <br>
    *
    * Configuration type: Static 
    */
  rand bit allow_slaves_with_overlapping_addr = 0;

  /**
   * @groupname ahb_master_slave_config
   * Default value is 0.
   * Used by the AHB master, slave, and monitor interfaces. Used to disable HLOCK and HMASTLOCK
   * related checks when AHB locked transaction feature is not used in the design. When true,
   * HLOCK and HMASTLOCK related checks are disabled; when false, the checks are enabled.
   */
  bit disable_locked_transaction_support = 0;

  /**
   * @groupname ahb_master_slave_config
   * Default value is 1.
   * Used by the AHB master, slave, and monitor interfaces.  Sets bus endianness. When
   * false, the bus is treated as big endian; when true, the bus is treated as little
   * endian
   */
  rand bit little_endian = 1;

  /** 
    * @groupname ahb_generic_sys_config
    * Array of the masters that are participating in sequences to drive
    * transactions.   This property is used by virtual sequences to decide
    * which masters to drive traffic on.  An index in this array corresponds to
    * the index of the master in slave_cfg. A value of 1 indicates that the
    * master in that index is participating. A value of 0 indicates that the
    * master in that index is not participating. An empty array implies that
    * all masters are participating.
    */
   bit participating_masters[];

  /** 
   * @groupname ahb_generic_sys_config
   * Array of the slaves that are participating in sequences to drive
   * transactions.   This property is used by virtual sequences to decide
   * which slaves to drive traffic on.  An index in this array corresponds to
   * the index of the slave in slave_cfg. A value of 1 indicates that the
   * slave in that index is participating. A value of 0 indicates that the
   * slave in that index is not participating. An empty array implies that
   * all slaves are participating.
   */
   bit participating_slaves[];

  /**
   * @groupname ahb_generic_sys_config
   * Default value is 0.
   * Used by the AHB bus. Defines master number assigned as default master. <br>
   * The default master is granted the bus when none of the masters in the system
   * are requesting the access to the bus. Usually the bus master which is most 
   * likely to request the bus is made the default master.
   */
  rand int default_master = 0;

  
  /**
   * @groupname ahb_generic_sys_config
   * Default value is 0.
   * Used by the AHB bus. Master number assigned to be the dummy master. <br>
   * The Dummy Master is a built-in bus Master model that only performs IDLE
   * transfers. In the AHB Bus VIP, the Dummy Master is required. The Dummy 
   * Master is granted whenever there are no other Masters that can be granted 
   * to the System Bus. Following are the cases where the Arbiter must grant the 
   * System Bus to the Dummy Master: 
   * - When a Split response is given to a locked transfer 
   * - When a Split response is given and all other Masters have already been split
   * .
   * A Dummy master can also be the default master.
   */
  rand int dummy_master = 0;

  /**
   * @groupname ahb_generic_sys_config 
   * Defines the ERROR response handling policy for all the AHB Masters present
   * in the system, when svt_ahb_system_configuration::master_error_response_policy[]
   * is not programmed; that is when size of this array is zero. 
   * In such case, the setting of this attribute is applicable for all the masters. <br>
   * This configuration parameter supports the following values:
   * - ABORT_ON_ERROR (default) Abort transaction on receiving ERROR response.
   *   Master will not rebuild the transaction.
   * - CONTINUE_ON_ERROR Continues with the remaining transfers in a burst after 
   *   receiving an ERROR response. This mode will not insert an IDLE during the
   *   second cycle of an ERROR response.
   * .
   * This configuration parameter does not yet support the following values:
   * - CONTINUE_ON_ERROR_WITH_IDLE Continues with the remaining transfers in a 
   *   burst after receiving an ERROR response. This mode will insert an IDLE 
   *   during the second cycle of an ERROR response. 
   * - ABORT_ON_ERROR_WITH_REBUILD Abort the burst after receiving an ERROR 
   *   response. Master will rebuild the transaction again from the beat 
   *   which got an ERROR response.
   * .
   * Configuration Type: Static
   */
  rand error_response_policy_enum error_response_policy = ABORT_ON_ERROR;

  /**
   * @groupname ahb_generic_sys_config 
   * Defines the ERROR response handling policy for each of the AHB Masters present
   * in the system. <br>
   * Programming this array allows different masters in the system to have different
   * settings for error response policy. <br>
   * Note that when this array size is zero, the setting of
   * svt_ahb_system_configuration::error_response_policy will be used. <br>
   * Each element of this array supports the following settings:
   * - ABORT_ON_ERROR (default) Abort transaction on receiving ERROR response.
   *   Master will not rebuild the transaction.
   * - CONTINUE_ON_ERROR Continues with the remaining transfers in a burst after 
   *   receiving an ERROR response. This mode will not insert an IDLE during the
   *   second cycle of an ERROR response.
   * .
   * The following settings are not yet supported:
   * - CONTINUE_ON_ERROR_WITH_IDLE Continues with the remaining transfers in a 
   *   burst after receivin an ERROR response. This mode will insert an IDLE 
   *   during the second cycle of an ERROR response. 
   * - ABORT_ON_ERROR_WITH_REBUILD Abort the burst after receiving an ERROR 
   *   response. Master will rebuild the transaction again from the beat 
   *   which got an ERROR response.
   * .
   * Configuration Type: Static <br>
   * Usage: 
   * - Size the attribute to match to number of masters in the system:
   *   sys_cfg.master_error_response_policy = new[sys_cfg.num_masters];
   * - Program the error response policy settings for each of the masters:
   *   sys_cfg.master_error_response_policy[0] = svt_ahb_system_configuration::ABORT_ON_ERROR; <br>
   *   sys_cfg.master_error_response_policy[1] = svt_ahb_system_configuration::CONTINUE_ON_ERROR;
   * .
   * Note that this is used by master, slave and bus VIP components. So it is required
   * to program this attribute appropriately when different masters in the system needs
   * to have different error response policies. 
   * From slave VIP perspective, the indices of this array corresponds to hmaster signal 
   * value. For example, if the hmaster value is 8, slave VIP uses 
   * sys_cfg.master_error_response_policy[8] as the error response policy for transfers
   * with thi hmasner value. <br>
   * In cases where hmaster value does not correspond to  master index, this feature is 
   * not supported. In such case, user is expected to keep this array size as zero, and
   * program svt_ahb_system_configuration::error_response_policy.
   * 
   */
  error_response_policy_enum master_error_response_policy[];
   
  /**
   * @groupname ahb_generic_sys_config
   * Default value is -1.<br>
   * The Default Slave is selected when the address is not within any 
   * allocated region. For non-sequential and sequential transfers, 
   * the default slave provides a two-cycle ERROR response. For busy 
   * and idle transfers, the Default Slave provides a zero-wait state 
   * OKAY response.<br>
   * Used by the AHB System monitor:
   * - Set the default slave for the AHB system monitor (-1, 0 to 15). 
   * - The AHB system monitor will not perform the data integrity check
   *   for the transactions routed to default slave port.
   * - If set as -1:
   *   - The AHB System monitor assumes that the default slave 
   *     functionality is embedded within the bus DUT. 
   *   - The AHB system monitor will not perform slave address routing check
   *   on the default slave port.
   *   .
   * - If set to a value in the range 0 to 15:
   *   - The AHB system monitor will perform slave address routing check on
   *     the default slave port.
   *   .
   * .
   * Used by the AHB bus VIP:
   * - Sets the default Slave of the AHB system (0 to 15).
   * - Always the default slave functionality is embedded within the bus VIP.
   * - The AHB bus VIP does not sample any of the slave connected to the default
   *   slave port ID.
   * .
   */
  rand int default_slave = -1;
  
  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB System level check on Default Slave in the AHB System
    * - When set 1: Default Slave checks are turned on for default Slave.
    *   The default Slave may only respond to NSEQ or SEQ with an ERROR response.
    * - When not set (0), Default Slave checks are turned off.
    *   This is the default setting for this parameter.
    * .
    * <b>type:</b> Static
    */
  bit default_slave_resp_check = 0;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB System level check on Decoder in the AHB System
    * - When set 1: Decoder check for hsel to be asserted will be turned on.
    * - When not set (0), Decoder check for hsel to be asserted will be turned off.
    *   This is the default setting for this parameter.
    * .
    * <b>type:</b> Static
    */
  bit decoder_hsel_assert_check = 0;
  
  /**
   * Defines multiple slave select signal feature for each of AHB Slaves present in the system<b>
   * Programming this array for each of AHB Slaves present in the system to 1, will enable multiple HSEL signal<b>
   * By default, the multiple hsel signals are disabled for AHB BUS, Slave and Monitor Models.<b>
   * <b>type:</b> Static
   */
  bit multi_hsel_enable[];
  
  /**
   * Defines the width of AHB Slave Multiple HSEL signal for specific slave.
   * By default, HSEL signal width will be 1. User can control the width of HSEL signal for specific slave 
   * by setting this configuration parameter. 
   * This will enable the user to configure different widths for multiple HSEL signals of a particular Slave.
   * <b>type:</b> Static
   */
  int multi_hsel_width[];

   /** 
    * @groupname ahb_generic_sys_config
    * - When set to -1: There is no limit on the number of rebuild 
    *   attempts on RETRY response for a given transaction. 
    * - Default value: -1
    * - When set to a value greater than -1: Defines the maximum 
    *   number of rebuild attempts on RETRY response for a given 
    *   transaction. Once the number of RETRY responses on a given 
    *   transaction reaches this value, the transaction will be aborted.
    *   - svt_ahb_transaction::status is set to svt_ahb_transaction::ABORTED
    *   - svt_ahb_transaction::response_type is set to svt_ahb_transaction::RETRY
    *   - The info of RETRY responses received on the transaction can be 
    *     retrived by calling the method on the transaction object-- 
    *     svt_ahb_transaction::get_retry_response_info()
    *   .
    * - Max value: \`SVT_AHB_MAX_REBUILD_ATTEMPTS_ON_RETRY_RESP. This is user re-definable.
    * - Valid range: -1 to \`SVT_AHB_MAX_NUM_REBUILD_ATTEMPTS_ON_RETRY_RESP
    * - Configuration type: Static 
    * - Applicable to master and slave agents in both active & passive mode
    * .
    */
  rand int max_num_rebuild_attempts_on_retry_resp = -1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to check that the bus grant is 
    * given to all the master connected on the bus.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_all_masters_grant_enable = 1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to check that all Masters have 
    * requested for the bus at least once.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_all_masters_busreq_enable = 1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to verify which master is requesting
    * the bus and which master is getting the access of bus.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_cross_all_masters_busreq_grant_enable = 1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to verify all the slaves have been 
    * selected at least once.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_all_slaves_selected_enable = 1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to verify all the slaves have been 
    * selected at least once.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_slaves_selection_sequence_enable = 1;  
 
  /**
   * @groupname ahb_addr_map
   * Enables complex address mapping capabilities.
   * 
   * When this feature is enabled then the get_dest_slave_addr_from_global_addr(),
   * get_dest_global_addr_from_master_addr(), and get_slave_addr_range() methods
   * must be used to define the memory map for this AHB system.
   * 
   * When this feature is disabled then the set_addr_range and translate_address()
   * methods must be used to define the memory map for this AHB system.
   */
  bit enable_complex_memory_map = 0;

  /** @cond PRIVATE */  

`ifdef QUESTA
  /**
   * This workaround was put in place because Questa could not solve the nested
   * foreach loop constraint that is in reasonable_data_width (out of memory errors).
   */
  rand int questa_data_width;

  /**
   * This workaround was put in place because Questa could not solve the nested
   * foreach loop constraint that is in reasonable_data_width (out of memory errors).
   */
  rand int questa_log_base_2_data_width;
`endif

  /**
   * This workaround was put in place because INCISIV is unable to resolve the 
   * hierarchical access to field “num_bus_masters” through bus_cfg in the right
   * side of constraint.
   */
  rand int num_bus_masters;
  /**
   * This workaround was put in place because INCISIV is unable to resolve the 
   * hierarchical access to field “num_bus_slaves" through bus_cfg in the right
   * side of constraint.
   */
  rand int num_bus_slaves;

    /**
    * @groupname ahb_generic_sys_config
    * This variable specifies maximum address boundary limit for a burst transfer
    */
  int burst_boundary_limit = 'b1 << ONE_KB;

  /**
    * @groupname ahb_generic_sys_config
    * This variable is used for checking address boundary based on configured max_addr_boundary_limit.
    * Default value is 'b0011_1111_1111, which selects LSB 10 bits of addr ie addr[9:0] when ANDED with addr
    */
  bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] addr_sel_bits = 'b0011_1111_1111;
  

  /** @endcond */

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
TfqR7BshG8cAvyuh+HZYjkquWXpHYi+qqTeX8orxvG2IXyckTibuV5uHTtcuhB43
rAf3CjGjBgNx3hsi2SS1muH93IqDO6DduKFRi5X68Yrf/GAxtXFyU5j/cM3HUs2s
xs5hsfXQPibnU5OYNQgsBmTDRZ8824fEd9ErpLioMNQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 10029     )
383ZBYknshAlEKfqE6j9kpP3MjAJMeTJCLc6N0k5FJEfz2TuW1+z958e6hucS6YE
0HpgKef5J+LxSWQMZ0GyLkUbfHSYvha9lKGNM0hjW59QjmVhOeKVB5s5SWrDU+lR
aFf4kb4YsSsPrOCph1ZWBXi+fgwMiwGEGx1Rk9g09XzBZL5xc5Kr1fNmjwQsb8Ri
WFrbJREns3NT9o/GgaSYnXYAecK7o30qN+LZaGevf2kmtYFmpryfaEBUrVFWjXJA
8r1jNE9N9981UYhCLr7Ds8PcRohHDkDf2AdBoLNxYaASEpKnyXe5KwueosQklqHj
xma25MiE1LK7UdBvutCNnrzs0+f7HfYjDQ6IczGx9lfZH2qHKP9uy4BlcDZhoxNh
U3EjoDqlabnC9DIfCq2tdCGyxTnNURN0gdgrs4gqhSFo2BuW1HOYXeO68Z6uiZzl
Iz6rvmR7fePO3GZ5ZC9htOmluK9rZj1y5gED3msIEKXpglkobF7R4Xkv49wPhLhV
GKc9zHoPWe8gcNAxPA5HO+CHE6wuY1ir+iaUJt+RZP8OHktbcwU7Wy1oo+taAtEV
0KWMDj17QPp16W02b2l5V1ca/k4mNvUq77mHFzTzhTAyTKxo6/fkvytthvmIqsio
lT+/XKkA0EnbKxi+CvEMh2OD+8A44c6wCcn6Xz48jUPQbIF6rH3I7daQGt7cmOjW
/qRWiq6WlwsqECBd1yUe+L/bEIkQ/W6mw4r6Q1nNNOWTTQt4EGrah5XXeMghrIkc
ZtjTyiegLjq7rcPFdWzZCaWiTNd/9ymu/5IdCEcT/gmo856FjzQMsTCHu03GtLdu
1pG67grrYPbOajopcj3bAXop3esFR1jHzTgFr9tDCsBGlHaAkSIRdevymHGt6TJE
gRkzvm5CGrKinObbFuOeQZKxFwKKd0HO4N/9+jP2U0HyEfi0RhTfApuaUiuqXn1G
jpBW81njJF845LpcMnJHAi99pNqMbNWEw1kySv6raDBXZdLiYiKMLEHUoxG/oJtT
j2c2Y9pEEatZ2H8iQYpl8uPMXdaoBrF+843hgy5q5dM0ilZTBviusLjRtczFho/l
Ld7EkjEqjagWsTzWWispkzbOqDPKu2vDIOt1Mjnf5RG9/wecN7IQK/uqZ1B9l64L
WEZ2H0CfH+dxsJ8+2GNeqDtf7MtFw2bTpc3IzZtWwiEKK1bNfBdqjEad7jq3UXGy
guf4DC7Xc8MGZ44vLncHXws4oU7HbQnjbPz3jUFhcoCloGjQN75x9PGYaoNaD8ZF
AItV3UvQ7Kt5hmdG2EcYnIMowxBh0SdPCC/R5X7pUads5HradTm+LrueqA7bXl7e
pgDtXF9kyqr7/Zjw10z2fi4mEwp4fAeSwYpxN/86ZwMFaiwnxaAHClCLKnTBuixa
sSBgHFN4S8A2nGbEciuI5MoWF+8me4Grj0jXU8Zf5p4XaBoIlZlg9bIeiIVm3V4q
z7wfQ0R/EYnloohtRVGDOz2wDsypBstnXdVHuD/r++IlIVBsdRcxM8AUB2j8T4EO
5vcUmxaJua9vxrF4UgCylG3QQUyTMhZ0WIoqc2SC7iAtRjRNkPkAHa/C7mqkEjVV
D7b7Ky2EBzHQkRFbR2maiNPDLUzGED7LbOujqb6eQG45lsmQvD4yVrGCsuaLJYvz
MDzHXGBtfHnTkhLTQwjdZBBm1hHE10+jm6KxZ/bNSFk3MvQxCHeHJ42LvHEZm7EM
mYwNNeStRs/1cbyEIO/9jC1KQlX3/5ruI+xXpQlgtQKoCX+G+sQIDE2T7q7NpqEM
QnWg3z/gofmo609GUiJp8HbCLhtx1RT4bC4oIe19EHNOKpYiFFJeg4gzYey8oxpJ
57eyPMKKkxPqWsJ1zDykqXMf7T0LXDi5qYXUkMumzR038JXW1vrBQFoxRgvwyknL
+Qfm00fP13/K9GO7iYVra5AKl7nHqHkucajSozF+U9wMTfvZeTY3fz9OorPianS2
KI2fPP47AJMnCL2VVElPSsFo7E9otWT9XtaPFOC2zXKPBxwebr6l7LfwliB42S+U
f6X6PVV9W9MED3yNkT8C1zul3LBoDhqWHCj2CoU5J8oIj/he6QAypzD2c2HYQrbj
4FzRFA/2Yo1s/MJ7jBFs2EGau4g9gOTFy3lJimdwNxxtKYiBrXMVPhmotyizQp2+
bcMyoavOy0tBpT3D83Jb/C5wMYfIG6PAHGFzjnT2OrX9ersB9Tmnu7tqI984ctrE
e8Mkjb+n83/J7/C2rbhi3NpzJsxhQHb7/c1PrpOsQ1I8WJwMEmZRy5OappsIq4S4
ezKwZYr1SK5S1hYvTE60m3NmeBwDr+yeti8kJrM0NEaQs7qaEtufsjskCt2AW9Kt
ebP+T5dmIciw5oZYafOc/nl0Futwcvl6lnodVRL/ubFZuZeh/8MZ5WMyfMIkwmpL
JpeaLkLmB2OrZU8rdvAzoKp27wrHMWKSUwqbkteh5UJYx+YT9RKnfMBjR3sjSVYh
cJQPu3NFs630/7KDmML9iGPJrzpON/Y+Fm+X8v6vj+2wtAfrTl99jOu65SS35Kot
LDU8TLyXGRm+m4SuwTSAIW5Hfg703JWoJp3ennDyk1EgJmif5dR9KE7ol9+FCxW5
04e95fYMsjQdJKdeZDco20e4F8X3xDTj5MmUxQ2Pm18442Zi+/bA8mVltFpv3uaX
cycPDm+geJXkGXxtZV+nT1P2awZtCv69ztOl2QLJycFSyZUPeoZuS/v2XTgiJ6NC
PYmrJL7a2pd3bjTbe4i2XyiOHpt3r/+6OddlKuK/Yyn7yZfrxsPnrYoOxFBsgsWy
HIMnu0DeW9Fkw0IGefWLu4JnTVZ+wC5hC4hWCUnrElx6OmrU48PNhJA0pclFBPSV
2dg5ACqZsG2XTBvLL8Ha/ohFpQ7+EwAj6PRAOkcvkdtjw9qkUNOS8szDhlkk/bqZ
JvoA65LEEizmS6/mKUxZSa+r0EfyKtyZwevUmUXYIeFeSAyTXr6T+E8R9vlqAYZE
iQW/f5HXx1s6qO5aJKBuyfOGkX6yha+pDsCFwM9F3c9yArM3avlfBqE3pB2WzFC5
bRj36LhJYOm4SY+f/3Yo08LyuBYgIGO1Q6+6EPZYeI/5hZ6V8C7T/quYX8ddQPag
CWV9pjSPYE8ZLxhVS4/lRplRGCCqwopXybIHZD3ND5q9h5mBnyYZ6MYJWJvnlgb8
HxhfF30gT8uvw5ndwlroDN/jDOlWPGbBQjASXZ+wd9zOBOuISe8aWD5s0KJe1vJo
5/yGGtr5k6odbFDEu/OJ/8wX2PBitBzmGKYBPAISsf5vVqxCv9C/DPPuMPbzlG5G
NltjHVl2TZwQHntgVencrmsstdzg1agBIr9oxu/xAV7JMuOFiM77ciwhWf/d3WVb
7+cJIu84P0BokTIinQ2yJLjaqFC22xutXROWx2yKKqyEgHvpW10CvS6VHI/bNs3x
BrG0y2+zOUkhz6swInAk8Qpdw8yCAsv6sWVBhwSi3PPwAObH1iymbGeC7dEir86Q
xz/BKCqOudvYxtXo2S07SSdOKq8szq6xga9ZyfxPQOnQlXWz4uu8F4X0LPq3mp8S
3aTrY6gSCUfjg8FMOi+AigfR7N+9CCnYafZ9y7B0OZ5Lm9xplZEJZ3I4sEdbyT1B
WK+U8WlpZi1PGVg2javrWiOeDM58b6cvfGLgUTSYoJiojejEKsUfFi6gsNfLo/rH
CdtYExI7VmLJFJIDM4Cr6cUta/7AqLD6mdUomvLxChGVaNBML5fo25Pzp1OE2w/Y
dCOO90wcgX6idCoA+nZ1ZdVjwfoBv0kEudI7E40DHOw8HURvx45E2kYrYNop57xD
cGgz5aak1ZuEgaCvEoE7m7jHshfkleHKeA8nsQtV9WZYWIwgXGbcvhR7kzesM5eS
S1X6BOuENJQ90bKAAS+Hx0atdkzcNzTYMLZf9eYQ/VDYh1YCDJm9XLrcOxzGoJPV
WD0hDMJzqntbqnXCWpM2sN8DmjGdSjpmmyLyGKLFWQPZUN+D6buR3m/Je8/Q9j0T
QNz1qS+DV7TD53QbmHNjypkxZwOFZqd9DdYZdZz4q8I74T8Y4ujUYVGgkceQEZ26
A3qQ3TaUMu1Yjatx9ZLnMjR3DrbQrPYq7ujKxsSHDZnTHQjkLgwDqalJKxdT7qBt
fb6o/xthZWY9WtuK5HEXPMnxtFJukMm7B8/+m7oLmm/kLVo/CaMqiqdASgVexRuy
p2J+f1c4oyXxbsqDlcAyZVp4mZkGjQBitXCYXhwyEYUt5ZsOsUSekEDwm1sjZhyJ
pjtVCq52+gDM135kBQsHBgKFWU+uDyMtZWuCRe6o3FsAVLb0BiQJ++aUy+d8ixf9
3CIcWbkanMLYVMbo5d6CIcsx84qgYfRmfZ/gOJaTFDG0K6fu1tEXKvqHRcgdVbiY
HE/zUbHP+v9z4qPnH2623d5axhDri15OlbtIj4ohSvX3dR9usHxRjbHOf3cYtw+O
K7WcOGeEloMWpeyXH/BKRfNGv/f25+0L/X8i5F9lJl6Hl7zblfY339ZOcjB3X+gW
LohSx8/sWrilwMbbC3XmYhxV+fEgC/yKmWaWM/i617NxvDTh42+3NDnrH7WRzIZy
ledEVOvT+WfCwN5NqHsUOIN4Uvr/42nXC8/0rV7xrPJ8r/LMLSu3CXTWtx3iPbQN
B+TBWB5MHiJjWXCgl1ekOS+3ccFm55XM+TJxqIt33GaDSfTN1j7ZW7oYbBsBxf/B
q8c9SK7wV3hVOazvvD5ZNp6BaZo8rDUBc5gLNQNOfoZ+zW+AIEvHsyoboG3VVA1+
E+cEe7FE6DxBkUHucPJevfKN5Z/kwPVsTYX4J/cTXpzFiV1hH4nhwJVcLQ5X9o5y
sKd1XGkphHGN20r81AZK+RkO0nV6IzwK9ers6bbvb4ZDTVOnDmGTbcX6DnRQmdiZ
oNkhnLa1lI1t5QslG43PR1nWtg4Or2zqQ2UTYageL5Njme/zJBp+DVSYKrDkoO3A
nkGsUsEhRgSvslrOKvFFSbpHJeWYfB39Qs6VMu9eGhstjF7m+lOqQr2f1jfA5E97
eCoBf45NuwU7vwbvArYYDcAZg693ogiZlHGa6kGibXOVbYSHyujRSufVqV6h2vHI
KvnRyhYSUWxGSEohJy1tkPlWL4wXWGhkkB47qhpqWMzwqWEzzpz5EGbMWir8pW1k
TOYNcDq3VlFl9AvS46TX0ntE7yZ9i+m6Bn+H5j8NQWWOpN2Geu+j+ezeRnoEndFV
ciJh6ukSpChx8+qIC95uyk7ElYYjp/ayt1vxsnVaf2sYLIgig/5ntj7Y4LzEtr5O
e28j9n6/gf7YRobtDc/rEMeHj3xTiH+TIfHdzpe28j9g1M4lpQ6PSVdd1amZPH/e
9H2YjdkDidvGJJwj6b/n39S84uOS+QtzMZ/ZqE+z+yVSG1m+ySqWoxzcYspDTg2s
j/oKR3dfz/oz1CAS1gDJ9Z4F7WUSZ/Ci2N7i43nlV4IpvQ9Pq5T5yXVZYJyC8hzC
Er1ubeM33cIdReDHL6quoe7b4vjXrs3LyBdVnjyQMMLp2Z5BcIKB3kXcEd4wFoW7
uy4OiBlokP1A9MWwguKy9RMyAe0vaKfZPoNk7OixAXpjD8UXS9McISKrA86RqQG0
ypEB2EGKdst6C7aDONnABk0oRs9jkwMwEIQWJ5ULp8bpLPdQp90sStUOg7DSsxiD
TFLijkayvUDAAnLI3Oe8Glff8ZAlecYLhCIv1IurrUyr0gQcukRZXqvk96byoE+M
SiERkfZiMHa71qCkVAhTtPChsLEH1mcDW66NCCArHVMJDQicSR7XpeHxiPZNWTGv
KYth4DMM580QG68fG65kC9iMJgN1PERxDid2ZNiH98NgRwWorW7CsNof3sfP2v4n
fIuNtMq22Ux8zP6mtJ5pDt37ky2ZayLEUHTTc1VG6IRri09o1CJZmwix+UzXZN48
gSNibfcAYFm4/DUclCeWQN7FdAZjPCPZJGaFMDE9Gob2azhP4QRgTGVRoisTvD3t
LI6iaR0jsXiCGs3WD5/A9aPag9+oyn36CSp2GDnm/eeG2rmYxv+3eO+4nkFDHUH1
YA8HPG2MEWYmzDMolhW1tPybDSX9E+SP/c+rKC1dSPGuKBBGyovLqboX6YK/aitc
YXS5FiToECJ8c+VEJUDTnqZsgp0+zblpvB+JldMsH81vgwu7fWPcLbqfhZJ42p9Q
wfyeTSAHt4u2DFEXqDJTotAS8QkIV1hQMBEAzbtLzYv6f6yns0o0Yt3JY4uVRPDM
smL02WNt9pncQG/CJxcTCE/pvSrQ0lpW0ymU6h23RzKmHy1TYYB43zA2kdOttnuL
sM+g0uc0/oIHTlyj+ZyxKfBM/Y9kOEueTbOStnkLKfRqUhCwBlBx5RoQRg+0CDdF
Q9LCsghkJ7aOUZRyChI0QsAHaPh23Ruc72cTVPxYKO8w7nYDaMH6FtzEHY40W+7q
VDROSHWTFK5xezJH0MBQVOnAnoxpu7/ZHzGPLQulgxFsq4gv97YfaVyMYjTMHe+/
LTJBdWoPWZ7FKDKKRfjq1Q2/uKP7yebLgasv/m2Bb9dKSiwvvv1Rzl4AEmRLhGn8
lrikYVcNhtUlpneDOKC01QsBKVXVfCeMmZdsnE9sFvn3YMIsdU/v93tkZYpqZ1m1
eLfYvrRLTp0f33Ai4vbB+SX1QctkfH8t3gIG4BpoPbVjmhZpBOUNNOnZjlJt+5W1
OQl6g6em2WjRCikOwQM3pFkSh4VD1zDAhP84aGgdCYcTxasj70malNpqD36Oxojl
1clOAHVWrsoOmf+wP/IlFuJwEAxxKvlQUxvRaZi7oohvRxADfex96Yhric1yTbZ8
H5EQmF1oZjX7ug38rP+u5qdLn5EdVFy63rxiWkZ4R/qx+jQxSi1/WbAc+bragH3N
sfEw5kKaLigOa7z0xlO6zEkffRfIzcX9u++i1sGMHUo+tyNKfmYROwNf4Bntns5n
irZWqPHI08mfBLK6XDgXHk3HBFsbGdWJez46uPxQto7d1bzXqo8f3RCW297Fh8B4
v6ErIMoToBMpjGJAxIR5Wi27KRBOMEyTIBY18l3werGubUaPsGisdFn8aViGqz20
uHjqbaWRm4Mp6jHF9P5vFB2S/JhbNORgVxW8UtVf+mImZVY4Lpsfisg7V4mjH/E1
osN+Dhacd5DjjV+gVTtiMOSGoPF+w4f/A1hhBK6NjOurYHSmWDKanqH87V5g2oAU
7GarxwrSiITe3l6iB9lFC2gnLw/qYY1GRpNyLOPDfaPuNy4oVwA0+LMgJgRYZStL
of+eJjIoSCHptrMowNY8eb48AFrxbwV5/ts7AmrScnT80bkD17mOEGkjljr+qokM
mH/M9F9BXSCURrMWPqGvboJ5BIeD+yQ1mjx9uRx1fbj4PxP1H5yaCgzPN4F1TfHU
wmrtwcIL3DSgKWVwkV1Zn/LYdP9LFvvDbTc+tOoN93ApCK+6U+wXliG3DlPfvbF8
Ec0ZbfXL3zGgfqVhgOG8LeUpZhIuXYd4vMwwT0L1N3eP7WZ/XGkJFZ/Hx9pgESZn
FtbL1JDVbZN1EcN1ljj5XzXOv7EVZPGDhK/37CtIJjBPRM1aAAIhMS5uZL2gqWhV
ykqKIdikn3Wsc6FpTf+J6JkgiQIN8ZypQN3+6OPTDKSd9jEU9pXQ7+Lgbe/gH14Z
HVQ2/ayGRNvjFbfWdTB1LqmCnDUhsOp91HawvYINYtY8MinEcZW17INyRr8Y730E
ICSxGJh+Nfj7nFswiO6+ZWXre3X1s/Jv9UaJt73M9+WvNu8kqUpOxNSIKfskRhRI
12FETNlc1z5KGMXzN+lyN3BoRsXeHuOsTft0TW64MDFSLs4ve3SzkPZkdsFtvhiG
uYeQfH7x4J98BbVk35wGUiYU+T01+YYJqgT/rDW7OWljsnIfmEwrbQnmefVoJYu4
PW04Voczc3VhHbbaaAibUrhfzdlQ64ZQoAfOPrQAM1+0BuMPWkOnKRD7KYX56wxV
Ovy6DjcuHBJyAGAfTjNHcA1IhHPqndZw5YW7KvDrqJgqPtdNWUKY9gjOsnWO3klG
j2CC5Pq8v1aIStxitMzDDPUjiXJx+btSoGzgsQr5wKp2tFS6OQYuxw4n7qHf+9Yo
r3MG9Dz4u5mM4xszG5IuTVSLr5pzTqmr8P8kykwFj1m0AS0c8KPZYSEY3TZUiSRT
abMKGiSOqJnWwV4oLiNY4y26cc66QOVoB2/Ziba8AYKDh/WoK4cHycbvMPsWeFQH
XO6wfbBsa1748cey48Sd0rYphTrMHXOGOBveEVOXjs3ROj6AXtFr5UpGlr/mWsOc
KjQLNNckqkNLoaq9ubn3i+xGNYsSn5J4tL9qOMLI0nd8JTUYr2uf4tdOqQ/DSYx5
/lUWz/ijuLsQApVJxp9dyLPj3Lmlc8L8iBv+Z9YGD8UC24kqaO3dPmFRGAi5AsWB
3Lf1GMawTvegIABzqA/1uRdH+fFXbvR6jl+zfMylJJThhqboiC5fNhRy099c6TIp
9aYCJnGPmN68jAW1yW7Vq92ZQ4cUbzBTrIxavQSJzEhhGHeJXLmSD299jQAaPP2L
3KbRVAyeokF03oA2kdtd2zm1LsmM5jayFEDXV/bUGpG8Vi+mvw8bMNIFbn/ZdolG
8QfDmStSk1CUYL8bBKzSkUuaGkjio4KFQffFO+WrkiV5ruioLlg+tb6hWx9AGUHI
5Qnfb1qG3Dq8p8WykKzFkTgZ+38CuNTETyLe9/LfqDvdu5+ybbsYVKrLE2m8b9ko
RZyyAQSZvZSbM7hj7ClIcA76bWfFsbLbAkT1KFGK3c4aEJyx1q7Matg5n5x10gdP
sSRQd/LKehtV6RHEhHZUFSEUu4cdfeyjiDQaTWeWHrXeH+nQpTiZHL774QNMU5nK
fv6pVYI6ql9Q0Y2g1MlF+l0SSDVO8F4oY3HusqHliIRYFzLU7wjop9URbUknNy+4
bEIwrdTaP2k/8KiWp6QZ880TFAFI5nkNoyRdYUfEmlU4Kff3RIUVZLVJCGO/6HK2
SQ1dNwaIPNoUMdXd7KmogVWKzof3nd1YZbgPEmwpFLDhUuwJvXsVUHkzlKK99GOF
POicIKJiCcyxad4fpmtp9gAzTByNiXqBjYmjjur1OBT7a3N965cEKxVE2yqzVKKj
E0elVMZxl4Vp08Zx/iLxc2VAKWJQHLld2ncKxlDSypa5DjIDMBrjtNJMmaVAzN6T
9nTr/2r6HWHTGXcX/RBdaxzQ6lXcWfbtLI+SQmHNraCOCMfb7E1kTTBdPO8oR7m5
hEF6ZLLc/PnP4/TILjLu1ECo1dpdTYNGUzECDvwj6+3Y0DHesxcYXSP1hQ2TBCE8
RuT5DCVV8d1Xm05twabYQr8T8+X11k+Q0WvSKuzzECetbAOpHlIKw2hudCFC1txI
HxpEeNSzSy0FCzwqbLuJucRBakrhCjtowTDJakXOdJ4Vq87JaTVH3fzh0abGUbFT
JW3kRdAaBtmMttqAgP2G0Ys4MzYjJX71yb+8TiXnISrFmpQdv6LEvIIip1sbXUSv
D37ziGfSWAYDWTw4/PsbYHL+KO8/7FIJ7hklNHa7md+SrM6P3olpS9dhWS8VIkff
42yZJSH0A8pleR+l/hAPKSuUmZrRAL65gCZOAkdS5OAy0KP2sciWSP0lH00YBcMC
vG51zbI2oca3cJoOC2YVoGwdwJV7gcx6tBoh+4tyrVzP+HQQMgpoU0a6vI4FBckB
qb596bSscXuJ9eji9py+Dk8zBefQBydWqW4kJHPO4GYgsHHdwxRdNj8mIPu1MMqO
7RO7HPGiF49siAGdbhT06rrNMj9v7dZSDQMUZXibMp3Gi9C5qSjCWdGcB3/C9kC1
4kwxIregj7Q++JPR66COTmpy28rAQ6w8HEEU2+1xDcPcu0MLNTpiDpdE0otWaccu
mlcOV/1C7viomD3J50DUhvazlMGbbQs/A1Bf6E2s/fguwSqzJKLoFKF6Eouv8h/K
dCNdJGaxDWEs1MAJfuXzASpOBdOlZE4UCYgumJ4VK2NSF0lOYLfZuX5mj9+qtsxK
2IlKA+q6cL7gEy2F92Sk1l0436hBylNFm7ta+gTAxKonHSxLFuNwmuTJ+4ee+fYs
AFoEpkMHad68nBa8CHm4mhLSXRHH7TbGimAGtpWrZ8DbUbskty84ATbmxS5L41mr
lvhiBgJZ4dzgi+IdZ9YlSiUh96FLHqWL63q/nFAVxTkmbfIu8hgFWr3OfpHeuu7s
NSZOEjnGri0JcSilpNuXiX1kC8w0WM3VQMVoX6/aP1Do/Y5tQjTYOb4ti/5qo5UI
CX/A/1e6t3hF5/SzUzQpACoSd/yPvyILQ1IlW6UIYaNtCJpwBHxZG8atK7OiEwlC
700fIv1ptSe70y0pWmKQzewz4cmGmnPrGvyVbtG0M7CjXQQ80SfiB7kdoyO1jJ2s
KfvZyxqRk/UZ2cqKHgMZzno6XjUjp39Ul1MnkhaSiS8Et2B9iohaQHb/jDB8GpGt
z21aPwkjltrvjfdQrlOOpLnX1rVyzZgQjOuFxUAdiU4gFDU0yS7XBhpIGOPr9GwS
uF+D3QSzcSimIT3E3LzSgemKVYbMKGKqYfCxH5cBjMHyjG4AEzHGjP1LU+M3u1+y
1XAGSferDz4aYgcwkaSZ12jgUdMakTx7P5Y7mcWn7/SBxfrEspoVueHxwH+i1hKm
edIW8gcHPOUkeJTsc84jvNjk5wugFfLhXq4FxbDJb302fxAlEXD98IJRAGS3YZ7D
oUKp99pmCZ9sTTjM9Qx5gGtEdHkPO76k/TZPSuMtojNuVTD4ZHDMpdMYAmobuiEP
bDhdclF5sBDkKO9CXCojPIgy5Wsb8JmSUQFpb9GfBZjzadsd46T98dOQGomYfeWl
Ft/JugH9TYLrC3fGEV50Z2Dqawj3obE7Lm+Dxv7ev1Hh/I4Y5cMShL/gXsDD5BJJ
kPApIcxNOzfLAnXCUJP5a6NfFYVr8OhNuBtsA/XlwsK38lhMAx1O3rHAx4RU/0s0
UE/Y1/K6+u17gWSQ3mQ+JGj1IBjipYnGcE/xU9UEpdmQu3mJ70e951pqg3mjtK14
7hSYTEZ2G/Ur2sT0iwiSHzlE/8NUtkNNy0KWArodvojuMabzBLwPu0wgJFJGaT+O
h+EHmK4j47hFJyKYUy6V1j/bDdqD8oP3KZOBEWMoJmf6L631Bn07H5YXCC2CZWHN
+wRK/o1tdggZZmgFiwUR3v3B93yFehvlMdoTNno1gudQCx0JXZJ/h9PdtOqAq4Dw
LcUaBrPtZzB41H8bDYlrgecUx2cBZOrSACwjzfQvcG9XLkJ5fWzweWkVJ7vuCMs5
ga0xAUTAV0tAREYUbcVl4YNYNOHiPf7cfNrcnL1JhEfAWqsU3mCN+pmzfBLpQi+j
8C5azy1G3iyl0u8Jl4rSPYpKwKexkX5slqRQfeOJ6EVOEMEH7mvMdtcChaE10JSM
QuD1PtQXUQTHD7+2u1hsVOQaC/EIF1dAAwGoZBzF3NCCuhbDt79xAncWm/y1rTU/
2t7jnjlD7/MRFBPgE3+A1dDpBQIk1kEzkdw1FP1Fc/jwO1xEW7dLkO9+SUDLdjSE
BRlICcpNpIfZ9xeRN0Vp9yyHJFkoBPqWg0YrfWrgUKJbsB1+OqNerCCLG/i/7u5O
PjUNelr2vizkch6j/1AKtDJYLk0I6iGuLtWwDOKxy1A+Jz4mUu4WlOAYbs64KY79
cPZ01mZEzEuYg/2jvs29Tr+rDLEruPlE/JZ0LB8Jgl1ut+aF6jReBabS38jbuI/V
LSVh/HawALJ3GdSeuks5X0IUhVsI4K80wsYH6MYY5VXWj3JK4YoMJs9xEBQlEmO/
t2ji0TZSkPDI+iVQmTjcSTNfE22lKDRx1njnyh5//5brCUj6vE+ig0/TWtrnRtUn
bw/dX2v67UKIsN1G+FN4iAl5tUC0EqRgz8ISbkydYnQZGAcVOVajzFSe8Fl0Odn+
`pragma protect end_protected  

  //----------------------------------------------------------------------------
`ifdef SVT_VMM_TECHNOLOGY
`svt_vmm_data_new(svt_ahb_system_configuration);
  /**
   * CONSTUCTOR: Create a new configuration instance, passing the appropriate argument
   * values to the parent class.
   */
   extern function new (vmm_log log = null, AHB_IF ahb_if=null);
`else
  /**
   * CONSTUCTOR: Create a new configuration instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the configuration
   */
   extern function new (string name = "svt_ahb_system_configuration",AHB_IF ahb_if=null);
`endif

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following:
   * 1) Allocate master and slave configuration object arrays
   */
  extern function void pre_randomize ();

  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************
  `svt_data_member_begin(svt_ahb_system_configuration)
    `svt_field_object(bus_cfg,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_int(system_id, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(common_clock_mode, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(common_reset_mode, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
  `ifdef SVT_VMM_TECHNOLOGY
    `svt_field_int(ms_scenario_gen_enable, `SVT_ALL_ON|`SVT_NOCOPY|`SVT_BIN)
    `svt_field_int(stop_after_n_scenarios, `SVT_ALL_ON|`SVT_NOCOPY|`SVT_DEC)
    `svt_field_int(stop_after_n_insts, `SVT_ALL_ON|`SVT_NOCOPY|`SVT_DEC)
  `endif
    `svt_field_int(num_masters, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(num_slaves, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_array_int (participating_masters, `SVT_NOCOPY|`SVT_HEX|`SVT_ALL_ON)
    `svt_field_array_int (participating_slaves, `SVT_NOCOPY|`SVT_HEX|`SVT_ALL_ON)

    `svt_field_int(use_bus, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(ahb3, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(ahb5, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(count_busy_only_during_hready_high, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(ahb_lite, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(ahb_lite_multilayer, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(allow_slaves_with_overlapping_addr, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(disable_locked_transaction_support, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(little_endian, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(default_master, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(dummy_master, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(default_slave, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_enum(error_response_policy_enum, error_response_policy, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_array_enum(error_response_policy_enum, master_error_response_policy, `SVT_ALL_ON|`SVT_NOCOPY)
    `svt_field_int(default_slave_resp_check, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(decoder_hsel_assert_check, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(max_num_rebuild_attempts_on_retry_resp, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(system_monitor_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_coverage_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_all_masters_grant_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_all_masters_busreq_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_cross_all_masters_busreq_grant_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_all_slaves_selected_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_slaves_selection_sequence_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(protocol_checks_coverage_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(pass_check_cov, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(display_summary_report, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(display_perf_summary_report, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_array_object(master_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(slave_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(slave_addr_ranges, `SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_int(enable_complex_memory_map, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_array_int(multi_hsel_enable, `SVT_ALL_ON| `SVT_BIN|`SVT_NOCOPY)
    `svt_field_array_int(multi_hsel_width, `SVT_ALL_ON| `SVT_DEC|`SVT_NOCOPY)
  `svt_data_member_end(svt_ahb_system_configuration)

  /** @cond PRIVATE */
  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();
  /** @endcond */

  /**
   * Assigns a system interface to this configuration.
   *
   * @param ahb_if Interface for the AHB system
   */
  extern function void set_if(AHB_IF ahb_if);
  //----------------------------------------------------------------------------
  /**
    * Allocates the master and slave configurations before a user sets the
    * parameters.  This function is to be called if (and before) the user sets
    * the configuration parameters by setting each parameter individually and
    * not by randomizing the system configuration. 
    */
  extern function void create_sub_cfgs(int num_masters = 1, int num_slaves = 1, int num_bus_masters = 0, int num_bus_slaves = 0);
  //----------------------------------------------------------------------------
  extern function int get_num_masters();
  //----------------------------------------------------------------------------
  extern function int get_num_slaves();

 /**
   * The method indicates if a given master's index is participating
   * based on the contents of pariticipating_masters array. 
   * @param master_index Master index. Corresponds to the index in master_cfg[] array 
   * @return Indicates if given master index is participating
   */
 extern function bit is_participating(int master_index);

 /**
   * The method indicates if a given slave's index is participating
   * based on the contents of pariticipating_slaves array. 
   * @param slave_index Slave index. Corresponds to the index in slave_cfg[] array. 
   * @return Indicates if given slave index is participating
   */
 extern function bit is_participating_slave(int slave_index);
 

  /** @cond PRIVATE */
  //----------------------------------------------------------------------------

 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);


  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static 
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);

  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif
  /** @endcond */

  //----------------------------------------------------------------------------
  /** Used to turn static config param randomization on/off as a block. */
  extern virtual function int static_rand_mode ( bit on_off ); 

  /** @cond PRIVATE */
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );
  /** @endcond */
  //----------------------------------------------------------------------------
  /**
    * Method to turn reasonable constraints on/off as a block.
    */
  extern virtual function int reasonable_constraint_mode ( bit on_off );

  /** @cond PRIVATE */
  /** Does a basic validation of this configuration object. */
  extern virtual function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);
  // ---------------------------------------------------------------------------

  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);

  //----------------------------------------------------------------------------
  /**
   * Simple utility used to convert string property value representation into its
   * equivalent 'bit [1023:0]' property value representation. Extended to support
   * encoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit encode_prop_val(string prop_name, string prop_val_string, ref bit [1023:0] prop_val,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);

  //----------------------------------------------------------------------------
  /**
   * Simple utility used to convert 'bit [1023:0]' property value representation
   * into its equivalent string property value representation. Extended to support
   * decoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit decode_prop_val(string prop_name, bit [1023:0] prop_val, ref string prop_val_string,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);
  
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern allocate_pattern();

  /** Gets the slave port corresponding to the address provided */
  extern function void get_slave_route_port(bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0]
          addr, output int slave_port_id, output int range_matched, output bit is_register_addr_space, output bit is_default_slave, input bit quiet_mode = 1);
  
  /** Gets the HSEL index of slave port corresponding to the address provided */
  extern function void get_slave_hsel_idx(bit[`SVT_AHB_MAX_ADDR_WIDTH -1:0] addr, output int hsel_id, input int slv_idx);

  /** 
    * @groupname addr_map
    * Virtual function that is used by the interconnect VIP and system monitor
    * to get a translated address. The default implementation of this function
    * is empty; no translation is performed unless the user implements this
    * function in a derived class. 
    *
    * Interconnect VIP: If the interconnect VIP needs to map an address received
    * from a master to a different address to the slave, the address translation
    * function should be provided by the user in this function. By default, the
    * interconnect VIP does not perform address translation.  
    *
    * System Monitor: The system monitor uses this function to get the
    * translated address while performing system level checks to a given
    * address. 
    *
    * Note that the system address map as defined in the #slave_addr_ranges is
    * based on the actual physical address, that is, the address after
    * translation, if any.  
    * @param addr The address to be translated.  
    * @return The translated address.
    */
  extern virtual function bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] translate_address(bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] addr);
  /** @endcond */

  /** 
    * @groupname ahb_addr_map
    * Set the address range for a specified slave.
    *
    * @param slv_idx Slave index for which address range is to be specified.
    * Index for Nth slave is specified by (N-1), starting at 0. If a value of -1
    * is passed, it indicates that the given address range refers to the address
    * space of the registers in the interconnect. The data integrity system
    * check does not perform checks on configuration transactions which are
    * targeted to registers within the interconnect, as these transactions are
    * not targeted to external memory.
    *
    * @param start_addr Start address of the address range<b>
    *
    * @param end_addr End address of the address range<b>
    * User can configure multiple address ranges for a single Slave as below <b>
    * Example: consider following address ranges defined for 2 slaves in a system<b>
    * set_addr_range(1,32'h0200_0000,32'h0200_FFFF) - Defines the Address range (200_000-200_FFFF) for Slave 1, defined as Range 0 aligning to Slave_addr_ranges[0] <b>
    * set_addr_range(1,32'h0300_0000,32'h0300_FFFF) - Defines the Address range (300_000-300_FFFF) for Slave 1, defined as Range 1 aligning to Slave_addr_ranges[1] <b>
    * set_addr_range(2,32'h0a00_0000,32'h0a00_FFFF) - Defines the Address range (a00_000-a00_FFFF) for Slave 2, defined as Range 2 aligning to Slave_addr_ranges[2] <b>
    * set_addr_range(2,32'h0b00_0000,32'h0b00_FFFF) - Defines the Address range (b00_000-b00_FFFF) for Slave 2, defined as Range 3 aligning to Slave_addr_ranges[3] <b>
    *
    */
  extern function void set_addr_range(int slv_idx, bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] start_addr, bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] end_addr);

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Gets the local slave address from a provided global address
   * 
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to translate a global address into a slave
   * address.
   * 
   * If complex memory maps are not enabled, then this method utlizes the
   * get_slave_route_port() method to obtain the slave port ids associated with
   * address the supplied global address, and the supplied global address is returned
   * as the slave address.
   * 
   * @param global_addr The value of the global address
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *     mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *       indicates a non-secure access
   *     mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates
   *       a write access.
   * @param requester_name If called to determine the destination of a transaction from
   *   a master, this field indicates the name of the master component issuing the
   *   transaction. This can potentially be used if the routing has a dependency on the
   *   master that initiates a transaction.
   * @param ignore_unmapped_addr An input indicating that unmapped addresses should not
   *   be flagged as an error
   * @param is_register_addr_space If this address targets the register address space of
   *   a component, this field must be set
   * @param slave_port_ids The slave port to which the given global address is destined
   *   to. In some cases, there can be multiple such slaves. If so, all such slaves must
   *   be present in the queue.
   * @param slave_addr Output address at the slave
   * @output Returns 1 if there is a slave to which the given global address could be
   *   mapped to, else returns 0.
   */
  extern virtual function bit get_dest_slave_addr_from_global_addr(
    input  svt_mem_addr_t global_addr, 
    input  bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input  string requester_name = "", 
    input  bit ignore_unmapped_addr = 0,
    output bit is_register_addr_space,
    output int slave_port_ids[$],
    output svt_mem_addr_t slave_addr);

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Gets the global address associated with the supplied master address
   *
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to translate a master address into a global
   * address.
   * 
   * This method is not utilized if complex memory maps are not enabled.
   *
   * @param master_idx The index of the master that is requesting this function.
   * @param master_addr The value of the local address at a master whose global address
   *   needs to be retrieved.
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *   mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *     indicates a non-secure access
   *   mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates a
   *     write access.
   * @param requester_name If called to determine the destination of a transaction from a
   *   master, this field indicates the name of the master component issuing the
   *   transaction.
   * @param ignore_unmapped_addr An input indicating that unmapped addresses should not
   *   be flagged as an error
   * @param is_register_addr_space If this address targets the register address space of
   *   a component, this field must be set
   * @param global_addr The global address corresponding to the local address at the
   *   given master
   * @output Returns 1 if there is a global address mapping for the given master's local
   *   address, else returns 0
   */
  extern virtual function bit get_dest_global_addr_from_master_addr(
    input  int master_idx,
    input  svt_mem_addr_t master_addr,
    input  bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input  string requester_name = "", 
    input  bit ignore_unmapped_addr = 0,
    output bit is_register_addr_space,
    output svt_mem_addr_t global_addr);

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Returns whether the supplied slave address is legal for the slave component
   * 
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to indicate whether the address received by
   * the slave is legal.
   * 
   * The default behavior of this method is to return 1.
   * 
   * @param slave_idx The index of the slave that is requesting this function
   * @param slave_addr The value of the local address at the slave
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *   mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *     indicates a non-secure access
   *   mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates a
   *     write access.
   * @param target_name Name of the slave component that received this address
   * @output Returns 1 if the address is legal for the indicated slave, else returns 0
   */
  extern virtual function bit is_valid_addr_at_slave(
    input int slave_idx,
    input svt_mem_addr_t slave_addr,
    input bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input string target_name = "");

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Returns a valid address range for the given slave index.
   * 
   * If complex memory maps have been enabled through the use of the
   * #enable_complex_memory_map property, then this method must be overridden
   * by an extended class.
   * 
   * If complex memory maps have not been enabled, then this method randomly selects
   * an index from the #slave_addr_ranges array that is associated with the supplied
   * slave index and returns the address range associated with that element.
   * 
   * @param master_port_id The index of the master for which an address range is required
   * @param slave_port_id The index of the slave for which an address range is required
   * @param lo_addr The lower boundary of the returned address range
   * @param hi_addr The higher boundary of the returned address range
   * @output Returns 1, if a valid range could be found for the given slave index,
   *   else returns 0
   */
  extern virtual function bit get_slave_addr_range(
    input  int master_port_id,
    input  int slave_port_id,
    output bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] lo_addr,
    output bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] hi_addr);

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Method to determine if a supplied address is served by the default slave, or
   * if a valid slave is mapped to the address.
   * 
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to return 1 if the global address supplied
   * is handled by the default slave.
   * 
   * This method is not utilized if complex memory maps are not enabled.
   * 
   * @param global_addr The value of the global address
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave addres.
   *     mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *       indicates a non-secure access
   *     mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates
   *       a write access.
   * @param requester_name If called to determine the destination of a transaction from
   *   a master, this field indicates the name of the master component issuing the
   *   transaction. This can potentially be used if the routing has a dependency on the
   *   master that initiates a transaction.
   * @output Returns 1 if the address is served by the default slave, else returns 0
   */
  extern virtual function int is_default_slave(
    input svt_mem_addr_t global_addr, 
    input bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input string requester_name = "");

  /** 
    * @groupname ahb_addr_map
    * Set the region range for a specified slave within the specified address range. 
    * @param slv_idx             slave Index supporting multiple HSEL signal
    * @param hsel_idx            HSEL index for the specified address range.
    * @param start_addr_hsel     Start address for the specified HSEL index
    * @param end_addr_hsel       End address for the specified HSEL index
    */
  extern function void set_hsel_addr_range(int slv_idx, bit[`SVT_AHB_MAX_HSEL_WIDTH -1:0] hsel_idx, bit [`SVT_AHB_MAX_ADDR_WIDTH -1:0] start_addr_hsel, bit [`SVT_AHB_MAX_ADDR_WIDTH -1:0] end_addr_hsel);
 
`ifdef SVT_AMBA_INTERFACE_METHOD_DISABLE
  /**
    * Function set_master_common_clock_mode allows user to specify whether a master port
    * interface should use a common clock, or a port specific clock.
    *
    * @param mode If set to 1, common clock mode is selected. In this case, the
    * common clock signal passed as argument to the interface, is used as clock.
    * This mode is useful when all AHB VIP components need to work on a single
    * clock. This is the default mode of operation. If set to 0, signal hclk is
    * used as clock. This mode is useful when individual AHB VIP components work
    * on a different clock.
    *
    * @param idx This argument specifies the master & slave port index to which
    * this mode needs to be applied. The master & slave port index starts from
    * 0.
    */
  extern function void set_master_common_clock_mode(bit mode,int idx);
  
  /**
   * Function set_master_common_reset_mode allows user to specify whether a master port
   * interface should use a common reset, or a port specific reset.
   *
   * @param mode If set to 1, common reset mode is selected. In this case, the
   * common reset signal passed as argument to the interface, is used as reset.
   * This mode is useful when all AHB VIP components need to use a single
   * reset. This is the default mode of operation. If set to 0, signal hresetn is
   * used as reset. This mode is useful when individual AHB VIP components use
   * a different reset.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_master_common_reset_mode(bit mode,int idx);
  
  /**
   * Function set_slave_common_clock_mode allows user to specify whether a slave port
   * interface should use a common clock, or a port specific clock.
   *
   * @param mode If set to 1, common clock mode is selected. In this case, the
   * common clock signal passed as argument to the interface, is used as clock.
   * This mode is useful when all AHB VIP components need to work on a single
   * clock. This is the default mode of operation. If set to 0, signal hclk is
   * used as clock. This mode is useful when individual AHB VIP components work
   * on a different clock.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_slave_common_clock_mode(bit mode,int idx);
  
  /**
   * Function set_slave_common_reset_mode allows user to specify whether a slave port
   * interface should use a common reset, or a port specific reset.
   *
   * @param mode If set to 1, common reset mode is selected. In this case, the
   * common reset signal passed as argument to the interface, is used as reset.
   * This mode is useful when all AHB VIP components use a single
   * reset. This is the default mode of operation. If set to 0, signal hresetn is
   * used as reset. This mode is useful when individual AHB VIP components use
   * a different reset.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_slave_common_reset_mode(bit mode,int idx);
`endif

  // ========================================================================================
  // The following method must not be called by users even if they are public
  // ========================================================================================
  extern virtual function void set_num_masters (int num_masters, int kind = -1);

  extern virtual function void set_num_slaves (int nNumSlaves, int kind = -1);


  /** @cond PRIVATE */
  /**
   * Returns the configured error response policy type for the provided master index.
   * If the index is not programmed, svt_ahb_system_configuration::error_response_policy
   * will be returned.
   * 
   * @param master_idx Home Master index to be used in the lookup
   */
  extern function error_response_policy_enum get_master_error_response_policy(int master_idx);  

`ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the APB SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the APB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif

  /**
   * This method is used to calculate addr_sel_bits and to convert max_addr_boundary_limit enum value 
   * to interger value which will be used to check whether transfer has crossed boundary limit or not.
   */
  extern function void is_addr_1k_boundary_cross (max_addr_boundary_limit_enum max_addr_boundary_limit = ONE_KB);
  /** @endcond */

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_ahb_system_configuration)
  `vmm_class_factory(svt_ahb_system_configuration)
`endif  

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
DxOcJkwrNekTWdxGdyB9UJGt+T5hdYDFVeOdAOwoaDgKeRZ3yUftNE6JBIPfoDGS
wG4omWtGqDR3AawPPbAM0XEK5SE/wv7O6Yy6skeP/wSHu6yKdwDm7gwwDFtTVRB2
iD5bo7W/X4vVSvfOGB1nUfXXF5PYW8x1hhGX4xGgIyw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 10390     )
/D0CJKLe/XNL78nx+cgtjtFmXC6hSQtAvyg7fvrg/AKI36JX+WNplOEUIY93fSmK
L7/Mhu2bh4xfAgqbhH4EWhwYVsF/3Dayoe5s/btoVoZeK+LjiMaCovzpGrQnqxW9
OzITEUr2F8EZ47ZLVMv/uT6JvVlFzAghGd7iEUjiAJmqjEbrqbt2Uz4M/ULb3c6+
07jJ8iiPsp+mpnNuv+/v8CykFDLUce8HppYpwQPNERLncPG79Dpfhtg9ibuG6Nzx
HW8Dk473rd0OJrOj/+nbsRfmHvbPqFmf58JbYIjErcwu417w0ppC0i/gjMhDCTIe
zSaWTmcoh1bAvR6mhupKaoBjt1bINmaznNaunrcKtJFUnXW40IbkQeidkrn9rWY/
AXvgKzZOm1TAdh9fh5H+OpVCvHpWBqdLhlkTGd8jjbqYGc/AU3RD3l3+AEZ9wgDh
O3m9ylEImxSRAkb4OtpR46RgFeQE8ikXfx07SREH2Z8=
`pragma protect end_protected

endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
cHSmVgSQsGOnHA5zEq9u8xHGR+Az+O1tpRlI+77tBWp+iInt+Px68eF3IIA/Jx/B
s0foCsgVyUGNKiM1Bt+jp28mxvy9pT3WwoqNfXIBZsjyeHgDRgRsNEV8Ex+1b6yG
D27l6GdHPK9KocXa/vvFUkyjMHJSqFNLGthSFaRDqPk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 11170     )
FhowGPwGLlhtVzJb2SFfyBXT1FUOu5O9vC9hNrHes1biTABX6NRjMg7p4wpVwGYe
uF2gFwy9n6Vha6ckw8lBlVoArbMlW7d3dyNJSYLnuJlAsjezQVYP3ftpHNBIxLfj
0wELVq/CrcZdBgayqvMqHdaX8eGQ2+vHjpv+XBq+Dc2swJh9811NfvZE7j9kap8d
N0uCyB4XjOwa715LQYt9bHxZAfCeWSnau4MvSFPwEZfzkDNp7/8RbjCnuT013UKn
N3AXyocuO82m32GfkLXIl7PxACb0Rhg+OT01kg4RGENLwPOoUGjOCnsfHyzCJK3c
NeYdBlKM3zleYhS8xyxTy2xu2qslt0LHo8NQBO31tC0KHPgXmXX4mmu+qlMbiv1h
WhrtWe00JFMdkkwpsgkPr8/IOFoeOtiEWiWDNAavRY2oCpWpE+Pba6+xS55jZUjh
Rxc6xH2jo/C/K78EPO+0Oe6Viz+ikztH0HR9ENx7WX4iCxYBOfIs5FMzSCVft9+G
jJobbX1YX4ICEJpSN9mdEu5+EI8ta7wilg58nTevpmQngGjaNiDyKO01j5+7uhOY
Wi46rBm8c9VOjbTIucQqPwX0p5KXFd4rw1Ro8M2/A08GWBXNMrR8fJdVWpvPIm0C
m7gdMRWeetP0yWUGTKd++adnVDVkVkUC0ynw1iRpaJwGHe24ZTam3dYKh0yqBedS
up97+O7jIkMLf77D0cvbuTxUYLfjIcHR9rGjl0oKUvDioF3Xx0sq9/QM1Oz9bGzk
ZGL6tKNiHnMfCRbUJVW8mU+FooKlRI/F3/tNALg9lgqwPi4ZGUW3iQvhH2TI8t2O
SGw6roE03Kq6ZtA7wu4iJLIAfHVAg45rmgUEJ/W5KzOQZt6GZ+h1oISl60sLDb40
l/QCvZ1OnZBBgIQr587cz4K+osLydF0uIViYnQCRHvCFX8MZW/9wOiXjzJCz3CYw
sWPf8CNKMzOR9ahfkBtIiGnAp+0ZBiKlfbk6/yfCfRKW52GfFpSvHtnHskFkwgqN
xu98BixGlODUOGI+wg1knw==
`pragma protect end_protected

//------------------------------------------------------------------------------------------------
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
iQqEk3Wb31V+7gtFlMc0xFoYT6yQVWdxtrPri+Sm54BF6NOHWNkLIEeJD8dkujyM
kaJ93KhjKqPlb6clgf2s4xXQitKtfNEtV7fgdHoOfQI5KYrFgMGnoxRsN+/pLZSz
oPWwlM6H4k+KyvCjsU4KvdxgFj0KkbQG4caadu14DEc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 11672     )
y361A1JP0sLfRpscwQlLuWz4YD8fNhuf/3pJ6AS1VvnToDeQcx+I9Nw3Vu8fMbue
JWj3Mv/UmZMvzJ+Bl1Qro5ABRUgAeTjVLQBwHJK23SfI83AgmQ5hrVQrYgbeMyjJ
dhS774CpgAT0xkGNxTAGazXVXz48um1CX3+CkKlHm2Ca+T0mcWzRfW4eaOsLbqOv
6KpOO5FgecqTZ0iKzlU6/QgSbtDarhTMA4C7LaMO1JFAmJE142jK5ZWLut+ZhXLA
AD14XaKW9MtPdk0qPWXXmxk9FXqAueQQ7JHf8HxcQ4b6k6qnaLCmtNoDdQmpt/HV
VlpvAzNOp1TObiFWBxj6/Gp0/IcLj7fdXECHr/qI8gCdSRXq8ahQ8Yf9/02lh3vO
8k2H35S6oYsvblEuyAVrVqYcJf/Or0c8sm2GIZ07QLZt2YJwkzCmGKgZA8qBVYYp
uId9fOxmsIIrI8MxCIzTzc4vjnNaxUkS8vSSBag+1+eqInoaH8to+s3ZaAAYb6oL
rEf4EX0ozNVjn3Ej7EMM3FjBmC1pVlQg5J7WSqIge/ndef/N8hJuzIvMcV5Tmwiu
aFWBiX0Qaz2qPS29uRRWr+hMEitGbRo+FQC1pIxdBYiT2JHu8yzG1o++WpzXMZY3
JiYd2ltWMisX7Ic7q1+QV7A9BzWcdctdiNRVd4MJsOo=
`pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
eHqQdmg4TEg7RLVafpnHN3WghekOKjmAbYrQZ/eoy1jVmyJYFlFJ3UzAPMxFbxEV
KRqkf5Ch/yRVULdMyibDjzIOcig3HFG4QCFH4JstAkl2+yi34mmXY6JMQBXzEiUs
EaFsg1dw8sEsbE+NUHRrPOD30nFVqZIvGYaRWwSbMMc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 130791    )
vunna6mm70Db7GBVma9vOfOlibrCO5OapDECltpeq7nRlbSco1Tn8ElayO6jobXr
IUxixGLK1L5qzYVXBWFElnh0M8vL5nUOaEv1oH6Okrdx3yh8nD/ZSETXrymy8XYd
9uFduQ89cieN38y7pYWNevduCYTyPQrwdTp6zjf+6D1/bsPlPbhzbmbYlO11bV6u
kQqcFkv7BQv1WnFNLrgp9J4msebsC2VF65h2tR5kiRqY0kovG5wReqOph0kgQzNs
aevRDyl26yHepQ4R2rkOu0KdtfZQyoCfr6MWRwpQ3Xt0cWpafkQlOmUVBlim13mH
aktNMbhC+B/oWnQJkw5F+UOGquN+9yCyn10LzJ5RwSn19CUPVN5GSOtNZ0f89hAc
vbi+sQG22nEGFy6aNQOTNIU2AJopBnL0GTjEUjJEn11L4/EQPo1qGk3nnwxZX8I8
e2kD2Jwj4UJq9CoMfvYwg7Z2/kv82MG2iG++AF+orqR/q9Pjiq3BU73oI04YJ2Qu
b6g5u7yJ0jpA+SCwZn4td3G3uB6AbRYrhNWqXGijpcjrFgkr7fmMPJWiqIvCfNMM
qOQ7xX0MuyO0PXfD7S9q6p6AIOvInOr1d+25YgvGa93Vl+x9N21HvXJAlw3N2sU/
Q5vdnmreWICpciMdNvKhDE9Tc0n1G0YwDKciG7QzFD+Gt6KXED3yZbHl1tp8fHHK
D4h+j2gjsDTzq8aZdpKi0dzL1Zs9DSs6l4MQtEBqA+quHxLSc08L8UYkMzBVtmgy
O8hIySLbpbFeyHtwz2K4IPqAsACRUYpTqZVHI8LmuY/1pB0Uf84690ogyeT38I2+
rZBhCou+nU8DhjNWjNWWnyNMHWwn/O2cr8oykWFys+xHPwX37cMEQcCKn7r+3Zn0
e4SrsUJV1wInqNlktBW/lYkR2NYDIXSobJCrEV/oR0RPJ2C5ZzfhEG9mwGcZvhPK
BefQBhYD71An+QYAPgWIhjrBQscBPhx1ApjBa69S074LcqwzbTElI3FZG9nZcCbL
fckaYPd2TRZG1C9kxESyKFXua2VIzSbSkDfHBMMUDjYti6pKTDnXbpT3kDBlcDXP
vgStyDV+7Pw55sTObtNpgzOM5K5jebSqV6lTptyFfuAVnl2tJe9E05L68+C4A2cS
5+s6loTQejViPsJ6Oxlk5iARbRhzqHlfFRxXfApWNGKJWE0NXxU16vnQPBLkZDII
90s2aQS03UHsbkKxcRDZtZAcccXPTylEg8stcjaqWa2ir+ruYfRwH2A7LwSQnTbV
AW9LE7oZeEJMgU02WUvfCCPJ6QNhMMApGhRlP0o/7j60v/O+ywYkZ8MXDJVoYK7p
VJG9Uevejl5FN2KiqTmhZf1op5SXFg3t76VAeDOvdk6KodBg11RBzMx+WQJ0IPk0
c8z4QCv1Q861Nxqi3yrlzK/jdfYhr4phKG/hx8d3xF8d2z6Y7sYw64Tc52YEJp9L
JyYtf5P73DdtDqj3YpTMvehloH/KY9XP20Ar68fR9vlwwP0VcwxIZBwE2KrfHEK1
8POnRTasxaoCzJhklY1u4PRfI+JJv8roMn+dJQqQxDwvwt0M3sPyHqBTIdr2JKyF
fPKGhFCL3s57pPTACbuU3K1tbqbH1OXQaS6EwGsWqMQjXysWEs2GivDoC5i7nPA1
IMEt31gRBQSKMQhgeVfFNMWmRVlgXTDKdL7vNnJrkg8JesNGi4P5Kl4GhsLGYP5x
XI64K7Ft4j64yd9YeTotzqdAG+bLXmL7RDqKEPt3tzE1hKJusVPmKJ9HQ7IJvzvO
7M74HuNbVrbHxauEc2p/Rbbmm82w/KVsARlfiTVDwx0YI+wWFyijBw0hK+UHJurc
0WUo4fotwtVKEzoajcg0sRbrmra1PXj+k6Slnw5uxNasEW/k6RTf15yWFbl5T6zj
ixpCtlJdBq7dhsWcU0u/91/ZYcfqn0wfVQyYXksA2tYuw/9eKgUNLYBxGPHc+meE
RJTkzHh37CWs5oHqXGM90abhWQ+XdTB4Oxw4uXMtmNTWzxUN54kWtdDtjx/0wbZZ
L1TCHKVjiihOHQLwgGDVwo5r7Onztd7kn5t2is8DaCtO07ZME6AbGIyluM1wuNr1
v598fNEm6KkA/KL+cx4CdIJP5Xjz5pimVJDTvyFypoFiaYa4mL6E8Drpl75j3bBx
wT55hrHOHp3tz3dAICLYTaf5MNkV8pxfzY4xLN4Fwxfoxwcin2fq9EyMGYDoBlZX
FJ29LuKxG9KuEfhoTiKtC70TT7oI2iRB3AUhjIhojqE3DPoSQ2ydVeAMtSH68RtN
TgdR40fmih/TdN20q6ROxJ9PNk/xdT7eGgZZ6UiJ+olVEKSYVpxHZ7m1oV9lDLem
q2zcCXBkU5faC1ucxG7G/u6l00Sb1pokj9gaZaNrVgMiE+dEXjjjRlsa9L/Al9fX
rexHWYRVO0YYaoDGHUm63jVcqMyr8Os8dJokHbK58J9RUE7EKDVeRZU/o68GFl3R
5XOela9NpW4biL9OcjATRQmN2CoRsFPFOHke/M8zwRZ8rk00W56jaILgdn9yj/k2
Ya8HWQqBX6cN+a2f/rX6Gb832KxWgxVIek8VX1bwcawWwZaIrBuHk9uI5EDP3g+j
SsRCWXzfGF8E5A2Yl9P6An5w0NBvn6eoV+7+Vfb8B+9mCxkjbYSTRpMTpdf9ETLb
zpW4PXx31cjoHyeFHn8MGlCqO/Tl1+j5iLWeaXWnykLlVcTwFP/vxgcS72Z2c2m4
zaTxsdlICAFlUBgGAErJo74mPPyVy365k3uwsnjRnD1EZFeCUoPbZ3H3ea7Ejc7W
+YDwQASz8laJ7VqbSZP+NJa0rgvyjtFensXTanK5a+T51PHw2vei4zkEeU0TiYPa
whNfolTSYfmUOfTJxMggdZKJvKynWS6FlT9N1+cjaEtrQhNFOpEArMNxmhJZx+ca
1D0QWkgMALuGYVw6EiwE1uo3JTFUxuoYw49qe1O3C28cveQQp3EyySV7zjbViRfo
BB1Sb1CxO33iFtybiMOmVVDvTo7+Y077ypLRneGVNJCPNsZ8JGHnWrdsm5O1XO8R
OT7pTuoklOQCTzUGcHrQNultMJEi53am8YPzks3J2bx98QfamEFUumlE7m3xcAWt
ucTVS7+aNVEVnwZBGbzBBRDqpsooRfo3ZruavPqwni5V+gIylUJB52lG5g0PVBgV
9qIqIQfPvqjzcVANNiHfu8nuezHQk0wQ20f5FAvIDQSWuL0xkGQZc2aTt6hQSTYQ
dV8rjdG+lqarV3djC9GYNwGPZHdfNLHvoiseyYf6HOL1+iQoH6mdPzPWx4/WM2FI
H0oKUnLf71XHPiNn966tFmce9PC3MxLwwW0KR7sMATzvb6Ax7dZPU8oA49T+osWP
0UBmXngTexcunkHKsJNijs9HNk8qfrtRDfvbdMIdDFVgyXhBEusgRlNzzMRifRr9
/DGquBURb6OuafOZYKCzRSMXVP7xpgRtpxiPHjmCJB5hfZBEBZIvazIuVTCEhnyJ
fvFAaPXqcvJPmS0cEhuM1CHqfKhRc238kf6Vx80IW3oirEa4nuUUTxmEXMKJgLca
jj1zLPaV/xDPwm43wx24rswcusoYGOU7JdUiVe4n7XiZGd1Vs5Ev/jfxdT4EmV59
wuyL+D7iiJY5jbM2DnebEjBfab+/5lsx4uwoKAKxE57+SFKaSBL3MQJNmxhpjQz5
9pXQTETpPFe2tGENw9jwcY3KNui6G1/f1jEtoRcA3PC9J94bG/ao8e2N33kehOzN
cDSmyMb7gpwzqYVt051L9n15fqpXnB7GV0YLQLsOs3WvVnmW4Urvr0r63suwQ8UI
T86HCD0Ol9YJNAguJ1NwpRcLpBSN/jriGVMa5CRr2b5VLr9kg3oDbQe7nCyJ8QTF
5WS9l/Hmlj2E9oc5WKinlyEnLKO7Gv9peYyAamXOFRqmhh8SePp3QC8ZPdpYLKjH
3X2p1jL5cUDtjc1KSpb7ntu1Z7eLB8/yNvW2ZKzOtnwwpS6kZe3FkUA4fakz4R9k
xnAwNuPY1nToz+WsPVKRGNUJOb3dtWddMb3FiXk0v91wSJVPwQf5x9fEXu1kKzml
X1ZNDcmWBhfC6E9VaLsCNXjX0oE2Wai17YNFkCWDdoUIv++zqdPf7D1lUP4tfiiL
1bJW709lu+9li7SUtUo2QlW3WQDPrI69p5+zRnd7pXwrshBUwDJNfUrtyIx1R48I
NfxjA5wcUxkoDjuawf7GleN8nuCmF7QGawM1xWC988cvp8hC4Z0HNIjNhcA1DF2v
SGjtxhIM2/9X+OSzAYQhHg+2VBwv2I8YWkhUXUh9lQheGWZVmpSDWyaUKeOog1sN
ycT2pgp0x1YVuWqthpbS3xhNvr2xYP/s6hWDKOAVSl46tr1QoIsdqNcKVSOZcZke
8v/QBfqIzLdLFwXERBf2/0hNNVZS8cYRAokoT5ZUIo4fzLwfOUDqZ6tqFaQ1kd3Q
tGLvCJNfYHQzwjhdZxzKPaB/UYziMKRl8ZQptSAU+nGraXF5KX4WEMt/y+cz/UtR
MZ6G/JznrJXJdNXRW84t3t6PIW7KQX7kLY8Ma8xcgesa0BNUCqimTnEoqbwwouWm
hTjEVkhKZyhyMbEJSyi7jLZi3/idCO/B5TyCEl7xJyyLJLV1OhlrCcpDxanUO2vZ
zxnOjf+T2fYFwjR6Vfy/HrHyA38C13wW/vYpxnifLXix35YH+x1n960B2hGq2gPI
sPBIYvSZsEewjyhdWhFjuGxZHoNhwlpJA7ely2xngvuw4ClRhmenQqJV9TKgUM+D
Ce0ABMWnEfw61wT52T9V98FJLhfLHSD8f1F0cZbkx/10c3ZrctsPp1aZMYbvJfsM
9mWp3noTZclr/YeBaJ2JYNf8L6hSOgqqMIzXNAwVoRHaEo1J0wkQOZeSSqbKmu+v
nLl6ug+ektuScLrtgRx39ugX4fWpsYDqMAX5UWJkVVESLy1Uq/fYTf+2kq6FPzl/
4WbYa5RRI5kWHUU8w4BImJCPIfKC93zmRSGxvrnAnqbuhG4GjEjcpdhKW98KcTUX
CGfOankyArQuFeXDh5zhVGsMoQ1qHKTBDoggyPUcDuWF7oAgqYqAsvUfjp6ap9Iq
Alg5Rcu3C6DKqo36NyBsdwfIfG7g5Sz2phXmxx+CM4MXIL5aeMIzR+aLiGh0fM3J
4zeNH1J7eJWZGYA/ygKrXekpzzBpkMyq6qTnobJrKNh9Jpr1pKMXQUO08fGz3j3I
pKCqzWyrWOG83ci+/Z5fhEL98g8cIz2Uvh6iEncvewI5UyYkkwicpAmrm4Y2N9f7
uoMSpgr1wwPOCAltz28NgeERfEmrd1d+oJnbbX9syNMIoF5ZLdXu+YB6ITYeXFyh
HNxywnv39Lp/IPCP/l9N98sRf6IcXXa4xOs3eoblAA0ofBP7GGipS7yfFPvRcmUm
zuZyibJmtAYbYGYrJS+N5j2W0/8xbBGhOypdkOLNVFhFKtOlZna9J7E1xyVFPBr7
P8e0/7rf/1bNsFEvoA3axL6TSl8SSOlIEVxWusmfUV+rDOo5jZHGs2S+C7Vvws7A
qkISv0Xtu8sj8MkL4czfxYdz/rc3WoATjRUnWXrWpO+olBzKCXcGcaUiXxghqOo3
6xHYglcW+tPm3qJCpHiT7pgBwQMt74JLn5rVBw/uianiZNqdwanCbE5/s4t00VnE
6m15M91A1XsKmh/jZwhFCIn6BUeis/QXHeiP7Q/l42Gxyp+n+Mo9WA1xXw2m31kM
tKDrT4IxNi3v3lNHR8+dyrkO4VpRmo9Mz+xqiTR0KMBTjc2KwubyOkfw2pIx4dMs
keEkJplGMtjrm8wA/SAb+n/rbHbl9RT5R+6/vZ+VWvw8pwNke+dRItYzMaEYp5N3
r9nokN3rRfmI2FX7QFPvV56s6TG23CaCHK3WkFMu92ez6nE9+3iOhwfe5iaWVsg4
08dd3dHnBGG5T2ECc6M0yP/1CgnT23ene3malsjriJGFPD/DLlfNo9xgHqjYImrW
GdGz7dBjaHvCKmgquq2SjpwLSQvnKBHiMQvQK79AVuIu+Vp1SEnT19NdJJoXfG7C
nn6SJazBtuI0agqhTaLfmtfcVOgBZEXl9/uKMWAh1yoraqojVtSR13c4NAF1aSHZ
+YcgV3vlMP0wYeGTTCBchnseOPsz5JtZ3d/AH/5jp3Pe9GtZnJa7+qCf9mfU0vDr
s2jYxU5NI2unbf9DdA5CcIO83/sX8lN95dErB8fnnG99IMm0dFo4xzWdXi9iC2k5
/Rrt3nG4jGw049yfZgUw9JpwrUCoCBriv42prf5nWSexEo/iyjSYTBOr4YIIpK3K
5PKv7wRgMtaUskxg8QRGZAkBvqhJq19fvHU85Vu9hRJOGL/COYhQdtZ0V6/F7bqw
eYCRUdMMnng2XxD2A76AM0Y8goFIMOZ1AwiYWFK0FHr4jIk/DmGHQ3mNzyb1Asv2
iIBj/fE3buP96FrZiyaq6ARd/FcUbDOKvRJSW4eKBDzAva8UztKfrK5qFiexco4a
MO2k/n957mGogXeuTYZ+2jyV8yez4ciZh9CJYzcqeYmLogA+ZKoCtvpqcReXGlHZ
B6hI1vx9tJSyIDB6TljqYNUgI545PXCEVQ75HTrBwHKwXwSL7vGrTSXPaNiJmdHo
KCACvtGnBkX1csqlvssS8wYA/4dzf5AdoTIOgKqJHJm6yVMBT2aWjZVduk6/+65h
YaF9FcPInp61goPNp282YSU+SpLESyX4ztIzdeY70b8qHpB7Ji+LUPyt3XTJZ/m5
CfzHGx2kvPhcxxLP05NDNcJFVFnDvGxFP2onKmJM6PXtExzHraWMmilc3d0dF8yc
Vw1e/gkhL33YGUpzSp1/iblqzyy3bES8NsEYlhiL9YkY0eIWGF12XfBeek+YA/Wm
C2cFBgxc0duDwNuel54JxI03FqdJuSlIkMvWVOJpFyA/Hb3SbS/0O1oxJUrfpu07
kumeRkGGx7usen08z/IsD6R/UAnU+OUoeus3L6kmhA+Wxl1r6dt+hMhMt134RLIT
vZA/C3BtIFeLcYhXPOrfHVwfI+wyA9byBZNMZSfhlKUSd4O5xHSw89HPHqJiSG3v
Ef0aC5NJykJMiUALol5SQ0+Loggqyx6kkDIpagTMRBXBYMyi8uuJEJyVcsTj4YKN
LWBqkMvTMV3w7SQ04FR+8Dg2aIU8/czDImsmPAwSC+KzmkO+drKRkc1PvwUvDoTC
yoUapQR/fU0jLBIO7y/krEOvbHq9o5OSewKidg/IvcZwzMN5IOMxb1bCuPuqSmlR
Ftx9J5QdEmviPKicdo797jrBwDwa+/RZBu1N/KuYFFbee1JsKefJQaa7eLfECpzx
cB4RSPLZ2X3I4INEWpdCRVtUmnmCXZ7GYeDPQY9BkMZ+2slUkOI/625amm7oanpU
dnckbq6g/tmrV/iHmMiwkiefTvQRII8kLKqpH0ZRmQhZ3KCLeJILyYXwBgoZOsZ1
WcyxrQgXigr/6xetNe/Id/1+V4gTHIusfoo/9AWF1hgfCnWP0VskWz/rshqrZY+o
VlA6kD1gTvV8kM0p9igbwMmCgdkqq/Z4jG5+VTbLfl6ZG1VN2nLXMZacC9Rh1NxD
jBy9jvpHfX+1D9VzUcow8LPWiFM55AgyODonVZ3Py7OGhQRrq2pyEdfgHUe3bqeY
G6eVIFVrVZ7vqRz54r8bksHVG8Tjmj1h7F0xlIH9gQi0xoBFe7GGqxXGp8tUfkp2
QuGLgFUcuMcuLjXEIPBoLW1Mk4I5MvtITy1TvXWtXx9MVuWCTYVihOOm0o3jzbzx
ICKsjn+c/XXrWEirvC10NX1hBlabDlsm/m7sx2cL9g68S/JQQ2KC6dfD+RqWfiO9
NuorVbWX4I+3b+64RCZ4U0Xf/9/EL2kfWa+b3Y5tslHJyNuhQ0za2UwR5RBWtLtA
a6txa6Tew2+hXQxsyCg82HNeJND9THKZSK1ogu4Spz9Mo8S+LJYqt7QiXj3gJkIm
IGW7QDNjDfJfuOVEPKJXXXLNS3MtPQjwMg2rg3cIjR9yd4aCS+dlQgXZctgVIFTu
BtwiSHEqmJAS01p+tduGF6xLwLZpifPBxpmHqr0i+qLxjvKVnSUplT7pYZxTT2UR
MALwCQ1yJ7MEjTWDU0/z9KifbIjxTQMDNmj1fLd1AAenTzwTHg4HCP5gxkieJcqi
n413hy9s+XyLL+NQBNNGMbNSgd0Rf4or0ccBQCfNFQn51JbIf9HwCbqhHE6zG+wy
DUIKNRxyko+sxPdU2IVgBzCKqPOLcWuqGR984OMEzXPnrnzpPZLPkJnGyVilesAU
hlZkrJf4vVGjzd7YzWe9/6YiiN2B3YBwJRTTsIvs7YVA1oBFQqziYM9cMR7Pwwgb
09JarstFlgLmUrDWaFwMTS2TrSM2F7mqRWHP1DQS7MYOqXxBFX+u1RVQEMgloo+b
kh7TrEuResJOlLNx7J8IbDRkSy7hfMaCxllsy0Kcydj9L3wKiWTcZkwqQxNIGMU2
FF5egmz6KabR/HpflsQJFzm0BrfhGxSkUP8e4rNOSgGzOSO/znuOYYtZIwbJN3Cb
Sutk8G5/FjcBY27vrZ4bXNoUtNbscvMD8oBiiCNRTeu11ky0nfptPBn0BcDx0LF2
ggfYXyFM1PL54qeaX1zjSmIp5n7Nw7mVgX3hkD2+ws+O++i1CWmGCIxW9cwYRH8f
+R1m4QT61Snss8CGyquvjlDHYGfL/xVTx8n5Lr7Wv7fqCBM+3QBSAxp3XB45wyVI
E5vmE9SnCuq6mI2Kbq6tQU4rsm3vw5hFsZ/hy7mDRUXTwAKkI57ptVLH6m+iR3Bd
9Hv+px+yIcV+vu2oMSsjaHI4yyXW7y3nmXInW0LEpiJcUfugAxiUysJkZ4QwIEO0
SR3fvRNmve58P77xKnDH3bdnNfXmcE3Lh2byvoeY3uWIxmL95RTc4DMTOaGsFdUm
0Nl9jEt6/xRyUDyghNAW/XjPnVN87qGd43xkTag5bi13eb75XT8W6UbnPlP3VTnt
DRDbzGMfvOaIFLxCdYHOHFiQjDZEdnzLOn3yI6dBGDTtRxo45hmmhJP6ity/Q0Rj
KNYUoD1p9tUBvPBMdi94fXtJOeoSb/ffkA9CZBvkJsrAwvXBfSqtXLWQQcV5n/qD
8JAsBMEd+/AE1BlwrRKuxQSIjc5d4nOhWo2UjTEKXVjfR++7p5MiMGVOfccBr1dx
rZC40ZYc1n9Tyv0bf9sLnz2edPaDU/eCrQIsJJ7r2YqaJcKm6la4gVAXC1zBC6pH
//8xPz4eK5ASgj6ERZnG/I5jZy3xZShbOpzNpKTkHmJZRiP4JwxOCxt4HGnTBJzz
U/5D5NRXo5Pf5H5Pl/ZnpPIjsT6hV/byJCFWwy92tjxZr6+IhjUGt9Rbnuhi/Pcc
duTUouBKvVkG8DlsvGxKtmGq54LLtHyVq3uFqiER2YNsWsY0gt6IipfK3ep6rHCU
E4tWNzi4M+7FX9Sd/nzGzNLOeE7JW8lbhPtl6YgvwxablxvCKLjYlmpMokkEfFqt
SE4m66VbB1bkybpR5h7LrN74PQ784BxdbdxyB3t75XYAyMdC5YBHlxcijO6nWO7Y
9Wdt8PQhFRGwUNJ19bHb2vgKFEu6GfoYRa8vquhf58fa/ItxA9FEsVAxNp46ztHD
5sJe1lhJj0O57zdvky09fXfdQR08U6twC/l2+dZRCr22WEfct7I8RYAiBRhH9C7x
0nB5zBmSJBPWCHwSMcpdJ95WkD7rFaJJ0+8Qb6D6rf9fPj+MWkYGExX3xNXBy/bW
CCnXsJ0OVheUtfD81wo6/X7sIOAjy22ieiGr7v5CfgYYqqKoKZgPWLlGr7hwqPR2
RTc0yKo9fLkLwIAV2c4GhjRIxPUGI+neELkeAVIN90HLnXUTGzXVM2pfsQH0tYMy
YWa/wR41DtxajihQYBZ9zzaXoBN3FANAcL9WoNF7ticxCl7T0xmvF9oA8S+gbVBi
IN80TRZsSeZYPSoWN4Qh0MNO6qd0ezrTX2MQggln9fMdyMzQNEb2LDa3hTVkjQLi
s9obC2ezmxh9UElOrGWETA6U5y5xAXsZ/D3fP3JUY2LsYGH86oO7Md9oiU15EUEc
uRxyqqxfhDWxm+6XsvaqBuQ279id8iMxp98ehnFBtzI8ptPu18xgbTBo87DMbkgu
mnUUZuPR/Z7B8BFZNuVGN6N8z26FrjNUd028c6Sixf/Pkh7irHtD8HzdFLQGcO+v
gApb3UMIrrK4HHnz7/qlSfku0h6zZQ/sOquqQ6FV15tKSltYVn7UiTy9nYW5hz/n
wP96WyBTZ8pOlWGmOcn/Q39ofLY1TimYMgyjrxyvS6zlccmeEvUoJsWjnfEWDnCI
erRA2X6zuTK75Z3C+KFotEK9zHhuKJBLPUz+45hO4sJCsisP1q3ug1l0PYtqKHhD
RHyDOIdOHgsSyyFJk1tz2CVnS5OfrXZlD6ro9mZVl61byIXYbZVEOtuR06LYXl4R
yMklAq93vzFUCi4ixqgugnkvN2+VaI57eRlfg03oefO3RevlFpCT7D99yXdI61u6
IsOcjNeEcpZsEuFpnWzNGoSZcQ/K7fX7TZJ+QzMk7o5S1OunRDkJvD5Kc9+CkrJV
lF9csKM+AfiGwdjpbFwIii4Xop1tE1RfjSMGQHOlT01aqJd04i+0SQDy7Izq4c5z
mrd58BykA0UFVagSmqfyKtGSspFZLlv7dDVIzDSEVLnaw7fPZDT8tjxO7LfnR8SM
CqPVxb9AYcKzGhR5phTHBynx19Ues2oZqzPLTKjxmwhGtUIRfdrzthXuoB9EMEKM
i7Pt4BoH9FQxqVo5ZZd3bzQGUc0ekcdryVrPuYFzOMGYKhhtfzlN3jmYi7gYBrnd
Y0axIEtjbXhXvOE8TN3QO323+U/KpLNdIFTiOQRSvO0n5Iv8zrqP+g+otME5NL8q
iNWAkEqjbC5OXabr+5CeHKmqRe1RDW68csNjQzp/cZez6w99qP2VuskGKXCr4xTL
I1LgKJIYZiCvgWqEFgGNDslE/bggHFL0ELo18y037o88jC7knCi0Qvp3bm6rGS4P
cwY0buzJ1z3KqvaAmCZwDTTmAl4lA+BBNLqL5Et8l0mZ+Lite9TtR2YJ6e3aC46l
sLoQZf719re/hKCI7z5enwah56ONAYcUeknoNcRQZpJRQ06E5gNAv5sC3iCEL12w
Ffugn7C28ttabcXYYRpeex61PGMYFpFBvVv5LtH8Q6oSICaU5Qj4jQuoJx9Dt/Uq
VqRptHhCdvqfdCflPE7I3fYt0KP4S9AmU/1y2qfbssqAbZPekkR4rJz+cQfwzsFc
EyW0sCZwQQshdDas8xD21UsCSIdl0tEQGzo8NE/jClh9mcZiQbBcTjSOq8XRuJSy
uI5KS3/CTF8wimWd6iS6SbrAgKK96XMhlZyogRCEBmZWHzYkcFLa5WUnodczvZkr
OefJSLHfjNMVAh574zmgEGCqXt1zvC+l8u4aw//hwnkZuGAbavDdCA4t6mt9xgAX
pHIx2LtSpvkpvI8DF+mG+A0dtoReZONO+F2wUD6nANlZJRiPM84lMWmL34JW/Emf
0KNjAufSgYU8oOpIc/JBMlkhUCW20J9Ov2AXoGt+iGtfFYkD3/cgkQaApV2nV4yp
R6wAGM6Ik2khztim02vKH/VLLcnZ/3SiVGjAmiKMvvJ6AuPydm9lyWY4EvawRa3P
jXqzIGYfyoeSJsSSW8NSuTaPLBOQpY/T6O1sQ8wUUQ+giuThLvaNewPfe32/Npfn
bitviyFeYcE8+uUl1xMEHifvcEpVkOOQdYgszcG+ZAXY8tWi6sUwIdwSqWQ1aR1m
rXUyQzEyjTIH0yn+9DNO5gfr5M0rBqVm9vHusc/3u2shP4Qmgw8bq1IswcG0yVTA
2ny8oA7/UxRiGAELBHwNb8vaLVwqE1mFiIdxmguUxnc45pRBjHKs07FD0N3eiq9h
G9sOK41FhYKbWryto4wT4KfW+vGTDnJnPFflM+V9WCD24ePJDqnTMHT+PUDzndNr
f3aiQDlLryMylDyieJzqFpdJZNoJauphneAhH9Rrt380I31ujx10QkhIpHO3XPcO
FduGWZkAKoogAMe2vcOx4jan5Oqolx3IDMYQYhbGpnUvHknk7uEU4guRsQgKbXiD
x8wZOzifjUHPw/iNKPoWAOrCbLswha4WIJea8iHBo1F1z9evB0DV7beeqIy4UMXv
KKvtC9EpUD4lOAxQuLHRtzgm32tdcY7Ms6tuH7iGxlxTY16i8TfBcXOFED9FLZ9A
+Rc2Kic/+jgK3kSkTNeqzCqsZydI2WwxPjoJooeWbo1p0SsGMbrlGZKe+wYgET2e
13+3QC1IqdEkQigrgXertU4kEyvMdEirnqqxZpO9s1HyCUFU+1nGf6wWURrkFsRC
tT1/2i1P5Hu/qzFhOfcE2Gt5BOWRzQWve7nDlOpn57623doMYFFjptOdl1Zo1kxG
Pc0VeewSi4xScUtR+M3s+/2nl/YS00xdvbmmsZTKDJ8IPPXcreEh+c4kzfUPe4TK
6/GIWtpvY8qX04QVwX1KPFW7UKK6qnvX8AJV10dbzPHAFEiu2/LB/vF7NC/V6ud0
//o9sjrZ8+mQ1mQz8akGefZ3OwVPVNtqdji0QQXv/Xo2gBtxjclHMNn2H3h0avkG
aogodMPJTRTmE9ka+EBuIUnz3Oeq/JolEJ8qkEBK9faPJlrli1PU7rWeo6FrDOU2
xfPjlRyYMJhszMXazE6/nRvQOW3/xLakc7xlmEhIFNRP8kTV4YgIVzK8DMc9jLSC
vnlByEmvEpA/ywwzMfkv2IcFCdTZe0PxC3C9laB5x6o6DA4O81hHPm5UFpf1D5Gk
FC4gPAIhXEgZz+j0l5P354hMP+fWudT6+LHQFb34bznqXqA22v5qaAdyQDs/V4Ge
w+ynYujSfxlPnCcjOlRAQUH2ajQX/5iBWm/Ht8/xBpnV7KUwnmfWetk6UeJ6lrgY
TIVZNqKu6MVLxzEksX8gTidF8rjMkYzwLU7/chqPJYu4TULE7Duc/YQgn1bgCZIe
2HB3dWoP31PZJZvlK40vdou2z+tPNnLiHpsAo7uXpF8ZRJMP3MqIdyWYi6W0VRMr
amVS0VniJgv6rX/H9gpgxMG7vllx7QzYSBLJSBjDVg5BNIKZ5ldOuBIpiNBQulAR
nLDvmIlxmDQymTfQCWmQdXQ4sEvqmpx6Kz8QK6Ibh5o0tZ2vtAyOK6kcojYHeRKx
lAqgw4KnydBVkw7tHqpf5fZnVK4b1EmAA2V67lN8yW1gdYGIlG/RNRHv/mMym1KH
ZcbzYUOddkmfLksLnqkWlES1YGHGFpuaiEqJ9q21lrDJN9Ptr0LyehKHJPA1VlAY
jCXpZg1hFl+QpThsRn814NJUllqFKFsPXUi+o4YHnz7unuQ/+D5zv55oi812mOMk
+jk+CNIKlVJP/I7szC5aR3KuPqtsAZLFONPUyE6JRWlzE8ZFVD7rynnGdcejvIBb
U+J8XZoxFsl4A2ZAINthTNAZabD6SvX0KYYOgKxiOqYDXA0nj9AHZOlIHIu+vbW2
RIinSq5lpiH4gxoeuWxEohO6k3oRbSou57mOwUGgtSJwKidsa6DvOZQzrjNAQjl9
Ak1tN+Df/Bsz+Vq1lSJIDiFhDyk4hoUuJpsZuz8prr+PquQSrHv5E1g2+Xm8DupB
X6QpxFgy7eNOefsKTkgKaTIzI3H3LR5Ml7pp/y0J6QQkXQwXMOfu+DOxTuCAa1cC
i9bjPfV51v4gSIk+u0jvESAZ7u+vjyZHvMzzHzdG9pgUKBu8OqTjaYSwAU6Qufsk
FNcD47fI2JpXvntILBBIY8ufindf/dAwndFDUiX2b8cSgVbclqx492NI0d6IA47v
hG0qMoCFTidESyUlzM84n3KWM6mzqjmEutbgM46U468c8Zag+skOBkmaCLPJphwu
xkiGYgrEjyAsxLuJhJudwzfTN42dAUvQuyXffWxAX8g2QQ8gj5WlwDgcnqmDVIsC
9DV9Fw69LOb6g1n8kezAjd2hWKTCNA6mJWH2LhHPxTdZ2sMAyUf4NjTYQtvV7IX1
hf9F+/7lP+uEJNWKC5xsI1J1CHSExQ+f9vcAMWOXsXfRuQRhInWGo405qqcGd+vP
78UQUeJru39YwpVMH4ZU96XSZhAI9pOheie1o1LIPSLlo/+BOkMf/JL8jY++xjWI
4I7wM0MYOFJWyKLhgI+SecW94uZKg2l57nd6qIobFwErpR9zcMmfbOXazdH6vHV7
/jt2QAQaNAUJNXFcwtkSoAksPJZR6ZFVyZh5fMLjmxT9+cPNhRDrlD9WLr7A3huA
K8u64Q4SGPdHX7FgiY6MkrpXTHGiLVNe8xZWeJvYsxffKEqCfC4psCo2aPRiVqmg
4hSa07p1sQAiraZVAR4dwHtJV2akW7asud1jGv0jUzR4DX0+//G523CnVo1tmR9O
KCgpqdpgqsc5F6XIZCGvCzBRqOLq48dleHvUXYE3AQVUDi9VzsExEuCHSXzyq02V
DCzDt/O3FjE16qkV3rDf1huLTO9bjaHfBfVubGomqaf9yxy36Dzg168PGj3Pvxe4
ZUJqkUQC8tf5YVUKfaNgnCk2KQIpf+ZSy4mzu/+bhKIH8uJHFfzBDaq2Wz2Xts2Z
dCsTTiIi4O/R9cj9VQnus5KST58kYhyVRosJ/VzgWt6G0pRw5O3GpkRYMVzJMJH7
Hm0Mp2E8ae01HCbWMq74d3ma8nP38L6h9U/uQHylUlQIP8PkV54CBFcAHiNZlzk6
j9eC2VOruzM6cCKtD64KoaMNfDzlNevjoRzVKnGiVOCrJWVPfVyP0OM4fLV2SHmc
zgQ80aqulNnKLokRc+lV7fDQ0b2kw5I+6r44cmEED2qTI0KDMh+oUtK8RE512KTI
1LplVZ923cpxMOyonZH/kPSKKkNPX/7jekEc/1XAZm1JfevZ3KzERFeKA7cfo5tm
yQ+jNBPAC2fC5EGFW95yhsoJ9riPBYFPPKQi6nViLOVR+4FIc1dgt5AsHvNSXunO
FmcJGhntJOJ0OgysqNdmOw9tBAeNZ5OIrrG0g3UfB15RvmkhT0sRfqFes2a4oF2n
aTFQASRwlHz16c0+xbXALCbk4jU1Ds1Ux7voQcsVilpw0DTeaGexPaOKTgD6nxt0
XsZ2W5BlTSDpj06VCnaTSYk7lioQrfctEa3cwrwuIYawj/a8EBJcNqVh7hav/XWN
+yaF5hFidv4zI5l5Mi/ixDNQXlIuQGoDAnafLjJBy9q9cBBstW09Y5ird65f+4YO
i7ou/fvYMOLq7g293M7r313F1UgpR5aCZDdVZPzrvtLEKvjrL6PzjfuVpKd5x6xW
o7G5c61Eoh4/sgM61PHv+8vULTByq03RzAQGpTyzSUnvJKr+vGYCkRk99mcxLhlI
4AFO9Bg79kWPUX28OsGUyvEmJatfE5Pjh/VrmBw0aNWuq/ZmZDTJu6dvsIi6kPQ6
wS19u5QZPXDNjS30bNxrux6FQ2qlqi+ejeGPTVnGtv1w/XNsVyWZZwEtyLjZ+NBI
KnPqWIThmN+RunFIClPwon9NHo0I3yI4RLZActuSQgQC+pAo/8vtncUp6esQbkX6
OIsx7AegiaIzMf2VR+g2NomVNB/2c45ijtjPd8WE9hD154vsWrQzH0BM6qJ+1KB8
J1nNntnQfmB6if61DA8N54jgUUbIbaHEgTcEbBhSivJ2Tx9IbN4ckJnI+Re+AWYu
pVwFodtwXuEcUDiHxx7quPq3G7cL/S0OE2BfACK2ar5d7GSOWPBrd0u8yqtellVA
84IUAApY4eTEALB8JWbpja/BfcDzT1ePt4mMl2/ZFyl40FtQbNWZh8JAuCelcCfP
ysq15dTckNo8/+rtZP4fBZOWTqR8Ks+kyIw9BZw4cEJLmkZM/qrn4++OWIbuQJRi
zd9KBoabSbvxgD8bB0FBPPGNRroKCPwESFEkQ6LDCNzMY8nqkMOqchtUpkv+av6C
tA4zHC0kjPorJ4qnGWO/aCMaUaBVZS3hRL2cAGarzRk/TqwMAsxh/L3sPMe7D0y8
UzgyeKitSjWt95y91Hk2rQsfz++Wr5hOuLdjb8SO20dEkXW8dty/4kjMKKE/uoUD
gclqad3gYNtsb95EhAgIJkckV2pKkIIi1wnr5FYaQS/3FszYotaVgaPaeA+m3yFQ
X1mDX+pm+WZctMO05GTwJFVk4qsqvJVL9Pyky83y/BMOLOwCCAQRRNaLIbXUjjrY
P+IrgBvEOFvSuwNBrGU9mQRJTllHDZzmmZ9m9kD+/TRxASS+YHWDiP+T0FWBQ4OC
9NjA8vi8KCNTBkYoezojv/yLNFnAmOiWPLEX5TahwC17w05BM21vCU8yYh8uyxBN
VWAjopT3bDK3gnpfKkcXHgwu8NrRTMbPJSzZFSX4O7WWKCPGyQeJlMo2LCSvBq84
QzQ1lkDwdY/CSXUywXUpnkajib3z5j3YO/yU37NRBZysoqibpBOiLcqFIA3hyFXM
meIMb4JJpzTneUfjRKmtKd++dAucHV8LWG1yq7fxWLv6hTh7drUNXvAkbq1HUpUC
sEVEYyf3mXspHwQJlAwr06uwciETtqzTtkfCs7RJcdQlNyG/56dr+hJa1xs8SH7n
srW1XDQzX7S4HmZdOjyubxc2yLlyfuk93wl+4bOvpQx8hf0CiFyjhLmJJcFCiz/8
daUtoo7Ned0LkI1thzfVD/GZrQXAIHtI1wVghLdHndu0Ms46RqId1YNxtFwTCXy4
v4bLmVJovsgyz4+w5Odze7xH+8EK28bJv9ahb2uR6MFFYHO0dJC1GQ8HsE7zncp2
dWHlXcNFlx2XoIJQUZlRRd7QYZG2JzD10gm5vSOc8NSsJveWLiBFZm/9P41x8jwC
Xgf656N56QypKmd6KYe5Hd3Q/0+4IWm4iWx4ma8/VH6JRX+6iCx5qyhAA8Z/8qJ9
PX8ZPonxjrAKrJ8vREHj7YiX3HIBeN3wpntoyWE9n1F0QHA5clUhYPeSmRLRfXBL
V4HxrhSB8HXfL5xrpmrFwd3J9E+CKweI2ZerQNAwoxeE8VYVVcOPDQjyPi+sqnQY
GLhHWEZJdvbT6/aGKaQfLtqn5L8YVV3X2g/+jDsy2uzqAzG8w/n2YleB0mNkcJ0c
cUnPOXGUJzWiU4LfpPdh42i0nWIHQDCpMhWvxLs3EcYTqBZEeB+IMIeHHVkkKcgi
FN9uNBgn+9K0IBZIfzVZHaOZd/MCKHRJQCOyQM6mFLRPOPtnLLOGhYvH3fjS0JwK
WCJxZykOA04Ceog+1YFMeTy0G7qia40gj0op47Rcm8zHYLXXZOT4/gsTwhFSbyEv
9RW5D37YC8/W2KixSHBrfqpfdPIF/x0BYPrWFlPhkWs/BWyZQdmswT1+OSPSjxeX
Aej6ccYfqb4Qzs8YnouEN+AJZdQqlwUwjQW34TaCE3kDfSN0fZRitV8kiJ6FspCH
9FGDc1sJ+rvkA4ILtpq6THY8hz+gSSlsX/EEemPo5vJeMMnJxoBB8xdAsSqAn3bs
pocIJI3hiAcvsq2bI4eeUekSSCZLGMXR7rZ/OAsj8vQzijZjMZGnXkXMlNBOZDd8
d0SvfmIkxltAeUwn6IbXGsNpHgIwRv8BYqSK6g/OP6oXV3L9Qa/3qr1nafYI1gjI
ij6rLVKSTbICIF9i357BvHJd2ov4gtIiHCDSvlsvo1nhmTQ2f2jS//4UyHOUewY8
o1M7zLfhZlZTqu76CMTOMvrdhtyAcLsZnxjS4Rh8iFpcJEjT3o158XyIzbevVASp
kid6GVwgWwwcvCb7GvWL1CgqdfjA0ox4gUswZmUlfe6oYrpw50VgWUIV1pZSs6TC
N6WIvYA47uofIG5WYph5Ip22VEYx47NgmzKE94r83xtBXJp/ZR+3vbBeW6qKVTIh
l1MFBLaPDIRIj91fyqJ1TN9eWjRPjvoBhKzVMqy5tg/4aRjZKZYrVFez+wZ54H4Q
THru/0arO4xJaNlgP+hS+tOCHp31MohKRKI/uJZSnQIKbUegENdi5UQSwO2g92FE
UnwZ8zy1HfTl+m7DvvjZJ3agN6V+SnJNVL7QVlUeDrov9j5Rrom4f5lyKHUAXb+C
s7Z/9bOsyU8oq6CtXcDrlQNqKqX7Je79a6UhKNmFU5Q/z3x3p2QcOXl3KNRyB4Q+
0VWPyBBe6wzzH6IWz3qBjWLNcvh7ZpfLcba54jFPQDISB7w4w3Qx20YGYMdXCW61
TEnuSp+/ZCFqncAISf41Sk55ARk4j4WcnkfcsYgMqg83RnQNU7u9BjtCglBs4/ik
nBHIvu5uvnf0VCPagBqNG/pzIKdGOCsOcPe0Dt03VNzfeDvzsjM79t5GtVlJQ3xE
gyzpdYc/wcYDGK+vBETj535dKPJ68OHzDgSdepeH/Kx7xp8nyBEoLylDyTk/dWwG
mS3W5p9fK7tdn9Zc2LNSdQPavR0RSrDVCKwhUbTR0f4R8CIRLKfoauRN8C1Bidr9
TkZzNmXe7ivvVoQsY0iBvBcGfWqLzjaGVoGQMqduO+PHgj9sm8J69Qx1eN7oERM7
FMpImX3J08Z89cFxHeC7eqKbK8/9DtQqHHizFYGj/NO8FHZDjTxpPzfftsKZs0tC
crvuJvBG1YfgjtDo5UBVR8dT2w9qNLyqLnLGm4fqg6E0rUW7rOQ49qu5BqYqe5ea
7HqEg2qNIfNAVbI3yLvzhU3EwXoWRS7Sp8vs05vEthtyuGCI/ywr+GhY9JW0/D8A
m7SCIWlYmJhBH0PKKCgpenjK6zV2itLFzQOqXk7BvCot+GQlxKcYKUtl1wssZOm0
CCxD0MtzyixK1+Tt2C6Np+JPro5nzyq9evc8u0cjon9/8x9emmaPd57vd/El3GKP
ocAOQFeCNpQrSj4sFLNJyFlg4kWGCUmBGkDB1qFjaHVlLC5J9IushB5l33ZOigh2
ZPHobDzY26yB59GMA37tG37KxyD8Hf5dYwr8KnOmvkkm7Wv799ETdnmslFQlqW9l
X0O/IsUX/HtCpSU0h3DKNDZjmGt8ls1wa7lOhkaFcJnZcstgSsvfV6OORQySKuZK
UVBegoVhdlUciXcFLrCjIsPUT2ggUZb8VMudNRO66K6zcKQ4LOKNxPYEF0mmB3qZ
+g4TuDqCEl2xl/glB2HlCtmK3Lkwa2c1FbKBd6P4kEQkAUxZHkWXY9+6u3MMrTU5
FoZuWTLK20bSlBCa9GUQljOXHZgv8N2FJM2j8UpGIso46zHKxZWtoF1zOtgmobYT
TaSVjriBEzc1Ol8+oo/rN18/mWCfTw/11tCss8YsgRfj725b+dpCeh+PNANLLtoP
AfF6FXFQciCWsrVhHlkt4Ooox/HjPiXaLN9HB16xZPnYbhbeGjp65/sk1BC/hBxC
zBOBu4RPGpzW2/Hy1hFn9XH18lAcwwQwwGE8MWepWaWiOx1eEau6HXSJdAsQZAjN
B5dJ/FYbOBs24D4B9x4TaGQEvdHrg1+t/gp985466DzMhcONdoSdtY/TWrJSZ1a3
43CjXKp6mmiXOp7k17krtmrewuQOhlWTG0UlnOhldei60ihvaKT873FNXYoC1lxC
ZoxY6MZD1exSRiHhkCq9SITrQtQxJkXjZE7FrUxPiJYM9oNfnvi2M46HBJQyuPMS
vFIZ7Ylt09GJCUhB46O9KiE/cQuPLOeWlGizl1HmFQxLrQ2H4uJnLFvpzlOXeARP
emHvx5Co4AITxAoOP1ZYZ73VhUiGUUrCyA4ftQuy3g01P6q4zLllYt0swnL5wJUz
lXdgtEGvkpU7v+oYMSJD/AbAQa3SGEBGR66BpG6QYemhaAOU/xBReqG987n4vLhO
tMonm6Nq2g9PPEu7JzQ8Px3ErP5bebSkiL4diaQ7vla6Kivu0GHl7qkhpjLsLwIl
BTcQbqvXCR+96Cf7BEtuXen9S5ur2q987IAW2fORQUUYS7pB0nrzCBtumGVI++jA
dAe/OcD26/zp+kxM2z6k5tsIYnwzKSBHMxMw1MpaYOPW6UK6sg4JTxwJcnwD5Iti
opl8tCGlIHYMFsT4kaotdV9jBTuY5UXdZEOhoX4fZvQc/ZELa3QOIG8doiNTfRxk
imz5OSg7KLRUCWHXICrgS/89NOKVVA4/Zsgr+F6GkQfogIAQX2E7MPNJCdzeETcz
lsEGQQkZ378Q2iEKa3IIFgnBz8XpAIz93cabJGrZWIL7Sgk0KRdxIz2ZhWXcg4ix
gpEKa/CWT0LWTwtJ4DB4CEQzC6QZrNYoiqc8S2JQewdUJhLvM0s5O+xMyeJz4kzD
KBUOeb3Wp4hsmzZRMKy9lAgrvtMTon6DawKY6XGS41piuzdGwLgwmXYchv1QTye6
FkOKWdWZStbgb9Lm7eoNgQGH/h38ZwaJ0ktyz1Q1LNGvCzgm9GEuZkjfoocao0n2
kWmWe99gGM9pMXIw81Re9+xTrKl601x3zrffS4NAI2QEEdO6okVw87bzDTUJj5rc
cGdEPT88dn2oc3bkh/IEf/ZP9OhRkRBDZBYBMvDXLaAKiIJCl/qGFFmy3wXEyKhG
4VR83BH5QmXmtCiCHtrIoJbTv85IiBo9WRuiBUJipNmL4rtPewW4Yzw9XxyT4hlk
7hVKBCoKHbUGxUtWfr69V3FNwr5NbbJvZOCzpi+BoPFgWSsUMcSqDn8T/n5dJjn8
zC/AJ9Krl1K0Wt0y5sc9m7G0OqlDoKABfEWBIxCNAiC+Z5VTolrwQ5wYa7mJ675D
VGne6yvAjfPqY4udXvPE8i07GH5DHOTdhK1YIi7aWERYIXK8Z6vb/bYPlonNKMfL
ua69616DhGPAXl9qHtre95RfTcvOl/GmbgNTj1k9X8oz946dm8GaWHmL77knPYRa
dHRwkKW2CDuNRMg8BucHr0dvAC9unPnGgrz+6OthzOiW0EPzOfDlCGWxpR4kaKdu
M+R8e3sVWF54wmXTMuwuHxU2c1XqVUtjxa3+wVwmxmPoKUqXdUU1hkhXt5Ce8HKe
zvXY8n5fcaCSGegi8B8iRw+5brLnZ33Bs4q6vTUP61qXunUoVbFprUuUBOjjmx/J
AIL4JaxXz0RmbfRAzd6UYPJJ0e5ilbKf//I2u6jqzngFPfHYr/3ck6oF8kBFYUZ0
T9IAcrouuz9VRRhf6hRgjtGesglMiG6CDN59wYO7tPUVju/fF07piJtc+sCIpic9
E+YyqpSYMkvJiCG/HY2fRxB3y8ZjA8qbgjQtFCUOTHopcsvzxLVUnyiD7agTYNem
r13TETD07t1RisZiKzqnrTwanVJzw2RdXyQC1wNHQD0V/nUexOOA7V76i6eUlVPc
jF3aXecRiNGMjOteaY5I6otPLQoyjB28VOuKHRoZbdC8J/a1t/sA+jpvegBjRlId
bH84Oy3CYa6tk2jaTlr/fHjXIabeN0VwZp+aHKdsY+Ilc9QZuyrWPev5AGzDQ5ap
4NHvSEMaP3ZREUdriy0+bDoo/7o8cx48x35OuU5MzQgoksfPykG+7FMrhQ7Dk7UK
DHyLoY2B77IfwbesVRdlHDdkjO3e2O01M0kky5y4p5M2SRDoELP9FhEVRXVj0UK4
cM32XYQObPjFkQTxFLiWHP1WRaTVxAGNQnhAD9IFEnEq9ITQBYujTI0SqEiA3evy
B0Jx/9cragYeNF/EaPep4s/6VH1atzQkTFLtRB5YZ9F+XkUnXuwkKZAaMbA0nT/3
pa7+OOvk3bY+8zfG3cwS4tTCAd+lJXr3nbrk1/r9phU8UhIZ+x66uK46BAJn6FN/
77G8py1XrdUaqxK8+c0T3YejTExuyl2DAU2QY2FXJWf7FixatT7TZCgmT9klmvNs
LftIpZQ/mJpspQZsazlStHsUiufgY1ODiwjuc6nBQhjg8US4/TTnrsJsjTOqj9D3
YEeTn1sBEKYCKc1ykDiFVV8KuGHOaI/bsysW54UM+MDqhg2gpboDd6f0+A+8aZcT
PAg1cU1INDONuFlPwRcFAnOpcFGAWPsFYVHWjLfJ1g+aXR/YUYoAmzaIPd/SUdEf
3eZcTRr0jPycd82bgxPMJ1Km1oQrHLDjaHgj4uRZQn8WF50bRjkXNYZgcHz3uUDv
T06dznKti4o/poe2zOwaQYWyBZi4THcyV/j7EFjrMBT8n1A9dE03fM7r8PX/FW3r
eM7urqmZi9kfKotONyP4gptIKjAOp7bc+fg9doO/3zltaW+/bcD8MkBIoTVVteEd
3eCNYtBsrw6P67MON8dh4neOw9y3jGySubIuT8JWuQCKd6HdubLrKeqDp8gJZSqQ
gIC1uu59kGaSUI2vL2NAGcXKNDyayTzch42pe0ykkY76bfPSL3a9utROQzBnLp94
A/z7sXaDCgS4fGS/0aCkWqMHBOgq7tlj6coHjHOIjlOJ46eVV8TCQvxC0bWHvA2O
rVfbgprUFJSJjeNCeyJesl6Ok5ldf+qDH428ZqijvtYd3VH8g3Hf9bayz7pvp1Lb
E2BrbtI46mX1ggDiCBmswgULqv3L4O5ojVVNA6ByHfE6tBHsgZoPYE794PHJuHiE
NhfMPcJHZa13E4+10JX75ejSYDif0o6aLtqvrqL2iHfz553oe5h3a9doYDziMAXz
8tCCTAO5BfEVtZl2vRPlmyaLj8fRs0N/7TkNbXJXqIoQOYJPAFQplEePz9vy7C1o
DaSf0dGfEObC/eeASO/5XT6bx9nJn0Y0hnYLJn7lYhSLtEekwC6La4FG8tCT1iDu
/hcFtsR/EOxVMX6E7xR2XTL+ROczHzLvdnyGm9TYsvCXrHt7HfrWXNpa59lUimM2
VHPb9LGWOto5xEbO8KA/iCx15TBtm86txvNL4uunrzXN+sZidLyzpOF8Or5EScQj
myEqfkFpqIRuiUCy3X7Nj5GLiG7uXa8J30bR5JdRnLH5RLhk1MuWUY3fz+0yfOtP
ztfLYAJY6AkAK2D2M/+PsH0zzP1YGlZ1RcWlA92eTU2SgM9ctJ3Y/P2GGLYGBSDn
6TDbVej4xOTDL9kpNHtCtRRvOGzpmzoqC+wrREdd7Y4XvDAGwKgT3m5M5CAHSemd
fAznoUojkkxa983+CrtjbgJHKpXnEKOOaEMj/Z/Vn6I5L3NpaVxRCU9kQvdMHyru
mCTFHgSveYfsz3LGREDAWXzrBp7JAWTqw5n6UQCzyyABV4vb7+RmENIhg8ps8RxJ
lmiAyqkiBiRpsWBIvCOS+lxngIdS16mOfISGkbdhnRWwhBYIu7HFVWeZc1KVryBY
If0UKCDDWe/I89pMAEzfQlgjHO5TBOFPh7RUEoObUKG01YKbbkfVxiRYw9rynseR
4BADBs8cmFE855grtH54KXCkJuItTwPIF81AB3gCSyPKgxV1acl2Ys2Gn7IgeCBK
0VKAnSKDt+WuCMA+kpC37kAzeC/+Zx010+a4A+4411x/uifbflEtwoPt5lRX2qTX
OOyrGz8WCiSh4nv6Y1ad+CHIRxFxFYi1Q9JvI8snJgJD4UGoFqdFEuSouQg+2XGp
0D1Lfjhl1bOdwYun4ghcY9P+/z3uurAglBUmAP1hR9glOYXrLYcK/W5kT0gxIMmc
4zgu4liQN0VvuoZqm18+eCM2snJITEorXCppjMzO7gkTdCX9vEGe/55FQTIe6Re5
rYQDoSe5D9pRD+fddOGIzGFCENNM6Myt6tshmXE46DR8F6qEL/KM+ekpq5UNY+E/
EcfeNb9Svxnd1XB0uYoiQ6jP/CoZkUBNSe9RAsrSRVRdW94x8QGG26zsEpBw496N
WfCjFZsW3E+cELNK/k117cxnHUbZZcDpnu/gtN278ib+njddT97dC0JcP5psD+jU
xXaJ/SDLV7kPuZy6SUYdUM1EfMitUEGqCjyIS5HxtKkTTQDc7vvJDvPIg00DbTw2
dL0mbmT7whd/NmDPC+NgnlEay3vQuzSLWyn/q8LYZIlMcg4ZJb7APpGmN5iH4tfz
ry4vYSF6f5lLIusBRGjdaLITefccS6iz/+hpcfJPiozvbWllQNpXXCno92DYT4q6
Sd0mNscy0luFhF5AGF7K7UMgktljpBw3KcVWSsavWMKxq88F+jbo+pNPcfQaX7Cg
Q3jNoJObajyNAppBy4oSM9avLN1tD/eUseL4g/Ra3NEzP8IRDpTGTGVEZLeAUYHB
6ybYK7xTO+TnsvjSIwyAgi1c2U2DbjScpNk6tnjaOjCwlDh+258HzgO4/vJjWxZz
S4RwhToZtCqczfyeH0rW5crU2iq3TVpWRTa7s9xu3wfNh4JPQdoLiWNyZxeqDSbA
/Ze3tkpRqAWTSsIqxRrQ54LQtok13NrqwlMhqak6lCnL70dxQi6ZoOibEWC30h4U
ljo4z3FJcS9Ei/e4FViH1zT5bXtNicdVFUMbiapM/8YaeLzeijQGMyBDpZyWx/ZF
0m7r9WbwWTowQTFoAL4XnsWDIfjm95Gbz6lYjhZuHcaUqcb6+IxejvMgWQcqvwqb
JCcl3nDigpgnsdvjYTJEYH441v9ETjQsD8ao07H57XGtU3AtE7Z/xP59ozz281BG
daBjhTQKFQsi2CDJ1Q6nJfkLlXKzJGQx5xfFgKXTaPe9/mCsnk2HI2a+X3ZqDw1x
K4NfU7a4YSMZiG76WVOrtpZ2XGYGBnFCDi8w4eef1nB1qYHJ09/Lwdozf2BD/vgi
ZY9B92+IX+uptV5ueH9gH2xP7mVlFuy5ES+24X/RdrRvXAII58QpUuEciRjsiOVi
GOGFzKMMIgxBHzF2eIT8hGFOAwkgn9+2PkXuynYjaJhTiQ/MFnbCgUUeZeE9Qg4t
KooR5JNwgIlJuHsKWdWSnefZ5NGJIO50h0ELuVZB5ItYZOx7MUdSOtkQX+BtBxzQ
cg05u69s2aC964o7a8V3X8pTDchlDCPgWWnTHDKjIbNXWLZgLTbt3Mzk9OMiAsMs
p81sHbCiXfSdpHDZzbLhD0viBwxEKPTDcXOVlfZw8lxx/aqoIsuWNgaFefCbC6K9
KTy8tc0PHdHEXkb4tZQ25y58zkwgQwpG1VrwtO7W3C4dqB0R0TPB+S3OFFT5oCmA
XfE2hWcw37rq+a8zfyTalRI2t1cyag/y1CzfB0zTxOs7/9WrrM4lTva9v1Ao42Ln
5/0+UwUV/0Q81NZIvBNVLKt4uQH6XeNtlDlOAUQSbq/974kpWG8wHyrfAnGcxFXn
UeK+aunQHXQ5Dbco31bfKz2QmuzwB6MVXUSf+5gRh0KqtnkQdTCADFYdN597kR8v
roeodpmHZ0E260lkmZ1RBhZXmPzJgcKLirAQuxnb2z1aUhRh1ukggN3cxA7k1YDt
SM1rCSrUUwl+r3fJsTV1AK38fPyR3kzXpk2HzVddWCxH7U9JSIYMlQL9ulRtilRR
pxgVxDalDzcdocb++0lLsrV8Cxztn9zYRZXbnzHTjNU4ASeJU354PHIa/KbxNGOy
zx/E8QbM3NEglgo+6g4Oauvy9O6PQGXS9pt9jnVWIsYuIUBef7h6neB+FLmQ3fAd
ye/rbIv72gMp3rK7CqG1H7MLNW15avUAKbnAQWK2QieDgPN0ylHJvDBPNGe8Hxlf
MvLLn/CBUfAUQqg9DftqCMXGLLSOGkWlSP7ttlRsmbaFFNUsTXz+ueujPAuNOjZd
Es5v8AY0Qp+vc/i2kOtP3JhyF3nmJPemyG1oLG+wkbuiXaSR61I2JrljRZZTravZ
SBos+x0iU/6UyZfOMJZVkybyqUxTyw3pZ34wQ+eoAinzOql/02bI3V09jpxlCFIJ
YrZbQaUyDSmv8E0/mHAKsHXGCcj6sNIq2m9gg5D/GBTDyrz7xKYc17zB3VmV7MUb
IoeD5vMKXfbVusU2VKUUZsRiRJ5RGSB6JgtFsEcLCMQ/5E+AkY5C2Sc9FzyQc7RR
iY6n56NLOO69XinR2WgT9mTsqw/xlL0eIECdxN1jTX3Dkmc6oRZNRIkuztLEogiM
T7H7ajn36e8bsKMss6OzjH/lbRmGb1exuqf0xVWpmb1ScBv7mWYE3ekWnwOo7RBj
asBpI0vps32NJ43QtoHJlhsk1/Jg7TIysN58qqR9POh2ce40RExnD8jZKTOz7LnY
mynIviQt3Q8d2jZvbSyHzB+sTaDPGPU3htlOY+omKhixkTqLC51zZi1P9vjInqbV
vfSR7xdITMUUAEmpvHNgqxA538oMpTaJJXTgIf7oo7vnW6+ME7O7ISHJc8VCw5tc
9X0fHCbfefdMTtbSP5eifE60++8AkmX5UQaTQI/n/wPEox+GVfIrNPTSi4nv4sTc
voxw0zSWPdkhnSBvj3Znx+t7q8c3rmltZ7fzugvH7tJIeYDjM9cRwc3cIR+CsyOC
rwZCcNv0T0lwJ/5zNxIZweLvbBIkhHzY7z+m58wTI2PywdgnPKSNaTzx46vrUh4I
FoALMsJUxDdCHmcn6mQVF6dRDh6LwH/zr8YZ81RWFUgep0+pg8EzkU+E5327qkKp
J+sjqbpbfEfQBsz/E6qzfAMxSjNlLDFmkMZV2zsykIfUJF3TdZPn5uUdi+4Milzi
UpJSvIsEFYNhMzFqOCdetwvEGZtBW5yyhOgNhOZRmkrV0ofI+9ooJdB1q+ill/Bb
bwLNR18WRiOvJJQQJNkRNSbP8XPGGkbP/QUGhCoc81vVOaKKKYD6VROqmPC3FxUx
CoHh/uRM6NMug5iCpoJ7DfjdDJS1fFv+HnATvxuB/ZMwnencQBYId8dOrxmsid4U
UTJsyJAnXO1ewHgxUxymzawoJj1Ty+FEhHU0SwPXS2M0kv8nFJh63qQP0EhMQ3K0
Rhi1C+iHatHKoHv6nFkN/QveEtfYjF/jTUhFyJHRx7XV9pouwlACnXEHn+PvZS9Z
bXnrEAt56Wvn94+6++l15EkMVgtXFmwsNeyDCY3WWdPmwFyYsIsBcle9NIBS4Lla
g3LyADNEaeT36mIx+DDSWhXxB9NFEuMMoN6CsyjC+L+Cdwt8VFvQrnAYRAm/sLlm
bFbkn1UrokwTbumFjogCOpsFsY/48uzVvSBrhOuHzlq0i8aFOq+rpJHSt5Xi07lf
HMGzx6KG9pYRC3WXJceLxoCVNAlraaS3If5pq/8+tfBxF50Sxsw5Fcv7N8xeSTfv
uI31cXfA7duHa1PO6eJdBoVKOvJUwX3jq+8jSu7nDOqN5zSESsu2JQNqP4DxnFJy
7Pdw8arSDB1eT1R9+kIzepCASQcxnYKdAroptnBt/eQ9MnhRYeMKqlbMWRTYG2e7
U4YnDDtTYp++u9dQR6Ss1FWVtPOut2Ur2nDi15Fs2lqUqXLLRtoZCFUyPzLXhE9L
ZuEUMn1NLQCQmtqLDdlngMfvKIN2qFD7DZ17Md/pV6uOi1Iy/Mi3V/oMJ46cow3K
9MQAfD7LL5i0E8I13W6402jccYdiTx9NSb0WjxIsIO+HgID1NvAz2ByiJeAWQIVl
XJeE9tHgRn/KZ5G7xIHfTTXlylhgNVuk5jw8ppIGknJ6TT1QHSbbotbNCeXuers+
NlDwo2GH6vlpfi3c06G8HT/0WYmjc9Khhajw8VsuA1a01X4iXKsrr3gO6BYf3VFL
mlVaPTs01+yvc29czlxAP86CDqjZ3HVKUnbgpgiTEi0BYDih4xsNY6TFK0hjFN0A
d7sidR3O3YOIjNdlmOLhZr62F0piyBXQq/hFordmQ4ZMjMPoNsrAIMamOVSJNJK7
xr+GMQSfL/bPXL8IUiekgja69o3Wp5IhPUnfCTXjRDsoNdmNSnM0P867www3lL1Q
LkF44p3Fk56uAnHRvrBcXb9iT10LRYZuH9w58Vr0pdNWrAjAJLt0eATmnxUH7sQB
3chEfIVa12X6/rvYCe5FQ46IRWLmd5ktqrZAmfOflGIEWAwr0sQ1MkysXsESSdHT
q9JdTT8q0loil9wLdJ+tu3pV6/5rZ32HgPv7zh6WVxssrqUoVpyBoIgS2dfmfdwW
cDFFaT2t+U10oTOJ6NZb3MmpO6vdZ6o3nq8lova0yVVafyQrdrGCFa4N+tIytbxs
+4BJTZfUz7vlaODOzOG00OzqH7ogeWDCzwc/g7JlZ2kRK36fJLEPudehSzhnn33A
q0RcoSH1nCyhEqEgYDClCdYk8KTzs/Ch+IEYAbKjFWLvS86fVVjKlWFaVMvWA1sA
PyO+AsCVZrG4JtlZpvV+PJ6x7NVS8NzgjyXEm1rLm8N8Ybj/6yk/3IxgUBD3H92i
8ifRY+DZkiyD7I+9BqqQNIrL8Dwu87McSuQq0Z5CRkRXDi2pFXEiTjLhlsHgJAsH
+WH2jvu+N5l5H/t8ZCJ3HHO3HPClezft4pfah+g+TeOwZ166utrWiFREY4u3NAr0
mF7Y2BFLn6qWn7C7SGSi/ZBuiKAFwPgZs/gCeTCn+lZ8brxg3yFJWgKgk+7Erv+X
Ohyd/liQxq6rlzPlUNQFRO90Vu8VwTykRfl2lwwJlYzIrFPEdEuaSp86X6iswgKt
zYDny6kifGTzFryFqh0Frq/QzsQl3ycHRUULlwmaAZ+710Maqz2IDr9B82H5rbxL
cgSD3aTiDNAhNvJgrItT6Ogzsu/OxffTPoz4LqqSX8fXG/kYk+oAYQj/66Jk6tIZ
JoWIWIEwPI7KEqeNxBG3NpgsH4FBS/CFmP7mR9l+D0rOhRly2vZDRoDjSG48bZTz
hUQtizh9fjKrGk+iTGDdemu+Gsj/V/qtlt4jLpCo39Hyy/xtNDS7f4Wu7dQnp/hr
RrVhyYQuo0P4YhXt9qsM6PPZmWyfaXS8OBgNjXSof7BJqmHYXLG7WldKiLYt/b/+
MDg8rSQ/ZXgU68RPuysDgW+o8y3XwiFBdhSGE1yYuZjKzTyCynoGvU7+siFIl3nB
FLec6wS+YdvI2a1J30u55uJjgo4rqef1rmX04M0YztffdwYt7wPntiMIniV7OYhX
F/XQVSTvyfrqIzh0WwPvtzEy0dU4+NcM0cUtJKSojiiGb3xQ9r/prPkLswl+Sy2i
qNtgonqT2jVF1yWs7CDosQ970rkU/ynonoYK7VFQnCRMixab+IsnNDenxHeiRiHF
lyyrIW1bL2hxqI2RYoeI//ZMdJPnO8vC1j5I8ncx82XZRiUdcsMTd8q4S1QX+vae
mRctf9fhN/2Lf/6YhQOI0x6m1oEvMpxW+a1f/O0irbL+KzBhVRTiOkND6Vf6XMnm
lyHoncI50Kj/RrrHciVbRY1NmPD5iymJqTEja1L5B2cRqUVE+pUxUNNgy2quW6cS
p6gk+BMEH7xAMa1Y66JXz/f1h2CHHUo/3obuCWOtQ097feXEDtYNA19c6nfi27R2
CwtZ7V9FixixtcyrM8d7R/S3Mfvt7+bcFge3hAqDc25GkgStCkqyz2loPR0a4G5a
e6PnxTKSYmfkAgQa1+4v0m3ZJ/HIX28SbLfhNwLXtO6u+n7ICSXhkm9VOvs4lGAc
zr3y/1wtA81b8oAVJ18GzC0aLRl0QPrZv8H6NdbndMzvETLfDi/NGrkgucCsnl8g
nJkrLSWioK8gRWAEDLfNc9fQmtkr1k0LlU1L/QXnI1ckn8PpINebz2uC88QOwZtL
/GGDyUJ0y8IyJj1FVZ4k38zq3t4HlBgfAbdk1RZFtAqmnwRZ3rwnP6Eu1XZej4Uu
pNg9Ft8K4JfQ5J9FQSWpY08JIz+HlOn0OtymIwA/51Y8ZAmvt8+1LcyEvDbV/BYi
2u0UCbekvYG3TgDke2NUimkBQrqypZPqjK5KJvIZnOP5gJE2YwsyIhewcwzvMVZz
APP3KWXp75+0d3ICxzk45nRMqxId5AWn+QoO6ToNh+luCqiN/AElYf2sEu6tTg9E
9+8FPof1dR93rFG+IlCuhW5sH0hla2TWhsDhF8+ZGQavq3VFLuCpYIJyLElbgwHI
yNCGoZMae7c8Cc5ILptu8Dv80yaOWfVDyl+7hQCoAZRypNd12vTynuJn0xzLy1zr
7mfmxdNIPhnUI1SZhHPFr5hYFsuCEaj8L1y7Fv76cBSa1FbqGHDv5MOGa91UoiEb
5LlfioNJIHRE8o1U1s0EVe0+mQY1dkVl2Ui0NmZXEjviEszjZSyqwzgjk2wfIo0Y
OPA+Me2VttDMHDcZ/lT6MRBdxMV5BpFJIBAoDQuCIZcumpH8Vv+WV8XuJ1SMKcL/
CvtzmWfj04QQCPEhPfUVar/sDlnyoVDVY18efATk0LHBD97/SC0oFfbExgNsYzbI
SBdcnPGG/WjAZN231FGiiFMJ0AS9zZNU6O9846Tly8oAv87rKV07kxIQhRkTrupW
d+bLy6UYuXs1LspLtgIpmkfxn3hB2nzeQo61/EqGnoQDtx3I39Sc/qSZSsvJs08f
JiUC0quqLCRSWFMaEj+j29FlD+DKJz5hhx4IJjfzQwQFEzbrA4CXdVjxk2eOIQ1f
FdFff5K4396GhaEEvRBMnLe/u5iWM1QFtCl2a4/QYYn26pEBC6ijl+F4bWnAxuL2
/FCg+m1ZRv9rsGAceTjwv8in1Lb91O7g6vPswHaCKlZxV0Q4mqNnl2RkVc+izrew
DM9/0zGLDT2iBQUpI2AvWJA7ww/5+Smnb0+KIAHPMvDLKu29omTxWBKbtkhWPqJV
/NLPgY9RTjBWh6MMswzmY9SA31eCMuxkmknbPgG53C26Kbk/Jhga6B4z5tD+VX3x
Ai2mstmhiKNfAE2n7UTvkcEoH5ZWDrRIdytDzyRSe0455ob2HNZrcvVkSbsWg9me
ag48gKOagReWOy0XQY1C7ADwdvNtVOYpI1J4QcqxyIGxIe5lZJeQ9EVJ35A6TRRQ
FVh93AzOz9mNCK0iGEMG1eK6SV1BVRYxtSrC9gm+Tx5aJ9Kngocaj3NV0pyg7X+W
BzNGhhOx/8DcJOs9BlFrYIvIKMoxp+VE7tKF7HJURKWsvBTlBu0tbvTf9OaVAv1L
k2VhTNmQV0cxP9F1yshHMWxtLr2TebxWJnwydRBPP7vtCceyAJM0nuleVVbEYVLO
XMQDXFVADpiuZTWHNkTzTi2LwY/agiNk+35ukHDnfxQiozKrPHUX80MdobG7qJ2m
REGow9wxqEwhprDnfRuggqW39snDGhIYUxSmiWylIbdhJds3AGGBIeND0sa4xbJz
R1spXm+Adk7Lisk+b14yZW1ivfBgrxXZlfI8KTrfsrO9TNy/+aOttoJS9kychixU
eBw+7PotIiyeOOVZ6MGFZXHfm3hNP4sODhuhAQSZRTQjgXz6v8vi1jsRtObhskGO
9Szue+5pJsrD3wCXmjHRABITtvWgquh+HOXWgJ/kn2nD2FDO0nQErrMz45/PNUO6
KwIe+L9LiIyov76WbpHGiS0ZDJ4I/oWho5xXUfpJ6q22xR3YLrXw8PpeIDo2l+kI
1Qtrmk9RJejucQpMVTt1724YqSb/NnkG/Zzl57TgivyNNuWGWbKOwwiWYn8HAn1U
Hto3ucBeVd7Uy/oiYKkWUqo/1GfblOqQjR4rgoX2UDiZ8zaM9aFv/aOeipMrDt4W
RiWVwT9B1F+5W42YLjBCZTYtZfxogbec/LxqkaPau1q9Z7trBXMbXp+FazzLLEwq
q3xns8SZoLPezuoBlf/CqaP/oHSM/nwm88t/bOJyCUyOiAT4Wfjq+AcVx8ckEjzo
lBQxfXiWv5ptG73W5Ook0Z/T5tQHWnkf3Bh+kwZRdMRmZNcmwVlxA4f8mW4K5yTD
XXFtj92vZwVWnDDeGCgzx+pbN4Qe1R/uL/e9EBil4XBS4bkwBwEUQBDY61LQ/53T
n+LoH7IGp8+xerKdL5zfgaJ7LsvayMW3xkVV5FZQZ/BLM2Gt/9SL3VKCJguJitLh
r8nUMvAoWPW9n1uEK/obJ6LHVScV/M9r0q6G28a9gEZQ/gMRHnIflDUtI2RJitdp
T0FHMAiiz3JBvpyHPGKoJeXmLAOmvyoURcB7JSL33OZGI4otpXlBcWy2VAKHLFze
iKtZNYvlS8vGsttf054zByfmNQpPinPMsnEImmQHPDDexOiX3OFWEEUSkrY2Qy24
A5D+SF8GEplUldyxs9O9wD1LSFWFEUzlw52j1JHhLtORhojVxqPnosM+ARBabWXV
2R5muILcb0nLcD/R5/jxxBfZaHQtxjsfJsVR7vWMuPMLTHEZ69Ix3L6BlemI+bOC
tqx40LU7NnQapw4BB9PATXpy0u+hFr36FWCp+osfFb4We/p5AY5fGBddnF4K8hp6
166tegL9sZXKzBWpq1H8uYLjRQuQpcF29j9FzqIfCNArMAt8Mktn7qMoff3QbOYZ
kFSHZEBghQVmtQSL+q5Q2dcUVBYurRvscMlSGCdIMOuYaBPE9CvM0gjmce0C4rMB
Bjy6liNCoYW0cbBuBDauviUavyS/Vi+fhnAl7Rci8FMyRo4v46/XQxw2oQo4P+k0
ncU4wGvzidf2n76rvUReTdcscxwxCzpwD/ZrEkiVh91LCEuT8BFAp/II7/W/5oV4
q+Tar1NrbviH2h6x+ebIUjp5TlJbA49JGk52pQzTFh0sP5CanQFp06awyb9YvbVu
8QZhS0xb+ImB+KtAW9RHVjuaV88/8tWw/iLy8kcN66Owb8b8uKCQjq1LoUiZoVSj
fsbPH96b0bbIXUf0UFWhLGJWZk3sKqvzerkWtTrpyD07jkFvBogSVun/X1R6mxvf
uIL0s1lCe9SVqEMHx/J6BNlcG02ubRdaL6MF6ZmArb4CY42EKfx8L9saMxEJWLu9
fbIczYJApKX2rgaqHrvn4QPRCetGRqSqX9QB2eKss1ierxaORscfPk+Ua1kn2eOF
PB/Yqzao3DVXBT9mWxzwHy2yBWVPmmSB7qN2sa043UB2KBao6grtHOZgY3QGrQux
GMnRpwYLmDSW9bHY/bTnY7EpmnO/q8J9s7drC/G65xsaJh1uUVOcEZ9xzHJ+zLb7
IU8YtODaytm0jLRxU+FjvKfCbxlK1MEc/gQcrzSavR1Sf7cngWP4jqcBx7/8/GLM
Y47myuBLuleTsdrP7cbORGaorx8kAJCJ4ie6VthRnEJNsS1pSrV6Tbpg3VULX3+e
oNPP9WK2FNzvj41QdiullySb6wEt2e6dYGG9e47xNFOghQ+WZpPx5IDB0B9fJ6E1
lkeiLc44joz8KubZ2fAUspsKa17d1U87C9Vt86vJwMM04V8IXsDb+3PVtZ7SiPXv
h9ISnI1jZLnnG80SyMCC6eDxMr3Y5SHYdAb5/whdcJaMcl5zuqFz3T7xuCVETnWv
EdxnJBiOtuLdotIyU5Gnf4aQdjvaMsHDAG2baeKJlRtMDQ09PM/1QB8+ZAnp0hyF
kbf1LBtOJFoBBdX91PpPVdrdb2PH+6P3w7jmqLNYIcF7OX9IbKBD4fLniQ3GBlyN
ECnBMlXVK69kTgQvOEkptYVFDfHbrX7SFB9t/BFj6piFt5yk/gdCpDRDlWym7+ds
GRmq6SqRGNaVm8qHFPrq04G5lu5SJKzrCgFZQTXVQFzPKX0HMBJHJHeXZz//vx0W
Lo1OjBcMaJb95+fnq95A195CKFyoM4eiwJVxzrKvbfxYsGqNMdMUGM5BOw+on6CX
jsV2q+3+IFATpC8S88KmwWwqTrlocX7K1/JVXt+lOE/oCe58bYni6/ZZ17w4Y9Q4
0fm3+vB4OAfVgr04QEZd+xJ2mI/pJ4ZEI9lvQZe81QGj71XAnhNfzJOSWYiWA8uV
1yKqu9ieGqNSDL9Wq3feh1SakNeMRywbHIJyaaguPS6tTd6aPVY19K+m+AO6FYTn
BkUvxLBjW9BxM8Dn5iYAFaoM6ktIV8wubobnfdKKJjmr899v14BFIKa7BYMP2kqn
WmpI+N8WEgyfKmmfIEqNCwCvYAJQCLii3vCAI/77qVc+VDX6Dpa70c1b4FGaaOiL
ohQYXa2yM/kNGcEQMIiEWqcipx+0067ett5GoTwJFaQO878Huhm4u+tRze0bsSJg
5RLA+XsEmJFYKmQlOCMzB0/gVfSKMmdXNn0UZLP4zmprGWC9mSBguG+fRUWkSTNI
QcRFTLLnMGq5N5B3AZJitWUq/uJZXMKzcZXgU4DJ8hTZ/YX68+/Q4YRP884rMhOw
8w5uEyjSAPUDHquZrOWuisFPJGww9yqJ08soR6PGVqCANFeHmK7EINkGUObTInC6
DIZ2jCYEPA23Qg/UDSrsRpBaTs7IZrgk7c17JVVMFEjl8aQEpPVXb+VgQqJUdOft
wx/nk/sUSDoDa41C6TIa6hLqZMDRoE8v/L/zd0dovUJAWqM+RuQA9BUFc3P+t7PH
Bb9oD19HVvkKY5ivTx7DzgDoWBee+yRJd1JSx7D/BaO8/U2rTp+948R7lNqUaQPD
xQ+gzMvpqG9yN9MNyxVGWlo0sGhSA5TMosT2HNam7y7DQTxCopuScBABDJ2gX5q5
H8XmPIpWzHVrvEei/8hIdpso5XW+JVR5XGJfio9e6sZF0zUcC4CsjlsBN2lP/59W
iPx4doghkln44R8NiTgihI3euBfKQy95MI5DwrFmK83OX6bzIsf8TdGxU8s1ZFQ+
QIaursu+wwM03NOWtpKnuZCcdAhl1w8jNmj/Ro15Qqg5eoooSmk3zzHOmS2pxoUS
CcQ0x3dGq6oDCRb1zkg9liQeRM6cDB8IZyacE90/lHSUSNDKfzF7f91+jVQo94wu
QqKP5LgBNFvHfa1LQod8qmHkfyyzt9Be8zOTEpawOFpsgIiR1X7FzvpD1Qc++frK
LJqd7GSm2PJFN0zmHAOmPgJQa7ojLexDsemSeNBQdKVcbjFnXggaCWG2THgAfWt6
5DULUmsj/yJV2i3kUvujIGQMFcbe3vodbTU58qv/PPpxkNM3dAyn6tNpbp1J7hIN
owvmjD0CNkrNj3qzJykP5HTtzPry0ugAlYpKbGlDlGhKS11dTJ9fRVxqKTH5RqRL
avEA9K4TLmYrukYNb4jwpISybukoYCmWxTmcDj0rsLrDvF3YHNKxT/942Suwr+r6
hTvsp55WmR88vNeKFT86Lgt0iIYCA3ZRMF8lCDvQPeIaqV1AFfIoSvCZQZ7SvMrz
A6CIRftZajAbjCND9tfcxk1qV7Yzx2xAlda7krsmC5/zDzmMLsZaf4YhVXhMZ5pC
vko90Fa4DjkRVOPzLZHIWqlsEMzD748m8uxm6TY1IK1sZd91YlgovnMgmCUfcIyO
ZFDO36rm0PID2D8ZPWV6u1qRM0pbr48vpWxCrpIAfEcWSps2QlZEDN2NbNI9A1pd
Je0cIG1hrLMxYmwoJnN0TncOiR5ML5xK0km4Gn98s8SJoNOYRrTFlxC/uRph0SFm
gJNENLoEuXEClwx+zrQJfeHrR/LN3LOEVDOHRPN43WVojiXMq07EFAeXEmfA5RUR
0u8QYWoAdYYYwmvTOOdwfDOZer8mQO3V5jqbp1HZjB8eHuH3nq7ywzgse2HFfS1/
ng8PpJW5iktp/Hn1VmjhIKhZT/P8NDlW6DuZww0QitgzOJIDijOK+VP7T3kwLH4z
73lAL+GKbClceJdxenjfJSNXHP00HeEB/G4Cb+84m+h1Ysk+yzpkkDJFsfqGaM9h
CR6OAG+XqR+D9lJj6+w85dagJ1jpwgkNRsviy1q+dxUTd1m4HQvLbODiPZ4wXQpS
tDpyQ3UYMgUp7kAQHhbL53rt/Ky+rVetgS2eTQ8FSODO1aCnuilmc6/a9ZTpOv9J
WbceD9rRGMBhtNILnKHG2+i6rmlA6qn6RhTuRnN4pFlZsEhU9qPeSmehyVmoTVPT
dr9pGJyyHd6nk+UMnA4pRiTp3lB9bfhRlu69QhGR7DtmXKMbEp87AygVKPfx4olX
mtKdmzpiIpewsoaYqxlMQcBo2+0ps+ASEW/zyigaXZs0kHD5L/mONQdOlRDOvSyq
GVRWxrA4WYiDGyD2sp+IY1Ov+sgMrpNtAOVEMG0W+NNWjwq95ucF4fqWfXbXkLMn
Rr9C2BrDWb0Gnt4qc61AgczoDW86jLSmZfkSyjJnvfck25ze4idt00IUkCGj7pFQ
T5R63peNCeIWZ4pkKXVAKutpP7Elx7iWIvkK2jDWIuk6GrkLrmb7Lgvb4ZWBAGk1
H6czEVQxFWp13jSXORmgjBeZZTxtzQN3+hMRvaXpfVFUlrehO3J45EY5h+7RL/RK
/yB1iuCfDmxav3X0smfSzXNW4AgUl2ptEvNXM7lg28qmID0Y/ttChYbg0uPGGxW9
t6pDnZMMm709gn1NLOtoCivAVImEnPS0SnNqb0ylYK9YIb7o520HOw5lJxLNUTaa
yNRnZ+ETWjFH8BBuYV4LEE3pB6hyjsIVDsUptL1EYTRHR5fbP662i3nSy1aw/7Zx
0EE6OVr69ywsULAVDv6Qo7aMwmbcPklN2GvbgD7e5ZtD4pFrwPDIVyt1cMzhaQCR
d3wNtmvuZmtCCQSpJnZOyxWiGCVrfEMKBOg0748poiiHpekeyMiOGFnKZPQl0kuO
0IkcjJKYuak+cD/I+B9CrSWQ1U1+bDH/+GmlFIEoX9Z8o+y0cWYcjWberxXANnc0
3XZPqBfyBTOUGyV9yyV8G8rWVxMavOa4O78CfV76CuVEQ+IOmNB2t4v58IyiHS72
I66MzsAlYR9E6Lux3a5kTtHunPHjGfkR4CWLgzCt0rzs8cAzGcQS6c8z5zyNxNz/
eodE65S76Dg7Ph8HhbXmYfAsumcJD0ydCV2nAnJqEdeWkEmjCULanL+N3lB6R7/Q
1sQxEYX+E6h7KIDsxb7xhmClPjicvdNXNcUjAlAsdisFPqv8x4DUBbsYIbSUNRF0
TEOpW9U9lIT4aVvTGEVM/ePoitAr41qOB8ivYgErEtRM/p5RaqHhzaTJ/gWT++Rg
bQaJ4RQIYvbWA6N5/IYntJ76WzW9N7rVBO+DGVbsU3M8zubnxvJRXLTzeo96CTMb
X75c9l8asR8TLfmuUwqSc+gHadfOl6AftZEyakinDaZtUwSzTg7XKR/M2U+4iPKc
sJqpJoZsUGFys6f6LdaApjehTOiPsXQnHnBiT4l9+KntIKwymDMUckKG6pCdpviF
ZyQtPlM1V52aYwPF29D4K3gOf3kk3DxAMtF/LSqQp3bm585fhFgpkmzixNKYLpTO
xraAxVYc292K//L6Q4JZSpNhGVKLfC/fyuetKBf353s9Ex1maUILbx82FhjMoeP3
PqqDobUWM1/+kv0m9o1AfGB47ME9SkDDEHwntDN/bYF3dN/L3Yk1J3Sp7e95hS9c
Gwye31a1uDyAF4niU8ocpswhm1OQMGapk2iZ8aGE6eUmzv4l1RG0IjAvW6tUrN25
LXSi+9aZGYEFGLiRcQIvO8Yf3xKqBUg0imUjbJtoDvpiuH6t567N6w5fX5FBEnTD
ea2A6OqBmhcsWkU+so2Lm2d3gOfzi0LSiOSANoe9KlQKIaEdil6u8fwJOqzplKbR
iMo+Bld3lVQeN3V7AUnc/TVbdPYgEHrIbva/afm0GK9xLDSv6BbH5A52qeFmZx04
xcQPYwT7Q6/fQ5Yynm2HOFHrdO6ISOeSlAxAZf/EKALvYsY+pMpVVsVD4O6i7KU9
/mu0LUOtkTIH7PiS7ZOU+xfNJya+SopXut6vpKo25U4gl5mdeYe3gVhFKaQfUAS4
aF1sRnhwh+ezAsE5HenOOjHTaQieQP409k7cnNojYNK3DyTAYKqTfppViBU7Ya47
tfy3NzQVhQD0tjTuUC4QJw46XRfJuaSFPzsIL/hpfFqS8YQUQ75d+AZWyrxX8ci7
11uyZNcJGsn29o5Isa7NtB02qEEhSOUV7GDREZuYAYnD2n914xbbjDRrL7iDY/g3
MGIOWp/ZKE1BkTuvYUMfWHz8nXVw1XoZp9+zXqhicH5HXedRWn0+S8gLw5SGo/in
UsCIrlW7wEt54w4ANSSkJ/KDjGvw68xmpDrm4INb/CZbThAZHrZFjVMs89pdDG7j
eCTIijBH90T0fo7GCjxyk/oSoljen/AUUyUgsw/iJKOrHUDaoM5IQ82ikaw38P1j
oM60kClkIdhqOTAdnopf4d1yqD41+wj6b6k57vc0kjul5LxH+kV+TvCgFSb0g8y/
p1/ZnA1GoK196QzTIQ6Oa7Y3SMwejFbViVUCDWH/vkxPIszkhnZ1zJmbVud7bh9P
o+RozREzQM6RTrJ5h4C7GCX5w7rItS3gStXPWALWtMbBApyd+srK8rEK24U6eb0V
DV9mgIZF5klkXZaQphlfnLgnVb/1d2L7D31BYfIlImhIkhJ6Sooq4zGF4WDMmnOl
pmguwyyKPycBbtva4o+lC3an8WsAyLFdcCnd0xIGVTF6JTvDj2jELNx3FKF0GqKj
lQtJSyxoP05YnkcoXrgBwZtqbacCFt4/MKzXNn7jYKukNACjuvvb4K9Py5XuhwiC
F4aHkziKK2puGhdu5JtMlwkMPbxYIIeVBybn17VZhuWwr+foq3ZSozaMotk6cmzs
5L7a5x7jOYnsoqKW+7lAquz1hNDJOwIiAnAkwsbjH7jsrTZ7/BUgyxxv/pQD70Gp
tHmnzAMgPSBGCKus9A13GealOWhE4rDhOLiBMxJQ8wA+izK+wyI3wHkDdSE31//r
mdniTRD3eDSEsq7czwtLm/nAGOLb9mmLrcl9S1A5stgFQ4Rwk3OdaV+bvFWwvE3v
5s/Yvd8hdhVnN+fbNcETA7A3LqT/gqc/C3yJRUfAr0crHQ3MukYX8YC9QksYueKy
Vd48UfIyqjiDvvwhuQjWVDwwCuewk6J8/uOC+g7Lmcx62jOL+eqKEvMTm3g75wD+
ByQPcAEB6GbrQIWbYVcj++beWnwTr3fty+suKj4se9vTmtD1Rz8WGh+WNKbIXEVl
ud2vHOCttPK4oAOdKJWtABlC44zLKCJLWyIuieEiA80gdWHyWaemCe85NfacRKh4
voxIk4oghCBpQhAfV11VZiN3bi7sPDDEj1bbiO5woAraAvw2Zo04xjGhG9XqqCrZ
B8fwuMjw4mLF/8F2wz1NEUWun/1E3ysJ1VslohkKkukHo23h/6spO7YVv7IhD9iB
uvfYAH9hrmTTRIYJTv1gAOG0rwQV16uVkQhUgkYZTVZiHiQkkMXStpRvAC182zYM
g2WiIsQBMP+1y93OHnZ3sp8TQ8BsFYTXnjQpe4m3XeVMRQ58PJi3b3kKERYvP8FM
ejx+TiiA4axMz70CGL9+9SzXg8WgGAlzQm7g9dYNNNY6DFEwhG4Rv8+n7hnVeo6k
ZVUsLHlxXDihspD79nNsor2yp3mGY3IDUH90gjopA5jhcvZk+3fjiIe86xDyvPY1
mlMa/BcNgdVTcQeZtv7G4IKqnZ3ZlYJPhQoHsj6Cy31MkdBNEDV5XOWxNNs5bQId
UqlgEfFet4rY/gDCTFNdI1+rur32Jbs37AOUJ5E+0J+aGKIT8/ouoEjQ2Sx9iSuS
tJ2l2guTFX4Wago96cR170JAye9R5KSKuE5BiOAR3/EwC2OCYS2fVj5Atnb5kizS
YBIX2trStR3Z0WF2u040ZK9yFtcOcQvsmd0GSeMbefa1R0tvxgxU3/2SxT2mUrno
iOLUYWGEYOzFJVzQTdrI9vY/gmx7vssKjhPLNSfSUh3Fe7q5+8v/Cg78nTEuYedF
3ouqFG+5TAfsat5zhT3XXXoZ2+9hgpbjTQnrEEeGnQQDewnBJU1bbaswNpLB7bfZ
XEidjvu/BJQS+6B8wGs676hTtco2WqGdKrQQFpLP651DG/8BfI9siChO5GG5wbnK
znifotU3ry0ivfR9+BcyTXRloJVsW0cpmbAUKV0cztRwnJp1uc3a21SskS4Zga6p
rvM5n3TFlK5DE2rc+FApMybON64VWzKWBbqEunZOi2K6Cq5dCSkj7WYd46iJTKD0
x9nIQhZXntLIHJaMDu3ipPwntOVXDEbvvGRlV2j/8rBj7UIJn5/H7ufJjJpHcJW4
shAieSTkpUMZJfa0bL916fH08swjz9FFR8owKCE6hMoLkwX+EbraUFqxG3eAhcvy
C/93ZvuHkqiy0j98nNLXA+hsIHbv87cQgYYSBBRLuhr9dGdKUs8Xr+ba9cLdB7gr
ZigPJxJMRHFiA9fH4GSkeEwx3JroBNfhZAiE3aPmnl+tZNj/Uz5ag0tHSykYS8It
VycFgmeyVMCgIzmRG3HJFLo3bp+ZqWx1YvHrlGyoUo3Oxb+biuC2/cSAuCgoS9Vy
2Tmj4MOcejRoP7CpqadLCnc9jO2N9I6spnEv8zzLyu1e5DS5774ge47Br+KRl8Kz
Tjk+Y07ykAB3D0Hc8Mu9dQ3ucPsk8Kd8twuMsLSwE5kDZ5X9P7DD3Pq9rxdZntVw
7j+3AmmWNbZ1+W9iNqOzp5L9UcIeMFF+ScmFzSFqEXwTkNSPNytgQ9KRWsp3LB3o
1fec5OYeGRPnACHTzD3qvuqOdbF+EPN7zsruLr0632t7l2JCULdDi45sZkBSioQz
jLn/JL10D1NZP2GZIev6vEcNlXMjC32xbrd5cF53DqBJ9Iq8dBMTq5iORprqtJ/m
ZOJuoziqK6YFiYkGYIqVv832bN434bCmDcM9qvDRoLm9g1rixy+hXVjTTY+sm26f
JbuVIfWPdas1iLHgtHdbBOejLtlLl7MKdPoPENf11wgv1uL3QdFqC3EarcVeSUig
jyH5Ju3JqSoa1YG7zj+uczjmb/FaxxK3nRcl3ZZxlQpD7VQqJKlCr2ttz1BBYh9o
lVs3OjduQeStGBp04p4D+gjtMZHD77yv8QB6Zw1A7JTLVQitRjivglFkIaCNMCiy
rASzeWBEnvlMF40b0z6X0Lq5w8DuzTsYA/vAOb5VFWnfkYzD7BCAbZiSs+77MW+I
0KM3nKqt3od4Ux+aJrNhNUqARsQTlj75EIB5iSjz2XYa5cYxuQzbsAU1t2+8T/xq
A0c6KdFkp36+O//gEMGW7TQoMNX9mkTI3JcxIx+CBdaNQjN2nr1DIk24eyIBIXag
0bqlwugGw6Oxt15Dm9S6edUn7ZXCWRtIbEkBL1Kyj7ItbXTTgdHiyo8RYOE5/KCg
kdj7Sl4LWqgqoOX22Oeo0US2pEVEeZ+uYrEMdHfy+056suWMtN/rAWK+W4i02tzY
P+2Cgqu7NILhdA/hLtbbqcd7SMEjh2inuVpxrmE9SBblN+IXsk3SApjZOR3ESXdT
7NTElRepaem5bLiBNxAXpQAVkofLGSgf0T5GpGrLqdga+HfPBlO4rk4PH8T2rUns
Muq3Tq5FFncogtp66yB48cQKLZBScY1wSMzeHIAEdN0I3kMBhYUfsaLqNClZRUiL
iTMgtioXAE1GoaBaR3h3rzUtGDPFLPolnzWb0p6PWtLqUHOqJMFhghp31sGNyZXC
Y57j+J0+ARpAwiVdLSIbqdbADJdnf3ItGKs+f+8hqcxSaM6vHngImB3YUZHfG9NU
jHcAclE7+pgTIRI++6jNc7+fduyVjswko0c1EVmvWpx/jOFUq0xLiajJWOAd5jad
aD8E4qVSfl3wJ87G/KCmPZ1g74GKjukoswDkq6oy9CN4exrLX44SRGztXkjzc97U
1tJWrSNTb+x9s7WHW0YemGJIOsC8lO0vIs4gtmAn4PSbSVtD6Hj8evddQWDn2Jja
S+udQ7rUnPLaPjcbnXoJSjjWqKvImTso3qqOPXLSUA+1SZS5EWwyXGfd9/wTloPf
XZSjAL5lq0Up3NmnexJL2rsayeNhJU543h/LF6oka5Z8LeICktPYyPWUj0i21xUe
5aWyxgf6iUkjWkjumSYFB4CfZuMa2Va9F42pP4ri74aFVJ/E0u1fhpcKKLFyx4IT
9TRhR7BiaQEtqlOLkyHl+kL910bFeeJanAhA0uzWkE/MkqbDPtzutIvmPHfLng5/
w7Nv2EUw5gYu8wivYPup3khiutLVm0NRTryEYupng9DCQGK5dCsLFc49hPLAMoK4
DG90KXStSA3XxjkLCeiD2Voktcul8Ox4lngYXdkzwvtZbxt+qRdDOc7CVZ71rKva
U1cX5LFJ8XwuDiJzdJ6FuC4F5GouVYhlHHrVBYrSo6eLKKOh75y3GQ+hSKNhbElG
Gjvceg7ahn47w+Zd0Rr5hzO93d2A6S8glEnSPHBvVOsKKMU0tI6j7ojkkHrJyD5+
Du4zCrVXyiycgAOnT3lf4wzwRDf//HgI/1OVu1UTfz7syZ4U1wGxuQm7Cuey1250
XOcnEySSmBagtyaQkMFTPuuBDhBTMp9jejuiIrO4Jwb3EHKCIOC/egXq3GaIEHff
VkcQk5JDkp/Y4LBTMPj9zaRgRKPzaScxQXH+3uNGtaoWYZbXgTaMW3Xfz9HEtObP
5rYfmYxoXxvusbPynXJOIXTfpQpjIr49H3xV0uenlDzqlKNDB+fXt7G8WwbRpWt9
u+noNtsYUAlDzqZrR+F9zUeyIlumcKIrd+/o6H0f7DBRxDAZWrLf6MgrXPiqgmxz
Z4qCKUZYQxE4uPjR6rBbwNo1YQdphWu2OFU60lKRNKW0uBKKQjgymEaCbvEMukqQ
z2K5bEX2vyxAhDlGCp5AwSiOzTZiaIGxnyNrBxiAwZsByBQumqqV55U5GPzcA8bi
MmK9GvCdhM2rGh9VMPeciXQPU/bawMIE9GBdLq+xXpId8OJ/aR8C3wTBKEOBoaQu
MsYciHTq6Z1z6uosd6CaNzU6lgQ2cVH3DWzcxMBp6ffahpdJBG+IIhbXKaD7Q4AV
NYoKBgpN1YDnqQMyKF3VFw0j56ih2Gb/ekY6lU8mSIQqIRZV781h+gJ1giPr51pd
2aAfbAhr1oktuzIVtcPUSA8e9qNui/o2L5fefpGHK7p9+mltXh0BXa7W4cGPF/kh
mbxJsxJj1zwW2rKS7PSANgaVsoXmExnwj3pq858bop7lcVX3MAVEvsZ9ppR2Ne4W
pY4znfApZnTNAiwmRSKzi7PgDHRQmABkF751kerA1HpFfT0nbWjkanc7OBdogPeP
dtxjJpE+T978AsAZ7ixBnHtAPLeXH20gEHyBWca+m4g5v1l75W6OofiCElSAvPcv
3sSWwtawaf4uQtObDqiNVGObixoU2LkmuZaZfhkH0kSQSwSazdpKeYqFWAOQ2DKZ
N+VMQclgb5nLiaI9SYOi9JdMW9UsiWsUqS0YkDJFOfwpP+Mu8cnMXbBOL/Fg0+1W
Wp1Sb3lTlNQkSD+NADivykXb+8u/ysANKfTBjSqOHaZfADgqWNv5an4VAmW/KpYv
RVkwtEyjUcLHtO/blZfPrl69UPkGEeuXB4lSl6Dm3HMFxP79MhBK208SuLRlrc0y
aEsRRrfU8K6Vx0o38JS61AcgAp2i/pnCJww3/YGBurVtm5WSPTcMYli9DUGm7kUn
Z3gVoiBeyIj/EiIM9FmXi+m0+nDiGRJ6NdNB9jJ5UE9WKG3t9L6ESllFCQuJr3RP
9kQW066vk2bsMNtrjPxTfFwB6wyDxMUVoht5qsgVhluu0EKnrvcK2+/ekVtNnwhh
mXV8qQKI2oA0x4cdlbc6ryf2YJHdRAny6qdDgI64IYZySt37+sgibnaPVBFYcD3n
GHWdaawiAtyhENd8EUoSarotHWYFSeErCZeHIUTI5JeViao/Cmx/YriiumiDuXka
H02w1kv2Q1VF3PwPAX1JAJPFAztCrrAurnYUPHXL+3+hsz3WjxyFSUXxs2zB7bX/
u2WPa83htUTjGcMh194ADHE984pBLGGg4Jzy6vMj0+mMZops1shbxlYKMVVo1bX1
EQVSjhPATGkuF1nM17xH91dcCUoquZpJB1Cg6Lq4hCZXJH5EOqX9qaD8KXn4eRdH
RXDmK6wlXXArlEqyZ8tJ7dJ3qrwAkg3+ep6pe5yI9cUYQT973yz96LyiUMEaxvq1
WqkB1yCh8H4SFnASxO7AKLPzPYvmeVIinf2Pjdlt3HE0q7CBxiViF5m42zUXi7p7
Ie9YDdPz2EEMuv10wr9nTRdz2WftZNI9V2gTEk/QAEDDnDk6sHbaGQ4cLXk/0rw0
8HlaTL0tXnC0z0KBS1O5fHnSpyWkLOnYuBcuFAvTnEQOWJOn9jDwGln/d7VrC++M
HSDOLZm6/YyAtijbc3ej+IKdGbeY6LhCNidBIhpw97BJvh79pQZLIeWyhbG0W00T
Gc4b4NwP2xAQsCV+hOsGNZN2m7OhMCx0l2dkhDaHPusQTjZwM2WI9Z6nwtNe1ftS
HfVaejHjB+HYLeOAJ16YSaBj1er6wSk9+747sd5EOep/9/kH6UW2XMB5896o0rpI
hWHJ5PmeAs2uv7u44HTopSApNfoLISLEiKdK0TpHRGNOIBKlb3I/wnBnfBTf8kN2
K5VImno8a1ELJ7n3WrcxRFXFbrgsKL4HfPhonzirCAK1JosZLxgPZGMCe7ZmZ0Ya
0jvul9dbMEjRLKz/c5d2C8MZStqbRNmhvOP4kbpyYQVNEpSqr0vD+ewcwMAhv8S5
SqWwRLqKDUoYM7Ku+f5BqG2nio+/rNvPPwacLHrqlF6U9yi3Zjz4IuPX4iE7SRv7
jjirgxZILlI0ZO5B9MnIEN4pEXQKIzKDruF3qui0HZQsTDJ2pf+is18r74GWBPxe
XJ/Q1LYF2eGRDg/a3Fd7DGLb8jSw2pKKAUt377cNV02q7FfQMbvnWUZ86IVu2ps5
Cy4DBmXLysnFWRWSSwvY7AxUkZlERgembGfKzWWFXZcecXPCOwFPWTE7H3DfrQDb
lb0a7NOH5BIzUGSGa7SA7FwBzHdV2E4T4rd8ls4MIuHNOiplVmfc0YGiFpvdqaHm
c0PvHyaUgShTWbxvvdoll2D7T6LPIJ0NTZeXEipvdKR429TSYJorcCipbI+fb3PP
qqX2IjuqiUxKZOkRRt5qBMkHAgFmTHf4J8UFTUdyWk3gRKliSFBUeLJuVkc4KpWi
LSnrAavJZl1NKm5cZmV7hwRhzZjaxWlkVTNG2qvfrXzzxShsTLF6H6DDYmIbkzze
kclPmJXLqUSLw2ch11vHPArhPTDY114LIQwun2lR1P3bwwxgpZBWuoNs84e3u41h
E5KqAbmsdHmyUJSt/UWnmV8OkDSkf+UOuuW0YGhwVwXDK0aYoLU+46IVSK8TMim/
R/A8fO3wF7d1QYJiKXU9gLVcaP5hvNKPWKPiFOtI/12dSgIjdXlco6aDnnB9ccrb
3tvPEWJD7UnA7+h7wZu8XeP3qjHEjaDIrPGA0DkTAR2XEJrTtnAe6XU2GIqeIHWp
6ZG2FfbqrTy6V5aiyARBMcAoTRp0SdmBggLPsPxmj2EdN3mlsFNww9DRqRFn1jSr
zsw2YYPolBdp4au4XPQs7TaWW4soAlXExHAfW73BGn+kpAnYbFILpx8ycWCQIFxO
oY+WExuRgtvHJ89YwshtykOCG8Pae0qT/QGR9r+dydxjVWCuXkstiSAQK/UyD8jV
Av0hZMOYraAReLAVZRpvAjV04bAbtnkBwMCAi/APXIx5VmaAXdklV+OVZM7pQreE
UdBADT5RbgAjbs976HwNXOYgIzB3a0fZmtbx4PkvXJW/cI6FwJVSrcTL0ECEripq
5RgZIKYIWLvmv+vDi/T1mpYaPpvo/HK3vOlMH4s1S+QS5DD3tpndVWLRh0nlgd22
3r6mEUIh0xduf5mn/v7bozPxH0snsqDkXUlaY43kM9qJNdUpvhZXfByL+cPCWHdm
r/oET1Fniol27VI/rDMJEuUBTzLwehHqpDH60qQx/STETxwPjcHxhDvdL4J25Rut
U5jd4DhWep6d5hgaghT3TTlO99y8ZjqSVQ28WiV7XRvIl4y26Ac+t7P78qvNGvYU
bjvcU+gt8d99B8iShP9VJKtk4wEYs8JU/BVMm5ESDNxiZ4QYFzVhzs3tf7pnUW9g
1mCSVYOP1c/8ixRJ1NPHJVEqUP+Yn971Ftso1WgrweNHTFeghCrgydykylUy4wPO
/pfzSkNvh7pSMabDbyyOyUrvXxgr2S3IP/PW04d7IbrvLdqrNhA89F39JHd0WWM2
HzJh/IDrSjknMJ18tOJfImSmCAQMqg+024bmuKbBEW4trDVemQx98OsT5W3pLepe
/0NAFlZR+R3x2O2wwt0k30segqBLnQIpiYteryozCz2QKXNhmyjN0HV4yJYUJugd
JOsfBuZOrfsHxIlfrPjUHPS17SZwLP45EItrjh1agh6CoBCL3Ev3SYLiVnLTrCyR
9yTsklqrTR0Shnws51fxrIcNjJJRawN6eZziWdJa300lmyBTpkoYoisw8cSLHaeX
SgBwarW/QKfNhYjrNehYEMLtaCnUj2GrSG+1PxBp3KfIslgCoxY3bTqtgCIqDlxW
r2gmPDSTGnY3SHgx8J6xSsfqDYFA8lQgkEHigZsUJlPy6wnxraiLxRXQR1E2J+yH
QNvLeJOMPtGtSc/6vFZPbq+Cd/pyvFAN8j0WYmCw+Jep71CL1xQkRKIqtpuNz8kb
T6iQO+rWp5960KNzX1b3Tj0/VPtG0TGnFjQupyUApuEGLgChK/Nhr44iPuVH/ZdM
YECxt2erXNEJGk3VDmxwqbUEEa8qrCrJ3+Kwgs4ht5spvql/+pZUnuJcTaYJ6TLJ
ggpCzCZWSE8AiZR0h4SxwawURU8XG1Jna0xBex8yHucnOL56bdpUV9WDdHcuoiI2
DWxYsIH0Wzqje/XKjtskvsll6ea2e+jWpJd6+KL4a/wUYziC1Rb64nBmGjbQMCPH
2QyTQpPKLdkLwEyGozdkC9LhWSIwYuQ0dwGlDoOqroeZfca0iMwpvbwL9ZTi3rLC
PGJDFd0xDL92Yrf5tapKCJShY/CIlzBvg3flTnJbApuZr7cGWOzDuRJGKxGOhwYn
X96xHT8wDGUJK/sKunE23szvHnA4Gazez6/5fXEjmBK6iUe4mXWtq/KS3nug7aY2
6PaJQFCJMXwQ3SSrHy26iDEK6/Z/eDWvK+8g6y5ioUoXi2PqYGleoAA5MEwzHlpB
MV7qXJUe2Lb8MjonUDH46PBUisrPLzSAHLbsOGCYh2bSIBphDueXIDuTYzMxkTzj
KTTIv0wkDu9YpwLq/+KX6NrbCHInfJnxc70V1Rwcjx/9yE7HECbCCe+pqN8t/ozk
e9Nzlp42g7gFO1AgzeqkRiqRub8N/RCo33ADjzWxdM2fUdJMwV1o4M797BWEQIU7
ccly7a+u46e9g9RmfCe8wrPgovUQ6eIoXQidkDGw9+xemJDc1ctkglWCiKJrkp/l
8vAragBFJcuMzsMSLTSQz288Gs244PS4sUUV42q2Gva/uU6kmgPKoJc0zhoH6yiI
QHPXG/ZzWW8LOMK5HniG+xi+iO7GFx14wpo9fBiPI8N/CGAybC0h3tsjRj2t2kog
kxpTFWWy6yRPw9VmPKhNb0z+QCRHqSq+TsJSmQDEVJeXitb1AwizveMz2HrFk7Eh
cEcD2oQnFJkHWaEhDhV3q4TrfZRRLKdRup6ffaKvkTsm5ChX3N55E/GAEWS8MWdK
nxjG3dKBZkHdc62hD/gFD1L62/hXkcvhrUnK2qHDyty902JiwRvYYaLYmYB+l87u
epEJAedGUG+aL5buQFxr83Z6W2oMBBe8Qas0f8Fedq7Mjd5HZb4qFsxH2SK0HCWF
AK07GASrPPFVTiwf0pqALqGr2M6H2bgoxSIRHVs7RfYRSe87K1pOH1JXrbuD5X52
ONnlueSuTsyG+jKwx8OYF63gjYN4fVbY4fZ3h+kaGhgvVG4DL76oqQPOcp5SCDlL
/ojMGlNVMi/iU/AKBNQNKSfoIZskFe5qvEhS6rJ+JGHRI+9EDxJNuQWGsyYOlncK
sQFOKKdkq2W8jbvYGRh3LJWbUyvmvuo+CkmM84GBQ+zTcAPxXvdqviG8Jw18WQkc
23js7SfzoLigXFMUu96ZVy7GAKKdl8EvI9gCcuJYWvfcmOwshUXYhrNt//X0j88k
SAtmLvptB5NXRoglT8y+7cn8nqZ/PWut7+Jzb3CZQ0RGCwVMxWQvIRAZvdbYFPnJ
lDjF/du1LIH7/4cQJ0mqlK8Tt/9j4NyZmbXk1tGtwy02bPZZB9VaK6gbFM+dtp5V
c1Lv19YWaij9yvy9Quq/Z5elyh4EY2vmfmiJo9ISq3VZNbeleYHiIRx5jeVDNpR1
x608f+8khTB0mkgzr7/mFuwRbykd6PSXEiTYczusEjbBFT87Wwn7FX1+sEUypWjN
yVORmEw42BxmvJhXuNsWqc3RgwPpchZBOt/GpfWwg8Lbu6xFVgWhYgy54n/yRqnm
R1roKbrqBkGof5/Ccq/L4q6XSSyGYk0ORO3aQAhk5Z70+K5cNXhDg0gTkYmCh+oF
apy6lj2I6SE0OqHSVplpvDWZlzRRe2yvgHqNwKWiFaCXl3XLQMsb+kck5KxNZM//
I8rLSRYJSE4dr8Ld3DO/K/5e6xCKrNG3O9u+Uva/iGaXD4jZzooDWEAc4V1i4i/M
Fv6hJnuKPVNARJ2qL38Sqh9u8V6NOiPLBMdUX0qbGSfgP8q0areacG5Nqbb69Gsr
OYY1QY8OtUNP1uK+a76Ivu96v7ytQDFqpPBBvQ8wiMumW1g9ex8meP3JWPMtfNmB
WFkBkRfPPgQx3DZkLsBlYmC3dD8TwkWmObDFKvqDtNzjypqXFM+S3JM89dEJrVL9
6iLeIk+Xv/943EJXjgRhklohF3QTImeLmqrR3H1JZ/JjZcM3P7euUB8J4uNplU3h
P3yBYSsLbqBZGu41+qlD2tTTBZTAWyZJDOekCIyAedt1WasSdHcoaaPjtdTzh4cQ
wgr8bEMS3bCeDMYNy39tGAKxdJ4TL6wToE9X/6XwBA0vcToJQRghkyr30w04PMiO
b4yxDr2MiEx2A/R4WLs9LJzDXyHjoytszkwvrfBCCh0LzR9PVfQQgx5xMFcIuDz9
RHiqzoOe2PPoC1TKwJV+WxIuf/6CSc7R2GJ17GM85ZX7efz/2XUrk9QqJiBaQ2yY
0lkmWF3Zd6s/9R09v7RFj5wKjPC7uQcAjOaPxw4op1//AidLLcl3Z5+B5PyFiDyU
8ILk3tuj+N5Q33RT+ZPz3UIkrGFXHpv5/Ss3njBp/C0y5njXyieKNeJdMX6zAfQk
gEFRpmwq1lFN4vWZ8CKm2Wsdc5wqn5wpZeK5nwA0MVWM7/j91WCpHbwant0TfifU
n0zrhTSfVeWoWp+5/WRQjbDjFUf8kP8bgwY5lJ3a4TwVmjg2w4R21G7nYrHtkTG3
lzRURHZxGneS/nTkBg2esHmJ6zQ3ilnGo/MRnKt0gecYU9ATSRZ2y0IulH2gSHTr
TJ0FcEldOmsbrEVLEg76jPvW0xNbrGhpGOJbYdvJJRml2Cofr3Mw9b3BaghNvmRE
YNnzBoGCpSnZUClZYrh7YEiV7DTN2mw7fy4rRmA1TXS91+qS7fR+A2uOf0Y7pRvQ
k/Ayf1L/cRSMfe9cVnQqb2kpVsCp1hwdmBY9rrMGzk5cmtlz56IOWiUdmWPR9W4P
H/vbxURUbIhqho5Cqbu/A1izOcjcuGZ7JYDdSbO+kzvBKclt+fnw2oi1Sdmr3v4J
/LFewrUk2XXwfBtAsDXONaMO/uhiUgWQkUYaXZjWkTJumQxeO445lmmVPOV8THin
2TkK/ezzC3+VSRWL6KGZbbBW3UQNMKXa3lhcTeQEsqZGMwADKduZHrE3Jd6xMGUQ
NGANUXSAyjfVPCsnxvPp0Wg2/Y/dy/h+E0pAs+H17prURLANPaqMv5E69yM+fiaT
zdPZ3skdglQBqh3rPmVqhqX90SeGsf4KQLSd30ihtb7CcgFJlz+SbvxN+cQoQOII
U0R6r0SlxKycBYFAq3FY2Y9yZAmGFBCv/dFmLJOWjkMHKn0abWjYtQ8iXG2vUJlH
UpiwQlytoOINmIZ9iVnxuW12AZ9Ly/gMe5vYC7e23sXMQnX9WBvscoCrhCiOa/rY
0WDQL6mc1SfhE6RIwqrr1q7Z6yale9uqoWAgeBKhIDWRH2iGRsdacdIv5AW2Ng4C
0acWZuAqRFTNTX8YVsIqpBSQyXjzUWUsM/K/JAywVeKK/uhd2zsEvEBQX3h5UFAq
TggIECD4+V4aE/SN6tkr5VPomNqXb/mkbWsAWii74HaOnv694yQMmDGmNTKj0ksa
3k2pfC6WkH0FVlCDG/BIkTX9P2agBq3w9VDPTWdTFmuxF95DsIROIhAdQ+a5e8et
bj5/Pda8NzZ0mApTVvdUXJ8IjawYl4tZfw+64jkmaVsrLNV0jE7nbtHbEJELEnTl
Ktw+u9QDoRXX5ADm9zzCFyEVJFWs0u+yET8bg5GkkaJhSwLjdim+XKF1123676KO
jumiKsB4ocD0ElNW0KKRZ6lVhFBn69Oari5bk2HIn0oWzvr10EZpVzo4IbgzlyDM
NoyATeO1sVjAfODLt+IWiRkdC5LRLztkA1qDxa2TL/Sk52Pqi0YtpWmIDRH6aZZd
u1t2gjYIlTN84XW0SCdwGykuxLf4LLzaLUAQGLLucO6NZbUbwAGtg6sAV1C9SL7U
BL+5iIQ/H5+CPKt3LuP7V4iywbewEtVtdCVcYyTsmaXAU3H0vzB4F2YLpOxDgUb1
2yLzwLPxDVNr/lUnKrN1AqWPI8fhtCF2zUHyCf0DUH1VAHzB/vqmsjSIT6TW1woC
s/H7GYjG0C4cDGR+VyLfzyuXZP8jI7T8JTzl4m3EHr4oie4vBKityXT454DIwx2x
DfbvpKf8xmNLriyv9IKx1dqoJghVyGhz+xFODT7W5BkdTLkm7YyGaJNUkYrhixgz
69M5pjwGsMLMGpaalZS0Je9wIC9M2aPMy33VNlOO18K6i+c0hSlFhqUZ2ms94jWE
K2DU78FkQFsS7kZG2cNNWAGBtDuSXaiMZUkhQFw9EUIeLMZx3aYuYvqORb/jrfQd
71MXMLLL6TzkIB3thTeLhRWoHNsWsrRgUYe4WhqFO/1/ZxLBgCemh88j3FFqulsK
GjbDzAkw5EcadfBcDX5+jaOPEtzc4wEye3/6/hPWJnG/bJMaktP2CxJy3FP5vDgT
SmBb8ExdcIJXXpgf7ACtVKRqJfj4cPZcsk8c4W5y4MsYp6keKN+mhadPkUbk9a4V
rGUNaheoQkXBFkeEAgoemGrDIz+y5Hlo3b+ozEOKfQcbqDyvckBCO4zQW0DRzBhq
UfqBr32jEsyX35zXSeP39QdGP4dNBfMvHlL9BDFExyOMitGK1ACvxIh+C+eVrIvz
rGXQnJNRD2YGr4l7/ElyZriup1RDQpfjFHDQReVx7TIm4ZELjmaF1OVf0NA/r1Wf
JKXjzeGbOc7M1iV3lMdfYYvexhFP0sBT9Oju9xlbnMlOmswGzhLaI6iCg/jq9ntv
6J2kPyP9uVh3hWW/abX67syccWsWZuOBbnZZaBZwqzckVnxMh0vjoD22ncijTBAr
a3tfe1JsKob8Pe1UMSqOHK7zDw5J5uRq4AVvN5ckLTeBnFTEwpY1uiFlV0PZNhzR
o/mUUSzvTkGoyrIdyIqhLcRHRhCfN1hpxFhfN5PRQYuJ3uQeJKOwdjfx1iwV28BO
Ok0shrHWGh6q09W1dCQ2HTeZv2CrumjpEDDMK4WcPvda2jQQaBzR8q1YkWwD/mbf
MdW+KWBcloYeVpe6txR4B/mdps8ZUMHjDldz87UTzhAqvSBSeqIdxocGDewtJnLS
x7cCjXGUCaCzqba/noKCBERwubxquncfuG0e8Nf/ozAj+OuQptU32RUslXgVNci6
P5VA6TtCK9/I1R1w8Wu2ngMNm4o4Szf5EqeiLZt6ef5hlqn0I14PY7D2yPzLiS47
jxRz/ghNgY8pZiQvHsoC7txNlCbLFOqz7oUNoYpF/StsfVMcpYfh7wJyUCEkuGcx
/lJGjfjdGybAJefJokyj1Mqbhkn+0MCVWglecgf4u10rdYvbP22cvXk0oI8H8mHY
BgNNROO4fE4vNFOsmYunzsNqPM2HCQNMkL4cbCUg3QUz5Xf7wV6agNSr69EhKjPn
/Rj0hGmGYoCyTvbDuLCPLzq1k/X017Flm0MOVeGeBUuUa967+wrsoOz6sKQZPVdo
cKvi/vfpe1d0LflWUCz9kdISDHHdIJ/vIfpzI1lqUkG8efkK1VfVr3UaepWr72Ac
iDt7iH7oG40q1HQPqWm7I+xrFTdNxS29HjGJ4xm3rcvDbW9YAQtz+p9aGOTXutMo
eoZ4Wg+NSnWlCUQtvRzb4gSXDmKUISLQcQ0vfCvlRRfxJd5fE67gejuEcJTcwizy
Q/TnThlkzGPW5F240sBtysXzkJY1vmwXZ+u585uG8DVRhfZP0mEnBon0T4wMaBpS
yfCbCNmNkma8cBczHCYB8U/6LBG9M9A6AwToyvmXJ+JdLHdSKNnS3AU9DZ11qeJk
OfEZX5ntQVcHfVoGjP0AQG7bzswr2PGMh2U5wMcYAfIGm0ZmNemjg8ZjLBbK5p+O
5abTGmn5C5UgWQMk6bzOJCFX/jjwsQEdcpF/gMRDDHsWs3otuWlWGoP9q9Mef9v0
iWs0lEt9ZqM6YEfALW14+CQd4XILFi6zaJe/qswW+oDLPsOts0OrrE81/5ilLwmV
MGbfKidjxqA3I8HN8MLnH6TQRoEM3sOEyoBvnFq/dldq3OSQptknqaYCVZFq9f3n
iN4Pfn/gdbxXfXLOw3tkFT4byOaT/fWd6PTMi2f+vBqkCSN6JR1sQEb/SJpQOLjw
XkC+bZXlgSZinE58/5VKy68sOiJn6wiEUMTW77edZfGIBWvHRI8LBHIGqoOYHoB6
j8DsSXW361WunSM3fBbjcjSttK+dUSnYtg+37krjb+lka4qyIx4MKxD6ZFo7CICr
83d56B3TG0TTkG+qR5OSUl4vE+POPPv/MYFCz7S6MiH1V3eJlGNUm2oW7eprVnt2
jL9CMCwL28f6YoAq2p0BakdbW6gpuuXbV5rcdY/6MxqXaTPa1zKOTZXfriVA2io9
d8iDPCJixQEfg7FuPUV6NzGEqJR1R0PuXICXRag3ECeFWp+Ob5y8ND0VuOTfqF4V
Nzt5tprkjOUvpSuteViZ9Bo/ntCU+Qpdmf6R2NsQlkklqPkbWwVQc8/jFKl1O/S9
ozWSQiPrQ1mspYuif9qmo2yLCpKRMjaXCCU5WAMP0xC0j1FDV5s6gQ62e0hcAN5D
4PoezD8uyjCf9PXvSRhFyYjFvM/6qgYj5Uon89lrkCMkZPydYlRDjxJD1Uj15n+f
boUY9iczWTL8AJrbx4ZfgUov2eA1lFI1LdfUKLAWHHVxI6I15+sU815XCRktawn8
viyzY60My98THa6CdXGdLx35CUv1MpEfTVqtomKqfFhRwrCEndcWdaaDI+04jZBP
96K+v8KvEEiNYIP4MLZC7R9xGlQlooXsVQTc6Ii74jamTb4NCN1kVtLse7QojNiW
NZUR4XzVt9vSQiAgJJFy/M8AKacHbttAmsIpZ65IWjcuaT0O61nDQ2eU74All4j6
H3j+WQAuzrqV3cwsIA9YCRlnDWKPJflh4cQKgVUTnHNNtAKWci2vDsdhYXR3x8n+
pDUk81cZM0s+rjytSqbb0hBykgi0b+KlzNR+DhwF73CwmPmBpbxxnI/sn1VjMYPx
G3APrp0hyUF/hvVTbCIxueCEFCz0f21bytoty5CtKKq80Uz0hevtQUaY8cx/XHQE
JoWo898syzhRbznCtDuOc69voTOgXn5k6UJ6OBvg2l8/ZwNRgmiHAvGTmjFemvZy
gUeFE9HoS3fYkUuuaSPhBV67skwKUyOCgzOH8YECtNmSSw8DuxFM2ixyhoSIHSfw
ujFuV53NGtxpu+a0dfsKJ8gwybXhnv4G40pJB34WIYfyi32TOYAuONfb14tC1YL3
lJ6Fav8jWC90R1q2mq1BeQhKviBVUW6Va6FWm/XROVO3XX4AmxaEFJaSeWGe7O/l
nNt361EsZsrPthr/wO00Dtb1ThMJ5HUCasIO4s7Wbkbl+9q+LJ1NBmPjrQkprghX
OfwGvylACt975egzTLmHApR02oXaqrKZZAR6gQKdf6KTay8W6ZhUIJZehLyPhk41
9fBiYf7lXkYmakwUjpjRSxNK+pxSN+A0i3rhOo6dtXzQk4e4u4wvoAeHXBNZdN9a
AFvBd5M3T2fdU6n5xr0VhwyQrUSFgrDJDXxP7Hce5ddJFX8YAwkmvdL6PyTYepKp
xJlDPXuajz0ky0KNoB+7MzV5JZ2QEkYSmhPg1zDfC0WPDHIb/SXBtg5qx5wAnoeN
YUZRVr3qoRtn9OkW6ExAv3VxBmK4AI4ZJ+0Zb/Ve6NKffuI6ud4ld0OaX4H0Z7I9
NhUkpHM/S+5yfyy8wCw5d5TWSJfueXVzC0P4xwluHAxKACpIehFiIwVmgCwgxtuE
Qyvu+Loi6Sj2IMi2tn9YrYbKQEJmDLZ65kQojeujLJ5uAvlVBAMbfg8gXWvmwi44
1bKI6/qOU6VRpW7i+vmPHr82nQyUQHa49DIylG2WHYOldI7fw2FwU/6uXEVxZpJe
5owTOTEjOGqL6/KwThQjHUMXWJlAEhsH5dAvB8qzmCgAZorkyQcbsgJbyP3I433D
zH2PakIcLv0S4/A5a0iXu7h0nux/2OdzOb37TceGTg4c6A3hDFIU3X6J4oxgKTPP
Ai/T2V6AWF1eyP0L3ekAmrPRMIZZCHCjlxpJ65Pv1R2Tz/TeSdPaK+1Z9pIHtst9
zbe6DzuzRVxNwI0kaECamfbwOM5/+QzMg4NBryrvNaoxguvGQbpoK2zrgxAbKNqA
B0xlZhn/BjUfkTsxKi/L6cfTgbeeIv9uhumSqBaMYWrXQ6kTH27Xpf468MabU/B5
xe/ZsKu0i/I44jMzpUd10Q/z2Voj6lpwNGZIOUb/pszi3XPeemIAXM2veNjBwCi/
rE6cUC+BgEtmK+ptiGQFIzNaHPnw6HAGFzcv3cue0w/VqdD8XGoC6mpy22sXrIq2
zbi6m89NDnTOE2MYLDc1ybjajic8iy4/2mMJagBrfkTTNA7zXRFvwl90qEocRecE
wPqVCUiBN4DGJa/FaSsJ4ldIZqwR7xZAPDTh0YJ0vkC3bguv87dUBfd/DNE+br4H
JNemNDS3Y+ZJ3t7s6KVZmcZXEuMlVS6GOhbprFo/ICKaQC5fmzeJQ7mfK/60eu2g
7TgzngPL/0pL9TcTKAcuABnkvZooD214thsf4Dwygc+I3zfKwvQ/UrOS68n31ZlC
e7AUjC2FK5sGf0qCZHb1ej+hXDXzugbsL7ef13Vmf/hXj/0JDn+PJIcMAi2PdtrJ
CmZ+ofS8dSvkNvC7AadlrHjbqnZIQXg0MNpRa8ascO7Jfda7DFuOeakOApeC5VS9
e6v7+0nspqnXjzE+UcOTYDNO+ubswdNgkW2gSrQNoYjaySIc6HeXbk8fAvKWEhI/
InZVHLmBzplFvnAC8jufjTkdIu7rTZdZeNp9nDy7+mXawcmjJL9DphrC6uXvsW9t
+UwKAZareyz80SMJO7/nB/OghoUSBp1nsEbwMCTtvMjx1QkegfWbTSA+0BX4wDSU
PXDUYp1f54vqitCtm7+Vip5CR0McXuKmcDyLZMihJH6pem8BHq29cuNoJcfBhQ6m
A1kY3r/JKaiVgcm6i25wOGrMGlAwStFLiHXJAj4RSnj17gk2TeguF1pue/19bVU+
+jwkMW+zF3m3lnRAbW9HIRFnjH3FyDTUFTPuYQB0Zywu+3yGHNTykWcY01CyL4JX
fl4eISdhcXb3WMV/D29wTNkjsvSGBAm2w8cwu1g1BnWcfKVaGClxFpaplJ7bQp2E
MatQpfW8to51fKw3CxFLaBwrnZ476h5NFiAhKJdkpI6skuuZr5eeSnVECdpHyQcm
ToY/7zLYgOcg/mxVGY2RlG5+Q/EgsqRBiaguRpkwCasS8D34niqdjbsEQTNJ9O/6
Au7NaVDaSnAQsgFjkQ3kVCgaq91Zu/xzkn7iys2350XtqA6d0WKSRPdl8BC1G3Wn
MRbl48FgpE+elotLkBzOfoTwFD+4vV1zk1rQjcBfxePHdCZoZ/bIYkpFyKBe+Icl
iAp/Y3jIxZC4CCcYWU20h7mhrRwxzSMUMvCI93ifymaBRHYvvAZNY2k+YCQF56Z4
sldfJoew5jHJcF79/+5jwC49KYxPZw/5omG7Uw8x9C6HwenillXjZ83nIaSDuBsr
aYEHZajou3+7uEYMq+uVyaxK/IHUGsrAL/skvUeYhKnPptWWV4jGm0bwcTvtwk9k
FtxmnnUwvfisDQ48HlLr8mDdFNVISPS4z6Y7znQDzWkxsVYq1nsnHSrHPnyC0vjt
oSZbDQRBQwuLqUxqsA91HM8tyzeHXdT9WfBzPql2wVYijeO98AIqJGm0TdSLOzev
m/r1UGeWBXK0SGM+5frBLJQz6HadWNGC1pGnT7V12zSy1ZYX6ht5/tOjCgTysliZ
3/0HvXv8RgpTMF9+7g2FFuzIGbB9EMNz+KdQOgtqN0yDuikWggeUz04psQlwLdUe
cXWjFGMeaQkggD+EyX7tA5aQD3SFYyy2JhnkpQooRkYrfZ1zYgAj1oCGc3LvYu1I
H+s1Dis+NsLlD/klSeGTr7+iSd2qxSBa4UR2L+hTpIpS1hjv0QEpBibatdkzcySK
CHfbEwdbU8+CMriYsHtrX6I7N3O7m6g5ux1PtETdRtLX2dtoPYoE+KgUueifPgkK
UToNZP5CqHoR+umEoza5QRciCrutn13B8pTkjArGuQxWyiUTRnalELOmIxifI1KS
3TOsC5aXIp1wOvjJwDDSE42J3JM8lnYbttKZCD5hJMhjOAuq5b0JVCDBRGwtwoYy
ssf8phFcMVwKrvD04f17Js+MN4jllbDGJ2aXIFvCylaIzRGiviufP3kp/48RYBJN
BxZXX445e9glV0brfLgMoO+9Glbuvzl7ZdyHLXTNfDvjBPrY7y/xL65S2ghgKf8h
SHBC4/EDy6DShOkn4qjq3oX0qtKKGvFr3HivKAfdQPq75iNUM/SVKyXuqFbykADw
D7Y7tA2v+WcC4HRbB6mPEhmcI+mg+EyB/a8FpXkJrF6fNtDvqNTH/cbm0snheXO4
NnsNnvCNJQ2sDDVoAp4ZKYOXIn4xy74hkM/WyFo9SnOfMbxHlWDliz78pJ+k1iNE
aU1JJWTXny6NFRnYRjNN/nXltOAzBF45jJwO656Ii7vDumeKE6wBBNWDzVTb4ER+
qNH0w2avQCxMUFJ8tVmDxlu3VSfwDJpD6m0IlEHTYaLwcBRIhVS62OyHViZr0Hc6
7tsBdeSD27Qgw9u9Sg/5T5PwnBuhVpGa1bQ49XFreM6UtRodJYRHbsLg/YJScsFL
V0DMWi66YqNzRZT0cDnfeJsul0e04EewYisp+ORw66n7ugdq9YBIgSSnSnJVeVNZ
WE3r2+rrMhc9PAiG6Nc/ge6a/vLbhRD7LcCFeykmB1VhncMngu4Uqrm/8slWxrv5
LoYqEVZ6Qs2EhcTAE2F4EJ3VlpnipJBiZK+/ZUVzIWF1Pebjz/pLl/iOKIx1Tu+y
+8Wj1VU1ObGtujvZR59a+1PgyQC7nz8c0A8qdQwKcz/hHs5XSuZi1qtsTxxKw9u0
KeV1ABvVCAsJp/z9ixX90mfP/uaGV3i50hcimGKAS3cHjURWHzCN3VtoKrQ0DA+S
DaAaqzm32xNWAZF9KQd3bZWXi+hIDYzpo4Hy1shzKnx67mQJzuGJGHKwR0PS27iS
lBLj0wqUuGlSaLpp0ShhGnD/afREwnf173CRSpV/gxygkuItR07+mz+eG2gw6Vfc
PaNv05SsHLWt+qU5CUjdO1MAFqx9IXgCudcug9dC7GAww88rKiSLX4cKBgxP7+3p
LVumAfaKaKd3w55mdCHsxb2sI3oCRdEOeqSCjw5CRs+lASXCCjN/8JLg3yZdh3IX
jjHvDPu6/UeIkH0RgP/ZEjLCi/ZfPT9ohSI+2ocjxKhZgaUG5VYnB4JXe0B5Au9b
lJ8NGyI8+L95LXRCf0cjy+RpieV682Cg2FE8cT99CCq9CnERqBAYvoTX2/rm7o5J
6UD/AMSPnuYpL2HxwVCn1sQV03UZzzjH38CI+6YQbb11OpMs2HVtOE6eeVbNsR51
ErXNzJMA75924+ZWyMhu5VhGHSNYeAHiAN9xeifUdj40Jk4rvPWoeL72XE4ychir
g4948nEdpG4BLYAzTPOVetCrzkE68Mozq/oZOiM8NAVbi4x+XJy/u3d3Oh4NxFo7
jr+JDZDG4TxE54twguQbnlekUulUsWqpSOzFiONqrxKrt+Okkb1vJH2nyRq9yKa4
5MGUSCx1uZnCtfpFk5AW7pj8sPKPkIDaVyROkE1IsDhuCNdAg5q2/ZXrDkbtJhfF
KH7kQpFfwHD2l39jFevNrznsGWo3ZFL5PjhCn/OMeTaPE0yyxApPX8c3BFlqAufi
w55m9UXksL0uEP3Q+VAoiqavgs3okrTeCmJGLflJn7vJObb6q4xD+qYOfoUnUziP
TshXt3iJdJhclXAeNCPFAxrQZ4nfL0GXk+lCwt01p461EtJkI1YQv+R5H1oFKZ8/
tgM5/D3GuV+MO/Nltwz5oJ41idQyUctUr4UQVVubupsHbZ3j1ghcCUinoHC+TJdO
60NsUJ2EtbaWuQREFVfGekoi0yiLVKehcUo9e1niJYKYnJp/Ex22ct2svmKQIct1
c1faUd7f3AeVyKonutkhjNajzFhqS1YQXHPTndxQIKpvPCUPx1PMhfgBpNSEH2mD
svUdwg6rTNy+3A170qB7hWgxZAx2z9dPwkeMsbzeQuYx3jNNLb4l8HvFGEu4RDvB
IVEXdGr1kG6MhleHDF1RoapEqm2M5QO3kTdDlFycLNCD8URtQq23UWTYjZdXKLE9
LtP9n8rrzUn3InWVAOAbQcUsUtoDC67r+7yQpTAG1J0r1XTrkahZbWr0kSoX+yZ9
/BC/WF3uBEoZCiWSn9nJz1Tjxz01ERBPk+8IoGkSSFp6o5h1kj0I8wDJuN9EIbI8
h1J+iGg3Tkz767Uhz1tGeDugyv1pFHZozDzcBS90ycTwCmuKB2mAquIwkfI5dKU8
Gcyyy/9AuC8Oy5C+8kyeBUno3jNwjM7d/KsE8xX95b6LRIRWOviRXRqzO5HdRRic
gSuAs3lRs9oG1raEB8yqXQtFTsE4zLkGBxBHBB7ZI5CN/+GJp9NfPok+88iFVXtu
g/V4ELrsUZE3zsF4Y0ABx6BMrhiuTGJ71Fqt6CoYtR9Q/qwCtZaYgpAR6YjVVCVB
pKhgoqMZ8orHlaQxVClVB6SJdEKTTHynMDCq8drA/P4vMSAlhaS8dkhmHMYEvozg
MeXKxDBGyoLmHjeghBcoDnLrtKE4VC1j4PWPW9qxkZGzDrpuZOalXvWJVeHk7Txk
PTIVW9G6J4JewqdRiQICyvK2+0qIhR3Lx6s0EnKXhLt8GWEfDdaiLDC+r1KuVMdN
GCuvzUJl0myhPir2aEafU9GAQDKanZv0zHaOUQBtHfPSumTUt3xgCD7qLDm2RPyU
Vt1a9n6PJduiWF6fdzWxUz9k9DL3Ld/2KvbzwUdfuObUDWq9I2DUvAZ3wuVyLhh6
ZivVkn5X2p+ZYSOneAZYLVN/b1AliwsfK5HAUDnTnyzyBVQSRfoELt9bCrjdwY5V
Mk05jNEMG3+gy1IbXegOPnrDafmVjhwLr5S73OHhhnHZsPI2H9uceB1hRFaQ8hkC
+HNH8pq+q938adFOTR6y+bOmmjnsUJaRXe+6ENJ7viAh0xwxTCRK8Wel/lgT2H3t
mH56QxvWvCiwgN+NBlEAVe9JkeyDX7Z+EHmCD3mvlZQJ/7BYq6IGf7VZL/dBJ/me
Tk2ms40g44lidW5FmzWLRm6OF2rutFQOv5KRvwPMLsEGxxtLh6ZmIJzPZgTroZ/f
PMJXuMvX3iNzz2nokzICs1Sns6sK2H5pDm10dw6y63QlzHgKGit3zPeGEsTKeKwu
OBCISWhs9rKxr/WBlf528zKu0QiIwUDMANvvKI0wvj0w+FB94fRbBhV/pwlpe2gf
i/0KyaiQwiwQOqKlIyj5H3uGj6cB0gcquC82fCHoTfLO5FNepGoT/w9Q6Z73PsWN
IoIdO+kPai/iPpu0Jr9Z/Zc/5gR37tVIrgtKAnihkRG0o1VonqBWMk3Gnu9tO9tT
8tCcQAT+E0NAjj6WV/o3bbPWLhrPVXpCYlpMwbqu8nvCWPP92Dw/Vf+8d+5dOC5x
gCdvn7/khwtLjaMaU5GzE2kXKU6o9yURfHj0/VlGcDB5hf3nBHMgwQ9KixeN2wBd
zPQlP6pbB415CbPgrQa0+XjlQoKSJ3zu1gWWIJYKWVXN4eMxtc0/CyV5RCjl1vPB
qyCadjb0+Sq5oqMwv61B8odSffsQN6kRf8jnxqJwJysF6Qt8uTK/K9FfImgLgnc2
0fVAastHbuI8KEVdUyB2t6t+MHwpOdHcDC8JBLevz4RYmZLplbfHBbiwFEnJs0r3
xwt78P6dk2UCo6NKA+yQs+FdKaeVZ5sJoAcfYhTCb57cbIo8QFiBDbwOe1ZwE5os
DkC/CfjnV++YjyQFzuXc4qWLC26JjiQk9dP1esK33mM9FI0WVdLLmseapeUl6wp9
o19nQOoGBhQHn3jTmkH67EKsVb9mWKQjJfUtT4Vj4Uh7EQEQqRBshTA+ANwOhzxe
1gPp3mPSjEKkvY4jPObJ/fsFYnSa998m9uNs0ktHFWL0CCaAr3VUMVkS/c9WX8Ig
Vmdrb+8Z3y6RgBhwe/c/okOzB4imhzp2heVq0t7VmmOD8XUuwSyW8456X/azLdB3
ILwWYXiY1uN3WN6f8f6+EcClCE1JlzK5uws7TofNVsxjzc1U1L/ZXc6n6mVdc/mi
aaSUZsMOZXh71kkOPlRXrqd0+BWHF5JlkmpZ/YiMiKb08iC6muUQR0KJoCb1083g
PecsOAlnkIvg7i31weLSt9r1jCviwYAb7QZh6qkVO/Xsq4vGfYzEYFahf8/hy8v+
6anOHjd2uaddt0lZnAHHIg+eXfdunIivP5/Ygl8d7UEWqlQQenr5qDLV+KeLvL32
ctVx4Q/PA5jAQ/EOnpMjy0ouzaQ65R8i6sIZbrxlWqCEnKYIDCG3ob6ssDwOEasd
9qo6f8B2qZdOG1XA0PWyorph4+mJJ9M19ms2+2tLWVnYjV/Ja49wu8zXuYoFvl/f
R+MFUOS9QN5aaVnDyODV/emkOlAXg4gj75G5q2VOsoERcXL2fiNBxOr1UFm+EUp8
Mo9aVBNDP6XujQGufrCwTVtpXK+EGG74S/Mu43rRZaenqUsjKGCIO2j/Qyy3JKE0
MmW66o+k+cxjqC3+nybJx09mrIwYkoOqO2yyEpfZPki591FjSP3Flo0/RRSxo6To
TjMuT5Sdeq7bl5ZS/FLpCTPa0ne/hvNCXSc40h81VHQiPWmSO6n7pBJHyF6/qqwX
pJWey56I0EDSFk9M4ySfNDOKo9azNzJA4sA7NE0aapFlHbhc1L2qYr0LKlhFUUQH
Kgsynkl9+BjmkCwN0D79u68BDmEs8hfAxvJ+3yoQT+3kuDfc72iYRVIUPP4PxNyl
Pf6QFOBjcowbvY5t9i1ahzzOCUlDFzzLLo2ALjRZDcydxwuPcpnLLfCoAx+TJJGv
Y75pwc2XHxfN1Qtx4Sg6agHfXZUseww+SDxEmp+2+PPCZte7VaCSawBNOOuNxJ9P
5k+kUK4ihLkM4yp9Z0ZCvxJC7Tk+pw1w++9/ReawghpM8HMjD4pf4xK+0a/ZmgSW
E/eAxglU3sK03hKyI+bzy6Me59NzG3m5MX1/zfSTwULU4i4mIrBo7kydds0HXj18
CpN2L0qDoMdrnRQW99kE1c+YQvL59WVaN8TiwEWQbMbzCJPSzkj/bTjkNpzXPX4n
2JDR2lLSgZVl4dQbJTT2PPPyKv6hh7S+xKoCGYCAXsOeKMcK/PenBuQc0Icl/NXr
AL290L/56PFVEhHoycbsz9z2jYb7QaVWSU0fe6tJJ0k6sh2i7/k9hqp74UxRKR7b
eDlKOda5AFdTeK9od2ZE8hcrhwPT/xGH7HDl1Yu0tIKqUWDAILt8ZAbc/3y8FzEc
ltCGEYmh0/Yu0/ssxEj5+CKrYfyh8WK7T8QZsiMO9I1H0WufSwX6FOArpvj3ODqy
93RF2rr4lAU/m8mvVr0cJSOin5HrmsiODVdOjiQCJ40o34tiUTQiojrQeo+Vnkhn
6Krl66M68GEI+w/J+naHc3uXK7i5RBDRYtYm+j7VJEwRh/s3mVr0Do3rWkXh2on3
e5uyne0belJEduYboLU34xwVXcStstq+BvxNq8Ootz/ESZGmLvmq/Pt7xEiDgnEX
ysVYjPWcDcfs+PvS7kuvahlRVGQBdUh9DvqXaT3EXGt5uoVXFsvIu2ySTQiAJyIR
lIo9hlihxZw/hUxa8Xf0JF5nu1j/mkLoXr4LgS7FqCuFrcvRLi1jIBaXoO1Rjaqu
Vf+r2Mi7+8sA9eVA2NMI+LV/glC1wRpehruUtG8KRQ5V9mZhgA5b1t+SZrRpRhtA
nOrGHJXw5uvrd424KBOCAJG8sK//Rrsd/BlH41fyg0fdJK1RMzbLuvylS4/bPcL9
ZjP+XEW6+oW0YRnrfid2yp7GWk9GsPT1PiXvtId9IMtfGyRw7ZV1i1k1Dr3O20xn
XrPz0BejgJQm1ZG35bCcos+bUukfAMdpHAMEsQJ0o64XKAo5PjBW+d/RCrbJgVyf
hhXfnzXxpMgRWBmlQK/gWqyXpzayZg/B9B0aUL+h9yuR/2kcE6j5MF2GHLKEsPlA
Cpjv5ez2qo1Sti5/FoK4aE59v7+mkhAqEMfnziWfnzHEWAF/sxpxdPFTlb31ecFP
LbMbC+ZXrnChRgZ6GgaT81U9cP8TRjkgdFPmljndS8afpleZ0n+Jz3kNbLplzrz+
4t40SPVu0vSHKD8Xeu7PUgRMLIuv3BcrnP8uYDm6qZu0DI+9et/BvOD5L0UyohrU
JESULtP/F5wDdkazzLBqr3tHCBPPnCWeF5LI7G4QvpV9a5SDuoWgC5gi5OY7GGQG
FPxJF48tF+soIyCC+RtxrFa+F+Xp0IhhFx6SZakNo1nit5LHJ/HNV9gQAyprCSUA
Vc7G9NCr/ipCGKhVo+KSElMuV3fMTnke7QTenF1eRMHCxsGmzONZAgCo+pOyPEOW
46iIZrOdmaB8f8vhDETebW1DJu5LPovppAP7GsGdrkN1kMv+1VK08WqhtliH7llE
JHgs8NBHnPXwd8GTMr6mjDiu5/cZU2x75cJyC1w84iT2fUSiAEX4vnZkwdSdKrgO
Dh7qLWzWgPKiSXd6thiutGfCUlDjj4HajQ2S2PialWlON7Z03txZRZTRpinu2V93
FFt8vKj1U9lJg2w+K2Gvp5HKi9fHNvc8T1izTUR7eVPhs47YDbrbt83ngiLBnqgE
1IOd0B0DE2zGNnEkpqunk7rPhyYHEpAJSfkbqvKXCK/NfvH+RXiDMFkf8hT/lP6+
lt3RZXLPPcAaCtwoFTc08EstzMN5LW4Z+A76AXa/bh7CqMWxmds7cRLEwp9RtGPZ
qUbedje7xMwhVZ/rwauAIWh/d+kdeH+ocXGJv6CZZazhHuWFzmZAZ5X/N0Snav0o
UQ51Sry6xzcr0QCCYoD9VK0krrsUywX2xep+yjOuJCl0zw5m2/sh3EFZJbR1oRnI
EChVGTWd/2djVQ4ohjEXyA2XQjuYJQl2KvquUSg20B2fzQW/kIUxnSGSB3oYV+6x
zsfVnZTX1+fsK3uVwKKT3BgnRUoKyJiVW78EmsQ9XdrQHye1oWuo3L1k1L0VmtmJ
+uMK8o+Isq2/AD29oNKCs4r8MKvmu4eKQOLGXguJb3lTxOyOcPu+drng8L8WDfpm
kg1X1UObsumxsHU0ryVocUNWVDmxWGbH+qVz+ppjA4bEEFv1aNs3qm6UkkHG1S0h
lqMZrQ3ROCgj5GmQU8m38kwHxfZkF+KgxHNRhYxbiiCpsWlmzG4nYmF1kTO0RcJB
7VJxh5ycXMCGk6vV3mWdVyWgH31Fm04DW4bVmFQd6mvcQTKf9JRZrG5+ceD6LORD
JzfhJIraDVUMbICXpAS+EJwI1ahwtV2MQGV7hSGB0EDLfZCsVoO+8ze7/sJeFQqo
UeYJbs5Rv/WPORkDhUZYOuhCK1JZ8SVc4hGevt4vxIil6+VxSN5jVUlqsJbBGGWi
n40S9HXpcCCSxnqvDtdiMtKhx4tZNBDJwsTVSPcfv3+m+tBfnHX5vOlUtrjEASzX
bqYZ8VWfX7E6/2iH5lj2xONBucqD9l+4xCvW5FqXa6zI9oIFE313KNlbCDM5e3CE
bEC6H7rebnW8txGYvHhbSQdarAxWA6S7C6NVhz8VLXk+NyJm9lBWhkOENUBh7mMx
UtZckJNkOCKK2v6J5hvieVA5q4nQgcTD1vaSMF5G6O7OEc0dspFSF8fKRF6+Hgdu
FDYaVLKNne1bp1R9m3NB3mezXO0TdoD9gfM6CoFBl2uYyzhgAVnN3hzl9mNCTAFo
XEMfX4xJrqNVqoFBlhjdQFKJrP1yU6rdrOKdMCwzfpY32knuEDvFC5wdoR1Usi2E
P4XkzdAWso6yYAJPePhL2Uzd7JyuDBLqOFr+VjLd6GzW++JYXFltuDH6XPpMUS/2
r8RevFuR3Ph4G9qrtRKNnxeU9Ov8eXTb6PQFvtPMtePJORLepNQVOAKyU2uQb9nc
fZ0C0ftFygmNpPHLPnMdEmqlK36zBN1f9NR7QoMayf8YAsrXqfFIdGcidBUleU0F
3C93WIVAwV2Z/1JS3HXBoe2j2u8jn1AhChLt9JuSabjkEoDrpFpI03FM+o2uUBMt
u8MiSDZET12FZBBMA1zoGlJ0rnIQ3kWX5YbB4h2hwxd2ADP6HdichG5kUexTx1s3
Dy1uccI5Djq1WJHD7m8QpmmFkDJMceqjBAtmWLwMySLqCVv1g2amu1vaSZmGBbbX
jVrLkqYjI91J68a73/tXI3J0Gwg7DLJh+gxZ3j1NpkQsIiTD3qnR/FsnxbDGZqQl
1yK29f9gRAEcxGV11mPd5+BULMK3oLlf8Y5yScwBwokOtgUT3npGE3AbLfZGBJke
eIS3RdI70VYlMjgiZl/MZgpWe84EQ4NruqnXplfvIPK0YpgRkerNbVUK1yGM0mAJ
uwvOfpMdsUT0idrR059U84bW6pl62UPgle1gtXsxeE9K+AizIRdCuQG7i+o4Y7dd
jaXJszP6o9M1QzStuduBN9CA1ZDzeU4WCD6RgJvePtwxg1lV14VXpcFzgSR3m8EN
lDu68VArj3EiyU2sMgjH3pudqwGfG6bIfM+dxYQC+RbJfPcc57ucuvKyybdEiwR1
VJ2TjVU8pDhBeSWvFdSLujDz6SDId6vaU7eZEnrd6tx99GNHqIJ71UjiGz8o1bno
uWXnqqxAXUSHwYS5bUAFoarf0gdEcnFLFhNkIQeEwQtWoboC5ueCT/Orwf9ZCC29
DBeR6NWMhn+WA+E5yh60B1jWmJDShJXAaNjEhN5awBnP0zPx4mG/+dzPQwcgmxlO
Np3lcKzEWZ0I94xg+CpWT2W9lqofO0+YBdNwZoa/au6AffB1TnW25Z2LPJa5MRoC
S2fYDmvhflOPC4qMD0p5xnL1bfv+VftH39+aXF9QX5z5Uwh0ze60jq3h+uVdTFtB
2zjFVgYyEfwsMAK2Ez6w5hFr5mQJ7B5MWb+/vXOTvKNON/upzuN4lvA4MOrzugGD
suY1Ao62z5YVZrjNGbHYMT21I3Zdfs/WLc1yp3eo4t++gV5pX7Igxc1EmDteZk2s
p/VvzkuvPEdNMIIJb9S+HJO1j4I/+MPRcAGG3rlsFtL+Oa/8vcp36rOv+orQF2aJ
bo4veEprsyPEDXdCxS6LLXbUrQrYoh3eJjagjb3/TJTFA1GoLkHd6CywbTGj1OfB
NnfrltBAKDkQ0+gpybSM9qtyDLcTiCtRbpY8LrHvje0JlAVw5zoFbeJXaObAhbUA
XKZ8gXPAwQmtL9DuRvrQEgcX14hJNKHjM0PrPbHlYefM7BaItc39d9O1YwJKf3Y2
TnB8xiauqOPbgbsHH3ok+C/46iIXMHxNVWbIIO8SLdLY78XE0qqzf0YqeN/1WvNo
FO4INM2uHMxcSu623F2Z4D5SvAOZRH30C442pQUudy+ZG49I35xuqKyPbI/cG6IC
okczE6QLFbpmAJR4+q/WcCv9Ugwkbw7trfiyvGojSJw8x+R27duM5GX8awdmSqAa
Y1YQ+xT7Q2gQx/1483Uo+wfuKzueUNR4Mm8+JOd+hVAlxHKbFUw/pqF8pkH3aKPI
dpyBFkD07yQ2vFUrczt8g/tnnF3u/yTGt9iSovw3UOPCsjUADOkUUZ183wk5L9Mb
f+AspUztsjnZiUDEyFpH+leyrdptabG9Ve26vvHiKFAo7rkwOE6RTKbFgj07VLwB
lBqlbNCJ6LGNC+VgmktIE26kl3zjtbOV3eBb2yxgp7/REbI+tIVZ90ql2gRfQvcl
MLZ4uRMw2il69xn9rm6oSsD95i6gIL2h5bJhXB5rRSCBApCpsPx6RAwFmVdsV4xp
EHZsw9doilpMroENOMmGvNQzFbHHyZex3JDrP0/PtcD3DsVbp6LZuap02SSq9uo4
TvPwELrDW3S/oQgiftNWbW/AUkllJav/XIK1uTqQhiJAFpal4g5zz4NGdfw2abig
y79xkrHvgTLCRVAFiMTKql5yPtlLOu8fSklEIhTEWB9cv+e6hNV/zPFxAey0FxQ6
hnJx017geLJoKctr6dcGsxKcvbCcsOooJrgm/dWt1yF+lmjwAuPCKkQkhS6eWJbp
zRBWlhauqXRJRQp/nCtxBpu9cjvZiqWjnhYCTw4HtvQcmMrXJdGORAaXsyBM0rLC
vKxbeMVh8ZvNIx/rpfrxARxEU1JFBqbnmfo00c3Ts6A24OaEEAcvHxXY/1YQP3JT
iSrdiPrsTwi8JHXPIum0V6L4Qy79TewtrFroxRjgH09fB7W9JR/6ZiXDZmlug4Vq
1fqB3BxRWWNSIZ0LT+jvHSsC/QGSPea2kvE7sX4HbK3QKnseQIeOI+45m5BoZ9jx
3GSriVBX4rBvSGLClWtESJL58rji8WZ07W8vvySDh3bHSYEAsImvhxgLOpwoo2Zz
ZdKribAvk8xsxP35zLGCWiCZ80HzdNKmCMdO+Lm5S9OZWXgGwCJRYPyd5ghLh3ST
+tisjz65BDCo00QQH+x0uH4+Bnx/pxyMSI+/qvQgGu9mxqtAHiEEesUbzOZqoNff
vlupRmCrbU7kd5OeJ2nukF1Ke2IB2oGNNjJ02e0lYStRKr+A+qWd9hHBn+nh2J3o
3mpMwlu1vD4kxOnTszu+YwpOWu40//AZBGx3ccyFWB91M6zMxxuSKKeGVbhMhhdB
pFrzesaZloNvSrjpY5v5FNrAFUTWP/fvJZ6jjHDTd5R7cUPq4B6Tf13qfUSpiLcF
RWziHToBCsLtdmFj+Ck1oisJUefDewHte4RF99Hj6Y+nLapJFE4WbWUmRL7oF3PY
91gD7O5AwVIE5jQSKxoiQ6Pvu9PW5LbeHCVKHVtCHVMAJ9AhE5W1m/JRu62blx13
sYRpgxTg7CMjuPSA/wxbRNdw2gLZRU3ZFf2djpMxDQ+jXT8U6sqhPloaNh2Am8VO
IuuxJ1jaMUau26lheaJYuSFg6XQ9IwjTlvK/DmjJpjIGQp6pkMhfQ1yIGuW1N9B/
TuqZMKei/jwWWWn/i8POModGVy+/hHxtLSWzNWU7em9dUDHLNbgKLGlrGaYqxqqD
OQaC4FmqXT0r/x2m4ieYJvYNsrVucbKtQ5Y5a2H0in2HDivRTN8YuJvlVP3DduGV
i6dM7jTDPPhdbkKicU3o6HPj0svsIYnApaQQ/6/AgUNON+b5rujIz3z5a7aIDW0W
S49Wo5GqsYpxldQcXZiIMybICycx8LXLgbw5Pc8PT9kEOO2mr3NgaO+pMg2waGx9
k0DVFWAlL/YRzqyEubRO/JenLN55hIK6GzEKxdxpcUj1zYrmXvd7izv7TQbru/q1
cUDPs/+zv6DV4ad+AOEeY2n221UKSMywIuhK364YSlXIa895eyN8XWy/TCRDYmPd
WTIkImWQYP/HACpU6Ws3Dgcuxmk2cz1JNr2z+PWaug4pM0bIgnn/Stf9vKwBH8Jr
IX0XSTNQjTdwZGmJI00L2hUC46dumSnRKU4r1OsEqt7g2zuhXd9Y8ws0Wjfbd0SV
4V2Joi18X/2v4bJJ2eiIRCzZ99IwSsTuKj58EoNlOgDrB3H33e1h6Y9zG/qv5mEA
TKstsp3elOz/tIyXqIFRhgK+tTdZTY8JdsDaOldSaA3h0ZT7J8R+vX0g7kmeUH/P
lW7aEHs/CuStoZllckmp1uGABrp0VXrfKbXwhUEb/ZnUfhteykNluM6XJ7reAMgh
HUeNvOq/Q6zQ4O5h9dvOGMvs3EdCxWJ7VXnDq5FRGf2TuQkAeca9qbPYlvS3ZIvU
97tr48Lip+I5JXh0Oj/hM45f/04TE2MEIbBPsnFoDf3ifX6e5RkuEHVfFG1bzHTg
cOLAOOmcnsWC7xyvd0rARpo0RPkZj5LLRiGoyfOqTAYQK27aunRCYaZtRdtIoUQI
+tIGChAKL1Ho/Lf6rcQZ2p2fomQsR03s7n6ZpjiwO4/94lSvYwqfBkbxQRpMwJeU
GuKPnehcfyevT/MsnUBDqmW/rCzt2PtV4mNlchVYSBdkebINDe5R10Jd7FbhIzTh
blBVEL290caX6dyi7m+Q2ZnoJsk194tk9o75aouSnpcMTaPYyYd3kb5fadbUupse
2CRyL1lm2/BdCaHp0arTy2qQuanJGY8IDqDUP6HxMPIpMsrTr1tIjbOU5nCd/KTI
BbRE8H/mrrFAnX69Iog7HDguGVaMMsOEK0oOaLNLnt9nPMF/GhCkH6X+juwSqbLR
tmvPDS6vGMLmlq4aOlf4PbtwAoaSHv5u1XiD9LyE2Rh1f/VNvGQb3J/qc2ddRptl
fNsTX0jnhwQs+jy/yZOkUXVtICFRVRJyKzXveVOI7oc+nI3eRaTO7FT3zLM1/cyB
twe25nJzxlwAJb7bFblxbA7y2I0qQhxJy8qc0iyrkKOwz33OEctZlXxjXwI8VtCF
LfK7GWDT6n9j/VeFtNkc3ouErMTFJen7w30AFUoQbnkasAxhjoYN/1qosnztp/MM
ZK5WDA/yPi4kfLNHLUI4ZZO04RXQRVhgcBSX8N762KPbFv+MkvbgCsnavGyVWbun
u1/y18AX6JFRQM4PO41IvVHkcMu6PtcDxPGmUka0VQ4c/LXVjBc348C8bY0vHkI2
9hfYgCcuo6jgC9IpXCo3MFeKAZT4S463RRLUC3AXUFV40PYo5ugps15HxACZztOM
hY8g0ePfrd3V2L9Qsw/mU86kv1Y6KwcCIp9vT3pW4Le6b2Tlbt4E/H1dIeFo+6W5
/5d6HTzn02pdi2lJAIyJZ7NjpfYe6XFBxbawRG+WJzNYuYBVTOavmYOrlC9nrbgB
NiRcUEEfbTjsMj6w5pQm4FmJidaUHycy6hy3DL8lk5lG5kHqMrAUTrn3dAS7H2V2
mfgZjA+WUIrrOOmZhUMVvBwlUh2IfqdDfczGomO7SRUKi+uTL0z+LS5ja5rnhy+/
aQAlnyNp6xv+twgfxbe5+THBclQHWkVEdAxcb6DtHmR4/+sTEXL1OLa2ZGjmp7jn
Yfb6B6SebUhzoczR8uMKtvEc+iLcLy/Ai/6f2rsos+GvF/1SNDJB6X7id865WptR
fkEvxibWIUlLpmPr9J9SNXLDxe3yDpIoaqibarzWfTfITWy3QuG/sq2hJmDagwFA
unxN4uRFYv9WgtvWijEJvyh2TGG7nrZOyXwQMO2CG7Tw0FNrFo1yQSh963X73gcR
6TldfqHK12/toUOWUAVxCjLMOdcKGlA/Ce2kCZ4I7ql911C1v4uztGoSDehM9Aki
UXa43JeEJkdNFGs7cAMkqKVqIurDH4H2BZkUcLvOXkaSdW/4EjXYJeX+3z5V3iev
mk3I0/FVKyZENfMactfvIZMl5d1aA1goYfTsfS3srKk837Ajod81REJUpn8naP67
UFR4Z3MBe5UwhZ9iVoodqCqT6dQsvvXDKh2rnH/NzPlNLJsSC1RnLQ+rE0sjoOH3
cGkmVMIkt8uDSYxjAEuNjj2+Bso6NJyOaaQ3/C9WTKJpqt/oQHMvLYf2faIqnwUA
3JcLx1zB8JO+T/+wQNMC4cNgIKo7ToTxs4ZKQKq/G4isXCfICsXzdNdDHd4DqYvL
H/MgZjUocjHaTY15DgE6NP0j2KtrhP/2XzonOJ8g4WQeX4pxu+NwoOc9j475aa9A
YpQeJLIpkPWU4v+gSjj/WC4+nHTgsE3HEwgljV+oMnDgl6J5STsa7V1JO7wG2aDk
YzNKeqwF+QTvCelqHYvu+j4Js7sriczzLSxRHcY/qQwY/uUDEnFf5uxbHU/xaKNG
kJYAInFYcbdCCa2xwuk8wFyoApT5tXSZvTdl0h1nUx/10hgrT3ZyGCV8OVBzfeXs
YzV9iLoBBeVDUTWkMArlKTzMIwaRynoNfXZXcK/y4+G/xp+PGNmprEbf2L3u60Kq
wITXKI+ph+Wap91qW/I7X+I2fcfFPPTCkT8muCyxWYvXMzPuvhCGI89fGxSKQBYX
Nh9JhXpucjTLZfW6WyfgB75hPt5VuPoqcD/q/U0mWYua+54Q3zYOznv6fnHSnj6t
+ffENvvYiQ7MUAglqBCA5zfjKD8mSgMaC7UVsSRDW2g6VZQ2q9oKj6T7shLAErdB
3Mpef6/RrTcu5HiKOqGzLLWZBkpm+pmjFK86gbGkXflUKV5wjd0ZkiFp5CRysKHi
M08tymK+xjciRrD6nFf9e1IbQELjpL/zX75yEvXYcGQJmQvDroUxrxkHl8Gm7nNK
shS42Y7w7mqBBSFdwuzXkz/0D32M7IID4hzwK0ZHwNl0pWa5SUkXmRWwTTCzFJdn
qgWJoh06BGzWVrQ0RJIBYErTksiBcCQ1dA6boZmJhDgEu8xiqRIcmv1s2Zt70lm1
32N07mAdYhK8n+1rEyOdJcXwVvT/wwKlI6PCokwsMKEfh5CGhiRYxGO2z0N5Cmix
DdfXOm9TGicOa2pwxnJJETdN10EARjCmZRbUtTXSCK7Iut7CpMWKU46OARpYHHIF
CRglKJOKl1RnFaxYptdf/uyvRYUO3TwZfEttfB8FhNAqEinnz4Gzyc3awWSyKhQF
XbnQr9G8Wp3IkUT0w9ikWswwr2Io+AvpRAIkTrC3YJ+kib5IdZkLFwm1LwnslYfx
7CQoEL17BUOaVdRI9QLKQx85bsKYylDE5CeodbDthpPLIq1LLdyNVUazbxKNMR2m
HYMJY30qYJxpivZTJPFMAVPXMRGtKTylwi//xnr6fyH9D1IMKF9F709cjAELaCL+
hK9AYlEdJ48s5gd1QbU9vfkJQ1s3l5cG0zjGAY41MgSwYoVJm71BhwAQcb7oN9eW
QYlNvM7Nwm+cgS5AksqaGXjEEiqL35hP3IUVpB11/m9TpUfio6gGTkUXQXiBVZew
l4h8LAIpKatobErfSyk990scWFOWu2USksKwuf6elp9XQ5xpo0R57gADlnk+WOVZ
asqUl+CDDlylM+JDKH9U8zPCqMUSkOp4CcOnVh70tjHJAoIERWA7R4aIKKFjkHiy
gyY/jE+c1/yjR/KEVcVIldO7GV86n5WqSCIUOoHPhbbGqn/sHbZziKx3u7eVvqjl
kKmR83PwcMcM0FEJvEC+D1PbBBjvH0wcKGQbdrss9Hz7aAnfaLiJ9nR7xlAiVhug
kPPeTcdMrmr3WEbl5RiRi+fbEy0IetrXGfDdgHbAtOgS4PDCh3wq9F+n+pQWkH3I
Jjx4DK109XKJky6a9nBoexIas1ao/Bfo5J4WjNIUlkbhX/JGlP1rGqxNn6LN8A8o
8fIFd3WZAIx1mlQ1pEXH+bcqBVUhffoUepMCmsXoPW73KOdMibJYVVJSpb5cN5Uq
sNxBNVgUcrQjspQH5fObdC0Q6WPPqCa1bGfZvUfh+iCrZ//o8n7KdKJUbqN6gx1+
GZ7jdvj5WKaQV0qn6C1lcbiL9zVbr3o0O6EUm29ywAOGXllB8cvQm4IN8K+xK+EO
MpB3qZKUfTEESd4CVChwLpOpOXx9w8EnYFwEx+26ZbHXauteLTr/pk4UtoJmWxuO
i4nrsgBhQ9SWDQyrI1ft/MngFk0yavN/O8Fy0Ow32zmsAWvTtALUJncr4RxWnSJz
kl2+xiFGzMgXH+vR9FbcQ0ycmJ8WKwyjhj1O6On/NYIjssyGQFA2o+ral/kzDz/j
PWv4ed844GcfwNnEhIPUD6IHue8lGzIlkJJL1JbeTxQPaqHeh06nW6a+M3aMSZc2
CJXtk1RvjLx+B7fSvufO+5b94C8hvb9bqS995VthwvikEkt61fMNCWM0pvsX7pnz
F8L9/FiKxw6adYQcUb1CmPjKX1PaWlmUtB5fholw8Y1iNeXIzDpMea1U4hay96Z8
O1L9M1hEczLN1UFaftGdjAygVHhwK7sM3KEutiQcXaYP0eWKfgOfGybRLBGvXaNx
T7hVSy9CSMfOBdNIfKu44B93uzN0Tsh33gEJMPAiej0fkbkdNqwpFnqsGaoZX5PR
+mK9fmz6JEDSCWgPXFLwUKeQJzDDFn4L2tomzJbE2Hi9ugBbTPcHv26ULb7z82Wz
HzeGtKHX2TNnEji9xwrRhxvdfI79zI7yg8ZXPmitLjGcFoTUSwqR9nVgiET3OcG0
EkulXS3JtnmnkCqMBBpnn5fEtJcy31hyJ3SPQ4ZJgx99EY8f0upyF4LTaUXqxn0k
Mx5X3J+ob8t+HAJoAZozGFycWaNcyGztmRgYZ6QugWzMYnUrfbcW8ekMX/u/5A/5
W1/bD24vIkEI0JNGRw2BFEHs4J0hIpTTMugdaUyzAsAbc2OE6s25OfP48/EugW/f
8EU1fTKv/I1WoBPGTeLIlVff2LLoU1FcLhsBAFRRXcT1Xf2gwuNjciflLxF1tGur
HcZkVwEgo937Ze1yCJQlPQ5JXYeFoJtF3zYoVWjmLqNrKr9hQnZhM8b/9a99S4aR
zIYJFzTsj7Q5hIVmZwzXCflnVeZ983zYi4dsfYWfqj7L2H6CH2bRbmC6LzBn29xz
6hrX//4QvG1gH/NxrEzATERaaf+bz2eh62bKdz6YCNvnFZG9MzpqpzPp1qdsytk8
386QbpVcHLUEsYhjs0gYl1+homhEAcXMkTO/79X3+FTjkqr929v3FyAAFFljhfWo
QHCuSi29/AHGzr3SwbA/nsq1iOsFfn9aoIaGt5rBTAy65FcttT02oprWHfcVq+Sh
MwNcwsKAqfiLYluR5aCo956SJTqE4R2xyh5QT5odWjhEk7+XJsPdOmoUXFUATl72
Mvg9zvwGHnxGnhpBak3fqfVwXaENxomaWH6eefsClRX+t8iteMRLO0/b15FQ6GMf
cbnuwduWFoy1ujpMW8vKJsRFoJdgQqVpQTW3KVncts8wPnYqIEOEun/h2RKWNn+D
Dte0xDrFJxwCSuCBj2yOEAu8Jiij/6c3tbs76ur+528/1TIGwHNJQjd+xeI+BXgC
4VJR9cP9nXBN01TK09fqN3EJhQUSv58ZgMHa5UkWUCVpoxNRmIGz4Bjphw0A7RL9
d8j+YOCBeanEvfFXlJj6iWMDq4lG37WMhfbdl+a+FIsdQvlj5ELaPYkkD1zJ5wuk
HdudVDZJh1C+f3ShdJrMYTOlNBy1cTo2nVR+GMGcBVlBgbOLBeYOgPw+FoPoBBHc
0Bkly6Yj1qKVVQzXQcawyxWRj6tFMWBnPPyr8ELUCQfaty8a6LWAMhRKnPQfcB+A
Tg/lEaqISyOraA3Xsa40PLAGBCC6yJC5/9vxO5+91BQeOouuY+7bNcWihDWpaj/u
v3eMyYudKUjzzTMxjzeoZKXk4Y+UnBMUj6RDkl88pGGrZpbY8a58m0s1C7fah+Lz
e94R5JUpiEZLpH1uz2hlbdwVhK0ARRGuaRKUk7rvoCjeVvqbOSRCnqsgYrJv+iSc
CKvqnCKtWhHwea1VNqWHp6UbAV8NkJLKDvZlPYZWWP6svdX7py9abB6eg2RwLHKf
zkHomLHcaOxm0StSdQxrON4Xfh9NpCEZmcENwk6bcLQH7EHljCpMtbCvtG7kEw7P
i1aDwsTD5HIxQD6Mr74upDDfrTUg+9jQFrHU1TN+Qgkx2bUwdYjJ2EuhB20pIo80
Ws+wxJc9OQ/wL+J2cDXR+QK36lqyiI+4inaq1uX96LgscWWRcDFy79g6fluv2xIW
+jVP4DzNEudRS86+Oaq8kke1rc0bVSOiMZ2fOru1+Fhm/k+grgwTjTZJt0RHbTMR
V7TkQpwz1q7WvbsixOB5WgdYegr0pvxSXubLhZm0jzgDgnmq/4Vr/wE94k0jQojm
AhEErTK0y/AIknYpnBFCgP97zoMLfDdx6wzcxmDjF7IFcGsoyVIYZue5jKjAim+0
qwt9v12C1I28pLsspyRso2P3HKi56D3OVYQ1GruOD7/jaB7JG5xF5Y3/n77glTSD
CmhgVJRMPhlRkyj8uEvunCX67Hw8kPQXT1HDpsj7AnjBk7QADzTAbFqecq8vrfnA
dRwMVyp8u0DxeTvr1k2oYAj44X2xrnZVQDhCtNIb8kGwKrQrz7VgN01C1G0Skxsk
6pFOqI9UU4VKJeq60AsNb/ltKmCQASkQjWeF5PRbprzr2wXthS3Ye2g38QyOUVS4
JabDZmfHFL/Dm5ZyEiHt/qPPR0W9ja9Dc9mRbn/Lx6Vz/ivRjtG7Nl7xwLAfsAR4
ULoIC1wc8X1QqvlNJpkZn4hBbVdD9IW2PnlefVNEr4Fo3w7FJUTrpryRxhgn7Fmm
2/9yQ+LLZfA6J7LR8GlZO5Y1p8dI2uefEDJxKr8YHwHvuJalvWbdH5z6gfDXYI6y
lNEJQpim7W13K3oxXq+QCPPs6REDGaim0g/RYfOkorVBbElw9kHZdVAxBLZ8snns
pzxZMMC2KWeTj8CITQstdUw2oTAK3OIc0z103O9WmtJzGOikqoSQzrYfUdylMHoA
O9B7dti7DLod8XIQQzIpFjC2OPXgBqbF8aZpE2GlwYukkjBWrb25eHh3b5iz5ZKc
8t4ZlXiyrYh7zo6BxhNpMctpsHz7XM7+/1/ZUnpsSssZjYsd/kKtMYRx21xpZ8c6
k+q8m78ki2VAAwSQU+U9IWgOPxEJDTivKoGvh2JLQw1o2aKiviyDaYlGh7UxKIMc
7A5Da2oZDbfydESS4OO5LNtqbUv+o+h3/Uv00A6eAeyoaz+5hTGKHR0HYjhLFUuZ
+QiPXJrwQ8Fmo+88yT8GFIk+4ANDpPjNFwdMjmKVs9LWwPB9hSu5sDaZRNT7yTjy
q7aHOQ5pAehePOIgFsuOzIYMtUNck6Nvx4vZr18hYsRfGXSloEL13vX3L8hoQJZa
zNZJs+DDc5T5/flR6XhoJzs6FK+3A1uN7nxMq9I378++fnqq+LvpkQmtB5k8gOai
LOWRFaZAxgKXjc16aCENfp7CtQI6tU1x36pPBvH+0qVa8k2+0Vz+xTb22LA7TsMO
r064/PWmVaNfphkoK9UESiacADHfNAh5QYnf7071/BRzXNHUARYcC3gAfJOPsHsj
O/tW4XnAzTAeNkxWWu3X9qTCi/bloxO1ZE4Rhbs6aqLo7sa1up8bx3OGwiSnDTZ0
8kH2HCwA2krdZFu+l7AA5vTHiwrRPLZC1jmJQZCHjKSWreLhOv/U+5eQVJX59dfZ
sS1J1DqwlQvHbSLTqdBbp71wjsDMPWFRg0E91JFMybH20x0pOm//T87FewdATSMB
F+ORGY2Ov02bwvckUHxah5j7JNXWgc0UsJGwtnLVk4UHBsUdJVKnB5XCYt4McUS7
72HEiRc7+QTC/4hBXwAOWbJ/4kk7J09UQpeQm7SdEeWVVKQZltOCmtYtyhae6kOJ
HjF7Af457/i5Lwu2w4paXviVYd+6lpXAdHGBNeheQmTMFEhLTQypMRg80uMu+VVl
s8pbHmK8pkbu7S5B36P3oCx3gSlwRQcYTp8naWI7w5VSOly1GLgaNfrs8t8T9AKi
82qsU76/GvJlSY24r7iSgb+ue5VUvk3XjydIBT5rB86BAhZaAFFGRtV7piHWBZuS
R+H9ZG1HeZdCJ0gea0aVw74UjnrWTmc8g5aYEwdMgzvn+TPsd/2K0BqNguuJKDrf
bOLOY2s3EhJO7cOqCm8Bw5xKfajgT7aY22nFFsDfTVPGMZf8++UGvpJJ+lBUNt+7
NmiASy+NnSVSXq4ncsqRBejgT1yPQSc/TCRErZNqE1tbJw+eFfASeerJS26QPzbk
SnyNkHQH6/o1hcZB12e6dCV6naM4VgJeyV4W8xbVcM+O/S/xKu+WQrAKA+P+lNg5
NIf4K1Eih22FRElNr0Y6kUs7OSRvGYWn61BhomVzlqiZNglsOkxuHgTh/ULaCXNz
YwMmg3R/UucyD5QJCeVmKL2lly0L5ZtH4dXIojFJUcGpR72mx61Vx6Rhl54pud1e
wRSmtKoiuNiFB829uVdo4ZGfsxqCwPxrATj8GGcbs7evXbFt8IGg6XAtzY3YoisN
BbbBpZVOtrt3z0R63GsYIo+a1x1reqUL9XbgpXhZUomcOVN6KNbxc841OiGf1oCs
riQVdGcTillfscvgwxGb+JfmwfpfRj33qwRWqzpkOSpC7xcp/Yl64lK+3BGp1Oou
vBLWPXlkPWPJM17WdyLpi+5NjzHhcLIbvV88XFITwWQ+7aUmje5MRaYSb2AQ8q5E
JyEO/0A2bMNuf7BVETkCUIz15LCZ98AgYyrPIFFwvsw1YlML1QB7GRZBoCSDz8v5
b1XAkZ7IZroGTTFQy0fxmV873li0gMqsketasXXj8LXpeYuOLuEcXG02ZgQ/A8NU
2Zda7rimn2hjMCa3QmLfjeuEc9sfOlF1XBJyTlG7Kj3bMYsnklqkGaG2Z7i/SmP5
SUE/LgAWVraEiGQtuTyeH3kWr1cbs0adUmMGJcNB7ZYR+03eCaL7ezSoH18hWu04
4kSdW6jREQNoj0SDX1aoSv0UMw/J9HVsQfv5la9zOTBjWXh+FSmBqdNxYumLeEJD
VwSZhL+P0UExoTnnWU/WJA+ey89XqOZx8jUAMqAFSgv3zceSQaguddys1/zPnmEL
MoDEsRGhzEEseQfkFklbzeefUy0EU0w3oOLG2a+pDIaZJus0u5EJZpq4e05nZ76O
tB9k8j0kwGMvPfWtnhkkzConiTNC1Q92/GcY3z/sVe9AAYKU2gPoOoCX5qtN4IYF
IyG7hkzzcBLHpS1NJSk061xAxlT2QdouBhYGxpgegfwIAoouGsOx5rNEFSVpzxz7
wPvQvmzpBMJVmhoS1ot8BhfiKDBs+WiHXUK4rohkceVCny2MfJMvCnDr9s8k98Lq
Unv6hKiaCyKvYdy327rP2R9xoe+QOTyMWwS6628IOExZ76Ex+H7RnOwwYZDjC6R4
y3g0CUVOf3O77Wj7rw1LoxHI8Po9Nt6CykJzEHBB0J12kJ32Xsjg702a+dzinsy2
FtZw/f/s3EyB+evt0uFmtqaxVH8+QE9bPRIhWxk/AcZOfaGxlhwPXS44TazlehuZ
aD3S/42s3qThcIzxuTzFw9LnIbXk/+LRQW5fgyPZ0kQDV02tBHlIbpRizPcQKXjD
f0q08VM6S2p2O6c9zjMQls5FbxjP1k1/2O0NaVqYiV8b+xWse21uf5gTpikxBvur
gq0Frfs1EZmjemTWcsushddk/f9fI22s9iiQGVP0Iit9md/RE+jelHMJ62MeFBIw
Ztt5IOKnsy3+jv3lWp4GAZRdq/sgwFxU1g0iluhOPybtY3FULmf0JC6VgGcuCb6w
7VF2R2HPKxUGFpFrm5VCJ4A7TERcksB14LRU7VjjiaHW7DaKUzuHSUp3oGcZoRMV
3B3uM18d0yhkVMoA04In4y67IfXX51aQpWn8g6caQRvO8TFcsCcWma/NUN/CzhZ7
s+3fk9epftQ4w/CzoHIe3iYMEz0wtZkbuQf4j2MyCKVw4f+ue4Di3hSiTFYRCT42
TIKDmyEV5uUjuMXgGEmKPnhFyRAaVqd2OjEqGq7ZLQ+CLnwtyJlF8817m4Ho+5yI
UzGlrhMqJzSrQ832PlAg9wVRWDS1alQ/IkS8ZqGCdgR6U0MKf2twpKWGPwwFzC3R
a57kUWQkm87vHTuxWZAQcI0BpYYYPLFwTyUBz4IklYA+FGysyeLwR9sGPstl+XWE
Ci8n8/pYilBKWlml2WxyPJ+YqVVstDm+NU4wtdkMTD4UjXVzECib6V3VG9BjKxQH
1LEcOV2xwQFIoBAkRfzTt7quQZX5ipklLXJXpmWQlXHvo3cLH5GBv6fgtNmLFuqM
lBkDtA2AABA1MiHIy4d/hbD+h3LaVvCpZb/EZdg7/4AjYRpqd68bnTg9zohAtsai
nonbr2QWuhfNiOfNBagvhnHUXvIvIm1RXnIjNv+w+LrY1+IzMelUpGC65pH3MNAJ
r8RSMz09dKGPcEwOWjPhMxcRF4iyUx075dRTO8lW8FusIq95ndR4TCU8Lqn+tRBY
SQ46q8Nx0eh4I/GhnjpszHVN3HStCPWm+z7mnbaPdlpgdG/whz2eiMvBxZLN+wUi
CfkguzviMRZGDWKlh2c6HP3wHbH3+cI73IkNpazgiN9ZHF5iTFyJOCiHZgkOQUsm
/0SOn1+lKogvVbQFzM8YNTlR5Ml0Tp7hsREZIxvnGJSJMZY3vq2PznO9RYFdnlOt
o2ziFsDfjgHpvB7IGmCW70plSEvxLB3s9Q+OlRkfiePYtvS9lI5XcJwfTX0xde9F
DI7hxQee0dGdjSr9rGoZDsXyi2R1TAHSc7iNLfj4MT8lSU7kx40yBNiS7fgLjZfP
kZXDyvm5XbCXwpiTfFV0dHJbHZB/6FxVuK5cCu/RY6N4md+0QvWiya0JuK6dr9iw
aUMQXn1pE2wzAfZuOFN6ooFXqT6hToD/tMmJE6G5n/gJx36odqQiM+WtR+Fpgxbz
lzofEUrnIEfuJNdansKtINrEDZgUYP2ecPqEcRbe5kfvFmdvJCtonZo4qUZ1+QyP
5Sb6ljdWdHQyrQPO0XZCDScbvs8OMyQxew5Vx8d354tV5FwRNkBKMVXoVNoBMxpU
/IQ0eJH7lfKLjWj/3XCzlNkwrF3p4t+vJl67pua1xMFoeLh4335+3dnjkJ8kCcnc
ZkehGW1mBaWz3Qqso5hx0AeHL0bynC/hgZZN9M6eMkYLEIWiyCj51ytOwEOIr9H3
FLW+y9nGyVWu8O6VJYuoS3/h3kkUj7vNhMOkP9w3+cKQKhO5+6wF7QlBYZyky+j+
bbb0z0y6CW4FNZQS7bZzEO3x5OfjtpPUi4PNWrAOxyF4GC3da/7PAQ/xcs7ITwlx
1WbV18DndVBSaYVHtHN04iPh6BAVRDBAkmQwuxzsLvmuObrm5nHPnRISv9Or2PME
zWnA/4JFsRmVy6A57FGrKe0CVUh1HMwWkIqtTj8C7+xMm8cercN7VCe+9nM7B8to
G7Iut+Jt7/A7LNCOVLXviSYZHb+ppi+z7ixUirHQsIISMR9ScGFvpGDgYUnkszl4
zYVtVQpcgBc6PrckS7oM2IXm1bI4mFeB2IH3X/ZWa7sojYC4G8rYsoNJYi4+Nhai
oWcPd4+CMVmio/Ad25cLsIi/mxKS4QgUTLwnA/M8pqJOfMhxmEJbGAGnHRqxf1jY
mTJPin2x+SeHLECg2ymVmzt4aII0orSZ9OCqIqhM9+CgU3bVWHJIyylWLMim+7Gh
J+DXYHFJQA+2SEfTYO844yATnoluyNcX57xoW8lO8JgjEjMJOdKwjx9MmHar0pBK
lvXB4MWWpJJX3iPco8Sd6uBkzk6UYGe59BCcyol1LEqsr9FbBWOTpHMnBxieggTY
bQo8BPhqOmUtXtYBmctg1+84b+qXb2SDWvSAZnuESxmZBzjljUP0MhoFCwuoYmzI
rfuOimmqLZbJoDmtnhuVsWwNrKh79ujHK0a3zlriUVrmno3QJSBaYMme1AY6ELri
WpXXvhAMaEHheuy5MCALDVuV/VTtX7WMx74di/QkiRM8bFjl+QmWf/3sfLsx+NeS
QCYcit35Og5rhXVKPMiIu1uR4JMjmuTid5aBHXMlHekxHFz9rQjryLVahUw6UiqS
ojFQVBXuHVxQWODjvK4HSvKXe2I6tezONPVLlWk5DbZekKDtV/GXIsdes9NbrBA+
q8H9luq1TJP8FUEcW3D/H9chWDk2GC5XPPx9Vunaq/9gri7t73NM0c9JFbNjq6Qy
HzAnnhtj9bPhNalApDJ6J0X4JMbXLPllyLmai2dBZqdjlJx5T+snWLrV8tpIvITv
Alcg7Xd9Ghz74VmoEOMThkDV6JTM2bFD9+MCjiLzuPcX/rTdi2Cw6RMIfdJM9M52
JBqYV0grgZNOofp9dnKSzQRg5RaQC96xx7kzsj5GSl7LDrYFUmmBaXxJEgbwV5Nh
GbwSnBtIxSYaYkBIRI7A61PjVbbPe8QVUX+tJYu8m4ycfxw+Ja/0Lhuf/eGlVcYX
kaxqRckjKUTjQOLOjk8G8lK4rdXhnp1iYdzy0ZGofHEbadUVwlFD4+H2kWI8sRmZ
3nEZPW9PrgULzq8yORFfYM8zvbBIv9DrUaq5DF4XnEYTxKKMBbtWx0owxa8Xh98a
zcSQSrt7eGt0qb2Lh4a5/0DdYqEX2h37n/I1WI5G2YN4Yaw+pDChzOU2/0iF1y7u
w3PUI3CvGHJVpPehUIDXa6cxk4DhipQGNwwqjxwXnROXXCZv112Osj4IB08R94a2
sINBwlACUtaBopKfRTMAKNXVZL6paPMPzH+oRxTwp8HuFq48ctz2eTniSJ2Xe38n
Fn12yS42F/46tEN5lbVP8tBBSRMhn14wYpqpMeLhChBgWBJ9+WlhvG1zBDw/Bvsv
OI7Mby2xSf4HmKR8xzQXeyjuHqy3JsW0xmSy3SjwaX/nldnxxUhEVLElco3tlAfz
qxO0AB11Ja4PCNMnO3Q7uqGnyFhyBS3ucmEQzmbRl6DVGM5ohjC6clck35IYgjGT
jtKJV0+Ii3yylqEhqNR1kxi2A0uf4+RYRRxw6Sfsqxss0WdMirWRorWy/mBntpfL
Qnk4ZPIZylP3HJvALcKK6oChMmgkOVjbRGiMnBlKUXpeW/GeTLwk6zVQwA+9Jvpg
y26J+C3PVKH49pzukTcUVP0Ru/2fi2RT0lrIn3Cvd1GpyaN77Ig/eFYgwp2ViEPh
WRQMD4I0zluW5QtVVNWJDvgpMu23F5pJRoy2SRfy6a7UZMC93jtsj1c1dqy5HUJq
290FYYV5t2+KslVjwCP2TGatl54x0AVBffeMIQQEoVkIEvoeqni7mNbxKAdwHTw5
g1WfCKmD9ZHjM7aTAOCloEQTGKXteQ3zVzaP0kL8ZJgYel1BdxUPKwyYjD97TPrT
oI6BUGFAZw3eZxwZViqa8Lpldm3BT9dj9P4aOCIhuZ/a2nls0ZP+fOAw767Xx0VT
bzLhhtR1zQJR6IwxrLYqH1V/YBzQ7gm8miHhKUCdwy2H3dav/aUD+BLJ7D8LFkyi
QguEpIkNfmbVqvrOwzZWM4fgW/Vlf1W8YMZUpjIQH7wwo8xD2xWXwotLWSbiUK9P
POUd/nlARY2JnWsBCdKtdZRw5SrsAHcmOCe+znUM8hFohPtc7jYI+BYz+i4zaxTt
z3ubuY1n0FU+ZSAWNtm2RfDKQ2eapW3jUDlVtZGXiEQ8eKZLKlQ8NnvZbZ54xDCG
Kb/Jgz5croHYD8PoiMQZcLEzpfMa37dM+VT0xIoU3KyON+v1vKqvU6XH/bWza37V
6j+D82Ik5eC6flAIHXw2OfUmSqawU8wbq5qYwngusBMlsd/S6H6OepRPP88El8Lt
7MO82S5iGOWdQK8CNxH3TVAqGHco3FOIZSH3O6d4CaOHmBAfiQvDjNqc7O3cep7g
sWSPfbSM5l2yZLYBnVEGcuPxbDsst0T/NHWSiF5sQQI0y9oPy0S0rUs9kCX+/ZH9
6XDiCsLfE5d4NemS6YdE8hqiZiCSBb2F0xXJGXzcsH7qtyRD/BhaCzfQKtsxFOJ0
dKZny16k1g2KJlPNeSoZ7HDpUEmdaUNHSSuixL6QSgjviM5I8IdN3384sMyw6qDE
kH+PMCJ2Qp2NZehQQVd89ZMJT5bb7CHWN9c73rNbnNtZ/rWxIfkEtdgkP4VQBDbn
avL/NlQz9lTJK77cNKv2BAwYmrusC+Y3ubm/mRSfaY3lQiAs+VTc5PLUyIfc1zkW
qCJxbnGEnMZNEyxU9JGlqD248LR0D9EBXs6LnrsC1GEbgfkVT2DwCBSx1KIThir6
TYRSaemjurpw9Cf4ghIa/xFz/UqWSS96jonYp4zBopLwxVzwkEkbxOfWIpYvNaHS
VvKXFjDOtSgJZuaqIXM/rS99jpn4BHOWQmYY534TiGUQGsPyQwJJCvXgfAzJ/I7U
GXaWd6soNKGsmud2+mIOJfsVJOxE6390L1C7d5dUtJKkCs09NRjPT4jBE0drX+1A
3xIkbt56kVBsz42P5rYuJQeDW6irNqn9g0luUlMRFCu8D6gvyHms1w5YvpQIBi9X
Abd6QRCNSUR2qRanbMIet+uDE+8KKBCXpe7lq0TJUN5a0VPKCCGsDq+Aq7qjzukm
EcTjakLWvM22mlkL20DKz+TAqwDIypyrcqP5cweZSrbE1NEh2P1BJ+CCC8seGKxC
n69p3uEpouGSjkIrfq/MK4SBd/XPcamfywUGtOMaPokdpcI6Rtas68pEnrnIwBBa
a5UfOgX8uhvjgrV1SMEjgOLTqeSP+hmvIi5ZPWhNEWxqy//Hd0wFmP7+UYq7is9b
ITT3MtLircZM1Vg76Ct39RSJpv04sV3H17rB0ZImQJiB74Ixnk+HK5CBJKtVRT6O
IFH8mozg0pb2OX3+yvWS5TCOEKf6xhYsgfAo/BjDprhCljSp7z0rSMkRhqcF6fz7
DZjOJRmVWJP4DmqSreFYWY1G23/q8tQnzgGjzyGP3PXoz+r2KggUHZClR3ZJhPlc
b7CdGIZG/XqPooDiZAQBkirhPmrHj10C0AgCx6SFaaXBhBXOjsBLFrNLNtCwUk7G
qM80oES49ApKNebKfvFiqwzTXWkNOBlmKHhYG8WuVwj52AdGmcw8DPahWFLimk2z
ZRxityeOB5CBlf4S0xUJ9VPsRMl27koT/XztuV+SE4riLI9qCFjc6UIXgBz9ZSOn
wk8I5cw5u0ZYRaWEmZC9K/qPxOrc2o3yn598YgGASBdBdWDgltM3DzrKmvy9m9YJ
oFQmDh7pOXExjsCk0jIoDp3EGYed/GL+XlH/dK453yn2owbjGkpMD0AvhPHMcq7C
EG5QKgWSPtZSAqW1nzGqJnlWOQDIxrK/jLE7/+iryNjSIFm3D2yS9tD1LMD29sk0
yjIkgBvE4cmQRYArIFd63cjGp7QEDcWxv7xyOPfPgDpOgytJslLGBngaB/xskuRD
JcDsyFqukUUAZkR7fCqnHZnb054mvPqhQdCp3sHSVnTgVqtY9YT3SjBi26i1opOt
Cf6hx3auVQwGOXRShyS4Ak0QnQkcNJaXv+tc5b/gli9mdiwmIz9fzYdfCNrbnQDV
GHzppTIn+SdrLFZfga2QctsCCrIIru6j1TvY8divaUCyd2eQHtd0TMq7tWJ96dLi
fwHbRWJQkVHYrY+mwrmP4k0iPPmDqNDdfN20DIHugbjk+gfAHwMV3WXrca18ugTO
il6KYxcxdwyd+O1T0BV7fqlNndEE8ISf7joEKXcqmq6LY7S/EGpwKsgya3+SYMrI
udIMobOIybvxbZBmIgNeArXGKJbogyiuIZ5QhrfglYU5yg3lYvBrT5F+n55jDgFQ
fXK4X7EAuBWm/1oBzY9TKUwH4YeGMxN+Lhrj2DfXzArPVBP0rZttm0PZv8dVUaqe
WWv/I2vBPbpUjG+zXinMBFxxlCe7S/DbCYI1CEC/EcQwnXZZWXWKS/saxtJUXeyn
lJGgJutT6ja29PFmfMXspiEb2Dk+voyhd9BQMGaMNcxd1PudaNtmvAMq9xphfQRk
S34jlaiQiKBdlffoG5trxMTylC5QSpEuUVyTwBlzW77JftQRu5B9f9MO0Y+pROJv
P9SRVoiltBhxgw1GAdcAXV7CLFugM8L+L3urxRWcCSP8ujG41NjCWwB0v3XJSmgm
RybMa36iqKBnwsLduaMCGMJ6P1ICzPMc1C0C+O+pUEuaoqpQW+37RDp1yJIjswoQ
vEgaNPOF2uIh2zEW6o38AfFLi+ZajuvKrlLE+pUBS4SGAg/28y3Ji4WSO8NRvOGy
fXTvZUVS0odWMm2sYuoM+GdWf+cGVhepJOLpesks7bnVQVJ1aHGQ+uB+8mQn6/kI
MKard0C8xnjlL56kQ8LXxwWfrfaaUz76lBjd4ttW72Rpo68ELu9ro65DaL5U28o1
hX3DNVqOfhPqIUSpG1J6/IridN7tkqzLnhJNG1xGQNcnr4HlI0op13DaqNoTqvxK
3Td0zVQ5OjfGCnD59Z7CUfSjb/i0nI9M8kFeKgBTBfLxPFTr5J78dMjdufCLCHU3
me5csVs0bQqDg/6ZiMaaG0YsOd57KccFUkCzBA4KpErCn+pXN52KDKs368bpbV+T
r//n8n6eJ756bgKuhzuVavr/IRN9rLKZ2vmB2eQEbRYRk5UgT+eB5KQY5/ZlkPU5
2472Sr8E51hFDsUXO8wjJhWNl4QNpapm1vA1T069RNr8wvDcDClqitbeHMxvu36L
lNQZFnjOBUtGvE+KylXvk7ByZtX4DNCNqUVp/jgI0e7PJ6CkCJ07PEd9EH1XxAOZ
FwANZOyoBAYHgp9F3NxVaq/3j2lQlVto10AY6VvhWZYhUzbdWxRke1uR8njKOlyK
jtTx7RQHtQswRnm+zQtGYq3G5DNKVc85bIie7E1K5LweGIz7NnBGW2AlKum4ABIc
1I4lXI8b5jXpbgKviwI2Fvx7UGOhLI0p69yp7FinRuaynuqtRDMB0bCTH5inYaQ5
WhXRBdpWukIOLxIx0wUICuqAJTblY+9MpmNBY46NqRnX49l5zsh5NmMSrmww1OeN
L61cPTgF2ls5+5jEc0cH2Pptsai4l6syEdCJ7ys8u96hsc1ujIOsOr3Ngk5DFWg0
XhwssEfunSzLOjyzmE1lr3CdLZWMPzeEhwrpdFcvYuzRcFEqB980vP1PX62rOgav
lPKz8kOUBxYRLXOro5iAm8dJ21cIWL3AnLS2Ij/OaR2mt5as5G/tbo8RHIV5lGu6
YdfDr+T5VVfv4BDchioZG9mf+KF5SkuXEyCZ80SaF+IuDusMkrQ00rDCUxc1iX5g
AlgaTIP0aaRkCX6ymOSkrUNnLdGLzxZ6UHDZd1R9K8Ys1Qss5Vdvd/SV1hDpp6Fd
zTaMI52SW8vZsm4Y7zOOeyCsml8TB1lPJhP6v14rXikXsFjogM3DJ/5Ogf6EgQyx
kiSdJSR+flEZP/q6+OhLeeP3HW1ATXQostL5UkwEHC0ek9i15uVedOq/nAFc0CkK
gKpBNqHDoqvPaj5a1LYomO4l8DouEZFbCna5sgPF5gOf/k0AENKAbdn+6TKgUT0u
jomJQJEip1wbrIupK8zdQ6RKRBdxEE+a7+nC5jIq5rpDkUqYFn+3RjqvW0b7JBWe
C+izDeIHlzNgVe1svhgKP8vHX9sX4MNU1N2t3tuNk+lJZqqoh+B45a09Wm6ESr31
cY5qqoefc4QHbdaaPJWmkBfZVyHhEEAsNuoAatJU0KCEOR1yW7Lhl59fTeL53msR
9bw01GHI8kjIMa2h9JqpYkJw8fCdJ3oxpu+as+dSfxaVDvBExBFM098caOhkMRiF
jS7FAwhFqceAAkeOdVGIJCsww8fXVPbLsaPmHCSlasNHj9ovlqh0I/JSLmuS2Krw
Jn8ctCMqhHtfcNvFJoNDeqgqw6J89WkPR5cO52WmsrxpOvMzXFDL0xcr3ZmCScNk
I3fa5hv2ri+AK9q2PXGfkycFHHhbXQVh8nLcrsntCoeV0BNexErs4iPr2GnpdrDt
8vMLYxVkp3nd+kNVIyyrzXjv7gpWCyjtPW+iozJPwrBwhveX1jiF2bPOLc3Jg+++
trVyMA/4Kdqa76FIGA2zzxxaOSMJnEyisc5/HsKzj0tNrBidHzFiy8/sadH/fWGm
RIbKzelI4O94ms62Ooneq3SUTVXHwA7Ex0/uk+KwH8z3AZg/RHtBgGTaX9tbUlmj
mneFgPRiMgedurnj38JE0XtZskM5Rqs9NByzJeA047ICWz6+JEVzfksGG0k9MTB7
h+5PCPugDFfwEfvO/+7h85TZlgM6ephqoo98ltBFycmzArdJOhrXC/8rZm77Kj98
G9kMO1PKfnrz+dSkE9Ju1gDcPe7GeBGy8ils4bUf3Qw7ZsAvUmZKHHbTF97N6uv5
kZmCV8X3Yn/piLot+8xtcywcNQUFrbhzVnwmJmXT8s0ubagqmS+rvh5+Ou+UlYIw
LRJwBGrTwjTCaoKitsQsldxa+K0tLNZH+Z8LCD7f9rdc9feMgCb9ekHFCYjT9PFn
UN4xAtu591eunu6LtwzrOkA3rJ3tsBObsZ9sVe4aADRLdggsl0O8tpkNqZ7/BnqH
5vIR3iegY1S8uITaTQibXl+hznjpsNu9MV1PMzRqYXLkKdl9yyzUNqbqq/vvyZHB
JEfNPEIBrUuzptT+0R6GBL3ILW1XgfoT20XPz4CNiqEwDJx3ZhVEpADkMo4YKEjh
9f9fbIgQM8tKmYR9ytdM6XKfk+ueT8zroweFvs95RwWaLIzJ3daKWAE8b5JVIaqx
alhIsC2Y11ZeIEm3xIBoyKOekQGZWNye1kPKpr2jMgG4mE/EbrSPn/cTmCDbWDqm
k6i+GBJ3Mas96vgTHc/U3RsGkO0sk37hfTrfLxPkdWKv/fylwAp/jp7XFRYu4aKa
OlKxlV2oqytRbB12Dd98e2AaLFJ4HLS3Paw3oUvv2QntUjXy2pMgLy3+FQEOFQOl
lk7eqSkUWtGhckwWnXPufJW1dUoKzm1c6X3fTug3pqIisBcuqIglblhBmE3vcVAT
2bGmsp8J9UT+MKEiOroQFGfJd/cmO40l9uD1PDPafGqbfwsksJEXQ5X7bh5H+LbY
FT7C+ERvj52iBODKitg7ggdIHC54SZz3VK5Ki4yhJ5GUsG4IJmsVCFjhZIEA/Z/i
4lQ0defTPxpAlfWNotpRagnfvaOOzaK6Dm3JduP9uLfhqCTSq673JId2ST4YJe7a
38vMJjhB1UhXksQr3kJ43tTk+JKQxqvsH1T2yMI8H3CJh/f9U8zG6UczKqsxHvAJ
edOSSZjD+V4TX9qDbVDXba9uLtpNLRShQSiMKbDSi1S9wTicWunrDRKq2Z5vYoGV
u7bXyT76lEVWXyKGHBSXBsETc7VvM5MipPcufdyX4NLIKw+rkvARtAsXPEyQBRbl
ui76+8WTiL3Mkw9IbfHE2Z3Q0Xior7Cz0Q0Q+zpfZGtEst4xPuQ6jGU97DGss8Y6
dKL49o3YIzxbEYNbksVDzFYhE8AJzY0+4MeJBD5M9J+R0SBWa4pj1YxqoJ2fsrDm
A9n6vSc9QPUxNcj/aNKZoA3hch6/7tWB76+T8K3tzwoEWImvWhZ09SHnfWDDO4mX
ssTClQRGaBgIeHGCdO8z6dxDz0vdzLhYpxi1hr6WwJZAU1gov7E4LP7sTYf3dFuG
mLo7Zy28sm6sxV19zTEEGmCnnvTa02isDluEmCINvQbcWRWt7aKzxKO7X5XYxu7u
fDOsleWKUz6kn55PL/N8LyofjK3PLPOVK/zK1mIirOOZttZpso1tSmdt/xSukJBJ
eTEHhIS3AJbfGBfJuAKY5KN5A/vXQIwOBZabJHwGrdxzvY/AIHHbUy7mYa8mgt4E
a/mELNZUMD1GbFHQpEJW5VB35IG/D6mVpyOZKPj5d8iWxFRqcSeFsdjL+psSaK4V
6V1qeA/kGay0bHVSl9hDFI/zXGoqYea61pTSldJEehrnh44Hn+MlGjWbF57oAQg1
sPoYUC161qlqTBMowJjKZULfm1LPeyegnIz/Ad48p6RxaR9D4H2yXG3jgemK/NZM
21Cc6X9JOvFEnH/CtgpY5/OMlRN+BMqw8bX4McPNWu4ochsWYxznaVzsl1kj1n/D
atAe6TF+oxVfX04VjWoQmtBkBTXlMQ7+ooj6AUNoJfrcUASSJUOa87nehvAeY0D3
wZlyDp8MJwrmxhb+ogLKAb6skeu/yFcMfs/m2+O0XIVnFBeCkD9y0abk794d1kKS
Ml1GAW9NUvJbvYLcI2jfNn5WiuMpUTPrUsLnlM3q6b8MJtK62H3Cw75ahMnoz4VZ
RmYY2Ndxui9NnoF24nS2LCvvAor2Edw32XYOMjQzH7QwqwP/lp8ALynuYga+pvzs
LKDbG5iMknmcyHnultJlKoHiMxi8pFJgThZsr8LxPwLyzdrZ1cida7yY/SKOnDp4
TKFu6gH6z4+tMU9UA7AUcK/R1rqznDwyFFvbZ012Ut+FsaZooVCieRKAWPK9NXZN
6gUz+i9k9zl4GqoV98T4FFRekiYddga/FMrF6TPSLFKD0vU030ag5+UB12PoX34w
gwqySvXVUyte54eQjLtkfJ/Ut84d3UICWF1SmLEQWurppv0GOG6HdSqO53ZetKTw
BJ9IN1CWi5dwgPFCu2pAfEIlh0XH46F6ZW3Mai6gV3TBapQUpLHSeb7feIWbwVjg
oFs+5jqChu60w3DSktq7ymkR1XKHFcJMGlsjZqPQXuiqqc0qS1i4LWxsVwO1zOkD
VaosunTAxGdyHTUS2YeoEx/D56hhoEhD3cqSvALsNQv2q+yr/YEe4WAzSwfQ+QQN
YIbsFmAuT4EF58iJrwoS2m0dOkzJISqiIMvmKZaUxUPBx8gB5lqvur0bW36J0wNu
KYG8mzv/OwI7S5hScCqG1YBQ1jYu8tYqb2ly/zid9hERFfbsJyizJOy1+eGdsfx2
IiNoYAhRk86ppOvAdXcXqpqTOpFxZ7L4dTyuwnI42BpAyF0ua8BvUeF2wLlVI7Wg
e1T6ko8w0Koi3Wf6wBE7VhmS9kMGncGfFwzwTVAkOZShrBkqioNacvZ4BvUFCqvX
4AcrlqKzk7azKw721c5AY9DRRm+/aB4k8ahEZA+5tipKt3x85lzIzQZQ8p0WSDz1
wn9LEEgu5ejvhMpeOqMk7EHudd/9JIM1pcSC+YgIuH3aB3yaOontw01d7BQpS6BA
K+R3lfAK1IMOJIOcEW5ByIvtPYCsfZ+FwwrpTqwKyz4KaMEfOWugQ7Vve5jwETEF
nzhV1GMbNGaRnKUwpVK30Nb97zgghZPJxQACu/5/bg5Xo95tfpGnDdoqnrsajKz/
27bGyH1PNYDAp1SqK2lE5uUzTR/Wfq/7su+o+CW6Nbu9oW+AoL4obqTN72JPOA4O
cecewnNclXClQl2ZvDwn17LPoAwypoWWmQ313n8B8yk9jdxFAXUSuNQ8E5oOZvGg
GWXP/m9nWoZ6w5ecz0/+9upmEzKUhRE1P7x3R5Jiq/jNeJMyKCmmhpLnj3dIDpuL
e0OkhbjHbtuZsnu2FBSD/7XNol0mpVkOmeQjjVEnqSmydcbUX9B/8qqNt0uWV196
tmb1Cu5uHY4MQOXNejWjVVTRQkJnWx9kKDNFsiiMhLVDWOqpXdsuE4YfMofPGoiB
zcwlS6hvU34ZZnT0zamwFSZyb4eYaVbxR1kWlEOLjPj6Sg0nHm6NEhW81GChktqv
sqL8g1g+eB/OdoywznSpD4fi+RT9E38j2s2xf7RfJp9edMd3LZmjXjYFExI6fsrl
vr2W3ENDxVrY18Z8ChnAiyaMehm2BqlaxIi51HL1fNnfgJXW0ARPammuQrGeAm26
sFtwtw/SMKFjATkbx5JhbqDsL08Wiryk9kyQQyiaMrsKyaLL7DQ3z3TxKn2+2mU1
1O6Cr6lNg20b/oaze2f4bms7PkXvSaaL4H/Gh5e497GW7M8KLYNdA8KfSNqcZcHQ
QIC4o1/Ub1jBGmDwx4AXzbhksh5htyQZH5pNO07uGW79BWR/UAlJD3l7at2QWHVS
LsRsDMT98/xmkswQk2D11VZUxNQG3ecCoHRpybDoYPNVaSU6mpXQDTSaIaXjfpxL
8ZDziXNaDv7fX9SmaEzlIoQq/DSNJx2DQo+6I+4WWCzLnLOWRvblZ9xNAjd+5Z7k
M7Ff3KbltloeO2W1+Ye4w8buUX6EKJuL9sUVlHgP74lJIFnbtRfz1pYaB/90QvjZ
/+q7aPAW5tKkxzTHwp19DKxX72v/CfOrffMX8ep/DXZbjotZ3zoTbj31gU/xsT8B
oWcZ4p3txygonMVnC+IEngbxoZo09yDR7jXPl4fXIGpGSZr0xvw/T1G4xkemyNPR
4zQc3a/ebUl2QPoOAjdZfAHfPitW8JBJISYzM2FLLDThJL04oUOw4ePNixs7RBRb
30nwvKTkosBMTpl0Pdur2g70G3I00LqiiESxwDkgAZwS9nCBc+hB8T31yb/Vt25/
jcXv1Py44rwHX2lmXVgR0mHJvlo3uJGEON51VDe49asRfx+GaI7ONmhM3BcFgnSN
N7r8ALAMIccKD9qUmjw3VZSFbsE752a1m4PhykGw4y/Ym1yRmzvIrUdHIciBZZPz
AMYe9c9mv+N5YUn1QtX/owOQjHZ8HO6c9wjaIDRCNopv3cEGqD1AblBSkKl0cHne
trZZp5e0JlK/2hJH3XOEtG2gnSblDDSTGGgle+i7GmspAt1QddPeDuPNY4bhYBI+
cuY0h5I9xt53rVMu0btxEb2z4HH6Tq1/WOD4tVYHco3TVXe2XqJ0868w03mG6mDy
44FMikU3sUMVp+OwzD02fyKcc7ci9DN4N4/vq4sKhyO9rVlAOOveAF9LzH1pi8AF
u6LkriXI3K145LueBxr2V5udT/K7KUgxcfXeN0vH3twTstuMwOJphyogTQlus1aK
FKrnGTVo1XmS+xIgeUcETOUHwXcwL7mQULb0QRXA4Apw6iD89QcFpbI0YmOv9PhL
t8SjpDcjLtubqJdsClo813wN0FLmLbiBLbN02uUCL/wzvytKFHuJdotVhf/WagVF
aiFKTBeP6gOrdIIsl39t4Tzx+LG8wTMNybeEw331njZ+BgO/omuoBXEvvAEZ/ivf
Q+REdKHUEFkHXx1lT2E82JMJ3ktuwr1Rl1Gd0nCbd9zMxA4zwek9KKc6BJkCqcKz
zNmJDs5GW20wXtINdqnFhs3Bdeooo2mjNiDVOF/2dU079fvOdqbzmsPO1EfCwKB9
GNMHeom23q296cbsyAOPZ8dP1D0/80EN2N/VwC/KYM62KnR3px2liHsT6lsp+PEp
PyEeRM8rJWqorDB0319TaoE3HgB64TrRzQT4Qy0ZF/Cm2NKJdtWpMZU15PSieJSI
2w6Uw04mKowPQFTb9Yvs7lImaZ78W9uk7UuV7ACM74AEtt5miIKmRxEQCRkCi7qN
nCEP7d+sxO9XkPjY/oulRDwvqKt0Juq1kyqSe+LEeN21FGc6W1wTnQAtS6uX7YO0
uk8MADkJC5o8RHzyTpNl3V05s3eOzDnZM5HIMO33mfd6SgmI/HfeCD3Tfchn0khG
WR0CH3I/4AaSPPE1Cz5rEXkfnIAoq/gwfZRM8EABGwkMpUzhiqm+RGNAwvzr8Vas
3s0cKeR6Dg/l5NnrKkKuG45HWhtgOpMxTjTbqzf90XObbn5ss/LFqzF5w50Or65x
/X2SoX7zkIepPSobKaqO5xHu2qjonVEh21a3D0dts2oV4LLPRgppQelpBieELknz
ST/ov27XF2M4/p3h9qCbWCEYjm4U/T6DhQERjAcQ90zRr38oxH/2FwKBUWRa+ZaX
Zvep3ctQdDiLIZiXIZtMh4dJ7OwKF1A5Cygu5VFtsGHYa47bgxgAR71FSl5+S2sI
7UKtsUe1tcaXNHlF0VG5uGVFf9TqobTjncwWqOfTmWseoOaFSmp8LiMi04DPEBEl
zV/SD3rYRj5ps+9mnfqHdsgPbicyqkdPzx4ccxOaw7EaDOWrGfQ++DySPdJ9wmZK
MBWEs7m1Nd6J0KANLECQmDm7da9REYc8WU7qft7ePnA9Oz0U8DH/nUByEXbtG0pl
og7NcGUr+HAPFmbPXeRogRh/plyjft62RhsU4IKnVo6xYbp65SfLXm6zxixl/t3d
jaKJQhg6huSSBs5QpNA18FfN9R3C5tXnzpRiHd9QmpwIMf+WeUHLFRRCwmGY+pH7
1bu1BStmmZGXUXgxCbHruB8ZKxWI9XvqgYiT8nx5+grIqV9ln84gnNtM+Y2nzz0k
p5Gkx86I6Enpgm+5HrsrAF/lwB00Goa7j5iFNR2BEEmU7Lfygqxh6yavOBJHi1br
I+BpcxYe63GD3YyiRf6pEsLhwKHTw0n5Xh0H+ovpteovgQCvEOYNUm9cQV6HrDRD
Ba30I02iulJCWCwJnlLH/AmjOArt9Mg9AkTABFIv9xOevyalPy1w1GpaQXdqsYmJ
jvdfGZBN3/qZZsWj9tgFYnN/5bW2LqMxd0dMJA4igft48egWiZxyS9lJbaClPUrI
MIIhaY6VAxkxiBapUzjNfjQwwhHgYD6wfN3f6wPE/fD7cdst0F2lzSbaART0j8ZA
t2878VE5MWggEKBpNbtMH4K0yIxVw3hxtMQ12/7+Lbgoz2sjMZf5G+rCtw9rv6m5
8Qn0kzb2/tOEdPYNH35jZJNyAnoWuG59ft5aXEnsgQn72Pqo/6H+yG283hAIm3qX
FEOnyXkrtHR7DnoIcV31gZmupabHjr216s48BPo61T8TtoCT/kFiN5l/kxOkqHjH
klf0SBCZdZ505iVud2mFX7z7HXn0tTt+oReWSI0kAtncnZHuN8A8zrEPURTztgx6
T8k33TXfJ962r9O8ZyW2PKPJtlQFGysHZyIOd3a5CUHydeISrxE6Ub4enaB7/5lF
PoV89M34fOdwQRET1qhhb8BNJdEPBmJ+EBfCyF4WgR0qc+4V/JJqCgeiJI5uGbFm
k4nCkr7iIFMtRDSBap1bTOm7mO4CdwWDaFnrRQrRZnmRsCFBu2tZMJLF5Tku/jSy
Yx6NlKUobONz/pc3kOqC8BmDQI7WfpPyxx3oAK9NBW4IygCMQjBOu/OTUybc8qrw
Vn1epls8xq6VYwMbm7v/8HZp8F4NjMouEtvJcDT3fEUAGa7xseoX8nSo5HmQHCGi
UJqB7p7N5jJAJVFHXV6/6HGyRRr6Ikbw46zryn0ocJyWe4121UT8Voe8W0y4JjQh
j1i6WoUIaBfrTNF8gNKer0iOEWuVrUuVraVoTIk7PVyuSRuMwZm5HrvvXte+52s+
+Sq342/2GnIp7GqGvsmx11jY1VzyEtg2ug7cf4ki66MZYP1thAEr+CY0WlPVAkZH
9y7Pququc0HA8CNcHB64OAngj2eeScJfFyEARozjedizgkDsO3kN97LFCOBHMSm9
yCWHiXwkVCvGU7SLHRHRSV38ZdG75xRsCgDqpjolAuxgm2b5n1NKKjWaBvl5VQvI
JGkGvNLU7XQhe+DHWBRMlteL7RLvW2j6LNi+/1WxAUwxsVyGFrBlsWv5MYXkVMhm
0WIOHvPcVGoeAB5gdc0qbm+3ZEsbi0uy54NXJSMmK88tDf66q+ofa0GxGYE27W55
owOlSaCWjpAkKm3nf9a7B3l+7HK1FLJErC8JWtMSkoaLRgAJpH4dhP3FTxn3TR3Q
bYC+sKycVT0Znwjrxohy7nUso8W/iF2cVxwkNwTAFKHTQTgA62YI7X3dYbv9uERE
uZ7NAdMNUJMLngv+BkLavj8gvyyOxeaQ60JDKnz8TatCIEIS1lmfXX5WR6YDwab+
i86Ut3qDeUxcf02F9eHCcWDzHKS6Uy+OB/m3rI2+I5L6XrvyHlTlC5xtPfN4HkRz
kBJGoDHkIdK3+Ostp8ieWIyanqp88a+SnOlj7ojHTveYtraRDRoIQLDtDKMUuxbf
iBNUuD0oePW/B/BO85GKVm3U1Ks4i4a20mgoXCKiYCANH6bVfSrAXdV3RT05+alM
iDWc3QM3VTnZT4smdmf02X1M5/fV0ZhoWqNtKjJUMbywCNHeNz1pSLwIQZxMr9ZY
7vR9o6/Wmyf7U+taeEeYNeE08KF7Y223EokmNx8e7LXGamj2bjT+Jeo7L6BJ94+L
Ii8I6Hzk6SDdMb1P85VJix9AYduo97xCOCtfTHtFHLYoGPlCqxK3Wjg1z2YFQzyc
x0rgM8UPnLNjGMOvwBby03+X36fEVM3SyiGgsBpL1T2+nzwnxzA7mX7HaIiOTf5o
LIfc3C9kwuZSFhG3NqiLTaCfb6hHXP8S5xWMGxwn4aB7TMRsKPbrOg6W26unjBDM
OUfGBl//9Mfe8kgOUdbuMFMghxmnJcXSvrrFlCGghKUW16Rh6V08d2ba7fHlAKMt
Q6tMtWyylqaLrc0wIWDUmcx/qDTRK5S4VSazbjoGSokaxi1fubRprHh8KpqTnpww
KqClRe6eJDXE/NI2HZYS1Eb8ReByeIQwB4Yl3PZAdsipiwTKRA+QTsgGwVSok+gl
FUjfug0EhUYgYRQXD80Kd6/0FRX4SKD0qHIf7GJyub8rAkwDFsyONqjG3ZqZdHeI
0wmdYNW+b8wK/e3qXeeG1jF0XthLRu1YuXOYKuiDDwbfabtybfZMl+EXIywGdgay
Omn+rVrQWgBKJMgY1oFSuhmDAS373tVd2JQXoH9tVQNVQeoSwsOJyl45wAI82joC
GrGeh8tU/qOCqzCRVGZ7Zy0Zpoxi6xFRCAZ6An1vcz9Jvkmx+EUVywQTkCaG2cAZ
4yMhofEWalApUwv3szxyiusSKLEBbWYpEb/d+fCKtzf9Zl7wir0f1P/Nuo8odQWG
0agI1UKmTiwkYvDcakWRv8F8UYHPdG8Q7LbnC5DvbJep5w+cJrbUslfOmjbF8jdR
EOPwtI6bKlduNwmXVlZjvD+FQO+9bd7dNpmZ5rknAvQnS8kmH0w9wrl1G9DBiRWv
02sqdH25j49/UT/TXVyXIpUCrif+C6Xj2Evno2izhM3uXlBpX9APMR5bdCWLLRNm
QGdHL3oQ5KIZZ0PwCQBvdXrIsvfsRx7QNzUJGy6VX2Hy09HYtVLyzT/Ib3QpSvpP
8bC6dr0rOOvFbw3rydjVdSLiJi1yt33xDRjP59/k3SSFfINfB23sPupAMhxtmAsf
ZPfBY4huEgWgW5kO2/JIMrfyO+jKyThWVVvFAPfWhXUJOCxfa7Jt7fkmm11LnXcZ
cXx0nX3PSrW48GcuazYde1xiOMkW9ICgyLvps1yn7nsEEtUbSe6SLTZfnmj8h6TA
kolSadsWKbio7XjA7N0NGAoynLm46mNy37eeqM3yE4sp4jHuhZqvgsGeLOOVmOPX
3Fv4bN+OqzLh9GRD5MJe2Fm5I9LWPH4njPSItdvYVroOEIyzhI3Lq8ZI/Q0i+LsK
FkFL4uLcwpB/0m7ovGQdmEgarJrBsO5rS1zTqS4xrByfUCSPgZnSEu8PrWAFNVzE
JHN/HdO3GCfrixGDCrNcqtdK8WnW3EIXUAhc8I1y9/1x8k84rz4gIq0MAqZQgWft
UQBrPHlEqRbGbHMvVbI8vIoqMgk35vMtiFjFWDlGZ4raqj3P/WQ+b4X8gTAzmyF5
AXIMq6WQ5WkTHo7FVfPzSz5u0pRiFqv7moLyNXQuLjfZ+DlByES78FJel9CWJsaL
EFTUGwQ8C2gIr6UAyypntCycF+0U3xRuS1FOz79WQPJwzON73+U1F88WOQKzWztk
MVS5bFdZoV2K48BWiZEhhp0Yl5JbgKObq9WksE2um/xhZ3ZpLYaE3MQAO9onZBBd
nk/Nf+5XSoAiTd2hP0WIGKhyV7CDKwK5Bu9G2h2XoesXgrjlJmxgKPoZrmGTdSIc
MubmonwLokD3h/HdMyqGMh7MCbe1JiA6erEnOL248PHffHQPxDu8zFKa7fLN2YV+
qYg8l0rBU1ciawLQHNpX6kNcYwghruF+R9UZ+YoamqUrMsONHWyRANv63v1+FJVP
9TdMwOz8btD7Pmcg1d8s2sLkVPSezJIAldI+FGZOBXkisFYxujsmM+rXONmmPC7b
K07UXfrkUYzrS6n+1utke/RwOc+bYXDe8LkZjumZAdYTy/VcgAfDPXANvVI4lnQu
EKHyjI2DyXZdhZQQqtmRUR3gRho6Nmrz7S5ZOK1r6DRvHrlXyWbMzbbIJYH0nlzu
ghSQ9GlmvGczjsb7po3ngGmIv/Y9h96LHde+VupgUJGwfRu5sb3MR8qcjBoaww6n
EwBN8EU8YqmSf1VvuT/A3siqLvrwBIEa+39CQd8DuJuh5gF21PqYYSHY+KTlMlcp
orZlXIGdx4LECTOexFUXwqUH7m+wHwSuOgWxs3BqFaxvmE4RbM3j9toz+/jq+Vak
/NKcGSybNa3uA2qsxGcJY31L5ukSUxUWi7iYLhCKyoPHafPx1aucJ2beKMCEwGSG
waMgD8H6B20GYR48+rjLbRAdUkNpF1M+HdrSWFXV8UBlmIlHVVA+IAxEC5J76juY
Oi0YYLVlmZMTOYPBK7RXPdKsmupbdGv+oEZmVOnQxyYSERj75o0hg5bL3yFMDHJ4
QF/WhgkZPcd/h/s/3FWw61VtC3eqnQsuB6+c90xZDfsEylyFYDGbachV2vYcv1hR
3eo+SvYbuRHtBkfROMudr6fIp8InVelg/+gsZ9w6QY9ZMkuJTB2d5tSIiuF70YKv
ez5E9gIxgo0TUqSZVzYE3D4uhPNYL66hWPuJICpJ+cw4S/7jjzDzI7VnEkxf2R6i
v6peJwXTiNc1ufNjQL44MFV/sXDUXoVfTSoPurQ9XlKcFZ8lJJHUIfC8+f0hih/N
JhZQ479dG42Y14/c8ZPfGJihZ/Ri5eX3IiDq/uxxMFNFJXSNjqnl0/sXZKx9I/D3
8KKD98DRNkjjf+hRfYZNfTYJdg4OBHVCBST3Qu+tttyYbtN721T4EvnXrBol7VOq
GHsQI1K7/WtKvgd2SJtaATbzQbfq82LFSJTGBTferuVhbVCtlM6zFdRwlj8V7gIq
d5L0G8y5dW7Y87lMtkL4yLjRa2Ocjl87nxQBinAdbSPfNAAFD5OPS97dcLe4I5ox
ImmujSP10AhTw+YuBaxRdHdG6TIn3h4hA7v5mtaXTW2MpOnvIvAxPdw0lIpBAMBY
29zr7OVuKwhLq39ck4VZ6tFcY4/ipm9/TJ2WlymeTujEZqO74c+FDMT6o7cjjZsN
YKU9Gs6/lsB733QLlRcNLBsfCvjoh33UlIsiqdusVNzaMPEd2kzUsD6hZWnR2T+O
dTPpplohE4uvmcHF58a2TMZhfJMZpv6CM+7o3hMbAKdKC+vCo4uaSWCFIoPPyao6
teSNELbXYumvBJLoehGKuZChdVKXk16yRFoZbKxpYJREzY3Mo8aKH3AzuqQSYikf
l/dq41I3vVuD0+LbgKDUewAHVmRUaFuJVVtlcMctoWMHS3YNyEruIH/imskDyceJ
AnsLvsHUau16wmTDzX4QKsgDFyDUC1c1OGYUoxk4GhSsCTUfuzOIHqUdRgElTg/A
iXF9dw/hXjMMYimL8At9NqBhOLdbXepViphiuIB0F3yTqDBl9sbj6MsYK936+4Lo
YKk1jeL5Uo8/I3uw5rgrEflPHPhaaqCoYaa3PmWXWWV8aH7cDZZ1Q7b8FXr4InGc
vmIU/5TWJRD8+T++PGVOFzcezDI/NNJgklhRtqwoEsJvvYmg9uUdvm0DyDUFr8MG
oXRqmV5mZsXZHHubAxSb73cH5CPpURYjiVwJnH44TjbjpuBo2rVmO57DWPnkEQit
p1moF9NT7DtpTZTlWVl9RuNTiuIX/QMndEQxY46z2hFSwEcTdTf1hxoHTevYkE4R
ODI6om8OmapsYzxuCB99i/aBaJ47lYb18GKBbWblek8HjKiLNx8Bytbs+kQm8Y8F
DfWmUPnq/DPRaCiaTVvapwjaiYg6Hky2U/fe+ewYBjT0n6sYSVkho/UHgn7+u0qL
oe6ad9IiQyTuGw/9OxMxGC54xzdyqc6VxHggO/yQ2DDNvimlzh0f+QHuZdtGy1IM
yThv+KyKXhvq+iELxgwJHvnidbyGKi+iN/pxTKm/FJbMSmOq7S6GvjHj1Xwb8dSm
+ayHs7E1zbI2Xuv6AOhQ408tNY4bCMCiKFazbUeTKGq28ZQaUO29EeXTchN0+3zE
yCvUXeCk/x/FQE3exlNvNO40iRolAxu8rXfBHMaRjle1Q3A4YRDf6h+Hsw+tiMhY
PeVz8C4rOHM0pHjRfS3hBhz99qPvFNfeN4UYgcHokcQ5x1AP6xUDBrVMY+elgt0L
zq18rfdd/QzFpFbXAXdZl6nOLPoYXDXEbOsge6OkHSdqszCRc5m6yZ967ldN3UEK
1Ky6TFHT15PYZms3VcdINKs9mwNhpikEsBu2ZV/MljeZSp3S38w/24U40BVO8p+f
x1pC/j6+enb1GoDWkz1omn+uZh0KRLzRRkG5iie/rmkZnp5C/oigYZh+RdzdFFvr
B0Kfi+GDXQ+oELUHconCsqtiuDhXYby2C1z851jNkGJWebzSrGco0pVw7fV6DUZ3
vpoKLjaCAVgp6vcpHN3iGa52If5exfO+08NBTkFi4lYUGrwhsLze3AbDnWyTE33u
BOtj/IXUrCq8iITaTWvzg896Mhhpn7uC0gyxdvn6V6Bv5KQ5H8kAVyU2O01uITXK
gaKc6iU1W70FXQKJ1wQt4rqvwNeTIwmjXarcUpixOGLPX5NGP2ji9ClXONxxLTLT
BhnRC7+KCfdAuAFNjGrJmWi4C4ouODK8R8WA4OTStvirO2HdNOflo7u0KgnpfUWT
zNgzPU+ng5+f8Z1bE2EsAgdwfIyKpsGnFFQXOM/bA3bZQx8kJRrt6oxk4Nvl0QBH
M8TbWAcyWlfq2wT8q9p0oI+hY2gzVvy+zS3AZl66FrvpYLkzJG+WtAOgoWak39Da
Vi3u4qQ6G5mZSRYP21kO4vjEZbt8wfPgHFflXoBlbepR/wEWfreBZ5LPkIz4oGHm
H/44FqJlIZp2mhgGoIhOGn5ID4hAJJ22KDrbIc7qaLsfrsk2Mxdo/dnA2bUEE1l9
94KCDZyc8Cg3Sdlm0FB2WdwmBHSIvVxS7uMtqbRjbAtQiUjfBCaxYTcnSESipFkP
7y0hajx3Chlg0p9WevlcTpFNFguI5RVH63nI9gta9M1IxKEu8+xwgehCQA2N9vBs
X0EFMx9ZYHAVJozgSM/WB9LK0aM6/VsDbg3Z5/f4seAxNNEVNES7EXklXtCOH2cG
a1CnF9VReY9J07JsyAtMoOovky+0wwfNH45FlAeLIynrflR1ROK88BfIkWdYELwT
FUatRcKim86J8L4Agz2vmTlIVzzrYgpClW+b1Pcd4kYAjx4MmlzBLhkM/XFwsorM
IMaPpSjbDs5JaFDXZHCf13E1sjeRzbs1R+5a01/CCX/kMyJRx8Dg3ggBz7MGmgyu
DXCcAsNZCyX5Sw31KseaPNAebZb/kwGyIsfKKBZqhhdFBxRC7iVd09eOe4Ele1nK
QQvDyRccPcImj6E9OxgRhyfHaXYaV/Bd8dirfQ/FPxW0Bvk1nrPAmIwn5LAdQ5JU
sWwGQaj9mNQQ5/iIFfqj/Abn9+W0GbCjzn88ktVUMXEmb4DKbRL9aRN7g2z7eTkJ
qWbB/ln7SSvLCCbAAk9UfkwQkiYyKTO9ViqUM/Y0SzC56jL0c5ZDq59LcjnNBlUc
6caIoOChLjq711/ZhaelfxgUSjOaxUUkA3uv2oYFw2h/Gc22fc6of550xQHJ1PMx
SWc3AM+C7r3JDXwLpRQT0DClvOqg5kZWqjgT4HpMCUwoI3bLM+HyJyLrY5TbFOCj
XI/P9gwtYgQ3DqQb+r/dCEbR+RTTl9TC3CuCg/VUZFW+XnSJJ+82rTJ97WneGcTX
ZKR524DRsfpoQUNmUvDO1FmNye5Rp6qkxLQx5QixghxD4TACuM/AfvdDlkhN7pmj
hIcGvXHB+LGKdzZXLTUSDRQWR59VGwY4Ot8O2tqWokANJEQz0bjM+vOHNR8l4j8e
tgI0LrtkgSMntPhSk40M51BSz4tNAfWVQ2b++JeN58RNr1njWGLu2omZXIBQLwnl
aQFh3z7Cnz+XTJyZsyQAOsEy4ymlCx55qBgF1U7L1ob1vAbUeOcqmwOJkMap1gvx
d7krufLDCe8bflUCL6RKJWyAGyymA1tnPim8bbPDMrL5lqWwu14IvccgTnInHRz9
gTdscGrffaKaJwpDt+M150d+vm6bysSQps7S7rRBzIDpqgcudV78f9QgA7b1Y7E3
AlKOwGRNDGY9hHg0H4yHgum0fJ+7Vzld/7vEQMTs5ufjzZ5otiS3tPlydFDYKAtJ
frpB4FN/ge9Xy1bz3ss11nFOYTUJ8RCLgb12v/kx6jlBKPm+7abnqsEZoPaKR9/1
ovMWIyIlioaRnKZMOsOeHwc1nI9q51kzA25skQDYcc5I2PGU+UI9xH54nsmxpdJC
0+J2ns+y9oqbVzcmDd/zW3j3o0z9k6bzqezkdY28L1yWAKd2Ny71+CHzkRaEeM3X
gFXJ5wmwdpqYEHxlhloQ0Je4tSGtKxq2NULpzpN4rbkWT+IpiqwIW8zd7HrCGv7v
aePE3vXoDY/6M5izddBFv2dNNEdKAiIKhlcI0Kwq+qv6jNM8XrjwjrWKq1GS6JPB
7Rv7wC/DdCKE/DHKYcmTnp5jNqWmYfG/uPlmI+jYGPbCAvzPF0hyK1s4BceYSltT
nWPiNhbrSPgXbKKK3T1aS0OZobGK9Mb21BEQUL7Qksrb7TyW8+Vh5mvx/exJnD9e
8D8VuCOYzr7zJmP6224+NIGg+vKaoiRxo4zNvKSczQqGwQfRMCE52AtgLBMTC4Q5
ylWYlg43OKg+UUs+JzXtB8diT4L0mxtdOnd42b955nzDeRzGs/qVL/A14x3QjFCT
kwL295giAPQAMYiIgG/fHk9yya30o5vvxLu9CjiMV7jvck/GiBizYqVvw/5P5Rph
cbN8r7dKJDyn5LzjfbIA4vWG9jdyQbMKkhOPxiNa9vD2fBF8d4M3UnAEZsvtPHI5
3Z12kF7D9T3oFVXWENAJaI0SHmS2sTL92m/D+HFU9ME7VIoLrySWw5/PqdK6qL+D
wrOB8BPHJLIjl/atLa9K29xjpmG1XxFayFh3eU3xKUQY1EhaWJgSk8A308zPNo0t
vh8ndR8RDCb5ZpneZN4jh2iiISK4rUvoQjVvlQYB6PBRrptb2jde0u16gwHSiaN3
Oh2Wc63iK3/BKCp+2c1E4YksrE2T1dV5o26E6nIZDPa7mW14q6UTppWMYWg+Wv6K
ON/2vkKkhZvJN1V066me/w3ZRCRrk5AIC7s5KNH2+Vm5+U1LmRlWge0aqyISux6R
DRm+f4nde2DODcHY5EiXDGpi1L6vwp4ZsA3mRMbBj73KScK6AgtyvyLtMRzhjEdC
Git/jy/z888LHCzL6XEKSf6riiDuGGjgZrpIGHslR0M1X54hy6IG8eaSLE45ciMW
GrifzPVkXZq/zrfNuOyXBtiSV1CM4wiKh4xlswbSY/FfDbV6RSqHABu4+g7Yg+KR
FsNTg8uq0CSt8q8YJECQXm+W0rCkb/MUYCZS50CEeHZrWZSB1BDX+SXKGHDoNy4Y
FIyCqte1H/3WO72B/WmXch0C7Oqd+1p5L2imOtSyv0ukLxnuu//MltZb43AKLyb2
3LOq/Vql6LlQ5Ir0VxuqGee2GEy+xvz4xY12u/mS1JccRfksrn7tu0keoQIbS9BD
PKN74pYF4mfF2shp1pEBACbMjW6Nyp8fJL9TpT82d2ZT+zlbcnpNcxv66FPOS73K
2rJhiM0QezQ4Ph4hJI3f8Q55b/6h14E847YTT1Mx8r9sXKV+Vc0vp2DEfCEhcJ8J
fvGTomq3rVoiPqwjYJUpHN2AHUq5ZVzulTvY7S8tdBPasP3n9845Bm/nRThBfT1E
063kw0cTe4yD5RaAeWYDDaHNm814d9BuMoJZflBAyFeBwctcbMf21uWaCbDtSroC
DdiGedoGMSC5N7GT9dddn/HsMJq9aVVgKL53xo7SED6eTcn1rOhCJW8uBiAGWDWD
Yb24go1C3nA990sHWXqH+09CqjUUaKvtD1YermUMhAxMFi+mpoHp9laQINUT+kVn
2cYNz2A8yKF+iG+f4Nt6BDiPZNIrv8RaE9hy2B57x2+BkjY73q3iVDgGg/Bi56kp
CqTSnMotoXmvFTCW1gzTOMakCscJ4YYhYSKLE/D18cCcyI6LUswkx54mD6qvlPVr
HcHES9Jfw3GINqdsEFAhconYXueMG8eYXh4uOpr0kWKM8qr8udfU7KCBaOt5D8x0
5Xtday/zryV0k2xMTlshy1c3U8vvfiRLMzCdVTHUnnLera7Xr3su6+ugUGSYZsLd
S77WEhRyRKoQm1jHojHysIWsz3dJ9OyTXspJ55NVvMJ9Or8/zCemu7MDHljufIfo
L4/3LV+svID1vCMsUdJEYldgvdj/jGlMy/mLkmK3S12e/IO5ACotEUF98iQgZp1t
ylSjaZOFeMnN53b8lkwi+UWiy/O6I3sk9rHE4POwf/Ae+RXGNJ7p/k+vQYDP8piW
0Pc8X5Z2bum0Gs6bboWPAPA47XsxvEbVmgZwxzV9PyfiFzIKY0pD6j/oNBYNZ2TW
UR2YujYgqqg6sWrGfYVkgiPAZ28gZH81H98Z2S50ipqC7j1D0J4bLr47noD7Od4k
eKvwFc9QnBYJLDar7LUHIO6nmF8jzWdJBvWONAPi/7Bltrp+2H/NLjvg5d0lnt/6
KxA0GVf827pHiF2comg0yX2OgPDNXx45w/7phDrdeqmAEoDZSI8GT8PLwC51aTCf
NgpBjjSc8DSyR9dnQ9/rJorEUznkdxGBkGYpJjd54JxKKltBLcfGri8sn9673Gj9
Xe9WyGSamO3W2bt5I4/YACXWjbxzlrt45aF5K4fM2eUuSjK6aDJQ0PHeK+DkXZqX
dWf5L7UnKjxwIHbE9uokPvo7t8gyCrkoKQMjeq7DQR0fM+sl2nEQsC+pTrHMl4Wh
VHctoOCYVk93soikH5FvuhE3u/Uu+9FyUYgAr7orw5GafwcdEAobLy1BagSEXsv8
4OQcDuFhOgE1fMZBqd1P5hqWNMx/CRhswxmJe5nZG5yf07i6a/SdTTTWJROy6T/I
qI4EGExTA/XlxGt29cu7xxjSDuHEPy0CMpIEvV9ksNNnnof/fYgGYvBxB3JKJX3E
g5qPMEL+pYdW250CgKYX/0OJxljXGPZMs/H05LPHnQDD7b1V1ls5/ACrq8/MDNg2
+I4syy4ncKBO9QuaduSUn9rM32UaJRASj7ZM0G1RyrJu8F6Px2OOcIWQOwVFpUZz
Gvuxp6qitlGvpq22iEYrf6NC/JMQkJQ/7J1IPXPXtM+oRXZDdvJA+Dv7SrlHAEAW
nT7pWnTYBzDaHD9P340BhG5AdMMYYfq6pC54BybRDz5QTAMOqGXATf9iQ98/8DOd
Z8AuQEwUVu1KxQvZyh7ldMrl3Crh6eNntnCxIMTv5kg/gnlXGaDTEILJjMiabhnG
Cx1REI0twkQ+eI0BnGDrX61af0JGG9pOB4Ci1yqlcUzWhoTqBuW2QKgtGE15NKTZ
D1TLeJmZ/zHJPKjaGfM8mXrcQNqox8insPfw7ZMV79a3EM1TOB1H4HbavNImgUnX
1ogoyCCE9flwfK1NFVWluXCBHxE7MiMXdBTozlHyNMd5GBJuhfRE+1XKCQjyn71+
siorDuJ/iIUytcgNYgJXdG6iA0G9OSrgZsLNy+U/03R/A/JiuYBDQ2SMs5kfT9kz
Sp+4R8fnuQC4pVqmcTwg64yGRv+jQrs5+HBTn626ZkTBVC40tX/LctIt7+aEiaO4
Uh0jqsUhO5YCfHQebo03Qwn+GezXmO/DSR+ZDjwIeCx/wacD12s4D8MEew90s7xz
tz2svO6YpLckE+vp9IIFsi3kHJEqsY87k9qZ3lkQKkF4fsrbuCbdpxvuROJiaMha
J8SOp7b2396IjXa34kIv5ndAPhZMAMsjIsA2SHq0yNJWoy0D34IUPy+HllvvoY5T
srbsM/u94uCy8QuX72/qnsSqEDP4c+iAwEzFUzQRrkVF/STnXG3Ywc7jyCCZPoig
qO6dYHhddJS0btIZZofDFcMkgfqc2nrOij+OCHJftn65wtbxEQFVjoo+SrVWIVWT
ANueh98zsMMdM/Q/LB78XStH+F1+2g8KcIIybpR5szrfzJ3x7Rrcl5lqIZn4hrJs
6Cz+bnewKttIlFj/qWHtOYLa+4ASV+hJ3bgayzVG54hI+01Ob4YxBZS+ZT+lfb6j
i0MJAvv2l/Zy2sQN3LI4gZcwDZRTy7xlhV7LMloOhn+5ir3Bge6kSCU0HhMYYhQI
xscpncHFugrFheAL9GngK7YFFlijjNLv+gCfxvquMOzJQ2QYTJHxqkFpFBWTXWFJ
WPXiIQVCOZXw8wfKtNl+i9R/Hi04u5JdIyrbLNh6L8Ic7bLrb40kvgK4jzGB6XAH
QJhFzo7CBdn3DBBZVmr+amXvUy4vZwFiY6z9Oex4DL+yyiOGtPA1HCZ0mhpxF7tI
RGGF2/n0HStaWgNSRmEEpPKjmbd1z/GsnoJW9qxB9uCxv2PT4k3byQrimZ5WMFn+
D9J9FuyqphqjhFhWZzRdsh1ucX9fHFInjbbw6DN9hY2RmBO+ohcmgtM33llG+HQB
Z52coqp0EA7+oTnsn+ZS9VZtkznEa54jmdEkRZ0pCWv4dRzAC+qBwvbbUGV0koqJ
e7nAAEDtQ01GGQwdHQKCkwfO5YUfxlBVIKm6PK40WLzQkSZzRliooQF3kKkZ91vW
pCHLI0aW0DANyhLAZtKl38nN+hg7Nwp+lpn2erm1NTrgvq6jLa57xbdciSQlCYAS
NVHzKgIxQwbHM+6JA+joQr3LhOvc4/XVge1w9/oEoTKezTmr6Egh0KT7FLzktYGV
O3CQcAr/UbYJk1+Y5J6u2FmE7v0j1WIfH4Bf2WCnMeDBIliRY48KnRN8Lk5g0vM0
nz/ISlFQqfruSNIxU/dtMyPe4fRF8L4EfJ6rHm9nsyhiMJ83RueFs1oaSPtay41H
rY5CxvTB/RrnvCJBZUI7yToziZO2QEdFh2SwVPK9zsyMMg7kpb/BevL5pHTsh1Mu
yEImfsYlwy8+j29DRo6XqSsxlBqMRAxq0qLqJDogxQ1lOEcJF6nYZM1cQbzRvXe1
l7pIRNc4A1lLZMtftfHarl9x+Aw+FiJdHOYWd30oIgxQ47WS6o5IUWG+FoMricp1
IXLyiRSvBLOm7lbvOLkhtcSmloVfouuWk1NOaq0W9ZftGMRulJGdk86oBoCZyo1N
gJjhmlGV4ckQi/q1f7ZKCni8vlSzmAKtgjCqeUe5aO+RqVxnap49QEI+I3faKwuP
QuukKoqJukr31pPLIFJf6AWMoZwPnFYHlolUdJd229FTaHgO9mJHiy5vlr63cqhK
gofAtWgNlQw4gRPXmHslEUJ0doEE63Lp1XGw9x7sC2vozT/VWLA/o8YAPo74S+yr
+owskwU+igPSoIrL20VNMMew198NKWjO/zFjH51AAJNGRjF7LvW7xl9V6W1CBzn2
gfxucaOzvbkPpN87sI6E+TgQEN5ruwn1oIxivTrJ6IYR4fh4rjS7vsXcLeHX/hSV
ZrMV64V1zzIOS3ycXsbxJv197QDSTrOrOLUTYhPQd3S75GKStlgHzRG1hJ5Qhce6
W/ZNGOa52/wRlfecx4oPiL+xU11IHxXfAR0p5K2MH3xpwG38rGhCrXzFwZL6ds27
dXpbvaqXrWto5kbosL8nCUXAkUdNvPLSwyWFFqcpz+5uBPBWZq3EG6XBTmsLgBe+
Zx1EXmWg8LNlLWwF/zUg2wQQHre92kZUZAN6j4bvMmYIPF7K8OdRwMExKakWkGF7
VJrp+fhMVSuydaQcwddVMG0pcwOQ9rBITe9Jeif09to6HSDq+Utn5gqKbvDVncq5
ySoW/L9SCQXzB1T+ECB2h350W3co5PxzJo7NcFvMgoKQh3QRMlKsFhphkSzKTQfO
iWUPBlGncVquAnjSMePfnwWpWOR9PxNpBTAhFVbGMjJS7GaQZGxcZ/9IsZMwAGus
gQLr/8/dfoNukRbiexmWYaeihvo0fxHjrrYoehFkopeU4wVmZ57oapRB4iqsDkLm
H38u1/ylGtK5tuQUkI7Y95EokZp8ztlXHcbEqvm3iFEVD1vxyQN6DDsLDaD/ji43
qlnaI63zBH3OqlYyp0/g8PLlgnCbyYzmFaIwVR+NSe7f4CLxi71Lu+C7lC2Y+ZK2
e2IgpFG7OVMh1L9B0miacufU8YTi6izpVyCT4SpaSfhbliVytm+MpvyG079K8FNH
DHEV1ejvhScPoDWNExzmB0w69z8xgX0vA73HrXJZAF1KOaI35FWC+clnCg2LIP3y
hKJnoG7+teJPymnLKykfc9QOMQJfT31GPsjL/J4nWABL37Hjpi0Olee9Di7X1nMG
X+ra0XadUTy6i40wrLfA0BY0Dkb0IdoIvosDtBh3Z32OaHtMbftJQtB90mYGkPV9
PlybpiYRlm22R84ZeAYDt7vDFT2fcKNyOBSgeJ2tlokXR7Ay8cT1xqR7sHUaPMo7
5LxIkZAZ2erc64LSSRU3KndnUMRbPzmUuykzAa4ax1ZR28bjelOwhDbh+JcXdUnG
fOb/K3FwrMYxuqxDmjuZ2TiS7/9uZB6cyT9AS1YdS4NZIzYgbSDu2ibxNeH1ZKV6
a9+0wITrAghiXJFdq93iJLgdby9uvmSfWGOJ52MJOboFJ0QkPcb0hZVRZX/X1h3a
dRVtATXlhUgf6HR9LQgWOhfpke+t4N6G4Xypbo2mzZX0Upedeqxqv2gx6RyJQWOX
MtOA7WXVxOWC6oGHCZY/Aa2ZD33kZx9zCDcgJ5N2/KAnU1BPmAaSDrGgDJ+Focey
ZTeALylQW/N+3kSFKH9LaVVopGEPqln40eo1P5dRONL48OnWRwC4s+gPSHP9wzrQ
BjoY7o/2kjMkFsICvaDPuVB/C/e8q9xvHgLgo21DFKhveyrVDd/7EFBbGpPwQoom
gOP9R72esuCpQph7E/Zqe13xAEF6wEvR3y2wLAKzerWeFZKBuYd0IQKB0Sw0vAt9
M77hPDks5ElCpFfyYyut288HYTS2KzoyiVKjn/8qRqhjHlPlVd6r1ElHqFoca2oL
acSJWF3bqahNoksjGZkGXUaJDXdlys2XYXoIRdc8y9JRpgAh3oEK5zW/iZiJfFmb
zQ3M8l59bfvQXSfv3DzMaLiYDs7t89qliUGHm/+9DN/NemBngptPPCy93VuuErVd
Och1EQPt0erG58+jKOCiHd/2CJtO9jA0CpXIzvtZJPMFyHCAMC6ulZ+7eCZdUaxW
4gtcf5VK+XQR1hh9qwzr4oW/6Hnx+DQ9NxAqnhQZq1Vh76WCn+btcOFGvAaZmGTF
lqYviGNNp4HabPGkg30jlBumdMqzPrcYviwwgIN7kRvRDPtGzkb49AlhhRMQ+5+1
IfTHQLCcynMF7yQBT3MQ4Wj9G5C8p0A4lGQM2pTIOAO/Z4CaLCpLJKP14dMCTlnv
OyBvVVPSawaKSrcjHQ2gZ27/M9O2+Ad6fImy7gCvO4kHJ8O9TzQYMQ465hpwZL5b
ALwsNIBxFLn4zZVbA9hPOnR5SAx15MaG+VMzKRI781YLtHxjwLVELXrvo3N19kH1
JdKTak9g7myAWC8gyR0iZnoy7x4q9zPOihH2YmjQALvYY+b0DBl45wHZyXZvKxn/
LL7ydkEVqz3vNAhxVXoj+Tv880F5XKcoSPmZTfqfUBFPdirjaQYNAoBZ5qQu0InM
eZAaFGLA03djbGAr+PpFLvun8/GeJwCNhDl9sWdcaPR+ZE2BZBpt2XBtrpNMaIGf
hit63Stu6qO3ZeKSZ0eWBh1KuVPvBeyq3jEW5e+FwSCu/fcmH0jn1dVE4XNNlaJG
K+B3N8qnbRnSfmMAzllp/2odYlZMNyNxT3YpyXlMH0z6QJFVNX1D9vx2dvnRHpHa
+RKVZESahFGqjN6rcVNJC382JaB07usvuy6KNi28CIou6V4D3ZwxpoXoauKsS8Kr
LUrT5dUZcaiX543gT7alqohMYMb0Svnk5uB2BhYPC62pbFvFJEADdX0sbH3nJ39z
CD2gV5Vfj4Aw+fOdgZN1rrH5to5RLggT+9xZf1g/ien5dfrqqt+WsqKPNVULjzGa
BDYNnL9Onn0Zs4QdU3QBnp6VopN569wH9oKxqJzCpAFKr5tTVUGBlzrRRaxHEFVx
v5qnl2hgn+QTE+FcEjm6PnpSja/M2EHjTNFjf28zuh9rwGsokMVktGOXdrwRpYeo
r5QVjb9ubXz+1PCWwd+avEmXiK/4BrA35OTmEPc2sgTrJz3olnANMWiKmx+4iznz
Cph05YfebwWJxGjTYwGlwrLYOLJp1nagv8MRCjX9tDwNQRQqCYp6Di6ujlnq/q3t
VomloA6sz2s7PfX8k5Z2DDULcjAe6z1RSbd5jN7+BbsgRNJ6KkhBczNcVLhiGAHK
FcKpd5hjmMn1n3aAW0456zXwDyiZ93Q+odPAaM3WeFsWTs9iJ1TfxKTI6O0hpxFL
68ar9ueWjbk/ILuMXJgiH2EOXyoVZryrVdxQN+lfLkOl+RVp4lPvs0ZGvrGMv0IU
AwuStPQah1KgDgchJ5T3UspNyuoDWIcdHHE85EnNDiJ4o+xK8IfQqUL+VjE4trZH
MOfMH9ypBn6zSlUeDnaNbJ4ukxgo6a7GjPs62rVrov47ZXBOtiCgRB+sj6WpA4cV
H8ceuktcq3Du1DY5yp+U/MDgqVepByGl2RbM5z+u8vgipakDwvPqYddns/iWN4bY
A6hLNTFAMM9b3qWvJ+BY0cgDEa2fSZGQkp2iSRamXM9Kfd8eotyWZkmFVrrV2IL8
5aQD/ZrmrBmHDEnN6enamN/040cQiszIK/7H8PG3fansGtVKV07Ilp4R+A/0WVe2
BfAwro4CkqO1+1KVjYk60btuSFAZRkp58VW8OlOAVc4fsGL5xPIBHag03DPVKaJk
yum7XdiBQ0ogRWCYJtrJCH9H+GzDiOae7PNb9V84pfue7vaxrVKsOY8Ge+Xdxotw
82E0TWlAONa0M0+1kn1FtfOaB1/9QueXEX/V6QQycz+LBwZJyuoGKpcUKnG3hVVc
xf+wRNE+QfESV8BHWj8FuT3ApEIOGfAX6rjz1A4/Sok2hDvhwK6toIYRlZwzllpU
sDnRdQ3YzmAnXmWrTb98oIkvkmuV1zrFfD2SYcQhKtAeuoeT/2FUwOCzCi+7+0XQ
BleTk5a08g9UtDLKevMKD507RbEV1pLT1JQ0ckBqlsETQH/SwqW9NweWlYIkQ5UJ
R+cTod6r/ruyD7jF3tjTTfMCTJLbUZzzMrJBd3w5i+g6GNFhphFP2xWf7vRtpQcb
tFL1BPBLmmn8Vpsau3f65HoM03mILyudLG5pB0DUZtuAlaRF53femWrYvHNhgy5Q
BBMWW57PUHhsQQHGHtTLr+YkpzFC6QLNqrDAYC66XiYpT3y+796nJwsCEySd5v95
QWoIlgYJLi0G9fu76YiQLnMJRLBA0Ef92bFJ+6v68jwVIUpDAIrBC5JY91XjWMvf
ewZxVXbmhVf2XT3UdmzaJ9KYju7a8drvSWK7BrgSetchhUgw9KS+B6BGl6KAXI75
HVACWtdS6YlVoxAjE2TOTw7g6q3lTfGvWEnnMw65HKQ6IB01U1tET/zminYXRDn3
nzZbe+IzgvnyRec+Btj1ks2CFhAYTzrwvyPpycjMCHQiFilrWPCCaHuGZ/U75kvo
TZyYGCVwNTJyd3iHcaz9EssGAVUPwXGhpyMp45hDCxPxlS3dl/VGv05OuUu7FLRV
KgdFi6X8Oa1xH8HsUksKZ2FJGac9RsH/BPzA/NX1KtGSt1mNw0x9U20S78Q9cJ/J
o4WB2jFOAON2ckMAM12m0EamxstOQ1eHpc6zx+LVuwD143zj/q51sKxmC5gibgxJ
kvgDisKqtKVv86vC/kBs8pJaVaWF6MH+JOQNIrIINOGKqSDty2pyMSER9N+AMCj2
OFPGqVSoK6XEMgODD98R5Gx2rCy7RBsxi5OMZVIgefBbuuIQG+iB241D6t3pyzbn
NiJBknPqurqlh6KKJkpzZj7vStAcnuCdWkupvFjF1g9lgPPcmQFW342+OYj0KfQP
4oLKIBrxP9IZZlvMp2TgoXKbC+gUgeCkyfFIHG2iym+OTztMVZ8HLFBptteX+jYL
/xxjjagrmRGShnxL7IMxylIj77DM8W25T9zUlMvEG92SFZ4eOipib9PY9AjoKEEc
dRS3fmuKQVAUIbtNzxlp9bZPqHcQoq7PoS9Rh3+1tap+uIsq0iAcxOWmvw4LW4rF
rD8DE2Ll5GS7HBqx06W8qfrDxekzJsnz8UiCFrMyQoBttrK2rqIrSM/hLJeU34R4
0yZGCR5NmgHimoSwX8DWrUdRdimtKDAr3WtqaR4GhZkk7mEleeVEdN6RiwmK/RMD
fevwepXite5BB6B20L6+1RkD87VpYsoguqa7tRKuQzdgXl+jqSnNR79xYfxc7Y2S
BW8Av0H50AxYnol3a2D0do97zy7fhmvuICsB8A7jEWnwMw4Q9ZPB0ZLrGyTUpYTC
iQyM9r79pTpQ5OHuBoDOq2HnQgRQAmJyHIKfpGsMg+CNwmyBo7UoZHjvIjqon1aB
1/ZWTQn9gyLvaKt/YVrOZjbgbjvL6h+Wv6YXNw5xtJv0hzkimHX03i06GoS76rJt
fMnq8VTW/obiCW1DPvnF0EU/hjWCPgxbuwyTvBRX/b8d9QcdeI4ReDNwjB3XuFtV
LcAW9iJ81HCQzd6pRL8juTfpBsDIqfFYKSkABM65LLCLR2b6l10No18kTvGQZgx6
14QYEb6FRWj2uOH2Jud4ODoMCbBC+shKVd6xERKEjTkSY7wbKVIijk+/pPOKZJCA
3xVq8P35QAXSYcKvTykO4/O1v4XiFWhtachb3UrFQD/X0RtU86YQYdnn3zKbkMt8
bRiMMgfL/4Ao5f1+V+i4vdbE9yrkNRao5upYBrVshK8zFmbc6/lSKRvaZxTXxfS1
hkyge64j9c+kYOzKu5WqjJUcZcsNOVnhW0Ctm4kADepU28Qr4EArDo63u53QAXIS
P8vPUjntjQciJaUZyH/FCz5PGgWJ177QWP1Fp8r+WEN/YvIUE8ZRMjBDO9YLBNK9
JoqJvqrq/1bcHA/tjiuuLrchrv7hxYLrWxYg/+y3tTbKPwsvshovD/qxKIX2vNcl
dhLQCmpdJJtX9rKF5Elu8pXZzXhTcpycsgc0bXTg5LitW2tRg5CkbvUxAhJibns/
0CxTDO0kNjZ9YBN6/EZbX/vIub3RWmOaP+G4/R97Bibpj3KLDIQS3+PMqvyKPiit
ZLBtktpr3FeMA6QUjGb6o9sn/rfQx099nj7JwPufqi1k0iJnI+iuk4rfYSmpEc3N
h/rX8onYeWAia3+i43XcySLeroqZI0/e6mMszxa0PGOzdjwcyMVmpNNIE6RA1JBs
xVVRc823WmcBF2ojk0KLvQr5zX7g9NmIwdKdN8yfFKVYhoe370/I6FWDCP544eR7
d4pBcSF7C4wJ/8hdW0a8TfEIPGk8BQ2tKOU63C6kv3wzUMf5Ea+VSyJNl1BPDVO6
7Z75mgCgADd/DkqGU57jPawx/ZFnuuHlctUCwiU89d4s/EmAs5VSq7PyuWTJ6SvS
RlB9w8W5zhgR7rugmhswT1bYVGOLHtOy1O8eWKgtjIPDSfQTHI+LLo4EU7fbrFux
K+O7WJsLO09YBEpUeOnVRUKcPijwGJTtABTBKd2xg3kEa8xVnK5ZS9wySHYurq+/
GGcGalW/3JDy6h3bNJUs8RKzfavISAsy7es7FhOlEe5dlipcwKs0BtoYW9idWPl1
708McsX5CUFBz0pNHjLmNNugJyARk7LMPIQqwYYp8iR8P3hVzb8W+iBc16eIZjpU
GKtwk3y3F2L/uifjOLxqu5oZzuQA/u0gzt6LxoBlq7ZuI8wBMCYsr4UK5+c2hPAd
9BlQEjLXWXKxqoawSRzvay8Ptjrm+WntdVboNN3zHLu8t92tG31OQOuLbXvDlcrx
LiGj7I5pRiRpQnt9d3EbZYO6KXxwpZXJjxihv+c1hNYa/BcIuAPdgbeYXcgJqhjw
l1m0xsqsIQnyeW0DASdnssOt64ogYGSoerH0F1aVs42bWuKtdKHAxi8JPshdgWze
CxnFgHR7jqH24tWXhbWJ5xuHYlnJPcHFzPftVMf6yKeNk3EdGv1TKUvLpl9PxrOS
YPZj5tgJNJTLHjcj7v6Ql+pDES+cJ3l90ITj80f9MbkBuKz2Hv/g5SPLatkWQMaH
aUiilc8NvRXYsOtw/fAMAAyW3XllP+Zem3jd+FKioZMRc7qFsY/x7n9N59y3v/8H
L/o3qTw/rgSS9oPCMgoivOtqZ99n7S/9QWVnSRIMvqFdxMDJlT5AwnRIKZ00axa8
lLhFyyZt++RTvKN0MeRyC3+0aVS8oku4vAKGyMgSKiK4388W4DrjzdcV8k4Ffk1J
uoUtkAKpjGmESNr9Ilz7yQMjQ4ndcE7vMUr2QW/2bzrEq+le+J3rzEnnM9n3VdzZ
TUdvZKoQWNspfYvRY1pFF9YhYD6oft10Y87h05wBkmtL1Cx2/dOJnwCFIuBKP6sF
qI6GSEf63U11wrZBc9qxsuxcN0ez37fAWANhm/fuy7p9wO22ok7GwAy+e+NrhjmB
I0AqMCSCgtI8qWfkKYccmft5+I9c09POFpVLqQdWNSdr2pK3FtztMpzhZw9MJN1r
4Zt9xSfw+ai0apsdleAFhgkPFw0uDfIvafwIJPI7k6MImOAxkYOsSwb3AHTdWfrr
y/pSAmP3pLCNIZwmlEJ29AtbIEjfnw5PObXwHYsh7ANXYUiVoZTOEYvVOnKvo0lC
YoINuZy3dd36VZX35zrUWI8TE6wfksQHVmXOmsIA0RwFxLstyjgCLiWL59rqTtKP
IxTYTl7xWB65V5mAd0BmCKEPypyW5wAWMGkTVnpXA05C5qsV8SZoFktJ8KWfUFB/
/ExEz/C+bXXIT8pXIf36m0Kr5zNiKv9ToaqX9AaPGBpjHwz5R1sTMiANL3h5qsax
utZkgY4j4gn636LBT+QsYcW1i4xgMcrPWUTH4HMynILEEpBqQ8D/txdRQ5meOzDC
CPBAi/RMuu0bHXkLaYlbMq7PIVZi31qynedOuq6H8nJo1Gg9dY31HwJY2UsEeklN
riU4BZ+1vOgtBp0V0TehS4lZMQ4YZiBct2HGAqJP8flQZq/hkwWf2WVSDAgSdNWC
LtSqi2rwTzV6nHHBuPrLfpfIGNT/Aa383PqUvqs0zhGek1RQcCCQfTsjuit8cAuD
IuJJfNJb/kublWawleOcvpmbu63VIbncN8SkB+ZBE6UPnJpGDh5vqRTKPgvNiPlQ
OsghA4TsFYOmxtKxCcrTrkQYcgtu+cnbJz7AoCqIHo21d1mk0FYfV5rpPqkEWQ3m
sDE108vzMsJOql4I5wO+M9giuXM0C2eu9bZkdMf7rJSr2DhBK/vJ/nb4xNcJm0oE
0PKWW8U71dgC8FWulHPgZ67n+yOtHoa8bRswAYwzV8VZxZ4o8kPd7sEs9W+aZMJq
JXy/7Eupm1MUIUdHuOMbNSMevMsEQq4ugSeiBsdu33hO3yLa7/LF1lmPfyii9c7E
cihLmP3lRCoHIT9hg6lR9O4cU2cl0fY84fUmmKniRc661YiyRjMOE5qxI9weemDo
Wdccog7Xwtt+2iiQG90TSjPpaov3Xe/N2UdnK2+sU+yVs0yoNLNXusXpSej24UBd
xsh7WG3chKIStBNFy05NfoS9bLxYa+RbJevlYC4qYmJYA9CUEOwOMPjqaqlJuCls
binbnpH4FeMoT2m1gOq3fuYuJmQb3ht/SaEj7bpQ0h9c7i8A0912hvuuJr2GOl89
bPnB6OvPT8hvr7v7iqixTW0RhQZTB80dvBUcxSD8fHg+8uCewc6+m/+UYR6UEP3k
uZj0EheJau7ukUebntyRy00YD2yGZZox2Ih2UcsBTSBURE5IFH4TuBXr6YTYZLXc
PQfz2yx+imNwBtZ/LG0AdkvKj62xSCKU46eTSUhgwXAk6u/fp87c5MBUjJ40Mmkh
qeRZz2RmPzqrITPVXiuE3JV5vep5Z6pcJ7mMIqzd6hZqGWNgtkdExNmHIto6AzIs
AD+J8yT6qrz/GkWTYq0WZxanbG/oBqPqB8wyobR+uAQmay/+W43/UfcaRm0Dn3tK
m+rQh3+Ur0KLYayyTdsCvkObHQHnsr/Ogs2wGuT72uBL6I5VJXhX8DL0JVS1WSxG
U/ifVBF3pSuXTGpK3Np0zl2Arvyt98s44e4z3/hkAjC1CHtVSY8F8FgaX48oHPsM
OXc9XNvhrOCNNiJy89OQ5emR4m/O+nDrdYcyvS5IVqEu8nBrJs7joRekUhSgPw5k
mczU+GbAf7qQkUmaeUD2uL4j5RHiHJpQjJXUk2xiOoaTxrANUGoDD7cT9sKP/1yg
KxtSCjFE1SR9BmuEwGY6RmmP1+7oU3POhWPt4o06jORuSEg3HtNBfzKQOzqE+kYS
veL9Luko0A5UyMqLevsP9JAqBIY9f1TaGEm/Cv6M447Yk2edGLsjE2AO6P3TEhIs
9N2+kAidXgbTcCkDGGRzztcd7nWYH6J3Ae8p8id77iH1aRIRZy83FI+bFmt551f3
PztyWvjXIekoNXKLR0n7FYlFfID5sXN/S56+l/JNO7FAf4y3+pYgwGcYMMwXXsAx
k9YncgHsQ9+YG5efer6xLOrPBOaeCamsykOwBiBJaMiIKKFFUhIEQnAbRanJwI0Z
IiONQmvEj4+FjFfTvbaB2U3xrSK1xyWgG0m3ByQdafCnRWwQohnzmqXMZDKSErBy
NkU+hsjK7gy+UX2EMy5RiyHw51sPgo4RvhvU0Eid/8NE3rASloJiXBb5Bxx/Hulf
a8buj13V6mHQomAaYLjiXbC3721nReoGW+SrYakaY9M0pmzICtEu2srPNbOsllA3
hC/bFDzOsLIe90MopdzhzIQIjjm9saIpB4YQm5pXbHSJKweOau6Ki9QV0MRwQU+J
11ONxvm7tXVw3BebbstowdRbioG2wppd8SfwSdupzk8drCSnmQz4PhUpTzN0qgW5
VfhoPnqNu5DLLXoJQQjphnxluwiMpG0U/VOeLCXgCCM7EdgIdficyoOVSkXA3Jeo
73ZaKE2x3n2URCWaS1diowjwScteh9lDhwiQPBIMTkPioKpJpLx2k6GVARMbXJCD
N4frEUoDF5PbheSpRgsaG5hrXbU4e5jJGdssVaRLTjEhPPGQE8es+hcuhTTk+I9L
0V92saJzcY0CI4gIfLUKxtPGTfpjUZzC6kHPgYvg7oed659VLzMKXAT3w/HPM9ww
3vDHRvxkidJgAOHIJDB3g8LK3lhhDJ3MTKNeqllnqkIkZgyyF+T4Gy0Ex+r/Z6KZ
I7xc0+oA8sT3ghDdjuuRMxPeegAJHYwNRz6/Kg6a3uJ0ke6Hp4sRYT4PaylrGYtn
VZwIkRO5/sm29qLCwxT5z89IM9XKdmtU/kosJvyNGzQpL9hPg7nCvMq8zwB38lEt
BDb1bR7H955XhLcSy8S9fhR0S5e4zN5HJFXT3mcF3mzCzEIEwL+aDU2ujBV0snSU
L0/pXNg/IthtBCiCbbkg8bg9Gg9Jz02kAcpirfM8R/k9K7/nBBUQHOwx2hWDG+H4
D289Pzi+SiStGyR2vVytQeBSXvbVezvtrydf+g1E/2M5lvnqy+4X+ld36sKComnn
dHuPMdJLw5G7UhElVR2R15HgEQx6j6Y2xa904LbPbrx+hx3w9MFzp5VZXLLLtBoC
bg9We+49mMeJJF3h8t3sVjn6CoUF3ygrv1ndh+XyFE2CKhShLvuHoela3jsRhWDI
GihIEtDDjBW+QXZkXDG8CaxHDgJP1RUsmD097mJ978rDc2/Nz4Dnw2fby8ZyVBjg
oYcaokP/S2vJIs+QUUYVq/O/5jvYfIaZTTNvRPXXd541VDAtEfR3b/ZCimLtUNhV
gZcO4pMQZZnFS+Bi6G86gQCd03pHAl0zi0EIZUNRXBAkK9egNo6gBRToHP5F92nN
bDJBHQ8TlWWHoltY9Y5bL3ck0Z/KUF9a++w5RbnVK1PsXbqFNJ5Vjr3ujtEsFssf
EZNH5MxV8bUB++7F2UtgYv8LesdXGCJzFumFr85OWSWQjtlkMZkUBbKk5F2Us90L
FQU0e7OmAn6eD4tTVlMrmLlpjcVlCWnG+BQIyB93wcA5JiM8+WHvTPXXByulT/tL
qgpdPaxEyznAzwEjFXrvE2F9k11ZHA/vWDBKTUiI7/2KWNH2RA5N1ojZfp2v8hXu
DjeFbGAJRKoNwQGvTXpuuiT0NH2kiKUJ3Sye1Z3nZ3arTayDHxzWcZ/9hb4Z4TBc
yk+4e0SY+qx0+ojxZ+QUfY2rMC5W8YpBGMG3FOEkBgnkug5NXwmHTTS+Pxa+z0Gc
oJsNumcyOf9LWxgzK5KIUKIXaSSiZlkbj8NcY9X9GGrcPAg9Z2MROwlqYI+ZFLBP
TmDcxp4ZoyvzkfI4xudoqzo/SGUycuPHmJtddvb1Vev2y7xDLc0APDwwcfVV6qQN
rat/TSViyW+xa4nxrmQh2RZTcVvoH34RLFCvddvusy+DltsYhNNwmsXCekG5cm0q
ybqkb6ZHMnSahrNDA7sVSOvQco3ptbOTFsikEwC/ixO10+glWhCRO2WuQWseg4T4
iMEQniWZLPYuTJDsQlJm/EgMkBY0TLy2m1yl7yJlmEJWv8pXEdXeXGP+wKSTaTxg
mV4eAISOQNoh7/a4jZothzQ7zGIWa9u0W1XlnRoS77qWoPfSWgXQeYc7GZTABz3H
xdq0vqB6NT1wJlBoKY91m7CCU1iQQDG1DDZUezq2fFMltFqF2dVnh912XMlJJAOF
ULil0Owu1fcCKBRR2PF/LAqgbDVfP+DG4yn6+zSND0wmOaBibseNUWPPpweARNYg
5ZHlyg/7Lh9+6B3eOrGkJB3NrCIrV4Yy6nv3R/GxV7fGU+Lnt0ZiFRGsT/9bgaFe
1FLJ9A1OV97MICG3mkJttV37TDLXwPc6IX9taVGzirWGuUmFJeoG/M40yCl9h5uC
CT+r7PpynERK3bwfXiniFRqnUfVFJrGZow1TuTs9gfCDsar+9ObT0wPLexKPF5KL
m/cwrDCovRnBFND9MCna8+CsSStYDZil04S0IQlul/wZYSDh9KkRy82PnW1C2Pum
2tlHhlxNKUXGGP7Rm07nYzmga3gw1XOFv9XLb6/NgDuyHudyDDbrt3amgBAIehjR
YxlG90vVqiEelMgzxFu5AM5Sj2wRS8yJMGZYMpN14qUoNLKFAjG8FJtpK8QZID+n
ygbn1tRixAfLKbTNQ5+yibTtC5UUi1ZlwozLm/6eYKsYTdTa9TumGdtIiJ4Op7wl
cqybzMcRerEl9lieXZr/GCd14wmakOw5sBCLf+zbvUIMxwl8M53XwOYE0dXzvsKW
wxTR/peu/0vEjmlwgM3EjyV1wslkCCPRIBsm8uXvOcK7iphBnKdJQF/Wz/04o6NE
qh2Lkd5gdaEzLwdSYx/52ys7KwGM1xVEnAaOYs3EcKsgrU6hc8bvb2G6uQbLpfBW
7UN8K1rtA8qkE+492sdmuwLl4XbrOsCmOgy1xqZh+H81PS7fFKmIsccZ76KaKRCE
K5O5+jt2Xs0iwCNBLugbmy/LW77Kd0Z6NQSa3t74w/pFQyIMdlKzBmrEDqavMYl2
5Ce/kqLc++DtD/YMTuURaVTWl2ivJ/jx1eN2MSiLj+KgbQaMFnM3KJt+tJaNYlyg
oLac37NSBbUVqNBgaOYP0RqM8u0X1cFRRqvuzIW312Vdl2/nCilB10jxa69ZJ80p
+DDVMrGm8sUcDgsO6giA2Nayj01CwQm4FRcGnXDWDdBqv6z+6NlqTbiFFxsaMGXZ
T405JIanppkZVjDdP5ezx3b3d5mEVbRoksTTWqDJIx5+lzUgJym5thwknv+ahtSn
+aP6zv1szvLcSg0nGtyOZczrnSrqkGzlcwLfD1odlCkjqshloDEzJTWC3OWrQijL
vlD5/SN+7ZCJC/6nTrtxcaoaz5XtiBkwovo0CnvaPLdv6s+c8XICELiM/kvbjQiP
R1kv/F7PwVo6VeiqFzv2XnxFeqTjfAR3saLaIVm5fePM9ZIxdqWZbXGsqm6MT++U
P3S0HsMcQ9pPV9GJSzZcrXB2KzLOnf2yr+b4wbicn2GldPiB7T4A09hz3KZ5pwkb
uNEf2eS8jq0E4KY2+jHqhZDiZI1CALsuC68ERFO2BquEXagp0QG5NK4CdeK3uKL3
CUhewgAWJ9XMgouhUN1cHOh59MP/TBj4CEhz4KXZdO2QbZoRTrdnxrDeTB6Y1TCa
Q6ZDLM+MRr0AGG70BHXXVdcIb3y4tQs6fmtZ0oBFVX4sxQqAgxRMN9ujZbCHQWa6
VwgYq267D+O7TA5hx5aQbQfOSsJD4Zm/CIJSlQCxQ7ScaGBWGXSSk+u4VGWFWy2e
HC78gCYt4se++ohiHWXO9Vnp6jH+XfzwoBlg2tfM3mGaeWDOLBKHc+73K4v4xBIW
FcN7oHorFg3H6nF9keIQUN1ewFnblOlvzy5SB+AJ0f7pnJ3+catvtPRUFS4c36jJ
kmf5d4zSx2PLuGYjQ2KVzFRcCf9ENgB3Tz8edeP+lY2UT6qL4Dq4BU14aY+hilWg
X5ES7CUChZDP9B0/5KgPiTsoC1TTW5ntTWfpEh6xbB/8mfaaXBzCWtISg5PC6kBx
UkQ15sVE8YXJ9To2qA6hzgyvtaJ+XTsybI6YsV/eA+fne4MRdeO7SUSCkWWPlRlA
RzLjhRzmCkbJNUd7roaeg6MeedmRX3srJVPWfdPvjsaOpeaOhHVB/J8Ha6n+W4ZE
twB07iNFmSV8NXYLmDJ5EXz02i+gG2oZ+sn2UP/yPVANdUpHnVCWSwo54OH4GbP5
ugkjgWOo3i8I6lqYZFxJzEM+66OzIA+cNsLgVeENkOr9es+lDZeOKm56dRZZvw59
qgeJLWKAMtefCM8uWZLwelhc9i22OLDAJ3pAbBHdU0xN/iq8zcKuQOAcZqPutRCy
xtD/2uRpZcWIyyQ+cjepZpJylDe5IV3dwmObsOTRb3oL1PbZ7W4RfEKZTcVN9QCF
+Mg/antbnfzZPKVGlNQtbin9be4uzANGHZGxJ+k05CcThd/otO6wdP64U0TD7WV3
CsSrSPhSt0MKEC4ixsnTDYzbHyjyY3lr4HR+y07r5aGYwo0FkBHBRoktTCUe+2Ud
t3GxHksQNav8DNdE3Ej2smf8LuuzhNTW8c/zU11n8P4cHt3gpZlJl1EypELZlE5i
Qn+/t8rW3kHkltg8H5Kc64a0oyFwYqKnrKqiw96tJAFeqq6xorASAROsfrJDEkhK
kwlCQ3Ya0AOtOOapU1wJ6LyvO8if1vyIxk8USrVCcB1c8FcIVJIuA/jM9WpaHOnb
GqQ7iyPbiJBDjcVJ05ZzRqAIKQ895Rz0/Kzf3OKbFs3naqzxbefLqKCLYwWxPtvI
GbRAt+mzwje0tWHno7ge5wbDpZg/7xFTOamE001mV6Mng6MsDSUkF+6ik7CAThgt
WpmQONnNzaMO0Y728sXLXcKWVDG0jUy1Z+nD27248rnOYHi3A3rw7KUXaNyu4Q+6
dsCxHwT7RsMpBMrYlQ5y3LYtEkRh0FldBrjG9DTZy3kdx74n1lbfsyNjle2uXkFQ
l5UKkqq90pUio7LwIAD0Dbh415ccagaPAbj0MC6jeiBxYHRZHaGd+v7Z7NaaznLN
ewlI0jhXsuTXraoRfz+RCabXghpf63cJPGYYoZTNJ2Kd/r6JwDbur+om2t8HjqSc
+Buj0PaHPV3NuJqcl0rDQFNNAFZGUeq+GbE4nWDlG/TZMJd+/CnB6NqoaWik+JBf
8ygf7tv7+sGf/08kuR0h5wdfpNKLLnVDlHyj2WMrPERjt8MVsO9b7IwwMhcsIAvd
C9S8H8WkHeL2GzSXbkhZ0h3cy48MhzSqv5VF+5WR4kwVEzSy8zQPF12RBlg/n7Ix
eS/l5Ixat6bDmMJGYnRtmNsB4cYTI/LuUj+NLzJXJF0wPAlG15h8hPGT3Edqclfm
s2ya8s42MAi4qvWgQ5I4LR59t0TREY6BE6lX8q5Evz/qVUuTmWsFw8vVD7eq8mL2
d2O3zyjzGkJVkkmaYoSZJOXZdgHDPR7hnjDGpeZ83By/z1UBWX1j7F1OfsSfDsSm
uI8p5ZHzw3bAbMbVrFhfSmNv3HeiT85neLNPi8kponxZGOUcneKVls4J8uuxVoo9
sibmYA8qngcc9m11zPeTxQgrOHMJr3KjbMi5/SsQzCL/xbUHnByvqtlOS/M8Zhxk
f3p37FoQSf8RplVoLlnAMWVnh3XOCrA2WHhbjaiKrmuiah0X5GPmMj5aLCI5O/Gm
SLn1dfxnykVRL5+vO2+rixjejCzZrLju/1lcv5rF4NifmzQUWZRqulYAWTkXwRD3
ZbjUk2JPy6v6OjH6VQtqbs7YZpG0/K8UTD0BeWK4ac4ml7k9DRPd0aaLAEoGB6Rh
bbKDE8/DJK31vAVI5nlhISNq2BRUXLJnBsCjvt7G9s+gSUpspELYSH68SV4jYpuR
XPW6SrmZ3pc0PK+yemAqd218J1YoXYf3ATRe0OrYKWTPgFMZ/adI4xz4odsUbFno
OJ/Tym6PF0O7UP2kPuOwI1h+w9yKSR7xMqQF0wN8rNMFTYjpU7gVN5BW/lc0/pI7
3EREFk2bp4ca0RH5Ll+m5pl8bNIRYNfHaVbqeQLxzYBDt16r8Lng4Umjykly6Qzj
3Sgy6yDIg1hQFZb3qnucnEj5AL4uyDPGWY7HytqxiMF3z6oU/BE7CbQeUI7tWJcn
hReUJC+9wIFWw+BmF2V1bceKN8nQVWhiqjNudRvKDdlis1ZeQQOqKptcJOe4LKoc
ZJmesupjSOaa7z5oBMvUnVQzkifRQMdJdG9n1FJP3wQzBM4AeZ5OKr5o6M8nwPwI
SlQHL8EIABtj2de6YpKbxjtZ9qp8ZyRvKZyMOQXvQNncKKScObXGaTbRImS+HlmH
LMwRGnlw/BF8Fa/AMJ7sFki7D+rqFyScJ5Lbcu9alQLLLjXTYkNxLAVPb4XLdxi9
MTvY7243W4otp31xfkh4TnGE8s5IPy4ffGk3KuAp+ITerHrBuseRvmae2QhRLO2o
fP9iY8sf4Snsp1qZOy5sSotwQno4Hn0GkRZAnmB9DhuLBtYbqpehYoaMkDRo/zlH
EQoqvk0s2Jt2Cusmw05xQ6vroikAt/fQLNsSxV8TMDnHR+vdDPe/2bjv/vgiisjp
ZkIuwEJtYRAufE1YR53CTaayT85hvvI8Aa1hnVw4qF3njRV+6j/DrkDRpw/cTjph
3Sik2vhhVaqvJSaVQty0C5dyF2jjpEIO+3PuvbTG80VL2Rt2e4vm9eQWOafLtCSc
4M9yVGOoCGZ6wJV9fV4dAjIM/fdSjMi0x4S70ir2XY2lk5eRmUmX0XURVxLiVLov
1/yENMc1aJQt358Z/K+Spzi6/dL4l7q4WHzKoLcM68zXcu0iYTSyZxd+3zmf32xO
HYqVbzHJig4PuVgFb9YCk88/gaAGVfBK0iH0IoejhxsVsxG4CBjfusPdHUY3KrDh
DedBN4XetN7Hpy7V5TvoZwHUpMIWNyTDYDLhwK0/TcdE68HcFFwBfBum4aPf1Gg5
0Zv3XhWyfz38DT30msR18GY9nT8X+Z9Rnk1AyDxqjVyw3t7OpuWdsXGkzFdUXG9r
2XCdPZ/JZjqOoCBMy3z7tagyvaSlebU6Z4JSxJC1PfEL8x7BGJiqHHnOoTMjKB9a
RW90i0E95KEmmMHJidkwg4OAkKsk0abCs7YNw7JyrZEo+SQYK8u0RjQX0Hde4Bxs
C6u54KWEQL4GPMYatbT9cvlBbOtTGV4NdWnMwByj+tQtluT1owqIlmBm/f8twn0X
rJcVSgOo38afn0Ukfuu0pXIEYzm00gwPuFwxqPmYLJBnLWS2ZFAZx/U7G/KEXjvF
QMTI3oxoiQxSZc3SQrMqORM5N1CUKDliGXVlTMK0GVAY+jxyfJCMcEb2t3/H4ilr
26iN21zXgJbgFMNYtibnOGMu1Olz2VOBWaJGFTTnrbZqopcOBSwty/XI9nBhIc9w
5TCsLEiZSvcBpUFM+cecl3nxXtaVv/l8xcCvWQXt5V0acOrY0HTQRpEtakeZrHwN
kvrUF+s1X8FDs1iJJgOw452qyCmyPV8sjCJmmLBR1hKhq7oVyEpKgs+ZoZRUzege
9G+ZAv6JgYgvRoULMKqiS43/BjyfizQTldsRGSdYZ82UnSEHiiJ97XaK/o+MXB/N
CZwk4FgnlNmQqBDs2+PCesmi9T33jARvZSgkNar0Fw0MVIPEPYP+WgnwaX7DJO45
MRJVe2D3XctuBY247wcBaPGSzhWGiZrparO62tn6+wGt42cqpnzy+8zPZ+dBXbqs
tdUlY2TkImq7u01gOelXYiZNKytARiOhHKPEP7KvaGYGXl6kYVbktWNIQE4liroK
otSFtMdlqUZxTrXURJRtqFGTttZ16yTbw83ihhYNgxaTaxkRsomco93tBqD18IOm
9w9P7xVWAr0v7LKRrn1zRd47gDuaQztbHouYb28ONj2defFNnRy51wau7RxqGa/0
PBjzoV7ZmNqbvY3kwsve/t0DiAgnezfNyL4kxJRBIA6DNpJbV7tbFxwF37SfD8Fk
Dj85rmaht7rl+GobTlypKyHRi9lsjFkFQqFyCyBI42/2MT+Wi+6vACa2iwl1LEnJ
flIVXcYtjT+uPN5p6BJksn+Ki+BNLnA7EykoPI9SF46bri8O5tliEN3SravFQTb6
8rH7qKz/KUqmzNIb8ntBV9VjslMqtGlH1KTuG86bJM2Izpvq8rlkBmoSbvGMXCO5
k+Db/Eu4oPOnJXBAWhVBv27LE2EFjzQWaUT2CJWw4lK556ep/26Vmy8ZzkoF1VOg
dwJh02TKtAQjlLYq9i47j6yIF9xhfvc5x/TemLwshK3peMuOifjpxGPXRqe7mweR
vu9Z83RPZ6La4gRBKnHzbkfTeVFSZ3cx+msV/e9zTYvduygsZ8boAWRwLIKhEt41
MxqqFQqJODm34fkP8D5gdIq4kJZd2T8qRmGdTyiChv30t06du2npGCOfiBmy9qN+
qsfHtfiENiiBkW0YwA29i01xxiRb+Go5a3591/3SK/iIlU4w9HsH7W1SKlrxuG80
afAJoM+0+31VQIL4ckn/wTmKgGXvUCK/2GumIoQok7iX/1aA3vmzKLhv7aVuydpU
UjSuwLCa7Ub2pMcoN1TcK7c+tau7/QeSM8K197ZZvLBptEnMfUK63Hzdiv2s/Fou
XmtFYInApqdxk/N5hCTHl1RUVLZTqyuRMQFG2spxiJHjgEPiKtA0CydSetR86ZRP
hjWov1DmBtwJvLiSWPxwPW33up8kJlySaiFJ0FDCkvQ/ODWvRgOLuMziT/W2EV7u
Y7qAbh0oREEqBH1GCioZ3MDf8hnTa/CZk9c7yjSdQoLubTHGdv1Xm73ww64lkwLJ
BI8brvG5jlGLC4/n2i92PNGi7f1Ui1X1E0aHzjhzz+k5s4StBHDy62JM5+X2sCv7
6Vb00c3quUJfHIEskfMkw4hlEBm15s7vmZFHHu2Nv0DsDKgzTiZPMz5qnckEhhmc
BImXlPAjWnA3lw7pdDziD+kKajGKWbXMoa2W7lnCnsBPGDefCjfDallWh3MUbo5z
JNRX83Gev/zxtX9lp5/Y+0astuXvYL4nURTr3C0fI4mCRY1MLkdsl335glxaT1kn
GZhBHKABlFunyIp5efDYcBP0Ap7ZDfwORksaMZgy5QTqwJLLzk/QAZ+udMXyG9Zx
4owINExpqgWdTU/aa8N7P264z7VHlrTqIu5Y4jGjVjJ1Nbk2FldwackcJtiJgMC2
/H+8jwFrWS5ymVrjgxWAzuxVMnO+AUNasEEP6jQ3b+MFZ66VGwophl6gZhRJ9CYE
IOFJPIUaWujNPiy3eReYekr/LF2K9pI3oLKA2ZZRfkHU7unrtHODM8WmEpph/KAp
5TTa62p9/RuruXO80yPwY33FJTiVZtruac8UIJlR06dKxn/imKsARZUNeOcFvrHZ
XG4ivz4soQsQdoVUSb94lUK3taCApJiO7Dd+X35uhQSFWoLv9W3BgkncAWpI7zU9
p2tGELDvwRHUUAc2Eo6fVszr3v7Ql7Uw0w6oz6XKf+EJuTT6OhEjrFJOKgj48aV7
9Ofe/2DwxRcoHEEnsVHgQw7gjzv8ph/C0EGTKqF01AqK2VwNfseNZ8DdrGd+qnHT
1J9Xuja+tZifMM7y+xUfDfYIK5A2SsEZWtuD/jARaO591I9jJpIW43np7Ft+psDN
51aXFSNfFkt8fOPBZlCyrMpTNfyJqSvwfIGFbAmIagim8/UXz8LD6lCNoF8pErJO
Ob0hNdoIUHSWzV9Hnpfxb3BE9SXx9tOEPaYX3qVVXNNx8hizEUHp0ykb+T6AZzsi
I4Wx2qr9eBJzfMIoipDUAMXQrjm8QByOLdBzkZHwJS7DYGlp977lC7llzQqW+Mau
o4Cl0LKIzYs9lsvVh2l5INNkq541ei5Ev1NDtawCMz+2IGTSIcC61t/FY3ekKSkW
6ePQz4AQxH/lIOU2QrhCMC4hahxxq0DGoPDI3PBbzS+Ncns5OncFjy6udeYmL8FS
Bf+xuWjLwO4oIuhj5X5wOEYWU3UrKhsLUoQxhdpJ9U3mINjnGFUTQhSx93c4iG5w
qq3U5Z9xvSkw6hcstxQgJ67TCGYOHr6z3rEVGPfaCJtNX8FpQCidWqdpGFV1u8IV
OatmGTpqgoXfCHQAn7mptAK5+HsZLTUmzeJQSvqgDbim8biX3jwXVasAKgDXENOp
rkB09ZczsfzNP+1DB5Kl+SUcoQLKKLsu7IVKskHkEeeCProCBglMVgZ0UEzWhtV+
wrVfAIF9X4jsyoioY8LXkNfJMpQqAQtHks3HpOeCF0azmreq0tFNmUzt4HVKOc4z
/CXEj/ZeVxSnYcJalnArfCCXPluzk+HnPcUlDvAYaZB1XUNS+oOA9ni/r7mNFyAE
E9cen9+qcedxgGICIXhdBMaOuvVeanlL3UtRE/rcMWYHGlqpJluOCt1XA3bw41F+
+xagQIc2xtkrGT1M2oKnsaDxKrNvd5WWlLsMdkg/e/HBR1Y4rYe5ZJHoUEF3lG/I
zDeLAxZKrGCPYbmiNHsm9nXUu8DK8/BKMBig7CkK8WBcVP6RNeP5OMVxKRm4amiz
NTxMc3R7NCKEI9O+dXZG0YlSDOwrZjQn4SD2Fhm3nx6RmVTVg0I9wlPaA/LsqftM
geQA1rUfayGV5hmQAmtuJAUcQt+ye03sZMsS0qAEoGn9uiWd1T5W5KSHJVDTNKEa
2AfU0JoKXLkM9kfYxHAytheEls3u8sKXkUGsmh7lrP+unweegB66sO09HTYgzzMF
brJVDXf+q0MC53J/JSkvjRjIwKTuVJelKCZ5fmTWZFOKg3JAdqSsvHTrQiT5gROl
DPizdv8DJplgF0I45Fbf49qByE86FypyS1+TJ/JfNZ2eqglha4u3BihNUbvqhtHT
4SegOIVXUbSUOUmuSpbA3j39ByeO0EZsnZlecGFVqtxbBbsDWUgEJwQDyAr3AkVJ
xlsCpMgGBtU+vnOxtc0lf0PjO+YAQ/StaHOb4ZfvayhzvfTCVlv3a82j8nCHcsBR
CGR2JHNt3jPp46SYd6OQiwixfXuNYiiTjy+copgEVSb05t5Kis2/7AMi1n1PaS5k
TG8dqmhYi+HH7UDALuV2U3s6wnANiDGsr/VRW1vcEQBLORXlYDUrKHrFnpDoVz0+
4Ddm4tduYtlMuecuMJ17D37g/MCgkiXI/gdOkqWsfMuwC6pD9P5TiZJ3tFon11J5
jbYutYUdhkd558tfek075+gIUVa/HU/Y2uZ1q5m4jd2E1jsXouFavJoPmhj5+sJT
8fc/CboKzXrKFD1OiCEk4CRD1yVrqEgqHIJfdA+GSoRc888DPBaLBGWSiXzb30k1
SfJBGC6yYqQ/GWOipUsErSbgQJgsf2JFjTFjJTPtMlBXvVC+ug+y4l5YgZrKG1ib
UeCQ843JvCzQPLRnZ3M54hhTXCRlIk3CF55myLkLk3LmrN3x+MoVf9PqY2KRNAMu
HqjzPEwI6Yvb5LfxCSFAh6CBSfLVq9U02pJH+ksy12tzoIroC9GSUuwV1Pg2Uccs
+mKkE5Foc1DMfGqgXpHYU+AaaETgcpWUIR0HVICH9FEJ/wNA5MRiYY4pvIe7TkXJ
c2OpVRE8x8AmOaROheSFrOeR+JitbpPZ/RDA4G0WPtd35q6eyeKBasJjlvUKkgzw
Bxv7P4S6oUOc8E3AVvt4rlYI2j+XovSgTP1dzq4v0c9WiNu1X0mA6l9mJtZhhZuh
nmz2nB0BKB3CrQZG3meVhJrGqdF7bE8VWQKnm8OWyuS48Q6SXrBqfm7adryXiSWy
ZaE1aBFtm6a+ycKKDF3ACGDXxZxS/CBVa/JaGr/+h5MMklRy5xujbuflbDo71EJN
AAnlztyBUEeyfYNBYyIvCnc9BrU6hO4uL5BXdTHri0CI/gdogNl3co8lQ4Zq1PGM
nYuysIOlqiWvCbUqY0jA/ip5tQgKG9ti0kwy3dzxAvKyhVT6hctJaT5OrEtPe3lU
nuvBrwt3b4ePU5C45VjZVVoolG+L2/06zvw8vUfvONnC6JmfUGxZlLPhKjY0j+RF
Ewuh5v8vW+TigEI0zCcb4ZM69NVjP0hTseQT/a+t0HiYvUkWJd77wKu5DMPVwxCP
8eA+tOOfEggixnXNY3YWgbW0TzStRUywDyNUoubCQDA+TGHvhMwLZEcInBJUkTuq
4SJ1B/duyuXHViBBWXBiB9z6NnjHED+Ysm94+5korz493Pjofa+M+Cn5X0aQTsEq
Q09/D2ptY7GUqYRFZk7agZlDvLrSWfxX+Lv9pkUTMrTXI28TNEeJp4gHi+gN+tJV
aZXzhfGTYm/hy7YorMdgQsnmtqtzihotdTEdeWWQB8Zq/P1Ec+oSoMz55m5HS8Zt
VJIoVf62+fu+HPzlfXpfjtFZET3cfrJhAPTU9nQU/JxQpbQZuYh4JStr2Qsycz3i
0STbf0W9RK9CVcEOwFaBS2kz05TyRy9vL6yOqNDKsnK6+QVYC9bzLvZr/IiNgUku
BcSCVRAFhlH9ACo5ES+4Q6lwYfOtc0suC3e4JEJrC50YEP8KoYn/kpLV7FlVpyPw
EexFU0w8YhkMeCcy8XBbETM9i82N27liQnpidLZE8hFmEPSxnPcmR+SDcAqsV/qb
Ycmm6vx3ZJMXC/cmVhuyYQqWwZ8GLcxICoQ3WxjZP+I3EI7Pw7QmI0xpncHnnizj
N2ZfVfvjpPnWck9yV9C0h4hhuix5K2UtxQGXao4ZU0VDGEnoSmvYKbl8GEm8YcWn
yW8rDZEOU7NWyhfMec2+Npa5ZuvmKKOvbb490a+PH2VcpmU5ANeVBhdSsJHXoHpW
qqcUIfbH8JVGEAF7GrD4Q39KdhijTEEmL5NmAvMLSsWHp0sSjw2V6jZpMPKhfNh7
0SA/CdNdPhhGbDB4ALxXYGm4Ia1BnfpH2nkL+uzqzvgINgMLEcI56Ce7JTG+w8gm
jasKn3NSVesko2bbBgzVsfsydl30WsKtM4LjAgslH0kbCmpTOG2P/4mJhlvb4k0G
JAcQn9faMfYRQGvWSVIw55R1S+ssnayq8OmAOBK5SkFhJu9461Xg7mXOuzayWYUl
+nmDX7UpUW8vB89ACE4/b81SDepxMXV8qg/KyyS4wdSmfhfhkjwdwuFb2uvert4X
xi6pLV48m1g666pU8m++mSzTiyHhW+GO3/gw++7v34XHK44Vm7DONncvKgpylPg2
0ef3lARvpPT9LSS063jxWI5lo/QxAdJCeiA3UA1F56tHd5dm4P4d9YP4Dk048ZqQ
lQ3Ehf9aRKrupsV0YJ5EeBL3eGKzOfq6fei4rwN8VtoYK5ZYizotTNFKx0bQAEYx
oNbRXj4nrCE0mPGv6Q9trSFWP1CF5qPZeiVQtIrOgQ15Cu3HxAOlINJBQrVFQiyW
i7/haIv8ZtRyrlPc3UO2pMTL1xYvwZAEY7RmVd5Ti1GBxBlpiwEYLMYpTUB6J8hs
AE4+fcCybo380p0KiqkW5GQdX6urnpXCQ1RXgVp13yETUfVHLHLU0mcQ1DXQSr9x
kSkz9Y35L/fSnAkZU78hJTnb1OtwyOPwENtGpYiG6HC6WWJ6TeWdOBfH4lOkaL/0
tCbsH13nucszVFJOUkW0m9vj3X8MeTT/q8jqaOP/0g4aTQMZDe/tqWZS3UagIe6/
70OvT5OYyWRojMEdc2VLXgZfLPylcqgM0yfE9Hf5XmO0zdUAQyKBi4QJ2l2EGZSf
pCjuoc7ojGJq5aHDlacs1a/O0FzjYJpI8+smEFk3tqEpmF8zkPOoqr5m8x5drtu1
wTRtbtxFHodOyNo20rNObjpEa6c5DDbOU+2RHQVakg5t3jhD4197cO9ju95cv8OZ
zhrFfQc+g8wxZNHtiBLMPYkBsJnYaLiuNf1pQdIoiBQPG+x8ccN1QqtKmQy0v+Cs
FkEGY8AHJepY5XrlfSCK9zFrkfQhmhud4gnI1n86dkdHjgDFKH2iuvWqEplpymY+
ovbovqme0qBQVQJKliMhgsYQuJjgaUyBB8iT62B/rYfpU6NfJmzTD4youefbJdmi
Ig+YyqL1ax67XQmQS+PZl88ksmfyTQmdn9op+2mrRx1i0w1L0tIKTKdC+sfstVp1
LHKDzBK7c1G52Al7I8WzBclAGJqwe0lCn5fJufHmeKwiBsRdxvTYS+yX6fDooY65
S/HI1vw3WK26MtB6HDZuZK1oqeYu9fof3WRKE5HQ3rQBw18/Z0Zlm83DcFhvNZ0t
dDU/q6ag0t0o3/hE8RMBOEd2mPE3/zf1i/X4tb0LEGhsDcB1BWNa9ru9RtcY4yTW
qcbyzavQQyvwpRFTYPEfzi95Kadi+tymdNTpCkcGT+wtP5jTT7ZEgSHuKOzzNaQ5
fXY12cDpze+3jHa4bMNI1yx/T4EXAaCw08ZB47qNQM4d53A8DcShQkaucXv+bVeJ
wsSzJuWUHQl1FNg5mTV635WW2qSdIbKDXwAUAVDaueBnb73VkZUfEW8+q9XCf9MP
amnPII6UyuskrHjcDVybIKVMRtekqgmX9bnBZDj1Spf204oFTBopgA+BUemwfeku
q2rYKUw9FEl2NhK4jegJYY68YPrBj2CJa8yX13cFdLMDyvI+fq2Aq6H65cvrTXh9
t7ZAltUc9TVnhGYVbMcbUzoX3Q0MMsbbUA0dAQ+lxuo0/r/7KTg6iC6UlADCyMp8
TzHZ+8oIKdF9HynJxmpLR1kVD9KCH+4cU/zSNLT9PmbdJpOBYa3PyrJyBGuUtCvU
naaeVPlciiDZ3i11KQU1zWz0iU3Snbt5iGN3x9rC9RoxhmGJ4AGMNhxHUoKf3/Vn
cRZBGpsYc1Y1zMrnRfhM25cpXT1/7Vxd8BwX4CpNZ7Vh6G+7xkA8ECy6TUNQKl9M
Mfiw4FhEXS+B7R4ZIzW88AWSISSimiCTewf9jHiRL43/QZeKAJdZ4XmfgIkh/gTt
nHpdmyTf0Vn5roYe+EwvkMz6DBZ/7xskwfuLYt1ApopcFko1uhq2pK5o2FDLAITs
edrecy/oNY7vhCSKT9NS1EKWmhnLosYNrf0BIp9gDa/SL6xwXxQYmRSZ96O4tHwu
GvuO/y+TcssO5NugkVDew1+VH1RMUQ+nMJVRS4vUwr3snOSOPHniFOcooJFtPrKY
MzHKp6aJkGgVG2BsqECBOobPaVIq00rVy8oo1AM/taoOQmnMHN8Y9/l3NtpMvDTa
4WLQp+keSqlOrx5TkebJiTyHW2xozBTobR9A1VBJC6KwYCxfIHc19TOb9ySaF0vO
0qrh4mGwOCTDubUnRMWoeQW9BAPtASQGJWmgFTA92o7n7knqN3xNApELz7uXnXzk
3JOOwLq5d17LGgYa8XPQk6YC18qRBlcQ6V30hj5/YCTCeq/WJC1FqsP1vt6xjZnp
P0f2NFO/3NTaf9CUUf4w+wcjYjHvQpEbrG4A/Q8iTsF1coC6SngSCJWY0pPGAlRa
boXdZjHAYFsRhGiKVZVWB7t2pEtUOLzqD4cehRIEbBmnNNp1GcKzG6JDrP9R/73V
HP17H0MWxt0U3/DhyUxedSs4Qa5PpvAKi+29EqxNUidDODeFDIFd0NCNrZ1omeBl
YBzMgF/PvTXH3+tf7WTex7lf9ypsF5A/Px1VaLXONkY0d/np4zPSRBifHlAH92sE
taKLkppixzH09nXRykvjk+MzQ6SYfJlDX6W4Xix2vZdjgFH9tryjxo+mVj9fIhSZ
Pq0nLA52yCT33H5PbqRbzRde+XQQmD8qWLhKZtOcpOsMT1xpYO4s6Cn10LzsAb/j
Nao5BPGzXIvgpBMGjjo8v4zv7OTCLk7BAEmqy0+AQXX2Gj9a7SWj8BHGFMv/T/3T
ZeR3FyDF+pr1XJmAzS2wH1RWvIbinuG2g3j4WPjWkI4ZrUhVZgKe1MLZPROWvtVH
WLqBBLUPNQvssn3HeJtaMiixkRX2w3j/EaLvtb+ibUuaCVccVnfVWuuTktRdlxkl
/u2zzG/QWAa/m9ObyW/doDLOzzPZkvmh45PbCcYT1DfspF+cYQHTJz0IifZZqaw8
goXgaUC/XwkCNfns/oe+c/ZcI/NtWATDLqTiDsbr39k+4Q0ZDi7Ckluwuv3pE5bD
AWCwFOQjx+IDursBbD53mmltbsSqMTh9mjCNwstE/cqLGyZJxJbHquAm6xB6J4KI
r20JYNRNnyZh1HkcdxNY+0RkJ9II3N471fbWLg41W7zym1nqHioO7w7AiPciApDN
QShtKcpM/P02wHf/Ml+IddiOoe7Za+2oiOiIIdTqaQEIiQB8fu7kOMFet1w0uZ0M
eUxiMeWYU71JVeUoB1ARpHKcMHgcKNsoi4qRAX55ZHoNcnzxh1utWLuVWhb3zdfq
9cP1ZONAI3SotsBKz9aHhLZ6xHk9fFnVxVrIxs7dNNj1whS8waqALLH328sGfof/
kxA72OZJ0iwGvnS92IRLvzRGMNoupaRU0rIKUf0rG7/ScAsGlEgWymZR/6lJ59+P
Y2kkfhph3PqfBtmy9IT6Hp+92sroSHHDDVsOCVNSLLUrRSeVA0wYrk79JIOo1DGQ
crQNlTKW/mwNmJ3xHaR3fBHvh6E1zXLv3qyha/owFCZ1CM/s1NzAdEgyD++6syxD
as1kJyc5a2O2gvytBpLscUFF+RYutBRVRjSHf4w2G9WSZ5gCg862j8q7HKbDPvIj
WM0NAqu49aaQ1uxKUrEgIC5lCuJSSXhHe2rIeJru1rFCKTdqARHpvJAVzT8vkuzY
RLvgENUGd5Vvy+Jrs2xJVHKUi/VZV334o1hycL6ah+VXWb2LgLWoe64jRkU1Wc9l
nZTD0v0UrY19KOcSsiC/zhwN9IHPIZIGTWGijrDhH1r2NWakD5MnqwOyLDOBAdxQ
1ziIsb/H4L59JY2rRwNLUroutdPVS6EKUJX5Iq6/q4+xgyxoJ3cFhr3+ZoEydS46
PyaSw+9s3eFSXSNZD0m5NsIUHT2fwGkiADOn13wiXO2jqFwcVifbBWu5+aqTJKJ+
8XvQrp7/4qKJ4ETeFvv4oDAMDfbn5svfCgJlHWUPAwmPHsDhWxX0JcZKIoF0XJyS
CAzVGtdlm3wGnnBc+GiYwJYpcVHHoH4qYZMe80OT2aoe9odgudGW6kig2VxTCLB6
ojDHuPvu/T+J1lDBSWcdOR31dp5nIrFBWTnKcI3n7kydv6LsPQEvVE0PT2DX6yGx
Hg1StReNetPvDlrMbi6uHvQeWKE0XSfYB2lC/PrprCpUpwcN7u83PdQPobn9Rd9U
qh5eDdqaf24OFh4g9NWTcBXolCD+pVXbw7RNjksYscQxKesATqzaRGgMRNYfdh4e
eZc7ZvVKfVS5R//Obz0vlHDTTfjacM6fkh2YIYS6hxsOq8uHitH2K6lsoCTwtsfI
KZXY84ky3DU2/fkx/1iQbJ8zwhepz8mFm1asXL+pz+SE1WR0KhG3BwiOy2dsKe7V
IRXH/+LhGOzEKM66wf+QQMxfr2IYyHItukFkGFmSqJOzHVvF8Z7qR/+EkBNFnG1A
pDHPvJGxb2jOOZCr0j3+MJsr4YbnhgW9sVRRNuYrMO4iLFRH306cMaFqfZ/tEEGm
k29B8OrnOzAfijeZAYGM9vNq+nZdnFQUCQaSmmzAm3eo+UDNqxpWm51xFd0rhZq1
QK3r++FCrHiC/pKPKznY1AunHTpiE1F4PzKqIjq1hIWfdEJThEQ52bVaCZHwXjOK
1mmEr/yhtLEXNr5RJjfgVHz6eDTj/kCaqVjOFEcho2P7aiXrCvOae6FqxQbV+MIY
biOmDxY0wmlU+85zKXDx1qc72IMLVDKCGPdy6ZR41bshChdzGyQpIED2DdorLH3b
bh9T7lDJAbdTxH9fqeaibu9lqNjvVK2Z9bt9CqI63nZfGMc5W9wl057iWl2+BkA1
m20vMSFGbNgsrEVN24U3HHrK+p5roy9OjZc1/O4F3+JUgTfk3Iw2lrqw7HF5qaMc
+hgozl0wfk3Rp2eXbJoIxZnAtiGuEoZnRSIhef6HzlMSH1256ON+RE0e4qYtNsyN
Jk7ACvPYia+ccu8Nq995uofbfOL82LLhNrfy7HyMr5yqzkPG143uHr5eR8NwsMs7
FmO72TYZLT+tC7TRHuIfzjfMgBLuyKJ1pqyaLHpQFz9jkcyQPz1TwjKHdWcuLDXK
5E6XDpMXiS38zxwFzuzB39LawuHYa3EwfizstmXoZEnOrdDWkzvtBvS/ILmbbQtc
6ZYORgmUPQSGBiL+8KsWUc1K87WMhFT8I2sBeuYmm0hg9Ha/+lnb+fABrRBd33a0
bVWz6wo7l21hm4s3ptkB7dWy/eRWDHb1KADDtGbqg5HOcSZChcxNt2nYebUIiVNl
TcouivcAEAG5DSkeA5b63i4s7dOuzb90joMgR8U7hhbUdm72dULaYJvH77UKDUUe
0Z7dyOivkLaoyj+I3is6cK6SoyiJLA9lv9OA9bT8vdQKHoXc2TepNz47alWI/gIy
oUYdDTvDo2ip+fa1rZp+DjsIDfbOV042ygeEjzRlaYs1w+ojmpuz8dZtHGANhQQK
mNzLjUarS1cSL3VH0mC/FXlZwUnRZGdnOg/v2oEjVD9YOXyG0+TycQOaMgFwTNhl
1yKkmvDThU4S0j/LQsw7dTYdSXqm4U+PTZmPin/17rMw5QFpJjWu5iiHdEbkwRJ2
AA/HhHs7fzF35QVhq0FbR6VhCoUlK7uazAhu2mUip5THvfpyy7HQxMtdadh6XlSv
MNw4OhqFtwHx6/uPzEPHVBFJiy3XJq7Axd7Sdn8vRLdXUGeYGaYLYfKuY05fgfv6
izo1z8/1C0jjDbOn+0zNcTYgkau46h7zR7a/vABdq5uU8wRebpFQWlL8frNpig+M
C5vxno+yq38WVkux3qDkR6QfA4WL0aRR8mupH2XGg1wI8j5yIukHBdCiOxr1jQr/
u5FeZshfvXRTh57LZiJW12KOWsFGhmIS4IiPzxhf66LZ5jzl8jqXYQIo+qp242Iu
mk8cwhRbGy1D+rQv/QjT7bT72HttCFIIIi8bajcjv+vCRqw/J4Z3sK4vnxp/VEVn
bmXM0A45afc0POSqlz5WcrODT3JgKxTsI4QnhalG/Z7Et3ZpExp/yDf28s0ncQmC
RQj4AuriCoGSyC+ZdQ4DV518KZLjKNW1w0dgFKaYU0nVxXZKIgPxA2eCtYoisIsJ
4FkfhJZis77ls7kOFDyyKKy0uFdQRf00Yu436w8oRU3n0QfvPBXTBduKbNodZxrg
uq8ejsRn5L8FoXDSIvVirQ5Jt/WlfgvX/udbVXBc2Fgx3YgyHv1F8C/zsAYo39iF
gcyF0ypoI/dYQU1HYIc0lsZ99G4PvOyIHdyKm9HDymQYh9HQqiu3gSDCD0k2+GvS
QTTOg9ZG486EnA42dUQ+WXxqK+mAki2R/tzNQsawC/RYis+B6ObzvgsL2FrPH1NP
eaK29G4g5rCNe/bhHmg7q/ercgkQRmFuGMo3EH9YefYwZLusNMSNmGIhve1gJcFV
TIqSc4DxdxcQMhCbvLoyerg6MhAO30iLc8SD6Cpb39A6fpu6fKFh0mSw2sDIaRAS
igXFRfpKWYNCIUAVn07OraK9oVdys8Hl+L+CNuBLXnNgJnEFoxCABwR7EY74LNTl
vfYdhlQmoV83p13DnkIj5qmq8yw/OS1qwIs36xn7Yv+n8qN87w5mcvlmvupADP/P
CUaqDcYRK9Ph3iDjlT2+Jp1/2L8uZYe+YVOEsNi0n4y3W+8G4yVxIoUbhdTX9RTD
ESqmUTqecs4wsw8CnOgxhZFxa7E6IJzXm9XoL+BE2YnYIgX7wCTCOFPbNdDJ7rip
J1gwJ8JPD+v49RK3l/ui6JjBsaTfwHdMC4rR9kJRY7s/FjL9BEGnMyw7W3Q92uI9
FEwvUpIfos5VZ0Ol7x408hRugao7ijsavg0/F/i9LDnqecquxlgFdrNgSNeg2tqo
6Wd7UvD+98C46SSVnEy4Vx1qcaBze1QivrHiEB8fzaV7MmfL4ZBpgTm5ob8//3yd
QRGOSCuN6YDo2X7gExMCnFCcnzt0IRQy+i1/nS0w9yBTkoLpefIj9CJjO8Ql5xTJ
sDfjXeAtljvS7KEnP8VVlcWq6c5f2RUkP8WoXcPtjGsnwxmnuED6/uV0NC6gpkUF
ccwOFN4t5/AaRR4eA2JkV8uxaBXC/BuURx94MsUqNLdJeedy3m3Puzx2n0ttR2RS
5ldgYYtPRSI9QidH8ulTqjo8Mi9J8fUeyP3PNqQGrVOQb+ylciNUZgsfc/EV6fdq
iE5mBZTNjX7U0yZKZ4SF9jNsOvs47KlUJDEFXAgOhKCGiNE7HCvsAgGtI+bxldvt
2Y4PoscW9csdEl0ZeSPAFUsMkRdIGzt9Vkw2tNm0Afj+P0ijgLittceb4aQj0EuZ
tDv2Pz2Gv+NkV/DcCIiokr9s6dZ0t7xl97wwlxlhBooMVvQhap2IEpTnTW/14iyS
LL6q+/8/6D5LX4VWmtUG7ou8iwMLXzJM9JKckBa0hTpFLquncndf+vXD5gNUAJdr
NkIpZbzFq7YWKzO09iOB9VRXPF3BeQSnIP+mef9FSYb81jb62w99O96IdFuEGe3m
S19ca1Rqyq0fjSvt+emdgkz/ahIoWiwH2MwsEMjZrDFr8IyI/MCqt8tgm9KhoVtj
+jN6IQV6sNph8doJ1/W+3qIle/oCIIIQRkGoJK3V8bSMyiEoMVxwnCcEEABfM0bY
M8f3eRY8dj16ONByffp1QuQMNUCE4CJOaj7ongIEMmJK40tZ0cV5AagORsHMqejD
ijhngZGsL3rK4KtzNKN5hKCVD1tFutyBywgNkJ6QZ+LD7EwT5ucYjMyrqvIZcbbg
YnvHtHS0X/32wh1X0GP7j6LOqhELtnUxVTbIVu0dWtDbmntdoViOa0gVGY1mjzos
2XKUOqeABMLoRfQLNvotiHVGlsnpmdohGNmdrvZObMgs7/KpsApmmgpn5MptgQ8q
SFdZx8oqrPzdFf1DNJZBOeNkBciCp0JVV6tzCGGQNh5ccbWHHlKQQw+mLfPhSqoA
bbd0UXhKYy8zyLnkSokMNzzSN8awNtywzay5K3Ns+ocMbC13Zhv0lo+cVUN+C3xb
Q1e4yY4JQDRci3LUWYv6ory1QxujPaTR4xUE32oLCzFRHD5xZJfYWyKZ5Oq/8W+2
95Auv5Hmb88f1WqNpl1uLaw51fBF+j69Oy/wJirtFGH9EiTVAHvd78Ztx28pnJfF
uVHxPynO1spr3uqJUnDDSWJ+ZQHgQJa8EWSCAGiQ3btyTWwhkheCIf28N3kxiHwj
21Wai6F9e6l3jJTSPrPosh7skHo9p7zAgfQ4jgqb29HUugSYK9HbcpWlq4quug1Y
6IVOfDC11MrwAuVb+cbn1zT4KY5lLnWHH0/XGw6S9s4I8ctb6U04CFcUVa1Udp4E
9W2hmtY886I8FaTAVzLI478gU2jP3nu9kcLyozYpKj0TAfEqJXRlcS6KDpT6EyBz
NjZ/8Pn1fXmSb9fpnBtf1a84bWI4UvzheP+PXxsXsrI9AtXORv4ZNuDouuCJEqyL
4h+23kRastjkDf10b0EL3K1GTklz1/eItdReYNtMyFTpOucV7VNVkp8cAYmgYy29
naa0BOdepaBl+zFJr+VLDmdidNj4rN3Qsfe48Lo5lJT01jbxfVtqFikn5RGrXr2E
cHqLfbXdEN4skBWEGjT1NRaaBZwjNHaofU0+8+h6Lb+cHi2Z7vcRL78te8SDYUhb
ulH7CC0SA6iMKEYO4rdNCUlXdy5lBmH/8Ca15jvG8E+7D6P1QRrlj/E/SOsn48Ub
PhKZBwEb5RNx8pcXo9/nGWF32PhxH1SDS/HBw17d/XRCursoh6BlufrIjdP8LpM1
1qTuLzGktqA833mV2c7YT6dICQ+KXZFw+gs+hJJam6VY4V9NeqN2up3byogGkYHB
ayiFQ0bLhewOjAQ1UoF0M6/H3iz3n8vmIsDjAjsyTehnEwpx+oora2o+E1J/ZelY
fnQGCWkw91DJoCZ2uiOjJUprWufe/vE2Z9ek14vlsQEDSWmDJjWq9bma+NpPDNlx
Jpuv8w8e4eOhWBz8OSRDL4LOd8NJSp/t5Ov35eGLzx2ZnY4AKy2TSN+fak3nYGhd
vibAZEk0NxKGiCnRsVALP564u48fcbKwEFYIpKA0qBkksmtEfK23SeQXL5Q5qW/1
Ru/ORoqzKkTo8HqXgN/hXTZOuYl8QlBwi4nSpcMHmk7JIdHk7MssNXdqvZ+M+4X/
p38waaJ3LjPat2KKXXfVHbIDnV/anQODC5mVWbTxa9KVpLrCXzACku0sUWlJTQEI
mYUmZlh3Iq80SpTEY6kDA1saw1Lh3UYbiuU53DaAwuFFW7d3ftBMnHsDbqwSQFK+
6Y6hi9POuUI5UvE2KCuZoKxprNz6AUU2X0gUKSnFqRU3BHiJmw61wD2HO+1+I3iu
9TDlH9lYHdklPUtzYditUB/vxfGcc3mJ6zK/C9WL4OBHmNAgKIup/qDusPyPnG84
t5HwOW0t0Zu+4EhQePP0S+/Nw9U9LwNTuat7xoQVNGiu7p6n1znAa+qds8Mi8lsG
5RVIAz9Hg1c67wnvl07kwgcL1SIk5bfMOzmsCMsjiawKC3M7Fvl/b3UV2lB26JY1
xzqJwH43cV6hGiWazIDq7dRoRUIZ8HZyB2AyOJRLwgCzeAH0FoRsUPiKtQ+SWbXY
TAjXdLyCxvH8R8PRSk7RuDAmeEIlI4ryuTx7B6yB3bEbcTpLBLh/IlzLbzBgvQJi
Wu3CcFr0IJxVgciQSzOdz17lKk9ZD2dKC14qaZy6zYlxAmpp9x7eUCjSxqRec03z
tMpal+k9eaiM2iJEzI0XFTGWBRUEqDL2uhsHdIn5E3+m+UsEe1mzm0nxsC0xOstF
EdfT6BEukD2AHjKU2GnP1WSYyOG7bWQ8m1D1ZkYOjZKShZpbaoQeDy4DDtZDbTR5
SzUh0Mcw1uHZymLUEDmBYhvNTm7Yr9OfRfYT46WV+pc4+Hqeugx4IFzfB/rZkjEp
woO0aruVXV607O+Jwd53HAq8c8RtlL4awxLoJSItm9irjOPZZt7XNzx+UUGl8DqT
/Ch6dDNUjNAkA5fSK8+f8x3X/72YoanCMNy01rAxu9fVmJxV2S3BIZmtknsgT2BK
vpdKd3jCwWAn0spIrI91GUmRyn5sl+f5R8bMMpEDDyuniKuP2ZI6Th38ToN8Aayc
pVfhsRv7Ek02YjhZWxUchk9dkqzg7h+M/JXKcCbtu9TyL7TIWQMYAgaAXulzSvKO
Ycsv9VjOqPNdWZZK7bOwVFUNH7HbiuosvMmy/YVl00TdNyIAFn3zJP8H1s1jpb6q
1hqQRf/B28Bn3PeoGhLdFZh8xIJvXBqUpi+WtpZiY2lfp4wNbFISGCDaKU0wTg7V
hqYoZgp22ktKzEm3mzPzwxMISa6dovfCtJdY6Flm9BhfL1TuA344PXtgrqrIa2tW
wt+XCWe84aF9FlAdR+f+t/SZGzkPt5dUOvWadREqAICBYx9D6xEmKLCBJKVUMhnF
MCyCjmg1A6hKu3f+wXrIQyK7z5uT+lVz/DMnFk3s6DO9YoWCXjwm489M15F0hBBC
uDjlyCUQXeohXA628NDv1KbV4Q4almn4lVP6cKrOPFIEkhkBn8nqRpPn1zdmRD34
e/wJzUdLZQ856uqYUio5/buShgvoezm0n4MvR+Tr8Az2JTCz4azx9E6A7hfdY20y
5v208q1jgPEz1WFfJLsdFIzlCIA45Aq4OEqbUdQPgP9CaCNeDvFm8a3SZSUEK7QZ
Pby6hL+sfwViXQBHgq6LntvyWBzCUTAqMnlf68D1XHO0vb7y6QpYfQg8JaRXxYer
5EXggdrozOWm/q2XY8gxEDRoc/znodcyfma25C/n+qMC82/y6mXnSReZ1IX8XL8X
sO5jza5VQLmbxK8p/6WUm+2mAqRpNOBczQbWa071RFgYf8H3klfQKGychFojd9S7
ecPsoqi+xNZHgOyrTnJGZ9HsYZzBc2c3V75G16DuflYp4GaV+O6WK1/VijW7V3xF
9scPAxZgqNev0O4tNv7XACA/vV12DIrysSzjRhl++769TFiWA5UG65JK7Fzz0qql
3am9d0xEkBmH2x7PARGizBzmfuDWtPqQKL3TcAtvuIvGX38ciYih0Map2woLEMEe
THyTjJDgs1Iv/I+rw3mB4ehuZVTrZvcjAvAUS7biOLvKsZ50U1+MSdXrbh7VTnb2
y1b4s5geCj1DGuYeuX+dHzLLZQvGJfzycrP8KFjK8oRtZRAyuokMyKD5Tn6cU8Ps
FLJJF0Khn9Hkt0td2nKwAfzrlmoDQ46JCeIoNAN+mcrenHKewuc2/pQEy6Kk4J9O
rRFWEPbvelMsm1AVOIPk9ewXdx7e0faAFDIIQHODNaZYZznotF+wi8QweolHjkQT
R2+VQbJPYUNxy4nXL7ElFNA/KgvYR3fTalVH1laKnzA+aBvd3znOXVmxCB2kgj2Q
dvTi4cx3yOpE8t8pKjof6R+X8XCte3o6D6v9AgUAdGyIPoa6w6s8LAL1+iIFSZ4x
BHzIVJZFB4N3oLLpfzJzNwMcMMOySc6VFWFPX433OZ1i9zYc3uVjktN5ictZ62P/
Kasb7pf9HHN/ZL16X7HfPVLL0fP8kmMpv4+nA/lfXICGWzToF7flGnfTlECQFW0d
lcdCcSj8lvwiviF4wqvXZwNRghqjVsPFvBW8siALDA+wqKEEEOIYzQZQcD/m/hwk
XLpwtxZQiSFHJuon08WqMLmP1J/xu52l93rqGH+McHWaZlYQCYqVlDXAc3RRT6eJ
ixOiMP6mK0H44rSQwRe51KgADddQToOTXgBEJEM9hx3nF3TrYk46WwYW9DkYh36J
iZvkNUehicnbGmF8+yHJY/IEFK1HxnNrfUzLojRT75pAZRCKcwiYESrxilpzQOOQ
jfyBXxvbWXHSt0w1vip5UWlUmVyUjI3nrXJViTFeATc+aT49D5mCWFftKlPcenNi
w1GxNpjQX9t8HMMXi089/YSGX3a8XY7wutDDWi2z2JQqpSJxxwkViPnnIFQv3bim
pp/6b9szF3cLkXDRhWlcEUSYEtCz/vZyRMrAcySHfojAfuQ/tAY2xk6WrGY7liCd
G6IlD9O1873gCmnEr4ZINc8oN0a4CxZmIjd5pyD/f69H/5hM8PMRg57O6qmavjTf
oQQYySzOd0Z7V9Oe7WjGJHmC3gQrEwRH6aKOJFrvf27nF9f/6s9x12hjujX+NXSQ
O/81KkVffD059erbD4XHsBabp/FX+iCEI86sDEcLXYo/rcbrW2PxvutV4VvogVgH
kpkGWwMpUU/o/PtyDHZL5tA+jskJfsabiamOUL19gRMr7r9b52cSzUujX3EfJtqj
JDnb0q+ap8MqFIgf1dOL8Y3zquobCeHkUgr8x2mdH9Iy0u6BgLFzP/HcYQ/23v2W
1E3UCw3h2l3H60XUYIQ3ipznLzcq2XgIUQHZPXUSXfOFLEPvu7+ArtAsyNO5rf+H
YkGhHAaUauiuq+nMNdVEYDfSajWsH3oiHkisMzsKdriYAqcU/kGQZBTu0r0G1aJX
8H9kSVctUs5qzpfkb8BgfEAXQ3mYibDGZNrGAeO7K5tarBtgrTvEWh5s1Lk11v+B
x08wqqgEs0hcEuExlG3eeuqrWczV85YJm9hjvpxJnVL4WZ3vqNTcpwi8mtuHLZUB
+NKp69yesOSgRqZLHmLyLRzxlu+4IXtD/ahzucBLChb1L1I3P8JPdrD+m39cVVBr
Qr6m3ClJJxrGIelWu2vbl4IRNgU4Au/it3VQHKpt2DFhWym5axEY+u4D4A/0+Pyf
J/26lNUrj7IOGyW13i/RvQHSu2dvkg0tseNoo1EyQCu2fYROevY0XD85YNst2Lj6
a1rYrwWk/X/G0kw3nDx400EnkU26gLNf60Ha5xMIYfLR6B2ShFX/Q8qBs5tJa5Bu
SW9J8ZeibkiFcstUOtMZJ+CSgABKxj1f3D3zFsSIOYKH+wFW2Fsxa73LK92poIo8
Y8r/swflhNIAXAR3kahRvskNumfjbtib89AGN1A6Rlb6CyJwG8ST+OphzTEfIKoe
B8oyEOgO9ZZECcYWD1PAliB3ltDZO7c7DQG+UodyHyzs3fM1mmKWibARre+yaOi8
/6eTBMEPbNiWi5qQmD/KKz1wPOJeeEOxtpEM031nkvBESzYFrKkD+9NeIvWDBR6V
7byuI8TPyPz/lF1CSs+18dRKpH+0AL4AlP4MRYW8FWCc8/6CX1zcJRYsCRw//SgD
JaoQWW3mtNsY8fuF8f9JVg92TzifRAiojjPruLi4/r9PGJb+hLWU8WUevPfLjfjL
yCXPGnLD2KvNA6O7i/Qng12jwloZhBN27GfPT0mUtiFmVHLi0NOXpyu5bcRauknJ
xOSkcMpXrZWzp5ZBvDmDVmql432tRnGCahv23IfDAF4aojbmqoTs9alzujtnOGmM
FtN+cjkNGApr/pj7w3Y8mt2gGFO4s6TMqr6ugvN62TU+JANyHcWo3pMOv8pLx6U+
lHsOb7gIULo2qgFIykqKZ4gwQFo+u0UwqTn9m7pdx9JD1P41mylddDJ+YOT2XL2Q
kUIYUtCVm9rkaoor+YJWi8pTbm/f9xFqs3l+MQa8wHVHkNLV5KEbjYl7GSPBOqTG
NABQP2J0ltPyFdlcNChZtwhRQRo+rxTPNqofOlK9SMqfffzyxTQBt5y0OqHML5IJ
Sbn7DaTTwjrOJ6+NeHPFJXOSYwppShP5g7fU+5LUsJBQoX3XwGm9NPR1aEI2z2+G
5qobRu6dbWqX2fs+dUxj1eJQdyd5JbY+oMbSGJBI8L9eD4ySBkwYWay+oq9UnnJX
b5h2TcMiYHG7o9TRpmvrBgIG//ouW0KpDoH8Njbs6LXlbtY2p3AERmy2POJqSkKb
5GUlfu7ez+CNO3v7R09BGID8Xw7WmZXgP28MMUyzPFNnSyyEDQ91ps/t6tsRa/Pz
RXq6p5c58OnqyFVRnkdXhV9lpMdvnapwXhMevAonTiIYwZCj16bTrKf1vAhA9aqv
QSpftmfHSKRiyI0PARMytwqwp7HeVvC0ThfyCLgXt8OYjgxI7gRzZ+LczbDiDrI8
cYamXIlfGS7R2epv3WxJJ+NA8tok0GhzSOIdkaE36FfvHNDYXxqSQ4DIriuGC2io
Hu7D9Ew4KHbjfmA5VfAdMRe+MaGXXxBrpFIpYtZEQXKA8L4qS0mOOTMclYtCehpd
Zc8avQCrcseE60v0EBIGl3UI89tjPfq+DXhMrUPp8/7Vkdbx4cWMYp3+bH5yFy3n
QDO1DiSUJKBv/HTSetEsyUOzq8mVjwJvyWyBqLEwF4e/iTVXPsVXxLlkL2XYtpxM
rKEC3TuA84DMy4uFnLO8nEwv6SCLNFx6B7mVoeZ5SGmMPFzDZRjISA1soYJtzeEz
jy/JWz6O//eSYw35byfitKgT/oTFMVqNdjVlSyDMKQp+ewZHG7GnEqL4hSLxVnaM
AahI1SoWfoDlNmiPYdcXGwJX6TBAmBAKkaZr/IMaKPBK+IvYS0gbdXEq0w3eoTII
QA8QdNuzFJ6eEsJRPEjm/s5NXB9GFXtA0mhiFPdukQmSAxmi/H8GMneferkYr1lR
kBoOKDg+ZOwjiLW/DR5wC9fhPdIOcsYFqAxNYeLraBPBqOziuj8rNFPl5hbLXuSS
A1LFEV7Mh1AqCgH3K8qD6hQmFTF0vXZiEScBJMoQuihbgT4IjrcHdX+pbJi8iqbn
bHvZv23FoHgseUW2gAMen3DxF5dM9Gw4tKT87Xtv/4mig7G7x4qTLlSsCbn6MIHV
EvfevS9fpuyxFnJLNf8HYPHAHs3rMasmM47MQnBKIWeSANO1Qd0wpkK5S/scWLwZ
O7eHA1xjK+PzucAIJ8jv6Rj52pElnOykNYQS1Z0xA2asJKMWCpx9cgGVcrGdjxqV
oI1EJ4xayyxJZaZ2PkOTiNVNz5uFPshcXJ1NOZpMNgRZrBSMoJmJbZedGJOdrHZk
t9ZCmJ18cHYDKwq+XYCd9wlFajpznndwdUH7sRMI5IStS+dixW94GhAa+NG1JA1l
tFJ8SpCs3UwwekKuq2vH6nYzYMeiKf3HaGwmxBT4GxFdilCwodHvM+Z0ca009SSA
zwuJQPs5z2EYCQQFmLNV4eV2LRt85rkJ/su9ksDZUjb0uhVJeR5RDJBNAXUR633x
vVeRCLCx7wfSv9p5E8rcjtIH2mMQt3bUZxqNnvJZcxJ47teJn9DdNqng5aji/ghw
RDBksprBcwNxAjGvjdyCPFsz+k0Y6XXaja5EMcP250u11quNSaaPG6JCqVwOztjF
+RkgjKlnJQG9QA+VAw/LZIsjOEO23A/80gyGPmNxfsbkUvhLNKzcQDE5iThC4Tgb
ZQadKtYycW4XU+vu8ulIYHliZFRV3EFdXSAXmLjuomhLONSPY8hhGzZus99VEj6P
Uf7ObkwfRMS+cnD6mv0Jp9DT6kPQUzp84vCopoN0B2E5alNbeK9l1JW1TxXsjx26
L24AbrSWnWA6CAVlviYjAyGQhllZhSgI8hbGhj2UKLdXwQE7MUaZh813LqIy5E9V
Eb+77Pxgc8J+8HGb9oqwstkIRPG45dV600UAEIaG6rd5LZw0C2Vygw+TUSyhYhmB
yoCjGJgJMNFkPLnavJiUW88MK5K3Vi7oJrE9S1pUOE+KxmCjkA206A8d2lVSU9BN
twyFYAWcg7DJatjHEK8A2smMOIn0BhfaLIteiVQXswbpXuqwD1HwUgLuIFJqHPbg
wQ1Q+ymzfwJdE4g6F6WiDptyxclJRoZljIyi6TpcYrFnAJFHomQdy/Igou32sT1G
TnGh4QQkHzKVLJTDtplMx9s87d4cRNbpyP+jw6R4/BHjgstQRrGTCEMvKMWcr4a7
+j5ihw6IsnBis1/2Ir8BOxhUmIVMOvlv0T3Mh8Seok7uiZHxu3N6D3ninYGxXywv
Q+A56+gPd7iR0y7aGz5C2RBO16cS6QmeY2zOYE58ndwwlm6+mgHU9JUeqszx/G9b
xsOseBYW3VLnNcQcfNKgctFP1MHyRx4L7AatbX9QxHa6xeN8IIq0XLPdzNTSEoOV
JvAF+ihwKqMAAo1zAzL2Fo4puJ1ekK5xe4UUekqUUtBhhgKm2cusymXxAT5yViWl
zJ9rwP5Dyz2oXPbtSGAdHBkcUKgS3v95LONCxTOkf1UfHNXpVT/8sqopQL3TDskS
TxbceTdS3vZeXyfZhNI+fC9k18V6FygCMj5JQFIBtCTcvwhDll/WlsCGdMKgBwQE
cbklyR5wtuzbMQJCIFxtj4th9zjtAZYvPvIasE0eAlSQkmpOhBpeG2L19tZHsEJm
RAYhgryA8aXXc5r3n4uaZAe8HrukI4qQ4awtjnftTzcn1plZWIsePeIvCbPdX9q5
5di20WJRSC5JnA5A94EmB1Ku9LuVDAuoPz/mhuUMsJ5HGnt5L2jMof9MtKR8nAUN
6oLfXMkGSqwz1GhdGpnera8xBmCe5Tfj7xoXQFfAh4M6vxvlo+zYLWxGJXPjBRd0
wcmedOoNsbIxQaoeoonCaiRyDH9OzWc/6Oc5I6rdqdi5QluWz4BLSupk4aHfbjTZ
xlhJnMJyCR2i+JgUajp8d7IounzP9hOV8UwQyCCZKUINM5jeYys1Rt1Ia0zjmgyc
f3FtaP1bSs06m+LiQi3rPBcla9Sq+YMPe6NF4gF0htxKeBwxyCKmjdospR5TMkUM
C13s/sdtgvXcjiCls07uLbKKK3I2JW4+JxOnQ2rspDUJN5JzpwfHCPZfBtp/Wejh
fSolnxqwfO77PWg1SAUk7NfBOMabvlcMzNEowYPfvvLNeultyiLEfetCFlf2Q28U
E76hWj7XNEtOfHxjPVlz+MVElUzRPiV9CJqWdl42L0it+Cf9z6G+LOCrMuDX/zaZ
HQqx83S4Fd9BMeisEox9jLbjQOqEngb5vTcCXxBI6mgeXFayDT8tsdOsl0D1mhYu
/PRn8r9kCU8iEnNbCBgWv8qve8BFIMgQn4FtaEhtY6TTupKyBVpXZnLJmJblcPig
m7WJNfwNxH610p3CxmJJtBB0QXxdQipH1flS8AsK8xgb5cv9VD9pYEKhWCY4Uy/u
ttAsDv48EUUHoWU8FuNm41S7/JhfeSEE710Tk3OPYc6WASld39yOce29uGI691/m
ASaJSTZ1hEaF9ozUUD3DtbgP5XMRTfEMUg1BBAkOTowpS+Ou1B5UuA8KRTlZMlCr
ZZH7oPT7IQ5y2m5VKW2yjAxMh05Xh40g8DrHvR2IUqCyDonNR661JxAdhosS6VFm
m2+tDm+hpGDngci3Yjpkpu1LQ3nVhaRFuPBO0a7vJre+haLas4LoglHOAtRvudm3
wX/o1kLFXcmeJCnOI79DGtg4TkgJOtns8dg85HqUiigrVgWg+d7QzRJTS3v4MYCU
JbkSVnlaPALzoeUkdwpxNVnsc2aEyAV0qOQLNno+JOsqQvnUD0ncnpUh+Le+WTpW
KH9v5bnocesCLnUrufyPdhj0r14v3RCk6axlen8QfN9t5fgEb0KuUHF8pZk/b7TI
iN2HpIKZiTvbcKE3zUuM8bX2WXlVSOXBMQ4yh3vf5WVW+4iY2hUqwkQ/6rjzZYEJ
3X9K4kRAUiQ5kn6F/e4Gokb5AlyOqhGn/HKNZW3SwqasMoaFwtXhPIbeuiuF62W5
OKpW2mxyTkyAiB3TmkW5eav3f0c/ZPEwNOYlFJQWWHhIKklvXj/KZwAcaJBBc2i5
prGGboIna50gSPmUCCYbs5cu5UVQ6I6wtudXYlOIHadN+syHeCcrjA10kEy91BnY
OfQS+QtCvwWyRU9dx8ryIuve63K1FAyQbu3e675T/vsl57IhnL5rmGws6tTHS6Fo
I64uBw5zsotagqc2RXFoKN7ZjBXd0uizJQprrjx67BUuP1iuiDKjK5RVY3qL02xt
uuV2C9LsorZikfaKkgM9f/WFZyNCElGEb+M3PEroLwNk1ipiK1qqWjmW/DVN66zK
b0QwjEtkxqeuCdwLF9/31cU2GoKPXywi0QW/RMVHov+HK6UP2dJLk4rBS/f+Qunc
hbPwgTotgfiHyOEI1ASsR8JTrSxrDvlPgpbOPPEnKboUpM2DAIamJ8qyvMg1l/ub
DHImHH5+NLcH1Tuj3fvLKFPH+xIawKvEM6D4vrKOpFDGYxTsX9ZM66RvyiTYYRhc
Bfx6c2oBJV9DrXLNfQhMdtFn8NK77VyfgrnEUcvLcOSKONdmJ4ju06+4LFdBj/Uq
fKBrBWck3b2MxiBZqW3l59mg4SS39WKPRNmIDeqDo9Uo2+zTGp92um3T5dv+32Q/
7haYAStXFeQyadA3G9eE3H7kAeNouKps7KWZsikaEl5cc4LuOj4F1exaSKu6qHfN
evhTs1Zg6KQh4NoJm2ecDupiyd9zDlF4fuoza3StCVylmOFRQDpvU+o6/vQnKehp
hx9agSntsEKlDea8rtb7RGwYQlvEJ7fHsIPeD54nffEiYvAm8MX579pn8DSkud/f
AlNGXB0pyd0tRwFlpxU3IW6DbpzfS/50/X8ZtxnKxLc01l4iMtvjxMUZl/Mt3RXX
yaEh5gkAleNGewkhZgSRshDLHkOaiQ0bgNK5crKuUZ0CddBA4yJLPxqaQuUwRFmf
nGmIpdIr8lWKf/8TevL/ipyXzrHdGmDwYpPM/RAO0e3sTUGQ8TXFyaL2LuV1qt5y
wUnkdarmnl/Fly5UPLIe0SuE8XhIEnWAWQGmSJFe1b9WKzjJf/MN0vDKqNIL9ReJ
rxTbqSu+RLulNuY0s0jCK/VBDPfoAOQwUOvO5t01eWuP+INc0Q0Rk80BINaiv8UU
8NtWx8TJL5z44OZqpJfdnh8Y7kFTYp+eU9502EE3HOsipOcHFKGCkDWTh2MK4wLA
NxW1+1EX2pj0ZE/TBoyLZW8EJukZbX+NqsLQVawlqRjhi9rSC+u70m5JUSeD+sEb
MH8gr7bMKBTxXnbvJO9FgznamrG+mc0MQUmL1qZJ3foc1tEoboOYHe0vsziEgP2d
cyBI9f2QJUVgqumaHmatJkWDcC3nYQvh15GGZJD5kvhVt45bmSWcnSoKUzhuzB5+
5nJ1GpE/eLa+2YaDlyv17cCrsPn1m3q0id3w4GkvQQB4XHpF7KqmAmUxzciN+yij
K9CcGtohpgKFMdA7Sl/5OvP3BwbjUF0eM+SdV0OV9KXQdfwxlU6lFfhV3h1JJbZg
3l/V77ciF95m41unlnWJY/Y4ON7FtXI1fntXU9BSFh8nBTTUNmphYSYy2u3uf4tE
y8Z3Y2VUJJKlmvHkk1r1mUiOzygMp2VaV8vGIwb8RUkCE2/paYbPANk0ObZVtIa5
t3s6H2LR2o7vqwC3dQw1MrRJwiJU44fHTDOVWMsI0cEX3zlDoqs8wR2zAznLaILc
r0oCP6tvIIvh/nszlmFsTZI6Q5Ji18lxjCoDraKiDO8ZnvEl5XBwPYR1q6CVGglF
J582KVKJKofS1HVKPCy/jjtmCEAvckC8zguCa8KrP6cqW2jaCAPf0AYwhBAopsSP
PDcp1eM+gacs4+dl7R6Ey9GVunKj/WaYRX5o6vgCf4pso8iysUEay3xkiJA0BgJ0
22YcwGKrzsfJEVZLkxn8rtAaTtHt6meayRqAqH+lmlSyhzVtA3hh/pKH+P5KVF7+
54ZIdPnKDMBaBI95/crISCcKXqWFPXmmjcYoxMmwfQsOEUt/L7xNEy/FxHn6WxPj
sPZMFN+Y5f6+HyKzkI5vYOCIaAkYVLPhl788HjKI+oYuR96yv9leodYMXRCc1qC+
kKrBf2P3zscJrzFTwUDU4F7TxKDNebw0cqf6axmbDJMqHJD4vSJY921s2vyoakGA
zpuEZi90nq+7blA7l03nP4a/69bYVkiFrxrJuwIe1u7DTaEkpxdsYPLQFIgDbq9N
M7OquMeQetaDNDOOwAxFiPHTFKgQDsBUNeRlzpLHS6+WglqfBieHwNlss0pE1CGp
DGl102jmh/N5pJK+wWHgm62fMZ/nugbzx9AnEGxv//O+8PAl1nCxTatlQcmvr520
ZA34Tw9yPc+9l3b1Jv3LZPEFXminDp/l1LEqRHF9OiTSa1Pq6AK/C9j75S1U/eSu
nvlg6MfkJy++q2zYK7ya1rv7LIGHr11/0DOgjpWx+RYGgJcqdBu+NlEm5dA64yVO
EwGaYRKNspmLxxSdugr9iDQv0sWTMZ/fYknMuSz8YL2e7Y+mVNatfYVLFaigv+dB
j+IjVnTOwnrBbKsy4HUaalBVgvIYNmSDfVHoEClm+EA9ZT+BIEkMEeGhzZYUzC4K
BW/WJ4RiY85iyv3VBFUw2iJhgquO13RDrfIrE+XBP12e7eLUEMPa1A4m1Hm1JsQU
8km+4YPg7dI7v4PHwrOKR+SwW7B8jwU/Shl/8VfZU+gOCf4ORgHlOiyeGlYwiMcY
TyCSI6X/gNchAkfXXLLWLR5oLPrFcH5RfQ/UKG4TOXGZdv22D0y4cUavuJPnjnf/
UKgXUFG5O5AiUFE7h+2IIJdPWd4iFCJrbXBumwMSxQI/fyDydkPFu7n/iUmxTEPt
TgG+p5/McdH8lGtg1iGgcMjMx8mlnrjwhAxw8FRjybhwvPI83fiGzKisWVE8BlJt
m9LSnAWW+5RNv+2Rz0hbEg3/x5LM9wUebJDv38ow3hG9pgBp36eMzKvP5pEaDwgv
QLUWLXsFn3UbGlcqS4rm40opxM2iEYnoldsX9mSXjehy1DNm27e/Pbt7YVQjSMyB
McEuYesC4BnZhGVSW44PH9LfrApvJ+0WBoto1WKD8n3epwc1v8AiO6r3hFoJZ9Au
CQn70whjtuhVe/zcJ2EO7re3zCgN+vfvid5y86kIXI8WgveF/wwGFvdm0rQQymgO
wHX3ZITzTKci4g7+9JOOMlwOBrVizMw6RGLA52G9LeQs2lI9d536Usg8UkXB3pva
AsE+PLQszWjFcmwoYlW/JQttQs+RwhV9pPcvvEudhrq+O8xRLZjYRMSkPE7OS5u0
h1ky5nlMQpxgUTRS/DzczWybOAtGEqLj7KepfQJLv3qMxTncOXl20Yq2Lay2WUmC
Iin8hK+Cc76/+6t4H8PhANrFjSpOTbPBEnSwBm4/2SFdObF0k6NRUGf/LP1XkABp
kvzkGOB2TQODnLor7W3igkQG4KV+2YTPplEWslayuHB/SmzYbIyk/apJrdlMdjdW
bdsBM7umQSuaaCmaPzmRGM/b8hJGT0F62i6NqO7c5bk/pDxpRP6f5FmP6z3s31ep
qr4s38LbxMYkEhtv9xmQzRaUwmidfuSB7Byf7/xh6s8Jawf/T1/mzbuV6M6sO8be
nMlsHVFaLnKVFloa3ezQOv8pSBDcYjSaWQxM8m86XGJ1mFIysZpZOhs8L6eXH78B
lBoQKaARixRpSSuhuJOCYE2gOZaaX2Sq29avFQLES3ZEMPC7uGgNYfadNG6dD3l3
UcR2ZoEuVuM75WQeg9A3/lr2PYpWh70lirXwJWYTSL4S/KWAnDWBDjQcIbIMBT5f
I7QzoIPgvf9jY5ENplLQk/pzohLLqa0ZzojbyWWuhj4GIDfqkOnIno2BMl1C0raY
OBqWjBxUurFuxsvOb9QMtEgWVfuByLbBTXTSrVLl58pSux9G8u/ByvWlZXryqxU3
QvXGqKnsE2iPy1sEjt4ipgaG7HIpQ4A5wfpfKWTqvNEkt4+hz7MGZk/ujFO4gLtD
uKeyGRZ1HAKmB4JZP8qG6huPHyFPjoh622+eVvqv/lBAmN/x8cwxxDxO/DBDUd/+
CGfrVjx7Py2Gs0kz7eHmSKqXymhAD6izorjr2fq3LI82kDk8b9m2BZePPdwomAAw
eJB47v6tYYqbU26XU8Cp6yKJwiXe6yfa1CXp7r23GlaUes078KJwAgL8nBA2u7m+
dY4YUxbhl4EYB7GaeeVQP2Db4HaeaXGGZr7ua9Tby/V/4NPdIoVD0S+f9NX4V/D8
/q6wmsWlg5XrbdXKFh4UK9kxhAKHQnru3GT3GObW2CgnxWPb2h5CB4y+wH453EKq
e7nfC1W+gUC7zQO78GeBI7WEdDINUpFa3/gZXov7HRGAxdknRJwJae2MN5oOajYW
KF9vI92csuvolP74BD6X2nfnYHQoEaLcBQ4sOPppJnjwhgz2It4X76fJIW7DbK9Z
23ICeZsg6PhtvR9WhFeU/wCfHQOgnwFmx4CP4sonlSb5IG+MdBpqt68NP0iwFBsO
wOSkoTroqhmIMHoEvOqj6Ze93axKhnfFB/YH35atnGM9vbcMAKPVxM9ixvr+eKwq
tfQ3O5n9QAj4fga39EA8YOrE9T/LvaBi82nAKuisGrST0YwWxIHwINJGxTHQDvFI
HNoooyxWRMTGB1A5LQa3dT7T3GQNXvE/SZaY20ml3fEqgEkT8CThD+trEBHJohC2
hl/E8k31OGTYMFru+QAJvG4Fl7yyR2paWTbmxEuc824rhr44ZuJpJhL0cClX5e1I
DaDcVH8arHZTzEu9vOO2une5KsqBMXzbBY+Zt8y+btm/xVPnz4XWYJeodxdcTlyb
S0RqovGG3gtFTrk1kq+v+wrLDsOClDS2b6j1QzRHnzFEWPCXcIbTg43gaJnVtEYU
7jTxmBpQNsV409hr8fOz3OjcLan9nr6LGxqgbtyAMd6/rlZ24iXCO+LLDXCDufOF
3C+epL0zFTk6q9P8QAnmGAaDppzTBcgVj5q+kIjnwJNJHwbsyushIFvVyCYeJ+p9
rBQxucKgJDuJwd6Cx//TqlG73DFqoSAZRBOmSchcGsCznkFvQQrIxPuNqvn88rFv
WXuoyyQjGcGaI/0KFQNffD/9DX/fgH5bVUMyYJcp+hFAvr5YTmpWQkW02GaLPOkl
taqOfN/SXKiVvzWYHP2yDO2rM+xJfRPg+xwrde9/2xMZtFAoVblzsf5KaD+y+TR9
q/v3pXvyLaVee24fR5EE+QgUsoT+gh7uVjxZsNaGQcjRyQsFKWS4mmWGumlhInOn
hSz9IVeyuSLW3Vq+d8lxZXxbwLc/zSjVqbljDC5xAWpXZzXGkoUVAN7VCqMoUqiP
3ADbolSik1WfGoIghpUkswN9h9Mfa3P7PxUdPhmIt25Ygn09HnhAldK+mPOorghm
HvYHpk/Bg0yBwSQiDb35spFL3HS7u89h3ZnQKi7RiJM/KuVkFqFXk2MI/JAD3myG
OdVQ1Jo0yuXWwljX/XVSjWO6t/yV7U6Lds/hew9REaSXcCWJZryZT1zGlsbsrcSb
yU5q+i9Oh8t8UKasXLkJAx8y/TPnXqa+ylORVSB4NRbZVqZ4Nrp64gXMQlx0dpvL
vZrB3X/stus4w5LKPA460s1D0olw6iMdeYotnOGlVS7w4iKtb6wIhd64JubZU2tG
dAYWIUj8Ls1i3mo1OxqSXDFDKGfQ+sWjyEqKBMR5cn9hPaPRux1c8L0+btGN2ZB+
ptrgdTuI8TSfd2wdNVKbKnBaHhiUemyaP01yTmKRQqjcgf1SybsjW9b7SblsABc+
uSNkzJWrzk6CIJM0qjq4kPPxzZov9GI2yL4kZPO3a+1ewEw4/0WS6zvnsZPdGeI9
0pkqmD4Ag+Fp/7vgRJZKUIn86KjF5bMxggqH3SCVcqrWmnbu+KaW4xenBlIu7Vzg
bR5h+l+rgdY7YZkSPxgblDM/h7UaUEkfSPnlLgc7NEa/7O+KT7TL68976Kk0C8tN
+yIu4rLeVAgEa/ltCIcgDvMWqGSpK7QuIx1vqZVOo+UYDtIcpVFlUed8jbRYZNTj
mJhWs97OKvYZiXCqX4wgUm0GY1IoilJYQOeolYpQLM6/t+eYkOXn4egbtBOczk3A
/TzW7an3sFbDpBkRnW90FuITbEczzWbOGs4bkrhMjct4lrASkSBVle0wiy2rcyJ/
L15fFV+6wXZRMsdbC3duaKcfxfpIyQGs8ZPU7lTqazZqN0CgBcEuaQH7Jguzvwus
8GFcUVXhJPfeJH5YLDdQAfClbyY2nCGnUPfZNUrLcfe5RkbvO658NJZBCMUlCpRw
+ImmbmoYybZ97ALvOPWbEvR3t6JmqUnxy4x6yn0Q4iHJ8VcbqOSI5lDfB5ZyUDE9
dp0w7N9I/4X1kaqQTl7u3ylPAbi5+yEgw/hTusNFAVrrn8qlHeiIklet210H7fl1
nZI9BK3zYcbfMmAFDBIc01q4sq23gpiyXKqa7fyDeoY1xt81j5wnvblqI+QIeV2D
zseRZkGEDpuexHw/u4q8SilWzCjhqlt/XILWgbEp/xBuj0DLbYD7NyYGVAnoqSSJ
F4oyejKUVD/9ODIa8RqRKR9uKm0sSuXPp6Zc9vmjv9pMb8KpqmHnhEbnnECXphIs
vX1sTnDWE45AuW+m76BSDAl0KF3A0FOjP2blCLLooBZJ27VagLK9i7F3DqHkxVZW
pCEKWE+oYSFIztuj012VNkcnHgwj98utuQAbMuBLK+wP7jFTZhj8t+LVOQ3mXqkp
3fa5nYOYEzkBMcGIpCbGvLA9/H1J1ZrWdxLnCYoTSM4HKWBcS1uG1pCASnxt2Sye
+lCZxl1CdnBskRrXLGduGjCiQQlevROaJoGLhvPnI9kzZsWCTC0LA9r8ikqYNuiI
f06th/zTMcFQkUtNzqjDr7sIMagoxVG8H+VOjKWWQbdgTLiB8MFym6NGUFTSXXM1
x3NPnz5+OsIZiYTqIKDC+Gqigu/OSiNgGsLeMKTcktUSL0q2Ac8tVGUmC+pYSLJp
7jwiiDsH9cM6mOLiEx9nd9u+yPboqc+M/6XDb5q8rO3pJZVJ3bSQLjvA8JEnY4zH
h3d7lewYEmrqX4uyjXShe4BUF5672L86yd71Oy8rojji/q4s5It7olA+Aj2T1XV3
vJuaKnxqTCMDG/PH9fnlH5/SunFrEqHyKDDo4npQVz8JXFwk0XxG8KPsCdrKSjRX
6rSqFg9EH7vokdloPJzLIukF11kspiMYEUN/nGjnD17VhGMNQ3d5vhb9XBFjFOTI
uf9+w2IMH8pdh/nNykcQIB50QxsdYzR4LRRtGg4HMoI4+sxRvndSX6v5yFK+5SEm
nBPfxMqNiqu+59O06rEM0Hd2QCt4Z1rCu2O3zdw4M5hwCpAg+K598URb11QnxBQ0
kG4MOWnTjorzAzDegHl2uiU/K8hIQi8Wp7NRXcQfv3iFPFlhC0w4p8omjSd5ov0o
j9NDzkGONzEzar4yNJLo6aZCe90X2yQ9MhPW6izcLcaxo3qV04d/UGdFNFZy0Usz
FcuTdmHGhSZO6YbDA2g5fqhCTVIzTlwhYytyX6jdND8YLRgunjt7xIFLN3M1bBk+
cv4CvUu1mKsk9MDAZa/D1T3DofR0HHrPdvBE5y4EiJpbgs004qZj0h0pT37aWEW/
NwFqz+fmjkzDsJHmdq13u1I89nEg7HSu7CEskD34cfoodDVSiji2ghlclN2yJlAg
ppsC4mSOwRUIgU+72G422RUXlxHDYaJU9bf+dRzD0v7WZv/BMFgUVmaracNzZExr
o/764lDxQTfUXOOQt2FIgsm3G0YnzDjZoWDwGI/PQTQjDfF3vdv9LFafU4WSVtcO
dzQ4AA12nWiiJ+Vi+MmEteV8qcK4aMr0NLYa7HYPSdqI+HrDtiWMBjN5b8CVtjok
/skA835Gmubmykhc/I9W3NzZh9ttskVhZnnALPN7svJk8ni5DKbYRu6dZpb3KoYG
huv2gGwc34JYG7gEdVtVUADGH/1rwo55OzhKjj4RPa/fdiw1xRwaSj9G8RxPiTW0
UAAlnAKjLP+sOJPeB7Ag/Ji+Wg59IP2HnBJWvuUDQfADdY2cARkiiJFTulr4QJav
fCmHbbMNGbv1T9PYcxUqk54LlMOcBnutTKMlxaMDd/mg37ebJvTAv4fW8DKGZ0BM
lGiLCIgqNnBu/2G8VZPpe0ftHr4Yx5L5oylcglHVnssi1Wg5qy/+ATssPymvDRlz
AIWeyZ3P7oCz7r3si1l+CKxC/JPlkVeqFB2zdnFNGC2sQrWa/xncX4vmePIy5tks
Jgin+j0+JX1k0xmut9ujrX9qt4ikbCfttPmrY/cDKX+pwjd9ErYXg5n3kp2M2Xn+
YzIbMl6wqEIbgmD86K0ldX25tyogL9e2QF2kGiElYa6AhGlbopdzy1xCw81Wj5Mv
LQ12Aw533nU/mj6F5flZutDqR1YpYnOxkdDVUPUVcOti3wKF4gCluqw5dL0Fhp0r
uDBaCuK+6b5zM0zBaEVduQqWsTyHDI/0KwgUxqKHedBH01d4i6N16piwqk9+2rRj
aQk97POw0U1DMzaeNm+VY/S7Sfn0OoAduq5ho5/Ug/HzneuAMNLvKiSSqu7/O4Gr
jTHlSzH5s0P7/ARicFLNmuAs3xRZPBwiuOGBnoaDlrSAYS8HY1oYMt1aKaVqgVT3
6D65F/0chyVkkForpGmELF85aDsDXY1rJx552auY1ldJ8AwdT9xmaweZkJyRcPqI
e4EwunZGgx6Ks6rjOgBBR+TRT9FvrQr3/cDHhqCb/RAi2VNxe1eGVPARD8cXqpu8
/x333+sW8uIzWw/GmjRs8TB2FQN9ri/9hPFDxR5SUB2dJDXdf6uQhnEsbiAL14Aq
7FyHXVe8vb4i7BgcDsq2XxFhKy6LxnDmEXJthBCebtjZ3/8iKwclvKTaRW7Lbp8d
dmYWp8kmq/SjDV6cqxOLZWzDX1tQ500oEljvmnQ+4Tjzc3DvyLfXIuFhgFG7idQv
aPGN64uP0pU8nGV3O5BxCbvLboJJr8t5uNh9QdR2fgSMIlEgPAnzIQtdrGLUJlku
FeTSVKnf55BIOaPjGJRmjk81yZoLCe66ZCOhv9YnQHuuPPxaYRdDFp1EYmV72yvQ
ecir4GG3oDZY3I1xsi2uMzHajGH7DLLgiMSVPlW0gLv7aCXSxhP7A5hXK8WTT3PA
xnwxoB0NlAYAaWhthjP36Y16+pLj/n9fGC23Usq49sS5GUV7BfrhV7E1VA4UwQ9y
XL4ySywJNZRfMr23nWTU6INK72H6GlP4Z8ZIXjfO25T3m4b65+7c5ezXQ6ZuGOD9
9Kyiy37LXAUKoJwdMIz8r6XQJTh6tNRJdqJFgwXzMPX3Nw1c4ZKmvL3XILR/Xq7J
4W+nk1Cv4x2nfQtA+VTH51UTKy2H/xY4koHFibU5dv/hTr6WR1BxRNYWZFhxgTpt
7JvRCZPCbiQ28MygfZ6/Cvq0FIIwDq1kqXOuKz46y2xxeji8Mf4RQu8wA/3rjsef
zVlRqF3y/dbrJyfkqrTIPXXJMlgb5M/vLBafSixUEKQEKS3Lct1+wh5lYBNK1xDd
ZlU7xUgBw8Sw/OKdxom6hNESNOZy/X54LgEjFqH9IN27tf8nrCrNt/HWvlDevIUG
4bRn7xZGd6PEvCbBmL7x3yrHUYZ83a7VyEkez/Wo4rj/OSeqoR1cCY2KzA9xGQmy
JUUmQliyrWLUr8u79/d7PSkw2TnDwXzW4uD+cSLUw8neccQocF0x242vhFdIVvzu
A8HSXfTGDBEWQf0afMAmMUkn5ZbCw1kZ2agXdSW9YyivOh4ZyD/mIOFBF7t/A6r1
ebbhxdwlwTDAxIGw5yk28n6x6c6GKLN5rfQflmvD1F8195Z/ACQgTuPc3qQGz3MH
cu03NdY/HC73z/dhLFRMcWsXdRg26041llAGfE0P7szkCPEDYzhr1EiSO0uCnCEJ
tQB7Ig8t6xrPWNsYse87J+mU0i69u68S5N1r+fa653udOLuoN466AiM7bhCSddaY
Lmovf0U2nhOJf5zuZzoU0Hw0zK+L/oiVYKCpSIXBP/Q7vMb81oMuoxhKTdputvo3
VcAP1P+vc+dTA2nrs9UGG3Q4FTEm7c588tMFwaZAuQOHnfZWjU6D65yGTFF+akBh
cB/xfeU+3XyTemJ03RW7JUyYXdDWx+IWLO52bCWnWau04tH9Em69TVaXRlGdaJKX
E/KUJFxmJ6ZoOSxS+QfK6+2j1tqgC/nc3WsFqYvgunj8Nfyn1C0AOINvZq1OkdFP
i8j8is66t2wxYG8BcddhP4Zd5P+YMTEkg6DAk4KQFqUkKY+0MbsyUR8EEAsnFLJM
Q6jPbnVpjDm1zsvruKuw/OoBGubLm6OtTmQV0PhYJ+x6JMSpKNfT0VMd1bnyXpa+
3RTjlveAus/ovSlgp9hEjUIFXDzdsIfQJgz+H9bBhGW1s9aN9fX4bT6kh4i1BW76
dFMSST9ftzh5KNEnpk5EZSPWumu7H8oOl3jUHH1p/JLVYe/L5osP66WkCXWe3WD3
udF3LrouyuBunPL7NlDo39myNDDbJrRA8F6Kq2YngPnama4jFSVXotx/gMWtyhA5
NO33sGA+Ag6N0rp3Qowv0iy4BPmHfEBRzqYot3pIcJ2Rq4rHyq4pufhK/pkVShzm
tETS7YXKfMttSc12NYWwumCFa1CuFL5P0yVEK0ZOH2JcFleqLkoPrT+Z7ejXl+iU
JfOyPV1K4ZLEDfhQUAa7XpEK/xIfYMbEnK7uqN0xaTJ8QX81ct32I5A7qJZWngym
z7jAt0Of4iM1se7xwbDOZn9JoDxf3kwsCeuqzVMLgVuJDNTVIacH2DwlO1f5VM2e
igzDqj0bgQ2Nm7f+dgdOrbu9uc2uHSnQRtfntfbj/9Z8whwgNuKb1CbxdzvjRUyq
IlfdVCf3cmIzo1EFxdaM7iG+/PihLd1t4vqxRIvQ+aOsubX73lLg9u14tWgichgo
/aMrwQUN8pNHvbMPz1QygRKfGFRaa7ohdzTjpy1XFtX4q65YxRoTAkADtEkx5N2N
4YyT6IPU2v3FlhOx8vi/FNIkLUYY1LXhxLV1qjpdrcev5Mou9guC1yol9p8yZYZW
QVZoMl+ea8q5g9vaR5xCEI+Fxcjm0roT/F6jzl0XtGveaNChizLlKjGJIDtLG+U8
tdw1ZSo0JN3MFMYy8FFgcEmaL1hqMA5bRSRTnwQ6boE7hU6nc+vykulD1R+VkW+x
599A9COEQLdS3W/ZGb8i3LYIvKZw9zlgOAGnNFvXcBLm5pzAAX6aqiQNmlZ3LHlw
2iECvhfgIDvUfDfNZ4aQ9wkm7jIAClaEduHmlpqVsXSQQHhtXc1Spl56X6mUowfW
rq6de0BoMAT8bCX0999aLFsjF3nW9whofDcOguyc0xBsXEB5AIiFNLkpTFzZgs/o
BGNQ0b0xKnRGfb0TYP+CdD4iwRaPDwYUbd0vHlHVcFmkMOCYkUacncjju16eYfMx
g9wkvsabnemfkSEjDEFc2JVjIwTvjK0EQ4DS/EQHVmEObWaNtxMKP8f9RLthXEIy
imXpmkhZM4QihOOVWw1wXL6CUI4u/u5MFo7epPXbpryNpUTJJZWB7GmWLlZ9pUCH
qVEOU35jfml9QUPcuZbG62Lw3G7zitb8yq6P/n19NJ/YaRuGE4q2Ep+JBAms8iSs
5L5Fi7nrEW3QolpkHlykdor5jo3ZQTcUpt3sZRc3VAUjZsy70PcOjAejqeDAyo/D
hHuohpI0/EGu5k8prC4BNeXot8wifvzl3ohEF2esHcz8LWZJ1rdHZFTotb+t0B6x
UYqvMEmSioDaY3xhlSnfsHikxdfFEudWxl5b4RBXpx8TuJ8yOIVnB/Of7VhLR/iJ
BRcRQ89nEdgqjLw7F77HiwOZZExO8nqtEK6pG8cyojF4AsqYe+8Kx9qAJuO6QnVb
Pj1QyiYcLA1Cf2qlx+Iy+ESOXDHUVNVg1mHzFXoRKdXgU15RvK1MngDUKqohEb04
HaQReJNopb5O7NB5tmIsb5sLX25/QSFObuPwuE7A4kiPnH4Shy0ogcRiDBglEzFD
8Jpo+dw3Uu5FCA8qaBfD8j7P5f1Wpwn+IxsnHfdio3ApC/29Pqb9ewbPVFxINPWj
SzPpe36S6wm4kNTfeoYZ3z2UrL9S46pXGbUq8OXYvP/KjpSxGIQoQcVP6/C/YwPW
hv3WtMf9HeeK+u3JxDZ400RRXwoEyqNXkmsAjaO+Eypgm0tgc4GGzcOmdmSupmpV
hWv+is7zwBFJ/iUjJPdz5AOx0gBujnBAW0TwCuWTffl6OzKfMZw1wMTWMm5p5ecK
kURRgTO9YwAXu09FgSll3Ky+aekfqPhvIZRBXkIHJTIMk5rS8k8l2owcxQPWaTHG
etx1T0CYqx7GD0Gpbxh7mrPUzmYrxZFUvOV4lwUzcIxHK04Kebk+aIbICxrKXCD+
fsMEdijnQ330iaGYJwBO4iEpRgO4CfMU9dqwb0jalx+cduzsOnNkCr3vJvRhLnIG
88OiC5V3A2iibI+lO/xWsZUhlj4jGsm4jSM/a+vbe7QehSI1VzUXAU5JTGbIb07u
pTU3POPmQyg5Ss+8DoXCLocQITvaLS1v+KjHSfheinNQNRmNR4ldZxUbBfEYX6Mb
OG7qMMmGqUqiNCgNdLLPY0mpAkfaGIHkuCbDeMypEhvcUyjCMEfnNSBTI67LxdTk
LCIuLOKkcG3VrMD/fMYswJI5Uus0l4Auy4Qejzof4Vc7WMtyHahKbSM7sC7ni9mD
RXIESE86N6pTWYVtwZ8sraWuITj85ujZ0rH4W8Jmer71kW/EiGWnEea8EZeb46rT
ExlvUMrrUCKveBRY27tdAiamkwpt9XGT2MKGoD/qotTJYjshUrHkz7Q0iPFVsR5o
cwYP2SqQIxM8Xe0XhutTO989qvbwFLHRTTgBYHmDz7eC86ii3oKUfLtjlFcCjws4
csUNYlanVj5qe+d7AFXg3MFQnCAdQ0/uStJpO8Q8s4tip0JglX5y5USVygsrnwTr
XjXp4ZmgUk3r3R7yrktqf6RL7YNXsxZHY030mwkYNHyyPmUClW3yCsp1j48cAopS
XJrsGLb3MFiXNbOiGvLZ3oPSJP2bQLRhGAPvDCsiINUzsSVe3eSho8QiZifH73mQ
rQnsztHEeaypILbfqspBB4MvPd623cmHJZB1KFlAVnW7r2DjEHYgq/vx1fJTU9xS
vZyakt8WGAVGhxnRK2YXvq4lYG7YHnREd+HQiBx1qOeioB/d7/E217cSL1vSnJSF
b4wS/H/8WQdLD7tXbftM/kbGuWZY2/ihrA3SuqzrnJsEayz/t0F/BmP8ut+ax3Xh
ubz8q59Maon3weH4y+lhUkpcSfp0IF+c+qWRCAOxDFuZzd654GwAARHGDN90l9yv
3w+MCMoBzijR9YGj7YT0prR2BVfGRWdWemc/a7QmXXitNPvjBMEYu8Rc4xcAQH2F
j2a3LV8dp0m1dI5JzmxiRVLdKv2RtCA0xblc+wZTXS0=
`pragma protect end_protected  
function void svt_ahb_system_configuration::pre_randomize ();
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
HlRc//HZIyFpUVfcin6nUGDBXE3KKPlr3y9kF7xUbCZ1F8rgJndDylY+bcjzuaeT
nw2mOkwofHE4VEGLj5Q5cZhPWXuSo7uNtZEm+E+Tg/3AaN6kRwTxx6dQqFUg9mbq
KbFCtsUTqeUB8LFYoeJ+B3ESaWShtaACi+FfDBGPDqs=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 131131    )
mUl2pEqr1qjyrPFN/lRZsL3qTW7gOBDobtktFPcVKN6KbbXcRT3niqjhqC4cBRqK
LX8d7feM4uvvsvd5wRaIFgT4tXS+rA/5e5q/SUmRKiB6SxU7GL3p1BKPoYkg51Da
5Jlq+T1gRSZ+jB4w2gG9ICwmOAmdOAvu1DS3aL3mXACQsUjP659FIt8Y/Yx6R+Nk
flAH754rfkMKPORduvaZZurQxwTsZG2jMrKaG1GCi36tmjTbU6m3wEt7FEE004na
9IG5F4x03T1llMRCL0S2NnGgfOSalYU/stJlPOrbIKUnrdC96PVJcANh0/PVMdp+
3UpdxehDwns22SY7TTFb9pVBwUSf/d6OC4qlowZJk+o9aLyiE0wUDv6nLcqsha/p
0uHknbNwcqzltb5vPyKktuNPIwuy2jwELXGUovmUwUH94Stvdfp+3UCma4ZcK/Hk
wX/4/mzpQYPY/TQtUoUBHg==
`pragma protect end_protected
endfunction: pre_randomize
//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
mtTj5vS6ti2ifH4Rl9ezO+7S4mVvipjlC9LBrxJ1OTFKzu7wtx5x0WkSWfbKVlbQ
50PW9UDu7KW6WWiLdHLdLc7CuKj/OvYioZU00ytFYXfIg/i2t4DgAKEp57cA4y/6
3eBRkZWEFvNwmgnjSirW+SXc65O3FBeMmw6wD+O0Kpw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 156753    )
d3autWorWDyW/qRCuOoOVU7sFjbdR9gTzytlt3AxtoEDmQbnNlrEv3ga5kEntnKC
gBcXb5t3ee0daymsmIaGfHZK0kQcbD8NVLOOXaGlMr00NP+h0EbHFEu2imcb0qAl
YZ7Qft5UcxWsDClm1RHvLx5zSK0zvukqOX+RaRpyyoAF9FoqaO/Hl5bfZowqgLsf
5P35X9GnUDwbkFKtQJQEr7LgxT1oG8FqRCH9CEv8jWrZxKPYapWI8SdVSQC9F1Ha
wFSlO33UtNHXsU/iw0kYppKAjDUl7Ke2Gq06DCRGiLx0HHLAyFYyrgKsPSVRMtlp
1oN3yIBeBTwjPpxertPigWRZiLuh8ZttqL97f7wi8PKt7DXuPfEmhuf/ZpFZJ0ke
GBi3rxVKUBo19slPmrGjpDG1aCmkQf4LCH3FY93uVNipn2iaTFw8u9jqjvQaUU7O
BeX8ODSSnzcXklN8qZcoeYJpHJ+T8rcdMwfbHs5IIe1Fv3B/X6aJi5ZQFFzosP0m
GJBh87P8mDHXmPcd+C4uoPX/BmTa2qF5SjmuDnfmGrbxHCoSbRURckC7kPQJPgvu
3H+S7nf1NGp/C1c2GfuEUQnmfpliaOPVuzoCjgqyu4q3aUxZsMS6hLrhu0in/7x5
H4FxPe+O2d8r/cOXcEnjiZe1swiRhYsCkW4jJTvoFdUlC5F0C+Sdl1O3xx2Nv3ZM
axAc/MHWE7/A2ycdKAg9ExY+KzoA8C9jAo1so7mGmxPD5ZU6U0vsmFVhaeV1ykA0
jJtRqJCdnphoYdiYC0LXu7cs2BggXilhXH1Mkmk4oBCWvUkB8MVZ+oCoTHNnx8Rw
gQLHXl2RC92GZeeF+vhIdb++++LXkPrEAgmC80jRuaSY4M2tX4vNFeB1I0AULRzz
UEUiw+yLwazj8NehkbGvoy97/NDNqhiX0baTUQm74XacHeqz6MA9owkv7NJrxjYy
h/qQR6u8SPwQ8HvX2vRf9IrbX9rpGkDGOJm2nIgSrI/H8inCtCg4zhkpwhSe2ZAD
Hb1WQo/lL2hcwNgyCfKt8ZgMDHoJb4FAlT5BC+qpPJmJjolV0qUbwl31XTgZQIqU
fgqb8z+rfE8zqYGBI+gxSRxLH1HDi7BULKtTG/OYnTcHgiGxtYfKdhJCVGSiOKY8
nhZOs6ASeMZW8UiXYbb4JTrDjHv1vH/pgkYyYhHwo/9idWRo4f1APC6hWZ5lkaK6
fpBrc0lvliHwduXx6QxNqFMmjoSJ9DlXL1nBKfstXfrTKqstK72bcyERHqBbgtfI
vDYqJCS/48Bp+AXcX/xyKAGmDoC8BDokdIH/uD/A7m8APadFyjWNFPkr1UulIQ+j
S1kw+Y+/9c8qp+vqzZa+Q7xuBQoq6vu5gmhU87C5tl8JHixUttF/YR81J8LXCp4A
xzJq1481+wfZ/3xo9z7UWZy8kLsvH5MzinFw3GArDq2Ed9r+UtvXJoVnfT1AVFaG
leYYT0oQe9I3w5TZKwV1rQiS9eOfc5MyvJyGiRhE8D0G/B81F1dnAbA06j254D6H
nD9hqhiHR2wPG7pQzMWVpExIG8igSBm8jXWIu2qJuLCHG+uG+I49ZNDhPCMOh1uh
t70Nwq0n6dNFoMct/iRqVAbaWA/hKXP7Ctx/rue3wfprRmKwcQgy9bALy54ersVT
iaG7p2NRX9er8HEkXcuey6DmF0ayNqRSrvWnCM3kTHX02AraEXgioU9qcdRt51IB
D3exURdG09qpYdSxSfxtWP8A5gRQQYd4wt+Wi0uXDFfM2AplD1ZbHY4+IayBy/iC
uKZiniR15zXR1KG3OLWdwTSSHR4OJNcPccphlZDuukuZGK51SuEydZ4Q7LYWk0iL
xUvcYBXrGPaHnxg21GAV23e2xcg7CPRy54Cwb86B198iBlIptSPh81SHjj7hophp
LXr9E4Hl2aNyv54jLG/96sm5QF6TqgyypMLEiiqp73jYo193GlQqWegG6+gJaEKB
7JbtNuhlJABLDjqZFM1IpPl9b0PEEPB4BwqFUNOSJBSPiTLDrv/uf8+H61OCs54M
4WziGmyX8B+MlSyJRWXqVs950qV8fZfm/lCZ/S5CqH/aNlF91gfBUyxkojJqcyRV
Gcnb2KwNn7gimfSg3Qg8raY6kQDuGvdsDfdjdX1TcW0v2nRL40QkyAuekKw5R4HQ
r0ci+XyrIRQZboL+Qyjlk4U9Nr8XzrjcajmSPd3umb91YsA7lNkk2n1cL3SblASx
pSIgZMXl2YpuQucBlbLCr7D9m/94UKy+pfqRpR5ccJXZqqibCYJ8Lx8QzFFQVIkM
DK9c55exBMaReD2OUK4uSudGPNzAjAWmj+QDpCOER3uhDc4vO2E9DN44MSPZlN2V
hvbFI+xkQyOJk3rFfsGRUPXFuK7bfL8QJ0qP6ftb5k/NwaYckDEpFj6F6vng6AmB
ufd+WfwCfEMVzKLaC+gd6UKK5BncnyUIqVoChcqO8enc1U2/C4hsJ+8V9kMKKU+R
A81KZ+hM+E2lY8XTuEsLbg6bu+W5u68X/yagFKT7BQwfMo7BvAAP8zJo0JO1wqEO
Yw9Q+Y7J4kGTPVj9bwmsD22byIlu3YodjovkG6thJQVUJ2h5Wyyp+lOQ00Ns98G3
g+fCIZj9N+JfVvd+X7HhzusMpFfZqNylQUiRuOuZxudSFAQeF/6BRLiwZX9ccZC4
Ol5Ee9uOW4G6Cwhte/DsFhKVRwXms4XFl9eUBLeaeK1oa4zFi+g2GbK9y5PIi8sy
NlZcQx9btctyfGjewEtJLQ8E4szVUIzLCjVv8QmA00k7T8HE+s2mA35y7pt1niKS
wzSu8yPYeMNwIXL+2+rv8SXPVkLmMHrCASuRdBIC60VcBvXlONZbfI9YGJ+6d++c
Stw3h4KgJauq7otuNgq7xUZ2FtRE6zSL+wYgV0dtaIsuOtVWIjCurXMWuWfTxfTM
x/pfDUAydkYWG82rXdeuSK9P/JE2LSmbY8hPx2nB4hBBQV0Dh7oNjLJ22j8no4CW
oe+68IR3/Yv3Q8MkrLYECyubCHJVkm0cvWa+ooO9i64gwH3aKaQeR/cE0FK6hZgB
11x9fA9lzcFscrtiiq4cTanKxC2XJgSG0XwonlUmjQPmOpwzmklEIQaFNJkUYfvv
kWbXRo7llZbIiahJXaHrejN+eNYtWElbiUdJ6LuKKlDiJoTAyeEtR7jFdRUjOOvW
gEJf4HLhmptr3gMMtdZdczCWYek/o/gak1OIdoJJi98oqTC76efkjRW/DUSRVj09
l4gMKNzS4mZSaelw3YFILCUBYPPC772XDw0FrcOeMfkyL6t5u33od6T6cuuHu78s
EdOuvcoq4N6+uay2caQPrlWFZc+f1Ylj6hgmumT2sYuUbxsDSKAuXkkN4rNmIv/8
bx7oN3MncE7QWui82xjeD21Gr/024V8jvXSw9e0JJpT76pgSaUyLi6FhARaAXJ04
FEN9I8hIdz+CoD/bRndOscB0Mdnwe4Y/auWPKj21EEZ2KiD6ksvCNJ41FhYtnwQl
2RfPwgMoj9KX/1c0dlQurw2Z5l7LiUaj8SJyt9g5h8+M8P8wpZx6CRYLWwMk5jSC
nkU6yeaCE7izDMY5sR3nJC9q/5WUF7Uudj+cGPbHiIjPbRjjY1blrsyZRDrRM3Qh
HiCypHHzreWpcE0lnLu5EgTR9ua77CaUbRag05L+skZfEp/qsj9PX+19lhGpnnYU
T2BH+TXolnf8puGGiLyq36zNRO32f1l1QEQ8RPwNDCIbjI6wAQ/adND9H6JsFAla
pXoth1EcSNQEvkGY1BTn64hPOcE+ib5w0YOmlZyhZjKyUDZY5xzkdrMq1BmEhtwf
UEouVr1a4RDSjmw/QrT0Fa2fSvabRaRLHrqvuVMfZ4wvqItrLJ3K0neHX6ld34am
daQkE06XRhdfNnlGev0DQewt8rfslYEKA+zv1jqAiwtQH87jmTLgYEshHcQ9FKnb
DyNTMGIo1hqvJzDiIeKmTK4iMasM1St47kQvfzcd8WfJbuSASEAAoz6vwreQlQgX
Agh3SZCb5Iss81kja7nmr6WrXG97KNvMfyAevAyz401d8A189FLvVvqL77kHK9fS
Q3V5za2LlJ05emaxGiEVeaoeYSDY2MnthSE7Pfp5vQtX6+JWfrhfYJXtpunbcGio
158wV9UtrjW8DSDu3ZIqGZuhtCcLCo1EFKfZZft/2l4GEle6wTyQiPFEprTsAI+o
TMnmBoh05Nvvpa4ep7Z2zlNYFPChFehqd70EGKSE86laLDQLZu4xYRNRzJIflaRB
FLwl8WUrL+FApXRcAEw2++DJaFF99ypp9WVwUq3N6H4yt1DICh5+ob+Btj5eYGg9
OFpvQcFMXeQxzAzH7ootcIO0A5oIMCruoZ+1DyR1VoZEhkzQG/uuTOJvMN8YuGvp
QExMeHsxk4eJGKsCpdUazkjkIt62Vb41GRR4TzmDqU1GhzesarfgrI6oV+AG5hQ7
sWpBa/jBGFpaotaeNunZnhp6oOilrUGRQx9xDksEDSb+X21Ifl+yWMhp5UVv5Tts
zQVzWsP20k6RbMCcOfhfhk7RZg7GT4AJcsP/WH7uDP+imvbzOpilVcgIXtbO8Gr5
F0MAcFaqBXDyUMDDpYc6GIZCHUwc6Gpn2NuWFsAhGC8qPlkOzU2n3f6aTLZXmQLH
NJvRIU+be2EAtTXw1l3dsibFFn8GtESNw0742WOS81y84Hna2To4sjov+JD4Y8Vc
g4VLzykoxcjvh7NzNt85QgIun62iiHUvXYP2daUhTG3eAaVWNMxE4fIx4ObS4MfH
AigO3JKVE6K6yQDjGvl4Fr+M0Eb0BFHwloI1xQuGkDRqO7XtgnZxhYyTgLG35hoI
H6LD74SIUnb0/o6LfO7kGPKEpV/WAYwZCyVTkJdnCafHPhMJmd0qAmU2dcuYzX3B
8Rknq0i+98MZlev/BoOyKWDKm+f2GszFCunp0Rql3nRV0pO3yMTIiIQGAO893hUt
3oOCPnbqeEYK5U57iJO9KHLWgzSSzjMm/w6AYx1NgMIcDErT5vq1aLjO96l0GUq6
De/D7R3ezd0cC4xB2C9sJLEjW8Y6CE/vI1kDwA1ZU/2Q66TuFBd6aW5WsVkQTJk0
D06xHxj11LZ+1ifIxujiVIWYe5MplhMckz3vHyUR3GxB3fkxURYdvV/DSA5V34Iw
h93sCZyqobChIy1ss1SWewwFB1pTuKyws57baZ2D1ROvQXzyHPoPizU3yfRkCdP9
Ue3mf3XF+AkfBo74OQ8wAl01AaXdgdkqRvnNCz4p0Wxr23VaioCHV5ZFembj8VjE
ReZK90743LK+XwJrhgcrXvLpeEa38E9lExIish9oRbaP8lKmzlOpJm0PYo5449/v
qWSoE3l/f8EMmvfic5hjQSHmbW0Ejs0iJPWu8RVUSH1Bks0NnmZVjc9ThsZWiT1Q
uWF6MAhNaT2Sfj0BL6I6Sp8knihaOCq9RVkl4lsDZmEMatmW7AYCc+UrUxcTrK8W
02sZKvZt3hnebYJZ/cdwS1UTuggYBCE8F8MMpMx5DHkII2GVhwc20TEuH36uX3f1
vaJqU64yeVt1F9LG4Za3hUvsF2vEEchqCemQJBnL8IxB25GveONdmlVfPxmNOWOG
4la8GakFt8TnM/otcGEE1Qg+5XYZ5daYrEExMaJHGO8Jl5jLClVG2kPhY2f2vrei
vkOkdpJBaedsw7JT75ghnX8zyxbcgjgQLf/rUMzxpV1nRv6JPxEvsCrbSNsdIvSM
jeN+pdqUIS+4ZIpwAyl0g9hRC21rtNAC1OuUBxskuREnQq8rFq8d2ePGjTXc1mWZ
uz4SjLDbHBrLyzkdVOBpuAbBmFYKnoSG8vZs1k30B6buOhc0qbP5l6zFzNMpd6oV
LGfeCTptUgJV04eiKD93WJ8v2cUiJFlCFmp60Fr9/gdby3785laQeO5Q0oe1ayfQ
57vx5FzhOhKpHK3EvZQd3K3cCZj2nS8PXFfMXoU1uF7lK9r0gKxS+FRufTG+zQhu
imezxnz2VI8MQbawyf823nMHuZMJI6gE/290x3oJpQbwL7IwdH/bHYLc2Xr6LDmy
mQ5gYywvjLJTcT0AT+qfSndHB5vRkk38aJFJ9WFGwJPEfn5ReyDbakmA0ZrO/1Um
OfESwTkH0kO4grMDUVw3dk1dJ+flxlSMeCZLxQqPlt+TZR+GMglj39lX0z57L2uW
DwS6647/HeoWvpInw86aeYh14+iVbRTR8m3BmuvxlPXTG95wYLx8Lac2bY6qW2ri
4r48HGE7rNRtwmTUdE3HZXdDgYl+Qxme6HYpqfSAEif83cUNI3HDKTiCMqTs0tyk
xzBGiuuloFmSqxjS2hsrlMv4S92sT8ECRoRl2CFx/3/Mf4NUDNnXSFECNn6A6PqV
oaPnKfNUVJzcI3zczxumWOfZmCLqfuwtFfnlcJLCOwowK5zIFLeeVQwMlbgcA9iP
bxqDY4/U/xn3i8YoEH/pDb6L4D9jKPW4Ln87hRrjg56WnQuYMmxWAU7/flnrmiaT
sqIrD95UWON5j/kUnCx0AyCWGdaCLu39q3u70zE/C2eWQ1D66rnERg6mXFpfu9U5
y8XdLi/d9bO2WefppatmYdI5eDVU05RTM+nNVy1f90fgwq/F48nz/KeLt01xehge
QipThpMbum/esZ4SxdLVCrzg70HGafvfMGkqLYB6vAO1EFSFZTbjUsruK02M8dL7
fgrsn4xgrh9zFc4OWM2D94MsV9gHxlEt0T/gNz/BXQp9FQYoUfwCStqsV+c26jA6
y+3A5MyGQyWdzp1kv1NesobwjgSDfH5YfA8GWmVjV/zxreKnnwpfvMp50FlTI3P2
gTAix8W9mvr3aWTYBhaMrwCCpl/s3aFbP/Z4Ol9oh1zEBa9JmiYt338kjGvcv9I8
hj4GQLua2NmdIXW9mgrrL0jm0hwm7RHJa2SBPV8vU/3XJ6T5lPbfKYNw9vmFXcCA
Ks34/TiNBURQ89WPJo5/vG8SghDCHfeTAlCJBTR8YtaVZP9JKKBCR9GxcrhwiLHM
VfvsfbyjNm0oDJ3fnCj6zufR4U1uw57AVZSlnDAIxWHWskTU9XcsPrYWHf2HxYFj
FIfqLPfA1tmATH9T1P+VRHfZtTym5K0m2pLwgPjMJg80YfXfT6a3kUTnI/DpQcve
sUwvdkAeeckT1hKx1xzXs2hGNXDV6tVXf68OhJs9fAVyNRim/THaL9C7tj8ILXy6
fwtnUuxP0Ipsd6aMhBZy+0ykJf+rb8tvGbpXhp7vzY1qkoV57mtpfE5AKuVVoP5Y
lAfxTTMm6QQwyCj3mt7vP1EozojtPyWbzL/2fNxji5T1NJJMIrZMhUUhw82+pK6f
gIKoDSyhBUEzcBxZPo74+HS8BwAwfH7tbMtAW+j03OHRwPHtPXPN9NGVzenx0kwp
Heibue2p3rMLOdwORWMTZodDDfSiXDtkQPvtjGLFWioQjmcViHxwKD/9kXX7wih/
wrhtirp7Xmo0ny2hns6fnqX0OcuIokO8JdWQN9yHi760Qhcn4GHhVboaKovJxPj6
4QvUz+17AHPkG2mFOqNxuszllwnxTDjQB3p3WCinl08teZcr3tlftJdXCuFT23SC
66TxQyrNeR5b0QFWH+MBInIWhIJzOv4ux2a3O9Oc4gI6gug7Yrrv6WVoPVMEsJ6N
VE7gbWYqB7UShYFP1y753TEaw+9nbJB91YWkG41mWm79Ai2Jx4ciL18Oo9+ZOvGD
ShXeHTw7vdpfpeCwid/fdDiRVHz4f3uUpWBYIqCdhup/5h9Y07c2+mVRccnhTX4D
Ck+XZKtDnKpynwkt3QietOBN9c5nzfAf9JohbohapXcHdCc4+4zEWrDBzK2b+dIZ
TGB1TIIPyy0hlOimwFbHq1cXYS/ewMxReUeir8VfjVHREYTs1fvu/n0rY1ZJkWfx
kDJpju3QET4CQfeBIjf4oBJjSpHAIl6vE4li3piNPEwMl72DjMY5LbMXXJYdD81r
3hm/fitrcso8visaFaQXhoIUWBLyEBPIbqfOzN1bsdS80g3XIqP+b9OhR32HzVDn
7XJErMIc/kv7meaK7V57BguEOIDRZKrWGhT2Rqr82fcXhTxfkyCWG7p8kGwXTnm0
DrY5xFNA6KXamRi4MPi4vTHXIIVKdDFCxe9ltCpYbypZ053mTJfa1sox3pHJ3NeK
EBqAccmVE6L4jB2uL1eTalhyFJAqyroSn1MvBBLrtPpi0THj4rS6cP+etjSFN7n6
kNvvl/3ZCq7chV/r/mEZS0r3W/iMBhI0r5AXBkQyGb1jGGNlKcm+js/OaQriyBRn
xYHjijKxI1zSHtLFd+8zberGgagmvRHsSYJfAd3820I6kj1AeKAUuNILkKCKFSEo
wjN6MAdaLXyX6Uk7cCGiN5ygCVuDWLhudTkvRqv84ECpE/51YQg2xWkdMzFH5Pxt
00xjp9JkTYsqrL9KHcHV5uV+XOvDGQNAh+8OkltFP2by/cFA48x29E+GsfMl9PE6
CPqHrCnx0JHB0qlNfGKPVrTNzmMF6ui9onLEu4vhudxV5QvouEnATGspFMsTfeFk
3LIIptxGVA2+skWRYkHjEiM1a63Ia14nn3jrOcsHtL8qNvMPf6wJoOE4YZ15UCNZ
61Ci5kQBhkliE8XkTJksdZkrTF8fP4ajmuXupSQKopCn5n7PIvpQy5oxpsrHxwd8
7yqCFsIsQ6IkrX5rogtN040N1lXLo4HdYQ+QN7Fzcz06LspMowuhTvRQisUZcgRE
IEUi9yg/TF0EQ01kjkuJLhB6sX+CQ4vzQqjvptW7TEC4O50ViW3oshooqsdQDpXs
mKR4ctjK74MfDumXMkd4HC0eYYtaa7NVf2EQnd589LmePlrZwuPXvnlXNwPYysVB
ZwzykZn51LMvClukMi8qIi69YVwmwGwMW8+f9THASYJfw5oVNpx5gjc40usu4zTp
IjoRfpckbyfPtZLIlJQ0xkDYp9iknOAEtCLdGpUpI70u7zG4FPb1y5rYGpFgBppe
57J1/GhBDeojNMEtnEr9MczzCv03oE2o+llIloLxbDocbtl4wviZy+r2RCfyPBD9
pPVa+2XeiX+QPeCBHCLFBr27ixUx6TVHLfcIHOfQ+CUPS86/qjnt/AxC6Mz+NyMZ
5jGLACJoetJUDFQInZ+hsdtZoVoFGZkGy72/2Rb3Db3Oks1jhyNdQpGOtL7Tyh4I
aUjs9bs907dsMZ84D5XDoJXY/jaCSW2yNkp/iOkCvF0WcL+eA/uqpO56pNuPcgyo
K0W3UcxTgSnVSEMBtV7AOYdQTXRzUm1cXGqO7Aq/XBoKTq8VpbArrLSG6qCt0oZE
2T3na3ASnNTyrF8uwD9ryvzumCZxjIozwv7JOjE6mslOi5WIBKnX2PtEplx5bu7Y
IYnSOUQC80qZ7VCFCHost6bG1hxDSIY3Fv/z6XCFo2XN1DTA8WZ9zRf1sw++nUpA
McG4tgQ2fuNVMSqIEWHy5rLxc7iz9iRUCKITGIa+KF2DQExD76d2Qv9NFmTeford
EVWqQR7sX7/BHAlL4cFtQaOnXUx3elPoizHu+OlHH2aXpzZeH0WpMoGYKXkusNTN
g12eK/6pLSTv10ZCKdNkIjpZz11KNfkG5nSKPEVB5hD2ERvtBF/+Hb4d2Q9Lj7mt
byX3jLOEwWUsYQ1LY4xH6kQkcHQqr21hYx8r/ff+pbeQjyOEz9BMmmS3t/d2iyJ0
19UBtDxvKJ9uB8l7O/7ZgJfaKMCNKc0EWCTKQgdi3pt/Xeyn0gu2rsoeUhHTYHZF
5Y12jWc5KrTcvAXHP85cMElIKGME27qxtDUn5zBzzoDuKvoeK4gjFWGu+NvrSLxi
ogaSF9/cB9ZAIo7oEylilt8dV4TNA0QALx9kfFvKKNKRI9OBpPjo0MlClSoo9izC
8Jf55B/m2WOvthWqWyQhBPsmJLeK5sgoYefuunM5TQ8l08PrX1IBM2LWINaAsHMe
1TQXieUMrKRijyqPI/TBnfUAW4Y85U9ZeNc8bBUban4dB9Dy7HSPqx4dwNz/HHpS
HKJ0YpOqSsbaP1+UalbkbFGUelSpKYrSRnGD5ZZq8mgmYP2TNohrrR1hJmONXAxc
G+UDKm/gzWQF8IvOUIlKlrn9PR/7rLZRpWCl42qZVo+fWH0DX8DOBuF4SV592wA1
6o9NdlrxJ5e0NTemRJGj2I7+1B2G6Yazqh29lOealKvWf+fvrfIoDdRSy9tf9dUI
I+Q7Aed5kkuxji8YYwKjkcxZedYPDfA2IkGwo4CrUgOx7QK8iG/K+WSk7m04HrKE
gjtSFmwO2twO0cDTI/wsmfA+dPLghtOPaFRpoyMJbMNcCSCEQxcitLzFeLIMz4Jd
2KDyKUzteq5fwLbxPhaEYquugRSy8kCibim5zxNPG8pk++fam+zeP/dyhqZ/r3vz
CWcS/8gzpNQI0akFi3VcynDu2QO8PD8p1qNqSrQjZRy7M+57a9y9uwAgU4Pzb/3F
MLZ+RSkC3ZziQSlFX+osRlpDLCVPfRmmVCG6n7jYMtK1kesUwh2oW1Oxwsmr17yS
8XqtabpjsjvEYSm8IafuaxaX4+I7YoDzJKMsgF32WAJxr8lHSvX1PaGyZVXr0BXm
B2XvNzyrPZU7jtYs0RQIWk6mrMbH8xgMN4Mh42aEoy7m8aXiUUcerKdjX+6M2qRA
RW8n1Q+rm8gOW5/9z/Fr6+0d1IzKRU3TJ1yT8sykQRDck1vdnz1lJsI/WSwCxJm4
KVmm29Xgt11SAsiOtwcDsGzxp/noZX3RZa7jtlE/+MnVzdgG8YYIXpXpLynR+azy
x5wFLogtl1KAdWGma2OzYVAhm9iqKppeJJTGOD6i31Ooh+W0x1DUEq1hSWueSh37
HEC3D4s5sCr13r6QXMBgX8p+YYEJY1T0ApxEvZSi+PFOCSpzfNcrB5dgtZLczqbZ
ozAby3RVw5nT66oN0S9tQs8wcajmv1pzO5uafpDz0HWmabGzux5tYiKLbnWPyTn0
f/DMh7KFckKAyo4L/YwPmaWnXocbiy2zj/mbMUVzwoUnAloOZwEo8OqkXu/A7tXZ
KFVipFfYZygm1DI/YQyP78pGTVY5G21m967AM7UMW0OW1sUbfJjkLP5sHa7iJ9OG
oflEq9GwA9tmxhNAepLzmWDPHocNdowmzfIz+EbTtWfL37wAonApbXID/ZUZ7pA4
mUAFBu7Es6UL6hkz5whBEIOwWso6Ewumk4wPAvxI0vy0WyeI+IjuWwZeaPikOJPL
eF2hO9EpdPczGSqyGWCiYVaVHxnPuVOTvYzkaYg/MZDlwrtILX7GfTTtIpOFJLVQ
+iTFBKejz+/p8Xoq2moOOj5uWJcsp2ta2eLHwMhag25A7fENPJb08EPwzQkvshkY
vxTBKuB4u1F5dOld7aixn9R1yuZxVEVy+iCpUGsovF8s3hJodi5O+ncUDpUAQr7c
dPgxjrYXXlSJgIyjpkr7XvcREPPYXyGVbEod1SL5NOPQDsPeLboqW9xWXJrMIA1t
OYUWAI6RSJOtBwtg4NzW6abcFJuN5iVVPRcPcIX48QIig/PLhcjJ1h9eQ5hiTFBt
Zw0nlE6tV3k2Taf3w+VMVWJz5TiwJotfJKFLeFbEXz6M6q53RUdTkuJrzB38XEwU
gZ02jhZXNznYSszQkmOjH6xyg8/EKt6BOx+1Dij2ozLOKnzXEhoEPxES0GrPtSTj
3YiikE/t7aKhCPtg48uOHz8GJG8ejt9SyivGPvwbaecwj4B3acXBcPe4THGujsZw
Ccks5PVRS1m7GIyUHOlGqirS/oiXbZkzLKNQ984rR6RIFjtjbCp8yGuOChOLn4fW
g2NY+NPJSnWhlkb5C5NYexd8rWNyoFljKt54JxXc0jvv4dJXKy+OYslFbIDjWhRV
xNHzXartH3CBEiymwgPUfx0//I0o6jLsVqTPm587KYChqlXU+dQdLpfkOUu5/ZI5
IW2FZl6NfRY2KjO2z3MsD/m00TAb7XddBIzw4hi+oREv6m72/3JC31nVPzek06V2
YZdNrPMwpzPhVvNjzuBwFo9jZ+7V5fxTtdbgi0JFxNMiTHN/vKGuaKeEMjnLgd3Y
2Ee7k6eXyRfwKj4cE32OEaByxC8yb9goFclvHjRO0ModFE0jukX63KnCwMvsHexC
kHYo3jydcGd6/tPsM/gtCQNNtbEX+5HrYoBQXggZr6lp6zqkM8WWhXlXYUFJGzEA
LlwnH0M/1plZ/lW4bkYQwIcn9CAe9GV6Ojgd8+2FZaBNagIvcBZGv4e/7wU+my88
tOS+Ss85SvgFgfe1O7tcDDtrvh5kUmJLlP3El4rIzso1vlotpqCjOM84ZVG2381q
otntTmYcQlZTWnZw7kDiqcG589hzAJYTLOu4Gsi4cUEpFbIuA/rUBbfUqM0FGZ0X
nNVVMwLB3YKoPrVXE1AHYoHHtKjeqckGjUSUF9V0PX7FajgizvfnVrMyYi4NPdl4
xFw57ZP5ZlCi9JyH8ftciO732oKB4LtIdSKVvMmMkNs/udMAXVdR/sYsQsKVTbSb
UMBtk2cgWObUYmi2qXpRUN5W4ANFMlnNJyyOFGKuJybEDD6xvIecPLh4bhGbOe6q
q+K4RCfw1avJEAOZnQZuywi7KMfnzD+vhSfR7OLcdz8PSiwHlt0afOKG02irIqc4
l4QACYSHO5v0UxmmHKqAjfSqfRtpLp3azX7I3UoXvCbd3zB6KMOeD+pf0JIiggnc
EDIfCmyf3JjnvP9fNFM0MdX8xghVmhHSKnckraesjL6z66UuE4Id2xWDQ/m8ETq5
vPlmiZfz5Hv3IJmZS5z8wXajOIfxA5x0xJSHzb//7PlNdgJjMOjy407YSkJ3I5Wd
HpYvCGTH6W88is0YKI79xyXz0QoWvc8ev0Qgp/1YYG5DwKZMDWLcMTD1nJnMqeyU
37nQHU6tYcptvIqJBMDiaEDQD7o1/X3j9qoSLPQvzP8nQ1PPqDlrfnWvT++epwwt
u0nhZSzEwboYXWM+msoYv+JHEfo4MGmH0EdTpSk1pBhyGqzF/BXiSWL/q46c8UTE
eF9istZeUCumn/SjLBe81T4n+p7RFvRxHFAKPqTmNou6gTShLX7tgGe4pEVkh5Va
SdvAYMno5IZc4V0F+323n1K4JRN8brg7oKrJUeCm1isn3ihlTGNKLuebsNiXGjaE
UkQuM1rPe0CS8aBCFyd813yS3HuloPnpwLSxmCRZlYv9TraMFyOWFOmNTi+ovi/S
H9vXpVdKx194jSIrgIIkMrcelx+gwp7r6BWxfeI6MOzg8BhaTotmhMDwQIKLpOIJ
xHyv+d8EWW2CTLygGzelXHkhGmp+4QGYPwvcQ9XXgdbx7XQhyHuWX04tz+wOJtgk
o7XGO8/VztIUzKjVi9cr7qi+KluhDyXSp7i5gr02saN3a9ucSnV7OhjU2X97f2Un
vuNG9OPbR8/WOg96u9IPWd+byH1ShzRlTwV4YWoPDNgnJxFOQTDzBgvOU3ba5uZT
aErxfl3D3d6vy3J584FEqVosOjE0pGXdAKLtkKzOEeDJbHyK3vZkJCbLsM8fZyhd
5Pd0Xu8QoGaORIZr5Umpnz2mkL32YfBSN93RiHUlWsbimm/95AscHfY9HLlsgQ6/
94rDgFtK3nr3eAe5oJ5rJQkvZnmDk/0xkXIp08vstq2nnyRDxtQN3yAQu/wveGLv
vw3FCAEo4xpPpR1/kZSncbhA7uOgi8aOv2RJSAjk1chcG7E3k7JrpGUlnwaOFLqi
apJ2Z1I151+Y3qMSm+zZHcfcwsebo8vlrHGcgNnCfL6AcacovkwRaUfKhXM1iW+G
De99DufXEdf9hzCEDEhqbGivQmtE5H9JxslyVdiBd/ByHSE27VaYci65H4o1y+PJ
AXP19tVUpXY/SMWeCfVTT94JiU5WOpk2VsmN2eHzGb8YLkCFmRZ3PGxG76XrelwO
xNh4XXNGEKWSuaFNICDXuPgs/9yGunRbKhRSIEVcIBvbDGR0KX5YPzVTrVCq5UcP
uXECpISkhQXXUGVT9uadUrsbOaz3l5y6pyNinddhdifA/NYEL7S0Lje6m1Cj2GO5
Zi7Xub3AQmuFlA0/M3okND0CxzjP5NTxwSwheUPciXx+0/YmzqikIQA9+sBd7mfL
UsSSX17PUjyG7ywaA0ZJuD2YRoVdwg12zb6fCWihni0UoE9c2WyhzoMk2hzGEHKQ
8WQ8YLguKAPJlpE9LDaIGBELGZPawnnQM8qNyB/J/pBqt+I618rDTfB9qfthr4i0
6IFcKtSzsCw7T/J2YYRhMuv91wwxQWJrO78NsztWgXehLORGXmWCNzDzwMmUgdWp
NDOIZXXEkE6s1//9zqUDGpuns77v2tGD2OUbnIW9Hg8hf8XfBmu8c9/PcG6qXmEL
6OSJl/oGpZ0xS8JqMHhsafrihUgSshx96SI2v5ZmEnwEsbkk/eSBTiPQUNB/Od7I
C9Dl5DP9odFSzivrj/j0iMlv1L71xbSlbF5oxEnSP/EeB2PIOCIb7NEn/Vg5dRbT
9vkqNwzAZyjFMhSombZVeiZQ3/Jo8w/bQDA+OY/T8UFPx61uVGTORbd9xNDiSBW4
Ri6HcoxJag3snXMVoGqyRtKd+MBupiMNytUT1lZx4w1LIOTHmz4aiypiczvBa1CQ
3/NYIR7OPIbHGi/L4qoRHDu3NHRwoHQnG2qLEEX7Ot5UaA//6aTGIy3P5Wd7//fn
MXg6Rh++XIsigpuyMx8CmJHONaTYwO463o2RKJ/hMdBotsMO2h+peiJ7ntiHmc6L
5ORSvsJhJ/JFwXoJzGF+0l9WIEoUuReTnstrMsBvxLR3AVl5OPVteOcGD4TyVeuj
Ek4T6da0Z96ECYVWpuh3VMPxKDJc9w+JPo/Ruo6IcIyNODUI6BSHuvfa9by7eYUy
H2lZgtw7Rfok30SJ1qXFWcHiEbM5F+8m/whHvtA9eD80rg1dbfHUv2ebZryNcgtK
TYsK1Brc95gHigSYXLrPUjIOT99nkWMBzKsNahNisAZKeNMZ1uHN2WgMWTJJehOW
kUhc5ClvEmu9/MwU3CCTFz5vecX01E3PyI4p/0NiK6qgiKjXTY4Ol8Rtv0GVrDUh
HxKW4T8jlheDdTc4Z5pQfNbRr1SRIkN72fD8SwMapDKyzV37jukTucKDFfHrWvPU
oGgqTwuFXhA7cin31naskjusVkLo2PP3nsMdxnfjazVT3iSkd0FcF7zg0HKCkFUy
BJT+c0ZBaXQGaaP4DV41PlYJ+IjiwrTTL2Qs8CA+3eHUP19m4w6DFITNZBd/hcC8
zg1hknLNymnU75e6dphhAcneGOMpDVCF6mBmapv/M4l9IDf22ReDCKdWxBMdl7xB
qh+fgra4SR3GoRgBwVkibZoXnczcMNevTlMF8uVxapmSkzjD9GQdX7MQoGnhyEuO
BQhginWrRIjL00wD71J7ouF3f4fw7hcXUXtTkc8+PuP6ujybRp6qiwNu/yojjgi3
i0wqry8dE5P59giLe09MPxdguqw2ZUI/bG9jmzL3+fOtYXsksCjACvfhiwzmIU9n
+kX10Dj8ke7kg6q9gbYEuMELX3aoSo9mbWyBzuSCSNYyxF0ae9L2lSD1f7A3z03T
HJGzp1aUv8jV0AITTGpsl+3fwbajv9dIzDSatPDGx06lUm+lWQRqTGzIvALwspEQ
UuvERehtJVP0nVJLIOym8K49Y2qs66GELaC98lv8NvwNYfopq9/8fvPYYhFeq6gi
Y9z0HhMmji0WiTmK+onbCCEH88NODCfxGNAHF7KHgt2nab6ARX0UkeJUmQ8ZDH1W
as0SvVzlvS55tHn9qZkTz3gpO8/GLUnV9G2xl2nqpbL36dB7o4E3Rbjfw1c+9sCH
Uo1SxIkAoByGd8cqVf57iuIOvGvxyQvDIKf5q0nrCnhA1UxK22MDSDva+2fvJ08z
Q8fEc7OO2zqWXqxo2WKfE6xYpfpNofnjU8nIu7U7G0hMLTwWNZcq22evZeBFzWmW
sAbHbiDbFr8SRr7ULuglEVOZzUIiCqMUYJRPGAb1ZV4wDTklXhcDZk/aeyB8qKwb
GERfyFRSwdXSCIU5y/5h9GrhA8Cuw1+dHkmulb/r4IXLNGfQqPHF0wmsd7r0iDR1
4PkWOwWP/Co42VkH5FlS2G4aan2ixyK3DpP/n8ly7ZnF09KV9VF7FH/n3tD5p2V+
Vtu+2N6CNAA6ogJjCfNK5cOOG9AwhAjh7tbjmixYX4eEm5MqfaQNW4HE0mm0GjaI
+N2qlJ3RatMSNuEWaL/oXSVW2QxvKekCu+Vd0e54xuZuAGqZRIwKUHe194qYU6Js
1a1V5dYT6oChlcFsbY4Se13SVY9za+z/RVvn7W0/eveAZQkT3KA3Ce51qg1sgu67
WnlnOlfzI9rCYApuk9PysbfyTiA9EEG097GNbR6qwcPv6IYmfCTGfxzc9ONrMOEH
7t+zai0E1KI4bkZ01H76/LcZw3nHNgHCSrfaz6RD1VOzOAu0S3L+VLAiRqEqhiuU
+Mg9XvfimOsWQiagnUITbZErYS9GSVM6KD8xyMcCfklu5Zs8NJDXTUkrr6PKscdH
DGLpfIrVtr7M4aWs44tQMYN6l3VOjB5G5IaP/1ceTvIXwXfsnJysKcP2/nBJg5bN
0IKi7hDBJ1M6EjF9FpNLOZSpDI1QFmfTH9n994hS+++frEst2XSMHEleuj6vuwh4
7hVxtNOv9VAGU/Q+3VSuhwtjiutrAYNP/Y46Zwo7SMeS/SL889qjbBsf8B+XeIRV
gN56QjvxaNIMMhsilZ4uS26tR4LErOc1pxVWEc9dJAJOqJF+Je2v5jtk6M5MqB//
Nu/uHy3p/gL9/H0O+UJXtqOpi1fsG0uZLT2YFfUI7Sfm82SkEGVqvegDCo3uxmGW
TcRA+lgxCA4BWZKw8VU7Y99ZgUaq4ymOrQva900QRGsrh9cR1EJADlJ4M0QMQNaX
s2fVytcd9lHIwayNK25JhgCsGbI6LoBJKpHJ17KjTHhRgB9Yob8aDXCB2XK1LH7y
5p1jE3xNZvXPAriE5GWQ2wn+TkciifzREMZ7INv+KsNI+xpn4YoUENSi9lRdioIj
seOKDeuvYb0J9SfeZ123aBtsGSgRUL1lym9/nQRyP/grAlTbykg3c1/QidGuV4nB
wWyMbOZutJDcy0jn8wGNegWGStkx3CxjY2nYbsCD32TIO/Trzqi/otSsrk1jn8E2
KonCTirdSz8JLlNpUQ7O1VWkhazkRhSx10Z6Whcfr5MrXGZojdgL42Mi5q3G0KUc
0S7YGuSlSAG0DWz924EbWphEdo2wARTMoxiCryBJqy5WUaAR4U5eAEda2fVbyv8W
5ckUk1h526yNoiE/4CnPbLhuoslZ2kUPf7CM6e6LOcSor9I5/pdP7YAjjzHybVYR
WjXxmfjpNcBhICsVV26fNUqBvMr/dpFqz1xbWscVRi7H86oPuQdug5zk4kvEIbWg
Z4zx+0lojSWJf7QivBa9+OTmChOQCnT99hOOuqmQSIH6LM5QVIMivI3J+vmVK93r
OGDMkrA321RCdlL0Nrr4bPklKvAO8U1TaD3UtdzpeHYiwLMAz1EFLNEAhdwpHU0j
BlWCAyhkGn5A7kaeb04LDea1kwjOGgWun4lvVWowwrF7PGzowUJAe1SD9n0n9u2x
ketzZUR/RCIRPqU4TCJ/YGO92HIoOHx5EANqXliJOU6clbLUi5DItJlgvfA7JOPT
fQyDK8DkCvx5NxwNv0O6Fk7T9TdzhILnoHhLlm1RBwOnnWFRu2XZtBTUaYenMf/c
wj4XUgi/cdXrIIFjul8O29DuRbEGO1kYpUn+L4bdwUKBe6YJO59aNALzsV6F3Lke
OyRlWtQUW5r1hVVq/Pk+L/ib0sswjKcuI05QPBhxZxhnTr6yE52O11GFAcCjR2dv
ewHESLuRhfRJ/wlorxerHvjNSUmswQ4XmVOcOW6hdx3PPMaa261Qy9clly5z6ybb
cr9d/P2hnruYxl+bdQ2Wtp3x7KGzri5jkiQnNFsgw8H5LHYPgFsS82vLKWVH73mh
IORuB5YxFWW7+hzxmktHG8z5ak6Sb0fjqRo6z8ILMB/Oc2y8gKZdP2s0RC8tHgsB
EfFwsmR1Jz0npu/W5yfypZc47fJD9F4MEXX9wrneF+dQVBOVWcjchGZwZzqZmhei
IItBTQzX/Uf/HsAH5cY0FvQAiJ0PYL7xBCfkVI71MProXcesK70vcXqDe46xPuNt
PD1AsylGCwwu2GZkaHhK/Nda/GEfvc+QrBC1uoMD3xaC0Nj+F65vWX2lEIuv0x+5
qr90zNaoo4KEaKY5tkqAXWfTOiT9vXGxpAPbns4XwIMGHXotxZ1zDRXZxHArk3hF
fVggAlRz5e+d7BddSZyQuSA3Svb6lr7HtwBHOVpXfEQA0ZgjACKQ8Fjq3P5ZRZd8
wr/4oG/0QiSlrALZ0Wvr9tX3kIdlJMN1/11uzwz0WpBODThRXTI3Dug6k7b4J8SY
HLvhJiuROUKTq/xtgqe9nbE6IITkFxytg+pEZI9Wu8WK27siC+gWQrz+cPB3A+hI
CL9Uma2vDSpg1HcjqD7rq2HwqBLVafp1ooxR0+2lNVRU32FnWFFqrkkAUixNjRW/
3rZeAbggvvAGde/8DgK/CyR5A9iuXpxzcksZ4jip5OihCgNSB4LE/RJxAApWxCXI
+y3dVzM9zOyWOw8l5w4g/sShoWaMr7W8k2i2ltwBNxmwUuEy4N85VOyUtJFy+bCp
WUGo0ObClqIPuaxmoDqQrrIUph/VEffqlkNhm9Fkt++hLqRUe+Tv43+k+GyCd9FH
j/tEB9BiEHEHFm/us4CjxMBONad6MOKQKsRQrwKH+uSuhsDw58tuUJZBhtwRQUU1
aoHDHAJTBp1ar2qXZqXe143HUrdtr41LeUyA8zcJBQmbdLxcqaQsaZCGJygXXnRV
4W65cKkLziZkH7R/3+DC3NB5UdoCGWqJKgIPxH4fr859up7qHMAq1fIMRN3QE3d2
rFQofZ4BJCulc67O+4GINjU95vG4YOY6VrLQ8veJTwMkHdasFErWV8uMNKygqDIT
57kPld3LwTLkXdCmT4dcgg6QkPJHsYwOFwSLTx74FfT2pv/8JfVnZFejdDYLAPgo
kncwDuQHyd5SPVvdRwPKhaYl0fF4An8afshLw/ppC0ihAJz0/35XOn6ZRdN3WTxF
7vVoZ1RyyBs4NXVT5Izq061kk0H1+hgy1gSWV3dOnIVV9QarCb9860n9sozB0pYL
8j721u+4IhaQ50Mc9o8bF4nERWFup5MYAq76/mKJJU4zZL9dYjaKT9m+xb2IbkCJ
aQG50kip3hU3OmV352lFetvSdr/dqv7a2z8408g8M0Y03V6tG7wU6cPVeiBBxmfn
PVYi1l7wRwDGbvJy463V+ydwIQ8SS9zp+XgL/y17hC0wh/leeDps39LdMM1egXHz
BGJF8HALzC6EkvkRjZtFAjmTWoXGadp34eKYaSnyWfTtW8laTfaE+aQQd7RZY4JU
skUw7hefM+2tM//CIrotoVG9Opfyvrm4JSvqKTYDnXlXJmh061bOCntOJcjZAUYK
J5Kmps40r1twID/ojse9glO6hn2vpLqSrUrOrV+KA0IxnMqbzI+tGkdnmeOX5zYC
cwPtHzzWHNuoVJVgsMTA69fmY0/ObwV7ZIp0S3f/9KtE2rz4BT0YTLoSEeiNC+DU
W/CKrVWhMP3YIg/n120sw7eaKypEMgnkUzsCZxEq2SQzqAV2YKy4dtKeWm3+tdre
rG+6uf/81Fq03DB4Z2hOA4MP9bo0ujU/jN5caeZIlfmb3p+t5IoqWIyPU/44eLS/
dT9Hsyg4h53nGHAzajyVoisDAleh0h6y6QEYvkBgDHciByM1eb6XGLzhZmGP3xRR
RAgTHKZSu8Ddr/JEEN9Q5jh952iGRn73W/tR9TrVZQk4HCozkkJBN1oG3NqBWN5A
BiDOR8iQUsFcbUpGKJhfSxR7xtB+x97cqW8hhK8sbx9TSeghFgS3dDWTZkIpkFWI
Xjgp/bwsLwbu6P90TcYzgOSjOeXiWaBXa0u0fUg4BGjik01cEKhdv8ceD9LOi0Jn
ko3Q9oKh8lE6M+tMJBSCthmAbK8OjKni8dyWCcUYCjSPlFp7bNXEeKmu+WBo3gu2
3wKBJ7lZ6SrDimOU/txmbjvl02wM4p3k620sce6/G4/QH+IThkDKbhqypS1gBcuw
GXPjvOZj5Qf7rGxCPawQ8klxSRUKvt6RKAK0e3uymExYnS408Jd1PFPKhmo/8Z/7
Q+Npgym/GXaAisXcFXZQA7w8MymgudAKvfYf33pnJE2iqUzKcqd27gRFDL7rAB5d
aDX3iARSiB0oAXDJJOTkvOicNVc1v4OGE9iBEA+mQC8RXlWD0Wg/+24sEcHIvbFg
VetMYpDoq/AlLu40dtcT7fe49DLq89/Rr0Y4V7tdNP4wym0DsEq7PlLn859ocQfI
6J/9JITN4X5hfhq/jx9mcr31hmPN+trYPWWFaAIOIOZSLlMdrwDHD/MKdgTxHpAS
pFMTqrkx7ZnnWqX5Kfo+UpG71v85sDmZ67v3bxG4xktYU9pRRvz+DFBuJBPVB79W
VBcvo4XRxGRcKxalTqyhTNUt4xlUBzzzoHy0FrJr0KwvPx37yLtU6xQFIhOEfUpw
/kBSRaLCeeRGPfV1tRcNhBZz6nzKYaesY4zH9rrDhlxfk52eBdbG3/IZTLl6CJMh
FNg2yhguwl2YLQeWa6XnPdN6+JCMRahQwjUVcSbjU9nIQ4Np1QqilRfPYhZ1ffeM
9Gjyk41/nmib5VcMurUUeF1re7pehD1H2BZeAMp5dm77VQ2sSd+o3vBaKwlRdDiG
YR6GrMAU0yEkpn4aXNoG0w9ilK4VjwfclwG9rpzb5QWWqAe0CdgcKpYOOsKdM8Gy
omXF8F8PxxMM4UreqOmGPH8ji3VBFk3/xm/iGr6ZDgZDpNNE+JFp2NscSTsUZ4uT
xBAf37PSBWcbZx15684v8rTEY1vCzoSkNJzt8prmfxnks3ylqn/yAaxvnqe8Yz+f
nF46xPgWIw/Vsn4rUGz+18lZBMQnuPu1axRkpB5lmkacdO7nUUyClEuPoSn3M3UD
UboxfyMs04sPPTPMwb/QJPw8PVi4xufEvhOVAVV16BpIFQgMq0T85WRDAPaNBT5q
SWEcqcXxA3QwMb0uUFdUAv0okoaDPR5NHjVEMtV1pGJHwjC289581mkkHu36iqJZ
aEBMquaFl7zBqbJmzGQ1OL9taq+D6LkBShe6ZE7YR/b9A+HU28V9utgydUCqcTLW
BSfWy5enSZ0A+Q0xhq3daI0yW3xdGGavn4wEPwXkvPi6MYUUFP873FOwI9xz2G+F
je8pxTsWxRRoXEYDnK2MSUw1vUPhNHud/zEOdKZ/abuOiokR9VLF08rTjsKLko1X
nZYWw3G9ZawCh8DGfHnT4I7JKB/qjplMGRCLAIFhv3IezzH8pxMsx214fWTF1Lzw
T02cQltbkctCuyOZLQsJY3eK+JFJ9sEjWn9nKz14UDW5RsFxAlIytFGD5tLtBJuv
0Sk3mEzW39rhiaLbiH+NfkFAHeQDz3dUaZlUZQtsA8XHpYjdIL3YmkSJbs89EOMa
lBezZMwEjzN38ysZgwjtNMyERYxioycVKGTucvoomVrPkKx4UaZuKHhL2qkTDeYT
ffoPtLKacisYUYrGyca1/bz8ZYp2TDKzgorFkd6YYUWyKTaqO7zTOY/rxY9GtpPB
n02t6n2i3JX42vNQpAfjU49fXV2rOx8ZIg+XH5jOFjEniA/W3WtMVRZSk8lkq2WA
/jnVxKcHN05DuMg0SNGOZTnO+21a2w7FbI3yXrAxEAQT/FsCvmrdCaENe4ymn20w
ENfLIESl3+XhKRXG8h5rdUBJ3ttC32RhJC8HWBYgTcbpUzu/IL6Jrg/kCQUS1Ita
mmfUGguTDR7UocM8AZAvrxNfr/Dy5Vb60phxdt77GNyhi9i4gm6iff9APg03ZusM
O8rVHOUvJ2i6fptmxb7kfPpny3U7BK0Qny6I8drkbCKcuT7I8rabr089PqQ23rYx
jgksguH/zYLIrTfFKS44JWWFe+hrHGkFPgUlEYGdqbe3ae+VaP0mmzS5EuLr3Vv6
CEQKlVoOKMw3cv6a643t++6d9Hvv1FiIM1+uqKgPYyl2F3rhlezTsN9qk16K76Dd
bCgiF+5+hqeTUeATVzqTIsUY7AOcA9TKv8RJyowfuW6hrknCDQi8SdpyWzPo4QCI
JbGUXrp6XYaGpU9u5MweAeWaeG/IiHhqLa9grlW6MAPki+aCyPtdr+Zde/v8RyYT
WivE3HLGQX3papy+VwnjAKEgLSnLFXMh5UAS4mBdaqKwfDqTQwCEoF1NJ675WwCH
p74jaGikBamlLqPaHCjNyXKOcFInuJhzn3qnLJjxs7RkL/rrvG5+Fq0FepM5OIu6
ZLK/ayeSliLb3TCysRpD/XyPxmS1clgBtNw33Wl3Kxv8n8lXD/3lK2Y09CCCSK5s
8FXiqsLjFg0sqpu2rUIAji8CIGl3b8J3yVQ7EDkSzB+D6PzXJ4ZX8mXgPRE4/tqr
6ifBxgv1QJov/5Pa9OcCuCWNB5WzR1pHvgu1ERtNNniWOhwr4ba8pFvmwXDZD5OO
BFWF+BKRa6KYh3dliGc/UGpg46wn/zMedVySTbL09KYoxubLYQHBdFhTt4kfHZYh
mUKOhWszQLjPViWDgULWPaUgqFjtGPEp+6r3vtcsAS3/T0A3gjSevdQXhdxoFDzE
yNZhdjjxANwbi4ikRtSkxoIlhhIZrDYSAy+vc6vNlc/BhXqu3EIeanvnvW00OCuZ
bNjMaeFsMz4Jo1GO/9ULczYUtsnkdJw2zOfnEsfs9Ya10sW+gOdjc3zAmbOL8E54
lCP/3v9pIXZ4uIne0WUGqzFrmNC8VjeBWkRIrSuPInJxd2gbv99OKUTDpcp2zwlK
fFlsOSF0hDEhOGUEQ7ZZnywA/MjQW2BW+yiVal6EweBRWKYau5a0hRG+/RQMoRLC
U1vp72AfYU7nRkrux6mJo3h/4m0acxDw70XgiLWcvzMcG30K5BjC/IZPDW30mxex
mjrXgsxUIiZwVxRkullD3etc4TwXqYKt0eu9vQKi7FN4GMdBRcrWFT/JqA1S/gQ3
dY9VH0n1RZ60hk6AGFM416ziu04QybtGgMxhiZMq/3YPEnFdXyllBI3ccfTRvEFR
t0mtq8cz+HLYn8NoGDCIg7arnsO2NYXxXO+RDk3ZjbNhxeKzdEoZjZQwBjn78Qiq
MGPCmQ2HeuYWuDeMqQKpaBULB+RV4GwedOwHQLu/H09fKAVJfO35j86vDRi8fSrf
evGXkcWpSflRPk8q6IfKoiDk3WGnOn+21Xom4pzbXa+Rb7KGtAPU9Hmi3ZCFCf5Q
1CLFWH/atszw1OjQa/DkBB6mh2tXbvQLV+BCmApLCWlvlJSjNtwyyY9wCuSQHq/u
/M9P9T4B1/IgIBOu4OX7ItHxYqBlTHViWp5QYOW+gN9R3DeOHe3swAgeVHaC6FA9
d4RuHGx29EhLpPRlPzCWFqo8ljpGDJ5qOlrE2w6str7emCPRIcXEH5EutLrNi4Kx
aovTQ3G60nRuoAL232MPQcmy8JdydYqsnrsKa95DtjGITeAayDEIIc+LzxpOWjSm
OR3FsH3HMvRTBP8/Rs2E/Xq9eQ+AklXPZ2YWPCDaK8UpBJVLCy3S3vU5yWwJgeFd
NqkqzZP3cHIa4Q+xUTK8RY133H6H+DZFteSDKVNu6Uv/fajE9nnWR9qNraPjt90O
bmnmfhAE0KoHqe4pQqWZYGUzHSI4riXdHjdSkmFtE6fnSk2BQmgE9Emd8yfYi02P
8ix0n7Ac4tz4wfpXHQwmuuZ7SChIghPaCzA3cP6+FdO/Z5+x+faAjCNf2IEWcPJY
rLBrZ+r3KwAfd/v0AEfpbQQQjwWJt4+FeiZgIsNux//5IeEs3ixHumo3B3W2xASJ
InVpPNN1nG58wLA/GPx0vNGFnDjSzhyYyEWXr0L0A9JVqFeV01UI69Q1MsTcoIvI
YpNSFf01Rc0x/jyyVd5RfyhFzrtlejBbJssPAMh0SqXNeqRxXBfjQEoTD1GeW74r
T/Gh4ugjQoc7IOUX/i8k6lso+zjjzILjWuNr+JVlczlBURbykOQnpiJZU4STEdOr
MmNH4Evn1E62VOsbWrrEnUomMKuk5bRCjKcRNcYmWkvbWlvznMut9VSGBTT8eaGX
V3som/p/gEVH1e/niQfIqQkxNkmzCfrv0KjuEf/LmsCVehx//06rDG0RO3gN1Wgs
3ulGyBPOAo8teaghCt/d+h/l+lIccsEwgivkK7fhBEHhW6wvZIrjhAERIDVcit7Q
uPINo4G02SL84bmab7ikrQL9esGYg2z55ETASY9smKCL1Xu9UakPaBgy5AdJyit9
CCWgstqMvUYb65yx5HB5sXQT7pmZGipCY9b60HGplIbViJ68njRZHNJYPLs7zk0b
7tL0Xb6iVyCbYt0FZNMoBNfHJuJ+wePCElLod/D2GyDAZKC10u602A++GYqYh6Ry
OQum6cXDCLyWblKhl6WLDfZ9hwHjKbiaO07v1dY+RW4d8Ki6ebXHmYoNn0rr4vEz
rRJrSXLGbxYpfesSkZdo1MQQWy95LwCJpK/2uQOrF3KEzxnzbUklQwc7Ci14uSCf
CgxDY9mWfTc19kjmNHv+xlnsCyg8xcK8PfpvnfcClcFSM6oBHpKS3npxL1fX0GHa
Sn3VUUYjJC6aLPAf5upy5zQ8f1ZeXMZ1BwEMSZ5OVE1ctm8W09lfXl2LLCFGIavH
OkDia152xJqqaYppyoKvo1aiTjdLWQx07ggM+mwDoP3IG7lfC7CuZrtpcFZi6hI5
hJ4Uh9+Bot3MJLGQcIyd55w3bRr99KMv4RXK1Ogw67gzMjMTaYqMhYqk/xjvw9UD
3aI7XTq+PdQwoT8HsXSuISIyC+UOtPgrXCJeXTQoCJZUh7+8aOXhcdxD9Wrl7pWL
9hHKJn9K8Z6hLwx2jD08BvirAvTAJIIyp/dG9l6AyNmwIixBtHdXPqxBg+rmvb6g
7iJkyR8ZaFvP69L3ACJehhG7+1rHXxqL174VjrlQDVe4NhGIlTMG69EcMIKQqoKM
NdIZNhj9sEJxbN+cDRqPNFuokotyOCdGR5Pc/c7cYP7vYwy3P0KGP8jpJxhKjSli
aAYyvqEhN+NtM98ShbGNbLK7IS/ypVzfzoZywurtJ+Wy+ILm+odeGtHxh20w+1tn
QaZV3t62ZCQs/I4wIsPUoqvbnylc4gW83Z4sO1+Rp4ISB7ZkivZR4gwT74oVYQPc
vC9rPOoIaZPbtqjgpZnuU1Ir1jaA5+EaosgRTOg0hcX+ZzsYEET2sZIbzaqTieh9
+WPIw+R4at23xsExZRwXx7f7SSgi5/iInp9emFCIhjlO2F4EUSRugQvCcxwpKi0y
rkSSe1OI0ru1qkBnEDzp/AN+n1z7CVIIeaWXOygUCUItq9jhMBE4VfSqyIn/6fds
rkj30aRLwMBsSuI3nZaSzD9fwHbT+iGGXSMoqObp0J9FHHO83bHGsqAT1osjt0ZT
HR4S1XZHMZ5pKoIibfTsDDAqyY+G6+Qo4m+o8TkVwGMeH4CHPBjaRGoV8cWyAB6H
yD/Zd2GRTlgn9zStQfRq3heiZKtsFF77MzvjUjJpooCO2bfQo+TuP3Pxqp2OFlwC
PeokQPxAlvBNdV5/llrHwc3dqtfMol/uN7H51EwjrwIdXlg0ixx6Z40xYgRYHxeB
qNy2VnYk0d1eb2RPjzbD5A1CxlxosXCTzDLklALmDqJ+w6/mTA5mWY+98iZvobrm
MpodZML1SiK3onk2QpiuJNHCIuN13vkNaGTm5fZESpd9gv8WxFaVI5Lp6HM5riB5
5L83Loi/KxU/qSzx+deRjPERfj4L54lw3U1IKC8qH7R4rzNtujxAqCvwYg3c3A2C
yRZmyY2nv/o5gtMtinmYZTe8VR5laMshJNtiPGramjplhdI2KvTDCDSzkh/58g3J
HuJ73401Ja9ljyPyxCzN0bl75l1KNN2Zre0gym0Gp7bWzEDJUC0ArTA1K3auBCpp
5LSaXbGpbEqDO7ihD0MJGo0Iu2pewuYa0uaiWewcRONSFsb4/hycmoAko7f2QWz0
7B/kcMAbbldclTYklyMEZSZHaEXr1KhoJm93AyqiOVW7bVuGe43zVxqEhhiEvhO5
03pr39N6lEDgPx86PGc8m0zWPRNDUyebEwSNa2T5m6eqfw3NxBNznTXGRo6WFqxg
gwgPIee1Sj4AkQ2SyBaULvDucooic8kkMzd88XT8vsmd/nStlgryaS7yK8bj6XJG
Z4ZR/7tu9hC4FQIUSQ29BDp3U8hvAh2J68hEAG7nWnHNHwyOU9otPdxzZbf7gDZj
mAVdHe+pI7geqynUyVsVEd15TT/7r+aiVi29K3guqVhO2QU/9ctiAunQ0guov1bL
zWUXa56A0o0exf0cnfdA4DUiyxlzYPnFPAxP+v6uR0l7QwZlSRvCB/EjedzwzGDU
YVxRwajG4OaC7RFk2AYiV12avI0VJLu/Mg/Qgx0JhQ3xowCLTfiuVZgB086oPUgR
2fqs75yYPLbye/+0/gHqCEcsBdD3d8IWmwxN+vUbxnpfF1bo5MtQlEdLmCtFOy6D
LKDvfvMno+C80BDLyaw6sR+euNOMRVnCeA1Ya/+d2dAcV89zOR+hiYt61aTXaqYS
ATYtw29IK6J4WipYhHNbJ0YNy/S7lG+g3yE5I9pyrmvbxSC2KPUy7S/ol/iXdd1a
q1ohZxHjUU0ghtTIEzgueN9AWlxsqqszshqv8ZhCWQp1Bdr33xc05iJk65oHQmaz
5g2lMReyIBGmxLfD+OvW07nhx3cB5oeGoClgsVRXdDvR/ifcaFkr0EIejPbtDkJg
M/rTBRWxnbXj2WJLg0pOEYGLmS8Obv7aN1dpYPTg59S4UVzKNsVqbzo8IrulP02Z
E1dO+EI+ky7mjmDYxW9VDiVwEvuk/SKhw8ck7JgJaE63gz3qHrTD9b37JF2HyD8c
a8wV3itnEAr2I97CEWWCREV1oszeCJX1G/uoPjQXlceb9mal1NLlcC7zoQF6mhr5
mjPkVrxmj6+HbzOIo65HwpwFS6bxFa2Rk952Nl3gLxLZ1Al3EXqvNUdhE1LNyUWI
xkp/d9p1zSGH0iIaZgFOnrzIWiffebVz2DUGoqqXPE5U/q4wgzD7mBeeHemANICN
cOkRPkTwZ7m23tHoY/fIEJjHyD3cDEbqX7d7OmgzMQgEYCqOE52ulrPDhpph+vo3
h7Ph5drGS2TrrDyLbpwxyPRSz3LzhBlC8ixifu8rKQ7K28SmzmLOekyXDIrL888X
I1l/R8U2smrB4yN1YjMGNB/E+9ljcJibZtoI0Y8OwJbvR+sZmoEmRyUc7ByiP86d
IoHL5EokX7mgdp9t0tMjlb0xexzcp4IzSaEP2fHvmaGG7n9elrrT69ieiOoDW40N
Ae1FejxO0h4L8smCqHOQslfumiaSTx4dwGIuky29aG/7h6Y0fa1twIqhllpYeklm
NAm5HSpwsf1nQ42AZg3yEyFhOTEm4AkeREgjg37zkoNS+jbrQnYBWzfp+hdu8YS2
u88wDNpK9Vqxxkoi7dzuoDchGw/Tu4RkoR6BMnhhMQ+MGxLBDQUyqSMXq5m8bAiF
2vdJYlvJ5ahG+ez6QcEM13gifgy2d4kVuhyVZgZhvPTKevpupgf/XeITOIhF47UF
O1sWMtHkhFickfcuKWhZ0DAjAjoFip3Twyd81ImixP+Q/458mT/JZrJkcMAQwh7O
1eHyMwvsxLSLvE+E21pZLi+0K2bbcuOYXc9WculBQ2JY5TTZvlivzlYRHoq2+/ed
KgcqdCEVjXGLrzZPwNpOTbZtQflFjqbhHrYy3Zv2vrdqt/1bqBAxpLm2a0u3aU7D
/dWy/eGTGn2SflvokLB+TmhzhTvZ98+KpWV1XuGjNkjytE0cU+Dam8bnKSMEvdCo
7TWXivPe5+uBK0N+zUqf/bENNtPsRdGkthPCYzOqd3af9F1HVfyYnUGsKFWVAmkf
+btaQPAIFqIBxGFZHLC9kXP9vAR5spy6c5v57KfCFZec5cpThzr+OcwOG6O2LKjy
wI8rbSj1pEP1Odqf9maBdUD64VsGY35/Lu6+EZ7Zark0lJzFihDG6QeBFnqDbWYf
rNWVv9TQaWEuXV1pRcniF+uifR2gJmTrdSYM593/z5fcaPItRU9IpPmbK6UUdAs7
o5YmPIPvhsB4NQ6HX6ZczEiErD/8JNWz27X8tIh+KgalrfeJzsSk1k1SmtuXx4lP
rs8ZUqDb8xPzPZSKMytWj/Jq6w5scSqco77QG57m6chYvd/ArFdZATpRs18HTQeH
FKm+vD+J6gGlVxGY22gNC6Y1mm3PsjRd8KeRYblOvWMB8xr5my/Bh6tXfvvnmk3a
QpyRiyFhYeEgoVLJO9LMvXBAMib2H9GitnZ57ybit9V6TMgEqoEjwupm8Y0dn4rO
8ILGzFdtGRD2u3w/r8J3TRy9bh9P9Ay2pWW50Lv0kO/CfGGNb3QRdjOZP75FweDL
h/3bIwdb6Bb+MfT9rniSHZtJ5ppavmUgRYEnOBan6+PSQfkowPcNeOoHIDec6tVZ
M8XNEuDWXeLA3xbks/EBPDMhAmcWVxQ3PYASKfJ0/DFpnOJjgpMR7RZL0f1CyWfv
8EeZIdOvB8SElcqWfBHwFa7gqYXnbQHPCMB7H1HXVxz65gqt2eHUB27KX9NZh+zu
PldcOTDovT/5xeaREN0MWLXPGkz1mddYBXdxcaIGa0lBaioEQvfdZiRFTVI4P5Y6
7yaaQ+IRqRiNhm4rqHq/WFOqxZJIfwdv3Dhw159HCa6cNf1GHp3lye6bvtYpdUBd
12fhff0YEmMzMzDHh9hYn2suEz4ipoagn+gTlAzUW/zBkJNqR+BQomJg4GjoQWbm
kFvZuVqJc+EG1EFMsxNmzA7r05XNZF0nthR3DdAoAlkd3XTt2uUXwX4n++YsvVBA
Gx246OPRZPbvrotFZQN/Y0drL2S/D4pfYnEbN3TJ9Fkoafb6jLNJ2mQC21nQysBL
4B14MXee216prSqpRCuuP32b2B2XBH+MP7oR3mj2uIbEmZC8ACrnPjrL+7FUcblF
FsJ3tKPcIIOfnwC0x2XZfr2YsTEZa9BtD45vkbF/UhBUUOWIB0IBa+FAtnAtyooU
sgHYqTou5yfiVx6rmCI+/FmyLkYAzfmyTalXE7M40T/rf5qZlxbxzEg0XKN9ORQm
PWTDkY6VcmmT0lPUywmbAadU31yFKxjM8AMzL9utdk8aof0xuuNszxkRuYgNXQ+3
vj/1wj2wZ6LqA/Q/OtnPMRYvppblB76mZKZwJs5JTTf9/4uNVhETS0J/lJglqJBf
LTR8Mp2KnrlrNpTpIAlpSL7T3lgo0bSPsxPZ/E8nN35QA+Pb2iezxTdZnFTebBrS
wosdbktQlYRHT+FNiEL5zDIxaQZvBt1WygQtCpqjwbNn5kx9U2fW8ABgMt2LXaqC
OX3BKyD8JLKqIQ5/z342xjz8QprTWOUqq7c3nNz/MPXt3c5EpbL0ClyqvAGUVCcA
PTPqIHwnJhBWBVQOfMNwwH/NoWMNqPI4VfjM4vUgYRucNn3T8gP/S0lET7F3hglU
+yUTmkC9kk5TEEhBC0R2OmSlQO6/c80HDKg43C746OXQnBldiSqnZzC0SU+vW2J+
3R3+JhUaHCwRnTGJQaLL7eBiWXUlijo/JHZ2V9mxTEyExGUBrcQHYttfEU73ngjz
9ry5WL+C3KiMYSpPO9zNe1H/lb2Y8t7C1VZLP9SMYoUvo4DW9OVj+y+O4Qy/rO8f
vm3bQbZym8eLYeEaZAQKRhIKRVrmz8TvDLfY1xmJO5FP+lG6vS9uCBEgaD5K5hcy
n6ODMN0dVPyJrh9Dw+ZQoiiRKGleWyDyveuAw/AYNy1YYb/oZ2+HXUDqBxv2BgkY
kdBzZNhAe3QhsaF1eRkmuTesz4NQb7HKaEBN3CrcOpu2lZRnOuqF3yAwIbqStWM1
EhNePksLjJLI39Jq0ITuZiexrXSIN039HxPWBAcuDyqJy3kAvGa/GtWUJJOl8SwK
M+UpDrZ7SOkUeeQJE9Mmfh3dvuSOU8oPOM/NBszh+PVHesaBnE/38Xmd4H8bZKfR
ftcrXng9Urfc7yagt/jtYYFhm5IK0g9SeNfUU2S6eYaVQ9nousvlm4zfUFwskLik
Gon3diwqzEXRYidhtaHceXmoznyozMIwSKaPaJu1OQoU31/HnaQBpsIx21DANJuW
GWXw2QbeZ+5GYEZYVt6X6OE7OI386iSF0O+xpUhcsKsYw4yiggl1WWrJL186jJVE
R8sBRMzTHeDduj5lVMb+IknB5EgCNAUsOeAawZY1DComF7U+V4Vz/puHgVEF7aKn
I3SxLUMrjvy6kbtPTWG4HUP57VPstfIxx5mtV0tc6WqEZbNXxjAFD9aBfQaQTM3C
yeW7iiX59a/ZjSSWi12NVOcjbRJSV5342/N8td2EK2ktx/XM+jz7YCVRoeOnBOVL
NMBcp8IsnwJz4kPyesj3YO2MD3pAQy4Gk6AOb2xP3oS+GAj7s5SdmujXIWSv+EGb
AiTSFSH1yY1/fiLhVuZuk9sxtFnKf6pvVsl/gaRqHgHYXAJmFOEQpng/ax/sIHS5
nzR4TxpXLXE2JiMpxH0Twrd1gGASRJ7fgPa3K3QClX+vfDvD87lS1QE7PskVqSCm
ZSxf+6Vquxfc4gusQ3B/LnlD/UlfajuJTYRdl9YDyaMmgANWI7ZVqIks3d0UgAf9
Xf31knu6hiN0zDZ5t/jidgYEqmT+5K5RdKgx7w+GY1lgEnc07/69hQQK6QSR6b+M
WxBQj5RKFr5ChSVKLg1SIg1qo/RU8ELUuuQrjfT1SZmwLF7/an7FCyOpsKLDc7jJ
WLESQnZ36N4IaGdNlZSSzS3o9qgJR6/KmOhIM0l8xJrtZR0HTZTeGr9SVfqRYEZN
sUsoGtVchbXi+xuqPmvL78j+29b27Dzbs1NLgSCLxpNqQ4ea2D5qTqO8kee/AHNF
smyzcD0izvbqdcUrMS2ID4nQNq+5oHA5mpUY22+2TFAK4R6aAGCNrFZD6sSKsl8K
ot6wm5ywQTqM9G5KxCBA9Dw0AJ6z0Yh3HciS4fqzUyMpm2xUGB3KAzwYST1gUY4M
x/I5PkZfXF/2ZBWoYOK+05I4jlDE9vv4Kff4Lss9dGI8UtjR6/Bzm3gSDqCD5H41
Zv97Ve6B3VM77JBmIQ7kq62RhNdOanNnYv3P5C4UjiSg+Jv0Xz9F9JxnM12Ek5cq
JVAYnXtZjUAdbo6eMuEOqWvP4agHaWUTYKOpF7fqXqCQvNQOWL9Ti0ONbIqmL2xH
RygEy0cEQYbuKF4rXeEGHUOFEFyyacJxE16svi0MpQ4RjGfNHhGKifQVRBVzIzn5
kBpRWl8XdzQYy10kvKAhpXNiE5ZH97TZEmcMuEgRZCHo3feACy6twX4cmHHCbRbk
QlPGqX7ZoGwswX1xuYIQu2XZFzwyqm1lBU8YoHfqMstByqOtSxLBw7qaQdYG0fqZ
CyTIztGI27luD4+8dWyD2Ihc0YJqOu7moUssOUDJMLmiWQOlPtb3CKIQU21wFfXf
d8v1V61Ffg0hqYECAdCq0dBNvcVuc6W9D24tY9J/V9y98QnLTwxIXKHjbw8m/wpU
X3cMB0WUIZtkiYBLHxVdK6LMdd5l3x7ubm4VR5iHY/+WGHQEhSFz/4loiL9wzcaP
ZECI28DmmQfpDk/3p1TP7N+gM7S1OdyFCxLjVgKu70VP3lOjsrEinDx8pGEMUOeh
j8B6Sc47OpCr03yqzW4+ufMsvmmyPQZ3o4kGBf009Qs/SArAoeoVDrYGvGnHLhVr
wWFLChch1pKkPNuI+miQqat0Tz7B42097GlSN4eCPcTUVLZ1uem2EzLen68ZhyrB
M13zaejLCtMl95q6lCc7z+AthMvmEMKz0vm3bTzyXmk/wOd0mlPlSvjtU5pe+GJE
SqFLDvEn47GSnojxEpxl/DrDS5IfJPjP3OD0TIFAPp341N/HwAModWjGFefxHBuZ
CEuZRsGfIAjF9FgVt3f7FCu0Qc1BAGYgwjM180ZqbXGG9ideyTFRjhL5W8bCVpzi
4L/LjQiNPurduREhf8rPTATaWpwx080ZA4HyqW4iAli0349qQ7NXTCjG7T+uPr+Z
APCsYa3BXzVshxkmEQa50JIWW90dux+a7ZFMHFSRveCXrnMW30rkVs4+PKDPkJHR
t8LfynWSBeeqSSv0bmX2Pn5ThyrvmYK7yVh/pZXT4pv4JtRL1GjZcXoCHwblHzYg
Fyd5WBykBiwEAlhk4d4dE1TN2zt9qx30Ns2zH1kfNLw6iUcADrqfrwoYP/5pz5pK
1j7g9EYxMZghOlfElmK35jZIqe2NPJyEWqaKASCCvFSR85ajTvbX3VL2RVZ+SmKb
wAHyWu/HfO9SrPJP2ZyzTlICGL1W7W/xnjssQ9qNjiWUq8IaEcc7zowQ5KckoxxB
RW8iFBK/dES2/NFrgq7xFnR8597nFAOCSSGAasOG4s47eaZUeQhogIqgwKyI9ghb
LY17UOXsP4TSP6A2qCfe6ElZ9EcuI+1Zsle42CieV1vMTSpav7vXWJO4UbV6k2sT
nwuW/AmUHOMQ3I47XV0oBpbKx0Sd4h7hWJlppIH9Al7wa/d/CEO+3UD12ZTmKZGu
2+6jPVK77BYchIw5ulIykNXGNZv5jBRXaT2f6eSuR7tDZnVB8ZQuqlvxVKwQ+vCX
AIzCbvOE8QiFPcsIQKHHrftrAAGMzpDZt7dY6ivWT47nreyQMWn4QawL7U2IGIWw
x5a2LbowZNy5M8hmNKEwlpLq94X0bcC9uho7BEJ0+WnEZmoNqPGp0VK5NnQnhYhx
w4BprZfotDpN7/d1JdyEGJBmUHt7MLtGOaN3JzZbcQE+tljwptk8RZflA0s0mK+M
z5JEwKQTcHCUvpm/MUk3QZpj8ToEawBGBdiQxy6KrgPPkNszCCzT238DDs/PAn/q
lx/Zhr76tp5Fal/E9h74ujZy1GSUiZpICsK/Fq0F6RZ8MQKDYXitCGynAl180BEt
kf2pocTfZgWGUAkRzKO4lS4t+0Oi9AuJGDsTgUZOgEAO4umc9OvUL7b/HdLu97sS
83FzA3wARwBB7r+BgrNdO0nSc66TQVFcYlhTrmKkNdPEgeb+d8aXQFfUizd4AJhV
CtvN4yaEVnw1vpwWOZo8A1ZjDD2XrHTTB7pvR35K7rL1Lpqi3QOKQnzxmRUcNJFw
idv15Yf+F/Ra+XVAN3Gn2T37+RXs9sXhq5mQWAH5zMLIlb9Dag5vN28Bu+1MyNua
hVy3J4jI6X7pzxhhBWM+Y65SM6sELGOSF1E/8+MF3ezwMI1i3wZxFCmJ9Zf8QKt5
uRvxZnbCOjxAV69waHFMvNa5hQ7COyInPhKIYedsYXifixoQfeWBZp0yaMZJb2SW
zQT+CFUWfV1ykaN68TjSgJsYmPHWyUmGQ8Ig3TgupVn1qNvzIhVW7nBE0KO8/RrH
hBJlzjhonXoFe9N2NIp1jv/QYVMWM0JXKT9VaStAlAawPKVzUkWPOhYlN0SMf7ds
o3jW3gfp5KhsujzfMTIVcjPnFkkaokCeG1frbIMyRgA74+tynnsjpeXCeapffhFW
ilOA8woomXaAVT5zplxZ2OoGKqYWL+GZE+PsWfjmqCnKXN1CpOXBb4tm/3O6/FKi
SsArgxi6/yiy1vDR+o0GnPzxxqYfN0jIxzQlq8/JGibJxXhq/1wdI97vgDtCGJLq
MCQVrNuith1uqysWWl1Nd3mh+tMOTi6v3FHLQEFWoSB6pxPAaV6hRAY6+B9qkBqz
kjkHsW/soy77lK1/lywlTM6PF1freNBwv9tpziMll5GblTObUa7NiAOHh0IQUUeu
IY5lbERvEfdHdiEw3lBwyhNbhKAgbeEaJnPgmQvz7EmVguIHlfHVCG6bEIBYqX6H
mAoQYB7kDFSPGj1kxU+KeZLvsg2x09rqg5QNwmPx46LfZEPkuKbtQfYQG2COMPiO
oGosGXxs4g8rFt5S0HfIHI9DmnwRBD6JREQEMFEOHkQd4d3mVEzbnAI/6E2evI9C
`pragma protect end_protected

`endif //GUARD_SVT_AHB_SYSTEM_CONFIGURATION_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
UgaaTpGxvlZUxetkX5VB2ELYpCrazrmKkF6Eob9duirLObXFCdeq2Ts8UsZrqEjN
lrcw8WLCm3tWVXACYEf490LtvP9pGkFi/F0pplBc/5xE9T13Yd2asKTURHb+wR+Q
4qIVj0o/HxxFkxAU1feUeMHV2uINzCFrYj+Jtlc5oXg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 156836    )
lwDP2ZSKjMjJ4sXRuDMzt9cJXsgET2f3OIoAXHLMCw5YVAWgSuo0ntTaPDhi7/0U
Hez3nFs8M3VzNnQNFI0/r53UOh2wJ/ph1uKarfzzrUrdfSKrn9K81xBdB6E+ypk5
`pragma protect end_protected
