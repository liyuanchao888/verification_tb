
`ifndef GUARD_SVT_AXI_TLM_GP_SEQUENCE_COLLECTION_SV
`define GUARD_SVT_AXI_TLM_GP_SEQUENCE_COLLECTION_SV
/** 
 * This sequence generates UVM TLM Generic Payload Transactions.
 * A WRITE transaction is followed by a READ transaction to the same address. 
 * At the end of the READ transaction we check that the contents of the READ
 * transaction are same as the WRITE transaction 
 */
class svt_axi_tlm_generic_payload_sequence extends svt_sequence#(uvm_tlm_generic_payload);
  /** Number of Transactions in a sequence. */
  rand int unsigned sequence_length = 10;

  /** Constrain the sequence length to a reasonable value */
  constraint reasonable_sequence_length {
    sequence_length == 10;
  }

  `uvm_declare_p_sequencer(svt_axi_tlm_generic_payload_sequencer)

  `uvm_object_utils_begin(svt_axi_tlm_generic_payload_sequence)
    `uvm_field_int(sequence_length, `SVT_XVM_ALL_ON)
  `uvm_object_utils_end

  extern function new(string name="svt_axi_tlm_generic_payload_sequence");

  virtual task pre_body();
    raise_phase_objection();
  endtask

  virtual task body();
    bit status;
    uvm_tlm_generic_payload write_gp_item, read_gp_item;
    `SVT_XVM(event_pool) ev_pool;
    `SVT_XVM(event) end_ev; 
    `svt_xvm_debug("body", {"Executing ", (is_item() ? "item " : "sequence "), get_name(), " (", get_type_name(), ")"});
    /** Gets the user provided sequence_length. */
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(m_sequencer, get_type_name(), "sequence_length", sequence_length);
`else
    status = m_sequencer.get_config_int({get_type_name(), ".sequence_length"}, sequence_length);
`endif
    `svt_xvm_debug("body", $sformatf("sequence_length is 'd%0d as a result of %0s.", sequence_length, status ? "the config DB" : "randomization"));

    for (int i=0; i < sequence_length; i++) begin
       
       `svt_xvm_debug("body", $sformatf("generating tlm generic sequence 'd%0d",i));
        `ifndef SVT_UVM_1800_2_2017_OR_HIGHER
       		`uvm_do_with(req,
          { 
            req.m_length             <= 1024;
            req.m_data.size()        == req.m_length;
            req.m_byte_enable_length == m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] inside {8'h00, 8'hFF}; }
            req.m_streaming_width    == req.m_length;
            req.m_command            == UVM_TLM_WRITE_COMMAND;
            //req.m_address[11:8]      <= 'hB;  // 4k address block
            req.m_address[11:8]      inside {'hF,'hA};  // with and without 4k address boundary crossing
          })
       	`else
       		`uvm_do(req,,,
          { 
            req.m_length             <= 1024;
            req.m_data.size()        == req.m_length;
            req.m_byte_enable_length == m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] inside {8'h00, 8'hFF}; }
            req.m_streaming_width    == req.m_length;
            req.m_command            == UVM_TLM_WRITE_COMMAND;
            //req.m_address[11:8]      <= 'hB;  // 4k address block
            req.m_address[11:8]      inside {'hF,'hA};  // with and without 4k address boundary crossing
          })
        `endif
       write_gp_item = req;
       `svt_xvm_debug("body", $sformatf("waiting for response of tlm write generic sequence 'd%0d",i));
       get_response(rsp);
       `svt_xvm_debug("body", $sformatf("Response of tlm write generic sequence 'd%0d received:\n%s",i,rsp.sprint()));
       `ifndef SVT_UVM_1800_2_2017_OR_HIGHER
       		`uvm_do_with(req,
          { 
            req.m_length             == write_gp_item.m_length;
            req.m_data.size()        == write_gp_item.m_length;
            req.m_byte_enable_length == write_gp_item.m_byte_enable_length;
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] == write_gp_item.m_byte_enable[i]; }
            req.m_streaming_width    == 0;
            req.m_command            == UVM_TLM_READ_COMMAND;
            req.m_address            == write_gp_item.m_address;
          })
       	`else 
       		`uvm_do(req,,,
          { 
            req.m_length             == write_gp_item.m_length;
            req.m_data.size()        == write_gp_item.m_length;
            req.m_byte_enable_length == write_gp_item.m_byte_enable_length;
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] == write_gp_item.m_byte_enable[i]; }
            req.m_streaming_width    == 0;
            req.m_command            == UVM_TLM_READ_COMMAND;
            req.m_address            == write_gp_item.m_address;
          })
       	`endif
       read_gp_item = req;
       `svt_xvm_debug("body", $sformatf("waiting for response of tlm read generic sequence 'd%0d",i));
       get_response(rsp);
       `svt_xvm_debug("body", $sformatf("Response of tlm read generic sequence 'd%0d received:\n%s",i,rsp.sprint()));
        `svt_xvm_debug("body", $sformatf("calling end_event.wait_trigger"));
        ev_pool= read_gp_item.get_event_pool();
        end_ev = ev_pool.get("end"); 
        end_ev.wait_on(); //this never unblocks
        `svt_xvm_debug("body", $sformatf("tlm gp xact ended"));
       if (
            (write_gp_item.m_response_status == UVM_TLM_OK_RESPONSE) &&
            (read_gp_item.m_response_status == UVM_TLM_OK_RESPONSE) &&
            ((write_gp_item.m_streaming_width == 0) || (write_gp_item.m_streaming_width == write_gp_item.m_length))
          ) begin
         foreach (write_gp_item.m_data[j]) begin
           if ((write_gp_item.m_byte_enable[j] == 8'hFF) && (write_gp_item.m_data[j] != read_gp_item.m_data[j])) begin
             `svt_xvm_error("body", $sformatf("m_data['d%0d] does not match between WRITE and READ transactions for sequence 'd%0d with address 'h%0x. write_gp_item.m_data = 'h%0x. read_gp_item.m_data = 'h%0x\n",
                            j,i,write_gp_item.m_address,write_gp_item.m_data[j],read_gp_item.m_data[j])); 
           end 
         end
       end
    end

  endtask: body

  virtual task post_body();
    drop_phase_objection();
  endtask

  virtual function bit is_applicable(svt_configuration cfg);
    return 0;
  endfunction : is_applicable
endclass: svt_axi_tlm_generic_payload_sequence

/** 
 * This sequence generates UVM TLM Generic Payload Transactions.
 * A WRITE transaction is followed by a READ transaction to the same address. 
 * At the end constraints and write and read data is compared are checked at the PV slave side
 */
class svt_axi_tlm_generic_payload_pv_sequence extends svt_sequence#(uvm_tlm_generic_payload);
  /** Number of Transactions in a sequence. */
  rand int unsigned sequence_length = 10;

  /** Constrain the sequence length to a reasonable value */
  constraint reasonable_sequence_length {
    sequence_length == 10;
  }

  `uvm_declare_p_sequencer(svt_axi_tlm_generic_payload_sequencer)

  `uvm_object_utils_begin(svt_axi_tlm_generic_payload_pv_sequence)
    `uvm_field_int(sequence_length, `SVT_XVM_ALL_ON)
  `uvm_object_utils_end

  function new(string name="svt_axi_tlm_generic_payload_pv_sequence");
    super.new(name);
  endfunction

  virtual task pre_body();
    raise_phase_objection();
  endtask

  virtual task body();
    bit status;
    uvm_tlm_generic_payload write_gp_item, read_gp_item;
    `svt_xvm_debug("body", {"Executing ", (is_item() ? "item " : "sequence "), get_name(), " (", get_type_name(), ")"});
    /** Gets the user provided sequence_length. */
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(m_sequencer, get_type_name(), "sequence_length", sequence_length);
`else
    status = m_sequencer.get_config_int({get_type_name(), ".sequence_length"}, sequence_length);
`endif
    `svt_xvm_debug("body", $sformatf("sequence_length is 'd%0d as a result of %0s.", sequence_length, status ? "the config DB" : "randomization"));

    for (int i=0; i < sequence_length; i++) begin
       
       `svt_xvm_debug("body", $sformatf("generating tlm generic sequence 'd%0d",i));
      `ifndef SVT_UVM_1800_2_2017_OR_HIGHER
       	`uvm_do_with(req,
          { 
            req.m_length             <= 1024;
            req.m_data.size()        == req.m_length;
            req.m_byte_enable_length <= m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            req.m_streaming_width    == req.m_length;
            req.m_command            == UVM_TLM_WRITE_COMMAND;
            req.m_address[11:8]      inside {'hF,'hA};  // with and without 4k address boundary crossing
          })
      `else 
      	`uvm_do(req,,,
          { 
            req.m_length             <= 1024;
            req.m_data.size()        == req.m_length;
            req.m_byte_enable_length <= m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            req.m_streaming_width    == req.m_length;
            req.m_command            == UVM_TLM_WRITE_COMMAND;
            req.m_address[11:8]      inside {'hF,'hA};  // with and without 4k address boundary crossing
          })
      `endif
       write_gp_item = req;
       `svt_xvm_debug("body", $sformatf("waiting for response of tlm write generic sequence 'd%0d",i));
       get_response(rsp);
       `svt_xvm_debug("body", $sformatf("Response of tlm write generic sequence 'd%0d received:\n%s",i,rsp.sprint()));
      `ifndef SVT_UVM_1800_2_2017_OR_HIGHER
       	`uvm_do_with(req,
          { 
            req.m_length             == write_gp_item.m_length;
            req.m_data.size()        == write_gp_item.m_length;
            req.m_byte_enable_length == write_gp_item.m_byte_enable_length;
            req.m_byte_enable.size() == m_byte_enable_length;
            req.m_streaming_width    == 0;
            req.m_command            == UVM_TLM_READ_COMMAND;
            req.m_address            == write_gp_item.m_address;
          })
      `else
      	`uvm_do(req,,,
          { 
            req.m_length             == write_gp_item.m_length;
            req.m_data.size()        == write_gp_item.m_length;
            req.m_byte_enable_length == write_gp_item.m_byte_enable_length;
            req.m_byte_enable.size() == m_byte_enable_length;
            req.m_streaming_width    == 0;
            req.m_command            == UVM_TLM_READ_COMMAND;
            req.m_address            == write_gp_item.m_address;
          }) 
      `endif 	
       read_gp_item = req;
       `svt_xvm_debug("body", $sformatf("waiting for response of tlm read generic sequence 'd%0d",i));
       get_response(rsp);
       `svt_xvm_debug("body", $sformatf("Response of tlm read generic sequence 'd%0d received:\n%s",i,rsp.sprint()));
    end

  endtask: body

  virtual task post_body();
    drop_phase_objection();
  endtask

  virtual function bit is_applicable(svt_configuration cfg);
    return 0;
  endfunction : is_applicable
endclass: svt_axi_tlm_generic_payload_pv_sequence

/** @cond PRIVATE */
/** 
 * This sequence executes the UVM TLM Generic Payload Transaction in its ~m_gp~ property
 * and returns once the response has been received.
 * 
 * The GP instance is not randomized before being sent to the sequencer.
 */
class svt_axi_directed_tlm_generic_payload_sequence extends svt_sequence#(uvm_tlm_generic_payload);

  /** The GP transaction (optionally annotated with a svt_amba_pv_extension) to execute */
  uvm_tlm_generic_payload m_gp;

  `uvm_declare_p_sequencer(svt_axi_tlm_generic_payload_sequencer)

  `uvm_object_utils_begin(svt_axi_directed_tlm_generic_payload_sequence)
    `uvm_field_object(m_gp, `SVT_XVM_ALL_ON)
  `uvm_object_utils_end

  extern function new(string name="svt_axi_directed_tlm_generic_payload_sequence");

  virtual task pre_body();
    raise_phase_objection();
  endtask

  virtual task body();
    `uvm_send(m_gp);
    get_response(rsp);
  endtask: body

  virtual task post_body();
    drop_phase_objection();
  endtask

  virtual function bit is_applicable(svt_configuration cfg);
    return 0;
  endfunction : is_applicable
endclass: svt_axi_directed_tlm_generic_payload_sequence

/** 
 * This sequence converts TLM GP transactions into AXI transaction(s) and sends
 * them out on the driver. The sequence gets TLM GP transactions from the
 * tlm_gp_seq_item_port.
 * 
 * If the GP does not have a svt_amba_pv_extension extension,
 * each AXI transaction has the following properties:
 * burst_size == data_width
 * burst_type == INCR
 * atomic_type == NORMAL
 * except for the first and last transactions; intermediate transactions have max burst length (16).
 * IDs of all AXI transactions corresponding to a GP are the same
 * Other properties are random and can be controlled by the user through a factory.
 */
class svt_axi_tlm_gp_to_axi_sequence extends svt_axi_master_base_sequence;

  `uvm_declare_p_sequencer(svt_axi_master_sequencer)

  `uvm_object_utils_begin(svt_axi_tlm_gp_to_axi_sequence)
  `uvm_object_utils_end

  extern function new(string name="svt_axi_tlm_gp_to_axi_sequence");

  extern virtual task body();

`protected
2U-S-/<T0AK7.\(J=)&a?,gX,4X+Qa_HYRG)QT?CI=V@U@(fc=3d2)T</bT>3ZX=
7WYVF<)8B9>L^]R-Y:/;V1N?>NR[=Fe2;GTgAMVFKB6P4PXX4ICD>?L_Qf1]@7)6
1d@8Z99BVZU>e8,1]R<0X_].)C#I^aIWe\EeM<cSA^W[2Se6K[MeEAa^P9.T_I.@
e2\#-YC-0_Sf_F)-EB#CL\^:\/G7:9L9+CGRd_Z/^=4BU4G+O+ME-[RN#FWP=HJ2
&WDI^\3SBR2@G)ZI5a6M5H0e>K[:LM;M?-(YR(,8V]XaS=.,-()95]\f0ZI(f74Y
W+UP8:OK#O,WLc_2e4N3N]gMJRLD?TT5&A+:GPF(^YJ)DRT&J17=-;Hb<SgPD[Nd
dbI13B8PRF[_FA;PNfJ[3UP[/K::cY=2/b@8<A8#[BX5BYgL70^16+7DI;/(BD3]
/S2f>YQE\#\_^dLV&42.c?#TR:3U:[<d6S(;37QdW?BU&EOP;:C];T)6c7/BJNg#
=6Yc6KcfN<9)M.gec@J;B(;6B:3O\a+HS(=5F=?UKY74IIHD/Ye@f\4^MC_HL/)JV$
`endprotected


endclass: svt_axi_tlm_gp_to_axi_sequence

/**
  * Reactive sequence which translates a snoop transaction into a corresponding
  * AMPA-PV extended TLM Generic Payload transaction and forwards it via
  * the b_snoop socket for fulfilment by an AMBA-PV master.
  * The response returned by the socket is then sent back to the driver.
  * 
  * Automatically configured as the run_phase default sequence for every instance of
  * the svt_axi_master_snoop_sequencer if the use_pv_socket property in the port configuration is TRUE.
  */  
class svt_axi_ace_snoop_request_to_tlm_gp_sequence extends svt_axi_master_snoop_base_sequence;

  extern function new(string name="svt_axi_ace_snoop_request_to_tlm_gp_sequence");

  `uvm_declare_p_sequencer(svt_axi_master_snoop_sequencer)

  `uvm_object_utils(svt_axi_ace_snoop_request_to_tlm_gp_sequence)

  extern virtual task body();

`protected
eaYdf4eG>?@A8-3XJHGR?_6f]T?#>)UL#<N95S@(BgV#VMBM^??c7)N@I.._WWd,
b-5Ha6+B.=NbA?4U:<R94G:Ke=2?5UgX3S0=,66Ga[<N0HJ=-CET5Z2bE//;KICg
R33#1(f.e9d(7gVL9ROTL^[&NIabPS9/(Z3Y7DQ_+FL^L@,;MeU7f;fND(5S.B.7
&6=\&d5a,=^:^g=]aV1R\e;KV76BIMZ&D[\Hc4DA<<(eFYQaW=,a+9>B:Se]bZ)3
c8b-S@L?Bb)S&>]J+3M8KD:Y)9\?8,A9IAJ/:;A@c]FS?g>B&42PN^fRSQQaIHXR
QM-)D4UE[(^X1aS3:eY_F>,@FEHSL)8-6HVMG7>b)7SLT[JK7[E.+3SLS2^O^\3<
VdN;AJYgSg<UR-a?fPJ8D5-IN:3N_7-KPW@YMP?Wc9SM;,::_,:JPRgYa,+?E3fF
g[@ZVV>35E7,=5+f9KBg6a>R3@-<OE7dgbd\0T]aB@W\M.W?-eFc1e74Jbb5CH^F
g->KN\Wba5@2(UXGfV.U8V^[&^70H\3bfBP1L,d:Od5c&&K=P,Xca<74P$
`endprotected

                                 
endclass: svt_axi_ace_snoop_request_to_tlm_gp_sequence

/** @endcond */

`protected
+BPA(\=RT&(UZBO-QANgN<QE0+Ngf8dMJQ+R2HZNAKNDYEegFC\Z3)PAO]&g/\=O
E-.Y9VAFJ,GI[CK;@TKW^#&MC]ZIRf7K\L\a8F.b?.Y_>[0b(aEPHTSa#^6QM87a
LE+L1-QY8Ec2cOB4e(G<L=O,_N?VMP=0&R^7P\O+EH7[8KJN1c_BM-9g]3P585/^
g6OS>M&+&Lc/^WCF9[U#&&7(3&_CGMMaJ^ad):6M5,Z8?Ib1dRFc-N+D^7UZ\c,<
+SQ(cW5_Q70HKY_)GJ:aRRB;GGAW6Jag&M;^fK.3KHDAZ6L<J<3Z\0eNZfU@e&H^
2^LD+>/,)K3-bL-NZ.Z/:<4cWE5D/_:SbaKKJE8DX9:Z-RJ8;7-,a2/5PQZ/e@T/
S44\BFNW0XI-WSc9U17)e9CRbDa7g9>];VZfMdA2>d.2Q?(,)IMMIQg#Y&F1BZ)a
F(1Na[dXI3:=(1-aF?WQQFAga#BJ)KWfNL?Na&a^^ME/ccE^[Ke,TdBH11EB.ec,
+g6>17^9cU./eET1e@I,/W;](61a6fg8[BS5\2(4&[cZJQB<UE[-<;;Q6aV9KNDF
Q8EE?Y>W.>.-gB9,G:aCO(3@&3:8=6]3V+ZDLg9=UdJ:3e6Z@aYJ=HVDLAE/\8gN
0;FY2+f-.\W2?C6H]9#cCfB1e,7L(<Aa8gP/O3D4dNe[EI0I=2Ua0E.g2&T0HMR.
4#9.b#)C)8:Q\ITYQad.68D-Y/E&+=VJ=2KH8KcE,EQP73^E)?,(EPC[1ALV2=37
3A[256gZ+8f>_I3W69FH&#3JCV[2N;-PUY+H0W,:89-7b:+ENQTO,S]a(PT<A=G?
Y]=QJ@W,V[S,ENb,H/,3bW<TZM;:(L1#WeVM^gD1&&A?^1<7VEI54BS=6c+)]CFe
CHfZ-2NNK=KH0c)M.IN]+Gd7c)DKTAQ8T:O80)6c1BZ=)][F6,KBB9Y+fRLd((:a
V2AJf>B48g6(76E2:57FA:9TM7)dQGKC&ab8#L;gb8T9)R@T,)]JYfP17(b(=FA0
(GN,M]44;;gTgLWD=JF<+5^1P>FSXP&5P_,/ALe#U(b]8b@DEWB7X_2JX@<LJ=CL
.@VeUR[&ZF..PG#?dZ[#?&?9:>I:R(GUB<,Y9R5O?L2dC=#WY_#EB[.RB@])1f4R
,,]eO#QTeg0fB&OJ82^J;=+I+BPKK1:3[gF3-P\@HW+Q>gIM/TK\&2WFQVE6Ug6b
,Eg^#6g5\dTdD<0ZO?eU72e+4F4P<>4b(2F9^ZcSNXP0<GI]AI).N>f(Q\T#W<>g
bgFcVNXI/DH72:LRT[[L)])NDTA_@1L0WS?^UeaT9&S_58&dCaJf]-#fcTMULKFA
HQY<PGT[5[3W62TL^-YYGD[D;6e3\Z>CVORg(PCceULgZ17?BAeA=KA@B8O?dA?/
(HA)X(9]_1G9&X);6&Z.^<AZKX]8?fS[L=GL>&ESBfb\-Z0:H.&L]5MD34YH1WSL
B.,B:X+Q::K>=gUFB0@>2,4[:b?6ZdO&==Jca1fY\,D:IRFP@dV/48UBIDg69GO-
X7@KMdH]dY>P].F87)M2O@Q1F=fbGIY3>U1gNbHG^dFSV(O&GZbHfJ>9H7R.X/K,
LF+a3Z?A&]:#E=M:T\N^\-5;U]B_G;G7HS1[4ZAI)C/_f7&;C+:D]3^WX8HZ2d8Y
0aJ-N??\3[G0@FN]:Xg@_RaYRFTbC<G5.98/eNbN>Z\/XN;e:d#-F3N(1&_?Z-?G
bP]KQJ,UNdA25P[,,\5]+fC=8MA@20211RK@c;&,U6E#,:=V:DVI=D]J4,8@JS96
+8G8M]TK(09bQX=6A1#TcaU37?88U58?[M?=T]c(dOg>))dQ,V&HccC[>#:5ETU5
126S9B0>)MC5/Re1Mb,De5&QA1GWIZF/&b.FL89,0^O_K<?=LLY692U:cY^KA>C9
G4ae.M6bD^_Xf..#8Pg(_]R&4Z\c4<850JC[T/cWSAZOeV86LTXC4gMaCdQ7J._9
<ZS&J]7->LBUYWFM/YD@\a^-][I9XK/dBL,G/<a8U-M(XNJ_M)UbN]I^:Q+9RB:>
Q)6WI_[/6-Ka0Q:55WFRZ+#5;]S@9;B8SS<T_bM#eRQYg-NX-MRFDI?YN(N>L+SX
1HT.>.N8-#W>X?RC?CTb=8+d[YT#(7aP2]fSKbV3?4O8DYX&OC_AEg&/]R^fVPK?
FBdT1aK[<#<MPUWUKM+I/[_NDX<]VcUa<MTT89Vbe.OfOF62=>7\9WV/IU5;7Ra=
O-C8X&Q8X_gWc(?^/U=R523cVSNKfGZ3V5:K03dRb?YIebHC8D4W.fCN1O1HPR=N
\XSc=LDI04GX5@Q@#ca<\\9=G_E_C=e<4<eL?/7B/6CBc:/9CHE9WHNLQ03KSTdf
g5XODRMYQB1+E&34MHJ;/@[QD@I&4VNf11?.AO\J@4.6HL_.TU3JJfgACWM[KH_.
92J1+b?eeQ_ZY1BE)J5A)L1bga-0PafVNe=7LQA[=]XUB35bCbJaZ[.8QP;<;de>
-+\]=??7_A/4Sa^6)FRb[MSVLJ[gQH@Q]f.AOD\FOV0eBY(8I1eY1:F/GM,Y#?GU
3>D1,T5(2Z&6eER(-?_[d[=\Dd^4YECJ^>Ce6f^F8#F)=,W)I?N<7dbb>+Z#AGIF
Q@3YJJ3VddG]&(,ORH9<bQ]7.)1O6N=2eFRcgXR7-D2BQDeQ7[(#Q_F2/#X(^RdS
1Se_/Zga0GeWQ6=<O9),&,H=/eP4=9KMCd\V4#1a=:K7J6;E_TE:_3TC&/&)TKbJ
dN>MTb+HW4Q2;7LHF1_2,T<D8<H@KHg;?aJ2HGIA.P\/RPN,8<^U3IR5[FT_9NcK
3.]AceTZ+,.fff^bGXc>VACM]V1Xe,a28()eP6e?1U><^3aMd5,B56WS_)Uf\\56
F_[WJ8DX&XD.9#1-QbC^KUKW]JN@aK8DaJ1YQf>WQ0d\Z>5/S&aS1Q_W;gDZYG\f
YZKT\.-2Y721L@+X#8BN-4TX01a801@>-bO<U-T873d[:gNHKY>#N)cV,OE;YM,[
4e9NdO<.>-2(NgU2-gA-R+>SQ5E85M<33+8T:J5GJPe6+/\O)?H^L-Q[]MTY7&1\
9NU86L_g08egC3Q./K146XECJM-3S-69DdGO\2F6:@#SLEJ7,#6V3AWJ9[^F(7X^
.+GWCfMFUgBR[U?&1OaTQFJga_&FfQ:f#JNEP9cOeQU-2ZYF3G>OZd0I<#<cH-PZ
GF#,CcF(M-9,0=(E[EW^Ag638+4.W7[AXJeER1(a7L.Z<8ce;NcA60bAQ>AU^?Q3
1V9>_IOX0;)Y@#R.DHX&Yg&E#_J;SI/N):@H^)KM565O#>^6;d-JXSF)?&W[9.Sd
eW#K;@F2D)>S=/MQ.\5aa&-NHAG&(8/>gdZ3RVFV(RNIYSJIJI6BJ^DXcJ#LI?#]
;(FQeBO;Y7ZQ;fW0A6;IZ3BZZ#:a8718K;_^aVJ.96cI[Q:0.3f1APO#86\71NJV
&UT<J#ODT/PE?ADgYNP3bZ,,#2)NE32RZ:>URI[LQSG?\M:UI_LS+^2..C@R_V0e
#Qc_D6\NOP8QMeTXRK:E-dS6GRa7HgdK:PS\X;I4#J@H.M\&=&I</NY58]::;]68
_K@g5/./S([[,f7MA2dAM9L(fdCXS;G/8S;UFg5e+3BCL2?]TN^):PAO#9ZI[Q;:
)><8d0WE7MJF,9BZSUE6Q,9Zb&3_7OV)&^T@=<f@\7I^WYV5)Z12[.b]\T=-EY?\
,-4R>D?G>+)_=\(G0^8@W@[#8NZF/J^fb^QYa>X<(P:^0EPR[H0d>98ITKB4.4+1
+J.>CaK[/4-[cD5-GPTHQOPV#JHMf_[84A3&\W4,I(b6C>18HLda1WH,89F.VO7:
I-_-a..LTCCLA5Q^Vd.EUaAV?>d8Y\.Ff^\2ETW6>I/[0I>2T,bB3P\EKKIQ9Z7S
=[[5,)-CKMBTfBV/.f(b=HEDKB_]Z6W-/[EHQ:C)A<4fT>;K);>/+@[UHc[GZR0W
\eQGeZQ0,LA1>/V.8:=V\6LP&09MM#XXL2-aWEPA^D/HgZ_78J>]d_A;:/b[L\b=
EQV5(dRGJM>1EG\\.32I-[V1cf(,LZ^<5E=;M#cBS]Q.3QUZXRP#MT[J9-?C>4XX
(gRUISHccCMKBPNDbEacdP9SWHFH3HY9->2@dPGD(34XT<(D1\cSJK7]TYcFP7fc
)D,X-+eF5I.Ed8V@:5NPcL&4WaQ&NAM6e_A9,&]gf3aY(F5+;6AQ.:J+O/4b1ERD
V:/aD0dR=O_L?9<^@_I3R]&H8;;ZT<C,W:6/Gf@X2?M<PYe4(LH_eI(Q[6?Y+?)f
Tc?g11R]ZX+aB\<UOAG^8X1+K]eP)70/Yd8(Xc(R2L9-f?_X:6Xd:B,?C79:Fc8(
]Z\56bWZ(SC30&(/Z6;B<^\BMFN\]FIcAfH6?e>5.Y[?([E&Q_P>^1G6b46-7&J(
DXT#)8@93?I9D^f_9aEabRI8&M>H66-\EIJeEeYNV.NAY8BAE^L\Ka0,:EG.F]bM
\.ZDD_?O.<9PNa6X6W:=SLf=O9S,.76b8Td<-INc1Xd(FGb0+4VG7JJ:?LVO.@6P
1/100)ID=H.GNFgX\7REOWAZ-ZOgTZMG6aEb>U&[6NMFNZO7dRMJD-<<RO[dMRB2
eHYI;\abZOc8g5S_2\7;d5d2+WCC;#G>H,Z2-D0]C7YY262ASWYE7G4-P&7^M_G=
c_,9EfFHD+.1ad@B-MLZ,A4XLFTX;1?dSIXDba0F,8J,@[RCbd0OTLbDI+fe7ZKX
g:A)X6C;eBTCO/8@]4>?<bDcccYK>T0A2_;JcHgH9^_+aO-0&=2\2ZSOGG(_EE&L
FT,<J9#1^1HDI=[&,f62:Cd+c63?C]Y6Ga4WXfW=8W_]19Egcg^I4=V7JVP@(#g@
3.e8IM7:/4E+:>@Ba6^63BZ\]f;dB+M=a-(.X+d>@NbM4=<[gR2F+3dBLO4T&Fg8
/2Z-aR#Z&Y5)2&,BTR@NFd+;RX?0YJ+HLM2P#=\70dFQBX[EU5=cf5SH:gWCeA;T
L-(;A#SE#8T3GZ\ZW^]T],X7NWTd4f7M[L&UdCMHbOWAHM=?,YBN(MIa2g]7JTcg
]T,>C(T,N1eY^L2.gB?#Tg-.4YS<GX?R2=[4W;I(/^M4@&B34C=cD+cPeE,)-12=
#N4^PI#Z:,Z^NC-)FMH(cTBc8:/<[;d>f)-0E(/L)BWE]YQ5WFDO[;7I(O^eb^W3
CeO>P.8QS74<gZU0R<TO=20HQM)g[F#2:=-1DLa,[.I(9g.8cV=C)9QDJWA3,813
_=RC&,4:fG\)@BOSY^\<Ae&IN[,XF,6FRWCBN2^Q:#:3Ib:a>90>?/E&KA-VSF3M
KFFIR7,_Q@)bf/01aZD5X(8\IN@O;<b\4UW=X<;a]dPI:,XgedbV]ABR5W(:9=-L
EGeF/EW8H4YD(GCK(#FPYD^bD)O_&HY3/K:aOP_>Qce52W5_=d[b<15GYP3^9Vf^
Y-aQ5:#;VGR0Ia#K_Vb?7I+F7L,=^bB3W:<5L/_+]GIOJc(V#TbRPaB&Z@(IP_-U
NL[(aWHICQETZ3)cP;S;B#?<@3MM2?5X29eYIVfgVJG5fS:LGNcD+/g:H5MGec1\
?M&J@&U=(JRZg&_&\P\)>KXT0J>.&4CNXBJ.1R;BSB<]080aQG<g.f<6Wd/\F#.H
D\EG)#.#)^@R6FdHHGP]4)-7WI.FJ.;ALQ+eO<)CV2IF/52f&a8Sgf)Lb6_L_-&a
-MIGDBM77@SI]2H4XP\_@7YNKXa2I,<R<IS=4;H:E_D6Z^gDZBK4RR9TWC]/#7>Z
/IK6XOQ@7(3>2FK/(N5@8GOOB\cePYa<(WaF?ZT9Va?UX6_-,)_dRYI&cT]:IP)S
G:M<@<fW;RW4(TXY)RER#82YM3\I0YOENa[-gJVVSY+_U<GC]D2a?ZK<:B:AIc6R
H\#-U9.;44OP&]38B6,NCgHCg:[UV2PWW#.5/>5^MeO4/,M+DbE,^S@41g3cdD+3
VA82T^22Z4^Q8^JYC&-@9BQS?08GWeAb=(XeQaP,\OANG[KM:;a:P_CG9/[@^Z?/
fV?-Rb]SQd=8RZFTG?a@KNS<EgYQY65gQ8[U_)P;LI\>FY>:Q,2+#AaQ#LP1^_E)
L-^H6^3(>+517P;STdZ=eSR)0MDBN3X^1f5P2O(USbN-L),NGKXX9VY8[3d]K?f#
1D6Wgg;0&3b&<#c56HJZ[N8baR7:(f)9KPY#_EZ3XL[4R&,RY9])&_=&-FH1H\bX
bWE;>+MJ[#ZO,A+F-Cc\/5]ARKdR9.@I_PL_8+MW+2O4Y63VYF=;(??a_,[VCD,F
EZHaV)F3[#F[B=9YN#\G>L]=c?AU\)>UCZ;U:Y<g5M0\+TZEJAWJT,BU1dV=B:IG
>g54]0)I]8(6f_T;#01S+I<H1<=9=2HLRWP:gEH4c)g;XL[fF1K7ZfD(7==OfZ]Q
MKWZQNae?/V(Y?UDTIe((INa&#R][c0(Q5.BT/,b_E(.O5KZ)K6)NH#)@_8c@LI5
H?(^-I&^Z=7;A/^2_eG)6gZ:\(P,4W&+KVQC:)2,)9D^5+G=N<5a9=f>GJO=L<V-
3^O?Q47NO;Q0<FIG78JNZX\=7JJ6K:O-)@:F7;DcPeb([AU&CdDQ_.30LG-fdL8G
>OCEU/<d./aNc_W?M>AH@W;\Hf[0FC<P;QYY>7<6+G?e2@g]0T2;R<E^F0^XU,(M
Y4QdIE6H?/&CG46:&d)YfPeDQAJI6>2ZT/Se2g+5_XgV104JTS6<O8KAc[UX0#LK
\e_LF2[EaN5OG=LHg@4AR63=ZMOU7I\>A9g57;;HHb>[.<XX>H]Yb;W1_,&\QW&#
]#FF3#0V6S)Ec&#6Uef)RUAgCH\,-:34L,B>><IG\QUG9=+=-)TZQ6HFPIB/F2/e
>(BCHZ8MSS:HdWZD>B^5YP/YNacf&&AKYUG.F6FXPaW3T)080)EYF/R.#a+DCB]L
dSd&I<<?/O+0HP025,Ofge4bV<BOO.M;a@2#GDNKQ-N(21];\AD10\M-_EadQeXX
B+9@ed?bC9eGSW42/Nf;OacWS2^,>V^:CFg4DLA>P=?[BW2/=KRH:I;:(334X-BZ
?\=OII0S5OZ^RB\f\S.:9I5V\UCMUX>F-EI3T_V#_S]#^,5A6.OURaNNV&3#9M#d
HRNL^@D;E9DPf5OWf\)102fFab<835Eg4@fa5<d:G:P\0TcTdT=?[KFXQF>^gdIP
5FZ=]_]-BXedd_E@2=&V:,95FHcGf\X<;HPZOIW=#K,VaGRHNe\T1,LWa7:=.:\#
+J-5:Y4Q.GR=XE.T=8RNEY9K/g;c+3>6EB^dUI,95R=c=HA)ge)6U-LH=KY5R:UO
+E@GZ]MX8?K\/Q7Bdb?VfJ&\M]2FbCBg^b:.M;;T>,UG_.cIGJgM&FbF47&Q&Mc&
C.T=B@DEZcETRCGa;0&8W@E5TR321P3,-fV1QQI+4Ie#+2LZAeMYV\8L_E5fd1de
YDGQ+B.^3UQ)B;7b@WWVJ:IK58Fg@&HQW@YUO5WHa;AQ0OH^XdG,T#Z(/H#ZIK-O
A?&CZO,83;]gQV^>bf:KBFWM0_(V3=?K2_1K?+0_O+<MW8+8G(BIGS=&\>fO<ZXD
<>4OT6=^NU[/Z79-:<-J^D<0R\Y]U):Kf@^-^gB7C73>XeEbKZ7>J#^-HP)E8,]Q
/NJ5R0@>N+aL.cAaKdbT^4(J;([QXHPA7c<RYN^J?FF@K><?C:UA@=IPX[,<aU/\
LB[U[fJC4(bg0G4+<7SKQDOPX+(8(8)-+e]R;bJKJ<ZQ+)=)fSaWHeIH@(2R=Y&T
?)gNHMB=W&V]LKQRM;S(?1T0.AAB9=DD=CCASR9E@Gc&6DIf;A9AF-JYFSMU/#7G
eI-65KX#&]1\PJ+2IJ_)a\XKReT3.E/cXg(81<:B#3F.7\4=HfTMHXMMSZbf7+1[
bDUY5CH6KTdL@K83ND;4[P3cHKef4RI]YU/PU)37N2PZ5E;bbN9fT+Ecg>O(c>V]
,YaQBBeOY_V#5XO6-X>#(5Ce=-T=WK>0,MQVJ:79-^IL/[Kb6a59OT9@AZ)/Lgc2
:eF<X^6TJ_:<b(Y(F-82+=9@^Rb,@M8&J_Y4U31Of.d^=,Zf(C^@L]3M,.13LedD
FEEL=:69#RB3M(L^9G]5HB&(QL6c:d=23>FD^BK/Ig@\@6Z1.:;gD-fN73W+.[+1
b-eHaSUO9cf/<BB3G+65&&c?.)9Eb;aHL#C&]/A6J\?cPXM7P,P?A:==a)J[VG_,
S/K[,B<bR;@19NH2d?-]GOa<g<B(CE(BCc_][^Z?c_0_UCT^;^V:2<E)36+EJ]]\
-OLUJ-J.EO84CA>82@XRHX>(EBPH\Jd7_bPN)O8RIE[0G=:O6NP7c>NWeI[KQDgK
A)LGJ.DK6>;]WeC5;cRJ5#T=\H;Id=&A4/-Y^X4WN5MU5_K@+IFbNUB_-Y>T<]&9
Fe--\6A/b90f<JR0H+A<?[/K._/ABQ^FKPC>RY;5/bIZ26ZJ3S\EIV=MN8g:TQR)
TVO.53V=3#CU7Xg&JAXCKC>I5RIO#/ee-=+&4MPcE[:87S_A+(1TN-K4E-J:?+E3
2fgb@I-d.DRDc>?))eV(7#+TJ/H=MgV@VK:<cB6UKbTS>0c?c?STJ;8>-ME@HCdE
Tf;eO8_ZX\#8@OH&ZIN?&3OY>6-A416R(9UTJR@\H&7P5X72:,PIOZW&Hg-3>]c_
Y1IU-H)2?^]4]@M]OP8a+]6LUR#T#aLRAZcDJc&/c.<2cJ&f9T\T_EZ=/ZQZUVOe
7S]9P9EZIbFJ[JN/V]?,9^#]H^\[#H[Fe25T]A[[NMe?,F_b6IZ_MULb.Z#WK23J
=99K@f>BH+-51(PROJX0?_EYIIb,J2+#&MgR;c(A(S7LT[^I;JOL98Bg]4_+5X+4
JH<deaZ=d=1<bc&@&(^QQ,B@E?#O)g55?@fAgZMW/dP+56E,5.;3EQX,GMNbT9#f
LJ347FC_.d-c(a<QLI;b7_@>2a]28?3>H]\bJSF+V0^/c74HG:S8/O[^\]0TD5K#
Y1;^=aQNW^0bZ84^?6C5CL5^+Eba+X)fS,MG4USN35AZK8-+-].,T@FXE]H9A-N(
=?E1(Y39+bJZO88d\#CI7#<Y\NL?6cP7PJ@Z?9FSQ4--017U75YG\FM[UCCaVcCN
H(=9cL]LG4:Oa7_-.ZMQ^IF6]QW^AJ^N/CYC<&NDJ[A]NUH#J\X0BX2GF#3?^C&N
I2<I&=G2DY@XZ-.R/:ML]#V6c-5XTJ^_c=-UW?f1:/2g6)Q+4f^XC:Le6B6_&C&Q
e3O6^R^]]\R8C.K1NTHbHgBVDW<8ab;(/I#RWZB]XK.&GIaD4]&8@P\J[DfY0V.P
YJN>RSPL/,,X_Y^PV==0Jd#U9IC0e?gGFDeH96I]3NaXMZM<3agPE2(T]]7U2KUG
a\CDe:EK9S11eTda+342LEbQ9UA.RP6@)DPg8#6NbI8EGTXIQX,-L45(b31,V4JN
E#AWIO;1SR^)6aT]W_XfX7]:8):I+Jd25(2@54YWdd_S^1bWTJg6CY_T[B=gNOaT
eWCHDP3Y\32K2g_#X4PFI]#0,SB1:VdaQTUZG#3WT&#>=,PEZNSg;V&-AOFg/f8(
5V?bYI[ZEY.d)3K1VW0D(DNMFH]3Z<52<S_,SH1/[417,?Y?0L_=3HSa<BM\=A&0
cJ;>&bJH68c?U,TAEac97IQ8U\X_AY;a9IMGMJG@[e_])=5V3<K#+RUVg/DN<;eM
VD?KZNb_eKd@XXAWPT7C\,AEVK:(D4:cT7KOP-W]>U?[gEQ/4(5AD8+;d99e&;[.
L8;+;),;\WS0;D9)NBM-05b.af:Z8PEB(IW(NLV7H89Y-@GY@.@JM-OCO]b&A1Ib
#TW#dKHe\X4+0UcNb-YLG>G^KUJ4)/8;181S=Fe6TQbU7FP[;\SN1]KRMEX:1bga
c<J4&S/R<D:E;QNLa(Fa8RK^L]17fN;W3G]Pc09/g5>cIE7fYBU8gKME,WK=:G0Q
X,0ZP3-]@OeD<LL?8]VP;JYbcdQGce3>A7eAVLB5,dE^BGC4^X::\J))d8DZgP3>
dGE2_Y1G;Ddb^<A1>_RC3>e5(N>FRX_.(FS3PU+M]4b]b&)A73aK5R14T0);=.Ue
:_3_MLgaLgE148a>TROWICA)NeQd\GM3D2gdV[BE@Z?9ZaN[YH8_J1-@(B6&R9Ud
E>]N2:KcZ26L/,\P3U+DE<?e]GR;2#Z(g.Zc@@c+\@9W9eFCT;fO#ZMgM,_He/Vd
g&bH.Z)dM<5b5(/\+a=\/Q.]/8LA1[fZ[O#JA-7H=)1GJEL@e5TIMHI7DRQ[a?OF
3#1Z39;R66^=4OQ]2df],eg@/g0e0JDH5<FdH<:1C-U=gMf8?(+b<=MS9G[;?&\,
+9W=If.I0++QXZ,X9#e5]+=g5R8[I5A+&7-0bdC)VcRX>(:\SdAG89Z#_ecKc[^f
;g4Q(9_JXg3]RcA7E6gd;>L]Xf^O(E-N2\7D=4U[NU=S4WD4RUUU[1-6,7>M)@cG
;g\[^3YDY,?f-7+F+^]YQeVS0NUD9[G+#cA<-@ZG3,H/?G/c()<#[gXYB@6?4X2e
PSX\,GaK)<cJ:J=<eX7QT-,gSJ/H4K)UK[03E__ZLX3Y,SOME>K=MCOD7+;YBg?/
K\ELD(c<Zf,2Y]>@\VVgIW:IL3:<EdRQg]d54P.EQbM)AcX0C/d>N8I0B^WRP^-Z
:&-OdIMEWT]O]\g&KSGV;Y3VY/@>Kb2/g]&SOZ_+G<A+:0aLe)E+E5EVZ\JJ67f]
S]TceRCP()LCS#^(+PWbZN[+TZ;DJU=I)FXfY17+]:=(g1OQ()3125bc/JQ0/6+1
/6VZ82TH-3NAg+5MVWC\&XfUB[3XQ=JZP.J>B9NfBY]cK+-\<d437=GTS)-#&X=3
A.AfSCPa\g3.4,Mbf\QTHX7/[VQG/&4-/cRKT1U>R=Q+\^F1:<MC]?KHB]G,6_B)
P>>)XPYK?2KKBTV.L5+>361d&9O7IACAKZN4YGKf1ZDKgFRSF)S9([LPfA:KI2/b
HT.59@c3ICL;La(WJC8U>HOceL6aUDWV+,G##\-4#2?0H5^:ZT#D)PT<g;g^T.;7
d4F<VW)-e>4N6b\Q&P\9ebLG4fK1DCUYY=0(,16(d63I^f#5V;S0CM,<:dQ;,WH;
cBP4T7eRd6O1Td6&7D+c4UE6?XQ4Qf@f]MTM7_AaJ?\6_1>5Se6YP7_[]cWH:QAM
VR<0BVBcNK?2CEKPaM8732)7RSTLN;^D1Z,IL:G0eD,KX4Ef4^[&6AOEO#5R1dSB
-.A[\HK./OJaF2>f9M;UOO(W,(C8_Y&_CR:8D&?QbO3#DP62HKMJf@-9N\,c=8FE
c[YE73?<EIW&AEW;D/2B:Oa-REBb^FE;aF;?VDPM_cX]>F?H28&0?.W_E\F/XbL<
ZY0&G(-a-#2/EHOQfP\4cbP6KPHZW9,_0D[,/3UT2[=aLNY,b<R.N)(R74\3798Z
\2/@+b/0,#>-C)UC1Je?7BI(CSE37G][g@G>H@TE.1WJ)Nc/\J4JK]6CWV8>SVCH
Ea.OJH&<)@CfR,e1XYFLd_TRMf;YV]=(K,VM8+X]>?g4G-g]&Q?^2HOBc9bY[8S&
6d0:\+AJX+.4C+XObH?>/OQ+^Q+OA1J47Oe<T-W/1+2#U5\-FK@[3:bTF14;Y[^L
7PU_)[g&N&WceN1VX1@gX@J@=T_)#3\\\5\[?OUQ4FX341I-5<.@VTI+GEc),\Pe
LV(V:#T+&R:K9OB+J,^9<G.&5](WIPdG2ECTXa^F17P>]Cb@IP&)H60G+2VB13&@
+TD]#RVLa=8?,,a3cG314L3^8bF[GF9FBWECa\)g\+=#[(6P(H3_+[Pf3>EV&0(W
26:W05V?NH7^QKK3gWM^\_PQ/)/cR>a]Q24)/b>[)C3YJKJ2S,2(^[=5EELVQ5Ed
E^;\X(OcQf93WVgTOcZ0SS6&1R5([XXZb+LSPN(Qf:DJ&D)H&_7RG()E6-]6P,A#
ML##(\],,e0+&:e6+ETbR/-be^AB>()d\gGA3[Hc:Ba4g7W&_=>D7&gF9=DZCFA8
0/\^JCN0/_K9AJPCD0gLa658g8WDCO.?fI>[XX=e^d&MZ&Y[\QHT^^D84KP=?5H=
D&8Z,<U0II=@+=&CQ[N&T;_BeAKI3WD52[4^#S^SgdECOE,YT6JWNg1Z6???aEF+
<gb?AATAa[;F<XSVQ9U:)dY_c^Wa654>f2Ga6.T,3GVJHTV?:29J#2Y,f7KC2S9M
LP1E]94E(e6L^3NTB,^GCL@\_WP?FNL.CgA[a#R@[9U8Q3MY/?]=/F#:ZMD>3)=P
R>6YK/NPBIRP8)T=0OT.MV)V8eV.,78e;N-9J5G3_e/6[;HJOHC5+GKE]?,.5E78
T-Y-(?40E=1?Z5<<&NMSB>@CBHAS()QKf4f/LCA>N2(L99PAAO<=^S5H;.QR9V_M
T[d8c1#Mc-FaG9<#S;FA9,0.\IM1Y=<Me=-D5;BSW[=N+0D3A-e+9JVg5ITT^/c+
?;;VSc#5b+8618,]^K\CCPc(-;VcOE0d>:#A5]gYKN&[=FB4PO?;9M1eAN6>NU74
PW\OACeAE6/Bf>^2a_Z<J^GOEJX&H(]+aLD)A>-5B_.#VcM7-=,\]-Fb-<(O3ZO#
L@DIW6L.g;Ba&,bVHD-MT&]<5eER]+eCQV:.\?Y^UYa])D5,:b5U7E63QSPE:P_b
0MgBVdZfM@.&/\\\cO62]HV4IR\16Z<E;CCMf\)W<-2N_#P]6^W0#/.e<OTZ(+:^
)/g5^.&C-[<Z/Wd&86&<3WR8eE.Cg:(3RA-=BRV),7)@4_G81U)&(OO-?[+0d^b)
CgUgNdIIBa/0=81>S)VcceB+a0DJgCC#[-.-&3fAFU)JCD4WJ,[[:3gW&PO)#HT[
#Zb9<QPPgR.:,^5,c=92NdPBU<,\M:;(OWKb3;58F20Z:C>LA.K?SD4N2Q(MCSX=
X-/3E;J]MLECVVfXH7e(5=^+a]&:]aJ=45cXHc&[&cW,[2;DeUg<8b7bLODYC.H,
S\07^ZZ[<+S+S]];JW;2EB]T[MYB<2g[f\;RadEQ<A,-M,4fa;bL+.>^S/O..P5P
M5d4<6@?aXXg9FCGagc1T7-6J(#K8O90\I47_4YF=5#U8QV+.c?C5UI?[MUc9ADd
BOaLKaWCO.VIID,O0B6?N5AS.[VRGF.><FE1D;IfD@?+D5@?^\M(^O8F@QMO7d]:
ae##M)9d-G8(A+Y9#B]\=Lb_bJGIb)#Bd=c/g-[-ccC<8@<VEW&:A<:M2EcK/T4c
1)JP6gA;]\gJ\5aJW4(6^NEWf5?B@611,?W\T:(TY/#>TOgg0/\DE)0>8d.fF_FR
Xg]F72\;([A>DZAQf81.4,/[6DPZ,\4Q+?=A1TaKAX4@)Z]e-Gb&X3X0WP?D:E(a
#a+V;aB#KHD:CJUJ:4W=H#8_DS9/cKJc-0+^+5[\aT;[LD8J:aJ6J,5YGLfHMS-K
+G@KG]4Z1\D3TU(:WEHUTY0?2MXT).O(C#Q[(W/,=;8Jb9O&LZ/(CMR0DQMFOLbQ
Bd.fYQ;cJJ<[@LVe(<6+BC-GQfc#R?H-[AH;4g=P4QVN_CIC(G&bX;VG=S&DL.R<
9\I<,UfEHN)4]\T?aW78.4;V?U5f_;7BJ-aKe7U6#S@CSGGfPQJdae?Z+,Ke_+[(
[A0@\e]V+TO4U#3VE,WY8QgAS\3cK+12ae>:I@O2]BDQ31](7@_8a/>T13,VF7Wa
GVS0UL\PDJQ:@QW(R7J\G(C80IIOY:VDg)8]#?7;H_(Q[7gY:11]0R_6g1CE;IKJ
;d5&@5&:\+P&Q&PHI0C.g@QCLE31g5&:K6YGY\g)YB;OHVagJ#/R2dI&a/ZA#<R.
e[]BH<\V&C\JCPF,FJ\?C1WW5]DGceL,+CHYDDF8F>R;3D^9/BgBUO7>(4NdFV2K
?_1;7-+f5F>B6&A5@D>AF72GFIgK6W^EOQfSaBW;O>9MU1I>0aZUd]C.DYRA1B;,
b<g>b;Mba\c@a_VA[O-S;4g@VLS[Z9H#\1DV;.CM#a(TW#CHI_S)EP?3Tb\+0&&>
S?W(Eb^CT)N(/BNUXD0BE^a:9C,GQ2CSf#M4H.8f<W5aDOY:LWgV.&Z^UXW7dRP\
;)^[fEM20eDWDB8??=-1AZOI1Id,+?T(b-<-]MeVL,)b6aeX-MU#8LgB&]S8MK4C
5KB6PI3-LS),/VGV@H[U,C4H-(TML<N#M1P)PTa=];]+bSXHFUd0H29=WaTPg:7G
QbUY2I40=T_U[E5B81__P1Nf9bJFB8/I#Yf^4@+K]ZJDR&5K;Dc7QQ.C7aF)D)]6
NR;:8DfF#X^S#7W6.BeV+8=agA5EE>^GYQG:VcKR[W18KH@?R1geDQ2RN:M>@S=B
BT8P(MM5g[GJ[E.)]e&8(#\BAZe:C5YC:G?(PcNP]^M=&.Re5.fACbNe9(P0JcY?
NBO4Q+/T=X=UcID=KM==KOaPUH@MV06;)=SHQZUgeL)BW8B)1ce>\)I84AKWKI?\
L-HAe[13XM4c4,W=,^aED<3+R>aO+0AU([N4WBFbbe54VPRYC?W02P(C/1J-b<?C
?JH<@2&ORR=3)+9aB]HbKf]K&\b&a+=;/;]G+Hg@EWMV^972A_(8;b<(E9U6CbE)
49]:U3:>6SPK[4gW4NET\Qc(>H?[RS2?I:.&YJbeYY/([->DFeg:?>5B4,?0Z8G2
[Y+aJ;Y1^XG]HR:ZD<?-:-U^W?#I7[NUC>Y&Xe<-Ma2fCIA2U@#Bg6Y&.9-2TDP6
+)4fC7^T_Hb6_dL98\@8N:JN&W<BTH6V>a][RN7N[P_8RU;RM6f-#2G_[ZXdcQ:P
:SB#O1IF+CI&\&K[=)4>/LHY5T.ffJNREfXO)CJ2&KHGDU.E@gaG6?4dIQZLL\b7
ff1GZIZ;&NWTGES5_3+@(3X3X_7<TY7QOLMCB<9KOVXXd<RTFX\=Qg@Ye(\Z.T^4
Vf-\0eU1)]b4NUcIU_<V9M6BUAGK0\GW>@5B;PS)U:WN6S>B8HSIJ=C/fMJ6JA:B
cAfWH&LJc:=9^X\CaY)\Y(#&(=LQ6_SJR=gEJJQ1;YWfLFcW66;eNWH#)[44DC9[
@9H+==;cf-Z>F1CP2-)dOJC.R@\M8YP4_dd6MWcVc-c.YRU3\F0W?^W4<b>R3#E)
:E&+M+=D[Q</,Lb/caGP[7bID24E;&LF#9SV1I;,W_B]W[fBg-+L8R_M,X>&U(aA
WRJaAKA0[_e?b2-=+\\,.L#<IQ8RVA60#&g^CLV@e6bg5K#9<[_J.A\Y/);23\U_
9,?A5,a)c&BJ@W?UIdH].9_3#-_R)g_dJH?\0^eSS7ddV9@52Y[;dP3:1J/[-Y,T
KT(T_-I70EOQ>DH7;X)=YDV_>R&?Y:84<TQVWG1P8<b445ZBG:2DOD5f5PI4Zd>P
=DBYEZ>F):]MLAXF;DMSO3YN6/aS-d?I(a.gDNC2SSQ:WaU&@C2.,2^9VA[G433H
fMFLQ\5NS(fI3XB+K0L\?FT:>]0CW9@K[<g]15;(33g.T3c\7XQP(5X3/d&Q#7+D
7\5U5f8+:08CCIRc:WWO/6d7)OeL#>7Q?aJ:MD&4?51_6d/O)>8Nd:Y)HIJEdf<Q
U>U2M56M<&Y3#Q<X&89I8<-U.::A/NU:O,e<eU?M0ELYQLCI,U<4:]U<:H:W(I>d
LN_&I.B=A:c4+.6RG\4Ge(Aee;R;^T/K#FeUa#FgK+bA7?S5f&I1?50MW<daN?=:
GZ+5OG01)A+36e(W)+#4+DZOY_F;YcB74Ff-XbL:8cVd#DLZ&LFF/EWTG=.5e\LN
EV:,?X28[+:OE<0X3fI_\[;Q#S+A&U_TQg<ZbXFWW;1<KD(KDI-CHIXKEYRM+T^X
F:AT3QTTM\G/-4VdSA][-KZTW/AMW?XA25JA<KB4P^W&&?#cGdOW3T1C:3TJL^,Q
[+[5C\JY/.6QMC)I26^1c]9W6\/0DCU3S#^JW#I(GWE=g0.Z-O>]Y8=Aa)UJ/_45
&V9NaB@-B5KLF?Z4ZT[=8f-DMJ-I6@VY7?WAI:>FQb_Oaf&@T:J&3a5#c.-M.2.M
>^N,&MJ0ed:6AM?9:C7TS(dGDR&,-6;J7FX60RX?65K[e,SY+RZ^@6-d@NV;N[N_
T(WJ<&T0d1bS8QV6N.V71Z@)AD5]UZ_S6@MgB-Cdef\FH[U-(9EKF1T6AX>[5K>+
?6WJT>(a,BEX,3g6&;,R]>XJL[N1g=8=&Ug&D@cR?(8YR-\+Ze4VUUGVESb/7\6X
)W8KQ@aK>6M6>>BD]D\)&IXBa]14SC_]FK7G[\)2Pg)]E]+)AR8A>B=^W7^&E4#S
O0;-S[f=2=(51:5><HM;R2W0TZCV^e<<F-#3E4]MUJFf>&/R@7,B(Mb.=[_6+g,Y
=BbdU-FWc9JDLBVD)O+bW,_#ed\#c@S[/ODbcAb;=EZHS0OX()1ce1N<6eFY,ECM
HW_U2EEWSM@OS<cGJa2FD3M_[gBT[0bEa885-Cec1MeHC$
`endprotected


`endif //GUARD_SVT_AXI_TLM_GP_SEQUENCE_COLLECTION_SV
