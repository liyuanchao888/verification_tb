


// =============================================================================
`ifndef GUARD_SVT_CHI_SCENARIO_PATTERN_SEQUENCE_COLLECTION_SV
`define GUARD_SVT_CHI_SCENARIO_PATTERN_SEQUENCE_COLLECTION_SV

// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Request Order Write followed by Request Order Read
 */

class svt_chi_req_ordered_wr_followed_by_req_ordered_rd_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
a+jSpZRYkKI2y5VbTFY7VbtTAaZds2w333/zThpF1IEESiyFMIifwv6m61CBx2DD
tTkcdhF1/EhWyMlzE71IOYMkhhVDeGZw/We4n0maEeVwOMRH/qnC6cDXMzksBFLP
KB9q/nzBDYPWHL7x5j5VosbhaqevRnWBdIGkZnN+mqM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 657       )
cbv3taC5C1/IYrrAdHwPA6bbwEC64YpwnH3BqzYWQP9N6kuwAMqfLYxVz13xJRr6
+vlaEd9PwmIxe7BFnGjNnSBR4/inLHHdpd+rP9Ut/6q57GGGH9c7E0/z7gJQXB2v
8jBdOzltKwUMxvhoJhuN+JjGXXZ86z/heXAfhRheSblfHwf/jf7z7JtCCAxqHB9S
16cNB9mpbHs+bbMJzYK971TBNgvbhnmhdT+OrMYKTisHG8VK4IW/v7hmu8DYmawt
vRQE33aM1i3yuR/d8lcDSTBaqM6TCQg9kpMoJWVbd0b9U/UrSlHvhKZx0SQ9ArnR
qrDU4JCDwGVga2zMBwgvsg1Wp+fE2kSb+UtPS1zCCeECmosDC4p/rmyr+FAfdNs0
k30CRvvyZlR7hjY/cAJzcSipWXz54N3r49YhDoxCPNsImi/ch0/8kimUa2OaqAiI
FhK4AQFC+mx8/cieEZ6kgi7QTp5OZHftt+tYKgOVoNPlRnaNBG8j+EKc1AfnwTXq
R+DfSP4WnygI0zUdnHlDKhx67UFiaj2KhFoQMqO4TIVbl2zm8dH6eDBmmqpxSG2g
YrjoRIZXTPCFI+w5l1IkPtG6aLO0O3+InNHtVQiDGO6GONj/OS0vZZMqzv9jX/6R
bujlA2xX51GOPVBLd2xzsp2inc8+TDA8JvdxKO2E5oEqFYCsWbSsB/AKX7aX2U5D
IVLsToZAtrgxnKqPMJvvWiymxx2YtrPUjDu2ksMxFg9MYfP0UOS7O8Dsi3M2zW5q
+lxCElfC9HICqb+Y2vDCVSil5qPZc1+r0qllUYxfs215QHT7Fr1HnEUwAD0TjbZz
zQGs9KmtcEKc19PTHU2XsKRsaeeyPOnth+qgJUeFbNuGZICTYTNrH/jiVTiP5uXx
`pragma protect end_protected


// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Write followed by Read
 */

class svt_chi_write_followed_by_read_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
f0oLyp3QvZi38bgfYNGcPtDAUj+zGNCnYFl0x+qYCjtXMnzRtgSmM9hICdg/fIOo
gTzyibZWlbwZf/tDgUnaJ+NR7FNmzJ9pLhN7XAfPMusMWK2fd7UuOBj8a+EDYJF/
9T0RK4btggbvIDV9pIf3W0/RIWKYEKT3vYd71XX2hT0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 1101      )
YQTwbBd3DnhalxMDaLKspLJZrSM+RWAgTcJmgk0gXzCOD+Fx1SfcsAPcEIKNE/7d
/Gi/hRTOQpLkY+l1sHr90KzDCOY8D0Pu0KbexaNWptk6XWoXSRiD41EzSCSgzEWI
Txq95ioS5+b/qoQBaHBNxGVkWx3PVYmwIejwrndsK/dRmcXmbYZgDivY4SGROdwK
yh18EYRr+yPP5YrtLXFPl6j6aAj/vyRSz3pfN2Ck/A9wlK8r02pkOBXc706j2cv2
Geu2vNOloI15XyfKdS4cCxo0pP0jumeMwF6zg5uVy4mXdvighfgwcAGxAB6aedn7
ew2nj6d+IT9YU8FUzAT43eqhSJbHX3hUaoYdUobV2lbiGfkLbvtwBniYBhxlw1x6
STNFEaS9jzK3K0R8izpw18Y0aDFmWRMkbVqUHabY/odKWj8WgWuQF0+02K75u2gJ
eAcP45kBex+fNKM+8gPieoKOLAkZ6OX+LFU+25GIQMDvvshQQ71yhBKFqaeQ3vTA
bHgIcy6d5Wz+vn+TfuACtdqxqGNKMrgYi84dKsDFpA5lnqObHEGgBoxLVSxsa9Rx
UPv2gQRV3xMkxTiI+/EBFQ==
`pragma protect end_protected


// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Write followed by Write
 */

class svt_chi_write_followed_by_write_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
FR9mDtDG5YCcAH6UP8D2B//xdFOxus8X/eFfVSD6yi9Xl2yKqy3mUR6a0Hqq/4TG
jr7wbTY3CtmDmJER603pi6JtdCIkSTTijk2jR+4fQIBE5jVazNNUUnTOMXtsusMg
zpHU2p70jJlpGrHM8XIJdgq7cFa5IOj8pnU3Pl9QoZI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 1549      )
V3Mudq7EOnQodhT+oX27llOL/TGvAZQLGAWPY+uTne+tQHCq8u00hOfg18chWs0c
G52bfPYXH/GvhzKMZixwa1dC8+MxkiWmUQH/D9WveCsoW2NseNPrCwKQWSpTv68J
vq2RD51o4X6a3rehbyDza6w2gQsthEJ4MuW+G7rUc2Cqtb+KVvRvwf7hiSBNTARZ
zwW+/phIID1lCOvtEL63jEdOZLwxr59BiQTHCeOaSni1/nxTyzH90l5V73foQRRx
IH4jFLOvihlATJwukmYQyYG8ryakcBPnYLmdfFgI8Qh8moRBxuw8KVu9TTg+vaOQ
eKtxBPsHDrB3n1DbH8qCmihqcXIccW1Se9EONNbDdXg2r9vpM2zjAbA0id028phi
u7lFxNXzC6Na1D+6GrQ+Jeum9E+LopTLnnvaVh7C7fMCD+GyP+yf0XTy4S+RXksg
n5XVW1GmAqpegzi5OwLCKA7Omxn3NT0coRsdn8NPZBpBNio+3+yKac2+6Pzh9KTp
LkPrP+9SQyS9+9I3HTupdtIbboplaexMEHs1Zo9nE9fVGz5PFXOroB6yaC2WWtGN
go2NQkDTsNt1Bywbu2DhlVvwY7VEKoClLkQw0zH96Z8=
`pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Read followed by Read
 */

class svt_chi_read_followed_by_read_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
nq1PFUaXafv0KJ1s9JFFY8TBm5Oliwxiu2gpoHfbLlK2yrNyW+eOvupzo89OZ6Q3
VTLemUqJZY2xM4s81F0ZOZUsIoViGjbK5uhQDkAuPXg1/Wsnp68YuDZ1HrpX/Daj
MNFzfbwSWYODKEXKTP4KWZ/6JplPkF86LEVOhaw5Gek=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 1989      )
eCdQtLBvECcLmOnP43CDXPQ+nq0vv5bD8qN4ddQZMgJ1oa0TU0VrTf0XF+i0goec
a+LizmnSAhgIJ3m5XR50EcGqBz1Z6EWUsN+ewfLMq+5RbvcVRuZQkIrMmQwvgevG
pdJxDfANMU03uJ5Z0G89yhf5nScSlq2Xxi/woMXQ2bl2YmuPw0pLpjPcckunTzyO
Uix8VwP1vpD6Vu6S7H4kC6a8m4Ti3xzN6kZdZAm81cI89jHdGdtFRX6lLncw7kbR
XN2W0IY8uXgfpT+Wvhn0a6kWHLX8XtGtQW5YelQwhlcWf8heN/DKpAXSTDqUgCTp
IOGgUQt8Lid6QOqsry+JoxiUIk6J72DSuAY1p3QPNrxREYe/Ha5s6LSzjOAPJo7x
1tNfRAB/oUco1Rdx/W4rGbvLeL2qYwSa+Ycy3KSzBfw1F1bNUpDRW+MQT8N5eAHS
TLoUQUIPA2iGqWuiwNXetGNR3lRVAYfj7AvmYpl3V7Ji9vh4Ki+b4ld0v9pmg2bt
ShQQrJmXn6WLT3Y6IBWDE7QjmMzmu9F9j6CmB06vGmauwAq+JAm2z66lo7RoxIPn
LM+gHBMeichd4r25X5agHA==
`pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Read followed by Write
 */

class svt_chi_read_followed_by_write_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
fEgLXKOY4nkmBpqvyiRlKEThqu3xL177cyo2dnzCc4ab9sFbjm5nwi3+jchbECoa
XApSMAd9mGICtqYqwq1cSRnlNFlYWcoQhFaRuq3zPIw0FqQHiBZNCA8x+aSTfuec
8c/qcTbe6CRAtsYMtvlTk08UYicSmmp31JAOjxdVAKo=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 2433      )
QRn0Z2cEzDj+vHwSGUBG3q8NkRt+wV1xtxBYad6Fwnwzy+75MencpJdz2uGazOG7
u1XgxqEncg2pF9XrbLFWxB8q+iVt//bp4TcTkowLnb83ddKERHmRExiVokCFIBWY
bhSO1muyIfpf3eXtqoXai5nrPUTpqLUsh/ov061DGLG9rKl0WwtwROLo8p847Orh
yx9FScGawD/YeYR5vuDQ9NimCjN60ArchTZDjWrdSrTYMYMtCoVEhILd0Zm/EuGF
3zalucoCeH+OaAvTOLqH8LsOv81PNehNL6guM4XfZgYnmTlVHjaEcPvg9Vp6GCw4
+FfdMJLV/9UrH/ldcBkOwn608vC3Ej0ZGccPiFHoMLGAHDs7CDa6h3HFXvMgZZxd
gw5mtd2+qyIVLE1lOH+8x+EWSJr8Hp+a3v79B+SDpZRDM4xOsk+P16llRzVDCJzw
/pMyyUXPjEFyX4EL3QRDOwqErgSerAA3ivX1BA6/tzRbiIyI3e+pBcqBLwjMdsbg
GgkQHbsftpxxOGeUVy1EERd17+BNSY6/GLQlsHqmVLPvUbChIptS8g0RO9iM7WyD
Z01/oZwJUUypelOzLBo1Zw==
`pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * 'N' times Back2Back Order Type Transaction
 */

class svt_chi_back2back_order_type_pattern_sequence extends svt_pattern_sequence;
  extern function new(int  pttrn_seq_id = -1, int unsigned  n_times, svt_chi_transaction::order_type_enum  order_type, bit  match=1'b1);
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
m4YVt0WrPDY4D5Eq7v38CCEaW8svBFFTNXMvpZCHtjf1WnyVkL6E9XO/HDWNCJi6
+2FFfNBPbtenXThuT24PlM4gsu+sw6PVUC9a8fZ69Iheh9hyRKsyLpTqP0hEsVzD
Nyhe6P6HDVqeYlh4/TG8bVPDcEe9bAqwJASdDlpun78=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 3207      )
jnG9jrte1Ht2O3FmtlxnZVvWX4m2Oj5Ti2zX9B0FHTN8XOLpULnWuZ8bFhj40LnJ
onx7VTC7jtkWvWK05I8tYgjKdZnhyBrmhThT6gp2seVHzOxqK9GiWu+FwhApcgk1
W4faRNdnG67Ldgtlxz+2ERndad2cUB7CtUchqG/29VuIeZRIs1eP3BgBNNXBHMJh
MJR2uWxIM+dBTCAKM0Dic/g9WZ/lLnj/dcGSK+RyVQliKDOj+jJ2ThbreRmTYNu5
JaXo3C9LeRJqkPELvurTCqCgNQgOSTrMnVT4pd1/2/jNcCP4xyFusauNVDxPzPFc
h9kjTXo3mSAW2eInX/G5Lv7D3PKSSnh4O6uffj+PeObNo7MFSA6uAbn0poIuYl04
WwG/XlOkvfXxPLaZC6IGt7X45QyW6urFimY4c8GqeJNmShybNsuE+wmtq1CP0+dq
yPA689/sldmbocFY73iH3fAxAgV7CNwkwAwHsPjxp2EUlCWCwUeB8ERbuZbnSOaq
JeTQa+WN+by3VG9Gc094FB82x9RksqL6Av1d2dL3Q4gfT79f2iQbMxGajBQSjOYx
X0LJCD2OPYZhKMFYpJ7wN94GGzo6B1HEyHPs1WXWWT2BsGypdKUROfx58YJKlEhL
EsFzvi6tvenem8h3Uq1nY98xgn+RgC8VqwO9g47DanqksYYHxy0EAM41MYjCtE0N
+NgoAek1Ete/NM5ZjVywsAabOXsopZGr0uHhtq5FYDqKLQ9nO6F7SOi91Hh8FF4+
M0WheOIDSWP6WwuKZaKA5eD3sQRtHH71BefF/WCZRdVtD0s0EIpvMTqZQu8zEYfm
QeJ+VYqrWuSUDz0yyiYMbKUFJBSGbwxkHM3BcNG24h3NAzq24l7deBR7VWCBtGNm
ANdbQlu/qs4zq5e8vcxh3N6aqdGUSqH5/Ya5HdCJ41h0770VfwK3IMsKtynMA4me
n/qQNfl98c4W9XAY/KVS/5KTLnfHefHYsjCFRmlxZlsTI7YaMIadtRFrqmgmDrq5
jdC2XGhJttXzZqy53/9OIQ==
`pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Non No-Ordering Order Write/Read followed by Non No-Ordering Order Write/Read followed by No-Ordering Read
 * with Same Address/Different-Different Address.
 *
 * i.e. '1. Request/Endpoint Order WR/RD[Same Addr]  ------->  2. Request/Endpoint Order WR/RD[Same Addr]  ------->  3. No Ordering RD[Same Addr]'
 * i.e. '1. Request/Endpoint Order WR/RD[Diff Addr]  ------->  2. Request/Endpoint Order WR/RD[Diff Addr]  ------->  3. No Ordering RD[Diff Addr]'
 */

class svt_chi_no_ordering_rd_after_two_non_no_ordering_transaction_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
jXs8aRGjjWFYeSPd/4o2w7LyV1NG7IJGRX8QoTdh7mdITc6x+NDNIDbEyQ8W68GT
4c09DweBwsMQRyHh1tT+CCE6XEVMRZ1vLeR7l0XiAZf0eEKdv8Xuvsslxpk767P9
bvl1IRZjV0raEGCE/RhgDC33J9me7ZHIeUnYWx5SMFU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 3984      )
rnietU+1tMHBxXUq62As5NyBYJMnNhahX7B5q9D1uRBwK+xcNKR+dW4jDKEPCB4M
aGBJOL97vU7rs6JeyWttmMXiAaX8yvs/9Hd/eYifiJ5FkYK/26bkuMo8PPy0lI+5
+OfII0BLAf5f5z4Bdsf1IXVQdUAA4wzS4FCmF2PAb7lwgmGAwHHKnaGIOcK/+n5E
s31QwIyV3wJQJkBA523puPU/P1WhGfMV5o38a03u2GCCO2uCqnLJcDnsEsBdrUeU
9tz61SmKe6XE1UHwSbrfRYOznIU60sSnTi48aeeVHrWnOrLpwu3kKp2ZTf0XdCSj
Cp/VqE6Sw5l18zm3tvG0lztLL2qrHh7mO03aJyUv9edUjKyPgtjXrL2CFq2PkOiA
1FTD4lL/hh3sYrNtHOwEzY5sDfOJ0oOERJkqykKfv3go02BbBWZ3YaMLwlZJtR/y
XZft6ohBt9Pu2wDKxTObokFzcPU/eQ7qCIP/p0WU2qsT+pQtH3NvHgoieFViRVxs
2xRrXM7mPzQYjJTSXBR9HVbZMT+rOAr9JecbDLomqkvUwT8HFwgDpNHP2lHjmHde
NGZre+QHVr/jXampCen13xbdn3ig5ixom0GXtUll744kjBj344pfu9FN1i9H7+PZ
Rk+l6GODqC/3bS3fJv+KeOkFGqte3flS0at5z3nmMLShb0R5agykE3RBhAm/Yvme
ei2+YWSWwQx8QKEk2GH1/GbLCSD8qHrECAFTKVJRnZdCBeCIKUedZzwhvPRD3c0v
63V5QDYSty1yE6UR+pMfd+ZIFGjbDDCVlvkkbgUjaeii8rkD8a6UV410PBQtr81k
bGjr0REMC3A8iiDiZsQ+sFWgxGs7TK5C2UC4WRMKciyNRQN13fKn5acomUkziPDd
XnCf3sYF+wPzM3EzHxy3NvwPTB1Qp245Nm0n1I5oNCKetkaC6TeeK4pcx/IWGD3f
LTSABBwgpJSvql4eQO8VgLiDwZZoy+VYktgh69u2fdQ3eqIfqcRsQzajLdkJqmyY
19do/hWcBJuR+Pjy+9/OZg==
`pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * 'N' times Back2Back CHI Transactions of Same Source-ID
 */

class svt_chi_back2back_transaction_same_src_id_pattern_sequence extends svt_pattern_sequence;
  extern function new(svt_chi_node_configuration  cfg, int  pttrn_seq_id = -1, int unsigned  n_times);
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
i+GqNumAQfxA5ZSKbAYZWvBzLLSEoAgqUDRV+WD3TM+A6Hc6xVaHkLfSbm4V+yxX
HvvZ0YF33P1YVd2HxFfu6gxogK2ltriHLNPc2lY1nAszAB+fDUwmlEDBQPHdU1dS
kqVL/mhWaEE7MHy0YUc29VOG5cJZzQosK5+jxEr2L0Q=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 4940      )
YoL6efhMQAx1iYNa/84Q86ZyvFyZLgtLXZj9MwFdwo1600leikgo5nubYVkMkdao
+jiAeCEPKVdfEVqXODamjfVtUoEI/VOIiSNM56R4sVRxFYGF//qt4EXqVyiHwno3
YMtw5pQM5wVnq/HeOtfRe8o3knmJsLGTERMgNwUhyf2QBBj89VgTQyAgS3lLoUXc
mug28vDCVLXGNoNmEYdiO0aWTN7xVOGZ+dOftdB8CUg2FX6ns6nKSlE5LqwUGMu6
eblHUmwg5/mhUOBmfW7z8eXDjGF/hSuVzWMN/V8PS1tBPxcPFxEEhCLinIK7/deR
NlSX9rfzbulVDMwvyY0atzWi9CBQONA56FuTNxPaCap/ldcKdGtTB7ot09Ppy3sE
hKstpxVqNIgswR5Md1vyDEK0sjeEA/qVLz8+TUyXBg7LwdE0UWQ9ZMEpIPV8ym9j
G2hxf7xL7mLtgo2J+KgwIIzNEHVPIdSdI8XjYz5VP39l8BhzO+PLc+Cy4yiM7pAz
pj9IXYKPSE2cgtifx9nO/a+riMCOWv4ENSK1B2aPSvtCKNTXR5x6mBYs5izYK0WU
Cem5PLmQQM+T5vJPEP1tCqHip2rSrFS/fWE0dZjtvYJS7a/RxTGr5PwMH3X+euvb
2g9yPNvB0VAFIXkHsi+d4omftmG8UlWclRZl5Y4veyKfVZ/WWKtRwAqN1Oekr9Ug
s8+3N0jAkZXQ6KuQ9ur9yGEaiulkIEV7BCykOsvny9IMax9Wy5Sg9DiE3zN3wFWC
5rbCYgOGWWc5nG5SRHnpdxNCWDbVujkQsRa6neLgVyt8oAK0tTfNlerDHtaD+A4Z
nwcieOG/YDT9gFYD04K9XaoTpyHYUGUo2cfM1o3F7ML5t2zMGSqS9kzUsvfbA74D
CS/5XmfM8UFi0e3hWnjNA77h5BHDb5kPpCL8qf1oLza8fCdfLz1BpvhJbuouVdZU
5CSzM12MC/ItGJsryUnC2+oqoTD/EYn3lizJHrOyIlYCVUYwdF5u9GFtrnfRv6YI
i2G0GDCvlqx2OdNlrYnzVgGl8Cox/avLKSiLCHd9IXA5UnJsCDtqg6rFA/1kU+60
drwxTrKeEM/YTiT1T57z7pyAmTgvPT7p8/YvAuNJxCVRqWEQuEAbxC9ChGx/2Hbf
M3OXRGlxFUIxdz61ybn8tOVqTQ6AEGP7RP0sP1wzKa//Uhc7q8rmQ6+o3PVVqiY+
lVmyq40ne3PaCP7Ahmx+I7CKmrpv1mfSQFPqn1OR0yLxdUbzUiX7dSvNNyW5J6yV
`pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * CHI-B Spec Figure 2-23::Three Read Request Order Example
 * Ordered READ#1 ---> Ordered READ#2 ---> Retry Ordered READ#2 ---> Ordered READ#3
 */

class svt_chi_three_read_request_ordering_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
J4R3NA4hi7Y2EvvyuhqkC7KZoC6ePMamw6rkjgCJaw/P7yh5a/7zYZg8eak8OuDQ
QYaeUNbnifqMJArqUtte68T8CokjH7eR0IoBGifZbb9Icsy4vrC3FbUsDjMYXtbu
FVmeKLtUDLu7B8nu7tnibEn1UqEq7w0s2eIOQWUQv0E=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 6112      )
Crv6B6NwAhTVTIEGp25F9a5ixUwON64BsrLUMldBBrS4mn/Udlo7f0Rs6F3Oa6Ws
oWXVTJ4RY4DBhS7UkCWEc3T1oMtNChMdhbZLsBfhjIhg7BJHX4hKYwt25dUo5I0N
RvTk7ZUm1GKq/a5t+TcV0nAqbYDvkmhoJ1QKRpnua2cvmyW2Lz9msy5D3Yn4oNOG
fabrmyhA0Stz8gsOHM0F3F6vKCi4QZV2KhgnGurXQ/rWlX3UxxVrdWQ4Jpc/nwBT
lE/bcd3O+OBqT7BI63U5WVzLL7O4vZruUryQMNbU8CLjCvbzGWHNzjy7viqjStK6
7XhaWgIndwW60ucERMfGSze8DYtUOE0InJju7ZSvyTZmUrJ8yeUqqrJyNYKXD0la
AcCE078K5AOCpsNwnucL64mAItt6YuMATNeIBLPiRgnRfIDzLUkTC5v10+WjDqRQ
xTs6T3vLY/uSzhHr9mtQ4Gq5Oa5u70dUgKQmSUBoPXU6POIJBpJdy4BNb7hJ3yOd
TT00vTNP/wlBsPsQyTK+MPaaGZr624476qEbRvYdeKcCYIms1/kFdDgRXIL5hJX6
RHgTAcJoLmBx166dVGOSALxpEITWPSZl0osIjgjYh8Yg2CCX6uVt0gP43cR5F+KC
h1o8kowCoYUl8joQBSF2iBxmkXQAnA1VpMkY5ViKbNPVHOp7vEEamGWojW9gkIdp
OWJiAGkVssy5ITCFELp0zmBPNcHTKVJSsfRirpGI0ukyYJbZFD+oQs8LOJkq4qQ9
+jqOOFSA9nzQUyC3FjZQIXUlKn74Z2JRi8rFsPbSdMxhjHTQ8bYWkSMXe/BBrQKW
MWEoNJnXkwbCraRCGuOK186RJNOUHIGt9UHJ6nCqK8PwNo7TIIpOiOhTYJupHbDS
8PhgCdUjL2AumBGxlUM0+SdAov1edrXzBxdtg+PY5Q9OsZ9aCjW1bJVdCn243nJ6
vIZ5uVhZXDoLAHdQ7a9aniCxDyokQKW9XZXwStgLlyewhFDoEuYN81eTm2asrmUv
K8aTrhsIpNLOj6oTTEqGLhi9j7i0MNfk50ncpNpvCXtqFSgJw69LdwrCOCeoAoLQ
nYXjc07bhSEZYw4xhnZKXD0MwKjGo0lZfBGquUZ2OevAcCRDj0wPRC2i1TezDLV9
8urzL+u8QzoJefVEoMXMq6Su5k9ZLLa3dJ9EFVKRNN1UZa9lYlSVyqzVH7xYB5nP
xhFpX4clObd0RMh1hdEdnusbNG3vj4kgYu/zD/oGwaVZnvu2vK/Lipyg70yHQuCD
Pi4e6eNanUDmQh+ky5i30g9EboaCPYgPPXXla2gAkediW3bLjgOZNFLX/P3i9YVd
nWNz28o4y1lFiqnuB9bfCWzulAENGQLn/gXcFoNqNS1pzN07+K8vwh492LKsavem
mH7aUo4wDC3K64PyANDR+pUqFOo12fQKuI1rKTO5TN/h7zm/dyJQ1SwSTRBec13/
wowf63Ir5to9yjW+mN/kmZertUTGou5gi2zcCPAZ6VVGB9MlVbEVtJqykOdePykC
11JDWapP0kunfuT9cHhT+WMYmm+tkz9aZVBbLX0uvgc=
`pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     Any Normal CHI Transaction#1 ---> Retried Transaction of #1 with same/different TxnID of #1 ---> Any Normal CHI Transaction#2 with same TxnID of #1
 */

class svt_chi_retry_transaction_between_two_normal_transaction_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
OQ274kfWYVDwFhzPNViOvgBLqeXlSBYSLF7yjVR1Kyn8Cg8L6ktZMMCbCVlx4xfE
z9fo/xds1azSlPha+Z4cqa1XsB5GLUmE2bvnQ/v1M48SO5c9gaHxD1ycNOTtS5p1
hllKuuInqg1RxVFQS3BA4ilec006OpF34KtvqnTEajY=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 6670      )
HuVASAYPZlM0GMUHd5gzaHRBgtbdNSm9pyt+ZOLft9SKWm8OWsrHxGPzrF6xkziW
7Ae9Xp64eE6XxFQnWZxGQvFUG92e8KawzTFRA+3fObSlDGVgttsBwn6IFiK6RdhU
Obp84bsgVrM3aHJc+ARZ6xf/gCYErqpgDT6Rq9fNmi4w4h5szFvUMOXpAnCNC9iV
kUUl/Jxl5xQ1z+ZddV+kZjPIc7os5JTzXn2/1AYlw5qoYlGXAfE7x1FA5Z4Q4HYF
HGIyvg9xkJeHPWrDeyDwn5ArSbq/Ic//sTnTUIx2fLUwP4cAUanoAg/pRoBJeVlK
ebknyLrgDwUu5ju7k/luwZxFBaYYs7g4jmKiIxhDhIDeZE0VKrVxwWT5plMLjiU3
YhjlXg+JisCPAOiSjTRxy9rfuEkRx6q8dVaMtY2exL2CM9BAHiSYiHb4E0d64RdM
jvedYFvbCd4fYAnfQ+Bl8/5GKyQkRoO+x9d7m+MVwDeGuGlxiVq8hSvkVjxvYX2y
V5CxdUwxn7v0RRW6/8QqF2L8bD5aKFSqN85qoEmxH9pZHL5ediiqy7GCOqG7RNub
w5zLuI3txtWcCV9iTBKXyIirvS2L7/0mX7RC50GpJRrbrM++HC10p9NeqpQjaqWs
kgH8wuGB3qPdAMTD4HPHp9KEr7g9meM5HvTrnP0IIi+0clz89SNPshatjJXX7vZ3
lPH3IvbYGldDORd+xuTp6HtBRpecnSjZg3tfTJ4lfCE=
`pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     Any Normal CHI Transaction#1 ---> Cancelled Transaction of #1 on Retry Request ---> Any Normal CHI Transaction#2 with same TxnID of #1
 */

class svt_chi_cancel_transaction_between_two_normal_transaction_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
RbYQzNeXuVJuv7+Yb4D5G4UcBo+jL7Ude+RMC6zg3iDVBxkLBlVhPQd5wf3kvPhr
kufBNflIRbS+Fm0yNZ7cPfz0xwgYh7ObzgnBlxuZCFNeuTUr+S6UVDr+i0ITaO/s
u4maPedDvtNU9RtWRRLm1eefdN16CadA79kKkrqGV3Q=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 7280      )
pyvFIn042enLKKrc1yi521bjikTDPcCdnZHG3ZnPijPq/YXrabFqH5F4W+W4Al8t
8WDQtjZ8EHEnjfJcTbVuKGrlX1QkLIPuhPJb+gwsqV8XiX2ipaHZVndBoanz9Ei4
n2jOy5rzY3t8BRc9mgqDxuEHcPd/svNdhQB59OeLuhKeCAl/89xpb2Gynk8Sh9zW
SjJwnVoxbj7OZVKy+isj4d7YUa7yRmBfEeEmQkMsO8HiHVGNFadGU52HTw+tQZPs
SNkoKq3oIiXlIC3JOl3WDnarluyq4QfPBhW+D9XnfxmODyW+OLtNRvAuIfDFKcTM
Ij8UYJ+5LP2x076cBaU7/borR9Cl4J2NhYtBbfVq/YY7d/K1s1pSrxcV0OjKrCuS
vMZwEeu1Semy42FnRlDOBWQFFdtH5ZnnciIsWW2tpKlujMU2XOfA2YH7z9gGVNvO
qkf9G+HiYG9gW449ZE45gPH91pNfsoZqrhmDYtGZ2gepds0z9p9Oa/2ris6pTDFX
/95uRSHdZ4U0Y3Qb57hj5P3D7+fVuifp0ycARe5mUKp6NrqMALmGJLLd8bT9PSoS
4Bc5eN29T0URYU29FyscFjs4fR3Oshj/wm9Sjbbcsq2H0PMLLPQne/l1r+aGD62n
4JpN0sdGQialORdM1VyrLAkumDYCd0oWWlHp7+7Md2ZYLAW7Ll2v/2HWca+6vkQf
LDONKQrb2y6NoBdYpSMb6a98E/U+YnB9kWABn7Fidin8xrtdNNAg5SaNT0IAKaj0
cu2QC1rDfORJCd5HvhTowI+bCniO+zz1nxfN6i6vgbPu97qtv9VfeOYLRLlSLlqB
`pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     Any Normal CHI Transaction#1 ---> Retried Transaction of #1 with same/different TxnID of #1 ---> Any Normal CHI Transaction#2 with same TxnID of #1
 */

class svt_chi_retry_transaction_after_two_normal_transaction_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Bd4PZetG/TvF/Hjn6zA/o64+RfONINV0yZuQHd6Z2OPwIMaYyktia05Od+B26yLi
XOPCJBFLHvG10R3ltV1V1GpMoh1tjcSNVYiabOZAdAehCr2t2aJWuqlZIw0YkqVZ
7neWHZz7Lg7e1fsQNeDaYVLjUJ0cFXPydvmRCpkIvaI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 7833      )
122ecPdgy3qW/v7kt/wWbSe5o2D6Es4YkWY7vWHVAJn7ySuMjyWfoBI5LZOKgIFW
wvlWD8iXoRkN8Kw00flWQuccCad0bNf70pr96BOTo64ub/Mh9Kvv9jbYfd3lc61d
f8oRBFnGivErDVwNufZJADoCwvtU18AaTNoIvS+0SBWMMl2ywEcIU40ggO0/l3xq
F2MBwjVZxeePdUN4hq2nWkFpNv2w5xxOSHf05TPCP+T+Q+c3ohyfMKajRbUIf/CF
1/3QZ/ITivnU3dZzcnq/3BZ/pHfs+jCNnHAbqSqW9l1bfrqg8mC6p29+J+VVRNhT
xqtv6zNDl1ZyyOH7f4we+mFvL+r/aedUdHoikehlpQ8Okkb/J7ZnLTLsb0rnnIcG
k6aRJAY2z4eLeE8JsmFGvb30QFSk+n5/w6VXck8Wwtserr83uAlK1SfJgt3ZMCZx
QzDmeivUKLY/tPerURBjh+xAfNB9hsOFEeeLIvqauoq9wa+xPg1iGVztayFF6Eky
HvgKMa4/Dqpk58nToJ/MwuIjYuiUoyUlS8t/oBZctBsHyZa1UAMuUHZQInUkwYrN
gkJqX+YXQThYv3i3VbzLbke1OJHFI3nOJ/O0D690GMmkOEwQrIsAAua+S7u0pqv4
kCTS8pK4VKqRwxEwu2N3jYFhuzR6pZ8nY0ZNQToeadTNLOjhqu/ASXf4vn0HH+a7
0CMMq9rgTgRKl8IvwIKdWLelH7R74ES4j5E+RHwcqvs=
`pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     Any Normal CHI Transaction#1 ---> Any Normal CHI Transaction#2 with same TxnID of #1 ---> Cancelled Transaction of #1 on Retry Request
 */

class svt_chi_cancel_transaction_after_two_normal_transaction_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
SxhwS4ZekwHGC0/UONgKD7oedNYMxMb60vwXI7HnmTta9ngDeG7nd9KAOdVwmE2E
qhA4V/o9oy55sHle+VuR11c7kzH4AKis0a0scba4lEQ0YjEz+njPVko4mTXpifMC
DeznvX1OW4jQb/MOdQCT+IGqktNZZ4M485rPqCpbyTo=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 8437      )
TWr06y3GoCi6MUO7QROpFd28IsKg48nyPRcWHtp0GCMV424RTbJqemkFENP6uTTX
viK0oscYUFoY4CE6JZuaXbFZkoVH3UxiTliRvQRjDqwQT4n3TBrZu32V6KrJ9kJx
TSjTY81cFovNqRXkIdISp8ks6Xg0vwfXWrFw8QosMREIYrEpFMS8ADcB0EOysB2j
eIdoeUEnvyLVXoRR8Bq6amh4Hz0hve/XzIN9vwk3b41WwA1A/Cf9bc9Vf0biyzjN
1Do+jcYkXw35VQmv++pL7uW7kzbhdP0R74RRSfcnyIrTtN1jzHFJrknjAju2WLRr
A5eN01/a+U45KePBiwX1O9wJlHs/mQRKIOy7O8OFT+oQVAXotj+sNef0KkZVLrYe
5O9LEfOfwX3gaLtxQrC7gXqCBmSdNlVBYRpokC3+CptZS5L+3Yl+rf52ML6V/gs+
j1kVjLA15cLg729qmLO3que/KKNRQ838ViZcOx5VvHgcoxRqGFCdzWrLjX9086RJ
SXWLvm2np/nYCPAuH4CnlwIoXNGX2kC3wxKfysKpYAD3y+6VZTgTPC8y81AAhtdB
w+cusS6JOMqvw0iS6PJG2AIrNgRF6QR3wm1Zi/kgN4ea1poUbcux3DJ53Q4dt1RV
Nybp77v/wvZWjw13rr2W/AqsVQ6AhmnXYblcZ5yOpqxyrXdmE+DyVmMYGUCqE4O2
ZjSODRvVBTwZ0V6biVBr30Enumjhnu0Q57oeHOR2MuBWrUPgSnTPd9BhdCVvqvdl
kRQf/MdYpW2C/IROSifW+UI6CMkz+WouMO6ts9tvDK0=
`pragma protect end_protected


/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
OPG3EiGwNm0noOshmX+rAIqTkp7rowhHKc72HUEthajThZ894kegPTX6Z9gVSeL8
hsrg6mGbbzhWrSGoeMfq2xBj38y8f+Pdm+MRChe1d5bARlLXm9sLYpiTsOsKbAm6
ygZSreek3r4bFTems0Rrz7pTYz4pwJb9jsGb6JsoQds=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 9077      )
5pXAP0+57LymS8ZntFhCRd/cB/ocykZpj+J3gXP+v76vEqudyw7dxoVBV2AdDSDT
Ok9Q68MPKCZhTzVNpgR4EK0BUKYXfhzObwyAP4JZWBbaWBmGQRn4JroGn6xrtnvp
G8lvTmipI51IlJozjKsIeFPDm5uSlJUNutupy6FeXgSvuZnVJbgWtbvA7eOXdLgo
dpB7IDVKFBdFykbEKPXz9Usr3OooiNLTG2A3VVNoKy9B8+4Y/Yb2U5rCxbCIHIp7
Zy4n3pf7qGMJ+qj3igHsFWNSClxk7+24PQ/EErccjwX7k0GnUFxg0E81TqebxYyf
l0HoaTN/SunNRIqZEyPhphvgyAwGu0pZELoNafj4hGGDiCsHauQ7FCx1WHULbHXZ
TJUNGUqSn47WZPnnj8BFahPOeEirUq/TANMUesaOI8BFciiNeoe/q5QJA6UoJ/OA
7lFf753R6WxTWfJGMxSv5Md1rJklMH746NQvh2LNNfdF0cr4sXVTG4qMTiNsbYRp
hGEdg6yZmXEgvdQU887QEsjcVOMyIwfBHSuMLZY+r2+nBrAjcdITXNjAA+J/DRrz
+y2jGEcMkgTYZaSDta8LbASkzTGQ4TDO5VugRufoiI83iSX/pB7Bs+WRU/Rx4grn
KRoR2bAkrVcOZKgI0NX2l5CvFB5m8UOyG8cqwL0DPqzSGl58IDeVKgR9efV7lWOE
NKe4+CDs5pD6iKVsJaMaQlKSwpAPrCp2Kitf8uwytSKs8mDX7vpgWRAry+QNk4fA
sPhn8SCtwcEf0Ntj1IAbWMj48w9As5xkzc3fSrec9611F3/Er1oEJHHT+k4XLQV8
JM8g8+JMuP7T33O1DED12BQhGf7+IHrqM+1IeskJD5k=
`pragma protect end_protected

/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI outstanding followed by DVMOp Sync followed by Retry DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_outstanding_followed_by_dvmop_sync_followed_by_retry_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Ob02+93uft67VVaH3bLSGXUFgJGM3JM2riv1W3G4WhX5i2+24nrgy6R19POFTtTc
ME1bLBeljot2uJZIQ6vFw9YyzsgJGyDmzkZmtQ1ehs47LVGWm53GMj3igWjJ1WvL
QdoEPiEOzGSXOXKLSFJ3zpP+Q4HvAsZoYamqVAEPhhU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 9858      )
kXi5czGPw1mfAzrMrSmIsUrGIUhQ6Nr00sr+LeE4m2/k+z5Cy8J0UJiPE9hKnk6x
/IPLTd/a0L/rk38hi3kr69llybSGujByT1+3PUtjWt3fX1Z2aFLribda7g8S1pyP
HBm5HiZ48ajuZNk/kUyXYiwdMvdNQK38MuT5FLvUeoLCuaSC9zs1A8wuKeAkJ/O1
rQXLCG3ETwyCv3WNFVVscYhAA+mSXj9A8q//rTSNIGmemUC6DyJzykr4OIHxTwET
kbVxU+RvxuhGlkvqwnyD3U2K0hzeavyXL2fWemL3DSLR3Fmb09fHF8QkhMjok65G
P9w4Zb1bKooQrxSLzGkp3uiJGB8JLOY/J+iw9Q1sfbKko8FabJ4ZaLlYjOtBvKq0
pHwP25oKEtXAEJVk1zjV1Xzw2XB3ugJipXj0qFJFcszGu9hkOMJE7PFnWJ28VgtG
zq+ek39EIL5AnI2mdpfaSPU1O+ZxSg5ABfogyNnph4AvmXWk4gAL1/lPT0u8Rra+
8p9o9mQLx+PscX6w36JdvQFrPQYhDk6Nsk8SHwbEz7WwpE2fK5lTx6nRY4QeH+0e
7mW1XK10Rn6Ct34J2EqQgCba2wuhntBGhTVZPERoTcHLbiiU3fPNHwYwMllke5XE
Y2CdInnaFsA4F2RLTLspzmU/QtRQ6X3BfeIZMuQE/1HkjntTDZiP3dJzNyEZ/6Ds
aS/PgHAiQW+zcAKFOfhJCvSyd2WU4lKPvzJIKFGZvceV+41H8cppVyTT7vbuNfRS
a/F79eEolUDv24gcSoduqDb0tc2mrBt6xj3VJGQprBU0LOe3s1D2iKTC+lTiQjwD
6lIoCdyRYPma0nta+L51Hra64P+oUQrFIPbMVWfZxbjvFME9tOTuohCEPjpv20Af
z3VidQAKKwZduz0tpSP+ppbQalEObmkBUns9+Jg1HCMnl9/vKFwK55q1BKIVzk3h
cr30Jed/fh66eK76ACp8A174OYsosHP9SBLwThq7yXy4FrKuRh0aAxr2X5a2f+ZG
e2IC98XTEVytvPc4uSwTvA==
`pragma protect end_protected

/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI outstanding followed by DVMOp TLBI followed by Retry DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_outstanding_followed_by_dvmop_tlbi_followed_by_retry_dvmop_tlbi_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
QT0VQgjSa2ZkatMaah/ZL9KDegpu2hHXRVuJQfWigVYbM5kH4H3YT4zcQRj7LH1H
kkCH/EuGk/dpTu1VQdtF9S/mx49a/j8DPoTec9laMfYRPTZNzd/Fevpft3asgFNF
ydu3mxp79boVAUja9sa8Y0drn5tcVCBMxpdLcwFD15U=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 10751     )
eHuIMw1ngwCkDEjiC9UQF9vbHAdOppt6K3Mdf5seuaaUoPwFFBiq1SwWTYFv4ctb
OfKZhX7pyffa1BviNI56Nz97Vzs4aSeeKMwSM0P/Jd0P2Lf5D7lDoc1f0yVLjxre
S/DAGAOhFHdX2/zg7Om9pW50e2X61tqGq8hTJFeYb2y90urhO1WHid/E/1EvZ6fT
ee7zp9KYykSXG3b8Oz0lsCy25Rd3Cn+7msO96FBQ0UDe0gcmz8+b+BqIRwO9LLAU
zR5POr7IaRojdkBTTiWxBIOfqhUbXXMboDU2J3gynG+rLeoeCDjYH0wO00W5rhs0
jqiwLyBvjsSuUNwLAqazrYR0aY8o9mK4poYeTteGE8XlNr+d+3a2xvrJJS8F5IWx
F8HtBl1N95exi5NPQP2ZHOCMBJYoUwB5FMKxw5swv8Xwru/uy6FAtrohhBclnMVI
ZND2zJo6C78VZJ/EQmqhiq0bHUK8F5bVeLyuEjKv0CaV6quPzaDlmAgjGIpSzVz5
dWiQQPdjSC117nTY4hXtVB/hbrmSOzxhIuPBPcN35rkPNLCah4Ya6gRJ0gF9bZz0
8KbyuWZt7VSOEanuT+aQd0eOckYtVs1Q9tlmJEMR9wpjbaeXHqnqUChG6Cijvdp6
3JLN9CxE78FgoAtOD7umbYFJKTC4d9zbe+kwnWEXBIYZyY8HFUDMv3QlhDYkJ+Yj
r1DX1gqycomjI0m3kkL2RtqTg44TsblWuzVYPrCaVYzDa+bvJs5LRP1QS0wM52xg
8H7sfoHnn+wimj+iqNgNMKYwaTFXluJYLQbKhwDEsHHTLtSIFFn3hvtXw+xpgD+X
ZrijaQoWeC83I6RPr3Yq+kU7e84quMBt6h9IUqd5E1CTifDGdWUq6fXcKG6V9OVP
W0YHtjG2xMfm4WfTGzpTnGxwipmQkEHm1+0Nj6jwpKDTbCiV4/Ud6xA2RSPJMHFV
MoIKb21tUu0X730gOdkJZAtTP1+whhVh9kjLCRGQtU0ksQdateYTHJ7zcSijPC4q
jb/rITUvktSdmSUXXjgB7EVlc23c/2GwftIRZP9iNqep4jQaiYdriMni3EPqJfTS
Wwaqsuzx+eXPKbq5AW2wYXVmdkh3BVT3Gf9OFM1KTN3cn4S3fMHlhVt8WpSHpnuM
HdkdMpXvw4GJJQ+1QlEv7qtIjiDifnIidsOnQhri8a0=
`pragma protect end_protected

/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by DVMOp TLBI followed by DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_dvmop_tlbi_followed_by_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
acu92ErUdn1rV2BXWrjNpowABVpqf3MNVCRscawu1Nw5uSJc+0npmBcJI2d16VPS
cAID0M5rP/t7IBb6E4Sv+DxQ7iZRKFLYYjPIaCm48EaNiQRxD5558SZYPpsImW4I
Gp5t/VDzHhUt6/NZw1OT+FMZNx3DpMq+e9uAvH6reT4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 11637     )
DHB94YC4ZEbnXotQx0Z1dY2emHOtj14Wa3j1OGmOoSI9GVbHllrDIm4ZajFtwbbh
9t0epFItVwNvlynxGEce8TrxqoNbNDcqNtxm443mCDc5TjhIkvU9gJAhmOgLvDil
+P3Q4evVe9PaabXBFr8BWn9dIL9/g4VB253cIBjPjWdGDvtUmTzlDdppEBWGZsyo
Qaho0fgomSP8OwwAqDcIg4S7kZ1hbpmP2L4ozAfU3exP6jMk/KpPDOd7+sNGiaCb
7xay19Des2WkMAKfgl6HndADgKsFFPVI+N7H2t2j4ChDIXRgeNdfrpXQkWPiok9Y
ssgt8YPQ9nQF/EDUd3Zji2UbYlz3y8u7Sm7cqgldEGV+6m4QH9/miPA5YAyeN5te
oaoHgnkAAHbQHPUD3Xy5AaQwYe8jK53OFx/I1Do3iah7QrSlweULK0JP0mw6LKeC
kgkPSKm1AmGg5LVrA4BYxryliCqINEJOfJZVHdOLmEn4mAarFtz6cnCd4R5OiHx7
9eyDseMWjqQGxdYz0Xiu1lua7+0Z/zBqKLxo3eHCTsNibJ+3D90/j7IsKDSR25cU
hFgujsyvRn26RNLLLNEoweCDYMiCja0QFgAo5KEWUY2b+4/9GIDLODZYpYGrvm6V
zODZiaN3WI1d9F3fhKcdyn1qEPZpmxneicznBA1t9nv2+lrf3n3xAGuETcw/wWJr
U2GzuMTB4VS/t7WtZiD+3f6CrZsmi7U9zmkGvikxOnn4mNVHv/3gK0mMiAGDCvxB
wmG7pdtJsNW+Ojh6vH+OMfS8dCR14yVP5qzvflgUTv5XqLYQ47I+6mMmUlXSfpTq
dCKPAvEs3jv75tYvS3016HDlO/VAe+w7JfX5ETM5F3IMJDakUpN39BpABdhsEVFW
F32AkcJKniJj9Lj49UXdwG+/6xViOWPE4LHm5ROHyymFMeI62TOhSQoYaxUq3/ri
mpBRc/YFaQUpGwtAgkaLh3ttPClYSuuT64m/8hDU6W36VrMXGr1UuNKxxc42BYT0
leuNSwmwch49W1V8Orz1f+B6tJTVklJmdkgHmwgBJ0Xq04d1e1z26YDLZ3/tzOrb
q61dN7ptwcMx2gmig0LshorhJl8tTayxGDgWd/f8+HGuzvwceKlMnE6Qv0eaVwUI
DktvxGbv0GLS21qEZ8KD+Hik1/ckPX9QMqXknzUL2ik=
`pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     CHI DVMOp TLB Invalidate Transaction#1 ---> Retried DVMOp TLB Invalidate Transaction#1 ---> CHI DVMOp Synchronization Transaction#2 ---> Retried DVMOp Synchronization Transaction#2
 */

class svt_chi_dvmop_tlbi_transaction_followed_by_retry_dvmop_tlbi_transaction_followed_by_dvmop_sync_transaction_followed_by_retry_dvmop_sync_transaction_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
etFd/p/3X7TZi0C+7/rvxLW5AtEM9LCFkUow1cyOjHrvvtQF+xwy3W7pR2ebkmaq
tM9FEguL4XzisrCpsZ0LlomauGxig9F2vVk48N1PacjDNn5LIbWjLQnaHpw6jSq6
2h/CbPaODdL+KgHzZOTwJMQSXwlGn/zZUSPMkVPeAxg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 13053     )
t/M6WdqUffEGKu65qMlwBNUIIyujZUTKZpTGe5e34M91+X/usWrBQZZ45/Qbw1//
vcCmV9vXy5GVN7oe1OWHX04HYK2kZk0OMI/v6LE3tyIDgYSQeyG96YZH4DU+eI/9
kshjO8TZo0ywr49kciszAv69Bo80lf6dOvODNTAy7txIuiXnZpqiaRFYUopZm8SV
IjtEXWsHd1h4GwuzukssYNr6519TfcNz3lE8PFnuWT22CiV1c02bxFOwZhupx4QA
ssI2i2+NYwsssLMP2rnE34W5z3QJC5zm1nI4rhcOMjopmwu/BiNH2u65UgRLR/Gw
FGAb9Ebu0/CMaQkhnw9B7rAWFfe5H00zD89/SIvZj4hV8l3qjZRBlbPPCC0B4zmv
ADdbWHPYGDx1X80mo1k/N7e0+w1uIH9y2o56UVRvoR8H1blJ3OgSEv5vc+3mLn56
vyRzgITj1bM5nl02lyBDtc6bBrp1LLOtgc0OgZ1d1BczablrX4MktC+fq4dmye9o
sVUN8CbUNKTcd63lIDMls4JPMJq33PclXevEvCY+dXEsBhdEwTzOcIqu66ALuIVh
V7pC5YD2wY2YNGdWo9Bg29XKisWom2A0CaHJR9tG/Y7/2oqfRprtZFbUipUhWiIW
9jFrTCQkxf1WDGoMkV5ksprTtJlagWwrCQvD32rPpHhNHryxdSUSBIlPOj09C22f
LFwbZUjAanT7uSKUIK3SUzhc2l32xKiw60Go2Tku9qPSJPIjDht4oRCbh4QWu+uc
9qQTQkPvRYOA098//+dquIcez1eHX5VsiKMQoPvs5xuDEvq0lAuHH8RkIM+cVZYw
EmvhzbpaDxlYyekf+rlmggRCXeEalSYGP4+2elb1EST1f++mdcBkfOPNIWHybBvG
NOxdq1ihIHicIsDqFnWRM7F0WE/6kE2M1tO05k+f6Dsov0FuwEjIqyXDQUWlMJK6
ndDm1ZbWK45HOYzCBLVySPQGBLNNi6V6dkbZ+LXIz4SuPKk90JXPwMten01Hy8Qi
8pM6W/t03gbp4mDZMidflLqGalG+/T6k4smLX3hDNatbY36kLKGGHiEzfbn4vOJL
fvieF4906cDBCOiVq+pq79XWenHYrVyBT1eB220D0ztyOmR6VSxp673zwiGQ+flF
VtwHQYpAtyrtYwLgw2tJq9lawyJB7Dqxh+P+iizbU6P5J8Rfk//t6zgVZZBfyy0H
cykGAJh/y0DzIxfMLIIfFiDABS1+j7rdhrIeVg9bL8SDInOj2jWFRuTHGTSkEqbB
6pBBDAl7bExI+wiLiwiNaiq23HNJ9eOJ6g2su9nvVYZEi/c73yZ4uPBJjkQQPnjI
d8uZXdDBEl9jqCOpL+/B+EDtQNt6bb7lrqDo2d/NoLzq1E2qb85nIBt316d9ulxd
WlWS/jgv9N4kmv2O/3wnnxwV/tOICSL0hEQbKM1X0dQ7UJZ89uJSp39juEdwD9tx
FvtQ4Mpu+/Cf188slJWTETN9qki5/li4kkZk5U8QrBt7lrlCe97vQPoNKBO5lPhf
2uRJyttjho0R6fNDQfqopFiOtgcR+4QNc3SfUHRZn/CN+OGWikrCcj4u1hnu6J9Q
pIRSsUu23B6ogeT+23FScKi+Ei+6av2XZ8bOTZe80w9EpwjM9ErCTOpLJ1OxTvvA
NCjOXiuCmmM9/Gi/1w7i/8XcI0t1ADWkHpPnKDABCXqs3xIKdwxCOxyNvyJUkKs4
CtT5NjlmcB1v3zP3/vNgNpJNuYDMAjlWwA4iQenfIzWRAUyuA88gTDj/MjE9uG6/
gzmVW799Z6sgTxguJokkTqYWkkLnHjUymNSLpmepgjizN1lVgPFD2bnnX5wDlma4
67sJdighDZvGy64WFtMJrQpEx1O/APbFB2P+rZMgeIY=
`pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     CHI DVMOp TLB Invalidate Transaction#1 ---> Cancelled DVMOp TLB Invalidate Transaction#1 on Retry Request ---> CHI DVMOp TLB Invalidate Transaction#2 with same TxnID of #1 --->
 *     CHI DVMOp Synchronization Transaction#3 ---> Cancelled DVMOp Synchronization Transaction#3 on Retry Request ---> CHI DVMOp Synchronization Transaction#4 with same TxnID of #3
 */

class svt_chi_dvmop_tlbi_followed_by_cancel_dvmop_tlbi_followed_by_dvmop_tlbi_of_same_txnid_followed_by_dvmop_sync_followed_by_cancel_dvmop_sync_followed_by_dvmop_sync_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
aMlic2O7Vf2ZDDn/m90EJUxgS5YmN+Uh8uNN+GK3R9oFx/P7q3RrV2iWDszsxkNG
9AdCnlBzh+tEPTWLzqv6PaaP7zbPfbj6HWLRJESpQhTCHOaDHBJsUOmw5LCdnD4+
W+9QaSGkuh1cwnNg9qlEKmfL0ImDi8JTPf7Qg260/UQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 14856     )
Itzql+jHOUXDJ1/AqjqI7I3ORcNxkqHBP7fKwyCM3pTa6e9m9tFTCvTSysy/mqhI
ms3G1g7w0/mdWPrtab531fu/NBNELxwXPf5at1cQLI2fyHfc0w2oDkJmEOntTzYH
2Gmku/7cbeC9diIp94yLAahUU+R+IsF5Up+48WDZ17hGuzsCL0DDGO1O8TFeFDem
xNzj6ZLXBhZI4ElPiQBwratu2u/a03pdIGVyO8ltAEf0D++5nbKpB08Z2JmtffQS
50YCltxcQzmwNndmZticxOCJ6gXJX8kdC3ekSbEaeSxG+Xs29si8UI3xe9LiYYYE
h8HEco01RSoXz+wFR1jQIVs1Kjp01UOTtQJzCJ53ea8gl1GNoYAbjMfBizS8MrD/
P2gJIH5kNaxFMMyp/GVayC+nqUCdRahbNrHRIxzh+UG7LpNF42z1lfKgOuUKlxX/
FUUvLLGavPEUsLMbiN93uGMFJkUx70Rgd7GjEuBFUYxM5ujkLxH3bXmS21rUMozB
2bKV/uCz6JCHvGRYlzAFAlH5rjo/DIh2Nm+FSowdZaTTy1CySycKffpyPA+bQjot
/zcEdHycUjM6iDq1wUHUCyqpitT1Ibpfp2ZlHeTyyax7tiywxglKrK8K7CvmE1dO
fxKXaT8gYYPn7iffSW6z2nGTLDVf9kp39mO8fZjyMpJ6InFNUkVNjJQNowWPdejC
zj4joEW/KxgMScQePxjmS+tObR371VuBLnomRmRWN39uOa1IGnsr0fQe50Y8jDBU
hFW+v4tOGPrykmko7ZF28IIAk7nsftxP73cgI6Sz8LaSkrHsE9fNNVoJWOlj049g
7biuH3TBH3YHRzd9CbkScmgK9HlWcdt8QnoOmaQ+sxCCY9z3I5L4qEt6aYk2eF3J
dXS+ofyjRI0gN88+xF8NxwNU1qIA3Z4jGKUCQw95Jfy01vf8zEGFmEeDdVyXcB9H
DvtCwvmDTh3NfzpZ9EnkLdhk35qw6itncpFO8cmiqUCXxxhyLIyD0BZzE3xW/Jax
qXEmnuiqAH7M1h3Xmg+ExFLIVqBEdhbp31LQ911MbpT7sOKFh8IeKFSzjDZ4+VAT
22FHSsTYW5l4HDc65UISe6oVxR82pwyZU6rtn5R7pBd0sV3hX2X83fPxpbAfIAkS
PSHBlsXCZ/xpjtJawp0PRx2SjXpG9uYZiFEO/ieNktHz1yrIog9+acRAq2GDgVfa
CVvaX8UArgztpOhbJq9wRVsebgTSkPheWadFmf844FsinwWxHy75mnM9h6P+RP0c
RT/S3L3DH85z0b4I2l1O/64HJSLo9+27z0pLkzK5HcZUcDQs1RzU9WtunBiR12uo
LWiNTLO67r7Ss7FyJ44BSY+qOWqvMYOxXdWoqXHrXopYO5pYyPdHd3VrH+HIVlK4
oaOju4hk/KzCUMl2PBkMdPYkgas9Voct9RRX4SaqDw8GnXj+rooBRjtqchxP/Dum
baHlK5W7JVNxsTy6rxhCZmX1u8lQZl5r5hMHYgXSztbJtj0Zy7TyHMVZ2LuFwECU
6y4m1OqHF0QogI9iQPnYYk68zYDGxo8aWKZRFubulAYjHcS0W/pQhudTvPnWNiQI
SwgpWaRLWnuu5vpyEEIg3hRBX7hjlPC2fwyKVrBOdr034mIC4+2h1DENEEplVB33
JTC1Y2WdhlskW/lRhAQary/qF7sVHwHv+NYQhLOn2RGl7GOElRBU6LmrErAXf4b6
lKhEyrAZzJUZwP2dz2uXTJiAY5YWP8xGcA4eJbGYxqmExkwTboVSXMoJK3PDjgjE
tIaX1lG06iop4uhncwUsgyc6t6LVWqePLr0zA2dcMeL5xpxrctMbRv81olPGIzfx
wJcGiBGBR9+Xwawn+FZS+mFqj7PXRhcKU5SAa4heG2pMVvmouYl7UgrYuYJQR0Gl
v3dULWgrtEDeh35qxmWC2K/tO1/xnpuMhTALOuLX/NAUTsShdl+mymrxEg26IhiB
Et6c7Urtj8PJxpQ1BA3C3Tnm+XwGcfYP/GSPqQRojHvsCR0cMuQsRpPzS2VU3QGu
WOkJKdC0jQqxa2NZoI7uVxUKPOOyz+bx0/hotVpqX2B2C5BakFWQpnE6Qlx3Rtx2
bPgBezqc/SCSfo6D2GCcqy27x/69Zem79VnkLH32VCxP5oNIBkn8L50DTWx3A69V
i/JN+A4G52RLV8XmZXc0mPV5UCb4IX+YgMKNwZhZi0ki8mvd1RrPk/MEDgP0+6wq
SSc8MOTheWEa4KGdRIQOxzQt09okVqPEes9QW5+MnID+NZ9/S9/vEsZr23luIBHu
jthKBBabl2NKSe0MZp04zOZOjFSD2L8KFnzoi0is6m6+qJJLePQYPFZ4GEneyufY
RuzOs1/fiTTyDmy+pQNxmhJQcmAXd9McRdUSoUslkyg=
`pragma protect end_protected


/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by DVMOp SYNC Transaction followed by DVMOp SYNC Transaction followed by DVMOp TLBI Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_dvmop_sync_followed_by_dvmop_sync_followed_by_dvmop_tlbi_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
TVcnAL2kxJE7wVLiXppUcd0ziQQgJEsG+Wn+xlVPWcfBpNI41tW1B9GGFvV2ZdWv
3i9rm+UiFpAnY8NrD52KRx6qzIlpUTCMeEJ3ZibCjfyL5rJFh0BMu65GIBoi+5Wn
Y3QWVbq25+z7HDP64MdAkaTPQsMuqMGaUvIW69ZRXz0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 15978     )
bL1uNBrXkWCLwGnqD5Kamv6DE4usvZcZI6eximrh4wxNeOreiDfdbNnrOJG2pvct
fHmvjelgnoIKf98Hl/PdkNddXxi9jXtHtm4YTxM1y6rBUZbNJBbxKqWT+mj8n7JX
3qJTUT/aH/JhClt4pkpSWUOGtrgOxzkcIpDBoRKb+DqELZXlMoljljpMP053y76z
YoerTDrxNPaURHm5U+VHl0AMWEwbCiqQqoduXS7dhLL0UqKZMZ+phvh0xBwPK72/
VqBwkTeGvqO/1agH5uWir+2Fsd5AJnt6O0O8UkTEt9T/51XeQMbqM0G8XaFMtyTa
UJkePatMxrfcmDi7ki8re3jym+BHWA0iJjTFfSHatCB0lxPzvzIjWDb8HBu8n36q
SRiyvQsu3KA0HPosjHy5K56IDPpyjm/i4wJecBP69C4CuJ1VfpPlj7WxvtDpLhmY
sAWb5Hk+IgJhHkkoG48gWw1Cy1h9CNqrH6SgjSWeB4v5ra9eckGCL3FUoujFMUwy
d/vQKrcQRUWyDXpdHRUGN63NOvgxTqRScXayL32cpf03KB6vPHi0U6HiADKYRcdl
yvgV0sDM/FTALICBD9u7gOvI5BU26O9jUJCP70/UBEqCLFV4+7heO0x+GzgxhneV
b0A7yCzUMz3ZQZjU5Oq9OvzhtVWLCz2NlYKGgTIY+diAr0Onfsx1aBt4m/wqLEGS
/ARTp3kdgOErtDMeJoivP8/4Om8cG3PsL6+zqvlm0OFXYGr8s1Q9wrozsYzhdokc
j1sCyBOBwXVpSQiFkI/i//ZlAgCodsm+ij4Ch38TJ5FVH5ugkjPtQu4BeBykovQF
Thi9XHv57Me0qB3A11l4Y/z+kbGKs5V4xoFN6sxXF4/o1+8+bvHU2QjzfReBiHwA
TfemfK9AXL8OA6msRCrDRQ+2sEUSPELhO0mNrnGAPBeeVvpbcOtX2SSkSWXESGPY
8ZJqbFAY51w/O8QlOydgWAB1/9Rgnq78OYPGO6O65VcgPfyJGfY85f5dTnJZKY8N
27sadANwszU/k0t1F2PQEqMVLm2K+VPGMGCBu2ave9QYC8Ni7Ji8xYDA2rBhKj89
/VuhnxT65a1lco7OmhTOYID7mB5m1t1SbWIA9/VXyaw/4F8TAzo3sB4lwnaVyIkH
xpsV8lgZ6n5kS5FxSGVsfkBS0N1WJ6nI8l61Dve/rIbnP4nKUea/Cg+NCF1j1u12
t1TPuQyK2aNs7yz7pi/ax4PYjOc7kuxbM7eA5kT/A5HPM1T9DOx+oOPVEIAuVjoZ
0dhAe6fXdhZ/L8a7PEix2NbbqxptIKs89NuGQ0GaIAU/L4eBndK9TXXTFTUCvkWD
eoSbYI98czPeTmmB2XXPK8Wkq82ilFI5Sw8hB1TSbRDFg6XXS0V2xQTyG4kfX8vC
/afMS2xbeZKV4HQ3o9o7tRRJCykZ1QCF6ZK2Kkk/Am6BOb34F/vbbe9wd5rtrk6m
avRcSsFATOvUnowu0h+ZKnFrdTbQ5bJNIrMOizh4Tds=
`pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     CHI DVMOp TLB Invalidate Transaction#1 ---> Cancelled DVMOp TLB Invalidate Transaction#1 on Retry Request ---> CHI Non DVMOp Transaction#2 with same TxnID of #1 --->
 *     CHI DVMOp Synchronization Transaction#3 ---> Cancelled DVMOp Synchronization Transaction#3 on Retry Request ---> CHI DVMOp Synchronization Transaction#4 with same TxnID of #3
 */

class svt_chi_dvmop_tlbi_followed_by_cancel_dvmop_tlbi_followed_by_non_dvmop_of_same_txnid_followed_by_dvmop_sync_followed_by_cancel_dvmop_sync_followed_by_dvmop_sync_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Ac3hGiBOwEGqziYCMFNxrRVdJ1Ixr3F+z5/W64eNkNaZImIyKLFrr0g+gEH96KZ5
+VJw89dwT6oSLxVOZXMJNGN52ogYb6irFsyLWIr5yAgqXyj63R/0rYLaB2dlVEib
wdR7W6xayiaRo4z8fbD/FnMCCkHvoEbi2yt2/fYL0xo=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 17707     )
nvAJ7d93VVgyhemm+N0vv26PvmYyNIoOECyfp1c8ecgRMKeTfi7/3bjeRwMEauqS
HLexJrwfn05RJGi7MOQmcmrcuRFbcoPTflNV8uqLqy50cOGomT8S42cx7lhR8lws
tGbLqY/xSMyBl7XroPlox/XoIEzggmsxsoOBu4627Y/gTf4B8bauzlLdwB9UcIlg
eN4IMeG+C/nHd57xWven8aA298l9j6qwlNzw8f57xj2zCplG6v805A4LJftA1ZdZ
ug/DP5JiZ5nLnK31wpBx8rJFUf+VnM4eLeQY84DNiPvkTeXWT/KrSXpFQ4fhhDOZ
mIS8RpS94qTos/Wihrb+VfdFnNqCGZkjLAsdQwAYmFSSrSrmHUrUi8gS1m+Umg7T
mG4uzDv2XaAwtuX9uXqfFKq2KQoXsxwGsNmLUL+Ax6NhIzpxAdQG5JhHk1jKx7du
tSWQC7dR0WIRUa9i+PO8WoXu5Jdf3rzErbIIWtkmkkATn/yYFeQHoheCHniTAgMH
lHJjGnqIQLeEz6Cpb2GWhTi7qXhB2QQ3uDnhKkmB31H0AsCqSUkFVFl0P9WedLmi
1CblRdDp8q1E24cZyqbO1CHhF/1V0+vjmlu6WKMBuMmVg0q/p5998GbfU+4glAmj
d8STaq1785T9ezydi7Aq7xUyIXZXfg9uK42ckBtC+P0+jKTQ4J1repHuAIADwJwG
J5sFIiKgHi8kA7n0oWdpxu0HSI6R4X64nPEx5n/yC8N3e1o9IuAyEShq5xYbaKgG
9NjirHvQTXMOJHQLgo19L2SoL6Chuv10ANoNgU7zBsYqzpjYyYZHK8Lyl/9Bnqzx
EPnICBZ5wj9eCZsRIlLAmlzsIWlADYRNE5oLGf3vY1rdDF2LVbDVH9o9ktu3aNgw
okhyWqZ5ZsE65WHrzeCDNGd2wGcTbfLo6uwoXtT4mU3TrkLkMDR7n08d5lx6TcmV
3y1FqDEOSHRdVq1JGAW58f2rnPwlER1UimBO7+fHcoUQqDx30C1l+5p1yUm1MhsW
hJmmFcSCs6CNb0ePXbFCy0HMOaBRowMJRv/jNwHxXr9sxKUhbppwN/FnjNRJDfRt
hDbFggGR5JKADhMq4SkxMdfDQqbu2YeCRxcVsCwSCteqgRu46lo2J0OKmG4XrGmv
ZepLQ3Pie9FwUjNdhy+sufagtchATX4scI/vAjXGwDjBagtXC4VScImIt39BFWiM
tY3DlMU/tVAPTL7pQel1HlqFzLyc+Q7LwepkTNfmmAk0s0iavW8C8J12bUCD6op1
L3KJ+Wjer0xETJXEa3nTqESSoG6dQd86GIrlQKClfeAnVv99WlAoXujyQvlEj5Lk
OJsr/W8Fik9VW8sOpcTUv0NUTwqxJaQKEwa/pcNStt3IxwUdKW6xCJM4zOotw9FO
nMVvnNzHb2tHZDvbqR/H1n+MTdN4JcsTUyXcM5cOxWPupX2HqW31NwB/d8CNSEpv
vnvGXh25eG4kmXpwH9EA/h1pDcEVlJP115Cm7OpGr/jiA60dc/Ow1A0oUPmqtKv/
vkC18iNLEV7aCbhESYLBPh/xdjBZlAFOwkvSQ2JG1GDoLHS7QzTqMSmyzTjQ/yQa
8QFrH4myPwqKLeQpa2iyf/n7uYX1IOFYAxl0n/eIFltbZ7fEVi6FlScg/4sN5ZQW
wsmtnYHtBDnzZ3eNGN4y9ufVcU5LNfSqJ9bIYNnmSO7f2ywD4Gzz4Il8HN9jkBFf
T0IMv6O0T498qK9FINR51XcOF3egljibrLyOAEwM/RWwMau+ihnxqkqQhXLfScss
VuZlZUOfO68hXIPLLHQ8woQwN5w/t/ORbq3OkRmySHRNPohUCYYG0c5D3+z0vOKL
O1gRJQaLILL7Ul1dhF62mpWfwbc4Aug24QjDTsiMMeSUzcG0gFeVRi/VWRjHFhmd
RufJiuYUcwksRwDYvJ9Mk6cBHJaAh44PYWYR+O8kav3JR/QFzZqqctbb3ghgq63i
/F0l7MT257JgDJTmAkR6Vx5z8FrtzIL8v7WMlc5zcN0KRcqCDrOBgZZygh5pu7pi
fcNZysvz0Hew7Tnb/eanX9BcYpN4VNWNsNKYB3mO+kAtbMQr+nAjTdcd+VXfCymb
T0OrYd9x356Ia7f7XNs0WQgOYnqKsjv8evpBTS5yan00fh26Bo09fB6Wpl/xzR3R
fb3D0koeK851Dh/LkUQ9JnVJInpK80zhll3aJdQPhgOnjeF4rysdnt/EEwQap+uc
ia4XtGzvNKExqCNplT3IVQVRhd7JjAqe2F/JytTeApI8XOVxrqTQsBr6+5ywCtAJ
LG/AtTuDz8OR5QuSmuQGjQ==
`pragma protect end_protected


/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by CMO followed by DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_cmo_followed_by_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
RXI0xqudnxp6NGJ02MftOkoLcOfQmcSrJHLj1MGjftZs8/OsYkgPNXw91GqyL2PR
6fqAQ4/jcYGYQiOCEcgks6BNvWNsyi7YO6Xx+cK3xICLMI/k8zRugtMjoJnREgVj
kboNbtNYAYLa1HM2LQ3gsATzLivCz7vblojBbj1S1FI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 18491     )
0uJ+S4VUynnwilRbpUDkZNI2XJNBv4TKkT6xoa5AgGDkUpFE65F9O6aP7x9fbGEt
W08YoUN8RbRuv1WN+2tGzQTWwbTNS7PJF9DlAIwBeFcwyb+vN9WNs3Og9msSxs/x
yp7kXXIxVnV1MZUM77yhWFFzk61+ov0uqtndnTyulQFZNNZMJmCvqMBXeNyvKp+P
eMI6mc3qBe6mHi3oVbvAbx9Isq1pS/YfhukX1fsSwgwLcWNybLpa7VBmldIO40h3
eo9gP7Vc0KBMlH3Ou7ZXvlI2r/Lui6T5SSqng4lZaazfqEbdTJMUyarkK38IGhSo
ut8D3MiFE2D+Ocg9yHUxrBk56nEjhG/OGu5J5qW4GpTQUjb6tf+z7vf6sk/K+lVf
5ZnbV9vHd2uwSYahGhqxjufJpuvbeb40yGvac/TOiHYmOWAq9D5Cn8mhrVw2uKBS
Jkl7oy89+rBgWOZLZI9ACXE4LkLObzKUyKriNS8NZy1ktAUwRCA6ZVO/Prcs448L
bldUHgyHjDYt9OBMOhwUDGHNhkCLMQB9jEhgxvJTeOwxrUL66Dy7nWx9EaZYvOl2
h8buXU9F0RLLmcicE/E8vQcExaNNJArllj5zGNfE3fkRLzRqn7BQfc/dRjB81vcd
uWfx43AbGsiPPLv5pgoF/5GvzA0L1dv0pTVHuArlMDetNemTBoEpLIyEeGTA3DJl
0+MhDNucgDJH6aVieCxlDQdwJk7Cq3mEGEbc1Qlv1+9blVRbYJdiV5NPUfozvdYv
sIhce3JBZWxKveP1nbD2ErFDS0u6yk4vi1OjoWssfxy4hz2un73EIVU7iQ5wBeLN
uXnplW0HQUcId1Fs2xXDGJxjtWdUcRrfXDrJgRScHbuXQLzmyHEJ0WL6iGbF+149
udYIW2SjLm4lygLRdzkw9/ZzO9m1cpMUGCIRU1BKV47X/ahaqYhHuhWLPWb9FDSm
4e0YBejEDxRKzrcyiIZT6/IIBYrrqGSVKLjP4z93eTOeCHi+3+zbWmIpIEqkhBJn
Z3Vrmzye/6+RfHMg2IR2Afdr1yjGjbp0U/RlR3Qz5lY=
`pragma protect end_protected


/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by CMO followed by DVMOp TLBI followed by DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_cmo_followed_by_dvmop_tlbi_followed_by_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
hhcP1psRIWFxZd0xu8B5ytmup+wuwIvDV7uOuT3lzVKQ7Tvm47t2SZkD3mN902o5
2z1y7t0mlDa82rJO+O764OZ4T1Pw1mWCqsdUnj38ZkydIr5HKenP5EAFR436KmRK
ylb7Zzzp3FBWOkejdyFfsq/k7hahXuXQu3ErgGjZfqE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 19513     )
tHWaMkgOKNHxesTJrx/Ce07VN1S4qHpnEoNiFQV1lmKQjaF/ayq3Vidi7BjD7C8n
8SnwRfd2OnbTz41L+sokH9Xvhy6CKfJhlWCbFv9KxGPmA5V5g2nveP6lhwEcCN8d
qJag3p76+3qdlOVtoqszHqzAgthQyEVmp3BnKk1V1X5/J77DM2HaSroRSkCKE5Mf
Nt5VEbOchQWP6bj+mNllT/aY2O+HxoH039qJBd2TLYYmr9PDssPjXvIq3VZVX+os
XSNMUFWH12yZb4l5zPslyIX6Lgy0bPb3uy1t7ySifuWjucelbr/EMh3AX6AzdZ5T
h8RZv4WJ25RiYqc5oJoGRxikYnf1XV+SBXCMqiN+GyjHmBcgtmfl7LWSpEhwW/EJ
/a3tHLlISY0FSN3ZC7rp0U96ID+3Da3nzOcEhbISryaS9u0o1PemDjOMspRkqoIt
+AGKRUKUxFE7bsqjD2AyveMUAp9496c3Zzop70vcSyu2qF4s9pfexvbHJUacrqqt
8h5gqJ1ZqK6UqHV46yjh2CAU1uevj59pWBANkXlJWErT3Ry1m6g4heTivOzOk6/5
55D4VaR29BwZIg+lFomppOkn5Cj7Jhmbw5wDpBc0N8DDNr+ibqzGmTT0XBvQYdH7
PNi4k5SgdfblreB0X72LHlPXBe/mgmRnF8X6AiGkOPco0HHhehSjhmp2SsFfjiSf
9XumVIBHnuOpmU3trKsboOuoClkaI0bjpKNQ45moaiXAziP7vLgI8pS5xSgpMh31
XMJml34GjopVh8mImJ1hD1Ti6HVwb+U9rPHY1/BDjfBLtBVE2a9ixe3FLRXlQNqL
vhGYAM8OsKeOx12HPO2NyQNTMD54XHTnVnAgBrrxIy5HAiuDhj9u0+3ZUvhfSMln
Syt84TUghxHnw+jOLDTi7r1n08ieOP/kUVObU8mK8A8wjCPSzbolmzt9q/ax5mDz
P/oUGaX/y0gHUu/qO6l/PiuwG6i5Ebmm8gjdn5s8jYq25lLIcFdPyV0xXxRu13eL
9YeG946p6g6sWcCnTe9NHF/TtGOTjUM0tsB5u+s6fY1B6hEoZiTNGWQ1G7+3JAcz
EB7+9wD84KRL+xmozFRYy2oDf1BrGP9J4Juqf3qPFsNvyPdkkir8rBtYJhe3wGH5
8YS41mUk7ZjJ9jhJ03uGr4H/gmX+4jooXHJedyPvNs81DHDqWjXlSbxdnpc4aEB/
oBgzG91qao47b13rJ4SkOnRr4KNion6HYNtqGYlaQga7DIvG6R466hoND6UnKai+
QJDcfko6+wDjQkIHMbH+V2wSpCWn3Je03PjOLL0+5lJTrtLLY9UPRgeiFq1LzOKJ
/PHVcld4T88gVeiYmgKaEQ==
`pragma protect end_protected


// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Load followed by Store
 */
class svt_chi_load_followed_by_store_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
H35zBxW3WgpJxX24Ju+KPLbsypXkpoeeioxJeMQ46Kxw0viHKsA7EeF8Woj7w5vj
1tvN1R+RyvSxDdlDc7cMFo0n/qTnVubX/RipaCWVU/ApT2HFfoBn/Jr/M/xnJU6K
UJSutA9x4Yby74cQfxoGkB9PN2y1OecLbwoXjf9Z5RI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 19989     )
lDk50G9z61KoE1JxUmFc0xuTfJjijYEMXwToCFM4EslYCB4Z+kQlxr3eFmODRK6u
zsLlGjjquMtjE7PhLpHLgy3X633qkL+a4rE+I6qLRZWmNk2Bh4b7E6bt37qpGweZ
MjA6zpsH7AM+zdWS+aUf27dPRKv0534u5JG7ELnGHiEHR0baaeHt61EyCYjrQ2DR
zGdI+2lefL+m/lIX3uaXa5l9vAcMU5oJh2EH21LnVmDP0vQqrQAvaw5sdTotaplL
7ISV+nsjX+onXWI1n9j7juu31kZRr9L0cyXzBEqn2RtbnNYkT2Nc8vjuMbaWECyh
Dav4aZiDghSoYMee5acfFGjjm4EKfJed5a1j8oijSLIR/2FoGR9/L6+80+A1I9nk
clkhoXHcNFjXtizBWCtrcCWZqy8OvODd5gIlBHo940Dwk6jiobKl7YG2dYkoplWm
5I54Kgq5ydV8kvzivYKwawADXs3wRYv1BC1Ddn40WFLWaoaF8Obk/eu58jTgd7f6
y8KqwkozOv87c1HFxPV33GESwLUNSX+5U6AysBX9eim4M+pFc58gXyjMwnPIX17v
Rhn+t7U8mSd27/9gt6u99S7WE8m7eYBLnG9R5ThcKhE4LCT1In2kveVjfFugLSKf
`pragma protect end_protected


// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Load followed by Store followed by Store
 */
class svt_chi_load_followed_by_store_followed_by_store_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
PaA1M8XDl0lB6XeCWSOf0eDRpabLIzpQgV5llzxdj/G10DFDBlvHeJGQ10lacZKz
M27RvryjOnkYo8n0vwZkUXL7DHRkPjuZMSwcSxHfvHsTovojSaqDubUPJ3ay9raw
bab+d1iU6AXQ4RSVEOM5rzSLQutw2FWV60QWzWQvFMs=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 20626     )
G3Jrs5J+V1v/M3URxu/WcLsOCBVUGzqg8QCzsik4gmA2u/ecVhxtWaWH1p6dU8Cb
44GV9pyMhixeMW9XeuCpvap0dIsBvdVqFT1/oQpi0Q1rXzArQbKFv92i13l8d5/N
/j1eUr1pAxvX+jzw7aPjeMVIDHDGrWRzXG9WgdAaFn642wfWI7iEQuhf1hDNZuiE
1988akezkyOaSZTqrlbB35E6rqkDOQFFDFdikyUGd4wxDBJ6DXpb3eanAuVY/dTt
Y0c9i6l9FyaXbg7N5RBQTy/jXecoOGSq/mcsQl4QhIpwuM7YBY/A0oio/lPCuvmK
YSYgH5DLNOkE9c/7AO3VSuuJlO86kPprdvPN3FL9xqpVIIBXSPwN2xo8aC33kQ+h
jD58ojx2lnfdvx7jSnH37ZgCgG9Os7JKtg+DQFGlX5ihtUaor8aMp4KxOC/rhiE/
gBt8ScWrbri11SWbqYsfCvcp736R4imsJaCGx+DT18Lhp4EEYXQt9XOU5osnDPng
8rf6SvVlVm+nXUyBNSDuWtkQmewNv6j4D3gF9cgnQBO1Be1vZ7jw0EwHzWu6yXpy
6mC/FRdtr0n/F/OkjNZD/iF6dMETgQmocuFtHfIoGkbBlXOJJsR5oSR6gCvJUoiF
/Bc6hmiScY5DwsCeKMYCnyw8mUMFPRcpRC+3HoBIbDGr0jBXdJy819c83QdTWxyS
XORyoe01jqsjsRCugUceA8TN3myr2l4tH5Ta+Lu/lxXoFRvfOLOipFtEGYhJSpt3
jfXHBAyOJfQFcxc0z7sQoFVtJC0NS0P5xJKInxLg33xdlIBxsYbHRjFO1H4Pjva5
p+D679BtXSdbntDKtalQ/A==
`pragma protect end_protected













`endif  //GUARD_SVT_CHI_SCENARIO_PATTERN_SEQUENCE_COLLECTION_SV


`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
QO/DrVBIpfEfc1aOkmBqs1EmWROKnuT33vzb4rvqA8RYTTZ4UPONDMJMEMJ+n4gp
qyj1xoQ3OaNkB5WZZPBfuHPKa9ICw57e6dD2aRDYKK+o0buuiAx4eTtYIVn1akCo
8W1YntHjn6MXG3guI3tB17sIk6YBvfQqNetfiDvN3mE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 20709     )
972QCceQLASXZYX+4hjM0ogPSmigtDK3RBXmDu9v8Mn3L5k5TUaSkW09cXosWiyu
t9L22vyOHmN/kCmJRzDRe1M47uEUPX9ZQNEGrcHuEu4F9NOMSY/G9+tWnjTcAZMC
`pragma protect end_protected
