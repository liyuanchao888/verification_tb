
`ifndef GUARD_SVT_AXI_CHECKER_SV
`define GUARD_SVT_AXI_CHECKER_SV

/**
 * Class declaration of each of the error check stats instances using the 
 * `SVT_ERR_CHECK_STATS_COV_EXTENDED_CLASS_DECL(stats_name) MACRO.
 * 
 * Each call of the MACRO would declare an extended "svt_err_check_stats_cov.sv" class
 * named as "svt_err_check_stats_cov_<stats_name>".
 */
`ifndef SVT_VMM_TECHNOLOGY

//vcs_lic_vip_protect
`protected
[b=g2+.D[BabB.-cF[(K#eb?X47IHJ9VQDKJMgHVJW=2LRA7RAd)1(L4H.?5QQ<.
IFT;GU7FKMGVO,MTZ)ZC@KgK0)3VWeG)3HXG8I^80aQbb?0+G-aW7Z9:66=_FC)1
7<DFfg1d=430728;KQYZHR;2+bZeV>];QI22]O],BDcPc.O[#&)?Ig]+eUS?<)VH
@M@a,)0^Q>gX\6bO6]X:LNf,1)([8(D<<c5?ZONV.QVdT48@LT\@cLL9(<c\LG.F
dT?2+\JYI,CD800#91^d>H\0J@C+X=:aC9Of?Z0/?H[+T3I-XYDY\bY+Q_Q.GF0;
1F)^^1>UAL?S.ZUcgW=]_8),\Eb+8@A@=18c>(aA<<VaOT4J?UXO]Q<07>5RZC.B
R/_7[#Q[+b^BOgLY2^c2C\R5Nb.-EY]8;M#bgX697S0d\[J6#I_TZ0E3\1/1AD3(
?D#a5,5@bI0D]=D:=ORHUV_N^U7OG+[]<UFQ@1N#a-LZGb_&W0MGAI0SSF=6G7e9
47,#3(@593SdF@/+[4c8M8)08[=(&H[VD6GV)3\ZI30G3gCfFZ<S]XEH5SePZ@48
IHV#=,@#DN9-ZEI,>eU0bPe&R6;#^V+>0CaLI.fD1+^87HV2[.]45NPO(/)S04[d
e[&ROg/2C+V/fG\JbK7]Y#S]_(L+C/\U#f_N/9K]G[L/>:5P-0YBQ?1>2H-Id=HE
273IW[3HNS.+^JL>:4Mee7fC+Bf1d.bJ)LF58b;8ZZ/G;aN/Z15P_g(ME=A;Zd9T
UZEL=aUL7]XdDXX?S@/ZIZ]IV>-QLB6.K:(?R;fe[aY@)bGeF3bV5SegZ\1:NR#P
=5MV.cS#:I[_IK&060@94?:Y=Oc5&<7[K60,]@TH4Pb0SA(7X8WS62W\TEQ_.#79
Y@H]=U_f>N2?[A0@)2/,,Fg-HB^/<EcH?+:TCC?TD-CFQJf/FZB:8\UB5R)31@O5
>,Q40&2S?-F0W,a-/[UDbSHR@K97UT[H0(+2g+_?_?EUUT^?U01G^F-IPHeLYF0a
JAG:(N+SDHQaY<-AM,J#@0<>&\R[6:N_]g+PO5Tbc\\:3.RJ?IK]=QF#EFICTP[G
cK+?[Q>MUJKD>N2AH?K&PXfV-f3N6;E?/[,b+QeJ8^#MT1_,D7Ifg_/&P4,>XWP+
+Qb\,:Rb8<^<(:=GT9CKGe:M03A_ZAU=J5<OQ9MTOMSdR0D@99Z.DBASM\32.LD=
NgO[b8:aD2F9(@Y7I^8C.YASIY>EP_7PRP_8R1A/XH:BW><7e/KQ@C/Z-Z+_)0VB
G9I_<XPg5UGC76)[2Ief;65#V7X<XB.+aB?UO<@X4Ac5@B=M1A>@NN\.-1^S59-4
6e@]#WM\)H4OKOBQ&Gg.G,L+]=4797=3X#CAME=Gf&BB4Z[A&(BcWJ9<1+8#9]3U
FM:H)@,/gF67</_[M/AC/3c,4dD2M?=_N&UFG:RC(EQc+ZLTE_7f-#gJ18WDI0TQ
;-Gc&9e_a0e+Z/>O2c/N>+gS7WN8]b:\@)NRF?+a[7[VP).2#c.)6F&7>OK>^0I1
JC5Y1C0A6J)S(f;#,0N5W2CJ0cYY\:XS69W/3O3K;8d=0d3FO.9_.dA\5X#d=8BC
A3Y[<LOESGR^6S5\g_X6YN:3VHQ52\T>9(W+Mba]#N:9P3bSc(0P#-K1dE)P@LR1
U?Fb6&=[.HY5S.6C^H.:<eB;,GNP5Qf,68>&ZH;T-ZLR(LV0M6LM[&3bT&J@;.XY
AVK>QTB<K_ZSZ/#99-/G^2W+fG^=QK,W30_g1I&_#NM\9<f6_d+eH-SW4+26S_@c
2A)c6S^Of#bQWV)P]GN2[>UXO>,4,I]QUCZcYLG))(bbVB53^O;LVOW)545\2.Y.
RSMYcdR+eF&PW?=OT3-9BE],4W2F38g=,I^a=//1QA2?=G:R(EPTfJ(:I2C;fXJ[
@3@=-L7Tb-&(DHK=[Jf8G(:.d00OA\W.BFN7XMOJ7Z3IL@XTA9D#K)P75B]0](L(
+M&\#BE6[5C5ac0/gLD5E&C/Ab6B=4@X@C)d3/dYZ(Ia6@-W\V1SY+aLOT-3HUef
:9bE5EYWaR9FF-#aBG<PRg9[[T;NOSDX7,;GC8.ZRDQLKX5W;\RWAPXbfY,1EFT6
6P9RM7;=C<_TB8g-C&C4.7;75\9W6-aY#(?H;UO.E-2bY)/4#/C]S..D,@K(&?3)
_UF,4GFQJ,/@E:5<9EU8F+<JKV&1,L2a\3C^fFD1PeX#&3/FV>V#QM-a\OM-UV]+
BMd=J;a#;;:;R8R;_?(CZ:Z[F[ULeWeZaRWC@SQA27,6ZKTHQPeaE817.@EdQQ;G
SY9@,8_LN#M5<F1V<XS]Z[A3b4.(d9cH[c(I?6/gE\ZE>IS;Y5Pf:Q:56SG#@9V0
AUP[ZUCR,[1Xb]JX_a]^cV20d3V7G4=E;V&JL:cc;Z#(.6##[.aS6O?6@S&M?T;I
VLX^NOEbaFO6L#?J1gB/b7dS,53-RdI-SUH/+XEZ10B(^SJP6/ed@<SRZA)g5O@\
M):S1d?#KW7\d8;@A&TM<b<-G(e)-52;)<fN5)<gS+\D/L?X[R/^UN8DCHB(RcU-
EW3TR\Bd2BXPLZ7V3H[Jd)e&#VV855NaV61>7U5[9^\U\e8_a]\M.>MZ3W(20a[S
^A)S&I27[<A=OK?7a[I5eY8Xd&5OXI\(@QHPOB9(8c]T6O<K4a+dAXZH_=M#XU^;
M/E/R]445U;M\U2EOa]:#?c[>IK=L+G?I\M(X]cWMVG,,+1RKaR4P1-G0aA_gMDU
JPB8HN2R4WNILbOG9L85OQf>+/B(1Td.S+U_KHefRX,QXON)T>_P8L=E@B-8\ZJ9
7d38eJcTc1X4V8_=D/0Y&(9BO;f@DbC?7\(^_&)^-W73HF;c5[;)W6.A4.KGbEG#
POVI[bY/8#Q<\B)2T2_R60I8g^R:@FBg8Q\=a2R@?1/\_2AF#cdZ071-6P9VI0(X
AGVF&ML@f3-0Y7F;8].#8QS04/[Kg[.<dJ4cE/AD>+OEQS<f2cX/0J8VVYcH[G;;
71LV=cgT5;:RYb6SA[YX^9]?A9-WMM#R/_@#f<4G:?_ZW&Xc_\e;L#?0&B1YL3TE
eIVdGaU,:C&eH1BcD#Q&cD^ZIaGQ/1G9=C[AC.T++?CG>4IBW#AgQV?]NO3)/_?1
5UWZV(:)6R?<R2+2EP;JI5/@[OY8W,\gWA-[),0\LKP#^S30Z3+d4P).6UL-+ABZ
80=e]f;dQO\,P?+JR5M=?W^U,P-L9Ba98\gU4fba?=K<<e6GPaJJaPB[dfQP->P;
M2++OAe8XG[bX#f5;WBbYCV/aedfKEB)IGJC_F[=QecD)_&;QCe+SQ[WKd+b-b_2
HRacP&UZFU:)W5S(\YY._OVgX\TR/ZO.K&QCg&e/M]ECSf[5bR,&@e@7/HK:#I,E
7a<GB-BgBeT,eF3KP[\-aGb/K3c&\8TTM]Pb(,Ya0:AbM85;ND[H\]bHgN7dT_[:
Je7AP[=HYDE#cOaR6NLBF7R0NcP?6+ZE3M;B8LW8dM9LEg]e9\gg&?(?^NQ6;&BU
66.SPc6[PE8_aHO^832R)N>HTQYSSEC]9YNX,dc]0\6=8I.Y-VAd#UF_.IJXNB8f
S8)+Ub>LLP@ec[1,d?2Z\.T/@?LAX<bZPBa_Ud=&Wc#\#_71R_\<]4DceT>g;,D+
H@#=T6WcM;EI#b5A_Y;2EU8A&S(3MQ-05L=g+NS-gT;/K9WH4M&&:S[UQ9e(Ba.8
6R;:M:<(&>L,8C8HJ/[QVVNXYbfFL/;CAY/Z/+3gG9__KM1eDfUOX3^4]3>a(CJa
QRd<D5\.Nc3^.^U68a0,^//4WEPTO+^-^,eXT\;R([^2EG[+6[C,+,,PLGIJ&[Q=
,SLe?57O,RW].M[UT=&BE_Pf.QUCYOWZG&6S/SeXMa]M?]g.Tc2d<Ma;GS+gLW3&
JY?9F-<28)HZE^_CPS3F90[,E7_IL[.AHNE]AW)A/bPc=(LAYXIEM)@KWR=WEY=7
\?H1J8MYM;2:dZ_A?a]-&03#(fT20\QWRI[F(KMYP8F)d?VZAAMD)OLGH=8eK^Y1
3f-66WQO,]2HZ47Aa(9FJS<KN,0BWZ=gG,2X0^&;9:=(>aN2K#8,&I94fUYSUZY4
?MT/Y9eC-^L;&Qb<2H[8#GOW_eJ1dDZ+?fPeY<[5bK9^690EOEC&&XB5<>B23X-K
6(D>/DY<D>gS(2]J0G-7,L?G@O@a[NZV4Q8TW(=F0OQa?[?PJ2N[F2?\=JU^GZS9
+PSHa&b,4=gQK#8+gT7[4E^\Y::S0?AS?F5L5&Z:[7+5<KT9bY?R9_=C#KGO&;d,
.BOXNQH=?FV[gd54VM^Z?IF5HaOH:90F3/b)\?_ZcgaJ<6[OT[3#SV-7#+=3\Gg=
9)YHC4AgQ+1;/d/^.A/[85UVPf>JG4O]+QNTJd7Z,;8+(1ZA.BGd#N/dVaW=H&e&
XbJ&>ZGAPT5>Z=<9L,1CI0D>6.O9-\B\c0C\g<^M&.-\+VC/9<JYNQKJKA-bK?+B
&Na0Ie-(\SD)CG(Sd?:[U#25J\_+e6Ia@PK+AK)S&72PFaZE6@LP0#(3\3^A#[^6
_C8WA,cE?2FC=5O[AG<8#?b3DdK=3#WW\aSPJ?<]),HLU.Z41Y48dXb[EHbXW,N3
5(;T<aW#9R:XECaZS\f?\AN4TE81cTP^1M#V:L>4B)5/TG/^W/I8FH7Ab99aVJ?f
fD3NLB_E<>;d(J+P&SMEU2aGbC?GdPQ?QC9f((>W>b8e/Y[0/T25DY4c\3?/Y[+8
DdbXOfM4CDA65Q6/1/fPa1;D@3.77M>EVgJU4P:I&I]CG[bc;9aFY3Q;bD7]7=c9
F6938cFV5<6eBMX]KRbV]b6>D9<X51Q-A/G5DG_.DWPG]0@YIB&O#?&5G&0c1[RH
_J4MV/gYKK&;7d:@ONXSI=9+V=EQAdf/RJ7_-)V]a8>C\29Q<bAQ0GfI;/R/^;\E
_+@-ZCSN5^W;aXf)F(MJT[Q+_BFGGaeS?:cZ438f;TgO-U089-@Q5>CQ#:+Uc\)I
@Yb;2BMPZ6082+#V[BW=Zca.+L@YH.D,Qe[)9]XEI;3&9d16P0bIE>ZV-QH[UF,O
[?L+XW@\PWe&bR[fSEFU_&NE,<3P-KdC5ZgW[#CfH;<Wb[>+d;+/FGGVL)DbJZcd
@X-,,dV8EJI]^;/VJ.?bMYd?.A[ND.3@YRc6K=Aaf+bK6.0>3Be9E@E1Qb#V[0ZL
:14+:gTf[8EDf+@Ka/LIbHS948Rd5_JUH#AA0#PMZUQ_0aO1L,)09QccO-74E5IX
N^b^7#:TW9dEGIMSQcW_))TW9W9+[>A+S.;-WO#]AK)9W<eg6U\I5BO0U#?>?8Y;
Q1Ee.OAGN(2M_aW:4K/>4\H/B&N7.D\@4AHN1\KO3JeFZJ:08A,:B0Y9Pa:07E24
XG&_ST.?/,LXgB[5GG)c1)>OS2M/3T:eZM1;#@E_V+O#g[;2]]eK#+QUDH:,?S(B
/8TB2.TXdL_X4X1KGC^d-+fSX&?fa;#M,QMX.+Q=1eCHY-f=M7_8EGS6S0,@cY#^
:gPDZ)^80OO2EgLWVb6/P.ZN.[KTQ>,1KPd+\NQW?.^Z1.R7)aQA&C)8Me3TV_+S
caFDO,9^PPG+><)bNKY;L+/H76#A]K9LP);aCEO-/BbY.7U_^2OQ=5Fa(I&^UNVf
<C-1)c5-#K<;8EaA7g#7AOTOSf]IZ0K8^S-2_2ebQ[e-5PDTA:,<32P5HI\_B#QG
1C?F+]=X(\+J#a9FOY\Q=_UVYGFN(Y@._.@e(LG63B9AX0]Y]2K^NHJfH^\e0I?(
gU1+^NTQM^-e.\^0TeYPE0aI?=Q?VUecG[6=CKeD7Z9RD4(H-&7d/0-(fZ&e3/7D
-FI-C,A,U8OK]CfC2)]b24.(V;JD0JcR2AFG&C5HXAMT#?a\,&)(I3CU#[V;a)_+
OXZ9EY@999&Gf8\]P^Q.Q(PZZeZF0?>Z(bBB)a99JV5DL7VIJ9GABd8_7_A4]HP1
]Kc15V288QH6YMS6PLZeN_8F+M99deL/)EDfJ#U.S2f9.M4_gNW8(XWR4.fgZI?f
<7\<L1Eb0I(I,@8J=\8R#&J.V_J/U/Uc+2,BB>YS:6#ZHL,-5Y&DBPTNY=GCNC;T
RR^.0X+Ad2@I_+JD&/0@1NFERN[)9GZ^a(gY0DUDb)H9RRT<+QKGY>M/,AHJ_d=[
)7OeL?,e>D//#MaB,QA/)T9eM\cOKUA,B+(D7(aX:;7=09H8^]JD\U2VAAf)F9QF
##8&HfI55bKZ-Ta;eMO91fPH[?<VP[,/_@CCde8A41;-2YLRZ-LHC3EU/R79b)2[
YKX:L/bFS?8O+YHR>J8e^dBAL.9@4O#J\27@.7I)Ga2=0O8ELL.W,H^NM?4:gSUD
ZTff0A.)5]&Z+^176PP@P=VP=@Be<eK6K.31a:&6Qg^_GE#8AdO/&2f:<)PDcH-G
d98Y7gM38M)1Zb9\PX3a^B28\=VL-D\+6&)]RMBAf<UBHDb9UGVW:@0_N>I(7<dB
QIVPI/QBbM?>C/2.<1BTgJ@W&>F8EO1-e-SU^&696OWSN>^a25+b-F>7H(AI:d^,
69(cEH=R,N+NO.PQ&=9Pb@]322@>3_g)WKUBE:[F-EBb:X<82ddQ?K[4eG-JWe8W
Ra,)=;E^&+&[D>F=E]-YY&70>C=11]83gG1g:R=7E/Uf=[UeOLL105(]cBAI22TQ
Jg-X4^Z6J02>[WW8aGeS==P#8UY>1H\NQ]PU1>I3.b\;X&fEY@_4f/U16A4]I2Y-
/NA9R7]T1=70X53W[[0&V37TeG6&ZR7X8bG:dTe&O[2F8Ff9C0);DbC6KUgBCa9J
T)MGBX_;-2;<SAUE(N[b&\UA)bVUQ5b1bDH.Hd831.eTQQeEM[&FJ6\?:cJ;+eK6
SN-O1P/2(=-Z^Md^V_.3>2V1+>.Ze]U,COF,C7=180eKPON&6D=E@]LCHJ-Mb8g(
aWK-X8bJZQRV1aUH.+Ze?.37gGN_U,J.BLE1e+cM)3ALP9PKQ<I]YNIVZKJRK9dZ
C[?Y6\RRM4?]E9T(9JN.7faI8c85>VIaPJ@RQYf-6GSE=8#2R&I)GWJ\D4H\>BP4
FQbWJFTT4YgZY(YKUFL4)=0f8I<1?)TPMX^QKf=7(+HH]([TH9K5?^(XZ8):e,QQ
;UeG+[0fcJ&\88)=<JCWW.cbQ2M;0cTPUcKV:B,-f)3LX[E9VFYSA1J181dM<(\7
DVGa+65?2O(?H_G+.[Y4T1gT2(M@D4I_=+NdDYZE2BOUbIdgN7#[^e:5MZb+aI-B
@R#-^;42d0,eE6]5_#/^U(Ig6.C&Z(0bKCO4a4V8A&>=AZ_bEP+-NTbXf:G-C5Xc
^ZSZg)+F.:;[_/C@cG-A@.?R=8QWJbe];7>UA=RB\bY\eT+DFB1Fd30G4-N-;S9R
eee.#HWITY5_\QOeA/QE3?@1&)>@>1P.dD&IS8++fQO4VWBVLHbI.;74@5#WOF.G
aFbg=^U\EJ2YJZ+daTI,SeJg.<IA87,>C\JAa<:29UTC;GG_Z0TNO[aSV#1THCQ@
<LM=/S6;G_NA98RH7(3fNN_V0(3XK],;^U\6O0_JVMN#Ug#TaAbI1-/2/cQ._P@1
V),V.@Tb]5FY>Rf28)cUB62W==V;SIW;fBNaOKCT&^e<,VQKI)_#4c?G,7WPJ<.a
6.6fX-Cf50+Tc5Pb30=VaT=3TTXb,=A(b6-5PD^Y5X]8LKT4ZRVg-3J-<<7dYaOG
HYc,R@^.VSXggO7Jd06J@</.HDa;,P\NJ[L6F/7gEN5]\T/;8VH4IO3U.5Le\aXP
@978SCJNG-D(HHcUW;3>;eW=^55:+6^WH[+U-17D[a2.?4AXNBSb@]S<(OP[?N8@
\Ec?NBLg_OA,fXIQ<[M6IdYd/H5cGP_[GDa4.bX^<?N8M#d@0@aYHJ2E-B8PfP]Q
51JQ^/EC]fYRATb/f-SgQ]\CGfbWZ20VH55bNHL6?P35AN+YY7:1,ACRTWJ,V&5T
U&)#.O=g&b+-@6<^W5gF@WT.L&Id/g=\MKX7\#)5O@<>eXWWPFI8XDSEI#3WV2)2
6RGc4#M5c\^0LB^X(J3g5G^YB>D3c-X>=:e;HE]B,7>AON@-M77YP;A@NSC[c/[E
K^PORP2GS]/a@9)Qb3=a]V<79+f.#<cUN2d@4D-aT<3aD./AWWBM)SEGN90AW\I2
T=.H^a+2.#d?)</RKRQgL9M:H7dB/QXU2(P7L+GN@e@0I_ACb(-<T4P-L-8(NO[Q
.26Uf4X^,g0BYd3SV@K&EO2NR_#4(KJ1TbFJD&4#B?RA&WVE-;WHTSD_L?,BJ@+g
9/ggS&F?M??HM]8-,-Z:NK>/)b[G<c(P>U\=d#4+\A@CCTE#<_=4BBe-R([8ZJd(
b@g@2YY(b.PgB4a1GCW>ISdR-7f@2DQ]=2#?XIcJH-.S5B=F<BO:V3J8>+]TV>]<
:>>eE+99JNX1_)(6JD3B@I0E^1V[5aL?:SL:J()]dfV)J,fAY<BI1()VcbG\=DFL
\4]ZXE##ID@\:&OF@L7\Z\2B509S_CJ=17N:\NA/:IQ(.#KNe,<KLYU-DX&:DfNV
AAZ&#f)c8V2@6YAbc^&=O(I[(S\91?=cM>#H,@D,Df35+R(GQ_?G5e8@50SdW?<c
KSTJb=H/Z+Rea.J=2?/FdGRDfU4[Ve4_@?eLN,^SJPeDe:VMV.41\&DGU._A-WTI
>00T5S7LP#4_g4NV>O.1=>.f1<bLAf,FET8QX8P&.@H\\IWdH?Ic77R&28(cZM2f
&N26O8D3<Ub&5;=LX9#-0_6,VWFMd\--RWC0N_8F(=JFLP;C)Zg<d:9YL&?X5ZEF
NT0Z3QW#O\KD73#ER<-F&0L?#[@6Vdeda=VN:3[3ZECN;>Pf.cI4aX^\7H3>cCZT
FWE=Fc?[7I&XT<.3GQagS)J\/J:0&.U(L_G7g8e-_b>[B?,36_6f9:EWY/9:./2\
Jc:>R]62:;8]5<TJJO+1.-ceY[9L[?b>2P[.@M:;&Z+bJ\CZA/K0_Y?OIC>-Q58;
g4Y(C^1XO]1cFH)RIVKQ0SFb^SI&JR8g\IUW7H5Z@X#]2,.dT_;GM?b=L8dO>cT]
FW>G:[O=1Yc.K-AE?0)+WYYO,W@Y8^XX+T,,O/NI8,D7Q]9PH6]Z>B?b=L\^aa&M
:fF>AP[^.c:GSN\4a\f;/3KfQ@O-0/78C/UO=/?Q8^DTW)UM_g5P?cA8/fO>N36;
]WA>Q=FTJC4=a,gXTC)IM];68bP-D?U^X3-1?A00KX0]5ATXR+N@-K#7R[IFUEfE
aMKOFa(+4,496CIF(/Yd;MH15]=eJ:#:ASMGeENNfA[Z4/M:+<bSGPaK#Y\A3bP4
@LF;S;;XM59#IWU#07O4FKbc7R5[f^,_]4_BFL(#P3+.Dc.Nea\(,@YFE(S<.aVB
MQAd1cKBYNS+;Z\IANI/-<0+I6BN56[>:-KT>JQg0D.b3PFc=[+X=8MUAcdG.@?(
N4K+9Rb+00])-5fA:@3IG?Ld0I-GR]LNdTUS@)>Tg5\f4a<GG6WB5G)S,/E;,E.<
@>MYecQeJ17EY=bG?FJ\2PXN,UW-+K.K=a#Q[bb+PZZHPAM??@SR+3;CeTJ[(0/)
SC=,BP1YA220+;4cLE\)^/g.,&H^+4L]F(6:gPF5O<7#=DSH7;8Z>R6K=-_g)a4D
>D?G2C)aNW<Z-Ta.g>aKGKT8FU2.4C_&V7G>J9I24]7Z3:S;FNSNW-O50C7183><
2;,\V];>GWA&96H_1#,2[2-N0eO2\93LROUHVeb@2^[:.O(;=S>5G07)QUY065L^
+fgAaRU9f\]&Z3=5S@2WCa)5FZb8bFDIL\5N#GA&0E6IIUZRV1TYHN;0Bf>E21Q>
1O(@-\He5J:78Ge_Bffaf+bCgLde)\2(N=d>;TBL/,J3?#g]IJ0:B1^/1AFKS.d;
0g3QZRP#bS,YYY^WR?TO&@1Ba@eC-CR\E[O(S#K.&^ZB.@GM@MGIM3;ZY>I]8BKe
1:g^>+M_VHB+6=#0fFUbBH[gP+]28Q:a(OaHB>a9&U3HRYXES-8.^SGgZV9Q/K&:
L^fVCWN?eFI6^;Y3-AQ@]/2cS#Ne(e1=12YW2,Z,S/9\Z<Pf[5CEb+5H81>P/.:a
323TXeN[2ceXJgeB7_+-]74(^@]7=P>A,)\<<&/PO9e;YAcQ_^c(U\bf6Pg/V&HR
?HE1VSS.bZJ0-G-[_9W\VeN/0^&-#U?OT?LPU::d_EO?8a]+eb_F&CQXdA,^B-_0
2gN@a6Md#]gH8AO4354V(@Y[f+A(B/3^KVD-(3A.3=.9/&T6.;4>OG4#X]3:-EC9
0<9RY9?Oe[)#6S,>HH,YQ1RcOA^^Igf:7g5?@<FULU27ND<6aM4cW07_DMFL63T2
aQ3=]-^0YXM2TTG2?R[B?E>2E-5JKgb4.5QNTM.TF\SRD3\F)8/5J+5U5gcSZ-f#
FDbPg:,:#GLPN_1G/V^dPFJa@agNHNO)5R(4b9L>U&-2IHR^fGEP[<d((YSU3EN\
AfWI7O@d^+7]4e)1=K-cT\TNEL9gK9O5257C.Z&5S6eJU[CRZ;+aP@edg2bL@Q:.
E6->1L5@<d24PWbYGLNMXQ(H;cW2^.c7ON_K2LVQ:dL^3-OCBW;d,_.Z-bFE1d=&
Q^&W/;d_\,A+\a\<DJ9M9-B<ABa&[;U,Zaca71ON3DPXA:Df8[&+?GI7fXPMJY_F
ggR-GG;8fTfQ+E9eT[MBW==EA1,FIN09\P\&71HT>3G.IK.BE+#+:V;7FPX0KQ,B
.,8O6CLLO()4Y,3WgGd\Wd_U4.K(ZbCZ/\QHf<(3?).Q5N/[HP,&.L)Dg+X#YB;+
U]#<5E7W]T+D=[D_SWOZaTUH7b:A&I4,bOOA=J1Q(R]SHRdP)#Mb2Hg;9,:;5MX?
J7VMg>FBH@?S/64):1W=4Z57dc9V+T0Ze;][&A7?TO_(:d>=g9=HYbcQXHQL<8[.
K^9+=-1@ADRJSY#DObY(cJf\I/WB7d@6,49LK4D,4&JDC;K.5;P]#Q6E5LQ?:[f[
=30[BZGg+g:L>47(6OJSJJe:R__V(YXfPWfQOXY=3Na:04F67(@^/1,127SDK@L)
18B\=TFg/-(PA#NeL9e^UD:4aSc0LGV>If\2KNbMPV-f8T\X6BX7bK,SR+P(:(X&
D=Ke&,9^2O_3e-J8@V2BW5\Cg<)8IDY>Af782Xc2LZGb#b,E>0Da8-PdW8?]8^]Y
V5/_-b-F&R3NI@3Hc/I_I^G.J;07Q#dT4Wf7Kg-3IXTcN.PY,&+[R^c:eC478QZ<
0/TOS486bG)ND6VO]X.fZ?<b(SJb_A:\9E1Z^T=G2eTXEQ8AWVA8)27[fd87Yb(e
#Zg<Se:&7M/[PMD_d,R0(^5C_g\]TfC.AEH;<DZADR&/=WJP\4:f2@d;;;#L3O02
[a]W;/IZHUBg&7\+aE-fS:3^TLH5O]0Ff]1-E@#M]07g0b==:@d1:e-#(YPN_#<>
#T6U@^(E(YP>6M?J0?aEQ>^P++;PX=Pa(aX;G</S=SI-7#egDU9/@H=CR@:_O9F^
U4GY>:/U(U^C8O):Ac(Zb5DT=#6BcRU02.X6dT0gE5&RJ>8^Lb,/c8LN[Z8?7(4\
PaXHF_4WQ7QO:/C+PZ#&/W;gZ)?FU9,TaU,XXLK)B3;BAQ0bLW.a);bdP8MA31[Q
/fC^0,/M5c8A:&@4O+QC\cH2?3^Qe&=FF,YfUX(f41A9D+?XLFGDfaI[Jb[Pc5Lb
40K)#M.+47bg:Z#;^&+ga-b-WWYI+D^+0:[d,O:Qd\86]>#c[4cK#,/GKTZL:,RY
8g5@ZS+;gHHU9AM&,TaSNTd++8-2Q2[&a5;;4OBKG3;W.+_@?;JK.Z/a37fLcIBL
QUB:F@U_N6\L[R^-9,eW(Wf@[b6EW4U;VLZ.M26)f4]@KHF2<7Y5Q.)?PILAf>9K
>.4Q\RVTWc#?LK(:dU7eRF0MZ2@YPN(CR1-S3]#b.D\R=A_9XR-KLY#Z1dF/?:N2
AUFNcVC,]>U#(.dM>;e]BBLbH?;)8>g(-f6XdNgN5VI2&^(ESCM4;W(JgaO3GSIa
9Ma9GA_X#1cR1&ZF40;?ABf+E_[UJ.[[7aJ0FO1HcTJ\CJ=,ENV)6F;W&,b\4D9a
e,J6e(4(4+:>K\E=W^)O&ee\55QdXERaD;HCLG[&C@X@MV_4<g61J19BA@eSCW&S
4:S.eF-e9WW?:\9f2H?FK.M1-/8A;U8QFPWXMc../;X;4@(Z8AF#QD+&V6CTP<\?
32Y5X8DRYHOJ<g,[^:7-2-^1IIF\#S=W>=XDC8IY2(,#CZ(5+NR,6/H[#:UN_/;^
5-]/LeUOFX-?f#9O#^]H5EgSH4O8X1g:=U./GG8J?Z@@BW/2YJg13M<T;1:O2TAf
(F2,9B7OR,MYUdS\Ec^.ZO9.eS@5/ABS74<;f/MHJJ^KWN[UX:3U4HGa2U4daK1B
D7+D6=Ic.LP:YbdG2<#3MGDI1.KDQSg,&T496LWVEU?.dA(;d.5e<](4f[3d.DI/
ODcY?4K>e]\\fW30,R_J1QbS=#>0ZUGL6L8B,Ed0BO@7RfUeWWD:\K5>C,HKH#=[
LVYB2ALAPG-SKG[)TSKNR<O+ab1[CfFCQFa4[Hb:f+WWYG^[9>HEc>SRU)b04[L6
>ITd@>8_)(c5gQ]J_Rb\?B4L:Wd?E\&3f6EU8GfF3Faf8V&90_c.@-5@^<>;D-WB
?3KFV-(LLQLe5B:<4[?+;U=T[/4LOg3c0?Y\Mf03?3-ERf9P9D@;:A;@99+=1?]\
&CTBB<D,)<\<T+EWHYe.JYR5gS=0\-O.TUc#SN;MX&K/a?,\39^V_U,QWJ0S3QJ;
J@=(K]eSH)P;:Uf(33]cYGG;]+JC3PP0^)>7>X8TBN.T-KPJ&:#5B=^7gW\aO&Da
RGYUA+&2K/^:0/[:ESa6/Z<N55R)9\,LV9Nf>3GAfLb[D_3cCU_>T?KI#S(F^L<2
a0:CL=NSZ-+G>[GN7BV99:b8AQ+9J_aFTN#\BG8c3,_=/Qf9.=H]ef8eFGK+Oc9V
>A,b84G>S]?7F:XJKA\A2)TbdA90O.8RXSaOZJg\3-YLLY><E[<Y_)(7bCO=,fHC
1G>]JKWbBFTG#SAbAOg2)VFc<LC]DFN8-.HTJgE4/9Ud7:LgR;,3W&bXR-TH4IW?
W4.AZA##7efH(c#V;(Q^ZJWdabUB7TbEF&0aS[g47U4#I)SfUZ/DHJdW3cS(3=^4
4T9HSFQ#-X@9L(OG,.+=F@YWNUHB2K^(Ba>^fR=g4KN\\YHH5L4:/7^&/=&W2I-O
;BF-2[ab2:@/X?-^#Be0N=>MI9/7a<R)LZ?8K61<bDJ;VQ,5Z&?\ID90L^e)MK:)
/ML,3J(L1P]5aOV7T;O1[HXc;.b/AWDFN-7O.0]VY4V)bC);??BRK<>8Q:3bQRB4
O#f77d2g/AR5-(8U)#Q+#))#b45HN6TYg]DB@LPF:V:H8][fdJF7>\MX,Q+gP>VB
e7.:(T+;M6^@UK++9VEW;SRG^g#+4C+>:KZ7g0O0T,g2RA^0,D0VJE>CSQ.4RJVE
GY;?I6U,Lf:#Z2V-EG,Y6^@5e2WA]I/7L;TE&SgQF+=[?6NUJ.6L=\3+:MY41Z,b
\Z,cY8YI]=Y4C73H=3P-;0R\A(6Og(.6<7A?2CXb]^>V(-:gU3]1IAc[Td<La[V2
cREZ#Q5ZdNZ+E6NQ/bQDS#Y8+58Y[,^WK)<+^\5H46db8TV-P&g>A1\f:e3d//eS
6?-#@7bB/[L@(d7ZYYCf:gGT(2\I:AO,P179e/C?GS0-<DH..fNJ(4_cLX+69,?5
<I<Q2+F>^dd9)6\?5LMD1N/F-K/1Ca)[BI:;0gB(LG9^VL7KZ<P6NTE@G9OJEYK#
X2W35CgQ#W<8Gb\7#B>bV,cWF9Y7C72T4IGHM0Y592.71Tg4UA6]0#MTC/eZZR=b
/=N4Z/,VAELVJ6)S[<;-3(6fY[4F8V&dGPcBB]\4G+dH^KO^b[^XQB0c@GV[OJR&
SfeM,cC#7V)B2He1bgUU.7GP3ff4REH?c(gLGWBWCNXM..XYbcTfb9dK?R9LD#CD
D;3_^31[(>e<V&=S_YU-_2A(a+a9;:QS/E,IUQ>\CP71K7f6a@LgdW;N]PPHJ5Mb
Z9a=e:3c[8T0FcLAdKH@(#EX5>#G[dFg1R,<ZBFE1F-ZHA,1R[L_fM#?)d.QX09C
+G.c5XXWM-:JRZG9=\be^A;T9aU+Q.B0EB5fW_-\M(/CRU;ZNI\gC2_(P6R]F<Q5
J#]>e-#D7a@\513a-O8VN&:[_?A9XPfALZ_QV]61EKOF78f?3+NFZ,Q9AS<f+@[5
d;[A/2[D1Ib=(#dOg?T9EV;8JGGP9SQe0(6ENHdL4ePB3fFg&:0#JMaHG.2T4X/0
DTB;#Z52I48@&9?:D@\EZ&,e102:20V?2K)@0B7f>TB.VV-M]5G+&f&?b]B,RE;D
LY10O&Uc?Q8Y72UD(=Z=):GKQM9?-P[[HBe04JO4e@=<f3KXW#<V1dFL7I:,dVN&
.3Y(077OQL8@-(9-E05NXJK&:S@OZYR<,V&O@F?V.]a#F=)G9QGXVJ?U2dPe,HeK
@f7EIcIE3/cX3T+We^46Q_NH;BBe-SQWaKU2GV,J[)3MO.0@e1X=BB4FL1-N?H?U
6/Qf)fa0fY^L5:O@b[9/H^,-J2B^E,b+]&R33.VV?N^P:?=WD8CY8[4c;V)/b149
_&30Q>_,-F(G-8D;&):?EW0FZK8M:W8Jd=2XJ&9Q9Q(eUEL+E2DbLN6^SV@G/JNF
O&>Q^D=6WfHX3BaNJZ>UXd/Q8]e)818CD[fN8^e9TZ#b[,M+(O=6#g;/#TLQeA<C
)gXO@.M>Q+6RBa[9JgN2YIY:@4OX/F7=SJ<[.20@EXB(<58,0EdafDF@-4:b3Tbc
YFgY8-]I.dK;f2A5MXE@A592Y&B6WP8[S\H,d)MZXILdSI=0Wd93?;YNNO7V6.DU
K:LHQ3[)Z-1N/,S2>9<X=ZdC4<V@97(7]<V7.g2gJ4A;H#]9S0V@TgS<?EL@(Ia6
DX&N?(X)bXP=4\3.M9#8OMO89^g.TIS<C4)88e+GgW3UCN.E542#_JO-G@S3>ZBf
YB@:#1F+=[Z.SW:E6.b8QGQX<;J;f@bf-S-(1YJCQcE+(8Kb/?SKUY>UJ)H#WQA:
BL2UMb_<8FTOebfY+UU>^I:VRPeZg5CTgfLaY94BH@eA7/K5ZIcRaEf^O])72bP/
MT^B@&(01=XVfE1CKD:fNJFS[(MIXI#baJ+Y;<I05#Z1<ERBFD<>S8)O[CJG0gFa
bf_,--]RQA42\;dKPFGcg/-A9ZD.8DU[85TNbeH)+&[cB985)SJ<Q7)Z\Q4O)<Tc
>GQK9?eU\PX.2c#)V/C_c@Q2Y?X;H^W3)c^g[Q8//b-,3/e[B^bM9O2d+DO>-E@B
_^@574D\ZG8A7/^UH6[?4OX#EP[7SX6\@eZH5,d<3&d6Tg/1bI?0LH.:7@/^/MOE
BBcNN^)aSE3=L03><2/:HG2V:-=J,)g=1dC;+afUE1CIP?F)Y;dWF2T/KdG88bU(
EK,)6;PX/f,dfL36bg=SUAPYY0L)VS1@U[)3T&7=?#J=9-GRE,(c/&#.+<0+V<H\
+P/\=KE4c6EM:&9SCKL3?,d;>>5e3Qg@<8<^SE;Wg4IP8aRW9FY:Z1+&/c/^QU?<
&?<cSMX2.K]cM)F3WP]5)X#&3@5;TV7/F4>D=7<(;,-8dR;:KBbF),_KW82g]X#9
1c0.gQgd5.-IDg1K@D2@A;fU?cFEHN#GNKX4<7=X/(N;+beVJIRX=MXCW#MbGE<>
?\b29+e8?_KT&QbK0dF0UFO0D#H+K.CVg:?GZ.JBYOQQ[&5,=@U7S]+C@U#<EKE<
bRSLV/1:Q.+Jd4&_&P)#\C=UHb5N2V_+\EY#^Q;J6CN.GaWf3J2760>05KKbY6YZ
NADW.]&P#);V^G?R<V>7P:TE@Q^R-fTa?,-FYKT]>8^_A8VAI_-=5KZg@T6/5+)g
Zf=N>;19V[Pb,+T[Qc/Z(18\D5U/<0O<73.EX(Q16YI4=8.U/4+>:WH_4eFFZ>7.
Ue.&R<g)&6g62J-E/BY(F6a^8MIF+BD@LY.gYe&0R1a#ag3)VbCB+:WG\T;1A>B]
7;4RC?ad?ZTFd]2+I9#RQNTBE_]MV97Nb?UDD\,WJ,_6.XZ84GHS)c>ecG25[YDL
E?D8]\GU74eA4/Y_U8IK+a:]W^=3..,K.+6<Z4bTJ?Y\\);XI8G5V^MTTO_f-?&-
EZ,f4eKHP<O]/=,_LBV+/^.0#PDZ1ZP4CJPaUU2BQ]HN7e;8M&5K5OfN8059^H?G
DH]?a[6IY>9eVG/T6S.AZT?H;U/2(c/T7IP(]fAc=8:Z[K7X.@,TP,3\/N4&0;9c
B]6-0?:)H[>V<[@7\KR-E,<RO?(V>X@^313:=ZJM-L:>NfWZLc_]E\K>cFNZ0\6R
e?L9FfS,2UIbK-Ue.W;#F[aIVSF5(:[_?K2E>aIVW15P-0c45JUFNW4M;\Y+++32
5<ZFc@faF,@)W=E>@0SCFKgAf\JSH<@d<+(MY.H&KXdEL24A\Mb>J:f@e_U4-L1e
6?b^XDdTX\6b_1.W#7fE8GJ,QWG\H?7ED?aX8e>:e9cHBQ&3SPF0N\cJC>;dN,>]
(4Z&[DOFV8d?Z>7Q[Q/VK;C,U30e;;Z=ONOO&[]:,VI3&8bB?U^0:/V4C-.#CPb(
<+4GQ=C^[\1J=d5d\-)3T.VTXH3f5_6eU+)PQ,eE2D21IMZICST91[5/egR9D\;,
<g5?Q+5F=<F2/8d/1F.=0_)<E3I1cK>0JSH/KdVCE6<7ZYM,;Le05FYc7[OG7TMT
@.W]@DZP)E,X_V0U\3P7K7:e?F)0J;/3L]+1B_SfPUR5Q&:B?2QB)JZ&(TEI>GLP
71bQaWMYYT,^=@H_GZ,=QRSA#eZef=^L5D3TKc/+G2;H/KNaLBdY<WF,cIAVEWR3
CQ]IVYNQJde&JDT=F^bS^\\=fE>[Q=_.^H=DT\<Lf5;U85T7S950B]\A<0N4ON](
(CY<HdJ#IM42D)c0a<9:F4:bI&F?+N8+>5L/8aH:Ucf1O=0-4#4a-+#UbH?YH(bF
C8YNUP/VH]9/^/W.S74[M.U0=05R^^(@.<C9:LLAS@KMO:?=8U#S<#I9P]4;LSYZ
bb.PTI6KVALFW99a<1Ib\LdW\J7_MQ<NPXPN?TJ2\-P]g7]FICTM62f=F2gGUD)>
R)c&TgQSAGe]YA6JK)KOOB0=c,d+L1CcYIGTT4.I9,RdUc@L1,5@L0D99<I[73bb
RZO4>=Z9_X1b92++Y(Q;,HC,6Y?E7[+-<cfJK;=O,eNaW48cGfMP@VR9NQM[KMH_
6?,(R>eU>Lf&+RH:b4g1:&,//1;gI2R&a3D:8EM9NNL8M,<]4T]3AM6438\]dfe&
=N_JE?&G.KdE+>D5&Je?3:aK=B3K_C&Z^f3=+e+\P_>E5eL9MGJPM_AFf#T8-^4Q
/L5O9Ce.<)\<]V+=II,<QN@f:V76B^E_4,3V9dC>e++_.NM+>K.C<(0LH70U;9cb
NW]R3L=,6eG?^6NRAV.-;/f4N:A24<(aEgMc+[A&LR;XBC1AX4d1,#2?@cI8&>&G
VWYUKXJNf3#R#LF^/Xe@^U0Tf)\L1[P+AD=Y-2UB^1GY[fGRSLDaD<f5U805C4B-
>7=faLg\3gg(=RF^TGO#92G]3(.dJ3Q.D>:\UM@37+F3XBe6KAVg(Tce8MF?1>Q)
LdD_W?-6+#-c,-<cAU(?=2\F#SE=G.PYe2]D1_F:XI5^2KdP7?]Va:TUH6PG0.1]
c.-<d5WCB=5EXMLT?B31&],RON?HFY#X1bbJC\C[L&4eGVC(:8G0W_fF3D8TY6)T
(ZX_R\U.5];Gb+\Z/@E-Q4aLW;;9/I1;0eTHFYR.b,6,OZe&8e^CMC\IHVM>-\0>
8AP@J:Q-TdFPEC]Z[U@4T0F^gQ5^#Ya5HY4T^1<Ng0A/RTF50?>K^T++5e[9e1+3
/K@K2XO.NE?JR2HGGL@)EGN82]\RP@XB&TSIY+STKL(0>>(3H-(&EBXK,#5^6]<>
8<ZB.#079adE702KHc,_BUegAJIKUf?&E)@[R)OgJME,Z.M^F<&GOcF5O_1+cY[/
6]Y,aeHT&\#eBH46F^R9AN\,BaH)L_AMN9_;V>#6KJ_1H+Fd/,&RMLdCAW2E5UM(
KYbF>/eI)H,O3>Cf,Dfga(IMG#A<HHID3G^7Te?O<NFPTdc[F@96.=6;57b5O[M&
)]:1/4L5b<N^>VM=Hg4XZX>bX76;fT9UUK&DO_VeVOACA-@cM@8,L1ge;gUM4,79
GM4BCI03YO038;Y;9<0[X:Ld=d21OQa,;OD\5BRDYa1?\D@=AAYA9T09HU3KAAP.
C+I9agP53/R#-MLd>=>=<;X#9V>#>3.dJd]\9eU+B=2,@,(ef3.4@2RN.X#1>)H2
^K_Y(35gQ:87@[91^UD1.5Q/HZ4]RU-MW\4MA<IUTa=J4Q1B3b-_WRU>SW1]f=B\
C\e8UUe.JDYcN\Q7I9T@ae;2B-Zb)TFML2BdTRBI.b5&P6\V/&P9ZJA/M>cTUUfM
>#/G57gFZ;/OG_BXg/W0-\1SI<K-L5VUSD=:U[R4XTN7A#7<+E+VP.J^1d5C@[?^
M3TL?,;?8@-e9_S6>KSN#14>B<XbOZ/?_T\OM:/\PY86;dGD?DZ>5>H:R[=,a2@V
:5O]=@a(+cRN<#aMDT#X^QKYXXc127:I#15P=?gXRg2F.f\P0gCP/9<.IP9_Y)_+
7:J067QPBW)SLRKPA+VfbD&aTLVC.LC[W9CQFf2IY=>O6>[D/(V]81G1Rb8ag>,A
J[QLdg1XZPgNB95R.DD#B8:^9/MGTF-K)>eISAAH]Z6RWPP,#>.)=^R@[:^R2=XI
I,aM4eDe;@_S7J]f<Z^^DJc8SH=A?JPGCVK5TKD^XUZ@0YY6a,\\Sc0H7Ce1Q7\8
Y@:Q81bF99_6aaWLOV64.^^=d9EY,JNUKX75W)T3)e)&:Bf7#deb/0UOK#9/M=:X
.1Y1cZNf,9DfVG^?A;TU,?bfU>1P\2C@+e.8c>F@W3>\fF16F-PDKHd<BSPC/^64
db#0cHRN8@BCI<8F-,A21)0@a;HKQfWGa^dgK.6Ba:;1R8&1cL3I35Bg=A,X)7c3
,EW?d1YKIK3<,GON60/)JL7EHOcD[3a[7TQEG>>A7&WKVG7::QGg2<N?4@,-7O8F
:.JJY;+GXCf5&&7Z>1D,Q=REEVK^RHA?\Z?L?30CI)G(PCIb)K=B4PFY=Y<-1N<\
>I02>N&WKOK0?;@dO2Ycc:bNEAWV>S?bA.<aEQ[TQDRPC<C,-FF#=X4>ADBdW4ec
Y(g&e=:0)GWN-NKS(467=3#^=^[C2H(0_U2L:=H?W>.=FP6NX.:A>H[1;2:8Fe5Q
G8cNc3DEA8gI1\[U@Q:LNa0VM)b8Sb<L261c&>KXW^;H=Q)_;R2#NCEE<N6C0I^L
1c925JLW&FGP9c.@(-7\G>/4[5]U\8b;Oef.>HVQZVU>RbUHX>E_R@I8#:YJ;,_L
0LOKg?\#3XL+T_C(#=]266/6M=gZ(Q2cR/>dU7I@YI2V4&;^U(3IBZe349?+JQ.S
ATC9Lf+C3&g,3>0GTGVTf&,:OL#:Za6<6J4UL[_gL)G[gWK\:/H;-AQBb<bO=9.4
&6>#\SQ-@=>0g;BBG]NKbW:H]0T\E:(0E;e<=9D+R<.4:E)1M[X,;6-(U(BH\>gT
C>,C0VdC=MXWL+9LT]=;)U#XA(4CAX->(gE,Y0JA[bPZDKe/ef.=f8d&<LgOIS.I
YVQSa)SY5NBPE4DaS8dUCU75__VPeK?H8KB[N=YV=YN?<eM^00dc?L.+-:Z=:C<8
68YeTVb9)?7-UY9[a?2^?F9Y-5\_:F??J:D(cX>MP+T2B6I5E#D84W1]1]T9_@MQ
+ZUU)2Y02@>C;^da5>MBHWOdQ]J:W7):Z8QDJ,B5@8K2:IgR<25<;YK9\6S[Pf4E
F8U?+D9G]Q7236&3X0J0/,?]U2a[(]d1-X;1CUJ6S_GQ2FQ=M.gM.9LUS^HD]-CE
gE)I#7;K68UEMUL-4RfB?Z]@fXd0P\KdJ>2Cc+8^;AgSFDg#92.Bf16PP>P.R2D6
0^3EGPUV[LU3#;MfHG;XL8/feEK(XeaJ1:D,]C3#N9bfA?JA31E+;:Ug161+N#I<
?/7_40#0.EH(R1W\cU&C#g?_1IGd[LW/YfG:I:^(X+)611WG[<Y--BD4KL>>,?>@
6>?=?BW2Ab4R;VKM\_bD0UC-PE>P_NT+XJ5GD;AZX[^0V[\QGR:RN7_a-gg=TI:8
EN>Le(R_YX\,GGdPbG21g^0U39X.?:(8\GQ/5V8PP(I\0e<g]-+Q-@>Q)N9_>45&
6&[I+\&-2L2#3LR<?#(Q&f4827\CaJ@CcG@aTEd;E@))&;#H?:0(HbZRWO(E57]^
ISM2R:;egZ-c1;-fH@M=8SR4?\dLRN,/0NEGDQBHff2_U)g:;IT]TE#S;?1?AU.I
,KL01D/3c3M:R#H60NV&gFN^J)<aa2X1?KY7bN0d\SR6>0_c^fUJO?,^Z5R=9S0P
F_0b2#^f@1c;.-0L)>UQd_(R0[PT2.O+,,)\7LN(Ee42STef</J(Qf3DZ@XeO;T<
7,M0N\N0U^15Jf&O_A<2BfA31ZSLgBBZJ,L5,D5G<#56;XV@cFb5SI5Q?+;2cU.D
cN:B(?:O#X34?_9BL\WASKR+S.K+bSQPGSNLA4gNR02V0GUF2@Z:8DNCA7V^PZ&I
YVS)?;@N8-X=28YEQ.-PUCgQU_[P.):e)JS3[4?5.<2R_RQ5YANYa<R33Wb9[I)d
:\DBZL0VGHME5BMYfW2,V+g+>a4)DX_e8e9;a[9UAgJEA15OC5b[^8Vd-Q5-/W[:
a,?We6=bBDN@T^7Vc<dPNWL5\Bb[2,P6bD(TWedFK.1gKN3e[?9EX1f1&.C85NE/
&b9X7\0O:Rd9P&KSG&E:Z^cgFLN1OX8<^-_1CJZ)=V0LFc:BP5G6+,PfJE.4#1&c
6T^F=eDNH8[_ZC+:E2P.b\<5?NUaXTHgB[VW[T[;4WZIPIEX<=f2MM?1_2cdEE=A
(F-ZQ;d=YU@J)9&BAA)IQ[Y[QGQ=6QYB6R>Lf.8_aU@(S8-0US;-5R(+@eB.HKU?
?g._=PM0f/HXE=(&(K)Jg</N<H1NHZ,&G<,-[DIR#C>JBCL4;<g7-LU[M^#XXA,H
&)_J1AXZ<UeVFeEX&/#Vb530Le&a6WM,[H@CNXP+903]=9BB-/DWWbU.=g6JbHWW
JKFVdC<W@cJ]dZ;=<5FAO#?K1,NNB(XW5\0AZ9.dSFc_f2#JBENF/dJ?-E[:5<(R
=<V1MR#)g70=S&+0^4Qb:R2Z^fIC:HGRU5G5NNH;2_PIePD^W9>N2KHSNIf[M=b\
OK\YW6SKHQCc\)fEP2V4H<57Y_,8H>P0g5RB<>VZS05[BJP7#7:?H_Z=@c&8Q_RX
_<Q>W\D#M6PV5H:,I)18a3\/UfY:IET+61?KPGAR[(?a<XUA42#90)S4aNI8_BS]
g&[[9OP3+ILPD]Bf5)C&,-;PSRC)O0\.PW_C=Q8:WL.M)W3ZUTUQ);3W7)bO7f_?
f.R/@=?5,]I2#+&cf49UOB9\ILT2=gST@?@+#=J(@3R<I9QgcDA-:02-b2Q_5Xg/
FOX17?I8KP=N+E#;3[AJ=H?YGRH^a,LfU-X_;A/F;ID2/@S^e1[b#Zc:QE[a2B6.
,]c<K-])1?L),(aK,)PIfOR?0FR>/\1CK<D[S4^VW.=R,Y6[>EX6MOZX/VZG.)?2
8+=Q7R/OLKBTB_2Y2TfM.^K0F.;f#I(feS@C.(U+GB?#H<D@_I04\?_?dRFQBS8,
U^)1C@g7BER_K4C-Rb;eZcPRRe\,PFKdVL:B5CfFY1[-E8N;)]HBXLcTZ+9KGDc4
FU[]F[5>^/UA3bgcPNHGf=MCCM01JS5:QL337A:0I8VQO<,_;T@HOg)UFA?NEIS\
Q>O=OaY36S0M6b+6:^_e8X-.3)a5;HKS\^;e^5A3f)K=ROd.]dT:=LSIQUb:A2A3
D-[cD^VDRP\,-9cYZNG(?P=A^^//\I7=,e8dHaH6+?dFMZQV6ef_P).X1JbcLGf9
[ULQLF&+cC<ZU4,Ud?IVQ/Y]Z?8ML=A2<gP[L0@ND&1&1\I8UWY]7:M7#M5d)8A7
>)_DGP:c1AD<T6^8LF\<M<EHR)3FFe2[1K?aC5A5Ye)KGdOa=4ICO?XK=)KAY:G&
>MH/MgF@8M?4C=><./?1JcB4#7+DB9/0<7NgZ,gNg-?M4>@?VKc2)&;@;QD&46_Y
0@&J\@T^M&5:+E-e(ERBKOBf)Fb9N^>KMN:O?:&K,=2\](O,,L2e#UgRW#8LYDG.
U6&_KM?3LGR5N#)([+LB[Lg@R8JV;.34b@c<;C\I.U2;+ZOE[;G?Q3EN_)]6a\(;
.gLFBEK;_\#\1HaHZe^>MbNGA^D:.B=cT,9MON9GUK4a//b_g1&.N0b.&V3H3A(f
GBUgM_Ue7(9aNgUC;fMeV>QL:HTEW)U]g:Y=A:PGH]V6]:;/\>(T,#\c[bR1\Eg:
]4e33.R>gP]EC02gTKW(aaM2<9.,[EC9P,_L?7]aKUG+0\\>Y#4KE>@5Rc9J]:V[
TcAG)GSM#d5IKH_D^-W0a-MSR.BMGZ^I?WaMd6b&?Q:eO12:D0Ya<_SP0_&9\6aL
7ZOBYU16+<<EW?^:8X__^YB)#dR/0.@5O1N<,T#6f[<LBTXAHG,NbCF.Q=AJB3ZQ
E_6DOQ[&e#3L6Qe>g^[eVd8e<#4SK(Y(\bN4bPOc,dBC\RRMaGeH(H=@LYQ_?ZP7
7;X750)<ZNUf]:<SbONf/W/DD7D-?(3Qec^PI(Vc8]C<,FJLf>1dbeT-+eU4^7?J
cIMI4ZQ+8cfQd;UVSa12)/VdM6g=)3c./+-W3@W\2;DgVT(P;=e][^bJ3N/R3G[T
>9^-7^bJ).\C3T/JUN]X+CG52VIa3Me9]X;5S(#RO3g/00CDAId)fX2;,/\JX>3?
CR9d1C@^_>g4965,bQ8S[0Q]>J&Yd5PKfg]3-?+VH8=N[TL7&+2fCTaDg3XRE\EB
E31KNSHI308AEb01+cK87aE\9<4GMRLL24[+[6dGaG5bdW@b((7?6=7dHK]dK^Q=
QYC\g+T9F-VKeUJBO/14:;WQaG6Y;K(NFDU3><9^1CCIbM6W<[QTc/SVAVfbZR5M
bfL#-5XVMM+^^I[Q>,3cHLH8,&SZ<.970\g4CaaN#f-1e,TF,,6.1g[T^3UH;F]M
UYW>&F1gdV4FZJ.1;#FI<)O_cV)-,C^/_b/,FdF?]QP[ZAAETda_I4:9]N9PO7+)
6-O6N@?g;I#U?VDEb\<X\BP-K&\:7]?YdI]WQaRR;])[92XY.@F6\>+d/g2=_[.,
>C;SAI^M<)K_<e4efDS-J.cS0QNY]_eD_@?98F,R;;\ZBT\^cbU:_ICS9TeGR+eb
X_J65_486Y\G3):,[--4SB7Ze#19PK<Y-QOWHI+HZ1#9;>W+Cb.UO03ECJa@WE;D
d2OcJX>4<=Y,ETR_@(8L<OJ=?V,^.?46P5_Sf>HLIR^=G)afCa+=/A1/QW047_&2
U>/F]2SKTecS2CHA@RBZMf&=EcN#>EDFb7B:5=GZR-cD7Te\AS,Gg=^1O>b3(U>\
SH).+);d5dL2>YB(##A>D^.3aI3ED^#EE^_eAA)6W&bXXBB5RKI+R(:.R+>=P6KX
N(7[WC.;JAL69D8/[AAZB0Q0Q(Jf2>J0VB<@adFS&G<ee^?CIW360LWXB(IZ_+Nb
4Ggb2^UAF-^00dGYM^VPS-:FgJ<XVAD&@1d<S\@=&C+a4f.Bg5.5Q23V[\#eW3/)
LB+>PU\g?D+G8HBTWDI]IL^UKJO@fe&ECQ1fK==LMgUY<LgLI0ZFLUF+AfWV;/:_
bV]>Y-_EA]d[2KGM.8W8S,6_POK1E(7/[>@XK4N;F?&KdJA9;RaR0=O5<FK[gW:)
.gJd6)?F(APDCB1b8QT7a<0/A+8<8MOWTOLe+J?+IY_/A6TJ5&Ee>PaM>d(HR5@6
;XY@<ENNG_W1DG+FE\/f?EA2)fP_[ST=e1=<@Y@,&1caWRdAI#&G8,3)BE_RVNGA
TV[:)_N5Kg:^+f_=cQc7bBJJQ3UPV1Q@-_&Qb-4[U]N?,bI(FLH3):SHX8SOg?&>
K.G7B97M8BV1@P3TB/EZORQIDE?3b+Mb06:?1@J4T0\-O/<]-F[XYd<.MY&c+KR?
?:9#@G3<WT\B.OJ97B:S[6A,c)(<F/W:=]UHJdV5#;b.NDc2JTgV>@1^>+K_]::S
X>ZQI=H)SG6BJ@4Q20@433eP;XG=29(_)OYe5)58Lec+f;fZ42;_d_D=9A<T,?.C
A.R->BSE+(1+?D[3(W_@GGEQL[\K-_>^@0P?-(M\JQ:-?[O><FNDVBfd.L\0a.:\
7Y.H&H[SbT-aKL80QZ0+3d5Q;]AK0H@LaJ#@B<EYIfK_D\aYZ<0FR]TKS7)2XK<4
FKD\5E&.[RZ2C+#b7Y5XR9V+KIPD.b-eL:FA?7cH;_g6&?LH,\S#H^fL>(b\SUWT
=6T^d<Pc3TF+9[NP\/9:adMSI67XZPEYRRS;aY=KMW=,,/&TA(&G1N#(:T5cLM?e
QD-&KfLZ6S^Y>g@;:^QVMYQA3PW/7bZ9HJKNMBZA0SVgNUE/VYQ<.PDdFN13C=IM
M#;W&P[DTB&LS(8Kc=1V[<?[gS3H<S9S[d<+>46+4ASaLO2#\>:g=Sg50@Q9UTdQ
-N<X@cLT5SZIP)E,6U\ENgS;.))6a.O4;4;IfQ.P#(e/8;(d;;K>WTQ&[HAEP/1#
(7fd^3=/DP&#ZeF/];([/YPb22f,SU4LLF=MUTT42Y_1-#C7+b+a\ES]-2N7VUN5
Gd=?fc@6cZ:eDIL951]<_D_U3KC5_V;(JGbI:IGKV2LEAgQ1:C&=_)3H6\3+ZXQU
dUd#,3><PZK-Qc1WeF.K<D0#2PU,QL#gWb-H-/PWgXF]eHH0RYE^3B#R_H?/B2d4
1^:PeHGaNQ4C#=?f(0YeY1e8#B[A+Z-c_bDWCZN3:;K6OA2c4+/CT/3c7-14Z_EX
=DMA4CGO#c^Q.VLML>1,bRA;bP1C@Sg^QfC?J/B9X;)7ZT4bdC6ZOI+eOXe-+W>E
Yf[UPG6^aGZ^>8^T0SaIBeXT[I^=geAJdaaJ-N;P(.V,X?;73>O<,#dO>L&<\0O<
<>/;MV_GC2C3e-,HCVF)XJM/R7eF7AZCf-Se;<.AFJNG/6OLQ#M+CEHZf^F>?GFB
);0If1Z&;H+@D7&XQQ5_Z\eD;e/KU5Rd.4<EK;HW[W._D(VK=\GgBcf,:AG(SK2b
JE@DIbd:(H.):WN_d7SCd(?P-J5H318K(Fd:N[_8K4M=a#N_(90A_(=7_?<@.L4B
B:Y<Wg,,^JHIGN#V7a+,BYf48Q&C?.c9Y)CcPCZGP?Q)ZL>.6HQP)]BO(V+D:<90
aF&JY4f?2D./VK+392S29C?U1\G;<S><MNELKNC1XTS=97[D)\CWCTe=D=YAe#KK
T9X\;a>L7QBVI:-]#H@MQM)If.OZb]W:Pc=A7FE,^)/dbb/K@[>b#S8O^N53&99/
/[#(T_a5@BO1&&E#dce1<5Q[OSDY4/G?]I<,g,>-[.R-+C5212VJc+;HU?6fB<T<
EDNF-0XP4D@HW+c,)MCG+U]_7YF5T6dU)VYYG4#F,+E6JbgSb=bK6:@+&A,+/1;.
;C_cc\?^CWUDN,O\\b.fTK+f&R9GYV,c=/UQMUF[ZHSF/HWW?43[3X9YJ.\V[U?T
JYbe:)MQO+KdI9))J(2Q70GZ&cYZAGR@Q4J4EJ_e0RT^XN#M6]NMW/F6;1I/&P0=
aR+]&4OIAe?a_[C:bS@KO=J5APF+5A;5K_dd(NJX@,I)7)1&(4YLLKf-QX6BF)=)
.Z(DcT.W_K3]3T1>K_RLQNF,EUE2-?QS@.42\,EZE60>25,7b1<[e7g1C9Pg?LYb
:I<d:24FN[_PKVYZA#2_7G7TATU&g^UL]0&ddKKgYDgB:XGF)QXA0<5DQ#/5O(S8
)^J#VeV-,9&&6/(dYgZ6>&g6\_f__5LVbV3fQgHg)ADaI,=WKHG+11M<:.e2K?I\
U_.5?bA/)4UeH0IUT8#=XU(Y.3B<F]>DOW,(N>MH1K4ccgYP#T.@:9H=[RV/=IaW
Q20Z.&<(.>/&B7N-,Ff,X:-OSGYe=,+=C>5cHc6Zc:T;D\B3J5EB,^7&1^,YLXdK
dL7RGUY6(aUS/6UR_7bb@L[LR(V9P_CVdbXb^Z>F_AXSHEL^P(.?18/.g3E>YNC[
cD@\[)/M5M;,fZf,Y/dY0dFPQ9f@V3<8_&E5#X[1F>Y?e+Dag325VM2;5a/gUe_H
S.F]+c]P<#G#7TZ.+3S:K6-,/>4cDBDW<4+N=@YS=>KIDKE20]261;dV0]HA6\)-
REUAVg34ID+&=(2cOUZ5bc4b4800BF^9fIM]]B2?11fW^3V<J,f?=Ud_45BJ,OO<
1&,3F:.aP=+KTMU.4BTF=>Z0Z\5SQ\98)U(-YEWXdM6WKQ[O2;U79I##DPH.Nd<2
(0bY\MbR(Q\b18ZPbLP(Qg13:4D^4@[E@MWTfSO)HFfEJ^0CIHL)7-&dU<^bHdOR
:E^JB<f-bF;)bKJIMS14U&4aMG1Ze2NM+/2S>LM<@+b-O4gZRe@:.cO0;8dPPb1T
2[0[()1[BYD54Q=G+PJYN?D/0-.8M#_+\0-EAI1M0_aK/:36L#-)ggfaRX.1QK(4
3AQd&\5VYB)H<Z<FD=K9&G]_B16eL#6\/c8aR#a\VV?NIL^Ba.MFFY.(79I-1#(C
0T<D\TW]H;O?..4&G55.N]OMATKCgYfOR6da(SGOb9H\6OG2c8+\;Y]J5<,]9E04
[)Z8VX)Lc8B&PCDEWDZ7a<HODOdbA7+7HD[e:V34)[.eWaN@V0A(I^9L^W3:F+>?
W67>K=BNP)W\MZdGEM;bSHYE)P3<(9=Bc8]^Ga01KEW-+.ZYUS(S#1[-85K:D\FO
O-/T.3FL_8d0HKP/:B4D;\I2;+-1bG5@(#LOeY7XR+8UC3#=,[dMC?Q9P#1CgLLg
>FX5OcF#D:^2/<66@8JZ@GcAEf.cNDA3VYeVL),Sf]Rea(4Yb4/\03DJI>PMO/1R
[+I(&c.NVP;f>)CbDS<Ec>RQ\TCCG59(/L)#[84)V[3b2C&P5).[cVE2Y_PL<Sgg
0T-6U^OX\8-[93K<E6aK,^U@\4ZO/@9J0=.?:>cL93#?L]<GOMMJ.>Q8X?bC-N=D
Fe8^+f:.bePJ5]+d+972+IL7CWA[#3[^PMA5^&dH[<ERe4T1a)@V.</#?>.\eZ^H
dd-E&,^_fa+Lf&S[,?)deaNZd-Z1dU#16dYfUNF_K8.HR>\bI75N,,JX-2@G]4->
,M4C8240;&a,cAXL-668HBD]OSGU089Zgb_\:;W9G&(<[9/74UD<BEKEHa-U9Ga)
)80)^ELd#+H#Y<>d9X^]MT#:1V&Z;EO7QKNHcACA1?S9_JeT2K.a+4IK&R2=[2V1
N>7VL9J2Z&,7/G\GNcUGTO:1KRBBBcNJET2U+PTAM]U:g1beL+2D<@2YC+T3[EB^
O#4:8L:]XDME.]/5cXgBJC?O>cHW;V/HfF4BdBHLTUPN(?&M5@48-,^NG\U,>>59
@RIU>.JWcSGQH9]RPE.5I1?:M1+6>>^?[K_:,B4(90-FPAG45#8\AK.BD@]XK/;@
P[J5]>S.A;L,c[[QY^ff;L)#6SR?3+0I]f@@DM\^;aK_#9Y>aIL..B9[<ZUIf5N8
-eSAEP\:1T<Ubf]bRQ+G,3,>D17EIfMP1\\Vg<RcX&T+T.(,ebaEPD>,QVSed)&7
:TNd3[cdb]#0^aOKM,GZ->O<5C3^PSLKQ3W11V=OSJ@ZD&fMVgV=Fc9<1W>]J(](
(=<^Ff2DO]BJb:<JI]W1b:W,&)21@J]EW1ID/E4]G)CHIH9[T&@:17DGb9+__/Hd
c@&HD4bSA=5K]8BZX5;W554ce_@GX_4MV+0Hba&=,6D#&I-+R-3#V^1:P50&Q.J-
714fYH1OOM\?.5VIaA=)fW];FG9Wc?d1T[1]W0f1-e&X9V>UC]3(JF;BG#RR3T&I
,_O0eHP,Ce&BeOKXOWZ)d)1Z4AP9)S;4&S1d>7dNI?DO:+\<UMfY5;SRCVg=)I/Y
NL^)P63F82Wda+4_b,=T0;F_W=gY4?]/K>/ST?VEVBTS:)PEEg1>b\I5QRAMHfWg
^].d\4WGPcBLQ26B>G6JD/c8]H1_cFA(JV4fB;cGGS)UNXC<JcgY6K7BgU+VKIU?
A(F</d2[6[/f]X_(:=?d6.c-#YP-BU]IVeK0_./86Q_2T+b5VRZQ[DSDDLQ/C@S@
b7ab7VO:NT;Q9bC2?A8FT\a3;b17XHD:Q9KT=P,JDe\5;06MQ7O#25M<LTL-]#8[
Y\9c??[\0c-HPWQKba7)27UTR>Z/]&KDC[]PIWXSA)ATE[]Wd\VKMS#.;5T2O^]F
WZEWY8c:84d#]PA1AUPKS=VQES(U#>(g=+H;,;-,=N@;@DRW,;6\B6K5H:?LgYgN
GV/E5?>d9XE;Ce@\:T[M^-T0\-[9M,_2URd@1e&Y?;CWJA:6<9H5/]A_QG@F,,cd
FAK0\Ee]5.L+VV9AdC^0D&[G7c18Pd,Ngf8f&78a(J;Se6S3IU?,9C\&^A#-RR&O
?PJSa#LG)22D?<0\_WdJI;cT4N2I[aN2.1Z:JcK]SXaAaA5c2UVHdBg5b=QV85(&
/XC^[,;6L#F9-5-#cc:/#H1/]\U]d>O2Q;cBa)^A3/:M]ccSR2?NeK-J0_(gc@2K
J+27[:F>\ZW5Q9=Kba58b)WGX@N&RaQHOTEI\N6H)W6R;9\\QM;+c#U>Q5GSOaL@
f(>;Z+RX.::(TfZTK2Ef]((X9@.RPMTbd(3,=DT2RO<W@NCKPW0\R>HV:Ib=.b/S
9Nd-)G,<YebB/6(FaNHHGfEN^?Bg\3++c?@,OU?;E]=4,e,NR>^KPBLLOYc_ULZ:
G=&W_MO+.CZEGES0W;1XaG9V]0T3Me0L3Wf(Ka53][8_\\gA73MI.9,T-WZ.;28,
AKaEbP-G^:(A(4_&@/C[.Ob61:MOC,GB5Jb77#KX66PS<V]91QF5E((0EE1XbUVQ
_:(a\fTN;CJ\U/T./g/B&REP+g:J\=#_ee[^L>?gf;?[eLag;.b<TIF94Y6ZR^g#
9S&eWD:^OW@0Xa,&3@Y.VLZIZP<Vae1?N^0R6B-L0#Ig^eF0ff8AN+LcZ_#RGE?>
8V))d\LNVeWYAY6E=Vb23DIK.Q4([8a?aWcE<[6OB;50:SDX=>M3;FC=[#LFTGQM
(AH-2^/e3E8M8BQI(YO3Fe1aPNbL&cKFEE4_BYe_=KZf7(=.Y<H+.;()a41P>Ga5
bCM6<PXV,bV=[_=/KV._4=3+6d?KJ2]?D#1M:U/b)H:]?Tc.U-Z;7<YFG-0G48@0
(c(NY0PVcUXZ5/30WIM@(\4c^O@SgYY14EL#EGEWG+:-KdF8CeKP36[6af^<?R])
[]Rd#:5:@B,383B/W4C7CdZg:J47Refd2A(::C0H#Z6/\d6Q1?8W5:5OE(9T)H_.
MSC+>\<:,B2BG7-PVV(O7.CRNQ2PIJ@6Z7T>.+-U:1DVQ;W^a,52c4@=5TcHIM^E
c6AXXM-7PWHWQa^AEZ6?PIM_DVF4-O^(GHL>Ta4\]UKWJZJ=fTU-:Y3,):Y7,gCd
H2&YL?Te>E:U/XP#:7&ODe@0[V+UCF,+)1.C0UQdYO]LCRYVcgX4Ie[XaTeJgG@D
M6OQ=RX3JN9W@5g3aO]e1W,,cDTY(]7Y@1K[?^QN=SYS9W:)P[[6O-&YW,S4+8DH
HUO:0gA:6QgfM.)D>fed&:1GQ3IP7]Y)>R9C4TS>)NCe5GfIWYN.1d]Q[.V^/L\;
PQ92^F;,EMLHD)#TY@4C]FUO0YC]CaEQ5-=1GOE9E484_35TH\9Me_GGPHf=[VU3
(9#dBSf_G4XU]J/]@e9ZBK?-=QY_,F7^IfL:d/YM8Y1>Z6P1U2RaE^[5Z\QGM@II
8e0MYd\BB4Z80-_e1P2SPR;.Y-L6M#,^LEEXbD_O+?^DSE?S#H\GJcCf1&PKR]DU
G^5WP/_(_4;C290X4=D,?_dZ4--&JE^R1(P1P^AV+W-4HC7=V>4/D=@b8,Yd(S6^
7bUY0P6>V)1_:H2/A6EMREU-G:A^LR&dg;@PAQ380H(1,HWDcb&b1&UNHT#Z<C)M
P8,eBE[8)_-^W=(\<^CG;U#0McVL_@)H,@17/VLc4/DOO&^6G<Qe4+-#fMJA6\-B
XGHD:IK.\+.^ggW-ZbN,Ba.KLVXK#N4_VT]_IP0A810,>(#ZN?K01BVTbJE)&\S+
MO2]G:bccE;^Qe.f9OB?OS:RO#<)XgBM;A#1QI;VN^\^3N)-HbZ57Nd[/L&HH\#V
1EKN/_N&:);#9/3=79-MC\ZR57=^\6(e/9&?=I[7FGBfb/5K\TE+F-]MJ)NLGeKH
?eQI0N^J5EO(+Z9W>0HNL7(.+YAFd<D7f8OHCLM-++f6J8&@JS:FAN\UEHX8-Y/U
]]O]2WaY.J-T>f=8dU5Eg1[[&]#Ac53]W9O>&7>Z_7P:GYBdUH-Kg>O7)fIG(ZQW
TU2YMN9Q(>VgKb7eJQ>F0/e^>ZeURU4(SD7d)EWUc@DcaR;.OAZ<H/:E7&[TgCU9
_UI1<>FXJ6Tc=6#CKR<Q<Y-,7D4RZ5bROG#)=CH#Ec@.<WFe+Q/Pe8IHD3&3B]&K
)73;0.fbUC)@d8AYe7Y0<)T2?b75M,=bT-MABHXIBH/XHUPW3Z?c\#I9T?LS,dW-
cNKW[<DcAZ7^LeJ7N5?\1.eAG0E;YfP3UTY.^cGO<E/5WHdJ7DJ48L@g:HGbf/U_
)L\Lb?Z@GI,PS;KA=M6<Ta0^8(3(AdQ8c^5<\Fd>I/ZD?RBdb.Q4U>+4&VT3O6@e
5IY4fD,JUB>Jc14?XLTLL8^H450\:L(N-8MM8[2/;Fcf(2;8=_cc@[^O6VDY?<VH
[0]NO>9eK;A=>FRV:J)MRWSI57gbIBIPA+-R;]4BQTBg7N?2A:b>eKBM)M-f?;[K
<H(O32_RUO-8ZPS:Q1.\&><&_C8D\@_6ZJLZK#&H+G1ggX^c^?aM#PCHK>34CF3W
R<UZ3,.I=FBDDDNKF84\g&0&??>5L:JAd]gZ<(S/TH+V-g0.@55LK]DNS(Kf[T0(
(9[3eGRU&I+Z@bHF2>(JKK),#aZ;FQ&<YRA49V8;U;RX66C.R[2[#0+WZ4(gKdf@
1bHWJ]Yf+#Z6BD#=]F_.C<&_aJ&7+/(4b1WJ5+XUWO<G?geMA0+f),<>\?@=ZLY#
@5&e=UC,Ffg4Eg.eb@bA+J3WH)QH>bKBdcVSLgbHc/M;2:+aU=@3;_8#fT^Q)V:.
GHaaY=OSdE#A\>7(:dO_8cJ(4Y9#\Ld?[NEYNGZ@c:VbQccgLMCAY7Waga7X_G((
H)8HDOY5(<\RFf4E=6U>JRX#dd\#S@;^CPF#(2M4&&EA9W5/)?#THQYJ.XFaB01@
^FL.VOU=@6.=(S^LRcE_c2QWY]0f/5_.QcFEBI/cEQZJKT/45Z9QGOfg.;66@2<L
4\::&-#^6gN@.0D/\R,4>W3OH8#3W32?9+gW.7CM](A7f7YV&&c(L3A3T#@]GU0e
.[6G/12MR:AcL2??.Zf<.XTAH:B-CT)GCQc\2T33e#2e9e;Sa<U8d6f(dEH)c@[M
RNFdJQG.6T?^HHD_N_C@V/L[(=eUDb1;15_Z_D,2\0QbF8^-CKgC5#^^O(V\4^_a
TMTLC#>2INM_I:+T1#95)T1:12>9_T8YZ<J+NEXK:Q]N15e=D5_-SF(N4CaX.N-b
WA)B0&fbLVNF]DCNE1HP;#fQEUOe#8X5:G=;Sb]?U596,eg854N\RcRK@SHbP_0>
G8@HM@+_),<P<&LT[9<+G(IJ)B&TR7:?XVO4L23LS.QXa-,M\G1T1g\-(b]>G3+^
Q\8-(>HQPTO>?)Oa3?FH&UJ4LRE@/HSL4)aMNA)&1Fdf_(DO^J(&]:P^/fTPa3NE
)=0FDL72;g+T=DG],-YJ,KB/7/@OC9SJb?1E(/;+7(QAP465eeR2<>XNd?.G\C@Z
Yg<V0H80T=HT]ZB]:6R;J/.#@2fdRV;=[[a=eEZ0NLZL7d+7&2dD-;NSUH@bCJVe
ZM/=^6A#d;N(C(#98b?/PNc[7dE68H>fYA7O=67>3CNE=&6-,K(B^<^S=bRW4E5C
4+6N2B(HU70@+7Ia[bC?IA4^@I&49M7><3K/_;FA7G5bCS8J3W@[LL80TW&&+H1F
ZXfKTAUQ5;Pg(A5.ddTOIZ8_c[R8;<2?VS27.=FcdDce[1GcJQ;\&@1[4=\>N\gM
f4D59YY^E+X>_b<6K=e/_TdF)OWQ<2_f#8AfMWWA7@E</#B_aY]7L>,gaN=(@E<>
c(H;?6?K6RCVVR=cAd[CKg:]=N/J/FRJ6YA?FVX?2P-fLOSPG>UN;1H7/2?1Ubad
BCHX9M(SMFUc3+_C=#FT&^aAYI<1?+?;g49+=&EI>AO6O&4V0A1=b]U9&\]Wfd,Z
f0]/99_M#3D]W4AN3_C>29HGYSga0^DaH&[KA\,F=HKcS(B)_UV0UN5B.;^baP67
>C5FS5.]NI2<Y][I9(\SM<:GRMM7<]<ABUYV963Ae]=]db<_g/C(7@W4De^MPD6V
:V)gcYW1&Z_1T2Z::?8eGeL_/?D>.a/F2f2>3H8L[/Z,bV?a@U<TLZ9?L,@IGX:H
:U.^f(26LPO6TdY;D)_f&NISJ7/>U>I<#>M+8dN7E/WQWf+#UT?2:)9]bC2M>3R2
,IR33.\B^9[[c^HM4(NULE3f#V7>:E]1:GL4g_U1B]77FQ_PUH6LX4_dA2WC.^#?
V4KLC=:3ZT&QJb4dXRN=528FZ?KZ968dNg8<APG?-6d(9TCX?eQ09?-,1G&Id8Q&
QXC\-7S@\:=aHR,F#-@fU6ZYEQ1M()PM;4a0aV9N5_;VYE[c6_LU]R_EDIBRNYTX
ebTQ,888XSQ.UW0>fE#6MK28UcXfLF8RN_-e2+V.,=7#^UIJC]IP+QF+\7cfAB39
5bVT4LY^+]JaB&9BT(YI).AVXE7?,V?V@O+46UdLQ>QN&/?R67A@Ba.Y-^G12dc1
@K;MA;95eJEMZK(Q.\^R096/46@;GPNFNab2D&-LFN.LF\N8aNYe2_0>H^/P3^6Y
7.U(;]UdVL1F4B0JU?#_ZC79dXFWIG()4_CH6I;J@+6AF0;>1EJTB?5\V>[#DS:_
6+\G,/Y+0-_@fKe)PJVH1E_,L+1.?d2.f_[X::&C#1Hc/=J))VA.2gA8=1a]K3Qb
QF#a_?=[39G8/XbHfMg3cQN_eJReD3G(J)Xf#.;Y\?=+S<WH?E3[#[]<CdfNWYV?
:R#4&<:)R7HU)0LOSg0AZ25aBNTgb>Q.F0IN82QCRePg&@J:<^C4Ffd7Sc<4SMEA
gX]YAW-MO+e.+Db@61TO#g\G/79L;Z<C:YRWW(/2QcXb,+KM6>:L:&LX6+2.\5dc
9HBQ,Q.4K=g0^cK.XcC-4\&KJ0MN=SNOZ9S[H?Q0L7Ggd5e&?T##B3.XXBRb<F)O
OA:JB0\\f<0Db2A;1TQ8IM4bEK@cK=;a4VS7EWeJMVL9K>O),>=CG7G<HRG[f/AX
<1c(2Wa5L1]SO]Ud/OWM/8(QT02_?[Id<&=IBHW^dP2>Q(7?VeG9PP6c]3/L&bND
@_]XO;Q&F.+@6TL>f1O_Ic^L7P]S3<[OY4=]0:d7^,=O4dJ6F&_5:XZe^(_4aa<#
V[?7@)C0_EZ\1JHNf-T\6dADYc=-?6FU(\815^a@3<=0\>IfFaf0BT#S/,:+BKKG
N<&9gVce/AJ6K0F6M:.a7J46=AI,feG1;;9BXYV2KI<>-fH^EF\cCTFI(a/O7d?@
]LHfBQc]U_Oa#eSbOF_[gZc=#IAC#<#&-fM+>UG8)1C/_.#2TZd\?L2B73RE\DN^
>M>\3a#?>C/cA-:A8a5Z\]BO+.eNKL/LZdH3f/__]?C2,_6>:E:eKI8REP#T/cQ@
XJ,VI#PXaA=J3&D:4VQJZPYLfg>bMO<H^_N@SV?3T29+FJI5X(M035Pb2MC-E9YS
WD=J5F9:?2&/eeLHC983X+Q@A/b>^-Z#+<F0/U4N5?RK)Lg&MJDKICC42BI6b6XZ
T?Q#\0)f_eU@4PdE?J6^\8<LQ:SMYO1IAA4:R@GW4U.R7H.??-/ZI544)OJSPQIU
A]4+&LA8>TCYOfC)B7=&GXa_a<ZcSV?d2L+;2EW3=/^Y0^L/f<9eJDK.dF6c\Nac
dKg2HKBIKRE9=f;KCUU#++/&c29L:/A[FR:gOIV6]H&K=K8297dHKa7OYD6EZ/I[
9.a>F<3Vb?U7dDB@<.?626O#0C2-5E4Y-22LFK)Q]]d\TM_J56SQK3T1G[(7SaCP
CYFe(>KLJ@3X7E&M3(X[R_D,86<b4U:(LZL8??.Q^HS,B2&9^.Y1]&a>S:H-McX(
+3I4</QfX]gU),M@MWV4ae=I;>+;f<JHI2WH0Q311TcE9gI8LVaC?daNMYG<)Ud7
H9DF.R<EPcQ29_)/5=F>:QRUWAPbTW1[#><[(99^K9-[[V];M8ZEHX?KJ?634P)A
R56N00PR(_aS@QRI7b6.NU(Y0W(dLY6,GW)gHe/G[W<U#<b4f\]HWg;]&KGQQFXS
DQ?P?C4e;&#\1<1Gb/>[YIQ:YDN>^\I0[<Je#VN,\gA>B\[YRbQ0OCBJ8[CMBG80
;H2P6T1SP?b(&)HC?709=P6NQ]-XP7R[;UDORFMd#U_I]b5H0,^]<X=Z2HMb\(<,
FbND7>?TO/CO,)5B0T>,ee;OQ0461eQDTV<;[8#L&YdZ1gXe@/HMCgS+Q@LV6Q_^
QBF5gX3AQKJIJBaaG(:Ge/.Qf86,\DS??)HK?c&LA>8S-1_//^5>IeE_BT:^UJ.\
GUWRcOg[DQ,2CV+D.7F#XF@g?a9X[<TOKI9=\&^P87-8(K;IRgGf,N.S_I8A458.
M83=#FBd7ZOA]^:e;XW[a=\g2W-IPPf:]3,V?34?^B^5=gZ5VPVDZ)V0X=+;c#+g
18MIa2@R8J0NGC6,/Nb\LeA1/XZ^S-YW/:<[M&VORSM3#>3;AM4+YB]#ecZ]#7+d
0+3Z8)X7@A.QKZg?:-<eEaR4;196FD?Ugd_g,N;]#20]LKMX2/Z?J\](gTQ<?\8V
WS.FfW9aNP))cd5=AM#_(2:<FPc^]WG6A#KCceEVYP]:1.d9bA\1QAVP&9[8]]eK
6C1R+4EVA&?/^=-D9(eH?f?d]K^S2]JYV-:.b^7O?Sd^5:.@UZS[8f0VUZ4GF+++
RB])bgg(^B<UE-^Na99-88:a,O-M+52F;;5affMG71AIG(S1T?a/=AN_#LV[I,\)
OSR9A(@+9(G+0SN-gXK.XG6:cVc[SN_^?AGa)Kg<faT0P:)/J@fM-/7@VOT?5f?,
@dOWg8,]/G.DfVPg2MBV)D)L]bAa0\7f5HYC7;92].P;@F>=,A7a\F3#]MR^&O^,
;T8/OT#+5I]Wb9\]B;#]VFY.33\Eab6RUMbX\I,cbKMFM,0W2)75eg1c;T6Ff[CR
5DNeCPQA[?TZR[eQg_LC<=I0b,6KM6ef(QU__6Z,ABI-</AT9+@&Ja?;cO[Ie&L8
VAK]X;TW3^AVO@dME@/=\G\gS[:H/S3FA7^^].8H>WH<_GBLeCG-U=@[,A8UM81H
HEH?>4V[5c65(:213T_GJ:e<.::K^N79Z6-b?UU7.8]0bT3R@\G+U85;\8Q?VPcO
(X63_L^5A@DQ&@/AL8d)/g5FJbGHF9A-Q\g?ETacY#1.?51JZ[_R.PK1QCC,H?;&
B<DObPKWZ#2<V0D9(]2afQ#Be9?+T+UX9cIgR<@B#8dW2Sf&.gO5f7EE:Y;2_2Z^
?2Gg;30L[P&c8Z;]BdO=<U^141c<]/7FP>+ZgOcM9LHSU^_-@a1=PB)K?S7d+A<G
G.KI6;6fIH:8E2e&bgDF+.RE&)U>F[K-XP@[G/D5[X<0J;JUXX:0R2F+1X&>JS.B
D(I.&\W2/M_MCa@.HE=\fM&-O6MI-.ESI#CbNeDN=FK/_8c:gX)@4+4?,NOI6_-:
A_MA54:C^a\=/[[RN;:1d,]M?&)./^LPg^CY.BY-OJ14?OV^J/=cX/6X9VSb&]f^
,_VNEA_.cP#?+dQ]0;2VCJD0(\H?fY6[4<;>FI_QLJ0Q?@PIU#4W^<SJbZX?Q4aM
+IbG:P5<A)e2></W&DHSbV-I9.C87eUbSReIG-f.f<K.^e.SXHFgDYH+aFM=4R7:
6)(4,EN:dU)T:]<2E,+H2\T_;;F#9+@WO=794YRXP(aU1Z[QH.ZJ]LK/.KC-;Q;6
N_Fa]+8\IA7N<2-Q3gI,1N)\Qf=(GP@^.a763N_.?T02HdHc1A1C=VGPMbP@Y(TM
W>MRgX/[JG[,gE^3If/U-.2c&G5R7V0&(,2>ZC9A+XE66SJSHEV/3^gA._A;^023
-ERFeD/Z7??T;CJAO@:FL#61#XP^)Bb3L1OLNYEbXS,L4/&?A@J3?U4=)BBP:/2G
4c,[;QH>NIGEf@M.L(16/+KMK9Z0YgYg:G5Abg[^Wfb?M9@BJ(O[,ON=L2[Vg6cY
H&A=eH#XG#Z,a^(X#0g(IF#(L[;VGAU(T,V[QKgeT54TJMYUNOI4+?7KBB5+[=#9
c)&:a/AG:Y\K[IX\^_QY9>eO_L?(?BL,^9#3=>#LN3b\]&M<UVT,L80+f^BGaDSV
F_F:bMD(.L1CTC09X],b_@RY0=+_X1AKAb(]Ee,O&\AID6^&aXCZY;I>AR=F71=O
(^>.d[-GNf5LB+_<6K:7Q@6dc:bd?5YaZEXTa)&8,E[54c1G_94<.\D:Y;)326GR
+6ePV\FGWf=ePR:5+0.@f)VD=Ue:0XHW<YNG?Q(2aF^UaLC<0Q8KQQQ<)De0eB93
P+)<+_/96SI\3V]FcQ<fG#Q:eR>2W8:&VZSP4bS1-/_C?Ka+4P<2?D;GebTV4c&M
1:TM]bZ7Se]b?\?\KA4WfQUCE)_=?S\[+UU4=d]::;&/Fc2_;9WGG4TacT8,NNfU
@Bd^OPWU]=W.,\N:33@?Qa[2c;eWTa/6G3#9T+SWP8AU3_\HKZ7Y)T4MeUT6A,,+
S\U7=bg0FEb86:Hg+2Z)N#1&aVA1/UWE&\,bLF)Q(EDR]&AE\[\997RVWM(<J[AW
Gg7)ALb#.PeHb,YHKc+SdNbRDF<SB2H5I>IRE9QUZT_+OTFD4J7=e0bDGK2XO6dG
fV(-7fdGb?CE[&g@_5GEZ)>A8e<>>;M2J/WQ#@?cTQCN)AOK6:;KY3f^#TAC[U8D
9#g+efF)&RaO^a&DS6,fU3?bD]ZC9ANg=D=\=[-(A=4EYI6,)[dg9Id_XVRQ38Ac
/]e\GS?,C-?4b;_JbEXc3.<MFfGaM[8)>-^;5#[@(GLd(D_<\[Z^6NB^];IAK/?g
&I0.1M.a8F4YLGH@1@W>bH0AT7&bbMd2S?)>Ne(C5\G&GV4#Q\MT-<(8X>^NINA8
SBVHH+G<Y[Z?V6Xb&R5+.2N\M)EC^4,QASTTDgb::PAEPfSOcKQ(EJW>e(ZGHDIP
f(bFLN6IcEG)3Y9ade9e^S9Ic,J;CaC;eO3?C>DJf5VCVKeeTgA[PM,:X0P+F.,(
FHH><.LL_H7(IKYaGHOT):45DRVP5HA<P2W=R)4T8ESY6^C<BA>dC(Q_QG?A(S_4
55b4\K7XbJ.<^-=3D>A9B]JT#>g/6SP/E2=&(L0[#b;X;>N-=VB28C&:+>\>59A1
Mab/Z8c5[d;DZ_>d7_HcePLCUFNW(RPXEJ1-7+?G7F-?g]D5:J1VH+,@^;9)=E0G
=AGd]^=D^K=4K0V1e(B\aKWWY_>ACb6V\,U/TJ)&]AXa[NJS1-X[T4[0W2GG6.b?
ARB(4LLB\[38;G@a)-669P;gUONb^CDKGHH@^.;?Z:?eV,U7Q?>aedJ+N\4EgX&#
RZ+\CCdfM:1R64>U(6>=ZLJH757+DZCOe+F+Y&=_</EM2@Q8T6U.c_QS<,U,,<V3
+5KX)[S&N?BVWSCUPPCL75Z83P#H(g&R\/(8>bF8FNQY?EV:;?YRDD57O<f@CS/g
+YP):8-N-Q5&aY5a&VaZJPbB<VFJQ3;0I<0DR.G2GdK5?7Zd(Q&gDPI^f.^^\#IP
X3&T2JgCbAad<e76;S=M)4(#H@R,[&^,P\9gT,?1T-&WL:.>+Ud,d/MN,I#/S35G
MWEA)9Y5dVWaXJ__QKYHDM30FZ&,IPPgbVV-<R4fQ28CA+YVC[Z1M6OH7R^^L=)F
V9A(/63GCNd_YcIaDQ)I=aF3+:0.TfKV-9N.=Rf9F:bOW>S,S?:2JW)DGRYX1A]K
f9E[@#\H,HEZa?,]6R-H/XfVNeO)6Q1gbAEO.OYN70fT8FEX5P_>UG7@<,b/27bP
O^[9ecTaPG5_?J,(RH-HHe#DWJ0R,aU)Naf,&I_XD7d0AY].]bCG@f..ZF@\I0ND
_PZJ)/LJgc7F8c[FER+-@5.3?-JTLGOY\@:b_5X>+[FF\GP;KCRbZ+Z7@c5c-U0R
ZKK?Iec/SVFY^;CTMQ+5dC]CZfM7FVN=?4)4Va_3SQ[-7S?EG[A49BQL8YEL()+O
bEA&Z#;[)=B0M0DN,PS^;IQ42A3fCFD&ZMRW/5JBIA#66U?0Ra-^S=c:0c#E3ET=
G3ASCO2,@24@d)[f)>fc13H2F9>Q#DBYV9g+.I8.3-OK:bN0HAJZXE>I5&:OR[=9
d5-GbEWZ45?DROSV4Z8eOCFJQbL]994be3/(HY;P-K6]YcDXU/BBAC3Cg?fQ#2?&
T/cf9-AS(Y8XF0=G-T#8IaWNc)R;c0A2WRNg+:ZX,VF+@<XB]WK+GELFY,28DDFD
VGd6&OHg\b_5O>-.g.-8].R/>I2Y,.]Aa<a3_,cD<^\N7LS\#9H2NaA;^8/U6X=A
_Y>)B-@3baNJe?-gJ=V]KEHeCIeXZ.c0fec[a]D0?W)eA13g(D/:,&@X;]A)JaNJ
;-1b\@5RHS\J,<)D0f?&->5DROJ:I8S0V)dVe&VDN3^UgW+BH\#FNB@>M,#OcVIU
d>IGNd8V,aD?2N+eJU68#\ZE(<BK)fMb<1W+gG\[_>f)d[)3=&_M._.,44_3d6,,
=eQ]##+YA^EB3PXBZ0Rf<7DP:/7[V1fP/fTc6>U<B9XPgM/RA-3H0W/NH#:NZ(Q)
eB[,.f7OW5QT;<36:PI0TB8.9F)d,)B=S@^IBM_J#.C_J)dIM\T]MFH&PecO6edX
69--Nd5+SY(RfX^75f:+3)/N]c5Dd]AHECgE.AH\&B5S4:-8;_IM3aa@YOQ=(#7/
_^[T#GeXX]4QKH_Q\P0PY3bN0P87[,G&(HMb?U8+V-LHga(KR)U)FY6V+Qg&VMcY
X4NTHAgSIQ^<9C90BUC1UNAeZQZ/HP&;=N9ad4>,=IY0\78[-@WJL<)M=9K3UU^M
4>E<KU>UJEcU8V,M5^CbNe@+\.c\Z;D+8I;-FbId)dZU9e=[]I#(FXE>@&LKO5.G
LIV5:3I&.5Yda<#=9PM&0P416=]=5#gcD2Q0[cH@@S<@YX-5^159M^,W(b_1TY48
?]8?WM2M#C3T/;6?(\G1c6]#(OS9V-VP(0M#M#1G#P<eT9cQX^K;O3R&#&?[d>a4
IN&SM&.CW]Q+=;\OD)1:WC\6OGFYEM2].N8R@9c\1#<73AN=10V&NfFHVK0KC3Pc
_]S^9SH=@2ZP]<.3+,f0142<Q8=#Y.HGYBMO<3[MI,\^)eW7]c4D/&D94R>>\DT3
:3T_)F<]H\]U:3&153LXcGX#)J\,;S7EOWHa;PV;AWIRaR:JaI]fgeJ+/101:[:1
GfO=6P>0,\O:TNYE5I0)RK8AaE2F23OHb&G_501UXM6QV8Q,=[@.Bf8K:]K=GaF,
TQ;][J^J&F@)L&URBH?Ra.UG85-#(/fIbF76FIa+^VBMNg/W)5e6X#MI1aH+fgSa
PJM<U[J+<0+Y(Jfg@P>5D_:\S>.61CQ<[N3@_IUMO_(aWbHZ67bG@&f[56),CCaO
ZX5c^UKP/=IT3W70=3cQ7<+7edP3&[4047U&0c@P&@T7aBFVK0a=\6C<_&eIN=Y\
MdbOD1X^/U/Wc>f+B<MdLJ[Ba)a)(Y>dUW_+,?F5_]_NL+6FP8G#7H<&F_(@1&^/
\1\.J[60HQ3^\T56XfKTbPA(=b5@G/.[d/AV#+V.7aUSU#8JG8WJEVeSX2eLPNZf
,.+9C6UeQ<b2LSE-+_8W,XMJNd:OXc@EM)eV6O7#OADV4&^3C3(=VcG);3(Y:KR9
&P?QKM?HRGZ@+a:QB^?>JFZ5LeL]X@BegBfc]M,8TCR3g()(F^=(1I:_KD\aN:?a
Y=\Z&1+X:W_Ke61\<8C2c>Sc@\BCDG>@#b[R]O&Lg1@C5L5:(@Ab.[Ie5)-HHBB#
d&:Yg\=1d^.DJE_-5<Lg,M4c=e,F4//UfIT(XG\>OWT5WMbOWfPFL4)G;NY<7CbR
cHTDe5.U:EdS+?V7I;Tc[URad..UD@f\-?E8H@W/<WGKNXfYB)9Y)I,6J/e61NFC
@)Xg#NH?#<<8ZX-d;/PSROCa]&_f&SHR2a>V\Tb<391F6&-];88&K>LR4>+[O465
\U_,-fR@?AZCg=8A5C40E9;^FBeLgXE@LOLVOTa-HZ;6SZ@G5B,H)TE=NG6,EKfH
VCY+@I6>@b<1,&:7O>78+X@6Da+=Y-Q&?PJYW>7\XG3PURdeH=7Pf;MRH[a37<8+
WW8e1G5WRge-a#e\<73b^gV^WE>X01Ff]O_,)/9:LdNAXX2_(?@L;+6?Ee^M]g#H
IFR_6W0>=cN6QZe_LF)0=E[UO/Y4D(3KI&Eg-:KGU7Se+E1=(W@F6ZcE#dQD2f#>
5X=R^BEc(ZPZ<.01^+47K[S@<2=B)UG7NY2=Ea#-HbKDJd>;(cJ/b<g#R@e:_M0]
3HFUAf=+:2F@5L^0>8_9B_7C90]3U=J&D>(+=;A@(E.62Cg.S[1,ZF6N9If<FQ.:
c)==DM;MRM7;I&\@DW;W9.&WTa.?<7+BB/Xe\R/7802KV2>014bEcTP\Y7(2DZ+S
D[JQ50KMgcRdM>;)7:A)T.M/<Q^IJOb)^Gd9VSEFD8,e,#<,7]2DR2/?4)37+I.E
1-J>BBA:&5H.8@[QS4e.-=b,PH(U:I-02:X^UWdJ?aZbVgU&.QZN>0E.Xf>/93==
L;@NIV9AMKU@EZYg,DE6^GTWCZUfZ9B03_-T=&R8?GT3Web;TgZA;.6(V.?Q7Q^\
-?fa\9X8cfd=U5&-1=(-XYCBgPFc8eP>/E7IBY1cZ4_Y]A/8fg3[)Z_M()8_IWag
R.W7bKdfd5S@;F#G75T@Z9dA(\WbQ,HC=d_b4EN<Nc,HY6dD29PJ<HT1EaK>aN_Q
,]TH\4Y<>C=^@#VK+ba_NI46M625a<I:VORHdUL-&GWG52XE;2<Y=ZCK9;,Z8&(7
\;=GR?f:1#cZE^8QII\N_e+P2c+J#ga[=P,Z>?1E&]ec@MdNc_GPcWPe+Y.5C#46
1JR=eZ=H32T/#Je5W9B\HFY,J]YbSeIf(I4b(Z_d&9E51_M)3J\FcF/2O=)&@W0_
Ia.#2O^QN(DfdJ3W-)XE-J#G\/3L,6BA@E6Za#<H3R6NV2f_V4_\fAg@aKeKY+Tf
bMI1T[8:eUfG?J1R+Y5a]_0c_@d:S54Je4YS;d0afDQDL1=e56b1S_E_@;>HI8<R
VT_+F9QE?XK=<HJ:R4))_P/LW^A/N[_&=:\X,6FO#9)2/M=\8^FCW/GXOa8.d1\J
SJQ.RBaQ^_]KP5Q090c48>VCbF>6N@Wb97@5<EDeZM/5O,)S@A3^=-L9aN8ULb(\
@WFbd/E^<da(Y9c6J.I@:._dI8@2NdFOK:Wf5>OA<b?A]\>U[KYV@N\/=a6#_Y;[
a=T9@]W<)d^5<FB-.[Te/JO#^/(=J]2^#TeC\fA&^<dO#?E1.>Zd46UefC30T9eb
S3:OX?D.PZ[,>8ZJdVYDB2eR^cR.F_Z;^RHEROY:0(f5<VH>Dd7<>I^E/8[/6>E+
I9IKDOG>>5[NFA2=KDXZ?/QR8LSXAA3g>72F?HSaME6JR;?fEI3T+RbV(ZK85:9.
,-\#f)OD)NX)_.&>e5=HH:7^@C(((T=a[_^dF^.CfY^L(JCc/:WT,B\GK:@W\-7\
N&(CIR9V^\YHfF0328B=[P4[P\HGa-)(gXa\T^(P[\.=(J3LHM+AL,)P\DV1aBMU
#KVWV##,PJ70ZW7YU;B?0V0OLYaU,13HC@#K<\V?V<fDW2a;J94fc41UIVF:4e^P
2W4])G3NfO@Q[aSFR+BbS+e\RM8J,U@8Db.U&;d<E(Z>BWRICVC=XDW)R]110V?6
RYYa49SI@d^90B1e,d@+SVb7I0D_=M(OHcBPfZ>>E.0&^,KBC/4ZVN7^5BCD0W\6
ICBIU&9A]6#ecHTeM75;#/FNCcaPc1/[9^BNY_^N->CSP&c6(dQ_D]37;XM+eE37
[9dXR_SQ]c9P43O\X#N>eW+R>IKS?9#G#H8QK7K\DUVB-EGQ207-6I]>24HgQaI]
W5WGW<;#O/GG5U1fXZ-Q/IOe]Z?L5AAR]]X5^MQECGCBb28OE@AJ??G>GRfATc^1
V^S?[<?.U)M>4Ze0FcC21R3-P9#WD3L,QTIS1&&0?)6E)g0,aI.=0)#BK4.:T^1M
@8V#b@)OPF(R1bH\+S_[2BGDUY@&OA]^.+KbAfaIF.1X2PH[^L7;@GGIE#WV&_QM
Le(F>1#5R:8XF#H9)-\<:#0M@.BD3V,FHIB7=fe?Yb>4?<J,4TdTe9^d&BI&IRPX
1N>\eD?4+U,dJL:d5R,<D/K,@[EfQLSZb>M2TWPAY--K0;AM>QKcLSE)].YbS)M@
NGF7J.7)O/-Lf5S8,6^K+V]99Q_JV_91O9]3).V?FPX6A8EJ\-fGY^)5<E^.E],O
]bA[.P.1NHEAa.a3b8R.M0-a;_F1J7dd<aD^L0^gM@&9@>dM]]]-TP^5b]]Y22P9
C?Y9F87P>F;S<E8^_+M@L9\BMNcVI4#+W-aTED6XEM;M,6:,NZ-T=SLbRf44X,N\
BB\bS/(>eZ3_ZZAbJe&e2W(EM<S2]-adOX--FaTYO7<N4OU\Q62aLKf1\CGf2VW6
C>F9?GdS2=Pg_M<F]7P9J0RA97TM7^_Qf-V(+&XZR0B_+-;V,eU<_P])OI_WW72&
NcJW6,)/YW/#c\X093fC7-29W_T7<#24&TRZ2gK+]]R3JYK4Ze]J2N(TN_-==9;+
g>P4HJ^I(>N?[I-1I9:N5HX^#4FMS@T64_O^/7ZXF,]B?f3B]B4S\N;d]XL/E0QU
d86ORZYef3V)9Ed1QcZVK[e03M(<aLP_aa&8(9PZVB5eBIMP?-K#1@):S><I.0e-
K(V5M=),7([0I_<7VE<MI9LT=X@0G#Ue<AMD6#,ST_Q9eW#T+b#JXAEDJ[ED=U=]
4/>a\[G7fUYZc)/>BDIO(,?9&SgA)U&+<1<2Se18Ra)Y&e,(/4D7QPHYe3^H[5AD
=+&bb+OS;K^18&<d)b>9]?FB41]H8DN^LR\aOB7P6</e/5=K157)#IML1067e:E?
H:O).9YY9(-PI:Od9<Q-_,.N&G06g.?(&N2^[0WC:4]LcY[c5J,+O<P8)QfVCCLG
+;SCJDfE??^7EY[gcZA^Y+H;1E2+I83ZWUZDOe^7gL[U\5Z+SYNbdL>Sg;<JIDM;
#):5fA9c<Q0(8?EP^SB?JE&(W4gTL##)@gW[b?2JC=;&3JOOE20?&\0_MVca>VCb
9@J?IgZfR06O8]KHbJA(19&\5&E^F/]]CN(8UOJIJg3b[(F=2De;\:8#S43L2CYA
X<Q7JJ-b?cOa5BEfYKaXd/ER<Z=?N@gEI8@:KHA85+CeA7B]KT58;==AQC1N&GJ:
73Ued2Lb54X#G[1S&PFORIPJ04a<2:XD545A:eRfIV#])11dVK[5^MUJ=7ND0X,]
^_3F:.WN6Hc.4,N5d)_]d7\0D9U<edC9^.3B_b+M)f-0W(e8ceW7[fb\.OFf:_HO
2^&T:.7bIf-L/Nf#>cc?SHbgR@IbRJC.=R0N]^KT=;[5;KBBO^VQfTS>6_bfS(7;
PKE?_eZ9>MV2C?.LIU4B>e1eI1+,fQ8/eR]8c(a(UP]Ja=ee1/.PZNB^U/9FJ[60
0>-ALHMZ-JPaL.B)c:,]-N-fJUI\;+FSJUb<X8d#1:Z19Y0@<C=@/_b,b@<M0g&/
cQ?M7)L,WLROR<K-ZA?O=F4Y(L5]S80N[5LXa9=c<@YVd[##0Y3@=IXDZA87ZR^:
@Z_&N)U3=;HbI[+bC[0M<6ec?)9Oe-39JW:;aX;XPXV8?R7/O9A/P2(-fW.2,STQ
(2b^3d2UBDV@\GQVFRAK9f>ZaVL(;H9NH53;V#&WQT4)3Ga^^?6(VK+7AE;9bX=[
.\IeDe2W[#:)>KZE8A3<.ROKe8N+17.B=/^/;MTZedNW]?_+F1Wd-1\b2,_a)Hd2
OAU;.1#:F&U[6=OQ6:I:bXdDe^M_?8GG0(SK7MV9C?E&eS[U(:H81fg.CDPdQ1<V
>EAT=N))=]5BE^O,7UgMAQ>T0P+>O?9Q;)31\LH2](cZ\GDBJZ&(SAGg/=8O-9HC
JYI8T9A3QdcB.WM0M37S_;#)3+AND4(^-5\REH88Q<ZHQ5SPM7X2BVbZB9ZH874A
6GEV^0I#.aR_\-HB;R\R^H@4PQccJ<6YI>K\FaB\@1VF?==^FJ<d14eAN\KbcI7B
<QFS:];WCbXEBO0aB_IG]2B=Y,f_A64aI<GReO/5@[OB8Pd2Y.d5,J)IYOUID<KA
J=>XXRNV.>WQ[786_--G[0T;J=;@J8V0VEaPGI-^=RcA/LAFL;)OeN]^93g^&SaH
;INQ-@@.^_+AHG:Nf>8Q#LW[,-_(>0@=T-[UQIgd,B;E;3B=SP;NEC,01L(JCE\^
Jd\-C\fMc/A]Mc[0F3O75HO2(R2_9X_(X/3C\8:+9]QRd)0-RgI]L,9NB,\ZgcXd
BJ:G\=,&WcdY2&dY]9(BIJbD@-gF.QR_..;]dO^ZX@24:P6gH[YGaL69.H5&;[Ld
9cFFE5Q[.FV<]e7^-Z+IH)+X6C=d2:FX?\Ya0>41:[3)Z]O#P\CM.X;FV5T<gI_.
J[A?K4f23MA(K=:aM85+5]^#Rd#5EWU;bN@/C]_<)9.(7/CNcgM1f9fC0G>QefV7
EEf<Pc&fT\f[gcTgIBG^B1;(DIK=+FWbg@#H?J#a&G[>5/V>]a6:==:9?;\-e/=>
T:a<#W4=,9RKRPcO37]FT[T52ELHe\6e@8;73ZMW^]6g6XS1TDG>336EQR/KK<fK
R>_CeBa3V->8gWM+N+:.OP?T;5QH;#LO-RSU6M>T8()R.S6Y,3e3gZY&g?b/T-QD
G91)<WdWI<^IXZTX;DVfU-Z^b<0;\N4BJg=b5PTYHM8-,#S3GT+[J1RJ__g?.1@c
=7QB8?#A5d75>#@6P44K8,(9g=SMb<bbC\Cg>O,V?Rg/\Ua_S/Efa^>,D8+A+SLb
WLNaZbQbI<1N_D4PY7c3_M(B9+D27D:KcCeMdYMcJ52d#V>DC1.F,[e?Q5Wg/YHg
)5eG7c8\V+3fK4-&FF?)d871_,4ERC&,QH=@41TL;3JX-6\12E(3KU>,g2g&gaXb
B8FDO<[Ne]a3cQY6T+g4;A#1]GaeF//M_YaUddIf#860Ff0Xa74TRO8(BUZ?A)Y4
IWeZW^[HQ+8TX5YMdb:C;M1(A3H7VEc^B2X4ZYf,XMTH-W+b0U6)N[=36L9FIW4<
E3ED]5A\IVN@.^XO2#NG()c0/2Eg1ZF_T]V@eZ_@8ONPB(JCR4J0^W;AU6<,]O<<
Z2(0.1GS<Pf0QXAZJ1dGMbb=a#@U:_U59=cC+Wbf&?9+Q]:g2L\O^L]aX:BHI-6=
Y9LY@TWVN)[,EV6<MLFH&@3B9d]f=SN>Za8OgU#ZL_RI(E/B:3#F+76MAQ352JE#
3T@V/J>AJ;)Xc#/PJ:Z@[c3#U[;/3WaYZc1,HPDf4a3ZPMZN>2,Y+3BP=A]CRQ[#
FDXc_aPHWOZbc.LYDF#QV2;CPJ/CUDBg&QKO3PQQ_:=3Hf/g.LaJ,FHFT[PcG?QN
1PL0BIRe,CH[\#>g4]Y@B?=I9BVd01Y7=Y+(LU9\?T:Y-/+d\Ng<V_bgP0ZWX1:?
]G>McIH#S/f=cD(Yd-ZbO>SP8A(O1YJ.=&V.@TK.7E>5^24;7JAX9UJ&FT#GO6DD
<5W.0Qb:d/8K:,YSJ9/dH]YHaYR(Z^a1c4a4Q8GU]FJ])=Y9&?6d7F<&BT,_WM50
06LgE)UZ]e>[4#fX9W[0N0#I=P+Y6(?KgANN&]O8gPKZ+gd(X9e9(JBOKJZ+ORG<
F8V<_C9I[fJ(,&aZW&I2Wd,WaSU##bT;.2Q+0#b+G+Y)b@BA2X?gN6+S5Xf?0/MM
)5M^:TG4Qe1Xe6[VWdg.108I22D+5Q\8:5Y6.;]^;FQ36(_^+>]2&P5Z_^CG^4DO
OE#=#^NBd\M[3DG=)f9++D;AEWJ0SY/H/g2P/KF<BS]RL22-J66_A(E2N-e\BX[[
J>U^7Cf<<8LV2fN[fG>J85MD4Mf=V_/_P31=>O;;4E<I4^LBfgC4g-a2_./2,e4e
@X2]6Zcd)c]V/b^0+5B75R2?[@QOI7g;/bFPfHb,3WS\O,BZY9Da>0/0>YP95]R5
#+EcJM37RU7W_O/g(.=K0/1.E;2AQ>U?&TK/K0ONZ8fSHFeE,FM6G@^7+6QJV6TH
aLD#MYYQX+TX0@_JCZ)UN50b?YAC.T0V6CIfAK3U?L:^S,F7MMY<c&#AF,V+CIME
5Re2I+.&gLcMO.<T>aJ?f;g5Od0SBS8LA2(MQYJ0VSE+7&9BQf@cHFPfcJM1Mgd7
[^X[I58=Q1/W3/a3#ZV)1.[[/OOJ+5SGU5]6ES5)&O]Q0.fEL8><O^^gT2X=]+#P
:AF[U9Q]O3Sb2;T1.AQgLBQI[EBYRB>&OUFM;]4#EbZ))d9=..JBbBCC@MB=6N<5
ReU7-ecS^5ZA/;JeBL1G(2)L,G(:2E[]e<_\8YDHK2c4e>=-Sd5F3E;3DJ:(4WAY
ZT7R[\eW^N/IPbLfX?035]b7F,58cTU,Ta1#(F?C_]Jf\R_1I/UJ;P5<8Y&/c0WP
e;^1L^NKaT)=/6VcM-GJ&Yb[>]?FH;JKVP-I\b<5B80HIX#;1:M,SO=Xe3YZDSRH
_XG,c.LI?;_&)P^O@YAO+;HJSNP5/YFG_E?0O>OS)6e-R[HU1&7/=/<(VGTJI?UJ
U/\7J^N-eg0>ad1L8IP[MDgff&5UD[EG;A\HcQ3UJ+&.]#?b.c,+2^BaA-,RZTN-
:-:U7:04FHMMFf&a@S(V;U)LBMMg8=1T8YRAW/^/[fY;8)2E7CcTM?(dNF9CJ[fG
[BCG3\aPW9d@]5U1]4g^1].F:4N_fD4e.R9M.=<X#+9VP@2+V1I0/^e42F:[</4f
<EGDM0JQDBY-U_S]-DYf^O-dC,TV,M+53<;_KVCDOgX(d=O3@W6dF-#D:4#\PWb5
:ZL)X.Q(=LL51F9\OP-e3)GYZLOIU,LL1b>P_dVgb0QNDVFG&.2##R(2MdK0gI,_
eNF[3JY4SFFKT;fbB:_VQFQTgCZ=Y-C)R-JVXaKb07O]4dD>/@4RBN0C[K/&IG^W
N>d[<-9H9P;dKY=YY?MD1OT4a>R-\DZYF_,GedXFJ[<PK-<^P#c-S\KbMX,>]KBZ
<49M0)eBV@^(-3?>8.J:<G65@BS&GIZE];,4)Y2H1_77]ecbWNG:2>0WY)FTG\,1
Lg#4R6E9e:I?E1(W.&<1LJAA)?940G.HF&G#2ZHE=0DO0J/P@&c?Y@7^KBAW:L#,
0F&,R[f)<cRUM()OaFWN02=)4K=&18],D]5_bE.5&0#3>g8cTK>]?YSQXY;26>)B
BY0C=c#3IeCQ&[F6(4b7.U&B(WA[62WSg][c/dN_78eVAE[=1dDT5J8UA@M@QYO+
7<JPdL;3_.LJF4G4VN76?NIMF3)]EI80E=35KD1,Nf7#?_Fc?)-[?[#PH\X.6XYN
#c#1>4SHB(ZCbN?5YD#0C>3EN.QFX:<Ig<-FATF_cYUZS?fW\SNdd-1GT<BB1;&&
TaO2Ha_59<X8AIVf2D+-H3JOVW;aPMg78)I]/-#,^U4]]@ESJKQ#NfbT)#2A+5M8
UQC2_3YX>#.8M/VY1Ce?_4RU/85(=B+]D05df[Dd?G1G\F.6f1[VMPC6fCO:U6@]
:3CW)S_c3LZNSV;=Z]aa@f</NVZLMH/>4OD0/T.-U>B]1<];_#Y+Q)=,#+-^N<2]
Tb3KB[US(>-WSReWS3a:)8_&=2[c90=@TL@&R<aF\LOGecb3<GcFOb[>[\_b19:B
6^G]H2__O\L<.KB3,d4HDG5PTKN]DSFEPOGgY_R)<4F;N+4X#Pf?NAYFKIM,F.WQ
>.8c]5RNAN;U1D\-O;bY/XDaT^fe8_[_VE<\(ZCAcbX;3-0]9,6X3a&bP,Y1[K^6
5)PdQMB7CH_JKXSgYPXC/BcA2QJBd7BXGF5:O#U6GW7M^8H^dR70R5N7G[(AT^dV
S)1K0D/+3-L:bML?cSU+#+.VS.GZ<bTIV?XadO93802U(:#GK1>ENUd^^H5JPO;O
ZMfcb\9<KSFe4AfU2FHQ&0Jb:Q5E4<33c7/D41&PYJ3)M2DNB-U>8Z#LOKJbQXE?
JA_KaWe_aQTVd9PKY35&;g:;;L[GX/C=SR8IU@afAeN4V->5\?A():_N/>Z7V8_d
cW.K#BbFREK&AF5:HX&A[_PAa@C2]MH<S0?^-U:[)1_bcCJ-1YJFcW]Q?0,#UVK>
WKAAWb>+@L+[b98?-S6\ea0^cA?9Kb-)bb8,#F]>O.#a@LDf59:9]0WC[5IZ&5@^
e#7.,gRZ]N<L]=O+G3cQYXG0)CY/[@f7]51EPQB_O9X_/\HeK^&KW;;6Y(I#b5>M
9;NAg9fSaEGeIM&MT]+O/,2TUag+Q5BAL8Q,I<_e:U_D:?;7_ba2<?=++;<1G4L#
36Oc),2+8d.&HVHL]c_1-<W=;a)[G^.fN)RF&-Z_GHcU78ZP?>PI.5DFd>c[,BO@
F:<Ceb9VW=W0@Hd85Bb?>K7f9BOLOVHHL>75=g853[:66(T#X(TKD9YF(DRF3.ZQ
]-?f96&Q7:B]/H7f:aPc+M=5S#EE\3IG\<N[e2&2O?^2^AgWCK&^8+B40<1K:65L
=J.][gP5E+Q_3.?d1VD@1?+2/[Q3BJdS-L>cdEHZ0UO5eX?/>2T\TF&LZbWVBRF(
5UR4Db1CDFUKRO#_&fLJN3Ff&\Va#>A=E(&dU>61Y15WR:17F8AY-IM_Y1d-+ET^
::BWa<cKVdSO0+RSE29PAc/3Ce\_E#ZN;W;Yf-S<4U@0L-aEB7X50,.3C.[7>c33
bU^U8M#DZKKb8N1&VPf]>f>]F;9O^FQZD,<B-X4B8RXNQY_LI4:EN+=6FQZbL-SM
fX6dE>Dd;AE0>gS8b->Y<P,@4+/a?2FBF1@9ER/EG0)g0g[.QV/<MbE;+J;U-bA2
3U20-^BETX:L(fZ8920Q1HgDO02.L1R&ZdL08PgfUQ>1FXK?>.W#F63a&&M1&\9D
:+Wa?DHXG@D1c8(De#P1/Y(D<K,@V\f4JT4B^<fb0M1?a&P_AaV,E9=B4cRgKR69
76G32(G=FSbP_AI:PKT&9]UP,aUMN/\,CAQTg/E^<C#Y^Y6L1K)95_&fG=B)T^R4
N#3f.@MG#HD9IKN2>ZZR63,TQD2RJIc[OST[QZ3ff9:(#IF,C,9aMOZB35<#0R<D
E<V6M1H+A;RT27]YPR@2N+<:6VObT=#8Ug0#@V9VSTUV_N3Q+dd?A<4DBA^GST,P
_2Ic+(=)ac0#9TX2IG?_<2C;53N>]#8ONM,&9+6<X&^@#-BRFJQ9@U1BNe2ZZ+&F
+&DMaHO5X^SG1A)AaBdV8#XB[dbg&.IfSKT>0UI:9QO7Q8Q0^/.AWQQ;^I#)92D:
PZ/O[3-HX]82Mb/;)F&GEc_HEY5XW4eZJ;;e0ZV)f56]?#+;OSbfGT]3fg4FUf/E
MOb^BRLF@9f6,+SH8AgX]-1#M44DWF1V4XN,\FdMgGOC^TLGZeKX]WbXg/aR&_A:
(X)5>UR=0:L1cWE(D3F@Vb3X6RN81?_0_YSJ;YP/[3:NHM<Pff1EA+YIaaF28JdO
Nc[&<RO[[2:+NO2b[#QNS_?UC?91:OBTf0<L?2,bg]FS0H5@bg>7e,\J-0M>Q]T4
(CXBDFU3b;0]d+@.fKZFTT2&bQFfO6UGMgZCF;#EIZ9HCK08BBP?Q68UVgKJ/>0\
e@T-/L5G:,_Sa<[^TOUD3UW48:_=fIgL0-N[54Qce./I&]7DK<O6;-2R[5G72NX(
TP/38#4,2bCMZ&e>]bG=^-@GXW<N&a+Q7GLYH\eTVI8MO6O)GNN5aEXB-V5V2/^P
]Y;9e+2CK>-OAAUNWKLf:/B+e0&\Cg:FDI<VdUc9)K--76QW)ME][cY5&]OUW5EW
BBGJV6fH+ZZ,e>GXO6##ZUJc9CFa/VUF2T495SQHMTPSPH6b[HM)<9&7\M_g)9(4
Y/(SGb0./89S::0[Xa.5S#)47200,1/_gA5-N\37JPIC7UYL_7E<F70W.BP+XV)d
H.:SO?1XHX/XYHReeE0/U81@716NN&CR&A>6c4f_dbK^@C(MXd^=a:33X[PA78d<
<daUCPWWWJd0^+RS;T+&/\T;-?UOR?H)PTFKb-,EgMKfeB(?,4)-5CaHK>MdZAT-
#UJ7faM^KCf8:AcOWBR_cP^3NRRag?S5CL,R5=e18Rc:,C/G;eMS:4C3(JI+T73E
)[>S70<-MD8eKK?KMTEd0/UfB.R&ZXBI?<J+3D#3\c<5J/gYLd+Z[g10J)MI5EUE
TVW7F0U=--95GW=0P#]#&_#9/,V-LRS]f;A)U-PI1R@3=RM=5DfaUSS8gJP.-\]A
T#KA:Zg2B&<D4]_G=U#PUK/4eOX[\gQaW^W;XYT4<@VY=X(N/6FR>;JJ;V4-[RU:
XV497A3Z;M8@D8/?HUXNFc#8#5gF,CeCB,;L/;5#+4W2\HB@<IcWO.(F_6FJdBXE
=\SR3X\0=1;D/=;1JeG@[V&#Mb]K[2f-2?G7);&#GXe_>P];_8a[G?U9AY82e55a
Q[H6:ANK]5(#a;VI3[V_M>4:.4D;B_OOfZ:;P\P3a-H&#3/M[0Q-d7&>IBMCS&/I
A&EP-X&JJN&8U,5bME2e>DA1+OWZ/faQQN8dF(W,..\5#c^(ZR/J(WA?Z9cND\1+
R;;398a/IZK=+d;DXQ53C?E5.6/M>1BH#C^+3+cc+33.c8).ZG>NDNBG(C^AfN9\
&(>ObKN?=cEU1V,dJ=N@RVS3-c)Ea0MA1&bd9a/c1,:7b@B6\MJPDbM7.&G7;(;b
U@Rg38RbSIA@-d5ac]=3eK,98<gIU(W/5_^f5-620]979fQbDWZG-FTG&dFA^+X_
BC7F]ZY2ZIab(cd,I?dZ#EGc+5WaEV+3cMKD(/,\B56)PTKP([XW?BL_D,P:/OMN
)?_L3E+9FDIPHP[FIfXGdDA6S=aL,IeI?Yd/=c#a6-.g_I7K\<b-3^gH=S-/-IdM
e]g?(>N<4aTC4;,S#B8I-=FKJ:_Z^Fe9GBN>ZV=#5(_?bMd>I>IG+]g;&TR@M\IN
Fcb\7/NZ.VB+_5[#._&a,L[/LUX.6T]eZWABPeGOR4gVI(4bLOcK0bcHGXNQ@:PY
:_AD2b2()A]2#6T/cc([:(TQZ<WIZZ5d8QTCd2S@P=^HbZ5&&A?&W\_6?+W+6dcM
H+/I;#cHbM45RSO,\.X0;+>#g,\,Rc^&K=@7fc&J?GTb[cd2.&V(JF#298[PIfX4
#>:/>HS2<DAB49f]7Oc5L8C[=<#9+4GIBFVa3S,5=NbI;PWgc[:<?cP9CP[//9K\
@(A0D1.8eO0cPY:ZFeeY?)--DWd]PKXS=Z[\S&<WF(0<[&-HY_UVV>3>=)2]dZMC
KLU/FWbAgC5a?/S[5e.T\#^:32[gI68+QB=U\)E?).bf[V&7Qf@Qc[&D-YGJ;7)8
D=:CbOEgT3WDSgAcC00=-2GVGb^[4@60,-MH0._gP.QfD?4F>/;<e>W?(2#b=T:[
OKQfb2F=<:0?;g7[3)9#_V,L4X\AA^#2DB,K/0L+2[KNe&3b_fg1[:JH\1cf2,]X
@(UU8TT(M?YTILEG:OND9g./(f]MJ85JC@)8WHDHK[DF#;^O(G<Uc][8G#Oe44E3
97<5T+;^a9#OO00IOG?fHK@(KTe1?]=<VE&>09+S91g?V#^>?_d9Z5#-OD]NK63D
A2,/UPAc@OgE+>[[C+gM#AL?f@QF\P2,TEX@HVaeD?M3Nc^954KO-M<6aU#G1G;E
H[7.f;L5PQcU+/20RGDbUW.,QaS_Sg<:eWd(E;TDTdVGc-UO6XR8EQ9>X@c9-D<J
#=](Wc+HQa=.6O=L.O/dEFVHO4UWYIfKVBg=.E/_5/YF=f,<)f=:fI9FVb<SY.FB
YBF/9cEZO#W6FaX1Y^=EERTXN,8,(^4(TU)ZQMIdLPYTS0:8egJ<C3^1<L4:Z2.>
ZXaada3<L5c4R65M1EgeH]dNaO-dTNM_M?W83O+R<@WF//]Pc8[&IO&5gHL#_ZHB
_)ba8[E=<+f(J?QEdG+gHe@6eQ[^SAf1-dGVL]/3).;;63/&Z+9:Y@B]77ZZdS=&
dTQ.:aCNE\^GGL6ZK>P,:4(Xf1K/;3TAeXHV0cWgX<eJ=8[<=K;ZNT0>4db#f5bH
XZ9MV#L49ZfMTRT+\;-9XeFAP4^Q+QV0IY1+@4bW#?UPf2CG8)EQFFJBdF6\1YT=
ZL42LC/2Za-[#a5?PP63edbBY2KEJ-1):ed;XbSO,Cb1egPWeT90P7(+f7:XcFT(
+1H[QC&F[3Ha[^5E95^]#10@>+bX,bS;dH]D=//+/F8PX,b:C/=Z)]51I;ge@A.,
#:[F<a#]>\;fW9N#+e[Pd+KN]Y.\^IT:TCO#G5Hb9+QQT3Ra0CJ@W&MBC54E,B>Y
\LXB_Tc&3NJb9@_=?>].42BZ[_13\b:U?Q>OYD-&F+GP3J/@D<Z7ILF#&\QB2g^S
gBG-A,EN5Q2J,2(W&Z:D51K9F6>8L14;+TK(I1>L7AI??@F=H9AX,-U_6P)cbTS8
=;Jg),gYEYIN0C/V0AW.U5SEGEMbAX,&]L3=H1SI=8VK_,B+Q?:3Y^45eU\[I[-K
e9X4)M34(?QWY@88eeC;7?4_aOGGePbB9[KUC2+9]RSPW7&VZaY/SYU/4g.Q(Td5
^]5;NZ@8O\WY#_L<=1ddQ70>X2:L-gE1b>^fBO]dFNA1?9[I(KG&6AYKU>VCRM5=
0SO[@b+B;_2;OXa=LTYD,0Y0Q9=,gT1F+e.fIUAI_+T[0bB(JMPUAQMI6/IT?8M=
2Y&U=L7GF?B&=cZK[J8&EZAWRUZX[S)7[^7O\_<+)T9A(,NEf&^BCR>S95>Z:.T\
P0gKZ9#4)1-\Q?(?FOZaV<-e0?#,]dCGe)N?R:OLS3N.,F7[e1-A#O:Ea&:B4YY1
^1d9@8HRP^YLX(5dZ]8[_L8.<V;I-I0&9(;S^A/--c2Q;XHg)OX7<BDI=DeY.cFg
KCI.[HC+V9b6WG=gD#3MUd;]R>.>]1fK@&]+330eMdH3b>8_Vg<J&SB]8c2#FOO\
bJ<OGDX#E.(IV]5O^ce6VTNY8[A8Of77d\IDGdaYQG,b1O^\QY];?8Qe:8VNY)f_
-L)\AD;@WZCa_52eI/WVRC8aM+)gEL2OOX+4?fb)JIe\WZ?:Fc9eBG<J43:f/H)T
F3).-+=S3;.REA3\^A=M32CcBW=dU4Z0a^99FXIT6UF;:BBC9>DB:^D>XEOT&D_Z
U&R[bMHA?8(d:B?[a6XD++((3O)MI3Z)N=0VCdb]Q?5f)Z^S2W)\7:V7bVE.RH./
>,(=\-F,@K_Y8=#a:a3<7X]#1W>5QWKJ&O>(-8N]/D+I@QA.Uf@(G0525[/12]8J
VBACL749YTVXU7M85&aD+NY0BC4BaJ2^.Ug6RSRFLXI6D<>3e(e,P\#OMaXbVW.@
D6N2>_<I0Q2Vg&P:>Vgd.E4O-/.[b+X:Ig]DU7c<+B,Z-^=9#eE2QOJf#)Y(3Q(4
.R/Z^Ged^dg2F+5;W(],Df+I2^__RGH931Ag]D2>D34<.eL9a_T,;L5ETQJM[OYb
34AJ1>8D[XY[MVX5=4TA:f\NB+)?RWe\93?RBL0OX\:[XUWeI#O.XPLg4<D?D@T_
M.FbRA_VBWK[:H_,5JLW;TQ5_##g(CP0WeV+6K^22cKF31EG?Hg&FA,S567&d76J
6]UMW@,6_G/;@XU-QC=EeDQEA-e&+@T=+-HSY1XJ&3QXXEP#cYEaLDV&fVIJ7X>3
X80.^#-RIeR1aW4E6U&SP=S&N4YYGM0[GE_e.@)<LeHPf0_RFBUU2A)VAO(G(FeK
@c(YH[0-B4WPZ_I@f1)25EZPQ@JU+fN<X7bC=gc]7#W--<eHE\6\3?O-OEDL[7Z<
?.ZdA=Z8^LQ+>#H=,aHVWLUE#JKgCLcf>SHC^/=N\F74;/?a8U?Va(^F8N5+g?8[
/9dEPgJF+UFf5IS+1WQN7RYYLL(aU(S^e\CW#=YdU&GGaKRWHS&NQ(V=1,Q)[^^A
b2=<b,;:Qe\g92Z2AZU6,c[@Y^<cZQPMeRSB<9XL[>\XD_R(INBA0YY@^Dg>;K[7
BRd&1C@=)M#3/W6,9Q2#PdeGMV;SOR>=\,:MEa64L5Cd5^]IU[ERMdUTa51OUFN<
U=.X,dM6,J?,Y2)VJ11KK5RS<BPGMYXT^7ON=W58eMZZZ4IgWHgY@X.d486FL/(0
QDOP=J0QZd7S@@;IA5PHe&&=Jd=^M_a>M1f;N^I(+0\d;?ITF8,B>-2AH1TM-Qb&
a.^d1)B?:MZMMD).ZZD6B9>48;J-YD-\=G;_,fFd;,N9+(=O)&IFAdeF^-VG^AM-
2\@Z2#gTdNJfMf8WQ2:7.^=[A\4I[CG5cZY(=PaPX?Re2-M>Xbf]#BMIGE76U7LP
:SU@+4V0FH=C-]4:2,&=gR@\5D3_eN/[HA>^NK?J@&(9\9\O.GZ&9U=^a.g^5#\>
YZ+C(I9FMa[H74f4V>E1:\+5NJB<f93LBcAEAN@ecHHQQRFCNIMWAMLCFVHY]-:N
&f9]5GQM#=LN-]dBX/A8(JME3A8Pb9K<OCL+,E9C=?=eH>IO5=T]T.N&?=NfD?YN
CK?/0GR@Y_c(A:eY#bT[+Fa.FPFS5+2D.K7ObW@#?,42eR0\c(1YD<&&)QD\5Na,
S<Y]3V)7]BAN)5L;_>9SYdLBAT-C/D:/V1JU-\V200HI;f807)9/V@Se8S>YL@7@
>33<C<Df;eEK-c=NDF/Td6bQ@,Vd;+Y]=NF)9]:^@Y&B](2:?bB,I>YE>H(#VUPL
gQAF8-_KX9B]P2P9,:7FWWfg1W@;6GP.SY\0eB@gR;E>_YaB(S3I8-DGM[@FK^,/
Nf\F2B(C;XK>EIMK#KG??;MC(V?2gP+2M9KdOD1Z]UbTgdS^.D1XIaS3ESNGZC4P
0B[S<&57:799W04)Of37OZ+)&3)[/,\CA)dC#](_b/RUGN#S?PMZaEC/PW7E.\J9
=(JI\O.IdbI/L9cU^P.R;?M::B.&_Mb9^)))@B)6H1KBFC,Lc>^FQ)ZC>JbZ.F+&V$
`endprotected



`ifdef SVT_AXI_QVN_ENABLE

//vcs_lic_vip_protect
`protected
MNE-&_&G6]+0?WEPbD3^^AS(K?dF:E.+&Q4BR]\UZc;A-E(/L/916(53(NR?bC&&
D2YGY@/<Mf-OTN83+aGCXC_df29GZQ)MER+g;CD=bT&_Y3Df13.dVMBL/SM=>+3&
HIH-PRRFGPC52_30b[?DZ8S&0)5D=LLVBA/#/e/04;Xa6O:R@bOefM.XQ2TcY8=M
^UaDf@6+6:f;[9#;DeDOe+Ab=_S4Fb#.@:LQEN[>KOP:_e@Md/7>YWA+Z450)/:B
L)64,A2R?#WeTLH[+9g/.:)e5ZW/\T<-851D#Q-LX,CaT_RGeR5Z53S+:^/LPI3B
((G=\5J>J+0gXODCNID=W,ZdPRcgb1SXLa^R4+c</S0R\0I-@OQ.;NTNg\:B8)b\
9CU:\TA[=0H^+Z.XPZUWK=A:.C7V5Z.#84QF7MKgAV#GFKC-+BHcNb]+#_R/BYZD
P>.S,\(KVI30P<8Bfb@N7G;X]A1.XB?1AZEQRJgCWV<R,;(ee1),Zb0UX>eA<YS<
09KA)-\AHJ(1N@MC_b5fK]M9V6)b0&8KBSJE>D6C\f3-?P\1Z;&(Cd6WNBDHU]2Z
-VFNZF>[WI948Q(d#@]I<f+AJZ1dI.:C/KQ@3A/4,G/<S&K<R>]33-ZP/:B0Ea<5
C_>2T]F,[:J_9\P0GY\I&+;J+fG\AUB>BCf,CB_J1Q;/0SPRVN_RCfK92R-#K;VX
FIB/^O59O]b^GOHRX?b9E7)X:S:&\QAIZ/L+aCaaEfL^2997KMBM><5R(d;D.BIY
/P83P/Gc7I/PDfRNW:M[X,Le[L#?b#X,S-)2^<cN:ERS>2LR#[(QWWFEI@X8L2)1
SNeJ6\Gg(4Xddbcfc(EO>:TM_-=V>cNH4N&gISR:8<d;EFRfO7&AQLV0)S:N0G.L
Bab;2@)\&S/7N[6d]aW5,G&V<6VQD-S0Z[U_[?3;3AM._C]4@[05/Ad>;PM6[bVB
XEP3#VB^KgF#2<42&K#PYEJ##7CM1]F:N26a9#c2>&KTXQ7@_U,aYMI#XIGQ;-RY
#0U9)dWc/TDP3e/(?3Y>(>e)X>,TaEeZ].PZ+PG#fA_\7V2_]A8JaFBY@OC89M.f
&I]SBO+I1UK#8M9MLSH9\c41/,H>AA??X+(&f?G,;YIN84C+GZ&@ORE<LZ63)/B<
Z\8&/)AJ9YL\3O>;C4QB44R&S6E,3B3aUJXI:/S_XE7))H4JfH?)3(&.]RS9F=5F
;9BGeM:;/);#D)5YfFMA58L5ff[#L>1GQXgX&/NG3<V?A2:#=E&+7;SQU&.31fF?
\G=X92C#,B8-L5BCJ\-;+:#]BR@PQN<BEKcZA/?dSF;E@QeBD@>Hdg.TQ;]]cYZP
A]^1JPMUZ>C>a@eBGe2K6IdN<D8=dTEB2D>JgQS8[ZQ:f\bK(=,&/[7b6:2B(+VE
?8WM=<=Y4[)_.JdUC+/^_6M8I&6S19FX>+K>JD:6I6-SVa-;]=A.[E?>MVEHJPG4
^)XK8LIQBB;R,\P&2J3X(BJ2B#>@8FMDM>YO5)1LM\=5[b;==CTWRY);+JVHQIgM
LS9]QT,KTQ2d)/V\HY5-YA&K5N)?U57dH1cT/Lg3N,2I_HTE9FG7VKY4DCg]X8XR
W;d)\7C(K;YSg4DNS?F6_Sc<(?S@Y+A-fVaG&KgF^WWd+\H&WZPO@K?<2@D::b.H
8+?E(L>FRW;96:-Z2811aLQa9S1&K=]>)DVARC&HCa?Q:?D0W,<A2U(1T/XZfH7g
DWZO+C,-aV7IP]8BeaO54JNHXCD<<WH/2^c^9>3S2UBS_,(8G6(6aIgN/5:,V)YA
I7QQ/,MU=0WR:4[<V7\4<RAIOf1SWC[[1dS:b>X59Y-(gU0fNC?5VFRCg2CCaOJ,
]F0U9d\EC70c.-g#(&YWSSG^0b[>]>4,ePFg64+QNaCE<;D2C8,?E^MZ99ZK>\9;
edP71CDI6P,,@DJ@J9LQ7K(IMIOO5f/+7HeNJ;ZVAWAZ9)+9BPH4<.]SXGTH]/a>
02T5>/^+=0?V,M4PV3aPaDF]]#N)K0HL8T0\D-4Z10f9YB5fgDE#3LM^Y84\1A/6
XP(54-RH7XL5W-CG3A.f;=FR4?VPUb1Vb;GTV6B/_,#?=A;O[>@?;HBaN;eR3Y=6
9I<Y;I.GXb,8POB-Z]/>](8]g4SOC=[6A@(1;TXN\.7L&5@L)eH&df[?3@F-]FI3
9VR4S8[DUTWJFVM0Faf:0bO1VBT0L&G[DJ&DB,b.5G6]ZZMY#0K3((C#K<,./bH4
98R(6Qb\#VK;K5(g+R1SIB_e8be]]U:=P83Y]99M(52B3R?E(I@]T9cT,bJ(AXPJ
DBDQ&8/U9=[_dGUXWVYLeI,A,Y2VGUCTF^T+:T,DT[^&HM(=U:4:HU]WCU_1g.04
OZHBFC8)TeLDUB><#b:BL=Z3)CPI<C?5&.3U#D<W2e9KJ8I/T7#_GG4:CKQ#GH36
UX,6F@6B:Od#&CV?GG@8_Y^CJMS#FCU;6ODXON2&BK?1?JF92cX40b,f/T@G^(5W
&8?Sc]cH=Sb>1L-de9I_XTY7?EgN)\f4.CB1DTB2Ld+OWDHG\=CKcJ,Id)Y=AX0V
X#W@:&fUaDf;71IB>LL<M6M3JU3gM5+2AZa=.[6T9U,&d\aTO;T^B5D8HJ>Pa;(e
0e[+-@eL6D1gJa3FL0@_aFJ)A7eU+FE)VO-\5_&\E-gb:W@:96eXR&D8P$
`endprotected


`endif
`endif

class svt_axi_checker extends svt_err_check;

`protected
FE)5V_QaE)H6F>;&-+6]I8F/VG:M[58Y#@\C#V8EcX(X(e5^0#F,0)]EIf#R6[//
.C+1KIE&YN^6/$
`endprotected


  /**
    @grouphdr port_interleaving_check Port interleaving checks
    This group contains checks for port interleaving. 
    */

/**
    @grouphdr trace_tag_validity_check trace_tag related checks
    This group contains checks for trace_tag feature. 
    */


  typedef enum {LEGAL_TRANSITION,
                ILLEGAL_TRANSACTION_START_STATE,
                ILLEGAL_COHERENT_RESPONSE, 
                ILLEGAL_COHERENT_TRANSACTION,
                ILLEGAL_SNOOP_RESP_FOR_INITIAL_STATE,
                ILLEGAL_SNOOP_RESPONSE, 
                ILLEGAL_SNOOP_TRANSACTION
               } coherency_error_type_enum ;


  local svt_axi_port_configuration cfg;

  local svt_axi_transaction barrier_xact_queue[$];

`protected
,</aA&R-.AFE6RcUF.S?Zc@bRN.A]W&7T3g.Y\[5Ycf<T#:Zc6:M3)(V7/-A-E)Y
@#O@)c;H:9eE,$
`endprotected

  local string group_name = "";

  local string sub_group_name = "";

  /** String used in macros */
  local string macro_str = "";
`protected
9/@O.E7;>1)#e,<S698=;,LE.SI\PGb\55(aDMDac=e5GE.6&8J40)NP1O__,dcC
U:4^1L\?QFB,9[<A3-aXCTHeB494Yf>8:$
`endprotected

  logic previous_reset = 1;

  /** Delay from ARVALID assertion to ARREADY assertion */
  local int arvalid_arready_delay = 0;
  
  /** Delay from ACVALID assertion to ACREADY assertion */
  local int acvalid_acready_delay = 0;
  
  /** Delay from ACVALID assertion to ACREADY assertion */
  local int cdvalid_cdready_delay = 0;
  
  /** Delay from CRVALID assertion to CRREADY assertion */
  local int crvalid_crready_delay = 0;

  /** Delay from TVALID assertion to TREADY assertion */
  local int tvalid_tready_delay = 0;

  /** Last sampled values in read address channel */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_arid;
  local logic[`SVT_AXI_MAX_ADDR_WIDTH-1:0] previous_araddr;
  local logic[`SVT_AXI_MAX_BURST_LENGTH_WIDTH-1:0] previous_arlen;
  local logic[`SVT_AXI_SIZE_WIDTH-1:0] previous_arsize;
  local logic[`SVT_AXI_BURST_WIDTH-1:0] previous_arburst;
  local logic[`SVT_AXI_LOCK_WIDTH-1:0] previous_arlock;
  local logic[`SVT_AXI_CACHE_WIDTH-1:0] previous_arcache;
  local logic[`SVT_AXI_PROT_WIDTH-1:0] previous_arprot;
  local logic[`SVT_AXI_QOS_WIDTH-1:0] previous_arqos;
  local logic[`SVT_AXI_REGION_WIDTH-1:0] previous_arregion;
  local logic[`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] previous_aruser;
  local logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] previous_ardomain;
  local logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] previous_arsnoop;
  local logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] previous_arbar;
`ifdef SVT_ACE5_ENABLE
  local logic  previous_archunken;
  local logic[`SVT_AXI_MAX_MPAM_WIDTH-1:0] previous_armpam;
`endif
  
  local logic[`SVT_AXI_ACE_SNOOP_RESP_WIDTH-1:0] previous_crresp;
  local logic[`SVT_AXI_ACE_SNOOP_DATA_WIDTH-1:0] previous_cddata;
  local logic[`SVT_AXI_ACE_SNOOP_ADDR_WIDTH-1:0] previous_acaddr;
  local logic[`SVT_AXI_ACE_SNOOP_TYPE_WIDTH-1:0] previous_acsnoop; 
  local logic[`SVT_AXI_ACE_SNOOP_PROT_WIDTH-1:0] previous_acprot;
  local logic previous_aridunq;
  local logic previous_cdlast;

  /** holds number of databeat transferred over snoop data channel for current snoop request */
  local int unsigned cddata_beat_count = 0;

  /** Delay from RVALID assertion to RREADY assertion */
  local int rvalid_rready_delay = 0;

  /** Last sampled value of RID */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_rid;

  /** Last sampled value of RIDUNQ */
  local logic previous_ridunq;

  /** Last sampled value of RRESP */
  local logic[`SVT_AXI_RESP_WIDTH-1:0] previous_rresp;

  /** Last sampled value of RDATA */
  local logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] previous_rdata;

  /** Last sampled value of RLAST */
  local logic previous_rlast;

  /** Last sampled value of RUSER */
  local logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] previous_ruser;

`ifdef SVT_ACE5_ENABLE
  /** Last sampled value of RCHUNKV */
  local logic  previous_rchunkv;

  /** Last sampled value of RCHUNKNUM */
  local logic [`SVT_AXI_MAX_CHUNK_NUM_WIDTH-1:0] previous_rchunknum;

  /** Last sampled value of RCHUNKSTRB */
  local logic [`SVT_AXI_MAX_CHUNK_STROBE_WIDTH-1:0] previous_rchunkstrb;
`endif 

  /** Delay from AWVALID assertion to AWREADY assertion */
  local int awvalid_awready_delay = 0;

  /** Last sampled values in write address channel */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_awid;
  local logic[`SVT_AXI_MAX_ADDR_WIDTH-1:0] previous_awaddr;
  local logic[`SVT_AXI_MAX_BURST_LENGTH_WIDTH-1:0] previous_awlen;
  local logic[`SVT_AXI_SIZE_WIDTH-1:0] previous_awsize;
  local logic[`SVT_AXI_BURST_WIDTH-1:0] previous_awburst;
  local logic[`SVT_AXI_LOCK_WIDTH-1:0] previous_awlock;
  local logic[`SVT_AXI_CACHE_WIDTH-1:0] previous_awcache;
  local logic[`SVT_AXI_PROT_WIDTH-1:0] previous_awprot;
  local logic[`SVT_AXI_QOS_WIDTH-1:0] previous_awqos;
  local logic[`SVT_AXI_REGION_WIDTH-1:0] previous_awregion;
  local logic[`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] previous_awuser;
  local logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] previous_awdomain;
  local logic[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] previous_awsnoop;
  local logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] previous_awbar;
  local logic[`SVT_AXI_MAX_MPAM_WIDTH-1:0] previous_awmpam;
  local logic previous_awunique;
  local logic previous_awidunq;

  /** Delay from WVALID assertion to WREADY assertion */
  local int wvalid_wready_delay = 0;

  /** Last sampled value of WID */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_wid;

  /** Last sampled value of WDATA */
  local logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] previous_wdata;

  /** Last sampled value of WSTRB */
  local logic[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] previous_wstrb;

  /** Last sampled value of WUSER */
  local logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] previous_wuser;

  /** Last sampled value of WLAST */
  local logic previous_wlast;

  /** Delay from BVALID assertion to BREADY assertion */
  local int bvalid_bready_delay = 0;

  /** Last sampled value of BID */
  local logic[`SVT_AXI_MAX_ID_WIDTH-1:0] previous_bid;

  /** Last sampled value of BIDUNQ */
  local logic previous_bidunq;

  /** Last sampled value of BRESP */
  local logic[`SVT_AXI_RESP_WIDTH-1:0] previous_bresp;

  /** Last sampled value of BUSER */
  local logic[`SVT_AXI_MAX_BRESP_USER_WIDTH-1:0] previous_buser;

  local logic[`SVT_AXI_MAX_TDATA_WIDTH-1:0] previous_tdata;
  local logic[`SVT_AXI_TSTRB_WIDTH-1:0] previous_tstrb;
  local logic[`SVT_AXI_TKEEP_WIDTH-1:0] previous_tkeep;
  local logic previous_tlast;
  local logic[`SVT_AXI_MAX_TID_WIDTH-1:0] previous_tid;
  local logic[`SVT_AXI_MAX_TDEST_WIDTH-1:0] previous_tdest;
  local logic[`SVT_AXI_MAX_TUSER_WIDTH-1:0] previous_tuser;

  `ifdef SVT_AXI_QVN_ENABLE
  /** Variables used in QVN token handshake signal checks */  
  local bit is_varvalidvn_deassertion_check_en [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local bit is_varqosvn_valid_change_check_en  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];

  local bit is_vawvalidvn_deassertion_check_en [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local bit is_vawqosvn_valid_change_check_en  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];

  local bit is_vwvalidvn_deassertion_check_en  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];

  local int unsigned qvn_ar_token_request_ready_timeout_counter_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];
  local int unsigned qvn_aw_token_request_ready_timeout_counter_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];
  local int unsigned qvn_w_token_request_ready_timeout_counter_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];
 
  local logic previous_varvalidvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic [3:0] previous_varqosvnx [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic previous_varreadyvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0]; 
   
  local logic previous_vawvalidvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic [3:0] previous_vawqosvnx [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic previous_vawreadyvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0]; 
  
  local logic previous_vwvalidvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0];
  local logic previous_vwreadyvnx [ `SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0]; 

  `endif

  local svt_axi_snoop_transaction  multipart_dvm_snoop_xact;
  svt_axi_transaction multipart_dvm_coherent_xact;
  local svt_axi_transaction        active_multipart_dvm_coherent_q[svt_axi_transaction];
  local svt_axi_snoop_transaction  active_multipart_dvm_snoop_q[svt_axi_snoop_transaction];

  //local svt_axi_snoop_transaction  multipart_dvm_snoop_check_guard_xact;
  //local svt_axi_master_transaction multipart_dvm_coherent_check_guard_xact;
  local svt_axi_transaction        active_multipart_dvm_coherent_check_guard_q[svt_axi_transaction];
  local svt_axi_snoop_transaction  active_multipart_dvm_snoop_check_guard_q[svt_axi_snoop_transaction];

  /** Enables protocol check coverage provided it protocol_checks_coverage_enable is set
    * in the port configuration as well. If enable_pc_cov is 0, then protocol checks coverage
    * will not be enabled, even if it is set in configuration
    */
  local bit enable_pc_cov = 1;

  /** indicates if only partial ID bits are considered for exclusive transaction */
  local bit partial_exclusive_id = 0;
  

`protected
fJK08B/+AJ<\[_]80X2->6>OD)A2J<>W3ccM5Z^IF4a\BAU?A@?#/)965ggA^&6V
?T&+IRC7QTI\/$
`endprotected



  //--------------------------------------------------------------
  /** Checks that ARID is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arid_when_arvalid_high_check;

  /** Checks that ARADDR is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_araddr_when_arvalid_high_check;

  /** Checks that ARLEN is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arlen_when_arvalid_high_check;
  
  /** Checks that ARSIZE is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arsize_when_arvalid_high_check;
  
  /** Checks that ARLEN and ARSIZE are valid for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_arlen_arsize_check;
  
  /** Checks that ARCACHE is valid for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_arcache_check;
  
  /** Checks that address is aligned for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_read_addr_aligned_check;
  
  /** Checks that AWLEN and AWSIZE are valid for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_awlen_awsize_check;
  
  /** Checks that AWCACHE is valid for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_awcache_check;
  
  /** Checks that address is aligned for exclusive read transaction */
  svt_err_check_stats signal_valid_exclusive_write_addr_aligned_check;

  /** Checks that address is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_addr_check;
  
  /** Checks that received write data is not interleaved beyond write_data_interleave_depth value
    * An error is issued if write data is interleaved beyond this value for Write data interleaving */
  svt_err_check_stats write_data_interleave_depth_check;
 
  /** Checks that the order in which a slave receives the first data item of each transaction must be the
    * same as the order in which it receives the addresses for the transactions for Write Data Interleaving 
    * transactions */
  svt_err_check_stats write_data_interleave_order_check;

 /** Checks that id is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_id_check;

  /** Checks that response generated for exclusive load accesss is correct */
  svt_err_check_stats exclusive_load_response_check;

  /** Checks that response generated for exclusive store accesss is correct */
  svt_err_check_stats exclusive_store_response_check;

  /** Checks that master does not permit an Exclusive Store transaction to be
    * in progress at the same time as any transaction that registers that it
    * is performing an Exclusive sequence
    */
  svt_err_check_stats exclusive_store_overlap_with_another_exclusive_sequence_check;

  /** Checks that, once a master receives successful exclusive store response EXOKAY
    * from interconnect, then no other master should be provided with EXOKAY response,
    * until current master acknowledges completing successful exclusive store by asserting RACK
    */
   svt_err_check_stats exokay_not_sent_until_successful_exclusive_store_rack_observed_check;
  
    /** Checks that READ_ONLY_INTERFACE supports only read transactions 
     * Applicable only for AXI4 VIP
     * Passive Master,Passive Slave and Active slave will perform this
     * check
     */
     svt_err_check_stats read_xact_on_read_only_interface_check;
   
    /** Checks that WRITE_ONLY_INTERFACE supports only write transactions 
     * Applicable only for AXI4 VIP
     * Passive Master,Passive Slave and Active slave will perform this
     * check
     */
     svt_err_check_stats write_xact_on_write_only_interface_check;
     
     /** Checks that READ_ONLY_INTERFACE does not support exclusive access  
     * Applicable only for AXI4 VIP
     * Passive Master,Passive Slave and Active slave will perform this 
     * check
     */
     svt_err_check_stats excl_access_on_read_only_interface_check;

      /** Checks that WRITE_ONLY_INTERFACE does not support exclusive access  
      * Applicable only for AXI4 VIP
      * Passive Master,Passive Slave and Active slave will perform this 
      * check
      */
      svt_err_check_stats excl_access_on_write_only_interface_check;
     
     /** Checks that burst length is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_burst_length_check;
  
  /** Checks that burst size is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_burst_size_check;
  
  /** Checks that burst type is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_burst_type_check;
  
  /** Checks that cache type is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_cache_type_check;
  
  /** Checks that protection type is generated same for exclusive read and write
   * transactions */
  svt_err_check_stats exclusive_read_write_prot_type_check;
  
  /** Checks that exclusive transaction sent on AXI_ACE interface are
   * only of WRITENOSNOOP, READNOSNOOP, READCLEAN, READSHARED and CLEANUNIQUE type */
  svt_err_check_stats exclusive_ace_transaction_type_check;

  /** Checks that ARADDR[2:0] for multipart dvm xact is not other than SBZ */
  svt_err_check_stats signal_araddr_multipart_dvm_xact_check;

  /** Checks that ARBURST is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arburst_when_arvalid_high_check;

  /** Checks that ARLOCK is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arlock_when_arvalid_high_check;

  /** Checks that ARCACHE is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arcache_when_arvalid_high_check;

  /** Checks that ARPROT is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arprot_when_arvalid_high_check;

  /** Checks that ARQOS is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arqos_when_arvalid_high_check;

  /** Checks that ARREGION is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arregion_when_arvalid_high_check;

  /** Checks that ARUSER is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_aruser_when_arvalid_high_check;
  
    /** Checks that ARDOMAIN is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_ardomain_when_arvalid_high_check;
  
  /** Checks that ARSNOOP is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arsnoop_when_arvalid_high_check;
  
  /** Checks that ARBAR is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arbar_when_arvalid_high_check;

  /** Checks that ARREADY is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_arready_when_arvalid_high_check;

  /** Checks that AWDOMAIN is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awdomain_when_awvalid_high_check;
  
  /** Checks that AWSNOOP is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awsnoop_when_awvalid_high_check;
  
  /** Checks that AWBAR is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awbar_when_awvalid_high_check;
  //--------------------------------------------------------------
  /** Checks that ARID is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arid_when_arvalid_high_check;

  /** Checks that ARADDR is stable when ARVALID is high */
  svt_err_check_stats signal_stable_araddr_when_arvalid_high_check;

  /** Checks that RACK is asserted for a single cycle */
  svt_err_check_stats signal_rack_single_cycle_high_check;

  /** Checks that RACK signal must be asserted the cycle after the associated handshake or later */
  svt_err_check_stats signal_rack_after_handshake_check;

  /** Checks that WACK is asserted for a single cycle */
  svt_err_check_stats signal_wack_single_cycle_high_check;

  /** Checks that WACK signal must be asserted the cycle after the associated handshake or later */
  svt_err_check_stats signal_wack_after_handshake_check;

  /** Checks that ARLEN is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arlen_when_arvalid_high_check;
  
  /** Checks that ARSIZE is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arsize_when_arvalid_high_check;

  /** Checks that ARBURST is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arburst_when_arvalid_high_check;

  /** Checks that ARLOCK is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arlock_when_arvalid_high_check;

  /** Checks that ARCACHE is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arcache_when_arvalid_high_check;

  /** Checks that ARPROT is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arprot_when_arvalid_high_check;

  /** Checks that ARQOS is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arqos_when_arvalid_high_check;

  /** Checks that ARREGION is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arregion_when_arvalid_high_check;

  /** Checks that ARUSER is stable when ARVALID is high */
  svt_err_check_stats signal_stable_aruser_when_arvalid_high_check;
  
  /** Checks that ARDOMAIN is stable when ARVALID is high */
  svt_err_check_stats signal_stable_ardomain_when_arvalid_high_check;
  
  /** Checks that ARSNOOP is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arsnoop_when_arvalid_high_check;
  
  /** Checks that ARBAR is stable when ARVALID is high */
  svt_err_check_stats signal_stable_arbar_when_arvalid_high_check;

  /** Checks that AWDOMAIN is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awdomain_when_awvalid_high_check;
  
  /** Checks that AWSNOOP is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awsnoop_when_awvalid_high_check;
  
  /** Checks that AWBAR is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awbar_when_awvalid_high_check;
  //--------------------------------------------------------------
  /** Checks that RID is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rid_when_rvalid_high_check;

  /** Checks that RDATA is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rdata_when_rvalid_high_check;

  /** Checks that RDATACHK is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rdatachk_when_rvalid_high_check;
 
  /** Checks that rpoison is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rpoison_when_rvalid_high_check;
 
  /** Checks that RUSER is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_ruser_when_rvalid_high_check;

  /** Checks that RRESP is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rresp_when_rvalid_high_check;

  /** Checks that RLAST is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rlast_when_rvalid_high_check;

  /** Checks that RREADY is not X or Z when RVALID is high */
  svt_err_check_stats signal_valid_rready_when_rvalid_high_check;

  /** Checks that RID is stable when RVALID is high */
  svt_err_check_stats signal_stable_rid_when_rvalid_high_check;

  /** Checks that RUSER is stable when RVALID is high */
  svt_err_check_stats signal_stable_ruser_when_rvalid_high_check;

  /** Checks that RDATA is stable when RVALID is high */
  svt_err_check_stats signal_stable_rdata_when_rvalid_high_check;

  /** Checks that RRESP is stable when RVALID is high */
  svt_err_check_stats signal_stable_rresp_when_rvalid_high_check;

  /** Checks that RLAST is stable when RVALID is high */
  svt_err_check_stats signal_stable_rlast_when_rvalid_high_check;

  /** Checks that sample read data has associated address */
  svt_err_check_stats read_data_follows_addr_check;
  //--------------------------------------------------------------
  /** Checks that AWID is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awid_when_awvalid_high_check;

  /** Checks that valid write strobes are driven */
  svt_err_check_stats valid_write_strobe_check;

`ifdef SVT_ACE5_ENABLE 
  //--------------------------------------------------------------
 /** Checks that stash_nid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_stash_nid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that stash_lpid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_stash_lpid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that stash_nid_valid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_stash_nid_valid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that stash_lpid_valid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_stash_lpid_valid_when_awvalid_high_check;

  //--------------------------------------------------------------
 /** Checks that awmmusid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmusid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that awmmussid is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmussid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that  is awmmusecsid not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmusecsid_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that awmmussidv is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmussidv_when_awvalid_high_check;

 //--------------------------------------------------------------
/** Checks that awmmuatst is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmmuatst_when_awvalid_high_check;

  //--------------------------------------------------------------
 /** Checks that armmusid is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmusid_when_arvalid_high_check;

 //--------------------------------------------------------------
/** Checks that armmussid is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmussid_when_arvalid_high_check;

 //--------------------------------------------------------------
/** Checks that  is armmusecsid not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmusecsid_when_arvalid_high_check;

 //--------------------------------------------------------------
/** Checks that armmussidv is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmussidv_when_arvalid_high_check;

 //--------------------------------------------------------------
/** Checks that armmuatst is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armmuatst_when_arvalid_high_check;

 /** Checks that awatop is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awatop_when_awvalid_high_check;

 /** Checks that armpam is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_armpam_when_arvalid_high_check;

 /** Checks that awmpam is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awmpam_when_awvalid_high_check;

   /** Checks that AWMPAM is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awmpam_when_awvalid_high_check;

  /** Checks that ARMPAM is stable when ARVALID is high */
  svt_err_check_stats signal_stable_armpam_when_arvalid_high_check;
`endif

`ifdef SVT_ACE5_ENABLE 
//--------------------------------------------------------------
 /** Checks that ARIDUNQ is not X or Z when ARVALID is high*/
   svt_err_check_stats signal_valid_aridunq_when_arvalid_high_check;

 /** Checks that RIDUNQ is not X or Z when RVALID is high*/
   svt_err_check_stats signal_valid_ridunq_when_rvalid_high_check;

 /** Checks that AWIDUNQ is not X or Z when AWVALID is high*/
   svt_err_check_stats signal_valid_awidunq_when_awvalid_high_check;

 /** Checks that BIDUNQ is not X or Z when BVALID is high*/
   svt_err_check_stats signal_valid_bidunq_when_bvalid_high_check;
   
//--------------------------------------------------------------
/** Checks that ARIDUNQ is stable when ARVALID is high */
  svt_err_check_stats signal_stable_aridunq_when_arvalid_high_check;

/** Checks that RIDUNQ is stable when RVALID is high */
  svt_err_check_stats signal_stable_ridunq_when_rvalid_high_check;

/** Checks that AWIDUNQ is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awidunq_when_awvalid_high_check;

/** Checks that BIDUNQ is stable when BVALID is high */
  svt_err_check_stats signal_stable_bidunq_when_bvalid_high_check;

//--------------------------------------------------------------
  /** Checks that RIDUNQ asserted or deasserted when ARIDUNQ asserted or deasserted */
  //svt_err_check_stats ridunq_asserted_deasserted_check;

  /** Checks that BIDUNQ asserted or deasserted when AWIDUNQ asserted or deasserted*/
  //svt_err_check_stats bidunq_asserted_deasserted_check;
 
  /** Checks that there is no outstanding transaction with same arid */
  svt_err_check_stats no_outstanding_read_unique_transaction_with_same_arid;

  /** Checks that there is no outstanding transaction with same awid */
  svt_err_check_stats no_outstanding_write_unique_transaction_with_same_awid;
`endif

  /** Checks that AWADDR is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awaddr_when_awvalid_high_check;

  /** Checks that AWLEN is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awlen_when_awvalid_high_check;
  
  /** Checks that AWSIZE is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awsize_when_awvalid_high_check;

  /** Checks that AWBURST is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awburst_when_awvalid_high_check;

  /** Checks that AWLOCK is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awlock_when_awvalid_high_check;

  /** Checks that AWCACHE is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awcache_when_awvalid_high_check;

  /** Checks that AWPROT is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awprot_when_awvalid_high_check;

  /** Checks that AWREADY is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awready_when_awvalid_high_check;

  /** Checks that AWQOS is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awqos_when_awvalid_high_check;

  /** Checks that AWREGION is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awregion_when_awvalid_high_check;

  /** Checks that AWUNIQUE is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awunique_when_awvalid_high_check;

  /** Checks that AWUSER is not X or Z when AWVALID is high */
  svt_err_check_stats signal_valid_awuser_when_awvalid_high_check;
  //--------------------------------------------------------------
  /** Checks that AWID is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awid_when_awvalid_high_check;

  /** Checks that AWADDR is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awaddr_when_awvalid_high_check;

  /** Checks that AWLEN is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awlen_when_awvalid_high_check;
  
  /** Checks that AWSIZE is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awsize_when_awvalid_high_check;

  /** Checks that AWBURST is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awburst_when_awvalid_high_check;

  /** Checks that AWLOCK is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awlock_when_awvalid_high_check;

  /** Checks that AWCACHE is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awcache_when_awvalid_high_check;

  /** Checks that AWPROT is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awprot_when_awvalid_high_check;

  /** Checks that AWQOS is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awqos_when_awvalid_high_check;

  /** Checks that AWREGION is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awregion_when_awvalid_high_check;

  /** Checks that AWUNIQUE is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awunique_when_awvalid_high_check;

  /** Checks that AWUSER is stable when AWVALID is high */
  svt_err_check_stats signal_stable_awuser_when_awvalid_high_check;

  //--------------------------------------------------------------

  /** Checks that WID is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wid_when_wvalid_high_check;

  /** Checks that WUSER is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wuser_when_wvalid_high_check;

  /** Checks that WDATA is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wdata_when_wvalid_high_check;

  /** Checks that WDATACHK is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wdatachk_when_wvalid_high_check;

 /** Checks that WPOISON is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wpoison_when_wvalid_high_check;

  /** Checks that WSTRB is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wstrb_when_wvalid_high_check;

  /** Checks that WLAST is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wlast_when_wvalid_high_check;

  /** Checks that WREADY is not X or Z when WVALID is high */
  svt_err_check_stats signal_valid_wready_when_wvalid_high_check;

  /** Checks that WID is stable when WVALID is high */
  svt_err_check_stats signal_stable_wid_when_wvalid_high_check;

  /** Checks that WUSER is stable when WVALID is high */
  svt_err_check_stats signal_stable_wuser_when_wvalid_high_check;

  /** 
   * Checks that WDATA is stable when WVALID is high 
   * When svt_axi_port_configuration::check_valid_data_bytes_only_enable=1 ,
   * it considers only valid byte lanes of wdata based on wstrb. 
   * When svt_axi_port_configuration::check_valid_data_bytes_only_enable=0 ,
   * whole wdata as seen on the bus will be considered.
   */
  svt_err_check_stats signal_stable_wdata_when_wvalid_high_check;

  /** Checks that WSTRB is stable when WVALID is high */
  svt_err_check_stats signal_stable_wstrb_when_wvalid_high_check;

  /** Checks that WLAST is stable when WVALID is high */
  svt_err_check_stats signal_stable_wlast_when_wvalid_high_check;

  //--------------------------------------------------------------
  /** Checks that BID is not X or Z when BVALID is high */
  svt_err_check_stats signal_valid_bid_when_bvalid_high_check;

  /** Checks that BUSER is not X or Z when BVALID is high */
  svt_err_check_stats signal_valid_buser_when_bvalid_high_check;

  /** Checks that BRESP is not X or Z when BVALID is high */
  svt_err_check_stats signal_valid_bresp_when_bvalid_high_check;

  /** Checks that BREADY is not X or Z when BVALID is high */
  svt_err_check_stats signal_valid_bready_when_bvalid_high_check;

  /** Checks that BID is stable when BVALID is high */
  svt_err_check_stats signal_stable_bid_when_bvalid_high_check;

  /** Checks that BUSER is stable when BVALID is high */
  svt_err_check_stats signal_stable_buser_when_bvalid_high_check;

  /** Checks that BRESP is stable when BVALID is high */
  svt_err_check_stats signal_stable_bresp_when_bvalid_high_check;

  /** 
    * When a write response is sampled, checks that there is a 
    * transaction with corresponding ID whose data phase is complete 
    */
  svt_err_check_stats write_resp_follows_last_write_xfer_check;

  /** 
    * Checks that WLAST is asserted for the last beat of write data. 
    */
  svt_err_check_stats wlast_asserted_for_last_write_data_beat;

  //--------------------------------------------------------------
  // Checks that need to be executed externally (by monitor).
  /** Checks that ARVALID is not X or Z */
  svt_err_check_stats signal_valid_arvalid_check;

  /** Checks that RVALID is not X or Z */
  svt_err_check_stats signal_valid_rvalid_check;

  /** Checks that AWVALID is not X or Z */
  svt_err_check_stats signal_valid_awvalid_check;

  /** Checks that WVALID is not X or Z */
  svt_err_check_stats signal_valid_wvalid_check;

  /** Checks that BVALID is not X or Z */
  svt_err_check_stats signal_valid_bvalid_check;
  
  /** Checks that ACVALID is not X or Z */
  svt_err_check_stats signal_valid_acvalid_check;
  
  /** Checks that CDVALID is not X or Z */
  svt_err_check_stats signal_valid_cdvalid_check;
  
  /** Checks that CDVALID is not X or Z */
  svt_err_check_stats signal_valid_crvalid_check;

  /** Checks that ARVALID is not X or Z During Reset */
  svt_err_check_stats signal_valid_arvalid_check_during_reset;

  /** Checks that RVALID is not X or Z During Reset*/
  svt_err_check_stats signal_valid_rvalid_check_during_reset;

  /** Checks that AWVALID is not X or Z During Reset*/
  svt_err_check_stats signal_valid_awvalid_check_during_reset;

  /** Checks that WVALID is not X or Z During Reset*/
  svt_err_check_stats signal_valid_wvalid_check_during_reset;

  /** Checks that BVALID is not X or Z During Reset */
  svt_err_check_stats signal_valid_bvalid_check_during_reset;

  /** Checks if arvalid was interrupted before arready got asserted */
  svt_err_check_stats arvalid_interrupted_check;
  
  /** Checks if acvalid was interrupted before acready got asserted */
  svt_err_check_stats acvalid_interrupted_check;
  
  /** Checks if cdvalid was interrupted before cdrready got asserted */
  svt_err_check_stats cdvalid_interrupted_check;
  
  /** Checks if crvalid was interrupted before crready got asserted */
  svt_err_check_stats crvalid_interrupted_check;

  /** Checks if rvalid was interrupted before rready got asserted */
  svt_err_check_stats rvalid_interrupted_check;

  /** Checks if awvalid was interrupted before awready got asserted */
  svt_err_check_stats awvalid_interrupted_check;

  /** Checks if wvalid was interrupted before wready got asserted */
  svt_err_check_stats wvalid_interrupted_check;

  /** Checks if bvalid was interrupted before bready got asserted */
  svt_err_check_stats bvalid_interrupted_check;
  //--------------------------------------------------------------
  /** Checks if rvalid is low when reset is active */
  svt_err_check_stats rvalid_low_when_reset_is_active_check;

  /** Checks if bvalid is low when reset is active */
  svt_err_check_stats bvalid_low_when_reset_is_active_check;

  /** Checks if arvalid is low when reset is active */
  svt_err_check_stats arvalid_low_when_reset_is_active_check;

  /** Checks if acvalid is low when reset is active */
  svt_err_check_stats acvalid_low_when_reset_is_active_check;
  
  /** Checks if crvalid is low when reset is active */
  svt_err_check_stats crvalid_low_when_reset_is_active_check;
  
  /** Checks if cdvalid is low when reset is active */
  svt_err_check_stats cdvalid_low_when_reset_is_active_check;

  /** Checks if awvalid is low when reset is active */
  svt_err_check_stats awvalid_low_when_reset_is_active_check;

  /** Checks if wvalid is low when reset is active */
  svt_err_check_stats wvalid_low_when_reset_is_active_check;
  //--------------------------------------------------------------
  
  /** Checks if write burst cross a 4KB boundary */
  svt_err_check_stats awaddr_4k_boundary_cross_active_check;
  //--------------------------------------------------------------

  /** Checks if write burst of WRAP type has an aligned address*/
  svt_err_check_stats awaddr_wrap_aligned_active_check ;
  //--------------------------------------------------------------
  
  /** Checks if write burst of WRAP type has a valid length*/
  svt_err_check_stats awlen_wrap_active_check;
  //--------------------------------------------------------------

  /** Checks if size of write transfer exceeds the width of the data bus*/
  svt_err_check_stats awsize_data_width_active_check;
  //--------------------------------------------------------------
        
  /** Checks if the value of awburst=2'b11 when awvalid is high*/
  svt_err_check_stats awburst_reserved_val_check;
  //--------------------------------------------------------------
  
  /** Checks if the value of awcache[3:2]=2'b00 when awvalid is high and awcache[1] is also low*/
  svt_err_check_stats awvalid_awcache_active_check;
  //--------------------------------------------------------------

  
  /** Checks if read burst cross a 4KB boundary */
  svt_err_check_stats araddr_4k_boundary_cross_active_check;
  //--------------------------------------------------------------

  /** Checks if read  burst of WRAP type has an aligned address*/
  svt_err_check_stats araddr_wrap_aligned_active_check ;
  //--------------------------------------------------------------

  /** Checks if snoop address is aligned with snoop data width */
  svt_err_check_stats acaddr_aligned_to_cddata_width_valid_check ;
  //--------------------------------------------------------------

  /** Checks that a cached master does not initiate WriteUnique or WriteLineUnique
    * coherent write transaction while any WriteBack, WriteClean or WriteEvict transaction
    * is outstanding.
    */
  svt_err_check_stats complete_outstanding_memory_write_before_writeunique_writelineunique_check ;

  /** Checks that a cached master does not issue WriteBack, WriteClean or WriteEvict
    * transaction while any WriteUnique or WriteLineUnique coherent write transaction
    * is in progress.
    * It automatically checks second rule which says, Complete any incoming snoop 
    * transactions without the use of WriteBack, WriteClean, or WriteEvict
    * transactions while a WriteUnique or WriteLineUnique transaction is in progress.
    */
  svt_err_check_stats complete_outstanding_writeunique_writelineunique_before_memory_write_check ;


  /** Checks that CleanInvalid and MakeInvalid cache maintenance transactions are not 
    * initiated while any memory update or shareable transactions are outstanding. It
    * also checks that CleanShared cache maintenance transactions are not initiated 
    * while any memory update or any shareable transactions that can make the cacheline
    * dirty, are outstanding.
    */
  svt_err_check_stats cache_maintenance_outstanding_transaction_check ;

  /** Checks that WriteBack, WriteClean or any shareable transactions are not issued 
    * while cache maintenance transaction is in progress.
    */
  svt_err_check_stats no_memory_update_or_shareable_txn_during_cache_maintenance_check ;

  /** Monitor checks that when master initiates a CleanShared cache maintenance transaction, 
    * and receives any snoop transaction to the same cacheline, the initiating master must not
    * assert PassDirty snoop response. It also checks that when master initiates CleanInvalid
    * or MakeInvalid cache maintenance transactions, and receives any snoop transaction to the
    * same cacheline, the initiating master must not assert PassDirty, IsShared and DataTransfer
    * snoop responses.
    */
  svt_err_check_stats valid_snoop_response_during_cache_maintenance_check ;
  //--------------------------------------------------------------

  /** Checks if number of databeat transferred over snoop data channel is valid */
  svt_err_check_stats snoop_transaction_burst_length_check ;
  //--------------------------------------------------------------
  
  /** Checks if read burst of WRAP type has a valid length*/
  svt_err_check_stats arlen_wrap_active_check;
  //--------------------------------------------------------------

  /** Checks if size of read transfer exceeds the width of the data bus*/
  svt_err_check_stats arsize_data_width_active_check;
  //--------------------------------------------------------------
        
  /** Checks if the value of arburst=2'b11 when arvalid is high*/
  svt_err_check_stats arburst_reserved_val_check;
  //--------------------------------------------------------------
  
  /** Checks if the value of arcache[3:2]=2'b00 when arvalid is high and arcache[1] is also low*/
  svt_err_check_stats arvalid_arcache_active_check;
  //--------------------------------------------------------------
  
/** Checks if the number of write data items matches AWLEN for the corresponding address */
  svt_err_check_stats wdata_awlen_match_for_corresponding_awaddr_check;
  //--------------------------------------------------------------

/** Checks if the slave must only give a write response after the last write data item is transferred  */
  svt_err_check_stats write_resp_after_last_wdata_check;
  //--------------------------------------------------------------

/** Checks if  A slave must not give a write response before the write address */
  svt_err_check_stats write_resp_after_write_addr_check;
  //--------------------------------------------------------------

/** Checks if the number of read data items matches ARLEN for the corresponding address */
  svt_err_check_stats rdata_arlen_match_for_corresponding_araddr_check;
  //--------------------------------------------------------------

/** Checks if the number of read data items matches ARLEN for the corresponding address */
 svt_err_check_stats rlast_asserted_for_last_read_data_beat;
//ACE CHECKS//

  /** Checks that ACREADY is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_acready_when_arvalid_high_check;
  
  /** Checks that ACADDR is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_acaddr_when_acvalid_high_check;
  
  /** Checks that ACSNOOP is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_acsnoop_when_acvalid_high_check;
  
  /** Checks that ACPROT is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_acprot_when_acvalid_high_check;
  
  /** Checks that CDREADY is not X or Z when CDVALID is high */
  svt_err_check_stats signal_valid_cdready_when_cdvalid_high_check;
  
  /** Checks that CDDATA is not X or Z when CDVALID is high */
  svt_err_check_stats signal_valid_cddata_when_cdvalid_high_check;
  
  /** Checks that CDDATACHK is not X or Z when CDVALID is high */
  svt_err_check_stats signal_valid_cddatachk_when_cdvalid_high_check;
  
  /** Checks that CDPOISON is not X or Z when CDVALID is high */
  svt_err_check_stats signal_valid_cdpoison_when_cdvalid_high_check;

 /** Checks that ACREADY is not X or Z when ARVALID is high */
  svt_err_check_stats signal_valid_cdlast_when_cdvalid_high_check;
  
  /** Checks that CRREADY is not X or Z when CRVALID is high */
  svt_err_check_stats signal_valid_crready_when_crvalid_high_check;
  
  /** Checks that CRRESP is not X or Z when CRVALID is high */
  svt_err_check_stats signal_valid_crresp_when_crvalid_high_check;

  /** Checks that ACADDR is stable when ARVALID is high */
  svt_err_check_stats signal_stable_acaddr_when_acvalid_high_check;
  
  /** Checks that ACSNOOP is stable when ARVALID is high */
  svt_err_check_stats signal_stable_acsnoop_when_acvalid_high_check;
  
  /** Checks that ACPROT is stable when ARVALID is high */
  svt_err_check_stats signal_stable_acprot_when_acvalid_high_check;

  /** Checks that CDDATA is stable when CDVALID is high */
  svt_err_check_stats signal_stable_cddata_when_cdvalid_high_check;
  
  /** Checks that ACREADY is stable when ARVALID is high */
  svt_err_check_stats signal_stable_cdlast_when_cdvalid_high_check;

  /** Checks that CRRESP is stable when CRVALID is high */
  svt_err_check_stats signal_stable_crresp_when_crvalid_high_check;
  
  
/**Checks if the Device transactions, as indicated by AxCACHE[1] = 0, must only use AxDOMAIN = 11.  */
 svt_err_check_stats axcache_axdomain_restriction_check;
  //--------------------------------------------------------------

/**Checks if the  AXCACHE and AXDOMAIN value are valid */
 svt_err_check_stats axcache_axdomain_invalid_value_check ;
  //--------------------------------------------------------------



/**Checks if the  AWSIZE is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_awsize_valid_value_check;
  //--------------------------------------------------------------
/**Checks if the  ARSIZE is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_arsize_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWLEN is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_awlen_valid_value_check;
  //--------------------------------------------------------------
/**Checks if the  ARLEN is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_arlen_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWSIZE is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_awsize_valid_check;
  //--------------------------------------------------------------

/**Checks if the  AWBURST is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_awburst_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  ARBURST is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_arburst_valid_value_check;
  //--------------------------------------------------------------

 /**Checks if the  ARSIZE is valid for Cache Line Size Transactions */
 svt_err_check_stats cache_line_arsize_valid_check;
  //--------------------------------------------------------------

/**Checks if the  address is aligned for AWBURST in  Cache Line Size Transactions */
 svt_err_check_stats cache_line_awburst_wrap_addr_aligned_valid_check;
  //--------------------------------------------------------------
/**Checks if the  address is aligned for ARBURST in  Cache Line Size Transactions */
 svt_err_check_stats cache_line_arburst_wrap_addr_aligned_valid_check;
  //--------------------------------------------------------------
/**Checks if the  address is aligned for AWBURST in  Cache Line Size Transactions */
 svt_err_check_stats cache_line_awburst_incr_addr_aligned_valid_check;
  //--------------------------------------------------------------
/**Checks if the  address is aligned for ARBURST in  Cache Line Size Transactions */
 svt_err_check_stats cache_line_arburst_incr_addr_aligned_valid_check;
  //--------------------------------------------------------------

/**Checks if the  AWDOMAIN is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_awdomain_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  ARDOMAIN is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_ardomain_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWCACHE is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_awcache_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  AWLOCK is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_awlock_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  ARLOCK is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_arlock_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWCACHE is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_arcache_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  AxBAR is valid for Cache Line Size Transactions */
 svt_err_check_stats  cache_line_axbar_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  AxLEN is correctly indicated as per the Cache Line Size configured */
 svt_err_check_stats  cache_line_sz_eq_alen_asize_check ;
  //--------------------------------------------------------------

  /**Checks if CLEANSHARED transaction starts only from INVALID, UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats cleanshared_correct_start_state_check; 
  //--------------------------------------------------------------

  /**Checks if CLEANSHAREDPERSIST transaction starts only from INVALID, UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats cleansharedpersist_correct_start_state_check; 
  //--------------------------------------------------------------

  /**Checks if CLEANINVALID transaction starts only from INVALID state */
  svt_err_check_stats cleaninvalid_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if MAKEINVALID transaction starts only from INVALID state */
  svt_err_check_stats makeinvalid_correct_start_state_check; 
  //--------------------------------------------------------------

  /**Checks if WRITEUNIQUE transaction starts only from INVALID, UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats writeunique_correct_start_state_check; 
  //--------------------------------------------------------------

  /**Checks if WRITELINEUNIQUE transaction starts only from INVALID, UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats writelineunique_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if WRITEBACK transaction starts only from UNIQUEDIRTY or SHAREDDIRTY state */
  svt_err_check_stats writeback_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if WRITECLEAN transaction starts only from UNIQUEDIRTY or SHAREDDIRTY state */
  svt_err_check_stats writeclean_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if WRITEEVICT transaction starts only from UNIQUECLEAN state */
  svt_err_check_stats writeevict_correct_start_state_check;
  //--------------------------------------------------------------

  /**Checks if EVICT transaction starts only from UNIQUECLEAN or SHAREDCLEAN state */
  svt_err_check_stats evict_correct_start_state_check;         
  //--------------------------------------------------------------

  /**Checks if snoop response has data transfer bit set for cacheline in dirty state */
  svt_err_check_stats dirty_state_data_transfer_check;         
  //--------------------------------------------------------------

/**Checks if the  AWDOMAIN is valid for ReadOnce & WriteUnique Transactions */
 svt_err_check_stats  writeunique_awdomain_valid_value_check;
//------------------------------------------------------------------------

/**Checks if the  AWDOMAIN is valid for WriteUniquePtlstash Transactions */
 svt_err_check_stats  writeuniqueptlstash_awdomain_valid_value_check;

  //--------------------------------------------------------------
/**Checks if the  AWDOMAIN is valid for ReadOnce & WriteUnique Transactions */
 svt_err_check_stats  readonce_ardomain_valid_value_check;
  //--------------------------------------------------------------

 /**Checks if all transactions (other than ReadNoSnoop, ReadOnce, ReadOnceCleanInvalid, ReadOnceMakeInvalid, WriteNoSnoop, WriteUnique) are required to be a full cache line size */
 svt_err_check_stats  full_cache_line_size_check;

/**Checks if the  AWBURST is valid for ReadOnce & WriteUnique Transactions */
 svt_err_check_stats writeunique_awburst_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWBURST is valid for writeuniqueptlstash Transactions */
 svt_err_check_stats writeuniqueptlstash_awburst_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  ARBURST is valid for ReadOnce & WriteUnique  Transactions */
 svt_err_check_stats readonce_arburst_valid_value_check;


/**Checks if the  AWCACHE is valid for ReadOnce & WriteUnique  Transactions */
 svt_err_check_stats  writeunique_awcache_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWLOCK is valid for ReadOnce & WriteUnique  Transactions */
 svt_err_check_stats  writeunique_awlock_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWCACHE is valid for writeuniqueptlstash  Transactions */
 svt_err_check_stats  writeuniqueptlstash_awcache_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWLOCK is valid for writeuniqueptlstash  Transactions */
 svt_err_check_stats  writeuniqueptlstash_awlock_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  ARCACHE is valid for ReadOnce & WriteUnique   Transactions */
 svt_err_check_stats  readonce_arcache_valid_value_check ;
  //--------------------------------------------------------------

 /**Checks if the  ARLOCK is valid for ReadOnce & WriteUnique   Transactions */
 svt_err_check_stats  readonce_arlock_valid_value_check ;
  //--------------------------------------------------------------

/**Checks if the  AWSIZE is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awsize_valid_value_check;
  //--------------------------------------------------------------


/**Checks if the  AWSIZE is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awlen_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWLEN for INCR is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awburst_awlen_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWLEN for INCR is valid for AXI Transactions */
 svt_err_check_stats awburst_awlen_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWBURST is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awburst_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWDOMAIN is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awdomain_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  AWCACHE is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awcache_valid_value_check;
  //--------------------------------------------------------------

/**Checks if the  Address aligned for WRAP is valid for  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awburst_incr_valid_check;
  //--------------------------------------------------------------

/**Checks if the AWSIZE x AWLEN  not exceed the cache line size  WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awburst_wrap_valid_check;
//--------------------------------------------------------------

/**Checks if the ALOCK is 0 for WriteBack and WriteClean Transactions */
 svt_err_check_stats writeback_writeclean_awlock_valid_value_check;
//--------------------------------------------------------------
/** If a snooped master receives a snoop transaction when it is has an
 * outstanding WriteEvict transaction, then it is the responsibility of the
 * snooped master to ensure that no other master can update the same area of
 * main memory at the same time. The snooped master achieves this by delaying
 * the snoop response until the snooped master has completed the WriteEvict
 * transaction */
 svt_err_check_stats snoop_response_to_same_cacheline_during_writeevict_check;
//--------------------------------------------------------------
/** While a transaction is in progress which has the AWUNIQUE signal asserted,
 * the master must not give a snoop response that would allow another copy of
 * the line to be created, or an agent to consider that it has another Unique
 * copy of the line
 */
 svt_err_check_stats snoop_response_to_same_cacheline_during_xact_with_awunique_check;
//--------------------------------------------------------------
/** AWUNIQUE must be deasserted for WRITECLEAN transactions */
svt_err_check_stats writeclean_awunique_valid_value_check;
//--------------------------------------------------------------
/** AWUNIQUE must be asserted for WRITEEVICT transactions */
svt_err_check_stats writeevict_awunique_valid_value_check;
//--------------------------------------------------------------
/** Monitor check that all byte strobes are asserted for a WRITEEVICT transaction */
svt_err_check_stats writeevict_wstrb_valid_value_check;

//--------------------------------------------------------------
/** Monitor check that all byte strobes are asserted for a WRITELINEUNIQUE transaction */
svt_err_check_stats writelineunique_wstrb_valid_value_check;
//--------------------------------------------------------------

/** Monitor check that all byte strobes are asserted for a writeuniquefullstash transaction */
svt_err_check_stats writeuniquefullstash_wstrb_valid_value_check;
//--------------------------------------------------------------

//--------------------------------------------------------------
/**Checks the valid response of EXOKAY response is only for readnosnoop Transactions */
svt_err_check_stats exokay_resp_observed_only_for_exclusive_transactions_check;
//--------------------------------------------------------------
/**Checks that if cacheline is in invalid state then exclusive load transaction is issued only as READCLEAN or READSHARED */
svt_err_check_stats exclusive_load_from_valid_state_check;
//--------------------------------------------------------------
/**Checks that if cacheline is in invalid state then exclusive store transaction is not issued */
svt_err_check_stats exclusive_store_from_valid_state_check;
//--------------------------------------------------------------
/**Checks that if cacheline is in shared state then exclusive transaction is issued only as CLEANUNIQUE, READCLEAN or READSHARED*/
svt_err_check_stats exclusive_transaction_from_shared_state_check;
//--------------------------------------------------------------
/**Checks for no data transfer occurs for a CleanShared,Cleansharedpersist, CleanInvalid, CleanUnique, MakeUnique, MakeInvalid and Evict Transactions */
svt_err_check_stats perform_no_datatransfer_check;
  //--------------------------------------------------------------
/**Checks the valid response of  cleanshared Transactions */
svt_err_check_stats read_data_chan_cleanshared_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  cleansharedPersist Transactions */
svt_err_check_stats read_data_chan_cleansharedpersist_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of makeinvalid  Transactions */
svt_err_check_stats read_data_chan_makeinvalid_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  makeunique Transactions */
svt_err_check_stats read_data_chan_makeunique_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of cleaninvalid  Transactions */
svt_err_check_stats read_data_chan_cleaninvalid_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  cleanunique Transactions */
svt_err_check_stats read_data_chan_cleanunique_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  readunique Transactions */
svt_err_check_stats read_data_chan_readunique_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  readnotshareddirty Transactions */
svt_err_check_stats read_data_chan_readnotshareddirty_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of  readclean Transactions */
svt_err_check_stats read_data_chan_readclean_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of readonce  Transactions */
svt_err_check_stats read_data_chan_readonce_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the valid response of readnosnoop  Transactions */
svt_err_check_stats read_data_chan_readnosnoop_resp_valid_check;
  //--------------------------------------------------------------
/**Checks the CLEANUNIQUE, MAKEUNIQUE, CLEANSHARED,
  * CLEANINVALID,CLEANSHAREDPERSIST,
  * MAKEINVALID, READBARRIER, DVMCOMPLETE, DVMMESSAGE transactions
  * have only single read data channel transfer */
svt_err_check_stats coherent_single_read_data_transfer_valid_check;
  //--------------------------------------------------------------

/**Checks the valid response of readbarrier  Transactions */
svt_err_check_stats read_data_chan_readbarrier_resp_valid_check;
  //--------------------------------------------------------------

/**Checks the valid response of DVM Message Transactions */
svt_err_check_stats read_data_chan_dvmmessage_resp_valid_check;
  //--------------------------------------------------------------

/**Checks the valid response of DVM Complete Transactions */
svt_err_check_stats read_data_chan_dvmcomplete_resp_valid_check;

//--------------------------------------------------------------
/**Checks the valid snoop response of DVM Message Transactions */
svt_err_check_stats snoop_chan_dvmsync_resp_valid_check;
  //--------------------------------------------------------------

/**Checks the valid snoop response of DVM Complete Transactions */
svt_err_check_stats snoop_chan_dvmcomplete_resp_valid_check;

//--------------------------------------------------------------
/**Checks the ACSNOOP reserved values */
svt_err_check_stats acsnoop_reserved_value_check ;
 //--------------------------------------------------------------


/**Checks that for MakeInvalid transactions a data transfer is never required */
svt_err_check_stats snoop_resp_passdirty_datatransfer_check;
//--------------------------------------------------------------

/**If DataTransfer is asserted, a full cache line of data must be provided on the snoop data channel */
svt_err_check_stats full_cache_line_datatransfer_check;
//

/**Checks for readunique cleaninvalid makeinvalid illegal response  */
svt_err_check_stats snoop_response_channel_isshared_check;
//--------------------------------------------------------------

/** Checks that CDLAST signal is asserted during the final data transfer.
  *
  * protocol checks : port level 
  */
svt_err_check_stats cdlast_asserted_for_last_snoopread_data_beat;
//--------------------------------------------------------------

/**Checks that the FIXED burst type is not supported for shareable transactions */
svt_err_check_stats fixed_burst_type_valid;
//--------------------------------------------------------------

/**Checks that ACVALID and ACREADY to be asserted before asserting CRVALID */
svt_err_check_stats snoop_addr_snoop_resp_check;
//--------------------------------------------------------------
/**Checks that ACVALID and ACREADY to be asserted before asserting CDVALID */
svt_err_check_stats snoop_addr_snoop_data_check;
//--------------------------------------------------------------

//--------------------------------------------------------------
/**Checks the combinations of ARDOMAIN,ARSNOOP and ARBAR are valid and unreserved */
svt_err_check_stats arsnoop_ardomain_arbar_reserve_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWDOMAIN,AWSNOOP and AWBAR are valid and unreserved */
svt_err_check_stats awsnoop_awdomain_awbar_reserve_value_check;
//--------------------------------------------------------------

//Barrier Checks //
/**Checks the AWADDR is valid for AWBAR  */
svt_err_check_stats write_barrier_awaddr_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations AWBURST and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awburst_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWLEN and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awlen_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWSIZE and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awsize_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWCACHE and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awcache_type_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWSNOOP and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awsnoop_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of AWLOCK and AWBAR are valid and unreserved */
svt_err_check_stats write_barrier_awlock_type_valid_value_check;
//--------------------------------------------------------------
/**Checks the valid value of AxUSER for write barrier transactions */
svt_err_check_stats barrier_transaction_user_valid_value_check;
//--------------------------------------------------------------

/**Checks the ARADDR is valid for ARBAR  */
svt_err_check_stats read_barrier_araddr_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations ARBURST and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arburst_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARLEN and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arlen_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARSIZE and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arsize_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARCACHE and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arcache_type_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARSNOOP and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arsnoop_valid_value_check;
//--------------------------------------------------------------
/**Checks the combinations of ARLOCK and ARBAR are valid and unreserved */
svt_err_check_stats read_barrier_arlock_type_valid_value_check;
//--------------------------------------------------------------
/** Checks the Barrier Id valid and unreserved.  */
svt_err_check_stats barrier_id_valid_value_check;
//--------------------------------------------------------------
/**Checks the Read Barrier valid response  */
svt_err_check_stats barrier_read_response_check ;
//--------------------------------------------------------------
/**Checks the Write Barrier valid response  */
svt_err_check_stats barrier_write_response_check ;
//--------------------------------------------------------------
/**Checks that both transactions in a barrier pair must have the same AxID, AxBAR, AxDOMAIN, and AxPROT values*/
svt_err_check_stats barrier_pair_cntrl_signals_check ;
//--------------------------------------------------------------
/**Checks that barrier pairs must be issued in the same sequence on the read address and write address channels*/
svt_err_check_stats barrier_pair_check ;
//--------------------------------------------------------------
/**Checks that ARADDR/AWADDR should always be aligned to Atomicity Size*/
svt_err_check_stats align_addr_atomicity_size_check ;

//--------------------------------------------------------------
/** Checks the RACK for valid response.  */
svt_err_check_stats rack_status_check;
//--------------------------------------------------------------
/** Checks the WACK for valid response.  */
svt_err_check_stats wack_status_check;
//-------------------------------------------------------------
/** Checks all snoop transactions are ordered. .
  */
svt_err_check_stats snoop_transaction_order_check;

//DVM CHECKS //
 /**Checks  For DVM ARBURST 'b01 Burst Type INCR. */
svt_err_check_stats dvm_message_arburst_valid_value_check;
//-------------------------------------------------------------
 /**Checks For DVM  ARLEN All zero */
svt_err_check_stats dvm_message_arlen_valid_value_check;
//-------------------------------------------------------------

 /**Checks for DVM ARSIZE Matches the data bus width */
svt_err_check_stats dvm_message_arsize_valid_value_check;
//-------------------------------------------------------------

 /**Checks for DVM ARCACHE 'b0010 Normal non-cacheable */
svt_err_check_stats dvm_message_arcache_type_valid_value_check;
//-------------------------------------------------------------

 /**Checks for DVM ARLOCK 'b0 Normal Access. */
svt_err_check_stats dvm_message_arlock_type_valid_value_check;
//-------------------------------------------------------------
 
/**Checks for DVM  ARDOMAIN  is Inner shareable or Outer shareable */ 
svt_err_check_stats dvm_message_ardomain_type_valid_value_check;
//-------------------------------------------------------------
/**Checks for DVM  ARBAR[0] is 1'b0 */ 
svt_err_check_stats dvm_message_arbar_valid_value_check;
//-------------------------------------------------------------
/** Checks for DVMCOMPLETE the valid value of  ARSNOOP */ 
svt_err_check_stats dvm_complete_arsnoop_valid_value_check;
//-------------------------------------------------------------
/** Checks for DVMSYNC, DVM Operation the valid value of  ARSNOOP */ 
svt_err_check_stats dvm_operation_dvm_sync_arsnoop_valid_value_check;
//-------------------------------------------------------------
/** Checks for DVMSYNC, DVM Operation the valid value of ARADDR[(n-1):32],[15],[11:0] bits */
svt_err_check_stats dvm_operation_dvm_sync_araddr_valid_value_check;
//-------------------------------------------------------------
/** Checks for DVMHINT, DVM Operation the valid value of ARADDR[15] */
svt_err_check_stats dvm_operation_dvm_hint_araddr_valid_value_check;
//-------------------------------------------------------------

/** Checks the value of  ACSNOOP for the DVM complete */ 
svt_err_check_stats dvm_complete_acsnoop_valid_value_check;
//-------------------------------------------------------------
/** Checks the value of  ACSNOOP for the DVM SYNC */ 
svt_err_check_stats dvm_operation_dvm_sync_acsnoop_valid_value_check;
//-------------------------------------------------------------

/** Checks For a DVM Complete message, ARADDR is defined to be all zeros */
svt_err_check_stats dvmcomplete_araddr_valid_value_check;
//-------------------------------------------------------------
/** Checks  For a DVM Complete message, ACADDR is defined to be all zeros */
svt_err_check_stats dvmcomplete_acaddr_valid_value_check;
//-------------------------------------------------------------


/** Checks  FOR DVM Message the value of reserve address bit should be zero  */
svt_err_check_stats dvmmessage_araddr_reserve_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[11:10] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_hypervisor_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[9:8] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_secure_nonsecure_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[6] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_vmid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[5] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_asid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[0] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[0] of DVM message type Branch Predictor Invalidate */
svt_err_check_stats dvmmessage_branch_predictor_invalidate_supported_message_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[9:8] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_physical_inst_cache_secure_nonsecure_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[6:5] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_physical_inst_cache_vid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[0] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_physical_inst_cache_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[11:10] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_invalidate_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[9:8] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_secure_nonsecure_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[6] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_vmid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[5] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_asid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ARADDR[0] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_addr_specified_value_check;
//-------------------------------------------------------------


//DVM snoop

/** Checks  FOR DVM Message the value of reserve address bit should be zero  */
svt_err_check_stats dvmmessage_snoop_araddr_reserve_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[11:10] of DVM message type TLB Invalidate    */
svt_err_check_stats snoop_dvmmessage_tlb_hypervisor_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[9:8] of DVM message type TLB Invalidate    */
svt_err_check_stats snoop_dvmmessage_tlb_secure_nonsecure_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[6] of DVM message type TLB Invalidate    */
svt_err_check_stats snoop_dvmmessage_tlb_vmid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[5] of DVM message type TLB Invalidate    */
svt_err_check_stats snoop_dvmmessage_tlb_asid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[0] of DVM message type TLB Invalidate    */
svt_err_check_stats dvmmessage_tlb_snoop_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[0] of DVM message type Branch Predictor Invalidate */
svt_err_check_stats snoop_dvmmessage_branch_predictor_invalidate_supported_message_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[9:8] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_physical_inst_cache_secure_nonsecure_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[6:5] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_physical_inst_cache_vid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[0] of DVM message type Physical Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_physical_inst_cache_snoop_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[11:10] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_virtual_inst_cache_invalidate_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[9:8] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_virtual_inst_cache_secure_nonsecure_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[6] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_virtual_inst_cache_vmid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[5] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats snoop_dvmmessage_virtual_inst_cache_asid_value_check;
//-------------------------------------------------------------
/** Checks  the valid values of ACADDR[0] of DVM message type Virtual Instruction Cache Invalidate */
svt_err_check_stats dvmmessage_virtual_inst_cache_snoop_addr_specified_value_check;
//-------------------------------------------------------------
/** Checks the overlapping AWID of Write Barrier transactions with any active Write transactions */
svt_err_check_stats writebarrier_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks the overlapping ARID of Read Barrier transactions with any active Read transactions */
svt_err_check_stats readbarrier_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks the overlapping ARID of DVM transactions with any active Read transactions */
svt_err_check_stats dvm_xact_id_overlap_check;

/** Checks the overlapping ARID of Non-DVM or Non-Device transactions with any active transactions */
svt_err_check_stats read_non_dvm_non_device_xact_id_overlap_check;

/** Checks the overlapping AWID of Non-DVM or Non-Device transactions with any active transactions*/
svt_err_check_stats write_non_dvm_non_device_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks that all transactions of multi-part DVM operation have same ID */
svt_err_check_stats multipart_dvm_coherent_same_id_check;
//-------------------------------------------------------------
/** Checks that all transactions of multi-part DVM operation have same coherent response */
svt_err_check_stats multipart_dvm_coherent_same_response_check;
//-------------------------------------------------------------
/** Checks that all coherent transactions of multi-part DVM operation are sent in successive manner 
    and no unrelated coherent transaction sent during multi-part DVM opearion over AR channel */
svt_err_check_stats multipart_dvm_coherent_successive_transaction_check;
//-------------------------------------------------------------
/** Checks that all transactions of multi-part DVM operation have same snoop response */
svt_err_check_stats multipart_dvm_snoop_same_response_check;
//-------------------------------------------------------------
/** Checks that all snoop transactions of multi-part DVM operation are sent in successive manner 
    and no unrelated snoop transaction sent during multi-part DVM opearion over AC channel */
svt_err_check_stats multipart_dvm_snoop_successive_transaction_check;
//-------------------------------------------------------------
/** Checks the overlapping ARID of Non-Barrier Non-DVM transactions with any active Barrier/DVM transactions */
svt_err_check_stats readbarrier_dvm_norm_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks the overlapping AWID of Non-Barrier Non-DVM transactions with any active Barrier/DVM transactions */
svt_err_check_stats writebarrier_norm_xact_id_overlap_check;
//-------------------------------------------------------------
/** Checks the receiverd RDATACHK is same as the parity calculated from RDATA in a read  transaction */
svt_err_check_stats rdatachk_parity_calculated_rdata_parity_check;
//-------------------------------------------------------------
/** Checks the receiverd parity is same as the parity calculated from respective signal in a transaction */
svt_err_check_stats received_parity_calculated_parity_check;
//-------------------------------------------------------------
/** Checks the receiverd WDATACHK is same as the parity calculated from WDATA in a write transaction */
svt_err_check_stats wdatachk_parity_calculated_wdata_parity_check;
//-------------------------------------------------------------
/** Checks the receiverd CDDATACHK is same as the parity calculated from CDDATA in a snoop transaction */
svt_err_check_stats cddatachk_parity_calculated_cddata_parity_check;
//-------------------------------------------------------------

// Checks on 'Sequencing Transactions'

/** Checks that Master does not receive a snoop transaction until 
  * any preceding transaction to the same cache line has completed
  */
svt_err_check_stats resp_to_same_cache_line_check;
//-------------------------------------------------------------
/** Checks that if received a snoop transaction, response to a transaction 
  * to the same cache line is not received , until snoop response is sent 
  */
svt_err_check_stats snoop_to_same_cache_line_check;
//-------------------------------------------------------------
/**
  * Checks that the if DataTransfer de-asserted then no data transfer will occur on the snoop data channel
  *  for this transaction DataTransfer, CRRESP[0]
  */
svt_err_check_stats cdvalid_high_no_data_transfer_check;
//-------------------------------------------------------------
// START OF LOCKED ACCESS CHECKS
/**
  * Checks that there are no pending transactions before a locked
  * sequence starts
  */
svt_err_check_stats no_pending_xacts_during_locked_xact_sequeunce_check;
//-------------------------------------------------------------

/**
  * Checks that all transactions of locked sequence have the same id
  */
svt_err_check_stats locked_sequeunce_id_check;
//-------------------------------------------------------------

/**
  * Checks that when a master does a lock transaction, it does not target subsequent transactions in the lock 
  * sequence to any slave other than the locked slave
  */

svt_err_check_stats locked_sequence_to_same_slave_check;
 //----------------------------------------------------------------
/**
  * Check that the master follows as per the recommendation from spec to  limit 2 transaction for the lock access
  */
   svt_err_check_stats locked_sequence_length_check;
//-------------------------------------------------------------

/**
  * Checks that there are no pending transactions of a locked sequeunce
  * when a normal transaction is received
  */
svt_err_check_stats no_pending_locked_xacts_before_normal_xacts_check;
// END OF LOCKED ACCESS CHECKS

/** 
  * Checks that AXI master and AXI slave are not exceeding the user 
  * configured maximum number of outstanding transactions (#num_outstanding_xact)
  * If #num_outstanding_xact = -1 then #num_outstanding_xact will not be considered , 
  * instead #num_read_outstanding_xact and #num_write_outstanding_xact will be considered for 
  * read and write transactions respectively.
  */
svt_err_check_stats max_num_outstanding_xacts_check ;

//-------------------------------------------------------------
// START OF PERFORMANCE CHECKS
/**
  * Checks that the latency of a write transaction is not greater than the
  * configured max value
  */
svt_err_check_stats perf_max_write_xact_latency_check;

/**
  * Checks that the latency of a write transaction is not lesser than the
  * configured min value
  */
svt_err_check_stats perf_min_write_xact_latency_check;

/**
  * Checks that the average latency of write transactions in a given interval
  * is not more than the configured max value
  */
svt_err_check_stats perf_avg_max_write_xact_latency_check;

/**
  * Checks that the average latency of write transactions in a given interval
  * is not less than the configured min value
  */
svt_err_check_stats perf_avg_min_write_xact_latency_check;

/**
  * Checks that the latency of a read transaction is not greater than the
  * configured max value
  */
svt_err_check_stats perf_max_read_xact_latency_check;

/**
  * Checks that the latency of a read transaction is not lesser than the
  * configured min value
  */
svt_err_check_stats perf_min_read_xact_latency_check;

/**
  * Checks that the average latency of read transactions in a given interval
  * is not more than the configured max value
  */
svt_err_check_stats perf_avg_max_read_xact_latency_check;

/**
  * Checks that the average latency of read transactions in a given interval
  * is not less than the configured min value
  */
svt_err_check_stats perf_avg_min_read_xact_latency_check;

/**
  * Checks that the throughput of read transactions in a given interval is
  * not more that the configured max value
  */
svt_err_check_stats perf_max_read_throughput_check;

/**
  * Checks that the throughput of read transactions in a given interval is
  * not less that the configured min value
  */
svt_err_check_stats perf_min_read_throughput_check;

/**
  * Checks that the throughput of write transactions in a given interval is
  * not more that the configured max value
  */
svt_err_check_stats perf_max_write_throughput_check;

/**
  * Checks that the throughput of write transactions in a given interval is
  * not less that the configured min value
  */
svt_err_check_stats perf_min_write_throughput_check;

/**
  * Checks that the bandwidth of read transactions in a given interval is
  * not more that the configured max value
  */
svt_err_check_stats perf_max_read_bandwidth_check;

/**
  * Checks that the bandwidth of read transactions in a given interval is
  * not less that the configured min value
  */
svt_err_check_stats perf_min_read_bandwidth_check;

/**
  * Checks that the bandwidth of write transactions in a given interval is
  * not more that the configured max value
  */
svt_err_check_stats perf_max_write_bandwidth_check;

/**
  * Checks that the bandwidth of write transactions in a given interval is
  * not less that the configured min value
  */
svt_err_check_stats perf_min_write_bandwidth_check;

// END OF PERFORMANCE CHECKS
//-------------------------------------------------------------
// START Of STREAM CHECKS

svt_err_check_stats signal_valid_tvalid_check;

/** Checks that TREADY is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tready_when_tvalid_high_check;

/** If tdata is enabled, checks that TDATA is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tdata_when_tvalid_high_check;

/** If tstrb is enabled, checks that TSTRB is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tstrb_when_tvalid_high_check;

/** If tkeep is enabled, checks that TKEEP is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tkeep_when_tvalid_high_check;

/** If tlast is enabled, checks that TLAST is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tlast_when_tvalid_high_check;

/** If tid is enabled, checks that TID is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tid_when_tvalid_high_check;

/** If tuser is enabled, checks that TUSER is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tuser_when_tvalid_high_check;

/** If tdest is enabled, checks that TDEST is not X or Z when TVALID is high */
svt_err_check_stats signal_valid_tdest_when_tvalid_high_check;

/** 
  * Checks that TDATA is stable when TVALID is high 
  * When svt_axi_port_configuration::check_valid_data_bytes_only_enable=1 ,
  * it considers only valid byte lanes of tdata based on tstrb. 
  * When svt_axi_port_configuration::check_valid_data_bytes_only_enable=0 ,
  * whole tdata as seen on the bus will be considered.
  */
svt_err_check_stats signal_stable_tdata_when_tvalid_high_check;

/** Checks that TSTRB is stable when TVALID is high */
svt_err_check_stats signal_stable_tstrb_when_tvalid_high_check;

/** Checks that TKEEP is stable when TVALID is high */
svt_err_check_stats signal_stable_tkeep_when_tvalid_high_check;

/** Checks that TLAST is stable when TVALID is high */
svt_err_check_stats signal_stable_tlast_when_tvalid_high_check;

/** Checks that TID is stable when TVALID is high */
svt_err_check_stats signal_stable_tid_when_tvalid_high_check;

/** Checks that TUSER is stable when TVALID is high */
svt_err_check_stats signal_stable_tuser_when_tvalid_high_check;

/** Checks that TDEST is stable when TVALID is high */
svt_err_check_stats signal_stable_tdest_when_tvalid_high_check;

/** Checks that TVALID is low when reset is active */
svt_err_check_stats tvalid_low_when_reset_is_active_check;

/** Checks if tvalid was interrupted before tready got asserted */
svt_err_check_stats tvalid_interrupted_check;

/** Checks that TSTRB is low if TKEEP is low */
svt_err_check_stats tstrb_low_when_tkeep_low_check;

/** Checks that received data stream is not interleaved beyond stream_interleave_depth
  * value. An error is issued if data stream is interleaved beyond this value. */
svt_err_check_stats stream_interleave_depth_check;

/** Checks that the burst length of received data stream is not exceeding the maximum
  * value allowed for stream_burst_length defined by `SVT_AXI_MAX_STREAM_BURST_LENGTH. */
svt_err_check_stats max_stream_burst_length_exceeded_check;

/** 
 * @groupname port_interleaving_check
 * @check_description   
 * - Checks if address does fall to correct interleaved port.
 * - Valid when port cfg port_interleaving_enable = 1.   
 * .
 * @end_check_description
 *
 * @check_pass
 * address does fall to correct interleaved port. 
 * @end_check_pass
 *
 * @check_fail
 * address does not fall to correct interleaved port. 
 * @end_check_fail
 *
 * @applicable_device_type
 * master & slave 
 * @end_applicable_device_type
 *
 * @check_additional_information
 * @end_check_additional_information   
 */
svt_err_check_stats port_interleaving_check;

/** 
 * @groupname trace_tag_validity_check
 * @check_description   
 * - Trace tag value on data channel or resposne channel should be valid as per the trace tag 
 * - value on the address channel. 
 * .
 * @end_check_description
 *
 * @check_pass
 * For Write transactions the check will pass if:
 * A slave that receives a write request with AWTRACE asserted should assert the BTRACE signal alongside
 * the write response.
 * For Read transactions the check will pass if:
 * A slave that receives a read request with the ARTRACE signal asserted should assert the RTRACE signal
 * alongside every beat of the read response.
 * For Snoop transactions the check will pass if:
 * A master that receives a snoop request with the ACTRACE signal asserted should assert the CRTRACE
 * signal alongside the snoop response.The master should also assert CDTRACE alongside every data beat of
 * the snoop data that is associated with the snoop transaction.
 * @end_check_pass
 * @check_fail
 * If trace_tag in the request packet is set to 1 and in the spawned response or data packet is set 
 * to 0.
 * @end_check_fail
 *
 * @applicable_device_type
 * @end_applicable_device_type
 *
 * @check_additional_information
 * @end_check_additional_information   
 */
svt_err_check_stats trace_tag_validity_check;


// END OF STREAM CHECKS
//-------------------------------------------------------------
  `ifdef SVT_AXI_QVN_ENABLE
// START OF QVN CHECKS    

/** Checks that VARVALIDVN* is not X or Z */
svt_err_check_stats signal_valid_varvalidvnx_check;

/** Checks the VARQOSVN* is valid when VARVALIDVN* is high */
svt_err_check_stats  signal_valid_varqosvnx_when_varvalidvnx_high_check;  
   
/** Checks that VARREADYVN* is not X or Z */
svt_err_check_stats signal_valid_varreadyvnx_check;

/** Checks that VAWVALIDVN* is not X or Z */
svt_err_check_stats signal_valid_vawvalidvnx_check;

/** Checks the VAWQOSVN* is valid when VAWVALIDVN* is high */
svt_err_check_stats  signal_valid_vawqosvnx_when_vawvalidvnx_high_check;  
   
/** Checks that VAWREADYVN* is not X or Z */
svt_err_check_stats signal_valid_vawreadyvnx_check;
   
/** Checks that VWVALIDVN* is not X or Z */
svt_err_check_stats signal_valid_vwvalidvnx_check;

/** Checks that VWREADYVN* is not X or Z */
svt_err_check_stats signal_valid_vwreadyvnx_check;
   
/** Checks that VARVALIDVN* when asserted, remains asserted till VARREADYVN* */   
svt_err_check_stats varvalidvn_deassertion_check;
   
/** When a master sets VARVALIDVNx high, it can change VARQOSVNx proir to the slave granting a token, but only if the value increase. */
svt_err_check_stats varqosvn_valid_change_check;

/** Checks that VAWVALIDVN* when asserted, remains asserted till VAWREADYVN* */   
svt_err_check_stats vawvalidvn_deassertion_check;
   
/** When a master sets VAWVALIDVNx high, it can change VAWQOSVNx proir to the slave granting a token, but only if the value increase. */
svt_err_check_stats vawqosvn_valid_change_check;
   
/** Checks that VWVALIDVN* when asserted, remains asserted till VWREADYVN* */   
svt_err_check_stats vwvalidvn_deassertion_check;

/** Check that master must only set ARVNET to values that correspond to a VN where the associated set of token request signals exist.*/
svt_err_check_stats arvnet_for_existing_vn_check;
   
/** Check that master must only set AWVNET to values that correspond to a VN where the associated set of token request signals exist.*/
svt_err_check_stats awvnet_for_existing_vn_check;

/** Check that master must only set WVNET to values that correspond to a VN where the associated set of token request signals exist.*/
svt_err_check_stats wvnet_for_existing_vn_check;

/** Check that master must have read address token for VN denote ARVNET, before it can send read address channel transfer (Except for a Barrier transaction).*/
svt_err_check_stats rd_addr_chan_vn_token_availability_check;
   
/** Check that master must have write address token for VN denote AWVNET, before it can send write address channel transfer (Except for a Barrier transaction).*/
svt_err_check_stats wr_addr_chan_vn_token_availability_check;
   
/** Check that master must have write data token for VN denote WVNET, before it can send a data beat. */
svt_err_check_stats wr_data_chan_vn_token_availability_check;

/** Check that transaction with the same AXI ID that are are sent on the same physical link must use the same VN.*/
svt_err_check_stats same_axi_id_over_single_vn_check;

/** Check Before entering a low-power or reset state, the component must have the same number of pre-allocated tokens that it had when it exited reset.*/
svt_err_check_stats pre_allocated_token_count_at_rst_check;

/** Check QVN token handshake signal are not asserted on unsupported VN.*/
svt_err_check_stats qvn_sig_asrt_on_unsupported_vn_check;

/** Check that slave component is not granting more outstanding token than its configured.*/
svt_err_check_stats slave_max_outstanding_token_check;
   
/** Check that token requested should be granted in a bounded time*/
svt_err_check_stats qvn_token_request_timeout_check;
   
//-------------------------------------------------------------
// END OF QVN CHECKS    
`endif

`ifdef SVT_ACE5_ENABLE

//--------------------------------------------------------------
/** Checks that ARCHUNKEN is not X or Z when ARVALID is high */
svt_err_check_stats signal_valid_archunken_when_arvalid_high_check;

//--------------------------------------------------------------
/** Checks that RCHUNKV is not X or Z when RVALID is high */
svt_err_check_stats signal_valid_rchunkv_when_rvalid_high_check;
  
/** Checks that RCHUNKNUM is not X or Z when RVALID and RCHUNKV are high */
svt_err_check_stats signal_valid_rchunknum_when_rvalid_rchunkv_high_check;

/** Checks that RCHUNKSTRB is not X or Z when RVALID and RCHUNKV are high */
svt_err_check_stats signal_valid_rchunkstrb_when_rvalid_rchunkv_high_check;


//--------------------------------------------------------------
/** Checks that ARCHUNKEN is stable when ARVALID is high */
svt_err_check_stats signal_stable_archunken_when_arvalid_high_check;

//--------------------------------------------------------------
/** Checks that RCHUNKV is stable when RVALID is high */
svt_err_check_stats signal_stable_rchunkv_when_rvalid_high_check;

/** Checks that RCHUNKNUM is stable when RVALID and RCHUNKV are high */
svt_err_check_stats signal_stable_rchunknum_when_rvalid_rchunkv_high_check;

/** Checks that RCHUNKSTRB is stable when RVALID and RCHUNKV are high */
svt_err_check_stats signal_stable_rchunkstrb_when_rvalid_rchunkv_high_check;


//--------------------------------------------------------------
/** Checks that ARSIZE is equal to the data bus width or ARLEN is one beat and
 * ARSIZE is 128 bits or larger for rdata chunking */
svt_err_check_stats rdata_chunking_arsize_valid_value_check;

/** Checks that ARADDR is aligned to 16 bytes for rdata chunking */
svt_err_check_stats rdata_chunking_araddr_aligned_check; 

/** Checks that ARBURST is INCR or WRAP for rdata chunking */
svt_err_check_stats rdata_chunking_arburst_type_check;

/**Checks that ARSNOOP is ReadNoSnoop, ReadOnce, ReadOnceCleanInvalid or 
 * ReadOnceMakeInvalid for rdata chunking */
svt_err_check_stats rdata_chunking_arsnoop_valid_value_check;

/** Checks that ARIDUNQ must be asserted for rdata chunking */
svt_err_check_stats rdata_chunking_aridunq_valid_value_check;

//--------------------------------------------------------------  
/**Checks that RCHUNKV is deasserted for all the transfers when ARCHUNKEN is
 * deasserted */
svt_err_check_stats rdata_chunking_rchunkv_zero_when_archunken_deasserted_check;

/**Checks that RCHUNKV must be the same for every response beat of a 
 * transaction */ 
svt_err_check_stats rdata_chunking_rchunkv_same_for_all_response_check;

/** Checks that RCHUNKNUM must be between zero and ARLEN when RVALID and
 * RCHUNKV are high*/
svt_err_check_stats rdata_chunking_rchunknum_valid_value_check;

/**Checks that RCHUNKSTRB must not be zero when RVALID and RCHUNKV are high */
svt_err_check_stats rdata_chunking_rchunkstrb_valid_value_check;

/**Checks that the number of bytes that are transferred through read data
 * chunking must be consistant with ARSIZE and ARLEN */
svt_err_check_stats rdata_chunking_num_bytes_transfer_check;

`endif

`ifdef SVT_UVM_TECHNOLOGY
  /** UVM report server passed in through the constructor */
  uvm_report_object reporter;
`elsif SVT_OVM_TECHNOLOGY
  /** OVM report server passed in through the constructor */
  ovm_report_object reporter;
`else
  /** VMM message service passed in through the constructor*/ 
  vmm_log  log;
`endif

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   */
  extern function new (string name, svt_axi_port_configuration cfg, uvm_report_object reporter, bit register_enable=1, bit enable_pc_cov = 1);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param reporter OVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   */
  extern function new (string name, svt_axi_port_configuration cfg, ovm_report_object reporter, bit register_enable=1, bit enable_pc_cov = 1);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param log VMM log instance used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (string name, svt_axi_port_configuration cfg, vmm_log log = null, bit register_enable=1, bit enable_pc_cov = 1);
`endif
  /** @cond PRIVATE */
  extern function void perform_excl_write_addr_chan_signal_level_checks(svt_axi_transaction xact, 
                       svt_axi_transaction excl_xact, output bit is_excl_wr_error);
 
  extern function void perform_read_addr_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_arid,
                                                       ref logic[`SVT_AXI_MAX_ADDR_WIDTH-1:0] observed_araddr,
                                                       ref logic[`SVT_AXI_MAX_BURST_LENGTH_WIDTH-1:0] observed_arlen,
                                                       ref logic[`SVT_AXI_SIZE_WIDTH-1:0] observed_arsize,
                                                       ref logic[`SVT_AXI_BURST_WIDTH-1:0] observed_arburst,
                                                       ref logic[`SVT_AXI_LOCK_WIDTH-1:0] observed_arlock,
                                                       ref logic[`SVT_AXI_CACHE_WIDTH-1:0] observed_arcache,
                                                       ref logic[`SVT_AXI_PROT_WIDTH-1:0] observed_arprot,
                                                       ref logic[`SVT_AXI_QOS_WIDTH-1:0] observed_arqos,
                                                       ref logic[`SVT_AXI_REGION_WIDTH-1:0] observed_arregion,
                                                       ref logic[`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] observed_aruser,
                                                       ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_ardomain,
                                                       ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop,
                                                       ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar,
                                                       ref logic observed_arready,
`ifdef SVT_ACE5_ENABLE
                                                       ref logic[`SVT_AXI_MAX_MMUSID_WIDTH-1:0]observed_stream_id,
                                                       ref logic[`SVT_AXI_MAX_MMUSSID_WIDTH-1:0]observed_sub_stream_id,
                                                       ref logic observed_secure_or_non_secure_stream,
                                                       ref logic observed_sub_stream_id_valid,
                                                       ref logic observed_addr_translated_from_pcie,
                                                       ref logic observed_aridunq, 
                                                       ref logic observed_archunken,
                                                       ref logic [`SVT_AXI_MAX_MPAM_WIDTH-1:0] observed_armpam,
                                                       output bit is_aridunq_valid, 
                                                       output bit is_archunken_valid,
                                                       output bit is_stream_id_valid,                              
                                                       output bit is_sub_stream_id_valid,                          
                                                       output bit is_secure_or_non_secure_stream_valid,                              
                                                       output bit is_sub_streamid_valid,                          
                                                       output bit is_addr_translated_from_pcie_valid,
                                                       output bit is_armpam_valid,     
 `endif
                                                       output bit is_arid_valid,
                                                       output bit is_araddr_valid,
                                                       output bit is_arlen_valid,
                                                       output bit is_arsize_valid,
                                                       output bit is_arburst_valid,
                                                       output bit is_arlock_valid,
                                                       output bit is_arcache_valid,
                                                       output bit is_arprot_valid,
                                                       output bit is_arqos_valid,
                                                       output bit is_arregion_valid,
                                                       output bit is_aruser_valid,
                                                       output bit is_ardomain_valid,
                                                       output bit is_arsnoop_valid,
                                                       output bit is_arbar_valid,
                                                       output bit is_arready_valid,
                                                       output bit excl_read_error
                                                     );
  extern function void perform_read_data_chan_signal_level_checks(
                                                      ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_rid,
                                                      ref logic[`SVT_AXI_RESP_WIDTH-1:0] observed_rresp,
                                                      ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] observed_rdata,
                                                      ref logic[`SVT_AXI_MAX_POISON_WIDTH-1:0] observed_rpoison,
                                                      ref logic observed_rlast,
                                                      ref logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] observed_ruser,
                                                      ref logic observed_rready,
 `ifdef SVT_ACE5_ENABLE
                                                      ref logic observed_ridunq, 
                                                      ref logic observed_rchunkv,
                                                      ref logic [`SVT_AXI_MAX_CHUNK_NUM_WIDTH-1:0] observed_rchunknum,
                                                      ref logic [`SVT_AXI_MAX_CHUNK_STROBE_WIDTH-1:0] observed_rchunkstrb,
                                                      output bit is_ridunq_valid, 
                                                      output bit is_rchunkv_valid,
                                                      output bit is_rchunknum_valid,
                                                      output bit is_rchunkstrb_valid,
 `endif
                                                      output bit is_rid_valid,
                                                      output bit is_rresp_valid,
                                                      output bit is_rdata_valid,
                                                      output bit is_rpoison_valid,
                                                      output bit is_rlast_valid,
                                                      output bit is_ruser_valid,
                                                      output bit is_rready_valid
                                                    );
  extern function void perform_write_addr_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_awid,
                                                       ref logic[`SVT_AXI_MAX_ADDR_WIDTH-1:0] observed_awaddr,
                                                       ref logic[`SVT_AXI_MAX_BURST_LENGTH_WIDTH-1:0] observed_awlen,
                                                       ref logic[`SVT_AXI_SIZE_WIDTH-1:0] observed_awsize,
                                                       ref logic[`SVT_AXI_BURST_WIDTH-1:0] observed_awburst,
                                                       ref logic[`SVT_AXI_LOCK_WIDTH-1:0] observed_awlock,
                                                       ref logic[`SVT_AXI_CACHE_WIDTH-1:0] observed_awcache,
                                                       ref logic[`SVT_AXI_PROT_WIDTH-1:0] observed_awprot,
                                                       ref logic[`SVT_AXI_QOS_WIDTH-1:0] observed_awqos,
                                                       ref logic[`SVT_AXI_REGION_WIDTH-1:0] observed_awregion,
                                                       ref logic[`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] observed_awuser,
                                                       ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_awdomain,
                                                       ref logic[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] observed_awsnoop,
                                                       ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_awbar,
`ifdef SVT_ACE5_ENABLE
                                                       ref logic[`SVT_AXI_STASH_NID_WIDTH-1:0]observed_stash_nid,
                                                       ref logic[`SVT_AXI_STASH_LPID_WIDTH-1:0]observed_stash_lpid,
                                                       ref logic observed_stash_nid_valid,
                                                       ref logic observed_stash_lpid_valid,
                                                       output bit is_stash_nid_valid,                              
                                                       output bit is_stash_lpid_valid,                          
                                                       output bit is_stashnid_valid,                              
                                                       output bit is_stashlpid_valid,                          
                                                       ref logic[`SVT_AXI_MAX_MMUSID_WIDTH-1:0]observed_stream_id,
                                                       ref logic[`SVT_AXI_MAX_MMUSSID_WIDTH-1:0]observed_sub_stream_id,
                                                       ref logic observed_secure_or_non_secure_stream,
                                                       ref logic observed_sub_stream_id_valid,
                                                       ref logic observed_addr_translated_from_pcie,
                                                       ref logic [`SVT_ACE5_ATOMIC_TYPE_WIDTH-1:0] observed_awatop,
                                                       ref logic [`SVT_AXI_MAX_MPAM_WIDTH-1:0] observed_awmpam,
                                                       output bit is_stream_id_valid,                              
                                                       output bit is_sub_stream_id_valid,                          
                                                       output bit is_secure_or_non_secure_stream_valid,                              
                                                       output bit is_sub_streamid_valid,                          
                                                       output bit is_addr_translated_from_pcie_valid,                          
                                                       output bit is_awatop_valid,
                                                       ref logic observed_awidunq,
                                                       output bit is_awidunq_valid,
                                                       output bit is_awmpam_valid,
`endif
                                                       ref logic observed_awready,
                                                       ref logic observed_awunique,
                                                       output bit is_awid_valid,
                                                       output bit is_awaddr_valid,
                                                       output bit is_awlen_valid,
                                                       output bit is_awsize_valid,
                                                       output bit is_awburst_valid,
                                                       output bit is_awlock_valid,
                                                       output bit is_awcache_valid,
                                                       output bit is_awprot_valid,
                                                       output bit is_awqos_valid,
                                                       output bit is_awregion_valid,
                                                       output bit is_awuser_valid,
                                                       output bit is_awdomain_valid,
                                                       output bit is_awsnoop_valid,
                                                       output bit is_awbar_valid,
                                                       output bit is_awready_valid,
                                                       output bit excl_write_error,
                                                       output bit is_awunique_valid
                                                     );
  extern function void perform_write_data_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_wid,
                                                       ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] observed_wdata,
                                                       ref logic[(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] observed_wdatachk,
                                                       ref logic[`SVT_AXI_MAX_POISON_WIDTH-1:0] observed_wpoison,
                                                       ref logic[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] observed_wstrb,
                                                       ref logic observed_wlast,
                                                       ref logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] observed_wuser,
                                                       ref logic observed_wready,
                                                       output bit is_wid_valid,
                                                       output bit is_wdata_valid,
                                                       output bit is_wdatachk_valid,
                                                       output bit is_wpoison_valid,
                                                       output bit is_wstrb_valid,
                                                       output bit is_wlast_valid,
                                                       output bit is_wuser_valid,
                                                       output bit is_wready_valid
                                                     );
  extern function void perform_write_resp_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_MAX_ID_WIDTH-1:0] observed_bid,
                                                       ref logic[`SVT_AXI_RESP_WIDTH-1:0] observed_bresp,
                                                       ref logic[`SVT_AXI_MAX_BRESP_USER_WIDTH-1:0] observed_buser,
                                                       ref logic observed_bready,
 `ifdef SVT_ACE5_ENABLE
                                                       ref logic observed_bidunq, 
                                                       output bit is_bidunq_valid, 
 `endif
                                                       output bit is_bid_valid,
                                                       output bit is_bresp_valid,
                                                       output bit is_buser_valid,
                                                       output bit is_bready_valid
                                                     );
  extern function void perform_data_stream_signal_level_checks(ref logic observed_tready,
                                                        logic[`SVT_AXI_MAX_TDATA_WIDTH-1:0] observed_tdata,
                                                        logic[`SVT_AXI_TSTRB_WIDTH-1:0] observed_tstrb,
                                                        logic[`SVT_AXI_TKEEP_WIDTH-1:0] observed_tkeep,
                                                        logic observed_tlast,
                                                        logic[`SVT_AXI_MAX_TID_WIDTH-1:0] observed_tid,
                                                        logic[`SVT_AXI_MAX_TDEST_WIDTH-1:0] observed_tdest,
                                                        logic[`SVT_AXI_MAX_TUSER_WIDTH-1:0] observed_tuser,
                                                        output bit is_tready_valid,
                                                        output bit is_tdata_valid,
                                                        output bit is_tstrb_valid,
                                                        output bit is_tkeep_valid,
                                                        output bit is_tlast_valid,
                                                        output bit is_tid_valid,
                                                        output bit is_tdest_valid,
                                                        output bit is_tuser_valid);

  extern function void perform_slave_reset_checks(logic observed_rvalid, logic observed_bvalid);
  extern function void perform_master_reset_checks(logic observed_arvalid, logic observed_awvalid, logic observed_wvalid);
  extern function void perform_master_reset_ace_checks(logic observed_crvalid, logic observed_cdvalid);
  extern function void perform_slave_reset_ace_checks(logic observed_acvalid);
  extern function void perform_master_reset_stream_checks(logic observed_tvalid);
  /** Performs checks on AWUNIQUE signal for WRITECLEAN and WRITEEVICT transactions */
  extern function void perform_awunique_checks(logic observed_awunique, svt_axi_transaction xact);
  /**
    * Performs check on WRITEEVICT transaction that all wstrb signals must be asserted
    * @param xact Transaction on which check is to be done
    * @param check_all_beats Indicates if check is to be done on current beat or on all beats
    */
  extern function void perform_coherent_xact_wstrb_check(svt_axi_transaction xact, bit check_all_beats);
  extern function void reset_internal_variables();

  extern function void perform_burst_4k_boundary_cross_check  (svt_axi_transaction xact);
  extern function void perform_burst_wrap_address_align_check (svt_axi_transaction xact);
  extern function void perform_burst_wrap_burst_length_check  (svt_axi_transaction xact);
  extern function void perform_burst_size_not_exceed_data_width_check(svt_axi_transaction xact);
  extern function void perform_write_burst_value_check  (ref logic observed_awvalid, ref logic[`SVT_AXI_BURST_WIDTH-1:0] observed_awburst);
  extern function void perform_write_valid_awcache_check(ref logic observed_awvalid,input svt_axi_transaction xact);
  extern function void perform_read_burst_value_check  (ref logic observed_arvalid, ref logic[`SVT_AXI_BURST_WIDTH-1:0] observed_arburwst);
  extern function void perform_read_valid_arcache_check(ref logic observed_arvalid, input svt_axi_transaction xact);
  extern function void perform_write_resp_write_data_check(svt_axi_transaction xact);
  extern function void perform_write_resp_write_address_check(svt_axi_transaction xact);

  extern function void perform_snoop_addr_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_ACE_SNOOP_ADDR_WIDTH-1:0] observed_acaddr,
                                                       ref logic[`SVT_AXI_ACE_SNOOP_TYPE_WIDTH-1:0] observed_acsnoop,
                                                       ref logic[`SVT_AXI_ACE_SNOOP_PROT_WIDTH-1:0] observed_acprot,
                                                       ref logic observed_acready,
                                                       output bit is_acaddr_valid,
                                                       output bit is_acsnoop_valid,
                                                       output bit is_acprot_valid,
                                                       output bit is_acready_valid
                                                     );
  extern function void perform_snoop_data_chan_signal_level_checks(
                                                      ref logic[`SVT_AXI_ACE_SNOOP_DATA_WIDTH-1:0] observed_cddata,
                                                      ref logic[(`SVT_AXI_ACE_SNOOP_DATA_WIDTH/8)-1:0] observed_cddatachk,
                                                      ref logic[`SVT_AXI_ACE_SNOOP_POISON_WIDTH-1:0] observed_cdpoison,
                                                      ref logic observed_cdlast,
                                                      ref logic observed_cdready,
                                                      output bit is_cddata_valid,
                                                      output bit is_cddatachk_valid,
                                                      output bit is_cdpoison_valid,
                                                      output bit is_cdlast_valid,
                                                      output bit is_cdready_valid
                                                    );
  extern function void perform_snoop_resp_chan_signal_level_checks(
                                                       ref logic[`SVT_AXI_ACE_SNOOP_RESP_WIDTH-1:0] observed_crresp,
                                                       ref logic observed_crready,
                                                       output bit is_crresp_valid,
                                                       output bit is_crready_valid
                                                     );
  extern function void perform_axcache_axdomain_restriction_check(svt_axi_transaction xact);
  extern function void perform_axcache_axdomain_invalid_value_check(svt_axi_transaction xact);
  extern function void perform_cache_line_size_transaction_constraint_check(svt_axi_transaction xact);
  extern function void perform_readonce_writeunique_transaction_check(svt_axi_transaction xact);
  extern function void perform_writeback_writeclean_transaction_check(svt_axi_transaction xact);
  extern function void perform_axi_transaction_check(svt_axi_transaction xact);
  extern function void perform_read_data_channel_signal_value_check(svt_axi_transaction xact);
  extern function void perform_write_response_channel_signal_value_check(svt_axi_transaction xact,ref logic[`SVT_AXI_RESP_WIDTH-1:0] observed_bresp);
  extern function void perform_dvm_snoop_response_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_acsnoop_reserved_value_check(ref logic [`SVT_AXI_ACE_SNOOP_TYPE_WIDTH-1:0] observed_acsnoop);
  extern function void perform_snoop_resp_passdirty_datatransfer_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_full_cache_line_datatransfer_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_cdvalid_high_no_data_transfer_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_snoop_response_channel_isshared_check(svt_axi_snoop_transaction snoop_xact);
  extern function void perform_fixed_burst_type_valid_check(svt_axi_transaction xact);
  extern function void perform_snoop_addr_snoop_resp_check(svt_axi_snoop_transaction snoop_xact );
  extern function void perform_snoop_addr_snoop_data_check(svt_axi_snoop_transaction snoop_xact );

  extern function void perform_arsnoop_ardomain_arbar_reserve_value_check(ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop, 
  ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_ardomain, 
  ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar);

  extern function void perform_awsnoop_awdomain_awbar_reserve_value_check(ref logic[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] observed_awsnoop,
                                                                          ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_awdomain,
                                                                          ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_awbar);

//--- Barrier Checks --//
  extern function void perform_write_barrier_transaction_check (svt_axi_transaction xact,ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_awbar,
                                                                 ref logic[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] observed_awsnoop);
  extern function void  perform_read_barrier_transaction_check(svt_axi_transaction xact,ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar,
ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop);
  extern function void perform_barrier_id_check(svt_axi_transaction xact);
  extern function void perform_barrier_read_response_check(svt_axi_transaction xact, ref logic[1:0]  observed_rresp ,ref logic observed_rlast);
  extern function void perform_barrier_write_response_check(svt_axi_transaction xact, ref logic[1:0] observed_bresp);
  extern function void perform_rack_status_check(svt_axi_transaction xact, logic observed_ack );
  extern function void perform_wack_status_check(svt_axi_transaction xact, logic observed_ack );


//--- DVM Checks --//

  extern function void  perform_dvm_read_address_channel_check(svt_axi_transaction xact,ref logic[`SVT_AXI_ACE_BARRIER_WIDTH-1:0] observed_arbar,
                                                       ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop,
                                                       ref logic[`SVT_AXI_ACE_DOMAIN_WIDTH-1:0] observed_ardomain);

  extern function void  perform_dvm_arsnoop_read_address_channel_valid_check(svt_axi_transaction xact,
                                                                     ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_arsnoop,
                                                                     ref logic[`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0] observed_araddr);
  extern function void  perform_dvm_acsnoop_snoop_address_channel_valid_check(svt_axi_snoop_transaction xact,
                                                                      ref logic[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] observed_acsnoop,
                                                                      ref logic[`SVT_AXI_ACE_SNOOP_ADDR_WIDTH-1 : 0] observed_acaddr);
  extern function void perform_dvmcomplete_araddr_valid_value_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_araddr_reserve_value_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_tlb_invalidate_supported_message_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_branch_predictor_invalidate_supported_message_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_physical_inst_cache_invalidate_supported_message_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_virtual_inst_cache_invalidate_supported_message_check(svt_axi_transaction xact);
  extern function void perform_dvmmessage_snoop_araddr_reserve_value_check(svt_axi_snoop_transaction xact);
  extern function void perform_dvmcomplete_acaddr_valid_value_check(svt_axi_snoop_transaction xact);
  extern function void perform_snoop_dvmmessage_tlb_invalidate_supported_message_check(svt_axi_snoop_transaction xact);
  extern function void perform_snoop_dvmmessage_branch_predictor_invalidate_supported_message_check(svt_axi_snoop_transaction xact);
  extern function void perform_snoop_dvmmessage_physical_inst_cache_invalidate_supported_message_check(svt_axi_snoop_transaction xact);
  extern function void perform_snoop_dvmmessage_virtual_inst_cache_invalidate_supported_message_check(svt_axi_snoop_transaction xact);
  extern function svt_axi_transaction perform_barrier_dvm_normal_xact_id_overlap_check(svt_axi_transaction xact, svt_axi_transaction active_queue[$], bit execute_check=1);
  extern function void perform_barrier_pair_check(svt_axi_transaction xact);
  extern function void perform_atomicity_size_alignment_check(svt_axi_transaction xact);

`ifdef SVT_ACE5_ENABLE
//--- UNIQUE_ID - OUTSTANDING Checks --//
  extern function svt_axi_transaction perform_no_unique_id_outstanding_transaction_with_same_id(svt_axi_transaction xact, svt_axi_transaction active_queue[$]);
`endif 

//--- NON - DVM Checks --//
  extern function svt_axi_transaction perform_non_dvm_non_device_with_overlap_id_check(svt_axi_transaction xact, svt_axi_transaction active_queue[$]);

  `ifdef SVT_AXI_QVN_ENABLE
//--- QVN Checks --//   
  extern function void perform_qvn_wr_addr_token_handshake_checks(logic       observed_vawvalidvnx,
                  logic       observed_vawreadyvnx,
                  logic [3:0] observed_vawqosvnx,
                  logic [3:0] vnet_id);
   
  extern function void perform_qvn_wr_data_token_handshake_checks(logic       observed_vwvalidvnx,
                  logic       observed_vwreadyvnx,
                  logic [3:0] vnet_id);

  extern function void perform_qvn_wr_addr_chan_sig_assertion_on_unsupported_vn_check(logic       observed_vawvalidvnx,
                          logic     observed_vawreadyvnx,
                          logic [3:0] vnet_id);

  extern function void perform_qvn_wr_data_chan_sig_assertion_on_unsupported_vn_check(logic     observed_vwvalidvnx,
                          logic     observed_vwreadyvnx,
                          logic [3:0] vnet_id);

   extern function void perform_qvn_rd_addr_token_handshake_checks(logic       observed_varvalidvnx,
                   logic       observed_varreadyvnx,
                   logic [3:0] observed_varqosvnx,
                   logic [3:0] vnet_id);
   
   extern function void perform_qvn_rd_addr_chan_sig_assertion_on_unsupported_vn_check(logic       observed_varvalidvnx,
                           logic     observed_varreadyvnx,
                           logic [3:0] vnet_id);
  `endif
  extern function void set_default_pass_effect(svt_err_check_stats::fail_effect_enum default_pass_effect);
  extern function void execute(svt_err_check_stats check_stats, bit test_pass, string fail_msg="",
                               svt_err_check_stats::fail_effect_enum fail_effect=svt_err_check_stats::ERROR);

  extern function void register_err_checks(bit en = 1'b1);

  extern function void passive_cache_check_post_coherent(coherency_error_type_enum err_status, svt_axi_transaction xact, svt_axi_passive_cache_line::passive_state_enum initial_state);

  extern virtual function void passive_cache_check_post_snoop(coherency_error_type_enum err_status, svt_axi_snoop_transaction xact, svt_axi_passive_cache_line::passive_state_enum initial_state);

  extern virtual function void perform_multipart_dvm_coherent_start_check(svt_axi_transaction xact, bit drop_xact_if_error=0);

  extern virtual function void perform_multipart_dvm_coherent_response_check(svt_axi_transaction xact);

  extern virtual function void perform_multipart_dvm_snoop_start_check(svt_axi_snoop_transaction xact);

  extern virtual function void perform_multipart_dvm_snoop_response_check(svt_axi_snoop_transaction xact);

  extern virtual function void update_checks_on_reset(svt_axi_transaction xact = null);

  extern virtual function bit is_current_xact_multipart_dvm(svt_axi_transaction xact);
  extern virtual function bit is_snoop_xact_multipart_dvm(svt_axi_snoop_transaction xact);

  /** 
    * This task waits for the last transaction of a multipart DVM. 
    */
  extern task check_and_wait_for_last_multipart_coherent_dvm_xact();

  /** Returns 1 if only the first part of a multi-part dvm is received */
  extern function bit is_second_part_of_multipart_pending();

  extern virtual function void disable_ace_checks();

  extern virtual function void reset_multipart_dvm();

  extern virtual function void reset_barrier_checks();

`ifdef SVT_ACE5_ENABLE
  // E1.11.1 (IHI0022H) Constraints for rdata chunking for AXI Transaction
  extern virtual function void perform_rdata_chunking_check(svt_axi_transaction xact);
  extern virtual function void perform_rdata_chunking_num_bytes_transfer_check(svt_axi_transaction xact, logic observed_rchunkv, logic observed_rlast);
`endif
/** @endcond */

endclass

//----------------------------------------------------------------
/**
AXI  port monitor check description
*/

`protected
eC(LbUBgOX]?Q066?PAD#UG_0#A8Y9/HMG.H8#1UUN-9WCg#BM&8))70^V^HD2Kg
7-g(6^a5N/d+FgP8\f0bVX/B?V,1GI,2I7WV[c5X=7PS+]JB]RQF\]X6WCfF,KFZ
8CE,JC.]LJTX&WfAf-(J0XXE9#1OY3Jg(;gg(M2DQJB6+JA0ae+7\M-:N5a[J?0D
4GJ=_GN0g[JSYQ#;VR0/66NW29P2^2][9@d)0Rd4=M+QaX-ff;f#f9>AeV,RU9^?
=L:GXf7J<(1c1BOQHeT=62=,7QLVE5SG15?eY=5?GW(dZH5ESd\\,UZ1eMXV8c,:
47,/:Y810IZOLRG/gFcK>C63WGJ>7QS=fP),I68e_>^E3_e7(=gd::DE^:^cS1SO
O\(M1[:>DH?=1dcP=@XD[+d1><-^Q-TZ]1AABZ]@NM)9L/M\N.&TNQ7EX#NX1a40
[I?_.C,XB;a&<cZ5-Ha^Cc\UgV1K@X>-bQRV9g&087f[g#3VEVONfc@>((O>C.ea
@_+F42:4MEF?0Q;Z^6=\CJT>P\E[=K8>NFGVK])CebK^#RZTDP;O-:34^.N,]G6+
QdTS7?N9=07QCPUG7K64L^7=]3a6PA_W/YW2PJKM]^QZ&1X\5M_T)[>QL8[,99Tf
23_LXI5?XK9(f\>+TKE)aQ7LE4@=W7Cdf^26=KU\-)FcIfR4IV7Z\0<KSC/?D^+3
:UCKSTUc3@LI0US\FO5[3U&XPaEU?>f[+N/\^6\;Q4TFSXVWS_AMYdge8(7MgYbN
+Z=D:FJ-aT(5.Z?3T5;I:90C9,K6I7@VJAcL;DMd3U)BR(fBY&J+?GG^DX=C,]XV
J(6-DV-?B#\V2.4J:I<bK6]O>C5FCf>&)0=>_P.)YWK/:,T5[2#[+<cFT5c0]KdR
)=E[78FEf::7e>,]3=@72^KgT8L/C(AS]0DV\HIX>fD.EUR/=?1Q.]0@S&D--EVb
)_5LSZ-V[7,W3V,P15/?46bMY;)VCBO^D\Oe6Idd<FAF#TJdZIO0dI6UUFXf>4ad
dE(a((6#TY?EZ;=@L4RV@gK7b[/P7b@H(I7VY5Yf-3)YO2S117ed2;ab[SJ,9f]2
MO-1cdQ\-7L\K=X2C/=L_VGb9Z3;M_^(?e:f(d-.f94XGFe1<@,PQ+<4[N,.1bOE
c1<I3a+G_0.Cg-cOX9>c,?S7a@#I39HfgFX4<e3e.R[WOXTL/FCX/F\.BMN<Z5M2
eL8:=;?R/9LTMBB:c/1&&W)Q\51WQ]WKT/(_=dGGbHL15G\f&PJQ7@P0)G[>Z84]
Pe4T;QLdI)E5\H81Y+N>(eG??IWWL;[QF^+NQ@118JbbL;X55YX=3)K3B.Ce#8MX
EFWdAT:FRM?bB6_[-[M;=#NGIR#;7KFQU+BON7KVd=N3LO2U1-5D<F_+90>NL.=;
f&CC>;56.[61AJ@)]GLJ_\<CSNFAbF,^[SFDbUB[2Pcc,,Ib(><LV7WgHC:789\+
aIJLd87F6LH=A/[WQfD9Z=Dg8KEI\ESJB;W+F/Q?P<NR:4TV5f6(RG\YXQX]IaYU
R\K6E[:-TOg-(<6(D#/9F01I0#E;0=R2UeITZ#\gEK512O:d=fS-a,J;2AMdfUa=
LJ9eW-gXQF0YZ.c.dE]>2R7IU1><GE,;\>2Wg\BH^CZ95^0]>e7ZF]6Q[5W<#RWZ
JAFWf3Y.6[McJ;LTBKKN\)APc-F542#;g=H9LJM7=902dHFZYJW1]O0;T(f;\RSC
=4FYC4a9<IAV#:<Oc&@cM5#RaYIB6P9S].-8:+CY&KUSW?Ug9,)eDF<;gMC=@7.T
;INbGE7;GFVK0C5a7+\ZT@C.IA4A#DXT?(;J_dV\[ON7SWGK(R^,XaCP3Bb]TMIP
A4LJ[K=-+KBA^Sb);Bc;I:Xa+])P_Vb;E?1S&0H/VFeH#AN;5AOdCA-)D,Y2fDDR
H+-<b@+4:PI70R4V&BE7@8WE0?S6)cWA=3MHKF@15M=V^f]WEGBCHES/SgdI9BNf
CD-O6#f]\>NW<gN=F2<F>+LKgLY5PRbg<BFLI)9aIE1F=BQ5aWB/I&A92/W=7EcC
LS-JeNf8CCLSO8Ig]_\aa&+aDX0>,=e/FBN,1#44,0A+9[c]^K=9<=22&b#\PHDf
I(I6Q3WU]LH0-R&,F1O(]c_X4ed@.Vb_Y[2&4ED^:V6I(PO]D)d,QFULV8YYWfXV
_/@\TI.LbaWV-S(6IS4WfZ1f>Q?IVTJH46:gGBNT?HR9;6VOM29\C[37;)H^Z=fY
0bAF22GY)Y[P_TQ[d>MG_bBfM1^d<H]62(KJ)(AKR00Aa683g+@&=GDfVB,[&-Y?
Ff<M^?EILPfFK3K(ceOB6P8d<VS9\,96BCSZ=XZQ8SH98(8:=)(cGdD9+6M-;,P\
H@I,T[dDAc.5\8:6\ZQ(Q3=5=M5LSO7GPKBXX[Z,\#JOW#/PRb7R85baac/)?#P_
c-4#M5=1.Fd/5_WE11C)@7ZI0UYPO#-_S,3M#N;U\CT?N/8eCMS=eLIa7fLVU>;D
R]#IL/BK6V5]I#Bc@4?5cScGPP3TM</_+VgdaEJH,3Ze(R_<#KB(A63X0e#X6,f&
RTa9;Y#Q@?2Z\[--PIT9LaK:,JUB.TP&@+:^S-/K8Z]6^7J9O#ObNIO.QU;&M82f
YC-AQ@FH>NC/8I_@PGQ#VYbJ(?fNad_JaLZ&C+EAbU#94(?XaS]GHB[.SQe/U/?I
FZ]=O+KA[H;&QJ2Z2Dg+UR;X37>GLBPD=GQ;2bc0eMDaCY5#LQD09V2)FOa;Z70b
/.X9fC.W@G[Z1U7/YCdTe<Q-P1HHC=LLQ;/(;X]^=IMOG0>4b5AXTg[\R5\F-e<Z
EOg9>#6?fFc?,GI8O:ZYUJ?):C)_b@Z07Z?T<2[<2[Oe9+.CNgd22^B;MFML+>G_
EdF&CM&KX2=\E#XROf:82Iaa_W=Z_.]A^B_W=.XN4E=)O)G&Hd/GR9)TBAF/C&8/
)Q;(BgT_URD&\e?U#(?A=Ie4@/g_/VYC?U(8[NPQYI>##d,(,I;a=QI-,gS.TCC>
J<Q=A^O?2I1;.;RVX1B6-2W/XW=K=I1d=6f_93(WbOce_@YMDCbeb^6SWI/D<8XL
.HeLKITP?HQ:I>/E[NBeJ7,c/F.7H,#ee3//&50g(NZJ:Ub@8aa?#:W9GWQVK35P
,TGdF/E]&agG8<HX?9=@1B@.F/gTD7T>?):UVA+N0=:#,M9TE_7AX+S(GK)Tg&ZI
I<MJ)Qd8\J<_(\??JKf>Z:[:b#-S2H+X^ETcA)AJ@#F3PH6EF1A[fWVe_Xa1?Z4-
7;3dNDDB>.<YI\T]a3DUGV6E3]Z#U<f2dg4X(F4;dP:K_)1/=/cAe;)42IM(+9d8
A>\aZI-G946SQ\f0_P0;6DbW3Be7M_NI1M[EPZc:7JVTP8T=DH6Z#)9O/EGQeW)#
XPd8fTU:/9N6X(F^Td,>SNe?ROMU7R<5QGJV)#ER4OH<R?I=1:&9HDE&C]PQA20F
L]5O;eU5LED@5DB(T8cTBP>fe.BTZ7:+&#EYN:+6aD#B>^Bg906B-1b<EN@d5Z-U
Q;0,bL+<MC-O=?LU)dR@:;U,\f)Z3G->#FWFU0V;PC4L]D?Z@MO1JW+0R/C75=6K
2G+^/#Ge6KST]/]4@[_&I-T]D6.-af]0QIFa6Mg7S3?bEGdA&bIRCA5<TOW0/eQ>
YCbY9IYW(&W=P06.M4298=2.^(@>4G-g3BKW<2Ig6c5Z\T4H#1UCKXA858T<-Y?>
J&=JC8.(L/4(AbF)ZRQ?b;_Kf?@4+3I>3^^a+IcS,7L0Sb19YG25A5-QDAYIGJ(S
,/LJEMQK@aPF72]DO_1+_5=CR9AW=V#RC(FEO/BT1.<Pg<\X/I6ANCb\>[aL2<>e
8\#??Hd._W?/OcQS9NE_0@3XCQ_44X:c#F7/58T7K2-^,?-3M8K4&F6@PZ(O4N2Z
/Z-3P5:D-f:IH@a_9?G^AZW.-<aEJbNbLJ,aRaDWG4X5+J.7[W#RU[0CT;#F-D)_
@868_N7Ac+?^Y;fd3e\\d\A5fV6_-VVM4TACCD4\F^I.QX-G66>.8CdFZ5UD>/B;
I-?2MK<?VMDU31K4dXB=ER[5#2BaC/XG6g@COA6,6,XV))e:#[V8<8JZ/=I7-Q@Q
=Qe(G^F\ca(Kd3R(3.D#(OQ3A,A]--9QC)b2,9:c:a?f4FN\EVeC^3e:T??.A>3e
/^P(U^-F0,cGfc[LQ0\-XOU#17?&#O6P.3bNFCKdg#QPLF;TZN8Y5R<b6V>&U_JN
HK^g?BeMWM#B;cZX7_\eSRQ0Q6,dg:9G-DG<-AIEA75LWL/]e)T.IdDbN:f9]VK0
GUY\-XT)B24P2JB:1T>\?7/<B/,_85<g_(@M3O2NNJCBBb?-K=IBZO1L\J/0(T;;
QZ;eOR<JPX,g@ZbgbK?\?ge.8:e5YQ=#Ig?>1L9YL_3^J&G,VGRF_LYaJGb2AI/O
Z&F>2#FB0aR3__HFf[Id.C&HB51S_g1_@)Y]#8AP\fYIRW^_D2g+;>L0,,CTBa\P
M]CHDO9:U-T;9A[?\OI5GcUfg\5EBKHM8(:4JB\5+YWF8/bc7Y<gd6-ORc<U#MTJ
5R5,EA55O?M07;[[:4A.B:##KM15JQDa54#e9MW^<fN>cI>&gf<+[c[#8._)a:72
UFY4FA-f=(:?_WZR0.S0/OPG=;P:SacO07AQ3_6R\-I4K:ERI#g6G+DHcNO4SE9g
/2V@&#d3\#-#INN,7c2MC/UW6S^DG44DNF-91?E5)(a/X4+NFV6XBMQ&:HYL6=N>
TSAU2A&0bS4_-L&=P<03/XN6^>A)O&WId]Y1?U^5K^B[^:(KTCbfQXg,((,32GX0
f)J#Lb4cGJ7b-9f7^P/g).:+Db\Id0::MDS=9Q@D-5T:bT:,Q<J_GZTBBZaT2K>+
17H?A2aKAdEH+K_\=28TfZ2=Hf-IF]ZA88Z/B[-0)GdGQU8H243/Lce)X_.PXYQI
I,PR6[aY@#[O]IH+ALf+J3YbbV;.WUDbSSBI1&+(Y=VN&fB\N,YI>-b8H^Ye/Jg6
GRIK2>3NNH0P;gN;f<VR99c:VXJG]eQeJb5N40[fcUdUKZ#6:BC9TPU7E)N4M</D
AVD^3,gM(8^>-5D69,R6Y/B^R<8A=M/J@4/V,[+^@DNSg/U4I5HWf63Ka9OC4YIY
T_M&bR:D,H@)H[Y6G&9APG[5K?61.&)\KN,gfeX3b:Y@PCDR<\;UHe9F3@H@<+=J
9\a>fdOZ^dc9>M2a,>RH4])TgY+G:<V),&AHcV51L^YfQdc4HOK.B[Z83]9(B?L4
gE5HE6FLS1D)8ANG6F0><]FGc(3<XV\^7MQ.L&.,_G2N85Z).?R3?P:/U7[6=?R_
IFL?,16T1+1[Cd]<IH]XI3^1+ab=RYA9HeC5B;#2JG#L2G/?./4O7T;>d0[QU7J6
c5.c0/?SB_1gAgIbFTQNa\U5dEJ?fN#S[eKLVII/92+c2<6P@T6bP67=X:I)/4(_
RTF?7W^[Y/^,gN?K2YLUR?d9B?,X3D27BY,9c)1#QfW0Uf+JeHDc(X8:T_1d>7G>
.8(XP0,<10=]3&^:3J_,)aFTN&PO.bUKW5aN1F#&LcMad=Y31KbL&\\:4F(RU+T]
]+]a?a#eR<Bb<P^BL7ZI(@6:83W[OgaKa+eHV-&#:QR9L]0^LdF[M)F/DI9G2&#M
?O;N0&Bb]?ULXbb.QXMZ)CA[ZHX_,<)RJO\;Z._2?V8@BSXB8P>3D7_MZAW#EFDJ
6#99>+:4Z5]0XgQ3<a&4<5[C@OM;=\+1VbD27)D[dDgf:2M58dV?<S1SFU+4[>T=
:U&FT^QY#Q8OcEf32<0P_:BQeRE+STL>^Ba>]I,,e7>D7+WL9a_eDcYI#&_084P>
?_,/b>M+^_^K8&9,PG_-M[#<NHURKNE]Y6=VK)fX]BBWMT9cQ67GW8AYX<UBYaF2
R)0-e<@1L@fHT[D,?dNZ#J>gQbb[S[]@Kc_TTP)bfXH,&Y,-dE/c[7#N0+5_9<)U
T#=Pac(<P)<V=G98e-FK6AE.]fe&e_ff2g]Seg/=3B.Q,F76.)FLO3,Rg1D=HP89
,+e.3e1UU6[g=N84>L-1;He933P#I]IeZ]G7\FL<YMM_1AQ0gS]4g2\LcZB<d<YP
#PY6Mcab9:)4^_2U3L2DgP[QLKTT(3bS]H1TS[[.c)M7A6C;\KV24fJ^B=;]+Z/&
0]B(&5Z;2g@]:W?BPHHGfb[1NA\+3/VV_,37J&(Y[J\X9Se\42QeC^Ob0[Q\XVFT
)I]P5T7)T/9V_?cB0P>Q2:B:N22,-P-T11_.D(<c+Wc/QL[ADcC&a-SHA+Ba#e+?
d]:QS=.I-+O&RdR/O&+E@_/eF)3\@.D(:c>d^UM.)4NG3SU)_OeWYU1Vg7@5M]EP
^T(H/_07d=ZHZ&8>gJA.K+OeLK5::6IK^N+0><+QQ^1J4JfdcD,G@X&c[P)9CZ,(
\b@?T<YKJN,7aM6TUE0=bYBQH1[?GUBBTE_J?]XK99V@3>C80ZS2(I:#Q+Zae22K
/f[DIRJCd7M5361fa0?96@1AOYg?NGdXGTW;9Z_UgT7UNGe++)efNGg6X@_KWR?-
1V]f7R;>4.TF7R-DADW@eM6V3eg(FbMW393@fVF7-gZM]Tf<U^=[ZG2,cdAH<@O^
#=(e5F=,KQ7=g/2fX)a?2SWTd24?8=N/e,QbFLHFX=AHYd4@O&)D95C[4SRGb#36
bNVCI4Of+GQ3(/MTO766IAJcYT]f^<UCDN>MHIEU?1<c54NK];cNO[M@37WT(Nf\
faX]FfD](L6=20H5ER1[e+cR,.:bc)gP8-OfZ+?1:2H.:[;1<-@LYfK@#NfK0G-6
^J[.J1+:49CF,CD[R6cgVT0g^1B1H8L2EXU9H-d6(I542f^K7&1,--TM3-F+4J0@
>H8GQ)QZ&e_(,>KO1;NeY-+d+VOE8aaDL)2CI/OJ-@-;Q:/)=E:\Vf0;\2Ie\SVd
/5D=5#PgTS1+#g21D9AUP[=6Z5M(3BS6I(K;&dO8I\;B8Z=IJMC9V&,:g^RIYFJ(
Z\\?#b:6COKb,=@L_T;f>fP\:fOJ/.gQ.#8B<RK1?@KO0<(De.X[gXea&D<ARg<A
aSQST@ZSHI2XIO#CY.>@.Uc-YCe<G[W27W+SM?>ggS39U_f\0YeAY:I(1^gPB.Y?
/.F&=1D^><URBg3VW;AO/4ZeWe^BQ5J5+Gb;/SB<Qg=6?93&fA/Z[(6F=aP7+X/O
7c.8+,/Q83>bNLTSZK]KR,PMS4<ae/^K;JAN,,@?+\?.>3&aPe60>FP5VEOc7.IS
^GUFf.O9?R]W7M[PJeOZX\,/gGPeR,M[QaYf4CKTd]gZdH?R=9TK\?ZP96]cP]OA
H9WdDT47GQ_-?M_(P[>gF9gI#<#Oc;9gOEMN_V?0BGZ1VaSd_J0b,D8P;9<^:>Ce
-PEadNMU#Z^;<UOMJ&(A)ONbR7fYb^4C3_;SMIRcHL;+4:9C97Gfe[C#VU8D[I3[
U?GKR@W&Q/-T7;E>Y?-]>=&8;^8(@AQU8(;=2b]K#?7BY9IN/C@Q0;>,#fA>e3<Z
=Qf28>bXc-aLMS0Lf4(a_JG_7Z=-T3A86VG)KM;P_T7L^d)QbHIMUU1af3:^Y&,D
8+M<c1+f&:c#WAGF=V\YG&KO<>JHT..,CgR1e+X>d7gEKT^ae@VI;P5Q@60RXg&b
AGg5?7/EOSbc0UaT9dSXIHVTd#/Q5./XE/+LSVO5O,Tb^^<CeT?4^;d:&<P=[7G=
;9bL<c9Hd3G?TaU2M)D&Z7<9X(@AcdIYB)_a,R^3QLDe)Eb>KU2<TK[C;;3)?K_U
fRUT1^A^==)VN4Ga^IfR2@7O2cY4S)VCS5Kdf,]^7a.+0d/817DNde/NYP-.-Z11
A[),BOU@EP?_JPf.aADAc-6+BU)ALX:-V0PbX(eP3>2RKedPdU_(P5^4a5&8/?c-
]X4JS2L&Uc5B@_)XOcONXV5K.cML27._a#UOB8#2Wc0RB$
`endprotected


//vcs_lic_vip_protect
  `protected
>YAQA\2TV]DLX6&UXbOGT]<,R;E2:4f@R;S6M[]YBZE4/JMW=CY@,(+)8_fP-=[d
<R(M0fgbU;fFKL5_bdA,OK]fK3Af07Qd7LR+\,MELGNQcXT8^^]WV(U-_[aT<JBN
+TV#Q]U>F[(@[OK;79\O=fD7AZ1-eP?O)]&9#CD;G;Z/^Y>bD#P6G:bH983MYSc6
X<IBUCK+7QJX=\\)W8=,<]^RYgB]DB+fZePfV1-2gS\XeX>GD.a^3\9S4.5/O_[X
DOb#2Rd2^JeBe-B[444:BL]7f[>+TY,PVJGY@G[6+cQRDF[a>S?>E=N<QNJ.ff+;
U[e5B37e:Na-O&JN=bS(G0[^M3MU46#BXW-aM?E5McDRH_5AOE&[a41eU42]g]CX
2&\<fIga,H[1(\UZB:M&,f#(SU7EVD0F#]e/:bdB-VOD26<N-+4dJUf?ScHZ7Tc/
UW47/b.UYdc?d]b/;T)0V/]+fYQ15OKL^7eN0G/g:9U,/9<]f)d0_.41R[[/ZCE7
J]QH&Kb#6R9;f9Ff+aT_0W]76^=,+<L^dOaDRO^JGHGG8KX.23@C[fe7]WGW,[CY
QP(=PPNa)@TcfL<^+Z00S\Y<EZC4:W(/4ROCI1fOQ@2097G=,0119LG16+A8@Z9V
c#SF48DWW?D(Yc7F8N2:_eZfE9Hg;J5\+fGAZf6RJY0(7?504KWAb3Cb;US;4MUF
7N__a^KbD0-Mb7<PHD7@F5N3CE)DeM^N^LH_]BQ]B((OcQ9SYPGV3(Yc^I,73F,<
)@,.)cXDgI@=MUULLeAK=/]1W/;Yga(DOI_b_.9R#9[L.Ff4Y,&3cGIB]AIFX5c,
f:Y_1I4,dgXPU<c[1Rd:NCO+UF>5Ae:5gA=K^-d(?#^\OZ-@TAP;,f493/1>X.-Y
AN]GC_;,[9Ng4593RG@<ZQA#DD8VN48B@8EbCI\4fAOSH4G2QTe[I5@O:TW]f\#L
Zdbd#T_;:>gOVCNT4g#1ZeU[USJM#;E:(\fU.SAEgMX0(WK#G2#PP?A/22?;R\\^
+5X_-@+G^4[92+EG]e^ZTV1)Hb<#,=ZJI2F4-YFEW&+@c#_QL_-6VTVb?LLdXd8=
#e8EC_dI_6UTM7E_JLOFJ3fITPYW#3b1&JD5>O,C00>Bd3LT3?T=[YbJ:YDg,U)#
Z=K5S:RH45-a2]=D>+2dSJ165D9Z[&<Cc3,0=^FI.?4?NO[YA^M8gd^;^5DC)(bW
3<S\=G@,HVA/Q_/B,,(09Z][ZT>&EHab_^3MEU7gMM7&#,0V,:AQ1..dC;?E.MKe
8]SRY_SOS+gI<V?GId4PfPA1-3.LdWU_fR6@0J,B@Fb;[_DdNZN)dG>WJ(Kf@SYb
7GH37BLEfQ?=+T)ba0_BE(;#d#56RGPCbY3gEX9fN.TTAN>If]ZdYZ7IaS9B5PD9
PIMZ+\=9>)>0Faf#<?Y]S38Y]>7aB#/8DB27?FD0TJ@<:;@<GgbB;@OXLVN@5U;0
_[L^9I@K;^R#7Uf.daCX7G?HHEXO8<P#TN(]T,#7Ie]OQXR.DSLDSVPM/-8XPBO_
.\Q\;;Ag).F^Jb4[-46+:IP>G0IB93OTFR?JKLKeOaWeQ;6SP5+^[bMTI=\H1AX>
5dIa=(NUe_X\-/U]F^]F0]TE5UU=HZ<];E,S/>^fGJ@9@dFb<7N,OSHe:e:cD1C4
PSLJ[#dC_-?QZ[@89@KFP+FZX4Y5c&a7<#0eT+YY?f9_1K40W2DB6<c.,MQd[0e/
g]SJaH-V;M3_\I:JgM@@U,N.]@3VO[F#C=E9-I[TG+X)fJUR^X4_V^>A^^UFA&10
:M_I:8H1ZP/Y#B1OcAfQBVX7)48#aHS:b?FR@<gZSM8M;KX5K?8b(_bGE@CR\c:L
+95cF=N^SB_J(/7/_WR#(GZZHdL7/7KHa+d/WFUfeNP:+X7g6ZGDM<2?-I=QMA<R
e6<\9C?G11#C2Xe?dH_P\<S=B&++@_IgMF+1Ce:e0)+TbFbC6X:,PB2PO0Vg://4
0,<J2IC[S=PKYUJS&COC5_gK-3(3b(IOD6Z#HdaGQf<;P4^B7+?#\X9Z=VWZ0g5E
+f>g&&2]YHX@O)ZY>E;[YEI[?O@?<4I-;OA+@ONJ6cED\7W^AR.NI04D6?T>/3Z2
bS]?d)cG9UeI^P->PI8NH]7-;^10B^=7Z9=7c63a^]5d^7XKY]#0.FfeZ-)&JO91
Ea^RD/DKJD)^=<-YW9Ne7PQ^G0^H5g1W68Q<Y8JFeN8,)g^WH/&JN<MK-]/G==EI
KY0de/?J3c2@e:]=G)4X3I7gF-Me&:3RFSLa]eWD7N@?\e/E_Zb_#C35UZ[>F/9X
T5307=fAd(LUQ)eTYc[QW7a\GC,\1>_9TNZQHL\6:)PYOU,F.3eR.D/?4NAKI^03
L6Hgd;a?gM,b6-C+LIDAPJ;6E-/]5V[/#XL7UTD\QcC[K..DZUSX7c=^5^gT80@5
/[Z2N8gJJgd^Rb9+)9V>-P7?536EH##66+\J[0C^0]VI3[OKP\Xb:.Q&LHXYSR_4
@XQ>3N2Q\6^.gGZCR[gOO?I\R-YN^>-F:BI5ECMV3dM#X=5HNS6>HfY+KQUb)&]+
ZGY?X(&4gUNJW6O-1B[Jc[O<+6,d<\MHfUgg;5/U[T>HS-U<Sa&df6W\VM[IB/]R
A]I=@M=Z#&RJF#Sfc)L9-Z9](&A.#9TT6Z8L2aHN@X5@de4D]8CR[<K7H,<Q/c2g
DLP:181Z;>a:6:@WN\XVaWK7Y=N0).T\V0O6W=8fU+.N_V2,N\PZ:Z6PFXWY<@,.
;FM6^1SC[-fJ_.6EFPKf(^f#b?,(W/,\+_YOf;D?=4Ke&_G/P84>Wb9O.VbDGFcW
6(g>=4)E@D2XN9,X;Q2E-_KK+)LJ9dSG-3??6J8FMgH8,e44G2TJKT<eGM]SVAJ2
/S7O8/8&IT@IB,E]8TPC88&.JbWf:67U<5J1ceY&.G#&(QgPUB2ca(6V8eabdgg.
edA=Z:bW8GYH_#N##B5)>\5Y3PC51-f@gS<6&S-1J(IQa0:,69VP@SbRGa+V#-JE
.G4Dd4?YfZTYZFTN.Z)@RF4e64]T1,X[(XOe@;CS\FM:-Oee]L@-7eOW=BVWUS(W
+DGA(6]^(I]c]aXD(>f>e1B,I[7J)QH35VdYA0E^?B/4e-NN^CUaVD_?a.1/ZeTK
=^Y)B+]Ed(F+,,[3C2=.=Z_;]==,>:1e&^-MDaM;c6f3dWNVEPK+BPC^AeC_@MSR
CT#8R/GD1(S2C3PT9,I]9?MAOE[VHC4W#1]=129:TF5^8>9edfHZ)CUf4B(aN[/L
ePG+gd)B#2eX1+AWJ/:NBQSe<.ICD\,P?HK1Y<]KMaFe?MF27#5\3DF=OJYKX-W;
<+>NZY-<OZF9F78:+9[dDX=M80_g4d/GGK+>cM@+.2Jf\WbHg/f5<B^^U4#.c9NJ
4,_HUK68,9PQ&ILXV>41H\c6O(b++RZcEY0<XVH:YgZ&&fgF>J8,<E.,ETRPOa[(
aHRSL^W#8]WP4K0MeGJIf_SUg]^T-?E#d?YBY=;gK3/)c]](LNJ(^CP^f8ZN>7FM
,ROST=5CFT>TYdM53-f;PGbg4V@U]O<8#&]]UV))C[f2V(RH+6D918V3;.dQ[OIX
dO)P]WT]4gHcf8H=75W3.X1ZbZ=Q;LP,cSV?&cUD2/3+ZP<V6K7D0&]#7RG]O;3]
(GY3BOa:@]Y)eb8CZd>GU;.C[ZO#UNFWH+4AId<#[M0D60UEV0VaHYR(K^K,d\5e
.VZeWUX2(9;Bd#gR]=V=aa?H&=)UEX4=Y4:)[a)?T;G4C:,;),F-6^d]a/]<.WYA
DPNEL#B\#:c(eDGDPf8=J.aQICUSTd1a@QDf3Eg:dgO>Q\aF22>&fB+:GNS_-E^6
8YbdOYU>79Q&)?1ID[M4-3KbPcdMXHb^c/Y^AXTF)49UfKI357BF.f#0H<2QOB?f
8]#><IYL\T>K<@eUd)V].TTUY=;5_3]W30JJd<^GO_&-].fKX?PeY]=I.&G56gB&
C3X6F>)B3Wc1>b\FMX&P^TD1fVZ.PYB_Rea7QXO3;@T[<[H(9RJ]^VTeUaCFANM/
-A[J/7M3bcK;B7C&BfDGNM<\RH;K9)7a70gT+fC6R&P8-K7>3<8YA7O+&LH_]H3H
7&F@>.dfS<\7&Y/,+J4F\_#(@;O6;cW7#]dP0?C/L7dQ_@8N.JgQfP00/c-<9/-d
1c6.+#G,K@Lg8\JK>NdFPMM=a(F,MNYJ\beba^A8V+#T]X=>I6[4O=H2<AT+QWgB
_B3CeY7]-]DP&FJcSO/@B<(aa#P@POXJa:QIeF8/O]?BBb<1Hc/c+-cVZAXK+3T;
8=c3@)F3bX/W]:I2O4UGLG?_DRWU+//?-Y9VP9N,E)^(R,)c=QBBeCP:L;a.2TId
TV;RQ\1F(GDJ:7AORW<Q&T@L.0VP-P6=)F#&TDb\Pfg#a&GX_Q5O)Y-;VJ6TKgAC
M,/6)E0D;O27P\L),DYf,0BAOW^+NWR+8FEH>U.I6\272D+N(Xf)-5]E@/@eP.Qb
&C0N,+(=_\\R)TSTQP_a(.-:NaUUP7RZP(D^GGeO.(,1a4-8Lc[Qf@g2;=CHKRB]
K<>Z;d>RK=1H=YR+PIeL&8B7(H)4GN0(GBa6Y<A[(79XB[9Rc-#H#H-.ULA>6d;e
I]RC;9a)b,6/5/E.,47#<EQWAY^=ZN69&A-8_\ND9QV.1J@ZUb/2aQO6.1fQ;NK[
N,]/?U;BgKg=[CN.0,S-PUBCe[8\c(<)[NKR+0Z^^6A9aU;;_GN)5#.]+&9.[aIO
DL.ZQES<8,d]=HaPXWF.RA=?Y<c>)8^&,ad_5:NQ)KOeMeSM<#@IEOJd#JF<\H0E
,E/#2XeAGb^+QH;ZBVDe^9;R=M(Z<e1]KIL,7a_7g<3gZ-ZJ@?]\e?GW-+K9[c^&
-BF@^(V1.NR5F2W/,T,4]R>;,@)K=T9/FcB4#R)YE_4;KPE->f^T/#5SX8c:O2]D
/K-g>d66UUF7L3LS6N0:O7:B@IFF3CT5..=3Q&&<,18G,QJE<RNfPY5Lbg\<3[+7
UOCIR6@IfLgbFIGJ=-?LLO_K3?030bcC6_?GK?&IU-ARKIY9Ge\32DaG7Q<R+Zeb
0-B0edS/7\3Y-W-+I>9OHP^4XGFSNDRf/6ZIKWK.STG^;>2,.S]HF^:f1Cc[:,0#
5=TA2SLMY/gW/:B1Y7c4d)A-N:=AB6W(DL-d4,a]WN79]JfB5.6I:EZJX2Z-I9W6
S>I_GOL,,W&-+#fD/ALAcAOQ^SMMCB-ZW5N5XgcICSV>IG#LSR[MT:37AJ.PTaQ.
]-RH(#_?61<GT?L/F&JFJQISID#N#a(2,M5[J8<?QL3A=&LgQED#Kd6@P+(B,<N[
=CNKVRA5K=<2L5g)I0D1,W:I]M&+V0SL+:APSH#(\TaAOW;W=^G/NAccMJ4(.Z/Q
CUQ;Da\1Q2YLT:;C7GA;Ha6TER,)#_^TE@25QU:#?9&IW41DF-:T>5A2H@[OU_5.
H5C-L]>d79,?X73/GOC#@<#=D>?dD6Vb&2-(IQNIVL;0D&,?9V[dHPC/(gR]<YZ6
a2(-(8a/2c2W/SFKd@@&,US^WT,(5EJ^(3g1EUV\)eO]gf4RWK].HINNT:VDaJ6X
Sdf?IQVbBNSTI?4JG0?LQ]=3W,J59\?X+6FeW@KQIP7UIYVT.7?<.PYVCKOO=H[N
=3TP(Ja79d)b2\>HMJ?aRS[]F^J^1-GI&/:^W:#&OM?b&@ggO]A@ETC/MVD5Z(H0
#O7RH/U6CW71YE>]20B3/7YQS_[#ZYa#KU;3T6^&dbQ\S+fITfeM]URI@[SS)CR>
g@N&WRcZGPQ-ZUg++IIa?R[;#6aSUAE1UFLfW<Rb5NK-T6YF(_@2b3:1cNV3\_Q7
I[/;<SWdD-=Z@RPZNF?URc^W0G/3fLM;(:R<)YK5C5Xb\\&3;;Cg@M&DR(6?#.5>
WcH&d4g4#/EZgJ@Aa0PNc,?/M?9K4b+8I]c#df9;_Y_.D6^.fY\3@X^&).g,?L>9
Sd:dVTFaO(H\ZF94UB=U6IL&FgEe\T8?@.]Y?+4>+eAc23+dU&FWNOP+(IdX4_=Y
QTaa1,Xg5a^W7(M622CXH49-9,&[(G\4)L_M0?]N\-&4)Z-H-1BBTU1M?VWB6QMZ
IXH12T/A#2D1EP<R^<ZI^,/LUG4P;&F_T73GE.EObNEaG8U9eI\6;H;)3=.7V_[9
fQdfKKIAHc[d,W;fe_LL@9BO52T2Ce_&<;Wf(1MJf_=c]S)1f^+M5B<JU>H==0X?
[(QbO:,GS[LTM(NU0AZ:71MW]XSREB7UcH8af/0JD0Q)9W^b6>E;a8YDKT,2O&d]
bg/2f/K.PdF8\5RAVeRWVE]OPO)/\3VMd6;QIHORQE>/_<Z95YVTN0\@ec2):/KV
&4XY8931-W6a68ACbf@)&a&9?bSfIeKgNG_bZQ.KgH(D7Id/GW@??L^29-b0PK3>
;HS,,@A&3+/da)A+8;A&ACH1SK\;_8?FFeN&>6;#/1WScDN_12VF2e;\V^\S#fXW
]gR#>A>K\Y+>=57@.G&YG>/O?8NeIZ2_>2?5D16@9HM<_T2A:MX3CdR2d4&HD?SW
D^/cY/269C;5D?I;;HAgeZT82BNMTN9/@I[;,>dXJ2S)1^E73bBN]EGGM;?(]\:>
YIJ&MRCK(.@UXIZ:afOHZI6==WS86(+_D9/M&YPPA>(^3>B1YUG7X8I:^,9YF.cK
/(CUb>gKPGC/2gTPa9FASe.]TPZ[e<ReHO@?)e<8_RH?cAX1)2ASL4K0IV)cJ.)?
g94KP(^UC.f#Vab>>:E[7S1,(?UJ7KB,c;Z]N6:O1E)@A_;)61@NQc9=]Z@K=K:O
2cCR8ZFc_]PVVCB@QM_R2IXN4<5\06&CBD5WGEUc;/;/]IIR,P^dVOaXaGc:Z=/(
SZf)]3O9-AU>0,_S7[Ze7/\AaB)[8SZ]S(IW/>P:@O^P7a>SN.JHT@.6^cPM[G^4
OX.gF0QN#fUX9K,MO0MI],-/YH;H5MbJEI]FDWO:c;&H=Hgc.LK]gYDR(GULf^3?
<VP-(U<>VNBd/,N.]/C,Q#-/Q#^2e=6gVI3>/C>6.Te96]J\@<9KY^C2D9>AK1<\
>;cV:P0)_8=F#?I2L(+)EL.6UGVHZYe^(J#=M#_4>E)aH_S]YcWC[e+,MIe..d6c
5;:[AO4cC8H<@PJX1T2a[0=f5+TeRbM]g8?fUgK][RQR1feU+b,9.>c.64:^da[L
L/N&[gJ(,&ZA:g=bSYaK0M/8)aBK9gF=-(>Xa;^9bD#IHS8W?Hb#7>cceBS-&2[3
7gYg6#@;(P#][/>)]S\[?,H#EK6QVQ1b3D?Z8U8OL?,B/F2TRQd(T+HPGTGD:#b(
X<Z?.Ed^VB]U@@>_3TWX6V1dW\R>PDK73U=WZb8W@)@Fg/gVGWdQC)M6a:;>\V+,
B2^PPY/W<BVa7:=Lf<ZKU7[G3,5\_M8+L?/Q0&#W;B(53L^H?2g[\geLS&e_/HP5
(IK7XY@>T+JBYJJfD09Q)1PDO0^_724]-_Y4f_N)C-#I]CNRH9VN[(]e3-6MB-1R
Oea,R@2&I^U/>CK6134@#P(/:b5JUYO3#@O)@<U>LJ0YOSO,CBE3@?4ObUD9g]e4
1((&Q77\aFW[#<FS@/5NOB(>M@-Ig\GGFH;NJfYI_5NT;S_8C7Dc6/9A:VX,F(Z+
]UV)3)B.bZB/:g(-Ke_Yad7/INT&c#216NF#KXeMU1UM6KS#R9^f7Fcg0G/H9aJV
UU=PK8\(NKgIf8-(#&^c1F\OA&/CH1+<<3c2J65bOW&.Z9.@>ZPg:?;4XK+44/))
Z5TE1QPG+Ib5_&T9.+QU\\T9dATKgN-#E<)CI/\gc/PH<]V0=UKO?(g7O,fA@RMK
5W:GDIa.Z:0F3AeY_@ZAL&7bX=4XWI#OOK&-LZ0eP;2JBV.\1?I;>PdP7)([b_bf
;&U)1&LJ>Qg?;\YK/HRKe952XKE<3OM,\U+?5U0>O(:b@#=>\@YZbBHeY+&.X:b<
-6N;geSWHeV#^X=J2PXDIN95R<V].Q)X0K4C]S4Jg9)c]((?,@C@&e5_3#>]D[;P
K7&GdL\\J<ETYe&I7RTSU6LLU>CLVH=G+?#19K=26d[]UEJ12dM3T-5=V1a?a0)L
]X5FC4d_[AeW+[GYF5(Zfed\::D/,:.W_N7Y,1;^7T\Yf]CAG:34U?J(f?X7H7UP
LK4,,N]/Rbgc2L?Zd)?2&1ZFYY^RG/A9cKDRecE;6CD1JK>:W),7QGXLbQb#LM9&
dO8c\),H@2-b0d&0OBELLGKP=,<R6)_VF[?EHS<Q1BcBRZ-b[2P\?1NT(V\J\RTW
UOU)=)KdNSTd;J@,WW6J:;ab9X.4Y3DR9/6aJ5<:/<)6&EFbg?f@=CTIb55?ZEgc
aa<CHRX:I=91_H-;LF\L9(1c3D#P)B(:8WgTPS[\+IF4U7X&\IEW=;-aY=W_Z[Q?
ZVEGXReXIFP>]e#LVObYfB7MNFd8JeEdWIZ#E7,09U:.4@@B3^bTWWD#7RbB]C5A
<QRfbJMW^U&1/CSaX-1g-:4<HSWZ/dRS<L8f+,@,gTT6Ae6E:deegaEJUK)23eX[
YU2-ZG87#RH[BB11R80fPRDT3/)G3K\WLU,NXO5)X8H6S\>NY?e<A7ZI(dV7.#RC
OPP8L1)+P?1Q#Vb]eP])+:-Y8f4c1-T9S=fg[L=]2QUN8^N7cG\aCUeJI8IAP,J3
a23GEE,)>>+)K9DfNKY:(6MVVROL2cJAC#B>R#,-NTU;W_GLQ>BD-V2b0Y1_g=>Y
(G73:#73SGA\S,b#\FD(#g:35_B7=bC\O?+A+Z=9c50H8?dJCAH-fIgKY1UXaKR=
&95OB_(<YeQaZ)6<.T7d89bLWX<ZUY3W10B[23Ldc+2XIW#[06P#d\;44a1>Lb(G
GE[,^=R]NA^X6ET@<7N)3BO,V&U7_2YK9V#^\FDg(<:[?5:d.E=#Na[bZ,X?Xgd9
W86IX&Z,NEM,2aHOJ@^W8gAd(/54[dW=+JS(cCA=#3OX0_#MS<89NJW?KJ8d<7.=
IJ&:U+0#+BQfZGTKJA>.^A#Y+b>O<)^a&V-R0.97PDK?BW+7>U_EfH,#3,a;-XY(
2KbOE=J1;Y36S3(F(A58.Z3EU8Hg,3G+Yg3^N_Re<e=@a/Z_G3VB&Q8#HK&PaGTe
>F_ETE3OJT#&V>ZE.-15J>&-aF]dPQa+36bg15eeD65f6TW[CJ&]_3cg9WL__7Oa
aObAB@GL=8bdF4W(V7_OM2e,g[\BFJ.-_]=V]+8(<P)]bMV<WJWbVCcDXQWgAW]Z
MH3TQMP-4QMF&.Ma)O.#OEa.aC4_>G7N/]H;cB<d9_O.YOHg:)R6G&A&;+JQ)]7U
7&9MfVFc1OH=C]PXM38fJZ+&DFHga7(076df212)Z\+3BUZ0U7=^Z5<_feVc+8J_
V\7#8?Ra4&&\,9G0;\&CF^a,3g8[86D<+YM)e)BGO24G:=-,aB=)RP&dA?[49D:X
#Fa2+IMf&(5Q#8,)dVD>DE,gQ1g1<2d&HRCcG#@[D41,^0)#UO49\V[(TRgX0CAV
W:Z16cYNW8g\]UM8YQff)U\/Ra()H1ES<\f4=LVe41^H-L?@:?aO/AF1O+Z#[L[e
A]<bAgf(,#VN=D@A(T1GXUb#4HE+OI^?4IO:+>D4Qa@M6BNPdWO4XQM=aa/^Y\cQ
>5\8M6(a)/#<G6>HMO;5C]3^/O;U-:9FWBDU@&Q+89U;Z#g>S:9[@2gI7XO#dXZf
1K3)8O<7.?[0)L7^W#CD-ZU_L\@/)OTCUAQ9XBG-G4&+#M)G5B5K@_;L^OLGHbVM
8c2B]@KKD;5bS:8OGK\S60,+KD8T^fQ7)\8?N2GeLA68.1WPXcaXXc,]/Y1NRPKU
>X(&.5XIb12J.GWf,1KTeZB,2#SKT[<<^)FBAZ&+UN.<L/O]OGC#DA=MM#V+)9UO
:Q0ed+#S8dKg3L=>]#UAHR;:_:dQ^gCc]7]AK&TYEQ0e\fV3H2:S1#aSWa3.P:ZH
27XYHQ7eDG(AQ2I=bA5_/8]7I>,4d>(;9J6])Q?egV=;14S3-V.<-.L,X3eCRZM1
OH3\LI8FR#QP(dfP+(SDFLeMLX2ITQZX?NA6XGAHVCF):5U=e[LS[Pe#1E)02b2Z
QWG3^09N-Y44XRRQ&-M\.IHI)ZX1aV&+=OFGag.TUJ\=](2#LW>VK6M.e34_,#H_
Q-+;b=DZ_1XgW(D#@R@TfBC(RNN1/CC@LJSDM[f4=eS@B_+[N?9FK_aM0E0+Pe6(
e.^KX(?UPL)SEa<d\NCcA:6)-C7H<,DR?b.;4#UQb:7E_QXNaGBXFRX\T#4X3/<E
,HRPWa()6X4MPdK]6S9#9+MZB?J@I)FY=_:,HPSK0VH=Uf-2.?=4<d#[,0(7]TH,
Rg80f,C(IVA#1;Ig6\J6D^G#RYTO[HLG:/4-0O+]--;9V<W2(P]<6Z#\]W#?:dDS
B2T3^H.(]Sb4AaSX&ePJ>5T/FWKF#gI@dVcJXY+RS^g-X]:)Ld2/?C9)dM>aUKL,
#[_UVYCX7da)gT1QQUdc4NGE+>LTQS([[CMA7;QT;b6:+bZ)1@J-K<7R?)9#?D(f
N4RU-Y@@MD0<SC]7dNg;QO]W]\deG+4-B(3#XX1(1\UGKL()8YJEGY+QB)D&<WB/
gG?:5bN_&RRY;N,d_H^FfVAeUC2L4&gJJC8\K=P&L3&T&SXGaW4dD,FKC))DR+7,
dIdggIT4-&JQ5P]7UT#K)3-FW=D3@[.1<c0=Ec3f2OB@O:M#+#R\YGF#JaFE0([B
6_K[ZO3?RF5YH8WNJFdb8Xg1E->#>gH+6PDcaR9<=:f(5UR70VT9QGU3]913#g@^
#<cA-&R1>b#:a-,Q+a+IXaHeJ/>@.T#a,0Z=8:>.&ZI#b2-(#8N?T-WJ/]g)Ha/;
-<IX.I,3bE>==ENeG72F:XL)BK],E7.DS<G?[2:QKCV5BW5FA3ZP0c&6Fd(Z+?SA
1BX0EJ1:=J6a#NceeQ@,(XKe6M5N)OPJeU0RLE2ILV\_1@3@>@Ea_aaWN.)@GUYc
0bAWZKeR4&(gD4fXF#1IBg+;AOP6Z<E4NP5e43D7H\DTK,QP#<23ZB^a3<5Z+PX+
;L:e-69P_\4II;f_KXOV.Td0KYT^M0EH\3RVD54QOc4V9<E43=Q7_/K1B1MU\(dM
)OUH88P,S>7U:?3IJO9:eAGZYH9JTQ@O\7d3K\6(KSEdSc\BM7fRF7G_;]6dWeOJ
X<4)bF2O,f9NXCced9LGJ\_Ob(dRVMMVOJXI>U#S^/_0aef14aM.OCPWa.)#0-B5
@5b)U0aUU.-3/4XagXT_14Y2AE1D,Rg2/LBU+)N7L7&5]#bY?O^Ve\a:J,)a;+BM
G:L[C8U7Hge#A3MPg>#RLU&D>Y3@ERfM]V^.-)R(c:+8QS7,9Y0O6&=:S).-d/1Z
a)2>-MTOGKOWP8eWB0_1gZW,.+>-?deGKd\L@.E(FB-\-\.#H^7LfG<1V2[(VH[c
+@?ZUR8,#G-Ze[&[_-Z#B/?LE^df[Q-=@VV<Q4Z;11/#_Q2+BfZR(L>^QE#,-J,C
&A6OSH#7d4I#&O0)T#<@\,LLYF5,])21N_5@c-6W&&X3:8/AS]E19;Z/b>Z:_N\,
>d-^^_TEeN[HSfG&-.SJ&=YX/7J=/^]G((I9EV6bK=c(N:gQP0_8>3+M[(M2])A,
\Z;ReV;XI&AV4,;g.9GD5@NT:b37NY.)#Cg[/dW3f?<4HZc65HW<B+T6YUX_8,.c
b#\G6D0P_AF<X^:E)QBF(W1S4@/EdTXN&:EgCaEF[IKYWGPTBC]cNVYKQH<FfIJd
e7+b#)SIb^Hdd?5K^VUd>\0=FIcaEO\LT8+Q+</[,2LJUTPG;6NTA<.)(-a&>]JW
a4b/C<0H3P@67/,[+:MSZ:YOCaI3L<S4c;6d7H7.==WXWBe1Qa?_?/I(B:D.:cK.
Y9,_T3g)2V74NgK@GSK^fIN2]3#R1G^+SZ_b2+fIA4=E^DVfMYQR.M[F29,J7cgN
9P/AYbN5;^LX+M)fZI(a);.WMGa\B5^F4@MecUJa-+-EJOTJdGgQX(<>(eZ<f<E^
9>85FTUCeW/7CL;g26g<>L1IU;<X3?NL]X[+7/R\S-&YA]W79fNOc+-9ZI4<#XUJ
_1EU^\_6W@O_/NZ3(40\_2WecK4P25]9g\1S4HDGg@baHB4&J62=R.E&&9P-HO.S
KXGe9;0#GW[+)#X&CC32ZcQKe^)E;CgX0?A_+H1BVO1#4],HfDR)JPa==.I-[V2f
E^XWaVU]J0C#.R<W192N;a^M078,c<4@,O;LU-.ZS1/RB.b9Ec4<8XdRfB23\H)E
)Y>U.K(^/dH#1Sc.gA6=<<_6/DN(#eU>#NO03.Z&9:\\7V#J)BE-ad[6Z_#_dPB1
0<f-65V\8W\--fSF\O05Q^gDMc@[JXeP-22)cJ\7R?LVA4J2#3SG91]3Z0f67.(I
PG9SL,>:>XEFN:683b<CXH8:<BOFAd,1NdbGU84G#_9MP\4#D<H^ZbT+YDBB_J4J
aS2c6MPT0)E^\HKa8SU>YNEB<^_UC27\<9ANO:Ld+UC]]=5P.MT6W9DOM2LO)_XZ
O5;?D^\]&F//PI/I[<)@8ZH)_d.]bg1Q]:B>.a9:_UI&JX=L^BW71b1P[Qd#8XGR
XE6JB9,6)V=KB,G_T)9@ScFVd.C?[:G@gf7/ABW#Y@7\f_A3V<2a(,7@g[C1TWa1
CfWROFd4B#He@MR56[gCCENF0C8X1d4S#eR-HFQHIdGO6BXUFbW1R4@>[K\OC3X4
H2JD)(bPK^?87/I[b<NY+\VV6LJbbX@&(>6H&<+(7QKO6aC>,7OcT[4[,J:#HFFK
XS/ZY(_Z,MUf/E?/cZ]EA5@fC@cS^P)-39cR4AdJTU_D@[1.Z>/?K)Xa\./3)_./
A08PY[7^C.?J?\(3gNc=)U:H:]H/^b@15/P=3?,+&fZc3b^O]X37CH,e:9dM98,d
NT]+B=3a7N22@Q7=1X8bWRKU6g[,MPUD1G<NfQ1)1N5Nc\Q#U>64]LN87K-YYdF)
=2<f[Je5,O2.dZ_B.Se_f<f#;3B&RAULdffcEI0-AQ;,2V^LGD<^QG1DK(1)<8/&
7)SE.WeA>B(&^Gd1Y?2<HW5\V/bcY&3FJZdK0MSOb(4B3eK_W7]L\0VA>)Qb8S99
8.5d3O,30IE8_H-POX4gGIJD0PD26@4^\0K4[+_W2Me[bKNXQ;I@E&d@&G[I,2\a
/d:Hg__6>LF5)Z&XV-2QWDCA1@SfWMc5U_L@aB<_X3g(,Dg+LNX(ZP&3CN(0OAR=
,2T]?\J<G5d[E:XQW9006I^VeggK,IJ_A_HGA9NgSO20McF_?,UM-YV5<C++/Lb5
MS\HPD58;N-B,EB2Y<BV42F@<A4MD,I<<DPEa1@_D,QYZ-bOCfcRNSd7;abP/^TX
d;2-@C_B;PG@F<:OU32=>X>EYG_UR+f17f405-CN0b?40JK7;5@)+4FUFB1]PWBU
cV<ESG)MZA;.gW>V=NM#N=AcW_M4+VT[NKf:#UAYadYTVGLEK^&MFdA,[#MaWPFZ
9J9UV+I(Zd,M8=JX@=-&4&K,cUENdAG5=?@6D9g-LaMR-WW=_eG>5I6#&a:IaYNF
0A,Y8+:I2g,F^O1@)I2KAbZNIbcgF&:EE.3T9R19M#QJRT\NPZ/V,=gK@F)?gFM[
ZA7CIXCY\FM&bTCdE)a2bf47gBNMEMCM52_T137-\M)M9Qegd79gI@=UUKN@))c/
b0ACTV)[+EZaAfG0/gZ1L9WA2B<3TYd;=-3;5DIbeZ/O2-#JC;O6f]1ESD)D#PYc
+B/K#f(ZE.=[#Q_H7ReI2@70EL(V;\dP,NQJaZ7H=94@I:^UbDe#)7M]WGWWgRD#
VIBWf84]5,X.(EdG+Xa;OHb0DQ<,[Xa-]7GbO(R5U+d-\?(-]8P/Y7fN7BA81g-Y
5-aZI25J]:O.XHa?<Ag&#Z);T@,\F(25.-;#PS=ORg<)H?7?+K]5?1b1K_>0[9U3
L6VfS(Q#@U#I=0eFWaQggX.Of_QD\:d&a[@3BP9ee=A#5;FcFPS<g137OPNIQ@5M
XSHRAD^Q@HG=QV[9;K\R54OC)\H\75(b>ZN>G>/+GZA\]P03K5A)02M(A5^KNZe@
WPN/(NcEB6MbB;Z_>@9a:VQX(CQRdWO_4^X+=T5&WXC.LVX3aH)^E)P0H<>(=C^W
aYe+VS;5-VFf)&LY3N@[ACPJ0USI8L13<ZO,LJAcG+M+FT=ZV>4N5U+^YCU5A_@4
SVCP_]L._3fAPb#OG#eV=DJ\S\5F^:U)aVIP>QXM+I[,BK/-=.\TGE^WeN^g5WbJ
K9OAEDUQZWJ?QcY&3N]Se\bU<0\eIX@1H&9M3Y1/?]/(>a/#1Z605#FN-P)WRd0X
(+S&(:#NDKf,Z^:VJ\O:Cb+K:&J1ZPM]G\[<3>#UHIH?GCYKCP.a#Ld/KZS3e5T6
OId,Q_@I:-](=YI9aEeRDW#+R2V:<O]ISP0)(+.f=<]29d8]9>JWN.g_,XeA0+CP
aPX1BJSJ=4#]F&U#6./;(L]7/>MS(bIU4dR3/\H?M@;VF3S@)3#MQ^\6?Q5Wg[PF
,5gF42K4@U)8M2^.6PXa9F;)b^e0]fRGSSALZ.5RSQ-aB4;##BR9a=:Z9CRU9G5(
DNY7B.VbLI#3:G5GY[)]RB4,#OT_P7:O?3,^WdaD,TNX.d:,SgHf)7??H<M@7^9F
N?[ZDL/?I.8beJ8^1MeD^.cD+LTYf.WCCDdAYSMcDNOIYUc16E>O]6;-&>8?#7bB
=0[:9TW@\8PFe8:,f8=WLV/-J0ZG>;M<0>G8RBP/O:_=/U1[de@.<O7WQEY(^MR]
)G]&N&=:MZM29#V6T.gf4dg8A0LH6-_HNSX?4([7/a@QXL[QHc#H)NLOP-b26?T6
>3KOIYbH.(1M4PdG=14_M1#@RaGB3,d8(D/>66RR41SL_N)ec-6R;&L5QA@a#<,Q
V:X0J=8g->,f&@+6B/PBb/3aI0=P7)1GF\?ZUYC2I50L(#\7CKFA8BEga->[1E6X
DgNTSNS;9aS>IRU>C,@b^:f<?F,aRfLZ&/Q.#SKFIO(fYH3K8OCbV6Z(QF+>a5]d
WYd)&0->ZCY_>bY<YJ@)2XNUHC[J7T5\V&H21Wcb[.:-L.ND3C+bH-f:IBVP;<_2
:-W7:TUb]T6Xg^UO5(gU1F5;0GKXLNZ)[H7IdE]_6<JY;QGK20U0\P[IK?,61]X]
0a_JQA7)^.dX-?D9T(YM]_c]0AK4=<-WPJY]A5VEW---#A0R0@.gJMI9V=B)OL)0
&H@YIDERL],I+^A:?5AT:gb/6]M=O_<^YCZ\?_V<A2F1[Y2TF?YGSfF1-&,0W6Oc
bUYV:LT^bI(CJ.cD[PIN3C8F=a5HU,:;ZCfJ6SZ/D(Cf0Ifd,B-L8PM@^?;P0Z[2
,B=CB](1O[dI[d@[1&\UI_Gd;bf2L7C>?BOT3eN/1G3#N5_B^UL#R0Y=d90A&)UU
FSQ[D,Y(N_6,2I0E=YVL-PFN8^;K6;2)=cBV+PEL4?4J)GBLfSW2VSQ.4V-S&#[b
PQ>><QH:BOc^WK\(1>@)7@\edcZ7@A]gf7W^^]?I6G6DEb[&&USe#3ea1>WCcLAM
a^(;FJf#^IMZ,dJ71fXPRF-EbU?cW_(Rg/N)H^UK,,YZ9&T<R.H97]03D-A#:Lg>
6?+IOf@[c(>f\OGG)cYQZOg]Z,Df28U5;JcE^^#:.WR(/JUC?Ya]WdfE9YPL+=FY
J/#@VQ<MUPC^=N;#,]_Mc+@WMLaZ\P4W,BBU>Ig.\I5Q=?A;QG#WbX7L7176]@8S
N&N@PE8J/PbZ)=NL>NP90.P<<4:)VRZ916MGWH0EC=K/0K5<GSIVAGb9](7NcX+J
=VMJY&BT:&3;W33(H5R>SXYI6P<6<R[>ARIMT;5))0(;8CX@]6G)//?.D?MR18:G
7I\B]<+eB.GH[/:e(fbE4JY5f)IWETUL,3Z[7eC9Z#X_8.f-eIU\C.1YNDC)[X6P
I7Aca5ec-S1R36?6_UN4^@U&P1YYV_SN^D8SO_T#<c8EO11KJ8Mc)@;@a0B8LLT-
/WSaE7.]B7XbZ6ULPceWV[)/-AF,LH=JOD/6REB_E^CW-Kf_&c8/\T3gT4<#,Q/g
G=de=Q6<F18C[/?c):;d_VE_43-&UGQ\N&fVdWT(PBFZ]Q<V99?QS)-C^]3E3G;&
6[&c@G&?_A/@<aR0Tc+^,=Y;7N,dC4P8)VV8>MA+_:FV8UDEEZJXP2_6Y)/:g0I)
(8#U0,1KK>8+;_G)7]g5Y2.A\CD6ARWPW;eg:S@fL.CMNbCHRQc3g]4<b(6NEDgK
K]8<aQD?O2c5=@W6WWL#cKUcB&+_KL]@/,AD0<ef@P^>MLTE[WSK28Xb&ZE105_/
L@SaUe]<(7W[d/I?dM0/S.H?MH8[0\cd2+[]^[Y3W@X?3Z=>JX4[9N+&3aSHV45P
d(fYW0)L6DH;[EQEfHRS4.6c;QUeQe&==5=9+\I4)PUGf-.&b[e+[D7ZS_a6KaEZ
X:[0D@WE+)W,R,Ge1.X2A4UU>E<D99=5.;Y_=(Q+],HV\MT(U.QU:d#CJA#D27^\
;NbZ]&#?R#-V=24U;FK+Ie-[E(N[;gY7@4e_#@INg/]CW68_Ff-P71_[W33OR.>K
<JXHB+1QHa;L2YAQY_NLea#Fb/T6AZY7BOP;7(G+0c3BHa0b)35eR=;@1/d#KUgX
)7/B[L8d2=&USM;3d@4HC\9F?K07R:UX@1360<FUfSV1FD)U?^ZA&b-H^/6QECJ^
L);B7b(\2,8L-f9CMb]/;7<+Ma@b[CH9aZXOb=HJV1bUIP>,aX\Q9;7<-ZcfL0\/
T,>J[;aX^N/Nd[c^YGR)VT:HW6f&<_)5J];E8/I1BP3MA.Z-G\<TI6T1U=dTJQZa
I#dH[/[[bHNL\TTZ=QK#LK?N[\5H&NTWN1,])Xd]]5\FH;-a4H5LR4T-bS+S.+aA
0._:TM,#H2VeZ;0>.;I:QJC/>JT0JP)_)aVQe?_cIX[NZ-_Yc1cP^@5ENN@SH(gS
&OWK3G5cP7P9TXK(].@\N.BO).;@G=9S@3,+V=OF:(SLaRUeZ_TXeZg<HL(ULgBY
d0[]GI:AGNf^R7BeK4&b)\TLFCP@=e5HN/3>=BB+ccDbZVX37K//5e0>]X&+83FF
)A:-GK5WM+F,fcb-5-LECaQ&)d;edD8:SPcO5I-fHd;c0.REPJ0T)1PU02&WN^Ag
YB94P?eAZ-4d1ECF?TGg[7F2C=ge-P+L;e3&f?;M85#_/1H3),f>b0a7(,:U(6RV
V.bC_eg9a&=\[Vg.5b[A^>fCPEMQc^G6J0_a;E/J?+1eH3.,^(=NW.:9XWfQ^:Q7
d;D]a@J-S.D4B.SJT5F,/:b(cSN^QTMdZBQ@@)MCaN)59)CG+JfPJY3C?N@.<)QE
II]DFM,c.KLM3Md_U\H2JBUAg5.1ML::LP@ePdS.B]P[R4/X;@T];AcX)(>De_8L
,?7V&;T61\.VNF9dL;SK@DJ,<a/Z9\6>X6c9)CP8UP+P51#T1QgN46_(RS-&+;<3
;NaD_691GVUVd[JU#)b>cXe:CRGETd1&FI]gJ8<aCT6G>;IE\D)+HX,5VY8OZF4L
g_A-#(R-4(bZ9J-OB4g:Q8X/Pd?<PJDWeN<?PGa(@#7cAJQU=-I4LD5IVB=>J8;a
f1<MB:#7U1e=98.6F;_Z]2-<-b)a<;aZE75O<?7^Df;Y]77(c)/5:?7ge6.?&[44
@Tb)ND@,=1QLf/Eb\<dO;O+)?M=Zcb@5M6HU?b>P3HT;f_K?-S50BaLN@8=:\e;V
DQ1+KHB150d2HG_0PK@2HTCU8_C3DZ6ZA)SU[]5DKAVWE^S\]8dW^B[:\W-2.OD(
BTCFNa7W18<,&^ZO8TLR>@^>HNQO5?D_=1Reg.:Q6<Ua.=>2SV>KD-3SgbISS2-O
MHP;e;(TG>8)/8a^ZKK@MQEJf4O49D:719>c:UR>,7M>V@8(:LdSWE9^=39E+g,U
?GZ(E<FT\OAcab4066I\/@Bg/]U6EYZaQKZG<cKV,9dG0X_>H5-UQ+9/495d>)3:
<<\cfSZT7L5-?QUE-.)GdDJ[RLEM)F_BYLQ2S1#d]^IT)RT3gB>=F3V/18MJEZQ4
\::/5MP;RO(c[@Q/=C?a?#gVOI;]GcBV>eNE_02Q#VI04LS4-&Md[^)LTV.HL\0;
<@G7dHZXb>SU>0(Q+K8:&>0gN)HVQC3DQ54@aYAU8-;<YEV^LMXDI&=NbMKR/V6Y
]WP?:90FFf2K2Q.Wc^985b;VYF#;.=VggEM(4EJ_c[;P\-2QYf#^0<&W[MI]15SQ
HVKRG/)8=AL[06g>N1NdAZ=NBVWfI8[D__I)Xe9-PY;5CV^^G:/^CY)1Ra^,GeaS
RCT+EecOG0U:6WB5>1I>S2)YR<L\HZBgg.ZLXR?JA)>4K=VFJE?HWL4M&=+L0YP(
VE1g<<K#781/J,ZdZXd3P]XVeC__G)DaQ7_NR9()RMZD5<)21GQF<]X-=LA0?Y7c
QFSSA(,VH&c3b,\R]=#(LJc,P+^MSKWbKFJc7JY,.:K^2PAKA<g>g8DP6]/ER)Ff
a6@C.#g,QG6Va?9cEP]A\L1:,ZHAZE_N=c_S_bXc8GO2&A<LA&:,(@2aJZT)&<<3
^E,.KA(MT,;5=QbJL)A;e@(K[^g:9Jg-F<#R1D+e_d<2cY?=MJBeU]NIB>g1SN.=
Z7IfP=DL<^9I)=)M@fc_\E]+=GJHN.BC:=.0K?:aVLN_e?NY59.^<+,E?U@CIV_c
-f+e+T,EVR6DId2+,S3=GM>DDJN:?58CZBS6eY-gcTA+<>VOZ\[DOHM&..#/MT])
@^_9_AD?[BYdbL_S5H><<(cdGFGe(4@MOEU;_34)\d?)\DY(ZG?CN52]?A0,S,\0
4fZO@7_5?M\VSaBIc3#N1e66LG<-/fT^X8S3Z>d=R]2PF(TF&7bXSf+g]_9LLGE2
cN\b<]2[9f[U.+YOG\68bNLURS>LEf:?\L<)Lb):>W\=W-Of_0FX4gB/4BJ[D0LZ
.W64CQG7<]^Q:?L[_P32C3UJ0N_]EV>E<d3e+A=Vf86^44#8^()BZ@E,:O7]V#S/
TPV(@-D>fHW_E4aT,1SD1eVfO_]g:_gZ1=69^Z<EBcT4K+3GaX.2/(aKF38;/ZgP
TY@Ca(2Ka_9RdQ\L=2G2BVVVJB+#^GO\1O0gK#N1P;1X8bL:K]bQWPC16Yf3)XQ>
d6)GXDbe5.1b-;(I3ZNG))#L.[<L2IT)_,;S7JA,>@gGQd04F&:OFI9d5L,-07EM
&1Sa=d24MI>GD)L=)A4B\7dI#a(N#424:8095X.\Xg5;3H?R<fHK/\U9bSTa(Z&#
\PR=O8CN_g;&594HD@gcFROM3=APNR-<JY_@(=I3K4BKZ>PZCYHcG3[7eO<.E))^
S(63?1G^1RLQXf^]L<\ge_BUCPf2\S,d&O>RAYJdg0JZegf9DKB;4a;CFJ0FN(/\
L,d.c3GL0>^<_)d6)bM;78dHDGa^:Y9AE\8)3c_:&2>.d;W.BNN+BZH0LedI4AgR
U-6;e?XE2B7U3\^/.#12>WI901:0T6&\+ILH_]?dce<)B>MgZXNM0K^^aH1?,0Ue
234)]R(AW\D<8.e108[=eCc?7ad4F4#]8FON_PA\@R?f<KR+ORK&Z3-C6?VSY4+C
S3J_4EBa\)2cH)b3)&<>IV,c^2QN>I^D[bEYF+X_0K+aTeIVHZa3H];YKW@\;RWC
.a)SYSHFfS^37bf0ZOcb19]G9ZA\Z)ATT5BOef_ScI027BBRI)Rec9Q9=0+6/FbK
cBKfK1M_]ReCOa.;]3-/31aW\Q7+[#JHMQ07cdg?Dafad;;)IL\VI34f_R-V3X5V
?]c+ec4c2RD(2WJ\UC60ID&(8E=]SggU:27gP+\(KMB1c4L@eY0aA?,\aJ:1,d)b
J@eG/[>XV9#C6bC^O:;YAK:/D?:5Y=JLCA+^\S45G##&4=FQHEM^]1V@Q.UG#MS3
HRE+b-QT_58&\aN>RPV+Za=8L=LL4W62aE<1.L04=JQ=N\EY8P>\DWaH>6T2US2M
b?J>G2LG>HX:f<Q:#WX&Q^7E\4U+JQAA.YMBaIJ#^<&bJ:JUE5=WW\27SPP]b7@>
e6I?[59S@,_872#b]W2E.JFaHX<[&;2CA(aOeNOFSQ[aN3E;Nfg^7VHFa^cO_[X9
\G9Z2L;2#RIX&350ZH4KSDQbSLIJBCQf#O)^d4M+0O4F\L=K+VO4.64/TDdf(J:g
#+5e#&[81,CR0C40fX)=F:OB//L@VGX[G?^dW(#bP^H)]VU;28gC3L.f\ZG&R(3D
:J4>3V?()31IO\)U,)G_&:?N_P:,70KIWC2Wc[5W;7+#GbJ0DG(7&GA]P5c0-Z-U
a)S_0f/]2R3Q,@f8X-GW6I-:EBN2EOB-9?^5@[Wa<S+<J\UOMAW6cO9DgBUZ1_/9
9<-W=_;YdWIe-4HJK9P+-gRK),2b)eAJ>Z?HI&T80/_E0R#.G)Ed,N5DG[_#bT_Z
A<OcBXa4FX?-I.AfC.0dRI<A.6F^;,X#PP28D_dALA#;;+#\K:7Y[9@J0X)X]E77
8a\dQM;gWE8<YB[Y0CY<a67ME_1LYVfTaC7YRgYf/8<fW2]>;[>Pg4M?7)L#&,;U
-?9\3N(#5HK\M+<62FWPNefe->FA6e,[XcZfN<:]TZXZ)_=/8DYZe]e[Z[f<M0;8
)8),7,F(H^4BK\:E2)[/RgfP,bL8gE-/O?\[Te#D@bZL&/191\_V=XMa<+Hd9O6T
5<5Y;#9.Ue6]g^=7/R0959c_Af3KR_)9>)4;G,2#K^+U9TCX+[U(cW/dGJVKVT==
BK?X39;=O:ATf5<\JN;TUGETW0;L_K_EYN<K0]Z1++_>D&1fI&/:b@aFSI8cA30@
S+I9IQ#IQFdC[gCVN#0b-)6]G,MOb944LL_-cSB5Z<7O/Hd[Je2OHBM@bHHZ.0Ha
X=Za0.S-+O>MS,SeJe>453OR2FI77G.IVV0(:D9I8,L()759eM[MESb01C2Ca+4<
\=QKa57bDWbD.2SEK_>2,;3=]K_&SgD\2JNZ4S9BFeGS@SJ/DY20JT@3?5V\K?-6
]-@b<dbB(+E-#X8+4OD18Z68-,=N=XfA=a(g-K<b^0RfHML_G:gUSCS09PVL)/(7
fc:(K2,J_E,?>.QZW=3,_B@AG++aReH9XaG>.Id5dA[U4d(2J#SC]H3M)M11X6T4
5>V,#>9I0I.X_G:I<dd75]3dZ6X&dZA_/L&E_a_LH-eIU6C](Z)0cgNd3109+_5,
+9cXa=)X:<FCKKECNT:aR8.Z9VODQ:WbT2C<5[LT[5&:]5[T347[SS,Pf2QQ:I.[
d(\<@B#:>ZR?=FJ,cPF?fW<G:N:&7&])=[4W=8N:AV0^D4E0+TgM#@&2W76)EO>C
R_6>5S6V5_NEB24a#DJLPM4d[@-TFb2/O)2eIM=BXH:NQ#7BS_JOO.GDg&+Kfd@W
.IHZ(c>I<O\[0A_@5aY<55Sba/gWKWD]&N8HfPaadS#:g\Pg&g@GX>CGR>7=Ka[2
NJ03egPEOK-f7gIP<C^&C9>1:=SS&G\T//BGFJ[Y2Ie^b)PAXU9;/RT@0dJPEXS9
VAH:/O0K-V;T)9)3Sdg[d7d@If:&a+4#V8cO/9F5d-@:3c94IUAKFHR#g0K,L[GJ
5bQ-77cC[eKbNG.)KaKTU.IS=9fH^V[)UJR)0\;c.#2;>?KG6D.JL7(f8TZ:C:Ee
:^Y_<IY6T2(C[DG4aDPAAa+N3@KW;YGUZc(D_gE.M(f518a\WS<-ae0D-FU/eQ\-
e5>IUYNG7:deIFCT\0K7Q/B[V3<79;;#&RI32&<9f:Eg9^9?\.9<@G:_A5cY=#bR
b0K)5:,/O9V#gP:.&U[85/V.c@;(.L9):6:AQ=;;g^0e<dB)A#Z4=0+TNdGLaB)\
]aF^QSL.7#&CS##C,C^3,0=E/TBE3XdbVMJ88Re)K<./]\fD[BKf>[RW8Q.UX8\(
J9]R#+=&<>&gHC#9f<#BdRY2W/N38E600GG7Y5ea=1+aZ-)cVRQ&>Se#57CJc[5d
:eNKe@T;R^J=_-^b#5gKJ_EHTSH?OZAA#7Y2c2+N]ZRg3FE:K0QRfFS&V,Z#8_Ze
2<.A5(KgIc0NW\69CE8/SWCI9LD4=KI.\MDH&bZUUNCM24HKgMfE7=YcbHNJa2W7
;F/Gg[#GaXPRFMgQJ67N]^^:L/R6]:eW-/FRU;GY00c0N/?J?SR]e&J;,)c#+N&U
1=.7Qd:a\VfGHM+W0WWeQb\-YE28[K).&[9/-F)0QG=U/eVN]N@)=BFN;3>X)(_2
91,8CS58?.d;ce-Yd0G1a)G&N=ee_bV(^X3-YHYVgKe46/)Gb6S/CeC7^N^;=T21
4J^H&XDOU)AYS+UM5W&3cGg]5@7[F<2U1QGd_^<)/W6E^N;KE6SKF>#0-E=#PD]]
SD8]6\X@^=(:Z10P-ab4a<-R12-LLM;X2)/3PORQL+W<bH4OI43ec\.6^?E0dLc#
,FUg/L:MK?&a\W[?9aWRFB6LdO.JTQ=RN/)4?ZIYOV;^]5Bc4C?I9RUO+9G;>e4^
E+S:O&R0FVQ3X19X\,CF/[V/1D/EEe<Hf\\(#DP:ECEMP>.8E3gRY<H&8ZUgHda.
;c68QVT,>(]RBMD8YMV08VZ=J=6eG<]_V[?H\C2AQB:20Y2fdA.ReCXR/87]+:_,
P6G4:D[MXH0c4LId=IT8,68=Xg[C,,T?,[fO-HKD?FE5M;?9N1E<I=5ETcE?XLVI
KV&RVB\K..TC:C\]Mg=TDV(YV61UPU9:4BP^75Q,W6c:U.CVU,5RNPZ6A\dU_N4A
CDSND2)DK/DV477UG_a1?DW)K\d@2Jg+1S_C?NeMF+GTM5.CK)>>0CdDb=OJ33]X
,RU-.)gK2F:BdbE,\:5)K3JY\6\g_M,I&5W/1,g^L@EOI4;f]=WWYD#E,Z4MF<+R
,3IW:=6>PO(5cF#S9KGTND5Q&b2=L6I([LG/9fMEPMS^aV@,J?^A.8TgdMW#A>D_
OgLR]MHDHR=[?g<VgaET\+).JGKZ4^CF_\/9dWV6-\NGJH1U<[(8TI);0cd&&_-B
O/ZQ51FbDg]]e:2fAaVaT)7c(N[0aTP@JaS_B+RY]\QP^b59?>Ocb1_/Qd[8RQgJ
0.C)F<bBce(d41A2JL+:PQb,W<AF_,R4A8W)PDH0-?T<=;&ZdQd7Z&<7db@-?<3[
IS^[XGd+6[^3W?^;aD;Q@C3c57,4fMY_d5V:fIDAbFE&QBL?)EMVZ)c;_L?-<QM7
&D5c\d\XXI[bR@/YY^I?<O_@f&.QH7Y?:RdM)<6OY1#ZX,FXT@7(&U?e;gZF?7V=
0Z4#d8f@\c)N81=LVQS/8=.CV>0+.g6dL3QW6]1VBZcT88(Ne8=JKG,=Xg>)(UE8
5N>55,Sg>_PPCPXP[CX6DXGBD89.Q\Dc.8;D6b8DOW#DWF\_^G>)Af[Q/>>2fL8G
6MGZ##EL18\EU)HM]SV3^>+B;2bE33f,B.g#]IS(6a.)a#;LHTYB\Rg^D\DYMR9J
P49&J>?J/Jd+7Q#J[(RP/Q.P@[=B)8VB)9]c,WO/L^]c14@\e]FdIVf,3_W@5aU.
77ae0E]/U07-)U-M0g<f_#N>f?4eW,8Z-W5AANN>eJRU_^\G[;Ba=H5\X(JIReHM
_Ze]a73NZ<)_b^aAY=;=#fZ-#K#-,1:eA>^:\>11W#D\NWQcP)SS;5M\A<b71GR5
3^@&6MX><VYC8g0OX&G@Se2VJ2Q+P3c4>H2gC+[5V;(/[TgTZI[L=)]33F@)Y=gV
[@(bSa::&S#0d(HCCR-<c^]d^b-?LFQD7F?50]O?(Q=d6,NORa1,Z,f0DAGCDR6#
]S,=4SVSfdV#T(EQRO7_5QQ9JY8]?4MN(GcM[BfI1fgf1c<6J\218ZZ=1@gNd\6=
G(5ZTW;ALANK@+g^JY27b8N]XJ=>(NB3C0PM=S8>T964d#@HgeAda1..cH,_PAK.
=_6&;&F,WL4<6Z<-:1e6<^M\a)S3<g6:<f\3-R7:BT>f97-(0V/e^#3YFJZV6&6a
)U6.D4GZ/O2,gEN;PdC(G2NZS2RH6f:;;VES5_YQZ(efWX7E4:(N),A(&2TTJ\d?
>OR+dfOdg8N:E@FG::RAKRUMV^[;D0GE1C]7dEFK<SLZ8>=3-:1_R)54O]@/:G:R
N+9+BFPg+R)3<)2QD7\(XH.OJP38#\Y0IDVTDDDHYFJZd4X>(g(aTH2\(DR?1G.?
e//aOA2,=4/6OTK.Fga-c+=;WcBWf_15[)LAGGFUd&1>Z)NK^?F3a;_eY]DF9[-A
,2[?[]QE;BVO&?DYT?5fZ7JJ;bZ/.GL9RQWV4(KP7<5)#@,-f,ecKH#=O-\U(RXH
T?&Sb#6NbRa^O7Yaf=PeR&7-fKEQ;^;4Q(MVe<T@W?(8e^(&4bJL#P.0GM_LPTc,
AV-8@KF^([fK(5>=a@98_B+VL><Vg3e<X:M=4D.+0^aPYF()#CSL6M&#S?#U8Q>:
W68J:T6#F5,U-dZgF)W^BZU_F#^e<V3G]FC,=]\<gG#8T>T-18>FI:=FNS27AP8Z
PE(_-8_W;c@:43;5C?UX5@<4U+a)Y65AK)UKI-8DLf,6aQ#4QZ5(a4]Acb+/<^db
5+/9A[UY:Q.#W7a(7@MCQ0g],V,MR,a?7WeV;aDJ)YV&#KVBN=<GNFN_BE=6b/??
RBE&L.3>HdIF3S4Db-X.TBAe]P?fT:3JE[^&D>b_=&EAfb0g/W,L@9gA(,,^b95]
?dU8U_LI3F,R+EE74SGI<2)AK10fd;>:4MZ+7+fcMRHdI^/Y=Mge]/b2d\V1K=Ka
@KC7L1JQX&MIIVJ6A1Ac2^GD/g&RL=0bZHI4Z=Mf[^41S[.AG];TeYMZbeTOLC^R
H3f1W[E2#.T_Z+NZ<a72BK<KV^#@Y2,,&R[gbe[\\4SLJOF3Y@NMWYcV^e6WXfC>
0H>7DH<4T]A]OUJ9a6<1(BXWE+,HD/)5,&C(&_G;07cJFMcO[a=2Rf]d5e=3FYgU
4aX1@g#P5YHV)#;N&T6DYNHa=MHXZb5ENb<g_f>U9PEA&=2E0b6G4A[,fG4aWJD=
Ve;758[XL6MR9Ma:bMC2Z<#YSaQ0WE<7ZN+P4P-7gMC][V>/:Z@X0^L6=K@bbX@)
>^C-VQAPVMZe4UZdLF2GXe>OO]:Xd(N[OgQ,fVAYA\bbXP?.>,&X:aH@c0^=O+0A
;@<SF>-9XeTcE.(7cc-L+(SVKL(L.1=-UJ6MdN9J,0YY(-V5&Bf?_5FY?bB)HCQI
493c:33W.8eJg\O6:Q/^>:cG7<g0Q(+@9/edAe,e=B@G4ANI?+6-=1O,\,4Q?L<M
/8>^ITXg#eNA\[ES<,DT^,OC9@7&-_)[JdQNN:?ALR-CAd@4L?X<9RH_ScAT_bLG
/,<#Ye-NTRA]P3UW:=gaDLL=KUDGV0>HOF[:.^6^_-g\^3S(H_:6DcOY?bG4)72A
A<EW(=/=V[a,,1\J4MC@RJ;eS=8OFc<[=1(_)I_:+OOI6eNF\L;GYE2(;Nf_UFGD
S[T78\C_SVbD#K(QW/6]GEf89[W:E-XcG1(CZ0Cb;aaAG\:g+dJR=2-)gG>1&M>V
.d(Hg;)d4[T_<XSTb,-bYF<E,9Ya=QWeJHfcO^\Y\:)MI.HOfR:M&GH,3g;#L\K+
Z/CPOJP4S)S]@VSeS1G;^5A^Kd=-?(6,CegYc>.HP42=Ic38bQQGSD5<G)K<NReH
2SVE4/PP<a26=,QMA-(L,eB?[Ca;3:UBIbaCAd)4VFNJ&FH)LRJ)EUfd]F5.7dE,
^VecV.;E]^6#McAaKXbNX?9CC,0[Y@Xa1:0+7PHKFX_N#5_8/F-+ePJK.&PK&(;7
HH]GaK<CYB,OZRK<EU7eW0IQS&V.33T/D(\^F,#K;:#c-f)5gTPfXeD03[M188:.
9S0=Gg#V:I.1TJgP\01U0GUDU\MZ9^&CfO;181Td?0cPKg^X6ZH;3AW)FI\Y[ASK
?,Wc>&GG1IC(eRF[AQ.)7ZBW[>&E9V-S:^-GI)BdJ5#e5-+X7@9=Ag/C(HLU@;a7
#OWV@N8LfR2DQ4R\R-NY?E/gR)8J@(&a7.D26]_^]=\-TgLBE;ZaM?:RD]ZFX&5<
S;;#S&[^5ZT>7YR1Lc;8Q9U]+=(:abEZ0]8TbQ@W:f+.RCB\..)199(FZ-bE>KIH
=C_0YP1?NO/<Z)XQdHC^MZ71_.[Qg118FC-&I?,JP&ESY>8+deO/G1Dff9A@7;b8
S;(7Nd):U?Sg\R3].#=_B\ZP5g6KSOOW2XFCN#HV#JM5=LfXF)RXIa2:XeMaLFR+
EG@K=P([/+)K<[8gfXU?7>T.R.&J1&&Y29=b.?9;e+d5S\e5@AZee,L;agg/F^]H
?b,=S/d=EM@JQTK@0MF6FAY9U:eggG)@E5,=YW\?0UA&#\3F121OE)-WF3JC&SB-
1<:dF8AQfdWSR1fK:?P7TLPdROY/Ua0a#f\&cf@J:9Tc]daZDcY9>?/:WTFL2AG#
-GI@c/_E7U>G-cTgY0@GB5OCb2NW?=#HG\fb_>3H6-SN48MTQ[,c&e46=fB@gUT[
T\8\BDPS3&MH6M;V(60PeA6V,_[4\P&c3+E\4gF(b&@)A3E/T@?Q>C[?Ha.6cJ;f
;C1EEKB-=/2PEFKU3bI>fF1&9(I\bc]HE4NO32>CAADM<8gIce[(G+Bgg.f3JD++
NXE+O4B&4Xa-F>eHNL)MWAQRM:GF_CRDR[1g&Me=2Sf3UGF-VY?Pb)T=EENWCJXa
WR(R[.:RMSN9\I.Z<a\>H0<>415]7T71-(ZXa4\TdL82&&TQN5g)C-cCDMHML5+O
]H@V:<(AX@FgHeROTL49;UgO:g)?YU2GY6Z/M?b\5C4;][e.77T+0PNY-IbU+;4>
=LH2OP_<9GN5HB_&\gc)c_.JUWe5?O-0\PQDQ/>@4@S]27SD#SLDW@Zc/_7fDgB[
WM)/CPJ(.IJQXa(JSf@=-#>=2;9LZX_)8ME,8B(N3e.bK6>TR(#QT+.G:,<=e8:E
bIJ,L?<e:)d=J]?QI&0Z9(X7GU0[.3G1:d[SIA/LA_I.(_@Je=XI,G07@<U-.eBA
JTA//3GB?RX8aPeMP)^-6EC6X2E_e_e.;Ne3-9AE]F18DNUb4>/4HE>RbMW(UWM1
aFCI3fRCTS^6VX^a7a9gO872g4+@IIaTFCO.Q>=Z9DIKId4UYN>9,EJPCNBZ_KL7
DA>a)[U\O=c)8N5,RXZCcTJDCD(@/9[-?DJMU80M^Kc1+-S+QN=RFD:-JM(AGMN/
GCHQ:STPM\7APY#NT5NbN@YNa#GB(D&UM/8cG2V<PE?;?F?Q8GAf@/,3ID@ZY<J^
DM>YOgSKPdOLDd>c)<YWg:bU7.PWOI&7J#]KTAAK?#074/Sf&K9<KgV(E_>N3gS?
;+_W]&EQVJN:BKG8ZMBB^KD_IX7L1_D<]WPeK@7agHGO9),]+VQ8d^.DONEHFYN?
+RLAcDQN<b9>?^SOC-AaBR(R0C@Z21@U:FV;b<:0\Vg&=]gPW:;?=,H[L#S]?G/4
R3QE3&&L5<A_BPV5A.\Y?N0-C=,2[dQVQ[46eV#PMf2bZ98D:YE&:]-18eDKB@Rd
,&PAe-P3]XEeK+HOQH6E^,@6\R<1/L16F<K?6a-@/5:J#G<E62+C/B[U@EfP+^8X
Q.LK<)E77EN)<V-KIQT+K@5SZU]H,+9H3)IUce(aZ:S;>I.H]H60X+#EX6OIT9-M
UaeaP&gL7WU^.KHfXFJA&P?[=V#H/_)SI&E=+cB(K5KDHB:G?XKS3eYCNQ9-.g:X
1:.WeUF^dDM6GD1fZV1dSHEPVC^-(bCa>@Z3WgN@]H[(&U>Y7GY7&E,WTe<XY3]J
@\AS-RagJ/3FJd.>0BS0edTJV-NDOZ8)6AaA>/N3(G>JR(VY?,GZ?M9@Kcf?X6NH
:M-a5\<+_2M)WZ(NQaeZ5-PLORaATG/;M#Y@)3aURE(,Z#;GR3IR9f:U7Y\c@]L[
\eZ?dbEg)URDMba523SHIL1P,Ga<#366_g82b-H7PHaIQ4;IF;P:)=P99K>A#-.3
CQd+,,LE)(e;D]HW+7dY]<7fRa/6LS<(SWb\@C(JO>)_FN<f9PZ_QK^3Ma7Y:Fc8
9-9L,VbLPO_:84=^[EA(Z)8PZ+X90+Nd#V0,)(,P?]WcAPRWP9Kf_SSX:E/4)g@D
2PFa0X1ECGd:#]2KZIVB-R#)PX8FIbVBB1[-5\2fQ2YFfF^>VQ=G0.f,3DW443LL
dXXA,#2+J.\\c[CY+VA0YRE[FD-.]2f;<b;HW:I#b?XQ:Xg--e0G]0\0VdZWS/Ua
eM.7J=gQ[;Zf-/81e2F.5&_e@5U]+NWOM_7:=+(L]>@/7abC&gO5NVYGGG#6[Q,H
1(WHMQQR8\.^.FK\JA/^9=)9B1FcTV>#YcR)BY@Pa^R\P.>J/LZKHY/99Z:dV,63
X1^=bCbOQQ_EG5E6+C/P/T.a7(BJZTG&A3,:<De:\e9F3RPOZ@3+Y,M5L[/Q81[V
N>OYgb9Ya6PLUZXXD?9e@aWZd\S)Sae/e&M>]P>=#N@.[JVUPRLQTQC2^GX3S+,K
Y\@E(^:;T/_Y<K@-L.GKFR&ed[#Ge^He-=0W#FBbUS,^WC/SXg5TBcaR5dVDF:U1
+(6AS8f@QCT2>5J(SV1_^0,A&H)3)V=F&J:#27HS[G9,F^0JI[7Xe#cRB<N4)J6T
.4ML?</AEMP;G85M(6-1W[SH53<f8\O<&SA7GG=_ffON0cK?51?WBYI6/48;GeRe
P&WA#W\4H;#d7b<TN]XdMSdH1DV<[0g)5R[MFCC:4&)?ENF;P-+AR_@-D+X(D?f^
T9Q]3?G/#TC2)&+[-6XIQ5A(Gg&I9ME#8C-HI[9YM:2(#ca0J:FR4SZH)GbEbeVS
Ogg=M.T4>>ED<2c.?^1\g3\>T3/FQGd[;_VES(C_NJGc2F&L8aN#-RgNUR7))(>;
H-b,6.YIe>ID]X5]=TCJR(f0;Pf5^N:O^cI-_FeKc+,X7MfAD<@&0Z;X(::e.P;R
daYK#5\NHOAa3D3^G^M45)HFEODce@BbIBP&JaOfMd@S0RBU86BS0BGY&V+L^TKW
gZMO[GA1)c;#VN&e][(2Ke68G-ZUMBRJ0ZEfGRbcG64A[4IV=6:.eC3eU3aL8<)5
GA+(3Mg<T7IR^UEg&OYYVI6QA8PaE^J3d6\:G<>(YJGO@QQWa;N;Q?FC1</-KZ2<
>b\YMESH<#FI.04XdO2g;d^dS3ME9HZ4W@[5K9gVIE<)96<@Z^=,(@EVb58?OMU7
>8Ue@f^DR6G\gMX&]<?\C?ZfM9fW_66IX3UMc)C(7WE&XWA(O:Tg@Q=9NLWHM\4\
#5dLPOI8_T>7AIY\5a#M[^12bV&a/@>c0_YKIE+(JdTW+/(=&Z.Y;,?N(/1fHX.:
MQA2955KFdMZJQegV2FQdd5DN+_EafPZ7ZcK626dXO-:EK4;9&8C.aN/W,V+0PP0
c0?Z,O]dH6X57f>f6B#dB<Pa:^C&7cB3&2-1N-NBKWgM1.V,>S#,ORQ,ZM@d/(/-
YGTJV^BXg:PK-9fe.Gf+9AJTDRQVJC6&5<M7WHK+<2\A\99=CGL16GDfdT^+cG7I
I@>GEcZ_I)N#^D[A)<Z:[(fB<EXf3T=W5CfQdb&8IW4SbAO9VM7LJc^7:UU9CFX_
2788W_gJ=5;_Q>C9c>WNZQK,[#J)SZ9;\A-7P\d73\&VA56[K8(OY,6XS8C_L[KS
baafgeTXSF)</6[O^9V?QS)R.+OQf]CJ(,L,OMPK\Y@[:P^\&E4YQ,QA-.T(A,0_
U]:#aPF8RbK1=3L)E,eL)XcObE\R&<PKU/[7FgHYb,aJS_+ca^-(ZP/3>g6a)#74
6G@E/095=RT=3;UgX50a2YK>EMN2CF_.e\<gO,E,J5GFNP=#&2ZP8?4afO68I5fT
F\3S)80M(Q,fGSgfS&9_,^b/Da@GL<Y-19)=S^Y<6,f>1E6SHaDQ)8UHN,J<)2]L
CdW-O0a]geR;SF,2V27aAJ<?f2EXVBO([eaH9ZKLX7EL@R>N(LeM/5(?JEeQH=M4
\eL)G)fC+@/a&/e8Wc4(Uf58RP(@gV#>YJ)2aacBg28:(04D>.F>8+@54L9R[GS[
7VX,KU.?^[CHN,_8Da2EL/)FJ./P?))0)D8E.J4HE]0TUKV)9(156L)\[PC9ZF[;
O-G3f+WBY-DW-D,1fBS:TON&4ZC6bN_?8RQ^Ceeg2OLJ\WAag&)#P-Y?#Yc-ZE7F
Bg]8[cZ+EXU>@C9.X[&W-+9(YHeM2&fHY6\a?XJN7&C[]:[XGBFI9-YXbB<f()EQ
ND4)5O(<A8JZ-aL::-+YbILb()ZDIM8LUF:1e_e;]McQN?7>#+QTIdHO5(_SY^N3
ZM>N_D6I::/A^_]UT2__Y@/d:E:baSVSZaTHI.Q2([P_FfXg^g&fW:,&XW-^_]5M
c#Yf2>A[ZVaB^50b45CH&Yd[+_LQ7bIP<?Fd]+_ICgWZRO6;;1)/eL(YA0N(-J3\
L7Y<J]b-TVJYHB:gK4T8c9??&F;DB:5Z^<Q@X[;,b]+Y12#C8VZNGT4P0[N;U6LV
b;_)12I_d.WW@/D?/E3C:F:6F;gM>TJHb1KD&@NL-KRJOT&6()KIH8+cCfd4[Q44
LegcNZ6&W3G[&Z]D-b0F&T:BRS69=L^9NX:?FI#ZW@\PAQJRAZ0C[&ET3^#.4f(N
:KRT.&ePeOe55dQ:W4a=YDC,-;&HU[YS:MXQ@Cg1&G4Kg/)@GP-1YIY8_OdLR)fA
TOeg-YNf.8B5#=QLD_dP]0X657CQT^G-9;K3gb_XYS@B@5_eY2(M:4=eTE=@GQ^e
#+M@V5OGAZ]JeWN]O1(^Cf.Z(?@CZ70D^Y+5;+@aFP84#2c=PF6QDeIH;:KA;[R-
9C4FW?aS<87F6MINV=_7LW(QGb:]a_M2g.bZ5Q)])+b:,)1Nf532^/I#V56S9E9;
4P,-K3>LQ1XO4S5X6B<62Nb@FZRDH>CBJa^aE]GF475f>GJJL,bRS+9,QD\5(e5E
4;Qe-HZYS^A1cG><BJ;7KI+:A0^Fg6WH3^K4Ua=DN,7^_?H&]LE,7(C<=29Y&5C-
3VN[(P+#G0^Z/H7Ce>BU5QQB(TGZ0IN28F5>/Qf.-Q4+#5715NE18JgN?V=R=ZH,
SMWYH]=eGKab\[]MXEdG/O>BgZf099e6I=6<84,1.PgQRO-?f7c/0WJ=O+F<H_5S
VeF[bLeW?_cP^fdU0^?]M_\093&EUT5M[Fc\[V.MbG5?R=?>0:&YOK[-3:Ta?Q;B
)ca0JbJCG#-#HT;5=W/^@CP&NT5XEfKa8E-7W6-ETTA2];D00a&=&36BUF(F/eV8
(OAY1:D=:G1BN..7T9aQBXI<gaI8a9>Z#G7]2<_2:8I]U6<CbVBT^@faVDWW;bKC
P7JN9&=@a9DeNdNEP2C,#HB?G;PVg(XQ2V_^M\BG37\I4dP^/_OP/@VML&SP\JO-
4LVY+0A9N8Z@TO=Y^+Bf_;-0R=8ffF6X/N.]6bJOGHC],G=>(BFDA.DHA2F&L2GD
HRM+G_,G745Bc9B5.Wfc3C-=L;0_9_A</X-GS3FX@V9PgZTC50CK8aVd9K_-,WV]
W@=@F(CD,eLH7.OLIWW\QccP8Ea;gM6Q8g,X>E9b^04T,=[,MUH<-T=3T_[,IJFK
5^P&WYX+=T)(E,1@aH?&;1]4J+/YSYA65Q0X+SHK+c=;&#0;Mcf2,7+-?Qae2SK+
3,&W>/.F98-&gL-eP?-N<#gLII2DM,>J4F(9/E7dYT6YM2B.:81^:B^0#3,+[NSA
GX/9F.eYJQZ?M9I=eP&&WOUG]JPIDb4]a(4W^TLNd,.CYH-5@/^@ON1XCB,D;H)S
?8A7E0B/\G\+OZaA859AJFT+JdIe)Y:I?+=^aI:4ZgGdL9c3B8f:bM7TAL]7&1b+
-L&K_FfC&afbN_H]Fg^#G7CM=GgH?MUPDJIM7.<T&H8NOS0;?IO7dHD(#H(TH3LV
0ZN6I\WD3R-OFc39CZ5T^):EQ>ad-Q@OYDN5e/,\KdK&@9D:CMW=(bU@&MP6,3KY
c\F>/&<M5REbN^&#ICgXf^cK[(-&<U4Z@_=JC)/XdbW.\ea&)JQ,T&<>1-K9c]F>
aXL]1<FH,KL^4R#LI>cG?+a#Z>UdL?X^]:7;KCD:8PdU:;W;7V6WI,XMfVd;1Xf>
:V5@]\#)a?\d&d8>]6VBTBP/6.^Q:+FNM979[=#f3>U5gYH08([N69:2P:fX3Ub6
Kb657F0\DG/6eN\KL:966>g:-]=GD9??b73A[2+-FBIPeZ3.#cFcY._BY<MP-D.R
S)Cg-.8_+M3M&V+L+XB2QGAJ(=\7WB.QQK\4/A^DTKWW-C#);G#8+eH+aT?HdP;T
-;#W18K?SML<7_00#U&^a2aO.,cJdMELTI-+M[GQ-NS-F60Q#<9-=TF-U)HBA1bF
eP^C=ZVe&G2O5Z[e&[BIP]:0K92UfaX6CGLCFF4=RUF@1dICX+7?HeODNFVF[,L?
:+ZHFQK=06LXa_NBI1_8;]=9ba,-]Pf]I\VLOP;AWWg-Wf]TKc7T;ZD]5d#?e)Ie
N,5>O&ddc24dQ(XA:L.c,NaA>H/d?LU/48Q,7d]=R+a?aKAbO3NO9T+.5L@WQYEP
H]/DbHY=e&D34?:eG)=2fT\N^XE\CEC>ET/FCeQT[6Q3YI[WSec,U&gN7B+^:>9R
8NF=T?=?919Y)UG2154>UFAYSK3B)^3CS1--.FIC42<D9Z>IOS;FX,F3M/SK\14S
eS;76Q)S<5AE0)<U=(=?W0aZg<0DdNK)1LQ@>Q4-8QFd[>5TF2#4NDPNc(63:a@P
-D8O<H9-=[.&S@2TaE5HH@NKWFBNQMCGg^W@FU4H@R+4PNDZ,&/;dN=79^F=ZWAA
Y0P/IUY@_KSS+]gL.5dWR/JTDXD0G)A1Gfc?>TCN]W#SSbG#H-Y.1E>:EH(a+A=B
IM,;JdOY.U[Qb9>O]LH=<F=gCMYS0UYX?J5<#/g7PFPa6OT-R;CHA5(8FT+G/4Q7
NR2QA,L1)5<XA@YX_b,Z)gEK9(+R+-(46+7SFSB0R=D8]].(JD9+,)W_dW+=G=P6
4YJ)5@DWKYAO9;gNUe38:MNH6P98PC9UP>1>G6e?:(4CW67T2Q8X<Y7N3NX4;6C5
X.D=dAI#bfP0SZ8;JHD&<H\Z8(1B126LZ+5=f?6e=I;J/ONX\C+0<52ZDfM<E=7Z
;0H(GaS/aLdO(Z+bTO-,,d0c/MYaTb42IYD(H#5SZIR]I9Yda590b^<<0[^VTcaE
DA)?ZfaA79FbN(a;^CDg=1?@<gf@;8G0KQQZg&L<JgMOMVK]+>IF81[@CK8.c2Eg
.<8592/^.?_De33#Bab/(3GH)T=,cBYacFMbW@1[SJfC4[+]b,=MC\EddJ9,[Gg]
^.<;daP1[?<-dYC&(3@=LJ<aERYA?JC62WPO:1VH#],bKM6M9NC/1WM->E>D+&:X
-CUO&&]]bfHH7KLVK#O=-4_I>(N/4E+:eTX&@6Ae,[I4+6g4,V&Q05A;&&AWBgR7
/]8H8U:IILZI3FE6V-R;FQ.3Pd5CAb1XFbNIdUGSS,42OI@fW#Hc-G@J@O+U.a>T
58IJgEN+Y#V5gc)]H\^>fEdUdU9\/CJPOD(02=CCRHd.ANP(=)(GD-)_Ge)K(^Re
\cIMSJ:P5<0EZL-d&,-;3<IXNg[003,98^DM<#CK;G6/:RP#A4Va4,FTaeKNBXB5
_g?bY9K-N02ETK_(7[^(U=P23>Kb61?:5A<]U.@;C7d//V&7C4D1#bSG(Cd:G>:c
1@FO0=f0]>f:BPS2TAeJ-fMMcUHJV?1e9AZ4gDf(Ta;b:W^e3B]8MeNW3_&J_D(O
NSH_c2[g[b24&5.DI-5M#78/?:5ZcSG(ERDcO6XGCZ\.b<a0-a/HIE[a.SCe[AZ=
OI9g-YaH@.F6[[WX0Fc[@UC9=(X:\>F^U?UPaXdcZ<3cMVHQB@dTL^IO5#;d?ZXA
2d](YI7aHe.<5)G^@@JT?RGKWEFgfd>_NLM8Z=b&FfI9=;AUFGWL5]d?(+DPRdY5
.+A=V0?K0J?ZF]8O>98-,\-&NG5fgBR0E\_M?B8E]VfIeH?_Dc),-#^WQKHX)RW>
KfgWW^KaNR5MdAF^ML_8&QPeMc.eRK99B(G+]aJW@:\g++Y0H3N7N#eXN3d5?5X7
1b=5Y-d&7fUG&_FFNK:TKXHHG8TA=;P/^8KVW4<W[?_0XUgY\MY++8SIA#GcUeb5
BK)\E:-aCW(=DH:]7aOKF,T]#W0HY&+U@bYWW^1dc._X<Q0H\;37SeSHDMJ(/0:,
L,@N@NC(_@^6gO\KC(G+Hc9Ne>.]Z-K2D>2VA(QDU7S6M<1P=IB:OLQ2d&]&d@F,
>XN._cX0cQX(bVE]+\Z+aUN1+3Y43M-@Z#5+-Y&V,H35YFC<4R+dFQHT9;cO,<dU
9Hf1&K^C26b)L;:8(_Bc)FIHKK3+]&&(F[;Y>]2V5XFd8@AC^NY;9@NO>;1dYUD/
J;[=GO/-a[c1SD<BaG6HOTY9OX#3#@3=3^A@^DFY(N-)K=a.)8ObLHY?208BHea7
PGL_?UX0e^cEa2;Q3F]bI9RH9d3VM#_GYN?@G^E;M9\MW,>ZN2,_#;U)5ba[;.9J
-/844&38D2?BPJ3C.X<9BO.?D]/-D;(D[^M+JR3bT8?&?cIBeH6?\P;/A)>Ig]BS
VYZa_QY>6-3CR/>3LF944@dPF14[(eIfE:#XLGW3M@dEX#Y<O_<OGYaA&d-cVO8&
G&NdH(_HZGOTLC([bUQ1?TdEB#-_C_V=>SJI=YOBOLCG:?Z/#RW/B&?]9bbC/4OZ
FGcaTZZXW3S97XD]c2g].L(e&8D8#B:A52/S+)]3W-7&);+LfCC8#1@Le\5L3)1b
;;L>SLTO,H#14-8JIXeAGZ7J[EQ=T3SOR\Z,:WL,\1,-Te>/g;BE+.\[V+IX<CdE
07.?HM=X==M=.P;/11Uga)MB(1[COe0D/^N6WDV<=B@:GYABWHI(^T?+XOd78PW;
B:EIeW@\^?P.cJ&WO9;K(be[H@46ed&@Z4B,\?)9_&.F>]EL1:XTADCNPE+]1UYa
DaV<b0/;QUfPV6]USJ8)0\1DKYa4\<EI:B[BFR#aL?)CZ9Z?>B:4eGRa^C4UEY=A
:6#;,)4=0[Sf\=[c8FQI6<77F.=^1@0a&dD2F-K8H9GK6_4BD0;Z9PH:GE8@2WKK
-eaRMD]6Hf1@M2f65ZccgK3;MGH+/#AY0]7X-(FF/PL#EE?H]?IU_bcD67f4<2e(
EI5965eA@BE7bFE+V;W[G4BSFLKJaICf@db>0Ldc=a_R#9d2eTV(^-Xd)=H4LaUf
151;9dAB(,KdL(c,B7Z?T()ZEd;\-Ya>@_-&Z>f3a)L_9a6HdH3GL#DSW@PF]YD=
W(B@aP.@W1ZZ?RU69BDOdDMfA:ADeGZB)e<Y[e=U6=IN;P3PPQ7B:C=aUc^4^3,R
SX@_ZIN^[EF166C-9G6a_ENdSE3YOaR(CT\)#F2<Q.WQB1](N3EYY?;=)(GOBg#b
gVb7aB[F585.N283gSa>SX4889V;U>#g8/+gD(V,(HWIFa,[aNf]@QD/W>=2e_RQ
&JK>6RT&6_&M5AFg+Gad;M#.>&C/5CRV(W-3LGJ8eAb1.YW6#N14<I_<3J,ED@e3
&=e.H0[&V=c)4M;8_5LNOeZ(L6,:b-X3BG:KHg:4+>V,f4MgQNTE>J&@8g20Z[ML
MYGd>]@IH>X_B#a0d-5L:;/-_2TAdeaH^dId<\\?57TJI_(</,9FQ./ZSS^;R#QF
.I3<)&b7aZXP5G<N)74&2?\@\?M=QfMfC.(IZQC\V(AMFD.W\ebM\e8[PFOPc,0-
gNJ=7:?aLCD\Z++G#L/P;eQ3E]HeFf\ebPH\>A-YCgKe;G5BH0,6(GgLG)Og0)]d
9<0894=E:FX6Ya]aF0OIG?+.S@YTbRTc#PL,8:H7G=7gD9_9TV(O=[e<066g0E0F
gcF^XDe1_;Re0gS9\E5A<73R3^2@:cC\OUEKcV2Je3EELXMM/73\>]d=&FON>GJ;
MRIJAQE]?,@RY7#SLK88^[[cSO6_@&(-Ldb9PQ#B=6],LR2SfWR./+Y]/2d#Y]5=
NZ\FCSEE#MIW2Y-Q5#T7bSI1S_#78>g.RCd1GD;5^PO@7=2RfX77MKDK>0A^0D-a
H.A^8a^,dCDQa+9d@a\b-)QBAfZb>)fG8ZP&Q4\Y#/cGT<8XbD0_LZ)Va(R\ZD+@
:7aWGKPAP72(K_N7?PgJ-:HJQC=e_I:fd._K&4;T6c/9D):]X]0E?YXLY-G]@-]S
AZUJMg:.DJF44YK3>\Y^Qb/J,C>ANGNO5&59GU=?bE\N]eX]M33<=[WB2.<@PQNC
eDNBS7@.OG_1MLMS>]5&cQ1Rf9S:(P^)WG>YQP.W1@SDeU-EQE<1DEVNb#)P82I7
8H08;a3\08^Yc;Re4L))UO,?NRX7D(Q6:A<ER_T8YEDEd^:N62E<)c6UeSSb6.MJ
@FO@@M(NP+gaeP#?E&6[5HUJ/5LKDSVg>TI?.J61\KJbWUE_P_@F&b+\EXV=CMX(
gNMQG1]64)fVGW1PQ.6@\V_O2BQf]64:,fDZ:/ZaZeL>HQOY+CI&X3_g]Y)aWfP=
YA/H3cZDDATQW?9a5K-H.Q4fI]>>7PM5\FH9+Z:=M5@04R;,_-D,fAJ]f^CfGG1E
][E<N:VJ222Hb78CfWcA4+&&HCDgK,b(J8Y9gGN=affX&N_Y3_Rf0M.8GYAe^J83
\A&H&<]DbgTS<G^45gI)?F5K)-K6.7<f\#d#=)&LU+Y^FG807&6WKS_:TE@D<gGe
XRE0_La)/X[QK4-UJN>+9/><L+>0V)#IR9)c4HM=UTeU_PfM.f<?))d2A+7Z]RTb
GOb>5.U2.1JD,.17HW=.b_e3WG<M#fK4U,^/#WQ/+[g5;(A(03cRDG@#Q-1)3a^R
5MT&^Oda,)^eZZ&^SE=Cg5d/VfeE&Z4FU_RYKU#+1I83XYL&fV(/d7UFg5cI+E#Y
,VaeGO&QbC[7P_K_.D2>-397Qf&1A?&U\T]=0S=8c.A,[YU.>\TAT0)c6=1IgK]@
[?W;1CZ+/:LW-V#2eR,-_YG.&<]#02Zd\c)3bg8D_Bc\e[J>2NKAQ5TYfdCPN@Q@
ZBH89I7>/)@BZcWVO3MHb,5_Y<J93aWQNA_:^#M/NE^8DEeJ@]@PKBOb3M@1H8d=
[]&cHV;7+7Iga^bH&#-_:FfY&EVd,U_?MVSfKedWR_#c=4004<E[:/#7FZL?d2DJ
=<>O>e&N4K?+?2U?+c]C-1L3#.c26SD.R+Qab>NM3&/;4:RaZ&KeBW9.K#Sf2^N:
@AFHXYVB1Ha\A:6e03W<P\UCH@O+\/PZ9>U4N=>&,L>;Y2S6T)3CV]KX5f/SD>AW
BKP[#YIOg213+bN]=;[=cVO7Fg]9QKH_I0JG^PW]-cUL<HS0F@CZ8./f@/,@[#XW
FZ37),HF7MF](6OMP9-cEKN#[]D>)K=9X(RNC:FL-<E?&g(1gUD]20;)8\AQ\ZD[
fP:9BAL3?\(dGe_^0G<ggH.TCf/.5&V<[C>[[=(J&WcI?2fg#3CeUY2-G+g9-9NU
=G62I@3(N5MHS8X-Y8F:)g3I_V<VFAaYWA)=T=bU,>54W)af+G20\b2SRec^bdI2
O)V19R+75JXBU0UP0<PZRKN[.0DJREdYAB,\-=J@0O_+?:R=#UN.O-<Sa9HK,K4^
)N5HN^RQ4I/,R5A&:da,9]eX;Y690E\cVg33=//.OK5Z_YUDIP?#]6M5aA8cbf>N
P.e>DNH#2G3C)WV71_^_SJD0E&6J@20&BHEW@Q25eC2UZJ>^)[@^0Z0FgW.1P<MP
3TR\5FA8L[a4#L_T@1,d32E]4,65=9>SAc&^<7=;8=CR<8SAY01+f0&5@4&4b;.&
0=G:>IL.@,UQ_gH7O[/R>ac;GS>^3X^](\5DJ0EHY?D>CgUc5a9)T7;1?+RM,a<X
-TO1W5,DR>9ee8]f+F0&F:O9>f8S1CFAK0f<DY@-I@5Z77<?F.:0=f2+VDIL8f^d
DbG/IHD2Z4]B7bO?Z>eY]XS_aI/Y7RSc5Vf<WEPb,=^K5_E^MS<+7EA;2&VU\CZ4
YW8.1J/Z:/,NQ36P,_;Q?G3W7F&,C@1N==IM6++0[4NM5ZKLR-e>Q^/7F#<5<?:>
Q#D\91&#L9)AZB[O)L@0gaE^[bCJ#+GK[eU4aK3H.Jd3:aeR[[Q,>I1-.7SNP@)V
W&4d+&DES9YM)N#B2:C9>0(,FRJ2FNK.bA+QAUX2;aB0K#dB#>P3[@X>XL^Qg-E?
;dc+SG)8,V<XOX6.M9SROIUMeM0.)8?G94c<Fc<ETM_f=W0.TGOCTYFP/P.KFVg(
6Oe58>Mcg)/>WVb@<LX-\/04U,_.g3Od)DZ8MQP\HO6,1?5TP/McZUd[IRdXc(X3
&(LI=GB((YT<]W<+fge,K4Ce^GL4#V>RN7\(DTIZ13)L]4AM;7X4/abIO/bWCAXd
5DfFU6_JVN#+ULU4UNE1cM]@\^GL.<:<7TMd</c)C/(Y?)>+--IE@HeS@cP1WXY7
-TXKXC)b_/Ha\P(5TdY39fg47,RVM6J=VYVaf<Z35F,W+T_UM;:XNZI;)&<<9^Lf
BA0#(Kd/816TVbT+.2O[23T]2NJ0;1D^Md9^N37XI<E_Q5,C7BD<@M.d:1=-8@V(
3gPBe5d=?a3H9M#Jc\ggd-LHU5Z(@+2M(ERYT&L5Q=,07;KeJ5V+Z34>cBJQQRMQ
FO0Ff#XS4T]=.ECWEG6^V]Y?UTOK/\.@4Jb&V/bS,,Y4=S9g=QK6Q#(\=S^b14\=
\7.67f]GRH@S7CZIKdQOW<V[cE-Q&E)#7SC1\,AW=.BBCC<5K\Z_;0cGP89c1gE\
<XCaA-#+,X(&5d@>NN^_P><<R]II=W?[L+O/CT<JI>3?^(cfQOO32KY1QaNF67=.
:WO.2\L(JYRZ>-323C_,_UQ_AU_1CC&\Mc4S7:.\W6WegEWI-NNYF_HL/MJNEW(F
P_X3GI+C#_J9KH9J<,^9&WdH^M7#4H&:DaCbR_J@,6H>SaCO(=gLV.JF^<#94.>9
a&E;7]EX+AH>=[F;./bI<:;?0V7.ZO[.+0WM;\d)_Qg<5Y@U6C4CF8L,0E;=-;c]
J-A:<35d\FQ1#E-A;:K9^__c-9_S#I((??dN_8_Mf[8/1_O3M7cdS5[7FdS1Z\JD
3DH1Tf_;@be^D01^Yg@58DYX/6NR3EbQK]43/H,cK7#S_&]4bI@#=NA&W(T]XE&V
S^F>&;Fb.=b200@&Q)3_&A:fS)WI)J=cG7+N;Z.DaeI7^FV_-A&3J/:8.4^RcBC9
^]K53f>5#](>?(3:G7E+_@,/V_UeUC89,=;5K.6>Z@SQI5RM=\.4;Q1)f=Re?QZI
d5G+eS3@9A[UPFc++9&#Ae_;f\^gQBC0+10^+;ScJO@g>=KMBTF@U9d9R:Jc+<Y)
bGOIS<Ic[L1EI>6H/Zg^((EBg2NYf/JGR(EWT(Q#CS->FD.NIH2_6N][APG]JfJ:
S3Q;3[9ZLXH/-+T,?LLd7/9WQK]G+FJ.2YYBEQ@]P,TM?#14bLVX+c+^;)\UPVUB
W<D(,cMJ;DFISZ4bf/YaV_(^95)a0f7cGD[F=5\WRPGIDP)\c^SV?GfCI^M>7,S9
<C@MWOReM>OC+5KT04U[XX+P8,94X7?EKSaOF^;_&f6&7@_44^1cXfH1:A61RP05
8<a@Z9#NMI@0_L3,@NSB26M^P:&a),U,CPV7K_5-9BS_KQJENb3CMP&4X9?8+9SE
<M1SH]Ag)McBS^)fG>T2b/MYa8?]CHNKcZ/BFW?4].;L)2Y9b]\O\XUALdUVRROC
?=Q9WW6YBIZZ_;&6OQJ)[8/dA.OZKg1fO]B._3X+.U0+=[MZP0ZD_T7aW;JTO\+6
FVc+QL/A#e,8>;OWI@9O)f)HeG,(a?_GB]1)V:D2DS2dCISX\6(XBA]ND[IFJ9W7
-(&DXAO8[/#:(1:ES@O4gMMNV3O]gU9#X5>(H<KNS>g],GEgGa9887C:FLOI6&^V
1ME)@LT&A<c.V01FXEWODD=aLDTL=W(>X+G,g3X(GB2W4cN5K>I,LEd9&U)MD<]f
?:B#(2&4dCT8IYPU0)&\5FEDJ+V(a3ND+_)&-X=]TQQFY,-W2SU:]Z#8AbYKW(EX
+LKf^&W>M6F)9O2X;/;1b+V6_TLZaQKg18NIZBX@JAT=J_,Z(\EK:^JEfAW3MW&R
>4YYB2Cd37_\fZ1X=Uf,BNQW_Ac8[3PRX+5@)CB]_PK7<6X.#XAe/BVaK^RXWIW]
LF,GF:eg_SK2MI_<T6aO(<c3EfRHDK9(dH(3-Y&S;-VJM+J+)3/:f>ZI@)660EL(
DHWA<I3ROR=c3J&=36a9EGUK^4:-\fUa9cSY3MZJ0)5K8VRLg=fU#WL,8UFW4eQE
Cg1g[e1U1W.7-V#V=+X=,X2G^]FTMWOPT[CG.7XEHV.M&5,0O:G/->@H,,4#PQH4
P(fb#GMNV?HKM[d2002PY)0OZBbfO/?YPG=FIP,+V/-_I<ZG2e7_BK2BK+#9Z_=A
B9cPDEf?1=@)RIN:&@GIGBEaQ]0)7O,]W>^]d([0ZA@N;CdD<L-B[_\AZ_a5BJ):
W.J]OUE_?I^C=He#d@(SK&@Ycd2X<6#eFcX6)G2YTP2P<VX&UdQ)^><GR.]?LDWX
B9^YgILT^G)0[WN?NbHX[_TDS.6>0+OB3UBa;BO25MU50W/YePP^8Wf0S6^aQPKZ
P<3e/\3VbUNc?ge_4.N14O]XIISX387TDeG@@RXWU/?aOCOBWBfL=g?O7D7>I>f\
&]=25<PB(BW_?EB)CM:&[#bIGg]>:X)G>)J<^Tf#)>.+_C@2MM2S[L<KYN:cG,@g
+5<ZV>KV(8U1Dc]#0@CFgPA2b1a,L&4E8?M2[=P74N\))IOUM<Kb=F\^]Nfe2)2A
59R,#[B85<25&)c:KX01O)TcP(#)ZeOaI=?D=5Mg_OR#Oc62F(ZBDc.(4]R])bLe
,8VC3@:L79+7]U],YgSfQ4e9K,2X2R2NW&c/;OG\=>V_I9U&CVPa<G\PZ.3)dL,M
d?T.Bb,ZWc3#H^^c]>2O77MZU6Od=e\H)3#UK#JV)<11cOa_bVW&M<]R1NeFJF3T
OAA\R02@G\1cQ/2B0MTOC^O2/RR>]0fE<>cMK)Q(^/1.;OYAP7^cNZ&2Q03Q69R4
KGJP6?a^DO71FOI8JPg#Sf;gQ5=(.I;?54Xc&50H,6,QX_faG<D=f<.SE,3Ee_W^
^8]=K:CdEQ]MJ=C]Qb=a(Q#I:H4_&caGL<g&694\1#?cNQb2Y=CG7DQ+4:I+MH](
4H.fK,&DFOAGQ(95.3?_.bVVAQ5):-O487,]PS6=[@gXEBgP_142+Y)J16C>J7@7
W,bBcTTKd]If8ACJNJLJ8=R^HJ:;?HfeRKQVNMGQ2=/W&^<JYX60RJ?T:\D9b<DW
R=:IPXSa2]P;1JDLUY;_F7QbO7=AHL?K5efNUR(FRR5VRJQE6K9[N0,S\C&Wcb<(
de?c4RUIW:aO^CbFM+;2P(<gg^7f\Y0+(;0Q]^YQM&eM9gD4PWSB8=&F,#GBg?Se
G5I.?^UBf3),9/.L+Q:aI(J<NO?)b,Ze45>^X8LZ0<&5(5S=SVGRV_1gH/MGJBMF
-]LgFAE9//#@DE&56fLaO<_eIc,TcP-7:T&gFP/#W:GMI<>104RdNAE<(M[[FX96
391&_+005EDaIf8(HEKa]d:bLN\VVZA#QM7GFG8&IK55\CT<F,OQ-22AZ6?DF([:
F/1-)5VVJ#UeVeMCA+e&?X3XEORC/YXDF5^V2IdSU7PE_Z]#M+c3A0R8gJDH6#<K
Ub#5\:+L20)2Pe<W=_=D6F0H//\#7+JIM84DT3<(]E(Z4<B6IZ>9?((Pg)<WGVTH
4ET<<+3>d^GMQ,4B.6,c2geEP1+cOY#;VfKYe5X)+MV&RF+fR>M?c)<RWTL?aM^O
&P)ObK8Xa6/-4TcVZa)B_73XdQ)dI/9e3G76B)dBBe-URMMG,UfS\8XI^=:.46Zd
gc\/C;EKY=g=FIAHN_+@4WHR;L]eZOSFVYI+H8c]THH\K.56[HeMAIS]g,CSA;\H
9B>O)8aRZ:.c1B35;Tc085b==)7BB;gc+A;=bL:,O^+\d</=fB#+_f2gJ.).57;^
A)2).(D37>R#b4_?/=EbSC2_KKDPI3O>GQ:.I@&QZ(6PIIVfHVTbWT3)1#R@8QM6
0.b5#F/Wg<VCdf7R:a?R(Ye04G7IDFK3UE=X8C.XO055W6dEURU9I,fHf>7=JU3G
>U#,e?+dAVOW>3\?XGNc)eZ?8cK7T9KY9_?Qe@Y,:?<,LR>U&-)KT_EGd\&?V0VY
-Q\OX]M6@b[/,?Z_PO@?>3>N_Y&G1#>J0PA_P2fcY?KI8D;4IP8JLJ54S5#3?UG4
;16^K.(XTa,<cf\T8?#>@Z&XL+4IPE5T9ARg)A8AbID<V\1284I&a:>:J]OE364W
,5dRRT)fNYgeXDS4)?YVeSKGSC88CAY;9R;FP>L<4?d3,CI/&E79S=5(@MYD?&(_
g>WcT<VLTF0+[aY-DP(LFeQPT(NG&[RfQLC^bBQ^X2_VZBL7CU(R6@FST21&-773
/.C_QX3ETW(@/RQE#12OI=--U\;.KHGT&K.?D::9:X]dQ>aGLZ=T49\PMd/O9BI-
gYDQ_ROQEDQAXJ<HX:1T7W?AdE4&Q+>HfcQJDeI:Dc>ga10LV8a<Z8JAV)8\PTBW
9L3SY5X+Q?H>eJEG[e&CMDc1Vc7I5@;a4-2B(5GV>(f8UNE5^CeU-CYG9<_8,LUL
ZJ=HL]GA+K2e>H-Kd/E#b0#Vc(;S</=_fBPL,_<7H_4a2M7ME:6<UOa..b;.Z.A0
DSXS))(@.YW+N\aFOd?2@bGOW[7]?<RaJXTKffCMKQ54;gA#_gNcKc-#e:X6;B09
,CY^K17OL3Y.YP8[NTMBMX&3f-cRN=^JQ>QW-M\/3HO7,_:M?2)?aObQIg>CX#Pc
T9,3798>AIT5ZQdS8(_83H9/)[N]Y\Gf_73.NY9ED/6(f.]XP==MbPL3L[3=CZ^+
Tf51#@.I4:BeRLY=^0OH-^A];2QCFcTA&b#a.MTSP-XFS1?ReVKDHPQc]<#F):NA
V-fF;DKaU-=&=Jd#E6Q4H9N,ee^4+^c12MYN-.O@+(bL?I[6gHe7F\MZY&\4e[U#
;M:TPU8A=XQ;c:#Yd^e)X@AY2Y>_F#O1#RJdb[QgMb;&EXI5M^g#UVBQO[RZ,UQN
KGM:6>;2)GR:)E+M7,<8&.c(1eM=?RC2R1/.V[53Q#U5b&b58FbgNg>RcNC2gDYH
a\P[J(gf8Y#IJ4A)(Q_<0IY-4^I12U47cBAJabD5?f?9#d8(4Xc5E;9I([4\)^U9
N_TY++[I:bSLV5d]NS=/AG33W>>A;TLY7D00X0+-_2f=/g1QH_U,BF]\KV29+H\V
>b/2X8Y\6:=+g5ULQXN:V&G#)X&TEY8U^?HFfJWC)HDV83Q\HG0?\g7]0^VV#gID
?0_1,1Z_8@ZW.^P-FcT^c:5JRJ:V]1@^6>9KF7@+4X,XWcWe;GC:WA/M?.QPU\JE
R<;EdPRb?&.ELPa[.e^cWE/\<NVg0QG\4@S<F6L6GL3LDD;]//[D_\)IWN)We1ZL
bOTFI=_cVL>?HS@]=1?>\.8R+I8N4V.BG1e6W9,Zf7X^T^G_RNU,(PUUR#W3BZI0
c;M?<#MfC1E25=X++?9\P4NWH=T]RFf4HP19M:S;aE(Z],#^5.PaXW(@Y[FO#a@M
^J-@;@-A[?#EZCRg^-GH^N4M:]\67.S4+\<,X&4U,^V/O6JD0@RI.4F/^5)dINYY
#a(9KUA.J8AVUDI25#8=:<Z^H9Y8&G+>ZHd?4)[,SXJ0_K94K:>RLRP#S;+Y0Xe7
ZEfKU)HU_UMf##T;[>KIB@EDB\a.T^bdaLZJW&<Oe;?)B5&Q[PL-daJ1FN38@\Xa
cD:DLN-\W,Fbg)98T;9?P2fQ[MU4;;R@(RB-:EZB_F]-?]a)XB(L(@OXa8#^1?:X
.95?QF6AZC^YUI:CB^#\G+2,MQgDGg4(D5H^Ueb::4&f/[RF9QK?fV<7OQZ^^?b8
2MK>@D>eDe8.4/S0;5ZO,PC.[.Q&ZQ1;Df>>S?W\[84[]4cBYQbgTVeW?IXbbYXF
YK.I4/eB-^aLW1+U4^,5CP,g\V;MNS;##ZeRNU+6?WZdKME<R/?Z0(:,XM&FQC2#
NgbV70aW=8)0QG_O6V+UAVLR8Y_NdX-G0RGD3L9PAc4OKUEd(8\T]?BEgTZ\Uf.b
3+;:6#7RWHZ:Oe5ZAe2]2XK;CV&]3?UI2Q3dU;Ed4O909;ORE#.@0W_IB9@D^T+K
YR;K2<Y:?eY^7b6;D#Tfd(A4,T&&)9HLA88,J@fS18)fR3?_c7b.0<9IV(5.d-3H
3S=L;9OC>()VYO+S6QL-aUE6ZR@M_<-VG66K4L(@I&H2>.O)E@:GNeHBbC&X0O:W
::0SV+BWgM.4ePNP<OF6:D9RIZgX73&NSZ)UZ1+?@-b\-G#f?/Q.@)a-P=XP8IP1
<d/+fTN1+-PY>OGd05&A?<fWbB)+0JVKTX-/:c_4/1.(LfHb.@fPS9CF=.b496@4
-K#TOe<EGXC:b6X;aI3NY4=2a^H])^-4IE]D[>WKWYe/E5UNU6dOd;B&T^J)9gXA
dPL&;RUf1-a]]OH?\J5(b#8]2ZAXafXUdPI<OJ;ga^G+U1Ga(D&ITZIA^E;]58eI
WWRLB_<Ef[,+JZE9.Eec>])T;<G3^>.9RfS\3(&;/VBUO,?E]=3V-K=<7TJV4X,6
#.:/SaXSSEU71,G</5BeBXbUB;>KJN]HD;[d&?C&>TYHC7>XGF&d[TKe_>Z\\4+[
=9QUR>A:EJEK,XC=V-@7U)4OR9IZSM@_N)PDY21>40\-YXWU,C0C]FPfFP7M2KSf
\3=O#6(2Cb.&^D_X2]AF?,.f4LL[3T;<,X3#+K1BYbX?XfBD3G.L;c28_JIF9UHF
eRI+T/;7ABTGF<HE#CC;I6F;0V=a7J\aJKJ6OF+;_[0@Y02RQ:=T#SWM[f-D#>Q^
-^)3TTD@0#DOOL?S_FT=eSQ_BJIf7NC<N,(:_9;LbL10eS0,IE=GP;L0,Q-/f<,R
^8MW&UZ3BFX^URCM@]V:FO_bH2CP&Kdb-\>WL-1KD7a\;D1TL),5d?=>C>I)@_KP
-,23_H?G^R8\BA1O=&?Y(2,B<JgcNI]1+,:XK:46V,C4E3d1@N\-NAYUM:K+>)8O
:]&?#f)F7Kf>RIE5IF#3SX@2Gg9?cc#L>>KQOQE+N/EI,C_4YQb(OQMLd<ZN36Mc
@gNUT)7.D/T/GXL?aDdCL6_9X@9\4cD/)NHW4e1URHdS#@GE#GQbF=e[O#bKZVf4
<(R&5)a?-e(D<<.91Z\5b[Z(A&^^FIAV??g.bO(06<7^YIYAJV4VO+d[?O/dDW3M
.V:T5HK4VR2Q=_U:2<8;_1E#M-DH\3@aUd\5L/M]aLbSD+b^G:2D(Y-22JcJ(WDW
\GDOI6AU]IBKZ(N8O,.#)=Wc5A)[[?3W,O_3RCV8:1b2b&,+H6@^[N5N98PKEX<#
Q.H41ZAe\-ED>XW;SWE1M;e9UMLZS1^&&YR<ZV;Oc+AE=O+H^,U=##@8aP[0.VFe
LJ09=F(0+_83a4M0cW?>OW)R,C6L)1I5JE?2P7;@WaMSgIX6Sg865(aN4<3(9^6F
K02XKf(^-YU4>&T_U.dZM_H+Hd?8;\Ce+c0;5A2g\AE&0#dE;IE;3GUR?SFCXaX1
(6-g+[JC2,_R]c,&5ee&=BOYZXQA>&^61e(C>&56C[c99>T3^aad825d.,Wb+T/)
WM9Sec7a:30(U74BOOa9bWba-JDW-Z:HBSVf.<f5d7A?/e=0Ag+bU@Sb9M_eeFH(
5+N.,N8WNRQ(,VJB&U:g;O6EB7g#)<YKRcD8QeZN\TX4_A/\E8<0EJ5\e,#FNEZ1
.(IPNT]K6cFaOS;)WeVS4Kf+#<&J>TSOe]g:2H=1g^J[SR1V:MCWg#(UcBe7.MMJ
2,bH+1OX#8^3JLIVOFDT2J30<+P@+AI7KKg1-#Va-?9:H(W_N@_VcY4.8B49(8U<
KBY(ZR(FMGPS6AP.6F[:,C(T7EH2QL3IU(=_>)L5c(]\T3>3dXV@.-(#cVf.ge?Q
V68[JG#+=(W;;OP8UWa^QP;Y3]d=LQ[KKTSR>(1A\(U73WMLaMB[H+&AK4Lg=Q_0
EVC=V)R-d800L3LDX[E2<&fg#Y:8a0c&0__0b^.A@MN+2KOeVVLU-N6ES^=^[^#a
EOX2TaO(U)QVS+EBP/71F9WgCXUS@d+:E,2EAZ_+;IP,5Me3;)6GaOI]RZ,27F/g
/)dW5Y]IJ#AN0ILZ_dK?a5K[L,N.9OZ0-FKO)>.FLZW:3U4C.A1,(F;PU9P\JJHM
N:_J9K-:>caT:ZBDCD1R:g2.LVa^V;/Q+I0)IGD?B6PQE0a6PF_IcO@cE]5<b[>/
E-EP(O1^L1CWF@<5eS8gDccb3.)(>SMEcCR-6CDZ_ZB;7@d_/SE8de7VF;7VXb)d
=b#bSKb\Q;a&Bd2(H8Q-<c2a^bLZ\ZKJ7OePAPX)ag)8WZcE?,JcZ;[;)aR[IZ(G
71Q4/>#:VJ<)d&Qf:XQ</LQ2P2XK[87+WC]gQ\Na\)-GYFfB3Z8Z.9g(&_<[c8d5
8_Eg&>/H0fVRT;Q@NRGBVUA2L_DUaZ)G+F0@\O-BZI[4F(5EIeLN-TEWABb97T./
L&?I[LRBS.[gV+IceTcU1;]Ee\@eW>)QTDcKR8HfT7DFI1Y>_c;2M3CZ-M_gNHDW
^bS091g?GPf2A_8U^O?2b:b+g<V.g.6bRI(Y/6N2TZ6YPMe[/,eJ0Fc0EM8.YPV+
?;A(a]7NC8;SW-]e]F1:#<HH_9bc#IU,/8dU9[VNO];+YZX/bG4(0HFA/f]HPN+b
E]==D5DNRF7<&F=(A3<dd?=UO#J0.XKRYXM1VQ4/PWT\ZP7(XMC^I-/)c9N.:1Q&
1;M#d3QJM6D>M3YMJFb#g6^eBdDFc1[^L^WGMCF,YBK1C9FJ\0FaB,MR[@84WaTZ
L29+\T>LNM2gL_c/D1G);TY39bf_(1/f]HS&E@(RS/UH.G?NZXEG=YP<,D>R=_9T
>NA4]cL@&5cQ]V+.&2):(RYfC/=;>VX:[?I0c,+==D+^N)FXYN2V]Y+(X5_8HAEI
N8?VCCWI1]T\/LE)JY39,U47=(@Xa;MRK];<-DfKdXW3GOFaegPLWX98C6T[^Y,T
(bRPLeDLc1LeBOOfV>1g?)_eCZa??G^RNgbNO-gV7YcS<4VaLM_OMR29,&#GJ>eJ
)CQS@+]3,Z@XZ4<N3+H(A0J&X[NC@C+S(T07&[.4AM,RJPPGN:@N^\JU.[KWB402
>=+RbF5GD2Kc@;VgE,O^U8#0=]U=4>QA?9AN2_fUXTUY<57#:Y1IK-<);gI4X9)L
\9Q[_fOP<(7-Z1N@4)4CU=H(@QMT-#D47&6?+fDKQ<PE9dXf-PdXP&L>D85@YcZ?
0(Y-D[V<=\R73(b:M9X_,:5;7Z:EU_W9\_=aKQH^IC=KaI0.D/QR9(U^\c.]51>+
Y^7PK3A(X;2Me@[Df&0>&T+U)agKZ+83(RbCe7d,ZTSe<NPQEPAaE@WLVF_KMcaV
5d7DC4<e9RK+F@Ja>O;C=)5O6Q3-Z+JT/]EOd42gS[VRP4UQU/P+1XP_I9gS>UOW
aW,TWB=KU:6K#+-?gBNEb>1fLN5>e05L27eeF],<g&3)9&@)ObQJ#Z>,^&<R0C;U
SDZI4<P0F:WKZ]7NT8(;&X#YM8HD.42CdBZG4cA)O@JbI4\0(U9XN#7N+ZDMU[&,
YN/0\#MB_+B&^7+:<=1PDI3TO/,GEG(X^Oe153FFF(Z/GI&Cg7]Z>P=#bf8eEXFf
W6@I2WWWI<\7]]\[GeCfGP\Me]g^b.#^X5\O:>;RF8CES5)RE;O@(KH;IX/TFT&e
G-NNY71,YG)VVRO,I?VL^W[/A?c,#)MdV&.V(FI0B=Ba8C[@IE7\\0@:9c0J7O-.
?\aCPM\^LUJN-Q]3\J7D1>eL1fF3,EE)g,];g)Z;L_53E27Pc(X,<(&Qf&V@^R-:
cU-(WVd>-((;8c/&]]g=1+gbK+WHJZ#OT4cQ:PFT?GP^<=Ufa=K7&^1ZJRfY\0H/
-2&&#^A2/]QQe<6\D^WG=e&/MVX4[@B+2M5_P>:,I/PLOGICS@L8YGA-D8/HCY>7
2(CCW94F1BJf[c]2^@38#[&9QdTFFCW_AI2IV^@=NA8M8Z]f62,aKDe<I\BEPa,S
98a4(_9O9QKDXLbQG:@[2.#gf;/3Egg]Q@9CS):(&0b6=f@g3]2-]@R;ESQZ]=,O
=W/c]IMbI&RTX8:2N\;3.-7XA>X/fYGYW^]2.X&.=0GR5VPfS0a&M?K.PBPI(-3X
E@\O&,17@4SI#YSO_:#CO&/I<DE@D7CY[T@bE7\^#<TUG0C3202c5<#/7JCQCR:3
0JRe#Z-T,fU(]_+eVAOaJ09()=GKZOEWDbf.3Q+O(/aV.&HBA@^5(,B(Z[9#XY_b
?&UD30:X0+b9WYTJC.c)GPg9@ZNN2/.:621MeSA9(c@PYBL0[@^_QJ>d&=RcbP,\
A\J4aC5XJO+Z4XD6<daP.,81(aX;DMSK<S7#X2^.aY3=;55<.+BJJ/,e0^U+9^&U
V^OPT^;/\a24fb_L2B46U7T<9I-[.<HB,HX4:NcQ3da]MBF&U#+QXF[U3>>):JFD
QHZWUTgd#g:<N+_0GSR.;1Va4MJX)?O6JMLD-J2+&Kb+g-b4>46=eBY-fBN]MW_X
ES@MTSFVCMJCMG1E&]B,0.(eO-0&D]a&)\]+5?J9[T]gBD2S7Wb3aa?SL9,/0UbG
1Z(P#,g.+B#Sd2,0?.>K)WI<>9KLXOB5WWSFY3E3e9dM0^@H)b8\OI5P>9_-Y/OX
>1=.X<CdWM:V,gY7M1KB&>eK4BI+KQO8^__^V)ZVN4LK=0;U^N?a17[J5Ug1]-^Z
ODa6#ca61T&?]9R_&QHM+-[,dg4#U=T^IFO07VaPbK9:>E?e-\ID3BcZPDQBdgI3
\3TEe9+bDPWVW#^a2#00LTKA591+&:SN(b]S^JNA-dG]a[R-S.L7db07CE<JcYG=
DLL[H[gZ@JYaK(?7\.#Y&OU_&._JJB3f=:ZIb24NgUZZ[Z[:DZe.ER@T]/UCg[?8
f0]Cg&2+<UWHP[KVBR]^L@6cOYgf5EZJa8_AS(g77,9ZYc3A8I<9H@M1F[_S5E;8
LC8-gd)I5C#=bWb6Q@NaO9[-2DI\+,<@.0R6^/[aNP1JY3/L.T3eAHS&,=bPb1f,
5DGMgD)[+=IST#<@1d.DT)\65@#8J3ZG&ed?b[1Q73[fI,YO,9&4>#GHReW0EP;/
4&[..L??T9.g+a#>eFIPDU-@#BGZ2,4L1N\bW_e[]C:D):7K071&OUM.(ZW)@gM:
dc7\5.VCSWL[NRA:)7.L,F[.JI6<KH[)42G)1IR_+cC)-5B.?f?B)9A,^GX)I:;2
XBX]+I>/_E&b.;K11dD18F3:Mb)R\Pef=(=f=JY=BTX]?2M@N+XXb>cOR9@_.-8)
;?JgHLF5WQ,6;=LL_FCWgO13AfQ3d7C45YC5;NTGU.c.-_B^5I#O1>3fJaE^8S@W
eg7+P_a>PK(&&8g3WN=_CI(B(45[d#e7IE4EPaS.YQM/LNaN??@:eK7e1N?Ba9;C
?Jd;\O4=Ja7)BXKG[_W9YQ=VQRONBCb2=.b+gC2.[B5Of?dJ-_>3/c#L1d91ZKWL
S0b2Ea1\=1aGI//:g29ME&AJFNF^K^999fC2>C(K-a4,+#)0AFAFPaP^=-S.H)41
1<[9bEX9XW5Dfg[HU/E0Sf9GHZUB:K[Cf:?<A4B>Qa)3PVa;2)]-Kc)1gI714&<H
KF;LT+,KR1CN)I,Ed(J37KQ1)5Gcd_V3(=WBc8.:E+J-]=5&U:N#EITB@HC1\DbM
QJ)4G<I=JC+YdW?=;.X;47,AUM,8-PN.GN;VKZ;NH))C4^5-^R42g&ML-WV&26RP
g>e>B9_V,e1AO(:2c)HCJ81.a4>9NB>I?,9)a5d1aD&E14U30F]L.WZf&[Y9\M,a
Z#ZO/R[@<SRSOI[cEP)+=LdgWH_5:aH?f8T^dc>M>a]Z=5<5HG[Yf^3)UHRC<1_^
]2f1//^GL#2J^,;14PUS:,?QE.0RMR7KD-fDAEVV6=:CG5EWZ@>XFU6Egb?F\@eZ
O9-L(_Ic^Kb)@9\KdbB.ZQ>,P+EONH][ZMU?ZLM->+5ZaYX]Qb^<-T6G&KeSADZB
-0c3O[11WH]:0?I@W_IN^I:;Ac2fa4&2J73;#A;eacT+J=0XaNc#,I9<dY//L9\V
P6#DK+:efK/e.gfGf8YN>1^MVPd:eC7][H#]]7dSD6F0]1T@Y41J:PM36CRI6^Ic
_WLWC6A0\.c7\ceN-H4QY-MN/\QY;M4EZg+3+0GOg_KQ,SD3Ae]e8FB[e64&0XdQ
&-+gQ-:0]JEbUL05Qa#_Y3]/?[:VZ)da_ZEMKLg8-<)O]Ge/<1=f-]-T/<K_U?/N
J#+/VCTa:#F]c6V>.(^Ya:8^Z1RcZP0,SM8[EZ-F01b>+YS[?-N?,R6^C^LN_#S2
NK-aDOY.C)6&LdGZ\8+^97W>U>[A7:eYbKUD3@E09._Z4:@3K:70T1>[&NO5Y:@_
->G:DB];.?=2XBAL[Yd7MRHWP256+R#,8WQF\TW__DE[ERK/^/^K<)TV2]BHQ;IN
AQ[A\:&\VO)0)B<PF8YUA@,;K@QB4S\:d<,IUSEU2e4-)c;PH>b@#V_AQ_44A8F.
a5.LaXESgD#ASbY=,S)N2Tcc9I0IVbb-G.B4Uce0bGKCb<^HUM9Sf6R2c._X4PCA
,;WKG[]N_5SCYGJdYgAA_2QIe9+^;&aE.e0=6XTCb>;)d67G=QQNUYedGZ+B\d>=
MR6C>8LMJTE6Z&fA8FZ9W:5(g352F8dd_=_:IGIF)FL&LPe_/WK^Y^G)_>g^WYW4
>R,Y?Q@U92@P+^9=TJ,gb,\+(/L\:3]Tc]AH+&Q:[e6a+?R6?@TfE<d^-T+c:51C
7&8)P6fdA,SMI7b+KJKFbDT.N/V^/G=A/_>QCBgYKP;g]_JT3HI?BdO=5<D>D]/@
[&4>BefU=(K<?6#N^0_L.a&WQ6bEDdXPZAM7+D]Y5eM-ZQ<]P16DCW9+2g16[;Xd
MZ8OPFH(TOZ?Z.\aD/(eE+BcXLb=0f\/0:6JBXLJ219T3M_>1Z0[7E,_Y[<2N09B
3?b6#R&\KcILf1.ZP3IWI-45aL),VM0IIDS<cZ2IaJ[64Y,:d;(5LQK(:8>6H/9=
B9X6;&OCKR>15;S@^WW/VT1TU&V+<3>a>+Z_^.L,f_PUM_+BLI^IGW>aH3@L6.R]
ZXTSFG<-S=Rg-fYO9_,@UC-<c+UNK-08efR,A\^O8XVM6F?3UV:@fX_8..@c:S0S
,[S,:L/NUWO]BbP5^M_NF#K_&OI/6>/?NWNLW1,]\RVO5>X:IXgDLFULK?5PAa_X
6)#MVeb3VM>d?6ZR?6Kb#a+8^R&H1:PGFDZ32a(KbTV&R<UQZe(S<E5[8K/_ZN](
^^<YB7.]T9]a,f/KFeCDF##a=,,HGEMNC3B0AgdQYL8F@JUS0Yg[d?cc2:&POd:_
)_8>[UKS\#e(X<W+cNG(\+Z_aGM@e3IGW+H@Wb;PI1\J9,#&S&^,&@SRK-,0IQT#
_5G^P^7EZA,D?PZd^65Z-8b&L_PYBa4ESZO9ccU?)DX-\f>F=e9^<>ca>8V/+;7#
5:S(4RHHG?K:f3K77E.@F>IIIfOTP+RdL3RMP:Cc#M@BL57T,+[4W07;#2Ka<LQY
+M7);1Kd5YAVME6ASFS0N_(HZd-;XMBdA)6P8MF34R(J_G#+7a:[MAYe+d4J2e1O
-#\D14eNYd:dcB:^).AcWSCRQ9@Y<aY?U&-]Ab]7L_3],)G3B<VeQCD?\+IZBG2a
_f+FBZN[P>ENZOOVB1:K@eE0,/P+E1bg:Q@L4-Ba,Q<7B@(Gd#J)BM3</UfU<\[#
aUS_6W&(H(?gA+\9R4L?>76c55O^T4O-I21WU<T^1)HMLN:<5AU>\2CO8.gU2B7(
0b(\ePCK-H,OU;,_NbR+gEZO&dPc0.AAT&;DU5bYFV7\.((SJ\2)BYVAe=UU(#2P
1bCQ5BB.S)(.B+JB7?XD9IZZfOBIAS-D:XG2Gf)BF(O<Z;O7MOF(aT.3#.2:V3bH
TF\d=WW8&.QS..<\FgGE9MYC4@<-a5D78W]YeU#(=\_U2XZ@>3=cG<?O-2M),7>M
NV3g9Zc7.<8AP4_PE-DMgQ]G,=T#1NOMabId8T4MD;-CYPe@N,,aY<XQLB#\d7&N
KP8?G>?[I=7U/T4[<e,bVYC0Qe,RH57@R#c68c0>U@L8b4IfMgJ+P=X6fd@G3Sed
#Kb<V]c-D0(3/SaS4<0YJ\ZZ<c88Y^2]?QV7;RP0QLZT3b1Y+L=[_EN@fMZ8^-_Q
]]MFPS3>_CPa^E;S6EHb\<2UMVa+6=g,5D>F>Vb@0:,7;ULC4VP-EL/\Cc[W_N.a
cG.#Xg1K/,3J,AH,&1_V;-VH>Nb5ADVLV-cMAC,;A\J&-APBH0EfRT84Nf,.?\=B
AMUZI54ZV89H+6#Yg&V\FQH+@2N8SMX)C0TJZ5Z=&/VZARSFOVO6T^Q=\;I4],VO
e0DfARNHB///NL+HD13+#V^7)K4S0.4&J1a(7f&0:,<2/TL7HG2Jeb;/Bd)O1C:8
JGV<HGZJ9(,WEA6fZ3-IH:KO<7Og-4W^efDV7#.4daU2[gMN8528_2X49X:3c:>_
Hb+;-Q/YE)f7N?d1g^f2^KJ7Fd/Z3g@CQTX#Bd_IN31e:_F++I?+>B^/696AR90+
gUSOC#J(F-/A555g?F.^V5X.QXECXPZ?;1HgdMBBf??@HPd&5?F52=He\VB-=:@f
^[,b1HE[#;EM7LN(>P6Z\cYR;-44C5e&L88E4@#Z<@V[6_L;H03LafY-(J(Q0N-C
?.7Jb1^VZBY=<CC6FS/YUJ8C1/0P99G(GId#70>?VX0(VQ3P(6R8)+2MLdRF97?\
)W8?V5<(f9?W.HRC@37\.K34K)e=b92/XSIE47@<,Kg_L0@5O\28.M\J&B.Tb?T9
^SE1dW.DUY6PMeEJ2Lb_O_Qe-ZD&+#9PWHD5e-IeENS2<4+C;KPF2^_d,NW=.(?W
IYA]WMW_^[#ZSEG/W?3,-Oe/d(bJ@24GcCQX.<b(_.f4+E33BBE(a\^6dgHZGc(<
B\ODD12[+IN>&5-eD3JV<?TH?b+/fR2IVT788R^WE3HCVM,=/(>8__WLV0)K@)Y@
A^UZ<@gZ;Yf@>99.;46=0[YHEIN1\:.46BSYW>aLRB?Te@IN@\DFa[JF7;K<6>a1
_JHVPbTCY9SUd7F:?F\(WQ-@/N:20DCU);a(3-Y6Y/3O2>,#;X.?8eeI>)\Mb?b[
cd\J[-FIUd&(_&&af^.a5QZS;P;X[P=<68_1+/N<D7]EMdBb<G=)18CB<K)5eW#&
CG>0?0aU)MD)dJSB,+d>31JTaG=<Q1c#+DYVDdE]g^^_K0(P>C(E.Q2^\2KNO9KB
6GUU5+b[KJRb=1D^,D_+#Z)b.PB+BKW]SS_YdR&]dVJARgCVYa<JPLAd;0.5R-,F
fc?bN7SW</^FIZ9Q^<MB+N_TB+RSOd8ZF7Pd:]^dagQB/,:GefSJ^C39>41:9Y&E
[c^DJ38=<9;^;T:416PUSZ:S<MR45+2>,9HgGM=35Le_+)A-&H_F1G)+\.I>0,cO
eQ:SY(>PdgaL^)^7Y(.0NJ6I@Z:>Fd421&Z&N6&NfbNg^&cW,O+@]RLUD<.IPaIg
fM=DAA5P4LA4J[WU0=(]B+ZECH)Ca6&EHVGPRZaBIU=Y2Z7WdQXa/GB3F].R_bGP
D2L)C3IC]QE7<Y.O_4T_L4=Q0=Wa>&@QHJT=7;^d5UT[O@[F]?=Ye&69+F=SAW&I
C.2=:7YI#/6-1cId[W#(9]44Fb>ZDX8YH^=3(VLO^AAecMXJ].ZfA.Ug\,/S@819
/CR_])OJQ[]@>Z,3eRCRB8,cVX&D_L>E8UG-d90S4IUPeB.MEGAAYM2=@K9c+>K:
E6>LKb>WgPQbE=/_&.SeS;JdTMg+cP2e+5Y+-(AZ-X(4XIcQ=Y)9^d?#BW71];MK
gJ-J9C\[aCa4NQU>\DCVBg=TbI]cXV4,>>=-e@;cc;g9e_U?b[)a\gISb;8Tf1T7
LZ+><c7/>;N0<[7(9\X@/ZES#Y0:b(&@6;UVEIJ)U+TW)J4_[@-1[#4JA[XXe&Lb
[:BELFQ70EU_Z[.N[S:AZ?T_4A5UVB0+29M1)a4C&B_c3GW(.b,#^0^6Ua]^[UU-
S255ZE@,e_g37N3<4:WO6_7S\RCX_D[9g<?dYf-=HBX,].KG/NT]WEY0);gK-<gB
A32Eb#addRN<)JN21>ga[QV9(/RY6.]D5>a<^[=QM@7DVCYT4^)ODXITa.]5-Z?9
/[H16-1YX)6METS51&)g/5,FD=QUM1QTDBELTe+bBS#;3JH&PGfacQ[F#185]#Q>
c74aMHC(&ZPB-b1OIJ^UU^a[ZE(:c[.,;UQ49e1=6TQU?KW9T,,QQHTg4=320e=H
6-C>I\4e^)&GDJJ(WFT9J=(Q.8-&&ISB0L_B4V<E-f_C3a2FQ@TaSJTN+c7/PE6g
PBHWP@f=X0X2PD3ZP[\S5J32:@7LKgDbRa>T2c(<AFAP+IT^I>WGD3Cf5aE/<XbG
O?_cB-<.@A:S#HLaFb@,XgM8BPN[F<&Y(M9.,@2K&7C(5DFg[;^PAWW=83\_BQG^
gLE4Y.(>C2&VfC=<N-X36\@cO(_R:QZdQD.c(79.KfGN?YM3TKdZ+@J3]C.:P)6Z
>#d2@B=NH.S4B;I6=K5ZEZEBAM^<4Xg-\f&@84(R88A4J3&dBKg(7YX1V+RdEU[K
S4d#T>&UO[K?f34AZ8(S:^<_#b7>.QU^3\&6)MJgBO47d(\-OVc<90cGS;Y;8DC(
MUL6KCO^&WFG]O[c[S)e:N2]<,cP8JRB&b&f>:fG^S9OW60g@OGOa1-O<]3fTU12
K0aa5ed\&I;e02W@#CAdR?bR9<P2OZN,C;^8PCOedb\71ZJ76a5K/=Q)4DSA#RKS
P\;;.8Rd[?&:?+)d)G0YK@H3/3(H2g@-0P]Ea];88;Vc+Q\0(e]1.8a0EN_[7RRL
)aNe&G9XC<MEM:X9QKTFAQMHd:H:(N8^-QDc+W>1GY0,@Y++>/B<f&T,QdD<+<Q>
e(3>9Lf)Q70#+6&+E;7HOY+\XCZ:7<W:\K<:R0DRLP0)\UM\F<)39-[-/6-T&R7E
K^-MWT)IV1E-LQO-e[[V5S29b.+5B;O]+I\JVCIIV(YUdD:RJ?_GY)X3fObYaI@P
3K#YJB_COIS;CK&9EI6U[]VcMH7=-;.NP5LCM1c\2-0:U7G44aaaB5]WaF[R(M;O
KNfLD7\1&#[85TQ(CIA>Lbc>JYOLB:9WX+_.9-K36AA@8=NR26.=2#W:dYHM7)aK
beOTK2C.;&WF\4\#W@:c)P]CI>:T4F<?A2V^:AZKKBM=#2d1afVJMS,T\W99>=(A
22U?69C.E>+B2>>RHcA8W+2G:6(.OA(fF&S]JO@XL&f4X6NHYd8=7N^RE698dE4K
]/3^@_RP>LH@&OFXN/NXH/_,1E2\C4IQ8Me^]Z6YR3#2++TRI?OH;4<HW@;NR8gN
(.@ff__^9\VX=]dX-_3KCeU-eX:\HIH?d9WT?VTD&?49_>BDUdB.9>1DcfJa@BT]
O^M^a?B4(=DU^BPCJ?DP8T#I:HU1,WZ(EMZVIbDN&X[J84YbdBJ/SL6QYU;1O)AA
d32128QLc5D]:0CTJ-14.2g[aVa\J#+;LW?_OD0WZ66M0I<(8KN;#,;a8=35ObK^
L?SMZfTSFg^N1\aW.9eg<8A78PD\WdW(3;+>T/K(B=YXf?IE2YHJUK(JX8Vg]P2^
:2#<NC#gK&<G@O[1\@.OBPUX[>UWd_7fJgJ1aU+HUH#PNFP:]>L)+f>aV23KG&->
I4YTS;JdY=;V&4UeA[-7]@FO06KR@AF#aP7B(KZ+@Z<I4QON\X2M#P-?ZO5^DU\/
\;VbYAA7=bAE5c3;;BE#[aVJ@L1X?,719DGUD<89@>[<MT0</F^DR90,S4908cbD
+AN1N>IIeRO@ORHD-Qd;D69/aWF+H:5O>H@MA>7<]HU2c76=Q0WeG&2A5KX)T)d]
7BL3&IH#4BB&_6g4KWD[Oc=,&0SSLF6>-[Y-b).#Qc&&Ud&f7^)=,#OC]V.JD\WX
]OR&2W&_N4,KeFY=,6=Z.gACTg+]=VVT[f;&,6agA+<E9gG=(:>/2d[DPM&_AN&]
>KK&dS2E(;e=LI]V^)RV&VKRVY>>_/O\-W3bQe1-0I<VWVW\IN:eg,66LU7A?+=-
#XR-F6c@IB)TbDWGf@U^/NcaB1?9Se?E<W2,C:ec:NaZgLX:cZV5-;FE2ME#^#9D
6=//Xc/;3&C^EOdMcS+/]=XU/:dZ4[\6MCb=CNA2-R:RNgQHH+TN.J.2P<O-UI\C
=DM]aOIbSaYXVY[c-Qd]=HB\c84Hgg-C5@L/@M^?B2T_Cf9[Z//U.S1ZO8^41OfS
WC+J,>IKBEP,0,T6#-9\F3;H_KOFVe6.6?:>F(_YYD.8;T.fYF2F^VML,KT+ae/U
S\;&46LZ2S>:TN9>QFaP_2?a]@1(/Y-,abUXI:_\:[F\<.<d_9:/5W+^=Sb:Ga-]
L>NX@OK^NW)6F]DJEeP>[H^K:QbWH&LS4[,SL]\?_\,,C49?+\1,P6;20daVc5P>
@&WO7NGNG9ZMFfE5Kg[XJ0B1AJ9GCg7]&T@+LBeYWX#VG:d^\8QHJD#^3cAYE)Ea
-P,#^;CaYNY/RO=1LWFK;O3CZHWP/Q#<KMN:O13-LF@6OCB9H33AK7aR>>40d3G+
)@a\PgZO1Y@-+S@X.W@8dCG3g019e5+=aUZ6c)R7^]_-:YTca=TC\6V09?Z/]bB;
99;O>00OG.AZBT6ebH_JF3[c_dE\c7R2B3><1MM.eW@N:/FZC\I?[)0EO=4TZUN;
MO6KIgY/Y)FSWH.<N8_N+/(ceBMXU=_WWJ,#WZd7DcLb-(gPN1?FNC-A2K@MF._8
(51d4#cXX&)HH,F&+BG91@<[X./P6[gcYK)Z[2>c;:5C=8;\#EN@60<=-.(ZV5#(
83e_KWR=\gWKfG@9YHc5b0PU)E/#>/Q#QW6_fE1Q6/=^&7dJ=QNf/627?=ITdUX2
PTF>ZJUTRH>C_)/,,GQ\MY,1C9PVC-ad1]A<L9Z4-8EfSZU5\YC]_O4ZabYOTe:f
0M08b^3PG_a0@GP/:;K5SP)#?S&R\=A5>adgBCP,WFSKd]>b?3d1>/TGMM#N1_dd
96XWG3?UJ6cd#4/5\7/XbTY:0XPT/PKK_EJ)F=B-2gedRU/,DWAR7.?SRO;NH,+&
K2+#:;gK7d8bKBUXO#OE73E7LO/Q)/RYfS,TF9MT5RWUF][ZfE+KREN8YJ(VY^Ma
COG:dXV#>gL^Idca0#cRg]K?/7Y)]&a68eD6P8KXL_(N-123+WR)gZaXgH:<.\+d
81=2>+dS-6EK+4U(.5A@XTU5-MTcAD[Q6YA)6/.JP?6)M1efB=VK=-JX+Z:QgC@L
=2V)&N<ZAPQdE#FgA3<Y4<TDF]TfZ1F?GO1>E[4ZIRE?=AJ9@1b7T/ZO7(FUEC>Y
AV?C]B6EbG(U07W7).3KN#5FZ^g[92f\#aL=M1^ZE(1(.g#0aCA]M)2Ze;[c<4-B
T#Ug[?8(F<,BAYd2GVMHD0X+AdVK,OA>>,5N\D^Y7#R3,7eVdSc>+RCS&\9f@6Je
>QPI#;@BKFKeJ:8L0.GREW84K\KWF?8AAePW+C0&O95ScS1#I?RR;06IUe-876@d
+#G0AW_9BQ:_9TS)>U?WC2\Te5EOcX8e?fF=#,Mb.0/2:f]OWQR<=+.C_9R6:B(H
\)IMN2f=2e6RPA/Fdc-V@WACB>>#Ng-62YZHHP8G;3QQ4HVVNe/U>c+XCQ9-dV=,
H+7e7@#eF/bF<6Ka(L2=B:BRVeX?F05b>@b+?(K(ZCOYA6_(?dS8M.fdL84CI46g
,;U,/Fa1HW),^SYO4W,D@^SFA=KN,-@-eF]1QN@:8YCR>VJO\6SOKMfcLN0?M@P2
Qa_?a3?XXFCN:HHG1CHK3HV.K,.+F<3a9,EWF@/CGZ+YPT@:gV.\_BeN,->DFL^0
@63PE<A@b.NJX1Ue5EMM=Zc0McAE;RY#I<Jf-6g3O[,0=YH4I-@/PY(]1=A(WV,.
J6;XCZOVF5.aW6Cg[ESJ:6<&^b6::b,U@W5)EBIa+=(>Y0_\aQFN(DM,;\-9T_&:
^VN;KXe-f,(6+_E6]ILO.^PM\FW2>;LaH9X=Of[H1<:Zb:&4&YU-8NU1\BYeV6B[
TY4Z2S.\98OQ.<BE.0geYE(<NGA4O,Q5(P5PJZ/W::dDd_^fN6NMd8#1DC;fc0Q[
B]f5=_,^PHRQ33/Lf//_5Yd\<K]HX+Daf\=Ub?&/MdLAd^.6=H0LN?.>2dd88eM.
L50[B+8Zd;W[GG;XP8)0TRYQ_DQW=EW)S=?6BZ8?+ML.Sc2A0VICL=O0&bGc>=0]
I+[K.+f-fW++E<1ATQPDI@G[;7//)-.dbW^fOM8Rg_b7ZC6b;,=CUO.?_&9-0F6(
d:T:GK-AMW,QZQ9;0@<bSEGbb28Q4Q,RCaVD0B@;R#C9aMD)/[[\3=SAQg455C<c
@<A4LUfE@\dD8^V&9=<N1-EcO)39QB+-gRdc4M\-D?HS97Cc.aH..3fbYWLBg.Za
caH-)EagQO_=^E.@X[XQ>:_ZYeET<_0:Cc3@[FLQ-Y-R,^(S:QHU<S.&5SU;R/UX
>(_\&[RcRfTaR4YRVFCC,S;HfX8JK#f)-f/1YQ)4?-fD]7Z-?\Wa<cBVM,8Ia&N=
1M^3]DU34[g)3DQ[8e.TA<:WGRCK>cVEC#4:(&):B3H^C#NAdM.@4\4[]7XRJS3a
A>-1C7LPRVeW0E?E31Mc9B,NT@U^U_=Q1d593V]T/CeB@1Qc2:7@M7FN[HeaY]Ra
f4MgERa5P[gU1A2F_)=d#G<bfDQ<8P)T+JL;0DN_9Gd.)=W12C]8fAPM2b\\9Oe5
Zc?=KJgCGc=6359&bUVA?_-\-2(&C5;UNBTC@\2[#a9d\9/YB67FNHQb?)YEaZA5
([Jd99QXH]78]+@Z[44a/B,c8[2YJTXcNgOP^1/3.;TYH8U2<)Y7YYH5)@dK^H6E
9DM0f:R>.Q9+1[g.W(@:baf(46?I-Q>QEV6fK0bB7(eUBI)e#LQG[e9)X83g/P_+
,PIgP.WD\E/817:D&bI&W>@]RNNA29;@[99W,EI@8_<O??>&3K-b&DB-A<2QN^T6
\=<b#I=TU(&a_YHQ#dE>KeS6341)BC-[HI5K1E??Z6.TS)X=;SA;,4[QG?Bb>(M8
UHddI@GJ31X8?d.dNC[Y^+EIPfd1gY;&AM2]eIaP/OK-)^7GKLed+G@FaXbI(NSY
.1:JAf(=P(P@4&Nf[OZ7Y)75_=2L#/MY>@54G][.Z0DBf#Af8gC5]#I4GE.62^-)
F<Z1-)b:<aJ5KSd0<B,b#E#C_Y:G8=8\/]ZBN//&O9(4=DLT,f(?:SWYUKU;2#H-
H1-1Z6>5J6YY=5\0.K_@P40?8=^:dA6Y[4OG9]B1a/aH]3=eHIgJUW7_Acb-f&3J
bX:S=8KG<fcB\8O;;Ie?GDQI.(#6:d;2HY()Cgcb[]ZWOTRK[Q-d/@b9T;\^P[/b
-38OLMARX3R6NJV.<&G0NPJO8JP4P732=M.[9@UEcfQU&K,caLW>DTUB6QF#V)M&
[C)gZDcDV0;QCMgP3V8cb>>;f;b+3(>4>TJLN0MG#V](JUJ)KLd7SD[Lg[GNYV=N
G0\LQ[NRYWE9Ac?82A&N<#JI5)5F@:Q_J6,3Y;7ZR]<A#(4D?E<2T?\LaW16-cbd
IE.YIaa4Y:?XddUC.TaSQcVHb-2OHLBeQI3cNXD+QLNe1VP0BUP=0\;V,T707e._
V(C=AFS<85QR?TV[eVK[JQc7@?<XD+<e\YVK]6J7WM[D^W3:eGM++<WD/YcSET=N
MRLTBPW;>d@KHG6VeP\L(6CH7+dF2=D^4YMdc3WK>0b/9RPAS-L[ASQ)PRFJ1J;U
M#d_,\W&SEJWW0<#/50M]_ZH,YZZ2U/\J:b^(HHdDc>bS/]2Hg5O\FdZO9=+<X0O
YIA12LD?PC=.WBO/.62?B6K@)@RR+-A^84P2YNQF=Ff\dBLK.^_]>\78fA?EgE>&
3ZJJ[/2dJe7;0<?>FT_XLSO:Ab0dJ,\U<PYBOXI3N=W-OF(d8WaE66cU5cG02E1N
#3YC7cMU_P8I0KKIX?RR@\[,6Bfg+3=AaDa^8,cDJTFAd6&aK],&_DJ@1CG&;H_7
@2,7:H(FB6\RNW4]UfQdXFP+&gL6U9;bfC3OE[W(.\U[Q>K)-RTW478-2fU7P-9?
8eG+5YLC0QF>/XLJ;(MeOZg<<CS-=C@F/-7.78H#_bd-[=.7AFY(Q01VbO[N3S1J
c^8<T#40_):5Df@/Cc2<gWQ1@7(WTU]g(E^CCgaQH]dc8a)_1K/AEFJY5=Wbc-T<
M\FJ=?bU_R>X]][S3b9K8BaIbfFD)GJ=6FH=L][[/(7d1_01AYKdNOG+8/g&Sd24
/\W6R)dO+E4W2L349eGB&+JG<O;1:@J5]#1gDLGMD^RO:?RR_e3c;c/N,@P\VLEO
UI,6,CJA6fag.QPE53)0+E2+B?6>=.J^#3MT.C]HY.4>B.9_[^/;IH?@D:?]47V?
U^DTc/SB1X4gXVE@/ETLEG\;##9S9SO65/@a]]B77?IIeKa#?1)?]7>_KgGM)=(9
ZdCIU5]?PH:/LR+bSS.W#P^GBPFEAZc:8#I97C@Y<ET)^^STWAO0,<Y=<af]B/NH
;.#)60ZE3B#RUb?9eQ3F_[0#gS\f^d\#Z[6,I/82?e5d=]>.4+U3V#)HJXK6b=DQ
H4R(WU,O_9OE7W1FI)UH5^=\E\gCYHLHCEWeVYY]Gc;GgMS8GB+gQ85>S\Vg(gbe
HX=(O)HAE2DV:AY]C8;MI^KX;ECD.36.PU0d;#;IMC^\]dXKE1+UgO\OI5W5R3TR
HHV<[gbB_]^Q(G69[@Ab:Z9(A.YM&32?b0@<MNS_O54Lab)43Q)<(:T)C)H;Ma7c
gUVK9,Zf_.CX7CcZaA&^92:AJ397GKWg=E>FMUM,;=,+&Gb4K48/UcKTA(TO8_Ka
f3[8/NLKF1FNJc#2S?H-RYdBe=c4Q-f99MO<(@W#1<40VSb@@V2_M1U-H4^@PG]O
+#fOgE)]g=+0UX6VD>]3H#FD5+]LO5cJV1C8RZ:_<=NcLKJ21CQ9>N4&N66W0=9;
10.#2D<O-]^?,]d/Q\4B4QSIBdBKEN2[^#eS_Md;(L2Gd1ENZ<V<0Y^6]KU2(-Xa
TTd)=ND]XSH#PSF)SHMEeJ@.JFRUGY9]LGNGb0KOL#3d]4Y(5E-;.L#8XMBKaRK?
]/K&U)]0SF8XQ/X1L7VS<,/?-5^&BfI-WL]MX0^HfL&OeOLYIB]_SWOXZW9,bg#/
VML?]d6JI7HR_-&=a86KaJ@DF.TCL;F.dZXdb^NU@0?VH3eVd8K.XbZ=.HY3^/?e
17L_0^3G]K>Fb5@)596]RH9PI5c_A31J8AMM,bM7QM5FZF7,>fI4[aZSYaB&[DB.
&Ld&O6M&5(IgYA3O7?[Q40@;_-Y2gTG=LTg8F,SH5YI>?UHQ8EOI6XeNDO.g,WG5
.a]>7O3<S/eSL[CX9BG>RZgJd<J1S^8\P6F@1#O/?>NJO:@gJM-.DJ9-@/9GfBKL
.;\VSE7e6-IA44=2=L&0N7\B>+;K0&\S>Y6:5eG6J+-]KAG1N;R4AK>A@5,M3b5-
;DGGM^eMP(69@:@_UY1>-Z&^L5MOL8#K@9]?gNMJKDMX<6@JCW,D@?6N/6d:4J8B
Ye;ZcZO>Z/DZ4O?8T_A<OX]LPZ@1Z7)^[79[aPaDDbNIMNXDF77_PN^E0e;7/B(T
YQPH,CJ?EQ2A9af4/<Tc4=beMPV:MFK=e=/.#MQ&)1<^I#gDb>?&,WO8(4X<OM#;
:X\DW01Z&V@KI88&.23,E2,?8dQ-T44;;Yf7XV.NLP@\;L1dR?5UHbK5&Z?SCIG^
I?[,O4f.&L_eM8),)(,X(:FHOL.XB1BK#X,RZX?CU1AAS=MgL/b2L(Gf=N<_W0@_
gY<Y&@.;g&]9?)U[V7Y(?M&TX7fYBJIfO-.QfFaROd\P,I&<&fR.2K+O,=fHYT^e
gd&KBKS9U@Nc_8N_G(GX;-?P:=R9Pf^KK6:9M9]JfQ/S#DDd-N.E:@a]<Q@geJa[
M#/W;,A\64cI7RCE8?7JS7HQ1018=:NY=F9N0#/^5M^=)E7KZJPL(9c&RO^R[d:<
\O2K6>_(I_[XdD(-C/PIQHT\V>Y:g>-ZN8WC.-c\\fLDG=LcN[.14YNX39YSf[O^
I@A=O.LDR(?35NBf0[&D_-=/XV2Tc.=3/]F\:ZP]LgQdVGB9=KPb5a:(=I(L,3W2
=]?6&F,DU1#a?b&(Hg7bF(#7^HD18g>]&[DAQF,^7TDFMA6Y=IY-:,HX,-I_QOB9
W/63L9KL&\Ff6A5C3HWF@(E](Q3>^J>1@+6AL5U\VIV]Ub8E4U^L(O]<(T&^VFC4
2T(B9P?<fYA=4BR>/4HJ1EX_7_=,H\AND&=f<GaHYPOOc4AL4OTZCL;[UGR_cYIb
25Tg8H#:Q_@\S^APDK^Ea./)S>;GTV;Hc2_OJfZBBNKgZ2J?W1(\I\3d;VgWVC1@
,\B4;7K]]00@JI?8bZ?U+e(Ja).^&HE:9,A)\^9@0F>LQRfYb]<X/:=4UT?A0ZFC
2R(Pb7/8NLB3d,?)\X.-L=_eW<;eJ-16M5>G^a>\N.Z(g@\>N.JR]D1G+b)WC)^b
Le]AWd(BZ1V1\UDR7-P:X>^5C#T6PLQ;9MM7WgCMdK<D>(6DPgGRSgaXIJ].:[#6
OaO:@&L;N(NOH<648N:)09?<XSbC7J=]I]4QO:8fa:D&)U:6:HSdgVD]I_,3K7/?
EB]UN[W[:[FQUJOI1?SITYe5<dcW_UNV5,H=\U_25S_F@+9\)]GYSZPcYIbT>C8;
\91P6Afd4SL#P_]4Xa>]f]H4;=-,7P+TbFX<&gO-Y#(eaCRK7>Xb,#[H>J,e,(KZ
:;=U<Vfc^H7@O7:P6RKU_I,YU3R#D-K?Pd&T6a]I>QNQ6Z#E^ZW5^@4f?CEL4<W1
Dd4\O^Y(/HQdHOVT7)G\=;1#=<?M2R5Q1/5fHc;fX_f.TQOU--F9(U9(S\(fICM8
A((EQ)^&f8/D]VP5>Y8/gMVVO\V=+0PX=Y2LV1d=YN#T3E+Lc-X1Y8]V&/de/JL]
H,M94V<R,U.G22P6/.D/>H)6S?CS+6K@#db&HU6VHeTaH^-O62)^WK)WQCb0DOT9
Ae5WDPN3aee]&>U6+3Z3-9.R6&#4^YePQMF#)R[_XI<\Y#,Md(..==WAO5.-&?>2
g<2H>1+[ZPaKB@1__WBP5PKRDW73AON0Z]WK+7_B>FF:33ATT8]bPY:?_/NZO#YZ
,C]g_:K56O8CN)]G;Kb<>):Eb/LcHJ4M]3QLX-;T_;dCAO7fLH(FYJ&bTc/&b]X^
6NQK;[;OJZ;Df38L@J;Ye_(Z6PJ>1-dYeN79MOU1NE<H1Pg?9IS/K)[51G\TNLLT
#,U[&V:2(TK(:=H1bdX?^JI#5c[#aHZ.+\T8?TW_7B-I;)bK)^-:6KAVL&W^b6,Z
JL1&a;[DbK:?;SKe)+fTY5GF&AXX7:M1I\KKZZ,I\3/<VJFb]0<^,>X6DN&U@C42
IA-D-U?gWK=ZO+WZ\Y;AW.-G\8X>AR;JM;J]T).-X#:99EJ_PMa0Rd;f.Z(,TEIR
))AX\E^#VYRWYBX/4^JUMaOJ,f@6W7>]P)cVRAQT0H>IY@8TO=dC:W#>Pbg.=N21
-_YgZ#<)ISC;G^1][6,VEDQ1e:>JTN<SZ]8/UDAL:F+CK>M3BQIH5EBRSfSI8I]6
KN.TZA=5F>&BMgG\D.2EU_7JUCab?(MHbE:VDcME#<9_,C\UCH?=bFBY77^M6aM)
&-?IZUH/#V]UOK\2c9LMefM[-M087^^_:bMEKTfO@c[HZS#R0[L/]MEZG./@U^^?
UE.BCZSEXU01GYL(.9?LEUQ9OD,06T\M0G<VHeM8;Bd]>.NU)g5f._f0HZ5B@E^B
9c@&Q#,^/8/2g,VF5<)&(X)<VKX):K4F7MTbE<gW?@<PR#IX2+cHQ>N1C]ec6MV>
ZHII\M[IX6A2cGX&eCa&CKU<Sd+OX^B\&a@5LD4S).L=[832O>IT\+YGd1b#(+?F
;d;MCJ^E8^@1Qf?[NKEfN]&086Q,4OR65WHa2>2Z8EH0I4dZ<<-.=0b+aTQB])GU
(I?0P4>85MWLW_H]@PFe[+IgU_g@XSFb\_943gB9Q5U3O_&ZPgT/Cg_C0]cdTE:b
I9F\-EfcR6X0J7MKbEeP.)/L\QU^X.N-O@I>C=MC4@\QaQ_\N]RN>^Q/cJ23HHH>
-@]Y;RQ/aCZW=P>JI2M\=7c7/G1KJN?8Z1/2RW]XI[OBQf9;0aQc&)Nd1TAaa_S5
F#RG&<^B.SSRXH[UC+-=9-;<+)Z?@TC->S&/O2#/9^,060Dd54YI@I7-@f/V\X(b
>2_I))JgXaR\>13N(J^7>01BTW3+.d\f6X/[<<e](Wd_7<:b#TNg#_0?.;N8<S=X
(He;Z1aaH(X6cfTQ;\Se#5Z>.JDRW49[ZL6NUK7>9O7cJAA3HcgC17X;V370.ggQ
4,E^M7>=&G?1)\Q@DZP<V4SPQFS#X2DcSVb\=E^TXC/8L,d^CQC:F3SOIU3d[e<7
SI@3cFLF7T7aVGJaQ5P5/[9aUF.B:ae9667HQM0MO9d^T]HWfZR:-6,7Yg20(EED
:Dd@@T^eHIKPa=(4#Ca1Sg@gcLdN:f@\Z/,Z+&1MaW)OHa^FFcC<BM(bLSU=M)0,
g<:^JLV[\GKYUF^WX+Ce6dL/V;40ELf2<bQ_1V??M;]ANP\>8Xa:BA=2R&0/<eV/
THP7NaW]5T9=TSVE:RO.+]<(?&>AR:CW0Q+WVR@UDVTAc(/L.Q58,L]O840dL_/,
0e&>f];Ygb^Se[5[2G1f4<0Q5(/#(1?G=>X_SUIU43T)7d0@/J.YS-3Gg3+]#G^g
QfK&(.&&S]4C+O)<VRI:R=6#Rf3,aF@WBZ_?;<7W&@&5&4=3?H;@[MgD8.(c8_[T
?6P[RGLUR1]=S(VM9W/(JH>XQ4.1Z/0Q3\;=f4IQRO5A8>e012PZd=FT6N(,@,ZV
1&1Z&@K@@BP^3J_CB/F/FIT/\MEZYf8X?AdD.f>2.2-D98&9R?+GC5(S@G9UKW/N
^(gV9N[+79B>S1EZ\)d_32@B3Ya7[cK&#I>13Ofd(Y<QV@/_[L,C(M&]#58PGS8U
g<,4^BD3/=e;F7eP_7fg(>5]&D[5a?ES5VDQ)R&>Z5Q+.DWZ?;:eHdI?3-5(:0dD
g<1MWJ:@02ED0MTJ^MJFgMAR_MGG_?MVM5.D(:eT;UP2-YQL^J\WPb.]7fS#2,9I
SJ9C0(@?LA;0DMCJfXM..+bg<06@7W_XR^XY)S-G6Q@[70K(^.4a#fWR._12DU9a
:^6HM#G<ZSW=A)67U#JSGJEPbd=PTVaTdO8-K)[V3bGL[Re;YIE>TS8,ORTgWJ2c
X>dTGWHES_-6BOJT&#/3203&&R8Mc\-cgX&^37fRZ>D90&-@-8.B>?5g,183-/eG
DN)[d-D8_QS0]NQ344WcT@G,>P?J(@0[3:CA4FGdA,)P?:OBe?Ca+N,:ME8N/4(f
??g<@Hc6aZ+(H&[3R&aGFA_Z>[=TH)U=L;VMWeEVD_,HDU2N3IB/-Z;P3-PT5SgP
:^R260\c)5,<M7\AcLeAS[IJX^J0D6AUP=AU@d8-A8LSc?-Vfa8Z6S:>4X>5AM:F
,/5>&YD[?]&MBaGb)P>ZP0V,]^D@5#VA[\4#I2deDJ67?#4\?d)T5P;LZDG#:X#7
DAF(-@8NBET;=0D5_/Nb+L(faF#abX9@..>_5L?A)3(aUUL(aNYB15GAQNMTI81L
MAI(H5-O0#Q8^#=JV0<a@2R-e:-g@29]_</RTf0KO87&I(VU5[8N;gB<QGARGCa[
M@OGUE5CRe@a1_P3>_2@4M?PJGTLD_M?.RYS[6AWPQ.Mc10Wg#DN=dXRQ(bO<Z=F
XfAf+PZGFR9DB6@;9#bOPbAW^3Q/c4L-[.0\VU:[)e/A;Y0R:<SJAHNJbK@8HTP;
?#MbW_=LV6R]NgMLJW4I>R]6I1B[J&e-BaB1##T>X&[X.:A+1J[C5[7F:0Z6/MC4
a<c@g7H-3U,G.-e]VO^#.9ebgKgX:]Ad>S)LZ4GSS3]KMOUA93V:9g4ZCH_g^:G[
eDE9ZH0I[43K?^N/3c[5<I,QY(_#(UbdYGHf2f/HWT\)9Va=]-;2Z\ZO=V((-<8>
8I,,+dHW7LTgS_HQJI6P=8:]-\=TTSX/-910\D_]KL^W7FK;7U6,,SE)CWN.eTf<
aM1G7=V6B@^/;:IN:/[LHF@bYa+da;O6C?+fR\>4(@g1H_Y=[U>)d>Zebb@IVR52
22d9&HC<EQM4B;R,:]P)9391DQ7H-FVU;9-H:0N.VPefIZYA<Z)LUe_eE^;&0SZI
1e.OY&5[]_dF<E;KZ;1D,SeD/Q7M]/,PZ:-O=5.Y_=NM3W840.HW&R85D\4_dZ,&
FIBE=)<A_Uf8c/VbC5;;>#Oe^#,UH<?ZaPO+(J7/<fXAPSXRdS>P\XUeS1a2]EWQ
NJM3e2@-d),7OU)9X+EQ@?0J)T[3C-1X8>.ddTc>@eVcK@SdD18.-6IfF-3;5J2U
R.@^WQKf#Jg=g^0=OE/?T#E^8Y>3e37E6Ie=N1fD:3V-=VG9HQ#)QY+cP?MKW>@O
K5)G:-YFOOLM&--bNLFa)8IO_2\PT:Sbc91+RTG+=_G-29094M.TEffL+/QOg<C-
++565/:]]SFU2AL2Z3?aROB8U;SV-Id[8[G]M(Q;Q7A&G,)caCaGg)J+de#P^\LS
@bC:C@#bEF?+_#3&95M.1W,V=,J&@d<^G=[BC)K>S[Y;KJQL5M#PK^f.3aF&6.)M
)O+9E6^0IegI+CZg=PYT=\OU.7F=1f.Z&SNa563N+e]?RVUUUA2W\E6,S,29Yc&0
Z]^=-;\-EK>:,@)2,P=>W\,+/5Y,42L(9/.[RW1@N(Ic#1<fE567gBU7aKYR6e:V
<1UID&7=<00+G1KM;Q]37^I.PE@AE<YBNLKU&^.1UOZ3B@:59K3/MOK,X:=J.E_)
:e2_D:;A[_V(a/D<-A3];6)eXe4Y8S^2O(/F\RQc#=X?cVg4B/W(ggG8_>P55B:@
@C]WU92@7,Bb\EcEF1FIKWXb^R.DZ81Q&6YQI-8Y&6/<8J-=SIbM<W?)(WgJ-/d?
_#6AS+L50[/8a.AUP)6=SPC>Z/H/g8)J9O@YGM.K-9=Nb_fLFNRUB)eDcSR-Q0@U
[GFT1Cb(,9EN+9e./Qg_I:F3Ja+We_?[>8YcEM5?=K6cIEBdX@>fQ]fP]fLYEAZ1
,,?)fRd#U(?L-\[WI4QA##YYb<OK9cV0ICJbI@GQ=]#OAN(T\\0:J<^db1<P\_M)
OCNO155_<CZg2ZJ.YDRS:W@-)Q);8e@eBHF18Y3:AI&60CH\VBU@^L@>@K2;VGb?
Z:@5^>@QJ,1-.CG\XD#GT&F^\Vc#:G9GB=9gKbYRc(M3eW18,<5^dJ9@9F_RF(;\
-^]A\U9E/_b?^MIZZC_bcgPQSM/ETZUJE_9[YEc]N0M/-G;TX0;@b^-KYDbY53AL
=;J;SUG4KXV[VX;=1=bdZd5(P/Q#FOPSU:Kg\EJ4?O(e4W4R&DX_4\+9R=\-B6Q0
_^^X(1F^/DfDBb<TC]RaTRf<57V&#)()LA7b>/Q[--b@.TD.2aYYG93YT2F?J,Af
@M>OfR@G.L,/_YJZ=-g:W+,S@4]^4#K6.L7ED>#_7^A9\>TNX633;XZJGFTU/_BU
-<W@A(:?.Ac)-g77N^--4CJQ.JggFJe#ODEM\9cEMA[cV8I?QS\@fH/0Z3f\dANQ
^D90TO+?0OUY&U6b^+b-RY&5>E47NC;>RNZQ0Z;4;JC+@NN,MRXKR45<2S\T8C62
UNF8LeBYLH36#GegV@-(#_4]<FdUUMW#(WFBX^W-bd\0J03+E;,;Q0KVe)AG2aP8
\8[^L(X#8B&KX>)\YLBIARcVOK/f,[Fe#,PYZSLg&\3gP0gP^OTFDVQ:C^)f#5#R
@,?3(bYP,W.g-M(5(Nge/ZWb16TNMG@4+4YY+7F/E5Z]ZdUK8SbK?B9A736:50?c
K4-Nb<eg[5=+DY?Rc3(32Cb?SX-OfT)ZXDRXeSP[/b,b/OeIY:VE?1[JC6X[3[-&
[IY5ASAJ0+64]7bF89&B.30GBZ29g:ffeaG6JfCK0<XUO3^UcaF0U]8DbQ]5d/b=
X6g[:a<MTI2Q&fX,I(WDgL-S[=AO]XK^VCL,FH.UM:D9=+c].f>b^:MJ(]73/4cc
MZRMSZ&GDc01F0I0<5aU)9[V,fQJ+@&X=J0YF.YX<U#1.<B9A+E_a8=CgXb^7e2+
E3J@0f8K:-KeMMA,[^?94<c6-c4)Q&@#OdX44e]._&#XMBT),^37TXc\9JMJ]b<6
&&^CRd=#PU,0(3M6K&V@e?SI6/fL=VBTN:918cR<7IDegY-gQ^[6DFTZB,DDD7V_
T[S,)O5HE(dJ2PYF;\?4dd4d53b7cZfB;B28YD,4(6VQPG-2@-68cc[M4]Bd^NH^
^fZ=L;&VQ2abC(<8T:;NLb\2TAegU9L=_PB)XGH2(#gM),&Y&.DAE]+-T7e;1Be9
96QY,PU?/Yddd&dNgTYgf)d=PRCeeCTNgUBV@N+5+[e/Y(QYFC;UBM,Ka=]/X35H
K.JQSW[eR<adJG1,^f8(?_XMNX>;T^W[R.+JE_IK(2a+&I[T2AO958Z#-&e_c&_)
_e[X98aLVN(_U=Y83M[>JL_QG3I>0N4(E7K>4<@(DG+SNSM44Md6SX&HPZ3V,A4O
QJ+3Q]f<;b:cL11U1[P_QKgXIF1@&]B#J,M<AM@7L12Ke;=FE0FB:XMeA[O9,BSJ
JHJ<J#9Gd>=&/J+9-8(.ObfW-+cYC#VG8,VLc4^VC09^BbPcEgdO6[e]IWTe,=+Z
beHZ>5\)6]+]c0O:\578KAbMfHU\IM8-)(<QDXa@.5NY:\@B\WSB/B:#F+Ya&gF\
W<LJSUJc:L9@3UH;6.242LJc/V&X,NT+C>eQ/[LLEIEb45Q<F:R:S-N]+:(HHH/9
/G:d^=RBLQc/ZW=Q&-3<&)KW2T1f<Z?DW;2Dg<5cWIM>SV7W]@e2g(c;S6bgBG1V
)?Z)CLJTFfWM<d@Yb[L:.5](KCd@J@/d7NE:4MQGH1ZdW8S9_:Nf#5gEWD:VHXF[
1_aPaY-/I./7=795C:0W[9H1PC)OEfICbC<LL:8-Q?P/RYU(XRMEA0&@UC_LR-DR
,VJ,@Se_,dORXgdR)7?QMB&TKCZZ,R\(_feHK;O0e0J]O5.LV3&J8NJd6.PV1EJ+
[dK_(A=(Yd7HPLT</>EKV9@ZJc?<4:^X.LF8W_D,P8e)-QM?Z;6c^^eIM33X6-@N
-c4Z9](.)&2)12<4EYfZe-[K;Z0/=cTKY^aH_8f/e;d\3A,2QIL\eMWaDE:[&77#
=.E[8#N^)Df2Sb;)LGSe7HKD,YaOTH7aO.&T.cTV5dbOL#f5Pb,-b):c3cb+LVWH
)R2I[_321bED1.8Y07BN=NF8)\fP=c2YE4GMZZQN;N)5G=8@(CT[97e+Y07P.>>#
88;?eJAR&OU2A^<UWC._Nb8])?3^Tg0H_VI912NB?g03T37M7RQ2#;8X@G@)g4c:
OA)2Q)R2^W]4\U]OV6cBQ=<CIU;f@BNN)[HdD1VQAd;dWJ,g=4ObN:9d\J(.44P=
N1Y,Q[K.bP+I:J<@E,E_H,3_XIS0#L/+4QJ.YLXSb5S0NY6^81<,X,V)FQ+-&J-d
FC:BL)C4F?_bKM243EYVJ9F?,9=B6G3O9&/Q;1(3A-D@LK:V4d6R4M7E+(\&5<\(
[_dO&KJW<)L2^0=FRAd_M]=]XPU-M,d2O4G5gN,6bV>NFCI&5I)N=&FJXOB&\5]U
6F2OW+?DQLD#)T#1-_aCJ;g=8^@ZG[^c-YXU2;V:IF/LYM>@;6F;?+J\/dJ7\U+N
[70:IT<gLN5NVe_D:)ODYSU_9/7g@/:IA+>DeBcQ[T[56#3.4]Za77&8_XZdbH-=
<UVB;DKf;.DTFJ?b8DFEPAX5-]fbO&_OSJ9Oe8e(2K2,We9.>MK(YY4@1&CZdL3H
eT#T:Na&:b#(#?,OKc^&PA-fGUeV.[/D<RN?&D9gaSN<7AV4b][PXW<G#0Z0:4Y\
CCW1aXO^<+LX8S@=49d8d]e]OTN99(L++?[7+\C)1_]_^7C,E(#I5Y:E=FE,2Q&C
9WQ4CWODa[=5ED(0c_N-O_B0/_02?Z3;U<R\=G6QISAWE[EJ?fa=P1?\#:?HX@-)
QP]F]#Q&Af5bVgIbfceG>LUO13T>:7IF:_+Sg6+&=OH\DC52[891--Tc/aNT(<eA
NED1FcKFMIe;<3C^0YR)7FUR#C(1a^@;Y)9D/0AVSe<EH06ZN33Ge1;c-b6e2X@&
/.D//<G225e@aZX,VbPE1<Rg7MZTX9g\K?Ia]c2Eab86O3,JE@,VF_P)^(:,;7[V
TFA04BHH2@a7D(SAc[AGK87#.21fF@Z(6P#Y;R?-[TgfT<KcB<2E_J(P57Re#\.8
UG1S)eCT#,X65+2+g]:JW<AN@WD&VMW\Z<DDcZE[_33dC\Ma5.>QQL3\;^U:4DJ<
V]9CdLQTW6ZZKA1NA]DE^372ZY#-G-E<U32Q12JOf[V0>[<a-dJd9dS_:(C>)=d@
Q3H29WHE).#=F4WCDJ8Gcf>:19]QLLe-86.J4<[IM]2<LP+?b8McQKN]Z@[FI-c7
0;+63ZIP#JCNV(4dH^0X\YYS;g0VU#L_@4+fF?Z#7[B2UWR.AYd=@QMJ3Pd<7FZX
;;A9Y#TM,>FY@g9D7b=J0-2cA;gF:g4PEUWK78/XE;KKPSCF&(JEaL6]d9A<GY>R
dMgOI(;.2I53CKg3@-8&<JE6gQQ45C_eNWdYM:;@()K.1=Le]ZL+T4c0=@MZ#R&E
aVe2g3#CQN?I.JdHTF&_)5BSX:-:<HPYHAY]]?\I[U1A>f=_c.]W4=6(D)fP/37H
L#=#:]@7D8CL@bWTH^=NSKK?C-@;9XFQWQ6MQe:>SAA2ac]:\_L,92ED_+e;5;G@
,D,XfI=:1XPPTCOb2bBYbNfW&b=YJMJJbFMN/C1MNAP8NY4@JTS)J7Ue]R8@OCCV
g1G_6b4E;3DGNEZDGOg:JF;.]@+\(R2d2LN0K.fEFH6(1<-2WI^.Z:bI44^\4?:)
T1J5/+FJU_G[?aDM3W]9&U(1YX)=1-CHFW-JSK^V;c&-e3dAUT>^N.[@E/@,f7_a
FeXU=6Z?6/fedU=US+VFN[Cd\X&<I-FE>fe#YMT5]OB:P\1E>,-_X+(BbAa@XJA^
H<&L]N^eK./&<Y-).f_JXTX?PFT#WL/PF1Z)A2.TNd7gOJX0]#S@P@WE?\3@bU/1
5E/.O:=-7FQ_<:cN>_XK>J2J,1UAEfe[QAc^+<4Ma;=>Z+C6gM\IZ-3HB0=Qb#W=
\bWM-W\=W-^CM&FZeb@:g;5f8b/c-GR@4CB_V0)b>Z(cAF<RA0PSJW)4F\T1M<&X
#dHK^9-dVF2]):V>U=6^)=V,VYg]8DIg1ZAYeAJ@1@0bdKFD/?=ZQBKI:W.RBYU:
Td)Mb;gN]F,CBgBNU^-:(B9dGA:P+R-#3R35?7&#FA2HA[G\#b]A-@KM9G8Zf&B1
eeAF\H;8:b4@_YW1XE54b(X@9=eb2&EZd<^YgB@>OS1XG?cO1\Y@-7AM020G,6HT
(\e]BG&0aOTG\V=IAe4g:[J_T?[a:8EeMAeFRVeERScW>5V;._#<#LKaSf?W]T\=
8H,+.SMPJRb_4RP6bbLS_R@_C[:2N_#XP_OJ2;20-^+c;6d6SHAV65a<I_#1b,DM
NeZ0E1@,eRL0[Q+1Of:V&<4YdH^MZ0M1Y0fDU_==\VUf9P6eLL/;EHP8fC?<@D6?
4&5IJ1C?7ORBdR](=dJ^Xefa6Vg]XAc.eER6f6ZVUP_F9#7REDdR]GD;IXPVGY8L
a)@W-408f;^-].:D4Pb?EQ3R^QGHT#aX&-R7_^7)D&?0Tb+>^#&_Id:5Q:REV+Af
caR2S?bC1[F(2@8bYH&8M1]fD;[&2b,(<WXL]QDMe0GfJ6S#>I[e+\[#Eb16.X]B
=?TZbK[OP^#2B_d5_7(SDUNKBO3FMc[+&g/F6S,gf>UB-:ERV&OA;6RZeNI.O<gT
2Rf:KNZ5gRPMO]REDC_D1+#4U9a8?>V2R_4,0NBJ-S0YIF?PF,LfV6R_KEU^@#WY
b<+\W_25=<N\cM,eXL7MUAN5N[DVM#23>fLVaV>>g,W[H56<=3W3Ha&Mb#\96CF>
P5Re5W/<Y8/Vf=e:/S=Z1Z3)1JAfLK,J^XW72]K@;_;J7K-4Me#.MG.83A)>@EcT
@H_?.2[;2AgWH:AY2[[[9PM0_EA7^?a>/W<&2=/;S)Q2PHPf?+A0KSN:cS^KCNdS
gFK0a]>b3]:E.CZ#6Xa\3X=LL6Oa#X?]6dHIb2NG<6V6,YA#6HfSU1dWI[VU9V,#
U0X]?C0cLS^(g:Qc]GL.S1^;K]DOTY54bR)JP;R#>W@KW+Jgd4RMXXE@-U]2WS\1
,g2?KVR]E<NQ&A8b5.T(HQUP6<J6I@;Z;;)C-6+PDea)MbO#VI^VaM2<\g;0+7WA
=Va&&>=284)Q?c:7?M\[32WDQ9J[Xb705)3&4aB/fREM#ZFc<6DQKbGX>g]49g@/
AV;Bae,6P&cT0Mc29NFe7;J19+Q])FfMLZeN+HZ9<2<V#O+\^=b\E3,49AbFD.Q_
3GWd=c#LXA\E?TJ9J;Zc^.^)eU\g_XITX]AeUa0I,R@CRde[D:cPd0O/a+e8C:_0
eIM5TYW@S()M@U7dF#&NG0^M/eF;dMgRca4]NW7^D^?GG\GW\HE1:0DLR7N]7=#F
HX-R5Yd,,-Y^,Z_>e8Gb,V6c9,Y-GGA1cRU(,B#Rb0RH2B&X/R/QK-dI>I:DPf\L
RL9XP^NIL8A)GX),5?AM;5SFCZ?gOVa:A/E3S-8^>?ZN+eNc-^WI(UG(;IY4H[0A
<W@GD-gXL3Ta><>E5DdOSUACPD2dF>(QR?9G_I&^(We<7NX;+(C3CcA=\3Me?P;Z
(+^[>M0:fPc]W&,(ZU+XA<f09G\MB6#5>b-P#BUP5S-#AfCA8ZMCAg^KbZ8,aTC2
1^AV@,VF?e[,TTHb\#FP+a)3YET>bZ<7+NL>B(W0bDfWN8<_)9P(E\-Meg[7<ceB
?Kb2\gDXF(cL@R4D#4^E14ILFEd+6^d;I^N>K(fCSJ6\#a8e#cC_fK@K[b260+I9
SDWICZ>1Z@:<AQ\O-RQ^4?#T>1?W8^a-Af:^4(G];NTM=BSg#I?69:/QB+M9BeIA
FX-Oa+R91Z[,A=:JFS#H(FG4^AVV])2E.,^,-VeF7<@V7GcMBA2cDY5N/KN0[NF>
P,MIYKTB6ePQ[<+2;-)g^L:-KX-_fXDfZ)ZB738/L_M0KH0,cB#CV=,7=,61aJ#L
SR1&DTZ4]ARRf9eZ)8EObL::5?///d;H^B5W5S;40EKEf0fOOO8?<?NaW6_KFH(Q
I?f^EQS]4H=JL&)3gQV:Z55-;;8@55HGd]KLbbZ0fM?XUfA.KaI=]Q#H60U9.>OT
FF/@.Tb\I[M_4?g+D;GK.H&5_9=AE-L^ba&\f+P>7=:,&YFUaaM?26TcE,8ddT#Z
@E2d[;6X4V+A8LGCcOAaL.E#GZd]]8KL822T_e=Y2?c=/K8-C1P<];2EY=0G48@9
\AdQ74]g@1Y)F5F-(KXKC>:6H/)B0.6O2fa+\1MH5AHC6[>:5HeBJ[FN22E[[5b8
EIJYg1;aX@0HgHQ3\[;EM\ca4ZX:Y:/L.6/+)/CQR[NF]F4=2--aU_d4G_C1d6,H
1I/W]ORWd0?.&YQ]NI[033N-[9aH/@,5:H_e.@_7>a#JA8#@/L163cM[>=.@e73D
?8_gJc(Bg(V4M2:>:JK\TfNH.a0-X4Fe5K@Z+T&D-LagVYX#5E?Eg0+8)g4@GC6<
M21XXe/QOA+fDCQ/XNRXQ7KDA)H/I4cUBJ_#PDLS<2dPfJS7fT]LD2LaUGN+N?W\
EfX>Mf-]2UD\9cS<.c)A(VWZ46=fb907Yf+:e?LX<9YJ)Ib[bBd<4HNHXU-OaLNU
a])25fH4E,=9/7g&W6;f63:=W&7VI(R=U4-@42DJ>_/RKW]6Q7S[_56#6;a&H0N^
gdV7_fXdJ1^UE]5Z-\f&K?@-PaU,[LOL(V,&<,0,ZYf#1f(^A)A,DT.(FO.,]K;?
#<]XN/K<2J8>:-1fG(]GXJObD2C1C5BMT49/,M^fFLX1R4](\E+3.YO>:4fP,_de
(WN.#>X3[_\L)86_70.]E_gG^/-DR8FaE20R14EMY39MbV6^SJ\]1#=bDB@Qd2)I
Yb+(7(KQ7+-Kf(R55C)0.027)4>YM(@1Ce/?@g<IJK=,D#H)XKQH,<&EGf3<9(JY
4.g9O+AbNKYgbbZUY=TbcH)Ua)ccKecE8fcW[(1dTJ0S///c>5O-Z3Z5aK&I9]T8
:Y:_P@Z6cOPX4KEab:b75=&>\Gf7)8bV5fJ.M;C3JN;,#<:4gJVA@&3/GW^2V3Ka
13Db[_IN(QOcUG:EbULdOJ1.;I?D3V\WPT06UDe?].LGeO1O7a.YGY3c.1bI7]L8
\THF5(>T_F:(W+E2J]XMUBfaX\gQ@N:fE53Dd<3H=G/E4c\D<3f#>J-/:<baYQI(
OLN:5b)URF_&1P4=BcC69SJ7X122bC]T8aJ2.c@aW-0BT^cT[(:N=LG)[NU20E^H
\_HOM)G+G7UbSS#LNCDA1<U4Q_UVFM;(5@,)2:V(VA4.0&6YXWJX\:[fQ)-)K+ZL
MeNcJ1#.-H42Y7T5K8R5FF268WQ=.DY)U1G()\WYD>N2Xg-8f+9e9SK2CJ&<<9WY
BD+NWNM6]L5Pc[U:00Qa-T4T3c#H/&Y?4fU012M&P\X.BA[VfZ-F4,5c[),4WTb&
D5dHT.KS3C,f1D93312c79;]IKK;cES6A61XK,_1KDC,A.+)d.,>\Q=5Pf6#L(eH
,Kf=f);5<g)>aC?H(Re0)17?+>HcD;.;Vg106G&HefeUfQ(?J-1&MG#SGN3R&U4I
PCO8PIZf8PYcE=a)=I,7fMAcKWLTFP0?O#cH?UJ6M4dFA,#2R7eBd=SQ-@[V(=WP
^2+IFIVKE)5e:/FUJ,L(Ge\G9NZO>E(c4#=IQO]V(UC&WRfT/9/5\RBb:,cZ:d]E
-KC.\N?^@<KR,MTJRaNIQ^+5bH#;]X+=a<WTGbV25eVK7f\W5AEWWc]8@YZ<5^32
X8N>)E91c-4-#<D\#UgH6?S6Y3(R2>,@A.ScMFEXZeRT\J9O\1F_?KO3#\^2Ua2I
1YE(a-IB8gJD&0]^V4VbV,b>>G[5?.8,B];RF.>TI.,H]KCX#Qf?Od?4ZTaQN\]V
-DKCB29JBeBAcIMbDe,;W3,&VIT(]_Ud^#/)54-/<D2J.@+K<5e,g]DC(3A=3>87
U[AHc4@S2.=.LPQFD0P?#3WX-XXe8gJ&JaW=W?eBTM&,bC3O[[KN<M@<,<8;.+42
&C;:&NUeE00,R3X#N]9e7LPB8&>4UVH>:fD<T)53=,^E+P[LWg7Ub45V;QSXUW56
9)>^JdA351ZMb&8\],]@]T@/>OIKf.0K4JR>V.&Z(Z&Xa)#15B6,Wg,X,9>(Odg_
<)&J.f3<R^JFUE_D@KJ)#O;Z7UNdBS2<XZbQ:CfDXG;0MB9e/_@BcgDX-gPXKA,_
<+W+H101cePVCIcE47/-J-&[TGIRgcM-D,F&BHY=/^c<D=<\P2MTZ]#NK0][JH><
V1Q(@YAR^T?:73XJJ#N;4@[Q&?3X=Z30)-0O4<S[[1\CdW\5:-J:#R.e_(dRS^93
\&AJ;6_->_+f>5)Z&NM\].VKQ0E+4:;F(?g[eV@XHQBJ&g:+@R2FSLMEINRAC,N1
ZYR8?Id^g))C4-X/&#gEgWKRM?&4L=;IeeB=]de<OJX]BES0(,OdW5K4(.fX\=He
[XX;#VRg;EQT<VGEKKK5N)\1@eSIZPBDV@?_Qb\@Q9K+gKKd;bdL>cJMGH#S^c86
A/[F4&7W+DAX-d\D<:&+4EQc,dXeG&^1+-AH0Ef3MKCB-?4]JQI]T(E?H5bMMR.C
0];PF4JGbD>_J@,D,GS&E8>R=3@7Ta/:NWYLM_7.g.-X1[5UHW,eE[6,d:3ed8HP
SLNCPaJe/4)G6\&fSKXS6gJXBG#B_)W3,GaQNB<WU31?(;,B)?CL:GEV.XDPVA<\
97L1dV[gPZGb4_E&Tea=&cF0MgEXDgEEMW2a\#9P9c.KR^FbG@JF/3=T5Z+:_/NC
Cf>Peb[cM>0^HEYOB@)A3]#&?:@=HSVZ#4M>)a8.eJ:I<GH<-)QYTA=Yg=.(-8)8
EU0g8V;_V038McE=]J;ZAgPBU5\:aeFG?fGWY47=[#YE_bVOWeI+:0T#/E6DbU7S
:IHJ&E1YWX0OF+#E:(dK741ZKXSD#=90@S<34[H48O+2<R@eRRA@L23Vc[fS0#PU
N/,=W5Gd.6NN<-WZZ^M)f8_CaJ+BT>EKN0,_@,&_Q/8&?NT?X_J,O8W0BDTT+>AR
2/Nd]XOAcTGaG=JG+4)UeGPT8gLC3OJ39KfBg]J3(bZfG<Z:OJHF3_E1HP=+C41/
)JVf9<XLD/F+3C;3AEd8e/Z5?XDPH?Z0L9:cC)g[,R>E+_d0SV2.L9M/UK,5gd;7
D]G?.e:EU,2VJZe/<O)7R#D;43G9b5b)d4\2FZ4(-O[E=R6dHYII(b7,R(DS5W^H
68FEHcKJS_GBP:SHK9eA>JO?,_6L3]XdgP-<Z/\6GF2JK,QQ-d#4d^6+T#,JWVEY
)>B@@QL^Z[R:G4O\9]Ne;:F/G0(>&;YIX(3[#F)W6X/.eFB<e/J1OE?LLR=b=:I[
ALGbPdd2V[[(dWVI.#4J#=^B]<)d#RC3cH0,8A2>dL&.LA\\,(egK[I&L(27(6(>
C<10-IE2OgGS98C[WH8a04Dfc18QY/UZ(gA]LbdJ=Z\2-XgGfV^\3C\^#,=2cI)2
UU4ZGb[HOXGESR,MIc_[Y44We+81_>Z>IWSJ<5WTQ/8RJ\;b6fPJ]g-7&?Cdb8C1
/d[MbRJV8(gC#bF2Z;FTe)SJ:N+Z2WV]-9DF5/]=3-eVGB<K<Vb4+4CJ5fFaMU+T
^+57OAP+0]CgBGKEXIdD:W-H0JF.<f;;A-<(^:d&)+8Q#(4eAHP9NWS#^GKPS6U[
#48^MN2fH-AP6KaSZQX+;P)C;?JO/^Z\I2MGYc5-YBF&_MU)-JB-fBI<&2dNcOC;
1O<C7PTV;JP9,6Qg&cXd)-XLf-E;A^.S\B9aB0L0NI)AY[<F\\O-^OGJO.<fc0WG
R<eUBE:2K,.c.F(LV]T8BRQSE4YWYGDD@9\F#]bW735FbUg54^^NMR>:6QG(#KY7
PU@^#M7_=Qg,65/4PM70-(BPKUHV=,T.F84FC,9L_EP=_/@Gd;@IUFc\C/I<GAP(
XY4)-Q@766:aGXSM&6@AeZ[b6FS;;>(a69dZ-B,B2UF7#72)a9@H@#\L&N^V.C1d
QCE8NHAZJIWAO0LVDX4ME&7S?F)#EB]3T(Y+bL3MfX&B-1:g07>QJ>I,GXH\2;E)
WL]Jf5(f4T4UL#<38Z#H1+A:A6fPV+9BUD<=GcO>.6T)Y6@<NR(_)76JP9XIQgd8
@4H05I\cA9W07(1UWI_Y6[c)JG;2KZ0/9(4ae.<N&@)?_999?\e?YB3&9#ESN?V1
dC?J4(^B?A;K,(7K1,AP?8:3)KE_V)>-V9?c]PWL94#Y@<@CC(@ZZM00d-&K@++d
19,CIE#@0D1TORO<90I_/\,(33U0XRc<>Ub[+T=,QcCDaSaJ5[Y3M@(<2A1O#_fa
Ac0;AYY=aIM5MOI0N703]aS0_Y2MKeB8P@T#cE79Mc).,)H2g]L3+YS6[\#@>4bH
.-cYG=Q6c)T8=cVe_X9J,Y5Fb^-#&J1&XSaX>9fF(A<c\_1PD?@==_M>7-Q^>;]6
8CD\LHfBPQ@?;B0Vf925Y@/gc?67Z-LW:TY86@e-,,NR>PX)Q7UTX7LC5c&/(#P=
a0?]gLMW,LOTW[^G=KaHg[,W.)3)IVOY4FRFO#B&(0]P#1U&CIe<LM(CGeY,?/,#
:NfA;BZM#>M)&B?9ZO((-b=)9Z.<aQFU,418LOX[?T1gZXEK[-&U@D+9EeZX+-@-
^<(O+&9B\9PUYf3ad?G#f3b(.1)<0\NfX-b8^;L/SY05f;5GLKe_7OUN<3eg/ATg
^cM_[AgABPbC9KdGcbB-J?9XT4XJ\\P]U8?DH-bJC.G;2H6Ff8HG&[2@19bL6:EZ
7=DW8>3N.N97NN(<TbM;d(^]6/>9S2)ERg)1]@B#eMRb=Fd#eIB8JJQZ@KL6WZ;B
XA:gcXfM<.VJZ=K))5O,<]#WK#BM&D.&/F@O3JX..;B2Q<_JSfXMFUOfZV-K#cJ]
@<=7PODW9T/VS+?\7T&fc-W-O)WbPfZ2c3DHS9Ne20^<9-48,Q/0.bFT?+fd84G3
O<R3FM2K\_7deTO]He8/]ZDYKReLST.H60AXG=,eR(?L[4F;;3UCIe[<?G&@b=3e
C]1;9\L>T2W2A0=^)DLbS11dP=HWA2CdP7_,E&5E1\WF\=NJ@F[Y?Z>#7a;9)_a4
W,G-D><@_a:E_NF<U)P_^dF^7LT@0^M\#-@64E5dSTZ-R8>dZR6\a1;+&A^G=QAD
PKSS+A#E@.JJT7C4G_3KL)Gc><SJfLZX(5NTWfOCFc5IdY@9_9cB<:dQF=4Z.cEI
JV3b+R+I5#8\NZIbVBGg.;44#4[dJD6ZI[NK6C\G7a&H0_G-N&O1e7CF-ScIU?6M
2V.D2Z;6?>@6Rc@[c4&.0O66XCP2@FU95e8^ZXSG4VD5\9WKf@a;aO[90[:>-\>P
gFMAUc<>7[Ic#5K(4)NXdCXU/NC]-Q4+ESSG6VV5W-D-SF57_4g==/\:S&CbY,X=
2PaX?=;84dUH\^RB-)L>@-g\OK<N2ZDSg2e?6V3Y+cU/;QM>YL01Bc/YY+=,b2RD
8d8D\\]&2O8F1Bb4?&Ve:=U[]?#2:>TcRJ\cDe3@L24^dFF>bK9<X@P6CeRD;/H5
O#=WQ8Q?gg:7eRa@NA>_M/1Z6_bH;ZG(5-VL_A22g5?H9[0WN,0a\C_FH6P+7T^]
QP,LTHb_^PY7SagRe?K+gX1f_g,TZ^N[)U7O^a+a9e].:V7\1.e2JL](>@^eB9c<
SM-AM1#E.\75D-_/W@(R6cA<Z;Ke;QIKA.;ZDVY\4=GD7?QGeG_87e/.YM^&@G-/
1@^_RRF1:W]).YX613SE138[U)#g1a@HQdA1Xf+A>BT.4cHTQ5(RZ((]bI##D/R3
^AXVA>-@SH/C4ZW.GSJD@@YV2N10N=\D\&VGDHa,QbD/gaKfcdEU5_dgW^Ke&TM.
@?X_/583X.)O][C@cW2V#72UI8M7McPXg\H,FXU8V0(:SH5U&7G6.6U(OM>C<[LW
=YBb=,6?>PQC=M7(/ECJ(?Y8bBg_?YE4^ZP>_\/HV13?P&e/]6[3@_7G.97(a/(:
\O:J<I1.4J&(\8[GOADK&5=1X4&;XV;^V]H&)6<JV89^cU=dcBNMcAYPeeNJ6GVB
]VN<L]M\MHH[1U&IV135\-d4<UHKMT=(7,^J3[4a4\;12Vf#]Y;:]FL_05d1^L6(
LQ+R==K_;Cc>STJH@5YQ4:9A068JOSO@K\WV5(H7V@DD-/21bIc.K?H@6)?T86--
cb(Q>_M]L\OHF,8</c>YJ]3WD4a^J#=O1P[X;)P^gBD<#,2PJ#fC6@;@#eg4UV.F
?fYCWWK.KXCfFW56>-d5T,,,N7R,EH:g?EM<LTV,<IJ27)YA/)Y57Z_d<U9L;d21
f\b^5Q=?Acf^>IG+H?FbK+82g+/W2@24EVN_</OHg32YB&aY)O[fJG^XB(Df<G=B
OEfdLL#]/P.4;WP9U-&_/-@R\P[9eG2>XO&V+;N^Kd/aE/D1,LQ=?V,L;NX_@Z7Z
O.BRFGbPLg@AI:]&C?N0.XOLAa]DeMRag-<U6\bNMf:gK8FVF]CHKLZ85SS_)IAH
U,ba_Z,D5DgGEJ]aCaafZ7D=\_#_Y..#<dOTV(.eYJ4090/9HE:4Pa/O6&1>_3=7
P8>Ma@],JT@,]@-H,^E](e5d\M_#O1LBE983@bC[D>#.e@.T<gWPNcC()IS;U4<0
TG,E@Z9BBS#@;Kb60?)4H+?D5.g]N&XM0,&ZUN0(Oed#-ca&0O5/U.&KF543E>XI
#\,Cd5V&(]a\<JJ]FI.ZJ=,VfU@1<)#.9A\/&Z6UAXgSODG5dJ<ZX<GC.RZD-_[N
\/8=+gT,9\&4e<VXBQCPR\F[b]bNS?9,ND_WfBb-^-JQK_1F.UHL/KMI#Ea)P9LW
3^@PEH9_c=V\I[&#.7JXK345>&CXDU\8F6:2>/c&(-@UCgUU#:c;Y:L-93<;/M,[
I=EA3PXMC@E(JI:MIB\\5YFTC:-c8F:[dYTHc\Gc)[2Z:<NF;P_Y^KZ=Z10@MagO
e5)BGQ_S^R;8U7VPCdEHB5&dY)9bNUZAS6)<ZC6NW3;U#&&^P-M2YQZ50[+W-_[-
fb1A+JDV-=dc0_X+2:1)1\>NO3)EB8dZ&<#1KVa5EMM-3P?3T[T^f_EVUA=,]XTb
6fEP;&Ded)]G6b:](gP]VES[;80S?bPP/9-Wc+0A]H;T+5[XGT_B;\ac.O3#]DTV
K(aMWc#a9EW1CZ3R-Ue4U^_457F+JGF6?W]I[ZY@UMX,DD=_)==6EWGL/1VS#.QW
Ia@g].]MHW,ed#^MJ>.K=\MVZ4(@cXIM:R9+e[QDRA;S=[U/fEC_FeY^_/X?DSR#
#aY3D?I;I+0@39\(3-<,D;8V21835R&J]6a?:SeJ5<MO-??6]/O^AI0Q@,+L?O<+
+&KAI(,Xf#TdcI3^;)_?Eb;E7V7:Y+c6d<f:FNL,#W\]cIGKXSfM6_RC(b(a9-.F
ZMI4B5eBZ,018O0JI&Q=NHL^RI\>^YZg5JF/C32EY.BJVK;7e1[XQ53I@;&F89gH
T@#F)8+fI_e2eBL,SJ\F5X92#QWU8fGf5bF?LQ228TOA]0K&ATNefR<TN2cQ?bA2
52=^/gVT1/PX:^4A..K:)>L-b>D51U))JPX1:3>1/ET)]F(bI_\./;D4.5);aKC]
K]/48K>(=(SAP?;SS^X;.QNO&SOa@.>SGY/\.4()8=D.J#JJ,&,0[62\0L[E\L6T
g,c\@QTW1cQ]=O2<],U8:eeF2Ba<2&A?>/F>\-S(OJ/\I6dT^Ld@9aKHT/U0X46/
(X8O97Q<RJ@^#FIL9AgMG73=a#/P8a>.d>T;cdVZK9NGE-94BfORZPODcIL3cL@,
_(F_A5RY^M(P&Z5&5[9IIJU91#g&L@++6#PXEYYXf@QXJCDEIB^D8fCVX]I5cHLR
:/I2H^7NZAY(?-38I(1:gCVTKFUJ:OfQZ0:JE&GQW(X]&EV>ZJg-<3)[MI43V9[_
O\O@M?PgJVTR@NdU;9RPK]:^T-_]_QN3?T3b#SF-5MP/]_@e)5C+cL@P7\J[9;]O
JA:K6_=S3-<B)C]C=RU3Oe7P6+IY>2;gd-BAIX/JfTH>(Z6@V?<6UcWU_\.T=H]B
f+EJc&;:]0JKRO-G[40[@QC:RW>7/\deTSbB_^Q_aVDJUO7(MXKc\?ULQ4BfNPH<
#_fMTK[=gG/O0.FNf9Z/\=+_]HM13+4a=EH=I2G#@547/6/HZ:L(+I=FWFH7&5e_
]FBJ-DP-8a4G7@]A+J]</SJN.0Bf&\AL5OL5L,=GbNC:+O5#UM_0>gX5ZdY9Zb]N
ZCR>2;4&2NJBD(Y?=Y\,<T+K-7EePUCE8C(1=>[W#)>)D2\<b(UdUO\R[;IeO/89
gbG?FYTVEWXG-]d#V;eT-<M9:b5<Ua2=D6b\L6HL=?ac?B)cW\5X/E;ZT/)ED:4E
(@E]&Q6O/U;::(R36C/7X[9eYB[P@L6[SA7(2;<+LbPZR(I?&)IQ;RM=/ZGTagVg
\>XP#0^3fP;SDP-gN@8+Fc]VI7SVN^.aSbL=,]&&^3A_ObZ=\;/WZVcE3SQMM;KH
gM=6GdU#CId=7:_Rf7&@)&C@/^g-eP17G\-5R9@X+:MM2K(8Y,AW6A;VX<B?R)R0
Y2HW.)f\6=,TDcH1^fPT#>Fc8KYJV@H01DE[)fcgP#LLZ5PQ_.b@@f_,8LA?I[+f
c-0LSKf.;NZ=;:D[E9[J3V=>>POACJ>gU(.Z/>a&DN:R9b0\>[CAZbdG5gME=PC)
5_?=@C>CWJ2;4(fO4&ffYOI_0&[:da_2/L7EL@PDO(9fD&0+51f[OEAc:;U;_NJX
,A1d?4d7M&8-[;68U-)]BEJMIF/8AQ7Y_:9ZD9ZA/SQNZKb3F27Ac=Ea-^[e2T/a
,A5D,VTM0=>1VK5JUZcI]+&S=[J/>UO:WgJH_#Y;@Q=L69PM#F6+P9EVg-TL>^c:
;<LLJ+H_gZO2+Q,8.Q@PJPJeI]b67?:91bNL>SLRBT^8,CEYBVCa>ZSRP>V7.AE:
I?3=.E@c:2Ia];0I/O6?2N8B7;OH?.OI<MZcPg5C[6f&;?1.7N(D:]dKe@D_a]9H
,92:.7YNLC2TB@K2V:3509<HH8JHX8C6<25./<<@Y=&_[0:bbG#<4fUQd\O2P:b?
fRKLU2)+5gcGX+LBG(2R/6cbPIKRRX2aT>(UT4=&M0(aaP&=JDc)\T1G/eQ8XUZ0
DSC,KBU40Jd_FN?cQI8NVID=P2/=F:\FI(7BaGI9c1,8004DA2NU(MWQ#8HY=\_T
7Wb;=K\R1/+fE&NP8&<^#K:Fb,0,S;VdW+Eb<.Q&_2N(UPB:Q[^=BNFa_JY>671=
:RID&0Y9H_(B>?c?;=C&Jg2F?>ND_#LOHLGYf,-(CABUJO/=1YMUMD15KAfX+C&#
f-/:Q-GAQG86ca,dF7NU>?(UFb04W.;cTKG=5YR.:TdIWc8/&5\KQY@#)cC^dA)?
9O@?B?3dcHa7K0A8a0+TZE[a4;G9YUJHd/&D[Y.+O=0fG(e6EVZOFBB5)?d^dSbH
^F#ZPNH9-b#R]#\O:D9YV04;CJfTX>UAD8]+L<ERaHWaF=bE8(QF7KF0B>QSaH[=
g[ZL0Z2@/??^G=+2H=?U&<RgE9E()b_:UM<9=07&_[>#-WaO7BA\e^9[eM]B:PHN
0X?/6G0N6bC9QOHA#3XRHK)gWBWGCd+(1./?2D9=:cHOO896WT7McV1TgcN8=M0:
-a,KaD1TG9<#C;QHV#[599.a=>S-=6A/)F,VEcW]I81J\>._9_bSgRg1,GWJ)a:]
e9@SFL<1V3@#I6.1,C0S)\6O<K[04O+HYX2EQf:FK-JO]De-NM,-)2^9D>7KEC&7
LD@LZb+_[e1TTbXOa],K4R6J4J>#,I.AE,e13PZ\&NZN&0SbDT@4G?1c;Q(8b,]G
LCR_4N&\6#>a2X,\fVF@ZCPLD\G^b?2PU(N(?U^6=R.]M_UP:.Xc:D&fRc.GD]2X
-\fVHA2Ja>538#@O/BbN([J_<0?@2HLcV18RD(Oa)ZLgcffgY.+Nf763/FG0:;@D
N>9/ReSfVEa15HK)XaA)6d/<[5PJQ43g&+9Q2Z1/BB]MGJ&,X>R#C9Ae@P[Z+6T2
aUX?.S==&-9Fg3SeB_9ZG1NVE6&?W6O&OB8,QC.270eH4,DD?<S.4IKPJ0/O4DRd
XU1bd7S?E[#5BJ-<[K0ANH_TBAQBKLRO0N7#)=@/HVB^f4.<bJ<_4AX8QJ#5;f0K
1e9159;K4B6WF/8gV0bg]1#S<Ff)CQ6S=5:XQGUNgTGb8X+2ZWQ=^WU5KUMZ-fT.
OP>aaB\I]23;L6/,IL^dafgWK)2&d-Q):?.<A4+WW<2c&IN;LVRJ)#MDMf35\#dT
.0&7IL7WH8YH?J#H[3FSc&+:@)=b20@.Mf9&?@4_,6cV(Z2eIa-ecQgB81A_][4Q
aK19JEcY#V4P>>RR.9+@F;G_;Z>1Q0:Z4D\OeSfY3.B7AUHdA-_gbH^D,3L\Bc:b
e8/FN<d.,:.[L2,O)>]-\<_Ydbb]OG74T.c<3<F_^\=A10;5?XNe.7:)K21]&6[[
@+3a\QU@>B.BW92>B;G-<(QLdaQ11Ze=O@6dbK937\TMXQ,7[F5G2TAF=bDbBFe;
Ke6)D9#2A.&g6KSP<.4@[\K>^VOJS7PN:+-0fSR&@Z0QY:D^KQNM,_,Z9VH_[g2b
?7Icg3TY#>g08#8,Q62&54O5IU,fgZ8R>:BcB7>Nfd]CfILEecP:[PI_DZM_6CX/
bL[Ec6^@JDZ=aGA<F0XE8EX]F@-A[=@T?WW::AY)G,2Ug^[TP@&;LB(I)P\.H<B]
.Hb#GfQIHgA&1[^fH7QY]&+N/R^1TM;#NH&D]E_YMEJV=Z=3YHAR.#&K0L<<1c-L
H=IYFZ3:<T9FJ_L2fPfaJ?)-VZY#Q)dZVH53+]g5Pc?Q>4:7XU48-O=g9/H\f+g0
a(5<b)aB[HX9;3.D8@O96a:Mg=9\>YRTB]BK[+#](+/HJ&Z9fa29?NW;[S0YEg?e
0+BMVYD;O2&.&\W\P&X[^SH(I\5/?-,Md#f).d&d]S=D?I2AN^,.ES<=Z7;c9_9I
5C4224O7V?Y>(]1][gRH)=f;T:EKfF/b^;#>X\2+X&QJD5;A+B&F_#Ie2]W&;H9>
;_/&LNN^/40UAR#IMg?D(F,\W>5aDZB;P2XMDAIS4IC,/QgZMHWC?F?\QW>>?B]D
+c&:GVF9905)7AX9EG^5g9&a3-W>3.F>DI6T0#X>:NM:KcH7?g56AI/B4A#>D_42
:\;Y2WMHId?R+&2A^KSIA6PLJ20WA^><CS?M5)2dOKT\5N9,W?[&+Y.0[:<@=(6A
3UGKA4RB)Z3<HZ7VC.(;K]8@7aLDIS51ALD?FX@]NOKT<:+5R8M0(P3T-RRAUFZ?
O5,7,Bb[GNERV2We1-VJMG,JGFJRb3I1OdYPB)V.?\27FN:aNSC>Yg<f#\]\])L]
We),fM?)5ILO:@V[fVLU,6R>)#B(T:7;WS-[1Z^H7;\V5G?Q=UU9<7)\NUbZI_F_
aBVeMS80-=<FCD5,<Ed0dSFg1HW&&(A6cgEYI.3]OW(;T&]D4Q2>NPJSQ>35aZ^e
(Vg#4G=X-AF947b20,A>0^U<#;OT?S/+=P.@GPQ]T61c=6[IMgaX]BTe8g0dX@?2
>cGW4gE@]e>Tb5BHQL1Y6.?NAS#@H=8g(bfMA=1HD;CK;&=aKJV(=b<ZAU3[YfI=
)<03b5M5Y&::>SST+AMWB=g\7Yc?WJf+B-6_UWY9(U3Y6Te5&XN-E-QdPfA4JY?\
UV5YDHW;[STL71A-3C5c<eecY5B0CXME\(179+5GP>R)KacXG.COW\;&Z;=X8&<S
Q/UJ9N;YBZSGR2:\X48O)0./)2GHY3.Tf[XJEa303bGT;a\E5/HUP#1/BfV>1?V8
K_QS.T96eX]-&SeQTXTXg&-8F<[#55^c;\&0T0.ggD<9EJBNa7YYVRYTPR&YW6RZ
dBeRAS/\&+5<1F5S#KQ/;,1JURYW8JDY3C=.2&;>gTOaA&5-cf3-5E#]6BPU3CP#
Cdfe^dO>32[VKUBW2H/W9,7<IPZM@=D:.>7N_>MV9_+OSUR>)ZWVb4;<b1.2DJEg
3+c]<HEbWKSXP>UT0\e/CLNS(MSfaX\HLHXSBSZ>HF^Ac_5V7b^eM84)P9+^1+^?
JIJ,<^]>C;9@eO+\W>,?6@2\9XCFHNd25PCYT374E+T)fG^NTH9SBMN5ON=M(SZd
Y14FU6IJ3UO/Y:Af\DD9cZ9aWbcMc]UZZVXCB9eE11a\N<9@aeZIS8?FP4ad\96I
EQQ;)IIY@&9HY.9aTX_0WAQM<5N,^=<(]3c[@=N2^)S1#HO=,UHOdDB@160(C5C0
8435T]gP2JFK/ZafRgJMeQ?.Da99R:cNVO>g^^WgJVbR[JP-g@3VeU7-HDF\?GIO
C5]R<S7Y^-M]+MW?H[;<K(Vd+.48F[:FQ?1>\IIT<;[\#8N[)SgJ,Ed3F\fY<R(/
0/RL=BOG&BP(VT[#73&;5[H[X0W?50/YXPQE]2/]KO?[1&UfJ/[?EQ)81^DL065@
Kbb5,IIIK0+7+3-YDJgcY)DYG>-(+3KZ/X@FKFYH<LC^[4#D[8=c)cJ60Zc\2Rd=
fLf^e;eJ9:Aa0aFd-=+MYRI>S^a36T(6FRTg&7A_>dIOL?B<9DO2H7fY(/V\EX_K
(DP:c80f=^LB+=7LDMWUY[^:1T,AKJ;9)3\NQ(+MXKfgF\OU1E.Q82BJbN#W=[O@
_=W<E8[-G=?4<c63MZS9GcY/gJaL@A[_4P&+?Y&[@?34KR;#T/4=E0R4<c\ZaMe0
/,WcY)_?QM9OUY^c&@BF,3@=aD(>+JYUQJ]NWLGY:-[9.U=K=K@e-Y4HR:0EV]:9
,>ADWaS=&RCS/RX>:_DF0_YB)JcDW<IBXF@L.f)<I^ac?/T40Xg54c4XbUGdPXY^
3I4Dcd0RHDJL(gV/7eE<>J1Yc]+0&LUE+)cU2E-9]Z=TCZIAQF=c>)M=;X_aI<_<
K2DWb617ODO-?CYSZ@.BD:/B&cDM<)@T>=8,Z>9DH-LO<[C8X>c8<M&T_,8/@J<M
@3,Te0eT_J.ggc;JM#1:QZ..(]IW3,_)aB#@BJ=R/#W&2b]#B(AFb.(NE:DEROZ.
2\T<f@ZbMRg71WR[2AICBDTVK1U];#WCB6WYKOf4HI70M+1KGDFZMgR^FU>;/&g?
Tc:9@Z.43GZ)f?J#g,QMK-a8>c?3M>7W^7P4M5C=48/Yf#ZL24(LdE0W6-/>A-#>
D3ZX0892RBa1ZWUP.b39O<0EY-W^C/RYMNAZ-<Ogc]#FKVbc#PbdG,CYOT_^_+=C
#@#FBGc/7<B;PUX<K0b35OP8X[E]aee_YOaHZ-Q>-R03KOFUJ:Re;Vf\VZ8YT:R>
E9TI&:e8([PQ^<)@I&,_\e:\V_ZRgA+bUgM,J,#5d.W\;a-Z=+d21-GZ-B\T(&0(
(A^#/Ldc8F6MAf78(7.01NSN-1SN8dN.cKYH@NS#X/ZX.Z7D7^>/B9Z_0:aU^[fC
E+UUIQ.^TCLa^R)66X--+2KHGCCJFOGK3RaZC7MTba?_KX\OUG<,C&0LLJ9&Ec0B
Q9Pfb+GQb=+I54^7N&(OFVN,/f+=.6(3?_P4fBL]P+:O#/#__ER[C21P5BEc8S]P
X#;0ZU,1GZ<=F\=IU#&=ZO]P=^B/Ba\a09[&ZZQ>TK70cMf.@RF?Xd]gaUKWa?c:
S&JOU.&H;-gea61@[]2EaY7/JU[dE3bSSHG/\UOeB7_?.,1fYDZ-82CSbgSM.6P?
L<U&,KZ<I#ZK<9TTTG\T,6U]:G3-\E\#1?:BgXW:f5gW)(2d(&g^^PT3#YQ-FFY2
^=-:R6?dFT&9?b+gL9PCfU@H@b8^S&Q(,_,Q2U6R8]PbV?]-=;7(DI9EP+QBGK7S
#Q)9LA-O1?-KGf8X^HcK2#7,^c0BMa=\9HaYZ>II\9.;X)aOHKIKYOYX4BK_XIe=
@I8U6AS,Eg#^&D0aIQA=3AA^]EQP<3LHbYT^dbF[/cVN-[/WNH]Y&V4POT20[(=Y
\TFE.>+7>XKL1fW[3-=YB)8O;QKLJ0HIXeDb]=76E8^Z/6O<6Q86BUJf?.9HJ-TB
WL;Y;<TNaL+e6-R3O./3VAAR=&/NFe_H@&_MAS\K+>_E/=HeeB>1YYOdb4-;e02>
&>Z6E+U0S2#/3PU?-He@>DVg9A/.P)I]ec9WA(aJd&6IZCL?>[94;4;,T_H0^O8f
#4RQCfHGO-,C8HYZ;KT>&#/_c+E^OKHKFB@gO_-[#WB[1?9M+5<KQ^C5MI-;e6Z_
cOJ@_(Occ:d9I\CXB8e6T^][7?=03V/8.TeN^@=132Y:TWaQ<S37WfF(T8AbRHY^
)FASXR]Oe=8fgIMaG5S=WfGNXNA5L.&8DCa2@IVV?5E^TWEc^5<X9P;[7:)^)Nf,
b-L@LZ.],I&a3ILb[=:dV1d.6(=e7Tg@5=<#P<-=H@T8LBK_S:eHAae24W_=,OU(
5,S6T,:2CJZH-J,GYLVc@O/ENgTZG@S)S6W?]R<DbTd-R1Z,b7c&2252OO65^bV:
6_<DW+NOcPLc>K24ddVg=ec-Sc::>D7B?C=NH-1#WgBSZ=U9<R01U7P<3#gO[1LF
4f.7PeY,[UR7dc93gZ[3][U;O32X_f1<3/?<B1^dF=?]Y/5BP0G>WU+_XgLO[U/F
CLb+>BS:7_W/8)JWMQG]NP:G[XWHAGIF#R8@F[19;[fICY>HQ.6)SITZc@9)P1a1
7Q)4EIW<1KHI@X_H;)#3PS?GLO5Z<X5&>^ef/&LS9RC.XGP-.?aXe7N-3@(,Kf>J
CE<TKKI^^YNfSP_2K#T7KEU(Z5E-S7+C=]^[02JUM#TORf2Eg3T4e)[&G:IVdLT&
A6GHXI37fDIXQXE>,d^X6U.HD/IG,.[C=+LN(,5g@SQOgEXbIgbd=aKDPOWW64)G
S#^:IO.0e\d9eW<0K4a(,Ae3fL?R?N.JYY,@,FT,@X:FN.[X09Mb.>Y9e^]f)4TI
&L[4b7Y9(C\JCVN;<f2)VA#8[R9CK>N6B?:M,&R=_C[&,+-DGTJcP&B.UA42A9EI
O\Z9Q+;@=WD[3abM)7DD(#CB]<A:,:RAbTa9aJYV7,OF4W6Z9HQ&S&,N_B,/:(a)
U3)&5)WMA23LGO+Og7A@,PP<e=&UMUTB?\Y\4e1ZaP;6g)<V_DNf.VL;N>f/I6.&
e\g::^PG+eI)GQ&-4C;VKg23T#8gO/=(H.eBQYD2OTCG-\&c&cLUR\g:Z3?4_2S7
Z7&Q&.1WScW@+]IZ4;a^EN91#BZ1#N229G#a49dJEH3CRM,K-,K72eI^UfZ[Q?Fc
(U6X+YQW9NWND3Seb/[Z1M)W7J\BS;D,e>G@33)c/7#J^QWCg3P^,WbDOQI.c:J0
MR,8Id.;^CD[aJOM#b56UddMAbO>Z\/F<KT&SOAT.-_\E@HaTQ0+#[b6T\AK>#Y=
g1-SK&-eFebQCP\:4]-&.UY4(+\>@?e,Z-B&:.X1SSfBE>b,JHbbfDKfgV3c6:M]
YRI,KQ,R/@1R=0-17ba,\7Gf:O/c-AL8D2DUTOb\BK9^S1Z)X#A\b@cL<acDUgX)
Ea@[L1?N&SQ8H60W\O14)()9W@1c7.(Nd67d:DB,26E406Pg1GaHdc^EFbc@fY@b
\ZPZ)9LF;&)C:#F4M/J435-P7e/,R.c=:H;3R6_b]3f,+2W7#.]ID=NFK<4&?O<7
1Df5g1b5YKC^:0<&_e)_8dPb)&G>f=:P1GRIYS&Gf?ZL+PgDE#Zf@A8-YZZ]CK)@
[@N&bDf>#Gc:C^EC<Y4AML;SOVN4Y0;eYJ/a7RdG:<WR\K3Dd8Cb5ZCfY[6;3Y0e
@E18>J+J>QZMb]H@;A/\&13Y70Z^g-ATD5R6,^B^^U[DJ8G9(,f/T_^R4,/\JTT,
NVQ;TP5#)RB8c;8<]f^6=-]-8T#,Rd^4+Ge9_6_)GJH)V)ZZ9[)0ZAQ=9aRfN[IO
71@aWEKE:GAMg(D4-=XE>AV8#.?U(^B70VTU+4^8Dc=0>O01EN5GReC,E2WJ67-T
S6_QTe8;YP]+e7ST3TZc;DFK]@;aCA\@R\^JCNY_9&c\.]L6gS?B16[A9&[;<f\a
.5IfHd0.8DU[_;MG7_1PM2K=f9U9C=^DYGRVTM&/>+:.G/>QF[F7A[J1bG6:_0e]
+Nafe(&NH,BQAI=;L2EXFT3ZJZNXN;/Q+_L+0cH7V^5VRT6+U./9cTX]c1BP<<\W
/,H_)DIa;a?gR8^ZCBa+3S&/7>dDTR?,90.@+[G(GG#AG3__J/J@S8)76eY4@RH,
f1SSH_0N[\OTCLC>GSETPeMN62\/(JIG-_FLN58,[_:8&e5+?gFX6I&P]Ae0Ja\+
.X@83][9<A/F:ZC,/7B9X,QLI7\K9Q0J6-P?)D/:=C,=L\=[0S4,\_7ZK&0F<8V:
-f[1/;8b8KXY4U0)?2W?cPK52K(DE[2C6Pb:+.7\a<EA9+81?VI<A4O_V+d;YBST
.HZ\0NCY9aZL<aHR/H-\LND)E<TcP1dbW@L27-69gC4UKgSH:<LbJ>bA[+SSZ]\(
9f0Ig&S?UOJW90Y+=4V1?CP&5(R\A\E,/dV_/[S@;T(/H:^>H])>86g_@WW,_#M]
X4bTAbF)<a;P,^B4:@MBT.1Ad@(,e-[2Rgg+a+::FT8E)[;GB/Yg9>aVA-84Ueg-
DXTV]dIQdV98E[<@FV:;aO[ZB[8LL@E8I=J/@OgM#],EIP8OEG>5SIbF;IC54,4f
-54f+6.1+>CUN^W>.[D[/WZGCa8bObDA7\PNY_LT1g3LZC@#</[ZS>HNH7S[LNL\
EF^&aG/+P5)+)4^(PB\,.7]Q_K[@X)2[Wc(@&dXV0d7T<\3U#fM,GX08TT_Y,FLU
7KM1afI8^2X[N&5>d,P1[;L(:I<d[/\XZEIO-?.DZECC;[+OF^E8-Y,=,VdGaD1O
BEYO4G#e=Q,f44LdVa>)3aA/We5B2S#M?&<=YP1>0DaS)J?dM^6\-J@29CH]48_2
He?GG_/9T:4LZ[I5;b1@Udf:6P:f20.J0W.Q2\6?7O#)GEMC#_0(EELO44?L=\1I
ZJD+EeOX+I^?,)7U7(4)X\GX.d<\KMFON0#fg?]DXA[LVL]W,9KaO3&[AeU<6c05
)36GDV0=W_)X9]cAeLBTH.Z4ac)2aXQ_O@M/4=OVe/Q7f<<Re]IR0Pf)Me9:dfT&
2\;C.+K.<-G9d-CdSSA<6GT3)-?;N]LH[99+VK15#Ac,6UBCX;c.5<ZR_-4)-AaO
Z=Bb;/8XCf[a#H=HET),EDGU0\QQ0[cTVDGQGY8>/O45@LX.:gU5+/75>>B5(AfO
5LU#4O;[0DScbZ-?FW9.8;FA,/2+#9<.2]F.9W:B=M,VO,UBgIcM_K)7@1R?#1TI
+&1:g4^a)SA[,CL-15XK975a^MX=2;S8I6?J@KJP1?.Z[dg>=9HdGcE=YFbTG/B]
P<6ODc;R.(d7JA4BJ5:NS>1/^3@SgC.G]^R-T.59\[g\D[?GLLVd,66>S\/fHTE.
XALLb,4gO<)X)5EO,0_4WM>LgJ\<3DWE1_SfF]L4fIdA=LN:I-c+3>8FYNKS_9/D
N2PIBd_<0I1&9LP.^JG-P)GX\@@JDbg+M.K=#Da:0#,WLII^:+:JJQGQ.@86Ea=V
:_1MM@GW,bf]2AD.&44]O40U>C[DN8-J?PSYG^5cCCcX3IecDC:-471[C0M0+OM6
<_&EG(1PUMbEbHF45FA^9Xf&+Fe/)+B^.+HRKW00G1e+2_fDR)gTQCQK4.QM1,Z)
WK8?EOfR^R@_:Na^<.ga]d]?fKA]D?DVF<C>;4g<Id>DEV^9eJae(++)YQ2c5X66
d:MWK<:M7GK<>fUf,(AA_LUQ:\b(SZE\2:GcMQZ6_QWN\CK/RMGda.JB2;E27c_G
,<2784U^R;RdTAOPU)Qe6@AGC&/CI<?0.S]=fdLM9\9]0ME9+FW@<\VNe^)Vd?\a
@Kf6T>PS(+?9@e#+:CaA?-4<S<4O#6,&3eRU-f9ZGDP>RPfb_H3X^M.HQ>8YY3R9
aT2cG@/(^(&YXIb8QdbE\FbW)N;DU7>^P1X2b:1bA40WC6U1B_E9(OESP.Od(bB@
H6=PE)66D>d.QUZAHQD^\2H-ee3-7L=\@b?Ja?5>bR(b=WX>d4&?=502)&P:2Y&^
T#cVZF5CZURU_2[dC&(aF:7X-.)J]VFaSd1MCO(KBQ3REN/I>b#bLBJ=X+//)cKC
=39P87HURdL9[)==U<N@=f9,Q,@H7IVL6fTaWZJL6T8P_F]U0#)&f^XO\VP#42&#
d@6>Zf^R?3VKd_#8T1fUBNA\^,,g<c8D1g_LX_^bN&+E?GHLaRZXTH92D:PdKH+e
.D90935QU=4]\E^LO<,)7dOV2+&[NC43/B]T4PZB?@YPN@@RSNP^Z)X:J/NANPU=
N6V5(.&-W?VG?.NWHE1cLU]9:fFd^9BYa)<BYBI1YCJe<W=@Z4R7.^7]g\_#UM:f
L<fL0+X;G+=8c]589H9#Mc668SAUV=6=5J#aO4TO#)UL4(ZgC,<W_\<9UEIESXaL
-QU2fCDG#[dP8-EMI]R^;XRfX#,VTG>OWK8aH-_5fcf/N2LC#P5]d&Dd4^]F:21c
8+FJCO@(O1b;/;UY;TI3@=V)@b+g6O>Lf)gDA[):N9_c?JF,9>[@E?BWYe:R#Q)g
RI]WA,^Q;TLOM3^#/C3#IeJ9F;99aeObZ60E7_(caXf7+XTQNbT_247gZU4F+(,M
S,eSLUbEM[IZPPUOM+1Ng?=3MH284_Q.SGU+AHUOOf]OQ?1SC,aUT>5+M0?&>b8G
3@A6S&[MF/Q4ZEa7NLP=B\O7eR(NWQ__caA@]#E=/+JL+_b4Q..P/-1Q6cZXW=OV
7:X&_4B&@?W47C@c?88H=T=Rc,Q-?P3AD1J(.N,:BbD41&ACfBND0D58a04d/NeM
\Xc?R.cOLaGc2_#9A9#:N_I+BX?#3#G?e-&AUXC(X:NWT-;/U(Z&&LY,S1S:/4O/
adI.a?(WHbM.e@I;BO?8JFO=QV.P8>L\-&LQI0Za^L,=LL@JbOK>a3>0ZX.dZ_8)
@N#\cVO4\@a]KU1JB=EP>H/PP9]H6(dX,8GID.[]&#2&>-][#g:NH124PWaQ;AAU
/:X29B#[KCML.OP7H;d^72GC=/c2^UNbOGP@+e^OW\(@_T:+fLX^^4c;2TB[#YJ-
\R0<AC5Md=]B[#EX:.U(P=KIbS=LdF&;,R,VYMEPN)22FDS+S,>B@.VM4UXO^:1/
ATVKT0,OZSdIeA43.4Sg4d\N+TDeMD2;T,CKb((N4D-=I2J>aGTIcX@+LKTYATeB
T2388RZSAI4.:&DO&[J]99-N(=[^D4W5f;8,]5[QM).KdAWSdP)5d\&4a=K9#N+A
\]E^Y[4A6.^.fTA3<X7^._/BR)0=Pg<2VA;#N+QE;_:We?^.Ub&JJ)G0AL=OJP>G
aLWDCbS4ID55A[U_=56]_6+N#XF,T)P0NKaf=X;e-HS#AHI\7TK,E\C=B6\ZcR:U
aP@(7T@+1I\18N0[I[c<5/LJe.62^:YPfV5JcGLAIg+Ma=K69bZ)+aA#dc.1Q[OT
?E;RS_O5F7&D-Z\.&PF-R:X71J,F&D(;gD1Hb=[&aH::\.d.IY;W7X_H,894N9DI
fd/YIN:I@&8YQ:)G6,a_J4ZB^=8_J1Q)U(-_26UObOR9Ta9eZ0Kf4/(G#&LI^(VL
+&Jf/]R&^M]Q<aS-Z]GaWd#/DH_:4=;A(45d+PH85Ba=e+A(-967EX3.dW\7;B=>
LLbHPgadBB)R\aa[.V_eR>6\KfB=(;S;#XR>E_.0B.IE49e;<RLT4ZJ0YLGf]FVe
B()MT7,6>UH6Y&BB]+J1FD2U&4O6TB7)EZP[,Y-98PI+Qa=<:>7X-Fe\E[)(e-J5
=)G;O_YV]0)1YP:I+J^BC6R=gVK8Q>^e6+0)]+V44(aDO[:B@SX;BQ8ENHR;NB,^
,@OE].<B;<>\Z&2,_IW:;beG.OI2?)Na9RWdf#bOP3f1(OeY/?:HS+J]e<1NTUKH
Of#5<=R)8dH[#CG5&U4f4SfGPg+96THI.KVOfW8VTFbYCbTN99gKS8Z[UQdVgZc[
H@VcCEgcB&1S4aD4<LRWO<T]E<W3RL2Y2TP[Y:H7F\5fdX9;N7YQ;9Q1DBQ)DcKJ
=JX8<eW+QE-/Yb]bUa,J6cK(5DG6CU<HSe?B,P+;18(ZF(C]B:T-TGcWcgfWJ2K/
@Z660P^?/6DRTQE)7eZ4D]Mb4-1BF^F<WNd0F^:E#GQgBL4.M_E]E,A[6K\;?c>E
E=7]LJQEe5>ZT4LaH3TNIJbSQ5gUL0//&)JVdbV;KLAQbU7fF/a_ab6f&Ld,]SV-
#OY)9-Rg9-JM6DS]Rb;N^d8K:a?6KF#ZL?+,+8=?>.LF#Y>S5bHT#3c&6a]K-&WY
O-U)M7N+fSb1VX><^0I(9dL5()=Hb9CLE>V1>fKHVBG>e=(:2:g3[&GH-61g.0OL
aG)]=Re2O0Y123[[V_5ET#-:Sc&=cbC>WFc^.D&2b&PdI:V74/3XZ^T_3J:F].OG
GfY<CL)FD/Mb;3g<R2O>N.O\I+R:a46=_)B@+cSCN>-9Gbe9-9:Ib:84MJIB8A[>
?L5UXX7\DYF[fERUf;LY//a0+<<^d0-a?=9M,3f]/faO(4B)W\WKOe.+NVS,Mc((
GaJ\E,190;MLFXBO<,5+>Yd/MU#/Y=_PLb=f^?fYJBb<>576NK1#0?-Od\X@D-&g
SGdaKBG#A6OM_?f:-L)7>IXg]^?5]^g3fLIP28eX[><7Q&^-08:I\D.^^_Mb(22+
:LO:K1L0ZYc,A(#BEH;]g(<0#=^0b]^<Tf&?gST,cNYcaQ(UPeIII(gSU4RFSgVc
12>#S?])0VAG(<8Q86TfXARdL_LR/&:1NEg@Md\KPg^]>]]L/961,?O724Q[Q-(?
a+=#fS/U)(H,(L;5-]^;?,;PBNL@0<<gL9?S_F1F+U;R11^>6dA[OK&=3RP@)W52
\gGddH,AOQ:_8(U673N;.[^aTfFT\f:g:^^Xag5<I&c+Yb+,=BJ=-#XBEI5Q:f9^
YF2_/0&R)EL<.C.0FUcZ\E^&C2P)(>=D.=#IEMZ4853:6I(&,-+^ZAQ-X+PWEMcJ
?O<E:HCXR\<f6Q6_R;UCE]XPF4.Q9E@TJ1eZMCd+W_B?2Z=-_dVY,a+@D+4PCFBQ
>B4\^&M&Q6AA9VFGafe#)(58SVgV^X,ZF&O8P?L:DCcUCS&dKXGYHKa=5?.HS&RY
d#0Ac.@B9-d[F;VP0@YK,<=P[^,6#g]8JdeV[2EIA]Mb(.AZ]Bc4Y^P0OBYZRRCT
:.[K3\UEDa(3:3^8bH4VcY\,H(?T=4]8C;c2TL>GD;+0\0O-([^4[X^EaOT,P:gO
:MTD=SL-IUE]Eg:Wd)C69_IBW0PF#J4XIL6IW]c)BK:P9>DfS.bC]=6L,cf8b^ZF
,SB-Y#)J3+J@?AW,gC7b,O?1(?T:3#6#J/4A]Z]U&Be3e?dDUO/1P,e]^F/GAMP\
_C;5^2UI/S,[;@HCT8[^4Zf;+6JAg3I1@SV9&eg5[YC>c2QPX+&=YYUCebb>#g6I
Q7+A<d>U(PNPG[4d>KA[bg5(?C,:X:SSFcXDJ5[88<BD+^#]6=Y?92(VMJXd_TbB
KWF?0>bHQ](I_6M\e17JM19\(5Q:&M_>(\Y.a.9OY)^T^FU8,ERPBVPY3:.:?B36
4Ucf^P<-aU1B/?QSO;BO3/e/5/fKd550@Q;B[A4E7^AIY:c#@HJV>I130.MAbHcQ
#W9<OYeK9Y_9DX/6AW_Fg32(PbCO.1DH=.=;AG]C1_f^,>0BFRSLA#X82d&T:E,W
P^GI:H#gY56A;0c7+&Eb:BY5/,a?LX_&5E4NL,\6ac:1Q]K.+^dZ#690dQP2:7D)
M?5?I#;(-C0DbSZV86]AKE6PX_M7<;Wf#UOb<RIO[^[6PIT<_EMT(Dd#9V3ScHf]
LZ#g:PR]gE=+=V>4IRC_(N4Z>CWNCRX]UO3D3f,@D[[]6(1.<S.49.],LZJIb-O5
?M1,[aO3553^cd+3&3M:5LZ]5FFdH#Y@FF^<Kg.RSV:?-Vc4ZJ@.R0C2d+UKY+YV
HH[5\]3JQLH]<).N:P+K3S-eG;:>XKQbLYCaNC;?/7&R^]K<T592J.=_^^fC;QM3
FKZG\&KNGe5T7DcAe]ccF74;R,A1G3<H+-9/)f<)7FV.X4DR:[A,,aPX[<F[YC(B
PXd/1Z>:^a:[gN9?/J&+8bTPT+A\7T#0INX2d5,?S\B52fa26GJ]JbNY8.C;L&f(
(B[+>MLFFPI?e4EBFE>DTLKOH?#N)Q1dJJc72:?.10R&gc:V4W8H<>Z>]F7RIcFd
PJB46f)LH,:[;@b1]G5U>QAZ.Y(2UWW2<-ABV7e;75;QegW^6+SF_eUQebbPA)eY
4f8C]\+F44[YaNGQ<LeR(G-(QINbXPC2SZWR-\@A5:f+Z6<@g3cL>U5CMG7N+,B^
d,--9#f<)VQ_=e2P:#.2<-@?Z5(73WCNU^eD=eXHG5eH3;;e[6ZP:\gF#B.8?ZR+
GF?2Kg>Ag+)#8B3dT68(A]DC0S/]=TXM9fGLM6cZ5>W<eFD>OI2=g@^9Qa\dFHM@
CMXB93STcb:(\=@R.aV&+/gFF7QQM]K(Ob^/Sf>P?bA&@S?,7YXN7HK9KI/f5RK0
<EI)YGU:[-IK<4Q[AKa8[6Z516NDPS5,GJ_YJIJc5C2),aZ;DY::_Dd:AZ;9@<WE
LdCaAb;CT,]V94/</<OPC[,2A\WU4gcIT)/[B-J>bQ4XH=bb=D4&JPV7G]5@3E#d
(P\g8+<12ZgIDJ?_d#\1e>&;-/[Y(I^R5.aB;(<=L<V;O((L#2@_T9@FIN(1C/\8
g93T-Pf9BQV-,))If8ca<PZRYJJJ:/_Of3]:40]5f@9D]MFRgVXGZ6Zb&ZU#N,:L
P>\N/>0+MZ^:<D.5gCPc1bJ@^YF3bBVP;M.FK1aL+fBZVcV>YD/C5JJTGPRCCZ2P
3X@1?-aW_=ZWGcA]g_W2YZT]XE&/ZIQa]?I+X_\FXg/LW1&<<Cf=Z+3F&>]LHW#C
B3JI&O)@>8.Xb4ZVB\R#E06+:@MDcfdO[;VT;8QgdcV5/]##bS]WR<RCL1eN]92S
QX399dRf?K>/J?C;YM:T\5A/<QBN:CFaa1N<]3a1JbUW6\8=GMg.6;+IXWB=[Z-1
[bWPU+EEPENIbY#-,^UYDKNO6KaL]fFXS>0&;(+bQ#?@6.9Ma&15PVb@8d-CJ_LZ
c:5g9N8A&3?LM:AS@53ZgGWa04P^dK4.7=D,PbRc@/[M]EYB;_I)6AAEf.4W7ZdE
MC.(Yb1M.^I<\BF(W2LRXLZIX>I:+HG5L[D.S97KW:L0T@@BfcYT:S;3U>.WM>G5
Md1_\1KW4D/+VM@Bea2AfE_;11C,17C8)KL70f+&5_WcMgRW_A#_]E/JGEg(=M6U
5SKMOLZ\ISb;(c;O;6A@YNe:d7#/K2AD7W9\GV;5M/PdI?^G\b252H+S@1LK)7UR
ZO3K)KY\5bJCB>Q;L_<,TK369&:1gae#aV0ReW2:RK&fW4Z[]-UL=O.N5Mc=JdWc
FI61&R8?O>XADHHB\#3gB,1<&0QWT,<S]ZWGVd02ZNOFF_]#2+G2?cPZ8AQXXT2U
LDJ_.)RUCcbeGHG3OC-ATC3+B-E7&aRGBX.L=.(H>GAYFT,YGV=I5L<,\=dK7:15
cR;e0OK97\0+(GVH<X;83]-TQ0UF,:YcLgU2[-FW\QQZKYdF1FRCgg)&QF4>9I,d
5aeZae[5&eWJ]7aGTU2XPA,gMYR4f]RRE87]>=BG=K-CD<4B1:eSUgZaAU9/ZK4e
N)=N,9+=922M3]&cT(J].9ReY\HA(S0BL&RGZ(4(EDHL(:<g0;9FS,QID/YF5C:#
]^dC;T.BcX)?eX5Q=?)R3b-Cf8E;d3S.(?Z;=TQGAfAc=CYL7Y?-U.A+_aDYF8A9
8HYf#7YYXG4+DBA\d4:a3P^JUE-2RS&P-HgMKHOW]>HHfN/OGHOLD7ICJDX8CCVU
Y^N,b7U:5^4)])(AZ17.^LLYGD<_,\YbbN(]3TaN@?cW>@M1>QM^KF_IF@,<:UM.
CgTC72]4+.L\Y\NA.e#D/6D+Q-QEDQIHc^)Y.L4Z\Y70@TP=3Db,XP,SgR>A2.d:
TKCI&LU8c;-?6>L#J([YN@WS\<c?4;)@PCJZe#;]0IZ2BEN2?J2^5MMaJPD6e;aX
4d8L3gaGLC#=]g[L+CBJbdcQ<1GB+E3c[Q^eA=D7gdIf2\dfVUZSOHX&+4e7@G0)
QIPYIEUH<^W(1B;F=31KeR9V-GLX8AL:(_:e[@^MP9)TSH9]Vg^+^QJF9U]BNII@
8Rd)8eb1SJ93)4-G/LXQ=5Pa1;Vg2#<e8--baQ]TPYNA8-8U)=<J0)ALSNd1/H^<
CA\T\VL/.0/G&dU&3Y_]79FM[FIFYPI3eZKP864(2A2Zd+a.&PgPLEQTRH=O5I5F
\F7F;N?Yeca.:;g<?E(V(RL7[S7W@AIJ)W&48-/Wd[_d6ZPW,/AD?3)ebMGO=+b4
M4^UO[^^QQ_c[1@Pd:@4/+BM/W3e:0MbMU_-;fF2X9HU/\U/5BI_=V_U47ZD+&S3
59832.-8M4A(V1gb]1&baV<X1ReTI4ZgbW3L5<@L:.CI5aSEZK#I?QW]>#._aBY8
\4UKO(F#3MS<-?NW\A5;4ag597]AE2]8Hc694Z]3LRPb?>F+N@;9,D6J-T.F)&Q5
W^Y#Sf+<3^G0_D]>5V-F>;MH4IJfKLNAHcY@@/7gY=W@-=ZG>G^/:GUJI3MI/R/d
Q_8P<_WM6-R3>2@8J:>MB1T.34+OHdd+fe.>[4gE_TDM?+6c>/.eD:,N0CKJ,B8F
^fb:f/>CXTL7AG#QU?7H#,O@MN(#G6A8gca,B5_d/Y7AEb>503X2<d\)YBZX4^7^
A8SCfM@TBZCF4_[?S2;g>)D#;^bA_&ZNAR(IB67;Se9\=M:1L+X1_L]_Z^R.J>5d
5V4VQEfLYM;]N=PGgV;b8I:7^cV]B:1+JS7SAW\?>\Mc]g2IaVb^f3dSK;Ke_a61
#gP.B.IVP5//=)/N_Wdcf;>=:5VQ,LTN9db/+>d?\W&_fVS:D=/ARO@06E:dMM09
;N-Oe9ae9G;]210_bRYUZS#.1X#7f#Pe&#fb8_R_Q>XW/U6cHKg>7@G2E1XIb1Jb
7??YH&T=M,<..aE\F38>S@12/[]A0S-J1J;S;1PE0ba4W\:9\Ef;Zg;^Ra?4@a^0
g+)1483K@71O3KN[31Z2)#0W2B3bYNP;#06@8KA\0).0.1(Ff>cfS&0-52Wdd4+U
d\\^<SLeG6EOHAQN2eJ6[&eaE5g6E2X?IFCKGaOE_?G9]I=@=-__bEf]UfffeVOb
&Xc\]R5XYWO+;beLdJ1@D&3Y,]We5CD>AQGAbN4eON#a#93-&;1ABAbDKWY:9c,@
?WXC+8N/^&e^W:WXX]IM#I[/LN.aXJGO8=^aG/O0A?ccNQ=c2aQIU/#/H:-44Sb+
+WF\\0;@]R@_<&^EOHZV#,9Z_eYV/Y;bO-O4,6,(X[)?bXI9_fAe^2<g)-?_MEYe
)&B#:fFIaQK#gPY==6U4K]5RWKRNHT1NOZ_<WH)\=b8e5Q0L18HG.9TZc#8R1[#<
WVP1T0g(FA@[Y25EYgP8RV-bF)S/IZU<O348;@CV]O\S52A8OJ/-RB=A5OK1P+QQ
J9d56[]BOUQ-&,O,\IM3S9>\)>+>YEPDZA^-(>5E0G[A&9@IO[RceSeD/;]/.@E&
K1b0QGZKB9]-+DM+WbM@IQW\T4EOZ:6_L-=WZ62e&>R:@_b/g@aLA@]E_3](6IRM
+;JKBd(+]@Jg(g68\_a7MdgW+=2N1SfQ4AKYYEV3YU/52&)KQU,.9JfVWLQUPdZ+
b#Ta28?KA8@&A5Y?_a/P&>c-eOD.5_J]Y-Qe&BMa1f_>7DP>LB1>F-1DI,]X@V[5
U+g+]Cea9d3&b(gceZg5X=T4M/:Ia\X6Rfg2b#.A,?10eSQN>NXH(c+8eI4aS[=\
\1+?41B(A^gVKC:EC8UG&>0=EeaVYK&H2R?T=D+5G?41-6]B8.<JS3SB8>_NP#DM
O5XfM.+32&,3SP@KSU6K)McfMJMMb=.d&^4M#d&GB#ZcF-38)-0K+4_fWg=7?FLP
.OMa+ZaW2[[IC=1CK)NXUC=SGgU0B,4d_b\/cF#1)=Y8#3I.QNe33<10H;C<D<EA
OCb,238gR(92DdB&JF;>CH\OU&:6V9TTJ+@+W?]7b^Kac=(IXJ^)RK9Cb[)0cFUM
gZ<1D3J:2BJP/#\BRJ;c_QF/G]UL5(AN)NGZEO;bL&&Lf-^NDUJ&)BedE^.IeaeT
-\J,aLYEMSZc(S2Z#]gXZX.,)SBa+C3R.8+V&):d3N[_6d@SS\)92)KZd(c.JBbM
LPFWP,<Z<W#X.)_Z6\bM\/K9#P-,G1H?X7:6)JF_:2TXN<U^NQ25dbV?W;b1)=65
[aO7A9F+7Z;Lf_-6Q[:DKg958FO=LT&:H&]#.T4b25G=]VR4X/_J2HR-.SR+;ZH&
F);b6FNGZI32-g,G^XYTD[IV,_f::6[WODHZ0a);5.AcN;]@GKcOTN8LRKP]:3,D
gc:;UHa(4.>OL>C&@SB2Def2?P@YEHdJDNZSg-W+#7bD=dM[LMg+JRaJ:4>M=-)d
S5DRgg0=EC9abeQRFWg06EV0@+(aR7M#SAE,7)cD)T@[98:7U8O@f=6&+Pb8)4T;
5KW2VH[9:P\D-CZQ-.EVgFaF)DQ?HR(5E?^1CRE&/0S=]3JCY7@@ZANeF)9F^0MA
Jd:LOY^1KG.HZ4a@fdCNaf(:MRPXESL8_ea[^NXBFe2,^3\5VeMS#f[<IS.eE);d
W\d6^[97K9R)0UO;I+W:W]D7577>6Y9Y;,9>H+^b.E19PXF1+LM<?)&)O7E1Z^.@
ODX8_Y8JY;aAcB7;/QVMUdX,)<Q.LF\0]G+Z]4ggXKBa]7Fd\JNUg8d1b;CU-5+d
)S1]=_#V4109N85<O0@:VVZ6@bES#8)Z^=>MNXQfE[BW6&37E&b3GL7EZUW-FY4d
<]OAC]/]LL2U9:)[a5#&)Y:[0PW(1=+DTeU2b1+>B4^<M.-Qf-8N>B#cUZa,XBV[
KHC8]MZB1(.g\.QbKA,e<B75\:;96FaRC62W=<,Y=PRWZME1d>b6Q;X=A8&Y?T<M
ZE(,6BFY^DQ-Ad4U-[1M4RI@J.V0R.:)+4SYc-,^gG5cCY;VE0ae?84gZ#D4g@/,
4+Q\Lg_-T1cH.<gWI8Vc=c,H+(+UcbGDWdg5Z>X@\0f;]>_=M_3DWKRDZ@CeGZ\(
/#/<S<XNE=7J-<THUfU\3SeOb\ggO=BNcKE9]S4V=LZV4YeSTa<RBN@QKMJe?0FH
TK@7MYVe0REN?FQQUHIT>8Q4#IJE(]6ILM).9O.?[\2e^JgSX4e(c_X.-N/(5[c6
d5ddV_^B^)#[H3e&L^OH=a<PJMggJN&]F1#bfS26DAc_54>50e:?,B/Wc/He[Zb8
a8EJe<QcFBVg[f^D:4&F;#W<8FedIKCH<8:XC855<3g[C:]&,=4@E;b:\W7ec\7O
@M647HO1+^BYF\9IegDVfgY[1VV:EU@QKZ3cgeG_@7EAP2,[SY?^@)<af_Z9e.R8
aa)K]?H&ER:FRA[b>F)3^MGgH:@Y,#K_HEVGQQ2V^KD5&MeD#<d0N/=TZb;PHG?/
GPPV[J3GCeO/MSAJGX7RZXQO\Y8KI@&M=PM#Q;cFMc,g_fDOWP2@MYWTSH\^@@O^
W\]J9,;W(Q^C-D)SI3cO5<Y#CZ6L/4F&/>GFPJMXH1_4dE);O-9XDF9dc1b>FI5:
-F6c?F85X/@BW2a;#FbMG#O>g</O[fW8M8>\_9O[--NZ0e:Oe_[P5<#4BSOC)_[B
B1)<A(L,0@M8#M4VN^08GV4=Mg4D>Q83)aScR+E2RT))8WdWCY1>6^Z5HWO(T:dS
U2P-J^X.6T,1O=Z@d@L_UNeaXT,aLHN<NLZA9Yb0#Z,2JWW>WZ:9ZIcE4X].Y/W^
D2-[GZDFD4QTHP<d#c@H\g:@2K)g+IZfMN@N?cLPJM@;Me-?Se-=YId.1:@-f)H8
[;LAS7f:IBg8.@Pf.:&cF-gdcT5gD:=c7Ya(0NSKCJfP9,WSGY8@K@_^7;Z54<G2
dXgLadI\gMK-[^AR#b>-+V^8I,O-BR,9=ED#:d>Sd)7Y9\X;[Ed1H1^S)Kf=1Z)Z
&ASLNZXa\AeDbaU1.=-YL@a7]:C:DKLEQGg7-+#gUTN_c4S^FJO7PQLWfMTH\ATX
_T[3QNL?eD-e<10T_YgDaM>=(]aCd&B?dN\V=C99b5^\]#ND8;J4+LN:6OFH@0+I
YM9TP64?LJf-BDDSS1;_4-TAI1K+>g[O)O28N=7Pc)g]E1AV/(Y7XdD.-6_7IOJ#
7/<2fL[c]e17PdBW@TbA_,3C_53aQ,A[3>1S+@R@>/R?&+FATf_?D#/#NC&#5T2G
a@0@5[H/_WI/JMcJeJQ9)#dfU70f@->NUW7LT&.\,+F&>Y;M#g.)F7G.-e4VfA1&
6?;VGH\;fRXRGE0W+dG74^JJXeNO1E2&>U4Jd(R#VWM<<YL7Cg:SR8#Y5,YKKMRT
Z,@?Ng95KSOa-)QV(+WAJYg,;BN<f)3PV8fX_XH[HVM-BbcTW?,#c.)0S&.?&>^0
,Q4B<H3RbRP(d5.9@A-f[[dgd3X#Ve\#4JEH>[NGPDI?L&L)4=KY<dC657@U;0a1
G9UD/?(8R.]>J/3.&\.\S&NH)QDDCA8g_(dB^Q9e,&OcQQV25L[>+<:?\@I.HQ<<
T];[0fY2.)+>8BD/L4T9UMRf=<22TVH_5_FFS2=0,B3WWc<-faAYM=SD=.O+RVNE
ea=MJ_ZFd9))eRg/LX4C^QTR>RRHWY-#)b7K5AGF9ZK3f/T=-=6J,=EXPEF-Z=OI
7^:([X4@OLSEDP5(?TSB<c\TCUU&ZR_W.)C^,&]7;#RO^/L[d32G@H;HDONWB6ZE
<T6;,Wc6L3].RV-_B(EU-GM7[g\OH0]KC6V5/IT/gX[ZWQZ]LAa@d4P](G6bM5<Q
UH74T-&JSa.&^[;:2J=UFSSERR@O7]b#PN5_NXb()W752[Y)Sfb2]AVcI9=)Y^JH
:KQP>@;UIGIM\4=V-,XgZ]aKFGGS@MZ<.Pb.:f^??P7;:N.gUN-K76QL./EWTBAa
5HV&=,?K7UOBIgbJ8<\GU9,50fS,ZOSDWK7gd)QR<fIY1LRb]7gNX([FB6BH(#&:
=PPfO=1_FZIe/4\,#L<[Q?;=ON>V,FNB22#]OF\^?;1b0^JH:N[9+c_;3LU]6f\c
48\dFBE3?[^_]^4P,NH2bfWB(5a@Z8&9fRggfLV^4HU]8=H.HYHL>XIg(>=;JR?^
^^HCOC-f90F_LQEHK<;BE(4a<7S8;?A-DLRf,XUP\?;FZ#T+(g\&f<a:)f.R?JKM
CQ.@&eUf>1&KFf&f)PaBA95-98XJMeb75>89<B+/-.0FbH(Aa1:5:0c#_IbB9(Gb
Y=[[.^W+V2W53<#]04X=D=JOP^S_VIFH4@R25<,d&EF/#BV:GF3Y<EDV8V3=:@XP
&=Ad2c@[BJ\GR_MeO^[6c9AcFf#)@=TJ+<f/=7Y4W,23)UTS^;YdRAM=N]7;.<.G
b/LfVGWOLH&A_8^LZ)AO667E>/9bc)g(c,:WANcLKI#+CJIHIRPI7X_BB8(X5.]\
^:B3X,J6B,Q^F=I7.7.281-\g&HRJ(;6G_d(YcLWXFaa>#N(DT6aJBXZ^D.]V[6)
<Z\[LcN-?JS11@TTLF1)9W5QM(QF/W0)gORSUf>;70J55-(6XG>b(G2FB_61=Z0I
925]A0RQJ,+Ud]W)g^S6@c&b;,]H/:];8Nf)WRJW>AP6/^a2B\]\b6UIPURdNVMI
Xc(X+C2TATTS97YZE1QB6=2_9A1:L9gJN-CW6]\5K=J/F#QD>JE=NJWJI,NM,JRD
a<]_ea_8#1^gIbPO:cY[DP#]S_NBdNX-d\NV/Of]#PG\g5JFg5ENY-6,UJ3.3KbS
E^OQQ.eC.1#DW2&JL;PW;L,f_YGec<T:MNd[4Z(;&BW112M/5dZ=)+-H5F&0JUcQ
_eY,1-,)_(W)Y?XgC&</e2\-&\+&7L^C&ILZd<6<dNG;[a1V#_&g16D4KS88186X
5TI)X9WZ=5K+2)&a(YP@;X:K=:A-Y5+PEY]TG8H50gde+bQ1e(#.a@3;&,3.78A>
(68d=5_&VRaR=f.A9->+=J/E4,7F9>3BPH?#)MUD.1RQQS+Dg1KPg6R3c/2J-@?D
@ZZ+S_2ND@:V[&CS?b,a6/71.M.#]Y=S?B;:ARQ<.GbDT(-JL)Vd?LJ0/bSR[A.O
Q;dOaQDB:M(#UP]NR8P>TB-/JIA)F=:H8UZaC1-eTV-g3\Uf8-_M/]Ce7fG,-FMT
c6Q0JAg7A=]#U3_H<@08[4JO8E\KZ().D2-U,<V9I24NC/#bI9<g.E11+Rg;d(B;
Z_eQ[g4#0+.R&Vd?Tc(H(\YeVXI(dY^/=d.TDK5\7-M-I,I40JNHAaVf@ad3\HW0
FWd/#f<Z3X0>.8.CbO2V<.aN((02.A@(.WB>M=b&JDK3QL2A.eD:@>XR6:AF+a7c
Md2]f:Q:FdAPAAE>g^ST8/:M/<T1T@e?0:DNY0M5Zcg,#Z3dO+3:-d&Ua+X4QL9Q
^fB7edaLfZ?F;)+7LQdXaTefT&Z9-X3Z&+e50Dd.E><e0LI(eV17M-ac[Z8S@8fX
Y#;DDc?]Ga6@6+)IQ18U@6gUW=-1<ad]JXgEXTb8SP-WXS?#@I./.0^-.M6=S5/C
JaU42eJCXGIb;EdMe=97]R<gEZ6B1?AV6^ZARe@_UdUE-[67/F.C.\NEVePPP9I4
LWa\_29Na)(BGff7H1/#YNagS//#;SfOZ>FM(A2-_)e3##4FH=SYUU@VV<N,^FID
0cQN#1_gC(#)-Kg/LcKE+\,0TageF;a=W]P83PdfIMdFPZB/B&CIUQfbCCfD^SRS
^>Ie^9R-/P:KAIE01YSOU2S.)YL_U&f1N[^FNL53&G1(SA&R@e88C#@UaM,7/KYO
5-a;MS&X4+<7a7@JeA)dNN=8.0C>1?F6g]ObEab?:_e.I\Q(BbU>[,RWXY+?RX_5
V&Lc.=.Z9VE8>=e=BDTbJS>,_E9>7L(XVJ[9.Tb.[CcFJRPQZe2:GI9+_(\T8U2;
N[3OHUS2dc(=7Ha#QRc#MO&N56D>6MAg+_W.dN4eYHd32-55eN4H.ROfW8g#:PL6
4fJ+96@cc8&5dSW8(#9--F?JBWV0UPQ,(f0dXSS/.[(DAAI3&IPG:(R1I)08X+?K
8d2]WW:,,00:gCJ5@L,1+5-fN6TBJQbFA@]SdAL2Rf#cPR/C^Z?<KNX\DgCNJ]dY
A7+KKJ+J86E/d//6[W&gdg,+@W/efFX:&\+QH56>cO:_K>JZ1)KT\,<F;5XBKaOZ
/a,&MK+7<]QS8;XU/8d_:XZW-5g<0Id+a7TKV[1eg-+f;[?9V9Z&A5f>MXXR)?E0
_f]HW:YXc<]Re>HO[Z[W#UIeVcSN/8B_DB[1=JLTD6)IF12J#=XQM++=339V-bHF
FYMU.Pc;_-YaT^W(c&;CZBa>aM@ZN(4ZgS^N#/g((-]I/8<Z52eN,V>fG8/fJB_=
D&eO&SNZ5QE9?>cbH:?d@T4U,.=7bd#],Yc]7P#MS?(a.#/-D1XY_U]RU6\GMC=H
CB6[Y2M&A3V=M-W[JWET,56?dCQCdgc&4Tb;caT9>F:1=Aa3(aRW+JV(&5O65=CF
:eA/58>?R>K\?\9eOKHHGR_[fY^R^>#IQYM-@B^<951\@Y4QFf@E</@Ob;:V((,W
/>6b(<WX1WDg;I&:3WdIL2IT6MGA0C#XJHg+H#YLP86];FV#TN]M<R_Ob3IWTDgY
,67FXfA0XI1R1IIeCSA\]UB[IB@9Ccc^W7;NadS1NMT.)RA:.[Eb__UC2Q:2I:e+
_J3U^2E3/B&4]T4-A8J7U:Z&3Y,><GCc6LNU]ZN5/,V2O7Q7-&e==-4TOgg[CQaW
L04<]cU3WGY0f+LK7/f2;EOS8K6[.?^&HOgP-J-8b\=D2AA?K.CcaQ9bRV+WEaX9
Yc>0WW-Y3MAGB]5W9-.39F.]cHe#>+<a6-PDZW04S.3-G(#]]VAQ3EFBA4D#@BBY
CbQI?1UEU\+=6<H<TEgFR(:ebJWOY:4Y=6Q+I[EU]JSH350#LNDcSJ;_Yf0NOU_J
GX4N]=>9bVCR.3BIVd5WEK.b5?J\/.HJ63bQ1J>@T@&1&B_O]J[0b)4EW/(1^RI[
aO=A:gg/]c9Pf_NPJ^_IH6\:G80PJCP-QWT<\5A\c/&UBaAa8N;Q3a,)UVX#&R5U
4<_,2M7H8DRSgOI<3-CWT._3HYSLXU:=)HWg#\-)Y8L^NWY+=JQ.:MYM4[OONPC?
[..M7bD(+Kc.8YKfLgI@=D,,9/3[e4G,1a_N[N:,___,#Z8A.R^bI,Ja,;&?SHH+
?++S9T8;7f+^QfV=;]77Y8KdX<<gD1T6Wg7WD_Ygd4)KcOXL.a4/2P0>O7Fc4dJB
O+.K:90BC8N)\79dZ9.:E168=)W/<=G=dN27.VgTJf2XDV@D79SbZIGU5.MZ;/G;
0&BI=a,:N]2AZ>^0H08PN+;I.WSEH<Ce-YgS\-P35VD;[G):W,;HK+45@@1&1>4@
BH.XL<#)Uf&XDW(5?@#3PVG:,LJ?>B(e72)&2b@_@:S-D@@&D4O#J.]R5e#FW87&
TIH\S(Q1+Hd.#P==G4<#>WGK^@E5GOG23>Of8]56d>ZdH<BXe\cQ^)c,X.bRgc<@
dVDU(]QQIL1(<G7,PF11e)4]45G(^GQQR+dPL)9b3TGSH^?4aIfQJRegTa3CY3?R
X<IgEA+FM1UO1JFd[]<5:Y?435e_4S1^2LS^0G_9#f.6VP+R.5[S\5e<[_@aO3<e
,d+>1:3f,]RG;&)f+f3>FYG0^b0(Ga10-f_^Rc8@I^QF,&DTcX:9>Q=6Cdg#CP>g
)(3C<<L[,2/@LV)KG7S)X:afRefgY4gG8YK0baZ9CCM5W>QcNOM^Gd0<Y^?K?)MJ
,N)OFFf>eELg8+\fO06@Z)T=P8C>;I5@O@P;aLIfQKO&Kc/S^D+4ASG=J:>;[g&T
0RRbN2=/V:NVU7TNH@64FZG_Y\R=U01_EcRPB8N_+O\;)SLRB830-c>Id[CV/7gT
OXFKSg.eZbYH/#G8>G9.Nd#?41/8V)FU@735\Q.baa&65[H.L+<-c56g@^,UTa,9
]T>S>d-@#4g/-H>3=D:[6aNZLA&UX9/8aXD\3SUb)RUU[S0&T0Q^YQ?@gFc5,S;P
TF&L=BEF?BO74.RQ44^4?gf?UW)/6:H8#8.[S[^E)W[N;7>]Ge1-QO8^U<e7_S_6
&2cDcaM-8>(cBAW^N#LT,\_.TJGA@&\@3]YEEX@bbBTA,c##2<LECKPM>FPG-LSd
c[AdG]8NLXF-W39\T,?)-1:>P9?PU61L[f#/05f:X9FY8QCdM\UP@b7<,EQL0PO:
7Sb>-,4^VM+U9&dP-AA+:[70IQ>,L9(<1;^6YCb1LP_;FCc-=I&4G6.95B2/57(6
fd_8?.Y)TYH2<Y^&^K\K0C^cAK<+BKKR.,R^,=1NVQ(XTW/96+4Z[=BNT6e^&+&/
VQV[.0eZ_;7(P&9[H,XSQZ33;cQ79b@dV?<68aX\11@.PN0,&dR(TFD_\UI?(]Ra
QZXHfg..26SYHQWN&)bd1(3K2[c:I.;>?XeYK=LW/3Gf:aZ+WeE@B&@Z7;JG2_J_
0Y;K>/].DWAD+2GA<__=:13bE]b[=R\ME:b.BACP-_-^W,8]3NRJgCDd2S@IU@aR
_U,TCUGdfY#FYEAFX,F@O?JE&RRW9T,Z4Q\3Q[?RHBg]<d)#fQReg8_5SQD<C^K;
fS<=>U02b/,0]:VTLfJRc\MGDF]aCb/YHJ&TRZ\aT2J<Ef3Pf?D0LB/Va]=O(C[]
Q;a?0QEF]TA#S=]FVQ==-^?9/HN+,OK:A\D)>)MSF1dL:QegHSdOZ<Lf&>Z^e9BE
X1-NP;X15>6Y(^-57TDFSdR;A(9ZV,/a=V/<=\g>(1gGOf(IG,MMcGX/4U#U9CI_
9TBDbU^FS9]B[M8=(YHO,#F,/)LZ+PgJW&3c(TaR]d-FV=6KO^6B;G)Ha3E5@=/P
#7LfMGQ.4VCKLA/gW:12_S_e,94C?X&1[?ae?R@e4>)427?9KDR5dKT1CMQ1:3X_
;9UeS:\Y4[LKeEO2MYOSD+8_]:>7)(=e+WH;;W+X+:TOFP(P=)HB4Z5dXa@;DGBA
S,CX:=KY.PeFHg>_)2(@e)c0/3JI4LYAJTB#]SUY1_cGBYQUULJWFZ.;OfeQ+.g,
M^34=<=3)-&PFeVc2Bc<?]N9E3EZSe(1@]_F&MS.eV-B&)QbaWI[/4.&Z?cWf)Q]
8]TJSeZOMLPd7d+&E:.82Cf1I;Va9)JFOB.OeQPHeWT:Vb)417_Z:gLPVM^WRV>>
59RD^\,N-RNO1XTgb0-4+L@>6Y<2)&LId><,TM2B#;dc=FbQ;CRI?#)GBEUagX+e
J.@BF\6Z67\#LJ1D+,WT?52XTO;b4/dE;C7IIBRAf>_Q2XY\&(FXN/YE;/Qa[;bg
e[8X,COe+aDIZXNT]Ja36CU,2]f#/P6<Hbf[2M<JcJVF[K2<V[;c(+QT^^bO(_@H
&.D<#T47]W4a_^OH5+1&,DU&_/7\</;3a^6VLTFEa9N&JVAQ.DV7N@;IFM&VWZ0)
E&/a8eNDR.\6OM#aY:?BcYEBUCH7:P,;9?McX@caTggI;=X&907U\V,X.-ZAfPB5
c1=Y?d5Pf:1He:PDd3)71g</@-,Pcc>#)4U0EX-\):8U_J@M;T-;RK<VHO4ECG)Y
Zd],TLTH):@3VBWUL[F(g=FM@R(\cCX(4GdY=0@/_C]>cO30&2BbN;d\?J<PJOe:
\>W?2eWGF^2?.9,^O8X?-NN_c/H_Lf80L[RfSe^/4RTV7gVC2GC2SXX4<S]2H5,F
G[>#SBC.J[O0bH,0/3Xd2)1fK16?@G:X6\CIR^(1D+(K&9c:H)Y4R/5W=A5>gN#<
ALc-4V/F/&E#4e5X[FGZ]86GfZUV(\(/4)8\fC+8538:NMA,P.6+2UL,T8/fb/,9
R48Q)5:1E++;8,^UdDDPF13@\gf&RT.E)ZA)-]e@_JGcDH9XbbgZ^-/\O/FEERWD
;^g[^C)\E:aS#[J74.&9DQ]IH6+J8:5B=N;XK8=_c2b:c19A],2WBMG]6Se;M]Yg
<KX;++)_2N:1M<bLC><6)g?+]VJ^(HST+)&e[>OeHZ5A1dgKI/PJ5c[TQ],NA5M9
+\I><1d_Q,A=c+=5eO1P(=Y+>E0GDL&060YX=b3;dINB;SS/S^W8R3RKFPHQ8K7A
=_ZaE4:7eaCd::TDd,(-A^Y[Z(UV-eKFG]8fc,W9GgRU+X&Nf[/cFgKg,)gQJ3OF
GfUBOe3a1g=P-g4>bd,/4L6<P5Y)XU)VPLJ-Z8T:=]/=0>0_fYZ9WF(=\0dYT94.
c<-V&R:WP;IML/:,M:\DLFdaSUD[FW:XdGXBTJ]</#@ZcO-c]bdSQF4L1a6>Ke_P
2;&3LJ?/L(VZHQb<H?99gU1I#bKTNcY:\BP_>,4^./(&>CS[O=9ZEc,U:HTATDF+
1OaXI2HF\Q</B6EOGRM(cHddP?W]X:.A9NAd1I@[gDA6b(Y_G:A-<PSW1gJF83U3
?^G/JKL[D,]#bBO_;,Y6#3_JG+Sf_:+7CRB+]B+C1<6g]:=(-.dHVa=E[2)DbXcM
db5AVA/G>Xb5Q])=7d.-Ee;BF(ZgQ->C+OM(_(H1CQGgJS](9D0fZRG@NQ&0C=R,
]d?4Qc,NGf<:,SRYUD,3Z5_IF&S4(+/_)W)VCC#5EKCBQCOL,Q2)Xf=1TAH;<YPV
([c;AC0CZeD>JeCQT/(^+N+e:bD7WBHV31acC(EMgF63TO9c4,&e0,X(FC:W32K.
M-#1(8e5e[6aA,eKR)+@4ISYR-.4#U+#)eD_(QW,HJNPV(N+#CZ=aZXV3:RD^#g6
YR-P;fA+-RNZFf#AZ^M#?O@a/gSf+3aP^Ce8/EcENe2\g(7H.[31b0BIfB3)XKTC
4&ACPQ(VdYUN\9[CAa@@dJ7YUG.dR?9?Q(X1K9(\E;)@?2:QX]8+\,C_fNU#TXNM
\VC5gMSa_;#GRJNW?(W;OP(>3,JRSK>d5QX^W^TQY>QQe&Y--6)B[fR/5g;\WR[]
QXNNB?6IJe[#GMe[?:9cEeG0,:Ng<QN/MQ,B.;;A8/)2)e]F(V;b)STR4g,EbIg2
=8V-U8fb.7>ef9g64KEP>b:a8aEGN>E/MKZQT,^L63(a[TM+CT/@11;<dTZ-XM1I
4#;7H3BgXT(@UI<dSb20+]>OER<Pe^X(R(<Z_+C2\6J=?Oef09VdSRNXD.,U8#)B
,^<N19H.3_:@b7I#,AB6f].eDBeRXD/G:(_Z,g-ACA(A=(Q1]f:3656Y-D4WG(N9
>c:F9fWZH2HNZYTSM7>f]=U2Qa;L^0X2eNR1g,^=34O9-V0cWW8L&S-;=SLP)#5(
JTcddM-TQ+):TQ4dDdPLg<-#C]HAO7]Qe3]g4cNUD#<RJ>fGJ@#g.ScYKV:=#M^D
:/d^U^Vd1A^8H(H,:J2dL#8],D:d1\8A[aG7XZ>ED[AFN<N?Q<G9JO-GJ8:V-<+a
agI\3P.fO0T49:K0KWF,eB4.?c@5=)ZagX7a=W9Q1-UB.[5=JTH4\FRF:3M)723_
\GSXVX<6D,;a>A:J935D74D#,)PAGPP^>UZ]WEO(>_X@4[+)CO?=?Q+5d6Ga)E#V
2AOS4-NSI?&]=CV([+3[DcXc[=]4UUWH#g8bH];&_Y/MF:S894/UF.Ag&0_2@^c<
GIg.9S8=[S:BH]3EO78UZ.c/==X5U#/5dF<^Q11#YHdF&B[N]CX&HHc?Cg45cD4P
&[X=@<H-67GO;g^BX2T9.f+&5#1Pe)g8(_9De4\FU+K_^LM:g]W_<Vg8#@ag,.f.
&fA4Bd=f9<F)L:M1>3QE=8:YC^BAE;0NCZPB>:QOIf7R(6a[6B-IUO:8;/\_5dD4
4()]:dYIOE.dW@/FG5H4@VbY/J7bFDUbgV]EY,6Ud-]_0IP6MNbX2ZZ\S],/c-Ob
7+,Z1,A\REIK>UD]^bM=:+NLZI[V4H-EA(_OCO.U;^b;56H/_YF[X-If[TKAQXZ+
aX)CX:0^?7.ab8f\-T+F.US522[36ZedU?fJ&Qa;:/dL=39M0W7@?==bS^VWYHL^
1cfeYDOB,2?_Le=O9@d9,=]N-@?V86GL0Ac)3Zg3?3W-9#/@;g2S3T9K/NVY>ZK?
a64b(8&7d/\^<0REbG^.#^OC1>FBe(:I[?54]];\abK_41Y2g,N#/E4g#&8/]T)>
aKPPOd3dH6Qf#UU-A5gD4;ED-YN&^OHI/3fH,B@?A7MOC52]2[UO\U?C@,[[YQB=
F?D-6MHDG;HV:;Dg<c[X&C?^P83_91/89I5Uab<8c\6Bc2?(bJ(R\KJ>PYNC\N<U
N#D?.d(]dT1I#A/9HVFG1=1bP50K[UAC>;2RDZ>[PPa=D6:gf#N4@Vc[2cRfa4)g
0HaOVB>f:Qbc=dARSG@G]\/^T#.>8HGWT9.^RG1@0E<^TO;JYB4HV:^MO78^QE[Y
#GE)/9M]4FeHW:V#VU_e>eTBV2G?P=F:aO4IACF^aAA-[<C+Q[MZ-?K)W)SB[)]-
Tb>B7OV9.:>(S@d\.9@-]E=e8eb^4>2:G)\2;SUYH&P>^NP0?N#Xb^-(-HBM5=4X
I=\-[D1_cfBQJ)43Bd/AN>N#6<gGK/M(dC5CdIP#_Z?K_N:#KeT&NZ.<_?.+CP3H
#-#dYOE;Q]UbNW.#,38##37:^;^PINY.=_UG^^?^aS49X0[T+\.d3RWOJ<X2=9ZL
66(#OZ8/.V@KgZ72[0Z<d^>OdY#cL[E<gLHXF[Q+B+UW?O[^X<6AM&D2K6bO&,eO
_2#9?F(OKa^>IOV+F\a-FF-Lb+c[gQHAP?PW(DL6CGc#1,eY4I79J6_G29JKNgc0
Z<9/QMP((I?#@Zd^MK:O24A]Q<DK\^<VF100AS?9f;#U9-^2+a&ZJbT,6E:bH90.
-0\EVIIAg0OY)PKR11XB@9aA[_WM9/W6]a&PM-T6;?[/H;<4cO>E=aQ\S^VH[R=S
ca=PT?/5AVIYOaZZ=b?-&YE-[OV^RL4[@]YS:ESZNN7M<GYWR.9dLOLL-XBGGBA5
bL[QFV2@EU<)]WNEa_A==\9)X(D+bG(9>eY2E8<a3\>)ZA,=27J:7#+44]b-1V>6
F@>M_)D+S9;bEGEEdVZD<adgaPYDF[M21W95(R_aB+1]0V)M7>LY2E;N9M:T(_EB
DW6&<J\<8,C7#=>bb?V71EfKXc8U&HDYdI^9]TgcN+;-P9XVc#(GF#J]HBHXRH&b
5\4D+5L&L\[IZ33+0V&F.:C2JLO1F4K94@XcEKXPYB_eXee:_KCUC/TC_S//X/g>
M;G<_>>/BP22NdX+)99:I.V\gI;\3Y]YVH6Pa^59>A,1?1UOFDBT_;)S@ZK/eJg]
dSW4:#g563:N>:KG@XYU-ETI8.+Z:f6NSAF[+6MRFQ3[,GYIP46d&BNK:\)+9V9E
_&],A=F8HZAc3JS4)Oecg-+W^J+UR1T&aH<<GMBI#X.#g:V36,58U?_\.4?2,BF9
C2\;V:8RfbQ:DNO?)EL)PMQ-O^^Oe(#,N42&&=6[c3(Tc,dceYb@G5cVd:H/,1MX
0d)A.K<7J<UO>6MOWgB/;2/EJ3NL#J;Ob_RMa@<)I&(\;1:<G5(Za?>Ad5+UHYKa
a(5;PbESee.PdQ/X0.&YJ4.(=)+8)]Ma@Xd<5QdBcDOGLc@A.(C<7:6Z>,YQ9\#S
]dNS>+Wf=/D-)_B8H8676cS7BRULT0b3T#^X[OV[4?+\?AQff::dGB::NQ=Wc^QU
QB@X)<a\TI&D&^[B_cP,DX<.R)Cg8C[Q9:.]gRMfH/g=4;Y)&RE;EWO/&:Rc#YXQ
WZ,]?>?0HbRcWC?#5F(3T_6XGM3QF[aU2SQc#E</bgU.YgFX4<\Qf4,E8;_+>0Z6
<N1EA#UbX[OG@R(/J8RY_2_TR\d<ILTPU5d392cf9M&PXZ<U]b2@T35G=c?)YgQM
VK/M6E_F;AbBXI>ZU]46K\+32&_W.H/^[6X#3Wg)(\J0.eac&2d9]^MM/a5IRVa0
L>,YTf,dR(,P_7//^O:JTBKNA-\VKQ)Q0f(CQ;>UB7.4]1-47Gec/PXH0)]2_78?
#f=JR4H>^=GQL>dV9&]GGPL[_XO\B6(ELE#B3S/),d5[+e)GIHM6bOYK18B58[gR
V-DIg?<1D#WM)]=\RFEgbL:eb3T1&-OS?6B9SMSTO;:dU/7<\/cA-,ZKI]^Hd8(F
=+YE6(3f;+CH7U8VN2[P]#E/;D>A\df7._4F&d^2;C8H9MP^_?AMTc=4T-.?PdNe
5C@?d)+8N8/GDgY1/_R@9dI.57@&6LL0#+d4_8EggG&2=LRMLga/V?8_NWS=\E7K
V5<=]BZ;J9CgWP7CaP^9W@&08/eg=EJ@He5?6SdO1TI^K:eRQ@IP0)Na4TWdHZ0-
^5COXB)5:Q^7JNDfA&BKCH)aTHb2P?O5?0Q0fY/9XRP?U1EJe[<T([U_3<I8HEb[
OBUf1,Re<=9[(M)V=S]AX+MN<L8FY&gI+26_(Z8H(dWD&-c/,fHd<R\Q)f(YF7<9
a41dF,(gVX(\#fR)LePA#W)f\\eR/&8edIGQ,G1G1_#T,>CA;(8ae\-.TXE;>a2(
@9(1Z#@BeEKK<&Z+U[>OF;#3^L?-N;_UENM8Z[G55H?232BdWGE4XAONFS0[M;TS
Y1Z7ZS21T&_?>#:GW)]ObbdZ_-4#)O+X_?gOe&AgcW?_5]25f7S.GXUX(04cR-?0
e(3)/,BA):X+:eN,.f(C^.-GW027HHWDRQdV,0S[J]2V.F.G=^7GX[-_d2@,XLD]
_AJ2a=4-e279>QTd86e^YT?AN;&WGKF4Pg9RZO/84KLW21KGCWTb#6KCeR<C:aJ,
>gPg9)NUA>GEUPa\1\b84&Md67NO^D.T=Tc^;SEX29R4,:&fecUZB,EOBI1-2\1U
NRd.&M]K1I(/.+#4BHU:V[9IGGaQ-B2YA_g>PEI<N?Nd90_HZ<WS/K/a.([KTKH3
JH?:JZb;529VP&?<FAPAg1FB[<7\@NJ##fQ@#0.XO\+YH5\N./80N7a,3/g#B1E.
3B/M?Y0WL?^C:<<>4-_)E7#.N9E=Ta@])D<O[(N@>03#Z]TB=/J9>gW,._cWf;Jb
ZcRTT[HXb@W=G,4#eR34ZBJ0LUR+PQ5+1b&BVL+JY)OPP-.##\2&fO/6TEL@1,Oe
a-.558A?C+UB2gdgfYMSNZ7OdV#>&&+=0FK/VfIaR]C]:A,5EM&0MN;W<6+IKg4/
b#e\U7]E\C.Q-adGf4O7MPW5.b-65(6>Mgc?IWN=4&0N#)R(M=MO.WA43A0HESg=
MCP2CT>PYbYf6gT=Df(S[L<eR]fBM:DV2VN?<<(?2)DD.W05\c.I6),/8D]K.:gI
cfe/C8/D\+g0e372)3W@g:D/Zc9aU#OT;]+FW3b(?.91R(Z6RVP<9:\)gN)?;RZH
YU2aCO?8]U::KA#6B1SY&6Ogb38C)J3EbCRVHYWeVdJ+.J)[CW>CF<T>38g[1&N>
POV/NRX^T9X(L>?J:/9;=c=<_SQDPHP0B;]I/BP/;R3S:6]MI=A27N33RGfAQ<=P
_KdL<G\B17W0#dQ=?_7bH&V-(3:LgCSbYDgZ;)A[(WN](^@B)Vc7J@M.[_UQ3)L6
>+.=#ed1OAR>b5fa,>+P9/[CO-ag5b(K[B.UOPPW-_BK#J@/3B/6)-FQ85dY?<-#
F<Da7P&/]7M1Ke^+a3Z^HNT_CEBM2Pe[5g&]?<fAM[KeQRIO1A-fA2P^#RO#8,g\
f,\6T.T^#Ra22a,2O30;aG,()[CW+ae5;>GD]UO^T?C6VM(eBaIL<1GR6HG7&WM2
483W6<gUEA6W#RS\(6QTCFVAL)DIVeH(,N/b#A<B<^,eHO>^[#9<@@&/(2Z#X9F1
=V4@MGXX4M^IKECLA]T1cZ8VRVObLS/IY2@;8:=7P3dS3W/7AYB1(>J7eX-bI4^^
C:2)F]\#E3PIa<G#?,0V0]Q6\(HAb1/FfFLZf^)W2LAdS7R_GXcD-;CF50?#599-
g0.4]_B9OI.8a@MC>S)O<=FE7V:30WCXBN;R_IS1SK5fcP_cQe.&L9OGLP169fSb
D1=C4+J/@UUE>aEJ+fX\VDDZDVER:gEG:CR9#Q0_F0Y>PBfZQ7AJ<9G5LLOI(cLH
<K2dN3acUT>X5MbA;WSf[gA#PYB(=9]d&9T)\BVBO.F<_HMDKUH6>YC0SE(>I3]-
M7)/DM1=CB0>3+BbP>(R:7A&WEN1(ASGN6(N1=gI.E3VH1_HF[OB-/EN&/eOc6P<
T?MZQAJ+GP.Gb+6(U9-.OdQPa<<;=F>Y/A235[)T&-.5^=]+;LOef/Ld76GU^aIY
GYCXBF[WUW,0MB]=O;&gKd-K;&L.&F(IJfgNL><cfT463KU_(Z6JW.P;b9VAWd;Q
QdO)9MaMI=L5SD7AUeE.7+B2W)(:/Gb64AG^/YHG(VQ9[eIPQbV\G=[[&5H0::N6
V<0A2JPG#R(3c::1V8NT]\SB]C-BJ1b.:fDD:IX666RL4EXU4(d(XVb37E8:a:,b
WNfMG[BPHT_1T,fPH[>\E[AD=eBD7V@0NU:-4<94)(94a5Y\?bCdcYSCL>c(T=Zf
YdU1A(SaH2@:3-c#g7(2(fQK95a#0]:dTfP\>P-/VGE:7@IEf9fIO.4+1a=d,::Q
C]I(M=AN,5V>F^9K/VKB-G#aM7fFLOfWLS1a<X23(XMZMNCM((;aE/3B@/.gfTY<
2[++TcX=bHe>0M\9)4U)Wc5FbgI1+:5Z9fF^&\_V3GS3YL;:P-#ABII.D1KIF(\X
0[Qa?(5Ga)32]V>(V^;1C<WQ(ZZ&\b[C8H:MKR_F\Y]>&R@^#gg\J>PH?)>XaO:K
CQ-#)N8(g^M?3W^@(.a9F_;]VCT:7Z(#M-aQR\C/?X=U5HOEAdG)SE6V>d5^]VO;
WY:I_OX]?8Gd)GL@&,Ug0GEM(13C[6f]X+U;2Dd.BK.E1cTX#HIV8C4MJ45aO,^2
b-O5X..(Je#+,+T]deCg;BS3LTJKVXIJ8RHGV3GP>CLUSI)0TUM5SA]LU;MEdaC]
ISC1AT-WEc[K>eX?6XH1@;LU(661&bPgOEMBb_TKJ1bBb>X75<f4_QGGGVZRCX5E
9?ZRfdWMS&]KY6CM8QRJWQ=/[>@ZG\[WQ?Z2DB7:+N/RY(B(JKK?0A[bXTgZ-e_(
8TW=F_5L][J.?]H9=:L-7LbG)OY,JWg],U1:M<57;=?[4>+#G12e+a1T3I<BQ<5,
?TXfP.,(E+#fc?_(]<MPXJJBC[gYffNG+S)aSIZK88TV[]^AeUB8;?ZW#_TB<;)C
bIX7ZeN]3_R#T/_c24NZ.:PQML&]7>JO;W;;-O8,Z(LGU-e[0DFA-\;-+NMM-3&1
?59IcMC_4OA]UbBXCH_AS&)\?I2Qf+TY\8\Z5K;4\ZO[_1-_QV)PXRX\6eBe8;V\
<ZM75d=C8(1.dU/.B<e+E18:d7/;/X82.TQbSF_WF,A+J#5gTV(/6>1Y\A_[(H^\
X+F2eBN;aG=0f,4)R2^DeB4?T>dC1CAH@E3JT@0JG,8B-UL\T0C+AfeL5aUc,1Z-
L6R<]F(aL5<<+HG.VO:O>VSg[SH0ILE?Nad@JeR1LFV&-7VZ\e>1GHCG4OO7M[UZ
7/&E#X5NV(TEYacFYKK+RPLL?R5/(A<:bAa?/ZaHS7NCBV+)V4Z26IRQ@81_-R&J
&)9E(#cG4dDE.1^NTAOTL1TG8OHWV@U(N<J0F:UM/Q\P?Y4UA0B:Tf&LcF6PHLI2
aW\.g(=b,7U)dV1:#(ABH=6EEDZ+>:5>AbbFJQFJQ2/VGEN[STf,-ZY1D1C&]NaL
?GM4UJ3<7He(986N4?Q[60+TPMZ->FG?CaZ,(Q5XN76@U@.@SF5VWS22_B)=Jc0^
8gg<S9d[Z.#GIZ3&))E7I>?XD:>Q/T5.S4e>b1RRZ[]1DP<DD?T]=&ZXS1L\gaK]
HVb320BC,]9HD/<@-6U,P_Wb1PEYEaOcX>9P7)3VA00AG^e#02^,X?U=#0,2,VGb
JZV8YIU[RJ>I:eMISc0FcEWe9N3GJ+,b+eU\M#PPF3^Y&Q.GGgHXPBFc((cUYQU-
MbG^>d)=Z5KFDag2\QAO<&J?-9T.a1CL>TI=W;d.e,gJ)&2:;bJN??UgG[+46=B0
&ZL>#YI9eUCRfe_QgYe5,&PD?2Y64(X+Z7O1Bd2=&^6COPV<76;,\;?_2E)b>Mg0
@6+=(B443>2._C#=A\+C+dD93B);fC8/B,MaIbXW#_A;D2?OPc\e:;0-\+X;SDcV
WH21Q1RXK#24R<3OEU:PWQ4ZWHb&Z1D,e&D8+cOCR:fNX]U0UQ;-]Qf>^f0#+L8#
S6OeY]1WGS9FWVBM6M6#EC[38RdVA)d_NeI14N_FP_]^@L^)5dX:?^[X^1a2@EZf
?1V9g3g:9FIKfWa-33Zd)(&Q65V+Jf1:.7V>A_dG]g:^Q_-W]_EON[E]HMYe02)U
6:0aI.DN]Q]6NNWeecc@1->\(dU5XC5L=I2VISgF8;E,E2O.8L+E>YgMBF+J@C@^
;F[fA>^.;5^ZF(<+4KZA5)53Sd[X(?#AKI^FeV8-@B6_0BR^0<>8SY9=#HP<Cc92
J]4J^Z_a(d<b483]R?P]J@2VRe<).?NgHA;30PNHMW4,X;PMXd_S[BX]2F@OB>f_
6P,QEW,fR\F.\[QD;b[12D>acJV55M>KN68@,?dW;eM95b65Ia4,.57.b5B7:KY@
@_#Tdgb\^7,2bd:VX-DM=0?;.T>RYY^BE[]U)Af7C,e:Ff-LabK1OT2Id:.(_@ga
WTcG5G&aaGY7]f?NC(V3ZX=AI#N24^DT3,fR1,>Ra=R8E[Xa+@U(T5MCG;UX<cQ8
Db.PU)#5D[L43G:1+C>U[e=L@F=gBKE^:-eG_-W1/(KWEg@.I;+,(T0M_CUf;BOL
db/8GBX8UbY@A&PL]IF?fG9A3[_CG8I).Y<?#QW+R3)&fL2)CbA]/d@X7\6bA=aK
=&e+E)9W,RHZ+XL#Z19KWZRJB.E^ET=7:<S)5F1f^X1G:1#d^fF-C;0f1c0eWK&M
-LG_91Q.,b[BcfTYb?NOA#&RZI+6HJ6+2AJf@-O&[HIVc43S-GV6&;S,V]2U@HZ+
&7925FRE2U/QfJgcET+bNSY<V_Q.+NOX>MM[Dg#eH?K=0/@HI?fM(+4\XP3DL420
(D)=c7C@N3/dFY8:J;T=)Q(-R?[L0c:NLgVK.PGMA+^e0Q?MY)-R&O_1.Q)KBVX.
#H^Qd(1,bCPf?dCHKK=-X7[\P7c+._1:ddB_Z=cT8S&+QXBO8U-#&91egdS?QU0/
ZJC>CGg.JMK#I5PON;.^P-)>U_/aJF(F:S?We8YXM8>c^QVfT;\bE.#QK/a>.?\Q
Df+f:a=5(IXNa7O(fY6@>5CQ7OX]P[CVB9f0.Kb(OO)4,O3GD(F_^]2TH7941#EC
-&Y]4C\QC1/A5eX^&b/Q0V^Z4E?Z#?T]fgVU1)cd[(Q6;-O8_-19/4DA;32K0aeE
D9F??CFX/15Qg);+bTJYA/P?87;@Z5T:^[BdPB&d#T17B?MHMMYV#MJT+Ia..fIY
?=3HQ)G4N@HI:d3F<>WFB72JI[c7@:O=B56Wa)A/@>JeW^Pd2Y(9c]=LO.C/#^5P
^2DR5F.g>__@d54JMK1eH2P_(@_D5E4[TE3a.XIW9W/Y^7>FSXc4JW=U8fIgG@(Q
F\Q:G;eg,RO-e+.G>G63RI/DOa))MP[W46STaQ(((0>R<cf1eIM8SO7W@C6.([g\
TM\@+YM@JQLNMVaYW/1/bJK;Ic].c>X;6H](RG>Bb&JP8RA9dDT^YCX_;aC-II1@
a&J9CGg1#bbU@X/O7Z)\YCWD>YQaP+UcXAU:#&Vg_e(fUGK<dNS;APCK,7(L3@bb
@9HQL)VI/[A+V3RG\@L]aUNFH73cM+g0])aINXcNL7>FP3=(/fY-OPf?4Fg3=8/.
WT0K31L-AKeG6Bc&)U-NXeI>3VA7f]GA<J_cM@U//-FI1KR1@WGeJ6V(IaRYB1:4
787)4;fJL/MO2#<6YbG;;8(N4NObD?1fDL,<I/L4.aBXC;Y3PeT[HK(WT>^8&7D5
KOF32)/OaO+B#&Ue2+\\@R3\DGF=M[7cb=gRKE^B2MBWRXAQe>.<]2(a\/W0H3G5
&?0L0>UV)B6QBWU5W66dG)SaW^[C7MPG?Ng35QS=,cJ__DFT.9A@2Y3B=QQ(.8D@
NJ;VVO0;8I,O5\G8KgP7YDgV=K2+d.a]NX,>FHLLaF6Z6/A>WKdPb;Rc&O8.1FQ4
\S9(&,d=aM\>^XE=b/L6CY9.5=N<J+H:=MYU9Z&Of/>T(K@^:<Pb](IPLMCgK./D
ZE=C5QH+2?34.=8IVOWVRAf86dMO[K^=D/FJ+.<6H5_>KEHC5cIF6^4F5UaH2:4b
#+,AUF1O>#G2E8QTUGf-QO&fJ?<V]:G=1IN25UN<.2S]dR-V9\?:5&:S,^5d)^Gd
_M[aeD5aTJR3b\3gL7Sd4F<#SIbdV.(+31=F=TGb6N3#/F@]\/_(eZ&GEZg\[:U_
Og1LNeX\3A-:+f?FBabGU]9?bBZ#//H4Y0\@?0c@9&YC8KX\(6LBP8OCa@=TXMV.
daPdEWXb)_BFOFR<bHbBRWHVa\CVcK<P,Pe0;4AJU4b,>),b?CH.7>KA\gZHO6P>
G^Pe?I1MM+01K&_6Z67ZFAB8SHLb<I.@]O=^4dgdS-KgQ8T^a@5a,\AK:8/aZXBP
[c[?6g(HTO[9@A>:B==)>8Q,X-P_S&B@LaI7\CY#Z1\R:^2Fc._RYZWQdIY13[?@
IL18E05A-&U@UYAYeBAY^M7/J.@KEG37e+&JV_/7\-G,>=cDM37T#^DS&4(&+WaG
g1c40G[=06WJTT(<29N+,627-.4+[5,^?@EX]:7:bZ/D#ST7UC>+10a(dKI@,168
)S;MCCGeQ1H_T-3AOGD?;P4IEc/<2ac0EFP6T\H,b[P?2/e#96[Fg.\\1@Ad?H^D
5^YX4W_YD5\F&J>fBa#Q,[E>F/T5<UGfUPA?>U<Ha)W;0-Zg6gb6EU4S<JYcb<Ya
R\e?&03K+=+\;ROGKg)::T;Td;E(^Q8=0E?0O[Z_A?.]OVEYHAL95eeUWf;8ZJF[
?DaE,@HQ3R;G1cK/cCIa;HWc612A&-_:SS#-A;X_6^=>4D,baH3M<g;+_]QcbMZS
0]_)5,=X7#8LgS;]L\K]B7C,e&48TD?XI>9E(;O7&]4e3+PAITf3\UF:HRfS<+ZU
W?DYP8#3K,bN#Y.?.=Igee&c&+Dd5-B5)-N(XIW[0\OE6RP5.OW/>MXa7EV8+4#X
NZNV9^#\/e];]b@D<P:g+,&<2GODcQ70@:5;T>7^H6?4G@d:E8QZ_UD=.5T:f@Z>
=EJff5?N>_FU_3.C^3.+M\aL1ULK<@BD]-BEc/MC<SWS>B[3V[>FH]BH9gJ1eZ3[
.Bb@.aA:eXJ3YRUO4H6XEg\;;KC3&M-4XF.2?/M;/ga^=-(:Q>2L.VE:[F&F8_=1
aQeI5_\dIJ6]KWT=NT,;3(K<H11CZX\3^5R,N-4?IO7[a-b377I55>EKR3<)V701
ceCMP\[9H;3@0J4+aJ\NaI8/V(Cb?I,<-Q4+=.&8dJC\X&=><C4R&2aI@5J2cM=g
4fI&.9+(WRWA11O-(g;,_;R]NUJAOJO&K^VMQ=?4bRbG:HFUO8NKTf7g.3^]B4Fc
;cH2X]036dJ4e#(K80]0\JBJWH#e&[fR)P;:P<GEbeW)2\QeI<BGe^=He+4[X27F
WAH2T:c+\6(FV[[W9H-E1;;PBPS@TH6OC+e;IfL2F&^7(fXbJP^+W=:14^O+^6.9
4(X^KeLd.7PM8+&<I6X:^6g>37Wf>/PI8<X9V;10Y(O4JfRc5P;4c^@TIE042S<Y
.:/6[06QB;R[#R?V^g;8?0O+>a5PPVH]W&#)Z\PJ[CSC\38#QF@,R7e[f_1\FI4d
J>=>cYa[Ye;]3g7Ne.c660f5\g;Y[EG]+4(E_@eUZ44.5#(+.UK)F.,/cV[&U#6Q
MC:eB0\W6\G\#&H;4AegYcf5NS\QM-_HL7.S^_(/37_^edSQM:(9GCIT(/J=&(c_
IHBe^7]TQd?NEWE1eCXA#WII3WOUEMV)c&.YI92GFAc;T5d+EGSG=J@C6bR@/RQY
GRCg+P<6[D0H=]^3#VI/\91VT_8Y8K84.g\5.KU[ee^2dP>JTb>70IV491/Y<29Q
V-Q([7+P<_]Rg2&_76-2=9EO6&OFg(16)c8@OKcRG]5[cTPI6QY8:4gG3C[5G8YK
VD)<[6e8<bIQYW^FB+gY&_T#+Q:BULAWV^HB+HZe=WDJ/Z]NLdF+eXeD,fQKO)d[
4,F2\>DWRS.MEK.=aN0<[N010GMag_,SMIJLJMf6EY,S0<#cOf=29X^eF-]^8D:E
SI&I3-a^.\CD&MBQOD\gP4+)RJQT2=?.E=Z4P+g#0WB/HQS:1+C6f^PP_<__B54\
\H(4[K?V.ET=c4]3(D_U6E.MZT3\\aaR5JbT<a66;4Fe&_0<AgagTZ<Z>NA6N10&
AF>V:e^4e]B=>EeU8FJLPX1ZB\@1B_]B+V,&4^.ZRH/YY1MBZCVJM@MBB,3[,U\8
0:=9V]?Y<35OV2X32<-eSXeNOY3STdQ-ER_,[D26W(CID@SZO,<QACZ^Q:WJZ-LU
T:^/,W#YIg,+[Q)KgCYefH:J[/3CA@,a)/I-^A/HB?+BP+[9V.?b?OE:DO8R0X(D
FQ:S@->e0+BEY\@ff7.(B67PZN&SWV4D<F(<Q7MX2TN[T@:-e-[GSU/5V(2,K.36
eb24EC3DdYa&1U^H:KXFU@:LS>:N+SOf=+JUU/A]X?O9#I)6B1+GC[9K#NUSSdVa
PJX6CPHM4]&^eEUdZ,:f30J&?gG)PJYF;0F<XFS(JAfD<&\<EBa=f@;KfScTQB<e
(VI_B@Me=/QdK]4R>6HgO(dL^S8&GBJ?W&^6WG[aaK^0)/.=JS\9E7J;4a_MQ#Z9
4U+RcP]<PJeCPg=AHN0W=e,B)PD7FL]+EeC;T^(g97155^N\a58U58DT\\0HgP=<
0\3]60IF_CI+0J5^@Ta+[RQ104E@beN2&&NUL[<7VMeEZa[(_:2+75;J&U&_QHEP
5aB/1K#^:AT\+g]#Y-)#MNdIb=fWBXJ96Q\c7,\EBbR/GDe[7SQ/M4ECgY)VJ0QP
Y&B@1^M.I@3@W7TAOH&&.I(.J\c)B(X)672.+&&ec)@c\B-YA0W))VJ:@_4dBZSd
6ZYgR)d.:D&aPcW,00B9VU#NMDC,),?]N78LN@gBR/KHZKMP17IGO:J[.8aLfG?(
dG2+=:)9K-Cg9\(O9?g3@d/>&01&ebKVMf#Q\NG.&)]UePO^>R_KJHZV/-@eRb.]
Q7(;dM<];.;IdQ.K&1BI1?(AHUTLaEC/V\>9[g94geL;e]HY#R62)UWSaGL0PbFS
80c[],UAdR[CD^P/AN?T:F?a=/ZA/@:-=^#&BV/-,M_U/HdUODb)=)SOII&g9Df:
=bB;X_-)LA9e?F:+=6=@Y@ZCS#4POMR.dGZD1--M>VX5/4S_A4;B0P@[J=:\eBHF
Y,9@2ND+e]#Q]Y5>B4CP,8\(RI8YUI(>:f,3ZQ9^e?df]b?b><Bf9^,X[NQ>g<f&
YKJFU82VDV3#:FB)g[31(:A]=G<;Q+GXaU;R[W3@UF0[6FK6R&EVQ(AD#((Rd:PN
;4::UI+BFQHQb7db(/IbU:O19+J4Ub?NT,d><LdDIO^JFIPKE8Wb6X?]U?QU13SM
NV0e==CUbY-IT=_V5_VEdgaQG.7R#TQ(R(=I3CXFCE,)V,43I@f7B?A?CJ[Z[O-K
7^(M+(8IHVBPaP,,g.cPe?HNbI\O;[ZBC]L)d(8d3#aNN)M?=D)?H,SZ#4IZd_3Y
<Ub<PGN/L>A,_4<2U(de=F>;dae3-dIU)\X^:3@7bc#+TRM&L(ZT;BF5e))f:;N#
LD#]4229E0Q?R\6@;>Yea]A^A/2eZ=eKab=gTBg<F:CK=PfgN,U1EE-Z<_O,G?S-
eG-)(VQ:Y=?9(9D^M57\7[eR2?Z0g13/P/X+BUHecLg(R17Z=P68D0-=YKeOT)^J
,/82UML^.8g;MFc+9e?I94AEBI>VG(9FIYf&:fe&:6LOX9@4[:?b&7UMb5STNHUS
M#/MY^B>0UfeHA)YNNM#/d:JSY0f9_I7LI=bF=S=Q#HSS?[ge6g#7C8X?M9[DP3Y
R5\#[eP6]B;\L=SV\Vf,V^@K.G&.VaY&7ETI/ILFE9E+e[:):K_fc^6KFR&.^.OD
L4XBaT)UT=5W2Pf[)3X:cA&+1]ROc)4Y0bCUSB;DO0P.FZAXO;ZX(H.0CG7SVAMf
:Q2ZF-5GPbM<Y7=9876,:)?D@#TF@7>,YFLQD14)bPWI<?ZAa<P_KM>WYe;9>VNG
62OSKd2D=bOKUA:F(][#b.68L9P.:.7),#0\+>Y&?SSJY]WK)c06#N<bU&QNQJ2,
I.^#+Wc_U#21Z8LA_9VV]ET(1dVKcON_P>VF//e33M36Ba.\J0CQHgH+AULF6f7e
eII&DgA/2#;VQ@?,@H5&Z_9.@)CTLX;&UIZ;ScQLeQY1;;4J^GE2(^HVHR70#_1[
D0GeZ)JU=,G]Y4a2/7QgJg32[UQV4(RdE322?6;L1(5#CC&4e806VLLU&+e\f#\W
=A-XbW/a)@Z5=Y&(V@UUHZ64?8gU44Pg0XKLISJJ0+C#6)B=L&fB@?YPUHL/dR-9
Y(HD8_>_I14c?FW,(P,P&IH+[,[>A026=:_N0a3#/3G&,GM02_f_e8=;1N+WOZ,c
@7K@f:=5ARP0<T2(a,5c2Aa\I_P7g1CA<P-.TK1+c379F42OYWYY,b>CQ]eSSdAW
MO]2?A&@6f^[\IN;B[XU\=;U\;J5/IWLd+-BH0Ce>@OTSSZMfWSSeEYc:g(VNN0#
L:.K/-5UQL),K/V]?X0BIGK\@ME;P)=TQE\0,e0]LLM\=>7JNF7[W6LOO;AK)7)7
6(+[<1_J\9#+@V-9=31_?NG6G76g,D3a[+HgbXdJO&f:JD=HGc]S)0=LKJQgI4/>
1@(,0]27Qf[d9AS<6/U1<;<)1__g(+I;-U3<P]KG[?AfI[/19&BAab[Y0M080Wa@
;.<;M3#VT0C3aT_KXeW\2fUa8Q#7\[4bKSQ.\:0:O(a9;dKKW\a>^&gRTADB2)WE
^/QV+^5_U;Q+NY_J7Zd^;3AT&Sd?BQcdd](8ICT7W=_[1PBUF5HS+U_+c#a/UX<)
?P4[_U-&4S7RJ-:I2H82715D/QG@?[;PTK7PUK0>Kca[:=KP.f#0^Bc8\1;>?T4=
>KMK[SVHFHQ/X:^1dga.L8+CIRP&NR><VQ36Ea-c5B>0X\K_,4J5><)^bKK<\;b)
SI#d]SgGA1YS5Vg6:P2[-EYP@T4[W]VA/6,3G\/=_,JRK367@AN)7[?UACc.K-RQ
dQT<.eLGMMPOE+VK(DIE3F<0U9/2(be+)D]\=9c/00TTQfE;MT#GZ6Z=^aHPJXTD
:,7S>S6c]E1PeV.UPL1POQAZ_]cN.edBD#fEVaa&@#C>fLNIE+<dNf2ZdO9L4Zd?
[1)WaadO>=PUJ)>24P7^]bM8KUGC^9PWCgY89e7\fKA;IJ?+_bcLU7_)MP;<7Z<c
MUVNcLdR8:-U]>ERF,a]>cI#QNJT@.LQ6XGS&I\Z^RFB9VK1K@CU@Na<K6V)U[0b
\MC,LC:BIB09TEN[4T+2G?2LIBa=Tf0fdQ(Ce]X]QNQbT0AA[DMWB)g^+7Nb?07+
R?.WHU]=e_I34@V9JY4a]8:f3eHW_@7YTfRM8N+))RH19+\H\)cD=097)>?=\G(G
>d8\Vg4V75S]KCK-^7\N=ZI&.bL:ZM&@12d_gfObOb]ZM<PRIP[UW^3T2DMIa)RN
J]9AV4YYT2M-H[CN985CafX0#R_:BQI^0W123BIYR/W[)eKZa10-./IC;e:RIU_^
>MS5?SMUPV/T(]19IKG_=_b3-RW#<f\2&RIDJ0@I]G]E#@T3b\HWfD?V0gC/,2M.
5X8].?TbID_LJ.\5J/MIHLa>)T]6cS;g<)b+[Q[L[NB]2\^MX95:MJ=:1\U7+SEO
:2L]W\\V)SPD>??]@8)-Y<W>AcLXLOP?==U:a2WV<3Af0:Xf:F,PIHb<K)N452)]
A\-.,(A?a[f2Mdf70.NTI@bK>P:=]/,4L8:/@?NHCM>a,TJ-?QWTf^GV9?ZT.[:D
c2cJKg_]H)>5OgU5N)b,2^II;aAL>6;dKX);V3CXee=5<cG:NX4U=[0fH\[e)b47
NcKGP=8AR7)c474.^?Kf.Eg]/3Y]4UXd=H[ffF>VH^cF>ccRggYV3J4Mc@<HBb.D
VMW>ZR7^H6&QQDg5S,JFBHgM(VAO_@^[+,#=Ub;FP\FAY]Xc_bFF=cIFW3EG/[Zb
>0OIOYHb33Q)]g7GE,cXaOZA+;aZQ;JYXS-4T-7W(3<_3Q#\8OegWV^9ZP4=D[4]
I\JEF:?Y&W:I[DDB=N+/_^T-QeWDg1#ebaHE^&JABd9\]_d..@T@/G4FgT38MYK(
MR9Ve/M5KdX:?KRfU1R>SAf63#7H/:,SaRM:YZV.&Ig24_F<eeDZGTA2QV@7#[+/
6BF72L>26^Z+Ac#<0-OI1g2GCa-(Vc(TS7A6XG+PZ1CT1-c1SOQ,]@\P][<GRcHH
PQEM,e?=1W=PEL8=P73(#ZBID)U&_FUg_3Sf\8A)[HZ>XbY.S]b#(-090CN#&#67
2G]\68<R4WT8+>O:&=)>,9G7Kb&A;Ye0/V2BeEGA5f>@JA]E+c;De042eR_FQbUT
^D,L<VbAMK8:3.B^#X<;@U8.Vb9QSM/Y]+2N)TYae<_0a8Nd:[)CX>>,UMEYSb_4
R964=@Y#T4RJUa6MORIS][Uf.LQ;Fg1E6CDB\97Hc@:b#5B[K,GF]Q,PPLY^-6dY
C2K#f;^)32Q;gYWZ>_;+,_g6/)4ZTYdZU5/X(G<#[?4?S9+T]&/9&T)68YOQ:1a]
HJ:E=K,9<L/0KPO7NJ)G>#O9.\)ZF13a]c:8Ab)^fZ95QUI9>ObSBc-CS>JQX()#
UQ9A@_cU?)Hd]K7&5&e1#]6KD<c(Mcgg/FGP29A&8I<VD4-4PM&8TeUR6R=<<BS&
<KNDUD_>d&9\gODd5\Q->\W[\@>S?,4QgeZ(B8d4/)\H?E:][4@T\6>C5:,C@AMS
@XB^=KgC\@@]I;dOUfZ1\BIOJ+BT+a6;3T6#\&8DTSRZXL:/)dfZD0HWOIe))KF5
]Wc+C+ZGdJ/]>a]O7H>2R04H4@\\gW[V:\B2f(bYbYYf.-<BM^>352G(4&OdI\>T
TDb/(:I07f+_c8F6J^?1FB#\_^)@S=IO/BA1^DG,:KcI)e4[L=F5>V<7d^XE^+L1
]B.R(N&bd88E6.adI)#3(7.PJW50Cb]#@(Y,=bN/abO?WS5.]315W6T5D.-8PV6C
f#dfNE?@<T1=?1Hd0S<?_e(UL4NN>5AM_0)V+6eMg9][X=6472V<#WORE@K@ga/.
M+>B3bE0]0F#+ULNb]O5d/0A6f[Z)7Z(3N1==E53FU]AI=P2Z=YQC7+gf]c7#O+e
)T,Q[-FS;1-A52YDaGDdUNN=a)^CY0A@-6<+fQJTL4@DO?#[BIJ>^).;TK8.IW_Q
[63P:E,&#OMdZ18<g]8FdU^H8,Xd?W@#PT-7<EU65P/]>?4WJN2=9TgKadDcf(ME
X+B+aWfd^&F93dCB=D1@G&8;C+>T[\(UPdXAZ][bK7ZA<X^-]+3(KB-.19<9EA--
RQa3T88dXC:d^,L@eEeN,]4(-#\RJc:a1X-<A\:1])YX(JcX3&WE186XQ+3(NG-@
8ZS&:B735G.BW1e,MEUZ<8?aVd,S[H]Rc:-&f&7e>e8b@1XZdAW8PLdZdLS^SKQ)
\Q_aSG(?M,9W:NAOd8L=+16?7HYP<.fOg/bb>,_R)[3&1:B,Z[U@R#H4H(-710=5
^60J\:aM4@_)^b#T2G88D9)&Gb/I[FZ7Xd>4S;(93Ub9@P,<K<LIMSfdg1UO26S)
<=gGY@B-<=MIW[,a\cQY862b7PMb.F4?(RJ-+5dR7TH&ZZ1V#:SQ-B94aLaZI-RV
HAM;HU35#:&RL^1_=4Y.7Z[7S6&;>[HLSb8Q3g9b<BL<@a@gT(NNS#U9/a(B_9XL
1WBXWS/\[bM-MY^S,JPJ[+PX&AS([#]\L^?./G>H8X>51(aI_GLdf&3bN7M>O(S.
,7Z]KB@NF)&@aNEW,1D:ZGS)@(7^JZ5A^=P;NO83L?HZ;:OfbJ:#@V#P/)IW)+)^
5OaP7,#ES<O=5HBVTMHHAa-L77[PN5A<=.8F0=?^I84fE=dO^K57>dS4dI@,@@WH
7]g\1#MI#VQXLT&dLeT.M^DgF7Z6^?3<bGAEDg\O9)Y#Dd0ZZ5]&Re+Ob0A6\LA0
;KC4@V.d^2HXNVU#WcD4ac=^6H^e:eH\[0R[^88#2I)5L-a7INS/AHabC)>[)L[4
CO]Q2S=+:2d&57>#US_WO1)gN]Tc5>22efHQTaET7D.67A?\#=/TS7AJ8765>I-C
R&2^FLg:92^YR;>Qb#dW]J1bZ^JLROR&bO5_H)TQP]K]]/Da8DgU63R]4RcN+&J^
.@B[_&/e-;D@;CRb^>281G+4268\86+HR4F96=Q>SWc@UH?MTAS\8@WGb6Lcg.6F
c(f8bdSPG/a7;5Yf=Y-^c/-X=>ON/I_.G/[Ld3/E1gAXX/9&Ead:OE.X1<P/WT8J
fCH?]K-cbS8X91)+Q<VSN[D.CSb2@V+\e,7.(Ug5.DJQQAFI,3g3>^B=-W6IA&:P
\=VC=:X4[R7NF_<HOPSM/C+F[f#U@Y72P\LWe#XF1bIXc5;1d^4D\1I&\HaI[W2U
1:M3G1(\Yg;(&>3FPUN,E/JK,IPOZ7GXC[)J>e7H&?D87:=aVeRR]?GZDS,._/U#
#0/[/OS?4gdM<T,gP>OW:+I[VcL9?&./S^[J2:<e<A]B@@9AGKBYXQ.0D9DT489S
a8eM4\\A8(B0#H:bBI_D0WUCdC<KV0cK_=8-EM1GUY&PgXfWI_c,HG4F[K[YU9]N
0=:J)[AORIG;O?g&+RGSCCe5J1)Z__C6.]-=,G,J+BC]TZ,^@OE3<JOD9(b^I6=A
XSJ^-?GH#ZM2L-(T=.7E8;G@MY[\#U,S/&F7E=GKC4:#B,MGIRIa#(NOCdGE)?H2
H,]M,+)[2>I,8e&]HK1/C8DA]:<710SK>VGR+LWHcbPD4g6Pe5RN(71?XV^7>aG0
d3f3X710.R.=V>4PMI/<6Y5D-)(b3a&:-Mg.3K7U89A2K<#2@+RG=W.YCVP4WLZ;
@.HI9FeUT[&:4;dG(PJU\AB5RSHQ<-NP[KX31A+W\A6.(-1QOc:R9U<(H/AD;#<>
b@J41;X5;\>1@C)c5I&gU^QMONGT=eVZ&RFW.6_S1C:/MdRC@/1&P5Q1<>dQY<NZ
d7eZ.;I3W0>,d\+]8]HVb_GI[S4O=J5g?ONbX&L5;UR0[-[9#gRdP>7JU)AS21VC
;P-POWcHcPD0SAD_WFW&a-d2JBO^J9+/_GEG)A9:WF.IgX6ZWEa&QV<S@C:1:F08
&3g@e37d?_.U,/,^5e>8ZQVV16;BMS(Q5\=ag7AZd]>R96OXDcTL2a=Z^D5IBgBf
(&>+KT\d]PF:#LSYYLLY#T5C@XCV(>69RNQ:HOO,W/,AB4KL^d<:;>DRUe]g#gFe
dcDH\2XR6,c?,5@9@eH7R.>ME9]7,II2Z8g>WdgC1VUKbG+O9EQV)G9W:_d+NR;N
eU:_;9Q.JA1OY\VdK)\fc+a];b^<=54U>=aK4H-ELEPRGM/7>S4^af?B&XDXg/R-
:,TZRBWBW2fT[E?3>4T_RG\JXf:\aL>d67(>)H/(E+KDU59HL/14eTT<]UI(EN\X
fg1A5?/eXCTS@C#?aS(ab\G;cEFO1^G62(TXI5_S2V^\=1@C^PV)6TY.ZH&=U;)(
\;48(I+e2>dB/9Y>PS7E.eOJPESLce9TRf]b+L55AYW0#99M6?H,:^U;6APZ3</,
W@8<2eRf><[;bGD<;S#fg:M1=<R>+?>JQROV^T@K5S0Y34JZde(#?QeW-<?/=&ON
:+M&A5<OJ;LKB8d,5I9F6Z7@\P.b0MQNL.IL8RG7b(,;VS^7[E9KL4b6_/4dWf^6
Y=W2/>KMNKDV84#BPNAa-E?7B>DTE_U#e@;A^C1C)0U<JW),fdW&Zb-GIKP.,&BE
[bO^J)Q6]@ZXd#;&FE_KY77+9,UAC[VIZRFT,Y+?9:FUD<0[</<L>-K2B^bL2(fa
f^[g^NN0+(9)G/M3:;cJFWKK)eg:\SXT3W]2g&^dc].H)?BYf,Q/7#@9ZEK5,\R,
C_6:\S?XaF_.=.A\_]&gMC^#_,INDgCd#P-ZAe[Ef+9O7/+6;58U[WI/:Q0JGHB3
3=?.GAOE3\(eF&DbH:.G/:Qe7OGO0#1R7Yb/Y-.;=?;cZ^<ZRU=ARa]C\e/:P[DA
R#0a#-B#/T:-BJ>-X.NSMe:+(GHag1G[TWB\c\H(WFQSb?AP)KY(XM<&@HPYQJ&2
,1]d:M33/K/fU4NIF)_N\,=^,;5\8-ZWXaPSaRcV\_MEH1MQH0Pf6g4?S3GgMDd:
1,_KN-QHC11M.@+Tdf02CXDgZ&[,_LR@1^Y(\Q=T#\9^+;X>UKF.A\^H<TB_<51L
O,fWV@ARU.5UW)Z59CPbYeG7S_2Ga_F6W?6f;+9Ccf^eb7Re82M@>ZK9g,HV^]#F
#+_&<P9EJY/P<7b\URb6S>J0[_[TgLY85/-(9XD3;.]0=NeI/V&5>7T>-.f?S[)B
(,caD)Ed@ZC->\EKX:agMZ)fcT1V0.T_KOS:T=MR;b-+=_Z?NDWDffM?AS]@(]e6
(c(ROG15P44(LTQ?8]:F#_4\I?D9C&Y>S5J49\dLY?HGdEAO]BD8041c_HFa_8]<
4f9GH3b-0Y.:MWCdSWgWc&V9=I6UABe^EgMBdWY@&J/04]ag&_EYcIeKYOMM+.R@
SLC@9UJaW?c3WK6+PA@ED6&BFM_:c-1B,XUUcg6:cKD@Ua)c.aO4/LXY7CIbY3:\
^-D9RgdTP5LaEW[FHG.cNGH^#b0T/aO:Q^10VM+66H_GB[7ML,0-8O_7a:.NZ,)e
eL[aO8>&/3]LZPAEc98?N)J@WFP:3f2IN;b6C3K85P&e;ST4RBH79^1IV7AeM.;8
II4XN]O[?X+c71H0cIPN3MX6#XV^S,f?9gO.TG\I7;\[Q.TLNe,HATaLOQG&C@J=
Z07JR-H.CCabRgS228DCJJKNE@9Hf+J9=,75((8eJ_:PECEF)[3JK^CBZL.9efeB
1K>7,I^0G>NOK;F_2O)fNTKJCF[\4Y^7DE#6a29#g6.^DAX+[,(c=SR>gM5H5G2a
([(E1d,Jb#QW/OQ.\=ZfD4[G(5ZX#V<(.@2??H(aH&XA_6]HSedP8>1Ic#GI:]BQ
[4KC_\_CEHIQYYWNX2>^ZJ;]F9d<-&&]Df_U\^BgfB7HaFd?-40U4=FKRBF.PMEa
TP7&RUA]6bR&Q[+O?2U8d5M>d<I;A\65+3V1X)/PWH&V,BFO#07#57>MdSK#A?OX
KLfU39JL+E_6,FTP>4db+M7270&>VdK]_<;G3S=bAD_PFE)_Fg7Kc.1L++&<9H_2
:8gLB-Pa2R\EgMNK&?#SN#;47>IZLPA.ga3\OKJ_TWWd>?5V-^ZPdfK<V4?R3Of0
3OgKCI3XRd/BZe+U0W..B^9ET2JG-O8cP,P_O.UJ3Ve[H)V,6AYI@S;2MB=#8Se]
4STXR>HX;CP6C5cQP^)1KQL:I4M-(#JbfFdCaP[2GLTDKWMTUBd#K_\K_O4g8XY2
E4NQ,QUS0gMJ?Bg=]OgRO5D&R<AX^f:I2X1Q1fce.8&7(_V^@&7f]>Jb8Ke5\G8T
N-ddQcM=.@7eW3a\b)>B:;3&\(U-J#Y73XAWU41[LTe\dMLOD,Y#TQ8IQa>Q>J;K
>B#.&?0&<PQ?]^<7>&cI(d,0BN45R=AgA8U=#7NfY\DbWg&NW+3XH8P1F.S:XZAN
1_5G@:0X969SI#)c.B>@XI_9ZSZ<I-),=TUgLK-I1ZBHABc(V\884\A]F1OUN:<]
Vg(<L9WVST/64UZ@DY<(/a^N=L[U??/DXV3CR@X0ZRP1/#IWI)=\5)2)6)=OC[+H
F4,V5ARH0AVM3(89Zee:g9CG=:7YE<V&,)JV:0<0/J9JHcKG26gd9FCdM4ME6.7_
\LFSAKL\IWRF9CN@0eAd4cDK_XfGKB#W.<>T[ZW8b-,#Y)-IKCSK74=AMA\L^Ka<
-B3W/2<H4XR[D^UW(/QV90-)<O<D^?fA[D2[^K:G@P@HL5])H,beG)FY:>CR.;?=
=H83/a.+AVf.&+S1aV,0:PZ,d3_VP#0<@X,T1SH<Z4gdgXH@QQ;FIZYLM57X__=Z
>e&38K[JeT^-X-VE7Gb&LKM4P-?QE>9aEb,ES>ZBd:^gM5R617<:1/BWS+(M=:GZ
?3Q?[^D_0gR7d2=@V?[KU<e?,P;DEa8+gGHOOS;>,HV3K=BSI5_b^V#OOV#:L,++
WCDJ1KP/9[O<Z^_M4g)H>N_(E@:R5XaB8JD.&T<e^E?1]aYX#63(4ZY_OE0-3C\,
28(5VSWY4gZa\(XPGVBK[4=CD[EH:M]J4JCC+E.4<g<gg:A669,6NE^J3SX[;WdS
5[D0;a-?5IVEDZLL,,#)gT6WJ?)#=7P#C5dL+d5])X#&@G35IcKG/D9PFf@?XebA
fJFUUHOGf:9XO>(:BR0\AU1ZaYaGE4>T_-:d&X(U+/be+fI4GA(A?86Q(D[-?.9b
N;71YI@cZ;^1_g>O=X^4E(VdEad2gOB;ccS5;<DC;3+9)gd.M4eZ:\EW)RSW1UY3
)f]LRTf^2&35WKRJd<DQ@]NXPIO_F9TE/1a(e(=+26BT_<4#cfINaMARBf_YQD.1
D9=1ae2NbeYeW#V^N+IKMdaK_cU=S\AT\f8CT\46RRc7J+.6F;+7U.7GUXa)U:+a
1+_6Aa\#d)=AWF+NE/W)8AQ152BQ(M7Na:LJIR7_+_#J7&c:3^0bQRH,.RSVV6)g
4(]6f#aI)Y)@:YMY;bY)bIH;3.9fa;?0baD\\34^<H?>QNJHY+[BMbBgUV&W&R3g
SfJJRQ#fQWMH&MFNV>JGb5Hc02PVCB0R-M[GDPQ5V&CYN7H88P/?Zbg0TV]=MJ(\
Lf58;8,F^5GZ=[4.A7)a^Z5NYc;e0V<LP4a^a^4H8?8gKY_.V4QZ9_/J8&@L>IEg
\bZe[J3P&g2+7,IR0F4->-<0[D29XC4;7d[6UALfc)Y.Q>&-?^bDE04E_:8CTfNV
f5_=RVO.^5X9:.#CS?WP^7_><J8O9e6a=g+#QLX\fFR^5/HB028G8[I;4QgZ\90N
BH,g\]B7Z(dde?PZF2ePQdAb@</<-L^9>F,LbU/2\?:4&_V9G9-AQeB5];Ob7TS7
,/=X;K9M:Z]0#\b,/XPL\E9,TL(1c>/_/fPB[Z,QY,@4f_NOTH(Q<fL[QMdbdbSE
:_9\C0I<5Y:QMW&\5&=^D:,[)00>.]A]F>L=JTEfY>_W7cY/&-dDHF8J:+@4Ta(K
]D7QK]bUe[E9PNEU<cQ5Y<e7>b5R&?[6ecK@bG=-bL[8LKJM9d\[.bgE?9E7bBeA
#UY#MH\<c9RC,R8L8E9<Gd5P.GDUQ6(:[@cWdG@)&A5-:15=UBLR>T5_GBEIE9>K
M0YPU(4=8-5=aX,dN-6gTJX<cbgc2eEU_E]2^ac-_[OY#N:agY<f>Lf9F9acT:R#
&\^4^c8ZH8aUe0&8&^,,H7F)WYN7AHFaZ6)TSHJ@(g^N8,81.66RC>A#N#+#O7R6
2ZP+MdObcddVX)?Z(/PC=^g9RO=H&884\SBS)LH@T2YY+S,11L(5]J1X]>3EMVIA
:4MCT6MZ#VK,ANbQ/=R3/RA@>GgLXTDg+HcMS)(NA^Y-CdB9G-\b>D6E\c;bXO+U
/\b6+b15+<P<+=6Ed[YNV#D?#3>)DX;(\OQJcI\285^:R]Bd27:IQK?AB))@F7NF
6B^c(CA-YQ_\8AUQ=C3,(>.@/XBE\:D&7MGX7Vd,a(PRK<:LS3c#4:NH>E;Z]CEG
bT,PC<VNZa-+\IHB2/+RC2c4IC:=,&6R(faD^c_ZU2DWZR[g;(16+V=CZ3.F&&&5
8,=983VFM4H.I7NX<D9P88^9/392ZE4Ga2g).576]^?22[=]Z=XL6GJC\[e3+\fY
^POETSVV/Q=gbaSa562#Q,E0Vb#aKN(:(e#Q?OJ4b^b#93Y;7)K+>A\YCP3gd[J1
T3)Z:/XDJ=?HLFX966(H[X-T^Jf&b6J^]WIW_W1JfJBUY#0fAfdKfb[dgF\#5aXG
RE.&UE2(J\O@60-X[Y]CUXG&H(/f5=M5J^>L94?K7^\CU)8<egcT(6bSO(N]-WR,
I(?F49fMMc34,a1&>gJM=caAWgE5TL>GQAY1SNg,a9V:=?ff_BBAZW36E-&QN)e1
Jaf,LZc.A#A]8=@@<&RJcD1[TgI9ZB@+e;994b)fMV0>??-cZ0NeWVMOT]-Qc<a6
ORCY4b<Z_@@1NBN)A<_O<[W?U9+_<,gdPR4R,O]TU12B37TSE<MJL]MF:\(=Y?(D
g7RH[-3J]DBbL-QKP1Y>KNe6TOY-g3N]W:VWb15ZL(&I[GHB?-R?Ae-Nf/9c5[1+
GBb_#(MTg.OY#M)4Q-?.9Z42b9S79D30UBAf5_:_fP-U?DE47GQ:XIe^gZ]09DPB
3b;]G5:Z/@9O@GP0C[,>0e\4HfR-)_4NU/ZC0L@;FA6KcbY1M)Z=B5/:U28]LKNY
_B-1JfZWU1c25b(I1,T9X>^#X=:geE,1DX1^=T-U7)?4<ac3CD;:(,eQMHgO#EMU
/R7C9e8c/bRGKOP&d3,[.[;XX5V=bQ/7+[WELIFQ/>T5>X1>Q?b55c0Jc/,44fR.
Ze4B>&F#2,[+cTNK,9?D;ADD]]^K^b:I?5;MBT/OP76Z,JWYE/5dF3OD/+=dG=1P
D+E5cOU<JfWE]JY\\-;?6SY13@]_HI#f9HJ?=d\,a+//A8Y]7<AYN3FJc+N@3fQS
Kg&XSb=4A.^4;WMaUX#9Q3Q-J_Y6-D3P7>VXUR87R2_>HPWf#=g(1Ga3Ug(_H[f8
)J/77UPeU#SV4O].J,OJESR4S6/68.7U4g2]YJ:79c_caNdNMR3H,LXf1g9+FP7B
@W][,@98PP/M<VA(8A^CVSLCHDc&<WOaJ8A<d:04&E<Q&QNX^bAQW/5K[.bUL07L
BJ=:gAH5:0:Q8a]eDA9D4^#V.#BBUE-Gb:K/Ieaba2Gg5fL]7c-dEX9_Lf3TfUK3
D9b80VObc2];<<?Cb=M>Ka.-ZL7R=^VIK.0+L/EQ.aWHR@W2-XN?M3D(++0[7);?
?M>_)6],0G=5Y8Z8R>a8]Ib=#AIUbW&a&G&g/aZX^gTfYeAZ8DRB5=VW92SUD<O)
#5((2?[fRZSEAcWeD[L-^Y?YN#_RD1(WY<GKQMd5<C:c5b/H.MX66^1NfPQ>M:0A
:ZUM\c7fME>P?1=425eL;@2bYW+P\b&AE-0+C7^SJ8eCI:6YP+EI8=808\NcA=?K
efL,TXaUfNJXEF3.PAN;C4RdQ>+.FZ4H84T0)HMQ&d2gId.H\;.V=E>019PU21E]
HVG0g-2ZA_e62,KEP=,3-L.;-@XVD6>?;?+@a68)Rd1/;DK:I<\)(_GSe5<^1E<F
@ERFXZ&[GGH-RS<J#HgB9Y9K8Y4TLCR6R[2F/;,1+E][cL51T,4A)dN,CW(B+d\/
\?aQ^C(0FMUC.TVS2X#6:@g=3EfM[?;T2b961&G6[aYdcQF[]J#-#<d3gEIfC9g/
\ZD>2B;=.GUQ[(A^2Z9@6L.0=cKa\8#6L:,TQ84Ib@MU;)H9_517[Y<&Y@B8Kc>J
Z+b<KCWY0J?c69D+^)NSE2G8)V5MT&:#GNVM@=\U-a,OZ[/>S82IVf)Q9d2e\7Nf
=^6NEaWQP#?M4fX9,O;F?+XgMYGD.A)7Q6Pf7#J3a<UTfDV(,^)GdY=f^?O:G;-Z
0_R^?bU2Q]-+DfZV.:)f:[dD##>cQ?YZ@(6?9Z07FeG,Mb:KX]-cT?NLACL/a5ZC
IY#\PG+[>6)CF^[R>RWYF>#b:E<LLKZWF6;;J.e9VZ12?_=;-LA9Z)G7_5Q^-\Pb
X..4,9[3S1RPJGB^?97L].4\g1cDG-&Y6SO77O)a+=L^?0)HgE7C-0#I>N:PMWC9
a@4L-/_Zg(@.OECJ<;2->^JSbLbL/QK4;;IV2=JC;-WE^I+^V(:T^,SI1+,L,8W^
K>#<8:5++S26g&RPXNMA/OKfLRC>d3EP-O2bQaS-OXETP)TZE&DMP5RfT]2SSX5Y
MW@T54C/d9=K0M@aSA/(P6AW]8AC:GIX^MO@YKE&@e.\1JTS5C.XS]BBe8#]d\)K
Y&dKY13G.g5Y((DU9@0MV;DPU0S5BdM1<T?<DabQ@-gdVMV]62g^fL.ULF^Re&>H
UC9>F,.RB<=S?;UQJ<cW#N&2H#_fJ4Zf52;KL554>7?SH-NTLJcR/Ia\=Sd=#QHF
BY,,a5g4=JJQ,@]FdY<W-E+B;@EPSQ-TfSHFZ5P8(;<,)5BDRSO^Z>8L3]+cgd,-
H<a1#4b+UbHL\@O7TL;0D@P@[aQ^PCSFG4#3V:0ZV9KLZKE)NU@<-84FRCZ6>>gV
9TW9]L.d(P4f2,FC_]eC8W>=DfF:EX]1aFSV8]<;F(.D/W[GR-EV.>I?_Y=3XJeV
)K>SC@:>L9\XP^9BJ30aN/<)650HRA<)CR.5(Nf978a]#W-f0G>cL0O[,-LX)^2T
SA0DbL0d&RF838FR;#H0D^6DMN>TY5d#?B>a;d\V_UJ>4W\SM@MC&_d4HW@):915
#Y+CAF,Gf7YfgXeA\aRV18.N7N=RYRZNG:c1fA2##GHM6C1W)FDf6:74G\14F)6.
-6,>)SY.U\,TUM(&AgX9E?>ZUAM^RFSBI@1QY2-b.,,M59I=4CLDD7L9Aa_3>#+?
0c@O3Ddb[UPOD65^E4I?UJ9GXS#UASZP+T&N[5Rb&1QQ22000Yd2Y[)BUdSSJ5+)
[9[5.>^]6RdM9,^Y+?F38Y32cUa@8OA9XOQD1JfUS-==>+Q:ZB).\_WNRTR?UQfg
61T5V..f?=aF&S9&b>SLT9A0=Y<TbdCeK:7?4K1+F=.V(\=;16HCIe/EaLHZgf7;
4=FN>29O#PLNWe35Fe5/JD7BLA2ba=PTAY<E>?Y^[)+MRIX+.[DHUJ/^3Ua?)9S[
Sg-Q1SW)JQU:#bT<N2N^>15V:W/ZPR:2e[W,S+BGO2HAKI^HeQ&?ZB@M&&_+M(T]
-,ED=6JU#)I;&@(g2(1JO1GRSF[@^A:CG6,C9WP,56?Y<&V.:B3X_J\4=_(.E6J:
/12?b@Af1G:36)WUH>?Tg)=,UCRGI_I)F_8XV.&Ob0U^]WbSJ9N3g3Q8LN)-&:;[
(+7V]=QNS>ccg>G/4RR#?P+BGP=4.HJ]=AP4.G6E?7++.85a/cTNcc>SQUDX-39_
?)2DRS&\6JAaY+417OB9F_KGDN1>M91@FIMA56>bOfW>&09-,&PDNcf:V^\@>J.(
e?8b^4+?=2FeMEAG5L&IfC#N.OAK]Da/Q@L60GS<f.gDF)##E\-&81SZ<2fb]I>T
N;SOH#61J3M[:]QH-.EQ,-G@A8dG390#DS&H9^OW@U3T\?,PLF\+:@N;M9VR>F^@
><DeWZ:TKP/a>ZCWMTW]SZ__>E#[IbYRMTAZa)7,4AgPW<XLHW6W98BV<MgD<Ac(
Q3;4<BR-7PU6E]8\[>WM<@&,Kcfgda:#3MXK#)P8?B).:/WA>2E_.J>W6>cfRFQ@
<.b1L_K5c/SD>.1,:2(508B,&871FVV3JO9PGKRUW>-^;Df5O(+L^_S(Z[3O]U-C
I]+1e8^7:Y3XLEe[/@38gTCbJQZO=I:=J70XH6_?PX.[:/E+;,?[M-;V4@51bG2E
VUT#MVX\JZ?+@.BHN62a-6<cO-.0(e=UU[RLHeXeb@g>2QMdBg#0>>3SQMI;-f+/
L?OR>D_]G<0[]G;W5?3WJML5K=&1B))^=6_/XN/AN@g0+bRA8KRQecS0/K.>9(SO
SaBHXcAcS#:TY5g@cS8#>92Je=@E.fX3R_X+?cATe1#?T]TMQ[IKJKS,\8RM7IJP
N^:EOF=JPfcX;C>=HAFbafT6dX85)0=&EB&:6f-.11=?CP84C3&1>+G.+5@#cM4F
>--@5da8Z2>@=Y9=\c<2N3(aX-RBLAU@B=+]O,f7J3/D8(e>V[QD@?+?]@#S,,<6
6G9C&g=R+]Aef@Zf[ITF5dE<d3da9GGY/SC_,I\HGKPBeVI<&[LTgCO1<[ME=L:N
11Z#a;0[)3[(&ZS,LDQ#b6>ZK63gVAVDX#-015Y^H/d8dG]/LH7/E#7)L@X8gJ9P
YMX6KBUf6GJT-V1[.1_MgNP)W9beXTac=U.H30MT#(L3>bIc,FJZAW[M<]FG6DB3
K5.@SNbAKLV0=93B;SPcUd_#H_C])f?@7CB+?16f4>1-/E>Fa6I(e>XZ_d[.#IK&
f<bJ=+AgE_D<4\M1/VW>7d-gXG0Z01AZ;YbQ^)Tf67BP-GAO-Z6c_#9LY)>d]^13
cJ#U(fLb1C<d#]\(2)PZI8+Jd=L@2714eUAIeQP/&<F9d9g\KgQeLFXHQUY\#LNK
)U6RR7W6Pe8#d7AXB]W\7F2/U8b]eLW3Q[/UdMf6eGE&7PLbC3gWYI4LK<U2eBe7
FGIOVZbR(Xd<&K5+^4\@9A]_>/@DA8cSfM1/J8^X_1fA,K\/-4X6^Yb.P;BcC;3[
64#(9/:0GdNE^b9e.F\L_gMZa1)UPKHb3<24g/<5+9XP<2G.geL,Z5X-3+4QFT,2
Gf/WS]7SbOO3:1;/GZ9^72_T\L2Y@gfL/<2K.T6P1OJ56?3M?W?@fEEdX\S=_1SX
HaadHH5&CK:LD6\+L0^+7^7;fDQLM]0;E7;-(=,b+&)J>]=/.]W1.ZTCaKZ&bgG/
:2@V^,Y4.?MW0I[17ZZD><04M@.IX_3aX;[LI(DX\)]b=0@eI.N.+FT<<8@9KOQL
B0bW@<VgH966.[]:9?\)b\:00=KgGJKWF3A]aaI:8^e?=TYS84DFbP09+#K,WIQV
e0[,@:Z&gT[[_+MD_e6U;e+,@GfbbVV?G:WPJ,;3-/D4a3ZGIJ0Y_^KM-))@7@d.
^g7[_9E?CcU0-L,9;a[Sf2gb1J8Z:8T7N)-S^bIN&S7=#@\-MC5\@L@W>ER&RO],
)?bP<ce[NN[35DVE/ZYCOTK.@0GQYZ=X5?O;-9ea/Q+Y-O7Y:-S#c8HNPH_5.(UB
dZP)_O8VfV\f-BfNS>LA<f34RE3g,OAe<Y=[558L)97QZ&+U>)aL0G45TRTB@A3-
_c/C=da3)I\@H]2;G+8IW,c#=-GOX?fK9a6Y\#KL5T@c#OK.9;QGLY/6EeFKK5[O
JUB0-Ja7DVf#5\4g4\J#6-BJXI2;S4b,<(d->>^N6ZWLfM^b:1TfddASOT3KY2UJ
.G(MG\43,d3<[-QgZ2:KB+ML7b=ISU_>-1662TSg\<fE/,Ge[.N]O?G,Cac0M@BV
::NF5O4L.3g53G=43_8BL7T/]N1M6OIDDGf4?R72aXE#U2GVVSCEJ&,M)0P35\:H
=C=4E\F13\VBD40gc)6G]J=_V<2)ID]CBc(B1>TQd0gL@[J(aF:c;GeW>ZPg<;d1
KX:S0>IZT-e@bY7Q>1:O&gLX[S:?(4NDdSI4/FOMNU@ZZC)RHNd(4Y]DObTWJ:R5
T_W(XI/HEe4K:/7]R4)?U3e^#;RU>4^8EMVE^:+>O(;g+K]EYR.=(aH1\7P20K;7
eP@B>P.,cF[P2R]3J>]Xc7f;GV63MC2aQd&F2Y^=Q2<><@F>&RX7\(FT_VgK@Y\Y
@\3^9K@#&/_fe5U_R.T5_MPUB#R8-P7XU;,OT&dQR^8,[UUfKI9+EDaY]9DQC+Y/
5RU>&GYQ(JNZ,-O^CC9M9+BQJB/4^aF;8/>bBfdV?.8],gX9@@5<ETF(QHOPGQWN
H1/:>gL<+HYPCOQE\J&Ca.U;7J95cOWQ\Z9YJ(aZV:)]UM)M7\1a?bMT8a;Lc?)/
Q1\-XFF[fdWdZC5:^-EWU>ADNHEQX>ScO[V^G&Q5MC8MJIPJOB)bY94MR(G]P;;3
=Y58GNY-?BRRTS.AN=GP@BB(Bg,Y7R?RZaQ#8beC:K&=e:fC4817=E#Y=2Ha,760
WEWL9T^eP_:0DaFH5PIWNJXg.f#8?-cB8WNVUN#eZYC:bP?:]16AcIFT^9#Nf[9U
?a^Kdfd6@-Z/[#./[-4DLD50GCNW_U);,/fDd-_=N]KdL)MD@T,OES0-]<DB88KL
ECS&bZ&O^)T<^+FIR<0(gBaV@/PZ?<AQcRJ:&P_a.05CLXfI=B1JO0_VUQQT#<#A
Hd:4O(6d3)B<0fAdMF2241E/WNN-cN\S?Ca3>\SZ^6TNBT:;L,UE71S0>7aV0HD:
1Ide13g/=W[KJ+AJGS[:)@]dI)WWV&B3<OLBLA_3F)W-aR2WTX2F6ZL(ECG-Wd2=
1aNJ6b3]UZ2TBA]\@>MOHPGaEXRC(UQLDI?PF_=5.^eM7UDKBC2.\X)0N#S]+67H
&8D^I/S<@RgO[=6ZRHQK[.5eI#(@c,TH&OfVBaf3<7-7]bGVVFC<8^]+;;SLFJ;I
]LY,P+20HIRL_A^W.bDdI_LKWbD(NY_CN3O5?S)-T-3UEa:?#R(/:OOGab[RP61B
VR+A5cdN-\W=8/8TJ0.MFZ700GY1,gMUN+\2<+R4AP^=1Q&V:5GD.4/6Y@SRHfFH
.)\.[^,&d/-Da91[a(<C8/1)P9QJ/20\24_KTM1+XZ=WLI_5RU)PBJMJ;7:82BZD
#cXR@Y+=fRJc/?^1B/#[=a:ELX(VJ5V-Y9.f_I(a210;6OT+Tc(5:;aEg<KbTMQF
/T@3FWH/]=J.7EY.cSR7HgW:DXP;7dQVaE99>S(B6O\>:X]?7WJc-g:\88Z[NSdZ
.)_VPH@<PS@9704RUDdSFd1L/JNZO^2&2N0X+1FN]PB<?1<H/0[Z4^c;F/KQSP5O
b2H(.:LB]8+Vg#EW-U:?Ca,TA93\\0P11;Y:P0>DHPQcZ(S6E-F5.(?)NP-g?^8U
QgdUFfd^f5.-Q7(R3e;&LC7:J1OLbc_T_OBC_7C3Hc@T;_a:UFP@A+7>P^4>V@Y6
f;-&W\88+FEZ-V(W;G<)eM\^;=cZga[MM.S,E2;=#D_@C^DAVSV>^=aSN8+#F_+;
-^W138C+a>CZ?]fA?,.+&#SNH9[R?&X(YASN1aYWW;BL9=;XN\B-+\_SgP0M,;VW
SC?5I\-&3J(U@O<1F.a2UR),JV9(eD2S1W>PZ#&L=SPXZ+E0/SKA+>2f2R-bSV]F
/84WcRLSdDYfaVC4g,\(Y.G]@g.-)=KEUNG,KR\25A1W5dIJJU0?+&.e\]+S>4E3
WV[0TK6L[MA)HAf<@aMA\#&Jb(DNVL^ZgV0KY5\88U0\Nf^-1+F48=X7<ZPH6(=0
337D=I\c2R37MdH5B>/a6-,],RSATaQ/7\;/DI#AXecVb0ZG]P2<RD3(4fK4-V;N
\C_cQcI?DQ6&:[+K0K?BEdBg.;)7;[.5,A2_FQ.F>O4LIa#7cJKCP+b#_D#f9C;g
?f#&;8DMODJcU;[L-4#ZZIAbW;W>I0ZD6,RgacA?L(JZW5PT-<1B[8CS+ZO(?c38
>3PF^QMeP+Z28d):6>PbA>B=(-S-ODSB8]\Z,aD=#@,<<[-:#<,Z+((M=41G\(7E
;&^(1,U&EPX943=H(Mf5@AQV@:#3R5MTe9_d2)TSeM2YZ]NZ+Z&1:7OWCQK;D7OK
LfS+b-8(1S#a[N,MNGb#94R@_#GRa?PY)/RT;OAW,ec8Q^aC_^7<U780c^XEgYQ,
#]LP9:+b]Ze-WP/cI1f]47?Zb[FF9EJRRLA5/,S)ce9X@^;=(5>4LJ=U>;=H^47e
VdY0gP<KO^>f)PdgC+E/]RY&8UAZU=c6IA:BJI_20(@a6Z1cU[+12-4XRTI49gK1
FL-2_I7\4+P5b11(@D>JG:UMf^f:)&dPc(-e(gOBc-&S>b9,PFG<Q>#8T7_N35_G
12cE;_bBI/S2XdSF[bUL0#g@)SYB@/)G>RC5<LCaX33UL;:)?CJZEZ3PC-A+Q?W/
]XJ9H9M@&Z>I6_e2][H<ZU[FecO9ZSGMU-C&.bCf])#&I>ILX.H9YTB@FY/\g#Ma
.MfTb^C2Q@2H6NC]f:cBDP(L[3F#G(,6/^<FCF5^;_GN7T4/.4DN[OP:,3B9I.?R
#LTbM.dMP6K[5?+S1\=(]<&d&?EeX>&.c,CaPCSa-gJATHHSW-[LWK-.c8<Y03=>
fB7<1GcP=7Z8G\4ff+aHTV9Y@G7;PNEW)@Bc>BW=4NOLg([MS?W?:/53QFJ&=I,:
<]Z71G5WDa:I8.f@@.T(&d7E2\GQ&93W)#T?[eF&V27^c_?UPDU1]J]&1<_>_1GX
AX5GH7FWJTV?\dKNCHIMT7\80>eS8RW&QT3ac\]5.R/^6bN/7\7[/1-472Q6H#XF
3S6[YK:[.U8c#2G#6@;fR&1OTG[_4b]MLK#1YdUF@4U;18F0ge.BRAf?H)1EZ?WJ
TeLIAa=#9U]Ya?MdS>E]R,0_LeU;2EF,WAI99)(_/,#^70Ee&ZGA5Q<LbR+B3#A_
AbRV8#<KS:IgTH;I<=/\;5;:6D:MXaGB1.ICPR3MCJQMNUY6)gbE/Rd?^FeZC2Ag
_]JId6@G#aOCBH]3S#2;gX8g2G0AANPSL]gaV+#^>ePA+-P>8C,g:O_-e(?X5]d6
0Oab-?ODRBTD38a_/-8QaeW0fP4S?_Xf#NY+GPWD>/CD3^/3T6a)gP+PR44H.,Zg
[?\abJ2^?90C]T,9gUYOM-]]M2fT.C=)TVeE:JGPMO/a(eLSGTS.<5bTO9PZJ<W8
#<_c3:XVM8PFXO]H[BZ;5_D+I=(Qa2G1BGPg1Z-41F6a2a4J.\bZ>E08K=S)].CA
_bF<5]0O05INGJgNaV@ef?J0TT]YB&Eg&_N1+g[ZeDZ4O;JJ2D-YcMb<S7;d+WZX
#:><J3VK(MO?1O8[QPd#<X)FZ3I#LgcTIDd+eDN7J8B+ZdEL4H0_^QE.@1[7Q[75
0[Z,^CO0(.7c<FW<OZDPPXIADQ&^JU,F((_#U/9JV_X;AM[LNLP?<F(R(1MSbSX4
6E;[S9e2LC-NEeTX,[#c/QW[(QVOJG=O7R(P0H<Z^f@g;A9E>+<Y(LR/5ICFL/5M
#K:4NS]VN,a85d.[D-?-6P?OPLS#:NcS3KTM-&d\=bE0]C=P(WSAAN77?FZL:+d-
3O9Je#:gJ-H22TR[JHAGOcQ+R61c=:fegI)7QL?95Y<:]-K4TL7eH?2V=;Ff?23U
b<<Q9:50;g:8OE,VSKBR)N4<7-OQH+_FF@O,e[7,K1M]Yf5K?WebOB5G[^WP\_12
1WO4F76?UQZ/P/PYO4IV)6Y1B[aMfGA#I?]\LBdU>\;0(H7[D<^H^;BK?7F4__.O
<f);F5Vd2]W6P(9[+@<;agV>G]4DVdQcRPY-Sf7.4#5b5;IV^MDPO8I;X>#H=LR5
2IF<_1A?\.VIQ[,YLPFb-+@XOIE#I6[.bOCfdUV@>FbbCd_ZMd9;dV]Dc)9&@0Q5
@-8C_J_L9[)U0G)=10TOGUZ1B&-@gbaNL(NS1EU-0^e/N8\#8O:I85(d0f-80>e:
N8.5Q3?HI_/>ZRR_1(++d+>X/ZEZ;LM,<fQX<4XLG)7;<;F@PEQ,1Q#F=T:3WC0U
HSZSc@J0ESPa7>aP)XQZ+\#@c=.<bUHLe;<&6YV0?YL&RV9KRN\TaRAbGWK[[J,O
g/KG#A6Z_OZgJL?4&g.e?=ZN^M[4T:U:7Zg#a7gV9[:HfJ@T:X;[aBXD0FP.VVO)
F&>Y3L<QL,;TC5<YP>GNZ/ID/UABV=)+a@?d.MKZ=Xa9geDfP)TECP7fG-EWC_R+
CK+7SN?\,6Rb=FUBFKg?Y&UIW[1RK@TA\O_efMY71Z_eI^W-=1[bA1Y;dUf;W/UO
8LE=\;0LGgO+g0YOCa)L&(24c]^,\:T-4YWDZX#3^[6UTXVUOUg(BbgZY4gGZ,W)
JGb0CHL#Dg6(Q^G]C^=@FC)2P(BE:T@<@1K2]+d-E9ADQDI\f/b3G4^2:fZeE_(D
-)4.BFa;8;;)C0:2?#8>WK&RJAg]-?P>^NR+FRWVP?DOZ+[;O><<&eLTF8P,]YPV
9&6:8YD1Eg2E7X,GPWKRZ\60N]5Dg7.93B&,MN83BT#b:TMLI=V=D&(4AAF[;3QN
XeV?OH]b))g4J@#&EKYR[#+cAJ_c\Oc)1_6-IQ&.RLQO4Jd]Z>#1Y)_V6d0&B.&@
1[/EWXVOb)R<,J[)Sd2]QF=7B:6E]00Q1&I6JR;4:8f(5B&A=/&gJXWGd&2KWd;=
>=/O@;S1(?:Q,H3HN]Fb>5JIJ<(L&3S5)<a@1KWH4Ua.Y>ZX=gL67TT+bX7gC7)U
N[EUJacAf6@f5&5L#c3d81\]5XJ,5BD&XeWORDAVFN2YT5:f0F\[Q,40IUA@#8M=
(AUW=f?&05>T)T.UL+<[_YOBd,.<-Ha=721[UQIe(b6@GF6[H+Y#QWV2f)U>1_c(
8cH;Ld=SdS;ONQ?#;U[6=eUdG+,1Q(0F>U,d.fMMXTg]-gP@f/.cT^Y7+UJ7_OF&
,7K)I8Ef.KDE,VdH<]&8aT9c^\baVD^(cbF23/OGX#7F#:Q64e5,EbgQ(2=;@288
V;K^3/?R,)FDJ>g)89aa39KegKYgT5#L+=WPWS[B>/&)^F31<P=O+3)V-3G0RC_E
B?-8UD3#48)-g?/?VY,[[98?22SPIDT]69PTg:I,_5I8A)b^XD##7R4dD>Z_/bFH
RM/CGYP[P,H]J@2G688+XdO6Q5IKb1];K?<a<1Lg.J\F;#O@16\PWT.;0H/,FfDM
H48X&I4@7=II5Y(7R8d-D,ZDd2@cN.Y9ZJV:><@3C5-;gOfO&EFg+f38]Pb+fHSb
GM=W?g[Kda6:6.OGd0A;K4[[9J[WaEa2LfWQLKB+HG09.72-6Z7I<PQC@Z;-C_dJ
A85-BQ/CSP.2N<=<QZ^>R3+WCZ6@4N1Xg(Sd]bVfU&(&5<H^\Eg]L\UL3&0aZL,1
:EP](_.DIP2LHF1DC<.];/S))5LEY\SYU-2YcZRP8e=U;b8/XX(E/5XUafbQ594J
<Y9dSgG[N42+XZ/Da->AU4+STKKa&.IE2_H?#)WD=L/#G9IUQ3ZefWEL?Y1Y_BTP
fCK&7\CI9^]TYDO7\-&@6>JEI2aPY3,E&<O]OGAUAJOe?K9RK&1Ob@Ob66e0g5_F
9QS].-+K@8KM;3WM_\/O>QWZWgKc<<XgC=Zb/FBZX0HF_+]Yg5d9PcBGC=URW@O8
JH4^XA#@@a1TOc#>f=We4?c2JKWBEZFf<(\LPG@13+>:TJ.7>RY1X,d[G:JV29aQ
UB5<P1RC9g.)P5@:I\=gd69F(+=+aAK=0dFF(Pa73Z?cV>-He#<-O0>4]bVe30H0
4+RSUBLFA4@c/=#_RG_#P868/\LPX_?MI-R:ODHgR&&95RJ-Y63PF/>gRA=,P14E
9<45NKVaZ-#-0(97Q8B>TX618.KRG3cWfYNG,<7EAU;-(dO961Ga3Q?6MQ114cSK
#8A7S(EG9@A=Jc6f<\##Re50=M6_#9Lb4X,1YH6M&G0/M<da-ZIT7LA8SKd)UG:N
OF20&H@Bc4B_+W&Ag>[=844:_#N2GG450NLUGLRd?D^5_.A/^DU?M9(.#[(f=^Me
a3#bRW6CF(WE[gA-6-GRaBa;8[;C?T#?\G0\GB-GZ3GfIQe66^B@F#2>;,(?A5e:
]QB9DI^cg+cdd6\>:OJ\Q:1R2?Id6a+c\d#A4EDHUF\OP-&N90=@TD-Z;Gb1d,3@
?&Q&=_)T:<4b:6[-@JIAeRSC=Y-(\#H(4a.754KKG]f0GAC+>D+3&51#D@cCP31,
/ZP;H6PeVa=^-b\&cab43J<J(+FY16M2gdXM)-?.O@fWD39MHU.5YeX?DGN/2@8:
TBNc^J+(7E+^XP6a/#UB-8.egfTPI0?^6\L,g)/_GA]M\3_0JJ6]a+Nc:7Q+a(/W
3c+Z:UBVGTHcU,8JPg+R^NVG&SS;\7?BYfCOY7Q7a2_ac;U3FBMY5N63=MOe^GBM
)]G@Od2N/;daGGZ;)+AfIBZ0?4#ZWK[C4@\_-/4&&a68/aE:?.RSH;><4Qb;\0F;
7S6B@YD=27[;7O4J(H[-S\CUa&(O]6D35HN@HAL]ATb4+AEI3RFRb&bX1P_@f8Z_
d\\+ED/PD>LBO4#ZQE]Q(4N)#\517;X1O77S\a7gE1F&&ZeBE^,b1Q1C;+73\;XD
Z&g6\<TeAQXF+3TfGdb7[4^I;=/67VIKc,Gg,O(RY3:d[.F[e9Afg1;?P_J:O2_4
;8=GB/Vd])T:..3LRgZ0<9?H0NRPb<@H^4J3TY9\92W45JE&1Q&02H.[RMWG2WL;
9f9P+UEUC>(FeU:A(W-J/Z7>07N7#aA--@)7,bgg?;1Ab.46/;Y.R;Ta<RQG-/d,
Dd>^\f@6;aVZd)e,C=Rd,HP5V/&^DWHgV)85f/0f/aW:aK78,aRIH(EdZK-08ZQb
;]ZL9X^fOBfO5-Z^M_+GP\IS5;MYPD.QN7/Ge>e;^1F&Ra5^c1/+@E]IE;O+A?-R
HOLTBF8B:]Y;Y#,\b6R2D9+c.Cd78F1>6eQI->XR]M8]V2E5_2I.]+2>O2+dZ9HF
9>5K2cT^bL7<)A>;00_:R?)E+MRN\VQ9+95G^@,N@?8Z:b^ee0,G^-#UN2Ag:E>B
I7G3=/5&[@@d(,M^Eb8K.eJ8H?N<>>8RdGa=4ab4X[^FQ.:KU[1:H0J\)U:IE;L;
(R,O(<W/.WYIGZSS6:EQ?a=3H00#aXJG981/EHX+QCZbcUegS540#O3X+Yd#5F9^
6X@RQLf-LNRU,XAMQac6-=H+=/>H=S4:G5+B7V4J?#=?UZ&>W5>9JdLO06I/Z^;;
\f8\_T-P[MbY>g^ELA-LQY1_4]]LeO]H=-THUMFKUF5Q\O24W_S),+,3WS/;@FQ@
EcJ<D7H;F;=d,-HHBf\=@fF.^E0f#QcfS+b4\eSP8,gBd9\EK94/_JXb,LYCe.03
):DO&S<d9(5_X<7D&?gCb4:&I;KMA\AA7L.VGXI(G//<(KA.<.5<dN?DG\b7V:7+
6A<GS]d76\+[O4W18S.B7-Z?.EBI0UJXYG^c<(bLC9MWJ-Qb,)M-?@ZXPY^97b,H
FB:]aFFNS0-F_5I)ag)BPVN6.K\7f02&1(^7:4OW?9P2T>U<CK^d?LOZD<9bOIcd
5^AF=5/]g[[RgMBX4a@8A1>E74AgcgXgA:L/AISA><IU1Z/@>e1+I-5gRCeTT@[G
78\^gSCb):9:Xb,.-LSU8JfE^JQ=CT?Ee[FA87B5F0\4Sd4/N>X8Ue^a_fS2-ba>
HO\);BP.JD?SU2L@353=AddB=Y=]C06<e)?2Sd<LBNCPJ>Y:L\:RPC:.(I:F;J6[
Q:g=ICA3Ke9dY7W7F;g==YcL9C@?7,JWXD=[:O7<gW3X?dYQde/=[XK4>,TdX+&B
<F5Af_&K:gWQ5.^,)HRXRYgM?W-M3)532&I/f6UO^Cd26.bG&BOT4P30K6-JP1f6
<K22#6/VT4#84_E;g(AA/&6U[WX4#gUEK\+^C@)B1JYZ[b(TBU<V&QGYHfWG)QF.
PNIFB:4<6V=D\G9^a@\EATdR#Y;_]0W83H_=3dY1eFBe+4J:09@S]7Qe>geHM1&^
E3--24;7KQV=Y,J?&B6;P(C>N;VU7DcQ5:+J>[Wed32]5<\dGcBK;TF>KOND.ZK4
+Yg27EPF,>WER)]8IB6\g9?,XBd,^(KWQY3aT4DSRNdP<PSgHD<8FeQ?e8aYaA7^
5V_2&Ua@9(-UF.;>68P1MKD8@cdd:VOV&_cDb.RSPUV^5KZ8bPVN95=-7\V(8Q+]
6.<BR:V<6;4?fVEYC4I6dPA/J6Hd]eWSC(8HADg<I@?_XbZ.D+)NX&[.aU^=G\.[
D&ZQObH.JJWdH/N71D+J9M3GaP:;K9#?/#G::#^5/g^PK;H4.0bK-H+?(d4DMZ)/
X]Y/TJX;N+bN?T58LO22aQ8(TB[66><aRS9f)M^-3@d&]]ZgM&6LV?b;,SXDUBc0
_>6ZeE<7+@8DW5DFNKgS)9G<-)b:c:-a0aTMNKL:F9dbVUMe6-3LH/Ce,I\7\EcH
@fO[23:b9+.A:U>^/X/Y/S92@Q/4;,Z4aJHZc4U;./7WXY/IF7FMW?MY<Qa)\g\=
VHb2+\\4/M>H4YAgSY0A2/LMQ0XCMOZ5,CUc/A,=]#N4].S/b0SaH([)a<F8ZFQ1
+W3:[P@YMGH#>eTOB0PHD7^UTB5,SB(W<Mg1JDQ[5gNN,B:OX&J+\?VISVZWK5E_
ZL6B4X\?_;/2\ZSM/;Vc\N#IHGAU7PTE;FA5AH;V][YD28TBU^ea-&bNQ<5U5ef-
SS3_e\]K/0)9I-+-E^P.KT)cVL0RN1-2+P\Ed2W27e)V5J?-05-Qe]H]A#13EK,=
7?W=D1.VF&P8-/M^>CSd_)\aH3X2Z0=<+DZ2\YUaFfb494K3J_=(b95+6##:aQQJ
<@K1+e&.eZ[L<=8ORS?<GdT_@f^g09\>8P0]<P_0eY.&[\H06GH56-3ZcYPNW&12
:K2,W)?OSSN\&Uc+@/O2#.,#8]PG;5/IDVNS)N5J;,bD.??+RgBS(6\DLTe,DHa5
SI5SdD#B>Y=(.X0\L)9ENZ.8;1@>/([PU^\9SR4HQ4Ng4C0VCa6e<.7M,HBgG798
B(<((<__Ma]Cg.C/##TH(0;]bBB68?+/JO?[Kfa6bOaMU=59a[)&?Zb)32QN=C,b
P\FcZBMEg]2CGQO--Zd923W.:5WgR@I=SKd82T\:J1:]@A.<[(P[^3R<:4W8PINV
OMM93O1<Y)fN)3&RH:7cI48ZBg3(1CfH^+f;0I#,@?-I2P8/f/.5P9TZL;^.bf^9
_Q^EVMJQ8][7-7d?TU7(XbL28380>g<YJ(S5]>?:F3BAAg([B1#?ObW_<dFgFV6J
PAXOI3Mefb\Q&F31,@V@L+Z71I5@bHDC(EA(KWPYeX>@aO5^L,UT,FF&IKcKW0b3
]b8A@&4\aXRWJ3J7TJ4^[KC8L=XZ1:N5+C1aQ7S9+A/.cdUAX9YHE1>+HQ.EL/#4
]?+IBTgRcZc+9RWFabM?=:H[:(.GZD(59,Z[CSa1U6R[9K1Kg=P8GU)UH0_OU6I:
X060PU3]_S[-U77==)T6CK##J54DDQ=cB3F.#MeWO8Q\@0DAU6#])O]Yg@F:XWL@
WA5S(,g[4MZ<[(\g3D\&WD.J<&L-)M8<HM:Mg8DaP\bgFLUVQM38e@<:_5&&/F9<
3/KHTS+C&\Eb>5bCO(<FE2J9W.EOT=:HTD6P53Ma:dB\4^LM,3TL[1Q,;KL4UG@&
@,NdF^W.81aGZ]0T^WI</<I>6+>gP7NZ\[cH<F4CEG4?\6eT25/QafMSVEaJ[a0b
19??Q\=L#[#=]?)G=9?A+bBM9)2IC&&6SZIRK)[-9-F1Kd#\e-@a;:C>Q>:MDA2d
.^G/5KGVT]I6dTGacH>9;_R,6=6^Pa7+,J>FJ3:CE\)7PW;MZ//F1AYGC)^(#E:#
fKVG=2,d_G(LYdB5RL6NE9GbSFX6M.)d?G.Y7FX7R\A:,)P+Z4R+#U:&]QLeaD18
X+BFP>3?MSZW.b\S2b).^BM3]+HSB9B]L1CgE+E+)Ce.-GaZ1Q52O,AVb#&D+B[b
O\c::3QU##Ug\6/.V]1EAaUY2]&Q_e-XM1>_CZb7+K<Yc97cC9[CaVgS?SFCU;/X
(S-ffcaYV:QPUV35\NCEZRF08_RHNg2L\g-)=cbJO[D^_;4QIa>EMcQUG=#+43&9
N2aIXX.dWH9.0OZ_S^8TLHc,BWa,#EOEEB^AMITQ]9a6bGC:F7gS04W,,1XM^D5U
)>G(:VTbUdgJ(;69BO\G0dAN&OM(72:IZB,;19K?TbWNW_YOXcHDY)1[/T7Ae=G;
94[8FAgE>)KR]\-g2:\=,X5;+_W0:5H#WHdgGH?QaBO@]+Y,\<:>F^6W=&72-@U.
#=MJ.EK6;7TE//Xb7NcI8daEF(N,aON<CFa)00Z#G[>LOWC(>),.5#,K#AYZ^])8
S16cC#U-eA1.b6/JT,R:NAC,O8N2_43NDKJM<U-1Q[&83S^?VJM3LL.IAE;1CG9D
-D1K929I5ag#gQ,#[D=e0b5e>V_L\MH):IA(280/T9X5,P3J4XE;f\DEdD\W+)#f
0/)6?_V?3G6=JXZ^7P7J;g6Sb6+<P:cJC=+,=ZE]g@V7\H&SRgFgK0XA#U,HN@BD
,86aNCJfYEaCd;V?g7XQC.W[ZA-BTGc4S#R]7+HdY&H@XK;USA@.P]]#TO2eU+A\
QU8VLHJ9W1G_#+>)QfY0I_WR-0[&R.#0AQaS]fME1X7(KU])beE+VM\cBDf93VH5
/1Sd09EN&c.-.3@S@fA6CV^^-B[\aT[V0[F-5\]B[4QJgb]>J,bg2&SL<1R;)R]P
&<0RMM9.aCC.CP;(W,&;G7>FJ/66<-K.QWK5+<>M3+);)@=4.LN:d_U,K0EYZ7Y(
ZD=@IS(X)dB(/#KYZT[CPH=#g1&TV>e/HN+?Y;[3K4d9/8#F#ZDAd>T6d8U6Q@CN
Sg8SW)b2^+<E_5I.^>)J6PaBX3]R^eG:OcfC<FX(3G;WI\bR/W6)a_TFc<GSKF5:
\OV38;HCgUWK8cTGWcG]5NI?#=\,7M(BYCT3>@3F=<9=PT=_S^Q5D57J/8R.9HLF
?1E<+=>@OEC0f2G-)V,YD\9=EX6fYC<P_XDK2)0W3^:JE3ZKfJfg\5=65Wa1W3B]
P-VGJe;L\[eW3a/L4D4N->-;HQX29[eeBXM4>X\8LG2G:31_3;Pb3U5FPR[e>Z./
.P..O^-3/e.AX2?2IU45C<4GYcS[9;8F02(8g0O;gf\AMPM1R&V#bXa]X14+5CG)
FJ@f)_0JQ#[\^MB7:+@O3SC#@7#)3dSC;?@-9+D7gEDKRRXG5Za[VE.HLdUa#9OI
(?:HURTfD:(OHB8&6AS<eB+Q<:D0YXY]M@_58HedKWaeH15>N6IJ_+S]O6ad,7H]
)G\+>,H7;YJ12C@8Qc,L(J.0[_7=@0UbC_<[8;Wg9P(O/H@YY)[];R],?XC225O9
G^][eYD9)PS4OLR?9CY?9(P&KALYQ>;f.0DI?=N)<(ebW-22//XXWTTH;I,.A[&:
OPY.^G]@8A]\50gYd\=Z-AJ+1=gNGZXH[P66P>:4CWO2C8>,/TEX\IN/R?BdSS8]
Z+,?TcRaPR@IcELUX\Q>3aUG2+8ILROIVf/QY:X;,^/)S&cA<TP@:UWX(6)ZBNVa
cI#Qb3ND-)[9)^X)AA[[\.Q+,\2\[Eg5N5-bR,7>&O)UY4A,b\DA[gL[bI,B0[A>
OG;DDT:@=;YDHD=LQgJ.ARP/bP[faA=7-Q+0S#;IR8)5]]I-,^aQ?8R.]W+G4<.(
(K<O<S>QFK:KAfTe@B:cEQZBF?RAIZ_P1\9T[;16Z#VX-S^QIJ635&8Q5L(ZH_\W
V<R4(3RU8dJ,GY)1Hc]OF:JBVP-1bC9?AJ##AE1,b]C6(-WK:Ab]0bGccW[_2IWF
ILf#0=UaG:TQ3NRd1(?gRER&86;8#8]#F5EgW025&cb6I&1NG9&_PB^9?I[P;GbP
HJ6Y/&IQ1KVAX?dDUH\PH]F-=?2>BENSf1bCX/90OA=_Q3DHMW4XS_/F36,54\1_
D^B+HQ]A7-1RbFS;-MQ9HPLd]BPH(CBZ\bDF+.E?>ZJ34+IIO\?9G/@_MQJ+c#]a
D<2<a?+KYf=e1AHa7+/I3&WBUJX4FC\IXUDe6_Sfdb#A1J7c=^R+&W5U[;[PV96)
SPBFP/XDUDV>I(11?\5FC4c6RC#KOMfCLRS(e/H#MIg3AKgTW3HS2=?gX5_O,eW>
4,X>LYP\+3V:=YTA+G0L7=OZC3b[5V8C@157J2]1,PW@cGA<,4L26BW8-FS[_Y#L
YO?3bQO2(ITAWb3AB9I>O7cS7?PE^G[[f14+3Vb4V+ccG.IP-e0XLaQ-JUIF[V]M
@\)^a_PH:a0Ceb/8.(#-/;>NU1_T379TTCZHff60\g,YHfOJG6Gd3Z5]@gM7Wagd
#Ca_C^.GY6BPIHQ#@^9/FfC2AHGC2gc=4NU4CA^eg.&PY6a5I1.DPeM(#TD;3S;@
]BHf2_1PV0gd=cPC7(D,K3^5Rf.](SKgJf)e6H+.=UH(NL]])@:2R^DZ-SW+F]DZ
gJUA7a2?eU,(R_XG#H5f#,.^_?I:gV)2<TTCYI;P3UT3ZN7XL_7ZO=f6BNDLK)bZ
4E^4MF86P2=(;>JBFXbGE9KDFG.gQY-4KeC+dQ4fSY-f1dWe-\TYPQ,J-,:;3I6J
#8ZY-ddM+g<[F/U3FCDM-fREgV7R2<Y\J#2&g48ZaCa,(##)L,>1e@-+;4=8K:9B
/JUge<L6&LDEAUc2CQ2WGgPME?+@CGI:)0>,>I)H^S3d0B?DKW;C:CGeB(M;U9&[
MU\O+?0F_<63H8,F)H7RQL988:bPf&PQeB5Z<^gIgd<-ER/Q2)\5<YTBQB[E\SPb
Q9a1)U^J7TgRM5@E0CI0(\3.O(#g1JQ,_CI,9:=#:ZD+1RY(B6,d-Q.eg,?)[@Gf
X#H@<YG;0;C2QVEIA2V?)61?67_2U@3\];<bF3Q:L&0Q8S-\YXAU@OIEP]A8X+6S
M2(A>3MaK=<9a\^e\C\M2_JHfPSZ]LN12G<O_F@XcTJ^?cZC@?c>H]EK+)64Rc^P
RB,9CFOEKZ<D<Mff-<J11>+J=M?3b[W,22V<#K3?/YI]8S3J^QLKVe6Ag4e2>>,0
K&3.87cdHV-MOFYeS&QF?VC6SAf42K#B=.PO8T13HG=+eLRZTfXaC]F3OU(P2Q..
&5@Dag;86B7@QYgTL6HKF9&XL)G]QUC&W\E>9K3.Y+=;41B/4.@>BF?+?a@0e0TX
JI]9<Uf\DWN&]O-D7Qa=::7eMI&e25aDMDAUPLb+LUXCYac^6/,2L^ITJKFUV=\b
C/TZaC#3XfKf89UX,g(&G&PbN>0(KB4=EZIWM7,.07U82+e6MY\a:2T41a=I:a&>
<DBQ&B[gNJ2.3.U[]H5@X;^=_21F1ZacZGDUOPW[M/1.b.=J)IRdWPX#VC_/6a(b
DNHK=3XBMFSBd,NI?V0dYD?RR)1C(aS\J-:c]BOBZ_P(JgE7AOBJb]8f(HLQ^C<O
5EF;+^E]FW\WW\^-,^_+;I3&O^1W<Ud-49Z;?G_&\/4BH=L80dDFTU?.EJC-(5Se
@IZ\RG(QUB[6<ST)J=T?GO3N5ScFg<:Z:Nf=I[#afT?0RVe)RNf6;8+,2IE6:-0R
_>-LA\A:3Y16e_7P0[EZ@7[510:5OAfHG=MWR)R54EP,.#5(&TM\^f/]a(KLgXWX
]C8EcQVE9.=)TZCCS+;BHN)dPC\PYG_(YR.7046ZNVA3O1R.a\]>.BV1?N?07LOT
eGH\Q:6VR5660dKLC12H&IJM6[[\C/&/3]2M1IbaTdgV@GcZ8Z,LEa=a/;Y.DI)W
UBDJba)57\@>@3KYV1B;7a)@K#4#^eB.OW69a5V6/<cdO-VM_1QA/bH/&01<S=-;
P,Y+9V:I^F@5XBQKYbDeMcCVR4=9-6;T7[7QYdeMM,<Z[cDQb4Q,Xa>M#L+RQBUD
XP?Pgc0Ra\g-gKRR9N-ce)2_a6M<CG@P+/T:OL\:e=T90GQJMDWFWCM@MMe0Bcg8
A4/==BY6Y=7W]2D(X8g:S:6<-&7b;[\S8.dP_SLEL._AK0^EV?H7D?YgaN-4D/Y\
.5P[T)GJ]WE^;bZ[SY7=NKRESEd=(3fe[VSf=:8<V3NMM[SA=/06Z<XU[4C.6_#6
82=B_3VO53S-J8>YI0fM(dfY)cUQ/C3Ge]I9_L.]ILB@3b0+T(f#HN0fNFP8<<g+
9?g6CN]SR8MX6WBF&GV[0]0HO5ZG)T<\0DbVT@#Y]LRgB:-cI_-LCME9>LJ2Yg&Z
Z>d#&gYDS7_FU(59)Q#cd/ef<DK,AJD-TbOQa9Z)2-L-cD.:NeS;IVHSQc5-QDB.
J\7H^FUeNJ8XORT=>=>]-TX<[&eD&4)A:ZFIYT6323c_\V8W6VJ+cC<eH.\FW80/
CL?(-I#]X(<LH]CI<c64^W:2D:#@MbdC#Zf]BTdg8H.54N]5<CA,JB\7Q6IC/+0K
P:M1&ZGD?2f;=aMD?\6;Dc3UQ?b]&EWT8,\(A)N>P+E_8<X]G(F)0IeP6AHXTW8^
3_4NH,I9E(9)3=5Sb+c7SJLMc;0JX/eK#Y:8OQL0=Cc9)UD#Q;RH^@PcB>^8]R#N
>K8NKG(7ZQ&ELEa??.@EW@_+WS\ED:=#R:(3I?7KWUT9^PKDR+VE)eWKHPFWC?JK
P9])<AOfLBZ<9S^:77db_,;f\,9KBg^A]_4I1f?c9]8OFYdW:7]#RX>7>@<NWDgX
g#>bS77YBE]590R_]_9f]4]G]Q+?3,fJ8e&CeQ\(93MV,Z0]e<3P#YGe]_M>([SF
CE8-Af0#5<E;:TYI,XSN0<fS8KQ&T],J#,cPN>35S6^\9eDCGJ8.[.f6c8ZS&>,>
<.5Seb^fYfXCM7UD4MZW_Y?8R3-TX;G/B01&[b:06OZKXWBX4MdYC\JU&SN3HO62
+dd-5<KU)ZfNK[.&MJ?Ig&>D)L73d:,R/E0]dAZUgGELB3P]/G:cbZ:fGXEb\G/^
<)dg5>&9;(MdN7GU<+C;[/-MC-<1(67\U[aYNIH_][]+YgGB2H&Z]/K5Y?-Nd(g-
EV\LL\VM,1GA?N:fUM=HMdc_XE2aDD<<(K_KNB\P@Z8d)_=g.5fMcP>HC\JGOfW[
5O^ZIcB[+ag@DP<D5D\.Q2a?R+b49<FP;B11TMPPJDbLD?H5B/C>=I(^@R)4SXW(
,,PA2I6:UE9@OFE2\Cba&LaN)2=::K4QIZfaD?1,QTa>DT3R2f4;Bd16JdAfRZPN
]#e=7D.@1NI7D6-D:^.f?[.>RadKX2H:Z00f:L;1F0TLCd8=BAK(e9^+CBW6O/-:
N_J)T?/=0SZWa3D_gJD)09(1gHQBWHTN^O./5e^,2MJ>+,0XScSSH64YQ3UVaZQA
YHH17I1E0/X:PJ-/&aHV(J6c>HSAYW6OOOWD\F)JGJaA94fAR9R\=<<cH+9c7XS,
(DDcTZ_9,Qf_[=2c\)A71DU#M60#eT/Q5KeS];8WW#8J\,1K5#4T3<e^+.gL<d]=
MVUAU[]T.U)\3M-Vc5IGV148F+-QE>SVT8<:g00JfU#R[UNfQ]#f@WWGLN<GUPCa
=4OF>?^^=:[7]\g42LKOLNZHdedR,DID#N#7.<DH[^-T6:/cO.f-0WP)+VMP/C3c
CN5U?)3Kb<V)53GF^&VQHTT(XLKbXL#>7_(\(g.,1+EAZF,[TI8U2NM;[VC<G=Da
IADO?Eeb[SFDO0Wg[PaW?G_OQd]E3ANEQ?.:&Y=b5CE_E6D>&KXL_eI<0D\8]/K\
aTFcC3&F3VHB:c1</eYHE-d,-KVNb42HI0)LgF8DgV^P6-YS(db4Pc8KN2?3/0V2
/>g?Z[,((1G)@#/-BgJVA#DW(4AN/CbXPde]W&PQ5Z?P+7J32986#J3b;Dd4DEJF
RRYWg_T[/<.ff?7LXF.Y&;)3MIX?]S5dN#P5HgE)]JHB6(Hd1&?0cU0QG89D&O3D
U6D6P:&JNg^e>1\b7XP]AL<7T,KJHJ<eK(-WDRN^7IgTTNQ]HK;d;,CAgRETWXFE
U@a;+.\]c&IgZHG49,+U]2<<@:J0.FLLXPgEZ2&^V7F1U5LM6Cc]WIIK=<S,;N5E
G+Q?\5bZUGdbXJR?LJOgaRffc^:g2WTTVE\eIg9->J<EMC9K5<B[MF7J38fM5F/B
S].dS]H=HdMB2MHY72,GX9b>8)\F/H5CgT6-HG]1?-ZBdNf</F:\\4fO4Fa<JGE-
eB3gMcRK[]Y.bE>ROVV7L;_,R0>bKW=^eK@_A)HeWQ\:FH7JCN>9TQgRG^#UF1O>
.77]J^2V[;5W<;7-&)(U\EcD7;ARVCKSFTT>L6\WcW>P1b],YV6ObYGT=,g=S[CR
IG1J^TdDfP=bE[RdQ+EG_^5DB>Y\SC#N>SL@[CgNd_CdRF3U-]4)ODY]?d^Ha0S>
7+O0YBb26W2S^T</X8>8SX7;X2?bA7Hg2T&@CbceQ#&,ZRLdH^F\,NI+T&KOAgIE
V@_5,.D))L=-6Td\d6WK>^d4Ke3A3[<=U#]<&;1A72LacedI8gNJL@L[d&==CL92
=],.-C84G4&3O,T8[)08^]a0<c[(7&SWLZA5;=-]=aCZ:[V2HeF[N#@M0G?\G3XV
4V,.9=T_DfOOaLVSIB@He^GL5J&RR=EOD^O2WU<bLJ@H;]A0P_:)TW[<WT63)MD4
UHe[0a?^f[NBZAS;4IR=@_E/P7C>7Y59fb(eZWO#C72g]L,-W<N:2>_a\[3TX;+9
=AKX&UcFRcN^WI(JcSCgDPP.ILNFWLBLH?B4QfKYY_QT:Wcg4L9gBZY-Z7;#?=:4
@Hd4fTO0F)C1BIeFWKcE3L;,D&3W<aKJSJBE#/8QceX(J;Z=Z(4@K^\7e_cdRUb^
g#Sc0g_R@IcGZ9OZ_2\CDPWX79(,QfUVI_KfUBL6Y,[BX@28Q<L^VL3C(BT\/EK2
LWP47S12dQ,.bVF-XDaY_#+@70XL[.dQb(9__K?TM.[D_\aV>HLG+CPP3b5U]N2/
G:8.]gQb:1+4F+^A(@B+A;Zg;@[DebJU]-6D_P<GK?Y\6_AQ)KDJ5/A1IEJd_F2H
Z40;G_I.)9Bf3AFfWJ<71e/G2Id_#.=/gYAF?9^]12ZQ+A^:]/E+_]:82<HIUC0P
f]dc#O,Oe6Q,e^dL;)^@a)B^;Y9_#A3.E^XdA:9WXcNDEK3?>FDF8KLe-<0(F,F@
T<1#RaOV)HEP.aD(df+1<;B#WQ).dF5^KJ(g/Oa9-+5KM&b5WWD,]1g6HAJf-+Q:
cM><,6cG^X=Ad7&1JNTDLPX,b:>g&W/QQ,(bKY2?0PR6e;@>QF6&f0aadE1Ie]0a
T/UY8A4#OM:-2LUWJ]K40Od(XbA]0:dV.4FeAA^PTG3;RE()4PXb<.fPa61=-47M
9&[/3\P>U>>:Feb4DL;)de1SdU<6c^HQ(@8<P79FYT@B5>cUb3g/6:?/E93#IH0Y
,HY2#J,Kf&Hd^F8b<4MN[[9g?9I.ZLd#9-Y\ObTLYB[3M)Cd6-_1aKAL#H?g-+d;
E&^,USIDC=R6#\L9e2R]HeaT]c]X7afCHWZE08-C_W<^Z?&S+_6HCCg?g.A8(@AJ
_A<@P3b,</M[g8/JYYUSF29d<>QLg_2DL2@D._<)R-2Y0+>7JO6dH5DT-H?-HH;D
;;>07HFA^X6)V<4Q5EZ/M4.,^&STaBB7f)\f43S\5(I-O=T_\OSU(<d?]641,;d8
E9=CJ7L\RZMHGbRbFNXM31_-)X=Z.Ne/?1?<:E2C-RQHXP#3bU3^7^3cJD[+XTF;
5)\6J6/WATU4M7aHX/,JJ^EdbCP;[K^?e]OB/DWbMLNI=TXAYg:PSH8e+8Bb6W3>
43[R_[d6eC+3WfaD0;/P(ZG(-/+Q?Q2g6=gcB#.9T[X4YC#Q=A1:9@ObA_c6_AJ2
Q[RB>R>J:1A8\2D+8]?<4C\1/S7@Og4_<A3K9]>C+=],WKLYLRN4PQV[[O+NUUEB
+b1d]Qa\BEQQ<^8R5)/+>dA[U>JC0WNIM<e\)9g#X?IKX-SBP_PN2AVLSaSPQXX@
Tea,IQg0H_F8OXg>M7c(G3OYPEKSR.M1fA7Sg5+Z@)d?TR]S(9LGK:Oe2cde(<gB
eECd21a/&ZgK5VL=Fae551JS^^;gGFYD/9X#/Ve5Dg\G-2L^7d5D36JC?TGV5O,\
94B6C=>@f+FPLO:+TLE\^d2AX+9B@RT4^I;\1#&_f)3JbK5N)S+43#_72(<7V@XY
FX8WXF51,SB024D>?Dc+Wf-/b@DfDS3L760-AYBJ5I0#C]EPdA^EMWV0:\IAG(I\
<<Z#2V5A)V584RdIKA=;86eKBU36@;S+]VF#?S/^8a);BP?)O@ZGK6P60VZf^XT?
]d++Qd0M]9XZK8<@^YeYLNM&<1L:^&ZcR[MHIH@dT\/4A2B,T43O.T0Q5+&C7+[I
=cgJE0K.eX.)H8eY=S>P3>AV]Sg-cbP[\^FO75\L4Ce;e;Y8GI(V:JZFU8HeVaBK
/;O?@5ZBeHJ4fMGS-Y-,Ag-;PPX;_ce=4?&BA=W=]GAK9T31J5LGL[[K]LCHbHP@
:,4&8ZdZURX.Rd5PB<A7RH<_HWC_DT0#I1c;5.YAV5BA-83W?/R>=2f_[64,HQ,&
\)&Z>aG;@[Y:M,Z(0ROV.=^<;B/Vc^L=7Y5]+eGMJPCC2;)UI3[;T:YB0Wc\@a@K
J6TUb?.M6YRPa,f,#&U5LYGH^3))fW;E?Kg0Tf?ZeX9HTa>UdCC2MAWfFU&@P@G1
9fgUN9_f[VML;HKS^(<&\Ke#LQ&A.U(+L.2I[UBL6:B[eOKT)6TfL2@-3N/VG96c
TD:_5[9-+cX&:O8SHOG?CTKFWVc]B0^S^]f5&68Hb)0fgS>9R9H25_[1<.1#]AWV
X;?aF>&T_I4.;_4AN,=Ag]+BW>_gO_P@BWLF+bC+4@G(JVfZYbfK][e]>_\c7I2#
1&Rb/f1[PQM(,_CUF7XY4(J6=?H_-L?gNM9/]V57R.)d>O\A5.EZ0.\ff1<(MaSO
-WK(42TI@.[_a9:IAe.CTf_^K6\H3FC1]5)g,cYV]E65X9+IOB3NQd#:UA];ZV)W
b[0+V>LIdeC,;T6PYOS0eNPY2&PBIUKF90^P_<,Q+YG=FTLCQ@71?G1,#G/0RAdS
:).<P>,9PbHH7e9TZ@31.).MGT/WH]b-KU\c)#I@fObHVU^X6PU:U=4.1&J-U^B^
(\LQ<a>C:1N4^9+,MWYbBPI>F)BQ^#H]IV1a&[X8COS[C7S.PGY>)T[;[1e/FWge
fc=PMdE>60ES1fb/I61]/^P3;Tb,S1EIXM,/(>3)PN]ZVS>FC#=eBaD?4V8f2HN8
U&fDa&U@(?Vg(#Z[b__PM]R(0R^Ug@_/\Q6TM&Mf,7OY._f#7F?-aN08fU0gVaFP
cT=I)7;32gH2d0CPCaLYE_<Na+?\&:ZZd^-]]Kg)4(Z0#=,EKQeKWT:0N@#@eT/\
3QF#33ZJ8N]_#DYT10JI2(],;bO95)F(1AH_FY4fH=a_.<>HPg&H;74F_dL&@&.4
M_;@LV@7V1G)UG75Y&H7(^Z\>==-Kd?)0bNBB1ZcO]5\Ycc9^TKPc^YC-V,:dU-\
+Id>P3E[acgYAd_CRJ@,V[[]d7.T,5>8.8BgE<bf;39ZHJLINC8ZT<?Od+&bWUBD
68HUIFS;aG1dcJW\GdBO:8c.<DH6GE7/_b.dFP?-:SA<2HQNPH?+S7@Z)LI#GACg
2(W:;]BYR5&\18K91UOAVb(5\_/gcaEZ@I#A3]W>NEV]W/&H9M6Cg./+5VS0_C3;
Z/B4:LL[MN@.KH^SGB&5bR+^dc.]DIS@O6?BH4U3=GAgS/P2+F\R[OX&L.2UNJKG
X5I+S3)Y8)[N#SS\(L@DOODE0YO6ID8T8fOfE92GRK18aM4A\NDQ(d_bY\TV=d7@
(,<#]b>+NVV5^:55WCg>SCS=O3X11/L[4E;MP.&cFE@:=-UdMQ&3/-7;I9H6G2@N
NOK,ZG@0cDYX27)SM#f(3H,9<eG0SIaH6NGVb]RXS+9=,H,\,)+96V4(+)EQ,:6>
\^2\]^PL>DQaJ/^E79cNGBI(BF.WH):O[OST2ZZcSS#VKHXN7J;)?^[5+F3eM;;e
+81=cb<G-T3(:g]Y2PF+8M\>aSGb_5>NDKQ]F^2#3A8/QQX=:e[Zb;=eJ?18#_Mf
/8YVdFIKA2NI8PLf(+GUTO0GP6[42KK#eOWMGJLLWIHVHf<J.SOa?WL3+368Nb.V
^I/WM@c_.PEGC8^F()_=_W2(U9GPY5WYgGHM85I<0R&DO?:#MH^g<O4/8a5=&De6
CIJ5F/JbbJK#.4B,QOaGB?;@],SEM6LU#LP7&9=OUdJ42:C[_B4KZ7IU0&77&)_G
<DR/)O@HY8(WOOJ9]e@\,Nc07#U-,L\T14M5)gH)0E[HS]d_>X[PY<(-5=>D37XH
[-#OffG(8EI]HZc3+#/\;2<SQ?.:G,:=aDMB-8H@L+g>1JN2I9[)@gV&,f&9W_&P
ROe<\F0I=5_S]#3eYfW9DOd/;;eOBIX8;##VZV?YWFX6&Tf7PL/^3QUQECf9?U[K
aHEA?7+2d&F=QU-7-gB+@O=U_/&3b-c7EWJdO+PR#c#D+5K#I7?P3KRTC2KMM))E
X]:L2]?A6P&93YOCcTID@@0Zb.S<A,\YOYf_@HLeX7X2d=_f]4A&2US,)AU^6;6,
fHH]J1+DNUUF)\b^SS(,Q<96:X;.A0C[/B:Hb<eM]Y5DT1TUgK9X?)1;Z-FJ>;-3
]1Z6L[9?&BYHP8^THVIfU+X=#\A<NJCZKO.9TRJV</gRLPW8La.AOSgJ,:OF<&>Y
LNYE01-&+#T_UZ?HWcB[.P61/Ld,OBY=X3T;WPH#S8<U=B,.I[&gAF,QX:6987N8
F+;FEI,E]BQ;BRK1ATHS[:P[Q,312L6)B1MC,GV+3;-Y;f9E.Z9+0@?J.1Ya:VVg
a9J9bdBFN391a[QDf55d2Z1AdV\LIDg<&>&fXC?Rb#[\LV_KQdAH-\O20gE9)&KJ
cfbFWNc]V(bBAZS\Y:B5P<_N,853<./XJf-9J<_3d8c@,V4B[4L>\]>JJ/;KP&?1
bQg_cCN,D\1UD.4b_3;LN0_ZYXA4590P1=@SCQ(SQ-X,cXU?SD^ZJ(>#^2QSdcE<
DG@),FdR6(:2b@9TKI(X\)Xe\FJ?<0\TOaf=T?<CR6W:O/F:T[4+QO(&(COS-(LL
QJT7fQ/#+6JF<)LK>=dGMPeE-UbT7K.RY^D7.7G8PR]IGeVgfAb;ec58UR1TKR]g
Ree=KA@;/Z/46EJNQ@gQU?[0W80c:)N^?Q_NTZ6^=5[,B_.X-._=>fBQ/]R\-;XL
DN1YFG0QU0Ke3@4Y<.eQ:<P,\PME(7bQ?XBJHeGKMR^4FJ7A[fCdT5a0f22S+O(f
D=6(AO7e7PHQTa\16T1S4fYGE)GSdZ2;437M[#;6698PWBC<7bFeF[WO#(F(daKH
74X1L[1eHa.YXAK]K+]BPN/(B#/c[fGa;<Z09G+dgD[acEGcWO8K2<M-ZJgG;70b
J6=CJJ-C]>ORcN^LeJ.RF,I&G@/4J&^=D=VX98[,9@\,4SCEONa6EWKB85LeRINZ
Y@@,dL@DJ3^(M(8SZB=,Q)1&VV_^K^@[75<9Y5NW_aOeZM&@b8^,FL;NdA,#fgQ3
b<(#N7,,Y448D.BRX6;ZeL[9EHJB<3cg:<Gb<@LGV/c;]?5(>O>YR48PW>4+_ee1
-IG5QX5_/XEKM:gdV;]N3W&?cWDe6G\E+FA;Kf_T03GbXeN6.VWM;gY,GG(U;_I(
I>-Tb)DC(aX+V[,KH6GWTLUXaJa<Q.T^=30KPK0<3Z+bR@F_?B7#f37FD10Z=beP
HP\,TG#LF>#BB(@)>?C2M)UeCT&>JII6fSE(,-?9e(b,YJAEF]3.#KISM]XKDHJ8
PEQ=YLZ\VKANYZM0NO5PbT5L7g[74^(^F>]gBB&V.BT;,)\LAc4/eaVVU6E+M]LN
BV5^+-EK3&XZVD18#cHM9TCZTHI6+L;[QK\eKJ5N+X=JTgS:d#L=V=C\UMVN;W(1
OO;N#-cc/9SGHK2&<V@K(B\HT(GM\,8a@-3K=e2Q^=KANfa257f5:RV,3<?AEEQf
?cXO&7,K]NcAOE77^=5PI=@Ib/M3\d,)-=@=T0U]BT\HUW=6IbL0.PO86UYfa+)W
X<#V5;KTfHC?ML0/>Z7.^F(.F\57#]W(?YZXdV9[J.V@aYREI(WYHJ-(WO>11=ON
W51^XcW+G..]?L3PQ:Z/;5Q1KY(9F:B8Y7eU5:&ON/[Qc+1/0a19a&=@7O/5]24X
FZ(BZYO_/CM)gD7-X/\V\cB1G9Sg,Y@7M]=b[FL?)DWK??fQ:=/77^Q8B=^6]C-)
N(M;QMZB,:TI15b-D>,7O@N7?;VY6Q>E=9_M=TfR)bBDDPf?#2/[Z.(X]\QC^ZNf
>(B#X?bAI8=D-][Rf:,,F6:fWL0Xf3aA/N3?7-2KSG>1c_K-_C=:Fa#:dRdgD(SU
ZIOI=3M,PH+J.;fCeR8\(JN@D;H-gQ&a@[C&4FMTE\?f^9aKU_Wc&BI[De.@d-F\
<XMO&<&/2a8bg3Z9&5)UPP+>6I4\_<@:bd#_UgbT#)dZ,EK[,O</a#WF,[Gf??>6
)ZC80L9J&32Q^1fMbU(D[N&TJ4Q)P=0)ZK\aI3IGc\QH&JJ+]<ZKI#W#KRWP6<0L
[\2L/AO1<M7BM(K;Z7,b00D+C?9aaA?a6-eCOJ,2IS(He[:7UJ9Z,gC;UXAOg^H2
_A-C:UKd_2B/TXVL:+LW(K8Q.(?::P94Q1S_6T>A;DFV>>RFAB54V836,6MORfe5
bEFOHTD@>LXeI3)7#E-&7LOLc,LRRf^1D:8edS6-:9L#C&JSb4H.X@f+-<KL.3BR
IFMCfb&&SA4Ja33EFHT#^(6dY([MEUWF,>EN[D\>TCK,G[9_S=U,/W1HKO<F=6]F
@PDPE;NM3.252G>HMf[C]V3S6eTU2BAQ9\4#W3ZO3Ea2?A=2VR\E:JJBLO:c=O/S
9#d1&\?YYP8M3[8SfJC\R;A/5]ZPS#Y^bN3g,5ENZ@1TB-eZ831F:/G)G#L,)afG
b<KINR;0NfMKNMD,@8L,@12AXQ;(EY]d+=V7IZYVW+X&&X^KAXPBd2[E<Og+A;UY
eW+I^MV6d[E/\T]G)0d^=HC@I/TC-7O]W)D#V>Nb+e]#NZJD&78fN>#TcEJ60204
I4/(f1S_^[I\-E49JTMgV_E,J?)ee,5@IV.YWGc:MUeKGF]]4e/VN#[&KZ[7&W/B
U,@QJ-&EOWV<KX0XffC58N]W27eWIe?EYQ#VY5dI+I5a18fd4fE;F;U>0X#AP+^>
W:gSC7J-KY(<K:Ff;[@Z1O?\:<(2JX/3d\eeg8(>WCb,+PV\S#cA\;Fa1KR&^6J^
D?EA-MX(QM)LMZ2#B/f[<=GI=^HCWbOE7RJW:K7HM,R)Q+ZR^67B1Q-J[7W25.6+
VZB0gS82R4KEDgaVJSK?bA;a8bLX?5>H4N9&d8\WH5_1Z&3775K9^>LS,e5gB7_b
HWOg8WP3UI39EFI;841b?Z44OdF?C,=9+CK>YE[HZ=()UX-A1_2a:fZGd6&3cQ>c
?:Sg>[PI.4(V8?aTNB(PKLc)QGKfUS?R2B5JSgg_7M#>10I9]/O0,H8O@&3=KA(M
TSEYF8^UT#@H:Ed6\JOOd?B.->I_4Cf-E(YO_8a.IQag(2\SLHGE.L1,M<D\+4(+
^Y:2.ZU)(X+&0]I,AT1RZH]\U>#GAQDGCD^2H9X829]YV9UWaY2+cBfc\]c8NK1f
3:KV9?G#YagPXKI0T&27[YA4T[Q531_A)_La(+/S\^2LAQ?8\IJ2T&01e.K>5?4_
KQ9@PYL;(DS<;0GT3QKdZ^[MW8EY0CdT=Jb/?b[\g)(aCUXD3#+I.YXf>._FWFd_
^[P0PQc.dL_EKeTQ?e#E)\0+//HG7e0Qb\4b\bYKfb.S@V/cf(Z@K<_fLfFL8:P[
PSM9Y(@]0dPXSbT@7L9afQ2,+3Gb9(TSOR=[_b:D]][8Vf5L?J(^(Q5-J:@<>a=.
\=/HG7[T+A(HDd;&aOW>GV8#QM+F1>UEdE:]QZA>Cg+H.3:BMJ+NR/<MM+^V\.S2
\6SBGH7EB,S&I]L.C4DG6Bb=aB.UW/b4DC)OLfH5V4LR651XV-dQR^8g=c2LgM#>
W.8TXD@EaXW3XD>(,.ZKWSD#aEgU8GBfa0]RJ^e1A6-\JS)ASP/aW>ZgcdIZ(+d0
-[[=CK6d@,5L.]F6L;[2GM6@EPYf6\ad5+\dcdW[R->D;=3]E?4281f6/I>A0X;f
AP[@6F-A_RY7P&FF6+[6DgJ&dV:C1G3].I5O20ZV4L,SYaYW@:SJU)8HP+SAOPY9
eLaBSDf&WX]P5R23&T=Z2Y6318f_HF\LJWV.dLOc2cDPTF<Q.:#&Le..>A(HcIGI
aH>W88aN,Wg(4IZCYG.B.80Xd1Q/M3(^JJY=FO\U:V#L@Bd^0Q=Z6N.TdE(,ZJ8(
O36=def(bP?KGV@CPZa.XQB::_ITIY@67VH,GEY]/^9>U(J/)E.),H/fJG-74P1_
+NT92Z-#/+>_0LHJPe=Lf3-IB8faO(&#;>BW[E>[<T+3):d^<H2(9V_ceG#I5@J\
(&:1<V?VL33#L7-^S005:dAH\,-&5YD_^689E^H46Y5e,<Nc<M_);(A_b)WTWHFF
aG;BKaZ+349V?F5S-&.Q^a^Y?NVBTU+WJ8TC(G),g:/^UJ).9fCc=P-X:#;3gFXB
J0UcYES#+V8Q3WaLJOPgW8dIKHeKOD:<5(B8/cPOOZ4MZc>_e]3V<Yb,G)[O\B=Q
E8:12+5=06TK9a[BcY#,6.0ZV6940/?#4RWUWL;8#UFa4Me=G06T>,^T^f<IMZ50
MQ=bC_);?Z(O3KM^US<U,geZbDA7P?T9.A9K>1GLW8.3S(W/cJ=1dO=J3g.X9GT6
2#cbI#_d9/-;QR&/A[6O2,dIZ4c-X46R+P)+4NK;UGBX^U])WHLd#FIP^QV5GRa<
S@&9,Q8DZR#PY/9Hg@TOI9N&Z[A()/>#^EWMdWCO4fgW,>C#OK?.87D?&Kb\e=#7
F=HR9X#MN[6GYOP;OW^Pb@7EV@BW=6PBFHJ/E5ab6c/6fUYXV.Ae,Xg?5YV9VK+R
a;WeC>VE72\YYB8E3(bR2Nbd3<^?SaD>NTN#Q:&ZH]4[8+8afeKNOCPf[^)_.[)b
@NdDc6SCUaGI,<(2_.Af<4&c=9EfYI)[MTTBa[5;NXD5<O;Ab^=d/H/?QF)++DUY
XbYaF/6:]BM\Gb0\fT/&PAQ?O\C2@5d4FdRT5]E&;8GAIMUXd(=.X7K]11DH_9Te
+MHSU]Je=/R:7.FfXBd5K^=OeS9,((NWA&BHd_&:?TYaOM5UHP7A6R-g@8-QKB9(
e1\2R-TXI(G9Ad#;OA;\AU;.ULF:G^M=ZgYcI]F)eG:,1A(;SVN,Q#;Saa=b@?Q;
-+W+3H(<-/]SNF.V6F;]];U#AKLCZ&.^[8@2MRJ-^#@.OEV<OV51:&=Vf3_,)7--
QU/Z_-EAfg_dg;SGOH6#.,L8UE8[g.&QMSg]\_Lf)7agI08QE&252ZU_?e#+Ga2G
cZAV3QaR0@DN.70#6[ON-PNOB4@_J[cfI)]\8WRTKGLRKc8+V8OIYQ8:TH+UWgK0
GaA?eJcXe4&c\EgRUKG-^N@RN+-EQ^;AKZO#,Z)@fO&]=.-_O]@;]7=G(=E/6L8[
E>2;9NL:^/^4c>Ug\F^14g6;2D8K[R)33:F;c2K5TYPDV2RLA216UQ,QW8IZec_M
ed\VS2-eC;41[e\8PBJW^(9;+VI1Rc\E]//6R\ZOKgPPB<<J6YTJ+aR2#:@Z27:f
AcSb(=_)1D\R[e3XZ/LKW28Z-A?9WMZ5DL)JU?L/BW^N:73ZN5P3c[;-:dFfR4@0
,18@c+BTVI8Ff\2T8cKSTUYUg_H0gT5;:>25;/bgVe31M#.c7bB+M@;3Z>ZLDce&
L3f^V1:CDRX5\YY?[QDH#e)R\Pd<VgTMB3X=]_H=LHc/=OdEY3=5VX<E#dA]<C1=
L8N^cbbEKFPYacMBF:_3SC)OJ0V\PaSRN=5MP.-U]b8#W4fHC:<SfZE,+Q@^KY.P
ZN22f4,.1I&I7<SJ>Z>[SX9:9FN<QZ?^M(]3aH;=f^&[6bfC-K^-RD/=JNB)0KLa
1O=M3\P3LZ)bg.I8aba48f?dEQK7X(eXR/P;#CDV#13Fd&Sb,-^U82B<D19T85+J
74gB@TdWQ)MIGTaHAP>M4T+)#Y4MK.[L,83)6T2L#]XeAXGD-cYfBL(>]+,HcQ^a
_;CT49NZPWY2)WCP]G-WQKcVPRe5/4@NY\L]gWWeKJcH+F#bB._@^9fB_&9geb(.
aEX8.QcPX/9C,M\c[c4.>UX_E>OQHES>\]g_VW&9+^fK16C&fJ<)3a:cGf.+9F0K
M8K,aNa-HKRbH8A2g[;92OX/^XYFL9Q?0C_&LMBgE8C^JZE?7N?PSf@1XMRB&6@Q
^HE)2\;R-fC[>YaS[W:-g/\]eBY7K-5ROUgcUW9J0g#^aPQ6?>P776&T=NGQId_M
QZ7bX@aMRAef2,(/DBfXe#@GC;0#<\=E>+YR+d60#7NLH-TP,.CBTHa(HRFCGHA6
TK;VPH_B#+IBbI2A2RXG\XeMXdQMPc#0aQ30),&V2R-,Q=?CM,d1B39ZM-([:^gE
7WGNR;3PYF-3+a&])/+_=Ga@D6BUD&<CdZ[99L8LM/K4IL@O^g:[FWHg_LA-=b25
:34D0d(&d6<.ZQZ:?FE+DAfY&EH7,4+S6BI2I3I0g2g@&G]6QR9L>b/[7f/LVb97
_M:U-=Z0TL:>)+=CL1D9)EQKNBA^ZA;JR-\)cN52]ST.+YWY1JE<#cSV53@/c3O,
94d5FV-K&L9-E@YVZ4UNVUQT4fW-KH#1SD6K\FDfU7SS1W<U1a]Jec1OHWRYI=-a
(MFDRBJMT/73,+c16C;@XO?A;6MSSTJ>D-TJALFcA)fYdD<K760]eE1=LUB8P,8,
Y+_7[36KV[JW_.g>_cgZ4^K3:I+BCb^BL1HP7_-cZL,X<34^61P#(/Ke^C/+gOI0
Nc>M=g-=XF]Q@G?WKU:F>N01+ga&I0CGI?26:,G(da1@>5e.>G15?T-8]+-;MS+;
C#^2ME(ELYbH)52g5OEK:XD5X8d<X)YS@1EIR=:/fXA1V0-WRD>N-;agg;-;LGA,
g\U/CeC1\@UWb(.UBfe+AaAf<F=AE&6dS3@])#_VUGSYZA98L=5eAc2+2&)P(\dV
^bf3RGb4DcE.5+=A78U,)&=]-N@Ng9HCcQTW>WMJ:Ab1J-HQBZMg2dB(0Id_-<A@
6&D_VgG-[;SV394&1f](9:ZA1CWCU/O8-XPd8B\QFN-<#)U>ZMaS?M;d_9@_KAa>
FHQ_Y9]]SBC6C8)AT<1f,BW0gL9222Z<8ZDFYIF\e>I0,JQQ1Te5B^446WIW(-=a
gJ[D<A+]^FSAH_>6DgGA..;E.Kg^&@KQ@QDPbJJBWgdQWHcfW<#7CMPF5LE&LO94
TM&,.f)9V]82Z_8^c@;N6G=aPK#^\FM[_ESX:Y.2S6I3\&cHOCWZHD)U+ISF;+C7
#]g[;F_AM6^1+U&\>4<,#Y:XbE[&4=^KB7dIG7e1F<4/</;R<;:]##bCgZbfABE5
\7C,7B(IK_Te&P=aE:@:Bf_V2cB8-V0_RB:M7&&I9;af)O,D>8OG70W7-\-3_O#H
Z9TWf0J^&EU?9N1?XLT+b)Bg8J]Q]U:>?Ib>P^&G=L0F;0@X97FE?e#D>H5CU=9V
WZ.g7e(Oad7U]gBOT6-,]OJL\OT4cff1V/8DD0Q+;<E.,,5LU&c-RgVfPV,>X3BM
(fJ+G4eU9)g:CGEeGL?>bLgKT02E[IS)R9_87L0GJ[d7I,AG:afb3e;;DO1B7V.7
[?:=7cNL.>ZOg:&1C4W5\BeEG7B29VDYW7_-9gEgX?[Q6C0a9Bb7,LX96GLO)c:Z
]CA\d5\9GH?L:T?0TRSgBL>S[9eg^:&_a#W(T@<AL/W8BI/UAg-)f,R2cY<I5-\1
^[;\/M4Ra:YCeDSOEP)Z]/^6gWQ)&4,&)U1]:DEE7)Y0E57<4DegOP-Y[BU=@\R,
e(Y^AQHWM_9S=?LaS?6S2.#Qca_:N_V4c:(U#OK:2-ScH[?P8Z+-e4AO(RE^9&AL
gdf/5=+[\BA4&,/6<A\5:/P6-Y2:H4@c2Ha).6a_IRL8Ne:@/<K/SQfgK9_]c:HV
48aS:]:9<I;]@3:TDRL-^aOPG,BaQbA=?c:0b,>T_aUJRPUVeC4gQ6XJ)Z.M=]eE
DM61-b&CN](=>(+I7deQ^,?SSH,NZ5+2EBP/^,&4N0^54XVQ)_/KKX<QV=#S=?T1
+W</0S;#>&F]XW-D^+2O8V]@TYC.,U5G>2T/;V_SN#eOPDT?&a>?ZL])&>9XJSCF
FSB[HA+W>&I/ISRYadIREb45BQF0(JCd1Rb9\@I4N[4L2I:MWWV=,=6g,]KdaN?:
gW9<13@Ed3)).X/9)8QTB9fU;>g;/#W?B8-c<QKWTaf@^4QS5@1cW=447]^R,AT=
D)eM49H-FDYN/>Ff)M43g)]-g&HL@4be\_.\a>JQ2a__3[FWND3S7])g/A@D(GRE
(K7G\TI&D#B;&Lf4ce>3B)a=10@.=D9Xa0TKfE@BDW-P4F]TU-TeYe/6@<I7NPCK
D,c0<JFNMWKY>JM)b?>aTNE8.KId233W^),T]LXLB&.(?#)(@&M+ZB<Z83I.H#=\
fG6X8/=>:B2S6V:T.D^B=[4_VbZ7DeIUHeE8YD(,^R9Y:NY\Y=S[[X?0,fBSA?6F
B=g#C<X>VKS4ECa]fE>#Ea#BGJ>2&b=<TU)SKDd8aPF-b[V^CP[a;e/>eX0cG5B5
>&O]ETK2^F2.8T5(?Q3V1SI5,M5[_O_fJ.da.E\D2+1WF[9S^U0BF/f.+LX<6(KF
XPF>_2g<6@[#OSOLW(Z/UIQ>YTJMY>g8[I9_<_6WK<A8#(AUQ2LNL3A.ZP6;[HeZ
,SZFg3YPZ17[2;O\B60G,(B8bF.d)eE&D]VG.KCMB\BQVJ+624aJ.]C38^+^@TG0
FG4Y9:EY4_5=)N?#W^YAbfaQT;S8NYDX:6e_gY7C8e7UVd8()[FU<;5dGT[(_&VK
]RSAdRQE5B+#TD?f_,<aHM?H8/[D-TVPA\BE[b3Db(N7#B,g?LYJ(UfM86H9]dR]
/XL8INQ^>NET@-BJ5D[G@Kd9Hc#.,B;-(,..DPbZ),,&4_W#2<c@15aF64(Z0,BJ
Dd^&[G^<;.dL3(_8dYBHJ@B;;DL+9OWcA)R@]NPFLI^+6P9O7+](D+[=@47@I)SM
>R>Oc#aIQ?^Pg7fAJRd#eLYK<=#ZB\GPQDF:74-e2;+Odb8KL5<5I(bIAf?>e<S/
9_0._VX2AGU^S_-a0==E75CIbKD7=:#WUS=&T]-\=)e^>U.@.>a@0@I36Ye7W]=>
39X@?/[HG:M=KRK(V4[U-[?W4aPO@ccbYS1J.+D4F<&66RfI/5da\65I9V+9S=]F
SfG/-1+=K&_FX:O\MHWPAC-b.WR5X@)DJ7X[aG??,N,eZ_->)eE)M\<RF-+-[V>^
8BG3f,-<L0;_\<&dC+;^Y_LY_d&aIUJcN.P&+H\+I^;S;J(=#SF)5B;;IKZG6\(O
.WI/49Dd?HM5PXP6^gcY8\RZMCfcI-FX.HN.W1K-3f<YX-\K0/7dLAYb7@24C2C0
R8g4Lc8N9:]Za:3[NCAB-P4OZ3-_I&U;23=/V:\&V4KU40b=C70<.EEMS)aTH#V2
:8:WILZ@83C/?JJKGB?T5/G+5cJK@EZVZ4LDBQ?#O\+^,T1-01<MEdDbROW#PGMS
Rc:Pb?;D-)e(=<S9@>Y1dZG3)>T<&+7R<c+SUKc7?(96Ze8OH)S27aWa67UAC,O&
f])b(HU85N^^XdQ?F>0)>6Y1,?TeTgD)d17A1Q3A;2N5dPd&NM<5[8[V^]=JWYZQ
9Pc3_79_3aP#6[._MEMFYDH/.QWLdf]JeYeU@U-LB.99J=.O]bC@X&U;K7[+J-Z0
Y9CP0;^SMYFL?AX6HMS3UL;&]71V/GP?g(QW;A(e+]GW3NRJ>YM<TPCG1Q#gWe@(
5C:O;4?\T8E8?@dSB>^8\,,>2[PPZg3?R3(/=,V[g2@]W7.Q,ZEWPL[-),UTScW5
KY(PRdPbAf96?Vbg>1Y7adN+AX2?VeJF1K_TR&)+.fO&gK\#cF30O).]N2L=f09U
a2aZ[;EVQODT6O>&/[J(7IWZ:aB&c5-DCZb:)f/(48KQMK3bI@&.LV5gRTL<A[>]
.2V-N+dC9OVgPO3.?G:_\AH@#8.#O45NH^:33\?U2H.#=c[2-I1&OD^?5-g041NJ
ab#9b2Z>#H<GO21FQV9PcE?W[1ZAS>D)HWdX4e?;W;<^IfZ#F<]JTX)5/6d2A7/6
-;_3=^JKP1g+:IKd>9.[Of_2EZ/W3:^7,^b:Ha_A]A/54BOB^?&2#R]XdC>?RdCe
S_>JP8Oa\HMR8D)P)7(;LYa(H0;0ZEe=[4CIP).1)2L9C;[I7#-Z<bV,IRJGY#C_
Y;,SU4-UMdEW+Z6fM4>9/QIDOLM9N;SD@&>?DX\OID@-D/&BORa2C/;ELRN5M\QM
=<;=b/_[#C58e5467^Q]?IdH\+YG<ILHTN&9Ca>ML#G9/--G0C+WDc3+/3T1YE]=
K/OK01e\BO#]D783NQDY&.:O9bB/AAeEe^_5VJANbPH0.9M4ZJEbWb]L/Ne]IMF&
//b6(0GZ]JNPAf/6-TU858?8_7VfQMW@g]L<XG4:e0OE3H:,c6#7JO#4U\f;3[JX
8)#)NR,ZF0=@ZNUYdEcS,L1ITU8\0G\83\69J)3Y]HZHWY]UUb=8=bPIXP^a7K&>
2[gX^@URV]E&fDZR4SD\CUg>IQFQ5A_c2-1_1VW@MH14Z\+K&P#d^6J8f4QUUC4D
dYS:D&Q9I?:Q:TLb#HDbB0_7--fS4E(a-JgPaJ.c/&=3W.\I&YE3V(MXL@_96Q6\
6fITEH3gK&9RLVDB5)WdBR/AddLB>?UIUE@O#)Wg#4NM6e_8J)&c>b2R(]R_H@O_
][<1=CI+:V-[Ra#-_aA0D\(V?:;]]JKgUH5.=WJ>_SAb83DaXR-758&&=XFXd1e\
5J;PdSFM,Z>>R\dEBe.d9;@U1,(VFVQ&^5P0_>6+eUEL?PY2>#CQa(C[2JS0=R-6
XLc0O#;C+MY.L_EdG0S^6NHUM&AF#dL&ZHL;;TZ]<fU&B4Z.aEEB3aTVG@IQPAB1
7MF#)QWE><?J7_;61;>9cXS)635YJTO)Vd=@ND-G-I=c[GA<-6O1cH;Na.=0BN]Z
eY?dW1f/dba+//K5I^CIa@JG<fgafEM/_0Q:P/IQC4-GeJSP?S1>3c]WJ6-1880b
:<McX?Ub1c+>RcSAT16GOJeDE;2gFV:<?/-fQ8+VDK4\+g.\47+^V]YfbN4gaN+)
#^=,<^Ug;+@DV4SC/11aI,H?XZRQGPBQ]+PQg984Q_UdZFADgRD^ZgRPBac7cVQR
\=2I].+21NRS]J75A&)DE0B&E^-](<0KH3<T]3fWV<1<?FW[@@N3fC+fOG_3/]_b
E\1_,?\5XEYGERT?U^X+Be2^LVULYWDKJIcQF4S;XTN#2&aKea[AUN>,Q1,J&e)R
72@PM#\_L&LC(3dd&F6N9dG9H+_ga+Pb]f51_#EDK>fS4[G[T_HfVD(#\APbXAcP
Z_NF<2dO1,E=9g88X-Q.?J7&O5U\U5H/HD+VX/H;cO7VReI4-T0P\aX>6^6V\Rc<
NJH/@1/)LSc1(Q[_M[L[@?A@-QgCWD\M:E=E61f)?>ZH@)-=<N]2+PC[I#>#HZGR
c+B2\?X--SB]L=1EI/-/#N,XBGJO)/YRS/3>[@((2ZNg#;0/3dJ88&Z<S9&LYf7K
&-ZfX33F(3cK(4:.>?QS9?]C]_F@eNCc.EW[Fa(6I/]b.XI(ePdaK#,C;GBcB1W]
&;E0dg2_[];LA.C-7L=eE5:EE0Q;6NT=XIN\D6MJZd=A;WbbB>J8?[&,5^?:C+Ie
;?&217a&0K>+)@7^(gKFW#?bO1]-\F8GNQX+W93&UZ?3&3b?(DKD)]O0+&[92eZc
4(PTQ=P\Ug[fH+Ve86\PHcA0_MRbN/ICb-^\^4M,bY:F1GN79bE7@9)W(JWEO]\#
C&26b&<,)?1^2H+66?M=[S<Kgb]PC0P28P4@4S3+O/5a6I0Q14T,7:L6<M@=[#e-
/C9)-G@9>7_gZg=A[LCd^J8HG6)5]\b5]aLf7OEHE(c91b)18g[bC;C/OZ[E(<)E
HLe/]b:#\Y7KY@0/[EF5B#?;W8;.g57,BI9:U3Ag@+e=01W_<E+4Y9#IPL4QNe(2
ag&QRT7&R_?<;@+5Z;cfU^PL4)]Q,5fYX?1=9?F[V+)@aOAS#)VdMb1=R,aD]2\=
aVIPg+a1FEO(6Q[G(JJ+N4X?L74e(T[X=W@;a1EfLc8KC^:]C0]S]>(OEb(_NBC\
Re:Q_cPRL0f&Z0gENBgd6X)X)E;+#fg6=,IRRP60a>HR(]:/XR(.OVFGb-[6,B>B
2,7-YaX<.gD?O\PXF&@C0T[fDU]ff)9?;MA2&Og-.:Q\#;X9N#WNYf:AUZd@aNf_
5;NK41XGVfcJ-?VZDf&0^N7,3+c&HCd;@X>#F7K&EIg<GKc/cIO&Y(VT;V#a<gMB
]23R<begQUa0KQ_V9YS&dFPTcFcb/:7L9QLVZI>8_,M485=#V(#KY44a,KL3</PE
3D#/Z1UD2Lg7HM#I\dE>9=>6T<>>4cX6aS-[DdQG[gKJ@\MP?<+DA+g0^3<I&AZ>
ALH)-\X;QL2bQ)Z6>2RYJ9^I5WC.<1593VG]A-eET:=1;T1N0M87FQAYb[Ie=X<&
K=<#2@>L:&P?g.YPd8,UfE0c3:N8\SC4e>H^<5XTX)(O\4d.P,5:_XP,CM<Zc7DU
JO:Y:A=F9DP/LR@c:FJKJ5&5>/dE>e<aCBe=g]/S2_M9KId#5UK4#M5cV;M&ADXV
\#5DX,JXPG7&OJ1SYTQGDe4B;D4N5DO_TN=W4bH/1<C3:@7KT7QK\F+#KYFS80T^
3S+JgbE?&^U2/PE.34\fIL,-FCSN&G5DCG=,>]5(5CV]=WZIGK0<C-(=e/@XG-N0
(V)1:DBb+/LKRH(-LA=a2Uc#XD[Q1HGWfS]O_VWeCce@KWgX\N=B^[f.:cY2,-H&
DRBfddZ9^RVaeOJR2@]fb_VGU=P,FE-,H3.WZ>[a:J.W4,^da>1XRaaSOM>BU[_#
BOf+SSA@M\;\(OFQ\JL=[SNA;Feg;#:<RVE#.=T[D\A<M\SW9V_2;F/5_>\1+Q]:
K/+#EKfO.Tf0dc3\#eO-3(,]KY2D<PBa3>1Ye/8N^;Z<[8)4DP3O)NbPF/Ng&RNZ
+NQW,dOJ/(A(D@cUORMJ#L-?,YbSN@YLC?6fP+WZg?>6?a,=@K08AP[CM_I+Y?_M
.F7TYYR<&L0QA^Q,LZS<[)3Mf2eMND\5ZOF6TMI(XTbcS^@4\CAJ]gS[H@8>9bCJ
O&N;;),N0V\A4H668C:\2,-[[18gJ/TZ&>T/G=6IK,:O@;JaB)26^H,:;@<\5FS-
RL@3abLW,FWDR]L&b&G8()c_HI/14cB70eNVJSP1GNG3&C>H4f[/C8S,<3DaZgc6
64P>(]@)E_[Y>g-CC5H<.ReP)RCVGHgfM42OP/#Y#?3LP>Z=GEBC0)?@HKJM&_GQ
ONZ_0]+BcdB#5]IDfK2N1FRFA)^#J(U-WV3,+dHREDM_TK4XY3cS(0bdE)J&c52F
SOEc\c25[YXP,>Q8gTCDT;_aC:=VN-_9B,&D+7(BA3SQ.1_=1M@6X=M\;=;75H9+
A[3WZa&,)_?3)Q>4H&J,D_K:&PgBOLG/,@/>O,a.#//]1SY-_D/0J(b:@OO\I6.X
O?>/YTTa)5/e)2gF?dRM1=fWRS/DL#RTS<gUXVQ.PVE#)2A=N=]d\G?0HGBR_BgN
\C78fQ;P+V)#+C<Y2#dT4B_XM84[D:9E9[fXL41JK,YJAHP<)RE?QGf4)KUX(ZN&
eI>_ea+KbS/<1FF/H;>E74T13JG[^54COZ,cU<YF6AdK:1]+I43Vb-;d2J]IZ[c:
/F@KOP1#_NGVY=g0;BW93R0ea^&51.2F+RQGR1LL[WDE&cQYDdeHGPH\WY]7)7^]
49.F[5(3f79c<E)F;&S.L9XOcNH(R.1IPL2^c_UNC\D5bOgR()5_(.6/;8Q98NBZ
9e+\a7OD9B^@20#_+IL>gaB]f-N8f,[aT;M=H(<JZKCHK,O\DNQPLd\Jf+_=68B=
&PDPD,-V#/-WD//fDBd_S@#1;08=cW-8YT)TJUVBRVUg,3A]8]1-bYY:IX;8aE((
af=I@3F3#B4&-?OW+FL]:=:fF0PO-[PE]E1_6JA52^L(7A\@-HKb(aRAKFU-c8(A
F?C:P(T86XObUPY:(/OY,F[9MYdW:.F]DeTa<AI[M0DI,&4W1(/2_78Re\_(8AIa
[)?aeS8D+J\#G&741LE5V7C9)@0DMBXO,gb@c126Y5D7,?0KZCQ;_(R56bfb(5Z4
AAW)TZ4.<_CHNg+0P(_,Xa]6;(dX<^g#WY:U@,6d1E_((QQ;[]g-[>8>PPEZF:KP
;KN;1]PIN)C,-S(@Q#?-=]]cb<(g-(SHK;R:JK:aaU1?1.,-\>P/0X.3\d7/Db4K
XW4)^L34+IEZ[))+cTORS17cF9/0WY/5FK,9T?/.aX=AK4ECcO?<T)R_c/+11C7E
C^X)P&BeUBd>)?\[76#M>J:GRYZG^[NHRac.3?VU/=#b--g#N5M&>?Y23S=SO9fM
H/aA8_3>eG;::gEG\PH^XHI)7e:_g0H.TW^K48#?()]<N[P:2]f8.c=<JE0Ma&c?
DAR<&eD;O^IW+S^E][]_bW7E7T4=IB8.<61[3Y2<41#Yfe85S4)L0T,Mc?](Ld6:
LD1H(Z)&;e<b[L@[b,#M>F__HLdVO6#CS<C:<XR>d.FE-2:4XEb3W?X6J]41bcAP
JT(5gZ\F]6Nb0+WCgddU.6P)9@beDHGaI_Je6F6J80aKAdA48)[HF/&G(_,K\V\2
@HdF^X:5B_?]D1DWD89=[M26PcAIW0<DQa;?E[W_;c2ZACcD\WfI3X.Z9@MG)8\A
UQ0)XM//?VUG[ECKHJ.@<S/<\GC^:YPQJ6^,;7U._Qe:LUL^FU.K=7U/LL3Q<e&g
<19X+G4g\SVX3CD8-;),>]R>(^B@F@E\e5+bVgbd4>>bOb1B9DC)bc<@B.6FDF=a
d])Y7c(>.\Kd(P/(/FA(F\]_2#DPN]1BBS>J:C><]J,,-^3G-bOKab@Yb2Ab.BeY
ZNS;@/W3Se+MP:=+LI-<L\B7Z0bP9+Y+7^]L#APUa36O8Sa23F;19BVcI5R5VF>V
@)&&ZMFaF:MJ14-Wcc^4Ud@-N7T.S7-Z-8QD]]R+BG8gBW_&LN5+1S[P54)8.0a&
6aBfL?T/JRV:DJ6Z,_LZ^0#?BAfAT3e=Tb94-@dUE/(Q;g]@ZK7a/M9=2g]^4QT_
H[\g/HGKD^:75WEG)2XJ@W@=YIT7Q:])/#aC.L\<-@@\#?F8gD^,fZ<51ULVRO0F
a>T_I?6DTW?7&VO2CAO05&/^-fK-e)UZV?#\2\S2XVB2+C(e6bYD2N.K5>?W5_3G
/I_WdN[gP:Gd?BLVeb-V>@NHVUU-=+I=I^4NZ64XZG;H\RJB&0M^?M-a7RNSCD5:
X:ULKC62#_:F2-VWY^TFA6BTHR;d+YU45g0;_MN[[3eOMLTDWO)Q42XM[OMGEL&]
NY(SWAH)=KC:ecGR1J#GbTAf.25M9CSLAcU;V5DY7^R)R=d6TT3/7NK=>4[SPO:W
(TX98N_)A60)LC[NQ9CfVXVEceC-ZDGXQ>ZU9UTIU)7;[@dG6:KUb?AY6(9TANV<
-EcG6;Va&MJYX?g^VH?T85VU^O]C3SS8LCecI28[5M9fS];1P]MQO<DU:GL;RaZc
LI.7bTdS?V&3\FX+d6eNB9HY.,99DHAa/T7WEI)06/0W=7@]LIHR_bZ1TR2.;I06
a_Z,O<O\(<89KbKDJfIN7G_eM6aO(b#DN3E.HD<V4PCa=CYFVO^YK7C.@DOcB,NY
X=C\Xe)Q1a_I=N\?3D+VL9G;P:0fOHTIP@4E)+;0L&4/P;g9[B&G2##ag=MX(40(
=d[.+IT>YRQ=[\ITe7dRZ3<RB;_RM9X#8>]S&N<G3YB3O.?:^?]\QE&_RLQ.f?Q9
0f=3DOR9&J6WL3P/-+?B#L+4ScV:Rg^GH?b6S3\UQS;-]+B&8VQ0e?OZF,&N.(7O
,&H@GMHUUeV(QaX(^Aa7?9=(A<0Q:=&^5OP0+P.?^ZHP?=Af8a(_W-bdb.2&+2eX
8EgZ@<dWDIbRd^:g9_@=5CKPAV+5DW^/3\-Q^WT_2d<4V3OFV_)bGV_-Jf#e\RHO
HR+JZc;[Oef/Z#fXc;f]dfdTc6KRK)\@CfE<\:@1O3fW[F\>:C0LgU+&9#E3;Yb9
ZTA[6RTKYS1W2BIIU-TXHQ\:AP@TEBI@=]bKe8&d=M5(/f:5?I&4@Lc9)2JK&R]9
Y,/a)-2La]W>2U,b-b9&a7CG9\gK21b?fR_e1.6dAbd3A2(X7Ca&(fJ/f.)aYIK]
_dFb;2LXKc?gf7J57T8>,47-HHWD1>1\?]_3^)HJH)f3CUO0NN-O;1N;]d697KA0
DGKNQQ?U;3U:-#,JR.BG(:MY3GC81;:PQE3>;H1C(cK9P+1E/ZNU-WIQ:e(E076H
LVT)LCc@;.g2K_3VVF-EDMN=QB95JGX>.5LJAK:aM)fL,a;[;4.VG,4DLCa(>@7K
K@2IO61RNXQ>K9JQL.Jd0dcI?5R=1U8IK5_;I3SS,FLAg:M0CI?-<9H,J&aTc8&^
+&DcVY/f?g=:N(\1e+-J^ZcVO1_=5:.Og9:^JRa3,^/d7F8dSSVFDS50MO=#XR3X
FL77B3?Y^M#)@4eV]QR90M[7[MR--I2TAD5AGH8J/>L/&bfL<0X&UgOFdF3JHd=M
OfBY?b4UDLX7&&Q0:5B-84(M7(V)\D>1DKeOW44PK+-O]33@\@7JC/\;ZHLQ[R+P
D9=GVX5VCX:(,,FNU-ZTMQU0T.]fL6B?^7#e0]P507MXOU7LBH@W1RZ7_K0O@Jb_
?4H1.62\B9[JXJ5GP2)M/\_a#aF<OgK3,b:LW3cVe0eU/Ef>H9^[L24>#UW49&WP
18M,KK4aK/=0_&d);/RgRgKQ,]1RY=OY)UPTc:AFc0.QDTSWWgXN\<.KD?;MIA:3
9;Z2-Ge,JWVV+dRb/b8?a7TQP-G[]]_CJ<_C+8+Jc>e?Ta8M]CRNRb7V)+J+5YV6
?.;_6A6AcNFVc1bOZB/Q\?>CF#0:37UYZFW_eTSfW9A^.T(.J;(DJCFMDRW;6WW9
MSeLa94B&^<1?Q?3ZPb_>:KGaBN\<If<Q@0K.bX0#&UL)S\WW@+VQL8)^SfCa,KY
9fCJ\\K7=+]8]a+7;8ASN(6D?&1&fDTXXbN0eT\S:)G:L<LJ9a3A+D_,fgRLOM9^
#QI\M^N6[cF,L7TVe@5/63#[,F69CZ::C.O(&\VA<Z:R5fHX4RBXIWW^Z5R_,0[L
XO[f+(eOXS2V#19F8GbSUbEWJ?2E@40d[LRPfH@d<Od?HYMKF-&:Yb,@c,e66<5)
XUM6CU04G.8DA+)f;\CK-N-MTa;I\^)d@,\2cZJGGTAO]4c0<.@68>c,WZ?@U#=Q
SI0335/R@;d5++?f9[a^^.RWZg_f>Q5aAKZKDD>BKJQ+#6=DC\<N-+[HdH=dAdXE
<^FcZI],8(M2caEEL:)(QH&8P@C6_1S[JZg9M,.<V0.\4<_+M[e1^BH:dOUIQ1W1
;8_#cN,X,^3Q\ZV)HUOZd7e]M-UA7OE6)[[-OH5XW^DK1SZ3>>?a6V7LF]?K,eg?
O+<;\Z[YWGYGXO+-2Y;JOOWaI^^Ac0)IMGA&d29<N)]UA@I^Q3X/=T-^M^,8]e4K
8(f?FKY1gKYNW_S=MC7>afJ4LIgU5KILFcTJ#MV+UbM6#]P8P89/DT><D\-@gA^U
:]C0fEQ,&XWH4bFPd-\.0TbC#W^42:b(a<5>I4Vf7^R62d>1H2MTKKdNMJE+I1bI
)(DYd:.XD9H@\_D?.K\/bL12/Wa]^g.bT01+Qa8bW33f9b]DQ=]A\.TCf];3>Z2T
\U7da7K7C_+DOfSfT6+f2/cf6SfI.]ZPfYZVJUV3CE[0cOS(IH0RMED#J1gF]\EO
cAeX7J:7@9<Ia^:9&EeKL(Z2,.eH\[.[cTL+&861#/;#I.(<O&aLK]4\L+Ef?9EZ
Td(PaV\fTeX,BbVQY/WBV7Qf[2L\:D-KKWVB_:/E/GW>)M+XJY-;&757b#/MM23^
B0JUb4=N)Q-Cc56^?XLQ(\8Rc7R#(N[Mc;>]U5-@P/;+@.?.@EI,VOXWSVg^c>CH
2C5cD<@Pc_LX1&<@7e&9dWG)>)@H/EcO1/MW2]5(C-BOHWJ46L>^Vc0OD]/8Z?E(
MI]I>3(H5K;3;aIMI=/VF6HA4dEYOJSSTAfXgfS\e-]3#Qc&b;RRab_BIM)-S8I<
>.O5fEQ:]S-OCM[[_V@)bJQ22Gb82P_OJW8QL<2Vb+#Ra5K:@SO;;b;/cTU@SJM=
fK)eHV@dU#@X4;6/QT.fMc6=#MOX&>NNG^A.SAO5/0:<6?a3DK<E8-<4UV@+1?SX
^O<VRNFB4=Z6@c0(^DZ(YGLYa#VfW9gfgPN9HMH(Q=RI3;VZ0@MJZCY#T?K?>BEO
_FGVS]^8WUW7=[ST15MMDDLbE?B#4R81HA/CV1HIW[eCa5@+O;0X@#S[8C0S8YH+
gJ>_J9a,JOY3H&9S,VfQLQ=c]7#8G<]6X2>Zg=/4bFDPY#<F5ff7=DG0BQ8^E4.d
\(>F7T8L<W#PL,_DVGeXg;:03(VSV-EgY;S=U1XGa@C@#>MAVA/_+YIZ.IJR-aA<
T.V<T3Z0NFA&J5BKLN5_RT_BX,)U,5d[L.g@7MOP?e\g>7;ZT)QbI)L01C+C/)Cf
2FBO<@#O3Y<W=Z]PE<L-6FR1C)&23OTCZGAF-.)E,2N#I9=;[BAZUTaLF?PJO@1/
E37-#+-b:^QUXKE.+aRN)?CQ,0b>E-#U^8]IgM.bbX#NWTQL9XOU@_\=_ZESP_Pd
.a4d<JYJTB[>G0M?##7G)N0Q-/eAW_)0:BSEJM=9gF_a?HE</GVV<c@aS7[&G#N^
1&cg).K\.gSe?\V1Z/SG?(T^cAR[DNZ9JMT=f^cP:C.Wcfb[WFMBNL:8_e)Wf=VV
5I_CC63&YQ,fb0T5aa;W&cWPQNWa\/[e@NIA;;.H0.HGfNF7O,A&XB>HAA1]bZ\W
\dXWFT4:W=cdB(Yf/@bM6Qb)RbPGUWJ3:(4RWb2N+XL.0UQJb[aP7LdDVEZ)-GIK
0f+.;,A#-(@44VW=[5#-;9MJ+Z8H[M-;O8E-NJH_T@V/YdZEB0O^c_IPc32Md4Ag
07HLV@/EJdO)9.e4cI85XYA6FaMACL81d;TIcc-)AOF0YKMLJLg0@^>=(1T(YMQ[
5O9S5,ag>g8E,L&-;RP(@+N-=g7JW=aA-2#+VRI.HeeNY\<BOD>QFgB1+L1QaAZ&
J7L\_V_FeZZGF)ON#/QFJ8JH_?[TS>f0/C9^3N(B\B=Y/1_X]b=QA3C.6-BgXPf-
L[B&[0Wg7>e&5SX;T)GO#(J@aEQ\(6A=JJQHBe6B=:J@cRH5)QX;\D.a36e4ZYHK
+05aWEG\Y3cCCgOb/a+Re1ccHN>DEDXBRBB:;V&NPH1F=-S@T@,e>WL@+K3T@ddJ
)/Z\[Xg5UT3^aHGa(J@a?/<_9?(cd[5Dde2gIYHfL2NPCK.KD^IO#[V5.RG,)7PZ
dbg+WL#P[C@7_&QaRf.P_O^fL-1.<#T,9&3BdWTA7FcQOV(_,[gU]?]HLQL?YG>L
>3+LR5.\JbaCGR.TaO(5IQQb;PMN+)X-KEBNUM]BD;a<BdeQ]C<#;+A-d,L-cc>S
FUL=LZ:3>M(5J(Q4X51]-=C8<XS9]Z<Xd4Nc?FIBT;U^\\LAcJ4a;<B:&O:ATV4)
a)HK>I3NG[K,ZXI;[1D)/P&LLQ<J;g<Q?#cS[]/[=d_>bQ/UBY.bRTJT:HQ1I8;P
3R_T5R-5#B:)d#(S_K9#/GMD]PI(0d;A^c5O0&?@2-&E/CO@A3H)b4WI_bLE+6&4
#7Q3&EV#2AaK1QAf<C(5Z^;:APKba]Ue:9W.NY?2YRBN3JOF]2=[a8]+6):I6Sf[
2T+Na[DEHfD]ZDZd:C7RU0f\>+eDIXaR/7?6>HRBV_C+N?.EB8TGNSH,SZaAaQS?
M4H)D1>7./<.D-RU:Hc5E-(-#61>^bF?))&UR3d)LK/2EETA#(Rad&G,>:,2@I6D
4e3bMaY+/UTEC_agA3XC#ZY_+MeBU4O&72cNIgfb6.I:3dYYHSPd\ZAg/eG1W<-N
G,-88B(A/I\<1H3\Q#7G\US2ICPG>X@XV7RHBYgFV(&N@AVHT,_[0F,WScH([c4[
6RK?+D/6S9cWOaBFSR=9K9K@\g:Q66JH&VQF=VJ[=I09aG+CGdDegA7d(WOEW?Fa
5A?R<V#XS&@Q3f-:a[>TYMF6_3cd#bE@-0V9&d9I&X_T6L/Y_(Z4aELY>:NGNE&F
C&1VTgYOG;,JR@e[^?^dM=5dW7cN&QE]6LQJ77d_ZQ?39R-GXDbV7BFf3O/[TM#6
KWIaRa=d?4Y5==:17I4BM#Q^;#S3<K+F]d=I]Q:0]2dfVJ81b[V(T@X(-0#Z,-d&
UQM,?&R>22,^3BTV?F/^02QTNHDINA4P[&;;UNTfGLI,)g-H=MC9J]78aPUTU^Y7
4;Lb?-@-COLV,CA2;NNR,&e5P^&a^]I(U_4/VJ.YgUaS;MKWb80LfNc_3CRHIZ7M
+I\[2dAS#5KD@5N=IgcG2CbLB38b8?0c9dBf((PHQ#eaGGaf83T1Z+-E4,d&,R9M
;X3.I^;b,T<@O@HIL1;(2E6#S;S0e@8/aV32GMD<>79Ia+b6:AE0V@cVRBN;#O2A
Z:<G5>CJ0Z[\H(.>?-Eg3KaIbP)G.FSTE<4\/.A3_e35D/P-Z)Q7U7b/T.+9HcYC
?I8XI1S6>-/NUO@f?M=9Y#/174W^-+EYPcJDY+;(,^YCJ]H?=3VZc>?B+B6)U5QA
A^=W9YIYGFfOWfg\T:aN_KU2GGF^S(@>O9(P/ad3\@7WE9#5,;O-R0,gSc3I4T?#
=BRAVLV:[8XgE[?I0c^e32REYW/]=[g+^--b&JQ/>EP\4:X##=/GcU[7#\?-8NQI
;IWAKDGO]QP90AbN#dKb)WBL@J#,<gY,&.e#VL;bIVVQ,G<[J;95e[,W\3P>#-24
@JA<E7X,N[&Q-NK>\R;e2Zcb<M8A@F5M^5dP<R7bY6WXR.#LQ?<Z6D34W_g]-U;g
L[;OYNDU)R,7W+1_J?BLO@P\D[RR&eT7fG?,OFC_17a5BH#\I88PA@]EbO/aUO?&
EZ5)^g7@NS3./F?dO]LTSQ4HZ]C9+B]C@OfBP<]3AeLecPI.N,PS1/cL>Z=4cG>-
?Xf9@LaAL,&?Y31cE#T:U#OC(d1<YIa5E:D00b[a=R)K[3&>)V=36K8)3E].?FOW
\@Y,T\>L0@1cYWR^da6HTF+P70^eXTY;?=<<9d4=6F+&D;F=#4,YbO=cJ<&H#:YV
aIXKL_TH]c^OD/>ZeK<1KY?^_^d0?DCHMD6>K;KWfC3Z;bB0.9O<8#O7AN>)@[JI
2[OeVZBEW^2^_2QBO7(8YK+(&b+K<T)R+I\Y49W@K>8^Of(QAU0U@d95[4R;DdC)
dV-G11;0OJ#9#&>_[]DZ]f4IJ.<]L0b=C0GfPIVX5H2c0@N3[UbU,7^Y/+/?P^;>
B.>Z3#gLQf1g&/[\(^5BQY<)3NaP-_MI/ULMb@;cH+T1W)d&9C78(BN;_Z&#9g8R
RfY@?5&5/[\IBCVU\f>2AMKVK#><K#N\K@PYd]2F_4d+4F7g#Q&;]7&)?80TdEJ:
RgJX@RFGcY0d\YPb-K<1<^Ag?(X>9Hc+OP8/fT;=RT;#BC5O4b#0ZZKa(d^eAD+b
QDeKK)RIP;AI@P5RK;N;W4U7^UH5/L^3fBMP>J;ObZD/]N46R?f=L_c7>.&MO4X=
?aM2&Z285cb)(^JAg.=_#G5JRG.1=[1-APEN#4YK+gI/[<6JU\.+WB@g>0Le&-)_
?3R^_d8FWaO0660F(5HEYJKN207EW:3O3Mc9d=GG,F.6JEU8FO]^8Y3cf@<(+KcG
8ZVQgJc=(CS>gGZ+A+_Y#TQ[:@c)=&=150AX>O&>?AAO?&(T4Z_Z0:/YI?5Y6-K^
0X.O2db54b^3JFNa,??_2_CSEZO@N;,F2S<\]PC2.2bF_dAAbA[V2;?Q]8BS<1gS
052AK@FWPKCYWF5D-5X#ZU#\:9RI,gJ#AdT3#TXG+JM5>3>O:SRVTOVVg<E:GQ,,
\QGS/6@K]O=8LZeD2R\)f^Q^fF0@H5XT^__LU,^+:,C;^F\a?;-C#C@QT,BTG-5J
,g6gFRX6?eQ_bA/FB15PSHNbd)_:>4VE_GUOGA]E=4<3,1\F<P>2)7DJJ0c>C697
#)PIK>:0NK0e/R-EE==@^&-^Z9g?Qf76+JEY<6D>CWf^+AN?ZRf9IYDDW,O?\ZFY
5Z^9F=TcHPPAUf[9-VT0b)W:+.(Vf5K-O:&T:?=_fXa+8XMG[W#H@b@N,G+=0.df
^<TD@Hb0&&8VY>P>#P[&-(FcgAf.JF+4.,agM/&LK<LV&[fg/;D5.-L+9/7TN-g1
33Ld@&?.UKA4)FRI:\I4dH;]-UK>6dM)[LDb8AM/#3A+[PH4ED5N.SG)(QEG.3PD
H;XK78+a[R9dYE(UL<O\>?;+WDYea?+>HYI61L@>+QX?F)]cf?_a.KJPK)QE_H6T
4>MCRADcL-BN;>,]AVSDO:-]KQ3)S_Ue^YY2:f@FVV=HD1,ZWKeZ1G-fYUA_[V9<
[,Qd4gdKVe_TM?3cce,>+),+7>JaO<>(ZAfM)\7<9eZLDc\[7bGNYg<d#PMO^[XL
A(c^ObN8F/bYAS\0YKNT[N4(_cU#=Of]KAWT\1L)F?I=X4+&cQIJ@/).e44VYgOc
(ZcSW0gacWbY#XJ121PbZ:fHA6JJ_80+_2#.edeE=II],ET34BO^+YcR6@cBX9R8
TOeRIL&ECTQ&HU5b^P^U_\Fe<UMIZ)Q&8FZ9.L1XPH.5K/@?ZB&(P8-(fb6I6J:?
X5U2EW0IM#QPABC<<603^N8[?5=[f_JT.cK6Z]bL/R5M5B\b:=fOYP058O,b_AD]
/1[&fA9=FPfE50M?9:+YVG?/64OK:_NCSc#)C#JZg55gWZ2X=ag7QQ^4Kf_53/e+
[90.;8_E60DBCBT9::HS9^;1P3ZLH4&\,>L1Lc?6.c:>e_6[0>&&PBA#KF/S<cG-
KO12C_^@V:QJBD<DgW3cZ-afX7_)W&CEN0GFZ(b2,f2&8K_U<QNaC>,dG>Z4O3=f
(@]8ZQUD[5^I750;.,PXbLKWed(BAU6bdgc4(E5:+1/Bb10LU4F^]L<\<&..,L@J
D<-)RXgH(2f(2CSB>,Q:eLQ993CE/87)CSI9bd_CA]e/IVGG2U6+F\?cKZdf1J42
B114\ZM)0@6H_&1/RIQ9NWP1[FNcf6<#c&AbQCT#EPD)DAH#;WW=T+b(LfXI4D2B
#A/H0S/RKHSgG[5H;Z<KWg0FDFbLb6)VSFd14RfbNJB<H:&OBEIXdET3W>b128.(
HI5fB(\LD]I=-9D[>(O3-dN:8-W;3Dg-.V8aL]K&3HQYcRQf@b,A&aGWU;:KE\Y>
^IE2AU)[fLAc,V2MO[7b8cg-6-YJ<Y(6A4;YL:MS@a[YJI+#]58DFc\U(Ie]-090
f&DLKaK@RUHg-g<NW:GH#@@E-3QeaIA>DK.C2T]/@Ed&RYDbgdB_FW.&I33b[8LJ
6A?2?)MMK1F_6_96TCC16<0YB/RC-CQ.4;LF8,BDS=_KG0dVbWc)AY&/,SO^c+Rg
3\FO.ZX.Bc_gE)QE3V[f2LQ;feC6WLRa&Z[)E2<gOc&C>-(4/OWHAg5L4?C0T]/c
Zac>6KCF3CSB/(#4&NG;0>9V\8:D^/A^aF8]_8Y#@1#.==T6;0]gSc+WQEN0A[I_
F[^KH6+L7U(Q&WfTPRe@PK\;gH<b8,6Bc.?bED5+HX-90Ue_J0H[X[L<;bW#NX:3
XWIZc[5d/LS&5<?TK,1-^247<R.H+;g\6QDaYMN,gRD&-.<g0/HZV&&6JR3O[AC<
Tdf8RN/6g@W9_CgT;YPSW_Q3\1-2PG]+aE?F/L?2dL@IY0c_BWfX6RcWQg#aS\8f
6a\R_S:?JQVg/.WB6]8fCA4^+4b,^aMP6]dP9ecD/G/]50:NM[HJTbgYUb..+(&7
9[\?c37<&K?RJ#(E)?Q7D9BZ.-/4:.+XT2,e+b[21bEd5PQeJ[R)OURB<.K75&#2
R.f-_+RQPf4/a3ge:WS2?],V\fdXB_4/]U0RccH7@4]^F86e6;51)5,2dc?,7@\+
<RVG?>?J/O_H\\C[U&c:P#E7b[<<;OS3U3T&CU2abHb&PXgaER?22G\S5XS^g/1(
aXZ]H>8:7X50KI->V5LQ@8PI_@NMQWf/IdR4R>@HIE\b+\G(8UT@^\K@)UeNC83D
+];cYU4,CTC(:WOXQS2I5=Y]GdJ54e+EVM\EOEGXbZO1NASIOLgZ-O9PU;05N_XQ
04[PEWf-_]E\,CP+&b#32Z(d05H3,e)NMLLG=/1Z2\5Ng+>)O47g4WQ[G;N;H1X0
G&I-G^2H\.^7V[9S5R6RRf2KTM3]@f8GbRB\@@8b^\a_\.>3G(2I9KMO:,V\,J6]
\2PG0Q3M:U.UI(EC.PR<eD2:9W0=_9--g]B9HB?M]T4J9;N\/gO6-4MW5b9=36I@
/P@9-#+G1/+IGIcX#)BC?K1>K7;#2HV?8B8X7cZ/7631f/H?J6J47BL@fY<XXZDZ
V4=;_Y-Z51#,5Ig2/K8:JMUNXS2]D&22;40Y_F;8;c@d=DHO/K4ac7H+NVUD[P3W
5JWc2O.,Kd)(^)dT#I@R(G49>e&7Q;DV]d^+UVE<,.F<^g1;9g3#1He&a/ZHXGOT
K0AX4&:9^3^@;OAB^-=S?6X4U#P_AAYdfO]9]A)ZQ3[SG#W=-8ARcT=[,([D+1MI
8<,#N#ZA]BO[QV>N3cfD.H6I0NG\cA9@&=RAEY,M0CJO?Y>X&ZD?8g]:;LZeHRVe
OT6QY4f[33_M8F:&MF=bXf.B-<RL]P7MV>J[39,JFE_];@.gW1/X)>SfZd,eJ8IJ
(=XBPN(5P9e>E8Q5LU^2KUP.fT00Z2@>dF\\YHKQF&bA40])[=&WIREQL^AVc#9D
+4.9bRDL;I;+D.eS^UCA]HG5f[.YPa<NP-Rce]U:267WbE8;^TEbM5Rf8AP3S@cS
_I9c1D&FSdgO.0XO,Uf:d\8?>a:+>5S;1dI/cG8]?KCT)8,@\YF-.];LTG374XgD
.&3f<K3b7Td&e=4eHDN9#3EDIUQ:S@A/^]C@LDJV<^T;PM6.cXR:a@Z..,[4LfLI
U7MW.74I0,V>aTCb.GHIFXJ/^;g8Z5&a:X_OI6DN@8\?&aV&183O\[?G^.86K;-=
A0X#D6gX,.c1#f>^MVBEN8482P-Hb6A709;9@Q&gg,W<JAJ2;J[+d1?<27UIVP]M
[>:K@KVON&D&fMF=D,&RD-;,Xe&P19fR>:d-bHAR^50B.4^_d\EC]]5?]L1U^/[:
,3_b.2EZc>A=46Ge&91:S/H5FNeN_/-FCKU_F^T)(SMGWG37Aeg1DA@L-@VLEBd[
,5YEV-b-SGO4.cSa]G,UY1)V?T<]?g?M:(6@G@WT?Z686L9fgZaYO]\d[5dcd6f#
DY5PD8H.g.-0P0??N8;E-:3#J?1(PX^JAD33?(J,YHc)aZ23O:7RB(aRbN:I)2,Y
4c9d5BJCBf7G:)[=g3T=Ffc:54TcYS-H8TFXAcOKYHb[gFX#(eaSS9bQRL:eL7AB
7O9C9(FL32>W4PWD]:.8W?Q/QD3&6D+:-^XW^T+;[YG5OR_-4K=5fH;<VJT/T^EA
.b?A9b6dFLTNR[[B][FQbFR1_(D;[,R_J6cBJ4O3/Q&(,a=EXA:dZL5G#d&9O<S+
+2CD?FD7^G,fc<:Q?WNaX]#0)bdD>e<@0KK(5-5;KSYP)IW=:S;0d[^-.52\7MIb
]4?Q:@K^9+25>ZXFRd:CWd#b25Xa++YeXGD]d(ECT\4HWZ.W)b/QZN76FU1YQ?QK
aN-=_CdU=A[P)\)9Z(dgD/M4X]2d6>[5(8W36[B\_TdfXG,.UcISRCT3f(6BE20=
_,f41=bM<Ye)K--O>U,Q//7G]2WEE^]@&^c:XS_^eg..U(4HWTd<A>H)bAaCJCP)
#d-_<?AO)&69.):./9f_f^[8U406JdADJ^T:7dEVbQ@e[@N.2]F1&RZBQgD,<X8e
Zf?;FIZ&<MgE7BU0BbEMN?M^,WDV[;>?I::aM/;+YPNeKUP:a]ZNQ-B>?g?UIH8e
(1>_2bF10<HFZ+]#^SZT7E/Y80KL_&<N8gC+X4LFPP.DT8:GD&J&J]f7eS#cJ&Rb
ZM2eI_X@KBcPH@&CD^+U.;a,TC=1a0g7OY[]CP6fL-TBU/eO73aCS9-@9HOaU-PY
X0_N>FG4_a2C3M5]:(?9-A2CE^6Q+^K2])/6b5Wf7^7O.CRD&2DK@N@S2\,-C+)Z
H1HB,>__dJ-OC,^X9VEAI(74=<(V\ZZ;A5FHBNP+,4B^BV4b95f@V.0.Y6_SJ7K/
2Pc9LB<-e]c;CX6:)IOTf_[#[RTM1/>JMC)T&Wac/&LITOTW2+fJ[7XKW?b8LJ-X
bJ1#2G6)]O+IZA^317RY+?HND.8?5;/e]E?ME,)J7Jf?c,&/5.4H3=b(,8b?29:3
5J^PI&W2:.1Td,MYaTeUX;Pd&VWG^b2W+c_P&[&T/?Z>f6]#<.HA>69,A12Q>=QZ
,ZA<;(Na5J?_EeAKcLgBLff21;M(<I>+b1\e7S7W^Z1E7C:WP&YP1YXdNE(@(48L
VeVd9-1cN>.OH,IX]g@9_)/JVF?[8/,&OM1[JR-Zd:.V;OZ@3KAcU5)^8432/H_R
(Z62PBfY<c7gQ51.9B=4\eV)7)IRf@06+J7\<T265]BG\5@(.@?)Q)24#U#d5Odd
4TJFZeYc<_fC,,Aa6.ZO<14GUG#^NP(ET4@4a=)]E5US:#PCgD27e]W4#Ag\1X_U
8=>Q-cI18Gc=FP[Ub#]@\XRCOTX6,UKS7=R&K=&+gbN\8eMH>/]0Vc+24K0/4B^:
@A2+7MWP=.<)[IKNJ7KMR]/2F5HOU^XCBAe)Og@\UHJ5U?,MTc31bSK+?^,XZgXS
eX[3UUSI;La0-eU.W:,gLg/<()>FUD8(GbTGNd>R2_DKQWT0E.74&B;&FeQJ-^5.
9<\g<C3B\DFQ)8JgA3:Y+4-RB/PUE@1?\K[U(+Y>SBQ>g;V#CMbaKD-GA4gPU#Xe
7=]V:2\O.@]F(f+#QVW.^IG?=I;6:NUFb#9P2dN=4.CO)ZH0_S0#06UKZTB\T4X(
AgIaScWCDHYEY(a7H1bM7_cEa72)4^GJJ02Y^WYF&_+K?:B,7(FW,-TLZ_4@93A6
+_#E7A32QT4X5<(DC8a?(X5E8LQJ3@GT>^U7+8VCbe>E3JXaAdI;8e(9D?^D?F:+
/=f#ZB-c<2Y>#2M;4D?@JeC3=bR_3GLQ4)220@1NcFG4A9=3+&H#GK;S83WZL8M6
]Ha513.:Y0a0gUC_=d@_>;7-_^=NPXBWeQU#:AK0;fJ59MS2aJ7KM\L;?>8Y\1Fb
5F[/]83@-.X^V6U^Kb<^=^=63?R3F./,]#9OQOK<H3(SGU#fNGOfTW1:R4NXfgVR
=FB(/7a;)M<7:#HS<]4(3SQ#WcF0UGZc#G[O]JX2680:&&UCN9<T>d1Y2/D3N3;U
67aTe)g;VBN^CM(Z?b=G\:6XbADLPWZ56[LJWTPIHaU1F\[NZ3M1=.R?/.C100EM
_&+KZMBE+H[P=;.>ZNf7;D(65FRU8K+X&Q(@Yb8CcTO?)L7+[(a3Z=QHd@^GJYKM
(DD47+-O,EYc+^5JC+T:48V&d]^0OG-8-1EVf@17IJ-6V1.V3Cgg\W&g-#g:N&@S
AT@HU?7/QD.B/X90IX@[>MB#H[;>3#@/c[=W;U-e])4-:_Q:-<FWaJFF(FU1O9B@
_aC>e17)g0EEEM2e+g54_LEQLJ^LI&VK)X/:XeY,GH<F_UAUJEgg9=_4?PXc>_4a
V-#UG5Qe8;>,/EbHS1F(dMSaZ2J;[J7\;6faBF8F6f-KJJNe,TP>C5eCdEO=44+3
e@&MD20RA34gR9WAXSV#FETJ=F4>E]B2KJB^IbLg#4K_1RTR>)g:e7?ZN<FUI;D3
K&VE41</)YE1gO1>ZXH]+cfXe<(#3\>_Y@+c=T69_TF.cOD;?M?UeZ6,1GOdVBE0
><c4GF(,NS@SZf_/<_.5+M_FcQ)+0[g1Z.a/DOR;4^dX<@T9@_PfR(-fG0]7aY?R
D+G/R+]ND3+U;cg_6)VN=5\eQ+SQIgQ;T[1>-P8O4Cae4##A:SV]1&a(\53Q>fTf
dFY?.V+W,^+XK^3CP7@M@K&4e92#C^Oabe]NcfV2L,6=ge(+BW0B#_=)^9IIW7#]
/P@WSH^c:Y=X(MJT::-6J[\;I<M:(/R0ILF+gQ3==&.bF2GdH>;6M1OW4K=SZF,J
1f36#VA3PJE]O00-S]1_LFe>D\d1I/2\_0M-9g:-6C<J<cF8BC]5:XF+W.EUVSP]
+f7X8.F>]TB8LdC0^]0C7@BQ=56M?D@&_SYL;-Dd9-dP=@bV)V4@c026a\[a[-SU
@/J62D5CJfP3--3RWNOWfcQBcOW]ATd#9+ZYbb.5\c+K:7-/R639>LM@OZBSU+O7
d<V]=\ALD69Y>@c_Dd2O_MH1/<TC2@7&Q);Vd?1SX_7475>d5aD<Pd>1Q]#@)Wcd
BNXJKU/XWOE[]1;MNK5I]ZR9UV>]66,8V41I[I=23=B:If,W[eOgQVDE#RIcT0aT
g)+FX84]5DX2b<:0(IFK&THLNC(cY_^9d7VFcJ\d5:aNG#R.\c)8Y4WN\&;I_GeX
e(49X28g4KYZ88a8E2ML&T8Y+[8NCKHO3/:\c6CX5PAdOgY+<Z+PP(ZC^U&FITDO
QE\=-d+ANIOT66,,AHIW+9)R2L:\Z&?OSCTe[7R.4cQDbeL(W^>F?=2,6(V\/^F)
Y],Y+LN6WZ#3;PbB0/Q(bT_#;?P<9#)0>>(KN4TM8-LD5>2TOgNSZB/SXdHgfD(&
3b[f-AbR1#+gI4:C7RI1X<Xb8MU-M<gZGF:I>e=O1FbaUFU]M3dd+De(-g#6W6]?
[W.P)>]6a,4HR?5,RS4.QCa#;]:,S3M3JKBR\YfHI\=GD=cEWGIJM]BD0[6Xbe.#
ZE?e:K3RLfg5=&#H_PZ_e^,5V)/B_S[0>IJg=]BWcCfJaTNcKc2eBTEXD/^O&YWA
BLCIVE;8<&818JgRH9ZMOAD<X^5(GQR\I5M[5E[aTbXUG2eEF6])(NQWTXfBO7\)
I);?Bc:a&1;78-+S\fYU+1L>22HNZ?PWSM)SR/JB+f9RGTW@Q1MB5YKC_f41MU(V
2T@(Uf\a=P.b\.dWa(AGMCSI0#,AKD<65NBMM>CJ3-^PI#NZT#WK\HMQ5#6G9M?7
;d,(6R+VF>TPI.dP_P<P@I&[EHf+@<HPJ?].YD#E,B-H;JHD2bOL+M.Q<5[YB\/B
,&M[]YaHD0;CQH9Ug@LVX>=R6BBdb,=;SUF+<Q_00];J#11M89N,@GeW/;VLJ;eD
.8=O2K#\18eaJVPE[D+B=G8-<[b>ZPgMU&-H;6=:RRSab_H,<&3[+QW</+H:EU-\
H&d(;,YJ2eKRKO:fK_fKd9bF/ZP]dFNcXUaY\_U1GYWGBIKECY69G;]F.AT_O&59
8F0LEM?_V&8Y=T-OZZ<JLQC:J4H6#V<(4HYSb>bIG;+JT#/,YZT>OT+PCBE2P2X.
@D+CHN.VUOe=BD/GOJ?A\88XW,D29C.9[=RH@B?5dA:#).<7c)_.Sg/-ST:caH00
e/#F6/XEdF3&J.-#fVORNMR9DHL\0R[&dP3OU76FgXASQTMOYK5M9IY\L4[J0)P<
F#afRS:&XePc#YZ.B&.GbI#@?TK)Y=4SD\V(HF/C10c9[8c^9_(R/c7@?aCG&]IL
O3Q)G@CYN.E#d01OW?\2K,&De5Y1EgM.CbJa@eBHSH5WO2N?F)e4dA&(6/@1,PJd
5AJaH?:=EG2KbHJ5BAJZABD<NHLG57V7afRJ/<T^F86N,^0GAAR>f3J?cVP^4,FS
3DdaZWaLQ;LPM9H&JWQ,L<N8_Z+XPWQ<F:8_1BR.(RTNfeW.0],<+ZEPH8AN[c5&
Q>e8EV/^CBcM<I#B6Xg,L5<4\81=ZCZCga_HYHa/7?bc1T8N.:5?]F,32&7a5Y3+
3>f5>O5<#GE92_1Z6Y\QNd-9P\B;cU,LFa/G^7d;_>cIKX9dX_/B=9>7-CU(N).)
8KD:S;VWdVX[GF@P_)BdR,f7RL;cNF1-&PgO\A?e]=56Q)b.P/Y25G0dBOfC7__M
NPafQXIO-IEJ1?K+GFFa?,3<T)^MIJ?U#80CK@#T:Xa3/T6?4a0HEVI-#8@Bg6Xc
RYLG?:^7PIV41PR6JB)=QM)K]cdMC0)F([,H8f3AMW=UC56Ug?AKN(1>V;JR-_K+
\(>f7.O<Q7G5LTQQ[eO<K:bMHg<c0#Ga^9>3#4\0/;8@TX+C)O>J4]6U3O8K:M]4
U?2U38,9eL6GE070e_aI:I5#O^.@dUJRB8(IDCF&7^9R_a@BKUV/:cgI.E3\<XF,
:\#V_V0@X^W&6gG;^_KS,)F[5R@W;ZC?LB+LXYGGZ/R4bd3aLO+R<G6aUZ\9XSHK
=gZM86Z&+::ED50L?ZHC??1V=GC,>f@D-ZQ@OQ6H\,Hd&70PC0KC5]2[ab>-PTa0
5MIZ>aMO]_S4X75);M@eT23R5YAYaSbRHWVM0>?a@<NJ:(2B.PCY?G1F9BHU#]S5
\240N3&b^&#dN+BN&LB0Y@QVKBd?NY6Z=LaV=[MNU3LAE@B^,)AW@5J&W^;>_,91
Zf)Q9.LQJLd1NMe,#-DKS6Y@](&^J:CP5>8:)J0Se2=H93/e[_]ZIUIA73(5X&3H
24ZaTMNT,VJ9R\XH\7fQ(Vc#B^/PGePR#aOdgP((Cab[a,\:^V5^B6O)>]F=PVfD
&55=P1U[)f^6V)[;P>.f;Me8P96=)b5@CbW8QP^C&4;PRKaeV+gWK1C)WF?Z086<
T8b/:YN/)<7A<LQE#)]UECKKU^/_HZQ_M+=E+GU=gB)SMd6Yb>V0_HJQJ#HI[+WP
[9[YN#PT36bTN31J:b84GUX4UWKCN8gR83ZHG]PUBKg?EE(W^@^UW.SK=fHI_=/M
f+d\g);^Q;APXP^T\(57^]4H,52/fAMd#DOC\FG_QfUV#YT?0-(VS[M+EAXC9VQ>
dIbdLF(Ag/^+&SVfW&<>G#WY7R8RD(QR3SDc//^K=HKgNE[W;8fH+d32XY4d4Ab#
X@K6&=:UK2>dBb#gNYeP66.]UK:R.1fL.Rc[G.X6P4>T?XJY)XRX7LXMA5R4V)XJ
5KV3D1U(d<9S]6?5#VUOCC:]<&cD_+,DL[@H5@6)f^+[IgK0VSQ?QN-1,FQV@JKI
0U.+IOJ6X21#<8A\AG6\#[a0]DdLb&A9gK=7&54U#1SgbP<E_>M1=_aSVT\8#->M
DIL3f1+^#-V1XX+J4a6bF42HV?:#O.P<9L935\-^8+7/QG8Y22[2fF\20e4&Da,X
<S[I,].O+EEFJbVYYS6c,QM[?_][;FJIG]YV1)B&_Pb(F,@\2_#&;7ee[aJ>CQ^C
AH\22H&ef;-@&gYH46688HbeG]4T<Zg+38JZLb+c;e#D^=Z9+G:6.?9+>&e3^Sf5
T?.<2J6B1V]DFdI0)XG+GDY?OaD;&XPP-=GXIVX#(4Red]9EfVG@6N1Fg94?bHPa
:g.S:2/AP@)ID\aIR]Xd@-E;?UGcg+EE2RGY17HNW=J@1>@2ZF51a[\8:BgDT/Df
\)S6CS9ZP(;LgMV>#bM@7cOd(g?gd>V:F_6D5R+a6(W?@fP+#/)-K;&QZP49GMbf
Ef71bgIQ=K]^8(2H@;LXH@Lb5]@EO>XUAE1K(]HZ#aN3[XCX_XEX@:Zaef0g/NY<
Xb6AF+([dV3)]WQ6/bF6&0bgZIfEE2;\-V&ef/@6V,EQY>_XJJdKM>KKNM-=/P)3
I6?ZEG\?c=EAZ/GFU[c65LN;QQ<;#=9+Uff/84:TG;WJO825eGI(5;5D8D=BfW5\
RM:7SD<W\cD_5YSX-Q5#IO;<^RQ.K[07f>YFGE)6]M<Lf@[+46RK?5&IgU]=Q_b@
65UB_?@\8:=f3=^fM4dOS@JRZMg#;+:K<>FXCPE#A2=(7KR:N1b)\06H^gd4Ug@g
P82g>F@;WI]7e^:-\bOg)FJ\0C03QIJNKK9@T-ZQe__M.]e#(AH4OU[;LaMMIV69
8KF:e[\:4-J+.;.0Rd<7T=[dRYN(6R^+U#U.=4_)AIAb>2D/0XBLVga_H;E_ZHAb
Qa#\C#_OHRf\1.Pe0bYS5NGC-BUE,,+]]\,9L#HZ1U:dEE?eD7I8,P.&]9\V>f=#
:B[U]&P=B6H]Z&>gd^bZ3cU0:1)0F9fdJWZ^I)7D&;H272)(B?J4bLYg<1Q(^QgX
U1Ie#&.[)I8e)06+cb[#,1aXbE<U2IA(KIM+CUaX#)cSMd8Y<fP:G>B(/g8>cRBE
EV-QI=Q<KU+P1f8G;cEAUPAe]IV8)JYMQI+T5NN2+TX\_&.Yc6JB.A.1D4[;\3<e
,ZS]Q&Oaf2CK<QaS92)a>P(R=X19OUDa1[<<Y(VBL6FQABb69Nc<WTcc_R)K+FcY
VfF1U)J=D8?>26]=EQIQ&.^7X\abe-J&S;H\VUAb:^>7.XX+a\<f\PeTJJ=@ZLb?
.;K?X&<X9PYRX\=,;f@&W7a,#&bS-?&\O7<+2W5>0eFbEDad):2?SBEA8;Y]58)C
L&B-+@2F+50,3MB7&W0HF<LM@^A[aQc?e\G@40L<Kc(CH;(XXC:7P=39.f>b2=Y]
-;2[4GGEN_IIPg=NS>-F6)--+QHY]E\<bTHb]?M:72-S0dT4NdECgSg0S_bKO)^:
O_^P=@C,>GPY^c9(MP\,Kc4+O+3TKKV2Hb>D3O3gcD,=\HNAM@G])P-,?\(W@c\R
3dDG/;dX9V\:-2fEX>A[)Zfe3K.d#[/@:KGRS8B#(KLE#Q#fWSBD;1JcUSQ;.94Y
.HN\GV9-_7eRJCO4cgQgB9)MeGLW0:46d5XX:g,\H[M2YWWAY?QO#^@)_)\._()F
P)=+N^0<@dB2\8fVdcc_U:80-2_N87WB_N(B\0e_UJO)Z[XCdb#=A]J1&@4KAF_:
IGc-L_eWG5&CXb18:FZd)A9P=]:Z?(Z^ZMaBA(:-?\+bTA<Zb/)f[Idg,G_^+C^K
10&<(Kb\4b[YI#)>a=3</aJ?D<JV[a>:ODd]cfbSSBL3@9(Mc][1K0,S2([d8\^C
2FLJJQ?c+g3fe3&FP(f-c70-HcC5=0Y<;E:B--_&1eL0<_)^^HAQfMg9/C2FAV,6
=8.U05CRUCH(P;19H:E(8[GM[JAf[BCCcGZGERS91NR7/GAU;C)&KWSVc(XgI-SA
X(R3(Nc>A]:I,#+b]4f;aNXWSB9+CO4c.IFRgebCYSCD],^5>GM>WT6aY7JTTbG2
P=>dR8BV6IQB]=E-=P6D:bKU,IefeZ?4G^d5TDQcMI-BLM[T9Y=HY_/Q8AWW^J=J
:Y)c-ebf:/SJ,MHRVRSV@M8(EYGJ6IICfH[H<L50\2;5YJ82BJ+#DOJ\eg(EJ3UR
F/g@P>>J:0V[eAE0;(I]7C;IZ+U_;/6N-KLU=4?84SN=JV7b^WMPI)\AE7H#K-J@
GXRdb:_N.BO4BW)#ZgXHa5L,XH6LPH/-:ANfe&8VMOG)CZ,,fPYZ3T?>eP=03dc=
>A2d1NT_ZQH+gFRG_=_D2bC5g^deNd4g;&XSDKfR)cEX7&XA6H8TNU<1QEJ:HQ9\
0MHU0b)K0&Lb,3V,.1QLIQ2;(F0:6]/B/cDW7L>5;B7+e=.dR9#COP7)U)W<P/J,
BHCL)KeMPP@N:L@UYB.-)\H,-][_g?.CTIf?<KCe5QV1T>IMFU::&DPP_:?aaUH+
6?)/(GH9EJbLg96MIAAT7)5cFJ[L90X7.4K^Z+JQLUK3;TAVX?#?#EOC>+.,&4Y?
.d)EC;8dWZ(Yb;3SC;BN[g8P#T9gP,WI7L]8SJ@aO-/)fX&UN[)U;#(,/H.6e5X4
);aF9ceL2Q9R_+VY6.)I[LV@T+-IFf=YX,e7>7;E_;_AN\;.-a]-NSU/CWD]3D^#
^FP+&=4(E1SgVSC33;[#W<gVcJ,YM[29W4QECcg88==<eWAXdZ)?V(=)62X>)MJ&
QIC1C;KLAU<6=KZ6\(d07Ub9_@&K>&JbXBeM,DOZ<N@3UF0\<S[1VdTQ?U7>UD>5
1a_MTPN3PV^c#MA0TS1W+J1O<6e&]91b8WGQ#1]QC\N[><VUf:C1+HO]K.58cF1M
(VN2&e?P5(]3^;DL[J#:::FTZ,(J+R-#Q=@OW\<L.CL<OJ</6(]8/#,:;L^\172L
,XB1^[[G54<4T:f,/V3^IT\(LLfE3bbBZQHS3<MQSP6[g;3<=@:DZH3T#RPRL^V-
5FMH(-_C3=_IG+-(b_9L[<BZJW77LAf>3W>O5NH?PBO[(f2^/<G;CQ.JYQIE(JdM
9^+WPdO]&Y/-Ua3^03^:PbO(.6NA<=IA@DAUgD)ZAPE6c-]O<aPb1e82BG=Y6R<a
c<BO=FgECKa65dNO>>=20LM)XD@eA,dgPS^1bdI_S0+OHGD;T3Sa^XJA3,bc).3B
F=B@X4e8X1ENO3a=9ga01OO8IS^HW+22Ib-+dFDA:DdE73<cCW.\b9gFa\RLL?TN
>.Z7=+=+;USP(0@&S;W9BDf((\:bF.<gfJMQ4Re<aASPW+8=KAC/f9,=^OUd@^S0
UL@.#]E5M2H7=ZXYGgKUGd(?35@07&c[;\gLb25,5\&-UFQ\(;#IMZ9Df2gZ;c,P
2cf9C1g]3.HX^D/N&W^6]+QK=W^VF8.2.^OZT9MW)#+4J=X8bGF_CP?B:f+-RSc0
#^_(:5NW7?VeCHa<NbVI#93fSXZ6UdQF&faWSd<7>5AKE(PNC&BZ/QE&_BgS4V[#
NNa\ONQ?X+UHLJ?[=BX12CXK\+OJ7>]S@Z00EB1WV>M3A?DCH:9e]UZe]H#=d1e<
:3<<_R.MGAQ[)b/d15ZN48#W3R2/,@(2]>>1&1V>9QN,F\cQS2f4[IM6?XF.QbH\
<QID5^_[19<)YX3c.TSV([?>YHPSa-b_:OdE6,)]&YL-;f(fSR0NT6(6<?2Ec.#F
VZ)b?YOM.86<bEZ;([?Y]>]((Cc5M[^eD2c)C_(E?g>0<J]b.)YK9VR2_/@?BbO+
1aR>Pb964NW#@+]JCY0\P<TOMVVE\=ZaI+U3<DKg@gD57>8&82ILJKL77dF6JaFg
?P8SF+#T0_CCVb)=dF7;O8_62NSJJ)Fe8eF9S2U(:_4<GM]B_;7)[1c2D<-;_^+3
(AMReZ<7XId7CAMLILb,):1X-Q_eNK(U,/X&b1K2PU@WK\<cXE1A3R,bf;4b_L[/
]d9MU0I6f,53:E\_GSb_RCW9:<9-eYW7;a7Q2TYX1P5;BV48Hc_ZS(K]1;12Q:6U
HP]63=NU+Xe^,3#4JBdW,L5,PGITg9Z051]_-g0K(.+^:/C<)c,<U]VY=#[MFf+^
884/&O.LW&IB6Y74YSDL>eMU9e.Y810JN-Q79)B/0:C#]IF684NF2Z1dO0X,YbgO
9HK/,8ZJ)Sd2CfXNLU7Fd)PS5105X9aAO,H&7d]ZGMC;#QfC]X(-A+]cD)?T_MW:
M0\X_8<IT?X)DJH#&[;Cc5+,=3e[<&CESGH5WJdB0]#TXeD3/)=Q3C,IXRD_^0MD
8&<5X;?0UKU:dYOdMUA^XG0e5N4<,A/OMeBe;aL3HRbHRH>#AUCXS3M/P^RVMgR,
.\;A40Q,>bZU@BU3?:[b5EW5?G>XQ?J#<#D=0PA,XZHZG0RU59#ZONJLT=WZN^ZM
gS+FNCZ.6?^IaS46>I.Wa,cbY4<Q\<982,^2PJ;N3Oc<_6.V/Cb&5G-\6K2H>,U&
+-W9&b:6c7-(V@O-]#NC4H86Sc2UILN.EdI[g90A]LO6(\_a?W.6^=JJcDR[/C5+
R-eN)Jb354N#e6B;^1?[P:(=@Q^<HTZN7>?-=W]0E[?XRR/;g/HJ(/HA3>BaEFb6
Q\c1g8>3BD2?I(K#L;\<4JYd3,7#VIA58VX-D8NNdbK8;+]VdA=O_f\VHe6MdcRF
3]\W;5-@^-M#d&?MF?=:2X.ALJc6/VfW\7Id?NQbZ6Y+Y^:b9JB>Ie\\L09;>+.?
23ICQ_G+-J@^O232VSR:RU&71+V^?P,FcC#_215]_.D)F_@2TCT(/58J2>SJ#/ME
8VA^#L8\:a3SN)L?[2.YKf+PU-aD=[UGfD)@3[a+=<=;)HCURMIVO4]2T^S]9[gF
ZLL)PT23P,aEfB8a?NgUfUQgCPa9EYR,g0^-_]a+Z<5MW1=-JRfE&fHGb&TM:0e8
38-]aKN<?e?E:N/^Q@=.M.XG,>(&+WIY5)9GOf1>D^88;6QDC9=0@G/MXW@[WNMR
f2PGLc,T(Y>CH]_.JKTD)#FeDJ4181RZ6F95g,bK04FeffX36(GS75R85GAB3(#)
85/OH+[ZXGDF/6gHQX\\.RCc\(Q1SE]A_RZbE/0?B#Q]PM7=4YC]ZI\90/&b8.gU
F.Z.DKd5SADPc^,M--Yg^LPD-S>56UCYCM?E0XP4=;aU&3S6<7BXV6&/O_35#T:H
V;DUGgFZ8RTV=)AL;Z^AIMN#adH/+?fMDIDT]NUDg_1H/eX1G<Y,EK1@R6[-:+X#
HVXM11A<NTgW<@3YH<95+2XQ^COY?J649V]Q0,/,Me[dF<eM?T))A\TQ4VOIDZ,1
KMX#Rc.O4^X])P:<JKM_2:dZXGKJN58A6,.RY83\/M;._U[Z6B92D_E@+IeCA>NZ
E8Mdb(g5,F<b-f>7)\4Y8bOf@I-I2?_Z0JQ7W5:J^/<ALbP9<fZ#7O54bNGf#Y_\
S+]1Y;P)S?eW,+,5c:U;I](G;8G#&8YTWbN@cJP8STBXYQ49F>]A:&GZ7<bN-a)A
HV3JcW#:5VPQ=&=T+a?9>c<ZY0:T5)09B1BZ:NIT78DU15g:Z=^7L8d+@d:X+c(S
LKX_R)Z=d+NfebFc839[ZeFFg+0:+>UfJ9RXBC##74N8_@0cLbS7JW4X0[@&+-_H
aV[AeA=(G2M6,[bH<2DJHBY-dOL-G];:3V,-+F/T6+#=G:N.LRW(EeB@KTe1J;XO
[K;(f)VRab9d,C?/WbBHVO21Og7?YU0EeESE&RXd.f,H_)DQba6^H@4T4W4SGBX\
IU[@+[7eR(YOG37PKLSAS@9EJc>/e7ZcX^RC)0+6[2W<;c?=_9ZL3ggVALd1eR>6
FEE:e-?CfQW.F3VAR)Q],B#2XDTc3843(YPA\9TKAWe4\PX@?L,Hf(#1N(?-]-3&
/X>^Z30R06X3RgW^BI-3QS-YdUP8^f22A\Sadg<-<[d;SJH1NcWLK[aMc0M7PKbf
#YfU53V4@Ya\Y?HBEf<65P\>R,-HOZM9Y(]&FZX&D=Oda(P(V//0?SSJ9],,/:P>
UM6.L6b3.edYAf9B&8]9BRb[JR#E=Rc.^72U#?:,JN^C1OI5<]0SQSR?O(B9J/PX
[YH?GHC>U@ILJSDN<eQd&9>gWd(a/ND;5O39(^#(XA#I.:c]R:R#-d0FUJ^<OB5c
A5<P3c?g0:MEMKd6RJBgEAUQ#XW1QI:B3a)dJ^bA60SZdEa47f:8/YWRY9RS)P-F
;NC)FT/b]>(?[(P99,H3TL-aa/]g[A:E,@39(I7Rf@4EKCbIC9T6NN]]&>2<[RZU
+6+]eIC93aa6<cc0JOgTO.gLLZ08,JGX[1ADLb:M,5X)=^5QWCQPLcPT5Y>(K():
>?&[-J0egP>)IS0TB@W-)aYd5U5OX-X]J,M,Dg@3A[C##ObEUXJ_I1Wc9WXW).\#
D:5[087O5dPPaaH5+Me30LT2_)gBgSTZcV)/[SJW8EWV^N66+-+d/3QMFNZ(&TV(
aeDJ+8c;gE2M2B6WEg49(VL^f,&9DOL,]#&KHKIH4e:ZGMdJ;XQ1g-[5;c0NJH?C
-2;+>@:A#[730MH:P#0KQLP?>QQ8#Q<@K3;C^P3&0_T&^5a04#ND>XEPT1a/+\-B
?&V_,#9gK:6OGDB:IEa<:RTZQ?@1(=@\G@\39f?=1<#H#c+UQ2gaf/dBBa9<_<AZ
/cfW@(#:)U&c9IJI/&SZ:7X[Bc;dE,=9dB\ET-L=He[8:]J=+C1fXGW2=FPYba5?
C?SVaf?S/]2&8A79b?4,O/DSZ>/I&?GCZZaMRA:2[BK:)1E:.I[EH^M.PX;_-F]#
H]B&P3H7CAcZ1:2-3/7M)fg]2X064KcR_5ZcPYJ9MHB2a+_/bA8]C7F(^EWXSZ>D
R73<[^@&ZbNNUVP)NW,]OD/gb4eTR/RI>RgV&1:4,Y@_(=8Beb:#&B.[e/F@K?6:
XGY:2=G5_O;Hd-<+dY1OZgg[>5=0;>_>^LF4b/(bD(+]X.)#X;8=Y8X]>E[]@5\:
>N83A+fY0b:4JA88^W=C70_0FCPA6\b;KD-4MRN7=T=MA/N(5#2L)Y6XI#2c3FcB
VK6V13.ZF>7T5c5DLKFS6_.H(8;DV@TGT5<2)\R8U\TJ&R\@SD6d[_4NC#+&X\3b
Ze49\3CCD3f\Gf-fSO5OTS4J,bE8=(V>gG1;V]dUFB-,#.^EG0>]_a&..bA;(XU4
Xf5X.)CLLT?6VLP3g0TO:(TOF96[_V::#H>.Ad8LU<7fA;[H^]TN9Y\R=?[+F)<V
I=QFOc71?BT]NK-;45S3LGT.@N_=IV@Xd^0@f70aP^V<0V?[/^<LZe-Wf/K8D4&T
0H6+[f7#cVF#+]VV&,?#/BPZC6T3c)]d2NK+Z?B#>RT4H3_A^]9.[&F#<U[>O,;1
G#3#bTY?=-_QJS=&d^RQPI17EHf-DF#D0H>E_-^0UG=E#9GM[29UA0XZ=50PB94G
f2B\<H/Z^PTR>-cSa=bQC6XdN7[gH5/,6cI4feb?I23+8P@VF84\>/)O&47A+f1U
0@6b2c@K_QcT\HV_-Ha85+(Q8,4/\CNE<N02[?TBbVI)d,OO,F6>P6BFW^E+BDCF
1WYBAK@cFLOWOO<?Y0aAX;gS@@69R4cR,H?&F3C60dPJ8gXBH5bC.=W<C1Gc<e2C
fG95KN-C8A-B(#[-EIZG6+^5b30<IL@O/8&T)OK&bSe)_O)88PC@S:>92EcZH=<Q
c.-5E<=SHgZ(FKgM5bT7K[GR4Zg[S>8:P;b^0EIO/],IJR5a)Hc09JLTQT96)YY;
:X3S^.+?7C8[&K_87R&>Ag?_I1>AWQbX;3>^e/LC9Od230AS]O,R?fLA=_VF.88K
acJd?MbX6X+2)8[)9RTNA==F74LJ>NDC;&/e8=I.09(O+R\W_P(cVbHCS,MXQg&:
A(D,//J5E,FdE.eZUIHgd3AQO]9C7]78aTeg9=Pa(gaWB&09M//>J<3;Y;VS?TN?
fWI#C0:_UG>g:ZZYdb)BVAQ0[4]B]?OK,GM5WY&)RH.]+Pd##HQX)J+cgfOY,;A]
\V81:4Z?1763cOISG&Mb;^:5;6O<3;IZNGVQN;NSL@F9696(2c):U,(KA[/2<QGL
6RW3K.05ga?:e11^4gH3GLAA1@).bf+091e4/?U#C>]QI25:ZGeX\[@Kf\dJG0MA
RR2dQ^GCX8QPX#QBJ>7c/WUFSMd9OESc@g1^L5))Sf(EMBe,<P10:/_L^QZ6T?eL
gBII_/^3F=OJ\Z0D7g@)S#Cf2^1S\.PT^3bMEV8CI-_C6_bWcU1-WAGM0[)08E<)
SE2A[(:8X-c6Y4?@3N+:,>5@076g;Ge;08_<KFUbS[GUP+F\5b#LNUJU#N-BS3Be
C.._0cBI&LRHESDbR^aL=[=;)PSfTZJO7geQINJ7aD&(+7&aH?/=1Z>I+db[#)X7
O2b-M0MKaM<KeOKK9,;2TU5X=A#R9J79;]3?bcD,R.,8UOTF+PGMQVJ7]E8LD2C2
NH69;;?4Y[BPBRK=G+e<[b/L:DR48/]X-@3<2E0[7]F[N(.D+QR[]ZCM+=56FS4Y
V7.?7<.T,AfOL^<4f(&FB-TSUGL[G16V23MI60Y.TWH=e-QQP5_0#M\Q>UWbc5#)
UfP9g3SA)Q#E=CE-O^I3=+eE\/)P5CF;HPfA)9N8/=+_T.KV#LAf?@BA2S1[Z4XB
X&84V?&e6QXU+9bL5?3a3]ZHW&[@d_GWXb:@2&H.V#:.7](MD-[DCOMH::0VXA0_
@(H=__,f1AJBYZAdM-L;fY6L.C@0VHF5SYL=9^_.M6C2G#5BA)SPC[>;SMCB7IA^
<Ne0@WPO>96-3^d3X@a&<0]HPL><&RWg97YV+EfS(;Qd\RHW8)TCOXUOL0B)L2<U
,f]aSbWOOC1INdUI=a)gGNg/4gIG_LPC>,7W1ZTK.\6\U:Y<NIMddYLW4bBGYJ#W
aDU\/PXPT?4[J:<KM0<Y]Ub@6NT139+c+07b+b>RGU#H8_g.:ZdH2Z[6F@IS;Hd_
eL.G?]P@TH3F1#TP1]8HCAJ(D)>_KB(KRC(@._V<f0SD-@KH1?4OZWXcHE=bgdd6
LdUd2@7+VIUBHPeE.B^N]8.CX7DY53R@fM>[?RTV)]BUcG0>aNVG0AR&B<LHLZXa
.fG+^#[Q;[-_UV9:8)1R><d_TbI^>\LGPUN9]/eS,eQPGbB;N#B/5b0/[1D<0D<b
_I#1,:]B_RZaCY2N&QPFgS0^[8[9).4f,]a_SKQD]=)Z/cWJD>DB?b4,^]>f?FLd
=;])/TD<PKDK[?INK]&+&fc)BAF8cA^[J\/dO=(+TP:e@2>Q[62b,MF=16.:@M_S
;a+1)0,7fa>e\5[H[NXWcM[1^\GQER8WF1+KY?IMXPTd<<RV5Q&Bd#)C_[A0,GRB
>>(>UL(9_A8a\PRV\_fW0Q8=g_,W],(S<4/^[e-1cGKA_6()+e\CXb;S9&<4;/N;
<BI,)(ONYf\L-3faVAV[f8Cg)OaB>M^+E#N\JG)Qd:=3_PODP4ZTE>L3e[b]@?_L
ZCF/@[O4a?KQ44RCF0SW2EG+=EZdNeQOWRQ=f=N=>Q6)&862ZgbJRQ9GE705Pa^4
e9cC.\FgVTUY-Lg_S-8FD8R5=I;;#I4PBZ-Hc(^]A@G&<X54R7a[#2W?5L23S;>S
O(VX8ZO8Ma4D6ef\Yg,CNQV1W9+gJbNO:6YN6_1ZE6NAF/T-H2&&R^@7[]Q@5K+0
QNWc<bc/]H_;H\N4\3aB?N#gJ[+Cb-+JCc7fdF#<HP6&Hc@IU-J6IcH78P#,<PbN
eFY/L[MX[R7e=2-f+Z;Vc4M?d8^7Q)7F2Q(&F,#Va6:a4a6;83F<)XJ9@]YEEL)]
XS7O,Y<@Zb:=/U22N24g]+D@VG[96T\2e/SNCW412AN5\8eIZ7E50EA#LNUF>O9<
.4F>HTHKg97\JXceb,4KcfJY2S4AY+b0#A)^MI(DM,NIJ2C@2fKAJETJ=M4E7#(9
eGIY;cJ,0Q.d.WB]d-@.,:8f>TKBd3\WYe)UGW[Y1>U]DT_U0)3gQG7d;=IPZ3I7
J<eZ7_3+Je1R&DN3D9CZ+<cG^\QgL\=WQ^dXJ6M44DC:9Ia2-.\aGe)E?]+5C/.?
KXc<J^0I#3ODeM<?2P=8]dH0>4Ob>d2KF.a;^b^IPaP6]_;^<3SZ[C)]KVP6K;RB
G:C=<A3GF#ZA7,Z\&H]P[^;B=#be#YT#=FP7HUI)bF?5:9cMP^eaTN\_Z-KV&cQ3
GY;)=C26DTb@O\c;3FeZYQ;:?2?:I+86<B>F#g0-JOZ.W)\UU;&]^:X/J26P0&YN
<HQ&-2OeM-YdFN(U1OJ@X0OU](&S4C3b5Rb\<Z;2^:V0N;+2;V)8=3U&J>@+cQ,W
-,=QYVXg)9:ScUDX)\N<0FBd0e4MJLV5ZBFHWAK(QT)9I2[G5CUKEGS:^fUV^CU9
N7XP+YbD8<])N4LI#^@Paf<-aC.gY7+F6[(G^/@/0D;gUF56<b1+\(4g5VfJ86bF
c8c]K4.:QZd=)M5gH[>2\/XFZJF4S+M1K2]9KfHJ#YdeL=0ZaG(0SRFY]8G,@;7T
(Z?aDG/TG9RO[Rdb1G^5<?-6SSH)-Gf##XVF/?X9/a_W]d00YJa/\M11H3U@YL2+
.1I/e9b?,WM+bP8PJe/,EP4[_:2e?S_@Sc6,IL?^X9Q=JTOAF=;WI,F#0TLe7D>_
>7AJNTOdNP8)^SGP72Oe#Pg/DK3Ga94aJ,5fZ8Z7+CZ4YfbII^]?P.g&0^QD,0=R
QO[7#&a:cE>>g,MHNf&P5XIdP@(RRf3R?53W0caGR\NBb,Wfd1N9c?=gERedcXOG
<EMB.U,VJ_6:V,eeRO(0cZQCWHaQ?@#IY1J>^75C08@XT5dJd)0TW10R]/9.M?;>
eHdA<(MUKL)TV#-R7/If0LdQbZ73)+Y,I(27f#^g<>97J@#8d>^TMgV^0_UMBS7D
)(&/2J9#08,=P?]5B\cQDKT2(^]HQG&I@88H/<56?V.Q<U@RL4;:cC@K9eUW@-8A
NA:.c((6WGN90V;?>.1_GV1]NJ0COTW>7Ae(<BKJ+S5X0dJ#F5Je2ZRDUL;a)==B
cNd5LTX]JbeAJc251@eL7AJ&=;#HZ_CE>UM4->;[CEMaQ[L;WY\#@B<^eQX\XMD2
K[WRbgL\HbW7)NOWJ&P3XVb[.5P/Sf(C8=BIWfUCV3Cg3fW;e8^],H_DA@L;SK64
Y9bf7fK_;QWeEWY^ZZA6C8RZ#bM^)CQHU:-&M_\3IHP^IV#c[_;O]==8X[:YfVJ@
Ofe5DEK+K7>eUP+I2B-fG6MEM4T.M9BH#WHaD@R0VPE02f]CZSaP30S^b3R]d:/&
V=/S)[a_dD-7;L031/V/YDGcR8./QP#-LH4Ha\2^X(]d3THCe1_-?490MOMU<S>2
9T2T=(1A@DJCPBUDaVGYH8OT@ZaH\dL@AM.K-9U]=O@#]/D#M;S6LVXFF_8+-XNS
U[J(U@E,@gI(C?L8)ba6BO<L9@EE8OK(UHH)?XOEC[4MR0(ROM?C>8L>#&aX+OdC
+gK5=ON(+V:P)P@I]W8a_Z?CLDcCcTg5]-B-\bVDY&JP/P[LPI/dH]ffZ9@gZagV
7_6\dNOf88;?VH9KW.[,WF\A8U?RU3)-N+9TTY@UF?#C@gVXAL<Vc&,WO8U6W#8J
Ud..DLP62LV,PALc:X=J:8+S0/dbDXC7YO4/O42YO3QIYJ[M#OWN-eW]D9DV)[Eb
?JI.9JdG7/KA(&T(@EYf^)2SQT(Pc.SXdKM54\XXN.Pc<2GR/UJ\YDE=\8cDOVVO
O:Yg1JP<MA(9US[3:Y/VQg/IVNC=KVUADT9/H@U)5egf/6/B-cK5TbND;FU@ND]/
F&TVV)_>W.f#?X8(WX3=LP1d,[7>]40)[feLA9C]JCC4ZVDH((4@G^2^4H.X)Sf7
AP>,c3cDQ4^U.403EJ@e;gBM#)Gg=e6S,:eg0]?3\0=FJT5T4fZ_,2^b/DVG>_MU
,#87c##C\PGZ3G<CG<;J/Pg^a453gT>3fC-f6<B^W\8d(-@BNdY<\gZ#SBH[gEPb
#D3?^=)L7^2-OAg]E,3S\Y1[N4FI:_H)JB)RZC+Acca9e]<0g:FAH+/KCgJ38K2C
Z<Vg[P)Ic]acDXe@T);^);PE4LGT(Y+Qf:[EKgOI(W4/\]0FUU:/]SVM?g]#TRAI
a1+eA/,>C0_:C:Q)1(:a2/Oe+K)CLG(.b\9POCPMU)SV00g=T/d0NAbIRB=U[_\S
2QfZ/B.7LRFQa;E@060+0EBNMFZ-UHE&&EdPD4-eBSZ>c7:Jg.FKB)AfIEA\J7(M
@GNTg0[+ePGb(a]C,A)&\XHN7028?dE^YQRg@W.f;R=b)?K:QKB>I-ZXgN3DKF-X
_8629a<@V&b5-4Y<Q:]CPDI+H&WL(20^g9f,_H0gf3QI?5H,>A:[Q\;(..JV6\Y1
=Mf=Ec2cK8f54)P:)J=(M^LK6@cQVUWLbRVcO0IBMI(JCEVdF8D8NbEC-T]KP2Y]
,3#:J:]^cEfI.BFZ=)^8N+J=3R?cZ,PIc<IG<f)/T]45>^-XP)R<XAOMJ<U1fNd8
^7M=HSB>]YP_[U,7caZdUQ[8Lg3JXe32#?6L\fE^a8S#G,]+FPS=A/.Y5bLcg(GE
D5/)ABGQP(Jb[J2LGVC.<+UceZ-4]-\@89#g/Q]+;^<1W189[&M9IWQBP,L2OHS=
Q8370D_T+K\4&F^g)f)3b@COVUZaB<;L124V];<(G]I#^=D]Rf^[D;1g[>fJeE#=
#1NJfAM<Ce\]7YFZ/6D\G,S6a0S_aIB4?Gg.Eag;AK<-<d]I_L6OU[\ZMKZ),TQ[
baUgD++<CWA3Jc6gET>)8,JFc8g=4^b5fFZScT_DLA#SVgf+^g@0EVXFIGCG;1Z(
25K1fQ_#c^15]?K-T5[_Id4&&]MK&TaU])RL=C)EQ)YH\c:0A5ge+J>PQ9,WYV>e
1)Y;+D#[#Tb&@\L:Gb(:J91EK2OEaHT[)XK=KCa733F.8-L\:7^9N\.&g1NV1>Tg
3V2.[L;_BZfTD@S[=C4X6c\/>XK87X)(CaI#X[)&fJed0EU)A,X53dAe=OA5B.GD
)>;:B0IZa0N]W^3>VVY)KMK7LBJ-U?PK9K2=JZ(+#e9N45A66(:2a^cQVfeMS80T
1TW]^MSUK+1;/PL1>M2Y0b9a/7HV[91c]-A@2ESRb.V])Y,TR3fgTK\BZbg9E-_G
L#OZW,V5PW:_Ob]T5B=_.FV[NN#G+COggBa6:b#a#a/JVf1[II1cHA\V@#D(OT;F
(&20:Y+5^=ONP&fI[BHHR;51NN:CNH\2R_-QQ7F[6f:)fcDWcNF>(XR(T<33_ZDC
Hb7>PK31g?LD-<&3N>(=4OO)2JcWJX<S4;BRSg,YLL7C])M3^/Qg]I3YH2UR\C+1
VL,Dg9>F6NK87fP/O=ObDJP&R10KZa1]Z5D&/Y+R9J[@SUJ[=a6&X2W<^7&WLL4L
#M[@Cg)f^PM9,7=YC87=16TE5)C6Z.YCF\+GP?HY.BdPY)P-[H5RA\U+=;Y<[E;H
#\7W8E:,?1.#JWG.#9>&/Y(FfUP.=0()ZE>>QVS)/40@STg8a#-KfdLMRO0?b&.7
>0YWH=3LE;5#[MH6-b;d,LFF#1d]OE:b\.OKf&HJOC<FVR[AS)SVU]]cb;;cUc_1
5Z;KK8.?SGa(@DIGVMG2-FE1N(@f7FLIb=7WT>0V,4U?YV0GHIgXWaR</e#9P^GQ
=dB:g___aefJI2)eOIHHV^#V&)@^E:4:dKZ>TLUOE7GOX^57V#(866g[>RHF7GAT
4#JcKLUc3M1dPI=RK1B3<4]6_B-=D-6@,?F<-Sb6,CNE.=<4];DIMQ+&2G^D#gS+
beVQ3R^KHed3QfNESb+8eJ0[DU3D1a2N]3Z##\8)?W4CK0Y7&J5^A)12JZ_Z^=b:
9@XEIO1>#WVMHYPeBE;J+W@GPHSEM?CD/0RX<&]AF8>Jd:XdJPS5L(_#gdXgHJEa
H-[94Y=J?YaFRbE_[QY)VA8\DD8dccRNY4Y=]2AJRU1bG<S@d<JCRP05#eS0a1,W
Z7TX>ad&@9f=VUUUD(W^/&>S6OMg\)J6.HLN#TZ3(N;6dYe[93]>8?+EPEf5DP9b
Y&4+0BC._,^J.@]gD:IRJYGWf9EPE(M-JH)ZA1=YbaWNaUeTDBe5_eX:L>9=VTN<
T,Y<;Q7Wg6&G(9PDaEd^/@6g2bLGX.VN=V3gK_E00fF#@<]:0G+fYU&4C@V0gFWb
Q9?e;<3aZ3^Sg1&J=<4c]MI7))F25aXQK\]?1LB<9D]);O9YM40]fO>e?J<@6PTC
E50,I(SQ)AT(P6W^>4Y>Wf)Z7)/3+CcY5V2G[U9F\3f^7aXEaFL]&bTGD<>V0J(7
4WF.6ND2)Hd<SX/b?,bF8,UU9OEBf^C=ab&:=DW/.]K3MZ/>/XdAb>fS3c9?c2MH
Y>YRgaV[WC3SUSVa[M(77ISWO.6FgD:#VT+e9-Z;)?dJ(,a[]SRgbK-4^56I.#?3
2=^F#LY46KK?22-D:(G76T]d&YP/=W/bdPf,b)(KE7&1YBH&H7773WL3b/<]J^L0
D.Fa4K+]NA@ReJM[\_/66adWKBf[>eVgP[H#\H>:?f&(5FL:C1)\<\<.7bDc;Y?J
HH?,UTOCA0GO-UAg?aMXWa47_SK4-F.9>V0-G(&&f:7G3eDD2L]-:/;cc3@0Y7RY
]8\7#.FA4NX-1gF<=eMU3OI6?]E6ZA9X]K&-);;Y@gV1Mf/6OPIY.(.dc[/I?LS,
.FLb#d<ddaYW,5&\-GVRPVU-AFD./+_E@910&\\g17\([<4BH_CRc+aJ.4]D3#Dd
9E9\FH_6>Qd^BP:V9>092[_COXOVfc9A@<:OILZ(3.W&\<A3GWIUKP29#8;9F4FA
1K1B9CWQ3D0d?K:QABc_P)RR@EV<+/.EUHY.:7f3BQ0V:f\OO?/297+]e[YF.FeQ
8Q-&+W-K4B@Q)A^KO_1VZF;QET;R0TJTU1(J?]JI#e6+JJFXE_7^=X,N.205QbEA
GL8SXU=-G.<>cc@+KNF6<?d)-ZeYUf.@P=#Jc(JFR6::8Q,1Se007_NQB4aQS\ZJ
1P^2_58b^C/_3@(Zg2E;P@gGXVg)e9,EM\77>5ZgG;H6JK93HXD2(3:/@Z6I\JHa
PTMb9,ca56QQMJOG1)_<E[2\ccKY8BP9LcORf)CFAWN043:+c=9^CY25c/]]8<aU
B@fdYS07GTYd@>,,M;+GD_REJKG+]E=;_<T.Na?PcH2U1D5,aT+=\:NKc0&(b#7\
N:#=<_;^J>J\74MAe9\&1bP@L#G^Z.;B,R2L8?Y?U57/]RI.H5<&+[LV;14?EGAL
3<aWBN:,#fbB?4B79e_,V@7[dV9R>&dJWVTP^T##g^-5X2BTgcZPe43S>0_5-^27
84#:>NQRT].W09:.])A68A5C<_=DQ)V8<S?M+](G\+.Lf^:B)>P>5Y6ZSd?E7_=E
b8D78F7N_VT6cF)U5dPP67b)L5/_ZJ8[UdRO4:^XW8RdM21D4cXD9f>/6dWAFdFf
_7ZbY2C(FVaWfAVD&_<J84LGK0+(deFaf2eVbZ<E.S,0dQ@8A&ZM#TeLYJXf8M[M
/XN7bQM^Q4:[>c@[QQ[-c5bVC/RY_3R=A_3S@]PLU#d\+0T7>?]dT7?PV)a&=ZL3
V)K;]d)2O]L<]\?U[TNMP4>PdO23J)[S[MNc6[M]Y=].Q=RH>?H<\:R@6V<O>FfU
ZKJ64[R9dK.&]+81UH&#dSY=PZ+RHf^WIU@V?Ke:NfZN>4.fAQPO<?@.W<XPKQ_K
dOe7HFe-?FG=^G1;&??\7>J2U)(C7#L)D+8-8OJ:\B08<4M6.WD\cKfe-LcO.GS5
2Q/.N7eD2gS<HMS=JPbM[NM/gP6JaCdeX;fSB&?2OU3V\LISZ4]ZS279GO,+12XC
,0O2eE^U>T,bND8+0ag21R-#[-&XLZNEJB@)_P:N\#=H1T+IT03:N&&L^:Ec+GD(
U#,=#RD>^ce->L/1BccK3&a;IWW-.@CY:4dRQTfOd7[@.fA3H.NMHTC7<X8(\L]^
f3&[[YLV<S)8dLL)BBTP3B.)A6A>B3H72)BK1<gU:2]&01=^7+NeZ^0C6CL_+Q^E
8POJ]0N(?B]7L0SN>\FQ2Sg+-57V5^20T2_[Qg1O5_?+]NJYGS8B5W&KSc#c,eIC
-eQE@T&06418IS5=X[=?U+RXCV?g0MXI6VS4RZ^0A5,[;5#cN._R:52Y+9dXC12W
@@S(IGP9X41-MV_R)PR>B#fZ7ISE;FA52<e[0>.UMWS<G\1I,D\P<C;6J/G9:P/]
41D6CgP&=RKU&+FB,4YfQZ>&6/K)YF+aW=VZEM>HX@.[3ZZ(#[Z))VgWATO5RU^K
D6bYB,)4QXSfVVXCPd6TZK[I(K#0TA4c_@V/A7c==1AXD#YB)b,Lf_5H?Q_<2_Z6
-RY)\X95g-N#/Q5Z\;I-BJML/5?WKB)^KA9O/Ze671^H>CYOacE(X^0&80If&P,T
-EJ3+#J^O_VA<^Z>790C=LP]IJPcIPP4:_Q#Gf\^>0JB<M7-AFf_6e&]?6REdFZ\
acV&UV[gWe6FN5?e<XI[_Ifb06OI8Q<W>BObQPQ8:L(F[UZ;>XFHb9B0)^PXW<VT
@\Z-;,2-JKN=<a=MS&d4?2@A#Z9Vc(bZ/e>Vde8VDDM9I(3W];R-^IRQ--W<(efI
LG\V\D]a0OQ:27#&SW@80c\P\&P]B)\I00K#.,Y-^\S<Vg9VICa[RS9<-Wd6-\_:
_03^@aMef_PIW+H7a-P7)4&4,6Z-4f0;K2^N0/P^14]=6]cT\F_B@f,(,(1F/72P
)7<I7_-9>#-#XC17RBHORRB;+R:F#b0V:_@-AULPM]Z?G9\#&Y?@Ye]=&[Z>,g#7
Q,G3D-7aT.0KRRSN[Ve(RW7];9(BI_\QQd/W=f9[<a/O3DZOgVP.[^.6:]IO6?X:
12@aJIb3#8PNM[dS8D9K?6WU.&T3N+QaL>KRb)KR]6QOR+^M_#c+MB/#?6MQ+\4F
c_63:fVAULX0G6OGS[\PP;JDO7H/S3-[OF>BRYF;L5&S37R7&&0&d:LbfR6(Y]a(
0UL[@=6(Zdd8D#Z&IQ,7]OZ@Z/-J?FC.[0:V.)CDU,fP9HV/Na:/QC@b+eb=Q3B-
P2+)LILUJT4#=#)A4+?Y,1O[<^8D[NW_@P]?[>a,:O5^O.REb/.ccDQD26\[7E9[
&\e3,UfU;GFSQ@&\^0A:5@#=F8,(._V;-VW;bIZf@Ef?[X>fZRH7cagg3Q.DHGTB
X8&DCR9VdgSdGG.dU://J.BH4:E=E1IH6W/9KC@6_R5:c.-9NAU1ef>[-Q^;8\-B
D#KA/<&PG;Y7([)NC=-/VbP+Q,-27X^)J/#-&gDe9A4@,@MDJgE0XfDab:gIY;BI
#gPH)7fGa288ZDSe3^+:?FZgaZLV+F+(N+A+44E\]R^Sd>V,6>bgZU0<MO_?ZZc>
>/V(_#(V(J8)F\,H4eV<48=OA]b[;,6S(4QNYZV+-9;[Y.a8[7gM:[D0Y?b(RR+?
6IVcXCb??MH8NJDWI>cVd?-V[C4F3RD2(EfaD;>72MK9>STGC@bZ5X1VT4W8-,/O
I\#W.ZZcYQ<e24dCF-2;W0BI60&7X?N9_OTMc;;gI&JKXYFYC[SLd35PPc9Z7AYR
Vd>[I>6e7@A?7QKV:d)GIM/-cM,1^Megg6RUccSY]NP3OP<N6TaX[M7TWL-_4]>E
WXRUD:.[e>]@e\A1B(NPOEHW8g],-C3>,aI)PR&<L4J]LUc5dI4QNG.?IV,b>HAO
XI;S4?)_a&HT[L(^QP6@G7JRLD#(SY7=-/Y9^]S#2[d,;=1.d:[V<W[X7)MMD92V
=:e:(7aNZ^[NCCJT)2EFTY/J5U\?58ZS<@V_0\([MU3Xac=0]WZCMFd<&Md/Y2]7
XO@3#8B/UV5gS5GPaH>fd56D&CEL04?MZS5KK2_KCCS30O,\K5Oa+5GBH2/AJB-4
BTS7CXH=R@^HfUBI\a30;_#2?J,bN5O&BEe+1;#3UB[f8?H4/2R2#2Fg2?O:K7B#
g_DOH<9C5?O1F<-GE?CK6b;M;EOJ]Y2Mc6JNR4P5AZ_)&VO[f.WBIZB,S?R&U841
>Se4MD_H2N;)JR]b]]S&Z+306&cXOY?QON>@GH?515/ge.@D]BNe<G;(#5.@4?\U
#Z0HC/B<g>8=>H-]f[MI?0\eKf=.4fcaGK=Q>ZEN/X(9SU]3gBNUWdYU=4GF5&,S
K.F[J(b.1(<,,7@3..T8+Z?bB==(d>8C#88eG1e4T,W4N=RT4#R]DaCdeU2,9V[C
I@CJ_CZI_VZ,9@5\[^^<bL7Wc_<7^<9Z:\RY0I#>WG;Y?,((MAF)VN^/)PR,E?EM
,C-^I/NV[+WCF)g<AY&H4H(PXHPUBQ#E7-C;dC[>ga3WCC3AQd@-GEY+>XaZ>+P\
)]e19Gd8Q@L/eSN.7ASE/7BDX[BbH&\GDM4D0C@8?;#(<\^f:(ZNDQ1B=^:G<E:.
0.)K&)GR;5;3I\/&@aKa:I4bHB.U3DWTL.\BJTT-0--;WK^-_Wg[d.^Id&?.gM/N
J7+UJcbL3-J/),PJ9-7g(/./d+1<.4-4F_\BW^2Xb[8aXD6VED<](CF6VJ(Y@P9@
5dSMa\J.gRNIIHNVF70U_gb^1O=BSR1BF;M,U3BUKQM\O@c>d;^PUXV[&QeKVNIf
[c&5(2.N(FA5LR/K#I_PB8#M(Gg&DHEBQF=CD--J3TfJaW:R:3)96#HYb3/-;5H&
#(VIe=(THb@=fKE(]ZHGdDU(7<MGD9.(WN>CWcK--Bd:VEGRCY9/LD[O?2Z(7J>T
H@(.FBDY^g-4gcG&T_GTbO#.4QU3Z4?+fe/b16c0)YfaEB[]\2gNaOdO6&,INe:9
,\<W)V[0[M4,bQ4QC0+,)IJP(X]>PTZ8><Rc@?_7AWLR_(I_#Bc3/H2CI&60@18J
GJE4c6@2(c]^bMV[5P_O^f-NY54B\V&8CYUg(W>baKD6b[-<ENFTP26Bg?aWX=Pe
=Q)P=8F+^K]FRPV=A(7,/Q82#-a1e+PO_eTWW&#([86@AO6IMRaJ#77VP\GULDV4
_?AaPMZRd)1X-[/7V@QN9E\:?/JF:0g]a#cCfaRT@J6C?7G7aX,(L>,]HIC9\]KE
@5e9F?6>,<E/Qd1c(,)V_&:Dd4fVES/8^YY2O9\G<QBY2R+5&30SMZQHeLG1A+<-
:U@#=>B^-:]7GX<&H))a?Aeb#]M:T8D]F;dEQQTcD1eNIb]FST+ZQ\>^FHR.e[<f
>9G09+\UY-Wa@?+de&6<B>AD(MVLN.;b&Jg]MS;R]6A<RR</g+W.<Ug^D+PY4EWb
1YEJH<T]./C/Q1OE))5Sc&a.+ST\E59ZbXJPN]Z.X6]d8.JW/e(SeK.MWU3aQU2\
g-.P[E2.GR:36B_D@FLU5G+I.>2E.Q&L^;dW[9FP+]<PDIT:]:.Z/4Z4OJG0T8/<
[=@21VfE[=7(54Y+bGBd68gCL6(CJ0&c++Y3T-EW/.=OX8/<TUQ\H2\M+3#Q)Vf6
gMN0NP-0_WW+Q;Ff873-,0E?PCJ<T)AX.[02)O.WA5\OHAf96K[OP5Ae4PI?;(\-
^2T5YaTI\4Ze4#gT#8Q<T(XKMH#T9S8HdK1VD73;(>E(UWY[/MH.;,KcRKL<Od00
.7;QRR,TYZM@QFe53<eg8#6f,K>JG;.OEeIXe.dINX7ZLA>cJRR?9#VMdI5]<5Z[
;>\ggcW7=_NS4MY7Ec&K36_a2U(^Xcd]7#.P3NI]D]9SC]EfTR3+73<_,U,R:+[Y
:SLQTETAN:46@,AXO>-B[R,_NEMcU4a9=gc(KVO_9UWJ-YG8_;ABX@3FGZ;_80@0
;feK,JP7:K6F6\07;Y3:3+/1V3R+8J24]c+MFQLQf,@]2)gC\2.(&\F8/)dWD64Q
CIJ7X:<:;Q0S=d4(-[f7_PO.O[gcF+d(J]189RaDcF=\BKHJRMN&BKWC@&g(RP/8
d6cRB?M,J)67HGR=H+9a-aEW9<ag_R==T9WBRUZ_;<A8;_f+01?M+c;6DXVH//gg
MFD2g2#-&_)6:cPM]/b]B?\U@7FX[DG=[JeR.J?AX_.).N=<6]D=8(dJf_21Q[IU
[?#5BAU#R@R@LT0?aB#M1+I?>7baA-CV7^ARd_E?\Y.M7[c1fUQVE)?Y5YgAF[I1
,+3T[O/)O42L->K?We<0(MR:Rf44CG2_=A_Pc[0/(#;?JL34#V#V;P1H/CNG&G7^
U^a+I=5NNUXe4F.ZWV0B0Z1F(T&ZJTV]e=;THHQR_,9>V73,U6BbeLGQQ.d3gOTK
-7:;^8K<,6WKX2?FQ[I13VIBF9\V9RH:_7XBCT30&>XG?9\3e6U>f5/aI-FFE9VG
E,AB.D,PJ&)(GNQKN]6Jg)HW0aCZg)H203f\>WbE0>b]BI-9XN-Zf#SWPNR,1P(;
--W=0M-Nf3<Z<E-DI.C<I+I[9]?CC05;8-#UAfbV2(8NcPQGBZfMWA4HU-&H68aH
+:2KW\H]]/Z<WUc2_D\&GIF\ZC&,)T24[SKRDYU1aP?<B4DXfP_,Je.eE8<?GO@Y
RX]YEL4:.2\eR[a87WJ@&=VZJ3)OO0:JF5ZT;e2[Q,^W@DJ9&f/6V@7T^#OU75;U
Ha-ROe;@--8f<).&NNSV\-<P_A0L5Yg,I:A8BVK&;:S41F(7?NS.1J-H-@^9\W>)
-f@E4C0=AWdEGK\d.+g.KQKFGeaT/Q>HQ7Z>3U7,ZN/Y#KW?A/XWBeA.e)>BPdTO
^_OJ@eAU]GNAaO^3eT8+9ZQ@:P1B<LcfJBRZQd^)&3g=UX]DA:\I6X7U[LKN,@9P
7H3\/CP:SITD+W((a-W<UdEH\50HMKR/^D5,C;O;_NW_g[Id/7BW8LJD5Y.YbaGP
[XNe8>]ZJ:N];+C3NV@Dc^]b@S]VQb#=NO;P^)&-^GQAeB3B<9^/\;)Hb,-S1KcP
+8/I@U23X)L98PKAI]a6:N<QG]V/>ACIAC</9)P_e)B9VH19.5(Vd+Gf6dfZ8S3<
F0;-,]b_H_ZeE/5RVDLdgRF)MI8R;a>7,QR=JQ8IZ41eIZ,Y@F\RfTYeR30E-+5<
)QV(S:-g5R.Oc^g)^\e745QUd<+X(\D<GQ7M>bC>U0@#2IV(I__XG9T4R)Zf>Qg9
K+cDVD?6AGL=#@XCL9[]Z<LBX-d(EPXR)FPU^047E<03d3<6_(URJ#3E8J8WQW3/
,93Qe)g-?Af-^A;:2=M6M?6d;,baS=0U+?U,DPU@L)C[5)W&LZ@6de6X=2ZJ<[K]
:D.O;..G]JQMROU?85M?JCTV3YLaJKa.O6+0KN]bc^[.;D[M?6.EWPcCfHN3f3O3
cd=cBZ)@^M98J3I);;;XG7N?N;b0eGI:e=Ogc]F9>e_XFEL.-X2Q35F&XH:85^O(
60+FYRUVfZdF.RaPFP^DQ51dGYOYTMTX4f0CV:8IG;H/9Y4RL>9A(X@gf(5<6Q#8
>9GNE?B6.)g.Ye/Dd5Xf6W[d(e1gAd3W;cV(bZce:)8]>]2(T9b.TQKF:-\:fbQM
f4M3=VI\Sc]b=^K2g7IUE,XVYC8LRT2X5]KIYE^2\-,QR8dACQf7ZVJ_Y;Q9/\Y)
?00cBC\OPN&QHc\>V7S_MB5^FLS[M\-NC90F3Y#(G.&D>I2XWdN/.VS;Ud(aa3@H
.G/Me7KP;FXbMT4f]-+P]8FI-Zg37HV@]#TD;HW+=UPGf/ec2dcb9&]/WTb-BZ.5
:HX87/KZ1(LW.C8A9X?c;Sd,BfI2//KdcgTaC1RULE3PO&50@/:&\<]_G<VJ2-8G
ZM0c/0VcH)RFZ,.N=c93J[bgg1;P2fN;O.d@)5N\(EIV/26)gWF+K7PXB.J>>&)<
eGdF[aP\31JE[Fd+NG-<Ub)&_WKF/W;HeCREMEeR.KB-<I]3\=RD>O]NF3\e[^AO
f3CG@+]H+cB(:9AOIBU]=cS0&K>RI[7BFL8FeV)PV(0WZ,()NX6VEMGHC4M2eP^N
P/\7H4@aU02CL>6TCH,MG66>WF2>BJ6,FbP=G,<)D,7DbZ]O7aYBO6g?4&P0J?NI
a=W]<e2K4&(\/^U3<8YDFYa][AQGg\,9;F-8<9[g^]==RWFF@H[d2=Pa2H-1MO^,
bBQMTb-\<7BS<U[[+V/.fQR;O9b0e>]7@HF7<FY_4JG\g/Z,SF3\)b9;M6I;0L(E
;@FY(:V^=f_+L(d,HAcb;1#I6CCeaAX=@.H8>IB3-Ae=];9:1#\8W]b]YJ;)H>:-
5WD)3Lac]MbY/EE5:69=-Z2#aEb8G?=^J._R[CV<.6,=H&ANURSJJ3VR0P?JMfd6
<#\6bS=[4&BL@M2d+,A89b(G:4JYFHX.#4(@R\>e(9EA/R[YQE;/beISN3a5_c<Y
8LbG3(:+<:)NADcdZV.\FTJRGV9B:(5F925CYZ]E)YG^;=(R#]f+7C+>5AL=(,)L
+L>4)SM8d9-I>N.eKJW__;6Z)M3)D;+<T3b/ZKeb9@c>[SKPYBYSCC2YPF08^28]
(Q0JDIQKA@018F?+S@-c[_?5c-U773BWCb3<.,N7E95@T)]NDW<T+e\SFFFc@RRb
ZcZ+Y\ZDg0N:OcEcF[^d[+)W(^R8DG_f&213[H^_0_,NaQOONbb-I4VcN=)2;8.9
O8?60WPb<cJg[JVA2&Mb^LS4\=dN42JT6-7J9TM>,^ab:C+@=VY04SOT]KL..0Z(
[HE.A5U4,VNaXY@6=Qb:JR::X&E^LIGYKf^,9SA+0YNMbATQcWJHd6E:Oc?OC:F\
NOBX1C]2D4/.M2aR)VOFd.9\eRD4W2+6,f)&,1)1DF)53M;&]c;28OW0T9(U8J<B
8U)>KKY94a1fH<:-8PG-?_:.B0WLJ&c2:A6b;eDPd[MO/_8cP4V>1MNHbO[KDJ=6
]MYc<b//XL:ZJcI,4gZ9d34?QYIX0Y;,\?\G3\Z6]#N]#5B;BSBO=2]dQNQA4I@4
)9Q/YZ=A5[\5&ae5(P160KL_L;_?g,6Lg]@eY-J9X]>V/^/PIPX7DQMQ7E:bK^1I
X=[O^5=G.(fM8dYI/Y<W?a5BKETQF/K:O=2ZKFZ;?[00RWM)bfM]aZ0D>@CG1AO@
@G<OX\a8D)CYJFLN5ZC[JaH/gR5<.J0b&T9FMP=aT?g]fN:&5Eb,DR+A>V#IC)dU
PP0\W?F1=J;=\J:d;P_1a7W1KS0Z?AGAULM_7Y8NKL0.VbRc3)MWSd9Wf]/Xf03T
dM\LeC]Me.4&R5C)A0^,ECRS)4Q(DKLe//QT->L)06cWYA_73[.H)6?H646K/)ZY
fJJX)R5J=I(32.4XUaf.)b+[K;F]B44E:OeVZ6LeCe;3AQE0,Y/X>))5HQJBEJHO
\[;Me#;PLR)a-SR;21fe.Q+AeF59/?^ZRXL]d#SPBX?CZ.Fe[Jd<:M&Ja>\QHDV5
6/W,=#;6OQ,RW?3]B,UX/V_bDIK&=\>>43d0WHRd?+Q6_:;D&DB]4GM)AS3?R@-?
KIG6OEO-M]69Y6FZcRJVPR-Z#T-]W45NgQSX0:_CV3K;XJ0^Ae-+[;(#1VYZcEOP
cgSY?:<#68fc53aGADRT1.X9@#6X&9+Ug1dB3WcVf@dJKgU^,6DV3eAd[.M)LM0T
B)+H^LJI0M=4-;4OCF];44d0,^K6#?US<01=NL/V@B[)f:9/P&DQ6M:.L)J+(GF>
be4Q3@H37PWeO7eV(DXcDB@+>K(0\OY73.]b&3_KR_O1,HCR34=S=8B4?Ked#Jeb
TgU(.LbfLQKQ:\f#e7?>U8H<=>PcWa0VI@][LO93X7CD.JZ&KTWZJ-X=aNN(@Vb<
]c/A\D.c,)(AO?bIDG]JD&bP7\>G2F-QeRAYNSTX#?K?aaAD[dF2E/WJ#8S7d>]/
.7b?HK_@fHZ:7.D5.fR>-=7O&UN;3)YB]gIdcGMR;MYd)X_0/Q[J^)02f\9;USH5
[&^YePBJQIIQbZ[M+GPe3A\D<X^R^aKf62Z.0MROR,N1U1ID;TU?f(MRY]bg5Ye?
TYU^DPT4.6Y^&\I-I#^gK41(>N2dNVf0_&aDRdFMgX=E15&Ne_]LX[bbX+O>?SUF
f_gTcJ:ac)=[-BZ,OXM].VG&ZIF8NOV^9fC88gTdaWACY>X5YDd8Ed+@ADe5L1>g
=]Yc9VN5N=>dVf<:M?YDA+:VdD@BQ:B_JH66]ge8eR/+-cQ\2dG;D5dG8e1/B6YG
^^g2=MG:TB8^Y?S)NS.Q#1QA4IeDPeWcBf4C1ZRbbNH+)#C=0A;bR7DG3<?;5C5b
aIY2=-Y,&#O?>0]9CF7T\N#(CP[6?<G5e0:T(W5Q<3SL388d_ZgJZb9+-f_@=850
8E1e,L_/#@HLV-ON.Q[bR6[411EEH-5A3ROa=Oc_+H8,)9V[MgAQ/If6QPBFg\fd
8NU94O[>[5KYP8I>#K@2<^261F1CI=[Z(.)27Z,H7PH419<1Kg=<M0ba;;+-2QDc
7PTGYP&;_fcY0$
`endprotected

`protected
(b/0@.c/<K(&Y/?_S_0T?&:Y-#aO,_,R+#bN_F7@EC15T\OL&<)&0)/P8)gXVTg)
1^.;]@/Md2e&.$
`endprotected

//vcs_lic_vip_protect
  `protected
ccO5+0a;?1__3<+.fTET\18\c^A\M/Ld(WLcDF8b\GX=+HB9@>PD((\-9;HIFgPY
NX2V>57Fab93+?SPA=C(gR461G]U/,0I5@RR,3LPQX->+Z(8M\0BDF/-<.dc<YG^
g\UC3R6\dK7TWQRZ/:@QZX+^R:ELK&Mg18(Lg)\)aED2X^e=KRcU/9QH(Z9GbVD?
:(HE;f^3IJK);[:),gfVc02a22.Da:Q;G5ZIaW>5F,D[MbPT;g4dUI,J6-^dFW-#
/TB^c993XPLd;=4(/_7#;.<7QIGI::CW3P>Ad242D-GCZ1=[Ga/.bYENHX4ZGA=&
bX#gFC=L[9(:B0P_2ESXeMa_1O7&OT/a>I05/c(a2@Ed4--5M+MfE+[A?,LYX4Fb
BS@;<IF3M@#4dZ2)Uc[d2-110DBA;Ag#3Be2D+6._P+c_G.dES:2KVI9]E10F8ag
\A/-8(\I;PPYS4Mf]?3UOf\P_2,DaEfP^56V-6Cf7fa?9LZ:D>JS]7SFY4Z?>^E-
IY_eZ\Ua;Y]cU5QIC4I03B00GK-I_Y>F0]4J<EGf/MUb6\-KC_L(E/W4Z(CF3YT@
,Y(/:YDV;cJ?e>@:DgQ(AR>+MW38D[bXaNAXP-M(KNO\]01:)QQG6TP:(=E=Y4UK
</GKKS6IKD.CABG7<,>=g5+O22(,ANbBWQgZ5b,,3]FE3@<Sb]3?S]JF<07;;2D>
T:3HTB@A#J8:1&;Sd/UdX&3]G@g:?]=dg)&>7,fI9[]\XC-dHOAccY\BU[>=?2LW
R33H:b6(EFXARPHIH87>ffcOH@K8Z3^P#@J(\P4WRNSBW09b^Af?L;(AcD>G]\T_
V73A]Oa4LVe0H^d:D4Nc-;@BC#0eI]]\D,L,#e92HbeU/R:HG:K>c]c3PE?^)0@7
@&+M?@>3E7FYZI:PBM?e52_Q-GZ^cM/R(Od]bF(L:X9L87X7bK;eT3@2eG&VaT+(
FT&F&I_f#)YGY/6E-B^<.;5R[59SO/\O0<RB.I,\I-A&F^1gb0NRBa5DaI3B2FT8
g)G1QISJBT]56P77bcKJ\^[7dQQBG:(Lc]ZgDDDXCZ<@?K)T&\,8652OWd+#=N<G
+OS2eK4ELKG+8RJ9-7bd_L(0#,UIO4&gZ,:&If#+\M:Rfg,f43>W\KD](\g[aLQ+
VOgJ-b,/^X-TMMBQHEFT:2RDGA_ED.;Y34;L<[]\cM,?\ZC#P6RAeG4/Bf^EEaMP
=@;-+e\d+^#?J50dM:\TV^_T;^\?aW;N>0NT?c5CU#\e.J&W3S[RPB1g6fE(.O3Q
IMEfAV2J&S\\K_D]/05/0(L^9>f\K54OTaW;,#Z4?2Y:N<9#XUdf2[X]TeZF#-/[
[I+dX@INR(YE[6WXQ)/BQK[-gVW2(dYIeDK=12;IV95WbZJJVc5VHUdg5??)5H=K
9Va?FQSNT7GB50O02\9N+Ac0e9OJL7<U@A(C+A9[,5^V70Jc,MOT+.0fDg=QVMd<
H.-ICCXLW-E@ED7@[c<,VXA:5._YK;IaTZX?PT76+HO4SVS6DEP68_0AeIG>0?[+
)[K<O/T?XWDZ@ZL@VJ:b,R@(e4NP/0VB\9>QM_Z#7?gI2S#_KE0,;HK#TdMbeW)9
TdBUF/&;38<c[U6EYfRCC5CWB?e&dUA,PP@6b7NX4dM2aQaC;31=9YdL,F&M[,>\
^K&72+(Z&8XS<M4(5/.Ncd.20/\\;T9XZ([L,PeT6^FGME:]_4Wfa(;SN-:)FD60
c.KNF;B5:X6=b6V7#J@L>Oc-Y/RLfX4\MCFN8Ha^::T#W50+G@gMJZH80PR<8;c>
LLc=B6Y?L=LG7G^(I@6aa06N=/3HYRC4(9)5M?>dZg1F,VgQV7ZLEd:c]9(G6^f:
5^]6^5/;g4\T5>M629gL_-81)QW9_Q@GR.Wec_LC-[PSaPY39B1dU/E\MC(WKR_G
TP0\:2\.MW,NE3384[5ZQ0NDS[U(OJ)_7YDF-g56>BQc#UPSLZ5BeOb^)V^[,/^7
b>[T?3:L@-R;Ccgf)1/IWD0+-S@5J.001<NU;)GEN1d@d4H3ZbdWD-A:CO0ML]2E
1/NDA2Y0?7ac9+@F_T)1+@LF_(A5MIN-6&GS+B_BZOAb7CV4+\IG1V6U2I#_:+?@
EOYe[ZUeP.A=S[67(NPP_IC#\O[L<DVSWHcU9g\J3#QH)_/4Q</EaNVg0/K3b+f;
E.2#JGP10ZVbM5EBDB0;3[-&JKc.[#ZVZMRH:D-)[ff,[bbW&JF:LX1+.:T[D[NM
:?cd7+<G_G6_C<)Hg;&J,FLaQ(>N7K]=/52E<e-bOc:H.AV[1_4J#<WMYV+cfG1(
=3?UP)FK>J5^/N0DNbZ5?XH7g705:#E<Jd00J[WSN7Y<(M(B[:bG4F+QAHLPPYI<
0Vb#D)5>&-MdA.)52BgU3/A0M_SJFaTL[<g]d??b4_Xg)0WAUSd)=@beWE3<8NOI
]d2-.O,GA0#^OOda5FfT@CW?)e0^:QW&#<?R2G)5_FH^T4VE(KGN.P=5\>[S7D5Z
M\=6E6MJc8^DE<U38=GARRbNVK&TKP?^MPTAEP3Q?d,MW+L>-aU[=7[RY4K>6CVX
eC:0]gUgN]IP790/&)fKUd9A^SC:T8X-/8+fW]O>]>8MD=cQ-dI^J1TKHA=X]48.
:A3#Re,4J+-Wafa@_T&/cEOY(29/dW;^CR>H5FLcJ@a6>eDY;OKgNFP0YYF^UTGd
=3_a.eU4VVa:1)>(,M@]Va?<@O2T73LHg:FUOM;AB^Y6dVXf\0>MWR<g-gP/&\Td
7[EH.c2<f]?,/UNIR>=Q+E^GB&].3T/IAd_1&Y1_688ZLV0Ycb5[N(6dG+2;\[NB
_.JL&K#C>H9WI)_(aG#U?1T;IVKKFaMWf2[QIEJA#D/.^C<8&56F3+A)R;(/AI10
8X1#Pa)>Q:RgF(MN,cKCUB;;53L&\b5dN4.a;:?=)ICLZHZL+&_.&X7K7D+O#;YB
Ge+K.3HC4?S=:\f8N3A3UcSfC:4;D&,R:,R<c08^W>e,ISfR3F=dH_4D:GL+fFPc
TN6g;/b]Y8KJ[_@RWdB)fPf\aW2FM<^X.>:@[7..E.bM9D1Z5+E?_G.:[U641)18
Re3-Mc3]<,MCDSK6F&?+7I?TAeKRB9bI-U^d;/F(Qb2<8A.JVET3IV);B+ObP58T
YFK1,7A.5dAS3Ad5\8M1?O6<O7Qe,dPT9WX#a#C)^7g)#^H,0a)CY.&Dde;6^.S6
9YPK5U9bSHcA90Sg>5=J<\1^IJ?c_XLB)NTBR>MOKdN0aF8R+-GI5.-W?>e>.7Te
Y@AF0K&>^gBd0PS4e@?XZD\[T@/VR)J.dQ@adM#L)?TQBME1>_MHPH9^QY4NU:@6
5MTGDQ&F.W+\H1=/H-_[ENHDMb\I0RcND2OLBWNO+DLKa^XSJaBC7&?f<9d>/Ld[
P.Ab]Gd.&Zef?\=KQ2ZeSZJcK?N1VT;#bSOf0@#\2-L6,-@,d5;</MU6g<?Icc3L
SD2GY>)YdeHfKHH0[\8f]+CKFIR?JfR_/R879R/G+<=GN2P5L4)=Q=S\5).=8FfQ
YM6_(U-a^(Pd5\))?g/BVgJFS/6VU7^Pc,M/Sg930L?/]F&JQ8W00&0T>D8^;cf<
7)\)ED4E+\P+e9E6?gKMM>^4F5BgG3a#^2L@H;R1<8V(O;;7G(_>XYN9[E\1MC[1
.;4b<CNeT]?E.:.-]<Z7DOTb@C:FA&\R?3)Ce(MQ?LJ8E;OI^:feCY=1Pg5Y[?&B
HE)dMZ3-C5NbS^E\XS15K44K&)4AW)EaTFK&NeP:c:?M)LRaR=4P2?,V,G.d8QVH
?XR/VQN-K^Jd-d-1D1fO:[ILf?RR@E^G@&/ECa^<WXE-HgYB;gRQW\@R[MCV=3NP
O=#Y3?G^(e><]BEX9)KH1:a&V]NZ+PcB,[9<[fLCP=YTf>:&#1_b6E[/UBX4QXaY
HcgcF;V,;74;L7#P>6#@H7UKQN>V[8GN&g3^<EbEf;TEW<aa[[]<57Lc919H^TPg
1N/9:&>e?.aVL&gcK>T)<NRPY+bVGccA/G8K]UJ42cSDMd>ZLHATOefY9LJEfe,Z
3b.\M1ZSCW8:>V&)eM-EY=7eF->=BV]4^N_TZBSKX1]-=NF0CZWW+AO04L<?=SeZ
]/\[I:Z^b/d<)EfYEHXN(T]IMT4[5e7OKLEPM6^f:@[:=C[/@A8,1>-L?d\\MadE
f5\gWUg48;T+BS0VA+e&AefZ\aWagIO\(0ANS0IKGKeZ=]MY#63564C5JYI]T5OM
a<?\M9FCAf:81-+M,F\g[\D(4M8;+^Ia-_[Y425[)+ZX1e7#1@G;9bE4WXA;<CeP
a;#g,BYZ9^_d&WgETVQ^4EQD9E;>^^;c+OG&MZA:7=c+1,?eP/DBFNS<gZV4@8d?
7OeT]J>+CS5Z7)a9,PdK17H\7d3JD92BIU28[(6L0_caDN#3)0_5JgS?NZed6eJZ
+(adSI75X]Y@.Q9JID,)K/V_TETD+HP(,3)aPaSOa(>8[.)W1WI?LKZ&,b=W##GG
X7ggQF.Odf^f?A:DA2Z1U/.)([(d#CD=\MWCBE7)YNS?,FVCJObGZ<F35]gC=)ME
/@Wc?9OLe=g4-]4J^gJ()X9K2abNUN\T.,W<3\O>[+V7H_^NCZeAL(4)5KCW,=&I
T2Sf2@c59b_VH0XBHe(>INb5Gf4[_A&QSOQ?K.3CS]RUQ[^E^[6^a+:(^QZ4Jb7^
Q<7?FF/5g(+98I<ROZ/P)_0g;J_O8Xd84QF&[U>ca3_3:,9>WOPVg8>&^GH46[R4
#^BMQQ6P3W\.]?.\I+-VR9NU7AUQaC[D+1W8dMT4X.)N)5gH^BM1J7dVb3G.6^Y;
L,_1:>-#7M0^GH&7f@&1J,<\?=\,XB>EWZU2?6RI66SHCaG#F?fc>dK/)g@KK(^R
^TL4/8>+e^<XGF8NM<HRg3?SMaDYJE.U,3(W?XN)4BC@bUSHU:\EH8gA3W34^O7H
gU:0.9\&FN>Q_gWb=IL)JGS4,<:4d0>R\&U)&XH=INBG9g_Y9S^+d&7W6OC<2X.J
8>a[RgY4PFJ7(Ka<143<SHI?eN9[F:;FOE=?^ID9><\AYV6@TI/MNFC7?.(>PX->
?gRR9+FPJAOCee2Ib0X,aP?-_][;M(<<B/W(GO8)J]CVb@8J>]N#P>)9:f?58T?a
E<2dS:If9ETX\@:B5d)aTPRD_\QP_^4W^>BTBdL,/fZe+bIG<]QLD[[NF^@-Ic^#
>7b+f9-@9,,-B&+0(a-]Q?:7/Q/R_/HT32Y?OSd6[&aX9aI,D2aMW9U9+NHg9dd4
1T8H+JQ:EaBbVR)>5c8<aa.2FI27VJ;4R/SG3WQPMB+KNW@?Q_4^Z:8dPOFdEG]Q
\<>F^:Ufa_[f0X?YY4]3J=D,16+M3RE.TH8^0&g3V:\NO]OTF_JR5b\2MJ&)dRU1
#eNBgVA9f-DC_CAOD+=gHR8@3EFAP60+RcKVe9.U1L)fa?:L=B/^V\\^N2XNc]4<
4Z257G6^8L1H_MB;;CV_6>4CSQe?(ZgGU(_A2[2b6f[4JJZ?E36\D+?ICQJ/..J-
BdbP(Xa6bR)2&_?REJ;E6[aI<1M_;]^S.C\<7gWI2g5/X4)FLNJ&N(:dF;W]2]\Q
]97_87:#0^R)C-b;D_g-)@A.^YHTSgN<7+4\aT];GDZ&AEa6H>UD>(CAe@?@0329
JF\\-K@?<TQbgf&gWBb<6L7^E&@&K+N#\L)c49NIZ)Bb1P7NY3_aV]13dC=KdAWR
L4?d(g.8?R]W5E>3C@\;e;b+([(-DK^U<&JAA<LZ06V37,3O<[dM\AIeY[OZEB4B
IXB;7XGZCTIM<37e6F)>JV-5QCaF-eL0Kb;VOTg@#(FKAVXaYNL&F6:]O1a20]@=
2^1bfD]5dQTVF37I#6F-3@c?C0/9C\X4c=.B+#RL4IZMR,Da3QaI38<R+7>W;))+
2^Z])QPRYV9@>^KRS<37Z+,5Sa@7?[eAR@=,U@@[d-378/AC]0<2e_6LN]1?B\db
W_@&?3&00];W;-8P88#FfK([DS9<We5^ec]eFD)^8a/2S1A&EOH_7:;:b-@>,M_g
5N@&JT\MUA=-,Ycc<BI2@f[/[/]cIN.&We&Fg6S:T+8]C^JDLT_IJLBZGFd^_]S;
WM_99B_Z>(@SZRAAL.B2M4<G-.&=J4I:@@0R8DHd?=F1@Ce/fR5dOP9&)NIe7RUH
4G[gfaHN[1XJ02&OUMHOgTD4HcQXe1Mf8P)P5>9_Ua<5TG=/7K+A8f++3S4#12Jd
\OYI6-W5W6bGL-&O&\dY(7.V6X#(G.c60Y2aWW;S2D+DPD^K6)?-FT9(/EBLIe^+
E-f:O:cIMP)eWXKS8AaLadQgR<PCEBVKAX.W)NBcR99#Fa;a9SZX(D21S]8KbUW-
I]K:E.cU#/2=^L09JcQ92dNce&0NK69PT-XX4>,S&F=U\\KfX8L:2AO?/3#@3E6Z
ILH.R3_32gQ\PZ7Z1#1eF+I^>O6@5cE<6R=VZ_fDU1BY1ZX&ac\4g)1d&Sc8YG70
.-FQ_+Y/OYSU>6&d)a3+8/0W)=5c6.1BAd+U8;COc\JN3Q50;UJe^B\CDI7ZKb94
/K6V:FFX-d7@3T(<K81ARGO,cKAPE9NJF[9;/DY_/,c0S:e]7)VbaXH,0aa6gI.+
bTPAdG;X;OGL,Z.-MU:MVZdL.E^&Y\00D@^VCSX>^=(>I2P>YX<RMP]26H9I0QBe
J,3QS;+TM6AJWbA12.;6[-SIU(KG<c_6a&Z,Z+Vaa#Tb=)CWZ/FJFL\2C2d<@[\+
NJB=^b=Q@1_0]+VAEaF^L?Y[G0R7-X3X6ebG9UNZeNH6TY98((R.WYJf]gRHKVFC
M#Y3[=a1Yg1YI]CNEc1^-&I#/C8/=f=fXJD#7KR5H(#TTcB(C-b=M2I\OG;EX2O<
9Jf.,e\@>U@DC=B2B#X::Y6fP6G?@.&S2B1Y\cS9J7deM//L-\a(-#HCD(P._g80
AY:4^]d?]X\>@Z?O;/?#>[^XT[TgZ3dUS\eT10#=+Z=2Uf>b2H7C\1_a4<E[LEZL
N9F;c7JY=.VR6EMX?Y9MEF2a:+_<KXI2>Ue18^3JH(:\K8KS/I.RN+a2.21,]BG9
BeUNdR=1J)A:<\@OF?C[d@c[<e;V<T?cLEJ6KVB;0MI4T@KF7(+dG8@W:]Gg#P#Y
[5R,fDSH;?[^?eVA<]9@5_g:f=CW+][:Zd]K&;AQG2?-O:3OZ@7YQ.<W057G+f-K
\Z=Y-Y]M535\X-@-)U6A99/Z8M5O,<@^4@1@<U.fS3-BfD,6#JAJ4HBJ390UYG=4
7\H7M\(8a,,\Cec2D>:B3K:/9CKcB#?c8@Q5#L?g@9M<0g=;SYLV?PcE4(L=,V9F
R0B))GY0@gU,eXK@=L-b(M+X>8F]99ScP,XF3b)[W/[3-]a-XbLX8<[b(?/U-WSW
A@Ga[9BdBDU;:J-J(\Mc8aT>G[T&O+1)MX#=P<91RZA26P9gVTb-2ZTU-c(7P[/,
A-[+g/SRBg@?3;TSH5YU:C,20Mc@^7>88]_ENC/^:b^I)(ES>.Lf+TFMe3_4<,0)
604:KYNT^eBC(N<JW^P/142W\/ZFD,@&;=?5)?],&.IbCTH:W&2G7g=d[a=)c9S=
.DH=2Z4S4:LA)3,V&=]PR:KQ8;D#[7.2e+LGO^c,dVb/01O#7V-DIY)<HN/01&;#
(Wd)-4YP)5BPV,8&0I=ReUY^#,_9A4VKLTH+1#@,([2D0TUdK6;D/VY7NL,T@+DY
R++Wc)Y#8@>=)FOf6>)Z(Pc1S\1:a]0:;af>1#Q=7^cE)^=Y8^+bS_F:^GBQ/#Z.
g]72LKW_N:-<83O^O)<_ARECMFWNVSL9VPcYaHUC+=E6E6^R/a(F.P+[,;1&0fZ.
#fCXbL:4UK),R=GVPZ7JM6[Q:J+I)[(S0bCI,R>?B3>D:RDA[1CD-gTMPB[+9+cL
L4,G#D+>?O8Xb&.N#1GL@N:M^)N(Q<5.Z+cg>)bY+SD?)A,,LLT7.=HN:a,JccHb
c:):PXI=9<ED)E)&LBQLU&e#?)e\Qc1FKe(7c-9WX/X7B1.,.#7J2@/&G25c?QK7
8TWGd.=I\0?@5]QWX/5HOBgTR9HaEfN[M8F1d=]6Df949POUBNgPE1CQ+V3Kd9D+
7Z56>FcK2IBdYEMXb6A;B4,]#._-PO,-873&D84ER)=E)#I_I);6C[fM4JSc46HQ
>@R91d.)g+@Q8NTM2@SFFOSYJcDGc6A]4:?CJ,I8#H<[@^HB6e2L0-g,da)bT_==
A?UAdcW:ECL:c/D4AF1.6G7W8L^\U1c#\YcGTO#dgE;Q8E?,6g]QH4O]ggWMaLbK
B7P-6OS<0/QYLGZBU^EH\E3,.aUDYSbZ>EB9]XdN4W&/A5fK^,U(d-C]f62K@^:W
-bFKCW,c2)Q1g]85=cEcFYc&@]^-TMTT?7^U03?R3(4H]caUeN7PKcVLJCMg<HKU
B@MGD[+e55P;]FWV_gZcVAZ[(e_HS=R;(7:YZ]RV/@H3b8EJQ?_H;.bORZC?Ed<,
[,;[,>+6CBW[N@J,8-IU0^G#CAVfMA/B^UePRN_35R]Gd=V5g.F_&RL8He<MI/T>
;O#:#)F7J[F+cP[X>U#<(<g56.gF+a\>/2Lc#e.]9]8QD3]5ZW:#[fc)6HL3d:7)
ZJ_):10@WLd9A;gC2d(REVQ0cdeEeccB[3/+FfXTYK+18-6_YW_MG[V\4JXDa:(B
;a]J^3V\&/_N42E-1YHW3>WO#N4)PXV2=#?DXXc;4dDTCgDCMX#_1Q&WGVPW2DcX
#]7ZXfSWB)8Z9CC6[-b.D5T0+>9f<WWKfRLf<52),19[7O_(4X]9WS\9-M)f>L,5
.RdBaa8+,QY@8:G_T4IOJBEC7OAMXP5=&]dU]-<a0TGBC>IFJ>LbR=R>2_F:/=\#
EfGS,Mbc2)4F/(fX[8ddMLeb?8U)=)27f<XcZX[._L29W(()_&PRN6QT_KVH9?d+
?73N4gU>7XdRe8/YU:XCcaTH<PFR-HZ_A(gASTO^[eI2g6-J>a\2O:ILR,TaCPZQ
@=dQ=]E4FTfg.<C1_\=W2>eNF/U\355BedSECN@P>QL^?6CIbgXf\N?VMN##14E(
B_8^[(#<@UL#TIJRYBAH^B20FE&[-KaOLGR_[ecZ2aDR=ASf^&HYWEDf1/:e^@]X
8X;V52FVD:eN.@((1/4^8>c=<N\_5)O5K<Z_-0)J#3=10.1Tc>S#.-Habb-G4W;^
fcBfBWGN[CC3F?cOAC?f71(#faXPW_c,-59SHgA^Gg[TH<3GL\6RR6[XX>TRV/#+
ZP?-3QUQ:DB3@KF7S[VKPTO,3e_cF[g#eJ57AD[E5RSKdAa_7=e^GZb2:9P[a^ZC
W:EU1@[8c[Y2gF,B&KTKFSI<U8I6105PG8ZYBg/)=ZK+:JK=e0?VZg1-eBML@4[R
PdETC,;UYAV1JbS[_a^dXb^C54MV1,.M=WR2&a3?-YWD^afQX@<60aOcB_Za[+HW
;e2/f=/=0RE#B8(@S\KD]J&NQ>f?\D(O?.4#HK:<Nb3:865/.45WfX:EN:eadA+e
^-7^MaeY)LdRB2K?=((JUYc.92[,NSAN:]+)c1\TMJ8@c2-7FN]e(X;OKR]Y5-cY
BOa_?J7)]>/\gS:>5fYJBICgaK.?D8&=G1RdB@a>bMCD&XY2(P//DDHV92>gWFCE
+J=b:6dC,+M#DW2?D,C[\P0B)ZK24dG,UMfZ;R6\5X]+H6.e@N;=FLNV2MCO1FT[
_CS(WUEQI24MV9_^OA>V1K\9)0[M1RDPbQC,2WHCULC^K=Aa\&&X)bGEfX865\J0
N=5153#ONfYX5&cf8Mf=V_O-3;Z@e]L5KRO6@f+NBFVaDW)aeHY#XCHa82EAQ0T8
2?8_6\80=bX:9Rf7@:DIKZU3D?4]&Dg]^F.BCCBJ]E1ga::92?J@_VH>;b53HM<6
&BV>c;65dL,a>T\SbM3;]P^F&>6)MO^5?cQ7XYKZ.4EO_BQ&;9F=<B]D#O)9K8cX
F0A5#WQ^BT^8M8KgcI+O/U\\GcLN>4I1fb#Jd<1899-8C#N+XS;&&S5->9fCPPWC
]C&I(P#<8//];:J\(K[\6Oa>;F_Z_6[DaeX\_@e/R<?=/[fb5>^76Q;ABG@4cOc-
f=7;BDTO]U8PFTQ(S.B<S[<2WUOL?K#d/YUIeO.?DVb4>dK<6IE.?).8e_3Rf=EI
L7/P_Q@M&F(/)?AOfPd3?(FB.IU62E@g\f,#\.PXfRYAR9I&\#=Ia^F)ffdGQ2+Y
,3^Z)H4af>F1e:Dd+>I+(?DQX.;L;VaFd>P5[&bW:We-AI;O.C]9F&g-cad)83,M
WI8:)/CaMHcLfa7F0OM\?23Q7JMN+OfZf2MfISf?=E,2#DX0+CD499E0BdbRe(H/
d4GE;AL.Y&V6,TH9^K3eA(f;NR4GRJ2J(ZY#<-[MZb;?c1f7:OE+b=+[^3N#E8WZ
e1)LVWS#IX6=+e&T&f>X&0HeDG+AP((M39g@c@HD;Q+/QLcI(ED;=TR/<P47)a[1
0W1IDR78fF&dNSBT[S-TX<B62?g/TQ4V=dgMBE#1gMH4SVSZOAC]d;.>PDE63A=)
>KE>)Ebe>EZ\@8@4Kb[Z/];7Bg:MH4T3=L=+1^EDJJ9J0HJ16LLU82b=^8\W[+]P
)4D(fKdP+<.Y;JaeP)D#(TJ8;FU824_bHW0T]b,#WU6b<A4+.@-ECZDP^?+/c75^
Qfg>?YC+7-><NVKd@aZe5WL+ASa2G[#LZ#8/L8M57S<,I6fTS3TW.&2&5,1]8<]g
,@3>DN]B+f,2POYdV36W=NW420.baUD)0ef=FA6Xd38M>dHT>^WWQ2/4e^]QX0\0
&8f_\gWB?e[P/:7S5;=bZd,H>Xf)HF>P:?cJg#ETFR1.<XRZH1[7\#>6c_F)O86:
+=LM_)9=EH0B^c&_UH5cg9N=65@#F9U#T9;IA:5SL7NWFNEKTV7,B\+I+N6Z\TW8
H.UL=OO-NJQ@FCI6RWI=A;BVaK>Mb:&OL+Y.F?R39HO2=f9L[=HS(JKEICN(G6^)
0)0:P(;BLQG.SMDK/+S070^,ad,2HHf4U7\)H0?/V3LZC]a50EWe:>8H<dBfH0O5
fT&,DRaQ2NWJH#.f(YZRFINI6J2F@TWgK]HLP6XON2?/NFU/+4Qcf[>@XfLd-bFE
M>[=,ODNUXQ_(<:U-?J54befL+;-&TZ/7?XPeI@AJ#?4\YA7V/Uc[DPGNFI(D3OD
3fOR(<Q0DfRdD1UaIJaLN8OABHG8dA@4L>>D_9)-A;_W1P7fgWD8?#L\UY-#94HR
fPR49_S^0\>?^COU3T^TA:@aEgZL8I__<F5.5+P&;8@C6<e&L78D1G6LT](:-1O(
=61RHId]0F@KA_ER8JP>_e&<],T/7^V6c>@d[eaQ7/=ABD(5=P0KG7,_MJ)FQ7?2
Q4CC4.;dZM<Y&aZ_0HB9;WQB;H4]eO1a+D\Jf#1W,<f+A[da&U:D[#&&\d(F)+P,
]PORHRd[#PB/KF0\/b/IF_eX[LEL+bII_#M,CS^Z2FN&\L+]D5#LMYRF(MG2>MDN
&\UO9JIJ8WBd?TXXTb6_B0@VSP(3,N2;g?:C()RW\c@2U&13RIZdW)OK?N6]6RVN
]8VFAT;BU)1V])IP,T@A6dIH9fJ]Q--V]Q&2A#f&VTP\H01CVdS;Oc0>eU2@Vb^.
Z5G#^(RK,a0ORV1-F6J>FHaM1Y\,HQNDa5OJUK#N8@1C<DC(=-MC86#H&E3@__SB
_G6c?eFN9HY;V;-U>4a2ND\T(ZdPBAL^JC2\-DgBPF@.O75[JDW>f;K_YV+MLKV?
81B4SV:0:9bPH;V^#O3#K>4I6E<U3#5,OD@W]HG39C844Sb<R[,)>70.36@.\W?_
45TK^ZCdb838=^g:,O@R,?YWcR[Be10P\67f/7E]A0Ya8BQ=A81B5(eHAV2c9N-W
#X,)GH#C<P<6S[/^VA52EgY6c61bLTdG#-8.X34N2e40bZOGE5WB4R&:T]e,)+]H
CLLf[dA4IQ+M#<2)&KY60\SZ&6)T7]M[3R&/c==<,</Ue?>YT0)RQ[;2NAL[1e@,
:9F.P7C(\Ab(,WDO4##4\35+E4<Lg=9Bg.D;?D[01M27I@(T78UHf9[bVMV>BWTc
KJS;)9.P_;><U^^:6A8PIQ6&OEDbde&-DR/I^U^(PG++gP)UdQK)cOW,<a@-)?8?
C:Q;)-Z65IG7Xag=\a[dW0PQ^)&EJ:;2@f=42?f0?5ad6M,d-Jg86&[/Ng,e\.aT
/cDDP,MD=;8_ZL)b(QO#CdFMC9_:Z69^_76(SG3cVGO_SZDH[J=BO]__\=-S)_C[
?<7&S+&e>NJ[#[F7b_(TTQSd@S:d7GC5ZNI1DT:bR;;dB[\^(F5+3;Gf7FO91;=D
J(L,5@DE8D@@51URI/,/L.>Z2_g_0V6B[YCHDJT=E:8\<T3DaA/AQ_W898[M\=Ra
A#6#OL,a4BWc?P->>6DL1SG:a[VfHXGPcBgA4WS^TCV?#BeQ2.H;4]>fY[MTP<.^
cM9N#U6]ega=P\8:45?[_-bRK87I2,93KSP(05(Hf+AH:V#Jd#S1>Q8:4[,H37Ac
FI_SM,QOVf-=_6IUUQ0T4[[ZB#\./?eREfVS0N7LQb),>GJ\BM>:?O=91QYWSME7
=c9R36>/M<<IYL^.,=V3^7Ne)@V0R[\YKF1;1F.:;,Ga;?Y(cW/^>5S5;=I,-JM<
U)>[(^eH4\X=<#AYeLO3AT0K0.4IHXbF7b^CN4?)QKaH/fNFBS/GOc,X[2>_@Z#G
3M2g;^[_])&Q:#0Z-Y6B9V,;AI6:_DeBCb^a<d3,I/I?H[(Z9_SPA2K:CeJW=5-P
OO=E5V7MGA[8VM,b((Q94::K[\H5<G;7bX=af3K(A-7R3<J<0b:9@7Bg]U,Y:-4U
dM4&)AM31I>)AR.\A+B3ID:C+>5FN@:fI\OA3F@VW32<V^YS><;.R2SSbMB1\<PA
(91/,:HF/^\#BIN57cEBN?ZH,IE_e(SZF(J.N?fX[IPd;eU]B-L,/9W9Ea5WF)QA
#e\U_(&;c1OZbI/J#^Y+1;9NG@A(Z[ZTPbM5L(QESI7N?d1,LS8.e0&5]X/M>25.
RR,3c(bT)_]?ANF4X#\N;2E88S6O\:#8ZHMB4.caESQeQP5Lg[BCC01#T<NRC33.
HBLGR0ag.-C<b]I2eG-7C2GVGdZf-]8I0PLV-7Z<>K&#56B0_@PYe9gKgf2X88K?
[dSVS-IFQL-JBRUEMA3,L:MZ;,e)05;B8BSfV\b0?,K@e3;]]L?+ab_QfdR2@1E3
2-)XX?BGJV1FG?LQV6SX9MPX)SI1-33-#6:fTLL26)6384E//=Y8(W<71UKM3&@;
N5F32(gKHGS?)87B&#_:CIR4d:6PK51Q]a?Zg1A4.b4J<@VFUIc4Ua@MaY_bbfDa
XZJa6d1R/97LIO4[?7/&2_eY_H(F&HUC+gfN\ac16Jb>Za9)2700cXeJ8]STNGc[
PN+J7;ZeDLM[<9)6cUU)E/?MNa+QJ2UA_KV=C?g0EAG6@JJZ.2\VI2-5TfSG#(\-
g:ccC&W?>;d5PPS>(f:P/5g1ZeS.5(eM_:KX4DSKL;;82Q_1AVeRgO^F1P<[7+db
N:-6;R?6eS(>1Ma4>+D,3_[WI/,#_TRdY/DB)Ke#V.cZEQ[1IA90Y3D\MZ8]790g
U7>-d4g@D\,FCGL9]4NU^4\WE4U#Ha#IKbRAQ1XLXKV2;MGE,3,YC-3Xd[=?.NbE
0W>C2US82FP[1_aULeELC)/g(U<225#ZfIL#9B;Mc>:>IA/C4MDC/b0:N_YRVf</
SSZe&:86ES0,LCQGCQdYb1RI(f\4PTcD2V>+LcFCCJ3D0H9N@M3P[+XD1@X,,9N;
W?.f0VH=,?2^W@V^96eATGF:dE4&B2VUQagCDBMJ82-[#D_dcD=edEL(]V;ASSQ^
]OAb&aSJVGZ_O0TH_eP3TKFV-I7fC;PcA=aR&a677<c=U1+99??UeYBdQ9U6.[JS
Y5WS@1g/IcQ7,a)Fd]d,cXRc[;B5>&9KffOZE8[<DCP<C6:^<X@3cY@b&CW&3,dN
cA8f::1)BB:A9Qa=YH0]B@SX_2VCVbJFLHW:<MP=fTX8c[XS/bRPd[,Wa=T73C5c
Yd-H\=4LUUEHeGZ?DHT]),)>F3,N5cRAfD6>V[4P_S>,cJHddgLVP9=?H8YJFUV=
04K5]cT)cY;_&6FMDPNIO_E50YJ-Id7bM]FV@]7AbV3-cYeT9I&H2P7[4F,,C1.O
1QV^]E3;WCQ75C:XfVT,)#<#+6T[J\,&TW_]7UC()6E<+4T0#[3WW=SM=IYVNANE
NCP4,)8b/e8b8-#R^6GONCXY7NOM)^16L9=3>GeA14^aR7IP5aEL/-;d_eWBb_C<
I)5PM:g2#c&GcO4653e_L+A08#Ga4[LM&d_g?CUEU.T,NX@R/e5=a\Nc5=Q^:R+G
?(7RQW]L7\X-[YH8&1Xf2If7bOUTQJg;>)ZD(\YdC;CI/YIK(H-D__I^ZGJQ_#>6
BTG&HYX9C\6.#O\[[92EeO\534<UKF+R]dDIgWS<8/6[Sa^6XZ/6><1-?N.059dU
_,&H.cT0>9C\L,)GR>_HPX;WgLQ>CW9^S=<#:7T#?T64_Zga2+-_4[3B[Y7aU^<V
;aGa=<:#?K[BZgffX?FVB<f]@aUW:e7+NZcGb<++?A_K-S^dA8JARXYR-HbZ-fS+
Q=8G3,4g=Q</9,0/@JJ\DQ9L6<UMW4,>GPO^gTT;T?W7XZES?4bJZNS\CC<(+<b,
(^NSge@+AZ&R.Lg@.LdF&=[Qb_-C2J+?BOgA(g15#RK_#85Jb]SUQ79f-Mf-R4C.
Q<,715BPRG4RFb5ZCGHW>/W1DRNQP0)EeOI5([Y1;-((<GU/S4FNE?;^H+_^6IWf
0-NW4=928>,P-5D]9RHOcVV8#=).EYLHMH19X.:[#e,OMT<NTI[4LIaKE5P2KEcQ
ZYBdK#-d=F0F4>IdF+7V_A06d,G_J4f86W<[+7Qd3:&d2E>d/B^NJ-(QO>FV00RA
;N9A:<X68faa2,^&,/Oe\5_dT1P0ISc0Tc]cX^N\AP87]Z,]d:.3bZM;E,73HX7=
]WYH6+Y>9)Z[.Gd3A^D(?L+^6bEAVLAOG?],JZ6;:PQ6c<T7G;g-K&gLK=42fTPP
Te_=/(UTY?U3W6<cK_-9\Pe,#;c2NObd0O?@Sf<Q:NedAV#]0JL)E<E4=4FDKTPX
J4^Z8Q^,CJB1?3^_NR3GeT2L3_6g,IBB5cZ4F3&Xf=F&gKH5aBR8-Y\N.(c;:M._
Ege8:N3:J+EAT/0DP8-f#.CHf_;(];&V=Z:MO@D/@=<0,?dJI08]a(SA6NQFQ^/2
&ALQcHWd(7cAbUM:5K)<RDWN.YAb>SVf4C-BN3fS.E9,C[OG0NFgHe<<]bY6^0DB
JLNaOb:?ZX3/J8DI(0[/4//(4S532:FZO1J&M0H_99H3+,=RU]WbRXP;=N3ZO#3[
eJdf?0TeC=&^TWX72K2W]3/#8aPYL=6P>U#7C7FIS)/Uf567/)P0RK2@O#1a<3]K
XN,DW=RF(6TX[]5A<G&(0;O:68/]f]?/8B,J>Rgf\61F.gAR&<Cc=A4RW#577/2X
17M5FPA@(E9Z^[a1WUUI\9,fLIJ.Y///>==bT5,CRO/+UW#M@D:e)Q7bZ#Re>\Jg
_CbG_J/=LS<7)<03V(cGU)Q;:M.Y\IYUPQ<\fa68<F=N=?XPEY>W:EJN;:WW>[38
GT.?g<=\X.<(Q[RY^Wf8_KeHcHU/-V\dLc^)>\bLR):#T.(S(:N)b[(_3X@7J/L2
8ET^+:Ic,HWI1DAd06P>UEPPeL0IYY395=_\SA1Id&_KAM5.fe_M@NF^RRSL16T^
da4V&V0e0;cS6F9=8&)S3BB]+Q9U2Ga+6W=>R>?L1T+FaG6[66AB=AZfNdG#+H,1
Pb2TA4eJ^(BIcIC@_8&[cM]+V]KQ?:12d,Md4F<@@TO=-#bT&S:gN7bacS&(UafN
2>ZXc2^f(71)-#)<bFUe=CCBGFL9<2c(UMVAJT3G+<===HB]C2Ob@aA/.@Qf&EG;
NFF3dF>DHZJFb7Ja7&+S\)Yc0ZBaaO3b+\e@TG3H3UG\G<_7C#+)L?@I-3@#9:CP
;Qd1P6VcK4L@>L@IcdgFC&M2TQI4C.gGVgB._W(7><1dT_c2c#E98TP9RN4V79@M
5E/29gTH;,PX]9F;2P347J\<5>C,V^a-_CBN]3@G0,.8?=)9d11;gGEZTYKT(1-Y
4@+bGB0N\)3c:NRb:PaO;Q9K^EM<EZNV;dVaQ)^=?egV/Jg#2))8TW/:PJ^#_deC
HA2K_:b([,5NT.e/8Wf#eE#[P:/bUFZ\XA&LQG9LeZD?JM&<NB0DTb5;-G]VbZV:
@]PGAPXQ(YRMC#=5W)GVa[&R/_KT=6Q/)77H_>3+\QOA0Y,\^&T:KS5U&gU3^7U,
94,F1ZEZVNDGQDNf&0)^=>e5fKMce6.&cG7@<H(59g<^1dEH=/)R><6@TYM6A2bQ
T<2__?F1V>0_L,#]UE,fg.^4cTSFPG;\6TH1DPD<M:TW1g.,VE?FWb:C/aSa0X#:
B#g6BK<(TGggEJBY\PB5M2LN#dQfX_E?)UOa2C+J.>;a3.O+L7/>NZ=VZdM,faOR
XA[PC>PUUO9G@.eg9Mc919f>fRQ;+R47<TX1F=(W+^:^e3Mb;eLL8JSBaf4.6@N+
LD^+LZE[\TeP.-MA[fU&BN0KQ#Qe;HI[gA1_]-DSF@6K;)\7Og/,E(U,)/N=D-YO
FF;e]]#(T>M&81FP+()VAHX8-W<AX0&AGA<3@3_4.^+I+_W1&4UNc0V.XNg6177U
^XKP17H9&KI:Ff/c)?1;?f@ZP16.Eb_6P7Dd8\g)KIcL9\IPG#;Rb8>0-U2))SRG
QYXG;RJ3L[,.8<2\\HZ=._c^+S(>+O=Q\.>E]+V-<963SDe6)_31+<6CNXD<Sb:[
EQdEaTb@\XY7;SXV027[T6+_7.D,fgX5Y=-0Ze?6gKE=^9T.b/:Q/VW;]AU2>_#\
cN=ZeNbB5U=2.E6T.,TOG0I6fZHTG.6T-3cGbfIN.)J^+UQT_PCC@5dA?aJ8W)12
K0DR?LI<DQNE,WAgT?4fH)D)6WLMU]]OJVV0DMAZ9F3aMbaUE]>3VQ>T]^Ibd3Vg
3KQRQ?3B?VQSFVT[@cb_\a>[A4&+;+^DAVRbMVP(DJd&,,0G@g->GYS&R6Kbf(Uc
WPXVPA6@=gA@>-@HW.#cGO@5.aHKK@B1PKgRe-3=@aN;@TZ;MH&]f^ZW,+=GJ)fM
C1&5ZUIa1FQbG.BANO(4[>]YHAD@?#f?Q(ND2.9A2P(.),6W&M=g2@(#VEU1gI\A
-1=]/JKA3^BKK0H/+,bN,-^=dMb7#S/,g5RZ-e+8c+LV/eE.I&S/,<6@4DGNMWGE
NN<#1N;9-C@28a)c9;,(-F5W2f0ZJZCS#.U?K8C6U^aDef>NUV;_b:?0.]?2BRc5
Y>8aLg]B:9QGb:;4Q&_7R:,=ZJ/M#,WS>[Xfa+(g62^+)@-/@(cTc<+OdZ_,?ff.
;YTBU3D><E#[E.ZGfcIJc&8X9)B[2HbNOH0@;7K37.H72P05#()IB:H)B\HQ(6];
H96MUT?>E.&6ML-IEDL&TI/d?(8H,=.>cAP&1##/5M?N:O(aMK,.K?Xfg)?NTK7Z
U_K=agE6PE:T)87V970fdT9<]V8,GeBKag(e2c]O0Jb-:-(TA?^8G1P6dR;PO]7G
N]NUNX-FI[[9)JJ2OFg[7CgZGfIA<@cFRO].FT0:P0.geWKZ:BMe9J?JM37FJ(/c
IEfa4gJ#\X09\-X<O>HCgM?\15+-Jc.TJRU?(Y=ADKNZW>He.I)5a+^YE)(W)OI(
0g\7-N[VB9YeJCDN1a,Ec^UU6&;@<MaHGXLC?fC>3V5R#c/B>,7\a5P.+cS,(Ce:
g?ZY\);f./\/18QZ)0d1??THLTAQ6(g175XcYeT)M394S_CE83HQFIMQMVcb30Y]
G^4)L-7,JP/QKZf&e-8OWS,eMcL9JA8G<Z6O8E^/a-?eJKB31b)1>D:PB>R:<]N.
+g>W-2XZQ.Zd6YM_,:/bC/c_a2g1-FL,)=3^U=X4c<4-(8g/)7.-([4_S[(KABXf
1,L1W+KN<1.]U_V8f[Hb9-D0O5UTKWf6TebeMN620C#A4f7P9\L4^Q><4:g66-I;
9X\gA^,U3G>1Mc+J_RI:A<)3J>UO4L:I6[5VaJ,AcU,NO(0U1P.0@bYGGd-K,>2T
d8F?ZdY^TR5#cO<g[,M>3g.?f&&Dg(X1VbNRJ.5H>d_6L;)<-[QA6:XNDN(\^V#Y
d6ESP:^Yc_0ZO=g#+SDa:K9&,-=(#6USLCg7_gJC(X=NZDDI#K1->>8cS&/Bf4/F
Q@KLa49XH5H^?3791;<CABE_-f8^9.]3I)5Nc/BO^Xe.Dd.<NC3]SLOKO#?3W-)0
>4J/YNMX>HA3fQQ1gb8Xe><L+T^E?HQ+P\dSaXR&bd1Y@G?g>2I7>7IA[,7]:?NI
J;-UVfe1eT@=P.C+dKg1#e^FedY6XVSQ-?4D(BJc5MbagVGH[T4bN2cMEb&R)HUY
OVB9>6N3f3N&^\^HSKT2M7CZ9D](b:d,ZN)_e)()E5/8f_=:J=?dN5>9^dB_-,JT
QSY>+7NAFX>LLDA;W.S,^G[2;gX,982de4;M1Q3TgD::d7+W_7g1fL9G>U5Z?bPd
@R66Kg0R<I#+_?2U,BZ_a@b6Cac7Z508)WV99g6R&K+/Hf<^@:f0DE+./M-)=SZ>
P080eOHZ0TCa/RZd:2RM7)#YR3cHFJ]WgH#;_be=J(^+fTEECeg97[Y_+?4/b_Cg
.@LKIf9__0?WT&KS:8#WS^g[K&dV@R@0JTZ461)fC&(]A#(3OZbIA4G0TH][B@@X
CX#ERB1Sb@QX6SKG7528H5UZ.g2H4..BgKV26NUITCeS4+6<HfU#P(cNL_bF:_0B
)I[+Y1CV[Q8PS4\^OY&KXE^V?Z/V5AfT6Y-LgQ6Vb_16b#=+&>d]GTRE6^=;_L#Y
1YaW#G::U;F>(C4c):@/g?OUZ&\OTcY]+J4J_)bT<O^GH1=3C_K4-c-D?>FKIB^O
UP)UB@UObY<P<;@J]@HVVQS=NL^HR(/B9O^#LbW?ecX7(KdHT#4b,fGb=gAV&&GF
HebR?E(3\O-1(#H/=>T5RM7W/QI]K[/H5&baM6W;J:ZV[PY?L]GR8B)JV1BW\1g1
S:4_4RQ?JI8;]8bKJW[AFSTL6+VfV>;YNI\GEG,B-I.AI-S/H[.74?8bQ?#c^JY?
QU##GZ^I=@e<b?1ND+Y,a2EJZWbb\gefMDFV/Y\_I8cW:[)F=\=PH(cW]A()::YV
@AOZbUH8E^[=73C3];5\-28_/9:#N:a/NPYIbG/(=5,4PPNabS,ZQQgJ(UcQS(Z,
BR/>aZJOaaO(:].,Q167=-IfH8RF.ILQ@&fe/\V.f+Ae>]SMf3O>GMZAM2T2eAa)
BNN74IU]8fG9XWOH1Zg]@g\L\+1E.bc2IA9gPDIXZL69bRXEdQF.S;,)SG21T\1A
8.6XEN2E><9N:/.<0,c4IbN,T;QS@?d?015.>=0>M?Ibe[HM\FSCB_D8RPA:dfTZ
UMgYM-1@YPMC/A(^>>b\KA&W4PZXOYXF+\gN#E+UW/@]6T?R++;71>2([F#U]8_Q
JRPEJVTN9++>E9N\#L0,5(I:9)F/geg,5aTE6R&+6d9TQ0NfWC7[7]:CN+_+b_M/
I]1\O[PV(UWGBB=+Z=,4-?X[O?[NBE>I7DbJ[_0V/J3cfUe?(?Z+?K]+(>4g1JQ=
Jg#AfU=D4Sf9+UJ0EPRCgGB)&)JBMECd(H>S[d_U)&=c8:(/N]bC+9OG5G;I4;c)
cL7<@ZcD#TSc5.b0<a6a&P_=,JX\?7H00&:Y(VD(H\SXCWF+@]UTA0GY=DCH2I.J
22D.c&Ndg4/&I9&A4Z+[0e,f>:11<R5.a1)&-N7>2W=?03;W<H)[F?GOVR@)=DO;
P2I7?.\f2AdER(;XH0;)]RS5;Pf,L2AM,C(QT1RQ<ORe-,U8JZ=b]fHBPWeE/MRO
_]:eT[KYQXF3a:ae,+P_@,^2\E4ZU_gW&Baa1?)]5;BA5>Y8C9Bb\?BM2MddE_1-
ZA8M.Z(<GgU>gEBSBU-\6PR,bQ^f&S>&^b(NP8(Xbe3EVUYC=03;F2QZE>O8/RNa
LHI:Y6GgRC5AD1FXL5]U1GH(>[R;Cb;O:dK2,ReC/;R?[RJ+]&<8cN#<b:2]Z/L2
d_LELZa1E>6ZPE8,aa8Q5J8ePZS8,:X1KK\caZe;g;bJD/c&@B2YG&/8e_-+0@.4
=.)UAJ1/I[X67c[#0NFCM/=0)a1g<a+S5a@3,<Y&0EgSCLMQ/C+g,C\R7\O3FSO:
B2GE#b<NeLC)YMX:/:]M6JSKZKLOY8X,,4>MVAOKfWIc-ABdLGOMQ5gg^c=+.>5]
Ve>\?YN5.c+K<DSXHfH?S1&I1??M^<)?03Iba+<.DBDK+[[WT@XGB,<VJ=:])Z9a
K4ZB.AO1QBW=Q&AYH0A2@S(EJ,4EU,^I?Y..MN\f5EGP9<#I7NH(7H-YIN/?,JM]
\:XeN8B(gA)OJ3[(LgO7ZT6ca+;M]A3a+[>4FQUR2_D\JN(I/U+216ZBeVO4@KN[
/C#Y\&S1RU.PfYSJ#0V1Z.@Q[L\VR_XEdaG?7-3&&1dD5AgA1M^Kc[4=eIYL]b.N
EED+I14F\JJ7Hb)d0;ME33aQeT))0(A^J2_G7=SA?IFY/+Y>D:5-J&GVTdAe;N#d
bOM,>B0>a0@9b+,MJDY:P)U,L[V@QGQ\I;UGS<HT,S@.N=\#9I=F.16S+=.7_)_X
:]Qb?+OCYMHK9f4eHa:O5LgWA&?X;LHC4=IGYFXcc<7Ie.g6@IP^U@/?/5DO8#Mb
,RfFSW-KZg.@2.f@U;O(.)4&=W,V&>2UZ2;QP+e[TYM#\\F79@KP\#7O+91^PbGc
dfJX_DSQ:W17@(86UP:=7A6L&cX2FM/T[d(Mb(T4_F\VLZ6L+]G-XZNObGeXgI@D
8Tg18@e,\#M_QC8CH]\ABG0HU]4:JJ:H;GA]J,HC7&?01]OSDd>9HANOL$
`endprotected
          
`protected
Gf:7+f-5OIN8fEZIN?97R0R&^L(I_N5<ARG\C2FC@bIA,7V<#+O..)#M[I7^8X>I
HB+0O/9gY.HL:O:\DV_G/d&G#ge2#Q73MUb3)Gc=,K6Sd..VE[gYP8<T:\Y01BA^
#PRAYDJ<9>ZL0$
`endprotected

//vcs_lic_vip_protect
  `protected
PLJ5,]b_CSG3CB:Q&^5afW9X57)4a&&+?PK8gF;M\f?P@?\dY1MN0(>A6g4M9_c^
9+>8^@2S5P&UWX5A70DS9WCD/egBPL5[<=4Z;644A-PA6[;S9.WRELPR6.@]Hg-)
FXY)KP@^MDZ);-.@+;;=EB(HG5WfCDaQcKCePHCIJQJY.B2]I9].eU(>V7F&#(N<
dO)MYc:,fb68([L9^U36d\C\(-CDV<^HS^N79H:()\XPd(PDbS/BdVg0Q.P=a1+(
6O;OWaC=LPU5f<C<Y8VfCXf]V&W(egY<7&PcIa]7>;)YfLeW/2_-4INOXSQX,S.R
-NgD9e[He-AU^NHeA&5^UX8KG&2>:T_)7P<(7=e4a9T:]UdBU2&ZgLBOU><V(PA:
dI-_CeYD)&2c/OZ\WU_1V:Ace7bFJ]@#7.35MC4NDY,cNMKVaf^70?K@f2K@,S=,
>Q>^NYAW>D2)=3YA8QDg(WJ.U8-X9@HgKWYa?<Ig,aKS]/N,7Mc]E8C/1-UbGWWU
.#@=&23K9_[/1\A8+#YF6JQ6e]8ARHW2CF;MJP/fcS\U=II60ZGf=ZA=;@5b.WN]
A]fW=SB9,d0=DI4J#1,(PL5CTe[a+_QUMJ>2;F2d_O6FU.<0.@S#[gF)d\3RRR](
=@=-G)]33I5[(HaO/e6PBC+7+;S4RH52_NeXb:D=8M9ag_8b2,Vc.\N.S?Z8IKKA
K;I)bcK:_&B>dB^bW(2;O1J@<8#(?##Y6<VG/@-8b&>E#+#,;Ga>97YZYZ&,2?.(
-NI@U<:M>BE&PbH01&-7D2gXZ:=VgZS.\#;e<f>,?2T>A:c/K16b?-VMLAD-efdI
H4&V)Y#WdLUBI^f=]-9aMNf=1MEXS2Z]ga&I&5X+_]JU+P0aUF3+(OA472e/N6M3
D8=@Ff;;G1-X&D6J?+7(19V;EPO(,Y/b,YdJHXKTd&T4?Xf4G,><,b+MPT&G]ERd
@S:DN_+?I&9;OK)=HM8c)DJP.#KFD=[&L(0R-2EG./2FH\&_>#3.7)2?cP<]^VI5
WYXe.LV)>X;d^+YMM<;C&XCX6>#fe4^,G>(^,HBDC/8E+D>1Odc6/aR[>Q4QXMJ@
Y3=BP1:d[8Q8LN8OS,6+c3_62-e:&>J@3EIKHg1g=LW;HW\2964\d0_P0^I<W)F#
d)MHBe=Od5g.S\8G41+JbGRC89Afb[3T1IM--1[@9L6)]K.bNZ4+IfZ-4S,#5LJ?
GD/-;H2XcFVASQBYMc@eaI6MVge579SgJ:H]/VH3L@5cY/ffOT,]]]Od,]@Y_]\>
?AK8?R[&,99HBHdXJMFCT07c844If;@3^2e6d+=I7-N3)cO777N_APP6J/H<IFSR
>@:OJWN4V31Yb_Pf1U(T5?FJ:K?LEI^,HC=(QTW;(IO.[\1503M#RQC/b(TWYGXY
(HfICAg,+&Ng5AcV0)4)C)_@1-]L;@;=Wg3(C)MLPN#U=)g)0<5T,QCVE1QQZ1^5
\c@8b6?W6HKW,-9D40K6LP8bQQY(--4)B3c_)>H[WZU2Z<PXLD393/N77bTE^;_A
>?QY/Q07\DbBeXVEUCTb0N2LK8TIb9),H/4gbXcc9d8MXLV[(-GVR7C[a-DgW;)f
QM0?7[:RB_EHX8]U&M9GPL?;J4HKOV4N8cMW#<W^:?-9GSKW_AB7L-MB+-V=f;C.
/8)LW(6J5S>#Y#8@O_IB;PL7GQ<6fR=>/,:S4aRK<8<=9;<\A<E0L=.F+201B?RZ
#X2I@_BPDG1J(/HN4GX6&>Wc>eeNNN1g.KHUZ92RT.OF061RMA1S\8gV7(FQ2TT)
JXaWQId/5Lac[;^VJ4ZX8]>A+D[1I_K0Y1#@DB;6<a?2E5Q092d:H#:,-Rf>^SBL
]I1DG/1SDd<IE#:<>OAT8#HYS9J:2&.c@b2AZTM7>SI9H+1SXO&JY=[DE(-1IT8;
X+TG;HXYSFXc-&TLHRJ[,R-1ZCD=5S-H(GSE29bIT(D_>9IG\Wc3LVDg45[BL,O_
?A1e5a][eNAH-A?4X[-\</2PM7[K>Y)FLbW]N\aL_9<X+L#.NHKcPR7H7R<f[J(O
4?G#?J[55\P6A)-Gc.P2g\(<BC<#+edaD,eOed,B4K#X3M#=<6.XRP(aZK_GYV3M
6@;G]WZ<5X3]DM7cEc8FcI7MO)]YM9I1WXV5_)7Y7E1?3f>9GHB+=&_;c7/e.e&@
7,KAF_g^M[=JS:\F#,7<33/U:a<(@73;]9=6ZR(3GK/O_>0.+/01(;S0^N<\82#<
ZDN;+_WUWFcP5)>_WB4;]FF^2Q+2=;ZY8=B:A5.V\c>H#)X8d-;g)e96K3M@TZMR
[./^D.&+9g?E7UXKcg;BDYZ^aNe\M?;,[9B[IP)82<WY9V\-KKeW#42CWWAO6X@>
LYP7PbG&&O7Xf\ZGdK5eAH))RObc:@]9O:B/1(+S^BeENV^_O;4L>.CC[F;0\M25
bB/Z2g\GN[0.[G;<GdR;DDb2YC-96,)X[<_,GG@-@(UOC[]^g0^^^1;39=N/3)g-
I+UgdZ,J>9TKfL1-,I^V;5R#g+5@9>A>3&M(?LSf;8[#,.F>dE=_;;eO8:6E(:=G
\&B(Sdf@MaD=\g)#UG[Q3b(OI\b5CA_R0RKW4U/OU1/_b,2<N)^:Q5dN1Z21O]^J
,C7)YR@W]AcR_:9E_Q+<a7L&PO_;A5d:NKcASgeb2]VK5C=6B@g(Sd@05F>C=UKH
c@:4>L)U5/)7Q8,\_QfHgF@GgUQXTf2D+^;Q#f=TQaQA<FX9:eZYWNB?0?SQRIdH
BVCXBU/;IJN?Z<.EC+87C7U\T&SH5(ZGS<):E]S?)8faPX?P7aP\Y,40X3IT;1gP
M>VQQ9UY4Ua6<YI4Z]^@P2W]]&:XAR:,Ff?@XR-Xa67SWaGJ3^LBC:Z87<7gfbgK
\TaF7>OLF_T^V[\7/K_dR^@=dc9MOFV,E&\XZXG#SO=ceWD4#>J\2JO^];J-Z)Y5
1V<eXI5+^Q8CQaDSZEa].IET;1U#953WUZ\<<_:7Y;6KcE&B<OZ9:b6W6].N[,L=
?[2VN?\ZW6Q<S0.e15:._]4f5La:JJ30>;;P,3HTS79]Y222B22Ng0,HK?JJ\I(V
HNDQ-g#P5SEF78fZ3FXGQ2<&Z@g.=HG/ab?VXeZ^IYK.Q=2Y)J<V:UQ1=\#GNW@T
(@VGRFBDd(4G,=88@&XS)?+5cIJb@<;N)+d#2CL^H::dP(FA0_#XI[=9SQ+=>B6Q
[c5VD-TPP6GfVRZDD\Me;<_4:e1;4XcM2?1O-KR]FOI144??:YF7QX264F.7/H(L
g7WT=K7a8^cM_]\Sg,/g4MY-e.@O:XB)4FK_8<5FR<dM6cDG&(G/B@@e>6[958?:
,&D)^\d>0L-T&<CLMDA02P0KRc,@#S.:3;Mc#CSDL7USOGYYW@VOH]E5HbS1-RZQ
#]b+=Q2-[Xe/AMZe)Le>-Eb9bPJ:[0]]>(E2C8>=K8+.7W:?C4(G?-e.X[IH#LO\
AG>/O&(c;8c2I-Nf:UHgW4B/gW#Hd8KEdIP/c2gV3CQE3]FL5d3D:abNUe2/R7+@
6<Q&F^>H-VXGNZ_a:d[EGaNZTCFGMX\&1ddDRV6UP(#;44YO#H9a4DF&]Waab7\P
X4A<Sb(?:N[2:-TV&^P0fA(._8PKD+&(XeU\TN^dG5[WE\edKd/(13SG7#Z/[Bde
b8fO,P=MF0JUOg^LdS^N,eG:-M1IDbE:6(1RB/0F_f4gaV1D<<K]N50XE7ML]dS4
M292c@0=TO0WH#Tc5AWU:LI24AR+.R#-\B.L;-@dbM(RV(O27OM(YF73B8a=??<^
K17A]Q7ZK\F3U#?GO_;9adRUSN,IR3E18R9eA3A-PCF]aVEZG9W,^;\(g>8/5]#@
AL:QF<Eb9OGfQ/.E4gQ0/L01W[6e/\Z#PCWb;\3e)SX+:S2X?E&&51#A>7c2LMQ>
(9cI0g@H#-Y?5\#S16&TL_B+>Se/@Ig]0fBBZ_8[RVQ+11E1X:9.GRNH3gHfN]La
@,g6E)^B)dPFT<CQ^=@I6JO>R4VaN^L5#.]NP7=BIIaVU;G0YZV3c-g/0YEKGO9J
I70ZW4\CV@X7cP^A27[:C\1[RKL+ed>\Yg-=SeaQOMP<UWOR?PH90C:_&[ZgDJ1[
U,@C2MS0O)9)P;-9[<^d14<8)Mc.CKQU#I&#?^1.I;9DDI_D7O,]dZEcJU@RT.Y^
MCeA9.UN_K#)QZ)K]gcU>W8\,OJMB+Z_g9W,]9SVFJ);/g4XV(?GL@MXgZ6aaJ=3
KS7A__)dK/D^6Gd>Nc6UBe0/Y?.;cW\.bMR_^3G,cY2_fCP849W\]ea(G:>6cP#E
S=G;T#c.4>BIUTEU@MY4Md-;Q=aY74OK.VMUXT/@Se2W]IWB&I+RQ^7N@OcS=@/@
=-,2I3&)fN@1]DB4_;:<=9TIS?G@E&4F^74=7_9#Fc(QWW1VF-Z&)\HWV<8B#R-2
ge,9(S+IL;R;@QOOMS9.@.1U-.6-7761693IabS_e.gZPb&G.ZG)UZ>Q5FUSG)TV
F:;2ZFFb/BIUR@cNa</KUI^b.L@T6#Rgd7@I=3:\Q+N]GZ+S,DU4ZC<5WOXD)OgG
<P4L1I(D2,PA5<KKXT?Q;]fc],:/<IPI;+2#2W2g;-D6E#5T,XdZg9V+:-?/^B=W
WMaS</T)&FMV&MZ[bT6-agCE&UW.dB]CMK-+=W80-?IMBcZV^:7R][O>ePdH.DXG
D,;RODc<V,RV\VgPb^A=bL]e2XCEKEdPK_573AD,Vg\(0^G7NQ;?CWgg23T\P=PU
c3AccRcLVBEX;3UMAV:-3J0-SL(&I#gH[L>a)MA+61Q,(E&-RD5CER2_Sc4+7(AO
L?b:?e17a4PF?C\a<ge0U?JDe\cFR0;,NSJ.B5GTTe6KA9fc@2_g\#]Vf,YBBU9#
+-:R4729KL4F50M&U:^e2V8G.CUE82<8b_;J:6C3;ONGfD-g[Y0;c0E#AP_09JO\
7BMb/Rg;>JTXX_L^aQ/\\B]_dF^[S:?MFgW-HS#IKE4XJWZccCJ&#,O3I.YGe_;Y
&16b3[FYXagUO^Kd)8F-X]MN91XQ@_5^b-TU5KY,fI5^W[;<f&AXULD_[Gc;g.FM
VaYIFg?<(Y.N[BG3=XV\:--H0VN,+gT\@>(-c>b0bf2<[.C5IO#=NE)W4Jg=\=:H
Q_Y:QP:]P=RJM6/c7,4_KIA+](J^NdG?-=>8;I/U6/TFC[XGX1HYB;.05)\H@IQb
X<KOO]:>4/@[T5#1^<2&OKbA1_0K^()+/cc(Kg)]S0LG@3I:DVeZ<KH&Q#&KX,Z3
Y/,7:)K\^<;KUHK4@=8\9+g[<K^[.S#_XWHT9H&X<.c-L8#N#XZ1Be+_BUP(TVN.
R&EUDfdS\#BTc2G#7Z(XQL0WI^SHe+.P3@#e2N0M#DF5.)-6YRL_26\+FEGT]_7D
b::^S0N)@1XU4T.;]B\/P+Q0MJc7EY/DP#<Qe3]UaU82N(ZHTT,G=2V/[1F-#U9^
[5>UA_M=Zc.U7(\VY=dUaF5ZBANL.^UYB#F(POBYa)@6d^H?F-SaE8L^-.XV>4b1
a8D-(.#4=9^U)+BI2b,C;/Z.XB@PR@9K[8NWRJ2USYBa1G9\V@:AM=5[S^]2VZ7@
<J8_9bBCY2VST;PO#bY<FC#Y^0F<2FQ;T-3.=UUfRLf8KYEGK9&9THQ1ZSVY_?;V
1PATQXR<9Q.B+312@:Y2@aBVS<75_7SN,_^Sf3OMEY477JG)NF(=>bcd6X8J-d)6
XOP7EEfG1?SV1+g<e/+9fWCIU:/0M1-AQd2Q9.Dg/_5H(ID:CY\OMIIDH&<;dLB9
I>07KZRUY;JggLfU0<WFNC8<0;WdPBK>FE_54?AWTKE+&9M8=b2ZDKF.3.]@8=.X
RgW]L3\N5M[L(=,(Q[]?+IZ_OE4U]b@UYg03@^eOHD-N8(</cGRb-Me>JMTKKb<B
g(B,B0:9D6)d(=9[<g^Q1^E(#0Rg@I=].B=UeE]0B3]LG)7/Q[>O[e/88@4,ZeWT
=1d34#AAfdV(4:K.C_01/1P1C-8Dg>_gLL2ac,:K-2J(8_,H?+,CZMACNdT/P2b)
f_F^GVeYb(&>\FG0[-,JADQ[9<>J=O7YQZ+X\BMM<:2^-GaAX@)FNTUgW+._C/RU
f_-<=#4MDF439;9SPPOAVdJ?/T[)S[J^@(P&g]RCWB;KZ9U0=SSe2cN1U4R8HaX&
S(YV3D6&>>1\<=WV(@Z_CFI6&DDIJ.IYa5H4<UX-POC?TMg=0#fCQe=I8PfR@e9L
3TGMEeE#+#cH\JW4XA?MKf259dT/1Uc5]b9IRVXR(V)S,b>7Nd_.5f(=#[)Y1.VF
N:U?>cG@BA@=Q<DDZ>FPF/7)NPA/(P<_Z4bRV.QVBX<d4g(8A@S8Ie->KCaBH:)-
WRP()^PFAP_TGB00B_LAO-&B(]HSSMFV6>?f#V].@Z5[OQ@\fZ7U7MA)Z(TaWVO0
QP1NW]ZH7a&^<B?:DAQ)TQQOW22>^\VC(7^P0VH_ER:6+Q/EBJ3a38.\/N6R7Jc4
,BTgCcEH#680Y#-@]g4;]Q?^YLIeWUH6FL)5I^97)X-WJ#>R(^4#cDKe+3U[HB1(
P2JIM,K[;?8D=6=3SSOfF?d9:E+8ZHT\)1&Efa_SH&.&#2gOHNT;_aY;@aCbgO30
ONDARg8?gM:4TcaQ8fg&Q6H#9LSU@(P(_gEHcfFU3_6VM\Lf1(RU&B=J:;K\;+(9
X]3A&HKSR:S>TR53Z(ME<O&AD06U3V4N+.X(=BUNV\0W6+4,VA<)d/\UM(7L;X=O
](L?SOf)B(Y\5gZ#XHc(R5>a7)N/</K8MZ=^\92Z<09,RbfY>[;SLWH:gFa;6cHY
U.cL1_7S.H\^R@JcFY,]HcCX1_LV@,;,N9Kf1GDbE0>#>0EK4gXL72G+-C8\:RG[
6fPP0UXTB#-1?DJ5/R2)f1J=#28gc&<K[5dRX0Vc^GMB=XI^-=gEKZJdOG#+4<D/
I9K_BI/_agO.)aZ7/d[HNMUCPL6-@05KGdQ(XLUFP[_<W;0O.bSQIRHRHL[/=5E3
[+Q,+GHW3:=g25c[EO/M]MWf?1Y=a)fPaYK^6=HB5U92=VA^gLLdV@CVW3&(OdI^
M&L\.bXb<MPD47.3CH3V+//2N1EFR,POSV,_O7Na^2&B+_IKDY6bO?FZ@+46GC1K
C=/PfG;-.I.LeM4L[K,2#f)S:DZ45?\b--bF7XDM<dK]gNX]YXgc0b\U?U@f,g/#
G1I5\^,;EgWAb;7a-=22.Q9=aB2D+^W8Ub1:&D^.S\G)@UT8@J)<?7XMK90B2CXB
PU1?]XRE5<]X;AYNC7I]gabRW6PI0_()R5YR.7f>(9)(U2^4C.c/^PX/b_dHa9;W
Hf?M>L:_LcS=7\2KF;TFWPP[U)M\NQ5D4eV>c<AT?EJX=TMEWN8#BR[D(cS6=?K>
-f\=&RPIYYAW;YD5DB1<GEE-MWaNT>RdI9aS[cKbIY[,\3(9U05^I)gG5>VJY#Be
45#a2CI-CQP[CM<OCR&QG4;b]OYgSf\V96.g<64UbSa=VLUN-?7;V@6RHP3J.UK(
ZG+:(7+?PBAQK3BVeIK]]/3e?aV97<aG82K/^I>dY8_6#2J0<6[.3VFZ>P-c/&YF
\&6)J.-e0c92bEUDA^\bdYdgVN^a\N=HH)78ZeD<f9b)&3VYEQ0+Ggb@.)2GaB:V
\B(5W#+2UT:dbA?SL4ZNEfJ0G/D)5)611a[b&8CagK2<+)F&],6(=fFf9-QX.83a
/,GgC1>(WDGPW5ETS4L.+].]H4#JN(ACAC9OIaOTSGE<7,8g6\PJ=F5KXCe??.N&
X^[<:X.K?I&140Pf168Z9gdd2e#ZWa3HY,=19W)UA,ECT3>64W@UZ;Da7-14Q;W#
S=3.b[0NQgc.8K0+?O?:@GHY6G+=e)faUe5b0]C_b[<8PM,?#E&LCW99I^Y3H@0:
F/:+[+\(.&;T(N0ALFEfUF3LY\WFIT5[VU,G=2cWMI,25e>L[4T\?=71,;U@[QL:
SH<ZIbb[eD<Wc9H@_AFB3gD=+PBE1A5:?[S@E[:/a=?\(1++e/OG-50945W^J-Ed
Fg9eIbg??73e[V5MP&V[6/F(_=Tb^ccS#:)b:c)[FK[8SN&DX&5d_,OKB)&.@9KK
D.5?bF\.C+V_IPX2?dc6&e0\VCEIQ:[_/+^Yc@_#e;AX#/_=7RY+f=/gNXH4e2\A
SX9X,L5754#.D7\0\/D>db>C:WTe5Z==NBXXORbJI-a?58f;AJRB0bZb[-^Y-E0R
-]W4YYGZN^X[^6DTCaLMZDee[X77@>TC8:YKP]^WeW0KDC,L1Q14UJ3YG27J-M=T
1.1>RFXJ7<5=/UTLG9KZMgF:(84]&[fX0.CW0?N^A1b<FNQ67,#_D3@=VLb+aTdM
A)XH,E?Vg@OB+ZfKGfR_P0-bA0W>6RVALT2CIDCeH;IGJ7gN;C@4\f5O.Q?KN5XD
,g>b26O30VE;gEX-6\f>C5MA;FS]=3X.aQ=UD<a@B8Rd:Ug]BBTB:]KgU2-Jc6J(
Q^1Z8(>[)0?/dc.^#)GAXRV-b,#+6H,:5#:_#<e@63P]?gX1WYF_g<,@6+4]37Gf
U^KOT#9S9-5UTEC;eO&A[4fVK^DaF.ag2OL);=&N3f8Gb4(egb7&&_3[LPO#6F<4
f]V,2WU88\X@5SaJXL3aT>VDf#ENXCbV=eR6L0-Dd>/MS,QBd.=MZ6gZ;-NT=0CP
86HYBQBLfQILMS?aT-PR#bO6_IM\/F&dQ]T,bEC/f:T9>?8^COYIM4dFKH7QdTKA
Y:Ke&7f</G.I#P2\M,2WMC^@)bN(/&(6;CJJ@PXU2>WOFJ[KUPU_[J>^^MNA1FWR
LN0gV6Ea;WZ\6]JJN3JBbEbYG[7&5MFZGOK0]=Z(gW];IRWX:WbIX;@^KV9NY0]Z
W0>XF\#I0VL,Y<^5T8RUY5.Q7#f3/;Z9e0--BAWB,.9HAJ5gT7Q,D&6I&TJ5APaf
Pf/<@EIB,SD8;FQ\UR63@7S0)c-=BX8IE\@[^LBdBJ2-EIPL(0M><04I@.2c[\a6
Ff>HS?:(#3@B.0TcVIBNbUW)<^VH)/(UC4Y8)3eT4efc2VC0062H.X.LcXH+Le_>
DAKGJd@PPU9&,L3COOS>4D]D0cEQGTb.Bc8-.IWEd1G.G&#D=P;fA.UI>?ZLSb<^
?DUK>WH\>HYU9DC>D)#XN_]4L8A4L.=>BD<LHGJ\/PDVX4M(NQ>-&>.f2GfHTC>e
I>6(M.a)96CPJ[Y0T0OA2e^<)GG:4@HA-U]a\FGEd9#IWF)>g932SEEA_:2,.(,P
0;]C&271BZCe>g9E&OX1BU]77]YV48X4?YMUJc04.9/(9.4\0\U+d^/.Y\@HQL#J
\DC;f\f)9+QJL0JJ.[F2)JNd0TXEg(JL+3b[)#08E24Q6EG^39eC;?3R]b&FZg^L
=-+NG;HcKS(55^9Gbg^RO(&(Y5Uc^TQH@0S]eWI=.V[e1EfU,1E=G[7KSGQO>b>]
0ddCZMT+@+6<YP0+L4NVR6X^B?J7VP5[=:[;JK7,KSP#D4ZdBZXV&>:FW@Bf1S-I
F[JX].=H-fB9S\E5gS3b[UAF/fAW5(9A5([N<2,^#057=Hc)\OI\NbY5IDA>XE^/
b8UM&HBdfg5?5AFYP=D>AQGP7fQ&()(D#>e4,2VWK>L_TGPeU7F4Z0GG#LYa&\gW
(]?HC3a,4;fUd:&d0GQMFc;UYF[?eDO2WJUS@>HHFW;MU14O[?0;a.@R)6;)76c&
9\E5eI8V^NA7c1Tg_a8VWOfeQ4GQ^9aHQ1)LV6eRR51YS<U#>ZWU^.4QFDA8:I<_
7S7/#?EIY,,\SLY2cZSRK0CVY1KB<GXdYd<Ode:B-B+/Q;T^8[EV?DG@bSfQS6MC
6O\/86=]VSE6:fZ5()/a&C^QRZXVT<a\PCdYU=^OH?UYL=1SbZ@C(#P5.-&5+B<3
fZQ6G)NF[+IJ^<]D,L2#/b#--U:gT#+QTd+OKS]Vg7_0F#+=UB41;M4S419^]3==
0a?7,@L@V?+)+@G?M[][a2K+8WNeU)QBe=.@)L]D(C+0MT(&NXD(TNLMH66=^G#V
]NBPcZ?352_Q+g:[aV8X;.Ig.CG3-=W)D^[?ATO&,Ld:U(46J+41UJEPMcD//I;?
#D4aQ[S@b<P4.a#;JR37I8_>IRJ;Le<7F<]/ZEM_-<5/:I\-<B.[WKKARX2WQ<b,
5+:bX6<R8e:R=21.X;?-)b]Q[AbT)c/DT/I?C#H_LXX1^Sb8fg)U>.&^CUWPba1=
#ZD-#C6[OdF3TDT<I#Y6/6SX&+GYHBUeWC@_(0AH)Qa8\Wc,TD],K[03T)0N:DO4
F)C+e/K-ETEXR@74CEZA[<TOR?,1:g>3?Tg/EBefP@UVcK:]2=9A22bWD?.EGa0D
-.93#E^4-=AN\-EC^H\5V@M-Y90?0Kbg-X/,fQ&0U#MHIBb:PaT?f_,9)AHC]=-J
5\L[A(A21HEF,Z3dHB8?RfgZS-bSJ5A\IZ-,X3c6PE[MJG<FR6]C>DK_CYIHZP_S
E[MP]X6bLB^1CD\gHR8LeEbAJP-B2.dWX?P@NDA1&=F;,,=2L1JPY.6M-WRNCPDA
]30KX&J]7U5H^c\?YZ+7R3Y&3;;b)_C)aKe4Q_]N;SMW#63Uf[aU2^G.5@KY>1;Q
W@,:BM,7P8N&+)U5^Q2aM<d9G0)X0,gRD40Ac[4J1@#T=BJeMQ4B6e]]Z[W(K-Y,
U_E+a&g<SWE#WT(:)H@aQL0Ib3Qc_<0R;Zb19L.?;dE>.>[aB&3:1;N;=1F7dOb8
I/>e>:E^5b=2@Y^5#1dOcI,/XJB5.CfEGaPM4QgH0:#;_^C@Z_c>PYG3=QK75XNB
3aPSS<+Mc\9\MT,Ld63>TT2,9FIg5)LSMKN:HC//Q.J;M^,?K=XBDd>aJ[+D:?G@V$
`endprotected
        
`protected
I-B7ON&KFK-DM-9WFS6[:2U0I0_-K74C4O1Oe4(J]&<SMUcS7>WB))=a7eg/GW1[
6[&\WbD]#[JA7Y<#[aCIZEU02$
`endprotected

//vcs_lic_vip_protect
  `protected
+F+(dG(Hc(3eNd:eHE=N;05gBef7HM5K,G1K[M_SFAg/4QM;GTMc+(cZ^Y@.R>H;
\]aMd?Q<^&I-.;_P80O<HN-(FF8#KLcN#dZRK-7GP0cR.3_+_Tc/cH8Q6XV,gZZ6
;=N63<VNBM]&L;\\I99Tb8=6<H[,3dMZ.KI;3F4:Sg_>O;EPX#[^Fd3,GG<1L=cK
@D__IRCPWf=O+63Z1M4W<a0dc6WX2@W(B:T(.3[8_(9L>#gVe=MdCZ1I6&YZOB;/
f2.N/fT&BaQD.,YY8?eee_?;JZJFg(GRZd0#e>=BBS:_GS[;\D<Qg#^W7PRNL0-H
c]g>)0&O-Ie[B+-)UZE?/XC2dJ]J/BCeP>La)K_A;)YX)]ebQbc4-2WGRDN5^8/^
5_W7[:LX+g,G,>1\cZP)4)eQ5MG;V.<HL0\K_8)]Q(N3Z(1M49\76#:#QHZ.d_08
+O28VPYe1C+c=#X68)QS5J]_<>>^I]_fYg4SU\4@A\O#@746IUfQaDY/f-U7Y&1<
.,P72-0aB@d+VIXdSfaQTaQd28M(;=eg?5HEGDTg@;NcO.dK&?SAXMI+E=,@6C:B
BV@2Qc0F;;fBXBgK.f?5<#6?SZTUSB]PYQC-3RLGf_gD[TdCDU,5,TDJWZ>:GEW5
/a[[-B=H0LX4f)EfM6,6Y)X1V/[J^H-g[\G4[Yg7^6A_EC_V5:3Jf\OcC9TR)]E6
3[IXgd=S@:9R(8W/7<<LXBP1V)a1,SRXG]=AYP;_VaR#=+9(2^.E2gPQ#,943J6&
?1)/\C,Z\1Y@(TT<F2G>2:BQ3=8)3#d&eC87B@V(0ScFCL;Yba?]CZ0VU:ee3H0b
2C9bf#D5T_1P>QdH1ZK?aJ=K.@;O;SYN0=EZbL_P;XM[HF-+Y(BN#=3]^[b,2:R)
[cF?,5UOS?P2K=[58@[g?OI\=^AV==M=6)]ccf&(gcU13:5\./0.\MA>A/]a#0^A
2g@(2+&PaJ2b&Y.(1&F-b3JZXF_@af,^9::SG?8W,S=::)f.EFC0d/BFgA_#ERd@
FG_U1(deTVBHIfdS,>,MfQf,C1M-BeUeXEWCS(L&V=b\8d-NCDTb]5J]UF:aK1&N
FLXJf1Y(5Q?5-e)5AVgD)G<#8,0(^91b_8;;a)K5Q(O[(_&QY]8V&Q_=,<gc7L#g
MC>BVHNMY&K4MLIXX9-SQTL@e),T9MLPd2LU+Q,.C:3=+;&5>@e#Ua_)4fK2T:L#
8?=&:9#=O-;cLMXf[92@Ra(J))W#+LAW(@gSgRK-\dgcgUdQ9/Y5gZ[58bT[[TPZ
0,[.E<J.B4X@COZ.3@HJOTO/,f9D;+0OI-\C;7ZN0cDH>ea\EI(U^41f2.R]_R9Z
F0]MK_VZ5)C8Ld<:cQ:]=?H7;gR.(^fb;PH]-^e^MfSUZAZ-5UV+2J];S/bOZ0H/
TZZA-:\1Q-_2;/&E9/?fCD(_8)XRa:L#B#b\.]UUf-Tb&)>fUCZ25&4b.@?:3&]R
e#bB@Q=TGQYBXNgZY)CT@6BVXLb21=YW5SL>#6VK<Vf3^L?P(b>X^4WRDU\?(TIB
1]=dP5M8M(9,MKZ5\V]WW(QFK-ObEBEV\2M&K2b7cFg,\OC9L_H7D]B#L3O-cEP(
D-@U&/4E31,OR,>HHM/[]GZ\:^0F7L;AfK1P8@J;=eb69KQ>+@@YTd9M-4R(9\_b
S_\#BHN]X#4EH4PebVA(=+-:G4\\8.&&1aFVE[U3<3>AK650>AEI+I^W\8#R;d_A
N(:d[ZIMAJ\Mb_T&TXCc=eW9^[83FM8B]165&6VBS-V#7]\^XfOgd[-.a.&HTg<d
gZ4EN=SW;69C_T0535&#+40\OU12AIB^J&O71aT[YM2+dKO=_>a\Z,aC4f7W/\<C
W4T,^f10FHW;E6S</TZU=LdLL)+4J;>CcfeP>X5g5]:U7NICH9XU,f=[UD:(X#2V
#J_IQUMU:dgAKD97M@Fa_@(5>f8^-]=<_cP[d+:,[Y<LG3[\F8<5,8#Od/#L]J_/
MS[Q4,,(,8W#;.eEgfE9A@bGN;bIT\[##e:H>1+d\1f1S@89FE3?<Ib]865<E)Z&
6(Z:(>>J(+(RV6G/\AQdZV([IfJ^J8K?2A(+G,8Z(9d?\_Q97USa#J?ZC_eSBQTX
HY&;1E4/AI>Cb0\e#O5aQb;EYXH2+[UX9-d>A^Cd@U^fB:K9\cU2fWSef1c^H_+)
\XF[4:2_7UbPS/2cOFe[f5V._VEa+7-L77CB]@#ZH5fMN&:O&8+eEW4,EfHOMB+Q
Q=Ob:^V1(.&:]],:dMLT)#OOVcK&SI4-T&V(D[/Of]2J:UH;GA1]<f_<W4ebRVWW
aGP)T>7;U\6#Y=f+O7J+a#BbI?G#.US7<D1C(;3<HH#I+L\)03Nb++1fHHJU:/CC
].]6#\X80]-d4(EbE--g.+bOJT]>@e3/K2G4C?/Zf/OF)C4Y4VR).6;Pb:Z2HCKJ
0VF]Xe#f>G[A(J@Ib5\[^VXQ<R_MIFF(8,8:4OHId:_&F2K7W1O@UZ]c[3GPEF^S
1+H^?G<<SEQIUY:L)F-2Sa=S^N_.00CR+WP^McNgMZ<T^M^K6ggbF4-0)S>#<H5+
)Sg4&NW^7+MN.U9+Q[d)J^>+363WEe)[+_2ZHHdZ6V(=S/KOMYeA]N]8SS_gBfQ&
-d^FQZ.M]EKEF(FacEZ\)59;/05(fPMd=C8>gSa?PYXc-?(5UfTS3^I/B#XcaQ1B
YK:Z5&Q(F6eVHVB]JMA5(NEL)2T^5]H2[X(+(42V\4[ESXb?RIaM5K)9D_7X8bW8
C+UOWb=A3MFG\Ja)YO?&12EN=a8C84.\:.4^567\3]O(E+PaXJT-Y]b^A>fFWaT0
#)?R4+f]RI&@bJ:A9-cO8LS4XH^H?K17CQg\\BRNEe:3;IeeZ\0;N_5b+f01XRRf
:W_7OJ?TG5+8C_O??@0JNP/@-T4G?e;C#)KTf>QF/PH-0,CQZ>DLJT9W>?A\,I[4
eNRPVgFA(7D/3/>Fb@W)+<^c#Y[d/LJ05efIBL5Qa84/L]B,b/b/9/8C#Y;D/UX#
Zg[:180Y/NN;[2&B6@R3]CYP4R(ML:L5<24I/8UM76gd#3XZ,:6,>E>]NJfYcT(e
IO6>U)^:)PD]9CE(C,O-e74-N6Z_5LHZLeS1?0R/3YN_9gCQVY-;0<-GJOP/MWUe
7NGO5Y)aLD;(cS\=U?ZFaHc?#3TOULBRdLC0U1V)LDJ&e]f_Y=ZPG(07f,f9g7;N
[4_:])3Z(4FNafKT&b,SZ03]0EU^2cS849:FFI_+R1dge(^::.AQfQ-A/X,(g>0I
.SDAc#g;_&C>[C03dAP7G(eQ2=\RW25X5Y_5=8_5O/5-M9Xf2H]/HABXaMLU9FQ)
Z.)cg?:<SR8O0B2dK,07H3d_9DTO-=D&M7Ke3?K9(Ec07(,e2.Z&M<;MPP-fPFMI
_.&ELHU4eCKFfIZ7MX:(OCU2][Wg[ON1[]VL^JdIC;LW]VI^AZB)YZ&9Y+2DafM^
XcR)2b1-ZW;/>S,]L4,5RFORe]YSHP<P.-Z_6C48_5KVS277O#/7^VX<1a[VNNN-
I[(RST2dCWbJ;.;9M<R_9PLAJ&[(:SJHA\g^c6f>X<D/#E70aTN53LN7ZFLeU8X9
=EARf7,ac271P&-=8#\7:[8WKG2;8bZQ^];=B)R2df9YXX)-F)D4Cc7bNff;J13&
N?g9:2?3]5==F:@N:bG[S=,ZH&N1/?4:X2M<;T65)cA=VGQF2OEd0-fC+If#1.5D
ARO=@K1eA:C>9GK)Rb;1QVc^?:(a9)QRf])SR&[Td#fD-/EO&bQ5f?B9XKg-05(1
?Yc-Y,Jd4DMZFBH,#>RU@,_]#J.CeT=Y0UgEUIR-B0Lc9-MVCag.>=?X8-9Z\6-/
R5+4;:2U(D#,Y144f8:AJ(d13F2RB+B0+GR+1#=P0LLA#,-:3\0?6C#IG,4FCG_0
M08->e33VIaTEI9E,_19,S=\+Z+f_/+295(fb\b]#d6_fSTQ0<^#?\/Rf?(?VaMc
c)2J\f:(BT0e>5\U\,[Z_LdAN@C_B>>\N)gV_RA_.ML6;X/#-#&>=f=Q:C7KePE3
H>PU:A1b6UFK>8a2WEV/Tg8R5W4gO1\V;C4F:HFe/C<MFIfVMN_MQS8a93ZVMGR\
7[(DMYe.=8.]_QD[OVc#cYF4M(^FMga9bSU_BA,IEEB=GPQ7:AR2RHD[f618(C>W
MN-e&;?LgC(1U0>PFH]+VbKR^e=U@@YOVFX(LT(</1VTcb<FXF9T-aA-;PR2AZ:B
&#RBBEa8]PJ[gb.I7K#87#9[eeZTSf4]D1&ERJ_aGJXRSHg]1HUeMZP0c^dOb?B,
13WVdF+=@&X4QC^b5<C>4OY:.9eLKH)7&+1X)AH4?8/0@P#:85eB\6^gID@Y-f,X
(;Y<7D:;I2][(ND&4R;>8f0R=&35V9Z8BdKITAF#A5SGE_G;D[2P=QBR@bXTbX-e
0_AO<gA6;cZ-8D9UbY#:;eFO2T&?dNM_U46&N57@8(W@L^YFcB7^CB/:9IO7XR<M
0;2F:718=R-Zdg]EdMeUGU\^1D5@PYYAF0dH>N2e[.@F\0A62A=IIbN+&CKZ+(\O
e79]dc:I/L-4ZV]D)N](CSI<HdY0MD31adT5RQ_-T@TK(>K.R2SY95BGd.<QQ5F+
EDVNWc^aA#ER(Bf=Qd3b-f#Tf3eZbIa@gTG?<[#F)LYAG,.CA[04YUS&aHXL\a9^
e(RYDaX)OBD],\b17&7UgbR;GY^URT@K7Q#\K?_IBeOa-b^-@>VW7d+X=;505+KN
,\F#g[fc[YgRXT+eV#eM63VeQL@LXJC1;A>Ace^JV=4WV?R>^4ga<Y?)e1-+?Q02
(=0+dUZQ;Zgd&29I[#FO\L;,OR4K3ZJ>^NbNICgMDCRZL</8gZCfDV\f_E[C#eP\
B8QPB#WC?C\CWPKE(Hd_g@f^4YCZZDGdG/aDdUFXQRe8&9TI;c8CG1V0AI8=57V5
;^((d8ee-E9cU?7a.QE4W+]f0H-Yb).YQ_]f0^1H6V_7HbZ8UfVORb663HKA1E-B
aE&e=28@R0/(K>\T@3LL5>Zg,T2&M\X6&@c96O9TBC?#@;&V&JcIf)c+<G\28dWf
:_LbO/RQfK1#0-.1(T_C-D68O0L;DSKUf/KY^X00-:.=?,Dc\g(#&WeAFDM\fFES
R)XM0&K1HO7?>6/K&WR4C_FAJCcNY/gJd6QS+da2?[_cbZ]<-U<^2Q_/J5V8.b<R
B-9WO@>2XIVHL_4[-7?\-(g15b(K5Ib,QaWFef?f@&,9C[54HYJe]b\22c+aKdDB
3gYF=KHHKU]]9ZIF>-9c>B>B-MF.)_>O?J353cg=H/YMeT+-K<I;?aZNLTN?-QM#
?:/(.A]7EA]0I834P.b;5=P?P(V@MC8/?7B&S/:(H9D(Q4@;OW;72.\>HASfX5=C
P>]N>HU<EdT+S[U00?DcAd)OeW1FePL07WCId><?+=#)\1I/d[<cd^E0E&Q-OD+6
A+-V]>CUNG&/TWSQ))]dBQ.,bMgdKJKK2g:.Z-@QCc2I9,VdP+2##+=/EQD?H?DY
.=:,N?A>9eIa7TA49V5#P8T;ddSA-4M0@N#N80)F7bEN(>)cQ+LNBYFJ<Jc#_#:7
cF&,V=_]W[,4Bf:FTac4a@^b^?>LCg&6@KM3>Ke9I_B+#OGadc;:MU3F^Z1L?bDL
<3E?.-\^IRN&=@AFA0R\7=CXU7TF97bG1KfQSME^B=BXaX/GDabg1dU9^IQaB,&=
))>#D[B+,45:#/0g^0)4#?+c5>F/g5\:HWK\MfT,RfH(Z]TBM^EXH[BXSa];-4-\
d57Vg)Ub)83^8<1Q+^.3V[eUf4P]J1NQQ&\C>)R@DXCT31=6S=b>(38Cd<GZ2C-L
G3dU8\cMB[7FUZ_3G1Z.\R\5Vd=RR=7,cg9/T:d_G&Y97JY-=:eS6N#09OFJK6=R
QN;WSQKO)^b9K.O6/OR(CN/N9MeO\5PRC/BT4+KLJ1E=cF5a_XH-NU/8;&,V&]dW
d#(Cb<+@(#E^B\OIH-g#TWV]Od)4-b/B[?5.2/?[b)PQ3SNJ^I&P#eJBSd6<S([@
BR<(^@Pb1b98F.OQ-UXd-TMG:^6b+<F03S9YQTOH<<#:Uf7CDT7a-c.:GRL-/VO5
QLW_+0bXICff94U]LVCZBPVcC<<KdFDcL]LcR(1>,;BS1,e]M>.,N3SJe_3([QBH
9BXDEIQ&@aFV/dDD;N[[#^+CPSg\2)?_06\4VS8fRN+([2])0(f4YXQM6I]3C;e.
[4a4N;I&>HZdXK6-&358IM5KGTR#4?Naa4],f]S[YaLeaRUcRea(dUANE2eF1JH3
X6_GJVRTQ2.bI2Q?8)FB3;#ZFOJeAL&2Nd_7NN1d5MP&UJcR69HFKZK5Vg.bLaJ8
.L9E#)NN#fQA2GUcT//AK[_R7MVJD:ZHEDCgQ5X0VNI-/b9Y^V_K9K:B&1[^,MSE
5:F:f-^GaGSY.g=Z/\)GeKGXU5f##/;)7;-RA;7CP@A.-BQGIaPP4CdTU2TZe[f?
5#[HLUMXeBH)+afeP,+36cMXBDae2WI(>=/@V8KJSg(P-3P9f5PeU9eWM6-V5fKT
e1N[\_.=\R#;(+\X.1NJe1VLe[be3AdVYTd#U38E#+C:[>,f\cDVXL;MO=J[^:-J
/Tc+>39MX4^>N[8QC\7e\Y#Z/L-AHP11;\_d5SDK<;TM?GMK;EO>0+KRZ,JIVb#Q
&ZTb85/0X[3N:8UK=VXH],/DdTE?)]UGa;2<FNR4>SVAH:BJ@;RZ<88gM=4/g:Y1
36(I(<-SDMaOC)7[]<7d#KQ,__NA>1XKG#^Md_GPS=W34&FXKb#HgQL.K9e(GNf0
=W-X-79/7MRU15(58?JbNf1gf/>FK-#3XL)R;62<X796PKSU]L5^I=<-6XNID6]K
&^@5f8UPdXZYYJ-SQ/>6P<IS#?<&eY87DA#15K;)B?BY.W@81JJJ(HGb?IKKDH:2
]5\_C(c+U^1Qg[NW/.gFWcKYKVM]H/EK=bXWG;6)P,:Y>@GFB#3KcGf7BBb#+PC5
NUK-FdLTK8IgEAW/E0L[EP,0YR93>,/]@1:F><.IDBH,7feAR3[P:Eb:.H+GX@=]
Z0VCQBNQT@)G<5,.a52WJR]87ECL4?0=:<TP8VcI9FG&YUYJ][gXXCYBGZZH#7A:
,87KgNb#4+[YR<TR<IR;B5AK)aM,baMbgaJ#\UI(+B)&3]+?P_W9A?_H9V#A7c\W
KfKKfbIJGQCCRe0Hc/VAF17LL=Y6G[-FO4C]7Y2GYZ</EX)f0IGA@.eP&/TB5]N>
_#dJSJO6T;:OHG?HY6XTO4]V<=]b@13QVN^K5a4fGLE3D,+GdMQ?#HK&/KJ+WI3T
C(D9#LA3+ZW?dP=2>F#8dRBf>e11H4DV)?8O:?:=;IQMa1OCZFH\e3<6-d-#[5g9
L5Ea&dbZDABO&S4#g..K,I8&8)a8C/\1J<0KMeD_2C2.68V+?\GbM2=]E443B92>
ca/e2==)3YA6^V].L:U:IPcML:W#X;FDJ<:]7R6.MM(aaM6XaX&I1^^5=/#44[[D
CI]36@=B)9O=)ZE/W/C;.Ic/4C1#?:U\X2;DJGeO(E:>D[g^/=Z>HT@/FIWbG5f6
AI>.W/FP#3Q.bH7URW_MG,+cPEQ9_5Z0Z_Y)cGK13L/FF)#Xg39#H4I23?&ddNB[
A@5EO.a5C@7RX^HdI-WJV#^]&)aS0gV[cBBgFPT8&bFY3GBY5O=9L6B.+63,AA2-
8@LQH=Y@1G6<c:2Nabg2N5;X>4VD<:B2DP8;3X5P;B&Z+.]3S:D07+d3&\<f#T6[
ddMR2gJA4JK5YBT)[1Td>X2RE-</<5111.>\;M,S@-G)gfOC)H30ZMH4g@Jee,V<
NYSPGDTGOQ^.?Y?3_B(N2<bFY<R#^1Rc6(S1D9RXKJ?DA1NeGW1VL)3Y94,;SFYB
EN)?GYb@aUC:]5H:?.9B,K\4>a\O0cV?Z>5SHe>OBC=_Y)GX4/A.ZWf]LdRR\<.:
_+KaeL^UJf8.<I#3bLbEFd,Db1];&f/K:AL:0b#YeTI_?W9&cXcXCZc@5Zc/a#5T
UK&f6LJ,)H)aWF\@^3OJ<8BLJYDZTHcEggOTMfGFaHRQ0G(H@3@2R,87)]>6>>e=
[71cdDY:BXEK;fd_Lg5B2d#f0e5SEKR>Qa;V@0&)=UK]8:VUI[_<9bS59>/TQfGZ
>^1)].F&KU4UJ2UBPYIWBN0Dd_MaM+4[^XYSGa&3TC:-)Te@4X^W)E]KF)d6Y;-;
Ke//f#@9R9XQ[MJJ@2>L)@^^T=2;O1eAN-f4TdX6cYRF?T2C.;_RZ6=:I]&eX6bc
SQS-,5?cJX<.A1H39U;EDQc.H@G^de,8U-5Ke\WQ.ENSHJ00IJV:ZZ8&)AJ-KUDW
dA/U2=4c6/R,R8J\77f52bR>^A^)/EaO9B^)K]P^)_MeOUXOE8JL+9_eW6I=5J(O
Zf4#>7W8Ffc1eF1@5PS1,SZ.X\EL(#f=X,\>PFT\L=[TMP+;FSJ@JIG..;<DWGPY
F.fge2[(Q7ZDIPPT(HRZIMaMGYF@@?.aMS4VbJ:g+&QS=6d1\)>1&V^G0LM>]+?=
?a(61T#@^^VaJ[,P>c=UJ?[(=UV2E@^=6<&#5(TF\BeXGcEQ+Cafc?+X-=];Mc^g
7c>6A1M>#:V@b1=ee3cL<g_.f62OO.Va15J<2DK;/F3QeV^)T;5Z[g-]J2Mb)H&G
5d=O<I?E(8.47Q\eW)BU;VWD_0;6R/YD>9N8Db;f.W(#YY]fSa6c.Vd^I9^c<#?e
9cV6>3+e=7JT(Y6^6([MfO(ITd#J[L5F877)ZJP8P[.=;_^HNC\BWS0,QK:DMOSB
XKX-6e,?8^;JGdR9KD)AC1762WZAdC[5L_+&D(aHg82;QB_W7?fF@[=#PDHZDW7D
W+R<P&c^WB3I\KOPLR6O(1QW>SeeHDX/AVVg1CE8-/-XDN,7>C7WPf5daPX/=BV,
M](Lc>GaWP]]D/<U?(+c0,09DEe_Z^XCT9HM?&Ida21;=\9afE@Z5^6Ud#9f32+A
T.,1c/_NaT4?WX3N>:[86EaF[5RfSc699bLP>.VG7[+YAG>BO[2W3#_DM8#@:Z8T
4;D+e,6Ye)5T,A,N7D)#YH7-]MXff<c1IUNB4F?\3c#<bT./U66IeB)&6bg=b@aR
+Z8B0:XPe>0?3]=aIT=:aEbd2.PGWW_\(g0\b>b=.aa?T-Zb<K,ScY-<BaG62B.B
GO4B1SVA&GdL-QC&>WF))XZRW-S)X(_^^A#Q@KUXY@;;)5UF75.MC)6VaTWFCcQ0
PV;O(-;aZ]_cYO^V[c?]Qc&8e<g6GVFgIdHJR([;f./&:UQ+f+HS(DA#_I.;Bg?/
76M4cH0b2Y;R.SWA</[W;JXE?4aM)/,?5(_>WH#2[3@e19Nc_YcSdY,.@M@^]>UC
5RH&g-7+B9N@]@b7S9D77/>=gcQ/77K-.KJ/ENDJ#9X<V_(&.)]RUSe9//-B.\Cb
I:Pg][>e(5+2G?,a:\0-6\dE9AIHV/U7_3,FHU2_#d@:9+T]-IC@?YH#,E;^7e[4
7eKJY6X=L/b85_43-fS1_9..IMOJ6&=UDDL]7aZKS.5O6HI;O)&@a&/JIHB^=ec;
23TCP;g7JY/E&ILL.]P[P;UJB+M[AY@+5O7AS?>#0&99;ODAbbQe]G4Q)L,X,.A8
cc+]K9A7KYXMH<7fN)CXdP[]DR7HC<aBB_^PUR_-?g(U=L@VY]J^aAA1FTW7X5M+
-</WfAcWMINYA>=3DBPOfIWIB<]I1LV/OIEJ(^4,(GU<:F9Z>P9-bT[g(cd89/dW
UfCA]-L?T=X1AZZ2BDeM;8FcKP=^\_YM]ERD3N6E;U.GXX_[M)?>WU.#VZ16T>0H
4)g>P[6+RA+_PA_a>I.JDB#&1IcfS_QEXdW=ZIP#C/RE6>;&X9(+]9<c(:JEMD]K
/]ROR(@bNGR4=Vb,7X2R;aI3c&_#KWY\);UdQVXM?eCYKAgFTIeMS@a-3.Y;OBL;
J1c(TURY:AP[<CbZeg]d_Jc3Z9S<KPgO8RefNc2=UX?<PBHCc&XHX0D\A.CgHGXJ
?J,L08L8eV-\;7O,cM,656?Z[2EbWG+c_UI;g8M>=e_78LOE84J_c.J+cDJU_SLf
<A2H940#U?cRZ]JMS3@N@9U8e[YbS(b92G26L<?>Yd<f+AG]^fJ^>8aAQLUC:8>?
a3)/1][.\e:7^L)K(@/+GVTfLT9;2>Ac2e#Xd/f3&9C9[eXR7GAg/(81/SMK8Q]&
#6Rd]Q-TRZ?WWIG^=8NIR)Q+eZKBKX+fPEZ#-W\=CFUW(?.HP#(BR?V_81-1DR^X
2;?:cQ+N4+RCdH>,66SG@\\LQ=DRGLIG&eCV\OPOVDgf++9/W4d\WW<BYa+\3NGG
(.4A,0@@VU@b_IE#1^[W:H>=2VEY]CIgS4OFTIc\L]1e^ETVgJ:_C[-dSS:3H8C8
TTYW?dX=+NQKEIBdQa#NL37NZKQ[@8,VP1AVCa,6<(@3BVfe:/Fa\-4J-+fXXFB_
I?.b7#0TB+271=aP/bR#CGc&@=Q7bD-<D8B(U@]XUCKXX.G-aB\CICfbePBAU+,M
_]9-A2eK=HS&Z;fZHU7?K<APCe<GRIb07#-;2Kb>+7fA-(^JY/,W#BHL_f<OR[#\
A?N)?8O4#dV0)/\+T;HaU#55cOES<]\?0JEBB5JY)(RS+X@^WB;BG.W<d2C1QgMW
SF<[(XCeFR1,X7[-28Hf[JAW0bF];SK&Z3:I>Z..cGHZ(H]#_g<9?D__(5<Q/P1J
-Df=3H4MZCLNK4N+O=#e;6V2&>Q,(Q4gNHC/V25+61(.#).4;\&JVWIXRG;?5]B9
#VM.]HEZ(#[T0?=LO4-:1UIDJI/PT5K>+(RDQ-0VFYI2>FT2X&)J,,QU0HeEHR-S
O\Le\[QB[S29-6eNJU08#T=JOP85L/^];1U?;;+5N\JY)P8c\^D#O-.O@2NBF[gZ
_LB0YeNSWE?UXgB1?Jce=6>a;MJV&WQE6.CMDWE-/1LH+@],/QT8LPU&LbdXc6Z1
SW)N4YWWMB>.WA>Hg5AX0XY_AI\<=(:<;26C9ZBEXIPQc7:MS7HXY;7TgVQ,MN\a
-C8bSgKW5H@E3/,ORJcT5O\e2_[5/A4&@cYEJ96].^/KG9AXV7M?P=KM9?G+1_#M
V1T]5HC)?R48HXC<0f1AGHVEU<JLL1]<&Rcd,OQJI1R9,O3^;f0B<Z]?/98G\1gG
X5PVLcG:^_I3e93K.^f[;cFW22g3g\K8:C1((ZfMUO8?)1E_G2-2IECBNKEO<@aT
24A4^UH-d51^B1.ESH2B8VOIHFC)NcAH/[0>V)2_B<HJLL5<#UY+WZP-JS/V^DKF
Dad7X^@a(4E8-^HgMcFB=[^\UUB/e-&GBY-K4MgN\>+:<gS@,e+66FUQ84[)_MNY
R1:8?D6/dTQ>J&EK2O1CbcEW:]a;#b[?N2(#FH=7^+ZDIEWNT^AS#0g1E7dgd4#3
_Y&])VeTU,J&S(J<M86#JWg=/?G?9)1;P5a1F_OdYT^>B:3^ab)&&.49NIHO#bJU
daCd8cH#e(gAZ_e?7(69b4.0]SG&>:=FL^Za51Vb>f4cXU6b0/([.Lb2J[SF7DJ2
&OE4]c_bQPX/I9H&U-:aWPYAd(]g8+1T/X\1P9\QO;1LS;?QdH\.EL;B#+.GQ0];
40]a5[&Ld7\04.+SO1A?=5K3]a4AC@.ef7@C[N@29H>75JF>STI-]<@BNW3Sg;2^
-V?#Z8#b<4;9P/CE;=:dD\[OIf,UPSL;2HHB:IS&<C2TW61/?+aeaNKBT0]6U.N,
/0)O&2Q])RUf(Fa.FVgJ=&=#H;KL;_E2dgc<+Taf=@4S,8X04:D\cb,Uf)Q3(:L3
+_MIN^-L1@Y3L&B6L-NKM)T,2&&PO#U=TA657CA9aO_28eG+0,TQ0.c_C(I,90BJ
>#]F/W0[C15JT:2CE33ZA\3e;(XZWBF:8-52>QZB1R4TAF)U]RUA\6L_S.LD.X_R
J/I^5f[8B+9Uf7,cd8e4)5A090+^[H_53B1/&BCZKXff_F96<W5/B8),a0HKT8dU
)>L.F2F9H;X;CGNHD_NW--R;FLD+QYG94CdUE>Af@aAaZ70P31V]/);eg\/K))_[
QcbM[LD-g54C7YAP2Yf2K)^>:(BQe^7=D;W::fg,eRDA)2BWAEe6[5OGT5N>IJ>,
+?;JWP+.#C5ZK^,F(cC:6CU4@\.Dc+W]ZH.O.QeBHHB#7,\P@IF=F\^]/RYM<EMU
O7?)72M<IEH8Bc7_FP^)<eJTSKASB+,1A8=5@+W(LZVW2b^e\c<RZ@WR4a(P,=D_
BGEg,8<bL^VJ1O9@c,[.WeUL957QV1+JaUGHX&I0OBDS<Ng0\9WY,^,Z\3#:F0a-
6_-Qe#2<f6dG_7(ef]E<[B1bd#c=FfY@GD#GEgc-1WIJIF=C0.HP<I1;ab:Ncf2N
b+1YZ,.X?;4>)CM6FN7@D1U3:@U<D,eDJ#W,ScZG.cgWBWHZ>47XDV2e[^4YH,Y)
],<<JV>SE<Uc9M,YOUQ53dM#KY5NdIW3W0N]R3A7FfH#cP68;9If5^Z5J.2=eF@:
_#>#X2>8Df48->3Y2HATWRFdYR+Y=]5ad)=ZSM8g<R:_073(#2BV8OH&fY1AARKC
Q:KC6=-eIV(C3?\Uc=c0MFELBbUgLI6(e/RK??KP-TG<?d<@(cO96[bZQfQ;]6aG
cP^f[Q\3@TKY_d<077a-L1X[d,9\cGfFPK#<JGUILLcMMP@3#^]AD3\1?90V7U#P
]bMQ\D=gDbR&O@Z/111PQbg)a6#4_]\>1gb]+N[Uc>T-b,IP+NC>)V.B\\a3(S7e
S8-_04OV(]6)[M1PafH#B??DA2BL>F6W9R4fJ7=c<1R]C2W8:#]>B;KbX-G3aCS<
Ec5ZKWF(b-aPQ3QRZZ8C5<7QgT=-;;C/S/5BOO?B-d(I?#,9&UdQU;(?8;T:YZ/N
U->O,3,[.WSGY2JNS3R3-;a[^c0R;4&T(ZGV24.fCLZSb5CR[=^LgHP,9N[BRM#g
VDXM+Z&1)3&L.KW95^2bN4P>RA&T@OO7+9:>7NCfG37:&\.M?bN^Z(TP40[e<FN)
f4GcXASDg,QI8U@#b]#AF[1_G)(7G?(=cPD:S<)4G7>-O@bT)2?0cZg,=X()O)<a
]dP3F98U83M2_A#XO\QI^5D2Q/S5+P_B;Ag5IL3Y4d)>9^X9RLFV\.CLT<RT]\IS
=CVU_PC48SW35NdLIOA1f0?bb@U+<2eQR1aWQf\L8&MZ]d[./c5,E@J3W-?L7YKT
-4[Z8)I]9d_2VLgN+:(4F-<U5g?JGg+PD>bR#@GH?\&I9Y/C7BOWI0;NSRbfgA<N
-dFfLGKB,LVUXTUFF//P3PO.C]+:8D0_=,;a>NNORNC6N./6N(-gP01Q,PYeY0PF
SA?A):Q=[T+EJ#E[&5cDbDL7cW;/:\EW/N>9(F?VC(cZE//0fQdegWIM=5R4X3]=
IgU5d.#]G8]6,\QSf8c@?cD93#9@Z\JJNAL^Pa:WDaJbKY-5LWBd8QZa5,]3T:&7
2^0gfebAK0a39_++#.D/:a5G@&3;bSAA,e^X/DW;;NM;LXF6P[K6db+3#->IB^;/
=MC8RWgfg/HI13(g;\I]@:LX-D],dMBWH(@/b>-HH&,.CXbHLW_0Q(#Z93V7VM)A
+]:>Ff^LNcL\U(O5>?CZ+4#?\CV0ET]=M1>&VV9W=2EX6+V/f<[EY?f;,?7SP1HD
=?).9.I^OF.8Y<77T8EEPT?Y\?1PdH^C4T5;:f03.gJ26[<aIP<Q8gLYZ)f(gF8e
GM;(ONCHaI^,:)T-Z3VWC0>IV&Tb^F;F20JDB^GcT)Q8Z3F<C.34<5RFaJ@:X3OO
B7[9BED^d9BSP>.Z3PU64#b4KVI5,K45J@)#T+AJD,=YPE^;JD(Me[Z6[R3>CA]J
g3B8_AP<P6gV8Ba_QFSGE/cJX=J/g,LC&#C@3Ya;HLH=</eYR.;SJZA&\],=&OG^
&9C2IW^JX;c_9@(P19[J.84[7#?_N[Kf>d&OTKaX#)bb]7eZ@SC+4We;M+\CWE3[
cF7,_06]^?WB6[SNcF:C6Q7K#FFe[d_dHQ-@-g]YH[R^Xg>c[eV,\.fg6)Z48MW^
&B85G^TIT6>-&Qd;-]1:D#g1db6LNdAYD8(Ce].c9,Ad:W1Ka\3e4IYFLU,g=XF+
<&LeNag:Ug2E3g+VRJLS2G_(FNO<(4ab>GcaPRTA),H69Z10,,&ZK#^25&2Y1-XO
,H:-YZO,N<A=12YcBN)\E)-c<_.gCd)K:=S=46>=aS?8BG?#3NPL01.)0N^N<Dc>
D7CS:]_MH0(60bSee^XCQ)J,4eW&D+SVZ;X/<Ng&,\#^36VQCL1TA.Lf4,@)RDWC
Y_87[[NT2+gVS7cXSC5HUZ,N;W@,d>[a,@RCQfKP,Q_1CT8dC0D.)MN)C<7C,?Cd
^?3CI,T,cL=<@\<PJBO:Te3bR/JI[8WF#aDG0OUa@AYV<A>5M>\&6J1.T#YXIXY^
E,#9dIMB[_D#a5(-IU[/98HZJ4#gaRZHCU)]0SYA+f9E):\:G14G8#b(YGC#ZIL:
U#gIeUFdNL68RG7#L5J&ZJ+IAOR9?;@\Q-ZgNGS7#VDb=KN7J^;/LO[5JH]4UVY:
J)P#G1gb(O\OILUSc_dSVW>IQdg9\X5D7HfYK^D0QLH?+f>:8/<(^LLa5_+_8.7F
2J@J:21>W/KE)_YdR/.f8AN?cH0,1Z6Q-M+GG.+d@G7fO#\DcRS^G/_V,T).]_6d
)+(K8EYIT9LT;7N4.OJa9Mc:+,^N20cM5cXdRL50^#b8IT?)&UE]N8<=8/><HM#]
+:)>35F9/-FFVI0Q^dC=\VOPG53QT1.Y=0.TQ=2ZKU3349\CJ.B,]1-3cD2dPg-W
RUX=]7eT#HUe5FCUNc.NFS\./BIRAcZ)D)We)Pe-#[B7ZU4Ab<#L1e\K+VI1I6.I
#b+,U=.]<SRDb3f@c4&@_^(dY7R<5JB>->SMBB/eg:]YA08.;(+/I5PBdF8>cL72
96&BBI#aAO&VZ0e0I4::If3ZJ?-V#g9d8gIV&NNIDbc^R-22A5BG[U8-(,HbDUG1
KNSR]]#RI[gbSTL2HG0Q7@XI..\?AcLS]/@I]];2c=&94Xgd96.1;RN6eD/_4SKU
E+?_2(?DN>;43+L3#Sa)b,fZX/OP\HG,.^f7AC@dEUKWSXaU(,38#c+89H97Kf1K
;XULM_a?6E6_J&SU9E1.R[>gH]@_E]^EG>4JR=aI5C:=-(O=gF;a=OW(2NM/NgNW
[S4=gb/JQY+G#M7Y26P1[-0UHIdF7]UV^1.&>eYX\cGfC6BT<Sc/#15g\F</aKY,
?0CSTN/?,8YCH/JBK?7R;gb_4a_H(.&Z^Ee9.+JL=:^.XJP6Na99#8L(QXX7)NVG
eI4IU[ITHQB1-W#KXJ9;1\.P7RGQ>>/\SAE9d3F(KF-_\ZIN>SVd:,eZS2[<+.dR
HYa]@=Vd]F3D30ZKLOS\0/fM<N2B/#f6egF^WAaVHOZGeTZ\#P3C@9]a&L<(R:=/
M?2[4:S[QGQD53+KI<3RSH3fODYH#,.@;XZO2Egg<2@YaafG@c>[9gZED->D<\9&
OR2MHOOc,>Q34+,LJX.]\gKb)a^YM,3(FDSJ9X-]-fKN_:McDK]V(?^d;]Y3,?N9
_D4]2?NH/W-F,#B.A4&d#;WUYBX>HIQL+0UX>ZXfMT_Dc1B?dR_fF@Le07/4D[(Z
_F8LS@_-1.W=#0[[W]/>>N^/.R=gD4[S8^S[A=GC)Z/85PgdNN/R805#6@IAN2)@
-]WR;]cE_Z([/UZ>GC+(=UKfZBVgP)F#:,8++cc)H;+V@=NbN^]a,<X,U-1W,A7\
41#D:Xa8_G\+J@XQM:D8&62=#ZA(]6ZbSBFH(Y4NQ<:CC>_2:UB=K&FE(BL9R7^<
?C5d)@<&gSO9URNX\^MWaE+4S[H\03\<-#dZaPe_I],:[EL2ZYZaf.:SRQ2=>c;T
5=LaC8.=[PQ>4g82FC2CDMA)d:/FB?-E)RMaE5XYV9H62^:[A--TJ,0e[GT-]3ND
JE4-8P?+?,MH5bCZ5/8X]Ff)3L6A</6eeD1QHcHX[Q_,.0gZ<(VL5/0V@;cU7K[>
F2NQ42ZCRW9Ba4L@JRN\+,N\4K=\LJOW#\9VI1X<Me:AM/#T(T_@&(0OdZTXN&E#
\a5UFP<a5GcX&65WPIO6+QPLO1>BO@<Xd]=;D3EeNPS&)d6O.).a-N#@D[1UG^e[
F=G&1),)]J^J#b)^WJTU-03DFM+J2Jd](/HaMKVc>9MgA@b\cM24_gO]eFcg>E0E
[6ZAc&UIWR/1:[BQ.ef\1:9d^BWV#Y,RG426XCE)MD->99(<<RdT09,TRW3C)69_
@4aXLDa9OWK6L)5RIU_&WIU6FWW90-G,V2^66YZO:WZR3.b2^I-T(>UA]e6\)X;D
R#V4f(Q;A]8_X[[KZbR219]cMVeB9JaWaXM2OWO\Aa<<-F9L>S]]?.^1(a8VR&UE
QNL>9-;B707:4^T>14cBWLH\Y#+VMg6&<fSPN&Za-0c?,Bbe0UUfd5eVG#&F?=N1
:bJRVDZ36(>9-fQf>.c)bb=4#8=FfAKPM5TS0cf-MgI=QV?^K9XWE3OO;#+N::4^
L6BM6H([6V-FcAK1G_7X3G()aeWfIMSTZ<@Z^E[e5\a9<>ZPcEHaV7ZM)L.6cMKE
gcCB7X=4Qe.;e7?ESbSf1L2eWIbcSH)1XMX65XF&R89J,S;NdA/P8-c3V^^F\148
^A/1Lg_EZY<A[]Y>f]Q:NXP]Ogf\PD,XKcC.^KFBM\:M&J<W#&.H^&.\?<>NLJ8Z
6O<cK(fB98(?J8TdK8V?,LV6&1/#41V@Q?gSfBPQ7U=bBL26T\V7N9g/=@;]ac\F
E_/\(GT&A.aAGP9),b,):bJ@;.OLYFcbHgU)BZ)B8_+,-)&Y+Z,6,:AD4dL;SHI+
JI_KRb;UA5g[Z-ZRM,7.9?9\]d<?9gH_e[#B31cY&#;Ug041^GIR71:fPC3F3/,P
]ZB35#MagGZRPc1X(]bb(1TIbQ22b-YYC#J+.>95LA\R^2YA><eW.=TgC<)Z5>E-
&;Y:bc-WB,XF,_^B,_KR2Z#_VJN0Ac]#E(@0&?EMPOfM4?V+Pf@@E4@[^#<B3[N.
eg<Z0\2#d]eBeWE^@N8PY<;?dC0T2GA[/^7FRGE_8=]N]2WYL-e3;(Hc9YCV-1<K
U:c&.WQN([gd^eGd86M7A0C3)NH_@H^;Rg5F#IX#RVEd#IA6>I1e.DbZ_CgP,0<O
;S\;N=?=J6E@G.A@\H?J1CWCBSGQ98ZT<Qc<d<5LU4d&K2F8Z=J7P<7(aWU)3+?/
OR(C.(5G5&P@Z^5O<f\=&E?0<>2F_f_6#RUK@+dEA=6S(=DW)J)cQ(E\>C?fcYN)
48,/>9Q;e;7b5CA.PbAPD6TQBFG=I3R64g>=7->/P_:XgI=XE+>ZYF8UVf(6U_5-
2=G1F0W:YJT-@\ZZ4?+>aD)]([bPe:dN/CJ>aE[U^#=a<1P-W(N>UCc-A>?P+4eV
VbDd6-#a=BO(^JTWaQ^>PQ/KYTOB):VL?;P^H=F/7e4OWa7(L0J01J<ZNeO):X:G
HL,5T1W5>>-gF/Z#6INcG2QRSEDOXBN3-?H:F<GE_cO5)R#7(]4@-d6Z\Z]0^(YX
B=g@Y0][b]P_E#QfLE(_3(BK>94&0AE7)aX=9X.[KAEILX#9#&;/)RFSN<75)?HC
f[;7H=O7VI)FgaQ7A:[6cQDP)TIagZa81?MUbO^P+;6=1W=P9YG39;gF/QAD=-V7
ZB45X3@R(XC/G=&U<^^=B(^L,Qd,O80U<bZ6-E8#B@AU6TDU2_90Z(QU)]=@=Rd4
7+F>cMO+[aeN-c>U(22_?408@J=Ra(3V[-LWPdc50J;KRT/.#=B3Z1>00ZZFdeFY
U;B>KIW0S]eKCg[DLbCc3^-CLgX>I]@Jd]>+C.RJ69/3<[U:cg_V[W1Z#XQ690dG
De+32AVVL[H_f,d[JQNOd^c0deK_)TTHP[1ceEU?&R]XQBBeXGJ\9GY,J-eVVf.&
L>O9@XU=PXWZ.g@:OUJ-9ABRM;Y;IR7)C[P,/F4SO^/G#ZJC#_/0)b2FI]@QT(UK
g)B;RL,70R;Qa7#D,?e3Z7>&3S+9_.Af#GJL_\-BN>@X<]9<d0J_@8NPPYJHG+J+
VNd</3:3dU/&-POTI-C+P/;1G6L=+gaRG_CU4:]VgIY#/8<0RV6U2e[L]^(2-ER_
L6Q-3Z?MT;/^Q^TJB^Ra+\V\SF?+)^6VFaE5KdUH.ICA21cK(6\?f2.0@Q1JC\eV
^_+&-W<=).>I;aJa7MYQ.JBf=#P7V9e7^K+GgK70G@&Cf&+;^8=NCOZCYbYGe:6e
D(>0<V?Y][W^^9AH22AS&e:<WN-F[33(a:9O#)@N_7-[@UeeV,E?W-.YJK3-W-TH
<4T>NS,G49T8;F.fR+eFPH0=cLSfLT,]+>VBP5:W+e:gfBgZeAY1G6P\3E(a,EY:
58:?f&R)?<;@@U>TDIg8:Q;LTNQPYI.#[S&D@N0g8698=AbZ@^g@JCQK=I2VV_/3
&=O\;(EZb17S.&cN9#NE+HfaA5[0MJCJ8X#PSKCVP5]d#;,1dW^4IEaUb[_,]<N/
K3QK[gDZ(N?FW>e),V=VGVI(CD>Z2&\D2#._>Zf3_e#.C:Vg)I#(HA=X3XM(N@0>
)ZIT@1^RIL:4+QgODNZ4CUMT@9#gJF/+SXKVb>MA\+e/YEG>1760a#D/X&E2PTb9
7SV&c]7)\AfKc^??D[;dAL]&P]@)>#H->2,75eA#QEY8RL90A;/,G7=[P#KDe/Q:
BBgKQ#/?C&,:SA>#,JO^Q@O;JB+?bd\U#Kf22M&BW+B07U4f6DC]P/(:g<NI-^[W
AgGY(,\J8J^XS<#=cF6MET7ROQa40NHB=ER;:EGY1H\e;;UcX)B,SF3L#M]+E@@J
WY=f99X?]I=9HRadA4>.H=2=K)8f;^JZ?13c()JgD/WY:E=7/YU=f^<,1_?cDd7H
L]P2Z0)Y-+?Vf1W[[STQ&+:NG)6,/5bbgdM<V6.](H7T8fYIc_g;1d/[Lb3T7?-9
RfGEQ[#^J5<M2Id1Ad+\Y8MKe-#8[]:/[Rc>fT#QF3a+//9D<A_DJ^(G\7KdE+GV
2-YN#e?AH4JS--I&48MHD9]HX,LcO@VdS&)@3AS/.cH-[I>Be#+B?;2&9aY],g3a
X9eg<L.5PeUE:HdW-UE=#)D<.P]]HTIU[:J0X)6b^g.C0T8e@a9.5CR>KZ53IYFb
]IceI3d(&35f47BB;_<]bffJS(>P)ceOZd4R7<GVUX#4Z1YB=>>Y)3JL-17B4Q4F
5dK>+Z0W)(?=E)eHVE2Q);gb9aUe:DfSODeVW5e?:[F]-&?fBgX^=?/3:Z>8(1^F
<S?38b^NH&N,9_=[[C)5YaQUZVI@J7A.:E0CcM1d9@b-)Za+=#RAR-W?H7P7>=&>
=5a^>e-XU[Y[304/ZIKO2P7f>7RO7g<=c[#?Sa:5@ZT_-P@JU@38,)9TAFfZQ-Y>
>SedK3;MWa1e.UC^I6IGQ9.;dM\4R(fbcHQMf),Y,V+d:/[GDdOQ>RIR8J-M:+4d
&eLF4HEPPAI559G)M7<LC5TXJbQ<EcUS(A8/abX4])=c+@b4I-U&PUXI-UNEO&+]
;5<;KH)dS51_QRcSeb,g3GC]:F6I>=2,JFQZFN,#/7O(.cD?&_5[==]9-LUeHKOB
8=A7cbb90YO7_DNDFR;Z<N>Q-HcOe[_Q@Y_XY6(GP:N4G?J5&4XDMM[a7.[+WJ3M
CgE\c\U>OEePCdN4HdH(O/L>=OYH1.Y\1BePFa8=ULb&FES/U_NS:K9g>b6NSgeb
AAEC4/LLODDOA7WEW3EWG_X+GYZYaKONcC3.<Wc26cWGD)[6T@W9b7.M5QdJL+L@
bFHSCK#b1UTDY++PB(8__H[I-#@KJ=_+6Y-,_8bX4NF&;O.A^U1W3:O9f^aQdLTM
+&62^(4>>CKg[5AcDJ42;X7<=F6M\1FCIYTUb534cZBEES\[BbeOX.0+^#>6EDF;
3/0V9<4]4g,d<]D?=R=Z>B1+YbS(]M=552P5e2>RXY<e.+GM,.NYMaUH7P_c?f5U
7]\OH(K_\<=Db5cO0DN=g[H[@Eda9.,[\R^\0C8P9R+LUPSY2\S7V/7^7e?fW,.f
@TS#GZG?/G\N6BP7MWXG?5R95WVDYL1e0&NY?8>3dY8P(W?L6SHc:CVT-G9L:V[A
:96[MJ4]Ra5;[.HP;^4XU4@/@JF\#HSKCC+3Y/:@\^NI5T@]6bdZF/.gRZb5RZ(E
3CA><E6XB<S@.[F=Pcfg]CQ-WUWFIZB;(fJWbg\\.5SX&JaSV9K.2,G<M:Z@FFKT
f0>QWV+LeR)?,5OcZ8P_)B,SA+Oa\A9(MKI67B\_0YDI6ZS:P:-+DAWMS7;(S3d1
a<]^S);MXM?ZcGWHY<8aJO9;YTVRdgB;?NN.L3P/E>e96CB4P^P/W^W3GZQFa&b5
bE#3NGM0)1181bb@:AU>8QUUOK;?\A@ZMbbLK<NB4\:a=23UNH3K^#E.gUF=DGUC
cC\c>OQ124Aba.8+_ROd&^/]^^8&9[3g,=a<E&^QY8W(d^)1UAKa,3/aQfRJg7;,
X/(:dbU@V7dITBK,P7d^cRW,f;2B=Z7H]VJ=P@g56e,E]NWI8ES[#U[ESB/U2]RN
3dAJ7OR.LHg@BJ7Ced(ZZ=:>.41fIXZA9)[\g>&KeCIO;Df9N0EVA+F[g(VO0bH?
f_[+G5<:4AT@#0EJ1]T_&B3>9(YfG.B?MPeHG[?;04_(_@-K4W7IHG5_6F@eF5>(
6Tb:H.6FS=JdcICY](#P\\I9BMEf=[fX+,GRM)-MG)-dT\BL?GVFUb2<5](>b@39
g8aAgeG=2-#0OX.M2^6DHORd)08c_cY5S?V:\d;QSOU94BK.bH\NVdPBbSS))6<E
3S(G^ULU9gN74OaaYJGMF<0Oc^>\,2R_CEdKWV\Z3H)d=8SU>1_E1/7/@e&4)V]Y
#,PQ>3Dc1\aDOda3eYUL.(V+e8AJ9(W1KTGX]E35?f;dJ#<-PFJ3S70e6T4Z.N5+
PX?6Q;,g3]N6&.JX^Q,H.(020BETC9VO/.G?VP>Wfa?G5bJB\^af@TKa[RHEP1ZU
VJeEDI_@a5&OXZYfgXbKa+WXedcXJ;]T4#b@/Y^+PfVU>c[ZKT2N^Q3eg<\4ceQN
[eT=E+T3?LbH__+#RXNP;B942):W0KC;]ELcdW:-Qg3a:\+47WM5,U[,C06Z&L2;
V\:FJM4/9_UB>dg[@XG\gFKZ77dHcc<=@3fB3+9SKa8<ZgA\QRa]GZ</M1@eO76=
0:#fO<^-=S8S]eB-E86^5DXJaDEa=#^XGf9T#E7;Z9B>dgJ\gQD6\UUDQ4(+6>;M
OV^-fZeNHHI],B;CJS#A)X9Q&+@,84/-#R)4Q>>gV]&e;MI&7-#\VO:DDMINcLR@
BU#]f(3-VH8-^9@TA[PAM89&^#UaOBRQSC6LP5cH?R;&04OQO6ND<6;K(V(=^3dJ
d8CI37:aNU)cdZ@bAC.ABY@b)U#IY()bf3K.8GT2S@QA;C6SG=)_(=K3Mb3_==eT
U26BRLM<[2JV=B5gM=bX_deNUKL&,a[0fFBT[A2/Ia5+DL7FdOW4Z28aRUCI#32V
N#e87.IY-[,>M7fHaUNV29EW-EKAH:7S898/[;F07a2GbF-EMFDD/\7O>#B<?ebA
<YQN-)JZ9e[HX[LR2c0A:5\[MeTTJ75Y-78^2aJGDa2G>=QB0a:P2fAGWW<76^WA
6L;[83,7FZaM_^.#K8M@N)0[H0=K8_H(N]GE<F9D\-8f)3WYRWO]/a+bD9&WJ^EO
9Y#B(<2_ABI>BM[PP-LbTbaaLEX(C98?ES&F\BKD58G8V;gZ8<a9O2SaR2(?#;XP
9PI=H<X-fPY3#03<\gP+R[,8_e5Ac4C=.,?JV]g[Ie);=EIL\A4fICX)<)5b97FR
TEAP8VFG.-FaD^_g53+SgU#VL;5YNdS1/D>=bKEGM]PHLcQ(aKYAVTdZ)-Z:FW.b
ZV+P2XU0O[HE^[KH/\?Z/]dMPb]1<G9>1X#(D5b#1CXEUc=G,[J&I,.,AC_,ELOL
e=B9LAU=Od5LaK)CV)4N8AS=Fa0>>8\@AfVJFUbB./_g4#,YcSeG_SJ,(:dKZ:D6
;Y(E92W8egC03RV?HT4.UbJN-:NIE2@@QD(3SFLW[.+M21/@b7B[I3U8-X?L5OC#
DZ@gQ:9J5FY&\R]EN@bRD,?b3bYEU650T4[?0eLUUKG=V3++5Q>T,O]PaSR_RT)c
QL<L_L>6Y-GHX[HM.CJ_RU/P@O;+C;cY@S,5QI),SfIAW^T8aFLPb++7MB:PIL(.
ACgW])3Af85\V^@^aX:/^Zb_M3K>ZVX4gQ;[eOH>][T4K<-[CI&KB59MT+F:<c8<
3ae#GK>a&&L_HZd4[R^eV<CE,2d+&N]5R#(QQJ1,S[ZS/WZ)82Ac(7d(NQZU>O;H
K@.SL8[E[BXg@L\b0O0\E-6g[8;MGJdBF2=<.,5-V09G10[<?Z>3\-H6]>CA[H[/
^X+3IHPRLK3R0(G)Y#eXZA&4gBP69+a@,J&XXN<\29)E/@I_T\B>8=a;;0U5Q8BQ
QCVDD2<Yb:F7QcEGZ:C@/@3?L?\;#/7KO-d?a:I+6RdfaZO+T#0)05_f6XZ[_\GS
cM<)gSHH3_g++U@=[bdZ3SXPAVU11H;A96/f.Yf?C3LFB?+<+fgf<HgS#9[fE[U&
gZS)IJO/0[/?>CcCI=]17X&IF+0U(TC@&EIG)R,=PSVB2TR(>Z5Fe)cHW70Y9>(D
(#aP/e9O?_2I_YS#dRS)T^9^:NQ2W=TJbA6EY+@9&:[E[B>NBV-.?fbJeUf5GGQ@
9M=A1b\>ZC,JHU>U;XJc=H&[Y;bIWH56/[@I#fCW-Sd6g]IJ3Q8S<J.?TT.\C#WL
M_KTD@Jc;)X4DXHe9FB0a#>WO1TVd)fV&C3:2,9eAOK8O>1MM]\bNE1Z2gTJMM]J
5_S8C?/]LG<MXG+=E_H.#S774K@_P2:dHCZ]e.OF^+-;:)=?^1D>5ZVT453B/3Cd
OF6+&b-Nc[ES53eeE@/:]J[J#BX)[ec;@-WG]-B]2L>(=J[:U;M\+Qc9cYfD_@9W
B\]XIULSdZCc:cCA)Xe-;,_ELO):KYL=;V16M5@C\WaZ8SP^fP-WdWJZ(2PWN1V7
,O9OL7Xa&O5_TcJ?;XLCNY88D8&2=K6XY.>)D+:&?8,]5bS4L1>HHV3J:BG5MQFQ
dAfBJ3Q1fI0YQa^W/]6H<0&82I_-,=J78E-^HF:aVX&]S.G,GOM]=L^H=GFZ38PW
2^Z3(LUWB_LQ1#?cSf#.A#,c(W^N\>/Z5B]5d&>?K>8YYK]deXOMM8dABY]SL\5d
YGNKTU?NU#+I@e)TIXENb2V6F<Y37)KF(#V&>WaR,RR?7(?I\d5Cg&.=57-b+eg1
GH>+784cVIM]:KM>:)bCX#D^UB0[6U0HC8C@fY5ffS\gUFGP#X>-^1<XN/ZP5YU6
Mad<IONNB.fX1J,V#?V=UT-;<T@D3=,;bDXGO2MQD=XZ2TXTCWAcDE,T(,[DCT6<
,Z=gF+d_aOC;O-dI(c##R(_7+eM6B^D^g@=(EAXJ^1KbD+)/aS?T0,7MN=NYC-Gd
O&>6/:)/L0e\;0Na_S-DNE#R(=RLN=F)^E>5OR+/ac+[9ZcWNN1+8Re<WgMFFR,c
H4<+0+P9TA+@@.c3e4&ORU?1L>.5eSDE(e;S8Q,(I^)]7XBHI?7AaU<9AS(&V8OM
/3(N5E9^-LOM[I_4A&P#4=03[>P/0N(Sd3#/fQXA]D>.X39SaN3fWP?/29ZM2Q]#
/PW2)GTTHHY1];RZY&#\Q6#Y_g]Z9Y0<dPC37a;0gf8]6\4S=>1:FMSY7?9ae4Ef
=/[L,BOg1CRO0Zb4#.V?5d65C0<FUM-CW\?QE8_1KU2g7?T8P^,>+O2Jb,c;RQ9U
A]G-bIP32XYceRF71?<BGS7f/&#KeC-QWbd]<1(P@4HcPS>6G]][>3\6fOO:BQWC
d)Red1d9S=_KO)W]@V)15IO-,3f3M1[KP>)GII,eOd=AMOXTKX3AM5Ff5:)g>cC\
Id3f]SN\TC1Q[3R\4)>=.FQ_69a[.B,:P?1_Z](#4f/UR/FW)XL]Wd;4g0>]bCDa
I81<,0YX^e>O_d>)VJ9.=FXJF\K[)OfdU,Y;c>Y,Jd8G_&]fH?F]A7@M/d;0:GX9
WZ?K0-)\aO.SKL:?[N/,a]R#cUQSSV&Qb515#2FR/eDZSM?);f5bQ6]H/_T_6O3W
:2X9YGcDTW>TR78IF)NaG.:EA+G>T;fG^C70a,(1E+VVT@TKJ-8M@2Yg?8-T.CC[
SZ6\aaJ_H,90.8AB4(ffVf#gO1[BZ3MU<Bce4==;E+EEI-:->Yc15\MN@(H@50)[
\aO]O3,#HEZ5e)KaUfK?\NbZ>,b(Y[R7a+@e5O^2K<&1::R#^TR=Hb.A1;JG=Kb@
aW9;9K8e[cOG=Y4:>6<V5R=YCcH8G@Hea.?1/R6O8:]7TCON]gB::OHB.\c^MU,H
^8.dSFADUg0bFI;BW>26G@?65(7J-6eAF/>6X1<@K[G@Q=C(-=9X^BZ2FC^47Qg-
Zf2(<85CW3DU.[+STFUaZCV\MOVPZT+I?)eHeHgN2-O\JP^9K>DORWa36>)fD]^U
?8Jd#If[geE\BE.UZW3/cI.FL.9,Ab0b&?NJYVJBV8T;0X3U-Hbf5.9P@baL+)..
8DQ(?AFC.\]A05acHZD-VL^MVOg6]06,Vee8KKNc-ee@M9(F9eYCFMb5@C4gZdAX
-XZ^(b4<4MAVYZ]GaO5<BX(D-B#T2Y#XHPN#>5[UDGdMdM?J6[#OCcN683e;f-\Y
2L=UV=T162@g49)8]6JA#:>GP\Ug;O8K:b]Q268;#=-7Q/DNFBH>Kf:.QPSc0CC;
8c^1^K3TV^IfB>1fW(ONX<-aS&)WO=RaSHC:L>1D7]J+9CHb7#NJ_IFRZS?e]\O[
:SIB3c&>+VZb@fB[5KQMc@7R)(dRYHBM9H3,S7\08@6H<;A?aCC<,3&S&ZTeM?B4
W..:91(N^]I6[&[^)<CZ,^0\HdZE1K>c>:U2[KT\BTCeW/TaH_UeK+Q&29dP_6QD
-&V[&_]2gJeL3R(8?C1ZK_RFR,B(2)\M#2&\;.B0H0+,[BT8c+cDYVfLRE3-@KR<
/9)_BbMT7P;9A=A7CMD\)1.T6I((.P2F4UDB&Hb^3Z&-2ab:O9Q(2CeD^>+/UEX;
cX).eaM@5VBS[6X3&=8#[F)gR#b&2@MGE&EZZM4c2&<LH.Nba?YBXAaf=9V5+5W3
gGANCD&cD(b.Z\gHJ0@I+e9KEJ_<1&aS\[58?f^dVTa(b85LbIMb.8)L1P#7;d-e
KF0F\YbYID[)\IW]TUaE1TQCRQ;42aEIcB8YVIRC@d/;ALF84e[Nb=1]3c\W0GE1
D1H/.J.XgSR.)^gS.fO;-CWY;7:IcHD+E1bBVV4I.HKZafM>be8OL-FXA#T0=Ua6
USOg(,5&>EX_N.>I_R5C6V[;K(?,<,VG<.83Fg-RG2D6EA?L^^N?g(#b3-))=;>b
f-Ub\&^1,11(T2\]=4d<Z+;\CU5]^EXeAUWSC_dPN1HM_?#8fBeg4B#=L_2MQfI9
1&ENJ#b7A?[SBP#IHW?d.2@B+b_<?E0U3N/9FdO0<VO3AJ;&;4Jg&_4901/T386H
&H,P&N^H)D,33HN8H,TMaRfP9YKd?&7c?@4#c.Y7C>:C[aaO4=_XBN]\?Qa[)13X
-6A?,D;2.4^TTRV2KgVb^Z.c)6;U&&1.)4-39Z_?NOPgfeLLdbL;XfC+T<.[FC<A
,4e43GD((_RDJIKde\Yd/5[XEJ19QU#?g(gR+T.6OSS+Z_5,f(O3KQU2GR6f23d\
W//IA=PN7))GTHE)]e+\dAY1+H9CQ5cZ>\P)TA^)>:38Pga4TXYc00.JIP/NcV1&
^(,L90c00Y:I;WR8c4KPUX6CeV(IQbZ=>582;;)<MT;6&I=?EV>Md:Y]AFCQG9M(
1MaDX746^2e,;#J;CYBbga><MG9<-gP+>QSC#L]\8I9CO.c75Hf=SPV5b2]5WN>.
W8II0/C?)2GP_Q0DSZ\F67)4gJW=R?LdZ[abOX,]FZ75-(?<3C20=6_VPH,M_2Ub
V#@Z4&We@N\=P>9Q/DS##)e5a4FTX5c_c&H<UaCL-.2PX1f5TP08AZa9O<aV/EF;
AB+O(;&>cCE-2@4.1C7@Ic^Z(cM[Uc37\:@.C3@(7DI.JIE)\6b-/UW[DCFM0D8W
ab[b\XcJ@?;V_fe.9EHfK/A2bI5#(;HRNZ,]8SOeTC1^G^b2K2HP=LO+P(JI+^_M
99[NU&a]Q5e<7B+8W43W;8W<^9cLe(-[M&UU^G[5d[-RBME@N^fM?D:ETa)ZP_VD
4YK]c9M6KG<8.@UM^LSb95;E-BM:OIY,g)37fa420LAP8DM2#I>C4L;0A.\G0HIS
[S6C]c\LdI;;)L3A?#Ke=M1#<@CPO-L:fG42=>&^#Mf&N;P01:J,+fD)PeW[O]1,
E0RZ,AZObGCH=3VX[PUaT\](D&-/XdFT(E\S/D7.4V[LRT_S/AHCR]_AP_?d1Sef
fGD5d/.ZJ28,AZL5M:dNC8Q:CN6>J]d)>eK#5-4&)@=G_g]@Ye_]8BX@<e&eI(_c
?(ABMK(cC/E\+VP^&1dHKOXMY5[R-S\XJ:?\bC08<63IcALK<>:cN9XE^Ic9.7M\
abCH.aaWWL448;&FNG_Zb=;P97K]FKf\_N]PO)f/OaZc#:\460eDKH&#^#8]4LTU
7O@;bO,J?SVV^;9V\YS5,=&GYL_,)GKc7e^^.:NI5GL?d>g)b/V#G->U<bYN^3_B
)+RY?H-WPA+]3?b?5K&]_aSDOZeUZ0+DBYPAC+\)?]]<^e2<#_X?3\T/^2(@bQ?(
(?RMM4,#YM^NGFU#UO(5\cC@JSfNHU#89Rgd8OH3SQ.O5D4O^D\(eH5]0M-e829e
2R[d1@;QVOVPS84JKRP/?^K^B6WSVG+4-bK,?N^]U^&a-QZ5aAUGc?4J?WR27eWf
)@4Wd;Z898Y/fDD0]e6R.JBOa4N@Yf2egOaSI-+c;#<&VM2-;XNV\/=b\WR9+PS7
]NDW1,JJ:[^7adMaQZT)JE;@,+_4K\Q8)K9;)M_Wb=4<_12c82JWEaf/EK8Hga6K
/=_>))88PLQU\XdG,^/bcST:Pb.2eY96CK2R#5/H-O1c3?X[=-V/:<]/eH&WJJcW
gFG<FU@SYPWb:FET_9H2dRG]:@63,:Q(.Qe((49DSWDQgK.Jg-F3b85K?(HQR)a>
#0KK5<KfA)<Z@#P119MD]E+:,&(X@N[SX0X?F\S\]fAI.R_8HXNdN4Gbb2#aSW>&
ZH7_/L\I+<fgb4a+&F/00S)\IXRZ+_\]a6V0ZJ)J&O_97(VBI^c+5787^)EQ=9LX
8X:>,28><,\gVa[^[+>;U,M]b_(5Z662+_B4c6-:@45(OW;?>.P([O&I9@QE0#Q2
KD&7/dK0_+5#SB)^F;HRMb8P9_]+P-.:+dXBU)c8^5OQTJ]Xc=>R]-=#NdIef0N-
\.ZbEcEAG#WW6:\4NJ8;6P8MUM9M]5IH,C;=cRX3C_+TNdf_>]\?5>0P^W8Q_^Fd
X/UTYOF(E?GEJ(-(MAXND2=IJ3<-8E@(gB4]\X:<,)bcK^R>C(@gX[e8]_T>SZCB
-H)+<5Yg+B,^JFR8Le9JYK7+^7RH4>;XIL]3)&3X(19/>6UT5a)Y>QdFR>,6JFRH
[FP;PU<fPI+2WPU+DG0#_M;1N@\/cg[HZ)gR/X).f9N9S5C0Ad:+d30Z/ePL)ZPC
V_]7ANaF+3R6e3QVN;6S\>)-H8J,5)([<E[OS@]SV+O0eO3DI(&eHaX.eUCc<@K/
?;7F=G(=QL6C/E#Z4FF?Q^1JL;6,Y7+K9,-I]-fV,cCTNE<F8OY&d6b0S[G=dJ4b
MbW>@fbE4<HQ(d&<D_cDGYCF0Ad@9cb6S^2TW]2]TF;[P];_KSMaS.R.V,FPX\^0
:?0/fbGf&-.O;B+e+YH^-XCB.77P.M(81.4faE<MS<5ZD-+3c2TEbgSK+>RG<W6X
S7^A.(2/RC(X@.9PEaR+S0QD4XYH=0P:P4EXVe:7[Y3G.(H+bW:.H=.e.ZUYbTKI
&/OQT#.&&>L)W2D8,B,71:\-BOa6?S/_^B9H)E0d-I8dUP^=Q@H;a)[_7gga5.fD
.g:6Ubc8\9gN_NDG2?6X#(#FWcSc_WAF_I<M=Q2);P.XIIEM;Rg#[:\=^MaM>7)S
>=T1b[Z\0ge=\UbabBdYA5(b@cHOZ.,b7DW)A0O5Q0@=?41W>=c@(OBKHe/7EcKD
GOgVPg08C]<V8IG8F0J?#NQLUORO4ZA[8dO;EN;=1:-@#0>UZ4<LUQcCBU]R1dBY
C/=>T(+#OgB]RQ#]/dLHM4S3^f?a1^44XC#GM6M2NRJg70Y?=LM)-O+0-4gSJ3_D
_W<2?7J@gEC+AVTMAb)d<AQa-#Y6&Y0:[16HP7B<^J/ZbM[11aNLN=]S2ae2YLO>
DgUbGQH3HXTM]K#)R7H53SZ?2A+Z7^-?(UPd3a><0ZUV6_WDC0K4bgcf1S<@&<WV
.T3V6\QG9MGL3=K5XGDI9Tc[3X-ZMfCQGOPW+BVgc&WPQGe]0WdF).QZeBfR0F@R
0)X?I[FYFOW[T.O(/cV9@V8LLO\bXUb0FCc<.]YbPZBE+4>gSG6c1[(@e2@eVP.-
.VYRA,E?:#;\5@g310SN>d]Cbd;\7RLGc&Qec;&d_aNXE:6Y#4a&O?048ReE\0,>
=O1XHF&0<gPY&e:8F3d?Mad4IYJOP\(->X_\W+HRYCdLbgf=E(N]EbDM9dNJ:<R,
U1<)W88Jd(MI;VL);Q9C+I:I\@1?V#22WTg,gP<1._)EA)+Xg<3NH[Yg\-PR6eWf
NdA\S^?V&\e3RU]C5S(S&R(\.<WgT+S=b^JYTL;UK@TfIZ-Z_@5gKP]TCZ2(3I9O
>F(dDK62=Z]:[V9,XZ@1V0W^B[_f:-^0:QN?L]?PUMTW+<:eB4PO)H1K-0?ZY^Ef
+L2AZ,&be(.,#+7(-BPffMTLBJNWe:#LFfE-2DJP+G4U__X;)#M1L.X5V.TU\(Id
1#VSH>W..T;K/[aRJB69Lc,KC[5?T3)#DbJE^E?WF=NS=c32XXXK#J<Q(KOF+DO?
LN,K>UJVa#;#&N>f#C.+C0?9XfKe@gWPc,_g[1##44O83CW3E&McS1]B7VB6,gTF
Q]#ARLbUcI&/^;e20[L/>,Bd1Q09\DfHO<d&\IQ3:99&7XYT53[SaN<>]MEg=@V^
G_U^]VaZ)K;?Qd:bLW;RS8;;+]&KE.XPBHb8eFc1]&U+7c7-\/McKVP.?Xa(R3Y7
UEX#^X=R1U0WH<NO1ZR?L,+J8;&.NJI5YOBUJQ8Ef;8@XI7[?6JaYDGAGJKQM6d7
D()Nd+aEMgWS^cVcb352c337S(<+XIaIe;O47CHf57PO>WTBE++BI.@98&-V9@_<
=&c_FRPAMQ-#)ed>O<<THGXXJZU3K\7VfWN#d;c?b=-GO,-M7^R^7+@cAe?DGa,^
Y_AH7F5URO@dS._N?Y>7b<#@g/&f<DPM5F.XNe6Z+&-dIIEBO@]#Y1==[R49M.cR
AMIYY7(SK,43,05/CQ35]Pd+YK>P,6AY@Df:L/S,aS84AHEHF9fb2aJ8ScF2L2>c
?;LC<NZcX3W+J(8O88RUG9gG]0Ha=LF_PF2W&RRF:C94<1aaN=dAQZVRb_9PEOG^
R>XN?dI@,a\^PF&SS/IG6dD4)T[,(ZN9?.H6gc?_eY?:GZA[.9KSBd\\R5/6J:c)
&MdQ9<__aIKHae>NB;SbF4f5dJ;=X\DfRP+1&/#eF_MA4@_^8CGPQF^LLQ1(FFR/
.[WGW#>)CL02a3e95F/9L>72::AdE)QVZ);Xa[DJMM5LH+#f;EXC^__eE;#@NPYg
Pg-C5)H/W:Q1YR@DOWgBO.U>1W,5&H&D<T/dcGf[@3A=TcP?2)1#^^f4M8DTQFHe
\ZZKc&?11#AS?ObR/L[85[NSabU+HIVD-(.[2b_Q2J(&_)B@L[9>YUc?.1-DJ/I#
gPcK><_\SV<f<^Cc5bH3>ZT88;ef=UF^=8#90>C_O+PIb7C?MMS<L\D+.>f13]T:
VKMQ]?_LF]LO)_Zdfd>f:5.6IReX,DQYaRC=4dHYe<NE0^0FE7/)cRbfVLCEIESU
WK^>Q/YYIS;P&C_&:-[2_QLg?=)@CIce?Z.^11[R@\^/;FV[d2S4Q?NUR(:F66?I
M@HAZ[bUE^XCOT<+=X6_NNc;P_AZPQY.cZJ-[[83W^3c]4,7.ET^UUe-JJ#[_E7f
IJJ5UT,GUQV#aUS.01VR=;WP<gV,D2+M-3?32g=VT,\Q\9g5&gH_f?0KKQMe-A=-
bF\.HUa]I394DHWR;:,Y[>EO:\e(H-B#M9Md_XV<>EOfO5_5[3fY<,b:(Q4cAV]V
2:D@24NA]FP2VRJ4^^8B76@RD_)D.6Q\]LBT2H&DSD[&JX5<)S(dGV05KB<CRSCE
.4<[N_eK@,:D5<1AE,J\:8]^\X>\?;6.YY:B+V(1BQBY3_T[&]GL4&HP/OeB:MN1
VDHYK1YYg=G,H+4b\?fFZY4ZWXPV2Gdb_b/8(cU#;K,+\&fdMcZP&cBX@F.?O.>B
^UfIH.C&@+])c.TSOA]F2H^73R6\ROeJ^4[G,J#2K3Adg.8WEeHJ+gb(<P#a(QDH
F+_-<?K.-d6dD.AVEa+-dA]W2V87a0]@]-ND[A/1789(2Z1=YM4_KOW@/N_>LSO;
/MHJ([LWf?RaY^8.(SH+2NaK+W>.gL(+S&KC/>I\3(;Jce(H.0/;6b/?>31Fc2f>
,@7TT3G4dZ.WOSJ]U/T/]aG5S\bA95V?1N3[BRSb/dPe7-KQdQ5/@\DMBe877H]d
1<(#P6X6Ng>310^?.Ub+44aQgD&^<e8;:L]\L#-;DC1f65/db:HH[f]SWT[/f+_J
([_V]14e,@Uf[3YPF<MVdW5NcXQ6=L;6)P,g4FaD9dM67HC,3+d=Q3Ng^WXUW4U\
/)d?36&YK7#LAe>a#WCP(_A&77R@NIZF;??T(I<O17<KBTD4.#7=A_<cg#N.IYX\
/_.C2J?e-[CWP+-#]F=(Ud/8+/bcfXO\db[C_N]9(2V]42?=bd,G1V8M=@dF7Xc_
4.YJ0M,d/I/49d\:2ZQQ]0bXYIE#:\g06BK-QeSL\fJVBf-/6E:Q9(GA2O#ZRbJK
N\[<]2O#-Xf[TK;3CR7L32,(3.PcS26E=:.QS_6I^O?Eg=JQSJ//,c?(fD2CFSRO
KfR/TSb6S+<1b2[Z<\EX>4=f2O9[Sc0<cOB.OaP?TBT?+K3b0J:OEA^:P(CKM\=4
?\K1MR=3(cJW;AL?VaQ9/+&U_&=,P/X/8?(]=abRT&7LS=+eGgf8YJOd>\.9[20E
^)_#JdeFg^4BMJFT@E0f+//,,2QE/IP3Sb8cUIGJW]XTc4,(AR\^9.dVUI^U6H]I
O+DaL05?-6H+&]/ZN(EC3MJdAU^Q\aF&d:e#THUC()-_PNdIK+,3H58B,57a@gA+
:(?KV;5]0/;\.0^TS&ef.ACV#L4Xd9aM2G+16,.KBaC?CE[-aBfQa3a#JWH)&D([
B<VO<?@\SX5^SMdMgZFB8G/#DQ)fO8NU-(LDLY2@W:3C&UN6-K3]Qd;FO1Y6JLbY
6+=7gIVYB>FeI02P3W5F5ZAYcFb76?I8PHK]6]d8X7g+JRFN#,)dW6OVJC2NaT?V
BWa_NQQ=0@548cI+M_2T64,e.:>I0TfgI:eBK4O\cdF]e8>-.AGK&=Q:_3WF<f0O
EW#e+4]===\]aGQ.]KSD9P+9(Z@Vc@+Ca:#GF]QNU>f^3-LI]9;2FAY60+/83PFf
,E>O+;+D@b,TLPHC:7TLg?K<)e2X[2P?-d+HMa(D)#ZJ(d?J_g74:d43D#K(D=GF
EYfYYNOf2HeQ+5Q#53P#G7F7CD)NH)Kff?(Rf,/Z\Fe8+QT1A3VQG6&/+VDP42JW
N>g49Aa/ZT7EeC5RVH\?H\+.JDA.TT-VWf2^fKc@/(,.)57fGAQW+cMX,dV7JEO1
eHLK@WSP@W(9T)9->N[OX4]S9?[/<AP0Q#.;#MBbC+^HJWP;-H8Tg(?:&8:K8N-d
2ZD--\EJ0;Y,K\-2EgS,@CU2&)&XE0_1FYXSc^@7E@R6?0aD5^GM,>4)8&YL^X-:
7(D4C(Sag1H#V+J@:2@NPb#UHONFI-DI4BGZ-[d,0J?:7f1?J&:-?31TG&cK0@6C
&7QD\@EO1.^_WP5NcM0PK_<;.MBZ&[FS_UMd?-.R:5:@.)<O@(=8XGUEa1<V7>.0
3V7cBZ02bC@dVIC:<QJ@-8/4\[&K(74VI?H4),_aH,SV[:6H,<&3UY1[1=3Hb(-T
b#XX5+>/S()?UT_VeI9Z2:5W[.E_.T&E>4)eG14;96G/8ZS,V&G8?G3GBDHK;(_Y
VI;-YfV^Rd/H0.LO7JL;U40;PPPOBNQ8CRL&,<KHTcLZ4JX@02bffS(<>)D_DfM0
M1@N?ABfY4e#W8[].YY+Q:1>EPL(]bG8UDV&CY.][BMb2N[<L37;(6E/AQZN?;2)
)(\/;+>Z5XHE,+=PZ5GcIW^FeL4SVFQU&2,;d6+^cY0Bb=;P-=UV;HGZX)/^F=c)
WQ[V+1IJ>N2HJ3cUOQ</?YG=aB.0+.)?FCGC+a<A#-S@-.C=?]=a;K<+6^VT2BR[
d@_Y+U^KA<Z<07Uc3FD#SQa4HA^F(bZPZ0D@FeaHY(0^8:=>HX#4WJ8E+VT^g^BP
#VUR</,g);ERBfZ0I,635b6I:_2\7cdEL(9O/OB7Z<GI5G7P+((4CDC^LFcF0[)F
B,8>GDg4\aMS0NRIUI2L(RV_c97,Oe\V@./4cR&VUZ<eMD.TAOZU^[R;>7TUB]9X
0F_:f#_H/>OG<RWR-H5dHD5_f#\^VbEQ.&3)\1bUC5P8gQEKOLd)(,JaZ8,-0E[9
A8]R6(XL/cP=@TE1]+8>_-a&@QLJbRdLNO54#aQU(K3EZeUebZ/)D)<A_A:X3H8e
O-D_N2f751+B:Af1BT82fK5-IJ]bA^5>J/2I6#F9R>=?1_+8F9-Gc-CK/>SOX9FN
MSJ>#JZN59cE1J<PQ;PNa^IOO#RS,A];G^GX^Y7/.6gX#d_#^&f>ffG)8U<QXH>(
8E9A\LZTYK(?>dc<,9[@=HN,O@3:RRU:58O[N5^E^;[8H9=&HTf^QYII.:1OKQR,
>c<7XZ(Q[S2F<+O)D?Ba./b^Ef#9DE]SRc7^2H&F&2,O]-&2RB-N?dX;Z;^XJ>3-
=^dXPOT3cg<O:_MO5g,1C^>__K<S05gC/.bGGMb4]O:2P.>,XgEE#WNFN+e=@0TH
5J]+JT@Pe2g9C1+Lf;SL<3PM6CLBdL-B.Mef_.dDBR:^G6g&C=X&(Y<&]XH<669X
NL9g1c183NRCAL8W\@8Q5.MC5ME643eQ1K1.62&e:Z3bXbFCB(+TZ@([M+0<2L6S
G)P]I2_&UUG/:JH,X)I0GPJW1J@a8A48.BR#X_MT1I@f>&J:VggZ[/X&A)UdE,e)
0(Sg=b).3FW?P@NA&7->Y3NWfP:gcd_GRBLB>)P.I,BBG=28c7C4E&7(D\J,#TLT
C-LL]eUWME[>\Q/Q\Q:,8F;0e]Y1TI+TBD(.gJ.eJfS=ea>V_4<E(\PA5DY<G?NW
fD>7HCgI_P;bI0aQ([gMTI>KR;E>DR/<a\809=CC/?Ng&FaQH89c_2?PJU7Z@H5b
JJUd=gMZIQ<)I5W_ITf_=KCNV7H6<8094.6A3fG;2.8ECOG1KNAS.SC9fO/ZR<Y4
c5e:e#343[GU,4V:6E9_>Q=6542A30\JaeJ7^^4JO5?BR5A+^Q(XX[X6+M_B1+68
9&gTS-d08+;AdDcBU58Yd^agK@@TCT+)NVHC,C-Z2\P>&JP+WBc=CeV[e^<C:O2<
PMMO]4.L<I,<cAC]U02IOgV4R:#5.=_XR7CE05X3L/<.T&WMd^2S8)&\1/JG-O-_
&Q?^8.^\J)FSe&/)cJ#)82(#-J^gB-)f1AQ+8;90;MT>eE^RGW39?Q=d9WZ;\SG-
8HFgTU@OV4Ze:U]QK5T+aTYNZ^CWB/RW>5;5B]Y7]?8ae3&U9Pcd5(fWRb@;0,_g
Z:I()ZUdW@a80]0bDHT^SY1X,P)W54[)_:7N?0G&79YWcEUP-IP4-B>He\\aH//&
7V_7PZ?G;CM<W.5W\961.S&&+gL7.=f>c83PVGf_)3J?eZM.&cS8;>9?P:9BBc^F
N(bOBZc2KVDB5;VLbeeSC9N/&g,3fX^DF@+=?\J72)d_P29(S5S[L-(#O\:g+.[)
\VC+/337N#SaW7)V4UR=;(eU7C,&R7Hf+gg=U1)BUYd9/;Pg,_Y2)M^]F\8+^\7J
e7ZK<f-437W&>#LcN-7O9.2b\g,<<@)fd(cYbJQ3;F_)dK;dQ+,I</@N\<fXP+.c
AN8-QQOV]-G2MMF5/CV(4cF_H?R[+\1]d]HE7P\0NVW1MBQ3CbA6JgWY23Rd@G7b
;QXVD()R5TIF74W49Q\_/1U=\)dS&4bbYS50J:JbM[7#\Id9MT2N>A\L)O_E3Z7\
9?a&;H,:7QF]NT.6?e4[:_/1>HU-UHc&C5P8]R#PJ5.NX/(2Z4K2_0gb@J2LW\dP
d<#&SNZBXE\Y=<2&We;:_,7X9M2H(&Q<WBVc1&39I18^XP7))Y][D]eNE8L)W6d-
B_/MW4GHe2?2L&:Dc\NgHfC)aFN0:]fVW[6];N;#<&Pg=M0+\G18-;/2A/G=^G0=
)?C^N;34Y;P1)[R4e[c\f/[BH)cA)&(VZ33c8g951.)#V?NO37dgVI3?QLEMEM]]
76K>.N#Pg<=]\;#b<I+MN@F-#@+b]DIKPG7F?ZED0dETKRC\:+F3(R:>fd5@H:HE
5BD+cW6VK5)3[1cDSBZAUC:LS/fG;9(:@8.T5#:,(?>)/<4e)6+#4SIb6Qf\e5^G
6N-6B<>aP)\BBGbAQ1]Ag3<bW0#:aV2YPIZENgVE>1O.5BFaSDRHTA:&.=TN^^a9
5QW/P(S.cA75XJT:+9(+gW\PU5Y/Ce9dIE8YU]49._QbJBbVaf..)FbcP+()&]EQ
XG(_9A82g/X@^CREMWS9W3&A?8P+OE;d^S-1=_FC<6Tg.S8\?3A>-R@.;gTA(-X&
?0ERX\08K@TM1>.8E5J4]4I?N/W+11CN;W/)LVG^,//QNF@KCZ@([ZA=2)[@dK,T
,GQ1#3a3CP-\?&L4a\6VBBU=#3-0)5-0KV5+XF<QU&#B=/+EUe^F,cDN/8DDET4[
.[FN,K8BMW-KFPRV8gKGd[1a9NggSe+#(Db2cb8C^3dPX0T&c)YR2WZ,D&P:\V[g
/Q-HYcGCXd#1IXDLA/5T04RXL1M3BPMKOZE:=Z>^2\3e.fW#fN/I)WdQd<[UP282
-1G,8JC5Ff2SO##C:+0AGB^aHCOFWeWEGD\R8dSN]+(/dVb.c<c4>gB4HVK[O@SN
#[,-?U39gU\fLU=d.I&e@Hb;#>9:M4&-3H8)Q)E,2IeT^@6dS6Z:M?=&8/[4g]J9
VaYW6:;HTDJHBED1]#[P#6RK5.QA;.JK2PV<Eg0^N^\KLY+93_?\;;A@6@3b&&C[
N[GT92F;=DBRWY<[;SEG=V2g-K5RSF1<A^f-\M,LS.7DH>LJMa3BNSe)2.6\KLJG
9B/5):JgG+C-(11A1IOeQF:fOW^aL[[1BXc/4R<F63:D=Q@FU0O&)4=3_KZG>ZMg
dgTL2fL_&#SXGZ@)c&KZ40a@=X_6SE#I(\MJT/>)CKTSHHQeX9E0Q<AeVG5U(6E:
Wg-01&c78,D+/8DQO)973P4.YbZVEN@QReMcTMD[.<X^[,cKeT]11ge#)5T,031<
JL@<>g<4&+?O9A54/33=<[P:VMRc.5F0aE)@]F/ZU3d#KO8,]ADXaDHY^_(X74e8
Ta3@OKH4XK7Y]@K95XG;KCS=a]+03_NaQQ[YO+&OH/Ie2f+23B]GEUUa(]?]TA9a
R6TKY(YbKT9X(bdZYXGNO&DRg<(ZPVKbL[([S\9#H[Wg#<0V7UG>>RcAS6abbSM@
Fd+<&^gPU)cL.F>88FKOD+E048798@K6c<VAG:A2SL_SFK81[.-2Q)+0Y:,46;R;
-E,JRVR/RV@YFbUL6MSF2YC.7,T&VAHUI&T]6#ITA_BB@9Dg&P2]Gc>5g.)8-^<@
dbZ3AJ,H:514=[R-NBN+e)3JUgLH<R2Jc60?\DPbabG<./GL[&BcaA3(](?<X8KU
2eT&fDH.--5GaTE?/81_F+\9E,c1S1N-S:eE)F11d#QI)H[[0,1GKb/L0G7X,g3I
dTRT]5CTC4.1E/DI:QPeeNcfR-Z2KV&D(c7MH8#-X8O7I#/aSF3/[#NWNf;OD6f]
/dWAga,5YB9Z=T5]D;GUdg(&W=(RT<5-,))[+f?KT@aM/>8Ig@H:]d?eb/O\KHce
Kg.eYIJSLfJ[T22CM=):@cgE5)ac;=F)CR(gcY(V[BQZ3)3.E=OS;^CbfX=V\X+C
WUTG\)639UY]&BE1](72&6f#JKf7^C:<.DNf#VLEOUN/5DS8LK_L11EHM=Ac@d6;
K0Segb=_Dd.fUU08EgE1&HKP^40Q&]\&D+b6g5U/JT9ZI<=,79e4[P6bJR9BM6=#
X#bI+J[+H9&3Y_;/;@U[W]+)a;-D/V9d^6>R1.F5UD/^AFb&PI+[WXVc&fSV4SPF
PDa.c:80FA5/(W&LaR3)W2#;8XC;PV>S3aN26X@VCNU#aGKcTgI1[.>=V2Kd(N0c
G\ZPc,?\RggIW+0b9_\Q5gE+<[7ZGdecg;GG;g:QeDWFK,D24&cE,X\S)b,J0?Q0
_CPV4YQWP./RdB2F=-GJ@3;c-=+&Z:Y7YIZI(-3dJLd5;3<O9,_c[3b+N=:(4:JF
V83/N;4L5P64cB.d<,89QGJXVVZ_E(,Q>/,1U?S:]<,X5fO,X?TQRBK(OC[E..[?
U2IC-A#NI-8#_46R4>&)-b#G#V4-EbALd&M/[A\70WOgDa2MN>]9.fZ2Y,D]17[R
P0^0Id4\e5f1,,,WYK1Od3?XSL63GG-:,e5^I+IR.WJWfPR(3?c[\N4OeF[HFC8)
?L;7gHc:+AQ4+=?VPM&#>c..,KdM+L]IT_85gf&W#NCNF&G[RG)d.EUeHa-H[R96
3(7Z5e(/J7b=;/IW0#O,-fGfU?BDEQ/#dDO9SbT]LWTP_M>\M>.0W._57_CgI[A]
NO#37F&Te/-Ca4NQ3:=KO#Db]U:-<)F1;P_>Y\Sa3;?/de_AP\[Va(L.?E@WS6E8
YZE>U6Ka8B;5D9+W,^O#BFSQ1aW<#.@[8L]=-06_(@K]\B[UWOc(\D-O[24>JZBe
D?MIW(KHd1C=W5@f0G]R8R60]#)6GU+^ZP^e@KQ2c9]#@N_f8.,c,[@;1]MLE#)T
3E[R>+2NWN.D[HE#ZCKF]fcM,/,6-VJO8,3:_EUbIJ(cIeK33M>.XGA-+S5:gS@5
/]@IFU<300(7M?RO6?_(=D[eWO,H?-,eZE<+YU5.MHL+BQb^(1<0N6Z/AN(HELX<
EOB4e[^W=6gfT?.T;-X\Z&)B0/b__f)HO?T+AG-/5NBH>39)UeH/R8O4dE9QF.>b
1/6P2OaTV/J[OY&&0PEDU)e?TC79JHZc8H3KUa2\,aJ)@>[0WSSI8Da7S2Jd>P<Y
&O0(+3TGKV#,g6R,f]:5MR42.A(WB7SW_AeAQ8Z\@/@2?.cSDFD25CNII-Q]DP^E
6KE\N-5SNN#I;GM&Gea[gJDERN0_GZ,DT-V;5D.,<f.Y9dL/49<^dAAK)#24DTN<
;1<UX94VWE1TC#\M_?Qfd0_V9<&V57B6BW[7B7WORUY:\e),)NL9;F87RXZ6c,D\
I9dP2E8<)RGT+\-GRP8F(7/P6>NM>bH@08QQ0PeO#T58CBYD)Q_])dV=d2D^UGIY
a:<7aPdc\YU=7T+;S[C+<,b?cD8=S=8Ag):HO7eNH-Y,a2PTQBB<-##STcedSb-C
X60T0#gbaQ1<F=)Pc8XOMfKV1PA4gCYV25@@IceNH:Ie;/K/80aG6b1F=O5\\92]
eU7Y:N;[]YK2DU\[C4QHg6cRN[FN=V9dXaS\E)eaLXe7S:5V97&8-;e9UH7=08_R
>X1Bgdf>.Y+U3eRH3Zf-RJ+;>.BU[d-WL#ab_#f^CZBV31(#fMHf7gccXY7fMZPN
X>YL<gO&1-Te>[87@EIYGGCfL2SK/?L,BOI=G841D+N;@VF#NK&Q4(ZcY6<Ec@Cc
,O:>eLFC49R0c-35?O1HR(:CIIHPB7^[eYURTMYRL<QW>[dF1,0(I0c=W\J[&KG0
U[PVdQ]XNbO[?:a4&d8CN\E>N1,N?7Z#fL;W.;&/1Ca<Adb,Hf]9>-SI):U,bB-@
b1SS9g.L35c70+T2/=3:\9DPcCPEg1T9];A.3DDSe42LFL/<,@5D;)UAd+dJ7EQ9
TJ<8F(H_JegfT0Xc@=N#Z.,CQfIL?K@4^;DaX\=1Z^ZG.C:N4gL]:gKfIZY:cPJH
]8,[?S3GJT][DW+JIV0?L@b@?c(6<XO.FBUOdF-0V8:.#0D4&dXcDQZ=#?A8)WUV
NBGH[H/ZKB#-a6e^ZK+GE2AZ)K]G;_.7f<K\Dce98U@+ZM=L3]@9b3/>R+&(.)=K
0W(_U.P).VRO6\=]2_R@SLgL:RB3;:?WQB896TaDRB:\M6?AHePdb5A5gaY:?6L;
#B#==_1W=]a=fQ^+LG^)V)NMHAX#L:>5AQeTDZ^DP+a\O0^NS+EeC[4YG1[-^TZ]
>)V,,>;2\?(#EMc6b]<AHK0cUKN&4a[a,e@Y>>bNVeTBI(1Zd7QC:dCFFGDbS^7>
K(QS]S0a?e_UPTe4F7D/D6-VP><0-9==5:-5dc0f9D,e<FO?ScEI[9LJ7:S5Q@^=
EM7f9YO[,&;@Vb^ZA]PC_,N;[T&KOV2HA8^dWSOeMR=_,B8CP_R6^-f5CIg]gX?O
7c=,JU>_3I>0_LWMC[c?dXbI-gc\YP1CN:]^VLNdHQ7R=1aN8HI]KJ3[E2fB(6WO
^ZbY)Sb1A9@G3)6SHHL;S.S4_aBaBC.ce=H3+]YU?PLaE-eDKE2VQe5X@+)D[LM7
1[@BXGe5#@F8@-OX=#2_MBJ,NX;dZ+,:LYb[5f)e4MJSPDU.Qfe/@@]#:H\4C_P?
cOOb@)-#cM3T@/6GLZNY;+1]b.?PQ08,-XKEY;QZN#JF@(Id]fd+@Q(4ZDN>f><5
58DWI)<0bV6(c:.@@7af?-c3E=_3@6\2)D5(-KX>C\?f7/LE>L^S7[Rg+>,/A)?c
\?=;cc=&eGUbe4>BdH>Ob]H/UA+1f,;#L\Y\Va^6BIBI?f>?TF9SJG_UJ7-L-VR_
Vd9\]@fgX8FcCJHP[[G7a\5bK-CV)4O\E7JTc:_9V5eV(C-V73=_&5_LQbQBU8).
S8O[&KO5,5.<5aQ8c?a_Y,&HNe3e4JCGUd9O;@<^J3C4+\+[27K[\::+^g1WJ0+[
@7EaEf,cGL4<Ib\JN9\SPL[8TO@6O7b=YT[=1g&[5f)</SK7aY,F=QgQg-.H^L?&
+;>IZ7L(#gG]I&L?-K79?ZUg#E,H@NPILJ.SVT2]2-<-UES-eUfO7#,f[COG(6=?
(eSP#?b+#QORgeAP\+T(3eAHJ^Z,X,>X/]&R+)g9DA0\a\=9/eM>;gOXY>H>-J5V
ESe8C.,BSTG.?Ccg[V/:^=O8V;bXH[b14IR^2U8E;X6L\PT_@XW^]CZ[;:1AS^a]
M5,1<@/I[ZORXOYC7e25H4V@\(XX),C=0B&+/IDFLR7.EJ30CQH=IL8T1/^-g^Z0
.S>]3^&##c1KE>,0_gd994Oa4RUd7SCREM&;aGA3+fd1BeBP&baaG.P<&9]6NdO:
6(^gAZR@7Y0=E3<N#cZ4X&WgWTE).efEfV/3TMeH9G0PC^H1gf1X0.Z;3KCg7Wb_
aQ0,>7B>#6T.5QDZ5-229HKH(bYQ&=G70-+_&S91a>H#V_J\&0<;<L-ScG&O-dg\
e6GB[U<&EY?d3G3bbUVC^U,&DD@<B+38,[;2JA;LGK:3D79cX9[:N7F:A,#J3];J
J5BUBCNOa(_\V/U9fNSfZINUf2f=PAM&70b9E)EEWD\^0G76T2,?:7dG90U?U?VL
>SL6RD?Ig,RD++aSRZ?E;YFN-ILT\J#\KE=e<2()OS#5C55Q,VeU66+2P74[C,[;
U?M])GBW\c]Y43fN9UL01gDZC=NL0=B;ZGU-3,P),a@_5U]>?Q77.?[OR/,#\cWS
SF=J1aO+TaG;7)]19N^=H^#4-46,^Eb>6_#-eM=2bD:@78J?GFBd[eef=DNW8UP-
L?LC8BQQ#:6Ug;Vd4+^2_;RC+9e2[19</KK_2NJ-O^L(_CC+E8-.M1AA<PHCHPY/
9;f9c)?K=)E3):BbZ^XMTfVV)L?<ZaYELbc9.H)XSBI?b7(4:X8_BgS.QKH[5NAI
1df:TM(O_gPa&1@:ONKbHPOFM.@MV)SLE\Z;KWd\cYG#Z0O:,NN2]YMG24<d:+1K
#(=NVR;,^0VITA2@Yc+E+8cB&0eEU+0HOX.1JR6](A8J#.\(A.PgN4dE]gMFNJJM
c]X6VXSg5E3L+,]RN&a]BRW.F[U_B<;#a9b/O9d+;QVO[6E^?ZN-5Ke=6=?)ON(;
-?F9ICV0dT0.@0139F4O86WeSD&>C<F^_KAe8N2RDQAg6M2XG[TUAOGW3bea4f6/
==^:+^ZXC^0+VZ65O>e0fZ/Pg+J1>]/\g)f0;aU8d59^I9cC<DF<RK9#DS=SKP9/
9YZCVEK0DK(_(VOWPU7PBHN[aB_BMf?BPWD5/E.W;^Q;X=0d0Ib\WcWC)-_?<+c]
:H:@PM1CZ6@E^I5276:<<LA:5&@G=9YgbKSQWFZM_U5QL9[;GJ/#cK1&L<7e@B=^
7LeXBY-+@e(>YAASg[2O(Q\J6ES2_,fWHEX(<I[X[HVX^O=XJOW/J4LBLHN(L-9\
V+L]]J^(_1b2g>KbNEYELKD&c9#T7Z0>R3@J&BD&1FU_DSeQb>>R76H?A2_WA>7>
d;3LY&4S<WeMdPLaA6?.eU;>8EJLL<AR-G+0(18D42RN9bbgDYNOaLfaFO,DYI0J
67HgVO+IaUS=C?1E9:=WB4YDD-9V1VZf0Q<R^[Q\:I&ZCX?N0U3W558&^((4\3V<
#S@L9[/O2HWa6^\AQa.V#@VEFQe>=L)29,^XP41N)P0Z<\&#_&HXWYC8YXdHA)9N
cTe&Q;cR^6<&5DgY#cQQWB32=5V59IC5/OU1:]^V0=DG62P9Hg2)B8=U6(),Fb1U
R(BWL:A4eEP;a2:G8cTXYBFC3Q.b4P[X-Ib.^fdS>&E+1S21[:8<?A=UC^?OX/;^
egJ9#cL-1f+QA:OZ1GLO>0R\4KJ:;d3R7R2Z+YN2S?>.CKI<LM?gF;8^T2\O;GgR
@3)5&IUKI=\)B6C8?2F?/.S[TaL813^-46=)Z8V@DVWa9OEH[:D==;,.7&9:0K,H
_J&YU@H4aRU:8E>U+Q90dFG4gN@QU_Re7?<Xbb.2&6@LR:D2ERI59a,8M\J3^D_N
7=]Q^Zb&VO9Z&I88^L[K6#I8.K9Z?I2T.6B>JG5PK1\75XX7)X>+YXc1L1c6K0PQ
UJ0G,ePR60Z[g<I+f;Jc/=@_;C:E4GaZVTFZ2((Td.6000@_Kg^27C4)PM)IVU_T
G\eR_5cKY+24.-=L[gMVVbW1SDF2OFZZeZ&IEYT/<?a64JMdG7b&7(CK&9Sf?f15
Z(AO7?O(_6J.f<YN,[>9-=_>+4_d(9I&ZBg;E[>KEKdR\M;:]c_?ZQ[KF0P<B)#A
?4PfXC]IE9dea0Q[6M7bXI)X4KG7T1Gb(PXANP7(Q>[/W[NN?TGSgDfEWF:A/,NV
:IIc=_&PC;,cMb+@U.L8DMGKYJ8JFJg5F;@;,>\S++ZV1D;EcPdUcD9X)LM,XYBe
CbcTPALf:(LC&+M^7D6d[&g2MHdaQdTa6_JRFd#00V5B7KMJ35d3gNXFNP..U80C
S4<DNHVa5FUWU,;a\.(X;<TK-H0+dYIgG69g.0\MPN.S/W9ZA+6K&:T#Y_48-&AL
[L,482g:0a+3/,._a<QQd#@-dZ=S>O5[L[2=R5<WAa;7GPNF_Sd#geCBbgZAa0OA
@TRc4<-]9aZ)ddX?[N[a831FcR\.]8&:e\#24De<=,N4.\3B8<IO=bS]>TSdLbg#
V;.]DDW+CMg?N=R4e60X-YBa[BbVN;F#J\\)J>&)(@[E[GAHX_JYXG4QW+>6Q1-C
X<GKPbI>b-=82]PWV]^T_LCD=/2ZcL(SSLN[+?)LFD53^ePYRV5UP\f0B./O=]<7
,a:ca,^a=^<_[6gcd40QMY0;6M2+gR,]0]S;/L>Pd?38/#bPN@>&71AFd5MGH.F/
cDgF8NAP1ZD>V6JKf&)d/SE_LPI>6:9Q1V+-DU7L2N?W]d+UU2JM[b(3D#D,9.(6
GBIQUG+]]D[G+I430H8QZceLg2VR=,&@0,XbI5Y<ATJ5-(QB_+\fEM)=e+ER;ER-
F\;L.<(BZP^-+];1(=;fDRE7Tf/Q^M,1)^+deDMPW14UF4I2U2NOU08-^RK3C[\D
;:V<=]D;d(;^0W@<[U@GYV_43C3BJ)1BDYPX7B_QU2=5_G<^THa>M._?R0MJgWXe
Va?+JR19Id#:BZSIF9gT5EGU)]GA<9:Y55\=C]T,9#.UP?B;P5Tg7b1N&D)K:JRV
0^/3\O(d-ZJW)5^2SG>eD?34ED1?^4M>NS81UZ<\Z,fZ5^_<X2J:c]PIY<:M4:1&
ES71]E@A]QK/:f)]^ULKFD+3^Q.@Y/5OFGbO78Z9H1Tb7dVE,@c6Wd?(GbaG.\(Q
YJ1VHYQ.W7(D>LeNTe-6P7XEg#;J@?8CgZdfUZCIKOHTMWZA.G79b>Jg89+JDOY[
Od9:N].eZR:=\.4ME#Jd\2<.I@d>eCHL6a-b..e;>P\BASg^//^NU<8c[P1Tf^GE
QZW1J.)V[0XSS.V8d.W2b[45\c(#F;WZaQMY\D\G^QFS;,F_[;AO2F;_dAR__KQ4
UY[d5XfN89<M,b18,eQX573\OYJS\3C^1#6]OVRJ14)BN1fJ,\]g9]N)0Lc1+C9?
F@Lb0K_D+#3XV,?B)]0BP3L4N#)=OLWIM[T81/L,4W]Hd;W3DAJ2,L[^,CS58;&(
NPI9O<?0;#.)V8ZT4ARA1S><Y^Pd<1ZP4S0:OdR8N:ffJa_(/@+M0=V_^=:B1UO?
@B^_&cY:9#.J\dfdM(P(;T+N.&H6;^Ua3B1#d]K)R1G:+0fYZ6V+G?H&775,HY[]
1B.b9I(V@4cS2<OfID>JI:+;J&.8b>,Z-(dNX<X1)\P\WG^XPVZKE--4Q(5<#d9)
)1b;O^b46PUBRHGG_OW&B,eA?Y^FO3,#@MObdT;4W&TC?/N7B#-4,Ce,R\fQE?T?
eK5ce#..BgMB9QM4_YS-]Jf=e:7#W:H8JdGM:7]G<PPR0XO7R70df&W.S+R()8E+
FJHe#33aI>W+Eb96gONgcW+V)9DV2MWd2CBdM1II11K=C9\a+4==,S4)S9gK4:A8
Lc0FICJ5GE\#DJ)Dd<=O(+&J@0UP+H[B0+TJ/d4R1\WPE?^EXN2BTC5[NP;IYed<
.#6MZWFSO>E0a4U20?.HI,V5BCL6?g,ZYQK9<c@=^_=N+eGbKM/S<(2\f>W.,+CA
fHA,eT7Q:ZOC:,1#d[YXK)8QLcRP&ZXT#aQSeE>PITROR\c:Q-@,R3463;604@2H
2\aZAVPBETW.^&[:.Z?MS6T9Z<W=XQa:D):DaVSR]ePX(;T)+4K.XR>4DTW2ONT1
IK7(B<DgYD.]@(f>8G\E6c+C?,@/)SA.UJG.#PEGfA=bb5P>\_@,G3ZZf4LRc/5H
8&YDIHB^\2TY3gK/=[@Z?]I+aT\[5W_adY0.4b>8/78OW-)DL]QEBB]BXV]6b?bf
/,-9YU1E3?G>fA5E1IM&9C>GK(L0_&6MXOd4DHaQ<K3V,Yg=8G),&GCI#FJ3:7Ff
DfJc755\^^TY)]E<2.#Va^.fTCbPM4G/VF)g/MGW.:2E-6GRe@?UGA41,I3>U6Ef
QGR.R8,(Y?B_L&YX\[+DF:)5g0d<1IXM?^4WA^^06&2UC+2\/7W]2=.C(e8S9BRG
PR__8P(aS?T?9c01+)]_.>21?HL-_MZ?aK+f>S)7Q_+5#/TG7721e1BF=O-GXKa.
HG=>TB9?Y&ePY;>bAY3PGEe>;9?gUZK;:PMR9GNL1+:A:,Oa,OI#;P^;(bY,9[?2
aCP9^CQ+_P4Z[eeIORI@9&.FEWg)REc#NLQdaGPV,-MN#OgEZ29R7U-g(cB:.d&)
VL#GVSd7A31A7f>F]a/:CPFGB^f(MHd+\@RAAW3J<BD),.U,RG?f\ET&R@49ARXK
SbEb#afcC(bQ+^YJYg@(JS[_AH>IERKe\3:K&ZY,2<.QDa9+=23--J&VP3C#O,R9
P>7^E3NU@bOS@T0@bcMYP?PJ4P/:3R8>M[1RP9BScX;[XY[.50==V13/MRbSC,g]
]-+4C\X-XV;M@+IJE8-&P&aBK8FXeT3F:P)=,,/U^6:+.=FK_-R>]G</QS=^S3H&
/B,@JMLOH<VTV0W5+GYAJ><b0CF8YC:J#)<3,cg_-2YB(9H=8Kd]T1.WLcJ?cR]J
[D?&_@F(C)+=L;00,LK-,F>:]+,MD0<S1NQ0^-ZAV2WRQ>9Ub13dZXV]&SCB63a-
8:9/PeSZd#?V60AFS-?0f<.VFF^)@7#DO1N,O0T@<PA-1/EZ0<57-\[H=7@S[BD@
2V8\D;#>31N=J])UPO4K[18=Jae,189eed[,-UJ2RW=V<F<=[f01T-JUE+XTB)Y[
V)VI1SW/<]DEDWbA^Caf&c0@C+;9fZXcI-6J,ZSUQ)+fC_HWK>bSR^1MA4HPbJN4
G.N<UeXEM^UZZ6\8AU-[#f8eMQH0O[Y;:@P/1f/7gV3?]1ZR,DB4FCPWHN\PKNS4
B.,:&MO5[&Q[,Wa\541=9.^ANBH29YeU0WL<g?^7,O]<H;J7>X.9TV;5?c\=9VQC
B9NI9]&VQf=M8:0dDC<9Y-MMe/^3=IY_NQ&Z1HTX@b9KA#2X2&b>B(#d+K1.,[aJ
J<fF?,M,,&GVFH1(:\PT4Ec5gAYPE-6T;?ec?5f@9XC@Z_./OC;31A69(9O:aK5a
A?.\;/=2e,K4/A]?7--M[d[8-F@f&01_H^E5H_ZQ5>^-6G.g#dW4FZY9O603>:HA
8)IXVX++LP:9#>eJKO:UXYJf^I]EIRDH17+cXF8/dSZ<U/;^C\62Y]B:LJ-g/O,c
WG3Q&=;15]J78IC5NXYG1Cf5<g8faUd/&K8-+S]@SKDD[L=)Xef=/B..&4Z3DQPC
0\V^EZ9HARWVgfQN+@2WI4#GNPc20X@B9eL8&A(S6@698>-RJ=e?>]9Uf/U1.L;;
SVYfdfXNTbIXOKM7MY5SJ<&6&WRMX2f)_Z>\[Q^];=V&/;a70-/)>?Ibdc9B?Nc[
1?J[Ib)+L5:cLWCS]aE/(NW]S+E@&[X]A0#-ZNPZEe?&?G1(6X;8[M,U6:O-;X\[
J5<L86-^,Y9X9b_;N@HK7<\]MgDG:NA3@Z8Vd6JF-=Q-38?;\09.XJA>:E/Z1#Yg
Dd8ZIQN>@4EJUN.FUcY5^E[C3?IN91=OVC:cbP?ZTbW^./)82])C3EDW=XcL_;E.
1UJ-AL>N_)C[^]7(09HONc[C2$
`endprotected
        
`protected
,=2F-_UIfGgN?Q.E:<F318H\5R>[@32UTdc-@+9L\>fY9EbG^+_c.)aOM04-O;CL
(,K+gf\\_=+,_FP3+Y3IQ^H\2$
`endprotected

//vcs_lic_vip_protect
  `protected
X\PZ,442/VU(UR6:Y5L#-62&7879=Yb22A&>9E=YC&+@=CB7TSE,6(KEc:Y)X1g4
T3c_X[(33/<fMP@@>J_5P8X;a_4L3Df04@M4.ATfMf;H69BK>&We4SfIWD#O(eR#
Q;[TGRed+-a)8/#MM32aOYYA0dE,WfdULY_>P)[D9M?g)7^Tc7OM3e?Z;NbNO^/2
M;M>_Z+IVW>L+/JXg3T+ad_L]LSQ>(@f\D#+L977AX)bO.]L1&_H=YdAZcEW(D&:
A,DTaM2IWYb9E/K\-41bK6Fe.&R6(=d/X2A=+<]X2Jd,]D-8WW2d@>2Qa_.Zfad4
;8Y)HS\fZ^Z)>NJY.,E:VFcA>A-R;GeAS6fLQ\.5(/a+9aHV1aTB_DJ/72_d#4#U
=1#P0e+/^YHX,Pb;5WfES+.KbQ1S<(VY+;?AV)J?#?:f[VSBeAf8U.CR4X8T?&/S
:,\R)TKc5I<=a.1F5OP3W7SUNI1KcB-^@6./e\eSF+<<2L^a;.BA]ZeOL?X2DMgX
YY6VT87>P(:B8EVDZSg;^YcT..\5X3P-HR[D#a#O6FcLQV6cc1=a=+)QEa&fb=&[
2+-(HbG3c,b.[PW8Md-ZLDYFC.]5T[g;_<ET[<H^bSB0^A3MA-&WUQQ;DDO=^56^
1^0YKGN9R\173Y6_?g#GaRO<G+3D>^d9D3YSC=R,g:1E(SaVTQPN[;Z5GbBP]H0b
+M2P_a9BS0>MNS_<W+RCMb)C::QV/V#P682UXddYPT)386G+S9QY3+e?G3EJH-3-
Y\?MIM8OFL8.C6ONXYE7&f=5N7VW>J.=2c</D0W-R3:4HT?[F0.VYD)YR\S?_E0S
ZPTd_^UKH)Ucf8;TJRTJdCe4c->VfcZQ<f<EL.&>N.WNYI53[\5YV<ME<_#YR3]H
c&__>:=AS<IDHSGa.d+A:>YS(L(Sa/&+N0bNbWAM<AK4g-CSMT/dW)]B(U:JO,cH
.=Be=c\)1LJ1MNgZ&(LFJYaU9bEX:<K[>MWSg4E3>2Jc0E/D/EL9)>Q-&4A)bVZZ
DffZ/FSW94UA5&EFANVbY5H&+MgLXYd;<\U#?4/J/ZZ\eCD=d&3aHQXcBVL0c6Z,
6]Ic18[Pg&.+11VESfR;4b@T2+\W9S[0(LL<UCN]I?&QH&SBLB>\-Y2D3()0_3.a
]\XSJ:#gc1Y4N2S0T]#[<G9gc;3..)AW/HEcBbO2R1/;IQ0..]A)6DHcY:=1<&.K
7FcIU&Z^W=T>CI\;,,WgDZ94MIgZ=V.gV3@C6C?aMKG+25^GF<_#<^#&]HV)YT)?
Z02VJg(IZ3/SAWYN9DGL>;67:/1e;_29gX=e.]3YA6#._KZDL95^&7H6GR=?,c@2
]eeJ31fdUb2(/fQI<6?WJU>Y2-+KM\F2,]]U.D#W\#bU6&;7e80[D9<0Y_)>dRGW
B3N=N[-_466^Td6=4@Dfgg+O\8Y<]>0;DAJ>?N1M.VSS,MOG5WdQ5961).R^O6]Z
::DDCa(L\N0P:R4UOHa[.6IFb5:e:WPZA,S:5>5BcISG=1R=OPS>5b]PED;8#:4d
2c0HH>966J1<3B_a1b+-BI+FK(JRG7UNG>#Q\(_+6Z)Y5b,-\52^.)6O8&b:IR<T
V?O;7HaC@R->Ke?2]DO@E)^PM;;F&XI-UEg=7K,(WXVQA\-Y9dEaa=MYY:b#3U;P
KP+?[E,S/9)VZPTEd0>@-VTg,+P[8?PXKA@,L5<_MY4AB\/L=a[//_=Z0X>dJB.H
a<P&/&S73P3W4[ATY,8:ER8ASDZJCYa&<;(DZEPc.1<U3PW.^OBU\+.T@4V)BLD-
R)CHOfIA1[:g)FHeU0da>CDW;()#_\9ADW5#8EK[-a&MS8^KR?1F9:G5_XRX&4M9
gH1K-^4M/F4HO99GAN4a-^H1Z@72dgKa+0a>0UaTKJ+]S9f@C:.Eg[WF]\W>>;-2
fIXbMaX7Ae+O])8LMNge/=P4B0>[@<bA21fc0L6_?]:E>fAUg([6b9e.-7V8O#&Y
<HM.Dc)R657RJBdGA(L9][MNDU#CJC#:MNgP.SNg:eH@BQ.B6O(NPB4P9G>_(T2<
0eaU=U.4A:CcI;N0<L(NLT0UKJ.-/]f^T7-97#?bIK^9aO8:)>3a):ET?beR)eV[
AS,Od8>d]4OFd1@,ca49F6&1?f^E6D8b?_dWM\Z6f.7\/NN0c&8>A.0R)+e9=TTG
L7<S?WBg7LO&XWK1DOZK^2),D6T#Z)Oa:P@SaZOe.I+N<A;8RSYL1TZ\PU3=]:F4
CcT<PU5(L;AALcV#4>@[825?RIYJ57L?Hg,G[RWFP@PHB((?b<S.W8cNVeUHB#4K
/#A)^U+aCA9BaM\+L.4SD-O8D&H5<UE>a7f^3gF/TUAW\PRL5O@/0@)/@GWgUKXD
H_&,3:J;8g_gIDQ,_\c)#AFD5LZVB3H.cG4Z21.A+^3J.fIEE.58^?9:&-W5^[-&
S0P[,GZ3WPP+,\HLKL+\^D/Wb@F<5\(<D?49#6>]4B2E(;MX6FV4>;c4gWBEG]GT
Ag=Q&=7/[d0c\ZRG?eUF[=G&OLQSQ]3IG#7?9P@#H(WRI5F@RV3QRMb:0_>,fS5g
dYYQ_b)J,aSD&QU(V@PE]H@/Gb>D<-ZJEWOY<deZY3P,Z.b38+YR)@941L6<;2O\
A0C75:@MV#/b(7cF4V3@ZcAAPOMSHM8TBfB.bYB.&?e]f#RQ=+GbSgYe;F9PNZC[
;=3>3PK5@aGMX[3I2?bd/BD3U9M/L1e>?e6e+Q]+TJIG(d8cEM;bX.;4>UO[/=>P
RQ02R:K?UO9VZ+PF?7#Q\-/-EWca_8^JaN9],9F/V9Bd>YV249L7]+c:[B]Ec7=G
?NLQN(J70?dL77f0#?DS[^A]90YBMVK?7fO\];HHN0f<=JGAdAJ\&)ccH_<EUP;J
.cg1M1DB(=DcO7;KLKf]1B=8H?W:SXe(X4N0:;Bge5=RT:,X2WEFRJS^Y6\/]YGB
83D];UZL?KR[U_K3:VM3_;OaGga>AbOX_e10V@Z1b/S6>(XS9H76a0Rf5Oe4EdA[
,A4dJ;BYN:PXJbG1]0/6P\b<XOc&;I<WA3F;/-M#IaXPRX8[\7a@GZ]a^DGMEcbA
A;JHS3cH^IF:7RDebJ7CZI_QN_eM+La.TI^bO78?368<F2?/HEYb\Y9#<bN67BbE
V[2(bK@(:J)Q#D>&bH1RY;Y#_,V@H;PMb8K(\3>KK693698=7)(:=>cRH3GDK]gc
UcS2f&\N3,1N@TBSeN;1B_WI6Q_.0a3)=eTT]E5+#6800:+,d[S9G@\GXKC539(L
M-+6,7WWIZH5L0d:VZ1>>H8W6^1Y2R@^B;(=\1\_)(Q=SSGMSVKYPXKJQ?(\f\]P
/CN:603BMUWZSB#C&WQ<dA\e^[1Xcc40W9>^_)8C\1U(EKC(^)1R+ES4J[2S?Nf7
c:bS=YDJ/S)?8J2Ag2NJB>.W\PNBBH401X]9PZ-,OW0YSO<B,@_Ug)C5bCQTMd-<
2YR]\:T?JYCR6J2>P,ZM6D]ERI7g>N5PL6Mc1#ZZ_&-JJf&G6eG:b[e-J/1c-KYV
Y0UO?a__./LFN3fJ+_]a1Y6Pf_^EAK&g<3/)&36&4Y^;VWF\RJ60X(-J6AI(Y,SU
O5BR,gZ1CLUGS\bP?<NT,[c3P40LVO^65^92]>CZ\FOWc+5:Qc^AJeCBBP<VN>c/
.EYGXFJ?SJ_?K21_[539B77cZS[UD+)57PH1JU]SUNO8WVJ[fY-:-9#+8P9&fB?A
O&fVQ^Z^P-Ld6:YB2^9SdQY&Q+S:W2gX5L^c1G.</&fY[b#N=EQ+,-:C;b(0_L=1
@G=UFe88<;W:V+AIIc:8MT7E,dfX>/aT\0X;]G+O7==2JH[<HO03Lg:5OVZV[F#P
?Z=HR26\)37LCFaRVKg:#\d\C<M549_PS@C0FI8O10@PEAf+b0a;-1G>Db@Sa8YS
E:c(_TVA9cf8V=Hb7ReL_[XA<]2?4RY]g0/5K=a&<gHOJ:aCN4f&[Id9&gQMDX(<
<LMQ(c3XM_TJ2&-4)B(ZI#QVDO/bb)aXC>X8QLP(-YaN75.^TaP<Lg<,43/_URI[
A>9(Q>]B4^+/P^YU\&-E-6F](+P#OB=7>f7Q+[N[F5b^DePV#]A1\D[H2.KK>X,\
N+26SSK(ceH0A]EH9B>JE>Z^TE6FLT8Zd-gX&7NN>)X5LEDcI8K7Y]W\U04D&-)f
#V+M1>H0HS<JA16CGG;_IM&e-f;E069)[E);4g88E54;\O3E.^IS9MbX9J;7UJBM
Va/,O-Z,4L.[1T?FM<I:.BV(V(7^RLT8H]04\@0W^cgLW5\94DK^9B-CWCfKHL0B
Sd>CcOe@\0_GRH=FL7[@1N+NQ+aQG&B7_4_C8O/c4WUcKNC:1gZQO;&AOQ2E@bQ)
e36ePZ&):W7dXHO#L\[K?3-,6ZbJC#[?4a6X7TfB:T+1+6I4X3HJ/J8[<:/U2dXS
5(c3gMD&J^+53TRBN1WN(A6P43.ePXN.83@fIgTTS=+08bXB+NH<bF&V-dBdc3R+
[O1(?O9X.daM_Z-HUaG)75-YQ8V7+La^1a=#B2,X/B9b6WVZ-,4FA<NW_+-0;P8L
XD5?e<WFY^;?USVL#WPZ]GTZ5N;XG8F\IdS,@<LJ_ZL]91\5OV@fX).Wfe&2bA?<
<?COQcQ(9@c6#gZJW3Y)+9JVN_?+9HGI]9;R=<cCP2[agXEOH7aBE:9:Q>Z3c+ML
_(=DH^2<Na[AP4c3:&-<+WGBA::DX^75X\F=/WXUEcc><8,[3KaLV1?APKCG-:bf
:EGNI@&OFF066-.c<>OV#a6]bM7HfJc#I9&[BOIJT-,5U\VcXVMc<>.8\6)FEa;a
/6CW,03Q4a9dHTH0EN?G7V2.RIVC:[>?:3Q>7b#V.(X1P^.aCZLEbTUb^bXF;O4H
(:@6c(#>=ZPKR\@R9:;,1^K6\LV/;MDGEW1@U@T?Nd?XbgX^dFYD@7)M5LGJY=^E
2d]CF0.9bgEI6B-ONZ85+cG;G]_BOD0FOM_T@HXX_<]F)>EQ3N<>)-PQ)+#eM>W_
S&#JV/G:<\Hf7S:S1D:_C,/2(G]JWT=1Ga[Y=ec#CS36S<0TM:\J4LY5=VR>Q[LL
HSQ6SGbf&7gJ)&g79O.UM9[@7aJ=#Z<9:7_W<3HHRN1DC01#=ZC64HM1;Q:E2G)5
J5Je/=EO/F]Q/)#_F;#S(RM/EGOJbYP^@MLFFW@T72AV<b3_1AK51D;MgWSdSI[H
+9d60XZ8#2..[9JLC^+P.9dPWX#UQFg5&)[VMS^C,1L]f7V]P=-)75UB7&<DJOd9
7VcFDFOC_a#CaX-Ba,fK6&X-W):G?4e)8RM-#b2YeAEFP;E/FcJ^#39Jb[Q=-FbM
/R/>6,Z0-28g(B\I9Ec16Ng/:U0CbSOJ5K+5MTHN02f<Ne\.H8=dX&L-\[W+A_;+
X#c,K7a(&X:C.&T81WYD3(5NW9YTW>f1.<AKX&IS=\W,J\KZaBOP8_fRHLVO.RKX
BK^#e(B?5GLgW^.;7N?3/eb>aE51V69]+V8fFNf_@LNSH=]&MGGM9?S4.5+1#/?4
5KId+bIU(Y984OK=48La&@79@NgL0fEG0CU<-Z/FeC\V0@g73.Y2,C)Q/]:QDgb8
LX@2TK59\gKJOFI/,4()U;G?U]6R1>#Ef10[#6]/_[_@DJd_#<JT?A&Zb?3H?TMS
UV9JaVTV61SIKZRI)aW2#:.L3<Q&;eW?(.8&OOY-,]CE/4f#-4[P:ZZZ,^.S#d+V
BGX;bYKY\9QFD^:g8O@2V?8;^-0L]Ge5C]0R7[P5-Q?<d?():=MOODO1A5W1MKX9
A&VY4:a=_KL+L6M_+>ID?N3c;eTR6Ne.H=94cgS^-cB0\F/-:L7&V/T\&ZUIFYS[
F-e?/cNP6LOf8<W+I+U?MZ7(L]]-QdMe^^+#(bVBXJWW&)/>bOdEE:>N59?BVJ\3
P&0IU?#0cMIJSI/S\,&76^\,c&ZBfN3.GcU,ED9(LENT:)TgW\@@Y1=O^>VJ>EHF
;=B1Ec#H;N5cP[VKCNQXN,\c_^49BD]^>]?9(T6_ee5aUG]QLD^;6Yc2@fFC^O6&
?/#T_#BG8_@Ig/.LJ)0?1UWG\]6Ze4H)W;WH1_(DPGZb^EaD)R]d)0BU@B\8Ea1,
)-;^[,>OdBH?:+?T@5.Q?gA_O[UCbZ2)EFdV6.TRF/#eYB>=f/:d->IC\P#b552g
UI^]Y/XD<>agCKN#N95=G-HE#V?PP4eT_/9WF?41+WcW[/](fQZ5+Z[CC]#,F0-Q
U;>>.3g9[NH,?.A?6bd(Y3,MN&N?cV>]d9g^QI4,H+1<.Y9TA[OT0bPV6e<@C(SF
:#a0Y;0)4e<ASaHbT/>4ZM?Ya]-Q=4H5&L_/WBO0IL8H^<aK#F<4B3K7)bB54Ng1
dW.KXX9@<6DO(/CCDC.SYADR];?WHfE5fcPCUTVC_W>>2@H1A)9]:eHX[LH-\E:(
V;)=,:82VL<4Q)@>:N1-]RJ]5QY_JH150S4eM)(J[cY9KP:cJfM0U7PHO9^X>J^Y
^9(&T#/J2>6(50;+/GbT+GI>YKK90GbARUg;@aE@aE)Y4^60W2(fdg#^MLH<&7E&
Gd7,a].)Y>fAE,I>)LQf[J:A]16SQ?4GY6Y:7^Y4@36GUCK<@[P^Z+-N-IGb\?SZ
a0;e^.R)e#9b(gOVDJ46[(E>)N=_KfRK<]^GYC<03F=Z&:L-b3g),@#eV3AKMb5M
c<ZP>dA4JVY)CVLX6Jb<\]PRT(U4,+9I=[PA4,MFa/T4Q5O-WJ@7#TN],(/CXMVa
U@>\e;XH+3G/]LCY^0J@5M:\dWeB65H:EPM_AVdN,#+=U6IZ2fO5T_b3JUF)G;O>
)#S/(.Z@9&.FIJA)fXXOH@I.IQL:N@D=3U[JSX5(XMa2HW>G67TA?V]WfT:@1J]O
a)WBJ;(&:W#d;IO(TRd_CK6#VC2[XZB[6:43D<<1X38>(-:cgQ.80TfY=WdD\FaZ
TbAPD;D\TfTEI\R;VgTJW72K3(5L>38e)B]4c>M-.Gb4FA4^=;Q88P];YEfD\]+D
YL)WIN:-5EQ;4K=b6;Qeb-?KQ[[&;IdQ3>c\+ab(RPP(0b@77daI@NA7-WDg6/g-
@>H@JO,27_fFKVY@bWR)=_CJa.;8RKc]UR_8Bf_@I8^F3a1Zd3_cd42c^JK8Ud=K
bWgO5g)X\<[V6.H<RNHg:B9R>9@,K::M()XXHGT^_=Gb=?=CC^1\A];cIC#:Q..A
)1-/14)I<a(ZYMY<>_C3(bC+=FKc3E<\Lg#9-3&L^;(d;V4a877#VJ&#K\S-OdL9
_?E+FM3YJ>LN7LQ5YS^ILbE^]9LB3OE/6L4G.F87V^+c<14F_MS+KVB)UFd9=1XU
gLgYSO1^Z5>d\/\<O&>Z.B:e6](+Sg_[K#]c<)NeFAb(bFK?S?dNaDH@2]H3X7-W
I;GC)-/EC(5R9WAbG)?6[=.JYc?9?4=N)H?>TOUZ#7U23a3IU9:@8:R3dA-2dJOH
[0e40CMS8.8\D&C;@OYC.Q<.9?d^_9TYC(PNbWF@D.d]F.W:I]ZY_:f/.IT,6?C6
VUf9BBYHHB4&1K0ZeO=f@A3.CVEW1f9<5e&/E<LH##[LJgVQ=UK&FZ.MJ]=[C-dW
7E,(O18U@9Z(abQOa#X<Yg/08?R7T3)+I9(K25:H.6PQ0CF+a?JU<;&-SW;WLU54
[=-D^d?&6JW>U&KCe.]d@IQ=e0AE[KZFVSU3YK_I)CA7bce:_H5DW;^^U)e&FR4U
B;[Sd-/^QW-,8UM,6UZK]NVY-,,FB+c,>,eZ&IQe[[Y4]2:c&RgWK(;KP\2R8OPQ
I[Q)CCCP(44/TR&SNF+ba3AQONIA#7X[;I4d2a6,.DBGXPK4L2^ZU\<ZF>?&Q4K0
\\9SCSVbB5f<\L+VEK(Yc#QKc[,.>H3E7A0?g8?g).aTARA_beIOQ\I9EV>)8YgH
(Ba\]Z7H&L4..LD9gJd0]3J)^GaPdQLVMC2R,&>2.^MK(0YgD(S<J\A[WAGcU@H-
DV4\;VT.KCA;NT,?G7BV^G_XJ3gBQa)be,P[#S?Y\+6G)c[J4S<@U3;/b-YQCf],
QP_T,b+1GRM:;5H#dNW^<#H)]+N;^MY[(;](;,/54WTd&YX:4GbGe7.UXGR>UZ/>
IUZBaD,da@#dB;@(/PJU)S1[QeM-8??Cg24S9?]B5\WM72PKXHUS=PT//<b>.73c
G\<>Qbg6:(]NIXG02IYTAD]HK#QNT=V\Gd0NFI50/-^4c\:d=A,)Db#50#R1&Z7>
/IVN\42;,[7Y>f]X(96[PNfWRU:f,Z):#V>Z/1)6&)gYRE44efgN[BK.eOUF7e2g
AbO^-g\)1a(K=_<T_@1=J,\\9M?<3GM7L-Fd,R^1JSCP<(]UFfLP2=(,6RT41(YA
RXJY4Ba:8,U?MDV&cMUPOA:f/S\fX-^e=O;U7X^XL]X^+1@TF/ME5ZPX8GR@3.eG
Y9cE(<C^gV0I<)=P4T>=[FG;>ZJ)7G/-NV06SDEg]VQAJX7X2,8TG9#[QLF,_:.,
^OCHOHZ;F/C->,5L1M#a?b1US2@;\eeNO81D(&C;81#MQCPE>Y9.7HRF\f<]E[5Z
/G<+]Fb\=E>BH/KcaSOPRgN>g38G@V27_@.>HLVUd>-ME>C,>;RfbQ[Be)S(TK#P
Z2?+BYFMQ=G>5>HCV<=I2,V3;;G[IV\>20I^.NK]E,CeA,O8#N3Q&MR9&R>\/;c^
LY[f@)2LLRS<)\bc?:C,ZRL=&4XdB\0G=e.0>bDC=DU;9T@&,GJa#Ogc?a07@5V]
]Q=<QcG3/_C5f7+M0F+Y&[;YMINbBH0J#e^Y4b=b-S#4<D@adTT>/D@JcRL^0AK>
aN5,Y_<<FLIS(7S2E.].V\DC7fdJGb[;=6.S[IV29:g]:QZdbALgU-0-K>-R/\Ig
]MV[)=QYKH=UQ=g2f4JD1/2@_7?R]AD:bH20K;NV>]>KPYA0,BR8c[Y1dZQA8599
>Y)?AC,Z0I94Z\O3_<,34VV9c0V9PRK5]@^aA)DXY.ZGc8K<4B\7ff]/KA>L#8Pe
HM:JT7N,>#e#XZeDf,D0D:B>W=P/b#f4(cRV6<?881RTZV/PL>C0IPQ:<?g_PcLD
I#,4#f5ZL^;JJ7g\cN7dLbAc+f,#3/>RXE^>XV-<DRUCC&G<R:VL,bVYY5YJSLWU
TQH(3)#Pb]8Z&VJ75.gU0eURIB4K>c-[\#,.IY3;-.-4g7J<^NYF:9@&QCdNd7)(
7[>V2[,-&_eJVd;47]dO17De:TWI4XE_[1NW+,WMZDS0gF?:B/+cVQ0S=0;8\_31
NfF?:<CR(eXCQ60]e#,#Q.<R\^^).HY7-R,[\:DIMN=1C6(2b2F>aASd[D-\@H.S
W.;52;KdIVf;&.GU)0.,UdR;SZOcY6YVX:IdQ,5CU6?D+:=\@<P&[WPfaWZYfL1=
D6W0RT-;11^).LM,f4VS,1D<L-2&:^;&VaZ20fEC7V+KS>SX3(Z[d0/^(:?=@>dP
fO_:/=&23X:T^Rd0_6NR5@\/=Dc?@W,9c16(CS&>93KWg0-(;_\Y[bE96;,]CY_c
24d/-5C?8a0DfM<c;fa^d&9bY1C5XSKdPRf<EVGEVF/WJMg;1E:\cTKPIPY2[A;=
V1#,5=JcJBGH#4fJK+:F\_#=6>,O4)YIR<>BD6dXG&g1&UTBgVQ=AK_\=WSLAA&L
UY@7]KL/C)J0K(,[(0ddQN)-TeW4Z#F2Cee872CEHX>9?ec;-SMW\.HC(N]Y^0#>
>;:D;(C[6gQ3G^YKXJ>gb8FZ_X+GcF;^[@=H,a&H5Y;:C6NC_REc.)8<J+IYPF:Y
R79K0-RXX4Xa#5L3ORfa,IOBWZ?>GMXZ[#OR@WD7b)[RXFUSg@Zd>JOK2AL.9a4U
M;\M1HP#;aAO9,S3:#X+(MH4Y6ZN-0@;EYRYA2KS#2YF2D?MgW_1))gAY50A3)7&
9c6g2H.bKSb_1;b.P&c:(O]L<fRaG+=69Qa[[e&::VMO:MQLW#GH[)fK0._GL[8J
_+Y>JP>aH-)VW>MAN>V/gE\Q=\g@,L>6_9G\Td)=g-3SFXAeg]XWY(&BSQMYJc[C
2M:1FZfR:)d)#\cKY3NHB#W/X4af;[A8=H>ZQKR<VIQ[>J(bC)SLN2NK\K5V\OOL
,&9VQYEVF<Ka^@5@-RG.587)&2?_J_eQ\N_4QY-;a:3-Y&TL0QFI7[Yb_K5<01VG
Eg0-3C>-V2#d1.3bE=DOFYWNHAVgZQIg(,9M0M;N10g>>UG4.b-@J?57SgWK0O]@
^&cMWfZTO+FN-^KW6f\[AEdVXO5L\:OIZT4[0#g)QLI-T2I=9(J[,NHePI2J4Be]
7DSJ3UN\?b=1b^[/2JKdP,]cM)4a(g)(AN062ZB&?619EKXBW^0VKW=A(M\JRX?4
]W7[4DY5O:W_^[JX36WQ?4dTJX:X=I<2O)Y5NRX?W1FY9W3=8cV=:Q(X#&JNF7Uf
+O+776H0FH^F/=fARZ:PXTYYd/16ZAA1CPYe:9_UWfKb<Q#FEI[7fbLQ]M9(EEG<
#GE:<+);=810/)2MG\OISMU;.Eb.3c<>Uf<8ZaJX:0#=676+[0ERfBLQJ$
`endprotected
        
`protected
P5Z6a^LV_<]<1d]QLT^,,J[@9M\:H]^^a9/ON;9M-FfU2+]R:F:&2)@fV-+\L1MO
/\MF@JJ;]NHHC45VcITa8;KfT9;&&FfA)WO^4=eR\79RRW6&PJZU2\@fJ$
`endprotected

//vcs_lic_vip_protect
  `protected
^(GUV>e[X\:?55IO-Zg+MM]aa?e>eIAULGGY^:O=8a]CIBL#1^a?0(T6FHE4PJ&)
>cM-6fD>[U5AFe,Q04RgQ-9]W4G&S+aTcNfJ;I.1\L9]#5]4HO7C/FP4-_9[<ABb
/YH((J<NH]MS1D4Vea4[gKK&KYV?F/QY4Kd/H_:WGXB69.;CeL;>#KAV\A8fT>\2
gdWfGS+-9XN8TUNNcQ=F]<85cWP4NB/cGGW-#:)J9+(294^4@\CfDXdCGNM.;S?g
B/bS597@a1)-e_GEXUC+-^A=eGF_8I8>+QMBK(@b=X[ANfI)9f4Y]c-?EKfcEN1U
?C+F-42824A;CaX_J+AC]N93^ZFd,GYA,:_X0)?XX6(bK\N?WebOP9--_[g@D^-6
gJ1^/L+f\I)+)b(9-SG/.39DKJ,/38&d4P-5c^/SW@+46L2Q5[NV=NDM<R2bWO_A
SY#]@-9=[7DUA:f@/MQ@A1]_97BW5,R@0,E2Y:1QGY2V.RL_F5.Q:+E40,DaHY+Q
cR_#+70X4BF36?2J2X>848]f;K,?M=1<2Q(C&P>4]7e1L2O&J?MTbL2g7S;B>BDV
AY^@D)Va[O1\XQT^J:1-O_5,8[@&9Wcad97eCZX,5855LG+DFFLI1]b,[e09L@eb
-&NF5DN;Z&S2RM/V3,bBF2AOJ71,DdARME;Z(@(EeeEK:C3^]@F#29+HW:4+#B7[
EA>b\]YgO^+D-+9^+/GH3d:6S@GI:5MTEOWZ,\dL4GK/V#A@9)(<&LEfHR.VG^7>
ee#FZ=43?.\TY#/<0XDMgW^=;?ROL9KWIY>OM@KMV?&<\&6I__3,TeJ39OgfTFX@
[aGM-LVbXTGf>R7OM#@36g]WddS?6W2a,K^G0gQe2YFMB+,2/2.D5<E_CR2TROUY
.>:-a^S_;c=73X9XH8Q4NXf&/CAT&b>Vd#aGSQ35WK]F00Y+IWH&1EA=W6]NG54B
P4E\JJACB/L=#McTNH:HMJa@L#e84]]I1;\fZ]f-DWd/7L(NDFT](ETMeW)9H8_A
>fMfV15-)fC@@d57NZE?#J1QJcO_0DF+c9GKe:0D-/-?R8^R\0)]=3bRT_NHdK8G
/a=[&=7<)0&.)UVX36Vc,?._?+:Ra427YIBc9\&RR5N:4\=dO_Z@0=_]7-=B#cSB
NDQ/C=9/BPMc9(DS@QO^b<?<=YP336=/aG+>C9ZQW+D33_(U.d-?0PP<>W<O2_:3
,CC5=,QL45L=#1dV#8;).=eP3YTQ)EEBd35IYG\KSA7g6Ba&@5XH11dSdDDN/D,=
?,+0-#D@ZAd>.O^U4S08C-ITFHKIR3UNMWR-BM76<3Pd&QN6;LgAYI#Ya4MHN]Z4
9]e0?;Q<VJXfc&gO<c@2#T[9+FAR;Kg-N/E\a4(XE_-,=N6D/_]_[\GAbHFL8c;Y
-7.20#PPdE+?S=GWP\#RP,5^FUNbKW[ARS3OfK5:[IZ(&MQB-5HeKZSX8d)Z5eTA
,0E.S2]SS22R3/R/-1Z_VKe3G1__>=N<&?_fUF]_0\2D38()<1ZDN:EA.5+F9(QM
.:>f(WbF,b1I.L[]cNK<G/+OG8[K.1Qg]TG4]F6+K=g1f]De40)-F7_MBMbOGXUF
cM4bOB_LMDf+8SLR2N[c7^d>HD;a&W6;-7>Z#Z<Kc_Z-_S?QQ2KK,5Q\@_-Kd^3Y
H2RPWMdRYI9G21//<Bc]_cRX5Z&a;Rg&gABDJcN+.YYRUK(598\WEI=29+QEKS]7
3T?.O<&A/7H4-6D@:8:O?V0g7[eSeaO3./@SBGG1+Q+EM&+-a^#\UXBb)_QT]1g7
/>#H,5-DMP_4-.4](X>KH>27B\1>;P3.J]fcMVHP=16,F>,WaA>1.,\(02dCWX6F
DGIdXV(4I,_9;21E\,>=,R#EK;L@df;Cg+&bL3G^_<4J=RZ^adMa4SJ5)IdgWSJc
_(,A&7,?_+;EYZJKQ>L8]5E1U7.Ze9^d4dZ6\WO7A_X0BFLg\7aFV<ZeL<W=K]>M
1=T+/4Ve/1)^Dg9DD=;45.Tf7]c.gV;bCKX^K0D#ZgH56IFdLGa->Ne5&3>MW,T7
0^DPWVK(3QWd=/-3#46ZLB=9SVK44M^O1<7Pb83D(a>?JJ@?VfP\]gFA5OFNQcP<
gdE7gDT?aGYYTP,2ebL-->I.Z)CJd9#4POJ.;U.?K120_/VW\>9\_<f56YYI_a[O
XB#a(dNb?IC.9@NbOKf)8#N,0<ALO8,eH(O?e5/ZH\<GKKD1GECKS6Ra_12gPSQP
\\@H-8gNIJ3fS1GXJ<S50O>O4dA0<DWQV5#SJ.;BTRd190>S-+8ZLbT?8BbJH9IJ
GEf^[9ReOJg&aAC=<(;>=_J@-P)GRFW_I4)ANc^gVS-O(8Ec/)O[YA+?&9D(N,2<
3-Db;a4B?,KG6TY-g9SKUY-_2g1e,&3FO2>=&6LW8.U2]cJ2)MA7KG/T^&RGSAfJ
R)5.bX[:gc4?\>HHP(Y<:-W-?E(QSEA6f/+-AeV],Z2g#\C_Y)0W[(PM3^2>UcYO
PO@f3aXCQE>?O[=/LIOKH@2g&#DfZZ?e<(WCSbQbP.WQ2&ff&Vbd.^Wa0(G)[B]V
)@KIT<a/QW;R1DN<YMYcaeg/,#AA+R5a>=R45NIceNdeK2IbV?YcGQ=XFM1VU3RE
D1e3Y#QPAHB[T3g?CbE#bRR@08<WfG4,fdYR-UHdc-@/9;e[-<]g.d))?Wdg.1Rd
>79(.R3aZa;GPb<GL0c.]>94Dg6(J;+?3=GNYB.5VL3C\QWI:,._F\g\GY&KDg6U
YLDA\;/V)@]M</MJgdKPQ^VCZN9A=I68/gTLHKLY]0I,bId8(D876]41PSI)F<DI
>ZR;.Q#YCN?_2de5eL;OU65?;.6RbEOdQJ,g^/@Q-#YCeW+eL:F7cHVOELL]<2Pd
9+I_8](8;:PF3LH1KO@O]Ue_[I7E6H/05LV7fEfYA,<..ZeD)0eGM8c_A7;P7-OJ
(S0Y&L/ER+(RWVa0#Q]V@Yc)OIT0C\P-/EO>f,.[D\LKEY3>[C(EC@(\;]AR]eNE
#@[+W2bYgGIGHUSV.eTF+XZ]V>PW^g5b\.O,+++Z9PB(N_(cY)>-gTIDQg_PN[Ve
?LW2P\>@??HU:QFJ@JeW>0I,:fOd]e52?,aYL,VYS0I#CFJXfBM^.QEX^c+YW:a3
C^R#;5;efcKcI(WXECV^Gd2#H2YK65TQDRWX/F66c3bSbJ^VaT]cL9S3:.F\8C5C
=+1<)/3+S-TC#:(9,@,=\/OZI(IFF-+Z+:U<[-2.+,Ga?=H/707b:MZeHd_0aNR[
^ffNB=]._d@P6Ka&>U8@-A6?HLd)L&-6J\U<:\(5W=7beF4J2W&W3K6@;=4NKRKZ
S?9\gB0&MA),V0XLPX4@,8?Pf[0WG2V<gDcb1R7Q_G)H@)MRSC/L_[NcbNR&&4dc
eBPZaM&^F+]2SSRb:[A?R<bIF->;Y7&6]a#-2fITe31>C[(+Z6<:\,OA;EHJOR_e
3F_RFg]BC.8+O0SS8T@D;HKNfG@N+#096AH-_&O:V;./[S5R#7O@/Gf;:D704.a-
YY2f+)6^>KFb6PWG#R22F0KI><6dL;LF23MA9^S3V@-]S[]YJM0/@W)gQ03c0PJC
&.)]2-0SfVW@^4O@7>&AS-O+BeH8OA6I^)EOf./K,+>>a64dKGe>>BK36)e.(M1W
_\.I&^ZV8b;M&KeHdP4?K+NgDZWWeV9&ZSaE-&&PVS&<)X^=HB5R\aY6M^VXN^T1
aE5Bd[bF<R9_:,+71;IR=D-L;K(Q3Y;0],@Sd4)],E.d-fWMA2EAQCRV#[1@V?#U
12=OH]WEBQ_S^=OXOOHY6>4@0f;;PGbT:VE\CEdNe=423+T=PR<O+0[/eS),DIU2
;NR4<^.+=P[,JdF[&/E.]/3[WR4X@#VH@>I\(40aS]O4:RU7]>YSGe/.#0-S43\)
8F]f/3^QQQ)]^ZHg39N_PAC>AG_[WbS?DdU:)c_N)cSH#@?eH[d9+,]Y1[R8]56O
1JX1E)Y)LP,+59Y5K^d.d)C(36]:I0CD<Q\P4B:+C3[A,;RW;#d)_U>U9B0MU>YO
4GWgMa_\MD3KH.;_fHMb0L<_V8FfD71H&8d(/]dD8O4G9FEUN(+;>5D\NO^>GY.c
e]:,K#(&+>&Y5d8:4X4=RBXdLN1-gB-ZW^>=6:Jf^G+;8(+=0Eb<(AX;4a;B2MAL
5_dSLC4AFW8:H7J):^_3d7AC/&,S\MEX05R)),gQ\3f+;K3F=8AV?dNdK5GfT00S
6@CDAM2CdNQZHcg-J,UW>N=?1/ZMeI@b@(XFe>2GQ\LVLdbU>OLH-:De+^:OS/)^
T^CVC?G]?O=JF,7#.Qe)A30MLLI-d]?+.>:UX4(</A6R0@<2I\05SE^JQN\<ac<,
VL=E,/>U[B)Y(FcYa9WcP+?@85Ga)=Z8ZA&CO1K4M&@WEDS7Bd&2=QD6Aaf@D/E@
1Y,eKFKMP2TF:OSKF0RIHDD81JZ6;#,<W>MH[\,0gKRP]M=GaN@0T)QW656JORZX
L/MF\U/fOXbT2+Ocg>M3e;RGYHED-0eWY4f@+GLX9V6I8d29GgX1PXe6B1P]b6C#
23?DOQfAUK7V7DPW9&NcHA5PC(&D7VG,L3+1Bf.-TE^,I;2QRgPHNU#-Ma8P>T4e
1LGb?(U0:<XV;9BM\L0T_NSIZCT#@U]V#B=X^\7FK5U7+f4H0U-/6X(4#K<aa98.
B:5b-#CIBIH8Q1_UQg@Z1CdC#=M:O]#M&+I>.:4IR8agX2+N1F)#aBZM/IH6,/U4
Q\NK/-D80]2d<.c24QTAD7/@BSYeb>=9@8S:2P.d1dV/H:@5:5C?A;IVfP-FHDZL
98?DIgD_;E^NHaICSL3ccRG0b]AP>fINC2T10:IB4/]\<P&\ecaAY:=S,GW/1eFO
YWM6U?)D#+&TD_)1,7Ya5+1#[]c5_0/[?_@[HZ;M8UQU(dNV0GeW_;];)V85b]J[
6A.f2GBD0Y)<?:I<V579:6L>FK32^EJe3=f]HJSg<?eQU)M9=X88Y3HgAFILMf#@
&EDG]G-YbJSbJJS+PTaFQ.+D25+[UA5<<]>C\&?3+#@TTA=/^[A)/0^OM:LUN,4T
V1VWg:2J8J,\bW2HEM;(-V?O\NCdU/\7,[FO7DT+a\N]@-&O5J59^CZZXFA_X_H6
.0(DED],R_BL:YUgGObM.0e(6.#II)&=E.M;(&9O@>^QaL_S,U/8@J#)0&9>dLc,
1KcU:.&(@<9ZY,:N<D>APg7)JBL6YcfM^9:/L):Z(LQQYK=Q/.259@B.TeAbP)AY
SQA/<fL;#ecZMO@Q,4cfAgYM9,D@0BaB?b.,Te@AUG=A4M&DMB<16F\J=O.E8)J?
-cW7M>B9P7?DC+gM/(PFDe7<I-73gT1RWd[3^>]BXE8S-E8J&Y_a#E9aeHSMS_61
Je8G&^JL12+eT-Nf/eG1>;_e4V]O>Ce>T8@R,NQ-O-XLD>>71IV-GHF[(eC#;F-P
.;9QH\3PO-(XQF/MC#CB<2FQF<JI14R]A_db:8L?S?V3bLKbA4))(M\6>J>&&P;0
VF(>NN@6NCZMA/;E0=:SPQ_YPAO&,7cT=.&#b/;2->0.U.f5X@aaC<KWYN;LF.eR
K8GZb^[W074d>8-S.KeAFM;E@EZf_((644E<W0C]OP,+57X>NTP.H(c3^N3V+CN0
bF.C[:@I1>5YL(QQV-1TK43ATRb=\CQU:a;)O0;7@.F\ba)]WA7)S]&>df\V5>48
N:64VCg\1)X6<@@9P72fB(E4AXGd@5_#YG=OV2YcHTIU4Be<P7=?+c\SJGU_.M8D
;WIZL37O[bICP;P.4XDUa.9]8F)VcIY&ZTB.aa7ff/]OSd\dTESK1<c29(S7;Z)=
#:(0Z]AK#fR\6=S)=^I(Me@0\&(NT::YQ2/X9#F,c-D.OQ0OBI\.UB->)N#B9VF;
S(EaOa\,[Ha&B5KU04YF70@4RTJX74CeTSAefbb/9HE_BXfa__C_+ENU(a&TCGT_
N1g+Sb#E,AMER5F337Y_f8^4.KMSE;Z>FI(ZeS3;MO;e/QL5T?]I;f-MaWD\J5V;
FGF2WA1UafSZ@A4\HGZccWP[gdJY>)fA52Id@GS160;-O,8MP:6QAFXd(5-eH&7g
=f;?[)N/WL(F27\\Hf\_XNEJYPF/;0[<4ZO3B4F,R5O>2&P790<J<dU[=1^(GRMF
S-SE<53I2GT&7)aK10JCQV=8f;Yced)L:RZG<&W]^FMS<gf55#E(4(9X9fA@+:M>
Y-#Sg4W(=Rd&3BF;(?@=+2ZC_+3:fVVc8OA>3e8gTD@YN<R/?\+2G]>,@?4=a91C
1>3:EJ],XR;\0&[U+H/@S[1VZd:NA&_BD8Ra.c;@WC.P;\OY1LSecTB[R,F,7SUM
9>8N=M9^a^aH:23VM,S&YTcC)9MP]Z<N/>bY>#XOFUL?/>5SJ/SfeFJ#T[#IeLdX
:T9Q:BOXGV>_UHOQU;\^e#[>39X4\JY8acOd+ZGDGdKI43\+B9BMeOc\B6V?<f]=
KD=2Q9?ELJ7_^8/B1#KV5&IH&ebO>FQUg;_N,TeMNGMU#eTZFc7dH3&<MMUZ;SfB
2DVJ>]&3d&ffd1^aP_:]YLbdNN#I[BZ4J,U\M7@8cWP=,8aQ77PT,+F-9-bT@OfE
\);..L3Z6aX??0+7_,HN04G&4I<Y/NKS-V@Ce8eS)2NEUG+f8(MABRCR\<S:5XIR
C8Q4[9)-9O/bO[]B1((Eg;)0X]69@&V-C:.1:8HH5I6^\<b&0Y>,9.d[Hf27<41C
gg:.K+7GOY;[BW:>CdJVBV_cL844DTYH-_7[&5Q]2#@[eQ6W7gY(fe4^E14ddKMd
&JJ;gQ-f-e0aCdWEHUNOd\^4-SOV+8F:XPI7>cA\?OSF;/fW3&6[5]:1?[[M]aD&
9QUa?I;II4(<57;M+agS_-4b#XX6Q17_UG]DO5fO4=S;d5HgD6:=<>MLM6CDJX#1
dLNa2[^\B5Za4ZPOU_>D<;?RbV+G;>?(P9201Ib>=eXb#/)W.:W,6X&ON^-2<+^W
c8;d)aW#7+\3IC_Y@SY)7Y-:&Z3L@1:N97-M5C5REM61\-BGW?X44_YZa,<[=d-S
UC2/71(7+FK,9JY&1ETE.AI_/S:8?#_>#=\U>\/#M\GS.>@A6eI^AP<)TNeVL]de
/55:BY;LX)T8\=)6AQAI[bb]H(KUaN94.f1e/GFZ&[:V0^>0LgA(E;2EZPU?Z_^1
W2MP]@GQSRDTXe]e54&ZW^)\._),@5N&S[U-QCP&,:P/J&9F+L\,Q<T)bA)W@.5>
bI:&HY;e9\#DgVOQ/F3VLY>]=K_7L+b/gC]]Y1]AV;^[,_)T:&70Z\16KFJ(4LLX
=?N(FaRSeg(3UFcTaf.(@X;g0E[ROQ9/9gUE<TL:f)N[C;>)T6?0.T2?.3E@?;DR
D66Q7#Y8R[aPV]0DHUC.(>E(ZT^XT_:A?C@Hd+]1^5AB?NR-2_)G?8WC/09ZceOD
+K?24JO)D4IHS5U/cR-7e1Q^c^?3LJYU>&f0U9Y5[YYC)XR;Oc@MCH>H/8>4]_,#
J[?^CV&BP5F4(:DF4Od=ca1#LS[MR[+Ra@1GGAF\TN:X0AZT^NVC\7ER&;e:(/&8
34S(-.g1e-@&>3XX8baB=A8X^20]\K-d-;]A-[]W.-/L=5-@(<6/9TRP1Y7g08dL
4X-ND)[MUJcgT#/e]ZZc,.\XAHM6;dUOPd4=+\8,fOI_M<[0QdG:PV?VRG1&&PGF
V@J>WWAbHA8L8K9[gU3W(,1>)D5ON0E_KV.DZEQ6FI53eDM88]S9d_STU,=9VF\0
6:(--^..?,J>MdDLYeT[BX1aN+<A+0&VZLDF<Q/fH@cCI@=10:^JLCdF#ec>SJgV
F;/A4</E4>@C]M5b&HB\&INC&=E[OC[T0#eWZI>eAS@=/b8]KN[P]H7#Z)^4<2_O
-48XFQ+S[e[JVGa?HeM+gXABa1,VJg(,[Q<?70_>2X,=FE)F(^4NO(A\]8#V;88P
_T0dfRC;4f_G6Y#9VP5;QO/0L<VHbC/O<]1X7[L^bcR[X)1cd;_F?B0:G_@_8gH#
af_L?]M4BY;.IW\5XOPPVJ<]9BgC8E629<gMaB<B7N8/LU)Mc^#?_<=H0We_a:I0
MfS>)W/Y88\R,NSc+5g:,7H3&4YO-TN&Bf0AIG[]fM,TG3G^5Z;:0b_0eH3SJ_B4
CDA18dDNa\Ne9J2R><[V+(O+7(.Od9ER8C3DZ+E]e7@#_#fVQ9@,&[T/RGcg+/7T
T7a=MRTD>3IcCZP;BMa3EIUSTda/QX+6U[&NO&OK1,e]W/@95bHffF]Q&X4feRPI
-?W;B9[^<?Z0ZU90/@4<7T=#IZ@f&)SNJZd9:a1_<EW[GHMfBHCQ#@WYRH[Z+MXW
:_@1&dKbTWO.XT<]7[SCKN0DYH5E39QBe-c>Z_Ya-@/L@AAB_\NTQWZ0X,NH[BYJ
374V?e.,ZaI,LgD4)IO,@O&/3YUJ)Ff.&/GGT#R4dT@HEX&DPUUF9f70V:Q(1fD-
4T+9O0-N2[c3X/.MIX2>@HP:c.>F4&.CBBBDc(UVad/E3XUe90g84WfaaAX-1B.=
>H+_KD.MFFXb;E9Q0,R0GI#&Na)B<O,OIag<-F9]\ZL-S/CL[e<,&3>/N/<]G#G?
@D(UI3^gB2Wg6-0\UV+3_fgP1/cE^Y@ADPgeK1M@C?X[(J^?,R)W-RJWeec6>Z4d
\N=d\.W^aff?JRCL/G3NSW8:TZg+86B2E;?D4\\T3?7#?#c\N<J=DPH6+ZfD1bHN
H235C141ac33CRRLaCJa#Rd<161(EZCB-CY?LfHMFGI8:X\g5O)LE:Z8J7A&\V&c
\AF:+C+PZ^1d,7-F+UA7O8:aRYNZF<Y]YR_]QZAT;\X4Y]&8Wa?BOMe9;)=YNgML
#YHaJaLGaDGI2?:e&IT_HgNR>Y:XZG\Ua^;0VbYUa\TKU8M[=Cb-L^:M?H#_c[L.
,_F/)d)F1dH#5<cIM&-ZYL:dG_4/?U)gZfY&Td-]:b19U>K3(Q#:JZ55YYW>YMcX
W/bF<GRGPab:-^ABe/D9;W[=QOb\1>Y[1g88gGAAS]Z]M7>8)R<_e6IAM45@:dC3
I(:?AbJD809d733eV@L(FNQI>Z<\G_,MEbaR18Tg5D/<e9UW:[]T7JQ^)NFe;AF>
70//RfX@;Rf:W1CV_S]HIbdGYa\)Y.&-Vf>A>AN:5HJ2&9bA^&;3OJ;2Q-S[[f_L
KQ;/[:G_()9H-,OO5g5LcZF>,+HE3431\eXfdg>O\+PQe=)8]-8]+dea2SC045<5
K0Veb>c-1f:V\=Fg(KDY(4CM2Kgc-WZ#T]?:^3K@b^6#L-\5dfH06X?(@BAUK)<E
XT_gV#gaG#d_0Z_H,P,3E\VfJTMKE7GRXfRJN.ASeY+:cV;@EY>3,^Y=8A4G#CZQ
ZL53[TG+[;+<J15fX;9CQfLENc5E;HcDT,7ge0cgf(2U]G5(5Q,P;(^@7JLZ=L7R
?-Ga-48O<6HR(.8Wdc]B5&D(^0=2dM>R.S)#I9;J\-@>=_4?9ON3X/I\IV=^?0.7
d0)-Gg-e0&7MMGF:]<QJ5K6(F+/MZF)LL2=^:6;O/3<;0DGP8_4g+9bV?U;K0(:W
VW2_DQH+>4Se4AU.,T-f;O_PDL6;DH1eI-R;-;+7#9V<1L]8+,;E(65AcDf5Nc-=
c],fN@+=GRaSVPb8cb[=Q/JC7=_f8fFI+V\::)+^Z^ZRdKeCY;Zg-SFQb-7NSZ;e
Ge\4D69_])UBQ9CBZXfM;c@WS/8QgQ6-;558/TDUbOG@_]4S./+.))W8B=;,Y<RC
\3)K/Z0DI?7g^=dV^J0W&CBVGA:1R:\<5JL?DO)8FQbZTeX>LgP^9OBF[Ze,ZMYf
25UZ]UD27DF=1bD9>V>L8CSIFe43NGIP]>[=&GCA]TPaBX:[[-MVa^WMK&NII9E2
MFb295,ePYE.,K<,24TTYRab[aa,S7?IOSVYDYf_<K0D,YQ>P&/-aYP37#gR.G#K
\J-LUB8:eC-ff2^EN[)fZ4U7YM,GA0C6>EOFQ7f6_(g1UWH\&EJSH\.]@NO]2O&L
[L1=/EA3)5=Mb+QD>V8bACQY#-(I4UCT9;ONW@[CB&@\L:Y4[c\UTF(cJbBD&W\b
5NLgdb@4/WQYZN/T[3\3M+C1#bJ42TGTYGf918XYO=S/)=\=7^^:VV:=e5.C=6WC
cdXbLC]\#COVg<1SW:_R\J31E\EIbEGKHab+N1D2>#15KT[7BX<<8e:fV^<ST-cC
C<d9TZ(VPd8Xd5X_bA+9\eP>9<#W)bd<7W;eG_d9+_N1:=S;aSP,>J)CNUJ+<Dac
X.VZb9DTe08DOf7GV8?VYVRMX4BeF(Uf+5c2LGQDg5e5fL:ZAFN24bP)?8(T]WSS
64G\NcNa#N.F,?-4_J^-(Zb_W<9BANA+NFKLWY)L8+g[#F9CP6X@(YYd56K/_0ea
T/Y+Ba(dGb@+(Ba=X.;T/W(LQNE,0-XC[NEf&f4RE+O0MS^[DF-:Uc-D/W7&SfND
92@\&Gf49/-KZA-2JJ(Y_W8d0,)JF>8)N1C;QcLJH7VUV/]&6U7Z&[3L7BA65++K
V#Y>HL:LgDXIWbE.e)IU,QN4D^+>?&F862>U_<022T&gg(Kb/A;-D]5^6BT_:IS-
&eeRIO3c3-.19Wf(8:=4?UUJOI^9>#ZRRBWYF+Q1Cf)@e.-]CS+dI4SOXaOSQ,#V
#@8?g]1>:YZ\9\PFT?.&Cf?1.Ie+O^]\2RSA<UXJM/N]Z&BM_[8R9/R\\=COYTdJ
)GfD8IIFW/3#5c+=UNO#JC\dGX@).H4HPVR/U>&c@Y@_\N.#BZ.?BfWJ^[DCJ187
54a^B31;Udb1K-U-(K.;QHW=fb\VVOW04Hf82)F2N99X4Wb;+(eSLd>b):7\KgcX
CZd+>ZV#@QIGVTN6((@_CYUN#P#0AQSS&[\@/@[<aHHaM;22URO.fcTa_4.LU)#e
d@>([cD#a@,(KJeg31HaI^4d(G2U?64A03g]L\0F7STA-8FG&A7J@NF5U#()0\S&
K([-3Mbf(fN>H_eD)^@0dRAb?N[G8\.=/?Y1)0)E1@Y&VGa#+Y2T4/WA:D,MaT0.
I&6[g>CMS+eNCRg&#.VW8.+>->?H#&2B>#F(>.7?;,\2O#8>8Zd^XEaFDDEF;dSJ
JJ1FHVZD5MQ:f7.N:B_;f;1Ac>b6M[E]8g)_0A,H_2I-.;&ERdgcL)12;EJZ4Q_b
^.OT\5>FQP7D8KdCU^AR:46>Tg#Me2@(J;ZQZYDDf3gQ0\Hb#-)aXd(=09.<gT80
)^S92D(O,^5dZQ1bgND>,@GbG_<)3CMfUK/J[bEHF.C4G_STFE]>CWSK4&/O-DGa
>7PM[>[>XUg^K]TXEBDdDI(U/WUQ<fU#E4>@I@ID0>3-QKR?4BZdg^AMD\5e22=G
2:,c0:N]JA6f7(/1b>;Zgff1?d2/Y5c=_PZa6^^F);CH2:5+3GHc@WV7g.+M<3bB
c/&Q<7C(@;V5d2]XY3_S/@G+E4W=dFWK:ge(C.S>JSd[E5,NICaXa:;NKORU\\J>
2G/>HT.)b\;/[:<g;3E@V^U4W&WX&N(BdUI3+[>O\#P;J;P;6V\HN&ee=O5PKU\P
IeE&aZ9A:S?WIM7L)&?K)=MSeLKORX4AQL8;;@N+adR)M0W]SRf@X7.<K6[:]KIE
O3[C8I[Nd9>dU,GWP<U(@>MK1/+(_F\K-[>-?c8a0_E=3=;TA_T7/=TD-0S3V4T;
F1H^5.N2NL,gXC@#Bg0UG23CX.;d[;N59[M\dWDeQU)(W+6#HU_7<CKKO&Q]PaR-
GG(6N/GX-2GM#We@)f5f[H=/I<Y1T_.FfU;MZ57D[)IAG92/K2I,C>D;-@LbBgLF
Z1CXRc_4>\/L2N^^a.YXMV(XH6?HDB9e,5/+1:Db^JPQ@#(2.@0gG\eH0L@IAR1O
2R8BR#A3:9fSD70&fS:E]>@FEK32cRTL-TINJXS/;/8ZOM\-Ue&MQF_df<VBEJ>6
UWYgA1aRP[7eY5X31a=;Xg;^FgS26QV[DdQP5L<)5B<Kc.XUC;6=9QS(NQ.GRSfK
C92QOUG;+D(0;U5D^2cA+AeV+,F?48cPTgM/A^KND()Vg9>-<D@cU@f\7[GKK;P7
3O8gBXe@K)OEO7e@F[a=PC6c+Xd0QLbIcI1+MKB]D3(e9_JgRD6<YHI<(SS0Q6:@
;;V8(<HAO3=_PG:V1/BK-I3a?L0LaAM0HPA,]UWf_gPg1/[96Q_>fXf)CfI+20LO
O@23[88(M,R<7;[gPM2SMZUS#F(MEN8WZ.K81bc@:gI9IQ0@S4d2^:Y]TEMB>SP#
2VE]aE\fe>CB)JP3G0M\IM)A4(16\;J]?@]3+W>?ZDW9RQJa-0BIT+:&U?P[+V5C
Q8DEb7KQT_7eR>7^O30[BX<-_TMaBQ@+8J&,:.0=d,?D(bgRT9TGS]<e3Zba.5-^
Z:.[c>8QK^G6;_.4;\<BAGE+#N+4)94E1C?_)PN.F3JPe94T(7)Y(]e3bI_?V7IR
?+Z]8fHGMaDbZ0VYS^6]]<I_P0,F4HKg#)8R@eF(N1bFLBD<X<CgZe^XH[Y3;N\.
&=9NL=<5,>>eG\J+g+C:[7ABfM25KbEdeDeM3^ZC<2N4GNOUE\:/QUL[[UJ7?+W8
cdY/YZZ+N4595I&>;,NO)VD-X\G>aOD^d)U2^_gS;^3WLZD^RKcBH4a9fG,5C?@(
fa@V?/cU0R.OC:J6?A@gMO8DE+-?6R++MAa4c>ZE&eR_UHaE]T5faSQXNd<Q1J_E
##E@eJ>7KEEcg6-dKa4^[4EI6GM#KR=Q^KK3f,>[9AF#gSbXa,GE(c^CR@H5-)/D
IP_=<L5\#NY6dEMePP[Id;#]F:eFbQCPG2<Q^9(;O:S>+bEHAda92_R/9VP??,-d
ecc(@A6/RM4Nf6N1VS>FH(M8WX[Y?&c>SD,/BN)A6/O)F)@?AJg@-/eG>#<0+NY-
[EG0)_]3e:CQ3@8P#>R0AH2C#:+9^JA-5f;@-eYQPXEPFJ.<TKQIMe4:<;TXK23;
4eB/I=(99DC<ZMH>L26#eU[[5EY&db4^/PZO-VMMJ=])G,>b&([VR0P63)FV/-B=
CIaTBK.;8Y3>W))PM^)dI5+MHTg5>[Fcg@D:Q-0XB+K9^5&[H(e2HZUfaT2a@+PU
PbBL<-^FO[2BU632NE+U0O:^BJdK<M7)T/eXbB^GH<Idg+OZTQ9Sada#@\V.@bF5
8>L.2:>RKG+]J#L?-,KJHgH&<(O>]5&AZ0S=M>?-9B?WJYB#DKLOMJ-02GF&S-Va
H>@?(.Ad0LFVS?9MFdS#_][F,E^LVE)O2d390F_#C10FYI[N0d=:PQPD8PF\Q^?B
JAO=J:c/b2ULg(A-O-eX&S7GU2S063e7?AbS;\)=-/7/?8=F.&[H>W=X3\Cb-_DD
.>PKNXJR1I;ef>E\[I7WbO0Ng9P[UIKN=,L01/4cXF-3^L,R:0.[W-XCF#5/=>]P
bF0CP-Da-9WTYRT-_ZE_LLd/+8RRAP3A)4&^>9VMaD3EGVBSE1Uc<2(QUR,CTH;.
\(.f(W--(GT<=cN^Z:9L]McFeN.G,A9#BCI]S>J,V<2PO[-[Rd7L-faIMP1g?R^D
NBeQI-5L9)SW#D]9+S#&N6J4K_;3@J/&>;_N-_SR]+I2COd_.H8_74+bQ1_Y,e.a
ALBQW5/be;OF4b5M&OO?g1YS(LE.Wc9aa/DV0//?aW8[3ZJ8QE]WP-+?5Y=fFG)>
6be[Yb#F/.-##+F&S8cF2-fI@)=9N4g,9<O8AE,Q?g;/;;cQ42(08;8O[B/@E)TA
;0-(Wd1MZ=,@?^-<3CI_J2.+g--RI?6NJ^Xa47AIBaPaQO730E3FZB@9>WI>7,^H
,R;2O[P@H(=T(EgJdf#8H;fMS4[6RI,#&X9(cPJ)5caggd=7,MD:cgL;LVdSY4>=
e&+G5gbWJ_H;;K,(X?-KAHWDK&JbdQ(R49HDFS\QD(_PO_e-gf,L-HC1V;M=#TTF
8:,L=Z-_63S1E0NR,M4WO_b7Y]_^V]d6S<SOZb2M.-4KR))8KK<cY0\M[1WY9?9:
:?Z(bE3_ZGgW9Y-Y>;=b1^5<g/YV6@;1ERQJ5VaI?B1MRK==61L\RFeX=K/a05Nb
6X5GIE8,;7)OJ(Dg,e&dIb=#f1H@+GCN1AEZG--6-ZeT3#EB&b+I(WE#RO&(:HW,
#a.1@FQ1@Z9cSdZcTXda8L7&?;BV)]I9.d4KcB)L@#]eEORda?U1]^#S@^9d)R2K
<.;+;H3K425F1^WZa@4f>KV8Z)We\QS]2YYX]AUAB+6X5KeAZ]/._WF7/+c(<b9>
C<5LTNDPCa@P,\c<YCLgfD<3)+6^3)@ECZGDR]-\W:gY9\U?bVWfD+=BP#a7.g#:
NP,Pf]&M]6>15@UG,2#?9Da);8dBI<[T?ffg1e,9#/__1)L:T:4&BDfPT\.NN5/J
4@E1IUYVQ=a1=25Zb1&bOIL4NIR@[d95;fOV/d>ACCM:D/#6cNXPf:4D1R1R;+&B
LeKN_c5]+;K<5(_[/PQ9F<^_f:D/KMW?@fK#Q503P[FX(@)P>-6J;,+4&QQ(XUE9
/YUL6U<X--(L+NAYS,YI0aW(?@J(;QL>,]_8;3Zb,?ATX.T:\gH\H?JX:?TId-\^
;-:A0JgC?(R<KDa)7b..QNQ\b+e_&K4O34e_CdXXXN3Q_P/JD0W:c2>dNMI,C=[@
T(d46VW[cSc=F7_DY..da=1g0,&V93M7:1aP[VFS;d->:MA,]WT?XfQ9)E;D:#3>
A:=Z(9g[d81LLGA(1-FG7]B5FbWL8O>b4]YV0,B_?P(d-GOAC8YIbQ0NA_ZPYa\M
gVSUJ3H:J;TG#]_0CZY.19c^=2+dOWEG:CFAe8cYRW[7b.5Ke85=;,gY<SVRCM]X
CDAe@C9e+dLc+Pca6&?->L\Q\T#8,D7]Wcd>33#aQ877P^>V@XLbW6Oc/R3[=d-/
&B7]E6&VgK\G<4G(WHD[SXLV?I&K:[2O?$
`endprotected
      

`protected
gCL2KFU+[Q@]36SDKKMKU&^DGFAcV19OH?Y,LJ:.SJ2@.OPG:EW?4)/CF1QfVSR]
ZdO;H=EE/6C].$
`endprotected

//vcs_lic_vip_protect
  `protected
,U[\Y]JH:.J8+U2J1ZT7J75SQO&M6?VS2Z^=^XJ(2MLa&g[.O<dL((g4T-X_C<(&
B-V6f>]OK(H@Pg):-CI-IS,M)F2J6=G]0(/K\.ObZ;=IA)A6-M-F]ef>7?(dIOM8
YHVSZ/AJ0L+XFY9eaZ>I>K7#Y2FXYDc[^Q+\dU<HZ+NTDC0GCZFMR;3Oe.9^D@AG
J8=:)ROe7gG>4[SWbcWS-H0E,cRZ)Ie>EZ/R.c]69D?>gZ?_C(I-c7Y\SNe/2HdM
FAJ(QFVf7K3BF4Q10E?VDd61RRN.[56CFBM-K2V6?MK1gL]X(_fB.5-.>\+P&9gS
,YBSPPA&g(Y+OZ0f5IA#M3@#L?FT.KHMO=BB)LD6[>8T_M8IOK7^VZ.g/e.[GbQ>
P\gV9#T90fLTKe>^5Bc4E200:CVTRL\VBB1Y[82/b@Q46_K1V@E^O;TBFA6H#4U=
F4Q?P:;31K?AI6L59O;+BabJ?YAe]<A3PU<IAAU7+4B8&e=<P,R4YaUf6L<1U_))
V5BOU&g8WO5N?,K+[2b]3c,]KS49=Ke?LFT?3Z0,[2c)JgcYM#ZFJI6d[c51\L13
MMN4KZBP@URNF_a[ISBU9(\5bUT6OJ:L;;6MQH#)F^\7W8#+<?(c?=+2)OR\cMK5
HafU<N+T6N(-f2HB9P@L:Y&?#GA7S4g)7]4I0W7_WT_PB++[SVb:Q_@(ZXWPB[7b
,@-+26/+V0eC4OD@6]8[Y3W)M5ORK:KdDCSC5cfI_\)0-5/17\4SQX[b6IAS7eU5
3D#OG=Oa-[3F,<-8YD7=f\[/2GRRH8J8:cL?Y200729bH.6>32KNZ_<LB-8I]XCM
g@:J8E/AEdSN^^)[P\AA=ZDF0@QI@?D^<T4JB2YQ>=<@LeQ<a)]c#4WE9\6TGQ@P
312BKQX8_TR2=IgeI#7ZHR+(=1N?UVXc]DX&EeHK&Wc4F)C7HT[KH=TcE00)+^Y\
F2_KG96D/.ZB-L?06&c@f7+)W3U&W4XKHT=C570;SBJ6]7=O/&c+eL/GPE)6N1cH
/Z&8]fS-d;?\X<>SJSJCEXQ3PYUYG^PWZO8B<Z>^T38Y\2@7DQ;2-IP:eR4--,WY
@a]77S5f)G)/;?H7/=]2R)KN/436F<1\V8-MaM3/&G@0LU1-LBb1EUd4N>=L924=
>Ef8-[4,Qc4LI<f9X/^K;HbMa-])X0704&?0UNLdb:5:.@[C+,K@HJ@-f1O/<>)V
^1#?ZSd&^72d1J-f89D-(Q+[&U14)KMTBY:C#&8G5#gP,91,Y#T^S;&IS(4G5[71
R4@_+TX7ASXMZV.Aa))F20Y7L98O(7cBQ,T4aK9AXAT0(+)?:<f]G50A64Ha&5-E
7c@0YEbUa#FYa=bCHfSVaOFJd<7Q2[NT[TK3ORb>LN_Eg#;f8<FS@9);I6;gb^bf
4TCXK>0H:RL&@.dWQNF>G#-[(gR^.ZXBBGa0a2Z_77WUTP7LB,g=.B4_.[F&X7&^
Gf&+3Q-I7e,3&H9FN2_(U&)QGU45,/R^._[F]O([]Teg?ISRH10A3L+g?QYOV9VM
(QMZIUVJK/.bL/^G01UV4\6CRP#XL6FS=Xb0-+a^@6LbEVL6^2(Yg=J6J1B[D>.;
,NF1\XF=1X@DBOUa[/\4eR:3FME-E_gJF3/0O5ba.c)2)7E5)X#PG+&&8(B+,Ea#
]B@b>dPDO-=[9)D_Q(,1<08ZIHHXPe0]6/>D05-e3:A0IZgZ.H>4IGN<8#.\+ACe
cE/FB+CGE7JdF;]0a;9N;E=ge<E&/fV4ZN<\/F]K4JR3,ER47bF&ZV_Ng0(7VY:D
598WgM0eE-5#S&I]LE>^<L+e5T=#\a8I@MPJPXQW.JMA#H=WeGf@A_Y(6_b([-;f
NW,>9bXG-a5T#dLWT7>LT=92L;Q95(H.D;0B-IdHaUHGE1PQ/WH7M@^U72.6f04<
4f\Ac[GNSC4NB/#7B0CH0-W)13J-0UMNJ+0J;AbUZM>DcKPB_\8_)<L>C@JBVARL
;Y>LZLfGYT7\S1#Z5+;c&3148=E>,aLAOG,bT,VN3<+2P1aGgZV5ZV>X<ffNdFQC
UdIH-(?]OQR0V/3-9aLSQT3?g]DMfAH;#b#JbIS#X#/60be&5bP>e8I,6:ABRGSD
XA6AW+Zb+N,B]NY622eYVPT(a3FdeZ..-I28<+5RDFE>=_;E_.c2a[LKGS\2^bg>
/5D>/d7NT^gWgIRgVY?I<B1.\eL5;_&Na+\XeTJUVM>\@P@6.FS5#MIT^DD@9,:F
+H:2/4fT.;C>Rg@]BH-LHG;/6[KdCT=WBOI(L-RB+3;9I[dG0_A)#7P@Zg1-]PKc
D_f(5bVPS)P<.eZ-2X-a,a9J@g:+R/N_Z<@(#N1EeL/eH,CWU_7^KfF]/bI[0ba?
3B1_:fPPZ)CYdaH+D+IgWAB<+Gc1\b]:ER+c109:??9L7<D7_,S8Mb542#0P-8[+
.bg[TKUCf+]#HE6Vb5A:+=A1JLQUC33/7A3LGS&gK>\b[+5d:#C39g[6&1Oc9VOD
MG><+N]H17VT_JF@=,Ad):cF>+3bW840,EM5YP-H]/DL>cRdgK?Bg7VR_,X0#[GA
IgSD#Jd/T:8#cIDLN>0]_N4@O?MD0S/C0;#QV2cOV-L(/e(/.[BVCDJ7=R16HfL)
Cb^G#2^b2.(>WO3N^V(QBR.342aH9C<\GB79AN,:7=L;A?,GZ6c;V3]Dc7]P,0AJ
T2ZH(]XQV0\RK?2f[7>S<.&g.&XeRH4>J/)6I@-,[/]]>(e;&<I\JW2J,)4OTf^/
&f^9J)JL\\-ZgCY-SAY?&aP<M,3d7Gf)@EVHQ5/3CS&b+YO;.^c##4^<&2]a:QQY
;PG4],d(Z?9B6Bc6c@B72Y]CGWC9+U#eWB;99a[fR2bfUd4Y:GeB#JUE+d,Le)WS
bceg;RZ):K80172G.O2LBOE=7Y0G3E8(XBIM4J-;?QXBL)We)WdR(aD2YN0S4Gg9
,F8G:SL#7S]Z@gV[63;&aH3SBWcL:+?UEJ4]K&WDN4NO]&?bQEPS6?-,D4\R,DUY
8M]M[[TM#-A6bGFd#+A9[NHg9KI2gTQ\?C4#+_LC0CWZ,KH?ccXO5+_?4P8M@N@G
;38bBAG540L6;MObB)Afg93R7)86[(-IF/a-WcbGI3Z(Qfa?,V2#&bO;-[F_8>CI
0/(V@@]P.LRgY=ZR#>d<C?HcG,\:fb(cS5DN=62E4aQe_,<e,:.^Ee>Za>KFa#Ub
0J)&&-D@;]-_P+P34K3TUBS?)YVT^f<5LQfD67[/QS3,L5N5OA@6C202A-f,#S)?
)FS=B5.0(TZR(R][[NddI(P6:Z=?S<#9.HZS>]aYTSJQJG_2XC/;b:&M8DM3-.Y8
[0OJfAA=ZA\5X0-2JgLa75ELIfAKa@:B>/a^9&6bJdf))2f2K9V-e<,_B[94[6+^
YR7K-f<3EFR5.eH@>Ib6\.bQgF#Tdde+Z^67cNRIU(FXB\SG+;6AcRPHa3)Uegfe
FWY8\ZS\ZVI:70H-bgCf,Yb:E8ag75>1#FPe:ELJa7W4e_=;&,4>KWg2ISV)PXS@
dYP2?V#8FA(Ve-]Sb<A_ANHT1DQVL^gSB@C7ORe,5(]dEY^7X0\70Dbg3ZQ8gF?A
\.c:G-)Ff63)9SEO8EaINCXXb@_C/2\2,2>[dZ/RFQJb:N;4\^#Bg3M7A:7g0U?T
<?-]W;]6X3_XXNd^:SZ>-I>,8SC]eMWW3BVCGW:3a>6AR2;M4LJT0>eJ0NbD[:\K
0LeL7S6?0e\LAFFI<#\+UfI[\W(a;Yd0cD=^Ae+AKY,PZ4MBOQ^RPTdKDdR>de5I
C@?MEG_&O<GYMNFCFDV21YTb)aMgGN?)YK)IdX=/(_U3<:7>,dAB=K@)KJ&@31Ed
29B+/25510,DNcY&<NB\-dIUa,HTaCb&:c,e3S(=.>bXOU9K,UMc@76--=fFf>8@
g_+L8/#U9(?gFF\PG[a:;V#<LN,GGLBEaU=UO=(/5UT,Z1N.LKXOSW0ECcJT0a44
<J?TZQT9M_b49eC<_10[QcfDYZ+&R?;&^b@C+RJ5ZO,a]X\=5_&H[W^[+b4O/#U<
0YbO#7fZY8]RUME<6208a6MD6G.\=BU/W+bRR,R3F=PWg_9V11?-O@H(M^b07Z/0
La01S#EW]YRDB0?5fZBD.fg]GHGRZXE8,-.^W_f=;f-c9cTRf9JSTQ/PEf/?.;W^
NHK?9gOS&_Y/H-6[dEaIfH1,@G\\S95fB<Ncb<#+=ab8g7A;VSGfDeA(1J_ObCRJ
YL<(K/,^3KYGGW:B)9O:N^3]=,]B7>+E4(4dgH>5FKCJd;dZK0C@Af4//HTTKUP5
7Lc2O&b7-X=TbBgUd/]1]=8ZYI.XYC,[-+^T4:ZS3XLCWS:Pf1#)2]L2]BD,/JII
\E-@DD0bO]AZF?deY1NW3V,P2,FFL)2IT5BJ3a@cI.O15MaX1We70_:=f#a[N-Td
aE-QccM>2WeQ626<P>BbO-(M/V;c[I-MZcTG&>^8N#TN^AU#O&W+WWNSQOXET]39
0NS3H:25gI+V5__A;f#Qc#b0,?ECU5\;8SVYcWCf4W+4Ce7aW((g3T.)Z7C0S:B6
]+V/bH5M]BR-IPQKe9<=\C]7UDW]C.DXAb-_>;\D][09bPI6=?aM;J7_)VE&T(?T
0RS.-4R##e7])TAN1[K-DQ#\K&HQ=RH.&0a_3,Gg,Q=P:Hb<5L:#gd.UeDc=;Bc)
VT:9ae(,6W::\,Fc.LdRZYPQ,_f4IIg5HbD8)SO)1VX:.K^LA2>eU=91.;O\CC.8
X,P.dT28APF4:D;(:56B(AB5=MWEcYfa@0A-CMKLQ>FV2LE&EdX7gJBfVgF?X5:K
903XFP+a=],Q;Y=0>=<gOLV&\-#5+4^Jf?@dY6>I3<\?WbV]5X68HeL:fM+GB)Z3
12&8e6MA)L.ZVP^(HZ_:b,@LIOB)F1#)J1MfW>H;&5a_bgZd_0XPVH+\c:5VEJR5
@P]J81MH]>T\OVV:16Y-;V](B\:ESQ@?6YP6<?VN4J?e3TJd^a<YD#D>G&),SMdC
ePd+FB(_AaKa#:]/YH>]#&&?KQ;PQ?Qfb@\D@XH@dPTaLa/BKbREC3AE<Hf7?41H
BWA7D=\5X&UT7><3,RJEe?bX=2<SBSd@CUeZ/LaAC<#CE;,e0B=Ae]6M.+^@d2C3
IU+Y(NX,)Ud.[2fc7:R,00\)bI5C-TA@U:/EbZW0RPdfMY8e7\?EK/9H,7BcOHfY
6C1D]P7C@O/[0#+HVY0/3&405ECgS,c:e81>@9/@U\eaXH:/fX[0[\3(Z>^WHG@e
CGDW8_D)O@SP^+2cBHXcdbY2;9Oa>?:f6GUe?@NE<89@fOXA]0_U0Z?+F[9F0;6M
6-M/55JQ>?;BZRWJMZL]0<MU:[G8JX,DX^H#MbceOR14(7W3JJEIC3#2Q<&Y#FfT
I=EPOW/N<bNFgE@E;/>7/56M:6&DN9cd8BDNdI+Y02.LR&Q4VBR2F@Vb<@/LM9/(
.Pfg76S+#R&HZHO7NG][Ka(T+0?^^;R&H9g;^/MT1,-Q,Q_,b;7GYYDNgL]J@W(Z
[A;TPXJHIL4cV56A,X?@cI3=R<J@/YQNBdKYT=Ia@g8:EUcS-KKIJP<S6Df7I(E\
6UJeUT.a=d^QE+e,U@M4FX^0(MP_W/HdI&O0.[B]/G/JZ?R];c-Y):;16c=,H&OF
M4Ed0PZTVcM&Xcec:[LQ1RPJdA&f[M[^N_TTD^9PMVcQ5R65JeKfCXZUQOZVL9bV
UL2TS_.-_4(S\)QMM51^ba48+EQa2gK@B)&ccV.1\@0SYU_L0b2AR\L>LO.D&E&(
d-3OUD>/_:I3bPfGNEf[QHc3#H5Ne5Q/[8NC@MI,(37T@.J(3W7]I&2=Rgb9N/Xd
RUMC76d06(PQ(_9DC\cQ.aOaTdPBW7eD#CHCEXP)\eVcEcY@M4Wc<Fc=27>)@Q=O
=VZ.RQL2Bfd?<4])Y50R201Y]11dYGP?cX_H,]TB9.Vb2J4VRI^M>0)R;NTUE&Te
IMWb0eYXJg0Y9JB-S3C;B[IHXU,V8ee@),1H<8BCde#=aRWFT9,B-R6a+9>#d&dS
Z;&Y\FV59KWI1.-_+AQ[;X6f9\CcFNeCX/a.b0S>0#AA64D34;N#88-7,&9?Qd25
)\<&dSML6^8?XXN+;KQ9DTa,aJ,7L,_YeS8VOXf<#Z@==[VMHY8/Ree0E2>;U?P,
;Oa1>J6<E24ZR-9^U@8FFL82e(R?43<<,RS<^DBGU[Y^+_OXc5D2D<&Ia(>c<2H:
HDA63J51T9BbE,=\_RLQ@cdD?VC;UXPW8VFETDf)e0.?D,B&NA\^GN//=EF&F1aU
DgO_d;MAgP:B2F466,PB2<(Z&RO1EZ[&Z>0gF1Mc2O<#UR\A62;)[Q^<FPaTU^1X
7KXX/D2,aY3&BVf)X0fSZD4@J4fUN=K4]bd^<\7G)@+G3@C&b6g1?Y,FBgP4<X)\
A8bS[\M-05GG;:JD.;0cS>,OeWUDC#D[/eMWK\#9:+&/Y9IS1&X8Z@ZFNJNB92W[
MA#gI[2C27fD5P5M-#+<?R<DgE;@&#gUg+bEHHAN4-615.?>@&W(#>OF@Oc01-cT
cg=g&@B0JBMWD3R&Z/\.Zaa/I,M(<ae-]#KO;DHL7=D2KdbQfV,.;)VZBGG:DA<A
T;IDBQ8>fADW-$
`endprotected
  
`protected
>D7.,FK1Y9SQ-KG2HJ,Z@R^EL+1W7,RUU6WE]-+E40.[H\c8OSFL,)<5LZ^8]LG.
VU^/G_PR-a,Q.$
`endprotected

//vcs_lic_vip_protect
  `protected
G^R@>H8=Sd@O@aaRe=)RB@55H@5f\.\:@;N/YJ2N,P@H\.TU:Xe?7(4CJeID,OaR
G4=9X55R9>BZF.Z<Oe)>#>ZVI?9@aL9D7^d_+>2dMKI^JBDDPg0)DUFdJ([dDD6=
B1F_@\2E&Zbe#JE3QZ;=5I.THF[G^FL+I3=E.9^\<9C3]?2:B/ffUVKJ2(8MH(8b
E_+2c\\=e]I[E3J^JdcF@I]5S6GO8dZOAYb2;#cY06Cf?X.X05A^f-ZRBTA^W\FS
XA,-17C3?;(d,/HP)W_)1AIE<M>N+MdN_T-+#KTT0;XERZGEg\GbGf<<_N_27aC0
@6A#^>W@-FOb9MUPH[<SQ2\[ML?QL@@G=Oe/BQ[<LEJFV84OVFE(;S=Jc--EKP0A
-YJ51;NDGSUW+c@>4NN[55C)+,>T3P9eZ<NFS4:#):ST1W@2/\_Y<BR]V.[]Hb:)
\,:_J2c3-A#BJeUE_,LW?Z_ZT>6,78JgE=I@8XE>?VO5:?M-+WR@0?.VDC#A;&[6
b0gBN61\BgCZZ:T.BA[?OSL,&HfK?Vff2R8bOFR-;;:,@_UC6(F>0aN-@&.76#BO
4ggP/Y?BfaW?A?Je]/#47D.2bAfK6,gRX[=(4(R<,dCLNeNd8NK5#J_Tb:3-eV?T
AePEAV9,_&F>=;a;a4,bPG-_gXW@.LHL&1R?5O+/\/+SP+GEF,:eMJ1)gX(Df,KF
U<8]3SSbPK7@B+YYTR\0VH(Y;/?Y3@EZPRWeC)GGd@XJ3,F^?501bJ9f-@f/[AJZ
E>FB&]b(L1b+:DF5A)=&6_B;=N2eEc0K/<+N8Bf:24W.YQ[SZd_B9g8dEYf4RP?[
_Q)#ZX-]g[YgI5A[QHQCUS76PQKP-Uf7+ZX)[g^acXg>?a2d+.K,T?:c/c+LIPS6
<&9S9;?Q(W&71Y]+c&A\Pg4V4JQIf?#B<5GII=,AXTY.GdK<PA^AE2.f+a_N3-eI
4A,_d)VQGKXVBbDR1fQ\P)4V4$
`endprotected
  
`protected
6QUULLa@cd38I05ACU\I6]QA[J@S2,S_eFP@Ac694M;2g;A1E<RD3)aURTMJ,5B4
@J_:V<5>?(+8.$
`endprotected

//vcs_lic_vip_protect
  `protected
1^cO(\PZTF+]KGA+XWe,:8?[11CM>RVEA@A+BaNEL,/[dP+E0(Z:/(&8BRX5ZU)L
)RK:BSabEFK:Re(8+-7V_IQF?UcOB@C&#V,2_D^<U@SEJ4F7dQ@:cY7T1]4:1^G(
<g\(?aZL,&I]DW2d>K>c(fO0J;86#?N-GL9#@7>E:Ie1K7MI<dP3U_EOPP\M^ce\
Q<ICHW+QOP.)1ZJ-BE@:2?2ec[_C;?1[(AMH2J9[1J@BQ0fdX<NR4]A-3Xe>O(9U
^NPG]PMb>VXVTK.LS?K5W.2GP1YFegQZ)ecN5fUb5VI2=B>aC<gRAYG8VLHHFUR9
.B[1A(ZH;-BeKDCbMI[\;SBV,Zc7-QF\eb#D)>)1]Vc?CTTR0\G?NFb\Zdg<(^c=
=R^28C9>?6C(<gRR.?C\e,L2cMUf&a\++9+?\>/Oe2=UNfW2P?.\-cVXG3>MAL=&
OgQIN2Da>ELWVZ&LPPH>dFHWH9G+f16Ccf+TC._7#e_4AVP[RfGIUgd6]e8Je2/c
-QVG6PgQ7@1@a(SeO/5d]FT#PRT<R1-(cD=C8)ZQa9E7:4QaEbOPP/E>gHcEUI3f
(O2Q=PPZYa5>a8EB16X?c19-T=bK1+H(M:)L7&b>:TSSHVVC:b<9UABOE5Ha<6J9
2Q\5d<gP6-5(9RH9(gRg<#BD0B#WUf^Y@&]:[A:58#RZ[@CXXMO=Od^I1UX+<75B
_\_.1_GS2@>4\6P3N:bNTZ6Z?Y1J.N>O;Q5S&B7;cJ=^UX@--8+?d0_8UNa(Xb6D
47R@&R/fH:@P:MZI63<D.SJ7IZ(WXRRK50;YML2NJeRVeY,FNdK?KX=@O15YaDKN
MRU^(;5VgF6=HLg)8]B\Ufe15FW_2)1)@$
`endprotected
  
`protected
c01&;D?IU_--gN&R6+.]fDT8d]G\SU/\ddYMT2FMIV8ER\K-__\N()7Qc.9VEcTC
b,UV9\UI=g\-.$
`endprotected

//vcs_lic_vip_protect
  `protected
cCBPaIZ&,VDZ#?=9Fd+7PPW=^-/d)TK2G<PBg&K/)F4#0G;@F0/I+(#?bC[BGSB1
0K)D]B=cdOQ4Dg#T.;=M0[4RB,?R3ND5.fZ5^<b#-4Y3LU,Pb^E#fU<5?)TQEB(a
M:(8Ya57ZA8<ZYHMVFBVL#Zf@V-TT3FEA/O+=H8R?3<Y?+Bb/_14f-?ZUIXJBL6F
-?E:GFVM#\R;/gK,##.-D3<W&\;b>I2EcZ97a>31[&4YO?V1)FdSa5c.da8JGA+\
QN_9/=ICKgNd+5>K493YfcMQZBDU#=AN5H;2K7M\\:XLBH[gIBD-ZOF3&A8KD9OK
&;;D1-&T49-\--9J.W<fc+.1C9=4W2-<].)00@f\>PA;I^A3Xga+TG/YE(/SR(BD
7[=_c)QPb[DEcR)=)E50W@fSICT4,L8&P+dLE:&HU94dS?#.#G:AQ,=@b[4QH\#_
g2&^X^a@7J]@)8T5Da1F-bHZ,@e-[-Q/_H06QC<;HFF5FIO[TYL_JI3dPEEXG0Bf
Y5fGG4A;U6DU9^>D&LI21]0UB?\RL.)Q2>[BgWN\13g3AGT)D,]5H^f:91IV6O0]
U.T0<DA3>O>&[)P=W.=@YRRaB)9=EQ2eBLV1XBO_DBX;_fDID_TPA6JY7DJBKbgY
),7;>BC/A:Y(=EQOGN@KT7O3e:MLYdG+ZLa[Td^T_SdOcda-YEH&@?L)IYX69,CC
B7OU-^RO;[c,WW-]7Pf:NIV].6B-FZ21)@.,AIH(IX(?G6@LNC7UTe_G9@Q63S]f
-5F0#8OHH2=:J@0.+?EMH2N(Zf3)6X?L/b7ac&I5O6(KN5a7,TEWRQZbN5>KMe91
d?Y7T(FCB?^9\BY86;gR\;6aFE6RE#A_JVMfU(WSfQ/_&A=X/KZ2A;Q#7:B1XY;>
EH/bLCYA[]_64)cK.<WNB:cY?,6WAG=>aA+1W:TJ<fJDa\ZH3_S:.UG6@SV\0,&I
/+c=bb:Yg0A1H57,CD)eVH9[acbTL9E<2P@_&1Y;\4&ZWYK;/g_D47^e/P&=?OSL
:D=g=,?9)K(G8/c3;4a;2eU,FS0#J5\=]?,dfIJ[?PYL#:2-ba5@Y+@;g2)-(?g0
WH7^C&5:00JRbQD9Tgg28S8]aR@Qe6e@Y0PMSR5]IWdd6H-HaB^(CH#P?E)X64JG
Dg1<;8QP,#<E-OF#HC&1);:e=W,I1L>Q9\b)S<D)E7D@V82]<R2^RB=:A^^P6Q1]
AOfVHY<?M2QPIH6#dNX[F1Vc?+eDYW2[cL^QTgY.65cCS0=b08NGeLK.QA>3=-NR
WF3gH=TZ;Xc]e.f>=_eBN==UM?Af)_H#9=/CL]NH?7E-5e2?IfXd;H7eO>W4VU9+
/^SQ,9=0IO=/W2fA05F?e3BF,33J2b=;(e8C+0GQ01BcE54dG(#J4=Z1AT9:O=D#
QGPH_NfG)>6F?O/=:/EX)(HK.dCG,fIR:NWU=U(]#=g]g+4?K\<Ef198M(HUe1JP
#b:Ceg>1_5=-Y(5gJCE5#VQFGWAQVMB1\\O5HOSg#Fd]Yg68.G<VN?-FLH7^aba[
@(UL4,b4H_(^65:U7D2^((OB<J(C:1?&+f\5VaK?@S:CT;(VB_2T.4eC45A)Q+#D
6>LU<&6F>aS#OUfVOF-1IM7eE9ID+;cKNGdCA8fYAB4T]dN4L&gHO=F7J;:5gfYP
XKL#X+0L5U&B,K7)dHY5e[L2Q=D9_OH+8CXga::gU1a[+MNB87.O]c6bfXUFa<ba
+>XgAERH0cGNg_.d;:F&5SdA&S,KaEMP&;T)dI?Kb,&=C\c<P:1J;^([[NCe1VWI
LX2TS:DQ&fbI99H,>+e?FAC<@WYQM/UDK47MU&]+M;KL31@&VCSXe<g:>.cZd=S?
-6/#=ZH67+4A?RH//VUDI.70<W=.=W1F(Z[g\gKI_O^</&\)_\A\IJDA5I;^Ia1-
f-3+ga7?/6[^];LO]/\Z^c@1N#K_C5V],ccYE]be#eEIB@)I=ca>2E7PYDY)5d#^
]ZD01=FUN,EIY#<UZF:,9^P3=WT&ZaA/CPX?Yg[9OUbZ6)E-&Q^;eCRV+K:S6N&a
dVXV7TNJH8c.ZZe\U8U2<HTX._<IJN_9>P+NHb.XDA#8^Z\@5V-9;5V)ZC5f_SK0
C#Y-(5W\?OK,4XeW62EG]AEaTDR8L1][,YSI2d1I)B@&G_BTTEGd=(U8e2F;4,TR
GLKH?#5N,)a1a=>VU5P^#:I_OW\=#FR,I/\CS^U]MQM\bS_Ed&4OD6Uec_O_F\11
a6?I(-2C;8Va^VE9#e\>U_c+/J]cQVR-MV#+a25e>C(7a3\g.MV]4TP(Z8MUaLG]
PfGPe5B6<EYH(/>THfZM_NJ19P3VK/879B4F6D>SS_HeTd(#4LW>P@MSZJDaEOX:
9O+W,,K80e9-THW]bYA,(G>Nf+eRY1cdQe43<7X,Ba1@5QVf_UNGfIQQU+H4?^8:
\:4VGY]1A5UE^[VYGR6bI_=A#QKLVb_3)7)Y<6J?eZZAAb>a)L.6V5C.?]XTZMP\
T<0Ve3gc3_>5^_>)F7,?3PR.LZeID2BHS1L;SR6(G]eP[85eRFWS/.SK,H^1J7/M
LY>H(egC<7/W/G7GXgCV0bXTMQZb,;PHfC[cG?D2_VBI?#K<PJB8-fM33:&bL=cX
E\WU?P81+(XcE0B[<#LSB]^7CHG5X8LPf#8HT)eKHY[:F=XM2Q/3LYAHA3DZ625/
fgRJaR^OD\[PZMM-ZU9:Hf\Q;3?]H/JNQ+0OB7cP;\3JT0:R(N>^]<T3DQ\d32C0
HNMRA#M=e7M09@.5A_fAPG(A[T<QC@a=+WKLB\X/>I(C@VgNBX;/]aYHB:/56a^d
,XVIPf^_5Z.JAYeE;IT_[[2?X8]=WF9[V#F;)c7MS3.V251-;Gd6M(\.GM#cI+.g
40NB>7<(U\N=O0.BT(OA[:Z5W+aFb#-,86dZA1>B9[Y?=/QgJP=0;#)(TJd7K1(;
NB:Jb(I5E/8?Cg@<7V1V9Ee82PK3PV.6>ZSPAf6eSXaP2\/9OfOd?7RTCe-(f#JJ
855/bBA0F?Zc\@1C;X;f^1M+&\+;&2&2/QQ0^R8O5(HVC2#O0P#CT;A)C?E:bKKC
(H5EYM;0?d(_0.HI>a[9?@fGa[E5WN413gF[NDKUQ,XL,NG&W^9FgA<:)6WL@Q1@
I[Z-=6g7acdUL:G5_>IU8OHQJ4#[PXXEYQS863?.a=LDb@bfME3=bLGX:?Y5U_R<
7g<T-HO:4c(\4_fO0W_/BK)5d:^E,;Z(X,N_IG.3Z:TRF0B4Q\O<I=E;R(eAEC?1
29R[A,&c95SPb24=KPc>6>#fQMHXS2AGAXGNK2#\OW9-HIZ:bE/DIcI/JD<LWWK3
?3?33FgBfV#Ef=/L]KGF81.ReI;Q=HVbNDC<5JYg?@O;U/e_&:F/SA\5=?N?dQKE
bS7+?c4Q:c-Q7L/@11+=Y:eQS12/[6-VX=I8H?WG4Od(bdH@BJO,E@DJ;#McU.S-
4U/6Y-CN.E93MOJU.4DW(E-5Tcf#NI;CJWQ?bZMORRXV9\;MZY:_9CFPKT2?\7R9
@>1QR:gX+?(MYN3XdN-.<e=KQK2M&e;HC#2+WJBD^T:_HCYV(GV&@J4b,d]R9C(b
dE&K/9[-OZcYDVd\DbZ/>&97Ic2B_ZaEf&2JA/<FFCe::AR,:R(ZP4CM6?T1;WF4
dBG@a--]01=1D&09bPU/g7K,[O#2US=AJ0c)a33dL^BJbY^#]&#TXXSNe^6M_ADL
&F)_HJg9)dKd2_D6;Z8TgMXO=NQ[FaD?FJ9F;]_E2HQf2H2.R(Y8#7@dc^[PI_DK
_4GE7Hb4=:N0)Y-W(SPe:a3b,14?aTGI&J)^]LD16>d8C7b:+dg=GdRZb5GDZK(5
gd.GHXOK/KAI(PI[VX>/_WOKJZ4U7,6@O)c:HT:8R\Uf?((S]d,E/aec@?S@.?<#
/SaU,T5abAR<2DYcaD1c;(dYX,>&<.,W.e.Jf6,LPY,#_N]bT6+(?2ULX]+HaUOd
.&335OSTf>LK6b+NL_<C&Z[ZeSHK9LbR;9&P4_.0bcALcbHI>M#G9NHJG)\RI6V6
KPV_K:[STN[T]M33V:F9c(8F/RePdK=eC<:5ZI?db_g=K@5OU.=M@(_FeL8HELUR
c<.NGB)IeCDI;C1)YC>C-d1\^7f7X?YAaAd,:I5KYL/R78X<1FIUW8HA].4_-JT#
0e&M]6,4,>V[T7)KRc\D3AV(QWJ#8R[A8-GfGf#35b\Z3SK\.F_IU<O243L)^_)T
-d44)D.Y8(\)STFZ^CZ8TPQAAD=;C[4-?H-7^ZQ-U;aXXBfE0Z^NW,K8<Ta#+<g1
aVQC1g\bQ3,>CE7J@;HPY^3#VcET1]??3YD6aJ,dfQ4:-I-PH=LP-SbP7CH+RN]Y
LCCdV1FD)-d;F3VBE,^?)S+U=\\I+bWCKCZQLg648C.N0;963G4W9WH96?3NV6dD
-/J\N[YC-?#N,YX.:a@JR_22Vd=FRCR=-R62I1H1DL]VP>W9S_=RHI+-,3QX48P@
FABcH:DQe1aBg+X>AGPbMVf,WR3<cLBK6:R^HPP)5U3]??W\E+ZbD62Y,2@0]:[H
UUXB>I]AZGN/88:E2>Z/I]J@O(9ZE-T2&S)3.5)7TEAH>CTVc&Z.&6JeL3g0Q#]?
Nf?/?&ZGGd]Mge_8?D^>#PQNaCAQ.)(RaTZUP.b<@dS@OMC)CVGd7#c7AUBCAYN+
6KYU?8f=A)B7X(FVV)]CIWcU;LTQP1F4OYH63aL]76T_MI<XG<b><[?d/@g8f)LB
/>B)c@@Cb\6[L(/83eM(T[NEW#O0SP-&.YDd<6-&8(#XT;g-7VR)Kd.b+[b(T_YO
L19#0>]M^S(E#:KM4AT(:LN69KWG&9Y^VVd-J^J3N\RQOcCELR?:RKY^NWS^IbN2
)6bfI;_^5GI@G#,S0-N5GD3MCc1/I=M>[f4d;V+_2VS43gQU=+8O/,?/:Ea+JM-2
;VLa<X+:cVa>3+6;I8Bf8VZ_;MR)MA#5#)1I9PO-?BKF=GC<D_HE<6dd[2-#=3bc
V-DL2=?.D[f#PAgE>Bc)T,U8,48,_@OGNM18XdG/P0UK_b^,S8-?WeF#EU4,ZG?6
7M7ggHcSc\YHAQM)85Jg9CC0VAB>9)#\.6b/1A@Ia<^IR&aH3/UBCYJc@89EE#]L
T&@Be<3)D_YcXdaeUE;4BIK[?eJO:=cZ<c+V\/S7R8E4=>E\ILR5gg.f.)K1@>ZG
UV4&2b=#Tf#^=76#)A7+,>7IOV=/VTO\?WS+BWA/1+L&8fZg_#VJ5RUCBOJC@WN-
H^XCCN]C39S[Y0FAL=YN-+2:_1M[S2FfN2;FTRZ<1P<(Ye8a7]>,^>Z]W?9Ib\:6
cB,W6U=g0=c]LV<02D;7gYC2@)[+/S2<?[EfZLAX4B^PAAYIKO=G(,d9_H;)Z,2)
#0?:gGacRGZ6)SJW5P&UG[eFCJ<@BE]fS0f+5W_MP2-Rf:2NG3a]fF,>#;P849a,
R?);F^(J=Y#VQAX@6]E960&OM0@_JA??ZXA9?5[?JcF4GQ8#^JAMTL+7]5T6JF+:
Q;LT&9PL1R#,;LRMBg_9H]9(SLMVFEK&P^2/3a0,<8C#&LY.O@V-P4AAZV[4)<aU
VE\IQQ.YQ5^/ONJHYWYR;K-bEK637f5K>+SdJRa3^@2>@UfL65W-E38VGP2ZNUFX
+<bB.0MOUJcVUbCINgJJcMJd&LA)#ecMHMdFG>a&d6;;e5&Zgc0UPYSJ8L4-ab[?
_&42Q;=M@b#/=Ig=Ff>dI-I@-LR#/=;aAPB]WPCdTMfR1+2X6_89)e+PZYBA3NR=
<;#Dec(-D9/7^9PZ)8=2B1UC+a4V@Z?ggQNP3U<H-;T<UFXd/2ADKeXgA:P7R@H]
g.46&/Y8.7Z>-=A=KD+>R#ecbNA.QcT[P07XeI@3(HGVS;RC^A/^W+/Ed,<\U8FF
,Z7&_NV2Ia@##N75b#^b#Kf8:5ZY>Y1O?SGAQCG=/L;^SQ+=E=]C)V)2M?<_3(:Q
KPF&E)MLF267TNg,dQLbGH9HP-D/,IYc=-bH)#\A?F>8Af]1Y88,:0)WReUPR+NF
&.2X_SAU&^F)9C,P=V1b(@P6KS,eN1fV\TV8[_>R:?\Sa<CQeQJ[a+;:MU4.QB,C
&#]ded82(@]WGNX5-:L03+T&d^QE?OSNe+=B4AQ&I+YPNC1S5].4M:<BU\(]bK2-
>X;VS?Z0X^I<6NaISOW5S09)&>TgF)7;?QfBNB,(bD-IH-YDCg&?J#E<.K@:/F7H
-^9?W^N:\7>]5Z+);U7</f)8V>UZ-JXF5>4B>]+K^9MSZ#:(/ZX]@.YaUeF6NRIF
1UGN8NNR(Z7(.5:g(OY[/>0XX^b7)L2FRd>9H4@<>>2gfC).XF&Ia>XOKE-@=P<X
SAG^+bGSeVGbXXQ96_Y2A\YgF7>;bcf??A/?aKCd9NM,M)G4R+KFY\NW4OM><3.L
9?6:cd,acSQ@DZZ^.:cF<^e^,O0bfQR-+_UgEf&g@QT,eZVe94fC?J5&:O77&YEd
M,GIB_7ZTK]fedY_-7<89OTXce1Jg-;DN2>]=/D#UfJZU(V-.KM2e4_-cQRSAQ]&
_(-IP?RfZDR0OS+cZd9OX&S\/>a2c8@L\D1#;C9F6RddbHE2MMF1\+6&e;eR3&;-
28=Ag#[)WUNGON,G<66NI4W6a6>_)7U4-6#=R)J?&+9U(@3f,Ab&a\^^5H]=@43O
4=2\XY#R6NU79Q034JIaa]>/CIQa88H)54[L>H>O?:R=ML+C,H2/+K6J./^/>_]V
<P9,2\>QeLUK<&O0?cB3BEVbGX:a#13NZC^1GTUN\<?(M@D[AQD,N=F4?G=ID,\E
AKNEf:5B4#[152dY+f45D2YFUWN^PL/KTJ+&+@UK(a;G=d.FBdKY@eJd@R5fSX>[
Na.X\.^cbFR\Y#a4BLCR5f<_7Z[36YL_f?&]-V727XPD163F[R21TEOcWHD9G\;I
M@#C2PU>b9cbMPU?6GT5LOL,(]^,SRY?^^K9&ZA8+g4SWT8\aZMZA6?H.#.d<=e9
&d/=JK(#48@+,;X-AN>Ke89ZQU<EZ\:\Dd3P0b),3dPW1.a_YcBEf8@(AG=7\_gE
#eZQ(77UAD#SfDgAEN@^LSE>;53LcG,M?X2_L[G3dfZP.UB=L7GU.D#WEBLI[KBV
f^AN<6_8V<38FM/KgCNUPMYG[^cdXAZY4a7F&Xd+0U#:#72<NP361);V<IX2UZU=
YO8b[U<7KKV;c6K_5d8(:8ab&.J6:O5QW_[VR[S-6<P&,Qd6=\?f1-4a#;ZAKUX;
T+BY.(+1ME=QI2CX.1\2c3gHDEQ<AMe([?e,-G@D@8;=H^QZ_DO04O/c\8/d=9HC
M,VTA17MU)baWGgYa)WWLc@/\\e&g:Md]K#55I)2&@9Z;^S2/I#EO+-81:QffX55
;e9UU@V-#J/OKd@IZ&I-?4IAb;a(?.c:c>N?cFD3.QCCPcJ?6HEJWb2J17a)>gT+
VcfIBJ]MX[^+,-T)DT^eP[&M?)?)-P3+YNDOa0Z(GZ;KAOA0.,V>XUQ?+F4(1+Te
:_UDgP_B@?VL=LABY+dF()bC3BOEN)[dJ>.1dV_?d=B4/@=8:RA23d]-&GTfW^bJ
W43^Q3e.NU0PR-+;+_a2CDZg4AM8_N::0LPU>)Je->L^/cH6_S89N/A<V9<eGG[E
>2Wd5.gEY2N3F+0_B8(4HE[bH^#>=#M4\9&_6OM=?8<NMO;QabQC3E1(^_\9\QF/
18;>e<LJ>ZegJYGAF#]R7BIJSK6PH2+8,:f]UES1N\d5UBf@EE,):[S6:XWZK1=K
I[^X\(JbG^.R=5LJO9-V?<g1\&T2f1faUX51YJLQV4&7EUR^(?49^992T7DC=UR>
4Q-eNXdI<ZX1ZZOPc8>]&Q_eHF=Cc(#T8)ReXC^..bX0BdIM6Q63RA0+BOL/IY1e
7=\@=+R1\OOf<?d;-AW5JRYgEcQH9gGND=RZ?<]#R(K4Z5;;.S><TeD?/B:Y-OWM
?L>K.)Ig>/T]Qc^JAZ_LgK5H?(FbCfD0GJ,(.=UWQC#2N3VJ]47#V09#R.QVOZa:
6CVLfa4;>eH_^f[KG#I;_6>C-0b7J3:[Z_HCAXSZQP5V-/DJ(>0ec#MXDcFVF[LH
BDcR+:A#bbS1TX1V8/@M?H3G.]NQG@@,)1]gO1+E&\1E[/F5eV.9(GK@BCHH0356
0aRa^P5(2)b[223;RQ^:4GPFOb:QNOAVVE3.c9ZC5gb/28.D[2X.ANG1>/2c9O2;
171W>9<V\bV.cH77\.d>3OK1)6W9b]AN+6FE)5?/+X5-KI<dP?:=cg+;cJfP9VUQ
ARU6Pb)2^6KB-J#Y\_LaA9)f>OY6P<3Fe4F/0gBa\IPaDD9EeH=;-^<#c)S&VHda
WS3,Y/#<,]?G[XX:e@7\I0.fC-TL,8J^g);3RbZOJ/].I,c;^3C4VaHP1_PB:KOS
0URUbQP(ZB,,0=LJ8H\DRO7W;ePXQD_65=+88FLUCYaD8X)&VT,L?>eXY0/-SAU<
cFG4R5N#4U)_?]eb:5FLT&3H,/X([#RJ+DEW^O@V<A_7QX-=B:B2_g9g=X=Q<K)H
:d;8I?RZJ4L#G00fgRJ,&#BG1@XH&?a,0CZ[GMeDCE^M.D;P+:McX?(:dQ[L1BJJ
MPB#PORaM3K=LEcJ:Z)]G)O0WXF)]36-dV2H.c@UV)e\c<)<Yee/5.P&^5(W/:c?
D6N^)@;f(Y9[/7J;\D+PHD6N+O>Z<6?.^^+@_Kdb.RO8]g4(ZG@52R52.4VBK;[6
XJ,SA^--_2.#83da-UJU6]c<WB,LUgb+eUGe8Y^4^HNg3.?NRXcHO.HM#1E&+LXC
T2#C(7RQa>X:^dT#\ScbHA6BaSe#d3ZJPA?K^3N7b,P.#E6X=^])L]Ag0A8^Qa^1
6VS4eG@;0OL.G_@:-T+U,VOI-Y>))fCFaRed7PU^c)W8B:Ubb&\>_Nc4VH8+<J2_
D;F7fb#J(V7eZ.E+\I1I8?P.2OEa)8,@WS<,ReV5Tcg(HB5+I\e-+d?M&5\1>LYE
8_?1:6#IQ8fdTVO6[-TbQ&XO34\)]RWKYQd[1/[a@_GORcD/8_==),I^bBZa\2P3
dA>J^-OcFL3:^;AWF=\P:XV1,9Q]:6TLLQ]?3-[LdYO?=@74[Gc#cIHC[TG_Y):@
[G.M)=+6>RTb+D&&7FFTT6X14F30XZddY@#d;gWFf<D6O-PdMP)WW2daB(4PEWX7
dGD[B@H=DZO5B<.e#-(g?B3T0^(K#&+<M4aB[WUXf-=,G<)ZB67<C2I,V]V1M;:a
LX.+/&->:;<5.TFCL]C/#JIGb,=:?efXI7_\PHS51C[NLCOQG&6M3(7-L3:?EOg-
Q9b<aI#b9+6LA/7:?.L?2,M?bO:F+3=c_OI)R>&=ZG/>aUZ2g-1QS3O5BD+<K8A7
&fT\UVORX/>@8QN5]_FMOH?]HKZ7BSe)/]0T:&+)fcU>ZJc[.E;dBfH/\\K]QD_N
4(S.4&M,U3[,=8=3KAUYg(80-YRNED9F,:DI3b6++MV8J@5I7FYZ0Ng7OMV3RBLd
E12JNE&6T<_H,E2^7,8,O;Q./#8XL;g)K9(CX#aF7GdGS:AQQ,+a>MFbXgZ5J:>?
4a<2H83a7JT2Y+0^2b1Y[dY#4#2#7-8/\aBV7.g<LM-BU;/Ia;R3;94?:D_,L1&S
79W_(E&g-D7D;L@?8G_S+83]gXVHS4CA]J5::=Icac[-HDT>DDML];FZDS,-bO:g
f;:AKW>Y)MY[)_#ONJ7fg3;7K4CJd?[WH0XT:H+B]K<^AFg.S]b-;0.3[c;caL&K
+W:V+?6F4O,,]Mb(\4T2W6aV1(bQ_A3a6#VPG_,1+R=e29bHDK.3H4)f<QKd0bFO
3\EGEK/8-/-&<ZHYJQf(PX>d090M67S7T,,O::.M@2=5C;S9I_0DUY=ZQ].\VQ&B
3@8L#ZAdbg_3(L&#Ie8dE.7:9/ELO7)],K?98Ld>S:N,M^deUf0X;X_WCHa^,,M<
;;4VCG+/)_4g:?=bO9TN]-[8bS]:]R,gY;),G,7a,fMg_IJLD(3N4M;YVB<0DB:M
XNM?Z\0E;QXbVXT7KC09<@+&1E>DWB:D<McSdd5XbC_76=SC,;I=_O>]&T1&)TKS
Y5B^0.V9Y\<6OVe,(1140.@Y[]@XR1)QU=USB+VM+>\L#<Ib5)..,2B&YHVU[1Z2
UH==@.0=2P^7<FRBNg]9Ic.KGbHb)S;AG]/YcZ07F7Y?<DFJ-2)[3PJ;eH8-g]16
?QbSdH[Le+DUTg)d3U\T4?7<Yc6#M>=8D?;:CdQRLZ[FZ@#^S,a+L?QfL>^PF+QI
:E7E<+EEM;KO5::4Q[JUUd&W3]4&-,:(H,5Z9bQ6RAE76aX0H^fe9@]LE;e6gD<<
@,IbSdFg8SYZJ&ac3dV:g\LcVC?gH#+5LaQ0gYL[SD]6[B1MBDCgD1E68Z?BI7Qd
TG@CVW>TV6-6K.[5AN/K#&d:\^:UFZMC=9>R+I;9;M#D+G^<RX4CXO5DY)FQJZ;E
\[2X>LSUGL7.0X@^CNQT-4AZ)-+f>)-SXMe1D]\RN@a:[XB+Z-.20#,0gT0b08>4
RT<A&=^7>&JQ8^S3X-@b8Y0(I_OVQDZ<>a&(>C_7CJ[80K-cf:>N]&0EY;fPROOF
0=aJe]80)8aJZ_U^L.B=REBJbVf4U4JTYI5@,b(JV0HGIV14,(TI?C.RAG6[g#TS
\6f+cG<e</D1:9La5-R0N?72g=g8U9dF<5ELc,V(59DLP2CTJgZ@R7I[UAU8H9eE
,&Z8125cUM;:\]]cV<e+J4#YWGb2XbS(XfE#;JFe;C5I@g>MMXcTL]M4PCd)IaZC
f,#C_.g983(WFN@+&BLUa0UD9P02OJ]9PV0TGHQ+I:I4f0Re@QD>LPb2VT9S:aS.
6F@17UR32;e<f/FGUe4SG6ga[@YO/Lge-Zg+U6B[&2WCZ+1G[FcH>(C:[U#]UA6T
MJQGeSUSNY(6]DUOXHPSTIJ+/A_RN:MT[[[G/54e9<LC(fMSG0E>Z+#@01&(eb0X
K4ASeXWCL0\&B5-+_c42J<WH)4TfbGEHOQ_02V@N?WJT^1AR8_\N-_SQ9X4bSW(d
EcSYg)X_32H:6dI1:Z3X(S:T=M7:AN1#aL?^12+S?Q0e=<f9[ES>>75/S@CH?9Z(
\#V4Y5eZc5:GQ=SBSe-:G-M[RFG?Re).;[F[+7TJ:gWM73YQcUV_Z?MdaHFPf0X0
7:UX_Z[M6[-#<a09_APFUL/R,C?:?GDZ]dC=\Z&32B8<AD.5N15Y0135N\WPU6A4
69?N1?H9#MRJ_.aOQ03&I=@N,SKY/cK+EEKWcS97&JN_+gZ]>.:Z68(.F],O[/dS
POW[3HWNC/RF5RgOb.:BK+S=^Q^/P94?FcG]&)MK@;<O6-Q:A_1]YNVc@HD>ED\A
[UC&-.MB&gN,/^a@;<EUK;EMOVBH:GM?MEaKR:VW\+9X74-9WS[BOE3RI=17_K3@
^0=]INET1G\JMU8(ND6\&385KP9(,]=XU,=+]O#:>RL59J07FQVN&P9IdD3^L:<(
@X3@BP]9,90BV0(<Ag<Y2G8Z[U/LIW65?.\G:BECI9//_0X2YGHB&<#^,D6KQMZC
]79:69_1Z-N08BVe7[;]b[:S-R3H(6P0(]AfB+Sb4K,5;X[^-b_<_2[FTM2U[Ob6
Rf+d4F:0gc8ASBUP2B0_MV?V,\](Z+K->>N[(>/1J+HV:L[9Yff_7aV((?\3MaWf
f<W[VQ&I\_Ka-E)?9UUCMbYJ,d?T;0+8^4eUNM69(WL\2^QB8]R=3)&BAP,KOC7(
5M</?OCgD/gP8@PTRH8+IRN]OXPM([Mc[3L+K;KCJ/-AJBI>cgZDgFgX7#,P,1@f
4K6D@D]NcJ[A6^#R:[/YA\):3-?3b(Pd]5Y3WXb169^4U9YL7YfA6<-0F]O56f6O
-\VR#].D5L;[PBVfe#9cV-]Q1DD?]YN1A]6;X<Z<UIaBIPTG3gLO,Od^]9/>K_/]
Q^KSE<YCZJRR(DOM.N3#@DeY2ZI<BALP5fBT6DI?;DI]IY7HZ9e2S[;EQU2GL-^b
1/L1DCEM6TP2I6@g0GCRU:3I9/VG:ACOPBf(5)_(^#GfK4g59EVO>f.96cN[V^I;
g]-HOZN,Z74Q,DTdAFI[0Ng8?I20J/M.8FR?_UgOF7QZg8Da7/#YR;S6\5PS(52]
]8I?_,<#V;KLcKVTM2[<ULWYO]9a[T<QVeK)@-g[V:?)]@WA:TgAa1S4G\8QB:N,
Ea=19WXB=J.gK66N>19Q9S&I?1e7A&bOaM42X/H>HH;U0CH[.I6>3(UZRV7OJ7DC
JI=SUIeWf+SM#5cg_S#Ka4KOQ^)C>RLTL:JP;cI_5fMZXa@^MTd6+g/[R:,SITZN
WT0>2:_31Y[OCW=_Y(]DIUgXB5.(8RR4OC0ROHTP6Z)7aN_EdRLcV<0NN8J7gIT>
.N^(\<,/cGGCA=&;2aM(;(XDeAPLM8^8[gA2]]eBPL?(2,RFdZUPZ6K=M\1FgG&]
Y21G4^O0^WZAfWB[7=4(W31AZ1EGCX.\BR_(:N<KP5K;@,KG]GFD=>_OcgF4LH)[
Z^VdFa^?OXc^/5[.8;7)ffBC);@Jf.&@6,L>3KFWJJT#/1O2AT?AK;b=(Ldb\KJ&
-^<bXg@NN3^@?:bW;Z_TeDE<d_Og+YV[#PHc7R),3PNI5X<2KR@LaNZ[1Ef??dB:
1a9D+AJgLKGDCUK:f6cN+2YLX,UTJUJgc&G)Fa_<+,W\a&9)V7W0g\EUF_3(RM@^
LK.BX:8?ZBb-.U>e+\=IUKd=eHX95\(X;KbF3NbFF=W+V\_UG;),FB;#Gga4QP[V
WR\R?::Q;eG4fQ()^1H1]74Ue?gU+LV_Ff?XW=BaJ\f,/C\XEO,g1.CIdN:VV/R9
OHg:.SKFf;@T\2Gd1,6Be\D]Z\F8MK6f+R:(LOY&?)Q)</g5OU,dMLU5<HU;9UZ^
M-)1(4TY2[ggU-;DRVFR,1B&W.HgP82,;K?\J6V5ZPeB7/7WB#3&;8HOfJ5>MJUY
=U)])7>3AHV0QK-6[_<WQ6_.4d[[EK+@VWgSbAUNLB,&BL)@>4Ia.)(A]V48WG+<
E>8KdQRaZ^VB&EQ)K-(-?QAb>W\KOZ=5c#&f((>(L:bK#:X3gbZPE0.^VEa<JLFg
:W/Y.A4OR/ce[;V_IP6/UdH#61bUaa.-<C-CW.&6N=<XA_U3+:\PTL12F]5>7;cc
(+7-XEBZE9HYG#795I).]J0+bWYN40JOL@UeVF(Q_&X-A&5LIU0c):F_6NgFJPTW
LRKXJJR2/]@H&49DcUI<<<KDNPK&g49.[1RC:0BU?V(P3FNW>agV/.I)f41#KS^Y
.R^ZX[;C-WW_2._f?eIH1J?Z<IfC.;ePFDVOde2-2/H/6,2_KVRF;UIgbTA)6ZNS
+Z)1FNB-)E;BLSY5ORfCYbCL.+bLaA#<-?CLV:[gJ.X8gGUK-P9aP9D:a)L5XI]D
_970c2OdQ#T#6W-,2)0UBF@+WaPNP2PC24Hb@a4Re0]SPRU14ed7>J9_+_B6S.,4
-]PW>E((e0Qc>-4=5IB=R/,Y;C7W_OFXC;X+U8>3;a5C90K<1eL)VO4=C.Eb4O@+
BC7+F=aA0f?RQVIcd;G/E;91T1gTWV&c6<5W^34&A:W<b:X5B;3/GXb:b2@SYAAE
/8D+XB.ZF43,6T85)KMN\OR9EN7fa>.-AZ>d:V6APM;LcY]aY#5MR92M9>d:/<;a
V952L0;#V:g<</0K>D9+NTFOJ:#fZV_]U])R/0ZH_GK&-5;800B1+LCH#:+/]6+a
;Z&#FY9,/1L>[=/NSC+f:Q:F?0#Qa.]CCcJHR6N-9N]f/\6N:Sf6L#>8/_G>L9He
@GQ+OG(R54]N&Sg-aC52LEZI3W\&5Z\KbS=V8?(5TSPDO7TX]3Z)aL-eW-KGYF^4
c[)f0dcCeQ9#TR@Dg,A\,@[L<48F51GI[TbZ.g]9<YY<F=\F1O/1N)Y&;6T;G:FP
c=U06I68>)).;P/0X:=KR5M1[N_(,SZK8.:OTNMLJ.4@\^\VEWa4+_Ag9X&(,#a8
AcUeEKRc4=\4]476?;[a:c0VB_GVDQ-Y4;MP[)_[\LI5F#Dg)(KZ41e0XZ\,=fL2
-:0ge2D6+&#8C4T(?3H/FWWP2V76MYe5@+B3_YRAI\4MOVC=O_=C:LB,Xfaa2DBL
CS+-5JDN^E-OYC)=bE-SL+>K:5&H]RR^6-73QL-(Rb3(\FZ(3J&7F:LVYSAN<R[O
^X?,)5Tc0SDeeaWLUZa9U4GZfgf3<U,g&??-BPQ]B+LO,#99B5T]66K8T.+c,_Id
A,2^-]14#[W[e1?g73YWST?0[fMT0?(JZ]A2\)#AV2aYPM+e6J0aC-WI\cJfE1K7
<PI)I=;5G)5U&1:FSA?B;KNWDYSF^;E66968c5E-USR>.R^]H,0&a:DZVD=WVZHe
0>Q9[](<I<HFG5Qg5&D6LAO;6+W\77JbG_7Q7,S3QI2f>B[M23:1+UGE;F1PPNR5
PMe-[)3TQLAE<A)R6,R+6[IZ5V]T1(VECL3&W@@Lge^32N>-H/VRJ_/>bJW-9=Wc
_bdFZE+?fBaVPdQ3V^X]c7FdHN?J6,&<VGW#A(c>C1?LHg@Q-\;bWYEN6H]BAg)N
8_M9\\CVbW,(E,E0beW1L9#\U1aC871CdZNEC7^;27a7c],&K9;NU8_H38UgT-+f
eO9a)B,?>FP6E(FQ+KIRZ\dOJM(W+NEa[S[)T(7]a0G(M5M9;e1#IVR9-JEBQa>9
2fLHHKf07VV?>#0<[Y--\b6cCTWPZZP&27)@H4fE4NJ(-P;-64C22>ZP5PTHa,7&
c;+ebK93#;?EM^OZ&G.H0>4IaNR?RHSP?Y,(Q+S8CU;PNDWd0=):.5>7_V9?3Y5+
.3dRW/YL?.e:9>#KeD?CHSbTQ^MSS+4/1EF>?;,8:JKdDSC>3HE3gXEdGP:-R)56
O?dW</3gS/IHC/D[+;a&1@4[c^KC^S?3ceAP2(1@]PTXIRVI:6&&IEQCGI:XdNI\
QS;WLGNG6A(M@+X3.3.I\0_H:ZWT^/_5J>cG_SKc93[WY/./)94PFIBTY8H.6aF@
\_U,6F\eC_B?b\_@XFY.fN6^V\PU6H3V3P-SFAY;b2_.,cd6Y2eY06L94NA0X;OQ
X-7,1c:=#SfAg9-)K@NdNL\_0KVDC?Y:VcYT4Q.--UeYO6.3LMc?;2G_)\=:7#W6
SBAc[A])Z@[.IU<5\A_OdSI;BK#A_4V6@/NM7M>=Xg.^IO>MN8MS&BM5GdDeV&;C
MLPJPMKW_Y@bN5cX;=U,(N7WV\-WTWHF>MWFHHU1fb8NM0U6<?M_aAZE95_N-(IV
,fO,SfC>VeXL>d^=K?BJUG+L6@/,1ed(NF&=DS:&9Y^<B12[g+Pa^#R0@_+Mb<d7
a]&IA#=ceHN[EHH\Ke@9F.gR60.5-V7f_P3EL38)Q@6:#>JK8)Uf1G(32M\C+V^_
ecg9K;@-]<HY-/7Zgf1b&H1[cV7]MUE+>LYX0=-<&@eC2#UWW<f.+ZBT/TbX]@H4
A-V/E]C7:49/SLH3M_/US;RdTGVAcHB4E]a&4AM5(_^=47g+eO:V:bZ.aY;FDENI
1[C@(.M-:U)e77<6VUVg.bRZE-H-(Z.)@\2gTL^GXYFLQJNT8^FXc-F-1XeRZ=9<
&a.+GT_O&6DQC)=\a+I/gaDUFIFI3AD5Y,/N7\<,7FQ@=CV0LG/M9-;Q]/4]08.\
6,8L8_a=_<2Af>SMQeW2\>HYF&dX)A^6dV5Sc&VcT<\fR2I^bL&.\^VL22e[L<S5
,8Nf;;XdQ?]gZQ3^]?]HRJ^7TWEW]K36d9[dN2#bXLC4b#P(GT/C(6?L-XN3gdHG
_4T_0]c9/^c(Vb@U5<;[2H6g4;4Bd<\&I9F2V&@N&[T;/NIW.T,=gZ]4T>UYOB(B
5ZDX2:,/9QW-2d0=ddcV<9c(cbH1<^GJVFIg>a1A/^.K,&9]>06#TaI>,6C4(e[K
S_JV(1\EP44FSP,9N#ZgK5,<QNBK&=24>1D57YA4N:503.M/69a;bYQJ[/;SA\S(
CL#<0?..Wf,HX_9C-USF9/.&0)b74BS?=7,Q/MR3(-,ME2b(:TFfQJ\S?GGQU\A,
-P:]@[OHe#<^9S=P,])_-/LTOV^WC:E2\H^Q@b^;K.P_VNYVR(Y8O,a2>?-4[K5e
^ATR0&O?]#D]+J<dQd3KYRIcKF]K&J8_20g348b4CC=7K>BWR:F)ZKPX6DJ;^#B5
_7=8aK^bYBSf/;6LGU\#(7&FTCa:;6PdX,>C(d3?B08CZ(BW1\M[RTLE,YLJ+AI]
eY7KF98DB[IP1gQfB]a_;5+[gOd.@.1G4WJNb+^^3<.f+2_F);R=GH05]ge&eWA=
A+dK4@&6--_O.AHA^SDUT+2GORdP<FT#E@S^134?a;?9P]B0B0BJFe?e=Z.G]2:G
0(cC6-=XBQGJ9a^?2_>SOX5[Y^1@D0K;2M2((beHAa.Q#8JF_59KF3UQ.NJKcTfT
SGPZI:^GZ6.H#3VNRg];2&^XZT,56Q193VgQGaU71QEgXD\HJ8M<<XJA9\J-\:<)
M-Y<GEVJagO;ZXD[_MGe-Za3(eBeM//Q#NR/,=d^_0^Z#+Z-571^aaQDSa0W0BHF
8B3cBC9[)+=.[N7GC>1,])a36$
`endprotected


`protected
7XfGW7B<Z[FB=HJf/OgUd8?CO/Xc#1b[QI=MQc((S,a5)#S(F14Z&)FR\D-QY1=g
2^eS(7XFVd@B0$
`endprotected


//vcs_lic_vip_protect
  `protected
4c[\J-Y8H)Sf\])eL],d-<@]HeE\U-b:,W>>X?GR[=RVbQKc>d+I7(NVBOCZ(JV2
&Q<g?S>X#[F-A65W0g+=L52QFL;E[@fK.F30bKUfN.fQ8CFM=^G];+@H7\2860]:
)_;11JfNFa?C8,3A\,(Q]F(OBPV5/bW72?/8dH,,-P<0:FaFF/?g6T[gUM7Zf\HU
ca7GYOBD?0:4g8#M=M?OTbcQGJ1Y/c@fN9Ia\#X8A4fI/[DR.XFA?DXGKe;LK8<F
eKD,M</-61bC1P-=2U:4a&V+CY@K\Z^H?W:f3?UZ0Ob32\G/OYbc^H[NQT(JZ^].
\)(+O:E5/=NE#5:T1ELUTd4Y)C9/(-E>CR90UdY/YUEOU^MI3ECW&F&5,AXbg1UK
ZK.EH9N[,6-:>;5_F08DJgUD\bBT:g:-O6(\0-#1^@fL^fCCU)564=Bg5Jf#\)76
?b7;A,0QXAA5R3(Y.+DU=#)_0UH],,\I7M+HT&47M(2CK<4d5)6:)Tabb(FP-L#G
OS:&:53MYg@F343d7_32F/Z4JOF3VEd.FVUSfMI=LKb+O_@Q15)4/HS8NMCOc=F#
_)2\M_1SR2+[L/U6A8,([.T]^O@W1F(<_6FaJfZ-CHcC3/cU>I2>GNXE#a#SO;[[
FH,[KaRXfM4J=EV2CIU9b]RTB2fH)C]a^Q>dU(ZD#/->?NTb92XRW_P0+XM/MfD>
EO-4C>U-W6RFVM5>)CZYA>C<X#M<L74KdJ<bA=188Ng?95cYg<D8#66)g.IB>.Jf
VCC&]Ic<Y-#LVe/aB_?5WPM&545\Z3cAU#0gVJcVXOdW@[D>4ND@#ZBH;OR8:G&7
1MX[HE=]3>Q(G4_?598c_>)U>fKbdVDCTaKFC7V[b2AGJN_^AH5TP@3^RN@,^-/5
ffU_Ya)OPH3/IS1);Q4)CDP2B-GCF_)@\2&5MY4L.0UZ.Oac51QO:]M24=P^5F@T
Q.I@3FX=EC3(LNFX=;E=?_^V)LNEN#5a_&??,O&YN.9OAC-YITT+XX+@T?D..A&?
TVf1W)4>E7+4fgE3>8_1[.Y]9\,?gfB,J6.3)WXX8XZ.e66f0=F\4=_IPY6Ub3JK
^1fdP5_\.F__R+T3\aW02dJb8T&C2E9J2dS9UB[&R#:baBY/EgD\^/].WKIac0FC
c2BRfeg)9f-YWcI=g@]W/]ceK:<>SL#,fYQ0F4B9T.eDORb>e:ILXgBaUL@T4W#Q
>HVAL\1M,A6WS+H/]b#72)=P-3V([.FAWAd;@VBc2?3HUDBd3\FC73Hbe;D[^KM>
\e>9YIeOR0N7_3ZXC=7dcP0Re(,cL0gL85-I;.+_DO<5.HRVL.0HB?A&7gGCC[\5
_&)+YS++60<)O_P2LK]&/LJeN<BV=cLd]DI+MS,JYMg1Hf?@1/@)8[6e2+?=Y2>#
QRES6W-P2K5geEFCM?6L(b>Z,7(.NGKb5KO,c\LTH70cOPU?ME9.6a>Q1.3O4d7)
695(aKc2IBP].&7XVEXGaZ_=f#--NV_;9G]3M1VN<W6W#AJVCC:V-d6)Gd?B_.RL
-+\&:Q0?6NcW<a#;+WgP,0(_PRJ0]9WaBDGX^JU^T5f9P914Q,aQWW1:A7&eGI(R
2M2LPRHePK]g;g1LbNL1g529)f:WY7>T<7GO@JH^K6g1U#(O.R4c\]8Q0HUUE9EZ
(4J,T81DNV2YY(>=>>Y;#R.#86Q^A_C,[PJBNKA8.cMMZ;/.Yd#X5J,//=77Cf@E
FQ?3@GC&B:21[6dgX7?CAY0(9@AHCG@Y,eFGSPOK1(4R2\ab@Y[Ng^7b30BfFKgb
2a=RO[7SM(Q(O#9&b??YE:BRW&VY<+b1?8&BVgV/[\Ed+g=P>M]^g<DD,Q\E28Q/
FT,=G[RJF+eVUWT7ZIa2?EaaYY\1F)JIP:C4?@\7F6=\?GN9B5.YG)aE:](BWE)9
5_G?8TG4ARaL:D1Q2f)QIBgJ0Ea)F\G7@4d[&@#3N2ZP<?;&f>F^6PR70D<F>,bC
VIM6:66.-;X@)^FVagZ0,9J:;;@0MV1c]ddQTde1Fe51aSK95H2gJS,/9&(18a/C
T5Kg?_A:J(eTTCF89e4K-Q=593e8,]<X?5#4R85(d:)22H1P6;<d]Yg=(X#Ce-6B
e-_0La1dQ../P<5872)KB96R<:2FG0HZ0Y8AOO;RN8WRQNND/Z:\BK(3HCMF][aP
dRR#5[BZV9F?4O[[.0R:SI5B\V=V#L7(g&WN7V]Q0=?O.WB[H9]NJD)T[/5Xg;Y6
9XD1GUSL\/KgM85Y:/e\(6WU^V_.QF1CgNJOe=[E(]MVbTOK/B@fOGVgaVC;0ELc
H(YdU)D<R\UNX5JaO[P:Va4T536Y#DVN+=YTSPM+_2^RMKbJK782U0fg4,..)7\]
7:]TNJX?&M[@f_RB>.V@-3+PXObENNR;TXH4K@\U8GPT3f0Ea7[.d8,0PG3Y1O?c
F^/J@,<J4SBN&TAEP5LXG^]gL6>0>MJ].ALbSb^UQ<8NDWVWgfX[Ya)>;L4KcdL=
NeMI<PZK1X<2>cJB0ORHH,8B]S\WeL7.1>d\<=Q]FXH;X=f7+XAc_7dVg_Y,6RR(
JHa8=+;_.GFeKI&SZ2eI1+Z7(3(d.<6(-_d&:1CYD1/K2:fJf\4)7]U3=VMQ[2>#
FT..I6PbE2)HXN\]EU84&5]<W>7E;;72L+Ag#V<2.;@eWXX].cT3,.V&QGEe(93@
+>T^dM^0c=TY2da>6JL.?cb0&(c9KJE>@)BOaf9BNZTaCZ;J@Y_aXY]02PH5]DP#
2\H)EVX?=;\gH<J[[(/0YFAN;1Dd5;SYK1A<PMIO@8_VQ:(R5Acd#+5g-#fBL8>1
b8N::A6:dfV.W@DW8NfdSTSEL\W>A#.GO.O<UCG?702EX)HG[bB_fQ.;8=G<W+Nd
6:+(g\NaXMCCP\YgPaT[F-(1b1S41cdFN/X2,/gF))/IcQ>LTgIFR3OAF[.PfLHf
9,O-<VNgOAaQDQ)3gUa<_&+QE_aUP(Q=2+6]BJIEM^/+=ONe#Y:EW_OC-N]_6&f>
<O&1#AK5KIW]+f76L.4aKB)\P)+E-:WO(1EK/-3WB+9)OMNZKY&G.gO4S-ER2\=#
ZH+,f+[gRAQf3S+G,K3Q@B.=Y))L<VX>+;&+;acQ>gN=L@VQDVI#H.>IE4PUaOBa
I.=_#J+M3&BJ^SS^NB^E7H;e@;OB(Mc\LGN>Q))).E#1)fO->&P/6d:ef8&N(b;e
AZNTWE4=S+SUab49.BgOW+a)PSOZTS5DW0.R--NY-=][Ifd<^>G1UdABMT#54;g_
S1(U6VMK=gg2+72I+a2?-M\L[C<D0,,a:8aFFFfYe#E?D6?1?J]b7.@[FAGQ@b@6
gBUF/]7JJO4&1+WFEfTRLa.2b4WI9XC@5W\1J)\S<d_LAFV.9-&6QFZ=E7MQJ&U0
Yg4R/d2@)4P=(HY>1YIDB&IOK/UF/c+K]DOE>-&F95)22</EM&MICHefX0(FJK0,
dD]L3[/8:?gG92DgC<#PDA5([D8<JJ3/UJ)cICMETKN2--:0Q[8?F7TId;T4U:f>
4J&[cU96TNeLL^]419_Gd25_K4U)?,LQ+C&XM;Z\=NP;F.H+1M3^JG#?-NV)HZDR
QA=C47XP8)D(cJ#;3Z+W==fV>3M6AU9SBS-/+E;C6I-T#dD[VBIM[1QeL_3;USJ/
0ZX\FBLL88(d8dKPVTM+E:8cCWf6RI2cG35+O]cTPG=2&ILY4\>0A^I6^cUO5XJ,
HfH/f.)C&8<T_.9U8ZOa>IK]_<K0X:?b0S,R2.]-9>C0DaO9MWL,]B<(-/@=IL;Z
//^RZY[c4]8g^Eg\>g4ZK/dc&3&6U4Ef[bdDC8>DBJ0cWBX[SD/EPYQR:0W,HB)>
PTbTI1LL^GC89CH\D0U<5G_>LZAc?,?,WBU(?/,_O@7TRI\+_PNY?A)[KY-?EOa.
L4FfGNIUD0e/PFcR;YM2W,I[^CY6KL[\62Wa.a5MWE+WNMS98]>CBV/Y6g#(gV@O
bN;&Q5U^)DcA?N_ER3)I\dG-0d6ZB0dP[IHbYLU1cHEK?c-a,+G-/&+LXR@@FXX,
?;M4OX@A(,VL^c6bS;7@8de.c&(V^G@0[W^IVF8[RTb&=H#_;-K7G7e(B(_Ea;VQ
,aNJNIbC^9RSJ9O/E49,^]b[-V?-]aG,N6<_S1CZ1.33RNCSS)eUcS@C9VI+T4AA
WBZ=L+a.<(;2L1XL\>HM?(e?M,ecgB.8^JB<(ZXC]CH2IR00#S9@RGZa8fE1dE3W
YXgO^M[HOFW_;5SRb01[=2D7ZQ=T_Q^SGaW4MeN)7(O)Ga<SPa1G5bG<@ebE73AT
fB,)I)G_1JDM?@CS2DeMBZYZ[2AUVb?PR^RI^A#Y?M9fDP5>KZ)FCFU[V@1VPH7U
1RAg=Y7/I>bQ.XPC_^K#TV^TO>[H4ZZ0:)aO8<6\F?Z:+N^3,9Q:TZZB9\4Hf5De
R&7H?W>)V)CN[M<<I(Z;-g\cTfVY^[3e?.TH2=S(JO&K#GQ-b_YWK1^]^^bGV>Yf
(J):FC+>^8S2C,<#b0bY@-W&S#-(OCW1G#8=[5P5g)OCSDFYRg0J2[b)O3F..;;7
QK7O]XcL63e=Nbab#8S9FS:f(A3@Wd]8Ob#VXM4M9U-DY/3,YOaC.I;E]@IL=34G
&(3VJ&:(/fH>;#)1#>\PFbMU_Y4<;8V.K#?ePDMgVDU0ZYO&8\7#\L;0IL/Ub6>R
RKHc@M]Kb?:0<8BFS536-&1&)=GXW-XPP#\d5\BV.XGMRgc=@)Z>QJVC<G-a;.59
=TT5S7#LZFZf1_25U<b96W#.dQTXW]3#bQ03e#2<3HMQ.f5LG:?UBP>XaJ,TA-_#
I&Z)EF+EY9;:+#J#.P5_.d15OcLefVJPV\XU7eE<+X6M?V29:2aQRIZN5Tg]^?LG
W^>A-686R:b\6QFU060H:7;.0+<<Be1[XcUR+AHL)@9&>OW6M0VANSZe5:dg8&T^
KW#>IOg/Va&eO;OX@QScL.C([5QV:+B9QD?>R,2b?.\E=LMg\SV?S^.H,S18N,38
Y.]f]XLGR<eYOGA[;)9b1DV67^J5:H+W:MWVTT(K#@.=3/G4^/b+\>OVWS<DfTAB
F0:P;T,D7CO4O,;7D92\T&Db\_MX@g-DAGAa7\;2\\NJ.MbCGUCMF153U?=BWYfX
O_g(/cSL>IKTH.E@URO0a.K+TKHSP2MWX7F(8bF]46Fc2BA>VWH<]\>08G1Z4,O8
LCEYLf+Ib/WWL#-+IMPLU8dQ7TaE3HF+;TT#NOE\C;C[3+A+WGD8^B3(3,=LS4\A
-<gV;4\Z8CINcWZWB905HM)(M(O).TD/fK]PQRH/?VB5_\QHK1S,PX2UdT.cB[2,
]HK;T?VJGW[YO(&B.C5,+=)@/3(8BA<0Bd+<Fa<X-HLV1]M0Ae.b#\\/@S\O7ZfG
G-/a2@866g<==ZL#5R#W+Y-JWC1,)<8:f+36XeW1^RIAT>X0c_e;X@:0c>Q)Q..A
#WCee)DFaSd,[=0Q=Q\=CL6?#O&A]eMT^LK@1<VT)@a]W,ITGY@?5aN3Uac&H\1>
a/c/P(A\S&-T_:C:BV2\CMg,-4F&)M(H2]1M/0g7fA@7b[B0K)JZM?d6XWE8G=5J
0bYF&)TK><_2-8La<P4#G:T7>D0IV]If_#O(\LD;_F\X]b4#b84ZV09be]]1M-2[
\1ACXdKI\DJ)M\,KCR7QO\5<C7:b>(^^(dP>a++>(5Z50H=\0e;L4?;aEGKFOB(B
-=9/bPG_YX.fBIeKUK]:M(B1>O1@bZ\2,GPV[G\#I3bb?<)^ObY1F5<YXX:1d-_#
(TSN9f8P5WNG-;ZTWK_DDHGBa&JKID#2d[@UD6-H=aSPTX14D47c?4?g\.U=-,SX
eU)LOXGBXM12W8[7G-P7PLVG=G1:[\YYf-(.\J@,X#D;eg].?J-^/FaPRDV:FWKK
389;>b=N&7;:<=-TAOQ+2E]:L2BE?Q[A[]U^VYL[]8N_N-<d[gOJX#JQ3FS7W5I]
YEYOfbDHOADbZUSZ^&8^MH@PF5UTDf[Ka>)=VW0b?F@-KD=U0BI&X=9K-\^dW5E9
N,O5ddO(.<L(U_U<&\YH?L)McAA#<B2ac_-aN2VRGe8geJ8XN2K_JgEDC(:e#EM@
)S7:bEBD9J[TK6Uc8@-L;P>.RA[<adHDI3RKXH3(>\@A[(TV+NcQ[]1[#D]5MULZ
JZ0C>TT>Da>)GXIf&LLLX89V<G&4S=TMH(<+Y(gRZ_QU:-61TD3)ER/MHX/3^^<I
(]AQQ?.O7\LEH2Z(VH.fW.8M?+NQXe8]EC38O9^<KaBU1EQKa]XO^SV<^2e9[LCE
Yd3F0SIeOM5,(/gA=W-d8UT?5eT-G+HXJ48=G:>)C,OegSVF2=)N7a&D2J^8ZO\>
/Dg&CcC^^E+(S(V(-d5_;<7-1E-)c47]7@>-&:;061RZFOE,0+eM_0J&CeK<O3\?
a5+U5F<EIIY3:KAc\HTG-1N6R#ZKa.QfEGB-0HCY0<)YcQDZb1^8GSO;Q:\<5>NS
W1N1c(9?CO+T&JFg]B4YD,0b9RJg;+K7d:f&\;](Z#JaYE:>.DUgS<E+5XFC:b._
?/PBed2.RL(+O2P)\YW1OO7A6<RV0G_\1aZfJD9+>U;E#UU=^L,fE\YEV2F1aS7@
F@GL5:BRUX6U@Hef>d??\B)@+],8)+EB5_+\F2dV>GKEIA9D+N&:W/3e[+WZ,b?P
9a>(G+ba:@DL#b(cPD9AU#\N>3@RbHO2-IG3GS4AR4S.[RM]S,M3HGG4XN8C,SPT
BENd00<=+OJf+Z<+dU]XQ,08&eG_^^5-W\F@(G(Sc;8I=,)2FW.8O,eO3Y4dDZ4S
8L97]N#@09Z@-f9[W:.?;,W.-aUOCXQNDI<3AV+1(2P^@49:TcD8MZ-G-KefW^,a
=,gZ>;G.Lg3>a=)FG(4H1^4B4aKW:28GC-)cJ7KU?R(GXR.T9-V7#GA^VL3]@,>G
)/W>6].LGb6JSG#@ZN3?,dSA#-]BE7=9K:N[XN#;LTOd_6aS9<@TQKG]QaH4I[?b
Ed=2-CB6>LE-__9/X]bW.5e5HWE7UL=d\=&2;OP#\We4X[+OA/\B-^BFefW.67__
#67=<WNT9<)eKg@18f<gBEUJ,1,;[\:WBPbJB7B_L;O+F=cZK,^f)1_PN4)L3G=]
#^?;&Y_&,@T&=^-B@Cc[(^<fM:MUgEKZO]A;a)K2(.P5(Pd;@4C;S<Qd?YDa)_6d
^2:M_AWZ^-5R55YGG\cCQe(_D]/]?HH,V7=LA/Ua2;R05UR4321Q-/?U-7B6JUA0
@P3NaDY(:OGR&.CG3ZAWZMF7f,SQ@X-K@#+EX2.:H/JT^?b=]\Z6f?^HcZEc(#T;
#e&[LO]Sbe-9<HKbP=ddI@:((L4;W=<>TCVDTPQD;_dP4SUSQSJGXfZ1+5a]H8)F
,>fFgCR[bVPbHGWG&(>.GbOTRgD;>TKKcYc&aF[,,fC7O3_/R=RHUF?bUVWFYLCK
47?([a7A66I&JCFU.M/_Hd++3b\ACSRJJ)c(8SX)Df6:2]Fd(R9/[TcZ#MET\PeI
?^SW8/:E_:eV<7^.RIMHaMJ))H5@O)D9d;SfRX@9WO[:BYH&\VJSZ\4QW^B>4JV=
TXYV;]CTXLB.B)DCaD1eTR\;_U+a[S]A@1XdU\(--^7,JP@e,^8Qbb.XEPWdA,aY
b=W:P]T;K4+;Z&A>SW50:@0OfGR&6DQ?9>^b9?)-0LW_Y/O@?Z;9?H&LCS,.^25d
[#N:=QIW3:Lc@Q?fY[adM0(U[+bK4712aX[V41ENUQK,Nde=<a1O(^gSP=0Sc3@2
d2.&7?e:^IV(GCI+R?_QZeKAPVI;ec9Z6B6+A=HWJ5V878NcO8MYe&65;S7#bMD:
R65G&BRUSX^+;#K/H_e:W=V;GUHf/+c@E=USZKIJ(BU.;aZ_C_e.]Bg>TA]5g+HN
.2)WAHL;8+(2(Y-D<ZBWZI9@\QgO0>H7AacMc^dC+aA_d?JCJLfZ/PDadc(1XHN-
V:AGC]M#G_C&&d+^:0H8B\]OHe8P^/EK@))G-KMgK>g8AWeZeH\8+X-W@WUAHBU8
7G6)KQC[ZN^eS#1EI(->B>:e<,P_EW[0&+\=/DEP<V1YI[81G/X(BD(a@H[#6K;F
9@Y+@:V)b1(8Xd#=6;?;@J7^0e<A[TO-EeQ7:R,JQDM-.VMd4aU#Md4R1EG)>?EL
?=>-5F.,;MNG:<Aea:5(>c,NdT/CQLF?6aB6+2MYaSEC[R4T3Q8Z8YZZ8IeWS?I7
Ra6DdU)cYc<#JY5DY+ca43>X6aM>4bG4;<2S&_8:W#[(#]0ZL_1F/ZNGQP<ONL5P
@bf#NNB_C/W,K-?e=<]8U9,)QW#Hg41./__)TEQ?0RebO>DN]_a1:90KL6/WPKSD
-PPa./.BaSW4KJD0d04>XTPRdaLW,Q8[9@d)agNS[a,dPM0\VY0?cIP@,cN]0>PD
VB.TF+[U>\K^LI-7E3ZB?d:AJ\e6;+e+.G.(H[\QPRV+8[3,_(Xa6;a=Sc6BVfNZ
<;[A4(P.IXb_E@#8XD]&=]H99PL3B&NIL>_VCJa\bS<M&-,4VO/Q(N6((I]?6&+&
UN+e]]Me_0abC^JD>X@6@>BeKdAZeKYb\b_cZQ)3->I&W,<FIb:gW?g]_]UY]g<7
7=A@]7IO28IQZIMKK<>P:Q3e>^,A4g836b#CA1;&3e-MJSHg=JIDbNN(-I[QRaRP
K,Q2EA(_(,N6R#(g?D:PI7C]S]JJ>>\7<FI(FgA2ES9GJWb&&)_CQR(0Dg+V.8gC
G0-(AJ35(&&](,E;FO0XYRg@8BF)=0adAaD)Ae-dQI&,HD)(CSS:E9JXQ9+P@D,,
3d3J@_8<POH\M4P-f6R9_WK8QY51LQE5>=Z<)S,3ff109LP[cOV>)FQSXVTf>NM6
cF)NX-<&,O4R6^dWNSWC5]bO;QFBWSU5G[X?(V=@CVR4=L^A7dDG9X?#d]VBFe^)
R.LB8e_M7EFdBD>7b#4\M+d]D:C)BSC?E1K4PJ0TIN>DT[3,Pd:.c?>I<(4Z[-5E
64DRH)_7D8d&PYg]CK17?;=G8GAId?89X14DW<F#>-;aFQJOHI];KSI?3130a44Y
2:CUYM)D+,7^B7XSIc><B\N8EM-7X<AN2OB;EXSZ:2:S5Wc[3[bJUH/&YX6XF@\d
KFE.HIE>IV(g\_PJVKA7XKa<0bQ0F\g2LOYZ0fLS@<-6ZKbKHeJ.D^I)H^L+WP=c
N.V(B-:Q7NEWZE55/80>N7H]E7P<bH,P_J.eN@=]V;/+T5>-;72CV]@EdB#1XAJb
=Yea+\V@#>eMDgfP;),2I7NB(2BHa,B3+M?FG4ac-_/\5:ed,dEG8cX0[NYTH#]W
85d[4R2D2dZKM9,B#_:Y1YITb(SVMYX.c\G\.ZBLBbWG(MeWF<<7d[&OU6G63c8]
86]a:T@1P61W5<L1c3OUV8:A:D.P,(SMQ(TULX98?MPSXcLgLV2962ddMIG>@R3#
Z;>(.d9;K7C>>d)B\,/.>)=;bE<0)d01?\S#5/_J0M/SeY@9+SBdGI7OKcCMI9&1
6#NX<c;_8Ag>3E]/dTf)39)VTS\+a=455Ib6/^Eb:SW4AJ74#fS>@7g(d)adF(a-
cX0H3a1^891-WZE,:/&e]3?1<52G,:[-T)LTA(?A(24C+MY>)N4,1gV2U+S4\^)>
582_)[:(c<d4J6(2WL+UI<A7H>S5<,ENV(9[L&5\_VN03IL2P)_a.A\Sb=NE+Z]3
ONg;=f2d\4>=G.7[XG9Y?G45TJ1/[.f:KH^L:QA,UHC<(K(@]8AC9L=0XI/,1/X6
VBA.R-4.C,cP60[O\RV^LL++G^b;Hb,.N,&?,T=T??YDDM8[@^GT7EFG5(V4J(8<
Wa:HV]T[W/db19+(BRe9,@f/H_1?RPLU0e)I/cGM[9\3\Lg@0;OAHDBQW29-YXg.
VY>XM2J3TD4&^8BR)K^Se(-2GJO;5[N0+B9@KWgYg#BF[F[GFDeHD[92SQ:\BM<1
d_C:Xa\&d=&dI)..^J\^&gRYFbDQ:a>+:b-(1(HEYcVbZ4bJR/JD@&Fd[]C1KD-H
WbB&7>8PJ\R2T_(0;fJ:I7+=GCdgOQcI^=[W5<(LKLCM\N55H9S]D/D.?5_L<a?<
\fYU_Hb3Xgf\(-LE[ENNaE;:+))f+;K4PYQ<I51=VY-Af=Xa^,g8=64-bJB4#2-(
0+5X)c#:5C@)]?+I2&J^<,<AN;eUZQCd=3F]W&1-g;:B@&.g9],CQ+NKN]cE=Nf0
Ha.P-&;ROFa5@&C4=bZ^1&=&YO4cc5:cd\7R\H,Y9B1A[P-@:R1^CY8-Qf)NU<b,
#NEcg?>gU3+N0/5[TTY_fE)^?O-H/?:Q)MI(]+6_V&_63<R/I\7J5gWYQR8bS3_B
Kfa?ZA)-+&:;6Z,0K[,eT9.PKST-[EXO/U.-ZgPVfJ&=fcfH,(c(:6_PEdfg#>Z4
U:&#?QZ;>-\A&b_5]fb5OC0c)JMCY:_>:@&8VGg;4Za@aTLYJQ1AX^98V_C.7gQ>
7#4<F2&W3<[Ng9)(U/D??&:^UW88:JP[,PC>Z[R)&YBU2Y#F(4GO6LR;?_<]:0R2
NFA333VF(>#=S;DC,/gPeaGIba=0X/?48[,fU]QbA<5=I=eLVcV6/@935HWcOdDK
1Og(eI(SDJGN8:Z<c@6]Cd1SM49LaIN>79RE9_/40bg54I@/,MPLA]VBJ-6Nba/a
eCWB1@KQCBK\?T[P#(4eaI,OBJM&^]&/0257.3G0W0V=g8@,KPM[O/.+N2[6D0f+
Sc(.([3[1_6RbPQUUDSOeB.J/F)D3&__#C3f^HV9ZH/gX^8MC(LRcfSK]@[ON5::
0bI^Cd&Ufg6gL]/:6KU8+IO<=bKE/Q<[L.2W6K5H-X[U0LJ5#[@g(LbI=6gN+LN(
<QBfMV00Y4fQZ##bAQ@71@?<0R(fL4=3(?BR1&>I\1SXXH>.A,W;4B^3T)2]R=a_
VD9]P;/U:D[W\HG:I.2:6?RY/eD\^Z7gQ&9d/#f;HEKc&C0&f<=;EDSD+\R#7:VI
2:Z:]g4AY(ScMC&daUL/Uce?8X&QgUWG<N5FL&Z\:WXJ93.GWJ/^QKX\feb<FEOA
9^XPf5c=1Q9dB\51,=HUJZ)@T.L.;gE68K</8GU0<I&/\Za4@g5T8>46cL8F=SL2
(^<IfJg)>=)H9XEeO6<gf6G.N:E96-bIc<DI17W-+a+[dT=A05X^.-X?d.S:@+][
<D1T+;L+U-8_<BT8E6R#?d1G7>BcH04>638WdQ#12#RZ]G8OGfUY9&QF[+D66<GF
-XA\Z<I@+_L_16-aPSE2J_3d[8ZaJ5H07.N8NH7-:EOK)GD&J3H/0RbNYHM0G\,E
BLI,VRIV)G1TGB^A]f,^-eUF[FKFc#L;3X79FWVZAe,LLO,,?ZB>JJQ7?9M+FO=g
U?-DEM:94-7MIR:RHI_M+B,G+8(EL7?V_GG4b4&.W&=I;0Y+#ZbXaSN:\(XD^35G
\HFSJ#^U>:^S-0<c]9-cC>+@ROT1=F5\<cPa/0-]81N9\_>;E>_.DL_DYKV=0WUA
[U6a#\&4dg>1K(6e.+C14,WR1XK@5L\O7:S)3:[P6](-(T(cLC@I1LQeQ>Tc@:F5
01_+Jc-1+ZID)4>,IFYF,Q@NC;EYEB./&UPKMaeP0<I2B-B&ZadbP(YLJG(bbGE1
U]4W.76fg:=g1Y2)7&FQ\XJKWG._d-#GO+9?H>S[XHg8#_-T4[R^SbRC11_WG4Ce
[&5R33<>:YXS6[Z:Ag7C#;&G_R76fVSD@Z1YLb]eAYSC&L50M]A57>2J=e6+(T2c
^CC(SP#QXg,:,4OgaIa7F[U@E+7G;gJB03&-D#T#LEA2MdJ_NB,I3E)EbX^0\E<V
);bS;CK+QZ^9?#OEJX0(:>afGTWYQYB8(#=\R2[0CgH<I@1V>e0:8cA,5R;-KX\H
K58+J_<+UI5Gd::G&UY-VHZXAXJOAa2=6A&e80C1C^IV5?@8-#KB&ZW.1W+(UETb
+fD&2@V.[B@U1?f89+AVH4/ad1-N(..)FP610@5WNU[B8Y#7&;C.,E-^<MVZa4,;
SN(g0)R[H)>g,cg0@TV)NAd@43_)5,O]J),FJ[+D-JM\G42:R#gfJ-3K7=\O1Z6d
#,Y1=5;eg^f[<Y@91W?P=PDN<[1EJUHTLGN=H/PP1=K4aQe4fd7@^&]\;g+1^@UR
Y9L&Q#Y_0dL#[V][0N:GJL.1W5#RMCIQE[?dZaVg5TNd>MbPQ-WUCMdF1B^4H;c2
8-]DVEL=SW)N/NFO>U:,0FGY/90D.M5+8[;ZSI7Q9#TYS8P]gVZT@:HGRF6bK^L-
9KEg:TbMT^#S:VFJaH1=B7_7I3;fMMW#+B)],)cQ2IBL07O:)XL2gcLVTQO6Rg>&
/4?R_PU)DF>eNG/^2MOIM89YVTJG/BEB_+L6Ag]N<gKDa1Q#L+?BXQa4?9fd?^U1
4Fd;I,)M[3=LF\I<[HaDAZ.7S=#8#_)-1aI1QAKO<HXS.bYJO/bPW#b<_][9<X(0
XaSFS9/T,-Sa:+KH-U^gM_=GBT;]>Y/XCC2L.QF?[W0FQ=MQ)#_8B+D2@D>N=3=\
N81W2J[0[&VaW#TPUH=65-_D]I90DE4Q0U>5P/bgf^NQ,/WXKE(1,PBYP=9aZ\e+
_VPb+EV(>7cH,C[2FV:Od::#793FcG(_1_#G)_1JP&V+\4]#Z/<?dIW\D5-baFY&
6[dO-)&+\(Q]bTCHHI18\:6]?2^KJF&F3Z4(^-C4^)WJD-@aKXE:(2;9fc-<dKKB
T_Q)[)F-Aef1R6J(6Db9aNc?&-D4f66/?;WC-I21cI18_3D[6?5=e4NG@=NKSdW1
839:T2WP6<b\8MM#A7VM(B;Oa#_M&Z)FY3A5/#VIC@#I_B2MT_fUD7XeggAIZVcI
H?;B63B(N;I2Vb)fKF>_TBIGH9EK2d@&SMZ,X:W(6)VPE>e:,1Q-1D>JgHH3bO#Z
J03]XZaCR9W(3D:9_HNHABP&IR9SQ3Yc@;BUWZ:Zg.GU,36;^;Qd0&DCcf]AZ<f[
81<JG)3\S=_Sg_g^WH.E80-S&,?:]8H_\,]BM[bbM8=>FQE7M6BN61TNGQ>M(,76
T@(:AXWKII5Y(7f<@HIe,VN1HV_/6\Fa3EVDUHGP.4bFL+CgU-2]T_<U9V\EYGYS
<\JE34XdLLdVC_W)_.9K&4-SZNa1?DYMV4g/3_:_.S-f8><PA5?HI9?B#eQ,/-T<
V+LU<abM9C<af2[;QX/\0BSU[RdNERaED_L6A+[TSD7D[R(9;L<U\/cCB=5OH^bK
830CaZ-fEf8OQ@dI0eWI2>(6#7#dgU,FU;:Y^cISY22b+\X,=NEF<AZAPd#2G?O[
d:_>G@5V.FG?>62@cHEL4;+O#(]=UJdK.[/MDA.=f)O>8gT8_Cc4(8+JODDYRf66
Vd\_&PGZZ\_Z[/;0?62/#g?PM2bC=S&./>#GJGEa3^C8RS;ObY\DAEc^0ANB)(<H
B((]0MUA99W:gV/W,1:fE^7#&M5T\DZfZ[Vg6dE5_9P)YGMDLEHIZ+05Cb:QZV8-
7aCXAG0\6P0WY.?>Y:Qa-X\\eP,-SWgH0#)9I@SO3Mgc2(\0.QUBTZ3X#JO;(1P(
O.JLJ^:<g@LVHK?QL]75g-RBI^1ddA)S.M7bHPa#^,I-WYM--(&Tf]a=?(1d<??M
^EG1UY#/H-;[I#_32_-W.)E=GLYRe2Y/R\1]QI6+X#0ZJ&gQ]G/VLQ<.L9=@P):L
)Ne@[&Y<C?3.#Y3VAQ)WF#U<Cbf)?#N0R^U6K8W7RO&Ea;>Q:KUag+X13_^G3c:C
ET1<A-8V8+39e,>=>12Q)([Yb/ULZeA?PQU/M5N([gL)Rc7N4.=NdcWU#DCPd6J_
aYE(B3Hea72L#cMJ4&AH+WE)MBG6Z([<1;NgR4g3\?Z&S,)1=W/7XU4\K3\+bED4
=D561[8??2f6945TRSIEa4aeK=23&.;ce;IJ^4_Y-J+:CI54)f)\H^c)H(W0>FVd
80:/,17V=/Y9/M_OT-CdU=[:W&B)2]0a#G)I4)I4_Q#ZMEc?)E8B740,.O/2XJ5F
0gcX8KQN7ANHgSQ+_Q/XXAY_R_M=^MgWO04#>>7fBd0&6LMHd/V=:H^J6Z6?2A#)
.W57MC8/HAJXLU.W@TKVgB_ZMRc61IB(2Q[/O73X]7_JJHG0?-V;>>:R/JMIN^XG
Y82:DP^)^2T)?KBE6UK1DAW<-:\933FeL3BX.K/#gQB6eQ:,cM]d4SFc/He/8,0<
I36P3<#8EEB2OOS/93.6[d]:ZF\GG2AIgE^S6NPRfK+cW8IeJV(,JL:9L0^4#@&?
@Q[O\YgVYE)BFE^C-/bNXUCYXNgN[2#,:3HX?^O3)(KN^[fe0^4LIX/_^Tf)2GbI
E6c\TPD0F,:?Q#Bg?FeJ^BTbMOB+aRQGQY:(Ze3BA<FH#fXM/CW64^,>9dB.^:d:
\SYL2OM#?,ZB;#7.LGT3(.AfZ7ZfgGL^\60^OG26C:c7=IEK_B;64_+>,&+WC;+T
Q-1;,eX3JL\43YV&+10\eSIf#L#NY#FBc/,X4Q_FJ:)&H^5):M4O9/874VM3BWU\
3F#d#77/dA>LWKd5AJJ0^1;LVI^aDS5(OKKU&I1UHYVQYI2EU+W/@DCH675,/Y>g
e5\))&;6.WOROMBJ=5/>Y3ECD+AM7?BLdI#VR@U/RRTTN_0(W81,3XIER@a#[/Z^
#b&A4;G?O-TY#55CY0T],cGLPZW/PS-,O<Z#Vgf[dB,CIWECG^:Wg]OO]:>]PC9#
9])]/=)-1+<<95YM@>,7[bR56TX7c47G1Ba)TD[eA(;Y;&cPFGT/H,_eb#?MfRR7
)QdK7_A_G6RcA3YR>RX)#V//BQ.1E@Q@D9KBC;]5Q+R([gd_VO3fGTMIU.(DG@O)
Z[QDX79C&FACA12P2&EW\104g)8P-^;aDRIB1d269/CM7)]eAb8a[/5+9?d1_ZdO
J36X]WU68aK.#WKEZcT.05JJ7O(@HB@P,PG=XP0\E?[Yf(T,@Y3f[YX)54_H(I2g
K4=[\A,7LOLTAO&/Qa2R4UcA#NHIb0GRAT0;RRA?=.<^b29&d#,^TCG.K?2N<_Wf
7:3[5U4=GM<-G2C0TPA#?gL8gJ/b]^?]I4:SXFX<:ad/LK;6Ge4XQONQVS3=[01M
]9+/U7Af)#2J+>CNYPNPJAS9I7?S7d[\d8-[Q5SGJD/E44I2c^,aX;_ad[aVQ_dQ
WP,YD[.G7V_/)@7bNP<C=9V)1N2YHHV:OE,ZROQ6NGB/AK_[GLZE(RBc+;7<(_C5
RGJOd/SD]/4\4;[S,f]H1O#F?fWb[Wa/3^;R4:Y2^NIJ:eBU#a8=&6A)HL#+IcJ<
JbTKcGQ5=)@,A80^E.B;5+^XU/O]/U8aQ-CX(CeeI;.>MZcYW@HgQP)Pg)LX8]DR
D<PZQ??-JKJ8&_]]Y4>T@=0>d+@W\gSEIW,\:F?T(FBPWd.F(>3-4O?1U@:]VFe9
61;cbV+MD>P,cDD?+A7c_G(SBIc-,+\[;8CS&\XEKG)\GAbYNd<F:</APC.X4KM-
113:3XD_dP?J//GB^Ae_Wg[)_024\<PVe]F799d2TBL?Y3]Jd,8A>O4IPHGSOV_8
IZBKL[2MF\,d#>>BMRENB&YRf\S5Lc\1HbF.\eK?QeO7^52M&Ye=SU,GT_FRZC)J
IVO;=]WDOZ[.dgF.GJ0]T/]cVO[288@+O-Yg7Z[)dGGYKeNMFD1TgLO9DV)Pda(0
M+KYeI(dg+-Q28d7]9b^8Q1\dA6<C@QBf(FGZ42X)RTN>66L^KaJ-)ZGJ;+8SCQF
.)g/-f&X/(5g@#,8I,4DW1A?D2fFMSQ(fBHTfS#[]5+1&Yd:+aUZBaFNU+54<(IZ
^b^B.#?O)J5ELbfL#0;Ac7YI?V0SFd/NMH-I0Za[<?eF=VW+VV;_V3OMW]_cKUXf
[>e\,^ZXdZ__,bJP#f2g>VRP3NVf\USPD87;_1c;_UM63Z^K<A7[EMW3P@<\CMXK
&IO2?=C3AW1M<GfH4+N<FaU[L;_cU99(QeG?[4bb>Xe)LWM1K,B-&(/A2C/5b<aC
-<X3FHRSE\dBgZVf2J1+W1KTL;C5^:FVZV[Z<IEM\,MB.-@f(D7<YY_-:\/JJA9^
3:c<^7AQBJRcX[b]3[]c?G1cQE#X?Y-4Ve690HgA8SW0/DRA(?K+O6a/g/@UU<M<
S-RHN3B7XH57S8P4GEgUGI)9SX]MJ#XT(E10YV[A#)CT.GJERG&W,OgTa:O8c=7G
HB9cR=.Y@)0B=IYC;6e@a:/P#FRDV+;C4P(gT^=GaX@6C-@/<T[W_>JcV6,MT]a9
,XRK8=>/)-:_1R#CU)cKS3QQX2]CS#]A.AAc]/>-/WA6(@6CY/6&/7NO4M74=28[
HQR0b66F.46>#7I;Re^/Y?-C5/^?4gT9B+d5Pf[@]#?1Sa[/^6JJW+W-VTNcN67)
NV=?2Y//K5CV75aS.XBAXg;[[O]Bf:UCf,6eJG/P/>A=E3>cXF01;44>IZOe_28F
H..cND&D^&6=Q,f3;BgI+N#KDd6A+5M5C:-\6R.+DYX6K+g#=LGO-MBWOe:A<+KL
]Q8FSGa0:>>PWKME8C9L#>-22<e][)MIM]ZW&Hc<4=+g.TQYU\=-U?FcF1T47F/E
G4/.M>)<3Ec9J<bA7CEFTDKA@fT>+P(;(94X.^S1/^>aYH?D:TO1O?\5MS4:YVQY
35_IS85e)GW?Q0:W7,Hc)++?(a-Z_CgVF)d<V+,/2V::;Bac6:W=/28NF2d^+ZK7
>#W&,VKb?X-YRcYFYO;FA.?RG;c?15-&QI0\E;Q9@UK<d@.>WDJbf5>>=&.7aO,4
5QNWTLeK&=.C^We)3gNC4;&c=UVe,ON/C<b\5FLD-AH#b=H&A6fL2WMc,H:O\.7&
_g=@QQB,V-S?+25V4V0?\CM=Pe<&83^0W>7X46L1W](dU98;;1E<Mcc_KePJ<:^Y
SZdAOV=<I3ER(VC9O>FRC^>279]@P7^Y+_d,-4XVS(X0.<NUgQXZG29D@?9XN5,J
a2G,VUFK>Q4Sgd(FUN#@R1FX0BFIIeBFbW.R<QHP[[BHdcK4<Q@0FY\F1=W6H?,,
b5ACd&7eLX+bc?30L#Y(2]+=]T4#aaS:D#>EWd20,,/G7-+_\GZOE=?.SabM0UX\
]<B/F,@J4)YDcTJN50RIJA]2NR5&LM6D(P:JRLga4_f]PZ=2-9^OTc,&6TNVIJ.L
<]VVQ5TfUKG6RIXRJ=[E]@d?5NT)E:C8/PAcYFG,_2d2Yf^+Q<ReQ>a<4J&@]]c+
&[cfMC0)O^03/R+g:,?Ya97W;_]QU@V0G5Z_bA^OU>FU,M-E:T4=T]AN86gXMI+1
V3VJ(BQe>@G-5^XU:C.#JLE+,OaZB,/I)>;DdWUH[5Z?8^BK,15ZQREGW4L\)PT^
)g^gf;)//QJ\Ha;K?C):6,IWC+(&[+ARNMPc>&IPLSK(LX^H4Z)da7@.]LT2L7+f
.W?[P73Q/Jd_B=X>\AdUN6I<7>OIW56d@.2M7?gSeF/a6f]?)BI/[E1Y@5](@AD6
0B_S]9=&RM\5dVQ_K3EK]3c/3Z3:YeL>T(_:-;BEd_dB+:V?=gBg]V0R?>>:&FPJ
,aO^Pad17G4F>&NWGHfE_?(>>49O)ID(>?)1BJ#O#,(YbK;](-;=LTN;MBBaCXI<
2b=4eRF?<CdAMc/7()=b22f.>RO+Qb/b<X5&b96QLeD=fZaG@gES+ST)]W4,ABN.
;:-3.=6HSGS[OD<c(II01AQMBR_L[AfQK6FQ7\;B)M<Q2+91I^X]_8P_16UEI+@/
<;BbU_EI^16)-&]/YS]D(W\G69Z1E4R4)If+_Eg>f^c.ZT_+7?&4+?NL2=F:J8g5
9FR;X;;FEaa^6/\bF;2WS5IFZ,6(e;T^^[S@X4M395JZbEPVc>BdUG><F6eCJH7#
Mg:@<(EH2YEdPW3/c:(X2?9P+[<)4Tb@B<89HQRb6L?XKU:._#?4K&9TYM6cHNVR
Ug(P06M=^c[&NDY:V2370BDVBJAOEbNA_FO>ZOIbEY\>RY>M1g&3E\Y:1#2edAeR
OIUZH(daYY0)C.-U;?H)SH3^/Ub068]1I90+A/=]0(_P?XaMD]FdL47,?W0bED-\
;72O\fXBdDD&#<+F.=@@?.M#7KK\(,DeD,T,#MMQ[ca-?<]<cION]V8[3c(Pg7X:
(KF[e<a_L^R32&ESBcJ/5TAg@?]2Vb^ZA21-:::AP1>YA)W=Y@?;?WR5@GIU1ITG
)?DW6Sb9H[@-JNGTK_(94-P@RG>\.QG6,H(H@I7Cc(M2C\=83/XH[I0cJ)FS<dV3
<+;^0Fc<<-KD&a\:aAV4L9G=+=5VJ[1W&E(H?d6+27\((WRL2YSYW@]FI9&JR5L/
XTRTJ]5f>O,-M\ZdbYH;bH)O5]-[:>V0G,\=31>@T6)b&XC@^LG]&fH^9Y]>V8.X
(XBb+S/;)+()42P0\bJ/e>b@DHadC61<B0(HK^\V=2N0G6YQ,SLZOcC+R)I)U>fd
16bJO(aYeV:Mf@88H^BXD_S3bNI>D0Y4IKFJZP2Q3FO3=[CQ@V>A>()M@\W:cP4^
,^F#+R>^IK6K9>^b[XAX9Kd4ZVI_OZ0MR,_-OYb&S[&>V_.9]J\1aS)adY\,A5U?
gX#R,MF0<+dQC.Y3>:?/OF)0#(NP1QFU3gKcf;NHI#CHN/:aI.=0S;3)B5c_XSfY
IWbCRFI(dQ:+4#_,d2c)NC5+J^DPQA?VE\\ZdJY?&?]\7;^)8GEZ1Z0(3+>9e>BY
[\V2ES2E2aSHS^A6FRT?\DQN3S\A)RUDIRA5(E\[OC,DMZDP8I)W-O@c:\7T2<=<
Z2ZS,NGS-V)66M)1#3gGMf3>fDQ:+;[4G>4&6.S>MGK^YWUJD(5Y4VcAP=CU5L=:
9#X_0Ge3<Q[BA[P#:?CV3F[\[.V?c:TMVa#8&?3ON.K-ZA1\9>9ZgQM()QcSC@],
G)c#7N&+<;[F3&LWPDE8N:\VWH^)I&6b-2Q+^OBV)GP26O>90b#9a7CRgR:;<SP3
+@VNW3_,D6JWa6,-OQb(V_L44P,_#@(RYUH4-#9@8HKKJ7bLaI7gMV=)K<6](EeO
LDVUOcXUbISBd:_+3BVTTT(S?/H7_:_<@D/8R8U[1L4P#Na>dX=c]R4LAN]&(eCN
>dI2;1<O<3X.+CE0dD]#ga8gUUZ6HV2+>DTXD?PeT0G9R?LN46Cb-LaB0Ke1(4&(
P^Le;1d_Ib/V_WE<H];4;GOW18a]eYNTc=]_P/GCKgW43P=(]8D8;7=ZTc/T/.YU
-Zfg41KIF:H9=GN#=L+g>aJ9W^MD3-)60AJ>M&_Lb&J^1)7FF/S6PZ.M5e+^,U4Z
Mg,.VIgVIg+6CCSG<(,:3)RfVE=CV?6)Cb<TE?7MfB3Z,]#OBO,M[Lc.1QA)LgHL
16;XR.]E;F-6;.dd]d\eX^X.FW6P./FP5.Z\^+-H\F_EAK9C#=BE63\a2UIL@\50
<ORc01Q[NX</fDgZ2<46OURE#S6/OZUC03d2<>.RWcD??OVH92[0(+\,0gQ^?_07
#TONQca?W^NQg.La?9+BYX[<a+7\L\_UYZ,3O9#D&6JBQ8P#>_F..6fD-(Ce:ZH,
a5PTFaE[XK,GG4UZ:IJeeKJ+a<GKEFb;@@_d.+X^0OYdGOE&^;@=.7+5UePKWE,G
<2ORTE@U?\P@WBc&e=_P8;:&)PM_VeO/OLfJbLUIX)M^#2[Aab/>.a5PgTdF#_B_
:,^Z(.gBWCF0NKPP;4BL8DLd#c0/4=:P)L//\:aS/f9F?a2XSFKIVcRM2R48#H0S
WG2:gZ9<]FD1IK821cfUFSUBO^-6^@KLKYgJaCVFS=9()LOPRBaR<H&9JOZN]^GY
=1V+87._G7J0f9?NP98-L/eKbHQd4f5(1bJHW<8>BE[2ZI[,Ed0XWH(JZ,fA^WW8
3)[W0<E7]E2&B]c+B].WRSL#PZI:M_5JS7d=f<9PQHV9R8Z4S9GSZ_3>;MMQ1E_]
=20J#&SUTfe@-A3fNAC@3,HIJ8D9;@RaT;IT#ZNY3>_7.)<4-O[4C0NgCa;2_><2
I6YQT;gRY&H,H\-ZM:<0DAT4dX#SbE/4/?3?X=XAPE,W_[K#6&-ZGHfV;MeD#1R6
UQCE0gL;dHPNSR7MAME88]O,TAP[O=1\,8L=N<(,;b]Fc.[V\\2@=)/+EHU.1(5^
AS#9X_BEdB;[K335=&G8K.\C_XHWb=);b]b-04==H6P&bMf=.eaeNa=C8\JGG/9d
Z[G?&.K6+[b9RX=Q1CNANY>K^Q:S:1]1BF<:OCWYL[.:B4JRYQZC7=B9#VgPH^Y3
+UP-cK[HJd>G74NO_U#WAYcMdH6Z&2NRUN=0YMcAGM/O9T(XJB0PL3IQ(-66Bg7b
E9dNc3\G,3]V2I\>&Q6aJA;W9YUNJ;eKMI20@9^WA^IOC3f],:9LY.>0(T.6J7NS
5GHS3M/QBC&aIgD-gG.faC:YC>7\CS,[dTe=\?UAMBH;-fb\FGKNWEG;;&JI2gCf
>L(eY;WQ.ZS4=Q>P\9ZAd5Y^M\[,#\XgO)XV4bcR6Y#G/ddb6<6^;1M>G;[(b)H_
X..8YQe8bZL:KPCA-YJ&T&DP>^&T[BaX;Z-aHV2;dcgY?/UC4gRgaA(,/)HXA67^
CSUb#[.TO06H@6VUZPJ:M3JL[C5O4+aCF<UL(X\I78<,-RU.9O,4?X#T^V9c<WRD
7&_O4(9]EV1C<Md(Y@V^8F^2O?(72#[>9YdMC+QeV.P?NQ\LYTU8MU6B^UDPC5J,
HNf3NFZ))UP>B+cYcZK_6]d)dK-H\>]Y-DAU-R@O701S<7&NG(C(CQ,]Y,6V8L6C
d.U,7K#XI5U)WS]RL6Hg\KcFM\W+]BU)1VcD.e<G3/)DV<bQ(,KcVD+5;NQGY7J[
8_<>Z#ScQ>)f(BE2,W/;NLR5JE\U0A3R51OF=?Mc1c(CH:)]7dM(E[0:PbKccKIe
0P8XgDHd)^(cLE;F<bX?KB4B68)Z(VgdM1WH<FfXSG[Bd552]^E6J+eLUcUX/f_+
.TCDT(<#SYAEf54fa<OWCUCdJC[SD/EO.aGJ/?+CB9SY>0PJA0A=D)T0VV?&EZcD
;+c2I6[&aO_70C.;E;/8@[dK==G<3IZTHINM[cc>FWcS0PR]E/B5dgD0?c21c6=N
Od^V?M8,CZZ5MHLMH\VAZ/IT-Fg@8ZFU-0.MV/.0W9#TK1AKFTM\fYH4N,<:b]?(
aE8L29T-0F_Nc/_/G57O7[^FO0U&:-PID<g\,g61?a=f8=5(;2\0T.L92,+&2.3R
eH/(LN#XSEFLJP88<:OB:5WEafXbeMK2fITPIJ0(RZN.GJ:WS<KC(V619<eJ/4<Z
Oa.-V\RV.NTYLFZNGI,U3FJIcD2@/CWLBL=<XJPcWZCK\W,N<a3fe+A9g00.CX6L
T5&f5Q>MRJ(]:#Ac;<?3E]1d3W;EZM[PWY,eUJL(EH30Q9JeUIYdL;V#:/Y0-72#
>];<DU)QOM3OU#]BgT3;TG3d4eI7XN+.&UYBVC:NBD05#WX8M;Q&3c@H&QF^Jb2:
RZ?89Q256&b2Sc-0e5X=/JL-Qc^=;@]7/;@70K\\7DWSV[A&S>73G6(d#:2=RM/K
;H^G1Y:[14,6>9:.O.U=TaZf0>M0--I7S#6M,WcI(/U+T+ZJ&RI_&Db.W==d,<Z1
NJ=P@Ig+5d^NL4&8d7&<2>S)7C875UQ[&K>@#:2HMe\45,b\#b5RQPaEZQ?Y)F9,
U?_2#B6W?(M.b)X1]D0Y_fU4_@AHGZPMVfG0-[L,/T^;W>UHR-YR\\0=W2QSTV06
MGMD-eD3E+IXd+EC,K\L&L&\IX4CYWO^;+aR67]@GP/@1X=JELG\Q1T8^EV@J+13
JgXa;MQP(ZX5=)[Z2JBRV@YA.aR@:H&^a,#@YH9PG6.]P?;<@_H2C3KUC66VU18@
WffHeL_OH7R>8DDPc>Jf?H(?eU=RLF?51.[A[0D4;08\g:,Se-SegD6-9a3A8],T
:FXGR2(W@98a+4[TCYCP@f1B,VV.HVf)]N#U6,d#/\15Je56NXH&94T37X&D)>FG
3A);=P1QW)L@C1(,K;VNDS\,.@Z=AHME#4OBG;LR_U4?ILd9BMOD3XHI?/MY-J:Y
85-BYfM?QdG^1>;U7(/+d9BB:NS>ZCE5>e]_L#HWa4d-^L47R]LgGHR3+,]4L+OH
X7aLb3Y&^cN8c1bDQWGSYRg8J?)MR+/gV/Ife3)DfX2FDg@dVcU@WR6V&X.Z:SQH
=]3?0=.5a[aOaCQR66RXB--IS0UK5<6-PWII_@,9>HYD/&]5g,@,8;@0[];+38_V
V(/:)bNB<I;Cf46;T9[>.NFfR)eX?cHWA[+1=>;1LQR.-E2>5g9O,IE?:MXH?fLD
K>^dC\c5-H_eRJPBYaWK.5(68bTT^FRY.>V^P,5S2V7)LaVa8Sf9;[VNV@=;cJ8/
e?RY:=X=<QC^]7,#cF/JST(7Z18MR\:6A7Yf0KA>9D)QT/&3IFKBGEf5_d#N:@=I
ebBZU<d8VWP47DPb(KafEVN-JM<[&X\;K3>^b9Sb=eQG.bJ2884b76[JQ0&f#c:=
cS6XS5aV3VL#J/KWaF4YZ;+M?^WA_;)68?YP(+>b&(62QPX=aNRZIRVUa#+KNb&1
cD(_]0d6,TVEB86&NWL/G+E<4;KA2[4U>CH>ff_e+@72RK_01V+DFPaI8f]@@Iea
aH20X7:?RZL/H#/=MPI0)4Gg0R288<<^a@6(5NPSK\F5([L_7YSf2CW@C@W2+D=c
Y,/bCf;M\SNOH)N&P^)?PFFd=Z#G.;+F-XC&OD0?W4#fDQTEP4d7c>Z@28#edPZ=
D+9#-0EHa,5c99_8/E6c#P#WGVf/XHg3V?ILSAQ<<_:E&NES\0#CN:8OA(-RK7BR
aBEM0POLXgd^gN)QHOfROW&138LB56(Da48<Xa<IVdT+b=8aO#1(4N?2Q78;)Jd8
?R;FAN?,3cF1@N2C81:e1Q.Dd7EaAa0N3085^T#C+C6\Z&8U^&M@Ae]Z34b2^/7f
-V^ER2CH5,M1/3R\79=/dAcUR.:IT4+F7<Hdg[K.3Dd39TeW8/[36.3QA,P)(@+W
DcH>?E?=g,bK4_2<G^83-7)1RQGWOZc.,84JVPaXFRHPJ3#;O,N;^JX?:e1\MUXf
eA6BVLZ<&F5@;,@G&[)6\>HGA9feT#0B7K]OH@bKXU<VU-+5]N^U@+(H7cUEH)(.
-J6MT)5+YQbH-T&be(JGL-G9K:]/LQ[:.&XRIV]G.g5XdOdfNM+QV72^]2Jc3PBI
1DSQV_GgfR^X=I\c:=^TLL(\#4KKOFK#[SD<(Xc<E?;:F5EU./]d8];B5><(HWY+
RSL?3@>RGH?Q6YKddP^f076MK-S8Cb[9K4B.[D7]RHFEGVG/UVG9GULRPOZ7fAMP
-LN3?,FCVUM#0)22g73fJ[(\N08/>Z#.E[G4-+Lc^6D_[Z)FS]]b>XfU=AX[RHR@
HFUBe+,X>@Z-NUL,GbV1:0OW]G>26TPT:I,ebVJ[RJ^PG1@eG^RU@52TCb7dO_-/
L4KJ1VXa5f//H.H9>,G@S4-?^J_9>Ce/GbT9cB\Xf[&T;\Q[8=B/W:+@=)EZ60F(
WSVEH_d6=NH:;DP1T,GETbHWE7G1(+LK;eC-?fBYPHRT@?R:g45=\f()FH#HP_Hg
?YTC=L0Jfg_?>[<Pe)Q^?f-I5d3c@VW,C89JbaeM0KRSS\>H4eOR-A;WV]YG&03-
XN1aE-V]-JRQWR#L3OXWB6Ob]Jd8@+;=T+@<IO]Z@THCBCTBUO#Q22MB[]//18R&
Q)-#OG[>\f-\4C[B6eX#2RYZA36U&ZA.eKY<>EfE8D,8c-DA[-NHR?g/KBI86^:D
I3<L;PRc(K(1WI,dg[?E3e^I6M3M3S8E2F,]FRLgA()d:GeF7?AI=.aG7<CNRGc#
U_,a]C1JI1-&c3\bTe8a^E))-(e2#1+&d>_\U_5CKY,LWF8W<.=?^a:BXFTF.eL7
@aYCa:T]VDBJ_>0CW\+[(1G/73=8B0-R8T.L@H1fG53A>>d8=.Q1a9QXV/S-7R^8
=8\;6>;[LNb:NXN1.5=Gc-V6@5L<Gc(^WFDRE=9-^Y[2,Q_DeTOP1S09a/SPA#\B
De.QZP^^UYEAE7+1X#4Z(6IZ6=B(&PRI5C8@>,CJ_g:L#f3Y:E[B_VHZN^C6I;Vg
I;/S.3(H#3ZEA+N<N41IedIfgAMg^T++0O&bYBb[2F-.AfBK+a>M9>6.XV_=a@#R
)Y-7f7<4YZT@SC=e4gb4d7AM0Md9CBB84^IT-;99PG,[85+:\5c74aR[8;&J.#&I
@;Qa1A;^3WOVGM(Z1e5cS2\W&T3WGX,Pa-<\Q#A19/41EW5Y9R3?f.gW@B>15G,O
8G+DCI@e;:ET5G=H2ZfF5b22K/WDGI:MeVE&K;T,A.@D1@^.HLJ4XV2aK@YWQc&4
f-P99>e^X4LP[Y4XT4IWJ_C]-3/(g;84&.Ha#E+B6FAMgEEB(AX_7UW5JJ/bb:)V
?0^[W/cV@N?=)GdGbScfZYQU6P,<f8EPFYGFa08<RG-Y-c1X^<)KWA+@:L#eV;N.
A+.?^US,1\U#G)#1UD.bQT-?3)fM^QPQ.N0R@]-/]9Z5U^SCP\1KaUNed==HQI@D
N#:^)>&@2&7F?C39HYENA+4Ed<Ba[&&JfU,M>gLf:LDL.=:JDN:[T_4WeN[HT#2D
)5L=U#EH?O@-BJ()bA#]9YIIS(_<cJ(e=Ag#UMD5BA@NE=H[RA<LTQ#-_Y_1;SEG
]VCGNLJe@2&=8.3MO1)::,2.7R4TdeX>;DKd77EKLOLTQBNd_30A4&]1>YJ9B[K8
CZ]D,@70cEeAGGO:LHgX.\Q@>+bc&+?@52H/WN(=5&,09272]daUgPET]UO.D>11
BZ2V6:(05[HQO7P/9FPP3?[\6-FM5f]4SR[I5aHDeb=C#FFZMU.D:60N7K7+X5gM
P9VN/dA/.8PBLTG?D\W/D1UZY+Nd4X0ICH[Mf0FCHdW;aZgA/d1I=J.MLP9bGZ&4
g.51F/VgVd&Wb<.[V<CT,+CBeD@J;UGD5X/;DRF2[-S1Ae]GRHFQ1V0X;\C,@?8S
(0;63;e5#Ic;AW82.K_cQCVWJ[dL:YgCMR<LASFO3e-GB382c3L-Nf^Q/K)&WW]M
&M5Re))KL/;A_5CDQ3@MKBMaFe=S0KbZ51YG8G51[a&K6U_<.JW;AA,H[=]NQS&G
c2?U7>GJ/cU+PO>0P70V@)HAL/RdGZEM8=J8A39LQ+YfMU[[,#Z5S.,(XU0(?O>9
D68B(1,TV7-;?.D:IFH7#9XgVZDIXE9X;ZB(cZ1LC(M()gLT@GNg8XC.^);Q?6?3
AQaH7&C@gFH41Jb#/2@2XI30]Fb2La_Y?7D_.YRZ[;QDb78XC;KS?O7&g3P^GGDf
]3eg#dY5.CFM;,EV>C\@ACE7FT9ZKXR^W\/X(=;#A5DY</;3Y0HYJ/G4f9;TJ>U1
+:#R&>gBPI<)KI>a<Ne\J693OBQBI3X9-#[VW4YC++-4:<g7=3BSY3cLJb^@ePF=
A.BURd.4VP<J.WeUC3FPLVCH4_JbbXKORR4.&C>LB:>J70GTCe+5)DP-4a(=XKf+
D0G0-2dd^AgIeFcJ.-Td;)QI7(MBG(Q5Y?JYa\6eN(Q#g(FaID=2.R#F5aI?AT+O
fX9#.V1];(<A1].=GCMA-N)LCUe,DAAFM[DT7&cEW7:Y0KRK_I]@M..\\Y7XT@X+
#+?FXFS+ENLM)a9f\]@&CIH6@e.IE#J5;>S40C_61,H6XF/@G\#2=_;(O(TH?.(-
ge)d,9\&gS/YXN>S-M5YE@D90@[SB)fR+H2Q:[H<^;,4FGDS1:\^;=JX6eLc\E0T
7>A+\&/cM_),S&.PPX60+DT[LTYRE(&gb6aa#YObdL23cK(M=MAcW_&MUGA+VaZ\
P0fAZKS8gdMFI(.(5W6+bgZ(D7aWL^>4f+H2QUb:4^Vb./NWQL1fE[SXI?@([?Ac
4DQK/f:g8F1##S6Q4YU8EMP^Ja^AP9BVc3LJ=K89c17W\X15XB(e:WOcCdC.4>5=
L7NK5S60fLgMceUX^M]Z+?Z>V5BYPRP1I(XeF?:8^B;.U]J0[C>=PgFYL<13[N5X
aC0:AW[@6#CSQ@9G/G1D)cR5b]Y1HKE@E<^Y3PbNNMAK@B?_C=[(EX;eAD?X-DgA
+_.IcEV#V84]/XL@.&W\GJFRfUcXQ<59F+<[CQTH+a-L57_D>9VDBH=^ILHcSHX6
=O:30fH6Q,]_c>Z&H?G0JU+,+C&).37)FLWG9b8<[3f#6Oc0=#7+2LIP?^,)2bS-
fEg^0B[<Z4_?YR3R#WBUALfO8OD;07O2=H4A0A&T;;;?5ed>;)E5O,9>R73E]C(#
ON8W0C1(:(gRQ49Y\T,.dT#13M4L?I+0B^+^a)]e-Ng&?E:c<7AJ[e:D^[=caH/7
3DC&E(dA;c(]]WVX@R-6KI:?99A0RG\(geWW41c/N#A(c]&?<K\9:.]QbMS[Q7DI
9425O<^-6aV;GbXZJH\V6:fbTII?Q\>9+?#LB2A^S7I.AGGF;W8;)g7Qgde+YHTP
_3WNgAaH6/dZ-;6?53\K;a6b[@e-4;a)5N..#KJ\C)6IW^5gdR]PYWc2d9_Egg4#
.3_XWIA:fN-:c#\#G6S\F.2J(EM+H946HS.eca,3&52OJ7NFW[@1DLK=bfb9_4==
@/Id=\_;#K2:QS;)8<^a\ZVF9QKY._dUSQ)@GYWH/L67M]bTWDP.D0/X3W5[_VSG
Og:;_&<?\SgdMIP3RKgQSf,WSLPN+IMI=RS^07[P;g?^&#2V2ZF\40RI\JX7?@Q?
J;-L\K;?PNGSMWC+eQ]GdU&4A5G5ZAT1CI2]44aWJHa3]F\WQP#G/Q?HWNRWZPS)
ZC5G#82Q-[]^beKe&,T;7<]J[?F&TOHMQNLe(3\7254S?L,+cEN-6(NNR9Z^g<V/
gB]SLZ<+7b+^8EXb1^D)N&;D:XLD>a9a@[-[\1\fF&^?dTY/QCSBSN>&b]6=[f?#
@I_OS:f]b1&R<\W?]OLM/<g+N4dgdP08Z&/=OZ([7g>cZ?R^,^a;@M:AE:)K7BD+
S3-6/gTg&./Ifa63PIcQf.-Zf#OgIL??]T2<^fb@PPMUL?=Gf)Z>-:4W[XBSJW6-
2EQ6L?dYS0G&XNI\6C<SGTE?36^>Rg8K-:c[NV^b_U)\EXV]a1+f?A\>G(Q_,_f/
9PJ1-gaJNWG7aU#Fa>0<0,cMa:L5)^Rd]F,TC3Ge=W7dTEWM&32_[B1Ka[QTTTS7
KNc07\^e_6I2&9C/WP2ZMYX3-OKW@QYZd^<:QW3VS;HJR+U41-:)\)^1BcG[LDKX
+6NO/Q-+6]MW-UW0QC-JLA3O-9I5G)T_Y4bB:DHS.VMH-BSOWfgE22d?EQa4D;=^
2E#/B&+LMa^g]-4ag;B)B[&I;#d_0LP5/[F\Sb:<IM@G)GEg=,UZE19@ac<R77,7
Jf&3X7;BWVcD8:DJ_-H9(BOg_]D-GCDK+Z.d/@+.KUag;K6OR(d7D-[<-g?L-cZ,
7([cS##ZU1[.)-ba3L.^EHLb_8T93A3g&P5.FbLg+f9-@,QHdTBDRa1d,1<=W5SS
.D-P>26FI-[3]P+H4IG40Q8PfKEb.&Ib:JaZ,W7eL00Ba<EE\g5RQ>67/D0)d2<e
4S]JZ645#>=<J&\:/@SaW>\>/6]d,MagRIGZLOafA.7&&HLIT#]DfQG^LOA]_7cF
Z[.-4Z]&f,E_L\O<Z7bG\,YNEJ4#YX5ePOb))JF(VPfWgf[U6=#P6bNVaWaKD.[A
eH\PB52d#]HYH^LD:5.MVW7BV)PD_7R7WP/:/#-cIG?169[T>V,EF1T\NIY^]K5^
YH1/0#^GF@NJYa:@;?Y^5[K/Y3eXbg[3fHAY,,c(O3,=,UaZaRJZP0Q\+5I4+Mac
;7E6PZ+^.Xf+AOBS7S@__PS+W\I(1OQUa37<GbS8MWB+K]/YEIFY_I;&^OH7-(T?
N.J5]3#D#^W1X+3M[Re7e5XFdC>-:<dO5\&+1?LKZT]X.DMNRXf\Z#DM(FUGM]6;
764V\[D-LUD^-&JM)?4&SPF#bY<@dM#2N+&-FNfRWI_:M4?M?Oe1R@5=/Y=UJ]e;
A9WX@Aa;T([=fL#0I5/7R7XW997LYJ4_&OOV):U#;1G.M]1BV7>&+7HeP4+KaQ@Y
DNYZX>3Tf.C&7XUaOd&-aZ28GJKc79?C7S.5K)N9[fgP#aX)4UBE[YOR()5VKCHO
T]W>)U-X<]/d9<_6TfMXJ6Hg=I38]/b3+Z9^Ka5+1,/_-AD@Xab;Bg?N+VO]e=>Z
=1EFBZ5IKDcg2#Xc2&1<U+O=H(ULA]#-MIDD;V5)b\PeWA=4=5J0ZXZ19c\#=6/;
#.[JC?-,D?UPa2&/4a,NMIF<&H:[aH[G;,>6H;E7=K&00KF?K6D9EJLUC7IXE3M&
4>fD8d_(S^f?VMGR04_?U8ZWY756972@&Ice@PDJ#;.2WT9ZbA@8Pb<Me=VfHP]T
:Q;W_-+RW9cR-SC/WGGf\,4+J(/;;))RA;f]9-Vb5)LS_>GFL#VNF/RSD7DV)f60
MgK?#g;6f)8WLf(EEOac4g@C5/=E9)8_O\g;[8=L_[_UM&(ZZ&U0?S2/:O)g1E\Q
4U#894LdX^F\XOP^=2eY?8POOV530AgZ,51_@E,Z#@bHR(S4J5(eQe,^VObW0b8I
RA9(=3__RN.2NAXg8;>I<HSL8_>(;Ng7:YOaB.NUV&49L4cggHd8(fIM6W0?O)J@
cdE+?f/JX0+fV2g2(@dc:7&-(&_-I..3bJ8?8?NE>Ba3(\E&L>X2AD,Z&S3)GBMS
CfNbF&eVb9VeDI+Sc?8@a]+1XE_=;TFUf=E?4\1:4cDa<\:HMQ(^<d0NTAR_V6b<
B7GP@ANJH>PEVZ]QFU1[4.TeZccb]NNCTe]QK2MQa(EIM5ZDZS<UgaW52f;a5BJG
9BX4ZR=c5.5fXU<TM.D4EFTe.KDN&5NaSDf7HK+X;[O2UDO3.f7;C#P/FV<M^.FY
ZO?4:LNRH;3^<N-GX&?XT.#5,M:QY=J(J6[SbP/YRc@_W\4TPZaW4?a?M)bY1XL>
e_b9OFF\[EC^AJc)IdVFYLa<Ad[HF&,7g#[HEQ8-NRd(),-X/[WAQ_Ze7]:dK9(Y
8#Y?==@G[K@a/e7R=Ef5ZGZ5I.Y13DNE@XGG@e7,PeRE#cgA+ONJ5P[[M0YGI?@2
6Z3D-?aJ=)&^78[(U(\XR4QN-66bG[U3Zgc@^>>YMIfOG9SETKIB914JW:?(b0R[
V2JPd)HZ0DUQSM6>g.H]SRD:L<IQ3,;+Q6?QFXHbC.1&U[2a@2[bC:MegFO9[.\]
89P(;#QNL.b?/E@/1J1YAI&U4e<9[QcZb6@]Q9]&N:].KVSAQV&WgDW6c#3a@16f
AV^=YS-Q91E0OdUGc&Q7#R#8;?UJPGQEIEI\Z]S6G.J6+a+#O1M;F_WeG,YY;>bP
-C+_,CaIZ;+LTW:8FYFM:fDbE&[JF/7.]UR8\Z4TcAD=&J046b+6f,M^f_N,2OHD
97Cg=T3(C(JMG_;S61Q)d?OeS9)12SC.ZgKD2eX/NW/;OgJH-g1GaR?VH8-VA1AJ
N<CMe2@P_X.KDF6[TT1fYbV56O+0D\eNSe_K:ff6C8QXH2@OR-APZ,aURc,HFBg(
AZSRcX#BIGI;1;;#+TLA(Kf6gfS-R>YIK.+(:>2WNZ+R]VdU>>7O=5\TS1#,0LM1
Q+Y=>>-YN4cOERES:KOYaR?:G];#gWa/,GgCfX,S8Y:+^W+.?Ta,>_NW[U6&TRJf
]4;F^+c55cDa=HB(82]@WOY=#FU+YH_CUCaRDa>J9\Ee.)UXIA0agZgB#aS7(?cB
-F:.+R85^QMB7PR2>(35bZDBN@_E6)U+[)CA4R;M+bN.=M-,Og0O2(XL+W&Qb:_\
16gH[^UU].)JdJfGNQDPG46ca.0(K7,I7BDG1&Ud[TSb-Z.c;ef.>VKX?NZd[P)X
Wbc>UMfS91L5W.fKa^befRgPd+TJ>?ALMH7N@XIQa(8QT0KP4.P_.N\OJSB(FPV\
3P<Kd0R>C>ABeLDW;fTPA_TPebUAE_);0CI[C7P]<?R<a#-@;beZRfV&]\HaK;>[
BWafQN_0Q@M-dZ.IIQ7EO)^9^SacA.fPOB2CT>d;7INJ_WgAJ3XED.C5)a/PaO96
9fT?)4/+?SPG+PXNcEJU4L.Wd).Mf7T)I;Ac(WOCZ(fK75O]e(1<^>S.e60d/@fP
<cU_;7G8[dMZ[cb.>2]fAf]1Y/75M+<KSLE31U,U<(_PNTH4d-.&_XR2LT,@A#]A
3@=])_B+>:Q)]eaW5Q/a,2Fd&(8L.]&GFH^(1]WMM0d5f51:S:MH^8V=)<OJ-eCd
HXO=#OT;WZVB5++1@7[^D+aVEFgB;:G6DU5\ObU=SZ_EgZ]PYa\6&[RdUdKG/V19
WGM?SO,?Q.3Y>TcNfa;EgEI_<[L/I:L/-Y9YCL@T#(O/?;X&C\J(5V=XNcC<bVVV
N[9M/(A03L6KVE[7:.[HBYNEI2YO1E)5(]aFCE(RX.bDf=4R>a9b[99TQVIM^K=,
OQR=Y6GfOQ[&L:>]O;_f?,+8<SbX.NR4b,g3.73)0AH7.3^.&,O42e61&>50/=^A
U011M#df9.K10TS6>RLe:6/VPaSL]MTYMfa@g7Oc3KR=:SBEUg^N^:>N+8b0,IP/
Q:4:IV_]E=MDJLWR@]X;W1U^<IGA2@TC1)GRZ+X[ZQJQS=PJ27SF[MW\D813+?[1
P?65T@T27WgME@@d#3WO\V#7MF=EK.;S-VSf-Y/<B8AFEC(c+RT>(_cRSWNaC.NS
;85C/bM]_b//.Y,Mf7.^&=B\UAA9,;#,cWXHPf@^AN)LBS;,NUSUcS#NN:[#We]5
M()R&R_cQ^32;Od&=WIgF]6V559g;g&eQW2)R?Y1FaBP0#6N?\;XfYR6bBRPDc.&
1[e04XFX@bH[.:&_#[V15X2QT6CNdC#O<)#&bK+)ERbdLadC0Re\-Fe]CH8+N^[8
0CbdW95;].22D+I(&b0fE<I).2&2@XR.[NI3CD)b\<b3W^+,@:L_]^H\aSSCaJ-]
=,)>^0P#VM11-7?b]2XX7\6N)4XXS[>:<1VT?B0:JBE4\?2PKFRF0[MU8e#5IA3M
aJX4S6_d(B0Y]F53f2,)M2/Jc.e>6L?+/?+#)7(:,af[6V)I(Y)c>7-UVdHWKIRV
QXO4LPG_dWW32])/(7I9-7fEYMA0R(29DE9>[WTB78;;ZGQMSG<@SZ>\d/,B\4Z(
<N[K9)5].Sa?aWg><]/UeQ2_/EVUW-&8<=68:c5MLW;5f0U#>7FZG7V8cLfVf&S7
BcS=9X#68DNWLK@HAg+3V]b3XcgH>>eYT(GK=4O5_E]J7FQA]a;BfO=ZP\=8I\)S
4SF((BA8)I^FUd^K+cQ,\81-;>g]5F\<NS2BS/-.&d2;MI)\L(?g3M,&Tf0@UcA@
g\^&6]BO-(2B\f/J9R1I1\^(<:cO.,dL5R4IJ17#\Wc&=QWNeQ@[Aa46aL,POg=Q
+_?8@:CD7L?MfN]J4L9-g5MN24Ja@_a9VXc6G53S_3Y+G.E]TNW+334]HUd^CADP
7Z]FI)2Y5B@+_-cBXPD\@THDYFM(NHZGD+]TEaV_dLeNg0&d=#Tb3RW@129[D=:C
]U[-CbT>_d,-ef(W(Ge&-)[_bXgXA@97:NB:C-=S,QG.TKbZ/X8a@\O-0f^SZ;aB
fgR7A>8VM5C7U=YLO3MZ/:&b4Cb&BKDSJFYUIN=DSU.6=:5WKUCVL(.Y+A\\X^FW
]I8ZCT1A>b)^9.8U\Ic3Z8Lb-]c&Sd)Zf,)f3XR,GH7AdO9>190A<WJgS[:J61T;
dgD#^-O4GeANa5FP7[^8LLO>:\XBE=N7Fbedc[+Agb2E_R@\1K:&C?RA(VSAf4F7
SfTOI\J64a[CQX?W12C67SRY40]AOLC@eE._ZEE&E9ZSF+/L0(ECX76YGS/QAL)1
NWN-BA]Y.QRc+S2F/7NRF)UT@?cPSagQRgIRKI?&c;CSg-@D,5\aD<OE+e#<[CYE
XZ])2;T+aSa;ga?5E?VX>Y?_\#^NLN6:UKW,S/AGE^L9#_]fB-\I=1GIN=J\[F@]
4>GP3DGCLD)\@1\2TV5M9<3#Zc:W1^A[8S^P<UAb?@#KB\H8?>3SSM6df;6PS17X
R@)Pa.c?GY1>M><(;;Zd9Nf<4f+JdG9Z^CD234]D+)=/=fOF>f=R[.P1HbE7<\FI
6VOSU9-\2PN].;Z@6/U/fLE[3fO@dVd8f=5N(T8._B8T&WV5&1\)c,Rd]]_OW7##
-O&X^aXHOSW4KU.aOd53c104C1[Ig[=ePM9XfA-6J96eL<.2\F_I;X+A:Z9&>JIf
[&-;?CVe.Cb+C\G781(68M^K@g4)M(3I=7VH2b(XL]33,A^.SU:+BY<_B<5X^J<6
b(ALVLV2.,1.ZM>Z7UGMMLa6H)ZPTJ.[N28V9FI&\Ea4:[:aHG4-OQ;T>ES4e56T
/?<9O>]cPYVLf1B3=NDYaRCG[Y8@HP&A+20:=dAH):&aJ-MY)c>W]8_S=3MT=:48
_1<fQP#N(/2a4Y(GPF=H</T=;8(<+-f6(ESUGOdeO@BW96HDgcZ94#3dd,6OfL:P
dK62I?aBD[,1K6_6,P8/d)<=G/2N>J]fcJ]_^(&-(+MHN[>(I_aO;XZEO/,7LY])
(Y,4ETgPI?,^VM(FXXJ]:GKV3KK@,Y)<D]54DAU+34gQ/(<SQ:RO6HT_2edB85=V
(.;N.))b,-d#g30Lc7dW].VA]ee8UNdI3cJS]4Ka&5]^2F6c&NLOH/IP]JHK0-aP
8d<&6T#Q>]6)F2S4Ye[[c;1HUO<K2KOTHC6GX?>2_W?OKabA&Z&/QM2DC?ab5T2B
>WMNJMec2XXQ6aQML^E9:144O.==Ga-,3V>3B7T&U?,3+:5RHE_g_f4YOd,[^N6S
4@fTL6C?[.)8^XgQ#Vb\XKb[2N@CQ??5/d:\5Xe,WMTMb<(K^SF]N5VR,AD6f+dO
QZ;&=7b9USaWg&).-_ZG\PbgO[=KAb(a1XVag<5WUV7D&S[5[S,JXPXU4c1YgdZK
dVg2<c3<D5V(V5:6,JOH3;RG,1L=-V?<F5\DaY:,\(WB4e)5^D+E@V\+fN1SCR0c
73Z#?:-?;eXCTX<+9BZ(gH:BLX1MbfFQ#H5O/c1MBSN;Ve=c^HR+1&@1B;4[EP=I
H>Jc:R+<6H/Y=bd\(J:PKG0M+H_RLE([#E;13@GKX_OUMa&J(P.7#O<=96fACCFJ
Pce_1LOA#cA])/]F.5c46M75_JG:6dI=aG?.AHG<[_&D\;PQO>O@\]/\_cN/Xb2K
A+:G[0R)/g9EgZ.;=b<SZ=@D;8DZHI-aK6M(]FXEYQb9OSAJ:DC=<]R)+fIK_dU^
PWWgc08cJUOQ)>#O;>)U.]7AO>gaa</-26>JP2K>=\8-S6=+CIHUY81TMM=Z#(M0
5EJdBHD</T8e-AQQcg<3?P.d@<W7PgW2-4]&8S<HO)SX\Y<&X?>9^)>6f/#KReY?
7fOe7,XC:bF[TgL5Q@AHOKXI(D^05Z[_1:Q^6RBGdTT@SNT[=0AORCcBNS633(Je
_,1,bWVb]QbY\:0Df_5PYYMF1L+c09KI+[RVRZNZBX?c]ZJVIR@#_VLJ^fPS=OOB
WJ&R+V_=Q:JI>8N9^(IU^U<:TRLMAdB>\S(1W-#7@,cYf:d&QB0f\Xg#V9#AHV]T
Z)KY5df)#,O+@[G?]4BC,.>f_?NN_W2\HNC/T7]R6D[[I>;T:.AKD:N-;@LNQfH^
#-S;0)8<WB=3EF?;5_91NX=:NVAa,#UbXMK8^MO2>NM_FC-B?K\A&-aH2/#V[T5;
I@a)OWd#:G?(QT;M[>.eB:11IZYI-:7_eYD8=gLQ81R,=0>5KB+&;GGAX(X4I?T[
+NC1FU/5gG:V)FYL=Xe0cBI&(aPE#^?(<e=9c-^A(2@=B?U_4R?-)Lb?;0<>cbN[
ZXa3Y@[PNH@_QAFKM557&;RLS;d33?c0MHbFEKO/5c8Yff==D#aP#,TA6>eT?+aR
5(PXRD;YU+5MZA65(db0/_&d[)@Z;,248<;J#?:V.6/\Q\=AXfWK:P_6JYGB>Je7
;D.495,0-E6@A7@&6=0c=8VA^Y1&ZW\_3VZbLGC.8AEIY7G-6<=SKf8Y5C;U_W8;
2^,NJU1Gdd9K&O7);Ha5)\/V=1R76Y[ZA3T5C8fBJ<3@Z=T&N<<385I\SY6>P;?5
+g@9Vea-2=+KTe^=E[EQW4F3G/D3AbH?L??M]VC1UPZPT37&EI7?;L+cTU3BF?Ib
Y56Qec]4?3FCKZfN9RCM4V^)@4#)Q4FV_a08R0C7SML^;I90Qf?T2fMY3.A^3=50
8W]YE&g#cRXM2VU#20f4060@W)HWJc/f2V?bNM@g7B<dLD.726+gR;HcLCXCbGaP
+/R6T.JYf3HbgV_Pbge-NVG=AGSaW[.7?&XeFL=E?ST;>@FU98;6>Za9WL=bL04B
DEZ/-UN)=@&>^(788A0-H,\W(2/;(deE+ZWP-bZ25b(F/K^P2PGec\@^JW18T;G\
cYGcV:)JXD+)Q77F;KT>G7//=43O2OM0C49g[LY(TIa.758(]=NefAc^3GgQ7&S.
VJW8IE=f[3e7M7b.K(&J=R#)c3g-Qb-CO+R^Xg(()_#K^,J#B#\1f4FD-N:#d6#>
LDG]O7\U\@cGDPg^>112R+S)KeX.T,CFg(R6D5/OTcFDF3HWAL6gad<TQZP1OJ^5
XDd56[CabZM_.TVJKTC#9GORZbaQTeB6M>V&a#X]+YY^S0O:S,>(2H/&S>>FY[NA
KE[C4@8TbSC(809J.RAGVUQ1W+0/aI8B9;:7+\&H\bRC0V+Y9WD[?O?W3BaK./TY
J<;4VBYaDZ7TVggMDJ].+<][1#18S_B3+6+PX(7c/BW<aH3>5UT#Y2&[LIe9^4#W
>.-BK(46C]7dO&#aEb[K^5.?3XY6AA__7Q@Y3;;&64ZOWDYO(;\)8S2.1(fE55b6
NV]N#Y7U]++f7BJ+f&,aT?<&<U2Ocd1HCLI_2D;G?17.\+,+G5P)IZ?AH)XLVET2
\-PY)E;M=baW/H)\:>(I2(ELDQUaXaHA;T^T@fZ:QeNf4TUYV=X<L1P(/0WWa[f;
S:S5/\6+[5H/0M1[?f&2(PA=>X89Q/_CKd60#5A:INeJCTJD+-RfSfE,M(UP>_\G
#95dZ:]2b>I+[0LP&D^d7Nc]Kc(;UX@F#T/8HWV@P9SMH)BDTbESJde?7>RQcQS-
HC93>9#\FN3\N.a_;(c[QcJ##9F6MR4\SaaH?\3Qa^;8/b\BMMaFQ&<CVV>3/,3Q
N.U2<)\Tf)U,4_98STe.W/TG]8H=9R1LDC&YA?BD0G,3b=(1aVH.#X-eN?KL[bJR
DJ8>,PRHG-.1fRLE720,=DebTA2D=.>MGX\QH(C7cO&]U_a=0+G0GM]E8;5JDMOA
#GZT^,g,;G5bXa)#dASV^?7O&J_eG^/,]_(P@AL)PZMN4K\Tg:;,R..T02>fHQ]Q
SBcEZ039b6I_.ebZP)CgA.G@bQR,Xa],//<K5?/>##_g21NP,bO:ee04M[9\\UR@
KB@CV0Z^)AUUdRREFVH?Q8]#5dW25&(I8gc=\#6WDSAd<b()Gb=QIV9#LT^a\b42
e\\DZ.JgN:;K9aC,M^E71ZabVGe8A=>]2a^RN2Hg>_CdV8da,^#;,=4]^.WZBYW5
_;.CB0A?ALE+7=9K4[VfPO&#L6Y-&BJd5>)b;/GF-8]He/9=OZT\U?PbVg/RUGaT
Bc#;NB)5a&_0:1YP?XE0FCRZH5_UDd)UJC9,6T/KPCgO+GJdBUY__KVg.N@B5=6W
0Ofd]Qf@Z@+96&K[bgF>EA^DU]1?8)J75/GXUca)PE@ZG_LP)C3F#;PXU[?)^>J6
M\H0)_L-E-GBYY8F6Yb6Y/M.&L/Yg0CLURY?AJQ^J?Z^<X4[.P^YEcN4IYQ?SWf\
d+f90,MFX_#NU0c)75fTU=YOXLb;44[.LMY^#6N^^d^NI5>UVB=QZ,6gXgU1_YAN
QLcXI:Ad(gXYSQMA;e?_gSH16RP:I6FE)KNE6W,U18\IK^d.JMW=+3_WJ]_1e5C@
Q;&8f/U9RE-;:ceVH1EL+RTHTg89<QcR]B/5:+/M.P5XN8/?I>0YO_^S@IS1__S3
e9HDMG,&<g:cHW6Z1T8W>0>1KZ^Sag)+_ST6.#]a8-=D3--a3bZ(U__WA0[=N@#2
+)/E3.G,8UXIZd&4]G&eO#e,/ESegT<AV?>HaS=]c2:HESAT2#O#I->M&=UP7;QA
G5(S/_9.D3+TJ;I+AB3<RfF8>,)/)&/_M2)T?B,];+)]PA@feGWKO[JX282@0e(V
3?#Z)P#=b8B(dbMe2@:R:)Z/A[a<&W_.3?[_P=EJa7_D/YgEb-9.3/ZY;R/KH@JZ
Kf#OP.N+(&0)4^N3<;ZFL][L1a&)2>1?G^R&g/ZVX#^G\daJJ-U[M0H49O)D9WT-
&1eTgg;O419FVQb^XM79_@YK71A)V:@S3;1-5RfV7g_)/A<A_[Y7C6\#=]]@e&d]
9EUQUIX//T2K+4>+?I[KKWF5[b37YSQ>ERcg:E>b)gcFAYVNCbHGS9AP/]=AXJ6(
M=5cbG24/TV\=IYU0e;a.?MH6V8D227?fbRe#,3>f/SJb2R_bN)>0XEc3.5,e^U<
,2U6+56?&S&=<QL,Q,9W\I\e\c#YVK1K)+]g>^P330&,0-A928^U35JJ<97E\>EW
Og=^Nf>AT,_+5XI;&Y=BQ<ZNTDAF\C?^(R44I=Z.\A@a&QJbBT^[2RBUIL-fXUT0
F@P^2B9A+WD7C?2/+F),_B)67.VI)@bW,FXN2_4#B3[0_d4YJCNF>HgM#S-Y7=MP
O/Z0S=?fCW5)Lg/_EO3.EP=]C]W?N[]Fe_#L;,2R>J/I5YSO=_c1/#J#9bH53VL\
)-JZM>9.,_-d3g_3L9T?@Zf7WTXUb(;W42M0NE/fbD)K.6)[H<C/[>DD=FBaa@b:
XXSgNY6aDE3VA+)2X7PW]OZ&0?3GW3OaXSZ3,7b&&>a1SPP_\YF_WER--<SHS:/K
K2B-FK+/f]=V-bC=0V1?2([>(0P>dX1/:c4W3Q,&_3>O;Tb>gWYJU,\c=g+<V0aR
(Af>fAVaKR;SF9L1eW@39&g8Y]RM;IaW4d[Q-eGV+8\XEgVW=VBB\HT-ZcPG>+5+
58O2cc#4-#9aeVDR,QfP(g5S50T#<1@M/F@E]>YZe=2/\].,&UF\])3ER>C#HFBX
@7c:aO=_FE.F:LdcYU;)?-^Zg1)Q;N\C84UTS,U&:5P=HdNDC3#J>-N^@[2:QB5;
ePX3N)VY#:J=TU:Q0E+Rg_N^<W].^^2)AbG:\e5Z_e7g.(06Rb71Y;:dCBJY[.e+
#d5G4+,U0ZXU/eO.dY4a5D3-8.S-fV5Ya&^5XK9c)L-RPT>ca:DdLN_U8<Z810TR
3=26#(E&3Pa?/\4K(6.;b,XU#3S8TcMKaI-@?8X&a4Hd_(3g5+dHN20e.KXZP\Q^
-Ded)eQ=LeBF)WZLJb+c];K32ZNQW#R&:5D&RW80FZU.T?H,g4Q<[?aJgXCQaCUD
XSJSV2&Y@CIO87Sa3D+70L)31?e#-ebRO301A;B+MEJ;+K3-a+2Lb,1D\aV[FM4-
?0ag>HTGc.:9SK.\X_cA)bbce3Le43d9e?RI2FW]J)Z2MH+E:)Q1R2W)A2O>K6Q<
LXI\+)RTLU;.a;STMAZ>EIA\.5cDJBH2?6dGC;BdGWb]<IV35[_/#=8b8T#B;7O.
0?H7H9LNa=0G[g:3EFa4G#ZecC2MLfcKg9DLIURPROQ:)JH2=N:d/^US:;SP66O1
Z:#C(_@M4C7cU_(\e-ga-@IG#X._baN[@GgN/^96NWAH4I3Pb1B2>NX5-?OL7^.4
=\=(LSK0QOP.D#3We=V(&,TW]J+(KN>-DQ@.XNb[@(X&C4()f_(Ug)eAc+LR4e:0
J]@9F?9dQE>6MDW/bFa]I.1^_bZ;0b=U0@3ZG.?YVL3>B+U5TL&0bFYgWfe406JG
]5/a#[a3JV3PH(=O3F;E1H6\OS7_3a6ZYQUR):VK@L?/Wb@S-F<LA.X:[]g@[c80
2W:DZd\DCXC7XR&fGLP\+,#G/=WWc_D:M-&:;HA0UR:>gZf&>1T8fT\6^J,<d0:N
0AZ6^IS[A77U-\bW\D=?O;>7AGX@SJB#/Mg_E+[Oa@6Q(?KVC(;,AI7g:44[E(AN
FYOQZ:,?dVQZ2(UZBHNPK&,]9FNeYLO0G9NTb>:[BER=g9HJ6a4#?^0#0;Gg:/<)
R)B:9&K7a:45V^?54dCe;H;D)H#SXa8S(Pgae<<L?#BRYa;V,_IA/BPPLa\U]69+
>_b]98gZ2:-Da,E@#Nfd\AOMGCUPZ4SB2/1^,9[BG3__,EK:>AL=+g)DHDHIFZ&a
_>WU\:G6-AU#&<GbGa<D]b_KLOa?PEf[HSe7dPg=WI#GWUO@efPR-.^)Y;Qb@b&2
O6R@(^1B94UH8492O::(De1YedS5+b2WF9RGc@;c:6]MTMaQ;(/+[;Q.WN3<H3?7
J&&U?DTQ1=BOJ+2-&/]MbDgeJQ@-I:c[V&MWR6+WO?HMVOIT,7+^;J6F>a\b(EVJ
>\S&LJ4QLU(^,;,X45RGESa<?\TKV:HA\f+@?,Q(U4<0+:<[./VZV4eJ\1>47ZD_
L?QRbXAY[6OV;[QGCf#X.0N[7c;6>e5^WN6g7HQQ5Y3E(56I@2KX\(_]Qd_d)b2.
3,BPUNf3XbFE2I^RI:4&XI,>LeC8g4</B1dg:g,baWMP/-#L7_D<IX#)__\2d?b<
3d+EPR5bWBc2O1g,KNB-53OQP6>\34/aBB5^c?+YPd68?YZ#[>+BMQ[>PZ2e0ZKB
#_G[bO;L,dE1G#Ld8]H5&<Jde,adG07[T^KB8fPK3LM1+TR/\8NRH&c;dZ,(4.(J
L-[d5baKH>+^P@=F+2cC-^cJ+.6ZB_aA+Q@a^+g2>?7BDOP/b>1]F&7,AI]LX/]-
3ON3+KMC.7Y)HMPUG]8MI\&C]dZa5:5QGF1.<8P>438&J.DN1XRX/W(=WW-F_.PA
,eE<CQ0BXYB4HMa.40BD;<EM=GV7fS?fY,YGg>BF;@>e^-,[.]R;2&[<A+M]XB.@
+?d9/@c&O4[Ea@;SDQLW9KIZXNE3\T]=;4DXX[aN3QC:X29HXSQdO(,-#X]K#_1>
NQ>2ZbU)0-[[HWYgR&>TH-R+^#K];#(QA3/XVDW&0Z./)>K6_EZN3H9Sa+#G=H;^
&Q]=K_8:E;7/C-[U4<\\6HDNQR2VIR2:H.I1Q3bd9+#DRM4QX8;;OI5BK<e\^D@=
&AHJQ9^[=X;9PGA;S=Oa0PR=WJ3C58feBD-O,7XGAaf<@ebTO3a(9g=deOIDcd0>
#]b9WNR[P^eK0J0/F+UJS1>c1JQf0P2X3cf/X:Zg)-Z_XQ?<5+QA,W[27K<#@=Y6
Qc&1CNd+cUB@4M)[41:CV_F)#fKgc<fc&BM9fCL5U5)?9-GTWYLCF:KSE4^-0KC&
6O6GF^GO.G.SBb=FVI-f(e;^<G\A/R7cH-ZJ5c(JENCANHFVfA>Q/H3g]03E>ZP_
06.g<XF:?@6VFHIR741RcB[3EUd\Z#]R?c\gaI[g5Xb?(P];WfAU&NFL^a38C;0Y
=SRSFKIfO2K&DMCZDf2QRU<Z4ZJAO]&E=(Y35WO#3b^^,-?Y(9>X1XQAY-SQ6\TA
B(B,daVITLfH-Bc.c4A@:>fA548G,P_O=R;@(OZ[0RYc=3R4Ld#K&ST\0Tbg0?GQ
9X38J706e>0e1aKSd1^+&JE-GgGGdS1:&2AMb<]I;J(_KEQEbbD2IGAQ]cd1GSde
GWEdLNO7WJB/ES^LY3_LSOTPR?F,D=HbIU,NLg6Q&1,VT_U.d^-9>B)d^#V(2/C1
]<H^T,X4@S1#9&SR1G2Q<X#A@Md(P.EPTUU9_B#WR@6C>=0_.6=a3>CW#_D5AC.^
aTf?E(=N(FLOU.?N#&MN.YEC5]dQ;ZFb]eP&4_&;T6V0BS1)bD>U.b<^4f>M\[1K
[cL&V<(;#FPD]J\>3?44E0VLR&b<@A9\7O+R+HGbV7.)(6VQQ\NNC)P@N1g.#d3c
g:J[VUZ5PgCZ#,25#&E]>[TA\&<ZA;&?>^Q/EUL7R]0aXA@.1A5>)UYZORB2-:(K
gP>).EPWadacK9\10U4_QHgPCd/._O,?df7KYad28;a.>dPV[HU?9a0;.cU\)@U0
[d,/+N(31IA)=OHD:\&Ca=44GG)2HG?&(#YFLabF6C#E==],FCd5L#&//+Z<MBKT
N?A6=N9X21DTR&QZW0:IJNBE=9;-:5+85cWf8IF?A,F5J_SNPW9G(3>CM;U:D@9;
99DbXA?F2f8-Sd2TT#g<.Y#MTU,=Y([V9O#d\[N;I298=\I._d)e\U7+,.c++&6O
/?@-_0>WZ9Fg5RSU)&XI]C,/VB=H<O+Z4@Z\NDg4#M8X)\Y-g6_4VD&R2C(P_08C
,)^NdHCL@\^#cE>J^cE51=.^PJ#GY<c387^&AOIG,c^[,+aScIQ^^07BRdY?+51+
eb6Q/C1,_-SgA.S#UN)H;Q5bSQ@9_2(7\.E27C[RO;DT^?S^^1R.D/IHQIM.&a(O
PAcfg@2U_?g]?&d6]11aZE[4/1?403d,Gfd#/B.2^)KYPEX1Mf7X_SI868VU<1^X
N/bU?(&LCdQELZc./GVGNQ(V4Hf[2E;-gK(gM\0^S]3T&d[JdPf7V?E0&^]GRWTJ
\4J)XQ@RS?He2K@);2aV\--YX(854ED7-4STefe_#75UOea;L)XT4.&#C;c:B+_6
gFM^2)G:a4/bMCE#J@M]9[B,Ka-gZS\NK#_IK3#[GJ^I8U(VL2_]D/Sc,A0C^E<O
0(efHV9[VU:[OORbF;YR:QC?R4fYN[9/MN-c=G(<_3P4>N7S0>-YJ8d_MX14Q5Q8
\+#@7)K@.bKO.XOIDQ5MH:O+YYZF(._?>PDNgfQXL?@MgcPbNS5,(>O/2NI3gP^(
Q-LC/\]U6H1Z^M0.>7^3BT3>,MagJ,U=+/U4BL.6ZW,]dF=/0YH.@(bgcH,WAPfM
L5b)XLZ3(\@KTa,5GE)CDdG.b&d/d0(.?dcd-N)//e3\D?F3?(3O>5Xd37\1:0>B
5JbH4c^ZgDY#I_]C>)?4+aUgEMF]CBXXgH[7eR&VZT<db=T#8eEeF#)3+JT-&E.V
;Z]E<G,>MO,SBHAQKb28U2.&R^FZ7VBd-g.&7NKAe4S<(DCe1NCVfN<dD@^?QPQB
BD)ZP0PS&2<cSMXQd&Sd=VM0Z]aMA/c4I[W;#Jf<<4Y,WPL]OeT3dYU1/#L)K4-Y
L]_0EfS^[Z:SBEg@IY(;(UW)+,^(b=QQJS7>2e_^B&KN3c>HS9Zg5@V)289W<U-A
BZeG0R6_[gJ+VHFeDf_O\@9^J4]Ag#8?d+\4-N@TXa5Y/I&5eZA<KYZKL-#(VV)=
1(2C:LdGD_LDcH[AQ_g(K0:;,:SIY9L0e4@9#Rg[(5L<D&FdN-)RK4,dOM\LON64
\faO<V3XN5#aSaBG-Bd+gAcJGHN-<)eKIQ.?@51CU@cY4R#ZK55@;Vb-X:1Oaa#H
8<fG47.:M6(I[2aEDHR7Pc<U<)TX,NGP_\U4cM[:RC]gFRAWH/-HN2@A>W:g^[gQ
HW.2gM9;AD\f78+0+/FI\>>0ZU]P^?9).PN.FD0G[g5V_O.[eY?g?\3LI[5N0f^Z
D9E>F:Qc1735YN<P&_Lf(0#@I9,;Od=]=YI@;7T)J[-U\LN6eb>#32&O(.eL+:EM
Z^Rd3#.W8;d9P\BbL@4K(5M@DAE7e+Y;KYKOgW[IFO;S8cN]H<Z=23(ag/DIA1Gg
4T4&f8_1O#G[X?]<Ja2Q?aC(_6L4B,[PS.+<dNK[T:]A)S69/1=)4W62Q,3B+g3d
<7:H&:\U>MXR=&C+WfL1=SS[eV@<c:fb@/P@+80)63UWcFXR^IedFRD]X2gT,T,/
9eN+:10THMeeSbAE5B7g))2e^K=\daL<U4E3/,R^2UI#W:WO32c&g6O&E9L&F6K_
.C<60W\Jg9Y;+M#Ge.T=N=VX&4Kc_7^78gd.S8FPIZN1NC^d]=eg1+FRD+IZFGA^
1(Eb6:FfGH(_)?1:-TVML-3KUL8A2#;26\T<18T9I)ZZ<ZT1O(Y)+2d=&;^RVD-[
9&ETWL5-PE^KTe:?e+J?CAd44O317]5?[/LP_7HS324/g_(W2\>fA@N@)#b6a+(V
5<8_)d^3-/5C9.\b>WQ/5^;<>+5c<Z,6Zf<^Fc3=CeMZE595N75^:8IU@.G@gLR#
-&KFDcF?8d\U\JNOK?^6:Rd;K;>eYfa,+ME[SO(;a_EPA;caEIc#MW.CV;GK+F^[
]FAf+XLdJ:fOW8[\<7)YNU6LT+E\)&O3A2d[#VN8)fNDcF)O?<F^UefSH_P&YJU/
KAGRFWfc,PLFUPA-,eeJ7HcX95(Zc&g3:(O>faSG9Z5;Z^@-e^:I.A8)a^B^/#Y6
>ODeTb\L<_a=d;VL<5QeJL?LG6?;DD;2bbf2f@LfLPEN(V1I@-bK.GTL9(C3-f/)
:gOKG[V;]W[Jd>@gB=4F]243P1;0-F4#OKY#0d]Fe<2Ee\(@GJ:KYgI\/D>dZGbQ
SYU[Q(<-CN(NO>dG)63Z3O(#[WXJX(;^Sd9W7a^6Y_F0IO<3BRgC;JJ)?F^CKEgN
IFE]/2fJP^Z)MJR)1SW/FS>QD)=7f7Le0)\_QZNVUCVA8-@K^JCde:LBA4;<Eb(N
g-dZfIEOWadSF)3FdPDO>.VIMI_VZU-S(@6]1A.VF6DE;?4\76SAWR)DS=Q>#fDe
-Bf=gHDB^.H=_d)<P.I-gC?O7AGL4?;Fg7+LDA_Xf/--\-4.\J<V;PX@HBPY2??[
(X#7YRO2W=D03641Jg+W@:-,MW,5>W;cf5V@G(1b0bI.AEM&#;(4e]ZKSVNOUg:f
?[c^K.cCMAeQ&SbcI383G-#Y01K8)M-U_GKG-/MZYKX6]?T6f.G=X#(fP8IN,ESS
E??:&^g5^Z2:#7Sa-M.&]=O)HGK=c6_/Fa6._9\74>XBD/+GaLSFYUg&N0WQ9+I(
V[,I9&D7953f2R:-^f9./a4Kb3WQcPa:53SLZ_.Q2]Y1I?:UDK[?a7J@)XYXBV[]
Jd+,UN[ZERHbF^#70T16]Q]V7?M_9^I;JFC>MU;a+6YUH>Z.b0(ZI#>G9BUFeA-.
S+6WD9Q5W<DfF566gQW-ZYgF7-KB.?7e+Z@1QV4A9J)0MYY,[679eWD_XYdJNO-V
IBM>CV@1Me&BV_YgK]#<G3_P4cOZ?.W.<ML.EWF(_4SI#4,KJg_K8P4XR/]]<<),
H1].HQJcJgGeUg<7K8Q@N^S5S&ddb5S5]>VW87<EYf+_2-C4/3.-Q[W?Nd]a&):@
8WUbD5YVPb2/F3-]<0<2WU/Z.Z+YbcU41),?1GF3NV&1B,Fg04dd-ZTL0D[MAH6L
]#22BLbEb\H2^Vg,Xc4U0;?:?b7ND,]@H<4?Y==B2eUB8&M2;LG^F7/I^9C>b-#A
S\@N@9QB0RG[]Z3T\.dgK0WMP1E6#76.RF;^7R9Z4AU/>b)&8;_?cN5Z8V#TLA&[
>VMf9,-T=T2RIVDDO-JI[VZ06XBCOIH#da1FdMV0-;-5Nf)I0XON=.+AaO\gfaBB
aPdL5Ag#.2gFF&>=:E?4;S)BW)8L8[4<J+WW]^;9B2e<KG6g9;eI_5W8(8_ICB)]
gcGa6.1W^)3[/?@-3Va+2+^(<+-a4WPZ=+/(A6#0Ac(;\W>KH\KETPQ,6R,.?BNe
<((,gW).S+#9e(W6E12O<7]EN@BG7MUZ7;4&YIPN\DX;RJS=+R-0FaCJ2MPTG,(:
?C\0QJDJ\J1H0LRC@SJb2/\IX@-VOEFV)<=.V26-a^:W==@?7M2EPPT]C?GI;^;g
cfW2JR0;N5@][PAQ(]Vc[2\#0#F8LW6@PC>7::V-0WCS369B]?&O#,_IMLI)/<3V
U;d[9F4Q=T(;[++)&<OgN-#J/A\c,F8+3O/XC0:XD=:A;T\-c75,(#BJ(#YC1J6A
8?]-.gFe1+H:_)+/2&SI:Xe#2d(8;/YJ)3;]6:)L#;M4B=XJX5W61eQ,\0aGdg@R
aN:?URT0>MZSb<:b9<CbKWdOMOOgJ49YYW-Q]0+8NQ5F]UG>@BTNd.2bW.QU\1Hb
&QaVDK<&3JOK0?a20Z1@&+>(&gR[_aT/7+c(C&1&ba.3NfHb=Q4\B6A3VQP@d=&G
cOIW?V7)O5C+=aO90(g2-\:95J1FgScgXgC4+&dK,G1@=&DL@7#O2>f\B2:((Z^M
aMf+CcNIZ@GbE:[K2\OR3E3@M,e=]1=H:eC82_95X&/bWLL+4/g0V,Q3\:I.aQ?U
/XOQP4P2+S)H.E-HC&R9a]09-CPJ\O4Mg;:K7H#d&867Y>D,bf;7SU;cNA2ebJ+2
MAZ4TX4ZOGWE2Vb(MZFb48SZSNfI\D32DV^T=+IL^RAA5gIX,<2==Pb[?C#WcXf=
d#c/IeLWR##1+Yg4=dVZTU^;KSEW\KNLK(</V4C=U(eC[eT+]?4af(_R&H^.3a8\
\@NY?J)ST\LX.<\#V^.JEEK-1B@7HFKF<a<Wc-H81\F.fRLWYT^/PQAGYfI-(@:G
;,_TKMIeQ/#Gc0UZ.eR/+RJQ-aZ-eZg.KLeVC]9SU@0J\N+SA4IeTYRSBT_-dR9#
#5<G<TQ&:L5/G/YF)MbNVRKH-C,OVaZIdALGKS>-NIW;=GOREQ2DP5:>:\aIg/;Y
JP7O8AK301\Dg=+>#RLSY[PbO@Q1++bA9>[D[U:4Q>?M0SgK<EKI]DeOgR<;<?fC
VaV^3,<[QJ#\eYVOJZ]V<4(7Z3252fg8VD+Z<WX^=EAeJ#)A4E8(f6SF3F@4:Gb2
X.SW\\1#/8@3+f729(f#YD2EOZGO1&ANC3XE#K@-OK@2?E4_]G&]<6JA3OP/[BdX
3QP]B=FVaeWKaZc1?JdOOc05bTR,?>P,;YbCeb-4GRXB2).8>;,U<#[2?QM;Ra)F
.gLgGARK\V/5[S9-Y8=O>WRgP+,&/5FgB(dQJB,2dU78?:F9OCMYF#<CUH@JQT4V
_F?)U:,/48;.F(8T4O>aV]L&,e@Q^)#)^W>[bC0T)b)acUe<+BI(#+J__Xa?4^,<
./SUN1U;DMGFIXC\JRVEFKOMa)A?Ye.-7e^?BG++N#956cZ@)ZNM,,E76]G^-\Je
PW4)/Q#84(27_N;=Td_b_B&X=4R:KGHaU(/>f(b_=.AQ+aJ=_R^@(=K3U43A&/Y7
KZ+bCb,VIP1dDeKBQZA0>+YJCU^-=cD1F+9TbH\-T7R+6(gdC455IXSEI?9F/6[5
ga7E3VNbgWbLNaM7:+aHKd+<=>AN58E<Hc,Fd3f^UK5X8d.]IA=05g?fXF5OL^=4
R=J@F=d@cK2.VcY478;)<5@@7>BV&,@C6eYJL;^3MLcO;3IE^Z0T(/=38FP>K;O]
2<PMS=D([6<a_;FPTf4QR\0g]]@Nb1HULZ3Z4UOMJLe9KPT4AC0H1#D&X5g:F_P<
YQ]4QG8AC(O3c_48#S;F+)RR_=OVMD.=27LTTT?W\&J)W70a/(BG:\WVa96H#56H
+dB7Uf[1TM.X=90L@Td9G-1[,UM56N,J==0b2>aaSRV5IZ,Je_\GG<f0d;e/=]/c
J5/C2#8&>QVG:CNHZK,0A;e=C:Ue,8M</NU4_FR6^Q.c:?<(g4Q+X4,1UU)?M?#=
B<<BF+^D0\Z63M^A,CSER<\.4I\#16XNK0/Z@3FS7CA77Zb)T[>JHV1+)UC9H?HR
,=C&9M4cB_TQ8cZ@7)K+d:5CXO.DG\d7Q#=a6fGG78:=d;Z>CGP+d<W5)b95ed+<
Z6^P=96_ML9c(dVIg[TPe51Z0KJ^LDOH_Qf8VOfXGZ?M0>U4H#+79f^EC59;JQG_
8))6]T8YY3-K,K/A3U3(8ZPQDb<>&MH[L1.bQG]4eOG(?6DUD+bXGGP78F^6.^@d
Q_fZLaG;HB^0PK@2d7N8Of^g=8M+KT?+9+(cESK@7S]3<M4P?BY:I?(S(-?#VIcJ
OT7[SULP&;2OF@\PGT7=#W5&>.fVK2^;[8^NG1X/d,g/b)=^IECNCcd,[T[&JYWF
1b,>I>Z1C&.R:B94(Xa]Bd-,DLL0@fSR(D[CeZL#ZAXe0d?C\]N77KVQAgMNcbCZ
-.aD19M+bQP2:5IeM_>];I/(2K51Z?,IPVOc@J<eb?\Q>fW5Eg]MHgZ7.EEOgA^A
0MgBPgQ-?_BDIe5KTf=dPHf9Y?,7FWLCc-/YLRb4(<gJ(daS<:0a9J,AaNcSTO#^
IR(5?JWggY@E:Y)Q+SET#?1^GABN8ea(WRG]Wcb\T09BFaT2NO+M>bG<3,&K2)Md
Da,9JO]FP/P@e,.QLT9AF9[EU#]T(TT?]0ZRJ.,Jb[5L=F\<Fe=Ueb>F\(SNda3X
5A\C4WERA.[335<KOBO?^<6_[VL]TJMOZAa]B\c[8BOTFeXU-K[0#.]TRVIEW9IL
^\XK<O@U,GE];HYb=0UV^7c85@HB@5<[1d6A2C/FC9)NXUC]aFCVC540S><V)2cC
bDN)dc\f@\4TAX5_c<;,)B<@L(J-&)Z;3C/GBGW?Y^TC;b+e#&8Jb8T0L,K,]];<
=XZ[c\L4G>/@#Eb4+a)E[PE_PT1.KD&.P#Fd&1#aVeTfH);NELWN[[VHT2Kbf:5G
F0&4/gBB?R7b\QGLCOV[SE^OFF9c\dcd=^.&9X)0^gYL.K?T.eC0=@-VA]4_R]FW
ac0+H./#V(E<X[f0YVLNSg)F;4.C@V6d\>baI4:a=M2#OW12dEM>];U7#9E<.]f(
OH)cLbZ\-V+\^3d&3XVdNHR+IMD8)@gLN_D[A2G2b?^1@A:97;+^,@LXf)YI^S@E
c.,Q5/>IU+/J,c^2U9cBVHW]&4aU[^IY<fTfVGF3O+&+dYQED+764f.YA46MIV]?
\>)9R2W/(]9U:H)cS<BABXR?.=:QJ_dN)K#91Q]8Xb@V(KTNT#:@=>],\bce>G=@
KSH-_M1L#/VfT6eGC0gI+cW#UDcO\1ac]^d7W66<2g-Be02988cVY+cb+aQW/W&N
KIH7.V)?)2].TK8f7M6];WbGXa@0/5WD>Z>^H02\E=5(c3)(H#6_Vf9:PfT.e[2^
>UgK+O-c(1Xf<[0]N@O32&N-_eB+aPff;CDP3I:N]QD[P_OR:OREHg?W5IcK1f^M
B)H8[WGC]B^I8+JWfP/3ZZbKcW@^)R[Z8bg=8:(Y_b0K;b)C#GNEQF/VZ8JT:IB,
[FG3>D<#-FN_Y6:YOP6<=ceTQe2]^0#85ef9^_^V&#cga5CaTW2R_K0e@cG\eG0.
cS2I\186/+&E#MDHOP^G;>M2AM#PbG[SN@BJdEW-3LK6JP1C?\_XU^J43U-^9J\&
JVdcgMZY0XG#&TV]cg25919=NU9YMY)TWFDOG+\<?/S]MNa4FZ_89^S@T(fV<;LT
X)P5?5#]IC/Q(cC6K.d\3:,DgeZaV8-X8VA,@8KcMEV^X6E\M13R+gcODU4DYg6(
#>5^Tg4J[,:W=Xe/#7?V,54(_F24?U0fSQc=X=RI.P5bag>D0eT=>c-/VYLcQ.H6
]G:L.W>]<.0L9+J(<,[IUY[dS7QO0U?&SfMF_NMa@W;M(1>868:J,+3C2dIMO<\8
W[W=f_cQcQWXPg61Z0B:R?SWc>><;3JVX39OEBZ^JVbMPD+#5Z4ZZ3^d7cC,H/+b
:3M#RU0-T[5:0Qf8N/0aH0b9[3FJPA>0Z<G>H<B1(=#-@?SW>O=[E_NTYgLcVG,4
U-+Z?I;S)@OGYRG1+c]>3W8a;W\9deCC16XDM3#B),NAaeUD]a)QL-LR(G70M-_V
GZ@=C>fR^9T3\8Af<FAQgg3CK)LG+df70HbQZ48If/,#cQX7Se\=SMa9A7081:LJ
,G2B+)TZ3G22fO_?@&8-6PD#EA&f;[Vc+K)GP<YX;\+ZgGAXLe#\CEQd]dK[[>]E
QE)1bOG&UM-#RR+XN8&0&\BZ(12Q5FTbK5f/K5;AWZF;gb7@VU45J.ag)D<Ha\AZ
)c0R]OOgH9A=)8Fa(]KE/J_X.K,N70g^XQLdXHP>ggCB[:A>BdIP2M_(5K]J=Z-d
V+VDAYLLF)>R^/M1^<CTKU]@YO[S\]7QP[&]0WLOWM:.W>eg9PE9Z^[[XL60+Y:&
].@GeGVTCF?J=-H3QF#QO+Zcd.CD3Z2aE);#9>\\@WBA)Q(6F>2.76^g-^[/c]B3
N?8PgUe->215<\=b+7a9R4?E5R:8?=SM.B&d+eLDRf;OIU)[[BW3?=VYL+1MfEB_
Q4f[OV6V8PcTI5EH(Q/Y(]^1\F80T6RFGX]VZUg4YN2=g<_a6S7dEa=#:O4.K)OC
NO.JP]P_3+fAENN(gDa)N^-f=[TMP420Hc4)IPJd(.OI_8TCV:1(515@FK\Ac4D&
[UCCJ^M.UfW=_:L;;_.<.X]Z8>OMS-UM6CJM\T^?[Q94):5/^Y3,(-C0d+JVdZR]
;Qb.#LXJa=:F81(N8L04f<VZ2?U<R@Ha(Z/U@N8P\6;3QYK@D);QF2[P?:VNTHW3
^@@S,_J(S)76<?;IHbO0N4a75d7gAF#QA:D&)N<\(_M7EFP\HK97<ND#Te.MRI(8
eIB+e4g_,gL#JbV=SYY/3[.,SH\FFNeDbb]6]<L]?X#2DBc8Z02R1S6WPSN:a14J
RcB;5O7#?9aN:HbWU;5UXBAS;Qd?VKa9.B_[KXYGe@@fV:4d_S^8I;GQ7+WQ<OMQ
/#H43Q]61FE?VC/&Ff,?]d-GO>;Qa=4IJaI@+^Wd[(4a?KJP&aTceObf7XZWAV32
,CAW1GH_64O#K<>JAM^UO/CcMX9;B>+7aOLBEQ,6?a2KeY3RJ3aP\aSM\=^^e7,=
cEF?.g55J.b&F7G:/AF+^)0M?0>^KBX&7J+DKE[P,B06;[8BY&Eg1g;PD:;-=GOA
b^g/Y@3I4;NOYOa\;[,f)R8R.=)+7Wa\,7E1Q_E#GS>3QVC,g=dX+We_(@E<VA@G
]XW(\8K8GCCE]LOfNb<2g<+6_>b@TD0VK1A76/Dg&G6T-b)Efe5?,aB2RS3[>,BT
#_8F&PG8ME,FJD&L#Xg1N;9gX2+F84=.V-)-#gN5IALP,c#XQ<fA)W=EE]Jf;1<S
]#\6_+.[^Y=7a(X<G=JR5SK:34c=G]NQEJ:#VAXUY/aLD1W\7eP\-.RTe.A3Z+8Y
</c30T]eT,+WSNcI(\4X.9@&75EeE#A/MI;&C@RCPM1)LCLK;dO\9\f.VOCegS<S
;,1JJbV>D84FNBFT_VY8T:Fc+U8;CDD6T@S_S?@=\I1JJN<;G,9M2(fTZ-:a>QV3
fNU+>>\O=<(80P@\W-e01d;b-)T(ZEBB=.7&9O&6gOOY:D5V&/58I:L2F92H1fO6
_E&)D51U-YQfJ<F[c+0H7Y4bW#;#05\C/)VA.MWdHJKA<ac-)YH68#],.L7(1;X-
X[9VKZRM\-)8.:]GFYLRHFD8RRdK&SDCfGYC\PQ]HR/BFWKg+<M4+^2d9aJFV=K4
=IM:K[0PN4JL3W#VNeGgWM0:gdJF==JF(U]B,8e]9Y7M@RELKIQ)g5DHPDLNF<@B
P9D]UQ=<8d.[f?IY4WET3gZ<I^G:E6\LGF)c:D3D.Y1)7BacF^-Q3CF^LYH]U=<@
0)UH+aB6&/TUDd3+BJ.71I^G[Tc0L[)0#E]1^I/I(#ec(N&2b&18?dK\X5.<<f^.
TG/\B(@SAF0WBc]I<N#.(\I-#]@]RXfH&TMV_&df[&RLa;1c&;ILO]JZYS:8eXOf
9,QM6=adJ=aaVOF.e8,BeMNL<FP0&0#26b7^Ie2T9()R_d?/[H=W62_G6.7UB9?4
/DfL\YP79G=&AOT:W?)XfRUf;C5Ve&P_P-7:3^gM1;MeA\OU0<UEDZbb\J=X?Pgb
R(Mc0P]0Hf4KM,FQX72J&7g)BVEAAI.Ug-0gX2W9BK5ZVWQf?G>P&NQX&JNNLf):
Zb)fI>LdO?@_J\:C;A#ddbc,Z=d<2gR7fK[JLg]TbcR5+e.;>7W-(\&=LgJSed\V
IVC3JOYKb3a<:db.5(IPLgfY(X@REV^;SGFa4W#NRLSJ<#/b39[&@dPI<RGPV/c;
62F-MX0T5=H57BG27WETRf:eeOe;@)CgX;W<4_QaFBWaD//Jg>MI)OQCP^5B(dU]
DfgMTaHQV0W(Fc#f8OeJ<7YHGJcI:ce)02IcOMfE:[f]bW7D7UbNAM\#LH<KFb,@
LZ[Q#-McfTDU,T3g)7QHdQ;X3_e[Y<<43fV)[1dJ(+?G_[WF1C,fP.:U3S2Cc1Zc
K0#UgJDZR>CeA#KPN^^2)OC,8KV8#>Wd.)(8bDaW+cX&V;]ML;+3Z?cC<M]+79Xg
f[/.&^:@\-Q\d2C\K+S9L(A.1OJ1+<DN:=O;.RIUSUQPL@6EPaGHXaB[M7F=..5G
RWZ7F+AaaM2+a6#=3,VAJP)^VGU>+W&NE=\:Q+I\MNaDV^IC90Kd+(<0KASVI\^Y
4^Z;?^cLBHd+;.Ab1AQXg+SWQI54()@\E85>^:bTcNcAW+URI:Ab2^,S+.+]K0G_
YDc[/@Fc-Y]:ED9XEC3GT(F5IdMU:=b=c/XCYI(SM,5RbbH,DS.\&4GgC[-G07W9
FAO.61=Pd#S(JIGG.E[BPY7Nf[<.=&ZM_YU5)Z.V\@cOT190S8[KW-EN+,T?.H3C
19/2_YV:S3QcNNJJ1SUf1Xf4@9-3WMO.M-Vb]C=:.]H#_RP#+K\(d_Y0,gH55>J_
P5S=IXfIf#=gcMQTWW_^&fIA^O>2:bS:DNaaF[f,?eORZM>3N-VL71e0(VC4:a^(
Z(GC5->D1^DJ^[JbEQ,;Sa4[XP79]R:Va1]g6>D+?7e=7Tb8AGNC1ZFOPQ,Q5@;,
RK/0;=O(JcXWZ;?A>(g9W..1X51>L1]52eJC-R,),(Df?PH)Yf9_C;EaaN=<2?@H
6AeG6gO8K\b?cVFX17LKQg[e/NK<)HcP,]eSC8LeL#5\.FVG,[gD9AT;dEWKGZI)
cOK--#+#GUc/L:U61g1/GOf.1B1UU13.A)PHg++6TgEJ=9fPEEbHU;+UBM&>9#@-
9)_=cN7(I5M4V]fOad4:S0A?.Ra74VTQd\eAe]gM206IC0]+BX).GRgN\^ANd0#;
+dbBD0WTWSHL0KE@HeJ?d:\A.g9PF]OL/c5CSVV&]KMEeM6@KU\X5IF7-0Xa=O@=
.9Ia2074-U9KN4=XUJ#^7GBVW2(e6#M,F>a2bT\9@W>/^>BULYRGH(,W>P02C4H-
A6[DMdT;N&72U,BTaK.UK/@OW/K,KRTWB;BU3=9QfAc(20UW3OQ&21@;-LKKEPg]
fXD1=e+UgKZ/LP\2aP#)F^LSaC3-0([a=GLY=WD;@[3DP.dT0)Y=Y6^)]AT>BWbS
>NA([R&6_<<JX+Q]UaQ).O=aI\f)774U2FA/GXA#@2J;W+YX=JJ58a(92TP8:+;4
JZJNJ\.O.Q:Af6gU3cJeb;>dWg]]DC-QabY5MGBUU+ALJPX:B2=Qe&AWVE]3#(C<
FNL#\LD?O<;UdD<J/>T2KHEO><Q\>A(b:c-)>?K\d]/W8@Z-RRS2UY^a@,H\^3[@
;:HWAHA/=HL2.I@XcWBfN/V6-L^3N=WVMTT9W-eS)NEf@HO.-G0\U.MJ_3E>TWSR
S<@;7SfAC<+T1Fc&c#Q3?05HZKQA0)JZ]H/bF6W0J^6>^C<Y.<cC>+O^HFgMgDO8
(?a?XPC2-??W3Ff@/gW@c^YR&QO=8S-^^0O\9#RPZ<O^a?I_@c:S4K(bPG(TZM#5
J(ZbD+;C8gC5ZOVQIW02EN1UM/(TR558dXBIG:_eD=T)/.-_S_K/AQ43V:S<XgBR
eD\JU7:+N36<S\\+b_dfNX6Y2/R=^6A;G4ZGaQY)_5Y_H=89DWB3a75>E[a8D3dD
:>JRfS)M[F4O>fT;LQQ25Cc.GBL->?@)@CM&AW4Tb-eD9U2)-#KD=A(0_7C,OcE3
YARS9?<F:+@+HO>&BXc<5;PN8\XgI-2@K.gDTeCTH(,7(RE9G&Y+(0E7LB<fLV/X
K.dO4a\9^^=KT[D6O1YYT3(?cNO)=&;A1@-DW0C<JGHTKO^LZQ)W,LR0)?0[7<J\
Q?9b36AVgC6?=a:b-86^?BJ=Kfd<&ebf]DOH^e7IW72R.0e9_8-#7@O,F_I>4NAI
_aA#\P/-OMM,0H?Y:W8QCbB=@eTG8XRW3./Og<=U,=O/9J\Kd]L7A,X1;Y0_]7f-
]EIH.U<4N-<c@cYBT.EFLY4[0GM1g?WDBODfJSESWVF:\;VGHFQ-SNVOg+&LJ240
eRI@B:&3HbNJJUHL,\.RaRP@@RI26fF]NN+#)E[1a<>JF?&;Cac9;+7]\K8PSdL\
P<I#-JP=9EVPJ4+>XRSMKN=CRXO9\)]d<:bSdU@.+A8D8>RUQ(=,H(_=a>;eQHg5
8;Y,:@430,;DGg^FB_-/HR08Z@)d4@2HdQYD>.6OHLD=55WfKB3]F\b8QW]RNEAL
W._5EaX2O9_]XH45(T8=#9@L8.YK=2OA>2?c^X=7TY=\\U\F2X>CNdVO362X;#G/
05]ES2[3\aY7>cA,1/TB+=-<3\C7D=-d1Yb7aH,E+=/YJ?FG2^d4f>f0P)84]X1b
abAKg/X+C;#F,82X28YabV5ITWLbL:g&8gNcQ1@MV[/72/[f-V.<-CY/C\7[@\>T
K;U;+=)+FDPFC.=_(;V(9?;Y/=,2K4T)JQ0QNf<#;@R6PA.75H4(QYfJc)g+1OO0
\eeTFT2@Ma2SY:P<^G3F[)I>O1eS\L-.4EETVD&[\6.J8F:,8a9T2e,^M>Y7ZR?b
G-Ig:CV&6=_B>Q7H5PXO>O6f,8ZDSc/_B>DgDR[B(BO?&&7c>fFVY;c[9\ORO+##
&V/JWNF=fW>6ZIUZP9+0_HEYQ&GP,ae45,>[)YR8G65<(DfQQ5UE)c@-6.W-H]RG
Kg+d]^C48#UZOW@5^(]GKWGK[J3<2:R8V.L_5B+J;Zfdg1NUc@:[7,/W+3U:3:U]
HDSW):#D7)fP)eMdNA6S+=.KTPJf520B;?NY#PeHf?HJR4J?_,PYM=-V5CaEdK3A
F2?7IQ:f-XY<7Z^S3P2OM8&O_Df_6TfT#JAac_K&?YGaV+ABc8X3W&:E(+?SUHC@
@C]C-,I:bTQX@FA[#b^]6^^/KK=.V))SYOc2<H>ZMKALWTIABM:.UgR\A9^Pe(DY
(USA/#,c7L+f#gdU4_Y4TJL>M;<?W2:efO?IgJ3Q01Xa^FOD?c5<L=Z7Xc2[8.UU
7AY3XV@g4/bLOc8_Z-3d(R(<1[R.]SeWC#KC8^>O]).4FAMB@DeL;^Ng98>SZ[X(
=bN6#I.F=AM4,<M+25Y\M&_Y-?9)MXD2:6)-Y>Nf860#>H4-AKK9M&;.:JZYa/L;
.FX(>J&d_G\2^gT2>4:V5Z):R45YF#WVG?c<RXBF4PIF3Y\\5fL2N?7=dL;GIT&\
gU]YL7@fcC<_CUL9&I-U\C039P4RH@U3?UgMBV(3?[H3/LU:HMfdEa5JV^V4D&S#
7=Z<]AU,a8=&&C^BMa\SM5bJ./V>5,;YN6PcJPBTB[<32M07?[bCAG/e]Z4@=1K1
9.OV19LfRcDPaZ&](OWHJ?@ZSJY?Q>WI2;bV?Q/6\<-=?UA)AJZ\,2R=N\9;B8OQ
8R9Y]I33+cbS65)#I\R)7I2=gF:I[J6@XUU0C9<VO&RJ/>K8QKNVb<5<g7aZJIZf
e(/,:O@L3Y;7/,.YS_Xfd2DA1I/b7OW@]E#fA.cgQ(SYBNGE?/3]eJ^]4JTA:Z56
g8;gY;7EK])[9IJdTTQI9[EfBSf9>:Y3HAObB>;b5^UW42PVT\aRG3>#Td+ZU<A8
X8Y)TYf;5,=J_>T<NII5T>QL1aK01;9.Vc3X@+Wf;_IRc94g:a^a=7FCX(N+eLdX
XVdg7\+94?gZXb=GdI_&&G+NdOCD1BGN\[]LPT-V2&ONAC@g_H2@C:9O?N@5._@1
5UDe\<\]e\X^\&fE-,6OX&OYWXbV/0T9+/7^2D(=6@8<5N1A=[@H0cQdG6O_D;6U
4S3;FJTIaTKZAMK/<0707I^AL]74YRM1R@>8&O]ER?PVc1\e?/O68W_3[gT_-SKM
RO/E4RDe+=<KL;#a(K<)<,7-]-5QI+1\Yf6Q=J)aYN0:aF2.1VZ@SYM@ag2^XEF4
19BCI083Qa)?&1.&@4>--P\)HU/@eW:\+2ZbD\75Z@5JHHg@-1H=QIf>,+g)<NHS
\?U:-WGN(>\554R5fST6SX2IE0=KJZVY>ESDaFe@/K=ZNJ+4;0XX&Y5-BE&)ee-T
]\5&DccKUHRe^IT[;690QRHQdBF<,JW=0=A4;]cA=bHHV/+UP]R_DEc&R1g6F/SY
c#^S;d4FG/:](]Ug4EeWD]OT25>1N5GUDW.S7N.WGNbHHCEeeJ45VY8F@4R@HI4M
c.1L37.=:eCdVMX+FJP7GHbL<KK<#PDgUVLA-/&@?=VLLb8;BRQRDV@7JU;N[3E,
V9@V7FOUaC^5Q)AF>E6fgO1,&>&3\<P:S(2agFbBGZES:^/B:;TN(NKd7028#S86
9V#AX[]e/>HYcaZM8ZWa@Xg?Ub,]\83OQ0+fCUgFeO?W]dWQ.W;gSN9,.<80V-BX
-gQ1DQ3gV(A:MQ@D22Kd\]VL<IIeKVddH/3M5,VCg\S[DB(:fDT\c?Q?5@UMf-_.
>-c&>K;G_P//6D.2Uf95:08DL69K2<7RWO1a>-MT;]YGe(fZUUcbK:U)?W3_.+2L
dCAQWVUY(X9dMBS)]U:L?KPe<6Zg>I6Dc\QbZK#Ef;;dEYG@7AG(MZ,+Ec+/Ea,X
+L6?YSP7#T?.=?5F<\W_IPB2d18TH+(EPHE,0a9NRI])#ISbC)+VZb=,\YeJ6_.T
,BT#DfY_#;b2+O/EF@X5S?,N8BaH#]3aO^VeagQT#Sb&@U[g8MQa&J#MH+S;8N\d
\Rb(J5C39J+RT6AQ:2UIOEC437#9Zg_(Xa^E0BT(V&+<):O?EfCS[@aOD0/:R/>D
NEfFO;3HMN4cf4PR3C&Qg-H=V&6,;908XUFAHa>V7E0Df.VTSP_?U)F<&cd&F3RH
I(38ESP+R7X.+3&(R@A.1YacR+(@1eFVKMcQR6gM?T8WLRF:0OPYYO6=N5Qa4RRK
Dc(78<E7Rfe(+QN,>L7Ad0\VMUe>e?]RK0<B]Z-8D?4.O;Zc4N7GUA9W@Y2;DQ?c
0dX=6?QJ[[Y[X<bMQg-BLaJ#Da)()Jc:F+2--63MIGE=T2<J,[GYWe;K9/O3LJ.e
ITXB)^]1.g^O++3I#NDbd6.^,>e(&I(.A)(QFK.OdEI#G^PG3eDX)eG=S)0J6Z1e
bQf9eOa,/0J\&_>V6YAOW3TQP;NX^/TQ2+Q[Q[6eGKQR_JNUJEOGGbJ[XLM;EQW0
I]P+-QUe(PH_aZNJR3:S8+g0F>WAg&L-&Y2U0V[<W6)-TfK799DITcM#g;SN<T8e
)GbaA],;C=++\^8_01\[YJ7LgN#X.-:#6E@9dJ)4e04c4\0b;c+g9-F7W/PHd1ZC
Y3WA2B@]0W#X/&XcdXX8#YeVZOU>+?Y^&F]-L5<YeU\B9FK27[@.1JVNSPa@\=W^
5U90@fV9HA\Ma,O;TTG&/KLO=FF5Y&P]8(aW#71f-OUEb_NXYCZ7P2+RV2]B<F,J
&dH&JJ=H-P+5CScQd9ZGM+[<WSY)cJ.7L\6DeB>HSNBa/YCW06F8;ET6FKES2/TS
&6OK+cE&>?HW__=J4+eY/O]3X7N]a:-LD5Q]=GTegN4LGKVF3b/_A7>0-,LFgO.<
86UUXD50D&@:?M)BZJCFV/MVD]H;N2fb2:0Y2F-f4:UHF>Q5+A0@7:AA09&FBT;H
)?SMZ_OUB]Y?ZQ?g-]YLMXV5Q7M7d6X^a,c,UIM]@:TLd;M\66LW6\YU[)>=MV=S
Bcd>NQc3X1dd0>U.P<?V37^E-()g&Cg)a7g>+N12^4QTP:><_:gOYQ/KA#TEH(,7
--J+9,MfB_+]=//K[4\4&bQ86GI:7QRNfJB59P#NdK&5ECXI0P9XdgTVR[IdN+df
V9_SY>2;=c/\N^^KG&MdI(W(PH6e(0f<.ONR/C1-O\H2/4N8:9J6H=<gbXYBEEXg
Qg#MVTFI@e[G9U;5:=@]?I-0QUHbT3XM62Y9aJ98?L^,Y8a3[9HY9Q;_XCW&D8KK
F+8CQKPc.?/4#fNZTEP3V@Ub0Q[]4RM=-[)=:CXB58?I63VMI@a41dNJYW^=\2\^
//8B<9SNF-Gd,Y[_,TII3d6CT@5OC?F;>=\-LfN>H1@/A>,X9PKO6@TP4[DZ9\EB
^.cQV)fgM@R]XU=c7<PcIe3R7gCaQN4NLDgI=@)QbVKDLJ;IKF=2DAYJ<-,BHH8G
L28dbOb-I@SJf<D5E=:2++TMBR)VWFR=&W>+G]bUf#HB@42::_.-\a)&;SN7<#Z,
Hb9^^JHD6,d)T\?D=gPR/&XCUYJgEb:ISD=,[@=B+aM&+Y,MNaSZ494DU_H0T,F5
^O(M@T4^[,E[-dcaZcKfUQ(c,OZO_5ES,82.0D=0BHUB36@EMP4ER_UTOG2\dG@b
>gR3b;N+.#\I8Q=S;>G_R#Rd;JE@T^4:1g>(,/^[#[LSOKE<a_F@?bRJS/H.9=56
DU#g;\Z)NEA/]T3aI4Hg/U<0Z5SB+Y[YfKR0(cL^8dA/QcB#^5A5S;)K<b^5Z]GW
O0@PX,IW6W1cdd_7gWKZ];).]dGK\4(\Yba\cNF\.(P,]CDd<.d>4Ke6CZ[?-6>3
Z&0=33/LT3[D@\fM&DNE[,VRY[NDeR@:BENd^X5;_bWGga5]),E>?U@KD709AZHR
f,<PLK=?K[V>ADeaZd#Z>ecP:,.3a/#gCNGCecA>6@<CGCfUU;d\g4P4XR^T^H_5
5,U))U/D2dQ=RaG6&:_eaW9&XR=#&1.O<\.@D\<eE9)===FOXHW?&-L5Q(I6AJL0
83LR/)]=GK^<)X4/7Yge^DTB?RN]&-bJBcDJ^W/bERB\YMUHWO-_(\b7M4U[0Y<M
G]K&e[^8-_d09[[.VB;0#Vea/RI\EPfAWL^Z[FSN_RMgP.,#@.:8SbU&CG,);Ua2
6MD)\,OT]88>AWP<;UD?GOMGED/6&Y&a5A(Fa7AbbDT:A>M+7TL:C(Yc@XQ\9<.H
<@W9Q0W/X>MP=EJ.KS#C8FVLfGYbQM]Pg?M4AbXgYY)=/4[?0<.5^WUL15HbB9\[
FRbde=aU0Y1f9P4d#MI[H;=QY)MW3a=NHYMfe#.EJg.cEHN8gDO>Y5PN_gGdEc9L
UD7Q\KRH>X3b,WL?I]8SFHK?_H22GOLd=85NAQEe=ZWQ\Sf(P.E:_,WMJf-cXe_X
-I[.LJ+?GMB?D2^9^_a94\5W_:3_Z5fWg@S=A9#1W;@GH=c.5Ba<8G(XUg/,GMaU
+S2Qf[<NZ;-A9D+:I^FV0M,PdJ.)aUVcP84/b?F0]6H(I=B77F+EG;b)VN)4NE]3
7^K1b39L.gD5#;NCF02T@6KM2)X06e^MKQfS]K#<3UGDZU2f#F(a.WG<ZT3ZH7EC
.S&WOBG77G&MARKDNJM&()RY?Jcg<]HI3RX;b/46Ha,]V07@)JE^:V37ZGaF0WOU
_8;b<aa,#[^5]OW\c-.I?X\>I:CJN_ZaRNH76[O2+Zb@?\]DW0P4#Z#CdFL-7YD3
KCHZYPf@K>77RJ-AdecN#/B@+&c+?WR7V-&EPSdJ8.Oc/PePPf+^AJ9,,7FTES93
EA]KTVFQD,:,?M<Ib9[Y2E(IM7.]#d9PEd89ZQV[1E-4CaFHL]WcR1F\0G4H3fQG
cZ)UK(UM59Q<^(<@^2Y+H.bCf9PB3c2)S5aMZ5/U?dYNF@.OT3CF)>+;;G@[7[F/
YfIBX=)XcZ=/.\V[-9b;eSTD7-Zg0X6;KgZ0.0:Ue#[LX><.D;4N](-7>\GYT.B2
_D&454/[88;(\2Z-KAdQ:U;S[YP-@.TYd^)[R2aG=>MaTU-JSK6KgcY&;#,dT>4>
PNB8635(P9\3QODJ#.:GSU[O&Z:YNfKc,UUE0K5BX-5[L#DOLaP>7c3BO\eJACgO
UN=+T;M<Ab]H5&3#^@_HH58cZQ+/\1Ece<>I4/(69?7G-V0JYcQ#cO_9?&deRN\J
Dd:6C1)S-N:Lb3gI2T4Oe<;QOC\f)LE_fRV1#M[@-K?@d.a3eMWfN<S)-1Jd/2b0
A>PWE8fRaABPVTB:cVS7@+S<ZIKF,@Eb/H1cJ44ZE)M_8]Q?;eY.=\KTJS>dB\K^
\I/ReOgeV.C&/UK.V_L1-_KTC^ZHDAU5@Z;g@S;FC>7<.=C9;UKI0]L=58T-ReT]
X,E]8#U:DbOHQB2K(@T:8SCIFON:G.3JST]NDC5/-1f#R2B+A>]9L/=FGbA.SJX_
.cS#FO,Pe/#6)0M/PS>R0_EUbZ<QM8Z)VX\7d])@YL[9+Q47daM0[>JZKT2<,5SM
OGBX0R^XCcYMR9IR-JBdWd7\63;VG(<a]b<4,:A++:3).4\@1/+2?->&eUTFJ+9J
<B5IMZQ<&:L.@R:^BURWF:K;^VWcf84^)c&NgGER,[ZAQ5?@5+)+L(Y.T+aPKVTa
G\:J1f(\IP7(FJb9+O@DO]J<.C,f9_dI^0MDY#R;9-]<AbKX&NfQ:;VX@J&T1KU.
Q1T,_M@.H<ZZZ=.PDXBNDG(#O(^KXL,S\@BCA1X[Y660XA?LWZZeg3dG),)&S#:W
#N8VeUa9&5:_&DGQTPb^42X,[;BZ3Hb0:;_P]&&);d)A=b(GG\2&@/b^)6GAWC_:
P0>(H^.@7#/]Xf,>?FEQ2BNR3;2&ca=+]H5/N<SN+/2cRCFJIPe0<=\#bHA0K12;
&;A->KXQ?-\Y-KeU]6C#/H:I)fPKN;J/a#R]0;(2HVO\>JbM0NQ>+K:DRP2)GB3M
D>:e\SHK?>5U,cC/A-6F.Q2Q5R?]CJV+(g?N;(.;KQ&BW#NQ^I(3/dJ^T?f>/FQW
cI\PA4@#dL6>E@;7(V8#^(IL8410ca3[3^XB^_MW?QdD^NgSU5b>GLL#X-EIU>V6
a?;7KX:&?];ZD<,,[^[ba=.U^bd8[-g<Q#Y)VO7Zd>+,2aQCW/7895<5VYPa3,=P
ffYN&SZ=;Z^bFPD-\_/QP+8a_YT?QYKe:VL8e3JJLRZeF2]CLZ\d&-?Mca;+#-NX
KLVW7Q;cGg:MgPNcaX_AfJ?W_;RNPOK#S^f?Na(Y=@(-O98aMO2f9+0#V9_ONL.;
g/6&33T3DKXP_e&A&[46&,:b11UV4G7=C<K.,X8BBLA,C8BHVVY;(S2GLY,gM]aY
OD#GDf#NA&@<4;3IZc9c\_GVJ]WI37GaPbO8;#dP[O(GW[:0X=FIZ>R=)LB=+CHI
CQfE@6C>2[T;04?TGe+9I]]c5OH[6#dbR=4E:OWX0BHdd#Yf#8Ga#FR^4df1,a9P
9,T4IU;ZVN-+P6]>/5c=M7#/+8:JK1@8@DV7OGC^Y[GC2f;gHOK^49.ZbG]G3U6M
9TGY#PLQ/AabZ<^@Z(OU-IHL31[_L+[-g>X+ECbA;NB8@6/;/6CBaK?g[QbG7.#4
P>F59b\N#/(J88dAI\=IJT@XICg_HV[D2<b<A)\L6PWY,E-aeK]YYNCRQ0Q[eC?D
^]]8QPOg,UdS_VP86+,(a[)ce4JEFd&@0^L=3R-40K+:L.LW3L]3CW)]#7>d[^UQ
eQ9PTLIcFUC.92PHF.BfU>bbCPY:0[#]g^bBBO&)TaR+0-M0;^]5M1PQL3,IcD]Z
H_9=I1R:g@.?<;b>PKc.+eKd0Yd@42Qg1UdY7-^gY_D3fa?f-bO8e1Uca2F@Gg[N
fP51)L_IbaO.KJLa<XI[SWYE\1OOM-g+5V4#?dFRf^^@LfP@?g73df3a?21fM+6I
4T?b65b4BOPbVdYQ?W92]W?LUM&M&GW01_<-N[65^(aP26L?ES.BRf_/L]FPAaIU
O/C;#ag[10_<_K<]LS2-B9gP#7_PgHf75_79R_#L_D0V^YR8(:ddE(K;\WLG;TK_
LaT#aAOY02FH\U_UI:_fC[93L//_)E\+#;Q>b\8-8(d5(8?M.J7W@3age\Y/&9YF
;K<Ze:[NU@L@fA>R(Gb/+#cWP1ONQP_/BO,^Y]/YF-)Z01+BC86&.XG4;eJdE9D:
+^W9?:,K(5TaP6Z\90382E=FXS9ADSeAX#T9<K57VYT=^2MM7CFDD5MD3T3]&)=:
+^W^HXJ(@V>OG4-MP,fY,ZSZeU/d_TeV:OCeA.c7DJM=LN3^7YT6XDf^,-J9<2Yf
#C,NW7g[a:2:YT=SM801Z15#>#S\_GW_5PBa#CALFW#L/+dgTO6>52W^=Ad([a6N
RL\0BE/VG>CTa4X/IgDC:6])Xf6^.LXb6<C6<W(0A7C2C3,PUYa>P/H0R?Q@Nd8[
GMJJ-#WXV0EaTS27R=bB(<JLK>6dLe_@VANcNG,-S:R8IMQ:b\0+7&I&T#CHO>0D
-(b#g:QQ:&\c8@WVb.Dda-QL8MA0P(2,abG>cPM@#=Z&IQC_@NV5VIY#OLM+S8DT
AF-6NAW]^<ZG.BEHLQb)5>7F(R.[OTGAZ3=1QfHMW,W)>/3^(<OL)CYc-ETd2HT6
-6;.BVGF2S/86<9RU(3K@@.aV):fB77L)5RHZ?gE:8X/W,Z<cD7U<L5(4QIEZVM]
[;EYK;>g&86;D(\d)7;eQB+=gJAHVAP/+PC9&UegV)DPW5Z:D@ALRB@e-a74_@CV
ZB?:TL:(1ZXISAO=fXdK>54c<aD-D(>TU8YGDAaMR,BSJ+7@/+W=gI5cLH(;7eS5
cV<D+]L-:J-AHP8B,<b)PZ::8V[SOeF<?<&\UV\4103_Z(S..\7;bZ:+/SfMBL9)
6RT)OW&)eQ0eL5Y#H9RP?XTO&9FR)gYW;IG.VVAeI^ac7T1DEI0&(EHY36)@,;:#
D<O>(H8]6>aXaLf31TgTf)0LN73/>DaNG<X<gRJ^&ZbS6R&;S/?>M44@1_B^W;J.
abX9&)Z\#13>GU6(DFNS6+;X(.JPF3TcJB:X2UCc^2@QN06OS<_\&bZRC3)<4]Ef
=1)2&dF&fHQOe4NG1+Cf6/6=8@I\C#XD0#dL_-@b^90X-WKIO:;_2gePd6_W\^=/
gbf@#E.YAI+Cf&+HS6RN;M^_C>ZN;\#U@V=27RU?_8KHaZOJ0.g41VN1T(0^g>A#
&d7>B2d<W:PIg_W^AM]c8?)1KgE5&N6@[]7<53U;LF^GP/IK2,X3UT><S=<NN5C?
L<WZWWPZ,8^L3Ka8ABaVW><^6:#5MJ);OfU>G,dIXGK.J?&RPS@9+S=6M^K->RGV
c>]L=LX83BeXZIBTSI&/-B-;57EAdM+;<JX7ALaSKB#FWG5@2X^3R0Xa87gNPe#.
a+2,QID23eGaf^S]bM,a&+V\\LbCFQ\S_7=2,2+5=f>J97)8A,GeT)\]?R_6:786
ZKa(#ec[2Rf7dOf7dZ.&2O\d#ZSH.0BT6#(3>JWT//]Eg:dE[I,SEGZVe^acD19(
ZET5I\PgRBg&@f?_8?J65OXU()9FLJfL&gQb>?C(:g(8XKTR;a^LY)T=FAZ2EfdB
a7ADEJ(3a[]>+GJ:T:+2<PND49PMRR12.9HVg_A[[BUBf&dfD4[IV6\3+Y)\D9&T
.RGfI48?_Ud^[g5CIBIPF<4_:+Hc_Qf3=L/RYH6NSL<E@T3+>fH?.T#T@)N(=T>]
?Y3BC47U>COBf5<(><7fJJKUMc;/XN.a8[0(\dUOCRMD0QNf-7X6@1G@WSZXL20U
TPZ@Z;ZH)KF/c&P>J8A9XK<=e@Z.L\[@4V[2X>Wb.eJ,Lc^cHgOa?2>W#XET3Ife
IVIPQO4DRVXW+N)X3Q#IMT9[O^WagE6<D)XEESWO5J(fM6WS5M#NBF9#H;-RV1Ia
?g<QQI21JdVFB?&6<<Xdd1RJ+2_2aD<AcNJ<O9eHG;FgG[)gSE.0)3bMU(\_g,H)
1O,JGgD^@a5<:MTL-U7fa3HB]GM7dK,D<4F53HB\&:BKYX9Wf0[BY)CHU@(CI:]@
U2-.@0TA)?eF7Q5O?-,-,69\cFb@00g?3f_D&DOV1Q36A/==+)0114[]VAIM^=)&
/J2OX=F&-,GNA(P_UZ?(S-^<B+(,3QP;ZDQ:g]g>+4S7(MG.gG5F_AN,[WN+NY:O
ZUdX5[Z8eg<YLG(Y0&c/\JHb0ZD_aE#)MQ(A1/LLef3?;Q10<I4[-H6W?:EV7(g>
F]c,I2eLG_/?;KNE]:E]dJ;3Z3X);\^NSXgg1SI)OW53OR=]W?/R\I<XY7aMF>Z=
?/&E8H9(g2FNg@gEO32/@KAec8X2XOSf]MFHI\+eGOH4SG##VM>SVaC6V.6ETS@M
)M-F?QA;cOLJL2d)HTeGcHLN7/TV<R<Yb?B[2VF=9#:CCdM4PCb<X1+K@.\0bJgJ
S3.XWE:0SL8DV[_P(b_WdM4PN[J8U>;;J?\J#ORW8HPM^c9=#ZQ>c.#(ca[,ORTT
Z7OJ_(/><,Lb7P=3L2eESPTCT:A;,#JALGX?12\MNQKL[F2K2J=Qc5<I#?@GL6S#
NGE;K_0a.:=QgHU&0A#WO\Tc35?(F4&YPU=_4@.,(BBJ6^@I-dLJ46A]:/47UJAP
Z3[C^;3WS2B0V1N&[F@2.VW]BC;IP4DbPP]]\W&HEP9f#XYfS&Y&M9GM]+e&D20)
eFK[)Ce_F^MWH26&B\M1L/5cX7/7-WeVSR,d#@]\TOH=6BD8S[N,2)0Z6SBSV475
2>KMZ8cYT.ASBC</NJV\eU3e0W8OJFa5\Z&Ce<fB>2XZQVYU[14X41LWDeJULP6J
WNMNgTP\8f0OC<O18d9DEFFf7<I60:fXd3&Rd2T2=I,&FgSDA-[NB87EHMJ;,,?M
+QN9(3XKVW5Mf[EI^RPf:RJU/c+fIA3SF+3[T3B^Q;?egYFAR<XBKI4]S4LXL>Va
c&[,e]Y@^VT+L7SAVfP1c9=?AC8#TVR7P5AGOVSF5M67=)/d.[RN)7.:Pc<B32(2
I0Q6GN[G<LKY1aYS[6B&SBOK\XSGA;3+X&6c20K#ZT_VU71AAXGf0:Fg5R5M8DW<
ZZ-ac2XK_;M#=dTCFcA:U8PfFDNZDDg1:W+d)GU3X3=1A<c9QM)UNZ)SC)\YQY8+
[<;?6@&6O;T@LDYBeG^4BO+,K&3&SG_5QYX^\4ALQXDV-XHVc4[T0]B-4IQL&MF0
<5@bSg_J,YZ,<G6[4@_+&J#V#3W?LfG\NSS7C0P5++NSPSbHHI_B;9e.A_H5/A]5
PETD;-^+aeIF3P7N8EIR]>e,Je:H?-46N0aGUX(GQE^JN9IUU\FPT1bfY1a4_5J?
/ReI=^N\S@H1.T<M)\-U+9_5IJ#5+O)0250RCeLA2[7LG_97-W/5=[.NAIH8(;X0
;\b5P8)=gcY2(Ff&If<Kf\<8eA>g=UA+g5Z6RE&DT)D.KS\_aY+XI;-N8R+:R4Xd
eF)Oe6L0MD?\g(C)/c+;OP[?bM-KE&J&fT/5>5I02?/])DIY^+Y(B1Z6J?Yd+L2+
#a@_T023HNE1[YOUDaY[4EGNY3-MV9]XU/aV,HQ2bW9gLVSfeD2V]PG+_:c/)04=
ZYe[UUGSbXZF>Z_<-2S[1R@NUCQZ62)OF[/[HMd[aSEXCCaP(\T[A;fA]7f3XIL9
1+#&Y#CKRfIL^L?SAa,JV//aZ_+J2fac9+]ZVDfb5))0g>68/b=2PJABYN3f.E>?
dC.QO</8+A)f/AP;H<)MM8BQ937&5HLc709\6_4)Ue.P7Q^CNK\0O5W6WC<#KEE+
dCA,]&/]M9e_5+XL;1IE^WcZFV4Z+1[3fHSL;Y;Re]N9@4\#bR83^g)7DJTL>;YG
<ZEP=T[L\Z9HKW[FW_G-aSM)03AWPA8&&Y4<.2DR[>d=QIge4Y&QB9G,^:B_/WD7
cDV>T@_,gZTJDFJM-ES3f#Q5PND+c),?Jd3[YaN=RA=(LG/>OGAKW^9bW_?SUReT
#:,L97D>c\3F8OOa-YaAK0NaJ(+R1A@C=.(+])fX/b^&.Z^c6MJN4-.9)^0BJ?gM
EQV(G2R)?TP7ZaYeQ^]+OZL0/dDEC,eI)F8\=5Vgc7B98TJ-.E-;a6[VO&9B;Q7<
KCIPI1M]4=<Ng\6OD5/fVO.K2NCeE[5B5.(ZQbC)@QMCTO02BdcF-BBB80JJ(TN>
K.XT(7)C=AQIQ;X+&8gb.PW@&dS/UXc1T?2BeY05ePJY/N>:+cT?GN\<=I1)fF&G
Yb_K:@FQPZ.Abgb+R1L,J9R^Y8Y8.cJL:E[B]WY3+5CF-E[fIP5.aEIe&fLRcNAW
G?)6>,&(J_aB4P^B4b8B.URMZ\+H;.,O@OP3H8Y60)4)DcAGIA)=?GVK./?#N6<N
gWKJZSa<1PeQ?,_RL#);P&O7[>_=gC7]/J<RKDRT#-.,-N7f1O2+/\9AXO-)&:X@
>?XW6bD,O6U5gE7QLRYUJQF-=#LeAJ1+4JLb_e=GG>ad)SIdbb0Q9Ra0--#1S0(7
g\P+7@V&Ib6R#D8+DKKUbBN.I#9O9I8dZ9A6d5&Zf8bM?1,Q_._W8F8D(A1^N6E[
c:E^L@8d1KYQ)&8]eERBEB[JH<E3L&DT;<N,<[VN<[\0R8:,7\ECTN=SG4T]UNK;
<NS4X8+U.>N;-gT:4,N;YIWNY5/>+_KQUT5>Q3)QgNZ>@+MVUW+UJT4K7<:LEU]8
FXI7b?ggLO7cM2/&GcD-e_KgIJGd[RI/fZNRVGX7[K9/]cYP#f(JH=8Hg]7<-H)P
O/4U(2Q2<GH#QHF9B9J#AVgAJC5Q[UDERPHXU-R8M<LB>0N<_E4B1(/?e,@>SZKZ
AA@HPPT7W<LE8[YEe,2SL^c+V,:=fOF/R5J(9]Q?f]E,SP]e<?G1GR:#SIa3)C1<
];EEgZ&OdW]+:d[V9TcZ=P]I^&N>7--g2H0P&QJ&VYf6aE-Yg1;[S+e&;K6V,X.@
TD+5I(.A7F\Zd2UCJ1S.9(S@3YDM9=K9[8:CI<W?3<CY3dK?eWY^LH-_U3>O?VF7
Y9_-(#H#E/)VYO+]QFO.78AK<2QR\9\P@3X+0JYHZf79NBc8XXASUQ2eR[Z\(E]O
EDJL[>F1#Q3AZ=bfHE1;JDBNIW:S2bAZHAVBOKXL;7#33e-FSR^\L@Q4Af>I];Ad
7Qe]fNCKRW7UHLGA3^U)+bF7_NE[2C#dY]&;^Yd]Maaf8MX#8P#C]\:>1DWASVgb
7L=fC_G:B1VHS>BadH&T,S:,&Ce_#,APPJLO6X-b0XHg48>WXA^N0I4MK4=0ZLNb
X7IF8<cHHFd)@MMMX2(<bQ0g<)6?cTYGCf;.N<b&5V9;9-6GbRPg(1YRL-L5dT25
eK9WE?DcG4fR5Te(Z#;F29<(c-#Z1N;2JNWI2YfNJBdPFI#bY]]a31S8cC?(9A9.
dFV6[\U0KVXQ;\:X[KCe23-\5X6=1A-G?-QYKM+V\A&L@?SPAV#gU_^Tc9-CB[QW
A/?+M?a<YX4K8dg?(SP@)JAQOY#9((?1HKgI()T,8(:2ROED#7191W3Q=RW7[X1e
8&//7ZV;F;5d>#<&,6P+MZHT6?B^H)g[<,Q4_[XPa^61XF1[MZ@=eWeVa=7=XF8<
^M^?J,HI=]8)2^56KU8f7c>cTD)PXf31,<fW0)M\bK3MceDZ#Y3f:;87fP2DA,Vb
<g<V75XfPA_d2YIWZBUEK[C99/9>YE6-F)/-&S00>T69AdEYC/^2/.R:O8;FYe^<
Oa=W#f\;:fT.=^-;YfY0=H<d8,:?)/b+5N[NC&DY9EAU#1]]TES.\J#S-W.CcT/S
EME+?6^.#O5S:8FAGHf<XVN18(<T;eD2<1RPdcX1LZcOI?&(gSWDUdNN?OLI>TBV
aL-UdWQR-&WJMG&g&/,ZIQKD6H++,>L?,81:9ST<c_KF2]Ue\./,_c[1-TA,XL)L
Y3/S64#C_J]U,5&,XPDPZ1:&W25ZL6RC:B)PJWK_C##A=H:K:aFCXL,X>JLf+CYg
fT(a]fRG_e\cJPC_>3SNU:Hd2BK)C-]5:ZWfK]KYDG4:=7UN_U=Y>T(ZCQ3;#1(M
XGg]YVL#0V-_TN^E1dT8g3GWd,eN68([/g&cT8]K5#=:)Uf+eR[gK(1#,Y_a2eaP
C0W0[(706cefMg1^a1)KXLd@WgS&4Hg+d]KT0-cUFZ^Ib_8Za-C3caf2,13F+XSO
aDM@UY#)&a&J1GXI6GVPK_)7g/R)==YSc(3>LAL)#J1baMT#cFN&cU68/HSN\c-?
15,)Q[?&@,;GObcA7J>&K/OI<7<Y(5W;C?b?YTJ^ZQO57]b9cG+Ud4?X[bJMN,AY
U5^UZSeRJeGR<K5Q^R=22#\EM-1.+Sd2ZZ7@@/J]L&KGRL4]LEE3V0;9a248X7/V
[W&TGJ73^Y#)MY3[.<:#]:CV4R=E^#CQFQ2]bD6^/S&Y=d.6+8R[(,JIZGX6ZF38
5-EQVR)<dF2_-H@8bRb7L@.-Xd^?.6-83X1-8.6I:AENCUJLW6\,NZ4A)=d9>1<N
[:1ND.>^c1>LDCA>A?=7Eg#aR\U3fJU1/4b;#fHY<X#2,=c?IM5(+)#HO6J8A)<e
=9fT0]:a4YUeM+WIT6ba#<&8/>?UY-29^/Ec5dAaX:T_MIH&.b0]Q2/3D2,NUJ.-
0U^>HQf_2e0\T)>[a/;OWRSYFU0/#L,AcU-]<?RP./GD;(_:PU<[aeCH2Pa/25^O
>^/=<@R,(:?BWO[X#.f0PeBf^MR22I;\)fNS7FSg;WWgdV:CJaBA\,V]<F,-Z/+O
.2(7?^U\1)Q\)DY9a6e:W>4?U?#_BZ^S;#&cQ/3AFIe9XBB7c>>=IQQ2>JEOS90S
^QaSeC]W/(8cQ>G7#.HH.4\FOg.Ubaa@N2.8W9Ga6HGg.>T8H.-&,,B\A@?6V4Jd
VLIKP>JU?M+\N+/BM\eJS.LeQV(^Edf[PRfDLJ^_E)#b>JY0Z_^d/WQPJW)d\EeL
Q[L__&LZ8:d19;U=1C0210GfbL3W-:;AGO[&f\W+K0,f0&>Dc.M3=C;42HT;7#[/
R/^D=LYEZ^P)K#3O(;@db:PCM@FSL.Q-/)97(FQB[S@J\;cAfL9J8H^&.P@4G36W
M],a8/-3^g/NN1EIG9@L:UUP\J+f@[A4:+[?BX_.9,6V9;S<KW,/fFH1dC4F2T?C
b6Z)gX[OL?7dE2M\93(6PKd^Y@QZJa;P.[,7a7EB_6Se[?#@R>6f&,#_MFe7\&JO
T3d0:PE5P0KI0&\c08aC<@6:e7_]W&G;aZcF3K+#(N3ZJ@_U.?5;L;NV?GTWUBb3
\c8S[NFB.ZU&D#,)[ESg+6/MOUX1g9@]NaL.f_7<bP@g5[.#Vb2R@UR?D6AMa&E-
d7+P,4>+R:#LWR@Q&ee,Dcc1(Y8WVeIMMK+ege<)4.0OIA4gE75S9Z95.GLf(MZ2
d0cPc;CG?<?D6\(a>^1=2AU@,<3B0&@.6ZL6X8b<C?#gc2HW]cW+_AaT8#@McC>,
.Z-,K(D/4:+]0(?@B#5P_ONd@LVFX@,1:Je[K3@<:9L0Q-CV.2)OXI9#/OS6P84=
c5a)#ITJ6)=ZNFSed/L<&aR0GP^,F.fQE2O@A,VW#EH1Ff=/?cE=?3AZT2g/g33d
CcgA.BIVaFJEAdBd)N2_W5EIc9WN)0dEF402YATQ)=6OT&9Y72d=W9_RN]2/X_(M
X@0QQ7bW/:9a4N>^=TWZCMQ60()&E4.T4HSF?(JK:BQY:M<=-@/gX=-4EHMe=:5g
=GGTQ)_ISg?Bd712LT2Z(IWGgfP6@CZU,L^H\a\13)/3=_1+@,MA@gZJ5;[1,O;U
TREZGH97ITGDI]6</-gWa]XC?0L=TNYNC+3F)WD.fR\QGJCBI_^D6PT_C^[-Z1Ye
-C<DW8ZP>I]K41&2]V-+PD1KH3^1=(P]D)0B])fG7&D&RZI#PR];]R?b?X0EPW;M
78_VU,NZK0GUJPcf\,YEZ-G7YJ3+;^a##2H;<:[HM=S.RK?BE>+U/(0/LT((WFK@
C-Q1AB]@b=6((\N>N>)6Z5:+DPJI/@AKSB+(?FddSeV-]<+f90>OV9DB7P(LBRVE
a:BRZ-X:/R\9D>^C(\UOOcI.M,g#F?=/F#.I>KbCeLd:9Q65>\8>D#@I\64V3+X<
Md^I-\0W]^XdSUa>;J;I-O_bM+KKP-V)>c/?/VR\PVFM@g.@S2[V1#@F[4N+C2R)
g0;0)TB&bSa3<0\I:GEP0B]eGA\Z;^L-RGaTc<[eRY<5JT-.FaQQK<&ZR:V_W0=Q
J)DJcJ(6>FP8aHUT6N7=fVSAa]I+86G]<CC#Q.XI^D3,cU3:XC3B_D>cfBH6#+A?
LcLU+2.E(;1I857b4L#](<N@61L1a,NC^<.E]CfE>0IE[XZFC#Ka=?TPH08F=YX?
3I-#P?Y)_;X(F16@)McWO\NO66N#P4R]&SRReR&+[OX8#C,>b+FNgM>S9_cE<;U6
T[&L1c_@SLAXE6GU3H;0P;PL(HMX@:1(e(a#62M@^GMW#QY1YHW5.]g_1N^BbSP7
Jb>a@(VL/>.I.<.:KZa8Z4S/G,E@G,J78A;@[.c5B2>U[?Q^GWAMfZY^K(A3#U@#
,-+Cb[ZMGe8&KIF5X3WI&HJLLgUA>Hb#^98[;L\LdF7([3bgdg&&H#XE[+A9#Z]P
fVC8C-85]TZ_RDcg^\7LUVJN\EW6IQ9?E=X9aLEO),6I^CgGPY>Yc#/:eGW7<&MA
)LH/EDeOUH-=@cNS#5O10@Pdeb[\U+8R0<TD,_/fN8XK^L8_.V;7/U/+B7c>FK[R
I#>Q,>PB,UGDQf[)AaY6(VXW2Z5?)CY@Y@W5;)U=c]F0,N5UEAHYd43YDQ#aDK-G
FOIPKVY35-3MA2H(P&Ugd?BMOfZX(+C,=PIC;_=gJA,)2Gc/Y\T#c9>C>LA7]K,O
UIOP6\9^\P/_c,/38FF8?X#e2.NXV]5@0T3<DW1TK=YW.,]+\g/3B[QY5V1#M8Dc
R,[?LZ51HCBYI8Z?2&.V(M#I8]:M;&WBBO3JZ?I9-eaaUc\^AH1dHIL^6<[W+TgO
09UY#VM.+53JP)G3eBV5_F5+)gD1F3I\K9a.,FN2_SU6J2(YW)=,CQ9S3UYOYOEI
C,/fYGaBOR+;+LCN?3P;E=U#,WI:.M[U^a0_OHV.:4bP6,HJB])VCYGe#(7=^Bd:
9E\M]43M@;:-_ISR6TcDNAK8K-?Xg=NA9[X]g>X7ba>H_YJ879W,K08WWD-,(7:b
-+&>7-.()X78RUD3@LcE^[^LRPNIL#gCGKNR\(V=T;0HX](YOUE4SYfM@GV3SaGf
A.O>52RaI=7>A4E>Ma,E(71P@)TK4A:<UEXA3^#7AbT25ODZU\[>\6G6WMa2LKcM
&.,#D?(.;W]MP^0fR4(#gL(-AF5\2Dc2-)Pcgbdeb#XLM:W)Q]49_\E5(:8/O:\7
36BYCDF3H>dW2XUQ[<Z&)UBA&[:L=_L[RI2Y-G(^M=TTe4aS=5C=af>O1/W/1aVE
;)fZS\[?cL75F[UE1/NM/1+?Uf807T8#--8PcD(Y9,PZ./:6OJ8131#cc)gLW4=/
a4]N)a5L7KB6/c:A/dUYcC76N-O:(Z0JcA81>a(>gP9S3_\KK=>E8=UU13eNP(,P
NGeBbf):Gc2Y78;URRGg.BL2XKR^PGVU<CN1Lc3EVGN[^V\CGa5?,7U=;:,.XYdb
ZA+2@BTQ+c;H@]YXcc<d<cAUaMW3D;5[0FY2.a?;07[HRe4MdaX(;c)[^T6+bL_)
Q[(NP@=I81F.0-Bd\<O)6c,5cTB;8L77KM>a)RB.VA34H[bT95WLA0BIg\ZEIQ#1
&MWOaUb?YMI6Sg(@9ZMKAAHf5g?FP7JI253&AfXUG&I(B=d/&0QQ81AZ2)a&B,d&
-_P1g+[K7(@aeg63?W24GH5(3KTdebg+N_T2V>^BFNMD]AF/&_)F]U&.2[3Q_2QN
Y9\HV58=N7aAcPZI_aMf(7gQW8;;FT;?MCS+:7VWVf[+4B[X;1D;N)N(T_aE9UeP
d>\6&#Lc?GG[VVRe&G>TIR2AS)IdbX][X@]/3;SfO.N,g?RNS:.NGe5>-0_Pae:e
Z)g\E@UTH6G@&QKTN(TT7ZSG8^YV,6d]3<C&?dac&M7([V:cf<(NWT\1AF\)b,A<
dW[4(eg42VZG8;K?RF/,5R?&d3;_:5IedHS6,EbOKISZ0+R+;0d@fGSG1O_N<]\=
)P.IV&KBMQ0HS&8[(ZF><149OdI<(?bf,PARL]\Ed)<_A77bW=F;RJ_G9&Mb78,\
;:/&(Y8]RU?e^IX<W_W[A@,CDX5.X^K)TYJK1RBc3@eE8?;<0J?;,G;#<]8JTV(d
MF40D-6<#0\:a/WP2E^=aF>:^f:+M@#2Je:FB;YH1We.;FcF<23>T>2SQ[A3g:&-
bF(SO843bRbN,-TZ_P(_0;>6f<U9)F7]F3,:O1Rf?9>X50XCL\+.LI,-O[X.[\07
P=W_b-g3,4a,.;@&9&^R8SO]6LC#/+&B\L3e&B/f[4+fd]+CZb^ZLU[PSA<-T#7Z
4Q_MN[44B]e03B2(IQJC8bU&GAA/>-Uf.bX>C09F;c2E8L_TbLIfCGWYM9&AfFL:
Y)2?M^ANB@c7-[N#QcR?QI.<?1TF>L+<6f3L<.SK18,_@+e1L>Q3?5S4W5C5HJ^?
_MMW>5&GNgD2(9IX077IRDR\YWRWOUXd<-RWP(eJR6,fdAGQK_=P&K0cDF<>-Jg&
QU.Z]54E^3.@fg^+=H]R,g?d?Ua=/_427H1OIA5?_eS+RN;N-:>ba,MH&:CA,:0F
NJ&,T)O>SIR0]fHXfYf>=DA:;+(>+>?8.Bf8QLZ^]KOe58;gd\b(&/d9a7U=CC^?
^):MB+E21.<S;01MR8AC_=GH^=#Ma@/IM<:#B.G\Ld0Q#@0_AU:Z;F^7dI69gb1E
8[feA8H.?39#.]T8<dO1>#ac_If^Fe+F;5)LI/O?<L#[:]80^O>8,6A71WJ1=WEF
>b0C]HN@D?G6:A;f7#a>#c?IebM8WRTb+gG?@WH7UcE/\cS;gV(CPcHcIK-7#<[_
0cRN8(Sb5NBGL]0gQK39)F<O&AM7&e4DgB-<L+G#&V@?=^Wf-3?ATAJ/X)3QIdNc
E&KE]&,Z/#d)\(72bS_2CT4>^?Z;-@H?F7cPF^<aR>U#@LCcag11;<DRbN0BOORT
F18O)#AcA)WQ&@2,c,WgUY6]GKCW+-M#1Ge;M\[6a>B0W]SX&MQF5DEO]c6ON.:(
1@aQD>gZQWfeIV&D#31f;&,&_;GVZ_8EGAYPXA5?A7<B;B.g\-YfTf.+DF3Z66Z_
MR@.N_?KEZFUW<02;TIc@I9NeU.RgQeIV?\=E<_JJP=4;.=_[_c?RWS[3^Q_/Z#[
NG.cDd&DDZRG<5a;UbJ&DR-d8>TCN@Z#M0SB^W8?VJ96WN0)O?4Cc6L&?[ZR#>QT
H)=/H:7N^?IYdMW^I8_)fVYf=-Z3RC5XVLZeFVVba<A;8H\08D@A=;]6UcJ1N]SO
bfEH1@bgg.Y4(>U/L9=8<T[dKCZ9>,;REN:UMTb&TGB)PSAefF>_B9L9@JA2OSDY
=ELKZ69R]:H\bS&(8Eb9U-1P_C5/.I0?LgQ_]((9K^7)HE)F]L)FbCa9K/K,eO]E
)4@DDO?SJEG4]c[^IX;5U?A#+(b)T<63N.?I/<#b&C+P77<a<8eK.6R:&<b_3AYC
1>RF57e,]f<G49,a6cIGR4R9G>+09X9_9[/gDH[/PbEK5TJF^B]+K0MX@)]H4?3Y
e.8:F7L\a9;KXM[S6=US=.O4fJXT?[W\8+GJ2PX^dP;-]KJX_0K&S0:1SAYEdUfZ
4F=<\V;<-^8TN9V/S2\9W2]N\3F^_\CP5YXO+9=7&6V41\NT-K[>]@gE2d([(bT_
8D.C[ggE10_S5A6Kb8V4+2,(^CQc@<U0O3Uc4EJ_O#M.3<D]616C5=V@P+[9IOc[
UaVc\aY;,]?:HbC#INgEW[=VeXBQA>W;:T\]&1eG_9,bMI0RM#6ANcK4T:SWHKDg
T34CdKgB)NO<[9Z+C8XEd/VX4Q^MMW#Ed+XS[Bd\DI\:D34NOZJDaaH/)U>:a6cD
4UHb)BJLKBAH2<J=DWO25][MQE5\S2Vc7PIS.gS-):eIYTVPR0\01;O1?WQQ_V]?
TG>C80f[31N?=H9(DB8&>W(f]?-Og&JQ3J7?EI=Od+Tc9;#5,_<.TZ(),JWfXUf8
&7V6#W3&[NDHLZ@^7Ac08+Q5@W>^-TAcGd9a04Y(.I@8RCJZ[OD:JNg_3Z@OS/ee
MSfX(/#<.MD2-TBHG;Q,4OaBX139C+1:M^3C8Keb)MDMHW#c2^H[J?87MS7UDIU=
M-dYE7EP=.?.eXJ-S/cd.@gK8[_(X]^-VCa,?L/_M41E8@8M:R/WQL35L7_LQ^=I
e..ggQ11?#@P+[A;KR;UH35_@ZZ/)=.eA9a,=dCCE2+]^=7NAQ)<OI_B@VX90.2.
<WDO(bbI]X6Z2&+^UQ4)+c4Z;cYf7,#C>BFKTT,?_06Ycbg^EDP_GC2TTY)^8]d]
)Ld4Ye;B88=PN=^^>EGDER+9HfIRKbCYg2<fIcA5NM?R;;V^:+=S_aR]#fAKPDE#
<YeAAa67>B]<1:=:7J/(-&?^<U2=a&1KF6LVVBT[D3J79.c6RJD&7Y=LXHY<:(K^
VI6=Z2_=HRLIPR;bB.D+Z[F)Yg338Gf;^?_)Q=:4@]+9DY2XOd\feDUUe50W?<HJ
=DL)(7\9M3<]XQS:0;YP847\01G>I>>9+Td;&PCCE^-<88.-2))#eTgf5:#Cb4B6
f]ZFZVTH.WT&Q\JK\^AdEL&AfI?+cTY[f-;A/7PQHPYI7-(dX=I,@2(:#W<-Ne#5
\:#;R<[-b=<RR?aKd#,861WHW_^6KBTc[T9MB4V5F#gRYPcc;0(TQ<#^7PV1S-:M
X/#UfGB/+U5,9:SE-R3&]=P/g#XU?N1U^ef2/X?\S>]\<?bG/E)&/GH9\JR:.HIL
AK?W\(N9?A>SVSe4X1-[7BF=\CDePQ7,LKMN?+D2]BY&Ka(+M.(S/fKZdNbGL;<F
<]T(GaL,#XcN[:WSJCUVA/YdX70VARL#CO\?Z(,.49A,]..+]@.F9Z+2J5@F[adM
eZ3)_.gbE)3.P[;K8L,e;FgBB#G;OT>&_3bQ3Z#GQWc]DI_/9N@]aP:b#XF[)3B]
+)RHF.a[4fEa8)RE0.>:1K\:@#JIU\O1OX+,a_N&=LJ\A(G8JcTb.Ya)>VbLZf7/
6,/Y23<W[=c7/0?>5+FdRd/.W>0I8::08,K6,f(aCEgD\+M.D^LK?DXFNR#ECN\U
C<F:)g[-ZZU6@491\N-_9?^d-J)Wad79Tb@<X2f4C8a&@JZ9B1YCT;2S4CE,ZANP
K8UB7PPaT^/F(BP>)DBO-8@g<L0W,\gF4O3<ENc>7B&+8+67#e7Z(f4/HJPg,#+M
UQI]fGU3R98AJR8N,WgIDJ=<0(:JR@GLf3/?@[gF\UWBEQ8BFMP,)3&]I&DfeD=?
C7ZK\aR^D_^7c;J:U+65_<P7KZ\9-R^#\X/0/-H<S=Z2K[(=^Hg?YBQ;;T=4gb;?
Gb./.02WED5)R:2_C)>N)=)2UDFbZ^f/]6(RZBg#W_WId6SN]27<N(]K9aa_[7O3
LUQ#b8PcY11E1+.H(Q.4(.[I_,UDE,[4DMe&Bd0V)J5+Uf[3;O+:?_QRS]YA+3\X
>E@W)Z\#SK?,;567K+Y]M0-:MTb42J[)aAW7-gb)A]7+?b>(=#;VLQ<?a8R7=NHa
Z9.K-a32-D=A&\JZcX[OS=,\97/H.&^GNQc/d#AAQN).<^KW&O/VO5_^H@^?;Y_:
MWROTMWE&6d8?Q0ONOGVO1PbCb0O(A-Nf51[)8MC5N&3KD4T+eLVcP1][eaHE[0G
A?VV&)O^P@TXf#X\CV)T:ET>ERaZ,JB&aRQ^)QWUfNZ>XI<dZ\W2dW\<<\S6190:
;J[O8G-4U;2^A#a4=T0Y4aHQHB]Y)MR.d+F^P8MgUdDe5QI]5M7)V;C.LDNC;2GG
b>]2c[[;JJ^@5=a_VM/2\0Sc_0\5Z_(I29Pe@G(&LM1U5R+g&MRU.5-,.:Z&(0Y4
]D(Sgf;#P(T;g/9O[AMN7^g,.PZAW19@7H/(HgO@-UaES4Z:4,M^=#06N@+>cBc<
G@O/A,1?>W2&QE/@2=?WO\VFK&JYX8=IOO=c5):^af.L\JVM]YE1?FIgY#AeVTK,
BL9f+7(:4(bMIf#C-20,87QB^G.JbdNHaa-F@Sf5)bAH@5Pc59Gb([AKX8E^VXS7
SCX)=E2ac;_ZTf.Z1eGPZ,ef0V0;./2;e6Obge]bZ9cM19,[[=(#(V^K2YG2:/OT
.EHWg^@?;EB]YQ+&#7><b39IC_Q?;BPMD+V&(aX2cI.?<<NDc#:N51P1WL6#NO>0
e]_8TaXeCa7]U1NME&6EDV9MbRO6cL(_,@ZK/gN;I=G(?XHL=J8eZ:_<;T/,b>5M
?TFP_=&HC+d#[KSV:Z^IaCW)af58]a#5/eWJ=QA<6Q9b,WfURY,WU2^ZVdC>::=M
g1_SeS6E2Gg_99].GX.IEV].+2X&40),P@dRAadD;Y1fO@EOE)^aO)VNUE_gO[J.
>.aOF6Y@#XL4K:JKSXJ3\-&7]?7^6P[K,)TT^IX]F:DcZ8(\VY4C@7_-HV19H:JN
]E/T&cXWR2;H(S0:5PAO]aaA+X^DGOM#5.,^eU<CCd+WW<-Q;VZ\B\992YgG6][a
/[&+\S\JJPS1LP<53d/W<Afgf+S1g\H7EA#dD-V#U]La\?f[J9Y2T->B5,^WJ4+g
23OT4IaO,=DLNAJ)>5ADG<]8CGYc&&UXA;AGT3)YL:cJ0^Z^>aJ^e&f:#)gJ>Z7G
./OfF^I+NO00dX>G<+@NHM,W.-SRO-8XIQOG[@0MR&?->MV4Q.CZSQ:LP0.S7JY)
e\XT&OKG?ePW4A=>6H/+8)<@/?YHe;e88_Z(N_TU7;=CDRd\>>JRXfR,DO7ZTJMg
F09W1-ANR[WU[MPY;fJ;PO(ZbZXeH\4JK=^[Sf(<-XO,b;\)ggMM28X#G87CNW4L
P[>dBcU5]9F9GeUC_AWb)I5JF:M=.Y/f2(92;?aAB&dKA\Z#RO9P#Bb8+)UY>76-
FfI\_Ed5,Ef<>69+OFH#;EG(PSeC_e9_:YH0W]8018T<e(K#@>VLKY]EYbb^_AQZ
5<QcFW1T>_=R4FRO?GR]+PFUUZ<[BdfY4H@eHWIZ4IJ\]8bd0[]7:(2D+X6QgF2]
K-X]@eIQI9/A6^/&/D_bea066KBBZe+(R9)N&92VX/;87(A6T\Ee]+.@B8,?;aVZ
-T_S2IX_(X0F-Lb-6@ae16R5,HI92R,0c/OA#IQ#b?\CD9AJN:^@-GN:0.Y6Oc\;
=K38?VdH(37VX][L.1>CL[aE;)3MJH2a_E/MYEb?]\0;?KM;&H5DW31NN65M&\U)
QP^,dRbUL]aM;cE[,Q>Q[LG8<H8AccHOSM6WGJYHg+8B?EIbVO9dda)gTe?-J0K9
2J)N,(M3ZR7_P2(@C),[LEEZeTESG1KRYfUBGY/[f0>@Cf1>L:ZLL93gF8c[@5R:
W=#(#Z4+H3D>V=:N(2aOJI_F&fJULK5N;B&ZK?:MZHa4QN.R2LQ<KfH7HP5Q9ffO
>3R:,be@Aa.<082(0V262\aaa,E_88Pe_=c_[bN]XDFGeA&.>G=RbD]9PN:Z77@W
TbV(NGd,[,SdTRB&NSR0E1>_9J#A-T[O/^#IC5+Ib+dg+-]b7T(W,29VeZ2FRHMR
D^7=U\MM3]?^9#MSRM:fcJV[gK[c,V7SgQ@^g?[\#R.BHdaL0^9\:YQUWT_-I^C?
ILD@7-L_/N4\S6eG+C_\SXfe#[\@)^/P4IGUK,TKL8_<g2V8^(X81U7^V5215XZ>
dR7YORJAZSUA9)[RWE<0CC@.dNG]0UH)HLVZMXQ@,eGBJ].Y5YT-ZP<DZ<S<KQ)f
>7fgI4C[8Ce=IF72ZGO)QC1R];B4?),WV&P:fL?MU9)P\c#6Z,Q::M<DL$
`endprotected
            
`protected
ZRC3]<=1Y(b^6Y[<fA1>+F5^_-#NA\J4cI0NH;R=.EZMF4)+B:\2/)<dcQU-U(39
LC>Q3<YL(6#>Y=W@J>T)#_f:MO\_J_717\Na/Y15,;+d/6S+)[L^R_3La,.)=:X3
FLPV,<7L/Y2KZ7C^5ZOCf#V63U<[2,P^fU/MaNObEbY_7+MSHT8A-K8,=YL-bF4U
]?e;S1FC/ZA^g1I[+d<:;AC_cZSJK8E\Q\EVKZ(VGRG)28F\0O&=c8(f&BI5RZS_
I[T0UB3=\Z^,X[DD+<O0)gM7MdLe:T9UV/N.-4L4ffILCHdI2OcZ.N=8;a9bK4/;
;6>MA_=)DH(,-$
`endprotected

//vcs_lic_vip_protect
  `protected
?,@F#EXHcV/YL6_C1K;C7I;KH4\0I=2DV:[1_>[;4OdG@bWN,7/4-(a)[MC;RgbN
CRFGRO(M^ZfGI8&2K:L<-S9D#+cVO(?5XQ1O;#5fX[V?;?d]7DNU&\])dK:;S3:6
B_8EcYI3X[fM8/afY7_29>RPCD32AYT.bLHZO\/1aQ0ZAO7I#_=bdNe3M(9f;:e2
/C(RK,d2KS,<&1gSX(+N=<[I0bSN_#A2AZ_IL3E+J9KA2:O6B\_Q&20Cf[YH?#4U
H\ND(V585DRZfC0P_]Y.8?Y0YZ4Qb[X2-\:(<6KKb&T+C\F[JLE/HP(]MMfJe?H/
+cZW+64KX:4GU]&f.GO_L7SOGBVb(([Y(gRMDL0]L_E)cF#WT19?[T.H4;MDV)=;
eOEBTe]TD[Fc@@>#PJ.N_,YeYH2-Fb/RYgAf@NHRUa#>f35c&08-)L4&I0PVa;,2
&92MQ?BX1Q_7DN[GR]Q=?@JbFEP4a64)B4/d_-dO@gZA6(dC)A<IQ_FRZYBA]7fU
&OZY7fNO;bA9aP00<JT6FV+VQ.L0D)TN>3[X.XB=W]Y/WH6QC&5]5+KT:a5(AZY,
7A,f^g98\U7;^PI^G_LCL/bHP(RGTFFPKc.&=<ec9S3#.1B:Y]\W8:=8S\(bO.,b
I_,I424^Mb[f][#_G3;[>]-3RP.@4.N[?[U:I3X^LRBIQ+E=KDHGUWMg^,RDb,_e
6\QfZY,VZ:42.E91+(Z]d4<CFK91?<^78,V=J.8A8\GaD7W5H:VWgW2[WXA7\HDI
IYS#e/bGQRNIUC;6.D4M<T9Q:;HN?&9f.GS?Uc>5,2DV(Q:e:38B+IAIXX9D,1IY
T7gEP^cN11/40.g(/VAB]#C.J+0>K@29Mg;2.C-W0:J6F_=.6RfX9+b#-?+#BgE)
039]LX]_XK#,>6D7Q#&9<+g.\O<KB;&]#U;\U7,UG&TO@,4#XB)IfG6LVF>)MZ3V
CU=,b>/gM];dG((,>.<IKb@W<X6a>0\f&B6?gG38@a1R2RdNd#=dYJb;FCcFJ,8/
6EB_P#4=5[M2.DfXEOY/^N_P<+@1QO[T(TgQ7dMS,XS0:TAVN>W?UT5Me?WC[d@W
1X>QUKb-#C#)]S1b;FgK9=BI_:c@PDV8VF^5ET:_8,GGfK@TAcbN_MU=NPD(Wd4P
0UZKQATD)T\]Y@1UIM_?L2^)62Y.Vf=?_V/UFO^&3aGa)aYeJ0(P<R.@@FUT.D#)
R&]^A[_195@S[GNecD=(\4-&_R83P/<2M^Y:RUVPZ3DW:I7I?KS@W6g_;&WCf+gJ
ZG-&,b>Xd/JZV_a3&/^bH2.#:SS-:Z,W_>8ZU):AT;EEU:DH1LK+K:S>DWRCFK+A
=7P:1]O>3J=b0d/B=\Ra8\\C4>CMKg3/K//]e&c7ZE#&Yd2Mf2[c:Laf-Cf<[]&L
_8GGYc(A?+RL+KY,)]L]^7L-OQ2RLE_PY1?6/.]BJc7Nc<_Q&2L<3=LgG[SW4WNT
O976Ie3Z3g=R8/cE4(B?M/c?#]=HC<7G^^<3KLZTM>RK+K5+Q2^A+HN-=Cd?1OMI
<\R>()/gR5_N1H]SeWMU?HL?_JEWSI.U-;2G-f/gLB9L8DI/3>^/C^(E0T;ON,86
[0_+0W#O:Q\IUdg(V<>6[:caG_#G+\S+#=OQ.0\(;OPL2cXgPe=@TG\H/gf2e]2e
65\7[.bN)W0;=R0g@Sb.S8cRRF[AFC\CIUbRd=--[EEY^62K_^I@05=cdTeb>(MJ
I1#4/C7cf&:ge<QB@K:C.-F6](/;BfPOdFZ<B:R.b#:b#<+3<&OQ#U<#V.M3Hc?]
A>Q?G=f[B0EZA97D[d+/U;2,eKJU]B,[[Le4X&-?#V>fg#16R_LfPOF]JLA[62,-
2DI[f-g#a@R4dXWQ4IO#df6&SQ3dD<bDZRX<5#\)[HI_VQ-KL4F6d[AP(ec^50U9
;<CLNA5UObJ]0WM)4F?gf);@O+3P&Y4+]J&FUZDA,^WR<X0>0I6Y]F9cZ9_C;0X/
UK)<[a1KG5S97a(;&4d<#TCFE.B#E=de:dA0LA=1f2N#JYVR^-GCOE4R(EKcT;)Z
J<cVKFD..M:&<E1Wa(JH7MAa;Md)3BHB.5d9bdB=P^ca/+c#J4_B]edG8XKLWDC.
_KRgI(QEJ]g.bT;++0Lc,BO/_M2YYTGE_4(M912-.9OZ8Ta\c?@1C1ZU>76bD<c_
-F#dQ&fN)e^b:\eQ7U-_@1]2R\3?-5dEV9UXLQCa,9S#.#/PJOaC6caF8?1Uc-A,
7J73O[f0+NWX<.CDD^ZRQ=&c?R>&6g,?IFPX]6Ue@_B0[H+NAcA/>gZF4P6#7=@[
>7H7(,eP4G7(GcYa]a<KQ-7/UW>KNU(EBXN9O1e.EDPJZg[8>C:<[<0LW-DTgH_&
Y:=Y]ge#D4Pb=J^/N>U(D-YfaBQ3Ad-T,_gP:BDJe^,@H\14acJHM_Q4-1DIQff;
.XZbfI>^fSF)V:_J.&3];-Q&.EGL<=2V:EKDKd3R:I2F9Wecc7M&A<06N\6IEPdY
6;X;^FYa3N/1g228V_LE=O6_+.:P<@b?Xd>AN-8^_(-4WXXJ,FB];>eDJ=#OWdbg
0HLNDGJJ.&^/-:WA?B4UEcW)Xc48,_<9_45=ACd<Pb7QQRb>_K]Q6ZY+6W@X@_(Y
BdLObRPdJZKGPgf(<H7>1-a>;.Y.UW51I7bSW#CfX2&B1PgAK8M9MY6:eM>d);Z5
V)dLROH<UNZ&?g;MDXOT:HT]X@\[[af.\A_cW&D4L2(N;UWG6aKaL#8cT)#I@=WQ
M<(DfHG&(/Y<eTd:e@]))&4OXa4HG.JIN<c;ga2eK)da[,\Kg+_dI95DYf-eY4-E
N3&gG,&HCHd5?I8abXf#PcZ:\g/H]N7/OFEONG3)B^M+SP4Xa;IY9&V&&7/LS/3B
<^d7L=e6NYeJc)</C.VJ7:,CIPB\=S@#B/@C^@9F<Ac[]M.GcES7Lc?2S07cRJ89
2VcT8IY,WW0fdd=[<1N@Z11gU5N_[:gXK2C]<E]6.P.1gL[9[FCQ8aX7O63]=T^(
U?-DN66U54B5gK+Z-:@_3(:^?N5[V.[58,@=)(DdCE)K>/P1Ecgb05G(N4Qcb-.=
@#?QGQ((_BC,Q-=fa=g_>N;\S&)CMAY[.^fEPSK3&eF<JEc[W8c2g9=cA1E7.>K6
?;Z@R@UQF)V/L->@]F/^,9^Y#RLY0:^Bcg#\cFKd#EJBL5R9\cRSU/HJ8[VTb0J_
,Dc1(DHfe.15)=(:RMgM.#SAORMG9U=4;94C;X&L.J_D@:7W7:;#79&PR-NU&HYN
=0bN4Obb4b0K15QT)<dFg-.9YBAT\(D3DGEKI<+(=^G]4[?Q3:ZI9.07=#H5P]Z:
+ZY22@-&QG5#14+dC=gOO<1Gf;O\He]\S47C.g#6H1LD@[;T\^T6KM_3bOe7ZE:5
>e?6@]4^^cV4)J+AY.EcRMMUU<D3eUDEaBX#6WI5c=?fFFD2d8;QB>.ZFgfD+?f^
X].[P3V7=P]<F/=gb2#5b89=-FEW2>e0^[a8O:427X.[#Y-NSRT5,2cOQ-e3Cg>R
g#Oe4I6&856FFWD9IcV^YJKR6N>e2A^;/4=RZ7SMB:U/16K.FIG0GFb3M(6WUD6C
cC>IM0N^&33YeIV)3\6dKMF3VVZ\IO(Y+.U6:ZA]YV\K1@]5PeYdEQfG#eD]_?G(
eZT(?AL@JS)[Cd^G0bI2OG?W5UeD,QaMg\LEGY(e++3E0?E,Ga)F0YDN67:_C+e1
5D+9@EPY3_>#TBfQ\;-XJ+ZgY=95SeWPN)V[(#1cCbBd+\]f8.U:J8+f0U8KRE/7
WE,Y)F.g43K842D>,#:LcBB3<2Hd54_a<E93;.FRH^[NUb.RI)G;Q.]V27/Q0._,
?SU]K.3B/.U(;BIRP/Xgb#[NV&?;50fP3Z.QZ54HNIN7CcGO0c,&-JeFW?]<(gJ.
dE#NU^SXD=XZ=aHMQb;ZUcDa7bQTRLgKEW?][e81NC#>UVBKe>dJODBCI:MB:\?\
^Z1O3(@0cBRUK,JQ?c8AIU\^L.GRA1<0N:T>f3\-,@e,eAYBP&8T205TCRUE5bH.
,=8>C\TTRF>dbR7EB:RFK\AUeH1gR\_W2@0VTIM:S[[AZ-b+QM+-6g]FJSDV#cC+
QE5Q)&I9@Q.ZS4GfX5BZ.M8KXEWdE7cYW2M3V[B]2Ee?CF<0FL#)Q\OZF;d66fY=
]U]MXO6eBWB-<E#C80Y[QXeHXP[P18+C6&XBB;a)&Mf-FdUR&USDY/K<=7S<.5P\
IH(\0S--4HfI5_^,[?L0M.#f4e^_(0#aFDK<6)-Zg6-C\A;:X]eb@9QY0JR8#4R;
L6CNe(S&>W]Yf_^@9a.IZ6VPEbfb3MJ:.DF^9^M[c3dBgN0L+/>SW6JP;(WMdR8Z
^(4(g^BNGeWB-GfC]-GXF-J7E1SWfE_We=]Cd3+?AW8/B]9O2WLM^Aeb)Gg4),MQ
YS,4&PCCXN#H38g@/LfJ-P_J4]&d6,06#H?8QcXQ.1]K:\TD^aLbZ]A)<52O=/0W
#,@(F0;7O43T\1^R6]N[e60=JA<SN6..99_,[fc.M+G10<I&#R6V1K/9XBVX23Z+
4_)Z[FV:+].,\E?NP5D@9>H?X11M\6H6H#:-KG2eD0:S8_0]O;V5X@P^9,fd4>+1
6Jg?HCYbXM;b4aM[KN5H0fU_8VN8-N=YDGCcYeX4CU:&7(da65//7b&=gF>.U)OU
+6FFg<g0]R>O@I]CK5#?-MNYPH/8OO0D.bCcKQILAW5-531c0R8S-Bc.SdH1-6/T
S5Rb+);3?&^UY5YAb9fUc>;fFI>6<Ne679_+(_&IG__:BDbE^I58IR&cHT9\IVIZ
8MPF0ISJT]a030##T/]8#/)5((?e2Z>bWQF)#@[)[#9=TS=I+b-&8LOV/-\-=OZ-
=3H>/EX:Q<B&?8DdT.5GWI^\9JGC7Q8)Y0[5<?&8FJM6/ZdBPC9J?;f?gG9>XHEZ
g-QX\;NF[45g:.Eb2/S[@8K-Y;[f(f0Wea:Y91CfQ+AIU\NZN[T+5XdYB;31P4YP
F(fPM&DI2eV&ZCQWU\=YAQAXI-gAb(P?a>b,(IR)]P6AL7PDR;N)=gMW0-Wa6,SE
/)>/WbW#^Z;>LBe^_C>.1;C\IM5@LV.6[M[@F_J?C[eO,=M8YDDRbGR+J,\3Q5aZ
&FWPfNB2.Z2[O]8LNF_@7Q#f=V(HD(b0+ebG/Ne-Hg8:<S>26;O>T3-WJ5FI4(Z1
KF:YW3SgB(\M:KM#a:A82?F(VQ.D[9YbgYgZ>NJH^=5)dRcNZb,HPA\KI6gX+fdU
P<PCM#Y<D:P/McS+bcg:]O>;f,I/-:JIR#b\_#\:/;7(?WI)>0&237d65;WT29)C
]+:[CaE\?U6=[+#J-c]4.KO6(4YC;^X[Kf(gV)PSFB=7.fITEMb)HH-c1_P1^DH,
&M77V(\f_a,JBCA/CTSX)<6<@L9<XPdA+I=K22;7&S&F)aFW&.(\c2QD?Hf;?;J@
,92MaAGfW-aXBDDF>#:GLd(R-:N)2S/aLQ3;/BK\;fZS[PDd/1aOeGKH-]7_A(GY
YKXgH3N9,A>F(PS2dT@TcYBHCB9_E\9CN,]_13C)V]b&;Sa@BM+4E,32G8>-YDH/
+YWIJFD382Va/G.Y^2.cDg?/XF:PM):a(6R\OIfVGe2HSHDcdMOS+FV2JBHLeJN>
7IA,gQ+]0B+I((aVVS7YQ:a#.VR<5FLU5eOf3@6E]bJ]^&(QH@JA^@:H00RYBTF&
Q]WCHb<^TU9X.5+=Y44[J,5_^17HMTZ8IgZ=10_LZ:8;51TUZ(IF<\5MDc;\7_f1
+R\&?DOYV;#[@;5dJ#0&EW:#+Y.R-a>+>R:5C?2De=[5<]E,fRZ10&3=,7MUeJ2#
[RHG>06D)Vf]J0]D-<OcCW/bNSSSOc&I5/,<;P4^a8VF\9ecY)9@S\+2UfE#.>E-
e<Q+2F[YCP<dA@TA4/9K)</eU]5&^-4HaQ,:gVW54G-;G.FHB_Gc1abK:?,RJ7@b
JF0ZJe8J<LZAP)TSD3^bIa&W1DgF93gF=dY-BEHc7PV>F-P_W:#Z-D21.3]8RRWI
c1#^2XLDCU](HPD^?T08_gF1eH)(&g>H@#S<81.b(b-90[A0(7V@2&85XVL.OV=P
Oga.F\T>RZ5Fc87HE384^^?P.f^fd?Z)W4L2cW6=f:IR+EWK/SE/fG;4_\Yf-M>2
FHRS\F[5(9IF]42DCge<GLJSM_MV4,/9]<US.OB92AFH(@?DR9UOP;S;V89[@=&:
ae_&3R.-=.AaZf7&5[AYJK\S2S@cIc+>=&=4;?^VO<JW1)5A:d+P)X:D-bNT(;8d
^N(\6C9CU8QW]QAZ.aIYRF[3TE[3^YLOURb;^S-[G(YD&<RIT.aV9/Bfg]FJ92]A
/V_IPP>#\07SMZ24J6K1XWW_GOU+X3f2DfJK+;O]SQK33?<^OfgF,P#:T/dJ:-89
4RQ9bDO/3BMI>9BLLN]4ef3##K[9)99,YZ^eWX6B6)EbBeE-)7W;8R@LTWQ060PM
4E@6\S(0HQQ-8,,YKc00RSeaO9Ig(0d9\&Q\U3YAffOYgX+f=2F?_=^7U9[[Q+Y1
+J;W5E#G5NE<f:P14O#=Ib[e0LAeMX^_1T90gGW8D(-,T-M)WfHFOP7U1C@9.=JU
>ATLIeK[LLX,\&M=>D.4b3N[S>3)YPG^L6WYV?#fRg/RV63LW(IULb)/VMc:gGJd
AR5-V#Y@/8F3OcGa;(FKFb65S;_G6ADEd3F,UGPMR7Z?[Mb[,YVgRT<=V)I8<+C0
W)V<N)1QHcRV97XO-^K9T-VdXJZ;:3OWKMF0SZ4gZ5BZN5PR4.?[ZY2O=aC0:3IP
<OgL1WEOK,;AH+?0P>FJT1C5.R[Ae^:_F8KPV5CL&/P07aSAaY_&C3]f8ZM5774C
Td]0Zc9(FMe,PGIW#AUD[dTfD7:8fcb://5>+\.aV]aCU^1;WfaWG_OL60OeAFYA
@DM_M5&U61X9A-?&-/U]2E]I6;b9eXT2EHbP6g^N\H=#S&L[7Q>f6WGPYNEDOY^U
6bB,&:K6(F&H4GBCAaT^U9NDX-=BPfb8d+H1)\O@>[T=dG[Pc^R.?(KC6+QXEP?M
PHXI1_[XNE9DGL53;/CS<ICR9ENEa8b6UQ3F#;=O<fN:W8Bd:6faG4eJ<Wb8UY4^
EYNBV\F/AO#c<UdE7WP:U57ae@^9/@G>^48g,=SD;=T,KdQfAR90XW697^>aDMd3
>PDSg[2g_H8:_A0AQM&T95[#T#D3KR5]d2,KOZR>\34[U[7,XQHE#3g3HP)NgI5&
<H]7?=\44Fc4_U-T2@7=FX)@)Z,a#e8:T,[cR[\e?^3@:?8=\F\>,ET0-8JcK])B
]eeG_.8d8&K(F8[cdBV2I7Y8/@#(;0OC&FbN<I,F59-]_PA)=<)^]&A-BdS&A/L2
_\4[(gU,9?BDYcYaAD/8,Q@>1Y_/8Q6SU061bU6E+WS>_ZMcUZUZ-?bAVA1d,56W
5-Q5&6SEdX4d6[^e:J:.C2M[b?C@g9;H]g;FXb:ED3JBQeG/eH3aLbW0RY:BQDAM
44EG7^\LJaB0f8\eOE:FNIKd5P=/4O&aF+;QE9)4BfB^\0X5f)f5]Z5ZEY<e8gD)
=(3OT/&79N,b:b]V>HAKS\]92QG0V&I&JOLbHf][LI<\4TJ+7O;4U3)UGG.UA;[2
,@3FU-PA[5>DMVY5BaF.E_+YJYH./eD=L?@O,\=7(<>F&V?(GEZ?(9I3X63DN9.2
UIPBa/+-a.8S630FRd)Q85,dZ?BfW1:+NSR&e_2Jb#OW.2gR(MR_gWa\aK1e8@,R
U,OA;9#)ZE<(C4+c^Z^;]Y\E]ec3J<[L;_5f=/-3:G.B-N-Y.<e]fU7eXG5E.E]Y
S<O3+?T=/(^_R2AJZ39R5UXTf&]3JD_OM+\)48WZDGQFHDBg]-RT&GC^O0#8OSH7
VBd3CIKSC8/GV9?EcUB-G5:;+&[=@K&&>I?ZJ&Dgd=-F<GCJ10WG4^?X,&G9MgTV
_B,#6(-X^]Z/;^WA)>_/_BWVcM\O<1Y;Z98.B7JH5:SRJ/RQYB]bGLV939gXB5BK
/U.bB,>GB?N2PWe5N8.Lc=+/E=a1VCb8NTag-]IB=HZTBNC@TIH1EeM]#\FORK&<
HfHY7POX<.=_VS=W88O,^A1W3RHLgf<7bN#B,1KJF@N3\bJG/Y[d\#3AA]]#?c.R
:D-_ea;;:?<e<5<U=VMZHdW[g.E)fPT@[G3Xe_df(9.7++Y_O#g+-G9)]248I/&7
T[?I;gU])cRPNIg1NR1Yb6GELe;D;I_,d@SbIDgaD98Aa_CWY)K;2J7E86c>Z>RK
5G]2R8/-ZZHHTOSVSZQS:@YN++F^Q+ZSe-JA,@K>(MaAGg,(QDRU@:V2fPVQ7++C
feU\7IJF/c0f5b_+8Y\#=>]O>WW1T+&,^^)(8O>8B118S2-,C:9A<()<.gE^^]YM
.[TJC2Ged_.KXLW+cYe^045)\#?/R+JaaWb=Q@5A__d-bXGEIC_A1Y\N.H@_B2@a
L8TIXHVXRF-0MLWg022b1+)L5CbS.@+(/^bXeYa1:D;<_=J^/efDaC:d75<9YE:B
X/3>cGNA>;Y3((D?F.MFg4K,9XNAS]OV84??T4fS7fU^1XI=+6[UTX8Dc#2VTfCF
?FG,PeE8[eH],fSG;eDGAYHYXe>8I=->/fOU+2JT8X_FNObWVeS,RWd&0AL7;aC&
7(a5+fbUQ4F.e_<aE^^??8(_S2d/fVH8T85LA^_[LZ1(;c=fWD=(CM+BO/[1(K5U
D[7/1/>>EfU.=_#LL[@T8#;Ae(YX\=+<&V7.,[Q9^H6GQJZ#.EYB[W/=[5YeBa0W
.6PADa4(CR9b3c^,f)aH[,dQ\(.b-675@1&ceMG;ZeM9#cK;^AJ:L=Ob42X2f7.V
_J>F2\>cBHDRUg^0:\OR[YAc[4@Q4)#LfaPCf\2HX.AU:Q5:Ee68=GK/Aea+N#DC
g_c9QO(C\RNVQ6?1-PYT+IbcbRgP>Y2O@1WZJE66&2^62O5]QP8cXE-QL7R9PY)[
FOfM1K.DfODC?/LKBFf87\2)0Z;9U/W11QT.#@gJYZG]\8:CA1AE:18-BP1:OGa?
G.H8&?AM2_H7<8_G2Kb&Fg1BZYX^M0^cKb)95[.XdAJg.d.O>(+2QUCR+ddU]<g5
cZ6/Eb@eMc5.T_N-S7;#O@,HK)^7I-e(WM4MK4B)GXa_XE,gY_0-A+VTIf>C8UC3
A::\<@gFgB^C^;]IA0cAg/DbbK68U4<fa>HWI6#\PSY/<^VCE8L:D\>ce4JcZa+Q
0;c4/DTHB3((L?.DX[VB&C0:Q5KBOFGQUKD.[=g487N0EL6&M690@bJ8&/[acA5A
Q+WJG8V7_6MK@8faVQ&f(;Ff=Uf[J,L\Q)@9SP(X[ZOYA32aNQL]f-N.=5T6fY/<
VUPB;?[VF5g?N_5c1C6QUdSE&]QFCJ:6LTN9-:1[8^S@c5fN#0-)4L34S-&URb-]
d^N_=>,?H7Gg-PE3LAXOa-&JF)S;0-Z/MAZ6>a2>B<&)D@#5&e,70]eM/C<L6FJW
_a^d-]F+9:MH=&2?HQ+L^M/C_HXREe2]aR=PDX2#))O;PS5JY]9ZS+D-HDZN,N([
B8O.,d9c7O=1MHR\&/Cf\aHgL#\fT0ICf2d,3R-I/&QIB]=e;3XI>2LDaP&LS.=\
a/SB7SdfFc2D05gA5_XB);37@RJfb?#53_<#17ZUe)bRB[BWI@](3+.cZVLa>U_>
-N=M=X8&gA_GU3GR)cI8dG6[gE>0OOP680W)8CF=+AY-?#+_::LV./3UM&/@+&#3
b<RHFB=Y.#DAeQ83BQH9;P=5-.2(RA#Q]&[03g2)U&cS>3;.;\2&>GM?#(1GP^G)
&M02EB@9_)9,P71@(81aCMY]:?RG1<:4@-8R2GD90@81O/(EX&/d6W>QffP\ecD\
L9fGUgJ=CYbf0.OJ>_RbaAH5Ha_d2OK??6L+1]66Lec+7GPQ-A/DZf+=F^Y_-T:]
10#&T.Ce>??[M9]CHO(aC_E.6Y.HI=CHZFNgJ[EZ4YEMONg3c+H<G;4@WZ&,G&Y4
1Sb0-V4bT>H22/,=&f@;9c:_X?PUL83:)0&U91bWU/5F:(LX/><NUCT3Z>&V+DWb
\_33BWC-#_C7^T#T5J9TV8ME&A2A@X)f14+dS9Rg[SE/Y@ad#b:5N&ZI<:0SC6:0
5\EMB+c96W34,JTFD\QZEF;&VDc6SEE84HeKBc];+32/fN1+4>9#CZMHFB9]?_3c
1(Q5W//I<;(92RWVQ7)8OdX1^c)J=]E\\=J8D\=H?KIIQ59+^1]dgUY&g:74ZBcV
\H#,DcL6L0,E3VdO5V3RX^B9S<\L9\#IB@;]R#\_e.T)NRd09>E7JgA8TB+D.;+@
6d&2#I2VR5:<WLXLc#68L<;0QNUOW8f@16V4Ba1YV3/c:/=5b:PZ8AXLQ<b^JHC<
Ib-U,Bf5gENRSX1YL,fZ-,SJ5#g0^.1dR3I^S-ULgQL6A+]@a?7R&]BSaM(aI<UY
5_A+9:2e#7Xb>cTQa9Ta=YMYHP3758)7-SQ[VRD<Q]Nf[+8?WPIPE1Q61#I(LJSc
cQ(J5TFBBPEE/K0GHdNfFZ_f:0TNFd@/?=1D-V\HY5:g^a/>d0D#U>2;B)2BE.?_
_J<5_BZe/9SS:4f#5Q_?B\f?g..EDI2PO6([X+Pbd3]]f&7eE(RIT627W[cJRI?a
b&>((4S)b=N->BZ\2KZCac.e_3cK3-UZfS:3b4:EEPY5V=;ICXU=]2aWfTF-/58C
S/FCX->;bLPB>SYI-;>;a.Wa304+0=cQ685/PJVLCI:0+^2+J(WYKGcZJ4X-1Af#
7P,<F^2QKM?Nd8f3BME>]_4E[LeI0BWF@D3[@W\JSc2\b=Y=2R9-X=fE\-\8U@RJ
2PJV=I]19\VWZb4OUE/_4EA/ddJc\[XHf=edM7(,KG6DM,5K@S6,@\3I<4Zb\K2Y
UZRH3<2a+JA2LV=:54dM-FbCOU0.9Q>)#KV<>&(4RZMC/XCK6Rf\?Y,R<WHa/?IR
(O[@/7.I>5C0&gF_#YN<HL@MHHO-OMN^?P(Mb)0c/(4>(+@-Ba@(+[4FA/8T2F(U
>E?3._<TV=S=PQ]e7MEU,5e.S(/=THf:<9;.N.X:,[?VYeBe7H7JCW/LaEcE]Lda
3ScIHGAAJVaXfBN5.7U[JMQ0\Qb+VAbQ&G(S13[<aEK=#WNRRKP3<E,0g[)ZL<7?
dWORIM_W/NDS.cHR54]&RdIYgSE\c/),.)9,P<L(HL)1B=5U._AQ@VK,KPK,g:L2
68C@]/fJU998=EUUPg_VD7G#<2S_I[cMC/RD0=V7,UN7#A<F/bB^.NAD\=?+/XB@
GJ;T3<MB28g((XG,EX6E/-WcW.\1FJXSC&/(_(;(+8.S/)e3O[LfaY=bBN#5DS:;
d/fA/d2=D,:0TQd#1=3NW.Y:&,3&?<=@QG,gM=25)2b#/V_(-]-NNM_A5VH4?85^
=]&XDZLKa7:PH34cG-5fQ7R>^26C-_L1U.gMYRdISeE^GHcdXLZC;5Y)/TA8-7HK
XP@WOe]@0c86X=#AN0NXOH_bWP:2fAH_C&^92\&HTF^UAUc]WVVe,FQ#OZLPP=dL
:&J+Eb)>]9)e;\2G?O,QH4P]QO#6<#LO/<[M5<<AVf;6Y@Lc/&+4]C318f0G3Mda
N86+Y3@XG&4FC[Z@2C5C_T>N1;&8b8CWZ[8a&SVLS-<a0CC5F1/,Be2aG(R4B7_f
33--@JL.XHBI.H/TORS3b,,2ag>F2#<]#OXT-UD5VfIDJ-OO2>3f?TL(KOP0<PG6
L/((KM^#5egT09YRJ<#FS9^+K7.++(R^B:A8.M1WGFaF9L<K)W-+-aPJ1.Y+^.P0
]R->-L67-<]G@6AKf>\g-Ke=d7QYdR?GIV\QYN:OE#:IVMaWZ,UJNX2f9PE(D0:B
Gg9IBGT)T.RQ[b@M,dZ6(c0=IQPaD<S49[8.]9Q^Hf@@BOb5+8a9;F-JJdLS86g.
)QcT0M8CaRH38Z6_<O??,aS_C-@EcX+K<28[^7=9X@Fa8.PNa\9@AAC0.608fA2:
2,VS2:;VID\RXc5edb//.a1XZ+a63:cK;QI6JW@aRa0E+8[5LaXF>V1JHc+_c^;4
@;2C9HWQ]\cKKW]_?=1/HgCaI/06gD^9Fa<M2Gb[-D#EF8-[]6(VbcF]=U6@2Q.(
8^W;V..#H]4,UPI0HSSBLMKC(U\eY7caU,^7#[B7[(Q/a-N@B8<DZ1/R@4)3BQ)7
^K2b1<g-S+;?XKVMVHROJP,Z[?5fUCZ4Sde\S4UJCX2WDc;a8FV2-?5<YE&,RCG:
,W8-+CLQ),DKfaT6Ie_21\0.O/GK]P@\E)A#(57O_7V-U]+@/c30IbgDX-eJU62<
(dZ-XMIYT^6O58O>6OIeeU>A=CM^M&@9?>PM4YJFV^fNU<ZCC/].ee+M42fF3gL-
C@G/(c5M02>6b&5<]/A?).\_NE\E?N9R/^g,9V-g[-(,3La^@aED45=3A))OKQ\\
N:1Q2TI_6L+6Pd,_)^d#GS=KbWNW78M-@Eeg\>@_a\-TG&\H6\>PG?Ie4&T##d97
<&L9S0D0;XCU#5=A1YQWFWT0f17_U7[.^S8E4.M7N0H9.B,BT[eNBP2+?f]SNOR-
I6]<UHK@3MFc1ARET,547[,5LYCDZL84L:YJ;H>KW2c)G-)<80.A8gFaaZ7:B@LA
dHFM31a+YCDJEUAH,<HL@:=G0PF5ZYZe]E6FaRO(FE1,T_U?.Z#YN1<5)UfMW04P
F&eWfaHX;2EK1GfHb+U/5Q7dd^d2.LOTH0PeKOA07_]__G&JQ-.Q1Y)06Q000WUB
9<;PO6K_I\IJOF^EB<SSK-GfaDQ3+=f_?))E)<5PD=3?XBZ9#HB,#2M]^D[30?(>
9(-e7DL9_]_Id_6YY-1S+[a5O>]G<\=GUPL(@BbNfSP1TBbK=^I+(@Y9.9B59O=T
7d&B@U20#CFJZ:J6#+]@4A#WW,WNW<?8AEQ\@KfT/@PD,GBUI/N6Od-(8:T))X1d
<.H]7<Y??@@VF,cH]F:/SBMD[0=[8fA[W?^RKP6910BYM+a[FUMIGESf>(+Fb:(1
AK_M-ZF\H))BJ0><>;E:C\;UMW]7().Ue@8eb5+^FWMR&BUbJ;LdT?Xf-.ePObRb
HbE6D(XgSKOe4)d6g/9,[S4X+7?3GR5[,dceC\g).WQYHQ<3VEQSE=_9E<LX0PeZ
f6<EbC^1F8H]?Cg]5(G2]/DYHX)8VQ803g2:3KfM[=bQWG/+SXA=4:3_YH=B?(f[
+\,:^\D&=Y1^\C59KJJOgTM2+dIg:Ng(fVeQU7KU3G>ZVPPQ@Va9<f.RKP-FBfRa
RXPEE065IV:^?V\@0QW&NP2&UP7_)CV\#;ecI(8ED\3(.]]#]B[G+/]X2(5R@Md\
26>#;L9PPF@BX\8#[/WK-X)^1/W7;OdX(::.)HN8F/:R?OF9bX&Q6X^GFf)R<_/6
CddDYP,e9).<VF5&VUK]R0X8?JJF)_/KB1YP&EVE9:=OU@UG<R=((BX4)QTQC>&6
6YP8O1RR[0&HC@f.J47B9WScIIf84a=:cd(H)EC[=92.;g;+RgW79+[XVW/ZdNVe
^S7b^WKaUQ@@@R+,Q/?7d[K4QEK1U8N,DI2HA5g11A+A_K_(ZN0B^(&KMJ#?G6,E
b9.Y4^V(G6EcEF&)AgS7+O-HD5H3GD+f#.?^&Pd=9^V_)GWJc3:Z@90cBC:I-W96
R9@3-a_\:1I#5D<?M]ge\HBQ3D]K+)=eT45>U6<dDV+]4B88fA><_G(ZR#NW+2^R
Xe&)g&)@4X2gW]O.WV-G8dLK[c7&\4Gd;eB&I9?@BJ0^+[9BV+fFZ\4e7Y0/NP_J
]-G+SD^J+KG4@(04ILUWJ^?Ic/M#Vc?RQN;9XQXXQRg&N,J:#8KWAbdF]41eOIbA
]+bZ(?,3Q4;J;g^PGaIP<@XQZ9MK2@45b-bIL?0L\e>8&2Dd<<eJH4[Y279/XHg;
GOZe9[\W?58<MDO6Ic])eMBP29,Y(cgdIBff7WXE\U@1MNYZPOY\IE1cYJ34JFK;
PN@&+\R-57O)ZKXJ_ZaO?Uf&E#e?QAbBcEJF(^3\WS?X[<:[Z.TdTWNLeQM)bT_W
<A(\_:H_&(>/S7;Nf6c:1JR7b^-(eWf)dHfFL(.=GO/;[UD,25Y9J:Ne>1ae#K0;
(VXJ5Ha)[^B9HDSaI=QacZ)VZ.5V2^.=f\T2;U@bIQ]Hgf)gD<Me1&Va-N\JI;:E
DJ4/47\H1--K7^b1NS.FM-/JbCcacTY>V-?G^5\ef0ED3OWFRUbPX7-U@-5N0=\0
b/A\GUK_ad1VQ7ZJQYf;SVG?NC#H#(,#I_Tf,2<DPM+a\BC3L:=fWV_,7),QQAK-
+EU\MP_\U\+-5.,9a@L_>:D=0dc6TOdZIA.04RV:J=HeC&(Bb/a83O0KGOAb@8GE
,K.55K[I?Y;P.D+UQ]C&^_Q/O0I[;S<:1]gG=>U#e1+U>P9C<6.^(DHB/g:BRI(+
?D:c\7Q=VDJL86A.cVc#UgMP)dPTO>/ATb5\Kf<;1OT\>aE6+3Pa4]D]gNU?RC=]
)1b?H)@bFb@YX5.,[\^B/V.OHW]O\UAG-KZZEO\(&LRYa;(L_<E(f;P9V(d0(^;S
O[Je<JEMWd0MVV2IJKH24#7c8?D;YN4Eb8b?RK,MZ/_\-IBGPNVW<U(F3>U@]&(P
,gfWDcPQZ?8ZPF,#:>#>1GQ]0TV.FJ^^5&2MU90d9PV_GBG/2)@5G+[NIc0_GaB)
VN4Jd4YV#>&aMdgC]\M2]CaH,NI#F<Y#_.WZ9KCL#H.PMR9+XUN7VK2cYFEK>g61
OGRWOe@IWN0?708-S19?&;==8T25NP&&?G1>fe:BW\)c2@1BWZ=QX8U,M\<DI8NB
WDfH3XMTP)1J^dNeMZAWXf_WREe6>AS3TC[/]<PV#5,CT9V^4g0a\3)P5-U>MWW9
;#aa]8@b;SMDD5>,5B?8HS0NAU8[,E@_;?0U5@Y3UJ]AO>b1OBFC3EPN_8U.]7GQ
^^Kb3HfPSB_#cIKg083&)g5XBc\gC9[5I/[MVD&EbaQcFbIaS0T?F5S(9V#B/C-_
V7A5Y62(cH-?Pef868@bd\JOVB1Y&:^CO(6-ZRE0[:]6AQL1gaZ#5YG<gA4\cCV[
F(/DSg47)Igg+.=B=>AC,Ke52T_3WO?)S?N9^C93A@Cc_VIE=f=TKUbgfGe:0?U@
:2]AB.-GR64[D&9+@/U8d-0),ON=DPb<#GI+;]9^?]&C8c:c\;^,N:QeY>]dfe+&
EAc2ZNQI1QdgJ9d_6aa9>Q7@PK2^g;D[e7Qa0-A^V;aa[>O55:gRC?7@f0M]]EW8
/.(R4-.GDOY<0VD+(0OB1EO1IM#E91\e41@X-B^_/0J=H/&PNSMIWQ7K3dJT>HP,
_K+,;K:&gDF+ILcWaBJdFD<E]:9[T1af#HZfGfCLT@,6gZ<93JC+3PL[>&C])GUR
\[Y1U9_9YJF5;14#AP]&8(N)+Le0N8da&@^H>121GR57)MY1U6a7U,UgS9EC-f8S
dC\QO3I,9^YJ#>RaV;T[Jg@BG5_HRaf?W^XN]-b+W6ePC]W<\HL7MA?1W7.Pe;?0
Gb:.^B:V=9_[-SDQ7#VG2Ne3>1fb7d4=43NHPU[]2>AOa=AQ(6;35NWCU\Qb@C40
=cAafQ=V]PdcH2f9ag<&,Yg7FeCBc&R\9B;-NLL.EQXd&#_aU2Jd#8(5d&<DXaCC
-K1H38bdHY>a.eCB:B9NYOI^a>^^4P-AdU2KQ[HLc[0:]NP,HI?_AQSXg_O@B.e<
>NK,B4Y44T=->T3<\TY;SBdfg<-;f7;EbKEY]Yg&=\B).)[^M,4DI&9MI],Yc7(Q
-W@4/7#J@(:85,CPK(aC8SF+RDB>X4IdO@Q9@,H_5#WcCc(MGII]ZN1I>O?NFD@[
5-TcK8+Z8Ka:J9\fc;;/O-\T9UF_7V15f\=FT4XUO3PBA@)>)g,NEXe1WVQKXY8(
?dVW9<MD=E0a[F1X9N_U2c:(,&>D_9SA_cT#91V-E,QX7^&B3Q2/LHgDC=&^BM-H
3eUdcZT_F?=F6]=VZ;a(>I5C059c4b_(I-a9)215R:d-FCcf?dYDN)eVJ2FGIUB8
>f;dMXIbS5^Cf_b@V3@b^G3Y=9gLU3FI7;f<UH6#XWc?[I+E.a/L#-Va2N0<bEC@
SgYRbNd#+=;K:C>PHP7Z2L8((-HZ3c3:KP+Z\eREc.Jg+F,e@[KbV1[d@J4JR1?g
N9/N#:]WQc51\?Wb+^NT2?DQ;LI#WLOcg.G[e6gPZKb@UbF7<<5+YR=e=F>M(X0O
8B^g:>gSQWB@Y\C+]FCD#MNX?U1M>ZPQ9A#Q7R[a^,Z#(IYc-<.TU\[Vf:.H(\J]
.NGO\8cDAJ6Wg.UN72b<4#K>>4V>I5>URc&d7KE:FS8YQW0-_6OOW:BcbP-T:Ua/
KIDLe8\f1SeLCX,N(C?@3UML+@YKV:]NC6PHCEG=^X;a>P+#22_&<Q192P?ANC7J
CEZg7/gDMLB:d(K/gH]f8Y1[T\f9^0-A@\&>M_40G:gF/F4B>L#F)@,+4>&Y=3XN
f.Yf[46D3CG];(.EZ(4aO8f(WKg8d+SBI::a_+H,>XL\&?c85)I1](cfc]I9,eUT
g]Y4U[Ne9II7OcdCJ6L(X1<9=&AN=bRCSUa+c[>7/YUPEBcT3)<c-=cfN$
`endprotected



`protected
FORCU)[7a,5>M7+1DJPY=.@\ISYF=^c>U^GX21FQ2WKZOTAHN4-6-)gaU2IJPbNa
2c7,>OdOdd4-,b],3aBf=D@\2$
`endprotected

//vcs_lic_vip_protect
  `protected
&8BeQ\d=7G_&C9,H8b[J#Rb43]Md=SOc_LXC#-R)>fZ0c1_gE=J?&(>?cS8145a,
Gf_VQgE0g[I?UdRQa+3G1<WS;ETY7-f5c5e+\4Y_>cBG[f,Ma7N17b.3XOPYaV^1
]Yd7I=)455[WDGeIB65/LM]&RM8VI]:BL7eL,ZW2ab<U-BG_K&Z>Z9J-KgIZ\AbU
efV.I32(WFQ:^WTZf_C5S+dCY?2W4>H5(R3N--Z#d1fD4Ag7QIXRKAG<4aPdGBTR
OF^_;LP2f6K:-(,feUL]-0PBTM+3+XIfYLO\^U^4BL+QU+/8G#=V-g:RaJ5P:BM=
ZU5>9K]?@G/7&G_..g&;.81K_KdgJ<(1WJ9_=C<(d@/(@EU@@]6YWS\N6LUC(8A^
J&34GU#,(LaKK,8O.CETWDG^O#)8QJ?T\E@-K.Z9D8\;4G-ZVP8N,C15_F^U(K_5
;M:Z4#327-;09Be3A<N+f8Q=2R(4+([C+A\8DB.(G)PC;dL@M5I6>H\d<2,dbKW5
UG(DaZb:f(_R47MH=[B8ILRTc9RD;55AI:T0:-de:X>Y;)^?<XEA9<C[G6CTG,d-
5SI#4D1;VO)/2cXOM8J&5f5VP6cM;V2.V\:3V#-B:ORf:cPSIMM4&EBA?<._<6P;
L8R&]a<IZAQeWC5e_H;<\.?>R6(=/F@+C;?_6K+\HbBR4)/9T.[;Y,7I1[3^J0[,
E8K^X6\-+QF0]adW?)1=<(4^6.OH,egJKb+O,\:3Ad;4dE^BGY&Cd(9R?\f5KHbN
dCf]JXG956ZL:g<[V)5SSL5,1KY-04::<Y^6Y3KE5;cGaHd219W1__(-4APc+Hae
9;gZ+E)a&X5CK.X>fYD/b;bQ:9DZ#7#;9EK]1;[a#B5HO?[#5gdNTfDd:b@</\7W
(/GDD^\,\&Ja>-e:b.b&.VSWX-L<\V^J?(g:/YSJ6d]<UDY&2U\A\I?0(c?=&=d+
:Xb&Y\(c_g0Q.Y,9]c:gZ=9c=M(Mc?G>SgB.F?L+e>[XZ2)b924]=)>IT,(EV@g[
?29ca@KM8--GK:MT<^]W;P-AegMY:c/+T7G.VB>Hg(4a_MSQXJ]XKCLI18N/0b+d
#0bM&18(S8,)<NQb>=Bb^FMZ8gACfYWIa0-920MSA(4N=L0fLIAaM&C2D67Y]JQ]
+=/cAcW:XI2RS+dGNL1UXFc\Pf_BVS?<PbO@^YGJIL20@@,P7IYL:+U.1V7G^J+E
K<Q(YH>LFXC5:_IaGR^5O^^4/<a/d7FD,bVXKC83^S+BP7?7^-cPPSd,Y33MWKOZ
Paa(8O??#?;e?-;K@gO@F_,0[HXUR6)+A8H#I&;I)E6\D7&9Z^TUUE,=5P5D;AU:
(Ec.&&^5PGPZ=TE>ZB>f9>^I^K0>[EIM?;/W>/=TS+gZc_1S@)XL&P3F[#UDX&\+
a9Q&U=+V=ABQB\(D>8SU1-Nf7N3g/g/R[G,Y(09.c-V:=H>/>SB<Ea=PdLN>@ED]
?>,_(,;]QWL+(]_@3C)QM-71OJ=P_9(9Q@[cLES^2;&4/[=CP1GZ(_fG@YHgLgN\
RZgTe^/T=/1P&,1)+.P7IO\fB0L<cbMFFY,UYO7O2>)>J4P5_Y1]81b7@aFI8b=b
1MU^Ea8d<Y9H_>L(G+A79ZW(4;^5<R3KM33eDgab?09bN8C^Y:Z7Q:/9]1T]P#C_
@]1C,4,P(7F2WQDF9U;)MA>@7UAGUegc9M&J[e3<..YPL0WY.?X[\-V2W8N(fGK7
XD8H6A7)f(B1TeGOA(P)\;>I8I27DI6G/O<&6CbZU0,<Pg2,cHcYg.-]#d#-\FHC
JACG.H,(f(G,AJD\TVb[c)2XbXC&V93:WBC398eI;^I>IO#RgERB:<?:MTeEAFM.
OL^Z/cA=QZ3;^_a/(]5dgO^[)gaa;1WC/^U@?g#Y=[Ee?;8bOaUKE,H3D:0KL,7c
XEPICFf4FSPa\S:@,3Qd?b(\S3\-O2=Lb/2&I6JRYHH(4(.XIS@A:];3+?&EX_HO
=YN.91g9PQ[/WaIP\EQdN<7KXN&g_H_aQcOENM8B>LNHU?3;-A<f0cT.3<e,HZ#P
BWK4;I]fY3?=6@@gN]OXQE785_T4H5.c/HL^1_JgJL<e_I[Y(J<18d]]:d6YO7A4
]6^TV>OP[ZD&ZW\8RI&?-a)BJ=E7O0#>13@Y6QWb3/LcfLI:AP<YKWF9>#)N)1RM
7eJ/O,CQ\@^VN;+[>:H2RVN/9EKcMSMf7^EGc\LZF0<_SM983c[g=TY,_#Bb)UMD
fVOM&F(02IbJMF<e\b:LWAQYZde?G/:H<SGN-#\,c(5ab)gaW#FXFHFgCL9U/T>D
4a<13Pe3UNe/BYNQ;fSbO-[X2=N5OZF3OfK2]3;:f>SYM#RD,5M-(4fPKaSVASE7
GV6>1Ud[c<RTRJ-f;]\KZH0c@?S3T+H[?B(YBf9d+a85A,R_LeJ3@B4OX#Bc8=,H
#^7U6&_9C7Uc_0REAaTR#c8a/++K/]M86C0gD>ENLfL(N945Y3_X&=-S9PYMHEHX
Jd\+)_MY&B3=O,@gIg\MT5T;KU)QG79,9.]7@&YV_9CQIPH^__^E:4T6>SFYT06P
DG?)A4FU9<:G5QX;^12/]2UJ=.#UUX484+_4gML.91GTJc/P1Ig0\eaCP1?F.A_2
LRX7NcXg:7@O^\/D/A\)ZeC=<Y4;aY2Z#ODHc0K_]M^[g(SF>d\cWL(QRANU[,OZ
G;__e(g^J3UKd4&gP9[WO?JIe(5+e[b&e0)21A6OM[FA>dK1;O2\<G&\6Z:=M<TQ
P7SWb6<R)BBW\O=G34c8W(MOEf4-@@T7M<-@V+WJ5KQ?a387\eK3eI/E#XXWGP_N
NUD?&=)SV,EF:V:I&J#3V&U/R;8T-=?T.@Q+29)aWYBaU<;=a2QX7H9TT@UT>N3C
VJE&N3FHX=@/VN&eNHbWf2[0d6O=RVTF_Q?=XS8WQf#=/PL(gQI,TB>=-K4D;Y;&
dYR9eL&PQgP3;Q^8-M3:T@+FeO-+cB<PZc&OW/>#WTT\JFd@JbD-I#V=S.DKQbS\
?Q=Ud>8>S4gMHEN\74aH7_--WTIO?0TDVJ0+9<Ha:J-SHU[Ca=eFE:gH1FdR=?Ye
M6WUb9/_+>LVHK1G:]4NG5V)FeQX[FcVV&A,:D0cE&TU[@)M2[e_TgHNaEP/,:M9
Y8(Q?EgSd8T.=A?C#S2?R6+-B^,/RfD9S#2GGA^?[G+A,L:5?A]D,L3]RVH,#ePS
;LZ:O#;Zf@8+W#H,8:3FcIX((YDZPMM8>UBP>ZTT1JaF#Z5H=M;VP+,30T96U3+1
5Q3()HD59Wa+NLc.:c(^KO_1aLd&YdcKT>IY]@Y<]_9?UD;@Y-Q+We=/C:/)NgJ=
6L1OQ:eegMdFIe5411d/Mc#^T?G:?PJ##8.10,IC_2d&1Pd41Wd[N[14X4d_L[W5
JAV8S2Af11P.TE,>-gV;X?-Nf3?5D9\&FH(?SA_UB\:>DN5a3#2K.P?,4?FTaD_D
Sf5dA,g:2Y9\.OP/#Q,4g2((KWR#)3eD,:NJ(c?Gg^:##P:P4Db1NWK,^C1FH9(<
UGYaV&SbQ=349f=-IVZZB_Eb.>KeHfGL-8EU?H_ST8_0?N)QJ4>XAY5Te@=<OBOQ
2N9#(08-D1Ec-MAbEU]\HB.;\#T&eX)P(fe1MPO/BIR>87;6UJa?IVc0?8T.#_8,
?8RI=JM:K^YJ\SM@DN5U/B&#_D8ZI0,_0+U=FeLY/-.X,P=Z+cK<JF\cOOP[eIf#
3:dYR(I#3V-N7S6McS(7c8MDE[+=;D-#>MBLeWWeXQWR2e7F-IaDfD,YS>ZCOT.?
1g-ECF^9cX;(L=aI)26TTdf4((8#-#QMRb?K&JUY/&^+[E/:9NN9OB?A]adN8[BT
-<gQ[_cb9B?9@YX.4]Y?GOT5eRL2SRT:Tg2cO]Y<:\g&P==^0C4._W8MKXM84)1#
a4#Y/Pa36VHFIQE>c8J;0NfF8c6XQ^b-))@gDa0gfLS/d2:6+#Z.;=\?)1<#dMYO
GY<3K6<:g\(OK;W4T(X:9_=/2X&C6)37L=A92+@Q=<PT,6[U:\C,9g3U#5M?\6=9
LDY/7S[N_B/a.(-YXDZ=<39dMfI=6L@Qb:@Z=Q3H,?_3F\FEgU^Pc]33Ma]Bg632
&P:VFHX8H&[9JJ/(0&#9]0,^#gDU;Xg8[].b#0[4/2TGcP76SM]4JE;JCeLB23\N
.cW/53]LYcSa[2Ngg9Wb);6Dg.Y?H)F^)69PZJGU\<+OF.NODg0158MV842dV#dE
Z19aK/5:b=&QAB1E5B:Y701bLeRXR@93&RS]0U9A?ITRF-H[PN-JVP2ZT#9MRROa
0=1.]-_H@10PM7PB_LB8K0EZge>S<1^BS[^#+GL4]IIbf:Y1N]A;WM9=>d3C>L18
2E?9e?0eNI-eaX@+aAT&9@4=bJ)d/.6@(V03a(Ue>g2)ebMa]]:^),Q@d,^Q8_&H
Y.PIa=IM-?3W=P6EH:0\;H>2]&RQfR2@g6/T]GZ&MUPD-T9BM=V:ZMNWA[S;-R0:
7MCPVFK7[\ffJeA..XW\LSOPF<]K16JMT0UH#QT1P]0b_MW=A0=))bUD5_4RR=7g
\W]X[U=#=TGGE)bR)^@8F)?K3WG<CKY(>3W^#77A^Tf)cG/17U;_&(:9&J)MP6(F
GS^aa:/<#LM6FVd53\GK7+G+9aY@FLJ;A__JC4A)\P=20CYB7[.<,Je3KXDZR];/
#1<8GYY37,I6#F=dZ\>8_IEQ@L56@(-ad\VcdJ7DaAQ?1&IWS\(F]6ZE)7\.+,8J
70cO)CS]7R[4GD_SF_2C4XX8_TJ3UfB;@)@CKd^V.;/R^9<Q(O\>4+J=+MGccG7F
=g&@_KO\MN@b^5I0A:3GgUN\U0_YG834S#B_B9eU:M(Lb-#B8#3KF,2<b-Q7,1H>
7X0H(KX85;bX;afMXgD^TCN-?8EA?b=NM?ce,Nc:SH[MF]>:5S+J(79fV+D?fTY4
cGK1Y;@#a.G]e@F0d7/.ecaa&bUfZA0Of<L:-Kcg[TE3.9,6W^P:]FX0b8.LC#ZQ
2>gXDg3>.2f/9F=]651?JQB<)#N/?,\d?=0bP:=<Q(1GbTd>E,)/MZ#dW@T#UP5H
UR3RQgV?gKGXMa)D&a=g1P9Z1ZPQRO9I,bH:G>e/+^2DbXIg:NMg/N+436@5&PQX
C@X.(b1UG4gV,3eff3bW63?B]]#38^L@_&I_]cTS1491e]KgH0DF-E9+BAFaVHdb
,Y<6Va<eFT:1_+M4A2W2Z.7AD4O4VHO=_PY.:QYO,GF9(96Kg7H??b]P4V4b7dS5
W(A<9:;@RT)a9=W>J,EMFNHLL=<2WH[\dDY]W,U?dDVI11V?@Q-.:EE/Ob&+JO2c
Sc/2d2.20dC\BNJ.QHd)H/NPYM]/,<Ca;3O,g+7Ff@>A4LE)XGA#_;JPMVV.^bZ&
b8@[6F1VDWa_;0M1O,C6=Q&G:bFEVc?L>JaN30[:9V?NLQA(S]L>.eJ:S+N6>K[K
6Z,THFb.dJ4A&g&+W\DVg(IEJ^S+g-[+OXN&Z]f0(DV\f(G+>=F@,CZR9>d71F5;
9QDI[MKP8\-PT]JF4JSL?+ed1ENAS)#<1^AUO3BZE)+RU6K06d&QcAL;GJ/b;#:#
a@T,eP..f1FRC3eAHI,XEB5=dBX..5J,QR(11&RH7We4c]&/U1&7W)XZ=>5)SI<#
9;C-/./+3:GPaWAEPGSI76:9ST\BQ2)_ITN)aV_1CFGOS?R5\5GQCO??g;U+1JYL
AC=BTU]):@IaPRZ0f8_=\aX]&]#6RHOR]+\OPR8Z=>&PBM=&EW_EdHELV:&@.S\/
SBFJX:G#Fb)a>F6U-4<>76/3Pa(LV3.MaeW@#MO+;STg1@GB?R>7SDV41@Y&Ue^5
1[W1DaOg=c,(G3Z[G1B.EB3K:(G/&f+ATX;N:_P9NM(JTRG[fY6H9=[UI0UP^I\Q
_/3S_V>K#R5d#QOVYYA][-C2O[(X72AHbAfb#XI_-3J/Cg@C=3;Tf&\C[RF,S1\e
=aJ4^].PgV(_:U9-2eT[J0J[^._QVQGa>6,#e56.CTZRZHJC#I3)X.f>Lb-M>F>B
QR[O-9+]CI^cL#+178<TZIRaHJ,=&[&BcXE5=3f8\AdE=^IVQ?Q-K=+,1]AOd305
Z-I+FQW\bN050fJD?N3@bfKd]\M/3:,]?ga-L(JD_E_/e#>e2(c3F.9Ib<0Kb4dT
\F#^bf&Y^]/RS)M.L>C=)eBO)HA#a-#Z>\TK&UY&dAfJ-55)GZ+[cBOU:((C9P)1
G@1)Qc&[TTE>RO-L9>I32gQO0?Od4F&@@D^.-:L^[86O6g^UP_6?B7#e))+39[QZ
HEQ_#0_-E?fZ\<[?@Bf[>,e.[=dJGPB;UJD1O#ba:aa[YI@21cNM9YII8XU9[7+]
R27.#e4#]=O2d:X=E.)7(e0Y-/)[3T?d99DLTT4FRd//,[/I(8S6C&)&G?E5c4PB
61^:J&eL.J(W1+4DbNZ_K;;JB?XJWL/>KH+Z;(L5(,_Y:@/_4<#0]6=&]V3b7=eD
4R,K?RC&ZB@):R53I@ZF\ZcU.(B&=H1]\L.,]>(K>Kg4NT,ZMW@8/aKE_#f.7M[(
dEPJ_K6=KNN0Z[X.?1F2,[>YT[W\E0IY?@3?MEec:P-MbSZdf1&VPY/F560#McaH
\D#dPQICAG+4G/CVN<VKG29N==Z8VJIRUH3](SON#NQ#(L@[UPN[g7(.A94:JL=O
9II8f6Yf#N:#+9TO5,[.5OJRE,EgC7>>^\bMg7474.2=_(8OQX1P<fLKARKfM7-+
E4NLDde)BF?eFM=S>2XH(@L@IK#8J)9a:VR]Zd;g+X&6:e0TP/6@4(T,TN8.:5??
JOaGeST]f06;fZ?&QDRH&@./&]:54TCJ1G8]0I=P_g<EKEb&BXH?GaDg1Nb;2D)M
]J6+1-+U0gAV>>SDea&^-c7U15Cg]]X-1?V<b[]6AM3-Oa6XYb@0X[bV#F;5<eb?
.4VV:RAQ009,6CTVV7^9P1T4U>E5gK6K(9RO9K50(0MSQ-5cZHPN[3B;VKNdBKed
[[N,3d0A7cfI@2&gOF:H7,JLMP+Y0<4]NRG<L,<eRgYLF.c-2(#:Rb/SS_?5))^a
UQP8;?0g[g,LD3JSC@3aGL08HZFFI\>?\H#Z@)c(<_M]H:<SEWe8]1E3)@6@EH#&
.FTNJD];\0ba)a:XfX4]TG341N3=.></NF7#PX]f?:g\+BMB/_c&#L@eWI0KYVcc
a1R\>;[C.&L[3^a0bC:^UOCNP:cQ[V_eb?Z^fWJgUd9ZAX>0a6eB0/0^5Y4./6Ib
c2gB/[X)C\e[<QV[P7/S3<AYe<ceXPH-#/1I@S##AJR7Q(;F8FAedLHG5<EL;-=5
YZPAK^B9Zd)0?afEFcW?>7O=/HB62:eVU>I,ZDFa#:@<\P4&fbMSL?F;)LLVOFI-
]:g3:&U,0cFN0&XQXe9Mc@?IeL3JI]>7@LZGLUCQgdF_I3e=;\;>1&20LY22S)SG
aHId=6?2WW9A:9Z#<NIUYD&)_==^@d^fMPU?)4O>YY_[R2VZ7:M8D=6b8H.1:5M9
IFQE0CfMGPITG&<&/)GdCL(1(Q7)-^8a<9GdLd2&-7dSZ4Uc_SJUCU>8YA\Va+W-
N@(C=^ZK#cZKM;Fac#fTL^^\\-1fTPILV9#2BBZIKH\KF\\F1b@2YT)D:&40)):P
]_;\2gM.[&OOA#X=0501C4)PEb-GL&S(4U<GZ:Kc5-J=XK8O\I#SW[(83:<(5Xf#
SN9YVVaCeL_5Wa[5_WceJDDGOOd1>H^f<VdD7CSRY3+CHWPXB+)VffaeTSbV/N?;
ebK;R8SGVVQXO2bAgD50.F\ZWA,U3>MF?U)aOYF(:?NA+.M>_N&^Y=^Z7>6:b6Ib
VA@X)@\WCRPe:?OP7GM(]?U[.c,-&0bHK[fDOWYgNUO7\+ga<A.02UZgWO\+[ML;
>cUe#)7]R8aS7gXWcWJLP-G?FX/-&E:a]?fgQ.ZG,5a;+-eWPO(=\QFR]+g7ZCQd
g<>@Z3P>+NU<7.ICYbM1VQEC\[bI8N1A3[a5S?&NE914^C:@+eC&]&_M&25<DA<=
U2a3NK#R#Q2VbaTS\EKA+U@[)IQ-A2M-F.@g>B[A_ggA_Q/,[T;0-5(J<>YeY\).
DW(CCXG(93H:BZ&a>E^5)R4@ARd.1\AQ:45L,.ZGZY(T>U:\1[J6_CK^L^L;->eL
PdFd7R>:/./6Y2<_b5D//1O1[D&?PVOQ/V8=Q=C@F6WV?TdBcK^Dc-Rg_c\W/R@,
Z@8OESU+_4?E0\I8/^LYWRP5Jg4G5eBJB265f9R5WB1)e^\=2c_(XK9O]V+G97b3
)\AXPfa4+Z]VM,?Ce_C9<1JE]AfWN5NZ,=GN(c&DDc?8dWf;T)YY=)I?0&N@P(fH
#J&>JIG?Te]6[dcA/;Z+]?V25Ce:O&B[R0B@/d?PeUeZUHF<(R)C.><XU^.T@a3J
:O8\9\V/f[1P+M.8&/D1X7)1FX2N?[7gGecKK,FJP(V,G0>cgc0Z\>):gD3UD7T4
P8?;H?I+H][d+RO\P=Dg@;:V@+<X5-_9E,,Kd&U7LV5MLXF)Z7\G5LH=I;KP&eQB
#IZOadYYP\]^0d-4dJ_0Y#N[.YBEV)#N2VV46WOS]LT\G565Z^b;:@TA&\f^N[Zg
G-)73#aEC_XMF^8b(=-YZ&MA0YUR8=71:>dcPU5UFgdK^>+a3&?J6E<;6I>,GGJL
)Z:#1dPQUX#[H43N,Q(<6=\+:UX.A:#T?Ed)L7?:cM#S0e^D]H9eK/J2^@c5(4]>
gfJ##[PXY+3OO\9<c=,F/^>Q\B3L#182aR&f9>\EcbGCS\Fa,CYNH)Vg.UeC8V4F
J,A;c<aCV.RD20W+MR0T3d)Gc#:3G9LKKf4@gGM#U#S3U122Z5=ge2>g[8f]@OZe
e;2OH6#b?G2O+XP8;Ce;>89X-RaURI]A12FB3gMc1^F@U1O,4074@/G9VT4e@75Q
Xd^,XbGIR_BZ^FL@0TX,<[f+dU4>ac><g(C?bKX\d+eN&;V;Q_ID_TQ4_c;14XL0
cQ0&=D?0e1,:?S<1SE[C2?TWRY[)HcObVAbd6H?<77?f+O-aV4C9W5G27LTE<FJE
J-gffe1[O>U3)#aZ^ed^9GbGN?KgHJf(RV6_;EddNg;7S:.(:TX8c_5C(]VSCL[R
gYg6>N/e]O,M@FSDP#><\0#.Y8d_Q4XgPbC79OPUE<IL&54dF;#FCBeMfCTY^342
Kd#F3A_QU#=E1+ESS^<.BRaT[_OSfV8c=N(?)Q<@S.gNKM+[)[_L#Y#MDB^?0(5G
T]2,M0,g8KF?U:Y/TQ/A7A.]&FT-L8J3]5?>6g\B=,_Y(.32G2;>bRR-/>fbg2C3
g[5WMb@e(1#3cSeB6e+PGMV&QDF)XSDVe7,D/O1>>-R+75LTKJU&#VCMWBXNAKI;
g6=L/)2492<&PbK-Jd]L[Kb,g^BT6DM0V/=dfK7_+BY;Aff\H]Y4X1:;eS-b2G@O
ZUTXgWT,916^[V<_c+W\(/L;M;GSOJLBLY/D@:>ZG>g8ME:?ee;PF^aC&V5A)0EA
1[_c7REN,,#Ub;4be0MT:2-\P+PBKHS@5f4Z4BcEI#\8R1&063^8\Gd#KVS8.V=U
7UA64a).d?#QI]YYN,:I7/8L-e(YT2-\S]JEK(K[64;94MSP9?6g;\^KWCH;e6fH
4FXAAXTCTWT&KL_P2=aec8Rc>=d8Cc+C\:>gQ_.;+>;bQQOK>Kc<4eA)Qd[>G2F>
^=:S&E@P7Pb.6IbBc06AQZ:V>&K[Q1&ZAA^A09M8T96-ZIV_E>AAJQ]?6Tb[57Qe
(G7._E+GRD9+H^;51/^/T\WFV43+A@MXME,1[#f(fKO;eS=a4CKbAWC7;0T/TZc[
g&3A0ZOX?C2>GY1UK^&[8UWDfG2_-<&+)0=0>C^^gJ7/<GF<S\:QeWHS]a>a11B.
/C)29AUUDV@9K0+8gAAd7eS<4BBAUeKN8H4JNUG)HE5&Z:[J>JIa-1fBWY9YGc9P
M3&P/,DcKQI8J//W877E,g=#bB(XaMV2CJ2FL4<P>R1;4.(41c/gH4[>-E;TNK7:
8X4-2S]G^U@JdB>0J#WK;56J_9)LH=5V99,bBKD4_XLT4&]:K)_HTU&b@.SF(_)H
d_63M^c=_?1fBHEF6(YOR#6EBOU+;1-#,9[+Ce@]#,Ob0KgO.GQ8&e2Z:ARH^J8d
B]6(;GFEH430NKQYRUO=&FQ8(D=84MIZZ+0FT];U8XAT/g<:>&5>=d/c:Q0[WM2>
^=\H_&f]-SDJ6J9+;F->YR,EZ1E2>JFR,c43gMTK3Z21G/I(g91@^UNHTM@<]<F/
MU3V-(YI>WKOdEc2E<2R(a?C[>#.[XS,KJ:fCIK/AR_FT8O((G-\IYScg,.]_c__
#-O=<6S_GNOJKMQSLdf_46&&F;c>52FOBeL.6HK[I_R1UTNaOe8922^]bT@>3UEg
E-X0.R,0?T(16eZ0Vb3X775d&?.4eF)CcC_Y)G)NB#Jg=7+]#f_,FCfO7I5;MC65
E33L^XI+a-(-B:-Kf_W\O;,(DWRYY^Kd@=E\LDf_+d#=HQA-T>7d>F1HV0NR<GSV
IX5ZG&)(gER=<[X(\.O(:B?NVgD,NS,Q>NR.6aVbfLJ9BY,JA7BVYY/SS/D\:f\B
@dO4\-1Y5IOOYeb\=168?^A1N8GCGNgCNN81KWZ;GA&ULLAZ7ga3bK&J[49#/IW6
612aeQMb-4)S7J()M]<BP._UHG=D)RdTD8X/A6G0B4Wa]5\d?;5Jg]P<L@:T#)3I
T84>I]),G6A]4:7f&5=A,+(P+#;HE;ca/fb)4VbR?[bg/GL=dI0\)dD(YKZY(;D4
&.-_#S)?RB&AX20^O-44TD\#-K#0&_=17NY)F<1D<Y:9IV?bW)W7:;N#/&UACc3>
JEF/Ke3d;Q2a@2KUg(@]0X39[RXNP0AZA?-J=)[CH>g](KX,R_Vg5,K32).5)M97
bQ&OTYc[;-HX:KN,[Y)K>QB199V(1>/^&_TPH7M,9GIYG?J1R;F[1OZdXUL+4SeN
0,]-)57QA5U9-c,HXMQIRHY0X1J7-J(;XLZJ6@3?LZ)/C+G5I@K_U)IL,,?Ob(V_
<;1UZK4>>>:605NB(fgDJL&=J-ZK(b2^bAegc1S]75WfDAA@f&-_G]GHC^L8REB8
[Q0/EJH6cD)B2[I13LcV)V&P+2b\>E?+52cGO90MR@HHH16W0>I,8bE^ZC-XGdMb
<-=8E=/=FV)/FG>2e8Y3T+\S^G(ISSOP.Ba]C,0I@bb\a;Nd&&V?TO#L[/KG[^de
(^H.cEf_25c_;MRZ_Ec(KB+(265ND=0E56V6cQZgeG-\#(TA9NgQ@P95S2f31MWO
AQ3?8HL5c]\cN63EbS[EcB^7^K_:<X)>_W,WW=dJ\,8]@FII,6NYVL2(6P#R?>QZ
T4\4M?,FME9fIY,8cc^^2:YY\M_V\e.M&)(4fEV]f>0B^/I7AL8bA_KUQAZM9PA]
?c0a325aXR7S3=2f.M:-;)b??LBKK-ZB2.WGKRG^a4VD5cY(f&R6F=ZSRE6BWgOK
25VY92)+1<90>(4DdOXCZ+FV(N4AJWc-5W@6#WUf&Zg-\?cMW6g9Y;c;g=\_O.#E
ESA=&eP\5c3b3bbNQJ09VQ#^8L1d]:#M)IMa(8eXFI;5>[SgVAdEBRVP-(c7f6PM
FB]LS4P[?g=@[<gA1L\0SH2<eVMYG<O;V,8O0B#ZD?d[,[ULN&I+@#Ke<-^GF]_]
NP6)dT<:(R;b2-)-(M#Ig2+_N[#6]2B@ePGMLEDHIB)-Kb(Ib78O6-:4bZ#V[#:O
G8R+(VZ,U<)^:^GB3?JIY^H#aHW(+e@6>da@2MQ>fH\-9\d5g2>d+Y7566/aGKIQ
6]B[fAT8;@QKf2f[JE..]J]<YCVC&FMa0<YCY\;(Rc#Y3QTQ^_0+<B=9?<fF:]K(
^2>8\9RI5fSQFdKR3#(g?<WQa2a=f/LPe?2#36V^,c6^dC(bU:1gA<5:g1SYZ[Q@
C^9K5D3?RAQ,(WA\GR<KQU36HeW)b5Q:a39:1F:1<=,IcT[VDe.aBc;)O_Abb06(
_7:QUY2QK8,AVA[ATfVe=IA.O+4bIBLN2SDC0#90M5.^4CeCE.NEF_+DHEeMd>b1
1LJ1[3WC2g5:V7SbNR>fb00d<W(-@,BTKTQ>@[M21HgK];dA?Z(&MaMRIPZ9I=9T
380/PO_M6+L9J#40J;8_,>/-_+[S780->7Q[RS\Q.a^e^Sb=6aY+2#2#BMDV7V98
7XMgeL2XVL-N&8\L9)6af;GK)Zf?5a^U&/0#E=0U\7TS0G(\3BY05LZ<;+21;2L.
4VD_L<fRg2YAF#@63cVG=J5g1]8[G;E\:DB594BL0FK8agMX@<-SZcT,\&\bHaPS
X9[QZ<\4O;MUf)UURMJS(;baQ[V17Q4_[g3EZ=gBPCH>+:./c(MSECa7HL3O?/)M
X0[YaL8.5;GgJGB)O+Z>^P(50LF8C=TFfSd8ZA;2H/R+,DJKFKH(-/eI)S_QeFS]
.#abG3c,IVI^O>PL>W>B^&F:AS\^?A,=U<b>R3gRfS/AP)0NFQJGM3MQ(bb&4Y.J
R,HCZ>#OBg:+FYMa.>OdE6Bd,6\LH][^b\+RVc\<FdDbYH-d;B-Tb^aY-9:75TS[
&H=?WO.3HWeZ;Z4_Z0CRc\ce[/O560@3+5I6-1J]Y#;/]0=;<:ZDgR&L7?VHAE08
b@MWQ@44Z^@+Y@/e=,P^/ZaIDKB^=84&A12=eWZ.H,2-H,3X@4RH?/Y7eX(GSRG7
R1(bH^64UJ449MW41L?=+E(?_TO4@):JR#326,D9MBSOS3LI/eBWbRG/:,aP,)3(
&C/IfG.(b\Z:U?D7B[6+(U:8^g.AD1--&)WRYT3Eg7NgA#0.)LG70)M6FDJ-.<]O
J?[((C,CW.DOJ>\[M(?W,[2KNM(VIdE\U_H7,.+;(gL_VSPCbIAX0F=(?d6H_DeF
(<d#V-\O4bIU?,DRD7//Z^6VD?LF8@UFONN;B,HBPD/W;W.JaWcWH)\Q3EU7RcU6
A=eTg(:/@/Jg#If/4+,47(8P&NZ-H@eYfXEUE_/J.(dU@.9Rf_L]CJGXW80]GFBR
B47.90QK[_PQIA+?8<)\@HWBE7\[0J&PBTFb>eG(6A\b>R)T+[X6,Mfc7F_8Q\fS
CNXIDcb?0P/P;CgWab_=8UX9:6>aF01;DF.,Y-GK?(TML02W#,S#DaV5)Cd1CWa>
Q2_)(#OIK#a3M614L4N,+UcS_^D(WXBM)-.@@&J0L]B>:ZEgIMNUZdVQfUe@Oe/1
KOZ#1YU=8dABY1XRC?J,I,OQ\_4fD8JL[a)H;_;=6W:81&HeJ-)fJ<AP,BM)2^_]
KKLWY#_YDI^aZ8YfS?f@UA0I2[C&J(84d-(@LE]V#9^3Ya(IJK=GXH\G/CY(6+M4
=g890P6PR&]CT;0831=V_fWQdP/F9@FYZ_>gZCD<d=&Q6g8d==/QX#Y7Ia7WcS+S
a@S3S\1<9fM5E9#02A<.K^EF&RIgI@.&DNS\7KbXMK8cMQfK(Wa.E6L1(]DV+W2-
,9L1^=G5D:.N,0aacI75aUNU@(2963#G8:GWC[T17@3,>UegW/)[QI5?2[bQ;B<=
=&OPPD25eBYe-R,4.+1X&\0_>\5G_>c13YQ<U<,AKAUJ5&_A6g&_D.;[Q:X2DWPP
G-D^^[_2MPS\g6/9M(?bCf2R_;RF)/QC..-\ceS=a&.?dNGaWdZLO<QV#dA,^-cM
G[DU(QSTEE@MHJG[UNMC5d3K,X6Y?FV]IV_#B6+Z5/KYWH.)B,B3=DUGgMcN,ZaA
.Q/a]KMK#(fAB[M/d/aOQC1-2,RcFgLbKYZb^G#eQ0OYO(@P+Pc4G)aR,1+W_270
N,/2#A6dfE,,-M_TIV#(:H0^]aN;X4G.FL<;BabP8[;,7\?+-T26_d\Z[^5PDU5(
(WZBWLQH]UU]UUV@;f2T#JdY6B15?:YO)D]1G&6ge)UP5=Y2F<_Id;W4=I7FKMb8
--3[,N[2CHU4M8AZ@.e>MCV,,2-&W_\@65/M\g+Pc]UTU\&CRX98Ae3P45E]49He
T49]ZS<<X7HL<4=4e+BRJU#3A-#T._\5:I;TQB&.;_>fH_[E_2Y[;fQ?F3_.>&LA
e&;2_1Ha>UYNKP(18^;(PcDKF8\DEb4be:[V>#Ka^K+-)6e28]3[+X:^I;QD.efK
TO2cG0[O8050<?MY\6YS+L7#)W>4].1Z+<LL[T>YI@EA7FO613^//-K]ZG2-9^4=
JPP#?2A@8afKA6#eSJ+a@PK]G49T&gE0=M)QgJc1K8WZ0R(.G1GTC@[e4T1;2;\7
S=W-2MSIL?KK\VcOBcDIb8&RQHeH2;HNPJZ);CNP]<b7=XRGO]K,HP03EOKRXcRg
aRaX=3>OW[G#SXdMW5eLM1:E,=(f;)/.5=@WPRI2+)0]eRBD29gX3T8_]RRDZ_A+
&G3Y[_aA>VZ7G&7NY<M@7V\+c\QM4JYCZ:6L/HRZZO>KB(dDB1.18G-=BLefNVYb
DG<HWDO5@a+cL6/C@?^I5/bN<H(W;cT2A2EY2JQ-eB(Q877(113Ef@T^F(^g-),1
1@A/+TaAE30,A7]a<VcOb=98Gb7V1Hb&L_GU>[@;cYY<9(2DDB,=V.9aCAB:eA/5
DZX71g5>MRHJAL^7GfTQ>/+.K\fL?V441d\CW++U]1eeEEJ8#c(0BJ\(deAH1N>.
bb@T0cLec4?=C54&S-NP2(QGU/3J</HWV7g5ICXICQ]dZOZ<_#X1f@L6(.fJKCD]
O5f(9GGISS1gZ;cZ/>F04MaOMCQ9_.=,45AfI6g[f]Pg3)<@F(6:d]TQ1bAb8EcU
e+.AK9RC1Q7&c3^4GAbXHX/1\S_A<<6<#,C-CA#9>(SG.CLa05VA;:@4/_caGB[a
317QB@TH[Ga#\f]T;DYV><AJONEd965Z>ITP(X9dXGR\V&?#IPGWMG_1Y-S(:&6<
JL@/C(#&:6C,4?\,G@c;32C07>-V>@=Z)-UeY5&aOQ1@CQ&O<B9_8OV#;Xc;+C>_
O]7dfJP/)+/g0V,.LS-C8N6I>g3\RgW)e.YFaH+C,C/N)gF\&W=G>:8#a):8/6@A
Kb5]/+:N[-P83OT>PE7M#dR.RYO[3d:@IL_Baf=TPgXPLc#@P7#O&P5;T4NQcI;b
MW@Q--5O1F3,<T0Kf4AKb0Y_JL>J\fgb0+W<#_]GL:M/J(S]UD)C1=JJ#8MeP;9(
>bF2c&ZFHT=>UFCX;Z:\=LT[0\2.fL+/eREc[C3S_NIX5(I;EcHB]R9O^(L8T6W9
B3HZR/.NdDYgU:AZB3CC7-T-S8DW6/##99SJ@;S>G0+[Ugf)+2.C-,D2W=4Ua/QR
cD>e:#CQA?L^>51I1XWDfF3U19VA::F)P1IM+F2/+-A.QGB(AKZ=@\OO;cb2<5=#
aU#9>eV,)9b.X2REM=QWEc9:0b35JF_X=Z\QcYK:E@5M1.KLeJAYJM=-6b&LH8/K
BY10g)^:KJT+4X]Z^SOf[4&?2H:d3<Vd,/KRcK-^D)RIda1X]1R+RNQ]P>_]e9Lg
2ZQ]W;I:<3ZESY,8RKEL,.9c96G<_4#+Q?U@bf,K.EU(/3f/PO<AL\[J164NZGOL
MWL:;YPS?EE=@.?3NO.+DGF)APaA&<ZdBe],W0#=K#WB12&;IYKT5_7VC#YGeLEM
<&Z2&H6\U22_UD+2?O2>[>^NPB,26YOP\d>P\.K8[F:TfD8P/3IY39A_;4g.>=FG
-1D8J&)6HC]2\/)-__.c@=(IJJ)W+_+aSRW8;Mb>>39SZ<=JB>eR=eLRa/\,)e[7
8>?CR,Wa;7RV.Q2T/^=@;DE@@+]WBfFV=JQDJN4g9PDdWPM+1T/,<#aPJgJ/&ST#
^Te<AJZX&?)<^@&@f\@\@b3,OAIBeQPc\6WB#7BJ3ddV1f@P<PM2:-RI;5(WR,M:
OdE[?RI(5\Q,^G9<ALQ>@J-M14f0U1eT5#/FYbb(OgO#ec/MAHPK05;QN(dX>\0U
HN]P5,=0@Z_.cNgc0Z@A]-KKWeQ;ZY=5dUR5@G>](RW2]B4g)bHWbH@LPX_;a6&U
TX(VN^)85@6)NDOGW>Q+fRW1H>\MJXaBCg:a2I@T.>,8:]H;]P1^E_#,g6b(62A(
Y-SGg1FZQKB3OOQ8/-RP\>[EOcT8_M3]HR&WN>73g>Ie[[[/PNR?<gg(+(O4\Zf^
^0EIJX6>-DV7]RE(T([f^_cQ1;dGecET3EIKM@LZF1E(^+9:+_g+5095@@]SW#G)
fV(E_5#)N7(-&b);K/-1g.3Q_FED3Hcc02D8;@8P2OO-YX<+F01FAdeRHDJgKK9+
3#T&[C=)VNO.&P\g=N^;J4,/S-),\M1QQM&eTE?JNN?+Yg3Y2I+=eR9;;_B445.J
f.=38DZ#W/[Wc>fIUI1Bd1;[:2<@@U3>[eJS9S5H&]H.Q=.Mf\?b6/6>J.[,cg4Q
^f=P,RA?=b6O&e<P..;)ZE0AQE8fQg_RFTQW>MC=&KE6-FegS#7Q\BVa\Se#[_e9
,\f:PC>e/-YC\L_Q?eQRbNN&8V:+=P^E+@d]eQ\VfK>eK:c;QFJ9#^:Y1N8dL1Fg
D7f.df=+;Ic>T-09cR;Ye+OVBGKJ/#4fB:F-J3YUeA,]^0U:+(TGb<g4,V\X>>/a
7cc)G5X(:0:>@)^^&?YHB,DYY0DHA2.KKW(eC/QVH=f34RIKHEW]:VH5^LKGW8[-
VC8&&\gNNFO>.KXN\+)NW?5-]0IE7/eV@/I,c^,Zb^H6]8:X&UeK7Gaef:@&DaYP
,FBA1?BePTYYZT^FF+1I5BPB4QRT]R@e8J#L>[TF/.5:N0JcV/0DBWeCDf2KFMWS
I]PBXM#I;SbU\)O.YKPQBJ1H6JPULEFb,LcOE(,BgR@KM,-_@TWTO9-CBNLd;YcI
P.OJ+UN(20KS2JUaY2<UW_&GTWDb-))A^.@VP;>V)V5eC\ZfQ7LJFK8a@O6b\/6E
)ZaVd6?\90.LF.B6G[HedZ@S]e>b#7[[egFLQHY]W.]7b9@_R:X6;K#DXITONBg.
?M[JT4K/>O(b7[13.3bKQ=7_+=1Y#8JNbJc:+4\_UT(-:9#6L(OF-d<OXd\PARTR
/LM=J8&)O+PYM#@<PJ(5W3KY_?Zb6KYQGf[M^/b[C]X(;-&8(\;R4U,)0a?G9C90
>QY\G0Z+U:ODI#2cNd[6ZLM8VH5EK&R=+LS@A_.+^6L5ZYRd;QS:U=2RAbdEXI2S
;>\HX(5CfcUPbLeIR@?>7U=])^(9Ee:/Y=#VGLQVQeg)gM&UU-D1P<,017KU<-,8
+VRH2A\]J2&OT4F+9C2NNb6eb:3J4&I)Y1W4@>NMU8Y8\BOERP2&\d(#@YGS9e92
,aX\CS]HV7MJE\GC1C-?U#NN2HUfDRHbTPZ5Dg2f@d\\],+4,)T?cHM^R9@Ea2^+
H4_P#3-)=+1Gg)BUbI?3BX43E@C:>@=H:O:/\)I0?EZJK:Jb,;_P#+X3g\U9#R+d
1RW+:e;0-?[fXWD,^gP6A[RY\W16g3W#^JNbL>C1c.TUY+HZ,O80Z9(@/,O:H7Le
JQ4d8ZY0.XQRT-e&8Wf+:^^KVbGa&E5_BV]\G(K?eW]g^F4:b?-[Y(9E07a2)d,&
T:->-Wg6R1F9e(Y3cRD67.?,(1UM:LITCB&&2X7-0Rg.[]./0bW41d;bQ+B[7QGZ
A0/M3M:EZ#bGC=#fLC16eD0gYBJ]P3CA(V]4Q[8V+?Z8TSW^N<H3+5R=@AI27PI_
4b2I@4EbTS]?,519IUY,A1>)-4_@a2.I0;Q:@P@Fb:JWPIaKB<Md69X^<D6SUC##
ga];SW6d/F5-.f4+c3Aa.^-;,RM1DS2DZJDR)D._EU5,<;Yd@<.=feV0>Y=14B4;
BOEC1UEK&4P07QI92NYPF+a;5;WdF(+O,cI:#_>H(7WOI[d;G(FRQ93>N):3[K,a
@WX2K@SQ_8O.G]0/]F9822e-0=ZE<J&)::JY.W+JRM@1(>#N?+H=1#86R=>X:4R=
ND&>V^]#WSD3Z@^6+0JX_ad++Y;g_3R>O(MH&\.@C=+G;U\S@3,beO()UW<b@HW&
^@Z.@^b6H3NJ8&MSd19VP7Z_Q3eOdBM7aK44:e@QVJT3EI(H9[B3EIP=U+SXHB-L
;f@a-N>QYQdE:G-MbKd;D<PEKf#gM9ZCgUXcRTC@&?(0;3;?c6]SU#FgT&Z]8)ZL
94b+S^[aPH2R/SfA&8cgRPKLTH(HN1OH[AL&fgMS5E_R8PW.&&OHfH>#D1E;dXYf
c)B6e9D]Z2DcB>@I<?KE\M/N8=UL.?eBbW#BEO.IQ(1T#9V3Z(4=a=3ef4(R.J;9
C=f1L?b_-0]L.6BJE0+=WBTTJ/cVc5Y1>W;6bH,a=[2Da[#,&D:MH48+-Q2MAZJZ
Wd][eO1cHIg)YK5M6WP-4FCQEN<0QWN>f6,b5[A,6d1?R:HaBc5WSdV)9BJXC[FX
F>CG4=>@Bc4V4N@DAP-JQ\RHDb4S6Z6K+[L&NGAXS;[#_b=7Ma;D[dR;)eY=dQJ^
^DP,c/Qa_:2I060YCFW1O9+B4T=<5^>S-cLAXY4)ZYSQ3?7EK.9>(&O.+9-\RANP
d(?1KR:H<?T(Y#A+Z)cHTYE4J(PHII]:&(eGFB=:+(ecdf.VB[A4WY32SCK7fdaf
O.8P(c8?EQKO7FbGZ?\M2MB,Z/MYN[)3.G@b&PTD@2R0U2G#.\3J5].I0M-b6-Z[
Wc.8Z=FgdI+KYM3U6a+-Q^b=N6:a0a#]6S.@Ze=5;Z(:07JHELKFN7?UY+7/18Aa
8B/GLL2N00ZFG7L-(c2??_[f7,/3N](TE5JT8>d-4>&]6R<X)_9Q.,X]T>K[9KS4
F/X\-cJ\B/G[Bd,127568;&^U<GCgB50gY+&]KA9)[\W4@bNFD3A=0>AO<6f2X0C
.+9O0cFeXQUILJZ#345SXb-O&=UCV(<NCdI\8FgKA#0^#H=L4+3G,CSI.]:B.N[4
:8P];(&YO3)GI?]NM<R.@[K+Q:WP^H3T6c^GCEZ_DBJ^@5agO.W2)QI.P=#g\d);
P]^aefT?EEK[P1UO<&KWPY:3Gd>D&EB#f;3^6G=Y0O2cR[)O3J;S:FC@\UU/2-bM
-=@+J=a4+F<b,Z\Yd.VOGD-GTC]Y.3N.gXOb.4EPRYgfWZd(IR6gHJ)_bN_4)LDe
D>\&f/N/CFf\&\4Ha@aAX43/HO)7H\RWf/^O,cM?_J]5SHIV_&OITVbXJ97R3X_9
Le&AE3Y#eW6_+^6-1.E0BM\.1b[/A\3IOYFVf(+^0E+L#MF+#dTY?5=NgO<I7I(f
/51>M]c08YOg>3=Rc3KeW?0DUd:_BeOUHKG[/N:J&6MI=QgMEFHaMKf+F).LP:0I
AUGAb<IH.P#9a/65fJP::B\,&BIDDZ.Cc1RYZ]EO9F>fN9Q5dMZ,GJAX^H4,&?KZ
H&bFa3.:K#]\[g\.MX,O+H&_2LNVa=ADX;RL-b&AYWE/Q+GJdJOcfD7VgC22Q-W8
c;3E\VD.5B]IdAfS:Ne[2#>E&Y1RQ3bFfS3(4]B@>_^[L.:LYGJa&-.=XWPRTLD(
)39:=Z4bDTH9C.BOM>8)@3e:4G=,+20c/O,CG>c1[-EO&.L4T2EXMFBFS^TOW\c3
_I]c&D5HGGLgN?Dg?+E0;9WUL<^dG_&dWZ^>fY+JIE&J6=;5d^KKA=(H,_T-)d5\
I_/._XHZG_#QdEW_^,_;U8SfTV=;a@KfI3S@G4eVGa@F5R9N[12.NP)GI.2,Q)b;
YP+.B^#B[H/2OL+.CZT8)8,:.+4OY_MV3;I(VU#eWDQ_/V538C0\D1V:GcWP=Kc6
>^WMdI;U(^eaG,f#D3b(6gV]=SS^,^TBRKT+H91GEH1EZ7FS):eTbV3ME[#@L];5
GU+CMOSI&CQD7b<3f_7WB<RA.9601IG<==M^\e^[KLa2:C066QUOfD)@E4Y7:&0Q
>b9d8c9:0RN-Xf0,;#SF<:E>J9]#2@]Q(Oa(KQWLOPce^0.IV@3H6HP:F/Vc^9BW
#e.eGe-S/Tg4(IP0<9fO[S.b^W1TNf5-;W&1@3S9HQ(,;<Z3dZ88CSCH)0c0]WJ3
?B>PYFNc6d0MUdI@29f-ALc^KKBA9M4_/SX4C-1XBcC&_6]@SO#WD>=3N?XeC(AU
I^DDJ<-9&1UN^6\GfX+2?5_E2J10_2R/QY>)W9VHCF:L/.ITGC30-+E@/WfC9>@(
?6[F>HLG_7QfG1\8,?9?TI[S.Me;=H#ASKfePKB-TZH35Y\&HbHg<=>:U]7M^S2+
5A0\gLJ44?&B94E_EGd0Q:ba9G@d_57A9H?#=N5F&04OM63=Ma#6XT;9W-/ee:)2
AA7:VV03FL[dEd[QbKcHOPFVC^18\8/\0UU]#JeHd9g_.71L_()cQE(@T()J45O(
,PF)+=@4bUCIJHFC3QPaC/Gb[3X<,821RL7?<80I>E;.W^c8FCd-B6A_L8?H,&4g
V0W&2LM@@[4abCW@1D=R7<K&6Yf@<:Ncd;O.F&[VR_O.H,.4e@L1)_SB&gQ,T\07
0K9(UJ]17SU/D>_6(72_QRR^J9g;^+:PGTE)Q+JgWS0PKDC4QBA58T=^[;>J;Fd]
dc_[eYMeB>4?)>//7H[-:>Z:SESdPf1=E@DX&O6Pg6YVf1gSV6GTfSFDPcH.2T4J
<([)(W48]4?=g4AW3JgO(\:W=;<YEgNcDLH?eVg1_FD8XFO6#e\)7AE;B+d&SL7G
:gAObdPDN)A&Z^=&3KO&dCF2B^A]-BMO4g<CdMFT?RW3@3UX+Q\_XX9+.Tc;02JG
1W;WWKR2U3Vd,TL_)WX>b(I\S+f5;P+,465O(/.?EYO+:\/^YgM-KB=[Z,\:GbS^
L@Cf4?1d,gaIdHM</H?@]DC7;aYS[:@R/5C#fVNTZcL)-1bF2J,0eQ0,HZ7a=CTO
)5M1?A7:WBd-0^8CN46;?MS:-Vg#1A9+:?J?a,=e<ZGgX,a8Qb/NOJ2P>_<1YA:-
RV<-M?C2S?PVI3RbYa]HW0NI3A)Q5&0?M_DHJ2OX^1B:@BNF6WGK@f5RZTJ,UOQ9
I)_<65;0[@.DC,^4V^INXQPC#;(W:_V:XR-9b#QS29BOBZ.-C:L\8/Db\NNAgEb6
D4>O[GaD_@3LaD=2^LX,7+>N+M9dI@#NCF7DA:[&2MW[THaa@I8XJKZ+LNCQS43[
55UfBYBDHH+R-_-H2dY-^f;d&_^Sc?W72&4?\#C0ZMEQ-1SX1UC37RfJb03IYIg_
3@(,/(C3:,V,=J5NB&IK>(<SVA:,Q9CZMA;abO(/T;fB-/A6CKEMKZJFRCb6R;7V
=_0R4_SVYMR,6_6,R:+-W7H];-WHfE><J:4d4A\7#):NEHLa?fTc8:(_5=RLNe-Y
58Bd3L:MWP;(Y/L/f9aZg164fQPSa)Pdb_+cKB.2\5BR_PX?O^0)aa(W\OG7;&eR
RL+<.89^\#3^^W7(P+#@78D@<5#=;WfP:.JL76a,8UcgeJ2:1#]d^-bd#bdeEdA^
701226:+U?AQXYMH\EWJ.Z9YO0=Z@QVSP6]Z[N9eVeK34K)?EYK@&aHH]LcBI=[(
8cSKB\(1(>=RZGe_DO2A[Z6#aOd7:P0b.WTYSS6HRDC1K?-XHG](.f/]M(SIFD5e
ZR)28&7aH/U<TQT_&7DCIL&2J)T2f3Q7.K;,R2^2NEAYVS+I\7X-\:9LgcZBQIL@
.VK?.H+D?D@^SUG&PB3E9VabNP+6aBEH(GIC6_+6_b1\2<(#.>97LVd^>d]Qf#&-
S5ReGd[,OAJ_QR:^G,G-T-A@]F.@X4G^:aYA7N7SU5S@E9W_eNcO-fb/)S686ME^
4+&ePgGPJN:[S72TXcXQ3D;ECZPYNfFIY&3WE]f95b@63dNdSZDF5cOT:1O:>&,\
D&\cXb/LS-=+MR=ZgSaEfHSe5ZY)cA.-LQG^gG68c#;/Y4ED&YL=&&b<Zb1U2;GB
(,:@[J4eJ_FWc1ecbS]];f#RV#F]aSSI_.[N;0Q#32HA#H,f?4\7,1FaUd\ZLVP6
d[J>OWc=KRXea\RDI@4Y-A8Ie+S]5,B.3>Q<^e,;.aLC291Q2BDaZMXS:41)f>,E
M2Sf)3GMF9QZ^?YcfXXSUC8@BFDSUc3SU)J>D.E4?IR0[3^--gJFN-_JfF<]D2@R
9Z?OaB@W>VeH=E38D-JL#Mg\Rdb/[/J?)dAPW&_4O44NOQ73=5:L;Mf:4fCV-fE@
>abe1ZbF2X_;OY)JP.g7[SXJH@R5g=BF<NeAPgDg3CF8X:URHFTG#@gMBJE#T6Ye
g->[2ZI=+^38L@IP_E@]/2KN_E\U+<NH)X5+TQf2-YJB//dWD.+PR6/4Mc5_SW+]
6d#QgKN57/dg_+^ZgHA_bSZ:WcG0@g@/RDU.XOQ;=E26DdeFM8JORZJX37[^&]3B
PI)0G07T&]HdY/0Ad^gWT,5)@(OPQfY2.D]GW+f</@g^PM@?5J/bGFEK:RZ.+6=<
LW16bTVg].63)_N\Zg9X09\EP48(;K[/PGOf=INN#W3C/#Xb0Mf2DLLaUZDcZ1Vb
1:)0UGZ4GL5-_0JdL+2WT0Y0OfD8Y8CbA=P#Y]]&\JKD^\<?21]&@52NE(T:0(DD
d&A<(+/-AF92]0bd[.CLG:NBd\=Eadc64ZLZ<^<_FLTUOTd8MbI8PME<,Sd)Sg@(
PfLG_76?CGGeJAU^aV0]aM6)VXN+3(OR\M]Gd(?^:&/bBC@b;]>aVP-g^]RLBTK=
>-KA-WE7C.Xb+<d4,S-8APeTK3TD5MVeYgf@bIZ62878]2PJ/.e/./d..S-cK05P
]49\0ZR/8PG;B<P&OM.U#Z[HX^bP718DD8CB023G/V_U3)_D3bH8+5:a]2a=M]DM
dJL\(]F[BF=,SAV+fXe@WW&MK>^P=AC(;@<P4CdT\dFH]e]\7BRCJ5beO[A9MBTD
I5P]\3;;_7cOaJ#8JVYZe1G_?&:fNV72c\ISHHZQgZ;3^Z7<0[]c/K:JH7fFMSQN
G#@F.e4A+aScND@N1WW^64N2Z=\14E]17Q#RR1b[cK6(\3@OZ09cHcF59b@Y/].c
?U:(VSF#g_YaXPXe?a^Y]?X/DD1.MNc1XB\U0P^A)\Q=P3A7K<Y#W):gc&R/5_92
Nf39D\@5e_1:E9?CHg?6:AT@N8VASN5/SfbYV1H#)>(9CQD]dCEb6A.T-WD1?g=/
70=@0A_:.eMFZ22P/;[-OO7D7DRG0gE(@)3\)XaPX)R(-9?XdK]0L_>Q3KGV3B@0
U>G>6W>dJ5MN\SQ4PA,<5AW5+\/dcDJ@,(.EeCOBXfM_9,<)c35]S[#7&DOT8UNW
>?\/\/DOe90UGd[46SYJ59)c.63ZBU&+Te/JV/]RQPHWGXW5W+B#F=FQSWeX+-Nc
PIH>2KA;&gAW&YB]Ke5eM=,JZcXa]Gd[I#STbJQ=deQF(0X(M2\PVPYTD=8Wb[1K
J4bW>Q9C7Ge0-HF;:-X4NYZ]0OG/B^6CaT3>Ag]PW5)a&616N:EaPDF4^P5KgcHg
=D=PU^[#5W_)TX9/0+.<^2]XeXO>[()3J&8:#J.ZZ[77I0a;BCa;5U./-e@9aA2+
c8ab<,/:?KJ(Q(MQ3c^<&7.f):8g6a-N.JO-ge9SAdJTeX2H?FR5,R1;?X+SJDXH
b@_8VO>4IH+UgZ&Mc@YYF79,RRA#Ab+4L@.A4bFU_fK.fK<L_3Z-N:CO0T/X0AZQ
3FgB)[>FNQWd1T-#+N<-f?Wd;KI&QX&<ZI+P^CK?4Y=aWZP7+O-R_2;MCgQ2;.2U
WR70X^2ID>87LaWRCV\1.C7@=#I;Q6H>5eb?E/OG-\;V8JY>]^2<02,EEGJ2GT0Z
.F.4ZALeU@13;J3\JSB&1,BAOI4#16C5_YVH)IYW,C:OBBQ5U[=Q9c>07NQ0<X3F
SAE0--b;@M]H?+eSeY&UTT=HY.+5_GeR/3dMQWQeI?/e-M?K=\,R^;a>517S-S8=
7TdLHJTUg)Q2BIHH5+_KXN3aPfN_LQ^3(cdW=2f\/SAf[7/>+NXU.^,SB4VWXTEI
A]XG_a>\[;3VXT4=C,Ic-PPQ<Y[K]HaXAV_ZP)8P+OWgJ.S[U+WOG/gY.8deR[_N
K8JS/7;EfX8O24X?@B6\U7JQ5#/\;e]a)&\5dTA)Q-OWIU#Eb+VLI_DM)g5.^TA_
2H9I3<I.O,U?cbV&V/)8ZM?2-8W>1<-BdNaLE92613#c#I;>&-\>&bUGEV9V]?-?
g=,Y?^,(RZ&W;Sg7H:.9].T;OgI+82=Q7##H=>dJ96NM.8@6dTBKc3aaC;6.NT<M
KO:3[U]4<XPWGe\DJ.YFFI4C1ZdG^,(I8N1cB)f;@WIaO;WFQg6<Y46GQI6N.?/#
E6:1([\=A@6J<OVI7c=D.RRG47[#(&UR[\QE6NeG:b8XB96(3@WHG>U^BM=I<>\G
-[BZ,SS;OQ8a+7-1;5X5<=SDVZbPUR61.G(Xgb7EYD4b?T:-2S6_O1GgD[c,(:=^
S4YddX[SWMUX4[AUC2Z7?c_7FRFVdHCDBF59#bRZIMV-QRcGB#0Nf5K+0/+-A7>N
Y#ZP(MSOX6I2de:OO]9_#e.6-BcV<</&=8V&D=WXAc]:1g<V<[EFc\W,T=X.O&I:
V-^&:8cPIT]]V/:<:<\He.W)XTL5aZ;X]WIRP7)GPDH;&[2gJVCX4NM3S-_CF3EV
2L:Q?]WfUeUFH_ZF<),/F76Nc3EQ)f\1^I:CE=ZD(KX2/c3FI,e>6.\B[fC]M1\9
E8/,a8H^@LWb+TKQBMg75J5#LF,/&3^fJ0S.E<:(e903,T/4T<JY22K,2T].b+=V
W[Y?(,d:=(5gcg,Pbf.JCUg<E>7F[&E+0T-\eWQAgg^VaeHHYRG?5/A&]LcF=Ag7
[&;W.-IXKSM5-\@O5QS)><-2N>.6GbcY10AfQ8=_d1:E3C0)dM(@7Z?=34YSK;cB
MV/3UJ/D9aW/&,>CTSZe1aX;HeSP)&L.Ncf5K+:)KK,B:K\Z)YQN>beGG:4f8:\6
F,\a?OJXG#YNe8=\[bG:OUW8,3,7WPW5d/9EWQ18B\cEY?D;0?9^>Q=Cd-[ISefC
99_:F4;6/cI)L#7#KJc(W5=>D(^K.4aHDd1R/FGH.5:8IJHXILVC[)_86HR:0C53
]gN5X);H2CPOb@7J8LR?#^b)_AT8U&L-]eL:.f#_MJg,Q()M(QScT?0[>TdId_J,
a&153E?d(G1NSE&a2[]?:Q(Y2_I=TJ..>E6W-X][Nb:Tf4,?MB^X,S>]P1J;QSW.
H_a?<W?Ad4/U.3@#11KNLJ08#c^Z&CRBP<,:eC[Mg@1KIcM?2=V71PE/XV8NZS)E
,Lg?>>E7918G?_9/BeA2YN4WEME90T6c)>X#>b,^0_GPLUbX8Z/bS#WaNV-TOgY?
(L>[Z;JPe/,TDY;0TeD/:O(?Of3\:e\LZCcY4F(]1,/dDb0e?.IG<JKLLED-aP&e
_;\+aEU#gMfDe;/7)9#BJ=)U>O?_RMJTEK:@ZfJSM^-3-IA(?2bGP-7M5.D/R\QK
U+;2/\8B^bT/,ZAY]?e]A/V&+9TN+V&&8.\W)J,fPIc?f@6cN?XRL0A^N.fbcS]a
/&.M]#[6]a98YMJS#GG<K3gaG/dJ?gI,_K^YdZ?U(6a2B:US>R+L\9S;63E;42WO
0II,X(Xg^HS_ASD.7cdLCF:JR@.T8=B.?I;.fgX6b)48+B3_C>O^0VdIU)T\MW(?
#5NEEd??6L\JgEN2-f\48=6O-cVf5?TI3&FW35[=2&+A)I\/\N+^IJ.1&)9H7CZ4
+,D4PE.-LLdE8J/-DWV#g[=)]LJ&,XSORW8)3BHcF0de<DDLBE4J\7&eAg@Ja(79
HF@4YC0&UYK@(<QK>d4f7(G;3;Ed?P5<^_0DdYMUK#Z/D]2E_7V7e->5?3+]Z3CW
T>)V-;,+/?P>OS+g7eOK3eD;]-5->OGRPI0Udc0&9B/P+H0<&6b@K+>.T9E:7Z1g
&e4cSEXOM+5e[4;+?G5HW44KJffH]8-=Va1OESMQ.XIA?EMdGL)@a8OS=51ePc16
Cd+<aH0^e@M=I=)4LNe:X#WC)0>\F,\cW,9OO6\D06Cg#<W)c-VT[>d-_OQNN?]5
2YgNfY9&SWA;V)^&PX8F@]R(?VT[[Z;=e.U-2F^N+_+;9F+__<(Y3]HGCV+YCL?I
Tg#G><fE#fU8FOWUPCPAS-aNWLY\CTc\,NS0[[D2b^=&W]&88:3.cbZ/FRaNVJ1D
Kf]dAC\c0M:]MaHF)F1-/#)4(+)IPI;&=U)CIY+AaB&fL6<+ANMcA06(WX8Y(7d+
[_CEM9]71O.CQ1UBU3aA8B8EgWBIYbU5E)9GZ3L3;Y&#4dFB=a=_X@cBf)NO&f6d
IAW+&YW8J3U9G_E.LBf;HS-+E)^EF8Zf6NFDJU3G9g?Fd_;6@>M4U_a^/=MS[))^
X:U:U+@PXJL^@4]F(8O/6W>RNEe,.S/.O[C<3W.H3SV#>HZV3JO)Z:K&?/IU^a5K
X01N@?>5a(:9N8?gD55R2,0U<^T,/_\@AI3A0H[GA9)Bc0BMYKS2\C>eL#7QHY-X
e)c8>A(.,#9?3Z4O,[Q1C.Q2=(G/JH2KJ=CV9Oa4?<61K]_EAc[f:J,6GN79M:A\
-JB^HG=\:f>HVC-eZGeJJ.VF++1H]2KUd<[gC&[RY(XB?1^6<[P(I.,LcD<8)Jf_
e>MT^RX]+S(DgZ[1>6X68ZdL?B\e&?]NfgP0@/.T7.2^KReOVY1Zg@;=R^Z)+0[c
CcdR#?=]=]dcHH:?gE<67=TMY)_EVc2?g,=dU76\Dce<M,<VL2L4HUL\26)/C@,3
AZP7RZ/cLUAY\VX_7)?YP7Sa/H18baPB;45<#+10Z@/H#OM/_6Y[c6O6DU;&]5gG
#O237>6>;IY8C#5Tf5O(0/,MUUCX,>\&E3f)cN\Nd-N7;5CQX?/8OE&aG(XM2cKX
GfCA]6;ePE4FXe.5UUfP(AQF4F&B3;0]ZN((-)0)P:_aQF.#bSbE3XMg)[dg]\4N
\V3;:b3aN@4J8PZ\_WCC=Vd?=TgHE&JM0<9K6GLHVc#/J?2?#^&&+bCfM\<T/NUG
QUdWMXUBD^U[U\(a6\CIE&@CG38&0BfH?c4]g,c#YWbC-(f?7V-E@QBB&6c4<b@c
DQ319^DIe3GOO&7Q2=^AV(0BgPTA18PZfWJePd<H;gQF=UN33YL+=#LdHUf._9]M
+(eS?gSGE>JY+GOQR#CBUO1L<bLJ@B[#J#f<,?.O:^0G<a/8)3QfP[ECJW#Y;=b5
/bS4LRg24/3=T_/=BQZ2f6[^Ud+^&368c<-WA^>(CZFF/LBdeIO^.14Bd3N&P>9=
K;T+ZW<>K+^LZd(d;eJRb8DT-/AMe@(?d&AeQ/<\F[YB^1=D^)G-XW#<_I9K)C@d
d;UaVbf)<99c?-NM.&a[@K&\RD6)(52ZNO]=G1gXJ6/<T782N6Z79e7H.JK9;DN=
Ue&[)XC4S7_QRREO5-Y3+#H(Bg;Za4H[X>)]U?)L4E?gGY^>Z\3J_H0W.B(7AS==
T2MR<D5g]NAIN9Oa4LdBLJ\aR#bB#[>VcU/cLZF4E2,?LZ?N8.3b380bKHUI7(J:
TZL3(6\UYKd.(2X[;_#f(R<.b\R:2U:f11ESXF1Da?NETH_][FLD62Z6=TG[3Eg:
9VP<><6S9,Ia&aSV)@UIWa[g8GdN1c5B9+TE6G28>&cEeDa.df&4R9A@C5-K:0KH
\#0M3QeW2WCAR5JM5U4WZWaB0NE9]L;Tg5JdVDNTKXYN2KAHL1?Qc)d973L5DIW)
9\X+@f@,bK2A[Pd17-OX,826a=b4L2D.Q/91IM&WJ#+f:YM)OO[S@[0T-b_QM:)(
54F:RcgA@bH<OC^N.YBf.U43gWXNS+KJ6bAI&d&8FcLg5E:e0&SFM>^ZI<VZBU6I
J4.GKM5YXSE/#YU^(?Y#<gc4V>J0D1+/W<f>8eIPGBW>c:dVQ8W.@Bf?^<VOc5;(
MdC:X+1?+ffA2=(T?;e&&/=_FW]H.:J8)JIdAfXWQ.3c-AK+b?=I?aV1a/;#:42f
Vb7/B=E//Y57;KU<6a9gH3AX<>:H=a:DC0CeP&SJ/R=Z2cZ@>.GeGO94gJ/.D/Ka
G6FQ]@&eG[gOcK5(A<)&^SFO+ZDfJ0Qd[X>8?aT><EQ(aZWWU,V&&3@R.G[PUQQ_
SabXXKI^aA]WMa&2bZWYY6(a)0R4?[4Mg_XPfHcCCdUg>1eE4.#75FbcTN7/L-TS
GH\SF+\>A2F:B@GXOTJDMd<e=MY]R:2FRW@TQACF]_]=FP3A/U[PPbTJ,dbKT7FT
0R#;IE<WC#1fb:B9,ZF5gf:XR.C#e\R@eg,;OCV?,dQ-B+cX44I;@89/5[fY?+J,
=4cBdI4_b=?;R8;U(g&@H1P;8CDgJ?T;7WgHD0?[1F\T)AX<d14[J;,,UG<RKK?T
=3KXQM[VT>f3(Fe<Q7+1O#BX;-W:O^C)PPAG?W;b)<dc5P]:8)][;FfV-TUK;)Q6
R,4MNYC#Qdd7#O@E9c@b#I=CbY[6f1Qa@,1N&=W+D)@gQ0MBf6E/6@MWK.8HgYS6
#I1eCcAWLVD(A>OD6DBB.LdW5_@)g7+PgGOF#U-6FK@3c#c.D_,CLA4,>AI@00N)
/(^eI3R)SW5>0Kd00g\?)&6[F[b=F;cg#F6T#XKX^(;0XPS2GZ80bT1CEH1->XWP
P[cXPcAV?WV/IWN1W\M_C7@aF#[?N=/<CGZe=-M.b?[#7EL^(20PG0e\DV=XdOdN
>\^9ea4D]6fg\@.-X[;>X:365NS,E8-bRf]A(V-F#,gYC.FJ0G=>@6D^U1F,KM:Q
.W2=1KO81WCcfBL-)IcDP\]@eX_4=V3=5M>34A>\C-T>X2+.JV8D8M&e;+Fe0Q;Q
)cAcL)GE4=70AcQPJ>-0:P3H5<OK##O#>@2cAX#T6E\N:QN;(FK#N>1^216&GQ8d
GP+VZI0/#c9ef6V\VU^?X:6VGQQ5gf(9\K8]@JAK.+2-8OEVG)N_U5]_THb.L#+1
+0+>8#J/2Jb]T)QAL/\d&/d-3M\9_>Bge81a?6<.)6](Cdb)[>E.^Ld_[9#gMS(e
6V)dgg-04^2g2P<D?O>^:RaWH75SV+RN1&PZeT,KVUJAbVBA>QX]^LJZ5UJ=cPZg
.\.IU]P4XgfK?bXbV,F54<1U#57[(15DJ>_/9g29QU=EB]^40.bBDAOBJ=fEP9=+
e)^G,(cdRL&+KNG_-CFEFRKPCQ]44C_@^6[0Z9Re:a9\gYg521[B13TRUYLR(=R,
OQ[+PRFC[Rf,&)G^#fgB(@&=1c0EK<81R2=f6)F-FTeYK-d2V^&\(2c8X2@fWO(+
T>MO/.e=TBS?6U#=_\fW8aa&)R]3CCZEE:3LTS<YSS6/@CF[O[_/M9CHANgG^FO-
G[>KNXPfS?]7BIN=6fN#IXdD#J?H1:?O^P2_Z<U]_E/3<MJGP5\_NR/9fI^d:NB;
D2VL6EK(Sca19A<.=<AE<.g&XeJ>J.<_,@:==d8&[A]:cM@PQ#&g&ccWZE.Z^eV_
0,#_]Z^/S#1VTJW:.#8A1-=]SU&0:YQ5[]L_2bWU3eFF,ZdY\f1Z6.Q6\I=T<>&&
eLHB@;XO@>;&X1^a^N3:#:MaUc6eBe/T2#_?,GfA9WMN9/4Q\]9LS#<]_TSALF9U
^J7PYGgWeVYagd807e9C+aZ7RXV#5KLKHcMU#U7RdOcOS_WSFC&e^A/A1.Q;T.I>
IC?>CL;BHLA1]LPX(=O[=[GFR\POYH\aG7\<eg3gYCYB3g<^aLD5BbZ\,QVH+87?
-/cGe,L>fKTeX)_F\A.CE;9+?5\:Q)GR<1P><N=J5QSM+CXJDX4,(N7C&&^T5Q?]
.=L:D?eVS)-Ob&JS[?IVdMcH0M9OJHe8Wf=NSBU_OI#D0:XdI.IY#Q0YCc<&H6JX
KECK:,X?B+\_B8QOM[&aT@&2b8@>aAWX1#E?LS<;95]^g(J55D1/:CF,Y7HUdMFb
6.>QS5JALgRPHILG/ASB^C0CBUg&391QEQJb7+D__W^W4(e:I8[79Z@P9+U_]P>?
W^R/f.9?XXJ6H_=Qd^[e#Y7NW6,c,Qf1OD(UgZHd<&<_I.Y=LE-K)CdJ-)H^-1gJ
+<YQ#NR.E0\IJ&U?3AMdK<MLV-=(B[T.4T52<EU@P.EgSF382@g@87I#9&N[TY-L
LMV@OF4c4RUMR(.#c/3<L]1N5R?Ie8WR=T;3<BMZQa,a04)?TLSL&_52YVSZ;F=-
]4=]Q2DF=/W5EOJ_GG2^gQFgUGEZI+NN_953Dg9\X3DZFdU58K0<NN<a;CA+0:OL
)(Z8;S<JRFCZIHS(RBXP9ZX]1,SQ:.(@AIcbLJD4fUBQB,c7?O@&H/#AE[aR8270
W=BXf.[?LW.?1R?M,-O2JF>8A\0;,>I0L)I0a:dJ<(8.HZ5d76&ZKBM]@&07(;MT
V6eJgEO-U<@4=-NWg+=3)F(L2P5cXMfAJY<]-AV?TCTF<RGG\+fF1D>U.#N_N;7#
e^)YD02dWe+8Zag/V>0_.Cc+.NNY:)bAMa&([D;:Y_6XRZSX=+=c\_6G?Z)(S06I
ZgaT:_Ze:\gfQfU]0gOU\4I1K>6eFc\X0DVU9Y0K_=cXX@-0S=&7/De\4,.GK0/6
Ef_MQV(.KW-</aF4e[A-F_C7)S_;=:.RQKD+&S@a\c_OF\ed]/)E=4XX2-MDP5Pc
?LYb;@-(QRX()9PU=0SAOM)R[7ULFNIXEBVa8_[9f_/gBg.^C7&H).=1f+?TE>G;
QZ8J/I.?dLge]JF?We&5@\TX8W;ZGf&S:e<??MM1]8K\1TeM]@A[FT3.UKZI1E[O
6C=F0(W\3J@O#E.cZAOS;0T>:8.dK-1YW(N5WF@Jf]=g=2]+=UV,ODUHS2MK_0TL
b]5/e>7g/](d=K]A?.[S@f-2&U4Hd3eF12>G9>G0H@dY51?F)@d6V1DCQa,=4f7:
cT)edcg>59FcD5-ffVe5B9)YOJ?EbO4C3@]>gA6+D&@\?C6H>9087[eb]7f6-OY7
5JVSO9<bDVW:J=H\WVKZ-]Q<V6T<f;aWa@E-WBVNHdA[AR7G=Nd6[g2:0/)c,4>A
W;M^GT?IHa+IOHQ(9gD?\=&9D0]X/+6TCZC:<\QWF8=0aHgWbQ(.Td5e#33b2TQ;
YG/()Q(c1)GE/cV=aZIb4[>[1d1.X68CRE-;FBMNPLb)L-M;9_2b@H)PC?b=KJ&.
.ZKX3b4862Zf(2&F-gDM,YA^IPKDb_AWfAL+FX(V925a8N1OD@^f+T32516#9D:<
&6b/Qb>g9fLJ<@>&(8\;8QKCc:X-X;VG^79E>?L>0#&CR:a=&aJ7):E9;5(3cO@a
P6D^eKHDE?AQQZT4U(BC(eV7+dA8f5TaI[f0b:E2Nb].95#J>B\F5cBeE6JbMeFG
UFCef:]TO&cXP0Z]H\3>MJHGBY,c-X/]N\UQ5AHUC[L\QE#5G#-P,f2-]-GX[/O2
LZ45.06Qa&U\N128\03e7^_Q]6ZZ1e+F@[4A7?5.-HKJ7)@QG:^Hd+F3g90JMI:G
B.VAT??XU@&Y<RedEZfP((7=O7;cF[\e>FbXUG1:/G0O:\b]TbYFIOP]E7@,^2K9
\=\C(Xf6?WM98O>))VM-MAf=L2F4D6-e0N,WA\FTU5/,W]MK,-?IV95-IJ0SPC93
ITg,LK^>(3eSVdYXOJ.KdV6W0G6K+=0A/c>VT2Z+FALFbX&1VJ/>TV\:@Y;cBBH6
Zf2U(ba/ORN;d@0M+U@&9DE3RO2gQ.;;BE57I\N\T2]+M+4@Q:.:BJ>W,H:8,9,1
eQ53ILNN,=[D:#DVaeI.cgaDK+F\K\4P40(@,]V)]<9A->^3MSVGB.>Z_f0^YRf,
V4Db=fMXReQ>bQEB.aXdMXR^M8Ag>Z/33O?UaWR);A19E_=)D0&)C^^e.=dXPSSL
UfZP\_C=H:8_c]H5T?BN<>S#ZF]\+2+FT.5IZ?aBKMa(O[8SZ>)F]dKRRD9[d92b
0YMe8(5,4\7Y4cabW6dFP+7<1=GdHM9aU2,63eR+Pd)9]\G#Vf[_-WAV1FSAVf66
QXCA;W>E7NbH1TG_;=eONP@K&]8J-SK&e^@FAKYP53,RY:HQ&IOba)3LW&NfRB)F
DWN24V&:KOP4Y]A\FOEF_O5Y[W3L;bHgGJ\Fb[XcCcM2)PZZ8QVDAg9:R&KD;P=g
fSMH/6\LP9.864:e6T:5fBY)Cd-0E@6B0L)Cg(U(V1^G,N21M[UadVI2Z7CG=/,-
YRIZ0fN=D_9)48J.gUT4a78c3NF=c(D&f:IXG\K&.^4/aI>TI2(:R1Ed3,bN(+4R
?7F<:gMeZ5_2M=bG8cdP^4O8O#BNIK/5HX(9N&^AG\cSTM\2e)=T4CT>5=ENfGe;
O5?>THd:ED<Zg.+>G,D;-eF:,=P8?3SP\\(?N,2WCLW2=f2]TBW.#3SQM<LbVC\L
8@O(4M-,G/D]+^Z)7@FM9;@]T/\+?W1JWfa5QTeDJ36R&5OMWWX,P,,67bd<cG=d
)X)e@<B^,,_SYZ2bIc^Q6f@]W(&?60+1<,>SR?ZJ07b.[>;gb?-fY7E2&1@&;IC,
;f0#&MId:e5E:Y,>@g>/.&6_-PTSVcWUeJ?LfVER667F:O-6,?]:,E-LRY9J;[(\
<aXEXH3_U,RbU_b;b6?QfG-<S90F,2:d5LWDLBQ??N,/Uge+^?M<f>+gb2P:Oa-4
06I23CR^_=EQN9b(FB(TSIUN(=4TZRS86\MIX?PK/QWc#/&EZ[_F.>H[5J4H2OLC
7A<HAaB@,(4N2N7=/RE+KK+</RNX)QMMZXeNU=2M.H:K&D;/3R=(<].O](@7aNAF
EX]g2.QOJDGB3+88a5eCD[[]?OX1<c#4\2@7e1+,[0W[GVTD??f_M_dO9#TA5AE#
>=>]S/0Y1,15N#=ZYgO5Fc>ff7Z3^\C.I7Gc8Z@]REY9>,E@L6;bUN+2T9=7e\P:
cVMF.4PNJAYPSA,?7?d#_QLBEgd@W\g^B+9fQPX^24@fQ:HJN,M#]RRW1?;LRE6V
Z,EX/T<c;HWH=\W]SM;S&HL4O[RL7f=\6ROLGN1K0aS(N@b#OVWa#0;:UI(/XC;-
RP)5/YTUKcbe:a+U]](OM:T=([gXD96S/^N02))F)D7FT@Cbc3e_;9,>K#Bc+].D
XgE5Ug=R,cE[6FNce.(SLB[)8<LZEG;+LH&A(A3b+b3eIA2Jf@)+1,2d/NTeZ6/#
]><X&gWTI15^^VZ_ff8DPH-@FHFD1=5,8^++Z1;D[a18CN:51N4<WWD]B+fJ/ETg
f&YeBA[cIQ0Q1(eWPE2T6/c=?)HHAMJae6L;AOBcXRPg0E#A_BG@EWRLQ/@.Ld:X
85dD1AA#A_Q]DO1H&[6(<=A=HF5?L@1>,\@>-X_Y3C,1?W4F3UL:b>7ScX_AD#+/
([\J&fc>7=N)0>?.9WS&^Z0]6eYH3,;]98VYRRfI9:Y^CKKD<J)7,X[/SB/T9ZK3
1L<O??ZD/<59Kd^SNgOgfDS^5BB=+GZ4<DIcDSNDAF/G;N;00O:T-EZgU_R@DJ0R
5UJGX3A1BJ=];@^AV6fW8V]7V2M_3e\>XORSBE+B\&]H3I@OP\WEL15V@]NOO=fB
;g3+JH1U>egCI(^U=MX,[C:>ZC=]DH-(/>5;bY62aV5<)D=ZIS1E(I^7;<+HMRT9
D4OeP5D,[Gb4#b=9H\3gHZ,8FF1^7(ZeVDFS02XH5bHZW_9_N]?4?DU4.feU#U@I
7\#W^TUSVEF>;3UE&3AfLcW,gT)I5#E>f&E+V,]0P<d:>?PGDf.QAGeQ_aYD/4A4
(RH8c9aa@D-KZd#+53T0S<^+=Da_#F(O#B23<bK0Z:FD6OLBPdHKBT.b@Z>eZ@U_
2gL(W+A]I&@;HcV[T0W0YG.f5bcYde4Y\MTP3e:d?2R4>R-9>3\=bOd4M=8OQ;8(
OOJJOQ9KCC6bB]]VC25E3UO?T66BdQU-C6^;GK^>bF5TV#\>8OaU9^DAQKf7g,E/
Y6]6+VfQG2b96ddOLe87W[P]MTP@.bT9?AHZUF<P/UW3Ma4-TV_cCbWP@J;Q\IcS
&]X<(T-QG8bL+5RZTU3M,BNB:L&D.7Q,@[F]KW.O^5L##/G>YW(AWD50cZ;ESNCC
gZfB8(2F(S52-Jf.4C[#]JCFb))a&CV9_D&D=+)Hb:;(K>6:/#@CI:^8T@\,&4F1
#:4g98MKae3V:28],2#2gC6a88ZM49FPW_HD\GC?B/[Y6TJG@UePL^#+:^A7#_1H
Q5LY]@WGg9Z5BAT/=GVa8+]SfgZTAARL];I#37Bg2E]gH/(ZXYP9A.RIS@.OYfHb
2g0e4ER==NTbKcY]_@<L3=3bPBSdR_eZ1ce;<)XCfU+-.]@3W=bL(#CW/>+,\AH=
KcU/++;52V&8O(dPRTXE;?_O?4=@;[LB_IH68#Vd>J-_^HPgWeD?/WeSQM?H-7UC
SEcSOGJ?T?VCMD5B\HS/D4^6f^^146E\:+6UQc8fJ]&R#92>[>[;]L+IK)J;b0F0
5<.d[I7-R+(MEA6EHUOAbUU+<3S-GKMb=,.@f5N7<DP/@RD(+Y+6X71a-:,F?XKc
cP;,L&<Qg#,]Ge\>S/RE>bG7W.5:e?eWd6Z0([-.E[5DR=[-b6Hd[/:2YG&_@4ZY
TaMFfP3Kc(87I2YSUGLU5KTFaQ19f-9cISeL/Y9+;#QZ\AcVXM2eb#>82Q\,#>R/
0+RbFbLNOPX<\McAC<a9LGR&UZ=T2G2>([_A>M75/=K4RH0A8=TD3.cGVc+B/XA;
B&U,_S2acIQIFgg&IV:gOJB],]H0XGXK@0bD@2^]_RRfS9G\J,-6T.0DGG?SIE^@
TS??30CW[JZ\IAe/TFR\>(789>R+QK4FcP(-bN)U6_)S0>+U9c6L_9-5,<69Y=H(
-4Rd1P,,/ZD]Ce&7@GNOW)b9;G7ec6U_)0R,U0;F+@DdSGTc\QPY;150DH<V8WDg
=H5EB+)H4[EL=7eC\;&dD2/B>>BN92F;3RKIgJ37931c1P.XU3Y^-RbH&6ZL#N1I
;L(a>6b?2df?d<a+93X#/<R0[30DXS=gQY^_;G1b_WFKBN4MO^BSb6fP4X\]G3g3
5:<[##]aOABG_P6&M5MZ3W2#)U?#^eIHQ:WW.8BUC]d>2K[bH\F;;\ZdgCEU8MUA
YJ:NZ?9f8D05.5\>#PH&dLD\Bd<U=BY2;M,FcQf7)O2U:b#EK77MUAAHVgSH=K)M
35ORaQ>e36WUSFaK]ZYC_<;/3=PFWf-HSb0KJdE6,/;=\2P_BPE#O_#Za>S[/c,8
+D_MKEAJJd33F9BdR#VTE(7@;W9?5NV6NANA;ZW20F:7X\.80HUFSL;fZNCJfGE:
eV[Ma)b-[C5&6=ZU4g/#W#VM^ZBP(Kg),TBDNb_>Q\H7Y,/(W>]TAXW)DQ<_&Og4
V9&2]LK:)1=PF.48Q5H.Zdb<DTBH8M8NVZe1(<a-J#OXG=YeKW48fT@VNX&f?V7D
LEcCg4JWWP]T29.KUbFe[>bDS/1ACc[S?aZ6I:g05E?F@/>f#dCUUC-7\UXL]GV=
MXT\C8OZ2bSKM)IJdMCZ.:]UYd^dO)TJaY&DQC6Y-]]c?\#GeAaLCLf1JFTD^J,3
[bFNG#g-ME(d6BG&+fd6^QUPMHM.@HZ7b\6J2,QSHWM6d5>BM&-)]?XV^2N_88dg
f783/P@Ad1(?W#6KMW6R#I_N@COY8QdOZS]A&Z+2NA9(.EMA]DQgR;af3V4V?dH[
A;XO/VLV^a00_a&N\#+H,c,1;G(P)[CcQ.8R.]#\6=P]#OP(BU.Y>)EY\.Q907^^
C[^S&#(EH_/K;FUA[\6HJPQ/L.+[X,F^F?VR3=6P#:g\-?6Q[(PP?#3C&7/9?SMQ
^LBB:UK3(=Bd0GY=/+^&W3#df&Ad-B3a5f-]N>Hg,.Ld+@3I[A-9C?)JRdCB>b#7
U<BL[6+OMFUQY;INC/Q7E=?8OC7dJ9K5[NWM@)/=RC0E-\<9<5@0Y(:PZ]2@/12F
b->eHEHN?[EI9(OeV_\&2,S1J/2[M^VZaO+BN1.(8>Y)DM.),/+b?DaQGLW]bNfe
N,0YBR_SLL[I:TgMKNQaYbLe]/X+,IS5f9I+X/Z([B76@=fgJA0^cXQEIG10@#;:
(R(aUL<;[5,RZ0X]C0+c3aR^V5;O<9I[;IW;K[S0K#@d=UbdO:7?QcGU9DM\NZ2J
ac5QD_=U@^a@N/K<)O[<?QI222;?-63fQTD0O8QSXffNfa&>H:6d>cMN(&1A&cJ0
PGfT)a&A.8<1]AS+=3:3Gf@-faD@_E?)LBVEFW<+PFI\,F97a2Ce3<e>\:QT>=;(
C(fC/[,A#,N9[fO+d/;2DgZ(gX?e_W5.Ca10A@5K/V=QO/T;;M9\T(OT1Ad+R)C:
6((cKVR4Tg?]:N&6.Nd+ETY\&K.#<^CeF3PB,RG4Waf[8K<&F[Bg=FHG=UH3B:B<
N305g:aBLHB5ff-BX<CX:]3Na&X&AO,)N?>[9BGE40>QHS@TePGK/SN=XP46U=Wb
W_=?_+?^ACaCSfY+0(ObP@QcMbKc#?-(aX;#=a15\3#UZacN0=O/9AD@FE&V[&>Q
_,02MO?#RJ4H0a[b4_P,8)e=H[=7Dg+@3#-a0N9I.8=Q3YKW2Y/ZXZZ@P9_f(Q@T
<W=B;O4C2V:(G=5[;ac^ZN+#\JUFX4@Y&3b8cJa_>fL\P]\W-E9NeM9&=RW0A-7O
U>Pgf=c?VW[bTB=&U)0BR/PI50GSGYQD;L]d:PYTKIdXO5cSAXE(G:)e<+3#S)fG
#\4.1=_>PcNa?1KH54TC3<Pe<a-;EPGX=JD?XH0K6K1dP@B8Ra(B?HO6<3HPD(XZ
(eXD1ZNB@[CXFUTHW##XE+?g(84L(A,P9Y.#>Ae&-_2\R4Z85e#ZA[OT=GF;cTIF
3K>_MYUSFKb#-]gJ&c@QR0@/X0Z[NC=<(+\MW<F@GQ](R.S>FO?[NAW;7?;#7f2e
I\W^fRTM)PK&DF4UOdNUV:[>96(JO^d[SgD#Nf,PI)HSKXNPGVEUdW5023Y6FJ)3
Wf+-3ARVD<<BZO2X?.,NJ\SQ;2DS62&N?,R/cY+4X+455IM;ZdBQ;d=H:_7AeRFA
J2g+/F[Lf,WE)_7=BJ>]MIc]+30I8Y>DCSScc8g55^.=>g8U5W\22U9WZ[N#C7.O
WDOK;FcfA:[&-4C\\J@;YSP_]@_Pe5]=e2U)RCf.=3,=FH4D)6S9NV@V8W0.6<dP
M,C-]f:M@C&TN=\]3CbV:C+;[=g@+d)+P#4+[/)@LP@1/\M:0>1?IF[MTMfIcHdM
]S+?^?_LaGa0\J,:.eSdTY1eWJZ4/1HMaJ(]<[_-gG;K:I:Y_cY.V&@1fX9,XBSc
NAZ>@Qa;W/CdM1/CAPAZg[>)<//:C)UD6+U>&FgeZG<_RegDHQOJRP&)>UOVHfg5
3=M>@_;G33<5[OP_Q21W_c;\D(J_B@>A<e-be2WIU(06Hc6F7(;(a\3DdOROPS#I
3+BU_^GBS^4-IM@RW9VZ84XAL#Ma\Z((3L3gOZ][ZK)GE\OF:N5.:M-M>,^=Y8a\
S^JA:=)P#G)=d?bX^K-\C1(U6A.=SAf>RYK3-<[S/]JV5KPb?365CACT.Ie.GT@f
(PFCQ>H3#:_fDgR(_1+^]dQeETX9PK9XSRW[7<TM8DM32GHX\9M8e(4fJ^GAG9(/
@Y+OVS[4Y4<MESJGU&6e^JE^WK,^g/OYMV5I]da+U_[3^K>eNTBQ<U>d/H=;E0IL
Q/^)]U_Ke@B(WbEO0;+&)cLF>e=-;;[CFX5>X3:eaK1<OF&YW(4FE-a9OG&Nc#2a
Sg51W[>]XIN5#S,_CIB\;?]c857Y^A(b>&KBFID;86e([b@CaP/I6@Q_f^,Q?KW>
6DF;d1_X/5F#^O^JZ]:+d++a/ELT]&ggL:&Y47YJDK#GT;B71OYQdAZ3E2UC\V@Z
R6JaSA+4D=B:G_\0)SZb=F&C83(>bR\ZL\f?-fFQY0_;gUDZfM4?<BWd7(_:>5:(
]#^d,eSS]5cg1)gSC124XF.dSE9^@(/)[C&)F-BWUISO&_5)<CCDQUJ#F.G7f?IX
ZMURYSWG+C&(D0FNU&<d&cE2fXO+8d5O?GKJ/J#fZDUM234-O#E2C\..N_I0ef\0
?H0Ne#+I\)9f,#S4[<5=0WRNJ^MY4,>J[^F>eA#HLM+G.gg9^a1()\TYR@JAVgIR
;SJXY8a\[JW=B-OO9=(UWL0P&@9GU^&Ue8GN@cdL[c4U+N,P#KdM,FNM&/VD<J/6
S3a5WKXS_Y5[M)#,E)/)OJ0Z]eUAEc#(\RH0^Z(AJAf-3V:E\C_>^DfPBe[EO>T.
7[&3SgI].->P4LO-KM\8f=+?]2PEMSR#b>#K+MGE^YN]d:)EgM1G6+ee\8/WJG5,
?C6U2W5E=,803O^UY3MVT&CZf@]NOK4D8NC445=6L2TANCL5U-@/M1]#L?]0QMVf
3J6cHa@FWE)cH3P>b/W=]H=:SXT]0U0[N@C1DBD;TQ31GZ80BT&K^+ggX6((e:6g
fcMCK>TEP^8;(#]gYA]XUTFPgQ05N(VWQ>N0C[UWCK)R(:&>3^)>T:PFB9g.<=^[
e1(/dJ]QY6YRW3[L:JB>JaSY_>TZ9RN32&g^-:/WY=^H6E+Z?#POHNW4dgNe[bY0
bfZWOQ?@GE,cR[8E\[86(HH10,N7EG6N2+7a8A2Jafc\H9[LBV.AHS]bHMB23)QB
QC[:,ZEM=BSL._Ac5fScWSIT4R(a/&_U44MX4fLJHRN5c8C()Ud[4;\ad_UHR7HF
6aDa?/(IZ8g?(EY&V=6.0]3e_V87Ged4d59M1@;+6N7ab59S6f_4g_S?57>ANZF:
L>+0eM?c8F/5[dbK;:044DB6\O(WP=gHN2W0Ue\>W4X:\<TXK&?Ha8Uf)C_[P/+>
&.+Q#dV,SFMfCfXF/MC/6:#.FQH2YZY:4fdEg,9Lbc@&^:S16>U<S6P_+D.M1-O-
?J7[),\T[=0Q58[0X>Teb5V5eUC?fYgB1ZAS,;.X.b]^E(58_N50S[AZ\T+<de0X
N[dd5e_1/QR.AV,1[XOJR<b@WFM<MR,YRd(FEC8_JTZBU+-a)^b\.<UdHWD-0<cP
5G+S_?9E/ObBU;@=7@),Q[BLYQOLKUa)OAR:]JFCcP1_G6/G,&L,SYGeS^cD[DW1
PgV#(A>L:2-O+A3;O#<M+YWgHV&,U67-0a@N#JE/)9Df=cb?gAB,<7@/O,T7fSR\
A6JZECR0W1JF,WUbE9LA^8g]F_cSZIM<;F7c6ZN^<[7\ZM.FL\@@dbQS3@:AfIf1
#;L)7_X4CY=QZf]Q8AX-agZZgAHH(Ua>_>:U]LIDE:5@>NWa#0A6d@/SJ=_O7),K
C<>KfU:5XQ\eT_44_I=FJ]P/]VL(;E]I.dQ()V78P6&JYPX()HW8^#\ce#>Ed49#
dLJ6UXC.+Y(;\K&V+bAdc>/<a2H:Cb0>2f=R3S7<4/IVddLQNHedW+31G?&UB4RP
L)4f#T]\V5^,P2cI.,YR4caN04(\a+(Lb>472/80U1^5.KU,L-\4dCU[9Wd2+4b4
LLXLgL3;HU@cXI+-SgE:_7<aG2YUabEGVFa@9Xab3QIMK8@#61F,E85F:c@cG(^e
D16YU&+gc\Mb?&P<+UZAC+7@Z97dU]RS=ff\O]\AO\KN@0F(FH-CSIES1V&<BF?T
GgKcKWZCIgQ(]ffbWH_;/Hf:.@X>,+/UWL6U#H^LD2Eb^K9WU3U_C307DYDN0fV=
O-#f>FP9S3Y#QHNC72S<Q#,Q+RBJ[]VRD-./&9?+;bfF0(f4aMEeA34O?UBLM5e9
E^JA5+(\<\YVPM][#:\?RW..-RF#<2/.DKZ#P2:1ee>1A3)=2O^]_G&#)?H\Y>X>
M52Z@080P&RPX/:<(BYZ9[e_^#HHH\M\BgJGQK<<>;092\?D]\.(0J](ZbG3C=T.
Kc+?IaXR.W-5J4T9YeeB#_NIKN@AaM@3B?(LaB5&(#(,5b>^,G_JCc;J7&YQP&I6
=T6DN)dT^-c38\9<3Wc&TYVRGG@E@D]#OT2W9:XEIQaSP<Y?8]M_X;3R0<Of\01B
GUaCW]Q/g(#&EbQ.RTeWLUN(P9g.<//VKFL9>Q8-(bWOLLBf4ZV^))8MG,S3;2?K
U59)/g]gUZg0<f^EFA6#S[cZe)b1MSS-)M11b>7=R_=bA5S6OgE2RS9CQ:-+[LU6
gCcCYSV<.(1?&A\?UNC9/;D?/Tg?V9bFY[g;U(CObT_V7@28KRgcOaG4Y2WPOK4B
\\ZMKfDXS>OAcB@R;D/RX;94ZB6EP/;._7(eMK)f)1geX2d1=b;_&e5[HgfGc.g/
#:=]T(<Qa_XT:N#=QYg;[6(8;D570P<6[^YK1+L\02(:+&R=SHYG+I0V)I<90c:f
K5RLKe;Q&Y3[-:0dNFXdV=4,O\0R^+5)cIBLSfX&@M#Ug[E:..#a1[6Ac(8,V]G(
1=)/:RaB5#=e-eM:AA2VKb[[))f;M535(Q^PH0N,47MP3RX<]DZ:OKH/TF:QTBSC
,a0@NS_D5R.;_\BNS=7ca+G949N,89P&S.=3,(>@aFVRA,^Pb>;OHgfURE5ee[(J
>b..QOB@PgYS(UFB8?Q0H[E[>LaZRIFd1JbL6]MU>2IR,g;VYEQ3=XUc#G=fPW(O
9-45H[\4<2aA#;D/=:??7N0M/1bM)=>X&2+<4LQ=d;>7/]Oc;].<457=LO6@AVd+
QW(14VDd1KFfH7A?_eCeb9d5N4B(TTP3aD.U[9De2(JV4Xa;VeG9K2Oa3;Z<GG6f
fC@8b<:8([e69O<D[a:b7&S-U+1LHfXM-)^d8&=WY6Q/H;dK.-7gGN3Ia/3,Xf&P
;.;CCeCc^ED4c,4.gTE.fH&T@2G;[>W&d[7fHP#TbWL#:I2U3L:B2g:+aO1(8)dR
K7CX5TLg:VH,_J+@HT[#0F[HYIF^1Og,_-9UW<1,Z8W98OX1d==Ge&MQCHY-</@J
9ZXZdeRW1dDECa[GdAg21W@^D2#^Za3>WfZ?GWfL=:a=(I0_L98.>HF<V)cVUW4S
E\RL\:(8I&]bQNJVdFT<CdE8&]MK@=7/-@C3RL1c#O)8U5a?3TT;^917,VRPgCEe
>OI<F^<[<LZ/E(#N\Q#bXdRa1dV_,T[JD\0FTV.R4d^)0]YOTRB9EZ@(1c&(Q#;d
[.TdUWI5,)PZ,2[GO,d]L[ff/(@dJULE6MC.O1E25\8c6KJ]^DC<N_A3E[93V]dA
@>.f]H@=?Z8F_c];d;HJ_:G-&^F[V_;d^K7,R0]V,I_eA_Y=C>(TTO/c(Q/a&6K#
-U>]XObJgB^[#OB\+F&Q62G]S@(O;T(G;I:.>\19([^fZAT<dSG8Xa@L>#DW50&J
&W.43#/=U/Pa4+CS7#Q\_+1&+2<T:?;)25c2-6&&1/IIQK#aKQBE\Ie=5d#4+STZ
Z&2F1d/YeTEM8W/QP:(ATJUQS9UJ/9QE\9WgRBZ10R6103VbNbI4DaUaOQ=6#4Xa
eJ@:G97V9EO@J]VRYb1g)Y.:We_d4HMD>A6/H\W]OW-CX9YE>1ASV^PZYJ<VI8RM
M5;A<DEG^;^#HWRSc2[_NcDeYZL)ZZ>Wg-SG^]HV]4HDe>A/-OHd<B,4M>U(VE#Y
Ud9dUL.>af4>D[V[_.5E\(CLRVI26gM\T3R64:fR4<NO&8@E]8_bGI-f@M)5F.gD
PM-5;\9e9^a_fG-8#?^fD1?+KUg\8bfWL9+[-9/bFG)/^([E8g:X;P^HDQ=ISL05
4>Q6&Q-S@?,^H<=9d=IIZQO]<55VXP2+UC7T-5d8FVTbY9N)eG&M12;1)]LbVUS-
X)AEg-5YZ?AE=S_(]]gX-aKE#\LI2L6MW-^BRa)RP1KWK2SN5b3V,9X3O^V9.1M&
&T+^S)KB&J02>W=),;=OQPD:B([&?L:&0VWKS4E<>P<eW=].:HWd2)>>JHYY+Z)-
PDRHcO4[D/@[[67JG+BCZ&K7EIT,G1:H(&KZLH7EGI0bd(Q<9]9WDS):c4?N+11P
JB?[-)PTE5,0+)<CMc),b9QT.g.TWHV?B7\[^^?.g)=+g_)B(?](MAB(0F-+\WQ]
&57&b9^)[7;P[0#Ug0,M7F@fZ:8T2S?+7E5J57+:?3-6YT5d4<,GS_PT.H7MG(1J
Ug>T\_<^)M^MFUJV^UcW=4WRO6R+SSLb1B)ZJ1:[U=FT[Rdf#f\#O79U?Q7N<,Sb
NgKS4TEU&IT43BcXU(9Z2.UO4+=&8]7=H<LGT>e:eFR1?WCbCfEVg/0X<KJT[B/F
9WX5=XWJ9+@ST).5XVaIH<CagTL\^\_[RSX-fX)O13L;>LFFBQS0J-++]>:Q\53K
Ng:S:/@Bg<&2;-9^OIZ2DVF\:KQG2?CGfXWMH7HBb:cg@ZI@U1VYKW>_S&.#U?_6
2PJ.8XfAOAJB2A/gK>a4CC[]UUWYKO\DV4,5=+?.+b3R=+]cKEKcD6@P#8P5K4]8
#CT_c\II^XC.=&;7FI[9#EVSZZF9]Mg9bZ(7,^08\XSb7DK.]gKI?#6P1_MG9V31
g,TEBUH0Q(1X(9SLa+O@[:)SNcaDE)8F7]:D.^P;<\U,b1>(0BXYHL?1Ea^5E+B9
dK5I@Z699YYL]0_0O]6T-PHI)-Z,O^&2GGQ<0M8O^ZP)+MF3bdZU@[=QLG/9_O+9
g0WT)cVT?FW/T=PLd_QU@f0R0W+U+I,KZYRWf0=LMgZ@f1HE-JP/.#MY&KVTMGR+
I(NIBH&@=8JI1bEC5O(geGB59C85;]g&FT,&H<(P>6X,6[gYN9RCE.7)3H03+&(_
.U-F.G<6X,O2<FFA_\-+Z7=QK=-_>MgM3(XUK6+SB?gg32R(++cZP#FQ79F[fR4Q
M](),K9Hd5)C.L4(Z;WGAC1O[4R3>DO0gK^W/:c,?#=1.+]GVFSF^:C8ZOR3:;K4
:90[DP@>[?&</2UN3)fF&/V4<G^6)W-V@E\K[P3#)A^=:eMKDDY:B86(#TI^I]/g
#[8a=N_Z.VSRU^T>P/TWR8QAPEc0EJ1^.BNVOcB.OGHFef,_(7M2/7.KSGeJGcIC
@+LOPOc/,8-U]e\Tg,#XS=Q/D#YH0IEd?1]7a2aFNef_g@Hd3QH.g-6G-,37?MMI
E767::QY-+>4^G\:CbK_@)R_TR.M+&XL&gW];K7[GJ;;7MY8XV;LA#EW/H<CdWeA
C37OQ<6g2gTg>3/6?PK.VO(-b<N0)adFO)I_0dU.Ua;0e@2UNJ8gR:;5[=8DP:K5
C04ND.\=I[KHS,9SN88/5a;8g^eEM/3(.6WA_4YG>HTGOeaA5SYP7cBC0?3F)WT^
d)9(\9@IJ6@SUL\TZca)DfJBb/)E1DKUI&c?O<R7PD:&9(9+)P.RDV9RN5B^8OZ5
MID9\(gS<f_G)b==-U+KGgDW9gZK79A<>)cTQc&XI82V=Na<7QW8PZ#5J47I8UaK
Rf/Feg](+QK&+W4#<2Cb\bbDK@^_9<f;5TM,,IZ/DQRBOM50H61,5?(ad<?>?RY.
&dR\faeMbg&49QSX\FN;7)EXaTCdW8aZ@(IL[G.#,aI8-9E3UG\CY>LQdZK^c(fK
#NRVa[788@Yb><A??ba8QR7XGB4L>c1)P[@/aGNKJNDCc.@C8<(eFf<f5^R1LP,,
-Lc#&+M,^PMD8)4XOK[dg7F-dFTDeF@R+TeF#6I/Kb3]fSAX]f]06B)7G(a8B0P0
BCBAfG?&E[eZJ<CW2=XS16OgBD.cbVa;-<fg[@IO8_8IX73-CE#C10dO/^MS(MF4
&>L)?(=,=g8;[KPU3Ca.3EZCb0B9+9]G\=]_5/<<3QE;F5:L+7SQG(=9#]4+UdJ@
S\a<X/3L9:JW3<XH(=^(J6<2/6E+U/F6=DW:N3\&#7[A:F\8H>#aL&;3]_V1P0&X
C?+44=c\_-.1d;9WK9&JY&YM.UEWSeKZVH]K>b]EN?bTN(^/O\P#N^\A9E\U<)UK
@BAf=BID2OC9LN?He72OFVS-f2fBeVX8Mg@e0>V;<<?RU\WSRD(@=N@;d^.>d/+H
f5>X7J4&,]EI7;gJCOC>,2QHO(E:Ja>-W[96_WDZJWY>aY(GaT5R\E7&gAO.3,J7
YEeWX:VUg54TOUSFR3.PJ_9>P&WaW>43V,4<H9C.F75#NU9Mb+eXZF4:Z/,)[c7O
Z[Pb3b7):1<G[UMOW>SRIVGNVZ/9D621\E&=H2^3cP9XS^Y=Z=6RI?e\.EVNa.&K
997AfGC&P]GBe@SI?OD072VR\6TI5\Y&_QgBULVNRR)B8_W&]+IE_[>P]_3Z(8Ga
g;>Hb/S:OV(6aZAaV0?O=9Rf\]Pc^8YAB,_RPHb#F=f8#K^DbL]bS8IGW4>S1A0M
P;d_K^E(-a9eVE/?XK,W4bLKZP:_:/)W0+(FJc0K-?):=_SWeV^OA]-Y^2Z\JTQ(
DO#5)WA7[eJD;Mg;[J\WGb3>GBCO(f-4QP6/,KW@eL]]X;)F/@X23?.>F54PC/>5
SQfU3G,=?c]F5fTI72):TQ440U]/;1>C6H6?g[3L)9:_5a\:\(X676V.=9LW1OOD
7E(<F\]H58MTa-?;6)U#:WT(QUM:gg9?ES#R(L2Wf.fRFI+BVg[cW;d+1_I\[/K1
,NY>Qe]6c\HO/0)T&F^X&J/1:P[eRa_/9M]O&;TRI(&d).VX[#=^ARb<ZWOP,[)3
(9UVP6_-9d9^?8+@)d<c.eG(I2+=bM0KM=XM<)6>?M^,JfS=THN,^^[N3g\?HYMA
@87O@&[g8-L=B&L9fED)b;_WGPaNa=aDAXf^-<BBIeNQQF6M1SJQ8L@X\H,==XU4
-EF(.:fXMUd)P=OM9,4gTA@:ZBS:ET-2L&[/gKKY3B_Rc[2;SRKS9GO,6gW10HRc
EVTL#4KRI](.Qf7]D=(@::^7=1<,X?1CXW8ONDEKSBSb^N-C/V^D;_^7dc9eI?c3
KJf.IR8BN8@[KbU#GAB^e:7009/F,]Ja&^CP?X+,Z9OP?15JT_T3NTNd5G-)bZdX
C/_S]-^)V-TRAJ5C-Q7(2QB8)=I45=;,,?B?/N(XDSJ>FTQKWO75U,3b5J[dQcaM
&-@#I/AB:/=L=-SKSU8F./c&:S>c>d\M.9,fJXVCc&8FDYdBg0R3B<NT8;_^6E]d
.+P6@B,a7D99,g32TCe/aN60BbY.XA;4&29O\D>c]8BM\C&_>GgJP51J1#2):T_F
4:7+VP?aWVA,L^<g.c2UFGVR#V_;FaUG;A=3cK.IS84b_JR+ZDIIRa=/D<[g6-bS
1:_&J4)O];\O(:E=<.,+7U0[H<).KHBZL=aceH8WRN-/-P78Afa-?OY&JCG:dL(Q
.ZWffVX\Q>CVd7=0_4/W7C5)GCHOG>+CYg)#O2>T3>.?-19JHA=61P?-b>2]R>EH
T0a)Je?^,U[a@<a14P(Q8BCg]gg99,N7:4O=9&LYg,8cF6@:F6eMX^a>R^Q,S/<S
2ZbcA#FI9d[Jg?HD+\b<ZHTV5+S\5Tc_W(V7X&K,7_9&IA70).?@\IUb.=1U<Hf:
6IbN:H;aW<QO_baQ\]LIa)Z^XQI[ULJ/C[,0VML0]fYd3L_@V=5:Wb7PQT^?fTA2
U,UMedU9gdBPQ0c9:?\LV2@A6CF_9EYDc=+MB\+,fE(BBXTS(-TTBPBB=1S]6[Hd
8-A,YGRM7>@VZa<=WDR/V02fQCT=b(P746@0PG=0)L<\G6K_G49TG;94=L=18\=X
3)<1.gUP@OXe-;]D(V4,g-bQ<Aa72CB=Ib>_R?CJb4C8EQKcaSTDFP4A;+NRgEZ[
@=RC2JEZR?W4]VVM,A2<0d77S&957UF?1]#5.)FHABc;dLdE1,aWVT=-41&EFC6L
=5)0-8OJM\NEQI5Y\bgJ;P;?RLa,M,&W,_f<-=&^P#02IZ1):5\Q0gQR4a_B>UB[
)[NNPNJ33&EDMC]+_<]YX6I=_dJ^bO3</fNU<(af\=I[>b5&XbX9^6c8?U(29Ce?
6fDg,(T6:<=;<EGNMF=Z.EI8F9],YK@T25GXQ2<^gAZYR>X4J42ME0b9H]B:W<2N
>@VE,LC)1QL8e1D+@:^9R<:Q]f<F;,O8[M=8,C2DJ_;aaOF\HD)JbS+R51(J6=_6
>;fTcD#YR11#1^+[T<R,D<I,:?A@#Q[J)8#;W@7cYMBRS[UHU0Aa@7RZeT+eNc1A
\E:+4BM^DaNeQ(NcQEBW(5QQEQG_R#cT]H<1YV,(24]7AL^eYK<J<A<J0+2VG(/;
]_d/+O>-d/P[b\13^e6g^(B;?Lc/L)U<H>L.VeKJ9]D7cA?K:CBAC,8>CKaEY:K@
QUMYD+U+6ce/\3#E.;)<_d)aG5^ZHN?,LYG@/cYdCS+5f@5O+@cV./:@cOda&WMV
8/JLW04N9a>HV-\95Y@@F,EW6[UERL\/GW_VRQ=L1BQ4:AX=NJ<M<XOJ&\CKE[?V
N_37_:)^V8&6EOUBbFM?_A8^6=fH)AL(<U@URQ6[ddQX9)]]35=R7BW/4?9)2V<M
)(Kd(XUA5\9DP49M&TYQT\6X2<K,)9eSC-O#88]+1N56)>Sf0N@KFHL6^PbWG425
J]VU)(aLO<DZM24gIP9)--L&cL+WQWgY_<+L^,WA).eDNEHKb+aG>7)3DO?-0[P&
#PJDLLf/XOFXQT=PVdOH^,3g.f3NYdAD2ILFQ):42EDbQZVSgQD80]-1K=f@@+aQ
7fc:N59I1/bc8I)D=44b8ZB+87P\BXY)FDb(/KT8X+,^Q69&8H9JW]CA.F9J#4T?
Y2JMJ>OBN:ET9MRWR(,EO]5GE9>Yb?W(ZY@Ra[RXCc[UQ151MP_X:_O5.\PV,LTT
FHZ+Q]#1eC#T6;LWgX>(V+0IeDc^6]d&U5YE5I2@2]NLBaP?gM6E2Z7M]_)5D,#Y
W^TYLMcSX)dUe8N\[F0CZT5N)ba7J4T0X[;-a3FR)#D-;SScScDEYB0BRQQb_0L9
WWZ2NJ^A(PS7&?M:OQE:YVK1(XD&L_QDMH_+F1DV4?-8I6:;JVPB2KUB8;g]=XA]
JS0C;]:SK(<1UDJ8f7Q@I8]?UZU3]Z<CHC7H_1e/.8N1Pb^GI3[RCMg+S@AHO:g/
d.(<R.1dR7(A1E6BOHd-D.3Q]c8^fE/6Oc]Cg]6&]X2b&EbE\XWZ^aEXaY..SY:^
dacLKYZbYJ>dJY<_UE0_]7OcG(>>aA]G.#bR<4[S(\>IZ#TAZ3.H]QLR&1_DDW=2
6(5<BS79&QS?^dTWI9OSDS_=&R+/)aFSdSgg.53H]&9]H@fJ34M32#1\2dWZeKB6
)Ga&]UZTP^Q>6b-&.@_UCER.3J_)aNXgHZ<K@5Vf]W3/f5WOU+L0d+Gf>:&18c1e
\Te51]XYI@Z@9f\<;PE-M),gAFeY?]F-7Ma+gV8Y9WU]R7FV?TbA9cVXK[98(RZ?
&QTS?=XEM,8,3+3UVCD2JS4R#GR24EB?4)_e)gc_;^c-RU_PVdB83gC_TSD\DTe.
WD\SN7T^>FbgcE.DJYc@?>AHgOVHR.(De\88<B6#IT+01f.X]KTJ=C;.dLN2S]2B
?_4&g)(GG4T;a60C+cH6M;NfXCa/bbFD+9c<a\,>9^Oe>XaY@4[b1>g[Z5OD=0L7
-,61e3A@]d2dTX\+4?HM<N;1ccLaFGZIB4fQ3==WEAZM\8DR-Q6S[e5.-/\TGJJ0
DNXERIa?T,4.J[6VUFO(@200(fV5H71.8VK?[(>.U8(9W=U(C3/aF#,78]0:?74@
^M9^/17L:B&B6/gHM^\aFW,1A5-;[YL-+)3\aP6HbYT4BZMU56=5A_aA6B\4FV+]
&Tf9MD4VLdB-<QJQ0)J56Y&:(H\eX.d-gS(=#:g4B5DS</5^(HIHY=G17KQ;2V]B
ga\_DZJE0W\FE4=FSFQKEP8^;H&ZeB&P+Z=+W3N47U6Q-DN/[9BP5D_(UKO,HT&(
U&/A+e_1c4/gQ4LO17K_=(LM9,J]BV-LQ#W@SA_9G0X6ceaFE)H52Ee9TP9^+b#f
fda_:G1\SDF6.X7RVU.]TXIGbBIV4W/F[/4b(2]YaBdGF@17L=Z[e/V6?1cAgY1I
C0_\:?#T<_@[R#(a.YPM-e8J>AEQB/+=Y=PO^4=Rd2TaaRA[]OFRfeROXO5-ZG#Q
HEFGB^U/<WC.JW#eZE^c5(#8e#8/9E(+Q2baM@++;]5_d:B+\,DK;a>c0N5[PYP=
5\c]P,48[D,BfYU@:+V>+_eQ)Jc4g^[HR:>?\:d-gaeGFa\G[T(E7=Ka.O.8/ZIO
)MfJc5Ib?=_Z.-#>4R7/7,>]4;&S_Y@R=I)64RC7\@J]/.>1=/SdNK8a6P.TWWKL
[;W3dD^eTF8\C8)]@2@&9gB+fARSAbOG>a<KDa-<[Q)).e8R7+1EBHF+e3H7CTV+
(d)G?FL(.\f[UCeBDUXC89M;]6C,032KT<TMU^>Qc-,gY7S/G7CZ2C:fCVOX,8N7
6bK=#G^9CGeZ4B0-=7Q:BRDQcTdAW)AZ0TQPD5HNJ6<JYFU8Cf3)XHT8]76&Oa9O
OW,+19)(a\0EX+?W:K_[<b7G)GZg7Y?\^c,WMb,TW=>]_HB3:f15Qceg5:Y5ce3G
K23H;U/[?O#>U,GZLa#9APCN\?TN]T#^X(#PRgLb3RZ9Y#RN71RcPG04/1L&Y-fN
g[)9/ScdOLO)9+F5A33eSE:a50?J65R[3N#EOQEB4R]A?\51cB]5f0J63.WG;.0J
>RY0ZQc(1^)Sca#8WBe+5@,S-D_\Q.H;-+103OY>]XZRQT[TUSRd/Y@JE?O7)E-B
VT(SXQJ20.V7F<7C>fgIfaaI\J.c4=TU(,_MTgOgW1YU<C90&4?KIHcV8OVGHY1W
UZa4YY]M8McLaf[0E#_-=A+0S73;[L6b+/[G@?@?_B)Bc-12UKLQLI\07J2[4R&_
gN4F4,Og;D^RdgFg]#8=K&(G_MBJ;5NIWH/b@[;BQM#1A?>XNG[W9RdYI[YDK]cD
8]7ZSX&\BX+4QOY7VK(7W=ET9g#?],G^Wg1;UKQI#a2A;b=Q;#3.;,S7PcMfI91T
BDf\;I.Wg2Q/dSNY,=4O8-+_X8J<O9REWB]?DgTPXJ=D=M+C:NNb3N-G1L^WZDQC
3,R@Zd\Fg8-WcG9KfUN3e;bV,W&J;Pf(Z:RS/ba7:H3((OTB\\^gJ8)H&:#IE+>J
^0L25A67A+fOM8CMFOIdgDXX1.=I(F=W#7)9QedcGc,KXbXR6McK,D62?>7E#Qb(
M>[MCgK3N/D<<b2;<c#&VIWP7SR=[N^+bVS5c5==UQcO@;LfJ>6:WQD#@f1D0=J?
+\-)2+)#BBEZa(K#.<N\(Y-b]&@^_9NOc#&eR-g,E9f(Je8/\+HEE=C_B5fST3J(
\34_P0=:-aP[6f;4>J?<A/e[bI#AIHXfMdIAcFMOCdYET?,4VF&6]_-=DXBK=5M.
4RJX?)0WKNO?,(\+NbeJ^5bTUM?\aB:&:2>]5B]BW<B2@EK2I\MQ[_+3/)Y,ZR\]
<5PdSZffM3,+WYP[0:Hcf?J5&30[;BDe=YLVPd=b/6ZXggY:cR>=-IX9XC@,?,)&
92G,,a,8MYR>=\b=INZe-V2H0SH8\.WW;2VN^.b\[2,U#E+^YBX647.(VPQ3]D4K
/SI/)JCQ9fSDR7,D,)OE8@9Y1:6@30JIf5S+dgB\&M(&SGIgV:PVX/)^HE22N#&[
d@EaRe[gI\91,WPX70@@RXdA9VEe_./]2+QNCNT2+)7LHRbD2W->f>K:c=PT:aS1
P:Ha9;@M=f]0J0#IfDFB<YG5d9_Y01QZ,<:--/S\c-3XLMY8bGPY^+:/\JM4A]g)
JKDI+c]V\5HUVAXaTgf1SX.gQ<2e\Ae-IL26=8CG7[L0;,^f=>[R96<[XgX/\QL/
:g?OTA3]b7,7:ZU56>L]QXN@YRE+=Y?_.(1#0XGPGT;M\T\CeDJ_QUHD&^Z#-;11
:5I2(f(<AV+M491-<:+(N3+dR284N1XAKaIB;4=0>:a+.-f]L=egI@)cU;G4c\eW
PP&H0/S84<Df+Y^\>L1DH&04A@A]1b?O(86/XTcfYN[5MX1/QD0T4gJCQZ(T9,D3
.XG[>&dfG619<c7A1-,L_#9W8Q>[N<LU)6<,+7@=VJTLaNFJWN_CU+E^2:0,c?A?
;/WNKfNAD61_VVV5a/Q:Z>=WcaRg2R8.CJ,<JZgQ4@@#F2K:IXKGg+),P,4fL8(N
QBfZK<MdQ,@4G480T=TKCbC>M<Y<<VATK#2?)Y[]R-)8cE8L018WV3.2I@F4LU<P
3V?]ME_L_-E/U9>-I73SE>Nb]BfTMFcgH<L[<Q>SdMF<d^S_.DU3=IfFMZ/;dHS0
U++e-Eb5W3-\:HHe[]544:f&1Ud:9WMTC9HTA-G?a2d^4#W)W0a@&>;V:QRd0ZI6
5P3Q#P5BO+_OfC9f3)@DPg@^]2d(+UCGHORQ(4QJfJS?BB842,0VQJ>N3f@T-4KS
;TQ49\MeK&6bcVK_R\d/H(/2^L\fI.OYG=d__eD/;+.42#b_>QLUYFRBGX>933];
\)6P)4=^0\Y6@#;c9d8UXL<aICgL<F9^[G8NGcIfIc0&gUW/D)L8G92aN^@@BNB+
I]D[Jc_,>><BETQVMV5daXM5;HUDe]O-J,WH#9Pd@O9APP5JYg>2FERWRb=13M0S
Z5_Q=>4O0,WE6,L@DC/4=@(1&\W1A@8g0eW@U10gV(14WZ(\/OEC>FS_1[Sa:E9g
QHE2B4)E8O(UI6.NEa[Db75b-<,#N]TK[8W3V0+?M<dG9M&c^c68_A9L-=8<LL0#
:^#F4#^Yf/.?0\g>:A,:E?0/,QC]1-H@X[DU#Z(@gC.GD0<;C\5SfXCM\O5+V2\I
H6XECZJ@QbD<=&FD>UIG\PEID<]+bf^bN#<BRC,^S^6W9Y?1-\VULCdMe&3Z9g.G
BJedCFIRaTfe+4=^VH8A-(?)U(JJBE9/LQ<<+d#@#YZ,-5;:2PP5X0aQDG\R=+A/
6Q(O&>#WKB/S,Dd)+SS#U45P+)>)D,-@-R;f6-Y:Ja0PXVeVQ+gT>f)gLI1cIMCa
I9:dR,:)Qfd3gIX=>>4>7SMFOf@G5dKC/M#NfC&.6V^TAE]()HN-7K].gNe+?1=^
G].(H#bO4d_Z(<4&WSe\g42V<L/RMAd]0CPAdODF;GIWFcCGP>]aBD9L\)2@K#NR
_MOSQ15Y?I#cg2c02([:B+f86]B6P4e-)bZBD8ZR+V/W]4,Q)H0@(Bd6@aaKD;[X
9/<YSB.ACJ+[;Ld?.\#446bKYN7JVMCN/?VC4A9YT,,R1E.g=T5d,Gc3E9.0T2Z/
VC38e=acfLEgGfWTfO]XLYL4:bO8PaEKU@X(W\W9c0NEfK):,O7R)<-_f+RN.J<N
06[66<Jbe)dLBV##QRU+N7QYF.O=?P](XZ;4Tg9a#(<RC.L<;@+WTHRR2+UBTJ@1
W6&+6MD,(PW0S4N00U]\+OYLS__7,X]+)CQBd<[?JNRHO\&Rg+TRD&c>=X[:Ha-^
U@KdXW)J^<3\+SeP>7C_/G,ACTeZbF+WSe^TC2U,aV.3RfM7>;56QV;PK.8Z34GE
fG&W>6@JGC12\N17(]_8O3/b;_(\Uf:?E^f<Da8Lag=P@1;d\Q7UG?)K?RNE/+WG
(6-5:B#8f_@SMUeZR9I:Pg_.H+T<0a)FfAfFK0L1EU,C9M,.&W.d\C]KK\]3=+ZD
YJPP[5SfgPd(LM8/152F_I=G-65^5S4eBF#[9H(eF_<+5E4[LJB@2F4W<B>.XeM;
DNcGdKS[gI@9,V0K?&-JQH[H&6Se1^3X.5bABeCJ)K_]O7TDX:@6KgR4B191_#EM
UAY/70/4_OH8C_3GCU/7)AXBU3?gg]LI#JY6M<\:UCYEQS1(Q]/(<<F)NEE,>W>@
1f.eWI6YQBUH?9.:5OA\^U_ZJECZZS0UXXHZ((-bN>8VG,F&?>WE7e446;-(d@9R
R7YGH_YAe3VA?:[>I]ICV>6YT].S_FWIb;SS,+@#>6^SJ-;WVLR#L(+F,b)V+;\@
G8cO)L49eBV9NY_IUCJLCEd,f1#(a;(AVEK[&b12OgYacc^Z#;,75gX3FaJ@H(Q8
VW\,AMW6Nd7#cI<d:ED6-N&P+@F1D=+PP27IA)8EWM4+-4M5X,(X04eaOH+ecd3?
E<<L&515V[<N.DF1-U=DaI13I;OgZ::KH<c/A+INYJR:ae5g7FFdZ5);YR+b3^<1
>:/VHOVZ7L\[#/7KAd>])YdB]5V;d_NOe^_DU/X4afcZE>:eAT1(.J0<K#CAbe[a
KQDW^g1VWMMb7I?DcB^)7<C()d5FT?=>W1?BcO+7GF;Pf=DHJ.PMX5/43INHN2b0
+)Ld1fI/_V3I_Q[?(/aV32/8)6(D2A.+[?,gJ?@;F1R,6?HA;/R@F4DM3@P47<-&
&b/bCNQdS;0=]-CQHNF(Y.#B#R,/)E-2F-ZJ5#P9KI72QQfA\+g9A/3U\\EN]TX_
^FU&UMO<X/9d^fJ\M8S2I1P1<C(f8,_-/g(Y#b:+F1^LIgBaY/X,.@,5=SH7NA]Q
Y)SGM3E[b@_0G=d8<DS#0H2G(SKG:De/9gKf=fAJ>E^AW6#cSb7Qb_MD51]/N>ag
B55dP:Gb3:\-LaJ?:Nd#H=bRaJVQYQ5022J&@I:gLHC=FL9;1e=0fMN8?5,1Zb(.
F@54ZRCI^4Qcc176#11+:S\OHNS,b]a]&.Ya)DYX?.85S#d+D3L6[<R=UY^&=1W-
C]/.;/^3d_JG[V?M\J8#J(TZgNHZ+Q5;-O:Z=5b-@D^QNeGUHHU\b?69Wb7652:&
U&JZ>J@RV42A8X,QU=]F[b#V9TR3dMb^-a:7(:gA8-.U5&J8VfGWDLbcYNQ75XbU
==2@^(Vg9&fEd9^3+1VT2#cZWd[YU[d9;TRBW:@/7XKc#cU-)C7=9=H>bgXJVEIb
&>cI8/gfB9#ZZK8N&b/>)7W)91Z?TJb+/[J3:#0;/?W()S1F&<\;1EE<.@+aFfG4
[>a5:PP)J9L:250-_@<B3MTFA6fI_GH9#R->_#[D1Hc6RDZ/,R(65-5X@b;A4S2P
^Z,+/H9gLY4c3)F+=[6fV\OZ5&O?_L@W\Z]X\-OB(C]?-YR&U(SR;>[;F?@7[N\T
\AZDIL5UI\_[>C[>;YF)0E^KJKSR>/599GBG3\3]#c<W?a2EWUEIM8CA-)e8aS:6
d(C-2U(8./+ZY1V,94+cP)U8FbC5gWZ;>><#OD&P]#=)A?+[bcS)THdQTR>)#4=R
=I1ab0QLQJ>E-]9T??EAI0(Z@WD->gCN_INHO\3\gKg6Tea]^Z9AU;cBKN)0dc&2
f(&^]Kb[6E\5@NLf+I^CO5L2&-=Cd/@?gFUZG6I(#0[EGV9U()WZY7#:)0Tb-Q;B
PO+F;IPB7Dd6\Cb]=bI?CUA_-RJ-DPeLLe+V^2UFG6Z1eK:<_VMQZ@LKDFe+#?WP
8,EEbZ(AIM58+OL@--_0PR/6/E:LE#J1\+Sd@TA88IM7=HQ>@PX=H#\CeZbMF82=
RUQdFb+@:=[F<?;d)(4F=LdZ3AY_4[1V0UZ[\F3623c88=c)&?bP<WVaVZFB_^\O
M63V5LNX)4UM^EH#)fa)ZC:\MaY;=N(4^D#F-;EW?)Sd\&DNcOcGEAF/OW\-ga>.
+c8;F+:A0-a=5(.2+7da-.D;9&d1Hd8_b(8A-XD]-^H&55.D<0+15LSg,T5G^56M
QfMKOO,TaaBKH-c#/cJR3YS1/>;+7CIM7@7XC7(,BLc\6,)1FFUgObOBa)FEb&\6
aP:YB_?,OG--8W3?BF8LR)_&E&BBFMIW)R3,f@6.@UPd0LXDT?HbfGdZ>?H_&^R^
9b[fX)?F0g0458+1N<eea>NV\B=9[(XDP3,_=A+Z:aKD?TedA/^b.GF<c(TD(UM5
^?X>8[^PGRJSMY3E,dM=eDLC-DEf,R4^047WSSI#+Ed+bDdE@0Sg:0T\2<J5UgKX
[6:15R0>gM,T\?;1W#]<_6K;-,OTT0[Bg#NbEe8P+@=&5;0N\TO6A>0eP[S4d.J4
C(>H4G,)0fG3O+=MF,QR^KQ)])GF2WC09[9^3T40/;X#>E8=NZMgdgg:9f601b8T
PW@SMD>5L[#/+TD<I\HK5EPO>;2Eag_(/-7B&9-AM_9:c?ADM2[@T(NXX3==4VM+
a@.H30Ra6&P7AW&M3eYO@]R;DS3Yg8]JD@C/-++1IT6X7a<:6WMRFVgD<D<;dSZ(
a=7b&CIS)V\1aNV;5A;07Z)C4+EQbb0F3\J2OIG4@BE=4@@L3]PD&LaW)gYD48NV
^+&FUZB<I@4NPJ#,RYQW:FWYX0EdW&TN3dZ>18>OG_:-9_IW;@SO/QAS^(E5TYU)
)dM+eIJV_G8VX.<4#31PG-.<V#CVd0FNd\e\1#K?M/YU9[,bZMM@)P)]C19E&g=9
3@E.=c7QG&<3/9Q@Tb=4XJ2@\a=aM>B]1)H89b^Bd,<#>Y@145<[L+aJeaN0d&f/
V[bHe0-(^X]NW)c_XS;6F4,37gI-1JMC8a.#K(R^[ZKST^TGg\^2/@Zd7#9Y/W[G
Za>P6KLN6=9AW[<BK^4H&R@dXcNNW(JbSX,\#a>XP^9T\D_Rf<PdV+Gc7-[H&Z,b
Ae=d/FUQ35Tbf[1P_cG9\1CD+X0H3UQXK:Q-e:Z13C/EHP<QS6>I3&=5^8KWMA3b
_^E2eTN@-<-6dI_);<,g-d1G22#d#>1a:._\L0eO&b&O+E=AR:7.Z9P-?MM/E[1<
fKP&:MFTCQBSUQTgF.HM>dV=V^3fP6&X(G)(@/+,5_OQ/G2J5QJ0TYf->UP1a+I_
LLgZM0D&QR^GM?X(V\.O(@Z;9Z2^bDc9^9I.3^aNYXUG=&a)fKHA(&d(fOWaE7W.
8UL7,7863FSD2:>0?=8@V/Q@eG3PH;N.4-0BT.c>fa/VR(Z?G(d\BU3GeVL0CgYc
1U).55]+[S\Uc42f\>5RO):>?&&3Z?5F86+VWT?R^A4+835CC=g5G9JgJ=YU6ETF
@FH4=K6E66gMFab58&J4IXfRGV#9E^dTfYSF9-&B8VMf46>.-,8[#5\\YR_EY;PV
#:g5]ZO^>c;&E_SB-<^;0#Y,+QgdECH]I/ETK41CB^QGHM>,LJUV0Z#FJK0Z+\-M
9B_.AWAbaI,>2[QHO_:0fd7Pf^M/)/8Oa](,JO-,2dINRIC2[#f^AIdTM)?N5ZNT
4&gdLM84VO72;>VX#ZAP/FB>1GP<=?.Z^H9Oe5K,5\6V<V=PNA7&dW82c61_@@dO
.3.\IT&JS8^L/>N8=2RR/+Y0#2Og6Vag83.8^?;,UBX4BL]LTE_<9(T#eaQ<U=QD
Kc@\H7)DB2Jb[g#e#Hb=U#]2T()G0+1J;d5HYM[,g^b<1a6:bPNZZVIJB>;TgFU3
=CTK&0)K3Ag61^c/a]eeF/.M/6a4:U:.^/INLL,)[(7JK<(aSV#WP,G-Z/J+]7V4
+((8gbG@IP,0d>1/-8V[Rb/4OG99EJa/]g89Re(7K:L01@M1NgCS75[JA(X=NZ.@
gB9X;5LLg7f8.ReA-WEO]fKFda9)=dS/=0)#G9T,X7?c@#099V(8S7E+N8W?c)TI
[[JdbO(5;IE&L(fKWeWc\V6I:8;N<>ZPLVY@JY8XHf3+/fD.R3A2GXI<<MT:X7A@
1e-\d+)+03)SHKATP>Y2UDZBCA8/\]))GZ]CPN>XH[8\aG2g2:VY.>X?@2>SE4G6
S2aN>T[?LME8R]GE_]b]F:fc@XL.228L0N=,Sf]5F5ND^1,7=P+N^TD[9>f<&^N#
WYM].N:?B[,VF2N/B)EVP/[:4UaEe]I6LZTY7aZJDY.+D&RcUPO8_5RZ6f?K9-([
9aG@E[KRc9T&-(:=R.W=2GT+-/^]T7ON?=R@S--WOK@.WN3Td8JLgU)cH:>4.J\.
JX54>\I5B2:Z,/+=59;5aF5SN,(=WFHR;7-),-GA/:0.FT#d9RC@\g<W,@SD0N/L
TUQI8fG2WDA@K+\=Jf#ZD,-IK@#F(^D/RG>:fa2&2A8S:.FNRgeGI53G?E<QJP:]
dR@]]VC5O\gbYS3@#6TgW<BW0I3F_<?b]>NZ]S.cN?L/?bAB&;JGDLSX_[7FgRa3
-R.ZVfKe7L@40AR\M+(6gOJQXD7fEA82^6e-C0@CDMX==B/c/4^0g-53JV2A.@KX
M<:>3Z&W,37H]RPN@<?X9Be_##80INZDPa,bfDLA<A8FJ:.BX9B@?]CM48WEe<g3
]UDB1:Y-[1)@05T0M)63O(.OEHZ8a7O_-.0_YX7#W,IP,P.T=I[H\87\^\-a_#9Y
LLT#,PO0YC;VA/\Z1_Rb##2GaW&)<J<?GU0<IH8TG/BcaK>XE#7=^IVI_H8_a^U2
C4MH^;KZTa&]WWg=<U8LX1OVTMQH)S:(H(\IS01^gP-_CAR/fCcW=.)],\E.LJ+<
9B3g\bCbQa,-(Y],.<ZPGFXOQ_FD0_5Z[WH#\)SG4bB;@7-=,-+)4LQ--<2ecec]
D<7GD4<NR?\-4GDT8@5.5M0H3ebV@,D(:gGf=IZ(8KQ@=K:P^5VYTg<0U,5ZE679
S7TZ0<PMQI.O8&QHLH04H\(MQ#=HTD1(+,E]WMC8FS,1KdY2gA6c&/3FLB]&#fbR
[85b#=7:eK&Bb2eeF6We?+L=gUIWVA87Lb2J,ZbFe/SHI)D#]V:5L<FDJF3)BC+1
IRg@N>:EMA>6R#N59XV.3T3Z>c(-;>SL:R/0#[ZRFXD_?Z0HbT:c1cUW&<XO?4D?
bPW[NG@5)0cFJM#[e97L@R.I=FO?9>/Y2Lc9dDHg6CIc[)\XA1WB(=a0@K)S@Bc=
Y#eQO]A=^UdFbGVMAUa3KXWH\7#Jde8#caX0,J2+BWJ..X\6RPSfJB46Q6VK._8c
DbC>_^B,085af<\JC0SORS?HL^V8JXYe[4,#9g-XaBDXMOYfQD0FH2[JTeT;MX1P
4J9bfCQ_R3F^G-PQACZZX+52^?GL</85@#OX@e4_FAc1^0SDA7H#b6&1ca<A/6I@
F7dP;=.9a6G/T2S\f_^3._&M-\Q&1f/@@&38P(44-3ZPN9bK694)QAE]LXcLcI#S
06KCOBHfaZU[JJ;Q&D&(Uc,V4NR]MD->WfDG/IOLb\RTdKM=P.+UMfD?QU1OFCFa
9-4cR2&H;@&0-70g>cS1Ndd_b4(?&,gBT/\HK3I_gb2-+=EZIFZ;4.59::A]R0UK
G>RK=JKBGB\1Z#+2J.7KaH;O+T89fM;\<a+VdL[d#Kc=4(Q)PE>HcL=P4)T_47?=
L+<\4\<JDZ[M+gb715,\EXCPJ;9+LeM).JgGdI28cX^.Y-N.KgcGSO^DH\3QQ^01
>&a^IHf>B_O8P=<BfLQSdWJ6+B2AUG>9_b.TSC&>;CEA-7(@GD1<.gd5W+&6S.B\
1H?VOZE_RdDf2;O,TEI0JK;W090]X;3R[TcV=YQ&M&2,GLYG?E>OBD-3K5(A.9BP
b;8Xc.]5\<KaX.>WQ;PX53=Xe1dWP?J?.:Mb6Le[:P4ZLY@A:\/>.\=BRMGC3_BX
=0S<f3Z:K#gXJ\(N\KOWdN@W8HCb0K\D6GD.\#;d#]2C2HddX(:H9eSR<E1ZF4Cg
-2dP:3VK<b+=F84_J[QF)<Q=V5&8E,;DW&b(2JVJ/TSH_KGG1d2=[c,;U-0fYH/b
;6(Od477/g==g?aSCM7XN+6W;NSY0QB_&A,.L4I2_4.<CWdF16bAeRB>Zg3W=EL?
WW46E@_#C+?Da136#EUCK-H95W205W7&WNT//BA5c9L?(-2a1DW6EVAN7KZB.dOJ
MKNb.IM?cI^,VE:7B=]R>3VK&EC=7/dg5,=25HFC,Bf.<_dVcA=<5._2(e>&b5Y7
eH5ULYZe5_+1?ZZE<5-A&3-+(;-7NRbIe<C((&EPO#NQO)<\5<HE/400P20XD?X\
9P(_cg-Mf>,.,C0Ja1GK__M5O2eG=]VJB8_/)&<gH/,;eN2<PaVQQcY72e^UaPI7
c[YcG;E^0;2W;H^SFIb^cDgL.:MA:;2+UV)<S_QdBR+@3H4DFC\U7XBA:.:W^(AZ
6I@#).5(A;9a:=eC8bMJXH\N+^O-N+_WfMS_<;61_,APJ5B?OMa_f+e_P2@DMS?=
N:#TUSOO[[5=f^73>>(1ZK,PCAL5537=6F3A)J0;VCY;/KUM+RIAZ]<IP:,NC84E
8Y+1@9RQgVK&Cf_c4?^^-5gK9?J[a1+218b+Q^b:a.Gc7YL21?KQ(a;]3AWQQJec
<AQL-^->=3MOQY][3NK\CD+WSL3VMdN:HAN8TBY[B>VF=QL=-@]4:;6H?R0K_F9R
H1(bA2Gg1^d1T<McK29?77_FeR=IeI<W/;+PI+d_.d\^;8d;_)4,DF27XH8N_=K?
>YTef8Q.)f.JBM^EE/FF0c3TdDSb73a#&1]7AS>D]]aOd>]5/.@:XM5?a2YW3.)A
^?Z3g+Y5);RUcf15>F2=f8[&O[Q&K7)FVJ?cN].^YWBR^?LD<_6-/3YH2>@+Fb4\
^Uf>WT.:IA7_3FJUBWa?QCJ_C[b36Eb6^DNeVJ\06\P]/.eQ4.X-+0M:@:+P7=HE
bg/1cWN@:RA15QHf4IV,.ZVQ(d6UFP^aP-E6)Q[SDF)W->PceaCZ&#7dTZ^2E/a(
+K[V84<7)L@?=V\XbFC5C)MV;AZ=2J03>]XETJ4G_Q)[9JGZ0P;C2de;3>?HA-[Q
+G\L/EQA@-:dGI,];3+4:TRWIa4^Lc^(SA4K\0XU>6a;E+4ZJ@74-GgYL1IXISU5
Fa,HJUI@)1+2]Y[;,V/1UaG?3G,(V?9fNAR=1fD?JOLJVY@=<3J1Ug>:FaU<?^6;
4AeGMG29XR-&@EA.7C<D;SF-\>8B5-AEK^TJ]Mb8::deSQT2g1R0g::C\aYX8[d(
10QK)J<2JJ/OZ^&VW,C:<bQ/>&Qf\\CDg1#1A@,,0:IQN\2Z1H/(^-1d@cL8UYNC
KOePTaf,3];CGA?B&d+>E^C\_,#Q;X6JV;7]]L=QE.]BCC&4HW)[1E:.e9QObT[4
^=7K#gGBaN]b^-W4eA2=GEb0gTKf+AVKNg/MPfSX,fe;8<+bR.9K=eeI6Xc8B202
MAZ?438]0dCQSCIQ-LZ@[KcO.Ba?3OKT-dcX\@g<2.HW5\_C6-TUH?Dc82,Z=62+
/T#IME5f_d8MF>MD,U/0(.F2>,JCIe[2?4B1EDS^J9?<?]@1_9<MOZ2/P5&G\]@6
O@NDO.R8G2492Ag0RVWIIP3aWcU\(=_B1c#R8IZ@FV88&MN,3-_D?W#M@IM2>LFc
gaPgO_HDQ+=(Zdb)C?f-a(e:<D4I56P-0&>WADbbSX]7E1\:Z(2gRURR>&8(cX+[
&8GXR_cdJ>:P][4@>NYa]8:ICK<<g20Z-GMG^2,N9.Y]YbL3b4ET.N(=4557.0eZ
WJ(7:-Q9@#7#,:d]T@]MXM\=4da1_122_A5I_#YLEL6<4W.RF2_H)H1[UKE1F^5g
bg7V+W8^MQR<;YH/H7=T_,+b#@LC@>B+V_D)?[MK8VS;K9YSDQO8I6-U6S9;@,@#
-_)E7a91f^_P)Hc9_K64G)X5DT3^E96OAf[Y_<;B@MDOD#(/,@7+<-c/:&M5AGKF
5+E6Me9^V+J,1HPdDWQRHUSEILNS6XdGc.3UgcG-M/5C1E/J_-T#;0ZVUaTg#g=3
OJ([BP5KP3I:&BH_6d&2I.acN7aFa@-+S+4e929Q;P_U[>[@\>MAa45Y.F[Q09e7
];5=LL&+9?Z^V0/.3\bMQ@7TGgRbAf4H(?FdQ\;<U<(Kf&F7;[&2;gf@.G1BAR(g
=JX(:J;^P8@I7X:E[/_Fb0QC020EGCCN20fVNI<ON[]O_JLe;Z_3##0&;:6ME=Vf
T[(\J=__BJGc^80N7:>/8;/,Q#=RZ>aZB#-D;8S-R/[?HA:Ff-(-^bX#=_TdLKa#
5U,_&KWONgMd;ZXcR8-1:2J]RW4.;P2EG8(IeXJPeX<N]Pa7V\O^PddYd,P3[<9I
Y@c9c,O@F>^W<8CGLG3^ZMbW1N9H<>NP^+a\HLPO;<#Y6b@&^#=[&HdM+GI(H[_Z
Qc#Z(L9XF2U1=JYdM>d(O3K13^0_M+:+S0cH)3HA>0O(-Wf8)Je<KK?6JFFfDM>C
S/\&L?@GZ>^gV.^]<);?-?Ab1Y-bYaBH-;#JT+cB0MS-<Nb382+_+L<\N=J)AR7(
4dHMM6K:6-Wbe88OE[)G_6X\ZF/25I)fFG)/&LR_f8d96N#LUV[@aDGBQ2_CZ8cC
@eVKL/ZQ5P)1B#4;<:&&24LMC5B,03GaUUU6Z:f5XS9..H:8Q=:G[NSOP4RD@OX(
1W\g4OH,^)?BH_C5O=HfQ7Fc\K.2]R[_=W>dE&STRW0XX.F6ZfI0.(H4:8/dg=^8
L_J/Fd4#;g_O)^e[?/@c5OH6L]Lb7=REKOO3e<8.VC+Z3G,a/5U9Q_^GO5f)G=7W
]CcPHZ3F9L7cMTP9_.22Ua1[aaYX8gFY5)<</eJNRGHVYGOG++T:](^WE(7,MFb;
YD1UB6#PMZ7:=ODS#,?:X7#&7CH,MR--Y9L4DPC9KMLD]XK>G](,HI>Nb=<D>c?/
de0[]I]R/dJG&eK&d\EXLU>HK)=50R:E;3-?A1_,2@H>N&P8(>Je:AUJe^3LS6TW
=5R:OK-WG[fD[bPQOgT@+a7LU5N>6W1\YOb9^/AT68VUBF(BB#F&+A\A2/^MK=@Y
^U76(]@B:A/SBZM<L]C?-1VN^_Kf4fSa;TDH/1/6RRGTgV)-B>MA;)BF.+OM?>^M
W?^1C;A_\2[P><0gZ;P0MSYJ=,2W_Tb8FP-@00:E?4]Q[Qf(R5>RcA\?^P8<U=DZ
MHIVg)(+LXGXG3J\W-R>52+9(5(9DR&#>7XG;N&/XLaPFf44&(4V)-5aaV-[J(#[
C5]?.<(#B,B17-/1Sa4e/#-7cB[J+TdK2(F7ZgQ3.N:]34?L],e,MAfCW>Kb));:
((/5TL#aJ3[O)MD8TP5+.U^Pd5d&8=21+,\[+78dADL#<K,gd/+NFN3]BV5fIB&Y
3e;T#2@,W>\+R)YcX[=d_EBa_U?39Y_4C6N(5:cXQ?E52+U_O;1ZBGW+HP83cgBD
UM0_EZ9EI0)/;29:D\CHg)[X,)6EKRI,Y+?+UO<WVeg[GZ1?BIQ\(EgB@[b-+0S#
c3/:dLb(UT==gGS/AE+G#7A146T25[<=ULNT(JGJaD.=KY?J+E3KI?=GCU:d@>2b
4\8385Z1ZePX\[a8dA)ccS6a57LUaV74/;gMbO\.TN33SNDRM.8>eg=_YZ=2^B]8
)<e),>fE^UVSg:7X;44;bFB\#)V4,-5Q=3,2N+O#(RUMTH?I&R[1TE.bUb)H@FbP
N^J?H^[LK],XQ;H0//dL7D,/9V=-HNBO=62&\?Pa#-KH6/_(MVUgUB/W\)>H8+?I
-g&;(CK3fa9>]H4?K[42Q1d<VJgbP=6P_A.3=QH<6/=RcaX)0RW]\(V,CNBLJ^^Q
70WPVg:36YEX98NJX4R4>]:@_@@15Hc6K-d4[2W^<>\OeFMcV?70IbYKG)5C4fMJ
>&dfDf(&)M+I0[6\&g+Z\H\7Id5I2J.0&E/@WQA-<U5-ZNd94b][a)45g>B,JZ=8
#Q1J_?XR.(O7-LZ#b1R.78&L+CfAB2e<=f-)b>KZQIW8)N8-f^;266G3TPC<a@:5
f:&E^#^5Jf]^]22@0UISUcN:B_R^NZBdXaF#S+DQd76ANf8J<EgR?1,gAOX0/c)7
?K&P][,&K1,KdINJ=^c7:\?Hfd:<FdJD-SHPJ;+/PA8SOTLTHZJ48ge-)D;UO;UM
5##<,RZTbHW:(E/[4M^.ZZ;UFY0@<MLd(-@cT\EF##Ea][5?eSM/gIZT8RQdD,L;
UOZe(?d07=1XG9O-f,OYW1>CPd9_:KQZ[BC_T#UCef8Q+P2QbeU7Fg9Gb?Z.NYVO
U;JV/BJ<_I,56@^OP#XBGcB4LO?JeD2bB7/40&gZTWD>,6(;&OS^4NW//L\3B0&=
_-GLLLG=CTAY\W).b(^RL]DQ&aDYF(&Y:,M@;,4\8+0NgJ)Y](UgOU8KP?S)(X,D
>fMAB)P?L7)SYL4eCT\DUI:39=WS?U/_MM7M-A/(857DD5JZ\_Ng[+;d?AA\(0S+
U>V5;KV,ag>JKJ3Z33+/PU621FSFC:C<4Kf/:N0EG^b5UXBX#H4I:J\NZ5):6\cb
]TKV0RAfU_g]\aR>(@&N>VBQ?7U2N-\^M.]<+#-OAZTg@)?-SP7FED3OV&SaU[AQ
<GD90<-ZU.>aG;(D>I(<]=P\>:H.4JN64WV,bU\Q.8^L#E_OQDE03TM-gMK\[324
]WO?:\;=2UY68&gFC9H4;a;01TOMN?<g#9<\B^A@#4=VNgO?<899A&c8G8ab8bXV
(P::gd>Q\KZ+[K:X)>bcSFJHeJ#M?bI8_eg(202UY+(CI=+).+\b9PR6I#aW56Kf
;[>5:OCU,/G]I5X,4g\WfcN=..=+_BUE&NgM0WG[eWaY0EGKCM1);L^48Y+DaS&:
633LTRH/1/XV7Rf^K:V_AT06RIYYY2J<;ILK-K^dY2(2#g+fA4BGHQ9^=NQ@d>Ag
Z[UNEaW0.;V@.8KDOP42\)D>0Q+)9WZZ>R]S&:7#YCC<UF<C<0GXH\+ASU=61&H9
+T@]O_6=7gC(B(U[bP@85GHI[dYA_g0QW7^?ZTJU>gF]Y_UOd#&TZK49D9XdDLbL
O2BX2Lc7S)/YT^84.dJ,E&WBBE_WO.f]P)U/S>>>-Ma;POad;-a.7^<;\V4#;,dJ
BDAA_e<f)CLRK(1-XQ73JE2>(e#:Q(;@WJDJU#&_V/HC[dTO>>0+YFB@0DE9aVUc
G_D8W#Df0]eUA8a7#\g1438\;_gf7?>&/[=a(.]&_?=6[U6COGR^(T=,O/ZOCgU<
@=>4\MRMRK#/[MFRReSV?@URG:YBYGA0:FNNZWXPcKB8Lb3/V;(e,3F9W)#&&.[5
-[D@SMAaX@J;<#/M30<UA-b8c6#[FMM_H[J5Zc_e0GNf[XC.T\@<_R<(>ad=S&V/
[+W=/;[G[U(\G19P7CIA&e[__VYHDbBEX^20TM68Wa,eRX&g/+96aGKJfUFHW:]B
]-D[1VT>9_RT8S#gC.H)@cFAZFZdGP+B;_XOW5PHCHgYTUHJKTM-2;+gZ15^8,9L
-NY4,2\R<)7M7:JH8POQRU\HD/?dC&1FJfdcb6?43T>>_O\V0&fT-HK1+7::Pa=c
-KPZIG1UA<gbRNUE=&5;Y<_Md+6QR7OAZ?OL+7AK,(GDc0(&:;N\IN+]<3Dc++U5
0e10X[U.?EE.dR9>S-8bXeT91b5MP=F[>\+)I538H6Qa8P\?.\N+\G&3FCVPcB=4
K>THccLf9E]8>dQ6)=_+&99eLUF&&?UQZ2QLPSTdK#KD@_H1f]b.(>C^/^UY@/=]
c^<.Z[B4aeEW^9CJP67>X37#BE8G4<77?F_BC+2W4RRUAd>HWK6.G)]Z?;>IG<Gf
3U1c@H>WbcCL>H;MHS&UL,0/(ZU-YVHH@^&DT/]J17JIV.PAT//XCMAM._XJGJ@1
(QZWcM/aOgQa.0+25edfg8@.WU:[X<R[@.Q\8^bg2^-PA(4UIE99AR_)99QN>#W7
SHQd;-GYeLA>M@:FX>deD;P@M(L(EJ#X8-?;])b3dE\7gV>[JO+<X8+4)OW<VX4-
#W3_,BS])I@XSZd0-WHB)F9cCJE077<bdP,U_LH^AVH-4.O5KJ3YNL;]##VELc.-
BX8V7S:2IU@+QM8)/+:?#S1S-S:5N;G4;GT#[<NW.1C,e<B\TT7Y;>O<GX4K0V,a
.CP0BPQ;GZ_P@TFG@+&+\,YBZK\FXb&2,^9U7BgS\>KMdP])^5GA&7b.bSXUG(;9
U?2V^\a&09.S)K+aRaVGO+#e(ZWQWP]#O[aIY-(&#(e3=BI(-9&[1IB8?U?H,VME
XBSQ5>0=.HA.g8IZeRN^_>bccUb\MXED_g7:NNaO5)[MgNDCA.gVH\@ZUGKEKdS(
9[L\A\R2>8Qe:I_G),3RaV^_AF+H6,OV:da1F=f3(E#.3FD&B:^9\9[Q?GM;HD>E
D.bIUH2OC3g^9;[Z22GA-U=\Y)=.bKe[A6]DQbO9T[6@4MTGE56M.K-LaYKZcS/L
bN.5Ab(]/WIL:@RdNV@.6O0AGP2J/2I1cO)\+\\:T-Q[_fF8W-XGgDc9@ZMFU?I8
1V_[MN=C9gICdN9gF<>d,-V1/3LLJM<,g][0O1:X0.&RD<T,/,:2&9+5V21]<^P3
/O[dJ0ZT;=2WGE?b3F1#WF<E5eBAJ1WG.Pf3a_@Z9a,.GaCf06_#bRE?Y^6KfBO<
IOMS=/G756_.YTX=PDXVeVed;5\<--e8R^g>=C;BJH(&^4K6:0I<TJB,f#/AFO([
=7<L@D]eA[_R39f90CEBJ(L8B(U<0YV^+a3V@=)fH2aBQa:OM[FG)U^XQTJ\_\8C
-f\a\]W&)K2-G(bSQK3=-6PdN:,d11_.15YI6R<a0SRLW:P^D8D=6[K)BaBQ@J4d
46F#Ueb?4LKe/=1ZGY9e^_;D\5F>^Ma)[#0:[/W,A&Qf)2<1D\TXYOVBSE,G\YMe
@VO:Q++TaQDX6(T&9#(TOTN5.:_c1QEXJdHDF+N?1:2U[_ebK_\ST[fAZgb<&gVS
&.12=Z54)6JR\P<&4(/D;E/S3ALKN2POLV7WC2R,GEgBS;g>VJ9f(0OF3-&gLG-2
;eZXUO?]A)cK?[FY]\@/+XX5dJ^?5F4[AB.S+gJ3-ag5C:TQM56/AgcT-Y[=gP)>
aHaMTSDRBB23A3\Q(DWFOd??>,^3#,[EGW5-aVdaYN^3V/=#MKY+3cAJJ[b>]ZA:
5QK\cIN##?:T)WSb&=7AgZdI&A,)YVcA#LDMH380KA?J33gOI44U\YPVAAc2/4W>
aR.Q>RI)U[TUM)e.P8UBAd>+fcNc[(S8>E(W0IOY-MX9Of5^X=DTN>WHSOGLbX6(
Eg=<L72TB&,YB3Y.X(>M9FHP7^B>_1H0S6XPYGF1F()G]2&Fg\[L7TU81WK)8#;(
5;W&/W(gH?C@9QP30BL,+LfW\3M]\,BcX9T>2BGCO[d][7BfCc^JPI+f9Z>OMe#T
VY4-E5-Z&;LD_;3A/RcdB@[ZT-E;?&3CP@4W6e+6b5U@B?131+PB0g)-2_>6D8IE
56e[S6P5CL=#DE>C2cTN3]#9aP-L47E)R-^C-\CC]QL17d.Sa>^#(822UPN?V6JX
g([56.CaI,A2/faERMN>D&XI[UOT.1;d829J+<(T:=/ISL7^.WaSFED-E,U2f8?3
E)e-KbfNg2#T.cT>S#10C+I3&U;0ZAQR2TIAJUceLHg8)<g,BgL:(KM72:fD2>87
K0b)(BAT8A)MM_WA2NFT>PXb<QEPcHA(,R+.DA6<6_a.CQ8_H\SZQc8P>_W5>NCa
3,c^Y2(VW9;(b&4D.V+EKd]X4ABHe<@#C<c,(BM2?-SQI5EBM]N7bgRZgQ\@K+J:
9\3<J-&N0)-VaEMYJ6K=eX5]8Y-7g;>Ze>BJS:HWI5>BZ/SB/&HUW4fgZ>,PVg&3
N^Z_+0HW4B1@5&P,2ZcfJG:JYR2@4RA<Mb(X6gXTR?FdT6AFK1bgA;IF)A7-X)I=
:GJVI2aSJU2,.LAEX^3#+@SN0g[=3YgK7WG3NG?Ia,g,H0ZaV8aELWa:8/A4SZbL
aUbGT<SfP&C)D2P\d&GN(Z1eOQG?1/DA)SO_5GU\0;aN\VX0V@,:#,H\BHI7-,##
Pe6+;KOeRMOgV;55SGa<\I.095=PgL[I#,&M:AC6\.,&9X/M2UZ]@R;@X)XL]a=7
6#CES6^\(@VKd8Kf26V&0=eMUUC<<,f+D4:=;f.;298A?;(#&6@TbLJ4<egTJ#0(
gZ)6SEa6g_H49O8JF)BTEF&Kg^70&.eb.FZ@SIffBI,.a=(94bP<QOCK<KEE>F80
Q7eGRE:;P70B#RgK?WUd9,8B?)=f;IR4,;=\RdID;Z>Rg)K&XQ4g>d_Yf8DfRZ,+
M,R<9cFJ84MCW.:#8/.EBSOee[WbPffg+7?gF;Q#FPX2VPUHDU(XLT)H/J_^Y]Jc
]@L+QP]8WWZY=AIM=9bA)\6cR:fBQI;Y.Bcg>)O<2RG6\T._3VVc6^#3TWR1ZM+1
0+Id[T&cA<\ETbFW+J4H2]T)_-/bf@F@FYb8(9TQAcU[b61CJO)JCFCA5Vfg,J);
XRVVEK+,Xb5\J5fWXMQ60P@?_T:gV<YWQF[PcM3beZ:f8D]90ZU6f,WM0VcQ9;2-
VV5^O&Uf94LQ34&H)44=2)-D<(O1H-04Q.f&2TB<<\[[Q<35<a1_M-,M4XO0QfT<
/S<g0Gdf4]>E3(LA^KBKUJ?cDfTdCA/;ETJ]T-O3PS+5N5_/.ZD4f/7:80D+;b0)
@-@=QG_#H&?UbJ&<T@QTbQEf7)(d9K.@(XFL6XQcB7THG1#CfHPV:?_)8R(9cP.Y
-fe:9(;e5:_Md:=>#8.P24-:Jg^cYUTM0_dM?ccP04dC<fIXES#)33L)?WF2+Z[F
SIfU:OB2B+\^D?U5[eF2L9:5=6+>#F=4MQ@P_,+5@A?EBS3[9&)?CB.PZBPY2&YL
95P,O6G2f-W=JVP.[_)7ROA+/GIB[a?,?<8X()Td.ZXIRU]EQZW\b_c^0]fb04QG
Z2L;C6G];c#8N#/a2N+O43<ba<QF&Y^gG(I,OMN;,+D-[UZ:@;7?Gf<d(^7c+Fe(
5V+DL;C<?WFL,aSKA#.c#&HC<9DaS<(:8U(KR7SQHF<)\(OR.LgU\\&N.1679aIE
SOL]::[#772aW=V96/<baPH5LPGXW,,W+N0<5-4AC;@+NOP.eNC;Bd,FcD=K386J
-a/9LEZ\XSb7=AaC>YI-gI:cIBZeMM,]@35e?T;^JOYQ]PUdg]JK)WJ6gg7(WKJK
NcARbJUKU^5JXTMTFB);;dQ1PASD9BJXMb)6(b/OMG&#A\BBg_[FI].QF03W(.9?
?))<I?^e2(837S<FUDYR([KAHLTg?G>3d0H4GPgb4II^c3>GF^f&9:2aE+.5(86+
f26_LG+C81X-66Q1[&ceY7A1;/CX2?-0?:b#3a6:W@I(;KXAX)Q,33>&AgY7cG[6
,@3K4V@eHfZeQEN=SZM.V4F1A#^Kb7Ve8R1&KAF5QNFb7bF6AT20?dK581ZIZ@[C
;EZ-fJN5]FR9I;8C#He,AFbNe<a5HSAJ)V7/O@,:bO.U.G.5FR,B&@4GbHb_.CII
@(&d]H@1VK@cO6X)?U0=WP(0P.=M;9Y>c7XVOM7R7.8g+XY2fT.e@46^^Ga-+SdV
cceVE.HOPQP2+:>93([LD;,;MNEDe=gbIN]/G\IJ+=&D3XP_]WBeZY65gLbaTZKB
6A(L01W0eDQ(^WbW5FD=^W:-DHJ\)[(#.eQ(HW5RQIe6>g9S:=JN2)]U]4P(2#T6
dBKQ9/[Q:VO^A.e\LY<_2YE&^F>WXeLd)8KHNKVJNGMS?6>WOK^#4+MceCCEN;[P
b^97(_cU#3A;9CT7J6\fK1>VZ7TN0(EXMc5T@g1RHGW\5-HTGTe#[JL>^,-K^2#8
TXD:G@2(TXAe9MMbDP0E7gfD1W]RW+GY:@P<gV_B[>+/L9fA4Z1,97dH[@g4<+R5
5Ua7E\VMY_[W44&b5;2S^7NP4XM@>b=Q+GOcgMI[=XCe/9+eI[++Q5UBcI>c+B>f
PI_O5;PV,)#I3f[6#V+B(TDGSQ8#BNVdU\8_V49<M/=e(5TN7M\f3ZG2<APBD=Wd
.X>O^4]O@1XL-J0QZG:g7PbW&^OZ6;T^?_&F0;UKW7#d:64VVE7Q4I,?&N\7bRAR
bfOf1/J6AadI5F[O_>=J?J1N#@RIN_N_.1^;DKa3NCf\ZFKgH[>aSdWH0/75b(J[
H_?>QfPQa638K87]J?85MY0G(ENSPG\^9de]2</]:aId]S[d_@GPD5G5<JSYF;dE
-/5EO<HB9MF<<,,P1\8bWJ#)S.OZUD6OeFAJ;Z5KZ71L_UN&a/17Q?-JeF(e7UD3
F-L6T95.7R>S?]>^)(gIMO9ETE+=H;&7+QLX@Z7]K?UP_BB(_C_@.92?VX[]M,BJ
aeR8f?-IDI=[1V&0]&f&K3YJX:JH/8d7@_e?gHZgUg8)_NK64bBIRf8Q#EKfCKYd
(+Add-UA\a>::OGad7-Se<;0V:?3EW3<KHCB,HW)a+YW=c/9-P?ga8aVcdX(E7eU
@Qf)D,EG#IbSHMe??+2X[?^L&Q:D8,78cT+e60RY^e;D5=8#(Ca,MZ:fPD:JP4e/
JK7AZ5D/+f[3:X:QB@Nf;49ZI=QITDMXaWN1YVG8eX&+LW074+e]/GYWHZ:[A1?(
ZdaF97V4+G-:PRaWEE<1,U^[</a#RVW7I1#I]S](WP2R6HBEJ7KW:5I<BQ03[b-b
T2@_VO/MWSTeR=G+_L@6[SJ&a\8+9+72PA4@5I32L98<N.Lb]<I;@TQZ/3f3gUS0
0ee.DHgJ<;aNET7Zb4<L;P8(6X7L?>>eI[1L><S5NfZ-XN1<62<Q[[J&),CYd?Hd
a2F]#P_T4?M,8FKU0HGfbYc0eEDa8GKZW6KC22?RQQ[OK#^:TfV8RQHASFX3ULL)
V<4=7DgW47/G&2XDZ(WNG,96XOXP@K-Y;Y/9ff7aZ&ROZ#,VIP&3+D)d9RIR[8RL
8TYSU)Z.-BG@@-+bA6aI?Ye1e7X7#0TO?6>8UL3BNRf;[3]#/Q?_H#NCSF]+;(8V
Q7bR.IcL1=3_=-XI:b=W0,>c(P>^3NIdUU_R,&BU,)CVLP5G0_U+MOg(Gc?Jf1@Z
,@gEe;/5\aXcLA].L?#,K#K94X?,Sa<d6?X7aE=IVg3=-VdF=d5323+.=P(9(KL]
9fKNXZSd@(.F;Cdf@<f_NR2X-A.d+f5K.-XQJZILH,^GBa#V.fF:\N_)?:SO-:RN
(IS].CJI#+KYX7Y7R+F8?&2c[.Z#Gf?GSS#A(D&^Xb,K2HSTYF]2eRWdD#gEF9]Q
E2a]SJQ2ZbS/5+TDKO[)EBQMVG68V@Qc@41\7#9A;?(R=&e@SCE&d-Y19cA@]E.a
XU&BD;IVGeIfN5A3ATXfMX82LM<-fAY\,SfBM?BXbX9XD2.QMSd2LJR(g;T[A2fT
aD@^c\)gcUDHf/1-#Jc:76Y#\GGg<KM:Zd78#RW2F@7F;7+MQ@e06CB9O47ZQXVM
d0^]7BWVcB6@B71\;2JO^<^#e_Y:2;A3UXHO0)eX9Y)<^P[YB-P,O#b/.Ic>/F73
#-X7b&FE-.GNCTMAN,?)-K:RTFW:HXfR45eWZO0T.d(<=6=I5EWXOA[)J60O7I4d
EW]6&VQQ<W:T(4KbX?<8ggR-c;MXAKUZaO[WZ7R=79I+HI7QFO@L[aG^H<(#>K8f
9cYKAbA.I24?<:H57X85E,^_)-#5,2)YRT:#eYNQEg/6PdP3@RM,,54_=P)ReUO)
34d:QJH5Pc9cYQKF)\gO_]O?DOcGLVK.&F-J0^3cO>,Z)I]YQ/d_d7?O+^=Cf6X9
a)^\K#62e:5b/V]G5Nf@7/=DNXVCdC#715.^RWGJ55./,YBB550F&(4\1K&?;1Z7
QN>7Q[#I]25OeDfIXDW&e[]H?UQTAa\CH==E65eXPREQTUE9>0##c\H^<NCPdECL
(@;;6]WK@;QW]>.-ZJH^=0Oa<)ggE77@P?HdS=]b8O7I[2V>.H;N(I2JbMZRdV4/
ZaM1&EV@8#eZg#],R;dFUgf;V/2Hg__NYcT-,\J-fM8[2\TSI/MJ#)Cf3=R,6@DX
:GU#<+?1BDK6Y(L[>^X;2G\_,WR]VbFc_TR67YEJ9Uc2/GM74Sd/C--LYKT8cXRF
g6=NO8gW)ZdY9JX4T;IbZ@<TGLJ>-@YH0TEfDOWQ/,Hcd>5]5+\aUV&C2JVd;&+0
Q4@AM07fc.YU8T=S=#<,gNM8?&>.X5.3fKCf;]LeVJLe5ab7\2R&FA>@>QCN[R1T
HH<aH<bAK<S:M[KLM:=dRW1QR,dL(8A9M1@JVF9/BZ_0@\UZ73S^>X3.WP_90#BB
E2GSO0+=9e@MgA08>&O9=OJ3@(9J/Ubg@Z]?#cOM.>6]QNgSN3.CcbEHM)ISR@gU
Rg(26_<<aW^C.@7@3VM\UfL4Y_YD(:Fg,?L^#_SUFQ)-gF/PdI^+G6@<EU.WT8-S
WfD\?C9./3ETX,:4D\HF1&KSMR[@-e9^)[92]Y?&S.3fe.a86;YBUPYJE6ZYcU,c
T+Y\13G,gV.L3aJXY?8E_L@<c]6-9,TPKgW9d6EE;6dMV(\)-6bJ_Ae9^2gZ7GBG
&I0QIMN:X,=16A;aO?7g:H/YDaR&-a3Id=UQ/H6L5,T0Ga57IEE,L2=H#1VAd\Aa
>e1d]-b,O7WK12ECe_.LY=40:PTM9@2\C(_Y05&JS>L\@P4/FSecSMJU(C3)7\ON
UV3Y(<dF)XSO6KPR0cRF2MHcZRH@?@\VAN<g;dERgL.]T?@\E;S3SV>2ZG&AXbKX
fSE?HTB;G9>DG88_OX?:<acXPdW9Fe3::66;80_556?LAO5XVbW[7BQ:3/3TgbV+
,2d-P0E>B]]@C_WeI(]bA45]?@-Y\N&K9D)2bV5SC+Fc@@(J2fU9O<=N^P)FG#V:
?b/OcF;A;Y3gHOU-BbdDdM0+O6:^N,+[E:0C@[EBT<,-8Ad5V76fgF=2WERC5D/+
R^,SdggQ(O2JPe=#QF)0TJ[IXK^6f)1+TPR,<@gVH-PbH2],3AZb_VXB2:F:^PSG
I_SeaL\F8M])[?5NCT8)3TIKJ#Y3_7YdbdERXDg(f37<S&=15LTC+<A/O.]WC-UN
#\5?7f9f1P9>FbQ38@@_Y>e)ZQK&2:Gaa+J7+3];03Z+,9GHZD@bXM4/#eU<.YTD
bEK+\GM,a9c(DF(_cZYC11\4R3R=a?.+4]L^K=GT+.URS\Z#(b7M1240XH#/L.aP
E+OQ/@?NW=L-KW8ZO>TdFc(]&1V9.-/N-)\\R.01XX0=,)+UCH7Md1/P=JcW]aU3
K9J\JgUe[]cEV=0ZIP.Yfa8[OT]af4AMSWE_W8O<(/.ZY)C>RM5aM40P:_BWe[YQ
=2)5BS9/R5-.2N;+XPKbD+XJ@]@F2UNg:#)3<F=;#@1MaXI;CC3ZEE13L<T+4cHe
7FgfW2RFWCe7(576^YT(46b;PTd=4G[6__R[6>;;SH:N)^fHU4\R<T;8^26Z,)<L
]#3_N2B@5V;)F+,T:WB(DMaIO]=>UV?7->Md)>G/NL/K(81c?316e3RPe2+;&[]^
2[;dKD]fG3NLDPS-4Y?D-A6Q<587=Be3R<^(I-#9M&N+)&S_2I>Z?N1Pb\/A1NEH
&/QV+Ke1fFL^1QS6bHEefNJWUK<)ULRKGN27OT8W&C:O_1.bK^#492\;UZ,=GO]0
9D-W2050g><;@Q+>\#P_5fHGF4V55;<A^Yc4M.YNe;@5X^F@PESLS1]Y&La]K(gX
#>1V1Z=HK&+1IEEeUW7e6]JW6V;6,QFV&;,fEM/^/]B(Y&F]I&=@R1<T9X3S;7K7
XJ86L]DC.]5O?9-5M+I4+NaB,@I]\)<7KB#<&JJ<-W#H;)C;X+CNK1S3+YULV\Ze
8\-Dg?[6PfCaCFJS2U,g2gH,:+-Y->U0F5VE_=g7aNUf_8aI#aRE./dRHUBTN[13
>cACFT7TK)@&G=2[K3BM.B,=d\AH]eeFT/,L;2g9:.B)9QG-a_[8@BK#<M3e5FMb
>IS&U&0,00ZU6=GMd8#Ya=&&GNBbBgM+S08ORF.e\9@Tb]W:,&/+0\W9X9-g6B3/
(VEHUe_TYa^_3#W4YfZR.CV89QZX,>F:MN/3L,LR6Y0B\ER]aNM8_IY-eB@?4VbH
2F4A,/>-GID_#OB3_e.Q74.TbI>&XF3VEb]SebgN&b.532O?/Y^2#.7959[78O@1
L/4Ib:BIATQ>e7&?^-@Q06X8/CYP5P,.&FJG_L7>67QC:]T1;I^IRYWI:D/a\EM3
Z;ETdZ6C\eV2,L@(I,C]?4I1YV#O7[XEM_2IA[)[B+SJM,O[?ZH&,C0#J;2aagE3
.4D:2Hb6bU44EDK/D6X=b6R?MZO+P.V>B&I&dKZIMF3]MENH[Jd4.0(aW\.gd4a9
K476V+K)aV_#BB2;?1=#X49Q-:8I51^eN69M6^]:JJ4R4?&H/Y_E,dY<2W240P48
W&[YQ/cS(L6O4Zc(R]d(QJ]RFJ.6+@7UN<T#4E\[S:Kd-?=<TK9M:bbQ+2L.KGZ&
K4@HGFa).]M2F7g?>0KD=.>2H&O#@@&1HBB[=^[5a;YSMYQISSH2_8XdL>J6,]A:
Vf4Fe3[dZHMEXMW&)a3-6eA?dcg&H@cgE4:MY\&6D76T&gUY<1XRJ^T7R7e81ZJG
>.)f2<3Qb9f\U)J<,[(D8[WQ22SJLW=G\?EF92KZg3,&IM4(B6b2W=BMP0ZX6GV<
eDe:X//^?0WFGNP\X[_R-),WL2BHN:6XW@&9839<(D6R\#IPXPIJ1=:KcZ/6ZF:[
S&WFgTX3SUTI_-4B&UHW_dJd,(Zb5\1JGH37/GOYdP):@\W+>f]a@VR.XD\QP9?A
fPV2I@U^M1/<.,6:B&K.)]SA^W/=,T=b)0RMVA(<B5_U03#M>]Jc&>g;W&:b:C-\
(@HYOZ[J4BI^UMa,eF<#J[d)G#-)#,(B^6-BRHJ3eWZE=_@WN=9:U)8GQEVQ]J;>
(#VM5US;O8,Q]><;9SEI>.3eDgF30PZ/YHE1<(?f@7#&17#:Ud10()<+V1C.KVBa
J,a#L,dO>/&UF6+VCQL^YU,Oe,@<ZeB?=b1#U(PXgeNG8>)0W/&?0aS5H9d=+0FA
aKX,S9e@_W/)#B_Q1,;+(\K@ANY^RC4F3T#>dDG#Z,NM>ZE\W?OUEE)K_S:=9H?b
/.>SDX9WA(1\\OE^I:X2[(LAT20IT9&Pf9(aCOHB9)7@5DZMZS]8J#bB>TT/;,E:
_-fN08-25LK)=X5JgYS/T3#9;^@aC<&6OOgGJVc/S5O6:_,+M9PNNWAc.[BT3a_M
LPJagVR-\.d^[;JH44ab+P6QG85ZI.dPL?eD_GU83FLB[2Ef,J^/b]#T2GJNYdMM
H:Pb<M\T]>CcZS(R5[,>a+NLJ4M,4eB4_B0cKU4cB&8J89&>J@2:.Y0XNT]WH^@/
JX[1JND63_RfLN0&>df#\)fU&K>WXFOCQ+/I^B4P(F,VUG89.RN]^ZTN)ESKbYZ[
:<N7aG(=VQ.0YHc\W/I1UX<Y);@D3F2EU<d\a@8Q6A9AcQEEYaW1&V)_4I04U<3F
AKH]J>MZ3C1P:HA#L#L7F:?c7^X;JDY&Zg0fgBQ?U^.VJD;H)=eSSRG_-9=#9DaT
,CCS74LfSUKRF44YZF8?aMW9BR:FYWF+g&LA(<+XL^\HY_)9cCU+baK5GH-&HP-_
+fa;)E4@EPU^.XbNQa>3A.O6Q[#F7P#7]U<XL])G3DJE[U8(QTYEY[=PJ8@EKKfB
eRV0LHBNb(1KB<cbK8M6Ja9^@5T8M>Yd]OK^3MBV9(caeMP0aT:7PH&H230158QB
Q6G9X2Y:]_<NV0CAe:dd_++5T<K=_ZKS;9#W?)9<ZB6CFg)d2+V5U0=-JD^PH9@_
Y#B2@(0DeTbA[MX,J;+/6X/IK;,Q#ed)D_[S:N1L]@#\:4>/d;KdCA2T3)&MT98d
46<HDg19dJQ)W1:>Q^NUd[/UCTDc8f6V:NC<7OGV#?A?WF/=K0/[(][02e.#8)?O
P[90PWS;f_>)X_));gMP@Q([Y6=N+9O<f,9b;T[.J73:e#\R;gC5.8.I<GYYKf</
^^4?O65+HG_[AR&==L5Y2V1T<5cg,EZ2UN7;64Z:^^C7Q,Uf8N+T2FJ:@;)-,H1(
,:Q)\N@J&-bX/QE?\XR40UF=;Tb_IRegS202SJAZ)^N&9I=JOP\937MgEM<fYgRd
87YbO6HM-7b2c>>QM;=P;HWFKdS^cT7WfO9NG^IVQaC/F<,ddT7^<RdW;)>_0R6#
MRD-_Pc=R];F@#RC:YKI4bD/X[dB<W;2PMLI)-Z)^T8.;c3QFDgPBZU8>M6T7@C_
8H9H-_PY?^N2f>(RB]3&&,;Uf20c]Ve+M1c]NaF74M7f9N(2Z;?X#I6PNNZVG9BS
^I)IKI_+Q&5GZA[=KeZEL0@(b8(:e(aK]5B1ZFL,;OI)&[1e_WK&[PUP_?^>&_9&
:S68+/QaO<,,>]#Ld6AU.UT56K--OO3NeW)8KPS.-)]Ae.Nf5FW,;?7:\fDGF)-?
Dd=DFC<\J8FBURHM9g=CW,@XQY,g8CC[)_.<9XFX(6B)UR.Q8@T#JQ8A<0e@:@(1
.PeNbNgXZ/:G3_=W.TW1W6#C]:3T(5I+&IE6M<ES&47-=,7&^-Nc(N)7G:a-dJ4-
g1+/>c@VL0MF^Xd2Z=6,-S8g;XWS6JSA6RD;:cQ+D9RZ-GMP7Q_RUU+E74-H_YU,
2:[.)ec0WJ13BQNA<(BVPD@+.-?0(7O-U44I:>)>1XO<D@35Ub:P_&A&ZM^4RJEX
FH(L#_?;&fXLT6/#4F./XN2KUNYB0_;2@YWJRLL#;OUSa3(ePB_Q/9O?)@Q;gc+U
AH=R^PMIe]b4[7WEc?M)gb8NUDEZP9(7UQ<)d99ddG1L()BFJFX04DUcZ&_.SQ[5
W/_##aXf:K\AQ#aQJa,RPg7ODMA(B(_BX^I#R3D493HIM9K4+X?USTK38B4_L;5,
W93Z#6aJHe[[b+@&G(gU&4R0(EVW4I,(a=\:fXVFcE<H93[3>T6G&,2K(LD1UUBP
1QgEE-6)S)V5,BABfEGM(5Ee)bB/FId-Aa+QJW/K&AeP#C;<V0,/4+TY6JI@OPRU
6&S6LZ9I[SL-37U4DE=_/L)I,W?^T-\(e&_aL&;]EZ@LW:\M,RX:>H6FMF8SSMbX
bb4E\MQOGOUDF_6e)Xe[2fP.X\^Hd,R,bI\?D&aY(#N#ea^L</W4=6F&<LT^_KA#
1_+9-Bf&5=51c>84dD7:QKT,<T[6.KD]eUBJO&1#:8[:,0bW24\3D-#8c[#Q@-6^
?>agRgIOHOL.O[9&&CMTKfY(eZYMOceA?DJ_&.OZD60/d:+gU&V^--K3E6VeK1AK
NE2JME/Vg77Va]IFCIEDQR^)NN@cg)7I6.F:I@b[946<GbG)1Zd]+:58=:X<W2+[
BUV<;-WS>4\D]A=(bS^NF1fDg=^3=N.Oe)=(F+g8HTg+3QZMDcDHI8XDDee[e)d4
eL[>+:6cg,C#:]c(87M5#.QP(DH_8:PN#dD_X^ECS&2XAb]&AIe+5F3+DMXaQC-,
PcNFf1(#GUL#IJ4N:WRAQ>[D)J>8.Td7/N]#RO];Wf+29R+AO5^6#+G@CF_\H#,Z
V6:<Q>W#6B>S7EYbIHBH:E+Eg0.D^,+>3VL?KeED5cFJ1c,MYNC/Z<FTRaI&BQg)
[FCW/&/OVU#FR8Ie#=C@e+10[G;_#>[K5E@;6fT8MUb,&0.-A7?\M45Xef2VGTS,
?>I/+fb9P=>&@K)EK7O9.FUF^<,8;<#<HdP78b7MSc5R<Vg;B[D1/K,HaI5IZ(If
E14K.4=\O9&G(IfVZ)WaV@FE;WT>L\A)BG+KcP_].)V?2\a&JR>+.O6QUTI/TUfb
>S/.Y3HD_Rb=5;N9Z_000ZbELfHc_[SG&N+P)B@(4[G#;e_1IMSI;7H^dAgUNX?B
O3+Z7-2[6U(Ue^714fVN]G-4dcd1EH4Q>FHPQg?.K;\Y/9OQ(>@dR=74dIT#E7cS
]U0KD9a:2+H=eZG+1Y]7&ANO5)\5g?1FF1c\TN;RD8@GgQN3=K>JIeTcO+g(XP^#
;Q&dYBL3a>7E8KG??QaSEIJ4(adYQP&@,2b]EKQ^?>ZFL]W/g)T]E>cfVCFZ\\XU
EIH+e;5-^=_<.#J0J93GX_PXQ@29&WV(Lc;6#//Mg[XHMSRWJ@&,[1g]^3-TQ65=
/B_Xb]NgD3JVN5e6B0-?]Q1;W<L@g.de_;+@G82SO=d(bY.,BYT9MX:fX9MSY[B_
Xa\-/(W6EAI253ZEINNO#;g]3c>,B[PXA3)45)3_PBCSHeHS_5MGT?a--L=U[8A6
Q]W?d(Mg.g\d:bL)(4-b^@dTANgJ??N>-@9RW6=UcZA<8GVD\7PC&,PA&aU)-8P4
K/K(KR.[+a-ZA7EKcXZONR,^FaGVK?FI)eDb9\H2L=@Dd-F&2>+a3DD@/T.PQ1aJ
@bPEN2gRXA8NS(]88TcLPa?7H#7b-@=&Jb>EC\Y+dcKSL?b<=dK4>-2[.fF8-(4&
J9>@>J)Kf,E>,B=GA?@=O\0^a#+MAVMcf6g^df,JQUDXa_9,\U/&MW):e/AMQXY3
@9(FKH3C[./22U#G]?\P+aG(@f3MED\XdQ-;aPa\?#,a=L2=@9?<bRJUV.gJMgN-
EPdI3P^V.7O\NCQ;fJ1C3V8##HGKX-6Q>dWSV8F3#;_)WF1(EC;SUd>C4LH>WOCe
AIH0VI7/#242b0RXH1S]5\d[R]SdG4X\&c1aVgY2D[P-L_UOYEeG_OSJD6dJ>gD4
e_eU@::Mab55^]6,c@IcAE=4O<6A1]b;KBSD[#a.T.H</a8MLPV7;2,GUaPgb-c^
#(3</S.5&e&@2D,=b,;9=.a83J])[a_gQf#+:/c6X2JI0U61@fVKgZa/\PI(/6VC
^,f,33ZfF]XF7PQ7R8QgPC<]OVR@=W2F&d\?G9=]V0)MgEUFC1.-BS3O69W6,8LS
9IX+8TUL0B+cFG(^c#ML;T\O9bQ?\6c?3]/^J6?>Db2(a[+.;&U7GdLNGRZcb2WA
R?+3b,DOe[gN0OV?IQ.aUSQ\;8Z.aZ))5C9F7f<8fC2+Ig2^?F0e8L7&MMZKE^\#
gFGd#X9c(BT(g?4bF\+Kd<YE9Ybd0F#V^f;;9gI&\92>/396JDT\S.-(NaR,L/e(
SEXI@gZc1?+F5feeB8F@OTFU5DDM/3#+5QA[a,VKf+OeX0O-M=,85VWgY6FQd1<b
@_;<B^PC>@V^dTE]==(WU-L+Y4J(U/2>474g#VX5([5PM4-\d-\Lg):BGG@[;9MF
\[g3>C?;A848_]BFa/3#P59YC4N1M.V2)-2).]4e/9UaBQM,,EGY=[(4OPHD-gY5
NcDVPD(7D9-M[a\:,T,[KVQb@V(=(47:Z@U&MKVUIR)be6H)8>/O>+^UD35LbS[+
.N0Q9GITaTB(O\)Wc[R?d_?EaMVAc.5#ITF]#/(I:869FNC<W7PB3BTb\I.SPOMg
Y=;PHgO@__E9HB]e2IM1-)Z.3)8_gHJ,6,#N,[_&T9?&XgZe^^dc4MKU&F[/T4N@
(-4U#^7]ccE04Z-Ya5N;TI/M^Y<QLaP<>>HS3ODT^4b?.S+4e5(UN.)_4b]Wf-&P
VTD&A>N_M&E-:QWSIeLf4IK4/_#gOA2eE8FC))]ce8_P:7LXeB=_cO]_Ed>0TgHV
HS20LK2?8FN97c,CbYN:DQ.7TL@3Z0^UR6RMfc@1g-F_VWD.MG:BQJVU@=_=\#(Q
g+;H+aDd4Dg/>Q=E34WTJ_\LgN1(1JSbb6>2V;IU@MbdE(C58aF@b7JK&-G_dAZ)
gUZf80_:#Q9L/bFTFHg;/274H6F,K_Vf1f-DfJ&=QF4;]4@=WOg5)D(AM)>aeDA8
bXQ/W4;f(BU?2H@.CCV?T\1(=O&B@8B5YH6MZUR(]f]WbNU08dD7U&X[5Of\\+F>
)8cCEPg979d9XL,9G<[EM.67/634F.R=Y.2+=:OHS:4T+3f,4,?PfOZD@.P/M:V<
[(AH],bF[ZeZUC2&/L1A,D(@HUT.\Qd^+3d#>4Mf._KHJbW[ETC#_RW_/8:P_:D>
H_S86cWcbD[b4OD8:<L)DV[WON=-NW7PJ+2-H@gPd\32.?Y25O9Y3G(;H9>/D3&Y
;0&/3+(W(e(1CC>>ZgMY4J&.]Z/Od8;Xf#3/J=9MC+IBFc\Z?-N5?)g4[9(7XEL?
E6\1JB.@8REN,9U4L.5NMBb#C_[RNTOc/430gO>WUXD\/R>U,N7EcP+7<?^3KLWd
S]OdR<M6KdJ[I28\76,2Z3WYG^VVDP+3YWHbM8aLC@WH,SNJ)5A5?2L8[IC#KTRM
fW?&(>UHUXaV=7ZOe0[J(^)CEcS6I^LII:OUMLQWDLM/;/<e[@:VA;21RS^Z.[D7
R/J9GcXC7U,fAa;D/8fcD/_Z),EFRUb3<dZ^H6@gE@HI@b<Y3:UB4T&HbL6P1D;5
3J^b@.0=Y@eVSSO(N15SES)S]@0:SBNcJ(WI.ML.g(G)a2<:CE<W[Ge-LXNPG^7^
bda#N]ZXT4)@/OeI\B4GBM(?FSU(E5=(Q_NDIW1>FKAc,IWd)S9gV:P\)RP&9/E,
M1D,HG:+A9X?@8/fO5>P4,Re]+,2,+S>J:#F,HZ/THJMc9RRF#BU@XUC,L6NHKT0
7.3YT@+F_B?SN+2(YKR2fCRUU7?3L6C3@&T?dF-26NXHF2\09/[AQT@b?&GCKPEJ
N=JY#c#4_6L\@E&P?;fXEN1egF&c9NcYeF+NHM77D\@[=[a.egS(aR<=^+_8[P3T
e51ZMdT8L_e4a;(7e2,GC#4T&1(.L;ef-/e+R>:S6OT4gdJ79W(6cg:c)<3R^+;T
e37(W3:.faAN2S?XOXV8(&2Sa?-AaF]CCVNE&]TTC0<95gH6X4SG0f]NZI(]>I[E
aUCI^W;PU9XSEQMKJCcS<SK_Zbc4GbGc;[N-cYZ:a[D5(<f,8\DW0.fE4[](^DOM
Z_W\>AS(5V:SG-<&S7aE3gP?/F2F>;E.MND2bFHL:SN?D]R6O<J);g-&#Y6=<g+7
>4Q=,VTF)WY2Z@QZa.)f9._JK@Lc7QW\;-&J99+DE]1[C/dScEDg9R?6@5+A_I36
-JE#;A_-AE>A?_Q#+(-(B+T2MdW7]QaJ3YJ2WEW56&P3FBN7)e=2J+-&07_3C9F/
7bMM^__3c1GIIXRV<QT\]4:-\=4R/c<1LT2W>d/T,H==>G9Ye:I:TfH56fbLBN.Z
S,Pe=5/0_9fPZeEUcTB8V&&4ZY_U:]J8;<4JV1Z\K71H0][V_.DOd#]R2]+HGSO1
P[U/2[DgV?S#\UEb2Z90>[E3V<E^FHUg>&<=#]aZ3F37()XRS1(YFAa7#HaE2f\C
g\Gf;-P+;+gP8LKCBGQ,U=H\\2J4cAD3W_O6P2Rf(NW)bR6;+\H<7Z-]Y(1I+]MA
A1136M)8E4dD/(9eAfff>O&4PT]V0fXU(#TT3P4]#6K&HHa)]<A57Hf5=9A&@g:K
W#a[ZE9UG&+9W_,@+YP,Z9dJ6L1JJcP\&3G\\P5b00HDE):.X)2SYVO,V6Y=EY3,
CSI6QE7:+,1<S4O3SP@X+\9IYZ9<V^GFe-^RG];X2X)AB?D)<ZZ[I0-:XgYF8Y,R
/)7b\/DAK&BDZO1OI;[Nd6b5F>VN^4WYD?CS[[J7:f44444HgTMaGT4Od-V2CTGF
]#&FJ-X2>3MId8K[,DS;?2c,\)IQ@90^9.ZF+;A2<fB&TZMD+]X4DX/\6SDf0CB)
&@db&9gVF(VZdDC-,FH.0KLgR_=HJ[>]d]>7H@L9E-cPdCN?ccK]HYE8(-L=751F
d9BV)CAH?8AC<<T\bBJPPbBFLBG\#QF,d.fNWJ6=96IZ?bG0,W71JHN^W1=9O0XS
fPW@Kd;gRR7UfXf-]?H@:(VR[O4gD_eRgeRT(P(-?]P.5R[@B10FRDR[8eG>aQ4I
1##;99R>MMT/dSa<R,0.ZO>\^@KeA,.3c#P6LZI1Z=gAK^3.a98&\:BV6H<c8;1V
40)<fW/RJR7a3Nd3A8Y<FTMR)KP7HYJ]5DR2O,0)4<8GXEaJX<+1M6M38==22V=(
:W0OAe&(E:03C@.b:^VD(2F;XGIVD7&;NAFTddN-8E[(Bb?\ZIR2cN=B\7#62&<=
b9C]FZR;Z]XB7H?QC[UENF&LcKURSd>2ICF7:OM/[e23-c3K+/,[CU,B8(5674Lf
O_TBDCBLe#DUg(dac4[K>BG9/1O2&U/=SaOeSS^c9[P\-\_W6FBFeRR@?KE,<X:g
R1-2O[3VQG9]?&Mg7#19@Fa&>T@e_CE@+LCZ6GV^)VN7VKUL=eQ)FXa<(CgW<[V4
f)0[.M+94+bgIVd+6\F56]L&)g&?W^T@23(bT_F>KLPPU,T=AaaGGP?Z[YV9,eKS
)_)7HIA;]#c,660FJO#H@]S/L#;^=C(IY^X1P.S:5.a6AVJD55L.ZdI[#Cd[JS/Z
_\gI6a?cX8@3APZ?cAH?.W^-S:?a?U2^<7N&L?DU.6FJDXfea0-fEedWNZHW?@]a
I6H/5L\FLc\0U#Z,2>LG_J3J(J;HR^5dgO0f6>VWfH0O/(/SESC=^>/eV)XC->)0
:KX]PKV.e6T4#Q/2^=)C&Q7/dga3V(]g2T-I1CHN239,K<6&W<aO]dN]aA>/62NH
GJVHVU.GARU/>QX_@\3a,O^^8HJ.0=KY.Df7R_^AU5ec.R&GHLRNF,f_.=0@6^<:
=QKBOD?dZ-U^KfLAEX2T#UNSeV+^AZaXCP&4;KQY]1/PLHX^A6)/3UTVSX)ffV5/
f3bB&9/CH\&B,8.2L_Yd#?&HFV#M=\?(/N24b?=5^<F)V,&E3QaU\fTC_=Q&E7V[
B7FC)8_Bf9f^\#=305+X789e>L:V+U_L]SG\FFO@:VIQEPgGK:4#f8?.-<RbOI86
AQROZ7>3E:,4Abf+BbK^2/f0cgW[\1Q05Q.=J(Q2dE7:I3JZId+]ZR#6/&1Q(MO?
NDFTaa2PXZQ@<)GMf3VYY,-Y,_MOXH@2D\b7<PIL#F/4af,A^f[.\M@@PYJ@@>+T
7\.H0ZKJ7O<WgG,Z^.\44R:1Xf7XW@]6Y>7a54dYde,:0;)gF/MW/+=dAIfMDP,L
g@4ba>b\c4/cH;,>Y=W1U]8UZBJM?3>I?7.>efUS_0L^OI/@MP[OR6Ua\4&Cg39X
;[3Cd10,g\7#-HLAYK&I4VUf9HY-]D6SDGg1VBT;^74fQ]Qa\.LM#W#6.VAUV<]L
^HOM2ODR>U:Dg./M^4]c()AOa)+G)Eb&a?M\[@KEYXOTdS._D/JDYPQ1QeT]FO2\
\JUC?61R2<KbEZRee,V)I]8F;SMHOHb;+cf3?ITPS@M9JEYeWHf+eb(SA1U8gQ=d
g-1ae-Q:&1L44;ZCC+\J(OTe:MR0R0H>?E,=DE:U+bSWLOIKLf/a,6VG2+ZH38JE
g;U4)]_+@KD_\(UcQMg[c4ZK9&3N\M]=@S@@KGHT5V,eO_Q5#a(,ZYNOJU^bb[dd
(BTKMf6RGe[832N1YQYU0(_@E-6M]0&UX2-[-G#[&QC?JJ4&DN:J>/[&?b#acZV:
#Ie_G9ObNCZg9&^6G-;HbV(V:W6#1[b7/@WNV,QSBPKeaFLQL4eb/;(^8J#5>U-9
3_:7XdebI6^OLTdE#PWAe&6)cPf@A(>K(b4E282V).AKbHKJe-?W)f7JT>G7#SR?
L[6Fa+fADO>W,G4EJJQ#^^a71(+aS5=-UV-#2\K,&HVgC0169A:eWT4SE3,H=H]O
UOXF+7cXbGXCCefOe&cS[YYccTJG([-b_f\dA+<<Jb_J(bV]6ZWR;PMWR\-Rg.ID
0:C=_3SLgSQf=<KXW(gfO5XFWTG(QaQT.B?69&Db]GbQdL\8ZC&6@ASfVUfF2<\M
03JTOSDdUT96FDd\&8L+HIe-\g23]#[X@b;+#6aHDG35Ae8<NLQ]=;QY#A=;MYJ)
8LO(?Q8.eFNLD@E-.X\-M)YQcK-8,7D5BHM:UJT)ZH7c_8HdBa.D[8;eS[X8]e=V
Q,F6FYN#W(QO:QZ+[,A\R&aG2H/VZL(L##dS\>OQ\@.D7.?KZ7V/-:/?P8]#^UbP
Bd3A,V?Lg/C6A4&&X3^#a[1Cf83-UcCJ?\L#1ecg(8MAe,M9Kg:UN]G0H<WXJbO3
,>87O[Hg35cLB>@fP-_3>ZO9]Vb2XFX[RN&NHT-^gE7T9>/M>.-A6,8C0cGdQN+1
KdfT6e0OT+05G(P+OP3[G10Dc:1MGH#UcB17]Q-#06bH3<]M\a3,J=V&5TU2M\U6
]5^c^3.TLW.7HH1<bW=\#<e_./(J\R<?FS30>Z8U)_I)FND7\c(Bb]-^\O_f=5P3
54R2F][f^7e=GaRS(OQ^V4@R&2XRaO=RWXc=K]90OON/QV,0RaL-BULf1g6E=bU+
f)TTFF>FRZ)]6DKAJ#DfR]/LK2Q2\>G)9+6cB81c2LXG:TN\HD6B:TIf)T]?MF]I
Y<5WGUH,GNAg8aY)DdK[UF+1&Wd<UF8,51GR;9fP:8DYH59KUb-2G0Wd:J8ERX(a
B13AR0Na\Ld;fZc[7H<9Z.+[b\Z:?1?fZ@-d[RS&A#()31BXeUO_4R:?<?3[\3cI
MNb>[D2X2ESa1.b;65T=eZ8U.UM)ZeZTGSZH)g7I;5/RD4W>Gd+>U-VbH^&[E/TV
5\-9XcVS82(\?XR<TRB@\(^@Z\[d7>>7]I<ff9_B,#eC.D(cNNN3c5_@162QG-f+
\D9eSc[_8G8-9[fD0:>HE-#LLgc;KJLM==VJC623<6M&?W_M\/Vf\MKV<<Z<RJO_
e1:3\,.TdW2H--a_aKD.^SBBaR)QbHf8K7Q)5)F=,MQ<NHHIH<X)3EI@(Q1GYE+3
WJGO:fC@fKO=T6f8:D#C84d->O3fIbM2UB:TV;+\3U8SHDU.IFV,baAYXOWW2):?
U@E\g_-4YMD]-/bMTb\_^#:Q,KW.Z/b13&cSQ-4O-U\=H?7]:8G4GE9]9WI1a9_/
e9Mf_fc2GIEB<)@NR03TXG8ICYe:RUa+d@Cf:X@08d)?/:Q0T?;7JfAWJ:dd<[Z.
g:UIe(+Q&1<8SS5Kc:Z&f(0NHNX74TRZ6<CAC;DL3F=3#Lg?9L-X<e,&^<EEI3fK
e9gYH6_;G#R(P+GLac@EKd9;;;^S=-ATe3.(,f3XE46I)gF:+#J(45>-+7?]\f0b
<bNLZBOe2K#ZSY;K5:J7d0J[.=K7UdJXVg0^E4[.MW69gDG\;IX\V\69Va9A>&)>
I5W\7cKN(QB)#690:Ga(](R?V9\TD?>AQbbXE0+YC7AeUP_91LQ[6(;f:16L445R
2c?J<#@S2/;YfbTC@e];4?b&-1@fI#_b-QZ?44,AS#SJg(0E-H>P793Q_6dVQB#R
4;/-A6(PJcO/50\AE7&L(8Pe+)5dIfZ-C7+c\PIN;=&75gd.SI)2?X[c._JV)#,P
7f;EV0[/M^ScS.&8)/]:?EC+>LJK:51&ED4:/B/,YO2;\B92=N44?5>NX5J5Mf=&
105=d5_=;8[Z)&fa3CR3Q@2I7@-2+ED+XgeYf#EcK9^809U0Ub4PY\9=_(T0^R,1
]ZO9AF>PcfNRb-DE:DDL(aNANdfJ^@Y,4WN<dGGgBAfWOZRB6MfD,+5T+_ND8<[+
^9[.U[6ECYcD7#bCg1QDfe/9S7WR?=EC\-6Sfg<H?a[U,/)3TQU[LI__L\D\P0;d
TI_JG8.01#X)WM^=<QPcdEH0Dc3S)R.=18H<2g,(L0fUe9;(L1e38R?G5;QE,L0Q
(>1I6bWF6/N)J(,>:B(@1-&],6Ma?20\LZ5#2=?D\ZaC>@Tg9\&(b)dABe#9Ec;8
IX8#E)1SY6K]Z3LP/HJ7^E7G\HR5TD&5.<M9c,L/S#@?DPB&M;9<LSI@]0V(Y^G9
9SQ>R9)ABeNf1J30XgHH9Mb=(9T;N/+.[a2B)]AB+7^^;14AAM6J1CR07ECX;-&/
2JTPUHO6V6]>ffS@Eb:@eUD7Z8a8<QRdM6HLB(U12aH9NW/YcR</X[6V,A5,]e^D
9Q4A[A;>3AS>M1U[):YPdA9@&V@^?f1e]dK1D40L6?TM9Ye>5bTUXIRO?2e@3-GE
eR.[3>CXC-TV\M/ZE2&_1E?6B??Gc>>YBd)(YFdaU+AALQ;G]f-49:Zd,Ja:SVT[
);QFb(]WbDP3[:8:@/5]KKEYNFYd-A=OQ8PI2QPE=T&?0?K?#9_0]JZe/eBYd52a
V;gf95_#^;H]GG>HN:6T-5aZ-gPO>5?&XNAcLI,TO^?)+FQ@SP.)D=dK2e(O\IH^
-Z=WX\SgF#a..3O2a9,FT8Z4fC32a2K0g7/78<5FAe.V2_3)LfMb^Tb=B53W8&2<
>>&1UG]:@ZTKG?O(1X8\99+e1@c-O>2MS0R.I[GdMVXOQ[SCSE>c>eZ-=Hda](Q)
8(.JK5QCGY0X=398984cUU4L38-//.0&fQCSD[Z7,e&O;L6]eNL(2R#3g+MOSUMX
,-6/W2TafT-OHcQR6SYW/A#\,>^g9YG\AbYbb)M[NUP),dfI1;5f_4d-UCR>Q8=:
f3<;/<;(<4)fUCD>fG^4MH3KLHF/9YKcRN@RJ;D(X#M)+S.M6=@]=4ZYE[WBKcUF
&1M-0G/?W#L_8.3]2O+T5JF_Pg.Z4Y1CK3?)J+4_FLeV4V?T<+8bA4#2BJB;0BL1
GLQL+AG_UWS,3Ed?4X[eR,#^?aM:HU8##b?dF+Z6A9B;RP9PY(VN7Y8@a92Fd8X9
G@P9<LgB3ZFJ7K>ZUd,JR,G4C79HD+b?NYJEe2ZV8XbW1Tf6,Y-Yd1Z/RG^WP.G4
Z+/IV8(f<Q5/BY,d1\Z7LeB,7U+QGKNB+MVQF\]TG)AF)37P/IYVefJ>4T<1Z?>S
.BObeE_gLc+>9Q>6A9/Y5-Kd[ZSN24d-IL7K9?LT2bd/aDg17XYFb8?P3S@J<S3=
LR<DJX9MBB-27+AgYH9=b\\[(bGP6GgbA\O85@78HGC0K=MT[-E0(5<J9H6AI^^@
[:>\;<@B=94[KIM5:5U:>?1CX7R?GELgaEfQ5G@K()OB0JA3XeFT1)g_OC9\K9<G
fTf.ITEZ8X&/H?90OCM9f+)-R[.1V#9E,JQ,0>Y=FDL]4aU;[L3.@NN@eIB)?2GV
_6_5>c,c[_>[)C+0,CO8K+-+0(@&Ag?/2<Y3WAQ7?,4:R]HRM23WKD#-T+WMS/\&
:=Q.3<<TYeY?9DF>A@g2TD#-SZ4gYAW;V)W-A3N:M+RTXcJgbGHW<.AN1R-?_3#c
cA\XT9@d)8&KeZ5T1^.?\aP7G4I:Ea6386>G#CXUa^#7Q3#GG/9&N>XZ[-/WJU@O
]JU&I-C(9Ae/@KKag5_Y.6=>g?aH6M/FKg<^5R1Db<R15E)<gW?[N>eU@S+_5&\Z
^OfX.[4\M6>T<d2a1PJ&MH\JMS4IS5L)gT>R65_9,ETUNdN:a<^E1L[UJ@>R9&[W
W/Og(Q<.@d_)ZZO)K=@VP&d.RZ(.d\:XTcV-#[1L@5#]7KQRgF;aO^SBPT/\YB-4
KSAZ\IXKcKSX2J^SM0)16?8A.aI-]<b<1F&/2S;P7f5CVQ,(];0X)81IBJ#[1JQC
e&(?dRge>V>J>)^5J.)f-J@N_1X702/,eN[gB#24X_bNM5&c66^T;eLcWKGM=V2X
Dc]fBD,AKJ<+L:PZ@#R;3]X.[g:.&gFVfdAN+8@++3#D\-?751B;Q4IdTKG;BPPg
0Q)f\.NX4D_(e49V3_0#g&W;[.NP\[KEbENLZb=>+K7ZHXLVf_[WLV/YR^9e03RK
Lg<R#?8G#:R.ND4BgTL_?K\A0fWUB2f-1WP^S&+O/WN-@W#EYg_XJVNG;[70?d&&
CZ)&C#dW(0,MT7_A/gOf:bXdTCGZ9Of20,NQ>63YW2OHfDQJWHTZDB:aU:4.EOd9
M]3LF:&#\91Xg^3);1CG]QfdJ;^P6/,1(+X<5O6RTX?[.e?R[GSb9]VZUaR&.0&/
Y5AIb^65WIY?-RH#G^)FJT#+#7gCD8QYSI8S[,F(WB+eL\I87<Q[0FNYOFTVX5H[
Y\]De]S.)J[6Ne6d4[,>AZe0b3K2d/I55NW./0G?\eUcBOE0-<5JZJDZR\^K&:SR
JIgJL\c\FP_P?80HQ\6XAEMDYX[B<c@cdM/SET3:IP2>,FQ3WX?)dYRMbQc[G_N[
H54>NcaFH#GZOg;4D48U<]HY8I_S]Y^W[>F=bJ=APCGJ[H8\d1&>?LRY<1-XK/K7
KO7X3QL<EZ67XJB]CPe1Y=4B9+F3,BB>gI5KPRA[:8ING<a^XDPT7,;@>7H^CYZX
GDEb91O;c&;[5V7)ADCe:9UL:7Y=C]MfRc=&9S^]e#G>76M6A-LO0Z-U^E/Q>YD7
TF2(P?-,62+WEWcALSJO&\WK7a@S\M<AaZJ2=O:a5;0a8_?AGcd,,Ye4/34++UE7
HQ6&P]-J,#^59_-3GORCU7;TR#aNZ;E031J;eZR43K.,_44D:L3)BG0cVZKR)^0b
3L))._d1=aLF?GK44#gO?8@4E.0H?ZI^Q5Z)V(]:Fe3R+=_[75>b)fQ/RHCYX2eW
@XWb(O7X#F&#)?^)K-Y,e/CN7ff;73G/CJX6[<M?>CY?NC&?S-fW]G1I_WHUCNc@
1C4.E6OO,6U_aO6ZI<MXL-V2/L0a7JC<;@I@_5gTfBBVRCQ1(1):R&HH=P8PZbKW
X)8,BOR_V6K;8f6D;9=cb[BC2<1B-T6F:7W?=V,(]@>\ZB)cHJ;a_?UGV=\F/FaD
\ZQ/bI]c@Sd748JE;OLE].Q&?/XT>dHHC5KKG&#^+1W^BG8Q=/E,>,d42A?L#a6V
aMcb;VM64#Hce<8=g?P7(CK1M)/?J>I@4b?4BS4;f0f50PRTgJ@e000N#5dER#d2
Mg5YFWWCFL.6&f\@5eSL\F1,#^(5?9@:&UbND4YOR6]+\;0N?+--=2DFM+GJ[),/
0+:RGE19b1eO:?\=BJ#H(=;+YJD5de5Q,fM-M-T;/NB.C9]_bL>(IDcB_2Q4KMHT
&\8U4BE<F0#O.IO15R-ME<YIS6R8@DBDZHE[2R-9^:T64</ZD?+c3I47_QL0R6S6
DC#4WgN0(1Q\K@Kb2B4PSV:__#Sb1<6>AR\a#)?<_3[7[=N/]ZS]]G=[7bLEKO8\
\<1E4HT^-Bb>\ARc>@LI=2_)&fC&/HM)2F.4Q&DQSa(ZB[7fSX@J0g+[XJZgE2.\
,f?<JYL&8AMaBLgOV(@=P\P<[G/2b1)\L\g=^G7//;<9a]:^#]=T#eV1K4[)fC/P
_0PP8SfX;T388R,.UWTQ_QKH4:D6K57T<A>_#X->,?T@D,X=DAVS+M@b_:[<&WfF
;,WL5KLRO&a=(+P;UASFJP1PU_eLI?Gf21?>A:Y@<HCO:Y2TIKQ@7J8?_[KQ01.F
2RM\>>ZC(24PSOVf29JUY_&/7\[;(b,?4+TIf@&X-Y;dRMFe71<>/gSR)+8VA-/5
3<R@OOLM63-]f.[6^=fYC3D1@=UZ<AMI8?MTD<B?<TC.GWD<EFX3:YN2b#+Gd8,H
:40>CIT-6LR?ROIIbfKSBISZ?Va\R6JX81RVd/J8=<NX\Oe?0b6dV6NI4C^3,gaD
],8>@C/]LB32FYB15]1N(d,L)2>C71b[J2RH+f^S;fSeEM47g,g[]A?g>#+<44NE
H\<MJ.Vc86Y.C><<;]Q4?e?4;>e8(1L\e6?9,)=XYDNZ=0>G^M.?EE^U5QC#?7cY
gaW6X,YKO7F7De),^1bg0X5+5[BS<a@eL?bEH-\-BMJ/-AW2CL>:,46WOQ(e.GKg
_=0M+GV<4P?D7T:@(:28&(C=Z]<(e<aNaaQQ&;QO005KQ549K^B4=;N8H?/=F22Q
]DMc]AMSbd24])BE6+>dWJb5<ZaE(=IGe#YN4BC-@1X23eg/#d53ZGV2C4X3S:LV
#2=J4^7(Y]UO+#&eWP\(BXTd2ccB+gcV7FQ:PTcZNH2#d<-f=GM@@+Q70c9B+O5a
?Q+6+;<dK4@7RZA/)#DfU^E>P7^RQ1[NQIH:Qa9R\I&N+Y+\WJSc78XYC@a<[XB/
_7eQ<E;,7/7#@X?/f[2Q5/6>V6&G,F.EXZKBOWF;[6MH)I?7eGNJR/WN>3H&J^(f
>+3C__d6g>)IddYL@aVZC[U^,WV@T9L+d)3(K-<\;O(FY#DR,K2&<cA@)UVbc=Z0
bA,e-E)>^gbV_Yd-1#M53^=DPYcB)23-)46&Yf)EO@f6\TF_4,dIFX\_D6:bC\9?
FdW6gLV&;_fc4<ZTLA#0PO=8T:^1#R_E#@LH6_:O6Ue[bZ>5C74T@^7AE##Mg-(C
:2dWLFeY,FN\[TIVO\2be8T7@6G-31+8242.T;M[BRWB-)NO-LR8&IA0)\Ab+U?>
DCRUeXX2-7OUc5T9a&8eX@CWV=fK#1eJe>SU7d0.V5XG8)T@cERg6&2]Gd4;\4<U
PF.1JW1df@_B:(P,SA5gH>Ng3_HW\e,b[=@)F1cXT&>[I#4K:e8Rd89:K@<H#-Pe
/K#b0X]RbU#;+(8c50KT@7@=SCE=__@=f(^>e/JE&<TGFSSR]2-+>.>://5eBf0W
XbW>b<2:TQ=(eJOZE9<96g^ZAO13BD390NO&dS332PSfN:>9GZ[fE28FYd0c7Ub2
3O8@ON2gY642UTO;1UGMZ&-RR#TNX#TPW[TH&JCD;,XV-#T5_?][FN^a^+_@[ZI1
RD.5S\,PX(I_ZAfHX\75:EO&)B;bFXS2;)8G>.YIcdbGfIQW]9DL=?&V/;8E&;:c
\M)MN@cF]##4Y2KHbXK4U;5&>^GV7W37c7V4bYUGY0_>3;3,782[CA#7&5\:HEc)
3]^9ZY<g/0U+]))f3Y8.R7MWYH93ZSHJRCK<Zf1WT^<?.58:AO81=1[bb(cWbMJ=
6;=dF^H5ebB;,UF5LfP5AX2X@NR[LNX#\9I9>&1TZWP)If:Y+OS>XfM]F(>bG<D5
\)\RY7T2TG+KZc@-7Xc=B,_\(Ca2FC]#Z+E;<1WEgF;LAgC&FEO(T3&fA?R83U+.
?NZ><^>\.?<=dR];X(/L5Q^:Bd.W-=48N?L>0L5.[<K[[Q1:P8(&cePQ52g(U0;6
Uf#Y<>PLBII46dRT#JSgY_^@[1^&0OWRQ]>5.e[)Y[g5SX@08K@&&N6^]<+OFBKL
R[MRgCK\(JGC<C1P.d3.be(T8B>7cPdM#fNdX73\+a&;Z#T>XV)\70Ge+/A&;c[(
AXH9#CP3^6DS>&1=Q917,<=0W+Y+:I,fWb:VJCcU4S7RJ4a<:6^X@QWE<VdY,SUO
?((+[(L6FWXfWIZ<a1HXPfSJ=8FIWcfY:B7?1Z),4D2,=YPYebJE1,5)MF@J)WN.
=:PcQ,7[gb.e96?;L_7C/3QRX7Y6_05&FcO\>Se+I[//^Z<\a4ef<1\gKO43FL2\
V^HT\f)CN_O>>UR7bURN/.2(B.H&L(_#L8H0ccS)I\e(ZZ.X&;KdV)UJ^f.gGe.N
C73(,&Y(2G/2O#O^a6C\@6187NRg7XUTZ1P4NDbcN4]4JFcbG(#54QbNe0ZP\gdc
bbG\aC#5-RbYF1]C\1/-X(9e1Qg23)?S_TP<(7(;8-A_#;aX)Jb\O=E(<SMaX=\C
D[_0eOc-PTP4:e?IG\f08.EQW9([b)FUX(PRf)&B/(Q5Y9HADLLJQ&-@@aM9S)[B
cX<)=QI6C;=:5L9\6ARN63^T6JRLP+Yc68SZMB<W8C5;504U&a\(HS:2@_0S_>PW
_]P4)4#S-WBc69&W9c8d>\^-8aFbc?8,IFd4GR_T5HR=d,4g3+D3L?SJ;P>[T;B0
L\F,[-c.6KAYW6D\ARMH<4R4W8V@L[U-\LcEJ:B,YdE==]/<UB=bFcVe7QI+Oc0,
K7.\;T/BAE3R<ZB(WYMUGb:/)GABD]>HK)f:U[=EN^U5HO]bI(aYX\d5]53,,ARb
3SGd\I@RNf?5G8Be7=A&6:^#NTTb=)(/6:RgK]QHKW;HE8I2JI+=2)dSVO857-dD
a+2@E):@:5;DKKX3Ng_6_\d@[F[);fc@gC7bCA.W(CIQf+2AP[C-S>&E9H4NCZN;
a==P^=H++J1L.fdJ[<0J4&K;P29=:6]^R]=#\?P)a@(X_A1,Jc5MC_:FJOQ&P;NG
8gDQN<b_(ZW&d_<.0<K5R5Y43_P=5+2KO#R3[.W9+dLB_EGRFHDGQZQX]bSYUP)?
.K[)S0Pf4\f3KXX1c_bMNaDaZXBFZ?1A.G[;MG-C0;G:J)aFB?;K;eU+CVML=B.X
J;\T>7Y@<4U+aN?eKZPbS.2M8OD,+@V,S#:L_T\:-?5[;[Y+/YYR3@2VTY,#2AM,
DK^aB=d1aFB\Z5_E>=C8Q1d&8dW9fdNAC&[PC(A6Kd>a.RR80=_+RVcFXBa.IedX
g[+74KIQ+R@DaN:H?K:87;b@L2VXXQ+/7M9V<dONdb2Q<2PG:01NU\b,@(bF(-XM
f-PP9IS#Z[@S+HU.XG8+f/cD:Kc#(3336(aP[Ra(4NVb/<8=YZ3L-DeF.XXe1L<9
;N^5cFg79VQ/SZF=BT#O#VAE<[.B@S6,N=(-^NBNRFY1+P^K<1KC2UTc#7?LLbcD
RX?c-V:C@:g0Q\^eFLRQI<ECY</>A6ELR:+GTG)d5-MA7-61MT>KQb=M)Ee<J-P=
@H[??1D,a&b6?LNZ,KBdg>c4ES#eMF_R0VR(IgbWO?A([^P37TD1R3.+<f5HKe+-
8Paf8FV#I]2,NaaZ#Jc=fbcOQJ6R^KTG^)#8(GQ19JXH:VPKb4IH5fO;F:^AZP7]
UUF9Y4/?<;=#Ef^CLd>MWa-.]L&.LIJ)J.Sc7/7)JW5J4WRG&_F4#Z9/a[S;6Gb>
N9(+-S(7(gO87PTY;<4c9VSdGeR:LfS]88_fP49D[5?)a>^gEA7\VNQ-4UY,FLS-
D#8JSb4,^H&M/-2/bX)<(@H=9e3S>P5CSU+GZ?a-K51ESP]8J3Y5d1eK+:aFIe-^
IQEPAEBGfeC72eId-J2[1704=16-0bC6&W+<N]]Q&_RM>;EGN94W:LNRU7Zf(D36
=0>f&FHGO<H=Z6G:TgSaBWe+&8U^S1T3;1IT472)fVPN1^03(/2[M;28d0.N;]E4
DDeDaRd]:ZJVb6[bB07U5f@Z(-X&cNdA,@5N3G\[ZYIPb&KZV#b7\RJc4T9a.=0T
MHIc3db@U>YQM8Sa)fKM3#NMaZI:+5KJfFdSZ8HW@HL>ab9e[cW;50/Sd-L42RV5
c/(&/M1]?bD>JB8U)aV>HY+D0a-T5;+Ng,8cUZKL[_\N;DbIEZU7<J(a@PfMc(I_
^<2K02JKf2N&_QHY04^7#OD4OL<<O.cDKE.Y,\5VAF]^2)G^6f.(IF<19FKE/,86
e@45TJfg:,ZRVQY2?JJ=a3&;0VgX[c4.+UWc.Y8WeV.6(]&9K0ZXB,U4Ub3XGO_.
c7DP+WfXaUU(::4gJbM\=N<W@Y:1G\48;W>YV+FD1)B.FNZEc:b3OC5(GS;(Nc-2
2K4e1C^.Ic,QB76Q,@dEPP-SCXIg<C=S[BRaREXXNZ-6g;]e+H6Ff8>7X,N57dX[
)4BZWHF;PQ6AW]WHKb[TE:7HE+\LDI_2H/:)^g],d?5_S/TS1,>=Kff#3e5\G+YH
eJL<^A=Vd,d<eDfFC;-S8GZ[Nc=O8JT6LE\Q;.Y<#J^IfD>FB)>[((]GZ=f\RFN=
38TBZ&MHMR+Xc.b1c6ES,SadX(+:^H60/8=&G?T&NT\)c&ATSKALc#+UEGeY_SAK
4XKAd&)5_RP>N)^S8a?e+#<R3gLZD,D\NWQJUC;f,@NFe-bHL39MP3]8ALH:LD2^
\Y?fAOQ-[ZB[,JRbg<gC+AH2;W1UA;8/G^=P=F5#a_V\LQg[d6cC<@^:<&(-DX&H
]Ge,_I)ZGa)6O/@X>Gd,0]N+36(e;RZ\O49@[\/A9-Pc0G@>--caObCS=J>dF:HI
2TNJ)U47+&T4JB:O@?5QHDQVXZMHK6,X>c1?BBZ^.LNL>-K6Da@b+[aa0beH-7&;
8CS8\-Z=CTNW\VX@3WcB_JReEBM2eYD#J;]SMdXYJE<T_#4#>:XaL(=_c_S.]]E]
RSV(0\9UFCH02f@U)ScNfU)WTEf:-^C[a1^0&&;6Lc;a<S@S&TSYY[g4@M^54;.9
)M\<5b@6[GL#4E_FaY:acTCQ<V3]C5@?:#dP5f.33TG]^QgQ?P5[E=S]C@VX?8#V
PS=g.BV,,R<4:(?\<[Mg/^)_3VNQ]GbcfA(P2/-T8NEGdE[+-#QN@<(a^4[147bA
IYbccV33YD;R^6.KI7FM74KbH+(W(RGN&e+DKLUKE8Jd)=eDIM4E<L+\DU\?b&.V
TN\][LOWe\A4PS(]Q-IDgUNRD-,:1?.4^-GI5<FIN9f1=]A<M7N0Z7?),_SSUf6g
BG<@/aU:a@RO8c.ffIEZE&1T-2SMNf66.I8b?64O?]d4Z6D,g8\Y&Q^&(+Vcc6+F
0Y6H=-B6Bc]F&\eDQKd=,J][<85]W,@VGTP-[EY;e).82Ag&EgM7C.e#?TcMK9X2
V]U8Z@=BbF/F_F_I47(:)L29,P/9THVYT322(RGSKM<dc)D?C-WV]=\XLDN5T,gd
5_0@.WU\2_S67I_XI4V5I=>P.gc/>J]I4B(SC5/cIgbGH>RI27>Q8+0@B/5gE9L7
7;&IKN0Q:LHM9KVJZ9LG2=,?<2NNZe((+F,S#,N(\;cHC.;]:5,[-Q\SZS)Ya&U\
6.Hd.WWMG:?:?F9VD0=LbH&^^?O]_=aA-([[^E)^cUM<4@-@dd-OWI@gILebOKZ^
D7^.cHbI\Y+74963dR8e2:+AH,+c.:E4c#\JPI>][P/U)LAgWa;GYDV3P,WEU]dF
6/_&KG/,<V3.RXH_DHJ,,VG7I53B2<?J:+g?b<4EQ+6\&?AE_V1K]Se9e)(b_CJ_
AX=5H,g/SX\4VZf3N/dc(@OFW[39T67],/Na&_LEBEAFDWRb-;P0fL-W&S>+_][d
[Yc+Sbf;.?6CbON<E8IBP0,\(>P1>)11/f;BKU@g3]dT9IP8:>[+IfK66cY.;+=S
E)8D4NB.LGL=46RcV577bBC2;G_(YT/aE]:3MYJHL)#\CV&;=g],eQG6>UDH6eJa
]aP\N/d8bY;QC_]OI[dUP1S6@D0(JG6PIe.(,,AI&9?[.7^OK1bFA6IU7]M=ZGW#
ZP6))ffL7>dZ)@XYP.O+5e[\33_SXL[RZG:G;HdFC0#H(F_+QNM8^R-N@IbdD>KX
PaE6cC7G:JKdX_cHF8aH38/8Ng5^9:d?6+QfC:3F08gM7N=M/c]A\<Ib)[Ud07_O
5+A\f82IHS-cHO#bV#cJWVC(^8@;F9Q+^W9>gS..4KUFf[<?a,S)XI\ZVB[98JQF
7J@c\QPNO/0)@/4N:efP>@GEedJ@O2_#,7e>5YG3/L0dbQJ6D)H(I7_T]Z;_H/bX
V)(D1\0\NOX0:Mf[@DNF#64fI>4+RS^3+d1KI<Q)^8;60=.Vf_SgY,0,BAY&&\(d
K.MK&T/B=aS_c.T=@1O[H&7;Q(V3A616e:.Ig5ISY::8Rb,_=B]\R;2.f1>,XLCH
V@./]I_1C^3P6YS-C5Q^.Kff_;b1A-/+MV8L-I1_ed[JB\EFA8WaQ;\]f6RN+8(N
UVdTOE(ZcKM[V=T67@1aGT7bbCQ_[-L.DG0bOO09;4A#WdDD^IY]U/F+fP,A+d,P
J]CF4L+L\J3D:FMSD4Z6TH-dMZf]2GX9MJ.G,@Q5/)08/#[P4(VVaf@9]@KbFR1O
4E\Md/(HCV6N.L0HK.eZYUQME(JLQ-<D^G?6MHY>NIdTb,Y>Ca6S_,?MUQeEQHa-
VR7]ON0?PU2N7VI8f.]<,?^M\_N;,.3\.(^ZSME/]X-^BR9b<PEOE[8VfH=QR4>7
ea?I;I<55>V7b=4)(.Feg9^))[?7W4/J>UW2ZbQ.bDf4#4L2>_+Z6H,GRXOY)SME
Q,3X4RTead7#8g,.T:_+CY7GV8CBWgb6:W<#^AVSU,JBT<:HgC9C<_ZNY;8^)^9^
5@bA^=^61(2P3A6YP.PQ\ZaKYZ[F&G-(2)ILgB@fg,44,;=c(:5[RIa;3CO?<D)A
F@):JG>S[GD2b=3,8Q>bLWA&\3M?FA40B\K,O>(048EO8[E<>&8<(M]/+LUTN8@H
3/b5]@L\&b]cdAYfQZ<?J\MX\\6b@;:)]^/H,Z1=-7cgED:P5BQ-5PJBNCS_g?Ka
L9-K\dQBPJb60)=1JYGK,A0;MDCd\.M,AB9F7HUKI\3AJ,/)ddAY:<gKVNM;27IP
JP4-H]_+g7TC/>G=5f]0@fcC1fI.^Ae&EX-/;/@ZNN@X-4fAP-4IgTIH=QI^40Q#
e_K_0c:49IK;KDO#]Y1W_5,W_LY=H\SG/da_XFHd)S=>(a<5@d(KMUX[<DP0=/ED
(RT:_T)NT4M_ZC4f(]]5I30K_Q1+C[C)KeX;Od4NXUTA/\WH/2&UU1//68K,#/ZG
M8e3J/T:0)S4+c0eFd/B:7Z>OWZWJ+L4PZ(c?;W&AQKeH8ETDBEaW7O[<-Q/d,U,
&=W5B;JMHUdNNYVb3V#Q;M5VKNa]Ke5L,CcQN<IcY]de_4NP\?3a[S(c]4JMVNX9
-1Y+C28]N=>FJ]V8Yf99=dCS@Hb2OY3)J[0Y(9)/8Z-Yd<H/2I0gWKePbBa>#F84
fJbX5;#c[HaOb>Ta4=HfK395c>4M<_I138MTKJQ;?F7ICb1^QU_R)K^H1G[XN]95
@KMG.a,RK@Y&TJ,aWQ5^KNe_/)eB\>]gfg0;TRg>3G56IIJN(fI/X;(>W,H[/JI4
;JRF,TM##=5L<PG8XEM39b;XdA.>3ZVDUK#/-.727(C./gc:7Y&Q860<Sa9?#1,b
b-DY:[M[P#Ge+gMJIb/@]e:g?G23Cb;04#b0A=O9P<9<71N6-C2_2M>Vg&fH1b:]
]>@-/]E7cI1da??3]C=:&S]bBBWAcSPA,RMQLN;&N,fX/LZ>/<VP2=c\CcCW4gZX
M)T-^J(>8Cd<)CMLcBM],\MegYNNA?ANKTS&dU9]Va-R-fK[>_5DTdYbH?R:0ZV(
=N_P:MEKW1-eHRb(Hc^f63^5P)#56,:-gIfRGGTcK\N?8RN9DL8B=S;c9ZHIJ@0W
7c^,E0]EV+FGeN]RW)2:[Q8).#09;+4g9P?OfX9I?CaS&IC<VHV^W[TWeKJY)]D@
6M]S#aDA<a7Y78C:eG9]#1,:8YU#@9Q;[W&<b]H(fG3=d33&FQMF25RgS1QN<:8A
d)PHR@],W2(4c.>3LDC)\80):=B;A)IUIC_-@.d)b((V)XT5LV:@a?<\F^\3N9BU
E+&>T?/F.Z5B<3RS&PC>^S]@d.;V2TQ;(8eagI^#a6N8:WVgILU1>EGcXg^V[Y,c
XWJ^\1\M3BL-LV165X)a8ORUKeHX[7=;A84]096>M]g#=S;[ZY^URY38M2UY_++Q
;O.Q=Uf7fB;JX6dV>fWdLX4ISL[>B5\9f3E#ZQ4W,/@,W[@]\d;44PG8IAc6=FXM
M@)LF3\K;(;W1dLcHd:+afeUg@G7.>c/3Q;bQ8GN4GeJ.@gK\^92c+BU[+VG19,&
,IL1CNb\(,Fg)7+P.2PWfC1#MQ&@N4BF_T\aWS;\,U04WG:-.FD\<6@T/F]Za^0_
.Bf01)F4SL)U>.7c3Jdd>B928c=6)5=[=;LS@YHed_1\G1PJ\a7bMGS:HZ/PM&#6
_DHBgNK_IW+#Oe/3XF8?G6T=ZaXfLH<a>^79T)?^(Z+fJXd[X=.;#_21R/Qf=f\X
(;ZOc@++e;T(JWK;=E)Q8V)M^]_MAcQGNc<K#D>]fNGYB5(J2cD;cN\\,,BG#D8d
0?4=dPRg696#cPc9N1P#5F:Ra)8Dd=&JO^6O>6&8YS\#:Q<-EPWNX@)UG).cE=K8
R,3QDYBcVJ)7L,Fd()1)EE[=BgI:Jg#1OS1@C^4\L-;0()HQ8P-./:OVW]><aH-W
,N_)37KRFY][L_6R&+0^+Nd>VV+O3QKg8&/:/.;?GMSP^:RT.68F:X#R^bF=@.R?
dX8FGbTfZ=_>5W[RDK#cSB62C.?..>473W#T40c,83eaZV,3.&gZZ7SQE2?b/4Gd
FGbFO.X0DIDEE+7GN9bb-E=f8EW<XXK.576KM:5UfN088CB9H[I(2Hb?&e(<#a4@
X.bDZ_D[?^,RZWL[#1LRNTMe/QT\UWP=CQUM^aUZ8_0]@:.09A179):d&I=&KdC7
XFQRE#c3Z5Z>2<503cH>g7d5S(3_;<E0+G,#Xe\/e]g.b._f(c(c<1@ag9b5/(Pf
22<8J&ME1M9+AgZdB98(8DZ\9FOf1E.6DG[FYT:_cYL]M1;AU+3-f.9A,Q/;Q1AY
4J_e/-RfBBGLQ<dW<R;0ENYf0#4A)Y:&440)RP:)CX_64dGDTD[W2]X/F8eV^#W8
QYdeW9OeJRQ7OQ]QYV(M,I)1[RFg-L:#eZf3#KYT/BQ&U4T8#^=c>N&H>D7/6TA^
Cc4P/#P<F@XFI1G5)=?W&g6a0+WNC2eaS\8K+WA6dbVcGbM<TYW<GVULf[]YNPXD
8(1LffgP-7P-,6)PARO2QQfSg(^Tf1>T8DUQ6dcC94]Q@YMQc\^dN9[U27f,;:BF
3V-aZfKQFR_Vg/5ML0GZ5TO\MM?)K@T>+?;O-b\5_2&@Zd?<VCU)ZV.[@>&<O,HK
ZVN1ES0SJa<f4KFY/&7YQ54D>,TNMW>I:TA>6Zg0FaWP^\A5(C6NXJ]0cSf)IbEa
7@NEKb0?_Re1DF111:@a0=(SC?JB.JH&V.1N0F#XUa6_R79-fPWC8U;V6=M8E:/4
[L448JgT;.B@Qge\X&G+PR?,9CaUYeD]PN@ZWI9V<45M-:.GQfVC(VS&99X)=GDH
2XI_>7]e@PNTF4Nb\Zb2#N9)(SJIW).LS-CJ79>>>-Y>fOT9Ic(#?4Tg@FLRIDLU
c[f76Bd8a0&(gYS_;AL9ObBQFe-.]LK1;?0.>A&c4=O3-8<H[dRL?5YAJDK?]5DY
-(b<\+==XL./e0:>:.UA?D5=g?SNN<>RW0dQFeH(8PN]Z/3@AQJ9B?M_A_L<dN-Z
.8d/Ac,77>3NUC;]\3-021=;NadV&Ue>@=5-8#EBdg6[e)b=JNJ-=3AB)0L#UFYA
UI4IQdQ:FFf/J\>,)74,[F+O-_cR58+&-/+<-VMVWV[aIW_J;YSIgMf^Kd;LYfad
N^@0b@Qd_T_=_=V^:6B<Mfa]fIN?9a_HO]@Q>?2GBIL+9<_2&Z^>\e2g+g-XXA_+
M^K6=6/&2,BKRW[16[3g3HSH9RUeLZD)ZZ1.#T4=4P7T#JP.28H<NU52PB+\Sf2W
ec[DNMa#IaSGFD&2Y#Y9?_c3H&Kc>;B=[C^\EX:cd-?Sb7cVf\ND4@RHKHc0\/YS
XEL[g#Ab\0gAe@3+Z+EJDRdV3J@98@FCC@^5K=<O(aTGK@H6L@MK@SWPaeR8)<_>
bK^JaIcKABTD/c<FHZLf>NLBDRb<cN>(-])6Sb4Nbb_]aO+<J.->g9#5T#I(@=DD
?A7=H.>-2Rf=84-F5=XRU+NL&#X2:e)a2.L3)&PaZOA@B^Ya>^fR.N46^5g>\>AD
DgH=,XbC_T7TGLPRO1@:Bb)7I2bQMDZZ#9[FO[b(dV<aD3S.W,1VU]\#Xg41+>D?
L8)1+Z&Ma2F;BX.:eB-;bQdIE-;FF1WD08GA+3XeO3VEFLcfC\:^Cd,\\bbb+Y)\
dg0Rea7C3N_Zee]A;S,5#.VSD3--A_Jc(BZ(.FD-X.SB\Kf@5)>\3^U2/LXdD,D_
@@bed=E;A6eNaOW+J1DFeV4-J;@]B<M+<Fb@G(UYWf9P4=g@S_=LMR4a/5MDe-<P
XWHe@?bRI^@]7^LKEgZ0DM:f^E.T=?0Fg^(],,dJLFca,ARdL7OS)\dB?Y.=@1Kd
a9_GE9UX4\Q[e@0OI0ZB/0M,.&\@9Zf\]O\AR?[WX+c#XGD[d,_31bA,KJc]dU?g
QASN,0-[@\AM94/.C\O#1a5]L>:Jb5:6NHH74_\F?B>NO.2a[H/\[d>/[a5F0O9A
]5+1d>XX4eI20KO,WJP=5Fdg@KgeEeIEZ.a5IPB(\M_[S95U.^de]?4GREW#_^fc
7aRAaa&WGd4gY35+cab1EeA?BR@f6:MY#4@,E9&cBa>HN-<g-R4MB4=(E(HR5Q0E
\<7.,[eIb,7d(\FQ(+F\Y=2.C,7[P]3;fFVZWFTT4[B?CaDD</T;F\IRa1B0,EQ>
U^/4=,?L3F.#Y?D()?,0,>2Sd-2.aRWUBA7[S4X/Rgb>8S@)8W-)/>0;(e\fX\Bg
06/^#c+&->:gX(W/XgE:17B@UQ[^#L5EXI;YGE<]d<39)K,1#Q;1WQRMOSLB=;#8
EM1H;XPa:8XLcP-P]3Bg,X:d>cZ.Y2b;82HED4@.5?V__4O?DG\ObdNXPZG<XL]/
K8Ob_AY7dU9Wd9F&&XRBJFa3>&6SUUB@5N/+-g;5\eTb[W4630+VWY@RU3Z3[X_@
87,OL#Y[-d?#Y>_0@^_3VGca5SbC@1J74<;^IJ9;KD7b<NGcf+0dYaC8P4ZO+U\C
9KV[/c,KPWCeC.Kc8>KXOdKF@B0fg92g9QgN>^,VC0U3ZR:MB+#>fC7d?b67FXBg
eb/&Y>RF)9.<^eLC;SOI,>[?Pf6CO2U[(JE7,X97-Q]OP,c+5@P3,<Qe&4@4I\WS
>NFNN]&[(>R47a9?5(f.++=Q-Z<\92-bMK_#35eL^3@<N&K0-Z6@J-Ede^]HN#@g
d:BZ<A&B3fWG=bGZKD6KVY0,P04FTJ^..I>[OCZV4gfA6U:SH#Q^RaCfO2gBY_a6
SP1g>?b/[>YML.1H(1_^^Qf7BYN#F]A;F=GE2@f+]=.//=?bG3]=e0^J<Q2?#gL_
LLJ@4AUfOWH2@,WI2,E(LfP];de_Z\7_(B3#P4QaKOLC+W=F)U2#_#aM=O#@P)<@
I^<&dfcDS=_De2(gDaH;N17aeUN.PLGH?WMV5H6[[2=0CGc8U<6YAZ&H#-_)^cM5
b0g[^@K3_MN=[/)K3_&:)Bf&M<F;]_\b;_#T0#g(XeJK[G?^eV=1fF=d-],[)TS0
F4^2<5cWBW[B+UE.=0bP&NcJ#><aa?(]-,BMRg:&9=eD(-e5@d;7W)E#9dL1S@MF
&XORR4J;>W_IW=U<J6cC7c+O##[Z+fH9>:CS<DOHSZcU/XM9K/&[,6\>d^A]VXT7
/SgSB1\d)NL51#5[YU.@W+@fd#SbUETME(J>D+bJ_g0K4?RfJ6:_[1X>;VC6_&1f
11?U)C,UP)gFEbI4D]E)0&Z4gK6R2W6aILF8.F:;bQN6RY-cf0#96d59Y3.47^##
K-8VPa-,MI&Ne6^D=ZK5c@G2^#d)S[R6ND<2O^U&ISPA7L@S#PB/=_X(SNF=fJ8L
aM53NRK0HYG@XSMPeVc&&JDa7X3W/f\_4Q+[:O\He98_e.HP3\MdbLY/H&VBc>W(
PZ48MYQE6+e+K>51\b/W-Fg;X?+)]G>4JB>GN5:Mc3\987A;/)@fE]D9XcDFKf#L
>BCW):QF1>]c+TH9#?R1H?V#4(91?P?HP5[\AFJT.P?-]3FdC2_[[0ZD7_gP/dZ,
R+;^bHBBX_YQDfZBKL>+TJFeSE[D-gF^E?;9LF_&g==I<9e?;OBB;cK6]LA?b]XH
,Y&:ZKN<Ub4()U&E?[2X4NDC8S&e#e,?R<@G2ZXXdJ\a?:(AE#25[L_XIL^H0Z1U
GI;X1&STBeZ.AU7[V?R5RNgNRH4fSL86[NE5AJIUCN^ZI6D15MG>K@JUb]IF8)e#
?M)D_:;K/C()6b-IT9WE6N^53a1O96CB5)8/5MOP:AQ\YW85BX7C,CaS@V[(b-D\
P2CX..@V^7L_f[LXL8NL^#>bO]e&d_F&SK.QH^?]N,\+bAX[:f3JA9@H\9#I7H\f
U2Qb7?ITZ.@.5DPF]#[Q+N+A<-V(35g8>d?8--.K3Z=_N\[(\6M:_<BPTE,?V\]^
Z.PKIb4G20OA<^N7;gB<O#?bDGK-#QdJIQ?&KSJLLJgT-DQA^ddMTWebAc3:Y0_P
-H.CC<cI]b>])>.c6g@?4I<OW-?R=2\UHBX:4C97V]BY&BE;B+>[cebKf#U[gS?e
QMg2&N<a7O_^=DY<XI+)G#R&_0]W3(f7eSNI_4Lea:#2Q[E&[)X3>Q#QdT/>I#_U
Kc-DAYU^c)[Vb<C/Ee[Z[R:M-UC14CW]+E?23;[OC)#;ISGE3L_INY:2<-BSTZF9
SN.:8fY?.FNf1K\eVe>>a5c.GdMA[\,&gX35FDN+:<V&^;R-[S;AK4=TU]RCWEN6
U(N(JGC,TF)[Q_11NMf@L;8AR>/^WZWbWG5=U=gVQQ<)3LS?@^#M:NA<P<cUAaO=
HaLBDP0W_3^&HC.(B/EQTNB\<\.UQFf0,L;XRggc-:=EE^ge-\.77&;[f\-R^9F>
EN830@T;EO38WKV2XN</4>R&(CO(P#1E(&f\91g80Rb&&,8&XP51P]bOf7&&Y.OJ
[Y).(J-BJcb9A@-OS]96VQ4()WYacXge2??-0TC#>+;6&Y\f&V_.]:X[1O--GJJE
DN]cB5BX.9SHXY[M/O&aPaNW;bA1Qa\.(Q[F60D3c>]ee4V:Z@._V0TA>-[U\:0f
cH9F\?]WUH&?H)@\]CP^_c/4U-2,3(VH74)W<MEcN7GT?PMIW#03I+\)WJ8]ZP,G
N,./PN(-=+&@K\V=d357eNEZ&c/27>Rb.D>b/gYP^0L;-K#[S>50^&gN2INgU.Q.
3VH7N)ZEHP^_@8=CCOb?L)f.1ObH&T)V>JJ7<QYF9P<UE[:&D;YGc/<9T[HTcOZ^
dPTD^cHE3#<D:b:#\P/bfF](NPY=W)Nf7I-B]BXWKOO_a>JH),MOXNO8+N<KI2PT
NO2^HQc@C]48S&Z3\/a0LS:4=cE757J4X;>-9d6N,X?1:1d-F?=LB]]NXUO0HFAP
RLSVRa9/PFb:YJGQ^:RO6KRIU,BO]d<#bcM.JIP(HBICZ8C>TLY[5IT[f9C:2H,e
E7,4Y9d[Mb>->b-YLWIJIS<G5+\=B7Q4_;5eU]YD0N\[d_#;23KcCXSC05>R[OF\
8e;bJDaZHHV(\>2)5)U<Y;/d2?=:1[DC<9T^A^@FdH1=gQg<X<1JM2=]N[:;/<,4
aN3f4TQg;,#RE4MQ?c[W\-=R(bLU4W4_&)HZNJHcaBVJgF#_=.W^MdU5Q)4PIFI/
.5OB#&2<IHE1bQN,YDe30_d^\]TZ/HJWXPU(ONDf)J.NR>0BSRd^0b_5@C&=eb\2
Vc@#cA#,#]78NbDZE1ZQ\-]?=XZf3b=R6T.XRW97dV99J_Uf5Y]GOSMT>2g].Z/P
f4JF2F:]eQO#e,d&N]EB_3L?RN8NMIE<b(MHdZ<X:AC^Qg]GBWHL]>@ZTF_F<A<?
1G+3&b?/geCWg3eGeaO<>?@Y939_T(WSBN9\;fR-]SX7,M.@]9?2Ae8=8dQRVaV4
HS.HDI(N?5K<D4<.0eXYX0L,.+BJ@B_]aS07J[H9\C3FDK=/[3Q&YC?EXgaOU>(]
W\:@fUPbIB0KO\YBC0a0?+XE/+A&W(MI0IU\2:GIFM2ZAYFd&aLMQ&SgI3]fC;JO
R]NXZMeMA6bfAIIQSb_[LReL)GS>X8H99]X)]Ud8c@^8;+MUBCF6AB6ga7WW<f/W
VUUCR_gTeaU5(feTZeUCE(4@=T?b;eb_Vb;5VL3DFF>DM36d+Ia)OIZYB[4FNVG9
bO2aISeR)UK7bZ\-dH9e9<Ug.S@;_3a[S+V]H&]B:c\JbK-7;)^UL&Xe9#:4_##?
2-_dA_#-6&)\5Fb[):XG-EXYVK+7@f_VK?;\FeJQ)(6GJK#BQ;J[>?Kg#31,Q)#M
#:?^Ue2Sb@@\QA/#f\1LA=^-@aQB(T7+fgRfW(6G?<-eA[C^\2LP8<;87>,04?M<
7WJ9+[V;7+-CN96Z1?&MIO?Y8?Z:I)Y\I3NVVU:7^[(2&(fEHU(8P3I0GJNT)gcF
=\9&Z2QT4<&CAJ#&DQ2EU?OMU8c/K0[0IJP6W?<R4I(#YP.)8<Df\H[fTcWdC1OI
H6+P^cV(7)?<AMH_I([RCaLBH3M5?@7I)1IQOZAZ-L]a#CO,75VZ@LOR8aLJN+XX
bZaL5eU-.KF+I&5@fBRR4&E_X\LNUaYS&FSZ:_&(=d<,OG1e=W(UR?9_EaYB[dJ,
.R=H>0c+\Z[4dHX1)6WMe-[#C4B4<MKd-[RD2=_MdK)436[ae?bdCF8?<P[(\3&[
)H.L^IYVXZ-56ged<+D[-@X@UJ@RYdH89DG)LU>LHN]7[\<R=VH4^144HGeA:S/[
fb:g\.G1[WITJ,/cX>/,_8A+IS9A:/,?LC0fX<8H)8DHJ8TYWASQAd3eBZ;=.6B)
Z^I5EdW6&/aa4^]F._X-P_6S_)4/&Qc0BTRP??2G1VEZ1d[=DH8Ac@d3.C/Ob,<P
TgLJa/VI&[_.8ZR3TWA7V+TW&cW:Y#GV<R2-SBG3HX^.B0?[AX<+O13;ICFeS]TV
>\RY/4IVRAS,Z]C7Y#^XB5FD.MR&9=_,1EQeP6/05\;<Z0B\cA9Gd.T-6I/ZbC=K
WX7feDJ^Fg/ANR,gPd^Q5g4=X(^H^=eR[c28M9=YXS\dg,,b8O8K\NgJ&3ZKC79_
Q^1BGI91R=R/IWb9CD^U<_ZJNeJOUZdQ6W.2ZU>GP?.Z05]XR2@;EE[M)#YI\F=-
9G0aC1KV\#9Sf08AVY4YVSWbQb=H@9Qf8(+.GK4^3BO^;USRC5Lg&(U:B.>\e)]0
-aI>08:<=?WS:;=6U6:K6S;))GGd:62=U5>9.7,F&?]::14d.H\YNNN8+DEA=^/^
HbJJ4CDdUZ[g8GRHL<8+IO)XXMcU;-(H:C_c@9>XX/1LACMYTDeO#F^UIYQSJIXR
ZIITc:MO\9.&RgIMdMNYE#?/Y4#Qa.Z0C@bSa2\/dB3g.>)@L6cQBZJIX:BT3E9Z
XM)COYfHHLKN2[@4<A04/IS8CGMCK#f+;S\5NCNW(Ue5RX3@?<Y8\_UJD/(cB08g
>Kf4[NUPZ-b5Y7)V;\ZPeG39201[3N>RDa8e#+-W91=>./2?HGYL9fbW;RMO998_
.c^CH79e^Ga-QJGFQ76PcSHMgYOB=6/)cV4JBeJ.K-TRWP+<Y58K?H\8fS8?D]NK
),,M&1fYO)>Pgf2T5?&.Sa=0)P:H=G+d>V-WJQgag16G(-;;4Z46Q7C::;D)3:)9
MFTdeVG)9WCRXWV#CT7d>Ga[f]QaAHH>Fd2P4U/(T/_&>.0XG]DJ.6T;1](B+:Jf
<6<6<4efA<Jd#eGZAGaPQ(e5Z:ge)1Y=U-EXFBa_:V)S7PDc,2gbN=0>#MdMX?ZW
5HE,BFO7J/&.]9)7&O#Z:VH4g2Y)?/Q@Gd52Q[::,E#d&6/6X:E,d]dH02gdA)7O
QQ)MNdI\g-4f_IKB,@ONQ2U7fA4/889;IF)Fe16P,XIX#PAYadQ@P0f@;_5[V(CN
g[?/@@<deK&T72d.c>15:L&e.R[9;<-Mb+&\7>PA^767S,PIUY;UJO74?)9,I:?0
I_OV0Zc1,RUB<.d3CcEg2.UKJ;J:W.^+0](cS,W8I?(WI0cK&g<-:(:MJDMQ)XPX
XJg\>F@6+=cI+.bcd1#2L6E6bTN#X>WY&N;d2>aP3cZ2>Ha>eIYWNK-YWLdRWP)+
cDM+=-a+-^R_IIN/bE)M&UKQ/VWKP0Y;.?V?f3EAQD)N9K[4#GgM#2V#0T.9c/K<
W=8_>GJ8SH56O.LF,eSP@_f[WWQa.6cUW+W6;cCbMP&PDcbZU>U6Ya[B,2_&-]W[
RP&9-L5f;9-(+#D;AZ+JBLIUbMO#Y66&aP8BQ17f0)>L0SZ,LDXU6cKN]9+/:Mb#
#RcGC_2c@DUK@11&.&bG1</)Pb.bdC:V<0\_#6B_?_/72>DS43cd,L.#[-(V9NL?
N@HUO=8dP:9DJM=QTc&0<>1]WA<G-OJYM9V0.6\MFDCF9SN]M]CQH.]d6J9f=ANR
8BdK2BIK+^10e^SS0^L9eb8gf3FWa>UfZ&Z_TZ,UWVL(=Rd2L7:#GNf75g[<M9+U
C-AZI8;=gbYeEHK&EA#E18F#cU/VS3F6Q@WL@,QHcTE-G.I?:?bAa8SMa)OY=OCa
)>U;Mc//TOR[?I3IAf?#=XPQ[0Z-gV/<b8H-6NHOcfKYX(K))T_&PO0_a054//.K
_NKFB<]0,2e3dc[TY=#28SJGO]M/_U2[d1L.TM[2M_S,(-dG9VSUY-BFgG:AI_H]
IAgf3BA6Qe8MK\0@G]\LC-97eBB2=@,^N5LC)fDC8[7WBI3<;R5HPg6P:-G+F/+=
;?Ac2V,;)KE(7_>Fc@:0WJNBWT__#;5IZY@,5#3IfbYI._d4>\XIU1&O[ZHLQ^W6
4B15;X9A:92/Y+>^<.<SI,]b@:L#K<0NF_AU#+T7DJa.4KeeY1HO4Q99JdZOEW[e
R6\PP1EQcOCR?<NS0]KX,QB(_W)#G^_ScSfH1(?B@H&)GOcV66g,g.P)P]H.0Jd5
LQ8KI_:e?0Y69#D+B4:3S>A+AHR.E;-<E(C:g[[a6Nf(1XZDKE#BXKf>8S&?FD,K
/0e/[^He4?69B@ebKGA8D7^\->NaI),5XN?+gFJYY9&GQ=_I>])cXfdRHM[8)Xad
L>8&VX--eHI><6ad2=(-SVgdB1AL</2^-G&ZXaMeYCFe7,^\fF:((L+aX^&;N@.J
WCFS=Gd(:SEf\-).?;d:DYJ;,O]W6@=.K/QN<bJf>I>T<I8\98^E(W<QX6A&aVIK
(EJL]_2O_a<XD?\CXX2,7gMA\1;G#a1P&V6JJW;MS&)F_f_.M]B_9ZSCTU0],7.Z
dO2bH=_CeMI@>&>OW>A]fYS,+<R1VOJAeO5\];Bgfcf[+(J9c+Ud@U_05DJYZ\Y5
R]LW7[2gSNJ;(Ee:V-6T6UU<4LaRIeT<fA7]4-bIQ#4HMZE>?/+X,YKG<CeMJI]f
<NgCaB^M)6ER)^ZfZRd/^^.IIIRML\ZbMfd6H?].PgFPeH)S7-[8(Tf[A85SZ-FR
7:SZ#Jd;T/>N22Z[beX\>:R7B\M,Y2T/#+04f-YeCK:;[K^@^1\<XD2]QM:,=U[>
ZQR7)<a&RC,#U6UWQ_9:60>^1B1NPT?DL9R?9D;Z<;<Y?a.O^D2G\74LA_(?XY)8
?X(HC\^T8]LI4C5b]YO+_(L0ga4dGP[S5/Z1T[1EADIJX2\;5L[2IK?UfDC5(B7-
P44J0#@#7ARYP+U7HHaIK@dL38.USd3,R:VZ?HL=E@NFX_D^f9;_H4KB6Og8PQ>?
1TB6[&4O]<IaKH6S=3BOdZ1IHF,]CJe@OGY^11e(/.eK:>KX4J-HL#XF7>/^HY,C
EKG=M_;fKY_].\&SPR&QLT?2f=HM/G@[^WU@)g_O+3;]M>C2fFa86PQLe8e-7&+\
SgWde#4CaC.^/FJ11F&#Q9R[5G3X?S,H-0K:\T9[M2?GW1Q64AU7O4XD:;fX_PR>
d^UPOA<Z<_5MYJBH1CD_[bWWN+]gb6A?)=3W-8@?(N0.1K2^VB+5FcHCFH2\Wa56
-W>,40#_4J3B#YDV#XNgCXHgg/LVe:(C=c1:WHfMQ95C3O^SE0?EC2@<1(:Y[S.W
=TeLMH<V235UgXP]:-_BO>Ka)d1AR.a293R-P661[UA-GZ-H=4[2F1RQ@K(_f15A
)Q_;:][SL<N2g)5QWFZReUP&8f7c6PS\<OGHNccB<Zd-.JS67N5+U.Gg=3G/eOQ0
1d#B4FZ70>A-F(c_;6<JQPca)D3K[QMOK2L^XF<98-BX^e@A-.QRUSE3XY@M6(.U
-<?UVM.+O(YPE+6Xad1]XO6>K80[D-&?G6S<3D-eJK-QR?9DQKS+9L/6bCF9_7[8
0ZOeTY4LV&O>2<,]R74[/4]28^Hc]2VR=?Gf[H09[>GdbB3R#R?0DG^X7P2\<2G/
&,VAOJ8#Y;(NMc8,9=1F,4W9O5e8,IA?,ZA^]Z<8Td+UKAQ):^&]d]35]AFBI[N3
U]?X95([eJW(#.80)&<?XLV)SE;3C4(E3c<15@5IGRDVUL(HD#FdPZUZPO:DJ+WS
dR_.4IdC\,M8#?_W?BIE)Eg)gdHE-A<([B[FL?/Lab[d3H21F,e.AVV.3,]UH#b)
)#[Z0-;/IB=ca+Nc_>8F69XJWg][Q)c98GINfYS97Q?G,SGN&c=9FR1bR0:C&-bU
>Q3H#LP6^.NER#?>K7g&[IIPT6+;[eP5=WX+BPLLfF[0GPCA<1F8[=Z@Hd2WREHe
NYLc:UF_LJA1\_eLEd#+(-V@B.)B?U^Q&]8K<0U[F8-N,d+9Q+6[0.dB+;6:.GfL
1aE(Te?PX6Z-JI+2BUGU&&L8:1YQ_cZZaeQLf-/4Jg@aV=WdA1&=U3CUQQAX6KR>
H;3H^.b8EQT5f9DN1K2YU9W/O,D=]N5>U0^/QAEfKNeg/2H-V@YTOG0bG6aQP>X<
]4L@<493QI+SG,J5):-ZU\R5e)d:L+&;LPE.b-6;7b,:-d\6aFfT3;.;EUQB+;#N
FCJTcOCH:A4T#^GBDJ>HXG?^T7X4NDE\AD+1:IW@K_JG6dBbdMG>F9;OEYGSEd94
:;9.Rab4ZXS#DO(:\?<497SEOTdOUa917T:=T-:dGgb9d^OJ5c=O@<MV5&YV5]EZ
(+_-_,Pd71Z)fU#QQ#\\3_QbHdN=Q-b9+caBP[7bQGEWI<.#/)fZ\?;9S-CK0[#0
#9Gd:dX6)+,B9FBCO:g>HfHe+XHP3;W=/OdLJ_./,&AaV_V#K0f=M,;?@ge[,M]8
D\V>a<OOENM^fK;5Z?W7F2R\,4GXRG(_?Me/:XH1KAKbf(XX4Z9&dI[8GdYK/S&R
R/PMQ<[7a7[;B[AKM4618gOKT4fEfAaG_=^d<0;6654X=4I(<)U,=/bZG#??/F^4
JE@[b<H1>UYW<P)9RdR@=MS-CEW^NG:(U23&_:0&B>LcX45UQB5[AQ2;66g&+.7W
TOH\]&a.M,391[VT-XC]S6P-9(VS3cVN(/P]).67[P6)\DQI-6PAN82<=\1MUbZg
9<TVd,WdI@\:FD9>#gc/-].<SU5KID_:IbNQTM,+(L(,A&]JP4)F5_I@<K_:,W5L
VXY5>LL5F5#T--ZLHgKg_;EgO\)\F?G7Jc)WQ>QJRZUAO:;ROU&XM,9?&a>/=BSP
/F8H8X:51dGQ8GNZ^;E[<&U9UY\@=f3^1gJNFP((b,-VX):@#7\g0ZF<6+#P^3WN
,9:2^VCfHZ4.NdUOfLDCZ>L<a^WIL7/0GR_T+dT]Q<.L42K<4/^M=WDK4_>FT.86
H(3e^BEDZCO[1&CI.BY.2.[6UC?IMOKU_RFc86BWZ^L<2VaXO5PO/O##W;Q?K6fS
LbU7866LWIXL36/.[@LQ<d])<BO^faRb57gOWY,-:QU_HbYLe?CYBfOR^L1I77Ja
=+JFX;d0HV6#(AK.4a\YZTC..H=(]JFL>IEPd<YY\#Q(H<BW(_3G\I0APK9)bMBR
=:KZ+3gS#4CRMB7@-3;GDTSU-51:S,.OJEd\J2AD836AagIY_2)H?RQEa_7NQ(gL
<TNaOWf7,VAHVIORNW^-]cT9?]QL&-)?38LSPL>Db27+SYG+TD2?&8^@FOGgPG[P
2]dNI2E-MH1P>#QTHV]A:F6PQ,=ffea>,V.;GBMASc7e#HY8=A74<,_BBFS83G47
BOC:P=1GP0?E\7N[)]#UG58d-;B&08Q0E[UV./^E@=-B]?1W]K26eMc+F(7RCOAG
QIF3A-<e0C;5@0X&fFS4@J(/T_Q^,_VDBOfV(5f:2KK34]A/EN+Kg641B;>SF,;<
CU-b\IX[)B9U[:SOI-fLP?H]35KKcef\,76ScHGT/B(X[I+?M8>Z:2PR;:Va?P3&
=@(>=;02XbE(BI/VVZ6Pe5>:gIK[/&]M&8H?E3KT&3SS3N.D9-&+WJZIfbAIIIF9
A,/S>49SX,A::d0Kfa_e:U4<:6(RBVTfg]BKIP2.6[XY0a\3Q&VV85_1/faRN5V>
]O;AH5F6B7/O?DGWD+]?Y7^Z@=NM_f7KcW\A]BL;Xf:FU4)8GdgcR\]0U3<RdCeY
b+0@3.ISJF>SB7?HSK8MUf7^81H:_Y[5\Y:5&OBJ5S[YO0N56U8L;NO9.H(X<)O:
@</8&O][5fV6EXH1XCdZGdK:M>V3DMaH^IW)X8(LRSW\S&(&8)Qc:99aQ\B<XQZ.
&2MPD@.P@1?>K^>edGZ-^CM>N0)S5\b\0C>fNW0WN4]>^UI-3T]]/@gE_SHRPFd#
Gd&a]8e8aM2>:EF5YQ(7Q>J^-=4AHDLTg=&HS0VNXfN1g6?-1O?;L-V51LLg^[D,
@_:<E-gZC0_^W0X+#6#KMb[W1L/CMa1[E(PdbS?R32A&P^V3H&YUV_#@Z]0E01OQ
cFV<A9bENPN+\?VB5@c65WOG@U^][+0P^S5>Dd&gDH:_KdU70ZGWR9aMJ(/b^)JC
AP9dA4X7=^HL58b=WWHWec2HLK\@be:)96XKT+.0-\E@#KKaA]fZ,dd0X,,Y>5Y]
R@I4R;SLT]B:@M+UO853YaEDbB)-_GA[T@5<Q]L3c_V9KS]2O\\6&MCAaT6L@T@L
JYVTDAbO6#e?#[Efb9,g39PJVX8&X,WB]F3NLPNAKMd_N47AFcZ5N4(ea]5Da/#@
?dW-APe[ge-L9(aRMIZ_WS1MCM^PZIc8H,MH8ZTceU9--C:Ec)ZS80(H&c9,H3F&
SD^?e<5D=?5>Q(-b;?R#30WHXRP^6\DCdAW/fT2aC5;C/.P,A-W9Y7Pb,<O0RI@W
?dIL(3:NJ(KVXD;QVUNb8CbXK&+6(--)HJ(4<:Q?7^05e]N]>RE0<[]YR;Q_T^3F
VO)F+S)FXY)ODLgL6J.KGYgP1ZY-BAR-,Zb;fJ1Y5QNTU(+M)S]ZHP<QC>H9VC_E
RF#A6.bc(1WbFWP_gaX.->Z3/3-]W^BBWJZX8Q@a-?(J3c4F;4WZf#9FM+/ecd\;
(,gfV;&b[1BKZI7Ma3GD^IG>Q(FaPeVEcQ\:40.Ygc56Y]K@4D2:M&).@\L&,A_M
H252Z_?7Kb5-HAR\#ISFS<H]VLb:MVW6)4M(?)3Z\+g62SW]1WER\W:fP(dg+J[b
9c/@H+&^Z[deQT+#WNZ[<4g+5Q1[[<@.8_/&G>H(De2C2H2;42:2>G,]?15??@2O
MHRC_W72eUQCTc-4H1H\HD.FSWSb)eSOH)IT[e:3de;I^gR(N6U9TECUGf6:;>^<
3ZbQ4(?c]8eaAA.7:3g(_H(DIQc_4B@+bOZgaJI^SNVMPZ_d_/gLTg#00DBPXDM^
<8=)\&?c[<:5IEgDEKNQ=XU2-ga48d<7WQ3NVW/IXQd8PJ<B?XUO@g:#J#df:5U@
T]Q\G:\5X;]bJ/-6>5I=7-VS4K=U]bD5Vd3Q?9WYCM?I#@#IYL&9c2K<^FCKH0_;
GI-4:(9_O/Y;Ya6feR3Aa2e=f#Eg89LXJ&5P\TZK:(Hb(JEc2<OaEbEUE127;(I8
_;OBZb,MUF+g<N]THS\3[9)Y:UU+GJ)4Y_8F]+g3UWb;WKP+8DGQGN#bO><<RG24
W?0L>F1/bVQC=U,Q&/>@cF1aEFYEIbQIZ3&PAU9_)K6dS3\?ME_3&KY:;egBCR0R
-IWb4B99=,P)ROXSL.d.83T&U_^ZL97:@,8:0@Af<AU4^cASPP4e,MX_c&B07GdJ
\Z+L4XNM)-+#eU1@2DB6Q;4aCBAf&=KB4[8+JGKGX)CA)K]a9^:B?/#F8e[6D9ON
9cE@F8;a_03F_0Kf+cSCYR,L5.Cd&::W;.U\gM\OT5\XUJ9C9G,;bWXX#b^1X&M_
\[II#Q]=ZC)gCOV+2CUeHY3L;KY(LVbQZPEg+.CH0#OFQNdU)J1OF#_;2)X2U?cX
J75a=/2_JH46]L[(#RVU=&),4;34Q/KIS2fN2W)6^?C:Y7NF^AVP);g2))gOSX&2
M8?<_e\CH3bX5g[2[HLBcVaW;e^fQRGV[U]4A1Zbf:@gYUgD<)]caA3@S9WXV_^R
S(6.=\WZAe,PMb,c;-O4_3,7gf6)b-J]J6I@QL>-#/<Y:,Bd@.Ra?L8\7=8U4=6P
VXcKMC&[S:RRL?30gHT)X?B#[FJTO^,V/Egf;BdI2YcLS31IO+d#70SK2&f+d^1K
cT4NJTFD9BBYVcT:<S?A3;1_HXOdO:K/K#DUL89:d,NdBE46K#H[&@D1g<LLK;3+
I#VbFbd9gVB4-a7@6F<f+A#R9[T=:c2MY^,NA_8L#NEeL,>\SVH<+.\7WZ1P/N(b
fMZ]9(;)5(-.P>E4YXQG<ML>aId4G5^X9RW;;J:AQJ([G[.T]7gSP;EV7]M3c1/(
D15NEY@N_QD3R1d6d-^91>.E;=V=U=(ea7\Ud=VVRO)E]1T1&4>D6\:&=HH-0ZB7
fVLQFT#0GH95=)_:e7D2I0e_.6BNM5^UV=cZ:dYC)QP2>RS;J3B;-FCW]GM_5\2e
8PWWSXSb[V1_^YH@1_#[e#4RW\Q1C[cKT^)Rb4^3([[]7;_cPQ&;GNcDMJVfB0Bd
OX=_)[FT4S(;KJB)f3KZ@C8Kg>K1c-#7>L1]@^W([,K/38^#cT=G2cH4SN/9E8de
aEQcc8JE,_84\<)@0HW8V:Q&gL<4AMI@@,Z?bD,0@G_Q(Rc2IUBdYbR?c^_T^:4A
I99_O+XN@IER5U^A21LY49R_9L71+eDOJ([\@=BNG)T.2d3WaYBPWPI?#\#Q:C7)
c>dH^@EDW(CUL+d:96VG<?7Y8Sa\6E.^9?,\0OcBV\5ET\J]K[MXfCHZ5=b(I]J(
fYXEfJ8HQ32GU,\Gfcd,9<P9O6AKP(:/\UB:/,94\a^G70/cP6SIc4T<^J6K2aM>
]Z1:LM#8=5@&1JK.J>N^V_L)KD.7ZYcSWUUX8J4b6U)N_)+3Z)6W)1^H6[OGfH.J
L]?QM3^fdNG2AYUg;O\_-S(8XN>:551[Tg&/d05T:e8VR@L<A:6+Y05#^Y\)[1gK
DC.)Hb0dS@3=<@F8:.#4eB]6Oe2MA\HH[F-/P-:ZWb)caF[3==cd1OE1:F/7Ed&?
g@)aO4W2X3&RQ.G4HYZ^eg]H^G:I?Z8Bb2^1\9\).Y@=E;V4.)4^/fCD^/+M-]XG
C(\G7SfN6d<OLW_O=Q.bG\Z2e@PIP-201D@#6K&><^DI[._:+(WE1529.cRK.<>C
>[OIY7.a]F<44;fO_EH7;e(<+M12P8O+L9a/TWEVV>\G:+9W6)G^5(FCCF.f&N)g
MaZ^/UVF6^@0@)J=5X3J0E4N,Zd(fea]-_@?13ccIFBTf4-b;;J.61Z9=>eAag>5
;,Z_M/8+YUb,I1@#B;=E8aYI<Y._(\^.H[Ua<6&SfQ+_f#]<4cN_2P4X8FRG&XQ)
YIbBM(OFU-A.6U;Q.U<?TNI==gV47b:c8.[bB[A^;@?D(aC6G>TCZD@OQ&ZYHcZ,
[PG>EH\;4\LaX8-AdWH=Y]&UE+R:MTMXce<7F@<9aF>fUKf/;OJQ4#M=;A6d2A>1
8Z1&SL]M\a>eZS2e-a::LSe.eM24JeB\>2O?H2,6\d-RY[c#=5eSHIPeZ>IVDaP:
8,EZBeKd,Y4C\(AHagN6/9Ve];O3RVJKKI9F5GI-)_JaLA[1bZVDSTQWZ?OR^SW]
d=1V^e>(HeL=aL\6]I#/1)a9I3R1f2--\R#f2E9/QM6(\][::JgE;/NQ4L/G9PPO
XaW\,64Ld3fK-2EFDG@4<IMM#2W_18JLcJ^[MLH1bKa&I-Q+^RHB@&[L@gc,<[NU
B=R=XEAY>8+M(T+O-RJ(fM;;Z0Tg[E\=cEZ<C_g]JH\Q8N-BL7Vb-]4?:^>0<Z/;
@LCY(+/PdY/#H2a9<eL[KYLNJgOS<fN03R5_2:\#2CFb&OdQ=P0b[BQ:PgM4&3DL
,@/1S#]+3cA,ga9BcV\c_fad=P3>:]B#a<cS<:T(Z-ON6XbGfD2,EfE(F40Tfacc
&(+NFLDg_I4#F[\/<;:QO50V#f=VJ-9+),6_0.VWS7J[W5_3a(-&_B4>3IB)5O[J
8+R:56DY)aTL+.?QZ9#93+RNEDD/eS_Jd/fG7>8^5GR9M?I#<M7S_]M+=XYeN:c2
ALbSZ]N5X<OP^_HI<1d,AGdF[0A[5QH#;Zd\B<-HW#//I131VRI;9-egC;7WGBfc
e.1J2?9BBdW>5YBLP)U32bZBgSc0OG5GP6J+CWH-[aeJ-Z&cd^Hc02RBNIg,X=BF
K@6@?SWd]28-[A3f&X/0B-4T.:E&0==>dA#7600Of[:S(S^+FeP1>_,fF?_2N7>)
?Wc9N:/>,XA[7U8-5=N.:#/C#^C89=#;S<gX5Va6T#U65?71<7g.>ZZSO0#_S=I+
-S.c_gNd/NG..;P^88Z1][9W_O?(_cRE8:Q=WR/&.A6[K,R.+0(8O-Y:[EMY]dcF
;A&a2P3<.d,QQL30F,;3A&8.Fb_:GeIN.J+YS/CVeL&@Q+U.&\44FR@Sb]2[O<@_
@YY+/4B58LBTM.Y/BJH4L@P1V\40C@O[VX[2:H.0<<:+Q?)0Y?KC<GX;V>-0E#]>
U)9^QHV98ZVaWJEX:3bFF>#fVDVWW#R7KO>:O7VYR(^64agY=aWUVD,YGVD#]b\P
[J[<M#@MHbH0V8@7Z\1J-;ZQF]<[:2EaPG6DS@bRP9687NcXEV+R6=V5?eOX8g)6
FFMYK&]e??WIN/KMTbI_Md9d7eWNeFI22<,XKP\CEZf1H^cLULIL.aScSEb<(@UJ
7O?78+?fMEgD<Lb]QJ?_C\[I3870L\M0+M.R/LVcY]_cF,aAP/8ZcA7OGT[1.^Y.
f_YXZ40P,/R?dX,eZ=U?B&\Q<f4Z+4C79966\6g@Ba1QWIdb@Y97g?YJ(<dWF.S4
&cX5^gdQ&e25JPW&KKTa+QD,?g>J5F^/Jc(=@8e@0=D+G6\TdHU:a4(MT0L;I6TL
0=E#GQY,[C?K;Z-cI.,5OfK.<<WV/>93;]@[]HU[E4K<?ML#fPMJ.c/,YBfVC@:_
aUL?TggW[)N4)a-4Qf^EX=)[./C[R>W2N_I^MeG?.KXNdaO(+.Y.Me:9\(3OJ[fO
C..8^R5dCfXFdH02C>ZdT,F_>X8B419+OJa3^ACd7O:S.K2D8b;AUXT#[a:U[eW-
8]/]/MDH\b>b4Ke7:FB6.\7Y^D0-&+02Y77B]T]K,YZ+ZMOBF_4C/6Af9@=2&dS1
T9=0X7F9=Y7\4&N3g;B+P\_fQ0COOJ#/R2fZf:E210CKRQUbcQ+D/R,W@FA(K2?a
\@^Jc-(76M>;b:P>(aM?Q5YAT^<2gFR\a\>c&O3^eBY7C+YLK4S<G<Jff2N/Z&K\
/LL^5bDNBX9)TTFf5K.+J9J3RbGcM.97:++K_2Z8>e&M>&+?=dAUKa<I,,T?CE4)
)JRbCE;^5a<^;C=DZSU0>\^U?R@L[B&T:GX#[IZ7J2S>+J0-(ea<MG](D57_;A7W
>BI?<SV^1aDg]AY5#T)Z\Ud\6b/bf;/1IFURdJcNFT0.N\WZ.@?U6.KX3g,YR-&H
SLF465KJQ0_.(2/?H_.8ZE)dBS3QAN=H9d-2TJ-3>&f@Wc[-(#a^\/:.A-J[<I?e
0VA;#dHeBAGf#6/.9PLS1+?(7YX7dX&LRM&e1JK)D5GIXO17;^T3bZ;;F#\H<:XE
94BI8C41BgIP^,:D;-UHgD,#F;/O;ad4W4cf4b^d?QW:bQ2b[#7bAe];KC##fL,#
JP3?DLT/UKIS3NWc^J_,Cf#4)^;J]-CXe&((T5QP9ZLdKGebEE>AJ:g/JZH?WV+O
P\GVLB#D]e0?b=VYYKWB(:YVgXR]DgH<B&];I>I5C\gPOUEa[@CQe+VXFM=Kf9\\
>Uc[^=VAD[.aA<8,bQ;)..+aBZF@eZFZE1_K9Q+3<e0/&.7;T8P56MTLWg#PD>=@
IgF.-.F+dO\IaY7&GJ=ZN0La=0a^+Q05_EO7a;:9[W1d\AYI9(RI:B8-4AB6YcJ)
_R35L>Db73Q7U,09D8ULTCU;PB_R-KO.P&,?0R3N8OM9GfP=&N:<E2_?(e_V0MDM
d09]+<#[(^_+DD@>?LGI><eXMP.7[L#c@?(/^KQ/=U]F_G=,;R)H\+>=?MMCS[:N
[2DPN(bO8fP\fPMSG1Z@8+d=M?[Z47.B0eJQ7D]@:8)IV[LCK.4)JfB>a4#-dA#7
1],T9JTN:Rd(;EMA+A,G,&T?H@b7@8BXNWZQg&&6cVR3H(cPa4AH\^BVgPS7I4;O
PKQYLa+_G6e3LC5_S?BMaLM</UHOG6;S0Ud(fL4HC2Yg^Q#/#+>SYZ=G/;T.Ge(2
dZ,YeAcZ8=aASZ5PYgPLMO&<7YBLecYXZGN4]I2(\V]2=9@\aaO+>(4X&.YbcGWM
WQ]b\G^7YDHRa2R=/FY]EVPIN(,<Y<I^89>b#.d1EHa:+5TO2ScXd)9aM)f]YN7/
:Z]8cTgbSdA9)3E<VE/@/C_Cf)GXLg:R@RX0,:S<[CKdDbHZ4LP,;9bc<+I?6J7S
<d9:4&)bR#2.SVN)&g(Fc[Q&IC7@;89AR:ISIB],+Ne7SN_U6YLcgcE#B#;;5K>0
N2A&KIDWf.V,N:T>V,\ZP0R@BD(Fa(>^d6]N<[#S+Y&c#V+):)N7#81ddcK)Ac^H
\H+gIe]X.H#7\M:J,?G@FS2,NFW_,J;X\ffZDZ,AZNU(dUX2dJ-EIG\(GX?-Q6I+
c,BZ,<RX<BaQ2fe\YWX+)X9P56.ZD]0QUM)<]V)-3f&d+:41(PIZ5#G969[aVFdK
Ua[fZ)>@SN1OY:.+PbVT52McUUg@GRAKF<CP)A(Q6V8gUAX#;[c@+b4Ce=D5XP?<
?IZ1@(O7+4-MNH(PDb\RId^dI[WSS+O.NC^I[b;dWb5dO^6P51)06BV,^#>\512S
NM#ZL0;[(-XU#fI2GdWOa)A=^;[/5#E,@7=,,4T3S/IMY0_Q7dcHU13WKKe01>J0
(Vf3^>->G=:)9C?1QdbQc\#\fGKgEU\^YG1S(dEV\^CQT12J7,^1<U67]HUQ9+V9
f0.5a4dR^(/9SOI1\aeHG;SMa_:SLg]Y<N\A\F9TAg\5GfJ&,\W6O]/g6KP>\/\3
V/cfU#2NDe?5f<]+/DAWY<;,A,GA+KJ.TRZ0_IHA3ef?,[G-Z&-->6DB(,RHTUgd
6?V#MH;DAHH&8HLY>SDTg&<U<EO\5FJ<UA4)5U68MJ:(7E50LBBbCYW=PL<+X?9e
:0OYGRV.EX8K(ES[=N:^34>M+\RB2.;K4S4A^CG_G[9N2G(<^]ReBf#/#\S4HfZO
@N.PX:/H?N1KUGe)-3/c>9eD4gf]defJc;RERO1+]C6OVLHQY:7=MLX+D90PUV]G
@QQZ;)bW<7<DP8^-]5MZ=?B6e[6-SYWM8M()?D@^D2]3Z:>2]1Ne,M<<(.3aM4+?
.<4e^:)]a&@A-IY8MEaDY_(TGAQb>b=#]T.K-RMHb0ITPB=68;H;K>:BKST#^WaO
YM/fBW=4N)VaI:C&g,(:9[6AQ7-gM+3GU^M_]QF-V^NOUZU&?7P+OM?TNE3-/@\H
IeFb8HBEb=)62/6[B>[Ee#REfGI&E6\J-e&N(:^a4PTBG?>B@S>=W2#?9X:16J6P
<7efYW01D22TQQ#<<Ve+R]5&8KO<dW?)#?)50&K/87cY886L7^BYJ5FW39-4Rf9W
.?f^#)@VML3Fd^=-SX=d^@YQ?[;;\_4E2FO_g=V+2cL_ae[d6PK.dfU8QA<@cA(8
>,FB?TU.E?S;Q^9JO)NW4/PBf8Z(?T0M(=&BB63KfV9LE8LS3_ZMd_[Bc)Z?_2A&
[QQ+;+&;#aK#(WLDV0.X=9RK>59\^J:,E\X(E@K4N;\1S+M;2Q_Q3YPW:]4C3/2e
?c26Z]O(2Vde5<5<K]+U.\S96<7WYJ3H3O=X4RLCI8=PWW8P;EXeN-/AT8&VQ,g.
aeP?fd>Wb?LT;RU_SBG]EXJ\)\PLJ-E1^fa2V,+&+aDEc1-:(@MRcH1+Ca4PL1DM
?f3&aZ:[:BUbBVBTOY.&g_0+_BIcYNXQfOHZ-45#+=>AYHD2IcY,RQ3/BgFA>\?W
-5U>]eC^fYPFP0TJWW.0X2Ca[5ZK]Z&2W:]VbI=GR+RO,P1JOX&gJB)-A-0^)4B)
9ELIe3.8acC\^d;[b\/fW0>B.f,NS?eH@Qb#ECJC9QEgO\E&(XWBBD)>0/I9f#0#
f?(?b;-&NUW)(4<d8QB<bBKc03DE,PC8X=-J]65[fZ25;2FRZP4Va@D4HW3[M^b<
H#Pe^[\58g3d;S_Z-U9d12cE.Y?a2MRK/?Ob:(>A6SHSQc.PH\D8Y-#&A:=NKZ73
AZ8eH1(7/W4BbAB)2L,?IE<<#.-g\f9?Fg,C-bP-76AF_CS9BV+e:GJZC@?,aPB=
+LOfJATS.L]UQ)Z1A[\D7eI\K,W@BKBY?a-XI\I;1B.F=fB[F,1LWD6.BaD3G4CE
XgOU90UM=I(9.+D)S[]K6E.dK36bc&fYXV.#;/2McLHbUYf&W\K.Q1GNC=A_/f)f
g3N:LcX>bC/&fZ@d5L_?PTSLYY0WEU]PI73[1];]74Z\SG,Hdf>M1A>B?T#XX3<N
W,>B))R18f)0)#8a]EA-GMO8E5;URe1K<=3J&Q9ID5Z.##:>D8ga?NKB-R:P[_I8
LP):;]G:c,/Cfb\G6@2P]IUe3fN]0e/J0WW8f:SQbTSXGU1;9TLTeS<4H@/#J1D=
IAYRQ-[KNQV)4M^W9bdK>dc]cP,Xd-]TFgC\DHN,:J,)MJ4WIfD2FEVXRg<^R3cW
[MQ085(WQ=Q=+L@U;QAQVKYH84LIZfR4[V+ZR1CJ7K]ZZDJ:_2HDA+P=-2;#dC.Y
V>A7^E0(#3Z;N&74E4&,T@J,?aO\U&ObR)&<J0/6/DE7E1[(J;LQc3,H?5LD334W
ZX+4;#.3?a_8AK<)R/+gKZL[D6P1V8//gJ?ECg[EbM3Af;3BC3cDab<]UgUOC[,]
_ILP7ADWUBNF<:-]b7J#A3];LIBU8F7+=\:3SDVZ.<B6CY>;M4OU04.)Wb7UNIBL
=dYc<a.P7,cLR2WOQRYK+b?;TS/4HT1gK7--;(L?7UPO1SRYc5\BAL5U?[bZ<_.F
;dFNOf.HeK5.bJb8:eX]AZREGQ;>e&I-15&6:M,P:NYD8&[)<d4.DB1@Q9d2I=JR
<Z@3H#/4g.^K)O;fMBX[1eF>[Cc<>D1\N6=-&H[R-8^=_C/W\K_BRaL&9S<F<7Q=
-G<<<C8_.WZgXQ[-=N]WM.F2XOe84:=cg#2NDYf-K5,)_BGQJNF0#ZV3W-5CD\XM
=VU3I3,8\VIT3F3d9eJb==)-C,_EeF@QN>Rde4M,f@f/R-X^=S3Hc7cfW_LG-IH7
_B6G=F9dH-Y6Qc&Q<-\FP3QI@YQ5B:5HWEB\d]?H.OZRQbbCDQD9Zg_OP)d<BG#F
Nd7)gMCJ:V][4&]D.H]4?c:.HA16FVCBEXCDKS]+fZa?:fOda#+c_7S8B:X7Z;9.
5.;8^Hdbb-P&+8ORU#c/GPZ(3GUZJ@U5::8<a:,aa@/YDQfMbe7?9[84Te:LZce@
M5,VbF#10Z:;9?gAc7\?A^\2M&/LR\D8.f/9;UX^0_f:AS@9@.7B#C9EM:]F;eG1
CYFH[;@TCBK#Q>bRQ12:)G00I4d^BHC@7e+XMTE.I(5ZUP:4172Y,M32AM,dFF)(
>SFVLfO1)Vc<7G^.b6c9Y=_0[Xf,/-EF[@f3_9?XW-JHA]>c&IcPfd,]6[.fWbe:
HfHUV/9Q@MgW;Be.g.f3\N9#P236#J6:VS/g9?_T9W>#TH1ATF0M(\JQ7BT21=O.
#O@0I\\.4KRaIMCH1I8VEE9P@EdSKYg1,&0d5a1&;7LIb]6.Z7daHDeK;PICGYY9
GUa7@U^#PLN+FGU\GUZ(.,ZG##fL-JL90b=NZQ@IUa#LNI,J=ZNG_@+,X<g^-6).
[,>#:QTIGKF@1YOS#+@0c&.OHMW@7bTA3=B\D]7d&I&ACQY_C-Rb]O(gW>7,RE^V
Lf^L:>XSOXJVXLRb[=V;RbN[CfC/7Qc5DV#3C-e>HD6W<Q@>/]N)_3a]^Cd[;[&.
Pa#1M+75/5/N;&c?e(YU6Q;5g:/#^]WWBF&G\3DaL7fg0RCS7_,K:SeZWWA\0G<;
=UE#5O<_B>ba:02PMHK3b;R/5YGMT1SNNY)9=.Q9O/Q;8>Y4O[OOV&)^+8HK]Y2^
bZ;Me^,P5K_E^,RK3c2@LBX2;PV9J47N<6e0;]NUaBOXL#NZ9[4C[VTI,37VWfUB
\G@cg\a._M3eUX-:SC-VJ/abE,)QSO/9>b&&Y(MB(,/dc6gSA7+UKa>TFfG)E6I[
0Gb.51INaQWFAZGY7<2II),UI+,N=HHcDT+A?;:,883GOENM^.W(LVC_.RLH;-MM
VFB[UT4]OXg]C\3VC+#>B)5(J^H<8]1BC5Y5#9B(&=,;c^.-AQTMDcSdf/DYgC#c
5124a\MX:JJJ[Y#V,M2?Z&^=LZ]XMU.Y+4S_G08+g5W):@/)H/(D5@8eg/]A5P#B
I)&L0@bc?XaR4HPdE5-c_Q_VXI^HQW5fbZ+&:>(c>L3V_GGN3U-/O>ba1<1R,W-#
9XKS+[^GJcN@5eNS519MTKZUd[L+_EDXI-R#2&GSAAFXL.c(b=\U115AY5)=+(;\
;-Y5H)/]B(8GVO(D--edC6\/CHb)1&@RAJScP-NS__;[LG--7MUE2:9@3>c-e]fK
DB>S-JLY]/Dd&AKW_B\PHV&PO5&IM4]\)WF7&0#9<b1O:8EQ<=#:a_Ggb-:?+Ba#
^SCW^>RHe>EQHT/U:VTBK3@Y4e@/;NF\.K,,F6c31\d0VDB7/F>bD2@]eebb<.9;
BJ.H35=0Z[]:#8TUWddfYPUc]?W&CC1IY;39LUI,#A3e0)EY&S1>7;TX8,VB:(,]
deQ+VV2\[GC5(-WA@=:5NR6?e)FU04>;1Ab3f;f/FR^-OZ9cEDW]:da4E,X;)_[a
d_S^R)+KE7_&3-_@f@d]d;5)JN7J_M;/0]0a,XXg-2/e@R8TX,A\7?+(TFI>NMS/
<HLf>)R0=#7;PG?UFD>-]O3fR2AH0gN1+35Q]3NVK9H+[Q[?^?L]aI.>GT=\XH)R
[Da_(BZY\<d5BV[d<:J_,X_WL4G0((XP.PfG,7=D]O;08?67L2(G2BaU?)6SKHcX
?e8(:#7RdS5LG9[JU5;6,3?3[Yc40Y24D)(FR3OV>2\cc_@;[D20Jf=Q(QU[FS8:
#BC;RSW7SP:R&UA=/AQC=@3/V9[H]ZZBCf\RC7/T<U(b&3NASG7]_VU15Gea>:#6
CHE6ga]LDF^VC,?fYM/eF?WZMWZZF25-DU/c5/Xc4+LRd;W^7e^-V2AF&N=cU7Yb
8]]AR_>W?1PC^V0_^UOG<DZGOBgefXMD2V@+1FTPg.:YZL6?3)H#012W:GgaI^SU
cINc^1X]2F6X/B#BH51)#:<(7-:FYfYE[BA28e#GVDSXZ]AR(KP1PAYA<Y#>FK3g
;Xc_3a&(@+MB@e/6R[S6TD-Gb]W;=OHUb2.XO<SA5d#9DW<-3G&B8WD(2ZAG^aV0
g^9A9(WaY@)Ad\K<E(#e:&@LC>M51JS2a@)FASWS0&.P^P;SZO?@I=g3<)S&WQ9@
bQd80V)<IIEH=&X=0&(dQ^JX@PC#\A5?85@b:E]W8a1DV^aPe1dMd,=CC48Ed2<:
T9)9HVW5K/,K,,/HKJBU4<0V3\E/f[AF:_66UXSbQV+>Z6YPV[]WZ3QX-ZNN=.F2
2,UQPW0b54\SO+;@MN0./DJL,Ua=L2#&^Pf.P271^F[7bg2UGB5DA>]KfDZTE@H3
OWCL0_<fcWDV]&UMUQ&^cOeV65D/[5ZLb2Y<N5^<0>Q7_gS<NVbd<g,@=.-7Z?bA
@eG9M;#EBBTSI[c:^MICd](YJ#^^+_a1+/GLJd?2)C0JUEAC10SFI_fB,7)?C\K]
cA65T3^FfO-PfWU9(L=LeM/V:eW4HH+VNASbQ@X>4<[9K4@0.dg-cFLS.NEOYe2R
<BgD0@>)c/6^:#TF&T8IP<E;Z1>Pa@>#9-=A_1;dVcXLSQAZ\V(4cBA_Y^@/)VIH
Me=5N421=;HRfL@_eI3=C?@I-#16@I<D_NAKgg18;:P4)7W<AI(\H3.(2QS+PD^@
Hc/\LEX6H3<IQK?\0(=@E>S_X=6]SGQY8@H:g1?/B0O\a#c.M/:bVMR47e^E)IOE
K6Q)>D/Ag;EGL.?<40d\SN=E[XH:/]6eG+SKELK.AFLe.b8)BE)Ib?+?LXb5K;W=
.>HT35B[^X]+E:4=ZU9MGe53Z]2cM>4gQCL6A7;60Q+I3J_;&N.J-HT[.(3DQFc(
HBO4FKXJ#)?VC&;/E:EV3O#U5>.8:XIGM/Y]=FB=2Q7E[?X7MMce=V[@9XU3F4N#
;/OT4UR5:0K3==484;J+)PYZ(Q.ca1@->dH,ZQaG:VI5](Pf,9>K79HfU@J3+((<
H+#cH4:bg^@T]4e-QBOGIaaY.S/4E>VfX,&=U6\<JL@>2/bfTJ<BYI+91E.B^F]d
&]>=-TP#,E;SV\dMHM<A?J?)@RJM-2+L.a/P<S[5Pc7FY4_BSKF;NM0-LPH]ZJ@]
3,eNJeG/^fPNO;II]>90a7QW5^+_G1bX[U4^1F^\N&aX6[)LEg,D;0J0),(OC@BJ
::=WGUSf=-FW]0a7a.OX34H-2E9K>R7SMSaBgYBULg1V>\8F&W3D6I,DFZZ<<Y5J
:9D+8?JBg?M=1eIcU4a8RW]>NBf)#a2&BM<K#U.F:b/&8cff,e4J5,_Y^e)\?(8E
3L.gOcMF7^g?+#</^2bTeH8&YSL_8\0EFU[(7OYZ]MN#1@.eNADPWGCRL7S.FIIM
.4f=3#J0/\DM81DL=B[SUJ6a7OIYNePGC/g;6UT)=VUHQ1,dS(O-IM25&AK0@a7E
dX6#D-_cEec?Aa>3.+@.HL4@&BeZ61#NF[4aa+MF<R=<NOC+.f/L]8K)0AMe<+f@
M@Y@5I5XAWLE#+HIKWWVaa[^R;]E(SBfcgC#\0;cd4\NQ1D97EcN:DZA88O.5K;6
9c)#^;S@&5MP7VA-MIKA1bU-4__d<Pd#P@1E0I>bG;BLOF3LXZ+OP\DWQR2@I^+C
d/@O[T0VaLN)@BD5B54_V\]GKB[+KQWePK1GI=KMH0g,b,C,MYUC7&P?S.VFK9PK
K=&]DE?#ZaS-0&R#L,UN>2NRXCEO@3LZT/QN)Ce^R)fMcgA\>b4cOOUY#J6J)KJ#
MNCRQdNVF.JSU@7@&(]7.#_#eX0@W[PcVN&c7F5:f7-\FJ=3L)SE#,ZOXLDAF2GG
g)\#2/<T>O1bQ5VB0H[8)]KI&L-e_E-@0c<9]BGE.MI:b<NLbVc>&&Pg(N5=IdRT
W((BeC8-_;#;H<[b8O\6:@=LM_.)E[I@KM,g9cQVZJB^Se7@3fS3/>ZSFD]0g@UQ
O1J2c>[HX8?P&c(J>?JWUE\MRBDK]JT&=F13=N9,+>YDJB9c1dRHg_]S[2UTMO35
?_M-OU7Q9_8ROF1b_.c@.T]JSe.)WF5.7<)gF3IcRfLKa3&R=(J5(LHMS)9&4Ve-
#c(e5JY6Ld5^T\Kb8D2B3@L/6I_RLA5#5La_5RMb>#2<JT(W#1\bEI1bbEFSX#M\
gC4]S@#EMGP=@T?_KW,cfFN;Hb&V4VRBdc0DA4^?3[<:Q]aLW<ZLF6Y1ce>8,dK_
^LDEP_AM8<#eXd[_a.P61QH-W9[NY_X1)II&0_8#->.&OLf]<+C-D?Z4Z]dTeC_L
(X8M.B=AU>OK&11fJ-NG_KH\R#UIR^D4(VbT2/V5e:&aV_OC9X)0Y+;aZ<>/b,/8
\AHN.H8NeVbfC/&_C&GU4f.g(a#OV?[5=[@#&25115C\L=@O\1-QVFP=\?H,bD:#
^[K^f;VK>;FG)CTU=SPY;L?0Kfg[4Y\R,SQ::aY/GgG:I,3P?L(RXXaKK^cO[KYX
[Xe35+Gc9>bU_a-3<[)g8gJ;,X1]V&aL9&<(Y<>C.,KGc3TIfO^/_gEMKZ3N0;3[
?51+K-DaO0M[2U2_\[X+&ZY734-63SDJ?Z,@>M>A7.fK<ETVQHbJ+ENT]KW2c&OQ
Sa1K_@L8?T]6J:@LV@=]fQ(>Z.QC6MF74(3M-4IA9F;QL;^_=CfTA2KWV<_]e5@I
\MFb,TT>0EEB)S5@G_Y+a@-cXBGY+:DI.>8M3FF&H[cDH_<IZ?Qe7NK#FG0ScbGC
e9:eT[3VX>-]8JRgN<0RN[#-K>LY<=P,dTHCZM9ZQNX^P?&VMI.WBAC:cP12KG,O
]5DC(JY0OUa)MFWZCE9:&;_RH_+240BST+T_SK>I48cc@>IW7_?W,-6C);>:@?4)
BJe<3aaH\M>G>#JO0>HXI>]H<EdUE#^4F5_Q/-Td3OE(WWTA+b21P^JXZ;D7Q^3R
[-),Ge+Y[DX,MKfbKMI,Q)R6]RfF:\97_2_2cBB&\[>I+Mc8/2P3700TEYS(NRY2
;S._G,SE3L?\R(gYBT2g:IY+EV;@/J3;ebUSP2+JRM&7.1,=4e,0-(#_F6H,MFYc
SN#U/f\G_0EEG&[REW27#N;03335@bK722M5bHEbc<&DCE>H9:G2C=#RY6RBDXAf
5Z:eDBc0_-=/_M.>M[:Yb595,GNZ0dAW@>6<N@UQV#c@@NL.76dR17=3IOUNVA93
N\+?W;;Y(_1KV9aG7DT9Fg\JBI.^.gHVIfE3<H:J37a:8L.1)ZJ3H.:PQ6+cg)W0
JgQ=XV]E[Cd8;@X0F(BBge97.^;/c9XWL00c9d.MLE1603P(J[b\3S@U=<gf4TJ_
P:2.BU+PL;02e<1<I5=L8a/bD(TWT\G)aGOZgbELQF?A\9T;/ZG?S)[>Z>V6[QC^
^aH2P9\QQF#8g253<_T.Y(2SS<6V:A)dfIHZU2W-,3-:+:Cg7M?O=__0VI@:[M0/
^VL>e@^gH7fI4aYJEKMI/baP<<U(c_ObA1aGL>.+5WL/^d<(9HUR9]2_+e?-cH&-
<P\I.MHZN9a1U3FEDNL8.T]?+[FT:g\H-MBMMQ&J0aMVEPS+TEC/(>gM9UMe^?&/
/8f]FH,8+E4LH38@(S-<?+@gNMJ.OC<65@M5)@]-RK;HBJ]WWW9CfP[/5bUe>b9e
^)VGJS_082F,bDJ]O:MgKc,5I5\F>I>c-?V5B\+JbeW:P]86QH3PU6Jg1IQ[^5X)
eJ[N9=0>[Pb&dNC9<@#C)N_AA.3E56#[\9_A9NW1^5SMMNCE#U=\.Q.Bd1bC_7&R
TZXIEfb51TcOc;a0^C5)S+BU14gT(,X7f@W?NBYL&1R0Wfd&V:NbJ;[<<Va@+#fI
3VL8/P1WA9[a@ac:D5bAfSH?UH9GQT.VHS=:4V]FIRcgPTdC-&9Ld+/Z?:RQ1G@E
eT:P/0FU_\;),=D:e/,\Q(PM^6Nd,JIA)DL\BZP-@V-H^SPG3gGdYbT1NBZc=0J.
J5A;>?f-;>7050-8YG22ZXEE<-[Q><C3]dGS1^<U1Vc<&AJPC>0C/E+-<G^?1ER0
T:dK=O-]=_VMHT)C6#gO2QH]f2=YP#;Kg-HSHb=YGSFSGPRV/^))DF)aPS9a^?/N
87#YdI7g0X[6=H.[3b+HC.9_#OQe3)O&e3^#e2?LBb)EBGR@VTJN9SICU386.#dT
P>S4bfTC6ODIaaKH+,(VOe_O^JdR1.;5c3aB\-8]A,916?/C_EYYS[?]/FaK&^)<
^CI=\-a:=0==]dRJKM=ZR>8aVbdG+cHV&L/2BU3/MGM/72S[gC^CHRN0(dIBa/54
4ED;7f8@&_-H;Z15WG3+<Kf#8CLL.5b^ZCBH\7AIG8fg_Qb?aJ?GK[GR]UNM+=YV
>8V^a4T-WM>_U<AW]Cg-#>/^5M+_(/)\?Y+U;caY7bP,2.Vg[fD-VN_3_a[DT&#)
]4YI..KC>2)\fY3V1DS3O[ML3>BbN/gTCfA/g0?=H;]CW9(\2\ggULgSJ&#^b.?a
I>9-OI@R\C_2Z81#gbJaZK>6S;X(7FIYDPd79.7NY&K\Ma4^&@0+.M.)O\1455O,
&d&cM@Ua?\#@1@<RCK[)[2dID@e^FY6RY=@MZ->d5d>3ORO-\;1G0S[6M),TA[;d
dQ/GAR<d2bF>b<2^e+R59@gH>a8Xd>@R^bgEAc.C).OIYN]UZPE#VQDg-FLOg1G3
>7?SH-_]>EGE72K3)Og@^Sd41IgY/R5EAbZ@c+N;@g8-TAS-;Z4&WW+0_=XV_Eaf
6S=dYN.#a/)45_L&bPF@#6&P3P.E,&1.V3F<,e.XI\SCE6]4fHGS#fPgd\:4c;XZ
ZV\d]d;+:?(D@H4E=0e@6QY<;\T+.Sb/>1#L<[Yd[Fd(_dEQC/_8.+1MPP/6)-JN
5DTbMf,HL>RL&.e)JT=2W/dc>XZ?@Q9@=&)CBDU#26U=a6>_dYF6fK&.R?SNMN=Z
a&_U6T(&Yc]dUf@cf1O?VcUJ.J5@NH7GaI^]\O+)d\Z<SHFN([(,_JQEO>+WaJZW
WMQ1g+B9;W22R<MCa7^=LH-ebL/HCRM-NYBWRa&+DO_2UMMZ]aEf></^cB8D[YPG
dBgP.4HHYgU2U]NPd3=(de&I-bb/CXNPR[CE<>GS#U5)9K33KQaW=V@63@TF>]MB
4JK>5HX+YWRacJJTg+7EdW:O_[N?]8AA4.X@cK2/I;2Mbg-A,:9Be=N@ZHJ8G\Gf
B,c2I^:C5L/S-1\80/G[P2VD1:;:48FXbf3:>DT-/JS)YI<ZYfK;490A3@S\C[:@
N1JTN&;)X.b;.9GLE+?fHGaaeKF7a;)C-Bag]E^9U(9&[(=bLG_?5FA=4TT+fYWI
dbMQb5.N:9R\ZNLM?1H#+BR=RJ(&2&EHbF/)7,YJf07:eJWZX4NH_O.6Ggg:-@-F
eVZ16:Q9D6G+C5#f>TA4[Bb-+Id8R@Cb2MJ8B-5fW9gH)3,;7Re//K]]V&.-(V[B
N7P]<gIO(6A@]9=)<[QSUY5>,PgF<D&V\>O#?4?04>S5d:]2IJ\@<P/#/8>:Y&6F
:RcCb[U?G)02eVL<&,ab(.=3<9Sa(\QPB3W,0e&W(<R;91Ad)5=Y0c+bP2LK.HTL
_gaEE[FOeOPgLVQMRdP&1D.-Z5b(4c3IV.?a\c4_\<&TJedI>S?7-K<I1@FR78O9
V7@L\E:Ta1YW(eL63Nb(4C]O0K[.AA0S>J]/B#M&Jcd[1MBegeIcc+XY,f?0W^4;
R/VX([1-E8KZM:7QF/\_#(2&cEUCG^,(AT,\e,]&+,P1+4-G]_,>UYcI+W@2LZaR
P,WM2W=0=S<KfP0f9UC(aQ9<6O4LfK4KU0IFMUCggMF5SNf6]5Y;?Mf-.2\4@>1Z
bZc@K8Y[TEd7&@17LR-SbQ<H0]AKJ_VgD3285(d7#9;H7-[O=[(5=&@F4/0UF^_J
gB@,QJe#_E);+f.?/5WPG\S&3AL^0Mga[HgG8B<;JIg:]W8bBD+[/f?S-)]W+>?=
H^7P#Y&d4\6G2\;aR.;3f,L;,FgcGWcO6]K[G.FfOSQ/#U[c<;J>E+;T6F_7H75I
OYC65@4gG3IK@@J\D8-KJ>aIV6HAPbGf<8J;,:c<beCT:aXOIeYIS<\=J3[c=cU:
cIL[a0S8@\H(H8+G)2@(Wdg0G=CF\1G4.(2#][T#6PEG&E\49@EC3#HWQ3E:J0=c
B+NP>Ge<&6T)N6^E:[<?QScTaP7;aYVDd9P+Q^>GJ>L5HP\656R3HH9DMYF?dD+X
^(02HC-^>&WNUP-#fb3E\Yd3@+bEQJ&:[#&R:(:Z_dS^OJgD>&ff3?dI]B5eAZ9I
Z2O.Y6=2++,V..Q8\E:/39[b@7Af[bKF=aZA4+2&^H<aK?^VCfX<X/Gb3>/If1Ba
9:_B204SCbF0dK&,PC1\Pd^E:H=dWA9Kc8F,]6Tg?I=ED6D#eM4[dX0[_\;,>M5M
aX-::Q<I9K(f/:g0Q_5Q>96TYO2>)40g@O=SbP]c9SPW+;_4g@g)c=WK/Gf9G:,1
F.H0<;HZ<ERc:1gOZ5M:a,d,?>M=BB&[LMR8O>QVbe<82)?f>P&Y+]85Q2YYa@:A
K0g40R.aNg]J&&:]/<Q<SS5_K3\JO/KXR6DcW=++(L(B#+L4f,4:?Kdf1:-Hcd]>
6L0cN2)F/ggV^5LT#:RQ&^J[TM1S5a,C^EG5HB-:HT)U[\&_G&KIB3U.>HX-QYY9
=S?9dgD1#4<\/.C3W>CdUafdGBUVV&V#)9XR^fYK\_A=HREP(.05&2KJJLR5gX?8
,31b,f^K\(IL5^8CH_^&G)_I=FS3U?ZSK5T]]aa&5SJE<3<H85+EKEDK^R_+f@/L
GQ0HbCI60HMW>LH[MLa7LSP9_.XE3QIX5O2He>=W;4cY73?[0TQ#:B,.M7@G>^JG
72()a9gB]e,-EaT,e^6FZaWD[@T#b>bS/I@Fe]V-fTZO-C?JZWL>c]7_8/WW5H_,
([Q=:J.,+7YaE<LMO+UJ-g^3#TMSP?bW:@ZfdD]3De495DG(eSY6c#)gFb),@FAa
9QIR?8S@XTe-#@SU+(b4C>6Wg^>.XM9Y_b@DYBeGd+Q6AJHPgF_3ebGU>)J=e,:,
@:JO7@eQZ+/Gb-SLZ2SE^@+@6c@D_>ZS,^)6&JWZ]86E1^BT[A:.aSDPQc;FT4V(
40+W@O.g?=2_:CWM+V(BJ8;WL;0R8L<E_2KR;K]T=,-_#MSS),/)VaV1NBE(1WI+
@2,0R;Q5J/(fC[PV1QZ+,7XPc];Q4/)NAQ(J)D78(KaTH43D-<OP8DVQeQ2FZ</7
gMcPRU5FI?\:VKPc-]9#Q5VfJ2Xc4KCV+(XQM_c/gEV>+B\U+ZN6KN-.L[2^UV[J
[B[cKI3C@8CI#OAXgM=[aca76FM@^b8U^[R/(>(\?D\ORI80R5W]Q8ZUYOPEG,f=
82#7cc1Y<?CJe\KDf=?DTMdCC<?NKK.K28a4[@RYP^Q.V_bI:G:9S^W+6TeL#HeH
@>X]MS4M@J/R/:3]QOPO_#ASQ\+/N)a,SP[fY];(bN419&[BBQP-,;BAG?>ZD0]:
NJQ:4N>;5ND;2faM?H_9@#N^-P:RcK<C50RUZ/F+[U/MCY203WTO2BMcf,e=aR,K
OBV]a+#^NLe)RgYD78QW[A=LdYDU#H[PS8?PHQ4FTI(JT-)F7?fZNN-@fO2IW/G3
,8OBKGdXGTE7#M[JQ<c._L1HOLY8]d+(LR66GP6U#A8PX,_JU=H6NK:2P<QG?[FW
9T8TZKCCN2H8HSRZE^GMAB6@9JM6CQ713V<.B[+TDX<cE@VSA^f8cK]g>8IGCYZb
2+BC_Xe_8WZ2[3A\<@-8Oc)c)1R9JNC+M)3H(Y=GZM/T.Rf23=BRVg9)NI^?#&&e
egAW4YHUTWUOH[2SX81Kd-[K//,D(FP#EIF=^#IQE(I]_FZ>-8\-/-)1:)BUI>:F
3b(K3\Ab=Q^&);[FD^84:TacC9R24b^XL18F8P:XLf#=^F6X((B4_,aXbAb6&a,S
Q[I2V_YNf#@#B2,6K13V<=)]25@ANDHMPOPcFWOVLDPK[0?N][[#IB]4EZLV.HWF
/CIA=Cag9;.3VM,ER\@:Tc:8,;9A?.YbR(F/H(U/\U2Z09T9)b:VX6WOfYHPOJ-\
]/LM(5O>J57g0Q]e#Z/-1)40(7-0F]dEDS,1gBR7X+-aQF23QGZYT6M@Ef+>gP]U
+B(J>FOX=4=(C=(:EO>,2Y6Ya2c+8;WG-Gd=/+OQd4N?_BL^PVS+c\L>ABOJ0&Tc
P?,OKI)#](@509D3;HJ^UPOSC>)YH6[LXH6gZ)1g>bHXIIUg?D]];f-D/5g(D?DN
=/1TG4GMSe&UM.EQ\T/3HUFKU:=,)1dWT;)97-Q39bf29(B8A#&2dDB-:=S6Rb0\
/abe4YTC:gM1R&23./&CH0\H8b1/GX2+D6b,eV_dd@<<^eA/P^K7TO?1B\:CMB[.
J7/TG@F-5S#Beb_aC<EMaAD_=Q^WD^GfWP-&)=S[ZHFK;W8c\:dU]DV0cN8-aX1b
WH7a@f46.H?+;^UKK_6\7FR-GJIFb2F@eA=IE)J[/M?5_ec^^HUMA+<))(@7I8Y^
QA5T=VY+75]ER.=9P=Z39Qd=E3>=&+BKG?g9J-JP(BGV2G(3B3DaKf@QgR2M&5O8
0+Z]4Y1QE3FGD>_@);:Fb6J>DCg#/Ef8g;)0=74,J(4@gY3\69LPEF:2-VECY?;V
3UcW=)[WGV9\FB_d.TK-B<EXb:Te1[AS_WXL2=;SI]4)gHCSC0?2XM;HT-+]9V+X
8E2F&B)e8A\7>L<T8a8?3#c7RY4A-BI/0b?J9fda&BHVFgU+a:gYDYO1(?#2J+GN
cI05=e+@cM5.KE-9@K^1fF2GF1#(I+d0f\=\eOC\Hd^)+B7EUXfMPWJCfW59/fAM
KT^:e/]ZdWD)<#135]>\[aN,BZ]0L.Z:f]@F+N><\V:H;YS)d0A.TgM>/YgTS)#b
?2?GMQ/Z(N>8>7V6AB.#OUXY2.J1eAe&bZN90aJ]^@;5DS4WI_M1g56a0/DHQV;U
>)7a;dgL6X?Ec(.=Oe7IE=9#)BNE&FbHN,72EcFdCNA)>B+R.1g8KG4W/^b9Y/P:
4<V&Me9;7EFa)EJAMeUPG&Vd)I1==,0\ZEd<@9d7PF@#3X3V+24\^C=.&WQYUbO4
NB0?Ae-f@bF=Y6>MMA\1a;?8K0^YHcG&JN5)1Y,K\&/Y1>G8G4O3:>^gJ)bCNga.
b@;A0(^fK[7MI?_M#dHB<X\7OSSeT0Gf8:_\aPVE[PZSNV,QSeNQF<,])8;<AB:V
A47EeYE-OO@R7_KEK1dY5f8<2^H84c3a4@VB\EVS0SCS>.BDg_c]c^/WER[K(gMM
=FUPTC>\.4IS<Q>b:F9CRdB)eH(?FF.,82#_M#2@)?<@]^\.>d&b1S8Ed:7_7XFf
E:e3dL@U2M4KRIS)G2XYS_0H4Q?6,BVNKf@+KWTUBXTT+XLg:7:R5U41&4NC).48
V21574dH.==(&,_a57W+Od_fVJO1[O;WS&0@G>aU#<gGV/QgN)G2_7,_W2CG=2a5
E3^&aIX)]C5Y.0###DdVD<4,IgY?.&d/\.bd0eV(KR3.TO;]B,gS7P\WTF?RY&^?
&;])W0d]MS3WPO+T,:GYbH)UVD@A,Xd?Fa?=6B.L9LLV8c9Wd)(6/]DZ@.[CMI;c
CN[[B^\JQ\4Lb@(O(b^BS?XSIWS62>+A+U/SL1;MKAL/[4I-_FLRbY_N+_eEd5aY
OBY[2ER9T_)-_X\PD9RKM;b6W-(XK^Q;?5Me:/JVDZ7eCM^cd6Y7U=@0gFT<51T4
T_.4E]Ue@Jc\31G,f-,47W0@+6HJX0<>=Z\M,CL-3cA#IJb4YB[409:Pec2SLS9>
8,(.Z\5G:9I&D]?NWU]\[[(.2+F0BY:K8^LMb17]F9Ag-(>+08-4[;]W.P.d^1J?
9J,S,-K6bBO#_U1TERc/704M^[M+V(RT05R5GN4UFEQ[d_6H)<?gEK;&D^0O;J4\
GaEfOdI^E20PF3-S_E:>D\7eW@<e?d0O\b:;HHTbSM2)WOF]/<EH<gCMNDS.9JP9
bRH:c<>-LG#(QV>g9-,:5W[0MH/Z=aPKL?)beFDLQ1#W=A7;B)-6;[&QQC9c)aeV
dXWYB94H#GHb7gJ)Z+9f1#951.\JS:/U+M&Je-H@HE))R]9e>Z#HUP@2J_,>f+.#
J^^+c<D?VB_,FUXEN9UGeYLALO4=:S#@b0FfZK9[?B[ffb[N@Ac_f/2N@>63dDd9
1e3Bg)3gf3D#[;fXTC#VdML:ME)6310Q?K++f..b]Vd-bGQA0aNgB(3:=];PC@--
HLNT_MRf=3,JJ4/3.+C0\4dJHLDad3]S90^T>TJ:92T7BRCR=E(,<FS>S=X\S4S,
U6ca=/:10Nf&K/aU0S6RC5R^[3PMN4?I\S-YbLDaJ1(DaG)1b7M-BPe&-G?g>:NC
/8G#PYHNT1N^(GKWIYE_Mf2JA^cGY2+V^dgSA3fN(gI,.Ad/?1:_Q+6L4IfO]E@N
M\R>bb632EHR00,@cgYQ/W39RP5OHd]UKTGQ[]28JKNN<9N:9Ra41(0eN]_<3A<Q
@7-QcV1d)g61EQU9aH0CfBBC\DT@[Ba]KaCA=\N@\8G((_(c-e_eRf:^cH4Z8;6.
R3B63L3+#Y/](-B<KTaN#@]Od@=7QDXB04D<1UWCC86E\31:dQUHK,;_P:W,3N]^
)Q(19ag_f\a]1ZX=_\V[/)7]5:S805N4TJW8?9H(>-VeWO++ZV=cdc\]HD(Y+U[P
#B7,]BZLbfBWP4Vf9bG6U5?Rc5/2R?3#O,,?P2JS=A@/,&Sa,&BOX\/QUD)7>1eE
)C2Ze[2#/IWG(7IE]UE1SIM&5@F(75d0T^c_R@^+,N2F,ML)K1Wb-]&(7fD1WY31
RM#V,Z6749M&W4^W><g2R?JbKHK@=NH)_-;EM,#@b:6;+cV;)]Hd/1YSIBf(.XHc
4#aMGYc1=D]TgP42AFPde69W/D.a)]TFaP-TDbLOOd0JM[#D<G3:\;;[HU72ePBa
YY3\WbJaS>MB#K(J57O[Z>DZdOUEUB4()_c),cTc@;0&FF2AX&JV(:LeDc0INJM7
ce=J4TI^f>^1OD^9Ud&.7FK+\T1__6LW]4D3:2D]bP2dg^0Dc9OGV,S0d@a#fHR\
9_e,OAX3IEFa4f(>gd<-:FY9;M[&I&;P-T?>7E7IHHW@f/O\.dBd(DaT(P.ffDP4
-#UfMUM/-?5[>H_>Q;K0+A>ON(gSKW>b\9E\NScg1.TI#0aNM+:XDSP5P>U(LMgF
H7T;?NGXM-@b;X\@]@;6CHLGF5>M-[dB:S\6@\W:YC5^IOKSND-L10Uf)d=LVUTB
PCPMcP.T?1=RXad]_;6S]HI83)D9@IYDF-b-;M/fLKaJV]QX<ObN.=,K&aIb6\V/
Hc)FHge&WZT5NcKI-BI.(H5CTPQ<=]SgVdGg?4B8Z7;^@UEJ0+g?BLXa/1Jf8J.H
3>58HEc[0g](B^_=5:/:CQd9W^8-.a/+W@;8YAdG-5(f.B=PLC96:W_2>f<8g.]I
f:WEb3VMCPCSeULRUT\K:QgfYH]FQ7S020\7L=@5?cfY9FgaDeP2HXeG&YF@Z0W^
LbZf>1J9Ye:\0M&5281A@\9cO,XA1.<H:UfVQAG[-Z4ZTXH>g^b1D-f[.g^)6Y>U
BS=Zf00)?)XF9O3G[<B0[@@)E_AT@/]+GER[<B@(C<==KKP/0?11NF.7/1J8bA7#
UG5@d?W2V&R&>M(LU]3[^Ge^O0@EW]UN/e^cU608J/SG#JD>TWb5e&PgIC3HR((U
:1+8A5G(VGd?@>BQ^TWUaFHcU#LbP1FQcZ+4C_Z[[EPUMSOAa+=UK],(JWVDfBg7
PX78&ff_:?[8+//YIWY0P/(,cHIBB8NMJHU2Ea=KL?IKC[c5.YD:?80W>#K@0+B4
D-U()2#45M+H,SHU58fXXJC;RD-Tg6=W>M5HVW5,.:/IQ8Z1KK\ZE1PFUaPG=L?J
N7,TLL<5S&A+Tc+].8JP06GCI9WZJ+DAU&g.;YBEEZKZEX0L2:.5&)+Z?L2SZ1AZ
NKC@]U,VQF@Yc=WL?EKRZedJE/CG)02=V64R2e-)WU/d>VeM05-W9LVHfH4KX&_F
&dZUJcN3(6C;(.0[SM>9?g=V_FM3O\T1.D;>EecA84HeXeG,J]UBgJC-9C0K,#,>
,OEOMJXG5U3abR)U+;0bZ6d+D&;BQ0UO(R1<<N5RMR67^bgE(ERge2?&1#DM)0Kb
=O3a66F9FG)9<JBUKHc1@Q<)]Wf]3QGFfgX@<<XK;Mf1^^?44\VNA^QJ\E8Ycc>;
b&_2Q02FW5_D<J(4(AD^Cg>__KdAF@dd^L,B+Ff?X>@@PVgB2IJZ1950b8fScU_D
?F\2Rc1IZVT_e##(5E(AUWP-=R#X8CC@b=KK\,P/+,4H3C[VU>fD\dPLOX<0&eF\
_/7]+cR@V7JI7g4bXa+JUN;Z:K?FPaZ#//f]<CfAJ\IZaVgR1UPb,_dO3KaL?20E
IZQB@JdAVfU.gd]L8\V24^M#_^c\DJZ@8VOZI905_G;[Y6IA[,KVG#]>85b2IF@:
cHMQBUETL)dVIORO+,B?DT<[605276J)CbTVHI2CIEZMD/SYY_93:RA[HLaO_LB<
04>/GI6<Ud9O0-d=H+d)25B?MG4NdX1PU&PWA4FY((6@9H>G]R>6L8dI@AbYg??R
d,@.3bXSgFXE\>TN,\[I_:I5bIXb-ZUQJ+?BeX3faE0gW#NMKWTL5DI@YHc2]LMZ
)aU/R(f0&F1WDQLB2eb@fQ[,..Da5_bQ58OU=&_ZgZK8T,7Reb\DTHB+_)>[IF2<
b4Zc&P,^d@HG.ESGNEFIcgXdKVc:S.NO:7cA5M<-4QM+g&J#>.W_^7aH4-H+6P;S
PN]Y[.CZJ8A_8#B#Y<+e.SbY&DK.DYg/g((/@Y]Fd/<PT\[=@0C83Gc>Q+72OSRf
P028b^#O-V(I&\THgWd30.N6?,D233NS[1KSR_C]g\0B=QGb;R.0P7/Va?L-G3T]
E+7KdOZ0IOE/eJIYbe5ZNI.#DFeO?^X=#FURF.[Ad=^],U6A;HGKXQac#?+#M5UP
24ORR\90_E3b&MaeEd:A8YGVY?-:6CHDTdR1Q:=Lb[0KVE9UVT13Z+@](EfUNReC
F<[CEHdX7=),^_/BNK22ZGJ:c(_M[eH@N2Yb@5@-:G[\^\NG9.\&#J=XKg;94d3]
ZG3d1E.H5O^,)AD.+U?R?09-aC_GITP81B-gH4]cR]V2PQT7I5F?+P0AM7FM4]F^
YEJM^>:;V\44Sg#5-T3K#Y4B)-ZOgPKG#G>C@Dc^;/]Y<>BU&S<M^JN1@_Y<+/Xc
GJ/^A39Z;K2.#ZQ.0A(XVb@UBO=JCcF(FQ<-XI8K3K^17eVBRNT]Ng[I71/(LI1&
ZK>)[?PgM_B\6FR,GSa#9J9,_dLbdHeZ-E4I2P:D][O6[,0T/WVK60aSPD8U:,Gc
M&SYM6WXZ5f.?]P[5<>g)AWA&C?N=V0ADNb_K(@#A+bV.8/56#X:_]-aS#@C+MBX
V9Ua7.&686cK2FPS2NCZ:^NR8dTWLg)MQ6J-R@7P#;-Z^\3US+FI)/-49);K-6a)
NJ>@Pe:_0NEfT56L+c?PI//XV0@dGFG0X9&N#>4CBM,abgX(-M9LEP7WQ3=)6EE3
/a^BB^,e)XZ2T>11K3fDgZ3ZLL3fF1IU8:.<T)-7ECCbT7ZZeUfCSAUc00#/.NQ]
dKcNKWE(/5C7WL:J+Z]UN]H89D<,R<DH&7F<&JIWbM@Fa?SEIG05JJKH2\2Y):3A
5,J<MU,5SD1103^BEU:&^P<PaIQ0HJ)2K)3LIIJ;-X2JGId:/9<^<_I+5D+VKAeJ
14a23WSN&cXGK<eb3NA(,55+#A0Pg+^LL^DD0+YgC@f66C=C5DX)P122;A0#:X)P
&<BeF_LUYQB#]S\W8(C:ffPP@WU.NLf:D0N3<=WNEa)?FD&7?G8&?Ld+W10[TI]N
1N.)D.WS#(:9(Wa4[EKd7\0+d804D,YYHLIcP,^<]?#0,4YdLKCOXe1\OQM_;JS:
4C,DPf->Q-#Gd357]>WRd/acZY]FD2bTEJNNQ)HaXX@5DJ,BRML,M);@3D;\S/_4
@T5UJ_,I81EaBCcb]ZH=c)31,gceAdd>:USYJ7RIMG=)]La,g;LR+.J:F>TH/<>U
dX/1-8T4QZTK^_N\?V9#CObO>ARS515a>>]RYd3#+e>-g=eGKTH8]](K0@U2,4,.
3acab[_:0W2&#1\cA,.TMW;L<a\STBcMGW^K@5A@Ab63KP2^Wd4fI5ZI+ZW>e/T4
2_FF?@JH/@P=>:L7L(T7BK;W@a1+;T.g2\C:EW&:77/L;<WP.3?RE,XY-],4\Ye(
/\W.:5Rd?<.\W=;ORBUc?HVBEY+72c?fXOZ1=]9[&+PKENN1E]aE+&@G5_a=G09+
S(d3_H-D4(R^+ScWbc#?/FGFA9.6Ob9/I@#3(0Q9;YYE#CbG+V]I\3OK=6=aaJ5J
Y&5K\dR+ND]^?A_T#K&b<3S1FMIR=Jg:Q(X33L^?#@b;JNGX<QXMKOMGPQOXI?LZ
B@0796O.2da2A9P2)EW7^Q1_+R.F]6dF<EJ&\@28gcG\OY=Z7F=K-U@OXG]J]6BP
:OR;5ES.D12d.2Oa0aI1MCW(,V<S]TFZ:3_D@.L>#LDR+QM,U<\<O@YMK=D]86e2
KcA<&H/D9?969_A,CeAf2R6@\<]?&^B+d;-L>g]<Q/,=].b1PFAM/,PQ)>A[T(HG
dF,LCQ?\4d[NG#d/d:V0L(DEaOLcI[15]4a\K8f6_a\S2]L77(SUM^Pa/+#7W^#@
Ka/7Mg>-Zf8F,^W6eO5,..8:ECQ[KGa7C=e&2Y[B]Y,RCJ^cXLM>d?0]>-H?Ja\:
,5KVV+]9MI0a/b#>[^+Q23XX8/FA>B?3K0)e,SFC,abOS=61acXQ\IJ(O9d[.;_J
A9A>/Vb5g,>07M.^e1W=M,eNeO[@;/=d@TQTNUg,HZ3<?UYMeER._HDITB#0#?2?
)BFbd#DEd^ADE-QG\FV3Mf@bT&^:AU/G;.@IIEe3SG#(c8c26[4GB\+.gSG)DDAN
QfH&gG<R4=EL_@I<3FQLZ/,-OO@]7T8eYWeK;AK(Y+4U_L5B<#/RV\<O.UYN95(8
E>@A_LCdVA.\PfRdS&IX\YZ=1JYG&Z/M61X+geE7;6?MPSCX51PLf-7LA&c6[I=4
385I@_@NE8W?2D\#7Wc0@FMS74CPW,?,Vc4=/\fa^1F;/YEPPYP?@S(P0W)GD06B
.\:+:\^2XWdG.W0fP)Q?A+]+=3A9_E\@+Y28ZB=B(\3e7:)F.P]eRPLbW62@\,;Q
Bb=/4a5M++F7L1_;+1ZFTT]+LOHU#])V#/HX24IJR46V-6faU/T89:d6#(Ib22IK
1VPV=16=2dg,7+(JT[aMFBG,)WW]72)L<0TbVUMP_8W>DEb]S<;>C8fOD58UeRac
35d498PH=E9(0H17.-I(=Z:8aWDV7UIBH-)Y9QEHP,He(2Q]?D+3bL@_HA<bbMcJ
F<O+91WX3d/PAJc^<UaH[/Zb&Oe,1B;^A6[8H07H-+bLR<X_3:+AW[6bb?M>9O^.
B@OcI_47TacEgKM0QQ6,\&8VK@0aa[V0B,=M\2;4W+,b=SVW09=6E(7,BK.&ZKK3
9FI3OD/Z@D_?:L+:[b;#C-#)QH2KE+^cL_:;eFKY@#AWRBA;CG+G_0bKN.5\)G0:
=73IAM-\HN7QA=U=?7&LE&6;=7\C36a_LR3McZWg1R([)e_:X<M?,Qb.1I.Y#8ed
MUe>+@HG5@[PQ#O15A5/<N<6VfT3Lb8P(U@T^B]YFc6/_8YYYU4;^3CG?8QUAgVe
SP)a9:>3-<+5(.[BdL[b2T\>3>SZcL]XQ84?L(YP#>B.:&PTb8d#X=@9:MW.UY67
@UC8.b1=3C,,D]-S\,e#.@dM5>VKK#U1<e0--J+U6(LK1eaHW(#@W-eY?A>FZ:3F
3@9K<-QXNSJ;:]BDE#5K&.\^2RK0@IE2.5#eJIda0QE8;\VC:F1gUER1Vc)T5TFT
O=J?CZO(BQ+a2]FFb&>>HOgU=D7^eDU8,+3B4WKJ#ff0_@]+SQ6HP1YH,E)7^9@A
+_GC3/>FSVC2+//ICYZdN/g7^NZ&=E#CR:PbABFRT>=HKJL/W<X?XG>7=5b:T0E3
)C<8-PbTB^[XB8>]2_M2dL29AZPG/Z;VP@dAE+<_I/]NFAS1DM,P/T7>CT.:Z)cH
:SDO/##HBb=CV9;bJ=A#.2&XT-b@F&Q0T<WU&2]9.QD^>OfASW\EH;=AD3<K0B7H
S9P[-X_(YVWCSNI?cMCVCA\B4D:#KU9Cb#bDPW96HS/V=O4=J.gMO#/F4e[3HS[8
f7.?^_N<-@<FD^=]M>8a1#>.?+@1_3A44<]JQZO@:_eddX6>]aQ/0,XV(2PTZ-#X
F]#V[]J#^<\b-[?+;VLSeN5TR9U^-I^<_08W>Y)<7//8e_X]GH)=6-L@cQ_82;?Z
<G7XQ\H>4H7:4EYc0):cG1.4J=0E.GH)>d0ET/.T)CO^)=4&^]0^AR;WDXYdBDM,
S<J3E^cK6/Ye>)XQSM@XX^</R,VUD-A4a\[Z+DT46W[eX13W+LeM16db.1CUA(&,
3Ld2ffcTZ;P77\f>)HL==<_:+^eg^.3P;C;Q]RB,EIC.b_GZ@efPgR&+PTZPRV=X
D[-(c#8eK5P>Hb(YJ?X+8)T4+XU\^ebd2-[FW<O9+\1<Xbd;G3/Z6GBVE+gG/VK=
.60FHK/NgA5.P=PaJ=(1Ve^.f9Z.SaQ@L3Q57[AELU1+Pe/)SOb6DKM26M1GI?#H
\@BHaFKa]OWM(V5a6(2.KX?^ObM__J9+(?8)CZVY5[L6G]S-?,B329Bace?9K5XI
_CI_TCEV:g(;#faGK]W@]XI)9a@Te=/@(Y9+P;4&_6:1U^]5F,e\Y069[4SJ:-P,
58(6C7@_Wa[g4,]NFFOYBKIXfgU9-F->HE.DI8PLX[f&=E:@74I&&B#(B;D<8BJ^
<SVffJ55I3Lc+3e]\5=J+<PHWd^V-F?_@>?QLW,HH+5H#L_.?\]&&PM;e]K-F@TU
Oc1)<LU,QLb\WL9Yb-Y0B]8545(bD_3F4_#+RfSE9c7bbB>L8IAfa(V9>g-V)7T^
LfO<G#A43ELg;5Y>e+8K[PZOaT9N\<[KgQ8]<L][8FHG+Z&4d#8>1ZNM,g)L/HVJ
<8/IM=E#CTDLKe5:NYdb)ITLTSaS;V0GNT9<?Q?=E\+gPD:W1/(5J9d/3:LMfHAW
TX:2EHN[RHB^]5V9gfD.4=8IM@\<7\T26S:EZ6?7M-AdA)9FWS=d^TG,/d34)WU2
OJ<US74H;=XF?gOK;IJEc?5ODe>dW.PK+66F(K4TQfZDD(Q0<B9R,e#G]HSbFP>I
43\<^#H7/D?E,5:9PdOEUE9ZV.BA)&S)8\dP>]8eK_9.4I^2-3,NFKJ2f6S5/)I^
(aWJ<63Xc2@3)XY.7)@#aHeZICCF,E380eVaT=0O(bVC(1O7^5(OGNWDO7gQ^E95
<Z?1J^d\#<?/d/S?4=94NdM.d0X+G@H^KHRD7CK(7_[fRfPF5TIQE68USTT&MU^D
TC+Ag,Qbg;\<XXZ1McLP=#fRe&&7=^f)EOg.09<Z?H[@CRA@@FM\[e-Z),EJ8>PJ
)A(=d[CFWU:-2;<=+&EDO=_BD-13WVZRB9IQK2P)3Ag8I+>1TJC)C;PBa.5Z0QF5
__e#0@1V+CY===)O-eg[EE)gUBO?(c3NM709V]1PdSg6O(ZJ>fC-SM+N=\D2Fd+1
@C0]3gUUJP=R5)XFATfOV,>2A1T,FW9EeIFaWAS[8@:8;[MVEYb4Ld<K.)A26K@8
a83+LPZ\=EXB75a91c>fU[.PUfMVad)\UL\)b(A4.V@I>5[g:K_(YQSXG1;W-0.b
4R5S@)1GLVXR:EO-G65bR9:S#)b<@4^W@Z.541e<6T]Xc>VZW^\aG,bd^><#>6d3
?-c?8a)5^a)Qf[2;af)RZd8gg-bSNLJ4O/E1Cd7KE59gTWZc.8;T8TBKMR9^?)SY
Z?I,VLA-I;\fR?&,M=_&T]Q;.Z72^f<9M;Nd+4DN<1OgBRL=1#_)/b:)AV5[Q.SV
T<2;6HPBa,O#V4f:a1@f86J=.S(KC?Y2&>2R[\bfL;#eC)T]^BH;ff9^5Zaec;=U
PI:a,21HgFa,7TB^KHb@eF.2KV:[L7bL1-BXK8[8c3G/AgO]906:Y6U+]^6V.RU9
Ag3E38=MBP_5M3+H\Ab)A7/C;DNWK/#E#+S-5XG8ST(Q8SE6/&EVRG23URD&6B(c
_US5_V_6BISB^Y#U@5&>6JVWJ7RN61dR)gQMQ=.DYQ3fGAZ>IVM#1>:IC]J>_8O+
;VSON>_-P9?]__(AWb;PGI_(1&YF1@[0<2F>W#(0DSIUK4cE>O<8e3;TM_#7:855
e&.?F8OOX1HA^YFb#G&d6Na=N]CS6T?7)NN^;;UfN7g9(5X;4EZ@Y3C&\NVZ(c</
[gF+6/^GTff)=dM@>2b9c.D7aNJ1D87)Rb?1+UB?V.A[RM1#EA2U1E-R7Y]IZQYN
3?8GJD?:3;d&.=J;g9Ma@:XM,H3>34ES,DBN.7S+f#YMVGZ9YQ]I#7CU8OEd8^e@
&14;Y;O+?A34JVD+3N8Q:JPc90/OGAE]3++\ZgQa33JYD@A>E-_cD]G&F?8P[][D
g-I#d)Ab04U+0e>M0AT0FIAMf0/Z=NW^2#788\_6.\GUY0B@N^+WMG2B]PUW161B
\?OG3DYWUJ7XI4Q&?S>cDY+_[&f-1EVQ.>4O:WI\@,X/5Z7--;UBNe(Z,CEa;T9E
-V],+Y:-:6RYKLIJAeONKD-UCED0Sb&[W@),#8Y5K)S8[AXG7I84;CfH.&&c@^Y6
_@gg)BKTJ9?QE4Vg.1P?7RCB330NT728AM/e9^-aG/.9+/=3R9;HWaK89^,g60).
Eg_RVegU8fEL0E?L7HRZ43I,AZe;cO?#Pd&)TSB5)=\P:fN&H05=@T8gfI9N51>8
D.2N/=F_18QBb^23e[S@E=EJ+@[2D+cL>:V2RSgWMb.R^-Td0I[3V7;Y,G17dO>H
5;66TeAR2(g<^=AbMITRe?&fcZa-@9OX5^O.3F0TPG)W7\5-UKa;2T]:VZKcIFJA
\?&/:80OV+,_7MKaXbfLVU_gEC4^0T8W0]Ke)5:Z^a07P#6/d)8?YL[MT3U^?RNG
.J2HQe5>(/=MI&f.3[;03AeO:We0]B@K+<@+-AIN4TT/,?>b-AJ=JMd###C.#J:U
9UI1ebX;F@d\G#TU_RQ>\Pf;;TZZ9_\)F2#QF_c(O?O(NSgC/UYN01Hc1RTg4a\1
9DN)9,Nfc.,[R^N^ZLXUXZNKQ65)H=^Ta([N)JWM7A&CO3J0.36F?@HdI8fGc-0C
[-IIC[PZMBKSM/^+4H1&Z5]1RUZCL<RK<B6g-O4R^ZKM73RaXTU;CYfGaZb2Pf?M
LA8X@O>0VPPL?2^BbaB;E+(W+P[g1.cZRA^H+E;G^JL#Q1eT1M),B.=;_H6>AN70
2fO^V1/9#8:)K@VeN.D[F().fN,]KeSH=>VbU5+,5QU39Q,?C3H\5-KMf\\&_.^L
PHTc\K(V4X[&H=WVUg9Me<O6>O#g0c7P+G]>5\WTQ;IY&O;IJPOAX@&@ZZLCRJAf
=L92RUM+aB+S;@X;U>6cN=2Ve8E6<UfC.7Gb:[>aN_(5-8N53M0+bQ(BFGgN.:J+
]=c&[=2Z6#N\f^A\5/cAeHA[S+M9&-])<F83HQZ<21NBYV+7Db=SO(+WV<IE[=e1
.9^@]PTbF>71Y(d^_c038J?M@3J&I9?:eKdg6@;C1T&Ja-GM\(Hdc^<Jg/\DIOWI
ZXLY(,ZMBU2M:Q<>R7bbJ3AGVWBD-EFC/YHDF:(?O/6W7K-/KOeV1V5F5:2f2W72
?-+5(8;VAR160@XC<-CH</WKRH@15W-7KHBDaIU9^6?A.O69VG:P0:A6X.BAJ+f>
\O^g&,M#;78b&-X.7&GR6F=X:c2.SD>d^6I1FK^;5V\0HY35.BIf&QK?E\#KVU+(
V:;?A5#KLg/P,Z&/LN?^CZ>6_K4/JR&^@D4S+g8B2T?TGdMQZY5_7QZF\M.H/3PM
CJ=XCW+FC=@DU.>R4a<AO,8gf_Gd>a?GB)&FYc+bNI3&<&Ca:EMQ8.<d6L<#5fJ]
+WN5-<Y990:IF_Y8,R]U>Ca(VD4GceO(D6^M):.&L(OX624/\LA8ZE,-HIE@\F/U
#R(E.Lcc>I(f2YGc\b(PI7aEHTcbYK49bUZb6;6C07BcIbd.BQP<Q4L\[A.=geCV
(#-:+PbH:Y^[OH,YB,YJQ?A4M.3H_LHFBZ#LP\&<H.)[)N:(aYT62B953VAPUB>6
NKT0+fF>ZSU^]0.-EEB&c<_KcY+5ZfR=^fAI7b76e(4c<e.(#HYJe)&?&)c8g1I>
M6<XLJB@7+L4#&9d>J32b8I)1=N.BCU<9f<U4?QTb&0V]KL0^>9CaE8-bK?6c/?d
M.7DS+JA=U&;3933FcDH.>T6E8Zg@&@X1KMe8>5:5[F@QAg\c:ETWIP<+PBI,Gb-
?g-(8,<K?JKXK=(/V[X5e.PH[#ENa(@S#\WfC/J1<Y3F_O#7<R>>.^D65;6V-E_;
BI35SIbIgPE@0:3#?fQFF0e:AV(V.E\E/36@@fH[4PLW+dL@UKNC54A&EZ:Q)P.&
9,L:Qe+N+WH<?KJeeb\V8H&25L&XfT-I5>]SY,?62CLR6gMfd:VSF[-4Y;>UJ=JG
[QHa0[1KS8e-Cg9_)D]-],=cAI)39Q<GQXHUSH?]MSFA#8)J)G:H_0:gdG@FJZ5G
6(D07=PF\0BS,XD(E/4=-_C\;IcV)cDUIEWIK91X8_LTK+d:R6M=HXbLQ<//S<M:
\FK@5c<9W-NJDa-M3PI(OC#K[>@B?&P-Z<MK<ZC(X_SVMM7YZG:8d?&bfM6V(88>
dMaY).fDd6>T7d5CAV:JLP6GC7<RK:7OGc;O9>_SFO.GZacC53?.e<)Zg30E?)QE
cPZ15&+T[,62H3AaA[V>d6VL5M5D+9T^aY#,L&&[1V,#Ke2eQ]c9DTTNDKZ\gbS,
#S2g#+QQ.MAgf21?X:&56FG?QP>b)]@Pd4&-05II_XVYf>T7WIMa+ZF>XSHD3:+B
/+U:a&da??e8+A=WMO3QBW9\7c>^b[XDaJ+M(DQ9Y:M-8/SHQ,K2F19,[UEa0=@R
6]R(ZeKg+4M0,Gd\00U5T;4Qd51He7c<GVa(-SH^0fV:28>\HRA9bf\,899A#5IU
#RODbWHMH=/cL-_.QTa04NeHVHbPF56MWU1g[WVJ#Q=FdA&3(f75BcM.;_5XfY>^
.P?dg/>;Q]<]<&ADC]_#>Q),dEPL7_T+3aTbY9LMQ6K[]HCIfUde-&?_JCJR]+B+
5gLgWGAgdKTYA=,FM[H((Jg@P[N#,A[<=e]cJgWgdKgIE+G&]0IKUPA:e,\d0;+J
.Ga2(.LTg1G=ID>G594//?a/S@W8K^^X\#B6g0#2?^?:_[ODI+PL0SIKUfBQTHPB
RXCOW>934.Eed1Y4YBIEA1X-4-)Z/4HJ>1,+9SGeQRCe4a[9DVB,&LX]c(A@3-N#
b>BaT\Z1:0,<M)gMHd?V1_ZA=)<F#BPYN369,/.UgRS]B0Pa6NC#Z?/170a]+FfC
)c0NQdNSP/,?B(<QVC2f3ETIR9[1\O#D[eF/7YKPa\g:VKdD/4(>YPX6;<J)8@5E
eOVVEGaVKC@G[d6FLb-U>O#93+A.2AR#O^.D.KE8gSO_(#fFH9_@;FMUYa\,/RI_
dH3aD?C0;Z3g\d-gAPSM@Z;I[;F>R(0d6cOA[9Y?OF)\>)Fb<4-(fN74d>@2AS0.
#\QeJ^KB64;\.UO01U)d.Q+7VfTYH&2\d=VET-^60-:67WGAeHB:Ea5eH\fMQ-;c
ef#5KU2>a.=ZAJ8=:XNXK.>Hc+X6.^,@97S1H)7OJ2a)8F;acAP(Qf).P\MP/1Re
G+<e;F?a)H+3dKPF7]/eF>(VB+V#8T\X3.IFZIC3&+[L<+?3.KV^>ZNS)Xg6NO+c
@8#^-b[TeNJAY<9F(DMAZ4<LIB4&6IEYTS1R=7QSAP403YPJPQ70&8FIAHBD5d&[
gTCY+6MfWgVN3QI:4a[(#Y^)Lg:,K@I7dRXbD63Iab5ObC:22H91P3POJLSCL-^;
GPAc87)L#X:LXJ4&0H\cF\+[YE0DAeHQRH@:2U/(J)ALXS=^F?@?TG?U;JG0-D0g
MHAd2)b[N0](QDW;)[;H=DAS3JOM-,0R]XKFWK&94(dRT^5ZG(K<>K3PQYdVZULT
7<5M\gX9.I;7bJVYfDRcQ+A+LV)3XQ_P&](;@RLVWW6:Tf4Ce+(LY#ac;U4e?#V8
,7E9YHLI-OgeUYF;dW,#VQc5G<:.A#aMEcY69GK^J1.MG7/(:ZF##C&6R&(HJbCg
2H\VL,0g\8:cR.1/C:Z)7)=HFag#eZ(A?9WBIbe5,57e48(BTTd8+S(H-cfCU(R>
8T92/-7SfNYaU0G1/24PUF_TB[+-R,EM-[NBZ@(a8a20WVC_-3(K6@=FdIaFRHIQ
]2L=WUS0?(eI[0Yg.XS6(#:e+^Z4AF=N35^1B<a9=@72,^:a)FR^;eHb--H&=_9&
O;0c@VbHHZ#6948M><1B>_\9MZB+)Z9&dgO^V-/NL[\-;R#M(D18+ZfHe^T>CMF:
ACS)4PUYc)CR2>.XJ@RT9YRBQ/Q>(\.US01N[_?XT9K?H6E<W/cBbT&UWRG;LD7=
#=eK)/aH]]f0,?@.^D)2Rf>a(Lf=.;1)LG,d++X48b1A#5BER1^BDFL,D7@g3XNc
;8F)4FE?-\(R:Q8R/7\M)S/G[V4.7YBONJ00Vb\BeSgV[?]>^YcM,YFW2>2\IME/
Pb-/&e[f.UVeb-NY,5e74E)H=B)5(UGg[#gJ0=V)H]g^dG9\AUe8/_OGHT_HBAHf
Edg1K0Y?f]D[3f_FPK-9Z)<9Dg?d#[DR9/Y3\f3TY<bU_Pc\&8R;ONMdZS_D382Z
2IX4(cfTD+FZ5(T<dI/[J07M=4MXEL@9;C#3dDLB?O#,Z5(]N@Z/#.=3VJ(Z5dP6
>=QB7#Z@G@NI,:L\/>&+fI.a==Yb.^\G7=CU^Q:L^AMZG]H];1[F/7FSMD)EFe)<
HTe/FWc+5dCAA@cbOc4b(MU=&444G(2>D]I([CcS5GR/?+SIP]A?XdE7;;dacaI,
ZMI_ccWNGf1QVDU#H#HAEXH(NBg5c/-G8H=eH+8LF_+:cLE9-AKP[UQ##-HQgR=G
]R-:PKE1DRK\^@1\:.&QE6O<O0:Z<=Ob4be)_6JdFOd:VT8O_cd;3[NIa/D+VP?-
-1?OPIgZ#5-Q4YY@RX8B0TDU(g^)M[bEg+12(T(K]K1gK9?UJJcV=b0M()6C<9Eg
Ug31a24]-4R86+=60IBc,Y5A2T3FQ9ZY:E_a+[,+DB.LSFZE=8DVHF(@1=N:DZPg
A_:)dC@XU?PMX6P/3fbf-@QF&UW:-6YBEG))2AdJ.R??<,;3:ZF1Bf#F?B&?a<W8
.S89W:^J,#OgaGgg]P;PD2cOc9_1RF\J<3L)AU^^UDYKMK<0Z/[1cP^EbNDS\Ufc
93EFT5;(PQ5C&KZC4d4UVb,?#BTPEbPC2d#YFA>Zc3AZS46,YCLEZD_OY0^H-J1)
3BH4.69\V^(EVL9L2H>^VJV-Y.96\<KJFd)0fF&F;e-f#\D.WPG1S_e<5#CX0D2C
/P/a[_^)MH3TOR4Jb7];@Wfa:NJ[TSO^]_OPMg]#:-4e-a1=1GL,-\gM9?eENaIU
/W05BF@T_=YHU=O;fc[]9\e09[fH;NK(GB;U<[b8,NAWYK-,A^CR5YObJ)-WFc9(
c&U7C=bTJ0TBA_,DU4ZU_Ld6__P/e;6/\f?9]DZ9TN9WJHTAC^c_[Xb^H1_P-5dK
7d<_HK>3R.-4E)b=X>[4;e+XF9+U(Bb1G&cFc[&IbH3,?J-@F,(ES3EM7:/&@E/#
[#K:,Z=B>)3[a?T.VPGL4Q9,+AL.fC4<XACfV/E[:aFNSa;,0+\69M3OZH1V\GYT
]@&^aQHYdI+UC1>YRCSdH?c&NL+T][Q?KbB9K[BA3VZ9@U^WQ0b.),_]+TD5aY_N
R\_HcL\;d3)UADEZK7EQ-NVd(FY;b7/\YEVYgZI?1ME+CZgaTF>Q2S>bF-LL&3f:
43O-dW_dcJ>1X)[P;9UUYcHa.?LB[d2KR0YBEM5P,LYUS;AFb<8gdfC\WHW5+dP\
ac=f.Fe3\U[J-ZBZ<RXPZ7&]B=^10YbQ<WT+OVKQ5^P22+^&ENT11N(M@ADbREc]
F3]1SV7&CWA+c0XP>.2S#)agLag5^_5-0M^[(4G04dXFd\GP.cN0EabM:WMZA[_M
DfJ38K0793cOc&?I5VSf+QR[,_90Ce9KGIeLFg<C99P,6f;2TA:FDE57__JJ_Zfb
&4Q&0&F_@(HG2E^0g84J?c,ND7R+Hf.A_,/Y7O0f^b^V8H:P0C[)K[0/;=0e.:H1
fUR,)DC7>2Cc=X&,S<L(5X=F@_JdSfEYRHCP)@V6+H[.6#L_5;+SEPFe@0YD=>^>
RZ;2P<]8BDIOC3N5Xd-?1d,OD?OWC#QD#;g+gU+&>3^LdO6IRR+QF#:bO/[VA@B#
_M4dW6NgdJ\C@O?.R3c0]BVGXFZ]-a.K=)TI;^#VTBebDMLf?MA,U4bXGRbG37DD
d23P<]3_dcA0OZWF4R#20#GQDKf7/e;5F1PM<E):O873_(C/\ZLc</W68)^++Hae
<6M\@4X;K;#-<)06LAO:4^^-CLO]\/__Ud<+=Z8PB175_G>:_b761/]9B7WFZF3V
VDRM2]H[.GFfA0ZPVVVXK.)LEL#Z2Mfg<6/W,bY?CccV@e?TF5]V[0,R?d-b6<5L
]4=3c^D:4QQ1+5\F.V+aN-://Fag.bd7NdBdP2<66XG8:HeFX6:5eeb1UY13YG,e
(DNC;fZ40Y2N11K.CJ4=66&?GBX:71=PAS^+U4f\gF90@205)P@fG,6bY(^OF],\
1CGe>0E<1c26,N8FJYC(9:MbeWLfZSKHXLfEcR;FKWS/I.PP1F,HW6IXO#JHO5fX
ddA<:-+W/6,I4B<W6[R-&+<3X)9TCQ4;2C-/V5].)a.-;TD57#K@RQF4,@5:2LRC
=eH8M)FF;dPd<=J/J6=FNMV#PLNa<><F)&PO3^M,W7Pd8DcROGdJe?LR\SG/.8>D
R9PP]AA=9C9Tga\9HgME,2(f261)O6?R5_;)/58fd+];3]add+FNeJ_(BO>B6UK3
PSKI\;H^/c(^WaP#^Gd9\e@H2JJLKZ.)=C>;#T;ZA+;J_d@#[I9QFFP;R[6-)gb?
>[0X\g0HZ^?[HBe<7[ZH=MA@/8HOd[UDW<3SRGCfHQ4IIKUHNB=;U<W:TPTA1O30
,2)#[ZWeIN@dM;WP9UE88R.L5^+LfCZ,X-&0<3:>aN\?X_@8).=a[a4IH6gE(eA9
,6(:+?=TS>9Uc;P_R,1gYV2LUX#P_JD0XL.4Fb=TX=BEUJQ/D/^>8aJPWS^1b1^,
0a<T\bNKe3I+.G;TA<=>ADNI?Y;UacZ:/RFL/C#7_7Z99?5BY)SL2#UgYX/=PE\F
+GS#G6OBR^.J]gIbB<eGN.,ACG=fA#+a5W0CI]U)&=>fJ--<7S/D5>(RKUD+XB4.
a:EQNg\1W6.T0;>IEU#]Z9]DQSEN.XC@WD&O;X&C2\&fJ1RLK5Q(^Z)\)X0MRG-=
#+;+aT+FW@eP9YF(d@698:gY7\SKMQ<X,b1S560gALAKUA#/+GUf5QaDB<IT4+AL
[2&K)[aLR7C[gcS4JKX>5<f+P@c<C6,aPL:K##BS-VPa5J@B=43J=eMMS[^/C#f_
#cIF7K.fX)bTdOUMPCeJI?]S6-ZVU:7KLYABS?>1ANag]15ef],18SY5JW78VA]@
3gR8@)ge/<?JJB;DQ64A6,1g7KYC/M8F[.O^1L43FN/OgQ\J2Jg)=VJeZ8d,4@2+
23Q/NaSVU>)8X.HT,9,JE2+2<6&7Gg02/3ea9ZJ@+P?+],/2T-]FQ;dZQfS3^eN5
<&SH2gA=&[_.-+MN\X571L4AY&(\XVX[MDe>gS<B51N,U=P5<D=5(G_;:20YKK:b
-UBOTR6&d3e/LDK:/8)QA20?H?R)QI1\R]KY1W&ZYg07(DH5+16XC98_O2;9A8\?
?7+,70+fA3@0N8CXbPcd?N\-TT?f6A8d^^6dH[U&<F_=S&NY1=+-PS5S95<;a=9c
YNd;@-bLY?3^CO:U>5NZS?:X2<0:_[^eJ=B+52>MNWIFRKU[P:,d\NAecP/&W]L4
eYNLP<B@SM;6Q#-&]G)1?=RB8cYS1YXH?D(XaeGSR^BO6_&R4<cH@P_&gGE(g2BD
=.00@[XI+K)+#GGfURb-^<M>@?e:)9>#ZF+;/d4Id+,f3G5UA4D8V0+U=SQP#K;N
+LY\E^]#gDQH<>@:-c2:MW88[HdT,.OgH;)g])1A]66^@O+Da-g]b1N&8cR8C5M7
/B7W3IHGR^eX.&5T1#PX,V2.R6>-YfD=#&F]/L[?FURcHbP6A)N?@7&3c=C;@Za,
K\3(R8]KH?>,f#UI(?GCYe/:PH>^6CJ47c]&aFZ/B9C)S,1:55O\6:J+?BQ5PUHA
IIU[)K[.4N:2MK_f9I<H<MaY2#IHHDLf58SV:-/K[7fNBfR=>25E<&MdeL5H@.1P
@K[TGOSYMG/VSSNBVD8U&[2=1>NVX(2V6RAL(-f<W5HUR,d&#U5Qbf0Yf-2=OBa?
+X1aWOJA@KKHa[IIId?:?+JUB)9Ge(c#&0YL^U4a)75O:8F+5E;S>Y9fa)4FCN7?
0d@,X4MX_N;,8dJ1FQ.L0-_1A5S.//\5]Je07D8VE>afI0+;JEH4g@06E4I32QCX
(c^_g6J>21(CK8U;&XF][,acXX+6]G<7MJ[;S:a2.[KPNESRcVM6P=KUQKIYU(eb
N_C&Db(#)E-ZYWg+D_/b3I=AQ051c>eTd-L>B32c&XZ2NM(U6P;RA51S:>H/,g.e
cK:A=dC[Ud(@G;E4V1&C=X&KC5-A5O(AeDEWcK@LUZQKJ:&>7>>.?91Y0JVI=E2&
CcE5TbD^TTdCZK_54YZ\gSP=P+MQ+]CKB0S>M&Z:_VP4IXCV#+GK=>Reg(-IZ6Ed
EK.RBNeP1TMPAA[ad92-@1gDR/3&WY\=R9=79VFQ42U10O=b\?Red1KZ/1Y?_K4V
55R\;A&IaIBOHWZ2?[PLHBcbHbPL##9S;.J+6CHe^Z[F\CY&<1C38;.UT9D;9@(E
48ZY@4K^6@\D2bQ28f[7;^&7,59J3dBfdLJJ)0H10U.T0-G);4U.VL7bI^00b9Sc
5^7@SBSCdTESG-ddCM\DQ\4SSfb.cK_<;X=^]NJ@V+0C?Y5.SaMe-P]eR9bEDG8C
E@3I)NIV)DAE3bf\>KE90E:/X0RW3Y]CBVTT84@(4A\d9O)7R5D@g?9c[)\3@IZ4
?c@:DNC7\D_=<E6S[/=ZG-7(8C/>R7a7M,92=GEAZ,C:a462@R#_8PFP+8FYT?(1
7&AIaO])Ve_1:S#ReRIcCZU4aDbO@>]NI5B<a);MDg0[+R;Ta)<D2f[=XDM^N^b_
L[<51IRJ7D9g/8[b2=]]#V1Qf6C;>LcT1fS#JO<d_6dUHC60Y_VZ>Dc^3OaJU4&T
U3bg:66GQ_S#6=d6(LGFb9,1#f2S0/35\W3g]E(;fJG/H,6U6E]9^-Zc7/R<E]\3
]ZJ_U8A<DS03LZdc5@?],<>ID93DRJS9)?PA7ZF0a)AH3_1(3D>f,3([=YSD2BQN
3_]/Z8G4H.a38TJdeJMLA+QC]W&Q\(B+JVeQON.QOZV=S:R&>+XOHQI9[:>8Z3,0
>[7K1E:YfU_GIa3[&gO1NQ55-((41<CCfUF84,(5c5g0Md(cRMP5M]5-<I8O+DWX
6Y8&MZB6?SQWYM62Oc/SRAcY<38Q0&7/]NIcF\]-DNP\]+E-MLK(^>bVQ]=L_a8c
0^O2c)7A:K1C&#e1-?6/C-bE0U2>__ZI#4/LUSUQ(9O]?Y_<C&5]68>_&X2A9K\6
LEVMQ_deT.;#^M32AU<a<FQM00K#)4RZGeK&3M,B<7(8&IPHEeYC@)gIJY\fa3cR
eR=):gca8dG2#W_B,PcfY_ZgHaP#J&]U:2JC?Rc<PETRZJ0DRK>MA>UQWR=-b_DV
>GeDaJQfY:/f@<35SWGVO/^+aOOU9I);H8YZ[K6=U13YHLZ/e45S_C+U>dK:,X+7
I/bMGT_deeU;A&(1+117C-c+,-[a+T71&d/+#SQ=g=Fg.<3QgJb9GZHe[f/8W^T@
JDY7I/_J??VDCX8K&WP8DF\6g\\fR>YN2fNN<MC/#Q)X\1Z5_NcdbIH6FC-fL5LU
Z)UFU=H)HCTOHN>GEG]ZFIY:?/7J=Xb_G\[_[+6;XE(F.>dU,f\+>]24?[[^).EQ
6[+V7f+/-dFN\4\Z][?X=)Z_).e1.?-V.065FD-3SF]<DMGWT\6SaEX(UQ]<&W<f
S^OGK&Rd?58CWA)b-8X3>7g)X(-5-WD5a)bRX?(N4=W7E17,LHEDRCH+IKYG[2Md
C1De^5NYN.GJGBgcC(C&3C6Q&2e)fNf1@.R:G53g\0K(Ed_BRU1XT:g7;934:e11
gTUa?+:45/KMPJSL,<0Fb9@)M9@:;6Y^TUfF]U^IHebA3F9N5E#cA=-]:5aNET1X
X.FUW/3?N9)V@@YA;()CWRR,Ud=>>LX8BK@=\BP[&30G</Z6[@IFJcE#8\58\70J
eT3I(Q@F=^[/XL\D+5=,EKTVICJL,R;/VVGG,dSI(c.d3JMW>QJ4<X8N6[Pa:,4Y
^C;OQg7LDEZ<NFc@V:N:e_UcLa&FM-Y8:1G5I9#[09Z<X:Wa2(?BX(b[SSTPH<Ud
@/453EQdY=a1eT0;Be;#V?83NYWLZ6g+,1FM3(W4&(UH-:@TH@C5g-5&gQ2>ZR]=
LVQYP6;8(BX(955IW8e?Y=#<^2[?07W>K3]XOdS?>YG9-)MN87.8,)2>5A<<6,)E
:,e[1b[OC\^7F1c6Vb-M?eES:GFL:3AS03K722^PNPg6KD+RYHU8X?;#EgS1(4g4
Eb1ID1<Sa7-7TAQ5GV=S/Z.203TDX@AIO8TZ380-8JUd05c/aQC?gX//DW6(],EM
;Gc:^4(\UPRRfgFPQTXP89YD@4IXB;.=S=S+^>W]XM571[:W9O>A[LXQd=@4T;d3
G#;#&K9JC/K,Qb6U7J[;>EfA307SFZ(>P01Z(eUBQEBLW.D^.HAFJU^\&-06,[Q,
e[^>eB0^L>]0M2BYX9>^Rb(P7@B+;\DEE\;fePd^+Gc(B,S:3ZA+TA?&N3]gHDeA
<Q&DXRSI0&NC=<KOQ(F,6]6+V5UF2b=::ER4I+#42gE<IHL4.97:?0T4U^Kgb/7G
\LAb\BZVMUV&0PFM):L:Q@=LWQ6+M9J#.Tc\+S=GWFe)4V)PMC;V@S;?,,S=;Cg]
bSVF.DXY0X?^],C56=;]-PUaK1.MR9&fS=^H4[Cb8Y30A)O,fJ/B&72a1=<Oc,/I
e8+=S/fSI)HL+?<Jc9M\T\^7QQ([-(P(S(II2IHD1[e7KT8D1SbME<)RT\8477FQ
b\)c&>>XPD/[GDY[>6K8<@W)G;_P9.D<(9-BO(Ib[E<+:dN-@N(;1_J-96V3=F/P
GR2)_\b(Ae)I^<[KKg<M+2.M=O(,RH->Nd]T^eLJ;e09PMTH[5^]\P2UK=:6=DB+
-=,ONWf93A1YGW(O;L([[5U2A0=>CeCK_#LT&URf+:2\[;3^_[We^7(Mb29C?+/<
SVCK_9N^;76/H:;F)0+H9>8OQ/B#_)TO2LBX,[=VW3_L>.a=_;]C\,&WQb>_5P&-
3b^X2\D-8DD&,&e7W::/:#N:WY.^/b9Z:25Ba1YAcZ@XI=P.K(#25M<F([52#;A_
WT0Q#e-/,SW,=_dbd2LaS,(XaUXgOE;4XJ#HV&5W\6P7,C@Zc3=0D6Wf5O48+-)Q
<59_&=QV&>W7RbgA4c8d&(&-N/WI,3EL0FfM]&-R6ZXQ?^9\H7EID::[ddCc0Z0M
2<g/2BIY_\I@Z<&.A(1\8+=d@(7-ZDIg#e,TdQN@a]FWZZF>]\9TIS#)F?^V,Qd-
1R7Y4@>V(>F-7M<Hb#2Q@NZX;\F2KS?4AV)W\Q8EbUfB(::cBC/-U39,>VXLG@^#
]8Ya2D7MSfCW^0,L//]5d<?Y@73/,#=;.L^[BS3,007g9V0a&LN@J\d?A5PK^<;E
_Y8:U>8NS0N_<:>]O_YK(;Q8S=8aS4QNRM.2H\LHG]:f)eYAbd?K#Ra[A98D1X/c
.1T[H8_@4S_372(HGM];^H(]RCdS)68<FI]2cfRPO5UJ;27,Q(YT26RI[GQ/.dO3
U?.ZbMOEgbQ8X39,7<W:=cA9>?-(5_UJ\I1,)R[D^/^b(Z=]8.Q51M+35)5KF[X+
\e4#\2R:RK>N0VNW[VLF<g]DB,5W>]<F\@V8]P\Vc))19[./0TXOa)Y_D1IZ>B[>
DM36-W<<+8@@&UgM.[fKG811ec6V9Y,MMO.:1D\<BN&TLdRZ#_J/g1B<1J^^R._K
FF2YgS2JL7Bd@IRaR0:_NQA7KGY4?-WS(C8WYE0RHLAf7AHRXE3@,(CM_EO1PFgE
12&Y3^KYUNf@0aNJSJ0=PDB5#Y2#)TXe9eAMae>Kg;2,c80=?AL(57gIZ3?0]Z>=
eU#5ZX[V\T#;:^57G<?N8cHdQJS8,J.BcKRa7WV.A(J_<Ob7E>O;H/PTfMT\4L5Q
]3G9^VO4Sg?]@H-,F(Fc#8\ed(N?,?a1ZZdHTR&J#U1Y2KI(2cc63MB>E#@:QDC7
]g^fWC7+RLeF07e62dJ706@g54>6O+Kfa39EUg7L[BUeLW\dK([80a(-^FL@>&gV
@#.Kec:ULL,YdR&Z/@F)(TEaHH^\7I9gc;8eOHLQNYa7:1DDcaYY-\U9YcX)/V=e
WP7LER;BC35=1O[<@/[SY3DA#[WEI-?D;]fB#ae^-g+ScRDS7/9NJ#BXSDXc2Z45
5CP/U-<ND^B4SH,-X_d]Ge7:-Fa9W+H\J+-+0.:QQH,OVDcD?0)]Te57SP\Oa6P=
/A.Qb&IOeF.G;@E#4ST[b#B\9[AWFQKW.ad:KYD</3eJ_6[JdK.+A53[4X3TPHTQ
d8T?97NKV4P6#6(-;:J/KFc::@9ERE&]^Ed,^fdE\=;K1-J3b+UFVg9CJ4.&<6dI
HR.(K9b^/d9<LL<?AA&J7Z(4ZQ8T=9cU(gL]Oe0;cFb<5=S;HgSA]A+_K3Re2]EJ
UT\V19/7.L7JPNJ95FMY<PX@;GHPc_5]=+#1<TI5ZZAK]Z3WD5?WKNbWfXR2-V[,
Y/9VcIGNc&>XK[ZY1V[L\2W?GQb;<>WcVf2OZ+4V]V5T3H5M+72M/)8>cF8_]0af
=_-ER?U_VKfL#D7@TX<7add^[f2/@e<]K;fO^(P=<Y#BP5]V\=.\A7#K#J(eR#P7
VYSU_R?ZO4WXc.cVEcEf+C#S995@;Y9(;6Wb3@&cT.WI.dLN]^\J;GSRAILWC368
W0#PV#WTXHT+[6Lg5>6)T6CM@<d.HeZf0QeE(R06OGE-QGCSL4P<fSZG,e-;):N_
dW0YX<;&9Ag.&3/PB;K7B)RRg5KY6UEH:(K4d3<bSV>gL>&?aLM@@\:JB&GK]]2K
?;G+T041@IR@,B_&5QYf73W6CXHLN_/DDZV)-gV>88ESP)^23YIQ<+/d#U///#gg
P[X/:(.gaS(:JPCC=KJDY(<AcYYc+RQ7A8WLXTg(MS20I^NAJ[EFI#Qb4Q^LVJaV
.T);GVKcFc\/N@C:G_SFWG=)d9Fe1:S7:aIMXX(YL5V4?f5J/HR^DG=7&VO2)^CU
5[EDM)cgDMN.e.)[4(IYJD?e,HaK50LNEF6AR,LM\7QVdFSRBVG@[7#[8aJfN4&:
LA3ffMF+6T172U6.@&C55ZNMeS#=b+F_9?eff)</.6DK^:<;W@UfP(9R6\#CQ-FB
7La:0]GX?AM,C#f^-?g>T.O)c9Pdb81(3?71WI+=dX9^=D+L5T?=UIZX/V1H.?BU
Q>0\Y<:)#=8,c+7>O&9,Q1T[E:HGQSa>SPcQ+fFZK4b#K.I^Z=20bUC-KIC-@Zd.
7)R\Pc&H[8-NECfFN5c^OZI=YOEf8U#(>D4-PMX0]Oe;U?1&DIRA^Cf?V,?SVN.T
58=@SAC01[+.HHKc?-RWCf.@CG_^:2dJe=b_@JO)e8;DAN;/Y[E[RASEI83GE09,
9cM6;F?ZIG@G][0N3e)+G1?P(JUV9BZfJc\?JeVKJ0^I0+6W++Qa]/NFKIU4,N@Q
K^MN7C5LHe2T@G+,^M)>/,_)=I]0?1,VbYGZS:KWC2-#(BMIOH2U2+.X.ZPd?6dJ
I6H7<,=KMN2C+MT#79FKGVH#R(I<eggH_NM]@L=g]LC7D(?Y>AD\RT24F9.=):-/
Xa&H=gLb/O#UFLXJFRGbO?E<_X9O@834Zb-=6+T:g5N.]/IcUFS[/JC;e3(D5<NB
B-QW1I<K2DTg\P,&Y>6VYL4:XS?dT3X^,S?ZPdH,Te.2,LFW5c)f<9V=@E[9a_(7
2D0VZIdDV3NJEL>c#?I0?HF;JVG,UGC->@#cbFUZU]F/-d,57+C:]TEO-86LdZ8f
b#-<F50?(b0)0V(R_04c5dQCE^-Z^RTV&2)FJ7XZ4_J\CMQ8,bGO?0UASgVT:DML
H&:H7_0<7-K-YZOA_\\[f4F6P39IIR=]A8A:\a+LFEJ=]JecTE)Rf(7,QNCD_MGf
3c.g3Z+\B7^3V[CXY<X@:UC@F7>L73<d+5d.GOdE10Z[M.YN^>6UBaO=]#C8PHHR
?F@9f;F3H=-\L8WA)FfJUCTF++a32e1C])Y\Pe.6\\ZPZW^ET7Baaf_01Xe-Z3#:
S2?HE94I6bS(1a[-YUA?2;9:U4)I1eY2\+#-4a]CADfWK+DU41YCT26fV21+a957
e8T#B[dae04V-R?]UR1;edU=b\:]aKR&H?JO95=D41HcZ/QfQ.34QaP?QA3/1de6
5=ILE^dd^ARaRW2N;XM_G,>X+R5##J@g#dSa5cG.P4LFe@MHcb^=JP->:YeGTQH#
.e[TBbg3^&K9c(9KfSRLO.^-GPR7>@.)]gTP+R#,QaVGMSdXb@R#e,K)\/WB=[B8
E;D0?N-29[..Kb+@bSF;EeWZ>RLPPX/]+7?6[^9aXCRb2Mb,B4FK?@LCM<_Q:WfJ
V81d.Wb5CR[MLDF&Q5,.dL;?32E7c8Ge&TBd+#gWBC4V:1:0O985^[CV]7BD92D^
];:B,_.X.b76&34]X)Nc,9d3G@X7E)ETC\/[@54/.4b>47EOCT7;JT4)8HX@]@PO
)(HK99[>=F4de3c3e>-Ae89X(7UX[e&V@G+81VGgI)?7OKD>3+.29DF\,\D@/Q/H
\&K:X:G+00?IE#CIHBc\eGF/+L;WPQeN-cQ1^_?_?XPB:5_DSUMHKDFY:=F[],1c
#3,,ESW\D].FHZ,g:HG8TCaLD^Y=22-1[5</@a<C\G?O4#=PO/2TG;&UGY>5A28#
BQ4E[@5Q+D(aV6T+)3:c]93d6\57^8J=<3J1+[0dU88MVeFWQBDc.G^R-56aS63+
bT:H;?HV=7bcd?>Y1G0L?T.(/H(T@,:=#6:C1<K:-]8gN4JQb@H#N^IVc;TT0g;c
[aL&/FB+\IN.CXIM2\fbT]1D7TZ\4+8^2XZ8OM6b3_\_UbIe#Q&IM^4T:-^XAI;D
DK_XdNbUHK(3?SDK78TIN/T9gL/b3Ka\=G1VKf2H:_8a+gdIB\B;-]>Z69e#bACF
8Dd.C-<b9#AMJ4(>&UGbD-?Qb16;2K1H+Z=T.BSU(WOJQEG-A_c@C+W?)Lc8:7)C
g)_GaRZV^6XYBdT,RT4?VF?B-]dZdZG#N_a=M.7]J-&P]YYYP[-,?4efJUY^U6H]
e-+/V--+Sc@MV+4W?7[^N^V5KSL8[(#811O:KKX>P=3?X9Y#+&X-G7^865:YDAG8
dBYV)C&3AE&,7+T[E134<1\NGJ;9(R3C_5#@IIdg/.CM3E/MMQO]gTgDd3g6cX;A
HNI)8=>JO;SXY/6L#EJ[aFBZN9UO.=&UdOW7S#P;_FS\NP#+/BgSF8T42/(/\@]T
2^R(Q;_S(5(T=cE?c#OB/.D+Y[TDYRE^/LT_+43gLS\9F.[SH;HfHI1E:16MOUaE
@?eH-+eI&A=(3.OEceV<]G25WaBU\&(JW/BD=c;=X18gJ2002AK_(GZ5UGaaU9))
YOaMQ,F<B]W<-)#N)8;ZQOOCT_2,_d9fRX]P&d^M]C60Z5dBQ@ZP=.cfVTL2?Yd=
WQe?)0SXOd4bH-JI6A)R^&(Z\Q8g(6]I?+#/DL<@OG2GS435]N>-U1#)(9^d^b@N
H428/ILJK5E]\FH]S0;T=./,C+<#f1LMFbIgDGD;WP0>8.4^:aEBQ^^A2@R[[9Q^
JG)&IeU)7ME.8F88Q/Jg)\dLcU]1^bB?TCc[_,Y9ZKYU:^D]P\@G@VLA+V9c^UeJ
(<<TQM;)WdBEd=K/=60^)\WY)ROYE5E[YCKQPN[[+:cNF=OU2_O4L05/H.P96(M8
([gKCec&X3:dcP:]e=Z6</PX]Za21Q?+9_\9)+S130ggBcbWT@\GQ.P,=V78X<Gd
QC\DZAVUGe:)?L.\8/C)K4,6]UW)\7H.98EM7@LX@JcU=,4ACOAcB2N-KH&=LFQf
WYP=XRf6e+=@NLH8O;ZD8a929,fgEa<b>,#WcSXT^1WK.)1CYM=-</Ke0K#d:NCb
&TM1#08KO^@=W(E)DI@2EUK23A-]<A,RRU>Q&7B7CB>&B>SaSK[4UB/,=H0,+RC#
;F&L=SLe>F#W+gU(DPeddL6P#\>fCBIVg8\&,^TbANPB,I8g3@>(AV(:.R304AGK
Qb;Tf2Ea>:&NJ7PL:7[I[H0OF(4>N2ZSGc1\[DB6>_0bYbBAM>\2OI3@V(4[M;-Z
SN6=f):C;&1V&S;eV^=6e>+\aG87c=>8=\Z(PCOf1.<aCRAbYSKKLCK.3Z34=;@C
0baMTKb/84If7#=DD(HN7)Q/NcZ\HgaaM2+ee\X<HWBT&.,QY.OCgH;ebB[/Q38_
Jb8^+0XE=18DU?4&\5d2)-(8NCN2^/RH/A.f(\RQb@GdGJ^RZ/=XEaB#V7H8]cA_
LJg]UO/UKOQ;HC<O);EZ/9EIX8;ISeC/Z6QWSQ:(S8-R]+:2_4R5A=7T5Ba0gG8L
.DOYW+K[0M;;@\EfQ74b_&23)@7IA<4dcWc6cVG#3cNfX,=C42H:MF1K5Gb>N:O(
2b462MI1^&=PC8H@R17#&F>-a]g>X#=T&8)-/2=D<]W>MSR?W\bGMN_feM6&P_@.
e=MN]ZX=6>Z)/Le=bC/_S17G+ZCTAg-N3?F\cUJ=HIfdY[g89.d6=2f3MWA7U<J4
II;3\:eIcW&U9G5;GJf;5:\DM=O<gRc_P)TF\WQ0:U6HZOcCS4]Bg>?GPT9F&6<\
88M[OZ/#ZFb:9GB5b#WI2KI[-CN^OW,6V4Sa6O=91KTQ_OE>A2\TTgQ=_3JW2V<H
WCW/f@5D)X8QFM07]M4ZWJQ^c#&\e96\N6eF:7UBc2<\;]]OEFaNASb9TM,;2.e;
d7.]HJFF^>O?#)[)W;gI2#+#EV:<2EaVV_dY8&^b94K^G[CRTbcf/]@L5K)>J6@U
TfVIFfe1LD.NKFS]WXXVQ])b&b(9SN7F,;C1RI=,E.86a(YcNAVF;#3>P&1fX]O.
OH),eCZTXJa1;bMRg)OQKU2gaRMRWY\+E8O5dAG8g2D/;7-aQ&EH199?\_V(7T@>
1H50W_F5a^L3EI(-NBW.,9I(bIgEKG.Yb)f:O?ccKE1ZM,7Va4,/+NWAcMDK7BGL
^(U?.3BPXH8TD31RB/OF-TPQX(#>:d1I[(Ie9+Z_[2:59@J^A;W=,(@TAXEJH&X)
.20Lg.77a80:BAb(K+<GH:8,?OB?QPR7K-R+8a4NETFEMP=/R@b63U9=C:B\JT#A
HE),Z-[/>[M@AVQ=QB)K,:CREHXaZ50\KJD?YPG,PZX&92L[Z:[K-H9:XX3DC/XA
H\+SL752=_ZAG1+R1_^9?\2D\9fZDK39@5]Z#8QK#H^6KAHZ^Y:7dgRbY3WQUAfM
B[\_M+WE0N/VO#+D(Hf=L1(/K_^VN\Q06A4b,3OVSD6DKc(Tce+SaK9#c8?ULG4-
M;QM]?Z5a8dSB=c8c+BZV)H/0+,cW\OVKD[8^\P=g)N(S,\L3WFDG(K2ggZQS>[G
Zc^629=LS2FLSAZTMX14Q,0^9PNMgZ4K;^L8GUGKeX>@1#RDL=(<Q_&?YVS7TY8^
24YH^QWZ^X>aQfO(^#c/c7>8?S4L:b\E<J?DcZRLP;C\EZ22UGUd.YC#Z^I)0agD
&f&5eYM&U/]]Y(A_(X_&#IVfa_8.e0GZfB/N+Na>Ua#E1W,7XaC)7]T->a?GM3M?
VOH];_+<D\E8<H;TW-7HMeQa,O6T&W>>H^Baf:#V-VY)R>34XL]T:6Y8?Y<a?HgS
T;,[B#B0MND7DD2I,YYOP^&G2R[B4D]EdU#C^MgS:03&M0_0AgS9da]9LRF)8<9Z
MI;a7-4=,X>VOONNd7Hb1VbGUG]>_7[)g8=123fMbDNc+d6TeT3F_PgI<ZH4AEPc
+4WedJ_V]65.^9+/DOXU:VUW):eRXXNHG_Gd/+:dY^8[-=@6<9@--ePRGCK4L.Q0
E\_533fcR)>GdN>Z2^(6Q@TeQ[#6#FG;/N0FB8V_LV,bGKW9AH[X)H?dP)WANQJT
a4d3/28Z;CM@6Lf]=NL+\cXMN3@TW+5>VTP,[S)R)E]OS^KT^e9]:]VcZOU>bJF=
.II;]aYK<:0]M<@eLR9:C7=4U_c\6(R1eB#M-Z#UMZ:,8&+OT_NR9RFJYVYbN:4=
g?d;OD4@Z/MZMCDY7dU7c^I(9]e)DgAY,dMM=@9^P_-Q:61K_&a1QD]7,2??0?8^
#/BM,-R47-5a5e6W4@Y4TJL\J67#Y40>DSBgTQA7,.MW^M^\f/[8U3^/dcP,O9eS
5[/B(g>#_>V@GU@cd#/[,-cP\FS&N=;f-YQXU@dX@VO+M8:.A0<[H8A9_M06>WXB
f[&b8.Q6Fgc-7UQ\@7D8ISaRILP6gc?7;W0gJ@,B\L:,C;]]]6@1WcS[Y+(Y7SLB
LQHQL#Ec3@()RPL9b4&J;R7/H5+FY3U?E?1P<<;eNS4;WX?.+JK5#/[@)\<#TM]1
2fX9@1;V]/E/SKEKI0M/5_;1BbXOQUZTH?E^N32WJFb(a>X<fIc/?]@Z_YMaF90-
0-If)T/5a?4[N0\DX^e9@;G(6WJU\^g>>9EWCQII]420(G]@K?=(I>,cO7U?6\AR
2QETHBU@..&=<@aNe)&,8Ebg?GL)M3J:)c+>,R#D<GCg4=,T,KeO[XNdbGb@(YXZ
W:#YCB\IY_J5?ZKd,V,S@U=98+FfHYFE#WMJd.C#Z@C3=(M:Q[QZe9C)JG^G1CLZ
NaIEAWW/aWVT+c9VP7+ECAE\&O06d,JO&G-7g_2(b((8S@_(V+01AMB9;CBI?1QU
C:(f<H8L8_4[JVg05_#&<NGX=P_)I9X4QM^<YPb1b2Z-N=d1E9E,((VSI:9WPg.F
_>77];0N]]CDS.g13Ha<C9=M[VT92DK-bW4JNJ5;VHd]1D@ZD6LO.Oga(-@:f#6E
e)KTf8Pb>7=6DS0GUZbEd2B,b\?BF^0JY/>1<<c3?,71W)6_:g_d2R4XPFATREdQ
=[AJ]^_LZ^]I;af]-Z39>aQKeGKF>6bKB6Y10N;++L<(FM(\5Z#cCUa\?@HBFc,8
O)ggg+bG_I=JJ;aP8;8b7E09YgeB\S_I3J(T56F9=KUVKg22\OSHD-&6,ZQ8_B&W
KKEabc[GU.NXf@9<2fZUILL;7]b-R\7PFTCM@M.YOg+UVRJa9N4[)YZ2MU=^e_VL
V\W6FS+,>gPfS83I=0WKIg]Z8]V4e80R?abXD=YORYT>Kb&TL?d]H-U+[HFXIV]Q
FQ318H27XFT]L0#/5]3R5D92Y)V(R#G]WB#Hg55CH+3Z^]4N?F-)1\_UP)H(F(DQ
FG1K3TG]PWFGece7M1T3,fPId;?c:=.UG-,KY;5HSI0?.2fWQZ^[\3^1.38@-BEb
<&\\Y,XH\;2b,cZP2f[-&.S(g[MfIf:Lc><W\[DFHTaL8,Q1\-KJ]9W3WE7L4QF7
-JX\=4^^.VWO,G_RW/Q<97c@-[F(_O&c.C)>-/+F\SQ8S2QLQ6EUZ[(SG]^b[aDQ
T(Y?agM]O1K-DHbZ.gWdB<[E>c-8_<=f:BF=+f@VYg5IB)/E_P;UeBCVF7W=@&@a
RI30T1]S,;<dZ-4<aXNB;W.IB,f]U=-M1T1TXI^:M).cEQ]H76bCc.HJM\MF=7(<
R.AWbR5B]C;[H=1PA8eBIVT:e1WdQMK6@ScMVH01PUC62S,-)=Y1B]2GKB:TNIRA
YbJS:+_NI^K\V27O@>.<&S_:ZdWX;,2Y+GR0<D36202Td@g.eX0Ee(R1,e5GJK?L
P@ANRPD3(PHa_2HfgX8(fW3&Ld<#Pe]&9cW<4>O:ZQ3[-8KSKJO5(3U(-R5VK02X
3?YQZAC4BFS51PW_FO/CKY;;[5>aTNC,5f7/T4:0S3K4N),\?;4Ta._;HDN@8a[(
6g.c\6VbV<)e3/<\^KIQYOH0O7,;GQX2SA(6I+S1.5>XHS,OO6R1/b>Y2MNGc+@J
C<B77_9+<[Q>ET+Y>c3XLYd4aO\<N=XB(<_G76E-C6E+24.S:0=a705<\)a]PJZ5
C<80)=G4\2K\R^&HdR/DO^&Wf\?#->6>+RX)-A(_^+KdfP3JS13&B/]YJc4.A[G[
@fV9D6+,gLC3,=@7LNE;#L=aUZbL=OA_4DM0cICd<8TJ1FA=\6,76@aX)GDS-Z3_
QO6UY8e\V<PX/^aI_E?QfN@aE\WD/H0dY?A-VBR&ZcIVJ?8ZLT7=,6YaJ)gMcNV4
J9XbdQdPHEK<,\4+(H@MV]@\;Me&IUL+J9Y@;4cP/DR)G]#c&#8O-99A;A3TP\Ud
\gPEH:d_UGG]]NRA5^a^b_F[/C#<&K84@WUJK[Y#>O8Z1O:JLMPV4SdTMT84Ge2L
.<3I)e^2H;\9-E-JSV)M1U/#.(MWCC?9\8gC14-g<PAPU?5^M(X1B)3&MVIW5Vf>
B9A<UCF86JIg5R4I@a+ZE=4?YMV[d6H?V[)LZ=BT16U5SdcOfRSfTN)8fA?Qgcc9
(2.d].EQC[>:eZ3dEU?=_[:aIcOc[QXVJWd/>OE[4cO(<HKJ.M-UP06(#IX^g(Qd
IF__P?XW#9D0_]^;U7e+.DG\:XI+T>(+1YWR\@UL2V3fMO(YXcQc>07KD:ZP[bVS
@fHccRK:=@.Kg/P=e[L^RFe)46E;Q#,5UZ39&M=:M-Jb(aBBN+D2BPXACA41,ILa
+G2N-[<H)/fQA4(/b>W(.YG,-R)3)#O;_^[BN4=PQP+g\[+<Red/dW(+R3\R>]KN
d^8L)WW[C9Wf5(?Re6ME]GH49VAD.(_@NfY/,Q])SRb@a#GWLVI3X[@gD0ZXBLd^
94URFC^:V&-?U..RXRS43:SL61DWdXI=^H(K4BAPWAe-]8;<:eO5T00?7K>HgG;+
=50@.F[<8\T^5NZ8Hb^Ad7=)04)R)#<[f\43c5@&Y2^,ScM/#[:4^.b]RTT>VYX7
2A#CA0L]fgdE17:0J)8\B)EXF42I)0Z9Ceb.@TW)LgI;.QJY](B=_K;OHT6.07TU
IYe,OM4bX1C)_[32QE9]D(FE>:+/5]BTAMeDD[Y:IG7J_+@5gZARB-]F#-RXXA2:
MUMD\^DO2.V/;V;8D>JXU?Z:Q.=,>::B9V-5A&M(W\83/5=);(MfCY9\3DQF)W7Q
M^52edXb(IJBHSeBYEB>&E#.46g&GZVDX/aV)R&4>Z1JI+^.eIfgI=KSPgYTdA_8
PBd#=a5YeS<__b[c^bYT-9K\>daK-0#dTfD^0eOYPUdJ-dgdEeZ5/CBC]3RUO@C8
e=0.QN_?E+.CU>f-7+dB-U^V@E<MbJK7.9:5@DN.dfU)?9d9U#I7e224T,PA(e&Q
K7:2gTEXc^H2c-(MeZa\K\#YGV23=^>:WYNSeSNc6RN7I]YLPP2KGW4_0MQ>aZYb
&HXbQT)PR-<OY+Q#W966J1X]/@.Hgg0[7C?THTTF25g)d1L-A+A^7S:LH#-Cb,d-
EZ&AT/0?T;G8&LJFJV.A(;46A8S+b8(4281AMDB&6FaIQFbE0^R6)(H1D<@A(V5I
<);OgZfVEZVYc?-^]gB1Va7R/V)afXa_+W=RNL^C:&1SH@P?3ZWX/Q&PeM(0C5A,
E+_D>)I\Z\V>HLXJ-[Td]b]Ha85DD1Ka+f8:QW)&G>g)H;:AcPgVPCaO<Z0J/@YE
0=I.W;(-&]8PY<_UZ=)X86W0&&L=B:+E_U6N-.=47-^g=))O=UJH_.3-ICWd-#N^
(1I\IeV=4c?Y72f0Q]F<^NHB=b\25;>,GP1\=XSg/?32.K?YS?P-)BH_G7MITcFB
3<,10e3<bZ36ZE7KO2@^W@_1<(+-D[8??A8.G+PS:6T9=;#:_#JU[S@NA&?5RHT,
-6d>59RZC3;AXdYQ?Fedc6NSMbT:L=EGY6cH1:Jd5bc2Yd?X@2^18(;\))VfB40O
G(B\GHCH1^>-gO1DGU?g,&/:2)9KUfC-Z&PEZ?4RbMMR:[J,_PSdDQ\A3KBQ:GDG
a[6S3>_cFQR])8f#CT\GN=:bKW+E;3RPf498VL]&f[-LAZBMDRCE5RX2OVO;<B^]
\:P@fC=d@\Q)WE-PcRHGM,;UFXX_C+PY+;3^)DXQ-0PJW0_bW+6BTdRB08?5TJ0a
(SPG.@R_5T7Q(BHLL5aJc[UE&?PJ]9LQ6VN:IMZ:&HTXP]CD:3U;C\O>L\)CI2?6
6;+4:DY+#IXB]YJ0eE3(0=d827MK\LAV7#KX)UIA[#5\)+-BW]L_Kf>:f2LaYU><
XU>3_DM=:_+4\3:J-]Sb82UD2Q;-,Q:^=7).RQZSS</T94[&gSRY@PKHR)@_)E9H
W1K&/8HU6d;+S=W;AN(>KK#RZM;:,@,B[Z-L[GH(2>c^-N7ON&aWC]f+M4U[&#=1
E(/R;bY(&J=9U12[Z&Y9=C@CIF<GUd_T8dc-Y1TPRM4X_910eTB5M_NeO[VWgW\O
R\]+_dF#Y6/EIC_XUgMS2c)ZN8U8\0TTTTeYTL)(IN+&g+P/82abDcNKaG=_SG82
C0ICWa\(GTEV3T0S7O&bg&RBGY=c,@KWM9/O:,\c8Z&5<W^+S910/5I/=fVF1g7C
ED?MR/T\J;@Mb-.f]#[Q7+/b(abVP).E1CcM?NHJ=(RJ@0VI6(0BbL;cSV7PW)2B
eV>TXWaD/gNJU;KG50d]I_5bXBR,d(P4eNN_&]]CWS9+VcOW&P4/6F19]FFM0HfW
fF1UOH9)5[BG\[I[aQMdN2P39I_N<7e[CYR7g)&GHK8.Le_93,[G6/I(LB/TIK0d
JKcEI39;?B\_5fBX.-LJ44JRVC2?BF,PN=WQMG6NX9Y99::R1U[L=:4[,EQ?e0Y\
K1=^P-b,CO26AE9/LOQ\b\#D740V,AU,PbU8WU\DH>3CSVI6MY4(1R:R3/D_ZFN7
[HC[WN-I/7/13fe@L+_-8]]KN2ID81ECdePD_,)[2M8WH=_2LR7H>VXaIH;+TW_K
^7d#)-7E(Y\^GN5;M7c7]K?E6e[0C4\3W7Z>GSc+)E+NBdRK63?::#6A=Q&.DJ85
a#IH2:(^.\cI(b07?,2@2O#&Y:++V>3,(3_6b8OQDDX2:YbXXd6Pb[NROTLa/^U+
6O>aCU]NA;GXMWJ#H?5L7WA+,(\UU@aX+#R1d)\\O-&_L&+\.\.=Q(?3).Z)>Wg<
(U0X6^eCSS=@cQE>S3A]4R2<[<^K@U.VHKPZ780\Lg4N+cL7@NV0J&)++2c4)a>R
73\I#D82QI+2<^YS_M^_;\B3\=:EL9gL,fQeME:Z]IK0MDOdKG5Y;:5Z&@:^.Q@R
gB7OR.0SWg?NKY[[Y.=#>A-CZDfE9DHO@ET4W2bfH2d70XZZV?HWCb&gO1O20f7<
g4+NOUIMR1)(UN<bMeL186XcX]JZJ)eJHaJ0WO_HCJCJf<J8BV96=9F7Vd26PIBf
;]C6S[d46I4(f--fCI&F#[8:9J0;F>+g#Q]83a>W&bdbd1Ude[7?>CN6a@-IO?JH
dB#7&DaI#<QI8\P5=F-O?03^W]AWc/aCQEO)L:<Fd4<(XAb\/2dL[<Z)V07@SDS_
(OZ@<VK=Wd#_2M>MFdG)YTH=7.Ha-gXL._RG3c@XN59=NL,eKI,)(1D&Jg[J__2d
;:A]JV@UPf3YQ5X4/g#,I&KJ5U@Sb^;J7O>V_T-0)C-LL/B93+gRVK@2C&g4ETea
BJgG\D^4f-Gg4Q1<6]BFdNeZ3KbD-YWX-.-(e(aQ8PW-<Z]D/cCALJ6#>K9@>@A\
&PK\?Ud3&X@YB(-IFE6C;AA4Rf=>SJ;dHeaa.DM-g.Dad/3)5_810cRK5dDN(c8.
1-6W\5F&O>eWW\NcT#Z/D6>1M:G=]4:]fOC03e;7aY?e8/eR,JLO5T9VH:_RYE;T
ZfU03QN3Z+&0H1fU<aO>;TKFG24e^10Z,b-HR4CNZ5_LAI0@T3H;;dI&b,+:Rg^I
<)9.MZ.N1BTX.Z?WEF5U9R3G7280DQI<[UAb>][YC8UY5A8ebCR]>POB+ePUf/S8
c;)bAH4c_),.#N4[HG<AF]_.7[5fVJ=RU^DXZGVI>T=BcW?T@fK5,--892-ZTZT[
8Z3=^Z[20YQ(K;T4]8E_DeFJF7>026CCe8BYT:&?P3692KX,2E/5Q>?24?R&G.e:
6OH&Q>==I[?/2Zg<@>@L-f7dU;?Ra-D-0/L.b=3IIM(H/eB9\?\@K</F.EaO2T>R
:PRd>&_/-9U9f:[R.;6=7OQGGQ:;U2c:^:U]L:TNb@\&N::U,>LUY7HZAe&&TN67
Ic-@[)B,_>,b6:TXJgPPQNB6B@Ya(J@?VXD27/2G])#+8ZJGO1)#bg&T7eH8R_5X
Q]-7RLdB/34JJOA2bZ04c,MeU[B-/9QRE+f=<Z/-Z@\[AT=N?bXa52M_?35SAX7&
7VO6A02BSW1G#7(:HE>TcET#:;Qf,d];Mb-N9Ofd&JS5;3:LZG0U96WK1PgbWG3]
-2:464U#f]A/Ff[3-G(abR6M?a:[GY@>I;HW27eJ9fge+f&OKcV2)Obb._PF;-M7
0bd<V?_?=a;eEJgd3e<TL&4T=A^Z346:g\C54_?97&G4QYYO53>QHZXCMW6UM3Pf
H3<&G4F_Q.Ecd>;Ie+^]V5cM>FcQ?AM0S=49_YW29Ye8:436?F4LSa^3D96)U7#\
?;Z;eSA5XZ3db(]^Z/#-9D6VgN)5^9fb1[@XH-G#Y;)dW?e40B&<>?Zb>D4BXW)X
)[Z^=e;aYLCaK7_YZE;;bfXJ.&,MHdO_ECZ+0-C@C;M+6_A@YJB;6(D9\<aD4SB.
B?2+<LDU2?,E0AFY5ec^5-1N:9WGa)FO\ODQ(;J>Y68TC7:2QA-#O2Nc7<0OU.LD
-K/H8YfNMAA//GcGUP<7G4[YV9QF/X#6\8\N/RZ0HT#TQ77?HXI1]aKZ(U(/+_5#
]UN<CG8)\1L6DeDb&.W1@[PR)UD,LaL-C0QGUc]X7X20bAMQ_</76dNRV,]/Z87M
1g(VV?)HYTEH0SC;fQD>R=0HG9RSSeRP;&FB6JY[e;3WX99L8D_S^QZ?KE@0F,dX
9b10UOdG#)_4W[[9];+@,Z=Q@4?X88LY9=AL,QM@EV/T>BUE1-&HA+/7B_9M&YdH
bS>#1Ka;Y1I--B<NC1Z3<^>gX@3J.<g#0A7RPEa-Q0EFW/W[]Y^1E&7>KdN#X#21
IdCE#C]R9-NBE&\PC,+&X5#dXEW#b[M+IF^(.JHV8YC5H3L=05OTc<bFZ4+XKbgA
<9Y=_C+WE\QOX2]RWV@M?V-1LP++ZQSO9aVA?b<gM>5QNDB1D_W[>^J8f-\^9eA.
M1f:?F2LMW05:A(BUTG_g)=>6OUO;]O1H8NGaC1#Q>I?R6b3T^RL,QG2\.2??&Z?
^Ia]HP8Q4MA.51+^<Y5bTJMeG&H;6S,81f/&89FYK&5Rd)TYQ27M7FU5D-0]8&,D
CL)(,ZD6:ZcJVgMd,g:JH#TIeYM_[2Z(XE0BY]0BOCZXUS(3JdgeL5PVD>g6X3&f
K+gO\LMX:&(U2T7#g>+If1]NWA\L=g0b/QHAFO4]\dC7T;Y6@F;\:fH5]9PPIS^J
>4-W_V5aeMbRWGLL:K(a]dKe^U4dA9;3&)c&Q.Q[QA@]^2ZE9AS<TS.-?TE.)b=E
Q7;c+OBEJ\)V8(4H+GEKcB-e:RTPabgaLBTRZ]KP#G-Z2d@CR.GOCN>>HQ#LWTY(
ReX\Y9P>e8YG7UNY<2M58<W.[#g^0OUU7Kf,;J<KgQ>fF#Kc/f?\#AQfeaS].ZOW
)L7.1\9A+KKARCVR]3#W5-V9gR-XAJ<3BF3II&LKa_QLD6F.4@f>3F+25J2a+-)Q
H,;NW1?R:;eX7cLTN9aYT:N41QG[3bAJRX+ZF.Ue=&=\[BIa\9AgO6BF4#RB=[b8
7ccd:PdcM@^FGf_XE#4@bE(D6JPbaL@Te=/F\I\C-?+7FC(#DQBO?R&(>FeS4I@+
S+:N_?4E]81)c#]fc9c\?)(V.Ta-[TX0YeGGACIaGTE:7RC.2QE9]?aE>6,YU3\]
8>]f18C5)]6N1IbGKU:VE>AT<^=I]7#<3X:+;-TJADJ+R\,3<<:KgK(^17a#MI][
<87aL4(:.<7g[1[UY7e4E01eaG^V<Y3=6[\1T0@>d7HOKgX_Z@bDDNYHUTZH(P\c
8ZM=/?eW)>2&/XF>H5^M_P(&fJb0N1K47C,H)_&R_\f+P5:S0.cB)V>N^@KaXN=G
MDeYU-HGH..4YDFbSKIaCgTd.XHb;<HagD)d>.,18b)bZH90c]A6^XYNOCOYFQOU
a@4PAJ926I0@LWIOPTK>T=WHbFZc.U7a0.J[UQ3(RC]<,_T^4+5aNN)(JdJ>(\L(
J0Q<?K/\-,;X.b-3bQ[]-_[Q<RfO(WZ-9630[V&73Q.SOC<_L@28-4K.:;a99KC\
N<&2e_]0B6f7&3UEJa;T5TVBSf2)Yc&7F_b/@6.N^._D?5G7SPA)T]cf[B;8UQQ:
R.YT:Wc@@3PR@8>:93GZDAR29DSH3O\UR9\b;ZBccc/EP/FUJc4<?[GNe,@4.bHb
,.U1V&[E[g(L2b:E9\Ia.(F?1+3F#E?\NB;T4O(\B9ZRS763UcH8;a91.LVR-<d3
[[@g3MA]/G9A)-^<<K/PF[6D1=U(#8b#N8?SY5NW#:,Tf1EL4^&[E0BIP=RDZ.7#
V-1=^acbA\_#;G>E570BCLIMX(F?K^U+F1E9<QD.:RH43G9(G8V7V_LTA-0PZY;6
C#C6]OMKQ2O4->S<;;S8]T]T4;+S<:g0#,/(S3:MNbWN-;FN^d_4M?^_8/f@8C=8
;NB;5H77M\1YHOSbD:&3](dVaUGGRXDeB>=;]e\?6B/FV/.024(J0=]1J><__#>J
(56bL@GcW#&<MR2T#TA]^J[YMfNdf^[X.XgIN7NADEcA^0Y7<DI\.DMa5EWF\d9S
JgVE9-Da7I([c_fPQ80Cc9&MO]3A/#[Z5S@C1UEaG1&18@HdV?BOP.bXMDD-OWb1
cV5g5=O,abg?.7f]&9_8L#-Uf]H&f.gLb0,36084YTLacI#(cS&([@BKUd8JO[^V
O>?P>?HMWeGE;Sb:W[IHM^G_-&<<-:Ug[]:+04/ZZ)E2MB]9-C91f695^V]2Z?U,
M=[PEX8+K4&?^,YGXV3>H.U08;?F^,?0Se<HA#1MJAA;HZ4T=^g9V4RX>HHg2Jd8
=;/WOb5_Z54\XRge8[,57Z-D@(WU&,9#Id,9Q2?[gKCg/Zg?6]4XJ1?N^Yd2_eJd
a-A:G/f0-227O-UDR@;fN(EPFF#d&?9L-,^:?-be>B)CM/6UBRFTCMeI&@[HU:_K
)J.AE:1VcT>QW^=6?SX1>gQd=WZ>[N6JZbRBCH=U(F[7[6>T/CQ;=PaGW(QSFP@7
TWBC>2J1NP-=7ZBN?6Hg4X&;8,(&]4>,X\?Vd,Z).b[@aL.AF:\NVL[1Je)4D[cM
WcZL+&/#,K,;X[:8>^4bXUb)S)(AQdd0gJYaZ5\2gN/R&G>c4MV@QN#c1Kd=,)F^
Z^6T?>f@MJ@MSd]U4F?.ES1-X/QUe48RO]e<908O<Z.&cZ4.3I6>#RR((gN]gO1&
ZJF,#WHP)K2:@8<f)KF_E?B_=5+M^B[6+^M?/-beG?YHAJ[EITE.86G4,HdH:GK,
IP]/&90e^\#e,gL,AgVW4f/+K[2RL/16.L&Y/G5KHL9->#9=->7-JH&A&c(.8TD:
>J5I;KcW>dLN4g(1XR_KTL+W\aJ\EgM+3K=@][T-=(+W.B^Y\gZ=&U4](P=GL:=;
dcHT,fHd/Y5JF/Z08VSQ-V@-d6]DO42a<Tb?5Ob=[4G.g=a2TfMFcPEWdDSO/M?X
9e1GV_Y,SO7LL9?<PfYgM368C.)0_3=?4Bb<b3CL608-AO)^+)]c(cZ(M=(d+aR\
0ZC<6ERG[FNX].Z?Q]f2@3P/BLJ-#5<I5#L5#>N09;9US;NN]96#,QSE_,Ma5VcA
fdVXB&<KH(FFgRFC]R^b&7AR5I:dB9=B0ScISDI#PW(2H[O;Z55@.B)4bO&@-_gZ
QIWFND+ZDRS.ECQU)<>0<@+-G/41:FB0Dg.TN8;C9c^^],U^#]Z4<6LKW970/YfM
DCdcR_c)I5?VPb6a2+<7H7a\K+>3=#ET@ENLE\L_,AQ/eI1d13Oa1ETGfII3:2?=
R\Zb&-=R<H7X&#E1dLB@dd+@Pe507KN[#Gc0C18L;RJMcc-LU;I\aO^>a+VfGG,?
0I0\9ZGJ(SKD#XNWFTD.U-LW((#>]=.Ff7eCbFR]>Gfb0AI=WYM88d1fdH>^E+g=
Q+PVF;/60cKJ3JPWIJT[OYGJf,C:2WHOBW\8?HeFGAT-ObSZ;CZ<1Ma&_#9]=?)M
ERW9U?HKI233U8&[AQ<TYW&N.F\][4Z5=?Ge+ROSd@DN?HV,M:[eT9IVZf)_#;DU
Na)5a8a?f4(;+K,M>8+@PKH&20JGN[bDP,:XGWJUFF/A;CA0TN1#/]CRX#7-(]DD
GVd:P4MU&TS8CdXfYc@a3Df(ZKge(0XNSJR9F/P7b<Tgg^Dd-1f]?[[-(;Cf(9UV
S)EQ)<D\8:G:fO^LCOIS)6Rc_QI+7VQHCW0QE/=37JGG<#acd,HW;/S+Z#HQ^06^
?1e_O;g1;@&+MbUT3d,g^bF6.CYU2&+;f9FXU/8Yf9V_bQ?b-P1Q^bHd8bf05-ZO
AMdGFT\\EGNB7EZN@]75>48ZG^[?)8L\G]cX+.8KX@CE606R9:E1R^.99f4bVe)\
S5A0[,N)]WZ2&^I5]TMBCYT62T[\T-;FMZ29[_VZ?6(c&SC1D9:&3LH@3?NI/2XM
WGa9MS9<KgfQ_.=A99B6N^&BX(@)eZRZ3Lb&^^(GbR^8C)^87ZZGc4Ff)7RJ0V+:
\&E1&CM.:C(.H3S(8&FGK1G_J?C0]7=QH\SZ<0=)PQ5W@bW:Q=gB5?g-B+:4+af)
6-[OE8S]8YOg3-2MB++,V3d7P;#BY)^AbCJ(DFKE:(3=X<KZ;/YYK<#L)1J5QC(D
34+]=e.(UP6E^gB]OfVI<P40eg(9KRd<&S=SN?B?^D6,bBMNa&-;40bMc@@QQK=.
;[5RI7[^B_UT,WN]QF)+b6L)0>]/M2>)E-[/aa^IZ>E1L;BLdg=,(B@CD0?V?^TZ
C^@a-dKOEG)1JadQMY2_BM)I5SG)<8KER>ZZ0Z+7/D/;;_/fLf&LP_OTZC?f<f#;
O[1bO/J1e1]TD#V?;.A+XW8+.?@0d1/XX-?a-Cd>5KA:eUUH+]\Rdg(R\T4U&UTZ
3L:<7PR,gM>&V(0NFUO5;XFM&YcXG^B>L6:SDLOUNE3>5/514H4gQELM2)a4V6O&
P>8.7VcLa@2V=:MQ<8#becSHRX)eFgV0X^->P-2[?KPV<Y5Y86E3^WV(2@O.d_:]
(P+\IRI=EF<G#eE\B]0QVOV&.fM>;;_<8Y3PJY[BOFOFV3NRaX4-K]=4N/(H05Y+
P@&^G293-[\[Sf#M8]2F4,g_TNRa;[UV-,G\)\cZ6,&^?0FZ\PMPbG+ST3^AD\4f
BRTL_JfMN^I6FC=ZNJN03?d8C<G-1QJfO=V+CH](5GIF2\V0;]0?YgdF#_Cc;20D
S77@Pfc>R4PD:,BYegN#170K<@WIGUF?+,6Db3c+fd\f\#WbIa\e3W7S@4WIaMP>
C.dL7UO@2T4:d,<QM=Og3BK5<D,RG;gbD<)DT6WND3g1QcS]6Ha96W=bTW[#d5XY
9+fXL,-D9;KVZg-IdFg^QQ=@H;3ZI_RQMe2RZTf[6[WW6[&LRc<)8^?c+=9aTKPV
(e)QDS1<#cCI[(:N-?<157S@BB95)g57XLW6/_aPQR=1d-A;M]8X#D@_T-OR&NT+
/ec7(^9,Q+/-06Za^_fNU(NfEc6T1U0HV3W8;[@c/eR7<ZLA-40@A>J2;P8F\O5E
GJ64F;PS&e0SY;PELeGM1+U-ELfS-NLUF7EbDJNJ&bZdW<L<\]</.\T\IP7[_#U;
EbGZQAO&HKYY-=SJ=d8^W40dRJD5cSSI?1=I5SJIFF,XAK=+3JHD,UX2JM,7TI:,
9gDRDW?)CgQ4Y^YZ-#A,#(C.c81/>4.fc,?_@G]48=)O,2GdD126B,74#+F4]B;-
37#?Q31?SbC=(]>E):UeC_&_W>EEIJbV_=QTUD_A_M^6B&N^4E265fB,S&ZS#,):
f6E[^9c^SO]Hg+N1?&QVKV^4SL/5J+MECVVHU55fK0XIRUIIAaI-IT5IOCL74+7-
_,8HP6EeO08a?FM2W?9W.E[YW;<:_,O=&]a\.(6\)6IX;L(>9T1,7.^F(6MP.+<,
]b987ZO\KD2=3H3RW]D?A=g=/_86Z/Q8@7]P:JLDN2<5<C]HIf1dRQ#02LQ;[@-0
e^(K=,c+TF99&_NW@_(?<,\WWRYQ\W<e1P8d[AA[FD72H,?HHeK\D2P=6])(OOIg
[K+VOFbC#d0YJ>0YWB3W<6L<A>1N)Q;K9=]Y6MWDD[=&L+1L7(HW;#HOOIbAEA@T
L.5@5LNR3](OK)1:Z@?Z8?),0fCI_KQQ@=)9CFQY<f4M]GB8X91JCZ]a#/M^D?BN
LX.BGZ\I=e5]V^Jf936Ge;-T=L>2^;PQ^1W7:8U.ND,5T[G,2/G[#\d.K/64Y>cZ
ZbUg4R,KO784]Af6^^R4,2@)9H\E:7afU_J6(5RE<:eZJ\25Q][AO#[2O_e]/X@)
:SE]IA?8R\Bd@W);fO_\Ac(TIF]c8\FA9IBRCQB@gXcd<^eGUL/d(#?dSRO8J=eZ
,gR0bA=8>NAP:IO?K[a(&dHB>?#@+?B80A\<8K]#fM/4e5gA633Q[_3HJJ1^\X[U
;U/V/&(C=#+G-O-,</@^[R#.V\g9L]XA4+JK+]G_)<M)CaYY-HR&+R_Y(D^FZM\7
5NXTdG<1bUKeb;;ZT@HSbJ.I6.8K#-JM__3@H@LW8c2,Q[X41(Zb__^g]9Q2:A?5
^+P7f;>_]]dY^X\d#MccZPUDND&VA@bN6=fQJ/IaCD_2,14,c7]Z_FbBW_XUbZ-F
gV=A]5#2.2bUd3MMYIDc:#8M^e>Q=)K7/6H>HUQA>6.1H4C+9&==8\8?AWSUXgJF
:^:-,f.NB<8M+BAQ_O]<JGMTFV:\9?RM\;8I043&gY<fVLXGV\:/cB;>&9W4Hg:d
O=R#.OF?5NdT.a<I;/c1XG/gR^8F;WRQCfX;8g<3(8()M\,N0VVM,X]5M[bNO?7\
gd9GaIg5Nf<W>X+,XJ6?09Lab2O]SJB&^&G?UAZ-5TaS)O+5A=G?e;S^A7DY-UHR
X;_38@Q0UANL_NBQ.1LTAb?I#7Hc7\EcZ6MUf9cI4\LZZYB80)S897LW>Z0=WD@R
K7P=R3A9G,#b7B\:dB5F@@cb66L1eUE291.GX)HZJ/64)6_R:[>3;BGg@@b1LJ.=
J9fV(\cMBMaZVCP0IPW#&&1YO>PUJDKR,QPYbc&YR2]Z/L<^T:CR9L[QI;D+,6.@
IZ(?4#X_&JTccB>B;\#J0J),809b>KaRc.4]gY4AO0:aC]^H7LJZ6B#=<#93>ZZ<
cASOX?B3M<dH\;GMWYbE,I4#ZT9:3G-N+7f&,T3)MfJ-P)fK/c?><gI1>g=bK#TY
N4C56VFa3[Y.S+.LF)c2J2bBXJ]1/URBJ5>--\/7U>ICFAbIYLH0Z2;[-aW1a_9Y
?+UG,<#&1\(&C+.67[FUUONEd[[^#4UUb@0D4H7dCD=cH8g@b]>W:;^H=(^B^M//
DAS(+@04#NCf3.SQeOGPZ+:(J5b..1^G;bA/[@^UQ&cYT-c+.]8/gX75X?Bd5IHN
D(6;fHSY03+(-/NRPU7KeYRYcEbVW+,0<b5&B0@dZUEf4SS,f\F.GdcCN<6I?LTb
0LQB]=_be?;32IfV>6dOW(0d8Ac>9^.g.(@Z.T@Tc<HfWgP.E])57I.Ca@>[3H>>
9<R8cgb?>d,bR\_,HQNBJ#IdM;?+cgbUG4&68<[+=R[f3F_g/U_;1J4/^4]_\SH2
3^_W63DVRWCAc4AB,[KPEfSa,R+^=^5B&CPO+W:FDY,#TBOZ0G3+6-(J(9O89.6,
381/#9PD6Tg?D]b,[I;MKVFPI^E^O02W>NUd9c(P,-[_eHg6=GJFB0A__&,M?:J=
<Wg,f3JHMD._]e[GBC>>NN?5A:EB5B\=c\_(R8?&d4eP=a8\,M^1#dX8H](_,L3\
+LB#Xd2?K)MIB-)9MHC]..I2.:RB692LODM>+I3.4RdJ?W[+W?d8_OA+K@P+8)<K
)b@&],1V#Q[@?Y4A2Bc\JbD>N<O&Z#9O2QGQP;?eDCW?gY+CRAaQKAY:QFGJgHRZ
;:C9Nd[Z@9C=00K6IcPggA;-I&&=TPK/Z+/?LD>9fGUe;)fK8P;HO_1Mge_-O@W6
JLNLD^+(Mb4dLcD=9;<b5(_.NEC:+8R@B?Pd)^DSQbDAK3NO:<Z6)0aAM1edaVYG
TE/>HD=-KWLRc#95S-LM,&2+ZWNS8+P.^c]L@&Hg@.0F+U3^OPGg]Xd-K&^7CUY>
d;)MEA?0^G[],W2KHY>a0C:1>b0.L6=9D?W(_#H]O]).5&F^9g,H@@XJ?3;09G,[
7;D(V=D0.;FREGZ0^HRY9Ff4?&+U>QTCJ3Z:MYD@fTf1c4<#Q-;ae9^6L5(&-MD>
17YBQf.^BGZ1+9F5fZ->.[M2P>Aa^@a]80];8);#(B&;[018FBQI,UOP4<@:Q83Y
_7GOH(<]2<8#NT-F9DQ21Xb)YIFB9+aMC/E<IS;Y#Z(Q=>;d6&VA#a+?TY3cJ7M<
B?5XNX-TN6V8.QBU2^\#)Q&;TU7?\&83[IV?+Y^,\^.4<(dTI96/DX@IE?5WIa\5
E7)[8\gK+HXW?F3JN(LNgdRP+_QH&37&L@4AgKMF.KLBI=bU4KR&AJ/YdIcEHRZf
NAJIP/D6/0MR4THZAO04EA)XC5UPgG^E3^GJ)LG.K#=eNd:&I)7K/5D-E.&f@XV(
:L[+]00WHZ,6]:=e3dcfTgfMfE\-C203Y-#T>U[^d1D66M80^cY3JM&IDBLAMQ(g
RK&=+f7N6K@c3d-_/U)I&/4NX],73EAN86ESHbNe)4AL3K.[_cZ]KZS__./+fAJ/
1;[Nc<.UZS^(J.Q,=cNLSaIRWa3UH<P^^ba-a:8a#_8676.\aQ7R#1gcSS/6a(QC
K[20NeS,G2+gW;=_FI:;#d.0eIYdVgaWW-C</4\gK)g;+=XBY_0U(=:fO3P?88K7
^ZLJ66\b.^AAMcWUCAFT=bRa;_#,,?PWMEb)SV-3P)&1L0e5JZ>K18WVFfMe8HG;
f.O36OG8OH>Q628eWcNH3#<3W&cQ7TBa<+?3D]4fX(N<?(ML@C(;VDJ<=9M9T\:B
f^)eUg;Ke\BD,gKb<c7AF?C/b@]KI.Z6/0Fff\].2@B)_8\U.;-Y/5TEP=Ybb-,<
f-JI0SE6.TdJ\bV);d?Q[HMA_b:ba\3.WT[5OQK,DEWgDaC2SgD\?]3/Z&3.P8\=
T)=&R[a2.OD=KM&]&ced-2IZI0EcOfc+R[PPa9NSLg-OVgCUJePJWC9#>Q(ELF<0
-O3A?^Y@+Z]0#L(;dTE4LQ;N<YFBO9_+c@2[A,-Q^:H:YH4.@ZS5?\\\8-Vd::6Z
:?8BNH^CU=SE#PILbcVF2KJ88JaYSe0Y#,QG0GW/?KQ=X;?8ObGS;JTS&0KP,#OQ
J]:M;DNgFZQV]7g54cX<:4@H\GZD^S3C4XN4O>0CC;LbHKKXc@.>:^_?2Kc0KSJc
-RC94,;0>f[b3_B09O:Y#P@,4L5>IN?,J,e>&_U4^O-FWQ9)J^&<7N98957\1/BU
Vd(F^C>_J,\BPJ[CQeOe@JMG99#3eU+Gab<KZ8;eGN=g[QP,;.^abKM_,9R?L)W(
PF\-cAN?WL/#8.^LTT7;/6>g>&OVO>3W9?8IRJ.>M7g5Ed8LPSdabKGJRNL:a:]9
c0(T(@fW:^DV,&5S^FQHOc65-?bO?EQPWbF7I)7XAd>dC4#PWL[>e0?A&=^+d.^S
C\2;,:I;\JgJ/KX;UJZ>M2EI0UP?2U]2H52aG368@0.X-ER9J/F_V,A6>Ua3P[HN
3^cE6#?>.)OY^S#RHN__,,KKXU_4fKQ9;L?g0SX@G>J:@[2ZFO/[5CQ6,8DNUA^d
1MUF4TR9.MI+;)PV(QOgK5XF^F6N0YI5=SQS5=12-1c^1@G9UgP;SS1_1X[O6WSH
=XdZ8.#0QU/XGZZ3JD_,INOZM\]SI2UbDR;RZI,f1#E8ZP5^DK[N)g]-MD0&&fYL
>g=Ldg:^G=Ne6XXG2^R:I;/6+]T-B[02_LTG,0N<^8HK^g)g67F.QS,;RA-&&X_G
N#5ZC3E^df)8YRD&[;N(>G3LZ,CQ8c^P3S/)P0>fSc:<9MTcf3C@QC1.4\3bK#=B
DXD,]eX?b#NSI2GeS(4Gg2(@Z(A)>7<MG8fS_aT=/@P(PNE5GJM9@-@(e@,9W/1?
+<=DPSS1ONAR\1,@=UeUQLPMM4V?/W/Z_3fK0-.Y&.^_5W8HZJ#GG4>>P#aeE(83
(3B]0g8MZ6@+]=10Ba@K?([\?7KJ.14bVY18W&3UFGIY+8.5:DS6^IZ&EAQ/O9Hg
]I+bDQ(K#-QQO^+?FW3)]JAH++UZQf@QE:QX?JS)QD<QJ6^H&dL.J?8d55#2##K2
8eWP4Qc+Z,bf=S4CS]Ye+>,8HF0-M#;Ca2B:=FUe@1K[,-G915HP<&9@1&)_GaD9
0)526&-X[efVXDeJ+#5Le2Q<^V9::e>UYZD1c[<6M+0N)+,KD429IT^8>GWJ[WPN
bY^A.dg=FaD95/B9YMfV-[H;+]C&^6(,gZ69)NM1>N.H/3RR8Q..G)]VDHbAXL/U
R,fEWfPEIgA<-/?cAaP)WNE0/:&Re(?=gKF<2WFFN[F.]L^W,c9K8^CLH41JBTYb
C\AM>aW<#2A0P-RFK=@FS7e:Y&?QC+9g;fH8,FeaTEYeG=<?f9;e8a_0b):S]]EZ
6897TbS58g^F0.a+,SJF9Y?#D__4gf3Q?d(:DE5\?61:gFG-<\VbQb5\@+L6E@ZH
BPBEeZfGdT5EU\BGUJ3\Q)L)(TeeB4R]D<GH1W^575Y.X73a=^.d=QRD1C6OP8IJ
)g-PM#Z?Y70(ON1F\DcR_fA;(Ig//-.VYOX7CeCMD&U)X#^/+R.?KgZGH[-:TFfa
RZ0K6SZIPVW]fQHDJG#E\=f.&ZgDCY.-_D>:O^<V21^;fWL+-Z&3J8^[RCI\RRgW
f@eJPaGDPG/BH,QC3[#f.,S7]@V3V2TD,2&ZFM[b9.f.S68XM)IO);)>736;LIE8
d]<CB<@WGQ&S>L&=DBNeR7#gS+C6<IN/D<Ef77gB0O;7;?&@@S_3T)M.4[VQD>F5
TKVcU3:]G(WJU=QI8a0YK]C9GSUd)0?CbD_7XL/Q^)fHdG-CYbVZXAH+FDf^G\5f
</]ROcfD)]F4g:?8(0aaK)^ZQSce4^VNJ?8Mb+.<d;OJ8C>^7\GK66V[#\O;Q;OH
SVSP2+,XUe3B<]fcVW5ZLAS7N^D8I<;7@P=(;S1d;SH50,[7f8^I2Hg+?b(RQ@Z\
&C=71,g8IQIUOAeK_7Y3/+dc8?Y80VC?0BdBQ3L0dB.I[[D_[,dFe[g5]\==f=-.
EYHgXc/#5,Y-H.gg3Q:HfdIXD&LPWBOgF7)@S>F\UEc]408-NH@aZQ\PWXBT>74=
YO,EeYY:M&1g]G7bHPJYReFJNLKD3&BS#1#+2YPNK;U<f5I?#,5XT<->1W1U#C^R
GCf?8I\9.Q8#;]K3CT)3QY5S1)S-c=(I13b5C4fDX,=&6.N:MK#-_(Ab^7?-VQFX
-AK2c3>_#-g]RS_?T;\P9VQ:dLTJTV^b=T.Z=J=.@bH);H]#Z5-/MYURM[C(ITfP
_DI2CN-_+EQ=,EdRHS.G4?d-Vd9U496U.AC^RXGM;7;9IZ,,-07Z9G(DQ.cYO<Q]
V6HTISG5>HYX>BKD=1[A/C&;&PL.^ZBbL[]\6FFfg1(Wa.A,CfX/7KD>2E0IEbL]
ROQ.ceEJe35aB_eS)_T6:_#A-:Z:N&4;060ff>5I1411K?R\gSGIM]BaY-eCNA4G
(b0I<E01\LHF,\SF+BcHNc-[++>U?f;f>H[2Qf6Y_DE2cSEDP6C1W68H;@>fG2S3
cW7E4JT6)<H@[@#6LT+BfRfB+bIFcXUbd(,^N?YfJ>V>CE/06=UY<E>D(a[=&_W9
_WV9W\39I^STRSKaV(6YF@SJKGGQ5J+KI<Y)WaQ8?+)2@V,5e477Qf^:5]@/F<+_
/CLNA]=@YN-WVPHPE&d[dUfP#GI>Ja]J6&XP4-BAA>N8bS^GNPfWU#B44)\e5dc(
]@fX)3Z3O-QH>G4g@A1]8H^W&/>R_JaY\8-N5Z3A4AA7?;L5)7dVBf&X:eIdJ85F
0#03\e.JG?2DeU;cJ&>S(IeEabb5K4E82-4Z,/_=_Y]0QIE6U_<6T^=c;1^X]PHW
=-6URVc9ZMTS:@B:EU9KI\;/YJ9[9EAHb_IY3]cBXX.#2ZF?KN4VYRBQ:.^JF1g4
FLb6Z&M[;OG;HECYO0Cc#.,f;gVZ1[;aHdMQW]Y&cY+FMOF,eYIHF@UFHU:4CSfR
c]G:\ZZ_I>#R,1?aDN^;G4U#_,U^AZ?&^.\GU3[=.>2KRJ7Y0U\5-J:+2gU:4E5K
HIM+.3J6^3>C[7BZ+?,UTG,XB;(^73JQ:FCE0<cW7VD;^?;EDa8Q,H:Jg&1@.JgP
0ed_E\9ZR=bUK^/#@SQd.cDG/4?Q+6\2X<2OPI^:PdcN,_a:Q/3_FO=2-)(WcZ^I
<a(9U/g;61#>d7;G@5@M-[bHa7A3Z-2G]_9\5\H9e),?^<gX3@13J.7<G_f^a[]I
1/.4gQF]@G2TTD&S>@)1V/9=I:aYObb6/&F85/C;Z.6MCQC+Ye(L+Q:\;@T-/</R
c3(D7dJGT(:O6K,J&[51A54^>a&SPPJIa/Af(cN0)FJOMd>A73_/D1e0NMHB?>CK
dN\7.EWVYRJJV9G32_SM)1aM)<[JQ.-eE_GJ\g)Y170S.Z5CR;,QEOUPW;dReA&/
#]dJfaS[LQ/#bJ--LQI>&5M@\I&g#7.29bMDBU,R+D[L35-A\Y>FB877?Kcf#E8=
MDWB-:_BN9QHW<d+:JHQ?d>7#9=dX2N]PW0U22f^M.N4:GU0L^6QPM)4^.Daag1+
#bX<eVEFU.:?5Z<6(#cBNZE]Jbc\>YPS^VP#I]U2X8]_+H;/SB?_7aX6e38X2L3[
?ELf8M.GbR+N7]9f&.==[ZKaFa\@<9^0N3)^>b;RJf.FKF)aNcT7/SOIHC<CgV(b
_JfY]I7BQ3(&0aVRO)]Y-d9e@(+HZ=N2ZA;=N(=9.<VXBG68U-3;D4P8N+HQQS<[
M9S8\^FJ.da?KO?.c(TI.?[0>fW(@\IF+=G]?HceG]-(IFNdV33K(E4/=Z?Id;;a
QI:O&(U[@YC<RC2K8UQgg7e.57-(K&DO4+a+9Q>2g51c0D&g?Uc1]U\K.D.-,?,4
/+XR=XV(],QOMg(:0,g,CEDNR2OYF[PN@-R?XdJ+DT/(=^K/P1e5M[[6R<D1dIOg
LZ[HL24W8RMN5dUZHQ2H(M1Y8S/R,\\I+73gOV;;CL6AY]V)AG;Q)UCfO.:-b)#Q
;#?EUM[A((7S/=4^b&R5/9WIS.eY_W-JF70&/3D,VCXI?GWW2cV&R+9gg8CYCH(d
,-Q&G8Bd2HXYaM[e[A8MHCS#A@GYOJY0181;&O8VIb]Y.[/H1UYHDd1\NGSJ(@f6
3O@-_GW=KACTQ_8NNX3IL)#>e9/UQ9g<F+-3U]&V^/#Z-#_NOaHg/BL33DA>ZNS=
]F3E:MQ^-9UZG#,HIcf?b^/G23E3f6:FS3,4#HJ??(DR7^S^D9]5.82\A=Y2A-1\
9MBU,XK8/&NY[cR7AY\<M^LNMT?SZ>c+.W+>_51ZQg?F1FSG@f8>F\CbPg(Q@5La
NUAV54<X)T<eSGJI+REb^3SC,0IF=:_f9)S[QP?ZEG[?;VbaVF#JO7CdLQ/3_HVX
^6+#Y8LRZLHaBZ2U6AS40BOF\3a(=c8XZN@Y[086b+T,e@QGPZARb]<ZF2LK>DT1
KfcXb(V#Q3?2IDcgM>HaC<YM8;JL6cE,9&K/W6TZX.+L38V1-=UIENf<RG5/J+FC
WKYU_,cZ(Q=FC=RIN4)4NOF+a)C(V,TKObNT=Y0d-8E3;:Y_\U975[XMAFZ2>O7b
dWb(K)([F8OIL,7M^+Ig&>3^[T#8:F>^.Q8LLFQ+:=<BW8>2K,-G7AV:,0&L?@,,
XEMH7@9b.8Id<KbR6+L9&fH,,P:QF=3eY/ceLBP-6?EE8DSV11ZaNXFW?+[d[8-.
L6VP[Qe=K48Y+/3PP=W3#4c725>(7c.^.FNGEf&RSZS32S,fMXe:\8&W#AYT+<aD
O41fKeWHE.7bVQYf@9fb\6<Ub2HA6UB@D#BMYJ\U35@D+Da&gIB)dFG4Fg.H@4T<
;(ef<XP8FTc<(E#0,.Z;,Y7NTGVA=-GDXWER]4_;C\:R?_SCWBXHF1P_3\<&Gcb>
Y)Na#aOV6^/LgL4>=,#K,@b:X,9GO0F+.+2R6K\>Z@D]&_e;@<f,]BHD/3,8]cZc
M[U@[6<d:@92@U_H=VBgC?AE6(U@.&2:_6L8,)VOF[c.(7#aa\9>C+<M<J#_\cWC
=Z5<:TA3<>VE.IB3I.cNC:^8NP^JV,LMXeD/b8eI4>O0&5&I^NU6SUE:84KB5db3
6E52EUbIP^LP])Q3@-/<GAQ.E+_:TE<)C&&e/=K8X/ZB?F.BW]YVe+IbV2F64?_,
//\@eOPc7>f+TEA@V)A;L3([51XD[UK6C6Y#DLLO@CW?#[a4=<.;2F)XN72R#feM
>NU9bQB1.gSeUP=AE[H8KC;H#Y7-CB_.;e8<MaMR/1>7<QK+-(]AdTTZ40gVbBNW
Va37&[LG>I.B:<10C2U>#9)+?CYB5.)QgZd377NHX+gEV+5,OQQ<L3K7^B<@/8;X
b1IX]<E-&]e_.Z1((\:>BG(H/6<If85@@#c[):HdDABfP;IZR72A=.IUTHOYN0cW
G52/IHb#LCSL_0OaF,fE1Y;EKWM1X>05R2g](7BNJ;[c?f5.2T5@64?T(\YMZ?5\
3b_\@ceb2&@E,<:&2E>Ug>)([==]fRV&NX;OOaCRMaa5fI;/^8BX0YgT-G8;K[Ze
YX=7a@cRRD1EOa=a.N;@DbW0OL_-YB1Qe^S[cVN;018I^B>?+67DP,d5(C<bX52M
P(394PC,FJTc/.>OP8<2MSdLFP/8Zg5/DW<fK<8b71Q1U-=eTP((@76=MLH0(0]1
Q&M++9?@.F.E>&],LbJdN(cE+K:+0LG+-#U+DbZ#[ST-bfZ:cY3bCV8+@\CbX;]5
a6d_B2U?8#HP&N^B\QZSE[_YD=]?ZK:cFa+)bC1ea-IeS#Y04089]]9fNcO-[I3Y
5+Y/U:6:J/^Bd//2\5JNc&,#101H?I8YOM\H>S1eOb]:6HA(5LENe1<NVZ7gbU&^
F=WS^Q\&SFTBK>d6H;,)g</Z]XAKJGL6/VBU8_=_<S@880KG#8\C?CUd(2Og6/1E
A5HfNR8OE1A=B&AHdfPY^JF^d>:A;>M0=U9LC=EF=H3?cMVNOe&QOe6;U>W=B@OF
;3K1RF;SVH&8OR5<FdU-;82KXVM=]@2MeTNV4+GW&R0_eOCY.#RdX]Z/]g)_I6NG
UJ[?2-)Q#\-<Xa_@I.@9X8LHdaGPdedP.=(ZAP4)(;XV<L.G4@>13XILFQQQ1I^.
Ag2Af>MbAAa^4DX1/3852_DNWAZCWWWP63XQ\b#GbK7_TAg,>>L=VH.(3G>U7C=<
LBe3&XRTC8FQ=DLJI^+_(B7=][4g;1g1LQ+;_81L:He1@a>.ACC/^]GM#C3?>e(e
[ZX3_7bIS^.&H>\=2ga?FR(OUNP0YCXa>/8R7=]F25.OcfL=H(Tg.[,]:?FPF-\^
W/bJ_6N75J8R^[_f[-/dP.a,)QD@##M&=YPW02G#:@dD9Dd+XX8C(H,cb>F&TT.I
@_5dTLXQ.6#)F5C001c-MZdP9.IOF&f\V_Uc]QgfOZSDFd]@5_=CC_]<VND^./:(
[]&XS6T[..K/g-c:7dBQg>E5S^-O)F+-Q_[.P[)N=.@H&F1Oc42R[U]2K^BPeI1V
8IcUE2f-Ac63A<?2<JYWY,.bD#_&IT7<4cBM[dZ+3\PY#I3B>HeZWN<fA\9eebdW
_&]G).?+3EFa&(^2:=>c\;(N,d]0\EPbN[#U[9=a:RPc.Lc&1b2[^]Fd=R]O09+1
L<@4P,[bF7SPWPCEdT-RHeY)_6-cc\Z@fUIF<??Q9VcJ[-,##8fPZOQ]ED_4>^J(
W\RF#\3[gOM(QQ;;,X4A[I1b886S2&S9(V\=,=eC]S1;0:X>>)TJRY-?V@+aJK8Y
Zd,ED_LX;Ca^##5Y0g6TXA4LE[c<.4Re<DM7a/T(BEIL(,F./NE.WVI.2:b+eZF^
:/I#V6S#^BWD(73eC)0Z_[D]PNe(c0\#abK>X=QcMdK\A2Pa57C#Df23g)2@\4SL
K#.bU6\B_K1W?Jb9XPAP,>-Q_>Y0OR5)BXBO&D6RAbeIfIR]]IR0IN0M[KOHHR8^
3D1+2gbS:KMQ4BgL?P[_VN5KXb\C<AAL==Z=D/BU.ad@=<&SWA,GF,ga)T2&.9Ie
9)XFd9W4]2QT2C8dOP2H(6C^6=?4/:V:\6E1@0U\bYfJCgYVUT?\=&8(3Y()8WfQ
KKHWXLQGF5#X6I+>T9AZId(W6#4aGI(^gW-b]02U&1>VDK0&;_HM?=TGPHWL50)O
G/Z_0Z:HN(ENU_g[Q(98+eHCF;5_LcEe6Q?X]_PJ&)NY0OfQLa0gH9CB#+F<.A1A
/PS+-IQ&<#O(:^TcD]:Z=I&DMQHbZ3_2g1Sg1YC4QdMGaWJDV()=>WT>HHX@5>3=
YSHP;U.W.SQ&Z9;SSeK4F<51,Y-51KTBW+Q^d^2H:M=WXf^[CD-;>EH9+:QFF^SL
>/PJd\M6-ge<AG:cTQD[,YQKE[R+V;^\IR=]#aa3)@2;SY3BC[/URbS;]W0,ef5-
ENMCHLFNM133XcON;EPAg/61/KVSeGda<DI=cUP[-/JNf(<ff3YD8GEJ-)QJ((Lg
a5O+CRXK8(cMVeCNF@<GMc=I<BN6gI#AZK,SI@,\HY[60C?SF@?C>/a,-0+O;Q,(
DW@d+b];1+_.#,S;I:a]NMff5EZAEeZ-64T^U;;d@690@M.e;e0#^X253aSD&6S,
GDBHI)5:bSMEc\UA_TR+&ZV9+@5H^2W_HE]AP+9JRIZ0@D(\,#6OdSD#=U&fZd[b
U/5]b[f:N,BHQH4K6S)B2U>9Z[a[59I4d/AMNUZ&?#E<,?--bLc&IKR]_[^M\6c]
81dATF&66f[-^_BObeT86X=I7[-7C315Hc&B18[DW7c0]T<A/SS-KgfIbI&[Z:66
]S6?>[9[2H^VMVY;5OOc,ed+,XAVTSB;;:VT\B4@c8(9=D3^],;W?IEN9E.N?]\\
@SUMZI0+@Y^B:GPW^#IZd?4S#Sa&)bT5/O08#5?7;^>N8J8Og04=U6D=L/FUNPUf
\C<W5EIH&[X<Z7GE_aO]@,2A&]bCT]UcX9>@YaFaX,6<ReW.H=#SK4fOf]@HIYP(
^@.93>UQH5Lc:L/cMH8#DT2&RR_:>AQ&aC(^#6^Cb/1ebEFdgWJ5X,=B;:\e)HUL
Z8L><CP:8&EZTQT(/6ZM]N>)?dC81OT.\OdR1LB=JA^0gE[,-NFd5S[WF;DL()WM
@KZ5-JJ5WG&>/Ve(E(N[=Ic=,:X7ET.:^:-V6</H(eA?T5G5:_N+9cD8-5_8gP4S
;aD.02,L_:4b(eXG?0JU;TZb2??9NXCH#QF+AgbW<YdX4NWW:R>=H4MP_D0[+-DK
K2Q6US8M6V,AIP(\R;037c++cJN7)D\9a=Fc:IS72T0[8aEI@H5VR(D9SFJZCJ5^
f+EF#,LB#;AY?7U.&4:C5\6F24c<MaFW&De[Q@464:9S9NV.b:M.=HLOb9M<Me(N
HKDYP@N#KIC@?8BB0E6cbf40cM=W<9;-V@-^9I.MTU@_ZZbWeeH:1K5<=2II=/#S
,^.M]&RI]gSQI,(JDVF_+8)#+Y3L#CI:Z_AE,Wf-f(Q:S9FJ@NgR-YD3\DY3UK\e
=05CL50CUQ,HBXVZ0f07N[UB:-F(3dP;?6#RaL]G4df&(=SJ_&,;Lf[(LXZ+IXc<
572HG._@X#\01VR7Tc]S:af5G=d)A.\A<gYHeOW.cK[@J?77TY=(M7:I6NUc3KYa
5PIN?K)[f;ZF)aNAP_Y9C>O4G020e]]XML/5XJ1G@8SUdB94C4M4WE]2_OU:,eW]
Q=WX6L90M8c+KU:ag5Z(fLC4LB(ZBHR#DG\eU3:gLF):U]>9a9I[=XfFD;JO&>cI
=N@R4@Q_UT:OTgBA+#.fB4BJHCW:3Mc1M-&+5>#BRX)P;0V)G6EeQ..^a1V:af<7
QgBc+9:W8,&@P=+I,GJ&G+=X>NcT5IPR[fYR0D,.8EJ)TI9SPVUZc@HMV_0.cJ8(
f<KHdMOcCCC.)@aN=-6MLR2D8]Y)OVH9Oa2_:F317\T_R#8XBGX7?RKdCYSg_bQT
1Cea9QHUH[]C50_V7cQW=-14DIXI@XedA&cP\8E^2+\S\0Q6>63<f)OU^L]cH1L\
0D:Cb]0gH.^JL^M@#79DP&(XGMA(bAB95fMNO11UT(#U,(V)G7BRgV8)RG@RE-[3
E+7?>TQE6:1ZX5ZGG22?OHL5@^>b.f8C^7?^H)<UWeMa?4aUe+#cdfGC.@aWbR8;
:E-X4Y]=RG\d3>OERc@CJPRRQLJ=daSTSB.N]cYX.<T[M.SYM.EId7[>a+M9AB],
=+8QJ/QffAT]W>I7I8aH5aEAge99TNK4V&UX],58]dF@>IMc,K_@)SF@>CO,3W#g
3&#-8]Z)bAa0.9K;DO=gR><L0egRfV&=dF)\aWH>f&NOgG\4M<3L>J:f>/+E]-O:
0EZc,Z^YN+C&\,:gg#LGTC5Ab_[)1;1F6>WEC?T_0V-IVI@/CNVVJX(\PP/\8RKT
caI2B^?@+3)a6<0+?SVSaTHOd:Y/-2KG1:&@BV;9D&I)WBU(d.2QV.3fbc\-HK]Y
GI+NC9K&QXD<IbdBJH>5Z,R]b3CeR(bK/DG]5d_;2QUSTX(PCBC=eK_P#/W+c]Be
EeO;;-H@925cT8-=LI/03DT&;CV70^cPOP)dPQK^R=TX3=\:6/e0e#[&YTO-d,=^
R6Y+7eJHeUA9?+H.:<9>MH-;AdP]fUL@&9>;X@EXRONB.U&Y.R>f0fA;dBVbcYD^
.?_NUPQ2W^<IX.)H8HRDZUF?^JELb,LL?4IK0_c1ML91P28[UIRFBEB&]]<):91d
T;@:Y.V->bH/L>@/P?KKeFd2::U@7Y6PECX<\cM?J2T,Og.4g(0<1Cce(77]e5]J
eK1T9b@Y/E\K19+LP6FcPV@,NB@KJ,Z0NfM/d]b0J\>=6_]8Q.fa7)SX_#-;EZ;.
Z\gD#Y?<)VY,>3<Nf54&e-7IH[\DX9>](Q-UX8O#LP7:L[F[,V92=Y07I_4AT0C?
dc+-P9F\WW,<L/W(&&9gRA_Xc.T-(LE3ML(<J,VHMCf\L8#J,@;5a:#6(b8Rb[)F
G<T0T,WX>JI8A4:#(]cG.M:-6S3ETe?GB,_P&7^c2[+(<OeK+AT(AA9CKNcH+abA
X6S&g/R?0\/X<O>SI#cK)N3I^@MDcDK>8S#cbFR&1CV[ASNIaI8,B=]H[7gb3)PP
P^9K?\XNN6NKEZ98IX09V66M+g(>QLb.;XMTBA+LN\g3O]c=Fg#.I#adCN;Ef:B;
)[)Y-H\4@C\-Of_74-d)4gE&^/O?FYE9dE,?af>>^#=VQJ;+QWF\I.bC7U9Yf-c.
A^87N>#BWC8F5,XF+Q2M[X@a\I4,8<Rc\Ia670360A[?99M5OF(-64O7P+bGM+9Y
eR9g-EOA:F(Z-<>7L^YWY^C^P;DRe7#].#6DJOBO=3IfLD(/e7G^&B#7;gL[__RV
>VWBF(GF.Z^:f2ZR5<@K#1Qg[;f.c]<1+CL[?Y68PG#H&eZdgQ96\9)]g+G(a#=L
,gP/=fVQ251^U9P&<?>CTDIUY,,1<4RZ>A.ZdeB696AL9F2geD2fa8.6.U?&5Tb9
5cD\ORIU?\6H/P#c2RINg_V12>_6Q@=NIdMaF7.;R]/Dc#SMH9BXc[VD0)Q4LGPN
3EQ9&Y-ZB+3cPNU93a&cC35g^7V?5T;V?##CX(Id3aAW8:N7_A[LLEIg)@9VS#Vc
;B<,Ab@9_XZGRE,YZQTO(e-^UYWXf>/HVLVLU9TX;FO,BB@VC(LgRU(5J&3G:4Ga
HeE8^<B1ffH5XT-@5&FKg:\-1>#MIC3:2a^2K?U3(<R(I^EP0\:RYK</_/[Z)M@D
)#<833I9;cEJ_&Q4KL:0P.E)_GJ^XXgZ>QBQFRP@-WCLLPJ;Lg9]<1b]a3b-S7\E
KURK]ST((BJ;4_GbUf,\dK(\[)2WU1QA(#ZW?Q=D=E^d063Y#Ff<cZT5@,eefB=2
a7QQcXH2Y]bNd>L7<XFHWR<d.Hd2:GHP,Z/0.X[MAIIYd6P]-Ag\g-I3JB,<5Q40
6.:F9JSRKG=F9?CAG^d:ELTW\6)8=+6,C7V#5M8A7K..>?XOVKPL+9MF0),(^D>S
Z]3eNT+L/fM56T=;.P00/>RF6(dM@eKg\>_.FXDL_AEXF=BA1fac\67>:fOM>65W
,W>]R?^WLZ\S/JW?,]QK^D^,c:]1VgS/S^E_g/]T:cU&f(IW#-\Z7CV#TaK_F),=
J5-0fT7HSIObaG=Se1CB)HBB1KU(\KcZ40;R6efUfMON+29K_LI)&^?5<[Kb02OI
HOcT\&4QEAW:3YDT&B1a_(+Z449Z>C^O\_#P(8[6ALP7^^[PGC;)(fX45;&fg?7K
N=RT4?g;2H8PJ.5OfH;#6.TDC<-OaDH-M]Yf+N<I0\6bIBW2:MeY9RD\[OTX@cNY
PQIQUdGNW4^H818+2.7FfHgZVgT4O-GT5_&N/X._?]fG82(SD&b+7g&DZ[L\1SHY
,N2cSVWD/6(/Xa55KX3#](,2.G9O&QGX6GUHJ2A5#-NB#P9)8/e)Uf>_+1^L[5@#
QNM5L8fO81#f9(=W8U>bH=19,)cBaW?+.[#e>N18(e93F#XI<R]3XLE_M@W;c()<
96<4P&2F@N+T/=G=KY)3c5LDe-<3?bI]<Yc@P2-.e9WXbN:6+#[1?-F=?eI_W;6C
DWUUB32f?BFGf[A7CJ\YDFBL[DVMEYI+65W^+OHV)5;7;1cZA#CKBI+LCb6>GV:W
UP2AZ/W<8]XG[090L9g>7+SbbZ_F&)[A<GfQ18TO_g&F-T7Z5BP4.I;N<]6->;.(
MWJXb)[P;R&_0?2A-+U9MZf&cg,&(gP/8\4-[HPVF1QR@??\KM+1MV4X14+_&\.4
Ua]]H@V-B_WK]BK4D;Mf_6<V)eN#M>4:S&1Q-S0.TS33:##aZK0)]JJ-&^OIM_Y?
RY#fbLDZ8=9E]3V0OecaUZP\J8aB3\5=3NX?L/D&+9;LeVXg6(N5/M.1,(W.NLY@
9LK1Y5I-N;@>#TDCG((08DHdRN24DPc]0eJ\PWT?Rg.:27T&/H#@:[LATYWVKSXG
A^=7P&GSX=Q1F?EYQ)1Ed>,QOa3BTD?I;I1])6&Vf4(ea:Y.BYH4\\7@DGD)E+\&
8D)@3F(]df@K@O^]>-gM0b,>+,d?ZKbIc7HdU,F:#d53DP@.a037_4F0B&a#.[,>
\K]@,G[-Eg:/GEPH:IU<<4O/7#?d9e6ET_Z9_;W(X,@TB0S>VO.^U<f/__D:+Y.)
W;6.#e?-Q2<e(ROEFYDAPfZSP3XX,LYa609TEHJH038QJ80=fT3g#=&R@f#9,ZKd
:@4KPOAEQa3bQNL6_DYfTGUC8Qb;LC(WZKBa1;TUN^bg-be(9[Td:Q0EdN#;AN,Y
009d2fLf9Q_I/1))IG=+1(=VV\NT)<D]a@ZGAHcO9LE<b)gX@DHfVY/.<::(Q_/Y
N?\?b8(FT:UQGB9:JH8S4VZ.)/>.EXBgWD_D>Ub\be+c;0WSY=Q4cQ54..+)Sfb^
a6,4Q79N\E9UMZ1BA&=g72?+TRLHN>UWU&FN0fN\b\IKe^PTM1[18adD/[@bIA@e
FbaC81=4G@,[//<@=\?#/9>(a^+OYOad[f\c0-/21)^_\;a]4]A<&+38,ZcS:UYM
E>dS3.U655RTa)#e-=UR@07T/_@GN7]JD0WM9@#PQDVF43F:7)<<6\0E)8>Hd1#_
5Y\=>@?S459V<=XaK:N0D3<^-(@PZc+dXVXBg\Na&U.)_;M1;IS;472[PVP^4,c[
=LF[Q684>?\<WPO1G:RGRdG6Y;;VG+K;E4.A:.S8)4IX#FY&cf0bYI<a.O\=&Vb1
Z7KND+9_CDX>3dNVJc9gQ+U^WRUO-?NED\+BP0dO-.ff8IEPPeXKLGGZDW^H^V7e
(XXJ3Sf&fQF8)dO^U.4>C[^^[7868S.?S0d->VcfKU9K<AgaAFVaCEQE0=)5FIBC
](+Qe)I=9I9SYI0\>^d0.(3]L@<IU,0EJ)1>A\Qc_7>L5&1gE9[B/bK9.K#6K[7B
I?A@G5=;cdB\([F]UJ7c^b-Mge(++6gXXE#(PJ7A/T7]X>HPWYKd?S/AgX;ZJM[T
Q2NXO,)UZ)RMEg)Q-X):T\c+ZKa\W(fI]XP,=PT\df[[^Ia.7^M+DFD#0V.48O@7
B7^NWIV2aFK6A9f0DK_a)V,>f(:f-H4A6d-2R(cTNga<ebOFe-VeYMP;0C\RX^Jg
Sdc(D8?S2bREO(fM#UaWSL9P-7;;5;JO#&C^6QI02^/B9/P<3-E+S69+Hd+C#M#X
bD2S9e^\>V/ZeXdBNUXX]>7B=2/Ybc-ZF.,_5b4YVX/ER:f0N1RMG;(?^#ZW2+9[
aIWb>J(d-++b_L((DVR<+PU6dDa90[Y5fg4BJg&b4C+^O</c[QJbP=EOR]4^_@]F
+<>.g>ID3f]932=bN4J77)DJgZ+]IMWbX2BAGFX8MNPcK<I]gV7J?@FVL8L56LD7
.IP,,:)45EO7\=RDbPI:Kb?F;1^^@BBC_HPIOH#R^_01DGd(gf03^N>1T6U#5IR]
5N)(]=P9)V2BC?Z-eO?^5?QUW#OCNK;?gTeVEF.;a-P37&&<e8AWJ=0W,.[R->JS
27AQ>H_?C70KQZ<.;.W&\9>[eR,NSN@?LfR[C+;S\=^KK#9KgPeHT095W&M_:2,b
Cf[>.=;3YFV-(<dP5-8IQ-O7R?Q<K&3&Q_T6NUKMOGT-9SaOF\]0C:>=H3cF@SIY
RLC9[F++K@+W\?e<+646b-,YE^1Q8c>#FV+1A1S;e>X7F^HHB4=Dd7OAW:<;CHb_
BK7D;2Sg2NdT4-^G7PL[V>Mg(4:EfET+JX2(=#5FP_;Ug.IG+Mg86\<19g5KM3=J
A)[6DNc)(NW_(B0S7DJ]8I]Y8e@&bXIR9d&9NGaV][:-0A:Q.Kf?,JZEZ#/VI+GL
O\5L+abd;L14I]<&=bIRgYYXIea<Y,Ma:G(S3D;PV;Q(a(ZbW5?Y5J#QD6PRaVQX
93(b-3XXMSgJ(<1]VI0C_AVB//S);b>F#X0KR:DRBBIO\-H/3S:+V7PRdR^D&G]K
SDYCEWS+F4Cg23\(S[Ia&M=C):Nf(W/PR=d9AZN)b9TH7:0QfKc>g=Z[[895.6UN
R(Ce:U4D/f[O-328=)ZYY#+dTaO36Z9G&NFCGfXILE;Y##/KF5[GOefJZg,C/dL^
#8IQSI7PQ@L/dVRB+\N;I6Z(M/IcBLM_=1U8b-+c[QFH9BX8J/>9(=bd1.e1QPHD
Eg_<H7RX9\5?5C]CV:WgdQNg7.>M#-Bf84BP;R1VaU_EF,&@=]:0>/VII)G(f:H1
[\VR@D(:,K@M5=;.K,XADO/d.)-;aK3fO#8#f:<?2X<R.U\\e3\dM9LLT0\]-?AN
P/a:Cg6Y8>d3S8-TCW@(e9L^V)B7.Q@H30Me)FZHPcI:^>R(bP[W<>R-UIUK_?B)
3A=C#]6e)Y,V[cIb3>[0KF=J^84X^TP<6TU]+cB.62J./B_W4g;]/[S,Z\[RWRBQ
.1,0:Be>>5_0T>aU2Z>AJ?A+\IRV>bWO/dI(?QGc:S=^?a)JNL6V1-2H303LaV2+
:W:2V2FO#<^07U.Z(4W0T]E2Q^/G;?+g7U,[gK3N?&(@]77Pg-7FGPEIcIHRO^<Q
;U&@U#?+L(_.\#g^5YQCOY8c(UMfF]PfR<@ae.6JcZ\H8AO\BM9I<g)(-S,_1#@[
Z,#GVI-a=K@#FAO];P0[f[-NH[P]R@cH@D+dCAWQ7>NX8(5;7A]^X01N4LLK]cU/
\UY-1J&);O@-dZ((N;?M0MMVJK^-WP[MTBHDH=[V@Z>;b0d_FT[;(@X\:CCDQ48/
,OC[P3JJJ.UUX<C[+A6QaEf=:Ja3LdF5g2X=)bMf6\<c:Y-B#OX15<gY>EL_cbf?
368#?_K7ZHAHg?-9CIHa@;LcUA@0?THP9bbKXeVJT,3[[;T@6R94UBc84^/F^7]e
cAe^J_?F+7f4A@Z+FIFD1[a]aKgUA)fQgBAc]US4g^Gb3:YS+bdaHQ0>_N/UAPM\
\X^E7TW?gP3U.\Z:CA?G+)OR\8H[\JU5)_\a.L79]#gQ<gS-D2/4&GIF2X+^fI<e
4WJ2?AL<PI3[G3^^/V4/.GNR8<daRM;<@a1Edec5+K/HB:]M0@e</6K-BIA7c=94
YbB-AB]G-g&DgS+#-8J)=M=[O4&AKaFX)fG3\/2:=TW^6-EaFOMSB4M<IET:\cUc
RXB6UD09+dgb9T@:0#X[X-Z=WVL<&;@<:6Y_<VI7+TI,dGTQ^,53a5;0L;Z-A-^g
[X9/[I=1/9:1IcNb[U&(.(_eX(T,T_X_IK9e:7@?O/I7>JW?,M41fObdBQ9\/?3=
b2^^3H?//HWVDbFD9N?^IGTPPY^/=.<VaX?@8PGeE^b.e)fF(E2]FJEd>IVW/5]2
C^QY,&=JAW0>,(DT_C[3ZR8^P=JBCA<0f+N&.7U7V_+;eBeEeK2?9@_CKP[\JDBZ
6WA_=MF/O)KY(3/S[FA#Acg:?ZP]G9KAM>=?WU_A9=>F6_636fQ9>O=,IU>Y,IJW
Vb,W^&UN^;)<[Q(B.K?N/DQ5QR85NC8IcMD87F\@.84FN>WOXPgZST@YRca^/Ha3
1<RT+fM/VJSM:3;:=;B&eSeN1HW09a9,GGg]BAX/G++-Q,3_:]3_=gN#+E3+;2(?
FN^,Lb.Z]f0P]]/E:7=]#E-J,H\TU+M-(;-JRcdQ45F^Q;EP4FQN9?d3<.=5,dW6
7E0^.[<B]D]>3Kc@DZG7CE92E&Le/?@&8XP_JFKd.#&6d@)RF)6_^?N\G0\BEIEA
Z<IY_M[5/BT/7B7DJTWCf,dM4gE56EceZES&L_63UL6;2K^O?SA=/,X5U#AG:F^G
86H58\-\-UOJM0c:;:2@]JaIb:.:YX+P@;_Nc@9XZ37g8<d@bHX6UGZBV;(e)8WA
..PL/:?.:AKHRa6,.A&DPAU#KSGV1+e[CS1Q/7:&\)1d44&K9WF_g7a/8#dCc>[Y
<[A^3OAWAe81&,C2)RPC-AYJ(>gIXF>S8-FJLg^BLP:JFF5/FTH(2(0Na,;N@\F+
4a5D42(/F]W8E1e2O.CM)=D-\#N^PDeKIB5UcPfSTU1Y30)8gY,9aSH7Zd[&Z[/U
)A7.F1)2E^T],#(eS;<[f:>+e0^KMXaF[YR&^^_fa@H#[LDBIR9c515Y35#=Cc31
KEQ;FLDYJSb2=M1\+aS=,e\N=2cFB#?L(D5\3>_D=;1\[&Z548CPe(7gd(Q@XN86
T26E+VU\MJ:P^F,FbVc,-7BUWR=4[Y11Tg[U\;1,ggXH4=Se&?EAO2-[UP5[1PQ^
acN))/f)dI#D(c1/PE]_QdDcI?SV:Ia1IJ/)>58DK\]7H\(:PU-MEV39@Ig<DKVb
MI:5BaJN(\PT.5;N7]4OLY3M70fL@H[W(>WP/H<LWVXe)g8/_W)4Adc?c[.MU>f]
J9CFD)ETa1/0CddYb(/@ca8<WB,PBG.)\7#3#+)CG-J]EPR,ca+3X>WJ?#.;?f\E
d:XHCF]X0I_/(YA/fFP&,-::#bdKUV-cK6PcKX7(XgEg?<M[ETKR]TR)bP&I3;^U
FZ>H7A]]VOb7Y8MT,\U(6RX?cY)YDQ)RP]#]&D60PAV/\?)@e]UH\D.LdK)0QCG;
Y1gFA\f<gN-MIa88.?R1?7R0b/]d6S@?1;X.P0BRR(_N+#]JFHeD3]QNb#+a]?TN
g>CgZGbgEZ.UEf97S6X4@)4Q1_RWW3[?Af[-g<.](U9Q.64I<:R,G9Q>gEWA5SV:
L&:DHO#PIB]?WIDF=M.]fFMR7[]YR^5ZK;\&J]Id+Dc[O^#4H9cW>#aFc<a\g48(
]P/C9dLUC?64\SG76FIH6Q@H<):;c1CB1;4W9V&DM/_+1C=X+Z]P9AIHE1dJ?D6B
Q.#_OYQNO4/B_:0(CT_RH9)@R9+[5/?Y#E)>CS(G/K29U^><OaR.R=;X4:ggK>LF
P=UE:+ZZYVB9(WLC430E+R5IbYJ_6=N0MH92VP84<Y#M\L49:M884]=T@:[g=>2b
7JCg6;aQ+,;O.?TPVbeK\G;<2[SEUFO\bJZc79L3&<&_N^]>11\2X2:Eg;)F81A=
&DIGIeB[W25F+Z06,\2K]P^dXN]>?F=_3KML8:L&:],BK;P@/=UfG9.J2VWT,SEV
f]((9<-;R>#@POQ\-YF3g\QU3\-0JDM05Z<>MXgZ2[TXM^,N69g8f>>=Z[AEe6#8
,9Y,\2ZMR\fVQ@:TT@Dg=FQDVSf9S=8;MB.B6>6\D?;ee6N8LW6>(THY-:<9g_\+
<;]:V_#+4H7JdceSGNA/\88?6+.8W[E59FE71UTEZTD5(^USE:EcPI[HWE2@.+-M
Q]J+JP7-HWSWK:0B)fUIQd(F(/R/(O^dH+45,)MSWe/<0F)5E,F3QEJ+HI6,]=+X
7:,Y9\YcQFCQ\\QMg<5_d.H,2aHE5.GAS5(OOCI<aIXVc_Mf3-/SV0D6K0dbKWU[
^#9+)/BT^()+0\??HYQ7)CT@(A0G8+GF(_O^J2V<?UQW:0=6UJ^#B;5#5A5(Y47^
9-GA7Q+1(A,,c#\R][93]VU74FV)f5\)MZf-A,Y@87,0I9TB@c(d:N-7SK]2Xac\
MHU+BC#HZN<L2QB=c5+(L@^BX.0A-H_H9#3E2(OC[I4>L>;9\LSQb[b=&4M3=@)7
)5V=@BN,[d3++)=CO0@;b4^]:/K19\N28NOAb@bWaK^Z+;bLJX6V&W-S^L&+=,S.
PJK)YSQTgbg:WaN&]>TSa@0J&/R.C?,)E0^;D_?:L_==J0M++/)(?8,[MN\?_eDN
e9XYZ5=c3+_Yg)P]Y6HE<cfde=-CAO&OC)8+e,2=aS[,B&IQ0_]ac7d],O+ET>U#
0^8-1PX<R.ZCcS1aK@H<&5A[5@)aeBbb4?PPUXf9AF)0Ab-WT5>bdA;MRW>bR:Hb
;U4]-8e+UAJ(=H)FB<I5\F\\7Z3(A<U+QdC\[[fMF7W=bS5^S=V?dIFJ0>RE>XB^
E7F7I=]XRZ()L(+WKFL@X)f^^:@S4F46:bS#dTSOU5VOX#8UN)PNEPeJO+AXZ44S
3;d+_FZeMbQ)7?9.Y/Of;Ef9H/2?TMXJ[GgZTdHGRTNO</0<4VbTW0B#=J/a?:6_
-?0?QAd8Ae=DB+N^=S59)(.:GcQN^2]T\[H2b4OBO)f8/^83?RV?51_]MQV4-@N?
8(3JM;N=G-+]@<f\L@CR)3DfHV.RFfOb/(e^2bWM9,,21<JBPTgL,eD=.IP]Cd+J
ZKX4.Ff.gL>#D@7K_<WJfAMfO(IG^(TfVR@Dc@CA^g:V0_IHUBfFVOIR[T?=BNg0
1]2feXS]d7c>/eMTVS?MVE>dAZH.(N(==3[#7I3_GJ_aF)bBaZ\XXV#cH=MZRdeY
0OQ,a6:V7?(/cVV;]U.c=9[^LJUSSd^B(3X3A^bbJ9N><\[-c)/(9b[SVPf[(&:]
HPF;_cT.47AC=.;M1-R2>PUNdH,A7&>OS4>B-_8\RPCX>8<=/4K,g1QC3I.cLWE/
I0d@4PO\[#?A[.I-)d[Xc,f?[>CL-M0@4(b.:^2(Od/>AV-X#,KT;ScD\PGP\49/
fcU#L.#cQIG6S51UFHXJC@?[RJ[fRS(6X95JN<1[I=e:\&8[8+^B97Eg^_[?#cP)
Xg[/a.^77E;8N9=f9Z)J/\_BT0?Z^b#:cWK#TEY46R5gS-Ha/DdeE?F6c.9IPbK2
]E13?PTa=KaG0aCA&Z\g+=@?2]31OMR+I05/>Se,R=(J?#9A[YE9a3[0._dNZ9E+
?[A(/B>3AgSP#B4OQBTH)NgHFV/?GNY0LZ)X#<3_(XJ776^V3HU@Ea:OFBZLD;VI
PO+)g.DL#Ig9NVDTX:E^EV&c@8T#XZ??&UQ3:@RY>CKCSS1--7bd]g)<>+RLY#7C
R@OI>J<5a/[L);HUU;HX/[WSAKN^H3E3WSb>#:43Z>W2[#.F?,0=O)Mc-[8ESaI7
=F\];YVJ;SZ<d#fZ0H3PTe60HT3^Ie-<WF4f&7Z;H/7IZ]3-SU[KQDUed8Tf:bN1
.?dV:LTULD\)>10cW+X/fgJYH?E:B-aXN4G:0XTb0^RG82O&=JDF&;/LZ_+#7;HM
H&IbQgRZV_aRId46eg2I;<-2YGQ1=-QbUMH^:2fZO=.]=UTT[F_aga5ef,?Q)-g9
W8#1&=6HJ/5MTcP=,Mf,a&Z>.ZA-A<VQQH-44eBW@e,3@@?(bHKK9BF0-DTF=;[;
-.?)6Xb27eXMZ#/M=(0XPYE9K9RdU;@T/1U?QYNV5[R@eePCF=CD64)6IV9N:S@e
ZXT;V3BTE+C^S.U&I;CeT+e==;0-;Y[+-&330Y4Kd[&^W85XQ0N+W.Z6,(W-TK]#
5_TK::W_F:2)X7Cd,;N><WCcS4b0>3H11P&,EXNMI=)N4&NC/_0Y3K2LAId16Keg
:cY:dCQ>2K.L?;F=^LM=X-Wd:3=eH.071F3G7<WcKB7R0^VAc1L]&3C5Ya/WOH?7
87,O.)@[PFF/PTDP(&;;0<B0Y,.0D=/:b\Re+=[\0eG0L+NGKf+g]>1@I99Ie#c0
aHBef.86U>eYeI;?]]CGRB8gM#):)AO_cVT&LdL+5W[[X7__eS#a(B.1:Q=.4J/K
,2VX151XL^9=fW,M75^\AQK7;B>ZY:1?DI9D<9W.?5A[1YBV:T1O2DBbVaK]5/XM
.RB)NPaKP&2E?Z^gaPC0IY(Jc=[CD@&PS>VZG>[5Rf^DXc)_Kb>a+K&\gTaOPE()
-_^5)LU,613N76#Sc?^P\\2?B8eJH#UW;M[8</._4f7\\JK@.,/^7DJ5\V1LTJA<
228VN#c4f_W.9_>-[W>3&aY^Z^Nd)D762d5dLJS33B[#_JA;X4J19U_(^#I.XS:#
T[0HNKVJX^=Z.V7NC9689Hb.Q6:I+F]HR8327eDY?\Y;SaR[1@aL765Z[+U#+N&?
?A][:SEAad?78IF:DS.WOO6^fJg(S2Ie@@T@WdS@TeBPA1:P6g/5A7O?-+PIA/a,
WO=L?C=LOA&=)-2-<G/A:KH@KDI.5(F=REUQCLBLH^K)Ca=6dEX(D+XE27UBcB0C
_S\TS9eT57:cg_4C@0B_RgRT_@=U<OPZQWL?CTDVL?E90e4E<UNe&,)3,WFRecP;
-9EOd3.<R#F(<S7Ud\gNMgLVQ[Qd]LV0;NTb8[QUHa[d8LbXLU<-/THM<(R],ZDd
:d3aN@;@W4\M,:KDV&cUBH(8=FC)90)L__TY(H5egcBFRPGJTC5R9[[0Fa#.eg4\
QTIc#__ef\-JZb2SRLNQ,.Qd3Pc\V#<9N\\#J6<c>8DK,f]64aS8U2A52IT@RdcT
Y:+IR(9&>)f3b7U>5,\AH7.L&RA84ag&TPcXPQ-?cg&.-3VLa9Iee9J@eU6LQ\.O
W1PM>BbN+5^[.8ACYf>](H<cIQfHG=>-B8MJNSSBRcF?Qf098Q(#0JNY\0b3U8AA
(La7SS4OZ0#IMUIEc;329HHQdDOBTD&/K.SaY>7<H9@J/cK8DK6#fQb:[HSXY>+a
,2g5J/TTEK;E)bE^,2_0b+66E0V8HK+U=]F8X^,#A3bB=;;PI/LZ+00^H(#e8:6[
&6.D[GS1T/WZC>IX82[W,>=0,.Ef?:[.7QHJ<UeU>0&GM.L=4b0L&85c^/NI_;GK
/A4IKf]S)Vd\=KHXOP;LAdBf+=d=0eK0K4]1>CUBZASC8+Y+?9=+)3UZeINJ0W_^
b\2e9U5b9,;c&X@]#5)ZHQYPAT,A&Q<Sd/d]aX9P/1]c;<DQ_bTA=0[[M)a]]f@M
KYb/dRSdBFZ9QeVgCb1YLbZ#MX=8UE&?IZP>E2W29HI3]8@TMH\\,+MEebUUd,#/
=B#WD)=TJ60G0]C>-(a@fV7V#>K_#LYeM81N)L_e4)]ER&;9KUSP]ZV9H\VO_@:/
aN+_@J3e)2F&;),VcR#[/SYE_/d0GQ9ZVIF@EY:9d<[.KUg@@+R,b:2&=7[/I/S.
Y.I6db0=QF=D\OX7]BN+).AWc=I#U1VHWK7I@&GGE1S;Q_C,eA^R@PW>a;e-TO8X
C9=fM_4:(FS55;a2Sc=?4ZCB/(>AFA72#)b7Ja6fIO/)a.94J7]H:(ET\#)8^&U]
]VO?]XL?g,JH;.K(LK(Q__EO8b^8+SJW]G=2:bMK<PTNS6?\K\S:DaY^>BaSL6YV
Fc][\gG]AK?7.Q5X=P2\T87^VTe52&VcVM-bZJF^?ERXJgeLA6a:QF(6DZU>d;T+
5d1SL]EYL?Z_))H#Hg2,ceUL[:9VMXOGOY\]d<GaXGU;G7Dc^,.M-Ne1?/QUL[fW
Vc/RUP:e4<HK4.X/N1?8(;+^DRX558&7N9+9UH8(V/:Je<MFcH0)[?Z^D9>ELRbF
dZaGX1655LI+dMV-deY55,.-^BR.ffVRc_-MCO]A(VFL3IMIMO7a/Z?-0WH/5PZ3
^4E=a6N;cY6R,9S2IG2@-&6gcLaU&#ObZBUJOfS\5<FMO6aL;P9+RD)Sb=.02[5G
3PFd@:RB3CM9_6XdEKZbDMd?SKa\YFdL)QP/IJW1a(TaHJUd+:>bJ#\=MIXaBGYJ
;ST<c7]3;6DcE-&dH+=@QY13D:BWeJU\:.3E6>IfP.TG\VZggfG=W<6#/Y/GGV3B
-D6KGf@Z2@OWEE3gY@S0VP^7<Y#WO3OaL(9-,=;#9-DGA0b&2)T(bOIfK&(=+,(,
aG5X[^N=2PQe5?7;Kf3)?^_4^_(dT/b?__]#dY-.6PeO/X])E[#df.K8Sd9Y2C.e
EgH9;5Y1M<A3PZL\O?AM@fa)U6>Q[(W1R^=@(L3?V>+0gB;2VY>0QH)@e+CJ5:>>
HgVKDRfPa2cV+3ZLMD8K,ZRbb5CK<ZWMVXC?Kf4Rf3])^]TXf6)]WE-DDV)PHT5_
RLIRWG;C0A/g5d+[^GJTOZ6N+cN9H)d@e/MCLMSI-Ia44)-XfHgE,Vgg,0#(T_K-
&XZd(LQ+-H&f:D,,e&gI8b?1NX3Y]IVH]]6P.)Z;6Wg.&(ANW)345#NZA-KNM6gZ
+C&=>fT_0A,CV6]=FTV6W)RCLOF7SX]Z3BLY6@,MM&UP=A/W1=cFUIBFLc1[IUfc
-(21D).EgTT/,+7BSNJ^EZE43KK2EF92UNg3DfOH8EZ8]PI[W@F5[dag4@J6^NEI
PGa74RUZ9V<<7b)AYc;+++c?N07&b>@g=/JF/e4PbfUMPBI./HHO7]DS/QUT9,,8
R],)g)8&3\NaHWVL7G\F-=0MeeFDT6H[,Hd3AQTNE+2382^X\CZA:g1JX_+E)-H[
3\,ZK,FPWIP,K4^CSLO8+cW4S&d]&#]2.,TJ<YcaCHcGYFTd2_FT@JB9g[(<V#@W
_46Q[C.7=8FTY+39g]B_?/(Vg7G/g(AU-3Z&g1YVP1E7b/Le649G,,W?OWXd7YaT
c^=&0/;R,5]B73B/cPc?G2L>6384F:L=+=?S]V3J?YS0e23QgC9XZ4,W]4Vc_E6)
GJ)J:-M3J3;WJB4.^Q/WXGC\g..)7Ob^-gNfg29d30_-\d,L5A@5Ya[1?gC.7:XV
VfT8Jc=<7;f>A+A0:c</8U7JUZ4g0DT&SXfM8?\g)0gcL>LUKN)U7(&=XbJWDC9Y
8G1-DWM/76;2cXV:)b>(#?ICfN-,XYF&P+#8^O0VI<P+19#[1ONb@VIRO(4g3d/<
UJ&O)ZD(_,8#g,[==RAF)H)8X<@Jg&5f(0VSbCO#;X0@0\HN07/F@>^.gJ?YaK3]
Cg#f7fAFge5aL2#BM.7E_FDH+EZH\?@5R+^]dY>=;O=F>7,EE]139,17(O)^XRe3
=M0UN,::^[36:.Z>G0&GQ32B\W39OOYF+]9#0Z0_.8O4\DUaII9]efIE<1=,1R=7
FFN+;1fCR(RM53Ye?d:7+ECLPWXMPY?]Xgc9Z>0X^\D0#/.;?B6,O4K_c_LK<d]d
e^#BPA_WHN@U53d^GK8R7MV;?>6N<O#a]Ga,7c;e/fY+H<]bRN8E0??C-)c0c2_N
B@=JLdTLHWJ<M2PUIP/8&:.87Y>]/E/;@]1K8+O1X&:ZK)LD>E(3W71H8a;APT9]
ZV:]cMT>48VVd?>NBId85@L]7;:YfcJ<RA8db7[WbA67IVba/MP5fPHJ0JN;8Q#;
R1_[e6RRERdg+&\<P5PZ?O/&5,+0K&F0fAZS?CE+2<B1aVHCYId;3d>/7(-dQH,-
?,9&DEZ>UN#0bAg1NIO+AJa[QCfe\MBc:UW95C#ReNIc<bJEET@V2f,>4U.c^8JP
Y69ecE.MTe-C)/+N(G2IQ)BOK7)Z5Ea^7886_8>27/MR58<0XRDYB1eJ,F^X,^Y[
ENO(ODB0;2B:0CJIHcFNGQ@AK#V-E(RR4dA&:)<Vc/X2Ec#8MgbYC8gIL\6UgZ&<
9a[KA?7?:WbZ9)(,/4.SZYC]+fW9F3<8c1E^9:ed:&U#=0Vfg/e?ARYB]D(b;d?-
E?(GQG]?CSDE08[N_B<fOQc#HQI24=N^9D,<[D[[8\3//AWHNENQgK.-1E2aL.+3
C9+R(f88)MARS?+U6=5.^QTPW)[ZdP(CCR<2CXAZE?T=E6:C8OF+REZLX/?4/K1X
2=BJ/II@MY\NNW5275bADf>[DG^:e&(LT/)YWU136T_PSMEGaC09FXd+-RZ7]GA,
&gF,B1Q#eCMW:8UP_1W]F5ENLWN\U@(HMS7eD+V=?C1&Z>cZ2=CcW_dgS:U?BebP
K.)WT([58=9VL^&:89WP48Ya2?NfHGM25HRZ5E(B<ZVCFM6VP<00AEGaS@(R3T?;
WTgI&Q=2#E_XL9Tg-,Y=dZbg+BISD0-c^6<]/@GM:MK2-APYe^:>5c5VA^J2EJI]
cYNC3\-JPR]6+O6HdTV=:Z/\QGD&LN4+Of#TFK5AGG:7@fC4C@R1,]O^SQYK9?b)
W#&VaZU_F/2_K:3T5?I#9b7;OX/Y4TCDW:eWC,;>f..Z:TY@8D75&MC5g[eLZ<P\
C2<2A\?+/5Q)a][:8&a[J9P/9cM]<0J)g&U>fdgM?H;caeg8eW3Z8D\0X68R=L;b
1TRfa;IfP&).RLf?5/VeL/SdH-L\8?ZHN;OLVIEdU4+ZKG6Kd6Af^8@/6JI_b>NS
S-OW)S<gD)-C\MWHfbf:bE=7H3XV&N2A(8CaBLBH/IU?\_/#>90ZCfKOA_,2Hd3?
LbJ^DFN,9ZTa^R512SX7>8.cc5?S4Nb:;B3&12cT?L4(J^\Q#+P13B]gZ/3PV_36
eD:FW[WF0GVb6&QU>B4B-@1a?:e)0>eWI;DSZ-\W]A9,fD23_H2^,XDMYCb3c\MW
SdA6W;,S_3JHD7#S]/eH7+5-7-U?XV;^^13<T;Z&T=^J(S(D)Jf;GJb6e^c).]->
XGDff(><9G<O2GbV2MU82cS->V\<cZ0\a#82(4QIA8@&^1]390FL^f=b^MF+<_OB
ZJOG99/Dc.M?H60P.Y&AaDH1Ueb]U-5L_P0/11@C8W/SEga++=13J&HN1f#g_:9+
VBgM1SaAHC=0(RPB#5CGCSP7)#ZXFA7Ge,Ig<=cRcM/S.MLN51Y]929:,SWZTG0e
c(=e1=4(_?A3:.JDI3[cI_=RI7#_L<Y9>.ZI<KO75S3Q-N_-?X+81<&1EHX&AbG8
\(JW>&(]AW[W2OUH2289X,fX3bI\+dVS8]Y+<BTDg\=J?-#Ta:=@SD.:7aH2BM&E
^):UHS0^4C+_0G3b=[TBU_L7(#76<ZIA9Ia?N@^G9<MAT&75GW^R7HFUd#&KGdR(
G1\6,(RJ^Pa]bSc2Q2PS+>;\6He9S/=B+1-6V(>G/[B1a;ZZ=BBS[W?f)1<Qe9P?
VV=>I([W>eRH88^6ML+V=5+1RO5H=U@-&g:LPMHc>;AA.g19eK#TR0CgeH#gFG,H
B)6bcaD3]#M)+gB4Sd.:>?3.VTZdaS\U;:+bMd95Sf^WaZXP&\f8Nc4Y7/6TYGO.
d.L9V9]\H[Db=:M2_33?Df11NHZ)S.N[,)N.cU^#XHA1GSe7B=^],=:#N1P(],CH
&:cRCZ&Q0@[&=J<#af:@],V&XJTd=Y?)(-&0QGVbGM>S(IA(dT>E_a#LI:^YB&);
fT?9=I\Y<362dPeX4b&<VJ3IRefI?bO-MSM_(/>Q/a?0CVD9OS3@4NW>UY@(4USK
V3KDG60gg>0JP>0Q0:Ge6bb\ZUWK#g@MW=^JRZ(Nf067e2E.+=.^dB>D]/_EL_\G
5^9/Q<SVf)067>T#9Yf.XHY_eL<]KW,U5^QFf42-]M?L_IEf5]K=R?Q+G_ZY3>,@
1BLC.V_QH(I8D<\FUR8d?&&&UZ&G9:2WA8\P=T&gD@[9GL,PM#LT8I@P@)^\,U5F
f#\#aa5]4J-?=RV6F56c^^GH+@N?T.^QT:>J^[I4])8U[E#7QF[V+B#4@bJW<O;U
b[Jc\a&SP[Z6aT_1PQAa):b+,Y3KY)H7Ba#]+>U:PS^/Q,dS+9=J^&;6\Q\RS;\<
=[1e:Nf^O:+_)/T^@Y<HU)05_dG3AF2U8B<A3I7=RN[ddHIVBO;YOIQ24FTC([G?
9_/][3.?T-F#>\V+L)&B)Oc&d(2XHK7<7PgYBf];2<OZ0N[cTFYXDa\PV[c#3.+)
ef8IgM6Y?G[FUQ9D=/-a>LV:F&RR5O]=e832_FNAX&a:TIXJ19-:S:SKCK7a>4/(
93T7g((=S=DIZ<#QB6]<U#BO#E7@MO=J0&bNg@^EgXQQIaK7&WH>Jb?,Y/=BFf:=
f2M52@g_4ca>+YS+;IKb\3#=@&@Q;aaf8]]&\KgA5@b:;>3\SP9TXa(P+H[fPRaY
e3@C_N\9H5K3fWDLP+J(S5+41N>G@V/3#=DPf)f&+C>)7d4cGd5CD#^#AHcY(&7#
T9O-S6-JVTW02abNUSV9J4L0GNH[#Z.;^H]#XJc8)U4W1QF9QKM.;=?]G<.E4#ED
YB(DJ;ENI(]&]>[]IPJ>]S,(SGS]>IZIcO,_],0cY<Ug&4EA]LMVIA.>=^9N-?.J
TL9cV)/]EBaN7>@?,CA+FI..gS8[fF/+2541Ic;.cZZ+.EC]F6Z<UWN[]&QJfBaT
[eGKeB2M2;JK)e[IYQU?^HOgJMJCc)?4:3gZ7a#a^I]/Y8&=:)MQ>e&H>gW1@S/A
+S:aaC46<\C\GE(0?=daM97>a(O]YZDV_OSgW5g_K2ZGRPbEHX3TYT/RPRO,MF5&
(dXA/\\ERI_6YOG/>\10=/N317V,Z.=4LA#EH_8U9J&dGMF_,@<QBS5_W.;ZX>9I
GFE44;#XgD@KHS+g)@[S>e1f>K)d;fAI;Ag58WCMC=,^5aG\1V2N]IM(52.<8@DB
TfOU&)C)];=<3e=_aTfA4BKcaSWR3YZ^=FDeQ&b:AAf1AH]C=E\[4;Z@c#dRR_5M
\[GT4N+be>Y4G(2(?+dRO^CLTg1=[5VLa<5.B,U)3fP,JNEU#12[V^+e:]b.F&ML
0BWU78GDSeE[&gKK0+,1S:&&QT3Z=#@K+Cg@\+\5Y_H)XEe-AQdA]e_LZb68JV22
UPJP-S(Z^/>_Bfg^SQ:T@OW1_YM?/c/Z9e\?fQb21YELBe4&_>N707DcDI[CYeb<
e#7_.UKZIIWV-3F)3E_JCP=8[ZK\85Q&N^cJC8R;5QW>T;_P)BNIWG=5M7EF0<W?
;)-J9d&_?ccfD]1BTUb<EX.g;e.\K>-.<S28/V3K_OD(EW:Q.R]6T/0FG-@;9SU5
]FUER>ZK5-J>]TG+PN3#&6Sc-Y.0dK,&Td086Gc?dF8&Y2RSa[W(23J\R5:;\IC[
K6O;b=Oa#\g>(2+?5S2T478-^S#N4&8,7c=A^[TP(Y.XHK(FgfY8CeAS?8aP9T=;
4T+CAN62B(7DCO9Yc>B)V8TK7IY,B-@5c]K?<Aa,G[>IK/0DE>=0M/O9Dc4J-E)P
=1fE/[3]\TU;@cb6>G?@;]<>2=0VTCTK@V@[eA0IePH&0W+G-;QY>;^]g5\(R;0]
KD5&HDRY9-IRBYIQRLK4GV8RBD1c)FXb?+21KL>I:;ZdNO)/;-8EV9IUcTNSf#GR
C0O9/@MXdWI=62L]UY7K9F#O3X4^ZFY)Y^?^@]d)K1&E3@)=cV?L8G.Y99&1.BW#
eXV0W[MWCb8fSIa]7)50#KK<NaX:CB3bQKe^N5FOg(=^5R(E[9N&;;g(<WJ8XNgJ
aFac<Y3I_&;^,7F]/A)d?fIE=\<,R5=WZ7Z\DWB[TXR/.+WCWV)f:FEV#aTW0_Z]
PFdX-<,P(4Y7#dMI9M\Y(8O48<#-\(-7>FfBVd^P9PLR-#bLC+<1&F\O37eOa;2@
.E_ZeMd1-S(?c4(aR&.8A&MP5@RC/HGUG9R^2TI\X#&S6]fUL/JY&3V4A?VPe#[H
I8e5.LM[W.aE;4W/J.NQN,YJ?#LN/TSR[R+TU;+WJ_A3]W<=cNW[;LRN&N,7Lc2S
>FeAAeB:A,.RS(KaATI<^_@STbJ?ZDGg7&X8&U?DBZK#OXffD5L[a]?-Qc/4SH)E
TSC]?C<P(HeZg5];aXdALH=<TXIE;K?a;>>d&C4E=Q-.C=\+S:/-S&=P8U/IfM/0
T8L?d&J:0X2W2^.f>5bB0X/[I:BXb_>LgdVTJ=P+X=4FVg1N(:,a728GHY_R0FDJ
M;+_(.\0S@U7U2.K67P[fLC&BTda4ZcY,P=F@]8FND<9gP5UU35^a(K54:V:8L;D
HCN]eYT-=9b223:@F]_VK+R,W-#:J9R<D2=JP)@\_-(HSP2K=&Fe,.(91Rf&bLf9
+5JEQeeLReaKFAM+JP^QZ1KE1=2FC.KF\<,GBI&B]bJ/?UN3-)g@2I+f]GBaDTGT
T2HPM9Rb/[1\J.L;J6:Ie/c9Tg4[)L>Y/M3..Y_[EDO>Qd8bf#AODY)0gPQKZc.#
ESAe-Q+d0NObRGe[_7B#,9]dEf>JI<3GR5#aRDL)I+Z1#16_U]V8FD[@S7FN+GS0
ffLf2d?/=fJfeW59S<;C=;EV?aY=FTdV<aYH29KHU58);SRZGeH4OU1JXXXbceBF
5EUJ9IN-b4VU=\@18_[LDa2=<K3V6DCcb_LE(O7I.4BG<0d+VWg<PMKP+dH@CUZ?
,_HWQ/>H<?HHV\:+gT8TI5@53G&\0f-aVdge;SBa_GPgdgWPEJ5EIVVg?J4<WS7e
92S3Q<E_aG+=bWfG9YJ16WY-_A(?Z/AbbgI3VKCg@12YeL\,Sf8U9F8[WAeW)Z7e
7,9[/)FR1=[CEG7N#B(J(2[&EcO8(^+2>U=Dg\:&\^]gM;+&e:?UCTKWXOB59YG0
3c=X:#d8VVPPDU_/-BF6JO=POg4e;Pb2T1.FLAAL)Vg@]+OdHIE@L70PVA64_/&C
]Z>XZ/dFMYX#8]dXIb_C_/H]XT[JW(OGMG_ed-+,-Y\d2DdBQ#c\0;Q@0VMfI&P:
&@J&c\AEM0=5L&=-+L.KDABAODK2R;.K\[V4TTeER\]R((5fW#@-4Q+M,5]ad6R@
UAH=USA(01ZH&.AYV@-[H=N]U)LRS/MDU/KJRgZbP1-A26GHSL,0BZB=@9b2bXA>
+K7e]Tf7_>E^aU@J7#Z@d<.D:BbEE/ORE_+U9F#J2@S.F6e1UUb[[W@]acg9ScMS
[3RZ,8Xe91M\/7ZZcdVJA2=aVF_A&3YQ^7&aOd@<P0a)<_WV9Q(cbFP>INPf>&GE
TG2b>R,K7K_M>;9FN3UXT=\TCNC/gR0?CU_/8;I9<\FNBCET)4J:K3Y(E8Rc)(&6
cH132(6\_fH>;F..(OO-=I4QcMBTH6/]:2bQ;.AG9>,/K68WV-)-Pd#D1AJTS+>M
aT_.&8+Y,JgZLCfD_IUNOf-CR89d7BdL4DA@?-E]./35S\HTISD3[NdVI/F\_NR#
;HE[T8S?HH=/IF9g42]?(?=TCf79F#W/AdF/XaY>-B0,YdR#,(baO-SVAbE:T7+S
/\894P#)^;QP5Y#f;OK=\feB6;-=05aX#]F+VY5C^-Ib<TQ\Va3WQ4YSWEf6^>LZ
3Mb?&/UMNMBHePP,4@FS16O.C9\b5];-;\&c\M,U=/IV5DN3S[K1ZO,eW,&7U.MP
bW&#DVQZ#-N&6?I\.V3)2/eN[OGN]ZMAL6VIO<N-2,KEg\gK6=K[:eU&+25#FS-M
7>H]=,UdM<]_,=]PRP9^V#d5OdRAWBfZS<VT_QBQ1(;9K2ZJYP:AI(J;]?:MB@/0
^^XT7aVOQLRF(ga7[DBU+AY3>-@E;RT,AV.DA5]XCUJFSe2GF_MTIB)Qc5U=,PE1
VAU)CGNd@K;-H4S.H(3R;^RY6,Ug5<E6N?)U<33#a#D2=I]#b/++9YKW2aK6=ad-
3K?_c<3gTdJ#-=:Td(?.T3O,.g0JEX2_^87f?DNOZ_G9&gB))XM4d^K4#_T,.?V^
?@;NM6..P>54?e2]O@?62JCOa3??LC/#>3B96NgeQ2^=50[H;KbFKX60G4SW9>?^
2F8Z80fIJ5S5F/.9SDVAba5:aD9)<-7(R0S4\C=SSbf-PAY8;7):<[L67TDPOMZ?
(X^a+6JQeJ0UgE);g[NU_BX;e\LWZN#b3g2FUNMD/E._:S-7CC&9N+ZXEOT^=JS4
Hf3C]9/d<0WE[WL1&2H1C[YP\9H,Re5CJGY+<a5-3@F7@A\eSHI)2WF+J@S)HZS1
6Y[>]cFJ9OJPWUI&7)ZcZ9?E+a<?@BK(&3.#(/cLf-[<\MJf&cLT&M9MS>?a<+,[
d9@Y@2O_.E,F8d;P,28T9[TR6Yf1^H<WbMS\=L,DOUV/>3J8E.fP?ASG3><CPMQ-
X[cBK:gI8eGL-#aG\ReL4<,#[N]/&Y1T.@c30BG9O1JDS\WM+(D5AO1b/7(g#D3^
#P1=B@?bTMW)NC5LgC.bW]+.PYYH.1KU[cL]6.Zg/,HH92MT4TT07gQ9gN4;2SD7
UQJ_),:N&Z)X_/egPC<\3SI:)=Q>^81JdZ;+@c?DI;M1ADAN9f,5;-O5dg>98)gc
g&28V[XXW?Zaaf^X[E<M&UO/7+@T_AS+8N/]<c.IY_Y+&F2=QL?,OX>AJ^5/g2X+
>_c8b9[9[5YfZ2])0<0VWa0F00ITZBfL),VQK?+-GDQ+W2&#G+UZg[=HFWg@7MZ\
f?CJV]fe/AJ<LP_0(\O:7WgV#8KX=dZN;2PN6(T@T2@PC_]H;)&FUKF>MabD@8<R
abJ2&XZ3bX,Ff)):4ga3X-#3==Ue>W]5^U?RBYO3\O]VCFg;d;8PaR\+WQJY5M00
U1]KE/dK#;=N2W.@cBS>]ICL5gO_:,E:,g9N)a6DIE.4&a^/3<B?e:EEMPK&JMF&
7Bf0\Cc#Q>YP(=KPE@MA7\+L[#7:<Wg/c(]CB<576AB(^:R,LcEg].)P7Y[Q@T,.
SLV]#FU)^U,=e>NM81>Va,McKU^QQ0D&7YYS?;a,#IK-/-M(]^CL.Za_?+KIfY13
4(/V0>.FL;J9,QVQCJQ0M54Zd4Q#-bG91M&b7RTI8P1aDQ)_(\JFU)?KM(4FA1.[
#eGNGd>e&c&047HBd)W0)O4R9_KdNOKg70C3N6S:2,G03J;1AW+7g:^c950ANB(\
G-NPZ<cBb^U:ZFWLTf9YRB:aF)g9__c_P_]<N=?L.U:W/5>ATJ9)@a4:)NfC:26V
4d7/(aTJCdg3/[RP_bE+P72dS:6gKY=b[ID1YC4d@cO^Ob[@c6b?RPECL7f>\IbW
;/a.TXHVHF1-+]IU_<DPO<EZ3Q6_Ic+.Ma5^DDJ,5=JJ6[Z1-^:gSGO0+\E(cDM0
Dg:3_O,FGe1+W-9Z7ML49?_31WA\\:Kc;K8D[?L9Na2RNQXE]4CK:.]MROO^=g[e
]RITC9cZB+/:D#Q@D&f4UG=QEcP#D32^LE:@8c]MI@Z_2(CB&0JP@)YH;2>H91UR
5F7JM/^L>)VL&,gL:S71JbN_0&/KZKS5OA0^IGe,6C^-RCOO(4Wf9(E:dVD2T./^
)#3dE+M1LJfZ5/[P[[B7J/]:?.))\=3Ye(KfQT>c5;2:e/.8?1;_e+JUZ/G3fJHa
NbEA2EKIEg4fZgHVIDPIY\^@MQ(2.2^fP95Wb(W0_?[JSdb[]aa\KFb.;2:YAF:#
#\dF@@VMS>,XWO6)617S2[\3c@MX3,(XYLTCOe7&LDE3d.^DJ9Fg>&UG@e:-Q;DU
baT_fPaIR:002IJb7A./45<PQ:B#Ddf]:U0;)R@d)K&/K:EPDK\QS=B+P)>O5,8.
EbBb0V:V:-<[XIJ6NR@LTH;T<ULII=&FV\cVf:NEZ04Q)0K1@&U)?1;>\LTgD>3,
Va0+VM-02bAX&^8Wa&eLOEFaE5_c?(,M0L3IMf)@_W3<#9ecH2-M)++T,(^)R,&a
DD4Lf5bcGBIbeD:<R/@-\K[#[]9@)N#@N8NL:Z&OgKD-T0U[GNI+8LZUK=(@^?,8
<F[UadWdARf2P[HXe+0NN^,DRXHQ>X[-ZHLN[_a=RH>@D5ga^QbDf?/EF(H9]JP-
Yf<P3?OK:HO^f]K&@,G&&N^_7KKTIZI+J_]3VM[Ec\g)#PFeFb2Ge_DQYG#3(\cA
ECO83O1RC/UP;_=L2UYNG;dZ;#KgE?^RUL>gX].DT>,K9ZS]U:bMA(X;9eJRHA.P
D_1U+8+aLcdXLB=dE8?E_LcH.5(_5E+OT&@@]LBN3^bO#f6YOPM#D&fG.L;U>8[3
0Y[NBT9G2@,1/Bd#<e8&(:Q]PAP3Q_APF[VV:^^N9bL^XA(5NI4/bLHK7N(UT5V7
?=d?c\<\dR;>GIXbg9KLT3a<De#BeOXSW9]@8F=M2E4H[56K,^R^:@_HHVOQS5+[
H5;eW[H:][,aERZTNMYF(VbR-e0)PXbB/TYK^4_\,V\9VSUb3bBK:GMCSSRIYTAd
Y[bAgX))_]>8@4-L;TS.EG5<X)8,FCCS8M(33<BZ2c?9O8U5<IDg5Z)-#PDUDH>+
):D,H?2XFO1SVH=1L_JF7^^QdJR#_YT.R3V+f=FXPL@7APBZO-7OI16-7:&_CGGP
QFV=ITV;SJ2YRXCg;IN2@5.WMfK)eXVJO?9.#cEH]ddC4BOH-5E8^)3H([G\;P,(
;,SaOLg.>X8/S?;]Q3DX348XJH6R0D4\(;JM=DHAf??a9]UJ,b)P)EfX-aa.?;5T
:3>:_IX=d[Z[(KE+g>T@.2M->F(K0B<g_-NA?YfL.+K^^Z5<8<Dd7gL;:-R&NU_Z
.UR8L+<AUF0D7&J/I+fa[E32M/G+Y&:&/18L1EGXO-aF1A)3;X5a70?+T0^[JJRY
;W4#O>IbH?T5EYM=(S2LAKVYKbfG;M,NM[SO-6/g^e3,X1G3#&>JKZ?PV.KI@YZ6
cASNae[X#[]MNSM8QXY=D])Y.JUM-Hce6(DH]))X/c&=TeY0(A_XSM_&FZ-(>:TZ
HNdU21S]XMgQBCebNb<B[Fb8Y1H@M&S9(104:XNUBa0eREW3DU1a?2dO\[:/V^cd
4bEON:FKDZOMWP3J..S^Z_A5c,N&CMG8BG1;f_\^.),Og(Yf0>+TQ#OBQ)P,Ub+E
b+E5S&B3+XR\AbWD0D:aDD2P@g4e]IJTQG&dK,)K<26P@.7<7\FDe<N@UV80O9>X
-L2b8&UT6a:(C<.Za1Kb5fJ2O93ZFV:>Q1^J0CNWT;K7C4UUMT@OfMJF00QLTFJ4
XG+Ne,-Y3eM4TCV_TYR2(cRADBggA\GbDS-UI[)<gUT]ITVR3^L/7O]91>51KBT@
_JFfDV[dgK7/TR)Y#5>\?a8<dG,:5_AMFSF6QYLP/NW=F+#8\MHb:eEP59S/(KA:
QI5)LW+G2LZTLb0T=&W-?<d]I.J14QHATE;\GMa6)>Y11&M+5G4G45]C9:,/Zc8)
\Z?E3NF+1Y4.Fb0X/W=D:HT?C::Z@>R<<3[WQJ\TS]a?P_Cf7Ca5VO/X7c7.LZO?
/.bf-TVOaY2(R\)#I(;d&g;L\PO?U&MV9P8,3=N8<Ag?R:,<D)N7>J83SH7YS>JK
Oda<b.3O:dObY/:@-?_<\C;7W&R<>:\&38Ag\YeZEW9T@)M^74T@U)OUZ2:P=_<&
0TOg?-T9^H/U5e;9^J2]N1(C1.7b+AJ[G6DgYe>;^IH-Mc0gW;DNIBXPRWUdKSGM
b>CIC?&,O.[(NUG;(81N]SNC=Z9+bVGeAdO]1)c(KE.(OV4UQL]8.:^YP>GD_]@^
=\.HWOd^^H>[Q(@]F1]IbJ7U60X^8.\Q\b\a)_4N4cVJ\1XXUJ_EN6>V2@X6RINO
gbJ14TW]WXCDI-@e_a?QOGTOB6[.4.9)R5#fOFA?)IVKYY9H-f1Gc;\JB1N7@:e=
<(aM&W3dUN;S/C0efP8J;[:G/cM+Y8?^V.75Q,-UE[eabTVMPJ<H5E.CTd\=7QEA
=[(,?,LL]9172JMOTTBU2>R/?9&E_E<-:Mf;DM30bH9JCZ(cYXYW\OM#Lab?+be9
VK2380VRCUU5399]WE^CGWFK9.JASXK]7+9:Td,.[ZZVOc&M/&\@>Y#R>ScV..&.
7(E4D]YB+C39OJgITIJ,Z.U\bRb9LFc.UaSC>EN<@OOaQQ[Ce6IXcT9e/K7_F]&:
[+cE.#H\I+#)+;U6/1Q?B^\J@,#F-M2#7V^,V:J->9>N/42Z=N--7?W11?&\50Mf
@cLVNV#&1Z[X9276J0a7^Z2.012U[O=#/09V9R)[3R7FDPIVe17/PfUZ2DYDKQ,Z
<_S=7(Tf\)JFFDV3NcZ5>:,f#1=g+4GLJ17=X-R\S4_?aLfWMV],6JQ8dY:WTd(8
R;YbFbJFZJS5Q]K[b5:?&YG@RK6&3.+baK[FPU@M)@AFXW@f^^^WZ,[ZH#f]TDbS
,Ne(6E;K0G0dYP8+/Z[\GMLK(4/Vf4g&:JGZ(\(7-+b7?\d;@/PfRLd]b)_ENE:_
II6e;LbEY4Q2#Bee9#dEA1/c./OW?XU84]+cJW\:7&J0IT]SbAAaH\HAOd[[GbgF
GPV+]?<DeF7S[&feGKY0R@Ef]c6Y.5bO?S30PYD.7WGF;aJ?9g(>S=OFdL@H70Q9
?U0^AZeTAB\3-a^#60WKET4DR0g@&M4Z3>03]@=<EJ3>OKd)S)S#@8F038>_&2d2
;>E?JQ2/dSMUHU&e/(5I(Gb:>,c<,QSHUPN1XdCUM5^DaN/Uc1GZaB?K7_Mgg[]D
HPP?2cP3a(;IeWV9-)S:MP(J_LbcGMa-MS51SH[N3LB@<743S+,&25L?QN=Q5aU2
NaN-3EZ/8HSZM4?I#JS(0;HPL2ZD-UgU00;^@4PPZJ7-8b&eB^F\=F;^S_Ac@IEJ
SY7W_.48(V:V;)928aGE[X1IRKNQPK4SKRN0,R371&#,K.LS))S^=E++Y0@X751D
SDD#0-g.4H>;dLR+/BO)TZ7=?E8__]9C)<R\H.(Y/]MJ/Q)O+N1ULM-)bML+8MQ[
EHM&f>,=/:>c9OAGd_8KIX4LE,Iec)BL.@9=<dHS]4VdYgg1>N&R24>40J7B<6Z#
V4#A7@.?=)Qc1]Rdd>P?E6H-XHEdK]6f&]a14[P.VIS1EB6ZGJ9@O^.CVebP\_D-
>Q6IZR9&&Sc)]\6MW:gW\gQLIe>ET#1eb<H);)204:T(d#HOF-Xf],:A+P+3)-?D
;gZa&EP]+2^JIQV<=FAQ(#OW(<=0M4Y:_<QZ\Ae<<C)@E/[D]:ZC^@]K,6R-YbIQ
9c\B[1QZHUS@(Dg2Ve=[^6\M0&PV6dFPNLe]U9BZ;b)L3f<0RORSgefA/H;F)N6+
OP.8(76fDQ[62UPBb]bG)GbeRXb-6^=Meg4G1<9K7\R+TUD(dd1<DB_dU/6WCg9T
^?&YQM4B[Ae#Ie[DXMR5YAQ&ZC2=-YHfW.P,5f=U;3_O3B(bN.SFUE97c:b#3Wc2
HRAU16WV&\-N5)<JQaB2WT;/+d\R,/-9A>:3WT02798Q^WgOT0\a1+D2PQ(.)?ED
PU]R,O0FRG@aC;I1(]-:DfPGDX8KPL?URI/Q&(U_72I?^@]D)WbRRgU2T/fR.AB@
FZ-D/4RS/IZ/2?2gG1EG^?\\gE6_T.RC,#5T(fOI=d<0.]([-?62a6C9Hb)#_-,L
OIS]AaC\9M+6ITXc-c#0KI-33fUSbH7F4ZUO=0G@UL#SY9O:)M)H7:V51-WL1KQP
1CI>Zb,ZR1,fd3O>6A,TJ7)P(N?GI6--XF=J,<R&2D>0EQS:N)[+M<P5P_=&E=4c
G3F)B/OSGIT_A@\4FT>7Pa@^Eb?dD-^V#S4;^e+7/[L4<(5ZgaSK[dfcRTN&XEHF
GR@&/RP\P6A^VH0Ya[=Igb1F&8\QI-f6+@X(#A<L.2-X6Mc4]3/\HD\ES42(.[?]
9ea&12/1^B,6)[?bDW26gf3dAcb7bG8G+R8<BI0-SRb)=+-4]42/H@+[J(MP3cE@
\PWU8Y=aTNXd@]Q_:7O_9RK^FS1>d.<U6f9df8I^7NR8#^J[0f^-=IX?\a\MIV^g
D:2bI#e]A?D4H(OfH:fNeNga;aX[7W(JVg]E2R<0TPYXVa@HJ+:3GY0G<:.YbfT+
1DN+H<+5cK>37S2-+f^SC.ARDDUT&4;HMe.D0[]F/L20gO&)/Z=H(e33=+->EIP-
PIB[HcE(A;[Y#8U;OBYQZPF+VF@aTT&Q13@&U.4UR6aIG04+Bce#;&9J5Tc\C-I0
#:.e7B>FKQY#:ME-ZbI0.0ScBH_UXVDT.RM07/DJ3W>Wae3YATJVEU,_G@02Y^C?
AaJ9Y90Xc1)A/KL.<]IAK?8EeBNdSg^];6Q^WGC+:-eZMXS?0e(^b;TOJeZWYS8<
7ZQ84+Lc7a&=CW_(EK9<LK?Q3Qa9T+2b_?[[79E@E9W2L;;4bQKR9L=/JaTL1\2F
^2e5^,38U\2:=GfQ<M>1Zb,Z4FA.A6#7<O0&<J::&2:.\.W>Ld0STESXd_8>7QK4
29:G_9?6BUg3>O32SL+AXbE+#H/&#X3YB;3&?=9gK8H.XL/:0I97#@W/@+DI^-]/
UMIV16MQE]E5bXDUZ[=OS),(I22Bc1d27PT-dC-OO;fB8cX8]Q1-+5MG2b)\H@e\
FBHGgNIbY-_R?/S8KIGfa+=_NHE9=f1I949GUdf70:;=W4\O8K4)D1?N]EJeMcVR
WFgcHOPRG68B<B3/G2SOE1?cRD>KXI2+P@cS,TXAOU1+<UaYRG2R0cQ[E(>[NJAK
^23YLB_L1eDRUMY:0SYXDT&ZWeB7d+9)f0H+L)-F>\[VOP3^GYd8T)^4L]]JYMU)
70U]@2Vca/[_PYLC]5Q(:bbO;;6]=.g^AAA-Uf-A3efg\,dgJ\fef8KHW<IF;^9Y
,DU7IZS\G]>O#.>-M-3X&D4&P-&=.JHUUgTEe0AD<8/AY<I:ZV0]fV+>H&))VKMU
W<1EEX>\Vf2SF._ae[dFHDM]++O9]@WD_/TM36]J0eRY[de4H#-S#X[.)4#W06;c
C:,;MGEJ)?TL263.>@fZfcf7UcX;2RFS<XHAgf.1:\O&/#-XQdHVBB84W51VUaF?
8EZDgc.Va;-TIYR7PLP]QA#WaOT(GU(N)e&/D5\a#76YHU3KR<:=2N99gCNe/CbY
4g1TT.(+RaUCC#8KSQ&NGV1,fTM1DT]2IY_cc\.R^YMKTH4_3S.Q=ag)3#PGXZ7W
NaJW6g&c+^]&M#L=C;dA,_L(=?(L9.3RQ21Q472gJMRF<+ZY?aKN;7R04.b;Acb9
1Hc9U=?0gBC37M>2GKC^44V_7O@SS4d&EMFK)M#Q4c+(U29/L0]W/J<P&H)KAc;^
^O,L1N557fZGfAP0URGA/RV__dLI7)ZBH[JOY.&FJEQ0/;68-g2MK5C@e^8<_X34
<5U1/g];[#5/#3ME34[0)6KL6CYQ>JSTC,U)dcXFGCDfR6<,cRMG_K+0;)O]#VA=
7?^f44bU9H2KVTd.IWZ<YI#<:IPRI@]X=N#X#&Q>/AJKG\fIMA<-7BV\+9MLG,[_
UT@O>+BW@#&Fb0N]QAEb-b6c<Z/?-_4TeIQQF#F&PDZ<^.8a>UD&#AT892<0N/8E
Uf7C6d:DK2f,Qb/7PN]IeV2>MJY_BZFPEZ8W+AedWBD[R#<?:\QAQ]5>@,Pc]#(,
U6Z3:-DRPDe[LdJ(c(#@aM>M:,),N+2Cb/e\QKDcH:;?da9.;KHOAWPc[/7bc4[T
>0(eIJbE2?W.gJ=@2cXMIU2NDH6.+D?(;O4>D++UdB][8]Wc\[UZGK@eaF^G@-QQ
.OY-G?Y3K2Z8V\.5Q?MSGBMdNDJ,?)eLK&gM>OFY&Ua.gC?:7(WWYEK]]P+g7F:C
g05+3MEP4SH,#9LA4B4,<3dVJ0KgMG5E:>a7,aL_U79+NUFMLJfL@=FX^]N[6I7g
&H:ILGUNf&2:X(P-SSgFP/g1#ZXPL[2gNSK:L6.,T7+M.-BWbDSLYDFBRg3LU1O2
&e4HcNW9].#J6W8\RO?g<U+[8@@0c#R9bW6(1C]=7FHBH;C#>FNHKDbWY\P;?WfZ
;F(&1@Pe/MABJ-@4O>736W^a=N1_O7Z6a=^)2E&PaYSb,6J>T5;+&;M#OH?dJ+K:
:AgUF71O;XOdY=W]26:00>d@V^K_4)P4;7/##fe:2^09dDgc>L9g^Qb<J&/b_ad5
;JSDb_adaL:feT./;K]6ZR)H3I=>_ADNMX<]]MYZ8FRe@L7EV<?P6IBF#PSe_6K6
cG^F)P,B1W)L\SV:H6752\fS:3DM?7O0&=2AN7\J+,aZe>A^=3#?O_Jd.c3dR#P,
[=6\85+<@Zc(Q\L)Md[TR.8dFAHH(Nd@C?:aNFE4[0>?YNbf#a][6;8UYdBL\Abg
#Y\(=6ZX:>DaR&:BM7c:cC[JNBNBBaIeSO2b-[KR@ZI3X0\RQ\cbGAecXN6VS7?\
RRAT=20dT>N[c5EL16.1<(J^/SH7SS+H9^<aS)^KHLVa^\[^<?b,,[]cLb74K-d@
]8ag&_M./U[[=(bC..e89dBBN>6g^;e.H_T4=Oa&9,B)cYObdg#VA//1[^B=1-E>
72TFWbY6.J6(BH?-,=ZU^T)>VOES&?E0T>JVdN63de^48O:E^A9H/:-XR/./CW1P
g5]Y@X2].Y->C7\+b,IVC.MP69?)V^>]UCX/GHMLagU#BO)A[X<)b+H6/QOSg:[X
)DPeXG4BT\8,,CM?IZTQI^2Y898=S17<:6BQO)g3:5>Y];DWc?3Z7Y>U)SA\b.]J
a)eH442I80bY7Bb@=F07=M5W14=.Z9^eV-C=@NVac0gO.:AWF84B8LIG:N8V3YXT
)I_GR;f7KYfTG]@NMLd:9B5(ZB-K)BH#\CJ^Q9QgAO]#/#Ec1@?RcJ6U@Q6:J3b\
2AIdZ5Q8-_P.G26(\A^FBbRQ?-HKNBVI7=c6U>^:G&Gg->DP[9D60J]^;XF@#;B[
6&0Ga)Md0.+Y=#V<L&J1\2BaJ.LU7<[2YSWH>GM;@&C+;ZZeFX8:HK\BW@;XNdX4
d1IX;?2>0&E4FIN,OV+[?NUSNS]0aV&CGP?Lb>4GH^?fd9F(LW,(FN(O:HV_GfHI
.EWMI]=&1gO8T-K2TE;W0G-PL^&C[)a#XgV>YDR8YD=7QCb-.b/8Cg#RcfUe,c_B
8<JbD+I&bM/OfN,8D[?Yc;#M4E6+J2HXdD_e6Bf.GO22^.\\@0@7:a#e8aL9HQJd
.O37L3B>-]fO:4>:EU38ACJ:6c8Rf5036+aNG&aC:JU(<WI?ZW@(F>XULf]2TeV4
F01S:3^dR&?_,8^)AaS[S?&)IU(E&3]N(a&7L<WC]RUYI8E;0RL4>S^B+-dL=7X.
^1H&IX;#1)-CPN)M0)Y<aR3df)<JM38;#4]+<\KQ)W=^F^C]:@S;54R=?)EZPK^D
<V:XWa84PFAR2c?7X6D>eI<HLH_7eH\CM#K^30SH[P(K1JFgV9U,F5W0T@@9+>[W
gBWOFO4g;QAbU-/#8;6\>fWDKI?2@e29O9#412eIR26=dDf:H(4&[,L_RY3<Z)^1
)ZY84CJbYQUb^DBa[MKK+a7.]#J8OV.7LW-#\;ge1a<0;Q,F/E[ac9>KSHT86#JI
=VNX?L,d_e\AMA,5<WYWeSba<:<e-7U9MO#8&5-dRa;SfI#DDLDEV]NGJ^^5V+5?
D7XB<c1)5(?FH5\?7;f4JDF+^1DXEgDDIBI^c:-c6=L6S@\8^f.TfgN@?a(:,Sd1
.7_(0?-AUY65:CHVFZ#RSfVPR[16R@@@G4EYbffPP(#H+OIM\Z9a:,QgX,IDTbAY
PBd>dW8;&TZVT/UAG&.aDNGf=21+06J]_1OV1gb-Kb2,69J_QA?S\S]5\(XP-V8G
,\14W3Pc/18,76JU.Ya(PQIWe.3YEd0e_J;9#0Iga1aV92DG9\\VbA?4&=-c)HfR
=ROb@,YJ8QH=5NWQM=adCW651U\b76f,9,(FTLT37?NED>g3XM_&X?@7ED\#^DXf
RNa,eWR(U1-W:D,O1&Pg&>2Z+3]Wb4;06Rg]A.;c\>D?J6BL@URf(W.1+\Ub+@=;
<XRW+f&TO<DC(F607eW<^_11bKKH^a#D_##-P7E^T/]->a<L>QF2a5Q)aX1866V&
X-d)/\1b:@A[0A0^\>NPW8XDfX_N1g87<aD(^TELF;\dW)ECI>VV/Z#E+/cF[_M:
7;AOH?1&(LA:>ZQ\1aVW7C\2c,^;V.>^TE/fYeFUa864bR)#/?W8-B9PNL94><\f
()BD0cd;Z#2(a@]V?9L]V/&0gIHVOV);Ae_gLB>3dN^:5=T)30FX94_5JfaP&MEW
c?^#DScB-[#SAT^^=7AAD-R3bVN:HQD(N:-?B,@=KK@aBU&XZ?.@E]S]9D>21]HD
&3XTGI\3O2X]_H<-Q;-+)\U491M6^1^#JS#OH2U2D1cZ_;W13L&g9#7/&Bb#MD\N
D5AYgc[X-_Z;F#,4cGHPFgBag@eRbC+NgM<BT9)9FBVZM5CAMAE#NWe:C;L(@XTH
MD7E2(K)FAgZ/)]-H?NB)g3O>2@Ae)>,(FRMJ(=Q@MaKF;AY+-5XWfB&2E@\a6OK
T\Q^>IS8;R;Sd854\B6NY#H;c[0FR,<=[=[g4f4FE1d2U^LY&AP&+MPb:M_O08Ka
_12=Af]S.8W_YG+C0WC6ONNe^8G&bL^WJ>g=)20T?N#&bBX@JQ_EJ5JRQ5W/?IUc
0>W9,:P/IJR]=J:Rde6VB_B+RbF)a\A9VJ7A<OS/NW,VM+CU\NFeNR,G>&D,L(]C
?<e2RTEY?8T2U767PZTUN[_R=)cML:F0NOU0aAC5GeT);KV[,Y\OJMJY1]WOAF)8
g#E^6DcGH3QJX1cG6\bL4UQ,/[DE2S[6<:S&6<[7fX_Ua5J_&6Zg3g=g4W0#7b=F
JQ(9CQNRY(/LbE?F)T^<2V/.Z(E4TU,>8bPGdcKefLRW/K:LeY_;PXa(7,F)JCTO
9[PUWGYeSDAO_VZ[8@M&?B2/1cEPT:#CSDC)CS?+Lg+&QF5SNb592,UP=a^R90#=
0)4VTY?:@M1c2)d/V,YFW\68febH@)&J:9TL2A]YDJ7A<1>+UDGZPQ1J:/cE-^.)
Z0-YXF<Wba9,V+#7deM)UgFcbTN+/gf+cY2S)=aI#1eH_U_,4=S2.-I?d9[DcNQL
efK]/RI^,GaKf6OTU\7CXbaJa^R19XCfIGVVX.8f/#:#g-;_J9(#<CeFAaC(D?_N
46APf)@Y:P(4S67bW77])&/EU.M(Y[d[L_f4Yb_7XM:7_5K<VYVT:&7=dF<4gMDb
.=HS:\N6<#a[Y@dC7a)<KaZPAHePQ+JHT4=\dQ<a;]-A:FU.RIA)QBA\_BH>\K5/
T6]59V+MC#e\OUZL-[:dcb);NDUaK3ND)W:=Y#P,Y>_5>3E]2^<]B9cFN(LLdJ[\
ZbLc6f#X#PfQ1^9/=&KDA69ceV)PgZe-#[,,gMN@,6]=\03X=ZGCNZKN_eDCFf(Q
(QaQ]P\8_<B(b#g=P2BR91?WJWQ7IQ6gg&:[HdMLKPPN?/g1Qe:#+ORcX1G;]0,5
9OAQU[a7K<TbE0^+,3H/CJ[@)RdbW;QObcN\6<TT:bRUW:Y5eeRQI?QL[-6(NO0R
fBLY:09B.7Z5#FBeO=L1A.SFaB<FL[cCHBS:Ye9b0_1M+,CSJ^<AEKE.a@R1_X<W
BZBW1&g>X]6486g)[_b]1:ON2C2/H^A.<Q@_gfeS.+-+):NE4?A<9TcNHL&Y,]f+
SPYLF5:^C=O2c9c+aJ89V>R0\;(=(8,ZbV#YP036dbc:\U0@HZVT(20b8dK4#AgO
Pc#Z(Z1))&_G3=P]f-.+7cR,LOFc1A>T@@P#4+RYT>-0WgAcH2#KL[8BJ\6fR8Q=
A;)9#B02A4#0P,a\.[7H=?bVbFM6V=Y<ge5:BPdEMVb(S5&HcgFJ7)D=/UIK3318
<A/g8dgFY@3)P[?+3<0@6Yc-fb;/)-^8+eQ=&YPU5U;RP@.+ccN&8FRQTcQ\^S,<
e.^0OZ[?XOKJSg3MHQR2P>V@e2DAJDU4M+f&-&SKO(^04U&P[B/8[3b_L<RU)@)#
XfTZ0SXZM+H?e1I>3/IfaF6>0FL1S.;LX;7F5((48d4_AZOc32#365#_QE+.Id)X
E)V\F(dWD[PO@ZGR8).];01>Q/#MVNNc](1dL.Z:,X_\+1#SWO3SeCC42::-OB@D
\/R]c8A)ZD:;L:SMSe,@Rd_OQ13?&AcPELVNABY)NLQDTC7XTU]_N][CP>T@_,=.
4>48#D8b=M<EH&<e>3e0]4>>aAX81]9\4a]8T1#f>Y#?F>A>KDZO;_<V/:BHGXd\
Z@U8BIYe_0[Q9_]]e;f;feTT3Z>;5JK3UIG7DN&=XPdDg^af[f2f16gDTZ#I=<eF
TU-aP6gKR2\cV>5C56PQgC)aXdHDDGWRX3c3QKWZ<L]@TRPLOR.5<]00?Zf[<e2#
1SWB+M&B8Q4DVd-NL119&?F/VT=(e:ZZG[LXM3b45a54)K2X,?[FXBXDbVF=N5Y+
GaA3.XLYCMEYBT3ZJcE^UL(MbaR073<c3B=6YgW4RSBPT<6)&aYCY(Ha#d3SS@<T
QJffcIbCVERUDEXX&g2N@RH79H2\a#)N=KKK5A)),;J5TaN16]fEc:aT[<5SL81c
[F,BG;;>CN<d9YG(Fae,P:K#,F&XTT;e035CNcU41I=gg4]&Z[NKJ\Ba-MdCYK;0
gV\[.5INegf/\A30)PCMFZ69U>#d6@8D=Y<#/6a2T#<SR=[(@2ZMRWEYSIRZXFB<
Fc(dc.EH-NA?88)4IcWU@dDN#56Pb[[A>0.#5A0MOag)f3NAJ26AbLI:d)E?P]TS
/JF>Wg9_aW]W3GJfCNc8U49ad6NV./N4.-/>OGbAa=Q^V@AKD89HfVg425#LbgV.
F68#T(A:WJ?.7=Z3UeC&5^JKBb<Q>GHO(GS\X)<bbfg9A-;W]L3d8EEH(BI-5^5_
+G=RCL]W:UaU1JSU=8HZc\M8>C(4@Z=/d)(>[ESa[5G.I@gW&5Y8fLKXWST281]U
;O@GWUIDb\44[CO\5bO7QCd\;B?,/;<>aX3#)92HZR8:[/d,72=3[H[TQJZ8RLGN
3PEK[-WdF=\X<YYIcC8EfK[DVR^OVP;_@Y=Q.Cf1^]@B_C9UgU?fUS:JW-#B+BI)
?4M6G\Q(4P0FRR5X=?R3_45E25Pe)3+ENBWB&?)(-2CXZJ>S4bOJ--\_TE+]2(XP
=JK+Gg4772P^cHNL;/L5P9e71JaO?(Y@I(Fa08\&LTM+Yab=?&PYf[ES.WT[5U]A
M7c8:H.ddNI\O0QCF9#CJU,FP^+8OOJ28dN:\^(_53)[4JBGbSa)H_W6T8gaEU:V
4>?SeQ77W:J<Y#KD7L^cC3Cca0@;\82MU15f0<c4bV&LNLc;[aY\L9=B[9[KHOY/
L1a::&_JLQKb,)FU9G8^O]3G?)gI_3;eMgaSQ2G88-BC]@DQ=LFZU(a93/J&2Z:B
HL@.>9b53fD\[6=33(>M+-H05^fVg-P,Og8,=@+BQ<a+/_(S[(?8BV:;Q\\4S61M
a-cB7.RTJPd/4;ADFeM1cR+AU)CT(GV@b&H:6\;I4A/UDL5<bUHgS?5)ZK6M\LQ0
d4:X0c:3RN4KFWOGIbD&5&>9[2YP;1D=&RF:d8?Na>^=1@@Z+bJ:7e=64Sg[1DIf
gT&;0RBVR:=5&Oc5VK>IJ:f>c&-(R/0YU^2C,f_dD:MGCK4S_BeQ;ZRJfA@?Y<[M
+RU<(G7X[f5R&DF\8M4e#)=<):@,\Xd8.S[MX+H5OJ(3U4Jd.=6d:+N(g@0bF=A0
@7?K/TR(EcN3U,LIZb85YN>4@RfaC/N]<1L-_7-fa;g\)G(QM-f?5.NOH1TdHZE\
^7d_ZEgO0DHKIW?76Q9CT-B9cOFJSK;7/Se,#8+F40d&7TTO8S6d=Y/-4T89Y&7U
;K+gN95+4ZT/?\cdN#(/SIY50&gX-77[Ma<b+4VM\a40QCCCT&QBcJI[e.FI?.H;
SB@6L36R[O]&XPP.a3#OC#ASHO1>g42d_)fdNfZ-_^Q50FO:#5FeKLegQ,S&W&;P
]II_USSHJ7:7GbRbQ[6T=>ae/1^]._dK+0US&Yc+\M6[QZ)bFC2R?)RFD3Q+>L30
L)AP>9?Ia+b@QLX8:]N;)C=I&S&BJ5ETB/8g/SL;,MMcYO)]YU?4NI,]9GATc30J
Z:R/+,aQ#gff,6)S>-2?#C<#CDURQ.KM4/MZ12gUQ]CW,<OBU.bRZ9?<&N5P/P82
f2(^/-FE50#9D,QP1O@)3OI?b9b>@=G,N7g5YPMB)U1Z<:efC9X+U6Gd]O<QNZAV
cTW:8_S1,NaA81--MMRKJa(Z9.M#R;#CX3Bb47f]=08S<O=88.c(Q6^>#)55c5;:
9:MF)?.;6M;B1,4?WP(dYV.Q7</#aOGBNIK?R3EOSEO<7VH(@SH?0LgVb7SJd-P4
XLIGWO4JaS-A\-a/Y#.?WK3HBFUTK;)fg#2J;A;[D+OKU5KN,I+\5O#L46:/77Ob
O(KV^8>.Z[VFVg>_H?JI/DV?4a7g+7Y@efH&fY660A>U,R\SI32[M\/4cQU:C.>I
8D7=1T/0YYKNaJY#2CgS5V)d,=[Q&J<,+-SXWgNQVfQF3AcdegfHX=;^LZ8.=#1g
@ZPHEBH1@LHL@CZU\[>WM>+JHD:WOPJC@4c4MWK6X<g@MQZfM?^V/ZY\IgXd@W0#
VFDb=Fc4;OP3SMd@R_IGNT23RZW<#c++8\O:9#^_&]2R0fXJVL4<<?a^I12IFOE<
4Y>0AU)Z0(?eEC160AD=-M2U#39e;X^Z,27;ZP]E8[D.>bF=?(SW^6N=V7S,4G88
IVJ)B6/<P#PP]#1?M4WX)J(52<PRfKd1:#NK]f:P9L)C0,&VT@fN)c9WS68P<G-<
Z^ddX5EJ+--G(94FJ+_A)<dIE0_FcL\<6^<F.1WR_AVU(<8+A3/Y5:33><8J^S#K
XIK&>JH+ZQRN<X.B[F:T2N-?3@T5N>UY+0IA,SD0+U&;TQedA=)11-]5B/E4>?R>
R]UCA5)S>XGaa_BJc_W]RT[18IeIa-P7)GX0+#C@SC0.PIg#,343>GZW2S2DJX8@
U_VL7;WBSb6QYM]_Z6.ZP^+_,M&KEFK(:W)^=[SOF_(3.(Ua>43E;Z)U]a+:bR,U
]b4/:b<HV?HMBJXP8fNF#JD_;XN5-^f,P0EfT>@VD@G.[YEZ5_#&[bZDJ.Jg?Z+U
^NGYU=dcT7FR@-f=?_@T_^e_#]\geYK-L=<J#:Y\\D=2-bFOYLW6GDG;#(0ZL]&<
)TT:M-[OSR)3V,.R[?^[L3]#@L#c,Pa^7LS/,-]BgUX,WO<aR_bIS_VD@Oa6DM2N
a0;0MX^:1SdUF5dXE?T:1P=.3NE9+7<f^VNZ>6&@309gU#4CJC??_FOe[F>gNdN9
7-C8c,QT@LS1T]#[&1(He.MR,(KD(])/YfKF43e08G7]^\[T9Q0VXLFHCX(6/J\_
dAWc7c><D,J+&_Uf>-#WQYJ9e4d-4#2.gP[_G1/beT6L=D1A4&MBU?Nf]6>/_X<4
,]&M86U<@4PMNJO,B>H2?G>\P6-D0Z9PeFF98EQ]g#Y;Y^YC^R=_C+ea=#ZBI>N-
4DW,7P^a769;&A3;@(0&W<dPgeKU?bR3K35[<DL1e59-)GLa5VaRD>;1aSXRBUNP
IcOLF:@[A13<Q(4U,#3d_SEK=&E-RGHEVM@I81=0egKH1H#<=a8GVD_+C-Y<TZW\
E=c=&P#\[(U&ZCB;JGC#GJSPLE.Bd.[ZX+>I/<5F6(TUZ;?Dbf783]0KR07#.V2d
J^X/PBU7@)<2Z?N3AA^d?Qb08+\Q:PA5H5U#:c-08GUGdS>[P@\D04&f4/PLYM3\
OZ3gc)A^fI=_=g7eTgVZZ)E1N?+WTZY:?&@COM/Lc8&<F7f4b5^1X79c)X=)7/-b
Eb6@RS5JUCU7V9<FYKE^(ZRBMNd9cI3>YZ=-N8&2NQ5&a6D-V0IJ>5B\FMN18Lb=
56P#bIgZM=,?eKY_9Dc#HY1)9,FR^CX9CMX3[M-6X;YPL.=-K??@Q;J##2TgcfG,
3L;C#,N.-F36NP8C;_\]+F-=_J3:Z4H)NVY_D@CI15/F?N2;=?+M+Y@68=LQQ3Cd
f9:2J/4C2+O.XE#c\\fOaFHTI<47gTF.7bI=Ab0SM88g751)M0Kb;T=WXZ_ELNaB
=gAdHb=-QIM@44,EYHe3S+06LBA4g(0,ZP9+;c5MOC6b^]&B[G]NQ]/W)1)^:E?L
71<^MC:e:E<[JI)595B40L&DS+ZQ1>IWE>c++Q4?3(cZ&bU/)ES(Ne8<0#C,?QUT
FTY^A0FLI1NAY=C92NCX_a;H?5Vg/_;dETDaG.(==G300214@YF2U=5.07e6e(0>
A6J1<52A@=Dc/ZCNAT]fI/M:=&9?7VP#ANAgLEdH7FGE+FIHAJ8Y8g1;1cC>0f[8
M_=Z5d#EQ@4#93MFU4PRP&^=,[Z:<\J[><AM_JUZ.fN\D@b^BJAd+bPRQb,#BC;B
7-V&,;KU3ba>25.168\M,KXTJcVf&IN/;(TXB=@CI_JWd9<6^V<]X/_(5^_Q3AHA
I,+ZcKDU:cM/_]NFBO+,0&B.1I^0IN,(5,eR>DP=A1?@FPZ08dD4\b@eHe6WY:P#
bF&T1B9@G;NFT]b;\_W/3_eID_Q<,-]UX+UQ>YM7#HPSKXQ:19K3:b5C9O97ZVI]
2d3,gefE,<=/12?#<#]7^S>Ag_X2/<6ca3Wb<>O=P-CbDP(G==Wf&f20BV&>069W
Te21[N(E#&8>.E]Q5_#E7B,F<L4c75Z__T#\NUdXcbM(=UPaYd<-3Z38;?#cU8:G
(D-=Q]#cZedAQZVAdgB=gWH<(?X2PX@J8L-6),&>WdWeY/-;OJNbgY-;2-C&_]]B
<WNWFY27SJ^B-?>OHADU)OIQOK43;,UAU_MA]#=?V^[.:)K@E(#D8C<Q4IKXE-f]
<H\[>?^LC6J(_<VRdECB59:6P#g=PXTZTcI1UAWe70REX.I:HAQQA1F]F+YdAVJZ
G[H63V;(]H_NB]0YaIXB/S[.KSM3fLdTCK]ZH(f[(R&6:Y@E(I>YI2LgAC25_=g/
)I^Z>V+:ON:d>J1^2Y9G?=].M7S.F),+&1W0ee:8R#=IWZBbALWFL?6U?\G>WZUT
<HWd0g)G[5]P5ZN=]?35c+M0PdJ+MAb7DB)MCXTNBX1^@+P5>\aaC>Tb5fU<_R\>
I?IUd20bV^JB+_:HHX#a4fW0=KJPA=B6HBe=D#JAYBR7M]P^g@>CaR@X^&S/1C=/
9#LML#:\D-7/+N>&#Pb[NY#+Y:\FK-FWP3]c98SX=cWSQe]V:NENGf9-LD]&C#;,
O4aD9#eC/Y<]P.&NNc?abIc(L4GZ(PA;3;LM^/SI+9P=WaaJPGDgR&T7J#e^UgQT
ePUdIFg&6GR[\G2g7:/>+O,fY&eU,g2gON8-J;GJ,a\D&^.gM<dFe6@Og0C1R]UT
<P,TIS:-_N3L,:?Pb)+(@g(M6]b@SRQ;&136_.,aE21#TQGMaM/J[1B+2>O=A5;K
)02AO:VD:UXV#G&O,=_=f\&,LL)Z/FC7K\HT[cMMTEHS\H7dV7B)/5)GOMe5Q5:,
Q#BEEb^)8(ZY8N3V-]3B]BS>2(ZSWdQd/a,X\@9C,F#@M;NbM/E\,R;;3(:#P(19
3P;TAOgHCdM9XT8ZEeM^CX:;630MI^dLcJ-(MF&L)1BaZTM[^VV+95S0cSMKc3dY
.D5dVO\1bRP6CX^g](\K5(G[eB&\7F1)LNOX4LG#SGc16UKW1/2;JW)9)DE,@[^]
IERM-HGf0LMR(fHbE\0O/;6aDCZ,5=1+YZc8X@>cc&6\(Q1Na:W;2Q,QY.+]g];>
7e>.#cS6NHaIg9a3R,5(<&_^:KQ3ZI<ACEY-O,IggPLF]Vf^AITDXL^6S9XSK?_2
-XC[1<bV^g&NV4LM099QH-54Mb.T@AP:\(3MYWa,G4:VTB+XB]=bL1=)A#)@1fZS
gCSUC_@+,]B;TPG>#&<?^(^U(=LR+^(P2Y8P33>6M@\&R52f_0.DKT&Q2Nb.#48)
d27CPP41I5/3H=/ZXJ#eIbZYDN.CNb99D#86.4H:W/>HX(R</MM+1bW2,[^@cDMZ
.@d>G]dW;7AW.OPAM36bJV:dLFd0@)IUA9,F0g>0Gbc@SG&\SXB>)7&\^caV1@FH
_IYU6Gd5>&/aBccK_<)DbLdc=QVAa?V9]-&LdCRX?Z.3?QEC^YY8DBO1,G7eW71?
^9/,?N-35TMN:JS^RJ5a(=[EWO0d(R\0J50-WRbABe&_Jb8UPbV7^PKReB-c<DE:
&^V-Q6c+,(05B3.T>Wa.Bf3e8,EfH-<^UC3V@Gd)CP29#X8:>NJP8H9E40e<9.3F
.@LGO[f(:^B,8CQ<W)S@2SOA5S6fXFAE5/#=;A3GY)GgQTSZIScLP\M4UJDL(4E7
_(X9aP)U^N#DQb+&LIE31/8VCP&YfG4UI#:KBKYb0QdVOcI(H6Q+N[K<QVQS^QUM
OKgVI/Eb:_S_O@dZ/MQTS058_<@>1gQSN]&+AZHg,OBO+-2/+^^\aXMb]]U^<a8;
]CU66N?^1Xe]^I\T+HM=Z0FH:E_IL6b_SA+d;/((Y0XJPE5VP0W=4+L9O2e&fHB>
;e:[M;P7@gc#_.MQ-fOdNQ,[[U>_&@8@A,)C]4-:Ge_3UbQG[4)a=2b?&FK@HG[Y
FR>KEg7H-,C.HQGI5VZ+YEdJ4@JZ7f5/7USO-6C_\@a<&:_4IV@e:0UcI1+#4:]:
:NDQD<0E#0B0dRWO18TO?S5@R7RORP3@J)3K7(7\,#?dYeUZH5@Xc2Q(;d>S?2\X
6c)SG[9&Z2D7E):SN^@<Q@AC5_=214LW/03L2(2DCD<MGP6Ia0OOS.]M0&HM;V&P
VQb>39:=5OeeH;QQMQCP^Jd]Z=2V&e.U+dC;S1FFY/U5-4dL#YT,^JVJI=Bc9bHF
6.XWH:X5EI4L]11X8+B2/GG)7)+)S_gPGHbfQPKJbUBZ<9U<&GSSL=>OG3980B_:
^G2X(4bP3<_)U8)MT0))[E&NHBSSU3](\N@RL.bB@;7B;5P+?RB1?d-UD2Fd#DZ+
Ta->2eXSW>7;Q4AG/Z9db98#IU@]?cIf^a_X^GY3U+<[]LA5+d?,U,#b74TN4U)I
H/V;beFLZ#Q]]U./+7GTOUS7T0.ID(<)#G0@6\0UC&;7L2Od_\+T247ME6eJEIC>
)(,FXK3N\VHT].bF,SNQL>YTG>X9?Q8G>O3FB8^0H7V>Z(L<+DGQ+/X:;,UY_HWG
Q0T1HBgZ4?DR[@S<Z+]-8e)]C4W#(+GVF+@gVIQ6+d99=>-Q5/9VM1SP5H4b@1,[
^&RcSKag9E/:;TD^_.ee4I:g<H=E^Y9+a\[4[7JN4<5QVB/@LYbW.[<OBL-&^310
2EQ=YNf8<b#5M95W=.QFaMGUOW[][ZB2Cc?dQ4UOXe(K51E^H,T:b[I0WFIbMLg;
bFX?[4):+K+A#TFIb=dYYBP0Y-D,Db28Y0OH1D,,BFX@#]1/Kc)CdFMOM27FG0YN
1>C<>MQ[Y&><9XJbQAB1B\eg8ecPc/GZaR.(S@TR&MQ_V?]=4MKAe?H2g5W]BHWH
:UE_V7&4U4VM2cPU6L,<S>d]#S@gcaf,1^XccK-=.K/HP6PQLNIg6=CCW.W0?RKT
:ME1;c92(Z.EYUL;.[LMC[<D3S232SXWJE\-XB#KJVg-H=4R3;HAMN<N7.;KaLN3
Z5TM?#[^fWS]JF=53=QCC\E#MC1&V:Od9V^23]B?-##S]]aYPIRFW@>6aI7ZIT3e
3OeR9aI5c<dH,LN@-+cNTBO)<JL2H]4fB(M6/OHGe<0^@1c2;M/@HCK^LfLM0)/a
JY1#/gdd2a.;B/Oa/(YI+^f^S#Vg8g(=F9;dVOS1=Ae/VV1SP/IC/#I^8NVeQQWg
W#2<VLcP-=.g.IA0E,QYfIPL-TMaNLNN,DSZ+6<Z3ROATCdCEY>M@ZL?)&0[P&)L
(d(&TNS:3D7>-YdgQWI(A#L9-8YS@gII9)3?7Z\S,TbeSOK=Z3+>119&)N:W6A>0
HOfAA;g.XN6Ee[TUc-T2+RGWZYTf+=#c.&-AHN<JUZ,PSO6DgEDXa^>NSO_ZS)LF
f0_XQ.H[:E@#G]]RR8SN,f^_=bKC^S/cM#e[5GR1c(SVZ)KG^=+WQFPNFaR5#COS
QVU]FB7B(f>7VdH).&O>4a;6=1B@9W7fAbB/NaUF/CU9.WNSOZa3TI+.&5/=T1=V
/O.)Pc0PJR3E+^)146HT[a^MDMfc7_OIF5CZ/^Y+9G34;KKPE8bA-\[6_T+:A@94
JIPG?[HW>-3K]X0O@?QNWL&]ddWcSC5gK#eNcRAHJEK2f;IA]1H@cC&=dD^X#5N]
@E2bB1e4-_^=>KD7S5K_YXQQFcE?PCZ,_D#74AT1H36aLTFQG>S)FN._b<>2<fG-
/FIX+e/(.-c-5fb:?+TR@T\ACY&+E0e,[UgAF5=\YFff)aY]O1JIQD1<@e]9R=T)
J=<BTA0U5M4I27:dFQf#cI_+VU<]F;3IZgO2185e04:KfG&3JLO&(6dX+>ERW[D_
eA-2KGZ_.[FbZ8GaaN5OZ/>W]f?DRa@M5:D.8EgfXHWT]0\aN#J&=L08f9U5C>KF
WN2,J_TM3[e]J[-[B1_XBXc)a<9f.gQDb^^;XU19dOLC5UQ;S:(Y3f(@/H&2eTZ@
7K.(:LHC:GN9O3,bR0A)R)SCQ8;cI+e7>S_=JF-C?:#cWAT]dOFD\,A(E+:=]cLV
-be4<XeU#6ZZ,PGRXfb_IMFG4:.T2&U\ZP@Q5>/3J_4@b+]_8HC>+]3T,DP;Uf^B
GN4#O^NNd&P/4&@@WeU]KN_E+?.bIH+3C-5]0<Nf7e?Kb>I2bc@fK)<W:#]1;GN.
DWRNVU)3C0G&,^9,JfUL_B71=EBP<c\SJ@I]O)C6O-V#ef_CXR>eO[^caKS_d^a<
3-(?]08B@aN\6QfUOJJ_UZXC3_<=:gE0/M:S;W)4<K?[JdH(N[)V72/ab8\?=<ed
K,dA]OUZ^;:dB)R8.D(HOYUYTE/8E-)O^9g^K->/Z,\2N_/,a#&T-a5;O7^/L<3I
KOWa7-UAGY\<P29R@:B?IgPDJDPR-SC[D=Lb+,[+fe0(=fBEGSX:Ga,0+FLe)V/7
=6/C_.XXa.E6TJQ=,Tbf+DeGE^+:[Q1#FN>;U\S,S-C)2,)bK\6>?)&+?e2aI6b^
3HS\39Fa)A\f,N-A9ZOB=;G4,(+JC8NUg0cccCL/d^G(@KA>Q6Q:SOFKPWQg?N).
Y.<NB/d2O_Q87O@K\PY2?J\6F>854=7eDU5:b.S9N#VEBAc.^[Rc^=CJ7\Z;F\\E
?)UaI7gd]8LFG>BVE42dF@B<AXJ090,SgWM7#gI.3)3R8;^T\JD(U?]fdQ2EU:M(
?DA/[1?D(>=9fV&]L35JT0^MHcV_QfZTXEV2@,^^@U=(Z9P]=RaS7EN(R2JLC]FW
1MIIJI<W(F:<Xd9<,ZERY8#\fe6P#O;3Z[=cA[[bFW0?5X7(1Rg(N8X69FM,9FOJ
EJE_N-POf4&-31\P0<1_5W=XWCG];UZG-\2^.QE30+dHT(77WKb;Y8R,W:WFR[>J
A>Ga+=?4E1^>]UZT-AC(6S:2V,,9P;\50MIMd<\ZSA0J[W(F&D=Cc2-J/F1]d1I8
N^ZIfUUD7/>Ae8->,IRE2ET<,GMJH#;JAegXF2XfHe0dd>OMA([0LLO_R6Y\-]T/
/(d;g;MbPSR7,D(S]NIb5(cO?b51JIU0XScbHR2^Q&>?ZI7UYB;;S?Uc&9T3RQ5\
ERCWeCNGe.VUVbZ^#:fVC:NbK(P1:C/K]6HO@M?:fdN6\Ye=Q+6KFHAU60eD9@^G
U.3Y>_G--3;58>Tc<Z/bOHHc46C.:QJ6BH_28(GNG/)=fQ9U2=DJ&b,8P0H3cAXM
4(:C?>MQU=X(CHeQ6B2C1a>B,02/N/@^30]Xa8#O83OQWT3MTaf0BPPQ[O=[I)SZ
=#LF#,FEMABFL-(;2T01LD5Ya/9&6cV+d\3(PV=#K?/GEOWPc6:,#(8,:g_MI75\
)U^]8@I1+gEV,c,MX;#KY8cV>@M<;,L#51:[KT4O6TM<C=J<#cH)+P.X;3F9V^dP
.B,X#Mf-5S?c_4M=(7@>P9f=F:IQJ_HZPKa&A/dWc+=]^)1WL(.(,C(_8:Sd?NJE
gA83\A]>E()c3^BW;DOGF5BJ78KCFT:9FbE=X;&a2bZ_<Qd.CG:UNba9S_B94<N,
9&27-OScI8)+3-YLL\WBYXVRZeU,N&f,4Xa=+e7^YUSbDe8Cb)SKYJ,;T5bBgTDU
FG.Y4e:ECc[CMf6H/=gX^?Y[&B04b,<(2P96C&/a@&OJGfc:_Ad8-e;8:@5W.]^a
J9/F.,:SUROVU=Gb_X8=4XAU]]:E,6C9)?<7RATX^e+2.TC^T9ZT@3>-\BE/de^\
_6C[F=e)_[7UVY9#;&L)C/XL&)S=9bE?Da4gMIRPe>Hec+C6CJ3bdSM30]0L<)1[
Red0:=1>>YT__X1PX?IA,[];V4KH=6CG6X?&Y[TdY6K#MDQ[;&Td7IQ&Q01/4;L-
MBbXafG>LTF]UI.=3I&ROEO:a\+6=FecLPfPOa?CV^\1Q@EPB-g]=9&UU6e_VAaa
[SD-6)&c3]g02dE40F/U;R^GcPXdG;:1>\ZBYFFaFb@/FI^],e_3.,2V]RL8RBP_
f-?O,.=_6LT(;6WD-,X)+9:PJ&;PI-(^f1VeO.J^0cTcHDFFBAE/f9B)?b?Xf^<V
1@BdB8<YMDQQD4=g0;>JK+2U.fXe.-<@\1;_;N8[V)XWVWZ#,YRRRc=QbXI8V62]
I-OUK7+&=?0)1c39Nd;:I@?-,H#^)A@aIfVFCeY0c+3O]5AB/_V?a/B4CRW..VBc
/DV&G@)fKR#S4Z9c=2<A3[5f)^0&I)D6Ya^R_6-@12TJ-@(G[b/cNQBDL0JC7gU(
=@-L402Z2O^>PNS?g+\SBUYOKU=/ZD5gUPHK?_,.QT-cE#TSLb#QeQ_6_ee0X+W6
7eD-44aK(SU@0H@-[HX2<TP>NB](+<>^:0X0KFDf.^^(-B9[.ES@WVVYXSVN>UgS
=[AfFU/WE\EZ@;U/+d^b[.&.N.#8V1PV9JTggWB](/UbCZ,-:G\<.IfG]]A2TW/J
L=6D;\UTH6EO56[eI^fMW3Nd22(@-K-4@CNSbKcM3>4:RT[6ED;UI4fWE&AF.A\5
@F\F5>;:D1BSIQE7GM;+XMC5L=1_gY\E<O7ZN]bN3>.,TOO,)=1gP-Q(AZD=W)3+
L49R+@bd27E/dO+<_+W5=17(S\[H7OZQ_UTd_ZeRd5bMA:^?F?-=?NDbTYT(YLd?
\c=I&AKCBPYPWGfX_4X_0U](+,Q-S6#9LQ_UBRcZ\9&8:J=\QTGe&gE-C_)X-I9\
&PY]2H<^<FadJWR=S-KPKR/SO/?YDUUg&V,&E@c)6=gPe]]3^8@&,\=<Z&^)_L,7
ITb+Oadf4C+aZ_.IO,_/,H60ebP1cXX>eWRMSZ_2B(B-I:U5-^U>GeE.:#39HbT]
<MYU+KQV,5de-P9Z98N(]C,#JHd8,=?#Pa6._SXMQ.U54L:O.AEX=KE&N3DTE5gO
a7I2aaCbJ,/-VP@H7X(WCS8X\GRZ9A;21:\J84@_cd+>NaJ@dcINU6_=L1-5BLBN
3[3T:GJXedUF2&)1\d=SOc0WFV-cA9[;&?HI.P:@?2<3E#?Z&^0cUPS>)ZX3VNd^
7cP#F]R,X4&e^X^3\f^W2_V]QJeT2.:e>JNW[53XH]87d.+#XG\Y9F&545)4g-R9
Sg^F^+b37KGZ6>8Sf,Z&eI&2egB8Z0ROJ;g=54?H-E)E7fU4)[K_;.?)b@0fUQTI
9#QA5bc2aSc8Nb9RR)V9HLRb.&KH,Fg1_G0F:&]CXeDLZ(6:SLV6:JD_bfC?;g-W
8fbY,#fR[O2HO0f(K@Ae5RLDUTALEFf_L\5TVVMNV]2JF)T9<:R^IfP]@ZRJe..X
]-BD?Y>\cO4G]^7O[BAF4&2NAI/B+b0M::<+[,Hc(&8/QT2BWH8+,@S\AT.T<C6;
L[SIVKYP8#fN6SBEf2]5dO[U-Beb9NL-+e_?6Wf^L]K2ZBfX7gYDBQET3CCIVT[[
G&+QN+L0D+SW^Y>RGFVO2JOE-RY7efN6TG8Q\381B5>g3_e>NEX\9R-aM5Q0bfg^
2fB]-f(dER2[J_\^CeC#[<FJV]Q4G@9&P5(Tc\)8c4(e)5-&(,0fN,fUS7V7PN>;
#-bDQFcS8ATY)(&J^M18Z[1ZD](0c;SBE:_1YBfLB8F,JKJ<@34@7UfaLOH?9P[;
5P?XV++<QT\\BX[<R2BTRNG3bTK)[(,4YEU_(XdN<P=SDAbZ9a.b-QTBVC8Cf^C]
d+[GRMID)cf7@VX2,EaZ>(#);cHI42;9B;fgY/+.KaM^P?MM^^R@>QVCa-eP94RH
1D&.21].dDH_G=G]g-TO.8:LB2d\)=N>]6D>S:42Z6HA3<bUHDPcNYX+Z@M;d-36
)0O#[e^Uf5-JVF14N;#&C&b02@=+We^W?=d\1H(2<MS-7G1/REZ7Id9FH,T[C-P3
4YR8UT9IE)_9ZT6UX+DNWQLJ^g(E@CJU?\)Nc/#<UDe]^5U7b<#fIS0>Hd#]=J@\
7@Z:fIA]W<[a/H\IZ&gXE+\8^CQFf>9>F6((Q6IeVe^5G-(4L0-Z5Ef4_HF/78e=
?.dNMMS?U_KIVPONQSQB/F0aD&3cDZRK\Oc.I#WDdMaLNG6^(ag3e6RY5&fPIRG?
eg)IKb_1+.;5>/QG[@^=6VE<:(;O\[E4D+fcHfXY)g61_d0GC+[X:+X[K6@Lbb^@
\,+EVB9&(;&B8dPIA-SPJe01PRLQ2d)V0V.bdDKS).+GV\_=ROI,?+\9^K2#_-X1
H>bAZOP^Ef_6GUXHH\1<L@[eFdJL(GP:M:6SCfgL44(6&4-H5ZQEFQTN5V5,aKMB
d-+e>0=);)XQMF,Hf[>/e)E&O@Ra[QO?3FgE#@;>FFH&QNIBD>:=0WH4&@Xa)#H=
R#b#M]ZH7(3GJLX/e?gB((CRR,O\=#\=Neg#J[?9QGE7RT;+4:RI3gEKJ=aS7.c-
<7H#2f(,Ke_AMgXcX7aMAHL&-F?7;ZL0(61V/c)?Q15aY5;ANMQCVQ^;^.MP7UK_
>C(Q/Pa<M=,IYG=A-KMA1VaME&H4QbG:dNCWWPc,HbK5L.;6UfK6,S_X,6C]Gc;T
(Ma;E5\CVSF+>.K)2XHR@86Q8RQ&AG9.X#EUZS1[KK;<HEcJSRR\0f^1BXL2W;YU
3R5AE:F:.VJ)8dD6=XNVg]6I@Y0IL(YI]S(^RU:G2A-ZD/E3719J,W:KHef&=6C?
cc8-/T9N]=W6/SJBB<=Bg3#([QT<d<PFDSUg3,,&U_&.2ef^Ma8>b^](#[N:ZaAU
TGK^9cZ[bdU7>6TIWe_5&a)\P;:6^3&B9JO4XVIVCO>O^FL2L2)XI?AP^>UcIeGP
FS]KILD9JT6FA8?8;8CO?[3IgFP=FbM\EOC_9HacaVZXI&(XT4(KC,R+3BSH-85a
DWXZ]X#-.f..I;&SWI524-J_6]^_&NdMTN>J>F=;=^/=de5P;K&IWO=#>YB71;VM
4d^B[<L]e4d;]Cd;L&0Ga1WM5P)b6]AM6LM=Q:?cH#+3=]3-.g9&#]BZ8E_MXPRC
2?]OKO<04<<V<<AEd5D?aYBaMB1/8R:=)3)=g/E\d-]2\F/&5X[G2]UXBJ,2P\7f
8+Y97_JEbH;^,P0O9<.5=PFANYHN\H];#-eN][XfE(0,5a8J,B,feP&_5G8e4C_H
7L7#>YDXKbRf:&X][d,Z3;+7g_8>SPQ+,WJ=?5WF5./ba;^<4U3TFVb8<=]1^.&.
TD/WcaW&dSCeO>O]a)[S;54WO^XS>5<:,M[>64HA@I:YC?[S+?PU<1GJVPC#>HMG
23MB41:#6ZL4XM>YM10:(@Q+aaMNAZ(Tf]B=)^&H,c]<HACELgQSC#\aLVgC4dO^
S>:]4ca0X=I5KSQUWC:GU3&DMJL?SbFX2(6=)=c#,331gFQAW)UT_V#08-BGYS<2
@JLc@>(Ga5+YHKc2602dJI/3:L(AO@0I/f1WN8T=ede2BF]+7K:/2E>Va-186TXX
XX8>3ZHa_16#-d4EEU/&[@Z>eP<5QL8Q6UBKYDSBC)BLHMe^_+V>JH.f1W1KP,fQ
A-?=OQJgS_V&74BP/?E^&V10>:;ZTYAbBZA/O),?fbO158_#T>?#HONb0>7:+df.
EXP@)Ue]?6c78?a99K:fK29A_[+LT02f/(CB,:(K(cT5<\UF7EM<\1G,<86:bUDZ
RS,1HQ7\P9c:.(@.Z24AW0LabL.U(^I<b4U>)-USK_3fX2C\B>=Wb+e<]-EE_MK)
M(dXP](_;FY[_LNgYV^G9DP,T9Ib18c81W3Z4VY\ZJI(3S21W2?gFAL@9K@6Y=Ib
>+X5-2Z,EUc7FaZa#Y@a(:&W4X5Wg_3JJc?OMN5E\A;?G;e1KMZ[E:(E</P=8d33
U^^XI^g3YT(Y?.-^/Ad-MGc@LBVX(5#Ha06e^-5bA5B5ZGA1fBaHW6NXFZMWXY]N
BZ:a.OJ&OM?RT8K(D?UA^?UJQ)8=Vc<(R=3>^4NcS_>JMG?>S-6N\2[e(eX0?)#\
WYHPNMDUTeHWa6J)f>CG4ZF5IN3]C69O3;-[#6D.E-7/90P@AISRAK5X6CA3G+9=
3<;Z@8^TQS#&JU(1.#?3W\5/+cQNVL(7Q65SaBD:H)2=K098b^<JG^0CB)6^>]@8
1XfK2ISPT4O5Q\ec8=fWJ,EM,FD/9^5Ea=\S(L>6W4eK]?V#I,[aa+ZAEZfN1eRH
,DC_QQ^SLY._WaQ(dJ?T7TE4f7b)V<E^CG2TU/F4_G24fNBMgG)Y7(GI7PQHT))+
<T^8C7d@)>b&D6d(6:0@JD_BNIM&D^JD5(bA-1/KFV3gH.E_M=cK](>AJ4AL<TT?
59fcBWMcddc?QRTGO3^Q.RT<7QW&_cN^^WMg++(OXFC\Ye6TI@:c5O?CTPPEb#?d
Ue1&7aWYA+4(4(8QdZabBKKd@P_.+24#5eHg=C<Xcg.#\JbTgZg+27W=-)7d2;BH
TX)T+\=,QIffXM(4RIJ+1U)A\>P/=]<76+Ib.>3G+@>\+4.=.1>[L8[H\K6NJG)8
O@A/EY0Bf>:VZ5XdXbEdH4)0g60L:6&>PG(?S[X[.V[VB>7:=)@,+P7>+D:&46-,
;DI84O#5J1VA(Cc&4RLYX6HB4\E66<&.JX&f91W.^G:&A9-,YW(HHL)C+8XCE(6_
9^-\cSHc,\83PWaBYXPa3F0C41g@LW@E4:b5>\_YbP?H48dD]LV[F8N0f9JaC@#)
EK(e,H:&2<H:@8CM_adWZ#ZY?,\F&Q,;TO)RORK:Q0Tc\7[MA]_VCAS@[?4E<Zb^
KID[0-3VC7IQ<f+B+cDA?2TN0X0E]CT_UOV+&.Rc/I?b\V4IVQT2#Y<g;^6ePVPP
L?WMX6K=#.?HB@c5JN67GC;_R/;(XV_/4f#1XXL]GE3XK^K/U[.bI6ca0WU7@bFJ
YA6Nc\@b;O5^dTRWRO]W#WefffcFe#M6B2A.PZ?1fe^Z;FXC44<d5\+W#8.:Y:RU
P@)G>U>NB/-AHb@((V)?41U=14M-,6W98FO+]N_41U2:8A&4Z\cG4C.c;5db=45N
,>XF;\Wg@C5XEG;[S&\(XUcT;ZD=HM_[F(+Y41,JcaMA\Z:bW,8UH23.G41[O3CG
HgU\,aZD36?1J?&;f&7+60>K#IZU\CK#Y53#BA(Y>?\K8B[8L8OI?1LMNGQ\[VN1
JD68C_L<F\d-](/UA_QTb7:gc/\&=d@^.;9b_@#)WbRX-T8&B8a?I)@?Q3I@<e>e
49B;D5W?8GU,F4FBWH)7AN9M1<b\Td:Jb55]KLE-#OR#b+^f.O&aGT,D\CNXB>H5
?3Q1<\C5)<6]:HgFZGY=_Lb[@5gGP]AR3L62EM(]<M#dSTbcae[UH\^T#5[:><#R
2#@/BHV[]dcfK3?:FFbN-f@>&dOZNf9KgB]Q6QO3K=UXY4[70EHeU:33Z@(5VH(V
f<c]6ga?]]M?(eGRK4-#LK062b>/^UZ4aXWLZ7U/T+T(N88[&/c=?;W:KUQIGgC8
[Q4cQ^Qf=X&W3/8R1Ga]M0F42/4K4G9R7EI.MHc&DD);(5VK772EW\._4d3^@T03
cE;_=1.>cI,1\:+f&UdSE76:ZeA[K0cG@K\5@^II-,G6NV7+W#>-;E77e.;\c=dc
QD8&M4e)/=1CGBRNZ84<S7WM?Lb8+@N:e<R8Y2M)<2Y1<._X0J9bJ^H^2<QM&]CL
KYM:c];2]6R,SJ;/09_=_UK\ZE;5E>:;PQ<Jgd]Q)F_GQ+(\fSCG]]U#(-SX9K2g
PMG;O[5gfKE_-f6M:P,_<NPD0HaPedb#G8=WW-T\;O[d[P/cfUM=CBF,I:T^-0Y(
]YH1=)ZL3+8@OIee??a34,-]+>ZSEPcI4@X4W?776]4H9fb+e^KI[0DeKdeV9XN]
Hcagf-cYW;+)_PG+M;XU]PcD72Z4fO+(a#aE8^C\0<@\/K0:bH>MX80IL;FZ&0+\
HY2b#cX@Q)QH(#RgDJ4JL8L<R<+fVJ03N[FN?6I<6.7NVCY9PB/b+U?K75V.<:EY
;,-3A8JcM^c(AL9DMZLZ:;NY+17#T]23d_#g5/F&+CD2/bG1YV>BRYFe.dIYP.Z:
DP9][8@OAH1Cc-B;O<Ca_C,35fLHUdO&Y#a,F^\g@C0>-a(S>T]e67DADMP;^dWX
b;QP?FI@7=;Q=RZ:51/J4O=gA/>M<H>2/2CVb;UA6ag,CM;>NI=0&Ne>AG9IZQ.3
8]NSgLMG4LU3APM,b]JBaQ0H.?\6MNPaD)DVeZ^[[^.;4UI3[_/K(Q=cLEP1L3a_
;0VFZ;DC-JY=XB6W7\d_6SB_99?8IB5O=HP[/3,6Vb@Vee>Pd;;@be/+Y1,3^_e>
?3H]50.TLVWD9e0\c?X](.aT)bM(/V^MR)W:NHYE,=_AU#55RFK@585\M:89fD9b
SWJ.g7X?K2S9U2Z-5ICMN/WR3XX<^1@9@,,ZIe;T\c)9WW?C/KX=::bH5V>V8+e^
Hg4I56?SeA9=\,91QeQ941C[(LMTSWQ@:L5^2HJY;+^=.G2,O=0A3JGF]:75PO4/
_>NW9G3d<^5A)aIa?]SS#[TT4SbU4]75[g20C.,XE)YXZF4#,7:@#^d/50.B@UIV
;;ee@CF4@FUZX52XACX6V01^>VBb:E\N8a_8&Qg.;.G.C>g<g_^-YS&a.1HSG-O8
Q1+TO,FfgS+G+2c_FWYa-9K,Ub+OUG<CP/#X#C3<3O<K-06]^g(77VR:;.F):7GM
JO6\99ce4;cMDa=E9JeRCf>[<4,HMH4C1DIJLTN)HM9@YC3d?G@R9+7_)+-72bV^
Q<,0D>VZQ#-#O:TP9_f=XgG#CW/g?M]<K[CVO29)8WG8[3HS)Q.;Zdd7fI>-gK)X
WHbfL+_1@fCT<:9Y?<8Eg1PefOAQ18O;(;GCN@#S&P_Q/[g;WR;gdJ2IM5IM6NWJ
FNeOS,D-<5GF^1/UHDP_DADB6R^d(FScXN24F)1;eUdc0M>eGJfdK3F<KG/N:PW_
Ye^J4.-)))Z;A:b??\KCOb,,F@G(+AM^_cJb@)\cb1O[g-:P#RCK:YJM9fH?HEP[
&X=8=4R<MUT24-dJQCGPG>M1;[DT^G[cJ8GN1I.8CU/gYBT(5@2Nd6OL?7A_)[YO
/G5N-Z[V-&#YRDSY3XbT;1K;18fE:ZA:]@AKI+UB9_:/&Vg^(28BgcH]Za(<fM3:
A24A.>IHfL>STZ0?S)C:6\0c?O52VgB=B)aYBU.L8G4@M?B?g,a441YCe#6E,)XF
KS:1DR&)/A(S&+]=CW2IM(AYJ[;Q_L:+dZd^,RK4_HCZ;?PMLXb7H;61Xg[8X_dY
+MVPcb[4<JB<R/^-b(D0:&B,gRd8(V:O\9gO/;(V3W.<F@O4E&FM,L]#_93VCbT9
JP-HGRB5C5Q=eUNICefg:c((gd=\f[5KdLUVV.L=<1QHH2)7V339:2.P^PE2?UG:
LMU\d]LZKKIfOJH27G+Y04e53Q3L?PB7].b7&a\;+E&OI?FGc]]#RWR)]JXd?8f&
OEE2ZP;Q6)9W0cb.1HEV<8.Cb-5LOU&M25&8@==F6W\NQA&Z,TT]fe_,(@NL/-=9
-eW@\:;:#OLKC4?K/a^9Za7(0/g<9fBVE)Z:d4<D-/eHZf]1\3fg,b.QI[AN>U(V
L#92M-,L\O)9X51H+adIGe]JAA3/:0+g\dQVNFAT^db)<KeT8AOKB?S+;#b_GHET
/e.bU80=R,/C<[aUV=7\3-)C5\cGT^cL&CfZUU_MQ[#7@G?<b:+UfX-ZP6;]dcbg
PFEDfgXY/cV4MAQ:@O3@N(:fOYc7S3AB:N\F;-=aV\c7?SgWZf(;SD:;.4-]JPM<
E6K_D0bb\gO;-MP2^SW4ZM.eLV.XF60^bS,/T\-;T>+CX?YMZS9+U[N[GB@g./]#
baObAR/gI[^]ZaUC_CBYTI-0_M1L^[Y3Qb17d0C&[dKC^0Re4Zd+VfE\)be]^#g+
bT=^RP.K1_.TEf6B,U+#UG6_;N9cH=XJ]V@Q]<b@g.V#RGJ[<?THPQQHPV<NQa&,
Y,DP.Q=4=QGR=f39RU+WT,[+LOL(]JaId9ec1,?7/..PV#g(+fdAK=ac<1a&DUWJ
MV>29,de)>F2.B38N=b,dIG)/AKC.Xed7VSUC(F#.+ggB+CU;5PfF8Kc,Q?e8G>7
.XF?DRL97:Q[6:e7e,TJ0TUA8O/MC)0B97f0A;_@/DdZ+],8IX2cEBf>FI5gDUL;
+]0>TRS#>;.EN?dRX5dK2X]4g>3UZPOHg2SDcXeY/;<YC[-M//Q3:+16e0#ZLRW[
F28Y,=S/)-E/fP3+7c]24X5Lcd?;PFa2OVB#S+ePWKA&.KMdD5IIg.M?CQ;T/IV2
L)O_\_G@NJA0J#N7IO4)+:W?ZV.1-C3:([_S\@#4aMSJ126fHG\-?R(D&)1YBY2L
f^>J\]2G>G1PA_HO?5?/VCT5O@2TdJ5W\YNSZ\bAJOd#T_P181cH0gVFA3&=608a
AX?YdALK6[YRA/N\Q_L.L,GXD,A03B^;;J1XcBQf9WbHJ;89G.[8eSYEN=[?Z>JL
-7P16PATK57Ua3BVDKgPQ:+dM@eIcNc2,W,./4)@WcZK9#e?X-f<LaP2M0+==bWc
^;L&3N,5Z7H43^GN/A#T3FH<O<NQ9W#\<P=OWa-WLZUf[1&UYBU(XB&=@DD<M1^>
ULJ13MNcXCSIcQbDb&2-F[&QC@UUg<N>9B^C,Nde.OG)eM/=A&)0+5,BD37Y11X(
@CVa?IP9J7KV11OM1>9F6f)VS4U5_dYILR4IG74gF?K\Ucc7WX-8#67K,W]K+[SU
;7TI2(G[2JNX,IU@dKOR[?TFUO4,-Rg.?EX5CTRQ<Sa0,81.dD9dB0DB+FU(=RBB
BB1,@230&E\5QE:D_=Q(@SfQ=00R5W]O)X5B>40d/5g_7WX(7&6f+2F]bP1dW3T+
C1SaODLRKTg#f]<NL^K;8<KHe?&Rfg\+VUTDa2+cMK_g#T5d3Yd?b<d#LVD-VV1M
7B-\PGKNG9Y+&WDF4X6P<6P2=Kb].?5H,S9?dgHZ^V1T&V0,.;VZTX>8S;8DZ^Ka
5=Z66Y_H3)27;U-a6._RQR+/2O#;bNG^8;&>e6YAEN\.aK^.V14>O#732NBCQJf^
UM^8A((&I+/fRLAS:./..F-R>g^bO[I.4=6#<./\9U.=4;0:GHU\9BL1IIDg_=b#
d7gNdF9F.E<.<#R+LBc;U:L@#OOD,]@4\d>BF3[8cZOcZfSgS4,]O[1KUOC(H4EU
\gK.J[2A6aLZ@TF7/T[^2R4G<((66#0WDaIGbQB44(WEVPAI&PeAXcc[F)W[TJCR
Y4C]J<KU]]51;[f<fdZE-YQ)PJcfRWIKeU<W3R@e7=aM&50UYUT,:f5&\MWEW;M)
[PG?7,CC+7d/WN(=F6eB.^M-HTN]AfgBHG>4_I?A0C43cGX@fNMW#Z9+&NgT66/<
-?-S:?5ZJRcG^PJ(W+,>+2^W<+/XN#CPX(d4K#P&e=<I9YSbd_\@@8Z2T]NJY=J(
U.)V?.[UE,B()KQ<PHYQ@9B3a8+.=6fRU?/cXW916Cb;+e1Y1\IZaa(H0E[WX-4=
/V]Q0/d3^_M@cb@/+XR]-&K25+c-.9@\L7G1KH:Y)R@D+5SDP25EE+I77X8KY)>[
UPb<YA6c5=>b#:<V,>K(Lc3BX6A;b.AcX_:gb1.d_OS9bCA[3-[C^YAJ#DWZ,&e[
U\^SOJIPXPb;EKc/dMCd:A3)D-C,+Y\M#V\?<;2_A^&&J3UQ4\IA@P1P54DAJ/C=
_X+TLSCUJgGGCDD@cdCNHJc4<\-YBQMSfOc]K]3L:#BP2GX.&IS.<_Q2I)8#E#^2
=8\?bOUEGg_1;KfQ>.gD__7\0DVJM@8>b@^=O]NEB[[BH(=C@+fC2WWN:R\@80Se
_11A_QfN3cfI7XgRBX;)WT[)932@/WNUW.g.::WWP-6TO92G0dcQ._31/d0Z@C+;
)T<f>#\><DH0[#&>(\@?GJH>L-TH=795ebC+&VR21)XN--7[XGOe6bX5gJ]9X/Gf
R8Z.5XIK[Q_]JHB@bf5=;B2C:YM?]XJ>g4cCN:TObd.5Q[\f^9#4Nd7<AL-#Pd@W
R1P/+JZC0PW]<_W?T80f#3/A;Z11eF[BOVeddd3(WK\)Yf\U<JG512-7#,]8B=-B
;DBGS&)TQd,7QPZ(S2H#6GR;Wa<Fb+C^(e7.&_Q68R4,,dT0^-_Kb<?8P>-WRHVA
IdE<?XfR_DZaJ3b8F:+Dfb1c<f4SB#g9;KS;R-&_O0D;a20^=O^>P\C]K[N:4OKM
2EZ4.)g0DR_R)?J9P>ef,M:<+S87XB=a^^+[D@6^-H4g9I2Q.GT?8(__Q[Ogf40[
A^&D,#TQ?g[M4(92>_JT;8M-(.RWGKCQ@[T#4(OR?3aVBe2(Y7(Qc#XdDcLLQ-:&
;ZQP/]26&N>R\:=b;MZ.)dYfK&Df#RLK1-e1G]TXa;?2A8RcH7T?K7YAV#1BX:C5
_NJgfS;#3\bf-3J6XXcHcH)K4WVP)Xd>7?]L-O?8#B=JIgZQTGLCeO/?3L1LN5LF
0H8,S_aG2Rc5D.(44CE#,C.N_#+\UX5#41L^Ud+O?AC3/[Md9H=N7SbY6.VcS\H/
c54DZeYOW;T[dUMK@SSc_76@(ZHI+g;CR+7-Ucg_>Xa5Qb/F[@#c>B)CC71<@)2b
SUS2;K9DWJc&:4-C.+Q]ARKTU7G/J_3QC[(gc3)I9HEJMc)C1.I4Q<<<.#K=gH7#
4JPJeaYRP>BXMS,O770=/DRMBZgGcA41Z[Y.;]P;aAge\@[I)DY&d[67LE;NVB86
TOE?:DA]T>SG<C_0ZTT)K.XB-6,T-MI_ZZW@+3Y3T)STD[Y<I,8LBP2^Sg6[I[OX
7,-WT#aW>0Vc6#+V9fK0(cF:+<X3_G&abS.fIa>^X@LJ+PNRM_@GI7)ZdIa86-^<
,Tb1>SAJd\=TJE_>,R<]64#CXePG^Gb3bd:dSE&P=?3ee+aD>GI>4.D9aYK9=,;8
=;+F3Jb1G7[Hf/IM?S6NYG?a0a0V_K^XNP0Q::3,17b?.]Q(F>:BX^SF;812[05I
?M4g6/F;,WfF01U6SKEE^c?9.EV?,+fO_D8O3Y+\b3+c]-X/=I8&9B/#UHER/QYY
0)g=6VHg1M,]9eCY-L5[GLC[+=>e[Y/I3#\Z-gd90A7cJK8\,P^Ec-bD4@=2=>+Z
J6RC5TD9NIXZ:99M6NEb[CBfM]M+2+SMbb]O#R[/MY^RSdQTB5,\aC-5GVBedUF4
S(J=[JNOCBH(<dTeYW<,AJRL:\S]E3E9,IXGHLI+[XAL_H\BS4[gV,^;LW(OO:(7
B/2-ZZe]XAD?.X68>]H/Ba0f^Sb,&^[G0eH-@cL2#EAP,94Z#A^-cf@?\CKg3GUg
SQPUW:+1.e2Q<(T1<VBO\U2RaVeAXLQ6ZK:E@AUBO_SdFA&\GPEX5QGd[Z<V#KS4
fd&Cd-dJ]4]#R+H<:IGBE54HFDdNK4e=-d\_M2]WS3.<Hfg_^:g;@ac)Q+O\N1I,
L>L_8dWYXe@+18R0B?N;+YRDG/&^]\._SXFL>cSQFSY>T7Gf/7_BFY5GWFSE-cXU
4/8>)CKLU)2V?LG&X3[cZJX:QHC?A+ZOg3.LT74T4W5#FTRYHT0D\bODA.\\-Na[
b<O30T=YN0\6^U^YLWfE9T7B.YYA[eb]_/c2<=,]2U9g&N5-eGZ8EXK/eQ3Z_g-6
g=I3eWM#:0#0U&aK.C#McI:,.N:#V;X_A#;G79+;M6[.1+@PM<=V0U5?_K=8ULM4
<g^+8??<b]M_)8df<7ag]:+Kc8YD4GXJR</]D/[?ef73gW;4^@Dc5N@4O8ee>4OT
(>^T=+V?:P9@L)C=X4&a&<VEVBD]VO>B\OQ9KMN9I06X55QWY?=e^>(/]>/PTXUW
NOZF:]KD.Cac30\2ebXgX1(bVAcId0(RJ?BP5gV#>-;=;FF[b9cMe95Z10#9&N6I
/_BKS[N;4eeC3?g=A<a^WD3X#(N.FU-_E66DCB(+]#\P;T2I0O(5RU/]-O4&BG>:
\aO&7J0+S,adSWOVSSI+&..UgXOF7]#0ZGa)>03Z2AP?PYLCa97#2]9Y/3Q\A0UF
/B^,6=&_9TbY8[@7GYDAQIg82<L3BTJ^#;[<;QbFb-6:3b]S;_SgXAT#:^@HI,2B
?MA)[KID)T.>Y;EI<fdDSJ5&GG56T/g42-Qg8Q17];8@[S7YbBXBMcQ.=J^gCNS7
EgC;eGAEZ13VA=a1/RdZf?U&^DN\2<0;_&3X,CMF5/L,7NG(b9CSTY=@DU59FE]A
fJP.934FD;Z?Mb#DGKFPQ6QcQ\\Uf-_(1Tg+EF6HE6HKB\<X8(Pb](b7BEC>I,78
>>]_XM9b=]<#5C@W4T2+DU;N9b;VdK.+52DC.JK81#GALX/VN@LS])LV+L/@g#1V
[HNN<DG[2\/02951FY+.Ybe9dJ[gTNWe>Gc4(Gb&40&4C.&6@.6>Z/V[b85YJ[c<
AdSK]G+)5G44b^_HKPc,ZG0PZ95),U7Q_6IG8e,fO&3)fACS3;2?E5ML;F_+(#MP
de^R>UXAK)QQ2&0f45KZZR-P[:D3RI\>@38Y,858KbQCJ@1;AY-->H:>/bF9F:98
WHXC)9gI1g9DV+a1YK3=aAD;R(bX.=+dE=XI=A,X0DO6S0&M5E_I>E(41bHg+XT-
P?cUFHG,9]a>X@X80VK,#&8I2PJF.3MQ35KP.\)B&U(2^BF3&WWbW?]-3>e2,/F(
PDTEV9SM=3R71fN8,C:WM5g#c_<B8GT\-CRfc@U9ggUDA/.XFSa+8OM<G;[[&ReE
[BU<EF#4T;JGR#gDO/9a,F#:(O:Ra0+C7_^+UMZ26K;7e&25B[TG:V>OHb_<;,M#
GR^\WG&&=X+@P#?2#4XCUVKTZ5;]cNdb]B2Be5Ub5?2,X[/8GG7+a9Ge9D&.P=3\
_BO6P-,T>D\@_((IB&73#@&)CPAg&^RBf6Y0:M)G1KN7FT_V,)3DF-e@BWV7>4I0
A?_OZ:7Z-0dJVE5@4a</DTM/9EXOBaTc1^J>+VHY1>45N9.S-0e@bB+M\bb(1Hd]
Z1QP2GMM3O0Qc#:X]SdgY///g=WN))/8M.B4.g):.\EM/cVg0:N6/#5Vg^K8K[YJ
:E11CfJ0.G2.0gBWB?Q5W#d-Y,UH5>U<g6VDXF^34IbdBSSJ1-]W>fBQ0>#WeH@9
(#;E6ZC56;,W2J_V3EV&(A+3C]F-AaMUS5D^]+WH(MZVE4VQULXO.)JMCZ.NfJW&
Y6,9^bc4b/>[@H:P@/\gd2F(@,I7f+dPAX?6>1(DNTE?1SF)A[CASQ;4V,6]/CB\
CKMOCE9M:2CXT_[JeKd?Df)47ISdV_-&Q^F111-fIZf49,SNC><JBG#MDF&Ab53:
@RIOSC9#MM^^-2=;&<UL2C]Z>>C34)2)^5F#L-Fce<;9?+GNP-#HE3A)(RF#bV+R
-K(dTN,1\1C1\.Y>gPBMG8_H/Y=V[b4#5>,2dMI6O4=OQSFLC#@_C5WC\@T:TSb,
F=gI7FP?6gca(Q&-/6/1TZ4KBcSCf-A7\bI#ceQ2eO#:K;0/gd.+P72V4)V64.C#
8XPJQ;5ZD]PC_V+d]NE]e[^G\]<9Cc+LaX@3U)g85\LR2Xa93WQQI=f=SdW+PJdZ
8gG9d-5+9VZcBCG>EcQ<,aCDf3ggW#A:VX&<]Jbf#X(DAMH>LB4)4FKTFIY40a;#
&d)\N]BF^,b96J#W:++@,-#cW@aFH+MRJ18::=?)dLUDF7_YeOOfa6K+eE?2@<H-
CSGB?.@NP)@T\CO8aMQ?ge[f1(N/)eU195=9f[?JKAVE5)A3)5^4>?@2&6W\5R#H
(JMWXD_8UC^SB2LUT1T6GZUIP(A[dK>bZ(/4N?6?O^eSO1C;95Y:JX_)58Xc@C)E
#)50OVCbdeH8KB<&]@f+gAX;GJX5W+1=dO722<H?(-;ITaT@5:Q(R^>#gJH>7E3-
8Bb9dA[Yg.8?;AY0RX/B52IICR8_Z-B[)d872<^.A22WR4U/G&cA<fH:/TC,.L+G
1@H_/=Ub&6GLB[3OOc#D_>QNBP9G(<,824Fe7H9WbE@5<&-_2+[)9GN<bHF0fAHd
g2>_5Bf;32YT02C->85^4-[K5Z]I],A-O-V6=FO_,8,4/RQ2g0S#9F9@M@/?>0X]
AMDJH(004K,PO+D:Q-Td05C>]7N>gCH?>L/._0.eb+J&VV:BRW@6YG.\#41a,63C
[OUB+F46UJ=T\?CUBM?94N]c];@3W6BC94;Q><6J\c0Na8QIP7>90Q3HV,-_/<=K
+K1B4=[ZUd3RId<Gb<EUcE4A7SO2)C\B)CZQLL_Q]33cdS(I,bb-9@-QRZ<^7e.c
D=aN?gAYN6[S?+I++Y_If[E1J,+<#(J0+3,-UB?TLE:V5GUX^Q,NcR<0F;dD(>>K
J[H;_Na9>([I;6HSJ0?-@_P,gRgX&>N,:FOMIT>gb=bQ>86MCdf]N?]g;_.\ZQBc
&ZE.RA+J[3#>g+Y:C3b/X>/N)TNW3Ce1,0Ma?I#L4M)6QTP)d@OG6YeK3JNYYO2U
AA4^WON+0g,)b/c-U,&O>\I#<#6:Y0dNNA02eZQ^Cd-C_3J;._=W<,T3H0cYaE>.
?UP7+d&ZAaWX,^?@gV<Q?6G=MK?]GHOY=[g43^Ogg4?A&G0/9U2T2VV<&\_].)bQ
ADAMYdMPQ.7_QJ<6YR>/]@.2+^,BAH.0([5e1?B8IDYA\-VKX(Y9B>S9^=eZ8<=R
)9<AND;9VQXbeTBeJ)V1F8\2KdeLT.Mg_A@,.NQ9^R>L0aZ4U@0Q0Q3ZQ)16:W;f
CT):]R6)B;EGS[&H#)][f\Gf\^Z<R-VEH+V9c3AZQMWTF56_CXS-U+9?D.8]E<ZH
9;-7_\(K5.ObM-]<-\ZJ_V=Z6\_Z;DM0R?.P^375g(U0?6KK4ULd1_eF7OD1N-X/
UbU)75O\5-\IKU\?M;=;G+cYgMGU2a;6DUdB>3Y<-\25A?\<?9_RNDLZ\/4X_7b3
dKDg39JT&[@PXXW(VQ;2@79.H<dYC6Zd+S+^HZCX51^aI+4U[\-JA>&\[61aCSOF
H=+_YL4OT_/IW_?N\24/4C^E#2QBf8F)E<D792=(6N(bY@HfQEU&5Zg.07d)fHgJ
)ab?YaR;I/2[aT=6(JUB[bAIeCeb,g?dOfJ?[1V.aQLa[JF7Y^[&-XA=ITJUWJ:G
P4EZJ,_&T:ALX2dG)dBeWT\^Z&5X;FZb3;QKNCRO_M-],@g6@8&7c:dQG&4(T4IO
=0&O/WMb>MOg8D2SQ/@J_]D]Z_Q644.f3#+O#<L9]8D;;Nb5XN(3dVI0DPA/MEfE
_gFb6?R:G0<c.fTbg_6Nd+MVe8#^&0,&E1eEgM@:WbN^&@:U=6\d7)QH\(OUUF><
(SaF_e,4@.a6Yg.g1fAP1:0^ggVVdAeVadB].KFZ6L_LJKBf<EaWE0]@809F#UJG
;Y7Hb^[eEc/Ue=3D+Vg6^WI.g<TN[-.WNO&L3E>[)COdN\G8LNgN+@;SFIM[RS@0
H?(=D,?:C,]?3L)N/O0a[89A-e7MRX]G>$
`endprotected


`endif
