
`ifndef GUARD_SVT_AHB_MASTER_AGENT_SV
`define GUARD_SVT_AHB_MASTER_AGENT_SV

// =============================================================================
/** The svt_ahb_master_agent encapsulates the sequencer, driver and master
 * monitor. The svt_ahb_master_agent can be configured to operate in active
 * mode and passive mode. The user can provide AHB sequences to the sequencer.
 * The svt_ahb_master_agent is configured using the
 * #svt_ahb_master_configuration object.  The master configuration should be
 * provided to the agent in the build phase of the test.  Within the agent, the
 * driver gets sequence items from the sequencer. The driver then drives the
 * AHB transactions on the AHB bus. The driver and monitor components within
 * the agent call callback methods at various phases of execution of the AHB
 * transaction. After the AHB transaction on the bus is complete, the completed
 * sequence item is provided to the analysis port of the monitor in both active
 * and passive mode, which can be used by the testbench.
 */

class svt_ahb_master_agent extends svt_agent;

  // ***************************************************************************
  // Type Definitions
  // ***************************************************************************
  typedef virtual svt_ahb_master_if svt_ahb_master_vif;

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** AHB Master virtual interface */
  svt_ahb_master_vif vif;

  /** AHB svt_ahb_master Driver */
  svt_ahb_master driver;

  /** AHB System Monitor */
  svt_ahb_master_monitor monitor; 

  /** AHB svt_ahb_master Sequencer */
  svt_ahb_master_transaction_sequencer sequencer;

`ifdef SVT_UVM_TECHNOLOGY
  /** TLM Generic Payload Sequencer */
  svt_ahb_tlm_generic_payload_sequencer tlm_generic_payload_sequencer;

  /** AMBA-PV blocking AXI transaction socket interface */
  uvm_tlm_b_target_socket#(svt_ahb_master_agent, uvm_tlm_generic_payload) b_fwd;


  /** Handle for uvm_reg_block, which will created and passed by the user from the env or test during the build_phase, when the uvm_reg_enable is set to 1.
 */
  uvm_reg_block    ahb_regmodel;

 /** Handle for svt_ahb_reg_adapter, which will get created if the uvm_reg_enable is set to 1 during the build_phase */
  svt_ahb_reg_adapter reg2ahb_adapter ;
`endif
 
  /** AHB External Master Index */
  int ahb_external_port_id = -1;

  /** AHB External Master Agent Configuration */ 
  svt_ahb_master_configuration ahb_external_port_cfg;

  /** AHB svt_ahb_master coverage callback handle*/

  /** Callback which implements transaction reporting and tracing */
  svt_ahb_master_monitor_transaction_report_callback xact_report_cb;

  /** Reference to the system wide sequence item report. */
  svt_sequence_item_report sys_seq_item_report;

/** @cond PRIVATE */
  /** AHB master transaction coverage callback handle*/
  svt_ahb_master_monitor_def_cov_callback svt_ahb_master_trans_cov_cb;
  
  /** AHB master Signal coverage callbacks */
  svt_ahb_master_monitor_def_toggle_cov_callback#(virtual svt_ahb_master_if.svt_ahb_monitor_modport) svt_ahb_master_toggle_cov_cb;
  svt_ahb_master_monitor_def_state_cov_callback#(virtual svt_ahb_master_if.svt_ahb_monitor_modport)  svt_ahb_master_state_cov_cb;

  /** Callback which implements xml generation for Protocol Analyzer */
  svt_ahb_master_monitor_pa_writer_callback master_xml_writer_cb;
  
  /** Writer used in callbacks to generate XML/FSDB output for pa */
  protected svt_xml_writer xml_writer = null;

  /** System Memory Manager backdoor */
  protected svt_ahb_mem_system_backdoor mem_system_backdoor;

  // TO DO

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Configuration object copy to be used in set/get operations. */
   protected svt_ahb_master_configuration cfg_snapshot;
  
  /** AHB Master Monitor Callback Instance for System Checker */
  svt_ahb_master_monitor_system_checker_callback system_checker_cb;
  
  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
  /** Configuration object for this transactor. */
  local svt_ahb_master_configuration cfg; 

  /** Address mapper for this master component */
  local svt_ahb_mem_address_mapper mem_addr_mapper;
/** @endcond */

  // ****************************************************************************
  // Field Macros
  // ****************************************************************************
  `svt_xvm_component_utils_begin(svt_ahb_master_agent)
    `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE);
  `svt_xvm_component_utils_end

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * CONSTRUCTOR: Create a new agent instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, `SVT_XVM(component) parent);

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the #driver and #sequencer components if configured as an
   * active component.
   * Costructs the #monitor component if configured as active or passive component.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void build();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Connect Phase
   * Connects the #driver and #sequencer TLM ports if configured as a UVM_ACTIVE
   * component.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void connect_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void connect();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Run phase used here to set is_active parameter (ACTIVE or PASSIVE) for master_if
   * Start the TLM GP layering sequence if TLM GP sequencer is used.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif  

`ifdef SVT_UVM_TECHNOLOGY
  /** @cond PRIVATE */

  // ---------------------------------------------------------------------------
  /**
   * Forward TLM 2 implementation
   */
  extern virtual task b_transport(uvm_tlm_generic_payload gp,
                                  uvm_tlm_time            delay);

  /** @endcond */
`endif

  // ---------------------------------------------------------------------------
  /**
   * Extract Phase
   * Close out the XML file if it is enabled
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void extract_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void extract();
`endif

  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  /**
   * Updates the agent configuration with data from the supplied object.
   * This method always results in a call to reconfigure() for contained components.
   */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** @cond PRIVATE */
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  /** 
    * Retruns the report on performance metrics as a string
    * @return A string with the performance report
    */
  extern function string get_performance_report();

  /** @endcond */

/** @cond PRIVATE */
  /**
   * Obtain the address mapper for this slave
   */
  extern function svt_ahb_mem_address_mapper get_mem_address_mapper();
/** @endcond */

  extern function svt_ahb_mem_system_backdoor get_mem_system_backdoor();
  /**
   * Set the external port id and port configuration
   */
  extern function set_external_agents_props(input int port_idx= -1, input svt_ahb_master_configuration port_cfg);

  /** 
   * Gets the name of this agent
   */
  extern function string get_requester_name();
  
  //----------------------------------------------------------------------------
  /**
   * Function to get the configuration that should be stored for this component
   * when debug_opts have been enabled.
   *
   * @param cfg The configuration that has been supplied to reconfigure.
   * @return The configuration that is to be stored.
   */
  extern virtual function svt_configuration get_debug_opts_cfg(svt_configuration cfg);
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ezDxm7qMOAc9R/C4On6PiC+BB+ff4sGcJVP2a2zSWUp5dwDmvAPuhO0u6fZlmaOp
j6qXols5KNxrO/t/4PNLJSaFBgR4WrRVSMU/LcLStuv4kQijAkGFdutcwQOS+n8D
rRkKmXX/7KgEFpoerIRfca4vAw/LREQEzu84aXm4Wc+1Er6uajP5bQ==
//pragma protect end_key_block
//pragma protect digest_block
7s5uehy5InrH6YFBQXo2g/XmoVI=
//pragma protect end_digest_block
//pragma protect data_block
Ux4qumBiZDnLLogWj9Dc0evXEeXUCga4lGYsDZVYesRXc+pKwH9uzkl7+ru0FgzV
S9buauL59Cmd+CFwFiXRKHyEl7/m5nfODndRh+Lcy6z4NjN1Dmlk+oi05b4sXT5l
kknvmBadZ/bNexnVzSAzU5tCwMjuTCg+OVpsro+KCi5ZPv7jgf4yhQXQ9Zt6YgZF
MLZJdd7xpFcfMDBukr48IApSCBOO2ncpls673unG8Ow8gP7p9zqLYEcXg16DZk8L
PIWz43vZJr704MrCGvq+jSOBioyFHcYxGrFMRAqyZZYVU1Tk88/0VdpeyV6gEFaN
T6WV2qk6IuL+G87l24akuQqXxuKB9VeVsHVtxfjQ5vOEygxv+eQ7smbpv5Bn654z
uvcFQSCnoq3K3c784mtUqCuutv23U8r1rwkwiwk+JpwXMfDJL+4WFM1ouiUML/1W
U51Au3xj0bOu4Hp8aBaNH1ZlcdT+YtwSpPLAHObuESSUuIjCaH5DS/QRQNsHy6NF
DZV5jmmb//tSqCzlucBf4LxevZthYX5iMDyoJsuhn11YYeftOH4MZAmz0BLJ+G3e
6xmGhwcsmENJB3l3uvnR4hU4WemyWz/imMr4SmzhDl6g1QTTyk/b/NADWAkHdEPH
4W1StV/JlF+qjtJ5KZE4XWZq7qWz58A7fLOT04I+g5c=
//pragma protect end_data_block
//pragma protect digest_block
sRYU2EzIvZtqKIQP2AhQarCEwGw=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
xz/mqUSBxhVYE+PWEfjf6QZtIl/ApXGa2UNBqEsGix4tQY1609gKEXGlCen7oiSw
YCYTd/Gvno1rN431Hv4plQ96cz63oL91Ssl2ePiENlVC64Yv3ySHIxRFGG0hFlbs
D07d0KEp9YPnPKtfQMhQzWRn6OyDVaeY7lOWwCujM6/ESIKf7wD88A==
//pragma protect end_key_block
//pragma protect digest_block
57OyjZx0xILII8O9Y++5l8Ncdww=
//pragma protect end_digest_block
//pragma protect data_block
Va59nAP7W0Q0WevDMzklbAga8iy6HehkBKY34rG0LPOT3MEQZwuC1OabZlnyl1Qm
lNbtpGxv4/qriAc+P9+vQ1Dbh4Uo9TQLKb0x3PoFsyEPPpqenF91Y9u8yjxwp78E
59BH8YPgNosKV4cP/kUlO+UwEgtYwAGMdzHmAbPFuwRzmL3udNJ9EU+7NFF8Yqp3
XAeBYLWf5A1ni2poRKnBTfTM3ksDWIMa0VYToJ+cURs5ebxk4NQXaTP7JzFX2bqe
y0Pwfkhnj7k2otE5r+bfwG+3JO8/iPrW7iKx/ec52odYfYmR0HqW+shK2nwFeANs
tgnOr0RxdWHC5LaUeOiywm9E8B/e32pdJnyFiHfk0aZKskqClvRsOD6nPH3U5wzN
pAweP9mHL4vavdpiblUSR/FzLh0vUZT6tudA215zQXNnWPigG8Petsjx5zdWmVNN
aprerkZZqEO6oIM0kshx5Wye91E6KbblRgjiDsicLlXLrlAcVx+2O7quB/3lUE26
vyTqUIQEwWjvDE1l2fVu0bfUDVroB5xCEkIIy5rXN3Y+3KAjX00Q2ZyupxkPOUoK
JaZuTK2ow/W5Zz2qrDKFy+YcZd2aCNs2n5W0sCtbXKrH/2XrXQ4fECxBkjl7L/l+
knpXyl08mMGkZXhLCIle5ffTSvH4+gG8HYPnIQG7WYBK6ShJWWg7Zl1GgT8Iu7F1
I9ooja5JkSkCpDIwpO7DBLxLDta5CK1k7m6uTmjyuw4P7Runx2t/a2y19xsq4kBR
Ajc5Lyl76npJcALMfhqBp/eLawVhQZA9q4BSmJlyETGI1GTDol1nULoZqd6IeFKZ
xyzUKO7ANZ3q/uuvVxTzJf5nuYrr+gS2+0GmN1kQF9ddIaA91cNYHVnbc1nb0dlp
6PpRMtLhph4zeRToE3UfGOnndeMKDYrSkrxeGFKyDfSY7gBa0++RpHpJQYkiiX98
Mhn+LroRnoNTS5xLFgLvPI7TRPz2z18UEz4B6pkGRiUp3e8HAHTmPJNp9p9s3FAr
s6GzSOQ/k+GZ/oTlNCeT8Bh0Fdm675PjVH5CA+VwtcO3FsNzWOGjb8DYH+GAvxO8
PrVoNEr+uA6PutIOjNWoW5ZpENT05KX/sy+7QN5+2alA7IsgeeeO8x70Y5GIeWTw
HfCPmoj+xM3v1KUTj49hDUALOi2LoEsgCma1Zb2eM1LG3d2YDCFAxDSd5OegUJJg
ubgRk9JpL4j5JLiIk68023sbZNUSyzuPuVO+aEz3BBa8ogmgGfkmhNmgnaxEjdDS
MQ9eLHI0vdS3/gwR2PTd7aPPQRh4Ew/hUbHAOl7s0mX3KsSyVKBM8sv1EGxlYOf8
MVZwIWAV+Ljo/+dG7Di4dGuGpJ3wpy61TieLdxxh3ALa85jFtQu2E2GL1MYVbeuQ
HieClZSRZ+tQoQAKCwE3cAwAcN3zKlhh6wuJa/1Bi7pK34Vo8ASaoG+GD4EL+f/G
iVZWNTy+kYcvOxg2/q9fB2pq8rPiqseQN+h7gQRNlBnzpTAx2L/+vzCkteiFMd/d
4LACT/XXjsC5I+vU6mZUzIsOjX6umTTVsrhCZqBM2cN5wT91fcQ58RhID2o2X9lk
qaK63G0fpM1BhlhpETohxO6O3ScmpHRrksCsNqQw8h88AurawatLJd1vKIZc4g88
DHKZws8OUXLeBFStGkhYj5end3KHbFSzdeowbV22RxnQuX8vaWr5GM6PuuWwH32w
KKplpnwP6qBZRQ3HpKuAMQypciFGJfqDjZaaNtf2d4aOFbV8ocv0DlQ1+A3fm6te
JOHvX5DfHG0WPUjt1Q10DMsUCY+TYEUU1w2cfLQjXLYu6B0mM707r9PacCcMcxuE
P2tkj/LsyYumNvuPEXhZ6g1fNzQ15+Ka6vtA2801HbzOIzVf/mLqw7HQGDtQ4V0s
pbYXCzK40bYdoH6WA40lE5hxX98/nco53hQ1ZcqA7N7iiaqTxhJ4fuobsTUWTIFt
0+qI0V6yCV8r1jEBU3f0sRQwTMT/0EuMrvNxMX1NXKadu5NgBSkjXI0KNryocSr6
JgQk65qvAHRrgDXdQaN6WZP50Kql3yz0XXG20mO3SW9FT6pIClqAEu9tBxGZrLdQ
7hbrl6LHQdtok3J9hPOQClIBebjAbesICZQGQFSjp/GjypGlR0nwCcPfy+xkTq1j
d8+nVx43sSlxo7enMAjttyveuyMLvzOVC5oQY7SzlEqBV2m9ljuGx8Ngh3QQeE6E
qaCCCEYZq3ddXRpGHQ2pJ5aChXqZcYhfF8mW2cO7YFHJl+ttYWW+6YvOdSzP3vlT
ZhxuKrgUkx8+f7ur03x+FZddOW0NAtXKkzmPSVLIIj8qdF49MkV5WVWTIycmbjZ6
40ZzzD7JzVSqUK5LcEDanC22PrvHbmzgig5uF/S5WV9Roxcm+KJAVQ7NA6sF9w6k
7bzhAyoM3XAQe0PK2qOshxn928pBLHAVLSRHFEb93CyDHlz7MvdMlr4llIvgzAH5
P5/v23jART50ezXv9JiGKX914oxGZNH5SFtDeTInj+MzCSKK/f29O1fpeYR2piVs
iuQNH8ZBNhyJZwcO7XQ2VenJbGGwahDzv5MYG0CjfPQGJgpFFpkmZW0dt+FJwIx/
Ggr3Y6ocR50XUcDH7QzXm7FA3E3BeklX02JFj4WnQoW9xhlpdtypB9tbnOTOH9k9
2vFe/nBrxM3JnAx0UF4qg6rRCQMnfjdSWAF5nmkvz3PDnjOZtde0O1DaOl+Z9V5z
D1PXrv5t/eTnDWkhSoR0YuVwM7rLhCUuTtIqtV9lChVAvukcyh9VW6M8tyMe378w
VgDpveWysWMD3MTVVzkPJOnVC7ceavfnp/88StBzqDHdn2X+V01y0DPR0NfmpSnJ
pZ0zv0XPx208cIfF7E0J9sOWSOPkbrQTziIxjWdpBmbm/1wFiG8RG0x0uIYq8rbj
fwB+j11+VS6x4ZkLMDGZD8nPwFHdsfpmvI+Ky+XB5p540Z9FjEXGB365URUgJuLK
gsL3y+9+W8HJxZ3kW0XTB5dafoWngO7j+hjhps5Sy5MCVySroWCCKWDWZCo3g+tx
i0KTd8XpG6uwkKZNYvfVlB9Rndkgb+O8xCIxgQ+5OPgh9Aw+7//mFCmDhed8zW7X
bfN2ouN2irH8bA+SOhPtLiLbAizBOOn3M3VweLriUOm23uQkvSeu1RYhqLuiooCZ
IE2NJYNgH27rY0gYQYZKNE5+AeeBIdO1PgsiNzKYSoH7FdENzKXjlwPn6iUi95kh
K7j82RAQdhASrmdbOY+C7+rypU0Viee+JP3AbFNLTlijpkrp84OZoXDaUIF9hfKg
GB0Nc27ZeHE3HlUJwgLgkqyj9qsxgPK2bFB7VFur/hnk7Rf9pM0SAX7ZX770p3P1
5XAPmGcuG3LgjF+Scaood1cj5wxTC2aGSfM/1+BcSEfTwURcJxM/K2w7IxaRJ/3B
8iKCHjeuyYE/9zJsWSNpaUDfgOb+Thl0oZ/H59TpTLZx2Q/WrWk+nOGIE3LYoKiw
cvcBvxBthKuenFoKZLYYVvo4h6qOPI10X/qSbaCq9k0KvLc/H//Hpr9ivFzUcl2D
M4Frng9yTg28YPiQecJHWh6oc3bgtY8carWZCHazA2hqecvupCp1+Qt7vuVbi3gs
iXfb5OUufhg7CTuP3NESlwxUk0nB/AO/lVIpUCsOZan7Q0nXsSYWeWTBDzVi045n
RKpxQHi962IHHajFFtY0TuGTt4+/My7gEKMxjev1elLb7YewuJrPutBvpa32dfQF
5nHh0ORgJxD3rx4f0fTg5CYCzNVx6I3GeeKvby1nQ+Ruq2iq91pGYA9YIV0v5mVW
Q8wmTpfj9yu/rYGpa+oJn7SpJiJbq0x906F1njGePKW+cOOjBxI4N9tP71siry8R
DZdUcIQaROpJqhGV+mJaUH9g31Zv/Jdmwu34huG2PIA8mwjo+RkbQYXZV/COQh/c
x2nez4a0IJPL6ACfWaGjmylulI0fJvFmz18Mf+iZd9J2mBTAd61wgHwwg76Xpguz
iktjNJlfyl4rMVZ7uOzaNXqioaJJUZuGZKQZJrcK20PvIJu+dTxweIEE3KnfOww1
o61dkIy9V+zohhhRLCS1kamh92vnANyN6XjSM1BrMztETgNdh75BI7+lwX6Q9qCQ
4YskgKXAfi8CAZWDztjMVCmAVzKlN1P0ElLg2EBbOjwVsJ6eg2H2sNZa8+eoGMkk
JGl794tJmV/0OI8m8oZl459Dav28D0/L2TJEWzRJymjLKfPuX9ZxC60ggyifLUT/
Hh7tnDTQqLftLCaKs3YJo6I+uf/vJVsVaaqAPoAxI5wFD1Czt1SrEXI6/5+aDobC
3USiXhV5nz/R54iJBrkMBR1QsdQmGQ6/FSeNxHwDO1QrBbzynP8WnJ3qewYswptv
R6AC5mrX+xZE2zWmwaJL7GFEScoSuKO6a17XxTYWhcw/8ZPW4bxrOHuTTJexcylk
mvKc60omJ7J0OxLixiLv1iS3lPWz4f+NYtBRHIJLJV07Y3WB+20MQyGFcet1nWSN
ag0yIghXUM7kUil7JrFXwmcVxyCfzm/5W7Vhmq/gXUrkUoskYeGAqJy2LUH51fQ3
YU/YuhRiDfbo+JxotgufLJGgtH3sB/1WiViHpPF6kK1trVdczJuHDGZXikiccrxw
zY1hrls7ujkNXqQ4VWuof6lYN811/cjOB2k7uFjFwOQAfbcfOjz/uqv5tRY9AFaW
ax+dq0ed/7fH6PG2qtIz01WXmqsWjvo91NZ6UmWvoDuQ4+xiTBc9784FUrdeV5b7
Vave3q1CLWIoYwmy0gJnCI6y3Xj+ozDQ4daUDZB83AZeaEOfV9aqQLlIpmtYAH9H
0kZ9X2NWr2R3YiBFc48XvjZfr7sdprgkLipde9jPOwKoC8m0hMTbjxfnm2xPi1EL
jKp8ao37NAkbVJGTCz27if5qIXPnZZNjdbYC7vG/dN8jy9PQ7WAyxtVgEO64gIz/
LD4i4AH/xXYLvWVHKd+3z4h3HRJRNodL22o6skBgiBu+1RbqxLmPBggYyKf+9Sw2
QlilGScAym1504uvS9RpiJRSnYeP+pYlDhjInrXbKeiB/T1QwcQ4jxnouvJAUm7b
GzCK1Srp9wmr1vpLG/YdEdNLORCIi+vyB1Nk2885H/KcnftBai236r1/4+dhbPsv
6H/eyj93lzrmURRIba8D2D8nUat5Bjp13el3lCG5pSCaF6/z7nOppq/l1Sbvswgj
/YQfqrVyf3yWp2ByzFz6g7VD9vO+ZXTrP8UgSzWzIDx3wwd0ZbNXMU/rnCxwmY9J
NymL+VB7FOxYHJb8+5Yp+PcouqxSSK2pjV+gMzu5vrnQY6BKOA+mOb8z1ZGw7t54
FDqU+5SBxsVi3BjY7uGc8NNEu9DBmdCFGBccvbbEOhv7xmZz8vv9PO1gDIZhDLAb
tfK4AqBgqqJxFQa2g1funOjLF4TEYH4EbyFDeHkwhetAX+TikWnUR2dEoto+Hdiz
lpAlg3Aef6u2SuyUJ6THUDtkC1VcJ9qDAuJvz01kHYR5k2Ze2KxpSNsVOr/sSQ7y
BG4U7RcyabxYSf4WNjs5bFGh0e9eEXYUVVCVh8JIUoFApS8QAleGyBHXc+bxnwqQ
rst/2JvKZcyCMaFC+58xwsxCvrVyc3nRVRAsphxhf9GN/mw47zH50psLBix7QdNT
KIouudQ7tMvldVc+SfYfNFTWsWO2l5grtbc72DYHH7mUbCMczBG7A6v+UG5iRD6V
bVGP+qwiFbeP3Zl55fjib4yvjPYlkSHyIYLx/1ey5cRBDJVGUK8Jjxaz2nJLqzaL
iz8k5ZDrLMCPCwYND6smR3bEa9icTURDYOePW5U/YJeb4aQtChr2ACnnctj0VsaN
Ngbavwl/oAdEoiVM0IddWauBPj3df2KXRRbv6jAIxpj4iKVSk7lpPaaQd/9L3cys
k6KkPSOaSHZNaBZtGd0qBUVLzPtNmrzBC401a5rKkj7+9xJX+PtBIcNtSwkbiFNl
TjtX5fjch3y5BmxgXVbpEhMo5yKcg+C3iNm9SFE+uwXxomRP8VVWxWGVp74sew6r
vJo0Oy0Efgpc5XO+CTgrnTb9Umn4PngUCCsCAsdM6CsuYUCXwpijhdH29y+0bCIz
ZkLHUFMuY1rNoqckm5UULdC+WE6ah0ZY1TXdavJGHdJtglIinm1zz/NJ5WzLfQ5L
Ay9y9yEPPB7RGzxta2Ej/Ni3dzNgODxuN9/RmXkAibsQ6hEBoy8LdIjvxFTMjAcY
+j6+VWOCtlJwvLyEG+yqy5qFbLt53Z2lDoMyI/nwiIbh/Us00l7z9T39h8cbQh5j
X3izNCFLVL8lV95ja/yHLLhT9rnhCNdA9alucwV/VeE2bdL0dxxCUT+He64j1UU8
5118i4+6MadfDPZC2/xS77nEQESS//5rOl1t2sVL4WMZ+hxnoNLaJNMNhHP35CWQ
9EKy8yP9qqizg+yRsozKhUfIUmoseUUTVs7sUINsnZaLfETIJ6jHoX6ikGp0I1zK
P58XF5dEjwCRKafe+Sz4yPtsWq5+Tg/s4Snr3am+lDBDvNNtKX+mZx0npHUqsRbo
29C3cmoIEGFoydU6EF5KTfUxFKFPXfcswYlE6y5Taa5IaCZv8CnKvHcxw3+1dRnv
sjZNe/GdGzCCxarnLRty3fIKg/bL7t5sj7xAiCvKXSBi2t1Wf5fWH0hDwjshXmo0
Y58cG3bTj1yId3U2HKYQ+ThDC85lgWqlj2BkQvUO1m8tCz3z8NeJtmPhVyny6uaz
evqIKSL24NyoraspirF8m4kjCYtPRPcr80pXN83Ov3cRSsQQEj8M3duGiHDyNZDd
cH1i4uueLFZ3ilIDHYq7wqyy2yxRtL5byan+Fv1ZTzJ9TCeCymiA9NvZ+U3pyOdI
FrMPZ90Ny194MV5+y2cKZbw220A3U631nS5gQkSHGb405sd5QgW6qpzBf0ZwVrBD
4n6B+Di9CsnTEIPd2hu23RblX7zfQMcCfNUyRzYAmMl8rpyA5NbOrTHwshJfEyZZ
qLGSg4uDJ4Qb0tNGv9tWJtlEJuC0rerEJM8babE0lnIndJDxWre63EERqE4JTkJg
fV4xjxj4GUfwH4rC8MFSbSBCtAPAm/VnfPS4wfmmDuGnH4LMqW3AYIydQjoQ2YkH
/aHTXEz6BAqhN34iO9W+r0P8m1uiQaOlaibo4xXThVirvecrzlQuInnT3ZcieMdt
x589lJboZPvgtv3qUeBz40ECuMXk6Iw4t2aWoBzuNez7gYXlLOQwVIhEEfRiha9y
kT34wNidT3WVTTi5DBGh2sqzNZ39TmR/k9m9KMhUxtKKqOlLrq4qbkh/k2zCjgZ1
q3DiztVl8jRLjMYKy93ZZhl+xVFiPbfiYRJF5QlD8pjIrUx7ly94uBJ2G5w7pWDM
BabKAThgX6NmdTG5cOm3GK7xIjmURvGQFiV8FTuoIH4gH5o9k1PtDNnlPfCSLjWr
VvKW5583m54upvVhZmMIMH86+RRklrJXzBkqBAfFRKv/6GwmySnwJNQzGsrBEYoE
h4y5xn+b2tt6NqV0eE/am7OmWNI3K8tBTntYDFSvSJXPqjhsIKIOr3IzaHsoBnOk
FoatT0j/ex6jaWXa/QmH/jcQA3bcTUnCTc9oKb7cyoInMpzTdcpRC7i1VJrzonXN
ODuCAjsJzZsgj1WNvelf4wuvveGB16pCMD+hwsgHCpowszCqGX4th8+KUjGBx8a+
pp7JcbyY0ECO6vgaprdqFAQDFZunckLXhzWE4c2iZ06oxnIzt5uNao1MW+SBwSQd
FhxMAwF/n3UcldCU1Hj5PqAL8177KvengPHJHzJ7tFzsGLyMeNOVHZsY5wDE1a4o
WNL3QODdan9gKgDZzt2VBgW16rRXJ+hPCmcNco8RHR0Tu34yTh2ufrcvwLN5eKxp
11nfxTtDvHZ5D+rcSsgtkd1NReH9+iDrKy9ZTbioCvMB2q34/rzT+jp7D85uR2CL
S8vdJ0eONcFN1ql8u9YiTvVJZf9DYVZnX10l0t+zO/8aHwt050dd5rf6TCGD7bu3
7c77ZamS5RkhXwVKc1NKOjaSd1kR1WUyFRx8nYJ2tULPtihm98U4Klymer0gBWlQ
w40r687k3BLm+M2aYlMjzUrYTOxU6QNqWbv0lEg7uqvUh+yCHKBsvz+NARplD9W4
XSW0X7otEMY8+gVYkmsNxYb38z7Z7ctfUhbGxQvaXLD6/sJ27/jazGzcNT/TL/0o
di/+bzWmSRdfsubwvcWsPt8K10MIBUTFvh99K3njDMbDhvdOwoVi/ZWvXWML/was
ZZK3Pb2zaNVdEF8kVXryEUujAP3YgVh1uy3ctnKDjznDF7IWU7MdZWeoJYG859sT
C3QEcP+6jVAMuSqFp3xclR1ahAKFnu0h1VBUzbsF/RcHXxN7nJFz3J7RaNd0eoE2
4fJsKwe1Q0CQ3JGaTSSXXluOLJTgwwJb64+dDS6XkHCLWp9/eqqcJRtJ7ZjgoCWp
wXp//YvT5KV8WrYZsJJlQazNsSQjPKmrixnZK41OcYxxLJHJrJFaDE6ygcBJiVUi
upz729Ioo5g3wjn5zwzXMlXBOiBycY4/twSGWAGE7ed4tpYLwEV0vWbXgEmLJWnn
bwtkhk7t7YO/iDYP1SoYkeRPzggoOwXs0veCX4Rsf75V6zcvw+c7XnfkWIuVweo1
gk+p24Tp4+mdgKf8CuwnstTXMAVBzXfmQ31jf1G22qSCMKclx0tT8m1DniLKMILq
1UDs+mMW1dIXpfhowaUioUHvu7932Wx2/1cECKfUb/RrVJ8uDfG28ifMpJhiv0zs
IyMavNwDC7OCym+7LbmJq80mExHlrcksbK+/umYvijlsnR4BahWunR3A3pciJPl5
Z46WUOZjZ54iG7owzSEkoVVROCln7hoEvNLhlioseeTEHNxp1YfNwpLSEPhM2rO5
6QGeGXLrToNPSmLSUyXr5aiIUXdBNyKrxiDtCU1cQ3J1CMPqmeN6D2xoMmsljmvr
y4jHRUyS/5FQhgOOS5dFJSTb1Ry3tFxoDNMF1tSdYGkrhzQOGbI5Iikd46XdRmC8
f0s/cNVQcI+c1IUHV7MgVtlyE9lJbF+1VqdV791UW4j4AU9wxPEs9KE+2y6E/4Sy
begFBQ5wrvDNRmDckBExRB3xOHVHb0Kkftf8ErdxC+174lsqA2KE7qqc64uOlI3/
W2GyJ7QOxRmu5O7v9vKliHbyxvC3YSw1ZoN+Zoa6mLl4vXZl3HYsPvgYl9N2Tq65
tk5XzT91s6vMyVuUduUjCMUhvsGIJ2CFVxKyDBPXh4xrey58jBK+ZrmXzBv2eGFL
qZI5ONAx9saVXkrrxodjDkRiiFEAI6dY6GX2dZati1+ovJPYG8AMMlZ/gVUinQFO
gBqiEmf/cONsC4zSjrH7RKqUTNM8JhIGEiH/NRmWJg6VzfHn1KsvZC9UyVBBFlWi
4Khm3rExUj85d/yXdFY9U3pfM32CifML45zo4ngggBkJDIMXysUZMCZ/IUeZtazL
9hA/SoiOOhYmqToCMSnxAG24EzujdtFfF5eLqqQQIh7jrR1drz+o8bJJDcpU+GR1
T71xln0jH30VTx5tr0piZGvUWqid4tgGYoTLbOSe+vV+uFKHvozYqW3jih0DjwHe
2XGafcUYdVgxkoKmbWUmqUVPrEX4/jRmyCyZ6pIbCKL4S/tV6aOR/1TptkKr7V7N
M9q0LvwqbCTdQB137kA3+JUoyq3PAyeISmjBNryxWwe7/E9uT7gsG62ftKC4S2Ck
sRzaJvh3q2baXnIeSjVZeDVpjKpgzdoGmAtbYZ6u9vd3tQw9xJrtuMekEAh2lRj5
VZk6Rh2mqBaYRIgk6uImPrYyVSSqCiaxoho7DpzApG87q1AfSaVPiY4+hOc1XtGK
YR7Jw/6ADalwKzWT54hQrRligF4cnMWx6H8Fx4SgW4V9oJh2uvHMebkVARBNNEKt
juR8Uj6cA9Ig00up7472Jf1KGS3p7wAwQ101mT0a0lp1R3Tz8QK8W6rfPwZuzyq2
UmegGrCTDMFR5fX4WTxRH3uI/co740Kqt6R7IWcDCXeTFXsNrHVf58qyIW7XSZhY
Th5z9T6p7PzERqmMFl+Ig59PioY+1e+CarW3lH5Lml7OKNbILUnw/KsDkx5W/7WB
hDCUW4tEjBIe1ebh2+FNwm9HRsZ8QrSVfylln01x4s5wHw1tjMEIkb+x6SAhfNvU
W1SoezPTokU5XhfbqIupUz0BJ1ObTOxR0cW1ncH3UBIK5D5YZjyixxaxbK91dbsv
Q19qIi+mHnjMwo/C/tJKK63+EuBreoMK6E8FtY88RleriNuR4YzbpYo0khIAp3JF
Lb1MjOf4O0elP7I4Xyyydb+HYfQNWWepCKxcsVd81jOBC41vx1VIkvGVkhkQ3C1H
0GAAUzzMEBjDZdxWm+Kd1oc1gkMRt4rQOzkJEYGCOGJQ+uFtSFLzB3pI8uskX4SX
7LXzrRVLWXuOL2ze+J7LRlB5ronuUBBcMaJb6Y0K9/zqgT34lTFd+R6Zlx+CkRM4
yU8DWYqtSlOKWKGrBW6cNuxV5wOAMY6WIG5dw8SkvvSD1JVwBak24dAVc7VFMA8A
0KKIiFBtaY6KaRm0uyx2UxfuH9bFPU5E5wahhyE/PR49Hz1/9IqCIRODf3XLajF/
zUAbos3Bxvkozum/OGQN9jiMpDdNaqtu0W3aFL7QDBcnBfLeTnIwnVWe2lb+DEXY
n+LZ2aYUMKBqOWXLSbCb3PWzkjk3uMYjm+Pu//KNsSz+YOEDMcJRDTyNiNudbR1Z
WjDEelRJ1M9vhGs8N3vz11if7ZJNU5R0tvMQuHqNsCWwHZLF4BP/1wjvz5tKpuaa
mWk8/WTs9l9hripjGTyLoC9vl4QO4fa2uFZVHbGmZRA3eeTTros8i7EnDR125ULC
NZ6cmQyfNc+HBD08OXW7mEMIAKMkqPEnNFJR/yVX+4xNzXcNhBO3GUVzfMvL910C
FugekUxwP2RaK4QQdMpxjF5LHtsUeJDF1r8+tk7CUpj1KrxwWlNxfFIPKgwrrX5Q
Ikio6OPKAjyoAhDoykoS838fowUJXRSIEB7UyStTOLVbUZFA4vIi8pkQaRf/8awx
2swJdJYZC5AWyAMLCwl8uRqxtoMmGUkM+WYgw17y/hZXjubHZ3s72wWRORoPyU+I
V7adgPfLAEzqqMwLrUB5gmd8z2M1PFyi5cu/0cKPUDNg0QRx3dor4Ca7aYlansdl
fTyj3/a49rUicVhB8GjOABEskz7xqgFiuf0o/EoZRIMQQNwOsL/6mA4Mgb90CFHY
Tr+DMOX+8lROqHuaPc7b2h6XX2LcWRFr584wcauLA9hyfoiI8xB4yA4YbZdT5Sj0
i+76Rpsl3Yi5gUYE5GxWPcujeQ98QtEUilPNqHNH+ITJmdjP/elWfNqHya6eMH3c
VnIKiwQqmNdjbWtYo/1klGqEK/mJVEaO3paNL/HIXC3+m/5g/Alfw59p0jXGQuky
jLMDVrAPw57clGZVwnSNONrR1dK7bbVnYwWru0hlJoZMASr4//0GtvJE+B6IpYli
nq99QUCC3b6tdU9cAWM9kJ/7RV6Hy9m49aEIsQa58b8N25iWdQwFeGr+2+78Rs1P
7UQ5j16R8oa/4tgNO2jkKi43K3yHiv+21CLjqZp1O71frg+i2NlMowJmR4YXUVSO
WHd1JaUlGjq9BGodGdm21fnuMxOReLloH27XjxZdgdki3VxDeBNFOuhCJvXGSdXD
35eK9wMRa5Vr7SVL5A7EDq5uIZipqx/SHfKs/eUB5KURrRgsKKH5Sb97pv7Jx4jG
J0+uaAb3HK1wQQmGAYbpzun2Lj1sXkyOBbeQvR/dhZiDbBsF2j9eRopD0lg8joH/
CPQqgYnnTL95r/oa8dzBPH1/HAS+TUIXoIYeOH9/cQaHuFl1hDc83cQGNpwA8X+9
1LYY3DiaVWQ/5WLb2RdKdFEWuk5eW0GIe+zv8TqDEOOS1Ka34UHWcAW3pL9tZ7Ix
Sz8dyTwhUUX8J2Z4Ih0X0ZpADg8bbDqLPXoVQEei1u7MTtQSBFemtx+iJZxgcHhC
A4o3DKeO0oxoz3+P8Cib7TE8AeU9huXi0OQC4hbN5Z7iDJRqGL4S3c9kw9neFmf1
KQYpBhKMNRWLUNvXV1WX4AvFlQ77Lb2CcW0Mi88aMf2uZSKwb/cuTEpxoaHaeY5g
0H85CtDJXR0cRnRNwGUjmiyIt6pr9AMKpVQbNxuAPbcYNiXgHyN1F4xtFkYgMrwA
fIjtUFAUssjSkp+8ds48C1RAW9Zrf+Lnb8oiUSbRdJFwIPT0eeR51cjpQaxsI0Fa
vHAwfYWznsmQr97JRJShhQtSmijc1uIGssZ/1jhTwqA6aFEb5ROghoUUjiuB3ulG
ioMGmNuJibrpPICbjbtOign/23kmheFr+IF18SNWDhvF6jLmU7YnAjAYAUnYT/n1
lq1HGzwTuwl5BEwHRfao4GfjmhMBTrKtIs+rKZ0ev3ZcYV0NoLrkvJgq3ksYfnz4
0nN4B84YKjiK9UlISJ0o9n+6b2AbsHupevJS4XwdlPKS6K/caw27e6ezmZsnAr+e
RHa38a7x1rSXN04qwSCGSXZ2HKSuPdq9PFCNcQZPYmcc+uww9aDqQON26u2s0UDL
NrGv5iZN/WUu0KAFW+mUS35aNV//d3VmNjCvmIiu5TwVboGsakTHV3n6bWDXpB4o
9afsj6CaDEzequdDbf4izjLC3iNt9SIu8SJqHZK/LhWsC15p6ba23V82bAKqidrQ
RHBbOhP5weZknOjZVKhkaQ/TGXS4ebj0yuYbVzoXGaqOzBEeowJovNf+D7q4K9Fp
pwIC0Ip09a1VMmuqjZsG06yQhVQUGBuyApHSN9EoJrYlNJjsJSrgrVjIbCxl3QEd
2XkfMIIg3Ijv8f0B9aWNVboLJvMKcjbL+PwREoKUq1XKN9WekVPyfEoxKRUlfO8A
OumB+COH/cBTRypN5WNllgTCkKz4u4OOOnl9o0EfPnKasmkiAAq+uWe2hefOeDdE
KkpImjn9htxiIv6SSD4SY+RZCLqJlVs5SzZTJUJ4mHYVXc/sxkTPeDTpfZNOxFM9
RXygslaxTGIDlAnMZ1WPBd3/u3wWSlMt8OGVEgwuDY75HDc/ekUYOP3YmhfeMBnh
EAxjjPW6coKMOwEcOTP9SPMdJp0WOzV1hPn/E+TVsYrYvvIH+db4azi5FvuciKbE
hJqIndpcgCQlqaqzr8bZfFHA0Ez1LpUuOy2baM3j9mAAuBXEwQ24lDaJLOv13hSx
oGS7FQpfpEhYS8btnxiYPZIgBbqqlD5qVrkkxRLmYXRx/ej4xviBSO7m24mShCfc
40sdA5WqKyoIEQSpbMUgafUG3fo1YqsMa79mRQzYx23SwR12AziA/yRLQGKi65HY
T+g6NQPzkK0Vd7W8UlELGYB/oFDCLwIXy+FYvhEfUxhvSSUvbizHypsaoNWbKvco
gRq8EsChi1F2dKuz+30f0V529/VJeHUc/yufIKYyI49moSE+R5d6dzgenAkivUXh
TArvy2umETFFKdVAgZN2MXWCEPu6IHdpXgaYDX2MYkUezPDUN1L+JASarHsYsJ7U
ltyn8SaeW4QxepfppfAZiRUX1CjLPKFIYYN3tTUrDcoESV+pahH498SnHutepPV8
1zOquiQe9swZJXI7ovuq2UeeovUD21EbZLJ17zXynNWjpJekKBgWjLsWp1lzyk86
rcyPZXZN3Nqbci0SkiqUTolNcthi7jF5s+KcamUg407fzQWkB8GoVi8s13D+zA8W
VQGPL2+6w7FdkELSauT4dN/bkJeWUTLkkLY5UjcKLDVLfEjmoasuMB2Y8kTCtrSU
KkTb2I7IndQ2NGyCHXZNm0KqIS8njDGeilXMgSdTuiZ8jt4YIHByoty6yoEFEiOB
JU4k89VAJ8Kw3iHZAZAiTJUHf/TfMtXrGuLcO5YScUuNooGLoyd6WLel01blqH19
9Q3TrNafsxAa6GVNakJyZCZptB6DylQ4PJdBtXFR7dKIxhfYPnhBSXyT4kmpn0AO
p48FeE1EpnnYAtVJwB7OhXiMb/PR0bOfurAJbZMM/1RIbYr1SC2IM359aPoLvC4J
KrpiOHlnAihNKyxKDxXxQarVCJ/PEkCDM6Yy2mlPtLvAGPs19IXzVXDgBXPvW+i3
58GatBB0Sh9pmeB1ZdoCcJak1bddelO61oiV/nHnFSJ6EV4NHcVweuUShBffpOpa
nKh0eOmCOudskrlRErrwNm7GpC6hPPrn1zsdw0bB5GEJ+bxFyJorHiFr7rU7NmcA
mCDRsdqzkD6Q2+n0Dzn/Gxewbgad/zoot0etL0JIKIHaIf5ENRv32Nho6v3AHovw
PfRTiLAd9PuEv4F2wI0q/NAQChi37Crge8A9ee+/GNdDfJkiO23v2pOZL4M2wiZ/
nL+ZJ6Se4zZfwYpcByq74JjC2hBKRaCoVyqhS4uTIakV4/9EZv/tSP2AfET2Oo/8
s1Gc7QzXSs24DQcc8G2wfxTYC3hrhlO6CWLQU8+0Rvc0KLKT7NTp2zWSRLCvl2py
kpD71pApvfZdd3xohUR/Zm7kMz38pNAYValIPjNL2hkR34LzOqvJhzDuaVvQLLNJ
5UXrpoNkc9MfJuyNHnZjh6FSWlVxt3ZeOSZsazjtsz89VXMdXPTzTER8nNqZhF4Q
hZvu+TTLfn8GnEPEcBcMwC2MJ10fyleBFYzCCqRXSlIi7IhI1GnM2Io0cQR/Nful
ZLN1dLKEOXRUZpUS8SNRURZsDiJsdsZHPT9/ERprUczq5E1mK9WinC5LW+sRtYmm
q7K3HHwDwndY2+AD4E4CAXs8t35pcwjL7x9RudIjFbfyUtPICAJ2vOxPlN6ea5HP
AYRReSnQO3+x79ovUB7gfT4ovSUom0K2jVCG7i3XFe8W8c5TtGFmRxBCIVYF0dPd
V9XU0hZGFla/EFp+WM7L2jKqulzu+Cjoe+oCQnk4RfIOeb55YrgZBsveeyIPrcLx
ZHTwxGwCfEJoZU4azbtDKm8kv42ZpefvqXCqXo4XhlWO/Ddd3W5pX3wU4PH5xvp0
fIGkQGuX3d++Onp6wIHyfPTy76bSgZPtOyKWXiL2+Qj6x2fl7zbcM8Yq62gMAjNV
lXw1mSlLk9DVc4aC3SsOYdOSpGvPG1ASKZBpNHN6csMs61XRCYAXBBgw/7bDz2fI
NRpcu4v2xnbY7M9oADLMn0KVI3L5zXj2GPdd49ra5Jf0S4E8wQCag4JlLi6sYhpp
2dHCVOQa66HfVDSmydu3J8A4p3RBSgFfibdJtjdQveC3hodlXhqZW4J0KLOkK/Kt
qiSICH9Z546p1hfokaLN+LoKEKTZQOfeCB19DyKy7P7lPBaszYfriUSGHjjJti2m
cWDROH7i9MVl8jlfJW3Vmic85Pe4cbFMzrE6k6UWSvpBLK8mRjZgDbF8INxL2Z3P
jY21ScfHmp9A+8o8BHx9wIZ4JulAJ0Ax0IktFtUY27z8trsrlQ2sA7GW2zs0QDmf
Iu0O41Jk17zF8E9RiK3gTE/u9pT+HsLNhoPtSio0u0zMqOBcS6hfG1w6raSYV9Id
tDalodDmrvW9GK2fKMtf7e6EBjqenpqCEZMqqzdxQh3uQHmL6pxVQNNCPG2fxr/V
TvZmoIZA667Am28UlqXN/EzrT01hx3vHxlMfQSKvB3WooL9a9VD/uFkPoMqgfnm/
UWtalYSjtARW1J2GxLFV+ZPJSyzLNOD2PBM3bWNBv6yftV/+fd5b1hQvE5BF2qLu
kaN4mSndg87fkLuSIgU04FrMLpzLWQuNTAScmTkl7o5caUCl6mII3G7KmiT/G2QF
pIKr03V6T0PTjKTvs5/Ksj1YjRqKAkG8tX3aK/sfot+Se+hc+54OXdEo2NjIJqD/
O0c3PYFD7TxMJAxzmWAWvqFVeccarbUWUKUFK7+x2WI6z7g/frvtBDv630CpIwuW
exhOnZjXCnh3Uz8eKb6p4l3b/ylOLav2inmapfq+/WX1lVrja8M2H6ENigTib2Bl
jCtP9N4wqJ5rEMU+cLZ9sdzVuQXuyrgiIRZAzulZtL8pxx8aGnIwTBNLyT4Mmep+
MtBMVb+o9wztw7qDY85Q8U2xXZmCiFnL0vayV1VAekG0OfFpS7YlwwwvRCFZ3KRV
L60ZBtjvB7E1z0KtRBct7F6TGIBnoTsyg9cXjWilhX2DwaognLmwrp9MSy6G1/wF
+TtD+AwMM9k+W145Ca7KG+kxmOKAIMhlPfjN5MgdYtaOUKlPoecdmOviaXyhvsRF
m5TqSx9UbEfuBuMKUTpH2JZ6+pmwV3W64dfloaRsxntI4RnI52qDTy+TGHs8s2XQ
o+vIXjwKmDvUllDETmvXpHRUn/vsKpOsqbh3iVQVTSA+UAcnR5dDrAGRkPr+8tCr
Q1ut+yfqUJN76ar6SHm9uxplESy+nMC4RmCC3wQTHtUHqn30b8AQx5XH6kHvyjKF
rL+y5vUPsnA++Fhypm8KEVS0YgXCPkZNQmnEIVNKGg+scsXg45ZQPTIUtZctIWuI
UdbNwBYqAE2iSGV9bbDxMFe3+4c/IMnVEsCk2pvOWng9qBds2lAFezx/o7jALzzR
OsFeWIfhib4R3Qwh9R4Y6M5RnJnIil1/7zZ4yiQEh5Nm40vednoICYlc+teSPEFM
8A72vqiJ8Ww5xCR498z56/xVfZsAM5/Lnwjc6l+JZlo5lrLsZdOn9KNEsNtanMNh
VpyzF3yWTIPyNZmXMCIGWNP7Yij9C4F0vpgT7FsYOQ1ockx+q0+LJuMYOoqwBfmv
9cBIHzpZw/K6FQZN0Yhgt9mD8KqhsSG5qVvNfbtXaLMQJdDi2huLPk8dfXN3T/0r
dC65iDli+/VIPfilz5EFkhHzYhQtIIBI3eiFKTMux5hwGTl4O5DqxwAONe6WFD9V
vou43JBuHMJ8T1fywbvS/qhuD5A5gUjBeqHNUZqVEuyUS9+1yhRNQkOsRcCGtJMS
D8ArbXGasa1AzzYQJNPGFyiO65WYffrpw77H7KKg+YutljGHQuKh973PHcBeL3S/
WUIRUJIWmr/9DcDCojz0WSRWElfIW1a3V13h0flhw1FR2lNf33ODXoOxQwNY0BMe
FPxMJkvmmU51G88fuHwxmc3JoViD5gW9uYPwaZ7m/IRcmefXmgxXCXzkuaFEa3mm
Iuz+F8VVNJekNe8cYDWbgWsAb6ZSKkfCEFQbKM025k0ssVyOc07QPvXal2Aq7zjy
YL/gRB39h4af11i1JJkdO5/UHAdtVy4J4YhHWdaWH2lxWiz8U7CoGRJIeJ1Lp1J4
yHvUIuExNpadBIu8WfgddkCYKLSnt9vfbFpSKoHTQOvZU4UUmAZd3Y0sXlJqsNM3
6UtxUskn8Mc3umD3e6VMpBlEWHUUwgbK24+iQxok0hgjllqNIRtiRFyQPdxxQoE4
6Lb1v03NSGwkYTF/+TBOKH1uECmQFzkHQQ9V/GgZXQ3u+04aa8vkIDnFSJdlqpJ6
WCJp5NG66kNu4zl13j0krkRMV1GRGA9/7EuRUPG6QGvAxm5aOxW4bA+/6nvDfdG2
DGYTzzIoC4MhFAst9lvCMsOObFLjWuIvc5Wc6FojSopuy9MIAY+b1TKHH3YHLE86
0MEKnKxYGXZJfiV6GOuOKN1WakkZtSJD3u4ctNdb0Wzc6LUcLzWq9r9+dl3khqxw
Dt1GUKJxRP+LlzydwOh1wPeOGSc5cVDfNjS6L6MuYHkXZ+2hxd5+D1X2c22Q1Vol
U6Jl+qq/2L7+rMJ5d8Xn1YRHD/usQUKyg5uNyDkbq2x8+PmdfOBxKDmjQ3I2HxFC
rc/CkNe32eNCJELecA6k4JW3OWX5OWxKopJBsd5yYjziY+2KUc4wFBE9RJuPwbKt
AIHtAAhH/OxJr98qC4a9NzCNz1bEpgaUl/2HcnRH0vqIo1f78PeLUePzCNEL/rKk
E6WpznMMA6PtVNeBZKBMBjJE8iICpLZZ6b6li6miDUl+NCWr8jwTd2/pOO/2MqU5
rP1hoOw6KR/eHDQmd/8Xiczoip8vzj8KC061OpAlOKUtmvbHEvUAi73Tx3bXoGbh
FGE0EnFmTNQVpyogAj+d7iJwWzEv3TW3k575k0YSdeNeF+XZBluXRfD8oU9x8MUC
nS84xFOMLLnyTJ2zAY6xjNx60kuBxk0lwRtCQF9vB0XEkUDnV4362k2Qc+mOPjCJ
4WobSZwyns5lnFc/8zqG/aq6Sd1mgGu0GadZuC7w9TtukS95UzbY0pm+2bfAbf2K
3RWAsk3qbANxh4BGAAXPg7N8Sg8Y0k8rSFSAFmMFcX5Dz1d32s6Yg4lZn05SX/V+
kLbVKU+e3DXzX5cDC+iYooJ82lMyh0aFhDYGWx99Lc1z5snox+YCseiv+9R+isdP
nywBy5jxy1F7c3fOPbNwf+GxB1Nld/lHtas5SS0c+O1vk4F8hRIGBNQPuQGAd9si
r4P2kJfR7V1fnwIzwkND4iXNiDtbwpQoj1Nk6DYsOf1Qhc7DjwkC/ruLGUKOaxYy
SI6PR4VtwFxtVnOR2hZQZzW8BT2/B0Wx90qCeWbNuXGtRiDJrCToxCbT7rkF5WX8
ncbwQClq0kcMcYm6TRAYHOgAJD5UI8xBIY2hVYwwvDHOIXQhZWG5V7NRvhTTJxTH
2Jc8e0WaMSRV6+ONidRr6Co8JZ8t4X3wLXejzS2C4DyYmrPakAF3ZpIBmA/YQfzW
FXtJl3UmHQAJ0JQKO1UQGWjlx+VsndXZVk/QnUg/NqXqwmT26OxxLY7R3QUiVUCB
IHgX/Gj3xtvaFDGre4MwqCgCyMypwegTX8W8jNQrQKb4SCRpOaxkcfuIKt5wagX2
hrQhuosRfbMBNlz7B+awOtv/xeqXTlrF6deI4ivcpc6fh3zOxWMs5YD7lU5uDheK
xSJ9yLroUVVxACDcq3LE78LjYi6CrF7PLUN3l1ks0SvcTLkTQB88MoMH/JZlcFgW
DyqmNcNnIInzUi27ZZ4Z57MJCiGKEWETf62oOtBGOYk34MkHnE9vbQFqZXI+/6J6
v7R0rZM3MiJ+aYiLzsmZ/RzdwvKa2RnaVEdtdEIF5Gr5gd3LYKmNNETE9FZoBeVe
+Z/PbYDV8H2MbmJ9dCS4tGimgbHeOBL9T0+h1MQAPGzJ6pO+we9wXzRUzvkKr9fj
wNeypf8NmN2vTq3G9Z3uBz8VIoL7RfCl6xzTjGQQPlgC91mURtuLcI57zrei2pMd
ziZZ28l7DDviss3SVC3PC5wZoLXbMSIFoB5WFJqNcOmOB86cQkLUaM/6NPnRyIjf
RD7zKaInv8cczYjoRBNI2eWFCkgqe3SMcRIf/2UiUndSPpquxHa01k9mDhW2b9Jo
I4CyvRNQRQ9aU2XQL17nqTc4fUf9SMjSRKF09R5U2ntx2vqrp2cTncYPU7k1+DAU
ZwrkbvXFWp5Jv4qo7N4wkkepe8c2o9CeA4ln6I+i3RGhQ0fiBrgjbmAWp37YqJCC
AZkB1BJrLZjs7Sz3cURZS+JaJ8OaqMcJjGj+4pdL8AFXZGCIpDSX4Q72tqpaniCq
k1l7eeaDOl8Zf4n47JsyqkOpUpGamfngytMV3jzmFwIKFILw/voK5ekSwfGCI851
Zn+ZmqnNIC59eJGnqs82K12FCH3Vv3oU5wJhmG5RYsJvHKCGRQKKsQG62DfJ8WmW
vJ+VGLBHJYxPMbHIJZwIDUNclKb/GikataDuuwv6JLbkky1tEUZVdl2bYbqXsuAk
DiEMMdmULhMv5eGNHgBGkiYoRONd+dDcQyGe0RfkZcfhgmDSfpDlFckjjCMtw+t7
6qSk95HERHMws1UZap6vi4ROec2guhnZKc2QjDoqElVU3cXBHEI1rLrfConarwwL
wraRtugT3/T7LoWVBvaniMLLM0kaA6WkHp3Trx72e6ZtzDDT/NU4ePSQxSJBSCoh
Z017HB5LSS56Sbm/RcEF3bWMTXqJa3Pu2u5/v5TZl8bsK3h00hvAxsxR3aGYJN9n
gSwxYe4igtJrYB2FJ+tAnrRo+tJC/KcDoTr5nIk8i2fo6za1BcLW/MIps0d0u7w0
wCGodYyX2S0sf36YgHvMtKh+fYneSJ8iNHbsbMIuXRnxwGcVjeqPs8eb0epXnfjI
qFgNDk5JuhBJYEzC39OiqxbPq8uY062aQ7q7WrNe2kfQBFrlZBKrsZsYjqIloYm1
BJMBtBVcZCTUVgeDJgN3qvuwvilEA1gZ8+bE5OXWtWQrzHgdaQezMibVIs2gl5kG
fW4mIigldzbh/9WJ642RB1xKc+S1zl96CUhJfInHFh9RZAYMnQJJLVA7wQJWms+i
rBvsqxBVXSkQG9aJ6B18uDYLYKIpcTxdpy1HOHfbFZGbQGqpOrt+9fQ5bzPcdwGx
OUPN4XlOFOxsdlOByq9uHsCIatf7fyq9mlNZ8nBptl+JaDm+VtWnXATJ4u5UwYol
5EZZAHQswO/CBl/6QByBTCURmJUtm9A6i5GTl8d5P1k71oxuMH3sKLTLdoBRPBrM
0C/f5Q0J0fePHQP6vsXbxaJzflkqoqq2vdfjEAEL4DkSvuxS1dF9SEmGNKKfL4FH
+cYs/vDvVz9xREcAKNdiudma3D2qPQwfnAuRoRHPGunE6vwoom4PgLkze0zduIy5
ZGcCMWQoBodG9lE7T46JcMKgIowF/sbX6vnVICzO5df6ImpYzCQns5a60+fJw7un
xW9ngHmlrLQJYEEWIvujcJV7hTwybEzovTfZtNbdTXEW3a5OwFvB9N6tFyLpHmom
gxNXsG9rCYUNxHJyml1ND7BUiDtbVfnqOL0um3m3i1gpkz8ecrE9E/QisX3JwCxf
dx1UWWL/54IcydB0eEVdbzh+464beaxKe4Q/rfOqlnSWrzrlbdeoSPRAV9vwmYYi
HjUzKEFc+UCffPuG+p+sc9DmYlLokrDnpCY7ElKixzcnd8/q6qSL6qOaZoshSrcs
wy2xB3QNV9MIW0Qy17MlFvMZZKJdNr00IPeJw/n8yzoz48NuxLP1+9OGKkPPr9pn
EK0QFi4uqstCvPaI7qKJg8z02vuWGCjkCizWmm3/35jsVK6sxkwFhXcWUdbK7b4e
tQUWruC5QDxwmfhLPARajfJ+Mq4IWwcvcnqA1ytOXNZZRwqJ/9Mqqw0RNPyOWuP9
fcdL1fmNUzJp+LKHQjM1bSgfGjrRW19lZtfcCjynyfJGVKbeyncDnclaMo21F4og
/MQ5Kj7H/nn6VHTlHFGlp4PHa6vNE86mkTYsFfyRUfp8wnH3rHTICkA5Su/C0pDZ
J7ExByCJKDMxUNglVdcnXEl+rtD50a3xSkm9neOv4F62qCXYqUDVxdHm6iqx63XX
DPHB0G7ppizMVumW7dovMcUTVXdS3Bv5Ypfp59HNPNYtFjfhbd4vePayyryF1R/J
sl7A9bnmEps4s1qN4dp7+FBEZdau39z33Moy01qIVSkx5JQBAKZj4QwbPca1cDIh
NMpTcFfsIAUNFfQyq6TqyUpMk5j6zCC0XE+9eNBGXrcDaz2h61M9QChWzR08eyFt
SEzzCs8vsPLG7Nwzi5BWu2vUFU9MOMpgusRfWyQx5REQ+D1RlXuc3IQppNXD+DkS
jTUb85K6awI2RiEP3SuuDBMQOue0IHZgDHOxNlnNP5qREVTmsUHO+8fGG5eIlZOd
cy79YgfRpGyT+ebQQ8o651xgFNIN1iwK1jf0F3mmbsxLnhoLJVON3ebVGh6W+/C/
vC5FIzA+oENBIn9m6XQLIlzDPrL9KIvF+9tWRI86FE0cFld3DQvu2XRYpr+ABJ3D
oBOVBq7NYG4NP6oeYkHBc0IPxsG7fBYueevDuw6qyzvcK12q7q1VvIWSr4IgJdov
YxR+IhthAlJx8rh0m9ReT1jvXHnWUMgyZaiOGbebXPsd7zbSHQ1mJVm5Bv2/6bRP
Gcvp49tYsqkvwgecSskGNujlpa12V5lqUpcGOAXW0AspjltXCPyEmNMn5nTJ5+0U
0ru8No9wVqBO328YKIvd9e8IC9pOYa2ipteNkV7KxAusVDKHjwO2CkUA+uUpGChd
Y2TJNo0+0Avqrq/r9flAJTP7KYPAFp63cbwMgPe7TNnnKEtB5pTtgbefQ/qqR5O+
2GChzUvKYDHHTCQIENG9oaO53rS/jOI9wmQtZmt71QxFO4XLY1BU/6sEZluQQdvJ
SG82r2ZchVwklf9In7kBZpnJ5kJe5hFDR5Cq+0uuD548LnyHxHUitKD1FmSZQnwx
28SMXFoLny728TR7gv1+twZVqAJphCttE4OKGThg7YBzruZ4bxd8tLgN7cf84SRA
moqd7bgorEJo8pDwWcx+61A32yduLuLv9bIliGr7f5bullvK3OvrEpTtYPjiUOjd
L0zsqBc0Q+Kn25Nx9QkYc7Ikbmvr12QS/Iq7FWpSUMqGz3jZ90r5qZvSiBUIBCiw
Y9R/Wg7DmANeIYbUUVf/z6FddXU7NtqM/qS0uxClF5HTrZt31qAmL/xWGqEXB8gT
wit0RGDt2CaExtxxRugN7WiliPHDKdVZRyaJtvkg4oJwey6IM88O1ZUTLTu2oUml
1cHcRuPQ9D1eEC1IOWOPzFMAr6SBmTiUMuutzIbyz/vkYw/nkDOim25/eLGu1FEJ
/dZEosF2dLAw2mJcMPAobavowbRCwumO9zgiK9vO1tk4v1MfqTp2L6RHwYTg5Zz6
MWUSDdBLH7yz4O1iQg2CJ4mWs+IOSV9ddzmCMVXdl0EE3m3HNGAbzsQr2xo0lcEB
XbBlJQHXA1Kgd3XMcAZsexzm/GpDub7uy9ytVyKL1laSDvWJTHIS4RBxJDDRpZy7
Nb9Tn2irKnrz3vEqxd1LFw73JWQ40x9cxIc5BOwltK5YkSBykDQ2kQk6OF7RSRa7
d81qKJNR4h0gk0NuoGNKNdWZuJU4M9XxSf766w8wckPKlcHtRs4QuKoilMFUob5W
ABa2FjXW8vV/yiroWsJlkLbni7T5FMzRthiU9UZmelS6iSW+8gGH8m/TvIOQjj+r
jg2vsyrf2t32srESpSJlIt7fekKu/PtYe9IOL2BXJwiDX2MFza2AEftGOQBEBHAh
0JFP9tWh7gcpVIk0K29JZvGrKkeDv4JkghfEUu6zdNTNejHvb/5ZwQyHuC6N05Ez
4DspXfAb+ym5SEiHq54EdA2KdrIKtXvRzvmxm7oU4JxL5yZ5ASw6hf8p+xO0ozLp
iM3vD5a1a/J4SOuhzT1PG2Wn1add+nWGpE1CXtYS1YzWkloE3RnWqWBjcSfh3AVd
uxqVHLkXSV4gdOYu33pqpLdsBlRgpvuCwzQU3HKIfJiwnh26JeV9gfvtb9rMjky4
b736o2MvmpJniWBynITr7lmeBOsz5R1pi2E+Fb4jCtnDXkdXNlDXrTvMH9QHU6HY
O9X5ZVizt/BCYeJJxvtgNYR+Z6pY5cmxfkFEKO4JYrm2A8TOlY4zHZm7UbfVskTZ
8SO2uFUacrRMojsGS3zdGIDnLxGSvsaGpwIUqq/AoO8bLvU6QCkBOK4AVNlvE1fr
xx3r85v/Ls9dhcBlqDfpyBSGi00kW8VQAKxDSIIqcFwL9PLGsJ9TXBhHyGqG5dLg
X+/1ZzWzq4es8Kuws4cAyHPAa8luTLgsYfw3RolZka8ES4+jaRtMR3QHZ6IduMM3
4t0b1+1jHZHazosc5wXhnrQ8aiatvaZZnBJKAWvdphMDFZeohFRogL+T10DLggBh
1WvEkXSi77GCf63uUDOsw7D5b3G2DVZQQgOOmForYNaQAVwNbtxKv7Fi0WMh22w8
/rU7qPRXTkU8UJIrk80nwE/5tV6gziFWALtFXG4+Rh8s4zln+EdGvYtG/OutUGaF
ZCrW0RNjSwWk5EMCDnNaz2eaV9uW52Sgdvd+SfTResH0BY81ISqgU3KHitkJbmaF
IuBqc/ron4h+4hCxWXCINi5Xc4tn1jngZeYiibuSpD0Kf5suweKPTl7qVbO3Zv8v
mVa3NWhQKxzBl2dhnniAjy+yPInd4MAUiY6ff7+kICUhLGsGYtCzsmOK4Hpi/xIp
IIWsVcVTRzRM7/Te+XyXi35VDecxZZwJ6h3SkiMmI8IY1xJ/KWRtzXVbgnN+j+oF
rWT7hAH59MX2Q11cDM8o+OuOAB3GeTmw/XfLyMDPffiYfFuqtxAFEOVLF7OS1xv1
9U70Muqhpu/p/nfYIWasItL0lBiLCnFGQGcly/qJHdmvWJET660ghw+oY3DDmp24
OOWN9ykw6LezPB1f2alUknlDcryQw+08egAWBu04bsCgDQOo5Y2D9sBV806JeLBi
dyffTPgnJtbH50H73dsYAuFqPjmThNIZzWNPn74VYS2Zo1GZaW+dS5kr60tQEslL
E6R9qP/6yREtF5c2LyaNC92uS1B9Ls/S5YoWH34r6Gnuf9W7hfY6Sgk+ZW5R90y4
aexGBg6FPRXwwooX4kUb07SU8LbRBpgeUi67XdO4PdpXc+Y4HFErFbTvDEGhiRkW
uJRc8Vm2Vp+8lMe3TVHSQLvElAsw0lRuYFP6Z0+Fd6PKYlQx5QIz/QpN16Olm3n9
VpFTwo/nOxExmPXyUOx1jeAObREnXQOpcvGNmZcXjQEIX89YLfPxg1ZyP8mpVxTO
TiAMT8eMujNZLqKcQZb8vbrgsBwRrlq0UHL2dWrPH5TSusUId4qkp8vPvkaZvxuf
6ODjzE6vSpPZQYB7dhNzwMgJ165iIXk17NLVO1yxQm07l/rdZUCBUYoLfECaBVol
06nah7bFM3lagCzFNXsMkemkKwr2efRrfblq9lys2NTsWBxHknDJcw59KxwLPgfl
Nfd91zjeazSQnC39fZktl4uxxYmfZGh68egZpkILnne7LFGQXAS7Zu4eay5LuWN7
sFUQ49qGBZjiQItjJPA9vduhaNm0sZpUtZTUaxZUa8e8SmuSmP+2oKK6+KIfiIWg
jT4fVKMJRKXCW6jYlZVBAmyXLuJRBR61v8OxA6y36j3tT0vghJZ2sIKlDruIF1Px
fDtgGtxkF9ki5XcbikyrHMR8alsgzuGxyPYhZNe1WaUwFS6Hl540/FQuxpMXn/M5
G5vUdU25EsKeBn/IdE68tF/+G9V6xDqGO+XjZK1eptMG6oRcwmFn7yBM3ld8b6LQ
yIPg869WWWkaUw+8FIJ+tmu7rAWs1HRTz5jeTjlhosQ09cW9ZjV0+rxGSDLnbcHS
weRhzeY+sTj+Nvl/gjuidiG17cBiH5Y1TGFDNqsFbFr4TR1DcC0Bm+QKNI/1RehP
jOGbZOAWW23FcOCmXs3JvMnT2p8P3hlxxfdyiVYBPv9/dmvAsMOgijsU+8gqYUFO
Um2wsG3NgLslK4q3o8Y6l8Wn/xLOLeLhclg5db//mlEZbqBUyHDAk8OvaK5PNywk
9nvNx3AL0DBtePB2pAcuqcmzqyIrbz9f13ied6gPRZRATTKlXMJVRgWrWeh91J+4
5OvEFJgyhqxXjhajNsC1XjimQEo5WO1U9KppY3t32F4lTm3Nw3FMuuVjO73lCY2l
Y7pV48lbWxXA2wBv04CdIxVRP0+v6vfTlNwS2XJruBqYHpoEacnFDl122WEJ2ESl
MF4WZruGWphhP+A/GwLQU2dUVgK5iYl8Ev5WIzLUmTfbObW64AEG9h2klWLZS2Zl
och80DJfHihq8kcy3Ku9wO796A1m0N2qH9i7EPSi+zXtN/snBPCVFPYIjpnkqIf8
fJqPM26AnYXw+959BTZHWyJ1gpzNMtRMGSkpzUPaIMK7olrvCCSsrxizRF1TFj26
Rh7PB7rxD6FzP9XhG+5jH4AKo01LH5S2hdnunBX8XFC2ezCWw4QWxdHaMOvNRwG6
zjbXhI/Mp/YVHOozIRG1i78bFfKhRDXT5d986dWtX7gBp5Qh0LvY3HiPhr3lZvxN
FmkOpKjfNLitg1j9WVWlXPN9U5qe7Gnf0+gelyvA+GcpMQeAtRe94RhX1BOBqlSa
7vxXaDAdel07NZpyHmZgQKZHGwzJyxIdIESnhU9gpgMSUv8IhZMJSCPFCNwJ1IDk
wFcNlf6P5Mg2JILo1rUQF68QMB8AvXavyXXe00WssungnAjMLg2szX72YaubyMRy
KtW2HjPetO6EtOgCdNW9M/ax3CbUVaWKRUuwfG/2TnQwGOZLVAT7JAeP3e+oeUEM
VV8YrPb49bINzSfxusKhuK4MlMWm45dTYKoDOJ2j3gfOqpIcdEEDjB5zGJXUgRu5
Xh7O1jAXVIXAjcO2wQkcm2LFusoQxCDcg4t15kZOS3McBXOFZkthYqfa0QkBnwbG
c7iz8q4326SKvIWIKazUamh6tl2XnEpzERujjVH8fowWJBzLzBIYvbtl9k6YHBVn
QYeX4EAx20tcw4sF8dArqm8ns6VJOgCZvgirS/78MkhnfvojsiKCnI02CQeRb566
Cv2WzfIoN0YjpGHIX+AmvUpuL0EYKOXIjfIyb63Q6Z7fzK2SXbc5cgftNDXMs45V
SgNTyXRySkAX9/5piGLxhwhibB5P4TQvT7amucdG73f5wpTB9/N9hnnhqaHNfvMX
saY/gAxeaRMJgPcslwG5x9JXSiI07clhDpgIKjfsyTzzxjkv7tsjANbUQ0o1Oe1Z
Vt6MXPlkaeD8HnIOJXz84k8+NFxgavtxH4OxFGREhYlgz5e9+gQwbju3TMkBPgZL
rGRV9tO7P13OoEJZkZiDpJHUIBFgbHdtf0a9SQ54m6pHWtJc2O6QlBSFPf02Q6zO
AaETt8/uTUAVLIu+dvZiNFNkzpv8eijddNiHPp3N/8Uq35myx0qkvWTLCz6Y9y5q
Vo0ksEbUP1BgqN+WiN1YV8d0m4WAcUtNUGG4ADCZSdUjtIavrOGkXc9S8eF0QykF
e0EqxWWe1aleMqYZvgKCvxH7cLzM9bT5kMap3vzB+BWg3RKKSnH76EXtLKXuqUv+
s6ZPqFI8pv3AMD09/UaQe9lg1o9UswZLcquFJI6tPg8elHQeDyyk0MJbrt/Xuv6R
9r6WNszYIPg5jVUi++Xq3bW+KJi3YmCuA1B8G8CkwjwAQFlgeXaYRvM7JT7luFgD
VdNXSKAhVPOMm/OSxTuyRB5aVi8ETPSeJdfh7M7TwV+UXv/nMbzHRmTry8/tPaXA
EawSotbVxE6FezqW920FwZKnn0MJY6PLi+FekG0UKbAWIjZ7kVWuC+nDkSGoC6Yb
a8xU29PJpc+9+wsUO03zRqAqBVzkmNkAtRlTy86oCry7JghJwOEvAHJGiuE7my8g
RV2dFRJoZQNHdTGi2XmzfxM9fUpDKJuhfXCUvNaCKFzWrYFxgN6IGcEqJsavCwqz
fLHWmc9golhoCe9hjTnnEJtCgKYtmDgp2B4SLjevVhDVRgSxmvjN//pGPHRIUawV
nAn9KS1O7JQCF1uX1ZnFsOmLq8wkpSZmUZfnOMb4mHTGiSsZUubJmDz9LDsPWxdZ
+Yll1oyTv6TiTkkG36pUWRg44xlWMNLQ/6Cx5W8LKuVMoKKOCdqFi2igXEofJcWd
8ycL6NsA5h2K3dg6u6nirsg7yfVDwUe82hMFl5ya6NjKfuWv1g5+H1vpAfRQYziN
98Ro5di7LVhihKNle+rCev0pZideOtdTJ/QSpGwlIm9z6DodmVh8rRO/Ip+gL1gI
WjDkU8iaixYjVZMKGnCl97uK31HOgK6tz3FL7ilqtKBSNFIC/sJ3YsqFrbQbR7ro
T5sVN8mceh8RynXJQl1oxklkbEfTshbMIhEvapQRWmtBREZHpgRuePFU2Kspqb/t
o+JwNrVjN2FLdQ5T/dJKx24+YnF/uLzguoFnq1Sr/pAUdcfE1dxR4EMaVBhaFGKP
rWdQmF+c0IEiNOeMv5VUzIEwBFM3MfTnUeLyQVfnsCib6Tu8SaHGvIaPHCYx0/0t
f19HrxXBumC54toOWvQI+nYmlhKlyDF5Ezu86+CdzKSUxDSY9eAOtAXtLnQxJlMq
bbuA7a90lFry1W+B9bcUx8IgUYytE6K5oagzCyuDmWrK7c/TzZRdwDmeTN09o0/g
qe9U/XgXwLkHPlJFQUZm+VkDtV0o9UKE5cTqjCV7caC996lyNII230mpCzjKCdoP
77m7vbH4mH2aSJu0P/mF3igrRAXgBk+1KxmvtGkp8EgiAarkQ+FzbqJC+npTAWne
TFw6x0YMi6XZS9tUHz0jQ7fUgqa7XD7BuozudFauo1yGRc7Q0bY3YbQ9aEopxSsy
HmVLmI2s/74JAYP3GeTuveWPDdEgu1FxYqAjhArggwxMcv1/P2D+7kMhsP3LMBGM
lUIwQwDp7IJSgHIBNP6I1KeabkOgJHdMc94BcADo+gi9X+BPGVr2yakFs8Ha3x18
0eeIdUbIyqrq43cg1SJsdtXkXDwbIlwHIN7JhCg1KKSVvCuqv7eukzs0O20+OsXk
RlsB7NEIA249UhaXqexgG6mFanE6Dtb4/Acff0m7Q0G1+moEf8x/aRQNPPImOktN
rAdGnwvtOj4pRKpEOIm58IEnsvNzm6kbFwHLjCu+SaQLs6WYE2g2jN+ZDThx4pfp
/a2+MBNL9Ksq8mKnSAKqix2Dx8wj0wq0kywjqGPjC1Ob7RKG3bVuXDvA3W9JXEGC
u0kubgWxwYr6bJpEyFSSNx1xN0mBZ6V3TlzLwE2s0ncdv08V++60/4AjIrGMChqW
bZjs2bpaG8nU4KTEiYi2+HZyioRuMRJCAc1JV8qWmiJjakMKZHAYgA1VpEGhXCmd
U8iWndFtNpp1tWeO6NspNLSMcOJ5QJ/RLfT8kl8SkxSS+UvmMafKvs6LiegsFHy7
EEk4FsxSO02LH0eASnj5nYIsTzQge/N59XHRKcMAFzCElcIyldf6Bn9AMTGlYYEm
+j6ryV2V65YFjAxr1tOEXhb1l6FG1wh2AXQjL7GMaHywttkBU2aQ7V18QDqsmGvx
MDeG4aCUJ3kCAFqzgOZSrEAx7xwMZNdJeK2DTmtANOPpKqNZfGBZU2XZjKKKj//8
oDtR66y9/P9oSbpaK4ENmQnyTKwQ3QZnuk1DLKqTy+Tyc1Kkf+sf0umEmh3/9/Nj
j/bhwJiT5n/62xrwkk+O4DsOywaTIsOHsYhsPN57RUK1s8bwSEHKj3seYwnoYpQ/
/7H5wiYctSlmS8+E0r38R4Mg22kkiOylhf/3ajeBDPWFBjd9AMA+rqvGNj2tT6CJ
hFfX+vaFx+11s+G933Aq2MMJz68V+fjGzB6jBCi35+HIsrZJ69we0nFUKHFOgpsU
jXvgMu33oSkdAz5pRyKlxP9zXm7Fat7HnCHw8W1OSW4kSNcm/tuTgM6F01OvhP04
Z3jmofysWmNrF49fI00TveuFhMSd08T5T8npJkwiRKL4iJw5/8xfX/0T0IsK9dV2
chb95t9uwwT9gAmJnen0ddbdct3ytPwdjDVpSp3sGbrmgb045KPtN7EWINygJWsC
/02vfldITIijOlsRBukLrUGNFZk3huEDJqq0D2EMZ2IYrspwwFtZ8qcdsBUtMMlo
p1f08MZ8LSyfMXrpgwXFR498f1hDBc+GcHfTQNi6mN77QKCZPULPzIHYhttPTHj1
eUeX4XVjUIwItGUKZYH8FRq23tl41gSTq3glXWuAFPYYVpDkbKBD0lQL+9mtHi7g
4k/iK4yIikIeZycN0i/TRpuZMTl2NNBmYsJRvtW6xPOmi4HYB88d9oGGkjzGJgPm
QridX6KMRwgLOpLMa3e988UNzFnhOr0PTfiqJBdR41NhUWe2wPROCVBQQh1AzGLf
ODJADkHpZBZ7RykuDN8q4cAAqfY+cXAFpVR2/mI8CM3OrJKYelQ/CGrrjHJQ+vVd
zfo7W+f9H5DH9cq0v2aX0rUixiT+/7tGpWVbn0aPmFZ+yN7RfYftsGZRAcaRec3V
eHXPsf6QPMq/wLzbqD++KOdtM4V0emuDrfiparNaEyIizew3TynaPhBOGB/ixrUx
T/shq8Cu8dFt+t6+7lGpakuc4JqdmwHpym27jbWU5VVtEKUr9rWKbfI+jBbankp9
tjVZKPLanxDtU8a4fUbh5qSQHBr9GMiNuy/xecdYn2jZOojmuLHinvemwptATXA+
BobcDDqLG/mcFliegkxnxALbT1KBtmMkZLHvyqEBBjQ0kkLMLDZ7HyDJ/LVUWQJw
viiRzA1snnmEIZaOIVhq+Zy5IDTc7Tquuk9zb0hLXYUn/U1UzzocgOLiAPwVfPNE
KlKS82DJbez8rweKD76ZN9EyxM5d+gdCSHOapBilCk4z6MLzh265A6SjoHSRwSsT
sbo6FY2Wb7WtgptSqhkXD0lO+9R4Zc3c0XSUHyGmCvhhJbP9CpW/eSjve+5pbXJr
2Qgq3P4izXJZbZF+e+6Aisj3q0cRy9n1Ij6gd059brrla8S2nmtqQqkZCSlor3jI
BVlYRvnFNGBZ7UkZbvSHTnwsVjddyuemfronVov0u2xulk7wQrr4PojBUESpw4D4
kTRDEuvoRQ67rHAJT56BEWNh99KrY4CqGrPSFDJhwX47o5XzHeoR3iNtfY4lr6fE
DWxYcfWRspG42xExMe4r2KYzFdXxHzwnxx6pDhkleidECKJg8/pi7vRoc1kGVPuA
8L3SDolfaf+tc+wnQPRmqJoNqBo8SlquYps30VY13nfhhA+IrkrJJgKGOjNFDz/T
lX4B4qhBGYCsIIGLERN+/sLKd/6qMH6HIPvPOVl021Cg2unZLRgcDFUy3ss/AgL/
CUPXJUbWM5i9LRXpkQa359/l71NvYhH9FTIg1XKCgT3jK92NqM1uh6ZOP5uMs6n+
+x54VzZu0hJyPcFXwBAWd+kWwo08vbRGuOhurKdxJHpBWQehRa2ZvmCzrpwMzIrg
ieODzsBcAoEHdf/+L2onAtdhW5kHMc9eHpypRPrNNHrtX4/4iOD7WYAKIdvX/OZR
M4iJEeiCl7F6ia8K/y3UdtaROdtQ8i7EsHHgUM064EqbVc2KRTP1thm4RyZvPYud
QgncqrMsBoRjX3ML+SeO3vDDETIUzFoF5SXWUlrPmjFxbW/PfJ8LZOcrYtRFZmp8
ZkdlB9pzRTtxIHVe2w2dDxC5ZNryavP8aPGyebANPJqbTU0WGKaTYMQPTpBt2doY
kRbbNRopgbm8u7M0QIgSaA==
//pragma protect end_data_block
//pragma protect digest_block
nIa4PLA9YAf2doHHgn6bRNX2dwo=
//pragma protect end_digest_block
//pragma protect end_protected

`endif // GUARD_SVT_AHB_MASTER_AGENT_SV

