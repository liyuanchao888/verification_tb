
`ifndef GUARD_SVT_AXI_SLAVE_TRANSACTION_SV
`define GUARD_SVT_AXI_SLAVE_TRANSACTION_SV

`include "svt_axi_defines.svi"
/**
    The slave transaction class extends from the AXI transaction base class
    svt_axi_transaction. The slave transaction class contains the constraints
    for slave specific members in the base transaction class.
    svt_axi_slave_transaction is used for specifying slave response to the
    slave component. In addition to this, at the end of each transaction on the
    AXI port, the slave VIP component provides object of type
    svt_axi_slave_transaction from its analysis ports, in active and passive
    mode.
 */

typedef class svt_axi_port_configuration;

class svt_axi_slave_transaction extends svt_axi_transaction;
 
  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  `ifdef SVT_VMM_TECHNOLOGY
    local static vmm_log shared_log = new("svt_axi_slave_transaction", "class" );
  `endif

  rand coherent_resp_type_enum coh_rresp_tmp;

  `ifdef INCA
  local rand svt_axi_port_configuration::axi_interface_type_enum slave_interface_type;
  local rand coherent_xact_type_enum slave_coherent_xact_type;
  local rand xact_type_enum slave_xact_type;
  `endif
 
  // ****************************************************************************
  // Constraints
  // ****************************************************************************
    
    `protected
27Kd:^PD^V4G:#D9E+dOGY_^:#Y7=>ba3a#XN1C(5U(T-Jb?9fS45)E>a@H:Ig:2
dE)MRJIH&7_G0$
`endprotected

//vcs_vip_protect
`protected
M4#U[VDGb?0SJUH-OT530SU,7Y=P;RE-Mg]N+:\^XBC>Q(82.7#^&(>:G]&G<)U4
f^\<\K3/ae:;&JO8+0GAS-=Jg_L?2IX?MKIV.PIYN.I>RUPcSPL[079D#:1]JY_a
&HdD@QQT1HKaGSJ>TB#:9U&Sa+=RR+H#&5B\@A#R-0(9(eE9IIC@NINJ.)c]V4aK
4<&^ENcQ;;+NWG#e^UU#95S4WK:OG,J+aG\edV-+f<S)=)CBJ-)DAV/VLL><;S^f
:gPTAH4UGIAZc+=(ATE9;5PT#.NHUD,GA^=Pb9WP>LK324aZ9E5A>_\-E]g[4/cG
[^-4?[=KAUR8PMBG4=egd\SL,@]];IQQI@_\4\V3DE-g2K#:?[G9NP8?f=(MbKV]
;&89@#SeA\L_&(OWV(bd1OCI[=I<5#3G-Aa5[(QIO?]0FcHGf[d<:Q#U1O>Eg(K,
:aZ)M>_Z7ZW58WFV(cYAg&Zc-9SHS3.51#.8W#=U^JB,>L?][7Eb3/]O]cC\4?K=
ZVe0W(A)gY3LM:NF1b/4Y8[aT8>]^B=G4Q2M58CP^U^E@TL:0[9:6^&I.<QRdR>G
5_&,ZNI:?BDcc4))OT_MQT=aSb^e5T<U;809H\a-NS-U_=[c=H1^[T4UJR3LfBCJ
g-eeRT7ObOP?L;WbES,[ZdI^(GT^R79=T#?feE:S@/9bM.L[W?_BcN.Y8bQKS5GR
Jf(AH@3;Y1K+@dK4-S?K/?CPUIO<X4(OU7#7PfZBeA3.@/>57/H\E]A4PALK#\DR
?O?L8W-YV:ER]:O3.\??V5W_e4d():TeTF7?=#P(A,L&a0;V.cC#J3UWPWdcDZgd
/)S)>110653&DZUZFZ0WWUU45<<fKVV<F9:EV#R0UT[>dKT]QDNV<fG)TO;+T^+4
,(H@A1?T(@I]FS7b;XcF1PWFd?>DdM>6_g[<O\LY2GZZ6^FD=#WUbIAH#CFF2H>3
#15dI36Y-AB8e-6PN+?0-L:5H@Z3DPY-6O[a-XH(P;LIZg^YU2afP:&905IR@[(e
#US10U6bfc+Xb40AT_18Y<F/[3SE^9@[5K.,LdFI-];XSeU+UJ?CT?fX@U:c@4HP
d,:.<8)2cT58M>aVR0\8cG/G:7.)G3c86g/T9)/KT5YaC@SV4IgPR<3Ng0ZY)U:S
2S(7(LXDIWa:fV0K6SeFV<Z^N)da0<D9ZS.fX>f>AE^#Qg)?bOR5>X5#dX4M/6I0
8eR+P-XMUK&?C+]WM;f<=BQ+<KOa^^[=8NI6^&311Z5<[>A1ET3Z\P\;7=57SO27
.4M.<Q+@G/@D0;cIQ(YHNFFJPLcN>AOIcX]AMNg^/\5BS+EJ0/;G3@TNN#dg;H[Q
a[<+PRH4_I6\^(5CM1d@EA.PMOEK7[YT<[\VeZECge-I@,=YXJR1M>?AIET?9d>J
L&&.NP8BC[J.babJ(eHB\cAM<ZUM_<5FK@I:b./52T;d60@,]/MH@O<.0Q2GW)8J
ENG27d>H.LO<W8\9<a2(RK4OE[I=+)PCAJc=JG,:9P[&Y=3Q:#13e;&S@JXC8L,G
^5fHDg0[@U(H365)EW[_6,RSGbbfMT+E#4[)B#QW)T1)<->YFTJ@YF^L,gaC/HeC
)Y;MY35RWXRPF?>O8eE7/]KR]QdPQT:G),C()Bf2MV/1\E#4JQfM>6WWPd._?T<X
6_,Q,UcDQ=8F-:9DTN2A_&=4#b0;UHQ);fEIBYNTT_NOA2JAKON(^?IXWV?PbT5/
(gP5gWNR_(KGQEde+gYN/B/69#771=Yd7=9^?7\)g-EEL[UZf:UK0]V&>LLEGO@.
S3)G9c:E=T+6J0,?K7dHGSOKJ+Cf(^J4AP1JS1]\ScR0M-&_/fe1Dc#5-F-?8,#M
[T&,?C.J&X@554[+RKHcCL,?J3UZ>c:[He(\AN8])dc;8T&.[5[eWe,8TdR\/L^N
dKW=W=Y3b]Dg@Q1HgXb/B]&79^a9;RE(F4Z,;<^O[64DeAXPI+/EXDJSXO8YICI#
[M04>?D5f@6R)M5Z^@Q]7)BHJ95<9TIWIB723>,\(\OO32)VJQ/a/S2E<6\UDD_L
W>e11Z?c9WR;d5H?V9TdacNCBC.d\_,F9XZ+)B1I)U(_I3Vc))2#/F-:_)-MSN?R
;5CfCYHK#NF0Zg&?J:-,d]fT.NN^fWeeHSPY73+__NEQ-_R:TGQ>6I&b^[;fB72)
IE<91=&L-J7<A)B+L.P]CJ+:9610JB>XAgH4Ya](O1\9D3XL^WR8V#W#dWGXRAGX
VeLH2g-\^IJA4&#84ca0DbEb.DMBF\+gX1=SKcg670_2FeN;5Q?TRV31Td>=e05:
PU)UBO[Y9U1RHSXgSX#Y_./Y;0:X=S,X\Q?E:UK?GE/T;(M<#F[c)<Q>797d)@Tb
e>G0&dJW[bN\@a36&,[D>d-Q.YORZXMKY1XBS5IX?dOQ241-86c8a/IT^-E:b-U.
VK3(a(UgU([2b5(9I,P<6?=426.]G?e^.0H[Lbd2EYG-U)DMKb+PaQg<c1^E@Sd=
))4Y:R\-37U62J#VScg<W-d:bbg6:7ZJ8S6g(/@H]3@MYX#O>:D74-EL&7<K-5KM
;\^Fb)R[_Z@U)44f3#RJCbK7>e<\C],B^?VI4JJKMTU?1T_2LH_(a[JSeg4ZWJ2b
]H+F/<dK<5?#\X.WA?,aR78^TP2PeX[O+ABf?\:9TKL7eFTJUI>)28^gMbS<X)IW
=>PWbM4BC;5?CbWZ/YcCCZQOZ(5Z0A4f-A-;=2-4#K:3[@;a_/B=-D+E0PL(0)]a
e@Qd<,fA,CM-_X;Cg(A,f58/IBULZWMCF-<Ye@Q/[L>-b7?aFJ&aE;OcG2&+7.GZ
<c<IK(]KY/d0gc<OQ=9L^^[7.3H(V;C&0]<PFS1MMNPE>LVNGYJHZ#2[N1JaS8?7
4adVG01U^;&X.4)Pce)5O3-/C0YK[XP&4K?Uc)\MZ+,SaI5QRTN9W/QVZTcL9UF8
LKCL3K_bU:EA_BM2d^I3P.4K#W87c\P;=?TG^M429_/D&KD^E\5dUU4>-@((L.;3
3T-E1[[GCZ@JK.&&.M[eLOUJ^ab+969]ME.C.fL2B5Z#6B:/)HCd5,d4F5TWfNJ5
OXa^/D]]@B9&KUB6F92\+CCXKPRcT-N6?<U\0OfDO.S:af\BF=PU_Y@g^38I]S-7
SIZU[7[)GR@8b@a>)G<cecJ^+2GaaJQR#g72HAO/K1?C()ObR8M-L-R(8[NCF]M)
38=\D#^\Je9#88]\5BF/FD1W&R48#2C)F8N?NL[g1LGbO9GY<B5QM^-:bLN<D+V0
<.XAKgbPdTM<X^VP+O6HA8JOLQ5gB,_;,ISG+8MeAF3#SC\S0eGO8?[-X=K)#LGB
KR(PMT]49(?)9dK(57#\G_@G.Y=SY_:;E[gHVa<Q-EFJ>9()PX:ZVc;<<+]F]fXO
)OKf4B:.:?1aH,#-246VIK.=b/g0]dOV4LeDU<;/Idg\XLSMT<I,MUDW^):Be:<N
_WYXP/B0fOZU/X6H\&TJJG<./Mb;][?0,[8;2#U(=>W)G]Ie0U#?V(T:E:IYacIB
7/+U#R[UB62EC@5TaB3:PW.F>-R&+RH\/9DM:@)(bY4(AaLYUNDT.LL_H5Tf1f-U
Z-2ZBW,\U6-0cER8Ad#G>:R]<#LFQ,L.5M/NZY&=C@D2c]AUH6^b2D[>F>J8H01Z
/RXHd0RSHQX.Z;<Vf&;M,XY_+;B9f3YZ#SS]gagP::5#R)+SdNAU@R_Q/8;Y5N7;
L=UG(5PLNUSA[Q88TD1gbdc&(YQT1UKESQ[/7RQG2KP;L?SPb^-U(a0-aQ0Q_CZX
Fg4T[F@\EJ6K\;eQPd98UQ,99A#T)AI7I]E/YYBR2Hb>GOadFM.\34IMUSg_1+Pa
gAPVLcG(EZET-(f(>^+701T=,_4>4/[YdL]d14>^1gMY@QK2#,.F_Gf/f(AZ0[?N
4cg;4dGV:S?Ydd.L0@R]&OcU;M.=2ZGOL0[E=OXB5M=UaBE7E&bI5D+S,abAZ>_V
6ZdH:QKdV1bBV,fbCE27#faDOP<?0P&Q6K8G]^7?(1,WTMS1>4_@FZ=9_H0KMegd
2)OXMBQH-FP,9.TG+@-Q#YCJd:41E4N6]&.BY3T5Fd]X5+fE(D.bLaKTSb0faOT5
T]dF7Za_T;QV8aJ-<W@d3?XK[YPBBA6[-G#bUDF#g;aQ,IePY9b&J3R4/JJfK7XV
4#R2I>@Z+f;+:e5O9)_Z7F&>#Ra_/9Gd2:495:DZ<9ffA7NI-;V/M6[MRTb^KYI>
8FTO&SLYB,NR7?.()&\EQ8T?0G9c@#.0H<Wg@dH^L@fdV],X<9#N,cJA,3P..efL
\c\gQ&:LgcReRgVYV<\Q>E7+O3d<T-Q^a93EUG/8d(YRf0-.M+7C78FXKX#a4Y_&
.RQGD1EX4[I^>D5(\@DCCPN&7&J/LC=8\V-([)=,a1PA>C57c(AS@5#N1Yf#G=L^
-+<T&<(>>WGb.QHM[?6Q71#^UE0Q(EX/H1-D(Agd&,T+^Y-QYKXK9WP,:PXa<7I(
W6=cHXfB,806a+=TM^U9-2VRf]b3HS4G9MIfKBUE\4g=\I/_EPE=bX>f]Pc4Q,5J
63K1OfO_IFP-LC==XM,=AIbgf>Lf/+P3EY7QAP/RN1,]9=HEH,Gc,,-b[C4Ye(gK
;FNgA.CU[MMD_30UORUW47H6U#0Y)gXP>I?98>H]8aB?F;G<a#DWY8\QU9X80E97
J6IA\=Ad3G96<b7<WPN&C9I5a.LUeb\M^Wa-1bO\G?aFa76IG14YgTS2.<cNWdMV
c0(^U7^\c8U0FRVPGZAe\>/Z^d;F;EM#[XL#a6BafT5:^Xbd6Z=3U<G.QL<E#R+5
@6G&34JB8a/f(O^TYJ&CDEOGEB1(>(-/;)b+eSdQU3gTXWEL_2dFHZ:L)&-P<GI9
83f1X^KgR^61[331Z;=Wc6\)42N^DN2/@V85H(;8-^RTQ#XgfOe]bRfbH+Y[9[^P
.M#0<=Q2>[P/Z;B>-@V4:43@12Pdf1@DK-TCf\4VZ]JSQ^7GK[6PE[M+A:=P@A@K
<L5^2:.a#P].D]H3<Ka09L@Jd,(eYB,bb,d6:f_]d<]/5@[9HT8QVI(&K<7(<Be?
A3Q5R[Ie1dagCK_BPN2G?9)&QWSF(1_NJTARN2B74^1([LQ6J6/(Sb<MLd+L\bP5
[L>PYNg5M)/DfJ:(SFB95d.Q>9L7X[PC(@#PdRHM1UO:KB&X(JD[Y0<Hb0T7KGQH
RB-5&B(B3R8c(f>,b#cK0+W\5NWf7aSZYTYLO<ZZQI@7)TeCGFQNbL83A/QE0]NZ
be7M)f&65ZH7PLL;(@E6Be03_S<]EdS<JA.Z^dN8SFc-J_)P#[1;\Ng>JR)=P.Qe
VH+8g[PT?YJV_&&0<XH)Y.<(D8JG4O)5?5,K:+_MA9+G67\H1;K\22GVJX:I.e62
J:D_3HS&4Z99ZX0WF(]DQTLH?(>:(@Y5HKO3UKH=SZRWTOM&?/^-<CeI2aR[Q+.V
SGJLXG9X0D?AD1dEJC&cI9-H=>,@<bA#6a>-Z833/K51CUc]Fg?DD=HCX^1(BPVe
RZM2\H>TS3=VYLK<OdRA;H@52,T2P4Bg397\8;Hf=W>@4R+U;>b.[ZGRK>=,\(g=
?aY08JWIEG\=4G9a[eG\J\a5_0FJ#dd]DI-Q3N2QH^b4.WeW.@X(,IT[X]4:AHdL
-[81-)7U].[0@bJ5_F_EFC6F2/>M_dGRVXT13Jd]:X?OXKS^E7MY,V3Uea[V7O8^
0[6&@U4O9N&430?U\:D>_></W.fBT^f2#b_SgJ--H/FGOZG(]TQKaG#3LPOW<Z>#
E8#IEfXMLVI=XdDB4N3E:LX()Cf+W4a4=.U8M>a+[LZD1C51Z]U,=?d^J&Z2W600
U1b_5JBfZU#A&:.W/6FcOM/Ud],P/6Pf()X1_M3&)I&bBbAcKFaKTX<JG&[R,;R?
?#^\NO+TD_eQO0P/S/>I4M<gSQ^Rb),Q<a,N5Pe&VIfRV]<;8Df,CEZaTf5(c#We
Q]6eG]bfLI<C?D=d3U3QT]_SFWU5TW+6D[.)BQQM#S-8.>:KG-4\N80J6bZI@5LU
O/2,@\KO)fI^\]0KZ^5cE^4NeM8&acEg+5V8-bL4I7U9S]<3S6K+&69OTN+bOHKg
EAW+#BQdH64A5CN:MV8:-46QL^M\>UU8?b,1N<(J=\CSXCRU[bJR#ZJYW?[KeQ&O
/GK=EU?+3BJ57+1U\4#I9Z#NZg#3b:N<&S>A+DQN(:1;I0\Pa;[0>2V[fI+#/&@O
&5A94U&Z<fC>TWe,^0E&VLFebg,8Y\DM(We--O&T,Y>;RP2:@b70Z4E#G9RNF]5)
:-,6DTeB-QgeWZ@3M=WWFg(,(\&MHZ8::<\1\(IQEI_XVF^5_BS7((LcW@>6C^2A
,)[\0]C?Z=_Q&/WPbR0UT)CV\;DMXU9-GW4=Y8ZPW_HLG-<Z+#I:XD1DCSBM)IP4
I(B0DcE9Ef<dT5.OS5F9ISBA4\[S=PX<<+3G,dFBBEYMGTL@TN8K<g9C&+=D00#_
-Af@[#NUKa;c;W(A-8]Ld,D1OJcUGVC9/.#A]E>S#(W7/,T5Hf2DD/Qb#&Y,(BUJ
&I]YN2d9?1,K4,95b@X@cJg,2W,Y79M3L22YN2RI_,,ND[GPF+D)K_).O\O<<LE_
,IT@L6E0eTU#H,Vb?=f8[8f=N/]>F<?U]f&KE=Na7B8]>b@O<H#LgPY,A=)_.-;K
efOHZ++eT#.f.F;^(Zd-\>VJDIGJYAaDD5=>>5X]93-MA@dC&^VNF._S^N5UBEK=
Wa]X=3L:04K#E,L32d5K&df1I(F@=7AGfIBH7EM&]541_&SO10-CaKcJRT^JK^S_
eIY18Y1.MH0_937Rd__;V#MUL_O\_e]F,b:5XSWa@6I&9URH)e<DLLJ,e?K8LdbQ
6T:ZdRZ,BIR;]HQPOWXc_KNL?4a=RF>@481AGEdM.e\9=dS?G3+L#3a30+cZ@Tb#
NReJN:aMB7KfILH(7(AH>=O9F+<.&c-a-_8OaeS:LaT;8S_@.XJWP]1B1-KC@cG7
N#>65/G:bS[OfbR^BB0f41)c=74(4B5OG72>NGHU.^G?M)g>+3g39LK=8T;>51HZ
_I.#6+7/g:DAYJYbE_,HBGU-8AV)KD)?c+\.+/DW;/2^Og@/b==M#EITTCQ&:@AR
]IJb/:,W@W?a;9,IW=eC&UIeId6eO<QC_gZ4[bE>f(9\PR^3A7bH_GENMCV7YR/8
+GILVeSD-:6@6>eE>b,TA9d1#VQHbRL5]N,Oc8U]EP+(]LJ\L=fUQF&=9/;)LM]/
.PA]AI[W=,VQG9fSDUdDTP?YQ=G_FI?Q@:XcbEM9[-.GAC0PHC:\PDP-EP@2DT;S
J]a-/NOL51^gQ66#5b5M,9eDFHYI/&b)b/TW/C5&VE/,Pa4IBM6J#_f-a(1-RLME
I[fGN5L#4-J3J2c::bCKA??#Cf<aQ8^&,4+VJ+e1)LG^MdJ=I5/SX5fQ@Fa+PM.#
,<IR[fBXN+_XD;bOM9[9McCC++\F)F6^E,.(<]TbbZ)M8Gb:Y\B6(=R(89C;M>Hg
G1,8McB<-#aaNb:-BNb<12;9BX4W69Jf=8#A4J&)(8fC_@R.96ad,?E+D2Y5^=Rf
;eaS8GGN5T.E_4LAF.a_&E(e.BN@0VY@=8[e[X@J+;e?JZE(;.OaXgg+/T1@ccFJ
N0^[UegSBO##N8OK#T[e\N(Y>?IDQO-#3T]2Q]R8gcQWHa:eZ_^+LOPdPN4830Ug
L5O;S00BFZbV1QXI.EB94HVg62OU\YefU,IM0U:,VBgT#\CF4bDJY3R\]OHST;M-
6S<_^(]Le9UgbbJ=,#dD&:A1F@;BS?>&9:-G(^6a<g&9c8E]AN)2MSC+PP-2/4.(
-bZJ7^;:Z,90d(K\XM\SNVM4+40SC8(fNB2)R>b617K2)L37S=;\::IPH:>DA<^I
U:P3&^&R\^,gKDP(ID6=O>@J]PL7(bLb/a7W9&d;B/[:()/?0_\S)JZ.W[]9;1J4
LLfdC6BD-9F\@QHK(9[B88TA)gXNT>(N534ga4:GVWGU\Q88.eOCF1f+JBDEe/Uf
2R(f/Rc5/d;2gKfAc6C/ffdHcO,T_f.@DR0#3;K9VN[&CJ\3?4P.B1(]Og0<3(,.
4<ffQ1HK#Q;bMLa4gOBRS@AR]>@F^+-9?PdG=HT6H+T#->L/DNIAN[5O.=g(1(]S
Be>MFYC_BR@U7]^DKW)&9c#d:QPH@KMNB4aJYROKZ.#IHH^+?2D<F2(?2C]LFgG?
&I]=S\GF4aY>f6OT4K<;\U-BWd:@;4)Q;H)#]f>V29CQPV3e9>9_eL26JNY@0^/U
\\+Y4W[U/801GQZXMQ8UC)YBZ/Y;FS/cK2_<<ZG)^W#4Tg_P(\<NQL:U\/N>]&Y[
.+A_1BdZc;D>01+cG=W&GPLZK3RI7JY4=[@NYS?(dN.bIe;LE3S(QZ;/.>ZE>]9:
WeeM-4QOX5B<_XaZ9-<[dM4<L4-f8U,TU&XY\;/HA\Q-T<MdaA)@<8Ve&=]0de&5
]:RT)-49Q@6^2/&5EIZ+ZFBW.7]]^27N_;0BU@]=7&fPWeWcO72L-^YgZA?&^A<7
\d(gSN:-1B5M2;>A3ae;N2U4T<,]4WAX2/?0d2[f<@XA[WOJG^OG^F05)#YFg,&]
,N57e<a7HaFHI8;J_URJVI\5Y2((70KZ8g)[>X.6B..1LP&bN;\[T8cFR4G]Z/f@
T,UP:1[MILOPCZ=[NIXf1_4TfA9g@2[EbW.6AT\QI1RbMKY.^6VUbCXddac7S1NU
,fW8F\a^UPDFa/8N9YUO\A0)LVcU3Db]DE38;TVT)8c/W2aSA<E7@F4OI-XGbH44
^I]D#&#aF15,NJ[N9;G.B&1UCV24f0PT]:1YZ1\<62TC;].fcF6@>7.=/?QPNKOL
#=S_@DO<W+e>>,0@#THS4MWedZ/S,@U1P&<F2Y3?)F;(W^4@)b3YM5367+DQ-,SZ
O)/3T-9G#;\4@N5Z_,@=Y#/<WHY7>)SQ;/I690cG=W)=.<LT;baL73?E)F:.C&4S
LfDX85gA4F+;)Qg;Z)(544#-6A+-S22I+APYLTgQ7f?)A?8)M@(#6Q/HPcFY+@IZ
.];KFPC3(bJ:Uc48-0C&KcV?0EV4F<gZ=-6G])KCP.eG/2(SfJ@YZ1eXUB^U82Wg
;KQf(Q/0))=DFVNH3c#U2Tfae66QCJZg^:?GO38+(DVI5;?J@_734P??.R2U/QNd
LG(=O<4?V)6&U6CY7aG#2Wg36EfOYTZ?bg#>=0JL-\NQ_5+W(AGD0-C,\VIHML0)
6>2EER\,f_Ta\^UM1]@gX7VM[IM@Kf-)04<C34c>&@0TNAFXQ\(/+;20BZS&&N(4
H,C=C@\\C,b(M/:I\Ve<NO)]/H@MUC_Z\)9\G=Hda@M+4ee[<Z;AcB(2>_+\Y\&g
Ee1,O4b1+W4DP:-N)-.]RIbGc]Q66=ER22PbPU?RU#QCA]8O=(,?-(a=C_G\cba5
&C+aE^<.;M#I;LfXc_R)BLe;D<Vc0d;EDe+[]F96HgfILf\1^X;GId_1-1;S:71;
a842:\,/D[\T^.4Lb_?Mcf4XcFd:.MXLb]ae=Y)QZLQ9g4FHH_CJKJb4cMDWC\^L
->0d;bHQWMeJ1F77MA^UN=^Q,G,R?8,Q8<U+>N>)YaND5TKJE97[2,eE>4_85U=[
>CPd3b>A&JI2;7VF+YF^-X98NTg@+?+(;\\._.g\fPXd9<[/FK>2J^(6XH^XWEQ,
^/=@;TQFCdJdTOGR-[_VbC<.<X_d_-S.#2H/UV=\]EHg)NP/@(&fI6B#>_aK+U[\
-T[TV2VS(IWU(GG\_9YHW3CdgQ[W##U9e6\^\]LGO2W?NG\B>\1FR=&A5Xe4N[69
H,>5.&/@>_I>L:H,)ZBPH(P<ccUDXAIUG04FOfA4T@Z]ES)_<&0&D98SI[;5U0?c
AWR#gG_?)DXHGHECW=VKW25GS:XU_:@Qg>@:HX[M)VH=E9e_T=La0c3U=_-Y&S:6
6_A3,@KSBKQ]f6L;cMT3[HH;eU1b^M)>)M>V26F\0:DE1[QV<9F,5]?IW2AQS^1E
aaRf,M=#;.8GaHB]bW](6J=R-P>BdPMKI22O<LUd=WSf,@aO?8c8:6X>FOQH(UN=
+U84bOb8Ad?9=LfW@#9:^=@-BD8K37#16IITQ@UaGCPEZ3F_.I5c,Hd+.EJ4RK>I
)f4J@7Y<(<MO.CRV&90V7WZ<9LeU^2V\T34<=M/UFL@P0(c8Y)GC4b./<SR7:\cW
2((.28e3U@MPN?CTT2@KLKE33^2Xd&3UAf]=BPU0QUX+)KJFHCH/R_4\]]Hg0Z?T
YXN+8?EBMRC7bR=.>A1KR[YC;_]Mf4bK,3+^d,S7MOZH)FRNMB3F5f5aGLYL:bE)
6#>[J#bH7(^G0M1b)V6(Sg0g(_L+B8CI4+&)EQd<\A+#?W)OUNPR6QW>SVE>.BH?
21VHRC8+dB/ILLL@W=]A7G(Eaa0;_P.&9;N.cc#B(I:M,XJ([Jf;/e[)<D0/ML)S
?Jb8Eg87H>gYCfVU@M)9WPO^:+f,9B6^S,-fd]Qc(6N3(.cHSBGGgISHG7F>5SdH
E(?]?F4g9Fb3L?[.f_OIFAaQLY3?RYM.3Fc>:H5I:4O2,a>D;]gC#0<2=M:XRF_>
]=;5:4:de4^AB.>&]1]3G]HQG[SfbK:SNTY]IEH\4;.F0b@Wd5H@e;RC/IN;D[<0
W;[S=]QW;U1eXU><1c8MH8@1](Y17a]#P)-\:F]0&J6&5&,DE];8T5GaU?S<5&>H
dcDOZ+HPS2^LRH2;FL_S5N1N=JaU:]<UM<QFI&V)F;XE,XG>O@;X;T\:499TP:9#
fBEOU2=SG#S>KS#Yb0V4I>ROT>OY,5/5HEO#FUcWTBGY@+42-dJ\Fc4c(b_-7Ie;
SS/6/UJ9UMdPS@11O(2P#58VO=1LI\_-@&=\Q(R\2]/L^)LebNP;&8>2Y+:(YgAR
8@B<UUP+b;YLTPCU);]9ZX0dd??AM8ZB>#O2<S6d/NGI<,-b17B+?fJB&R28DPU\
P&[K7dLce@I,G3ZD_3@M)F&>aE<UHeJ<Y<+T@Z1fOFcbfRODNVBN^[4(?,&W)-#D
+L+QX#GD=]0^DRUND+^5d>P/<05:61#aI[c/fc3E&L[E=XVR6F6EAT_=M;M<32B+
=<519Z@BbKI#WGb;0?YVJ3_EgCI(;f]^_;LEO0H.&=(8^JY+3cJS#QO\3/g8a_NR
98Eg;.=V>YZ9+6\NN?,B_0\Z=06:Y]VU:IOQQX@K9SbG2T#?TFC-.9aF?<E&[L\U
I+?;KfgEbO8CG[5V1\:2T,D<MF-]K=J3ACaRC7+]WEfQfDNcL(\K,>/[RV]A]+](
1dK3S-4EAP@[;E<GHU/1\-_TdQ/K^aV[CX>V5Db)]QF^PcJ0(HT(@d1af<OK5U4d
N/3?6]F_@5,@HI?<;&X8(?Ab[OFADHeA2V?^e\-LHeDSDD9gJ(^SK&X6?@LTMAHF
fKg>T&XYca4=BBZB^Re=gZQ4_af\/3RW43]dc6fI<-ZYU:&)>6_,X@Y,0SEW9D]?
gb\.AF7ZZPB;14UI<6[?O1=#\Vf]gTM6A/RJZKVf2<4^g0/D0N4EMYX,N_[-05D_
bfJCb+1L7Q<H(cDK\GK(L&WFg1MJKMG@L),)8[1QIB,EZ?A[H[D-]-aX1E.&NWF5
6K(6<QgCdJ?R<?+F_72_2SeRZcMO-F04e/]]&DA7XZAA6.5Y@>F@d[g;d:dcW:.U
8QdI[3c/06KNI5^S#XTC#[-?d3D44?GVN;)1UXNGZ,RgWUCF7Oa>-B+/1K^@Yd,2
900BAHGf?-]H=DI?R=^M??5>(LMI[=0)OgQ;&JNKPAYJ<?Y,bNb,TY<U/[adSJ>M
Uc3=ODYCG7,38P.XJO&BAVe?e)^Tc-8&dR_:?If8@f=J_)WSe&>69;0LUbURA?0F
g>FVPC4++6_:1eKPZAG[)b#,AR&(V@Z3XC=8N8P8R3dQ/4T7Y^788#]:_8.7T@D]
2FVZ#Kf&a4J]?:EZDbWSC7cXgWU9PDf0X;0;J-O5OZFWXVL>U_1([)J^04K:cfR9
\)Z\1^<(aTNP2a3&6X2UbMY@Qc]0>aSW@XGQ3H\+Wc+<D>UY4aDP/FPOY[QN@JH:
EII4]9-;C+)TU+@6):KN/Y\2Z-(F^,ZV#gT>(K80bbZ;F,QVZQYDZ6QG42M<-]VC
J2/M^,I#A)(PH+GPcP]g1DJZV=\3,Y&B7X.e+)aOg-2/YA#c<@L([?V)>JG<L=E1
#ENVC&6#Ee]A3)4GSGUCZ1QgXYUcd27B8..aDBQR-G<<.AO,MQ3>0^3?-[W,CO\f
&HR:P?(5b2,I>=-eMg5gDGGBBROfV3BcSY,5a]>9<YA=O/f_,T[CVc.26\M>=3\8
R4]248O@8]OEOI,70IVT6JK,1,]_KFQG)L1S0#(./7[de-/(O>#NR=>>8QAcX)SS
9E_;>O1f[-1#6A24C9VMaT))-()0;\T&:80+d+3b&?Ng7?1R^4SGWU+_@Z54KO8K
eH@>1WISfLOW@?F;6+\BPc>406E#G5_6XSbGQH;RE8(OU)N^3<H5P@4YGd4(AO\>
O+TLQ\;54+)#>X(:H?CMYG3Y_XY0,2P/H0IAVce97LJa^CF2I_PWYNL+Z:79^gN:
+S2HDRX45S)aF-U1==E9?\_=+V7,e\.gc=4A\G\1(L?[Gcc^:@#?)R&08^95:28I
FYSYFc3.P:c7RKH&d#EeX>4,.0R_Q&/^]LPVa]XQ]e[I&/ZT+(7GGX>I#>;GJ:#)
E/^aJ4g6U(#Aa;7<fAb?@9,GRO#5@<0BYB=(3[ZQAa#cP(\P;<,Qe=cCXZdH(ba/
C^a7VVYSN6WX@S:CSO.)@/dZZeY?d3^a=5PMQA;\I1ccbaeGDc=_^/c[ST(6H19>
@Y^O9;PG<KE88da)d6Ca6HNV@FE3aQ@C.GQE5XK\7Y=51#IZ9+;(d185#d9,afHa
?a0W1]15K&(&Vc^LPe[a8c-cF50L)3C09Tg#g76JITQ-;ef^/34dD7W_ZdIEd0@d
KGEg>J&&?VY.cJ2:3@+3REe.(Mc7HIJ63b=d\KbKQF1>edbZ[(W116N(=3YZg2-\
g6@)=\E79a]0_ND0Ab_27d.OE3R&NE/1IeWeU:4=DC/>H9cZD<L514S948-/^ZUB
UcRcJ^GR4\Rg9CGJ+^O/#]E68Z6/d:?^R;6&1J+^CPM4,4+@5H]ddUEY8G:1N6+_
(^aCA-F_2E<7\gS0WY36/gVW-HW4;<P(D#FKNd4HgY]<c4,VI1e]gB=.OKLI3_6&
AT[[cPf0UGe6M_EfX;GIFb^HNKf20F\EK\b^)R]ZBF_LFd3M(V4&Q3TX1\K@>TMC
aKU5]<NKR99IQ3=L/J;Ka\#&^4Q>F^1SeV75R1\YA[(>A.X[6.:O\=CE-H6\&6B3
,G@KSDZU(OE(DNgLY7\Z2d+7T3Nc7MHOd]J(LVNVGT08)0+8d[_]ZZCFB5#X2H@c
/LXe0/E,J+Ef<_E1KYKM..C>B5V3_GD?YAFcZP_5bCcLcK;3?He_fM;5c>UK29d8
=JYHTYNRATa&4EI>L).B.Z>F<\.2O3bHKfZUJ:6e+MA/4cSVM](e=4b2,cccZ20E
fHCd44FKD[bJ^R4)J8<f3(:GaNeL_fV3=X?&ga2d#-a6NZbHUR(TZTK7fd8DT]Y(
F,Q9a;LE#fIed(&#=;PZ=;A6GN?]8]_X3),).QINg_R0OL(/:bQ<OeDX:QdS=b<Y
T)^11=d(V)[5T^^N9Adf]^U#-N7#ULV-^&VcH)I@3.ef=RS]/28=FNCTg/]C^f2S
+W17eT@&_Rc5Ob\0]a4\16g7;+>c^(#YLS>[GG6ECSFI^R:,EY#6>M1-XRZY#?;W
,S\bXFcMH8&,B2^/<=#SZ8CRW(W8@Z,aZKO&Wa;<c]gF-6=WE>^^d(bbY&3a_MIJ
8+_W.WZ)TbOKY_GcNDJ4[KIZYAeJZ>U7X3c.QR>Q;9DVE3\]f3V-e3b/_9/(:JB\
a2QgOe1)6\2eI^(3D9O+EIb54U1d_.f_&V\1],D3cD<\GSM<7fJP6S418edgG<#<
Bc56Sd35PWKQBP>a0Q:0X]RX46/;0UX7?UFgJR#c@KK1(]9[G<CGBN((RCMCJG;a
+4.8ZJQ/>ORfDQ\Xe=N^RM?b\@BR),>g2?U/>fZg^d&NE-OJW&HVL?9K0YE)#H</
ScN4UKCcT_V1>SBf8S=,,a:Te]A\Y7.^d.GN+05X57J0_[,AHLGd5G.KC&_SI1fb
aF<_E#GBTB11;e][9>(e-b&@Q=c0^GY;1c=>]@b.WWG(GScg&]:C^]\@5</<QQBN
Oc9O\B7:S2LB:+A4d/74d[?f^93P//#20Y\1O9^L7D9e[5G2M9^RadfBJ@/8OVV.
>768FXE()d(]5AEe[HaR66ER;&FdB(+T7g)[E^^[ELHDA#2g0&7IIT((A.5aaJQQ
8:<RBT,@-A?S@f\@=,5(KSD0aYSPW2ZaQL:fTN:/[c^E#ePS.=ZM0]5660T&1&c^
BH5;E6L]2WYdceI^7T<fd:b+M68KD>Zb0:71W&Q3HWN20N_1e#E:ONJG>4ZPE_[Y
,AH,FIALM:.+A5&3<SS>8SF35gQ]C>LO_=/-M&H9IJ9fP6=G0R4;,<G.T8GUeU-Z
=(T\W)6\M8./J=0)&FBE/U47Y6VY^\A_:4;6P>E_[cXgH/QC;/BE2d3b#KNTQBQC
91Vdb1GH0NF4,?@,,L6U>Y,9B97Z=f&K,87ZHR;C[[=C8MB:gdSV9\YAEWIP>X<D
](35E=KJRM#5ED&\@3PM0,Q2+(4&;Z,I_^O&Z#;Y6FHGfTCR8/dXdK.#G>c><LGX
_9g,20c#>^[(/R:0afN[,KG2d/CVV>AA2+cd^<:J@EQF8F)EEO[I(UR]X3ce[OMU
/dQ@U/GMJ]XSd.C]8\caS4>7Z??]b>:M;(UT(eUS6VS+VaZN^ET9fVIN4=)0#;f5
UW3.]\1.JAI,[/4eT,U=?&W_7L35L#0SMI0^CSI4WIL#;cS&30[@-1#/4(M]1g)E
\NM5GMZ],G+9#/5D+6)G[W;HXX(@LcNQ,\OMJ/RR5OJ.5_6L3]##\UYKcV=Zf[48
,aTg[K1S2\5C_X9PTdNY+7Z5_]E4&UT<-ZAA_Ob3:,C8eF1bEFARU)]5O>+M^YQb
4C4f,ab?QH@N(+8A7.?M3MEg37;C2]]G[)<R)a,@RG55(YGD[g6L^]_CWQ9ee8aR
^C32(J<XJ\fQ,BdWbQ#G,-X48g[LCV7E3A[?;K4&=.TQKGRX?,G16c0/)SSEe7G\
3dfQ;4YA30I2IEX,NFL8M3bO<\#WINC?K0D/Q+LQ^S5UbP+]#(]&LN#/3LKYaG0X
Zd;_3=3g3A;deffJIJR2c8+^Ic8+^HT3-b[G<@Ie1B.7O>&P9@Kg+#WfP/..6/#@
3Mc/bA#IfI,UX^39KS7HS1T7(HZVaZYe#8EB3J>0>V=/S<LO1+Uf&g50>.IK^FaK
4NCM>7<KHdR/5=B,Mb+G_F-eMd51T\\PF1YbJOAXDF</WQPQdU6AG370.VIF99Da
^7fcZN0^N58T+7NVPP08g<b>=F5_I40@P_2fVYTOJAC@^TS0<f7_<&WL_PEA[^[T
6XZ6WdfQC(ZYY\EKe=SFP:dfG@VFcZOeE68\,6F>=f+O/eVB&aWK=&S1B>J11f<O
B>K4^]eSQfTP0B^L#3MS+2>\c-9/-@E,fN2.^_R[dd,70&UX64gH9)HB(372e[]e
bGHdX3bEcCV.2?aY-,)^K8.O=S5b20MR7K_9_.f7<]acbI=#7L>L7+20.RX&e1,\
[Dfg\[(#D(-fGU4NQKPR-e9V,@,fB;(L[eOKgO[A]+9-D)</P,GaF9;FQB_YS-F[
5;&B&BLXHcQFeB[.MO-..KQ@?03-MW#7.XWKR\]1C\Of_9]J/ePLEd+eGeWWLVN/
JgYA3N[d8<UK(>[9OLNFWQBaVA.)AM90B1#[MEF0@;(.XMU=b;1f9HUa-O1IZ_g,
8Lgc6F0eFP,:B;KF\XAb<G,-MDYe4_1-fMfZ?CIQ=XRe?addbaME>Qa)6,#44E+/
O?T<H^S&_OaI&<12P\7XPcN>(_+@#:QE42_9HU.#O,.bE;[MMYNEN[,,#1Wd[9=V
Kg8QLQ;c)-._<C)CMP6RaELe6fV1?CG,R&;])g\dC-+.-SDB8;B\EHNe4[?YbWV_
3N6-3_L,/+A1P]\)MDVRYW)aL?ZI5Vf,QYW@J[5NPf&/R_F-aEY?3Fa_+9J9F2gW
U42[6D#>=G?#LZA(Ud\9cZ[;6N>1\8KU/IOd@;L<02ECN2\(Y6\>U\V>[JDP7,[K
bHR]@5TU&^KFLHNVf91><,caU40c)?T=>D9f>27P9>L@G91X6SGQ\e7B8ETdaJ+1
ENVQ)gLIE.a6<Z1P[5T.OLdg>5NGa,V=ENCSfY#We6N]AU&9.2RKYG?d6\/[JfO]
6(0XL6?f0_NBE88.[3T@#Q5,O.]S013=aU_<E):adL6dO?Aea0XX&/2f#LB8Bf>@
2UB0EKDDXSJ]L93AELZN#\WS;gN;(.K/M</Tf?/d()2V,Z#.._#:Q3J1/D8K(G[L
G_.FE]1M/O2[HK[VI5PSd8?P?I7[OgFJL3>FKA0aG2MK&aS54KVE1Sbga1^<4)#g
&J[O1LA)YNcI;ACCE4^RCZ9Zae_YB3[TYCZTdWO)0ML5=dJ/A<5HNU/#??<H^N,g
,)1CG&8P,SWA^]X9TR1&5UNGSbGg>&dKS4H^9DF#\V<6V(5-Lef2M=VQ=f3A02WS
GUEIX6dFa?(C/e+cU;U_=&W7(ff5gA5T3MWI>V+]9#K[RSC^HCR4R@I85-^cK8Mf
,CeC5)H87Q@D=G=:QFL)A3Ff0fN[Mg4CfC<c.BaLQC=MaMW8PaU_,4\=Hded,,eE
JE=c;[)D9&.gc726K@Q=,&P15VeKTQ/d/\a+YB6\F7CE1eEKCS^,aMT=A9FQaDfI
a-&ZCCA-P;]#J&X=7D]B05B0Md:P:P@LVBYK3E28eFGUTaLI5]f4(+Q_MV98K.]N
R\,9QMWL=>CO0#)a]Y9aE@0dO_P=/:K>J;#_&:1VAC?a&5,+^#2:MA.LBTYA^)=Y
?+6JD7cX96cG+7^N9DHXVSFV.C+AWMUN_3==WKbQZR0KI1^e=I2K4/LBffUM[AIG
VBea,S<_@=eN9KO52N77:A1(><LQY2WP.[HR^dJWG^X>65?Pc4?2.f/FZ6c=8U,Z
5=[5>H#EY973UL&dP[E#0CE7>K/E@QIR3DIY^I-J^a@bKS^OAfcgWW\0.=^:#gdP
ffLAf\eY>SO-<)J+Q.UF7Qe2RA?92_QgfTf2,\d^e3):[D(TR+7_^06e,3Fb^>>T
RL-C8SI,XZD:XA,Ud-F&cQ2?#G\P:EJWPMP&fJ@BIJDCU#K)TWPY8\/Rd4)=5BC2
[+=>F4[SdC1VV_SV>e[.W8??RB45RH/=DT0B0/UP.:[KM7d,O]YGIGGLe>-^\CA_
@Xf&8d41&B1I#&.Z_1>4-EMTE@I<2aQI].8:R[aSMZ4R6<>B3&9W:T-c9U;UX/()
E1@QBEC;cG0J95/.WVD++Xb_K3A;g/4a293/L4Y,(4I@SNZ6=F4FDE>X=MC1#69+
S7K;+_4H;3(4,64@+8.;TA,AW]Y-]7RMID@gE)B\dCNM,QBcPQ#b5ERKA--GReSX
RO^0EVZLBe_bfaZA;]6M>EQAIIRZ<(.Q]4S>ERTD\Z)JSGG-eL>&5ee:Y3S(eaX>
W()9/TK5fTWBJb^0):##RaBA,\]LDN6K3767KJB^ZUI-;dDE071?>3T8]EWSEU6D
=.Yf5UO(;^^1RL[[,Va(6f_E&(E3)cR<WB5]P;eNdOJW_#/649A5PaL47A?NEMWf
01B[SgSTO3L,:Z]^:?&4B?HOJf=6Y1CY6Qag_Xg&XaP].:2W=Sd],&519[(3N_0W
c0^Z#Oa&<:N.f-3gHZ(SKI0CPC[0f)b@(:SZ]80Jb1O>#5(3ZFTX:NbUgLeSZGH\
9PQDLD8DOBV^/TB=3U>>OKOe^VOa80JPJe?=fX,W-+AZ+1BA=B,fD)fAGc+M_U:_
7CF]S;5>M]G;.GU-CN6HaQbC/ATe2(GW2[7S#(F0?,<4<d8MCTb:0YX3H89UQa9[
M(]SSVSFQ\N:decc_V,/I[2aMLM[4M\T)LBE:+1DS39a8)Q\cJ-@aWU&W.LTU86M
_cS]g8WF[bS?PBI)cLF#LG1)caR86(TEYQB^Ra)>_M-(L&UZ2Z\37DV=-_Cc2Bac
dgMF<6;KSf6TV&V_dP;2FJRD]+4Q3#456.CKP,O_]+TP>IYG:Re);UMKfBa12X\P
9dIN^b=:dT(LB\MbZV27TF))/eg0]M>JX1\(W8Q[&^RU7D73.=)S(F1YL32/?4Ug
Q:)Jc@NZ[9IGF::>eZ=53DWZNN2Y>(((d,eg0SI[TCX0c3EJQ[:F0RARJW8B/.?O
<;>O0EPSV>CL;N4I9Ie15[?[;3XY64QPV4B=4P/W<013^IDND9:@P@T440+SKI)]
P@;<K6@Sd8.6#1<g3B[52&8<R?a0OAaB0Be4=-UY;CJ8_;D4_CDg]R9g<J9ECQHK
#BORATgD44L&FC0&>Z&IH7;UOa?HbCgD0&.K,e7<<IWAV,7D??B]DYWISOEab=a;
@)_9]FeIE-?[F&GgTc\fLXIcF4g/cO^ROYBZX&6L]X8=XB9c(J6\0Hd;U\:S0)KA
BK2;CQN0f]CTgI<[eC.Mg>6]ONZ_-.)Y^4I,.+A[gc9<9EM/IeFF2GH=GTKSHPTN
3QR0)7MK)-6FAJTM)EB+,U&L]QY7_N\e2YARdc-L-96)R:()B?##RWP@O0O/3I]N
AI^GD]Od[7@T_-_^V=),?N1G>3)0ICV59+T#5A:=@2R&Tf3>T5U^gN4<-@9OD?e9
YgCESD&e6e>+,IQ5<GE:\^-U(>a:SJ)GSBQaWP-7>R3W@=d8M74&]Yf9Y&aFAXTO
g6H_AfFN7,Z7-<.+?7?&97IV@B8=]4J4g?U+;B1A)NN,->dUAOZ+&dg;Q\PC[^C4
CdH_eK+L[\T],\:=,=0_:,5cf3.W6KTU\.<X.\=#:1/a9PSVJ7Z,3,caO/[3?:A)
TG;X(cf+:QQR+H2)Y+(F4S4RSI&1ce.a;?NbYgVTT;@Q.\fIKF9eD^P#d2YES>Y[
6G6@Ue+F=SS@J/J(I:d\,95.(PS)?#N#;ab[V8ReCgDd16VR3e=KGE<#bV9-K;M9
Gg#32;9(F_LS\ZfFA[MYN_G/YBT=),KWIgV>[F<0ZO+9+CEN-M4PdQGOP5b]e(&.
W-b0\&=@TL;94^356R1#Z39&QP99V;:G@I[W+^LBH]PbZeg34=YAI>F?Ub1F+^f-
2(7YgFHa_19bH+7dM.ZH+82&37RBeL]]#WR=gQgCHfH=4;W\/CR?>#)e/3[?&dAU
7Ec@Wd^fR?2\e/#937^g2><)ZRFJMe5Z(UYcK/_(&HbKG?.,1FIJO5Q?DfegOG?e
@RG@U.PGa)M96fRgfe8b_?PBa64ga[,G167T#R.-#MB3YE2UX44GgeU)<N7M85I?
PIP?25gM6>4=1\:=8Ucd2-?T__JbJ?2ed8^H6BEX7fU<EbaJ8&=&CIQ7g<f\PXdU
8Q&+a>aEMdGEKON.=E+T&BXcbPRdXM]^@K?C3CAKL;?N+Bf?KUOXU/9VY0O,X9Y)
^P\5<T3]5M50[g)S<18dO:L.#P-LffIAP<\([YgbSV.:N98QH7:\83#Hb;ad71&,
QBN3@6<E/DCB^(g^[O(a(U.37D[]<O;E7Df0<<LFQ&/5.8?XE6A>I//=CP47BA#F
PMG,?Hd5S)[BY+&bfcB>(..#&YdJ>EEAH6/VZW-S=K^ZU49gPM8XPV9f(3cB9?S<
g#+235K^O09=cI6HFDeX:1>]P]ZKd][,B8O@A^O6]QfAJO?4JXDIbE:7^COCcS9a
16f@2U)2ABWKRgY<?_Z(.T1/Me.]]I#WcWBL)Y3PS3>SI6,=H;IaGEW_(/Y0B[H[
6D(?4]CCXe=2B6+cVGUPB5[E75e(2eS4bH4C3WDGAWFFQ:EI7ZTgIR>&cR232Q7@
=?:(9]SEfe4XRCS>&9T(TFKJ,;@?.2NC-3EYCgJSVNOCXEQA0B8QRM=bF#TK7\.\
?&16GV>ZQE)]Ea=J\dd+:[I-[f[\4X,-dQP<@-37>-C07K)SAO5a/Q,CfA=H7,bf
e;RcN?+1D6PMSPPS;6Fa@]S<NJ3@,1,04d0BP(7QgGU;9-eH1D8cISaH-aPIa>5(
/\2M;_E?dOK:.gGRRO<J&J3&1)Dcb(OPW=+[OaVCET9H&VN;,aGbTMZBc1L-X-U0
U0MM][EG3d.I4D(0gaI@W@XTX@bR)+?+a[H@Adg\aV(/[)V/&OPL]/\33IcEF[=@
/bGEeX]4cAd<&gPAT;U:dcX<IVAa)eCaTOJJ-@T63M5+6N5XJ)g:N:B+c;:9XJ78
@TUN6K9#ZLSO5TTb?>GRY-1cg@Eb)YMe(J+K#Ud?@3:SHZbSCGC1#-aYL,=:YADg
APM?0U@fHR:+>IT.VH77<6PVUegQ<7VK8NRCW0GD202HD<R>fa=?-g&BdBU)e3HX
TdCW&9EZ:eUV]8L]:8Qa>YRF9XD?I:]BX)QaAPdZ#FK-J[R-f0e6FaH5UcN4-TBN
XK#=CW@cLP6XEE(8LQfX]N=c9KS.R]&Y@X:A>Z68:@:?5-]08FOf(53bICD/JV?^
>,9QU97C.fbbD=-@GM+V=_6&9)ZDIP484CN:EXHbJ]:\e-^&JPG@<_fVUV1L>ALA
<>ZeO\G,:3PA03^F63R1_e7L[MW@e>4fJNZWUI)9@#Z:2dAZG4ZHaC(dDBWcTf^Q
8T3,C)S)V#&S]^M?/@0Ze6^6&4+QZeT(38314:DET2IH026UU=aG7CR7E2g,NNWK
XQ;NKca;MLHPOX:Af\C1=9I]/6,EH.bX6+Xd6.Q.d8?70+^\L(<K89)8R_X(3DCM
/#.0&BYDH,#dcc+(g3fc:Ma3FS.gd79_:Be1D51U4<WTMOg>dW\<_YM9&?Ucb7I1
IGZ?J52Y/,V.Xc7C9^]GA\-IA0]O1#a88E)AV1^HY5EeUZCXMd8-XESeZcT-4S9V
8I8Ze:2H4Q>=E(.3e?3d:SVfJ:f^B0?AH+M(&Oe^caKO17>;[?.IE3J/@A77[S+E
HZOZGGLfaW)dg5(+O(TB=K<a--#P/U\+(V#Jb6P1X^,?dSE&\:<#,6X)_S3VfKIa
d&59eD=B=GV+eXZ+D+;FRP;c:d6H;@UB#(S7#2_,ffIaQ@JO/,20JcPA>?OC/.a-
aeM\YIb,BQ,>K2YL)c.dWAS:ZD^GQ3M+\AK#8aV1FIbOV?:6?@AE\=/+3c&\@<OI
&f4Q[O6YMHH:4=<6Z;Be=/862_I/F4aSI;9?[ZfS58908dFagL&TT+2^5B+KgH&3
^\(7W7[.7.(bgNAVdX/A@\Y7-C2\#T?U5)gdg>[f[4Q6.<4O.AVX8P;L2E[FR+Y<
E,D^^A]W/>b/eCJ8ROfN+XVAD83R53&&(&Y/54PB/_:Y[,&cU831.Pd9RH^QU_gZ
XB;=CS)E8gaSTV[g]WVW>CUa?K,OEK7/4.O_9]&P1\L(5S?.N4]>TdM>W.N5:1_2
(6A(&+BU/?].AJC=)6R<ScV:]=>P;_V_F@X:D@F^9g]UDE;Q,#C?V#6046)S./dZ
#PTLY2)6QK8d:NSUUDDbfg>0,3&g\<A6[.C/?-NN;/EP71JN#G&HHP3,SF_NeV6b
I<UTG?HN-?]EWFaV_?B<WE+T:5b?f+=F@=<a?:\4a9d81Rbb[f8JVbN(0WgJL<YH
C>D//Q:,;OI8A0AW;^d939Mg.F28.&gX2cGIPOUQR><bH=EHICQ?/J5Id(JNEe4a
&J.:#867]d9?TI;P)I#L]cD5\dGVbF+6c19+OgXEf<Ic3CH=L-]9)=e.T8@@,bfN
g^eZ7TG^,5O0fY_N6I0Y=g7P_Ig69P1Y<ZM8)YA()0QAM+g(TUWa:\BX31)=HS1V
bg_G=T-be&ZP>W9NgIRbBIXaTRaTVcB<<7dO#7:QE/c^@&@,G5^:M8GN96C.I#H:
N,8_g41-=B/K,aBBSf,A+:gJ\U0AJ-U&FMbWa_ME7E9Kb0Y5:d-]E0g1</>?G-Lc
N;&E4:b\0LM[Fec(<-;7]cMZH9GI##_D95Pc?86A@W:-7K?;\3@@<YV^V96U[e3f
XHE4:7T(<T7G0V/bS)I\DEE&;,?]UC=)dKO&a/AXfH_.](5H8CMO(8bgXdO-<f@Y
VN_^?Xaf9>J&P[Jd07ON\APY#f(e22-^&?YKWW3VbeZ&9EQY6:e96#SMH&BU7?K]
2#0CZ)b4c#4[3<]_E-15&:Q^f@=THXTa97DQY-M[O2+bKDQ1Sf5g?FXF?Bb5MG&0
/@c)dPVK8dCDTZR/60D6+Q@D7/ORP)XPf7I=A6NP?-<bD^:+V595[B_;?D6L+-VC
JM(ga]O;UX27+eA/8M0JWV@APb>C)Y8Zb+Ae1(b)bb7H((9=P8^(XZ6P35CC=#<Z
/(;0ASGE&fae=M/<>8NPBSJLYPOcCI7f:&VULQ;Y:Qfb1;8@?RJ8(3,G75e37Y&4
Ca,+\b_-B@#g??04@&=0S_Q<X<&GR5T=>E#:Yc)M5B>@0ea-2TV,]GSe]5B3;0R-
>gFe96W0#J/18@.[PfJ-V<IUQ;+]+O,W@3F?QIRYOd24GDQO0fWKeSNZcdVM#NNV
SPI:M?QB2DTHdC(E1I_?_P2(=(5[?Z2&3>.S5URV3+T#PN-A1_B3a(+<f=<;=KN<
9,?)^M(Qa#J->7V9=.@ALU9L3P.a^34cW(Kb&&eRa:6#8QQ\\#-5SHHe8?6Oe[EH
c5JM[R<=#9S8d).4U2P,6,D-BL&ecK>,+Q_3<eb&36I;C#+)\;<?:BbHOP[V\XCN
SE_QXe&+:H=aDS#.fM-0gF0#5[Gf;Rece-+^5./QQA?_,2.BGTfcRcfb(+Mf7XU2
QN0TaZI?bW?9^\Bb4=T?3.R?[=1RF#V6(_>:&I^<AM:IIMX6KY9CQb<?]0L-/UcX
-WgCcEO\Fd[(_^+0eQE(1We-G;6/;4TD7;_^DdM.F;YbNSGK80,@LXM^52eSbNYf
,]LKcE>_@C^-I0,(6+7I\2+QSafH>(Y>XMBg2;MNf\QbJ]W6MMJf7d3GKce=5_S2
\L;(M(Q:US@?B[]4M-EaYS/R)PO)5>:XcG,QO]a\-302TeBR(_I(4.?2aC]ZAfef
+S\)(>N:52+NZL<X0>3e&+/(N2)J_c_V^:_9fW#,/=#K?;c<=,^L\HA[g8O[?GIX
0e8JA)]DAf+c;f;/?[Q9C9:2S7EYW2(ZN\dVD,BEO\O<)=Yb]21+WDX:..BS.4AG
#4</C3KON46cI4B)1J.eX6F7R>Z;9#_O6e&EXSI7DI2<dc#-J@>L?LCY;Z09AY(D
+C>fFfeB)fZ7CH^4U[1IR^AIQ3M\+3N1XRY&C&^.XbH3dD/J#,J()3>;&>53I8.I
V6c-J=_\F6M55c1dF@Z:Y4L&[AU?c[?f-&G0NNOEgR<9G6/EW4/^=gO\W,=eO5B0
,BTL#T&/TLH9M(L_2^;VEC6W)=F(T:4;P@&aU:]ILK3^KG\[AIaE2OFHU9@<L#5,
XJSQKKL<>:&UZ4^@<7E+&PMZ5<&5&D-NEEW&-O0W<>^G(_&e2.>JY@@\V-)b,d_/
@:)856EVA+3\g#1ZD0SC@&e#38QVb?dYRS^IcJ,Q\\@RV22ML[_QB+YWY=]>Y<6K
BRF6Y?W:A(CHea)d\_6MQDW@=GE1SR>,.;)36@7\d]O)R=[PQf3BR9)4WI:.H0?R
BcLPC@JR^3LC93B8@c\f9-^C]2;ERf]LV8Se;D@>/2UcST2d&0cIH:8F,g.4;SF>
<STgH9\XaG]VZfU7[69/_FUbRL,>4e7^E.0+g\8M,K5K(f,HbP)M#6AXWb5ZL3>+
UIBc?S(LI^G5dcX3+e-E7KHH6.+D)KEJfHX4@UaW//8C_RJ/gOYS:.8fgXf\?D-<
CW)8gD6PfKH7YPOE#<_0@?K(=N&Q858EB2.=f#<9;=R=gR[Af+<6WLOD87IS9=9^
Q5@8Xcfb7]>IH1=H2G>MH>X8Bfb9\R>b@f+14^CKV595JH.&S\HJ)E&bMQ9A=VKH
ALKgg5F;b4Bg8c-L\9MN@f23FGBEOQDK76WfH7:FH?KgQOI_HCB52D[4Y+LA/F:.
cO&(L4R0[I_QT(W#P15Bg^VJL,L85[8I=4KFCPcM2/J[6+7X=M3UZ;S#8Md1.9+T
W)THW#O_WBIYeA/U5f1:;;/[WXUMF\Z;A77[HMHOUP+RJe,c=c4_G_??).=?+:-A
D7^AdIS7T6,a/:U--+B/.[[Fef(IDdHY.0;8[><M&X6[g@PF6N^.E-A-M8ECJ:9.
78VO]6B;93.XRO2cZ/I(_OUJg&GU.<Y/2Q;WC(T4V\c?OdH[?:=.JU&;HgYgB8Og
fM6B^E.)D/RM?(C<ML^bef82XcK.gSDN0@NIR&GG#7PNEf@/<^P+Ka3_dUWfVAX+
WR8^S/PODDC-C^#O9(#5]5dUQ;T>a>>IW@,8<S_5A.A;SeF+g1N.[C<=NYNcT0XG
Zf0bGDXY\0c21E,,C33,0fO,O+:UaJO?=NK];6:A3b99TXH4]Cg=[:4?7DV&O.fX
Y\[,UU_O&6Ye[1fUM__;<.R\gDX\CKM?RUV)@S49L/NC+@fL-7,]7]\ZGH9\Ff-F
H+c&YH\#eUX-4,?D-M_41MT,-TLSGL=O7Z9,76b80b_?_IU4HR1KAfE.BH\P#M5T
&cP3OG:ZFT&gYfDMV_:/AHGg/a9J+9\+1M&\R^BH</\RUQKT(V>3FHgL4f6#f1)&
[PHMd]_#-Ya>AfKHb=Ec6Pd66A>LDcYb1P2HVeN/-?R_RJ;.#^_12_4GXKSeE8]_
XP)(_6=U-SFdM1b([W@(DeDb9+;:HA>I;1Ud9?/_1:cF\@_FA<Rd#gV<d+7<O(EA
Z-1[X:+&Baf(1NeH/FNb:J;GQ+YHY@a7Z+F2M(6SVR.cR>=YO=)T+0QZ^b#TC-LH
F5LQ:<,ce8N3^MfLg^BQZUg.&>g:dNZZZ62U+=:bbR(XEO5bF-=+\Y0OE4,XJ[5_
3;6)J67=>?P9=&.??>fS-)DGQd0=X-7876bfV;+-+_gc0>XM#?]7&ULMX2G(R.IC
6+76a/PF(#4WE=33X9H(ZGZCIe==&MZ?[^>8KWdWE0BA&H78+1?1a9?RD[(+:_F;
df^IZ95E;19D@9>3JeE;ee]cQ/QBbC6A&RS5?M:6?THD0B\.I;.)K^Gb+2NIO+3b
+X1-M10GOJ1U?V<TL=,:EO_0MffV96S:5(-)2\8&U2\,:PEQPY_9@O6HdA@[,LcM
Yf4.GP#3/ZMEE&[5g2WE978C&b;UEdWXK?6ZQ.1RD0:a_F8Lf2_?N@E/A@+(,6.+
&/0SU0_Y#4;5egb&B]=K->JB+#:[_0@dOaFX:&g\fL1HW0g:DEM(f)QR_EQ)K431
_>QK,Kb27P.XSJ.7C]>V:W(dLV+X-_/e8]I2G)K]K7LIZXA@8?TJY-2F4O.>OGa5
4.9?IICeM?a]DW]:^:b<-R=BEA(E#_X)[:QG]+9(U8Y=<B;B[KdZcaLP1(\We390
VNe2AATZF@b=;X5O-:Y2V59EH>-3[O]EWMOALM6b6a/,A]7D.5,MfZG(2b7>MA]U
b81YAC^YVf3(M38#:1a,g5K>OSLPGJJZ9cWReFg,J/-5VXa=M\Z-N=,Ba:):29C=
9>7+)FLC3EfN8;,Z]C/HLYP]-KbGK7NXYV_=)BOOb@;d56=e6?14UfF4K;XM>]#&
>.G)1,O2Pg8@fd,J>eKX2[TAQA.L77D3A)D#D1AZ(4W?K,Z2S#HN&=F,^?07_)^G
\#Y0X.+DDB64Cg6+fD@/caORYTTWbPR:<W_g9-505W]RNQ_CRIJ)J1B;]@adIIRI
>a&aWA?7R=c?@A0EX:fI5K_^B#N4,Y32Vg&GE20ET>+?@@gUYGgLbX^KE<UCE1,.
H;V]TBO)eQ&;-O2c(\FGbBJOV?[\dE>.gUMQ&//0f?^<(19QEL(LFf8LTe^a,E0&
]&R,ELJJTOQ1]H#a/4PcT&7E1<3V?e(5CDTJ,3OZSS<C_^aNU-:a]5K#4^C[+ZKQ
#e?[G)YL4@BXdd1JB[cMYL40VI8<_5Y;8Y/?T=J,O^KeS8]GD]6gVOG-2)ECA?-c
V[:#7<V:dEY9PgOFAT4[G1B[F<dE_](dd_K2Z[aLW?e=OUHYbH>QdfMUQ+dUO2Qb
\[YXbK>&2S-VJY?8TFU^9QcVP.);Kg72OP<8c@ATO(UB,:Y:9A&9gY?#.R0MUO.9
HI5QI29.4)7.R^BH8E-_b<<Q-.-B7NaN)R0+1aa;;LH+/f<XZPg=H:\0YI-4=9OM
JWRPV=4>39f;K#D[NZAW?+]F\81Y1aM^S=c,34NTWf5_BXC3e<R^>AW9)]R1@PaA
D1a=V3e^G@>d,<XVSb9H&C;T/:W?6Y,-#\@(ZJ<V+G)/4+daCd-d&-U5-SZWOd_#
:RSPXcDC;/:N^(&BfaI3(O+g1?4NEZCAHNc-T=5T+W)&NGZY](:1WIHG_^PWK)bG
9;+dc?d:8ZVN>.4[a1?<eZCP5O/=G[Zg/P<)Nc[_1@d/\CDV@FTYU[cB(_Z:KDU9
IUG9LfU5RTEG)J2/.Td@@[TLJ=NJ\P3M^bDf\b#5c-UDRZW(]U<GYc:,e&/96[]C
F^8FIPTS0D\]E<fR#F)5_(1M_^?7WP1XE4Ee,CbEdd)78A0@RW5_J>(N-VZ]SVOM
LgVBOUFDU-RXU[>)U#@JAWAYOeC4KfGDgL?33OIH2G0WQe0DJ^bO;=/Ne+8UVT7b
<a9\aM48[]KgT4N7<W1;[5Uf[dZZ4dG3>6<1X0)HKMXR^B.+=Y?MADNU.U?=FLPe
Pe8SHEH-S0D[fHb2PY[Da27QAPN_Y<CN6_3RZ^ReK2E7B_E,GYSX.5Z@N5a_-2>^
TNIW3K-8YFaC^.N(=S#@HSSOBK0XGZ/T@(PG\dE.KeZMeSRYMPC:H@8.-9fYT?8G
g8D,eQU>cQ_0KB/+=+B5DQIf(3KCee,SN^.5I.eH,\XN=cgZ[=/Y2;5HdB/.@dVH
_5AN)]M.YW4S2,?#X6a6J^QDH7e3a<UPGP9Y3H6&OWR(3\E2)8UUZIKG#:@/[daF
1D9e4B&OFa9M\8d]/4)baD0B^<cI-MX\>cBQ43RK^++)=QZD_Bb<fAg>=P&3N7O9
aJA1EX#SgLMN6W)=M4Y[,=,URR2E6eY9gf;1(CZ4V8L_T)J2+SX\G^bX=53X1f,F
1g\O+Q#6>,-^?^7O0BKd/C=a1;RI6I^B77(O-AZ.QU@cI:ANaSE4(9^gKWA&N55:
ZU;:UZa/@5A=Q&cgP5_3dcVXQ<21J+(7].2f.\0U#E8-2eOCY/_-Z#WIDLK(eBBP
,Y<>5F,4.,#Rg<#,9LJaG)&dZ[e6>Z<L:G:P4B5V]1XAS;gHLT0NcK@,R,LWM@N:
Yc;f^F&eN(&@DM5;9VSY8-UW#S_c@CFVX1D6+_]YJF(U85WYY:6cHH@Af@ME8U49
D5VI&b8)9W9e?42c0c#@A\g/(FfYQO4R^bT5JaM[/RaTW)KO<68@fcF2_@GIccW5
_(:[\-;DfRWdGB?QO<^&,<E?H&7XR#0Z<8?9IX<@MZG2_>XPKXK5M4]GUDOb:Sc@
4d/J))ER67]V_IF^I\a:>QNI/3G0c\K>GH=FD1B,X73)TREa7+VegH6TWbX-=<T4
D+(_8Y9+SC6-3Z.PgBX;aPf:>U>PHRUX-5]/F+b;DMCdQIZ8K-L?f[[g[:MPIMUE
R11CA5(M9SM=>c_60\bTTgOdf-@[+]:LSSRg6^?[W<CJ],=VceYY-U,;=YT2d\A_
P(;<gL5X>I=e\Y1A]9)>6(K>(KTH-A>R9D3S^c1)g/;@)SH?e+OU_#a,>f>D]<4R
5dYa=@F6^IUMK)(S2L#XW(&..F?17MI&P+MY8aeGOBf?T.?1\^E&^1gCA>07PD^0
ZFe(0@]RcM-XO;#PX.dXY:Y/f=4;f3SSgX>JV/.4N&JD?EJOJU2:LW9PD[>2dMF;
H[W:?X_CU7NBF.QL6e>_I\DgF(=<7O2[YYS7POP&V,^T>MFf+<6I_C.(7USDg@g_
Fc8f<1KUbaBWT/4UZ(K9ef[,2^43&f[_b#fcUE-;)K8AcFIS7NbHYRaS;H\5Zg5<
&eS@6-@SV&3-/ZFL8;;Yc]F<G;3:+_8Y37L_5=<cKFDDK(f96</G/2S:85Q5_4dH
Q>CZ+1deD?I8K.9CBJ?AJ7KbR<&ECG9-MTFa;JTM:EF=]QgPC><13)+;EAZOHfOO
SHZJW<Sd)FN66EJMLKaB2:8+K\[72&.8a<.MXT/A5,We^eB<&2B>\#eM2OZB]C7-
gWeA1+V4;Vd]c=@LR\;e-Z3P^Y?&9ODH)ORQ5&RHe@1[Jc3G27]IF^[0@O9/=J3R
;eR[cR_P5>\GMQ9#383SA4VHfcAW+Y)a\E^FD<4?gV+d-,<O8B(f5=ANYX_?D<T\
Q7-^f:g7&,JC3^I60A=dCc8Wc_#4U/A1X5R1M9#&feQ#5eMR<Yb2?Z:;][TbV,XE
9/CFFOa7F):\S\L;0&#@OQgXS8:MTL[&1G.M:6/CKg2)O653BLf^(7d@]#/+IK#g
ZDVZYPX[LGJI@5TND#JaEPFG:##;YX0:X]ePEV_#Y_D1<MJMG-)250Q#LN)1gGR(
SL6]BE/D;B(U2NYC^Zg>L4,RYGQ6=BQ_/GA>HSHLIaRAS^_SH\c]2>Y9&J1V7cS/
ea8gH&0P@303)1Nd)?@Qf;KA@@;DJ_22eZ.9dTY9_9W:3^QH@-CRLTgc)+4NfbK.
dRI:a@8^D?L7HHH203@0]NcHc_N>g_bZ1+AFKMPX)345,=SfHN>>\LFO<+.N]E@d
X_<R5]>0b)T#.6F/g\?N6GX9IKd8eAQ4].24#fYDD=^ZQ66RFDP:.b3g#5\>7FV3
fI(KYVV)W:J@<N>2ZNbA]WH??S+YHfa=B=GWFF6AafaVO-,N)+UJ;,>_fBaME3/C
,bbbH-L6_,]@,J]a048\+3<)-KFfea]&A[U2g[V:9fF^F\CN]fT<4\Qf9.=fKPG.
bfP523C\-R(;]]+HgH,&UE,g^;L^g+#c4@)7&<)_#-Y-[00PS@^6[b?-//N\G8EJ
E<I=MM=9NRF&X+5E5F7]J-bPPRXO-,E.N#@ZH.M67VXPX>G;O]3>cK>UUJeWK]8D
cE1ba4B[Ua_,(.>_TcY3FB,Le4)10d@+_7Rc=[,XZb9VLP9Q00g[0QPVBGL2cWVR
3@]:LVR?Zg.2_-+]=D#@>@+Y,(48V80,Be^_VI4Lb5b=3@O3]N0e>U_XEeR3<F[6
<SRMb?5P>+@)ZF(G8eKF9;@1NBL=(KBUMJ53J=.aJcK\a14BV1Fg558(/#^O?GIT
HC.FFE-cH(<5dX1d&BP52=fQD.[F8I+7B(Uf34R3Jb2M?+2=.>EJPPEV>SVDDJ#D
4MQ0be]Z\RfM^fI;FJN]::K]6KP9LdB:,?+eFXOU_Xf6A>GaNE82_d,BNV;+=TM>
K@,;7C6NH6^f^d1(VUfbDcUdBD(34;9^Q]g\[E7G6AGS1cIa_Q./U]Z-8d2RI[R;
GH8agQ?A(gb8e)eZ3M?SAR#IQPDV+[\bLYE:B_(.H;6Q?W.?PXD(LV7Y+Yca(ZOW
.^(Vc1AB_]E];GL2@9Z:^E88VP9VQ-Q&NY->WMN8JOQ##N6;N.3(;OQ0H5&PCL@#
EKC/fK6F82;\3YQ,M;T74B2aHN:Y#H1WOE;[0&;c0_>FEfQ1,BKb[A&:MEJ:#>Sa
7ZKTS:.=>L0EK1aR-Y78DD6BB6VI)&Ma=>._;V?g37?Y,Y0P\I1WfafMe69a)I&9
eXaVGAe&d-CO2OXceQ.RA4VZY@[^+4+(>2J:Mg\A>EIeV\80UVFDBW5>S/_Wc=[W
D#6@@V/VE.V#4_dIf55@94f4^TOgO&dZ0>78:,SZY\Rd3-aR(,g1HWT>=b]0R-B5
IDTVP6]_eeTK&b=S60YY?23)M7CB_\4&W;4+b;cC_1>NM#_R8TN_CJ1QbS05XJ7-
;6<S3c@>L\,U\&?IW<IK)A65-5WT4O#b?:VCQG8/M#WXf3-J61MI^eMPd3.a/J2:
NY1,3;gKe.J#2Y6ZA0@W3b^=B(0#Q4fW?Q1S&dc@FdPfF@4T51Y8&KGE?4QcHBR,
IOWBcPZTJ>AeN>O,W9Z6LeAB[U].e1dbW/^(7H7#IG_&#6JI(:^?B/P/f/OG)X0J
P=T3E9N9OX>U53YUE#C:TPRD8Y;[LKE5aN/Fg^c]T@/3BC<_[)^3?_7/&8+@KSTV
0P7D;.PO-;IXBT2aXD+NHFIE:@#3(HUOP5GCCa,EW_VAJC1_;C#K?U/I5\UX:@ge
V7]<=^YaTC)_ee^We14);c-Z=dMTBg,GUL+R5d6BYIRIIPD3A+W1@1-YA:6^VK+C
6>g@@4922OJQcJM6IT><\7L>a8<LdV2;f=/G:b>P+^1^>Mg)Z=^->:]2JZg7,#JV
M]0=URb,B[dBWJQ3G;fF3YDG\;2(1FPa=HGg6^I2M9:G0E6K-0[=SP<H8+ZK\.a[
<L7I);T1,LZFU]\F@MZYY^4Xg1;^bZNEebF\HXagS?/0&8IKC;-S<(+[DEBNKUa?
&9CJ6MV_9(XL_.X3(\-YVK.)D=F/+7^^B]H29@_>a)8N)55FLK:Q98HLL7KecUNF
DdBMV0b]8H[g)0GCXNA2Y^b0+>25:PTbK=d@H[FV&Y^DWO,=T]:2Jfe7V)c:33C?
AY<1GT(aD?G8=A[bI^c;dF9HJTfA.?WM3g#7C)[XGFfFT=SDXaM8IIDa<;0c>O3b
-P(1dHB>_&be\DaOBUGd=R=0:[44PH;cRF3CP38/9fDTUG?Z^)2MJW7@[;GKDTYa
S_]8V/KN_O(6KN9)e2S/;BMO__E5>YFD-P(XU#L=VKb,AML/JY9VfR#7V1@aL)TI
&NV^MSX,T<^&:=R[AcW)WW.GeOLW@IH9=DMa0T>^WYV?1#^6J5QR+f/c^D]dbMY^
BSf&LNcaXF9aH;?M7P,78KgC+((gaE65?<4X@1.TO)X@>MTX[2gB)2fP;FN-K0G3
BV,F3I_7fY]61-MM_JR2UIDcSgdN2,T&#U\#D7(a=WW)V+\950^TYgK]12.KBPX]
6?;>:,6c3PcDO[fDM,>^?f\R?a)XZXFSdBbP/MaT)_A\gRO.]5eO]?SZ6S4,Q4?R
,[;K@[+/:/^:_0.H4@g4<<./ZZGWTA3CB-,V_UDKU0KfdA]@KHA0(&IZX\Z5b_c.
Td-]A?3UAB)2V0A2cfKdBOGE+XJ1MW)F4,H?DKZJdSH&N<DE&.;c)Qb487R.\A0T
=ZY.=EA=eM]4b,PB(&@(VLO7PSF^WN=#[R12bfGE-_>5/SBW;E272_^>[DNacEOQ
?17g59JZd)4:C=#RW>YUY@2:;CVK_M1ZWCF8gLf#(]b-_#+cU=EO?H\+/c.JNOW8
/dWFIa<^Z[@b^:\4YIS5&Z;(=2YYU^-=Db7QbM)XT09CCRR+9I3C/c>HY&_8JNLa
W/S2JDVaF1+=Yb6W#W8:HN>Wa6IUdCI]We,\WE3(ES6]082+><^X4<->BT>cO>@A
:FgESTg\7Q9^:,.\GH0.7I:-d\=DJK(DC\32fYW(8DEb<ZbKIT&.D,KJIU6(8@6_
3NMK@+Dd(XA0[[#0/_GI>g_B0\7D,MfF-1LJ#P?U[V0YUeI/&,(GI?Y5J8TBZaBJ
7/DATP5CC+YGKV;=GG17W\V6>GcCA909d<+963R2a(f3EZb8#G3FTeEe[C#<[[\D
:c;N<X<,E>2/&eJ?CX[WQd3B)6:(/@JLT,C2)H&1P/-EXIH3Re4,8(MO=9-,ZD41
BVa?5ZN_+#;[?]?3Z,U[A9cI_KFKcUE/6YDOR-JOB5ALPXT+Q8P^L@09Q8J)1(^N
P1;EcdVUd;/QAN>H23MRK;@1?22PG;+XIIDJ#c+A@M02bA5F&A[TD8<+A0S\YQI2
U_6HKaX6He9HGQ5P&)M,N_:U\We,&,0^=;[0a6<(^Ng7T^8Y;9((ZDTfQPd)PAMH
)CQ4^ZX3aI/BO/G]\XYa,FBfIJH2WH<(:S7\]3HXAT1&<R-Y,#JPWMRDUB50WgN0
6\17@)LH1O<511@Lf9dV>Ug-Y+:9SO;28@L)ZD[DIec<FA2T+5-9_^,[>W[9,ZM[
]OBKNR\\ZSHF:+38</CA<d.7@#=O\g)Z?P0;R7>/LPZ&(5R-5B(6d_U+@#O;Scb1
(82H@(;\_Rc7/&7#?M/36#BDMS3S_Y_);3e@6]Z)L=/Oa_-@^+_e3:L0;WbE&E6O
VPMJgEgd8Ue817?<SW/0Ga[c:@J2O\?T[/AL_dW&Da,<SD=V9\S^6BG&K5g8]MH@
LUfVb?aX@&@]M&+&_SXH5b(Mf&Q8G&0TR(9/^?4?>;/^3]#ZBORCOQFa?cH;WcPG
#I80D0L(\J@aC2aUa@E2=&U.MDK+5gJ)B-M&ZeZ4CAF?AUP&9W+X/\U_N2(K&[)E
J>Ra/77O^>DLE+2L3aW,>Tbe:G=[B>&[Fd22WNZEIPW#,ST/K=P\?[=SR4/89cSJ
U2NF:Ye2PGUZ/F:[2O>-5>YFNV.C:g/8Mb/C]a3XZ.LC+#NI-=#&KJHG[PcK<ebX
a8;8U@;b]B7?>)^8RVA<Z-MNKK]#3^TD4(e.RT.6#eV#PNR\SVKYR^T0KHC7#<1c
ZL<+eOS]A>OXIYRJ/XaKgXQZ;C)&E-PQ_I(6ZQVBR9f]T,8XJI\:P:L7,]W?7H.,
SO#M]Y:OTSOF,50b6&bEGMGf8FGEKe;4X0@M>T1FWc<(aN9b?\,5Qf).4QZS:8L>
^S7F6K6D(1EMgZg6K_+UI6DUV:8<_XY,@RY]&22CZ3SDCER<Ye51P/:ee>=HO@W+
,8.1\7>OH7:NQ+g^-OOC->UE<9@J0M,8RD><8XS(_FWeg.P_;:&9)N/_26P>c3,O
&/52Vb)V.3FbM6P4^cf(1#^P5:<<bCGHR2c8^,M\SA-7_LIM=/I;AG?7cGc;&dA>
KC)RM4=SLP0JPQZ?R?aVJYO+5_aNAN+f/8GD0THVEU,:I][N+W^6>S_,C8d&dN5V
9_D)4--:]2I5<9+P-,-Pf49b]Qg(Rg8S)g=1MTXd,JW)+BL.8a^7N)7L569-eYB5
?EL+M^>9caJ:110(GU-FaH&Q23,8#XN,-.-0O@/X:<;:IRWa=4Bd\ad0_H82&Q6U
L7_dW#L8b6f_?&C38Z70,3:c3BQNL/]7</Ne@Fc0B9I\\4@@O\f_)I,J.dZ6fOKA
=I20U_5><H(5Z]S0@V[[F-D=;/KX2>JZGECT4?I_IR&QH6LYUKHM1dR,Tf&/]D.]
D::Z9MI@SYOB13#MQdH.&IgPNC)dU>[VM\KAe^5,D]=NC/^cF[e_;V[8KJ2?BE?.
?N?B_OU@NJST[M@AaZ05:7gGYN8)Z=Y_7]e]4HUX-\\eV+&D(.AefGPa#/VQbg8I
7NW4W<(OOObS,5B,-<LL(_MV6IU)(IgJIgL-2;).&Z.X6YacBIE151J95=#)g<@-
efQANgZeZ&]FJ4cZ2,\7X&;E)\Haca?6P<L7+:4Rg1QHCU\@JT1&]PE1PW1g23<L
KceKW?GPEI(<+#J0KVQ=/[<08g9+6EX>2(ZX>0L++),?eO5&aU[J5/<=;8@c2?&8
g_FV&)f.FTT.eJBAZ_(A:]EfeL4UBCa;a5BCE5,SXXe6(\,[IZ#Q<A9\bc0dcT1V
82=8.ZQG?P4]8<Q8Id)J5:E&>Q7H259G+_cSVP1WX\IF6]^=dR>c+6@]-CM+=M,b
.?ZO+Q(gU&F5P<V14LQXZ)XQ/]^8KU+.N&aOO)>&FH1GW:ER-XDQJ.fC^c-A0/7T
eUK@_M/FRR2YMAcCA\J3/g<aPVd+b12X2JW^H88eT(6O<c4P,c]>CU^PM#e_.1U@
eCB\?F\X]d8;JRYT&=52]9/WFU.)GSN\Q8-WR?:X;YRd<_@1,S:aU<S(ILCOLdZb
B0Qb0Gg(>(Z[^^F7W]aCTQ#3W/Y\L.59(J9/6K@bC0GKeNd3fGb0CTPV(gC,AQ_9
4Vg>\<gLdDe<@Lg7W@K=GcCT&=&AQeN3IXf^:9;OZ]H#1=MU<0;07<M4G\YdR<_#
aEKDY]-=.@.8^CaK4Cf5+JH1).8=7:L/JKZNC]2Fe#@&O5IU+T-HeE19_D\HE3MG
Ff]6Q5_VTK&Deec5H\.@QY+1H8cFb3AOQAGGUfg49GQbGGE75PG9?=3F[1:YLYN^
9UDfOZaDO9H]#>7H=fbef6g9SFc#1C\&(dG:FUA+)WI,M)&G>Z<#d=ZWLZ0O;3@Y
BA>CE8-)L(LDR8TRPJF7EZ9T2#TS9\3,;H<9d.:>P[\c@a^UNbSHPaP5+\5V8aKV
P.X7;CG/eL?AK\\Y79^Z?4#,GQ9@<6W)IQ)4g4gZBQK[Z(g;4B))-6c#c(RVEU5;
,YD0>f;C=A#I/U9UU1fZ<a,:S8fPH2@V7dCP8^]W)=URK(-]E@NE6aAH,Q34HJN-
O0#4JT3S0F>;QZPBVK8,(\7.);\/:U:H@J95U<?EE19?fR;.0b406UdgB#e19d;?
=eWJZDfY:&J@??\3=d@T?;91,W8b2H&:RQ#&5(d;)DPg<0;c@ZAa_e>S_?dTJF&O
gI\Wc:.Gb\14YdU2U+W6MCdg<<_:ReJNAf_53G?Ub.>fG1T)S=bAgBX.;^J6YW#9
CJA\7:88Y:?VY<dIOGE22Wb(VfFB0F:KV:@Y:.,d>bR^cW\TG:I(R[\[\;B]1e.4
@:-.GYRdJ[J:U?5NSe@@#D<H+UB/NVE(gZPRbW:(.B6.B\+Qe-SSADJf?D@]Z0Df
_0=HR;4cBE,@Q0JXAE6]9??S)RI_be32+VJR&.A]_T1&Wd+K2UW)<dAX?_)OEOfS
+3RUS1\83QcOP?A@\[C_H[Q?LZBHYON3\^H#5F^R1NIMZ=gH^3@Z)6^dBHYIA]ON
QB)8-]A0Q+13F;434#a?T[<\.&^Ka/NBP3H6g^SQ-C)-0O1)6Za\P74BRS?@cACZ
0\b)+ag:c[)WRH7EcT@_cM#^/48UU]I7,0<T\a+(KSNM/eeVF+;OcFGAdZ7;f0WL
=G+_XP?5N2KZU\23Y^d,.^c.WW_0g&V_JABg[fd0@O5eEO@O<40(,C_.6BC&].[I
B2T.dHXDY9)bED0;K2\+b6JTJ<gBBDbg>QSa2&X,Xe1@YN:E06_375KMU5ea.-H)
A#HSH0J#64+UIF/#,)JV0A:g80;@Y>9&OW\L8M\ARJ4A./e?(>H5a.<WcR/RNE,Y
280G#6g/F-H;Pa7GY]:_bAN@eGT67O3GZ&)YgF\SJG9C2bN<VW,SCE)A&AEg^O#R
:+YH:C0K<-?PGI,<g+]7KQ,g^VeDS&1U&9+:@ROcF]BL4I,PS-VaS#9d>QSKJ3@G
W88aNOLIf;JWML9PN2eVK7cV&UJ4Xe]=aV?N.E0X2(^?d)U>(4OcJITb1>W3=O@N
eH=eAM45^^H2YfGe94P:](5B/L#Z,#R8>^R(C-_D;FY4M,QG\F.I#4ZXT:;6I68C
1W3Z<(V:d=-eN)7T+?IIafU(=&F/8Q-a?Z5d8#aPWb3aVZd?)#X8?D1-<Z[SP5ET
;T8I8Q;]PMFgdB(H4Pb\&K;B6UAb[d([A#E0EBPY^ZI+Y<9fQ.SOT,5+1da#_9FY
G;8./0C,&>:QUJ1Ff:)T#:FMRDK.-P-cf.C:(eaA(;GNDGge&-7I)7TLUfMD@KWN
E.adagN\eM:9;KB4?E/[\EW?c>.CY9BG,DB;g0RE/99MZ.VNDH).R<86?/1<.SEU
,gc?(L1YY@Y8XeA4a#[64>0c=a@a^)Jb5aE^O07UW_S?e48)EDJ:J@DZ:=A.62#a
9;0XJD/c8e.#9V6[72:eafXO3)LF5K_88Leg?@XK+&<Df(;JC#G,bCTOHJ,W&T:0
>0ebH+/CJ,Q#H^.L1B(efI5(F4-b-81N?HR5L2-0C3HLP-B);WMY]),R>XHf57(5
3fWZ83R4/&@b7,:8VcK[cN?a=0\2W\JV^gQNKCBd;fHHg,6O+4QNS]@PN[28eN#D
UA2V(6+FV^(B276cM(8&3(_,6U7dO/)7_7@51UY)IZL@9PU9XX?5K>\HQ:-;?A>>
7VK7bN-KfH=RG,f6:M(3UT^OPfHWRb:<ZV>-fHX:[NZ^A2C>bM5-fB]0@+1,^A=\
5aP#3g?2B)ON)P5\[^T2;Ze?^U>bG:Z\7NT5<)-b_AgDgT4#<2+,E-/CHQ515VL>
/bEQV]Wg3(O>+edG78D-cOH3Q<413Z\\RD6TXP&LOV-(-OdQZ67_HAXP0b1=2G(U
8/2A@eQD24UXTd(;^J5OUM:G5CR;?M0)c&7WGV1//<=24\_-,9_Q\6M)ga3>];/#
#\<,(WcD#a&1RPWGbf7K+::?.S;AX05M+(U68W1g7THD[a+D7^X)[O3KM?aXP.&C
<UV)=EU+,Ec>W\E3V\P6&E:X19ZM-BZeVJ1:=(OI7FOJ0\\VM65@-]=2\O;&/A&)
X6Q7)M_&g<(e<UY@[g9]C6g>L^2#>d^\L\,?2M7:\CP:WX5bYOGeWJ4<1,H^W1+X
AcX=EfZBSC-GR]Z4RG^?EI#g=/F2[1T._O^+Xg@cG3EBN#Q2E0&eCZgDDF<UY[)f
H(1749aAGeZC)HF^S3-4=HfV^^c)D7XbK_C=CNP.EFJKKI9TIEU<1>O;P62)DU>W
bg1Y.V/dD@T7W7CTbQ7/&[&JeUf>cOW/ZYJ39M,a?XJX_/J[82V)K^_8EU^6.I.M
e::+D4D@c+DJAdU^6)cL_<N?U38=2a-8(R,:7]a=A-bE56UT8W1g6X6@g:EgBIY2
&OT&I7AC\;N^&WEB(?]^/f(P=F(^>,=B[R2[\G#@1GB+UB5P@AI?L7BA/54B[RPG
&-EYNc0[:fdC(bRb@;g7WN0?,>cA2#X.Q<-T8L.Z19IQM#Md;9(A?^\Ga[T;Z:MW
=7V3/g@:P&[D(-:RQH/9M]O.d,@d<D7B_a79L>]#d9&gX@6-G<L^WXX.@R1]8g8&
PNB-31H.?faA=-V&C(aIDPdeVVLaEZP5F)8UQTBJO>MA[d\,ZWXZP56X7J<Z4/M@
2ZVg:8)9KOE?fL7bI:R9[M6[X^^BE37^D7@X?dF0<O?3AWZ++(e1_WWaWY#M04=8
15MeN\NddTc(Y^E;;e7(b)c7&K^[J\dFZCZEN./aTE[a0D-Jd6?QT(M1EZ0R]a8Q
2f8_[YV#@3D>&Y]2+UP>^KK]0(H[=Y1Pag63?;0ADJ-Q?UPV>OTNF)-8)V&)5O)S
[6#1A2^;5GG]I-?&@];@0@55(]ZOG,cSNF[7=&N<9&0dASQ+[HX/\dfcCP8W][TA
67:A-(TDT#8ee0#E2#2E3&IIA@<HO^5R1J_)8O@\3C+Z&@eM/.U&1WW,?;N_1dg.
,RW933<AScIVT6G?gV=T0fP:aDOe6d=MP#ADC]R>>VSXMP[:(J=M03O,LS56I?GL
<B.6aSHD_Y<&=,3Z,?PJ[:]VO^OaeE#^?LcTJ)#8_I:-8NCL=(MC1(=feF7O61.0
K;f,PU]bLe+C6^IOa5Q:B8II<JLG[-@1dF\R2WK^Y-PG=T/&M\)ffVf64/NW,47J
0E0D2.56g:E],#(3CbF>bLM+W/9ZXLbdR(.#+\OM_egCgc+K#D;-,JAL@S@@X,<(
L8]^YCTQS:/Sc\Kb4)/Be8bKT^B9e2HXP@.2HLZgY#].S4JC6?X;P=X60YA9Q9BL
0ANZeQ(,FN-I6\\^ZZ-__-T&,6FOAHED/WWBH_1dgac-03JC?TC7BU19&cfefKSc
d>HDY:9>#UTC>0NCUDa1dSQ@d&CfcS>:Z2OfDS5E:TAb<6VRO:>)RU=<X]bf.A)-
K^2Uf7L51=c:[H;-F7Y3c^U]<SdDf8Q7BBJ#,5\#^.&A(<)8gP_M]@S-2/F:ERa>
/f(K9=4.,N)4&^\+gc^^E8B#(HMJO-beOA>IHZ#2H^:J3>4#&IGIH3Y(0Z2.S,YX
_D3+Y6Q7L7bVBKFga(=#=R840GVLV?IdG,],^H,J[67Y/_J32,>V?I>HR3<UYZ;U
1IJfX38RLd/<BcSY0F/-3cO4H#8UP@Q#e1LOONAW/b4;-f:#B;.,QgF_?/>SFAcQ
P&EKAK5_Q0g7VL-/WIF,09>@6Y0Z97f23?R+GGDK(#L=;;MS62#5Z5LA/.<NX?D\
/O)-W:.TZJ\dW(-Z)78)80b,2Rcd-KE;Va4^@ag4YQMCJW:8K]R7-MB0ONa_5[,D
4)OL8L=\]FHB8S_=:D9?;b]?><IW\NY#9FF.XN^f<KZJLHO</.<8:JLJYV&.O#.T
/Sd7JJ[W,^8/NDUT[EU,[_8[bNP23BLME@I^JVO&_<F9\-Z/;D+E\EQ6&FaUU4V<
gB_[P?#caF.-&.P:-1.RJ:Q=#_2LK^H2cQC10X&A9C4JD7Z(W:I4KU;0CI)7?-,=
XV0R#0K.2LWKQ_X(f7/;1X0-9O3.edgC2O=HZ.L,+:>/@EWS1VQDZ+Z7d/=>E)aa
\B=Q&KFA+#9.FZ6=RFK19[VT<#QOFX14OIT+.4+??N/Q4:3S)@:;HXZ;][,A,0-c
+JC6NfHZ_X/&-O8d?Y9/F9IN;KdBbJ83FT1CQIQTU&^]6fO^4B)B;)1X/2Z)T?2g
D\]DN1?c<R0[<CgD;=gP]#QQMK1;50(gAQ1227\d4EaMG)PSDN765M+7G5-0\I&&
4-AHXaaOg:VTe/.[+E1_Q.XVR?WZK8b+V,FP,TY,4]4_65X94D]EOb\(,)5K/GV3
9DR<V0Q?7ZcT-$
`endprotected



`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_slave_transaction", svt_axi_port_configuration port_cfg_handle = null);

`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_slave_transaction", svt_axi_port_configuration port_cfg_handle = null);

`else
 `svt_vmm_data_new(svt_axi_slave_transaction)
  extern function new (vmm_log log = null, svt_axi_port_configuration port_cfg_handle = null);
`endif

  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************
  `svt_data_member_begin(svt_axi_slave_transaction)
  `svt_data_member_end(svt_axi_slave_transaction)


  // ****************************************************************************
  // Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following
   * 1) Tests the validity of the configuration
   */
  extern function void pre_randomize ();

  //----------------------------------------------------------------------------
  /**
   * post_randomize. 
   * Calls super.
   */
  extern function void post_randomize ();

  //----------------------------------------------------------------------------
  /**
   * Method to turn reasonable constraints on/off as a block.
   */
  extern virtual function int reasonable_constraint_mode (bit on_off);

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object used for logging.
   */
  extern function string get_mcd_class_name ();

`ifdef SVT_UVM_TECHNOLOGY
  extern function bit do_compare(uvm_object rhs, uvm_comparer comparer);
`elsif SVT_OVM_TECHNOLOGY
  extern function bit do_compare(ovm_object rhs, ovm_comparer comparer);
`else

  //----------------------------------------------------------------------------
  /**
   * Allocates a new object of type svt_axi_slave_transaction.
   */
  extern virtual function vmm_data do_allocate ();

  // ---------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare (vmm_data to, output string diff, input int kind = -1);

  //----------------------------------------------------------------------------
  /**                         
   * Returns the size (in bytes) required by the byte_pack operation.
   *
   * @param kind This int indicates the type of byte_size being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in a size calculation based on the
   * non-static fields. All other kind values result in a return value of 0.
   */
  extern virtual function int unsigned byte_size (int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Packs the object into the bytes buffer, beginning at offset, based on the
   * requested byte_pack kind.
   *
   * @param bytes Buffer that will contain the packed bytes at the end of the operation.
   * @param offset Offset into bytes where the packing is to begin.
   * @param kind This int indicates the type of byte_pack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being packed and the return of an integer indicating the number of
   * packed bytes. All other kind values result in no change to the buffer contents, and a
   * return value of 0.
   */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Unpacks the object from the bytes buffer, beginning at offset, based on
   * the requested byte_unpack kind.
   *
   * @param bytes Buffer containing the bytes to be unpacked.
   * @param offset Offset into bytes where the unpacking is to begin.
   * @param len Number of bytes to be unpacked.
   * @param kind This int indicates the type of byte_unpack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being unpacked and the return of an integer indicating the number of
   * unpacked bytes. All other kind values result in no change to the exception contents,
   * and a return value of 0.
   */
  extern virtual function int unsigned do_byte_unpack (const ref logic [7:0]
  bytes[], input int unsigned offset = 0, input int len = -1, input int kind = -1);

`endif // SVT_UVM_TECHNOLOGY

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>read</i> access to public data members of this class.
   */
  extern virtual function bit get_prop_val (string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>write</i> access to public data members of this class.
   */
  extern virtual function bit set_prop_val (string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
   * Does basic validation of the object contents.
   */
  extern virtual function bit do_is_valid (bit silent = 1, int kind = RELEVANT);
 
// ---------------------------------------------------------------------------
  /**
   * This method returns PA object which contains the PA header information for XML or FSDB.
   *
   * @param uid Optional string indicating the unique identification value for object. If not 
   * provided uses the 'get_uid()' method  to retrieve the value. 
   * @param typ Optional string indicating the 'type' of the object. If not provided
   * uses the type name for the class.
   * @param parent_uid Optional string indicating the UID of the object's parent. If not provided
   * the method assumes there is no parent.
   * @param channel Optional string indicating an object channel. If not provided
   * the method assumes there is no channel.
   *
   * @return The requested object block description.
   */
 extern virtual function svt_pa_object_data get_pa_obj_data(string uid = "", string typ = "", string parent_uid = "", string channel = "" );

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB.  The pattern is customized to contain only the fields necessary for
   * the application and tranaction type.
   * 
   * Note:
   * As a performance enhancement, property values in the pattern are pre-populated when
   * the pattern is created.  This allows the FSDB writer infrastructure to skip the
   * get_prop_val_via_pattern step.
   *
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
  extern virtual function svt_pattern allocate_xml_pattern();

 //---------------------------------------------------------------------------------
  `protected
HB+CF-C)O5MZ^??N85Y7b3,bVP1L(CbbSUWcM4XQ0@LK<#7IOV=80)QQ75^@/C)D
:E<(BfPaG[FZ.$
`endprotected

  `ifdef SVT_VMM_TECHNOLOGY
    `vmm_class_factory(svt_axi_slave_transaction)      
  `endif  

endclass

`ifdef SVT_UVM_TECHNOLOGY
// Declare a sequence library for this transaction
// -----------------------------------------------------------------------------
`SVT_SEQUENCE_LIBRARY_DECL(svt_axi_slave_transaction)
`elsif SVT_OVM_TECHNOLOGY
// Declare a sequence library for this transaction
// -----------------------------------------------------------------------------
`SVT_SEQUENCE_LIBRARY_DECL(svt_axi_slave_transaction)
`endif

// =============================================================================
/**

Unitlity Methods for the svt_axi_slave_transaction class
*/

//vcs_vip_protect

`protected
Z(69aKFZXN;5KUdcL=<W4C37WO(HX#P1IH\ff#6gg<U/Ac)NVWRJ.(b?9G7RH6R^
@#E4QDC)C6-OLEf:&T>1;9+=V1NS(bgB,.S,b>]9GN:d2@AV+Wa#a^ZM&aCJC7b<
_=C_N/NK=-&3;19(M.S;&BVacT<_E+c20^[\2\e+^R^>,YXCCAG)J^D&_>?[0+23
.,+J@)a3MT^G@\M/5V)J0X=0b2R5O8K+MR\4G\/FB0)]:50Y0B^1^Cae6LAg4>26
(IH]=]0^Hc,3G15^^[dP..T4aEcD::NAOG8CQL_TH?#@DQ6G[ZTSZ<DgdGb0E+5U
1f?II2?L5\GKOaF#N1g9ZHKNY^W1AJC17E9=BW:MT6aLS9F?2.H6B0UP:3ga8OW+
ac#HYL>X?=SKS>C#\9U/8;8V4?MVL0#aJAAVW[cPVN.>UBJZ_^R(Y/e8A7W_T,gQ
\\PZ?.3RAT7ed]fDVAC\a6L]<;fH81MU5aLd8aa.?4.KQ,HK/#c.?UeAa4\F/(SH
/1=/F/\GPe=T.aHg[:J-X-<,=8-\4>\Hf0Y4G90<>8,-U30H,)_9)ZNL?JU0IB;e
D?LZY^cYB8S)>d<P<dSKKPP=E\UQG3W^WeBTb)=(_,HRET<c3E+#4]&1U>TKH.^;
T#89Rc?(eW5cgB@JR&-YM;/&ef&O2@QA;$
`endprotected


// -----------------------------------------------------------------------------
`protected
AT9bI@)(7aP8V&HG9&\&cQTE2=+QDWMKL.-Z?X:C7NQ7NaTD?+Z&.)Wb3OXV8PBB
_&M=IA(D2\5&CaE@bGA,gKX,G4ZK?E227f>TaHTMLJe_-\_;E5F+/-3\a3YJWM3d
70AHJ8S.2+QKH=OTP,?9/Za5W:(5Y/P11)\X8,dT_FfR[Y=[_G,5AS^7@Kg-6&4R
6]>PVH#ENE#W#&AVE^YA7Se6N3M(3,#H-e,d8JVFJ,H2_(S5R_8^Rf3CeWFWFN=Y
8P:VbBRPY3QeO0<J0GcP=?JdZg0/N8Q^?=EcA/caK_4[Q:->2X;XRS640S[GHTZ-
R0N>I,6M]AdMdIf.TgWI^]MR46N<4^=b?6+]CaX5aSY>AaK2-_UJZ\(<JB\)1LAY
P:&DJT-dX8\=EO5HS&^[1FcXg?G3S;V-;W#-CTQ^0UKZZ1_eUI)7<f5?4K_TEVa4
S._g2@R(G^?@b6)YSB@+4B?D4R;d7T,8-PJgd6.B1ZJ(7Xc(U.0cf@.g;_AID\[=
YW..Cc)&ZMB#L^D_=3JQ=LOeTg7+ef55M_5M-+Te\O74?]_GXJDD5;e<ZR@KPNOb
CWD1VG>MBaVbUU+a-I_3SAa8Kf]943GY>_d9GQK9c2Wg>THN9e1g/RMd,S&>7H+\
OCNPe\[Zd5T-J?G:.\Q<VVBFIG,]]K(78T(K5P\=SI,K-.)62(PV+LJB@Q2#V(E:
L<+&M;74W\-6/N_J-S&COTX[9YC,&A9ZU=B#LWR,bQB,KBeU>^HQ&/^XRa61DM9B
_HL(g#a>I5NA5Zf+.]_MX0/LZ7>5;9X?AFMVgE-J8QSNY1aPRGC)P6[(\P;.Ka&?
?1A8^C..P,E<>^g^\/39eAF?9>?HEBM4@,W@)=4&UYK6+YMD6??0NUW^E7A1EQ3F
>ND<EO92#/,7VV]WLBVf@cNf)-YVBeO,f0-OXJ56WFXAN3f:3XMG,KF0P.a#2cL_
ZV6+FAI\6d7P7RG1B@TTIXS7;CP]_MGU:-F>gb0<9GMK9X#c)GSZ)ga3-W70>K-a
FXfT66I8QIePb-Jb\dAB9gFSEb]22P9,+_6/_+>H<e9eJ6TG#bOeK@/=-FCZg[8D
OK,&EJUM]HS5^dI74eJ)L2.P5W<5X]1++V90/=;8.BUf(FO2]E(ePeX6[[.HCg8;
A.WHDPN@>7=^b0;D^GDg.C51(?YTG>ZDLXW;EXEe<M]K06;=@1&4X\B?^B9F;LNC
U#T5f2/;gH;J3bHH>bFFPSJaPXKf];YA+_66JM,7JGIL/(ON()EEREZJcG^OMaV4
-Z.&3[-=DG_4Q6,(N/]Ac)F=^beH^R5d[FX=4PE65<4;fe9&_:c^6OP>JeL1.-2W
GaI;=,6B\+ScCGC(T^2G;d7D/V,VI7fb3.e&d=)G,g4970?_=1bC^fC5_d/cF)Z[
BK_Aa0ANC0-6:H?MS;#U;GJeC@6,/\.VE60:)R]A4W+\d5?+J+QbI+=I2Vd;RbJV
7BO@#If8gRBPAPY,^E;D39?BS3@Q^DLY6R;1cZ#fR>+gG+JC0c0U_-3D3e^;@67/
O.&<E+8/(A2VH0TWYP@f9gZNETb92_9L5KFS&;49FgMd:Pf4MZ]_8NbR(a6P?ZL\
d)9\&ZJXU#^=^?J,6aMJH.SbC+\IW@bLSZTP+.gb2DFNB(+QSH4XAKI^OAdc,+cN
gBY/VXYOP:GQY]b^LM,[&;#eS_SV@WC5Bbc@6I[8<Y>8T-(><#<X+I5&WM3..KMG
N9/cf7/C.G;U^9ZfZ7ZC^#cGQ#DXM-cH&_?aK]NG;CJgL)-3HbPY_XcX.RPb8.=?
([D.E;F<M7QaOXUD#K_JS8#S++SNFJaJYFa,Eg[O>c<SCAg-P-9?,MIL3<JUSU--
fQ[4W6]bAC,6VRG9gKSF)49&Y0)>T][=IB+VgK:A0HDO-8&;OQQ-#P91-I;:Ya&Y
]7DXC#X-)L39V?fP:FP-PS.a9:KUL(PU#H7aTRf<Q<QT0ba64:g++cdJ<UGg;ODB
7R>Hc/<4B-XdT_:G5&IJ[WX^<\gU-S<M=+b7KDK>)O;XX;e-5bf/#TQQD(?)cWRc
D;0/\ZSeRX+[3dg#>;6e2Ad0P2C8\2EG]>)W6eFd)?)4]===6&g/2Z1^,EaHP\+6
&e\?&ER[cd2M73K_EKJI<GCGELYE^MUO)6>^@8>0@aB_BXGY3?(XT2P5:\T@^RF&
)S3SUE70bb5FGZ&NZZ,FI6<,LNK7,+VSB-0LbJIAd^VZVJ]9N&N^6GJ:2RR5aI9C
5N_f@+a[^/2C\Xc.33=TTKKD]gU+9c<X:d4?e[YRZ04A,C0C).Z?c+c38Xa/J+af
B:6Ud4^10;P8AQG_QYUgX=G]KLc=&80e@P>bGIO374Lb8YJB846_5BSVK1FdTMWJ
_CH;=Pf:.PcR<:6QD\.ZLS>;=(be]:BbO:.:Ca.C0:)bZ[\#7La>G9?;)\+C4G0^
bbR?Vb\?eJJ,>;7P/K>GX2=21e1I(5&?K&=d^LfM._f:VRY1UB[:?O0S(CEKT:#f
40.LNeSXJH22-L:-#N8I=ZFLIF07\KT^)@0UEQfcA]Q@8).P68<9a(<.<=89ISU?
YN]5GfRW\4D[eHHWGG>[fVV8VDO81dUJ_+HQ;:;3C+LOABBH8O9^)G0IG7cc:KW-
RHa+;AH21d)e&LLY25<K<a#1@1geU3]@]MQ<.;7f9]MWSM2#GYO+S?U2;D)2()5X
#b6_d<K[XXJ+ZX1;K=M#deH7G>4.HN+^7G.dOLcbWcENC?/,Pda-Pg3W>5U^?/fR
FLb><fL0(VfO9E#L61LXRDC4RF=cXWR=I+Z,AL95U(a708)55+</+f2KX6;1JLT<
.Z=ATB(Q5<C,TXVI>4;>/PTFK=0W8-<=K<RT1N5&6cZJd<Ja/DP8Q--++Z&IaeLg
abd-[Se(8>7/E4T52>;)(-DL\cPRH99b8UM6Df3I+A59f?3<7AGeb_^,K23gQ[f;
_RWVV_[>-_MFEfQB-KCJUDDQ2>B<(18CO60,RL6N>I/4IcK02b:UX#=1<_SQBP/<
3.\X=@>TG@#/,b?OeI7>d2_OHJcBag1U=WDM0G>GeY3dB.JN8KL9NK?UHCA#1UX5
42Q2f>Q5EO0WHYVg,)OX^891#V>,YP3>[V.:J_7b)CB0G)3RE[Ne\K_(c+U+5+)Q
>MGNTUT(E(V@dIgH/.46N)f.QPYU@)M5>$
`endprotected
  
// -----------------------------------------------------------------------------
function void svt_axi_slave_transaction::pre_randomize ();
`protected
PYN^VR=V=0<.X&:?HE_,=0:T1c1@+=9/c7^_(eF9C?YHTRCVMAE@0)J6A9g-8</>
48KCZ?W=\b10:=VE<=FWM]+gfSAcKTVUJI(Q@5HDL:<=_@>,6ZC_#.K,R&,e^5G/
F2T<KYWN=Ud+c^gTG6-0T+O?4,W11?9._;J24@2A^PZ[a>WJa;fY?64e\DMJ]E)V
]<8)N4f4g+3SLSeAQ^>;RI:FT_[E-WeS4#2bJ5.0&RT[3B9Fg2VWJRR)@K;+4;4(
TUU#PNCHRU.3KA_YIPK-JBHE&01A(@@A=H8\J#4=<.a[3@O(NPd47Zg>H[b7(T=,
PRC>A>9@ZO43)$
`endprotected

endfunction: pre_randomize


  // -----------------------------------------------------------------------------
function void svt_axi_slave_transaction :: post_randomize();
  bit data_only = 1;
`protected
DSfY(a4;WGOK^=H);M_KPJQ[ZdF:f_?\).P[g1ca_Fb+4^9>?UfX(),9U5P/cW2X
fd,7#464^0AC20f514,RJU83?g7gZCPg2GT9Ca?Cc?@+C$
`endprotected

endfunction

//vcs_vip_protect
`protected
3UX2CTMNP3M5FD30a=R+(6N<UC6+e4B.DDOVVK?#0;c>#GC<TF.64(Z26A/[_C=@
KB]#:D78U]05DEZNfAE@;3JQ+:M>>(Da6B\7/=b>4,E/VCQgL3SCS7?])BC^53(Y
1[+VVW:d;0GNd\G_9d6)515+/b@fUT(Z0Qa15]T:S242YUOYNP[^Sb>(6#&L-PgR
eZ701TWG_>\;MR+4]#]N<ea4#5cD+@#0SS=A@N4aY9>edT8fb3@,4-aEC\S5AF><
T?3Z5G5H^g7SVYI)+<569_J4dWWC:FVd#2M<a]CZ]QJ)d#KZY95Y(3Z_FMcdV[:[
d++#)W:X0LE,8^]6G;)AL@&Z^789F#_WS.V3,N-\B_DI36@PNO9YbR=[;5G)dBc/
&^YGO]DEZWTG;#H9BXf>3?MHc]<E)b^c7_ab_?FUO[QNU\@,6VBHaR3AJ4S\?O4G
ee(2&#0[3a9WZ6:RI-;),5cRV&JE&_a4(,G#&2UK&;#Kd[9P(fA.Y/0bBd=6-7GT
A/X+fd.ec8XE+)9f0]TU;3fI7+U=W+\[2.#)&<K8,c\JZD=gcR6G=3^9eKeA&RI/
a=+a12gAVbc:gUaM2Pc#<dE6118&;Je<+UM<1P/eEf@gROeeN_B])Hb>S:?@#;5A
)#,<BJ(b.I2a7,_UJDLE+&EZ13:D[-\A,baga+UO;)^(U^B0@(NXCe12C:^4F[2G
(B(&\_gPK4ZN74d#-HeVSJ:M;FWLe:Qd_?6dT+?T^E&S(>:M_D]](<S@H\FJc8<]
^N^gcBHXcE;M2)8C/=Y[c;C517\F6Pf(S)W,/>OUK8gJ8a\QTc0.7fJLIA4Qc\RW
7JG8(9J/gWeW-M[IcYCF:K]NQ4U;>J:TUZ[:R+Q:g&<E5cb&U8=>-3=]CWA3+BR,
J,&RM1L6GGBL6J]@+eEX,\5a;7KX9D,ECLg@^\)KNX)&<>\Z&0SgXIDd_.IAgLN?
4U63D50B,fD0BC^ZX.9eg.S.)U=Q,HG;#dG:]M=F+cC,c2A0d\9Y,PI=@ag6^#9W
&<9>JcQ?)L6)-X@LTMYL?YX/f-J2\NUW>IW&8@U(+UV;L[+9KP#Lb2-=U&C&I,-_
NZ4L.N+f+O72__/XF<g.]f[f&D=HC-gC3FcR]X4e3GCHM+9@#@GC^>;:16G@2Y)c
&7NEbDJ-CE0=^TZR9>HbDBN0dbcf<5cPG(fBJ85,,FW3\6c8@4/?M?@cC]ZO06RG
K]fS0S[cL4;/Z;,4Ja.dW/g3cW+d>0C7BAWUW-I,Qe]XDH9\[/bT:W,/T.MU7\2T
&MaNbV1Zb4g>dUFU6a[13/G5e/D:_CKK?OXJ_]&IBA_JCJ1fAI<EBdMM#FKG/\0G
UYZ-0UQ\;\3f4YS\F.CU2VF>=P2GHQE[fV,18BTMA0_<H&TUWZ+WNdNS-T<[INeH
=8M3CM;+P^3]24<>O(:,0(H4O\+(DYU/\+2T_2=:BC37B^UG0/_LSSE_V9.R:86N
d<bZbc7c+;J2,:ABC_SQ4VE+Zf3N1#fD&-9.3K=NS3Bc0ZcUI+D;8&Na1g:6W4DF
W]48#I^3X>AT3\[H&g/L-c:G]6>P>^/Rf?K4/+BV</&8(b_-c+I[QD5IM=_-HSQ.
-Rf]aSfQ#?/<ca@YE]U?RgYRODb2M,?&1^RB+MUO70SR?&c;87XGO1:4(XAKIKL^
TLNR6,RFT.:>IfGH)GCCeVAEV\c&18+YWP<AS2;IZ]OY1bHXP4PHN-[ZGTX2Z3K[
+X:bH6811J;;7H/+D+8T#)YB8N(S151/P26JfE#6T:^FX1+4A>N2<]7(TDJI-TfZ
dWE;gHVT1L5.g<OfZUH+DCC,Y]KaAgd6e1\?-0(IAdd,G<<.K3^MVMT\ZC?ZU.K:
,HC[Yb_;^=?ZJPT9)H/a/,3]H6NTVaUW7eN8V<5DZV82UC1B\Z4W@W^GZ\CV#?QC
Q4AZ/YTTK3FZT&[3^?/3+4fU9),#VSRdcW0[XP6Y7,GJO])MJAL+J>H;MK3IZHcf
I9?W_UG]HL/07I@1ec>,V/8,U/.>\X@MCCRG0\_-J?)93@A=-,[UU/ROQ>W@Sc._
5DVA?CNPPI4gb#9U^f>>LS#Gg(5FYa^c0:T#0[H#V3]@TXYLCXDCG_>gbQ>8a#27
UNg_NTeg6fd]74UZN=Q(/#RG>_,7(&W2&f2:]1\1d\Je]4KYAI>aFMZ+DB[94D_)
A--3_[R@CL<F4^ATB:=/YDK?]JWKF\5cC=1f8;6Z8(]1cD>T@RPK)O<>FFefM8&U
KWU_e730=/KH3CGO/A3L&.\C\<&D_.d(A\&.2cgP1@/d&]:B40[a?&8JD0_;^@/C
3KV3Vg/H;+/?+^f\5e9Db]1c;FS(22[KCgZN?=:C)2ecL.f1]0H5-1QIABNb&XZ6
^(gD_[d?)+TT]@Lc<ZTM4TVTWX:^WFa<L/A=WJZ__OfEG7#N3#W5>M(TX:(eUR+S
(^-]R(X1_+6IC8QA5F+H\,XO6PfOZBS4RHNN2Ta3BKeEY76B(HZ=>a8+a2]5FVGJ
6bSSTJT4-PV+2ZgBc(g<EMS+Z0CR-.-^@A;ETF=bVTbeIZDK:_g?Lc?3+Q6bAT>Z
dLMIXOU_WN&<W>9Z]>EIMQ^51B&1,9[(]7Y>O3D,(>G5d44bMg+\C][93L[@6dMC
)?1d@.V0XD#N6&eD#BOGHEg1UBV;6&\ZD,3d5?1(W2Y/&C-UcJ4N7-\N;O3H7Z0U
==R7GO:N0<+/85fcCQ,\V(U@NIF):cOAaWC<HXLe&Ig>GaZ?_<NQ2ABa-E?4<,E0
VEHcH#EAEJ5;->LJ2bGbeG1:?+U3:Xf@-9UIBYU]C=)Na7+?4&1V=RfY1&7CVEF@
YL/Ja\<M)S7O=^3&>]HP<G3JH=NNgALH+1&3^Ag7]OVTd(=,E>/FS.;3&A]GQUF8
-K]gQVIE3eP-8B&a[DP.>M)9/_E,N<<[.N](3L3A2\;0Tb?AP8L>Xe^77Q-8N29I
bJ6LY-fgWGI+PZf9gC(fS0geEJ[gbfFdWE8[CC_:+HObRETFGIU<>W2A/RTV@M(?
Y>^bZ.^A<VZ.gG#\YB:^>.;\=E+(<Q3J=H,)D79.>2>K5g]@bN5MV2CV9_/[-gG(
cS_XaB:N?U=ZZ2c]EI48baS;?7U^bfM&&D.,OPJgF5c.-</Y0N>^O^g2F+I-=.)e
\\CR55Z)f;\>ZS0L<K5d4I?-^H?/b+T7g?J/+[[+U(1,G1&2^_CO7g2G[++<WJ85
NV_MMb7VS_#>EHZ+dBI\Ve;eR2CA++S22c?JEB\Je)Q.^BR<:^;SWd;OH^d6;]8;
MUMA,eU)H+WP5V8@Ig,KP^)c?#5NRPUb7QE:LgABH;;M=U?>ZVOUB(.3fNDZ/G1T
_eWVZgRe?\)^,YdDJ>72XU3RA+<.P5>DP>>MH\2,dP^ZLVBP3&9>70;<JgC<fY-<
4\I2X7[Yf#/2QS^_Q_Q[NDCYQPN5./ETMA#?/P7ReW:6X8[#g&IBcV/;d,)_^0@M
6S?g3&b<\K3&RFcM7cH3_HYO@b_Pc9_B>cR89+3U9HA5/+.2d^6Y_DbAd\LBe[bK
Q4a6<W+^e-fLQd(<f(Re1G:FP6?M?/N@Nf?5F\eHYJVAFZK6N>f60H7QcH-2>D01
VJLZ6M=Q;bU&?XW9B305Rf5-8Pf7\F&4CG;:7\Og\J6H/Nd3KK9,S)FG_);ME,T,
-8Dg[)BR@S8fbO00CX9/aa7:K;@#eXH?US5K&I?K_DX7ALAaZfAa=,WY1O\:54UD
Z28^_>DE_,LTUP_gL@:P[;OA.SE-E;5:3FBEURfadW/7,8\@I2Y3Kg/=;GG8T=T.
QOM:0f#eQI<PLJ5\LT=d.D&8DF1YZ20ZBDUdNI;e#VP=b1G^>#MMZZ?E-#RcB/b?
JMC8_IO)(SXQ?c5QNAObDMa-3YBR[0-)RX0+S^:F_-N@_[Ub..V;/cAXZH)Z8+5G
L?X+3Jf]NM@JM7?RT.0JEC;>,,VcCM=F3P>1bbR.GEAD(P/Q?ENYLD;fcZ?+1W_1
/>FN3U<I_GS09\,[Q9RAO6Sf=-)>b=>U\;?7U9aGJC=g6gIe^;=42,NfER)_LH4L
L:;5-21V+Q1G28Y^-\aLV4\)3^>DPGI7N,\0OB0\[(PX&g3d:5@b^)W>M;G#Ibb5
N<>gS<A62H?:HBAP7eRE5P]g2c0JUM/IeI1N,LX9@?@c\&3Q1=L/_:fM(W[ccZ3>
1ga82284K,ba=8)/;R>/5U@daEKaV8f)ddfN\+Q>BKW[].\0]#cKZ7A2DPN\95S1
?-NA,f<PIFbJH4=8XFDEf+(D8O=(XHSZfE[^fX>D&GAa]IPKSPf+[S<>fXXX2dC(
Z?7H1-H7XGAAaQ3??DJ^]C-6])UV[)I45.9TL3Z5H(JVZ0K-X6bF+&R[=)WSRI;Q
aN=;<c2@3gYgTgF9:eLQ4EMM/GI:85V?24ZTAXI.Fc6R^#(\0IQdAI5L9EQ,4;:-
JYId>@[P,:SYW)8KIdH,F:X6WXb\-gNg+044LAJ>/^ZN[F+A7T^)]9,CW.+0J47#
/L]fNU][7A-,KX@c1JG)5S&W?USD^L_G^H\TbY>Z-RM,4:=6LFQWK91Y9[Q\24UO
d+VSL>8/5_OD@T(;_HN-U#1=ZM02NG[BNHL^<(_W^?5XJ1VNC2-cf_QO[CASLS-/
1OYB3.\\+2WVR59=beATXReA;E<H=:,T[;IP]T+79.BN@A8AE^;eZ7JZf,-1,dUU
E&3g[97KW0&CUOA7QT[NbRT?MBLcab=&:e4e\.UHD-bP8HHb#f;:4T^ENS2ON5He
9,9P8,@A)P[TINOfJEO;N>E&0MQI/MN(ZUKWBX[XJ\Tf8.S^T#A?F6Na0_Ia96Re
T^6R8a=5<6aQM7>f2FF@+(GK2];LAKSaU<P@^Eg>\c:_V4E5)]SgY@F/Y(9P]P^4
bS@VfYE,RbLFA3RSg65S1FU&YN44S&Z^DHY>S#];]@aUYQT^AeN(_7-B2T7WaBdB
c=EI<\/ZDPfB=0Fg\.JA)4@P:?YDgB^=^9a5Q&>6O8g@=:A2cf&KC]Q?\.Z#@4KP
7d]T#<-0)X_d7;UA:EM&/LR;3g;JH+fcNd7+)8+g6.:N9DP+^Ye72D4MQgWeUT(6
>U-S?XUZ0(]Ba<8)bH4-0Ce@&B56/+9RD),2Kg>-e)b@\YJ/@?DZ9MNaN5<QMMBP
bY+JJg6<_5-<^,9a2bL2e_cT[>:6(5_GK.BbXF;5V-S<1;d,QAfO7fG6?7_353S^
S?=YZKg)#EYd,9_bOa<-6DeQR@82G=dCYJ(EOb)<Oe4a84SadPHENU^8W7IG\c<?
AUQg^KBOSUDd1>LONe4a1/a+MDRSYU&,\b]f],.9LLQ.K[-WR;(0:IEa3\#UF@UD
Tc:^,b7FJROCE<D4XHDNZ55I++2=WU@Z7;>K,e4fW+H3^GL>f(SdJ[Qg)C/2C5M#
=O7g)T^&EH[7(<g_A?H._,J?&3E1.M[M>F(M)B87cbc[_ULV4V&MKP:GVM58>H+G
Aa2_AW1_,/>XDB/7#g1(g5AL/6D/^>XVP#N:@(Q0>7V(V90N-(0]9Z#Nc=RI>c:d
67g1&06eNH?gL76UDJ#77<c)3(4gKP45[Qc>=&fbQ(B+Z6f(deHB<1;R(ZP_VER5
TC&B)<&c^7M[CH#f]fEG)ZMb9IWH4TB;Ja8<H0UI_-+aA,e,/1OJN^-XSE8I8MY_
;@VL4I(6LWHeObdK9@0La1>c=L#]@34=S7^I8WVTV&E__/QQOI(?7YQQ,Acd_PS0
C:Y9T?QW5\SL\XT6.ZDC,48bW@H133d5KG9A\I-2_OH>1,b+;2\#.FW&UIR??P#g
YQLd9N/b_KH>XC<,NBV#UO[/f:9OL0CR\CDLIBFF(XN18a#3MPA6b/CH12A5CRQ>
c5c7;F7\;[W7X?(3TMaWH#X++1bTRZTSCV0c5ZX4G..GP[G9=+8J52)MATYM/QYE
2-Xb#I7;>[A75;8TEOMa@B.R_Yf#W3GgaQD5:7/2:J]IXZBC[5>NY3D8.\&+H;[1
gR)?GBUL1b[3^W-,]0<?I#FHCD_fLRc0;XD[.=@EH@^CDHSNb,S5QLY1JD&Y.#@V
0GP59K,(>+87ZSb;+(>44Og^2?9\&H^=9HXbI<(bMP2Y/M7=#J8ZO@#(].NbPX]]
#6Va&eR:C+44@6AH]3,BT[_X^[1R9M_TZ8.ZC3aK^8E=dK<4V>bP,Ig)-9B[5EJU
bLPJ<@;QVXC>E#OSOW9Q<Ug[)QEbY/+4Y+3,5da5)<>RY7O:J;W1:a^SXK6_I_+Z
,F7\[M=,/cKX54UFb7KQcG<:1&GGGEDeJ_>8_GI\DB?SRL]a3RN9=I+,TE)C/_a0
N=OSgJVKX]KZ3NK61Y,>5N=OGc_>cFV3[2[YJM@Uf;_EGX@><6IOGG(JASB1[Uf=
S&&AA[DE(J_J7R_LH+BPA/]]7ff(D1e8^A#^MDG>,^Af46DK5.RU7c\;[C?+<>S2
TRbR1U)>aS.#R#=F<[&)M98Ng5fL)Pf=VVb)H&Y]L4FUHBN6fVM,_1bLgN9Y#9&_
:2b[cHJ+d^NS<EUC--W3H9T?-aIG,_-Y17R>>gRB56[<I\0[&,_3-e@AYZE(6FNH
EPX<e2_JZIJ#:e^aU?=.,[]]77Y-H4MIE-3+Q#JY>:R8J(9(W94SdZB729>MGW[M
c[QME5>O?ROC)S5<ROZ7JLc26URM?X_;5PB4W2C]>eZF?BYc4>>4)ZAD8)9M7W68
.9>PPAP@C93#8SEaN6UATN_d:H//Ud<gNd,c&DD]G?KTOFJ-TDY=I)M]AT2U_acO
<^e6[MC/f/N:,>V)(1V_Z06447RcdJL@X+>WcVaWD<?H_e9.I\0d9/&5,4=b1Qc7
K0_.SVI#-PY]AC;ST)ee&.@@(fbY19(D)Fe<E:(=&KDe7I\,/NfNaJ<P<\_KR^:4
/Jbb7XSf7eFZC57-WL7G56.-?gIF/ZMMO]ZB,e+@HOK63)3PQ7#TW1KebKQ0#Z7d
KZ>a[QV90WB9Dc/;&/<G,QU>&+,Xg(DbLO(0Ea0(-86-g>7QXdIca+>,N=51D,79
A5=8c4JY+a^YI+ZC#8>6U?X(b[gQ\ZTO&LDY.[3BV;^82^IObV^A_b]2W9N&)gU0
160U#a@):IA@5XK(RYO_Y@M:Af3FR.gPHVZ:V^CM20ABJ#P-]QU(Vbe/BKbF)X?d
+@ZFD_9U=,JH/RG_C1Y;5b5<1(0PQ/HNcffU&1L]cQ@#(D0IFDV4(3R9gVC)0.<E
UNF07Z,<_>.NX[FZ^bgIKc^0ZEQU9a[_gJER2?6P^/>7e.d1SYYPHX1O68AJ.A/V
-bFeefIAIM(6\4]MQAeEI?2D;.?VN5)c1e;^520);(aOY^=H7V_W;8B08706,B6;
B(b-5)U]YF7:TEU(7RC3O_;WFU=Yd+Y6Y_^948FI,a+@\5&&b,6@BRU2(YI@5Eg2
c]W>_0@.?;Z>-]E?BNH>9(\SVX_PZcUfMSBbI//@f]EWA)P.?_&eGW5BfWG]T>K,
\-U)1TWIM0d.\J0,^3dK1S=B(dFW)V#/5GLc;#&S27(E,@fHN#)TH;1]d:)4&f/I
548GO8PBW,AEL>NMZY3@7-P73Of8&5&_Q.[N^2ZFg&+U:K2=DbP)U#(3N>MRSXA.
0g01NI-bS;g[[T6H6cCN@2Z1RY],[+\fP&BHOHRfYJ?_5XZ+]85e=C#Q110>:6K?
CaS,PB,dOHK?b-DBRcK@3DOLfR#KSB]E>YM-8PAU4^DSZ#<4cNZKG[IWI3V>d-3.
R8U2=J<?(T=f:>>463A82eBD_gb^dXc#+.Y@EFOZJOC+,87U<[OU;N&T9AP\<AU<
bY),e#:c>JB>242TM)5cP_>07Bf_bf5W>a_D>.N)0;S#E+^Yc^,BN/H,BWQF3OTD
Xg#LLXEI0+FYRE4_d??^KL:P,-:cR_;.[OES^WWabPAH1JcS]CRZ3R3Y9&70e7D<
.\<42BR_MM:_#_I&UL]2H7..IKO<86ZAYgER[Qg+TQN+3BOc?ScE7)./,/(fJQVd
>)#S]2g@e/C+Ng(#D?B[eTW2b9S,dM\,^FY3F:cbYHS?.8>MXbP(OAS1:=EI6P/D
PA6HWDd3QdHG[)GPR2WVNYTV-60fPW_]IN2@Z[;85P?gbH=Ea(S-[8N4.8b@_HA#
=-FM1,YKg0E]ZF4XM:/FV5e-LB()H[J&#KB9FHC8<>?;G(;C;Z8X>BUP&+Z8DDBX
J.U&2Q4]?161=HIC8b-d;g#ZXQ0QdBRR2W]I-UcQeRbd[#Y]VY>/2LI^fJK.?[FX
MbZ3G)I)J=[8F85.TabGa7AaM\?O9[[D&eRD09H.[/?FGL2\^1.&(S[1,[(JPWP1
gC\:fI>EB1P;McA<@HLZFWT:EYZ3;F\0-)L-N\>ZbT>HAc@0Q0+;RPGVI4]HW&f/
3+^4X>7E/R4B\>aRK1D/g89c=K:X=47#,dVZH?BP<)X<c&ZQKRdQ0K^I6L+-[,2c
M-9E2)_D;^Ga9bTaNT7YNNLf^^MKSS?L#.9?JF;QaQW34I/<JPU<W4K#Ng\&TX4e
,H;PK#16BLf?R/5&K,=?T+Ce:W-X/M5T]EMY/>5(PKZVD5DZ#+dGY]U+7T@(4[80
EJPC.LHEP_#76>.:0A-Ub+EYPHT#9b1X.d1ecO6G8V/^TI<?JX0Ib;AHc>QB<f>(
79dHY7,(WU6OAK04?3I8P8-b0I3K9<55VFBRaLGLY>MVJ08=Y<:0><P=F4_&2L\R
T?A&UXe-_g2Q0G[:G(\)_WC:.<e=]/[?f?;N^<2[9,1MA.Uc54G=&;Mc#Xfa_Ub9
-L[HXfO-@MO9MV4])55,PUH7Ye>dNBEK[M71]_.E_Q;9M8L^FV;Jg.,.DNGQ6ZP0
P5DC)K8R0S5(EYLTA4W_dT;68YS\M(CAV/^OTVc,UZGJ\>b@GTWI\M^W0__S@gg&
a2;dP/3+0+=J:]FKPDfI01,;C>aJKOTL6>3]U0dD+(A\2fSb9FP=O0-^&SRdE\JZ
Z(4DeI+gT)OLbe:K5;^?(#[UHc3c<eM,@SO3VW=VGS#PIR;I(W@\&1GJ.;HY0@L;
E0We]D#099]-eW3=/\]\:d.#XIT[2AXOQb/CKJ@g;X8C5;(+;I@+\Db_H+WH591H
\c4)__F;c<\WS@I3/O0U6Z2QgaNYS#@90M:QI??FQ/,J7&4OWF-P5FKEA>#QF4HF
L[Z@Q:eNZHO)M=AK,>fV/^?HGG_P=TW=JZ5FZ=fH/d;Y8;G?H:._a9HF/e@H\KeH
NZ7);XABY#b44JIEPb\+:RdJIARNgV6H8HD:a2FFW+CHg>I,>KA2AQBF5]FCa[?U
U@,U//5a;KL:d)Lb]:2J8XRN)]8U.W:]/A3476REOMcGb@WUY[,;[[10H05A]J0a
5eX+QYJ[[\KJKTZ77<H9f.g8QEb4fQ3ZA<V:f>=a^(?]HK5ZTY?S[V5_EOSRR-&T
Y>P&#A6H6Q+7,_bYE+X)/E02NeTJ1<\)#_eQ@MdW1SKR]5.JE<V,I2X&&^#X#e:Q
?>:S@NVbU0;H>/TVR9g#=/OD>=gN?H&BGF11P7>N.T]#g:^2)_DXf6WG]\GcQU]R
5X&5M&P592^,KKOJZgEI3YC8d:/P]M<:LK\8(83CF63BEI9;W[6,TZ&7>]FSY#<O
@b_7dXPE^_?;QC<C=>3?T&7C36CAY9@&fU=\3F)A11#9R)Q#e\O,=P3;ecK&IZQU
1>EYC0:>:ITc0[]=\3DPPQ_SA[GO\7^,V1PC1O8([7ME<C#Ma_H#HK7<M337M^GP
_8>JM5W)6Nf12Ue7EED@(UC@3-?W-@?##QWUCN:FRH0IUbJT8O>D61POSE8+^2:Q
ZQD)(7YEV]_4Y+DJN45_Xe^/D(@:]LO)QOV4?d)4N2LCIKK/M1de,0GV#g3T-&f[
dH^?Q4K+58<ISVDJfPOA,aX9VeP0<f\TDe@XSX^E7g[f5e?2#);EW5KO&:6)5?,5
5#(aMC+Q,dc(X2H&D2;63TA=N@(+#3M);D7HS;F@S<ZSg.T\:H?0R_4eL>QO1FL7
[LR)KGAd=d[Y)3O&BA?8V(Ag(aSVA^faGL[GCb=Vc.:EL21:@(\H0_S/1Q@&)^<F
)#OUTD@ZPg#)]@3D#=7efQ]R:Cb):K)fEf3a8YGUA&&-M4AIX)ZCJ^],?.68,)9O
,Y6N+5UX;;-^VO,-a[A1]cSbgG<E/AI><U8[>D\;=73/A(#VNPU=<gB1Ca9;g935
e^3bL/S>K<U6KS:?@;O,5;NE/J3?9eLb[)[=<VM/c15F=A5_f18U.9Sa)>,C]e0K
VKb;&G5BI_f\T#cUOI(G&7B7HNH#H+O89G8M.1)8IBb&6?@>g6[M;AcgV15A1UF:
Ddf(1A_@)U?CB6;;5<5e,+fLW.7f@[bQTPUPb+1#:AIX3I6&XRa[/2_F(5V/S5-@
.&C_]J[XNKb?0S4HS4PVe,-HS?,S6RSB;<-)Y&4A(VU11;77T99B82Q5@fI[;e3L
4#9LPG/?gA2gTBa@,d1(a>TH?4^38FNM)]]2LH_\[c\7CN@&2^CCD?RFg5e:U<D+
5@9H;]]fS9YKL)[)2Y23Q-O3bW18V+/M+MKGSDP;VKFQFfEFMZ)c^BVce)Jg)SZ\
LeS^N\UMfa3YP&+2b(]d7[VS<JUMF8I#,MT5Q8O\_0KWR_04+[2JQbf^66MXcA2L
8S@+N//,FdD//K<D?C[;S_XJXN))bE^SY43MbZZdVN=,W7aSAF?&b\MB_LgCR=Q/
_ZV0bd:BSc\BAW09W2--;0KVSK&9+E:.C;SG<e[bf;&</TPV4HM;5PX1+X;#>L2U
#J5I/a7JVCe-a5@^<RLZ7KR:5C=4SXE4<8S^^FU<c<^SI#R\1c1OC0Xb5D:Y8#1Q
_)T->TK)IMQR8\(e@<@]e_ggA?;EXM-<KR26@LbS2+Y]A0+]64D_^P[_H)J5,VGg
6Ia]f=b@Y:>08EW[ST4PF)[bD^Z^W9.1LSIHBY@TW2[Y1fK:H<#?@FK_H9_E+L+O
R-08,[gJ0GIC]LaQ1b_Zd__75DGR&S8b++e@a[T?<GKCF1[5Z/?ZN6URF^CB_V0O
g/8>_eU[cU&3_^\\L;+JM+0/F?=W>(ETZUMD&--Q=_ZTU?<ZDGI0#EgN/[59E&)5
Ufd/[MU=I\[._,cGf/9d7X=g,X:_12ML@72YbFRVLZSTP4c8;L]+c-2F@BAX^-U[
;b#&SgL5:P2eNN\VWNO\b;EdE?H^PJOKf5,MgL+U@B<MeA8K,^DagR()FG5_\48E
N4ae8?@\Bf:J_M[CIFJ@.W=.<R+8\/Se0b-/10YIY+@K^[,L0b)UGHU3(^42J3fD
F/N2#f?1g+1(5,=.AX_#)[6W93C23<7J<a[<N)FK:R#7-7(26?QRZC5MNOFcN\ZJ
)\cI<67L/\43YFKg5]A;-bBf?FI1X8#=G>e&T/_D)4^BK=<-&Bd>KGX,[+Paf4UP
XH-#]-Q8+,I5aQV:0LDW0MM(PN_,RLgaW>ffS3JJ6OEaCUH/^Gf8HY?:[9-66:2b
@DPYKBdVPLZ[X0(/6a5UQ.dTA+C]_Z8Y#8]7&92GW7OZ73K/<=[O9D5MIWG??F;S
4>900&D9IB8>BC8f&NaM#H0:/96)g@RM;UcMR(N]^9/f<>1C90SJKd6YMe1][M6.
0MQ7caAE=P-e(0AHM>\N].V5+Q]Z\XWH&PO&3Y1<53CDW(C9\f[FbZc1SI;<#73(
H>\4V]V(eW=:W<:gO+#,^T7S0YeA)=,VP_J,MbE^?_][EZIJ:g4&<e2572<,@dAK
EB7E.3)>LTSdcg\&L+9gN8<D6T_f1/YTZ:4JL)8S.OQ8b5XXI4T?a@_9?#..1PEF
<Zb&D+P6(HcDT31L&aO:QVC[SS&.+0FU.)\N@d#gK=J=6#@XRdGJe4eC[ge:bL8;
B[/XOT>[+K8PKWZP7^9C;Sf)?]8#9W@\E4\.HO]VSf4W@,#TROI7A/VY:CSK\7]X
6dbF&bJXYe9TVKd=UO79A/;IUTNO[O@PPbYOCVA)8\Geg=G/Pbc/e:fMP,M/Bb[W
+HbcIYd-WO]2)TE3AP>dWY7E\FAI2cU]BX=^0)d3Bf]P3)(;U0@(0]:=,6g3Be].
I:#fI.da[&>E]4,e<_c=.6B=a_fZUVEOaXfH_KOZRDB?YZD]O_YR\]aLH[5HY^.M
>7[8_PAT)72.QWLC;(]9WV-[WLZLf\+5?PMJCJcQB.?L\4I1XDeJ0?F2&@KI_VbI
+&3J3VW6/LK?JJ1cM(;e#JJBebKICFH]Y8)V:g5b(21G5GX.,&]BSH;5TGX]bbLS
d2.C?HJ/Y;>ee&(I5_7E[V#LR(JAG_+-CI5LQ#;-3@D8IN3b10WZeZ1gH32TBJCZ
:8EG(e-;Q#NV+g+/IZ8J8SYUCE_MQDI^BA(#C67aG@ZOe-=6_,DTb<9O.C,+_MPI
(T8bZO?IBd,EV8c(eQD=9Ya,05EDJdAKJHU&>)M2I[@)=&MR^^9E?@/e/?Y#BZ7=
O[NA<^&:)J#\>RL^2b=EFGA-KX?fP(01d3N_G7/5U=3Q:M/-&0db_>GOPZbbK&b:
\0XVMf-e<Oc\XMaO4ac2R2>fDWKSTYN,-DB>gfcMIYVV9F[QNe_FS<=<\&)YaC7\
1JMU>,I]J#O[T=S\f>:fP)]f>E+968T]3d4f0L)JQCQ/0^>Zf9KKU#=&T6XV?@Q;
-VZcRI@^a/0b;VB.-IaA502J6+#8)_2H?Le;F/0F/WaE9X?VK[a]DaeCJ)e0N\f,
].=Le]@f?c^IbG4X.aU(HXST3R\g7Te,+I+I,U9a[=e,(0)Oc6VP(&1A]eJSG.IL
/LYN2cc74&&84_@4:)TV>+JGaG)PS._N\AACZ_I(P=HN>A^BdP35b@)9NI#bE#I_
=1;II&3L^9\](@dUR/.ICG>0R2A6C#^(A/T+\&FVC#S#NF0RM6cANPJMgd\QLHZV
D&4-cf0+=[dc;Z;b?T?#>WbaHC:1DO/77R3>Ia1P1[M6@X;+]>Qd)R8\?/[LKI^>
)8S/9S]aHQ3f9CP&=/be,:e&QUXD[a2TB6G7E(AIa2V.E<cP,PaI4^R^A#H6MWcI
QT5TcE51a&HO#VU1GT^UJAQ7T<fF4g53NeVQ)Z>S^OO9V;S(F]-H&Qg^UU5,.[K=
:^ATZ1gXPYaA1?EDRaK5.=\IZ2<DP-QKZ>B]NXQfLG=]/;K(C=-G(BJc:-cF]M+Q
O#f4VHA<W7@YO6(7[[.D;,b0-;)(YbQPX/aBOP#PP@f6]d&Z4RW(/<O7^RA097:d
4UP,gJL]CM6gXJfF:W\A^&29D/5USVBeDT9AI?W,_TGE.P>BNP6F9K>IAPNBd5_(
U/3HMFG3R0##-E+]/T=f.C@0.bL02RQF<]VD;DX5CDDH/Fa@@6E:H6OFD,54=Y^R
/&PfZ5?g@L?G9BVS>NE>S5B:Z_c6A4A7MV_Db<MYQ.X9DD>0fe3\U0O^:W=>2ZB)
K4QKA6c#[RYaGfZ/=b-d=YSPA4P>DfO?(X@U,9AI>.NbG;@KX__X[]ca8J;STU0_
ggGX=<[Db&^9Z623cMbOb:4Y#??^,?F(1g+&D1<&OVDAAVUJ6_MbVa-Sef88c8U_
^\LJa==6d)?eb1aB,<YZ9g&)^D=BTdTQ8PF9f=f;Pb(_12\,UH-8W3PcMC\TD-52
0VcZX<6;<c-61/c+3?\@MaSd\+HGCJgXRTE32YTL1.YX>J>HB8D4)&6#PP)D#De7
dc\G?CC_+,836dB1g[]cZ;F\Y\^X>e2<f)3E[TB,<RRRW2]I-GDI@UR?,2?E7V-6
aPg0M+eLL,_42J:W9-<b/M;G.TS](2]7D\Z=3?Lb_W.CM?I+JQ<d12HGU?MMJ?6a
8T?F:Hb[a7+;?Q<>/g:dQEOQg]d5<JL8<T2@-FJ;_P_bI5a>OdUHZ3#3R,bBbKJC
^e@G#VY&WC_\aE8IYAPdBb>D].MbHVOUP;7OG>3;P#g43=BK6->476[ZJ(R.OFZV
(A2KF81a,762+NSJ;/[3<Q2RQ[X+KMB4K&@9=.?YIJ>G/:58f0J_,Q=2Y.>\f6<E
XO?O.W^:2db_Y9g]CLJgVAT0:\=96g>AV[\XZTW0a@2FNEU#_@[A#6(@@_JYU5_,
?26Q#/>&bSP4CJB\V?,@K5I6PB#VK#Rb)(Y>.T<F3].eIHBN5:0^.]ca:geA]c1&
CP#OA45ND2EXY=Sa07)6Z_f\CARW3a0bbU=525:S1=:<EJfX2]gV+:AKX]a[_L(8
4II)(Y5C[NVHY_@B1A,BW^G]P]M2Z;EG\F&^<D,8d.CBP,QTAUO[D\fQWD4YFePO
9(Q\b)ScgdR,AMQ=MfT<B.R:A8;dAZ\HZPU/fFR\7;Y-E6/.UdF:]c<#F@729QS+
)U@S/JaIFSg9g3\Da(SUNGDf+(?BX8eD4&,AB7_.W#_\8C&)E+GD1]\0/#PgC\;J
E;SE?<D>P^SD2eO3K[P+<MQ)f./Bc6O?L)J:aXPY_O&KRLcd1A1Z2daP>#EJ96G.
L7Ce\=aPS6,FTXZV4B+;^&f47e@@[+Vg;V^9eL3S2c<UG.FNXC)YNZAO];(IT27-
&da,I<Z_:Sab7B]DfB1?I&.5GbV-X5@=B.BY0W90@bPI4B4BCL5FEU@6B.gXaF8B
J.KA:E3E&C[TQLg[H/^bQBW,OO;]Lf9RF8.V+8[1UY6,#.BUdc^4]FfaN+Se?3N)
VN2T#fX3SMU3)3WH?(M+8UH>>W@g:>NO_+3aQ\,/.DXV+PX;Y6Tg<U_[5<H6cLe=
cbeS7]SR8^H5(RaS?Fed#d?dT\L0?Q.Z72@(:QIQ\F7^-G3L]2H=MDSV-FWZIE[E
eZ?-+-^[Gf#RD2EAI9QYEcF&P?S3X,R?/?#F<\VQ=GPf.)_c;#AQ6F4E.LRB[Pb0
DQWW,g4=1fQ=U,H1JAB1?&.[<?CDV=]@.gGXFGND+#@N:?:W7dX6\(X@5ECe:Mc]
HI9X&Y.S3^V:13f19<S5dE+UNb3<&N(27,BG#D[ePG+PZ01>Z_a,_\>eGKRVW.3?
2G1QBW:WY0VQMA]AA.?&H?;N&cP,&;74O[^Ma,YWM=&1Mad5RB=K(8fW@(7[57X3
CRfc7V10<G1TI8>8HCF2I,.<+5-HF;_W3IE--U)\cL>B@E]2#d)+CTdCOd@V,RU7
ZM\bA106BcgA]6?[8NX&bL33=D.g:a9cCO\FFOZ?G->&TYDWdS.b78F4&4IIE3;Z
5S#_=4cR/b,Ye=)aXVa<YW)7)=3=.M02C(.N2KeM88bc+\Nc2?/Q_^5RWMFc+[DO
,-H3[W+?b8IaN[PW/[L]N/@C)Y,\-),.,g(OJc[(F21]<Y)(Y61-;SG:cd\F:9>-
QCP1Y\0Q_Sa[Pb&&),g-HL^_Y:IA^[T8=_&W7\fU&R0SO/(>3X_B+<)>384LR&9Q
Q\-8V+K]/55(<5c&G0)-B?(I3;&/[BU;ec>)c.?eDTK9&]6@PU@ZMT..7fYAH?/P
@=&OS;Q[;S7cbM=];U4(CD.2C+71f-G<7>MS&Sa]0KbHE6DX)V,a+_#S[b8L_//V
HEQAS3>g?.]Q=fI))RFF@,dcAaOJDb(^U)g7eK6].C9+W_TgaCcA@Sf6gf-<[&,.
e^:JH:fA6G>a)Bf//((?ZbW#fXA\;e3,97[fBcPWFHX&^1WdBHIB+H6YaE?HB1EX
U^LYg9<VKO&->Qg4fR4#=BIV/^\;c+:B\(([I?g7&1-ZD.eIIN,W#LYJSC44;#f8
0G\f+[eS@^?MPP-SgN3-d[FA:ZUM[HZ<F31Z@:#[dUDPS):AZ9/[Oc?GRe;_PCJ3
V5NRXHA??OPHF]@JQLOI/-S5e9_Xd7@R9(8g,),CM97F(12H4REN]F.V0=]Y8#3@
&=B6^-80>]W0IAE\^.)-bIYB=L<NEJ;M@_CEZ#^:gZ9a2,0@d5^.(:&A>[77M5R4
);<YWg,4e;[O>CeYgb:;,SCN=(5I&9<?GURT&d05c5,KSb<]P3GR_=&M/L;Z52)@
(@VMHO36YSH,,_UP;U>YVa2\#PA.8HMA6SJ+d15P9]<8GK8-U=LU^JQG=cd5RQG/
YaXf5>0RGJ[ga^@:\#7G^g82a.9BL1#8IOdaMK-YaFF:K^AgE?UAbDa:fg6C>ga4
?Ze3>]B\F=.7f.(:49HCCc0&II0CLL7AVC409Mb.0Y6WBa]bS-L)0H7?UFa0P7;7
c/<)dV^?d&B;/15GaWVCR-#38a/N\NDRE5YcJfET=>^IScKP91);&;(3)]QMV:LP
WPfF]<]FQSf5dCGY<_E];/SQ&,@1IScJ6(@0JU\I&AG_#9MVL.1.)=E-e?g@)/DR
)BN;.?)\LMO_D,^1a,@0VGUDOHSOOQDPIR7^f;[\G]4c)=5@Qg[B7T):T<46X+@Q
S>&VL=M^2-E#7Yg]g\a3]HVRge;BXEd&>.RGH1:Y,=;-<\Z=EO0H2<cK]R-M.=eA
Se;\AGKEU)VT0g&<1SM9>^+C#0:RLWcGHO8X&e>T/K>1bEAJ?Oaa#CMCZBZ<FF]&
C(EeaR,-Y63<5A/Y>=QIZPNbee0cgK7U_MX#XGFe-3f35Zeg&>g6A,/Q1R2AWUcF
7-;N/9d_e0G2\XY&ad<A6#H5g9Q[=3_d.TaUEV?VJb:-&6/LT>CSUV#^g)Z>K87#
5YQ/F94c/:RR<H&R314Ab9FNE(d0PWE,e8T@ZGYOXZX2JD@[HC5cP&8G+BD;RPN?
R;fNG[X_]_(R4SZP9X4+[-GSJ-(/0=LFX[X@f.b:X&MFRQCa^2?Mce,-NE8BV0\2
f[4Dae2930#.Gc8MDbE>UJ<?)_0?,c^P0/:4^/4I46L_?eE1T[^@;37ObO7S?cHU
:.dE+<U:9_Y\c8LG:]=gJ<SHMT(Nbc]3VWbP],HJX)\6^3-5F79XTA.9NOOQ1@f4
)@[B56#3SX,S2IH1DJIE_gOZLGMJ/&C?OG2FJ@_F[7H)C@HE9/,Z@[;8(JPEd=XQ
b1eM]5Ua+e(.D_+.PTPEST<gD_A1?=M11=a8NOAQQFNR-_F;0_Z?bV@EdHGE?_GB
5C9[^_-;[Q_H;O0YEfXU.DH0ZTL5WH+gJ2ge239/+DQ6;L\9UL;\/CGL/VOCOA3<
X-B8YH;<9K60L-A#&aR;bTY8bg\&8\&Ue2=>_J2CcR+GB<K]e-C4Oc55C86c_:+,
DD.BZ_R6E2V[NM=AQ#:?9]+\EGH#eKbP;)-5dB09;.@S&e:K/c_;\#P3-:;<=J=-
eM0F&WMF9,(<c&:LITJBb_Vc=E^AKJ8bJC5\N(7f+TNU,\<XVT=2K+O;[+JKcTBa
BSFI6BYC[WHTG#6QJ[/])\F>PN&]fD7R^8)S:T/LBD8ATRAOENHa,/NHaaAW[KG4
(0bJEIWM<RP,V9+PF=HQS\L0TEF^\SDXaf\HJ(1^d(N^X/U0S6\cGGUY0:N^=gAM
R/G)M59^XF-#JP1S;(B6?]dIf\5@5aB(5QMgXS9V(Y4+K+U]c1T3UA1XZXYGZLb&
?MDU5U@3Z8->Y3Of+ZK6_W+[YTVNF?@/&>XE6F;M7D7FWO+Z?:@88:cSDF7(Q8==
29#YZb@3BgLT:F<F;Q1eFA0HGc)<;5WEXZ?MJ#XDLaf1F93]0:+=fP@Xc#(4F5RO
9HbgCAc^fgg.9(:G]ccgLbf1QYH(1&VTF\&PVRWS(O-d/I+Pf:gR?JaY&=MFUY/C
g1T;3CVbUe13D]>UI+H0R(0f;>&R(PW_;bD8?DDM?2DO9NU@+4PcfC(\/I:)g:4c
Ya7S+0LUU^[;2H>><a,Ug=C,:,BSKJ(+&2cJ-R?Va9<)R]L1&8bM;5_U?/<\05IE
ZSO_KeH0-WU67=HD1QF#D<+MREa]FFcMQ^f+c0;W/AM:&]8?f7VgD2g6WK;A[1g?
^<]5HFZ2T^4,1f=XJA_?N<63GLK9:]5OESVJD,#R.=#_c2=EX9-fb_N4(/?Nb5IF
1>-9DbA#A5Y4AaWgB>AR#&?Z?.Y+?A1>g5TN/)L90K1O@RbD#,&)91dc=LKYG&0H
6;[T6SJ5FSF2Z,?L<F7b\E+BSTER8D?B&,.>)R;S@df2Q0KKc+P)fZ8^RAW+)6V/
AcRMQJ9EcTd1e4FLc+aMTA@.J?cdN27KAb479Y7?C?;@W[+cAC[NJDf>9]YEUYf?
Y41J.=-5f9)^0;M&ZRE]g>PA;9E<M+0=gUM(-WM[0)M18@0C#WE&MA(S8aQ\B)BD
acL^?=94EJXIO?A0bOd\D_;c6[SgIW^;b0cO8H/DKZ@W-N6R.^AX=:fb#S2&dX\5
[;aKF#\(\?MPf[a3E?HMbYC2.Zb;-G(WKZSJ4KeSPMRL/EQ2&:5N-FN4,L/6;0[G
U_:)442A4F4,JWd@)9R?Ibf@1@.S73MS_(.6gONC,?UT]c?a]GO;aZR<A7&).,_+
MI2CCXgV2?&>dA@dI6?OEIJ-+.SW[1^e:5fd((D49O&NKD@9dA&6WC+?;?G)I3X4
02Mc\G1L.JTN@RD:9f>X;))_7fC,O+2](ICT^GT>+Dde=ORTHD12N3GW@O14UDNA
JaXT)&VQX_8LC5@?d(_d+8)+g[^T>Q<0Y5/(A:bdA(=bQ+Y)DI@CIPfH_RO>303G
SLMZ]C]]LMA\H8G;]3^E6JS7@dY[<cR>e3:PY[Tg/PPYAO@gB4X>L\?^g\FIFUG3
SZQDAQ;JM4CZ,c_/-92[\\Yg5Kb(^Z77)K^XLHU?D3X+ISV56TQ7>Wg^P/8XFQ:B
FHS]2Pg1E-MVABb\E]O;9T<)A5:C[@1Da@b=YP3cE:-.afb3N80VRaI&,JEW1_gW
cI-I?S,1,9W6R:SL&GI]-6a#/6/>2AJF4?R@R-26HMHX)_?V[^TTc_Y78MC30:8]
c9C2&?J7901aW#e2R^03/S86QYg(8b?TZ(7AAHWeGMX?B<^+^E>YY37+,4.#A-cT
<U#\V64EET,(8H_L:W9VW,WHL6.TX8&;8FT@dEFH2OPg&2gEc&TJ]L9)4LFGa1=Z
;-HE_A^J5@[X^(JQG(9G1]LWK8=e.6g^TaUA;KULLW=,+cES_FUIBUaD/e>^HHDg
g-3acbQ<VS4bUQJ?P[P>C[d)C//TSB^XJ&g_88<9,LHALHOXZbJQ?@&1IG5f)8>Y
O]bD:B5@)()D8GKJc.YbYJ4??;1#(AAd.F<C1R(4NUX#U?L42)=<3IT\OWb4&9OO
W=#,6M/<SQ\S@S900KgEPBR:IDTgW]?;6QVD-7YF\F57gI^1TgHSX:E&./6?\>,B
.(19Ra<Q5L2BIbSIRT5/K[&NN621(6R+E/-6R9DB@+LCcBMM134@;[PPdbU]P)]3
33#PX]ETT/];LYNRbFLd_5)96KaE+aP>EDJ2Y/NI;L6A>#TEFNP@#DOD@OU[VUU@
HV9NX5&@?A@U]/8TO@,[3/_RE53NMX\E;cNdXHB\\=DNKdB44FaK^@T]N0_+N_VT
R,\M-e]&9H>c,DeM]Z5EE#adU69M8TTZCY5ICI#1<8](6\^NT.9C5OHP8+LLZ?\]
Q4^X6H&13Fa03^Vb30H90+<6Ncg5-&=,DFC(4\MeBANDcYTYE2,cUFfZgQVQ>IIQ
5=ZdQ(.)(TZ_V^d0PAR6NF#Q:Cd0?[MR+4ID/<&1FTKHDBG-,#b(E.Z-1<-4@eYP
I0=@2#8U7(f6@Vf_VT&\:.U(efO+ZAXf#R&T7BMXKEU39NUbCNVAgI6YHG5dXX7Z
HTTXeD+F?YY,+W#+f8J?OU^6X#T-;JI5:;&;0AWPfUg,,fV^9;5eXO=ID03_[,#E
XTZ\SG,f,C/1abFWF4N4OG1IO?Ug]GLc98-I(ZB>-1\(I5#dF6g<)4TW23IID984
F&0>-fe3VA5;1=<\GZc#L&2WXU+b)\&N>RcED0aK@4_<dc<9OcR28_cY:GDL<79D
WNPXG)+IP]<7g/=[5QE_ZdVP)R>P^,9:fR0AS+4AFSPIK^>a#Y\J^+a&&NaOcB9J
..c\_4JS^0&Y\F#M:PeJ#E=&WEaEEKC2P=+KHEAe-B3,cJeg]:#C,++KX-gA5R9Y
J2@?g-\W)1N^LcXW7]\>(DeZIA]I:.<.\@IC#^aK79\a+\,N=GV?gIdb/3GDOYF=
^g8(cT=d9EdN62GF&KcfCD>/6R4?]-Y0]F\bU/URd2P18]9A,T<9LC&fO+Y1ggfI
=IPZ/e7;/8K6:7I\W)+AJeP=@DZ0_/@4OKD@;^EE>MCO#cY6U9MM4:b^.0Fd_9L6
:Q.gZBOS)H+g/Y5G4OF_T1C9-PR2&Q@P.,6]K8VQZD--B+d]Z;:]PIZ8W-g26IcD
JUJ[9OM;NXA[FG(c&V]9\G9\?4Z^<:UJ0T/7R]T>^eQOS5JMeCIa]_/N/IQR-?Y8
+#0<HLdKWQBc:g#+5H)3_c9>M<3Yb+,_+=CPE_b\:+EA2U5HCVB4:X\JR6V_)1E&
J=M)2>HeWb_BSH[0fNM1C\3<MD6CBX51-&4QL]A.g(WE5:@Ra3L\+@BQPUF?;#^O
^EJ5+3[YVNd]\T7_aA-^1\9D6M5Q.H?5X4+<Z&?WZESY>U:K2\Ke/;<Y@e:7eR,P
0UM10cEW^1,:3DNRNTTYQ)-a7NDN-0M2XA=b5QUMBY;0.&6@d3R1KB._A>P]7d=4
()=fIDa2AW7bg.&/AG64>_HTNJU:Q;0Z+/a-<O>>A3<e6a0<I-D?KIR0/CB88,:J
J+fP,+]:B+@<KbT0cE_\J]>>d@F92E007U-gPEV<=[35G.J9E8N[MK+H:ILWA]V(
E,(a)R-CL.\Y-@K7gHSBd=57NL/0J>J@/_L9TB8e@U5g0PfG6a,C0e:E\_]BQ+#8
+8[J394_Ig\N<JTYdG(CbKA(C:YQ>N6HJ4<Ke.;GVb_d(=4N5=Y@QA0TVT;8#8V5
==F=&O#@VV/+(T8:TPRJ,K4)F25>=dgA0<B@7NcXI1YVH;+YffJ?HbH)67XeDd(N
,[VIC7UZbS(]Se0WAKX0)[<PI5VKUH7=1.gBABWZF+55S[);1<XBEZXZYc&0C\C0
a58G/HH44QVg[ZeCQ)8&_d2D(8>(S<)X?T[UaFOJ-V.P]&+O9JfZVg@;g+UW&.-?
:T5eT+3&Hf/GS<V&dUJ-^JD:YL/U2<FZ=V1f+b(,X5J6M[LLOBQAW5WO:\W@R,,]
QgHJO<X;e\?-B+FH#@+]KfgZbdIE.;QI:&U,6W;O5bA[2&7T)B)?8ZQNI5H88-CL
/0D>6ZgQ5+@AddEW2@R:?(SL:VVBd:]^<Z;3^0bJ<-3KI.Ia/McN&1eB[4F05g54
-TGI2,)\O;+c/<-_S4M)Z.5dZ>SL(]J_BRU4,fcKJ]A1F3@&\C?Q[9eB\R#IH#QX
^U_Y_URDe[d8;/[g37b0R@\fBP=C1?=Y\6N^]2DFYOXN\9W.@-XSX<[=PUMY>@LX
A=+1b9CL+eLMaVE4MVJaGE#N>GTKa170A#F>/Z2BYA<GW3X@Ic\?ETO)G@Z8Z<6)
@J,7&G3;(^C+>,1K\ORKC<1YUM]A+]Qf1IZIR=-I:?MPJS6CCMQN<NT\[HW1Td:T
bJNfg6P#=_4@QdM;K9_:^ZO;):08@1LOO4Wd?:B(]R,M)=\:(G?-\(5_=I71=X\Y
]I\A^4U\A0Y.,Z1(DV6A[f1X+PK[#96ABIM^,X\E:HBObFPa30X1;bd^Nb,KK4H)
O:[;H,N.IF>)EUCZKM&L/TF0H@,),CV?Q#V),U74XP-K^4\_A#K<^7O(/;;=.fHT
V)g02&)V?+JG7^,dFJC:CO?Z#Y?KY9E-:@aB9_6(@DN=dQ&F&DNO3/D5PH5+<T0d
J1JQdF/Cg2d(3.8Q6@JPaRXc_SEJ-A>.(8)^WKCGV=?&)\BI;PDI@YHA,#[Q:A6B
OcLF>AObNfgWHe@50g_USSW6^U>MeaTB[&]EcE3&</WI]RZf-E_7=8WQ&R>+#>9A
M[>-5WF:JVeZW49C^]fcJT46(N^68S6^R4f.:W>ONgS>O@4W(-=-,@22cOC+.2]K
.ZPU+)^C=IT,(MIF=@T&EY;OM\CNa==8PSH#1G)D<?7&90.01OZCGGCa468/J-^?
6C\0YDS:#T>CBEf?=FO?_OK8[\LD9OT&-?fX:WZ1[)>X-,fWS.OTN74cY(YR0A@7
0P6<fSL20>^KX#5)F;b/:\</bXR5SZT4C<\Z2gfJgbG4,ZaE_GaLQ>#S:F],>X@&
083N)>8=^ON?a&9/)<,cd.4f:O:JWb0IC0dGd[>D@,R-IfEN4[b\37^HQ7D;K]I>
B>gHAG&K&U1eD>d_5gWU?VHB93YbZKHQ.ENG8P_PYJ\Te\+RYCD/[<OU^(G7-8I@
&DYV)aGc\-VH_a)#Z1fH>@+2Sg.cTWf;Z16(D=U/^36X>@1P:J]WFMC,fe7&EH#6
5Uf@+TN38e+LO@VQAVXYY=TPMFHC:U>,R7.(6K-)Fg8WT<L9M-ddWW:Y]=]VJ+-I
/75^_^L0BV#e5[LAPPY2:9_X\KAOPF;06SBEPeD1(gBdb\bUddWS<YZZOPe&R)L/
\=.IEe)abH^ZO<?JFHE7A+05:Nd1LXdG<=0g=-+\,ZH@-CI/4MSJ2G3M5UCNBZ,H
442HP?ee,5+K8dFDOA>&G7GE<_+;P-fV=X107-]Z&f4#K0DNdLBP)bCHe)(Y#MSU
+N<]+1T7GTK^D4B5+490P8B@=WSAQ]NKcG#+0(;4^Q?[8N&5L;E/_V?NF&O<QgM>
5,1C7e[U_.@[6d@Z@0X7TD]A1O5?=dD3/(OTTRLH,:dCXXXNaJ2U9@2R7TL55g-C
1X/KUE,>[77([/Z566=8U9.YZfHMSQM8&1^X?X_D7gF-AX4T,L&Pc9f9<<c\VOdE
Kd3-\1;/(=X6T]T]]SBWX)1^F2=\(cV7P.>X^KYTD&VT-I_+>Q]fgFRRV<IQ#Ld,
5<C&;_>?A+)KICgF?UOGaDZ=8Y<\:@;L^6^+Z\d=#bHMYF7-d;.W:a74Y3#[4a4P
C[4.6GVZL2>]T_=b1#9PAJ+PJf.^3.-V#8VOc#U0\ZLAa#LK&+1EF?GbY&X]I0gT
J-EReS51T/I/DP728>ZFU4^a79+UO3=+\Ae,);KKEH15:daJ;E^1D8>?S9:ZNZDg
D196PRUD32]f#\2TQPVGL_f>Xa/_5N+55+08CEC61BPK8Z2e,>Kg&aNg51W\@1?4
DPA(^/XagRc4dR3:1=MGVBW2IO-affG@QdQAZb9Z9L+5MP#dJ+QIHIT<VV05g&5S
7O9@9LNK_=BaWS-U6BE\R2;UYB?0B6N.UU0:;LW0\Qg_bVCL)+C:=^,a9WK17.@N
J#6W.W]\QCT_cgIc)&#3^0EaW?[\F#(259(WF0B?YF^Z./b9=<,QMc=P=YLZ^)UT
H8#KCY>_\L=D<=Z2<EJ[)SbHL+D;U?R)FI.(WZ__[]6+WD2[PFa[Q.=c9@?g436.
PWVD1S_fU+ObPHFS>A,_3;<H7b\+)JERcF4V17K)aY&[D)c/fP,Z)>]T-&:\fL0.
GGUT-+,?D^2KJLBJXY99,)=f/OgPX\.(3Vef_;)ORB^K6:):#::)E)?)>YB]d\-8
PCDa-fZ[AJ.&gVZ4[E4/^S@(Y36I\3_6W-S7DA][6-]ccEY.99a#A7V@EVG@:\]-
RPCPI#P2[P^K8@TI(G#>L#;)]E,^(6QO]/0[X&>=]S8:/Ma-XP6^8gZ77f#XCZ=^
G9@Lf;DMObN4YB3_E+8]1#bW=IAQ?M47ad1?T>HN9_]IHSWHPeR)<3_I-\32@?-Z
2R,,ED9+=18<])E-.;)@.e5-L,)GCKY\,SdTc^VCESABd]@;D>,2_X_7OYJMW8+S
Z21dT/4L+f\C7E&V/[^-V8Yg+FLb>,_SG^+^]S@DOMIKZa3=1VN0&P2_[U(L?:bM
@I<JA#[E\\MW]Q)1W>_;#.SIK&)MLcJedKG<)1QZc8Add(^<NbNLM?<U7&:Y^2?^
F5I\EFYIUgI&2OAY7=E6H[5H^9I46d,G8DPKNRL0S@TgVI@S^6JfVK8eL275>2TE
58b9^3@CJR]Mb;15SZS^EW#SY[]dYMYD.6DZZF?PN]VgI@#Ib#,^C.&bK;3,,86,
I59B&717c<a[N\).((]K5:D7U>Db)(LPB8:?7#<V+@YUQ7:HF(V)@J4\NSU4W@-d
W7(JZO;RVJ-fdFHAa;:5A,.-bPQO5b,S\-7YOCfR4=/E5+;/5(F?<Z_2KI7D,[^A
1&QOI.&(.]V.8+,6E@Mg435GI(-:IfY?U_[L9cBdWI-/[2b+?1&ee7;L/-[d46bY
GF^9@JYD/:/S+V:KO-WT?MafPRDC,F(.B^2J2&N#VcVT<,?M<,:;J,^V]-;dJ2_C
O;CHA=IdU(.@N]:W]LVTS]e)XAEW.?0W-X[C3aZ6PBe@N^d.g0Y7PX3G,>cdGF)N
cc??SJ+BFc@5<Pef\G8A/OZ.#PC)f4;Jd&1-ON5g\VU3R);WG:E:.QgA#g_^cL)T
66E?NgF#[#Z?51bW4\gW7>7gNZ8HIJ((&W1ebbA6gLP&.-#HR[fV^ZJ)Q-LQH3PC
0A]I#d9=3QYBaa6QX+K4I1(#Oe/AZ1@MgQ:]+Y#4:X&?\Q)SKEc9M3e?XZNL_8\D
g0B+W0\H@.CfIAa)TKTS^gK,YEI+LeFfTN[_9-IO(@OS[b;8(E\)YLG((J0NH6cg
5),H2d8-AFCK3XXGC:@WDXPBOEF5]ZNd)UM^F)J\.5[;+>OMZ]#;6bYV4;<(fDKZ
^>4;MPMN>#gf/+<.8)PWa#W53<7D+d_?)E,87/K/53CLD=&,W6_P2H)U/fa.(88\
@:]&Q5(.V)#8b5[d(0U^Kd8<1SJ7Z;cebXH>&9+0dVM-b7e]4>K#[PF3fV2Ne)FQ
0c7,:R[8&^HS&?X3(;MJg5/5][I6B1].J@#b-HIQd_KW>FGV&.I)&M53,5fc.>K0
_/A0N\b_)Y1dW;d]/P+_Ad9VMNL+=>bL=?)J0Q^WO32&ebINLAS_4Y(7[6?U@2^B
cFEYQC]d^15=NfJeV=1V/bA&?gU<JDBec?BTSZN7AG/+PIN];DQ:9Rf;?FLHE;J[
f;Ub#U>WSdcIMDbH1Z1&U]aW.+06a^VM=ASC@R(MaOGX>6I:(@d8.:d<NZcV+3c@
JOCebSL>FM1,<aI/A=SJ_2b7efSdY4DY,Y&L^K,a3,#1A>02^T89TdK.8cUR]@A4
[<]AP1bNG?WFW>K06N8_]+_Z,dHM;eOSI927@?]+5_5AEK.=Q/a?;7>R>.5QOR+&
7CL.G6JE[XI=9=42^8&g<?7V?8V+/<Z51ZQd/2bVMT#AfD1aG?3<LHeb?b:6JCE-
JP[T]_)F^@>a4eVIE3<_bQEC6HH=FFR\1<(P;6WagEUZ/C[[N6C]WI9U#KYU.^[?
4I>b84;a52#F:B8,/D@c29S?6)RH#M4&=@a5cfC=DXT]=1<1QcT,4<OCd9AJ+2N>
PR;,dR92EA-BgdLR+>_595;Q^Od[2Lb(\;J#=XP0YW^5.eT)ZUU]fI32+CSP=Z.]
,6,UYb4:3\N.MBZEHA4EB6[4MZMfWXaLEW<.S3AZ0__L-=_-ADWfVSFB)?6:1JL(
5@\IM<>fWG#<)b/cJQEK+0EE1eZ@4>\]>/,W+d7R)1HRDAV].9H<#([??PM_b?95
Ae_@+GcD0AA.2S/CUC^O;aV083Z?d?G)::NXQC2A.^H>YOQ-1E6CCdEZPK_JWD\Q
TV)TVTX+<LIa:VEK.4KTPIe<,C5=,5(AH>8SC>&9EJ-,+<&W0\<eT&8NRFNC_,de
#79=FDJgUP+&@]B+,FE]Mda9d=dZcOO.^0_aQ@Y#923U<F2Yc^CCBB;gU)AYa];<
17H;<=CZT]H8daHV1D#DA9d9EJSHRfb_TDX+-@,J_35N_VKaD9?HU9UO,D,]FEcG
<AD_.4._dB-e[;6ZPWS&7YQ>+O@RC2DT_EY2;1A^<?P+[;Q+2E9>QU&LI>1VE+Gc
62\JNVR\UHeHQ60+=STTJ8(?2OD8\PFB-<9&RNE,WT_5X?3:;P1O2K5927&]5@)6
30V8/:7?GgT=3S.W#UPd9#UFe8I]=:POQ4N5;1QAbH4BYPWTM==#fIUBRCVQSVXF
M#Y67ggUO?;c:BI,MLgTg64(#ac3ME@cR>cGY8g6Y5Bfc/=OZcb+1^YK6Q+AEDKf
g^>&>-B(HVUfB.]=-)1,)1gQ2@f<NY=>O49a3f;K)9EO2<#L3;a6]>UR8Q@TEYU#
_L^ZA:cUfcf^/Q<,(>dMgUAK-JX[Z[fc-1aNS.g_<_<31K@IP+_;Z@]+NP2CfPd2
eT@b#A#<&1IVgK=XIKD0ITDfYS][)0;J,AWO-+L^8QY/BdJ8W\11X<Ue?^RaJ<&S
J]/O[-+MB^c,8>-M9-#cCON+R;D(<>8@A>eZ2-@Gf+R,^GL>S_]P1&Z<FSG0+<(4
#<=_@XU^5_fRFdG++e?gL1_\ZBVX<>T0KYeC(DP>=+Za6R4/[J^Q#MV?BI4B:=M+
W1/YDBV6:8_URE(.XKW.S>)7AV-6OP\[+5=HXYfdB-_ST;YL2RFBA:;GV7CPAW6[
OD7D2AUR7L)O09>0/(YZBIfWe6PgHRb5UU+,gFY28.BT[bTT02<40>,.L2Y8T8C&
_5a]=(Aa\N^QceIG70bFJ[PJ/JS#M.>1/N52>4_JLK0>]7C/2Y0NF#3@>SEgI/8R
a2XFCD1=1<X(Y3\/,MTD[CK7?[f]BP<P>,5TE/DL74GK/;IQZWg<-5T(OT)-6;]2
0<X<003^WF0;B>fda:Qa0)VC9JKN:>W2)M)KCIJ+;OL&8NW/f(R#7XP2F0PDV3T@
2H\XR^<TXeVD&UD\N0-b[\JFeKS)TEK=F>==Tf->D>::ZKQ9,XAe(dS192=0#f8(
/Z\\c218LMFd@9bb?Xf4;1d<B8O7UPTVRRS#40WY^R;\aJd^.1.JaHZe7MBMd+23
57cUSOCI@6cF>ef&<^GIMY<4I)NTB>WG_Da@fKHVJ(#FbfHEcLYJ+eTHX+W][Z\=
<M/A=COgG6L:&6AMAFfa8HJ7X:N&/1W[.Y,#FR?L0UZ4L7DM49.JZ()<HRfMFSG-
D4/5@\7GeNT5\TH3SC1A#6+>C;ZFVWTY<1.bNZ_c>XQ3P/5RIfebV.59&\B?Y3fN
dLabGR,dD[#]XWVOL3GPY5I](+]M6?e9PII(37[]U0H]CdMWJLc^RL93)\PIA-aI
g4Ze+1eCfZdCbIaUVMUX4I#:.I\C5ba-/\c<Q;=-0a1)O/]CVDeH]SV[CKIKL9;@
ND#>Eb?Jd[L#f+/eU/^M1c/\3I&#1=-F+=S+Ne+gC-:@ad?JZ97U7BU:Q);:KL9Y
2V<829+[bbG(Aa(KAfe>4A=dbEUVGF]G89<X21,BCF+DQ;cP[W79dUFPSeIfOR(.
H]+(+#(_4<#)a<:H.aL3_U@+4+((6Q;U;a#J0CBHCKNXCV2,F>e_.dI_4QQ@L7Lb
M6L-QE4&5G)9=33c=g#7C-6[V-cI]^\\8T#Z6R)Fc_T2C_0[YV.52Oc^(Q9?>+:2
AXUCeP0P@>Q,TKgdF/9:VL>W6+Ae7)4SbLX/H)CSfgMC\\<^E53C+d&S\/E&04:D
Bg-EG,J^UZ(HXA;fTL<CYSL5T)e&fM>7&-[9F4)UWeG0VHWebI\:H\L+^5M@D.8e
V(ggd.R89D=C+^)A8R1\[:L4>Tf2;M9gSbNXGY9X:YK\d36NC>a>3^CKV]4^_W^/
cJQAOeOF=]ZE;DFGM&fPVRD9)bdQd@cNObL.3dT7I4aKC-bQ<\W&#.f]?]TZKV2.
.@6N#,^Q+:PC:AY=J>bMCJ0I)\SNH]9-ePP;>N:5OfMIZ9(f==b4O7>E-&dT?0V3
X#SVgITOXff/@8_ZA_RbOH3UNL-?R[+9f]7?57J;TN.:]DgX@4=(+SgK@1R?eGP3
-3.g9<?G8TPUP+;0_.XL>1?&LC-LE9]H_cI?X0KL9?g<M)?]RTVX0(<>B\=+U#KV
Vfd6-Y8<=OXDaOQ\a4U9O34>X\3\eN#[HGVaV/f.fBANG&Hf8P\@G/4:/dZ-eNGZ
SO:B:H5cZb;0XUE56T8J^WcL48WY]B^-g<NT6<FAd3.8d>?22)XI_V]9DU9[LGD+
T@1E&f(B;Z;@L3?<STWCf=;4(DQ>Rg(ZUF=H5ZW,;]a2)+HS4NU[.W8e^[1fg\9=
.,N2[ARJfRLTRD\XQ\Q8R2P67Qe4SKI9WeQM..LEA4NWLUBX)#)ZB(;3Z=1>G\0R
=5KeSBDF-b8dDfM2[_<7bJ5M(fK:>a#-Y]-AEV7F)AZPXCHRUD2#;0O3aL5L9c=J
RH?e_V_3:O4TLTLZf-2>S:FHa=>:<L#S6BEeaaPMQ]HD59N#+8D6>;>bV0D:W<DS
)+/cJVLI,W>aSL(_EHIDLBbV1;]^>0MVIIQW@eYT1AcSP+L9[#EDE.Cf:?_,g1cY
(cM)P4IAAb:S9e5d+RU_/VfWYD(bWaUA9O@NG_=_HHSHbVZ.JME0/+NRQa1=,=gA
V7<eAVH@D0]C#)4)OSPG^<gA5[5PfT,G4.BdaZO73EC25LBBA+-<OZc5A5XKXg=C
<WZ16T\C^(R8WcUYO(egKALDK?5P[C;dSYLCX@X0<a_a6Y[/:+Q9gL41eABId3P@
+B7,.E-7CX=L]:9)3bJ)8B?f/MO6:970)Xf1RJHS_KOF1Xf.ZbGF<U98/1g)ZB1b
>6@0R=\VOLEU8BdCfJY(Gb)I?/e7eUS/UeWU]#]/B0e:V:fEBQ75P(=^8M1?G.bb
ZL<(7YK,U>\Aa,=.6D?AEE;U+gDI@)UNUF3K9c:aKJ0S6g)g<Q:A\@I0I,IUUf-?
K]KW7W,@-Rg)SQI0;WcNL[NcPddWAF:].f#A6Z@43AC]D5CLLZQ1XZZ,eXgXaBPN
-MSZYPG#O1823X;1;9[_B8J0W4?LH:@7?fKE<8^9ZaZ?FY^XSa-K]:SFK[Ke_]9+
9)TME&-HdXXVKJ\P(Xg@E=V^B.MQaDJcTJf</,D?>Y7e71,cOC]f&f/JT+6#/\6b
\)<6YV3KbQfG47=OHcII3RXaC;?cEa@I^^>#5?SC\0A)CL&<GX.\NW\<9NP@@eWY
:KIJ2Cb,aH>W^ZQ)<Ua?M3U0K:bGdTEc2HFL11=4;9B9dI091;;KAV/PUX&5QHQB
4/LPF71b7e]@?6>##+W3H91=gSZ>XC6>HeI[JU5]\e[3Q&dA:X(MJdfRH@512HX5
W_[c.6RO?\LDHULK80G^BFfaK+8O_#V7#[)FO-W1[=dL&DJNZS\X>9BS>0cG.+@1
CSC=^HJWXUC=?+JU0(Y_B_]H<V3aMa9U9ZNd:cPYf;(Y]1g&DF&,&Y2E_bJ7dXMd
d<L2KbB6J,;c,&ZI,J\F,\^>:#=4/ZNY^V,=M@U&T@<V@K-gP&Q@cWP+@;;X;b72
K4GJL,E78/6.FB;^e1S7gK_8b72+]?0>95+5FeEc#;W7EAeY0#9NUgMP=[N8-A]-
?F.&]Ag,R)PWGGIXQU/4HX&C;d8BT:5+8OWF-17&GQb^MZ)&a1&b.T\8ML):NXBP
_:J&I7.U_7IdPEA(127LA@#?(A2(U[NaQ6,dT2c)P7f/2OQC/a/M42+g#&V3=[DK
>e,[S1OXE9=4E&QM2P).?2R.Q:ODe1ZcgDZW?(@]NYICQ(cTL:C,OZd7MT&d,2SI
(SG-SM-Rd=+&=.0LRgSR96_2W],:U[YCHV<IXcEXJ0MQJY@URC;OV]QB?>U[3d2Y
\ZUeI>3JM+9W\Gc3EQQeV.QcZD.EdUgH[WXY)Ec32&F2-3<-S[F/c+P><\[H>\QI
/^\3.2R>eY^db0a:0<eW5Ac:f34H,TdWVL8QQa\7V&afJ.ILUZ>>)5VP5_RH9(3<
N)O^<#dYR1>N/+B5PaFRC83>KI9da7eD/EY&]?HDgVZM:4g_Od1?JL-afY6T&VK<
ebT;99[;O7)Y/+V)PU^4fZ;X&D]Y6AIIT[Q?8=?(1ML(?0R,(QAKcN^-,Ze/82f&
5ZL8M8#eV66,c&+/6^<H1.FO4?La3^A,S(E/^UDQ]N+_+AFCb-R;\V?PF;Gfb5>P
X#CP:\[a8[?b\U;9N4N&N]dC&M&R2-G8DQfNJSH/Q9[7.AF+0[83P/Q?9T0PT/<(
4_L-@VC@;L.R14]UH\D&f,?7X50I^,FVVe_>AHU^SB6RSS6171)4L\:68_NI,baK
fY_5gFc8+GDgYFVf?BR4.\@^#6;_3MS3]&Y7bGC&N.=C@3WEBe7Q&dKD^7;aMTJ/
@Bc:U[E3X5B^O;f8A;/LZ4C7b(XX]CVLC9:#a&S<5+G3)@Z9Y&c<@\37BZ_QI6YM
GFGXL#PQa6+XO0T--c5N?L=MCDMHcIR0^[RGIY>\9L_+IT_O85PR/T\+ZL]\MQ9g
95EQA]P^_5KC/MN=aW+F-C)U9GG6\A&@#0E-A0,)SDUHR1C^2>Z@SbM;3eM(2:V.
XWQ&AI>6VFea#^SG83PK4S?B:W_8V#50K5/R5QLfG:U0P2&R)FG+CF-C[?CJ;(R_
<B#;.65?I5fBJG<#Y<ZL27bNEX>C\PTH<O^4]]Y;J;TXT_,Lc;(/dY^Y0/(&E1E:
97BY9;B4?Z@:R]7E(XZ><V@Gd-H_,NXS^c-dg4;?]f9=d:@,BbAN?7--?A].E1U+
C]]AUX<G8M6G&^f[&_=F+0M8/9ZVfMTYELg\ZCL#)g36I_#<5fUeRJAWddDD[Fg)
]C+YWMZ#[d+@WDL(.=IH89Q\_@:a&YKO5Q/:MHTL,-8Qd8e>[dIR9J2,ZI&Z9A+_
8@LCFZQR_NebXLdVXW36<b1494H46FWD]Z_A^,-?_H5<=J^;V/[+YAEe?UK^)cY\
g:/-GD\+O9JM^ETP:?F\.HD/e(3ZfS8?9:WQ>Y@EO4@4+D_eDB45e_/V_SOQ4,c[
76Y<F^PBEQKc<f3CK7^Q:0bDZOYJ-0A:2G>)-IfY+/QD#AVd9R5HX:BSKV8#CBa&
^H95,2BEV,NHRTY0c@F9(5@+M.RQAY:8dHG/Z04ZHX4HDXWLD6#8f(M#E];aD9L@
)?g,MSA-266aH;FMO^>E3Yf28Q07P@KT<43.=B.PX7UBBA=L&C<&?WLZ4c5T8Kf)
7ZC4[MYS?W86>9AfQSJBaKfY&FH80_&P4,:Ifa@EY94,99:G?Z/+W>0WRA[UXLd8
T(5F_3:A9.=dfQU[0^Fec(f93P#]3K9.c,#>Jg>eAY0fQ0bg)P@bb(e]HEJ^F/Yg
(>c:<f3gC^Ca;9+UJg(\/d,72AfYK3>Bb-e5,\EBM(F-<X?]Q<8>UVS9BK5HdP+8
WfHJ@(<QK1cFBC6\7ES/]8F8NM\RI[.M,7)(+SGaW)I<[,1Ge>8PEfeVeN>^)DPF
d2EEB/YI68T4d:MDfHK]BfQ;\D7O>g3N5P1PCGGg--=_]QG;&LBHRE)P43<^+KP>
AG_1US,Y#CY.6f5=[>5_PVE?X_;683YV(2[<\.IVA.>-SBe0N#:\fH;Q6)TT1IB+
)WcQQU_.,f15g\]2K?@H,3WId36,F0?d9c:.G7OY6IX[0>O642AIN5TC]:+#6>)\
5\&YcecZ3^C_HQ_cSVTZYNZ/S>F@QU\_S-2R2]G]cW96E43@AGX&OcXX(47[5.8[
3G6KE7D#.Y9R+LbKY@RKRTGWNbRZ98;:3BJ-d)7O4DbgE<IHK\4Eb@_J[cT67feN
ZK[R-1b]EZDRg.#41-4&2J8XY2+cH(7=_I_8[F9&([QJaOfM8ceg_:Yc,,Q+@;f=
NDaEQ5g;E;5+>NbW37II_)a7FKO7O9V]L(_S3J-c7[JDQ@J[UZN<L;M2:)G/89&(
_/:Z\<9d-F4c=Z)@eC?&9@X8=S29)5PRYR0:d:GH&R9\OEeLXLfJ>-)aA<5LB3<f
JaQ+U(GV]\U2^HaX^?C9G;Q?Q,2d4.2,1H-Be)RB8Z6;T6CG+THZ6TTGQg1Nf:\2
-\QOC+0&AeSc]/WPW]^Z9JJE8FC&K-)(aU3QPd4H+]VE&&I73)7KNSIB5;a..[O-
W=4Q35_M@FU=6DLU?.]X:,BUE83)3aJ6[b36S@;7E5XgKWgd;?WKC_dc:J7_CP31
L-KeC10fE>H)2;Na&WRd@b,<ST2fMB[Y1?DR_GJYa>MAPR0@_+P2-fG[\@/XXa@6
LU,C?#JN94[7E5ef1,ERV\I,7J5\5>B/_fG-&]ce:)/N7S^bBb4WgOfe1TITJUB@
TGRGZ>.b/=C+FLUW&c20FJ[6#@KGRCVg(WRb#IQ;acS8-]\:UE?d-]eG^6)[K#c&
E?c-T0Og0gZYTO#)(+F>eS21ZV+g=3_CU)M[[HI,g3N2AR)SC5dU><VA?/R1D=47
71@WBJ^R,T7JEFMaR::?-fa@Bf(8,L)_VQ[AS(+VPH,D/L:H&CbQ<XGGFOKd)OL;
YM,1:-Xf(T1/6184KH0MZT4TgQCEM)VGVa]C<77>G#+6R6VZ,Q,:O66BEG(;&-Vc
C,2BUU<4.I(OC6#(K00V,.5^C[]6?;f0bMWJ6M_)f^M_^H#4FN5JbON2Q5J&[I9^
2JLdWCN-f>U1WHcBBIb3<Q<Q/1=5]&5:J-S,S4O5gcY.1gE,ZeaaL19&0S]XMLO^
?Ree0U4@_#F7C:OE.??L2M(cK5C4V>Ofg-F=Ma@5caF(\gEIAc)?e-R(3?Y@+[_f
L@\X#HVO57;X=>1fB&XW]Y>EF;d[:T+<SD,HgM+BO1(eFGR[].-/E+G7eNDPM<98
.RSF]CD4G_L6X]X21-_[+d8>HF_1dT.M7JXJ+Z5@#-U(a/IBQ]0eK13[^)Y1:L2W
cY8\bPA#(Z4X2-8EL1f&L+-dG>A52,?fJ2>d[d=K23FMc:#N-d??Nb\+0AGQ0;OH
,)Q)Za?2EXBg<;CD&Wg=3C=5LX7^&OHI^;#KB/agKbAB.1aK2FHT(;#N6egGD.7-
EACINX?@LcM32[+JBG+44+]&(\CJ3/K+Y9.-9BI:YD,cN+H1)_0YTGW;2aELbH3U
U^VWOP]GH2=?FgGQDP(Gc<N99cZ=Hd&W_:D5FCY1)B^e#I7T(L>^8f:=ENE\.=V2
[>0BZ^1>CGF)^-fVbH@7MR02JLIFH_6/,g9[.[1;XD4S:&E@e5[@LE&.gTX>H<a+
-.J0VQV;+U)0YD9G7Qf<#[Y^P.H1:@UFa/bF?[H1<_8S6^>YL]F_a<db?B]E,=g;
L;,-ZP@JX0(6+FXY)(gAYXaHGg^c^NJT;1J?\Xe)Wf\f)E463TP&LJ:198PM.b;T
86:E?G\P#+/.)&<);P:X1)@bGCEW8/V503^Xd@[2FfZ>-6=JV=K=MZE=-WF<1Ab6
:]?+MIXI8]g/G1fM&WZ4#C/A/RR;Y\[fHADZD1a08Ff@0AH/&?JI_PM2A99WX4G&
/3^)SMX43J83LZ<d.7>?IU3c2SE9XEN\<bPY6.WBE5WIaI375LbKbU.Ea([C@_?G
OMHVRAfZNb7.D]/(<8eMSJS6_A7D+Y@&[CgYA+^fKS?BcGXG=4I=,YXFaX>A+T:[
\e6c,E@\+/\5daR4U_T)XOb]PAc-ONg.3bKeR(QbYa,&UG)?fX:OSf.TNXWVBGU?
_FZ(:)MM7GbOIc0NH4cK-<W:&7W\-\4YVc:[:IO(;A05KXgCa,&8XL9:V#5<.UFX
86=_RX/F:G</VYCIB6_4+6S9-@;JRQ53JM^)QZ/I#4^93e::S3O[7)dSS,W]07L7
d,L6<Ze05,]9Mf/]M(-;RRGS?#PW^?I^dZ<1(3)3cb/7F9+<^<X^eZPU&=S8+CQ/
40].aB-g]W7d=)?L<37U2U_H#<ODZ-O7T1G1_P7M:B(LH#?&NL0XD[(:VI;9=>2<
aI#[TB8\A&D39.)7_4:2ZLNN/89\2.DCB?+YH1;[#_P+M]GJ;Wd7YC3;I^f6_^1@
Pc.LQ5K?ERBfA@2I7_RMgTG/g7U>8HDaf-:)U,-cIHS^?DDTc0(G:R_5QO6EJQeB
\d=\8(,3G16[dJSPH]:[BG25PGV/)H+\H.JAEgTSKCE9.&Rae7E.48eZMN=Z<^9\
[fRD6POA\LFT]5c.O7LgDT?&7\+LDN@Y=9<P/8fc3:DdP[>-#eD96-b;X9I_Ugf.
B<K>I6=L0d@J8W8?QL;)a>C9NQ_1_1Q&>#:?b<,3EX(g]J+,^MCY#1.A&/7097:B
M(8[Nd;8<dYF82-80#MSP5#V0:WY90NYbS_FA6\Y:g15WTQD4CbA9S6M>Hfa8UY\
H;U]V&F(KH0ec9@_&>:fI03V56B\[8I-3H=HLH16MYJF)\:HS?28B/bL5Y?Y(4#D
LT-TR&O2A@+U)7K-IV,5ed+aW<9+Zd9&dQDe58T42<BNH&/U1C#(?IXN;\:@Gd4)
\;MVT/U7#R(#gdZT1OBKZMR5H-)<T&UEc<A<A<-ABML\Q3c_Nf12OI-)D?+=XD89
F(TVBCcT5?T8777S:(eU,b1IO>BAX_Wd\-MMHT8deGTQD+EDdS;2cE+f6P3b8/(7
F?ND7>BEO&(5WVN+J_]YB^.Zd08F/\?>@Ofdf:8_&fgg^cQ=a(QGE\;WYe8P7DeR
+Dg1@)[[?.B]Kg;:(V[2.5-I[]OBBMG^#f()W<3A\?1K@cPYO&=]Nbb8V5]82)H_
<>05.J0Z1XM(LCBS+3^\<;gAbGU5>X8K+Ebb,;g54;&V[W?R61H@S7]?>Sb;NF@4
R2FGG9/,RLcDI_>C+6_@gUNaX^<K\C0T,)?AI_IZ1\_6?]VHb63G<AaagA50/?X0
GC#H/[)8JK=74_]WH.<NF@&-QC#DbfI#POWZ>UCS/#c6Sd&@3fV^C.-,T)=)?LM\
FTf\JPe+?W>]bQD^QQ5/H;L<^gdL(IRb64IM+Eg?Ve55X/Q+@8BJaaeRCbT(X@]D
R@=bW0Y,3@A/GBBdg]c:V:)dD3Z]E1\Z?,=#cQ0bcIC38H?PWI404aUE:L95bAg5
)TDeDEX:f]#R:a+X5L0[BV9[e239Wefa,6I<#HJ0/&AISY#<W8S]&Y23S(UGPg1B
?a(7\D<B#LNBN[g/>[X+6a\HG0E0Ca1(TGXbOfC8e-\,XD#^J(B?L/FO49=LQ&V(
RFSNI[[JHcZL/e9C18c)BJ)=69N9D/@7M@)/,IG;LDfIJ<<Fg1^Y1N_J7^4+>9YS
I#908T6E^f9)e(QZW<gQA?&4U[c&bXb8QgDObP]C_^?gbNLV:1HJ6ZGRSM7K#AEF
G<X+8KXL#ISJJ?:#A(7]^:.M^,@#B#Q=Z2+6A^L=Jg<^809R5K;U1]@_+]>9^[IS
;HGH0\DG3(4&6g>0^QD-a0cAQgV=SX[ZZ>545U2K3A?(^+JgY8IA>1@8HC?1_,E:
))-Q]72fN2;D78EgA5O[ab?7/5+&LY?fdaYGP;UPTCHJ-GG[5^dPYLRV0>2a;]FW
NCE=C3^G&(MQeQUUc-3HJZ,MN(+>\7eQDW4Pb&G5OY[L.[R),e7Z-OVK2fOQ^#K^
F5K2a4?C\W:,a9:H/ge328-b82(cXW/g=)JgP_N#FeHG_RC[)=/1EadO@;?5W-f:
[+N+],ZOd?AM#SOfC?U4U4)4GeXb6cH8SY?]#TOPKA795TGd1J\g&44;^U13Z+[<
(K3U42T1T/?a^<+NWeDQG36@1Aa>##OP2Q-=&NL:,[PO^3R8PfV#;LNXUAJeUJ(P
G4X=([2F?V/FadD?b)gFEQWS^IRC@N<D-89DdOUI0W3HS40?-TTVg4F]13=+>-W5
5YT_^:=g,FBDXW<-W5:>bG&dF3^4W[J=F&O.G]^L=IXIAUXEOU3NfO:[DVaeTaVP
f9af:T##2IUU6+\4BUEO&@FO\<.:[+0Bf2U&.gVS@,[ZI[8/R)c[MRSeCEVLaAOJ
W<?/UK.K[E>_=bU7Y.Q@1?B&#/gIWT?&>0?d2d>SFO05Ec/I3=,2+5=;MV0L?,ZF
&=0&VBbY(EC\<-d&6;0;#A4PcVWG1TAKY19)3CM?AdRE#ea>;Rc)J2_]Ka1]aT>#
[;L(F)NCWY9(g]E)aKddC(,c,b0fCZQYg>&7g);T<e0cIZE,30HU3+C)^D4E8V1c
G+JGW)@3f?GPd4M#d&T42AfCP:&,c33cC4_&,/E6I:2GD>fHU.,0^VPU8#_8b?52
#dV=S+0DbPX8cL(.5b5/#7C^?eDMOW?T/90>Y]PX=aH?<9JeD1G(Y(N22aIdLYTB
]GdD-V@G<1fcKMMP@,KK]&aO?GRUVW#?8<\.J>B@EP9)5Y#W,:ZMXb4)Cb5M=HA>
SPWMX?<0(0OMb2.XY[V-=/CA]5QVc?BN<-Q)@Z,aLTV.0)57S4gX;9A-J4gZ>FLR
#&^5=55IP,6<c)6>edcHXF-Wf;L+JE/OF\a8HGDIYccF]@G+H_DB[+5Gea,Ua06\
#M7J0>KN8ZS76HV2.D2X?_e/D?Yb6+I?(8d,?=^XP@>H7)K2<a,]WBQ:M^8O]2#D
_JfQZb>PB>fM(WDJRA;+g;P<0NM.-TL;^.#;)\bB#9AV@USeQX(34?+5)>^?.EXO
>\>e9MaeeLJgG1#9HaU^,XEO?a#Y4NA>ff&gdML,XHO>L5SbS5;9GQ2a^.B6H7WQ
/03cE]<787-g;,2=?c(QYJf0Y0B=9&V4VYQXcZQL;fJH(ff3KN5W=[8=MNb&&C=M
+1R#WgZWX7CL8TA9E9<S^PaV3H:[&_VGfgMBbOV6aR_9NGJS+WHCXI9V,HKGdZ[e
&Q[8f<D1gV4FOMSU.[,d2<]D&&(N;B5Z\NJbN6E7]-G+;&-U3@LE>?8(E7+ET:>1
V>cFJDT9UEK^@+6HKJODD4T-O#4],N_TCMdb:9O)gc[5JWc^9T;<I1D4W,b+R,ND
1M4UW=USdMe0\JDG-JCb1&@R30eLGR90[3FBbbSb343MV6#JBP[LH;.]FJA.=.c_
;98#Qa]3RL6+/=X9H,M>6,3C>eQe26@dI:6J76aG<R[BF@>,c8d_&?ZBa5/c)aCU
/F.)4e^YAS]..Y.We:;^Qd;#:K7N?+CGHZc/N<LYdGCdJV#EX)8P56HcI.-/9K,K
9eZFIaDD_,]M50G9>UT_,3]O+WS.PO0S\V#YeQEc3Z,PV^VGMHUVS^]ZUSY]<@67
1(/OI8dEd&\TgC8AdfcST@d7-R9\]>H/gQgV.,SW#DQa#7?2JXRNZAI+>7f:U(=N
6XHA;].(:@+HFD]1+JTgM[faa870#6UH970\#TU460UX1AOO4EY]D,XA,26dZGPI
<6e/1]85;d=ZHSgC-Abe8J93<WLfZR2W-^XJ27&+[.afDFL,JI6ca674WdBS@4U#
>/QYTUMa^Ed0DY:E&@\6N:-LQHZX;^^aTX6(,=1/-g4YF7KIQCd1M[\YFYI]&DDZ
,PKC^<+:X\8_WV<BS=^a@R:4O6(\Y21=&1=NM#D30c)BOS=AJWK[YV#+5YW+RB?6
SY-I3=WD@O5U,\e,BOU>D[;aW.:0#0V.:5HRL^3;R(/6:N(_050U,Q>/6KVP@52F
.X<.<5M<f_8,Lc9CeO#f)Vc,8N4.8bX[?\E4M&VVJI3-T>55@SF=2B>U+APc,2DZ
9+UF2_F>aZ]&#ZM].11BQ?&I(dXeAa4@VPDN9?FEC^MeS?bT9@eL0W-13OKaPC9C
9S[4Ga:8f?>.fTXF(7X.?5(M/-E]>]L()b>^TW9WbII+8?cOK1HA@7NFa3-74X0?
N#Q86H1UNV2?aH/(LZ2d#cL1]6?.];LV_N(,[X./)]D,.X]VY>]-feW/,G:P\d)3
O.ZdKf/:6A<3f8O_eO62U9#Z7/Q-,DS5LO;3J6/a:a&^/T,D+TRdZ7W14_8/Cb8J
D,9S5C<)c6aQN?F@&\&-?9UJ@4_fHE3U(HQS43S9KV#L8<<,OEcNaKP?80;C;<KX
W@#\XN0<_Z8?3@_Z<<>@X@L;#,N=^4dNGS/D/VRJ03_MUd2_-P/5L0Db\W,TD1[J
_[.cEA>.23411<@5#=/?LSO8B(0S.eIL^?Sd:aT&bW^g2Q]A;T-_TdH>U-f623]F
<HC7NDRa#IHU5++-#,YK#OJeS60TYK>7(d58J?)PI=3OG.aC@C-fZe1(W;2+X5e\
F@[cF&+=cXQdP&c]KCfPD_g#RP3C8I,TGH&4S?WZ/aPBGZGX7IG_0/B99H-0\>1R
BER4J3=dV=71@QgCd-KMHP^90(eXHJF4AQIJf-;Y+cKO45#&T05BKGMZZ)9IR9PL
S,6X#4V7]CI8(GcIca?R+DJEVK_b10c.;/LTN2;TQJQB4);YW:#1Yd;K>984#Y>3
M>7LbYeO9;LbfYL9+CWRY.d[6=7Ic\[T&f[K\bUI]2<O(IdHZ97>7g.bF76+bZ;W
9QB]L)]FCAY9W03)g,-.//NX.T7IID[bV8=c[NRCcJK?[TWYP3=G1I0VdKE?e#)W
#1>.24+2J8FF(c@D8<(D1-#-NHWJ&=b]4A=Q]T[4-OI-F]eeTVB^9<?GR2(9Q313
4KEd5OJFC\KQb.YCS3.:5@3Z^[aEbg=S/)FX]VYcS^=HYLZ>DP(7Wd,e]0L3)T(C
G\4-Y08gP-Gb(KJ(9]DS^[ZYT@CL,CJ>7Vc=-Fg+TLF^E>3Sg\PQV#M(_6P[3[21
Z<c&HD7MF/?[b^>HR1)U.(]9SBI.6NF+31VQeY1+=0#AUTG=VYZOa.LQ75F(&6Mf
/GX2?[cZK1023:JJcUVNce+O_?57ZB8cd/QHDbecd=TRP@/6)OYTdBRd:.aWc@/;
W?23BMaHU=WX,^VUV@L&SD(M-=@>,1e9.=,B->@\RWDW^dK#O^-+C]HH.FEX>^_B
(&]1IA,7M/A+d&DSBYUI72\,85KGD(6O<gQ\Q9);^,XX22)&2DQERX;K/_1W_W,M
)6W<?O?g-d@4GG1gC_S5BD+RL3^(R]99UD:];E[OT5a43[#6F]YUcdg4:<bL:&OS
6Q\IRSN3_Hcgb#7XY6T3V,Q7=cG&RBR\H(^bY1[:P^&S_E[?-[CUJ8N<Nbe58XI:
0:gW+F>&I/QbB>[RZ+Re?dU,Z@DOaEP;@@@WF1+]c\A1UZ&cG1HVgQ[4bDJL=XP/
:XWDV_b.@4<6+b2KQX(2F@8K6NEA,e<O.AJ&M(CS,+-R(YVJ9GCQAE7A38X0KP:X
<T=M+TD+6-VU?>&2Fg-Hb5:WV=;HKL.^>F1FPQ(1)d.1<;eBc/f9f9T\6@\Q)d6.
2O3AD^(I[L1,DYDWHX=4DBD<G_b+Mg^TD3=E:6ceUY&4T4OgZOHH<d0,^&9>:d/&
8V2LA^8WD<7MB4VI7GVP.NELDW(cWJf1]Xa]>MX0O5(KQ:YQ/AU]Aa&R/E4J1W8^
B4I<R556D=?(K^6K]/YUL6KD\3Qf@d/N;:NFHDV5,J^AP/dQM>RR9X6Ecf_(AX+e
QMdaKeS+]VN615P3].-eUI)UUBPDUA.>OPV;^1QG\O^VM@.PJ4QTIQ(6FO2<bPP(
9@=dQVQRA(O]>3.DR9^MIBe9NaUc.C28GY\4H6D47+3EQNH96D,A#SP2\6B,2QcJ
<(^@.bLfF33_/J?6.2fM(;dHe)<\==.:LVf(Ma;[>bEZZNg5Idf=,cQHJL],_T-e
8TF0cR<YXD>2aUI5L5AeBf9D5:#EY/\L?8@,/Zg8X3-#^4P29C-/M1OTCN@4.JKA
-9.7J9+@L549B38-Da(5^PO+(.E99&:_3C[FU,HQ5aE6#^U9S+7#P18+6;[NGa0E
B.FFGFc4B+RCbLQWaQ\T1gg3K+A,KLcI:S7I+>HO1-,4W#\)&cUF?8<(+RIT0.0\
:D2TWL7:;V4Gg&K/W\<;8>QK.>I33DD<;45@32=9Vb9-++[FBHEcP?WA9#=9b:[P
29[N+.2VOcG:YV7Z3#]ZG(0NMA3>-2Nd@>28J3&<UA(QPN+QN<<QR8E:SN(523VW
S4X70#4TZ[U4P<C9E0AV&:G.a6-1M](PPJPIEB&.N\YSTCZfEF<5FbAC>E0O77.0
GDeFG<;V+bAC=XH<YBAPbfFA(dTPL4<Xcc;NMcNJ@H7Hf2=#M8(U0M/;ZS_>+JT?
3IB=I,1=G7]D&JD.AZe?;5CD>=/XKL2(QX2MW./;OM3PF(EY/Rec3.gA4-1OKJ]S
ED9J8;H[\&.U@dbOHgJU++8CZPD)P?DR:06SW(9(bA2B<C4BYHYdLQYRHQ;DFSAL
(>_A+BIM]U=0TGP:>-XCT/>HUD,1:GDM/J#E[1OPFR?<6C(O8F4T?K7:<5309K1D
]d9748UC.)_0Y0653f?3UF]0W>1+FUY+48V^cHU0>N]cI-GF6\=a_16R3_bg[E3(
G7M>=Icc;671?[Z.dK<W0-JW[6\8g4W\@DBcaa@<@2<#A?[XLX=Y;J>E2g0:4^9L
23>2)7WMgbJ?=_0P1^SgTHT,/U3G]gT^=6DWEISR55=d:#?PYM#GTc048^U)aAL]
<2K]eV26E_e)eA_DJNL@-V0Dc,D7(E>SK@;.WW/]S5BbB#=65JM([WO>0F[;7d,W
@RKW=>gBCeYMVH<CPEN_IBO-\5M==O_[e4^Pe;?eI=_;GE)2gB7\e1PG.Q(,A&,R
XQ+QO@\7:3/ND<OKeWTg;<(L)3JOD&Z#G6,R=4_K,(7PVf,W,dbDCgPO4Ze(W0^Q
g-/A.JeHL_VYFXddB]]-TaT\5cW3eO<F#?6AJ<IMU\Q3ND[KE^C?G(g>3;0@+TeX
-Hd[N\RR<&-O_N)2e;@FW9JT0K[/0<1H#NO^fOf>P,Q)acCM[ZYCE&[GedI,:R5U
gY1g6-b\Of<WCHWK94WAN3:VfGe7MWaU;BH@dd,Oa3^<_e;>K\X>21;7b\G:00(g
C7K:8T@S2FBN7:P7:dRQ1RYOYeOMNJ_@2COIbc\-J]C6LR&I\YNRb<VccMZW=GQR
E#1gZIDe#+2+_Xe>,@^E]Z3&-0,-K2\+/@c?cVVRXL9g3(01P6B._BU=K@<ad&&_
81F]/G?Y?8];9BLd=]PHX6fcGbDC>77BYZ?W5GROC7X(]8D8()a8@9B3@5LES447
W-Z5CPTIK;f-,7e+7.]0[f;K;5=1(Ma5&X=2XIOfMVRf-(CEKLBDdG/<d_A+,ACM
(.WLF69QP/S\^/9,<3J9HGB>HAT=Ed4&E&LdO=;OOYM+T=]/O_);I;b=OcDAUQ3T
Le+FaWcYZ]VR8/\R#?TRS.c:C>3g)OYPEdDRcCCKO>O^S&AKUZ+d.+_,AIMDT<aI
_^e(MCG8N-e(D8J]03_Zg,HQVf^9R^6]5G[>4R-329@9Ag::=a91Z)M,TAc^GNCA
cJ?PVSfJdC.UcQ^H,^^eO+J:bO/E6JG^?HR@3-O;;Rb+\MbD[(YC#aJI81J;\W9K
9(L23TcQb0SAD9>?bN1T3A7YgCWFN5f)<HUYb98-WNaE#5[;VLCJ?=AW7BNWE[98T$
`endprotected



`ifdef SVT_VMM_TECHNOLOGY
  typedef vmm_channel_typed#(svt_axi_slave_transaction) svt_axi_slave_transaction_channel;
  typedef vmm_channel_typed#(svt_axi_slave_transaction) svt_axi_slave_input_port_type;
  `vmm_atomic_gen(svt_axi_slave_transaction, "VMM (Atomic) Generator for svt_axi_slave_transaction data objects")
  `vmm_scenario_gen(svt_axi_slave_transaction, "VMM (Scenario) Generator for svt_axi_slave_transaction data objects")
`endif 


`endif // GUARD_SVT_AXI_SLAVE_TRANSACTION_SV
