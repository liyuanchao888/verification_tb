//===============================================================
//Copyright (c): ALL rights reserved. 
//                                                                 
//  Create by:
//      Email:
//       Date:
//   Filename:
//Description:
//    Version:
//Last Change:
//                                                                 
//===============================================================
                                                                 
`ifndef CHIP_DEFINE__SV

`include "apb_if.sv"
`include "spi_if.sv"
`include "apb_pkg.sv"
`include "apb_slave.sv"

import apb_pkg::*;


`define CHIP_DEFINE__SV
`endif
