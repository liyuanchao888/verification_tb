
`ifndef GUARD_SVT_AHB_ARBITER_COMMON_SV
`define GUARD_SVT_AHB_ARBITER_COMMON_SV

`include "svt_ahb_defines.svi"

             
typedef class svt_ahb_arbiter;
typedef class svt_ahb_bus_env;


`protected
aCVJeK676bCWEJC9DX/c.^><@M-9(0]E4aOO90CA(G_6&cd-.^Zc.)H6G[7=PU-S
>6<<3?A?6AQ;<bL(]QI:e,;a>][98B_4,+E1KdCU5^Xg@[&0P[^f4MBZ7_FLC]g?
Tg;N@Z5Kc5/=4,J]>=FDIR->+;7dG>d2M#^&24.,]f905>[ZM9MUa[?aN2RTf8E\
]M3:2?Z0/([58&T1[YbU9g7Vgc-?2R:_UTTH6Bff8K8)99</ZO/O^:fK(gZIQ^Y]
a<Sf9b-/E?94]7b.):dTc8#_+F(F2(;_@d9F8=)?9e35X>TH)+eE52cP:RT2Q7-8
L8(8/27OQY/9^b>#=CBB(S:7VT]&Bb.Z+]MUZ/Ic7K(g1GEG01_91P7?^:G=4E96
BXbI/C-O:c__JCdS/N:1O1\_VC;B9/>[D_a?+fLS?5K.OTebUK(>+/<[O@2#CZ;8
-:X-Z?OMR8>,HXL_DS^M8VBfLNXW]^0GX:A5X-^eHO9(H7M]U^R4;2PC[=c,Q&0-
&FOY8c<)L3];3J)1MB#C9#dHce^?gM9Ye@g5^(AQ:.WSc]8\V/:>HV.CRF-?,be3
Q;+VTMZ-RgHGWF70QI^0<1GKbG<2:W_^fU<B5TB\][A,K5/G]W]DNc-&gXeBMT0M
?J<Dc?&e3gDBe;Y+Mf7=O3\ND/&#;I)c1Y4LBL^G,IW]?M^ad9@WXW\EG/.BA..X
MRBZVfB9_R>)a/F^PJWK^,;OPAY@)4BC0(LOOPc(g_]Y:J&:P7=]IMF-C09_L>S#
;CFIR6:gf8BR[LTY&gV(-_5R;=#37]G7PSb79Pc-A#S:BJC)7[Od)M+J3g-+G?BU
gMZF(J5+61Fda9F[0GNR+\&Te^[4<.U0F&&AT^@^8b@BXFD+N_-IbOgM^D#,^N)P
=HdQ+U?J[Q.\HGd;LO,GCb/QCf=?;WRBg&R[?:fTaCK,DV7UbU1Y,=U?^_M8BPD+
/>65L4-bO/M[?3HY0^b92C<.3P;&64XNCF4@8S3,6KACA333bG;L3+F76.FD3:3^
[YE&@&;8EfP(1))9EBOf9\T&g)aGSS82U=/G&=C3CL5f3LFNGZ\9SRd,;0.23</2
(>HTc&6A44XVRHTRE]#bI2>[-b);LRTYY:/.cN0MKUP)1He_gU&\7Xg:6O6&[>;9
:S2GWAb092R:-D0d#.dXP#B8N]OM/e;@cBe/84,fTFf(B.3[4M^GcbcE(?f-PM[7
>dG]]#R3L<OX9U_PbB3\Ce=bM(L_SbG_Q=IM4G0[U@W,>,fI=gQU[PCICQ:9W?=G
)YJ:>43098X_[Vg^+OZ8cc:G45ML.U;:_O\NSSI?&A\)X_:@,2>KW;RLH\WbU<^+
d:84H\.5H9OPOX9L0>8-7=ZV^SXDAdb1bc=+N:_@CSaLbe7XdgZ(&FID23e>R[aI
11[Ec#/Fa&e\b-b@DWAP7]8CSIa)W75._&aK,(+61Cgb;Rb2d:_+.;OB&6P7XW0d
^(Se7AcPNb?g#;04^NVY1fcBG\Q_IZ+]4.:RFAH_UNgc;7S:UN,B<<gD#)PPL/KO
\^[JPT6HLQd<+#6=M<U??GUVX@K4(MGMW#H83/^DP8HV712>>63cI9.I219T@&<:
P@J0ZGWS:T^8W<0ZO5033SA5>#+>MKT=eaURX//+&YAQ?]X:g),g\9QZb6f_N?M4
\ca)gKDX]Kf#4Y9UYOgV\#e:c69)T&@Dg_STE?1>4=a?AUb)RUO5DOGU.RFQ&=g^
DI9+a:SV(J,-F^S=T5VUY:[-7\\Yf;R\^a5@2C@E@edV<79B1XNYN2-Veb=&G4#P
Bc-aVKZ\ZK+\+[K2f;]UMZbH^,43]V(QAQ#F#>IHbXgT\WIMJOJGAMT(>QBPV.2.
LY\bAQ-16?K=B#afMV@bI_CgTGULD;G5_^(UN<bfVa8O6-)Z;69:U)dM2],5J&L_
EZLL/_<<COVgNWK2EOV67+QY_R1;U[WBQc87K8RD,dY+9SQ&;K+^7L.;6[,ZRa5X
,)X14#S+4#4>+EW.3U==#dIYAa79WfP2DL&OcV1E+D<D#(AG:.5]#O28>4+TXND,
9;LNA?#&B#)XG,QP.,A-P8S2^7ITC/?F;HYJO.8+VSD>4g-H1J_a([\5=6K-+[fC
+/5)GaNa)H[.AD@]238+K25fgIL[76@Z0cV+Z&NU)5VEJ.Y1A3Y8J[F68R#LJ^aS
]/IRJNY.L]8BE-A_?TQ#QSG[/0abd0#eG/:.5;QdDZ)Q//E/;K6[<^IQJDcZYIgX
b3ZWHV[@O#ITB1XaeI>QGUgC9aV<6D[BYgE^_AMR;_.df5bY]QgdUO4:<ZR;1FM4
C\.A;95OX3c-eEQ#cLX,2Ta48=:7c?g.A-N&A&YAFVXLR+ecdJ,?310fF3aYaC\4
@9_)NLZB_Q9<U8W.OZR4D-XY:&OO.8(5eD#@+K[JX-O-&_1R.R#UJAP6#&[c.52<
<>0EI;&[8+QNF-9,E:8)Z01-g?;\.#c3YV/PP4K\9M1@LW6;&R0/M\3+dGa)e)A(
ML@BEE^T4099S[fF]fBWEJ([E589P-R>=GeK2HGVX\-Z_PV,@RI\_PY&fJ;F?CH=
@#WL=J3C[S8QH&T1P>MX<<>6JC?--;)gJ7,BAV=^D.,DRA>:D_(-]e\f=D+H,&D=
8>W6U@&Q;SVO0[KfM3(S0g/#IW[:B5=/-faMNMKD1^6f:]=\6E[c/(>58Fa[2G\-
1-\ae5DTZ7=a.J5J:Y//Z1AQaX096c??\PP#O-177V/BJDX)eKIJGHHP)C_dIYM/
bCWTJ\D4C:N?P:dXE&@@9Z0VBZL@@G]f]9+P;ag(8)XQF1PCOHU679=C#0+PWU(B
DG?6LXca6PI(M]aUeN#:>5bb1&/e<+A.0BVW2JOM0^>&Cd+D9./(CTeADQELHJSI
de5ON-KXPC@.U[aN41JP_HS/e;&NAe?A-Me>_1[c]C6UgB<[N/D/1dKMTdb(fbaZ
.KTW(&S52,LW[@<gbVP^5@B:QX03-_Z7;]3>I/)\KC0,WB11VY4X29HS\MQ0a)3\
@f0QeABQc,B:AU<5.2?e-TVA;KX>=J.U#H)aRUfbB4Q5[H#JN2C]A6G:fS\WU#Vf
_NNe?#;I[NccVFD6fd6=PB?>bd74<76--AE:=F]J<Wa0WQB7+Fb6FQ&/c41HN,P?
T]S@b=KQ[Mf@fTJe)a/[gJ)W.8#Y/b7F^K5gd])6K<aY-2c64GE0L-E0\Z4Y=PT+
b?Z:e6N^e;FESEJ5QbXUZA&-M5_:++O<bL^951:-;K[,(Y>1J#)2GXM:QT>EFL=&
OgLR-YMcG#G@SQ+eY\O=Q03?:dHZ/_dDGe162(6\+:I>+JRdRDe;D\7K,[#IN],)
K]5:(4KZ>U+MJ.6:I(&&5PC)g1Ib&V>g+<>f5e-<;5+5H4Y3B])H\H\5X^TJD/Ig
_AD6@IdUJfKNU##)?>RCO4:Ug.611+dGI0Q&>U,Y4S3QLN-:e+0.K<VB&58b@9)Y
0aS3./[DZRPV=]G(K)=LXCTQ^VBFDN[94R<AZ5Rd]a71GQf3AdBQ1G[BG4R<YR9Q
::M9La@N+6OX_H3a)\5;gf+B4-)]b<CQJEIE;8Z6P?N()U,E_7,b\SVNH45aPI?E
:8NS2+CWY9Z4BM:&3TUHAb@gd-]DFL4SeTH<L/OZ__];[2K7Fa_F>5M8D20Pa9V#
5YO8?ZZ09=Dd6YHgKTK-7ZJ2MMOV#[-68U=bcf_ZDb;GKR#B:D689WQGL(;[)Gg5
/T6a1+>/(H96@PNEJ.,;cc3\fFb_[J+.:$
`endprotected


//opening this macro for dvt support
`define SVT_AHB_BUS_MON_MP_CB_SIGNAL(signal_name) \
   ahb_if_bus_mon_mp.ahb_monitor_cb.signal_name``_bus
     
`protected
I[F1H=/,+KQ2M<YM#T7\7IB]GC4[U4V;NBIJBW5NKBE4U<EHeZ+f&)IAbC4P27T&
I=5-SS5dQN0XJC2YeW1<-7P_Z.+2\5R.5eY)OgXP8Z[UP1TcaM1cHY@5c9)2TG#<
]d0fLD;=H)B8,-4SeaDGH&5(MeNNI;_>Vd)bDdO>0Pe]CR7[U&Y=+H3[A7XZDF(0
;(E)1D,;B)<R]<J\HK1VIgMcFea?BW(.HPUKCZ-bIG2;_fO(SY/bBKg3>]bK5-df
M5)^/EJ2G\d[O8)-T\W#MIA<.4EST7&UCMHYL<TAK)A[^=d-)HfQ5Cb#c8c/-Z;R
Q1M[BQS-7e6E-b_CI81[J]a\OSV&]?;d[S#9#7bU3J)WIZ_]fVgD9[?1.T<J6063
)]#G,>ag:+5AeZ2YP?NgY[+S.Tg>WKg^)aaTA/A8NY]]8&N.4+aNX7M8J?0f(^8;
M3g,?FD/>gS[7<[,1>>94e]RH?9V,4.:1:3;N:@T-Eeb^6OfU7?#8[Zb/D3F:2#d
X?_M)OEHZ>#Z3>A,5OB;.W&BV^UK5N.Re(48N&8gWG]JLg#]9cY#R;:cHO0f04(_
A_<:+2SSfDD8+Wf4,3YO61g+[;cLNHUK\&+JLVeKPgDEdIac&,S8/C>+QK>;1Da^
FKVFF5+N/cB-bcJ_N[\IF4S/9IA)P2;E0C8dKa<#;&9PeZVFONg^#NB2EL+aC>B#
,((YP]bOB@.CGeKY+0S]]aP>g.U/)^ZUfgF_=8JZM87G,UA\?[-B91@#5Pa15=>[
JHfA+M?RcKD.&VQ=?3B&]Q:OPUPL#B5^A,=AL;4(2V<M5_<RB>NT&.)&2P?Z3d,M
S^)Wbe;-N&8AV_#YH-X\)QgHb^(HeTb,Z.ET,0X&gXETg.e?+c++Y&)>)K3G@N?E
IFT^T/0UOP^<;L_5e_R,#W;K,MO8/g7@O(HRI,/_RZ&?X5SW&W,(OHC2&ZQ[02OR
gADRIFO-MbS0]5e.1B3TX&EN1-,K].,0+A5VMNdd<7W;9^Y3/CHd^PJOFSJ1:+#+
0b7VLC,FDdP6I?W3U]?GE6[fbb[aH:8eZ/3&F991\C7-=2J2BKE+N-EO[MNQ((6@
8RZ9C7OO_:@cT?&XV#5QQ?V0Z8g-?)8Q2M\aGLbMW_M-YeQ(DWVa;)I+Y_G35>Hb
W-OI08=.1A\OeLH#4Y4b9eaO0P/W&W8Q^LC.GPWR5CG)8Y3[UUN\KX3]OJTU7]QX
E#UCHA6LXE2R==2.W:D49NOF@DN6aLbA82@NH>DbI/H5G.ba&760TBA)ET9^?.RN
BM96ZL)@LV6UD&E(=]G6:KR>d^?EZ5S6TO[g=@7(TI+@/S=QKRLP]ACC<ENMXcGK
<d\V4ag4OPd&?<L06LPR3eYTd0_J+[>=IX&Xf8,OeOdJVZ(&1Q,NS&2^>[BO1EbI
JB0.A2d<EG?3AR)MF@R0AY;3S#X/dWGJS^(7UJ,OeL780\#^eAC<0\6)O<Z=6cbN
2>2_1P8(CPK)dG8OVfgJ/N[DTJ,AGJbYN@Rg5&/;RP[.Zgd:.cT+Q(<;2\M^WR<,
5:dKV2Aa0F@21?.^B/W8^b,aKG<[KQQ0gbK?Q;N_BXb6(M>fNC3L^c\\\N-7,BaS
-[gg,UZ8#[OWd4;,07IW4a7QAReK>W5f8_#)?8gfPM_K9Xa_HN?6^L8S8g/=+@8a
[@K-dQT7631,O(8D]PDX;N,IR+0A)TIJD(=IPM2J);)P;RJF<fH91<^IK-]ZN+TH
0cN87QQP=ZJf5XNTV@UZ]<-a#ARB1B.9M5KL8M46)f2Q?D5,I5,@IE,MJW(<UP_d
M&STQU^8g4a/Fc=GBe=b80(V6/e#6+f0?A1J9d_Rg-U5;>+9d#3O+Cg,VCbW?JSX
F+PL@9&)@2d@,R.)=fWG.X]]AKU8+4?]UOEM6N5^DUJR9IPaaZ/U)Me?B>7LH^cf
#D^X?ZB=H@=^PeR4cA?C@(@[H<Q/BZ,]dXL45?JDV0B?gKf/D80CW2aG16^/#:?-
(_Y;>AK6#Cd]57EEM++H7OORa,B4?HU[gKaZ_O@Ff-FE(]0R\6H85eFaUA@RT3C?
T\/IW59_VLXE[UbTYQ+D5,0V1/=TTf0.gE,64c;G4JS?@S&ZK4_2<CM7XTB;GKB(
EJ^@3>@6eT6]#2&)60V46b3f095_CD\_)e:#Z[-A#O0)>d.NLFWg)a-=#.>P[/>\
(1VcFUNNb05D\&[79TH&LbO2b87<5G&M^Rb0VBSM,WIMe8eYHA6E8O@\Ea&=7^\G
[91LT4H=QR&7Sc;Db-&<:51@\Q^[@D[DX\a+(.\(F;6/PKBee&5:BO>g+Ga.;f<S
[a89#/LJfG:PVE]=_QNJ-@cHaaSK>0F][\Qf3P6]IL:L\:(#dPZ7#g_FJ+YXK]<^
7HQf-L,]d,9<g:9LB#KJMGO8&b\g[L6T28GFL#XP,YN9.J#00QI1cDWBC:)=9NH\
8X0_JJ);8GJP-e+WgP00CaVFVbf6F[#/P70++?Z0Uf#S-O]AT[:/:II;TNWbfEI[
X+f)>R4+>6cQEJWK#=XcJbBFNM5(O/8OOP7,fGUH8P3C:Y#9.#HK@EEL]VBCD5N(
\C7[GO.+?<;De;:\WJJRM\ABHaIVMVD([68K9PD[<C5#,S+XD49S#d?eYHa-&3G\
C1I+H@J3d)MFDYA^D/>+@:;dSNA5V;Q)5#BQ,6@+Z]SU/Q=Dd.;(&]g^2K7f9ZId
3baE4GL9gb^L7XY7)^8U7L0)OYgQIVZL\9#39FdLEXDFSCgbQYFY)e<)C0M(O7)X
J6g2-=6MS[O(NHb4J#UC1_]U486b&91T<aHC:@K7?LFOJ:PR/ML&fe<2#RW&4>D8
MYQ:d-IZ7?]5O9X@da)_7/a53EfPVSc/:8##1+10Ng-Y6W71X8.K1:bX&>NMSIVJ
BaV^RR3a&NK6R(RDfaJO4:cJ6GHUP0;E]0P766\H.@)eFBVXD/D_3R_W:GED]#Qa
5L\GG103Ue.@O@/<+Fa,Kd-+Z8:b]HP:FR9AEYbb2ST.CEWDc&#]Y\gEWJ-b6O>,
g#_5JD[@Oe<1F\@CJS7]RVXDZVJR(N^00Og><ZcM;#AC6SN>d0NgHQ#9bdYef#c0
<:De36>OK[W10$
`endprotected

  
/** @cond PRIVATE */
  
class svt_ahb_arbiter_common;

`ifndef __SVDOC__
  typedef virtual svt_ahb_if.svt_ahb_bus_modport AHB_IF_BUS_MP;
  typedef virtual svt_ahb_if.svt_ahb_debug_modport AHB_IF_BUS_DBG_MP;
  typedef virtual svt_ahb_if.svt_ahb_monitor_modport AHB_IF_BUS_MON_MP;
  typedef virtual svt_ahb_master_if.svt_ahb_bus_modport AHB_MASTER_IF_BUS_MP;
  typedef virtual svt_ahb_slave_if.svt_ahb_bus_modport AHB_SLAVE_IF_BUS_MP;
  protected AHB_IF_BUS_MP ahb_if_bus_mp;
  protected AHB_IF_BUS_DBG_MP ahb_if_bus_dbg_mp;
  protected AHB_IF_BUS_MON_MP ahb_if_bus_mon_mp;
  protected AHB_MASTER_IF_BUS_MP master_if_bus_mp[*];
  protected AHB_SLAVE_IF_BUS_MP slave_if_bus_mp[*];
`endif  
  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  svt_ahb_arbiter arbiter;
  

  /** Report/log object */
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_log log;
`else
  protected `SVT_XVM(report_object) reporter; 
`endif

 /** Handle to the checker class */
//  svt_ahb_checker checks;

 // ****************************************************************************
 // Protected Data Properties
 // ****************************************************************************

 /** VMM Notify Object passed from the driver */ 
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_notify notify;
`endif

  /**
   * Flag which indicats that the address phase is active.
   */
  protected bit address_phase_active = 0;

  /**
   * Flag which indicats that the data phase is active.
   */
  protected bit data_phase_active;

  /** Event that is triggered when the reset event is detected */
  protected event reset_asserted;
  
  /** Flag that indicates that a reset condition is currently asserted. */
  protected bit reset_active = 1;

  /** Flag that indicates that at least one reset event has been observed. */
  protected bit first_reset_observed = 0;

`protected
8[M.HMg44e8D:TDQK:^_.If>&IQJa0F&]Ha6K00bP2EJ#B1g[fV_))aCDA29D8S6
(bSX,TZ\#<YD,$
`endprotected
  
  /** Flag that indicates that the dummy master is granted */
  protected bit dummy_master_granted = 0;

`protected
]HeBFMNZ;;&53>c=W7,H38DKPIWXgHFOJc_ZX3.EFAFX<ZV/d3g,/)6N6.DS=MS/
1eVE9.29+1#5,$
`endprotected
  
  /** Flag that indicates that the default master is granted */
  protected bit default_master_granted = 0;

`protected
TZPXT_,:PR7349[9OT5b_;CSb5fKG#VXEG\4L1B_?8cIaZV-LgE-1)020\[>1W/Y
>9)8T?_K#cD3,$
`endprotected
  
  /** Holds the sampled values of hbusreq from all masters */
  protected bit hbusreq_sampled_value[`SVT_AHB_MAX_NUM_MASTERS];

`protected
X\Y@<F=5HRQ9Cb[QPX&3FZ/K.IIAB_,Ha(#<_=NC_.:H<QKBFS@S-)M>+4=@R>.G
.(=Y=-E3dO=9,$
`endprotected
  
  /** Holds the sampled values of hsplit from all slaves */
`ifdef SVT_AHB_MAX_NUM_SLAVES_0  
  protected bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsplit_sampled_value[1];
`else  
  protected bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsplit_sampled_value[`SVT_AHB_MAX_NUM_SLAVES];
`endif  

`protected
O@3@&A@]Z.Hc@.ZINI#I]6TF=1d1@TFUa)Q)-A(/Q#E_<S36UfKK()&@P>J7/_Ya
gUdQf=eOV2Yc,$
`endprotected
  
  /** Holds OR'ed value of hsplit from all slaves */
  protected bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] consolidated_hsplit_sampled_value;
  
`protected
R0V&??8;LMUeg2dc+:][^eTdK/O_cTD#0,YB4:P3+3.KR4KB3;?/3)U.C3gbKfdN
,Sc<V9-+@=Ne,$
`endprotected
  
  /** Holds if a given master has an active split pending so that the master can be out of arbitration */
  protected bit is_split_active[`SVT_AHB_MAX_NUM_MASTERS];

  /** Holds the expired count of the cycles before EBT event for a given master */
  protected int num_expired_ebt_cycles[`SVT_AHB_MAX_NUM_MASTERS];

  /** Holds if a given master has the grant maksed due to an EBT event so that the master needs to be out of arbitration */
  protected bit is_mask_grant_active[`SVT_AHB_MAX_NUM_MASTERS];

  /** Event that indicates that tracking of hsplit from all slaves is done before the arbitration */
  protected event hsplit_tracking_done;
 
  /** Bit that identifies if the transaction is a locked transaction */
  protected bit identified_lock_transaction =0;

  /** Bit that makes sure that dummy master is granted the bus after
   * SPLIT response to locked transaction is seen
   * locked SPLIT. 
   */
  protected bit give_grant_to_dummy_master =0;

  /** Stores the master number performing locked transfer */ 
  protected int master_pending_lock_transfer;

`protected
GU=RZQJ@/CGAM,-)N68e^77>5]IaXfZNE,cL2fbHQL<cdPg>b)6@();3;YIANVXP
,=YK<MIV3U:A,$
`endprotected
  
   /** Indicates if currently granted master driven addr, ctrl info is valid*/
  protected bit granted_master_addr_ctrl_info_valid = 1;

  /** Flag to control the muxing of addr, ctrl info */
  protected bit continue_addr_ctrl_muxing = 0;

  /** Flag to control the muxing of write data */
  protected bit continue_write_data_muxing = 0;

  /** Flag that indicates that bus master is identified */
  protected bit identified_bus_master = 0;

  /** Event that is triggered when the posedge of hclk is detected */
  protected event clock_edge_detected;

 // ****************************************************************************
 // Local Data Properties
 // ****************************************************************************
  /** Configuration */
  local svt_ahb_bus_configuration bus_cfg;

  /** BUS info */
  svt_ahb_bus_status bus_status;
  
  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_ahb_bus_configuration cfg, svt_ahb_arbiter arbiter, svt_ahb_bus_status bus_status);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param reporter report object used for messaging
   */
  extern function new (svt_ahb_bus_configuration cfg, `SVT_XVM(report_object) reporter, svt_ahb_arbiter arbiter, svt_ahb_bus_status bus_status);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Monitor the reset signal */
  extern virtual task sample_common_phase_signals();

  /**
   * Method that is called when reset is detected to allow components to clean up
   * internal flags.
   */
  extern virtual task update_on_reset();

  /** Triggers an event when the clock edge is detected */
  extern virtual task synchronize_to_hclk();

  /** Method that implements dummy master functionality */
  extern virtual task grant_dummy_master();
   
  /** Method that resets bus info */
  extern virtual task reset_bus_status();
  
  /** Initializes signals to default values */
  extern virtual task initialize_signals();

  /** Drive default values to control signals */
  extern virtual task drive_default_control_values();

  /** Identify next bus master */
  extern virtual task identify_bus_master();

  /** Track hsplit from the slaves */
  extern virtual task track_hsplit_from_slaves();
  
  /** Check validity of address, control info from granted master */
  extern virtual task check_validity_of_addr_ctrl_info();

  /** Pass on address, control info from granted master to all slaves */
  extern virtual task multiplex_addr_ctrl_info_to_slaves();
    
  /** Pass on write data from previously granted master to all slaves */
  extern virtual task multiplex_write_data_to_slaves();

  /** Drive default values to data signals */
  extern virtual task drive_default_data_values();

  /** Drive write data to all slaves */
  extern virtual task drive_write_data(logic [1023:0] write_data);  
  
  /** Wait to identify next bus master */
  extern virtual task wait_to_identify_next_bus_master(bit wait_for_hclk_before_proceeding = 1);

  /** Returns the burst length, burst type */
  extern virtual task get_burst_info(output int burst_length, output svt_ahb_transaction::burst_type_enum burst_type);

  /** Tracks the num_mask_grant_cycles_after_ebt for the master that received EBT */
  extern virtual task track_mask_grant_cycles(int master_id);
  
endclass


//----------------------------------------------------------------------------

`protected
(J@VOMMaH.c^a.LX^M0Kg1_1GD7?5JgRTSX2Q-Fb-UgP1W@UI(_Q-),1&>R96aZ0
)CBL27_QI2aVfgbDZ0Pb=+JEMAf3e6aHc]b^&=80IUYaRUHaZ\X159a^/,FZ#-6P
a/7.UVb2&+J<)F/SX_#H(T.QNJB-3]MN/S]Y^,@)Wd4P;BKY+2VYO\[LUT01\[Da
4OS=#PId&c=(\#YAdO@BG>gPBQN:Q&&4I&\7Z;+N&4HDd3IVNGWd/X-Hg9O3YSc_
A-6Bd>C]11gIg&2;8::NWKZ99;7Tbb-Qf\=ZQ5X&c8[:1\9H7OZ4+01W?M,E[\L)
?U1d]d?a[?&K#SYL07G@]#=f6d=5E[bW;Y5&+2LC58N>bY.>BU;dA;8GV,<-IR;W
);c<-4LWYaeAR]4,NccZKOgK;Bd(@H39Q8XB1940N]Q8=caW>66=XDNW[D?P&0Te
10EH9-Va?KLTGaVN5/cbNS)=-7KE5JGd+1>F9_6CMN0e9;^TQC(dGW]ZWe>YX1YZ
eX=BKe/DASH]TC8.5,,T:JJR\KE.9&5AV@\bH]Vc3K^fD?g(OUQT8>0]aEC5KJC2
,AT4B31.UXIdNO>P\2dE./R7)R._YgB@:JZ8VT5&;,C(bKKQb8CM8)E.&f;:L#f6
GAf#I+WO;b4?,CCHA&\A-<?5CH?f3(PXgN4=,NX]\2eOR.W.=Pg1+<df05:4@,Oe
8N,(-fL(I57_#RMZ)[Z#/Z)8.6#<=<fU<$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
Kf:[U:f1YMX.Y4HKg-3,[K&H/KYFB1?JS:U3LJMeWRFG59&d_J4?4(4\ag:g>+^(
/HMb4_SC-eRgJ6(-L#&NC)(AOY883SCHVT0JWNG0]XB2XA41aH/#9S[Cb6Wc=]EH
c&O5OaI+Q\O>Mb8dJ728<@RU<cY3&bVUKQ+&Bd-a_N9.#:I/\9[+P;65ebFA;91,
H/9W/<JD(3I.7DcF9:;ERF2b.Y:@__;[V;\<ZZZ5>=DI^Xa]^:</-=/dH(GD/,2?
)S=BX,VUa1DC=R3I[b3&g=VAZP\:[KBfB[XdfK0A+gVDCVSSC#:24/#9Ga,Ua1b?
5@DO9W)<DK6:C(N2M2N;H;65G.YfJ,.(/cCQ+Y/(VA:N:(e-,8Q+@/?44[@e+fHF
&P#=W/9c?J@\EA:^>158XbTaS.1dJ-QSE>9&YY,;_Ec;:@=89K;G_&O=JegF#d/?
UbP?0.QXE0d]O,P1\SdLb885(X&[KM)cI]/dcSQ>WJMg=AD_dfBQ(1T?M8/8[9J>
2EO=_AQNF2_=B@TC<eS>:F#e?B>Q=ABT(N9BTTa>?+f1RKILP.#@6]S6<0W2a/4D
AeUTVIW2]IB56DWNK;ONa.(\VW66,#<ae?-:BT:aOC8&dE99L0]=3NCBQ<TIO(5F
N9X#>PZ]+IUEY9GZYTN7&^M6_7Z>+B#.[7_@J]M8SU#Qe_Tfg(Qb7)A_U7:=W6C+
a/OfIYL9@8_)/S#RR]A>UW\aK@U_4MR-3a<R=_3-cSTZe1J&H/[>;B^BBKOU;cH#
MG-#8^(ba8.]b5IJcI8-aYD,O8cCgKE7W5-V[\+#Z/+KKNfPVSE0:^HGbZ<\&^#<
ZfNG0CUY[IfHc7K(9[70KLH7B6GQd,8Q3b&B8\130PKX0/R26f?2Ug@#3g4=&TX9
&.,U.73:P:]3MKce:J[)Wc;5:1,)0)P]:b(./B+AKZ\^d69bfKXBfd1Pde>gX2AR
7NG#J0?FJ>^R/_6L.MFeR&/Q6ZKdF4_P+V_0GHe2;5We)b94R(aa8[eIH&8@QUT-
+8+7P=<7=Q_Gb)W/&G-./S.dT629C@/F4RIHL5?,A,c>?;HcMO+^E3=J95gZFe8P
a?NXK_R;c]>+GAcPg#NA?4bWVIfNd4:1K+f#7<EMAQM:UI]7CcJP>K=>X0&,e@E0
:/&Kbb:/1cBS.XR(\CV9K9.HRT]8BPDUV1(DP6&RLcF@0=F:gV0ab-4X/RUc<GXd
O9M/_9V0B8#F5:5-ARZ?@J^TMKRXa0U8&_Mba>bcPK@:a[8,])PSV4RB3+9UT10g
?^YQ5C+JS=XS(KLU/+d1@CNU:[-:cd-Q_HV&9Zc&4fYD>0_fa1[Wg5/V/,8GPBg=
SZ\S@W]>+:a2@9,M(6AdWGLJHSI_,8ELF=YZXCaHL@](L+L8OBL@QMZYf>1=)aNY
aC=O74aP),+<IAM95V),@UX/I?ec:::aJQ(FU.XR:-NK6bB&Z&ZOIV&T1/Y4)VR2
#=WQ3<&/EUD2f)#2S6R?M]\341d?JGZBe#9gD-#^[Og_A:.8D^OB]U1e/#43WO#G
Q]_=.8P5&-QE-C[[F+/32#\])KC?W>;LdV@\-/OUZfX6Xa]FXJ7G<2HVTXRN71I=
E5cV]@]69T3O<0Md]):7ag]>B.P^-A.TBED(I2^@CZ1[\SMQ[39AR;GC^,>8-g1b
N)-0><YL(LZ/Pag1B(OIeE2R([R2N4@b3H07A>FF,(0-M+PG3J^ZOBBaaK9F-].8
[S#<G6/;-5P]>?T,]?aGRd:),+Y#BLB8,8ZIe_IUS?@@QJe0JH^g?@&6a4c9Ia.Y
UI]N=D+3)e#7_0B.U@c)7TX_gba,KQf/5Y.D+7X)65dfA9JSX]4C&-@W8MLV;bcJ
A)@dUAV<MeV@<,1\#1B,?4bgZ?:3NZ=?aeJYZ\4-a@X62AZNHB(5B:1YLUg9\^V6
3gY)g.1>fS67(;DbfeO<b4Ze@(--^bS]EXQ,OD65/\C+g,B+:VO@f:J^BH4OG;&M
ABSK^a?[I+=##QN.<\-JD>/VKH19IGSJ3VW&cDU&N@097#QR#_^&F_CTANSI?P;Q
T0VYDH1gS6aS#ZZ;=FVfT(-4>NS#8U/eDe68-]DEcOf#EN7-5?P=\?NbY8;-3Z18
S+D/QYHEGOQ]7^\WO,#Se@RT_06WZ/Z]AOOYb2+(HLd7EP[WLP(0dQPdT\UHH^K:
0Y?0&.60H+Q&a]0V,^:8HG,IDDM30b91Cf+gUVQXG<I[&N,\QI&OWM78IW6#Ag5V
-V3;>g=;IYJ-,HL?M6BdE>(-^Y+UJ\8)?F8OBY/6W0c2.GEbL/O.9_K)Oc0d6Vda
T171feL?07XRf9SLI^RJ.N&,.;D21[H594VU27[NcYcZ575dON[X?.4.RW^c9bfU
5M4L;>2GBccXY.eGO/8[aIHJgd,JU3/AH=68M33JE+TbQ86YFgDGg5BCOF<<PZX)
0#P=+?\4=<7H(ITFX0RbW;VT1&D+gD7PXL^R:)L=:&Mb0?bYJS5(H.6OOW)_BQ\Z
T-]TaOP,UgAGJ51F<^S]2S++N47]J6.IG^6/5&KNOb97/42dYLeEY44,aH=>]B]Q
L^EbX(.HZHZ>]W#A-TRZ^bDC([\KXX71(b2/AYGN9];;#[;@_GNH80g9OD+Ng7V(
WYL<QgE]f2]XFYI[HAHFa-VC0I=@1TaLAK@5,;9Oc8[:TQPeG<L<PgYD;O/?\)cC
U0R-AM(ZE=M..T81?[e7G>9-1UaY]O^27U][-Dc[[+S9AW7c6P<_O(#46<e1QECS
R>^=gf4/dUDG81K,75^B.S^=2Ggb)./VdBYd8#cW65KKP6Xf&Q[<I^bZ92g6.NYD
?\\V9XbXOd<Z\I(FT#33+)@IT120Wg22^9Y1/02d6LN\#PL)0(=GW\f=ffNSBY;7
dPAIa?TaL<MS;3_1\NdXc7[ZSSQ64@W@Zc)?HZBG>aW89)gF_Hg8A+DTR(c<cD?F
N9-NGQ(1B_/1OHD/b&ZU\6,KBSJA<Fb7SJ^RZKL7M&cC8RE)aee9A6=0@9)[V^Ad
<WbWH9<K_C@-\\g5NUGTGC2LQT:A&@dAO@4@c\04??G+N]I3?3Q31L&\@>3SdL\T
]1K0X2J6:1Z>_]Q00WP#T]cB=0[LFS]0ff7JIFR[2#bf1<=;OMd::<JV]EXb^aA5
KPb^@L^&HKGMMJd&E7NLIX10@?/Q9+@ESBN-BCc-A9U@CaV(?N2+K71W/3/S.c-D
DgQ:-04C6><,ZO0,WcBfL(/Y#.@6A51^FFN6,bVQ2HUb(LRI#J(OEE]eC],HW8BA
VN6J#gW>g3^H6_44+D,6XI:[JE3+\69b?]c3#D]3Z#E0aJBCIB#X2+)S?gda+TKQ
d)AY.dX];F2),TV<2eH77+K8T+T+d<#KY6dWb8b:#.aUP[MPcKT>1NF5,(Q.9:47
<#0(X;McDM@C8LRL3=<5@/ZdUD&1V.ESMAD-UPLg-Q46E5#RVXLg4(,]H:&_4ZFa
)XaWVaDT>gBXe2d\BMfF(ef)dK0;e0]U&\D+/+^SV@L[2[AgTR,Xg.:RE5g6a3ZE
fdY;I<&cT/PG)AGF.N/_PB94^^E(\TG.OP&1K8Z^Eb+&X7ZQ5E+6@S@G-ENB3.@e
bSFYgK:a^b3>a&H&e?.0F-<cS-QG3YH((O9U(N6W[TBGa0,#Vg3gfWFU&03G\YOB
[:.>\/bNY,:Z0-Qf?d<Ac^\N+O,K.bUIO((]V4-=P0O=#O.[)/GWJZA?NJ/dDY2N
EC7a7b3)eB+eSWZ8[\a7LP0B=)HQ/5_T<>995H5g\NZL\VKBIN)+e8e\X)9(8OK+
;6^f[]IK3Fd;<1TCb/SX-WB?,@c>CMJCa?PY;ZFf#5-C,M\[L.]D])-<&.SG)5H&
M48b8ZD,[K=+#cO@U+A_TM6&b-bPY)FcRNZ)1Ye]T]LeA:?@FRV@46LC.PVa^7&f
HLH:F<^eV4+T84_dKL;:^J+OJZ&#0E]5H;<9[f#<O2HMBdfRO[4MDe5egEMKD7_D
e&6X2aLDC7:\U^RDg1SYG_C0B32aZHf3KBF^)ADNJ-e/(_8RZ7EO8Bc::V)S&G4Z
.26addQPJI\E.Ef8R:X&IHZU5(U@:Y@.XZQHVU)]H[].[G0VL.Td1deK=T-Z6^S(
T56SAdJ(Z2&(5Wg(.?XEJRZI]6L(Y3GTG-&.+#WLeCg3RZ_Mc=:E6O\N^b4b6RI]
@8#EGM5]5](_(U7LJbR_#]?M6A<03C3T01<:BU&5Lbf?X;aQ;YPL>(UD,.SI+7=E
J]BPTZ,39>?eZ65M@/;A]>BWG8BW?]T<=])@4GV9UP=HeXV.Q1Q57A-QO>/Z_^HC
P32/e?+-D6],[IEOYZ-B7@Cd6B-NQa_Q^5K0dPF<7IBFE0Jb6T+5Y,6I^B-cA>4U
=A5]&^M,.IG:^KcQI/;=.J#HVaTd.K<<WAZW<C+YIZG#>JIM58=,)d<g(Q7<==Oc
N03TYSMEC8Fd3:(f=C>?,4_eNPag++C[FAM:/=3g>-?=\;e#2+UZFW,=D=e>\[&f
Q:_+:Y5_9A<[_P<>S+a>cE3<[]PX9FZ6(WE^eC5gAFNW9_T/[_[EF&dQ:bNGV#3,
O5XKY))L0M99SVL/2+-/:);T[ScXgRb+bMD8NgZJ@->dRF//DJ&9\IYBH6F2.MM/
:=A=YdNSMXFIgI-^VPRYC]1NBFKI#55>IFL;cV74K;2RN&fWR>N;R@b77(S)eZE;
:CJP-1cA[H:H)D]gBK;EC_ZfL-fQ,5RS:4G:GFFU)O8F1:(;3>&KHf25LZC[X\^J
0=Ig.A<4.Z3S)JN;FeKE>IL(\?3JdS+QI?[XIA8X7I@]:)14a0ZWGF,Od_;D=TSE
cCD+N9U0<Y+c,3_\b^O<<FL1K/[OI,eSNgB@PXZJYUaOV(c&(G<,N#^,L>?[DRM+
CA?TP7?07;[^X,YHG2>3JB[WH1VYQ/P86E-B/GA.JN4-/F7Z1EdTUFX^\@Z6:e6_
^F:7AX^A8:\A7S6G:;#,(06f]3W:41eM>M4#4Z(dD]Y7S7@YIGYL[G0CT9/81YSG
Tg>.5DUBTLU1cP#F0g1;93EB7>BUc(S_/=/9]Q1OSVO-/eBSB4UFa,fG>0.9IR#O
N]MB1/+;1RDS5=SV)],;H^\KR>W9,D-9TI@+:B23?^55b07+-6TE[J:(Nc6>(NKF
;J<4H@NCEfAX.<4&+AR.#C\6A:JD@&UQ[BYa]9UQ>)^OB^Y4c/GZPS\gTbN]F_N5
e)=ZU=e9+>3?.97#WbOD;7;MU=g=b[d@1fI@aMH5:.6VN]?0?7#U,II3D5E80W#Y
fJYGX[9AWbIc3SI0IHbO(5BYKR?bEJW7)^TfdNO0V5ePScb734#>+aKG5&bJXU(A
Kd16.Yf9+24AIL2.L9S<+GNJeHQIQ+#D]P@N4QQ@]\#6G94W;S5)90G\G]@6R(=6
XPcL/XT?b2+I=YOGI#]&A+Lc>EA(3)BGd,eRZ7?6>c30WWIOP8EJ-23Me?0+=F4H
,#bcL1[&\+;a&??J3CJ70[-@C.a6cebB]T6.7N2GYD4c]OPYZ=4c=FA7&d<R1YDR
XSc9I8;J(3CHKgW-M7FM_?.a&X/B+LGH17^6EY??GXS4--Qbd=H(W@H.M.G\7dd#
^D?8VW2Z:J/=FM#Q)(LG7cI0,1bHWc&>JY:-6PTeK3)AH,(5[],3XeKO[_&3:eLH
dT215/321E7?+eK^(GIdWXXX==XGDBK5KeTX5^OUXCI4[Ba&\fgZS.&K5Ge10_/G
I:aa4;C=<<,fJQ]R39<44DWZZ,RW@DV?NF;Ye2T)\c0S8aLZg]&@8@H\bYC@GZ@#
1]#IFW0)QM#E1-3ONDBW;D26WWFLWZ-EX>aDM#W[=_&G-RJ^1QF^1(44[X@Baf[&
I6#AcQG)HY:@>YL@B14N&g5OS]6-g&>&MZ/>WKfgDFVe)[M2WE1;ER0Y&8e^N)H\
e:54;O;OVGNKf@T5Be4^,N.?8&QV\L>NNP(:3@YcY57U+;V_a.=-9,]5TIL/cRQ_
[F4(6LG>+cYL5?[ac=aL7f;/De_Xg0RC1&aI&7Wa&TW6_L=P@27a#DaZcZ+[ME_Q
S&bT(WDI^/G9L.+?^OTV#JMYA+V3U>+:YJ0JeS0B<F-M@\.VgXJC\;L5:&6_fWA0
DFg[Z,15&E.K6HM5#g^+S(6gMU^<ff^D_D9FfD7\BaOc,ZaVdc84)fI]Z>dY+2H\
(Ff6Ubd\:=ST-9#gVE)MP4=bA/_IWB8Ee=gg<a]SD\:AML8.(cTM(J4(<=\GNS#9
1P.8\DD:XWS?5?QJFJ/==8=2F7I0Y2aLb^TWMCa7.JdC>EBb@AH77(D>KW,=XX,@
497c3BB3-?<gE[+9b:G82(:)C3T&.IE(5?K0__<dO\dRH.5bP@XNK<VXI:9EK)D)
dV>+OJ^O_EGXMP5Z&f:V/D-&(bJd^g>.+#f1RP]M<007:?g/gJ\BJZ&Wa8VPSOY1
97M0_d/eX_>]S5R],],QNdNDG1VRZ=(&Ze^QbO;2F=.^-&R3^Z<A.CT.>Q-9UBR[
A160B[D5I7.J.2<,S1MfS(C=K41/?O:YdBP>-dS?MBSc_f?Z<#:da]&31P+cD(8T
:DfWTb7289I=.I\DMDf1]7OK94D+0NLLd2RCeXGS2,IM6]HO1984d6B2^V./O9KB
L=\E^cKX(gcNB/d7;UO8e:IF:SHLH-UAZU5-_))K6\95ZH6?Z^^:GWYa)9Z4\MLD
PY2W@^,:J\X1<]N0_SLT\]L^<SbH=K\44W=<T96KgGg-efPd0RXRSJWB>-]a;N<1
HY5g#:&S]2#@TC4-1</b/]1OR;#-8Ofg>O_A-&b&?W1UM#IM5>ea7&b/cU^e&66G
b-4T\WZF_N9dZV][g9=KZ:UA>\ggI9bCSNI:^LK,]P>?IK1E6U6Z(T?2[1]SUEG]
),g(-#X^FAA\9EcBV+.#_6DM[X?<L=F+19IF30ZaZ[>d&:C:H^/3<ZTA@(P;OK03
PTZ73;#KZ<WMWFQ.@&ga(c)P=+6_6=SBd1Q()R,5KCG;W2&eR,SNFWGCAW.ND+:U
NA_PXOR,88]^MeaK=>]&\\:L9-<H;6\6_Q<e75J.8HZ5VP0B4T3/04I5UdAb#g>b
Sb)&1]YP,V4VMe<6P.VSGMB7=]#Mb.dfN1e(<IC#HVCO@F@&/5BX#U^_Qgb(IG,Q
),PBUcT[AcCW^d#B:CJV&Z)A=MX,GM6gNR8/L0OKMAW,2V;0/<H,K98)0a6aZPWe
&A,JA3D[<\3a^7UV+>LB;.@QAA3[be0/R2SFWZWJ@@HDW/8,@;#bRTHU-,5AF;Lf
AG4KKA1)Kc]LaLTGU[F)I:B;A+4Y:3_B?#.4e[^Y,VKT-,1X)d)\Lcd1U@NA5FS)
?QecQ:=EGW66d]gY\e\.^@gEDBXP5:@/e<0@U,41=/G;78]\84>RAWPCA@/fO<&\
T(L,FR@\\K0E<a5>ecRFE3b01-Mb)()&?\:F8K;;C;>\06dCPOO=,#B#J[+M<6@6
9.9#9I4S,JYQ&@N&3L##UK+2T2&1125gY?21DZ]8I2-B0[<DA5gSJ&LgXRU2(fN)
-SSSW.Z67fVaW30P1HD,O6a;IG83Y?5X?_V[Y?=B(cUZbEF8Z,)D#YdK-UTKeIN^
cdFa>\aRL,R=2&DMdg^eY;dAT=]aD^g<FWVOT[-K[cHELPZPb6:/d[0V&45<6)c6
;+7a0))aR(c^@)?]c;78S8]<;[,Pa46Ye9V4M(OeV/c2SJ3+fTTZ&.<\@gYQJ8VX
5Q=T[2b,?Z09-=X6X8FG@BGTO<8Z,_4]I^FCKDR;NYHY\eaB8Y[NE;#V1W1Y?<,P
EEFHf\4-YZBe+&EVZ9C0PT-4T/J5J<M&DI&GLXeD+bG97)N5YO</0Hd37NFfe4QU
c?)Z6GDUb=GY-8[0S29:8)X4+:^T\fKYZR@LW>g#+V)e&fJ:BX>_?Q^DROCReD6O
JFWB,M)C@eLLK^BLaNRU--b?<(.KeED4T&;c=B(3PW&K-PY0,JOIZ5=7&2DDMYea
9C[E6YRcSXTa:/)N.PddO=4-7<.Z?X827)WEM?8Z8Y>;^24ZL71K9W1;YBEH]:&d
^cgRJ2a<8bN8VL;@5e+R1TU4<T#g4Qc<L^^Fdc_(=#]6DfQ-?_GLZ+U/;V>aU1O&
.g@Hd11:_@;^EHWRLNJTf0@?VE..=JTW)=A)Ec);,DLad93:\R-J#3:4JPAQSZZ4
B8aR/EfIGJXVe4VF2gP;JFGE^JV-4(N=3JP6F.OJb0g.aARUg::6/I.P/bZJ,Yg#
OZB#KIacP>ZJ5?004R_41_e+.=<J@GWA6FPPWBIHfP;(P5VKB0HDGNU.J9AaNDKa
3/>)#]O1W?T;HL>eIORffED6Vc5BaSK;^T^AV56W\7g.g??YWe@AI]NOfARCfMeJ
V,9P_V4)HKTQ?C/D7G-A#\N;N4eQD+I8?I]Y)#:RR<<CfZfD[].RE-&=ad04ZaY#
<e8^Nb+08Y3GY^DYL8S6LV.XB&2OX0We&BXe2B@a>Me4BW9e@KR>R/TOc]==./\0
C5IcJC01P(X&UL;.cYee(?C>K=4F.QDKf_.[3;,_Z7XMR.[OD-AH37?LKU)^=d8W
C@SY^,AF:+Zg_2B_EXKKHe)\c.DDVH<U#([Bf_Md4CI^9;SU=eJ>XM#D^T1CfW_/
:TZ,b60YcbRSHd2bX&9],]R_;?@EFK/dC=F[W..Hbd:a]&1D;2=:AC01ceLUCN^P
)8@a-<Z@#dN[+./>b4^)73BIOVH+52AQO#ZAaSH@_<NVH:2#eL#B<4&+W?;T]\>K
Z4M?I80K?e&#G<,H_([:OVYLXD4dg>4,9^_68Y)^8UB;_,T)M>(62^:<cY]O:9Y8
e])J2S?&>^b7ZW._-IHH@W8AO]G-SI_[89-\+G@XQY]N@Z51aFR,NSCIRKOUZQHM
>J(.aT_;C36g;RI6(D8A3KN2#DA:C9+JU/79O[-SJfgZ,XUIedAJQb-6=3/\cNMJ
CJKM/1Dc+</a>X;8X8WOFHb:,[/\f,C8)2K./d8D]0b3aPY:MJZ&/#]+eVC\e\_&
AQ<L.<;f-&4F^cgN+\L+fgIOeA0G[WK5&X1>J-VYX5W90N\/_cMebP-Q/5BAVREc
0NL<#U\7@.Ca5<7YXGXW,__V<QLbH2C2X++_DQg&?/2Z5R@_RG\bd?g\YL/RID[(
gA]QVAY(/TE(U8K:UYA?XP,=G-+aZZ)2C0)b4[ae;g,7MQMa;0<S:]d:=OU8Qf3\
R#Pf4QOS&NOYbW)SYf4<J@/Y\Lg[?<^5=/J(./6)?96<D.>IQeC/S6^+#OM:DSYb
&L)??02DWa89+<#1K9E@@3OGKTV1CbH\L8YG>QEVKV@M--?)Nb=C5&Q@AcR7ALV[
.A>Xb0@+_1Fb<=de:-g+6LdQfL9-E_JN8MJXI/3:Q9)ebe03B;_2/2C#9^OUfA8f
1-DcSSc<?0G^N=,.dH5OZ,.5dCRTB#D,[D39MUA<ZXMZ5(>:+18IOFLHZ_V+=J]:
JT(;B5@?R/dfc&[V.d-,0?@E]CdIDO6C]Xb7CM<HI[b9-c5QXQD&c)J][9G+RaNL
1?ZfQ(ERAGF[8g29Sb8WO?9M0_;QF(-V81VPJKaO[gJ:J)VfdJ;]3;#+IE](?G7C
\4?31=eeA1##7)(XPbIC5KHK@.>2R55/fVUQJ+G@_;-J9+?e&bDMX<NM<1A;.N8<
O(I93YE#/e<DMc8SQ@BL30S(<c.f?T;KO0,F7,5V>DEaBRP,CH0;:@0WOeUI&K8W
V7)Od9UZ358@@79?ePLMB]c6^:8_9eN]];?+AdgG/g/9I+a5P9Z#@\^VGId7^]K@
aGbUVcUV]HMR=>&1a1;/;Le/1.B4IUUfL(eVAg/?H.FA(:+K2GUC,/8B6OHY6:L,
6,DH_ZGKUE8:>\@T&1+3H+^R)1bW-D5),89=5#G0SS].TP=fRQ-WJH=@XLU@_DaF
Q2^_7M(:dBU^+gW3C3=^g^G^1[HF6?7f[6f;QKKFQ_d9YX-L+4/(Q9_A.#Y^4IJG
Ca[U<7.c=RLVTK_)Q@:D_DQ.4IUCER<F9UKWWW=3.ARVO18S-3g;45Q4^/O-2..V
B>dW_-(/)B^FWd.MX]BCT:9fMFJTA)??2.Z:\e+?1C-;gD9XbIM[YO0SYDANZAED
GT(0E;G<?)V8OEL&^<IMe\8MZKE<V8A@e?8N(725&.#7g.H.))1f<_I>BgJ_:8Xd
)[3gI&9cOYYKBfa&QZV(K8H]MY=\@LS1FM<-;,<SL\]M?UBR)V0&C,C5a>@]RY+0
5N;?YPIW9)C.DIQfb9/HF9BQ4R7GXI9X4G@(R9^Ga7f6<;0R[DOWF?,?7J)Q[OKC
F?JB,PZE,+1]bfZ35Q:1YEbf3.,[<;b.5W/gVW-8(UdefAfPd8R0_R1LK;TW)5&=
S6d&_RVKI#dgI.VGP)24Zg,25eGL.JIRcdP2;F8JSaNA]-c04;:_Pbd59CUFPaRO
8X7U@C\fVD7_#J;9F>Ed00f8<.fFZG)b3R8YD^AFf.@3EQSHbU1YYg)CVTWFBPF9
c9cVRPRIf<JZTgFRZ\[UY\OVX)MI#]##fIK?8B7W48d\1eXdE]Yf_<4dD:g\9\8#
;W_MUWKgc;XLQ9@aZfC\JeTb+;6^GG\[RLY2F;_1/1CC@Sdd2#/XDa9T==>WM8ZU
/TG]Z-X\bO?aU97E2ZV6TVI/W^#4X)RFIASSJbJ]WJ?3,e]H\@af882Q,SdUK@2G
[_)]E6+]Q=\=M(PR-&c/77DJ9a9GPXAGeH3>A]/_/PQ859>:A\&;Wc&S2A(e(e@G
E>Yg]8IUEd8^STVP(Wf6L4-b,(+aICDXIHDG+L0gf.B]>/9WZ-.6&A?3dEQ6#7f,
:N#^D&/45PM&E9-V)NU&b@<<O/]H[[(D6Y3(M0Dc#^E+dGPF/C?([4Q>2^L<&88S
C:5OdDHP)/Vfa^6-fd8)+^\]AUbFWAAK#WT<:./U2I<[Z58X5RS^Ng0U6QGf@,WH
4:e\2/PS:RMSWZ9d7E<:VR4&OKT\-+P1E_^8g8_LN=fF=7;>#(OV?M9NF]X&G:YT
4N/8#-<G6=-S,$
`endprotected

`protected
KcX43#g\B>;]@V<BISgg.](f2W>fZ+[3B^YEf]\:A]TJE:@+MFY:()R9Od<7&d16
f)LETM,H2XA]0$
`endprotected
       
//vcs_lic_vip_protect
  `protected
gL_/BH;5R=?/_FMc^WB;NB)T1MVPVI99)Z5M-)0UI6FD1W\X?dEG3(>Y12.4PDG4
8WX1-\M.6<P3G:/Tef:Iae#AX;b3<+9f&>MZY9&D:Hb0EP=8JN>,G3@<9MSXc]J]
BI:M.\5bGCcE36SN.W_?H_bN2ZJcR7;:\:Z&SW_b::EMM7PfNH(IOTQ0DZFab)SB
Y)27YTQU0[<;)^-#;I52+KbS6f(HF_Ibg7O_BCH,RRO?3S9H[?EN+@[]5+LQOaIa
5-G=?)U@AGcF50:&a.-(##30=D(7UO,FKDB?F&]Cg@gU^FSgPKIca#Ne3L]MaE2=
cQ,2U&PVS5>Ta@9T<7N;L,,aNbRd@E.7-@ZT;(J-[3DZ_0A596\<&6;40NJX-9+Q
JQXc>#a;g04WS-ca:C3(Z?P6TVTY+FU1E]N:1.&_2EAZ=Ae7[T2CR8.)H4\3f5S9
]+ZFRGPa2>?8QN7_J-,WDJ\:HKVHY8C;B_./QWD.8_^^7Ad;X2JQ2G/d3IWEA1Pe
4H:V57,<5G4:VTf-84R^>_U&U]WX^\eRcJX<@6CdS.F66OgE,-#52gg#0OGL)R?M
)_RJAZM4e1&R@5D^6]H+d?CP#>O^C#[##S,[()?YKSTX,bbK4?5Lbg27RK)#+UF8
T9dYEV/d79gA)-N<:X7[.,SR=@+>+4DG.V6=W6YYH86+<A4\7a/<.BE)>H&CeQHN
#S4gI]B6Kg__8-ed2EVQH7-/M6@g-/?LW1,@eFY9-39M,,^>3YY1ZefAf[.2Dgd_
?/S9f?9g,.IJ7D8CI/c57Y.E&c+AD&4CXJ8&b#F>Pf(7E3E#68UMUYe.C9+)@_VX
&>I[aY>G?=\UM:/WHZ59U@;O-KU7:V^Ze:T411c4/BNBe^Y)5?BM-47#T4Zg1#9W
eT8^4,H=?.MU0$
`endprotected
        

`protected
GB:G+b#<(@#?SN>ER:LEV^=<]:E4=GRJE9[O(D8/5O:PZ()UMe3_-)V@[D)c9b^9
PZ<eA5LKX7N?bfQAZT2ZOZ/VHHa76(+bS/S^QDENeg2@JaaU87?:U/\Z>F4S=(1fV$
`endprotected
        
        
//vcs_lic_vip_protect
  `protected
G2)Y(I@U#>W2VJ;A/PbX]WA#-E+(fF)V0^EVQY?KW)f\K-EE-I8/7(BCAO)>>?YV
#I2&Xa>a^ZZBX->CJL]&X<+,8\]2)#-P6.78M.]TcI0:KCFSbP?#:gIM,MW3I2=@
^.JH5;GM2Rc#,4M?>\-_B_E<(8=&M(RK5M2WN>#XGC1KTAbUVc6PG-@W8PNMR4U>
T3IEIg,GFV:F^NeA+(f5BFK6b?7,8.Fd2]Rg1GC=b/g#Lb,I6;K55EB.\<cFZ5X1
9f\&93(QBb]D5N6bZ_W?8,B@9d)ZS&P?4b][)aZ:XM+7Gd[^7)\PfW+RTV,f=93Y
1Q@fPDHHC0WfX):gBZ>[0(NT>=9J>WI>6PLcaZA-K?KB:15Je98d#S)[LOR0I.<@
bC3-[,F07XBT-9,H@AT\\B\M#7<LENZ3S<_8J&-@@S=\2BIBcL>&I8:OAIP&.[Nd
MMS]=87?.,fOe,5U2@A(F?,.cC8FBO[BQ?OL1O7^P.KNR8L[-UA3\S9[E,=(cE:W
R9aS0LZ&;8W=[K>0IE/Had_>M91e67-=A/.9g:Y#e=S#8@7W_\ZRL<0KCP[I\E)_
Tb^b[]:P1Ea==P=VO8:6LH7EN.O^=ELec(YQ=1RAgNBdCY>@aNZeAT3BF)\gJ=GV
B]GC]1@/1OE)cWYD1O5bJ556gAZeRSH\_cPRXO5_8_b0B[\L]:PTI[V+d13#,IAQ
)GNUJF-VRa^?eD4L.(;.T[<6J,>FN;<OU1FM(e_?;QRNY?KG?97U6#NA?DGFc,,\
8.D74N@aCP;=V;=,/,#XfF]A1Y2SOS.aD?9DNKBJ7KW>@GXY].MOTAIdNEZ\^a9&
Pf/;C/:G779NIB_?554LFA:_B5aFWZ0U,4+^79778)XKFA)_S>J7b(eY)<cYDgM-
7f-O]eOQL6YF/[[>OOcdM-@9398MX1<4Ef;f&YV>/89/bGHVd;6,eZ3116U2_..S
dA7\54K:aZQ06@U8)4NK\CD1X2Y^=fE^)6VKg,V-L?5eQcQASae^=<0?;9Z,f:<(
6,MFa9VgfNN.b\:d::NZ15?OAPd.-(:01P9-b:&FgaC\^B?OI:X@Y&/WG8+-G?BD
#7Tc28,JaeIM3_J?9A1&AWX2_41>+(8=NMYF_:P_V^\S>^Hg695/7V04T)X]#RYT
;dR3:/3[G&NAgN7H+?H:Z6M.W)_)CbZI93g_NMFReBE^ZK@KMS[HAK;2dBB81H-G
^32P[Q2+^dd0,1KdB:?D](KH<,Ib?@:a?d).(d57,IKe&WMS5>:bISe:SNI2S;0d
-06DgSQW0[G7<5fA0F@K\,=:P3G\+I^U&._QA&0:3_X+8JNKG3GN=#EE2&@#+M\:
5)2b/1T>8]f(<VCLC^T^?=fXDg?d1:;0N;+Pae>I9bW2(S=CJEV3Jf>Qe9VFWX,M
(GJ@KO&LF><@a9@&\L(a\QDGGE,7VAcA8?S2VeW^^FdWR6,^K:F)84C_9@>UA0)R
a@E._3]<IF>d@HPa#K2)gQe-IJHMEHH1<dd209Yb5W>JZOdK]KfLT.\1g?O;JAV+
H#Z?XD/4e9]8HgG/HT7M.I0LJM1_4S9#QIBK;a@P/U2MC(@1O@/EXDWO/]WeZfKG
W<aPFf]Q6;MPCWHOFL,Lg+])-;O.ZR:)MDFG[dBg^O@OVCC#[IEU1X,+W:-4CITI
\Gf=;4F]/VbbOIM.8?9+c)GF)HK1Y?\;WKPJBG^58fNJKF:<R=#BPL4_Rd7;MBbO
&OPWV2;eC=/\FED5=7BZ3R?79+Y1WM1JeM<]PU7[)R1F=VM=(TMA105#DN<3^J/#
WL99(VB,XIR=0cTe1K:96L+bHY4@0;^N7aAX48M]ACgb@Bc#bCdS+1ME[9aK?T3a
bEaN+))SgcFUENJ[-L50@[DbBbFA,E/Ie3VB[+.I)8IZ?c<)>);,.DFY\NU@NFZd
_E4T5(Qg@:K_2_b5)S6f>:X2AHfY?Lf-8S<S0[UdRLZgA<b&?7Q#I\fQ.b,(26\#
]0<)(KfZ9OC5ZI;aQCZ@gR>5#_89R/SI37\@0P59]?8db?LS>(=3Pb_:4:>,7,WT
,VH5<(N&Z/6Ac;BTM82JH/BL#K-++HEK7EEb_(.AV5V@(:.JTINEQ]X&.\bZ\eS)
]U5?dH/U=Ib>TI?.c09<IML5]ZS8cCCQ>[.#E6D0_4/U.&VT<L&569>]R\@ZV[AM
cP4Qe;Dg>L3Z#)9c[C_X(2G8BaMDbJIX=-#<2[M,FCKc_XF&1bf2&):RJ:Tg];R4
N#KJVTLI/[BdV4QVVf]UU_db#@V2-5][&W+B]JXJ.@0<4.@AP:0)[T69e4DIYQLS
&C]F#(]CSTa7P_ae>_gA@c25&+JT4dTEQ:b>bdRSfcHTN)\d0,SBH#BNa8+?8F.a
Ha<c:aT5f=fcQ?Hc_OTUSeHZBD1,2[CFTVaA2;(9;^Q?PGORH>D_8SfF5?[A_E#+
H:TBT(<@4\P@?XZA>.:MYE,;,)fNZ.<.C],H:g^Bb^G-,#_c)?Q2/#._NKFa8;OO
NNY:afK^=H=_gP)(WLRU,5DdA4,RGR,VNM@FU4Q#If(fPPE^NI_OV2V#\.fQYM8d
KSL7=E^K0-D\6:XT7WP7>RaFeYVCb#<G#EYRG.fOUaEKVaB7cC,M0L7dV)\J-AW.
5<#@K3=[2T)U8CKe>0-0IN8g06ZR]/>AE+cMC3P=UO65.1BK88@Zeg92N.R.M#Va
8g+fJ.FBRI-#]N\2I9PfbD1;_QWZ6E1-TE(]63T-UaC=[QM79Y6YK7We]=@,^7U_
<Q/-XY2-UBfPSXR4JFQbH3;#e6CJTB?XXQC6gVb/ceBJ=TK/Fe(8<6IA-KO:;?fW
^LWJ\45XJ00HUYd01@IJ@9&UY,P^/.2V;PbHe&<4M0D[VXXD0=BG)PPVU77&;.b0
^bQ^#J_SQX\6PGYF-#\NQI5X_^I9A+U1B22-c[d=H5U7<f+DFQUGMWLCVSea]c_8
L5;MH;e(g(7(5#ES&HY19VLJ#ObNL+Nc)fNKCX>a@LX,NN?1UH?)gGO\(>Ob.K__
X#Fb>D<e/BfSY6.1[5LI,,E#ZNgg1J:1(Cg6Xa0Pc.6;&fdD]TdG[g;0La0PWU59
QeG<G8/P[;M:XEFa5>7SLEJT/)Ad]VbQc3Z63BGaOaa/NM4PP29LAP11;Z<P1&H\
P_g^EL4b_@CdE8^b=\X6XKKY?+0:P6/4AWE+cUZQgbdQ]>(,U+g7&K02(,AV[bbB
GW7[)a6H_>FgU3NbW_YP__9547S+HTJ0Fg]6/>H#O&=0\.E\f^N]U<B\97c7:U)_
g0fLdUFHTGONa4g(?<GV@ad6a>R7L\NfV/MagX76FTOJGPAV;V87FUd;5<Zc3cBL
>aFD[FdAGU.A.I3V/Q90V47LJF69GD<Ga44;K\GafZ#\VLX7]b/fJMOE>;?+OBJ]
?<M.-V?BVb\HU6V4@R..)V@EJd#P<7e>J-03^)cDO@ZM=d&@15&YQ,)G;P7?E5CT
1MA:V\8ADeee<Sc:4DCdQ5&f)O:)GY\7BN@eD5AO)ZC8+3?Jg8\+9,A_\R\(ecJ;
MLQ)6C0fQ(.S-eXf1Ya]<A60H+765W-S]bZ,6?6LNZ^F/]c9WbX1LI?(S.Q)EH^5
0RD99<e;GRRG/f#+M,ae4aG&Lcc\P;WWT7FE:71W+b1FQN6-SCH(@Ld]cb;ND7?D
=_9.+).W>_;BZ;+f1AL]ZWCdP^/(a3TC[N#&ZaOC\;,#VRYUGI:NV\e:H,6Oa-YQ
890/a3C3S&6#>ed_)U+\Wg]/3Y(+6@eVX2,H>4F:Bf,_=&S]b:\&KQBY</?,YS<)
Z9g\KTWL1;ceL&V-=ZCD@2(1B<#FFUMD@<9eJ1OF-Y[2AA;9IH)4XNU-)_8K.=2D
8T5S.8<d1>#DVc3)X-c&dJ3IL&WX?P=?fJ3JPTZ)DBc4\V2KC]\df9_3F@T<]-ae
SSEF88-CMK,Fg[>KCKa49Y.-_1W2J:2@H6A]8^;IT\;5+8],c59d^&,Ge<<.,J?:
+-\HFYT]<dC4bSIMBU/?7&?/[^&_V,1c-PIAJ^:HDcAC?1Ub9e1#Q5\20R:geSSb
Ja2ME8;UJ@K6-cWGQ_]_ZHY,ZX8/H0_]Y^[O[.OBa6K)D/I0#6[6S#C__;d(Rb.O
(-&]TP19)9ZM0<7]4LTc].(d#OBg:[5ZWXHa;VWFA+IB8P@bP3LeaHT^355^T/a[
:GeM+ECD(I:YDDATP0WQO(a=Jc36VfTc3,VVe9Df@\)FQ<\;82^]cWFG28eRH0><
_DRcb2_OZGV#dC(,a/f=(@M[I=#14f.D?b)T7-baW67gE53BNdF^2G-K8>P@EN(D
6TLLOMQed/gFTJ,>2\O6e8eU;UJ-NIY-TG#7W=JK?G<-Jb+RUM++@IP&DYe&N;2O
;2U,N)G0Z1)JS.0,cKH#./O-_G>K94TBA1YK36\^339-@IbWVc1^0#(4GB6]?^:Y
,H96+[;YY(B[]4B&a:5N,D[7a#A=Y,);=6BR=HZd)RGG2?NB\7\7F2fX1QFC,[;7
/_?42.JAg(&<1:5begNU]DS]R5T_.60Q]:4=#+bRQ;HUeQYDSN,d).[:#W9+GG^b
CML:]X2KbG(7cbUbUUU4bWZ1^,9GR](aOB^?_W3,YO1a6>e=[e,.=K40RHC.&bIe
;Wb38G.2#(d#SQTML?_P]aWL7NVWf,I.K184Q;>E)0TTWR,Y#a7D#e&g)[6D<F2F
K1R_KVNG?B,M(=@S55G&gR<G>WQO:&g?MPYeK=B.Q>^==PMV_2b.5+9,U3E)F9FU
<,c+U?JE4NA5Q?=7E2A52V9e^&DUJS@Z.R:^D2VG30SQe4IXU6dX/GcF,YRS?)UY
\_V,&8+(,)g(&bZWHP8N8N8PQ6(PF/OQ^9@ZZXFX.@.9+beXW&4JVg;[AceGE]#a
((g,D\Z@<a:7\fUI1B^678U+cG0+P(D(9Xb+b1dW2NCMB#gcf?MC]J.\K4-)U^#)
E<0.,44F:>OLS=U-Z:SKULfF02Df)1.VQ@aP4\g#.&OG.&22O0FeVR]e0YJ&Z?00
8K1G(d=3AKRJ/JE>^#OG(@&2AKf.e&E_;gOOX97+\EN;?N]RQ#G@K\_\\E(Vf:OH
8AA^YM^_N?.H;[@K9<E&LP+:+&cGENWZRAaM[+fX;O:7b7J9aV0G);9CI7bOb>&(
IE8;K0?LLL,?T-?A--P.G][#+=X+,N81<,dRWA1/?2eMR?S-ULQDR(X6J/2D^5G8
\MK&?c)-NRTHE18P@SaKISDF[Pf@18e^bIO(AT\<.g_Jc-QF4dQ12URM(VT4XKO/
ZcCF,e9O5Adc8OEWQUO[-I^]NP,)5KFBO<=2^cEFDdX,TWYa2^[@_NbC3E+,J[X<
/8=.3VSP?ITS/_fXcB2>YgG5SC3C0,3UT]PCYRQf_a.M(18#1K.0-3Q8>NCM&dZ@
0PWg)\4@R54H@c3WPDS/K>\R_=2V-J6:@[P[cK2@YL3KF_dQ&=dFCM0\<Wg3O=A&
6Rg+0F+&c6;b-9&;BS=c\P:TWZPY3R\V9cUc9GM7J7R;5[fWA0CAM8C4([E_^b/C
ab]\:@[fH2P90FPI)1RMGR#f[1fcF1:KB8P4WWcO#C_2J2X@?-DF3N8eYIN/>/;=
F(JX/>0RGE_0M#Ce9<0NeE=C;6Sb+.Q4a,K6#I-Y=J2>M5OS:,FRe87DJ5,]F&/F
G?0,X\]ZIAT3OcN7,>MRQ^VbB>5[I20L,@8TLF)8WHLWL,N<ENGa7/_\fGZO:a9a
VeN1YL)57R3:HRADITB53a8@:/?SC;5(XHHcYXS\:F:&&?.#A/W-E1D)gPaT\PID
4@_g/J0T8Q15NGaY(5@/JFM@]EU-.<X3#XBb&=R[=JIH?SN^=fFcU)JUO93RS0O?
0W4T@;TB;C+[Z.Z=HK4SEXaPN[.IP=^Y.UP07MZG#N<V(e6,He5SX86=)@O&NeL=
AWgbSTfM&SU&CB;=X59&A,D#/V#Tg,D;VJC_d[DH:A+1OUX(,-WDMPXM)-?RJEYR
FUb>B)]7DK/MN>5dT8_]GN&USG\RBg5/K-bU]02F=,XY9\b\e(X<O<XYE5=@?6?)
IRJa^9K_>MOZDER:Te1AdD-XYL/DcZ5;5D@E_P:19d:E0[6[A)JT.^NNI=3c<O&b
NO+g09fWA26Ba^AV32_G<DU?/@V1TM@eEgOB+<,R>[&N=FC2^\?J]H?LWZM6\Q)_
(4;Q<;1U]BU@><e7L;g>I5fLgS?&@K96EU.@^VOc7aH12ATXLX8/gM2ZUd+ETBJS
aeZ/[eL_3dZS=S<6B_:CccYLGFGS;OKR5QX?M?PDK:?KEdM>6,e9]<P^.DXN1VLXW$
`endprotected
             
`protected
;eWSb:CNUC57GP8M<3924]f0U.&(H78B<R_CLg53bUY-RM1D7E7]-)3Y9+=&F51g
\/GUM@Q7ECeSaY](BIL(PZD5bGCdB\b[f(RP,HI:Y::G>d.4Z,2E]a3YK$
`endprotected
      
      
//vcs_lic_vip_protect
  `protected
>43Z5dA:(0;0Y//=g9\VFP:>ePI#I1g+9a&?Nb7G=b\)B>?,P]Z#&(PBdQa6g@HG
f/a_:RT8/E^+1bNa?H^/[^-K)Y<0_EKD+HBRXH>;BWD^M5;SQAGB0YA)+-O<BL\G
P&?<D>FW8:0&C=e&bZb0N.G@KO?;,?WT26A>bHKKEG5]F-^Ta-=>@2,OR/J&L6.2
^<>I9;Q\0#E2Y6::,J@fN2<?)W)8OFLeNTDK&;&H?gO]3RTRPU)X/d1cGVPeO.5(
O2<ecP=fO?-/WEPdNa(?[UVe7g528S]B/05,D#,NeM-2@U@=)ET<:f0Q77R[&Id7
A),CD[:N15f)?fLcPY-9S]E\B6]KMRJ?CK04?G1\Sg>g9;CM+0MUKaX^ZOWW@3[W
OfWe#_>)\J&6+_9DKLFg8<\^D0_eE[\R#SX0:c@_VK+I>c(E\57-cf:-5a.YJO&2
^E(X12>LDL+ZX;G<gT3C>5(W3bK<S9;#7C-A#UQeMUBd9d0ML9C735[[?d1g(]OF
d30-:dU&X?2TIQYC2C)?J&F\eZDHgIIgD+gWL=H3W9a;JVB0H9/QVZF4-1;JVG-Q
LGcM-?<38U;VOTM[46K)#1\QBM84QII0XVSK@Q_ST9_GZDEgBgM?8E)-YOW-SBPV
W(d?3,NGPY2#J44/7Sd?d:71MSLYDd6;-8dPeg5C&F#2I1ggJ:I/YfH=@L[&JY91
MeP_C4ZF(_QLY;ZQAY&bd0,fF+J:cQ/MUE+BH<1e1Xc:D&;NP].MVT6@LaY<HI;I
2UDP\@_.g:S=-Gfb&XgC]U^[bT:PBPQ61+cIbW5-.SHUf.O6W_]//.X8f1>,/?G^
HaNKE#6CU9]T_;)WYg=gH:J3JC23Q]Hea1/.\YB_?^f5K5FECOFH&T2\Y,](^f7Y
4&-Fd?GM1Je3O?)/VP\X]SADKT8B8Vf0[Y:N1/C\e]JFb<UNeM2(2Ic^S[SX9&WZ
L.LCR<OS/A.;.QN6Q#1QXY\W94U6YMf^5-Wa=0D3>?e7SaZLX(\FaMLQ<DS/D;;I
FfJRSMZBY[^6P3:g5SMaR9\RZfaR\^PA1J2[5b7e,M6:(X=KRcGR6Y2Bc)?JDc]P
._@#e/N,Mb7CCA5#6#GN=?P2b_SY#KK@;g0K8LVc,M=caK#1>?b2[V-Q&//RRf]5
8SMF.LO:OEEaN,X#/UZ];2]7@C:6Hd\V\gQ50@N-+LGX?[J2VZU4^d@3?9/DHO7g
N(7CXL@GL;Y\)8KMA_:fCaL1aK<[.Z>L,=3N__F#W^1dL/A(3KCH/])^NGDJM,OS
@c)G29gA_<DNHQ<ZM9H/;dKc]-@70aL)Ka+KR?Q5FaD:[EcF_S@8MF^NL3#(CWK?
O?;fG6:JR2R4R5WTAO3Wg7(MXc_TK<2O/0V9)@d(CXV><;LZUb[NE2SK0ZB#FIG4
Xb&;VR;c)@,@7A^c=)B4U3GAKK]H#W8/a8UC1H<ZN:FJ,3Q5Ob[2f?QD+7W,-@cZ
?2aQ-8Ee.?E6fV:LY?F#F.(LN8PZW8TU+,b+Y3S@JgAVH_VcQG<^SUZUN5?9#O.#
W6LY2(K1T<@A][[,O4EK/=dX6OcJ2:Se?V7KJEBa)ND:UfLeLNB(H_((dD+Mg4OF
[YFET.Q9.Ga^HFXZX<(@EDZ+D[PX,7cXVLML-10D9c?5:&OY^H=X,9R9;@F-/C9-
4:E<fgb-[GGR>C&7J)=L#-a/=GK^/)3e34(P<2_5dPE#aD8/DV_gE+fdT3g]U0OW
1.8<5N93HHU/4eM(CTC<(YW7G^^T@=0-0K?_374KG?E+.XJP-C=SeKI6C?#>OcP=
Q6:H2L]>T8a3eX/.,g>(c13E@IEZOX^3Ke,e-_?X\:\//Z,d+:egN1Z^6ed_XD^O
,#R@\4XDHRCdH2K;abXbaTL&-fOTSE+AQ=_/]gMQX^\0<gTf1^1L.#OUW8/\CGA,
45.C\I_,?M8cR;8f>(aUaX=cK\\B,,<:<dQ=:.;4NbHY,U5R7[AMS7M:JdB6b@.e
Kgb?8gLVOSfO(4[(A+1\/-^^77+F/0f#>b@?SD#YM/:-GG/P0)@ZLGX_4@2MU/.X
\T445);B3f,VYAFF98:NWO>F,V?ZYV(N&HMS^J1Z2L4e6D^BfD_)U65G513;/>?;
N-WKUaDWMb[LL27f3(BOg8Ha<)^]3)5DeYB]ZM?H,(G>1Ha)EfDP,24X-1CDQe,L
&)\.Ac;U\L;+1b5V99R7I]FHf,fY+K7TX:S?GC;Y795a):eQXCC;-eI-?5a^ae.1
:IHED&-+-3WB1&M8Bb4XWJ?PX0Df;/\P<Q<2[?#L)+7.Y&))JcYAK=V/2?G@V\.>
P@.<g]?C/E0&CIPL,Q+H[)Z9bJPB.U7Me&ca]J;VR-<,f&+MdUIad55U01Xa;#>E
5[ag]KMOPSQ(8Y(L:MgG82T,U.OcL+P3fUP^R/cA7&1V8P4Zf+e\QXT#2P[93HLb
FR\)[<ZE]f8)TY8f&[OM(P[a6ZFe13F4;3b1Q52[O95PH@_RCGaQGGE(+&OeaKN.
/b24)NT;)>=7FDO3-:W/QJ?OS\6eW8_L3Z-WB=6_1W]66S_/)6X#-X[L1OaH:201
bP)]O1@WD7PJ&Cff...J0AP[=:OA1_O4aA-S=R,T&)PDa3f6R<^d#^>4JcO4(7.F
_dgOF?O7NbUEf&&<><)V&ZJ,5:-226S-<#4GdN9+0GT.N-)THN3:aDL?N5ZUX_+F
]NDLbcE>>\BU;TSO5YH.;_,+NJI-RTS4[+R^GI6PQ5/g=f=LVU><EV/A9Y>;1-IT
+0N^].29+/X,R57-=BS@gFaN&D:@(JH9f)MFQY4/NQ<HEKA?;LL15=6@<S3R9W#H
[]=6aF4IWXdG]I&Qe97?E/LbI&Tbg5P_d83H_-#J.-1UU+::;^F7(KIV;aK.e5IK
.A+.QWae==4EMaK_0#a92YQ+7L<OG)-dCeJ^M^BH)X&&P.?:(4+I=55FHM-0[\1(
ZSgK0^\f-MZ]bSAW>a,VD(+4+I[g&(?758N_A[4G>8+YHVCVL5]WIZ]\()5P4Yg0
->0eYbcf4@T&L.bKb70F1bK)=Re6V80I?&6B::UHC1b3&BAQ2W9.M0+2)1cZ?-a0
Y6F,6N<LF7P+OC/(,_+)R3V.P4W<M_-[.bF?YR]?GX)6+]gI_PGR_B_bSY=K:&>;
#P_(PW4;XE0:f:Kb;G5eY,6e6QUJZ#HJDV3QIB,;A=Q#fYN.0S0_N+TNVGVUS=(J
[0L1WF4g6S,/2V9O\EPf/4@592FPLC:2<\JRLb1e[W)UgbX8+=#&fa8Q]<a4_Q4Z
OC9\f<Z/>K?b__#AJVNDZ66C&d4M90E[XOP8)Ef)g.H]I>[EDA<WA@(<CaA/:IS[
GV+R&S>GN3RJ,A4?aJV.K\90-:\V#0HDM3LWcf:3CbAK>?<VOUF,39JQM6+XHA82
?T2Q=ICQ^J824>JE56BT2CR&^gB0c(/&56B(0e6FLKSP?IKZVeJ.>NT)2OLbFB1,
,((9-,9-2Eb&a5T@FdA6U.;V>cAP7,7,Bd^a;HO0R-JdCaI^-ZJ,M))>2R)TTXD]
Lcd30RH0K.fBONPV(:VG=L<9K<Q,K&C25]\)fDF-4Y4^9P-VBd>f[Q#GAE6H@dg6
FN(1)-L9@5^Z&F?/42/_ge?VU<:\a;I127Y<.8cEX^^5bS9[S#.XQ>Fb5?OC8/a9
aUZG8Xb>>8d1CI8MBE9,1I(_2F01NZBX#A9/Y+OVgdSXG/Tf2\1G84&#E<RD60I:
JSDL;\V=X2]bZ:&W.CgQIB8cbA5K34#=X[VCRUIbN?C[ENS5WW-/C2_K6HN80POM
Z[QbL55C)0Y)\?I=;.92<aRK&)OdJ6TPJ6V2eVD>cDXE)AHPbLU-fJIcc=<#+QX4
4A^\bL?05ZMLe1FgJ(8gV@2G3e@XX?6VEI+[KFR8B4?+C\EU/9Lc&>CA9;DOCcR@
IY:G1,Jd_3GeRBT;-c#Oe]NNO[S@Xa0.T43CJ],8G855g(V_W;0@W23<G5)B4N/b
0G:#HT[2Sb66=0e:<L?JE5Fc;IRTbL6O],Lc<H59T56;ODNKg=9L;DJdT-b(g60S
OYcA,SbNPa)_Z.KS9JB5+@<D-0-Y1aO=^YUKESVSfLF>F:U+R&-P&)\P12Y,N=.Y
+cJ7c3E(#U1bOCL,ELF&P@C;94>BGES4.AM+\12<dDSVb<9U[\P9G0SZB^19<#aC
/CPN4Y+_,7NGJ[[]7>.FDIEXB<HHPNAXcDR>>:0Y/gb^U(1b_A7PQ+()eF?><\QP
_62T14QB]JW+UPNb+\d^-/2UYX<#1;OaB?<#A(Eg#Jc6U(DJ,GcO\>8+&M^P&:Z[
^[dN0M;J^g93A4/VEHM##\L6CXHJ57.?MGL3T)FI^FJ+/:9>OG#6.R++Cb^E@WI]
PeCG9WR[^45Dd-\1?:I4<,?GE5eB8<]ca<.<H9U@9IdP7@b>CRAI5BOJ(5X=;g:0
&8FA[=13B3fY457,HHbBfA._YO+K+N/B-O8Y\NHc&F9@W]UARC,J-?0VCD^M>Z19
ULZ]JWKG.O.#S[X/I_7PJ[G5\D;KOI/7B?LFO:MBN#,<0,>V)+1O\6H00N]E@Z0[
[bC&gPFUIJJGOV0E#J27IEB[9NCW,780E[BJYKBJ@&JaNS0MaX<0&fL.[f;9VB94
TWUM0c/J?8:#H:A)M28F<P2IO0/a;9M8LcUN[:M][@-#KXc&:V7;HJ6]eWONBXd:
JbN_#QP[8be,4W_Ze)[A3-f_>(8EIC2f\&(<@BFLOBOcJIFXWfd:E.CW5SSXKPJ,
H(=S)QIe:K0a7D:V]=3G:1ZB<>P1#9;CG>[99(Z13(eA5KI1-#b.YC):&?8Z2NcU
QJ:eZGLdD^CTI?>=FCM>JGNB(FY+(f)+1WB&.&4N[P=2\gF#;W#gG,,?aX\,SgL0
B:&ZZcVY7P+ZEQ)CS\T^M;FYZe=g5E\8g.O6POK.M5U_7.RBZ<MALY0J4+>CUYgK
+@U+Y5?E<L<:>.VK&SZTd+8d-Yf.WD<5C>>3W#,dW]8Yc[b21#_XMBW/PS,/NT-U
=HP,F=IGeTJ81Ta/::]_TBZX-cASJQSG4P0aT&PJ]/454-)4eZX+;MENM0PZNd<-
TC3(_EVCBSA.#Oagb+P.AGV6Rd=A;T]1K3@#F@ac+eQJU5R2T\V7U0?&H5_[RH@6
]R4EUI(_431TNABCU_(&@A,SR2cUS+fE5aTS8+54Wf1[F;>FY(cY=DdIV/>eE(7f
@A8=H:7NJPG\I,=a@S(@7S&O3V79__ILWa-ef#eOAGG@@+J^)7?S\N5+]&,EeJNe
=4XLE]F.OBLFL.<ZTG>PV8a)JcTUc]5YICM&CD-R;.XLAL=:A<T>87?c[ROg([BD
11;MJP0H3H>G<A_-#]HA3/?/0Q5I3D@;R+0HS5MUfdU.XP+a6?\I@D@9fFV<540f
@_1L.@QF^-K(b]>1MdTGWY1.,BQ61,SER0/>R3;TTcY=,Z3E[)H\Y+C\F3/8M9)8
:<X3>AEKXC)X@Q?,9QR3Z,D-T-OY;-[=\d;:^-KXKUaIEE;BG5eLcgaf4MR&/4E<
X1<d(7L(VYe6G(BPVC-?[=;[1/dMZ2c\#R5I&10?7fe#Mb.dg\RP6gH(a8]?+a/3
eJf_FCGE2DIE1f8TV\E1V,S<U[PNeNf2R:4C5:NbR0T5UD3^WBLe1/2TI\<TRW.2
8BdB<][G6)7XQa22HM]YA+gOXSKF1C.2APD>dW<#MS]UOKC4gYaRS[/IGX-&YE2_
1>1W6Q&Ze5ZeIP:L3e?:9E[C+U=5^NKgOc-Z^^;00=a)(=1ARR8Db<IcD@,1]CRN
DV,+?I>AVUgc>Y]PFY,^8+VO7be?Q.DTGX/\>.<P4OYVW<&:eWdc;J]@.XP/8Qf>
M+Ea3FK.--4?,?76]Pe<Z4e@4D>U:K5WEgR)a]-S1P/1ARg:;T3.E3BL2WB+(d_c
;H(3LfV<)LT(JaO-#,>fa5)WI_:4U<;[I1#TJPC6baVU>HVOZ[2SA.a8X0]\FeU<
Q;#-b>9TQ,]We.;]X4H767UPBacPP&0BDDbD[^A+0E3<.L2A9D:g\^RBN+6bb#7A
>.&_?MMdgIOOC79DKcDd:/??]e/I<G)2;39:66:OAQ3cG_I1F:6@bYA=Ff4WPg8U
[bTT;W_#&e/9dO[7dX+E.ONZ;K\P)@;U;LZECH9LSNWc:TT7])R;=GZ+9AfT/CbP
8G]dVD@E9@HP5&#Ye\W7P>UU4e>6.3dCX/3EW_f((7?Q-Z.EAg\HN8]C.7NS]ePH
<e[I-,eg58EA)8g1ffgOB<IOD5Z=Wc&4.UN0C:/\&1GMd1:8/Wgd&@bHC7\A0If8
I+L(]U,+:_&Ff+gMPO<:B(,=HO^H0M^Q#=DD5@@#cXBbEGPBSG>dW<ZI\A3J95ce
^C;EM-=9\8;MR<=6L:cTCeGdS&E]g=\23&MNOS\A?JVQSe&,eU+P>&+1P?D^a0DM
;I>M7c+ga2bS?BFVECNZeO<^FJ,ZaQ+=0XJW624J.P5=K6H\LCgPB;6]SJd#F<bd
YK_?23g832AWBZM&[BEW#4E6-bY5(@M99:XMYBM?PHQ;E\P/C3^<gX)faF#d)I<2
LPM(01KO1NCW<;BP[3GQ<-_J+-eY+X8I_E(PC:\U=Gc.<MZ/fTC\5#beBEPIU>C+
COLWQ;9EO(f[;APAUBCP6;>ZLB6I4HYda6CX8L:@eZ5?fN<XD.dX-?5G]^eZ0CB.
a26dX<S?FE?2\F:Zde0/0T0,+fN^ff+<Fc]-W7Eb.GM3WM7V[a)OU#+RX&8=B9./
]a.<XI[01^[JGA\]G#0GB>KSbac7++_L=Tg\CQ6>1?2M^+M-E;\-B-S6?S@dTa+&
PQUcXYK0,_RM&d:O1OC^IAe4J^X16LQ=?#U&50d3O[JI>(#Y6=CMP1X#5O,ASFC/
<XQT8?RT>Z2V3?FcMHfT1f_EJ;Z<(=@T1_GHC#,G#Ob:.(Z>O-^JYaM=W)M_Tgf)
bW9Y:4bgA@ACS9QWQI36bCLKOg^43HDg)M2R=1Na&,:e(KE(2S_K:UT1A8Y2V@g<
dM(CTU4/GU>?2gGcOd;6Ae6&(]#5L^[g+c33f.4C2R9ge=caQ;K@VQPdC?E#C;+;
;\EHc)@>51RULWB>+d1=L.4:8?<EDB2T^7U\P>=G2-fK<bc?#:T__YGa4P#_;1F3
,O@DgNDbNHGZbdF+N,c>9U1Q8R3b^3^4E?(/N>BY#RC:@Y(Oc_2@f<^,>E\P)f.-
D(0[^=a[B5_Q6?E;P9WEbCB((81=8FQE<6(?#3-,I_>Z3cVSf2>?^N(DHbY5;Y(E
1WWE\;XBT#dXPf]-HB3NaGJI\5I=;>#63M;O[E<0OF^)GL[b\[G-:Y,aT7\/aH_8
Q=PD=EWG5+\d/#a>4.XdXQ&+O:&@VaM9d;gD4?)9S)(8:2Y5.P3TI>(-?R8A@c?T
I1C/&G/LH+83SPX)X_fgJ;;/&I^-PR5NH].(_ee&f4C:>16=aKX_2gOB^^cH3b=[
Y],TSM=T7_AU;?R/D>:.&Kf:H4&cG3-(Xa+a?WeEZ4MI,6WV,Q6d[FcZJ&E#9RcY
LQ/6dF7H<[a5L69:@\/25.0@G9>?W)0a?O59_K0?9[bPRbE^H3>;4CDR&D5.C_#\
3SXa,DFH5KU&)Zg7_b[B-KCgPYSM-R9d7[OYTb\]AU#J7JP_8X::3Z7Wb[4:E>0<
[XXaDF1Wf/aZ(NJNd;M.VY-(AT\E:ZPf;Qb)M+8741::dB8.)]FQ;cf#&+U>>-=E
+[\Ua1TDFWG[/W.19,PdPV^:<3682;84C/1ZV=>U7S18]GgEVd_\X9/A^65KaWX9
=;[=3W:f=S#gY28D[fO#Q0,>C(#EOUYF0d.=fLLLOX)2<1^JY24)3:#Q\Rb2ZP<;
@I&8+[+CDRD56O74J#4^<E)?;Q6?.F=Aa1F+b(+1?-f5HEe8H).&cO8OWM1d\2@U
(ZZL8D341.+;Z-O^XgBPdI]8B7KSb3]#OO.:)F#J>7H6=N^AAFZ?R?B^V(@^KZ)?
0T47Q]9^Q.FG;eRMe>6BY40T,VQWRSEL0bCb9(VIW&6f#Y0:I?<OWTE4HH7e[A:5
#;=PAXcQYe6GecEReSH)O6c?^W)[I3YNfD(eOSYRacT;88S3e.<J2-aVHGfY?4aK
D_A9N/2X\=3^@S>;K)W6,a#KNW45EMU/U7b1A)<1JQa(S>)EO]]97+@4a3F]7G9=
);19f:e(I,^:OSS#<>FbH\KOIfb:DG/VZ6,QO8Jg[5D/L_7T0#S@6FX939<59L=g
RS0>Ad3Q6_4e7::\@(<(\MUEO6T\5::J.X3GMBU>[dB57;g#<\RfJP-:JbF-+ED0
N69<M)DJ2eUA:f=/eT+8+W\\]A<GXMCZ_+P?d>7@QP\\SRc>^57D1\C0b&YMCZ@+
,&OY[g?VbM/VS1=1#c^FPAP1[(I6O^@#BfZ@)=-JA(.1P@c8\+R_3F)eMN7O214S
&,=CPL7@47\]>>JM(Rg&W?\H6/F>#S,b\:[\a-;YD2JIc9<=O/,0]K?\g<G4eC8[
\1>KCDcW0_P,d^ad_Mg\M+4FXCZ6;>\b:]d^LMK@#[W+1<<eR3QH(B[[[6]6L8[9
+\Af^75:^HJde,,fgJVT(8.L[V@fM1:@\2e^T/,X2X/CN4;:N0(L;S>N&F:R07I=
MLLb-9MEOP5[R4=+>IDO4L.;AJI]F=D/YNb&f>;80T.27DXA85R\#P6T#-=KG1Rf
fR&_L=Q0DbZ.3G)>E,58F(bNf^2JGNW(2P0.FgS&4HE=DK5#WJM?MbO6H=<><2]A
I&?1]SeVC0D85P=@TGP_ZI_@f0/F247IF,E]g-^fNDAO8=cdbX+E98,aA<=1-,1b
FggZV3Ua6H7;8<;)MbHQO.N66aZ@eU7KK<_W]b[M&.a#WTZf+T847;:,LPC;3+b\
e/+@HWA/^5aVc&C2.Z/f<<;)H,28U]M+G:OKGRP7Qf4]),b,V;ZP]b^JN@/A^f9^
&-26KO0>IBEgKVCE+bQEXL8\=WMGWY/@QdVeLGWWUeSV5+4=4^\W9N>\.)N(E31B
Z1MT/M8O10O)8f_:5.SZ&B/#\JOKYO&-TLI\FT:1TMP=7-V>B2VTMYG_CC)\L^&,
^][4:YM6<&&089,DP]Gd4Q6]G4,8X-#/2Vd]3J0#,#1?5a144-\-+B,L&fXUb8E?
/LR];LXcSZ@ESg3FA\(352cS+ZeSSa^ZaHZ_V^YG\^I/WSSP)I,2UR9f/LR=JA3]
T?dK9R3O,QW#T;E/E-KHeB&QUKV^:GS]6g9]P.J,A6]&+KgPU-XU>CU:/X]37;X/
a64:P]KR&@S1&OY1bH?f2)W2PI0+VIbc90Z6I)R,>=9:B@&AW8=P//2XZA?1&0R.
Q;TK+BEc&Gb(L>)X_:]VGdTKSI5=A;950DR>HD](2Wb28.ZBXf5R_9TS-[eI,82:
JfU>6PJ:TW<68EOD)P45?6U+3;1^_K(S63)3&07J,;b_Y5c@3cdI+74.+aXTN:Rc
eL,LD]7;=-AK7J\LRO,0:?Ef:Qe(2-Cd[1Y@_M5;JQ9=W/=SEA7R[&SIOX=0A0GE
T</>-[>KWdN<La9<W)RZ[G)a,L_cH&Y]e=?2N;cRE00GT+[/Q^+bN.M+Fd[]2S&D
<;ZfIT[XPKSEB;3Ma>\MVZ_FD511IELH5_>&:WgDe#9:F_)=c?FJ/T==>FY\OQCF
<QgCcP&\HV^HaP-U]+X>He2;Ed/JP=H&PF:[R?J<,b[V.(L)a9:/?C0;M(D]:Oa,
EPGRg[&\E-^K;4PYOKLea[;Y;K#SRWQ+5ZR[OO<W/3G+K<7?ZDZ16C.6E,WcI93&
aEWcI?0f5BX0Ja.B;U[Q^;H,^P&/6VEc;;#L(Y;23\@JP@;):ZK=>CAB#CSaXFO&
Lb16?-ecU\&2e9Y7eV)Ef(4[P=-OD,>HXJ[9>&UXE<98?&=GW&K(I=[CPaTZ9cE=
+4(c@6GYQ6Z-N7g4R;2-g0^[ObC=4=PV:eSJ;=O+TX8R:.b8dF\/eT].?:)TW=e#
G8^Rca5-e\5.d2RGCZ6dYNBTUD-8/JdbfJ(Od+_]+W:+&V9B(46YYebYRV&4+8IA
EV)2KZ.,Q(9254H;7[K7WHN&g7[@e4EdQ,H(Z.DHO4]D=+Xg#d9Qc##EQ2WZYN7S
F&_XI^H]XXDQ>DUR=@MJ\1^](\RE=.57E/3g+8gP/XaK0DGPL;LP+>:Jcf[T#AP2
SdB]P9)B9Y(B3;>(b+(]BL+d3HEA/4Kb<J,cXO6>L8Yg^OWF;UaB>MgB8[+Yc3G)
[_,(YB.ISK)]-8SF].Z4E+HcN6&@JK/cO:I;c#M+G)7#6XEKYAR=dY82GUg#[g:U
6J^T59a7AI7=N)RXcDaL4G[S93_I,([MC_1=ANeO2#501]fV(<;YdRO<eY95e#M?
ce>4/ML28DR@C5GEJE+e2GN^[ES_Ye^b,[K:?^^VV2\BA\1YC-0,X;N&#R:^)=ag
;U[P=cJ77<a;EL\&7&>Gb#UgEM/::?](NH)gA/D0O^9fK#FQd<4QA)77::VP&=K#
2HT)(<T=.C4NC0CR=S-7<8ZQB<g,cZB[,COQ[N68,KCcLHRYP,HcgW.)OA:<&XG6
[#](W]Y\:1F=3Q6X(,WT0GV?=FG\KN.Y<9Q[bdHK@D]2dgKNYJ&-1(M@Eb1K_@/[
[?]N>b<AWd=EHOVE:PS3\g7JJ&]F.&,+g3e5.dT0@\3&YbVP_&BDWO6][X6IO,K(
b+B0_=V]L1E1H,\g4B;.)[CX-aZZ05)2C/HT)Q-SC:VN7>4a;>C1-,_0(IeA.=(Q
Z778bgLJ@9:4)d:\5d;?_N#:&Q7#GL2:Qb[0Q8;EK\5ILI5Sd@VB6&Ub)ZdNPLQ>
K-H5=NQ5G?-QeO+fI@845:]V@X?E:>MaPaQ(?O\9Tb_5N2C_VF,EZg]WB7V(Q2V=
CQEG(BeKTd3C&ND#Y?d?0/-Z=-5Y<M7,Mf(Y6Z[R=a)b&#2M4CL=A/8<E\XN&71#
K3IMF:G+#:2SbJLF\SE[;53:B.),[WNR)CeaEFV^?80M+F^Z-Db>bSYCED6\MbfB
9F[8Q[E;V[K6MFEU9OZV^FcD_3I9_P[NHKHP=1aOaZ)2dgJCM==e2?,Q5YbSPK0e
E\@6]6[?NGE:6Ze_,La3R0-4[_CfN_):c=14@+@4fV;VD85S\P]6HA8a3@#Xc]9K
\K0:A32<MGcA(<53D]gR_3&(1=dZ(\FC)2.5)_9ad;MC@QQSMZN61)-MMH5@Qd45
5LZ_X<ZZV)cP:O30g4^/2:EWV:LYHbNFSWZ@cdTTV,cWD6>L9ed^TB\Ua16;(-?L
eT;?e)+_#L3(YV=_@@US64@OMCYB;f4I/DCUGT\+K[6aJd_IUZ]US-G4HSa8&RV_
dO3/UK<K<<1OV4M=J[V/#O];D6&K.&]f@8=Ya_F]/fURV,0F=T3f-JOXNK476MW;
W=bZ<dRVL.#&E3?86\BSLSe;@^7QV][C<5ITHOV,(/A=&R@[e^]._;^.3T1>1;;P
GcV,JIAaDL5_W79Sgda6cY>K#AHOJ^OAG@:^7:T118L]4J?JWeN=+9K/b2MED],U
Q;+=+&AR^V?9AI=P#bUE0->(?9cNZU5XXMM&OB;;6RKcN.P84,bMK.KJKQP.,Y1]
cgDK=[82a>+A0:=C#5)92RS</\VF.N(YZg6FU<N1fR\^7I8B,8c=]8Ye2EQ\?FTT
&.-Z(1FTPF1AZ]1S2[Bd<^38G+Y>QSLX@-6FHH+N.BCAeU]_C#KH.bDSV,T^-a45
3,QW2)//3\L;U[Q^R7V<XL,\_^&YZ7gR,aH=^?eY@S;WY0YU&[)g+&CCWMG?W0O2
)HWPda44,ZdBYQ3RgN&F84W86N[10F]H;UKO:4a_D[eNL@Baggbd=CW#W^[527)[
JL@&]g9RGcIL^X4=7C1[)2ReDQ>C(W)fb@YSDS2_L\NeM@0f5g4;NXOT<:\FP7B^
U>S<[c(3#XE<5XPK>=B?83DT(WOFA:WI:@/?SABb?:&=:_#VY2:MD:^TG;]6QT?Z
\&gD;S1[ZGSeTca(f&&XMW5M?U1D7NLKBbc<V:3AEHR/Q]X/\c-,?2JNa1/@I-=7
TE<c=];I,VV9CC.:4917@R&\@&PDePD+P/6;UY)gZ5)76<;/N&&-#M,Z6G.Q(J5E
g38@.=Q>T[EL]50P>.H:QC[_@R-GKgY^EMb,Xe=4B(LP7D)@[:1&BGXFWL+M1a.Q
+8C=^c\39>8M8?M[fO>ECE3_Y+;NJ]dLC&R9e8(1R9:Ag@[c<#DD&50\]5Q4V1G?
5U:4Z#gGQEA\/U&ZCcSZ#^=L2GC7,]MBZV:40,BDd]P,FJS7O[>1WK)1>;a50e)<
>WDS2,,&;01bXS7JP7(M0LS=JO8X.MPAX3.2Q&&@3_PU3fT+[a+UQYBJdHOQPJ^1
<2?]>eJW:FAY>MK&]K6.QMS+:N:f4SK5b7KG3]VCE>32Xa1d&g8dR^&:IeVdT+?/
R1<Z=J:?&DXe79<&Yd>F&I25,#(6;(2RB[JC8.:[Y5J)Sc@[WV^]_SK8^#-WOAJV
U-_MKR(;>T,NbaUL<E.@>LX>>6(4J8GTLW4e#UBK]>U4BIHZ8)fA(MT1;1aMf)>0
ce)d^K5F4cBcPCeTA<a<LOX10>CQP>Hb\&_VWOCJg;a#;XRe0+ATe_]M:T-VZ9OI
-XKA-.J^U#g5[,Sc)a7_?PW(:,XI2TaI^6V8[-G6;)Ic5KM/08a(4B+M9F\cC10.
dHK9KFCA7U3^KQ+\:UfS50Bb04B&?O+P.-M/ggAJZFQe^RcTc3;eY_KG/K.KdbGM
Q42V.8P>S,HZ>fA^+Q8J)C77Zg;aP7fZUW,05cCVQ+Z2+5<:Oe@+(_#UHKBCY.HC
aefTV&)K;?H+gc(/W.LOE5=dO.1J_LW(A4=>##884DWL\fg1AG3?]<PFJ;\J/+aD
2L)7N?g8aH8?PQV<Y0O1(gR057:L657Z:3)f>Z+ZcXA_/?EN6AWX_^S[2?BT_FcN
W,?DH\Y=.X(W?ED#OW.6YK?f6d,Z,ME6e7+QZ4Y<9BdMb2bHSR3YZOc)8:PD3S=3
TI<X)[T.R:[aE<-I8\ZB,_RYZZ7N/FXO#_Z[]QX;87>RY-eMePU2V_&DUa;OUa,L
>1<]2KVJ)2A<^Zc-FT(QA9Q#+N+e3dA]C14Y&IC(U,4F[&IT^1:3IV7&,28&0GV=
=.KTF.O47JD2]Bb/WQd2+1Q7(:^;cA^-ONKa6VQ3+FOGAP>JT<[8c9>].B#9eCS@
I0J(22fT)_6Q<2ZPdQ5WM5A-/NR1)Mb@\)C##POSI[\eKO6[A;VB6<2&J^_,g6)U
>8aBV@3S;fLVG>9gC+O@XCGgcA7@I;=4SBLe>fVU5;N@-4d@a/&>A\W^;^/_+P=@
8(gC@T@U7c=/dNAE)]df;KcB8SHA-8cGYDT9gdW:JgC\50^_+6B=9@cJALHZ>R?:
VIg,&VX5^#H/H-1#_@FI>Ba(PS_&XOH=\_UT3E^MT#^A5=\UY\?ROLd#,\=6C6]1
bg5eO.S0_@N5GT5UV4>?C2<Q5+aOS]A;22=?/(?G7:B(C@JCAB(Na],>\e>//1A0
N:8S(CUP:;92+e\&P(VFK>C?cNZXVVW79::93GH;>W^7A90?g/_4bPD?QEaUEQ:]
T<GB-O+TWE5SG4JG^a?c<96.eI6LP?I^;F_M,VY#;J6gH[+57VQ=0JAU^RBIU-CG
@#bI;^R#dGZ^D<3e<8[:7@8K6)^YXMMc5G]AT7X#5?B4XQPUeF5/V(+//O4]L>U^
-#H[[<R_(@2()@c886AZ_^V0=I#D2+cC(^:C^geGI?E(#4GZVGYGa+Wf;GK3ZZDF
35^NX_9JM2CQ##)9C-MJaM[&KH#Iae&;)..WTY0MFGZ1PdN^P&cYSCGZMKTBd,DC
.S(Q?P1Y:TN3C,]5dAcVODeM1S+6.>S[f,)a_9:MK_=KKe]-Eg?,T86-4BH31/JA
?Y17-.>HP>N-EBgA?+]GR>;f7R;OFKE,\RC:)O2F)5,E[.1S2C/G6PPcHXI1N-G>
L#4;^3T3J-T+8D+4MVPIDX\>7.S.Z)[;fJWVA\Y]J8McNf0+MDNS:.8)a(=TN25-
cREG63F/)IKEQM-96FdD\3H7T+WQU)8RHc/R,2T:F5XV5_)SSgGHDM,P-?Q@[H,U
6CL)+G7=PV;W:[-M.XU=9U[a\PTN4/7X9a\VQ8\WHYV,O2d&NbfYQ=Uaf\OQgYb9
#OfZ8(VQHR_dKa#aU/:>g5fTJfP3Ic]cEL1@:VA6J[b>?<>aF=d+ZG&d(W\3+/ZT
b=\G+<KI>QIYU?40g[??L?VSe:@BC]XaZ.-(Ng]\1-(8aOfDR^9@N3cIbRP^e9eX
ERS(>_d6YEPe<?783cRdD9+@Vc6gL+=#EQZC?QRecLW(=\&IT\\M7<eI?0dS?A@6
-O?62eK5T5f8^R-K>;,AEcSZeG]PBe_:2+_MT.^L#-.g^&\T2W3OaH/5G.2K.#9B
\)03V\EXMA#,aZT&=507Zc[@T#]>>,&SP^ca]g7KEJ1VJ39GO6,ZK:=K,&X]2,^&
Q8^?cY@A07f]CBgTB9e03d.V.1OD5a7-@A(Xf7JWSZ8OU\(\7?fcdMHS5c0+5VDQ
#,B@,\AGWfZ7He,dO:T-UQ6(PDU7T8Y]aS<EG10];O6dK]F08<((3Z[c9YbOJJU.
UC\];?VKgI>T+_Pb7R0f+NDC2GXH#(<Z/0)7I,8FJd_9X#O=VR@W221-=:8#XP;B
<d01Pe=Q<F3#[#</+,_KUNTbNS52I#^/,[f9P2>YYeFKUQ/D14Kg&O;E+[DNFZ+0
[)MDN#(-T9P:bF8)7g9.GANKF>[b:MX0fK;S]Te^eeg<e1-Z/.FL#WOfg&..S&8W
a0NF2PB\>)04H\6RPf\R/H-#?I/JR.Z)RB?b:\^9BJX(;+?g_ZUd-/cga8]=/^#<
L4//W5b1c&JB+Z6A5=CPW4H=(^SF\;,aB9Me)?+,:N(CEXGgJg=;b2/[<.7BS7gY
4c;5,<#O<HVFCg-7KANY?8A9ROF]JSXe(:OXIM9NL\N9OO7=cRGZ1F;PB\.6?J4X
Oa8P(QUF8^E;a&SaYW)D<3>-Wg]c_D?F.X^8_.BZ/MF4H0\^:\X]J6S6@ZUF)a(^
2A2^&^;)T_NT/LAP8aaK/[gU@:SRe@.V4IG_LG.\?10I+7T9[1-Kd8R#H,4OF>BI
bdD1,144??2<^W(VJ2&0_(NUU\d)g5OKCV72IfID]7#6Y;\4/>67KE&XaTYVT]f+
fMWba;9(c\G+JHSaQ_SBH_aZ,3F[>]U)1<RJ5N6+XSE1EK2^?Jgdd[\BT243-_26
P;X6&edcNVOeLM1,/KJ&PY,Cd9(>FQb0a64(3\D\^S[(.O4)NNP\=;I;aU?Yc\<-
\_^.Z[K_OB:<54P?SAYHc,:dKH6=Xb-,E+J9&DD;5T0HAYWN9Zb>QOKDP@I1J__]
_Of9E5WR]7K3X+YRVZ1MN]LDRWDANC-UYbD:#K6UA2ZIB]RYW=GMeK=-XB4HfT4)
_^7T@8^IQ^0).7(Pc2AHbO(Le/XWg5Mb7d#6<E##Ne2b,b>5V:]#Q)9S-=SgXaV,
KY.0]0X_>]?f^+E+#^LRgM7WfFHX3[.-,4S<=.K,7Z]&WQ?>SAD5>b_]^P/M&BEP
0DU,:NI^[AOE-[RT]T:3P/)Y_18&AQ<U,&3INDW/ed,B):gd7MCYX=(@F)VK<M_\
dC+>6b)#;^KR=Dc2C@<.]YCDZBS0U#;&Uf.B-T0^2-5>>;F/gM9-NV_G?ZD4dcV(
B6@6^:dUBbH26V0N]^,3MZ2<(.20?\V<#CB=?/]MCCJ/J.RU&O\:SDcNeWL3M+^7
#c=-BgXgO#)3e8]f\8bgEPfLJ@(<H/9LFN?(4&E5@f_?Gf,faZ01HKX/OQ\>2[V)
gM6c,92e,-TNPQPW=PU>La[&EUL5I?4<e)^U)8/(7EXNQ5/9W&JCYOG^NEK)</J8
6F/X.\Dg>3F2b,eFF6:OPR5D,V:UAX>O?^B?[QdB#G2e25_](\XIVT12La@[AN0\
VL[&\XF;RY_PXXZc1=aM(LWQf:W5SPI[Fgdf[B1;C?9gB_C?_YH_6+a=SPR;.H8;
71b^0KDLJ,:_(<^b(3QOJ0dHTEZRcEdN@F/Mg)5:I8a-:@1G^0GYBefL]FZV0cO9
3E<c6?]f0#BA/-1._/[K]\Rc-Yc5+O7aEY;RHC&.4#X5+dKGDR?L1T45=MA#1D1=
0QgCPE10&e6ZQEV<L-a>K#\WOL8]B<\L^-=6MO931K0gb\R<LT&g,Re;N)-&SUcF
V1&/_:?:(E]a1S\4^2:C1V1JY->;:;F)45[D<@#J.?[C9)(3U]CER\&I]Yg.>X#A
[F\d+d-W)).[.LW,Z?:HQQ]FWT:4a\9L,R-8^DfM7IPe98[[?-^C8b,>9)]ISeSZ
-],.&)X6S&CAaW>#7L2ASS7@Xc)UBX_E3=0c1@82ZS#CYA<YEUDH.OcA]IO9A9(:
&+#^AOb1U.UdBDfdA^/VAAL&1=DSI3EEfOUUaA[SR1bB4=[O&[,A53.<=6U(761-
^0?d^P7:?;aeV?]NZd+:01(<Y44&Y]A(a-D\./<63H#0f;Q3ZLc=Y&1EefSJCY(&
-XF^_-DJW:RY<H<3fW9Kdbgc&K5<XMXX(+ZR=IZJE^a+cMFCbYFZQ3B3KPe#ZO0/
(>&SdM,,=]_:.<gPg/+(:(FG7g:WY)WK(;26((I,7Tg4;=:1A<MLJ2VJP7.P]a?L
dD?SaeK(1KGa@CaXXcAHQ25d?NS4:S\<7A?O0]\<[gA-M4H8RVRQN26GWfH@XbEI
gR&JYNJUENMN8c+0#Y<7/;0Z@NDfe\-,5/1=,2@^Gc:fAd&F@E+Nf6Fb3I7:>MC1
R3e2O7_+407(I4B;cMa[_Z/Sg2UD:b2b.T7LB@;N?D>;S,Y7/fH5SH\e#RHS^8T#
=?T2?5)=,(OBN:BVG_T+D@1J:U46gGf\]6]4VgOdTD;2:G,FRB;@0fZ9>\_SJ[D5
3OM4f:?IL/\+_6(;?/8YTG#/(<N^=-S_:1V@S)6TGcY[KJQ&Z8LSSYT.?a]6Cf;,
g&+IUA+X2LB_&6^,OKW9D95K:b[QW7VT5eW?GN1V-/\aP=-V23??+>I^URTJA/3)
8Z/ENG@?O/]OGS4cEf2NYY(-(N@LcWN720,]4M)VOeT_H=:D:][XB.2QAPdX?7@)
+;(DP\I/]d2EH/fSVZ8)\)b174ZLAf()H]M]S)cCD:TAd/2+fD9eYbG6aP(2J/#)
AHUXT;++IA&ZV,)O6->UBbB,XH;Y.H_>9cE41-5VX=be5S=-7YT;T)ZabM+0#HE2
<;[gD:d?(5>#Fa]ZH_G[?BPUPBD/HZ]VCJ6_a;MK0N>V/[W9.KTONL8N(.aYJDFU
F10Wb>ac;_(EL8P8RW=.gg38Ie]2L(Ha8BGG5)FHJEd\1J^AXGgN>8PAYW&4[[\]
98(TP9_6T1QafJ@=IFK@\\3E3-D._UT4-1EH61/6O<M#]9#50cPZSc[3/WF-LKJC
5&NP:FD(:78=FM9^Q.Zc^#+QbFNFN9DB?4H,YdJ#MYg0ZXFYOL09\^#0@f?6g&M]
2e[B2O9fD5;gDgEZ[/,-;GS]DC@9H,IUAXVd[VSG/C4HbN9\a+O]1\RGF7JJ/d22
F_,OR;10&T;Bg,-UTRITcb75Add@NZa-/5:00)a?7e=P:_R8=)ege^cfY#R2f_5)
0ed)9HLC07N4+bd+H?XWe/W1IN6+aO8.DCCgMf=@+[=7L5aR=?^(O90H)SE3Oa?Q
\L.aK_SHB[W-G]YB,VN;KC(#e4TdQ]K<?K=T#_6fP+)?&eL>(T.[JNGYSP2=_RFY
5/&?7c->E\4JE2/g5J_A#fEbd:L-fF9]E5O:O(J7T-AZ>KGX(Ie>I4.6[CF@R(fg
cJZHZI55aF2G)Y&KZ7W3EKdJBYe55557WT?-EB]S]4+1adfW\#R&900f+?DJ6CIe
R)1bNLPCW=ZX0OSB3/P+H1f4XU<fP;Z/2bC^EV\,=R>[U,;9[WPI\,3-?K<]CXZ,
ZZ+ZC]X,82+F48@08C?COef^;S\HA1IFHA?8Ta,Rf2=B@3=NSJJRK8K^EbA_RP07
N+-L.\^K(B<D##:a>-\(1:2)1T5T/a=LY4#K/&0OGE11;8NF2:CcPE/Tb>C>K1JA
WBJ75eK6RV,&2EMc<3Q#&S;Z91W27O3&T@Z;KISM\E]gA?,;>:+d(C(_TAP&1FP^
[5(,KQ\RXY_7DZK)0f[C7+aR)NT9A=bcY=>+A8a^SZAFSHGA6OIT6f:_.fR3(DFD
eSf6FFaHVM7K957H6,P\S_FfgV1I?KeaV>]cRB>?e?bEKTTK=>,E8Y<_I@Lg,Q4M
F3SQ4U;f.#X&/E>O(Q3R=Ee;AW\(^-F@2CfCb_;C::R>L5.7:3DG2W\^Y5V:[Pef
PPE-#67Y_LE,2gdd_c#1;dgNSaBLMCDC\Ia8]N#aC=&<a)V,-Z:[J2S[WCdeE<YL
5:d\O_e]?0:8OK<DKb+f_E?)XTC8)C1-K([OH:R?]C-WLdJGg@>2(+b)a=@cW930
F6afJZH/E[Z:U4(#IFM_H<XKJ:&LaIKR]M9;dUIF]J\L0VF--AV,:)I6fZY]Y&[a
eCaEXL93>[VeV]4H2]cD\+\7^?_#3SI>#IUOBTg=/E7DdH]P@.02]=>-91H(<2CH
8+BV>SQe8bDe>6g:Z=KL2/??&7HYYc@YN-N_aef.#^/&W]fSR-EH8\H+NBc@>/-A
)f:=R2aRQ+Y=5TdaecZI).MV6QC)0(.Jb@&7>\^N3Ub3P[Q9.@=\I;AF2P_d\E,c
0S9e]>e-B=d\1I[V^+T4]6(BQcKB/A,#+OE0-BW;-=d;^WKW8_cLEKcHXIQ2;Q0Q
K3:(g2^Z1b@U\GYS3=fg6:4KCW()fgGFICR(eXZM+;<0#_2Q0>d\\IE3e8>/bJaY
RA)+D1U(52cL\G,\YG9@YeEF5?&NH+2_I/2W_)b17\Z3J^6Q.aJUM-:\=DK,DS#Y
^VL<)@G4=Zc1^2^;/8]U@5R83a:5#)/G>BQ&ZBD\PTg?d64UB_Y-?BW2L@5WNg@J
:X(0V2?RW(G.M<XWdS)C8K@2>][_^^AL?<&[b/U)D@MQ^ITg9A;E2X>->UDef(?:
H(f+aa]];^>3/>3VZRT(L)[7=b;4FV:0LdUZ+N?2QR<BF<W+WT\R&NOUIf,WCTN9
c@L++QdPGR24O1X\GLYKJ7#cV)=bf?,d#\0.5g5_KeLS]g:&C7aE#_(-MX(0_9RK
1JF/gTe+8DFf<E18RP@@]F>00#5M,HWK^6<,&8U-V,=>EMKPYcE\g:RTN:DI^)9N
7SX>;F56_0a/O1M2#I^JNU64[:Y;8fB@Sg[=_,VY7BDfH>,]IM;0NDM>U(_?XI2N
.9UIe/WNRWU1<RD\f3O3=cNSU,<)J)STdO7Q_TY@?f&J4:AZZ[EY@4\,>>7X[NJc
W3gUe-:[b8eaV[]-.5L/Aa+.Q>QL4J7.\)-4gPD^a;A>U+^A=AM>f-:+P:?OdfL)
K,(A27c>D/U^=54bQK/bP^:Wf>SNV<N>7P@aUa#04HfX6_@\Va)F8Fb-2K:L.K[<
NN=Z:GXOJX.<JC^99SL@3].QAfZYNMc#<<>LQCHaac0MNV/@c-I^&#d5)<44dO)T
(S&@eY0/LK4MV3b1Q5Q6;N#BB7=O4ZAIb+>WP,@Z)=BQ8Fg78:[R1V(UDbB01dXB
+FN2d]R]_.28Pf>_OWf>6S04[dHeg_[?&CS8CU&f-cKV43V0^fQWgJ/_^4#e_dV]
e;M#8/7JSYVW/,9]-J(U9DY3SI,L_gCP/Y273SB1:9G2EP[BdMI79ZgV@P4aRB&d
8;IFB.e7gE^Ag2&S9K/VHcO<d&\,.5M\UVI+=-S.Nc^=4G7[R2LP&dUB[PHXE;-M
MM_5.2C8BA+Y-JMN(6V;\H?5>S/5Y#?;:D3<D>]I6Mf3fe4UMT/8B2C(V(FQAEOQ
MF05+Ne/HS[2I#@^7gBeg66JGeeE@/OBD^:b#8adHA?F&1U5PdC&\cO=72/Vf:Gd
c;HIRE_3;+F?&J,>^73aITL-B@^KFdNFMNVI)PQg/L^-L>IWR#?d5GY+MJ#<a50.
W@gEC=ODg=WSTAIIZS>CDa=K?6d@M3d6)]I9:;(bO/R)E.CA:L(-I[Nc;B[>ZKJW
SP+G1T3T=W6OY2fe0JBA[M.(\&LcT,9=4ADBG&,b#?@S,:T+U7(L97(@SeJE-c=L
X0,XTO^XaVTaL@fAMJB&1)DP22?GU#S_Q8,Y4,5Ua3@[2=4/6/LXNEZ]#_#?[c1e
Ua;I1DD(+F:cQ2=9/T+B#)H>0P9&.M&E5FgFFfB5S8Zc)]dLJBQV,UL@?\\JI.dd
0NV2K#S9T(/PGfK@:>fL;e(K-gFQgM_=?J6_Ga)<@L4TE?[>fK.b4YKeTYVV-7\?
H<O6Bb9FSK?F=S]1:SfW=ROE&4[aKcW-PDbfH@YdAKUc(;;<R5QT#+HaXN^Ga?g0
e-Y<RCJ71U-]FG#VQ@RO+7BWS9:f[OEZLD_#4+@]]_4>K=X?9XfD;XQOO.;;L:9>
&B^B>g3A3gV7+37F#9?H_KLXLZP):V8#DPWDZeUG&PRA&_=CAgd^f^3QR9bQH0==
I0[SE)HCe]AKL<F7)E36QUcbO:6:+a,,b(<U5HA;,+D]W#[_I&-BFPBZLG6U\C@X
_<cZbMR/VGVLeH7[8G7HQWLNGT>fK\I5.SC)b+:B,_.DL8>=.=aY;+N0[+3M/;;c
=bN/T5H9Le?V(LEMg3)9A/AKT;P48.]E@K(f3-2TN?_OaZHb6;OQC,1f@HISCQ?#
DXEc-,\cG-V9)#,<BZ>.,JLTF=;bJO+VR[,-MQd7dE0MJD;S=(d9,.&VaN:=eVAE
HMXb)AL<_e79YY-gKU6LP_HEBV#U6@^BQ\86I[L/BG)9_cYCAS1?aJO9cO9<&d:W
>_150F<D603OZLB=gR^#29)Tb,5;)IFQ__>]U1U]=DR,gP>)J[:^76@F]C]Y5DC.
D:/gI8CJ?aB7GULPM.-3;&^)c-X3BMD(UHCbGgJ3&e+_FT_\#6Bf7W_[YgES-\-5
DgbHPS8&>;&>g/D#H+N+N]fYe&]C[DGPH7=CP9V3?V0/(PJ#6;KdMF7ffE/L8528
NQSIPBL)?>H5BN#^J-V5KV(9R0a.)+)Na)5@-^J^-2/H+UMMNSPD,EAgKcf&PM=I
KD@6CP0?W,4P=(1Sa]f4:4_>CNa3?RVaR0:7<C[<NKKcaeJ&H3e55[=bV2Y3B9JH
RST(/0G6R[57E(?GRP4L_g:=^U_eFX8OQVS4F_Q24;PA3PO/UMQ2[_6Z0Y6#IeR6
C?H1Y_FE.IMa/ND351<,d]FUCUD]cS3Eg73^FO73cd.#AfUC3CU^B?=[6JFT29U\
1HRL;8DC:>0O0ABZ2@V-0N7BL1(dU?033_BTf2O;JRK7WG1ZH>#>aFD-E>B_B863
B7WVAM5QT^)b#193S6JJBK>cfg-O&IUZHD=AQ),)4BRbZK>HO2J;8V62A)bUM?Q>
U3]76=PA&BG/dSK,#JeR[8FQYI4.GH_I8/AIHF,<f?95PbDH=M@X777BS@_0G6E3
<2+1XJNMU&_DeSb6]G#B+G>d7&WL;E[HP)AbP_@e[?AW0QB3[ZKE7c[])[?B+<GY
G3\]^V^;S/QBd^/.L/f0M)08gQJ=H.R?[G0fbe_3eCGag)<M0)MA4(9d]\e2(E@e
(IM9N7DY@(7WY,3b-/;8L=K\P1_ZQ3I^#EAM[3-K9dUbHa#/f\/add]<>H4T4Xc_
?TY?(N_E8&:1]4@O8^H.RC\.(+UX]/70HB.X@7#_=).PLN26WI]W=@E?Q0[>Z-Qg
f_WQ(afDJCKAY9S-A,Ab3dOQI4GEOKSBS^S;C;Q.[b&[>W1#dRX[D=+W],]&R[_D
&S<T>=B9aYCMTaDYN,&Y4.g&+Od/V=7;IO6)FT08SQV)[-9EE#>REQ?=?TeM+/90
9T0QbQ,=>BB+]L#:T-Y/e2#SQ?Ng?..T[d5FPQ79_?Bcc6&IH,#=c-be2:>)6LKP
]OWPf.0XCH#OaWP0:DRNM0S4NWKL)F^:6DUHI6cAf?/\F<;?4_K[PTQ)0ERXgH;A
>g[Fe7Q8IgVRY38=2d<CeBD-Rdg+eI5Y6..CHGD>_4BSTgEGb1e(V,WAWU\_E>K^
VY^#XZ:?MP/4&NNA5cPLd/b(^?I>85K@9@G9-UP3,[4Yb:3#:H:gc=>OQ(^EW])/
A._0Wf@H<+Ne>NMG2666(=[]X=G<S\g9.HEN7]MU;>XCIH0#+SFBVYBIc;HcHSV/
ID<84OHWNfE-;ga4L:>I6M+Jf8,gZ;IdaG+LcXCg>7MDE^EJ(9E5>=>?S2;WRVIV
TI+cJ]PDB3/)\AfT:Ce:->e08\D#BVF-2948dLMc>O34JR,6@9-4_ITeHF)33<eZ
Xd,Z4.FZ&Q8a9NX2\2HB_VL.31SG(cQe]OX8T4gXGS/])3IeXI8,[U8dA50Z+Pc0
9=;5AZ:?Mc=SA2Xb,(;aNg>EZgb+(M;(I,;-)UV:V9&IV^TT@W1)8X;5b-/;M#6c
A=A6ODHc?8.I1[OHL979>()X>UVN42GKQGCC?2NQ-CMDH7PU8RaH6aIW29fB&&\7
>\?OF8cM84<[cPSGIc^IEf/-OKL2c_fT#KIVaPZRYdZ-f_U49F:CXA)BR>),O:4I
)3g#VYQ[(;HOg;F:/DJ8+)K\GW[-Y66,N4]3I2NEXeA=2LL=29Ra/[SU6K=P(,6_
Fgg@R0FA\KfbK=0(=b-S(Kc]ZH>,6Z\:1<YF=b_S(_:0M?aO[)C?f3AgDe&.@0?0
ID9TBI8KO\1TA&ScK+f[;ce-ZO9K]15>L_fJ.-,dILU<74@[/UBTYK#]/d1#A61C
HeF+L^JDb)TG7SN]6S2_b)WK(US]c4f=QPL,GE><U0;O&_f^=BEd@((Uc<C=0_TB
SVFc60+HVLUT[S);VCeQ&-07ZIHT7_ZZL7(2b^dJPTLg0:V(DV^HO(.WW/W;MT5d
a(GXUd;23LX5cW\S7@XV]@\4,gJU#^?G(WTKCQ.QOVL(aI>OG14&f:-T4VA2fd>?
DQa(>dBBYV</KaEeU?d=8NSG5D?FDXQ24M@#CSU;T3HaIR7)DIHDV+b._J#F-/B,
d]Yd:bI(J]?G9\b2NV8KDFU&7^;0_-2f+A@=_\f-0&.aEOV:d1:;\^58MT?Q\=Wf
=UcX?E5R0MQFT#08A[]-fREf#M:JBFH6QbP<B?0[LaA<<fJ9KVcP4Vde-1^7#S^O
?,5IJ&3=cB]]+<Yg#;/a;HXSA5&KA6,L4=fe36L=/7_Fb401g\&\[F2SMK#;TJ;B
O_eeg,ZdF2>J.?UfCc0@gH0\GJNVW+=M])b,[9Kf^,\O<9=VJ40F.G&]#BfF)G3/
MUUAdJ.7Ud]DK_bMCa-We#NP4(RKP^/_;:GW?OBL7^=_+5(VYLJ]NB9O0Q(MES4a
-MZ4+_L3@ef#R=?bFOg4#44FL705/cDaJNG26I-R4^:CIBI?Mg_Z\LW0YLJ_eTCF
+_;(CZ_K283IVS9/\WN>F/8_M-=\UAQ[<FTX.<b@W7P08WU\3:=U<V7>E)3Z)\#0
O,gZMYf=OObDd3g;73\-FO/X@ROV#L:?)O/&22).NPaC8B^>QN5/U0&-4X/FPbS@
QCbGFgaS518Q7gRE9E0(HW.:EXb0[I7+H2JU:25MRE)_-=dMDH&f-ZM/7)-^&e7J
)d899(3R2]/;SCSQcA^V,I^bf4CGQ?)gC^G;T^HY=R[7aWJ8&;>92CN&SB@:?M\,
BOG2-=B]:XT;>X300M;3fK4W&^FYQ\S_7aJ&;8M@N8D42V@A3]QE<)4U<IVL\3W_
X,LYL^H&<_54g&IKa[L+fG]AceOE2E?9a_[4ac52K?]4[]2@AaTRRD@77DUX1,0a
J@=IX7WeUa<E>\TAe4#DbDY3\B62LQgd>^16.[-]Db9^-,ZW[ZU4@KNfeF+V9&V[
W<\?/@Q(dZT@X59K5IOVL)X5^^/RZV-^8=;<e1F<R,;JKCS=Z=c),43#;,R2UR\5
M=Dc)EMD2e\669[WSAU4BIWZM@]J8)9g[-^+<,2QPc-L;#e9CG?D+#MdXeUKJKWM
FH0+Y:^QWEaGB]H.NUa78L>P1WX5cS+d<011AYJ@dEVQ)4PMb).K_1S_JTBX&6TP
><9QN]NDeeS_PbDKE&=KT?LXS3YC,=7CAVB80@c3Ob7]S,NKYS54MOFfF<#<G\?O
[QSFV./gG,NV+R\8-[K]0XZ59(^4#T<1164L5FH=d&GS6VMHF0:2.CL0a>+agAe#
OTf/N;gFZ3^:AY>D1b?Qba]).6ZF#e,Jg-JHCVD\B/^5G?c_^\_>b+([6TQ<Z8EV
+W6PfII^#_@=@F=c/P\eg89SR,9cER[A8LB90ZRICa.3d>c/)04]c>;RXcSR\Y6c
&L@#.LG,,S[?ObfHSg0]N#4I=\V.7[PXH=0)9K:9I64e0g@<G2+c^?3V+Y;Lc5R>
:-N.D1Z>T2TROXBMJ6BCf9\[X9aQ(/7I^WB6L17Z9c?-/?fK<)?OKS;P^2,Md/A#
21V1Ga09@XJ1<RMbVJ(..22];Rf:A,SBc(a/(#P\?[UD:2_/@W60-&\CA>X]^[(P
YTA?.FU/]3214?Q8,G[8I0,aA69+XgVF3MWAB;BBBZ14LYA#_3agfU[NWcXZA?Y.
69)cZ:OM#aA8AW:e>T-CY@.Q(U#JA9.^_JJQ-^IaG]9?9Y/V]K8](,-Y^fG2BA>Q
ZY@dY/67MBH6X:FR6bLL)).f6Fgg<4BM7eSX2?6K8<cGLW_AIRXeH.,VR,dKSJLE
HZX>a_WK=aPNL^8XQ#0:TXQMHX2F8,_c;_G1+8cdaW46V/)U2JQ:XEJbg[b_QJYZ
fI)HG7.,2aK7QZb0G?8]D=5gM4@\=Da_NRV<:2OFcB8/9=.(a=+I;4P,=L:,T]7H
8KJLfPdVJ@81H(_;D:BUQ.gWL8E@2;,A<^I3QgE5e..;OD+/+Q.?QN(4(=B347SS
\ZXGa9.g^0Uf1E6;b=/KWNK/F)[KML.-#4(-=\Y5d1;-HL<EAM>Ta#RK<fF>?0Y&
D3(FX,&.,dVFR^G3O(-Z,#c9T/\SF,GbRV3\#c.aM:U\&#7gbN#]Tc^cfF&47SW:
9FeWc1_GEY\3\)0E1))QKH/H._<5[CIgS]/Z)[M/U-6<#;P_<6b9PgVUUULZV17]
ULBfSa/-G<8_9U--T4R&.dKT.K:0]e[PUKGbTM>YE)GF:UAFKC\_F@:/BSab#9MI
UI78b+#KQeC]R1D;0J^c=eAY=7I86>#J/SGDE-=>+X\XJD@g4(]5XHT(\_/\PQVd
A\K8B6CV_Y)^=V5R+?^3<P.8].2/CH8MXAB4=,2fB/IF^P&G)4=:S?CE=43-Q.@C
Bg5>(46+VO0&41G/0>PXX(L[T;UYf8MQPIB=a>1>QNdBS^M+94Q0@,bYV/,P4RRI
?^Vg+1NX,Kc/V(O-IY65+:@S7Y1^cdc_T1TF/\f&J26Ne_eC]c.46P3F&XHZ5]AA
C6]d8Cf4S[AVQ96\<f<Z/FA.8ffaa(N.V\/10Y.B=N)2IQ-^)(]eX^>6;?FADOIP
>R^]Se0K;.Z]bI^OXHFR#FL3X[Z2dNKCZP<bREA&?<R=>6-9II#g9R(;@M<)OE:L
S<Y][7B_NP-HG)LG_8)7QJePX^_,bHf:ZET?>?+L\dRE^\_e7>P<fa9FPDRP:)gG
/@L3LX;BDF?^:HM^0]AW2I?-F.K9FY2fRLJ.B&MT0[Z5E6)BJa.RVR)>;EY@FF73
0;4@3(A\)]I,/B,aC=_D19TbFeN&fSF,Y2Y]X#\KW&(g>TP:/,cB7J..[e7L)V5Q
^cFf@3<OC.)M_0=>bI_@WCEb6@N&F?Z(4I>ef+.);@-VEHdGBSZ9cU[78gK.g62S
M)33[2<+4P7:Wag=0=#Fcc5cV0]8ZI1D?&JQ2aS.F?.cQ]U0:<YGNL#Z#eMC8:HT
B5MdDIP()J^QB)+BJXD&B<5f3e5@2.CK3]\.\Y8IB&)(/_9+VAN>YN,,Q=\=<G-<
,BX/?/,4E,K(<9D0_0NHd\B?EJ7e=>f?5/aWO-cdgJ]R+A9c/C8DdgeZgJa8?c4S
:SYgcEKc:3e(=?RR#.GR?#g2f]&_,b\P1PX.](U.6)&CC&F^Ug7&H27-c#E3+V9.
[ffX1O)L1_PaG-KDO7CR3-Pd-_TT3#K>TVK41V[8>_J-X0]5(:\1_+g]FV/QQ]PX
VT<>;Ne>Y\d,X#8[<D+(9F3.Ra/V)^E-=A0Q(@G,P.(8g08GY7U+(^JFY<?e-2PY
f-<N&,9?2^,]Q=&83YG[B)G\XSObA:EH6RR1&.e,DQA;JVLb4FgU=\5IZ_K[g,UM
5:]9J/WV-#7T5=UEFX\]?5@VO(-HME\_)79LaU.7:KYU(R2?VVPI0cC+1=2EcMSP
P#\)RDXL5K342RU9T0fNe;?LW&Qb+@)eU[fJ\H.+bYMRT#C5Z3K#1,]IDY(Q1H^/
T/\I1eQdEWA3Cd#:J5-Of7^?(>8\\7KDdMEK+0&O0[]=g1YB4ORA#T,++W+;IZKc
40?>\=3G85C+T)K@Y>(>=6HQ1U2,-Ta61VTV@9\M&H>^5@afVA6/GO9E)bZG)Vd^
BYfV6TT&D[bb:-19a-B>\1Ve3BIK5&P)O;#bSO?YLHP8IKVZc6R4-ZeWVCI,4R.)
0A)\+</-#C+MT0fG><X=)M5Ya)]4NJ3M&ZMd0_3A1?>9WC#P]RK0<IA.QF(f=R&R
[Re)d.f+@L5f7d.^IgAKAC;/g==1D#QRZN4:R+UW;L_b(\.&.cKNVc9.<WK9TK+Z
RAQQ:O\bQfLCd2Z&B?1T4WRV[.X+,W.C&b\/B]J_F;I&TaTa01Md^5gWEJHc)N/7
W9c\fN-d-d)OZ);/c?-g]L5HSW7KH:KE.db\H6f[<_1cN+X5_2-,.#L9a0<;##JH
dV4-/X-:.P&]?eZ<A,IAc(LZ8f.A=LX4>&O[ZVWM\XT7.,MM@:1Z;Rd4+AcJ1>Ja
O1XTa^;X@,P:(-FaO(TADH&#2gES1WFAI&:N@(_@[aO#(];]^DQJ/7X56]H>#,KY
.:A,O)+YXD#OX8D6J;H>\SH-NTRO):HRMLZ40,:-8g+4,_]OR#g:Gd-Te]cP,=CO
-F@,Ja46:D\Bf#eI=D#Z.T_+XP)XbIZbP8+W/d@=&\5.7M164:A]\]aT+fZ3U0[Z
VC@3c:=)PG,95.)dK.b7TY8bV(\C[]0f;f_-6#U3ODM)KB3O233SLD<9dNY<Kb5T
RQ0DZF+c&BM(HIMCN(#Oe4b@g,(=P>EN18ROJFB=1YS9BRP]3=]Y[.0L:>[=Zb38
@>Qeb;fHXF@O-,@3+=M^bQF5g+?J^/RFJ&A]IE<U]>SRGHTE^^8=CGCH2EU4T&Ag
9fDb>G&JQKFgP?=V=M];&eEI+1WbaHAZQ0;NE@U#/74O[&VA2N)OO+5GK;Y-H<B9
U412>Hg1+_<I6T,B,[;&gM;7/BTY/;5e6\H4]:LeE(e(XUD<PNHL1O:^PPVDA0(G
80^9c7YgKdKS<X2eHagdXHLIYaB\E#4EBP0(>N17#(5#TY_]J[5gXBLe2HI+fE?f
>d#3(S#(g,Ea6-=@=575L94Q2><eX?_?P-#I,0XU1W[M17N/+da4N<gQEAec>BE]
JRcC+O-M\#cJ9_H+(F6,ZSIRT@bcc15@?G)7@M8R^&7c4,DaPK;e>;?gD\(Z]DT]
ZEIWNW,cT;)eX?<1)F5-S)\EW#+TPEe?b2]<c[,@_O0ECMC;0da_S#:b7:Ec:6I2
1&d7<gYMPLD3G,Ha8[VJb/FWRG8E(//EEQ6WbI3R@(V0(Z,SeTIOg4.O_c.C8.VZ
H1.eFAG2[-I[-;?C@PGOPYLJ#[OXL/]J48=T5G]-/EG=dG?\7#;TcT_GaJNSB=ag
M#M)+#>A]MRg,9E=,S99U.<.8faSY/KZNCef<4;(1,S>E489b+5KRIVK6RgdLE.Y
)8_&=QX#X)WZ8#Pf&e\S[Y1NRZ3U?\_4VaeW-+]59ee^MU[fX/8@If50f?PB<BSE
0R;7^,cL^D;@X(PD.OH4N,#FU\SgeR&4(;U,9;dXd#\Oa50BdCNf=LZMP)HbFU.V
T>W2XN/&#QLCDF4(L2C]FU0+TKCK\Q[9NB>f/=SB=.bJZ<B90IH[60&S@S+7]S61
Q]P@[Q(_BdLa.N6,V1Y>PF6YJA<N^F:&7FN\IOb]9/7Kc?5D8W8cfb3e[+[EO]X]
1BEW?)X&>G:.T#g7GCVB1g9/&Rd,]Q@+BX<Ea3[,4aB6ca.aN9cZd\cVe+]2O#H:
IR5HeNg+MQQ]NcT1\c67g/RL4_X\Z\bM1fg\&KH2<-A:AGM.IMfeAO-/M>Hc2LZe
[SK.C9+L]RX\#D)B5BN>^c1b((g+dag)-B.W&?d7U6>DE4^UWA>2BS7e></<<&NN
Y;GQ0=bX^5g++20)01.-V2C=SFCW+^34==g)C\+8H0+XP:^a@5&Y^QPRGKUA2DcU
K<9KPA.e]O6/1U:CbO3HS;WB.=J?12Dfc&3WPNTe58BJX0H\0[+1E.U;He5])227
/&KT0,FXC=Kfa\QQ9QHA.OZdV3@aW/C/3:WWE3G6<WD/>PMUa,.B:NO)W:I)I_UTR$
`endprotected

//----------------------------------------------------------------------------
`protected
g6XN];&D^+-)Ag,7-GfXV5aL:A/.XSDVH-.ON;E/_YEa5YPCaB/N7)?WU(]V;W&O
V8)9Y33:5T;X3.g;)bJ0VCaL3$
`endprotected



//vcs_lic_vip_protect
  `protected
SJfJI^aL4LW6eUCSF\5]G,gL:MYe^8J<\(I26V83J<_P70XAB>8S)(X7P+LD6#OC
9]@05,;YW&\^S]X-Y;-X5,gI88,9?2C;b4EeAXd/AD;JQ@:](>P-VH\]b(BCBf?D
7QTDQ@]#5^E38JK:(gYRFg<fDVL(]:Q6gN;b,783A;H?3@_8>b]77SeLV9I&6H^0
+(\4Z39\M0ASX.,PXbe-Y[>K0/VDFQZ+SZY/OYH]]RT6U:&CU+.EQMf[BZ0]^FTD
g^@HB9C]^SKN[/IE8?3^2^=(929+3AaUHE(ZSXE9>:C^EU1L<UBBM(JgT3_97MOW
N:N0/B?DYE#Tb6C;>f=1/]4E:=3Y?:eGY>eR.)PDE21W_DEc,6^Af<]B\Q_2,DN[
.a^8+?HVOGg/0-b6Wa2H9RX)FM?e>.7T)2Y-N7=ZWA8,^YQ84F\N^Y34)VeAWD[+
Q>D]_:@=@XB^A06\4):Q@;:P(=&CPT9N_]]VL/)XO>UH@Y3@,2I]@a3_IcWR9=[K
J@Tb#Z1V@5:@gg65RKZL(9VU=PQK_3LQ&Y2@KG+@eO9d,MV_[GgH@RR#O3)XcQg0
V@e4S:(54aO>>AL>EU8?@Y9PA1@dUBQBJ>@7D@DMM#4SAH6]-MKF\YBP?4UEO/4W
Y/A=;aY42EM6PWP1@Z>3&J&@#)L:/4W6I@C]O\SO6]9@>PH+@fO(P9Y^.ZX@1/K/
@+TWOIC4WO-9(&WB2]MN-Y06Qc?ACC,TDKH37<X_fRcQ#eL[YfE#LE<7+=E,#39Y
WI:b6166B[OI-Ed)8fE?dVR?W]T=8(2AQL,2G:+8YR(VJ>F1&RTEJ:GAFHHH8W_2
0C-fH<])6G>PPGR9M:)CfcKH..g54@86F\>U7TYb#2KJKM;H5/5(3bJET1#+/ENX
>80;#9cg=V0J\@ULVPH3b[d+BT]=&f,KH,X1RSY=^]@QH9;\?/HGDb3G)WE^#@Sf
;?U>OG5Q+^N8.+,&XCM^Ha;[gH+_0E=0X2=_+6bZ(PX:L49+AZg#eBB)&&#AK-:\
H[I<7?;LP(M&e[)I9LOWSB=5:A/AI3/B/T#10DSFS7A\Dc@gW1X0dPYTF3g&aNBa
GY>cN-B=_DCZ<BDFF18T-YSPH;MS/^K<)D:7E/G]6CZR3^b7>f1;?ZIg1-R,DMZK
#fQ5>YffU9g_W9=(32C+,=Ne>G<64IX:PB+eJa.9XXU<QH[5(6NMaZg30/W@48W<
E[A9R-ILDa#D/XW6XbTcUEgAGOFec&O&gX>B9K1G/JVU\4,T-9>KXQGC1UQ/R)8H
G&OS\[aXVXF)c65TPC]CXDMH?78EaTN)7K>]ZN=(JM>R0EJEE)X\S6GJX6509\M5
N-[\_NGM/_Fd:\_)&C+(-E:#5(RZ0@0AP^IQc,B]S@C<1d&JB9cKCTc_J2N&;d(T
[T+c[J&I:gKcWJfE/YB_JQ47QIS+GWa85)?E4SG;L:UJ#J@gG>e:?0SFU,_>-3QK
FG?c>dWBIXYc;:NPS\S0JL2a6:cc&FdBFR:?I+_?MU=B>@UG4eLPJ;92,+><JY4_
A/IGCTG&]M#USWCF2GgMdUQ-SM)K)+X=:gFX;)7+.O=D-F_6>fPGL?TDJ[4:8.P]
I7AgS)F#<I7WdQ)YQS^PI<T#3O_P<6DJ9aM22/5JU_6+X==(T(_OOg-VQaH4-0P^
8.(J9.=GX+T;03)\RbR.ab+[N32&1I=3=3URC-d8=]1&D(\(C6R_T@S7F72Y+<?J
UCGP?T^[_]U+J^DV;+DY)HDb/G0_JA;Y@fb?ZO=Qd^NQcbO:_(dF_:dB5?_2E0<3
B==C8N<;>99:2:ZTAYMbUETC5^V&>gYOJb5E/=gE&KaXbBFG3c+FPJ19R6>MDQMT
XZeV/DeT?DS;YeOK#2dD./QgG#88MTF9H2XJWF2D9[-GRFDVbM1L797:SVJ9A0\=
&eFP0MfL[Q.>#WCM.]#8b.I=PC6K&a@AF)>P=\U=V[R6P9-bY(V-<+)W^GI98.M8
e/H,1B]^=:RZ_BBbG+2X>/S=E8e[[aT@VJRQ,g.T8#fX@[==O2Y5bH_D5R(EAILY
/-&V0bg9/De0Z3QM1dOfPGT+XUDKAa_?,PcWLd#-[RAD[ZNVcCI=,C4DZ6HTVK41
<:bR(?8fES]/gfFIR_bWcd\5[62KB-=F;HIae3[E/D81fOc0b,X4AHe+?:T^GfA^
\93UL3AF0?<,U_4=A=0Zb+41ZAJaQ^FUB>c<Y.2OVOT?DP#R5F].(C;9,#LCU.MZ
fG6>E5&>48_@KdWE69e6?:[YI9I8VXZ\(cBRSV7=-+.S.B\6UF77ZTRe5)_GN-\W
T1NZ[W)^EW5DMZUKeK@)Qf2_F-_OabU]TVT?0PO.E-=aCAB:(?NP(:SWNZAZMWBC
IbNS-<A1EZ>6QJFZC\)T7&_=cQ]CB;\1D,9K:7LV&&ff#[U=MeOb[Q\@&>De1b.)
g;5aa/XO&eMfg]#T8O\5-a]6F31F<N6_#>9^-b+UN<\:E(LKMNg]9C^_(;M.]dW_
<//3<SgP,Yaa_Pa\/4;BH:B<0WfdC92[F;993GY)&</-dMaG^;]6@QH.F6eS5.7f
fIZPQb_EMUXFXY#PK\YaB4]5^KM1P_2UFH2dBO)-V-fA8^9VN1WM0aGf8(Z@X&<Y
@&bMR?T:[MQ--II=bHf0eHI9727C.g?B4RTU2_;5I?bgG?d(<e>;/f:b.)^D&KO&
N5/4E)3V@.cM;;AM@-MWF.0bJI(1(F2c,2LcT?745=69;f7:VZGLNPGabS:3a[^@
2c;d[3)PdcWZ3ZGcR7V=J.+c2U7D0aBQGfIS]&M.c\_aZc2U49V6e5c2a+EKV)J>
SPK^EeO<UDIbP<1Kb1I6.ef4^^T.T@F^_=e7@3#Mg-K8)]@N[OBT:GTC[5(=PMTb
cY?G_<B<EBJ[[W1eZ1c^VKB[a1CBaUAYd()dW&O=Y#&UJ>7Nf-b0@D+WGNL[XNPG
c4,g>0_>BOfXaHL@#;+V_aV]C#bN]Rd^d^>aSFc=g+.e8e1B_CQF]ECbb2<<fW:M
:,A^5XUE]]&Y^BgF1?&d:N5f]3ZIK9\:H^SY6eM<TaP39@&TD_S][5?3?]e5^#5O
G<gPV=>F=/31dTU<\<PMNPUTDKVH+Fg)fQDA?-+-S0.QbGQ?:^;Df4JVb5=JEJ/I
VgbDgNFDaDBJ:S0M.c95+A/#\9R?YR8BK]#.0KdY-[b^]A_0F0II2Ef.YW>6W.a6
9fNeLS<+;+/)]PWGY,e:RRD2C__YTJdF2V3>,;\VKa9g;:_L#<V?>eR9AR-_&OgE
O[-K8\SP12.[O,,]P1@RT&:a2dFX+PDgVP;3/71F:ES7M_J^QN:8@1E:)XZRcYEG
ea:a.-#/DO7YJIOV3_G2KFEfSTfbV:.=Oa(M[V[Cf>,,b\6HFKK,?>&.\;;YG);@
e/FKU)7T-.96-cY?B5T.(A75-WC#G-adBZ?NEe\=\e\K6LL[QK__Lc\?S.b>29@e
c\-O]N02NgWE,L3]G;YES87:bI;gLI,DQPGcX0^QffBF86A0\8JI]AL[<VS8RRK/
bUUQ8-+X_F4d<?+gf15).O&d,CSG,b3[M>Ge:Ug2ePe\ULPXaJVPe;Re)d/2b7/M
J7.L_Z43HKJ[Kd8:>:8&aGTC9-Ea]FEVW);G[P38V(R1C\Xc\bN&\T&)/8.Va4WT
[9VT/ODR<V;ESVA/:b:-DPXC>)=Ob<AEY:Bd-@>[<DHFG9S+Hb7NJD<OQ+S=;F&R
B@O=-C.2\N3dXZN5LENTdDgSJ6f.>\g3T9:MV[)PX+7@J30/<LVY?7EK1CDQE0[Y
PC/T[1DZSEU;E:P.Me#FeFOge_bJ3M1.89,2\XUF149KPGWDIN,bT4Y6NLU8GYOG
X8#Na0XKH&\F24-R?D5G5)W<=@fQDKJ;10QU9G+S_b?F,C:1342KMI><gY/GZ3QC
5OJOe^1IeGE\Qec^\V&b9@S&+P[T+IJb[?;2UOe:-S)fAb5UCM#(b<3A,##:T.?G
N28(-&[X8ZHEbdR4PHL+18>1FC&TIPH<D5USaP\K3DH]Q^I#3M_;:=SOL4fG\;&-
<A4cMa50)e6YA4OMaQ3\cOQE>]@eT4g-He3?B]E>?g8S9B=O0+;/G>0V,0cdcN]@
X2+ggd6NX4)EH3db[J9(\14P9Y_d,T_O&(SV72,(4-f;<f/\86/DR@@.W_;,;):<
&V1Oa>eLHB;:g]IfZ0P[_R/JARcR#)CCQ@)V04a6EW68QL_YF8a-e)1>4@RP_+>E
d/X]60/:;Eb8#-V^+F^]?:QJV<T2AD>CB(;fXa9<.UW,.<?+:<_/2M[:ZZaM,/7D
]DGdHN(N(WR]WY6F66Q[C=R4VN)8c2HP[,[/Z/#(ccS5EK=NRD&G,M[_a5VW&>N9
VS4\?\8F8]MPV])E,d&(.?=aGeeC/eN=#P?=6caM?NW]d[U#g9Vd2aC57/c7(8H(
F4334/96<-AY.aSc6DB=\\AE>Cg2,O9KK=9JWW0:K0bGSf+5)71gMVf]a0/Q5IcB
[ON4G>RX=1_/-CWJ10A&M(L\:GWAGRHV>E]2JP:WL(98e^UYWg+?L#^Cb^91=HD3
f&+WEA>,J#9T6/49D^??HQ:,:d67,I5^:(FU>EWg6#?KaggbLMaOL/,0e29&9M)7
J&4G4([2/&D,I(P[BRfJE6S2Bc_JU.>dDe:J&4^O@9c]F]<;;Z<=&H0---+)OdJT
J;D:Xc;2]:8=ZR[1?I7#_;RdaU9.9LQ_.IR+2Q6],:WFZ)7;Q[7d\\d8POQ^-;:J
;D([2Z@BHA(59+S_F;dSW<.2N6B:9g1:<;TFHGC?KSMAWV[P#F(9P6(Q4TS92._1
>]YH)K>++S@=_6^MQc,?9)CG?7R-0.?g09.5LR?4cS@KU+W_=8@+B7bdWN?EF0X-
E.-.O]fR9a.=F#UdV/Wa_D:[_,)^N.g03<XT>7#E6_A[_f>0-2\W7,@(Wc4>g#&6
KbU8f?a-5L>[CPIO2gVf3Q\_P(^;bO/@4SG>G3WSWTV=eB&7gK7=)B7.ae,E5[[Q
M<,JDI8JI(/C^BA5H<CD\/3>ZFbDXe,J)<NFgO6fE&KLHB3CV]Fb&AQ#.f-9Fd3Z
9_AI5+O.]H_NV\>8+<02\=7(JL.A<9-GJ(\M<d8)R4CaM7<WUaC>4DfP&5M27JN+
FM9V80DNZc3dAHHYX0@3YQ_.<We=+JHa3)eYPf:CT.N7].CU6<4:>S5ISKJH&TO/
cgI3/SL-^TS;TCJIb>RC,J_U>@,PHK<:+9A?V)^;Fb/b_dRPI5b05];BGX^)S=g(
UUgU[<+R9g=>>_/EZPg#X,d_=#6>Vd+eKJ[Z7F[R-)Da4D6Lfac0^a=Q3ff[cF/-
afWIAGBZ2f]S:gZD5/W=H88AC)\Ie+\<&0N+Ld^(bc@)ZV8LM@?6:;6GP.SJ#/\a
H;8;#;&[Tb1eMLd:Dd&>31:SNBK-SOb/Y+Y(P7;EU.e&O9+,@+_R/E6)/>^g-PQF
L05ZJGB59O1G_#5M_KaM#VJg2;&WG5S-7T=,+)Ic_\K1).,J^JO/&?/#:5-II32>
:,R@c&F\B9SL^3UP)@HG\TOOe;fX_MI1<HIZXWCE@BFbXIfYZTFN.3&UIY54]JFg
(NS=+\6.B,;85?)7G/e=@(Q^XVcU=<e\^,W2[(N(d2ACRRNfRfRYTK@39S^e^8)5
E0P4U75J.gI[5gAg6=-9>Rd7PF)R\LB0IS4W\O>[H__,4Ub<5MNR.K=>cU.30@_/
FE9H&eL</UWbe=_RW+I59[,4NQ:ZOL?:(,98@3U+fQIB+aY-N1E8-L&VU/L>RRTQ
K8f1:;=0]HUJ#Z;B#7[K4;81OU)5,,-YX&^W]QC)NbPK/Z,629P:&WbQ6;C=/Pg0
g+\@]=4CV9.FZ0bACDbQV71)JT]^dDgR)_3<[6ZLO:dMP?-J>BEOZgMa[A&N]V[B
5_P(ZC.@PK8BHgMM,XNe+4+Vd_L=?-B_IXXg64_fTMXV26G<[eZ4-5TLP976(>NF
E9;=S886(CXe<#:C=)S:SX[C1Od-dS\B+PDH?aMSS,.(g4OYC\GDc3\dWYES#b19
J5]bJ4M4Qb)B\96BJ=7,M<_UD2NG#VTH]/LP3@P(B,,7K\I-G<2B4U=H=@W>YUEY
NAS[9f+<V.PQ=&,XW[Z[5W1M==_E-W#GFPUCHIRW-0T70M]OaEScUDS,LU9CeG@;
7_4]8:<b4KOLa3\/d?TS]MQ<+T&5U[MI&g1SbU)F<)e^<.G0g<Ud_?WLHVMH1B5@
9^T<1f8^H.>P-ZKfEb4H<eBFKC@,[^AL,ZRPS,12]ab(9CPe6?KF.>cUf0=4S2dY
c:[;F[](BJ;dZ=^3>9E7aD9)ZT:.b<-B=2;NGPUS6S?ZKDg6gBScN<HeFK4MO/#+
[FTb_Kd/fZG6c6V83YWK]2G@cVL.bAd@VTIX]JEGa+W>C@Ud+;f[CUc1@[_]3,Se
N?/0?=;-KFL(DS,^CDd.;:XePRPe9e;8OJ#)H?ZU:Df^+AG[4L<R9:H6#N<_9+YY
MgH]1fOQ;ORAR9\cJW.2I6KCVK]2@2,CO[2G4?b58<a?64PI7Y2Pd2e=1:f8UTF.
?.J4E95)7:G>FL+.7^^Of:]VV?A]]H_3FJ)P6Fe\L29\;>1?((D??/c1ea4QGOO(
_EF]0\[dJ.c;GfV./T:-<-&I9M^U:6YZc7C/&TC-X?B:^\L#9T9@U3a\D]OQ\5,7
-S3>B&=0eYV\;f^C:/)CH16aBO4cAMALgBe5+VZg;6gPOb8,(:=&[^^I_H^3bD8b
O)fRcbeN#1N?F9MF;3,XTc1\1FSd)+E2F_S+:;PA;3QdD]ONe?Y=8QY[e\2=>/P\
G?L>.8:gLEdV[dUTKGc1VJL2[A#+]g4H\/=YbaQ?\J/S:-RfYFeIgQU3bB<Aa+BK
0Wc=4268-1Af>S3+gZE6_1Z5A/EA-1];]X:8J3Y(AfI./f9>P@@eZK&#M\:U;62C
V0R14=-7g-MBZ&=7-EG=:X9D@V<;[M-Q-VcP4.LJ_ELI<P8][\QNS4<a;@UP#PQd
A;L959c<)1,?6NcS:+YQUW,2Y1W5)@?QAb]Y/aF3NDW6/B&FGMP&G]4H3EdH#EXT
-ECL4FD4:-?b=YJ]WMG)([ZB>9K3b@a)@C46[&A53]COcWGEQ6W7\00>bDRF+\:<
<F4E]AWR>B/[G:QT+<_d9:.CF05+>bEU2]FJ7ZT\e2JSB@3JJ7UTW.6<Vg=2cGI>
HOJPT]&9MAIB\gXbaEC2];\32AJSS_O@c@X1^OJQ+H&4U^PY\>B<]<]R6TLAgWNS
1&Y]9BWe^1)?Kg^J<3[-/-Y\IS/(;9];4IX=a6(#Fa#UcA1S&;E6/&D#1CfF[H:W
Kca9LD<&2<@&&I60WE4#GGS3^<7N;dO6>;1g#f28,VA:RGAW<H59+_^>1#R5-QYa
gKYE58L6e8KUfV,KQ/5V-Zg+4V?I5\D?gGc18T[\B#6c\1-+B:^HIW[Ue^&]a7a;
1C]-7+JX+/1?G\VBX&NFU_WH>ObXV9W@4)WZSII?B6fR==WG(P@?NJP#:+^Z]6)D
.La8T49639OUa^4bD_a4BYC1GIf#70EC4:d7Ab\fF<[Pb)P_C#BL^F63R;9P_NDD
3\aIRYCX-;:W[PQfcC#YM?PVAbCKGH.&>V>,acD1^C=AZFC,R_87])UKOQE;a]Q^
Z_7?KQCddSFF(S.4R].QR\=YdUM]3FFdT#a8F;PDNOOKaOJ3W@a4RcF4#AGDOb3X
=:J[cQPKfKgKK?XURXEc)KRXR0Vfc(Hb6,0>0KSG_0R5^XS;d>)E2^bBZT3E\FYS
=c\+O8-YDK&CVM8ZH[6KU(PQ&7=BY+BNAfF<8YZXAKXP=7+D0M^E:&+A),VB@,)&
TL#?,T24=R?,6?D<30NdU3gV/+C1>TQQ+V.4M-QC.X&/(V7e9:/FEK&/?Z6?4_F0
M(f+Bdbb2DY2Q)]9H:O\A+ONXN3]6(-Ea-H7AH<QCdK,GT0:Re[&aU&M-J=?EGIe
0<UXdV)6Vd^[..>f[W,IK\Ib^;^J3aI)L@0(->W?#<\A7SHc?RE&/#U4\2IbS7?L
H0:QGT#gUBX&&W0\/2bdHHBMSYOF?EEA#:-7MW;#:4c^H^A1GDbL2<AKJ-ST>8P=
Z^-4L?BM][Vg:146(MZ)HIVg12DCd@2LU7UI_dBTD2?RDG^M>I66;C^Xd<#R&L#[
]e:I7NUXg5g9OUKa@6&g/KR9@C-8UVECcX+a#,Y#91N2\8IAB:<.OVf=HJ_6XOY<
2/S^[/==a+><<94PAS?\d.&-eY2=;/TCb\_9HEE3>1@dgDbT/9HLI+;E>5:=Q^<=
E6gGSC[M\VTUUWQ0L^1M1c[+?K<HcKZ]3[cJ]?-QOSY5T>+-C6J8A,33f9e?Z&_g
E(7VELMZ37:6U&0#.Z.1Qf,Lb(@-AgMIC;6XH1.R:LG9O5)48#QWV=^ZZ55H_ed)
9gT=Y\U_R-;S,PA8MKBJb.V=C8ODS(?25dM.1D3+>YL]b3G^T@GOKM-F3+-#:L>6
T&?cQ<2gAdA,PK2)U1[#ZGeY-VDIZ<WIgHcKCd/d1;GfRX^VgJ38@8A(>&ZM(Oc#
a\\4@@>PCJ7,N+4TaKE2UW&>P_=>;aBCI07>B/J(WZ3aI&3^&613PZJfNGKd.g0V
4d>^<,g\,XF\62Y3ZP.HbJR53A?0YPIQLHVIV6KRXW>JTV_bT9S#;CZ.D@@DVA@X
O#=M9AYcS^gf6A])Z9ZJ,/8,Q4,-P)c:V;2DK)3F8HUIf/7/#/<?5bXY:BI1d0.3
R:ZUJHR-QRgYHF\T2W;?BSO)0X04:BE^Q0TT5&I=B35&F?F_FAZ59SV#>DO2,&1.
5&0>RcJ^1ILTQ/UP280UL&RV0H&Of:6FPcSWdbdaCKefReEP^:-41>ZbQ)=CN0>^
gcMNZ;>f+M<HW_9F=G@0E57E/98L-A)M-A,&>@MTAF(7.>(J].A4N&>]F?DfRaL#
B:2CF,A)L(1H8NG&9e,;3[D3X=0XP3cIRO+6(MA:&.W?8e4UP^Z)I6f_Zac)9X/I
TO_1SPc0>5+IIU^aCX>]N33YfWCE)9RV/3:TTgf^+gL.P)3fTM8RLFZMOa1PQ_M?
M.[<<?[7D[3X6\Q13NBJX<_9ISX/1/M^(QL[a>JY2gJ,P)4dI:JNcWS+TQVY_aQL
BfY6VES8+,E6+;?-NXWAIB^2]-\d)]1-ZLR5F^KH)aIGQgY6]?dUT7_&3Xg+2M5;
0ZJ^Y:PH2;bdcE958?JEa.9fQ5[2)ZB4U]T32X2QbQG@FX;(-A9[eG>Hf.PS_MY#
D,TR&4].1OQB+C&J9?QWI,0\4U9GbIN>.0.+L^gV,AUY]F>fR#Y<JJ5C.4CDEC:C
F51)@V;C2NI<YD?]V_3T5eb^2YA3.)?.(ZHIL<X18T1,HCb@@8c,aR_Z74M6gVGa
/)d:1[Gc?[MN,9f+;9/QE^FRJgZ4RQ;0>J,E24O0SCUfPY_49HM236_S\b4L<-M5
Zf.MBY/N-</JDJ/90\_FeA2N0&bXW]S3CPfJLE5<W;[S0Y=57XC6U+F-=d\I:3TZ
@BH>C2N<+GQ((1CdI3#B^S8I=/WW^,WNM^/GKTSf;9><M(D3fH,Jf=d&2g4FW3d(
4a9P7?e:)AH6C,Oc(d=XXGELGQa_geE;)V/S8M>#U@+FYf&F,aa?^M>e=c.+,bM]
7PMXXI9KgKS&,+(:V,A(,8TS]-[_NKcU-^DU?[<2abW<U9I-2cQ;4BHXEN_.Bf):
#^[<f#QU=S&8=.@C9dX3KOZSN07bAV12-2OUW#ab:#DeCLf8OJRIE[OI]b]cR-O9
PIP4,7]8FG>D^@KZHT)E<>]L30S)5g^O+Mf:ME01TTBgc;L(>,0>33SC-L,[X,XJ
&LL\W:D(2Y42O8J--+\6>6KZ@1g#FM4EJCAafTX,8Y81@F.;4+DKX-IZ+TY&P4NG
cN7VcZ,]UDG)/2I7FDf-OL@Ad]\fTSFOe>W]7_;g]S#0:[-Q&QbPV_J=(3O].3MJ
/TKdX@86M0=bUYb-)^D84=<8g;\:eH2Z.Z:a>g>09KW:@(,P;K^aV,Sg-;1S#Gcc
_ICdG4c7FJ:=3?ZHVcI@&IB6M(WTU^bRgYNWLaQ;gSB@Bd3QDPR#CQC8OFQ]1QfY
[M,cCW,d:O)HJ:.AWP;.a+<VWHMI#54[&/)Z.]RZgSdJ@@4dX#0UBU=c(>eXL=I-
Nb89/g+(;>TMHFeN_SQ=#e7Od+&H=gZF^:((=R^\=PDd\]V/=c]R2C,RNVZO#LZO
0e3(.XDIS3786?AX15)RWOUY[2-OC^eB.NX:caVCfEVbIb4G/L9>_.((@[ILSZ,R
ES(MB8Xc@=A8:FY4:c7CE>4<Nc8&XNPca02FJ8,U;OE3C05ER0<TVG:[eAcZYaC-
YI74Gb>?GUICeSM&K+I9:)JSUc+H51DM&g6))TQR]H>:53ZE7?e(/)eCD\(LK@6F
T=(g>M-&T063@Z2::J=BN;0-CXU>c-9([RUbG2K;c#a)K=T69a+eU@#c++QX;YV1
RW#UcBJM9@JcE=5H^cV>1&7HKEB)S/P-F6YRD.,[_I^2+Y3VN>G;??RP5POd9+PB
ANUgBeQ:0+>SVZXS72R4B1JYg?-+B]]^eCJ(QU>c\fCO1:M64CMd+7D4B\]#HJ9Y
.]5X(C31:-7A:&981(.\,bX7cE4FLY^7@V)1Eb5G0+>8H24<K,P&KL?fPG\.J6c;
3VMY9(#@T-U=IaW--(B>7P+0aI4R(Ne?JXNB\EVccYeeS__a7CUNW;;3RJ7fc.-\
GW94fD5OKCGY101T.L(RZf<SBC8+f5(Q/7E58#g3\U\K?.T9;gQSUXf0@97K+=gJ
VHKd)P8KLM+e@0-aB57cK=]=FBX&c4N\IJ.9bRXPFBeXf@5KU>b7_+V5&1fQ@:R(
>0e.0H-FEF5e?\H=RQcEX7K@&IAC,VaN27-0K;G7=+ME#-Ka<N3W3<N&0PJRa.&V
A6IA@9/G@/XU./bg8Z_675JOP=G,?0:XVebPBJWBeb2)X-G=N9JO7Z,^0E?.:^b7
@/E#?cR(Y:ML/d@e,7GLUY]G>@X4P@E]/9_N[13eT3S9=,O^_I1OK5+12b?071JR
:.>(8g2W)XCYWWNW,S<Mg[cRgVZ>]dU[\VKZ<:;1H#UG/3W[YY:X(^\>50TTZ.-[
BKX.OEc^,;IKH;Ig0AH_DcH9,Q:b[^a1K/J(Qd:5U:+dN#]]QE[V-P?gbC2PTe+B
-B7dA1Jb);[[^XV0cMW=D<;A0>9^K2&\gNAEfVAL4@bW[4]3H;LcCYMCAc7+>[OF
K[C(OgV)a<[0.,:4U;LXFNQ7Q5[Y.29[7,BMIAAZ70A0&V@7/8Q()6Mbb[1U?Ad2
OPZKgJ\\1U4WZe<d:?Lad:@[a-a]7@5EDbb<?4HM8@9KXQ;@ZT\^-Afc_KIHK[#U
(O2KP./(\)ZL4P;DN&<[/NX_HaA:TP,__&7?ZQG:+-IU,g)QDMC,F?fAB<+IO]&K
bTA?USS9I8)HQ:.5d5]2<eS6>58X,L7:^\bA]SJC&SQR[Q+?eU]0AGQ0__8ZIRI3
?Z2H?81AD2)Bg,e,1CDXD0aX#.)d<Ma6((?M^^9e#E3D43U29@1XIXMeM?=::J(/
2:,5BP^2bVZZG?LORO]\RSMgT0)[YeJW;K,6Z\KceYH@P)@.JF[P/TQD2fSXCddP
g)HW[da^?9Ue4Y=8I(Va:#aP\?@g1-@)KBC&P_,V=Me-UM,,)_.XD\Sf-+dIb7fS
2&8b;QV_KU-AU\#,<-S]4(PW#(Q]:gQddL9N]#7e<,FF3]HLT>)^e_+XD#=5f53a
13UOZ[Z,;g<A#DJL9&.?[eR,[b;;F,JN8c]\=]XF@G8M9T(J//VG3F8JO@)2YfZZ
>HI/3AJ#I(E]c9A79XH8&+cgSb,&fT-^BHHL8Ub/g^AUX#KL/KfA8\^:DUB;^fQC
I7C,)J<IAF:R(aa>(CK_Ad]O#SV,/WSa@2d/H/#Y,AVW7T-(R#:Lg],[Y3#O0F/5
cN\K^\04ML+A9R?KE7?fK]Gc]M0R?J0a@eC9<N.fHXaDQKG(]/84L;PNL^K8^E,A
J1A1-[ef9d2)?;E:KT3U;d4[=4O:EV2_/O\?T\H.\=(==-NCDg3S\V-)59]P2RFc
c1UMURCVHS2IOX2\2e,5BI=5EL^;3@B4-KQ(6SCE<C.G_^C0#-EP5:C,^I25LQ2&
((5^:N_VC9#;+8b/@,ALLJFVM,UFXQ,2E88cSEY575T=F@ZU]b9c/=5S\SLV<\2a
Da]<c0O@&-GFe][>>TPKJcMGW]_XK+#J2@<4GR.4/=Z](D7@HKWF]?3=4OX;L\7H
gJ?.#:CT56ZB(N@D&/HDB+8<cQ<E]]d)XTa)aF&e^\V,e=aUOeI+].P(FWfE:.7C
,eKcdc6R@3<^IMEMf9.gedA/[(aTENHZ(a\+?&dX[9>=>R51&ONG4[#PbTM<b.-E
dVZMMV_.g/fOA=<5EK&E+5e&U=KDD(M@Q>EYN)#f\c\\3K\6>aE^UL<Wa[Zc6^YI
R8\g#T-fNU)&.I;AVg142>c2AM2Hd\R8b]T^F7U/TXKMKdf@<;cM#aZJc/G;[:8R
3;_,QPF_V=60eM3-OPDX8dX@_[Dac1E<C./JOM8+dNU].d96)T,DA:6a5+:-15C&
QIbeS6735WIdQZaf(KS2G7SX1,1PDM&6RDaARI9UJF\]TAVVgcL7J#&W3FM:0O)Q
I,Y1XC]A^\[ge4?Ke@+H2:W](BBcTCNVPY4:WJeN)<D)LKFB:R]-S/9>B:WS)f&O
\,&Yf(aRKQ388J1M86BH=R^VM)aIPcbXI\/<ANK0.)CMU69)P_g49W6CYc?RcU^;
J=WTV]/28XD/\@Y<P<PJK02X-8<>EBZV@.;Z>S_5J>=1]<MVPI/&Wb_)TC.[O+M(
S)G01a[YXW64P^R0/MEVg?c9&>DGU9(55c>B.^7OFGJJ=:f+e>IE4G+\6@H0WW_K
,:ccF@>._^J[#U5G]gXS0E3Fg,\8#7:2+bY:5:-GQB(GY<Z49ZY:\7>GSf)X,FM1
H#VD#cMI_DZcL.QY1S+HOcg#1(MWVD9.b@L2<RE_Vf-cXK9Ta@/1ZO0KPP@TU,F2
]2QGK:<B@IY(f//K4E0327C8<:BV_UE=)1,4>Vg587]2eOE#P9AI(NF1deRYU4I)
1LGT/;d@77HWRbU8VZCC1\->fH[3QT1MG^K?M-?0Y<S<,WNF-bebKN1DXe[1:FTX
=_Y)Rf5e/+607\).[f<NQJK30=11#0EL]](\4TE(=;d;Z?.O44Z@.@M_2&N@X@P5
=+,]e3WPFg&K#.&+b0HK2::U,7#T?bG<8b8P&A4U&JX^(AAGRGAP2(1Cf8S2cQ8:
M95N8Y[gDG+OA0U-B0_ZYN6gD><OZR1)a_e>D#f2O5M)e-5]J.=M<E=SBc#V8I9;
Pd(c]KM[:47BTK\^SW8b;5O,(E5(CWHWDCY^+S,[YDe8a],K=,NYcCYg78;4L>?4
V\#HE9L_bd>][5(G3aKcgd>FR9:3+7g\N#H.PAF]9EZ[<,8#1VHfR5RI\?8VWB8H
O009Z>:7D2QR4?T[#=)_B\7P6>)\WU49XHbGO.7\eERS:R#IWD+2YH3=F;JFQ1bD
<F,.Q3AQO\)Kc@885G@-ERfIMVf[N<8-L>cY?SCJVJZe\E5.F5.\DS1Zc5cJ0FeM
(HYF_X-.E0Pea6O3VKNA1B(U4CZ2a7/,>?1#,,\]BQ@R2&[Yb6YE8M^BVU(ZFVX^
F;8#GW_0JI8\#XCB/W=TGG/,\\;.3=026N(M?C.[E-PW6I,->:88XAW9R>_e2Aa,
UFKB7DdYdZ[U]0HP>f+1L+a33?D_]RR<M^@@&4fN[P/)g3T872])5?D#4BGQN([F
\3e-^<BTV0agT9cEM3dHWRRQQ04IW@QKEUWI@)I.K=2/HgH6_O^OW9Jd38\4cg_Q
4d54,6A9\78W]gPJD4WZ,45FGW7RE692F3@>@GFb\5?0E,I2/UTS-QS@e,eS_,RD
O7]-Hg)2=Q&7B06/L^c+XK6Nc:1E(ON>05bM(;YG(;\2+C:8<>4)KRgd-P;FK5L^
#dVcf/5@L96\]3R7Y[@Bd_<cBf95ZJ9)/2AM.YZUMf+\H04XZ7>URa/(LHEU,Baa
O-5+)R/X2CLAc_>07<0SSC+[;MYI7d^Re)bd,C<O[5c-fcL(F>FJ^7_S_c[fZ4Ib
8P;L8dSJH>PWEHEEQ>R?T:KB?6a</SVHCT?0:A9Z69&]Lc;,@6I4/Q5S>Mb4O[[[
A(AIO6K0,:+dN:2RURc)344f_(+E8YcOLTPH/+8GJQ8C)[M_2ObIZH<1K8N3,^);
\_e\]@S41GS4I(SfE=Gb-4TLNO[--6)]28]O\g,aPZN9VX>L2Ed@dR)[WdV160C@
g.[<Ma\>3b&K8d<M2Ac9<ZZ>8@=1#Z_D.9HWC#=a@_d_7CS0TdI;[/]O_E;O8@?=
:HE3?A#2#8N<<[>)g(JE?@W@H@E7cD3g:S\EXABP_.Q_SX;GXX\B#74)35W<2dCg
+,;U>fNI8=EU4WXXbL1D3fJ;NgJKKNU\.VHNPDMH5MX.C/YB,>(FS&LNcG>116@J
8.WLNF/O^34ea,?#RC\?2WO7JPXRQ/Zg)8L2-3)XXaYPAeCX.][M\:)5:2ZZ[FVH
6#)&U]IfY(129WZHRJ;C-_;6EY,:D_gK4YP]]BRPVY[<[](SB;2SVU6c3AK_R@D9
+S_A6Y,J+X4>XJ\9-8>a_IX=G(bQJI:6ZIH(7B3O^fg5#[U,-Q6/@]:N52I<6;#f
TJ<Z=EB->BB=B@[_N.eSWRJ^DYYF@Q)X^&dYU]bZZ:/E,Q9B6OLYaPP0/_Ac.SP>
.AV,W(0d3YS5TUdEg#>>b,<C@-ZLT[EURV1_D;b@OAM+&<>82G;F\>_eTFL+eAJ,
L5Z_S]ZU?[5JF&M.Tc3CV]#efC/;\30:_U<=DCI1Y4#/J7bIK<;38CBEQ@C=9A.f
]4dc3,WRJ5R8S038#>_^R;,c/[?Q&(J7GfMP4;ed.P5+Q8.+AUR(>U^ZfS[EP2C^
OG=O;\f:23d;PW5H2Wd^H&R]5eQ&5?[Z\e98LI\,_-ZJ6UD&CJ6]Sg2PId+0<A[U
D<)HOEOR8G\)?+BKcVWgE?YW9&5?dPS^FWRgeID5J1L8<<+WX86[?4K1L7?(S>Rg
D00F;QV+SW-@gaGQVLaI[9(UN,a+U5c;/(aH9;Z]7]?EU,V3IH=?=O#(2YGSFWM9
GZ):0EE)G9W)671N7N+L>Xe#fV)H,a4KL+X)U;-=G/<DQ28&gd+TES8+VdQ,PH#J
/&F<[d)5K@A#_de0BAYRW1bE:+dL4^[IfW<>85?@T/F(8@Y06._G[NJKB.C2;7PO
VR[=,X_be2PKd+&+VD7-dECa#6MZ(KVFR\g_]@Jf^NH:OB@C6KCbN4Q<A9F[5,V<
8d9&6H\Y8KE;)+ZG[&GE53ZTf,dT(IZ&LOR?FZ?]#O:K_dT5H\X0T)C\ZX@G1He1
(U(IZW^:R8;OO;H@X(3@VNGfPDE5]0aW<<b:6U<IX@^?4^fd)cOZTXO9<5D+bD-G
UEK_:bU)Xd7g3&OaH?;GL_N-cea.<ZZ^UU]GNA#G0bI=#1S-P.cPK[0-N6cI_J/A
@AdLHf,)R=-KU]L.4O&a=A:,X[]TcGN93>9K&^W=K4+:EWBIe:O,,VaaAd^B])D]
50D?V2&DIbb((Q3b&H&Q+:VU1P(II)E_C:D^5;eZH)K8_)b5a<1J=7JWGDAb</@6
HA@6&X[40S>ICe<3N5#KX/cFQfa50&XBg6H:#1b5=e^X55>:.O+U8c0JCX^:R+d@
RB<-BF@d?#K,?7A^6]GF@(8OI;Wc2&I+-1=VP^c=SDF_RYTdL6?C>+CSIX5@\WI6
C[-[/528F\ZY\K#Zd0<()LX2\;WD2<R_)G\a>_QH8=?LJ2[35Z2c1#DdEP?U>-0N
=Cf<D\.[@H/gWBeJYF?M&AO6I3GV]5?[9MS<A(\:>9H2cY/L:6LU[Z?#.fg+A@5P
^X)g8^(b/86e9/P#4)M)<@CEIA790F?[;9[2/bO^,##Bg<GY)1ZH>([9?@;d=+>N
MOB7<AI//4#b#61Be9_BH2bI_PbFT9OE3Nf5]>bf1QG3(FI+O5HIC7H/?WbU4HNd
(>0M+:=GF_=-9A;VDeFTgNP#b);d-ZB;R5+eE[?e>bDK4_AUd=QD&.[?AcTId^.B
agH9(E(ATF<.\S/fb0XC6_TgG-PaU7bAWcDgW]QF<B.0B512C+Ea,4F/OIG&Q&Z>
<==BaL,:Mb+MN)JZHZ3N1B3HC0aI</D=edBZ]R:L4P.YXSH)7/5\AX^eB<3?df1@
&(+L5c?F49df;U?DJ:QIFX@gWF;HFgPEQ9Q?R,?F<FS_KL://F,(RQ&J4Y.(C3aN
fL5>GDHd.E+_O?6]A)U>1@JGL_/)GS-\H7gD4LG2=CN4&3O_P/87E>)IF:UN_9W-
J2@g2\GX^HM,Jba15-WDRW>BJ#MaU2QUOgZc-?46c7.G,a,Y=7KAJX<-@MH:e#/g
g7KAPDGeDC=]c2D-aHMYY?V@LD\D./+&LH2BK?BdIGO,T&b_WLC2]J40,0Le>L(T
b)+0A7gI1?AgC4d?>ORGQ^d^c&Y0<7F@6Z:BFZA^-:^ce9N]3QU-TYVaJXabR54e
bP0W@\YR>#b,(]];OTMA?0T_GJR@?RDAZ;)C[:>.J?)eEAfVRKGI>=#58=A@U5D1
;P>[-^T;&dG3<I&,L3Ic<AS-<e?9Q9C-NLF9DK>P:OM)B,L[Z0.c@BC-M(B=:\TD
<&89]S3-15LQ=#S[e0;bN47V=[30.2IJdZd/)ID]5:/L(US[C\KERI1;LHWJLR/I
Z3+:6URLf2c8X(5W&GSUOL,#U-2\]VXB@KFU3AR==;<]4E@AHYAKV010/]G-0DY9
(LP9F7HZa7/0)Fe.)_DDWMLfHNN6]0U80PI]GI+HTBK6A#K?Qf&Q1KH?;5>5dgT(
+)+g5Me5D[2Mfg_7?6ZX?C6URCP<)4>Gf[=ZIN4Tad_e(H]1-&[aS[=O-_ANcJ]5
I?-C@Q9VR\/Ag)8NF1KIE0KKWD/@PJ7M[)W75b6@7gV2>UH8Q3R(FN(=UfG=-QUC
H2/X1B/8FWD9QaIENM[>TQ\f&C5-)Q3H@\\V762^/-I;^4<JcDY;;QBSW9,#KS-;
DS0T+YH<)ZJN3>X3[+a(E8=J>5KL2B.0GPDN8VEcX,XXC+g[&;g8B/SJU0<8S-[W
bF&_W:^6;R4cKV(@6BE]4=G#eO/H\SY^e1X=&T7]2^5EDK^;\?\0UVJ6..(WHd9#
98aQS,c5GSPSLHaeF^6XVX-0^ITOGAa2UDQ@S3Ua([IX^-S?@LXFBN2=Zc+YL-f\
QA6eM;;;db@GYFN?+K<,Y\H70e1_N+-0TgUYNQV.^;48HKgM4d:WDE0TNR^F&Q/&
FVf:.M4Z7;/Ne)Va./P/5a9X[_?b1O5HHXbUL&]+(,QCMa9OX6bV6B=FUO_EV(b3
fD#DeZ<b-_Z.cA^8S-1I[\KF[6&dUEJ);GfNG6HVG#ebfY<^dE56MeL_9M0Q]ZTH
6fI9F\CCZIP.^+P&3]KKe??=.KfD+B\Y3JP-bLQWFX?N,#?XJeO=B54._ZNVTXLX
f(7SR+ZG,3M\8G(C-[#1a;FCYc^D+N.\PNT+?S?-9aVNBALS>,LV_1#5@T-K,R<(
9,b<_R.?V8bAa1AH)MJ3Z25)U0/I8R;56(LJ61X?P^Re40OBP<g.QV<,IK9GS704
3?RcJgAQdW?\GN)5dKMQE21I7]L5<K+K(4bBW;41=DXdL@<?EI<+)Ia+Yf(6K3gD
1M)?H9GH28MV.AZL4W7d=,#f+>fH1G3Sc0^49\RZ:BO(H#<K7F^V4=K(J5YNgH<N
8G+0F8;H=1N3#]S#Ye<Y4T#R[NWQ>7H<@6+9<d&Ua,)B-W^JBI<JeSG7-1FAB[KB
)H?6fe/NU23U#PNd.OBa[8,,=1ZgL_121^GFA?=Y8<MY^ZcF9MUc/\d+=D,?H)FN
SK6M[D66XbY1;Ba<9]J5M.\:f.AXO@Z@Q,F2dQ,:&.:77ZJeCS?:3+T,<25-<,=b
?MC=RWL+##D&\(a8f3^cZOF+M..]B?69#G.fF[3Y#g9:(C2^-.=K\\?&2C==+,B>
^Sb,UXDg6E:-+<BWbQBc1ML#?:fQ[VKIE5>OR[<Z=#f,1X-X#R4Kf-+:gU#_^+3e
f,A>VbV6.g^YEeGEM>P.f.HWAT@-K^F/,<7+]NBPeE//Ka@Z_?d\2?(K:7+0ECW2
;bNVgJE+\<LQ[:DNJRPOeJ#L1bd7D6?O1A+_O@QP;,9-fROZH?M#ZDPPbTSgD=UW
^VM#-1,7-SHd;_2@Z7.,^>07\BLVZ1MDA]XH)6?/9Q-&[/<_aGFRd0#X)\M\2.Fa
;-10A1CM@4S6RATJbbI(cJ^g.9YXG)>KPbR1cB(9\M.4L]2&-eAS0^-9H<_X/>L7
0[]d+DJMJPYF0fU^7e0<9,S_=_&-1.EL&(<^+VCVVK9SYEVdQA^=D@Z-J^,_T44D
_Q;&P;2\6d8N+M]<L@c<c.>I)\?\\9YZ7Ufc_TQ/(5(+EN>8RgS2&,?JF>XP?D&H
#6DSP-G&aE;RW28X+&U9DfV,5a,<+)3(TK@DB3\>YN;(1^C5V?YT=SD94[I?bY5c
cf>]?-H0/G#30;(WTN[6-LG@aTD89cC7.K989_-fRZe2QYVSD@KKO8d<eR#A3eAK
3J<?>N]3ENW<I,>]2NbCI6VPH5Cd6/02H:P]^._f;>^KIT8WY5I0^^VK8?EfV^cG
G],_<2eG]N[NH5PY8\2/HW=aQ&LS@@HX]ASbT<C]M;3-V]a\S^JJ]EZ\NMCWBLdV
gL0JE7F,;^e5bGU\DD;;cSc/___ZVagL,H,1TT#KBU#gCb26/4NUS&=[PGW)7VaO
TM7dTB2EZZK:Q[b5^W,EX3b2A>K&OT[-TC8GQHAU5YL>02B7[bM2feO2PM>DeDW4
b4K+Z\^1gHeJP(FDL8:1-NeNT(^0YE^Ebd.&@ec_<3/d-><>0eBM^]U6BK<2>Y92
S,SZC1a[S7]Z?N)J40QRd^HAeV8.ICX&]3<S]4(D3QOca-L:Z(d256O^,5eXeETZ
SQ5[DT19:PbNTRY_+Va?Q?+A05BJHQYMMOR8)=[;be\L6,>IDD74C6W]&F4C.O_H
PSXQ;HT@+40K?--]X(1.,d_^@.c?L2-]@GT.CEbCWcaZPY5c;(^GB\EDD_P;W9@d
)U?1@/101\-LcN33(0BM<eY7-a,9S.4<,aAdU7(BX-f4;8b99LNF40cG6-OON7/b
Q0_JZ(229c5)56c]MPV7)__;,(P;;GM6a<^gAbNDe>0#;+M6.#dD,DK;\MKR@BQS
^<V,R<+./.Fc.c9WPH)88-[P4=ea;3V=bSGP)ZFf05,NAAM-7.f/^ZC@NC7)CQ+3
cYc:+C[SdQ,\O/6XDBIK7T=R(#5,<LOH]S,/CQR\Z>.WE5@<.70W</fU;Z;G(@BK
_\@[-e#G0GLO2AH9:POGP4UAYa-O7X=fDKMYN3bg(W).?,<4<;Pg5./VF^3<cIcL
6d3D=>L59-c5E4SGTV?3<D^@Jd3:^)7/YZfHBWa\++^e#3f<@;@I)DWLJN?\aNY_
^/:5VM4LPA1cI;&?\Z:R8?PA.(f947/NKH5):a)49YfWXJL\4>L;KCB.#NT.,C>c
]b=0U)FH,g/^N8,5ge>>Tg6<gGH>>-N1<=<PK(cO)E,<@B/gL33R2U[<VKX5)Q_a
Q]6M^dD?KS5c7^8OVRZ-0PA49Lb)Mg&X_f5dDF9R51;\]4;S6N=].0B,6JgD[2T?
QW6CBY.ODGZ-R6&1b\bUJB;9[I(NFb=JTH+Bbg,-;D7G9R;?F[3Eb7DL(4U7\62>
Pe\WX_P#bO-DRAI-KG]0?\^YOUTL4:\b4U:9PTVfIg=e1IN8ZGEg#Q?A_X>9.WSO
?^Kf4Ub3PaW9@9Z_R20USaI_,Zc56#DUU)J@4MUH7<QfJ#7\\(I_:JUQUf)Ce(=A
dH_UCdaDZM[R#87?;7Gb_R.)/>#V)J7&A4fb-5HZ+HWI:Ra>/+_0Sb>IQ[PY-6+d
25TFW\[V7E8SI]^LE<NGc>TLJ^#6,.a2B5)Y);]I4=VcKV_]-cJSAU;DHSfTWQBM
eZQ0g2:a6I=N[KF+Q3>@OEQMabJ]16DA/d7;UZeG/_L,5bK,A&>4&9&->e-QEaBK
cJ:?d.P[J5dA.ff-JXX]A)a^?OWN=XR[)=^B?CM?=^GH:P;3<c3YAdIAQF6YL<2;
Td^WA&#[:<B=726[B7+EV(H:QW(48YMcK@NW>fSX+9\V28FRUg_.-Q.Y+K#cB-M?
T[c#O1(@aT^,/NUB4U+5_:M&J-fQ^[f;FKR<L5]X\IP7_P&I&EaSJ=Q^B>OGL1d>
H)5)BS7L^PR6^M:ZMRVeS;#b.H@>8F@BOM9#83fQX)0/MdNf&JPG;5#&12E<.[AQ
A:<:KLSG4JTbQfD88M+[SC97_<=JA#-N]/;<O37N1JI6]LDT@+?#7VJdC+16W]O-
:G?D3Qf?FN/=HR]1GF,Z-Td521UYBb+OKPD=IXJ\\e#aJN[a@]J.TRQ^;1:9F+(:
UBO1PHa@8M(+W1X[,B^?0(ZHO(D=SCTZ\f&7.f_O71,3/P,)S6aKf,R)+0V&/O9H
/Ka(V>/^Yd/^4bFWfRT(4@)QYG)aQHFfb5c_N_cbQZE\IedgDM_ANZOc4.F[Y@?\
54_YRBGGY#_/I>[;#QHaDYg))CW(H\XX#_@-4&,J3)?ce]Q7,?:ML\Se\@cA@TG1
2g0[MV?[D[d7fI=W\)POT]AfgJKf=Q1\_cRF)7N\c)JaA\E51AG2Q^RFS3[P2JX&
0Yc79?[6c?F2FTQ>Db;[O08aY^fJ]dCBBM1XPPH]W5a?&V>BP/),S378?.H>d?]D
SONb(J[ULF3db;A=>Z54;Y<35<b#\2+>PB1PUg/#:?Mc06AU5.T(V84-U[CX@PS+
4FUZ)R8H@):-0\6+6,fD_Af]7e=F@6N&ULAKC+.6]cBR>1bf:)HC(I6PRZ5KW#:2
cO(g+=@B;.3<-9](447c4+DZ8UC6;:XaEPW6T1=7B81OFAK\5ZI1<P0_P4,1/f=8
X+432/A/eA/-TaegeN+)7;SF24b4QT#36_aMFSH#^:5VX,(If>M_M?3^NU:RJR;?
cJUX:.#?X4W(_RJDD(U4Y#?dE6]8/>?9+U@=\VHIcd<YAD>A@Y([_PZU45]?W^,\
6_gS7OP3S?8S96WF84:?fWTTf@MX,;X(_UCAI[>JZXA1BAa^Q/](W^bc^DL\M?^?
H+E73FIU:[=QJ9ZHBd([N?>T/FRZF)WYg.c/-#)GK<1CO+X3:[;D=&#3JgJ@Xc[H
=B&gA=a];K@aR<I[@?&(<H=W-R586E8HRdg0UN5R9G@]Ad#IQCAJP6@NHb7,&K10
&4]MGH,.a=A]ZO3g:G^4;d5E\1V?W.=[^94O/c:,ONK__e@[(Hf6Z?F0=]4b>KJ:
R]W)F4@X-/AW7Z<FRR,&^G#,CfDV#I>(Y#(gJ-J.aT37OAVBNLG&^Eb5NGTC6@QC
;ec1:Q@>NU:Q=-#Eb[@-eFX<EgI&)/,-ad&eKDc=/MXY2g3+>51A]M(8APaAH)D8
_/ZD^JfOEbC>#5C17=WBPfG]YA1g>V6LX-Q#.<\@#2S-Zb3FFZ4@:bMP:G2&?K//
M8C<B+H0Y0^:\.d2S8Va:I?>eFU.ZB+LM2VS(BYE;N>+QgbF)L(VeX-/5+c_MOR/
>-f-07;WFaD;)FG[;:eZc6]?FWB/9D]PeXF3/Je<R@gF49=P0[EJ#Vd6&VOWGC#a
V0PFO=YFGH4>3NX4,7^R5&,g7CEZE?V8<Rb7+gOMRFP@>@2bBFM.>2A9a<gJeIRQ
H;/b9I.4EG4_(Q5GXEf#GW>Q8JL,CRP0W6G:5BG(+E7<DUeY2VO^QUW3#b7UOEbg
1Wf<3J;?[Ag2)5[IMA\>::4/K/=SZ[B1HUX/e:<OG(NdKWP(U37H9/L(#R4Y&CXX
&@dTP/X-J,(e4(>64d[0&2^QJ+5R,KCSUNc8H3bJ7O2VL4HK2MT<K52L[+;51KMQ
dcXGP-BX:;?+Xe.[c_>8a;cZfU9W_:N55[Z=F?:NP1-9O3.d9(1_8a(,b=15_gcO
@L;>QX.gff<P91YO,\EV,2LD9cB;=dbO43-&HY?g0S3L+eROW,+0ZJ/[Y)7f.ea_
N.6<?_ZK]#-QC&H<bGD3B?]1YJA)<?H9T6WCg5CdE(JS&D<A5-gN_4V1N.5/4LV1
]7BB;)g;QSB+()J<Y.BJR:e.5U[YX)JZ:d[+\\A8b6N/.PON3B4MQ#ITFKfQd0^B
FCHI.8WMAAYHPV3(52/@fX:8];T4g9NKS]@#\9Ie6(K_/<2fA7dBREX>&3=[Wc7)
6=FNOP=Z.<3geY4#^g7XT]R&e_145,2P\:E8Ag95BYIC/aU8H-O\7g86(fW+JacF
_Q4ffP:\QS:^ZS&KIY:;DA(:8KJS@XeTC[d8VU@OCZ8DT@U#(#Cb\e<3NCH])#[-
,^d_/.<M,[g23&Ig7^Y+(+^P\SfAf-0>c_>:#<UAT\-URd;/;8VS^YHN2SX\/Gc9
;@bD7(Y^-+G4MIA:=T]K,J6+U_.JEBTB7;)7E<cS3[JS^A^@0ERX+;<93Eg#CdWW
L.6IMD&>R)822B,#Reb<5K-]26[<6eWDF<A;N^A44,#VATTK.N]eg/=1Dd_;3K2f
3dTSXRRg#R/LN90RR19^&2eK.cS)@+I+Y>FYFd]Pb/H3dQT6?RT.+d59,/\C9I8\
c79.]bHf^fIA6OGYGAcALMa2=+9N>#3#]W8<)IgOE=[bA^UAAR1;^(X)(58Z5[R?
01[fXG;BSG#W6;Wa/55U4<JIV#0^.5f[d8>96GdM=\>-A@JE1@B:J<L3_;HMb:a3
Z>&<)KSDD+LL/ADE>VGO;K;\[9/W(<H^B0].JdJ4)DY\bLC)]<-1.XC+fKd8Pa^1
NSb?3O6UIH(@9QOXXb[4FIKIg>35b9g@4O-FdP&[X14@3]eW#^2U^P=,R;#=O.8>
H#.K=?_b;1/eON6bD.e?(>U2>\Lb>aZ7?17]L0^P;a])X;:3A=Q62DQ#._(.3\-g
5VT89c&VJIKG\09?R]KQC,RaK7(].)9\-UJ[J>#]..;\PDF:B=K?BIBO+#8gG>LV
)RU#A19E;a1gb05K3QG43+H&/YT./DEaWaB8#c^?E&CWW748D2-IV@Fa6E(C&O+\
C-5.eT8:B<)0@&&fNdA&U&Jg+15PbG36G/R#deHP?K>b:Fg3[AJ0/I;0FU/;3=UZ
)==aReY<S3g>&Qf^aA5+KM_75TP,AG?8KIHC>Fa2E5=R84=a=7/+-S7\e>I.])2e
;E[:LD.gB4-eeQ>_U^a)CS5Vc#Td8J0)I5?8ScI9A[U?ZC9>/HI:+J49AP([74/V
DPb<QOHON]=e_aKUaY7<0.NNOKaKaKDZK?J5e?WSC(Z.bNdNJUB>.3)6:;2?TZ8a
-WbLAME>#LT=cc>W6e5#RWG[PVJEU@-B^f>K>_IcDN#ABD-VO(_48]SKeU@M,e:]
SP([&W-OY(7F?SMT.=\d1C91WXH+49+HJ(N/2B9:e[\Vf];&K)^@a]_C76#9_D8A
[9g?adKRdB_(B\(g;]Fd.6T76#+784^:0TEC<NGD=_=JVe+5:Y-U?N;_1Y(RK392
eZQE\]D_IMN4f&Pd1a]Cf]_Z&2aQ>/YbaJ-J,R8&\M7/Ica+_f:0/-PJ,^=(^Y2Y
V2ePQMaP],_A7@ATPF,QH8LfTS38B)1N7O=G<<\L6L^c:]D]9(BBfP?N392:KUVN
&RNa1HV08D]1AW9g(KY_M1SSY,K2_#U8RfPUXL[1DN##d[@P)bDRW)/8G@bZTMFZ
TZ;dCRNI2Hc<,PILQ@).]=3A&W](P7Of+):=OEB10O,WgQ&gQWBFbYEQ=+If_7MU
R+(HRO#MJW8Q_(\B)3NK:Vf1NO6H73[+@e4B;@#ZbZJF(R(R]U[dEAAE9d5KOODT
1IH:BN.;L,N6/f(.J^C<DW]aa[Z22IEa#g4B=2MSaWN35\JfM17,MUdb+@C5:33f
QCDdIZKNWI00c;V8OJ^C=(0,Q[(H6CFT1#_IHWNc9(+-Ea@:Q_[I;26.@d6Rg<H)
]BSL7#aS.H,g)da8]SKc(UHc+c68eA(C/I9MEf2/=>7F+Oag,A#82c9,5NSZPIe4
UE8L8-U9.ND]VA/B#79??6M3H3d@N],2&dL8@I4<Vg6>ZGS3[;c5;HME^G9>4dMg
aM83VG..[88)/AOPcfP[a^D>>&8+QL\TZRP;VBFRAO9#HS(,GX)VaLZILF^VL&HH
=5T8P)2f9MH1LLQZOSOYc80&/#.#H_0OC@9@WD3-@DLV5.W(eZJWH.W#J++<B&)X
g;gg7S^^[3?]+\dgP1UbMa-Z^FQZ^Hc;R:VNDd4U+KXbX7\a428d@5d#()&V403X
XBW=8U&3fF2;7<7PG0V4[HR6/JY2-P4;Z##(_GR]JOc#fEV[S:RM^709XE:\[K:L
ODa3?d=N<N[8)()@:FSIdbHEVL)U,,->Kd<P4dKYeZaU30cR4PL=O3E;:8g@?ZgB
3b^9abMG6QP;)K+KM-c_W_A9LA06S=>?OeceC&DRPb;cC>(&.Y=e&Y^K]EGEZ_RP
0FPcZLgf_1d?XS+#CKYF9b+<ZMH1b&X>)fV3B;;/[6^W4UaZ.-dG<)c:;D,E_D0d
AMR5d.SAN?\b3Ka7VJ-Bc4-+S+Fd[2\]&-_S=+aeN,>QHV^+,=<R,8U^BdB1fZ^@
4<Za\D7((CO(d06,E[H^FHA:@,437cU)M0X5)RPTB(_V34,0IMFL@0\-CdLMS@VE
ZG1eOeJU<0A_M>(##\/+A8?,57/+dP0NA8:\3E?g(Sc;<U^5aIE(26Xe2@,TJL>f
8_9K\gD;AB3/Qg@g9-O460Y.D_)HO)OQ3DXLe^g+.gM5[\fJ01VUY3?#(V;V9\e,
S[J26:L:GX7e)T\8I[T?K@,fX;#[KLQHB\C6>JdA.g8HM0</TK]RJ)(L<9AGO>W,
HL8+Hg@Q6YMIL>P_EgP+\S/U,UAc+N@KY?N)L\):VXb#?7VCU#b>eKWJZ5&8E5SN
S8?9^Y\b>8NYgb8f-_UOb4eDE>f[KXUX\Q^&g&=M-/H/XFJ(:[(g4DTZDC9P@5;c
)LX4W@5G<]6SO:@Q?f9OgDR[:RM.1[We:OZg>0(DULb)+ZCceOIDU_De@],,4CX9
5EfEdgQ<DW4;/U5C3P1&W4P4GEWRYd>3Ge;K\,3f/FfASfb3QN1T9(23;YPY64Q:
68C>g\c:<eF&OA-X9,PecQDMO@AMA1AU\d[VIa57PYGWb&3Re736BM2A;&Og2K33
c@aNVfgO>-FSf-V5F\GF+c<N?#9RV0TD0XY0?K3NeY=c-#\@PU<0QLCG/X8YNcL@
QeT45GMEPNAg39=6CNc0Y.PNA]dC?-NZS(T_KNGS[LHI^N8;6OCN^1)]L&08EC),
X#>NN332D&>>I5#]C<+Y=NT>3-VEY)Sg+=(WF^WV@[E>]Q^]6d\WfT<bfLWbg&aM
42#>GcT05cgN^\>0;#Ba:Ud+1;3G#KS8B,H9L+B9b)<L<X9D,<4#40P15CLO^KKb
32-ZEVG#.+d=OR^T^gDPZ_LD^XO0&/7WgfH(gcJ^O@L>JYVF4+0]3JQa[#df7b=T
];J<#f_=3C.G]W3A/;\g&f;3\\/c^Z)S9/E9=MO-YL/B))L7((@)d,7K?e.c&JAD
J_;^bHLf_Y[/)IKb^eZG.bHZ\[+;W>BU7Y4HGY=g^+8dbQJ0dS/3#;fA(_3.ZD3#
VdUH?)2R<],C[/7cdFW:PN(7d3fWW(fLBS<]Sb>=>&@J@KN0FR<_GGMaR]#,Yd8e
[<[_UQE;(+:D?.M/(=1.;W<@1GR._]AR#E#G,0O7>YO1W]W39@T.+.B0VYd7LaHV
##KYFP[2&I;A#VOb52J7>gd/gYHg2fB^9O./(9.NUI5OAb/D@e?^TW=7G/A,e0OJ
07;S.(e3_<R;OJ,H]+LY;eGPPVQ=,Ja?L[NK[KUE:]>=T<O4YbOB>Q\?dQd9:G>K
PcIN@NZQL6HIUBJ7TL18XDGCNN;1bEPP7/&T3G5beO9GS7F[7LUAbXV;_/aH3&GY
C[A0e>.eH0&&R&(@-N(ZC_Za/2Z]#a9(ZS(U[T:G/WAN0T/APeOdcAbMKG@\D21d
Z<KU1Bcc?;ae:P?:eP#/TbEf)#T/@UJYE97O4aOYY>[F>01]JMab&-4P[5PfUb(@
g/f4gS^M^KF\Ff<3SLT?E39#8X-Q^[FM(deC18cK]b,Mgd#(3gB=8_TFX]F3C#,)
,8La0648H)#4JDYEd??eWMW;OSa:2O)LAN\9IfSG6LY>V?Pf&LU^WgC._N\[P^X-
G9LEELRKHG)V,3bB39\0U#a:d.:a?JNY-<06P_M^8<@]O2eWF;42\[L(@5W5&DLX
663@#\1S;Idc^C\QOF\BB9F07bMDY2L3B&3__YHLYP9BHT?/GgW]1_YV-eQO?:.^
7aX_3D?d&E9SQRA9EId)Xd-B<N.Zc&;;PLJTS@Hg989R2@0//:W@@+((]=BJ?=eV
\B76QMGAaGPf)_#N)N8TRbR^VZee=GS:cBddH@.[=T#P/;H]MN6g1&5&QFW.=gc@
6CA,;NNdFS]\0=UX-/g_HC])UPQF(a^_20U#fV4a4CG1,4+=d--GJf.M:#4cA-,;
@<aB)F&0E#F)@aTNMGCNQTRLgR4b=a<BbIRQZ3)ZFWRD(@]@G3S6=;+L&&8H-(0@
;YXaY7/LJD=N,L=BUKd_989P=R5<]c9a5f7.E/gKB4PB1dAKc//A1+Qgc6a28UKG
fS_S-2)E,I[Q0=AXFEB?116bebGXF5dE9)G&f1<0X_3a@VJNZJE0Q=/cJYcOWX+L
,35P:>.D7A.<4/QcQbB/Y[,1K(+6(G/DeMA.CT?-OEN^@9fS@KHg_4c>/Y(f_/XV
GDP^MF+MPS(?US(5XTMZ9,)21QC/&5]G5G2CQ8Y(Y>-(P@D9@D2OZ]Mbc/b^WJ;B
3Ce6Ng09VC(IH6L&=>(U?KXJQ3bc[W-ICa#0SF?0P;Xc6<]6_bHH^g2-7c@;DZ1<
d,RD_?aCA;OfPKY\O+/Y9]X\[5fTA0BUe:Df6+c)BGW_BJ8A)LKTSCQS?@LLHP@L
gT^QRfBGeS;4g9Sb?C1?/EDEg(-/&c59)4?:D>7XX1XO8PKTP#;5=),ZgM-,2fY[
O96EZD)c:NG=#=-L],EUM:dGL&==+c:&L9&g8Q[L-NcVT[(LP-4\(BG&YVC.E_@,
Q-:cbVX5VgUBAa9EG#@a0CZ4,XKD;SET5:288\]S]3R]:[ZdKc&TEZCY<Pf(fOB8
A^#.GWV3RDJ9;>R,U4FdLbHBJ=GD=UR;P5ZE\^_-V#IAJBGYF(KJVKK5X&GM@I:4
aBPF@3V<XLC@5#L;PZSNHagVgc6<d9XACC:L<]MO:Z/ca,P>KR&ZT_1OK>_XNLK;
::F>ZI+4J)cfOCBK;FFTG\[6b^56T]VMK.cC2O9^8D(\>17[^RY#33]ET<Wg@eXD
caZ/,C]1^.Me/ZY4^[BP7AUG)OM39#PT#8)/-H[#@ULBCgY>Q>C]T2;75K(E^]2f
[be)8#C/40RKOPCP)@c^6&8IM0ZBGd&<-5>5UWI5\[1XGOEYBBO3@A7fX9Wa\N4A
R;]bGHVN^R?^&g2?CDFP]F].E,ZR7\N7@KL9SFe_Wg]ZBT\&KDaK40\/5g8&&H/6
e1aS<gX,dS5F05WETc6B\6-7.PH/g:AP^\FfB4(I27,KYK1RGe>4=K(a=):\:a9a
MY@8<HVdKR^]aS69<SC5>:+d=3B30]ea37H).W,,9KLBc5b&<4M8DRUTH(@:&>g^
GV(9HB=P3[-_Wf=g3Z2c.J/ITCNI9[S;L;#G,@R^X_g+7cdIORUM6UAS^,S82=Vg
J028fM9H<QS+ED=JK)+B>/_F=.=Td0=94JTUZfW9+fa>f,5NBA(2>@=[3M0.9OG)
_2X3#O@J@#K4=J32_2((\fPOg20_E^STdFM\FF)Y4OEGJQF6?\JW;SfT2R/,RJ.@
?aSdVX=/V4#+:4dS2X.7>2;IQ)I_>TKV(Z(aLb>cAgGO@eY58:7K4JS,>,TUJ_T;
.Ke^_4Y+&LGL5EEM;IA)UO/F)H?794E^Gf5OQN_egTe#M0#\CNQ5,8T+MT8]aP7f
A#ZP6QJG)&CR3e12dVcM5I3,R7G:a/T(ERYHZ2.-B_L@WR1bYEg9d,05e?J,+X6e
ecK]bCW(73^(UK9NQCMFG-(/I1L7XdK4H4EUMGe;&Pfg;>U[.7R<7c0#)HL\bB[1
;NZbaN)Nc+gW:0,CRI#8<HT5H6J[<a#<2bG]@2-R[f\N3?g[C:gSC..:U\/0XVb=
QEU.6<]_V(WZaAW3N+77-_Q+c)B4Ra&?[XfZ/BWFP85N-TR3XRNc:Bce(GYMDAfa
V[<]PXA(FMTP0@BaLUK??KUY#Z(R6.034^OaP=8,O^d+F#&U,I[S#BJB,X&O=U]_
JAaHE;O?_,VT-NE,\0^[JYJ/BJN<>_dR3-0T\g=\7^/2XYR&d7FPX<_]FQ/CH<F\
(.Y61d0/X>0DfRL.97>U,aE[5H2GBgdJ?NC^]Y0&f,cU\SZA#;a=:eCEC?.0(IC,
H5AN2A9(LZ14\P&WF6(Na4I^3@a);Z?A:(Vee#6+YZ-)X/>a<LGag[UHI9K1c3#M
#dY6]faY?8>/+W]1\R2_1NBD)]#^&Z5;e>(XN?.dII7^Bf#4@EOfWDCa?8\f[8SF
NIT[M-=1TW\=VLF:]e897N>VQOcN]U+g1DcT02/;<e,R?9QZ>4>RRFQRUV,\HP([
fa5_N,KWM6(PTI[5A>:&&09P1E/#N.@VCD1g4#a?<5JW9G\V6U+[Mf<M0:K_)G^b
4:,B[:f.)652E;94adA>7S[?]-Y[<G8;^g2+NgRPdbC/JYYJQG#8df+8L,,_10S0
B,@]/J2E;(dM4cP>f6U+f)6GU[>g4&gNBQARY5dQVHEcbd&[J<,I:JOB0#F-cJU;
QVaJ4XGe6(:[V@EGSH5DKf>5@[YI;Wb@G9Q8UA?D0OCX.KY(]]XbOW+?cH8:,,?M
CIe^C7T8JS,f^J/^Ig?:M5RG6G[?H4<Y.JQU,\3FN-(F8GZ@PaD6BAF7/&RLT)c^
A;0gN+C@MD\<1&W^LKX]=aC)7O)(&^d\^-Q#<3YdACYdB)0#F-/OAM\IV4PC[XJK
&WES@]U>)M@GHdHeY_E4SLdR.EO^EQ#AJ0A)Q44>P58fAG,1ab=c_=YK(V+g\KA2
PQL;L)S#E8^.M@M#aF@F3_d)J^,2fOfOfaMR0S\aC(/aM23)H?4#e2AHV7Za9[=C
ABT>64ZX:AWd_8WK^g,8ND;+aG?@]8.V2L8/2&SE8bS-C:T:3T6MYaJB-R],<_<F
A1LcY)eAe].;L+0Y2/Qb>3-+COUZ(5T:Rb4UaMbYT_IM8c.4:]c:<d6K2XcM;QNX
##YN2BBHgeeS=9)Hg:3\S2;(C>G&Ib:#\1H-bf/gFgd_(A>D(EROGRI.KX6=d(8Y
))gWWR/.G9#FBC8[Y8T?f(Hg)=OUe9V0Zd-P.@1?Qb0OIO4>eR7R=.>G1VDY;4H>
KV[@\?WX,?/e#]e;bd;LKC:2<CEd)3[[2F7IY1Y@5U71^YL\JFWYPdRN5c)eQY)&
,;ZcQP7M5<CBE7dT)-1M-L=?FbA.(6ba1Q05YMY4>BI=#dNK^^E:5EK#.Z4&d;=@
Fa-_HPdLWF_c0I]MV@eTf[)b,Vg63@6-0@.PG#e@0(VZXU.0,_fb<&1gI>]?P1LZ
E0L/VHWBW84?O0<FPV&B[bfI6E[]Ha:C98C]&]#<HK\,&H,HE0R16=Ob0gS2SKgI
(@FLI9=2cE5\U]5c.:f_40MREP;TPKUH(8FOe@LeE3(G6/8S,F[F.gYQLUHBJZ>]
@=ge@^4e<4KJ40U0)V]MI_U&&.R0Q=DAK^JUPc0XeI686Z:?F<-ARVKH9fBd?c)V
;6&_[X##_BEVbe:)fe5BRcXP<)VQ-D@b1W2X1c#Y?S?e:M1UC2TD=VL)XO2EECJ0
(BX1OLEHL9cORH6-<B.<gUT3fF\6(JN5)>_(T8?EM[Y<6#8fITAB<KF\;H0/J#,S
]0&Q;MHb<=bE2VM,fP8/e2+6A_?0?&+g)P1OfZ+B[eHN&dIMX^dfM^=;g>[bSTRN
TVPQ(/ECcgF4DI5P25QUV8.OSO<F-c<(/f.Xb7CT;3]T>fA<5<YGdO?G[6:AUf&&
4VAE4c7A2X@N-<b9_[)=.PJS9U1c)BXQ(0&9PKY;I8Q#c^4EG[\I:Y=R9/[X_dWP
O/XH;<4?5(bb5dS-W05b>NYP:d,B_VdQ5QQW8((LaSEKW.Y[IBY>0#Z&YF:)R/X#
>X(_&-]0)3OGP^f/XU@&KS3c]]H:9B28[f(4GdP66ebXf+N]LMeN+\@^O_b&S90Q
YEa2F3_J6I5&gP2=-)MDC10_?5,W>;TTH>-9d&IS?]CJH1:J?gCJ+aVKZ#Vc..6F
IVdPBRU2;UaQH&H5X>2VH9BHP?CC>+UWAGX2C5J,VGO693:##U88?8>d1:PXf-Xg
bga,MXYM::8_=P<UAQNZQ=YO=-E7-92A^XUSL<06,PRB@K+=^&BdM@/V8HH>-M#@
4-b>AdKbSC6B\++Td9IA99NR,S)5V^XK5fX,13STVA?<F4Q/\6Y0@[0SGK\SQPPA
03Z1]c2)dGE(_FQfDFYQ#aQ>JVOKS)MQMNQ7Mg]N<Cg]6LKV8ETG+S4d#\KM)6\f
#C=A0_?Yc/F80)]4^FKXH5+??7CELO<F?5eBO?D#Rc/?VU<NdE[0=PXP&W-6cM;3
&2Zd7S3F8H,-C1YY=Q:#4b+0BJgSa=D<]T6876OQ,BaF3<D08L.G7AENC9_G/,J;
g5LWM.CPA1)DL@Y_.PDFSI6T3Yc5J-RS3YE.)HSK&5edQOfH2#P_[644)S)LW\f:
b/Ka9<3)gM>-Ue2\HQ5VT@]&6NQ@8P+Z;#&WCP3<,g-U>/D7-V?9TCdXX5gD.[S;
(XFFb_FX<K[WdR4N?\X_U+#>+3V(PeKD+aZf^&Zd]CK9;?JcCgaAVVb90^G8RRZB
IF):NXGSQI.+7Z+E>1Y7&3X8ZB?\93H9-Ve&B4)Pgg_)]+^;eZ]1fHV1E;bd&W+&
84a_-\K_-J48@Ze/K@.\_6Pa5YM1?SI4c0D:]MD6=QVCE994JPa8Sg]Y4I(1+d[D
B>#;E,4f98EY3U>RU#+TGeG5>^cI)[e[@O8(93XRGJ6+YJXFFO1Z;SHV&Y-6QFYW
>IJ=d)(L?Y7.gQJV-):cF)JUC@OWB,12:G+Lc,Q9U_?3?MUBc/g7Z/DSb>C&:MSC
<->IAVS&;dRH-/R/?GF6(&JEXg03<H#]1N7&(.I>QS[@X5F3-F8=TKX:ZbKJOMOX
J&]3eY\TC@RK4a.9Q9<FHb06JF?6#CYFg>8:V_#BB-d)>JF1BY8D&]=ZO)G^,2;,
PMMcO^A.eLUReY460?@[>SG&887W_V>)E^??4.3NGL&65eWF(C?3E0>C-)BcEa9(
,QPXILAX/0>-LbQ0(KOYVV;92Qg#d)fGR0T48F4PfKX?1_^4>-,L/F[D/d?g42gH
ZdFCYLe=3V<>I9A\ca5E<VE5V^O]F27C8QTBf:GTJW/N(O7KN9<W#WPLF<#MM^&N
V^M(5=I<Nb/&?a,R8-eAOUQ53Te5./JeDg9H:I)-,FN(a()d;(D/cbC].=PC222@
cL23SH^VWINIMHO(CP?GL38_\4=dT<b#gD\M=#@+QW)J@bQKIG8;4G:7gI,:;NVX
H0LB^2WeG.YI-$
`endprotected


`endif

