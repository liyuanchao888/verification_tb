
`ifndef GUARD_SVT_AXI_SLAVE_AGENT_SV
`define GUARD_SVT_AXI_SLAVE_AGENT_SV

typedef class svt_axi_port_monitor;
typedef class svt_axi_port_monitor_common;

// =============================================================================
/**
  * The slave agent encapsulates slave sequencer, slave driver, and port
  * monitor. The slave agent can be configured to operate in active mode and
  * passive mode. The user can provide AXI response sequences to the slave
  * sequencer.  The slave agent is configured using port configuration, which
  * is available in the system configuration. The port configuration should be
  * provided to the slave agent in the build phase of the test.  In the slave
  * agent, the port monitor samples the AXI port signals. When a new
  * transaction is detected, port monitor provides a response request sequence
  * to the slave sequencer. The slave response sequence within the sequencer
  * programs the appropriate slave response. The updated response sequence is
  * then provided by the slave sequencer to the slave driver. The slave driver
  * in turn drives the response on the AXI bus.<br> 
  *
  * Note that the slave driver expects the slave response sequence to:<br> (1)
  * Return same handle of the slave response object as provided to the sequencer
  * by the port monitor<br> (2) Return the slave response object in zero time,
  * that is, without any delay after sequencer receives object from port
  * monitor<br> If any of the above conditions is violated, the slave agent
  * issues a FATAL message.<br>
  
  The slave driver and port monitor components within the slave agent call the
  callback methods at various phases of execution of the AXI transaction.
  After the AXI transaction on the bus is complete, the completed sequence
  item is provided to the analysis port of port monitor, which can be used by
  the testbench.
  */
class svt_axi_slave_agent extends svt_agent;

  // ***************************************************************************
  // Type Definitions
  // ***************************************************************************
  typedef virtual `SVT_AXI_SLAVE_IF svt_axi_slave_vif;
  typedef bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] max_addr_width_data_type;

`ifdef SVT_AMBA_ENABLE_C_BASED_MEM
  //Memory core 
  local svt_mem_core mem_core; 
  
  //Default Memory backdoor  
  svt_mem_backdoor backdoor; 
  
  // Memory configuration 
  local svt_mem_configuration mem_cfg; 
`endif  

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** AXI Slave virtual interface */
  svt_axi_slave_vif vif;

  /** AXI Slave Driver */
  svt_axi_slave driver;

  /** AXI Monitor */
  svt_axi_port_monitor monitor;
  
  /** AXI monitor performance status */
  svt_axi_port_perf_status perf_status; 

  /** AXI Slave Sequencer */
  svt_axi_slave_sequencer sequencer;

  /** Pointer to common class */ 
  svt_axi_slave_common common; 

  /** A reference to the slave memory set if the svt_axi_slave_memory_sequence sequence is used */ 
  svt_mem axi_slave_mem;

  /** Reference to FIFOs in the slave. These are configured based on
    * num_fifo_mem and fifo_mem_addresses of the port configuration 
    */
  svt_axi_fifo_mem fifo_mem[];

`ifdef SVT_UVM_TECHNOLOGY
  /** AMBA-PV blocking AXI response transaction socket interface */
  uvm_tlm_b_initiator_socket#(uvm_tlm_generic_payload) resp_socket;
`endif

  /** AXI External Slave Index */ 
  int axi_external_port_id = -1;

  /** AXI External Slave Agent Configuration */ 
  svt_axi_port_configuration axi_external_port_cfg; 

/** @cond PRIVATE */
  /** AXI slave coverage callback handle*/
  svt_axi_port_monitor_def_cov_callback slave_trans_cov_cb;

  /** AXI Signal coverage callbacks */
  svt_axi_port_monitor_def_toggle_cov_callback#(virtual `SVT_AXI_SLAVE_IF.svt_axi_monitor_modport) slave_toggle_cov_cb;
  svt_axi_port_monitor_def_state_cov_callback#(virtual `SVT_AXI_SLAVE_IF.svt_axi_monitor_modport)  slave_state_cov_cb;

  /** AXI XML Writer for the Protocol Analyzer */
  svt_axi_port_monitor_pa_writer_callbacks slave_xml_writer_cb;
 
  /** Writer used in callbacks to generate XML/FSDB for pa  */
   protected svt_xml_writer xml_writer = null ;

  /** AXI Port Monitor Callback Instance for System Checker */
  svt_axi_port_monitor_system_checker_callback system_checker_cb;

  /** AXI Port Monitor Callback Instance for AXI slave ports of CHI System Monitor*/
  svt_axi_port_monitor_system_checker_callback axi_slave_in_chi_sys_mon_cb;
  
  /** Callback which implements transaction reporting and tracing */
  svt_axi_port_monitor_transaction_report_callback xact_report_cb;

  /** Reference to the system wide sequence item report. */
  svt_sequence_item_report sys_seq_item_report;


  /** AXI Slave Snoop Sequencer */
  svt_axi_slave_snoop_sequencer snoop_sequencer;

  /** AXI Slave Monitor */
  svt_axi_slave_monitor slave_monitor;
  
  typedef bit [(`SVT_AXI_MAX_ADDR_WIDTH-1):0] _addr;

  
  /** Associative array which used to store the write data check parity values. */
  bit [(`SVT_AXI_MAX_DATA_WIDTH/8) - 1 : 0] datachk_partiy_assoc_array[max_addr_width_data_type];
 
  /** Assoc array to hold the value of poison in case of ACE */
    bit[(`SVT_AXI_MAX_DATA_WIDTH/64-1):0] addr_holds_corrupt_data_with_poison_assoc_arr[_addr] ;

`ifdef SVT_ACE5_ENABLE
  /** Assoc array to hold the value of tags in case of ACE5 */
 bit [(`SVT_AXI_MAX_TAG_WIDTH-1):0] tag_word[bit [(`SVT_AXI_MAX_TAGGED_ADDR_WIDTH-1):0]];

 /** Gets the tag value from memory */
  extern virtual function  bit read_tag(bit [(`SVT_AXI_MAX_TAGGED_ADDR_WIDTH-1):0] tagged_aligned_addr,output logic [(`SVT_AXI_MAX_TAG_WIDTH-1):0] tag_word_);

`endif
  
  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

  /** Configuration object copy to be used in set/get operations. */
  protected svt_axi_port_configuration cfg_snapshot;

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
  /** Configuration object for this transactor. */
  local svt_axi_port_configuration cfg; 
  
  /** Common features of AXI Slave monitor Component */
  local svt_axi_slave_monitor_common monitor_common;

  /** slave agent instance name. */
  local string slave_agent_inst_name = "";

  /** Address mapper for this slave component */
  local svt_axi_mem_address_mapper mem_addr_mapper;

/** @endcond */

  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************

  `svt_xvm_component_utils(svt_axi_slave_agent)

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * CONSTRUCTOR: Create a new agent instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function new (string name, uvm_component parent);
`elsif SVT_OVM_TECHNOLOGY
  extern function new (string name, ovm_component parent);
`endif

  // ---------------------------------------------------------------------------
  /**
   * Run phase used here to set is_active parameter (ACTIVE or PASSIVE) for slave_if  
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Always constructs the #monitor component. Constructs the #driver and #sequencer
   * components if configured as a UVM_ACTIVE component.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void build();
`endif

  // ---------------------------------------------------------------------------
  /**
   * end_of_elaboration Phase
   * A local factory is used for all construction within the VIP.
   */
`ifdef SVT_UVM_TECHNOLOGY
 extern function void end_of_elaboration_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
 extern function void end_of_elaboration();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Connect Phase
   * Connects the #driver and #sequencer TLM ports if configured as a UVM_ACTIVE
   * component.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void connect_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void connect();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Extract Phase
   * Close out the XML file if it is enabled
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void extract_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void extract();
`endif

  /** Writes a single byte into the memory through backdoor at the given address 
    * Note: if any of the tagged_address_space_attributes_enable bits are set then
    *       this task should be called with tagged address. Ex: write_byte(xact.\#get_tagged_addr(), data[i])
    * @param addr The address to which data is to be written
    * @param data The data to be written into the address location
    */
  extern task write_byte(input bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, bit[7:0] data);
  
  /** Writes specified number of bytes into the memory through backdoor at the given address 
    * Note: if any of the tagged_address_space_attributes_enable bits are set then
    *       this task should be called with tagged address. Ex:
    *       write_num_byte(xact.\#get_tagged_addr(), no_of_bytes, data[i])
    * @param addr The address to which data is to be written
    * @param no_of_bytes The number of data bytes to be written
    * @param data The data to be written into the address location
    */
  extern task write_num_byte(input bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, int no_of_bytes, bit[7:0] data[]);

  /** Reads a single byte from the memory through backdoor at the given address 
    * Note: if any of the tagged_address_space_attributes_enable bits are set then
    *       this task should be called with tagged address. Ex: read_byte(xact.\#get_tagged_addr(), data[i])
    * @param addr The address from which data is to be read 
    * @param data The data read from the address location
    */
  extern task read_byte(input bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, output bit[7:0] data);

  /** Reads specified number of bytes from the memory through backdoor from the given address 
    * Note: if any of the tagged_address_space_attributes_enable bits are set then
    *       this task should be called with tagged address. Ex:
    *       read_num_byte(xact.\#get_tagged_addr(),no_of_bytes, data[i])
    * @param addr The address from which data is to be read 
    * @param no_of_bytes The number of data bytes to be read
    * @param data The data read from the address location
    */
  extern task read_num_byte(input bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,input int no_of_bytes,output bit[7:0] data[]);

  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  /**
   * Updates the agent configuration with data from the supplied object.
   * This method always results in a call to reconfigure() for contained components.
   */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** @cond PRIVATE */
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  // ---------------------------------------------------------------------------
  /**
    * Updates the agent configuration with cfg object supplied from agent
    * command component
    */
  extern protected function void vlog_cmd_set_cfg(svt_axi_port_configuration cfg);

  /** Puts the write transaction data to memory, if response type is OKAY */
  extern virtual task put_write_transaction_data_to_mem(svt_axi_transaction xact);

  /** Puts the read transaction data to memory, if response type is OKAY */
  extern virtual task put_read_transaction_data_to_mem(svt_axi_transaction xact);

  /** Gets the read transactions data from memory.*/
  extern virtual task get_read_data_from_mem_to_transaction(svt_axi_transaction xact);


   /** 
    * Retruns the report on performance metrics as a string
    * @return A string with the performance report
    */
  extern function string get_performance_report();

  extern function void reset_is_running();

  /**
    * Gets the index of the FIFO for a given address based on 
    * configuration
    */
  extern function int get_fifo_index(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);
`ifdef SVT_AMBA_ENABLE_C_BASED_MEM
  /** Gets the handle to mem_cfg */
  extern function svt_mem_configuration get_mem_cfg();
`endif

  /** @cond PRIVATE */
  /** 
   * Returns the name of this agent
   */
  extern function string get_requester_name();
  /** @endcond */

//vcs_lic_vip_protect
  `protected
/B@D-b/L5LMG#JE4(^\739Q6:PZD4>P7:2W1L)UL09O.B5WFfX?5((B8?-8+?<HS
UA2;=d,BNP;CNa;E])0d,4-8ZYGI5a6<:X<O,e;BUCNNI/RMQS]#+>7AZ]2I3>ER
6R8K:Zbda3V_2U/?Q30H21S=S);(GLBZU<.e-P;5)^YYc\3JfN2IPSX[5QD=;U,X
RF5_aGgXN+IT]NWU>_U=dD81Xc,CBM#Q//_7S#ESSVQcD9QC8J_a>\_(@(RX-II.
FcPMfc=Og:V=_?U0?\KXN3W#^Q5KWYFW(S-de;A>ON3<G9_7JN75g<\GW+&#:1Z,
C4BCb1Y)TIA.E#W):f>F2>+09)23(Dc;YEg0QDDNPf]?_S<Q6\(?3\&X\_I-(=.=
UY.DGI])UF4RD@PW)=UfT.B&F-G1O\DAT;=7V4NTRW]e#GI,:gbgG6K#Pd+(?EN5
L6eKe=K9S)cH815eEO<54eB&5$
`endprotected

    
  /** @endcond */

`ifdef SVT_AMBA_ENABLE_C_BASED_MEM
/** @cond PRIVATE */
  /**
   * Obtain the address mapper for this slave
   */
  extern function svt_axi_mem_address_mapper get_mem_address_mapper();
/** @endcond */

  extern function svt_mem_backdoor_base get_mem_backdoor();
`endif

  //----------------------------------------------------------------------------
  /**
   * Function to get the configuration that should be stored for this component
   * when debug_opts have been enabled.
   *
   * @param cfg The configuration that has been supplied to reconfigure.
   * @return The configuration that is to be stored.
   */
  extern virtual function svt_configuration get_debug_opts_cfg(svt_configuration cfg);

  /**
   * Function to set the port index and port configuration for an external agent. 
   */
  extern function set_external_agents_props(input int port_idx= -1, input svt_axi_port_configuration port_cfg);

  /** 
    * Suspends signal from being driven based on signal_name value. 
    * That is, the signal will be driven low and will wait for a call to resume_signal 
    * before it is driven high.
    * Following are supported values for signal_name
    * - awready     - suspend the signal awready 
    * - wready      - suspend the signal wready 
    * - bvalid      - suspend the signal bvalid 
    * - rvalid      - suspend the signal rvalid  
    * - arready     - suspend the signal arready 
    * - all_signals - suspend awready, wready, bvalid, rvalid, arready signals   
    * .
    */
  extern task suspend_signal(string signal_name="");

  /** 
    * Resumes signal after being suspended based on signal_name value. 
    * That is, the suspended signal will be resumed back and respective valid,ready signals  
    * will be driven high.
    * Following are supported values for signal_name
    * - awready     - resume the signal awready 
    * - wready      - resume the signal wready 
    * - bvalid      - resume the signal bvalid
    * - rvalid      - resume the signal rvalid  
    * - arready     - resume the signal arready
    * - all_signals - resume awready, wready, bvalid, rvalid, arready signals   
    * .
    */
  extern task resume_signal(string signal_name="");
endclass

`protected
;OcNCgV?2[(\8=OIa#_Eg;&8@/F1Ta?J[0EY73W8Y^D:J=68TR=b7)W(]VO#X3cb
]d8NcX(B<5^R(9TM:WGCJXQ5HNCFUE^)B?>FNKR?f2)ZHR>KE_JVZD6\YP3PFY8M
EZ:2P::.fF.6RD57ea[VFe1VH0D[MLR3F&+W>ZU:QcRQ@b(=7a6+QWgE,A)B<_K9
(W+DKGN&X+9,U.,\Uc.GIF>D;Qd7>ad+V/6a^a&Y,PNY;^+?5>CVIQ-5e=2F=P2S
)&O]UH&e-3+,8fD0g^<EQ>1<&6b1B1).B2,+PE5FGP1Nf:5I^M1IO[eXg/bb@=;C
+A6+#(&KPFUF&RP\UK>W]@^Hbg(,]:Q8bbY1a)e.JX^Td6WIR07\-9H.H.(LSIXe
cd^ZA63GZ4)MV?>.Bb(a)YU^LLZM0JZ5_#@_H>VT?=R[e>3#6Qf_KQU\P-=T7NK1
bM/AbSd//=JZPTVK4TZ@=HJa5M=<:ad43BZdG^aRO1VP],P[>(AVC+dEGHHS,[,T
($
`endprotected


//vcs_lic_vip_protect
  `protected
R;g0C2UW/@G22]5bQ-+4&D?BR7X\,QfKFQS1[I_+3C1EJ[+HGIW].(U4VLZ6ZX7L
V>8P?CcJM>)ZWS>F^;B3KL].EeP[S0O55Y:1D,Te-X)A4TP],B1#bG8]4XK;+457
EfRJ53[V2TLSB\-P.V[P=D(T:LV;0]L::.7IMfX,E8LXfYFHTM#Za;bN.[@\=gNa
bO?fd^R-+/I1eF[#aAKGHM?93Jb93OEQeW_6AV0G\36Yd-Je34BLBLbT4?2HaV.=
BU#A.=4KYM#TAOMJM>f1N>DfO^DgN>BaLfC\T@eG^8&0#W#=E6LF#/1K4MHYZ-S,
?HK;38#@3-3?>^d;f@,X3UXK6TQL@A]25f;9R=6XgC,<Q7S)GV5;S:-.W)XZ_5Q9
Y0^>Z7AY^HZ66GDWVXPbEdP7U#J+/WY0cd\[#XFY&Q2e)3(Y<3A&aa[G/A?U8WS(
PMaM0#8?\S9;BN7\+e(He9<LEW0AH3>0I_^([OWSTK0W[R;3,Z,ef6e,9:0>^a3U
5e5TA_..X+g];S\RD->M)3Be#Rb+YJU1M0fNB(LOQ<^:HY4=(I-B>9.F-/[<d>KP
=->FV]=<ZQE>M2])K+<:\(_N0-?Xa^P79(YD=+>-9eFGC]G^T_?gT5/^6-3]LLa8
)2SM^,S-975RHE[<74[(7P?YW(gTRdM[aWNV+K9;0Q&EV;E?Sc@/3PS._e45dc+I
EJa@IbH).B4?UGH-_>ODc_g2bU#\:DI&dQfCMO2D3/;Ib7c[85-9IXFTb,ACTJMJ
9>=b5dKL(Tf-<2QabX^/T6F@L.ee,;1(&CKUHNZF5IFf_VP#4MYX)FPa1TJKN2Qd
(,D@gB&1#7C/2[TZ=4OffCAY7EFe<(4QD&UVRb##d]@K)HVXOb&W.fNMf9aO1?9E
=XRB\TcS.,g[3]5K3fI[H,gDb8A)Q7L2<W,.\(Wf0S=S&5WGZ-?6-#(,-_.5c,SH
ZSMF/:>YT.Ag58G_VBX4DGWGZQCf\M)8RTIXLF3&Y<0W:0c<EX1b,]b20&@#SGX,
1B.EFdgeR+g)8DI.6-<[2B?LZ1\eHIeP]Od]eATgRL3,^FQ#)=AK[A(0d@]UL:.<
Z@INAIffQXF+-T^-FRGU/cOBYgcU2XMW+F<&J##OAXZ2^W;+4N<4fTgV7+(&O=XS
D2LGS\7JGCdGMZ]A+)M]eR+gX@/9-AX9;+b#W5WQ#JWJ_@I&NTgSS&O.IC<V5&A[
]a_+,a8KJH6P)()4B548e(c/_WT?SN/=/Gf7161J#Z+eQ<0HI.28F/aN^>8LZJZ+
7O_]dJ7D-647cE_AGY_,:.FZ>2E/DE6MD+\Fc3O17E+JgR.eV4K4;]^B4G+HJ]6@
2_ER)=LWYTD^@9P<=DP-DJ+U0__f?INe-I0cD&-Gd=<70BK,>)._/SX/NJC1P>T.
J.NEFEdPOTdC\JJ2^b#1SECR[4ED+TXbA9cfF]A0VU/&38EDJ?IFL)JK^@b>cVbX
YVX]5f4.FWA+#T/>NT\SA^Xc1[93(R>^UQaM9W:HI2^M_ZX>;M#7K\)RWYF&2&,+
4P/D4P7=N+:PC\B>C_-\D5Hf8KJ[H=4V;EV[cF(\:5gS_JC@AVJ;H#DcC:UdTY@R
;&-Sc=-[/>042&(\OL?5GMJ/_HI]f/Z0#T0P5Z]-CaZL[R\HR&&=B5C2Z_?1e@_3
O+e;=#]Face_-SOc)?1IOFC]S20d]Q9&6.5CXTR;VPY9Ka<fHT;dZ8TG#6_f]H&_
[GX-K76#XI@#[2@L(\7.OHbVO7bbFZ)[76J>W]6fHcO-N>U/UdEFL8=E4RdA?)aK
J=@M_PgCcH/>;Z1f?JeR>(,EA(.VP8.I)(Ra0]TdE5NZ.bKU?-X(DWLS9>DIgU9D
@<:GP>/VQERM3f.2>cY8X9(4IY22N/RcS[WEBPafVD&KRJPSKF,4G)ga?;c:4<\T
JALY[O;M#OV?GVdT#9G5ZO)-U/3Pf:B?W(IRC1PNM=KXL&W/WFK-.+_Q21-bYdL-
\3Ef7;2LY2>C@0KR=:(/9cOAY&PV4E(O#EBc.B#HR35C97^Yc:P1Ea\5X=bER<M#
b-[e3cHd/;N,\;b4a5)5YDSE6NOc5C-ZIB)]^1B^)ZJQ5_0X1^HCYW4F=DN3bZ+0
T6@XVc3L:WL@S5)>^JXODR3OP))4H>90-Qf6.27JPQfG=#Xbc=YG<(c0RILFf<SN
-QL_\9Z,/+=>^)5I8(U17/;4<Z:L9H^EegML2)H5T]N5X0gYUR^ZO5CeI,>8BJ/]
_)2A6U?eLb5[OX<)dI_H6?UGT1cXVH8(YN2841O[-^XU4W;=L\a-V1JOWAWSH80>
.0P#&]0Q4TQ^-2^K,9^Z2DB9S8<\_UD+N]+aS?STG[5F2,M>8/.2_eSLUK^XUJ-C
;KR:50QJNR,DQP]Z:BKD7YO_O2\.f-WVCRO0_[N2FM/FQQf>(#EP,U?H2FU]E<](
6J:+ERa3B+UeD4S@;XK^bIDR2@_@+NO-?:2/E=42>CE:.(?\P&?(&A-E45ef=Gb3
D&]\VWM?L]UK1L=)#a<PTcYWR#fJ]U:1=1_9&HI9S9/G@E9ER1T\,OV6,I=VI.?/
MAE0J5;AH1KE=+F7JBU0;44HE53XA\TB.=S.bWfH;@.W@&GYW;8J(dQ8?5PPS/02
6@Af\/&>LQF,LDAYOMe,P9MVDSOB765.[U3E\J#1<T6,/V@+YZf4;5AZ#;7Va?ID
#JA@CAZ8CJ+VE:,T>Xd,BUVPFJYOc(3H(;8,R7[>]&U3?^\WT+<:T#S)0JN[I#6Z
DGIaV?&)<bYELS_L5?,=_+?()TOeI+fZ_Wg#<[8IQfNfbL&?>9C2JF=XM;WcKU&3
5dP196a]B?cC9>V@eIOP-2ITJ^ZMPNc,<[L(G/Tc+Wf)<QJ,>MgCC97[XK6/1(L2
W/89ALE#FdBE[ZP&Sa9ag14Z8g(R&I,Cb6T[==LZUF6.J>ZUGa,^?;7L_;F+\G9T
F2H[gT]@7,5_AAa:AU_H_ZEBHY>14P0U()59c^<R.cA@&/#,IN3C<[A2GK-+_L=f
V+_UPf730D@8OeY=eUQS(#\(Y8/ZaZB]OfG:f9W;WJ<TCC?+9]W1b<#Y/.>&KNY1
XCf.A+[DJEJb@]cgU08V0f;W<fV486P4C?,4HU/Y?5aPLJ6(eeYBE_@_3#Z;KCdY
39=+4d/()V3)11cSTeN/M;JCF\,35T&S)VQJ_\b7.YME/@.MZ5Ab>E9#-GGgUPO&
+3d(/Z^,GT1MD?YSOC8<#0D=@AI]+H66=&/-WWe[J+[&\PHd(]OM-Q1698a)ZS4>
MCa6V[4==;Q<M_+SP3&6T[86Ae,U/2a8+45g+R^f?J@T4_<V\I1d]P[M]g__90>S
H/PYaF,&8^_d\Kb^0cf5]U:H]K<[(/b[HO)9#]HQ>7>S:U&PS.^(++EL?<#<4\FQ
B3cK5IZG_;.DF4+EW;1a.#C26@9I+ffNVVGY1.,H[_4.c]Y47QU?.IOZee<954/L
9=c&eWc2^dLPN.e7+2]bRK+];98)I>Y/BY=;N2P<V>_EP).;9^fcUHP:IY0=#+=M
K&#KBYDaML&,@=L#SC2&7OUHRbd:@IcF/KXQ3@d025=\G2YR(;1>W?-_-/X+B20L
.DFJ]?Kce=Z0HO1J#MV1Y+-7=OMX6KS^]YB[GN8HMNN?=29@e6>CX&?CL,KLV]/3
NF3,BVb4KL;:^BC5TB<b=JD]4Z;+/1/[TedfdLI>S<OU#fEDMU1G,b)RQeR(9[21
T.NG7/?+93D5<\EHX)A.SRE/KV0/IU@>E_;a7+]c:9XYIQ.PVYYcBDN[E:CXc/Xf
C.9]EY\9Md=U3)7/+9D5f0O]e9.#K\>=XW;[+#[fCGMOf+d=1S16/_Z8J^YSb(6V
3L6-K<.g]&:?BNI4V:],NZF:I.]U-U)DU0H?O+ULbH.DNCaEZXTP6L+A+&_MAOQ5
;W+e7+:+(C<=7OT;:PD.&IL]b=_=U@&#Hg\0)g(+W/a6).MWP.>>JWNb;34AGe.G
))_D_19UBI,-d?<JS0.aED5bIY.3=J[TBGY&5/W(YJ5Rc1.8dZgMSY_WJ23ZA5Ne
)#KE&G2:F^+3#]I5.Le([QPG4\<O5/M2e+TeObb^#c[:,b5](I]dd]MYQ<ZBHe;C
&Uf;(:SJ658MK]Y?U=^cOCZ\8JGO.&d:e:D=b5g-QYLIcPHf&QGI^LJ5^P6BU0KL
e:-VYL6Sc_RE&HG6[TJ^NE->Oc8]26(\>8=O?)XaVZ4+^aFH-7AF_?#B\F&:1fE;
O->]JQS1?e.AZd[(Q(J@_;-,#baJV_C@AdZ@EV1KQU6@238J&9Q)B\E:JMWJf@;2
X#,9A49TgeA:?e(:R@VS-f2;LLRD1JN\eb0DEUI?J&gR(N5R:9OA,X>JI+Ab\E+g
O.SV293-,=DD-]BB+]HA(c3bYSOP=6;.Y1#=R0DFDFJ;Z?;_4cAXc0<P2[8.f.FO
79AGODQ3^\KX[ZR,eDPV.;E]+APDdOXZ&445H22I5F(ZN,:3X8ZY)cG4G?;IFQF=
A]MW97D0e][34<OHJ[677(P@@7W5MYB:<LEA52ggT\fVHD]SZ]a_5.KDaW8Dg-4S
H54P_S[BHS&2A<I0<;5:bC84K>fb<g2b#U#P-9Sfa9J>:/X(3MJ,#RH,Y-+4WL9Z
+)[W7^]G<>2P,V7J&FQ7CLF.+X&4I&EFXFX4Y5Fc5\c0?e,Z/6&CNK6/a<879NP,
X;X^GITRY#\\_3<GIJf,\dP9:\+5D].L;QG-[ON.(A78OJ(XfDHUF&(PWS:6;2UL
[=JRYVAO6,KG<O]c/2Z4gF]_V@aYBe_,R1aM]@P+&7)XJ&e=GYY#Ze6.Z.(2?^NV
1LKa\N9=QgHg)\SSX(N/C(V&^O5M]^FWe]GCMZY-fbY=A.PTQ7Q<M#=EPH#&\=2K
V,JQX9[//#?bS31(P3635G\f27:BA81;U\XEZP<2J>6V1V0HZ/JXU:S)OU5M]6U1
+]I&<<?d.=g6IZ2f[YTJNb50L??E@dV2M,IU[dSQW(\NJNeM#+g<^NUP]-O<U,9>
YOAc79UcKAK:>@V>7E+E)3XSR/70]_5WTdW()4aW,L)YG-AYM,K(aJ/4F]W6e_a8
6]Q6R_8[fR\<,@JO4f?/8<cL-dG\2FE<@<g.=RPQBR+L)+DL0WWU^8^BRNV-/_1A
G9AP\:^)/@KMgL?TO0+3J6Y=cIea?Ob7BCZ<L1(TA]BQ=Z_4CdXLS8d?&W(E=6/G
]P_#;WP@2@W?#1G#J17:.7LDTCE\[B,GJQNNVa4T[3T21R;K/I&4G4N=d;bB^Ja,
QGHY8\8CMXN\-R+_4^T?Lc>264L8Bb\XgLX[4#Mc.V6HM2fG]?266DRJaP&,YKX-
&809C8&PL^0_SAUe>0dK.&6P@=(VB@>EVDC>L\^?TYT@H2&SOEIR[K[;KVQO/Gd(
R)>/:2FB&P7=a@0.Gf][<>PQeBQH=QHE6X(#_e=(R,HO:RP9Y0c>86Of1Y?bIAQJ
\>]R7K53ZG,@<dbUYV8.PL5gOd,V[c_dV#(a^O&@(WDA@#FI>A33C^g2@H6M4;=^
]H7g)dc]T)NcgHbQ::a6:.NA3?AW9W>]L@e76(3N,H5_b-;L2F:;@Y8R5d)TTHP?
U_4,<CGW(a0Z57Y<Q/DFfbWBdef2be<)#BU@^+@Fb]XAV7(D2-/4&TKTZ1C0YL]5
7WI&aXF4/6,V:X1ZKQRgK4G\1#[EO<-T?PD0X37\M3=:O3SQ7;H(0e4P&J;:Q[XH
-;+ZLF;7X>ASY0))WZS8Vf&f&QQ=g,V-g1(R(Xb,\gZ+Z^NO>B,(aQJ@H[LZ?5EU
0(K5)B##H?KGMU9TS\<a)e#D0+?2g?0=,SM7:=WaNEVK@&,&XU(]KEUC57@g?:OP
X_NI<-XK:d_#FY7AC^D5&bF.LMT)&K=HP:Gc2Kb?6.VA&F>(JR:4-8W9CZ::4C.4
=3-<b@#@[a.T)<G:V->IT6:K-1I)_@<Nd2,]6TW^O#H2T;?IFe/+^eX;Z+(=[?g]
>ObC@/D8@C7NM2_0(_G3>/40#A4&T(;AVFU)/=f.eVYbdJPIAG?Oa@(4W29CJe(A
>WI4Y]H\#9SR@eY\J1I6PTQ=-]F/VY-/BcL_/1Z&;O=#E,XY#L\<#?UX23_/fK>b
+ZHbKCT)Bg2F#W#,TJ^Q-V/K7?A:e9V&OEfIU8N>46#9<9[;_^S#bPGf;ee6D,4+
BD?XM>T70E,#J#<O<+9(dYUJ06>Z>c=#1[OJRN0\b^\,]2ATD&QF6.]e@4TNZF^]
#<@2D]4:@8Z5\>1JX]TRLR\6E-H&PICS7H,ggb;([)bC&CL1/K9gW@]_99T\]VeK
H6^bCUS;E8?bU@GCS4g9DXCP0(D92-2TP;P2\f@dK-GNC16&BT2NC9ALMAK80R9O
75NT](.dZ?7X5[eUg@S\NEcUN+GgRQ<A8:[7Jg;T_TgDJf#a@#ga:9&IgBCU0P7F
QVIb+#<&>@bO=G@81;^U#N5Z8d/XF-U7XN&,U@DP=[F+&a&NYYRHR9>G6F;FQ8/O
>RH9-LS>(5(aA\+\+_&F(.SIS#L)-N/>)f194#bC5M[_@_44gW5]e1.03<52a\gC
C?J(/S6N8(Rc<WYb8NF.X:(I)gaT-#+484ARRXMC(:fJ#(TSfF>0;aCCVZO6VDD.
19bP6&T+DS63T\WE>G3,N3D+T1EEM\>3XbcONEDHMZ_TBRQ)5a)a1:UgWQNH(R6d
]<@&gHQRG)bfEbfVV-2B9BaZB8/^6_225a.JGg9OKgHXBVbS1GDDV#2agEXc=J=#
C/\8LHZJTFc5a./=AEJ57WXP,ZG>>(c-Nd537#JVO/R=Rg\[@g@FS/aXQWgOB/,I
AW#X(#FEd#f&EJEIIf\50_J7e3<PLS8_NRP;6f6F/I]]KNEX9?)N4)?H9T<;dU39
+d+7(JXTD0(eQW)IST1?T;DOWWaNJF\a,VHSTLZSBc.O8>1^57af:bLW1=L+S9A5
S:@4e&QHQC,-SO?8gR4U-:&<aO&KO3f4L;@56UI^=aZQP,+;]).NC6:&W=EO)A;&
DL;M,M<05A6+aOMJ@JfD0AN>+#^4;I?K&TO2LNBY5)6dL/[e_^8;6UC?gZPMV-+-
#4?5:)).(FW\F)7YQ\GRY^7)9/VW>N8X\_YFdC/?+O(P1dbf8F;d?S8JV^,CO#U2
fD+e(\L>4O]EU<4QMSMS3JeTF_2:SaBSO<,O1LU9/Zc@8-#KTBc2N(,+137KZM^1
b9eKRf055A:2YE((QYBPV#>LWWA.Y.Q)(BAX3QT8JJC&K5Jf]2)N^5X/;\\N/U)G
.EU9c0?8Ca:XJbM<dR^fW+=U;0XYC8U]egOA5)W&>X2g=HOBMf+H&-P<W:;+D8Y4
<@E.1,e&g#,\V9:=SCQ(D7cM&K,&-(6d6FY]&.SBB:#&Z&0BR@e).#4NfY44/=P=
/bP/.C&L;5c;22\eVY?@g\aF?.]SF2]B)]#S7bL:f?&,@1NL=V5:@P;#&FBQNV)+
ZIP+_P@<58d?Zc-;a_73TKbQWIPIH4<IH8A31>YE:)<O>L<ZQFMUJAAc=MF?\=[V
Pfd29/[0Se,Zf:d@#V.92>eGGaAb\2f4/@HD5F,.M6?J/X;2DA9MY3MY8(^e&67G
Uc6XLS.8fP&_G-S[d>40LM9EE=..Aa(Y)L>\701\XS-8@<AK\8&KG8dSBZXYD#K]
&8[QOfT5];;&:R<MJ.aYZR5c0aX]+Lg2V,YY.fA^Z#TM(BNK07ZRGFaI74@?(U=g
T6W:#XcC?fYfWBe;UPQJD1K5HFO0@P#8NHJXX65W\Ta@4^bL//;fNg_JPAcB;VBJ
]YNcQ].N_-,L.PU#e=@OA/ZIc)_aeAVaOc-3fFcC@Q<VeKGbPY8#I&5/25c9-WaF
d/#X,X&TL^=XZUQ#QLR9O_QbD.KW#B\>eKf:-[F:EW/KI?[dO?GK#FYEMgT,]1f)
_[S&Te2Nf)fXdaP\97(LW0C)]LZRCD>bNZ:RL?8J,Y6LLN]UaCJU.-S]8-[a?-e)
]?;<2bP;<8=&;gK/@8:daTE8FIg.-:^AN^ZfaC6(&0A>BPZK=&906b6agf(bAFX?
b=;KT>A6YIg8UV<4e9RQeW]&<NEaZ6[TLMGM;e>HUUMY11?(4NZ/c8Oae+0>PB[P
HUSaVe.1L1V,-L3.e&F<>+.>CK-C5XgO+&dO>JJ6PX+\)UH64JNQUAc1Z9?&;GEc
(,:ZT-MMRb;-f#:8DB1@7YI:FdF[LeJO9X5#SOJ_W(8Z=^OJ]CP5=Y&dSeUO1^G0
.HZgN&>@<GI5TAB\e@6DH,(\B8FcK4ZA=W@Q&&MX/G5MO^@#KQTEM4GO,M=PD][I
\;V-==_,dDcI;8a]UAA(],67C1MR85VZAHe#NdWZWSYEQHQ&eV=;b]b9U3D2(:HE
4QGVg^M@-3@N8>V_F\J,HGGYF3?@Y=M1Yb0XdMR0YHIX/96@AOU4@=H0aBeg7G3B
O6NYZ:e1&6.)Y;5b1UYF(_<BYYHgLFXXN.gW]^BDUJG;E_[7.AL(].:[.J/>7Wa8
)MB.2K&[P@<R1YY31eZ),4LaHGb>&5ZEJgU)<A8@]U8D7X4=E=WMdTSMX=P.ba5P
\,K+K_O6F_Z;,HSD=U,4G#cD2N1B+fdHZK)dPgNXQ=gI8KeY(-fZ_1<;N:BFg&AF
^\cUX_fecW<_fPR<<DV>8,[_R;)bK^N#;/W(@31F7JU5I9PUH])+#+IBG>=;+1^L
\XcHF?F06UQ?_TH6<I2K=43R.+c/XOJVZE64g?QgVV,9,)#X:R2CE6;359G?Ee;;
EVM#Ig/L2c<g>.2@-&A6_[]#d8P8[MZ.6d4@U&BLUc^5c1Y#XCMA>fY;TR1A.Q^)
)XDMb/&B22E>B2C)(MJQ;&VD:;Ab+HZ)Z3_3&KN&345^7fVa0)d@ERXK1RP<2\HN
._&924J1XEWbDF#4d.dJWSbC;?S[1.\I/2gXP4W/&T^IMX)0\fc5EF&9#A2D[GbK
L6STXR-GDRgVATNPAP>6I0W^6N,8#M)?&3HE_aJ&51^-/c<]-0XH6?(J/MFaLg]/
)]O=[\(;W_5)74&0eB_38^P0XMWcgAO[YS@9M>#>gBc.6aFeM[>W36e<+I<8OGNU
L6Aac=L47NV5R0Lb[J=,.<OHg5G:TC6?,0VRB,U,cdFY\8d)+T6AMJ62OO=<[T9D
dWf/SN__AE1W;_][4;8cJKA=T#[-8HbBZ@?.OQK(E^?>9[AEBSNL+29d_5[3eD\_
[1?Y([CSQRafE\YF;Yc:N_F^<(BC938:0ZfL,_E.:+\?U<)V/)UG:?5X_5AMVG/Z
5BMG2G<_8-d1M^a4g7][SA.0g:1#.VcTZRY<RP+?WS/>b6;>YACa8aaZJEOVLCK/
2G\BVSAF/+NM75YC,&.7:gE/EK4]F..>(4E&C1#\aLTNG0L68C;g-[,H0d^+1815
K8I-Z2f4=dG;:44PV3f>@ZT->ddDPK@<N7YS)<,^@93AF\W(IX)WQePb9#Xd/@LK
5)5c,I5fI0Q>IO2GaA4.e6Y#P;<KEc9a=&M(&87]_a)0M5BMW>@ZJe)>.>T,QYBH
)U4fI8\+<]U_GPHg/g_??)=T3SY1YD68;\B_-CY>c\S,V1#gL#\GNV;8#)Z.gLe1
Z:[gR:aYAJ\U(Y;BNE<FFgPc4(T&L4F\^=@LM]7R;4UKNA[:XUeM\VbY0YP+#Y-R
S2I(Z=b-J6;,HBB0?WE22FgPS5NFMVN;70SZ,gAI&&C5-0G_=3(+7GGH6<cg,:G0
Kd\N@MUZB/3e0AQe:#O3Z#C8Lc)H9[FLbAIX9MBf1B@<L^g3(0,^eE(9fKf#eH=;
DLVP>g_9KY@7#/V\A<<+Q3H6+RWVdQ<4c]-b(>4DadGJVd0.35&[gFO]CXdQC(1<
(6,dVDWGTZa2L1[PIgO9,4E5P=]_:\DR@7471(Y[)P@Gc8,AUb5VFdO:^Q>>1QaB
7<T3IO#-FBCB_#EA[>I>.ZGG/EUc@5ZJ]O9a;I,2?:WE@b8WbV,Bc4J0G<c[1FTG
2M,dW?7f9:TaPRR5+d+25.Y;(-e[C0c,:6d^EeD./R0+#<T8EOVcKHEa-ZFD^U^:
O/BXO+9C>LI6D(Z0=UQYXP<-YK@[c<<\PG2b&W?_,NAa\V^M#)^\(@Nd;c)3^6+\
1c3Fg:e#\E]_LLdd:&aK_IR]L>,1aFV#4d>IVK6>G]#5LE+44N8FK;ZD&M9N,:J7
2OA60ZQaJV&dPWgEfCUG^>:0N-:Z[c,Yg9Y(C8bVF.N[.2A+-bgffW1JOC7DY,>&
)fWfTFMN:5N^Xa#=VUHd?15g2@)gR>,UDYF>4S&>Cg-OG94eGX22PH+d2,)3]QNL
@S,=0+&U5N\8aYSeQ4,_YA=-(N=PLgB/)aO3L]>aJ_U0ZE:W&SfS/^R^^/T9>75f
4)QB;W.WFcFD\e8MXA0RK&QE>-aVYI>UI>HOX.^f<;4<AK(cV2fbS.VX.;7TGNGJ
)aeCIUBY2]<RW=WA?7Hb67GT&eH?_:3SG[bFLNZKPO<R<,SI.0MBAU/DZU4e)+EY
X&,@aU-11KWa_S.&KSQV\4/_:7KAQ1b+COP+7EO3>NI_Y,#Z_f3?8N^]-\6QfKN7
e.g-,,IU4GF1]cO73bQCddQQH\eHcO)WNgXN:FWP3bCNRIA7c^Y<;0IJI,WY4XY7
8OB/I@&0,GX\(^/MG3e_-.:[4\H7FC-?d8bb:).@8T2Vc@NaL:eR^P)L7;HJU4,@
)>6(?/;QadPgH[d5<9-CU@+M?&Le2[]UVBAcef/A5g&7TY>RT1AO^B1Z_-Z-YEf\
?@<1IVP;J]):7S@dO^)U@+U?gX.)[?EB=cU/-,1OZSK&ZZ]>@c56dDWUg:MR]#R&
)2\b4;,gc@1CZd&d7b7(<D[ZOQ\6-)BTZ[5DE3P7Q_cG\B[IL7=/?N7SSNU+[5^[
GTLQ;[-/Y2ZJNaHUeXP(AL\8,HV6QNTa>608?b:>.YC_:R)c?CM1Y,eRQ#cbg#bK
F>(S-853\8<52/_6P4-aMEX/4;OH.0bQRdU,bbJMII/QI5\/8adSG3LRUE>:c98F
OV1W\(eU#&)FYRS.Uf+S>,&&Ifg7/S93_<L0_JU@)Ve/6U&b_K-I7,_Z?H,HD75U
1Ja/?D\;gB-b@L;>5C[L&CXRa.fX31/WIcE,^&_O9G0TXQDPXc^G#[ba/11?:f(+
YI4E24TVG(6T,d2X9-?D_eBQ\e)e5gWgAS_YX:3S23?7/G^b(Uc:I<P2QcN:N_J8
cU4WZbIA@b#TQ:WA_R;W,9XOQV/U_dS[gD@Y-_\0a.O/EAN3?[J)Y)#;QMeb/9,P
SR>+EZ#g=[&5bX8X#a(MAe899=G^d0O8>7WVWPU--R(ce1\\DW+Y:43#>S[OV3R?
.6b0@9Kf9OT80&,1LQc>e7gAHRHgd0UJ<?3-UTaJIR<?W&@PEgZ[W3A-b5?a.:4A
=0KY3BM\-91^U?V.-)G;da,\.HX1->,R&N]J16R_>KR9E46.U7eE:EgXUONA-@C2
8H4/V^Eb@,50ND.@?5M.,OU41K&Gd8<Y(3db/+XaJ/<B+,#[fQR+ZQ=D^Og,&QX0
R/f7CB2bI0OQF+328\fXb.:+C[&_EYW+S#@2gLOMFCU\)<=Y^H.cfg.bC\b+DSHH
J#C.(4O-GNDV9Rc;3/?/f\-6.8^Q#633L8(_=\WEBG3<^LU=YfM^dT5V@E<QADbJ
SANH,,L;[+.HY,df8^)7ZO3@B^?IZKIEHG3d#ML,N1#PD1V5HD=7,;O2egN3acIS
TA5WP^T8?7)D=YBHQ#,00)H_,NMJ9EQdN@8?3NQQ^T:M2E24HP#Y.#3c6b\SM,5/
cTPL1_Wd5F+&0f)Ld)8TF+F?HLF-C)C2@[@O8->=#Z&1bN7/RJNb3\cY^Z]R8:WT
R)(@dYF:.SVLHa)c(@3ZgW,#./4)@e5-E4FdHb9]+9S(?#9E0)TI>>V\FP_MT-)U
^bER=dYCW<I-^QUR+K,E>-S6>&CC8-;NPUM6C#(a.\bQYK_8gT+._LPL6PVbZ226
+(GSS:?_A@UU9Z1BYc]1B(&-<RVTF4G6DLf?a\\d)C[WM;2QKOQI,)9X<[S3QNGA
O5+T[M8RND]DHC6&TOFb01aG,Ra<;WGb8f68U0>XCGTEMTD6KRQBG[:P23L8d\]a
gI&/@-,[/3J+9PWYLf+aXK)VAYVG-LAS0S#ECA[9]/9b33@db#d&#Z;Y7N?4;aaX
GS)E=X2cZ9X9aY.R=RPe>-S^<?2KTY=T+PY=a7O4EXY3b1A#C&XGaIXbRG+MCaM,
-,H(:-RDD@cA?HfOgXAZ1Y(]0cF&;A^9Q#_b^f7MeRE;\/_D_-YP8>)WdZcCcDXb
?ZQB&W2XfCLS#UJHRLJ_QGd#<Y5&DZe(OFD.2;BT:CG7L)2YNOL^LdPVfbEW@XgJ
8_gJ^ZOITeRe^LY8e^Pf^41<8B0Ddg)&Q<V-6c4d&&^c9HQZ]Yd^;W26bK8,;VQb
)BXKKd)@E^RQ.X:BTP(+/eNQ\EV(/3>QRB5gL5e;66(H,[L4#ZfFG4Ab^d2H&Z5&
M9VTLSD=J1[c3HUN^>.H-6E]DMZ2T(2072,ANeS)DV8IFEQ-9?MQ@X>?OPQ(Ae0,
E2<PR?BO8OVYeM^d0Jbg](CMTHXUVN[e)/7HKMPY?,G7bLRVS<PY\3B.3,-PWVCc
9/&^0C00QJeP##G+3e-<&Yec4cWLS5;NR0[DA-g?YP\Sa#?_NBW1:Ucc-fI53.>I
Kc,1F(PF8GW9SRR-GTTd#3^>[a;QMgO0R1F<J-;g^-@Hb_P#Id84U34JKR69,&3R
QF=X7GAU/@Ece&&-E9Y7]>)&483G\C+,FA-NRd:g@.#(D^#KeM@ZYM0,-#R,/fZb
KF[3;^)Y<ZW/11ZEQQI7GO<FUU[=:,X(:#7cO>1AS&+\T]WTOX-c97@E#P0f2(H5
e0E-I/>bQOK/Bb#HJ\I8OLUgZb1MJ^c?P8C<85d\D6&a^R@2:C.2O;d@]?I9\IR&
7QFe&16KIYFGB0:f2eW^WH^HQOSc@60SNIa4YU.-\af,E1:VM&gY=G;3=)@Z0F^b
dV59(LXG3RgRP@fDD,)ad1d\G;HQdWQ3X3GOf)9RR->Rg@\IDA_,O.6[.cCY&_2N
3c-:Ka@J):)Rd6W&dc7;5D^_D<>6=9S,;Ge3K:9cG<UIAK(E?Q<=gJXWT,=>U1c3
1][_:@Q#)]#aBK/=1Y#CGCE3J]Ib6Mg(3<F<^HI<gV1eQ,B(JNBJ,_,\]W^;[7=^
8@Y@fN0]V]XXQERYg@.MNVN,UEX#BOW=G<3afWG&e#RLMTWSEA:E7c<RKMA@3XW]
XR_HM9PL^X,;_f@[WT\[Y.cFZ9A?H,>9+A#6gWG-G)9]C5UO3a-X#I[[\?>]Fb:4
1=aG2aVZM:fKFPOHE;U#Q_[4RY?T[?;2P=^52=H3Abe]deLLdYO=8cYF5eRecS]Z
WD,R]]PY\Y^HM/:;WO2]=6C;?,7f(Z-A.FF71N^;[OM/MK&:>9YReMSAAMJ1784C
L;[PdK@ARF\>/?MD32OU+c\(G[SP[LFYe?1BBd<_?E6M<C6&\(SFQd573R\(BPV?
<Z2X,I7)IH29aUBRfC]Xa<7=>7RDO[PU2J2eQ>&5-+_Oe?UA:PT.Z<:)E?MfeY1\
IAWAN:F_G-=:[6<\e-ad/g5M<I(DXe@)I&8?6d1VUYCQdT4()VG<YEGf3YZMJc32
_9aMCL(YZ0Y-E^14Q-R(Z@\P]SWa56I,II?b>&U>E-V&A-91,E>(#Z@>9U;^E4(2
:V+cQ1UNbQH^&R;9^3Z&[cJ8+E9/AK=55ag98+XU=-OL1Q]ZfRaKBVT.K+.]3U.P
RBbbAAXO<B9T1#7LSd(0@.PbZKN,_K(M#d.U7O<N31..>=@3.JJ9ga3=7Bbd,^NS
YOJ:&/L;\Z+&F(;,J#-^8QKW:SGf.OR1c9+3]P9&5SKS2XRT2bbS&?I>SN929;#H
Pc9+>ZM@9Jb<U,.+1:4?Hc=FJM2#PbTKfY^:^7\&WSL^_A?#P(;@[C&J:(:IbSe6
OXa+)Q(0fL)=4@fKW,_5;[0QH@Q+(4b2?7UZT0_?DQS2JSO,;PJG7^[X-1DJX8Cf
I:(BdKLX[6c49Sf:C@)S-<J[3H_EDN7<TX&P1BHASNR3]MN\]4+PEWQ]O;MdSF]3
PG@VAYB_IaO.)4ER)J]TTD5;J^1Q,E=-fd^_L)0,>P><,_H?&c,5;E.V(^4/]dPg
&b1J>KcB=BTa@S,(4=-=RM>XdMQVXg+g/WW/U)5=EYD\O,\D_\/FRNC?P@XH:4<#
Jb\VA9/NFK@D()U-@SDFe]G-b?XWM[1;,,5LDNB1TaaD>N80Z<PH.L=-BD5)Ufe=
Jb11eedO]_&6aB18ZX&gR:B73FOQRfT8J+,-P5faSF^Q+bO6[,c.gE1V_e,M8G(b
L;M+R70(WKJZZgZK[=7BYN51VW:=([FXMaN6:LEX(7J_4)<&S.XHIW50/b>0#I.K
[9R3>NgRHaV57]5]_+TW:IIf]P7#P.T(CYV]YBM5-D.-Z1]SbN/\bVKH8dTeZ,D\
^4H&+2<dHfabf+ENHQPdU3F4,&5I-Ld&&:[Q:_ScdV#VMSeO6P6V]CO/5d7Y<eB]
(\/:.TB)7HR>YV_gY[EYZ)+QF8;81&N:5X39CH2#R;KM^1F=;3R0H<N,?5,>4C&S
<G]1Bc1gPRg.dS+>Q03(9;B]7UJee&<F7<.(4MG0^f/#SbP92>QOUPABcZ/B5BNG
B_:YCT7PRT8bO5\.H/++_3?(QX1g)-U3CSHWYF&PO9.c&UD:(SZS__b:VODQ9NJH
X7518>AR9fMXSH51Y[d=+L88E(c&^+bDGb9U5@WMeL5P=dZ#)H>A93BFNMDMP<G\
MAbYGQKO=RW;gbO&0PY+-75S=,AVb?g_g9[0/=I&KPe)(6^[XO[dV4M)Ba>T+(MC
Pf.)dHOAWLe)?.CHX>WLHBQ4.I[;Y9D@[);DX\/?c&GG;=;d,&.gI0He(2cOYTB3
:EGYW7A05L4>C2@F6:W.HNdHgKZL6QA()PS#<L)Q6d>B\[8c.?W<G=[><+A[L657W$
`endprotected
    
    
`protected
UgEaMHHC>c(eCR8[+US,bYDa[VeYaUOF]#49S/cF.SHKC8^=O_(;6)2(,)_S_-P/
RX@Lf;)fB<Ye.$
`endprotected

//vcs_lic_vip_protect
  `protected
I&C0)^1:1]#_6E&Y_cU]?^T_1_dAVO1K,P1C@:6+NAM=-e55FKG+4(KB\VG/gL<Z
JKL+\-^RNQFJGA+L_ERA5g_cX#e\56=&;b45[I1ZOP)GTg9=8:MPd4C[8+6-^)VK
WQ>^#8F@>LCfW_N>ZHg>eD_b&)_:X3,/HQICUH-Td2=.Q6BMJV?N>/5;<gS>SF@8
4KLg/KI^J,EU;&WS3ATUG>9K2/CA<,VfTDL3IgK+I7#a(HQ+42R6]2cS@D.HOLUb
:9&B^B^16RDQU^=(,W[_P_Wf@5)PdMAg(JQS(1>FFC/GbPB>OLZP57fGcZPX@E4(
F?6UgBe]E1fWB5<QU0MSbQfA490YdVg),g5&&KIgC]BP,e&eH7N7ZI?>+bb?A,;\
VMW?Wec&VUI/g_WAZa?#G&AWMWP/.LdD.:,G:L:@=f57C+KLH8;dcWMfBKc:b-3(
f_(H434W,V7PZIJ\NN4&6B=D+N6;DSgGLEgM.,6I;f8RLeJZ7S)LN>S;Q8_+Y&-&
d6]7VHDd1O0Ec.#4M3:,._&JH#WL/LQC;M(6]D?NW/@)L(G3LNG3c8<?:;T?FD@7
-(0(2>?;(dL;[OE-OX+Z>GN>4)?g3/>,F<OeTY\<_,-adJI)aF,&?-[MIRe&\W70
A9,3V>]+N3S9LVA57W1gaM8XKOc)3&FSO.@R;],RDX;B_544L66H>7f[Sb.IT4SA
f-0fKIN;EdO0B;6]XLJBTQN04VdH->5A[I^6G6#\UbQ<8PY&8,,AJZUYA>66;L-P
[ZPQfgH+.OJMSMS2)-36X4.(\5.V,EN&4KJ/KTNF[R&0Od)E9;6K>10H;]I)>\a5
B8I^I03(HJC2XL>;K]8W:+1I#LBdYbe7CPY1PTWPbQf4]FZ\]2VIB54Deed]YPGB
Y.b=7AM.K&;-27bdGXaAIb>@cDT&aLQ-6R3f-c272#+1];.[/P:Xb)K8W>Q>.GdF
c?;3R9_V#AHA?G65-20N]b]&VJPa\:G=Y>gJBaF&fKXBW+NK\c43OcbU.5SDX)#;
J\g>7b,,Y5Kb,>;I#@G=aHcC>H[9VP[C6WU_=bWS3f;9I\],Q6EA:>=18d?.<#GA
Q-D(M@5.62Uc_-DWFT+bV8]#LDePd+0U<aKM+O8B>Fd<XNPI.ObDOXAL-X\16]UD
KV0W7QP8)H5]=:5g(\ZP<1P;2FU<CTG1@3\.T30^[1KUcUEWHJbB9H;/Q-)g&aMN
&.+cZS9faH#LcOF;#AUY35Y<KOZ3O\1I8RHO=/ZHfG5_+0gcKaYO/cR1N9aY^bM9
Y2^=S8R<XA,@=2036fc.G(gOa:<R4KEa:9aBK58CH5gVEc9+2H0[eXE^3:T)O8D3
_]?e@G1Z)fX<8>M@8VP&RcS/e?Y2DOE7<DeDXeG+J9]JQ1dV+T&4@T19P)9B8@J.
-:;J]GMN<G(,]4WBQ0;&1I0W+82@52GZ,LcO+^0bFB2>/D2P.BJXJ7DAT?B;;e2^
)2KXcPKOBc84LAKM.aRH75CY6[7YD4&RfD_-+DgV\f_b1aE+=g;#)dHbB[8J[7O,
S-7UW21IbH?0FJTOD?eOY8&7SVA5,\MGI<8f&]Z7YL1;,<Q)PHd+[@LM[D.\A9>+
/c7A8fEW;4Z-?ff<E+>FRXXRVf:ZP@cFKQSg<_VBAVDY^1(IF:_J\H@H\V)a_-0U
2fE.L^V?L@+ZI007D1b4c&g<AVXQ]8(<T9J2,0)Ld0.RV^?[S#Dbd/bDfC.7W24d
LH#1GN\ALX_E?.91F4)M->>HWK/FFA<3YBa#),VS?I@+V7.JU.Y&b8]a\=bg^QO:
9I3WTU,T+_Bb0+I57Wd?Z8TA2])ON^8D/0TEbQ,+;IXS-KZ4e(/TVcB3@,1ENA7<
+O&F=RNM?2gPg,U_>I&],cbDE@@(,:>dQIQRF:cS6=.5JU6(c:V_\;cBR,36MR;e
Q.34LRS[]Y+R4?_]LP8](b?QHXF21dc7FeSg6_c_6I?a\:?Nb/)-\U&Q\^c[=B-]
.T16Z5HDJYX0d.1SO6462EPR\0.fE/e4ad=1SF2.,1c>AWR2O;U5,a)A7d/e(HY]
^0MCgRNbReX-SU-A66)>)PZQYZ3Z@)b;+PJ\e3C?H^]2fbX3_G)7-L]TB0>c[=DV
J&&Y<6c^X\e@8ASec<X7\gU2T\<VTT3)#1HCK[[PD#e4fD;ZOSF^Y;-9ZIS&DbJJ
Nb4:ON\ESDfaS5AREQ<LfP9?2X5c1T:[:3,KN0d/Fc&bZN#2XGD3e6RGBebQV^G@
f3@=Kd_),Q[&.cM28efVH[aXUGa2L9cgRHWfIQE;#WI9,E2]E6BFI;-5/,bO0NFF
\:<&/dI\RS:I-V6e&TAHe_K-9eKS=eB@5D/[W\5]8J/eOL?G;bM2X5:bZ6(bC&WA
:GN3<R[Kd+cDgCY,G)OU^959MEGc@CJ@ffdf83?HUCaCWeF](H(3^W)K=OPJO0FI
9B,P5,]_7)^E/56:YBY02L9E4cVL:LTSM;Ye6OECBCGTb4LYL1ABT<C]=BW/RUJ>
gAKUO=SIV+WSPON/ST9Y1JHXAQSXYZ+IS3gP8:&_L\2HGCM53[G^3@BQX+dLFCJG
TLMKV#&QR7GC4Ig:2M]SDc6,@\?8Y_O:(0^0LV9H17gd>.TE\Z_QgfWMSRP8\9b+
?4S@LP(F3,?VYfT,Z.KgH[a^H2D[6_6B=49c5G92g(N;P2KHCY>cFTVZc0gP3G]W
U=2?V4TS.KT4+LNX[67PNZ)>E/)Z@Z[38->/SbbPYJ-Ld@38faf/<fAXDY435LEB
(:2\JS-NY=d^/JWFY7N/T9c#S(B#DOQYU#6TH5Ta)/7U\O3KeTZ^,DU##bVMW[MZ
9(ePB4/FZd05Xd<]AY2,fC3=7K0?IgP.bBf7)De(Z?(9aJ=7X@B6XRXJ@K1QY6=:
aFFJXK)3IEfR3DRg:9a?HfF,dDg\M8^V[<A<aO&E2^a1^:Ub+GH4ID>b.ZfQ>]/O
#B31@QAU4CbbNLF=c2=\3=B2ACfBM0TT@CV8=</O&^Q8@81FeDOEgb-<&/#C=4N[
:\f#[@&^@;7FV]1d@dPJ;2O&W[AM/WF^W,=/9Ia;XIGg8B\U@HWg81<>K/5<W<O7
I#Qa4_I^,QP9,CXfM2cZDER8gg7JNLWGA@0:ac?cV,\0g<Q,T:&[L-,<QWDAV[KJ
>/6KdgSgE\EWI#XM450c;)]:M@3<2-4R9@(P)e_/SM<97LaYWFDKG65dcU2\58:^
[c,&35&-=WY>PL4KbVRTaaM(b\Q;B3+eXIJI64CQ0(4JgEg76>WC<d&H=b-d9MY,
^cccS3A1(7MHH^?dS7g^eJWBg,?7_>P<8Y.G_,]L+X3LS=[&;AB,&8UP[JL/D_,#
NZPSeg:SL/Y&\I1B6D8<F?S3I=K6U?Z\U/55aV_>e>N-HZ#_1YAaNV2@X^7MA3//
4f.c7AeX&I\aJ?8FN(YBRYe&A4b,P:J3W27#T\4#aM=A2F@,5PSAf<;_O\97J5#a
YQ-f6gL)ICgL_,M6(f-YE(T\/.SFb>>@eTXR3L;_0JPE61S>VXKB7M2d\GBgY<?J
Rc6I+9RPWSf:8E/dc]HP)G,O\E7,0.C<\F#3?DDIB+>@>,HES5]07Id:Ycg=cLb8
)G-SD<G?HTHPf/#+A,;e2&QQ^+eb5>+)F&]X+O4)&+4:+_^6gY&;bTaX=+MDR9#f
EYN,S[P\OU/OEQ.G7O#RN&VT2/V,IeT)3:YE[;,3O3Q:N0bEY7E:2XHGHCI2[\cY
AZVBfJL#A>)g28^bFJCQHbfO\@EUdJ1_@c?aYg^7,LMP(Z/>MJS9dHE.3[>Z=-ZH
CW>S-EE/V2@NQ+T4T[c3cf(bU5OZU-G>5N:>ZAMSOOQI;Y.[RB,>B3PM5O&##aDY
C0F8Ed.B+R7(I==?]&&4YWW6P\=@d(Q3.fH/IY8McK3F=02B&Q9:<0/6b/6Y0R)]
S4A[<^3+:dSX@_J1@@_;d0(e<P)X=32[@ZaCJ179H9a7[+P;?cHK\bM3S18&K>-L
AD<L(I6Eg>,SDd_V>fCF6):K)[G-@aLQe\9C/BO&\)+Y@1Zf7A0E]bWESEe]HR]+
9Kg+S7\HKCVV);BK3#>CCe1:O7#TN80R\Y:9<?3gF@?ESF)7Vg,OGbef)Ag,L4-.
0Y302U?^De6UV/P^g,SYNL+#,@(@O#EOd&#E+f]]0E1.d,11\R400dSa@PZ_P#AH
=\,S[^<fN@ADWNKgc-KC9CbA1V2QX/;]&?&9/IXT@,[PcG[,8&R_;aX+Y[)#5,\F
J7+;@W/WfKfI^b@1>D<;4\W:A<=XBT?INd)L-\4.[@WIXb[1Q@]HX8//&APe1g6)
WMK/F<Kb3F?=WV.XYCP6,g=X7#Rc7/Q@EP/#&HB#eXG)@6UEB]6+G3]7SNeE@2/;
U\NUB+<Ed+GI(-J;[DG<I4HTf;[=:E81K)[]F=e0O=^+f?d)@]-DV+#<(SD2OBAY
c8YB^Q.dL.ca.:8Gf@Dg5=N)I4,a#A_>g89S1]YU30QZ[;L0[)152Y2O-,)GJQ(:
/:B5_;>0C[ZF2]907EWJMY=^WNN[?/7;OCbUDFF(0T/JfMS-Y[=P7WF0HgOKRY?[
a8JF<M9CfcH,S5e(e?I\-S]?<X0D7;a8)LUe;AMHMJ0G9&;d2HC(dG\Q5E1g+0RS
A_L(?Q&JQAD4;NK3Zb^<R,a[I-9X#RUH[)&f&Q;SI/2CR3I,@FXDRK1a[>e]E+MZ
1R/7[=b?<?.U#J)f-;A;K6(J,dfI&/.;DC(-7EX[ML(7]4YO0Y9>LcCO4;J+X;+:
e]SZcVP;XRL&#0+-EAbSdLK8THW44K[Ue\5T^d=N-cR\@=+1M-;>^Bf[_DSVHDXS
WO;-bH@c#\bI,W=5aa7-(]Wa>>E3H<+<R60a^a,D8+ag\4Y#f58;[XPU5GQ=>,JT
;Z4<P]S-&eMKB&DVa3&dgC?>3;)\L?=e,c_OK3N\<:?.Gc;L:1&ZfQZbWGV0MB8&
ME[?Og#C;(1Lf2\X(>^3YA?Y_g(/CRP1WAG7C=cPGY2?WX]KQb]6FNJG6BB/?5Ra
1.:P-WCK@&5UVXOHG+#DG:0fH/O]F+B59?INK<@OUX\TFH1ASbb?4eIDX[MAe1\f
8?U44>BJ3WHYR)[6O^BAUOO4\_aECN_<[[5Z,6=4J_(D?H5dD]U>NIKX:K_P5J1]
<c0Wfe=YR&?J9a8(><D5BG-8BP<I:/,7dY1S]^C?\)Q>/>.9U:0B8NC:J.Q\+U3T
dOd/B,&FYPWRGN>F,^@]8K3?HefDS[RQ?F&[D,g&H4N1=.)Fe#HARc;&,5Z3dKO3
HA-K(P+,/?VE53dbf\#1;MA,eMU;H.G&c3ZC](RI(aL7YRXH8:;7\[bd\cGVO?fF
=T9]cU,?:DcX)3N+WS&6R=Q;[]A2a3a;[J<_38@/\@\S\e9=N5H2VU<-<T4>([\X
:6b.6^K#[:GeMZ)E8\P=dQ9<)LcDU4+gIB>0B)-fU#ONbVc.40C;1[8@KaQJ^C#c
RD4AOSSB+B.OCeYJC^c,VM3f-T6g@6e&&O(4N:&+M)7N?&URCKD^I3/)^IEfKcTR
Mgf7I:ZZ:9W2,R1Z<6g^[;gB,XDE+AcW/1Gg2^4H+Y)ccP58F38UD[0UD-HGe,JI
<a2YBd?^#UeZ@>W4RI4KXeIF8;5AG_ZYV4+NUdJD<=#b(GYZ,ZVA7:)c+[L@)8C@
14#:./BQ^,?X@#=U-:2gHB5&R)39>^FSY#d<bC^cfIX#M]c#D4V#_Bd=OcGd8S0\
X<&2C2Q\U04].JZY6FU<>:+Ye@7UUPG#JK<d.cFF<f:M&X98G7HBgNSX.#1g0VD?
.6SM97Q03)RfK8:8.G<0/c[0P4FQTd1;Og]H?4.WL0VA+/W11Y0POQ52;-d?<<?>
1=2b\WReN5b+a4_Z+E(5OZ#gd+aM9UfOV8GF4FRa#XX/<?I@B(cX>[8POfN5LRf2
Kd0=(K4^W3Nf4KBaRN_6.5A;B0DIV=>,#DYNWd,M\f7Bd,9a62C)>GEI^HKb,E(e
aUQB=HL3U-O&9Z^3V2,RBUL6@U,I3GdH8Me[RNB0e=1L8?.LJDZf8>O(g;9VBF1V
=55I5S7QH(\\&4ZHEIBV[M_1d:?)8,4TO]:P4]FDP6[-Q-_,Af34?C6XWRR]9[7\
SO\fEBB?2VMAa(#Wb=APg+CBAe#KJX(+C:X7E6VDK3fP2&9^LWJX-#A(KLYGgfBP
+MR??U8LVJ,PT,D]\0&9F;&<c(3\4==V_RZ\VE4G3U#BNK=O61/-TD::Va>f\)a,
5B8,7Ra_U4O3M\5]5&#VJ^d>5EK/_6K;5e_?[e5e(_g6(,K1MZL.-7V-,\;KBSK]
LS54A2&]_1[41^SK+^4>L5AbVZHA<8B+.g(>2>,e?dY-XY46F;g(Tffa7T>RCSeF
2S=.;8.2AJN),QZQHQ45)F/I^#7Hg1RL1(9Me\_>F,RU^1adHb:Q:f8.\U5]Pa]Z
Qc6>7OK0()/Q<G/fC&WMOY>4fg[N[,gM/4&2Q2EG#8K_1)M4U[0bePS,ZF7#[8NL
VN5.CQQffAb?e/S6539bYAIQ\X#H8)FL93.[Yg\bCE<2>3f[2f1E9KJ5D#M&\=@T
UB\\,gG[Tf4_;[WM)@MOHXXKQTd[6JKUe4O[GPJV+W;8X-)efe)-X0:4KDFI3B=L
aRd.PV<UcY49YY<3\39<_+OYNHE<PfefP1-ba,(I4eC3<DWKb-c=/.)-3)<aG5fA
39UdULJ^_7<W2\#cbEfWMf5Y9/f36g&ZU-:J5AI57UM&NNY2ABb>T.6^EM,_N(8.
/Ia.=L[TV<DAA6,-&P5&M8RI)BMS6?]0<,U>0WH\#F5/#NE<_75,^^g7NX>=2d,/
f.1C?^\YQ\-3U0M_;KDI&PV5@,&^XJ^^e5N8ZIH17\,8+7;d8NFBf]T;+]N&2f^^
Obb+XL:Yg)+b,?c/J6/;CPbc1N@7##GRbaBd8T?>1<J)46RQ\&F2?RKW)[4?O3YL
G1Q#:S#PbCg[V@g.H13aG=c,&J3IgAg#4X5Pa1W6S2=:M[1IN&<_[g0BQb&9?0OV
PcgSUM>6>26;IE;dZAM)]_/LJfHN-F+U#dIPAYHDYP8DVEXLS2,]4JQO.6QPD-CS
)O(YQE_B^CS\H<TK#d(Qd769Z+;-L2/L4[a,DcXbbU26@_TXaQ(QPGD8)66N?2[Y
EVc/@1EFDA9QbRfJf/IW^&,)SdPZL;V\&/e._3]6():T6ZU8;_,ZL<U>gd,-eeYF
<8T.a9R)2X4cWG,e38WL-O&KHM4<TO-1Q;;MFg?6L@WMU:72OY3Y9\C?>6M1AEM(
dg#)GKSG+>V+<c6d,aP:)YVOX;)QYMJdfC=T]:2aN@9/FYX;<_I9/>fbYF:<g-UB
@A&=SVJ^bC:?\++D,QP[OG/@aK+<e+<K=cMOOK<YHU0X\#:]-3]\0=LB_U?@E^L_
-eF3>>eSfB:LOefCTUg0a4-,LT_.0@76AK\gW=/5_7@7O#K;L-1:4g5FM\PHE.ca
Q<3JTCX))a-2DK1;4#SW@[&AK3dd4:F7+eSgeT:=GVI)&C_KH?+B]GGW@URb],R4
;^LWW5cLTAYGWe9_<c(SV+^U#:@.REc&)6?I3FW==G_3(68W8]bacfbU@FDHVIJd
I:9XG>R]VNM1-]/1JD3##,>>-\I94W6<EdXO3)1Wg>d9&7A?-MEH9I/(:Fg3B_?d
DfNKd0aB3g&4a4eePSH]6S_/<;cS\4fC[;5JeCWRCHUW02#B98g]e[>fCdC2Y7dK
LI<e;C,+5TTZKe^_T)gLC[HELF/E:W/9,]4#0TUf5\XD7\EMX,O/fZI0aaCZ_^G.
#f^](6US4b)#RJL61AS.?T:+C9&+:7e@<BYMCY]\.U908<=MDfa]C?b+GY,8)L95
gUe=AQb]AK;3HS3bN0]I9/<TDXD3N=VMKTIfFVb>FRG@&D?;cPA1Z.6:1OC^f8Ve
fX7O7^7b:U?3Q8gEE6\L&M4Y<J>.6e#?(>;2&<NC+D)/MgMR4OM#>/ePg2cDa6CS
Pg?&_5(_\CfUY^34<M\G[RM9=b(_-fBV[16];#gO_AED(5EX6J<J[M:#SACWf.(O
15b9DWZa2@#XC@aEb()4;XTX4HKCE<R&1BegS,/4#Z[0HW6TF9>C@TPXZRT[A1;J
?5.)GX08YX]NU8:1Zg1WY?RXd3g\g=a[^YdUJELD50XRKZ2b>8HDVRB+9UdE[K+c
bP)(QK<NF<4cCcO>Rf+a+f3f?]KHG^T+&QP?9J((T?G=<>/XMIST]KgNRcO:M26?
gC;Z9RI@D,5gI_0U6W?/2g^A31VVH@0eLOeOI1+U=QX8)27(?7Q95DSX45TZ3N;&
WSN#7cQ83a[cP?/J6H,Y;80#FN(EfQ<?>Sg=I70<DDN\2>>cX]X<IK9;5KU.4O.]
X[8DdW#=)<SUVg=K7O(EMD(L9\OT[SX7c=\ERDXIEd_58:ZD:d?QfTgeY_#&A\Gc
K<D55/-6ODMT)54\2QJ[T@QfOAV5:2SYU>OGe58a7#N_CbG[62ZH-Od?AKW&#6c7
9</g5LQ(6IEa,;:JaKLZ>>)&ae)JR2G;:-&12[d2#+IM>57_(8MMaV\AI#6:-TJ2
G1/VOgHG+H3-8WYb>+\(UMcagWO-K=c^[Rf&#K[JCAGAZT7N(XfV<1g6S:&JZ;)B
gOa=?Pc]NT_NOWG:NT?FXQKWN/=-Y&gN1C[72]:5L7Y=dKMcL-XK,:[-B,[ZI@Bf
?ITEV8cb.DH(E.3gU#d/&WfcFZEX\EN?T<cQ362H2:@:77.+J?(^,]MDN<6]>V+/
K,;3:#++g#C&-0XE?M\e;&VGO#VM<(,/C)<5W(Z\C:DgbggVW1^TO/YCHMF/-;KF
c+FG[geFIOe3G0-6MTI\2N,]WcA5P-\,GaN#2b0RK<.gFC:EJ@)CQ)EOZQ;[F+)d
J5a5g./M#f8XRJde[9RBI;+:42&UKNG[O5T.J4[HE(0B/7KWP2/]:aU,@L4e87U:
V7SEfGL2+G-2adCb>&USPO^19:?FIA^U>#dL>9/(]W:C=^^GO+I\B<;0>gbGS-aT
9:9>XZPNffE4AWba8,abH;?/fB@g#W8LGJe6.7=<Y>_&NC\O(K-0LDEXeHYN:JSQ
)9]D&=#TV=IP3S68_aQO]2>\L@XVc7UXR#:=SN5f,a\DCCEabX^=a((GB1/4&6f?
@/8WD;H_e9._\1(1A/M]QG[RU?3#?+50K&Y[GLMW7?1GXSMI4I-Z(;77Mg(M&.^=
::OeA/NWaDGNNZG3JVO4#=1WJC)f+]4UF5RSI?M5^d)7.;#_SVOI<HRD(0+394YB
=KH]<FQN0>,CH;8^LZ^VV8fUC+HbOQO/9Ga65-S-gagf9R2^;G2BTQJ>5WH8TgP2
efWGJAHa@:B]Cf7-<=HbZN?(ZSTMSE_+3H4Y@1eI(I4^UUPYE0V/G,S1He/;c@6Z
];102E=4S&c/-E(HGGPUfb,B430>g&FNFR#21FB5_H@6ZUaeHW>/_5c-K\NE-]WF
YA?1XLI\8M9Y;05X^G3)Pc\-UYLfKggJ-,AfaY>B/W40M_BWMXEAYKaR<X;e1LXS
3U&A&HF2SFPd1WNS3VBVBPN2M^36GNW#a0@M-O<T=0=Ze-M-7T/@(/RVb.ZR7E@1
4QTG?9&(A.+[K+FX^d7.OP6T]_>8;g7C1gY+V;Fb>S)[-)>Q41=?=S54<bgd/\4-
N1IR-NE1BeVMZA@5@K=:[ASO24.F&H?edE]BRE</=UBad?0;:PXYU>^#gFMIIBHR
Kf).+>NDSEd#PfG\MWSacb;dLU,Y-)Ud1a-VX4:db)FQcCMAPK7-,J2W]>e>6,V,
eJX=3QC^9c9B2JaLJ#&1MPNcLb>df;JO[C.b@fXSTDfEZS4I]O[T#8WKNK+NQG5a
NO&dUQYDFcb&aIN1_<H]_EN=E2c#UZ>8[+e_CAY)2I8_Q4)48^W]-.]ZAMG_2Uc;
4>eWH;SV)+M#,Xf/I&=LDCe48cK3^:6?Z92PK5?bf#2HIW]CDMVRH^DN-e\V@J@I
N8aPOB_7^6IQP;YTf@H#dbTR17D5IK]gJ76;&TU1^B#&Q&&U_-_NFE+-Y1HQg#P[
PRA;.e&6c(QBbJ<_>F?-[?\1/a2)Z>5AgSXM2\/ON7RI4W90^WFP5)(6C7\e<\&Q
g4LYHL-[Ie->MZR&D;A@5/@_XWf\J4X#8MDV^VN^98c\7OT57LE(^M+(1f<[BZ:Y
f_R)6YUGY.H20[+OC_>RBc;:,(4J_8?X1NP)V<((Y(SL.LfNL@&L-f:,,Y1TOGVL
,KfBR>TO/]#^O\R^1D;MT.6+4L@H>R&LG+V1UI9DDUL,;aG\DTc4N(FI.[?dS<-B
,WP&XZ9-2(K_JW(-^L;D:a>\7:KdS:=Sf7a&YAI^OgS]8;eMO77ZA><JO0aL8T[/
B4&VX3&U4,Y-B=AE=\+\G9.NG4FWC1T5#\#UO(QUd3M1POE5<?fHU;b+R6+4M-GU
7W;WXYIRfSBR]Aa6X4[8-<JS4+KTWHLLY4c1[@GKaMd7O#:7#Ha8bUdO&\Z<-Re\
-&<M/(FI[VI&DBM27[;AWc))4S:d92WK=HLF,#1)0BF323]HK@D6P?JNH@.:(-da
UT+TVgY=Q:4P>6&A42OaHJRe+d5BYVLH)1#;[Ae0_Ge::g]6c&?8[(]CO,4[/Z8)
RZB(1F-3)&:N5QIMT^7KILOT]RbKYb\&^S3V_^1+#SGadI0)EK>d<HPI=fB2F^VT
[6cf2,FW;cV;a]]\@EZX.a4Q0HE&?\07&<+I.@0bN25;eFX?deNI>K,ICH74Nf)Z
.3LgJa]L;4A<a7-(f>7OB?Ia[(29YO0(/eKK52cZZ?D3^UY6/8+5FKfC.TJ2?9<[
PW?_[eN/6Tc7cG(?3BLU&-R]MKG(WVAPAd6>ZTa;D=5LB\d6LG[d9#QFIZ\(<G0e
W>OO.H48)X/ZJS,P6G_>78/:M-J[Z7HKYb.fXLB2S\)FVLYDG1(4<X:adHZ=H9Q[
YOc?VTE[9W//8B,/FT2?>SSK8\,=>W+S_1IGO@e#(GYJE^c3_O340b>M/58a3CG@
Ug,ZFBBB[0#&8.53/(-\)E-ARMWUAWU;;LMaJQJ0\9fdU88FSa[<;H]]d90WF+W1
fQIF4Y>3@<ea#L)PKVWcIN#.1Sa&?CVg9Y)ad4PS^5&B6)[&C?(+:H9Le>Y@1K]b
TW#bK9ZO>:;Z+fJRTY.1#0dVa2[<gO<MfQ64TR_O4X6=g2&Kg,d^-QHX@\>AO&7H
RDgb\K<.?Y1FX_JY0#LS7OG6]-4/SHYL?+.Tb\We1;0XR<bc9]JIJK#VC\C-)O=T
aKg(geY)Y-]LgHAZ^08LQ#1ACK&)Q+OJ(cNUH#,_FSSKaPSDd[d6-C&@:?ZZ(Qc:
O_HTQ:bL<G\P^aB.:B#I)11)b<>.-X:86R;0A?@_N&#AQBJ=3T3XPV+&[-#@D_F)
^-618]#91@&X@G2LS3;H)CIWB3CIY<+C1(D8_D@X0DWS36U9&Ib@L\Q\9E-b3aLf
VSGFG//g&&/&>LHa7[YQQS\>&WR,S?9gbebe3V<)E4/S=@NacUQ?5HII2a33P#O>
XT8WO=4+K6.>1\a3<#2#7W/04SH5#g:[<BTXdL0^24=WKZda_<65JO8-)\?b1Q,^
.]IRQ+/KW3(S_,&G]<?+^0fOc;AZO:Z=WLfcTcZNbA=>Qf>NYLf,b[E]WSNQHF]I
8SD:&CTJa=&LGC/?+\-aPA^QNMXHH(6P5/ae<Y5@A5DP\)H6YLf4Z8BW7=#Ogca/
JCC<:=D_Y&48PV4C/K</+L@&eQA<e?,&1gaU<OWeVeXYA6]b_dRR9,Q=HEOf#WW6
SDF<P)46(If5bZeCJgLTTOaOcB,f?4X1=XL3<YDXG8PUgF,(30BO^15)fNU^#g6X
;P@Yd\M,R[?Y>QX1C^X/C1TFZ#:1<9^5M-+IQYJ:RM6-:<GPTKT,2+X,<K@NP_E8
F>Xb9GG?EfA9SV-9Na@f<L6AZ\-2CeP?_O,c@cPTGac@CM(31JQ>02I<QC6I&A_d
;/QOU)1E^?/J+=?@cE@2GXPU5N9dbV9(H?^3_CJ:_+WGdIF#+B&P]ML]2EO^0Q)4
.FgK,0OIc9?VP3@AUPW02/E\T)4W_T=@1XE_=d^_3W2IFK(Y--)VRU/F33;6GYT]
K6,-#LefXLVDI;4]BR(Sc>#Hc]N&S:Q5g=ET8ZSQ/VA,6J1[R41)SMf-P9146.,A
/7/cca><cYKQ7dKe(M._O(B+/QP=][6QOd<&\V(MPCQ=e1;2CQ>ODS6Y=>;?<4-1
^aL:fIA_UNd#=>Of,Ce8U#-@?_NH##&DO\_F907SM(#eHVXDG1O1@J#69UaEFd&F
8@aW)REP_(aO6cK/Ob//QW8[OKdc<DbTL)KY+fbQ6CLg,C(\L#4ZQ.g3K:@f>g@Z
GIKe>21AU(#1UW4ZT+7^AfK,JPOK]R)FP4U9,V>XSd_cM[4H_/]@2P@D(V=gU);&
9C_G7SBUTM6NNP2]S07G1ELa)Z5Q(J@J,I4g]6:)B\PN3S7ZSd7:;O[0I[J?<#)D
NT+0=4;C(g)-G6>VDHTO2\^S,1CYOM85[@]Da]LJ.e+0K)KJ:g((Ab#C7\XIbE&^
:aF?ZS-[HB^B_UDHFa^JVDWK=>M>eaNW#CX48_UZ8VRW_AfBb@-W7]2D\)M6:U+<
C(.(;Z&JW[78-F)5;U6A:fHM&0F,(LTLfZ,M,7?R]TaV>6;G;dBI1RF7Rg-,MZ3(
E_ZLCG/F<V=](WZJF&gfP(,IfcVAEgYeEE)>O+J=A34>,eLHQ7I90J4QRQbIR2J4
EY89R+Y2^A+d[a^IcSHX0\G12+;L:E3A?N\abZf?a.^3fD<Bb?Y^^\Y5)eC.Z@dM
O(+-:,B_d\2X@G.OGFM3F=C:4Z]SV^gR7G&+/C7OE]bd;.?;-?R]=YbW1P&3J=.2
R;2[BZNQK9=S]&Be2I-QZCOHbCcU@d@1RZM?D5+OT?LG/HJ)CG]>KT/-C>O5/a5Y
S3E33_1d[c:8;#a&R,[\a;\D#>_Q5@fAQfAd0OFf?#V/F=[V2L(1IFWS303&+[4Q
Bg?AO)VE@&M?UP0_e\_VQW3K/WG_RYJ;[NWCUM)^\a=<1</:fVeS#E#eG5F-R,70
?Zb7:=b\,PGR]WeZC9&4+25Oa,X3.?<Vd0E2PU=KN4N^&+BPS]PO^4GML0\0ZU49
e6M[/ebb/9+cI>H=WT0^7BfMS)08P;-)Z>MRZ^2fRc]EJ\c@^c3b=;1979f:P\?c
8-G.WZ:>9IDfcg=57]QA_<7&>O^Y)]<9D6WM:Q12eP>^IYNgKebP0>GW2)&G>^[=
2(-R>fd.F\Z.:9KXHg\W0B6E2LF,CV_Pf)8\IU6gF++8+bU9D]f[Y<e\[d35-4.a
K+<,fQ]WD5=?/gT(#R([Y^)5]@#:\2P/SYC?=UR+]2Fa)P>[;ge7##F-FQIbgOAH
YKgU[a-CP@8dG;Ef3F_+M.B:-UE]WNSb:EX?Q9DLa+N3OL>,O#:2Wg<]f(5_UGOH
G_H1BB9?4bQg+:6.E5AYGf_(62PBaaX?>4(DR\aKY+[#3AL:6)U_FWf:T5_BKOU5
8T_J>+8X7d0)36S8AW2R51BW:3FC5UW,;>(8D;&:TPbS6HAP@P<9BMLK)^[&P3da
:^(9@=7@e#d_\91?OE?]b8US\2F4cX:Zb@<b8Y0FWN@gI5CKQ^^44IBb2)cZZIHC
/<IEcaF6]3bRXOX==Pc@OHA=HdX2Y6#;QS(V(&c9\[7G)Ca0=:8:=cd#7Y5c<6F&
ZYb8T1^Vc[W.<R0Yf&2>7X<L?DWY.ad5ZAL4bTdX;UAX]E=]H,d/fWT\-cE8Ta.R
-.C<gTfX0QgB?JFS,R\b:CaB<0#dAN75>6b]6_\J)J[TY(JO1[d>X@_K>Jabe^LS
^D8^LK&EA0Q-60RLG41:b-(AeY2Sa&2K.09e@-#72SR7UO>6e10S;-c2)B(VZ&C2
][;Y=W]NJ?,::FCUGR4)P3BE-I#HYFc5[]A,a1/(4H6#3OIT3#<TN(VPND@-0\@X
(1_Hf:56S_P&SM(7Y:KS@IH5Ba.06Xe_;KI&Q4=9e2[QECNL&8b2JN.f@>UI\c\e
MJR0UO(UB.c0g<]2ZBS&RJeDSJQ0G8<&+GO\W5WBRF>1+-O7#-D1Rf6J0=45M[fN
,?G>]0ZAV_W-V&ac#beXUU+7@JE//JO?>0@0]>E)1QLZD9T34@O</D3@)\XGYOIf
C:G:DOXP>M-_@6+O3b=6YOcDcNV4XbE^Z]Ag2B<P,FDXPA>+-I4J]S=:MD0Q3:BU
Q(QgB1b+4c08QQTBb^6Y9PP:QdTYcLfaCAY)X3f\A.MJb,J]bLY)N1ZN=[S59H#R
:WUB[=U3B17J]PL.d@:fZ9.:CVDY37UcV1I])0g;H5..@?^cNGa#P5.(BX)_B^QK
R53W;=/]:GBAD6\KR;C>-b<#89-+GS[8W9HH4BA[\Z&BFMC.BE-D=)5-XFJ#3Pc(
:<]1OZRD_T:1GdQ,S,&Ia#5)9R#3#\^TCAZXB7)A/e4(ad.1=EfL.M=WL)YH5aAT
LE(NC#DAeF:.ME@;+dB7@;GG]<59C9b&[D<,06-,U+/K<GH&?=9)LH4&MB_,1BB?
+4)._CUYfIdOU]@#K.@>?+<#HgJe_>LF>eCZ=NUAL21[T_+=S2?O\0ef?_904Dd[
ZB&/JaXUX95ePQZ&6d,[X0XMR?bEVLCDK&UA<7SXC__J;[;B?,Ta(BJ@[N+#Z2G7
@A,=CH\_.(G2:]OP-;:.G^L6fd,<Sa-QB8F3<B3;gEM,WeTX25;<0/L:15cL6#S&
XXQE3#0_A@TV-WdG_e_=TcOfNTd=A<X>=I@HW3KSB[0MDDDZdFJ)<ZC]8TR^_>LU
=eZ7^>VQ&Ob_A)(cPNF3(M06EMS3/U\O:ENNMd5C#7&BI&dgf9V?=DJTXN8X9KKK
NM8KVZP1)FXSQVf>I01IQ-K#Hc,T@6BUS(D[A&<G@FMG<N^3QGOLXGT;6X3@92RN
e&LZNVYWWK5f[42<C;d-DJ,.JOacK^HLH]CQT?SI;=X#C[1XORB8La)12A.EZeC7
Mde6AS61BZcG(A_T91d\+@e3S_Q3PQ^7M/fMWZ2-be[O9<aXE<g_2LS?,fTT<d#Q
aOUA73DZN,BNf#F)=UM/>>BHc&C;+V4WV8BeW&OE-NT:CW#9PQe,82@g]B/7XPbQ
X;S@L#d8aG<64Ne3eX2ab/ZN^B(4fS)4?c>1)HNB)4Y^:X7XYY6S@f[76d_60>)g
H,<Q7,,-B8S3&=5CUQO.&6BYHCdd\R;/GdR?A_AH+]ca1>R6>\+I(Cfe^cWZ@&.<
E=L<F9JGT7&K.IRFORB3H/88<=KT:;N&cTWI5K>Z<O-P[fNIAD-0fP+Z?GMQ4Q&e
Q1A5-@aP,)QfH@213#A/c[^YHVY2QXe)27_E_@&9J0MfA3YYN0Q:GWD+9#IAZf#:
f,J8c1:CaU=7AORN3X&AI>FK)A5#H=(YQ=)#/I1;8MFcGSP3?,OXUL4X4@JNK2;_
>BAA+:79Pb87-:\]6:Yf@g5?L(_I,b@CIE:<+9+J\UZ<O755BAb6<d_[ZH[CX@b]
b1X9E@fE&g^1]P_9><^)cSFH_^2.e:8(<.L<+EE^89G+PBKM,>XTCP)&d/CEE+G2
RQ];9:#O+Y8V[f@.RWZ_?,K2_TEfe;Ud/S_1[3gg#U#TbdQ]K<KAT?>=0_UBCC>B
c\WJYYOg8V/VFRB(:O)4<C28P7(#\IK;_\3R_^JHI5d9(\=E0F2>8_42(X.A=d(Q
&(M:DQ&dRE\>3P(R-/dbFC=#R,5,Bce[X7g#:W@<FT(JD8USA6b]67f\XMD_XKKD
D;:Z&/V=[?LEY/3=1[PA7B=&fW:T0#11?CdcW9bKcJ<b4;9a<XGZW&LLY8WZ)+]^
(7SIKeg66c0_7,7TSOPKabC1S7;]Q4EZC^@XQ;\c5[a/;0]VH.d[3:7W?6_<bF[J
I7AM_ebP2(_=&=N99?0,-R>>@,TY_0RE(;EQ.Z_;;YVO?WXS[4(;@de3\L24Fg)[
S](e+84-gZXS_T;TF@I@?&?]BSDFBDCI&+QQMG(UMTZC1HLE1(](EeDa#0S8aQMU
/CY6^FC0@4F(PP[4S^0F1Te+@N5//?;H5e^=JB.[;/P]6VPHRE]RY9)<9R1N/(ML
Vdf()=.LH_+@UO0a@c<a2D1KL-CLeQSSAA;2>A(E_-YZRGH1;Dd,T2U]()<a9c9A
J&KBT[\:4-N@b:(/WZXO(V]Zg;LgAW/0MY-[HVe9^JB@&CAWeaA(^E1-,T2):XMK
=@)?Haa(@=U&^Yd:..>D0Cb__VI@)D6Y94+AZc\7;G@=\8;)aI=Wg<1&bAQ;(/>_
3=KJcf?C//_IG<8UP]>OO(Q,@M0e8_>8&]-PAVD4#[aN./AKYS42f5<a8>LGAL,&
G</KHOIXE-:F4JSTb10^^W6c8_.,&<a>#IXG1G_fW,AYK-3B3,7:FG+))WV3c1T.
G&O[]Te-+QSU_8CcY7PZCBC[B^+ERU9NVR]Mf42/(_+3K]3e^-G5BYZKS^cL+,;Q
>L69H@F)W+V[C&H/<(AYBa_,-F=E\PS<G_J&P=YWN-EE.NfgaS0\LF(B<).c2K,H
1SB,e[fSbX05T1d=60[5OA;-K((6D/_/BDgQ_D^.>6dH8_b)BELEJ[e2CES:H9Q1
8@VM;.-/Z,MP@4^cDLAJa+<UQ;Qd/WAJOQ^[(7II+)T?O+&NZ0G#-@@99)QL4b#B
f@0Q/<#[SK7=GLW//NSK<e7-C-gF]0Me3A+TBfE=[9U;FP(R._KGSL3OOL#H#1=.
e^#?.(DHaLHAg]LP_:#)HZSS]V+/--N2[AOX.T-&2_aK#M]-CdI?92>f^8<@1M1]
)>e)VbbA_0\;H;-5Q&.ZLIXHE,48HS-,7([9]VJ7cNRMN[)4KRQaBE;9=gG6gW2K
5;:W7X/#8FYIX@P?ge9)FA#0\CR/(<XKM,FG^?01AW2&^NI;[&;g7a.=fW>&3C>[
]]PM[0D\O4#;LUAX/<1YN8I,D\,cM-Z&+aU,GaIRb@D)_28\6R>-:g:#D3,]PbAZ
>-;OJCDf#S9Y<3SaTAgUP.^W9(ENIb3YXdF^g=Hf_1F[(\9<85Eg??GR]QS&WQ8[
<>g@d^O1WV7^/cH01Od?#6/T-U,b62d;1:/YS>2U;Y^&ESO5KI>5#bHf7gV=#,eg
:-e=.]OJ,5gU]VTacMOOD=>7b12bNG2IK/K,2#b5LH87fR-0Z2ODQ8]HXaK<NI[N
[O_?;3<JSCMWDE9?/8Y?VS?,&aQgf?Q;#J],LIaB+)CZG[2#1VGLNX#O:+BXLPE6
+:T0@_(bgIgQ_1N>\N.(YNgKHGCb[IgA7YR;,>M?\.>VTR4SR+D@XX.L7&<<6^5W
<;N:D1A&<_Ma[B])1==)@VO_T5ZYM^fH-=cO/;L.HFK(7=-QZ8?cIO@4eF8XHCPd
XVaP,.#<S8)P-5da1.J5T&^/PX@6Y8RKVJ7aK4YM&9&:cW(Y&Rg9R:MA3@?PU_+a
R.2Od_(YTXB,T72.b@7dOcFYb&?-B5Ub;[OWNbe6[gHW^3L<Y3g\bXKgXGZQRD-0
#P.CfO=XR]dKOK9_3NNe6ZYCa8bZQb9H)X)\G@/&Z)Kb8J/c=N-CU@[R9K:VC>LD
Y@,=MU-:V1NTbAY<YDMP^3T=YS.L^Z(aE9a&-gM14Y;_d8W011QX#cR1ZgZYb_3f
)_42KW_B/]IF\DYKE(-H&?0QC?#D(FU/4/+ZJ>fFIfYLPX]]/Y.J^Y?C,I<JE-<I
>Nc]69eC&dLAXbW\4J8OBF0&QdH>PX,B?L93B9B5N2f?(2U+T?F<C83,#;0[^JL^
0.N[OgQS3^T7\U5(A6?J>7,8UBVV;1W^HA15aQ-L@R;?1Q@(YHRdO;;P>MH>37H>
b@+>dJa<,,2S-[Zgd_LV6g8@0(BG@R#I5N>;^e-?aIX3OdLYf#;-HN@59Dg.BX04
2/BCGPaB,D.O@/E\FgWDP[>Z]-g7dN-VMA4JJYfPc0c^a.M(FNTB+80a.:@7>\3I
K[AN^Q(5=0d]I<G.7.;26_7K3W9GT#CLMf28aA[VIfc+;ZC55AQM(c0Fcb4#=PU/
eAN=fKbH?F?;fT[Y<E65ZGQYI69:/X#2PLZHD3eb+9.WH&c?TNYCa117IB>4_3E4
R)ff(_ObU9TOa9?O<c6ZJI:UB@A6FB+,?)D:+.23P>=gZT@?XG)G2;-NQC8@A0Gg
MV^N-(84R-FaYK@^bE3G_LF<dc7K(c,//;AL\<<c8KbEH,O[[Q9.__W12SC_9:DC
WMUVOJc07M9@G(5L;?OQ@7;:J;Y,V]#M+?D=2/L0649e[Y=;U[CL.D1Q8cXU>BZ;
,)C/07/_-__U^4J/N,6XcI^)2++-UcZb6GU#A)[_02f3MOHaca[?]cB97G+/^Ue_
?3CgO5HScF\3Y]>)0UK>OQ5Xb?T=1,PB)I[QMOA^:V.?KaM]M_EeAHH@b3WL@7cV
BBE.Y9aF6<5C[Y0D[XG#6_g8(a9<RBgO?6Q0&+c8ZV4bFTAI>(b-a/edC@K4J-?0
Kf[G#GbTf6Nf^BUDVeJ6]e^d.]X2I)eC,BM_UIWW5Q^>BSbbf[/?DdP1,=2XF>.J
9JVN+]+N4/Gd#(&(WeAT4U.F=2\)KcZDBf&T=<8-BQCNFMHD_GN4#+GM(_2UDdRR
gd,)_^2&?ZQM/c=J,^?.SR9;2BA3+[R(gJMORX=LI:cU-(YAN\:<7EfLRC3/@4^8
+4XZ)I]4>+_Af0>(>LD]A<fb,;N@0=]SaTO^.f5C3]5_7]:R_f;BPfaNTLV]^_6\
O_eXGU_fa/d&<H/a7MJ;1>DNL\ba]ONUG_\_J,NfKRUYKNM>Q8T+P1_4KeUHQLUS
[GS>P<VWNA,J<gT61>OT_E,I27S8dC:LKWM-APPN7Fa6ZbX]=A(@fDR1c5[?M=8a
HL8=]+K\WM/^dPa^H4fF@7Mc451[)L.0c<CWLFC__X0a87S,,Dd3RAPe_L?._BA)
eC8gHN8?U:>Ig,/ERGJ/P4F&Z2HGDL];\].SUW5IKb9R.6fP_:1EfcS6DdPCbHW-
/,+f/#PN5aa5)d3c-B0gE<XO\6/09b-5DS)>@PS_d<D#-FCJ?QdUTRSPL?XYB32.
N;U=2J6MI:1FV04H[?M-FW8JV8^#X55+U539@<-(0)Da__d_V,JgYC@;:4A=+XYO
EXR&<K<75a^4FNXeSdGEB,cB4@HbX=QLa45;8[\b#JP4:[XE>TW?XD=B29H][YUP
?2JN\ZA9SO4PGKY.@_b-5Q5,f_gXAG-Y4UF(?<N)6e3Y4#U0cQD#4X#H99GD_FF9
I73dO41d(/Dca(Z+(0\d>5^BH><^52\_c&72Z6)1CFf9D-I6L[7D/dY5VY)d+R&g
M.fPO(b?3FTA9G2b&]V#4/6R@NVeUL^/:8_K;d-6SPeXO?GV?HO#;&[^:2XS;[7;
ZM_EKb5F9\Sc&9f4dLCB1L7(f5&-?-4La\Aa<77@097VPQ1+A)JSC1YRHI)X8?)P
#Zg]XWVaCCFH?JJ(-E[Kbg.KcB;\YKM,VdQ=15.JdF/E)YU1>>a]IPd6-^UA1@<&
WN]90Q2Nc\X9GVRaebXV#f1HaZf=d]R30D2IL#)2A]6/=A2@ZQXOTM3ZfNIdf_N6
c)]A4>>N5VC3X<[JQS;?#-8(b\5KB?PHBX?CQV.-AIK/<d0Y]CRQJ/6-8[K\;Yd:
R98)U+AKLce_WQG1HdD7dd,X=<QT/gH4AbH09bZJ5Bf2G6FMXSIT47+NgLb\=ODF
\;@)QfAYg_ZP4:f6QUg9NbW<bgIggW&a)Fb/[V0XKUB&&#fNDBbdCaSDeYQV0d4F
^JX#5D[0&(UF<3/SJ5(dS5@:_/a?M-MD3EKB:BTYZ(T[+:_[_G&&CA)6\_MPe7e?
ZI[C.SV5XcCc++A4?>NNN):.U)A,13P=/f3^3T[28f+@5[K4Ac>[c-0-_SX7EbEK
]=?N6_8O5+W]KUf[V._^WT32/(a(XT;YMfNIKIN>PDP4\7=CSGA2bGG#9MY^KV>8
M/RV:[^A-EEX8c4YCfX3-QcLGWFW5;HPQ_/&a>IF<I(P:P(AAZ1ZW#Q4KS#.ABRN
AcH+,V+1EESUB<dFSaf\9_I&BU?1c_c?C4-C/A4_QXDg2ROOMV9SF+DM)VP8-JAC
YW@@C^HL-:eMT<1M0]GYMDbM162I)FPG+BbcT#J,YdAa&BWfg&aTBL8RZ6AM_/:d
CE,Pf96\3VD\aCZ/UaMWTRLKXK_,6&^1b<5W@(\_H1H<Q7Q2R(0#+BG6e^GK6NJc
a3#\C#1/.]/UOHT&WYGPK]d;70C)H=)-:K4gLY-dDY7KX6(aVL0CK:bII&?/JO..
)20FCS#gVI_:V^f^8)gWD/Q(TH5M<RSCeU^J#,)L.d&eY/?F_FIPMXS>5,Fcd(Y+
ZL&X+PdK<NbJ38/f_>A\g.B(>KdSPNdd@3[)2UL3Y#;Ce#_1BR9X]7COHZ?\_g7]
CR&OM#?>+<_:GKdYadc19R1#9cW56VH8bZ]9\7XM0F;Lb.\;bIEKUJ>;UXG[OL[e
J?9I-_MA./QN.(aHLIT6#+U?])HR.aMGH]\7:L^Xbe8#4ZNbVE>S5/RPDUXAABVb
(+X/]]H<IGL[1Ld?#f:U3/f]K,YE>MaD+dIO[gG-X3dR2XM^b8WLBJ:JD-D78I-a
XLdLJP+RdTM/E?G=#_)DWG:Wd.-#aQDD_W)[fUKSNR;fBHI^TP0^3S:<g4af92&(
^Mag/(?9=SS([Y)AXf0C.+\dcaI_3-g)[&YdfLcZN)g01J7_IAFWC5c3:C#L2G)-
YKDS=(-[3Z,EL12&X7YeJFfPF2W^6LbP4T#MG+,=O5\1,])]g5c\&L9J]Z4VU&YQ
5BdGCQ]E+D3N#_cH\egB_./@:0TOe6Ma#5c#V7cI8\?YCU11VWPSa&N_6@KXA3I\
BL9HH]40IX49J]Y65L]\Zc23<X)[daE]dS280A8SYSS0#\R?A(LS/fTPNG&d\ZBN
TWGg:T_L(.-<+Vf@W&W:CeM3)a]6K7#=M10]E&b,0N]F;bJV^3)XX\1S70E=J#=X
=CQV6?JOMgLK8PbPS)LMTGgJ\?aPB;G46EY2Q;AfN]NB38N>Y/Ic]X2g4X1_J&2G
7J=6-=Y@2.09(@&K7[f&Z0IbbMda@?O=R.C8].Lf&&\6EP3<(\<A+f6)>(HVg0Gc
0+(CWdCXX^>dLd[HR=&BFYNE&<CQR=B(f13.-eP3]W?S,Z1D^YLVSbdHGg7LbCA1
,T_93ZYVI2c&E>)XE[9D2C]eC+E.F:XHM[T>5C30[L2=2+:?dM3aEeW/?M6WH;Fa
FbB9AH[2W=Mb5TWWDETP50ECHE])SJA>Q140g0FbACF-AMFd9AC^4=70QeQ8?J^X
]:,QK&)V,1U8a:6NaRXVBCZ_&gT[AWFQ./RVCa:IGB4Y3b]Z=K;,.SM1H:D,d+(\
?K&b^FESH1T>](;1LR3V;-/P3+5BDP@B]3dgM._gH=Q-#;-8;HN?XfH70Kf4SM&=
+.]7U3NAS;HL4P:Q=6DYe03HVG&GC2EOgMaQb:2AbX]8Nb\T6,IK@ZV\gZcMFVdW
fV@]>VA^LD]dKD>9/+/8fNcP@KQYP<&X@ZSDJL/E_P1#.;^:-O\gdK\a;.3N0(8G
(g?S7+K03T@+TCOC@&cNTENR(@R>1@V?>_\(Q-6>:OD92?baYRBS[;gL;G;g1f/2
C:O97P7/]9FdLdTa??[;Ye^RO<0\f-@>7aF/X<Z-OD8\aX)gT.9RS#&:^(6LU:Xe
)9Y2NZC#)U@=NGWg5GR\T,;BTOP,A2C;[SL6A@W=SG?3,V[G3/f3#8=[>RU/(eJg
Gfg<b;YA^O]NG[g27.:^N6Nc92IPNgS,NL(C0a)MZD/[O4EX?fUV<=DA9c-6U:;3
I?85d9ZW+4Y[JK+D.R#.dINY)UNa<FZ,LN;1Df2_GY&Nd(7d0fKGCO(WAESOg@0a
e6VM@bWOCNQ9dbZZ_2A<^1WLag::(DA,g/B.Y:_?@L789:>#+-d=#&)NbH+@=d<P
X\E5=@c:.VDCA27KU(E94(:CC.[4(6<RH^S:LB=0Oa1F:^C.&CA,^-a:;H[<WbBV
a44D@8L-YL>+6Q?+_DDIQ.@NF6F[@L67gYJM,[WX-NI8AL\U)b&\[F(]>?-(S?_0
=Jc4DLccE\eX(X2aX_O2NaC31ELePB,.;[E#A0^H(?NF[./BDW2>Z[EN19I7TGPb
N+Pd<I1+9TSM?V9#ZHY]dG[6UMZP.8O/G28(.Ye8+SX:7cO<_cW@d3RQd>=T,<]2
6<9)eeIN&35>c3NN]+_J\:@INP^9CSTB.Ma(3-#4aE+F+3L-?0=,)C&9FQ1KE1UZ
e^.N9ZYee(&52BLA-8d<?2J(XabZ;,\,W>OVGg6g&B62&IVBB9^6bA_ZO@UXE6f&
R>26&T-8Z4CXTKSKU/X28/1._S.YdQ>0eI,KMVQ?f9@W#GgV]\R,I5I76dS>ea)H
[BR3B:;UH9ed&[\L@2+DFXb\bZNLdcL9PR8=e#@8+IJc&+?RFXV.63HYd5XPQ+_(
V^G4X+Oc(gY8cLY&HVLE548YQ<>T9ZHR?;eaM=eBGNc.b1a>,EFd/#B_&Q:JAA[\
Z-?AB)1K]YO-/[DMVd#fO]8+<f5DQdBN2J32g;S9&35BX4)dX&:<ZXJSYY49YD(V
@JW;EQJ1,/Q6944<:\DS(TEa@,c,9,_QKM&]N98_ag4PG,JS=+W>@GLd4D<5&YXP
,@;D4EC8EEU0f2ZL2787N9F6JCBN)8_Y(a(_&1cW[[B?^\5,US=8[IF]=6O/&#SH
eTTF\U;&(3f:I9]ZX-H8KL&I+d9\?&K[R3gAd\6&L&U;D-0cQ+<@-)?9Bg5#O6Tb
8Kg?/_EW&9OeV)X.0/7OD#S4?M4FdMK613]bFg&9GEZ=L<C@T-TO;[SHI@S8L5KQ
Q=Q<W.^DRC\WJD,)<KcK-=YG97gP_8/bDCVZ@NgWVL7;f#IRD;dK.BX4;I<MDM]_
#4,(3F1[P&IYEAd>Sf0H:/@&I<@TYCW_FcGd)(\@^Z2AKC5SGI-a]R56B]9P^ZW:
X8&cR<=60#=XHgECLBV]F]?MOXb0MD]DZNeg7@[XHBVTfT(<:+b<]:LE596=+EA6
aB1gTA/(;+/TE&B^AAIARGX,UJb(95K(,O5)cB3M3SSdIMXe-JYX;Y+9<.DEFeM?
0U)-NMZTT(7WEA=./-B8A6QQM<]<8.#=[_&1/DQR+#4DZbJL;EI-4ea[[.X#8[b&
?6X]F8cI_6](eBfRBL(@#Q\9_.<:D[=H200OSVeR7+U.J?)@#@-3&&2-8P2W,;K0
S=-_P:OWKPJSBP[BJP2>8)97cN9PG\PO0a24[M+\J=^X_)1f#@L=@KRK,00WYEO)
>#0K6CfL8Wc)#[N91G+?::dSS+f1<:]/D9aXb=_4b9#7d&QR/Ac9fG?]QJNf=H;K
P3<8BF(U::/X9b-@VA.ff2K,/C0DK)=B\2ePG\;>8#?))JI.=@XfKAd+e-W2(&G\
^SGYSQ[P+O0Ng<G+AD+BD1IKBNgE2?&b<=/N8KFZ&#d#-dSeFaXWAY6Ig;+P&F6Z
SJMX/&aH&7\d;6@J(@:].Id15d5N@07N_:L>GX\L#X5^0B@@<25D0)RR(&N^:[(A
.W>\<d9I^WeH@f+012LJIFQF48-#:S+-[:52+PE(cDH>A,aG8D\B#IVcTBJg\gH1
PJ,<)d,..9C.>]2c6@1EG09F;^).9[9G:30FTM6,bV93OR?NLC:K&##VC:C0a<Q,
Kg=42cK=I;=FM.f><a/W5#C,@e/@IDcJH\_=#:4g-,4S>Re[2;bL@5T;[&gCW:EW
NM:RSDaK\O9E;2.W@88.DCd:4b)+RNYC7JKKION^XV4CUURO-\4#-1.WU#ECH[RC
Q(M\3_3CT/e3O)b-M1AIXH@]TPA?H29M0<a8JV,:Cf^MTRG6C)QdV3.>S9df?a]O
_04bgG.,2HJVeVAE;UGA-D.LS\#WUQdALKPQ:OcJGd\\?:</&8L#3CO&MEVJe97A
\L3E=440];TeOO]00I&S;MVTI)gP?;+D<MY]>RM/3c=C58YU4GJT4L<,1F?/]GYd
1<7Fb?J5eVN6UJ:J5J]T]YN02#aS0gH#Y#/4:BVOXIQe>,_E9b?TE1L.>W_/7dA7
R&338SedeG=M@W,P:dTYOMNd/F)I=B@(DB>;;MF?P<T[HNJ)V@6dGT@&(>J]CK57
F.E;&H];:L(44R87AY9_0;Y9YX0KK-9_-VKYcJXFJXLJ1&P0HGLW@GCPQ=F^S4M/
.9.DOe7;]IWUKH?GCR#IA=KE0SF5J3])EgS;:\;d\2KO>;6]G#Sb/?W>-0=dN?/(
d0#PXeT9A@XAM\CI?N,[B]X5F4U_X#>bLNDV::&9P^>57O1/-OaH@FWL,N4NbP>]
ePVX-B/R7J&XGgRNPB92QJZ?b6dOMJD<_F?4QJSN86Bef7WB#gcI@>B&4;];<EEI
MfPUKJ274a718U^_caPBbYe_:75=/>eg-XJ^T9ZNJCA=<dB[\5daL\8J,ZY^/6U.
]01)1[IMAPHbL5bJd=\UXAd&5>a5_@;@R.8fKd>\XORC\Ka+5YY^Y011D.CMG0AU
1?\FT_.2Xf#9)DEBKd>^4GCLc/Y[\&DZ=a)cUK-]WN4&S?_AIda0&IVf7C9+Q-bM
L8;N[0WV6&ITIRf>XQ0PU]W@O1DME3\Z]9:cb5B&O&J][b]M^PH[9(86=WHW7C(2
Ma6@=P9UPNJ7H4a-#@2Q;[6R/1Y3b\3-:g8DH@&aHL==G.&G\XQ#8]>W/P8]^PK;
^a):VI#\)KL8UN>0@23REKH2_@)Z9MC\.QFa3>9+OWU8/[-@1MJ),]2JMO0.b-)9
Y^DF)?_\(ANIO3:1-?8ZgcX>b/_gQ6M30DGbf3We^9?+Dad[0F[&-\YP]Y9(,J9L
Td,3-c<PK>KXG8Y>KeRTYM.(Od)SeV_GUN8JeVLF@&)KAR@aI/)ZBcR]E7CVJQO]
6>M34IQca:3SNbVJI@1:VW7T<L\R=9:Y<1H:Gc[,EQ;a1,AG/X2.G\E:e1TYI0,:
U5P.AS8DAQL@6]J#&+\AZ5V)5,RdKP8]P]2Gg^5/X1X;7D84@920_I4R.K./)34V
FC4c+VH<3Q^3?cG,GfOb=JV)23L,KH9>Ka[C@81H\Q\M5ANPN?e4DAc55[KQR>ZG
a5SEB:C12G>(59Q@gg]OWW#R5fMaCR-EOV,dJ@_Y+U1RYPEd&_34K:e_O/0-?\9e
\+BN.O7>C+_Df(8;Y46^NW?+U21X4B)<E/:.EN/_[3CQ9aK(afY&7R]bYQC]J#Z^
f+@G3=:Rb&7>9^D-B;ACG<f#);GF-WTP-^+bIO#a^\gf;0MWM?ZR9Hf2.[]fQYAa
6J_>IF6>[?Z;&YO8RZ>P42A]dU5a9[Q=BG_.d]5eE#62>H0-4(^8.;Ea3-YV--E(
QP>KA8#Z&.#cM87[=_OLf8ddG.O&-&;6V4f&G\SaX>NV_,7^OI/:^Z(a4/8:]Jdg
,9K71IBe2f9XB)@ZY8gTX<]BZVMGYaeIfXD<9+EDBV>,+Y.@_c41ZM3X6<ccd^T]
eC>WH)\c8eW_A;fNJ(g+5b_D1;[];7FQg6DVYGEEg<FP&C#WJI6\B:BP.BR-Y#H:
e?TWGaPeMg8J0-^EgU4,HfQATM^_,;Y8dTRX:Y#V<910@EHP)/)TYeWA^LF]5_0:
<6PT4g87P1eOb^^WZ43I0I]3C[:8gX?d0PY.D:cO.+D7=HMeCPA>bJd2V7TBB5,\
^\B>Z]@/@M2;&OdXIG9-9I@f5SBSc.;]D[Aa@=C:UgT+DNfATRA)F:e+8,IBaeb/
_6?2bc72TD,1W,86TEC;V,-PDRU4&:_+]If.&-WTgM935S?QQTE&ce9)]4.;.J03
,HXW5f:>25#>QJT]5>7@0H1g47CJ.;(9&EWS9#ec6.d8+1Y8:GWf3DU>/1D?A.-g
ad&TgX>^UfX+29:]]L/-g&=XV@f?YIdP4ZfB4[.fD[+FG4eI7=VDG]YJ1]MV,8R-
f&>,<V2WRgM:BDNeRPT:I;=#6eN[eCSQF9AH#db&XJ)F-+_>?-TOZ.P@8T\6BeUK
_^(OQ^6R=<Sd:0D6M5WE>\_df/Qb3W0TCFJH@)c<1U7<WIOT4DZ8gPe0O37XGGQ>
MM74dFcfQY9-f77Z@<YXSdW:R=/2da<<;\(\.WL#X^c3,IRe7PL#KJd#3?;J(RRF
I:=--=Ed7IV6KH[>N4;X=6==b[/23)S(_WJ:Zgc.)^:4W&SCfH&3K)O9\ML./OC^
TRDGE;24M,IM#\,aG_eX_LMLW40@^7A1fY1VgO>M;AZSX+9[F?E#(<U<bY)Wc6cc
bCNZ=P#Q;K,A5gOdEXdZ>.<9YL:V,b]-/gX+^34HWV-A&6J3SB]EBVY7+-FZY7#-
A#O_G1:0O?A5.S4b1;L?WW^Wae@[gaYNH?MAaO#+EBgNFUQ@(K&-6:2,TAO]E1K5
9T2I;H-CU\4+83#a)#[\ZG71SBP0P1+J/N^UdN[;ZcB:Af1CHX.R4DOJ385HOa)/
4E5H;<Y1e25U^YT>#CBTV-(812Od_M(TH2(a0BgcDAa-POc^c,a?M/KPc_+.0f3N
G<I^(I2Ubg;b\5_W0]89]@g]1O(eT9\dSNL))[UEUL=H]W]f245ZK4Y<ZbJCeY15
1P.(<-^,Kee.VV/eWId8ZM:F-2_^.6@/8?ROE+5e6U0V)[R^/8J8/8=.>().Rf(]
/5\JNg_=E35a158g>3gHV&\(He0<9ISL65(Ad=4PgA;EJ>6Xd\@0Me++J^SPUR0W
g3<V5EQ-AAWgQB@TeUEG6D4=OL,:5Y^3-F7XK&e.>^73\7)7X4EH><G#gCJE,>+V
,ZY[T>>&NR>3FO_BBfG]Bd_J:\)9-65+-<O>^G@cg:L30cQ)=:;:4-3Aa6B?BV;5
P&&5HMbM4[=.<K]b7a1(BPT/NUdfE&gP[R&8[d&NN;1-S-&IYT[8R^(gJNUSEa,I
X>ZTZb0[CGL_1\5D]#Eb[V9V@C>N2L^RXXC=^\\)A46]bD8QQ\Lb4bH;7#GAM?SD
MOA#622#R;>Y_^MPX\4[-X+gc;e(7MM@A=d2gY-K-;SL2Cg#/>C4BB[7aAKBHN?,
S</YP5KSGLac@7?AeW@/eB40/eO0X((.7X5\YPK1M64G^XBI11-A1R3;Z@WGZ2BL
<f)MfNP;c?EbH69/P1<)N_F-:EZXU+e(&SJ2Wf5^F:[&,PBVe_]Q1#I=,;0L95f_
8Z\=O->1D1L5&?TWQ5WNN#FYL+6EUNS5>26_bA0e(.CaR:3D^W_OQ&EBH16\g/B:
,4HgZ>-VJD?)@JIe?W/H6R[74</AI4eW)b+5)MeZgSUe=1cPON68N_-7f^J0F3?-
AR8+aZSP<NAME@T[9IgAAC]dZ?09I@9TPE5:aZaZF7,d#c)UGDC52a7RgIP?@.g?
BAX?fINIR[daQX8GZQ&)A<;6Y#GRf3M7V2B_ga6@6;#=4EEI;a_J<BY\C6]b[9M#
K11NF-H>OK^L@gA2_-Jb[C+;F2&=R]Z_58,&?LHP_G\JEO;4feNGWbL-]:EDTd)C
/[CUS]51VNCBAe(^B?:\\VL9[(Z^<&(d(;UR_5MafQXPaN8F4<HCJ0H-Bf1GZ?>6
\a2,\;K>/I&E4\7TY0KX-0+Z(]#5;JSB1F5CEVRSSg8eS;eRIXTTX-\_RbHB.V6L
.ND<P()=501Y3@7(2#8W#FTR/)Ig^7bd7Q[&0F37DQ:;D9^Bcf?gVaLQ_1J+,d;0
8U4KRA2TeK/eA(ee]UaT9_f,:Hd:/;/<8V)ggD6/PB@SZO,1+bEKf_6OTI9DBE?J
&WCS(VV^U;g8+2bDOcc&gMZ]f^^>D2<8G<^-(MK=aLW^cL&04c[<&B5UeE:[XaC)
:aX1G0fEC3ZJaY(S##/d:^I^g])TNRLBTg?.;J(Q[&&+)S27VVJAC3C0c=Y+@]D)
gfQcJ7\MAAG]ReLJ,(R.d(.(eIF.c27MHHE&(d.-M]RWJ.>3b&@;#b3NLH+=ffU+
,326:F8e\J4K2A(1J1T4N>,#Y5VQJcKL75.VB23b#/EH?^FOVbOb>UdTFHbL75GM
a[ce38TJUD)7YLMWcC@@Fec86O7Hgd.Y<N(ZKWO71?R#]WIV2,<?:MR_GA.GdI4G
CX/^-QEV3#eQ94:Be4;E-Yb8f9HM[RNfK,T@I3M7?FCM@06EI0g/=&/V)-X@OWU<
1FROTU?1KDSI55IJ()KK?/W_,RfeQ@X\:(Ce:NB64\;F2JV&DAA/O=-)=)(7S?5/
/(XXOA(ZRNP:V/DTG.T>F[T_6XHV7T&5^<58UA;#0#Y6E@UU5g9R:g;]YI2Te;e-
0CH&d;/O6\Oa)b=.;9V:RK@\6B[268UJ;B_bSLZ8VFGM=IEW6^P6JS<[Z0&RUVZR
@HIe#&dWaV>:L.=@_[WO8P)8S/H]OR#(c.[^Y/JfgaW/68SaX[VM\B>^0abWR:OD
c\T@/GKS_>OCW?<JS70BM4KTU02.E]_+B>XJEI1[/OZEFRWEH&NK/eB4/O[A8IE@
75dL2)X(R[XHFB[RUO&:@VPANeff43-_#ac=g<Da]TVCUa6;Ce.Q3H1-OHA;)Z2W
\X57e/F4&cGI)PICf&Na/cRJTY=UaLGDVGXB,K(X1(SbO9fK\+?]cA3B3^IY+@c0
?H]ZC1];.+4TT.B]b](:Z;::&/IJ(3F0W3(NU1=:E:e:3)+WSY3Ic9L7OBJ#\2Pd
Q.Y<=37>7?Tf997ZM[eceGb>g1W)\(N?FMR)+@^_^CVg>)Ug?5Z[K/>DIZWD>RDW
.]bdJDA:YKNP/bL2B_TWe4E9TC-\8:/:ER859<bf&3gSCJWO:HNNLNMXO.6P0f7#
G>B;M_]EJ[D)d+UKV-ADddWNQP6;.5J/;T8NHKb>CO]^3&eT:S7ZI(X-(+L<a#27
a?C1,#(4O&e#<cI)9I/)b.OOfO=F-Ng2PFZA(=<D>-^aM_#KZ]KbeOa^UEd9_#W#
H?aRR>e4]Y8Q7EeSL@]VXceMO<?IQ;DaXB2=_S0@da>(/]BW0=DZb<CY6fDF3E#F
(A.^EAHfU7M<e:eP-?a-+>]6PEc8HWbO5?f+e:-U#GF5VM1F(e00.,F,C[NEgc#?
-7V;_27B?41H_#g+8.G2cU.Zab[GNSR[f@A(>=J/eaWKDSXB(g.O1IQP[bM^@@L/
KHeJ&6XXDbH<<bTZ1SBO7EJYVW6SBR_f+?E/9GU/,Z+#9,\(1Q.QTD;O]IF;Z:^4
]e#1Z^4G(H5S?D),W(ITb8ZTdV:Tg3V.(7.(c2aA72F48K)-eY;Rc[^/&<+cNeNB
eb1F.P>3BSBR;g;L)6P]#^3M])G<ag_EC2TB(86_.2TQYW7OIb#f&0A\ZLDF?6d\
N1IL-.Y9HX\D1BT.])B<]/_LbV<c1VGSSSUdeVS:@AJb\XC(#eL8gH4<HB&eT2f.
M\^E,ga@7;4d7&DK;AKU+KbL#BOH0HXR+Hc=U@T)5;cBcM)::&.]J9(EJ@ZG>+#D
=&[@51/cE&P.HI8Z@@[K<e5F<GRPAF&9ILQ6V]UUH&[T<,>SQ<e&+\FQ9V#0(1RU
PfC587e\]bXGU4Dd;NIAB,]Z=TY1.I4e#M=X?8PXfL499[cU_8E5M9b.SG+<@Gff
C]0B(Ua@e^?Z@N<;36c.@>C<Ic,/cLK;Q8@0DLE&9UR85P8FfPN[7Bab;e[?TB71
+fK.&FHI>S-8^CV#]f(SUJSdeZ-0ET&-B6REGH6A@11g-d-/F#TF&O1GV8YZNBdb
M;]&5R2UbW3K1GE0M[45W:C(S7])RHNR\Lf#_E7G5^\Ce[:YM5C/&0([LU6,C[;\
PNe(0RU0UIV+QK7AC=TU9d(=2(3IN2dg>V_PQ]PX^\#X7Z[Y)NT1NDaMO2I_?.fO
<JV&<OLH:0]?#JKg5ZKWZP-#(fX7[fWVG[?H.J7eC-WH\eQ0WDf#+1Q]g_UZRZ;)
B3c[a6/b@E7R3_Za).G\&gH>C;EYLY\I/LK)Q8=IfN-MTQ.AK0@<RBKDPEZ.FZg.
)ab,:V<-\cD@KPe_6Z)eC[\VgM6e(\aG1W1e9&?R7NX9/?0;N^=cC._:bZ[>7d0P
0GGY7MO<@=(>/(cCENY<]feG935LQ0WQ,-DH:AA#R41#(_+UJb)=-aBK\O30,XL)
gY6Gb8_7([U@._1:KV4Z.T/9^;>^eT;[E>@c?D6+fKISf6ASB0E0#JTTL?GTJ4Y:
1#>a@Fg6YHLZT<:E<fMA^+].)]UbF\d3WbHB6cg6(T9/cX[dU#^[7PU6OA+-::dR
Pb84F\NP5Z9H#).Q#1Q,Y+;fMOX)8ce<L\c=@DBfD]<9:#B2VER3Za/.XT^QadUB
\RH3NN5].M]@2RWSfM+FZ,b,),T>X;3d\cJZ;bJ6IJ<>VVHT[\>;H,b6O2:;QN-^
(--dHZ&9=POgTQ^HDBNKb3A<GW=8HdX0+&Z04dR8E0eY_+^(,DLFC)3L<7K+O=]F
0<&\4Wc/-&c2IJ:V)YKdE25^\c46C-U(=7JZO4fU]9:T8[]-K2NA>K1(/4gKb55;
IR:7MbA&)TFI9@HY9]S8E+a=M9ab)_MP9KN##bVBKZHKXfgg+O#[42(VQEW>G3RD
(,-RSKNH5,A)dW@9/:@&K4[\c1Bg0MA92]\>R,aBK0b<?eKaMX[#ZPbd;BS7#D1F
4Z#NX86&5C?ATaKV((Q3Q3;O4DH9]5JEeILAL,OVNN,RS,4c#LXCJdF0_/=Y59(#
LL9#,KT2Z/Xb&]6PLBb^?_>Fb9H+g:HO]1-SHJ[+B+Fb^](9-_)W?0RITV([G&JX
.A8RgEcg6@gKbN9NW,:83@[g8-eE&Z#GK1aZ\7+#&WHBGUe9)79IRJOL.eRF7MeK
^FU>O<VJbFI:D@RAP^AB^[:4P@4]W7J7@N2g@EW>cPSgNV(-/BRMJ>eR7@6BeZ=a
SOSVLQAVCM+dg>(7-RM0Z)/E+Db\T.::>AcXXPPC_22I&<EBCeK>LW[aLQbOPW>5
-NM7:;F_GL5@X](6@(.BfCaURB95D)L(@C\c6Ke1;?OS6Xd_fFg61PJWdTSHP[f;
T4[CaI5&U9ES&<,CK1\-Vf&P^EbTX8K4:eCgb?MbLUX:?/)cZZ9Ge/X:cYS8RX/f
YS>4YRGON#(fR4BQ?H@LPUKS;)/HIF]Ga>ZbRcW(KK;a#PQ=F.6JQP4LWD#;::E.
?bRb?=BIUcb2+H2O4PG7Na#V:-H&7[(??E9N^K3//L9Wc\E>0K?R_N>dGI)QA4&a
^BOOD:43fPKI.,O<2,=O_TCeG7?E\+IC^RB&aHRVL@\d)WAeC>DT3A-^+[@-d>?C
:8:b5FN+[f3?T:g0=,[Ug)2d=;+UVfLEE0;5dd6FEV+#fgf[7(WF?VAE=K0c)_GR
@=SfC&<5@gL5FE8[Z+(XfQe8^bI0IGeR=deKf]A47XBEI8S=B,0.WRN=A4#Z1G0(
:H2YLbW4gQ>-?]MG_QGUHIJZd,]Q?XKHT#Y/Q&X,#H1^@O&7::<.[S2c6;3:dN8J
,:Tb5ab)bT2)Z=;T><-+A9c[^97AO,e2,LVA:3]QAcB/T)2AegQVFcW&RZ^>H.X)
4Z/,V>8\,V#[9+)[\;^3T++;(B]dTEWY@6\^LGXYNHF^YAcEMX@D;W/GOVQXOEaV
XVdX-99+W-dZ;A@\)^J0LHFd@J7fYSDV7aW&=FW\7NQR?73+IUeMg4[2KQKc:^JF
J9^#JS^FZ=9TGNLC=T4\.EfcSLHEP3.OFS.fS1,>Oa5DJ]^(ZNU<<[9Y8SeKf91F
;6MZG2PZ6LXT(3JA\G5S6XYBA:V/75#O\1Z<].3^\/TUC+F[Z#e?T:4YC1(8.F//
Q@-a>+D:)OZ?_(Y^<I/20GJ>XKTYFP,fF-d]WC4]]TU<V444V8ITF\;:-ca/8RcY
-e8MJINe0#3_75R:cW[B[JDVX>83\E\BYFZf.U2E\#P+[6A/5=A1=OfNKWRF.9:6
V](5Pb\(^KI>PE-X[MR_XA<-Fe6?0-^&VLZQ<,0<B)MU:K0J-gI()X3NfU\@ADgR
:&EgSH0>8GeB>g(61SE>)0],&1O9Z;9&c,Xb^?M44bgK&dFCP7;96c3cGS7bL\?=
7/Dg2\5HXQAaMJNc)fN7TC(F[d\SeJaH]42&PV\d.;;1_OH5aZSa;KR;]g9(MV?X
Z25HEU>/[JW7@>adH3R=d=0JU^/[T8\.=@GaB6SO3T6,OV(=3MJ5MY/]AL8^,1dR
F>KHL&_P#aJC_P/2U#bD2cP:]CMA\(AA)[@ZYf@)bF3c8CQ)Z7+e=_334/+7E),)
SKS-9.#;B-B_8KXf>92V(fPYHESP.>9,PLDVPVJV28g;<feZ^:3+g]a\3+:_7-0f
gVd0-R&]25;B1.OEf,P]c#T0-:MZUP-Hg]0f94X)U#V,B-bRNM1->Z)HLMDKS/Z6
CeDJS:L;(N<G_eWGQD+0F,T-^_2/<7O+T0V?L/&NS4OD<cZ7dN^B_0OR<+\Z._^<
IR&?Y#UTF^LD34fDR-d.WFN(AQ:DPOU@;V1eK6eGS7ZY1[BL2/:UfW5db=>5fD1Z
NFMH.3K4#G-R,^A7aK)B8+FdKX(g+],E09U(6VA2.\F,c/7Q[>ec#HWB)0L[MMSY
c0fV@FO)D3+B4#Y5SfUa>R0PR[#1dBb0>+?C&H/7Neb_eH;#I/@RQ#=J)0>,MT-[
5Q,=RF\2c??ZgTK[AZP&/[c5H5#<0)()2?3SeVTN=g)@e#9M]\:U6WbIc6d_UWRX
8<_D=L/cJ/D+0LAP9@L\C@BO<>7[,?;IN-9ed.7bZGI0EMWEZ>(B5G?^A=+Z38(L
QKIMEeN.:B6G]Y+@W.0?f2R2N0F(1/<-<=M)](c_=933(>2Ec<e?L;@UOXK;Z+KW
-G=L7[X=CMURA=6MYR;GX8WLWd\FOe90>,4bOB)>DG+G:W+294O7gE((D^>+KQ8R
M#XcH0dUG7J6@+a78/_+;M7&<[/6:]CE9c=82A-_gWFZaaCBZ3Ec+1IYA^R.N+Hd
Ub+/CcF[dG.1B4YfY=G<+8U.@+d.9bXQO-N=a[NXKP](P>HN<JBI3S[/@_@S9;fN
1S40^S5.[&Hf>.eZ@J1?@<(#R-OC8D4V8[@&4YYV]e:Z&:D)K4Vf<OT1aX]ID.=:
J4S^Z+AeTNVWFc13LU+&b6LD-:6cC2[4&-^<[Z<=+GL]U8:12[X,XSF])ASgWfQ6
CINc>#G@K^3g_T=e>/>SM(3A/.dG4QN>b?)BF2PYC64SFf;M2c;OYbS3UCGYbAHS
-gdBKYL:a6LW8#OJ4.8K1H4]VJMd7X.7,]ac?GU/F/O/H-;2/L[.e18X9HH_P1J7
K^#,>8_;&3UVG\(]=M4P]a.<<7,?]\U2E;@K6eQ+Rg,gaOd#1VX[X?bdB5D1PV2g
d]2FK+_?[C+F;1M6X:5U#2[fbVN<57DVH3T@:JM9CeLHaFT3XHRQ-ddRB^3eV\O>
(_g/0Rf3H:H9?:(Ta1=/0Ig#QQcKITbP[#0H[f?UCQb^[d]DeAF,^8F1F3DBQLZ9
Q?OQ:FZ]M-=844I<GdI[R5SV:bMC1YbL49?gRHX^b,,TONb82[<Z1L#AM]Eb[SB)
J.L\U#.X_gb3+\[@]E.QAeHOQ=M-?e/Wd<C-3AJ&MJ=ZZ).N#MOa7Fe/F(YAW0PB
4N?V==<4d]314<TGT3[LF7+J&/T#1IW;-Pd((R]ZMG7D+,OCZ:;DTXJ@HOF,B??R
MFc=<_F@G/YM14V[)c33]dIg_C>H\YF_HW69.+eMccD0B#6WT/#d;_JG<H]S_f+E
VdfUaTV]Bc/1M7^28-#c[M#XA?>bMBa2U-I#e3/e1I_(g_S2eS:A4]-,gI=V)##4
M0OYcEV0d66OgCH75L]N6]A7\&Y9C9(?;MFJ1M],6,_A;DNS,/OG#/TB0eC<)>UK
]/_fbd,++&aNVAJMKL<:b#KB4@O.CCMMG;1+)P5SMa4-)0R.(WH5M@c)##VE2R]?
:O5cK^D-8([fbWKK]+)M805H,NT\M_SH_e2.98]XEVD94DOM\Y71+8BAMbS:,=MN
>J,bX3(J[:Y]Y8,86Q_a6HBg?\7caS8L6O5MEF,EE.00??AHcW:=JKe;</,_?fYa
3abNLJH#bNbLG?]-cYH?=gK8gWL=ZRPAH-GId(FP5)O;?ONRIQ.@]8N&QQg;,EDg
]I:KTO:H^2M,XB=(:LZWJ0/,4QgY^PHPPM[HdJ6)Ka;HFJMAGAZ.GITf>JdE@8/Z
IEB6Z,88W5>73#W(BD#SU#^FU+0aXe0,O:D7?CRHdST4-g];+T9(N4H2,?Rb2HK0
]KeR/bN9<9\^T2OJI]K0H:IVC8G_KP4Xf4IF\:Y]X>+J\@)4/g+H=b.0V0)1/UX;
94#O8C)VICX.NV7Mc02)U(Zg+9B2]DJ?g/bDD5W9BeK]ZP?Y\)O^6#0K+:.eWEHe
g,3#&K)[.480-YI4_e,7E:5V+DK]UPFH63K&d0?7-\P6=CENF>T>F8.GS45)_0ab
@EQKg:M/3#c+Mb#@T16J>DYVX5g9g_G6?MPF?K=f6F22f0-CE0&_@MaN.6Ze#LUa
;PTBXd6O09EI800V08N@]>#:aM^:bT5g_f6+.JE;PZX56)8)9>V6AU5e9aF<,C&R
1FcQ<0#_4Pd#I?\Q,WDAA6#T]O^/#J8=7?C1;BNCRA/I0F\R0Ed+;U7UYM0EKDM-
5EMFO>VC?Y+6Xc<+(^T04deRCJg)O>g(I\I(.0)+>VUB8]A:0^.dNB>)QT,Gc)2^
VSE])H:\4Y^bS+9C4#?F]7bd4W9;f+MUCe[cX&UJ<=WN+K0A]9IGEAePG3SC?LcD
<]/Z-WU;[g34IZC9)FV.(2GPO\@?U^)PAF=P<;XdeUG;W,\4G2-V,7,^KV#TSX&(
,7[JQgKUOZJ:A<e;]fd?K:_3DT6V)YE\#&;51K\F+DEa2f7c6SPeTQ>]MO2W^;SU
HS9HIOJY6(1&Q+FA2FRZ_;ICbJef?B/?65)=XeFS3U>59X.Q=?K426E3<[@-bJa_
233/82QVL-9g:2WH@P3.:@2a?<5+@#^N-bAQeJ<^bR_1R:+46K>ce>f/OD:Ff]C_
ORc4Q@[,3-U<6^D<D1VZC52QU[Vec6\:-G<eS\PIO=gXU9Z-6)R]aLDAf+^9MM5d
3JK@U=PW.@LC]b>a#+:.<)HgcU?^N/M<KF@]V_Y=+Bc87GD>Rg/aW8>R#bRaUS7(
]E8@e?MfNZPEWc;T,9acM0beQM56]V6fO/I,;d?>]&MQ:TQY;3@Gf</.Q.49/ODa
@5NG+6I1d:#Pc:@R>;+^4/V^]=bR.4ZW&aPD<HB[2KV3(,Kg[+PIA[?<gAG>)dgS
LY^..V1YC6e7Z20\M:/a#+V[fGM49,/L;/;M,>4Q<U8]-L)L_C^+Y0PXZ,9BCZ1/
U(&3,Y/eM2F0)0JPD\8Fa=[b/d&<A5D0LJQ2Pfc53&0.Z3MA\DZ2_)d^/6;f6U+H
(,e1^EY/)5R1KO+GH;[K;42,W[UC+7R?GKAdGCZO]\;DYg;8DJ&_,SDE\#P0F]de
]T(c35FBJ)3P82A5c@.C\Xg(+IC#dK<aXHI-M494^.3Z(Wg/Y^&ZL-TO[_gV#3dd
Wg?(0LG\e6IS??:LY/=1V(I)8)J>VJU24.?K+eX@<a+E[N0b5TE?d=/Z+JQ+DP0f
4K3gS:HU#:R<J^.7NE:C::d0@ge)/:[dJ9\1ZV-P;D4fQZ5F\E&S;IR=HH:VKN1B
dg3Naf/EcfDK3Egc&J5(V,fEZQ60]Q;g#3?2>3]X[;T]4M^ZE6a=Q:?Ob<DS<SWd
I[T<MIScd4ICHbdRZB[]<<OM]?[@+?gYeQaE,<QBZ&WY/DU)1UgD).P4-f#G0UF3
18MaQ@S<<.(<N5=L2F^?cPAD1?e>=K>A24X\G7WK?<gK1E:4+(DDcg(V-a_G9eCR
216e[S/;F=eR0.25PPYWSH7@GgICL]EDe,PDVf\Y#W/a;d)d5?,N\JGQ.+RcXO[_
cLGE<5aM4]>PU_Q#1McYNbIUW=aTQ\=4^/g:U1,^EZ1))>KJ-)NHC6IDNCGFEd[7
9)YD;.?#?4HfAP:::7PUdT62@I5D4EE]cOVWL=Ea<2YN7WCXV[4.+(]9[RM/>IKY
#-8(+fBRdT.Ud5VOIbgM?R<b9A@LLV:]R/RM0MfgQd;+@;&f=#43C;aF:F^D=JLX
XW:GPPdVgYAN_AMN&6F),.]B/>BBI\VO4&aU?eOa>25SFEMcbL7&DS+&ND^@<5HI
D(07D]BSG?.DZ#UI@0\Z+__),@CX\\cT@e#bHeBR>X#IOA-LXc.(\U6?:,Fa<EZF
^L\UI03GS:=g2^Jd927dE&1YJ;S(c#^=A)bAA8V#6H73W(F9A0+ECH^[N>+eUfYR
XaQ_ZLGAW+IHFB+6HVCL6.IVIe/]_JYW7<4\?C6e>A4MOOZfD.Md59+<[^),f/_]
)Q)@3\gD\G]/&)S27R^/7K+b9[[[53I9Cc6CWJV2_^QQ2FRM(0g<L]LE^SIDe\N-
cNH:M^DGa?Va_c3Z#FU\_]aK:H+E\Ed]T(+Y+d>.3H]29f\Y\MF&7U_+ENLa\:+A
Nc^VJA(5XOc6FHV[ITef6;F)97M5(-F?8)dPRW(Z46:c]S?TMO[&EAHP/O)?6U]:
V2RIFY=<B/5+.5-LPXV\J?LRK9OE.GH;A8^]X0@P-Ha/g;Sa=EEBfXg^Oa6/Bba(
J0=4TVM4cC#K(]:d)P]Z5<<X8_XV/03C),[B0H?Sg3Z6Uf@@ccT[FG/=-<d<80:V
UR;XD16a+ED\4d8Ld<?WU1gdL^5YK[:d:1YD[-8#O+-ZC,>E6KK0+<:15&DR1P1&
6Z4>aPef<V_aIQKd9VTc#)XEK#?BM)M06@9/0+0->+5SQ\eObQ-Zb<&,eOROZ950
&A)ce=?0PPc)AOZVQ^1MN(:Pc.ZJX?Df4QS8Fe.G:&&,4eJaGa>H7-8YRJcG;=V\
@]FMX_V>Uc]0cC=eLcd=,E2c5e\U.6CF0:R18f(3)^]V5RITd;J_KHELO;H6W5R(
LdEcC4Z<TGR?/+F2&Db;XAKRg_a.SN]NB6(_;[Td/KWCQ484XFS=&GI]aP/=6^=&
:e#.7ee_=&dG4Xf[R/;+?c>[BGI<UF52Ce_R)^a@#\_B@R3OF@?<1VF]=C>A;[a\
TO=:Te>TV5TK]&T7:U<QLEU:_gV3,RW3eO)CF,LZ#=QC1\b0(BX.QLYZb_L4YO/)
-F9?c:;?g?@-:AUa/;IO>?,[(ENRbd6.4W+Vf/L88&B^3G2QO&JE#1>_LEW9B:Cg
;a>H:df@.GLILY.M4HS3aV\eY^5>#50-=.&:/E:DI^D9.:--#8W@K-.^H#N9cKdG
8Z)TYVO#=KC,P;EHV)8\AfN_.56=?ESZSR.2)8X?\cLM):I+:^RN1J@BZZS4EWV]
B_;cG73H^#a8463T4>K:N?V\&>39/DW0U_OUb9#Gbd_U(?UI4EMFBZ77+[#gef5G
-GXYBD0Zdc<eS[3:]+ff61GcMSRI_\Y]@S1f@R54gNI21:Xd5X(_00V#&@cOZ,d?
JPabFeMLAQLNd]#5NQ&EIK]&&)F4>PGC?S70C>R_3<RWS2O5LU8..-d80T(9A:B5
@9#R&.<^TR,0?dL)OE1;/&cWM_0I)J+;6/I\8Q=gd,:LJZ)L,^aG1RY]FR2eKL&7
04aaBPCUDLF4gPd8WRc4c(LAY1Y\[W:M=X]aX5^O@#d(IAF(YG?(acILfFJD&\Y@
OY)JVZ+e6CBZM.R)c3)TgdPI+[5,JY=HXZ7IUT]//4V+VG)4(I_^L1f&KGa?/N&U
/OI;b[ZS&[f(@O;M;JHD3^))Y17700XbZOFMJ/)d8^:X+05UA)QZ(b>,VB\,,LN\
4[KN^I0B\O(\K0QF?;M<KA-SHf0X8f/)1);_Zb/@:V-cWC0EC,S#QdO[g4Z4U:=4
eab=#C8>D#>9e@bMRKe:f5-YZA?O65_K>;=5gM)LG=YIJU\eUaO?>48PefE+/W4D
1fV?49;?(#O5BYU]C/[2C,<C-\d(;&F8;M>R?EVE^I3#LNe-_aH.PN;YFGE+9<[L
#5GM;(]^TL9Y7_\KXXYLMQ<0X-<)PJJPcP_:D=dKDg6DdLa?(N.6,dWcE5S]#(^L
?^f]1UP>N:OcD@/IUHH+B>::JXA\</E[G6/E3^Q3N.:9ONPS=Q]UG\#E\3#:.5TB
c[)@OZc?,;e:,T_TAQc;ELFAV_+1]4,-:EI.TDf?43^0?(Uc]BIWX=@T?X:XMVY\
+^Wf-,eM..=gY@c-]N4TLP\/9c?TR:WAIE\UefgHe@;:dBO7S+4TgT3J?X/,7;@3
U\e46f]&,4B=H-@EG+,V3OT@B>2+]HK\/N-bb&dS2H6fHMg<d+K_D?INeZTHc;PW
gJDG.d703@^X_6ZH0(4S]-J++<)KQH:@5SGBc@g08\@eUA+/QJH6X@7U;0gPZfDL
F\R9<,SD\gNO1OX(-\D5a=;FPc&WbZV&-/f]2JC7RN59^<W\HbU(5Gc6&>;1IgC+
dV2#aO^_SQ,_=gYTNESL/_<FO(HGb).Q3],6F:_/G(=H.WY7D,:aAG.O.S/1]S7f
+69,GK4YIY&F&NAR+Ub,&-8L;&A=)<=:C;Y1]cc./aU4@X2,[KKYZ7Oc?0[4;I]e
/NPM.01fO^<+TZceT^:J4F)OXZ+D,3e&AEJ6OcNAZdUOK2^7L;0f+AJ?d_2>gI1F
&K0BR)D9V;N?9JdfIZ4Y?#,EV9ZG1J,8X-48WCH/P;G)S]ES:,F>c.&I(7;0EV6b
T1cO01gM]T]./3HIZ_Abb>Y(2\d&)PQFEE[9Ud@>N]WY/GbM>#gT04G8=+DDMDWU
,M-J,+OfTO4I:@CPKK:fSeg9+f7R/BJP5NY-[F/CCSa+<A9V,#VBK<9Y#H)4:@\?
0Ef^(LVR<Q(H00^BF+0D[/6DT;_C9,NGB)O^9Idg5CEC&A8?&RcCWH@HI32UaRZ;
GfH;Ma(^<#-Lb]E/c.@F07LQSVVM1eR6a;b8F/P\;0/=K4)dV48K1+M5;b/0b9b_
EA^1-1XIfJL,F5(e3OeU-Y=/-ZH[VG0g[b)UD=N:]WC_1IL6NKgK05,(QH\@[5B5
L(A&]1AG^JQ].R69c/8#g^cR.HUO4S/SN;8[#4G/FEU6McN-2K-_9QTZ4ReCP7)M
C30,#PNT#.g3EY+EMaRW9L3A_&05aG6E&cF#]N,BfIZ;UV6>U[Ia7eSU>g;D:a,L
II10Z5HW0C]f4=CdG-VTXgC3,]\JZ9,T3bSRT@>[C^,B;GWcU^,(I@eJ_C3eGQNS
\>@^+/T9;W+A@fVN(&;g>.<,#O7-G0LYG(.5[eP>1)W-gcB_M>>g#>3E(fQ+&3_O
f4(f8OccOg,11#5&S_W;=4g=_7I,/,>KF/88AZO2L,U=VVKfKMTRB=R]?FJgfeOP
/)Ef@FO=#:ZE13P\PW>FE?gIdaD6S-3P(+-_G<),]5A6e]:^04QM)7Va@>./;=H7
92=gWJB2@T#PQfG5G+::OJ+:9V0RC:.HZ\A20,AK/\UC6C0aH)&MNRZ;@8N7&/)W
M)gaV#MEeK]FB/eW/GK9cXLRX\?3Q),VC#?f=3abNQ3:,HP<]RRBa0D;P.&>8gW>
VB(:)<&;1Ug)LKEJ7O/V\:a86e-V48b0]<7,Gg[FP>BWU6>AcEEZ[1AdfBGe8/)J
VRad(L0-_9QfEN0_)U^J^&G3F=b@6K\(:f(H;\_O.Qd^2A#X+1R3_I3cAQW=J7?X
d+TR@M[?ED<A=AWeccD>,f#..WZ)>]ZKQW4M(^\bWb9&N-<]a)6fe6KLQJSb8E8e
B_e+.==E\PQ:Ge2T;,LJ=LI4I>(I+NZb2IGd=O_S@W2b>CG0.UDZJ/D&X-W7UKP1
aBWP@/cX@GT+a[2]Wc[I@DKM>5aa9__2#,(7H8D<M^/AU3VCU.[g(J=M?/1RXD=Y
<+M=/geX\eH,HWPgI5d1=0KZWPR5K=PdSD,9\B>RMRPa;JH<?W1RMVBTY+-fC7/O
0c\,B\<-,Q4M-M9BA=c\U>9fB1\F5>:_6?gBbff.MU39[2JOMHDMLga@&81,XJIB
9D-MJU)ZR:1CG-@H)JW[DcFgJQHa\ZG9eCV(5X=W79eU,[.OWD?2=K]gK\)E2SNO
e^I1KdB?;69Ob/>dZf?GcdERX<9D,SX?c[9O)98M;/N>_B[]dA6B.R\\8cNfG5[)
fgXaZT&]3W.T:d0OR]]E9NB/?ME3;BbUO?ISZ;>8)PYTg.f-OH_HD#8LD<U\W+2(
9,/1F@H99fCgQ4?V0VUT/QFMcTN9/_U8KTINcP=g2cUP.1X@/aY))g,EA/NG+gH]
>QJ]JeLL1S<;T\)RUcX48=A:Q9@@60c5bQ2&IZ-5O^W>NAb0Md[@RV4YWe2_@]^,
QJ[gC+LKWT:#+^+MgcGN<fL2EMdOYKg50YP2J&&?bDQQ[3K_6B#[JCY?/A5.]L+D
,<P2gN)dF/P7.4BW?IfJH@H+,-Rfbe#GS<Wd1BZF)PQ:>@X0]6-g5W:<?\b,IL^-
Y#(dT&Q-#;:d-@G(U##X,\bE5PcPKeA7[RAN74KUc7U@4S-LN+fa]R3P(aMO2fbA
YK(5O\2^6R(\<.Z62=0-D.#9MT\c2L0L=^Fge5fQcZL[CKM?,d.=f8WGX#VCB;Ya
2B?4beN6;YSGT7Ca-b@ARb@L)#3]CE8]dD1N]V[BY[P3LR^N>9fg>D9I&Q@aN[7E
+H[YHO?CLQUb7._dAVE7K+WL6S>^_Mf.UM\L)JfXKbVcWJ;2_9g]&fFf7<X8R=:W
X=<GO,BO9<K4X(,MCN\EC)K3I;__0-F1)C6<&NRfE)Q98ScU.I@eV-]CMafF)Z5(
+V-+J>TWd0#8QIYIA@:0+HN0.<KA2:R4K#60<AZSEf8P7Sg7JZ;gV<)]\;&3&#U3
7SH,5D28;])Y1GPN?JVONM366d/Z:H(E#0SS_G_WRQcA^LB[&gUR<>]R#e#5]8JH
J2)_g8-&EHf09VB\L0.aTc4L16;#ZK29)Z-EOLNeXLN_/D2TJO?\g?YEC?9SV3:6
a[T6BX__]VFFgM6,>5RMUf:96N3</=SPL@>gE>/C,1bU7^P\#DA(RO?P.J0F7I-c
3\D\[Ca\(0EfdBf,].R_bBJ+\]1UM_TVZ,a5JH7)ER#HR?;^3[0XON^<E4d-K(.A
B8E(.6EJ,MI2KAXQ]OeGRH7.N/f5Q7gN\EY6/O>NBFWRPBGI\e7OAS1@1[JcU&(b
UgJE>c,/:38AFDP>[.9T95/M8G7gF1D=gU&3RW0;dD0B9HB5P4ZA;A&V[2)2?QTY
Z#8C>OE#F7&/\g8GPL./BLZ/EE,ECOILMe(.WX^6E<VK/FC,8F,C37dG=U,RfJ\@
3V+KI^?Z\PM\\M-<aFCd?9=__3PNQR/^4:3.::N_E^L(L2Mb4/(3fUX)O(,fcSD.
^X6LOT6LNT8D79GKK)P^<d5B]C^[/NYdA<,Gf2+Hbda3Q9T1@-[I-.]Y(+:-5dP;
,>ScV/e+)==\X?X>]JK8D(,^R4TC#M;O?9JHJ?<,IS=E?JZ6#[[Da;SF1_ZNc]Ja
8>=^PO/-9\NQ;PRHPU-,Q\OH(W[O,2(Z<08b/1Y_T+,MZGE2D,Q3_XMER;AJS._B
]?=(H8E&Db<IfO6S6_)KeDTFGd<_HC?EeP>J46-0KKFdTb^+GI9RD)cEaY9M?f9I
XEKV1e/QINF>A4c=:(K4e8/N@G+BLY_5@F[_f(ZBRK0PJca21G]ZgI2L(d5J]>UW
@1U2,C19#D_a+aPbK&3G_)T<Of<O.bTH.9C22A#)16I]TGC(99H08DCZMILPJK0<
L>B8+I(>2BgcU;3L98?K9DB8?I>S81B4-LQHYP6G-)b8#cL<+#[0cQHH8<XL:Za.
)F)E2Jc0F<A5]/7=GY4dbC:N>8>^2<d)X<+9(Q@W85G>.7B8^E+5.G</5L90HDW5
_-2O5(<F(TL4>@]G.<-;>9B[a8dBaO(f7^gHJ,2;Za,3@>>#bc0E+ZO:[5-(ZgYF
bF/31CLNL2[<:Y&Za-B6TTe2e8dP2CfN^SBIS(=UVF</cC)^J6W4B#7-V58Y@GSU
E@a+=,@.a&>Ua?#=EA0&]c+Db7\G=^0[aD:3G?/R0HCG]0eOH+TB<ZJ=eL&0.82>
65@Hc5Nff45D<W\a^[L#[EVYDN;)37bd?.\IP1Z#RLJ5g>?J?BW&H+^NBe2I&U#5
=22=:8WVKfZe<IH((4;=BNW]YV/=7OW.U)Cb_Z[JaP<RFdV9S1BM<UIU)XJaNa\X
f[&GLK(.,>MgeBeb0F1N#;97gdJBD/RLQRM4Se?A-Jb8eDYeE.Z]M-b-1:ZYUG/B
3T+L\8\Sac(d5F.=^XN=aBLD+47dW<3[QW149TJaFg-H,8>M6LS-,XMBB(WEdeHS
.7\Z>8J+HT/9D23&X-GAF3#dg9H<QC.NZa<a^#GN4AFUD]B.bC5/ZWA-C#AP)NV@
?W0.[>FNUA/)C\\[FTKJ8#<K>]U=9(<-&A:XUWge3>WO-1U;-=Q=__B]+H8VE]H7
<#?ANE40;[6:=7OBT^0M:#D&V833QXR>ea,?MT@?FC\fI=6JKV2G5#Q)[86db>^=
@SV3a_Oa9U#Q)gZO9)Gf2(Ze6V_R0S)aKH<RO9_A9=a0TJDaK.G^/^9KSaLMC+Q2
YL-+a5JZgK=8[#VRg8^)&5V@fd/XKaTD:gC0]cI6R#C4FZO>^Y:\ANSKD=8MPQ3+
LeefM#)KgJ6D[U?a)-@SXRE,D1181WB(C>U_ADI7Oc2O\O?HMLU?JH(8)8e6,CcM
A)1(.#IR=>4&=c8.16+:9K<1=URTWVC69,27a2</STSfGSNX6c7Y_94V1YYR/KC)
_VMQH_MDK-DU^N?]82OMK(Me/MA:I[B[>IK,_Ca[\B)cg3IM1[7X)7Y3>^0SBW3\
gT.YO39/B3KZ5LCB@27O)C4#3GRd2UQ0C?PY^JCG[.1VVU+X,70QC_FY&K&Wb:5g
)@(6,a2ZREU)-be[[Df(Wg&_>]#W6[/>N^4RdDe75/22ETMZ9P;1;>[Egg[(gbT?
7?LIU1f4VT3)0@_+9R:T0\c^4:[&7;W1SfL;]#PD=66_M[^c9D)67RSLNCEI;,0^
B>&?.bR-KN,0QO=YL-.[b5)9&:#-K\MK1EKOC^5eOBD(?[XEUUgI([dI+aVU5:OG
_B[fBNPfJ,&bRZC[-?9.-Z+^IC&^abNVd#>[8g^22=SRFc(#)T/L9=&BWU_//:F8
<78#^OO[a2(E>-W.QY-Cc1E/5:dH#\X-=LbAIAG]#MB\5;dMV4/fFfG=7C,FOO?A
C7eB)a6U5ZV/FD?D:>Ua2cI/.:=CQ7\.54@D/bfYb)]O>;N-\#>;]N>,HYQL./P;
1?R8G0H/ME8Fa8/76A^=eR_gTTVSO5[Ic.CMOa/E61Ed64a<>4+NOH#W0P^UbGcX
.Kb,EcMbMc@R#IcB@\/@HP?RSOXB=+DI^g-,<Kg4=K+N=gHa>0g)H#DI-^+1CQ/F
1a?Fg<:CEK.5QADGXgNTg5:Q;[gKAW7_61RAc/CKJS;KK3GO90W1XK5M)TSJB&H(
&Hb7aGQ;5\+FCbK2KUKI4,Yb_JHCag2TI8[A;?(QM\a>3D?9([DQ.@/=-X)1&b>Y
<e38L=L9FXa1)THRD+8P/CfXP/a&b3LY;MBN5[S2#GUE8B#V/?1XF&EB&Z4c0K9+
cNFTaDGUSMcTPM7PdH6a:F3)GKK0][</^BQVQ=3=_g2g^;1e..)P4_XF\9A)/7[H
g2g/+SbSP##6:UA86a\^OWDRWA)DU1LRfI99MeU2Q,2G+59<RXV8-7f7E/6)K1dG
U)P]_.NfG/b&05AIN[-+BS0F.8I[[e.Ed;C_KXQB8A6@Db^-?V\W:]87MHdg\Ea.
=KcPK(M8FMIE00LP+<X,/3dCbfTa.:F@cd9L:5>)TU4:(W?cc1KGf.8:Z;0[W8)b
C9#\GUCB#4M3^d-Eb^O=T34bQ?NNBJ(1)D4ag[f./BP9T?C@5FTY/eCDe&YR.?GO
<;V\@A6U,a;36O?a)&Y,PZ_1G]I,XIIXKJP?;KK9;?V_ADFcW2DfP\ARJ-BAH#T,
CcDGS/#b3<_WfJ49d,5SYbS/XKQ.Q^@Q0QW[c::;1WF9JKC/BJLW1ga/_/bX,VH2
MOKa-K(>)L,@?B^C\,POd;I-cZT5Vc,beV>=g#[FD6=-5JM)Bb()aH48I2c)CH\\
d1J_4G&4[.V@XfB]E0a\gQ3ge1CE>R?^B/e&EW7,^DYBA11,FF]JO/V8=HT3?H^B
=@N?e)PVD4cdKJ88DG70QQ>:TL#&QN=<&5Md.?;H64]3a0P:\9H<X7BfUX=d<b&9
c_aXJOQ0N:SAHKJg#6KPeZ6WUZ@\J<-L+e6.JCNCCI(^f^&.;a>FPc/Jcg?&.^W&
Q/@;O@3TG(O7[9A>ZHSOHLfJ_WWO^H5I<<GRAU:g]Te\K37IaHc=IBJNDA:^eFYR
Q+,MT,3bQ&FdEeZLcZN+H2WdHTT6C1PP+H;VV&+VdQ/,18N,K39b14:.bU>#J:TD
N4KCaQMA(3,/bcVb8]eU0__:+[F;ND/8U]?URD-C9F4]A?L1(_407\T(e?ZH,T/P
8WM^6c-DTP?ga:,9d2GA(](RZNMJ.b7,H()BUL4dT[X<\.d4ge27@?SUJCX/:cDK
SW>b8<a#^ERWASR3TFLDBM2@5bAa05_BGVMJ7Hc<0\6g[(7QBU/<QgCX;FfJ&52=
0NC8G=6f]dN).Q)N>]VId<-cO4UT886D=-7Z7@a40aL>O]_QU?Y?#H5f^aW:b11]
F6Cc@4NfV@_3cYH[>-;b&KfZ5MG;@]23BDe]=#SAX-f>8WYR-S,AHLG@fA;2F\M[
[cf[]faGa>PX2HV2-TeMO_YZTCD;V.G]CRPN2IgSCW/.Cccd8YEAc@Nd3ZR[JMg+
0I->&IaNK?Ef5H)gP.OfG=9)=;[.Q^F]B?;_a0-(1.G-U;^.VC14S.:e5g6Bg_HH
#;eT#J]fe<Y,eU]gT9VY.4[K,g>]&2UBW4W>XBU>0^A,Y8(U&@DBTd\Y-+C&60(K
8OTgC.00]Q]ceCX?=P;f+YQ#7?_c\2c]DK5M:G<CS,Kdab;(VSc=59Wf6GV:CN[5
JH=^B,D6F7,:K?D.a@=g5O_WIKL[ggf5Kb?eB6]NZ8fcfEC&c]g1^BE0TS;DB11N
U-IFZ+<#]50Y^+(.G;4^aBY(J0..7ILV&9AG#AB//gRF;\K9Qc=H/CI;<LaKXLEb
VOCa]Ib.Sd#G@DgJJJ0D+bJ[Va;Vb016<^GOe;=c^B2bWJ42;-V-(][JN:V:_3eI
NNWKf[d^cSe=+EIgW_]D&@VH^_ARF)<2VWYFE97BULX0g5>N,6:BedTQQ(g3JBf@
B1H8U,G4B?gQ6:WKE/3^W/LQg7I(K]&89C3HPSe&Nb:FUVIKZ5YUf;&?ZW.d1=&g
@J+WO[QQIRAM1515Na(9MZ;Ig#P:)^,B_#=dM?GeF0_][M4V:MFSc+1?2<d^)U#g
K19(e,C+(9H8g/4T-6I)9@2]5B<?6A-[/aK+c6dC.>,+Of>9&,@]7:RY(1cfO+Dd
=0SEd4^A0?Jc/]KZYa(@#0a6[17@XSQ)HTGZP#4#^/Q,gX2;YeR2X8UWW[Dc.<K;
CDf>.0U-\^=>eQTg(1<@\gB+X51cSAe#7LcK4#.HTgBZXM?KE#?14#BIa_O]M]Y1
QR4_L.2LH9WfMI\CM3+\.ATdHeJ0PW3L]7LVDWO]>M<H+9G]Y\;YC2D3);]T](X+
VA>7f23ba9A2&5Ia(S^()N=ge7+0?XG0]>3U>bK(6G4W=ZQ0O/.>4gR#CN38YG3-
-7H]O[bXC(a;B<=<F0,bX#c^)SM0JUL=+CGJc).bE:1?Zf,:3F5R)HNG,K<KNP1S
=K-WgAYZ9&;0\:1W]BeW]P3E^YgTN@gQ[=+W56Z[VAOZ0aXL6>8QeG?CF7=N^fQV
D??J\X5]c24OGg6@e+YAL_g;V5M9OP/S?]WeaPQP9VgaNVQGPU<G<=>0e-RTBIV4
Cb79cQ-GE#IB6;Ff]8:^/HG,UNY)W,\<-P4TY_YM3CAgNLB[d4WJ0ZN\HJ&H)L3O
JU-OH5R9N7IdNbCSZ[FRY-^@8S6Y>UWX)VVD_c7P2)2<V0a)++BABbg1K@I,dQVU
B;F>?AUGc5\34#^+X)H1KIGH9Yf#aEA=VMM1-KS+Me_6DG6d);gd8Bc)b>=EIFF8
:F[SMSGYebKHcfX.?Z0#868^DSg@W>-X7J>c]]@6KVf,;_E-D#5=)-@LJ_W965YA
>E2Gf]0fA.a5bdda=X#/#5Y1-^<7/NcN)Ag[<PH>RW>&L9_e@8V0MD;QLde5?3ZF
5EM(VG.8b+,[g=)FXT[>b7TaJb_<O<>GQU1Y8J@IWRV6WB#eANPUGb_[Vg@c6@>3
VV7d=>=[&TRG(bNP#[UP<L(V,PC0TD4S@+A8NHdW;R4I#F@dMbU<GG<3B4I5E+([
=JcC3[\<^YS@17d#(a3I3[M,EONW+BgPO#>7HC3UbH\[&5+?)OLQQ(Ca[&DV6f\C
X.\e<1.82784IG\UJ]5,ff65JUXDN4QYXS5;1FADdb[XV2G@>)GKH+d2-#Egf@]X
<HG(],Z#NfMH7X_):/DW<]/@V0Q^(#:4H4gcS177,F9IO0PbKfC<(<f1-I=C-a=G
CCD-_1GP4<\+#G9N\a1VYO-^_HFa88)g<bN=C9KT?1Q>R<]=#9JTZ52Lg1<_I:P7
)g0d3P\+M+c7eMX<L22=Q@WN&LEb0e]?ETH:/P0GT8YaDb_S.NGA@b:W9/FK:gE4
<SKb=\P,,EJ(5I=HO.d&V<I-G)9O^4g5:+/V#7N]/^FR#NS-;R?(6/2F>CD7a1I+
C=NMea8<:^CK)UW;AeZ]DCL#HOd)Y.bf4^9B8YCZGMM)I&aD7,Z3X&S^W-Y86dX?
T@HBO[P.BFIO;OcZ)/H<)R0>(FA:e:OFc(Pc<E&=0c>UGbG+],0:deXS?,^YU1ed
CcWaf31;W677(=T?E]=bW;)0DA0#M6.X44@:M1,H1(8S\BCCZ2<^Xa13@]95,Vb<
+bJ]WKTc+,)O_#,.HL5([/G+\.7#74gda&OD:TE#X>SC&)?9W:.U:AGAc;^Cg?-\
8;SLIR(;^4-5TO(1+JM.9VQDTPM,Z;NN<76cSH_U2LM^9#QNU?=3>A>c7YZ:4D_6
M4K@P\H87a8YN3FEB9+@)RHFBDAc@J59WS?OIc7:?/-1WBLb=\TaZM>^L+5[I8+P
M^&6([\]OOKYLW7;e6RaMG9S\OU60UM#dgK3Q[=(;ZBd6bS&Z8NcR[GJ\K,eQI]1
RJ(Q3Rac13U2-)^fe0Y-UVJE7YD/Cb9>H7)e#<@1_.X)YAQ0EUc#50]5f9W94CdC
2g10WG,ISTZAcZX20AL>gJ4^P65(=1WK1J^?\_@5>&0Y6C11F,-HG.MS,E+b@9.&
_W89bE,N^?/.:H&B@T:;(L]e_,23P2_6V<JMW95UD\#VQFC0@)IE2E6M<#&D),4\
?U<dX>RQf..7I)Q_^?EQKbdb=\6D[-IIDg,U<9MY8/ZUH&;?PY#_e0NW9Y\Y@&]c
RASdb]HJK_HC#V;8\X>DFEHM+T-d2g;e4&f>c7QX,e5]HIPEgeA2,9dRK?d-0.F6
E(8PWN/)&ZOGZSHD9:K<((TN+CaAOLG7e<>V-/+#)D7QGZ[c24/J5bOcGd=>3Q1J
K)<VJBeY\=,Z[6aK>?#QgE#]CMKgbJ.Q;5#UU[OQKdWX#3=5g2+Uc8PdCC8^7LM=
GZU3N.BZ]+SIM6G@<=E=IP\a^W7NGA_P&&V:HK)CfU#X+STXJYD6I5[)BFG(\/>+
Q.R>Z-XQPOWJc-^X(B(H@,cM0I#dZ=1,:ER\C:O0F&8-]NP_/ODT+^CKeB<WYg#.
2g+Fca-a#]XAX4_Q-X7<Q:A^JKeA#2>3e=&/65B_MUT_,?XWY<79R]Ge@WCJS:5D
b7.KH8]Ya_12&W3.>)8<#\<Y8LEQAMU)C2_E)K&c156a@<ec_4+IWW:=69C0A2H6
NGaY7QL=[6cB95_(M<MY?69>b2F[80BGeDB&=(cNX[9e;)@?K;63IaXf#XD6ILB=
]/]S#>V+,GFR-V#2.eH)dE0.J[BJ\W)e;bJGef+GaS[V/(Oc#W:3FB2UD[&^OaYY
.,Q]^,dW_U)<>gX6Y.Q&?C.]9(F962@?^a\MM[[AFI^,G]?QXX:6O]G4./)\D3T>
CMH9c]e&=<aUZ\1e#LNFG._(e[fae5-Q_&(:.f?8J;OF_d7/TdO>JD3QPTXaV=LW
.5>:-#a,DQb\dcL1d&3>:QDMbPS\JgAR@45_c#BOfVLREb441A)e1^++#FD2EAF_
K<G>BK,[B8UY;YRZI?WJ&>NgI(ON<:,G(Q]HYNGQafR^N[(<e5/ZF;=JHTU5IUBN
=H<VQ8c:,2g)S>NS<<G:Lg\_J_5LQ8>f/[VFAGF.Y#\@C^;.FFXgTFL7L8D<5RRN
fZ>KYg^;Y/c,Z9.V@:@/[L?F^AXU+O8(NG1&LPP/g7cAF.E[67[a:HO5PEK\ZI7)
eWE9e>(f2N\EF]RM2cAC^:\6REJ6L&c&<_W:M-V]2SSZ06_[<F@gSDE<OgYa=<Xd
W/X;DD094U0Z1aSGaJ=2Of)M(bZ6VDUEN;\\\&Uf=80fR>RL-P0S,MX.Ng)adJ3.
C12fW>/A5:C<.gS@eOAg=,5D74WbD\^]gaD+P26_VgFBOc9^O3a-gde?U#2<,.FM
=QDb3GCOZace9?Sf^228NcW8P(D4^fK/Le,+-?E024?679M+Sc/ed82dSb>&\J5&
&V43PF]&2X.-0L67e3)EO:gFWf_RTU9WD^X@)PgXQ?B,+GF#DL)KG@@WB?:+T0U8
B<#\;J,e.#.0.-Z;?1-5Wd[ODa/a<,T1F5b=/U4^1ca]g9S5e^+=V&WVLP7a\CTY
X+-:+K-#T9cLI52-,1+[MW@A;/]0&3;eBCHQM_W);;IA0LIa0XG^>VQ@4022Zb_.
PM[U@,)4DL47R:7EO+cfGe;-_=A0W[Z9G2]PQ(.HWIV08R?3YbgdH2YSc0.GVOc[
^F3)2KB)GSOJIT(cOTe]a1<E=b=RVaU<SB#ABP>.LN5.+;dUBg2=HaN[Q_H,GeI-
;@I&4eJaHY(CZe@b5Ha/4YbNM;/KcR+]@f_</40[)^fZH^[)LUH=BPQ0g)SD0Z=0
,g5-(P+UU\&^B(McCM=AL]A1f)4CMdg;#UGT_NgPeVHD(Ea,AR7:M\_Q2=WT8658
)RWEX1L5UUA9T/?6N.9ZRS@#>+cPfWO)+<)6g:#.d=7I_65cHAccL(9-;eg?0[&Q
4W=IEWb],<1&CG7C6\,JQPH[Y8=L6#.0QD2KP-SF<ccZXOE.]7B_[75^Udg>eVIA
PM:KA3J9X0H<KXS;R_g9P:&5<egAAR+&SM4PIDPK;5OU<R5HY+]f\P[,5YNPMPWC
BT9fb?VgXU-Y5d-FLG#aS7(T02e<@bg.2O<&MfGQ0:/^,<KARY6W>1=T68eUg/@C
QPg7>W#&-?Rd[XS\]ASY[CLT4&MO\-V5:BAf&Ga4#P7+DR<EQ-XT6^2/4KU_B5LX
^IO4+Z^&2/\gc^J&T5g2^1H4-[fbUBDW6cNR>W((.,6ZN,^<EVUL/0<&dLD]#/7<
LS4DgX#?VI4Z,#2SR9S./(]^/NCa>a?dX?RJ6[4P[F:@d^-9TP_3HY2._YF?\WMC
#\TEI^_a;;<+=71g&T331M6WYOK0&WW/<gBU0S5Q0,&&+ICLb9FD_9H>,S7)abb^
<5J-@02@H&)G2D72=SD92S@Sb/>bX^VRUDPc-6F70Ue5Qc4N<L/D,+cO^PE(^I)#
.I0?<OB/^8ac42DXfU=cA;OAZ?eW>Ca\Z?g2Adc:1bW=VOf4GTDc[V;eac&T[b[Q
BcXc\\bC>f9G(,V.f>U>\&?e#6_II&3+RJe;416NI:K@)=,A4\Z<U)XSa?Z3KdK(
8V8HXR[.H-77F[8?Bc9XP,:Se289NGBc>:-NaOG-VUdW&2BQPGAK\[;[(7::EQ4Z
1WT^0[ODP1_4]#dg#F@UATH;Tg6JTTN>KHg/-1VAI&ASR=NNR_/@/O1#I/DEE=2;
()SZZ5D4;J73[F<8ZALgSKRYb&]^(d==cL6@bU0e3:EY^VT7#f<HVIa:FLF(3660
PgbX1e#UPQd5HAYCD\Dc7fOCZYT/4X/G5E,1XX]U)OE\@<1bDZ@<HYD.0eHE:Lf:
cK_5GQ;[-ET-ZdF#Y<NM==;4U+\,US14>?1VON2:PdQ+=1CGQ/O4//W9+.dJ>WP6
e?Vg(Re+E9^=?XaCNPO?;b3FLGA.U<fG9E6Kef.=VbReWa\g[&2^8aS)KfQLbXg)
8_/8Z:dGA]E^fd?[g+RY53/Kc<48>E/?e\#5c+.ZY<43@@4LH.&O1g.Ue;>AU31Y
4/gN5gU=R_aaXQULUI87d(JKNCIdI&bB:Pb\_3Y9I(4ZG]/KDTR:V.3I:-G6FSJ@
BWS\f,S[G_QSUD]dHL:5C6C9-L</9U7LTfJEM2Va3M[4#Y3E&P,&ecKZ0HJ-7_/d
0fNI8Y7OdeaRJINPW@2EQ^H8G>G^1g[(;C2:dFB0cJ;bJ92+3M4b99f3RaH4^VXU
(Ra[JYGc?=W0+Eca79)XTTgH2O6R6dfOEW.S2gMH\9=CW[1.IbE[2a,2YPQGN/0N
JQ8^LafX058P+#6QIREWO>_82S7<A;EA<I_&VON?+e8<+3#b>,d\]0GH^CeVLSAS
QB]PWP8Pd7514E?bI#;JF<A6^&)8@E9TBGWE(?X.^6KME6dKN0V^9^.6[@:.DEC#
+FIK\:NV>3cS/:eLDYa3eGX>M(N@)B)4JC6G4D:AYLL^g6ggNZd5QWf21dN+F<-+
b36&bdP4;?O(6CI7E5:&K;8..U<dAAZU+@-e[^]4d91<WTd-;0YLTVX@THQ9R.:N
7#)9)Tc^JgKEK_\(X&aKM\8>d&UG=.NZHaDR+G^+fFWGW\aN-;^L0MSLGCY.4g#3
]G_D@a(]\H4:7C,FB0\R1;I\g\ZK=C95H_;)IgK6FQcM4[3)VTVESG)e?Sf]QdJQ
&4Yg,M(aTQf?d8PE,MC+EcT-QDYA;\^.bW<+gOL\9;IK5P^9,.&.82/C.[Y=;BC;
g86TMb>XTeDJ<=)4R/#?O)5HRF<AP/XXF[]7)B.-WL;L7EfWBOQ+]:-(=6efHgI6
V(bEP^H<e7F69V@;=8,\;]GT/5#8TPL;8+X&eID6BKgdZ:g)D<5:aWeTDK,(O@@9
>@#f_PeG8W?^W,;2S?;BdBY@C=C#3D.IGeaMb+JfW1JQ)7gS_:Q2;I)U\=A)CHDT
aPc/RB7;:>-=;(#KeMg2E1\<d-T?f>#1GV:8)Y.bfLJ<#K?]N]7ZUe93?U92G7L5
\e3T#)>DBa=1=e1U)9>].dING]A?(B(a5&a]<GSS/Q+NVL-f5@KV1XeS#UE;-AK\
@STAAT;b9#=0NEOGWaBT]U,2K8DH1QK_Z6+CG]e_W1JL>X[+S?fVD:VIQ/d\8)0F
g=X(.6fS#LLN8#3FHLZO>If9+UV8d7X4O[XeMV+W,Z63C-SJG#+8YMV/@_-4g6/L
@Y60M_/IFbLBS_+@e:Nf5;BWeT)G=/C=XX>T5(:EA[47[cW]dKH7KB4YHe+Ua#1M
_c^d8,_F8,<X<+ZHRZJe,dfI1>QD&f(]K55&X-ZE5GGAS1=K]aJ)2)EQ[98]H/7N
+dH3J3WfPfc)M>0B[V,9DCL@Wc=XGgZJ\JD_eUCQLNAbL/EZ^#_\3d)/.BDYF.03
L3U0<O.?6LR]LRPV(G3K+DJW<5_aMW;XGS]-W+/:^<+6TRA6^b.)fUWRWD1KJB3G
daeTMfTY2.cH&J=Mfd<Y0NL3:D8acNA.N+<UB=XPZN[1>>>f)-6a&S>XcSS+^(#O
4GJNC2AS1)CD&SAT4g8G_Y,T8622cU6-FdY\7\;=P0KN6924R]TXc9444WIW?MVU
62Vaf#aQaeIce<c;;ACW0KZAB,?->Q)47LU]d@(;RGC6^fcE?YOPVbC6K&_H?TQ6
.3<&f+<^_H52E=49&-)(f)f+8?NDFfe&XIB@]_SZV\(R0)=S?LRY[b=d+Od@bR^K
a#\d_H-\_Q=K,PKK0T1#=E/K(f7ULTee=U+A^D37ZR5R.TALDag078R?7^VLb/15
QRd,^9RY28IZ[.YA]AT=)C3CH.V/VKP0;<[IIYbbKLA]STNMe5FD/e]#XFJ<Vg;R
(7>STPGQ,(^aA/+?I1=J<g#VW)/HL[)L[8bC<&:BdQd,=<NMR..b1PL@7aFb?I#f
VF6Q=_/0Y3\5,NP;4-9]:(4aT@-=RcV:JA<)T#,@W@9T\^Mb5d/;d0/7?BML7H0S
G/HNJ0K?&c(GaaET#R<YWSW_X)DN@Gf)Ga0T#d)4^3Mb9[/(<BO[3[[PZCf4f.=7
=KCIR<PWI;M+73S@cV3Z2?(a=Y,E5a<?Je>NdGE)QOa[<T##bT-F4O8[S5+(QZXb
5H6^]YLc\5>SZ1KN/1N<;B@_\9BW=9C]/92993Ed4Lc2,XOa>XQ.bK(&c28F?18A
7_V9fT^4#L/[JbN-P?O7?Dd(?8G6N0+Eg=cRFB=]dOQ9+;G4Kbe>.Z]c?V;0>]3L
=)FK3(>DJXQ:c?#2H1b9eN=#K)00:2#A>WPS;,^g)42:4ScZ?>4L.2]\&GQ[N<ef
@;7MSM]9,6_UR_/O]_&/)&#QR[;W@L.GFN]_\]820YG=0\EK0ZOUR(Pg3S/[JeU[
(>aKE]-_a\4M/F&LWX?6JOd</;>NYaDdYF_VdV0-\(e7,:6]3H7Z=BJ-0>-V<2dH
0TS2J.TM8/Rb9O-cd-;D-<-=UQaTHLLV3e_S&:Q[H0H=U^G6YR(V0=Ed2(5gaT7c
)6(DC@bLdJ/d>=OAd;U:8b>[Y>-+eOSAASM.?S+ZX<)GfJ(@D(JK4:<_@].AJ\J+
3Lf#6]UFOX]#[Haa8,H<;_cdT,3B,+>Cd6UO+?=QAZD=H/3=:-dI:.NaP,8/)>[T
KTe]A^3\00/R[,EfN:e#C#&<-#XcQ,N10+NcXK4WH(f@+-H_G389^cH\O2Fc_06J
2:@9g+a(^0B5L_B85>CcD#gc<)#aTN:2>8:)5@/FM@7eWL8NAVDD3QEQD0K.D:DA
=cbdDN(.##IU@X_D8<:<_Y)<5>KYS]0EUVcXe/>GO^fc>>6Hd)K=?\I,=.IX_AS&
^?+17B7O=Ie(;2]AFI&GXO(#[)K?(EZSH(>6((,HQS6W;K)e^@=cDFC+)X8ACGFH
[H)<:A\:=^75>/2\5T)UHBF3F0F&DSE9W9U_#L<d</AeOH-:;Kb5.+a7XFgG><eJ
ZbCfJ\OKVLJ?M_A1HCeI2BaB,KM)c24E>YXV?O(UC6)R:&2=?7DVGWYdM3VOaZXO
B9W&G_ZM2Jb[MH4gE09-H/bg@EgFJ>:AUF@[C\Q??57D2GPK]J+VRY-MAc;ZH^XU
41Agf1D&=^JT4W3:=eY;Y]<c/ZY822e\;XCagG@/XWF-A.-XA@93Te2CJ^OW@D,9
KC2+cFbDQXGH]KagSEFNM5CUfHb0EM>J&f^)LT.U49cI,NJ223#E-(H]8ZfW)Z.O
B3aH>YW+Z0ee2F-c=.S;-^RJgDffcT^eMf5:Z#C1&^Zb@YgK/1=AF(BbF[G]c9Ic
J5\D<9?\S6E9e#I0-7OE)MW,S#@b/FJ4dGDN^_DCZNLN=^A3>:[68SM>=H7)[GZM
J]Y0A4J:e.GSOG=91C-V5b</9@c(<U22SX3]RB3[-(7)XX,D.AR;8&:9_,DaKM.0
09P@_\X5LC4J2\T8/0FA?HQMREXeS4FNJ5e:S,+H>\OK00PQG56VcPV:3cVT22bW
]N(4^?MB:\8eR546.eL:BNYITdX4L[^4/VbNTI<ZZVg,1<ePZC\6B[07f:]ZV(E<
5RUL=.XYec/G-P0WZF]D[54R_S#P#=78f6F^TN.EN=EP@7E.<U71#&TfC_W1c42X
/K4ZDBaL&F+MUAG@_RE_UBSd+5SD#ZW86b=fSId6E37,E&A4A_#VN/(Og=^OLb/;
HOF]^JHG_QdOU9)NSY4A.:8GZg<?1X,D5gaH:(>9><C:U]K(gf(8?G:CZUWUW,+2
+KI@J,7-c><5GB,-D=XgV^BI9\:acST&AHL<8R_-^c5B_dPHPdbYWc(4#Cf&A,3K
\;O?7B(73M/O&_EQ]R61.0H]6Z#-9\g5T8&8JK^N,.B:eJ66Q.U(C9FA&874ZQGU
_AXBBf\KJO5#c883##9&^GJ(F^+,XN1Ja4DX@Z9W_&We13J5^A6QKH#-CX,.HLRY
N]^G=NLV3#3JK?WO=XF-SWNDUSNe3C(RV6NZX/Cgb[f\4c,dNWVf\D]H.^gZX?T#
SB-LJUg/9A5W-K5UK.GM:e,:73V5bdC2WR[7HBWG.XVX:Y[=L(B>7.)RZ:;J,A1\
UVAWGB2cR2gQ-VW>&;@TE<BbCW=9J2)]G8DEC^_fe-9FA4B9e]KLL0:XAfST<[M<
S._791J59-FRg]I<CQ@fHGR-:8SQDR@.Yg9XW[g8T7/7Q^I)Y)JF_MfNRHJ>MYS.
5O[.(Kc9G>[6C_?eBU(0Z2I@_g?)XB_(Q?&G<E#DQL>J/+eV4;A),U4EK\AKO-+Q
&AVHGZd2T#dZ,\PVH;_Ed=65WLEe86YS[7<JKce=N2VIM:M[FKXECDVFQVc<0+]a
[>c@,bd)((;Xf]7)6=_:.5>-,I8P[Ia+cg^b(6eY-:(3BVCP^0M+b[B)CKI18dR1
UK3M4B3&\[/>+2\6eEZ6Dc?Kc;Ie.A5IgITa>/+GF^GS4Z&2INK9UPJ&HZQ8aTZg
V,60Q6\[7eWB+_J+.T6f]E#HEVaC7>-#H3#5M=GS#eBEMTID>=&/b)>OCQ?[,:KA
^_5#BH-;ULZY6<8--13OJMNTQV=YBVe6C:O\T(\(8DE+K=U:.U].1-Jc#N,B@8L(
@X&1H;SO&RAO#NSYK.5)X2LfT<7GdS]CXd)Sb_7^Me4B>I.g&F<UId&@?36@9+73
ILTY?W2S?;B#5J.Z63O5CKB0+UXeeeT;_abYZ=.:,RRX&fYJ.XAg:Z9=/#I3M8De
T=]W<D@B9QMO78_d2&I/5XY\&<>YCUVYMWZ9Q4&0e>OL(8X&F):?2/NeC5A_GO\U
,+Y.#Ya-P<],QbPG81/Re7fZN&Yg0BSP>C\>65(NPT/W6RIW>F2Fe.RCJ\GO1^=R
@c>P(/d[e[H(eCUJLAb?cQ<[E)8(d0;+U/_,2W5<7f4>9+#97cEfB\@3V4.4:)2S
Y5JDZYE>Ic7+&HOIC)8LRLK24#4UV&,;VL=MMcR]d;QUVY&;/EO?YFD1,_ggG_&K
M)S_KU=H&FDHMPE)U)@6CYJ,RgcK3?5\KBRMD@</gNFWRW&\f47Q-2;Rg@-+U+^A
)11Ec4aL+,,<TPfgZV@H<2cZ]f0JGPWMF(E([.^HPU5^)g0W241cE]J>VHMG_TO3
MPSPAU,CPe_B0+F\I8eYc<T]O[cQaOXHe#g3H+N6;Q&AH++c.C9S9MV-/I,;]IL6
XD2N<L#/#YE&K6a3PdOaSUW<9U.6=a,@B=3YAZ2c;3a#JZO.>eE;1^;ZX,.C\?;[
NS\8O@FZSKP@9ReZ9bH0><cFAK^_6aJ)MO[=QIJbTf80SgQFcF8HfT@<VJ#1_&2H
-Yf4J\YVEG:SG7,?W?e&T1[.LJ5F^+&,:PYT^ZZW\e(Ocg#0[H>12_?6>7WO;&@6
7^J_:V-B00H]SNd,TLBO?MI&ggO\dWP=EG8M1]D^Ad_VFM9GYN7d(5((ML^:=c#?
:MX;99Q?K_5X4L:Xd@S725/VT<R6>]U[78(&D+82R6P4,CO.I(aOK_8D<\dO-7=1
@g80L:@A@b5V@a-R38cZ#E_;8N=K.8(QU7bgB5WEK_P(8.f.,bJ[B?=)>412b.2)
XZ?FPV>TB2:04LBERL2QVW&d>eB9>R7S[:a,IJF^[-@G-_Dd^bF-0fXeJ2IeJW:6
cJ-bEF+6M(.O(O:I+?28(</GJe4a3GBI,IT/HNJU[:-d[QAcG7Ycb/-1>AYeZ/2N
2cON\^@48ZHN3cYY_K,&BMH&O?He4IILHNIg^?OW>fV?8Pd]=4_Q:UL=bY^[0-B9
<E9I;3;6K14R=&^_\-4&;88IH+S-2>^[LT1M]4N^X04219a>>G#OL\\KgV_C87SX
1f07:[X\]BLa:fE)Q)2#]=-8MYYeL]<^HO=R[0@:(77\H</J//U4H55Lg16\>J&e
ZZT#0aQFQQ9@VDTddH[KIgP:T2WK\/LA0HTRYY5JT?TV]<6UP&\E-#E:a..(d9^D
<[45UM&V6/cMRIcX0.S>H9]KbKQE:B8WF+,YLeA\cQ>?fDUD1JKDRMAGRd>M4^EP
2cE9#1+>eA;O\FGJ,]L#-e2+da>^.eJg-S;(KV#F[TLSTS):bX6CS.RB37gHG+M:
QB[HgAcC<f:YeR&Gef<f9;XDKHEdKS4;+[EdGXA&8g[D:eRHFZ\+_1C_:1ZC@;YA
KZ4JcJ2GdE5PEHV0>FLU[fMC[4-?]ea[P?M^cSZW_PJZMEHG=30EEAN^@bC.BVMM
#JU1VFK3CWHA\fAQ7:a916Z4=,9RL^,B<C<.I6(ZQ4L8P&7P]]^LQM73;QWGf_d<
X+WEb\<)S-@1e_]JW]I7MUHX\7\[R+9371Z,_ZUN+H__+(gC#Wf6.SMXPf\Mc[Z#
4f8(5CQO>FH<M-7f<_LXYFVaMA]9])fE]F6dZ@O-A^fc&CJ4:(+N2VH3VYLB@+KG
W51A0:XIb;UY4E8\:][X/_S&-F9#591;dc;:?>QW5Rd3>FN\_(g6cQ#XNdY]=H(^
76[+P8)4T6H8>f]W^eR#FN5YHC(E;HPUPOgR3T(]eB@fHSH0bV9,Sf&#X(^4=4G7
(<&.[<De,@1e?N&\+T8ZGV>_LHTT5^1SbI+OLT:^Xg&&1//D\NJ191geG05A]X=2
-Q?V69cM59>@4/0fA60.<XCPGNg-QbAY]T82TYX35(KPX2(E/P0g:/;K(@VQb)(A
,DH_XQ;^YeK3,BRd9?N)DA4S#<;5&NZEL#EB:?W3^63Tge)/[<VZ/ee.D@eff=5e
cFMSK9.6(P=P.)ebAG+ES6^3c5bF_Y&^YQFWVab&^:N-4efg:@B]W>^_/:ZeJW)Y
Z0F)J4gM3S6BACBALI3RU=?QP9;/g\Ra^46CNYVR(8YIPG,[4(ILEOVIJ0#KP@>d
aKH1[QI3;W/?CBeK^01OVbWG/,fA^Y<C]\C>F_G[(^C5TM-dT/N04CJQ:VC=e3&7
^/9S]Rc_52,:YcC[3)C+CB)XJ\T^f3Pg83d]\.L.>dAa#caOW-MS/g_W_2G^9#gI
[5ZDRM.ODVR.2FbfE;,e7.-9G+&>9b;0CfX?]6_5)Z?4b)(C;UW6&DJ&f,\cCX]g
Y5LOQJNZ,J6F/J7-7X7cA;KMAA373Eg+C+,9d,A36-7-+CdaO[I.N/4D0f32HGWd
>,3C82.02==OQD1BJ3_\D&IFNY(NI,7dOM8OC=(dPROS/>.e\;SSL7N;_dYXH.UA
4?0W()HECQ1^T(,PJ@>B5e>+ZUb3bT+;.QcDecD4-[#W?]ND@<g2BOEVgACReU1K
TR=aBQ44#(87+bVCDO5M321(?N^.+6#XU#NTK3=15=H[R)fWD;MKU+;C3668\B9_
LaMG2Zda-B<SBd6=GD=4Ma,;S41=4YED@U9.EF@e:<FDVDcQHKVFHb-2<96N.OTI
.<8a1BG2FMFF9K2W)f#FDceN3_))MKf65^Q65B:J<I?XIPTVGM-Bg.eMVTW7SR+)
,OS7?W8P?e[I&ZQMQ0Z@(4Y.Cf>.2@D)#U14[X=.f<U_\MNfKN.L]S6/4]=@D;+G
/(Tg&?G+\Y,@H]-Y#SK7CUc\[/:G+/)0&gKY7:D/(Z>;DE>#gJGIQa,dPWFU.&FU
0]MP=M9Y=g81ALWK?8U@1b3P<(&B\+Q=Z@^L0D+S<G45K;+d):L?VQ+58J]U1dO-
[;F?0F&3&@b29FVPSK7GVM7D^YL.)CaD;@bYZO5/]7S@^\_,AHMe6>6<+Rb^2S<O
+48g\1[.H6g\=VM:^J8WM>50):\I3R7#7AU_=WR#DQg_#0I=6f/(C_N9HQTDP)81
Ec/R<Xe;FTXa]JU?LVNC]dMU0,OP;UbOGINRW3ZD[3[3CW,1/.6P6f,Gbc+Oe>S6
F7)875?@UZDFXZ#?HaY-JEK4+eXS@V&H4\DN?59I>]##aI+0JI1eJ+;7@1ONeZ)_
A/^6fQ&6I^MY,]\(db\OR]X(59;9&GC//#L8U\Ub\A(F-N4N8)g5?W84LWdd^O-D
X@_RLM5#3UCBT8T=g-+#/7I#PD3=7K8K=/9\E6/AK2gZ2\\W6J/UAf&Q1PA]RIMG
fC4WOY)-47WfR3f#4LJ3WG3@-#6Y:bFf9cDSNC_7R-3RY4f)^7^O6PUP:=YI4AD-
[HOK/cSI]W0@9@:4M1/GV.,?eC6K258]+#Y?OJ/gF)&KeRF(S#1aVN;JK@5UK^=d
VBD.1LGKZQX9M_=:&JJTK5@I22Y;eKb:WFYQ[bB:JQ?cKKg/;6MX[;gO#SO\S7O_
cBeXZ[A4EEN3DK([Gb6eWLcV+7\QP=eW_eBOFPYeWDIHPN=K)Z&(K=CYPAQd0bcF
3fQ)[@_a<F)[]:R^H+S?fd_cD>LH3223@YC\4I2#X<#;e#U28I/P6NIbNXC:?a]4
.Y9+T#\,=\d+c?OBY<V?IH1^Z>+LaZ[IU:R1OCR@;Df3A)3WQJU2Y/E8ICZLUg=V
>N4BA<XROK(;>(AB0,.NN2?#2KZfJN._[&)g/<>b9G_Q/gIegXPX[GN/-E1BE6-T
Z0H0:S4Ef1(F3R7Rd09a)UPAQa-7/f=IIcF19f[5;[a<)-e&/b89H.YII-N.NO7@
Xd_MWcUZCBeReJQEbQ34B?IG^[1M_SQ2+L3&)YE_COQBbJ\V0c52KX^GX-AdD\D]
;4].6ODCf82Q<>5\IGaX33e:WJEbgga\H2TG@&8+>Sf15OMcMfCY:/-)aeVP5(WM
.H_PgQWJ]<=O;+N\(eU85S5[YKS3N2L@b]Q6b6F3X,:-ZFWJP\]\3S>O#AT@[dI-
1Z^7P25-_<8FeKRBR0P37+;@OHN-/-(T_I-DHddc+FF87JH4aPF7=A01A1>ZNf>U
VEe9cCR?[?,43CF/a(71T-A_(&:9c2PGVbD0GG=_&c&=..&d0f32:3_ZO[M@bC0:
#CS6bg@HUF]DQ7d-@_7MKWVWK7V&)8V5.:1c<\OY#g@&/>B[8JL]+?;1=gPULbN/
,BaZ5b@9I<bGU22-]ESJ6+JP^N>N<&?-[1ZLc+<O?9SOF=ZU]&#N@Tb,<;gHU?#Z
?UH]c:Q31MK1fOD0XPB=0_O+MGOZdD)H6R?&R@.5ca9>:^WS.<M]&Z#&[C^T]:>Q
;dB5NVLSDWNcgNHfRFeG4MRY2U-8\@LbIT?ZdA1->U@/9MFgJR]4.9g3<1.Nb=&V
E)J8@?@0WH79\Ff3KGB&V9\SeT6B[WT9XCB_H;;SNfCdV.f02SA:3]_SW\/NFYS+
-[Pg<VUbV\^4UU332F.cZ5K7M3598_d>T)FV\_5SF>#&4Z^]DQP((=ea_JSR;HLD
Ob).+Q>Ie3)Q0\VBAa6W=-dTOb=5eUPFY<Ye>bVLbYYW^V3U_0^:D2[,,Bd<0[9]
?O6;:+(:DR>SLXV0ZB41FBDU>Z)3/H.(/d+@^5>Y^_6J;1:?-N&/_>.E+S\<bbHN
:B^cZ32f-:e<RBUDP^.<Q+FJTKDBJ\=>6R<R6B0^Q/Q=9GGZ_4-a?55gAc_gaLG/
AV]dYV<0/L:.ULf<9D(L)cT]@>X[MXf\-5f+8H7PH1.1U/cSJ.1JEADFVU@J43b.
0,-GAZS,>Ye=R:,R4PH@.(\a8;;Z)6^?(dFJg\+Z8g=2PUM>[Qf[cB86R,TE>MF:
/3LC_T9Y-XS:X-K1EOA3fbAL1<f3Z&,d-c((Z.5b;_3dfR(9P<Sc4c7g7SH?0gKI
JIa+GXbP;VBA]5DLL1\e18)gcbJ-c,M:SX,@D[Vcf;/B.a2PGZ#a0XZ<4JQ5JW<X
^U\,b8\F0IQ+5KWRdRM.1_g4+R^JeUK&aB-f;4NbH;EMZ/VH)V0^@7a:UaVfV>-.
WC5?=X@ABA.0F3Wa?JdT3B,3d4Z.?M.SB4;()<V/EPbW-4PAY#&5,.I-cgf46S_Y
RPZX/2]JVBU@XZP.5:CZ<MY-Y,M][L\#RWB(<WIPe8Z8MTg9S+gUU[17;Ca69]bP
L8C5G/V5T)GRcN)IG9GJVGU5(RL#9&5,#.OO#K8U.919O5JB&f3]>WN;ae?T29B<
c_:75S\-eb-NCSNAAO8#[#R(3aT1_ES>SU1DG]\[#@D=Kg0Lf4>\4:dg++_-V,.N
PTA\,&H5b)^<;\.GR&X>TBg7+<9E9375Ld.>OCN1:3T;;M@9Y0B[V-V)H[O>1)He
,NdSWIZJ&0cOF1[a_6beQ_9G[(RSO_\:D_dE;9:B>P<BadHQ:H8#/YY))3)f/>K.
]5O#CO,#^/@_+)bc^32>G<e]O=@FP?)8S5#BdHB@VC:MS0Y^.)2;3dN&36@3g:c(
DP@-[Z+2(G4-LAI]P14L=H>A>6:Q0;D_=d(^M2^cWJN^P;2EJ@&ECG\eZ86&b,>:
3X?EB5Vc(@K/>KZ)+;K^T#g45UV<_)Q8A6.d59J9BKH6-PWG?6?;<IP2ZE)I\BB;
LMOb4QY@A\HM/<X<KY9aBQAVM_6JBYgURc57)N&R\NWWPMJ2C>PE->aH_?L?\I[#
YPHF>X.[XRc4M/@7HZJ7LD#f)7,GS&X;IP(ZJ>E,CdUXMVMcf.Y67N.O/7aO2Ag1
dBe&2dCURJ98IeP+eI;b0Re(P^-B)^Qd70@Gc5^^,JH0@=b?Y1A9,\#T]@Zg)HZ=
.::>A-C4UD[NEHN5<,LK.\aU(]6I>C^>:]CSMeJ22BH1QPAg9^DKZ?##+JMe@VC:
@Y5/<HWB4I2X#1fRX?7L6,F2H;fND+8KK(/[>2VT_L@UfS,E32(WXTB1W-Z2E>d5
b8Ad(44.9PW].]IBT=G(R-aa#V.,-[g(LJEKRMg3eNd^0gM(O7D.9Dg5KW/A(.+K
fBe,Z6[ga,D9QK.IPB#Y)D/E47H-5<XE^G0@1c4:T3WcY_?L.H1H=T+cVE3HH&(K
XU0]cPS1VW8T9JKd6/E)?]@aOE8QHD\WXaGg+bP.<XPA-&1490M2Cg]<P;e<,KJH
MQJg0VR:eT<<5#WLXfTP+RBJ3[6D;A.3Q\VQPWY#MAP1A+gJIR?=4e33d7aB0\]d
I,)Vaf4<\2-PY5=H0_LME6:?EWYfAQ5;\d,b5d]^&f/<gb(8S/@@3:<;D,5c6-.=
0D]3UD.<S8GK/TeY47[891HR&Xc[7VdIFa1YR#eA<g:3YX&A0<aK#(83TNIYFPbd
F99&)-8C6-e#GZ48\_>:B/2cdTGeOBDc_)S]&fMO\<a?1WKM&/=V5YI;cC0<N.O:
VbO>7O9&<6(#@^?PPY1[W.3@-0bRO@5.LAH)&NG6_-Y@^T\fD0=)/?[N6(\CUbQA
51DU+M4Gf2OX&@JS2DHbHa6NaOf[FJ&[N52R@B\[BC<8Ug/(<=YFT=UD=UK&6SDY
:\_^FK1Wf/.B>^PX,8EB1acJ[GJYIMVH,Z4K:e(XM<IMdEEc7.]FWY(_cN^)KD<)
Z_K8(KS&Y]NK@)Qf/>M&12?=VDcd4#M476#HQd4PXLRBB-)[<D_,^gTP<=72,9]a
#.K:LIH7BBdK^C9?/&5IF;HJ@(/S/e8cMG/)AbW/:<Y;f:0M8&+#K\LOgGJT<&C&
A/AA^/Ec)T#a_2OEP082_/EOZId6bTbd,dCN6WB;?>C\T23C[FYYLL.VK=L054KZ
cK4[6X^)IU&D5R<(A)4b6-dEd(bXR0\(;&0d1<5d#2PDKJcBIN)(MRNMSHSSJ_.N
/TH:\<0\QUcRF2/G==<R>Z0FI[-VGE3DFML,CXCFSU_.YU+aK_Z,0J&J?RJ(fCJg
13XHO(VWea>HMb=g>\Od.bYMNV)gDCK;f\a,QJ0H624&DI].]Wd;71+1G>HP_9BK
#0P.?LISB2be1&,de]T09f?(_-APJ@.CA(CKZ_;/S^ZG-c-QGfRS1AHQJXbMP+^1
M3LEX1Q>LDCg+_B^b:.I#6++>Y.3I_)LCceNYKBW(/((,4E?YbFUJD&Z?<M0fZ_H
_=6\VU^ZDe;f]D97gV/5P9NX]>MW,Y^,YRCAN-7D=.6[?_aaKDXE(4+BRK4ZD)48
53W#7fd9PaY?;W^[=I[\YRG_TJ9XISf:WLQX(B2g6^.W\A9W#ScaCeUO,EK4,QSe
&GE]f26HB#8fJ7W#Faa2:+CXeT64P=g@K-.H=2.:FZJ/0;#AQ&bG_gP#2T,4;01W
XgKSdU5G_@J:URHW=aC\a]UAR+<Z+;F=E(X5dV\?RU0a[Q\K0g,WO&/R[T&9K+(G
5A)N3AT+^&S09,R[a8+@4,6>Kf^d(^H(<Q-NE8L-TE]PLA-E8Ng(8L@\,C3a?\b+
IaG#fRCD]3?JE>TT&#8f&WL,J<d2_<c-S]X2PbX_]Ub+TY-I@3>gBW2Z)(&JIGc.
I<fFZ2;5.#F<H3eY)UdgSWcAFe<?b2L,+BgE]bdWX3M,@L41?R.&Of@63O5@G6)C
:EI6:AWLL#2a03/;]9X@bc6O(A>YIcFXY3^BD?D(c;242P9d>5RIL=Z(b[#.+K]\
0MW(+Q36#8-QBbMd9_DZ/+&]&TH9B4A/M,0ABf=?67MZ-XJOY88X1QN^gH8E?]aT
_DT1Oeg-\Xf,6^?U(JRL;M<f)@Z4XP7^^0:L^bU2)IAPHg6O_H>:+QWG58Fad(@)
L;@(U9cA5/fZGCI&[,bNZ=7cb?UAX0@aG5SC_CYS^,<@XY.(B9/a+YA+a]1<M?D[
HF#BP8,&D\)W5IGC75F2Sb[(5\Kf6.6d-Wb]Q[U]XX&eD</>(4eRL-<QFbME]^:V
/Sc>,5TBC251b6/5WI&G#I=FE+fEc>X1[6cUKKQ6bOS-1Q#O_++\,I870f#4AZ]D
?MagK6ZNb@1gDZ[>?#,9E2?J^a(B)I](,a83fGcKKR?ZCE@KI9_/)53-:g>G\f@L
^(Y^3.),aHWVRB:Y.K2^1)02(4Y)9A0:8:(]^>V<;S_GCQ,5=UJeB3R+(7JB>H<C
4D[fYRJA=@2(e/#^feeP6U9<VL<dgI-D66P?ZBD1Y9Y/\.@)K3@Qa)@\88Y<O_[T
HKOc?eRaF<D\-.dIOg20bJ/.J1+\H:N]U[SE>/1a(T]/B2-O[QD/R\F-7\651g8)
7YK-)I3N;8a-X&33P0a[@24@3]SgZ/N>BZ;]/F-[G9N&5XGW)MAXE#:=Kg3:4+62
]RI.Tc+EJIOdWN)]CC:BC+BP#B(-=(/7:B]W,R)b61[K\f]@fO+ELA>J(SI(B&MN
K1YTgG.R>+VN^DHD3VDCKb.&gN#L\eR1BJ66_X3T5@8Ba89T,4<3Ea,A2.=JKS2J
OX_M:fG-^d0)U#=H;=G4RCY.#,EN:V@:)6CcS&cW(7E=S?_cR(U^=c=6A&ZH])C5
6Z#2X_cV&-])bS9J1732A[[SW+GCHAC-YPR1Y)49bEUY1:H#P8bbP>3NBZA(+XUG
1RFW_6RAGP(@:6U,DEF;fD\a(H2[Af)D0XTFS^?TXCRVKG=.>ZT8PL+Y,@H305J[
,YJ=A\1Ac+J&3^0#cE<OSJ9-fSYF)5fHC/09S1VU0-DO5E.T:TVVSQIAO3F\>34.
6Pc-Z0[:#YR:V<<EaVR80DR49/7<e@7fYCeN0P1c>Ma[BC+<^LQW(V-A-598VXW\
2W@JKgWUaZePII1#?19D2IB?R5ZZb(Vc+EMW(9=EYJW<)Z)(M>8N[8X>;ag1X-5e
EGA/-M(?^UIQPC3:?MHH?,c/R&SW<BF)EZW;B3C=)=]/8+HJK43YgO16N71S>a-6
NM2+&-SN?02ZDN<?O?X7,a6KF>8aP1[@@SDce)/AO;Sa(PX8IR[#EDL/#11&K5--
H>JL:/-&a-&W[P+5S:Tg,\._U15K9aP^=[&2fVE?,RYQ1(Z.,-3:)RgRWAEA?Z74
KS^=EB^6IP:^5H0Ab7&E&#=6[F,W_52UgG3^5L2&K5S0@]W@O3F623\ef2K?@84[
:,28fY:U7?+b^RT;\L9Vd,@2S&=C:>]0B>U2E;6;&P4a@WNTQYM<SKYV]9I&)XLY
7.&0BFI,JTO#\,@<b],+CK,(<W.>@.f8gW4I:fN/_a7L.&LH-#fZe[cC?<#e#UW7
gBWZRS=P/6R:;1S=5E_/:8I^J7]]N5P?@5/0W21,8@WHac6V@ZZ]fg+QNWX5T)R;
=8Y.J=UHP/I\MX/?9g2EK<a[,FZ(^0>KGdM9&QBKeN.EF1(=^S+[2UOPL@KeXRJU
:\)UCPZ]]C:=f9\-WG,5._2R3S)ANU2^QB/U9NR5Q(VUf(_OPR-(b,NDU\P3&NIT
5cIK+]X<Y4ab2^@b<PU9=.G7e\Z1D(@DN^Z0Q3J)_EPJLLOHFR#;JKO6OeVODF(f
V:31E_J?(I_YUNOO<((Q1)TAb<G7c:T1Ye[M@(,;+8-/;f#O+O/N\9QWBEBANQ8W
P+=b.XRbg#dHI&Z-bURDNBO=40b:F61UQSCF:cE7CO[.OEIC[?UM5YRN#7/OIA<(
/a1D3LLTA-Q=LCCW2b[ZO&<+-aDJ5cbNg/V<HVP;;F@?1UB3KYRIIcUJ6??F6V^?
C4ZGC7aGJJ.S@\3MI^PG.WY>6XDdfeP=bD<:KCOMZ0_7RLPc8>7CYZOF.,_c39fX
G\_K55:6ED>6+dX/M\+-U8<6\+(T\4P7YUc.bZO=:<3BaegY[gAXHg^NM,)f>SEg
Df^b4T&LIM9cJ8)Y&?B]NcD^.770@[)Dc>RGHHY4I_+V/QCc4RfY4ZD6#Wf=B+39
Ecb>c\@J_.U4Y4C+7PHUg;:+S@CY89Ne:&,F#&c2b;f&=[0gP4SX1Gc&CA5V4X>S
K7+[1+aQ1BW8J&f9Ycd,2Gg\,XW=)+R-.IXJ),BGGa0B3.>;=SMaGP?Db/(d,?Sc
^=LP2:;4I#I/e2B.+B;&,4>>:GXMD6(<D(>gd86@TcEIM-=_W,Ve2E^G]@a=F2S=
bDY3Z5+_/O\?7b)=5[W>eMT7+1KeE8Y.<7N_I<^G?E<WNJg7L4CFQ@X61>=C07a7
PY@bO2fg+K^+;(5NR,SbfDdRCNb>F&3\:PVV=d,<d\aY-L,ed5MMF2\8Z6#V[IY.
77a(2R0GS9@RH:Mg7A)WJO^aI\K-NcS5QQ@5RN@3KCTQg<6+BfN8[b&a\70L]HKK
MH-4G?cI94<+ZRS:_&K6Xg:c>H8@dbFF1GfQ^^7L7N-bSGB6K/M3b.E[92@e[Va7
#=.KXE+]DfLIg4WR&?E=L3L\2)P)J4KC1<\9;bbC[I:OIJO[30X-E,6S;JFL,Q7;
0X:RXUN7C+QS]W9e?)J=-g0#Y>,@egW:E+<>>Z)DL@d_geJb/FY9g?OCe,:6R5Hg
_M32@?5V/[@E8Ea.Dc\=KTGUG@PCFN@\@_?(M;g/(6-0>&C@(2&IZ99TGFX+bbB<
QU2&IE0,5SZHR5)@]7e1eKMW8HD]+Z94eX73,R>#gID-V?RaJTK2>1>=7B\HU<]C
eE;cc&7SHc(M4DU):V3O;Q)3bQ^cgRM<-PTJ-DBOWS_,0d\&+<+_2E7.eCe,DJAe
3-8LeLafGN3=WUcfGDIZF.T/)CCgDa:fg7O?-2La@#,e@6+dMV03g0=PP#UMLRE^
dQRcOGRJ\-#W>7VUG@[]EaAc6\Ie.C_aK\:-4GW=>&H(+f^).;d3NPT4],OF\Y1T
#YTf-O&d)UgHJBP=6BJXKX=(dV:aAGE0M.AV.6N.-(=?(N28)#7Z#YFJGgbX<#d&
gC6EY/V/K\-0:_6;,#M:1A2Ge038XdL[0>2]^Ie+5@L1FE;;A.QE&-K^5gF.>_A+
&^LdGT^e0;/GBOEW#\EBgSe:eF&KL607_K^[d7;7>?G,TOFF6+4^+bP:T&BFS4be
J^e8P7BXFM:?^P\Q9N/5M07P)Wde#<R,;T=2_Le8^-EUU]90M4Nf,5\W#V_b0A-P
-2VAD8E4>[;KK)YbKG3ONE,^(<R9]V7/cDQ(7)K@F7F.U^^2>G_&==CLKI4NQ+ZO
2:,&1)-d+ABZ\TQY.3&9<O+D7?d+BT+Q6G39\_V/-F]PUSZNP=R^-QW\[]bOG;7D
F.c#><<V3-W@.cJA.<>A5cC>HZgNYMAdS]5/b<2-bY^gDMa);R]-[O(KWgBcg7I(
_AD80FP7<M9CQ@RH9:E\=\aTXQ+K]TT(IB=7WP&-^:&77[3O]PK<_9/G:=Z+;E[c
G+HJ/XQ,YUa5\YZ,>:G3Wef33DF1KA13daS,+b\NO>VfaFPSe-5@E#aFK7;H\Sfa
b7\YN4HNDS-W#cR77+&GZ/#+])Ud@5]g:a1?[J8ESM/&Y@CZTM3C9C7E&H?L1bF2
IOc4TEM5^S?;R=NR[Z4C/]7>>>\3+BgY?7>IAGW>J?\AdN(de^N:=^f[94Z_CNWM
c[:=/2?Id#]Z#<1QaLcb62\F-+VC&M@+L#1CJ^E\O>[-P5/DD:Q/MLIADc6-)YEJ
Hb4YWIeYe9.Q,^4N.^g=5f6<\YMV,UGV+7bF\Ne+ZU&0REO(OTA?\9ZO;d=99QQ^
J?O>e08Dg@>#g1O#=(;@\C2:;.4Z,XW><c-,_Q1<LV,N=5H?GKebc):cd]EKZWNK
b)-5dQ]#_O>+<M=+?P\4;(5)@aOO88E,AWU:HBYJc(FX2N@Q..Q6J]C&4bgXM_ea
^b0YA.=.Vb1f/D>E/C1@g#-/YK>XXMbE&35K84.P^VaOUBBdS4YHI\,P[XZYKc&<
ABCPE(&#E8..,/8.)4V5=TU0HZJ=3acFZ3?A--^-F?L]P.DaP+S8K@W/HG(XIcB5
+E]Fe,UZ-V^-ZHY.P;B?e6d;KX(>[f0/D:X^)ES6Y(5(GH1TfUB7HT6>f.7S==AY
CDZ8G8X3;aX-MVJ2KB-BeOcS.OQ?6bA;Y1(X@&:V1cR:.[_DQ_=2HO.eFdAgT4ST
\DH(E.DTY=/U16g7Qe2=6[\HL<TGVOS]U(cD>KN2SGDcVMM_U^P#1A^8=BIYD#@=
:K:\4NdLH;K[MKU.X_7b=fU/CM\1Y:dDK@fYaePW;@ce1dG9T(2a#5OQ9G_>,eY]
gF6-c)[3_<S8aAYN&[8^9<[#5DTdI)_:35&,7eT32S77Q#MbM;82^8Za75_):HD1
OZgRK^e^CI+2VJ<bQ,VY>gHV:J^\2WNX?T<1?Ob\5dGHX+TX.fLIfAPSOYLFKG2I
4]dgM^U9Ta7;NSdZA2Ue3c+)L-=VB;>_W59S2@;.g40Q0F6S.#_WSKNZ0>PJ)^_3
P(RZ+]/^?_-70GON]SZ;2@>#NG53AF+01YC)K/GHDaB1U.JZ)5_E3:[V?F=)X>>@
fQ8aD2dR7FJD@OK1A-[?/P\_f1R/PMX9eOfXe,EBLESX3Fd/,)G:P-C;KR]8;ac-
,)fZ>gf1Z+?WP0PXF^aceBJVQ/S;J=E)JMgb.b/9\_TWJ.&CV@B2bGU#4&QY:bf1
fcXBObA4R6_M>73U&&1;Z7NQ#(;?CM:8+P5ReO1-,P#@]S\eM5\,U<CU]#POK[HE
4]@bDe.FB)_A3DbHY7dfO9HJGF05J(^YK6]SC;A(CU#(JEc(aDX8^UREZTHMERDV
Q]A6>1I6)Zf^0cDQTW1FL17N;(P2P@)#@Oa+2[7G[5SN?1TaDY;,?P?bEC222-Re
A>f7/I,5P)UKD_gW)DEeTEM+#\A-6.bg+FO6\-O#,?e:-e8M=Vf.Cf2c26GJ^624
PFfKKVJFYBGaB@TSRfM^OBQ5=0:ACV0GXIF>09O;_7c36XHJfa2)((J_>RMd7dPN
H;X3D@LdO#J=6f(9PW4#HdcPQ#JE[@^.8^A&95G?5A&?-+=6_FF&2[[K]W?f][K1
;/@59U;(a?GC)GXKC@cR3QYbC-IUAE2W=A(06GT9QWF1eVJNbY^8@(DF\QX,G?C=
,V?]DLFcfA\4I/fgf^\[FDVW+N,<@J8=.&R4KFWA<0P;;/301(RKb2Z]F;13+e[&
T+L#bY<gf4OEQ:Z9ZUg:fe^-3T[dI#^M0?+f14SXb&MF&UH]A>9CW_R^F>VBZ))Q
[&geDG_WY2gb>2)WgOZdN7E/I+21NQS9;:P(g=,4:4K3gJ0O1IgS8B&CHcCFEeU>
YcQ^V398734bR,UP-)ES4&NUT<NTSQKWc4WE3[T7OQ.9OD^FOHPPcca9>gbdZXXA
@c9A@7>,cd>&F)XC-H#8:5PEgU3GK7f_SV0^=4#XIc_9R=P?\\GQ<4L[CXHC=(Ld
9\?J]eSM&:4:#<Z,EYV7]J#deECG6NS28A1)CYNTJf=T@68<FDP9#D?JcA\(+e.W
ZOZ_MX)\2gPb1A6U(D:)fS^[XAJ#eQ:LGJ_OQ@=YZP0U\_^>G1W-1^E0=@&)Hc#;
T/&DVA@,,O+1@2^42NMfIJ47P8V^7aIF12&1MQdN#aZe>gG/WbE6IedR2Y.]\-d3
;]LFEF-5^EU)b)^PSFDbg:0>D8&VLafT?_7C=,\-f)M)9<WDM>LaB(.b_<RNdeWb
R]X?4Z5V.#B0RK>&6W&cH_.[B@/^@/72M?E8?dfS@cZ@&\M>GT<VgM5BT)UQ,]bd
Y<FH8+gD3d=N\EU)1??;E:<N2LZLV?7Ad5]RB-Ne?D-_,9=2?OD9HY@20^f+\5-<
7TXHGFC#>X=Q^GIJOfQ7K.,ZHW/QYK6Z?df17FR6>H1Fd?,01=/<:bGafQL#D=4M
0?^L^<T9dEOAT<f1,-IdB4N2gX?d6?a5#AYdT#QcRI9K9LN1X8][YZ_bJ5g6\A0K
+A1W/IB^TM0#Dd#D9[f:7E7\eceI,\4X50@[V(U[>2de1([Z@#IGW_E<c.Ac3&=\
(e>fJ+N&ZH2\)ff&eV0b@Le:ZdMGb15IfSeAF2OJI+TP(UQf\bC3Tf/OP>02Xf3f
f/D>#6F@\b5KA[//F6UEK[fSP[;#0M&3G>QF/,)>50^Rb_MB6MQfD5][7d2E,DX)
=#7#BU[0_K2/^XG\K49/I#P/]]af0b1DW3-g5C#G3K?Xa;GbW48^2OHIF=53TR#d
MUN[cG>d,PBEI^X0:D<^g67cM<6WAY4RfUOJg]779D5Z\22;,ePC^D2g,?0Xbb?.
)P:[G-^O.MKV<WZ-G^.:,#IZ+2[HJYSKTC\+cSC_GX:.fa^^K^,Q)5?=ePU2dV;M
U:0@&7b@R9+1_9)CD2N2XCL\>UJ,X\)N;5:b2V1]]RH&>P/&I6]HESe\Z\6&gRCC
63Q5e,eHDUX6FG-&NQF\)I53X51CR[C@gZ[-2f:TS9QU_20^TQX2g3^#UbCDSB=/
P>(=&]QJ3&0[WRV?&.,-@+5NcaLc9aX;\@E<H#&-70fM7(9BBe(QT^QT\NbZPFZZ
B]-^[^?79cEe7,0=@&4G<R;H^XGK(-VEbFbIc2IK+4;:O0RcG+f@#XMC04F]:FY5
PM[)f,(3fN[Y;(:8:(\51cMR&DR2,+@JSC^J-K\61afN:C\_TcZ,]#I)=dT@6.5=
,Zd14K_Y750O<acJMDEN\MEV2c)S/:YGQ>W55)=FabBb:FZF@;<4RK0T(0JUN\gP
/56T]e=3.GbA[F^2]VF1T8e[MPJ\/-,eN-A+3^1X#_Q;C^DF7U9,T]PA]57Kedce
ZD6<BXC#\F89WN>B>8_fU#^+e?S]<7/+bA[JC<F+aeP8H4;b-@/Pa_c.aE4EMTQD
Y,S@,f+HWL8<GC&NdK=49b<eCD:F?HIQTQ_d^e1[_3&&d5CG8#_M-T]?]ELKLG#3
Ya>[?0SHP:05c]Q==55V)^U(ZW.5#?H+<L/fQ+S,D[X:+bK-C,6&Kf3c/H\9;-OL
<XJ]XKH5f@Rc1&,UF;c+a.[d2Sd.J@?8cM(G50MdENB(We&I,@EcAd^49KY_=G25
AT.=D/WLMQ][10#V&Ie9b2N6S?:-@7+IXW4<9WN8F,IcXEfFAF,^eSTUG0C)<XKL
W\:0DAeR6RID0b3--.[b05RaED.9GDAL)/4^[+/Ag3-V54_gfg-(_>TQ-((JPS_P
SHPdVbgFO.];H/ERc5WO:+S^ZU.bRbEZ/bLI>0YYYP^<3.7EV@>0EYQ[-\WP.b0R
P-J&.F_eCV>DXD2#/a4_R]JF@N?&J2#<:XB<:[P\c1^RR^6UZ\5,b?^B=6#gENTK
6@0?=+:&WUDb=&N&.-4692e->2G=[aA2#([c@M(aJH[YO[YY:a8QMcIeb^>W]-T<
V>Q0Q81TD/3O:./cWHg>OaI9?HD>/[J;)&[bb.=a)X:MCQ)L7.@CL-17E#B8QX78
f;^?@\5SYI9eb3<\5cI6(V,;4@5)?:d98^(VdCR6?dP7+NIVd6G&90\TZ^KMJC.)
D?CB>OaA8[VdJ&0E)3Q[DgF8_#_)g&(Xd)V\8Pf5I6O/?fHJ0fW#UGDB?:8e\U84
I6;]6B_R0;A<T@W,DKY9TW9MbK(TRJC>?DfM8b]:a_=W3b(6be<e)#=+IReURJe1
AdBKf?K^(Z\OV37a^bQ:9IZVJ?54S(J-]cJ515M.KK^(2Z8:3Ba;#I491XH6(Pd@
fHF:((Gg,\>&(SE2TVTLMOf&5AS+(F+@)bcN^&0fU:g=P7T>9X+,WOfWGeQFMD&I
E4FZ-T3_93&N/NQbF]PIJXc?URVHZ/.=M(CRTaY<B.4,]9D2.]=-<P0C>gH5]XLC
IO,QV5W__<:.[7KFb2@<3WNGKP<1Q?PRKT:H=Wg=\;BbRdRC=S2cSNV3dOGUd/Nd
<H_<2RS06YR^B9b:QN3-?OZ2Mb,:Y0H^F7KE>:K]?B>.CbeAMeH;8.?6(Vd)+_)5
4+?ZD.fg\<PdY?1K&25g9VF^5]Z7=F@#;ATO:::[.[#ZG)]&<&\b;B\KLB0@=[,Q
4;5J8<aTZZ++e;6_-dP3POAU5abe2JMfEJ@[4g6P+f7BNWXU\#b)B+;W6cGRcUMB
XB#]JVE0;;)VVA7E__2AgYS?eER<?P;P5bf475S-,#g96S32F2VP#gVfP8?OB4@_
1P7<.ZcV)TMA;[,c:;Ja+]21_T_#7N6_W?#UP_Ie.eeg,AE\V1gI<J/YZM>0C0?0
PN.IA[C](@3PNAR@FCK@Z]IIJ>.d;R8G>+KJ1D[C<<^bIf.+X&d=74HQ/_fN1NW6
W9LC4b=N0KF9aE(c?(9S)J[-GOd.ZO4&HKE=&T#OYT9dZeM4/H5>2[fOc96B;-]c
5RA(:,4@@L9V=C3:1(ED.7IDa3d\W(HZ<ELAO\F;<T8/F2F\g-TgW]9K<Ub8JH0M
B-f,<Y5GGRGE\T-5VK+JUNO,a3/X-?>Yg1C95f34=Q^ceA1]MTR4KZ0?,J>]63Q@
e+?KBIO)RV7LN7#H-O7I=4b4V<VU169J5TS.D[e/K-eEFZT@04MO]]^=;cSQR08b
d7_)dX>^N3HN/V7c&_\AD8)3KPY\1C;K5PcKRL9[2RN#\)MTYa+C0/#@3(BUATL<
T;6+/d]JA,#LF8Q<Y3daW)D_HSAfLcOD?\4TTR41JI_RDAI_dL0(DC,ZM5HS+Q/#
SeU?FG)A+H0@C6SEd[D@6dBRF;4Ud5\F;SRTOJ?SGP5KYdIe(P+&>=\87+02Z:<[
L,ANCEB+BW)#Kb^g^^gS8]d;6OW\?#YgfZ9Af?2e+QD#&E+I;<G3BIZ\eUGa&HC4
WQV=27]gH9(LH_D^1IJYB#e\QEfbB6C5JWf#;f?LJ<#2_0:.fF-Y8ZbBBLX/O0GI
RJ@UHBe@&QYKX(b].RaY;_T8FG]\.L6^SB3H[VG#QID.^J4984D]W<_/ULRXEYa&
G0c37B-#4LX(C?P@N>dRT>1B1Q604SZGNDYC>WIZSN(F?AU_d+:A8LDRT:ZOITBO
UQ,\KN_ReR/4c<9Zb:Q@3NVR6-)\W70f86C-3Yf?=4858CfHI156XD_X:]g42G/>
NJ&L9\RVHRJN,SZ1HfZI0XX]9WPS+_QQW;FAbJ2K_?FV#-:Dc.3IbCb4(+OF/H<Q
T+ZTc4U:#P7EK68TK]U]LU\Q\SPF6+TJT?f1:C50Y4PDg89)cO@2C)b<4aXd;dP@
]@LgTR36JHO24FbI_=(BA1):A+b.T/dJERK]TC(VbFf=abZ8Lbc-P;CZKBE5W\cM
J+U#J8+?I?ebQ/FRQ[[(b^J(LM<g6=B-<4.9=1]L:U^bH>-+XN\c?:@X.?1<=)S[
W(N(7M6<U1]TGgA9eTN3(3=4+=7=4;+7Y^4/#XaTAg2FP)#^Z784IN).0NgN#XZ.
][4L5AL+]DCTREW@+7R.>I&-RA3[g-S^@0[Md.e/b?XGCQ8RPETM>9D)Xb]?bP3c
5Q\,F\W#CLR;2(SP0=K4PAHNg=+(#&DYa(A?ET:YcI/WR.6?/#/K[MJ=/CPf^Kc6
3Ub[D-((9NY:TA?b=B_C\5BCEF6,cFR(8OTcQE\^J.bRCZ@8:RR?&AV[4/ZV[089
e1Q?VVCDbZF6W,NYE[@4LQ5SJD^4A@_S.[I&Z,7+&8Pe-d)F,UR/AL\=#bbc8]]+
>-PGb<0RcFDPH-0Gc]WbYI2T8b61J3U@+)U_,7[Z@d<EY9>2/HNU_Q&8N@(J]0::
_6K4@73fCL+e]M=>5Mb12.&-,X9BZ5)J[Oc+LAL\J:E1&=B3a8_C)8#T_d)FNET:
cS>IQ:KCQg6_O,]A?2gEeSc^f3M-eT[N;HU:]C43A9#2O6bC#43LED7G-Z])[PTd
[\KWHfGTdI/CWY.1IE0gdNE?FLQ9#:?/97ceJ9R.]:^eFR_DJ/HcKJ=;Q>=0f(H_
)]]PZQ16^/E6X2V+J0IPIN&CG/N2Bc_e-Z:MDC9&NTILZbKF(2+XC2&7JTI\aIGU
CH+H:WOJ4;L-gWI@31Q)20Y.K[YLTEX8SU_^,[GHe1/F=]b]7&5[#KP:_[B323fB
[WBe/+)#NO.W]W85<RS](WI7@3=SF/edGCO87IXPbF.K-/&^&XS@1IS_@B)R:R[_
0<O]I/CG;Vcac<J&DaIENcS-:SIUN4Z_EGYXY.P)d.aJ?1gB3W<2dZ4GAf_ZKOI#
[3cDKR6cfY(N(H/^T)Q2Ec(a(Z/1\O9a_67d>&^<+:)0:[VEHf<B]B]cE96fA-H[
UDI\QLbG0e5=AG29^G-AH;Ne7ZQ]eX29Q/B&]=TaaF<eYDUEB2CM3TfMaY?B<@Q^
[-a4d?QA]@TTeRXO/7EVd6I_60[G]f0OFW;//3FbAOE(N.OL<0MJF[=>]2MKO^I)
U.WC\eC[5:f9gUSI.g]EH,X1/MA]VMJ\6G<cc<.e?d617D.^Yc7QRcAe<E9E2/4:
<#MC7CC&@C&G04:D@2]+3YT3e>b?<_)cXFVU9Y<R]M4_63]aA4X-T5gVeaDZ_#YL
H3Id_J\(g))gLN47aCBW&fZL4G5\^WQ7S[MM>bL9]a1_^K^8VcJ[f\8c(f4b[+0/
0^=bVMfQIUH-2[C(Te5NCW=#OYUEeBb2B\O3,9;-P3-H/O:DVXH@;PJT4XPeV:DI
A8G_2I?dIS@0(N]Oge.T3;dTDDK5>=R;/SPNW3#Z0.cM=]cSHGL;4eKDH;Z#@Ufb
McEB1gGfRJDbaQ/DEca_?:5a8XDE^IN6N32\#7DTEX66Q41?JX(=N1[g8XQc1PPc
PaW\c3DM>gB7#-H@_3^US?A(]HI<(&C-HD]W?d_-[&G0)Q,DGJ0Fd[K7:PWYf(-W
CR4>FV?\eU3gf>VACTCW74>XM13;^9^Bf5SRZQAC6.S^cDcT?S:G)_0TVG:42&Rg
g4.72TbHXQA?.N;8eVE?&ULB>0Ub+DEbE-6gBMYaO<If3L-D_67]aXeZAZ2bc^3;
>(8=EL72]O;a7=A10W)S+f(J005b]@8;00K:;K3PE>Z-_e01H3EVT^OHZ1E3Aec=
EO8&4bROfIc<[4R&^H_:0Bc6>].ESL8_G4:TUIG^\fI:4@JcT;8&^&?^26R.=V0g
AaeRcZ/311=EU62\FZI/;4AMa>HReW/<NZN@bW0+[Ld361JeJE]VDB<(-&;&AOZa
.6P:I[g@d)(.K/^EQ@QXXU6Q\>EQW6H3#<afPdRFE^GOA#C@\G@;/L>/6UZ:W0E6
eZKCO2W_+RSfI;F5DAO8^6AM[5YD:^<2gE&S6M-VY>c[OW?([XKCRGDQ9NN>Y+b@
@b>=\(V<6E13Za4[dC34^fa29&_9C>RBTZIe9Uc.LZ]R4ZN^>GTb#1P86b[(_2^+
Nec5AIYPb3W-XI8MNE;^QV3,Pb0DR),K:W@RNG6,d@(05(TeXG6,ag@91=)Y[:-e
QOQ&CR(_DdVS9M+3UfL+.&YQ6DFFW_DD/68<bAZK2=,(>9+8\/7<cV.CSV&6gC.W
I)AR45Ja^#KDaB5@2d(TX;=a-R3MddNKLY5#XD^47\=PAE3RPeZYM89C?41MPV&T
-P&:S1Pe8/L.=:.&N#(4/Fb@^GgO6gNB.D@H)AQ\RU/K4[6e@U\6c(fW^M[gGc\]
4>G&Q1ESTV<3b;NP[d6c&#+bK]6J^UL15\<=+?=]KF;B#13SB@,@Y;2B?I]M(+:D
+(+2/XG(K0ZIYY?[.)\Y?/;g\9J8JDA;&ff.=DWR5LG4,+A>?6Tb1DZO]2O+O4FA
VbD8a9LgWX(^E\4\F=_c]W<gL3IAYPCb?16VOAID^>9O(#VL;YWD5RN]7E:9Q\W8
7eM<:;CUV7e:O#K\]f=O)K.g?L1T_3]FMA7Z5e11>.T@@-_)BN2L^=,a)Teb:ZXf
c=-98TT-IS<;O&X8YW\=6fe#:16G5dVN<]a[KRY\I939)3e5G/#9@4,01+XfR]g)
.f@=AYF>D<@/R4,aR.f?WQTG7FZP7@=-d?J0NdGI5G;3JRRHF_S99\QX1>A<3KZ/
f3D63eTPe=&05LAY+A1f64PB31Z#)9PYZ1CBHEURQeQO;OBbWD2E:g.bH+Z-(BYH
G,6MTSM]V#cEdW6Jfd)EZc_1VCL))]2#(_&VC?5^5QM3AHfX0@^N[TTCP<I]Z>CG
YPeI=,S_[JN2NDI0+9:O0YHM2(RU5W3K7OeCd\?NWF\1VdT5)BfLI1L@F@XMAU6?
/0@YcE7_.-TT)I,@NQIJSa)8S+0(Mbe;T(XU:D08])5F4E1?==3KD.K^LKTSE/fc
VH11XIQ-^6FJc,+V_cA-+#U7W6]^I2^cFF#@dW<BR>CC]A6C)KXN)9AM\20T6&+d
IH_YIS98V<:RZ<4Q.8P.1;5+EEK?-BHKXFf=c)YQ1I@,G;.X&TXX,W57^)UdH[5X
20@c&G]8O+Z/,R).fHc4?+c)a3^aZA4PW9.^2TIHAc3=.\.ML/D10:_>_D@^]J7A
LF+R);XPA67g\-E,=7)YBee03DYP?RK=c<JFGd880d&R8/6/GdP\c09bZ)]EKNQE
,A&+/Qe_6,.ga&c/O.7E^IGL?32>SdI\2&9AbM7TY_d@F:#Z--:TbTNJ6,;QKe3;
L]?<A,:@M=FI6e(4+&f_e1g.3_DPQ[M>dBVO<AC3g30:CHT0BK#10d?GO4==O]ge
<d[=5NXX6-+b@JX;]6a&).WC4<&S^D4P4^V1@Y-D,R:9MH29.AFCb4-F8#P).WM<
L+a58,fX_]>3@Yd+FZN)(^^7f40=>cUDT;;,Cc0W\LNQK3[IceI(HMAR#-Jd)J[&
+U\)^A49_@+/cXCG_.f_^VQ7WP5H0MX?VRB5b;QaP-F]TBH_7,WO:a/V.PJ#c))-
6_V4Y=#MbD,bJP.,bQ5&)EO6ATF60?5f2\@]]/9&)MBD]_FFCcVVb:1:YT3@b@P@
^PQRH]MB0Y)4OAU3HP_/gQL-X>b;=AW6>:O-9ed1\[7+YU-NMOda[FUZafSI(D18
V5\52CURcBSG8G+a)9?fCTG&d/9ZAJKdYZWO@BKZY1HVX-:<6>#5\=C?ZR\G1K7F
J[#DQMaH8_7N1A3JC]LQfI1:PSO+=Cd;317[0(=1O,N=gNB]=]73-WaWUE.UggJ@
B0+bHWT2:EGB]e=T+3F5RK4)g_1RG?ZSY3U5MI6NW4ERJJf+dZTdQ/HFEeBI:Ka@
E(83LT(VR5dWMZg(SN(5.\PNU(=a-XR&eJ)2@<.IT>_NQ;Dbf0#:9&#f=\KX^-TB
,D#&_.F<HE:G?499/e3e+6PQUI(;8+<UJ4L.T5cg[e8[0?RH;_f>:0d?_C8e/W3c
/XT,1\-&I)PbX^=V]?eg+f12&3bf]?==TfACb280c#;MVMEM<eA9e3UU,;S,]97^
0X@V&4d=C1)aV#8)R#dR#-Q]N>\[#-C14:NA3OX1]/QcA,d_XM0T/-Ce:,2M/>@7
H>-Jg=?aF?N)+9M^-3-KJGQV,g=DBZaZI:Rd?CgC:[2.0Vc(L7KEJ]c_)4@L\5AN
]RL=F?c&]WZCY4+HR-U3DJ@I(//ICgg1L,#?^M5&#L24;==Rga(d)8B8S5g58P^T
79a+7bf6YVC3<D@T=BKQ=dK7bSc0^AC/VLCLR?CHN7.2))DaTZFbTW<b.(&@9_PU
6966cP7AB_@bJ)AL-cM6U.C=@][=5X_@WEK7Og>?C;#AK5dZ\G]Kf2.[)YKYFdRU
Mc]P>8W6T63N8G#>=L:I_6bHCd<eb@DO?=OMFWPWE=)Y>3.B##7CDR;.0;Z^D(<U
?&Xg_R<_(P]#5L(K(QA4_Y4U,23g4K+KfceXg)Jf^fWR?\aB6ba8[T3=CB7&8,-A
;?[6YUWF.,2;A[Ad-P8VGIfR,V?Z(Q?3;IW8E4/&&XJ>e]=OWZL#B0c42@3ZNb4)
;J=8&#5d984#LfC:O:gCBbA0+e\PABGUV0/_K@;\RLJ=Z6ESX6J1ZaAMYb6#?=B4
HE6T2OF(>NLG8Oad/P\gH3dd-B0b,(.X0X)<XPd.7/LXPU/d1U_=LCJNU20SXMg?
1^]1<)4bKKL_9XMM&29LH(09-J9PdEKZ.4XE^HU(e[DX\/.X=NC^\Rg8#[WP99O;
M8+UC#++^^=/KCLSE6M(-UBc)f:C.T-A(L.(/U[f#aBKT3F^QBHY1)c-?:G9./fY
\GGe;>aOJ7acW;(Vd_O/Z9R(?8b0O1+3O3a5(2AIR_P:]16E]GB+M0M/(LMCQT^@
FbM,W\YVX^ae,e2^-.D+aT)b:SS^4V3CReYF#b;G4-:9]OcI3N<3@/UIP+WdI(:P
E@L(H0HW5ON;\IW=^QceEZ/aPe387Y#9B(G[0=6\2.S/>9<C(J\NP\K8@PB_9YQf
CWgYeM\T>XWLW+].17Hf8ERQHD>-C,A&YJWNN-X3_]PVKg.43(\MPN_OBFN1PBRH
Y-)JaK6X8QP,UU)&^:@YX==[M(3V._f)&RKO/1H7G+Q#))Ge=gYC,IfaTFZcP2e\
6Y<BGKKDFa/aBI.-(>P2M++BB\TVLVEO+8ePT2Y/L]g30_DHG7Ve^X:MF9<&#/+9
ONOH/?&OWGX)Kd+cc:7<#IEW7QFPK/SA5>1<UIEYDdH[RNZW^,b34gE<69\,81MW
[7bDS;2f9_6JI[&K&^WT/50&KL3WJ-<Gg2SKab&V)8OC#HT[fZM,/4/0\VRW.X<3
>5F_IVV-)U:?[/EUOWUKV)WO@:_HEXF<X[#=af&P<XGd/F#4C/eI28)]>C(TMZ9V
QIg(K&OYa1eb62Y=a?4[(Z@NWg1EUW8OCXK/eg\M]E(g)/TRg4^L5#^^9B#.G)gH
g&JUAII^-7:TR>V-5Y\YC5FV>Q+^+&>89=a_86;8<CL8&G<@eCe,7@&UNGR-5LN@
>OZf&@Z1G77M@=g7?J,-WO6_aHAY.>f]ZA4[e64(1QdW5Ne;H&fcbY=UdLQS-Cbg
Z@V7^aJf):N<:G5R:TD&H=>bZ<SGRO+KT&-NE@[/Z0a\QVDI<.<>Y8B9M[_Z77=1
I\)N4YJ&ON6d0@,519PH@44CMLB5S_H^6#9<,@[G4GBPC>]^a-?>PDJR]Ob1[g72
O<RXT&2HR3M8Z;(?>H=8(B70N=_=E9c_Mbd5/Y2JDHW4N//<RHMHI,JEQJPe#/=:
KeLgcG^ReJ3P-NBd@V_]GP>_Sf>#PDW;VQ;Q1R3R_HO_L(UO)H85UR])g4\EE)A1
/9.;Og/CS)W.^fQ31SQCgXHE_NUQSX;8Rg[]&CO:H830DW3Q)PREP1UVK8G+1_f(
A+=(E_7#N1e7/54GS2LFB>Hf<T&M8Id?-N)/eIDD,VXeM;M7#W-6JP[S^C1YQ4>[
adR[ELSZ)RU/OZ&cIRW,J\ID63T]2Sb/g_Ic1PY&JSSPD<8XJY#9d<&]Y6,N?I98
?/OaZP+:J91XZLDV.5&3MXX;>F=:U,V,(4,?C#SKPe]W6c-_#.;#e6W5g=)?Z#19
CF4b(;4Y>XJF2.:GG?DM#aULZQ5EF?AT(F586]?&?5_J]:@PIbD?+2<\H[ZY^>-@
#3fF#);FXZ[PgVX)H<4WZ9LF/WO7B+>)J^e=(N,()-WM>E/LbAU:b^XFHB2O8BR:
QSWZ\.D8=3O2A7(W:]]/?0cfWgO<8[cDD::=GBb;Y][Z7c4aZ[IO5_IF)0,D(/&C
U[XXJR:X.5[,(d;Z#R>NY39L+F02XMdWZZ&4&KR4]Ba1:&4X4[Z\_W&d=N:#^ObQ
#ZUe0->Rc[B)6aSe>)&e.M8:dLe:,D6e.2:MQ1#^c_Yfe\DdW43=gV3Z@6DN_-Nb
&QO=OKfOaZ_?B-X+Y.-@A&YKX;(E1A7^T##\Y^BG?MTMS_48fE<QB4EgVRKD1GX8
ZMd6^f&OU-V906MbA;ebE75]WHB>E5Y6G9aK()_W(X]NJCGRKY#IWg&HKPQXOEYG
04fTX@9F?Ld\9]5W+(&.(3:Pg(O2<YD</gZ5=T=F&]EIEVUYBE]DP-)5XO.Y9D-E
Gc.]eHZSO6LK1[g\&UP6ZUM5:I#c&=a.<A(5VC\;MD@H.dT/dd/W]7S;@@M_#?Yf
;&,[edZYIRN^7PaCR3Ad4HRLNUQ?L:.)aA>A>729(3&6dbT5/+G3S7YZGMK18HYC
]JXB9cI2JTBGIYFB8:>:2)d0533#ePYEB[.&EJ@3L(.Zcb3_Y>_c^B,MM-Be<M+=
/]^<#_J&]RK@YL[_DSAB&S-Jc.MaH5US_;&\DI22J1(bD,5JBe,eNKG;X[+0@>UQ
U6GAW)ae36N-2ZHZLGd.3,KI^KC5>3)]&JAG^6K&N=58T0a];I,>]=&E(>0;\2U3
KBXI<WORHW2OXb;Ea<ZULfD@IY#VCgg,YC=><B=O/7&IQ#(IQM9??34^6A6FT_;6
ZER(d]I4V:-a?4Z9F-B5^8O4A@fJZD-#Tb^GI<J:C8\gIJe)7]9L[_B@_,abfRZI
7ggc,\QFZX>(5:<XUMDA@J4\-3g(]P<3/L^gRQJH6G;2C=:^<#[69\QLBCe#]F_R
gVA_B^K^Wff?,b5RK-9U&HGDRGb&8bRKbdf^83Ge3^)DDK^G2)E]>3X#(ZM,<UTK
Z8b7H,BUF(1#cE(dBXg[N#;dKQXUM&MTcV4T\Z=<<)K;QNAI4_HR:]I=-_]2=X^a
\E[PMJ_JM@HV#D5B_PB4Kf7>>4)5GJG[H&E=_b)>N+#dMe8Md1R_+2DZ/4V^1DFb
V;XI=:B]4FGAfUdRS?LV]CFg9;7bB.e+.?)SU\@8\2W:_KI^.9[Qcb3:LX8FQB#@
6NP&+SHd<abceeYUfGD9,:(a>E6CRI>Y]#E3(I0f40N_:==(W(gTHFQV&3/KUDEE
O-OFQ.8c2=38NR;f:1J3TYf..e4)D(+.,3C1]EQKfA(-<P6@8Z]H49OO[1fX#C=T
4ZdSN;eF-&(GbIICa>BLa1]^]/K3W[CI&Za^FY(M_BFMgNH7?]@e=A>_#f0&T97e
/L1/&2S5:T<#bRDXEd:^Kb;TGN5H+bL@\6#7c]^RQacJ;T@(CN^8;]]4^3B#2ZXW
1MJ34bgIB2g&f,#3=Ya^VG<R3D#O32&K(P(,WNBbP54aURKNdKE&?NdcP8^N1[35
b_Ma=Q9#G590Sg>.9PT1SNX.LbH.MF)YYW=HI)MV\WfP.Z7@bHS^(+6A]]M@6L9c
>GSF;TVCL1[2G(#<JT1CYaSJ)I67:]7MU:_X[JB1[fU,85/U]&YWg_YJ-;08VZ>R
.&0UD+6Oe2Qg8?0e1Zb9cg<NRJ=^>2[=RF.SZ9Jb<1J7=[MFg>-YAFe5dIK&&?D<
&S4\HBNQVHB1G>,\.N:I-CSAD8H4LS\c0aG275e39WKG1058,?RQgVT[9I/Ja9O:
QF;g52W074S/]TF4U5A6ESP.OX2?]E6I68]G]E?V/+S]6aea[--0A-V18CE?-^^2
U.g]>UNc)8=7FB;d@:/7]X^+[BG#V2Ub@K?T>fWN&5,U&-W[8/&PVK_4c_2I&>D5
X@5MA^M^VF;=_J9W0)]PV61YHBAeb=HTJ2WJT8W+WDGe#dI;/dd(Lb5g;D33M<40
UEEO[a)HHD3cT?Ica>J;/U^OT9P^/>8^.-JMM-+/Z:)g[IR>ZS9g_=a.ET4P90/I
<2R9c\.+W)WI&+R6bQ(.O)Z:Kf;ZBSW1PR3J2YE:A@RYX9+Z4)/H/LJc1;J2TaRZ
+/2WI,L74TaLaCRJ86,1=f0H=Ud9+2g?&#/4:Z=NE-C=B,=T+g_:T;-_Q\f?M/+S
&&:Z?NA611e[50HDUP]QU&[8/;^Tg-)dZ^#aVPB>^^C4CC&AcdM>=&a/:CURL1PB
?2S4G9Z1c>VL^J]>F7XK3,L+O<Lc;8IFbPK26_3JV:b?J:^0HDX(#?aDHW4&>8DG
KP;+UX?BaAQ<Ifb5QBT3__0fB?QBL#JBC9.g,JP-Oc[7d84XD6_Ygb@E_ZQ/CY/O
^Y]WQfc0E<6RO\A[/+.H33[)a,Z_BGSHgZJT2NgACgb&O.PXX#MJ<ID18,:AG0f#
O48[T)<Ga1,-_#CF]^01K8Xg_)7+)Q[6ga]C&3Q\P.[D]:fF\JH_9,:>I6MFUIIA
_]-K52\6MdgcOX?^O-JIM6:+]:^BU+bUaY;7+ICOH2<S.L2Kd)\2EK2/8QIAYSH5
O1Q3BO.(dI\&62cH;EB\@R?5Bg]/#c1_0RCI96W.(O\__&DH4Z)O/dLG,gY&9fK<
_-]<W2EGJ18KQ;Z_2>?:#>8,2KdQ&?L8&_a_J@I<Mb4W9FGD2-TLa(Q@b;]/<2Ue
+\-)5(6?^P,?0&ZA:SSF^\4Y?QO#=BQXI0HT_56D^8YRCDWee\;<T\^;BP:Wa_/<
_(.Sb3J]IV(\7+6a_2Ha8C57G1?2ZYBTJVX9^\\#4[0OIL(_>2(;b&@W1+Ue;,FE
FIUQ/,/QdDBMQ-bf>TC1CPYfZ9:?P0L;,T]b&bXYO_f@TRa2DL+8@;S7^T4AZCR#
S=7QaH[)@Qf6#\ONPaVfQ=d<APROO@NWI#8[NVYJ]9N@^/NO,IT0NM99C[J9[23)
dWGAH,NBM:5VHFFUKNWM#<DL8A]5,[N>R@8fYY#[YWB^#U;\J,;&.9ASO//@;4[F
bHC\,,-]A<K,#.)J]L/64OOL-)QRAIZPLKW=b41Xf[DdOLK84M5O7(7S)H?;fPF5
L+[3/<OX;HfS=^G:f)KC4[7#afZ2TMda8_O]_d,OU1?K(@dA[4:3UZP/+T:g.f.^
f^fYTZN1I7XQPG)6\f)Q+ddKYb?_L/cS-]<<(HY>fE:Q0Md=FP1E4e[b]6YMcdYD
f=+/7PBJf[Z>4Z[UL.WdJ]F>bf/FBU2;M?:.2J0c?E>H5IVVF2=C:UEZHAV:[C3)
22BIZ_>]bCH;>H2C[(dB03CQ70_d26Y0>\/N,P@[K-e6X[bb_S/SQ1>L@S;G^FN3
4--+&(d(4H1FUCc+Hg=V<8DM_ER7e#F(85dXMbL=Vc,eaK0Q]9AaEGc:=K.[NS[J
=ML2M4UGKW#^a_:DgU6,.6W44->?DZ4AWg?<TEM?:+RER52ODHS7,Y2>_4OKXIN4
Y2<a&Z#@0T.<5f#)e:agUBH[_&@)XJNMEb<C)EK)B&>W#TQ1APLLG^VN9WT^PDT-
6?\A]900S59D3=ZIb@Z\?gd/]+F.]K,ISY00\+TEW3J:Ff4#Wa)Da\R>JQ0[DeI3
fQ+(_YNEJN.d51]74O1#M@JY<-S-\9<X\C+K]Ybe)BI(g/2ZI),bM3.dc2Y5J-ZO
aU3S5?a;HJ&S+R>dZ&([9=HPF3,WgEMMFaQ24I62GYSCI&R1,OYRWC:UQ?>/D^FX
3O9,6#cF.B-_B.DAUCN1U^HfM?c<efKNe\MRNQCF:0VWe3V=^F_7_ZV:9fX1&:&A
<1B((aYIV^>W@e003KSYM^d84VL36?:7IIgO4/CTHdWO+3G_[MgY)J^0=SVT-6MA
;-WOD&FQRBAQ&GecdCPQ+d=+A,/14&O:P)Y^<_)Z.dX[+KNUXL^KeWY\X1Cg.+@;
P4IHBLT2GMKVJ;##6:JfDROQA[ba)=SC(fP^7XLdc2Y(.(5Ub6IR:Q[_ANCAM\]S
;dJRN:aC4(T_V6HUQHf#[aUV2GW)T)d6)&e/EIBUINW25UJL<_KM.[Ee>EHSK&#G
^)Y9gG:N[BY8,S(+eObVLO<fKb##,;;AV5cX:NM1#XWG@:_?#M<CIQWg)0Y-HdFU
X#V@DFA#><7T7agcM_S-A(R>6TRGQA#G@VNXSCf=Qg[/FM6e7]<_J8\a=_Q1A(U_
^=O76GF98P(BC&YE.XG:259ICMH.<9#81OAF(5A-/0PZf@@O9MV-/XgJg#II6SWf
#B4LM4+ER2X_aYLEaC11faISNWUNSPZOI9SL]B==,FVV.GWVI/ZX5MCL0/PgZQbR
=7(0-0L&><g^UeR64ZIC\J,PO[;FfCSY:.>:bS,f&C_\+G9G_9:NEO+#B[7>&0_J
1(=\X1X@e2YbGP91ZOAAaK:g:L44V326,?L_[g]]DePC>cb/6D(L6;P)aPE-0Vc=
W+]BV#LM-M2\[SBLB]<P/+?.]16CZB<IM#_SU:NPa5Z@FFUbZ.eTYE36HLQ?Of5e
N^FPc:&X6LFBYT)XGXQR4:LDe^g[McUF2E5YQC2J[aSQeMe]eDY_J4[dUQg.B]UN
<L[5dP1FZ(HN5aY<L/N8RT3FGP690ASBbF/Tg(FE170#D>SK@GT.C@I3c)d.OGNL
3/SE&[+=ZcB5X[K;:BeZ9HgT@W>ES0g9>JY@7J0S/VX=;F[\,#A6RELI)5:D;)VE
W?2e^S0RCaKMK?4^\N-I,P)NY<Y4?7]g9<2QERBAKEZGRN5bf9EF>QdG\T8:FZbK
Q0GU=.c2.NWe45+SCRDLf):GLRcQ(Y=&/BO]#NIXL.X^/eIdW55W@PQWWWDY.W4#
2]L<V>b]]HXWO\eB0g8A<[4<,5&MNWC.YA4CC:<V@\7W6N2bKaZ0U_&cKP01O#eN
.OX8FHJC:_#IS9G-cQIE.UV-3CCd9_.ce)V4W1ga8dX0(A33\WXL3&Z.>P\W]cQX
]SP9U-D84(72[(E>G2@.32Sc:Ed^:daNdD#VUQ=#c;^(F5?dP@==/=3?(M/W=Y\U
NOFg3F=;0C\bPJMX3/^B>XG#OD1]BZUfPV30/TJ^H)6Y;+?6?/76bT>>Fe4K[PXS
E1b@[U6JR.=-gS_BUe0E,EJcWA=<^Yg8dM&[VM)F(VaFK<A_=ANUH]ZWVGe=JYDT
L71IGBaU252/9VOI/(7B2^ZS,-J_=a)BS#RT-KF9@.U22ZFX0\gdJ7OB?3UR]VP2
OI.<KG_RgR^M1E5L1P95EJ8.@>>(ZYC2;.3_^HA;LddNI>(79CGc+FVF0B1;?I)V
?gb,I@E6UD6=abLCE((DC,W6#E+OP3>dbTI06UMJJ)-cAI0ZaCLF<DbD4ISA4C)E
Z[?@]E=J<&TEI)QbZ]/,2LNfPdDV71LMe:?\V)3NdcPbW#K.C/Ce?YUMcNV@5_IN
&P[O_cT^AKEZbRTY^^Dc7/=<(GZP?\C]0S]b?3#PaH^cWNE+54+c&BH8SQV7\+:\
6.:PGP<;SgRFM)aaU_QgQeXGIB?;dM<&:+<aEQW+:QOZ),4VO,+e52Z3(ZM7;KQf
:L<:36de9,,-Ka;W/8?<Jff;I.0-RB=?Y3d4-S7?S#K(H#AeNK-.LPcg>5VcUdG5
/\d(M/_)CXbcO65d[d?4b\TLK80&fde.ZI)V#V8J#E_EH79-1Z)Wa9V1#R[J^7RG
J>8GR6,>YKFB]W#H?,D7,8R:X.8/Y+VFP;1BHJSIBWM,@(eJA]=SK4Sc]7OE>-O#
4\PLa6Ucdb@STfS),HLf;8cRA?fQYeO^J)I\F?e2cR+3>KFN16RHD.6,Te9gdAPT
^Y_(6T:O7aP/UF,B2[)CF4b2#::;ReQ=J5:W#:gVB+IBPcGf&4M4COA.6V+^UJ.g
b[E#FQHWZd=?ZWd6NL.6AddDJ3,:AJ,,bW\AacES;5]WM1-<<Z.PNNM.6fNG6C2U
K<<cQ7?8A()N57R-.((&C>P_ZM]eE#?9D=_:3gO;(bJ8WXd8K#HJ-,X4N8Bg5595
SG8,&T(>U<6/@4B)MQGScDGP<_Q]BG2Q,LILG^gDI;gFU//d7e@.5:(V&;WXOIA(
/FG(Z4Cc]&=1XU7gd2,bYJ5=(Ya(YAF(S:LPK#SC=?[GG1PCG/ET>=.>R2c==]OI
0G[><UL8(bZ-S(\RF-b@NDA<RA04Xb\MCG@INA^5IXa1^H/OL,LWcM/B[8Q;aaX6
gK_;[N:.38JHNZ(I\=ZLAS[bf4cd:PfPTGQPPQBKUB_\NQ3VTOZNa#5N2<NX;]P0
DP@RU)IB1O;B7=C,\K-E/BAR3N5d&6-0L3^WQceB8#d<.)3Y27YAe7LeB;O76L>&
OeTCbLF62(WcTA3OYKZNXYT(GVL]V2H(>]&^cYQHY\Q6JASL\<QTYOSLZL-NI;J^
HSQS8<9g(2;02O)RR+REC],.,GYVgIMUVg)dPHE^3HGES()I.\XPUgYA/2L&MILS
0))P+fTUY^,#/g=#^D[\b^_JS0J+(2e<b/<4X/(2)E6X+5PV80#;1AGVMO_eYWY/
32.H983=RMed-2:=\T,FG@4I&>,F9#)_e-dKWFW^bZT8[131FEZDAWLTGc<&aQ5A
4OJXP6-2Q\eI8AFfQRB]VZ\7Rae.#QD+cHc&FKO2LM1MF08HTd24,;YP^AZ.@N\-
58=PD8O8>aNe2+^eY:8CXc-SZ0>FFZY..C)8N8Xbg\F-/BXGfE^IF;UK_Z@Pg#/^
T(]O.,+U_fa_YN-]N8][VBKXY:[6Ie@K]T[&F>,cZ)Q)98^bQ:?J?W-B?2gYK0_7
/e:Z4\55@d.?Zbe.=d.-b(4;5[V&Q8NN&>?dDHV?:Y4Eg4FMMA#E&L[+:A+PddJ&
cD7ca:3H]@?]W42NU5.IeTB[0-eG4b,f(/TaW,:dCD<TCN[b>]00CFVFLX_:J(&G
ND2_[X1@;64T&;W@J+7DX?d&B^NWOa[.QR;Ng:a(N7/JDY?.UgP5+J5RSSVS@6Tc
[B5^AR4CK<JLL_1(X?cKNJeg/7]=Jd\6.R1T-#8@K\-Hb>P8.a-e1(QZ2/M8=Cb\
;=3DBV]TRLaTD=Z<V>;AR2FT7[V?(7UCc2^PI,cceH-F_F-TDF(d/-50g86\eUUG
&Oa/(P.D_4Ca,#d/VG=.KdI(-@=TG]OR@V1;e(Sd+ODJ286fY#)2[F?dP;O>NKZA
F:Ccg,^2P/.1eS&b?7Y@K8_8M2.G)]4dY/NLYE2U^]6OJ;9Y]K?Y4DHQQ\2F2+K@
O:5[K=[RK1A1I_(Sd_9Y?>XGe&?8<gOQP6>>CZ01gQV4/<FcVbegcJT0RZJ(UBAb
<\5QDMH[+#X4e[3\#Y4M/(W:gfb6VI1A@RT#V3VW)cASc+EV:K^&FE,dB,e7(6GY
XL@edGJ4PBD+FG5Xg6>dPF+e_=XY9?-Q:Z6;62A&G^;+=<Xgd-dC<&RL^O_;0/GE
+OST9YfE9SB>;NRT800FgIQe5E<2)9:cUDG#LQHdfN8X,RGQf[HO4eS&(a.18F\K
d4?\D6.EQcSV3>5C[J=3NISMHJ)XD(Z=<\H0D4J=.:JE)c=#[8]6Q=>b[93)eB/J
10(BQZ3ccU,B=fU#J4RVeDVFHM\5f4eI&9[Wdg?dW69WO;47_UBL?CI;b\Bc;gG(
]/.b[&Z(^6YTW6R#+(eQYE025A],f2_X/V?6-5B=dLA)CX]9EEJIaEDg-U<)WMPF
S4FJ=7E2EJ@+c&4DeI1=V7:+H]-dG-EL_Ved<<B1TcK:BMeWJD(BJd-fU5)F\#M9
ga-3Z#OU0P7_<DgF^HgRRP44_::7OT(e&ca>:.>HPT6Ie:O)TKg8Jg38KY-,/8<3
CLdOF5LKH\J4d,aTP05L,;/5;c_L^QO(VP27H]cUMbIeT[;RRHOWA)DU2Y?M=[QM
.N<N/;eCZK;QUSe9E>XI6+RWF[(-eVVRab:C<<0\d]gA)BPX/#8K5S2PAM.JcZDg
a12e;bO\Z>P8BG;-Q@6V^=c#b-/SBD8#eW.YRT<#+BC++40/4U\[gDQb2NEE1+Fa
#_6)eE>HWSI:dGYGMg5>/I4<G[^TAH&Ia\?YR?MI95_R,P=XRMR1W_6IAIJfEd]/
Q:<MXQR(b66&Z8a185>SJeE+9O&4C.1(Q2Qa6C#H]Y^)8R3CX,f3>#V=@7)^=OeU
KITNaA@?5J&P<&A1F-C1Hc&GaJ;AXIa][_;J^7+(^,/10K.YV=DM,L:d83T=SG#9
3QJ&C\GN#N<O/TIYdHLcPf39c>+.,cRDWd5J0cS9Y^IPVQ)N&W(c7//@E(?#_^bJ
K,Y8W\c#U/>I6,AWcWOH&#G+2H^;WHJ@V02PcN4O;82YJ2ZWNOgQ1AdH^W?6bVN[
,@=_dN8]P]BF.JA#._PK\#U1>4YCVMA]@5G+WOBf2a/(RICb>A^(Bc&/G80?UQ+.
U+@-0_b;/-^c9BYL/OffO0<aD5Z2)aRK1+0C3JBdAIV4T7/\eP\&1bJ+6R;eOIdH
0MY>?:(e]32,A4[+,P)UMH9EC0gETb4&7D-V\7_AUW[RG/+T.688b/)^=2MVb[-1
eBSRaF94UMDAA(UR[)C_agJa[M;4dQ@>PD4?bbE1@W7THI;fY]:]W.Hd?CANZ=6(
?M87TK/=/5Y)^/L,3<>UfW1Qeb[CH(J_1,KeOa77_XS+W,IQQU?K)H14V+VI<?4&
;7)MI)T#CF?,0&CRNeAW>-CS174NKUQ,(:,0AGTTGD_N:F/L/Lg8ZZ(Df&#+=9-G
0UgFHJC6E>UI7VNMa2=DYU<-cY+2&4Ub/JLSE@NG9gU,ORP?@^[/_Mc/SH#S^K;X
?08Y](<gNDa(;GJX^:dY(30U6<f1.KQVERZWB:V=_SVX8=a.<CfHbD>AZ?9IKRXH
U2TgH(X_3f8/M>/8T:UE-9CC=.#./:b_&5OJSP3O+N1,cPV5&?EYPJ3dQTXK&>V.
dLJCKULN/I3Y)TVQ&+2?E:bX@,g;LW_5NMD\@CL.4;[:,EP1VV]D00-7/.??J9&,
]#Mg>T[>D6VPCR3K5,94I27B1.)-EXfBc61=?<L(@40TJOgE;B_JT-(_F0J5:<.b
.MME<H=^>fNYHg[XdR-01IFZ,=#-QfPW]N=GBW&>HOQHN+45-H::HYUO/823S:QZ
1D/c:DfI)MHMMELff+</e6^@:K6?#^e3^5IJ_c@54GB;e#@TS7_OcL/MNT+63D>T
[Hb9CJgO-?+_PQT(JW=gC599,-+/_BSPCJYS9@_PgOI)P.S=7SNSBgU=PRJ7f]C0
;,>_C5^AH#4:IK0b3TLHUSbYYH4gD/f7eHFK^Lc&ceOO[7/9-OD9^;;4GQQ[;K9a
E=7P<d_B#NW>&#6\WEH;?]78_5e^;PT#SO90OIU>5Ag7FeDGYOX<N+D/HP:8VMM5
>C)19LZU)+VUc])\2@56A?<,=L2CJ?-Hg=88[XFL=/[)3PSIb7M<,@^04E:8KbLY
3Ta2X?Ea^a_8PZYgMN:,5bdM&7]9;aV^I\EZ.e.EK],[B3T7GUXLCFYR2>YNc>.\
Xd,PR32J?aN,Rg:J_KDb3Bf?2CT;L.8H=cA4Q#C5^>:NCf7.W;[5H7V5W164-D&,
^,a41PSbWM<fC\Q]PAA.2acQN7V/f;7BIP#g8&42-NSOCb.^9MNY.^HbO3_I1JS/
XNGgTXGC8UC_Q:#V@Z=)IdV-(Sc=:JRU3Ef7^1)\)5Y&]73+ZGZE:9+W0D-M[&SG
C,,N3RKfKN-gQAfd^=MM;&:@19XP0?DW,94ea>EH#0C0cMIL-fZa+Pa1Z-XfPcaH
O:N#N5#.)0S&A2=_?H,P&ZeYCUd>Pg3bc#:::ZNJb+OK?M1T:+865\^N[b/bD91V
_=@F(FYJ:RI;3V42MI6d].#eVV<I\a,eR?cH^,T^A#L+D[NT:1CH6X[c+QC\9JVO
-AZ/BF@]3+:3]d_PMfc?)#5&U@BS=Z@[Gef8OH#-G]EP0Z(HICFJfE/1Jd#L(MO<
N?P@FG>9AGcT:(\/(^(?&ZKS36S(?6?2eRUEgG\>R;;C=gK.>e^BI;9^44[N8N^J
5&L8_[,E\@<N0I5\e9@TD6[DZK#ZL0dW/#cKAOREGcCL)]^:A#OS5-221Y>e[8S8
LIIQ)Vb]180LESZ)Q;==+#H7XU9C[Xc=-I3cb#^XUa@3RfQ:GKUIGf_.a/-R)&^P
C7]Y9M]DSA]W.7#PFFKWL7696Sg^_6gWC?>,:[G3/]&#,-I,A_Nb]M1#,[WQZ&TU
V2>U/F@>Icf11ccJQ6ER?&2;6?</X\Q#5fV&7g=Sd#U[S7M58W-eLRgV1OFZB^=7
6B[+E(49P1\2C5Se/TPXb_X@=F4BMF)Wg1BG2H:,3[49LVFS?FWU8?X917f=,DTL
G#d.8B61EMc?6+OK)4V74<@UF0&I[1Rda@aS[)8A:EI[\TGG:Z0/QS].6?-M19N9
a55@GeIEZOF9WDT#f9#US5@PVFB(T+7BX.>[Fe4PF>?UX+4Og8=C(dITc@+=YWAG
dZ\@+=@]W))O,]dZ2YX42T\Id1.aKKH<ZLO+b92\FgFI)+f1FBeb7VKQ=fMdGJ6R
T+EZgP9SIK\29<V5A2:.D/6C3;:B&ULTN_6(^;LX?CC/+d/(S^e[91IJF(Y@g;I,
#WOL=cA;)?N@1?[M1Df^+fIA\aN49?9/fMD<5W68=;Qg5LJ]-c-]8];//GP(]K]O
#:G6:10IPI&g2HT&.>TH2\[Pf#3&TRW;@\P9]9W_>;<V34#9C4NFLR3&LScJQ.2P
:=LP3^>GEKRc&J?Sc(3F+@6K,:[BKRQ=^E/BR(]_V9CYA<>[7BK&I_QZ@(R;SdNG
HMDS2]<M]FbIIWEC.@35#2./;T?YFH3-eDfOG4.ESO0BVT#;LP&U<>>>HYFG#=6A
4-9)ZDW6aBdE\bR5=<b2MZc>P]88RggbfXPg2_W;GY1gRVX^,cZ,Ae[\M@W6^.Q1
;TbQ1Kg:UP(>ZTVD)PBEGR=[L3[,-DLb>5E:K>H.I+0W&NT@I)g>QN0<<YMaL1_M
#(TKJX:7aQe\(.9[SWEQV@P;^=S]NNV=c:F8(VMS&AZVYdH?G?b\&Z/(X?HTWgFI
JTO\,NeHA7+.G^[<P?&[@Lde:C5D,F?2BafaEeAf?,-5Nb>H:/ZU_aD0S(D^GZ[B
AY=)d\c3CIR)Ic_c^B3bc9#@aD7@dD()2MQ7dX=dFMO[/8>NAA[)\Mf8NCfDHIJ(
a2(0g2&?BLUE8,(TfLPF@H42ZEc1_f(PML>,]7YI+T0U6(\GAR/=(AOa2:<He7I>
]?X]bCg9-LU/IJ4TWXDf=]JBVPeVD9(ZJ[L\DO)N4JKC]^3VAW@,HMPd9NNNVeU7
ZY\OTVdb_+XNXOJR^R5J?U#X11TN7,?J.S^U:ScfCLX?VQ(/#Bb&,)M(Ld_(X@@S
>2P(H3.FFfHR^-E[NN5#@0_.Da>ET._S8+T4G0OdR;#TY4>OQ^Q93>fO21O11^gE
TH@2</-Ye1B8>W7;;_0(G/DO/[KVHB83/;JR+GI0_d##a;]cJ)NM0>@<V/FP3-Y-
f7#)6g2DAJg&FWQ@SM0TP=936HPD<<3V:>DMK+D4S7#XS.;gOW(VKgX^F-1&Kd#]
X_]D:8KP9=edIde])ZVY@O\\HMW;(C\.1RH7F+91[2E6Kb.0Z&@CK>TU7SLS=O-F
]4-QXT?#Db>TES[IPH3YC?eO9)^.V>3E@ge7^#g;Eb3Rdd4+6SbIOFAbe?aNAZP1
#N[K5<,=M&+S:ESVaR1#^<F(0f8gBXBDCPG<Z&:>EY++M5EA[Zc=I<7g[Kd_S#\Z
W4Z^T/,68B0Q5K&+g8SI[62F-^dSZCXTJgc&41Z+EWH50T7B>f=a\3]\BaA.SM;b
VY4dYZAMUd8QdZ?6>SMBQd#NSIZEKZ-V5;#,B:QZ3P8U]EeFfg]C07W,\=Pd&(UV
M75/Y7C]UN_:C^F4Q944>2IUG397RI.NgRA+;eXa#c5fX1B:1](60NKU/WIfe^Z:
H?PEK^W:3fWbJ,7IRJOb7G\5,1JgQ5\R&bA^/CS-X9O@]:T9/6?YPHDLcY(aR0\#
Q^PA@&YK8/B71&,6203U_TJ2E32EK;C036>8OMPU2#3YLV8c,^/P#O++RTWIe[3Q
g.6LF7daX1ceGMNPb\ZDWJ4fV-42^Q+++9,[CX@E_\2.Y#S7TKFU]49Id5.IJ\A<
:Ed_2<?L.d9;U^[@5K<,HF-&D2=a[LR@8J(P5dZ+ZcWL26MgBTV[?1BWXK-_\9UM
NKF^^g.IFBZAcK-IOJP\8ZOJ8K\[):c)IOcB(Mf1=&:O\6YLbOHggD29&C&4IL>E
FWEXW]V&5E^U2E^ec^R+;g9X<YbZ\)+76VC@)9^ZGFOK#,9D_3@9f^F:74(3>G#U
@WS[.M+).9EfTgd]0U-OebEKg<WAW20M7\),2U2aY?T_c^P+]K>a&IaT0JH2TCW]
[dVL&A8HGJXU=[:^He,?M)&D2T6f&SI4Eb-_e+M9>S.H)Ob\JR9&GGCeD(6_R<Sc
P^^WRRWW<3QJ<bee;8fQ>U&dg,1@U^dg;+CH:7K(Ta]+f:]4=OV^J:.F[D?L]d4Z
(6=.XVZa2[dcGFH^V0b.U]CBP6CBJEB#c+>[,L(T>K,MUS1Z>Q+Kd(&9Ya<H?gE3
J+_WT8QL2g3fCUIbPV&&FXS_5?R+]Y#9M>d)KJT.K/XgOgTIOeFN0J4>>\HOSHQ/
J\<_NDCG:M;07EUXJJ)LA7MS@5/::/9/,8)^X-=B2\dU@]#&XDMK8bVaX+#]N/8g
d\M396KdYK@R]>D;2Y[SD3X.W]U,D&#\OMXSf.g,K3D:16>CVYc,?GTA+30@,g1M
ARQ_B9+4DQ]_VA<&1[e>6SC]&4f0C:9;_)+TA#TD]4&9Z)KV]0.Ra=aQQ6+eNe?L
;g:\N<g],7&IX8]A8f3]5&QNB5(7A/PP\;b7./J.U92KHDT-A7)f=Ng8H:gI\,2J
?LCeLg;\S]cTVNMP49V85U2Rf,76fQWIRC4UKI3+11#df+MB?DeYc>-:>dZ[P0a\
9[7g2244\\:LVJE^OCSG3?E9MCYg3+;=5;BPXD;Gf1R8Zf<,9>3HJ=7&W(Q-c0&D
GGP,:3#P8SY(195SOTSU<S0B,PLFD82ObB_NY^(>IG14BJDLHO]HB5RC69-]R524
4L-S]bID85303)2N#;>2.b<W+G)g\2e:C48_OKNN/^?#,KeGV<X9_fc&[P;\c?N^
[:,O0[TK_]T(98(745\e).OS6I(,8XY(ZCaTHd^\14OZ80ZXHLKA-AG?4WFY?,PF
N24K0-V?)09b9;W=^3SEIDg:G6ZERbID()6PB)fY=(^68T8&RW9Ed>RWB[E,X[eb
&>We>1#7c3_bIe2RaF\eS=-W[NOO/BLI.M\T?b=Zd@Q4E^B==9T]5A[6d2),gdN;
8G;?T8J\Ge)-A[VdSU&[HK1<X+64IT0C+6M.LIVW7KL:ZQ:V[#T:d^M0)Xb=H=<N
GL6>#E8b3FJS?Ce5N^B+FHA(Ha_0&,7^T=H53-Rg7PKMC5bOZS7EYa-deaBH^&5a
^G@3;;BeC3?:aE)3dfVg#G0R;0\;7=?@@WfCd8SHGXW)XFP3&X\_XT23a2C_/Z6Y
YQKUEN>7W=_AV;[(e9-cSdL_cVK6(DdAYfT>-E..[b90(?K,&+gDQB@.IUZ#OGT(
N9VE.S[P\@(+:?_#66P-&@:[LW>Ec?;[5DP(UO<ac]LQZN3:JT>A_4UA?WOW7=?R
HA-d.gBV?_ZQQ4cQC1/5(D?df&]Me.DCgP/9:?+eCOLZJKX(&eV6+9R(LIFc=GcJ
D91Afg)L=b69C^<G9>(#_DT1eLcJN]bZ7Eb\Z1B&e-HS3&CfF6/Kd]MS(>H#[9S4
/EH(_bagYbB\O@<_6-T>+3A/7]J^388.>f)O&d.5d?E4>:C\O;P4Cc(9L6_Mg1<A
CHFN0>U--)M>fWWW#A40;40O&KQF?7WRRR7_b&[>3<Vd/<UIA6QAWPgdO(V1-d,0
CWFZAL7?e4@>dA7-598&1[J+]3)gO5?-bK<G&=Z+4[->0BgMX5V2Y(MH5I,@3?gR
YccT7+8-G^HO)N0e^6+U(fWJ_e9A=#/&G?5>B^9]YGELcSC@b00BT10IP22>NcI6
7&J]_e?E8e:#Jg:?MC>-M6#_STCR+8D69<Z0SP:9P]ZX.6[3RcH^gYI1bLbT@)E,
P+e;D)<(:I?WOFKbVX=1[.95-)c8E-R#Q6F(ZY3M-E/_/GG\f;KE4CQR-J[.f8RX
SHJNR(AAa>0LH8E#QL#AK)CQIQ2Y=9WeD(-JYB9\Ne7>(a1[[GfX7SJ1OQe#X[df
LPOP>>]FLed(>95>XJQ]ZV3KX/]b(;CTYM&FD-8HCJ=b,VXI4cf_QIJ9Q?V,I9&?
C_f^;K5>Kb<Dg0:ED/QI3.0O8J4C@N[D;D(N]/16MG\8Qa:ED#/X3H)g=b#)?TB2
&KM])a<g8e2FAGR[)?1#U4OUC0Q0b;;Y<PaAF^G#N]A@@KS)FLK4T[?4CQDQ40_-
^8eNOe@I7F1>a5B^g(<fAB&&JDZ5P(5JAe.9PFJ+L5G1Kd)G#@Tb0QF,[-cHTVEY
3NLPaKKE@EX//.aNBW(0/-7V2_8X4JKAgZ3<[M&/V&f+fL.L8<_1>2N]D;8Z#/8a
ZI3?]c<f\-ag[70S#>g^;B(CeKg[<V6^9P)31A461Hf1W85CdTFAS9\S8WY,2(IA
P+VPJ^WPEb]UdZ3[]>e1AI]Ia\]LX]L6_7P@,Pd6Jb>bKdIDYYd^4d,)_0@GA^G7
JO;ZFZ#RD/N-TO9B2e\8U4Fe[GaLb.Fc0IB8QcE5Eb]ZZb7=K40(F-AE[&]?>2OJ
F#OAY,R?^)4CB:A<>L7dT#K\gEB^e@#8T5GP4S[F?NP;RLCD5Y<C_-RK3<IW3L1N
9EHY&gW/9OGU&AJf7eP:CIRP[.Y#Y\?D/DB2=<>EW#?BDNAXPPB-f1A>-AOa55O8
L5SgIKC7-U1W6RGcb^BYNYddaFX?cS-Z3G^>K;AI0Z]BRd]7)7g-WGE&]C0:7KOU
NXf555DXEHW@57DYJM1b7;W?>B^I6A[NJJ7RM^9__P[XX87W_dW^(QBHI:^EYa;:
HMNE#I[H(g^D4U2MU_LAAM:S.282DX:;MdB\7.W_A)Y<V#H2Y;G^gd-VK^>V;^48
LbZV@5J[R;A7d9\Og@8\2SLf^T,A#OCdX:/5&14A&)U=CB@T+<f0_F<RESYb^c,(
O<RB^(8LbA.])12><#XIdC1e3e1C#c^4WOGJ#0AaR.(cTNKK1[,?3WIdM0:L,;,E
B<#=2J_J?c+7\?8XNDd;bYg>V+>)(3[bUCP5W>TJ5BegBDdMNg6Me?WOe&D6];Z8
OJ3.-J90<R.49BUU]HSRRUa?2W;/2e,-0+H>><Qa4ORU#B3#AZ_+7&G&d/WYJTO5
<BRa&<fCP8V<^A/G>BABJH0QBLH;Y@:Ve6MaV<6dVagMD313]fP[[H<947OB-:PC
P4[2b?IT9EP\c&LLJ:#(/OD3?L=/Qd)ZJ.?HM,WTV:IEG&V3HJ+E@YM7LM#?[dR&
DK=N4Q,R)9_KTKLX1]<(Dd/Ig]_gLHRVHfB+,YGIJAS,8A)[XP>Bd;Sd2W\8]\dX
7=R_])KdQ)&R@[-c2VGT+D&=DVX]LCPALP2Mg/@ac@T4:a4F=6:2;\^3?6#g1I0=
Z64aS2+#B>QXER[GTJ8]g).ZI18G[?Ua^N-6U)5gOacILOg15,[=8c(.;CZU89XM
_=+NVH0BB&GW[TBIV7&1U+6\1_<NT8@<C\4&/Lb1R<[#Y=_ABNGTK#HQb?2+a14_
8@acfP3-2X<>/35K2Z7)1(4-R0>\G#@\VEM4U)g[-_1AAFbAb7(VfUEF)P<=<IXY
6:,#0cgce@88[KA(8H26fI;;3NdF9V&BH3@Q1<LgT)2fbK-\_]IQ#8#WVXW;LKD>
/ZJ]WA4QN=QcE2-:/5UU8JgT.be>R00OD[N8S\\+HTaILM]9dXcIg<J,G:b[7/&6
A^8gH^O8^=#EYR?F@:a#F&5,^>\RCd+aXYNJB8P@[TE#D7<AFRC@eCWAV\[bJegG
S,2dT>gBa7X5W24bCaJJ0a(D-,N;3>#1]@7[;0Qa/&]7#QMb_V5V7C<a-\9#C:cV
LdS?dP@GBIJ;>/e@+OFfDC4M-9e[YHUUT[04P:O/]^4C@YA/3_0XR2X/f6/,[T#/
2=6(I1:Q;aR0C/#,(UV[7C#-A#,J25\<#5+J^aFZJ?SK8HOXQ-HL:;@.^(Z32MNO
&5IW4ZT]):P6ULF>ZS([</_604]Lc5NU@9@S-<g)P1Hb7a^?e5LG71=#Tb<baNU.
.fKY<Ob?:VZ9MSd?V_G7@+9+?C7.bQ+ET1Zd5<A?3F:e-<La>6_YIMNJ>W>DR&\-
Tb9B,@_f>Q=0ZGZ(/AHWD#MIZYU]L82UQfX=8#20S@]g2KD19I(,F\99CL59,OE;
Y_d.F(.PD<&RC/(D18KSDYQSMbK2D\_NQOOHMMH\1B6BMe&Z947..[BF+Sc,.D7Z
[F5W_KO7-EBJ22gM62[=/L<bfG:/BaBF11K7D=,>_#O))f02^DR_5=afQDTWc+EB
[GEea+Z0@XVbe]/N\TV@,SaP&7K=:6K1X.M4[7@JZ7M4bX;-G:9;\,W&A[YDZ0Z>
<gRRXaR:Y?X<bMD395B0=Kb1@V5&98]L[#YC[C4]5WFgH,e8VBHP&)JCQ9JHHCA1
,B:bc-?VO-AEMUT^G.>L6HL8CBa6G7]&I#,G/Q+4=Z:Kc>>9_,FRG_b:/8^&,I-&
].8O])280S>Gf)JfZg,RS6PG4e2,gEP6T=P5)6)+>ZaN\VB1Pd7DF79We])<Z-#G
Y)EU#R&MVC;=#^^=TTMfTIDS\MOM\57e;8WJ\88E+<d@g\N(DfO_LBBO/>=g86N?
A9_V\1SK25IYMbJV=5=NP[D6R@#[FT3^bTfZ5&A4e81Qa_\\F9;:)?9Y)V;UW2ef
+Z(,SBg<4+D:BfP;[186+RUd6b__K,158D/QX24(;X-cB#fCM1O8a7dZW]XG@#d1
/:#95H)+H?V?6+<(aT9g9d(.[S@F:\U#a3CAI5B#TY4c\D:aSd75,;>RcCB\/>:T
ZZGP;Z0gbIMII[-HP9HV(XO51X9:C;[]_;a4J>9?U8F]WD:cg?:&^I(^TCVUJPJc
ZB8O,&,A:BUfd,B6QM\.F&T3+YGSM[?WCaIdG3Hd)/CY_P^WGP-)=f+L&UPX,7N1
11DCB9[K+-M/d.O+]&c_(b7K5>36TRBFHNCB[7>e>b6\IHMK<8eB#Gf^gVK:E/M3
Y7c-A5+GY\+.M(7Dd;U7>I+5,JY6I&f@c35KU13E5b_eAAC(dKHgGY)5b[KY8La6
6)25R[6?Wg1d2E/2d0W.W&+XKCROL6Wb16c&3L>a.3FNVIW-3RY[\+e)>?^<S,4@
I/VaGK3:70R9#J9E3P?+=BUNBcJQ9[)UUdd-7QC_+,CCVM,0U5bWC1Kd91]O;6e5
6a]e.-+K^4/,/U@U_J,g=LM@Ke1\QX&A+M@55&KFeY;=FfO2XA8D0(g=OFOD[;9-
PfS^X(B.PE20<924/HHe.S7EDEI/\15XQME._5Ra36:C^.5@9fDg@E+8#.:2+\^U
86O]81S#=[O)&W\;0?F^ZJEgX&0@TN^K]CU@0Q)2?#VdBO->X>D5D@[cIF3&X[c;
==)TC0R[DF))/PH[45\@7I-Gd>SZ1^.J0K/MSL(CH:+[,f2EggMd[Q\7/HMP8F@+
K0gW_Ec9fVP?ZX7[@JB<Ef]M.N4fcZG-0YD2=aR_\1)-_82PJ@;+TTL\R^P,MDED
P)VT0AOPfNO.:JFf?6gJ>P0](/DA+V_1DC)^,S=]dPZdD),(9I0W.;.?-ZJ/^g63
(c[6&]<A9DVM#cGW@;&b>HM\gS8MLe8Y8d]5.M]O?b;O;7?V>TU=&6&c=D4/>Y]W
a;WB_fI\@+98O:)2#>,gg&L?6b\,.]8OR-PP]\2_-I6YQIK5YI/YN3=-9DTZ3(.N
dJUeGQ=EJ)&P<1K+]J(Gc+_?-:+5bYTg?RDP&WNa[e.Ib_+.FYL[4Q--O_:Z<178
WFeN\WRDbR<]/JY,Q\/+[52?T>U8Z+5=-Lc?9)433EH)<L>#4c^(e;EZ-#G)?GZf
b]NfLEcEIR_ZLB1:TePD_ZL)(Z?3-UOT^Y<0-b=/bOPZ:VJEVB)@[5J2SUERON2+
31L9?d]2/A>T9G1DE5-HgKP+]H+d4R3Q.P60]aA+XXcV7ZUPJ9BEc:OLP-6fC,RC
2K=FGfFP_b2:,>ENPAGR1W]+-PJ?_T[7V+8e4H[Lc__.V^9eG3,<VI+UQf=MJ8eZ
HFDO/2R^0N\ZIJ1S++S&^f@TELb;d#QS;0&H0eH):L>&?>8Y(T.FE4?4C6ERKEYg
Ce,.X?XWA+&eBcVXO#Ya]=-+b.<[/V46CX#OFY]7Ld)3.XG(V8FV;T:8^F2bYH_5
SNOS&QOHL?2a>Ve#@N/FJ3&Q\g^6?3#/>HI)a/TeM[Ab&)B1b5T1?HPG^LKe>d6^
@S&AIF/KX_eVBY[5f[89?9aPgc92>Fg?Z5LE)XNg9M]9If0=/MA2;@8&/>^e5+NF
A=8\2S.VX+IN#Wc3SX=D1<1cG0gg&=Y&EHR3.RC@@&g,V,aS<I>\O(---?X:A1XW
1A4G?/dAKX2P<c5Rd[2?:,-8V>^I,+;Yc1S#<U+Q)(Q2?&f9GPF:JYE#Cd0XCdVV
MbD?[^:2#OaBBL/YG0=J@H<I-PQQSg+LPMCJH&X+JcC]R]_LVQ@UFKR1?I2gEZb=
-XEC@OAYMTU4?&CIU2Q6CCSH,Fga/JD?2@V?C;f/#3H(APJ7)e@?MCObTdE1KF5f
fBcWcC:FB_Q#&(;L(MP19-?IAUe@>V@Y=>9P@I#-c[@dRVNE.HedBHd4b<M\GK3R
=LS<O]-KcR^g:_KQZKOCN+QHAR>+EcJU52]6_6MQb/PdJa7DYD9_Nc\;Z_WE25W-
I6JR03<K5ICH;JC:J(7HR>_AV0e/]NA8aaE1>+Q9L_JM\O,S<f,dOP6UT[=2)gP(
S\J@[=P&BON\O6H_\^cFC&=0=ERdCQ8K0.0dTgJI-/Pe.3R,g0:QLN7LHZ)A[N?N
7e87&S/NDa_K_d:69?cJO[2MJEQ\2?Xc&bgO&@Vb>)cM9@9Zf@Y4,0ILL?/O6_>[
&e&Q3^3[-=X+:P85[?1Pc6U[FP\^[f:8SCQ)a,3^#AY?F140-YMD4VVd(IEZD74;
Z=;^H,F^N]d[RGQKCL^H;Gf\Jd<XR2M_2XUG00XPR)PZ9=#R4&H@9EP0^\P^YWa@
fET&f.#5Td?V&>\a;P\46G<W3>?LQ@RQK0(3=@UEaT<I;J/=a1V3dB/&XeZcQf6J
&ggd0.d)-)ZJa/+@JK8V?TCP@X\OaHDEKM5BU#J?E;W/1C-77g(PB8-FK(EU.HP,
C=T?6<dWD0),NeI:DDX\QE<2@KEg8E?IX5<bRFCOMB7BF-,B#3MUZ;Z:d(__gZAF
Wd-WUO\CRa^<C&/#]1?&2KSEY+U\.J_c-gb9@/aV)LB)EYC53LO;QLKG.=I;2c,G
7VVfOJJS/,F:KGMH<G1<V,d>;_^fYES=M(6A9VHH14a^2U&QELE#\VX_gcaV5IU=
EaP&:N2A>C13+&9SQQ9;<X7R.OBLN4YdS>N-FDd83E(>W5HO8JSS+c^I)9@\NWd2
VZ]-2H1)#30]Q5)?3Z(_KY058AUMU05TQBf66EK?2gg0f2L>\@VCBV#BNDI^0MDe
6ZF_0[=)(?HDR>0W2JUQ3B/.,<4f34)188],V=cHNQBV4O;Y<?f\SNE[N\BJ,XT<
?Qb#L[97[/0Y:db9BM(1J3NJ;IMVT,UC0/5]P:77Y(XCUgR0\,-X)7B>;4Fb_X:b
bHJ]0_F>-_b=<EY\#Q0aJIP9c\6aYNAYGIIDV=+Qea>DM/HJHC24\:D^+;#\&WYE
?eZdI&K,(Na\UBSKc20b[QYKC03AB^3UagNKeb>#Nd(aRHOM,70GWeO?a^?;X6ea
M&e4.?TF@^3f&/+aN?c,O<TfXd36M74)3E0@70]0YES^+?fLI=S&S&^XB<LF9WR8
3ZVD1Bd.L#Tf\,;0O4fIZ2/4=e-,8&7Vadd6WV_cbg09-4W82:S@34KTgTCT+:PP
;c+UEPH-\OSSD_Ta?2OXQcL)/Be40KNI1g7:&>?TIcYL6dEP]2dR.]T,[a0V@2]V
98bQ^MfOc:64G+8=a,d#J=<H_Gb.P[ZVF)\VJS7M?/WbHX9A;Q&;O[:U36-SU2dO
aT&);>eQ_I5EP(=aRYIW?O<>^=QObUg\b[HdOLDZ]6)GYAfPP[+3DIg60]1W)&=g
8;Qg35?DG^,\d4O>]4P1W&1]F<VG:Jg8#M6W]^HR9&g2E1O@^WP>UD7K>S4_K6>Q
I9(JQ.>]+WNTgW94:Tb)B/74)P&+_).ADg^&F39X<GBFYZ:d-d3MJMH(bO->]QR+
dX;8UEA#Lc#&@/+9I)L5>AQ)]fV<dQZJNU[MN29-(R[.<2EJCCP&/2P&YCZQAHPX
.c(CUg.3?TBY2<YcJ?B6O2a^gR(97+#+fDDAGHeT-+).bNMMMb9<\Hf(]5A_Ge=>
:C?-:c.]5N#PQcF<c/5(b:@NG8ZX1IRG8D;U-B\#CY.,VcVNVe(]B=TX+)ES-+RS
22B?M(28).IME+8Af>9.N\C)XLY:bHcFO-:<OWLTSU\HMXA1O]OQO69ZCDKV=PMB
DX1f]/0H^a0P;[9a.O9]Y8[1XGf&e5KA\_Xca,)5E7)cOaN#P(DH.TB<(cPc1d)&
J_^a8d9XVKZS)bR-X^,+I_EIdY1+8\8HKF<X5[dYP5+eB@NHfeVEJ)@;[7gU[BE0
2Dce@B1\]+??[@WITCcS3;@78V4Bb6MOa\_D;BSW5Bb#Q.fd6#BI+W>8U,BW;ORG
(URS_,/V8a@a;7UfRe&Ad/Y.Q(M^_d,,WY6O6/9)]ZY:B0(0<6&F\W5<-4J;9&0B
;4(XT+#KfDaM\@SQRR-Y(:T(Nc+1,5UXa<))a#AgCa+PD(VO3X03OW>S]Ig@LGBe
^cQ]EB(6.aW&U/AK]51?]REX0<cRV7>([>UM@CZ:Md[6W0\Q??4_(Rda/GCLb[Vc
XWB:]:]dC#.a<(@<<?NZ9,^RJXA,P[:(YM4R[GAeZ[]#;AF)XAG@ZW,:Q/,^V/9<
F:D/&(8,.cIC)?Tc66TcE<?^,B8[?#<&SP?(Z9V1E?9Gd&(TTJ+R_\\KK)93G4;5
A>^9+@[<WJU\g0=3H-L;X/7O[7eD?WaHgURJVA_/0-a7X:2&^TN:0QS7ONK9KB_^
NPSYZ5<DV0<-#(8R)AMI_MEM3IVX=]NS?WH&T)VR)65OHgT1d&7Qa3)_?E^T&)X_
@[X_b63eVTX2D4/F,?SOT62Y37O6)5)J24[W@D(+6-f,e?O4P6)EF(A&VIU9-b28
TOKOXg.RaI2FJH_=5IIESEEgN=d4_PS:;&ZAa7e?2UIH2J@536+F55XQZT7#12ZN
PUX):\2=gQOIMUS5UJ^J;)NDB[CEJe_LeQ72,BeAAN]dBT=6\6OEM.b63?b-]X,;
8,bS&O&Qf.3Y)>XZ]YE4BY3R@NV_Zc;fB[&]^a24=@@,ZFPG-,W,Ye&503S39eG(
VPFP+.?T;ZRZ#BScYM65OB=_f<UD@MW]L8UW[J>FdL_+Q1G.0CQ[3D3=A0PCT7XQ
Z#YM_K)CND?\[78QB]@><DIU&KaY50H,_2>e9-QZ8VTI5_eH-ca4:/+c4@-X6EMG
b<bJLXQTGa3Ld_bK-1U#TW8e],I<;?P^;Xb4Ac,VL>:I4CCZEaUAVMCdGG?6K9R:
_aeFOTTg_RK.D)4a6W8)XQO(9^C#+acT0J(UBd5]&6?8:&Q47FZ3^<>E9C)[O&Oa
^^D<e2MJ=Q:BSZUVCD)I-?)/:M6CA2SE6^LH-eV96CCVL<R75dEPN5;L8,X3(D0]
Wg/cPJ62Og@E;8FUKA+WM\C_Y^b#9(3db2RVYE/8QF7dV.\4D-\K^\2WQH,T\+30
OdX]#1EbdQbO+Ef+DR@c1:(\&2/GG^48+CN12=9L0EUXD):I3@,#C.cP[B\Z\E+>
Z/RBeONgZ5E1?)B1/,Qg8g[Ec2(G6XL(Mag-)N9dc7feJ]a)4\C9?A9g]WQH2Pf(
DgcP-COaYY=<c)3@_Kb5^U_&YAWI51N\b]R>TG.c)_@VdF_EJ8-IK@P<[B=#?F>H
9Td@W-cAc22.])+;A58,Dc\3a5K:K.,?Ff=5IN23C0)+LH4H2?b4H8+)MMERM,@.
?d:ULgcX+RAD7^3;DWRCAFgV@#C87.-f(C@_96aIfK8V,\H(N4VTHJ?R.1)>?:4W
[X:FSRd&(@.MadZ;?86UG\S<N69-d,RUdYYP.74;3T\4;KQ^GGF[D/1WT9@cA[45
&L\gILB&FP?4gM8S7A_F<^9A365(C?b2.FVVB7SYYTC&c]T#ePB0+GSA,]8/9E=7
.:daNg^]_>.^V=QLYYV[&#cZCCH21F-df_E[.Cc4dcP8DP>B3.Z-O[O\<+7+bX(?
34bV4X/WD#>8DYd]VcfH>E+3HN+=_KKL6R]]ga-C-AC@82DSLQ?VF1BI7-[WDeR=
YS^(-B.f?9DQ@E?:4g#)1c+W8XFR(c_KC#@K89dKb?9X8H&RdTOMW1Q?7TYZ@d9G
)[Vb<[15XdQIUWH:eW:H,XaL4S5PKG^PcLT,<g:K>P>W;&,Ib9[F7\=?E#-M\YIT
__\XL3ZeQ]ED?=Z6Vg=\]gaQa__AEY(?9OW\N1R7M+>MS>R(EM\;MK?OEXfeDa2<
ANSO7W?8/_KHI[YC=9\]K&AOTPTLdOg313S)cSSd_I[Yf@&QG:LaBZ;J8]:)g>FH
3M[S.^K.aF<3(VDYVTVW0PFVN/6NKU]^eU^JA/<=0Vb4B.@WB#8SKXc+\)U68^B6
#eXWK]f27Ef5JdFU2FOXf^d.b+d@XN=/Y4O[,12.:AV/,EJ;BOF-/TVaF4X)ZeZ_
JWEa-M;H><KJQ3_fg9ZC=];RO>)OA[9a^1X.6@W09aM1c+.Z8N5#XGcB\CPF9DYY
<BbOE^(_NROMUC(D#]?b+OCY;Q;[?/D<b(8643_/BUc<e)6^Gg2=5GWdXH\QHCA-
[K[gS\QVEZM<&BZO#Z+YT0W(Pg79+0^,8L<B8V2R1>44HLQUeYX66W\g)Z(#O;?(
F9_a[XM.H:KDOO.D)b:X2686P42?PRN[Nf-^SbY(aaa^:>.a8P\R(eDc2PU&NJ2?
a_DYTPQ1d<\9&HMGU8=9TZ7)I(N.I9,?Y80B6P)[cc_GFBG2QbNWJ6))5g<#Jd#A
W1SV#0)MSd+@VV-3PF:c)7g8X4dOA56&\-C-REK43;]/JYVPG2bUe0<W@\^PIMd7
R</8(0^W<RY2FI)&8F>AX;R&Bca[M+7L5412cgXMW>:0\21W6J>X9@^df.WAX&.E
:^(1#UON>(aO(YV\OAc)X7^(QE/8+/,c54=e6>R\d2E]bP&@fL0<></4WDJ+g.>F
@8;N,XeK_]BQc[(P2QN[69ZO:f9@Bf3bA2;#e_05V_^16AUB>M3X>WE?X1TCXOC=
I1@#.7JYT3JBH?QEH#WQ?\A=AM[f3H,N_G<PD)Y6d\=1HYDX\-Md72F4=+IVg,F7
3BYE^fH\6N\:;-0K:#A]XBT(WP]F[740V:W:0c\FdK6T:)^LMI@6BagYA>OEK2J8
>eSV)]Z_LEHTG,[g4^:/c;<Je\EdF)ET(d=6AD0LN=M5(>NGQc<V-;e^UUADI+Vb
JSf3_#^JZVC6GZE76TUDY>gRb(862VaW&]gQ9<2T(X>[<V\><=]2:N2Pd[YZQ.(Q
4&+gd4_<],b\#C(-Y?egTY821,cC+GT=e0S2B.?cBMI+)]Mb3a#SAcgb@.(\\agY
_b+AaXZAcF6cQ:6S?4Q\-SA]A4WcFGGMfFU2RCdc<2?=4&B:]A&1FCR-S;A#U/1I
+8.S6T#TF-0B4)LEMHD)1H.g@5@JWQ7_WJZBPKRD_.H58g8)G.e5QO>fZVYMHfa4
6T>ZX+==8e+TQKJK3dK&<&O98TOg&UAE1MRVeg^3P2cS=&?BYQY.;g3_NG+/TEX.
XPC&SE=7^8;ZRJ+A-46GBHYC64deZfC/O<0#+K0IZNI@OP1@O;Z9#BbL5Vf1R<?J
Q=T)PO]@GaMK];;M<7bVEEVEP.f(8A34AFge,Kd)</\PbWOU5P>cD0[MgG^H4YH]
3/e1M<c&+P]EG)<7G,5A6V1^&-:BT2B_&.f]\>bS=5]6<0F8dD</CE?](C1//cK@
T]]-0fFVa@_0&7ACF3^&a59g89_P:[AN/@T</0)),4:4d+aA-Fab\<(C2D33B9HY
5cJ?];g^a5bBb6M\X6aMAVF=3,>ZDU[e6F#SC/71.R[;=:UN(X+V\eN#[7bWe?6.
#>2_bPSI7Sg^W4J+eXZT[g+]A3#Q,e;Xa3O2R9+DG\W@Z<T^U8c0gZ9GU>KAYPY-
b#,<O;d\?3>?Z=2_&A;V<,QgE;4=F8>5aJ_;GfTG<L[&DN/GHJ_g8..bWK<J_Vg_
[5VLE<MGEW+<D6?^)e.)&IXa8A]8ELKC=Z19)?0#UVJ.A[>M/=WHWM^7<TN]g;?]
9/7^-43O9_cdfUNN]=X#:U1>=R#;]cCC_Z^B;V\ER\&A&geB-J.cMNZFPEa,C@0d
bQ36KK]&>1Lb(+K/BXeE76>CY0^0/AbOH7<YL4M14B4_4/F:EF>9e)FdG\dcS+cd
?4L[W0?2?P@)_>\(JAEHUG#_gE)cN@O;D6Z1e\:P.>]61LE(_O<&<0=GKVDA=&7E
\X,WSJK6[aEEO^XX?&Xa928[5acXfgKNO>fUV(@Q^.ELD>b4NWJ#V-@a^2BKbGc:
O#>_JS/J[C/G9CS]gWG\_[2&EZ0L]5O?U6EO5K#V=L5]G1bJ5MdFYM54/SW^L+2Q
P#D+G>U;#]_L\CD48DJ^J?S80AB0f&E_GLQ7R&SSc(b/a[_2K<Q)(=3S-9DK_FN6
,S?G0T#Q7,EY_/LfH7G0ZA[_:LK?O)ZSUBKT[(E16\e_U8^\O4F:)-TW&=4eS<07
[Ya_N4HGQV[<\=DYYY_I6Z&bOY715Gc2\3cDUefbH2)&0T<CJT#;2(Tgf]SM&3O>
\9X9(V&1TDa@YSRT92dUe#P12<_NL1P7=E<.\S.YQ2d7IAdL;fA2X]K]SHV/fE/@
:e,5>59UE8\>+;dg\eFX6A&5V<4Ae/XA_YbN<VDB5]8@9M11If?>@(Y&9/b(O@Q_
(&27Z4c^#100d4T7&g(D]NJgRS1GVF@[9[,-^3>.L68/TdOR(gX#f&-99)HPPfF[
G>5G[>9MBO>\P.K^;EgWccdN.f9V#N/>7;MB_97GJK-fDaU&#_gWgV2eF+Ef>YM[
M&S.Se9#1_BBT/_1IC]K_?8Q\\9(f2f0WG&YP^TD-eZ/I@2fVCL?L-/M.GV/YG(<
2a3#&-DZFE9:QcSKL0U^a+HbYWBZf>+UcX\eaXR_T;^K+?dQ>aCa4_<,3LAX4;cQ
.F^W3-PBNZM#??3?YQ1bRc#8F_,efJdT3bALCA1RfO6:SVPYK1\OI(,M2.1MADMf
d>G#=ESe;(LWUCMNe=AaXSf2##4@HT#<?1T6+WMNT-0f;.]\,=7C55+=62deD?6@
H:fMN9b@OB.MXcZc]M5_29#XRc;#7.T\YNLJOg1WZ-O=O62fWaGb)[,[91G]bb?A
A8W8NYU5c^P(a4a2fD][OI]Q)92b(/a(f(VW8\W0_IZ8G7L/U\I1daTTX.H5cH^R
/\?:[]48;TfbKf/CgYCOVZOc-5S/\YQX.9GB@9ZCYA^ae&gG7#WAL.)Q=>&48dHN
]Y<Y70Bc((1+<0Bb2XWTBc0eEMgO=CSQ@gFSY0+D0D2W\4I_f.:SZKP/3VHFVJM[
,K?d]Da[PD9G-DaF3K(S.^?gKb+?:PE-d3A\)J0KHbSQ06X^1:/^>=X(@N=9]YT[
Sa&ZP40Y/=@=MSFS[HD;aUL_c8BaSgeaI[g;PgG7CUT@OSX.;@gEBXfO8QCOE>Q\
U/Rd>O+dRY(S20\>TM)03&PZ_.3=8SdTKR)?YS3Qcbg=P&>OE:11RaP3^7[#56eM
OBW2>S52TU)EV=-EQg:VcU#0U=g2c8Ia)]HgQ(LKd]^4Db<dIG-_ED\&[OZd(]=4
I>FG([Z4#?]_5;91g<6N-(^HNSO+W]g7JBGX8&/>6RfcPBPX1aI+?[_&2b8\PT?Y
:7b=BMLPK99ECaCN:5+N=VDVTeKAgF[F\a+f@Z6Yf?;I2=V3@UE=RC(W-b#3G4Qd
J+COO,&,/Se>)P>SC#,9Ie<N=7\OQ^.0C,\^YGF.->1RY?T:-OPH<SY0f)GY4F7g
GRgHSB-N)LC&bZWOR/+EI9[Y=/,0Ib=<78A_G#cYW/NgM9KR^LF:1(A(c@G2E0-X
G3?[S5U[Q-CB8M=2113?,#P-,\(O]MF)W=b[.:JE].gK,9MQIgAW;7WP8OWg#D<0
bJ,Gf-34KR[POdAX/^7CRUc\>E7>3_5KAd^3-=GNS1=G9c=[<KN]NZJ1IPGPPENL
ZW5Q,BgcEW\4)I/5<HG(H0>>gH#d>G?I&CG)BC.]OWRMT)(5HW4&Z@dTeFPQdIaJ
SHG_V7+99CX)WNOD.=P#1?[bN\)VSH9)gGMV58/V59S)#I7N;O:S.R+-)=<Y=ILY
1cfMbTg<-cM](-fSF??4>3PX;gbfMOOW&b@_cOH(>6e.81bZ1,g-L\5X1Y8,Bb:G
OXZB\FC72e_#Z#[F0MNd.?\>[Z8G:OCZN89&FOBc>;4W78V]L[2)9aJfG;@Za[G,
ES@5F-c+EV70FPPc[Q&B(J+ZV2S4>TKg#T,=\U<Y@W.1FbZC0_SEY1#]^TXOFB]H
I&;4Ab<^gc1+D\US<[OO=RTeDQ7+/2PLX0M)T3FHZfE9#&:ge_OU(F6W\>^ICK3b
[7=7TMa1VOI\A/ZQ<:,Wc]VAB(K\TA2P<aA163=6WX,LIW/+bJ9-Tc1\3AaH]<+Y
SY#XO+08\aBH/]ecI5ObE,JV.]Y&TS0PaUN]-,?_P>9B@I2;<#_UUXcf40d&#cH2
]V-ZQ(b,1@MUXPE@0e2DH;D^b[/N,fTG=B6Le^L2_ZW:Y-S4THL2e5GQI-Bd0+:6
+e.#4X1N?.L/?U8d+>3-AD;+)\e17)B?\73g+4eA2P(<,MYKU(>+g3;R7=B6Q38W
-@PQg/77g(23H3dG_9Cd#2-+eaQWD&7A.84/B[NZ\1e7gQbT=@LT.\HK/-<=KM]:
,BU2QFX#U7TM;<GHVGD:N4Y.3P3/ASP(20c,LJ]VTGU&d-01)&@5dRe;73FAON;T
D\XM82]<gE=3[)\UCQG:[<H-69N-KI(&d\MPFSg2-+-^F.SBdKd?-=9R;@(/=f_F
51fHc0?W9d52fCP2;dF[KMJIIcL\=d]WWM[R2<543Lf,1aVOeK/2f>,W.?]5aUYd
cJ+X;FKD14MD:de92LLJgg7T)2<LZM7#2MU5;^E+_E<&SCZaH=+:9?O\4;0_eP[N
MI6?fQ4:_?A[AG0.@W>;4V,?&+F>WN9&7(UJJ?53>dU+aESR<DL#WD:Tb1Q>Of3g
dZ[EY4Xd@?5L@=b-F##McVZZ7U\=S(R)X31?F(BJUc:d[[Q+EA)P(d57.CbX[QO0
()Y:dcD/4N-B[HF_TBS75Gc@2P#\L2+GGTDc?XW)LWDI-N85F^1MW<MNca=Vc=PG
ZLUAKc,Ua>:YFZ04-fV?3N_c;Y&B14_^MBEKaZBf,#>QZ9Mab&_2L^NG)Pg338,X
H0V)3&.Zcd8MN/eG/(Y^5\WYIdc<2<9XTR<??<R(Cb^bURZaR_3g(;TP?cF<Xc@#
P&+\cPf0E@70&+)bOaabW;@]N=;9P4dW+?]P;eQ66KReJF<SOFIBeDMM[L1Of^/O
1U^B(0WI=b9NYW_/2J1DM<#ILUee?0e[IH4d63V1:V)BG;A&4@/QWCg]a[T]-ZW?
7J>&CRAEf;NI\6T,<B7\FTZXZ)OJQW#Y)?^QPedgLM4>E+e5d607fKCe-<J2(W4b
FZQMY][2fR@aC7N@66,OSW\ADd]#U2D_<(,R+.^<:IT.M/#fAPaW6c(&,^=&O:L#
.D:0=9DE<5>LMW^d?O=6<a<aV-)b,PS7b[P2^85@K5\]H_F>)S_5@LG+=__QBZJ)
+gVIWaS#gKX<N,FGT:>7VV68c07-G;?cYHM#-&C45V(FL2168Af@6:bD6YC@SAEF
_6c[:01e1,+>2\N),53A6]CXEZ/0Me5P]4WMR/gH/=K46Z,5@VF\Q9(G[&9R#=I,
f3NbY-/[&49HS@C#5EGA1VC.]B9g[]0QeA70eGg(=8[DHVVD?>#7MeWH6<+-&\(]
9-#?<fYaSRJc6[85]I)Kb3;T#e<Rb6)+@>AOa;:E.f5B[&0fL2\(5T]LB_BAfgE=
^XfbN>aeGK&86>M&D=.?6;=fAH,=6+ACM:Qb]6:JUZS-Q9SbEQ#Y<;=T>:AfC.cM
FHaa^d0>\g/bafF/+4]/#KaZVRNM<HI9<e8^-WLUH;&a,[_c92/Ge=]X.A1=3HKR
VgN-NF+54)[]@5UYBE@[4Sd0HY)f_RAf4;39B:^MY-0C_a1YD\?8_T#4=(4G^8RY
^YDKa0L5Y\[C13gH[,E4.M,?&XS__H6DdbT.MN2KRTXVNcAJNHYCK;-Td(CWR<F^
<ARZ(4YN5gX#NVe.5?O5LGT;Y\E;:&@W\2f<E[f<]1DbL#bH)dCB,Fe4b0^,C,=(
F5H.G+HQC0WNZ3)-K_F85=5cR]eOfFEG[4aZ_FI=cCHYd-[8?GE31^KNR,,Sg?+I
X5K/VdIS>@8Y,4:<JAbOOD,B+Ae\g6\OGYV<;Fd0B/GR6_\fCKJ:fUFd39OH;]4F
#N#5;8E=cZ^fH12VQTaa.9:ad-SEP<K8bf2]^F<(&C_S<&OO?_VV\IMLC==&0O-(
:03,0+eE03X05W>-LU))BQ)#X;-Z4.<3@)_D#C1U@0;YUDL-?Yb#/dC^7,BU:WU#
XGY8Y62cVA1F51c>f8g1K?e-_>W0&<::(D6T]13P#3=DU?)FQ5I[WU6EOa]9Qd/F
Z&V>-,N<VTN=MefX_QB7_?=\0+[M:[&_c-a2ASaV2.a,3bFA5b&fegFO4&OBI5PG
,4_e<Eg_Ud_B[R>VYf^F&e2_fd5Q;M>74-Q;&RGFHHNJ&C?9d94&(2DI?D1N+@[:
S&a?Mc.UW:V53P:7#@f0AfG3HNg=dHB^7?L8f,b/3IP<91E+b/=Y\P#AGDJX#5Hb
T^,MQ,JND,U)7f,3R92E,10VKP^+gd<,c3;@D-IT7]/c7JeT#AZWWX508OUG#@:9
L?@7gBReb)MEZXR1:N0]<^<82FS]XVGBCXJ_\Q2.SAR,.Y7^@\-:S/I?H06J;.e;
<J;=>1A^g?#HO7bTaGO0a)=>;OdQH82QRB[5dW\6/::Kf52LIW(TWLN-JCV\\3J5
GQ@U1L\bVD(A<)APX7TU;2bWJLJd5->;8,=YKR2,X8#UUACgZ[EWB_<IbKFbecH?
]C8N?XL[[4EF]9(g3J=O5>e2))VWDe&ZZJ=IJFN78MBZeBT?6OEUVd8I7bebX.D1
,(&)6+7fK&\[,@f:(]3CDD+]>D>QW59+/_XBV2&HDO?QLIBJ1<0+[L2EJRdIO7K.
f6Yg&D72D4NJB#7e7;A3+/9O2Z8)C+2D/EA?Y@NR(,g^P?_(5^R(_.&HWfX(3EH1
,&[])27EEO8JCJYV83Hg&V1]a,-7W4ROJ1^.R.\O6VTV2:U4_aI<Z3=Rc3LA^I5V
AH9)@eCT7,7YS-\145?_B-:)RZEf()A:U0YTdA(D:GOPcGF_<AY+[-:5]FG(0e:]
CV)+3D>6fA8;fEYXfVH-3VOL.8^W1(=2K.dG-=+U75gRUG(7RLSPCA.T0OgNDUI<
7XB]=29CS3L(^cR,144GJV>&ce1QQTSP)L@285/.17UM?E-aQ_IcDTT76M/WQCT8
ZLAB1@ROGV6>H7a;8>HXP9?2ZC8.G94T7F,=44;V=BEKAQCYgQH3Je0;-g\C_f?:
586-1FCV>^g.3E]dZd?,f2.V[H4MY=@;H4<RO5-Y/M>ME<48_]@@29e#GGS<E?[A
[gR<e4ORMC#MMCPSB#0eA@e(fGVG[7);SOL.<WS@+&.+//cFKWE,Rc0d;+4E,fWT
6bT9&Z&]WPG^>=MUM&bKfP0K/-L2Z=>EAG/JVbOZ#AFf#PcA0Ge.H]91KGUDSS10
00W:E_JLcVXHKf?2^)PKfLGW.#QTGR+/g?WPLcKeBRR6&&3SY\OG1gc6Y8GQB,W[
+Q[C)>8NfKQSL^gN._#e8N=]UXOb-M75Yf#LNc1L^R\@,/UXLcM9OTL7Q3Z/;K@M
I\7P+I9RC,P[(;H]G4R>a\WNB<,e5bGG/5E@5R6UGW8OJ>_/:;R,L,7]_/+N=.6#
Cf<8J_I4^d48b-H>1WAg44;d)#/&^eQcP+]RCTOL:.5^c,NU5HVW<4HU=Cg@(2DU
(FP6\<\9fE^&NCRWHC<.^X-M@5@6V-G1?_Fc+cTTcJD4VON_W,13H4bKNQG[La2:
29W:N]C=Y.LE/^Ia)-?&;(GOWSLA9Z<@.[ISX8ZeJQ&,[d8G/UTFRW]M+<[A#2NH
TI7_^gB8]4D2:G\9K<Zfa.gg8MG]ICKCcQa.SXWHc7(=-RJIU[;bUXNP-;#L]gN)
#D#?:8Lf/?e>^^#:41.J\,0M_DO,6]9\RVWb[.<G\>WU@Q7gYZ933IA?cb0][+.a
KY;QcSZ-F_BT1V2[7FM=;X43GdNdCG2E2]b2=O<^CC]1_g^#NL3H@6dWB430Xd7,
;Y@?SW(<+UXBFH5f9@^UF1Ka1?2d-Wba)9AA_43,X[S(]RKYag0[5MXJ_I(c([)J
YAbc9HNd,P+6b&?PBKJOV&.FEC=Fd&XcNK<Z5#ZQ[,FG&HMFGG;#.K0JJe9=-(<1
9>AcG/,S]JcKL7e=d5SEV21C\e-TE:CaP9F<G-aTH54I6Z62U\JTM=-@dVG)-cG5
,6E-dVE>-b28g=4e-(5YCLFe&^c#IS7WA7+d5,f]7DR3.862I1Z==.UM(CGTMVe-
@NIRVcbB(a44745;T2U[fR[A79IEd>1/UJR5YA4Ea7g:Ed42]XZATV5N;E/_(YAG
4;VTYV>)6(?3FV>T2bC4E>?\JaGN#M[TD9;TJS:WCP7&RS4&a-<a)f.E>RVdG;V9
6_LZPb3+9ND;WSb.KV#TI74-Y:,?^P];J2^A&Nb[;F)7M_@TNE9>(1J.g(EMf1(W
]c^SPEGR6gEbbRfZ.EJE1&NK^bR)@@<M]B:BZT<MB)3g/\3AP39b+<3e[BgVKZ>_
&XQH3_BVg4XfV^KLPF4GZ7YP_4T3GP6:4CNS0YDK\S(]^(D56]F#M=L^a2P)gJC8
GUaGgXGYOb8HPB2a\+GV;Y:<M:-6#/ZgMBaM+&VE9J/(c]P=S4bBg-+0Q5.SJG-<
OfEQT\a&I=G70ffQA7D=HG_e;A&(W+0TGf;_Ne3WU8c?3CPQAK-ZH\U;@c.UDW0D
EH.&47&B92AM>O6\0R;3R3;>0dd,eYb[T>WMW]e3SdPR<:.<A5#44c[G1.]f=^dV
VPHg9\\X:\H5SP]Z:+b5=62dd1Wa8?19ND3dMF(T9S^A@cMC@_dB;>&\&:e1AF[T
[cC/51.HLd^/:D7GLDDB,.(8O,ca+>)]U9LIgBNLR+@gWU^7#P\bC+GBd7&_3.?d
gPF1=ZW;G-f+M33\5dZ6D\TDeMPP8:UX5-\TLa)3([A:U8C^[fTZI3/MFY+24]\X
<N:H<14\PVFga3OZBK32fc4eU9:(,fD6R:RBIcHM\CQa\HW[W+5JN;6([bY,M>)M
YKF<I1,22:,FMbX^0b&(QA3Rc=N]QK_Ub-Lc0]/S<C)e-c^O)XHZLbZ4X9AD-1+G
:V6L7C24?KVD1e<]A?\D:;61:#a1UE?DWP:Ue&,-egAM<cV=A5<:Je>RKFDIBbK8
&7d#]gEC)026G&_a^@:^NNeZ_8FbO)^XRe-E3IF3+bI7QAAd4ANF.1<<YRS[Q\gH
-DLF9RPdJ<.bC(P;3cZ58YJZZ/=]F6]R0AfM4-Z7eI6^6LB6)8\>5J56db]GV2SK
-+ScVSRS0db#cJLE(a\?8>G:XD-79)1Z_W@eG3>COQ3Aa()&>cb+3ZO:XMcIZP^/
=@cU]<N7W^>L@]-XVMY4,c49KG=e8&7eZ7GLTcF5XG5-L(E&AP/aL^+VJC#;<NG;
JO[Kg^LJ^&g1QKR0_aFJDJB22^70YS]ZBK>R/X]P.:[1ff(]BYWdc\TO?d3OYPO2
cF?/UR6<eA2/+(5&\SUBSf01GAB-<Z4GAMP8Ea217.R93a[b3)_T,RZ,/e)/Gg:&
e7?aQU/B8OKF,M7f=[C__:eY3b5GTDK>M?PDXX?+7Q])#<GXA+HBY^C//GR3U>G?
2R\[X(Z7(B6_Ge41A4I1.MVBF7@MEaVD2AHR1C&[FP)(Y@G76Y3YcY(8E?=b4\FQ
<&JVQgRB>9[Q>\10C>K(eY(]DCR/.=[7g5.INKB-:<^V93<&>GV1bAOH3=V2VK7a
;Ca.<EdLO@\+LF&A6/KXU([c_)-]d/@L^N&K=)Q9J[A@RX,Pd_X;/fgL>(S+6fAB
<-3,</MF7\GD0PbAf0AMg#<MK7MaHJg&T#(EM)08,XeR;\/J5Ye(VB+DRP=[XK40
N[=6=Hff65B>(0gB_.9MPZaU+T9KI+X#0XY5_,79,:SbJU)/=.A2=MP^VNA&3@=H
[<QB</gV0VYS9/^c=^70b)WZO(b?H)b/55JZ+A1#aWVf1;,^^_#:<_[QTRI0Fg^F
9ZebG0egc,^K.6,51?;MU5_YFOfe^QS1X1&TUPXbN_W8K-2]6cGG_7SYB,25GF>c
ONJW4JEG(/)7,feX4bI)NP5b>V-a,O<3T5JX2/IH>VfdcReg/7S#J^K,&7-1L^d3
c\OVYH6ADSJeS\HA8;J_X[:Q>[<WOU&TO><L.DV85cfd.Y[.EJJ+<&?CfU<dE9WK
8/BR91SVT_,]8+1bI0D/@][X.9D>Ja-a><HXL?(.^A[(4V31/Mb0\(,dUdCV[#.;
.GH(2F:8S9>?1T.dB6[K4#0Y^)gA^#&B:K75\Q6_KQdXWGU5T]7@RK;V;b(GY)S[
<+?6ARQd^C1=g[R40-\INN[<T:6JY]QH9EgfCADIUD2=I3JU39c;2N3baS-c@e5K
0;4@=\/OLP\=NE>_IRXWBW^9(aBfK_N.9[KfX<8XS_1;W^[OcHY:f.bW)XU[+=T/
.TE85]fa@B9?HM:0UFdH:18UYSK9c74T_&/B/&F4eVEVAOLCUYb_U\[W@&@_NX9S
7[)(KKHa.LMBVa=UIO<8eH+QT?d8KE,JQd/?\I]E.K81-7O[5&5TSYEC[@<?7a[^
\6>ATP]50.<1DQ)F-1E&W\_BH2WB[P=YTPM<e;JBVAeC6A^?UeZEMF_c#6YQ:MCN
dM-9YH/&6a;V;/XKM9D6-6;g,fYK,IE2.8MR43D,E9G:M(7=Z])6)R6OB5JQ@7?Q
f;.XJL+TgcFTVQYZ70+:N^&(R/=R]@+2U(g2/CW/(JH[MBAFF<A&6Za+R-KPW4I5
1[A<C,WZ/fSJHKJA9aQJ:N3HfOPT243BAB@)f6ZVE[>P[TgMU4MZA8/<=B3)23dZ
^K7KNMQ#:#MO11C)/eO^ESg,/:.Z,8LOC7(d5TE(8(S:39e(Hf(-ZMUV1dOOca9b
TNaHIcf+MT3,+]78QX@/RR<ZT_]6_abYZN.e-@Q:3I,](GSBZE)(E>QcJAF+=.X0
OJ)SM:8^T:fR=7bLb0G^QVQ0MH8M(#)(5\ca:G)G4CK:EZNgZG/DG0T0cBF,>1cU
;bO>A(0^O[cGCgJcM3@]5FJc&1TeUWXY8.G8bB6+d2Cb7Z:=Xd=:.[^FMgIYDeND
3O]C9:,62.SdL^#A_8:Z3?@;/^TcYL1.KG)0+@C9M3X>@#<0\O#LV&Nf0ZG#-8E>
(;W=?3H.\W3@,Se[WR=@BGW6a(4W4)gZSF8PA8HS.c]Qe1C0M_aL@^&XS8J#GB##
b;@Yc]^d#L2.8L2):CK4];\a\8)>WVRd<O.M_Pf:-ZL.52FGL[\,FP()5>5Yeaa^
2^\c&C;],H5:Gg1Ba\[;I99R@C.OLB:I96[(N6Q/D:gHO[9HdeW)(:O^8DgTZFN;
-[(JBSSHB4Q9#G_;fDCS2HL9FYaEJX==B=,4]=6(?c-+#Q7NafDZc9C))3)20;Oa
_0RJR::3_a40d8PGJA+Q(U\H[GBQMM,]X7\ff/4N6W9e@QD7Q@@=<R6_70Ua=2;M
4c<1:IYPLK3g-R<\F+CWQ&59K/fWBZcJU#2:.3d=[X3#Q)(bc?3ca^bc[B];Y798
;M>A[<UJ]J#8=9-UF5D7aOK814+TPbT5([4KQVg54X7f]T:2G5LE4P_g:B.KgWPS
(ADV]NDDDO(QR@P820\\TL2?A48V9=U-A0T^1]O,&H9\T0+DLce;V73NR\?3M)<P
UeAR-9I[6U^/O:M;)N]>E-a,R09fJY).9Z89LC67#+ba.7\3?:AN\4Ybd4I2:c=P
HJdK<KBJLK-2?;bTE2]g5V4(fLAOK6_R]d1FT.)WOC=?:=_e#Z^SC^Oc,(PS-c)?
X+65Ne;Q]3Dd&8fWdYWSL_^J^#_^=4_39<.DHU\>0c5^_ETF/;;:)H,2_B<AF3_=
,MPMBgI(JJ#9dYU.L):5c6\Yc)2[d9EPI2+8&,b(/Rc,f9T0N.,a0V_VOZbd^8^8
GQ><N^Se,@_/_QQKXD(gN=,4YU#0][+/393[J>ZEgHdZ_]W3<V7PV\b9X0#C/Q)A
KHGP1gQETYSS3X)I=2@6RYMZ-6^JW.QPGWIVUD[@;5=Y1B(+FI7Wg-0b6WU@?Q5V
75DW0TBf6DIF4\]ELDE1IgJb5>e6AJ.dQ[b>9Z5bSP-75>gH<RcF6T,aH]52bVe^
,Ye(MaYdUM6Y[>\;TE+6FZZMTXQF6c3FdIHR,<O#b)Y\b<[.H/(X52AJ:V+g#Z1@
(X_9.>Z42OOCLaEI\>CMC;7FY-fD)[9<7-G=:(KNC?ZDcQ.f&Ec=BPRH0B,23#C&
NQ?O:GHF7(8[R5UbZX0/+,1b#MFQVJ7<?Q5W0KgVFNC,>DZKN,AaXCC?V41.Q3&H
7))-YSSaWb:H\2+:Q3aO_;+a>]8CJYcc+@LSJ)?T.SU9_X^?41P+-,YPgYYXK/Cg
[Z7\;gMK-^(Z4TTTC6EG).L]1;gIA+e/g&/7R_7]NH>[>bQecV3/\Tb?,.(GY=39
7:ICd_]6]-2]]ffUKgbRMMSF^Y>/7,@>7]Ta_=S8A,G)HZYgR6T&1/\=E],K9\X/
@X5Zgb-CgB]+7CLdM^8)H>154>Z#b1Nf6<E9IcQ4P=Z(YWXW]Q7(5FdbZ(I1XWPf
_@3K&85ORK):-#Ib6[2d(Y1W^/\FZKZNDc^1RKO8,MDOX=#54))E0]_.MLaWRC][
FSN?:P]+MJYH[Q>R\8-3/OgF2.)eaVO0HB=W/OTeJ?HU@U;/I+OPgN-\4QGcU(#G
:c?]bAeD>Ye&]4W/[KSMJg-f47D_/VI14P@WF^c1,\NF9H((d.(;Ya^IY=Z?B=6E
XV\]G/=^T#eHN7P(S=H5&ED?U&EM^8_74_9G31QE\(I3GW[9bFcYQ)0beb.=?DDK
a#<7Fg0&1T4Q2T4aXZ/Q:5dK7Y_:V++02X,A,E=aFKP<UTD([Yb_6+X:(8Y3b:T:
cT<YDRY97&W4_+0PM^RZ([FE(J)5J;3RLH).\7.ddX7B32-87TA^(O)VE(;^B+6V
;B7ITDaRZD/:=]XQeS92c5S(.5M1<T)?<0Od4<5;]JFC4=T)FQO2[E<b6O2MVS&[
fM#3[B1cE=9g6>-5[V4,eb)G8&:=9WEC;Qd/H0#ZL&:S@K55=]E&<PF@R>A9bB-^
)W.BEaF[SIdK67JcJB58P5O<U;8Sc4B-D5C/6HV=1,Za.\J,Y?]LTW-ZWV_R2IeZ
NO[4<e,-AgG(0,OWSH]80V]1?f+C/U8]=4?9SNW#cDQNM@&WX9Z4)Ng=SaHSZV[E
a[V/d[OB+Sc;cUZ=2L38=]_J[\3A55gIYPdKOg\-<?Q:3^Qfd0(8ETQCUcVG9OHA
:S\U8>S/)R]1bMb&9f9Z&cR?8IJME.BCCQ?W4S1ZSW-/YK5EfR:Rf9T<22E>00](
,?INR^DF,+MdB^b5_;P8TL<GO&dDCQN0bK5RBSRc+?[cJD-O6V?cfS_d=?NO#=8)
BLdZg?ffgK,X,_0Q:W1cD(30:4>-FZX53)JbA:cWVEL)bJ2LOKJPaT+9BN^Y2/aZ
>26&O3d?D,IP1+Cb^(b^SOIcE3YUcAeU+O_0,BN[1FK07^@eW@^]1^<>RZCG?CIT
O.[D?Q8NO;@a:L9A2Q_QU<YIAKgaO#\K4:]g&O>5MA)TGb_?eNV8/Z)<&(L?OD0C
/B-1?Y;VJVY[dNEL?^9=F4M5+0?7@41<>9Y0Q)3)/6:MQ#bTPCC^^01&bU^.Z]RA
&KQXEL<fK@Wc&#?;:V<=O8IbT,f^XJNJ)E5,2TTZ_J8/LV<LFQMT#3.(=#:>S(NM
K9WP5^YfDS7>Z+=M=9,>+M<U\W=N4Y,IKH[,_O[ZU,B>JM(ON,CZR0?JMT9eE0G=
N?9/L1?^NQ>4B,YZM>L+3EPKUO6af\KfB;O<9RBIUYK5_\;V<c6]dY#Ve>EI)\Z.
SY6V(aW^IgF2>Kac5\N@RV=:eX[PC9&\G73;&VPZH58R:#2MV+K)LSb.#C/ed-X6
+O_G#-VS1g,.BS5C#D/c,\1>#[RHT.8G>BHQ33]:9c-7V,S0L&1EL^ba2TTeg4.Z
=5@F5@/G-96N(+e=/L+>PGTTJ.8P,52BQGXFT#B4:YRW.&\0,cI;)Ab2OGMZ[;c0
)>EB0RTQVJE2f5/Q]>g]4J/P@Q,,)Z)>>:;4b/:628K7c6-+^LE-2XLS_>HCLRRB
<1]6=/)1FQ5IcD2efd)L9(_7a74fNLAcTR)WKAY.CT>&7)H-2CbX+)68E;eINYX&
ZYI7NBY85<[+6d=?XQ&VLW<;c@/#_P#c&_JJL<d(2#>PX-C\@/@78dA<[g1dfg#1
-=]+JIQ:VM8gZI&W@(0S(/E;O]EY<G<a;Z)1K/IKXH)^g3K,(_>H)d_0[424b^@>
5Q^KHC3O.Lbe&LT=@4X_4e0K=F,9AD//aJGV&eNNGXcQ(d9[A._I\?CKJgHMA_+S
HM8Ycb_PFf;8d\MQMFL7OaRVWHfNdPgA#&<Jc5Y,G8e@OZd:6:SL<1H=BZ>/E^KE
V<#aRRS>baI?bTKK(?1\>BA)fUHTfMe-F9D,dB6dSB>.,fNF:UK4-=U\9QPE2)/7
cW<.fR?6XYV1TNO4CFGH\.XR-P2F3/9\50Q2I4&S9S+:M>CL;UU[JQ3;UMNOaYe#
9#@[&J&]+GT6L(+;M^2PSVVX:bb(5>5CW:aNAdSVUQ14(CE97.5ZQT<baU+f_?75
266&T]U&LP3>K[bSD^HLWe/V^4e:O0WgL3@Df0N]R)XBP[&:JGAQ7N<T9RM]FMb0
M1H.Te@J@aE:Ha,.BO5ABCY6H9XS3[/-9<[)ZV\B[e;W/@;#[e:f:RTGV+VA959=
H7c.@T&a5P28GBAbMfdbN(AO[9\FGW=G\Z\RF4K^:4SFZXM7_BD/Va:[/@@C5XN2
Oc6I]J7YP;fAIL3<a-g=VVF-HQH(gUXN;5BCU?+LC@c93T@KKO2eMG(?\I,@R[E+
5NeR7E1?K=)U3T-,EH7HX.^<Z[CfL8d16^PGcN/A(-c>C<L(LQW3IeDXA8ZGLAc&
EU.1]bG,:)/#LURUUUHDa7,>B5#<>ceY@FK<.L1+eE4S7Dc)N?dK4]eC#^9f.e[g
[P-3>f3B=.;\4Q><gF+>a?<),=cG0Id4<Ac8<[_X)@_2#b]^3dLe^K<bd@ZJ9.A/
bF8,]T0;=>Dg0@/E:XOcGRAH7LK4OF?d;Z<cJYaHIBPC<IH=HKO+>@f0/\ee66#T
Mc^++IOT]bP?,;cD\IbXFPWg-2^Vff4Y^D&WNJXK+4Tcb^SVZ;R[b0SOHfbFY+&A
I<6KL3;(C[66ggK@:Ya0027^JTa>WCN&P3M+:_B=bL#T\M?OR2cE_)LAYMAX+6;E
Tg:IcX&@YF@f&QPXG3WTfIHIJ^?YYFd0]Q^EcUJLSfR2e2TZMZcOPR\\SYL8>,06
e0(b(C4\70UbFcRd^-32\5M=_5J_dcf9-W@Y3,M1V]JVfQ4^;3T\eF7=DgOeU5UI
f(-fMP)5F/+#=AO,Z<;8WeSKA.N6&-BQX_+D.IHbFCM7(#KgZ1.2FWe3?6;F+=Y6
dE_=X5LJe?>/JTY#0e&He+eQbSHL#bQbECHQQeQdV)5bZG^LZ4U8^[a^(cX.T_06
VGQMYK^=?-:OVfV.U[4-M(.=Rb(,O;bUfB@\:?N^X[(),#:;aEZ)46&0+DGe^dd2
M11fbcUURB]&0N,dZ:UBM:WaEMV6.eI&J_+,S3AFgS^6:IK?de;.Y@6GP+W\-IO3
HBZPZFEf2B1LJdbJ0O_R;Hf1(]Cd@<>A/OB2]=dUY-fVES-\PCK2.e,eg[^8fGYK
#&T<KR#a,545O6&<ZMD_6APa]fOW<K2>L5V1b]ROV3:HCa1#WA.AfGU.e06RRT=&
7]>4d:1gdS9YKO[3c<2Q2#FQN2XTQ[.@7/X++^H5.RDGD\LJDH<&HbNaVVPfaV@2
E)]Q2D>WW-K)5;2>/;[G=&C=H)[A,b@,(O;^cg]U3UW_BQIW<-\Z=4+S:-E6TcXR
a@B.>(BT4;VNO_#PIC@Z=D35#2E0fM^0R_266#VMXJD5T@cIU4d,7?3FOB(;d:NO
A6XS8F]#&L62.O\)H)P?]HK#FH9^3_f@fb:3Vf)#;f0bDUYHW@JC@\>(dJNaDOcf
W+PZc[US?(,gI73L:KW;fW(UPeP+WYQ)FGRQVH6>(DY-FV54[FegQG1T@d#J=CW8
^A1??aJ/B@XD@Xa03S?Q,5D#NKYbROc[(ZgeV+5CMV^ceHZ@+ZV+#:RDb=8.=E(P
CS=;+_:f7V:RE:)[fMfQfZecX2R.NJ#T<J4[e.8>CF;TI[(/GaGPJ#Y;VcR:T9NF
(N3c)&H(K)#.,NG,]b.I.^60Pb:3BdNQDMc9c/([W=G4HJDa[,T:>[Oee3VG(9Ee
D)JPFFBGfMQc0J/I(O(4f>2@3HUJDe>SO5QN:GUS_K20gLZ[\<Y-dcZeTd9(UMb\
-TI0W?dcK;g>7OV]cbB5ed-fc;(26LVGIF.51NE7Y1P77)0I=107<^HJKM5J(DX6
EIe(bXfBT^=ICGe8CVT&K#.:4.AD3+6J2VYcNO)WUW-:]3YNAFM)-f76TAN_D4BP
;Y;?1gXY]_Va^3aPbS2U,g_SS+;0L9I8L_Ddg;\IfgAR@+)YDJ2DO11dDQEJ?M](
Z\FB#\X8;\ZP-1f-IX2@WDVE_;Ec8UKE]>eO08.1R:fEFPZ[A8=RAJN7DS#^FY>P
VJ,U7\KPAb>.EH^ZD1B]QUdJa4I(;Y[)8]fNWVb#V<]=#\B=Ud/VSA+R3&Kc273B
2PMU2X8FYR7N4?2RLEU=2aI^3McPKa783LT+EDRPSF?-.@HD?QUL?/MbdOJMd?_E
JB(3aYIS)V&?XcZZY00LY[1dG@.(@QX^a/W1-+S0MYE>0E(I.d^)@M#WLCfS]VaD
XY<\EVCJ5^WOUZD++73^8P+<=?(RSN/<0JW1^8J_7\b2,=X#0FCT7E7^AZ,[I:4f
Z7<,9K?I9bWA-DPB=DMPZDN8?1B4Ld-Z/eY9)Z6FA_>>DIG3eUa_XID@3X96G#TU
f#>4KQ^)c,DeKC8YM;/>_4.[eQT2W@M@L4];K>7])WT3&2>(eMWCIV;d/IP4&=PH
]a#@FTKU1fAK;ITYB<?O2V5fOVGS6E>M(VL^2K/TgS7P4HD@G,):W\V7]c6b=09e
Ze6<a?]Q:1&d>8ZX)#XSFNTeE^LWaf_J2H?</.[KNH))c;f0Z#EG&-;9G>\15^Xb
UaeKO>1WeN:(LY0WHdD(EecgG;)7B-[M/J4)\WQK\&Gf[5A/T9.J5N#E9d-,:GJL
<P&b:<=21V]&aa<Jc/G:fJ4>:)V<RR)<#?\?:<PDZEU?]B@2f.GdLe_g</3G,W(=
H-@XMKU(7#DFFLAFD_3?OL>BG#Ib/]P7P5-ZfIaGY5JZf)Qbe;?WVT=M)CTX6<7K
]d@d865UMU5=XXN\Qb?UeI6.Q+6VN.eQ2)4W<=-M?8Ud;50L?9J#WXR;Mg?7[&Fc
S)E-[C:;@81+81H3;IFe]3T+M<cQ;;4Hcd=R11VNA&,V6@eP9MB&48@aIA6WBb2e
b&0J3WdJEOfd0Q-9dRYUII0W&8#/,DAgIL2<41CXL--JN&QRIS9WEGVXIYDZE7_L
0^?EXB9S]8?4^4dP;@gL8[VO_^#A;J]W2&0TA,R64WJc82]DS#?@=P_QUQ.JGQf1
&H(cNFgS<=43N57(Y:VDZN:L-6]4[cP^#XJPDRWPMT0N/[dD]P;UH80G>.W7\062
S&KaK,+/#\3Q\.VU;FWS\DVO-H2[4-7YWe&D0@AYW\<A4W@^);M)24U]:EO82e_M
VL1WbVU&BLH>7)9)a&&.(8EB>Te:MJ]W_P)@6^VH]OU[48<873OEIaSCIU>aWI\7
,Qb:Q3P^3c5[d\JJ#-&I;TXLdN_7=/T66C<?bHdT8?E2[&eT/L@S5)13,TL6@]8c
(2BP&M;FZ4g\\N)cA-XE185L]=Baf[X+D_FH^-^D[AQA?5<18X\QA?-^^.bK;MAf
^E+Da7IaU_N;0Kd]1<^G,:T6Sa^VNgMPYcHcA#I39gU[)7&EF5Za+eS^_6(HKAYP
O9a6g8d#J(@6OR?+ddgdF\Z8eBg?/a[-[7e[6KC4b+J_V?(=VT?90(<CC0/_)_e]
(Mf<5KO/ac-R31H@dRC+KMdOYP7GKO\]>U:P)QVaLA9I6&>A2U/9\2acCd?g4IZP
UXgEe3;d_-_Ca4#@RMY?RZJ.?@Qd.KaICR^480-DSHXTa4?Vb#b:A(6?G.b;Q??e
H\->;&F6_b0d&J7MXXG_=9M6FN0JI:,#6.&<W-Ab.UFYEf^/,>D./9WB:6MSGN-U
A#X(]82.BGPXNdc/0-e2O[J302(-gSM.N>:3.&]aZ9Y.@EO-J])FYQCKca@e<Y^D
\=_=.4/aW^;C+FF7L#>.Tdc97].7&7S4^(7F&QX[=/02EK;6G>/ZGIMH-=O=6?QH
C_VGD9L=;geD,0_F?ZWO9LQ=(3DG?a/+;L_Va;Z\3R_2DeM7V4+AR+<bC@9SA(/d
N2fQ=RfD;M\&gHaNCYV(Mf3g>W3b9ba381aQ3cNQ+dS+dJJW[_5a(_fU(3H^K>4(
US&<@dI>Z5V:,P13;V4_U^eKR/YXB^O<+a,,e-K7N,[@+AO^?efSe??9LU5PJSaK
3KDRc&)>DJZ(>H4BOUcI-PW3(5R4OXIf3JAO9,=<^+K=Z7?F05^Cbe9Z.IH/]&/E
[M_S_Me5ZZb,5J]c3W@4C:Q89d_9U.2R)1<aC]0Za>8NN4Wb8,2@V_UFFEZ07;SL
&0db#V@d&FKSNd&AN,5DK/ObMd)SZC0)UXOaae[JMOBg[1Gb3#fKN_:5LQN),SKR
TA+I7#M&8AU24WZfcY3QG?YV<JebA)Q5LKAgD:>JHV.b;1[J[c;;Hf7-5d&L1[VP
,]U7P:#,/eUEK-f3F?ZMUHV+D<>7\@VJASJYHaQ>><<QOG>Y=WfEP[c&8e)HMM)A
G#T&<[JH5W(/.1HWfRWF:G+^?GDL7J>]e,2eOL28@-??SFQDc7WK;)26dQJJ=NcE
X18KN0S,+;dXA)=:>b=FF(R;.e@3N>5IfHb3fH&=N6\;FH:TNH9F<E42/O.=]H3Z
6_<PGEJ5:KUU2QXSKA;&YS[OE:F5W6@Zb(Z[06QS[.H#;D4+E&A^]C(QD;@I(4GV
BUPB8\64&d-4-F4T56B:eOd+D>Df9@eN98I\ZA#@YNGBCJ;^IMb\NP[=,RV<7N#[
d,eD5)1-?aHBe7.3E:S)ebFJ3:(=R<eSJ(3<8GJZY3?.;f[_UN6dTQU2W]<eF/0G
^1H>&d30)8:+BYHD5O.Q_C,W]YZ>BO@Pb0B^ODSaS;NX12BE8Cd?\SK@0CaH4KTe
>,Q9,U)[GLX:H(O^AMg;IL9\<](5).<U(Q[2MP(HBZ2(\VSMU#.AV8FSdc/(cgd.
(RDH<I8(eS/EgKgNH38,8S]2&7)c@&A@#<HW;W1UOcS\MOZ]5=/U&6&S]CJf\O=N
7N:?dPOD6.D#@E1V>;&#fJWEQ7JOEFb<41J\Z\A__<A+DB3<2.V9Z8U<4WI.^<-a
DGWIGK34SZ#,0>/9@PZe)S5K;/.@c1VTS71AcMNfVC=gb_B8VYAeS8Y\CVe_W_<.
VS1f&6:@_4=SU89Re7Qg]E?Ig_W;3g1JPA8F3f.Z6:41@CP5XMUdZ>UD=ZX:Lbf,
cM]KCd]U;.DQ,P4Z/VM&g=.U[5WSY[_.SMFf?)<CN@b-;[?cX(C4V0GP+D7@0bN2
aDVV:POVe6:)^a\LI,G/2gJIaVJR5HYR93;,:T^8H@a7ZVEX_d5S1a451FMSf=<D
ZBRLDeNKC3Z,/?c<W)5NL<M&.F=d_e_K3Ad5:\GKROM^Y55>QW/DA27D>&&T@SBC
&.(KWP?],F^7dN?G^YCgDPC)[][9NZ?8A-G1O,gS9[9\BeHaFM>gCKC#^d<9)&7C
KE/6BeE97a\SBV=W:0PD=^QB;S?I@gG);(GDRJ])FF6WL?\L(F+SH^?1DIBY?U>O
bK6M2e75/\c=-81F&BG6CX1S9?CFV]_WO.c]M72[/B/9OHXAG9#>6XNUDUL<3S[a
1LQQ\)UEgAUH>aaX/92II0:;/_[P3:e+eDIPLJ7[9F?-Nd0,);V[d4>\&EYdfWXL
5[BB&4/F5-N7gB73QANG)C1_(Hb:/LV@HV9W6<f.95@3L,X^&b5&_6aaV_O.:J[U
^ZUFIH--;D-(Y59)C4I+POgK&<5T9]UUTB5)7(#,PAC2N\QJLb7DG/BXX.YWUBBM
CMa7=MZ.:Z13>I@ec4W1X\fV3J>F7_H59:IA7IY+2_GMBI:#MP8(16(e]X#@YLZ2
7d/KdQ#7T5&&]>D]&ZFfMLS3(VC8@H;3Mf5O(I,^@KJ.&-bJI\XTZ_S^^e88g?21
g//VRP=Qf5D2,]-11D9cN4/#MfZa+U\_Z?[Mb1g8GJ7HQQ^H6&)8:UY7)]9R+aKc
KK_84LW1N+X^_]23N<d84)I7K&_XC\_,W36W-gaS-Y7X+M.f>aTB62VRAK+eJ@[?
gBE@&.0)8NT4cR-QE<=adKV>P.=S]E1\OAdFG=4dI3SZB+^0B&YZK-U_QL1HFK&&
[cS?T+ceJK?>+ELbSFN?>bf&R;0566>9Db<^(7SMVN/.AB8G0,M,&LB;)We>Y^<V
=Yc)67,Y9@_O(GK7NQHHLN1;&R/83JSfW)BT<MR@d++aA)4F]5X/QPZ;_#ZE[XO.
QCBI-BSGTK7M88P]=AM_+(YPPTB8.b6D-a.a.ESO>]IJF:]4b,J4+&fKY?844550
F[VcUBgaDF16g/U0R--?VD@4a::K:X209b77._,+;dKHZH>T,bZQ+UXa:fd0.CGZ
f.#P@]=_S10>.^L#)@eX##PT7FbgE44BWBZRS(2N.(c4/LVD_DN\/RaBMaY]2Vaa
B/e6?JB;,GfN7:?-4I>c6V]@<W5G/1QL_a;2+_YJ\;A=c(-?&4)[G6Q,2OWQ8fN8
ac\QN\ALO>V[Y?\/XOR_8G&<T1KE+-)c,V9:3\.+?CK:2RVF9Z(]/)XA[/7F0Ldb
]\?8[ZM8IH3I#5c<7VHTe3ZLV8],-S7((N_4F-8T40KVeAL9:g9P#F?-eVfJSP[(
\[BgY5gPJbUT?13QBOH0A)OY@1HII1QeJ\a,<Y8U[PbGBQ\cRT&IVJ#PS5WF(gY-
U_b92=T7VD0>&=d[ag-b)KVP_2V+V+B,.E/QCYCf>2W,/Cd>PKSBUR1;+),D>,#]
KZ[:I-cgG<@[FZVI\CB,)GM+L2E(=\H0]]-32bW^(8]gMg_@a<Y4OEC+VU\N+=9T
#[<QV&=JP=/c?0Q;;eR-0SI]C3)_L6]B4ZQ7)4fAIB/eT0&G]E\Ug5\B@>^HNaE[
4:Z^-gdeI9U3H,X=B-aD-8f1KT)+B3UM,e7g7@=TLL876@d+SS6YdZWV3Y0;R94)
;I<I4/U1;KKdJ/=M==Va)gLP[FG/BLJ<6;<Q3E,Q.-VFSaK;M/\;?VaZ@D7RCT7Y
_]cdB0OO@a1b7Ta0[/cL<VDd2ODT3<66D5)6XGJRV@Lcd3X/a\J5G[.\ZB@Q;]G1
d=\M>@fYVR)Y=Z>G5Z3g4?EdUF:LN_EP]C/,8f\60<>cE7MDY&eGZ>eBB0>f-#=U
;2\P(=,=b@I(6f#egC<PV]?cfR0FE<:DO8I6MA;cS;ADS(R)N;)5]cSVPH:?R(,F
,?Og1IN71-1K>FEUbHf2ZBf4,P[f^DO2SX0CNcE_LY?DIb>K(8A1VH@ZNR=115Q@
d_ef^e\3[HW+[998KL+3@A#77?D<0AXI1Je3O?.Pc2#KG38?WQ,Qg.gb3A(7B2Zd
8d;-XU3Y:M3-Z?c(.F.B60F;DS8f/(U+3VO>b>+KB&>2AZLN.KW#D;L,=AO0aZ0X
T[T@YDQ0cRbZ9C.=K&@[5R,J@0ZG+,(Ga\17#A9/YJbaCB1IcPB+98RV#Y1A051\
)+VM>-4^L5^=&^PU_\@>bI8\[7=(@(SF^STF)FZI&70]9e_Y;c+VHbH0#UQ#)@)#
^d9gN23><19;L:CNN4:RE<@M<I@^37-D3+gL]@g,_AcCTS&&W9?^+cb5+DcaLb[(
-[[RS[+[7MY[-C3DgW058+PI1#LI4QO(+_W;SFQ?V^Ze:B@0BT+;a^\M.A>g2#&4
CTX]1=OX8e)H5cf?WIJHYS0KKgefJe]&YNNZ)00C/(Xc&f&f<[TfO[=?LE_(a_J^
[&ZGf=5OT26@?;3]JG#V)fD0J\5f=<-:V:.>#Y=H^fOAKY##3AYNCBff@&I+MOA(
HL2=REO:;4RXM7?H^GM:N<c6@S,)LLZ&_1>^GOIK@#J7<10MV_3SK;TI&ACIJ([0
OXWC\/AdOM5R9E>_<_E,_7#?SQSf]-R/:TP?4@TSL/00b8K)[Q02JJe#Q)4Jea/9
G>(+P>O==BSd6SG[ZW2IALTO?JLe7?EeYJMfLT3?.VRD_[UH5)8)@\VFFZ9-TSDF
O=0_PH?7N2WFNDVF3#DE.3)>M^9>GdBM\MY:Q0\:FAPK+A#&YM1[]S#)dF]MKJIb
Ke7DN916SQ11AaZ#IR37QUdeG[8gIY8JNUe8-Me.#L:=,6V3KJ/FFbbeY5/HL@TE
RQ&JRaX3KKJK,\6RSdBN?W3&=3)QR,+gaDXAdG;X<<.44_=0L@YL8=U)>_dTZ,?<
HB6)^^\b4cJ_,=f7(-A1DFB#S@32M8D)3C9/RF(B\M:\[;aU98;-6E.D]]6_4eV<
@9]\W^P.]U8T7LVJe:;a1@MbFKfM)5)#;Y36dVa=g.RA/EC,P>HB9cC[b2IUH]L#
Ca5S#U)-8K,2Q?DPOC]E2VP.1d7,C5Y/aCgca(_g@OV=2M0:cW(1AYPWgc1DQ/GA
FIePDXYcWU0ZD]J;V?_d-C7MVXM72M(>W#V1eUZW.U>I+DNQ_TBX<_9/eRJ5gZ^A
GVHd>[HJ7:e?E<S2U_#;M/9^b=&Y\dEBJg?O(#>L<DT2S3FVK2C.LC4K:6K5d2,2
6U@@MI)R<gJBZO5RdF,N-EKBU+4X;_AZNEU0g84>S4D4.U<A-^\)J_?JGV0dZ6[:
(J2F;Y>A:EYP/0]XaBGC64J.NS4g^6fGXSBHU<Z]VOJXCT7@/>QR9FRgW7aJaBU:
I_W/P.9HTEO26SMFBa[+;[3e#@P@OF5+faTD3(\\GL;Xd#gHR,2[XBEeB+DCfIU:
,4(e7-GW3DRV7P/ZE&&@8.IH9W-0&<1(P75@VDMfS:64VMTd3K1;,47KCbd#SJYf
P\V^3<.T(OYH^GG#fdg1Ud,F=RA@K4>,,eT;cZ^7RcY@E-A+I8S_-8a5ZBAe(?-4
e60ZE.P=+c?CATUXX@B?0PaUFEEX/.g#3BW1]1RBgD(\AR@39[UZHKcK.2<ZN2R-
DAHLUD7Ff-EgA++GfJMVZ5770ECVA1<8MRe?06TK/5cec+HKdDffHT3IX?RcG_Q>
7JQ.KbO4P=MH&PTa(gA#0:B-2O?g08a3,W)<1P66QUTCdMER9[0CL&W0\^2?7eB&
WCORc4VVf-=BK<:_aLYR((Y0TWK-;B1cB^#UJ,QeLO3\@LFXWc-P4^->89be)T)G
FW+c[S3QA.d>4ZN>-@DBC5FS#FU>\OgH-&>(+Yd\,bWB1@<YHMLEL\K(W(#&2dTD
)E2?>CadVL9DEGPa2^?Q[(dE7B<,/Z;[QQG)d:O.A-0#+]d+:H-@,@CPULO:D1O[
+LSQQd+A7RC\RaM@0L0SY)A=g]g\ZD(3,D(>ge^#Q;+Nd_8D43GI:2>a\>Q#WBQU
Icg<PI25H@GLE.]I0C@83&60.0_#.2Z5Fg^2ef4/[+^?T9Q?>O_FP,(&U&\;a_C=
2;+=d:L0(HS0BfY]HHI6D--[8_H,+cZ>XMG=4N0ZADH-YP+(ZPeYUcZB28^dc>UR
&;YaT&6W=4fPY9O3NH1B1,]7K_9@dJOJX64NGCM)8BVE_81SfCgI^QP9e)]VX(aL
WFSB=(U<CJ/fd.[TKDc9Xd-LFU9F5)9KYTL]-c62M+87.4g]Oac)(@b7g\bK-)T[
;I(bg.?)(^8bV;Ke=3P4W4W-:,)0-=9&O+:Q#)60KA&QQS]UN,IM+NA:+AMX^YcG
1-B(+Y8,]9LPe>1K,G[L43B&;,A2+4U\Sg4+<e++;1S&)AURKGRG6DS@XKa?JJ2,
=AYIQ7#NScY2/SHf?<^ARQ@bcMV#PT0+<4O3gYWc;2[\]&1OU-Z62D#^()gYK=9a
NYQ]X#6?VbI]+OT<WZUbP5J=;)2>gX/+.OTUCC+beBF8ZJ;O_2G11,gcJBBG[6F2
VI(F;-AN<19f5\1BMZ8__SFd8\UHD3>7L97?+]Jde?55bB#^BbfNE-OgFb#@K13P
)K#X&ZIc+4;\@)IV,P^V4+a>3_O4?_,3bd\NZgT)^<G025@g1ET/Y1.P-M-X)ReC
>+E8P:4D9)8QN9\8(I;;D=)eKe&f@M(JVG(FH:L?XZF;8a)2HIKA5^NOF>>G+;YR
^T:J,+A<+)Ke3N(ZYe[P-4JcQORU8H0@7#9H;AO-cT4(S@GCR<Q/I0Kca&&d1-5,
8#&1^N?IMS5^>\Y3;K26OK9R,KRg\Y5G_TQU=W=+OA&7(9S?D426]gc;fR(J5UIa
^Ya]./YE@?D0E5J0/]a?^\dKNc30c3A>-8gdFM@YJ\_FfO>gS:@&K#g-7b=U(=41
;8;cAdN+>K3D6B:#V_UAE)=D4/V6SCcO)EgKDGW.4FQF(-#P90^J4J8f@B#NPU7]
S[3S90R4^MVIK[D<]T.1(289Q=>YFa(VEUKJc,4cf,d>E1R8<C8H.MB#-M+T[1L/
ID#&b=LD8R+(LTT.K6CDZK4>VI_<b/Hb(JID4IXJ@GE(A4<?S=+K8VZ=8FCTJOHQ
07#dF[Vcf>^#(T+Y1?R@:PP;D-73_._=#?.OIaP&?QOU/3PGZXBL(2PN(CDY>^;5
(9_d56O:IS=-eCe?P)6-QAgH5G&[;ZJd_5M_+Z]A4,^Y8:PaDTZ5=bOFGTbb8eE0
2/_A.VZ:GYdIU=5,/T.65ZGF85(gW\&+FS7C.Z3DL\M@/;_2ZT4M=g=SQ?A@JOIJ
P@V;d_+C>-]<D#_ZfU_8]\V3Y8=6>/K1.?Pc\E=LUc>1Y8XJG(#8Y261&RB&&.P/
d_3RV^^:P=QVJS0I;DMTfNOa)Y6=B[4?WS/a;RZS3K3&T]3,\WMX1=(88N.81ee1
]R,3[(T=JX/YUMB@PN,A&LRP+C((RC>RMEZ<C:P0)LP=a4USJgZ;Abf+S_HCbO#)
&:a2&/:fLegF\V:./c(c:A9Y3G84\?-CA<M>L3?b_-S^BdRD/?^c:W]T56^&1<+[
T#>3N2e+5>3g1)KO=#bHA+LY[+;D]JB>MPE;@LF<RD\UWgDOX?:aHS/1ag6KQ+;M
f0YZ1YQ9M=K-Nb?YTAf+A2K,23U]OY#/AW0ABccD.6&W20e;4&R9>05J\T>fg(>)
-cdNDM^aPg^4>Ga95Z:CO8EbCBgNfY9T9B>;bRRd.93ZfI>5Z4S3Z9F;<D3,0IXZ
MAJRH]=4b8Oa:R:c7&VXQQeOGcZH0@W4S:]baX9QdK:?+E(/CYf66GgH\S[RGM37
?5+F/1O>G;aEU:[LCdB8>A=O)?P3YaGPa?B4BX1K#X=C<U1GQOeOFIY+#-_KdX=4
)4#ScH;-HHI:4<3YZ(0&E6e,4(Ue[c=C@F-aNe4/SA#48BV\2JdY+6;E2AL,3M^M
NR9ce+],D<<E.XZVUc##L-+TNI43KUH8F;X8Q(f@E_RXDg8\\300U\ETb:?>=QYX
/].^MGf/<0OfHT?4Z.SA)f9IOCV90<9UcbZb[#L.JBgcH=UJWTUM&<c5K)AbK/Nd
PL^,&-3HE]e9FH.2-&2BJ),UW-X=98cNT02Ce);g^MPW+]O@FALY4YK)EXOXcCJN
0.VY#YH&T(IFUgfB&V7LBFM=Y=WU3\R=(PV>5GQQFQ/a?LW>2#_.H[cPbeDOG=L9
@2_;3PU_#J0[85K_)5M@Z7Z=@Z0IXa6+05JNdS28MD43190U.H;)WJY?d7_9Q,6&
T(?RcB9I:-G4.#G#f_HKX0XCR_[bOV\?GI\b)gW6:14F#c.7A04)1JZ2RgeLgA+P
b27;AI5PW@7FS785KbgN]=,0>E<H.S9]:DT(SU>F;J-c:gQQWT-IPU&P4L;eSRY,
2K9IWDAP@5R7/@00=^ZW4(S2/7dW6LeQ2GL54_^\XG\LfUe+f@,L?-^5ae93B.4^
K^EA?A2H.58cHgZYF6D&^HE8=8P<\;+6e4H^M#2dV+a(GBA1H(OY(Be.#Ae4bV0G
QRY6aWA?eIc-#/2ZJ8K?)2<A[66UKf5eQ,;Td(2IaO#1:e#dRf+TR>E\>T54-]dJ
GAY]c^#F029F_Q4>f<9,5#cE\bT.EQQV>$
`endprotected


// -----------------------------------------------------------------------------
// -----------------------------------------------------------------------------
function string svt_axi_slave_agent::get_requester_name();
  // If the source_requester_name is configured to a non-default value, then
  // return that as the requester_name, if not return the name of the agent
  if (cfg.source_requester_name != "" && cfg.source_requester_name != "mon_axi_mss") 
    get_requester_name = cfg.source_requester_name;
  else
    get_requester_name = get_name();
endfunction

`endif // GUARD_SVT_AXI_SLAVE_AGENT_SV
