
`ifndef GUARD_SVT_APB_CHECKER_SV
`define GUARD_SVT_APB_CHECKER_SV

/**
 * Class declaration of each of the error check stats instances using the
 * `SVT_ERR_CHECK_STATS_COV_EXTENDED_CLASS_DECL(stats_name) MACRO.
 *
 * Each call of the MACRO would declare an extended "svt_err_check_stats_cov.sv" class
 * named as "svt_err_check_stats_cov_<stats_name>".
 */
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
CMnnmuziiiGkzlJXTb3PnYjnvbfWXC23tuc89AwST1VVM6DRS3MZ6621XWDMdpDe
6t+fCdfmv4lDHno5uzmCQhAL0qIPrcJ2xYZ4wO7HDXqR+sQ0d4pslkzO56mzx17n
VHlxX4ASsdj2k164ntHxFx2YKZk8DXYZPywDgGyS5Ao=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 2155      )
3L90br3lcKLjHuS2hdOqeEL+T2oCcRceLXgkUIIeJkpIgzNzjvkJPBYUbxvvxcM+
4jpIopQxUtvWyvNyhvb0cwyDEBkDQ/tDweiOKdL/hN0kez6XxGHh21HhQUabzXIk
nsoLeYVzHbSwAr6QTqbu4A4Ckm0+oJtabWSw8AtgmbOgGODF8yDP0YNqIr52Tq90
l3NyfCb8q9SVpPqkrJfySe5cE9KpZpCbztIwj7CKzjwcPczwHIdZYVhtZy9yWVIU
oA2uXnnvKUj8iCJ+YNGIK36e9jpHa4e68kxP1gWpnrdWCfeKSWObF30YihGuNhVI
/DMxVFWMPty72CVOWM0zMqB+XazwyRfC64nfVwoAzh+1sNLFHxwCIqozX5LqwfC9
xxNo+KDcJvv9ONu/fYyvYEeijD9rdORgumgpX557XPiTvWN1NQl7yH8/8sJB1+Av
NaO+JIZI/gn3h0xkFM9laJd/oRDpCiMraC7aZFD+6LRa08uoIZAVSHvlEhhprz97
HngwI9Uwz9RW0/wIM+vHQ4poBFw8T+usFOTZ75iCxwGL5KCB+5Ad557BXQv7MClj
mUbrY6grO1FrXulmlkcqdXV9TZg3HDq/h4cRDKPvSwG5fPaI6CO6bBfpzwXxUg+z
ax9dEj976WSt1aAtFSUaeYqXlNwMKGl3qgyHRP950msbxTvyu0tdRpCw8zE392Oh
nrzBdEMZt2tQ1cS/R5GVwtZETiUrsAzcabMWQYzgOe38rmBQu1HWVUYsFissw1nm
l9jvV5vZ5RC7tBElewlRpcsavCHHrOLbaUhRec8p5hi8zwsZZn3CzB90z5T//HBo
eFUyM8uTNkP+1mT9jtqV5DT3UQeMLTkn2rMZl6eo+ziDLI3Qoo8H85vd2NrU4c77
apIF0FFJFcKJDKH1Z6KBSf+UhkCElfk9C1U3dk0J6blJ3Fs2uwN0PjPq+1dftHgW
7+RPlZ3ttljoeFreHZo/tph0A0owuvS8H+sgiqKo7ubRv7eHpKPg0tDNNTX9YdAa
vJ0HRpenUrCO7ImgyMjmoygGHutSgJgjShdFo7DAUPr7wVhdUORh3MMuMCQq4wgb
q55kIAQRbll2dIRxjn5/KvHc5jWzccOuX8tUVLVVmL+DKp11/E2rjQ3iFOfhqqWC
m8PztRkIO0GDHKLkXeQ6z6A2uYxmAi0opgv1nJuQ/19w4pmrIfnDRaC0uu05my+R
XnTtilEWK+iyJlETFhP8C+L7oe8NN0xMMGPQjMOCpamRhq5S/hwi84pt0lOdlRNj
jobSkAbDa2k5JfB7uBJP93nuD/Lg3lyjufs7bLxXuR/MwgZdrIiLD4tYDzpby3a/
xoFz/YPZqzcgFCWGvqKKUdpBGerOOaZzyFZKc1gefetZVD++CKq2M9clcoYLqoXy
sbdPsytR/W+MKDY+m06J8F3SkJzj+z1Y8Qjt/XEsJ0dQAWTr2uaB1h7GPtd1sH8p
w5tUGRZ3nAk6alpnnbaEY7i8UD8FCi3DkmC6PxCINWYJZ2Q4jZ8L+SgjHjMZBl1I
lxSRjN2nozYoWpY9MF/9YqMsi6hOGny7w/fqD4tnAAziG5TummHj0pfocdp2JouI
atvrEvsr31Tj6Azs0caWIxSSSLXRC1MCjH7ctRQdc4xJ4LFucOmtaVEpol0V3GcR
mMcb1oeroRuNsxkbuqzIMflh/CAhkZXESKhLaQmBcYhR8frOph42Sk+2r+6gh1Oe
Gibfgov3Ekw4YwRcIfI33bQSSMkHwEI744Iy8N3Xi5+AkC5NduYl9i/jZ+E1A+8B
Ub2X88pOBm4YYSRLL9zXfyqtf8bZctd51fB+PTiZ7KGuTTKkKabg5lrQ4QKGgHdh
/1kU3nE6HgDPi28klOck2owIBij6XpBS28XNml2ZMHWKXCR7TrytxZyNLSK37EWY
SQomBtBQ4cXThS39Ug+QkzK2vxvvlzFGLfxeLz98eIft5Gsthyc10oimCA7RwHUl
zYy5QE+yrax4SMIGrRQMue5+3iiDKs+eoJw/72imAQf6IVutgrHi2Tlo0ywh47aM
9HSCMcB5cxy4ltUGMwkMm1dt0WiQmT75qk17GZTJF880ddKT8n69hzsabwr3WhJU
VM5Aq9CkKieV5LWtsyYh6KD903GYwfT+qft4w/+OrXZjRsLOJAIOFLGHitCwJ0p2
bcPjNCrFt99YR2C/BsrVVBB/sJBcGyZln2pH3QYQ0Zs9g6EOP1cQN/+SE3giDw4a
SkqeXKN0CvpJGKwbW0L9hh7YJnirVIQZSXyvyQ/iqQRcnqDbzxKuHcKA8UQo/Wca
Z5Iu4XsM7N1casAbRXPQekrwYKFZi5k6c52IRasJheLn4ZyY+LbHauJK0TSDmbjS
y7hFJSVZR6KUSK+zHg1tjUEI8yMDWI91B3M/48qh9oM0CMY5Ygo6VbLVG4idijYl
taF1XnQzT3t88k33yN6ORAbJsStyqwTy9X9d0Leqa2xs39Xo9yC8UmmW94Oo9Ouu
c9hpCAPHg2AQMnMF/5bLgutgMeEObzSPTK5ofiPCqjGU1q5N40b5lzDkaaTIacI3
Cqe/GzUPvBgOC4GZzPYzkfHVKKl0mXVo1Xeaw8RwLXR/FKHWzBco9quUfu910+j8
UZ+ONtJzaSSeBh/x1wCZbsXVrwKh4DOb6W1MtVX2dKDnnLGWqTrgg7UdxfKJU1P3
MRDKkRGMBMxh1gMBFtqzU926XMq8x0MGTGv+NeiZjVMhdcRjgT/7k5BC+tV9dY5o
BRuSs84rVTec0TGX4MDmbenfJGy3Q8cGGFKEyTIH3ab7P2I+XaImlYhlc5ki5a5t
hbnN9Gt9VxUpqLndcsbwxwF2rgM0jFgiN3pLvrntG8peKbXV29Kyw2SqTjYuPkwf
`pragma protect end_protected

class svt_apb_checker extends svt_err_check;

  // ****************************************************************************
  // Public Data
  // ****************************************************************************
 
   
  /** Checks that PREADY signal is asserted by slave within timeout period
   * slave_pready_timeout 
   * Group: APB3
   * Default severity: ERROR
   */
  svt_err_check_stats pready_timeout_check;
 
  /** Checks that penable is asserted one cycle after psel
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats penable_after_psel;

//--------------------------------------------------------------
 /** Checks that pstrb is low for READ transfer
   *
   * Group: APB4
   * Default severity: ERROR
   */ 
  svt_err_check_stats pstrb_low_for_read;
  
//--------------------------------------------------------------
 /** Checks that after reset deaasertion, APB Bus is in either IDLE or SETUP State.
   * This check will fire if APB BUS is in ACCESS State after reset deassertion
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats initial_bus_state_after_reset;

//--------------------------------------------------------------
  /** Checks that following APB control signals do not change during IDLE state:
    * - PADDR
    * - PWRITE
    * - PSTRB (when svt_apb_system_configuration::apb4_enable is set to 1)
    * - PPROT (when svt_apb_system_configuration::apb4_enable is set to 1)
    * - PWDATA
    * .
    * Group: APB3
    * Default severity: WARNING
    * Note that this check is performed by passive Master when 
    * PSEL[svt_apb_system_configuration::num_slaves-1:0] is 0.
   */
  svt_err_check_stats control_signals_changed_during_idle_check;

 //--------------------------------------------------------------
 /** Checks if psel changed value during transfer
   * 
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats psel_changed_during_transfer;

  /** Checks if paddr changed value during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats paddr_changed_during_transfer;

  /** Checks if pwrite changed value during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats pwrite_changed_during_transfer;

  /** Checks if pwdata changed value during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats pwdata_changed_during_transfer;

  /** Checks if pstrb changed value during transfer
   *
   * Group: APB4
   * Default severity: ERROR
   */
  svt_err_check_stats pstrb_changed_during_transfer;

  /** Checks if pprot changed value during transfer
   *
   * Group: APB4
   * Default severity: ERROR
   */
  svt_err_check_stats pprot_changed_during_transfer;

  /** Checks if multiple select signals asserted during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats multiple_select_signals_active_during_transfer;

  /** Checks that bus remains in ENABLE state for one clock cycle in APB2
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats bus_in_enable_state_for_one_clock;
//--------------------------------------------------------------
  /** Checks that if illegal state transition occured from idle to access
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats idle_to_access;

  /** Checks that if illegal state transition occured from setup to idle
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats setup_to_idle;

  /** Checks that if illegal state transition occured from access to access in APB2. In APB3 state
   * transition from access to access is valid transition.
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats access_to_access;

  /** Checks that if illegal state transition occured from setup to setup
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats setup_to_setup;

  /** Checks that PSEL is not X or Z   */
  svt_err_check_stats signal_valid_psel_check;

  /** Checks that PADDR is not X or Z   */
  svt_err_check_stats signal_valid_paddr_check;

  /** Checks that PWRITE is not X or Z   */
  svt_err_check_stats signal_valid_pwrite_check;

  /** Checks that PENABLE is not X or Z   */
  svt_err_check_stats signal_valid_penable_check;

 /** Checks that PWDATA is not X or Z   */
  svt_err_check_stats signal_valid_pwdata_check;

  /** Checks that PRDATA is not X or Z   */
  svt_err_check_stats signal_valid_prdata_check;

  /** Checks that PREADY is not X or Z   */
  svt_err_check_stats signal_valid_pready_check;

  /** Checks that PSLVERR is not X or Z   */
  svt_err_check_stats signal_valid_pslverr_check;

  /** Checks that PSTRB is not X or Z   */
  svt_err_check_stats signal_valid_pstrb_check;

  /** Checks that PPROT is not X or Z   */
  svt_err_check_stats signal_valid_pprot_check;

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
/** @cond PRIVATE */
  local svt_apb_system_configuration cfg;

  /** Instance name */
  local string inst_name;

  /** String used in macros */
  local string macro_str = "";
/** @endcond */

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   *
   * @param name Checker name
   *
   * @param cfg Required argument used to set (copy data into) cfg.
   */
    extern function new (string name, svt_apb_system_configuration cfg);
`else
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   *
   * @param name Checker name
   *
   * @param cfg Required argument used to set (copy data into) cfg.
   */
  extern function new (string name, svt_apb_system_configuration cfg);
 `endif

  extern function void perform_read_signal_level_checks(
                                                         ref logic[`SVT_APB_MAX_DATA_WIDTH-1:0]  observed_prdata,
                                                         ref logic                             observed_pready,
                                                         ref logic                             observed_pslverr,
                                                         ref logic[`SVT_APB_MAX_NUM_SLAVES-1:0]       observed_psel,
                                                         ref logic[`SVT_APB_MAX_ADDR_WIDTH-1:0]          observed_paddr,
                                                         ref logic                                    observed_pwrite,
                                                         ref logic                                    observed_penable,
                                                         ref logic [((`SVT_APB_MAX_DATA_WIDTH/8)-1):0]  observed_pstrb,
                                                         ref logic [2:0]                              observed_pprot,
                                                         output bit is_prdata_valid,
                                                         output bit is_pready_valid,
                                                         output bit is_pslverr_valid,
                                                         output bit is_psel_valid,
                                                         output bit is_paddr_valid,
                                                         output bit is_pwrite_valid,
                                                         output bit is_penable_valid,
                                                         output bit is_pstrb_valid,
                                                         output bit is_pprot_valid
                                                       );

  extern function void perform_write_signal_level_checks(
                                                          ref logic[`SVT_APB_MAX_NUM_SLAVES-1:0]       observed_psel,
                                                          ref logic[`SVT_APB_MAX_ADDR_WIDTH-1:0]          observed_paddr,
                                                          ref logic                                    observed_pwrite,
                                                          ref logic                                    observed_penable,
                                                          ref logic                                    observed_pready,
                                                          ref logic                                    observed_pslverr,
                                                          ref logic[`SVT_APB_MAX_DATA_WIDTH-1:0]         observed_pwdata,
                                                          ref logic [((`SVT_APB_MAX_DATA_WIDTH/8)-1):0]  observed_pstrb,
                                                          ref logic [2:0]                              observed_pprot,
                                                          output bit is_psel_valid,
                                                          output bit is_paddr_valid,
                                                          output bit is_pwrite_valid,
                                                          output bit is_penable_valid,
                                                          output bit is_pready_valid,
                                                          output bit is_pslverr_valid,
                                                          output bit is_pwdata_valid,
                                                          output bit is_pstrb_valid,
                                                          output bit is_pprot_valid
                                                        );
endclass

//----------------------------------------------------------------

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Yp8VcVGuwy6A//dp9CoUFYeyFhez1wYSMqF5LW1HyzI8MXl53zIWxWK/bGtsC76W
nscqYpQuo9BEUdptmQ3bdnxsG/rtwdllNLd43yOe97IxBW3MizPZ2WsSrN1oxpRr
gMrPfWO69vOwuGX2qMooT2q8oU2RFVFOwQ9v5C2WAwM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 8926      )
sjA72G6+5LRwTBhI3kTEplyEGfvnd0yLlh991FO9VTTLLSvxrwWg1Sjca5yDSbDn
7lezIiVBQ+IusUM9xd6gknBS/BCgaU2AZ9n1mGZ0FIMLajscpYD/2iji8Byo5IAr
43nk77X0ZQYCS39W3rYFbuf/U/tP2MrXUlQvttfWzEAaoKq4ZfGJnZx2dH50S+ef
Rm5vrg6aBRruo9T5gXnPb61pPXYVNg9omHYmHnxio/Us72bYLHBQ9PlzSAcOYN8y
IAM00Omw89nGcaeEzh5QN5khFoVM/bkU7GTFaSCashzWABthag8p8aXw6efSwMn4
S0idOCBXCU5CBYFq+5nfAAkWd+KDES71tDNIK17cvXamUyD93AUqUZwLHpO5jwaP
erxWL9OD6daULzhSL6H6A0iIBujea3iGh4KdjQf36XdXT5ncBN0V4W+vuYsWHFiU
6/RunPErYxHuVlhLDEU5sx9A6N837izd9FNo8dPlBDkknJU72JleqwlD/Aq1FHi0
9wVlm0EOtItEYKoxoSl5uCw5aqthKEUW+/V4zDWtFwIWheUkfaR2nQJmjOb0p8Wl
rsV7F68xUDCV8V48NZ0UwOo1cRQJkFHXkmioOq+Fr8737BI0KS/1KGRqRe3BeI0h
qc+59Zu/3QiigiZxVDDZdAqYy8+WVudHURoq5ZjHJLA+1IqzD2AxFvJ0IknpGswa
WjmLi2zH1FNant/tzCk80UjL67AfGA/H2f9/eYG3Cm2zZgIIQaQkS0lIQZu2Rrg+
1CC3GiEzff07FMc3qlHjABBP7MyAiy/NHnUjDTMJnMXv1pU7vTTClYwmQIiWvzLC
G3r1HihAptPKHXG0IxVAJTHhCf5x4yxErf6tge9ALZYAqsZ+Y/UYEGY9lJEnpF7B
LusWBSNp0kmUwSE+WJPmyVx28+z09DFJgv6OETyn9EhKfDlAOOoxujGFJXOYW3kK
m1b2iV9WIlXM2rTddAlrLPWc6zjTvTjMmyLRbQivzgRVUT7jSZH5DZPfQNFU4d6r
2HB7T1oV6QZEIP9A5wO39QGzoFbBD0f31lCQz8UYdjtkXn+pQsrC00hVAxs+j820
whTgUxwVlfdzXIdygv6s1vEf3XhghKzUj5lvzZh/JR1EMRzfmyHHcBlovxLZV+Kd
7yx/R2xNKxEeJcdFH8M9Xr4JTfVVMEA8PiNBysL9MjYCDNEV801/C63x/NlSdEqn
uHTRSz8qtgCnBVsXrx+sJITqAB11UHLI+7+2Ts5cGUG2mDXH5LQpseik3OjNWU3u
OCHs+hi5oIW52TQ98spYsSxh7Aoi1gmJsXvGNoUpno/fjlpHqrWiihMSZxx6hAJt
WhLMwsLJoosOOW8J4kddPxHzeZcDgSv0pGuKmTbPYVwr7Gh7B4aK6NqlAHC3ALko
AXqYu+xoZwh4FpkL/DwEmQvvxSj9WMZrz+3ZQjMKqyxK9NgR8X18xeIFiPsvxPjJ
2V8OnlcvjhBMXcyzMM7WlByxo9qsEvqMP/HUzTeLLUaKZ7TJqzGlXbVD5mDGConv
3A5Zs9smOAla76dnRzGrxSraqaVPlU+XJe7s5tILhRDhi7L1pHdGA0PXXlkIXaIv
zrxT3HycxOcW/OJsY5uypKmrbghTc8olBWY8uXvBOsiDZ9Gc7bqJZo7yNwH4pM9K
ftVrlkYIzzt9Qgdmgsr+80DvI4O8C+R3NHwroiJ7Ml9sOeE4/gMw8C6BhIcXUYz9
4v0WipcOb4bDPvBZ24w6B0XiPXgLvfOndHFPdRPQ5/T22T1mOvyKt+hbmq3iDvve
d9bK3PPE0ojWK6MIcvr/7IO+P+UGcDbEHIc4/kjsYLRZKWJsxdRhEM0HvW++RWku
HS88wAkqsbpNesEZ1C0w8tc7M15slcVOL5m9qzI9cKRrXftmv7qB+PxAeiDliCp1
M8gatEneMdk5vqAPSdJGauY8Y6QF+SwoM0Hw41PoU78QvLIFaKCl6CNjifpDiW4g
CjAP70mSJKtvbcpfxsTw7XHIAh9mC6YDIpmiTbQ+xXaPXd2fc/Lrqqc45mi1xS0t
Ze/oUccPA+MDRHqfkF+wizODGNnK17qRFzTJgd7m4QtJUXZmx3E+vIzysn4Jn7+R
4EJhvVonJk8zaJuJayRAROho4QKcMVUuFOK9t9Ncnfb+uRT+Yn5iFZrw/0u5/FVF
DxG7seI8VJBHBazgrOY1HA1AZrWGBQ7L8lqrycUrZecd7oZ1miwqUnzJ6unNQeWa
BwrahDjbnb4qJ671/ewfPp0aMnSqALMLJA+4y1gktLp4EIQ3aq+zjwLtxNQGcNnL
dBNbXqjgXvAzn5XPkl/1yp+aS8+EqKuv5zKrrXsCtHa9RnOBcpbuH1U+ffKWnT7Y
PT8SuYVAFoTrlg6j6zxpvPCsYzEm3pIuLVGZcQRvNN0EN+v//B81VnZ+zSkHhRja
BoiYbzWDZb46edM2CAeLHu6tLR2/mMyWJ/0SGn4x8X3mU7KlWyBx7CwfwjKw61s8
VLkP2gtyrUQ4uyk6braFHSM29CGwCKj0cbmgIFEfFxz7qhviuQSvl7/Pd9PJILyf
CgU1smfQ4aLskOyziBlimIR/bk+u3fqLDYip+c4/A1yJ2LKZkWyzir4EJ2i69zFI
YFIbaUPAd/RRFNRqwpwXjru1q9+C9z8Iu76lpE+hxPe7FEUm9pb4srmxZT9PxomW
GFxf3qx/N/hsth+PU9oP/e2HLXxvS+nND3uoz9hY2rTZeIg0/vnoVjT2efVOr5tb
zfvIVKtxSyee5pHPtIbT/cn8YQhlgwA7OLbv8TEe0hViJ7T8EQxLtlAcbtSqzvxO
8oMsVhTCRkXew4Bx0MEBGSB/BiC2m/ZyaKqDw3MxGEu3LWiLmk5SfWt4z/8buZmu
gkn+c9MuQ3xl6K1wFKbAOpAIGmmsZIg0g8scDUfl6JfTtNYlK4I51L7hn5ppsGK3
lsjKy5z4XYE/rWrZH9KxeYnFPXaInWTmnY8BVGmixiATc60H3PYSL7pGTOkLEWI6
2nHtnnPqHBCiMVuLP/peE8JDUv30tMMMAh5H/YENIa6fol6MFg9VF4oImEk9HRHD
udb8Cq7ZI9N+uvygcm6Fi+5Y7j/IEbZjTuSNBlKEQ8I7hj8VTJolBNM2CHU+Aw5f
mkPoj9h5ddrmdRPJhThr4MskK4yaAPNRogiNz1Dn0L/6JI+R0GQIlwgCsGS4+LxR
GRmW8cZlKLxe1L+zi9qTbifPofBZIZAB/B8ssO+VZfRcUByWEWuw2mX921K9wc6t
cOggWfxUnjRT1IllEK7XJKSF9VDc6Bw5eXbuMT29ywL8PfOOpBscyv7dRKi/Z6xs
+tV1uEvLHGkicylX/+3fXVJypP571wJ7heg0TlbQLDTcRtoegr1I6TtpSTTebWWa
5MjPbzkK/cKEtuUcxzdhJsAbpTirn1KCF9l8PI7aWhIRVz4OMAqafJWUjWrCQHun
7mg8tv1ilKvWzO0DiR62h8vKFDk3coeBjfCLG9v8/RbkHjfh+NrRqDee1kSMsGpL
LvlOY3hTkCG9LqtWSRiWurU/oEvBwYWMJy6DzN5TNMIRx8H7zQwAAh2vcpie768k
t6trQdnp82Q6s+Enoced0IczBrPRBz7TfEjxpXJoPgZKm0KfW9FaW2xOxaUVeXvg
ywnDjdFFYaiP1mk22FhGjfYGiViK5dk89bUPRcQjjs0O/7bfhHPGPg0Doq5AEax0
leHaV8DtyIk7ZRdIm3/2lai0bQCvSqcSCgC9z2FvVmJjgl2YVAwdnR2iDZYYQD6m
Vmwd4do8JusK3QlzyCAFyX2DZhtmox7jxWQ+JghWWOI59Dldrq7/MkZ8D7+j0SeC
Vx1UOLEXHnJeGZ6lbrjO+uOZPpvNgv8lPFUYusuyBU9QUqactdrqYSFS+RXyclhl
H92DZRBE8yM1BrciwMlCtVPOklzNIJMRNuwNRxxRFC4VfXcdYpT3VSwkV9N4G+Im
mMmxYwZK+FRXNtDta3jRAk+4c/Y7lkuegPCzQy1I1/rEJ52uHJ8oPvBqRAdygNZC
aGpoXvFHwU3/XeOSx8vHLs7ZwicZ5dLH5qOyh7eSDspemjgNusk7mtiYJGHnNWK3
EHf5Clt1nKLAzR7/KzbqRYPszBce09qAt+DIk85PdxsXPm7bA9mdej4JW0MFJy9v
JAL1GKyZU+2LHojAVcazGf6qp0WeWlbCf4eBraAhK++430Ua2Twa2Pcb11mUKxni
1CybhytnC6slfVVktChljwstg5itEmTnozHfK3RXy2nCxSxofQkWu0wpZXxPXwOq
BYRhUg2XZXuW5Egl6rHBuKQM+od6m1zkTWNQUVadFCOu9LE9eBQ4FFJJE430GT3L
34JNRYuPD9ZJnQ0+61CXt3tQKZUXSGBpnTE6Sijfw083Uz1nWVAmbte/shCfItNX
7BVbaEm3+Bf0s+gd67Ro9CK4ktGUnwuHS7NyyHapGyutwJd8b7q7RQwWuISDAGw5
JT8q/aK5E/oH+bYHVoUbVe34oQnytn92GPxyo5L5bV8ZLaOHZiDviBGx3A6q5RLQ
d9Z3gejJXmUu3ct2AGrjnSYujkXndmrwkPX/2DhEuqYWDZ3A7z3ymuGoSdsieuih
uHVTzrYbggxESZD00mDDnCaObagLsIGPUmWlz0FfoY7F5W+V2l2tkFAPCoyp7Qhz
AIIL/NLVLh9lEXWm1B/fkDQLXfcVSDRqbbvcC/aFLQuKMdcI3zsMSFbTgBOcIfYp
MHi1BdEmvLz8OfE4j+XfidxB6eh+CY6igGLoLDuVnqsP6fJDVmJARmfiNH9th7x5
AxcuAbIgrdH13lJcBYDvSdUXfw+nqXVcFpKT/TXR0u1zHf/kHG74elMx4NUPWd1d
mdJDln8XPilILrsiZkAyHkg/5XIZLGQoczLYSSSI7ZM7pP5nO+LG8TBhXO/vHHhk
0sPwL9kApuCpet441OnxEXbO4DRbJJqwoZpsrqO2xF9pIn71qkJhosYX0eBJaZ3I
I8PVQ3XnAMDr81h44bSVUzMnNjpOow8GPvw6MF7JajUKTobP9OGgK0fOAtoLXXTg
UlBs4v7WXAOJj72zoVTiEs3HHyYyH1AvzJTDIWggUWn6exdSfwvR0dH33QL3oGWL
yLGuOW5KKFtPYCQN0eThg95olK1Jsfx2HXB/ehjd+tTsiBv22ShT2X+ab6xNmTxl
HeeV8WRaAIjGVNzfYXXNI3VCjrxd8S5ih7dWEftzP+ugB+P2kN4h+5RM/SjIIea5
8+56IVJHW0aGRQnbqSkAGWrMJyW5LfAuioXe2Q8jYZyra+V1w2Rgx+cNrq2o8NpR
D8ZP+zEoxhkE7IrHH7z/0nVLj9vK+ORSSi2MpnFLehuSuCrYHwcr5p74Q2M6/vfE
kI4uEulPSiFPuZUxKq5yf4IUiOkYFtoWxIeU5jHEQwdBFx2czb8DmOHd7TUGlacq
sQxYuVFG2gPxDFPL8s/FHlqk9xqYlXOC/78KXu6MfCfpE7yYkX68bs38mH/YWFf1
67sU2/9Dd/6qmVzmZks+0q4kbWhAQ9S2Uc/P8R3JnHpdwgJoLl828h+03PO3LGN3
AaZAA7Gf7wyNEp3fpzwlGopSbFVKM2W3hhe2eBJ8u85wRH2nSBNPfpSTmTkg46pw
sc35vPNxbO9VwABR6deb/lYxdoqOlrVR6uwCr3O7b6rTXmmHMVMk44NCYQnuw+zB
rVe/q/mHaZjEf6ExIigc8Cx5dqWQ8PN4/0jBwV+pjn+vsQw0IHik1vU6uj4Xg8Gx
+WHOoFNoUC3hIMEpRnoC7ouBbLsKO9DYSRxPSrF3Jk/g8aOZhuOXhcEZB6cxGDyA
vzn9ltcxorf5SxzTTl29iRImexwSiaL+oMCFkqQRNmb35yKEi6rq0vrPw3unfgpb
KaeN1IZvv2JWePfXp361vNEDFgQp0ri2ygUpbvWRTBRHqC7sXaSFVvSFFSI1FPW+
yU36gyGsi1LG8EfF7Po5FbG7ogGx/C6qsHJkr5HOpgXAoEVfnhuckX7wCEN7Kczh
/qBE2z2PyeY0mGogYkE0WcDH6tLsbjzLGdFTafp0o92wVybKfyo0svaMMnMh3OA/
KIwun6u7LA0JQ2cWjkrpGHAbFisIBt8SkV0FzemIe8CZuRFSUBVuTSW6pWoVa7Gh
kCYgesMbS3JW1IgWy4YQPQ54FsD7ITyI/FQ8z1ruoIANn6pudNRl8QoW/jjtr6qa
+fNXIWEui3W6k00cZeT5Ahuc/TTZBle0laAOfjtjiV/Ib7pBZzGxRAhIqQYwgUJ/
GnxA3ibFVoD0tntLeTlbWWLiHRZkjgHeZ+VWriZ1nfalouMk1em9p976cEMVRlMj
kd9u/ugJX9BTJ+hxRRqTzHRJKLsJWEgCVrl6r1pFWcUduo4fTNFL8iY4x9QzHPwO
Z+xgUMncHc1qK4db/+srLaHF1O1z3Uw48rE9sEHFdw7qmzFj3cIm236aXAYdyd/j
YLxdt+q+9bIGWnyw4sBc7XD1ojU9Z1jF6kwCshV6o5lvHIrgeSCx60Jz4lvZtro3
gAtLF55xt+P26k3LYWLOVc7afWmYMme3Soj/zesVV91rbr4ssqMMNMqK80pbMubH
nYenjWhOfFMpofnXvizvoIdPCXW+OjevsTItzVx55LiU29CokS3bWcz0VNaYbrxU
v5VL0C42kDPVYl/hF1fHxZE6SJMj1ts4O1RjY6Jm4FTsRmOXRxuXSVYYzgKvxyCg
q7A7fhOgtcOoOiuECs0X5jjJVZdy8nq9SadV1cTlqe/Qjl4M24mXlzKksDGQKOF7
RyROtRKpiB6zAgsyMUEIk8J1e39JDYvxcwaHmRARzs3u8MB6V+NwJN1sgZkSOHNp
Coi89VxPiPaANGFeci5QE+blfoPVQjcOyu0U82JbJqC8klkjiZQpgVP3IgHK0Az4
f3BZ/cCFugOuKNUpQkB8onNdzxaHNVPRP0ZojkBt37JRNEWoccmnCPRlsZ6aOYEb
ImFi9h2RiigV5lBTonKCzxl/e+3+naz3EDHhw7Os3Yj0x4+VoHVxmOwjTWYkjqE0
6b0olvndVCPYtqJGCiwgzYimL4v/ToEYKsZXBErYbUcA6lOIGFL7E4KLjmR0MCzX
HaLFAfcftliNDLHwZQQRQTXbctE7X1NRIK+thHLO9VxLsk2zjg2Cn4ndVTuDZABz
5blUkYSLT1yMlps2mA+GfcnKGpByk9wMytRvdJ56irMlltWLFYWlbp4+U347pdJF
mRdgfU6p+hlkZ8uvpwa7ctJj/bJ757GUoA0QR9dqywyJ0eRfSnQKYnhrDzPSq/nT
T6hx+BXmjx5ZlGtk/vPm7RBdUSajXuQg2S1iXLRKDsrqTraCQG/Ve0s2oxCXceeu
6oE1INtDUDwJPaOHfGQ7TR664qL4rH8VTei/NjZlQujKuUWg/NxvFVlBZRjwGA+r
nVZT3D3ptfBrf++/1m/cfx4X3nAUg8j9pQsc1qo7EzIdq/AcKFnOHZCp0rbfJSsk
NcDmTRvlmMKVopvuk+Ws1T0kSkQwNgGPfHQwjx5I3igukqRprCPc0u5Vjm34w4sx
UQCk/3dlPCyLw11v6/ffSX5xEWi+DnKRyh1VxqUiG1Sg9EF2491VY/QYCTSWrKXq
LKDKZm/Cy4q48HNPPaDdQu9q5WEfUpZZoHQgEhkAQvQoHLyrwz5EpBQ2mn4WSrLu
gvUbAiCZt9OB6l2+Wgcdx4X5IkyEKT5L4qAyFPSWEHUgUhFEV+CE1VDvCoe+p7Q2
6m4Oio6R3vq2aIy7XJ/VqGBPsLhtImTCnHKGy1jvxgwJB1EH0W1Wo6+0ZrhzG7cK
ngouflIhDyBqHB2fhZQVn9/4vHCmnLm26SO5htUjcT1F5CCzxVfdBSF50Da0dw4d
v2LQEQANXFs9hoGLK0Sf6UjLC0OK2cJEfvq4tlm1ywX9oXwleCZ2cIPAHmVw0jKr
mL8BX66a8QHMxCYiD76LJocHDH2F1ZlVGtTu8btZyzelz17fm8G4VSXmSAj3glkS
/rPobM6nnhZlMKac1QiiIanrus3FTYLzUmwMNh0DNW7ITpAyUH5br1/Ww71SsS4v
sUuNST58XOMX0QOyG1FRuCyfZeDo7S3znfgOvkA8fgGaffuE/tDHBvdkDMQGj63m
YbjPJfeshwSoF4c6lPNXreiEpf/UjpnIRcbb745R65sz3oMNjLaRVRNMCd0GDDA/
ko7eS+fkYy+1cVDJP5p3qDX52kBBTgcr7jol/9WNQJuTYWEaMMF5dh23q0Idt7yF
pa/VO7e6F6WOxh4IsA6VldpQ2terbgBoNoSaLwen84fn65q779VJ6DXJ13t33be1
DaU0z+yvcCD9RMlil5XrQN8v5GBGtBxrxHJkdILh16iSJOOn+HD5oH0Q3wDE3U7x
qb5mZ9X1hDjkMvPhp8ha74ZVIkmA7vP3RlA2J+ilwZAIeOODQzv8Tdi3KKOrFTLX
ScchQgQAMHnc0eP8+Sm1JHdSgzymUuVcriurw2BYVKzr0ablVM/dlifYYX8bOs57
GyS3czk2l9+/nuLvIzwx/Ks1D2QBloQhc20SzshYarrVgz6+yLVPrlgLKuXdiKWy
wpro9lWdKjs/72RPJylRuzdYm4aTNKA1i81Y4AjXpDgjSDERtVM6cfeEhsRtcEod
e14E7AninpoeaucJAMxCtq7m//SdEbqMWhE5S6lzxV9ecCG+wEq0dWMtF0pHlldK
ZFWRv5nh07YZ49qRwye4NfdlBohyBymzot+Q6JfUkk6x4E1stUjO+wbapCHCiDHm
DjVjoNywdgtlrT2SoZXotgrmLECRnfWcHeEhauFzlBTERL3fPpf0QKpfS1WiL/mY
QV4z5Va1bYjV7Kwz+cBYmFhpcN2HPlWxjcQ7Hzt4G6KFgdZiGtJwSuv6n4IkjGVz
K0wHfumqGt8T4qG2sHS/sYEYZI9KHuBD3crmmk40Qz/CsC5y0uDqfl55wmC1ZH0s
j6C59JV6yIvDrlQsh3SJerJ6D3fslstOEE2o0Ov37fOINQ0Y8cU6+LNe4+tm1quk
Lt+1VK31WfJRrD1bRhr+NA==
`pragma protect end_protected

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
SAOoyHT7m5KTXGlGiGTXnqxyCix8/bMNSSh6b+C0eMegkDoJsvAo1CM1VnjDkj0J
5pHnZUpgWO6MmqAlHtTyZ1Lq+qmWewfUlCvvO/CHNOIf4tAMybJ9tV6a8pPV0fEJ
vuCN1rfcLncn0Qo06h+0a1mGHZdalexs9SYGyrmjvVI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 16731     )
QSOEcLtFnK5NahydWPnOOvGiN6O2uTcfzsbF3w3Ta53BChECzN4oucvh9JG5i0e5
0Qsl4J8TKw1yCnqy8ARoksvOtQWDshJbqr2g4rhKyPng9xUJH99CIiBzuVlWEIEx
ECoubpBK0fwxsCklETJJiE56xJ81e3UH0RokCuNMSYsKGD8OXSqllSfJWbYIHsgC
AJtMoMabf/qPJYZVsad5vaQlqzbOhr8IYbZ4Tx9+rCYVg2ALczI+Je2iWlfjWFTX
ZH7Vd8aE5buZ7SX3WHUilQNyW+kFmmY+6/86XdFtRvk7rRb/TmKET3GlUp8BJ8ea
KwRqWDr5dIDz9dLFuR/EU7o8lUt3Hc8InhzBOiafB8gQOV2sDWgPiuyCmQf/W20u
LdjBYbm3lzDduSWOPx5BF3RlKqDpX2rhzMcdVJLKGtBwuUL/pcB6kGg4QkrfjgT2
UEADkb4EUEFkNvxqoFkKyovTJNAQ/VsBuKdzYhy2d9kBrvfubrAIAgftonVYo9Aj
bNB7pgKJyZ9oXFbO4CcYngRR/JqhjpyMkfvpvqJ5poipU8bGzrIfww3RSMcuSY1w
a0cMOD6iBPe/X0jAd9v9XcepxG8Agp2kGvS3H5Sx2xoPi4VMwCySbJffsNuKRJqO
fokMmwN4kVRuLNjA4aR9hPCFoEtnbllA5gCKl1+ZFLx5caz+FimIy73X62yJrg+o
rgN4mHFgkc2uDP4BoRC6IJJNGLXcd36Nd4gf8ybZs5BATAr2Tv4WaliPz1Ex5YSA
Pp35B1FIPLjFVvFxI3YEbHhteJwKw+upGzqvjhwy9XJR0UyHrOSlsIyUfE8xYwEV
ijmEmPzBzaX5nVAr84TcifAU50MrF+dYUIcMw4CNyGBtSLzu5x2y2pDlRVmhe/+J
rEf58soGXYlB8wqfx3BXCRHMbURRtrk/alnGHMAtPq1iha5zsNJCnoatbiB74YFa
MCxPNXIfUIeOIDQ8ImiDbEHBdJQth513aCPjFh90fWGJA2cAEIhqIyzYpa5KbKfj
SNz5b0qtykes2G8sEI3hKLVCJ0Gdtfc3SXgWV7MH7iVW/sm/1ylVx6EZUMXAC5GQ
HmRQCEt0kJJbPYmVvx6WmDiNUPA5GB5YFktBS9GN/ZbIkz4hX/u5wook2ADdmN4N
4GPXRfiWYgS40gM/b8XbbLxCpCM9JwGhyPlza7TrN28nCSBxgaNMo3GAkX5Ng+U0
UG5VILOyAlSS8PfejAI/v/o8or9uIEv2BXDc3W+6rr8nJcOFm1rvYqHO2AJ44Wze
OnMZZrGJ8Le2mnUpU0LsXGR8CshGjkl3I3T9FIwlRtghb52nu9pj+FLshhY3G8Qf
G5eMkAzRKjVK6bkas7jO1eBI1MEosXiN2ABlp0f01VAty6yQssW0Fqo7ZN9abrQM
4TQJ99Y04CYZZlgPTU7LgK8mTPzGQC3P8csxRN5DX11Y2Wf2kUfZtRpsGtpysnS6
6m94FOnm79ov/pb56QE2sUX8fxlVrhPtHU4F9znvz9SwUhAMRqx5YfPiScHOJ7os
T+yBzjJnA4EnThGWfeeHw4Dwbo+m2uAPt4HXYlZ4z4OdbI5q669ahrB078rEE9C2
WklFDkxR3Bk9WnsVIg3v1yitp4uwRuMTGioRyc3EhNt56sL4LHG2yiADFt2h+f0V
vr9s8uVlttX7lMe4MLEGLfkdzmkh73zrb1SjOJdatYqNwixuyoOIoUoqcxWZqICm
5WU6NHRBwyFIWpGclX/O+Ssol7eD1WIoTznR8KhWNHRr8LTW1KTlU/LbrwcQDXZu
R9AGZcPofqQBfPW0CbV2yclCYea0uF+79b4SssN/Ye0FWDhv0QtwR0Zn/TvgX1pE
llQB+rF6WgnX/Vgt4h72y05eIUzYf/osT9x9uGsacyfw5qdQs4OKGztEIpqdCA7J
Ro0uUeDmKD53yur/FWJlJmcMRfkijjwV2d8vStgazRqCCIhJUpjYRLOG9lx+0lGp
4+ESKr1B+ocYMgrrO0MKH4TNhlhuBXCwvPgMZ1HWrkj8KA9F4CCHECKHDEZs93mF
kaV7ELRgLDi6uUqYHm4rMFkj58jWgQD4PPs+RvREPCHlFK7S8ISoBQbpBFue5FqJ
An09cH95BwaET+eQ34y+Vdq38DLphfANa6vcl9X6rd/7f5rq4Zh3cYm4VfCqek5H
O+NPyQ0PNKXR5ZKlZX8rAIIh5J4li0YNfg/BsAqnImXyU8wf/0aHC3qIFqijT1yy
WPGcrEWL2HA521eSikNGrkq9twE1Y0D1fDBkPyBOg74M8dN7XqzcJundZANt+9tM
LWdv1g7/CAXPj3Ic9gjSkqUiAYbbkpaEN/sdBfQuoW5/o6dkX+MU58FVRc6fiHR9
GRVNbYhZYIJl33y+ABhMLipePG5F/ql3KAhmImDFebe3iVF7lj2iCiJaOahtTn16
cQE5zOxgAgu7QeXwN4idKOHQfL7Y3dvStZA9snfIFMEWICoizEKZ6Ow4MYR5pt82
J2zjkVCmRwBuEWVW/Hc29HpAy6fYPQCjSb7usD2pZfE1AQtp0oYukG8Pa5b87+Uz
CW6Kqz8l0ZqFLAce9zTuTLFWqIRSGbsZQCLA6JM6US0VhPmZqFQfcRJdANJw+aAE
yGpIBRU9resU31bmALn5kDwAv+C1UtMPcApfLabUktCIVY5VNipMQs1gxQaLZM3S
PQt6vSRbzq2Ki6WhWUijPVK9SMt8ApKxDw2Qj4oyd5LhBDX1g61hsR3K4bZZrHiO
bJ70IMTmKcQdwxfRtd6HF7wFC6/yVzvvs0P15Qu4ZFImuzpRerX3LVlU+DEmzife
9HK4kJe2nXT+ZXHJtBMvSP1+3Ur0ZJd+C8KUFXSQgUV2vjxWJItDM+fBNuYdfzOP
KASo2yFOpFOtnQeiypr/xRPgNZ+s/1F30JxIc0CEX2afoMr1givLxGZlRB5sLAFk
KfXrV80bMAWBS799TOMwvVDNhoxXhizNIX5WSQlcUpp+TygP049D4UC+HE2SYIWi
cpxdx+4i8IZZeyzxTSsteWQ/gycAmmPob93f7b6KeXlMhGev4dDO8Y33I54T8kmo
fpiJj9DDPAjhWRvKb+4cJcAcKxk2/ehQgBKbZOgyySYZ/SgE0vsBdtI95VSeSDrJ
S2PfzqfPEbpnluPg4im1rQFxV3V55vBGvu4W7lM62QzsKthHgcL86Fgy4VdrPF4V
R5MlazP3n2M5ISi7pJDxH00UaOpSlrpIq0vdwS8QoDHSNY8TjecyDymN3BfInJ4F
BInxdod+u23QNx/vI8QqsDhj7QHklPUmuAJd1WheyVXcqJCV4oy1v5K7IjmnrPMZ
a5yyMWBbSDCwmg1mq8k3FBw+JoKNt2eCxyt2ms80I+hp0Ej3LLRWovEamsWZNUYb
w5iORpjbpe1OOx8PfRYBu/lKiSUF8CgeVyIP+zaR8w8SWlx3wBg923XUZ+TCP1Xn
Sq3NQQw41/STYQ3yAinPtTZK0cdh5+9iPAOGqTc3f1CG0jvEK4SGwkwCACSxmDQ2
iLRNIG3x8OTrCYuw9vgoHw7SplmixC3Z7N2zy+lbKclEaC5Teve96VbEB95gYjaf
NvvKX6jvqGewD8hDCeI2mcsz06v3ZSwfhiRfLo1Q1CpV58A4YoMWeXfNCDGbUE/2
3IjnyOuSokLgggj1S6i6g4txVhxBaeLOFTdDic8vGXTMQPgA5OstHruI99u9HOQ+
FyOMFZvLk+mbphhvTVHotaDbpKAqkzDWofwGEcUjyYJ2jei3M/4D2MZuWWM8Dr1P
gbGTLpqtip55T2YEhHdbN+RUQsxrk82/HUx1jOwThEk4qi0x9j8+Zc3dMambl1ug
O56B6yyroQT7w2jBbptBncmImMEhOY3TlBs2aug9Njlc2m/i5VdsmCTaRllkaM+f
75KZonKYpV2Fh+PIuGvsRcYLFei23SI4mPRm90xEtTHHLr1ASGQJX/UBmQGjrvXW
KrNdF1q03zx8xmW9z6ufzuefc3hzrK4j0dMriRDGpsJ06Ys8kavnkhe7Gw90VWtp
pqVAuJpjDf/TUefc7O61XDk+H0xz1dS0NMIWGmGhPzqfGlqggpvLzrX6ok19IJJZ
BYAitDlDmm57eMi1i8fd571jVFb53VYUAadTYIo1ulxm4uzW1CElU0fjK5/kCLs5
0a3QAodyi4IGQvkk/adZa50h/6004REFWiu94x0tRXDFy2UYNiB9dvPCNxLtgFMU
WUVEO8jgSbkCVkTmOcYrYbjnQI6JOl/RnlMn3BFkXB8jaUd2JnhQWt9Gh+qmENTg
1pSvvEwU18y2sPYAZfS2xisLbw1lSlgwBHfXZUuEDNZt2EalhFbYfjjvADW31+/Q
XCvLjmiNcA4ClmWj7TBOxhvan5lwg9TG+6Wf4MmO9F3yL8O9NKP9oWoGxLoGci2Q
NmZWylhdxPf3UvBYMBYPwCSOC2r2MGYCrASHQUpnxoxN5XWkn0ZfXbhZDuq/uwYI
XlSQKWlY3g/5YcOrjTK/Ce71FaMT6EWsfBi68LaRkWP6N/v4Xpw3KW4BxcM2QbE9
+rEx0dZwsqeFGrpyV1iW/aCfj7vgldjy5tehGTWrqRAkffME5dMbIbsmJoWC8Jaf
albmT9ST3OJGvLnsxSUvKemw5oKpkvDDGO2Cd8v0fv71TaljAxeoEMgEgv8RT4TB
bdpuMkaBzCfLRziFMYYBqgjVPGFn+dW2XNPt6D7N5kqUZFI2G6gjeTH0GbAX/Vek
3IF60fxrzbBtRMPa9NUp0raIDxaUqBUx7S3n3watLAnkApUoPNooAsN03CspRsiL
S4vs8tgfTYbTfn/OsnIKW7RLLxNeZ2b0wJ5+jPNwPWqUNXkpfycvefAgdE6ED1Vj
mrdnZgpJEen404iJy06un1Q0jCDCWxilXKujXRMSNHmWqrLSwdzcCm/UqQdzHeGJ
pS10ytkLKP4R/4EZuvYP1yOj+KJFH2PLTR7Oa6bS3EuCly+aLAKkCgvxrUywwmty
4eNtgJVm7k9adqQ4sDBUCVTgx4hIdttO4dfYMgR0cgLBpDJyEoEBE8pT3CqQtMFz
vVXTB1p9lF4DhZPAkAfbvfbzTWBAAAe/D0Liff8l3ZacqlXLoOJcE7u2w1o5fO9k
qOFmkGUPStLYDFq9bAdvWXtXllFwLduvV2jSAK4/6HVoKnhLTJ/P91vKvE40B+3+
PLN75Cf5vI9rtDHUY6Ek2XF51nIWz4n6fi126as5+mRuNiUr7SUu7I1t+U5zpW36
Vc9y5NAGRRLYS0EOnQkAG3KSn+F94bbU+Nu5wo6qjkXWKnuGyczKaBcQE4NgSRck
W7P/8WtywQwRW/8eYw52OIpMPxUHZxis1c7pTdN0b03Ia9eanizQXwvO4YPtZW9e
4pwi7RrgOaK/SnVT7+utIQeW2yLQYnn4AaMdis0/2wdItrqUwi/ATRGKQOoWvRPq
PAKNCVEpj6fsRgRre5/yvUBRllSlkopDFeZnC/oaS3OuCZxJheGSJcfDmlNGKYvr
TQEmQvspTjzFhve83GhbdUiYXm1LokLEMZLXVnhwCkftSIPeB6JCcXixAFV2qrLt
6mF2eXwgrxPw2XbHodqPlj7dxVCOG35K838JQbqBwlACXP1pdn1wwxjxle/nSQMy
ziFy8m2O6XOabqMFzbJSlF9VWZ5zQGLysyS/IqKBlKfRZMlE/bxupkNc9dkirvEk
pGBDv45/SHHk0eIdcL58DOL6gI+Ci49gyIg3BVP01+KAuUIejdZ+j2OnEXb1OM/W
E688gdwxiG5PvTLgfR/0FRtfAt7PfX7PuAle0YlPGHLR2jVZIHhwDhVopM9OWM3e
lV8FBy24M4QWAEnE0CMYIQeBuefhEx/Sd3U6LBzbpBZ/qXVtBSG8hhDeuii0xir1
P166wiKCTZ2yrQAblbyxG6ieeCUw/STjoSxUXm7BX0J2FX5z22qKs7mfleCYuw1F
nG3RK3eNOvRYT7iHCyx3h7bDuKCS7VT+JzddcjzQNGnOnTdagkJHGWVcHs2Any4h
qGNwPU+JVnqfV8iymNJIFvuvjt5YdaDUnj+xRqpMaSa+32CYmE9uty/vNulsA3s5
LBZTmxr/i/c2ZMRcG6u8W1RgNb9MN824eol6lN/2PqAQI1SSKJ94a/75G+ZaY8hO
DCfoI5BeqpaDr8wAwzPRstc3m6mo0q59mlXKYf4eEEVYyIphf2d6rbRDH7clcTLz
RlA+A6hRXm+jS7HiH3AJUAtuy2XF64/XtZpJOnx61gHYwaZN9nnveDqGvZV3OGNn
3v3zMpNfUstRS7KiFKvVJ4ogLSCD9TJe0JuLixHNwmrF8PVuoHCWCgykZarkzWqY
Yvt3quqNt5/7VNyZrN87ItLoIBVUIKHe6ZZKt4Syxl2lKvoaw2AGYp6FSKh71dba
NnX4KQ4FTwMGzwdfEjYKizYRi6T2X2sXXZmy7mroB2Zo6xSIxxgjS9YVZadxAjrI
2df7094djUrsXYdHIRcdD9s2x6UjoFl00qqpdEA4OwpwrWdr3eeAweXeIXpdVgp8
Ttf/XMMHgyIDD+1QlmKkIoTKdOsMXBqKARG0O1SLpaxDB88ZTfL0DeLJGu8Ekg/u
BEDpGXZz/+XSyshK1ShmXaghmCk9GJNDIvRL5DErsrzCARSlCLVKuujvsbloofgO
B9ZiSuB4PQWdCYcooRkBChw8jj6qqDF+o+LQPLxQLUsFBF4Qc+i+Xbpeg9NAJZC0
NVyplQ1tJf2rf2X/MszgNUKHzlPqPNGgXxcYBvmyHHbn66IY0GI298PWNBqkj5Nh
fJqgcktw0MBARKeYRQxOBwbkvHL/DFWvyJE4LFjzQYHx6zxKnHlx6F6pZzJc1mlK
8Sw/v7o6GtQTcaHmnjpjtyOz9uYR9yAL6gg89qwAozwvfQzQDNygGPcydYg1Q4ic
opDDHMmi2pn/6VzOAyJidFk3aSKYSK+GUTqsX61i5goLnIKbFqA55Q2VLBU38X+f
O+wOKX/jIamCcM4Ss9F+CBhUttOisUozk5HxuJeFGdKOspSSCMVwsm975acSnSYm
1ZoGBK2ejeAs4IdJetRd2dOYI0UkcvtCGRuCm4qbzNO7qOP3FxLkxf9eGed90oYw
XDoYjoTFyJfiNB4oEFhAMPbFnT0mXx/iW3Ia/i4KwttqjPhL0FsZuSNqB+R/T6g6
mqN6OYu5MxKUs/2gpjv1DSp1/sZOPzUpP2NBHYV6xARyExs4OzEtjR2bUzZbfN2V
0E9fLd6pQ9QU1yKjpzDGVyZjUCV3gsn7nY5n0XNTRWyFrBrQ6+gsgvFnJDbg5z0p
PB13ISNSXYjZbmI5KrJxjqg5YBOs/yFaMydlQGaBLTqdOB1lgrTo+e72M8cbnIFv
/22chQzfrLgPqxd/dD1Gzyh+MJzdcrnE13f42cZVyDiqss9GyOUqKQHNxeJ0GU+l
F1BDrghyBZitJtG3cQS22DuVSTaUQEmMU4NJl9cC+dsS7pqNFzJX6vZoIy6sph5P
ibJdywgnhkp84J7eFqy0srexgIVWyBQTjdwH7G+laS+cxIhQ6xgVrg1k3y7UVtvA
4bWq0BzneDKE3RfQ7+vrSPeiK6VQykGWsb1uMtYWnoeaRw/WP6JnGLZD6C7/U6m/
k4g3xHl+CqPoQKIVaylAFooedr00RpA0ZvZ0mp7zub8qh51D1CqYBHrcDlkHtAUA
Pc9gzTu1JlEM/pWrWr626sICGp00HRqBDlXnTc/NI1L2aG/7VEn2R2WRiJUjmskW
38PTrsFfqnuTdQNChay8BR2UkaH4MsdIz9g1q+qxMqYH65B55JnNB3q6g6spyt3C
B/iWKUZ+9lIFaDexi+O4pIp+S/wghg43FkKF3WXQc/ihbsm5LAOQVRSagefOTjnP
3DJijIdqhYjWP7cobBHmm9i00m9k2S2lAeydEZTnaApT77wjk0VxYUsc8HnEwNFq
o9O0th8GU73Co6KvvFEA7qRCORFz2pMqgsa/Hk4GZ+jbvmsPqoQOzpTtreIyohr1
7ZWv6drDFUAZR7Noev+vnbnFGFk8ajAPhJaHN9cC76t/lZhoNmwAjusDEuVHtwA5
P6FBC1G73TaMdAOWD2rpwmDPPad37JdamHupDhVglpL3aVZck4xWbcNjImxDhh9H
qM4TQ/+NtjUnMLiPbP9kWck6rHZ0vmcpL1Zl4XyPhs9OS/fApl2oi4m2+1kxMYl5
ja51bf9zOluoMrR6uDTGQvmllPS8OALJK09Nq8NSbPSHkEvrSaQdVFaaBF+jj+eV
l0M6SbZHvvDue+xXOXjTC2g4UtPMFbooKebwsTUxp9mBJqvmCmmXNV//1Q9D/ZiA
l89lyv3Yq8quxa6S2WGuOXwGW/b3CvHvYHfHBt7qKAKh9poFeh2yhW+K62j3mnHu
Gv8vTVoDghAOKFwQYqWaOQd1fAVBLBnLAl2A/gCYqioRPXdrUxbTyDWIhmQsH4C5
f3CkUBftNYdbgRxGGFRnzPYotTbus27n43fQboRHZj31rl3mmE797oYtlzDiP6wy
Bj+PpdQsK0NOC7HJpOUZDqG30nwmwCKodhk2fR+FZILZZtdHDJT76IJ0qQVyp/df
LJUxi/yJH9RHLxdCO9LTdyRTY4i+xYT36bh9Awt5gNQF0gFWjBc56Z/mo7uf7nyU
rbCWrIbb9gh0m6apnNEJ4am+yy4/03LRRIKEsnuBSDyYy0s6MZZZ9xuYh4Tkglfo
wmXPFqSVkZTDWZxRrOoX47zVnm8fciEhgnTlPViHpjX0OZUfjwcV8lVbqxVGmuf+
mXHhpejpJOWoOzhjJFXekyYYQccJDTJvxnsYFMSw+41+c3YQt/5hIG/HIifrvf/K
yN8MujRcyIzQ9ICpUlW1OoAISwfnjbmSMMNlLuZXIkkWwTHCLHBDFansi0Kxu4Gq
6xeSzu8d2KXvETG2zrEgoe7cfblEaUavkBvPKD4Ku+gUqWHqPDqpl6JnACefS6lF
2QZ/qeJf7PBwD4C9rAxZOVu+jI4IdVziQqR3nT3E0+K8wjqfAuk7Lw3TuQCxoZ6y
g57iobmG6zkM3+4NAhZ+Mtw0Y2PnjjwI2m+W4/7hih6ci0GmQfGh/UrOfzjZ+c6p
+khmHdyvccYXv3RN7mpBgiTNerPde+DCHBID+UQlOJ6vZ/G0XfigOiKEeuJWkIz0
kjs8/bJbYza0MDQmBBNF7Sn8xtYoPzElvq5Q+ESP56Ysw/HCaG9uhv/p/5phoniT
QqlALpYJa0aMVm/kM931t1JlGSMikat1iKG+BT/VP4EBq9qMyogzlT3HiUyLs3+e
yadTAqmZ8qqOSLm8QD9xuteiyJjSnQv77fVjSKao1YRbuCkjOP/y3PszJAvqldGx
KXJl2fwhRcVXKZ/TClMliIVbvRe49koA/5zw9tGDXei2S0pUBkRuU81YehHOMMnR
QiT43RuySb0JlqK9A6TrVhtTX9+OU01EUMYncu7L0KRU8gER061KkUqe1VRjYPOZ
09qjvg7zG1gAkJA7uP1gAG15/HOileBajTQa+7eOaJ49SHvp+c1SX+ltfCL3PdJL
sQyPtO/mcNqoSdqbuwSO9qf5DiCqxhAg3Ws/t8fv+Ke+m9uhDSwzG9Z87HzpbQhP
qIcsHvxdekmUFXdPybWzxD0I3GgJabllECGgXp6Ta3gTZqRm0IcF+13Xpk64WpRR
xDNwZeIv4H/L8MT+ao6rznUbrWhO44RJ7d81D0GbbV5viJ3HPINHjszGBAxqPFKB
RGHUmdbB+MJVh+FohU7+vt4VHDMOXh+4rfM97SEADpp5JVVgsmIuFLEnt+NLuRft
4W2SgiJk7W53mNIaAvJDsg5NH2AzF6t/PAkmPs49Flso2wm0/L9uAQE13HW4TyFC
KtghFHQCN/LpBq7yag8EqL3sR9ALt00jT5AWb0Z69CiRS2onHoaBrLdo/v2XzLdy
Kb7fE+EFFAMItPovA34YlZSY/5tH0+h6UwXCsoTphX5Y0cO43P6+zIBDhk+ZPRqp
VY8Woyh5e3sKkkTF5G4likgcYnfXbfSKyfCVbshJ/mQo5z/5ivVtIDb/m0IuWxyW
g1FeoMvp+/ZP7w+5pqX/Ftzq+o0k4GjREi6Y9KLqHQVX3kjXFbVADwzxl+70f6xX
LIGisRFKUdnRG7xP0sQSQVhwerzMiE3wxF4iRUdTa4ZGbTEGkmmGnM6I48kmgRqw
C4scdavYZEVHVeW+jqyyTcLxwzwt4ECrpSHOSyJXA3xj85FEamAQGa7jxY9sdGa2
ZncmSe7m+d11nIvIcUo0L4MCDs1VZbCyOklr5/QkjdXZwR6/8vumiEObXNGJILxR
+o6gFGq5bicQNYNcLUWEydwGhyCzZ2XMY/C+EsQl5qnxdl6N2qxR7Ki5951UM7Ww
odsvFUhLGTzu53L6maa90rrAA8dKBCkZW0W80K7dsvg=
`pragma protect end_protected

`endif // GUARD_SVT_APB_CHECKER_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
XQfQokozcLL5H2v7kyY3sgh3wsF4eCnigB9mTud7cSszDID7k9uVnsdbv3jpaR0N
I8cIsVEuM4oUKpC0QYBIzd6eo/f0LKQ/ODLS51mhAdmUAa4NZO2fL9g+IlrjJzTO
ByR8oiuL4OCL71QKpKU3H7RHXa9RtLv9YR/daJ/Bbzg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 16814     )
lc9jrWXxery6v+s43QU3bPcbrYuefqXUtBob9cfhr4RSYcWsCCuLH/Rjiixk3ieu
3e7y4Q0hb1biVNISZTcbaeWAhrfwNxRD6gCC/tw9trzLLPM2/kZlPf3WIuy+woay
`pragma protect end_protected
