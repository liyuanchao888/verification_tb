
`ifndef GUARD_SVT_ATB_SYSTEM_CONFIGURATION_SV
`define GUARD_SVT_ATB_SYSTEM_CONFIGURATION_SV

`include "svt_atb_defines.svi"

typedef class svt_atb_port_configuration;


/**
    System configuration class contains configuration information which is
    applicable across the entire ATB system. User can specify the system level
    configuration parameters through this class. User needs to provide the
    system configuration to the system subenv from the environment or the
    testcase. The system configuration mainly specifies: 
    - number of master & slave components in the system component
    - port configurations for master and slave components
    - virtual top level ATB interface 
    - address map 
    - timeout values
    .
  */
class svt_atb_system_configuration extends svt_configuration;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  /** Custom type definition for virtual ATB interface */
`ifndef __SVDOC__
  typedef virtual svt_atb_if ATB_IF;
`endif // __SVDOC__


  // ****************************************************************************
  // Public Data
  // ****************************************************************************

`ifndef __SVDOC__
  /** Modport providing the system view of the bus */
  ATB_IF atb_if;
`endif

  /**
    @grouphdr atb_generic_sys_config Generic configuration parameters
    This group contains generic attributes
    */

  /**
    @grouphdr atb_clock Clock
    This group contains attributes related to clock
    */

  /**
    @grouphdr atb_master_slave_config Master and slave port configuration
    This group contains attributes which are used to configure master and slave ports within the system
    */

  /**
    @grouphdr interconnect_config Interconnect model configuration
    This group contains attributes which are used to configure Interconnect model
    */

  /**
    @grouphdr atb_addr_map Address map
    This group contains attributes and methods which are used to configure address map
    */

  /**
    @grouphdr atb_timeout Timeout values for ATB
    This group contains attributes which are used to configure timeout values for ATB signals and transactions
    */

  /**
    @grouphdr ace_timeout Timeout values for ACE
    This group contains attributes which are used to configure timeout values for ACE signals. Please also refer to group @groupref atb_timeout for ATB timeout attributes.
    */

  /**
    @grouphdr atb_system_coverage_protocol_checks Coverage and protocol checks related configuration parameters
    This group contains attributes which are used to enable and disable system level coverage and protocol checks
    */

  /**
    * @groupname atb_generic_sys_config
    * An id that is automatically assigned to this configuration based on the
    * instance number in the svt_atb_system_configuration array in
    * svt_amba_system_cofniguration class.  Applicable when a system is created
    * using svt_amba_system_configuration and there are multiple atb systems 
    * This property must not be assigned by the user
    */ 
  int system_id = 0;

  /** 
    * @groupname atb_clock
    * This parameter indicates whether a common clock should be used
    * for all the components in the system or not.
    * When set, a common clock supplied to the top level interface 
    * is used for all the masters, slaves and interconnect in 
    * the system. This mode is to be used if all components are
    * expected to run at the same frequency.
    * When not set, the user needs to supply a clock for each of the
    * port level interfaces. This mode is useful when some components
    * need to run at a different clock frequency from other
    * components in the system.
    */
  bit common_clock_mode = 1;

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * Enables the Multi-Stream Scenario Generator
   * Configuration type: Static
   */
  bit ms_scenario_gen_enable = 0;

  /** 
   * The number of scenarios that the multi-stream generator should create.
   * Configuration type: Static
   */
  int stop_after_n_scenarios = -1;

  /** 
   * The number of instances that the multi-stream generators should create
   * Configuration type: Static
   */
  int stop_after_n_insts = -1;
`endif

`ifndef SVT_VMM_TECHNOLOGY
  /** 
    * @groupname atb_generic_sys_config
    * Enables raising and dropping of objections in the driver based on the number
    * of outstanding transactions. The VIP will raise an objection when it
    * receives a transaction in the input port of the driver and will drop the
    * objection when the transaction completes. If unset, the driver will not
    * raise any objection and complete control of objections is with the user. By
    * default, the configuration member is set, which means by default, VIP will
    * raise and drop objections.
    */
  bit manage_objections_enable = 1;
`endif

  /** 
    * @groupname interconnect_config
    * Determines if a VIP interconnect should be instantiated
    */
  bit use_interconnect = 0;

  /**
    * @groupname atb_system_coverage_protocol_checks
    * Enables system monitor and system level protocol checks
    */
  bit system_monitor_enable = 0;


`ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname atb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to UVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to UVM_HIGH or below.
    */
  bit display_summary_report = 0;
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname atb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to OVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to OVM_HIGH or below.
    */
  bit display_summary_report = 0;
`else
  /**
    * @groupname atb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to NOTE or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to DEBUG or below. 
    */
  bit display_summary_report = 0;
`endif


  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------

  /** 
    * @groupname atb_master_slave_config
    * Number of masters in the system 
    * - Min value: 1
    * - Max value: \`SVT_ATB_MAX_NUM_MASTERS
    * - Configuration type: Static 
    * .
    */
  rand int num_masters;

  /** 
    * @groupname atb_master_slave_config
    * Number of slaves in the system 
    * - Min value: 1
    * - Max value: \`SVT_ATB_MAX_NUM_SLAVES
    * - Configuration type: Static
    * .
    */
  rand int num_slaves;

  /** 
    * @groupname atb_master_slave_config
    * Array holding the configuration of all the masters in the system.
    * Size of the array is equal to svt_atb_system_configuration::num_masters.
   */
  rand svt_atb_port_configuration master_cfg[];


  /** 
    * @groupname atb_master_slave_config
    * Array holding the configuration of all the slaves in the system.
    * Size of the array is equal to svt_atb_system_configuration::num_slaves.
    */
  rand svt_atb_port_configuration slave_cfg[];

  /**
    * @groupname interconnect_config
    * Interconnect configuration
    */
  //rand svt_atb_interconnect_configuration ic_cfg;


  /**
   * @groupname atb_timeout
   * Bus inactivity is defined as the time when ATB interface remains idle.
   * A timer is started if such a condition occurs. The timer is incremented
   * by 1 every clock and is reset when there is activity on the interface.
   * If the number of clock cycles exceeds this value, an error is reported.
   * If this value is set to 0, the timer is not started.
   *
   * Configuration type: Dynamic 
   */
  int bus_inactivity_timeout = `SVT_ATB_BUS_INACTIVITY_TIMEOUT;

  /** @cond PRIVATE */


  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
 
  /**
   *  Stores the Log base 2(\`SVT_ATB_MAX_NUM_MASTERS),Used in constraints
   */
  protected int log_base_2_max_num_masters = 0;
  /** @endcond */

//vcs_vip_protect
`protected
8L).3KW=I44VbF[-XB3X8EZ=gd.2GeNU)YNT:B^/5@>f>ScbS4bN6(f>>Z@I3I];
MR2,:BD[?2PCKcb=#.Y)C:U/?#>/2[,OLfMf9+eC9UA-,8E4^^Z/DHdaJ@M073b7
V6^\KQUDIG=LRGJ+&0+->Dc\D.W^-b6O.;;AUX(f=V5\BCZ;MV#\>+TJ0>b(L.95
Nd)UDT3.=U:Y9@bYE,CFG1427+]+b2NQ&YZ&.)MA.L6L<XabbONMR]1d2W:@1F5a
f<cIGO64\fJ)_U]9GYCW(H9)@a-08FA8RHBI:&@B&e;0P,NB#4GaA\R#LA:3g3Da
=;CA4ZUA5X,W#55)&X06P<\e/Gc(A+UbX@5J#NC</aQ6OK1Rg3NWZ+CWM[UTV&,N
KK&V[HF\c2[^<2<1bTU<#1GL;b(JHN<OC4^ENY15GEDVCXL_a?.8VD_LX049^J[]
?>GXLHT4f=R[RGA72#e(/cZY,.,ERN#2<AUL/>gF]0#XDJ^055]-H9a4BUCMZ2P^
N7M_5TW2WU2+^I+3f>0.a1)XG/(#cS]^PC7Qb(5,T2WME3+B,UfAGRfSD&9@)D4Q
=)/d.Ff_]I@gN3#bERE7PU_/<5OITUf:_KB0OQ5JL=_-V,\>DB&/a+(Q[77)&VP^
13Ca@@VA)>90S4V6<-g.HMCJT\JC^bE@M&ab,\3(HRC->YXaS>)@O;>OIGbYZEAT
bIS,XQ(W[U)f+Y)-JRMD&I1_a&FBHg[8O.K4=V5G<N>aJe3==D0.Q/.MYaJYd<TN
CI:2Vde:HC+]<Y-VLV659V=5(Wca:2F>gW7KQ=DWEa0S1;aI3;:/OM77>1DA6PWa
9;d1/+R,87E;[(+D&/FHgA3VRgaLEC]YTZMT4-/HNY3+J]@2MFP8S65E)2PVOeBK
G9THU=A,Y18aGIO[/J<RV.#7GDD>01JC1?N=A+=K--H&gMK(PN+f-#EcCf(Z7\XD
K72#[#I1\J>W3gW/MaI)S7002VEYcB3C+CGfD#(#:.52@&9Y^V_F6aQKWQ3,8S,O
&AJa2=J&IId]0,4VLaD-?DQD<1e0Sa0\EAYWaY?>.-DX.1QJ7aA,KPV28X:f.6Td
X@6ILR#6Ie4U:;:VKPP.(M8__[0W0F6<Vge0X/2WBP]bHSJ1.BY.(@8E(.SKX8@,
QV3g(APdc;cN0CDDN]bV=]X.D8C[eLI=MW/AMYb=IY]32G=HKEcPaPRIaUJAGV3e
8Cb<W/()S&3B^d@ceDe#18G17LR\56_.?B+H7Ba);EBZDe5N8BQ&9&V<,ZHC>)e@
B_0U+JHQ7)7=#Ga,4Td2^)g)Z=XXFDfUGYaEU0D<M_e3URaF.=UBU4@?,U3V&+YW
/CYY8_M\#]E2-_&-<B,WJOFI<W1&6A=6:AEBf;A)<4b<g[G:V^]#8]LJER+^A9AT
QGY_f4N86Wc<>O7<6\[7.1a+H)D:QWDRT&+]3K?@aG3g4LOYZUMS5c]7F,KL8g?E
4\?L10+#LK#H-CI=a2D#fgSZ]2d-#E&=7/_:,a>ODKL0=2@AVQSZ)[,.K,dT#\&C
6UcPU\&fP((EDcJ0?T5CMQP_E(fEX)44TH;U<b7V7]WL0@O5Q1bN?M:XGXC9aNPa
C)K-UZ=WYa#FUV0DO.XVg&\)FIaWa,b\QELeHFCYX04_QIK_;CGZXA50T_,QdI=@
2Se)HYCQcgE]Z5TdMAQV.X<J+CII+,7SD<^]#D250<OOe+C20dN2I52T8e>=_GF.
O^TOYU=0:JBAY\U7,&Pb-:eW9S<>MPZ#FFWdYW_,O7Z1feE#8.Y(a[6)gEI;G]GT
9@\^eAWc,;Z\H7N2+N,R^R>;OdL,5:?gQCKfWK(SfLEV4BeWNa.A\4W++cR)JYaM
)W6a&L1gVB0-8&EC06F5VZ5(54->FYPMI@R?+BUe:BMgIeBNK,RDB#7NQH,,g^CL
;OG]=71KTZbM7)eB4=bRVCOH,,[e;[aDb0N7NE,D3=)MP9TCY<,#eBae?9d?YGNW
LdJ72&#DUS/CJWD?81Q>A@4PLF-F6RN2C0C:Ue(LEbZASPGCF8X&N9b)5b/1>.HR
KE3d:V@/TdK5+(>(^M<6L^Ia(14&6Q;J;=3g2+Ja4.T)GI#&B9-4-=ZdWdPB&(=Q
Seg^VecWSN2VA]YV#MF@b6#:TMQ;LD^>9@LR#56DL6fIJ4d6L3W4b-Q5W8fJ3.]O
57Z+:RS(H:HKZ;d<L#.,K#RHOdO.[U([f]Ra.\N6>T:O(Q]=U@-EWM/WR?N[9X6O
/&(bP7-6c\I&f+W<.[ZJ^\6:B5:-&P,3-?<_e)3+E4=Y[FT8TR4J9,=G=53@U73&
XG;N,IKaK/LH-XM,\IO>Y3W6<YLD-E[IBCf+@H:e/W+9WJBN:Wa^dfWY?[BN0cWA
A<b<@_b[HB^#a4>cSTYY=^g2=X.W+HL\\dDg/1&TBQCN32SZW[0g7\)Q-BeNCb+A
6Nf:QBf<H0K5f6eJT^9M9^^Cc5\]W/S-)]M=MA1VBK_R7P.GB>Q]H8Z9/H>ZeaF9
7AQ&OdT;X>&BY]FUHLVA.gfBHb2586X<P^/@21)S=(R9_]T.A<8E)9e(WWdg=8+;
\=,A2.R^1D,:69ULN/;1TCH_+Z@OL=MYH1451M[?T:MY;EMY4;:B_2Y-+IAc+^=4
#_1&</.G2_A1=D#YKX5^TWEc.O9\Z>JEeAH8W^c<TRI<IJ\,B0\WML#X012&L\Ic
Z8f<@;0TeW8&fHA(50NIG3G<<[1MZ&>Z<$
`endprotected
  

`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
  extern function new (string name = "svt_atb_system_configuration", ATB_IF atb_if=null);
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
  extern function new (string name = "svt_atb_system_configuration", ATB_IF atb_if=null);
`else
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param log Instance name of the log. 
    */
`svt_vmm_data_new(svt_atb_system_configuration)
  extern function new (vmm_log log = null, ATB_IF atb_if=null);
`endif

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following
   * 1) calculate the log_2 of \`SVT_ATB_MAX_NUM_MASTERS
   */
  extern function void pre_randomize ();
  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************
  `svt_data_member_begin(svt_atb_system_configuration)
    `svt_field_int         (system_id,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (common_clock_mode       ,`SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
`ifdef SVT_VMM_TECHNOLOGY
    `svt_field_int         (ms_scenario_gen_enable  ,`SVT_ALL_ON|`SVT_NOCOPY|`SVT_BIN)
    `svt_field_int         (stop_after_n_scenarios  ,`SVT_ALL_ON|`SVT_NOCOPY|`SVT_DEC)
    `svt_field_int         (stop_after_n_insts      ,`SVT_ALL_ON|`SVT_NOCOPY|`SVT_DEC)
`endif
    `svt_field_int         (num_masters             ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (num_slaves              ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (use_interconnect       ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (system_monitor_enable  ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (display_summary_report,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_array_object(master_cfg              ,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(slave_cfg               ,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    //`svt_field_object      (ic_cfg                  ,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_int         (bus_inactivity_timeout  ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
`ifndef SVT_VMM_TECHNOLOGY
    `svt_field_int         (manage_objections_enable       ,`SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
`endif
  `svt_data_member_end(svt_atb_system_configuration)

  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();

  /** Ensures that if id_width is 0, it is consistent across all ports */
  extern function void post_randomize();
  /**
   * Assigns a system interface to this configuration.
   *
   * @param atb_if Interface for the ATB system
   */
  extern function void set_if(ATB_IF atb_if);
  //----------------------------------------------------------------------------
  /**
    * Allocates the master and slave configurations before a user sets the
    * parameters.  This function is to be called if (and before) the user sets
    * the configuration parameters by setting each parameter individually and
    * not by randomizing the system configuration. 
    */
  extern function void create_sub_cfgs(int num_masters = 1, int num_slaves = 1, int num_ic_master_ports = 0, int num_ic_slave_ports = 0);
  //----------------------------------------------------------------------------

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(uvm_object rhs);

`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the OVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(ovm_object rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);

  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static 
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);

  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif
  //----------------------------------------------------------------------------
  /** Used to turn static config param randomization on/off as a block. */
  extern virtual function int static_rand_mode ( bit on_off ); 
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /**
    * Method to turn reasonable constraints on/off as a block.
    */
  extern virtual function int reasonable_constraint_mode ( bit on_off );

  /** Does a basic validation of this configuration object. */
  extern virtual function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);
  // ---------------------------------------------------------------------------

  /** @cond PRIVATE */
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  `ifdef SVT_AMBA_INTERFACE_METHOD_DISABLE
  /**
   * Function set_master_common_clock_mode allows user to specify whether a master port
   * interface should use a common clock, or a port specific clock.
   *
   * @param mode If set to 1, common clock mode is selected. In this case, the
   * common clock signal passed as argument to the interface, is used as clock.
   * This mode is useful when all ATB VIP components need to work on a single
   * clock. This is the default mode of operation. If set to 0, signal atclk is
   * used as clock. This mode is useful when individual ATB VIP components work
   * on a different clock.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_master_common_clock_mode (bit mode, int idx);
  // ---------------------------------------------------------------------------
  /**
   * Function set_slave_common_clock_mode allows user to specify whether a slave port
   * interface should use a common clock, or a port specific clock.
   *
   * @param mode If set to 1, common clock mode is selected. In this case, the
   * common clock signal passed as argument to the interface, is used as clock.
   * This mode is useful when all ATB VIP components need to work on a single
   * clock. This is the default mode of operation. If set to 0, signal atclk is
   * used as clock. This mode is useful when individual ATB VIP components work
   * on a different clock.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_slave_common_clock_mode (bit mode, int idx);
  `endif
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern allocate_pattern();


`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the ATB SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the ATB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the ATB SVT
   * suite. This is checked against OVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the ATB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif
  /** @endcond */


`ifdef SVT_VMM_TECHNOLOGY
  `vmm_class_factory(svt_atb_system_configuration)
`endif   
endclass

// -----------------------------------------------------------------------------

/** 
System Configuration Class Utility methods definition.
*/
`protected
ZMK#A>^KV/RLcA#A^G7NWE(NRHf-2,R,SADCPbd9.5;IT.=D6F<M0)^,QH=;:.Z:
)RD9ZB;T.^.+M_HI2^7CP[gU?g)/I9gW5G7,BIGR#+JPJ\cc,Z?FMQ\O,b2;Sg#)
fHP>]5^SdY=&(&F#(?NgC\^F#12H,c4SJc9)IU1&U#4,8eN5F)d++,.6f?-5HJ1B
,LV2G)#;8WP1#\b7ddUXP28:T49a8aXM-)OAZ;BR4WOg.-ASQ1PDdGV;3,?,M7L&
GPZYA,WJ/gZa/8-XdQB2-)5f)2/(bcFWNJ[=QYI(D?TR<^RW4H:gD5J\B]88B0e:
I/JJdMf4YEG4BbJ_Z;@A&CKc^?8CLY85N:]4S(#2-ZJXe_SKF5SOAC/]bX(\,DLb
(B<.@333V0@^X(^W9;3\?01S6K.A)cE-?AC5ZBRD6+DF8SWL4RN1XPI>SZI&#,2P
FcCHIWD;CHWKP_,KL@9g0=#MbdA+gb326O8&GD>NQ\@.+VKCH)Y7EF]6YD2_?0I(
dNg>&8#.]g&QKIa3F^d>9:OQ]XAH+D2;F8_IEfH07+5895.)Jea,5@=<_[RR8dIZ
ESW,:\AUGbY[WcLeI2_UW=UZX9IZC;><W8Q&6LFYW6RMQ+dgd,=+Tf:3<ecd;4<8
4X9_cU8A=FVIgKCQ41YYJ?0ceF]W/+S;8/d<,U??7]4:V>ZLY]Pc)GLbE>d8JaLV
<:@3XHS]L0eH=L3S47C_5@LQE^QZJ##X),WA([P40,@X?CADe#_;EGA4X/dcAJGL
J5&MSaZ41B.:O>>,P;X7Q,TU+;.E4D=VA1T6Q0LS@)N]]?.g/V,@fgT;@9TW3/;W
-^<8\b1,L.;Nc0TKVY/BG>TAaPZZL#e_U7@>^V(E;IYcFKZ1[CE>NFRD_2Q&bWWc
:5ZN?J<CS7[S6JU0M)bLb,fUFO)2XR;ce_S9MW@.^=LB\Ng=GMF0#X5<ZR,LRG.&
IDEJT.7XN/\HV:J[ZW2b-DcQH4a5)AeI(HYYB?g[]HAWB_0WHTV2DFL5\dcGDZ_Q
WS#-6C..ZHIQ5BU_,PBd@bb<]8::DL=5<9#8J9?GNFe(R?6SH@A:D-45[bfbB0(IW$
`endprotected


//vcs_vip_protect

`protected
L_@\E3XHDG>>+8Q:QH\,<H@]\6c;/B&1-FIG@XN9P)NHeAB_8bFV7(/6,ZO+=^/C
3C8AC(>cI+YHZQKGMW6^1ITNEfd6EcJQ4OV,YVU07??[S?@[9TH/D2A.A<N\CVBg
Y@?2OfLSUaA(f^GT-aLIP9e_X<K]&PRPK37BH@ABPH&gPQ./0f2AMT\a+#/+U;(H
bH_JIgHS5SQD+eWN9B15O8^G5PAa5975dVED2=U88MKI16H_;1_KeMGaZ6AOUH^#
SAafd;2?5/>SgZL)e-HSY7UPACH5T:@e.WZ)I:W>K-[W:Y3<aX4Hb_TGDGf+,@?;
WdSK#96IMK)bC(=.d13M#9((E>RALZOWLa@K-7H<X<=-1g94^;HM5WW5\(TfIcFT
c7;&N8fcHCNCN(TgK@;F6]>T-dBZ_7F-I4>\L[1);90fIL5dX:-cF#\D?1C4TbLI
Rf;7O_[MDD?K<]J\\Uc-eJ\_(#DX#@bUG@/B=4fa6JaSU_[eKCJ0TK#CI8C3L2,4
[LN0KQ[C[+d2Gc.,C^U/FU>,O]fUHb/HF]eQ&9d,bD6(V\W(g8ANO(<-aW+P:J5(
<X9g]fP4[QHU5TJJ7[)^e_#8\dIXCV]<gaQ^e\3@+P,=?5\gfOa979G9,:UHLZd_
59Q1E0()JdaM+8JVF4WL#L@I3^fMQUMAXF.E^PC@G#(;4=XYZLV<(+U)JN3,J=Ab
:)T+<eb0[(Ec&D2BGKW>R3_^SBU_#.:\cOBZ13+g8+\9=N=QNJ:4:#g&B[2/Oa1K
D2I=A=bE>W\O[L^-#3C7WfIY:\D+gKV&QJIJUR9:[>_<)T\JUVC4G(D[4:J?G0>F
UO9[2>)/X]<J+RG_bB#DV-3TM4NKE\4-bf79YEUgX76&Z9bcb6Q]OAQBLA-E_aL@
1ebX@T@;3K+]^HO5AJgWYB;J0=PE7^&d7W>>=RZ^+DSWe=\XJ^?=_C.:]5K82B#^
)dEAJ:[N\6+eV&I=[,R4b[JXYgW=PcF[UU:/L?XL-PBK/5DA[#8RD#D6GM#>W8@X
gb)3LJN@>&,L/G#5:E[V4U:7V-F8_gf8/G33WN96ZeNOTB=&f>9GMQAdO9UB-)-+
aCANTGC:Df&LO&QUD_WB9X0-/,Z7UV\4c6\2(ONFc)DZNYTNd5]<\aO=>?.62;(]
TP0N;4P(Ve7TBOee\FBY<W0>9cfW>H3CDd[gFbR#1646K?VN.I2gEW&QIALfIM>;
ORDdfCI+fP>0fA_CXf;6-KA&KR&U?X:_gb/[9(Vd,bEUY+33?7<K)QD,=:<(\@][
DVWGWI_X+D:-R(N@A44?Rc(fB_7dc9Z_X#XcX4(N[(@]Q,-M9XPQ7d[FPL:>C;3B
3Ka;dNeT##FNI2&A+T;dU@TB<_c]GA);67bCR0#B;?2?BCJQeH7[3K3U0<Pb4d6?
XT4:ECEOW)c_^G]UB#<,3)]+gTfO+1+1]W7T,#a9#)_I9?HLM<6f26J+WEeJN\71
.f5;BaY/.=GbQ3NX)6D#)a>g)g?(>\OY]^L8BOVTW:Zb0)3SM6_dg2Wa9J\Z4YQC
SS&7QJXEE;C6>//8c:Y[0-</P;6,GVcU>eDTV6e)@J.\c:U,V275HZJC^[&aB)-K
^DU13aO#&>d#LITMa^5?X+a6IF/f4N5Z9W&e98VJ?+a1L+8.@RK/NC].USBNY<XQ
NY+T/6\TG^KTb)Ye>0/DI/Nc8ZZ^;8LaB[0>JH1Re3#J)NY5.FA[9PK5)M[A@C&8
G-8,PS\12G_M9&)P957D4Q-=R28#5+[)#=)<PVM1M<[G9&d=ZOAW:C+=O0NX.LWQ
-2OX-VDKM_-90H&#>^@[+#XP>NA)K#BLO+b/U+ZCV7#4Y,Y/bL6aO\O/UYWA?IZ5
(<A66dfagM(1^)MUEC@2T]-5K>JP&LcJ94;TPeP;J1)-9dNMPK?4_-\)9QM3M\J@
0RB:Y^,N9F#N^9HN?MW&7P+C<C6MU-af(&<QH;]/gc8Vf;Rb,BB4PQ(.GT6Y<(VB
>PU=5Dce9dWU_HLU)L0b5^_N_3[d_--KEXfff7QG&c+Oc=MT5LZ8:\JL[F-.de\1
-FK>=.b?M1HEXS/SSA5BM1@a#FMPYd\A\&Ub>C4cB/c@B:0X_]^:BF#[>\4B,(;)
U&\,^c^UWe8,f@Tb-G,#MH1J?+YD:aTagVO2UeT1\=4:85.U+6/E&S/:NGUL\7LP
Q-?c[H?@)@D6RbGc0GU>J\2bA>5K_0Mg9TRN&KWX,)G^&:L>RP?>-=@[\NZW&RP7
O]bGH>7OS]&]/aIQ[:e9))0NTb^1[SB;.(2FJJ:/LB[6TCB;TF758e52<K[/EVgX
f?L#f11]d&QK3S67F0d]]fUC27K^eZ2(KK:GZ_Re9e4^[)&BT.M^dJG)K1@\;#Md
U]2@;U2]eM30&O6,ee98Yf8Z<HeW/Icf84Dfd8E(5MdFe)aKbX8)B/fSDSMFVLTW
P9f:f8WF41=0G5A+eAZ7GcLeM<@J2?b;^dZd67YR:&V,6X6gGO;M=&WTSP;8UU+W
;;c#G?E-0_+N^A)/_D7ORb)4&:E^9</OD77G#5[Id&0f6@:Q;EDe\]T5L2]7;XNM
,M@30(7J_/g@/RF?BOaBgL)Y][M5V,fE<=0-Td#TD5J61U8fXe-7_gYX2eEH?Z])
L3.=_]c32O[I,XV\eK,@Qcg:Pee#6E7B@]<gQK9TbLE3/\/f,79,W0Da4eDOb\8T
B5W4,5)[<26;>^^_WE6a[2G^a5H/PIYe9FS)2J]+JDT1a>8X2D2&92M[X2M5;gb^
@@9K_K)6SEI#Ga=8[CBCG@M/4X4)MBA?6:CMbR^=<@O.N<^g_EdO/Y5P6UOb(fc,
9.-75N0QOQdB+I<9:bZJ?5P4)ZL8D3,7QNUa741c;OU]f-224S>)H#5b09.SL;91
^7-L&.#H-1Z,M49:;MNBR>[3#2\AMdbAE.D\=BEIO;=1QGW9^EA+B.++3(A66MF0
5T&6^e;C3bO583[Z4Yf/gH3<K93\6aBYb8N2K[H.f;@6=UM?T(Jb/P>6SY;FQX,-
Vc0aGJ+(H29CR>c2]-fFSV:KcH^SYAg.F_&B(P4L(.cEX>1DG938>HZ-Egc9d(aF
RC.AXDLV29Y&W6ZI>57Hd>5gTWb,[<gIF>_\Ga-E,&U+EVZ5P7.bSE?W#V;dddf:
S_A;X,=?TE:Hc]Rf]/89d_FE-B,J>gWK+P5F8EJBBJ9:APB_@\dU/e5JAHg#c#GP
U2a9/KO1T:\U]62S=39HT(-CKEbf;6gXR[]9cCBeGQC?NASTY0#NYIg7[4#Z,/]D
=fF>I>d<M2++<-bg^HR&AdVGE+3S#FZJNIb#EcSA4/)OXd\I>SNa@@&?B(6]BKS3
gCQ9\Se&DeK5-N=+[\;PZTU6&5aKd99NR>83_fe[YO,5P^0aG2<5^](KG5UP2\=L
39?Uc;^:QVa/X?-Aa6K2\0^2OBR/>MCMO2DNFXH2ZC9(X(cEIVC/<EZVA5Z]M]aG
+<3VNZc(b7L:]^^G4D+9>60>cccSd@[91Ab0;_a4[K?c=C568fIP-#IM)GKfX&IK
H,WWI57^eAX]ecFCQNPP=C;7>YE#]dEa476HI2Ra=RF=CdWBgd<4@@]LQ?2):&.W
@WD/O98I#ZT3N3TFOdZC2NK>SJP1fS.Y#L^]J6\aK=GCG(\8N@IL@<R?6X98d+1H
W-W?Ye+gg3gb1KEa&gcK)a7FY\Kc>]&=ELWC??O73HfD-(PO=H;C+4<Q.3#fQ;3;
,EaU^D.dX)WeQNH^<ePbK.ML3GL]@X]L]-PH24/+[O?8+MDG^TECF5\\b^UME3K?
:-?YCXXIXeC@0GD#IBO1))O848aC>B2)b4EL8\8@J#K5QM]V.CN5LeZ61S@eAH(G
ZK=bF?XLH6XUE7&;BPL#]&90.3UPdc:T8d2a#\&#.5SM<KP<<W:1&VW?I_=c^K-B
Q_N->-[KF9a0X^^57NC.J&e@M>]_&H;2FHPX1/AW+5.;eM_Y\.,R49G/+BE&\3LE
[Yf)N)SIX.)8L68GF8><5R(\E1\f<2c]4)MbM,U5.G&)_76\PV3M#SPDAZd[[<e:
\N4dTV9.,Ad^7+V]QR:48YEFGDbVA>eU+C9b,=QV4]dOFP^;QJ9];+e?c8QOZNJ;
X&BN-_>BaG8[b>K#>@AJ;a2b^AKMD<WC=2CUFO.MQXeEb<2gXMb,];6K(L:\CbYa
/N0dWT+U\LWZ1(<dcFQ3RTT[8B0:Y.W+BFe_=MLaZILF/L3F>8K)U1(44_SFfL&4
BdSR)E#ZWW6H:Y0b4C29dI??+c@eMJ=>44>#=KA,J2BB&J/DZ[?/)N\)c^>LJG6(
9>eD^X):?IZ6+V#CH35R^+R_EYKL.0>g<>@XN7>1#f@[]:,X6.9EET.HZSSc-#BA
ME>)d@+1+24ITT[d,&e8;GBCaD\0H+^613SL[IaNOGQ.F(fQ,bf<F2-66dd?U+Pd
3BMJUBF4<6I6BI@U2C7NL[Q.TH<W&9Z?F7(>3TQ7B/d5>g]6D7]+XY:b>D+P@2Je
UWQI>S>c7A9dL]NgUfNF/WO;R>;J-g:e.P^+YW^)Sg.H+/_.UGe;3X^NG(GL^O(I
YESUP)2H?F_C9Q8K49..1C;6HI98TG1#g<=JGFEG<B4P6a(61:Qe?IVN=3U(LN#V
[eHUV3+:^6XL5<Y[@^O2cXV[DX&,S<c1+1:XK-^R--Y-IB]:2;J2,K9c?eb>aT?9
,R^,2H6bXDY<=TQQ\DZN7(YWIeE)2#0.:FX?3(Q75_2CC?TOB_H:HW?#B@<eS4RX
W#[c>G[(^SUY3/-/-TMBAA3FLM/db_]WDHf+B)>AOU8X,1./==0@+b8+1)0]5QDZ
8<0DXERB_G5]NNBP6J&g5JbN0MJ(@b^+./FA&\F8fB[AG2BDNC7I4[#c=0WB\Obf
TD668K9d(MJUZAd[g[CH((QVN52[/F)cE8JRC[AQHL>JM?=[@DbL4^-I^?(DF8?A
O=D8<L<GKC=Dd9I+GM^:L4U<_),T8Wb@gFBF8e\QQ25>,]\_]04E4QR6>),fF3V>
b1MT,Y+<8A#9O/33#d=,/e.WI+DP<Q:AP@,b3FR?f_FcAIfB+HD96^#BFG.63]HO
0;X\Og]Z-cO2#1G9])8QH;J_>.T0OdK]fKG(B#ad^51.:_;:SI\<1R-c]W_aQ/SS
=R,ROM3AW(a36[ZS02:89K\^@23a_0AHA_M3JcYH6-F.K(&H2_((]g(2VEV0KFg@
=g90,NeY\EeA57gA_TgPJ^9:N]DZe_NI)J5VIbgA[A3Q/T2/MI6ZaD0#R;2gRA27
(KdZ9LOc6J.(\ed]L[]&ZJ5OX]@QN7f=fO1LCdGH1M3+LD=2eJYc#G]gAf?e9J>_
^,],YS/A-&1[+-\YRUa>=;TEA#&90f4O4EBX03I=0(V(8)\&=WR&\I0[I?>>P+P:
(Q61F(7Bb\^NI)@BYfU,C;)]2Y4eO.B&HM3M[c4YdVXPPf/6RAM?^g)@9WW,-T#S
+LR;O7e;;@1K_FD11IeTaX6SR]Cb1M:WbG,P&WK+ND4F,gJ)?G&B^_;C,YdZX]6f
2JOK)PK?3,+))&-\UL#gYQ)L>26KE:)<5LC0&:UV/(+gZHK5W,PQ<gSd]?E+0?RK
A)G/<QFJUOc_d>3JY^6gc&4P<S#@WURdd^c/YJ7H>]e=>NHOSNI);L#e:DEQ<#WE
9T:gG0DJ(BV_2^NZ;)?d#D?WZb1+6].-d^/Fg0bBFMB-+W+g_@2cRe4RY5>R/5Ud
;(5YW[cfZZU?GNbAU>,PA;Q:JWVI)J))[OH]gK1HOJVW,:P(=C#M55f;DYeO-d/S
7Q61U.#\2X,<E:X@M/-fLUH@34UJa/0g:S+I81Ca_,WEV1?HRWM/I<-8:fYW93PR
488R@UMJY)L#I430f.\d_^5Bf2+L<fI8R97B+GJ:eH1AQ]A2S1M41,R_,(W>X7ZQ
PeRVO1D&R:d>A]8/YO@OEPFS.BTI/b;(_T.eOfOK(/T^cBL,>6Ae,,\#bVd@PeIM
,0.g\1L(8^1>JgQIJJGT[[]HJFfgXFUVccUQa374_0>c(HQ0YL+MTK&NL?9dA3-S
=e^-0L?UC3Y<SO[b+WTW]Qdf<#3-5=AIKc-&)L.DJ;7Ia)JE,^1/FZ,PQ1=1dM6C
B@:e#Yb]IMF0.@-<fG+F0b2Q.=0aPMJ+AR6M1.64)Z2=GR#0P^V@QVY)S@4-H<@A
c//d,M_CbQ_]fMbM4>]8>6aa7A.F(75;3#Cb@V&?\5AIHf/>@;(I)+P,MCMZ,)/=
XY7)ggaMRP@HB=1VTWD80#1ZC0F61484KSadP2[[.5NLV@;2I8=\?ZSA3#D-Mg^W
^CWNN5PLK^)?g^5HSa.e_02I.95DHW1<>?e<^+@IE961M?T?#-5Z7gW\P5:9d_bX
:U.2(KN9IA)[)JRML?M6^#SY/[/Jd(<;c_]519:?A^1ZPHF:/K>@T@+1f3PQ.XB2
(Y2-:De(V2&1)TGIfRG)@YZO/LFEK]2de6F;b:a=?)+JQOJL75#C,N#VE4fQ7>ND
bE\VeJ9Zc9K1(1?-](O]O\8W(>TA_QQ1W.ac2W=YV.SK-M]3]2V_AB9Jc>#L((QQ
_HL4-O[9bV^HB-39Q0@fA#UOP]0I-#)4&K=3DT5PJ(5D<Y,32\_@a35LE]2HF.KX
S=B4/Od6/;UHQUI+,ZR4+G4Y>g4>>[;1QB4HF_;]\>1<AXM&&^cW?3(HUM&.K]53
\^JFLO5\T0f5BMMC]a)I2_2\2/P:L18,,\b55FN6;aYS^K)DXbK2g9:_g#O>[;c@
CYZ>/<_SXU5R<)#&a3EB,OGO6^245e/N)9424Nd.W5-/.]UJUf0K/GD)-\c^T>N9
P]4D@dM/_-;Rb@Z0g#,4(37LJ_e+LX_PDY/Cbe7Q-VK:g_+4VX0AIFfO137Bf\UG
>5GMIb?/f)T1UHYFVFP-X(H^&<FT\e2]^DZQcLS.90E:Ub4U;[]W1K=g5-GK(I2-
7H:&LSS1]b4A3(8Xd-cR1M4PQ#fDK;V\-dagC]YW2M<DG4Z<W]C7AA]c<9#^JGQC
Pa:=bDMfc)::f0A_A=,0CcMD6Y;Ef1YLY.3a+4TC:I0OU_O<2MFQ?7LQ2;&;^CaO
.<-+HVX>b7]C;5G@DU]83J?<W7347+39R;TK<GdF,H2#<(\KN]:]LdI-,//)=ZA6
#=@XFQ,b-+B]+[RFPV+U34LGc^)+^TfV?1L1&#ZF??BXOCK-]U)Rb^?2\T8YV#K.
5]W@+I3\/E\_E30A_J+L9I[.bO1@YOC8VUE#Vc\5081=PV)1@?AgKfOcA?R+G;/&
G??8gPZKg-5RAQT2F4,ZM\^>ec6RbN:(a1V81KK@\^LP)6/X69_JQB+/[D6f6b//
Q>b-M^IWF<b<:]acX2.(N5fH8K7AP)RVE=SIaXZBP9<6W9X0K/b_/QYL#)C3TX5Y
FV?bJ28<,B=RF]7T2N6d&IY]P)XIR?cFIfg?L#;W.6&CG:U:b@GN+F6MJ^)_8@Hg
DO_((^F6SIcN86I+e;f+[e,((-CUa_=SZCE7-e96E?+9@[KFG<OX=f4fNHX-K[0g
DK3/>MS,b4Ya@TT@-WG0g9N3/_BU#6Hb3;Y8S@C#(+/)RQ;ZV^>LafLc^6,-(Q-H
Q?O6.)&WKM3?JNCO^<1GRMgMgV2=,ZD<.P/FR&XN,a5=-Y7^#[E>)/SD8W?)&D7/
K&VaVC33V[?=aZY#VVT.d>UE\GSS-#)1PHa8B1+M3.@(O8LL8H92e2;6V_dO8+a5
bVS6FDaY+;6#dFA?cTNX0[[LS<K>-WAI=8-Vd4>_TS[.CgX(.XEBL@B>P.P>&B>7
YSddN[Gd>GY(RF\@UVVPHK^/MD.cDJ-/GE2S)T4e0X4R]CR=c[&RIAD]&d/T>6>-
c]9^.d;(EZdP^\V0<H(9,WW1)51HKa=aFcg);-+Nc]KOIW4S=(LX\32dPA.\02W^
,[00T@eKD=],XEW<.\6cT[cN]T4GE-^NBT[<@98<A?9W1#9<2f:aYFXJ>W-I^7:_
2W?C?,)4I6)L9gWI8B-/77LDgc(FJaeLK.GY7O1:F7N?ObP,N[64]\eYbFQQ8aHF
.W[Ma<C9X@1KL9\gd>==<Z-U>fe8^I,09=@@7@&RX-@IW@V;USaZNNJK2+O[=B+.
-G.+(QAd:K[5e=YE2L]937>F0e5NPV70=aU:JI9WH:=O?+9]1e_#cFB/,KZQDc4T
>.:I(PC>=<N(&KKCQ&b2FD\[&52Y]DJJ5EfP?I<cdNXCP-><g\gMb(X7-I+,dTEQ
\FcL\g16:.EQD-#5,&3&6)]8GGX[TH9Q?K#075^?<5c8M)TUaFPd5P:7(/88YUI#
D7DYRUU)K>b2BJ<;O9[3C=GF^5JEd8]ZZcdLb044Y_Y#@6^c4a](0U3H9,^08:0X
OZFDJSF^0_\_;\COd@bM0,A)cI.b,+79&VacbBN3F_ZaX>cC[KbW0[L0<IR7edRB
_c+^O0:&Sfe9d?eFc[T1MI#W\S5S:@>(E/[Z+:]/e+.2TL^f8]cX;aOBF,R,]7:O
(?RPOSF#PFcBfeJZ+7(7A(\Ug-]IUd);g,-a(>2S0WU6+5#=:Q[(cLY=S+=eZ4[U
I:&98RcdJ]W54\Dg,)gN_=^^G)OPBG^ZD?[N8<]T\:gUc,(3G]/)6CbIZMIQ(FKS
E]7EVV);\K_=S:4f:R,1EMTQUU6QY[;fJ38)[QTT#^=CVQgY+(PKHFOa)@@-#/f(
4b,B9#cXb&Ye5]O83L(C)XA.J(bdH(U]N#3,/<S-]G:c1ae7^a)>eBWEH(F4Ee/\
3g<JV9G]8KcaPAJ=0eQ9CB5\b>2>RPIO+DVOad1>.OOG39Q(&.E.18/@6c@8>bLg
IAS::D)E^N7:)L78JD\UA]#/09\C:Q[S@-D\Y33gL.8M+YBBd7W:[N+c>1)S:]?d
_RFTH.:gMFaRD(;ER=Q7[VNSPG0)d;J2eUg2<CYYHZcd-T_bM+_:=&_ZeI[U4K70
I^CW4WaYNWC8XZB,eAN/g]LC4bQH&VNR/GDHR2I.FB6A4<:@X7M5TfCSUbPYeUAX
74<06C_9//bDPT7/A\&VKQ-d&c<^?b.H4W0YcO80+N^UXH3YSCOVT;VOQ_3<S;1]
=bIdII.L7Q8-E&N](@A3d08O5g,d06HEE?d/-dIL5JE:7,BVFfL];G93eQ#g8W_f
Sb-X\LdM0-+GT..;47Fg2+g(JLB7<74VB#F,29),BNQJ+Kd3gb?CJQ)&AgP?)4N3
HJ:NBFe;CZ\fg,WJFRI1cb(=de2b92a98E^d>Lg+&.:S:^^M4RYML<J2@MMM?O-S
ZBZgbY:eBXa.2[[B9S<=2MO][R]eD5&J^O#81D-WBbV;2:1G0A:Z=FVLUadWJKa&
MA3(TS[.0E>(OcI>WX3JN[2NgT>@SLA.KAXE1H4H+fd+0#R_9)S_DWW<+_7^/Q3#
[2Q3(3K1LK)gYD:IE]@/MbKdRN,g[H/88;&,]He((e@SSMX@:PS0S1[@C/&5FO><
Q=0U\0N2].1M@P/eV5;QXQ0g=HYR62IJAR9G=a&#Y3GH_TJEg7RJfEd?@/(FFce7
TM3B0H/ZI^]eCTSR[5T)fbV<<H#8/fc8K7cJ;\IU:;31DKM)HdFDJ4+?g#?-Z,+S
]g_/D6cJe3b=,6C1b@A(dFFXWDWdKU7YGGMFG7f8S[UIDF.P-\U/.HEHdR9YJKX]
MS.P3RZeZ;B.59XP1XaU;&5;caME1eGT]R<EcSP27>c,c7C,?W[aH46X;OH;+f6S
,39aYdKA0acCPR#&dD5g.1Q^3dbMJN+Y,4Zf4NBMg6G5C3/.eF_XPX0W&5:0OKX4
>QW,1OTf[X3BC8G9WfC]<5NBY4(eD-ZNfEU#[(UXQO;4Ygf5-Y_)WA<Z7J<)(^2U
P]9J8[K1/<&-Wg\1BH13BR\ID(/CY&P@V14WRB^BafGEMFNW)SZgBAJLB.E>XI]3
74T>T;gRDf58CT&:BGYN1>f;Q^XOeJX>0OCAC>\R_=[=V[]0TNYPQ]O>2P5IFXNV
L;JdPB,]R(dXMReg3IQ)V]bI#1b)C(:YZ]8;JVMSX3Q/XKS3U4Eg9CYTYC=\Ke9[
07=.dK?0/g,>8U]AY\?dA#c9F82T9eNfAA/aTU[:OcP/Ed?05I)]@O+.CJA_R93V
bc(0/@^ObL921I#Z./-=H88YWR>gX[\O\3MU^8YC[/7NG-6F/.e5<-_J5LIE2:5H
2GBL8,+QYf=cgZ,A3D9b.8);IW=_&PgYW.D^dG_SILRVLJ=.94R8L?YRTaDO^#HU
TB8O>7Udc1D=53,#G,cBJQ_?2\2+0OZMC4/?)ZNEa4@A+Jg3GA,cMbQCB0AM(ZH#
/=SOVB8GC<V]^T_gd6C1\^IJ\[^?COOZG(0+\H;W716Z7Z[8+-UZ+DT6\@_\&b0\
#>:e><TV4@^dR[<2KU6LW2b-02HU8.1=/E4&H,HbQ/DF?.:M@DG\A[X@H(]M>DO3
4Dd9,>F(&B5E,&+9<B3@XIYGW]5Q+\&EU[YD+6\NJOR4#F8<MYe?.[HP7#C/C9cH
7N8@DF-[J[]8_=b/KUCFAa51-;/_L.1Y#V#Z,&KOIQYaG&5[#.>7\1HdC2(21ATc
Pf=c&T.&STM7?^(;1E0a]?g)44W@2E7+:MfYP#NJ/8#.=HRM#UZXN0efA^-;\;H5
,2R1W&-P^Z9XF0dNL/eFdVLH-GgKDeg0_2[3DG\aS47YCHAdMfY=HU[NS=G3<]X1
(3V&V(G,&^gUd[>9U7OJ&N;@682[YKO=6KCRR04aOI[\DF@gZJ/Z^Q9\d];V,G8a
JY92^c^5^bR0)O?>\MPO=IA-V=/N9-+?L;UX#V4g9RPL_C15F;PARdSE7JbDX.)(
ZT^DI<1A\L##f,Q+B)-f8EG.VJE:9UbEgH0LgKLBa-;Ec3/.9&:b8WbXeJR+eWN(
@J:#Wd[c?R</Q_#U/,dN^e&=AIZMeBQR),0Q#UM:ZD3D5H1>Lde.&/CY14A+f>,&
J>be;0fMCKI)L5?<>^86DPd]I[e1bg;;P)BF;6=VJJC/MBV\JKE__P,N#3IV/M[_
?,::<FCFZ-Z@HEc8Pc\LfBW/Y[ZB+.FeVf.af]O&D]@JIX)FRF<I:g]b:[.JYLbH
Vd&1O<?Kg\;daMTB9e_&JPK:_K;0gG,X36GT[D]SX+=MWT-H58=9/8)dS3U:9RNB
&JPc+B-[BCFCScRf=d.6N_F,P.N>KZYU.J76KRdSVS>=8[M&MVM52YWF>RYP0D))
UOH7/86dPg1T=;4<^AIRZeJbR(1,_1Y-I^.7F?g1XA>(DJ4B(.>_Y0NI1YC.9542
.2c\#J_5<+DAB\LD7GLVJ4Wf\6N7Ob[D>]]YOKHZ36\SX3LEWV-cZ[8?C5RcV-,C
>bFDHgR&K.b[bW_Z>S.eM=8]@,UMP:2_H+[##>YPgOf:I6]bAA=e/UK11@[V[:T1
H8ANCE[^(cNWe2ZN?8&DG4XB.Xbc5)D4?#=;D_B\(MK[V88TO.W=WfSZ1BR]F]79
FUg-\:4+R:;78EO-1/#=&]NeEQ\\cL[/P^dI@eL;K?K46NPZDR=Q0VgYS>>DM3dM
7KH4)ZC)J2C4SA(C())caK(:0a,c3YW]<1OK<f<+)(+:,H_);fEUQ:BBVa(RdG^[
H9L>G_3YQ6I;gYS8Y6I5+_@KfaU_IMX00P[<B8g_X2,U&F>fL/8NRM:gW9&PcA-/
fg],NgP\7aWM;9[.N8OVAE+Y9G9BRWF;^YMI/4I6fN7.76Md:H>Agg(d,g9L0W+H
\(4fK&E9?MgR]EPWDA>GMf.=+_IFa5]2C(=?.9(ZPA;(3J)HQ0cM8_\7?=H?RTcA
Of;N_&D)4@C:J_B@Q9^:bH=U0);.YB?gN\&4\\#UYDad88K6AG,;@+J54K+bO,J3
</4OfGKa)+0&2(YG=g#A<d/B3>/e/LeD)W4K:LWV45aCE4ZL_1E-&PMa^I>:8G#\
D#/FfDEB/CHF[5U@.=bZK+7/=<L0U4FCZ[WZN:MEU_TYS3bG@.b>DRS#-G_H\Zbd
&LbD>_A-T2PLEfMe;\OY5-b.=I)9GK?e2]Jb;,95,.T0P[X\#6&6#H9BI@b6(;N(
NZ.AROF0J3;3S58#O&#R<&ATO2U&a7]\I(N=CIF_M\G.XD/[\a\O,bdDVM\dAI3@
AYEIZb\C1Qda,C2Xd[SNTHa8Sd86Z1,/ga&gbG,P4g,cIKB]O;XVUQfa;;&#1g-&
(_3G6;Z?XWeT97X;^5:-QUWPA0QPOV;Y9>Ff(71#O\2bS#DL-<PI:/-<)#Md2WI>
WU\7[L4E?5N;d3#CXK43\WX;HYASfGT,Xc@8#WNRcHJ]&CU42(9PVZdEAO=S]dO#
KU7CMNA/Z9N]>b,ET8-G@Fe2T?GZS7K;.D+SfE3BX_2\5+O=C>bI=OH<FJ0&0AaJ
DIQ3VZ-e@c7+,MG)OO<B3C5;RQ20[bBaaDJH9./5QVE4#HT?^1PPM&QF()@WA<33
-N#cU@[J[FcAGD@FP:gKM_UA83#\=SJRXc/fOGTX&?U>?fAc<?PX4/8dSKg32fD3
@_c@URgK#YV+&5EDLgb=XW5(F&C2RN50]-BFWT(:2F980Cb[ZTC<ELb:#?.FOWbU
1DZ9Nae/)74SbNZ1N1]DD8IPHdPbSO>(:ZK#[DK:/O]/K_3bJ6WC+V<(FSWE<WN^
IH0.(13757YO/88=Z_<VBE3V,1=4J4>X=XL_/+>V.4W;74ZRUEDCVf.V.B&R-T\)
/H608:R2/G7dO]MYUH-UNX,Idd6=KAA7^M,<@7I\DPVe46BS2:2O977F=:0?3R7>
4ae5;1/Wbac)#IcJ,(2CI,3UgA5c5W3\(_(9_+LHX=0(&[3NfbZUTGG:,W;?^5HU
\,\K;CbGTXd5JW7Y5bUTTcLSAC1[@7gT3/-&^Kg)Re:[AY>@NY/aHEVF3]7Ac(A;
H]Cf/gZ;agBM(0EOedNCJNbOQSPW6cN;2cFdE76SY^EN:XF3eSgM.6^5;caUMIBO
<\VL-FZ^\<)gIAQ2#L)G91Y^]CZW[.g7M@^;?>c[=Y?\DO:d[FP]5LS.Ia,(J<CG
fGJJWaJ3;DT5Vd3(LLDSaOf;T5QZ><)PcB-P@F2)-e/f>Z92bJN0V[X1f5R(/N&A
c47(BWKM6aQaU&OR2K]4d=>DPe5<5_5Ib&P4DLVC13_XD>4Id:[W;U6U-V:,Y,XM
JGE2IG.c(BG1)/6OM_]QL,VD@+,-U:<B6a\F;\44g#0X<@8(TW4R#+H::WXFXb0Z
eIa?Z[L5\1=@#3[B,B/+c(M6C@b7dP1e<aM>\I>SVaP)<g5,2c^M.HS9U,\(-G>A
A:d[,6K/2XZ9&Y=DE7//^B14PM0NFG>=C?EPM87>NIbFG.L^YZZ9K3&+=c[f35U]
8TF?2Da[KV7A<SZeg\Y;YP<2J,Z8F09=J#1&31.g3,T)72A4U5]gb)SA4[^.dR&E
:X-fO5HNM)HD^?(0EaegTZ7]cfe#_45LS_6FMYC;;H\F(-(QYbK3Ic2Z^DQ#C9>C
[UNGP@S92MUd#I6I9:;N3(#[)R>5(>=R/J;b+8X^L\:079Z+NKD.2-#1V>Na)EgU
\U^LA;]:I:Y4(_F.a1HX\]d>4XBSg6>Q32aQ6G>F<^2YT\W;dP56[2_cS?LMd_&b
W]gEfMaY61:SR7/:O[CQ(]<Rg-gHd+/I8g>&QP;/@XETb/^9\Y[U+M_^)Q(4)+Be
>+^cH>gJB>89aUS(P4>HZX3g,\PLH(BeVaJ7\\H#TS6T0;[.T=[]6?6:PYcXUQ(Z
?5OEd15Y8;K5W;GF(N6[,eV/<a=TUC@ZY<Z:PH]F[L[^?R?#.)fg;KPNV/f;FPNB
5OKZ@(2C(9f_ZXdXL-W9Zc[?Ra/J1PXVSfQ8FBUS,3)?V/C7]_4e;X__Q/HbKLKO
;@JB,&U,DR]/W_S/Gb;TT61X5dgT?[H9^B4<Ng;4-L\4a@IB,Sc,eS58&#_ObAGP
3@gH=-\ZOK93c_1PN^KV\ggN@g[TS&O\FZd&Y1K<VB5-3gT#NV1\;E.9Z+T4WM>I
D.4b\2#;?;:YHaeI/SEF?]Q)0=U[0fZbV+Ag#&XF1XX5YdUWG0V)I+1C=+NXb,6B
P2YfQ@?4U>4Db+R?,<,F9=7&;/ZV\1M\@cQI#\7AKN9B23UYQ1654FVJ4#XXJA8?
H@QHUf4NNC?CZ^PQ7_,B8^+V-C/I4=K(/F_VZ;RDcFU&a33e3JeUQONX+M9XTTAP
fgQ7(O(9E]HKY10RaD/\DU3-5:QIA@P?FF<a>\8Z3:C;&;:+M<+@aH<A;D/F.eQe
(M:VBe7<aGe8fS-H&@A&XKe3aFV7#e9;I&8B2fO6MHM-8F<[,ONSF))0B]Q;Mca:
b3_R7Rf^@-9UBNKf8fK@1)BO>L[D8cN80bGJG,d[W7V-1cfZC\O6ZR(F4eZKb<;>
FDZCR:6^QP[a_R/C-:NA-<f;SC[U-BR<B>VX)OJ/QE_aK;=BaRYU>fBC68:1N.1Q
DN,O_eG6>3J6>IG9U6WTbB)9._W;J+I2#a,b+@DC\GO-9Pb(&YU6Qcb/N;)0SE5c
SM9>6g9Q.=>W<MBH0S4Me(bW,Y7SYU[@ZX00=JC1BbW=Q@fc:F#1bf=8SY>RWA=C
Q@YUOI\5(K(>J=5]RDER>F:0)W)D4TY:,7EW0-5ES]F;MGQ[ffdVeOQN-bg(Vc8A
:3EFX3AUUZJ&c1f5T>N9S3dG&Q:aW@,CB8Bdb7?5E&FR5^E7IeY1d?:Q\4QL@EC^
:T9YY,0=9faW1,/AC2-=B]+L,3P>cI1;@Y[<:@H-bcf(E^_)dA1^EPCVNfO@9WgQ
P2FFG\.GL@M]-#XDKRd5M?TPIfQEIIaX[;T974>)fM)-_Gd3XP_8=V3JB@8DRJ7W
bB)42]A?=CG<7/VA4M_Hf9(gN#TFY@AKeCCae29F+]H.ATf0YcUb_2QM<OB=?g14
BTRa^2T:S>TMaBf(46]?3[]Q1_WWEfC>ZMHE+=84a[HR4efL&_S/Aa/?Y::BY?(0
bBgG26H0OCY7G,[D,H7H1WF/R@IL)L0GcD]3b_9310>Kgd0IP2])W5(;d^P=WeTf
A;1;T:/HU#;BfF/P<NK+(@#5;4TN5bBQ\T72+?ZePdO]ef:eC)I=<NVN2UJ-.Jb1
Df_:GPJ,VD(4CKI>:K0L_[\10f6c>JY9dB7J-Hfg4Ff[Cgd[.U[e^854SQX^FV8T
V,0(;E3WXXURZfc=79_NIEgV,..NYK0bE;(4(3&F<,^U@PJ[N8@&I&@B9e]M?6TD
fR?]Q,09N,d97OV;26=RR-5>#ZB_.PV0Z]UP]1(2V?YcI[LHD7CAF91IG7c_PJXC
AQOY:_=M74&#fQ^DT40JW/HC7,I6OZc2&:;Ke+AB.Jde2J[2UIB\DP]eW(WS)f8X
5X4:CdQ1B0_(H&@P#V&[QU<0I<BAaV7NFSLJaYS3P[=VOOIRCWNWC(.[bK+<8P^-
--Z&NIBXK]#VAJ=RPg2@SJO+B11&]K1JL.5IG49X_)[B0GEAH>^CG=80VI81?)-K
We90TD(A7[ff/CSDAgI^RJ=E39=49S2TgTVT[)D@JBcK:#ZFOb3BM59(XMGc>GNJ
N.8T;.:AIB>MVNN8:N3TTYY5[af&TAMHIS/KFD5F?-,X>G(;=\+EHEfe57Ud:W_?
g+1_MQ5?BO&587^UITb,IWV<=Lccg;Se,;(S^SE47PYB4-\9]c9<0,aM=&^O_4Q^
&,aV+7LZMDe,E-;9]-dFV\Y07#d\c\2\9L5Q,/3YJfH0X]1KEJEXVAKa<OVA?RTR
^6:?=3Rg[5baOXME5ONfNJIS&Y(J:TL@X@U0OPBL#,_TWKBFHL+Q.>GY/#>,I+,g
VJ3TT4b2KA(B8=cF6>:QN)CR1G#<,1fU-X:6ATbcc@P4dA^STU6>8[bc6H9gDKRV
)JA9Z[G85bG-,d^\8A=6D6,EK2Y;HBS,0G(B)8Yd2-6bL^.cG1:@>(&,V^\584-G
AB)G_0FA5)cBJ+-YCcY_Ob/M+\P1de.36N[gMUYC+2^IP<.;[.EBE63c]=S7#>,?
Qd,8[O[^GM?=>+>OIAMQ^PE&NSX#Wc&Z5;G)53=A;#I?O[MaN867cJ9g_]:=6YX&
.aLCV;Dc#-5gIYMG\I^I:B./Lc6I,./Z/;?18G4Ud&+eMC45F:MS30^0fH,3,4SU
\J)#d=\;NgICR2F1d5RGWG;QASE#4L/]:T?B(BDE^\FgDda_#]7F^PIJ5FDYY&T4
P2F9UEH_Q\<d/P0Fb75Z.>^_>b6K61<I=X\95F&/+^gVO9JG4f1PL5_TY<T35/C.
O@8G#9d=L7(_GOTE:/ITZAP=^+f(?:993K(Y_:9X#JcTO2(#K#YJR]bWbGI+Y??J
UU81;[Dg/_Fg,Q>M6HV@BE9LgWJ[>D((f&_&;aG+Z5#0(5fZcWP6^@3KU=/ZbO(P
4&-HW=.K@1O_bXV,HS\4<\E#M+-:<:/]^6#3OL2U_I8H&A/IOcK[C\SP5PQ3RL+U
2F\&Vd#(-0gH=G[A:_DTKabO8B)DdM#b#(\OBNbN>J[#((T/>VG<\Z(NQA/T^H(A
&UYgS,3Q<HQgeD@AgfOGU<Z]=Sa+ZFG0IN(QbeAG2V[)JA8SbWBQ,UH\C:J?B?(F
2@]c,b\MANV..bK684fJf>Sd_V9YW6=]X92RXPdY6DOeU1YY-1F0_;Q;;_d^GFVg
(bP(:>MPB-LLCND;g#H<#e:[#GY\GTBN>e]E7)QAg&AVM8R]aET[+MLgb(I40Y2\
KQL/>-QLD3;/E7e\dGdB&(ZV:dKb4AX_YAJIQ):=(Qf]0:CUbE_e-JHP]>D]N).K
[.>ATVO)\F?^@:Z\ab54J;JWP0^g>g(LG37]5IBW;KZOcE.9.Qd_^S<6O0g0I\G#
^68X:UO1,3NU1XM(<(]4C4#ePa,^?FXF7-)//ad^UZPKF,H3X^(\/76]:D@&[3ZK
0@H>.-#E?K,Y&)1Y@<)&XH5ef3+a7(<>.T32)^fE]V5U]G>Xd]_E^.6]#\#N-52Z
)_JaJJA=7U7_CHJ6S3ca(1:.1La&P6P_;-EAF(QSaZCE1N4.0gO6R9B+)&].:J;)
J8.SeBL5KY>IQLM1O6IKHG(EK[X9F7-K9?[0Qe5&Z0J#-YD8c7d.1/?QaQDU]:0@
8=1IY7,[QD_PC(E1:Xa<4Ef/M&7ce(E\a^<,&,\XeWXd07Q(/E7GX?QIKV:Qd?;]
\FJYfSW_Y1cG(\g9FSf&KbaKcbD4(D\NZbQ2DD1+A;0=.&?[99E_eZ9a_,<D[9MR
+F;d3-0UAN2G?93a2+L\U#61TF0&B,>S7Q>[U7^QCfN9feEg#3b@P<2O3L8Z2^>9
OQc1C.<A,a;O6O=5_421ST(_P,>fb?U559BBa&:g;:KXNGFXdTU3FX^2E[(#CJ2.
UA0J7/Y=/KabfKX-fYc1J)@R5;c7e<JaF7B\H7@0XK?LE3@6g&Z,+#Q=aM.&#;X8
1ABAfFV7<?OORYUf@1<:U4&R\e\4#<UNIHCaKO8&Og;OE6ODJbB>F>+2<^;C8Y)P
U(7OQ5Ze-f?;00^P-0bN,YIFZ\;+XA+YM>e&E9@?W-1>/009^SC^RcZfV5&X7g#N
N[Gg5\/dEeFPJ1&7;39g<J80.d4ZIJE\4HR+\0^.NF4-[d[JMfIf&&M@(KR4X].&
B;.WS2.<P@P9>&L>QfQa9F9/;?0cSg8Z-8B]6/DZ])bVC>f>NfF7.AE7,IJ(EHPQ
7,+-,Z:gI&9W#HVdN9O,UP;F0F5Q41NM@]BSH84R\DR_33?d2gN<GfWE=MN0J5_e
>9??&#:SX.5,EF7Q=9SQD?3g)M4=:e[0)Ba=GOO.PU5bcQ?ObGVa,_.QXf_X#;0f
(4P/]:<QILABB@X+LXbY/bA<-8a=/K^e8K?;A?5B@QMQbID7&;e83U+cc_;46>1L
8DHWIM9++4S@>8AW60]BH#]CfA4edI2:9W@:Q^UX75?V1GH\X3=2RF,QC8QDB7gP
?ODHgL5LHII(AAdCdIP^AMABRL,UFY]4/IKD^B?6>5--I(aSdTGLC5#Ke]/ONFN#
-HN9RC+)c]J2;@30W],dYA;W+Lg8<+0OV=]C@MK9gT.).QL^Y\BODAca?L>CB9&@
>>^&TSXSL._HTR?B<Ef5Y7:P<Z^LG&WM_ab.F[(0&E)(&@<N95FZ+Ee;aU22fXML
NMJYd-)5N4;eZ1)PXM]:9O(OceDCASP<JU[:127aV:L]_:Ga6;0N2N\@dD?U5]]f
b,a-EG4K.HUfN,;@aYG&:/1_]-[9.RV]-cUQ0:bO.fa+4_#[-e6IdDII(LLTVga(
f&c-Da#W+;W2bV\[Y[1).^c?3@R]=F4BIVPFW/3FV->?\2:cM6VC]^)9>=(/]7Z]
2>X8R/\Cg/K>UReC@\f_\W</4<XS>&E;bfYddIL#^N-^Wfe)R:CNGgV4OgD[>d<(
_IGaZ76I0(8\2bSBR[S__DGg47#9Y+P#eI4Pg#D8BNO,4[e>^YEUR#5LI46]dGG&
gXQ[+J3+O?X#0064)T4N^;7:&Q^_fA?J4K7<J?45e+e?#bSCD)Q8F\4OA)RB2E8_
gg84K?@K^abcE\GI0&MeE.B_46+J_;EQ#SOXZLZG4JM@bA+#7>a\)W],=7WL;9RV
>GJ@WRUaP[<B=->Qe.:1e2+Uedc#;cIU31B\D^Pa<Mc#KJ,#7>X)##5A),55WC_@
XWO9:WD?Be?+fBbRO,_[DRf\HDO+,Q9VW+Q6e\P&\aV;KA.?b3=/1,06\?eW9OK.
MP.Sd)YN]+KVOOKRW.d0bY5__<]L+E4]HT26??AW+:M<Tc=FR&c:J(M9,G02-<^E
?b7S0+2.)c)G>0ef677ZfR>E)RS+7[Qd=f+ZcVB_f+,DU5Na)EKT.\]:b5eZC>&)
XCR9/Bd/N[Qf5+)9Y.1d_.V\/QCWK,/L+=,RHAag3[.+@QP,;]T4NMT8>XSCZN1g
a@dJce&b5\a82/T]6F38HYVH=;0I_S?2,ZWM+HLP74Y:cJ=&5XLT.-,L(6J/Jg^G
FW]8+Y78<V,RF>I6\Ge[B[;=a0M=FFJU>&9g.BT&E#.Y7X>^5ad6.+SFUG[8,&E+
7)ZNMS:GZ;FU0&9KNYS:,&IS:g>BgX;^&NRGcY62AHGVf]4>HB4XPb&D&P,N^W:C
/IOIf<OdU,13\8>L2=T8(ce]6TGWE\(FW=6T@\RQ:SLP/d;2JTfG)>OXZ5G.MD>E
=P(?=3UQ[W^A]=-:0[HN];[>5+6,E_WW[TaJGZ&8HM3LUNeXEUMT+/OQFe+gLS9?
WNK<d5@T6><5DH+GLO=(D6EJg:MMUL2;:Z]D/@cL#JSY9?<=MZ)XN[-f5_]g^fD:
JUN_\+,Q]299dJ^#g\]]S:bG4;59/X+&QX#I)NM]DD<TJM=c@\&</3]S4Y^,I?=G
P88eAO\CW&eG-V+4D1,OaN^<Og7fa0Y.D)E.YdQ.1Q+,JXBKcVN]HMHT3(Cd7\5W
,(4.[M9AM:.U\;+N1#a/XBURN=>V,2VBWH^e;@;PdS<GKG/QZ4@a3JeU(MZ@Z[@W
Q&KKJM3B+_R\AG^,,f23Z2^8?D+:1PeL7Hda8L2aL>Wb:@_ON.,Q),PY6CSWfTeF
Q7Y=0O&1)E+/2)=35S9JZ<Z^,4H1>ZVK0b3DNU7XA[\cC.H>E=c86UAL-YYG\&M=
L7ZVCLKRD4RbL0VFFZCa]GD8&Z.CA):C4(-a1KEVC#HCX:AY7#HH^QAL\>^KCK9I
1=C[X\KPDJ++ENE[Y^GgcHgGOMYg&<L\1e7HCfX1S-/BEf58(/Ic:a+\0Af9(ORM
QdeIb=3d&=H+ObO@;-]^YZ+A@d+8&b0K[HcI^L=@BP+b^bH1[D(4e7O9TI\_4@(L
,R_L5+aDf:V.>4[db,#=]9P+U<P7K5cWN^PL\Od8?NJ?ILGF_2A#H/:,G,SBB<QB
Qc\>V#K5V9Wg:TS\BH&>>SXgI3K?dX9FG?\JS1_c:8P[:E)GMT3]?,]BP;;;AF-Y
Dc5F_WY[W[=(-W=8e\0KKX1)Y;K=K^893U(f-.6JV28+I\GWed@2N3g<6A?3cT4D
.aQ<bJV9<BCL7LTCUX3,)V(&\_M)>0+3B2NKd\RRQ,>eON;BQU[/]1>M/f9d66a-
UDK@>2,e0-_\GRWG)Y=^)CUCd5[36LX;+I]9DJOe2a4<RK2A9Q<^R8-gHQGaO7Ma
L/=>UEgJG31<>/ea8(>WP\Y-bDU3FbDBQC9P6J_-);Sa.28\?MYEAN4K7Y?@:)1G
Wfg-DZ@Y3\5Y++P?NMTIJCLb+#c0(Ef\X4\fFJ@Q[JWc=#<MG_I#:JY6\PRLd4:8
)E+C_<E[WWQJYY7HS:L2/A1-?A>E0,^a2GJeC-dP242-MO)Ld_RIZ<(JZ9#T;caA
cARZ//&:((5F&0-c0E\[]@,+,d.[d>JM[VQ>d#[3UVHD<<Z/VMf+6=TC#AUF[7X8
\TKffS?AP-+B\Q?OYHc(,dPX8fH.4+/M0AFC+Z+BK;I/+#D+EX,CK[Ycf^3M<:?(
9CK\A>7@Q7W]ENO2EU/Z[V3<@:X(U,\f7d>]4FMT_GITQ4XeYbf/;RbA+QBX^<Z5
X-7QG+[8[SY)G_B,)1X?]29[4>\<JPH17#<:6gM-G:-11gESPM)KBI=6=>+/(,X[
\d-@C/.EN22HHg:7#39g&N&OcX0HP]5D=B:JEW#GR@V<RDBEdbIS<VCf.^2D3eLe
21\H5WG0D<=X1H&[TW1[T52RMHa)IL0FDf8XDI9gI2eL7-a&@4\RL(MdbD4#C.]=
c-.M?>/1L,[D>\/dW-68H19QZ/2;6-3cdMS1F^2a_dSK+1V;aC#2(UccB=>JZ@7X
J;UM&7,AY-a\7FTd=#M<O\06JG+:[IN7]GZ@KfUV0E(FV4G#_QaJ<FD_d+Da^c>e
VE_Y=]6=H3/+WW8^5__R>,;HT>F@aXbLF-(E.#\dRLc89;?a-[1bS#dd[cC8+?E4
+2,I-_4?7:RQU2,_>f#.E)7;QSdXT_dD#SOP?&NE6c&CLN^FZ(1D^2OL[Qd4P46\
>6BVQR#:^=.CLI0G_e?501eaN]X-RW&>P1;]O7SY]_FZU-&IQ)bBgU8gab.N[L_b
7#4fTWdHBKJ;gS-::US^G7[e;2#Ze-)]I_WP@NFHB)c?5B1L_GQC20JQ/BLC^-Y@
[T5O0NWaYa^WW\90[R_;NFMK>6/JWRJCB?1J,1eC(6^U4^f(JC<(<Oe;ZfQ8Q113
]gQ(_)dHg4TC63\g8gF6Y2?AI4)U]2aa^eKBPTVO\@)Q3?BbUP(E_H3[>^9A&ZYf
7T0b,S)A_EA3POY;CfV6:_Ma>-Ea:6:fT6#[0bBAKfUW6DXHR.Be/_EH5/=0Y-6_
0<TG)+JRL+8XXRM\\7,9H+a6^C0gFB1^&?]AP;\2H=6MSUMN99OQ7[-+:&8g?W8Z
f\5ZMgV][:))?C-R3,VX]3KGd4+aJ+7.:4gBYY&HdOTNaKOK5JdJ/bA#=7fDcELR
.?:8Z&ET47_D=WT@G:SWcU[U#@7gH3S>8[-d]Fd[C<@YWg8Gd8KPWZKb\cMN+.6K
a5(_0eeBNd)LIN#G4Qdd=:(M4ILIMa,]N#>>YL0OVf2XC?,80+66Y;0AX,=TVg(Q
-cP>[IVR@)#7D5DH&5]C@4e)?Yg)0HX]F_?V#EU8=#1cCPa^APG<,>>AA1@A+61V
&EH;d8)(C6IU;&GfG,39P.LF<?7A#e.&b@>Z7P10US9LC^LS+O_a=WfA#]-\(eYU
^S3::Y<(gN1.+Le6\6+PHO2,F_Wa;8V_7-NCI;VX>_9B4[/7<.6e9G[LePOa9Z,P
cI?c(X;PNDf&OYC82+?R&-0]N,OdG,fe0\K0+;Ub4S1L\1-3L#5BL+#5HB87]@b#
NB(_A>+Z+RLY2:_EY=cNKI^EKd9FW1NC+QNNWQQ_a74\/6X66PXY[EfDC\2206gP
dR[fDd701.[\&NPg&O/(SP@&4#L<SP@^7+9F[?A)_[HFM[<FbU,)RNaKJK7W^-C:
6VAOUXYJ@9.D@S#3XG(_AA;[Qb4?Q=1FFP:\.Z^,Xd&e11I)U;g=0)c2SbX83[YW
R4=Ra362AHGf6FJF6:FF)?):W[0/^30WI/]R9S6795V8^9d?>-PC.-<M2g6.^I.E
4@f<C=9.#0<VQ7D.98U#K/2G]f))gZcS7GJR-.MB@<Q6\)]NII;OW0V:T<cBG:#]
UTVbI1e3]TC]Bf.(&b\RGY02AR+O:DdOWIAc#JQe)eF/R3a-daACKX9:_847(fZe
\K15LId?+bP-4H0:KSL[g))>(Q_0=MQbI8_9V]5C.]_T,B)3f8LJX_KDCFIJ,A\8
1ML6\7##5e>ZdZ;>NOZ.KRBXT4?Y.5<92UD1#TF8CMXfD]BdSJ\E\e+<3&EDOeF?
d/=+X7NZ#QD?g8=9RVK@Y5d&9bO6DY;@<L2f_^7fOU=WDK8dZ<OS4A?eFF:PI7\E
21=X9)M??6E_@e-Re.]KNE^L=eQB\PaFg.->PSM;2f_:g1WY[De-[cE#;LJ]Pf;,
V:GN19ga+)OH,B<]CGI6VFJ\2KA)TC[5VZbQD78TfX6aQFMH-+b?XQ-5U@3IVJF>
2^#9JCXBC@\Og)3X_E+;_/8_Y.bYY1+_c5cLfYTWXgTECSUc:,bW?:2]1P1ATfN0
X.WAbG/PW1[/de23G6PE7@]JZ>EJK&Fef,]_XK\4.FN4XU0E]3d@2GH3FVeE.MEV
0:ePNBVS5I<UQ]?_VB#eJ^AVHNP7,4^@&+1Q1,ZG/L+7&7_:X<G(NQdLbWaBAF2;
9;V\PJEd[Q@cD-:WB[IDfK@F]2OeE17\f76Q4GE<LJ)M),@G_4E#g/87.McC>#)E
/\VQ-@ScFg=J<5.K,.7HU9XR.2@N44c/ZZX5WHe?F&P?f:B:7+J^0c#Q>YIY/Ac_
3Q<dR7PMW/D^,=VNE:-a/WU/4EKSUR[\Z=b]AV(FFYI5]SK6)_#JE-HEW4PU@KWT
2#[II1_=dL6OL_-PA=(c_/_/B/+-+4-\3>XF,Q\=:fRIB-BN&I4UWO]&[#0;TYF4
_6ONT,)@SGA?TE8f+BGeYF-eTKcJ\=\\D#&O/b0d6c\FV>X]Tg_b6O9Ka]P?c[U?
^4F1VOgaDZ-=WIgb>d_06?#8>JeEO#PP81HZGC/41KL6<[-#M=?ObdBLC,LLE/de
S&KKW>.=eUL8W5/8A<B84)/E,)0>V3Q3/C,=\8[WOUI?P0QLdJ^7C]72Z.gQ)VX-
@TP;1-aBQ9(-P+]NX^5ZGT&Z[15g7)dbJ#OCSJ8[/O9C</:(5R#cY9?8g;9)J[:F
B(-U9+#J:H3714O#-g2W>#HFWID7AL^g)K+3eWWU6N84E0J([/(Nf=/K8YKcU])c
=G?]Qc)?2f6G#V1e_J[2QMgI6W4Cg8:XN(;Y7[)\\W5g.Q/Z?O/;<Y94fIM<#aY>
Ma86=3N\K:L4CT+1^Q=,IV.f[e[^Nf5X+dR]62K#U]K4@)6\Qa8SNAJK6OH-cT?,
+O^B;@>YV&P-QG#63S+W.9.ef8P]LaJ7.Y9^BLKY/-]6K4D\+#KW;MJf;bCFLHLJ
K_270DR;bYg@Q1V8MC&@QH?DB>NTg7,S7R8C6FFUTSJBYQZ=_Fcc&0OFP7c)Wag/
T3PQK1R#Ig0E7c);3M[+_JZ@S#&KYPffVcTSBC6Hb/XO[<OUH&E6MT)4E(J</G@+
5A2UEBUUTg#&M:aG^@O07c=[:f4CbCgL\&G-8>7;I5D2/-SL7P;9(JTdcIMSaYb5
B\,:83G=^MH/YV/UKT0d53O=YfXS#[MHaZPOLS.L&)adYM2ZO77[ReI_U0P)gf.2
Z;1[)#CU[EeC5C:G+W0gQNeJ1ZWY?db0SXWWAB#0B6Q1XP31UFN^5\PG67bZ+]?1
HBRSc&aZL05:RV&_&-W,V@PS<\K\&1f7#deM_P2d];Z-4L]H[_AFBP4Y\B2Ee(a2
M#S;IBQ/]c#++-gW/]P<I3G,C+Sc8\aBJ>#1/5M0GG3X[7OZR7C]TA>;=&PDM([B
PI/1O.cT\H)/MQZ=Y0<D[IH#_&)=5/O7M^>ba9)TJC4QPcCUb=.5?=6bfaJbAbd?
CU\g/AVUDN/J#R1M4MLTWOMEUX5DPWFZ0)7gWC>E[R6E.BMQ(]bRW3.03e[K3>UJ
U#=_C@39=R>-,0?<X_1R?Rd.HL)@O47fF\7HRZVC_/D>E=R=K)R>Y>1^9cPP+E#W
_?#B[&B]1Db(R;=D0B4XUFH>7)dSf]]eV2/5Q[8W\U3De7gB[O@@:55A6gc#.f]>
@Da<6CeVFAZ8:XY;cQZb7F#FYKQB12#1OL\^S+M5K]^KD9NPJbf?=UcP]<JCc12W
1_WAKfD9C.WEacM(\J?^,2)Zg8E575=SYPE3T?4_/RP:(E-)@24-]O@JB#I9OUC9
(Y28T33CTPGB67R49#M\PFG:T.?^1KD\]d:@LF&,8M8Ga0Dg&\f:3MPNbGQC26+d
(?)G(3PG9?bb]e2=VSg0G=I4Q7IAZHB^057bXX7RG^-?;EfLBU4O5Q]7_-MCXOGf
259U29I)f2./DL__U&@:M^PTB(<8[_RD.<dgcaMbe-;=BeZ+^UJ8@1W(=BR53MM)
H+K<6YDC?CUg[PRVa.6/U:UW3?MJFHZ)L?ee9.</ef+9&Yd/]g3Bgc#Rc/BE_IM_
IG..PO\FU_>T]7ME,^(N/]P6Pc\U;EM>eZdeL_]5^a70;NNMP7TR)Q156QgQCT(G
/ZWN(M6-2/,&X;f^ZFF4741cE6V#AVBA=IL69ZRF?.Z=HDc(8#R+,VCI\99OL?bJ
deF8.607&XJ?JAgVM);0:HH1eObZDX[f80Q&1Lc:2;+DO3_D5-H-gX5I^g3B^:QE
L#X)f;@O0d?0gD[E[(K5:Z)?.dU3Z+J8Ha0-<#a&<R6cEWb/gU5=+PDe_6N=f^GP
QR=+E#&eZEY_<N96O#F>\S;WG_YT\P?<cSIZGZ\&gU]@\?.<>ISJK#gfI#EN&b4B
S.#R(QGE8JeT.[W>C1V-5SZ:QebN^H?HIMEW0Z@BEN]b6QS(_O^>GRM7dA<E3W((
KEHUFG<;b;O&ZHd1Hf&d9NZ)bUX7C9I&(TgeE4N.X.##)X)c:_a2WP+(MCE9ZNCA
dJec=I58a14>IF.4a=58B,.J(7-VP83=b=8d9_IaJJ+Fc6D)[de7Wad?<C8B&N.L
-3Y2QZ>?Y^5ZZ,J3S5-6F/-KZ;=J=c.cT]?VRTQ\-Yd<fAV&Va7>9^]/dD_NDA[G
?8ACQA+T>?)K;^CcZ<YLC61=]XM)O)JF^SHf4&XLDS4?GV>IOLU1F/3f90,aCA_e
PF]:d:cg?7EJ[<KeFe\UU@ITM3:La)E,,#C8Z4D5]3+OV>b@/=LIM>K0+Q\CVWO\
2FGC&.+?:\36RPD(W4;g@JTY/>;&K,>XN-g/EOY7R-3XQ\+#Sg0fDJe0.90AH.DT
GJOSg85-1dXI5>:/,;08^6:#M8L@egWH6:+IYFM&@Hb.0GMKN(2Y,]G<;K)bL&=_
_O\a=7d[N.c@b#E([B^GR8OF^]W8Q9;ZK>:];)P:cU8-Q@KMW#13PZ4dJf0X>=aO
,T-_BBAGS;81F+Y(F9/?8A6QIYTQaPJgSY^UKccY_I1RTM-f:=@e.43X;#/ZH>c5
VD0K\X@P;4Wc=bO<D(VHd/__08dS.8S^QbeV0P12Mg8/V+9b=EE(]=W9a;=DI>XU
/5E?YU\J\YOGUN7cFJE\U0DdU^NO5Vfc-b9]fMK1^eY>/W1?LJ?W/K6_/;&?7Z>,
-O4e&F9UO@GWcdYdeL>_\(]Ge^S<6Oe;@W2III;#D/1G&^I>,]<NV)D&UcTAJe>-
(MgAZfK;_L8B9aG+If1W3_>@<DWKa8O^>:<]4LA\Z#ZMXD#8N&GT.#\R<.(Z^Y]7
c:)2cJ,><=N[X2bf,60.B>e#NNQFLf7O3/MC#TP)GAc70D8F=,D1c:=[=2)M^N0K
Z2,5T_G@\=+fC6#R8X,Z923D5-FEg;/84dWGX8C\gaa#Y-c-AM])>=_V@\A=K1GF
S\bf4+?;_ZS/+OV98-CgTbR<g#7LPL<6(:edGG/3WN2)Ld6>B1^fPE);)>f_:e,<
CU81E-X58]#ECe3\NeP_<KCPR(6-2<d]gfOEbN+Ce[68MQ-[,dHE10UC)YSJ91YR
4Z9))T9C4;EJ)Q]>aB:fW.G.ZT3QU5]fMHDC=\-Q.KH42GJ8_43[RYE:N&d>E#bP
13UZ-;R^LeF2+U[^QVA;@+78EV\.4fCdRX[-B4#WY(_(c-?(BH@.WPC#;<C;\;IJ
aK6JC-RCPL2W\^LY7V@/</==CG\5OTLXQ,_.d&f4LPaT>3<#^46BVFc0RGg(R8ZN
Z8g=Vagf7<.&:^21XZHa2I4c7?aMf+IQ2@_@VIQ\9e7)=13bB>@7W?J85J4P9MLA
?2O\=8TM-N^@WU=35O8g8SH-c4]LB8eg[@Y3][=#I;/g&WYK)BG;#WC?\38(LG=3
W5P;KQ/]Z&W-,V,U4[29cdMG^G?\eQIHG&?8::.]c4,QPRb7gSEFAbfM^aO-,7\O
[Wf,D>;I+[g=WK)X.L[ef;.\Qd&^bQ2.Vd(8-4daAUe)VZ?21_BFIMZUN&Ba)BPf
Af#R#1Ng-EC3HRLI4_bX7FaHIAH-;CXJfOWXUM8J0+A2L4G_0C24.fK&\T@DXH,\
KE9f8TY_G>R[9SaWHAEU=/XAVI&,BMR,]0-7T/AZ&G8K;W=8.Q8AE.ZfDS3_S&G7
^X=9PZ?GO-4U31Q=+B8-Vd1L_0UcgVPaA&93PA38_?I7RHcQ=88f#RPB#DP1A_2g
aQBc]2EM:gAbPM746[baV)&F@fa_F7&(A@g@,<fF<&RcGP>R+[aTV4(.UV_MI4Nf
VJC1]@GHZA_D?b,7W<?ZW/>>]SJGaCEf0?E?@d&D<51_JB&9SPeJKcZR/cFK1M:,
b0QFa6=@KP8N(>&TPIYS5/ZXF\;8.G?\T=P:=?-@V3NBRA2Y#ROS^-IAeaD>TMb/
S59@8g2Oc1MfEH8[1/eVS?(@GGWW[?3I9M+\Xc?BI4H(-WC.dCbL(O\]3PEQHT.T
\EeNced;,9H&MI?1cK6W;bK:B=)MP?F6+Tb2cdO6V.<RBQ4Ib@W+.c(E2d3NMJ?;
>3UH&@S@1#Q2VVHeG/>[XNZYA:WIJUHd]e9IgDI>Wf-6QS<-WY-[@XT=\@ca8=D1
GIF1SN^5BB6Y/4ZGL\2.g32GQ#<+OCH6HNOIC7R/YIPBD<]/&9Ibg3M4Oc)IeE[P
W(Q[_9-XTZIKILeTI+)O/9BBKU[PKTNcX(DFa\O&X8D#Mg:2N)M7GJFbe\GWgaO]
,V_8>.-AJ>SOQPf2[TO--e_,,__8IN2H,gVKZcDW[9QVcEDY<@(>2>W@fABMWLB^
9GU6F>P5O(S^bCR]d/CY4]>af77+:X:<)Ja8a<J3FfYbI9g#Se):X4EWYSbYVMSK
07#<=-&<gVV#T,[:b4]Kb-ZX4C=XAUDW(54I5_J\<c0D8=N#&3F.8=I[-BeP(+6<
/VRT;J-Z)3197B6_P=8CCI)(dM(-a6bWfC)\X]KeF&@?FQ#:bK-_gJ<XDKU,9;8X
@W#c4N59NSI;.,=?Qg4)@U>@&I7BN:T8XIHBTYD)43_3N,J@8RdPH8-):&DU8G@V
ME11dD\-(?^,7=b;KY#G9>J6,[77eOaDCD<[+_B)0LL1c\d-6BT-KGG--gDc=]ML
E\>=+[UHEHG0V\P;/+LF/\IbLWgYZ2SU&JE+9-P2DZ&6ZO3#N8?(eHK(SR\G<87g
f2=^]b&L+M6XZPe@3074=Ic]VKRUNFHPV<[;4CSZUe65/:O)AFHHBG7DF-f(;Z^0
&A@f9a(e,9T[P<;c?+)<KB\#M5Ob60eT9O0)Wf4R<2@+=Ee32,.@bfJ>N8GIM>9_
ZS)cM:FF:]G&7,EKTYM)=.=/\[,@-U(@QO@Z);:SU,,D&3#>)Y^4G>6+N\B_(YWX
17H;@M:.W]&<<c8)QY4B_@O[a<PAS;Bb3bbPR=If4F9#e9PJFV=g6\#TC/FV4.L#
-0WS9>PCbb_C[@J[,_HX:LP:a/a30e<,)c+F)TR?-b5T3-gT<1G;]_8[c65=LV7\
e454b(d9E@OF(OMacC/(dV_56X]S?YSP5]d8b;XN_DLDfX1M[T7O0RRg#5cL^Ba@
<X2F;@V(VQ+b,Z&#CC42FGP=Y1K9#c59C?7SdGZHB1=#)2TXJ>BA^N/6X7_1&1YE
e.S/FTe1K6,;]@/D&6DRC?<>9(aSDJCOFH#OJZ0#IZffLg-^EBd]Q\S=Ac>P2]?c
[ZAe/-NZFVQTVR&/ePdL.c:D-P^;_])7++Q^]7BQ3]O4Gff=S(TR7@/E=T7:RB5D
eJgMZRNS&+G/23TKe>PK6#&;S7KV7\ET:9A-IWHfV+@8Q/BZbY5IM;6IM<WG]<M,
R-5;/+Q8FI@+JgX6_gOF<P,-;6(fQP^ce+Y)@1]3M1\HQGSLX/IL3aG_gC.g=LDZ
/\/;;Z5UDc?;..</)F)83-&-414VXfS->C7a^dWFV<6Y)^KSV4G871VcNNdW6]#T
_/QG1Z_YK:1T<XUAJ@D=R2Fg2,gO8Vd6AFQ<IJ=OKSc<-DN1OZPE+UAGb+NATA_D
dQX_&-/4\H\aDf8,KWf@+EU1X/&>78+L:fW8g#W8cU=<D1M>G^gBMg1(YI>3_Rb;
IBUTV2U>c/dBD(M@Y^#FW25U[)Fa)6[T/[W@>D3RFA52E6WY28b(g?aDP0fg;T>K
Gd_)UKKG84-7S_JFB-R6MXCL@:.?>.J-PbS0#@>(aX/VebFU[N-9[+a7>fNK;^:/
]B=5@4e8LG74<)c_BFF5J1PK))2RS^fSR&H@a44]e/272-f&VOZC@YaHe^;EZ&d/
L)gFJg,cPJI01&@BOE<19)(I137_?>.HbQ),7K.CPg6)#5Y94HdKEEJWM098/06?
cQ56eC+-,Y./(2.7[7ELKb2;O&0M5,.<(?^AFRbM&_8DO;-G9VC9V<c?QeFW10H?
gY32b/UD0e,P;28B+]D7Gc>.N5?a:6N<5.OaAZ,0)9Z<]d^VD-L\#3:IBEe1^I]_
P3L3X-B,[JN9_RgE;,Z(D((dP:U[1WQP^,T-HeF;?Z]F/QQATNe3Fb>;_C?JSPL9
VA_LN32UCK3<L6F/U,H@)+W<<g4)_D:3J\O#R/B]cA,:+gZCY,(7+U4+E>QX,D+D
P&33/,#K4bK_,JHQLQ5RE-^SYC0^Y[,IBH?(;FTK5T=^#VC66R;H&8/6c7S<AT)(
KN2=4,O->:266.C8-/)GFdV@:EA=ZR/BBgRK+VZ<ID1=F)cX;(BHgA+\b.+#:NFa
A>Ae1>WC_DaG[EO_@Pc?9;^(F-eQ6HL&3^[N,L?7U=5U0a11aJ@>R/;BMaU;a04\
5@<LaBNVE0^(]P^IH_<e]A7;Y4N#TR,K,/853U1JB+A;BMLd4ERge&6SZ0/LZ^I9
+caLUN<[2\+G;DgAOKfP^8>8@,=O.#Za1W1\_M89(9eT)_)+833&[cP(6C8UQ/2Y
?R;&7Lf^(]:_Jb8gCH@?8VR.^K,O]dF8?>a7Zg0(-^8:0@?D@FH)Q6GJe)G^]@,G
N>6J^.]FBJ5.,2dC:AHYKfYA,3K^X.gCa7IK\L&1S(>&Ua[YG-C)GG.;Bf;3R-gL
aF(4&H[12b[(Q6683Zf7Xcc0>9LPbf6\CP-5Y/KF=[,eI^TEHP64O?JU@Z_FX]OU
#K9B#SQKQ)/b_V-V0CK\##EJGN:4Z(0=]<faJ^9UGebc]QB=0HRVL8,JG-:fcDA)
68Ya.<7MJ(J&0W]VNMfd9_;J23DQR[08cW2:V\T^Ze5Nd3C;?K=@bSgNXK=S]Z#<
J)&A.O6;HYbZZ.K->)G,dCZ=90K/&<8Y7[3<7gB,.[?S#Ja36GgY=V)da:Y6U_R6
&?(_\J7Vd2(3@)TK4IMT-KeRCLEF8VQ\(d=HBU2W-F,MA483&._]CW-3:G[<f^?Z
KK5KW9KMX=K7aGa5&bCX\T],6:eW3,>4]MKXOFS/+AJ)S3=)bKT6(?gc-T7>@+[]
M6]P#[#Y)OMV:;8-+T>g&F58X6bZDJL#_[Tb,:LeCDKaU\\4-9UP-CdW0FH,^Y1+
/=>S@Q)3,R+?bZMV\NL9,N;^6R::==F&MFX>MeXQHgd;O0G<0J[XKBD,,N6(Fb=A
?>_fZbbO[V+5A2)RT9?HZ3=U])RW,#)S7BR431g+gAZJ19/[9HfaU^J-[;<[DA_b
;O8C9JR]/UO/<YDe0I_B+JP].]eg0R@5S+2B64IRS>f](5-5/;+@D)RUOMc.0+\V
aVS_J+c60gc14,Q,)G6,WWN)a6cG\3;;+FUb70A3(>.BYXC-WCR&1g;Rb;LN1_RO
]D;aE8<-)Wg]YLLe03=59/^C9O_;6ZGE,.g-F@.]b780DdNX(JMd/_-YS.IMRAQ;
].S[\P&]9]9#UIK5G2=>:DH/8W>FA6YGY&>FQ@T4C4G]:M?b3gQ?)/Mf#/^aV5;b
;dN2@d26+#8T2Z58C<L/g>3e;fGU),<=V@--X-^SA7/.O]g6[dd\\g7[=__.2LYB
c:fW/9dc]#NZdN?M-ea?+QeZ.?4ILF6/,DG;?UCeBQ6X23eLOHf2_eD--W3,X&0f
3Le<1:g^S1LA?MRCHdA^;MC98KV1U[<e7cFKX6[UaT3W=>;USY1N.gPCA&dW<,@B
29ZO)4?I;>G_08)J/(.)?1/=Tc?VP[G4]6,+BQ]TL-.1Q.Z8,2(WcSDAbbH#_+A?
Q(WLWE=>>9BM&U=(F>Jbe9<+3#cMS/gU6,Gg,8MaFH67&,7E6^3c+N/&-9)SLfaR
ZX[D70(@0<^c,1=.1;,&1RC@SBV3=2P::4#6Y=W0FK_VE0Ja:JQMY.;c-<Xc/B34
J\LQ6)6@4RN1WIE3R;M#93&D6:^/&XZ.4D;QD7a;a#9#^@IT#LP,P;)ddgGbaHU3
e_?EHa.TCHVE#JGN\3/(Z<)^9#JN?\N+1\#NQ=7?TEg3(QW8;2?;@Q(c>LGW2:W#
]D<,:8=_^/^:DPdT3=OXJGM82,4\eLdMXg]O]COZ_.57_RG,]^3DCb@8ad24e)P,
I:#U1T/e>K^c@XA&SB6d7WMG6#><da=dL_U4X66-6I[@H]EP,UfX])d#<U73B=KT
7a_1AQ_)Ec1)KV1eS8fKG(H?Q#FA-[ID#X@01<)@26d^SW>Q@5,77[0=+2Jf6,[N
HZUbMf-EZ_EE\QB<=.2HU3KbX+3Ea(.X@bgc_L4=KaT^AFF&>IT(QS<5YD7D<?T<
X^20OP8SDIA.HZ8.-8<a2eKE[ECL&KS#LX[;)_:0O_QW4QL3_FI_2=C7)a5WWFRE
caS;57-F.Me]+_Q139]?a#DGIENf.)Ef_Q=3.0?IIUG7Z,Og30G2B-3@(CcCHcVI
XP4BeZa:T.K&\6C7_AXV<Q9[TQNCK=e=?_Q0/)dK5TggcESZ8E8^c[PJ&>a669_.
VNcJ[ZXO7WCc<F\L@=KRY?Qf6OMG;56Y>FHG,[4BXM9R/dN<&2dO0BE#95/c4:e3
PCaCD+587=aLQVBS#D@O3-g/S\H9d)/LZg[2<a.GZC^Q8R],(,^OBGYabYeR#(Bc
-eP;W7(_<)==<\Q1a<O,ffKVJ&Oag3\TN8])+gBg-SaN^WV6V=>3T-]a&IV+O[-G
-Vg(f-3P3fM8d0ZJfSP,31<0@6XT#5\8[^S;eN&Z&8Xb2751U/MME-fJ?N@=X)7-
#FI_GT=a.Fc:.H&]_K8.1:CV/9VJ1W).XHYYE,f-K7BD;CLDI[2b-_ODMLU2Qc))
KF8/@E6SGgD=XK2gUU9O:(UO[g0Y_KN:9,D3C@;1(Y:f.45Y?C@c0>(8/BM/<54;
2)SRX3Pg)e)6O1ce\Ue189_9e4[6P2[ZQ9+CAc-9O-^f3[]@T1X@-9.QB.20C3(T
.HTOQ3VIDK[+-L;T7&b-:_ZFMce:H5cQN.?_H9,NYOZ(FeSAe-7)b0#IAZ?<Fa^g
>/9DL06<=^413>BZXQa[_CP#-)K&4XQWJ=2YT(D@Ca39]ZC6aDCIZ.4+g<e-UR@A
3)BA60bKCN_Nf#HW1H:@GK4S?O/]ZKOb>4(M-^U:c1>]d)/)gVA#SE]-Yd.WMK_E
JNFHe<(R/?_#STGd9AE@(AF4K;X)9f+S/:2OZD1Q,[1fEG6b23-LF._HXf-<-UEB
g(N<BY0\4&ZefQ)4d/Hba;\0M3<P)O\3>)Kf&)1LD6#=(;:)EX3g3d9D3:N6c>4c
^0SXfW3MW1G8/?)T[>:Y]cF7&F4<?LU6<^U1#@P_:SV(Sf7&c,H:<&Z]f(6PNF)b
?^L4VTb=@3?J3T--d5LJ)+M;2Ff;6Z>V[_<+P7R1:dI_-HfMZM\J=2MRc>F+^\)c
c@d?\>bZ#LQSPTbA#+ES^>+]LDN&/R/?NQ830>3fRB4:6RddEF(0f4S.@DMY5Q@B
X)RTd<GLCgb^2#bCF;cVAO^,?N\[D[C^>RS2+7=3[]_9g2#K)OSC/>AIL=[;)UfT
YH3ZZ4K&f]3HMQ/Q8L,3fL2d3BICI?3/fg#1>gUH52(<eBVA2Q[D?28WIa6C@F6>
6eST-G#^G<(_LQ\PSJ3f[]6\VQH5XUEe)[JCX8/Q6.2HOba.B-@QP2X=X<Sce<&Q
P5Md.&VEWb:(ZQg(4b.E80+R?6UD[CA>eb=::(4+;=9_1O01WbVDCK5XPV)1W_F&
BDRXLN35MT^<FX8-BV>AN_>CY?JXU=W8e8II2=bc9ZV3a)/BSd]N0]V^c4^+X,cP
YLUI(0_2QZO)^;.G-]#]840VQ3b@7-bG#K+6NT0DBBf]+e;O94IXSZ#)0K/1\WCD
-8(Seb1;O_e/QD6Y(PA\ZGS[[f,_L;[>[c/BgUcVd#>SAN6X++/6;U\7b28[@ce5
H5\aA5P^/BR.d8A@Z93^\,_F:H,W\Z5J3Sdg^0^D.L=ITB;,W\38^P@WYVS#5Y_C
4U9Wa,bS;5ML(?I+##>N9Kc>F(81dT=C4GEgE^aa5L50.:,0g8/[8ER1L6YIJ_Hg
S4O<@KCaOf,1<NE8aSZd:/8N[4@&a9TeDX(TaE7\I,LA\3@ZU4L)YX_R?\g]ef<?
]=1]V+>G[/Y49<2DHQg#?:P>VHfMJ]]fHPWL@YU<B)I]E+C47.3/1\SBR=4/f)[A
gY3^H-S#E4O;^+Xg=7PR04C5>)_6.XFDEbNX3g7AKB^QCEYeMME.gTAY9^)/,Y1A
)&/a8XQ56\d&I>J_66-XG;9O1Z-GZ776>BWS3[_5668UD4f7@aNcN87d:67D6<<B
.Vd<&ZV>[?aR&9J/BG;UFS+BeM63,I&)XR8O,)_,E_/NGHV,+>5<3SJPOZ<(^SFW
+>f,#)ce3Z-KGSgLNe>&1K&Y#@<-\=CA+D8@McM;/W./A&MZVUJ;b025+/?ddW:3
AD57(3U>8SfLLQef\&LYQ)I,F.;V+Rf\>^()?93OF/JJL8[\EL@7DX4,aPN>)eL(
JcOFEX_GM8^Ec,fPIB1&)fX5-+9gGY,_EAG#[Z3f]JQ#;-<L.eZ(a\KbH2\+QAO+
,&@2/H..HSJ/YYd=J4)2:)W&.B/)NAT-fc<46XM]@Y<:[WR^?=P1RO7/+T#\QE,@
ZZVUc)T\8E[NSTcPYOLH/);I/^AW[&GbT@/2D328V?dfA&5YGB@:(/9E7)3[1FTJ
.WbHWYAFJ,D+4LL3\FC7CA=EA#H<R&3UReSPIL=WM3R^A\9[gJ?7]]Ac,2.fE/XJ
W,T^)0SJ9A0-U//dAKT].5(\Q]S=D,ZaY[RbS(<1:d&1e/4IKf8=7f[_CP^^8V^>
dg-\YHfF,ZF_J4aH]](T(AB-Ae:PNZY4+b:BOTJg8K0T/SCA)eL,=6D,Ed6I2;8X
4YC@e_BMZ8X,-d4R5GFMdNK2/CH&eX@L1R\^c9Iee&Z<g3<\9e?@OR7CZ?]6/afQ
^0IDMM](W=cXF[D(TQ-f@@JSQ)G,eQG8-[BRGL>Zg?X+XXP=]KP#Ka1USJ5eB:;Q
>/Z)\LC?I/.Ngb7F1d]\6&,XB?;SK,CBD51fUOVJB09P2SVP=(KY1#B(\EG^9O.-
S=5S^4EQA;IVU8G-_=4H]5_a6(1HZ?->\54Q7WfMK9dKED]YB6WH6&+Kd.?T.Y+G
Ga)KcTZ-J:C](bW2BfdbF>HY;]\>-[[#XZ;bZ-F,RQ9(PdgaPD=A7<].GV@X)#WJ
OXZ:DZZG\dM3LcWgaLSA>O3HdNDDHJBX268C(62DHB@,,<If7I3SS8+U#KUW\fTe
:2cUVf-R9C8HHB75#6g[-OWKfI\PR-A:4c=/>F&.X^U[^.X?:8/eL3-ONW>=^ZK3
gIagDAdXZ4WANbYeELC#?78[(DH_;CaT:eYR.5dIJPN2C3<TJ[2P3WH-c9ZU]DG-
OEFbP::@b9I0P7H43>[C(Q[&,7UD1IU>@6UPY8LDYSM]K]6Y<=\CN?)\3)HE#]:a
7Z0[[#SM;dae363U4+FP:N[_+K.e/O=PAFOE);WEf40H;V\=;63_g)4c(\JA#EKU
3fI-3_=UQ]>9J[:HX\J:P<0Z[=O+C2AR]04QeE.J8ccReZ6,&N](&L<XJHFL8_T^
aA-HUVD,bVK<0TeaYOAEQ)6#M_2g>GQ>Y32F3YaS=-HD(bY7cPFT95P@:#\)_N_;
BZaS8/R3@GI3Y-B(;B+10df2L8[cYXLKScJVCPL:;,PC1,F1@61QcJ92B;c3;S>F
V\7cS[QZ^@3CCM]/fY<Z</./J=0>IMcMgMF60O3]<Fc6S4VfY.J0.T312[bGgS5(
0/B/J=g361+)<TLGNgR9fM(d/=.:_V1R>5G84S&)0YYF5L75e(OdS^OT(bX<N5^-
FZ)7CE:,[SSL?\.FOJgB84RV+cUM[,;#R?(TT#@3Y>Id=)-NXUE]-#F.[GW/bGI-
Mb)TM7>&f&R#DDgNY__F<#W=W4;3))M6f;L6POS+2IaW_ZC0=1WfIb-K#C3ARf@b
Y/d\R-&5R;g1X7G0b-\TS]H]MT[>TbEO>OdF[FJ[&d>MeV=<f3J@46YRSTgW+.IU
JH[6B@L+10<S_#KRcA.)F8Q9MXfgM7LA?8&ad3,J=O_]Z(Z<8Y\^1_:I>?)P[&[f
NUTU<4:La<a2V]6H6UOZL9\XD>KUWgU;[Xe@OX-1KYM;:G=,]XN:.26=[5SOKPFL
f[=)77XEWOD?g]YbPF3,e4Rg:.U1f[F4Y?L[G4&0HXX2Y9/H+Y[7SHRg/gc;UZ0B
M4+cIgKe1fJ8OC(baGQ[JeaaBSE66N)#[JJY/V<5fK\29TN9F^=GJIASY#(&3LOC
QW4M2WMB1+9L>WF25A6PKDbLF=36(R19NB-H.:G^AUgH7Z^J38QYReDO@^4PDeMX
/V311AJ[M=:T:R_Yd43:f&K=+1Z4D.O6UUX_BZBgTG1,=49+\dbM?/D/[YY7-O+^
b/.PQf@d/Z6K8[C&7MST6ccb+GgG?>aR;EE9?P4@68WMbWG_;.7<DWbG@+<BQV60
XD:]8O<eR9F&JU>HFbf-V(#[2VE0W5b6gYUR5[1bgAVCe.)eF3DfA)E:=XC\NdY8
IQ2FRJa#>SWb@O>5[d+_H.LFHH_4(Y9SK9bEfVV+J5gW&K6acIT?dT6b8?0e&)_S
83.e6.47WDP)4Vb.?dJaAdKT<&]Bf4D1/_=1MeJ6?Y=(7EIfSR:(^.Ia32EVH=SR
O,><JHa.f5@agC]GU?GRL@(W+7#J8OD^9E[V4TEQ)0fQM8L?GDZL7>8Y7;?#ZS[[
+DSS>EPga_9V5beb+_7M<+g6N;V^aU-3ZBWGgf771EBW;24H96RH.JW9E8JY&QCU
ZD161?2<A=,L_]\FBIN[PZ6:&UI/HKJ]HbcVUQUA3)Z<:O6G3@&#^0&&dJHfU@@4
/G4O8=[C>TE4E&2>TV@a0NY>GZT7)>GPH)9038M[bSPa[4QZN=1dF,V(RMY5]7-&
_8W5##)RE(.7f=AO9H&;L4KQCf(NDJ3BQXc>Vd=0]VIQA5Z.>CQ-/.SMO.<S?DMP
U]H^T:dB#D3?<Tdd276+^\a45d,K)d\)1:TTJ(BT])c_^6IV2JU?_0f__VEI-g3Q
bT2^^HM^b@ENKY/V6+1/c#(Gg#N\H?NG=P?EfA<3Z+g/N:+/3LQMe/)3K1<A]_Y7
)HT0e#K#BA3].-Dg>VN4R^<)T1(\Q2()ZQ>H]UJ24Z\;bB29SJQ6C.3HM1L_VP,3
^UD03ZD]/J-_[DLVZDaHQ\,d&:OI8B>DT7DZ.^^KMS/^.Y\<4Mc-6/.7135:,Z&:
eII@,K1DS1?3(<c1U1847\]0T#&.[W]]:I^Q14=Cg&Z@-><Za@_49<g/:,6b^0>(
+XMY__Wc:=#g:Z(U1PL#3b1;:a0O^:d_P7P#40E3B0KI7Z5WcHZ02LNc,^7)0WX8
9^0AaO)8?F?V7a6TNg6&:fad,--LJDFO6-LW9^CC68HZ?ZI3W@7JP:G)S&4#Y:P,
[]S:BOQ92KGX68UUSaOV+HL26\F,IKg6bK0fQf7E=f/DB0C1L3Y9#ZU<PQ&(-.+G
>L=Gb0^W]6(9P(.(PO?BXF05(Q@6=U.6J2f,7P=H,8#Z;V_5>G]00eVTN7\+Ef(g
Y@4_OL3B5c8)g;V3fB/G+STO38ePNFQ?AG42Ie22&/cTAS3ODfXL(Q^\F\5YM9/J
UdH/VJT<cLSX?MV25,>Z/GdKR7J+dIAT8F<M[,,+WYH<_dL[cW^7Z7/A9<JWAgJ3
U1L,8a^HL55=(+Z+X)#\?.WXWB7VI:EMCH4@+W8>cI#NZWD>T3VV;7;_:HLd\eb7
H#4I#A?XY(F<eS,f<bW:EHL7E4[XIO/[H@LHP@/XZ&^.:1A[_<N=T8&fegQ?:6(K
XCOGDA46BR4QCe7;gU5UXc687O)XEVf-=MF:F>/4fC@4N+08Ja;]Ba0,@EV,<31Y
@SR/W.AT<N4ZF2)&8?RY,EXHH-0&M+dT3GH2YA7,:HV?9+a>=LPK?]f99/0:aBf(
d3e#YS/-<0S9#0._Z95C\GX];@A27DE)K,eU_ReeZ4.eJ-Qa-23fM)Z0024=DPUg
1M.H/JVcX&PZ[-/10N>K3#ET(b?MG0@S/aW:YJ-I3+9R?E9QP#>1Se5DfJ.eI9_L
_&:],QU8aZ@AU.BC]4LE;+c]549WT8OUI#gKcR.JEQJI(L2EW0:^T4c9P_6P&1#B
b#J<Sc,c&+[/d7CF.IY3FfU[-ON-WcNaM:LX)\T>M],N\+N@BYMDMd\/2=[8I#BS
LfGO2;d:J###<.=/RK1]CAH0]DU:^f&[K5=,bORf8[YBgV_\)2C4KXCL<:E+TQK2
aIDCNY.AeNg9D>8Y8JM62XY(R(F74L#Z58^E^T+CcG/R)4[dF#&XBaVcU5B^.7RA
#I(?I;/J?b:HY/7\U)FgU\ILL#7RTWcUP#4=894[+=[U)^PMT_#CVF@]CdY+bLL7
7OFN,(1HWRZWH;X1HG..H=+E)>+Y<CUKLDIWg<9ceY13cJ[)IM7f_FIY4-T-?-0U
//)/>[[KP/fS1,a\4fD0;&1<7_<7.AgTLaP3;I[IXP/X?(EGE+;bR2c2;Q;4,5ge
_Z=/c[6E;\MMXc?T3[;I9b]eeIJWed)LI4VaRY?&^>G))E5dG?,.6C_ZNgF\bDO4
@b79C5CZ:B&eO[OgTAa]bX+;YQbGDdYSUIAAD/HE9fS5S([Z)BGDMB0[?(-Yc)DN
:cT?0=S/FHD1WLRT1LZVI8da@(XE&,/G.:</,f#;I/)4KOU9;\>\PL<HW/2SH)R6
]RgGP@0EDYZSFfaLNAbI2>^+/[^R9P4SJg[S&@M3?3OOdb=-g,]B-U]GZZ[;WYSG
PLXBZ<JIba^F8-L8N-@2Wd)&5a2,K6&DV7GUL/GdR9^#R[IU7cI8&T1S>EC/U@U5
KJS9YMA\?Z_WDW9fY3SE>C9fLbI3DHWSXMHM.KI84B/PAEK^@H3c&L_Y,-1O0dgM
1#?:eEd_>=/-.0@Rg\^gOK6FBK>2[Y/ZfFI)L8YXfHa8_GBT-9R;d+d7XV=&cg^C
E/)0:+K16cVb.X5X^aYe[(NcTg7FHe_T>)V87Te[6eIM4^/@E>,46SN02=2?eKdI
N_(MPODPY+I@,>,YD;C2@+>FFB@:+CQHeRc;3)L>]QP5V5@Gb=G(4\E9KZ0^?R&P
777,+(Mg-_AN>/]LH)<N[CZ0K]BdAW:=aK1EP]^\2BcI>BLLdCXOIM1cE/:ZdbXY
O@;]VN1_N=0A,:01_\?(4NNV3KF#+a#G,)/-UBaJC?_U+.P4W69E+HcLM,DSWKJ^
5^]eUK7X^P=G+^_-WNPcP@bO3cN)BFU]#;cf;1>:#gM9bfQ[&?X[FKHX<EFZ_(S/
aE\9_&bXNUWcD0ga^R<&8cMBNHZ/DZ[c=:@(7>b>0\c.16X&UTODcOCe[]FV@./;
)WXE;6K:>)>U/<b=+35(8fb3)UJVH8YBVAcD6842>;;B?L)\@6A?Zd\JfYPVP=G^
7J8Y.?^R\O;@#V77>L+F]&Ub^L3\1G1MB4K?gR_1?;AN)BU0f&K#F<>b[<6Z9?FQ
Y&fB+7UI<KJZT9M=V_>cGYc1^D@07.604SJ=B\c2KE2EG_IC8X2<_FLF+bf&QN>I
B3D,aEaL]Y^T)EBdKaN<//<\TVUAQ,?T1b;V^Ua=&V/E<B<Ee;04T#/=Be]B9OIb
Te8Jd_2><2W52@P1P-eee4E/,A;AS@F9Q2@J^IKQ2W^E557>X<gG19V?B;bE(eI\
E)?<R[X0de6RGD_Oa;29B@B@PQ(OL^=+8LJ^B8WK--X6\GO1?;gDFUE3^YVF-I5>
2<W+>>ESQcK^A\KEe+LFDSfB?:1KRZY;PVI0PK_:WDF>IfK-E-):W?5P1(0:5RW6
=VdINbPCDcdT2V;>?XE42-.V-AFJJcYBJA?IbfVGBMD&@D,CYRJ-4>e5fFC#EB-2
S[g^PHIMN4IeX9:<S[7KBQ,W&Q.(3K+Xb/#K(/0d@DL(,<#b@F4d<4b7fIHAAQ30
@f,Lgc#^X4Z5([MQ:>QTFS&B^1c-G+-_Y94?N\/NaW?Z#]ELg&^8.&U^@NI\#11e
AN73M4c_X1G0/b0PQCA=;83I5IGbAfFOC?59MVXC.S=DX#>&.LLKTP?G:G>]>W4D
P(:7679QeO0R_3;Zb6CT^9LU7OGY>E8ULBcY2B>6(F>-E/5^]G3bMb)8T4A45SNN
2BXSFb1:5P\e5-Mg>+@,dVQWX]I8L&A1&&<-8^b&2[@+.4Z1HYDG?@Z;MC4X/Wa.
N(KKOb)3IZ#D4W/#E7d0g9BE;Q4(HfR#^EJ#D=@gOId?BT-6((5Z1e7CUN>U^=-f
a6YV8_a#JbZ&KffSP^C\UZE1VG5g0O/5JWb(L]ZFPAA.&Xc2VPdRbEXG56>3AKIE
-]HD1]>gf2F1S5#+7eCL+]][;U3Z7fbab\K[HUXdP&8RA#YeR]fbIQ&9fKAe#9/^
>,JCYML<=g^Z-gN<\;M-^>SV?fENB9EJK\e&4)U5#)7\^WGQfH0^d8ZVW+S^:?f(
H3182E66U]1e_@G,R-7R/HH7-E5MK(;V+JS\H#>8>/F-WUc/Ia8Xf]e.fJC2LE,7
_:R5dHK9dc<aE)R82=<.O7-QRGRM,c0@_D86?gMWHJ]_RGA7bDb4=066>LM<Q;:J
bUQ-2H6F_5\A>KRaYMETCgfX@K9ZJF7g+QHVaZ6#b2E:b^;N)8Z5KPIN7.?QGP[D
#cf16ZZK[g2bN]b7Z[PM7\+6^UYOMYP[gX@b_8Pf@9/E9S,NUUbfGJQW,D^?74PP
Gg5P]0adD4[gH?a+IR)+_gM53JJ&4eaOK6.(c9+?H76>[Q[.:5182Vdf(89<J7#.
+;>55eE,aTK:?[>FX+?I3IM2C,;@]2LZ=G7F<-ZeC#&92^b+e6EJ[7\9.DKR)Q)L
/J@>H]Z7[01M8[g-1(9/gLS7d)-HLR;N;<?OSPV.=EUeS]GB@L>3-M^b.f=B2:d+
^U<A>SM#>GdNf4TZ^I0Q.#0WSXecV2<aXcFZK<4T3MU0GW\1_Y.V1LN3@X)L]BOX
1d,<g\,NGDDO07g+L;\()/]Z2LLL,0WN.[W<F\GYDIEU<@C_f&?>O]>8-4I1Sd,;
[#Y<<L2a6.?[YC9>?[;3Fc27>LKU/WT6-.DeLA1[LH4V5S[\V+C:)F8eH#B>QgXY
=e.bce7D3[I;U\M]N_>#7PK7(-<S#4ZcA18,^;O@,L.VV_G_\I-JA4\1:eNN,BGH
aG.dT3<=4/>7(YP6\2IJ#2+;@O2AL-4R_e9-#P(Rg8c3cDB,Xc0N7fgPIJWNfP6O
_QK#X46SJ@7_Z__[.4d7e[5fC1?[1]TE),5L?9CTf#f(SNG+HU<3NNK7TWAT<cCL
UF@F\:2?EP/JA@8E74?89_^g?7eZAD.cN5YVV.R=R[@].UcP9TSYL5HJF>c;V\,Y
]UYCQ&Z>[e/8SQ4GC_GH/P53g,#ERf=X8cE^U?6.5[A+A-^9?-BY=PBCS:+8\&BR
@eA+1HQ:;_#1Q\[H=NKVabZHB;eZ^Y4\@fXdLUMgE=NW3JXaa2=UB6I<9?.[G#Rf
[S5AJG3aIgfD,.IH/CF^>JB.bda-J#e+OJ(/0^MMV2]e+H#+(C6)YKg0^H@51@T=
635MMddQg7_V\YKacfA:,+gC9]<1+[\,MCaE\954LZgC7E\dK0ZL(c?.Q+@N)N7V
^:01(4AcLSNbTIZTY&B2W8A>2M&IICD7c2.J]N.5:OM(6A)1)>4A]_\2P2eA44S&
U2=+7]/\IPLR?3JfGTQ(B)^YNa,aH_aV.JJDaB=Cd+^F>JILL.?-?UU;dU-:<6/&
,DB@>+ITgJ=c>2,]??I8OC[_]1&^.@DR?,U020)ALf:9WK7[ME#JTQ1LX9^/M_IK
L,8F4^.VAC:[I#XbABVH=gPR6^UP?Vg:fQTbg=A@0==EA6D\_H_9<#])][d_&e_2
K8[K7XWDTJc2?f#:2:>e)bJK:Wf&V&d;_HMNW7>,H@d78VAeeC:3X>AfJY?F.aUK
Ra4)a562;C8/+f[Lg]<;W+R.?#V;7PP1e5PD^aMR-BVN&+EM]KIQe-9NgK2d_W^C
KU82V:JG(RP:V]c(9Zc[<H^R,Ndg]Le1,Mc0aJ:A>T9+V+b3[23D[e37.G(OAU,C
dKG(PB:a91MZ0?K/E#S.JXWJdb_BJKJV5LXZ9^@a.7?cce>4Zd#W\;:42CVG_cZ3
P[H<d]^/g(_(0Z67]3L>a76^@]a[>B0,f0]<BQJb36EQE20U@<=Na&CSbZYVY\cg
c,,I^RO/XP+Z0bV2W<_?#K:eK5;&fC1A^.((58&DY(;Z.<^OQ./#Me+\+](,IA:X
gQg0eD;(9^RT9<ef7=BE0C(VJ7GL<P\E7M3F[]Xb[UVU&)/C&J;:(8-<.)aDf5LM
9O?[#[CB:?/B)(T+GUNEZ7PME4J4IABJg[Dc/Ya#Ea@:GPa(Z-CWfM&ePJCdBH5b
Jf;deeWY,FZ)-eF5dG2XO:9WGSTC2H7MJ/;(A_/;&S[/eP5)gLScI&.dLVX>P6@9
1+a^;/X>\DdH,3Be+MHeHIQ-EMH#ZE2UQHXN0J..7L^BaJAXe/75f)4ZE&PA(HJE
g.]cTO50#/\J^AP=?4JUNfDB0FR/f.<D@N-\PP&;eR]O8GA37?\73J_b/NYVaX:F
AdD1Z>W#)2W:-7Q8;T_\Q_=O/4OC=?b]fL/Y\R/RN2W27C:YGd78\/F86LZOH9-+
:I:Qc_[V/Md4_-?_NJTR&F8(=7]]D3EcS<TGZG\d3MaP87aB-a#6d+?>UD5KB:Z(
#=EUUg3P0/_HR-2(a\)9;DPK_2[XK>c0EfJ,(V^KMW9.WXcU?K7>O<YK]:G[(&_C
=I^,:ZPK[#,;:@.H/b-J^_>aV2VB<>.M_<&J&?LW.<LPVNTK?1Ee5,&F)R8H[006
XU8EP;T-N0:LJDBAVeR)JZ;A62J(]\LX^O&E:A,_+2OO42,&b34VBTd/=SB2bDK2
TX2[2TcYbH;6U&.YecKPSAgA1gJfeO_QF@>TNPK=GE:\@&K:;\=cX=E8f2H)AQ?K
Ug9=da1=AJ)PEccFY&#^HH[OVQ2b:g]CQ2+:LcF_.03dGW@Yb[(d+#70\d11+@6A
M0.J4GccI6fW6P#cM;WHB)_c/Hc7[@X,aC(c04Q4dBd[7\0H+SA\ZaSPTe#G]]1W
60Od1gX8B@fMJ[dTA,6QTg.<>[a(-D[g@UD_I)DKO,2L;5#GQGU?TUL>DJ9;2(ZZ
WO>9BY#T4_D&e\I)>ULIX^5(\V2bf?UO>QB4MR&_#.[Sf?WOcd3R;KbT2OJ5/G:\
3W#FZ9>W&-J8_J4S\X:J8;#:LLWN)fNO#5D&NgV1C05[E</XS=V@4W/?AaI?b1WJ
\X1=ZP\Q9S29,AD<07>T@7G7[4@\OBWXNXA+g-Yg&a\M)J4-DZWC54M,?NHY\/6,
(JC=^)QP&_Y7F0]B#)7VB]09&7ec#Y2=0NE<+&?AMf6eG<8>g<65T0<]TaX_P(H^
7RSX;,?7SZBg&_/OMWTES7c#R?(E(JQ\b8R_R_\-R47W:D-NN.,OHf=V++FREQ&M
JQD^B1>1f0&d\Bg9>ZM\A_S#O<X[bfbY459^A8S82P@B?cQbC-SJYLY3#b^+Z<JN
f:I5I3]AFgTMD;ITIB-FH)SX@=.g0DE?eDZ(,CU_.3gUQb7]);=eb^V](_HPf&G)
]d<0X9-IAHYA9g4Z_[c8NL)7fJ2I2W[V4G&_dD1c7;9M)B.)V^BM4YO(S1dZeMU8
I)+^=/Z9Q4V42+=KZ7b:MV&U8XFSX6Pfg,B[?)VLUAbNKJV232]1[d^0(W71V8>;
[3dUg8:)3FAKIZY9D)N2Q<@Z&N+\KJQYbM9fLB,WQeGaMb+T,R>]XJ5H5\R4O22P
ASC2GFD(4VLE2L[EI<NUS.+fJ;>KT;WTf-6f3)8)P0P]=UX=//,T,C0MZ9Z&Kc2Q
<4^_[YP\V<:_)cQKRFeAK1Y?I:[FNEFcBC_->J/50PY8XE9FC&7<LZ7Da&Hf3U=9
O0L.+#)CUL6.\Y?_L:fL.ECEgP&XY#1?-)We1GdSFTe>8<(MB5ROP2\AEVbNFN=<
Dd+GD]4&2=JDCO85/Pd7Ya]#1[^c\\VQ8T[H-SZL&99?E&-7a]2(AMH,9#[7OX10
)I4YXZA^\5&CU&-:g4OUEUC7POSb?(Xa6)8NLA#Y_1(HZ:a#5@0EOPZIP0O5LGQ]
,ORUSY?eUYfa&J+_>bI;[GQ==3I@g51,5^0;W;([9<fE^M06S=5(4;IK9H1;4UMV
ZIY6YQ6[e9K^]aE37-VH)DT\RJDf6WPQ6BLYaAJaCEOE.EFR-LHAYdG<(]_NYZG#
ZJE4;A#+3+G5R4,M8=5fEK07QU>URF,GFHWJG,=AS_@aKAa.H\@5OQ))^@^K<>J#
Q^ET6D5\MSdSRCS,IbIVS2(cAR&(IHe,)1M-Fg\g;VIB<7<>=;.+2Z+FR,V2>-Af
R(1QeDXOD7c95S;f,7^.edM5X5GESL6CF7UL?EF2e\:f2](GQ^Z2#H&[I<(T<Y.<
2EYeAG6K)+,#Kf8<]KO;U.:ZOQVX?7&;SMcbfO/VUG1^cOI;H=_?_bUY].Z/L?>.
/(:KfN-&\7CY(A[+L;[W&\8Q6&YUDc8gFV=_(G)?0Cf(d[0I9]YD79)79IVX/;_e
SBIfS18O.N#]CTe=U/I9<^VHgX;,d^0QAP]e?#4W38<BB((P@S4OfIe(HdK+NJL/
9H9Rg@9[^_Cf(:S_\2JMYc[/[Le##P>70aG;?3X/02g\d(^C2baP\J-7U-NMM]:/
JbPQ#,O9HEH3F^cIEGPfCA[SI?K,8@IUW[-)NSAJT;\g9<F4@=N#TBbY;0(?]cBV
J83,L022^&:4HPR-L4-20O,/7Y9^H0F</#-e+IA^L-gRd5?Wd+IS0U5I&U1O0\0)
?7?=#.MP3KgT:_M=Q(YRa9-K4WFA=I-GPAa\X)a#T^/:WF=18\-D1e]K.#&\ION1
NJ:J))FaO6dXV6VQ\48<dKRd-Y#K=MaX5VJfW4IIgVg/X^TTCZC;.K]2I\=6:D10
38,a#IUU,#K(^U6QEO5_dA6;_@g&;29I\aD14]aOMPI&2W#YSNAH^.:ZZ=4TDgT1
EE.R>OI@?Iab2#3&]?0PK8PKa=(O58BMHP-Z?T.N.PNEOCAUa=+GZ32ONNB@8SfS
Tb6=QJ2VMEEYA@A/]bJJX9S.[)D<IBcSQ1aGIU(f>A/MDGM.+8D_A=bg70F?Z_f]
<7CCfSF7C[UT+0BE=P<XVUW_BW9>D)20Z^H7eg-,=Q\9X2IbcF:VZBE9^.2B&).:
9PR)8B)(_QZgdY/+<X8XYZ4QL>7.\?34>Xb&Pf>MbVb,4cUWc-aU@1,Ue0+:P552
6O>b\:b9_?RWHH,QQ?3N,F(E6R9f7Qc=3/?4+]S(UA]A@,]Z7E90)ZF\[=@d>:g,
[cGDb11FIGUcTB#aC=<^-:GU,S+HDC+F]Z8/-72=<L?-9dITYQ)4N+J-<=EN)O3_
(-de67;>f.EW>b-W<f8W_]LbQf#21M/S?P[XM:e(&^;:8?)08DOR@=M\T&b>6)1<
#V+If-4MF8CMB.W?G1+BQ927)JYN?KOV,Z-A#:@a][((K5-3PM1_;aL<P^@bgG3-
D_>8M#P7]@/Ic5TN@cOWW[9PeKQ?J1HOME47Wb&aS+#RRQZ?73d.4W#_WE1:dfV(
\Jg#VWJD.1Q,+>:Pa1O/&_;XcE4Z>9,g8=&F4AW?Pf2E+F^=Dc\dUI4A]F(586T&
EI#B73DH<aLe1@FC_Zf@FDe;MM1TQQ#.9<4c<eDAZ,17,872_>f711L7,J+PHGaE
EBd4_9WL]AYG./];6fKcMV4OJ_d_ZYJTNF]Jd=4K+/_HCSbaOFPA/LQd[^gFVY=g
BdEagK>Y0>SB;K-\O9^]3<_QY.&7W63\JAId+MY>,A>@<#_DI#QfWC;318DI8^Y8
+T+;fCH-OF(;4,fXWVb3=EP[f5LN-M>667+NBFU9>eL#34-H??KOE8LHR3Ve>deT
2HRX#1(TgSN?Vc=C6H\c?9F;g(GBc:Rcg\3[<?SOXSQc&Ced[YL?ZJ^)Od-UPD)4
?Tf\\H;KFP7@@YMF6d:WFO7N8F[(93U[[#V:N<1QY\=e2CCIM<<B?Q17/ZNg9\RO
Y9(+.EeT[M3#)&C,NgRR,b8WRCV>Kc1D)NI_PQTJeF^<bX]3.ZV^WC:<9]bU\I3+
KHe)5]W5].=ML4(EF4ESfg+5PJ=T3JK1?^RJ.TcXQTSe5N?30<7LCOVbaBQIGOaW
Db1\47N;A>dYA2:7T#.,^.NJN#2]fM9LRKfOC3GKSD[9AUH9TSce;a-X-SXBJ8@T
9aXQeFBY/0)W0ZD@)Z:/Qc[bI(O9cB,GMH4DY4NK>aC82<6K]E5FXJP<\6e6YHUc
S+[deHG6.NS/b(],QV<@]9&ZN7]0G[U)LJ<9?HW=#0LG03RNA]UP[?/C&ba&;TC@
8=;RD>+.\aCbX<>S=09SQ)M3>2D?0PcQIW-e//d(7Y>692+11&^#ed,(cABU_0#X
EHgBXM5P6_H<L\?O5d;-;./,gB_-@R8Oa=7bW71^]+I+cQ+I86JK\gEQDD(aN1(e
NZ3>c>18?TZPRE3?d67Pa+)U(T&\b5?<M55fNA,=+)Y4,RO\XK?7GQ/gE2UDXg[-
#OX/BYW/b9b/GAe:0MXaDL&Udb,)4]^<bE/M&Q([,fUeL<Z]>#6M5-gRbT5?CR5g
FaWW0LXg9[3]?YN?@N_M#C9M=5N];68LS^5P846VM<.ZHfUbg?^DX,L>RW]I?2H=
<dd8EGV_aC_KQ#/9,]Tf>Y[GeNP_bGb[+gBYT7P<8P[SD;f]XB@Z)2#17KM6=32H
:-4eA+=Ia24P+HR\/>bTL0\f[QWB\_1TBX6BB4K,BY20RSWf?ZU1?gP]d>^SHP]\
1XB3LO(^HJ7b/V7?FEP]^P94Sc0XF-RLF[Ng1P]FLA5<T?eZJBZTXV5]DJ#-a+O&
?]K2S<KS=H<64.CQV&+D)G1?CD_7\TRBTKU,(f-E85;MbX6H(A.L4@AdJaQBWWR\
b]ME>FZUW\YGD3d,U0Ragb.0O9H@4e-TD6GNI-K3CHAY7aK-O6AUd^]P>[0_6;.O
[L3_P;@^[-=<HW#RX4aN8+=X<P?-\F])(,/d0gA(&eG.R_J_;&,XYb_@GXV6\WT.
Z,/T35NM-c]aRcQ(<JU;A_J/F#.4P85gafAR;<?]g5bDAeG3U@A@:Kc7#I0??:-<
dGQS,cTAb\49O2-IJOU6W=C06e<9U&\O37_K6L9C;DKXY0M@,_IKZP1XQb@)1V-R
LK]G(8S:B)Z\#13E9Y86-SCR)TYNWT:V1?7,2VMX70Cd<1DYVV.C&ZR]F1&K924@
I_J9Y6LUXJU4.aO=+=<(Q7<\UWH#F3U4OAAW,8@Y[bZI7da(\T)<7]^78P5RL#@V
H#HUV^9^DCAZ2ON7QVebc09H8O/)TET)G>R6HDW;K+f-^1,_W6BeG7Vg[5TA[\+-
C>S\5PX=aQGZ9U/6LfG<Y8gHYc\PX.@J7,Mb^HTaN_5I]bZXN3[&]Y=Wa5&]9&e_
1>\KNf4C9IZNA+?K6BS.PCg=TcUK.AWK?8#WNX1T<d/GX&TR=L0@Q)b\M/\>WFd8
I=cJM?=fAe;KX?8CbG1G0X]O@X?R+eX59aI7;IV:N&]FFI\YIcZC6?0,+T0\cFPM
759Q5SNeIf=\6g@M>(ZMeH.,aHIR?#.g@3B?d]\c<S6BZaK42;[gXX2(5H,IG08G
]F?Dc0Z./^CgFG8_GS1TX+FCYgJQW-3d4/;.f(W@6SO&^OMgNc4@928>OSZHN&#=
X=J8eM#@a)XK+5R\3DK<LU?a&XS;GcTYB+BSP4]RN;TfX<ea_\gbJ+CIYR@^Hc7/
Y>OdCI5OV6eQWV4XM]-GKUVR/A[^:XZ[B[G47ZM,XPSU236b;R1VOF\DC/,&9HSD
bV9.8)g(1[Be],C,\;[e=>T3,XU6e?YJE=\VD^_,0fHDIabG)?=<GYX=2:ZY;6]&
bBSLI[PNI45E?F0g@U]R#FZ]4X-/<CRg>U-W14Q;TH2K_TXbAFP95,7OJ_(NS/3V
]&-R=d?TK81dB([N/<1K_0L7-]c(BWc4N)J6Uc3I8gB,bNW#T6[ba_ZZ#07d^MJD
78G.)cN<Xf)-#HS/SB:.KK>S-6GNACZ2FEM(>a5O#d\UcN2[8b>,BW\T;Tg&I&d0
]A0(7XE?[H&Xg]dba<UU[#OOBZ)A^)bf:P?R1I(Y@<_ZZ<V(;XAO9V=g,:@F6&N\
Ua2Y6<QK]X#+9[@IE7D^J2daTGDWE8fA19RPD99f+36>7d5K2ZGKDL<b@DR-d&gM
H5SG8MV]3<g<^8X(UO],HRTcA7&BW4\f0.C4K6ZN+3>a832c&:e(D;F6KL;KSXIQ
WPHI;T(TI=:\MOJC]:@X2(RO0R?YSV7Z>XgNHBd>)+0>/SL-9J?DD20(>FN6G93>
?;<K7[B_]=A=b)dP\P2cGY_KZUdV]K;&A;0A)6/U3CC[+Z?SA7.]H+MXQU6WC.,N
[.CEF/FBX2?#CTOaW+fMNM:<Wd[LOM)PL/(Ec+5-@JBbZ6.N8PM@)?b7b<cX)?Ra
;(70[=\e62<(4aBKB(TNdAQ2VG(9V2V?1Wg__gZU@XA]P84aNNL)cR^\G#[dJ)7B
<@R?8F[:5eB-8O]V&LIJHE,N?YD7@052R&<EUSRdTRVUa6aBB[Bf(-11W.6R)/N.
8J68L37eH-Y^dPZM;CBSWZ9(GO/57JKQTL<a:b&T6A0I_;XV-6]=53OG]P975_>5
T)6TB@QKQU,c/8)_DbX&dPQG]R&8TdD(5g_1N6^ZAFg5E_YB[Z=,->XB<0[d[^c-
fc##A4<Lfe.AO&U0]OTO@V)[f/dcf#=#eLOP])W[>#N[c#+FL>/Ec[Ga)+d-OPA6
HPS,QJ@79\EHZU=(6;P)N\e<>/@Wc6eX3O2J;P0V6.@e+GP#R_6,.EOUD2O+TXI\
TN5,cDIIT1Ja=YM\O-ANS6B#98d1;-E0QT0,4#3()TD4;gYFGF(]7,@EGeUOcY=C
&=)W_JIST[3QRXPVO@gIPMC=U^1/ZPHH]EK,99^BA/7R6&dSA\+Z)A_R9:HT8aaS
4Qb@&0XXBO3H==LfKTM3b^eOb.&?^BD+\c:#=(/X8fQXU#V??,W+@d.60HY^.RBf
5Q][-a2QL@&gJZ7F<QFfG1E)]<\YM3(B4Q,9O&8@4c?XY]:-bI@H6\&NC_@MKTH6
NRdBNJ,3.XCKO^3S,VY2+]cgUV8._+e.(J)0TK+,1IbZ1NJT_Fe0T@L5AB--G+5(
?T3bb5E]J54>05TJB?eM>227H>HSGF(IEUJ+c&NTDdKDJ0>a8Yf.WNDZM:<CA]<N
D;9-6H#,.=W#S,[3Y3D.0bOd5bL_>93HLS>8._4P.[8/@MF3YW+gEG#6^)ZJI1&C
dV0B>dDK5eKQB/D(+@H>A6+UbNf>\Tg(TXKCEggg39gAQ>AJWc?48PW)DJD5D\=#
0V.NE5@,EceC+_\;GY\IQb#dQZ:#YcW/.&:ZcBF93SHSJ&d>;/6Y1&RO@Ha+@:_[
I&V#UJfcFN=G(V-LZ5SYNC92L(_BbH?;+OW@>P/Cge,5R.=O5_bM>L\P-BMNBY?P
+UMa7Ef,>P8ceX>Zd3WQJE?YN=WB]G3bUAV_O:XY]\BH++F:BA-1YBfY5QeBNSAb
@7Wb,]Ecc6#Y4Ka[==(Ke+52.DcU^H-e>JRKIaG#.I#<7@ZP2HR?WCPcQD&DJcY.
J>00H\K#N&1G9?0]GgWHCR,dW<?-@;AcD=]\a1J:fZb=C:]_e@7+16M-/AQ^&VPD
d(DgdS0BMFM:B4eSRe,K-Tf@F,T1G&_=T9)HQ9A:gE0dV39XARR:FV6N70Pb.P+e
CMa?><Jd[gGC;Db3?)24>Id6U1[129?4VVU4aC1U6QNYDYYgIcNY6/.M55e?Ab>K
b_@_=UfY6?NCI3.((JG62M=8.2DUB5=?(CHO<?:\AXZ=>RWGZ567b8]2@Y89bWd.
MOT^E#WY6KQ#[I_56+Bd>->BM45D()\,2FgQH^>5@.eFE^(E(gSK/5X9USS^1(ZS
Yc3]fG7Q:GCPKNH38aF^5;8-QP;5/->V#J]UZ?+V.H#ZbE7aHf2O7[TJT/?eR;d]
^;0_9RV3\85.f=MT-8KHQ[ADS-R;[>cCgMK0&2G-1[0^.M=XO4_&4^#b&=>+XCD3
;P4.X4K;e;3DKF=[HbB+A5Q,M;CNf0&EQ6H?]Ba10+5NMUBRA#aWUeHJ8_F#MA&A
TZ4ATMI)NQ?7f7;9&O;FWG[\?,JR2[<_&-ddJg@eCJ(3]=5&eTae>EHd@LF1V:;>
fI<8gW.PWWXLY:]1Q=4f5ASRF3QB&3,,8IQegSOWG7:YGH[BPSV]57g+cf:CfOQT
4O:gKd4FK&DIJ5HBN(aQ7OFD0gYIT-:7UMF/dBEK.bUb+DW6EBb25&X@O4+#ef9_
6[R(Y3(2GXQgAP(9K-a>^<Xc+DTdW)+f_-,8bF\b?fePG&\[0<8=@L[5eLc3RFb@
6c8fQ:d)<-d]B-=9:EV-M(4KR8(5YD-,f-<DT>AHVM3QP/8N8Q4_&6/4=Y#\fVT3
.&<Q0L?3VJ-D_KW[L)[868GGJX:W_g:VgMJU[Te&U;fR==AC:+Q0dTVI7..c-d3[
KVY3J3d;JU>#F+_LPQWD,)4:Nc/IK1KY.E+50#T8KO+]dG)2F2;@@UNdHV@YBICP
RTZM/X30.b@7X,&JaZ=W&&V3U_aR<R#0\4g1\+/,0+H.&<N?O&b[M>TYbbY;VVD2
^dGP(F9BII;Y8EGW.K8OR[MNEJ.[A5Q@fFgf&c#^aZ\NgJH3eD0;000Pfc#/-)U&
F<V8^/I#?CJa?S@N7fBR^K&6JV46H&FZ2P^>E5D5Z@=N7&I-\B<@5&>Z7]P+W?[#
_g9A.\^0+^(XTHBV]NEQBDM<Y2];N2Z]7+eI8@[YeTPQD/AdMO>+b#0/eY)f@:bW
]3DKc&DKaM+)XV+L\,0P=d]_Z6D\DARE][McYG)[eIZdBG1(g:5c]@SG=CSSaM+,
2bOE8f@+c1a4IZ7A/9IMNN,c7Ab^0.Sg)YUWOB8aDRBDIVBDCaZC:IWKDNIFT?8W
J=9UUV,)FZWWB&XB?2WZQ>8)GM]S@;&99=/]3KbHAYMg3B]E3+2ZMJ;]\]aK>&1C
2P&0NEOGDD<F4Hfc-U?IdCUQVBccU&D&RC#;[f<JdG[cAA-J7]G<AGg32<\.,gd5
^c8>@0=_gGCIS-M<&1+3R&=ZV>>ODF5[R)[<gEC&[,a[P(R6JS30gaGXFGMO.ZI.
5:Z@fF-@(RU(#W(>9@bPG]OSA3(F#)>&QH/H>#RJFO/ZgK4+C;fG>Y5&;=[3=,8Y
4:HVAQI>Q88d7bOQF0#5)+SRNc=U_V-N7L(dQPBQ\aVB,8@JPVaSJA9M&a^H=,9&
Y.QH]D<D;5I360EW5Tf&ET]_,5.)0FBU7Bb_dN,@LU73O<e@,MA,OEEZddSE<534
&00X>+P)QcVPbPd7>Q02f+9CF+e<984SJ/J2I:+aC?D_^JVbXZ#/cg^-@GBZ5b<d
J.75XTeBa-SQPP0;T(L<KML,N.fG@a/C>LT<8@B?Z[9JLe2QS0eH:8LT:Y92>VLd
Bb_M8^&KJD6HbNf@,4[@YNRgH.MKc/.AL3UKDM_IfXbO:C;e[Eg?b8+d+A:XDcG5
K?bWXPY;c[Y)Bf\T>^=bWLc_Q:>c5WT83O2bAJK&2T88ZF4>HP.dAT9]IfZ7fIc1
\gX?7&c87<(&C>MKfZ=63&M\7a=b[bF@0/UQ.eFT#(/R,BUF+f:-)ISDHG#FEF.a
>Kc#@<=VN4)./;[S/5&/Ic:L-T[TX>cUW/((:K;+@3^PB2^W[^HNVT,b.cSJ?P(^
)gbK8._bRBbB&KP/D9[,d?\&XL4:E54=6W;6-IEI9)/Z-HQ8#Lf5))YANKHd0WSZ
;]bJZORFWH.WAAOGUO\CTF0T4KZ5_<Z9.U6#<g2XcYXW-LC6_5[@<T\=+Z,8BVF@
O6E6g]@\_3T;BdO:JHb;@^\_QB,1bSVc^@(NN/PX+B(./J6ae0G]?C#3<U5?Q-6Z
RZQTI4_28#GEBYS&I?SbRLQ9X)J]->eZT5+,WWcc)CQ@B=aZKb1[_+DN-2?12HJd
3ADHE4K>E&\,\NI_5X;,=9K\[.ELA@F:PIb=(7aFO75(QWc1K4+#66H.59JR)6a8
Bbb<A<BIB9c@b?.HM8]TEX)1=@7N#QF]]N\<ILRMaF0P,+CHTB1RV_?/+<0<aM)P
H/5^)\HMR;;Fe.98.@5^#c9)eLA9H(C)6-VU8:.=.eV\>&UA@F7O8DIWZP4?GDT#
T<6-6^B?/TU1C0&OU(M]bR:-7/;<c6:.);MP(Y?7cG>EHY#0K;VELS@:?-B_LECa
;QC.RJfT0X#;3,51(d<BX?BO6W0@_/_&8=UOfMf^(8Oe5]@XF=OgV_Se^b<:[REW
=e\dI86D3L(fd],Y(WFU3W#0cJUH_b(1EIE[ZJWR=^^geeVR&D4&_PRX80_,a:bb
4X53P[N/c;R><e[EK:4&\Kg,U<dL7Y31\dNe<0+,DYM1MIf[4>:K5(7[U+=e-_KF
H>dQI_+FG:.QZZ&01X;@N>)#&;9M4,aBc\ED/R9.EI>Ya.&<R]IaHJg=+EB)a_#=
1J?B<cVG@;MGX7#<6c2]0R?KSdCJK(1>P#H7D/MRfZ-RMXE7@/ST,>57J5YNS=G0
\XJ-TcHTcJa?,+DJJ1ag4;2Bc(T.C[:,PH[f?XG@(3bY[:dGJF4R?]E9;JD\[Wac
NS</_\/8d+YcdYgR4[(B2L+20<Ze1=2(QK1eXF9R2@8QV0&.9G17,HVdY(NJ:g]2
BP&E+E(=KF>.QM.C1#V_Z#fe=9?M>GXSgTG8.^=.6FWN-0F^#UScW0BUCV7AMRJ.
CZY9T\UF=IaU3A;K_d0B>Ab[N9K<1@-Y=dD<Sb0S2,[E6V@.JP@@CCCD]L3Y(Y7N
Ad1UgCL[TUTf:0F+c=<C=PNC&G2O(M_+WWZ/S2G7WS@:F>-NS645:Q+7ET6^<D0P
:(IfJb6T:@Ed.e7HSK;>O1cHSfR\aB290&WO[7BMKFCM)I5]Z/A-R@,E>&_L1RQM
P<1BOAUVg?D7?NKV&<_2gP9F]cVX&M?IUaL3\3J6-Y)b;I.VH:UX5ACH55L1/Ig)
f;,ZWBdACRKG:/[@#+O9M7&H:Z570@0?N=PX9=(?M6>I7O+14?=,EZ2-)M]F>#aL
Z]KTJI>1&P94](d<5##3ag63:GVOCg]E4@9M,N#]a+OM<b,e_\17TQa^?;;-f58V
#4;R328(.[CU,^A,JFFC_]9GSGO+/3D5B5R6ZQdC;]=2.d3&E_VAB>.<VU7+PH;A
<^EBLA0>0-ZWOU1<ecPc<LJL58)?Be@N\DgR75&4D:8X850H1S.8fU>5DL&X)dFa
GSeF\P59)I=N.-K@e9VT?C,QR_b/ENIHMb.2BZGdX69NA,AHYe#XUgF<60WZB.QP
3e#>OKA5_J,T>1a@9J:K4#@S-7393GRWT@B+]Vdg4-<4GIbPcR<D>/^-gd^f?0N?
]W-Y5RaCeK<Eb8KJ4g,/HNZ4;J:e)Y0Q3cUa:3>7OOMU,]M<(E@>=;B8AJRLH5>J
OI?A+UF,?UB:J3E3R4ed\KC]/f.]U1XcM[,JObg(<+2Zcb;cBQ#\ZbFED/F8?7f8
],C;L<;_Q#8,TGAc:WA1J>L^)RNAc:]1&I3Sa6C7I4F2BZ@]0B3G[@7ZHA0/C3B9
DQ;WYD-+TV]2J_YHM8ZK1ab&Kb;HB-FJbc)Q(?VHG@D#>M)V2A\.6<(3R7ILMM;?
C^Db\NB^,#,HL&.\_8IE7-51(IJE>6<5b]9S/e1c_,_=M<&^?,g#_/#fG(.W3==7
2cV=.d.C.@0RDKNb+PYg)8_@@AC2,NQI=YG0/1U,D:?BJePJ11R:ADO3FK/3P\M/
^#)UJC4c6<MY@V)bH#3HO+9g>IfN,4;BAQB_/eHMAJ1dZ:M&JP1]<J@EgVfMY::@
B7_Q84GQa,\:\)NcM8AD2PFMZ=9ad&C6YC&#6#C,QMW)NK3B3<cZ#]:MBC,:K<>Y
R0/#[dP1>YaLc9f8a(&1J<(KfI9:IIL?&=5XN_Y(J80b1bW\/f36K1FS^L^g:0E0
Q;F_=?.7,&C7cP^)4.<14.(g9,)AgN^SD2C82E84,b;P.;?]5[Q4AgA01R?a<VQ,
1=R0#&<&c[c.44Q9VWI<O/gcgK-Y[;L)d<PeE?/T0AdFCebM?6Z^+840_6,Hc06B
,^G8&>5885OMVe&_dNOA[XDA<LX-TX_NKWP#>97/TeGEe1[)a[BOICcLE#D2NX42
H1,-^B@8YY:g,=:=1&>bWYG_MZF@41f.@9,X76@16@ebE-))PJW,,+#bZc1(c44?
&;<.U2gS)MWF#]@/Z[+8]/1AF38E\]1-]95(VE>_Ab<EUa]Yf&O>b[Gf:4K-E<f3
C\6_7;^f4c@E+OYZAbMc^=N68CLLcFXBd:^Bd<H/&7dX80O:B_[.K)GC2A+()=RD
V6]^E@0>A5M5./.O2f1?:\NX[=4NbDZ9.([.6@T>+2f.dSb.0R5@YdA&Ce0MS6EE
+A:L8I;<]a(:_>Q,1>-(dK5Q\0,@76;R,4[U&L19)J@OV=)O=4?(f5@OA:baSW^I
]?B8X]ELH8A4^^P:EQGg3GFNIW.D@@g[;=VS)>U,b,CC/BZW0g_MJX&KJ\(2L5W@
]<KG<(4g-UP2NR7(-69Mg+W1#W=H2,D?(8b?EQb.EVP>WU/3FcK1[c[V8L8F=(E^
YYONJO-FQ#=HGX)]HX),\EK\6NO\&M\fcPf6P;O^\DK7GfX6E5L>-K#Ea^?6SaKg
ZL[#D#KEPCH5f&I8Y,EC/]/0\@564H?B))NPT@@V&T7KJ?E)=&ZCQC7^BD52SLeA
\FD1a:Dg-7PRA:2:8:H_)UZ1gPSU/,ZBB0JC+_b,#NQ5:E/YZW:f]&_>FNDGL/Jb
JRBS8P0F2NWR&6N/3^S.?,^2P-X9Y>[F+S)O7#7,W9=>d=c@RMW9D9W.47LSafa<
6A(gQ(cCMO74UHQa<;TR)GQc?O=A_WE+P7W,7N#/E2B)W]=OUcM1Q]Q;/>TDf;60
5\[,^@L07GF_\.U\]^-Kd)4C72]M+ZX&8RQaMRG,7ReR>P_]ZbaV#.?^EgIEJ\Fc
,K7=ZQZ\BgZ>0#A[Se>2L=OX6\>F)Fe=eWNcMK1(\PPa9S08ID+DC004X)&.BY+V
d#?e<RJ8AX?QTT93[1):KI\2UQ#^DH]?:B]a^gF-I1,]ZKfME7J(\ePRP[6I@5T1
1=B=+D3<gEPf4@VDUP]\U@IL2Q_75M82b^Ra5/7-?&_03,R&)Q>.G27VDMe.AV>A
X.NXJUB-/CLB<;Xf?)JD-6.b-CeJQK8f+cK2UG5dJeOYC&IdV&1^,Y/QcL+2g\#@
^Z+_PSaGR5cd1>J:31,J2;;HLc+Z#.VLN^</O#Z0O;53@73DS7B>@>T?VBEY)a<V
5IHfUXAQ3;\e]1c8=b642,.=)VR)C4]3?.NH5J:1d-#Jd/a8fcf.(8[eAS8HU1I9
C&]^7_2:F(V-?VEL+b..#b]Z>RCH267:G?#&NW6:AZN6-78e7Q@CcDK^90fL4\)&
0T]^1[+HeUN87.R>TcHd^PRc)14<g;CA5Z.Z]/6+B=@]D[9c#gY(3-5M2?.ZNbeZ
+3TRc.29,0[[5GKS4WJ/M0@d;+;Gd[Zc&&<:e+ZFCJ,RHN55>8Ebb5aNHdb#M66Q
f5U6)D8fbU^R:4Ue^_eAOW+#?JXISR9+F4d&^cO3b=)X;_a^LN)7dHGAUBFYXA]4
M7Ib]f[Je?(^KAB^>J\g>^]Y1OXANe(Jb5ARPX-1YU18[0cM5,(T+3-Y-;K7Be2^
H//bVOXGLgb#6I9ZF_8NG.GY))&@e_1A?JW3?P@QZd&F\#2??/_B#gJN@ADY]RE@
O[R[dGcOb]52@M@\O3)R^8W-V]1,JCB0CURUDX_ICT-]/)\<T\J3A?c_E2ZJ5Nc/
7.e7NIEE.,A;&,Db7MAX]Ge3f?#N:#PZc?W7HbcKQHC@AAQ5#S@S?1Z1HRDe=MGX
e-<[(0Y)1,KJN7_5#c0cNP<)5V1Y\NA;O&8O^W^7^4ge,EAdb?S4@&PQZ=@QO;8f
7aAT+<#<fZfOdZ&GL^c3LQ0A<]X2VPT5G.N=@/B;QECEG,3&>@8-15Hd@.IMea1e
1VYbQ55)b8]PYQ?cI\[(39SCTXEWOG_cJ01<gD@ZF),f\4N&3gO,<e33]+3_J5G@
.0(1\IC:AX@E-Zd&_1AMO\84LW&5FLLERGb:A.Tf+86ZRLAB1,:@,SC0H30)1_)X
aeC[/^6].eBZ@.A9II.QFPS#,58ed0#g&^H8=&,]KS(fR=&;#^G(E).^L^f.>Nba
G<#PHZ3YIST)<==2=HP<a_T/gEbf>Hbg1S^KL?I:Pa8RXTaM#,Q2)?c.M03fSF>e
Na_B4?a7833g\Lfd.ZBA#_=8F=_b;5\[02/fHJBb4Ie129/4FE;M(T@bb\J39^(3
ee:8V=<BVbGM)^aOX/@.(CLBZOC;R^O&aAUOCQ5(d9.1)aNTRgUcbBU<)AHAQS;L
M-2Y],D<MKINGCVOc(ebUfD+T+>B&AVG3VNgB=BFf./ST+ZK0L8PR[P?OY=N/Q1>
.Xc+CJfcAG.FVG/AG_/(JQb[#L^HN<g4]N3@4;S_)e/e3^^NeABB&RZG>Q[:[<dW
Ig=F)W#3ETWN(D;?#MA+JLR,L7?)/N)1[8Z\P>9d?_fPKCHLDS+G(WeeIH0Q2Q/Q
7[X1^6b:5&DV-A.ed3TgE9[g.+e-a.g=,GS2dY)^QC;Kc\/+YZ02NAQ4e?fcH34?
ET&[)+V^0<TI#&8)<FY]0^8AHMD+>H#R#?5dVW.]RQ5SJb;-+:#6HITSM:Y0SCI+
;aV48[gg-/,9IL](JFUc2bZ-U8McSc>0)/a<0<A=XPbO41/0GAGLbAdFP_J,aKWB
-06=BKfP8G0LJdT6g1K5ZOHZfX0,2Q9#G2LM58K0I]NDRJQd\TG^.I[RdUFZ7&;A
Ua?4D/8>&3Sd9;E,cBd9#+X+.1&bV&7<#2<[K);@Y6]1\#,K&a5\VLK;05MV<SHB
OcN2FO\#2Tbb>72?-VIK1ZAG8R)G[g.>&OQR05IA;G^RIEQfL/XK.[YD&IdQNW,Q
KbKbX@VBMUO4>70Bb+(#AQ<^e2KI\D5A+,0<,AW1gY\[M94SLHP/;5WY7)>/DM2/
EA6),a_XE7+-N4)D4c4G5S<E;Ad9:18;/Ff=94d(K6X>?Xeg5.Rd7a,:a:d;0?WE
0cg<NZ520?NQ,G0P(<LM\c-\?QeLDV=Hg9VTdQ.>U=PC_(0V#OETYO@Q15LFa8O\
@E+[8<D?4gWTf<K1->0O:(V35R5#(&CF\=?@.)eYA1#fAYe(LJ>ag&:^JBRRMf;W
TFLF_,E2.F.[aNaG[URJ0faa-N=]_\G]JeQ70^->TI]D3X(WH8+G&@S<;&,,/c?R
)fY@Ua2E@CKgcYD:cR9db^C;]EH3JI4#QUf5=>gER\Y\06#Me?W6M9<^f_M0]e>a
F9IFTg;4?.<cM06.Q&\EGYL)\@8R0b[;Z3\8D/A6;3a:GRGOYW5>UKWVU67J]SZ8
)^\7LRR=#=,LU=3N/e>X+14D;V+S0AKf.@NF.X^#44/(][W)EN6M?SX=^)N8(dBU
_UIJ5<#-2>Zf?).)W:/K]_4/P1?1f?M.bG96A).P09Lb-VGKWa.JS@2?B1MKVE&#
e?GT,A2(3@C@M:fU&E]7a:86UPc(-]W[8\cD]330#0S9TSa6JLRM?(M+01TEEcMd
Q.NKc)>C>R-^7PP8[?LG8E_Y;&HZ&fgZA2FdW<.E:C6=Vc2TIVS&JGb/2+9K;eMU
+CDaXYL_/>)?;0]U>O4P(?a=WOF.:C+T.+]&GT2?LQe;)f7Y]F+gP0/@I9[_/5/e
X+HX.B/0>/\XE#Rf_gKT^#EZAU)J1JENS^51.8-75-=A?5AB&)[<c5CQ#2d>H@76
;O<@-DCI/9bU\&DZ4^cd&B<)VEg;S27BMA3=ZMWNR8+I^JJGZALKXULSV,,^&7GF
VIcfB9AdO]ZV4(\Z3W4+DK4T8ARIX_,^,Z7(,2ZfN_&9)/bG[JGQSY14B-NXIW8B
B,F1=aIgd5HJUGMA4UFdR,7b4AV(f-\BJg5Y5\J#b2=WOUVXG/FTB0AL2T1.O38g
/gbF35_7L_Y_?,M><IXDb<1S+#C0_,+&:+;>O#-d=EVK)HdXK9^^>a_-_?O@RD/X
g+P86D+a<_PXb&eMU9ZSbORB)fLNeS12.M3CO1)P:/]cO0A,,fE_7gUO2V/gHgJ3
Z9f@MM.EF3+7bBR)MLg.gD<NNBGMVWKCGD0#d//FV_#BY6(L9F3>f0]@PY60MQ>V
Q+0B9_90g+1JRea\CE(b[DdM)PXfI^RdNe><[S?gWM+Hc6QR(]XfJ;(BWS8D.[gY
<6#OJ0X88L[f\4((P+(AcW00X,gV=b\aP8+;/IMbG[L.Q14KF@R:a\Kgb=L8Hde/
)efFO<U9NI(D_>X>J_QJL[1<gSAM2Y7.(JG;fTZ@=VI3^WB7T[g8L>>-IW>@;>c5
Ee#P/gU07@Y=HLc8P4)f1L(AVR=31c9#;+ac;:_CN5PYF&KIRSaO0FX4ePWNP0O4
2IFG]5[M4S[.F?CIbJSDHLTe.,G2S@J.T;?bf)3DUb7:)>F/EI.aV19IXTS6/M:_
b_a[H-Xd0439EVXBCd+XR4SYbT;QQJ&-]^R?d2J.Y\ec;_N:[^J)K;H_+.H9REgH
?YIYKQA\]?<-C(6ZZaK<(MNNYIN8dZ.d,,a-d4(?4C9c1=X,).X09#V(ggLFYdDL
:4^J?g8_b?-GJWL2MV=^FCVOB_5W^&8KJ@=,,WScX:RfVFVZDgO7ecKbSY.D]HQD
LcY>M6K^4ZDG.R<X][B&0GB+3E#>K\:RYfD=(-b\&1;>fI=b0L?aAQK(6Q1.>#U3
XUJ5<TA7@.M5agX@RY)KZY;CKcM=-NIEWR=9K9CdF<+T+#-dfW.:E2.JGNOSA;fC
BE#U+UE9(7@2Xb&J36Z^\]@FXOUW.1H,]FVOIYdQ6D/Gb>N?M&E7Y;.[1\ETEM;R
S-S#&?8SQ/KTW;TUbV<Z-BJUd?cCA<IEDT@B2LMXI@B9R,DA@ZJNQ1[D=422BK:?
J94&+g9#F_ATA-g6K<.T)Y>8GgM[T)FM6.K-3A[N82+e[]SEO,LGNRF@:Ca=\Bca
PP_)(S-OT.;@3ReT]dd[Kb&@g@gY4_V\U@]F9(;J.RYdH+E_LcIKbE&c)LeDc:/(
VTaVV;9@8Bg_=BEC?UKE>>+W,+>:1QGLJ.-b\])DNc7-g/)GBVTe6B:4Kf;e;X?V
J4QCAX5bg?F]]-3@3C>)dGV4]YV#AfW8E#bcOe_WZ)c1T>O@8R7S]HMIX3+ND\&<
(7V&?T,Da14G[42a558()H)\\C-)[=2&b1D6DI6Rf+ebJR1J.7&f&<;-0G(]YdV]
>K:NQ;(.cPD-)g;713Z3)Q2PbE0IQW?YQ+8NUK:aW)<([S#f768.+TAc+-]H:RW=
a+>2#0EFTSKaP=HfOPD59[_HY9C61g<Ub@aJA^d2g&eTJKa-=S_TB0La@YVOD(UO
C8fDMR&M&CJb:1gJ/G8OMB;_8C?9FMVeHLA<;R)H74:_X1ITVd2^&;/90-5-7ECP
P+TfS:#J#RS=bZc-gS@KX_bH0DY++(aJ2VS:#W[X#[0HNO+VPZ(IZe2(JI2;D.&L
OOE5UIU.IBggK5>D1/ELQ,>F/P&?(5@eQc)bV@Q@+c5SQT&3VE+(Be][dQNe0H=^
K\VPQ<<Ld?I2;e7RVNf(-@86,@J4=P7]Bf=_CcJ)8L#BL9@)QOee=:OZ[D_eIQQD
2\?b\+ERSJ@25HWW>F1/9.[/ZLUc]=e=;3g;=RH=DIb@INKAGf5Ma<S<O:ZKKf<d
G-&N=E2G>Q++fQ[)11A][X9T_IdF,2[Haf&-.4:I_SE,,B;CI)c059WRc\cUA7?+
Fg.TAW7.F+ROPaYR0@a7TRdM0X=\gYTfQ5ZG:)>;IJ0VTfgZDBE\PVgXN[W@NI6<
[PeS=,H^=VP[G0S(<eO,05cQPP;+42P80WbH0e]eWWg[.80F@.4/NAQG06]3=8V6
K>]HD.b].6WdPaa.WKLff#8<bSW9/6TDY(+1gBXN#Z&.+b4g+UJ)eZ?AeJ4\d]Lb
F)1H6GQ6LZD9<]8NA3F>R9:Dd8d)A_dde-FQI],KfKgZO+>9Y5;?bg:=(a0a=4AW
-BOB;28.0P&cOQb9c+ZaV2(&\DM-47NTd#>POAWJ-7+1ge+J>4=1I2,-:IdKA_W@
#,-6A8L^S48HGT0;^R^0M&e/1ELaA3/T.4<R[;O+(=NCFL^#[H.4#,Be:,+5(eL)
EENdRC38EXN-@LUI<,7LGB#G=.KLV#SXBU+(FYECV/T9A/:_];#:ZE+O03N-+1MZ
edM_6g(&H(#0+6KAQMS;432HYD>=SHd?::H<RY4#@c5>I,Z]RWI.[N;4Ea-JP+O>
_UI]+\M5&-F)=G9L7:RedHZ4YVAST+@G14:8G\Da1GS)T/JZ&I,9Q<f3f(H9NPXL
Z4,AMBZbe#F]/)fB7NJK/ad(^57OHF=3EI,@XVAcJQ)DOB:FCcG3)R.CRd576_b-
5<AN@6OMMY,I37HI-TR7.(5V&aLJE6V<@Y9,T9dVZWO/B?a^_UEfPUe9XHa>)N93
];&?]+&7_EVBdS5NP=?\ae7E]G41QE)DP8EDNeFC<KaV^)fI8,M>AVL@JE/5WZ<c
-Rb_TR>&]K[9.@aT9.ZgNgf3])\P4F<#)KNFYbU17PdT+-\fP#TUS;.T+5Y=D3+Q
Ig&.O)7d&DagSWA18H48^EW@fUTD[3(ISYdE:7RV)a_3c[UFac-5H?WQRbSYaYN(
bdb)@N)MKB\4c10];^#7LEG7QZ-4[7GEJY7d3AJU9>g()e9UVfDP#HWbJRAG#LfH
)_];-3e[#UfZFb<adXN/G@5gcR_V_V7,,1NRJ=7LHM;]6^L9SV=NMR0SffAg@7Rc
d&1/SR_4N7)FE:A18]+K]GJ2M_0+^CFLL].S[8&]dYKW>IU&LP65-+MM=UIf22If
3R@=gf0:b?1,EJFCHf=3V;fXM4]Ea:\bSb/5\QK_.cE&\7FXXDR5FTH0M7GPUR7a
caF?Z7Fbfg[,->;9dR)6+BeYD;RE_A]DY=C]1LbgTC31J<@OVg&2=/DBXU?R]P8L
_Xc(2c4e)bI:2L.GU@aWe58Q4I1f8&+M5e&MI=S[I^E1LG9J.dW^,SG.G4=Od.Cb
\8Y.,Q)DVeJK3DZ7T\TCBO@4FaH(/X^HJ0bZe7d7:fPD6Y>)C<_?=AHYa>=\Of1<
NUE]bcBNN2\]M^8gB8AP8QS2G[B[f0]Z>GG(e+f?PTM>G0QD+#Pb.<KDX6U:3<79
\0YeA4\BK/KL4f2F+KPBaJ]VLeU=8G:2RI0L1QF<:USLg=H/b3\_#YO7@FG/7PO/
W]#ACQc8,G]G[D7[/.TJ:)37MAGQOHRPAXBKPX<bU&Bf_L,;XDHZF.>/>c.\<BL\
dY?II74(FYVU)PUB)6.e+(=K=^@=468F3/&LdDG4ZH\2+cEQ_HI_fU6&3(.-#GZ1
9G]->.P-6P.B]RHaL3R+?1GOV90b\6TPNJc-4gcNF<A54>_ZdJWSA[-RZIW,<LTS
PgH4XTDS4TUHW#ZKdY-S[d@XK2=W.=9-59Q84RI?0Ub>.]WW(g#IY7bGH9-\5M=\
4##VfSE#Ob]8R7.N#D3acLV_2+,d\]@,(S_-8f]@+G<b>EX@FD<;gbUXaE;4G>-#
F2\G>:RCb_74E+^):S[R,9@\0H@Y;R+L)^9A\:JS1#MM;CR(dd(e?=g5?RF2OcZ2
)aBAYS0e9.)=LBWAQ(Ibg#9aLePc).<#7-OVXOeR2S8\PMVd5WR@:cE4BXgZcEaQ
BKPGC?-4Q,AQTPU73>L@cLQ6=O^E(V-_B=W_E0CgXAO)X:YcC239R7J>7W6WSMSA
4&V]?3+=.7R2.4H>37+WP32\FI[J(9,?V<@AGgJQ6FBcY/_0W]6\A_KYMXV2+4f&
HC<=F)OfEA^>e#UIbG+HZY]K;5b_FQI)@X+bGJ\F&[/,-)d1@11Y]aaF@XWCV(U^
M=4aG_E;JMHB?N_+>)R>^X^)b_,+25)D@0N6DE]bQDQ+>JFTZ>_?1#?)P=D4gA3c
&0M_<OO<3MA_GJdRXOS>O(CV)E]U/ZR]/8B:gW&+RR6[N6DQ3SJPaPUDBe5c>7^_
NGELFG,0S&++WB>UaP#DeR&&6UB33=Y86E]Pe>Gea/OC#AE7ALIG15#0UTUN4@KS
-EQ:^X>)bU6gPgbR:BEX+B4a;\RQ+;\OLIYaU(Gb+[P4=QO5C/9,g,VAg3.PGec5
8J)AZ_O2ZZWA7:E>3_E4_W0?AI7(gM.<_+EVI0#>^>(6620<FKGb4cX5R3]K;1U/
G;eMXa5TMUH[EN5PR0DD4,\Y5&e-L,2bH>Q>9#=;+Q4Y&@W;X=I\J9fY\DY2O5[M
#6C&f(-5KJ:HL9NYL]_A&P?_9N;Z+V90@V>[DbE(:.S;<JLe9Q&^^D\@V/:bL=4Q
BOfbSQ44YPL7\ONOWJAVGW9fe:^A6dNO125ePGQJ,g?]M+b&#+,3ZO&V649WSI5>
bMH7_Ma6=aYgF7OG@/Of[M_(QN(=Q</agLPN#MR/ZT(;N??ZRK@MFLg;S&IVKEME
.8J_fN5T5g[PQdV^N_8_O<RP.HQa3Vb1)=Q#[+aCc5MCZA(-(2ARTWR=>aa>1.TE
_6,N9HM5]3dg_MaIIZNb/=aZJ2RT[33;SI2B]I7FY;aADLObMEKTRa^C^N\-SHfK
1?e@V[I0f8S/WD&@gedJ;988;BW-)Zb9bX_,GZR[CY,G<>2bWC#583;R9L8X.=LS
aK&@:<&QeeP2,>PRS-DW+23LI?CC+2LSc>RWCW_,WG?107EW4Ld(;>Re.d+R-L:/
[472L>N2C^]WC=Sf=gd++-9I1I5#-P8+G]LfR9=g?:DHg(2dI]_W#2.0AA-010JX
XAE(B=dUO?b2-g\R=./O4=L(Ea9eDd37<A0:_4K.\GbL5EA]HgZ=HP(K#CgZQIab
GKc/B,E<NE_LRF:[;T_e212gI++UG)4XRAN-[00cLe&8:V,V:O;EF;:eK\U^=?a3
CgNbTEc+Yad+c<B2&W;\f#7ZLTf1\X4GV5Z3@7GB#GULC7F4C8A#]#_YYEUOPB_.
bJPeTVZZ8_Bbc-f0bcEA56ENOWV:#7@BAP]<d4>Y,10FOF&:5BP;Y)S32a/CH@;Z
Qe->E5FJ_(1b]C/Vf^>#)YK3fL)-[FZFZe<eZ../,70(93A]eLX39:;ee=,CcVJS
4AEME+];c2M9MN6.M,_6AFVB5d)BL.)a0X:?gX]_9/d[]>>4CbZGedE1f0\-?F;H
(;-d#B-^=\aP0F5.SD.C.4M<+J..Q59I8/[>I)\[D4OP3Q.R]IWFPIE:)JIN-#,I
7&>)Y3.T&BR^HM2aBRIK&C_6RNNUeP9e6?LbgSX)@#>4QII1^AJ;1EK&g0S;OL)f
@b-1,PgGNYE3:L_IJ)7gV-Y?A&1F0Z1,\(.R=:^1-WR=.,M+BMfLY_0G&SS377@)
eR[aMLCa3MGX8+0[D6]g.0^<5G]OgF1GB2&c-&A<QYYP_d+KLW^c\:N\AU:6G@&U
=DfJeaK/)Ea7-S022L(S5=cUbMLH9RBR_:F>_JH_MB<]9(Y9a]S&HS2(UG,9c;:-
/bV\aB@-.YS;[QAdPg14.<@E<3EX:N&6IWO+Y?RZDKG_<E;=RHF@1GYUUP;O3F&1
Wd,ED?+)H-T:+3NXg9aHb)eHeGO[7<gcdU2(C?fY:-DUd@8<Y9FGSV.T5.CY-]V#
/[e5S+WP.@VD9J(1cLA?DDddA477..70)g@9D_VRdKF:aFVIKb#Y1.)#1EL&0GO.
L@8D3U5J])/]^gLV]Td-Z-/YK93/(/=/.Z8Y6@VFg:8WP=6PK=MT4(C1AI/6,C1:
19YVZe:^PU2aQe<d,0VJ,L,+eO)Ta8<K8U#+P&X#QL=B]&GIK@9FR:2O0^ObRR,E
5BW+R/VY,UK8U,<cQBS\.aD0\TCa/[BgM)@?.-74A[fKASB;?If7ECTgeRH=7e_a
WNAL_ZN3F?2Q[f;)BJ:ce#Ne_M>d7TXc2C(O)#P-DJe5KBU0FFSOJB,B@fg&6_<D
SU;T&ZV0a]Ya,-f;_Of(8C0/b1DOdN2;1Ng?09BVAJ?Nf/-M]JD^T,IC<RFELOZU
;=;TDb8JVgQMCPHE,&@QB:<NX#[HU6I>V70SUL(9[7S[D?fa<UT9IAQFPY[#K-Y8
MY0bI??aH>3(Y0IA##1THZ8fFeTP_>FR3VW-D\g,)3L^e,WUH/58_Z\3>OM,0)0D
\\Y;S[dQF6(KALgfZ8ae./B-10gXHQFEO&-2[Y:1fFV5_4C_H<Z4P<ES>/0#d1b)
LN8W;LYD)=C#9(0T&PO5I2X8Y,W&LTgf+b[#3a(.Z)TO3><5U(LG/(?LD#JRc/<P
@g1LDG^G_7QD;g:?5I\[+FC3/3#[cAKD_+_D^B9XD/eDVA5dOd;Z^N&47T^-LV1;
VT6(6YQ=\/P7CBbbAE#FbdaT@H2N@TBgK.OYc3?#H?>TZR]IX2MS=W,;=(7N^&6A
(Qd(UDfY;JUZT>#eg&ZdPP-XD]:.MD]I^34SSP]Xc:,))fdJO-RQ#]JHeAg[,[?2
XI+KI+?J4f2\;.V.T=.]\/N/U<d+d.^T#\,Lcg>AJ^__8>Pc-OR;XH#?W13cLP8Q
a;(:?B#4D1^I9\>+B:d3UC5D)=P@QN2GY-I9;1@dE7c/OZ0A[,\Rd4bZZOD3.L4:
dQf9[JfO3E;C^P#(VE0>#^.8K_>/N0J;V-ACaT>;d\a]@cd9[W7,R5+W][\L;5=>
6]8XD?,S]/TaT4?9L+(BI>G6E5PK,^#EQXEW+21V[D_LdNN+<W+1I2HEOYBS;g7T
@WX3:B660VK#ac1D>&T)J]&M.Q4+XO)=(W&UW9D:]<eR,W)CD>0W(ccA0A]RM)QG
GG=7#QMFY-68Aa](L+40>U67WZb23K=c6OIGAD_R8-C(2PQVNF,^bRHdUa#UPK,g
I=UPK@VQe,_F9:Bb?]NL&)<CcMX\8429aF>cKcA?KD;YCW(M32G:ZP<VIM?-;I/[
C]4\0aSU#(4-&IOR/#QP<Dc<(#WOV0Sg#a07eMZX/0SW73Yc4]8bIWE/HPQ7,(2a
_eb6V9If(]1GaEU8aHMZfb6^JFCG:824OK;XL@LPF>Q(Kfg>>&AZ,3B:FN<WL:MA
IL(f#7AfgeZ4^V\BP]PA9.NTbYJL>C55?)c(JXBSVfe:\--B]UCe_<-1-B,X(EC-
,=T-TH2,A2D[POQ3=:U?;Y0#c1#Y0R65TXRA\b&[8B:9HfGEaA4IbL?7G9gVLBHP
S-7@EVeCWdJ0-,b7U&>R#7AI[b;AF+;DbAbZ.J.M.LYDUgFX:M7Y;;I/@dS+R=ES
OUUMG&M6#g3->FW<5QE;6M;A#PHDD^Y[O)GZ4K8K]B5G:g]J2SV6-8HJ>b&XO[>]
J2<?83_FY?NK,/=4):J+e+,RIBIe0cX,(0>0X[=,&EQ[a6,0a..Y5CQC5d3SWfF]
<9_&XTPa9E6ecdQ,1c^c7W-2_DCB6P/3c:B@.ITg#-A4..=KDa3^F,WDC].&DN<N
TN&24ZGXb?F;:U-&<0\KHZ6g<7[.U[E>D^&KC]CT]9UCH1UC^HBLS^W3?,gdg+^O
1b<d(P9(dFH6W?3K8,Qfb]H9M^8Q<ZMV+]6P;Da:U<^FG9de[NcQ3,P0.3&,5G+U
B^>Yg+B#_7a2b=-?Sd\F2-HaAJgO):+K+>R&W6(8,C)(eJ\AMWIVfYUTLC<BLDCT
I/74\+_EY<])^K2\c\S:.V#9gS#OK985,T7JJ_-V#PC^>a&C>cbI#E3&GX23Jc-V
Z01Y,.U/Bb&][cBA3Z8WDAX=483F].B[bH5<PI]Y^B.gMGG1:L6J,].HQc>-@:^4
[K@?8V[7e>ZVeBL&@9J32?/EBf3-\>b=06^88<H?^NY#S5eUXQU4d=af)/8,\N.I
dc9Pd8/5U9eY?NDWTE8DaQ)OVQB0I\1g)A#@f8[\(0#L&+6/SaQf=dYH#I+0F=?2
;F1G;#SA00+<dB&U:)FBFNBJ2<F^6eY?cIRgXKe)P7UAM6TOJE7(EOHU<8G4g.D7
F?2Yf4:/>KF=.:M43D^b8@d[8bTEc)GGT6Vb-A)Y7KBeda8>+B=M?NDYbDe_6+La
E-0a#DPZ&C1_R#02a^0C<1J0fW_>PE8^>_3?5Q7@G@9a9d2BJf[=XXb_T<QCb_[C
_.;&cCa8dcfAA3/@^;0]O_97\:Zb:<GZ1),DR3<Mc6XcL#\-(GYXggNGXZI8MdA@
B47bGdG8<7O1/fWF[eMf_?/^gMOB42YKcTU;+,XN.>@E6@IK2@Z\@QWI5R\>OX()
T#XW?A003//).W&#Z=@355O<^]EVcMa]P#KcAB]VW71dWBBHbQELe8N6SD<?KNOZ
A:AC:I(L=5aI?IOa\U@W20++9ZbMP<VG+>=P8c9SQJ]>fe^L7,cg=bUREM_M_ZF/
>KgIL)C:-c5G0IW\UI6M=gH.8:eKPHPN?d+GG6[K1\&2gQ2<\[@Z0)6:aKg+F/?H
OQfT(>4><?4.9]=XZ/VT3+[6agHSXaTT1T]/#82JSPP)3\,CV>cEMG(,Zd9SC^GO
=E4AfOMO(3[M/UWVXY\A07>.B\;T>E-2Y81.(=U;B;S\[IH(F5X/4NV&((=>X=&D
^K.4?RRG<,]1gUVK:Vgb;cRbBAbODfFLC/.\a#6)6P2YB57/FL^a8WF=3gC4(BVO
Rb,S:)H^#:@P>]\SUV04MR/W<7T7T3DeN+W<=DeR08M>Aa8(0,4IHSB_9+.7&dHU
,1D?1VJS1Z)?JJKYcFPN\eP46B3+&_]AWc5]_cd70VDWFf7]8&+/]NL8NG\>DRf/
EAb6XT05a@VMJ(><UCYTE64T9BZPL&U\YabG19ag[Ve2X7(^[DW#I3dSbU)O?]RL
TT>#4dGC1@,QQa<G(YSI7(HKI?O?54WO2UeFW[d96B5?LL,aM=R#KYKUSHI:/\-9
YV=SW:ODbb(45\8,,,ObH1OVSF;>gMgB3\9JB[R@ZT2J(U1+3fT=@a/O9JbHJ5S;
D[>8HCE&QI1S\DJ=JC872IRS1eFUaMe8/#,XX0@_e[53(c+a4?OH[.<[2H2?SFd)
EG)4>Ke1W@ZSUELc@@T@MS7@ZEc&8IBPaZ2-5VCJ(0+:8B:f/O,+8QBR&G;CK7\E
Rf&V:e=ISB91SObX0Z@[\1-F&dF+R],[C/<INC2DG6BG].aQQdIeR)0@_P]cJ[#8
3AAC+><UVU?1f\9Q32ZC#@\)a89)IgYaVE]#=A/2]-H2]P+[X1eeDANZ@)D+-@-7
AX).4F+K.K<UM:E2S?->2eQ8(&M>>^S_K]b3\&OeD<X__6<_B^IP=V3-R^f#TA#^
XL)_g68A1FgY]T/FfH6CMOI#fB)0--8CHB:JeMI?H<cf)OXK<94IL19FbY?1;I,U
,,654#&<_]>UHA<;5VfD(Aa(FZS=1;[dM84/V2-[I8c-b,#6KW-PU:X<b<6TKN@#
4aQ;[JAO+>bWYbD)_T,]A#ZG@PC_\#0H5L\_7Y3Fg;LJJ-PR6E3U#fbPU6?-;]/3
-M_3f;Id470D[,aT4aN.d/F>Q-^_9OGc2KH<=+PdaPIe/[QZ4=XS^LYV>R9/;I)3
C[cTCU&-_R0;U>WK0@1[@Ed>>N+F45<UM_=7gDcH=U7=1DOePHHMg]b/))&5H(N=
6/a7?K&\>)JBY9c4DIG8]N&X:)T.FW[?f;DLAZ4[NM\WX96XBNc5Fc_TPLM4AQ9b
7]NUU+O9U52PUOBL+4(bYIR(65;8b.RXIWR@RB9=f3Y4TGW88Uf.d\JKU=O]cHQ3
6^ZD\Y)J^g3)L>56F/7H9K:ZR4]ZaX_H7?-?g53L#G3Da/3K(20:L;)KPGQg&Y,\
5J_,VRc1I)gf&V9gg6cGGaY.MQYXV6C]-P;?4Z+^4IPVL\)J-B6TOa65I5YSP,++
X_]U,ZQ;5I5G+cF?E+[1@0bKaQ\.cZ3KXBFaQN5RPJd/WXeAa8=5U<CO#1T@ad5\
ZY6)]_)A<?Lc5CcX_2(fD<b3GGA^U8GZZB\dGDJ1_L70OK>QC<4b19DJ+dZAWHAA
BM-K2B=/0/?I>cOJS1,90gfCgbg4_5)?NG(-?00K/bFMdVEcO(4g9f&I:V:@6d[U
9gdHKN_RL)V;HNLB/E<D9dBYD_EODU&L2?egGd+9WW1:)g/=;1R_4/D8P,?O;55D
NWKQfU#c]d=Q1(-7Qb8(Me8fI,SY4Fc0<AEA^V\/N[FE#=F+Y@==8J[@TKaa5eT(
)g4Y<K[FaaBADLa0/7?DH;XK4DNB;ZE36]R_W0FMZU+UgMEdB;#46;:4V3R;X&g<
0SCf,a-gbVZ]N9<d+^Y1&^>=cHgZ\>.&.]H]3a-=4A)F=[ODM#,[)P#^;NdD7-R-
^F(1)=YX_64W>Fbd)aTY0-T44B;99&,bLFd<.:/,;g:SY^B?C=X8B1@b]FC(<M[/
G,?=(^156+/@<^YE.IeE]OWXe+<Z2]0UJG=TP(^(gTX<IB(9g#,8EZKJ;G>WWD;S
8;YM\WP0?4A3eSSP+\2+gB]Y,#F1EGZS1dD_\G,V#-(<YAcb#cB@I[.ODR4aR+(N
.T.]./OQ)OH29?C:<^c@\,J9cNSGbMHKRU4./\E^:0aK#:?1aP:N(0,gG4Vf[=Z\
BH5:OG5O1,fb4d:+5I<0XA@^.@Bd6S(-^gM&dU6/5^AU<ZX]^.f;Z55C6?OK&8fZ
F3_eYT#.aaaW,DaZ2ZHG89&;+636E)R;bY4Dd_-E?3SMH#(/gG?].J7Q7f<40>MG
HKLCA#g^VQcEg1[DGP(1C3g@X_(L+e#b39Z1VDJ\V#6HfZC,59N,G^aPW0dX(#<(
dagcU/[W>-FbYfQFHdPP4=L@1eEMWPTG;a61gb:ZPe5CDae^dJZ:aWG974&8B=:P
>g6-&GLU(fK^VUG+G+b>.VU>(GQB?=Y1IK34;@/]eZ@FH@XUA1bAE_(G+/WV&VeE
J,eTW[T:&cYAQfE)\K;f;a4EZ=]<e>-#&ODKM__7B5>c\A[N:76g.;+SNLcV?_D3
B5G@ebJ_1TMaN><P_c=-;95c\6#.@e0Z[C^UaTZb\O&.Pg8NMA.DL+Z<L;fQ<]dI
:),;:gR7N[RX@NUQYMe=UM/VQ]&+9\CfAH]Nf;aW>2W9:8D(.(7A3D_fbgL_9;,2
\H_G)B\]S:?.B1#-3M)Z/H,Z[I-+eUT9#NR0N2.2K-ER5@Uf(\T=#LRV/\QIbE@Z
^PS5=5DP+dA3]F,D)M+3]cMZMU,afY/.>db&DfBK1c\[,-O57PXJ7<XaR:Y[F]OS
Z<<AaBP@4VOIbSe1e8-SYWbJB/08MU5^\Xd3@LaO7)6/Y@0ONH1XR6b2PT:f;4ZO
S7K?>39_QcX3]f34,YUOL]#N(Q3]DCG,]aaE:P173D[BAU6_1eUJ?NG.RG22C9//
ZbMW,HSL,HEGN(M4(GId[T:64@=&A4V[S\V=P1M,D1-[;C8]\OOW8RZS48RGN[5:
)W,C4.6\NgEKcdd?-QFgAN/Q(\1WIJE9:M\e22+CV\>?c8JT-:\WH<,18I.JZbX;
QDPH43UJDE,K&OZ>d\[3;9IFg?4^e1f?Q5XaD?@SNNa0J47#Z88^A_?VbdX&JD+3
;NDPgWMB-7#V2Z1b=X(&Xg<,\[)g)N,\gM0I\+^LC0=ZAU_1MWW7>U#UJXB^<bb3
8He<?C@:;dE)Y-3543=[LbV=[=R0_YS-1eMec7AA/e/.6e:If2M2K;^6;_L0TT/(
T0#b5J>fX>C+,5G?eGU/#.=2[L8>WeZ;-;_12ZDS(S)JHg.1+G0FdA68Id__8Gd.
C#>=Y]AA;9e\-OQ/A]dHL9Da1c?NC659Sc#.f^[\RGfLHA09XW)5R_dG).?12>H.
Rbf_LcM,(3]+Od?K8U&SVgfK)F-P^<S52)I2\6BQ08ZLR=1QM-F&c8^WLB[0D,[F
08Vc/-RTA;CT5;4(@PSTef6]#\fcJF40&8>+Z21Y#2a<OY9/ee9VIWOZJ<(7]Q&W
&HEL9-&S?QcgVa=#PQC(3cZJ]JQ+^A4]W95>BD1Z>g@OTdJ1EgGId#W?][<VUa>Z
T.c@KE622#b=0?@Q=.N62<<)U=(#UFGB=bXR7VE<M&.bb9cGO0;HE78DU7E,WTFP
_E9[cG]eIg7+RT\K7AgPOXEPL+M7UTH<?Z+2[LQ&/(=R)d2>0b-\JTU5MSH4VaL9
[AQ(7d=:TNKJ2WZ@7f1[=_9B/U5_JB:T9Od3KW7#ZUbV<YD.LKfU=_Z[Q>JB1:11
@L^V#?d+674Q#<VVI]>K<1OeHbO_0^7#H@@L.bJ3(ENRY5_-.<4KZBXM4W,(^5@@
<g)3P)^_?;C;cdIZ+_:bIe#((;C>LF>D^U[D#R\:)K112=8Y@>dB#^U^DOd,e<_V
J_^VDD/4U<X/2MF7,=>Hb>8c+&WVC=NSJ76L6X>T+NIDSPf&YF]VaLN4^?Z@4=P2
&)fC.AC4F7^b4\\(,CSZ9P<T8d^IcTb\+-08-?#:Ce)4(dE08H//_VFLd,BO6(,f
.EU&P[Y>f<NYDJ;UR1T8X70Z7C3cdE9de,J@H)6BIUWO.CD+=I__BJBX2=PWPFWg
JH_3@gWCT=63Tf5G;RT]ADKAG<]0<2UY<Y[1RV:4.4E,Ob>W74I38P9?<NYaXM<[
daVe3#;?2Z&G@0&MRce7Pg,e:#b][:5V]^HFI35<N1;DR+#1:&(DJL:G&.YOARDN
3@M&W=[F&B,243=<ZAOe66e2+0(^L)8aUAg3R:N2(J>\S6])#;^K?&RBBOf&_dB^
YLg:dGB2f7O=[750_+6BS;PZE]#gN-G@@5W:?M8#\Wa1;Be>:ZJ/DHTc>NGY#AE(
C@aHB6f)/UCF#7<6TXE3aA[XXZ,OY4V-[@#)1JXgK\:^[d7IT(?M@]N2C,#ZcXCD
3E5Ucf0-]YgbaF_Jc2(K1A3W_BSO7]3PM:6I<IMW3[71SYfTBR(S0E2b^B6\.(-)
JO_g3dP?QSDWb)9]c4\HcIc3I#BTRLY<6gHeddXC:HTc,Y6-=9^1KBca52e\K9#6
5:Ta+Na1R6@1,PO-9UbN^>EYC)]]<F^7(,/&4d+>>MGH#Y,O7>/5?CGOI?4;GeaW
T<Q;)A=CO;U5F:c&^-[[?CeYD5TSL.#2R>/9Ec3_7BT01WgGZ64TPN>-[5?K]VbS
CIT&BC8.FKa270Hb^.4=WL&_?^,-Q3777X).^1NeaA2L_HaMPC9)GHR>XXU&&72C
XV/42V]K=H24Qe79377FD[,@#Q5EgMg#L];G1M9:Efd1M?e9ReGNRaP@:1YNH2Yg
;g:NL+F8=c/LYSF6VP]^QX--QUAPK(:6E/BbcO\0Wf@BGdLAG)QL08JR_WD21]/B
KY0YL?b[&NCXXX,#<&^fV9;?&FE/I5.CeCC=L3f,c_-#,NRWJ2B&.G>AH+Y[da<L
aQ(O.]NZ@YC=O2SMcGHaL0@X=O@:W-=fE.CQ7YRM=9/1ZeEEUBB\0Y?2K03L6<Ob
N2?2;JQ-..,A;5>,^WA3:d3^FTOCO,3S5@7#+TbMANT71?&;LAW&&A_3EP>d<K[:
8@Y1M@f?O;-Efb>5/J0WUH0I[4^+c#S6D0dB8,S(@_ERD4L6[QBPb1\P[D=Zf9BW
6HdRJBSWO^7Pg2PUbR?H/M0edFF^_HD1X4.-5&N#+W87_6LI3fC&R&\R&\Fb+a^D
gF07)f)F>6^75BXSK;cJZ,G\:.W]X_.X1@>e2,[ge1ORW(3\UGYJ;PBS,B.Hb900
?cQPB<V[d>gU6<DKa^S#^Z&9[@Hae@IE#8L5ZB^gd4D9/7;+cc.e)d@UGC_[#b26
1T(VS/K,O-ZA_?C,E]&(<9ECKMZgc2F+H\/cT;GIS@T?<W]fe(Y_I/eE_TP6cOY1
,^TDbIT&\QW]>gN&^)B6.^B+.#(&](HFe_WE-9RgcZ)GO^14<d^7?(eZ>(6&-;E]
c9L3PHeO/,^NJ/f0404V4__<Y?d#UJ:\^58=GE:-&/:79#:I2Q1,_UI1;8C5]U/I
D_0c7I+T(0XNRC@]?6Q+f9GG;dT1B=6J@71Hf(F8.Z?7#DH),_WQW=&PK0Z(//X6
L(.<LaY@I/^+W+8:\H4:D&^T>KUbBF5XaMcNK6Bd87bDd4KYgQT?df]WS,fe>e:b
Dc#AD@dJ.QfOW33/^4[I9QU9T,]:7bJ,[OE>-MW3SHQ1KZF0O_SIef:c\+_[a+3F
G6:70X[RXCT&#^e(Q1MKV3Y8IELD/c7Qb6>A#&YEcX:@+M(\G3T-g975a5BQb;-e
8E:5PDBX4OJSR@T:3dPF>A<U1<V=3e_S651#Mf#QT6BOa<4(?4+M11?RH\a)2FK_
gQG+X6cX5YB0^3VC)DL^WbCWX5ME?[\=:N3WFM>V0N@D4VcL)<W&NT6f,H2c=1e\
g=,3<DcUC1LAX.^=fV:R#93T,JRW7?cMU/:U@K@1(>Ce+[1//385/C\S6,2([gQe
b<PH1[:#d7FFd):eOZg75@afU]42TAQ8V2<W_b8O+M)bBfPQVJIeb.S8?[R[(.AI
g9T16cg9FM-0a&1T0GG#MKH4UBDHXd64,P:+Uba]8S&Gd5)+M2\a0TP.S9=7^RMg
DG/DENVU[Ad>\<>Z>N_>Y/N(;[N_4Ib(19:5IQdVIH#,RJG45N<9XR30.:4F9W.b
57<XFT7.3_8=ac?fYdN/G0W;Mg20@5b)0fd^/VFU:c1@b+^+fb?CT7SX5Wfa>OH>
Tg<+^>6b+[aOOZJRVf5D-+H5/bX[#P:0E\/D/+NJeJ78CCKAN\R7G.-@gN>/Pe>8
aR&cRY4)WaW=X:ZVCDfd3I/DM(0T/OH50#_bD9_1./g66GfE(V9)IACSB(,&fX9\
A,8=CGJ93P-C:>YY]#2He/PDMQA6RAAg3G<#XG\e)gFb:eVgL5EB3)6F/P?B#JbZ
b@?60>U>JE]=DF^W^3a:8J62]S#Q8Z&P@6=bL8@8^e>[/3-_S&B9/FA9\aY/X]6N
]O&;CY:K10P&?0^&bf@]J2dc;>OIM4?4UKCSTdX:dYM-?,W07]Y>J+A8HQWfCa@\
VF5>JAM.g/L]d2WScGT09(dN3]7.#=fH#\[\G6;e,>A(J:H[UEL90H4cSO88;)42
0c2=U,]5>eOPZg;<C:#<4R+f__8,CO7.WQD_JU?V6)\:C#X:7AO?^.CgB,^V:)Ve
5L@3#0EW<8=.IPbDcG^+V?c_YL:9LVPDJ43O07fFF;./RP4>#Ibb+>XXH+N]S8.Y
_H0[3FB/?P:-TAWg)ZO[,?bBH,UcM4Gf/U\4Z3EI70d\ZO?][H)@CV\3aAQQ4E1L
?Za&LJ3HFfYfLM9S?dHSb[ZL/KM8c;@O_,O]6;[LXW,AS9Y81]:OaV73Q5&;^=d3
6/TPa_AQN>_#B+-S8&^_7Cc5]Q(XX188/VLI90X&bL4#QW4I/gAIJgL2A8Z=JSc<
:E[02)K93N#YE/JHEE/NJRa9K-JJV6JCbdgRP4/[.]g?^3:+45BfH?2aJFa]0MLM
=^2BC.-U&R1\)[Q[.7,7,R]SM]54X3ZWDGY&6:-O(R4GD]YE8g+@=HC#a+.6ZZ<E
9)\Pc8[c:VP5XGX<WV]X,#=a4CJP>1gM4@<P0:A6dO;gfffd(MbD28A#^FI-:dWQ
.0YM@PQNLYT+.7M,<A;F)DA@e.I]1cU[8J)cQ0Z)JOT]?GH?-Kb6MUPBY58fd))3
=NF:g>R?FXM_<Z)EW-FE-\^H_a2/WRSLa[@EPL,A;(\5BTX?6/+M5TW+VggUN+0S
F]^DWZJ+J?<XCdWURMA1?(BDD\W^aZD+9T_TOVgRbNS[H7M;EFLd=CEAS/6#PI17
?>NXJ:BG224ARG8]+KRS<<X)HcaYQIg,T^GN[/=?0L1Rb+;AP1Z;=7cE;&X16bS.
GU<c[MdY?^1I\0d[SDHP@EJV0D+KY08Gge(O</C9:?8aFNMWXeSJ5MPEG+/c?=?X
Xg11XC\^6+KBcT=6?cWM8YQ+<=D78Cf,7<TcW+HCefCg8DZ._)HG3.&S1dYGV#;B
e1LGLBLD9JGUBG@f@DN15]6bW^Q\F>]dJdC9@D>A/(]=^#)QXS?^SgW9]6N(M5+d
9BV5W\MPY-RHe2P)\W\8aIX@EZ^JTB6]>W;fXae9S>)0E6AZN;:?L^Vg,_.:+Y#a
7(Z3J]^A])^9^]>D7LSQ.-Y.7:7EP6@cfFGK,S#3=O[.<B-6(Y:QHc];/:27>IH?
f&-+:#_<@e+\K<Wf_H9BGe[da75:(R_T?P(4)<&,T6B#c:TGUE376I)g5bI^PRdC
IS):b5&PR@^R4:Y>S1I<=TQW#@2>UPT^JS8/1_.M6_3:\b/@L(\:IUDFN/.NM-?H
DU156V(b5S23XbDM&<ObUS62c5,<I9E<X,ZN#M+J:C8P-@YCg/M-^RN2@NJ]Ma<E
Hf\?IgIeDK0)<@F@[Fg4^OZ#=2<R7/\)0f8+NRfMdBNaA@G2=AMG?2DDb]<Z2e8&
L3+O-.geb42=J1c9QL0<A^\.R-A&YZaf3(NVLM1<1f7=&I+1e7H\1=E2BU5)TcC@
dJ(JGdA__bRA5MAP1C\BN2T:WI7[cV1C24f=>C5KO#BLLb++S26BeL1?g-&HV9Q5
cERD=I^+\7UK,L821bd=#-d++).X,_42[7GY7bUOZ@LAXH:e[1EWWZ_7ZU;_^\&,
J&C7K]bC3^>5G)_?EA#Ne&g-:0NR_)?,?6?V.6c\Oegc2O(Nd].WUO70<QORJ)5T
PcT^d]Y,K_g<68d\B2;_(F,0C_^D2c)C,W>2NYd9]1&-CVS3(Q^O6eX16]R.@WcH
OcDUN@7XHedG=#WI3FALV3McRfC+TW^.<HIKB#Nc1;]RXf9?8@[>V]R#F\;JL(XO
cN^=B:3a.?FJ?4V]BfBN=[1Q4/V2Q1a946=2DXLUXYgQ4C5_Dc1f6fB5Dd<>:-;T
^@g.M;Y1e<DKK5<T@@2?AgA&/9TGL\fT(LI^dSJ&4,/L#<AY0Q0O<F/dCgE+7(F6
Y4A_WCcN8)Qb;-B3FS48IO=J)EaZ-)R-d25IT_]9[9A^B;GQ.48d-f4Lb^=>MYYE
>C^_cG[?;JYf&2:-GR9R30Ze]ET1[+@N)8T6N68U;8,dTTC)-d;<Y6SF7cKaTRe]
3O0+;^DR?MfA/B?f737SUE[_P891McWFZ3Y54&#&e:JMFVaSWQg?gCQ;E6S?b8?I
38R6M(N<53=H00aCF(FRLOGZ\&9XKF15G#:NB>0;EG]6T,^L5P[H9,7[5XQFQX9e
dS=gg?5S?79b(BWZ:DNR<7fe(HFU5,=[&TW^B(>V>+c3.gF2?QMS)&5&K]gU;17S
UO@>Je&:W46e,?-V7AU0IP>,cM8OES/.8b8CEF=HB^?d-6-6UEdL93PJ1(H^(&KX
9[YO,N1.cS^-8&NdGK.)H:O=.H2TEI_]T.G0/,#Ad\g+C-_RS15aS6F7_X_U8NS<
^gB5<FdeFBFS;Y3Q-EULP\EWVa03ODX4:A>_a6R(:@#Ed,5b47@<[3N1QOA^Xg@(
\2,NAP]Pec^[gV3G3P;4K>)0\@=Z<]]DC7;b5@0/>R#4R.(&)VQbX5bAgQX5Z<T]
VD6[\TVJ,^7:OLY]L\V95O+D78FeSBRgH;G3Ga4DADL?<a&;GX9(Qa6YUK?G1R,)
Ca?MdbbZ6--+XP]I;R?JAOPeOe6c3I;UV]V2STD0AK;/W^.fd0c&(^^8&3H?ZCaA
GZcYKeAJ+@MGN03gHL9a:66DAKfTD<e=#,2,.J0ACe99-1S[.f8E3_+4+Jg+):cY
1X7_\EFQND.:-7/ORS>Ne-=BcCD(W#)S7Ea/MKCL:(U^g[TC1Z4)NA@1]3&BadUC
ENHD-bf4?@^&^KX_#M,b?=PQEd9<:J1[FX_\;.@R8YP\;M+aR_T,F/aGDfKE;KaS
ZeH9A0(VT5MQAPG#FWR\7RUCI&,C2;GG@S2>U4dA4:UJb_eC+JUQ&TFYE[aGJB^5
;:ZC2IVf4ID2VO5cQFG]O]B88K_-Y-a5Zd16_a0;Y/<U\K=dHU23RP?TZ_9J+-aC
^5XP4@E7::-R]2F,?bc>]\V]A8#SUaa<_J[J\-)I36CJ<[M/fgNWHBLMQcBFN<A6
BW_[AGcYN3&Q^S@3-\ABIL]A739HN^#2+VJ7dKK7RFgW?96g[_>O=DF4PW1;Kg4?
+USJK4@HUg<^]R4V279BdfWOZM4S7:;F<)2/59_07ab^S,9PGTC_B,[[R(_)B=CQ
f1;7@f^R-UY?>HIGFT9e00OJGFM?(S7)EQL36S=4^C9FN>6;-^OV1I+CS,<4@[-F
O:Z-0]&_SaDbG++HTS#O+b?2+K?^dD.N#=/:ZXa_P\?Q=YZ=]P8KT?1S.<T7.]J9
4Rf1Ff(aHJBD4BXff5a61\@aUe7HRH-4NcA?-J5A,6B;,ECYU2OR_Q,\=]6.QR^c
@+7\OQGZLZ60DW)9c9Y/9-64WJ_;G2]1OGO=cI)S1V2C=(M<(6db5BQWZ^a,2\gV
Z.LQ[d#^.aaZ6e&cTdT?;5N;#SQWT]XHeNcNaf?#O,,RcR6;]d,P4N\O_=L((JdO
.)F81Q8<_A.Ae,<TbGAB,R^H\F36ACP=&N,-:;Kg:GP3;Eb4XdW)5f:aB1Vc)[:]
]4gSG-S?EY_8\_Qc_NCd&BL0I4_:gJ+9g7(Zg]L.S;d/-RY8AF8;;XN6LTfg?AYC
3\9G]]>9dJ?K<S4Ud49,MUO&A55G4T)48J>:A9X6><XT(7<=;/Ug./WB(dS3[.0N
Z_\c8O6Q-cGc[eF_Z?:16\-DQfd-HgKOUgSCNEL[=,]8(B3-=,4RZ0,X<,_SUPPM
_bQGY;R_1WKCU)ZN>/L^;Z9IBcBFR7>/X+CQQPE42[V5Ee(LNB3US+Q1eR2#Ag_(
J1485_LGdXc<\M5/KYTb-X_7(ZDNA>T>&YCEG?C&aBFD)8g#5g#97aNQYJZTeIVb
Ad,WC2NOg@;R&R[X31\dCdd-?H8&IBLRRIbc_a6MaVAa/5F<Jd4f4NCB8fU#4+?a
3XR/Q<W<X,]:G(:TBb;U:0GUUR1A;b^-JFc0,)gTT8U7]@<@CWCW,A#@agY_d9F#
GEW^;QE))\RI54]3&[X,^;00+Af@\M_+<7EbGDf8X.-:H2GVA/AgdgfM<<?U<XZ]
<_NFX7#.Y39Q^PbVL0>_PD^D_V8T^5-EW>P@3\QM6A6MZa]XQ#QQ:Xd/UKf?.C]F
7N&(=7c8U]W=]1Z9W(>];OOL][=_MBZ9Z9RV4D@Q56U56K@3\K#(HI=dG2Fd\)Ue
K.4f6,/+#RV\8R#6WX>#[:D0719=N,,PJQLP(KS?b>fRbU0=Qa5M0aKN@c38]\>G
7PU_D#P<K&3VYM5MW(70Bb0O=,Q=P5<-G]>KaUB:fF#WfHS5=/I_<+_+5-J\b4SL
25L11[GQfE1.@f:+SU<f8N\:S)?:^D-Q#S]);Z1HDaQ9.WHK?7d&YbLN.YC@D;20
D:/7BaX\b2QbH_2/9((W.Y^d22f@bC&IHR9RO\QU\FFTe,S\UG5OAX;_=GIA_+(W
dJQGH/XcO(be5[4Haf6IIMFe4Y,^(NBLXQ>/5J]4eNfAHCXe<B)GC2^E.TNR0D5+
LH.e1OFSH#YJH;&^&5XeV+DRg_26dGJaA9C]gg#WGJ\F)>1?Q=/:BVN&;M_ZH-b2
bWD5]9&=#(G>^(WgRT4?AP<(L=,9LN>A:QH&E[)8D=Y_K4E4>]bdJUL<C<VbGTDR
SVb&f/+C\Ta-CSH08-b-:@Z))&9>@V2\4]F&T<IfA,8JQHE.cABFTe,Nf-S)-La5
0&fR+>L(E7]\J]608c,NO,dM0-=d.<;&7fD8)P@I\PC9b#Z)^N.HO[H9^\QO_58R
PeDRA<XaMN8AbF=W?)9FI)3^R6O>JK]b(K1OEe8d3H\A>69V3_#\1<Q-(ZWWR;b>
1:4+Sc&S(#4QU:Q1V)#,8.EP)Q>Ee#K8WD[^IV#S:24U3T1R2VP<Q?=]49-PIe9E
8PS?c)MJ2@.8DJO:WK]WI54WgOe@.2GZ[B06@V?.Ke:SaJYX^d9<&cVIf.KCGO0O
@8U(E5(G1.\5a(1.F21(f=VY9T2]8^?(;ca1M87Z?>+BD,57\,2@J9D,AM-9_b2g
E]^c]M?YN&V]BXY_-V>G@Df>d^VAFCdKX<.,/L<T3^W=V].c)E.5VL0@F-:EA9,A
YO305c^SDFO]Fb:1YMdQ;;_;?gfMA@B3X/.5gT_^9;9>[AIJbC7RZd+W7KET0cNY
>D>DY@eA;2UcTQ-NKfMS<X2D<EPc)Nc>-_d4W77>.HMDf7E?5Y9C>I6O#=ACfK1Q
^KcP9AZ1;<gF3eY8Y0B-f0L/f+/&/NQO,14e#DD#VNTKcZ/HWGJF9(_,SSI;Z2P(
Vc:fS3c8:#<1\c=/d=-g\W64_0f<OIL.XG3EDKCE;IW[=f()@\3BPbY+,Q;V,2C;
/SV_4eIUJgP3?5&aMM8Fc]TJQO/=;U8_3IW/:7;7;O.\\A@RQ7^JIMRIc0^7DZR4
R8=)ZJ_TffFZNXQ<_OfE?B]+,^01L+_^G.W74LcRd8&I&fdgMafDF26\&VSa-gK(
1KAGGG?752/67cKgeIMcQbN8c5bG7M;4(TOG3JHNAN/MdX,,2Y>XcaIZL/K:X_Pa
.gg>Ic_c67W)>\BPDK?HHGR?62<MPIH_?WG9/BU__]aPIEd8/8N@U@1(\W^b,gXX
]6bG,<fc#/Q7R(fLYY3@,=Y?C7&/T::V(Kc#Q<IDN+aS(5b76#KfPCQ;E)Q8U2bB
)4ZSSgA7O#/UYC^1bN)&CeIXA=);H&CTNF(LJY9>IfQGO6KFda,(5&Hcd\IJ,?.e
-0X;.:#K\GX>+[;Ff_V;D6ADBO<2K.6[CE1/9X5g3R5,H9f[d=2HTa\+&51\3OS2
><54Cb@EU69E+97\C?S5-:DY4/SOeWN)X^+IJRZM:gN+1Q5#JON/JUfW0cWJNCF-
=HNZH85H&.W_gY(E,(GV=OO=(2GEFIQNe+OA_ORRF?,5@,94([/Y5ea0H6QgBfE6
dJ\.)4?#R-A6+F1a9U1La2)aK3CUeDOeLU\,^>eOaV6LQYLf^A(FUE=AHZB)D3c;
],_N;22H8F37(O-2J@U:.6GGF5\MIc?c/@OG7@W[GI]((+2Z;7))Z+K=/3S[AcLZ
]WQd,55b4<XE7^BbcDQ4CL7c)HJ=1NU?/#<-_,3Y[<P7A9eI3\LAD)T8V8[+T4;4
K)^8T/)E59AcL5H4\Ee^/]=3O-B-2-:Z?(?M3cKL8fg^A_QYgeLK0[\PYVaV_cL9
G4Q4@<6;&eec]IMd(EIQgSOW1c6AO6X]Y2_.ce/VVHB(g?-SFHaG6-+SK<O_dST-
/MDZcca#9^R^/=1AV>&FA=+44R;SB@?S[\DTX2<\@Q7]CJOY=Rf)(K,MJ.9^5;I0
L8]0f=G^JEH&6d?R)#Mf8<<OSb9^/ORL>N5_-a2]6[&F(]_+BXLR_ZSW)-KL#0H1
c8e<4a[^P:7]2e]^AH51=92dI6.VBV0aA9N>\BR_d)80&Z\<RV:6_N2a^7aFd;65
GL]cc(F]f&RY->SI+DfA^IN5H@0B.HSYP/8>2C>EH,6D.(?<F0;27)f^faGP@61A
5;9MMdDY<7/G)BZP7_+&8)AJA>:6EN#e-^=&X4SCA>9Y043ZAfH5)M<7[D&;TP.f
O9a-WXP#1^E-d2PE8<S#=97/-91071);VU[QEFN(]8+U3<fCd>ZHP_U?&<DQedBa
]XON@21MOAF[;FK;RE(+edT0REDMIA0TCZ1>^?,gG/1BcbKBK1Jg+6_gO#:FZ:_f
fY-4FCG@=]>;&5T4L<?>QJbLN?Re5/:31Ec?8>UC-D>KaAcZbO.O1-1UGg:\&e5U
M5]2dBJ73N@[c?HBB(3ff_:HG?0N9Q[QA2b(VOU8ANHb750@+J[LRW(W#e8)\RQO
Z\@&b9cJ>I2K3B\g#W\E1Ta_+=9[([8bWAJQN+cK3=K=]Ud3<O0EC2</]+<6Uc^3
2A[SL9HP8RC0<MD/EbJTO;[32Lf3g2:EF\S?#2+-4BWRCQ,X]6)L?>K(HS]F(,5(
WfM^15VeT\E50NO&I;R=-Sc</d5V&KFP.Q6EQSb4,/g)RO>f3(FC>MC@]D_K9&=>
ELZ@FA=4[#.0,T]50;aKOf#:RRU,_I@JAQ-XGAFZ-ZZMIKS61DDd7G+HQJMF9UOZ
I80NFec1+@]8Sd^&KX#LP<R(36L15#YaSC5B^&J6Q,IVN71WT\N9^1#R6P<5AN&b
V-&,P6U?:\1@3b.)WG@7Td36LR>#[Y-.&\)Y+_gK,@_]Ea?VDd&Z:20UNNf+9?&5
E1T.1;7W+IS]L#NAOLD(U?cBP31C7291GNOZZ_C=Q>&?AH=X^-O#.7KDL/J.7&1^
I\K#>9\;X3N2BD0_U4=81())C8^4^bEMZ4)eg1>8-XN+,4:K2Rb4#a>X7Of=7500
UI2gDVE+Z&-a<2ZZLG2J:31;H7202;_,[Y48^(baHCJd,V]-.1WcIdQf&]W>?2cb
C1?HT440/&>RecbC3W7D9gH@1gAGZSU4\fB>W0WD0R48COQad)#eT)5LZWXL(O:V
6+/&>G8I;<LPec)2f80We7#J[G3GfO@Dfda;=&RTS+K,BZAG/N1#c0@/DH1_(Lg9
T+4>]Vb,ERIcP+),:K3#dMgEL3/:N](E+RYRLCdZTR>]dL;M7Y>69[RdYMJVaV])
9(>7cE=\Q(U(37+:EZBfRe<ST#XY.EB(9HKg[A</KI2N?W/U:1]G8X,MB0?PX>A#
M03MBJ8?EdEZ>)4H[/+W&H^<(^YTK/dcXYR3@c4@I=WbFR)9\/D)9UZN:Eb((91;
c+DV&dC#^/?2UX>V9.T:PX(9/JT-#3:Q&^+QI/WUBG5&NUORPS40,6DRQZVb>g&8
-_YS@^&]5(&+C:ZP1Zb8e+2dc[/)37D0ISW<VQdJ>0;>))7D[Kf^0K.S)78SZI\R
:UP\L^)19U0B^-QDPJ(8+H.Ce&3FA;S6:.a:Hd[7ADLPQY[Y;E28YOJY&MN_C#bP
)C8B;+T6TYO>8(S\@;H<_[]Y6P8P0eQf]@//-[](gNCFT>[:FN./\c.)<_7]A.#Z
_Y:IL3=1&^.K1&+05&[PIS97C]43W@?=Pb1)EP1g9O#P;OSTgA?QaD&/:-=K(<4f
+4[_N:F@H1ZdFD,=OFE=fJDBbO>XbXIF^SF(f@>^9S<-]g5[:7#NfbI7/1.N-CYW
2e+C[<\=U]KLVE.S7SOg.85_bY?5W8dF6#)AL8a)TG1?<3Cc0N+FdBaLb[G^QAH7
]QM\0J?1[Ec1[]HAA#42gCC>GOObBM)-4N.EVW01B]W<^^;8]JQXcRC,FM,)Vf\T
8T_J&?=>]cV7SVN7UOB>]-7_+AWIebLdX_-Z/aV[Z58;,#^.fT6<9<GJ<2H+5^OP
I0H=U@F^0>XWU<(\TeCTP2?DI:CZ1#@&f9WGC[I&V8RD=&X;+@4?d99#@XF1RCa_
OS8D<0SL,R_DV:-UVX=#>O14b4g62gEPV5C:V80#XN#W1_fgd<0aE-I4EV-E#)4=
.68;50D_a[=D+D;b4YK_6?]6cSg^O^B>B5dW5Of/_7)2=-8M&>X7Z/I_84;5JJ[3
d\TV#5W(G\D42U3)J<1C^Q?fX_f#=bYc,7V8f>LO3g6OMd\,cG^>/0UNba;EaTVC
a:Z8Z:D)8f7RaW+fXd-2&eB8eI@X1/.f<\2X,=?5U_g/ZYO2/9AfF&UI:a0@V<#S
]J@S<C+EV@e/EY?5)T#3dG/_R),T]=WN&)f+^TX]Oe2TD,&\5:+K)[;,0&1MY/.(
ZJf_eCQ2>;?N7(_6:5HE2J(EKQ8IODNF4YP/c=[+EJYPfSJM:]SZZXJ=\0/3B<gT
&S\.#1?T=Q]](8Ed4EB[\eLWU1@3OIC8-fT4FaTFZ3&#VLMD?C<+f]ZMdHRQQ((N
I)/)TRU60)QF]SEg2U5NM)9J+],GU6PE=EbA=W/8]0&^b,][D<Y&<N\<;gf?;acH
8#&Pf-7g3[,5e+>f(XAN.>C54Q=7B?6.PRIEfg>FOYG&/4?bG&-C@>]/VEa54b;W
3_^6;6\1bRV:R.ec)#G.fbd3[eQ8WQX;=5DSg;,XB>AVS+?>ZC03GRC#^\Z4]4AY
a4T=]LSFJ2-DI.:IfGPD]S.3?+AUUbNAA7SK:f@G5Y:MC5Y2Z9+8[aa?UZPT:IV=
ACA)M@2L9dd4I2AGPHe=YT0+:I00Ug=6N[<Q[G0N]5&&\)0c?eSa8L:9gdM@_YUA
)QAST[?2YC+@U/J,dU5fUW2;g8gP0SFT2JZ#:X<Vf+cc9.M(gX7G)F^D10T&_MV&
>G-7#A^X=1G0)Bd/>[FG5^-##A^;7P.GG1<I5&)Y.f4F8A?b+a,8GZdf^>,H-&@<
J_)X-\2PgXMVCR^dHOcH_OdJ^bfW-7VY/QV7CAM+,a4PRP=8U2BdFVa8N/C/OVI,
f=3GDcOX6=R6]eO8aW.9<&3QAb6e//K(]c7[:O7MJ0#BJ]<U)PB;KeRCLV3?US&A
[9-+e6K(f,03+]Sg9C<@>2ReZ0(A++/]Z+5ALa8KggUF/Y+6\&+Ta6G@18eN,LO6
A>XX3R8EVg3\DW59\VF_E=C^?ND#g=^COB[f>g1]@31bNML@1O]:ec#C5;S;N\2)
5)EK7\#14?=ILdLK@7c+cXL]-,.GTWR3#A&.WHK>B8[;75Zb#d(+Z/)dYSH3PF61
X6/-;OCY3VI-()XU0Z?=bZCV3F6SLHXHd+7:GgDT=g4?@g>?Ib>VI(TMDV7Z+59@
@&+c7#3/YeFXUQ@UKP7=gQgA\1\D7g3Uc_3R/8J^b]:=e#_d?7Re7440\YQ4Fb[&
W4ZGA.fL#S_1Q;W+9AYU4/W9_JZe^:De#N>T@N>Q-9.;d;dfac]5<]SJA#6FF2EX
@T&U5Z6#-c_5GTeQId,E_/4A,ZIQU2RQDXI4.NS405\1&;1V?.56J5c367]>-KNd
F+7VAg^aEOFOCQKge?_9=Je<YG;JBT/#Z)C6;eG2AJFN85[XK)fE2LV@L6/EC/3=
eQ:-Cg6Z]Sd<F[IU.QcC[00\/[F.2PE3F^a?2[Z]P/_1SA]<PZdVb;Mg([_)N?IU
-a?EZ7)c@/MNg_T2;GGG&>7)IK2<8RI\1C#f/AE+#29L>41:MIQfH.+O#DO9Y;OC
;\DBTYCOM9EObH)&2Sc+WP8USSU;5gbP1W6A^c\_B.BABPb^b0+X8O<CI1:)gVD;
g8TUfcZ][8+>1FTa^EQ>VX/4LM8Bg0M8ga\8+_gH)^bQ6P.^f<);N)<8/;/#FKTS
/E]gR9V6YJF>R96LES,GWUW0CfTgeI,<#_/Ng;[MQePC@RO-&+C>3YGJbeFA^T,7
XCO.0C.:,[V5P?.JbXPN2XP0B#M#Yd#_N9CMaKc#4\>W6Ue)8dGdG\L,J3\BBF&2
3?T]ZOI-=TE,WcbOUF:.?Q.0Q:Eb]g_HW<U0Kc77V47VZgJCfeI=H1BS&d0#R_dX
^_M2KdHT8H:HH#D/6/f3F&B<RZae.W5R9)#fQ#I2:#R&300U1P1STRQOCTRg8QW>
aJX8TFJ9<F8]WMd_&VZFTe,48#=Q\3YZ-/V/aLT[HaJU^J=KL0:QUKVLK/:N-Ve-
IcR;N+f9<-LV96b?b18QQ/M87ea1^<&gVdNaA]S]P:-_Q-K:X@/6L,-<U(#>:3K4
;V5X[(.FXF.WS[I99_\^;XfdJ#L9N/74VAOR2ALN?>\+)b-b1&;GJA07RW_/H7,G
8_(L1@Od@B]<G3-(\#SQP>EBJU/cR,9g4gf74JQ3fF?8EB9A3g/)@A[)-WA.\T.c
H[eH?MgZ2fF8Ic1JM_[f:MS(ad/TaFdJ9];dE\3ETaS9O;BE3d&MF8N7./)T)XZ\
FLS.1XW;NR^<&]:@^/+-RX:7Z.Y]CA446eRf\([@UWfG?Gf6XCcAG>:e<^fH&/6f
=/2\(Bf.FdN,>J9NTS3#.3/Q9P7(:b5W-Y21/b(AE1H_L58>OdL=3/a:62@^0Y5H
V.MW9D0fbOA,.$
`endprotected


`endif
