
`ifndef GUARD_SVT_APB_SLAVE_CALLBACK_SV
`define GUARD_SVT_APB_SLAVE_CALLBACK_SV

/**
  *  Slave callback class contains the callback methods called by the slave component.
  */
`ifdef SVT_VMM_TECHNOLOGY
class svt_apb_slave_callback extends svt_xactor_callbacks;
`else
class svt_apb_slave_callback extends svt_callback;
`endif

  //----------------------------------------------------------------------------
  /** CONSTUCTOR: Create a new callback instance */
`ifdef SVT_VMM_TECHNOLOGY
  extern function new();
`else
  extern function new(string name = "svt_apb_slave_callback");
`endif

//vcs_vip_protect
`protected
VcHdNQW:7@96>8b\bfRa(2MIF<HWd?\1>_>.dcWe2#3Q[3D<6=\Y0(/@9J-&1C6N
.,;K@Q@<1gFPbEEcff=_3@aZ[Ig,K,3MMB)KLU&V]02@9S=W-S7e>?]@L]\5R6)(
))\Ac?\Adc?6Xd3+Bg&ZZG7B_\/065OH1YGYA:,f.?1[,.;)GALP>&;cLbC[>#cT
HLQ8EgJ9>K31LB38B/>-@d7WEg:e@DEDA]@/\IUKKXadaTATB,dBaPH?VFZ>6cK&
W,\g6?UMa^FeJ3VC)39<V1NaW&8+3PF6Z^dPM8^]H6da]/.6T&F-21BYO:[YRMGa
gOa:5=7_&5535(8d6<E)d_\d#E^b18CD8VVAE9>PT\P#;cOeAD/:RX/+;<BU2S?V
UX87?63CRZ+:e3A1\3>Ob5^WB(7ZY:Df?U2@13a#QPR?d<[9aS]A.3(9E8_D@;68
H@+:D4RJ;HGJg>>I]SW;33B:;/VB,c5K@3OC0F4D;+B#4@:dSSd?OgI5V,HZ)W2F
7BSY#=;Abd67SS9B?C;2UK:M<0BA+G[Xb0geAW(GZKQK5ZO/]2cKA^RJ\9+S/@0N
4:90efHTRca@UO^a?^7>-#3edPZB&2:ZE-OYGP62NKQ2a]A3J+5[M=7&\V8J2G&T
]NHLZ6Bg4cJUF0+P6VE47aW+X:=?(U.W39fB/dN3:]G.>Ld/597HgZ[;LPbB(cd\
:US0:(VG^dGR:PN5KAMgS\1&5V..d,[E)X[WgE-H4,,;?&4(Yd\=VGWcUd(IN^)F
aE/6gfgH2SK>KZb[_1_#H:OYXHGGO+-;:6_JN7J5_bUOK0BJT6HWC>f.J;LdC@:&
>U2;62.1L5=T=V3=4eJV>f&=XKXDK03C5FS?]P7<g,G:S@J?[CCMK+DVQMS0TI)J
Ea4>WL8-.<b2OA_J6Q/aQ?19EAYPA2_-K4DDXcG<34O7\Q]C9PBSbf5,L2MZA&:7
gV^;2W&;gT,X3/GT40G,CM;7;0H<Hd1d&L<,NRWQgP2aM^^L7-_OHID_<Qf7-_L-
0aP<CX8,\EP,H<_2.D5DNKd7>E?6O@DO9A(/<?a6&\=gXC8+C2-B/[LDV2&>Y+5@
8]5M],_8Ge(ZUN,4KP0A+L1ELf4-?3+K[&TNa:M4N]Y04^N6Qddb4DXM__#M9d5B
,4XF7#a9Df]g2gJ2XcW:J5f.,Re:2f:J)XH^)fG&=.9PfB^;U4CQFcH++&<Le8=L
CG=Gb3B#QN&+#GbU_FD?_EXb9#^>e?K5Y&V1(e\Z\EKDKNQ]eNgBC0VR8X-5V(f3
;J=#@L/L;8Yc,JZK^.:C@8<M[eDD4Q:=Ye,MKCI1.X7111ZF_,(aG/2.Pg\.42VC
.3>9bI9I8S/Yg=1K+UATTcM2YP>a7]MW4XC,,OY)1UR3fgM-=2;#2?Z0[KM[E#>/
=ZCaM?N2-#P&U<RPe6dQ8O)O6E>HXAQ^,f#4:[=JL0>Dcd;TdIE/[LOR_&.3YaNK
F9S#b/5Z;I7a,@43Z8Tg\33[Z]/#_,F>XF;L06QMG;N>C+00g=3NM7fdO4P<P0,?
D@)#.IC/6QU3Y+a6IW6=F<.LSUDdU38G3&c-VCd2,eR5LcD]J(SRE0ZYeJSNSZ&M
V6ggJf1DJe:]S-9&W;H?[OXad7Xg=DG[N</?HHZC.UQQ&N&:AO<gRZU1#Mda4]dR
@ZPN7;)dV0Z#]?)Qb7EFQ[?P69#C;7E+a(3;dOJ953eS+04Ne_KQ>O5IZQA6.-c&
RC55WSQ)cF4(f=(A#@?W6+F#Xa7^NMXT6)/37[5S3-5?e22Rc?BHdIg>B<B[6=E/
N?4QZMOT0_e1Tf(8RGJW2?a><VG_+_^bF[=#1CW]T:987MFe=>@U>BZFP,eKXN5W
;ea+Q31]>XY\7NPUb@NHGHV7R\M^fJ>&1J)Wa(=I+VD9?Z7XPO_e@g?Z?bA02H)(
K5O;C5^@W];<V]7I_?.K@+5--X,G.CU02\]GW1Mc=D5-5fVf-#O,[]T,dMeS7HNF
^LDF[M]VIQ4)Vf2&U4(ZL0c=W<\0)7bJ<64Nc@V\<8RPSCUgOb(c+-T,J$
`endprotected
  

endclass

`protected
/I&YZ<e>Z-@8C#RfM\IaO+MA,b,9d@Y?>X;CNYVP/@F_+a8B>>G<6)a@+MVa+FXE
TX(70U/(PdMOXcOd9fQ#a>c2H#0(e_Y&Q/W#1gPD=KH-_7.0cE0T(O#Q3SW5F&VN
>U#NNU-JHf1/4U,eH8VWKb07-Z8d1Z,<EdBU?#D<KIH\OC#FB\1F1EPE?G.H=^gf
9E]g:[>2NC)(U(:U9W<dO./A+ZeG)>#<3M@edAb)JYWB.c,L?MT(a<CYHBN]1=2E
Qg4UJ8IdP4]cANcV:QGNSO9^0P<#P@F.?<W#B;GD2_,:I,0:Q:PAUY]KMgaBH2B<
RR:)^8KfMW:N(I\,_WFc(B6Ff6UNXA9Y=$
`endprotected


`endif // GUARD_SVT_APB_SLAVE_CALLBACK_SV
