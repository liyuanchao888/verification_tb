
`ifndef GUARD_SVT_AXI_SYSTEM_ENV_SV
`define GUARD_SVT_AXI_SYSTEM_ENV_SV

// =============================================================================
/**
 * This class is the System ENV class which contains all of the elements of an
 * AXI System. The AXI System ENV encapsulates the master agents, slave agents,
 * system sequencer, Interconnect Env, low power master agents and the system 
 * configuration. 
 * 
 * The number of master, low power master and slave agents is configured based 
 * on the system configuration provided by the user. In the build phase, the 
 * System ENV builds the master, low power master and slave agents. After the 
 * master, low power master & slave agents are built, the System ENV configures 
 * the master & slave agents using the port configuration information available 
 * in the system configuration.
 *
 * The user can specify whether Interconnect Env is required in the System Env,
 * using the system configuration. If Interconnect Env is enabled using system
 * configuration, the System Env builds the Interconnect Env component in the
 * build phase. After the Interconnect Env is built, the System Env configures
 * the Interconnect Env using the interconnect configuration information
 * available in the system configuration.
 */

class svt_axi_system_env extends svt_env;

  // ***************************************************************************
  // Type Definitions
  // ***************************************************************************
  typedef virtual svt_axi_if svt_axi_vif;

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** AXI System virtual interface */
  svt_axi_vif vif;

  /* AXI Master components */
  svt_axi_master_agent master[$];

  /* AXI low power master agents */
  svt_axi_lp_master_agent lp_master[$];

  /* AXI Slave components */
  `_SVT_AXI_INTNL_SLV_AGNT slave[$];


  /* AXI Interconnect component */
  svt_axi_interconnect_env `SVT_AMBA_USE_INTERCONNECT_INST_NAME ;

  /* AXI System sequencer is a virtual sequencer with references to each master
   * and slave sequencers in the system.
   */
  svt_axi_system_sequencer sequencer;

  /** AXI System Level Monitor */
  svt_axi_system_monitor system_monitor;

  /** AXI System Level Checker whose checks are called from system_monitor */
  svt_axi_system_checker system_checker;

  /** AXI System Level Transaction Coverage Callback */
  svt_axi_system_monitor_def_cov_callback sys_mon_trans_cov_cb;

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
/** @cond PRIVATE */

  /** Configuration object copy to be used in set/get operations. */
  protected svt_axi_system_configuration cfg_snapshot;

  /** Fifo into which transactions from master to IC are put when system checker is enabled */ 
`ifdef SVT_UVM_TECHNOLOGY
  uvm_tlm_fifo#(svt_axi_transaction)  axi_mstr_to_ic_transaction_fifo;
`elsif SVT_OVM_TECHNOLOGY
  tlm_fifo#(svt_axi_transaction)  axi_mstr_to_ic_transaction_fifo;
`endif

  /**
   * Fifo into which transactions from master to IC are put. These transactions are sampled 
   * from the scheduler output of the interconnect
   */ 
`ifdef SVT_UVM_TECHNOLOGY
  uvm_tlm_fifo#(svt_axi_transaction)  axi_mstr_to_ic_scheduler_transaction_fifo;
`elsif SVT_OVM_TECHNOLOGY
  tlm_fifo#(svt_axi_transaction)  axi_mstr_to_ic_scheduler_transaction_fifo;
`endif

  /** Fifo into which transactions from master to IC are put which AMBA system checker consumes */ 
`ifdef SVT_UVM_TECHNOLOGY
  uvm_tlm_fifo#(svt_axi_transaction)  amba_axi_mstr_to_ic_transaction_fifo;
`elsif SVT_OVM_TECHNOLOGY
  tlm_fifo#(svt_axi_transaction)  amba_axi_mstr_to_ic_transaction_fifo;
`endif

  /** Fifo into which transactions from IC to slave are put when system checker is enabled */ 
`ifdef SVT_UVM_TECHNOLOGY
  uvm_tlm_fifo#(svt_axi_transaction)  axi_ic_to_slv_transaction_fifo;
`elsif SVT_OVM_TECHNOLOGY
  tlm_fifo#(svt_axi_transaction)  axi_ic_to_slv_transaction_fifo;
`endif

  /** 
   * Fifo into which transactions from IC to slave are put when system checker is enabled 
   * These transactions are sampled from the scheduler output of the interconnect
   */ 
`ifdef SVT_UVM_TECHNOLOGY
  uvm_tlm_fifo#(svt_axi_transaction)  axi_ic_to_slv_scheduler_transaction_fifo;
`elsif SVT_OVM_TECHNOLOGY
  tlm_fifo#(svt_axi_transaction)  axi_ic_to_slv_scheduler_transaction_fifo;
`endif

  /** Fifo into which transactions from IC to slave are put which AMBA system checker consumes */ 
`ifdef SVT_UVM_TECHNOLOGY
  uvm_tlm_fifo#(svt_axi_transaction)  amba_axi_ic_to_slv_transaction_fifo;
`elsif SVT_OVM_TECHNOLOGY
  tlm_fifo#(svt_axi_transaction)  amba_axi_ic_to_slv_transaction_fifo;
`endif

  /** Fifo into which snoop transactions are put when system checker is enabled */ 
`ifdef SVT_UVM_TECHNOLOGY
  uvm_tlm_fifo#(svt_axi_snoop_transaction)  axi_snoop_transaction_fifo;
`elsif SVT_OVM_TECHNOLOGY
  tlm_fifo#(svt_axi_snoop_transaction)  axi_snoop_transaction_fifo;
`endif

`ifndef SVT_AXI_MULTI_SIM_OVERLAP_ADDR_ISSUE
  /** 
    * Fifo into which transactions from active masters are put when 
    * overlap_addr_access_control_enable is set in the configuration 
    */ 
`ifdef SVT_UVM_TECHNOLOGY
  uvm_tlm_fifo#(`SVT_AXI_MASTER_TRANSACTION_TYPE)  axi_overlap_addr_access_control_fifo;
`elsif SVT_OVM_TECHNOLOGY
  tlm_fifo#(`SVT_AXI_MASTER_TRANSACTION_TYPE)  axi_overlap_addr_access_control_fifo;
`endif

  /**
   * Port through which transactions in master just after getting from input
   * port are received. These are used to decide if the transaction needs to 
   * be suspended because an earlier transaction addresses an overlapping address
   */
`ifdef SVT_UVM_TECHNOLOGY
  uvm_blocking_get_port#(`SVT_AXI_MASTER_TRANSACTION_TYPE) post_master_input_port_get_port;
`else
  ovm_blocking_get_port#(`SVT_AXI_MASTER_TRANSACTION_TYPE) post_master_input_port_get_port;
`endif

`ifndef __SVDOC__
  /** Common file for routines to control access to overlapping addresses */
  svt_axi_system_common system_common;
`endif
`endif

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /* External AXI Master components */
  local svt_axi_master_agent external_master_agent[int];

  /* External AXI Slave components */
  local `_SVT_AXI_INTNL_SLV_AGNT external_slave_agent[int];

  /* External AXI Master component Port Configuraiton */
  local svt_axi_port_configuration external_master_agent_cfg[int];

  /* External AXI Slave component Port Configuraiton */
  local svt_axi_port_configuration external_slave_agent_cfg[int];

  /** Configuration object for this ENV. */
  local svt_axi_system_configuration cfg;

  /** Indicates if AMBA level system monitor is enabled */
  local bit is_amba_system_monitor_enabled = 0;

  /** Address mapper for the AXI system */
  local svt_mem_address_mapper mem_addr_mapper;

  /** MEM System Backdoor class which provides a system level view of the memory map */
  local svt_axi_mem_system_backdoor mem_system_backdoor;

  /** MEM System Backdoor class which provides the global view of the memory map */
  local svt_axi_mem_system_backdoor global_mem_system_backdoor;

 /** Arrays to store the information regarding system interleaving */ 
  local int num_ports_per_interleaving_group[int];
  local int lowest_position_of_addr_bits[*];
  local int number_of_addr_bits_for_port_interleaving[*];
  local int lowest_port_id_per_interleaving_group[*];
  local int system_sema_id_for_interleaving_group_id[*];
  local semaphore system_sema_for_port_interleaving[];
  local semaphore system_active_xact_queue_sema;

  /** Queue for transactions from all masters with port
    * interleaving enabled
    */
  local `SVT_AXI_MASTER_TRANSACTION_TYPE system_active_xact_queue[$];


/** @endcond */


  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************

  `svt_xvm_component_utils(svt_axi_system_env)

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * CONSTRUCTOR: Create a new ENV instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function new (string name = "svt_axi_system_env", uvm_component parent = null);
`elsif SVT_OVM_TECHNOLOGY
  extern function new (string name = "svt_axi_system_env", ovm_component parent = null);
`endif

  /** Obtains the System Memory Manager system backdoor class for this AXI system */
  extern function svt_axi_mem_system_backdoor get_mem_system_backdoor();

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the sub-agent components.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void build();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Connect Phase
   * Connects the virtual sequencer to the sub-sequencers
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void connect_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void connect();
`endif

  // ---------------------------------------------------------------------------
  /**
   * End of Elaboration  Phase
   * Checks validity of System Configuration
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void end_of_elaboration_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void end_of_elaboration();
`endif
  // ---------------------------------------------------------------------------
`ifndef SVT_AXI_MULTI_SIM_OVERLAP_ADDR_ISSUE
  /**
   * Run Phase
   * Controls access to overlapping addresses from multiple masters 
   * based on configuration overlap_addr_access_control_enable in 
   * svt_axi_system_configuration
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern task run();
`endif

  /**
    * Extract Phase
    * This phase is used to extract simulation results
    */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void extract_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void extract();
`endif
`endif

  /**
    * Report Phase
    * Reports performance statistics
    */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void report_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void report();
`endif

  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  /**
   * Updates the ENV configuration with data from the supplied object.
   * This method always results in a call to reconfigure() for contained components.
   */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** @cond PRIVATE */
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  /**
    * Updates the agent configuration with cfg object supplied from agent
    * command component
    */
  extern protected function void vlog_cmd_set_cfg(svt_axi_system_configuration cfg);

`ifndef SVT_AXI_MULTI_SIM_OVERLAP_ADDR_ISSUE
  /**
    * Gets transactions from post_master_input_port_get_port and tracks transactions
    * to addresses that overlap with previous transactions. 
    */
  extern task track_overlapping_address_xacts();

  /**
   * Returns the requester name for the supplied master transaction
   * 
   * @param xact Transaction for which to return the requester ID
   * @return The component name that generated the request
   */
  extern function string get_master_xact_requester_name(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);
`endif
  /** @endcond */

  /**
    * Enables AXI System Env class svt_axi_system_env to use external master
    * agent which is already created outside svt_axi_system_env.  User needs to
    * provide external master agent handle and its corresponding master index
    * number. It is important that user creates System Configuration including
    * the port configuration which is supposed to be used by the external
    * master agent.
    * 
    * If system env doesn't find any external master agent for a specific index
    * then it creates one on its own. So, it is important for user to set system
    * configuration with correct number of master agents considering external
    * master agents and set specific master index for which external agent needs
    * to be used. It is allowed to instantiate some master agents within the
    * svt_axi_system_env, and some master agents externally. User needs to take
    * care of correctly specifying the indices of external master agents to this
    * method.
    *
    * @param index Index of the master agent which is external to the AXI System Env
    *
    * @param mstr Handle of the master agent which is external to the AXI System Env
    *
    * @param mstr_cfg This parameter is not yet supported.
    *
    * Example:  for(int i=0; i<5; i++) axi_system_env.set_external_master_agent(i,ace_master_agent[i]);
    *
    */
  extern function void set_external_master_agent(int index, svt_axi_master_agent mstr, svt_axi_port_configuration mstr_cfg=null);

  /**
    * Enables AXI System Env class svt_axi_system_env to use external slave
    * agent which is already created outside svt_axi_system_env.  User needs to
    * provide external slave agent handle and its corresponding slave index
    * number. It is important that user creates System Configuration including
    * the port configuration which is supposed to be used by the external
    * slave agent.
    * 
    * If system env doesn't find any external slave agent for a specific index
    * then it creates one on its own. So, it is important for user to set system
    * configuration with correct number of slave agents considering external
    * slave agents and set specific slave index for which external agent needs
    * to be used. It is allowed to instantiate some slave agents within the
    * svt_axi_system_env, and some slave agents externally. User needs to take
    * care of correctly specifying the indices of external slave agents to this
    * method.
    *
    * @param index Index of the slave agent which is external to the AXI System Env
    *
    * @param slv Handle of the slave agent which is external to the AXI System Env
    *
    * @param slv_cfg This parameter is not yet supported.
    *
    * Example:  for(int i=0; i<5; i++) axi_system_env.set_external_slave_agent(i,ace_slave_agent[i]);
    */
  extern function void set_external_slave_agent(int index, `_SVT_AXI_INTNL_SLV_AGNT slv, svt_axi_port_configuration slv_cfg=null);

  /** @cond PRIVATE */
  extern function void set_external_master_agent_array(svt_axi_master_agent mstr[int], svt_axi_port_configuration mstr_cfg[int]);
  extern function void set_external_slave_agent_array(`_SVT_AXI_INTNL_SLV_AGNT slv[int], svt_axi_port_configuration slv_cfg[int]);

  /** @endcond */

  /** Obtains the Global System Memory Manager system backdoor class for this AXI system */
  extern function svt_axi_mem_system_backdoor get_global_mem_system_backdoor();

/** @cond PRIVATE */
  /**
   * Obtain the address mapper for the AXI System
   */
  extern function svt_mem_address_mapper get_mem_address_mapper();

  /**
    * Adds memory update transactions to system queue
    */
  extern task add_memory_update_xact_to_system_queue(`SVT_AXI_MASTER_TRANSACTION_TYPE master_xact);

  /**
    * Tracks active transactions. When transaction ends, it is 
    * removed from system queue
    */
  extern task track_active_xact(`SVT_AXI_MASTER_TRANSACTION_TYPE master_xact);

  /**
    * Gets the memory update transactions from the interleaved group id
    * of the transaction given in master_xact
    */
  extern task get_active_memory_update_xacts_in_interleaving_group(`SVT_AXI_MASTER_TRANSACTION_TYPE master_xact, output `SVT_AXI_MASTER_TRANSACTION_TYPE memory_update_xacts[$]);

  /** Gets system semaphore for interleaved group id corresponding to xact */
  extern task get_system_sema_for_interleaved_port(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Gets system semaphore based on try_get for interleaved group id corresponding to xact */
  extern task try_get_system_sema_for_interleaved_port(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Puts system semaphore based for interleaved group id corresponding to xact */
  extern task put_system_sema_for_interleaved_port(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

/** @endcond */
endclass

`protected
AZ1/bY@P[KD:,XHH/<S?I2:Z[PH^H_a9UPS)3Q@DPTc[TU]>c3eM6)+HV.>3^DID
\5.IB,PKd;CX<[X&[;2;ZY_#4POM^626CED4/&L.Y.-b<ebKT\=XAM.\6TF4RMN\
6?NeD,N+K2\GTgNC-f)6&(;Oc@;A]X,D/]MGI<C=47#N.SXTE;2>Ye+XQII1?>b.
.c65c2DM7)V:EB#g?>d(DG7R#\T=DYQe+:JUZC+T\6d?\--:e:#Z.]W5U@S>Y,,#
6@ZL<S:>42MPeY=SB=)P1F;-(H07K:_>C6TQ@8E?AV](Xa>2_DM&FUOTD&L<,K(&
aNRNV.b>=?g+^We,6[TZ>+PL,gKC4=)C-8PTcN]XX=90bKg]DX;BDe4FGc/Id=&B
1?d1]G8;PV4B+bIZcbR_[+NO5.8=ZHY2/3R5@=)c>)GQ<f9P?CLcDN)IN+P<L]J3
<RITVd<(3]2HP.d[UG\-+ZB\^a]0<d\-->.C]gJ[@T[aJ9NE;=Bf5FEZ<=?_WZKe
,FWV-&^&_2.H/$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
:<4YO5(9KfLGW>9_<Zf?^X,RV3@e:4g(?T-=Z^J^H;P6EXb176US3(G^SC8[PY)#
&Pg05EJb)d@W?L<U?f(gH-eXYc38_@U8COS6&&CQ(V2W&a]7ea0.JAP](@Kd+=c#
?=a3Ve3[O352gK8a76<.5SR4,=BI3VMa:Z^#eN[18@KcMFXQ[I-)Bee1fA2K]Q^Q
fa4E:ZH:G1cH(.VRVKD/38Yg6;::S+e51GOc]GG0cI;4-O8K6[G+37(A0FI(5ZL]
fgZ=4G9,[M<+HJEc4W)1T27TEZJ-<25M;4.fB+QVYR_0[.8;+TP0/20Q)?(-MJ=G
W/7(W].KCe1#2H]bJ8->B1d+<IMO70:PTJBRCOND3ZbG((\+]^43W2HZa?3<Ab<D
@I7/,7:./7ER;[=[0I24<_:GgZ]04\+OM?d6.FX4fZ5AO@M6.IJ@YIg8gg[?+FUL
1dR7Y.Y2NR&^H=ZSg/#1TKfLD)Od].7[a)_d0NY3QWe:[KJNNA#C4KJbdTK@GA<<
&MeD>LODLBOD)+A2[,@IG0fL^EEC.8gY#I[M5I0CdgRWSUc5U)g:?W.LV)HKKVAZ
PRcD;UQ1UbM(=E_<AK>L=ZJQa5LM^^dL2a.H6<JLd7U,HS8X^+&(IG7<Z8c&a#+B
T&C7C5EeA3VF?;bfFPcQ5VHbMOb.]@U)1\Ne3XL<6VW7+W_\SdB>cN\B=)-M6S_Y
SfeZHF32>/^XKNBM81H37O.>+H,2.7AeR27]JS3UXFZ_+3a(CPbJ-.[fMfZQ5#Uf
QGXe33#K_gYH:[Y(?JK/Y#HRJ#G2HJ])JZ&(5QeTC>5G:X-FGK[/P\P+M:1/,.;1
V,R7_DLYM()V_]fV(A#B@>c8e@+.Dee=YH(NE\;@^>(1^2_2RHB2,7A6KUI2#2()
(S^0WVe<H;,@C-d)YC.^5F\@CfC5Mf<L6fD>AT?[.7^cAgfg+f<fXA/)M^B5=.cI
TMK^4?1dCaV++eNTIDdSZE[-VOT:SV=J[3?b1D(#g<:]#b2MNBUg6=I0B7GN0XL:
O5,S5[^-I@EBVG>+AE^W&6?.6,cN30/G?]ad;.a+cgEe+[_KLQ,NcT@XJH.;XY;b
3?_0FAa7+9==^\4F(8F&R0P>N#RJ_b,Qge8XMTZDL9D4NCH&22dY4V9=I#OB(cC[
fNYCNE)8O0)S2ZR9;e;[)c,;3g_,A.e4_1#Z[+D3Rf^[gRa<N\:XYB<ZGbYaMK_>
a&=bKM8.&YK0#Ad2G]@VbU++LWg,ULUE:(--g735d&45IG7^5a3^_G/8<5f^gcZ2
?HHd.F4eH6.\&4Z)PZ.;58MXcK:4X\RO029?T&8\78)QW((RYIbS0&DEB34ZK^W@
U+fdK>RJd0LW7<W9g7e=BTJ6^)b>Y]gB+HHUYX4=OBHE1bKU7b\AdFE&+\/(]HY8
NNI\aE?:5O/gF/L[5ECV+d/QJ0QW.KPFSXE\5TJ<eOKJW.^RQU:XN7@-:0P.VXU)
#2R=1.8bBK&a02cX;9_Q_SQ<H<aZZ9Df0Fa)X8M7-/>FZMRV;EA3IGQgY#,=Hg#T
f5EeY-4&=3UY<(X^EM^dc#IK-H\B.EJYP@QN0^Lf2\5/)WFSJa[G@,NTA>^4G.M?
6UXM0<=Q,8#9a#Y-2\79ff]?cZM\Q0#f?EFQa+a#EGf/(RAc+=:W\JI&X^c3\+,J
U6)623#1Ogf85=B;d15&;0VK@HfJMU4NR=JP7d^ZP+1,V2#739cb.]:,RReH8KX2
YBe4JWB.?J0d0<5]Jc_)Uf[H9,VPM])(41(VNcXO&U3XDBN?KR)BNC\#=LBP<C:=
BL@-<e#?R#E>M.eQ_JLY&<1b-P5HadX^W:GK>cG?-B(IYe>-B-BeKURb@EE1ON]_
-@2X136UVFI/0.V;3F4dJQ>LPU-/+H)YB+[^Ea^[39=42:bR4C5]=eX(1/=[.31F
W]2@44JGS\BP2,KQDE.Ha_W_T#0YNMAg65TGcYIb\MISgd[]]cTACZC,O62M9OE-
Xe.SB@feV]/_1==EJNR&[&Fc)]b<;gJH=.AXg+JJE&J]:dU/GaS#/IeO>^WV]C#e
\BK?MVK[_c2.WFU1N<JW8UDX&M0?T1IfFe)1/<B(=4I3;];a9C=3BAAeV,XF[EB+
Se^;3K&P1.S4P?=2X=.[@GSdTH,C#]DW-N;LK8c[fK;IVALUPQL[,[47L/01\aZ(
DBV)g#_?I67&Z<#@I?I0Fe8O^/Af>eIdcOL=(g57(>d?Q,A+(+S@cbdN2cMKG2K^
,3>AVD-eEHg1ZcM]J>Y=?/9AW8c@SI8Z_^ge\g]U[(<?7e3Fg:BIU+@WB,[+J.41
B#/CeW](7eSMd&=E2=_N:GPg@2XFB4DeP/G@2BB629LJQK:\F3D^Bd8^(&QYSg7#
5-]+bGfE9T_2[,-<Gf75LVF[/DM>[T,ED9eUQLMg6OMUM.LBg)Q@A3&J8bLAC)5(
A#AB13AgQeKMARceXgf@=aTT1Q,.G=Kd1f=g-G2Wa]Q=b61b]?;C[UA,f=R>:CEQ
V@Z/-B<U-1V2]/b5L,RL7MN&4.U4K^Z-3KR,/PTP[SXV:/?#^=9V=NIX?(-I19];
=SYRIO=>O^5#C,)>&-/NcQ122=>E,A6fSW-8&a)0E:FMT>dJIe8Pf>+00ST+^M#>
K&K^HB21+-9=64D..8W(B@G,5FFBcXdKOf8F<S&^8D\=_\^TM.M?YB]b6_?0JV2X
WGEGK0#Ue.X1e-D0G[5DITedcbIAH[L\8b?+daC8gDcHP),>W_?a[Df2\_\21BL>
-::gQ3H]3<^<7XP8&=g(E=H/KPQ<a>?LI>/<]Ua4Q>R]c2-BD<VJ24\Z\]]g@HWY
>LEgND+g\&Q9dJDa8<&2:]0=B@,fDPPV5@?_FbN6:]0]N/5f]4L\@9:(g0O?8:<@
</@[X?R]03NZVEO&:Q]H7G9+3L)Bg_<,Y_05@+AW<(CIG;E.&+(aV&7]GQ=T86B=
2K0)Y,I[:)ZM.JE)FHC]-cP/DS]f.?#QRNad[0Jd&\PI]>&+>fY-&,+C3b=<#WT<
=4eR;WeM+^d-ZD49O+\caMDHP#4C[N:>f,b=fbS3IW2<S8aS_#N-I1gfA6V4-dAg
ZI7:7RTFN>_4))Y3[NF=Y]R#g3#X)?M8@.IX[.C97GfA:<DfVSCL6ZHg^70A)5XB
<@(34bHV9MW:FP.f9f1c#@:dVe9;22]>(4Rf9H6JR(Kg&;bS16XSX)BR:\2+?OUL
_SNcU]SfU@#NJH7RH[K)aCB51fRCS1^#W4Z[?)K+W]16[3#=U<b]9)BES1b(V1OO
MZ/&Z]#.C1LXP=XHb2R3TH/;8L5aZ6?JT6/T]UO6,[P:0IR50Ad-cDY-9KfFFZWL
7aXCVBD<C2E,ED]1K02#>-L)[>=bJ+dH9OdJ,1KT)YT9E[C14b6Na#<K65G+\B\R
A=.IYY=R[CUS1Qd;9G.D?7K#_I&ODEO>-f=6K6NW[c-R.GE@aMV:V04\M,=1MU6K
^X;,-ZEA4a4L2]H:UA\Rb/ENYZB8D+e_<<_06UO+@Y&+BIGa\??,.GE@.F]VRPYH
7EI-Rd1c)LbLPZGd8HU?7fA85LXQ3.#fA,0\G9N0a_3._ad4CJ/N)F9d^f0\?\;[
6TY?b14O>9X;0)Ad^XfK6G?aX9()]Eb-9:[QF,8W/K@:XM0C>YBRD\.-WBI]4(JZ
B>S_fe7gZ17J_BU,Wb(7/KJ]LaL/QYM39X+1.?=X-=]O#Q462&.>1I?PUe?<NI^4
AUW^3DgYO65fG[Z<)PXAM7Db6C74&97T.FU(1,M21c.G8SW=)N?dRg2@)OA\]0_G
c>],G5Jb(AMa-,^&IM@PPdZ((ba4,9^BLdC242N^GCR+VQ5_X[2dRgb\Z7P1+cf]
.OF::7K:eQ]C73<BYE?J@eLPF7LJ@HU_.VT[&6:-F9.A+,2+7@]IQK<83DY1I1?F
_P2bX0G5&/5A>OeC-L.E[?f3EB?=ZM2WaY^cNL0GAPL:<>^O-P5WJ@YL]/,J2-QB
D_FcFC275BDV#@:/W#UQ<9H&\)&1[fP.&WN3-7X;X/GH#)46;b9=(#MQ4<b#f=2B
S:7c^,.F./b8<AKD[c0CE&.S]0S&Q,9e<CQ#Y/9aMKb6:2B8@b/\,LRE8cB+_^0:
X(Qd&PQ7.2TL9aN##)22WC?)+T9J&b_V\.)49U/VLVdf-4c8:Bd-#2C;\cLAXbE9
.6GDb;3g3.MZE9/#=Z&Y8UVJ#HN=\;YIF2QH4_@Za.PE>K;,gDF_R3@)Gc<T@W?.
7I1fE1C;;88BROI)FXGe0-83?L1_.L.;a9d.b9V(\&GTCFcO>/-R<W[W.2X3>Q=+
c;Q27eYS@50P)U1==O)DH=IP][(?Z\L\G-ATbG44E]fgaHJ_Y(-Z=,)4)N,;N-UE
J3P:[-MVc(T.JR;>Ag)4)\]Cg2R+a./;634Z(Y.We;0KeY2R5_&F7A<bG#e^18(X
^\)Y4I>J;5#@c>5bAM-NYES61a/P\\H>L5?U<:g46c#DMPBGK\EEY\&f]R]<^@<9
W-SK:,&Z@c)I3HCS#C_J2e>A6Yf+YN.c54TFgZ?Q[\8@Y7c;40FgH>+R;-7N2\L\
GXSIc?7<\b+YWWg+/4EL\#H&=G@D2=KR^EY;Z#P)V2C2&6M:VgN_)7;8PESFf<=L
f_LW3]S>-^S/B:7KSLDM<UW-GX?PdfCN--5gg2g-A4bO&PJL+OV-HTNXa8TTPC0M
b]cRO[>:Q8J>>PU[(/:HTZ53d&c#/Za?YS06c_QSC?.Q=&9]LNVU6R?U-6HA[De/
bOJ56Z@73c3SX,eQ.Q&&7U\\@QMS^@Y99Z==bL2d>VH<f>;[^c:NJTbT,7>-b[JO
#XUDeAGRgZ#TL(VJ0dKLQcMY0+4:_:NQ[Q47c)P?[C-FAH[1OQQT[CA@81\Y1c.K
]MKIGV>E9O:&YVX)EN2fLcSHOdZ,62P4:1;P.HG7?X)8S;B&6(:e_N(>5+54[2,e
@HMDESf_HC\5eQUG3EH4ag__J9QSPBc5<f:7/R5Ea>#FP9D\HR)/:LTH@d(-\dag
(1GEMM[<WdL#Z.DO#Fe\g_e1T[]3FV]MEAMff;)868AY3]D<,>/:eNfBR1L_66T@
bTY7NPE-HW\=.1CX&K?[DR1@VJDQI4Lde7GOGaLH4YHgY#\WY-ca3)/?:]XH)4WB
QUX02E-;2ET4]:X7?-92fB1^8/H)g4_,b-.<-cb<1>N(XgZTb:RY9a8W;NP)LaD1
VegM4W:E):c@988.)3a\aWOdYEgA[;.-F+C&[4VR-QO:5>+MYD^/GL9T3<ANUf]L
Q,@C7.6bI\5a[+(eb_#@ZEV7RTbE9,MBCdYf+T=bc4X3+P0733Z#bTF(M)cCe/P;
N&^,g&MLIO&/>J^/E3\P<?S1[]I:;-)<YMd2.J<:db671/Q5(QQ]^M,JcHfC@2:U
Y-IN]OKHB6=V;g),<D[QLB)f3OL0V]4e&+V1>64a[\OVZ.Na_+_LVA>KCA?cG_FH
J,6EbOA5D#-.:D,M^D?Wc1GJf_2F^Y?CeaNT6=^.9G3S03-14^2^gNU;9X-^H9&8
<9=VMc#MYWN\-5.U?R(g7JE=SQ;29#L+\<IeC#\1#^CP[L36R-_1HfV)H_B<1.CN
-;CL<b5R>?)B/2=BQe,1cQA5dGG#-\LO@QA&A.Z6gF.16EC>TcSHaf]/Cg0(&?P<
NIK+A1&bgW+WI5VdfB;K>=R?cc^<dR@_?aEM3;-&_&D(/_:.BJ1[I0#[^6Md\I8X
E+QY>G/S<G.MP,31c:V?(V]3->,GNMBQ#H+YBG?1VG]I=W(Jec\S>+[5b3E_<FU8
-KE)S.+H8U&^V.2UZdLOT.Qg6IOG+33f>3g:SS[H?OB4<UV@43dAL<C-XREKEf@R
X5#Q0edQB7S@DP^ObHBVMB2+ccR1#HUBUOMDC>T+I#fA@15[MGgE&+REfI(<MNV=
>T29c]H;035:_,&Dd:6MM>3J9RU0+]^\A1EH9d?<dAZ,U.Y;J@3L3Tf+)M[]&SAf
JKXG@RL,I>SWJ9f,=F7Od3PMMAX7/)7T0/,SQVDP6Of=9BOM&9\\,\D4<&]([05d
f4GX_=8250CUf9eMd4/]eSW;+b1NFf>ANV,KF.6VMY\4).5c/BcPYID8ZH^(S),Z
0OR>@W)T6>KU[(GR)QfEd?Y^L@8\=,38WgFI_]#GIe.(>3Q\ST9GE5595\_^ZV.,
@H7^2Yg0[3aPWYONbd2d;VUQ59=8F4<]gCVP5N02<6C/ZHDd<\BE[\/RON=KXD8/
.4dT#ZK9\BL;c#OZ<Z<L8\>8LA#Z?(H_5CE]5Wa-C]DdPET.<3-DQX-HCX_;c>/V
)0;f0dL0Z(02A7HeTN/V0MM?_[SU9@66)/[U_(Eeg;Y0(0.,)3KL4O6NeX-10SE(
Ze/^\Z[QJb.c_M(IO>1Y6//OeW+6BN9W#DS=_W^9/A<_ZE;-a/GI_)+]6LCR=9JI
f=RPCVT4<<&A/gJ[R[@JTE[.LTRPG02L.PR5;T@.=ZOPQP1bF8KVKG(DW/JG1A6^
UO^O6@_>gL;2/S+FIB>(WbfI4D?D;f3)QD;OQ8B\^0U,]_]\gL+4Q&CdS8@I^UL0
<V:C_M;9)dTC+LXM.^C63JH?JI/2JcBY21YKPW@VRF@Y=P-@HeP/a-P=YgET4X@5
USY@+#4Z.\&UeW;=g8\#cAa[@ZG)J9,&4KSg;=#RG\[T;M<NT=N6@BD=,TW-=T@R
LAQWac,:4gcK]SSPV(:9G?)bY2,FP9U,RZ4.HaM+M_L^N=BF(b?Cf0Tf-ZSeUMB,
9g)G6)N1P()W3W+Jac\4__J,A4=XP7THDdA)<:ZY0fL-KCEL<,K@Y(&Nf-EcT1YA
VC<2b.-<5S\ec7-fQc[4JTQK\NEI@=5gW(R4(EcGcDCe3[3aI@[NOE<edI<7J=9^
BOe2;fT]C;Z[DI8Z51_Dca;V<PCUSY0&VKa[?@:d^OI:S,D)3P73@3g_J5fe8B)+
\QF1=5@126_VPLOG8AGFSFFCZfBRA0>[2VOM>dRPa(NU6Z>)U^2QVed6&#c6?^G9
a+UFNKV:N?1)RX),(=ZY/\8-H4fU]>Y+O&14@]d.0R\2RPTY-bW4dLD5dJG@^18a
26SM/?B,I8?1T[EDO(;_B.Q:\IVUMA@ZC>W]aK_UHI0>F.F;<8^QX,#ZO,M7<8_,
EOf&JY-TTQ3JHdN-H:/6A4C:cg1^\+Off7^<H=(JTHeSUQ7/eH&C#GPYM(D#B<.M
G0ceW::#Y_FKa^,1G0]IL2JVD;IV.GFCOAa)AUR:<,+fg8#I8ZGD\I[X,,Wd)2.I
7MAc&Q;4OSabOTKg&_+I?I]:36>DcPHHe#GB=b9#a4Ce0bJIV3#>]dFXa,c0R5^5
3?fKQf+W\0#aM^S+A(af//bYI0.A)8abOcRC0=3GX\4:XGPR_[^L_.0LVO837@Q&
JZ(-[TEF3>Vd5X;d8??=8O9+c1UDa8gS8AEb[ELIF>50?T:8,?0fc@SZHd93YM#+
\88U)SgJA.^4)&>T#5fU1L9@=G6LI,6R3(-ZQ@5e3@I,f-A9>eb)7J0NV:aZLKHG
IBZ=gX<.;N0)&U#A:4>:JF(<<eFE#:++c-5Z8Q[Y3XfgSR0TA>ECM29?eYH>H6)Z
dYW<L8PM^OA;#Y>\XHXbV&b(;A@@VE4f:Md_<>VB)GC7(6OIUU:^3\W.VJXa[f&g
W^EL)b_V_TZ?-WKE?ILVaUDS,WEE6/2V+H?.GQ<cf,+Pd@FC>65NRaFN#FGZAI/<
#5T.cI3;dFDUY_1L<e\gG6U+H)dJP4=,#Od-H#EJPB+>ZE?O-PZ^6aJR8ab]9.?2
=,39BfJ:_VM2AP;R#T#8S(RB=bX/=a4_PQOHR?)aD[;-aedc-PJ)[,@Ec3>Z(gI5
?OA(Oe3]]Y4&ecb,gT8O->O3I]H9gAV[]OA4[4S2X4O9eIf,M(-AbD@aIX4LfWT3
;G-M<U?YD7DIR_2<XYf)5@Q<L9M]VJN(UVdeVN#R>>4:1e-B&I]3aOeJ/>e1.,YF
PIF#70ZGg?X4Kg00-]+a[gAUgQCLPX;/CQQWYD,Ug]&;2cH0MSD8W(\aOSKH_,ZN
be4ZD\.R+I?JWS3fXVf^A:ANI[#d-H,M:a-ZQe./N_]\AI,edBC.4LBH]UJ+a4a5
&e?].,\_.2Ua=bGWK9eU&&/eLE+R(ePU)b[+=D<>g49(NI3;@/A#H)8+VMZ1?RV:
_<,&]FYTI02?Q>9YgNVf^WCbUD_4bVf2J2\<R^T@W-VE[P+T8bV,c^@c??1;?Fe3
(])&Z?TCVE&?[H=F0_H1PFMGEEP&c,)0A3CKQVZVE?OL.g-fRbTFV+(/IbCZ6Z;=
2/LKH_;1<+^ML.ZVU&_0,3KOeP;C<7gXN&6R3Q&A6ZB;JPZRS4IMc+__(^gLN44(
#P&=/fgSPbI[gD,9#dB].F-b6Bd8FM==YL)IO3^(Y_AL35,@MC3?_4&U/#PG,Q)A
OH@4BX^#)AgId)VX-[1[?II1SV&7=d9QQTLd2@1IL#:Eb=e0D50./87S=B<Bc<gQ
32=)A:WK[V(9gT87E]9C]FZ.OIY_+]97]J?D[UK0O.>^0&V=bTHIY8[HFa8/-X\<
?88BH96?AWaX(aER+(8@6:BO4&YHAT:-CV?I9f_VJN@H7ARQ+/TA38FYEV5@Hf1<
dcdRbB2H:0??\b9P^Z6/OT8?.=)Y-T;N#P3K[gc&cHY2H:2Y4f7US(]=YJZSEaNP
Qa+J&d@-LPE>^E6fY=dN)c#?O)PT^W-[&cdBc+aSA2L#dM]9/??9_,WXA]G#C@Wg
W,R(J&&[,?M+H32HLfXQ@3E#(X50O:GDf)(^N713B,#&T?9#?M_#C/RC,2A9C=,4
;b8+cDHM<^RVd>[eC\JM,E121OMD)7PUWY5Z+YMBAZC].U>f^(b>AP6+.\AVYR2J
9g&.&K(KR<AF+P.RO3A[ABS8]Q_Vc=[5;4#V)O\gI.5gGgN?(5A,A/9GcLgXBWB:
T=XOW.&M)Y30WHQ=7UFe9G_@D&>UGTK=g[EG[I1>e;U)fLK:=gA3:X@<<IZC]FE#
#&V;:_^VTA&eU+M-T9T^RU&OGe/?]8b5]Ce/[b:Q-K>L^JW-Q6C<_?([.)GZQIM4
BKSAc(E?[KFfbd,F,(R^U+O0BTIS-84K;EI<WN(M3;WJ;RZ-=9_FSKD0b/f5d5CU
/E_5#cgAV8N9WHc78-Q\\V6ee)-^530ID4I)c?4aQ@<bFG,:&32UI?@@K,ZRO5#0
,cf7?Z>9-\=T9TNRBB[UDAEI)=B)VK_:OA^F4?Y]T5U1[IRF3Ac4=:=U0.T-2M&9
-&9+0\JCaPYC6c)c]X\CVA\\-TZ])Z7Ne^ARMd?EKU^NfR\)[E4S)C#1EU-T8EdG
//1((X,g^D4?FK3ME7SF=f66ROO,FSQD:82.BL3[\4gJ9SgJGQ7[.CPf?:KEJ-X#
g\g?>).=KVGVdSQ65ZBMaF&&3;;9MHS<W+bI,P/V-CS3^cL[+SO-#OD.^,^5)D4D
PDFN-LNAPWWP,L_0QYJZQ(?KH=2J[04]OOD\5UV_V3)\6.-;5E8S0W>=3ZgRbgS7
)QM8F#6.E2@8W+PgL3Nb5NFP5d\_T//V+4+A^A(ZBg2Q6=Q<EcLD\>7O,L3I-41^
@E;_ZfZSTeC=HO)2&JBM]];@XK)4HcT8T&gG?,b?(;B?V&5#d[6>f1W-8RH&Xe4^
.7E>Fd^c?SLU>24bJ.)P([1IYI4,e-0fZ>GOZJUU>LRBaO#NK/BOPb(/3@/:NAVH
TQaRK3@._4HffAZQ6=J._.-86<?]&,K2K5,O[2.Y1eYXUB&UdN[J7B=&PIaKU.ea
__WXY85]R5CPH1\F<4Z@EZ_NA.N-SEge9FYC5ZA=7b-D4e)(<8A23R&ce[;=N2G1
ZfXV.C.UKP5;=<A^516bY/3YE8<[KM_Ff:S+28b/&;>VYd#[]S::T,-:<T,H0[/1
c#-B>,.#.L4H63Q8P27ZU+,V:O-KLRFF9ab4F20K@2@X9#\X-)<^:-JcL.E93FQ:
0L&B^P1VcK[9c\<[c6^IcGf6MZdEWC5@TSOX_6e8fD0\V5,1LGE6LY&<Ff4,GA36
2@dVFS(^9eW3^\+:1-aXEENC][>aV,LJ)E,FO/L:EVTL@5IEV-N[0+/>,?EHAb#5
9:O)Md@S.U\Za0cPB;A>J6_cb21:[Ab0BZ[O[<INI^L#\:/5YNCd6MMKdW\^B#-?
<-^SVMU>KEQ9TgL)\bDf74#SQcAKSVYH72b)Tfeg+V_FD^NcK2fRR;F<f^e@M5EA
?@TV9@A?&5=dGdYe9M\HZ)Y.-Vg]2V-VaHX9TIE@CBb#QR,#WM_::VSNAZ2^BHg4
RP;ZE2eOXO41;-]:DL<^=(?3fD^^-=8@JCG0b8;-MPS37/L;gD@N4?E;b+P#_^BV
RD.T93S=DG9<a=C@:D6??G9c=1#35e#)A9U6gSd;5AI#2V_FZTA^Yc,O@U?B4e8;
<,]<NW7FU9AM?f-FM\N63MRWaYDNUd_&XA1AK/B<gCTN?beX.?IGY?<b_,1I)F/3
c]4PKO6:TfO>+_1]/FG7#\PF[.UVB7/f&)G]DZFcZ/36,c[b9RF[XfaQ&9cV0NML
A0Y2HP97X_31.Hg>WI(S@(&(9;0a#?A\Y78M53dNSbHEf^2PD/=Fg?TOf<9Id#V/
ef>LVWK6B0T?([LDW_L1#MAS)/L-d/94\^[RD>eF=J\0G^DSOOOKR#a:@Yad[?[]
RG@9eF\/OH=.e8R;XZ4,8A[Qf<g.5@aY(+1ZZ\:(2f_R4VK6Yd#d-SNK>XFTb2ZN
DB=8bfeC/K4PR[bL#)bB1&[<1cN0bHYCZ&CJ\WDgIAX#\3#F.&)<+@#)9,XZ2f_U
bOR.Oc]J.ZLW3ID).RZK:?c@cYJZ;)d.OKY30151:1?GJ/01;dCb+)c)@C5KHbP6
dKG;57F#bSYH2eL:#>N)+C[<bD=G_S9&N]Zd-;>6I:_J5GSLe6^[,VZI>#f^)d>X
]Z_S<5?)-87@:]T@ABagW2.HGa.IE@a5+.d?I/F+4NY8TULeZa-5DO;.S<D\<bVL
YYUR>YDDOaM25;gGO&2c4+)@GS>6Ng/#B.f/IgH#g?1\cg2R->1Z(]KOX<MH;X>K
SfK[?UDGegOFZ\U=+#X_NW]PQ+TeGQ^G3R@ZOV^T9WDRC;QW60Vg=K1RSO)=_4IH
U8IA^A:afN]1E8G9;F^R:MNYfT8^\WOd/>]KCEZZOG#U43fd#8;<;/F:D0<gGbV\
R^YQLZ(;F<Ed0>>;e367VH?=C3AC&Hg,#:SRIW6F;+0YC0HUI.Y2-AIZOUA.e=[)
E:4Eg:IPI8g+#Z\Of)X/I_8(COG_@]B0ISH=/f0\#V(G0X4.=cX-I0LGOEP#QbgY
EL.+)3(8b\.c_FXVA_4/)B8KX1>b]@WJE@#YU@UL819V](/^J7,CP3?#E4L?dTI8
.=JX:TW&aA9c@ZNG&>\YXUed4#<gc=?DaNH05X&RHYF^;\QbSaG8\VGbYOWK\9[Z
6]=FC@g?/\&cK3^<HRVX2Ce:;&)]Ed?dNH7[e3(CM6(,6ZPTU:MH[/O,^OaG\+91
<1a#.0BdfR=LH#OFW@Be:#JUb_C>>:4LG,@]CL>W9K=DNed))J^7;Kc.BFIc(+;H
/gaW533OZE(I.4bZ.F[aTH;G,4;T;XWO3\RUa)_[DGJ5TX<eCa_d??6Q^U^<6(?P
YP@_@S)Z[I=Z)GPDa,/4,#VL3XW0aID.gK6?9&@e:3g8L#&8cHHLQQcI5f,IM0;5
@MFN<7Ng.c,<5F)ae=;R@#:8Z:9+XTd_29]F&?=)^geI0XN?1=AY^@MA/dfKg@2C
IGKM7=[FBb8J\/2g4]cfQD:,&H_H+,G(]\1Eb:LWadK7LH8V@T[f;]QQE?FQY;[2
=I.F5\_aG?W=aYSH<)0CE9:@.Vg->B\G7)9d@-[9/Kc#e?_4Y#FAeG(e+1TaE_)a
5>LLFfX7eMcFA\=WBc?=B0\/_2T=Z;Y80RAO,;K:Q&RHRUL.48V.04aFe&P)aJ./
?S;X0c6:J]ZU>AZ\aFQM(-Me0R9g06PK]XZ8AQ,]e(X,Z1>SS<a[91P0M]GC^a];
d6457V:\Xe;R6K-8(^(#FCD381<E,=#COAX0QX?.\CK>K=BB9-:a->U=<BA3AV:A
9;e&a25<[I#SVGAV09W1<c,U&3YY0M]PYddG.O17^(UZc,(Uf/=\,UFY[;QN^eDN
/R]<T2O+7d.YSVAARM9+LXZeV;Q9@/KN<JB/?E9d>=;[ABAA<-e-/FC^VT/1)#[-
.g6C-=TJ(Q4,YHJ/dX1Jg;U6:0Ed^_cZME286&>M?B3RfJ@]AL6g[Vd>RQ58J4>e
D?TY+)Sg)A3TCA\DB=D<51bUR2+,J7#K?YBP,39^&/D?Y0FNK\=[7eZ(TcaM\-^N
E=.(>H@]Y[Z/@K]c&f&5^]&I)/Z__G&S6V:><IRQ=SS&)TRV>6ES-21Y.8C,O&Q/
2W=+;>LMT4W=7LBX2)dXGG1R);X_W<=:F^DCD9ZT.[V/O)HV6,SY@(ZNcY]](<BZ
&Q&)D,-@AWf+)[G\(YHAUFa-T\]If3,+QHXeZ@=PB[5CE;G/M^UGdO_;9EEHe<J@
f0MO]^S.J-2NN7?Tc&YD)EKUOcHTZd3,XaC+^U,;3dSJ93MX_e:R/-8<)Yf8b,/2
B=\U?\3Fc0-1>_V.9bVQR=QQQIUK>V?g,CQd5^M&UEO,YD)9V><(KEYbNHd2M07e
U0VKEa7IG#c\&bc:E,U]?41D;.YH</EI)(4aBH07HEEFTG\=F5/4A>F4J4EPKQ;7
8OXe@,Q]:42U1/[7OWISV_(04V1N>aVd^1@C8U?OXb7=BUB0RE2BX+N\C#V;bCHN
;f).Vcdgd@,3UYS8-Y75R5;6A,CUO[-QDcJ?PT#8^b#9fOBPNY&<+=ZL@fD#F=2.
/6LA9dZ#5KR8Q/6.9.1Wd\JE&g7UMOH>#HWQ_7C,22_b8?O^>OQcEN234EO.VH7K
c8&HI7@5HF&c,^AXB<&cJb)Q(&@[\TW9-A8&0FV1F<>#+e;;F&cbQE]BSSe/-HU]
T?d/UZ6FV1<dg^fVX_.29GH#dK,42@/]>;3[5B?WcK74fF.L>Xa9R.76PaG.?CKJ
Q-??8JAWgdD#/2;]T3J(NE+5J.3B4[+:\@4@GF-JHVMg\0EYF__>NAFE=4XS>P^H
?+eZPWbM(L@=\R9-+)Q_SG16NOI]7L:NG_=1,3(U)?((>fN<7BWBQR:39-g&>U[B
dB]^8Y]H@]T/F?I+(0ZR+2JCb[?[D;NUd&:QGZZHDCQA\I#GZ4HOSTI&QX^fc)<8
6RQNdITM(U/Z[G9/b2Z]HJ?WfPK-gJ](OIPABH97DUeJ5Rc;99>/Z,16Wgd.LX<=
GY)-=Re60V8+5MWg.<8=#0JUSfFOX5f).W_6W)[IY/35<?L;=D2S)](C.a@Nb13d
TK3S?8)D6T;D-)\1[E#eP6c>#?\@G[F/;-Mg,Q.T4;;&aMYDZK/\,F\X)6cJ7aOZ
E+4B)f>[X63b+^YFB:gG32fCM6_)D>QI3b)f1M:L19IeYP5J;I@LI>@>XXW?,PH2
V8@/[I-P1VT6F#ba1)b6[VSSfJg\_3)^.XU<agFNBb6U8fN>UTDPC+=AG/KD1f@F
;P#/>8I1]EP;c@:F]9.QLH#YD](25>F?13Tb]NbKE;SD;a6F?FYR339dcLgV@;7M
MEEXc6Zd_9CMXIE3Oa4)+/b1^05d.(98V>58b<Hd=_g,B.R7>]/94cZM/20gFeCb
3cfa,VI:c<BEW5UAc>-Ndb3N0Kf]\0Z9g+TQ._\XTET[X2AaT8#JLC.;aU(FR^G<
P?AE@b=Tg1dN>30MV]V@Fa5AHSUBO;^O&6EUNd<&[NS?BeMO=2<L/N4-MfTDDF_E
MGKO)2(O)b]I]c5A,\E:J39HMFT#-KNS=D\Nf1E/VU;3+>f(X4TT0b<=^[#XGgMB
L]_,_:HbPXGOTO;;>,P]67_e@(;-[6RXc[R&OBRXG=Q>1@;.K,A:#5<C#M4C?W9)
\(DSJda)15,B]NSSNKJ8MC=B6VJ\\S92^ZC#R-[fd92=EC34[3P[Q@FIW5;T#J29
,KA>b;5<)M(1:OdAAec>QMMC6^KYMKZ?-3-=aDW8F=#@:bAV,8@XHg)]=H4@X9=J
Q>Ma[T3@-[KLgdXM132#dI>V7MR\aZ@89eC[aCB0(0C1R,8HROFE\0J]@WYGPEb^
A1:Rf;Zf6M(+Xe1b&^D/W(A4=HJdLY9-2Sa](>1=1F/,JMBB;(H(&YP\GMbR\ZGU
a_Y@>UFNX)(Y8gAD(#[-LI^DL,([TIN,[]eH;?\30\Gc>@=X^\E\_V/=f=MQcSRZ
<SdY+@_,.CC7VPb,>6V+Z6.6F_;Ia<VZTc_g?1\EJdEb^F?KdJ2;bQM<GN(ELc1Q
ID46d00[RD,T-VCL:2(TR)R&Bc_6UK0D7\7M<9e?LJCa)RG<?39RO/Je+XTR]5S8
ZGQ0-J5aNFX]E=>@>0[f^BG8^)]DSZMTaY+8,Q74&aE5+;,7KgH-P&\FF^+==[Z5
;M\J:XM[OBIEH5.M6>44#DcX9-3U3AL\M)X?,+S(I\3cGYBM]C-;&DBB629MKV:2
3UG?6Ze7g^<8#TC>eQ;B40;]O+41DHOGI@L<7/WeJ9]P>ZcMb+E?G9F#VN\L?N;I
OTG+^Fg;.O9S-fA1&(Z@=Ye,Te]C(<N()+6&+X-,(?--G4/S+gVKBSK>RH;,XH&R
ZDN+;Qb+AaV?T3R4D-2>_E&K.2I1^8#GV6Xa)#5?3X0C@(T9G&7UP-.8K)g;72_Z
aWOc8?BJ:HRM;W\QBU\dEO=+H59\?f,c.bN2@#AO<9<a-AFOa]E@?<V:cf6TJE&]
#TSD:+&9^/f&R7LH\@bL@A4G60<<KffRdZ<9+UYGPZ1-,D=K9SfXAfYS=CN1e]9>
IW[aFd9^7U)4OfZ9@3GgT.9:.W[U^5T:>OA^Q]g]A(=_e)49@#PBMJ5gE6dO>5;e
.QP1U=/R1\<&3Z1+0a&DG\[1IPECZ7S#1><;e+K;IIeX>K0BNKHFgW@LQ:#;ec@P
Uf]KUC#/SI^N@,;B>KRHc_+4)F,[]B,(SDY6:AW5I:e=<42IYV(fS.RcJ6GWWXAR
eH=UGWWJM8.aDCR[Dc[TGAec72:CYZ6JHYe#CL1AD^>8\-<#\+O(X;Z5BIbBEfKL
;2&P-QP\EE8[DS]16U6d/fJ,F>M0+1b@8c3)E)]]])27Yf=3+UZaGN2PG6ZFPL_\
G6dF(_1(;@YfOXL<:93NJ)A45E]<[W9F0aF>B4A_5RFB.?b1S^/FcOU_SaJ-KC,g
TOT0&S[:K(CMGF&4LUY;(IcT7;QV=IQ58?PG?0]I,9_9-CMeE47cC3XC[7KA=>K_
GE^f\=QH+9XYD5V,d2A3,NOYe(=W-0gP\0_cI/-<O2VMK0_,+MgCG\(_N>5:#Y[M
IQQK>E+>Y5<ReMU8YOA_1W_XVaGCSgWf=@UTHcU6VS>WA/KeCTdcG?<3SZ3+5LTB
8Teg#LK/e/&2ID4-IH)d.beaaS2Y),<=+:]ZOd&NPRLg^DgHDH1CFT\W]4QIYUO4
_;3;RAC0KTJ)//]XK]3&Y[aN&dbGW:+6FXUCXNX(0#40+3AVD8YD=/Wf\3d,M\ZG
a;9-Q#4S,\#WCd/#M+R#,56P/_P0FT6TE@P)a/DdWQ.BTe3VZ34;>4XQ2D\eXgTN
K0b4aN^[.0;9G?f>O6-P3gb/6XJ9=,NQd4bN[IKMJ?T9(G0MAJLgA;@=^LY8E0f@
8]=eK7,P1F7(0\6UIT#MP3OP6?J-bgf27MH=LIdB;VJbF?X]1d=HDgg1fP[RfH8W
C+U=&>Y8bbS&g>c=]YGANSQ^@.eJ>J9DMA0A)D8J,g+?e_<;>EH+=<5O=#+(gY\H
:UE#bC&+b<<JWb#+0ZKfVd@&YW<FdEA#T/2L@Ng8Z0BbA;@>+He2R_Td?3NSW?G?
MNSCE]P1#-V1+,cJ3Jgb[NW9UAG3)TV43<>[BWS0(B;X?Y:NV@?<Ud<d\Ic&2EW5
Q40:gM</K,I8R+0),X(2YT?13^Uf8bS=N@DTGFLdB@9E[+WYGQJc,@T3]VF88IO?
@EeV2P4H1:eNGG:#(I63HT_V^A<\W&8)N+X&b?6.Q:N/KgTOF8,V,G95)Q:?/+E_
:a^2F.D:[P,4[7X6de)/cMTCfd6GBbY,B]MXVNE=N?2CFRT.<Y4>D_@H4K4+[-0<
c+P(QQHDZG0M1IBZZc7+/\^OCG4ZfD@]QY>MAPSN?dM@2WERV)bYQN\614504).W
,MHAQ6KPV-3#CRF+_6=5V=0gT&1I_0g&80[DGP@VFMgBfLbK+HYUGACY/4gf5>D&
ZPc_f>15J[O(@OJ2HV@U,V^S</8;.cH)W7VcU#+C1YZgXNF@e-OO3#f,@d:8C#5c
/?6JCP(I1]=Y-b18IP\[/0?0\5^)EE:Q2&S65AVS17dBf_@@b6D0e:7]\GHOEVg6
5O4#f[Q/[511_X5=A9]>D<,GB(:O1NVgF<O;AH8G<\E:Pa=Z;c(3aXD#Oe;ceW[&
WKRY<&+M#cbM-0DKCYQ#Md+&,,<7Q8+/4Z\9)4K5@e3O.J90IIE/?E3gcJKZ3^Oe
+T8QV8P.:HL&5@^)BA87fH[.4\QM3H9<IBNId8L37YMaN6DGND;EN/Z08JW=_;2Z
M+#Ad@6OX@=T:N\(U9(A[NbS?I7O;.RCe2TWgYf80X^[9dE?DWZW+7KM<F<S./Gg
bK.T+aRZ:KZNMWD<[.B>g2e44d^&T8Z^Ea;a)VKdDAS7.B9&Q(B3CF&H#PI[Q>RX
??_c9FM^+f<.Z(g-7O^AUEB_BSG(b51HZ1CY>@,8TH?@P+[6V?b&d>T>#/OOG5I&
8QQ@LG#\7SQgHJHJe??T\8)@=1FaLH)@^I6STF-^QGAU^L3I@[)AH&)RY-=F#G_2
W&8X[9B=BI8OHSb-]-V9>?Z#G0M_^eJ>T^>PZAg:4E&4^4He7_D/gA(8U&#A(.PH
P/;,/-I,?9Y1LNU)0LOSEI(XE=LX<T.AB5.gX.7;:Y;gU=b]/WLF<?-(/OPW.:8e
^?-9a?eYT-R8NTYUeO&2<>->3B20cM,C+2+0N9P8_,]ef/?OQHD3/15b4gX1,8YT
:=b1Z=bS;N<ZBeCFfZ<\a\[IOAb3c:P@g5:5@0:?34S=Pd)VEF679/H9c/X0:Y.3
ZW+3B@NV[8@+2gKMb:G@JCD=3_(C6,_Z/Te45O>d\MS6:SYYe5R[Y^XL?_U[UHIA
GM8,?&TV8SZ?CX4CMcCW\b]XPH;/K.PePaNH[?TR61HS)_-Z?[_Z0:6(^.B9[bLd
F=4=?c_gIP2UY>UIfAF,PV09>Y0cDOT8JgF=WHSWY?E-9A(+YcI(Z\5:^@289?aP
S<OQ.>e^X\JTGCH?XK,a+Y9GT]+YMCT>2?\WIY.4J>NH[9.fPBO>OT2D8^[KdA<Z
J7R0OgBV.4(1WMC;Y272B^8NWXV:XDPb_P+\?5#g2+O]LS-RA];fOEP/^C[(0S(3
52I0#ANAH=_\=)-BdGUB;EJM]8RZ[f&3A6\d(G;C\L5(8^V5gQK#-eR+\8@0QW/4
@G:3Rb+-bI]K7S9GL]MWLHH6G52I[JU.@F5.CE-2(;#45405IXS,^VdY;FP]3.c@
<&/B:M0K7>U,[@&K1_c>9RC.Q_W,V-d#\09#9N;8@;e-ED2Tgd8EIaVW#-A?ZF<\
.28=EW;7_&fTTY?1E7)H+S.G?RMN7W3L,V?/YDH^@)P]Rf-Ec1YAQ;I3M@A2Te#L
#c0cYbQU;e>NW(=.0_68F5P8,<FR:^SL_[NUHWUWZA:W-+H3\:g7TJ<eWD\CQ8D5
C9.6::MG>gX8N\.&)PRY_a@D&Y_VfE8-\d71>2R,RR6YV\KD#(:90Je2B,YNN5;(
7FO2d0e?6P[&DeQ_[cD_9S8Z,Ze(5I,P)M.D1#?4MG,DD7b?GN.V-^dLXC^3QcE-
5[C^NDO=TA[@SVYa8>L)A/<4>1&+JI@Da^BQ],f4f3a1_PJM8AYZ.M[8DfC(9KE7
)SR1^/WQRA[\DPaaD(:6-I4gM><fXK4>I71A_C];=+eXHBOX_M[.K_ZJ;IEO=R8J
R]F.0>Z#+f4?WN++H+6WI&X-NcK3.KFPK9WJZgB,e?[T1)U1RVY\a<H_[0-QC,<.
&#;VQ>,57cK5b1XIPM2&.7(N#3V,?<J^T=0cU9G9?fAb^Y7+UJ;>?e@XAU14a)R#
KUZ5aC[?U83_)OSCJb)_6;N758-d)7_R?V2HW/^D_-D^@YI)&N([Y;W4KF>##84_
aQMgS5.#=H6X4LdCT\3=fVY>&II4Z.>d5MA&T?_._(f>Q_dE6b6+55QI<]5S4O1=
L>M>0>Ab^H5?G]97(_]YTFA7[U3EQCeIc7\D1ZfNKE\&#(Q_L--U6@,3?1>1+A6B
e&A6=CRYT^7BS@[1gJ[?,&\5+Q&)cf/[\g-gA7ag9FK>X(/#B5<aV2IXQ/aP4.\T
M>)XbPFXd45D&74M:;dP#EG38-]A]J8@/ab0PE8Ue?LHV/^465KOR,Eg=G7Rc&7D
M54S19C:<gASALYL@BREcZH]3D)F/LB:;NHeQ[K4f_;,?@/>;__#QJ8STPDU.6YU
3VC-5(D5#M3+PAO\//>eF,FdAQ[#(@B1\K<DcQ;ec^41g_PHM3T+LLU(NV>ME#.f
:;)@V6#8VLIE>6U7(g+ZWBZ8=?Xa2]P=BF-SI=X(c,8cf/#<@JLWO6D\N31W(XCd
;U&@)2eT_S;97HF3Y#VW0-9]gFP;(F4CH=5TX4CaR@+I1FJ&-X-aO:;)@2XZAFdM
a+@H?)d^6??[Y.#<,_OA^dg,@#?BQN[\+L.[;-X+5Db=N-@,)S&3M_eb88.PbAW-
/ZKTUIE3d)074UZ<W.9H>9_3@Yg=;Ud\]23,&6[J@&g(F4].]7B(A8IBUff>Q?5S
.1&[WF(GO8?#RPP4L78HP0:#AYNAET7-&UM[edD])_?+(#?GY_OF@3[Z<c&HOb6.
G;88;HUJQ?QcZ>V/J<(PDg)1Mc2W->Jc3JNR8CID8N:?T-NKKK0d,3E:DZ?aK-V7
T#M@B+V<W.O@;[H9f)BUF9Kc[?CD;/8P(13BRfHI+Qbg41?F3+b1eA7M(c:K<[VD
#gTSFU3NK/:b4)TMAN2=Z.3KEE6H<4Hd)3_&;4,X8LX9^Q)DHZ^b;]6U#L+ZA3ZN
VU[R7O<8XHB^S-V4&WcBF@SAXOe8[3WNUF1]@M)7O3]^_J(V?M-B1PX@05MK8+EW
T4+AKP#2G<WAAUBY>DI@9V+_a:Q;MOe33HW?=f+:;.LCYDHL=O0LfaW3D]Gf)@c.
G>:6DKfS)7FTb#1+\WJX+A]R&e@5cLI0]_)6AWV<\9Y8G?[\>=Ye0D@#0aU7YZ=G
YFd&C2SCN:M(e9<Q.O20<?7T>OSPD=:W816\YA+TGB;N9#36S#[-6[C=R++KZBOa
bE3^D2:M,M:0I],TBH?0LP,R.@5cIOG@\RdeYb^X@[:ZHQ2[URJ,OacDGI&XR1dd
WT,E@?L#O8Q@R2[c11O#3gHG<\]d#W#Lb@ZR_:)5P.8(EfHT,I1e8O6g3D;U(R3R
U_R=IGcVaEXZb8gA&#dEWB6Q2],[GU+6F++#R)^>ZZdYf<+aTJ:D[B-H2H#.:UV4
>(R90;.@b.AeXD7?TA?/g+HN;L:6b]U[>D1ae;F[#?VYXKJc((2KFbdWI^[T_^IO
O^\0FNVR:^f5+6e42X]-U<,4Y8Zf0_UDOd1:^efe\Y>Y3X;JgZZX3JZ7e\?ZHS#H
[6P1)L7b=>R0>BDSJ1b1Cg@QHe9bJ.&4dPe73f7NU8JdMEA6/Pc7-VRXgg3e:ESc
?H;AcWR?L3W\fJK]6I16:R>J_KdFd6X#M0b\@<)X1/E9936^YP5EE4X_&J)Y&b6M
KT\0H5[FS?dfXK(2eL]+8>WJ1BW#>#MT-RZU,aJGAK,=5(_c1+?7]Sga))E89C)e
OS,^)YfT,FYHT8Q;93UVJLGC<NBWeGD@P^]a;\GeHA0RG1FL4Mg0/S)EW6LL,5\5
HB<#3[8>H7g0_?TI-EDJO/;SE:>B^H=Dd&gA?-FA?2;X;8I:,U^RH[<];,C0U]C9
:+WV?;9)Y]UXQOP]>0\I78=NQbH]N8=5EJSaa[TV:EgNM8fRU3Lb1LU^@<RS;Z#&
A.60B182,9FQ0H#N;,aY(9+8^\^/K2<QD9O8O5F>3BQ6BDL7N33Sg+8dRK,eVX,2
/D-@VK#^B_I4F0\UV1Kc:K]DXb>9Y\_GXQ9/1N(bL49<TaO@1)OX_HOO=5]/1&J.
8f;.HXK(.#K:[=9]</;dZK</NTX;],^1aW_O:9\(ZSM=M@>/6O)J:DUE0-H0@><G
^f1[NLZ,d[TH/;B4E9NEWXBD9BX_KgK^dM7\L:W7^2H\<c2SZEHgYE5A)N6E/<&3
gX<FE):0I>OFd1CDD53gST/;,aR]Q[>VLL@/9T/;F_1baf;#_YT-Uf<&83^T>7#_
#?IS7#]3F2(<S+@_?44^=H\CW\6#R0<[PR#fWg33\:MCFY.?QHcDD<.V6>T+Y>.e
LO4Q)fZTX?<^E56GT8M[.WUABY:R5[LX9/?T?U,M-)K1G=[-XQA)W@D9:1BNA;M7
&gH2I+0aM9g2C/7f<f^>J0)<AO8G1(4^U.<cgIL-e:K8?<T6Z_#/e_dIE61(1_>9
YMU0O#/@aPT;67_J6]1X1H?PTfX67G,9b7;b9,#1BXJ&??QT[(I:ZP\G&:OBFR2;
bGIb1(9XMI68.-0]=N,M2Tc=P2)4F=>OC:E&KF3e99JKSe]8FR(1BbWb9g4O/^KG
+FH_\;69bY61#f6De\27T6CNV9H52bYKB[N3YU8[0CA6I;A?==FH\HP;?VU5a+CF
->0]>W1-,7KH?X2HN9+7XgUV0)8_O&4=FPWDS9(5V=_U;6#&>JTP,3Pg.&FacZa=
<1dD5[Z8/CEK12LFX.Y7QYO&I@NBXHLe512H3.V_e>#B[Z18;A)U1]DGIQN_#^O(
O,]RWB>L1<>JL=#e\\)?UP92[2;Pc<fW_?a[5?EI/[7FDc&efKL0A\Kc(f4JDOY&
+:g..HL=^CJHSS)ZRbXea@_M04XcJPZg_WB4V=cW(1O1Y&PgE5b6Cf[1LA.&b98D
-ER\ZC2>QY&.QAI3f4)Xe2J;dU[#=]V-/d@eUQa9T.M8H08SV-PcXf\7^5_?):>I
<I0-D1)395X@.3BSAPR2dMHd-F3ONLZNFe3/aUFKZW@TeSEQ@D<I<L.^.:G^a0e/
334N_c)C;7Wf.MfYL]U>S8FI)==eO7N]aMA-:Y?c7\eA6B<[,f>[/_LY\FC.e[31
B;8KO+]=8LHb]I:ZSe?&VDDZ?PX+6_FY=KO0Ng>31]ANR?ac=LZI&SMNO^Mb;1]4
=<ef.?GD#-Ga:c:W;b&A6IT28?M#A@SdD4.#bIH_9ZM-/R/J[E+;&dN6Kb]<O;/J
E.=dO(?=+<0;Z8QT6WF>b?)4]W]NCad?5EB<C1D)0e(2QGC4LV./F7/F,Q_NXT8P
]JY1C7-Xga-N7O/\R=/F4--.0OZ=^33-N,BSM;3-G5b2R0YFA8DB.X73HK(D3W5]
.RQEG&MW,/X7N4.+f#-bI:KYBUd1.&b,9+:I4bX,81e[9,e,d<9\LD;FJ]2Ba:@U
Zg[4SfWIBEa4gF:IefbF[c>-G=gC97XOJ\V#3b,gXM;G2Xe+YCX;^A9T+S/D34/D
WVaF(=V(c^N_8&P>#:fb6>+XSD>?N(&>90BEU+8@?QPJ;)MEUNOS5;;_FWeUD\?P
@0K>9#_f)\Y=GD]^WEZHIdV\:6.901JWMB.G(7]c8/)X6U/@2SQ.YOL#M[BX(UZM
UMO1c+&#+b12+1eQ4_+g(AW1;I_g_HOFg4,?e3aJTdSIU/-9fD4-HTbJ)QZP=_If
.F8a#,7NBbB&^>=?CLOgRc&)8VSEV80gS.c5;@;T]7-+0\@15O&TgLc#d,^:[W^H
6[>Q<RIE]1;\ea86RFHQ[=A^S3DQYPEAeU#<HV\R9W-DK/aXR>-52^.]FO@X/C@3
H[5gX].g:_L>#I<)]c,3=,U;LJaT6?,a>PJ=4A-cC@\0dNLZF@\=9=>bB5==78O<
N#IdL:NB7([>;[,5T+MHU)b#aZZ&T-R.M?Uda1T69^8HTNa5c=1M[=A>?1gG,4Q2
7?=?[;:SAd9/FaM8M6eWBaAdGHgO]S[0Tc2d_>,SATVJd/fe7WP.Tf>c-0Ae+[DP
c-KA[BU5eDB9+a_A(Y=85.?a.Z++N-a=)1UOCaBYC>P\:VCVBS[]WGZ5e78I]@16
,d<R8_]U7C]PUP6bTBZ,W,;Vc39#5_?A/g_.:c?gDSGV_9QX:]\[NADIb<]NR85>
0H,,0KT.Yf\^AP0,QRI-T9;:<P+MTIGSe32^2_^#KU1&HTH)9+(Sb<c[91A0^bD,
:WNQ^.OOb<6-)aWU<NbFG3/Q4M<,>T6BZcU^8ad@aBX0b@;.)#Z+FT_6MUM.K//g
cdM]fC2Q<Y?[X1e,^eDTKQ/]N=X_31&P6O^(=&)L@/AC(HK&7,<JdO438D:RN?.0
?G5#_BZ>fV6Lb,/(BPQD.-EM,8fU):P>AKIKT7T^0Ga+/cKH/C.MfcC8+WY+]<TR
##.JG:G.C?H64KMY;[^[HD2DH&.2c,9>TF+DHF+@AW<Vg_0HIH,@1Q6;Ta(7[a&&
NJL+bFU?N#CVLS\W7D3[S7(QR>O&^G0cLV+0/1589\GJG)BY;P=?T(XZ?.5gG<VT
[A=\&=NTBGFX,+Z.+Ca(;A(Ad#M&X8/[/AbMZD\fV5F+/.,C(IX&8?Zc,:2SdTE=
cb87OW+4,;KU59egI=Q2,A295bTc8K]VeCM5-;5:[4;N@[?GASJ,d?CK7TP8DHC]
.D98P-aR6OB5Y&;Y2>_7F)cb(4#N,@)BSbBXZfDBNN,C:5J2)3^T5?cM0ZK54;+c
]\0cG7BZ?E3JQK-O(C?<VU.P1I+\&5CI4b)PTW_I)5:f/c@/(JaA:;Q1dRDXJBW<
.TJ<.6<KU0++4c=eQ)(]+V9BFC#.<W/W=C,]V#(G567e/)(e,7dI=6EPZKIfAZHJ
aO]QR-U^GaLB;G<Q.^9=D@X.<R@^FNG0\=?)A.)30TL#+PF-T@?5Z)K7QB)]BJ7H
<DZBTV64g9V;@(YT.H=+1_N/X5?I9QN6ABc4f<6T/-YT:98E4J:+-7FHN[/N=TWf
)0O-O&NBXQ43TBdA5#/E[A]#QJ_CeN1C8D--->OW=1^)e79_O&,c#g[Y^(D8b0FI
JMEGBbL@,-g[<>MS):(Md@RY7X\HV\PAXBYAY5H+=V4#Oe_D0OU&7;HgG[PMZ#Z&
3:][.N+8,S,F^@G=9#+)7R3R1[a0VNJa3[e0?:BRa4OAEg.665dVO1P4A-TR@GP\
QKP/+=a1c(20cKDJH;fa9-;5^Y[4_WLEC&RH07;]AI<_a6VSCY-HB=D#7aD<Ec9:
+C;5EBR@)5T7R;-e+.5ON@;[RQc5WDN[H3970C19cf9E.9-Z3@/EJPH3.1DM/YM<
HZ:B90-3=2:Ra3J^eI80WAd]Q8W=5(.5_&.TT<.c<CI=YM+A7:A<33._bGG<\51G
6Nfa2G#ZSJ\G/08-1X>BYc(4NMZVV_fGETE+8TW@f4B[49B0F[#d;C74EWQ-IF/R
V>>g4gLAN,?Q2:gZOf^V_fH];6/a160/LMOUW[/YX_/g]N?]=@GY1ORVZ[SXO9Y5
eDcQ4V5V2Uc\IXdC0d^O:H?eV&V]GY87fO)KB/(1JCWXIJ9Q?MSR[c[5#.c@[JeF
G(9025Ag[f_>-[L&E.CG[/A/D9&NMMA@59GB+:,.V:=).dRKR+e78;ECO-RaNHWG
K-#;P[RULgC]c_>VeEV<Wf)6#eL<-GOa\[X^C\W@6=3LBVJ^?QZ+P=?Bc\7,#<b,
C^B9S2[7H#bf,8I#[,98Eg[^961OB9K1g7C>(@d_1(<8;A=M;3\89-O1NRJ_/-C2
#cML;HFAaUGYPDHA89&6+.TI>H@Ub#-VC>f2YK+EU^+K:/HUV@(g:57CPJM,<L5\
T2,8J-:,Z?e.RHM\FbbL=(86cO?CYd;2dE][X&2WN8R55f.4V]=AZR]F&=9:QK\e
[Ya,?dda2V64)]@Z+^Qfg51+MW.\K8I]A_>4BffW,#H>V80>X>-I)S/VA=X.EfbN
V_&>_d1_B==DSf,N\/TN:9b31>?:8P)@-gKZ.gF,TcMI?J1AWJLCQd2cT/QNW=6<
WYVg6(:]Ub,)5JY(126BfOec987JR--GPdKHO1#[SI[P?Zfc4^-G.A3FbVcHef2C
eDV=e;.:fXe1;TEZQ452NG?.:-7)#@/Y9.CO8gT1VLH\EVD)O:Ad]I>BaeQVd8UZ
):ASOHIT,IM6YK<3A6f-FT:-aS14?Y29L\+[N_9)=I_6D,TgXE,_S:g:b>TM6QQf
00Ze3/&SX<,AP5Q0_,SEg8/(0FB6Z-7bP/Ma](E:/[W_2MSI:BPN[5b?V]R(S=P/
)9S_a)-e?b:Z2FY]/F(1G4+cJ^NK?f8cLU0-K2Zb\NKB)0XaZFD6B6)]N)R7#GW-
<VLP)]+2LRJ]XP9XeO#TY<-,1=A+U0R2e(0[YG?]:_QZ8#(?S^0?WO5ZO-OeRKE)
8TS:;55DL.3UGD;c?5ZKK:?eYWJ2FQSZd1S;?UH\94RR2:Jg/XWc5L;2F@:+D?g;
U1L<\_1P(IF+36Ea<4EZ3?@TSLg_O)3LB[g6)Z4J&7a<:=[6;Ha7UEH8_OQH)/H?
L2+)2a^[:-,9&CWWUYY?\+-L34CW?_JC8M^N6L\,@=+;?_]GZ1K]/8UFPZMY5D,#
Y\K[-II3K4EFXT8R/b.g8+,fQ1B\&>1C+e48BO]<K@L-M5<M)+_@\K>J1BI/G?.8
#Z.U<6e\([e)NQ0B,XfU51MU]=dgSbQe5YO?g3(6TY7Ae4W@)I3VU^a\;MdH?]OF
b);R;\bESa-&4V;ATKH2:0+1]00/e5V1^QQZ_<_T-Nde<gV5(;e2N8C,J\/SU-]<
0KbXLJ)#E.G_J4bXPQ<#C.B_=5X8Z)@93I[@A\#eE07O=J8-NEGac.RbK65JUNbC
[4>:3YZM:V\3dEaBJdW:P87\J4)A.NaEZPQ+4DN4GaV5+L>XQeM1c0&K\JG4F#-a
QG24Q]Z_^H/7P_.X.JTRc;a5U]^_4Q:+dPe-.ATe^3K9NRL6fD.ab_#=2:f;GY5E
Z_BO<##?NRYU;F0MT+Z16?#8RaN?VXL=098_[K9\cD#?7ddZ=@FG1eFX6C@EK=2c
-HbQ24eMFRKW@1(Me,;<:gV@=UKOISc5Vc9e7:P-J].KG)LN+H]I_;E>E37V1Z#f
0gOUAD,V>P;cH++-?;3:.(G.H)1Q^[bTCC[VGMYa\=PB>\LE#-_:\Y((6#+)3[eA
F6)-.0CWBTJBdC_[_SET_6,0\C5C1>YPdR,BM>0TE^\A).2K+]>Z+/5eK?QR#-:4
b/GFIMD?:-#KIAB_4_;B(Wc3KEKMHG\.KUKc_LN,3dgDDS@=dNTVSS,-:U[/CD<M
O9E?V00\I6df9M@(X9P-d9_0&S)UC8X,ZR0ff/.]>&S&OP3O(/,SO.@4->C621e5
A^T,^[YR2FR#)ZK-OZ(E^>5>1=D:B1[=cH5QI7&SIQa7Fb;Hf@eG_S.<Y+MGUBKa
E=(Q4.487W-dLFB7Md0FQ?]NN3N:b#\>D(R^+/(7T_D&cYK-14a<b(E)5DVNL-;Z
342WU4XU#.cMg+L3SR)8GP2..^d[?RI1PW_A[11;V,FVPF@_-;T03Ncc81A\PU;Z
gF[8g23VG/#R=;\R^B/\8H2FKN50;O;C(M[e60V(<6D.M?Yg5S\R7KdA?]Na(+L/
Ua\X^X&I9O60@.a7=-J+a@QD>-R+W._HH\:@RANbDN-^I-F1c,R0TIK>#>?MLe)J
8CZTWY)A8DY:807J/Hd@Zb)Zg>[]P(gQ5Ha]+e4RHF/#a/)K5HF>@BRLJ.RV/8SW
PT.b18]abA8K7fUcNO,Yf,#&T8>[VPAYQTIgI(KbPQ)WZFeBdLQJ/A7C5aTZEDE\
WD^4[2=RFT]5-LB9QS#gG-6EE_(,_R4T30]^D40)7G(N-(Y77G,UT][NZQA1JfdX
9cQ((^=c>O2G]7V5+c8bW0eLD6<4(;^07MFd>[H]VTX3Q_\eY5HeSJY@^HJES9K(
c5NU2K(CR<K^L/(-VP;LTY2R;:5]5e^2BDGR>@V&SUe./MHQHT6OENO4J&MBRMG+
LHN:@FU+)T)Vc8fJBCL9)<X8Y)/e>aO[[OJ>N64.C6S_HNG]52&KU/O5WS//)R^P
a+\1M\2/F&JOeHB:75L8OgID.eH5CMBFLDQYWDQ<P25d>Y\T6DgY\Da+,OH4F]_@
A0\WP7YX.#CLFYg(?4>^Q4B?E4_PU0V;36Q-+WD7V48MOeJ@2\H)YKE/4=?eJ?TS
](WY)cW(cD[Z5?#6@QCBUKPPI=1RMN1d2?b+>43C1.\:5@(a[3b#<-8E^6:QDW2-
QGgPF/IP6BYI3F6E0WdM[/AH6&KR>[?1<^:.gS3EA5-a4VJ8E4\(6_JebOEN5]<H
)1#&+5LL<=:81ZWD<12.0T&S\9)2]#\B0+WRb)VJe721[H2gPE#N+XF)Q;YNY@eV
Y/cJ>SS;_\N_)7MQV>)G6feFdbX#CO@&I.1)ZPMdXgY9UdR?PcRH9;#J[ORa,Z\T
cIadHD@d@)DO^B76f#UUD#63<e^O?O#X6A7#4944KA@DT^U9AU+ZN_>fR[E=6WH\
F#d(G7AXE(Ae<U&fgg^,g8YJ54=WN00<@RXNd?SfO&,#X(HW>ceP2eW7DAdGcIV1
Y5)2MI1CG@[Od+IIZJ+?-,&I:J5?@>6-.B6@bX#-=6BOOPO:NL7C3&5/Q8>D^NV+
.FTD:M:Mf(fGW(dRD)H8]&aL-AQ^-:R=\^L#3W39bffI7G?VF+(+2X/@bTAC+b-&
DCS;O&=V7]0@5)gDbZ]=;HTW1<V]W8,;=]/aK/QOTN&PJf[44?>EH+06=;_DI(W,
,:;/T[=A>(3UH9CE44CQ]8,M&V5,8F>OC06S(,CfbIZ.F<.)UPg]]M#6-M9#8?@O
ZEG;47[N;Sb</T1=_f10_fJ:X-eUPQV7-2Q0]PfOaY>ZC<]EXbG7[R;Y-5Tf8^UM
g)eC+[cPQOgT^(6W&WI>HK1EIN]P]ITI-40H[D1]4]d59cV9[-,MHR9B)N5a7VFb
TRZ9cTBA7W7R_O2TYL7beSge-W9@O>TAUb[WZOW+_--5OJ2]ZETO8F>7B&(CPfUI
8NIA[M[6aO)H;YJU85TK9-)6^A&4COYS06^06&IRDIfU7_415JH<gW169CKcDT,d
N5dYQK.9P9/[:1C)Y_L_7/?d3C<_[4Q3-=6eHB-MWV#SE_\EY5/+KW[NSBEFE#_L
:GVH9+[:O;H/NEXBVaD<V>-411)7<;0\-<ae,.-GTXH+Q0:I&HLX6C^YRe<\HA_9
C.eJM+1T&d@/-BIQQ^E)G.YJfd[_^=Q@3]J1U/XE]EPWF\(#N1Y@Xb?D:?TL9+\O
X?0#VB,EfcF/KD4bf9U#773Pb2Ze[E\RV2T;.S[[<=#gN)XLDFYD3)85F\b?^((M
5;;+P@1B+9><)2b<.&IaF^]X-+-[Odd#<)PJ:>QP@ZE@6S)d#;@_D.32^:1Cg6]^
VYH@V47SW;+Q1:A<6W)fH_>,92B;e=AG1O@9).9a@\Na.VB3XVDebK(TG2W>)9CP
TK>5MN>2M50H.X1MO0C(S[SWB99Id2A-<#4#EHH^HFN_@MCQdET?(8\0UAP(Ef^\
CeZ-_0O,;b>^TO]B&B:J89_8+c[OROF5;A3TPbN\217P+gL8&-PE13[#3=)-&;VO
Tcg?WVTKR<Y;JKVWT[FWBY//ZId/K@(JC,e5<Q@<U#8E)FFVRH=b:.L;#1]AEF#W
11)c>&]0,8ZMUe-eE51D0Y[-^-X0,X]b]DdW+Rb]T2E5BHdIH>V+03,3SSD=/0NG
HGfAY/UO/&S24J>I_0b4Yc-5=V3&T?^,JZW,>GTQP&CALA/,4aEePTd?/YA0)>]4
<]]@:=#2;fC2(BC07B]<F\J>75.=PPSJSW,Q@IO^[5L&2P\TeA8YS?G53/2L>I/Z
gUT/^+AD&V4JcBa]YBJNF)=>FC2KC<BPFEaQRP363Q(HY9UdG>7BG2_D#K2XMH)L
/fH9@^:3S(a7,6WWY7g.S_-L:F.Afd0Lg8(+PPL]PAU7-CT5N+aBI:G/:HPKNg/+
LA.fSBcfH]UVPD-_1Qa3.],[DE#aKQRfEF8a1N=H>AT8Jd2Y,1Xg:8V(8F8X<N.D
?\KI.+M44f,FX[=3H/YZ-T=;Y/2Hg&Lc1T7/gO.E6Md21NLU8M9&L@XC&f1J@WHJ
4&/Id.M?M[W-1RY<4dC^V^bH#gHA/O2PLKgXG>@,&aBHD^/0e_/ZOJ(1-]#,b<RL
;#J70HgFXEFKF0a\WEcDf-H-ZQE5eb9]2M+b9OPf[>?WCMdS8X21#_03<-B]5=F#
^)+6T.WH^CgQc:++4?9TY3;T1QED8,+?TOEO_K87g>YA8POIBW[Y1#^d5#.^<)X(
<=\#b#EfV)/D]G:FcD8S-#>f)GH;?GJ/<(/<_=F:WCHKGc_IF\UX\]J=gUH<K=^U
XBJ&@=S\Y,MR&;d,fC)<==]V6U0Ba<8A+@ETc4UH;CP/ab5+U_QdJ>@.YT=]WQ;X
N@[Nf:^_@F)0&>b3<W].LU<2=;d#??ZdU#Bb77#(/OfQR,]-/NUeeg-BUd@&X;UD
Vf3gEeN=LB0cH>M9:ZPf##A@c\:Zf)7^JaLT.@FGEH>^Y,Ub3/,QG+C;N:^8]fAc
XG?EZ##08S7[WLa2M2fGD676K/7cKe6EdHIR./Qf@dc]N&J<RfA_IW[ZUR,@AH5[
6_=93,VCX,4#^g(@2(2=b?WVB@e.G.+(g63a:_7D@ef6/fU.)00WKA3T_DBCNFR1
[+-8V<483.Haf47U?C3KKO6L&1XF(+fW)D[bK\D],N\b9.I>g5@@NOUcD7DNY9YG
6gCBgE#S-/I7#J_bA77B;(<=]RQgf);27\=>^TEZB-(DVd]_^Ud0JJgB;B8fXOO_
]G6<^NE>PX+H]1,/A->TQD,)\/#V0B,F9d5L.QYa&Q8CXBW(:&H]@LRPLa3b:6AQ
UEIJ[Y4ZZ43gM0Zg,_D=:f^TSY72N[8=,1+?EN564X<W9Gg?KV9_OG9c&M9g#IJD
I]a1;fF(<Bf]]YN<L;88I?Ydf@8\a\baZCAQ9e=J.^@<:a]SU08(-c,5>Df5>cbT
K1PG=Dg2/0Tc.X.U4O\+Ab\T?O/EKE:/G=2J.V0E-?.7JHcg=HALadc6\QLC/Z7M
a@f470Jc=0dLJDWeH(.IE8cTbS#>CG5[T5+UDAeO2K9HS9FQN1BTT@\?dT_#&1S5
F&Mg]@de2.eV83CXdHSW</?\a./RL(N:;XBK&geF1/9aIL95OS7e7=9DBc&@>G_Y
KNLb6c-=XWN(dO6OF3c5_>V7gY&D>b7^_C<BD??8U:4)_c\>WNNP0J-4d14^A&dC
QMR]+d,17-X;07W,5\-[a\I-WTE&,5?6D[0.B.a&2A[5@K]R<39[b;aU<5\79Z(e
8O_]eP^IQ^9@>4T4Q&@162^N0S[CXSS>]ePbS.^8fE&#,;K@/<;aT-+T9FD7,YC\
8&K=/cCIQHM0.7#0S]NeY=O1)eZ6FS5=_WVbHM;X6N;F7.LRZc5>1?[4Y,(<W#+e
I6V)R/B\H^[S?I#]1//AB^c61IN^K5^R?^4Y861KQbg/EQ&@IUJF+P=eB?K.XOB_
T5>.85Ud_MQ[BMM\W<.9]X3DU064EGW97MZ]JJ,:IFI@MZg1G[R@KQ#ELR#O^dBK
#W)b4@XH7>/R/\J:U52FMSHcNb4#_V<9VC+VDM^0^C(O<WH2N)C+^eM)1EO2T/7E
a(T:Q(,8S<T.SA2,#S7;dN^(d(fERL/K6N><-V4\,L[OQL:;ae0C:a9N\N,72#[S
:3b.#+7)LQ5f:Vd;KN(4#7S6=>A?D-d9\+;aROId,L4FP+JMZR6/QP<<)T(fc3]]
gW?PE58^\CaY1ZQGf5Md3]/\2R8[N0-(JVWd/74JW)6DKX_L.HE&Qg@bIFBS-OCa
Z^-dA(YGQM+c:JO;4S@<FA;#\Q^DAd\-50Qc1VFN]dPU)@JCfN+a9Y85^QVMe271
H_U)Y_U,gc;JV:YMO(?Y+)-J;MDKB;QG=[ZTBbe--SF6Uf;2[V9g==CLC5P,gec-
]VSZLXFTTbX/AP?^I,R/E(,2d0eMV<fYN-@Y\]1LHWLE^5X)>d)E#fCY6-MOW]>I
@;d2+\,-\2^B1R7F1I6:RWM#1[S.&+QNV_F/BfV)W\I<Nf<&=+B@2MVN4+JP^4L&
SKP^ZD#K4#)Nc<2RX1?JNA-&TD^D>XXFHC@>]RDU(>-)KRWW=dGPL;CPeWI/b(P<
G)H6Q2IVf>7bBdU0Q,;.eT\VTQ1OVP8E2gQR<QH-#6LK?J.6@H?Y?-0c.K1BB50)
_<ER56AMOJ4bdM/[Tbe_RI,9c+?&T)@a8+&I:L/?+QL3XLA3JH([Z,c=aA6_12=?
)]]UE,,Vg[8O0LH58I12R0,/>0.L[5QX^^XXBI)<_KW<+LIfG-+#IF<5PD(Ef\23
V56Ca<8f08SBbK#TBd(6Z^@,C[]V80C1[ZRbZO8=aBFbR>#1T/\EdLDQ(JTOXH[>
B1FU2;#g+d\FIQG1L8//fGfGg7^@D&::I;S;^-)T>WSC2K]#L\OT4]8ELF04WEB_
VYQWGBDOf7=,fXES(-T14F+Y1:NA<LJ/Y1[Pa1[TE<11@D_g\WHN7#Jf5aG_G_9(
e:B?=5Z[[IV2,N3BZ017[(_FIO?d/TZ34UK>[4<@5e]13-=VS>R^aTU.CS>&(5Vf
NVRA(KPIZ+[c<#WN^C@#1f5QWB6SXOI1Ia,_4ABU0:Ie+bI^PAHRa^CQe&DK=F:O
8+_;YIV&RMXC@PKe\F&\/0Q=2HHe+H:VKHeEUE1P/SD_]24P5O.c?B3TFE;^^^^;
ZbS6D@B7X7+B;#EZ-a#LX+Cf(M;SWIA85ZAN\@L@22\1bYVZUS2:UGC)dU9A+4aA
BGX-C_^)f4Y^\6.W8b+(#.Y(bVM0TXVS)e2,QQ)V+>?J_K#<A:41-8;OQB@;J39X
J0M:S?LZYaFa\#VJGc)1ESTd5\e2J6WF:BY\K=<<]KbG-JZ@7Z/]_R)+O6<M?LRR
\5_+2TPg7g0_Ve(LO(a@UgDUNKTZ:.TMV;F,NLTQU77>c48S6]7>W/&=^[_)2aOJ
+>Y,Z53f(\C/+a&;&PD#ZRN8;6(VOFAC(6P,:ITJVbW2;?UDZ<:bO4eN&>Z8OGKf
K=A/V_6D>#fNBc_VP/fMDADO,TNM@VLeW24E=@Z)K1_g1:Z,G5ZT?.0\+E8;I)8&
bHaJ?X-JI4CCR<b3b^-aRQ9fU?>CP(PN>F6.LXNc,U&2-#5_&EQ&NBLe]>g-.PNc
)(&M0W3ZO/b(SZO-1A>/=(eaC7WKM?.Ug5dJaB5&_E-O)S].60@cY<W1L(OfY49I
-&,&b[TX0caQ78N>BGcJ#/H;b&J^I[:gZBKAb99e7=bW>FdC-@F73/(JY#@/GI^C
;[>1@IAXA:L/gOTW&UU\=K(RC@g3;Y/26c7C,[4@0KT6FM^\:A8?V)0U+4DAB^,G
Z)(bS5MQAS.HbdbMG\RFBFXI;>A,(Sf^<5#e;MYOEWJ?3KS(Q]Z9>C<>+P;1R_,B
O6bA8D<_Q3.?aEG=S@\Xdad=IN4LbV>:+d=WF_HPR6BIb]:_+A?PSP)A)C-HU1M<
g(>=&H=FP-\8,;dM1@ZZ&OHVdfK4\=O06QX_:X+)(Q_b074ae>a^E,BLI82JT^\F
F6(@cOHT;D<J_#J1#9TAcH40@XJ96Z4B;3VRUeFJCG[HU9B&[46,N\P09?-.P\X@
YTP2Tba(;L\H(eCcM6XAZNR7N;+HA+4NRAgVLIN=fQ1)c1HD:;8-76DQ6-#4I_:?
3a=MU_:HKY]A;M;]9[^=;E#N>AbZ?_D-ANBM1c9:[[F[-Fe@2c1=7L7@)IJ9I5Y@
W8@W;[[S)I\M;_bgQ\\CeWCZ#NfRL3d&MVE[+&AGf.:\OFgM=B^b8K8>I-[_2,IC
3L00F)/R>Ve_7IY/JP#a5cFFZI,<)U=<_XA71<^39b>T6,&D&Q@6\Q/TRg3XR,P,
E\2?g/PD#9B.V-5:L;R],MceUEgAM;3\b[-Pc48228c#PU].1WNB6g&PC5a&UO_T
P)a4S^3TE?a=Y<#>cO[0#VK6Ie0KaB@bd2+[8:X(g1)BaIX-<L^<WaceL/PD<&A)
,PN5YQIAcaACIN>P7&R0/LA_NCH5:LPO>CH5,eM3a:WAQOPQ2+MM+7DA#T7Y=cO0
<7++D_d0L\KSB1Y5\?UKMbU4UN73-dE1-aL57A<ed+.V,@8Ha/dgKTf7W^(APeCZ
Lg\I&<>B6/_O;f6BGUMH_.4G>QUV0CCU87dV]SAddS3Ib_18]d4:VCcXHRK?b(W]
-=d0,CW+O/g2KD9aRNVR^d-.-5Y4E:Vg:IPg6GZ2@Y-?\KD_DLDD6WW\H=4OQbA,
K\.14^H?YFD?[Fe3bLN+3.L?/T4/9BY[TE0X:_N3X#;f/)RN\FCEI-<K+g3)>V8f
9?&[WVB(M=K>KD^:(1^<3:K#99YDgfFACWb5PBQ8<=bK[?VT6=:aUa801&\3GdT9
5V1TE9FO3[R^fgQ4eFZX?FTNc61YNZR@bN:#fZ=\S:H6f+^>-eADdIe@IVQf3T7G
3G[56]<4K<\fg4=^3K#ae2g0f>GDdO&de@#E+g:P=aE/<[VbTOYEWc;-U0/O<?&B
&fF6F,5/.4XI(QHFTeMX@N3;Yd-DQP__/6TIP=NI@2#7D8L<&:;OU1DZM#OT.a)e
YKdCTG]87W+.C72\^=>VAN3d[O5FK:AOd12C<(3MWCS6\(cQ=LF4X_0)-H/Vg3LX
cbLJKRRCCJ=f==dF=1U?><Z52b=PL16cZT@0Eg[L#:3P]?9d]&PHFbZP3KJf8gE3
N?/HGYEE1N(,4TaFPVb]f&I:R9+F[9UEKe2O6-OI#>W//SV9TO9-?WYBZLcU-3Bc
8Z17ZXD)MLVO_,>J>gc);OeJMd3f@SKF>UZ>>\.cOGb@B\@LYg(Z=\+63<Q^5:>H
I:P3\,YT@EK#Q?\6,(@3.A>/LTgTdQf+N0Za4E9;RUFKH+HcR2TNJSXP7dN5IZM#
@=3-RMR2e+5M.4Y-6OS5GVcc017=Y,Nb_7[gA=N_:;BDdc2&&O8e2;L/JR]6.C77
5R9Gd1#=Y@LT<4#)G:LY563\EY/&IJ+SPJ\RJQ^AFC,\N;OU\AWcKZdMZ4\W-X>P
/AR2=HU8a@b==(Zf2aU/.YJ7-Va_PZgLgS&Q[@<MP6EC9UN22HQ9A<De7_Lc0I29
0I#YP;b,(;J)3,e?^>>MfK/P\7=;^Y:a>e8)a4^K-P3025)N/#B])_daTB<dAbSD
_8=YC2F/295](,D=c^),#Y18KB8ZaY-#^71=La/5HJ8aXJ3E#@D[GO^Y:Q.7&^=S
E>&L8VUJ+<^bgZ1QIXc,46?>TK(G9X6KD82,2G?@cd,f&#EX&O^_Jg<RH\@agJI5
b5]1E7[Ee=:X>=?<PMOcXAb_S&DK&^T,-LNE9#86dVI,@-A5;YT2N<Q)F,X.4X^A
CRfM;Y4@c)d=EGKBI<a3FRN?@b)_D^KW8LNfS&ZC/@Z-0CK=-He//LEWT7H(0Q/5
59AXALgYX[CXaC,)#Y&T5/T9JG@N=dD+T,(;eU0;DeFPf0>0Y[7N.&-+9PgA4)e^
,?c(Z-4dN@;2/<.?>H5[d=@TW^A-NXVKCI>QHce,JF&J,/QMMP?1VeQ2?cQ(FJL@
:I-Jg3Z9\N6UdIN.Uf+Ia9]-7/0H@\9973\PSSbf?W=2gMRQ^GGOMPLDZU?S0Ua^
@b4KAJ^((62.d,&ggV5LE)faSe:P\E_ad?ICX1&<;QZ6<=:3,36F.&7U05M=^gXB
D^(2[45AHY.:#533K4/I-aP@e//,;:>?[Q9<(R^^,]0LWF(AVbVZ5@][5SA51;@D
0Be&C#5b[_1_a/[T([5<cG+V:N#SG_(?I.aH2X&9,<d>#@K.=L6=8Y7Dc,>6:B6g
fPKWWKA(@B=-^>A_^0QP.X6D7)C5T)J>e>/\gQUU,gZ_c4aER_eXPO1g4+fTKMe#
3adP_:4]Ig6)JOdHC01gb0Q@_0)[GK0=_\M&/96G+NfU/A0Y.J?1?1JDI->,.ZZ)
g;M>5ML+>H>^\CIV.H[<K,U<e6A;\TcG<#XY11cKG_,\.&W;^\OadCO#eDJ<F-aF
-U(0>)8IMS/Xg\@V.X:JRf)PdW8]WBR2Yb[M&eSWO^eM>.<Rg=D=#S;@/=>[C;P#
TV/NC7gc23=XW/5+4Q3>,\HY0#/HK#6J5K9fCO4bYQbX;5O3_+1>#X,d@NBE2>CQ
:O(68B,H]+3MaIKKS__\I^,I3O0#46PIR[EbSUQ[VO?_>eEG03R3&dF2W)-\X6N2
4F2;ZIT:K3M0DFU8CN@4YGLI=D?YUO\P<?G/,dfOCg^PgON7RP^(9K_a\_@.EgSP
XY47DY;<L1@804^cWZCc7RDM[P&IYgK6.9U2c#IEC,Rg6G/GMIF64HBTW8<1)#cC
8DP\U1+d9<dQ,43VNV4Ge=CMfN/VJ,-\+5#3I;:E-C;<?2(^;/a=DXPe?8BW1/R;
\:eT\Fd^.@F0+PF]8@.2U#@\TS9J>GCDLF,d2V39N=5(A8fKKX14(/M+[K4./AV(
_G_/YfOI;0T9Q6MBXd:&GDUV]Z@76Jb]C85T\0<NA@bGM:O4PO9S[9b<1_?E\BcG
N78UG;PCLJ\9&[?QDBXeF&[_Z@R/=)OY+fgIH)PF=(.@Z:L=M..-/Y\8V=gKHSD<
[;cF6LP<#PE/fN@LNSQC][e]>bJZHU124+?CBY^D2CVfW5Y0X;AT>A;#(^CRAdgD
Vf^7O1W40cVP#3=23g>T>\<dVf^4N[N]IQAa<U^R[fK5:A4TRe7^K,HGT1GM_.aI
;DZL9JO&(E6/R_3Ig8bU.3)=Q&4<P_dESOfa^-N^YX<FAb<^:,f>:OX1<LMBQD+B
PJL)[1?LZJ0KES>3FbEWW0L01;d5[>F0-VNU-BC>A341U#gE-b=_FOS=]X)6?bKN
N6g+CT_aHD5<N?V74M&4X85SO6U^,[+M(E=G1C.Mf<AJ3@9RK0Y,_9Lg7KI7CGAM
E>TbKAD\g:b^S,DYL)8TA9]b+8((PY?V0CK<cfVLB,ES,PC]+&P3BQC@>fR80.@T
7J7YIP3:e3KIgFa23Z;N@T5,LXIRZ#@&]:=X+TB<A?1Z2aI1>N7_MI?#F:K0=32Z
6I+:SWQ-R^bV[S39#^XCg-FA2WaG;KXX?:^gF:@da3;\^G-_>#[IZK[\1\/eJ[Pe
]d>PSFF5GE70c\/Rf;;:+,ACMUL]VfLR_N=ddYRB5Qg\E$
`endprotected
  

`protected
,)8Nc-<S:A@<@Ub]4K4MKID@7GHI#-,)2dF8.W88FO<2KL1/K6=[5).WN6QcKZ2?
SOR[P8T>ADf4O50)MHHVKYD@5$
`endprotected

//vcs_lic_vip_protect
  `protected
Y&JI>AY;7A>@fd?P15f;2P\=MBbVF8:\TgHE8b:OX9b75+#;[_F_6(XdE+dbR=LV
_O<Xf8\MYdIQ:>c+K&5c_[&_-gbTN]fTJ@V7C,QM>H:6P/efC\f)9,N[NOR5_933
7C@#O,(LC.?^\5WP#36^N0)RJ)]L@2O,SL:f5&<fcATd&>CMP.:JXNAVTdJ[c<6V
)[Q^2SS+OT@:JP+[N@>2=/PEW_6e#1#X6NO<U8DFd@+>@LEBTT6PHaDAc?1a8<22
T3IRL4#&bK4O9d][D9Ia3gNLN2VN5\_6?\0ZJ@@V)d6-Rd?a-f/+G0-7H81WN/Z;
Sg#:,]1E3;M\ZdfVSGNa7T@d0JdKN/4P_ZbAS?Fb1MVZ,Nef=5VD#UA@C.<Y1#[B
JX^&1HTOK6TB(b+B@6653<M[1W)BU#4<PNSUT5.T\<+U9dOB;9g-3Kf_cGU]XW/0
N58R09g7\NdX^,?#C^?Wa\Sc)N4,=N.4#7<KF5S.c1L#MeUCA1?Ebb:O_1e]Y/5-
LU?T]DO5Q\aDT7NFGd24<Ha6,_Z41-CJTU+9C@aLA;VV.<L8,TDH[;O65P)<7DfO
1fOWb+S]XGfE5&XF,N,R]S<HN/X+G;0ZT)U2\]K,fT3X17,MDC9O:c[<O/RY.JF>
<aK4#L,H0.L6JQ\SY\S1cZ7EVecN4/)Q@JCQW,b\PXVUJ_U_IF7#gBbY_+L<PK(G
AW<@?+K-eI.>L7,aN(c\F8(7Sc(IWN?1:FE/^OM9S)=<HI<80&g<<:\FIf=#<Y&?
#>7+<&(D#0,e]Y<2AYH,]<J_J=aW=/@^3?9fEB4Z<G7//<H;TO2-e7@[>MLJG0H/
K2e2)&,^e^Vf]D4H/2502#VUHS^2GLAYM;&]YB\D];_C4,I\V[+.,V8([T;<I\Wa
^()^DA;MB:Mcc6:M<eC^Y<:2;S@8N)G?R--,G>BK)Q:I#2FE(;FM6S-=.).SKf(W
OdCO)C5Y>VOEH9MB_M/ca90NCL/Xg5D[UCDN(A:UQCX<5ZeDVA24Ua7)/XB7FXB&
L^2^Od9(;D^?;UF31NE#5D7+ULTUX-DYQae]#&F=-MPP/U#PG\-V1GaHe3>;S\SZ
K^=0JB5^>a/.P]f<WL^L1_fE/aR9H>[JJXcX^cc@[4RA_&g8C3-G,aae>dgP/Q0>
c-&_4SECB3bGW^G+7\8g)WP:VWKc<6JE]eD]AeA54Y#FD)R_/Y7JS9Lb([2.F^.3
d-Cg8N=3-gDZNFLUd7INOZ7&9FeXK;5T(3aQ=ED(Df10e\H<1T+U6S+6AZO^a.Q7
OSQZ.FG4VKN\M+1F9e5W=VV20WA@K=,[e6^1HU8;4PHRJTI]UG/O7D&YVbg[><ZH
FMGCDT-b&5J2?##3d##(0TFAc2K&^?86\>1N5X&;_JW3db:#QdS2eBW8Y7R&):>U
/KUZWB_JPRP.>>JA@7^^BMb0;@/5(/4Ec4KQLFb6?7&cCJ:;^=N_Ae1c,RG>fXLF
@69c9X7&A5IF]4N)c&Hef\K[L(BL_Gc&L4=B57:TcMeWKD:De^QY,E5<gR&39,7K
E)+7H\.BSA<_ZP3MC@8BAE.4Z?eK31/N2MM_.I5DKe9YUJC&DXWK2#(aU5We.\OQ
[-Z^4_e_U,caYH00_BX5BC)&<MGB#QA=^dWP.e(6E(aB25JD8I;Z?_&#Y<_N9Z?R
Ob];QG64P^BE#.<(,O>?/>NWZ5EZAXDfVf,f<I5^YR2<37.73[X-T]8#19d7?3\#
6dGD+A>c>GT^&Ub51[W_-&^fGa^@2:?Q=KWbA6E/-SM:461_[ZI=DQSgag<[0^DW
JaMdQ49ZI_cX&G29Z0LPfO>NHc&C#AFd;7^)ROJ?WEZ#0,RbB_?Bb.ZFC;/Q-7;?
YfDG/^,>C+--c,+c3UXRWBSX.\8<OSS+^4?OWDOM=Q6>1P_24&=\;\Y+4fcL7La0
/=,DRQ-K=CE]-3K/&EGCdM6<AB35W=gF-_b_N6f-C5C&gS3U<EH;PcU6/e&,.D_(
)Eb3.+T=T^9#I&\FC8ILKCB;<a+fDBMJN-FMcNf;J3.3URfe[\[@@D?[KJg5M8X<
#feONK[\?AFWI0=H<HIVZ?Bag94WZ]E?7Y.UYS\WMP2bO[TRd8LMMWWEQ]5g=&@^
:X0Z+?cgP&e^<=S&P+,E3Lg:WU#Y?WY9Ig@e2]+Q-1e5IQU976ORL[#2SO86NRP]
1LZQ9G[H)edJ_(#DW-A[RYFcI(TG\>\DSZI:GPH#;<=B)<X8)6RNE2MHHJ:4[bHK
[KGHKN54d/KdGSSV?=;[Wg+(RWI_ZaJ^=;1KMYcF>FU(>C38B#:7U@]@8-#D-&4U
b6E+>[O^F@7V6#cK@E7.dP/J@</;G646P+V<VbFD1N70-d?E)7bH3b0N.IcS44N)
1UE0(\=I3B56DY(eC^EMXJeF;NGaVWc:7Y((..Kd-=QS(O&F^c@&5I<PUfUD9:1J
3BPLL<T_fb8@)9?/;B\A&9E9O>S=)fQUIaJWOP#UKVQf,RC-IXY8d8^Qf6A?W7_\
<;L=9ID^;^0Q73X/9M[@^(HV+d38=8BH7[^RR(=Y?09KG0DXL&LQ,IM]RCJ+a#_W
U-4\<-SZ08+SQZY>?HP_S?YcQc,]eV,,BD+KS)U<_[[_0c[+_6A..;HJNAe_CK/A
Q@97;;G2BM\G2,/Z,^JGWEYP-CL2&PLZPZ4?0>EgQD6,LbfKP+0JBRBGU/E(D2b^
ZP8OV/BYHT>cbTee^gS:,6X<fD/Y6(D.a^2](T0ED_?F<TN;Nd[]B-cd,BD8\U6@
B&;8=?3U>@__5TJLDJ,F2E3]Q>6c]5X8)D_RCFa9C?<L_<.0a:4(N27d_TO0R,-b
-U(NC]K)AD98T6]?5b]-gAJXV1?BU+.E57L&g@;>E>L:=+S[KZ_9^N=Y+7Q>Z3=7
.1]PBWWg=)5&-R]UY9eNPd)]V]2:GaZcbK#1UV0[BY5_JGf^W#6:A\7HOB.e1Z=3
@?NO^)UUaE2dQZQ-GX)c^I1#Pg;EK&M0V_TA?E[=-TU<:./\TQ--ag+[>e9Y&7W1
K774ef_WTg\=YVR1.Uab_?Z>,:2Sa2_gN(SXN6@?]9-C-M)G\aIR;UST_LcDYD<O
>;dX)a#I@2DPTFK^HE)JFgEU0W@4G+X>5FV\+&6TAR?;gg)DSY7]ET7\3(/JdW@R
=RC?;KfKU81A@6:aPNA9ea/CIX7:b-dQ[VaATP=E8(e-.MVM\c:\E,<Q^.5HIQ6D
,KTRc&C;&-<Ta/5G5,:6-S=e>=IfV^VS+V_G<-TD2RQe5/@+egA<GfR3#SQRW1T[
+e\OW_]4b5K,/_6g7ad\g#5:8BTK+B;:4CQ3?SZVWJT(;F5C<=e(RTP,NBb&AD4U
.BLb-85LW+GTCRTM.D,W(NZ&)6(B5?IZG[3C;gNR\.Z?T<260a98[<R>Fe2dFAD5
1S?YAVZ>M3J?#T+U\0#TX#R,F,U<G,UFY_[Jd&):?3(DDL+D61(JWAK+U=KR(SW\
;BL17ENM]V.FLbSU7f:MF@aD(6PaMVC2B0_VU0W1+>FdDO:Z<.\c<<dSS9c5>7C@
+[P9+F)T#:[],J2-E-(NOL5<AL-+]De<gD<W#ZN()BEE2S\7UE(aTReXI9I[+DaU
Z-R^=F(0^T2g47X<e(\Z)FdNB]=U-O)O7Kc>;eS^?6V6:YSbL)ULXV#+5UNKA8aL
^K?#g[(#Pd#^[)/.@0dHc-ad=HZ;L-YgNS&G#Z+e]LJEE6V<-dOdL>0;692g[OUE
=O:RJV/^T1E2&4XC9.4HEAaVN8H6&0P>Yg6dQA>/@H)/,OIVdFQUXZ=9aMB:gWcZ
,]7++BN;VV1]IS=8M;f&WZ]F?8bP<1#/6cC>>,#AJ=;NHP]:V4gT8KTUHIY^59#@
Z5/E82Kb4d1\@;d1TCc?T5.VaR9].aJR>6[.)6UUYU]DbgX,>)Wf,DP=HdX&68A&
SOR)QQMIDe#-\3(AG@RU;NUNX#NEb:b<\6?VJ&_RF/+?A<(CX>>PdR4Y;I.V586\
S#b:OKb28]66M&Sbf5,:ZHG8^(fXaS_@]@I5/UY>9FYPV_,Yf7)2)b84OY?V<^&/
dA\U;@0[9SAMY]f7KXSXSY80E_1:FQ?XJB9+.g-7BX#@V_&DDP,8-_2]aFOgC0fM
H6\J@.CE;S94_d[+D9&cIa>Da2#JH9(E10&=dNHcYL]A]0;BEHPKG5fG23[Xc7+g
0c:S-C7;K19P[IP?LJ3+;V:H9,7FAgbX,&12VOC7M.RN#58A@bXT^QY^[DOXLAJH
^M(TP+@@d8_,c.ZEP6e?>3.b(8c-S,UD2M7KR8).g6AJg:)/63+^P^>Y=\ON>D]X
CO2R.dS+P8=(-22(>=Z<E<GH)==5G=S;[:be=[e(e2egBQMg\<]c@^/@<NL^9&_U
#3DA,@-0#>RGR.JgT=,]+L4c06X=Pa<]0^RGg4NU_47#TO50Ra(\C(XaT_-_O?,.
S7J)7/H8(P6?Z+DRAI4=K.5XU1JNGJB(@+W@QMK\CTY,=^9SE9G_2=]cU1_a1Ob3
23ZT;I^E9cc)L#0+UP\8b^2-5]TT=gC>OWA&DS9IE9FYKf;E]>M+1KfVbNSNH&<Q
fI_9-BG+OO;Z6;CC^)bHfe+@Q[Q4.:VHT,_N7-GLe\E-Q+.9IC#+;Y=CQ6&RKYWa
9@SYbg#:6\6H+/](\,]dIX4EHP<H2BD45XYSP(QfcdKXf/P^K&E-,QJDMR:RR-NP
VIZ3\<07YT=CAIT8:>^N;.,N&Bb?@c4.3]680b1(L]?0dfOg6/[N9K==^BNE>[-N
V+?eZPWdDXU4f?JDRg^,XV2Ub?Jge3KH@?Y]Pg3DfXJ3da\08@cONd;P+.N(/dUC
96I+GKa<RF)[@FBg756,#8+<X:e3H.#4)G&>?6CX.IGN4[;3b<g8cU]X,GBB<)7S
9&CfODH-0cE\NF;8?cB4]d4eSN@O6]bFJQ-YSb+#\^2-H@YK:_NPN>5OM,\57>:\
ePQZAR&W^\G3BFCTC3?LDgD7AQc/-G,Je]00_;VKICfSNDY?=;4P8fKX<JK9/&EB
8-(Kb+e9f1S/YPP+cNa4>;K_+F/):5EbeHJZ+MW?Gf8A]C((#g&,c0S;6;Y:D[TO
a6eS<e+g2@M:F7VOgdYc.AR,TG_TWE6]^^[AJ;&NH=591711D>RaC34CM2SgWB^N
D8eQ(Zd^IITECLAS8S#8J5B4<a4,dI^<F_U<cXXLLL#8_CdDNOPV-a+&9XR/G95K
\cJ/-BTQ>8F=#K84+[L(U0-1R0;L,2\bC62Q1#G+TMTJ]dL@).:+f(TB4NYBcEU(
H5,UHTEO\G2UC0^/5)COJ6=K7J[:MF<NHT:&T100g+d@eb0K0I&c<eHVFd0AeW@9
M9ZJM=42K2+7S?U/VC14J5bfee#6P&HCgY/bVHgV(EFC#3SBB>]R-;(bP5I6W&6H
SID1&YE-40a7g^R]RY=3LZONFgT4c:I?VK,;I1Y9[DJDD4;P<W3J+D(\P8VDT3@1
MO^JZ[<ETD=FaYY:4d\?dRA12DBIZPUg7[67F1;cHLRH;_(YEa_D=5g0@g^5?a2+
,HR?H+/dP&82=SBL4N>#MZ0a^<K5fF]G&4[N.,2V<J&AOC7S,4WDgT:#E]7:SM[\
@A(7T0<6N9>c5EcW@G,N>@M5=9\C3d:;fO;b,R^KKS284<Q?C?QRX[UN<Q?d[:P&
49Bc6b>^b38MAERKa=[IBB(6YRY+6[)8\[<RQ2>VW>B0WQ]S,.Tb+c&37aL-EM._
3]ZLK;YCd_P_NC.=b;aP.J@2b)e7Y;;,++<#9:&8>;<=N7ZdPDAY#IRX)#/&c3<d
#=24WRBHP(+,DZf\G,.;&;6J?+fWH&\ggFg[1)5d08<ZQ;P^BZVN+S7:63C6H2;:
O-KA4TT3fZ>5H\bLf-fINS3V@\58QJ^8M:HK2^YLGQO6f;AD_SgJ6^Z5FI1,2]c<
gM7-;9]JT9#RJYg[100;0XU:609T2RI7CHeZ,/Wd^M]:KeG_R;1e4?b>FBR6e]Lg
40_CWc.4ZWTW-:78SW0D1QB+bCL+;[)bIADU/7Ag?D]ASPZVaY<a3A)B3AbP(XV(
GA0QUN@d<,0ZBdNN2Y?b?:(Zc17eV\LOKYf)3;aRNgf4WK3YcXZ7eYW]970ZG[N&
AORcO^O_O]9M9GX7[aR5eE(AL4ce:[AYP+Tdd(>990cZ_WM)O^SQHLF=a;:UB?W@
._/Tf3]b(gg=c;TRD;_4^UeZ>0Y6Kb@1?X-]2M[]aGZHX<=eZ(,bT+?..7D1Y3A.
H.65^/>QB\1OE4W(W?,8>Td83NK(B^FV,#_D)3<1fL2=A:UCBHKb.NADQC_^ND)T
_6H.eRg/Q>?Y)2WE]&@7,J_eLAbXTN^AOgQH<05M[J2e:7]>7W90N7.C^:9A:C<S
A[<1ZN_,L8/\R,f2f3+PaIV>._GG,(>fFYe72/NJ@WU_T]<[_H[&6E@.Y^^&eN=;
eS3)DHfYdb=G^\N,7ZD?L.978OEBfQU8JABW]+<OQFaZ?.)4AO4G^:WBOG-P,C0?
I&LLW7R2EO#MFDXD]PVC1,,XC7YSG@3RWM1V>CP5Te0I_7a\&,J#X_eU[(E)IaF@
[LAHO4(S]L-)K1LDD88]?_Z&BBNW+BH\89LQA0\8;I6T0#NaHDbQ+K1>5J<[ZLA_
A^4W1X>RKAL&<AFT\JS5d2#RL&X#6ER3S2eHPV4)eHM9V,D05Tf=[Z.#RZ-d9a;\
b2A1X;-Ed1FMAHg\SO(X3T\gRLe?<:)R^L(S<4;&SDUGPLT0-GQ-\(QZ[)bGc438
N0c@W_1/9aggg>=T)AA23c^DXS?FR-W:&#>c(^U0S6gU>+GR<=WZO;CKT6L+,XL:
IPO7b[b+N1WeLYg)c+T92:0MP@(XZG(+H@?a8SIID&?;FbNEe]IGN:9a1CTHGS)7
?8,RHA59aVN-1R+E6E1L)?\5^(8<g/#fK+a8Vee^PGVF)9gE]_QJ#c):#S0R;f0+
BL^O04IKI/UeZd6:7^T&>^^[?bB))^RGV#EAD\?&?D3>H2>S1VfEB]0KOZ)3?PM=
8P4YFSW;K#Q.B4(eKg1S&NS36F)Y-BIf3G8YRJbKP1K4QXb&OU.B=<,J_1+[\HL(
_FXE]G?O-2MDZNeWd3@>+S?.W^W2M[1TCFQO6<NCHKHUU8T/)cfb(1FFJ]:O4HNK
_aLfIPH&QAUe+]AEZJPS6;ZNAD<?B[9EV94[DbZdE9(+_KJZ>^^8\9R/d>H)28,^
&GK+OF.S;,+&cV_N<ccM/O95=V?e@U7&N/28/^?XK3+,UH1Z\KPDIGLF8=PD8H+9
74Q-T9]Z^#9\R_=?#B]F1SHVf3DJHNQ>QEW)W[8;CEXQKb;O;N=aKeHGBKWRH-T^
1?BRMMC(L-b1/SXFUeA.R@_\<:WI1.>UFDMT61W]6\JR+.><85MRXYEJacG)7#XK
.E9VB#:9];Jc\+P4:(T3CQ(LB1]LTM&B3+JXY2gS:5]LM()FdO_ZW-gPRCCJ?<AR
N6^[LSX>>:6W+cZK7)F->UaW@U>APg&_Q)^e4HZ\]8e]6Hd+VONR336:WG?e2cBU
MH3T^7F+KLOcZd]_S>T-BMT6Z>2/.EKN#,Y&;.df2R0[)2=4EK3=\N3#-Y]EUEB[
]S(ZZP66-@OKU6;LROYRG5PWYCG=1MSS^[)ZT5d6#@][G11C/\+f65]S9IZBHcQ]
c<S<Pc&d,BDg:c)HC,(Ig,0JdL/75dMPf25T=T):UNHH(=XCMBCQH(Cc3JUc><ZW
[>?90E6&Jd^[+W\SD5;EAM.-[8552OWIee85B-Kg2a^-GR>5+LcVR#:P-+R)>1gX
5O_eTa:3-B\/G<#/2UE5:V1_>,c9_4MUcHJ-+NfDF@c9.S67O>)^X_(AMXZ+bTV\
V180^Y2cZ+;LgP6#-5W818:FJUI>6T<c;I?FUZZ[Z(A5-@,c;>dT>CTT+5/8LN0@
9[LaSGNG6ZCDV=&=3<CH)09SC#H^RM>9Z5W<a=KAP;_?SYCG9g;]P]=&.9GT/)>H
e2E,;<e]b57@ICP-9=&26Z+Ug&OOT/G5_KSOHV2^a]Ga1.dS#(12dM:-QMIJ5PU\
][54a6g6&IO+[g6Qcb;Z5QPQ:PJ9JO[^2JE^cP<]J=2;-\8e[4)+cc)24H\Zd/HC
]YF3+SCXQVR#/GcAY4f13RUSJeGPMO76A?g+9SUfP;K[PbFZ_E\RdGM7=3):Tbd6
\JafG=U1MYFQ0F9gR92<)c7YFeBcJd#[[g\+.M+c93)<JEX(<OLScEJUK;H5afO9
^/)+AIQUD8]CXLZSg<6?WSP@B[[YH.^X#W<<<@(Rd4N;[\gJb9/Ha@#ODN^\+OA\
\-A8D3cJGNI<J7572[/g0\4:cQI\c5F9,2<]EFe_:RQYbfF_QR_W9BJe-))FCMgY
a.4XHY?BIaCb8\511d@O]c,YfJTaISF+9P,5I(1BL7QQB/C-K8T,/15=cXIR,NV_
9VA/a)b676L+gW2.##5a\VY6YAI-39VdgH,8/e+H59U\>:?:ge3;X^Yc219/E6._
9c&M;,@LEM&@16G:]52e<IX^2A41gT]><;.XQd<\CB0C/T+]WYbAeC=b)V\BB_-N
67Kf[c7>WNOK+I<0X5IKUE8PU:]HF0(a;ZI\OFM1gVD/_@ZHd^VW]NK>VPN]A6N2
/2/)_@g6YE#deeK6#f9@fB5:8Le/Z99+EeG-1:ZOOUT,4HS0SNd9FFN;TRG\:4;P
<gZ/EcaD0CW.V6>5N#Sb-T>>SQ\W,9_6KV<7&cJ4-FEfU/7g@4DE0FM/:1J)0,08
E>S1Db@326gRf1^_L+)#bD7XB.G5(V2IA-CffI0\FF?SZ\PB37GPE,7cX#5GZDDX
6/PdD)1g2WA.fe>ECgH=QRUa;&<8@K_Q+3A-6#>;^IdHSg?D#U;V]X8\+)K>(D8[
FR-<U-3G;]@.YeV4ZeH>GS@E-7-@4P)M9@+^R[P9L5W+7;4,,J>]@d3]9[YVf-4J
/0AI(+:KbL4Bf_1Y0a#P1-:b7;J,SQfDVRf-J@5d^T68#ZJeB:^3;dcU_8H/?4<<
dfHb6+G><f?RJVad2NQ6U-TVA;O-)X7:/9L1?KDbOc=6VQVa:/+N7KPS<+2bJ@C3
ZG\H^O:WcfBR.47=QS=BLAZ-N?HI[&LOYQf\-S(Z;9e7D/Pe3c1_AC52UR[+Z@IB
)<L<5[B.6-:CFCg^M@J#/+B5038Bd]\cJ])bL5>/13d,4966g^.RfEe/BN0<>=dc
4>9.0+0DEQ,7&>Z:]K7D^R@+[8dJ?R^^5)YcS+[M(G]Q])UI))#6-A[(T(<]<#eM
MS/AT1\9J,_Me0KR;_7>XZe16(J.MO7ZTJM8dI^G]0FMQXRg3@9T&aFf2C?:+T:&
U.7Z\AYM+VIM;+-O^_g/9/H8IKX002_M4RBU:XED927/C:8c=S1Y)Y0c63]P1<R0
[0]5LD4A0bW7ff/QI?Gg[D1?e8#RTL[Sc#@V^/bG,I[XPPdMF/38[BG7^H]0)PDC
@VU;_[_SSd#g3:CH,fK>MPEPeC^B]aQ3(+X?N1RS?SHOWD0>BSIE.R?#:XZ[]J)2
EEFd+[G0K/9R6)8JdC<H<_IH\<bJ+9aJe_)S+9gCbWW\:66CR^HZ68YAa2<K?(7J
1[KO;cA>FTOWU<0,Z2)-N-&4?LOUd;76^aE8]bUJOa.URGC>WF.W65,)-ORa]D/:
@.I;IdD8(RTJ_/-U]C\/BY6[G&HZ>JJ=9P1QYAR9B/,E?Ud1_>4R:KWC78gGQ9ef
\_,.c13fOV:+2:P7P?bYf0K9,(#P^A>)0;,(d1&76K#bg(B6CORH3e_^_Y#[B]Jb
7=DOd^&OC2;gV?0><a8.1c+/a44TEOHVN5dA,BJgWg5PD(-TFCE_]3F(YGR68@>]
7]CS^d?@SSXfYK2ILNH,INRB>N6U3=gaBdAJ[EWO&]6ZHAaW1\-a?(SYA:[aV+]@
R0Vb@#V#H=_J#f4@d:3>K,FA6_>DIID_<C:=[Zd5),G;?>/F#G)E7/A/(SM)f8:&
\^<)Cf8NYbgPe/WB00GY</AOO4^eMUA^2&UJF7_V#P@HAYW>W79?U=9(7&[_OIU.
&Y(.f>:HS_0eK^TO&af<U5=L2MMH,RY^6d8Qd0>6EIFH>A;<?K9]3Zg\B-(UI21)
PWEB];7_\3NXZDZ._E;KL_[9,CKWJ,DUR9RBB5PI.UU6SbJZS#H-(;CX,g,H;9L0
(dZVR@5A(1R](Q5O6>eJX&@B1gF?BEJ5M;OCU(HHCDOg>A@_MS7,Bb)08.LNZ+.L
>=3VE7U22V1;I,dfHUL#W9B9,S:<TRW8G)W/C+I@G;bK&84^16bO-#+V[3;TV04d
H0.S13,b9SgI#b;cO+Q6<E[APb&3B/(:#cGUdQO_QL<>+OYa3/K>;(KfAH\Q^^P6
C.P[XED?>+:[#0;g\_L5H[R/J3\2@<@=4b(B\@d8T+Pb(cBfUDd^)9,g2@a9bfHJ
5XPUXF-)gDIKb@DQC.4CS3@X=GP=AFg;S^NQY+Jfc>GC#Pc4&YE@ZB3J7,4WSV9f
1ER<M0SNF22:KZ6AR.P.?783K8TcTMFc_54#0_IMYKUFJP50.F2Ac-V+VVWA,@fE
G<R\PS^fSGB9^5G)G^Ie26KM:V>RLfddaM&S2_(-H^K#?C)BG(VPRO5=(SFHEbE#
\=S1bcK516Q&=b>TPbF5P/Wb_OF,F0I?,FDe]@/HOYUI]E98C/VFV6-P^)YKEf43
Y&::(S&PHQY#/_/W=1,c,BUJL;57C16U^C#Z3N/7F1)+,T_PQRfLW/9(.P:@,V_@
]FJRBZIQ<V;RA7Q.@9bNC)AAUTYB@Hg=78>>KS-:6RO;;3C&g=>\,Y2#I1^;E_B-
KR6Qa;)#<06WPHN5VZXB.L,6<T(GWX(LM#JGD]V/KZg4^G+YPL^ISU42FRP>6PUY
@?SdR_I(O+Q7FM(-.VWE[WJ/P&].XCN,:42d@Eg@&AE4GJ#RN?(7D<85-)S=IaUR
Y2D>AcGEYQC5)=;6CO@e6S2+0OMbd?d[cN2S+e9PII7&#?K5#U[V^5Cg0F824S+;
S:LGgN)UcD7gI/+dGVE;XYJ#0b&b+EQgPD@4b;9=FRV@^OG#4QPNU=4&61Q3fO(<
5cT3MVYUYdR-fCc_c]^eIdf]\.0[9#B]BU[bGc4YAPb5:DBJFGR.Y:W&c.AMRa<>
JfIK.?49,>-PM8NJ6\[\ZF_Ub60;13DYBX2Z9bc2Me=BNKPeCc(9aFV]XP-03RJ@
P7B@<KHQ3K=B)d=H^d#TM__T&CS3VJF?dRTZ>dWC&Y>DUdOJ[1V[@L)18JO4eV7B
>/8f4;KKI4^eP)J9A8<X79GQ_YXaUfMJK8Kd83]LF#MP/-+GDb:gRd[JVd7X),3L
4_\J=>UE;30P&+?ETZPdN(TGL\F]A0@_P.NTT-)QV9dG01C^e>L7d--Je-+.YI\W
]\d3M6GR:U.YF4fENP)TDWc./=cbB/+RVE8-8^JG@RVPa+4:PLL@<A1448FZRKD-
R[A/ZgD<MX\HJIWN/Q+>[R:)W#JCEQ9WLe,[,g9Re^d_M(K;XLXSY+P.@6g.4TQ.
^.:Q[2;ZZ8c9<AI7Z4EZ[+?_E6Ig?0,N;Ree;;U7J^Z7PG5S&c=DZ@:NC5K6H)T>
@^/JM1?EeK<+-2g=Vf6WHb(a<\S<IB+D9_Z=^6Fc<:ff,^.&=)b.J\+FC,0L?/VD
ZDR1I]H6N)cHF>ab6dB</Sa(Y3Y&[4N::G3H/<I-7P@=6CF,T-.6289_gZYOaVUK
JJMIM)?_SaL=7#3X@f]AB-?8[:dd-<Cf90\2]>]_eF&VYGLEAR1&S222[V)f[H<Y
2]E&>)RRe3aV_0N97<M:6E=IdYP379Q-SM8G;J)T.GR]BQ=KXcGde_WT:XNLH^;M
6)?T=g_gg@V,:CENaZW,(dV,:0L>AP-fY(ZP2a0:dF#7fWBOP<a>1R+2++GVG,81
T8/A&CTE+6LN)GLLYU<J1VTd=F_WK1cYd>.d8T/90:(0KT#_12_TPcLHQ71<FaIQ
RE3SVCea-0[F1V)^(=)P6GgbR\8bWGc5#A3\LS1+5/E(CD[5?>AQ)/L&F&4LTM4B
1B/@V7Lf]B8g(&cBRXAN9cXfX7&@P_dO_4,YQHSfL.&Z,+AT@bB]R@:T.H9[3UC0
T]07&5e3?TPg4>)F.A8(1eFNL+DWQ5&>NDgU9<[;Yg9PNKZIZT@CE6E8OQT;(a;]
d/R,-dK;27HfT/OW;2:Ldd#1VUBURG,1.:Y;4\9O2UaJ,Z>G=R_;#?T_9H<Mf0&U
WI]e#d^g+<H7GN(3FGIaL3W)eZdMJNg)=M,)HBUNGZa5gBK(&9e:)EC61Z<5KZE>
>CH.c?9/(2056NP^=<0a(7Vf:RYROSaYTf&g=TJEg9L=+4N8>-KfO+ZCOF/M)2.f
Y,]&5)A[ed>8@fM9fJF3>=)dQebbKF+>H<S]LV,R(L_H^&P^3>=(T30YU](3RJ,?
Se@[/a=84\I.3M.G1PRA&BHBY1]QCU9gUJH:/+>_3P,(TTSf(ZD2#2/UD.d=Da(G
e94J2Q&52(=T,_gV==RX^]&/a4cA0+]_>F\.#HL:dZ+Q>F8SY^W96<b/ZX-cKS3g
^a[;B@If0#@\N5H45S?Q^d#D,a;(>S.:\-MN;\ITH^a(COG,?/=dZS+F\>_;=/S)
L?-K/9/NbdJd+bRb1e)=?(E,f[aY(T5@MU>6?.2D3YMK1;7[62R^g-.PO)e?O/2G
&\4IGM(UZ@MaT[31Cb,(M2LL235P&B(Z5-LTREZ(/.@KG640-T[[=Y/0Ag/U[:4\
)G7IE;WEUQE9Wg^UXHg?:N&#a6N>9W,7:dH6RDbF+AF<:R43V3>08W82gOL,_\Ca
;0Ee9_D?<B.>.;N5HQ#[D,##@bGEcKZg.TZ[Wc4=5DW&>]JVcZ)dEa;M(PCAREZe
2XeO1=ML[.JKEL[?=PT))bFa3/V3<6-<UC<LdIILD.OLb_W,:4Zb,&9+_7/(:T2L
a,#QJFYR3[]90fZKKGQ5TC4P0K@I&MaN74EO0[SAd^7b?0e,GAL;/U9?1]O[BUY,
VF8^a.0ZdO_f?X)7.cM>Yd:GPBQ6CBP^WB.KMW(a)(BMLF5V4ZJY473>G9&YWKb9
.RIXL=gWPb&1RV]-,>05HS8:Rb]HH36S/?UZe>gH(eWQMBd#2MQA>OG:Q))ND,FH
dZD2H3=GS;5BM,&0gbbZ0g9.SUVEeX=ecdTQ&X#CeeMN/5QN.:,1UO+b9R(Ec1B-
/=b7Ae.VWL\DG+GI3JAU,P#:LP2H3UVcBf0RR[ee5]_\IS\]&ZD5\9QD5&U\g4df
WcHR1;4;&OYS^87X,ZDLO4(&f#ZJLT[9OP\ZH/>c4UI&XOTC=:dWF78W^DYWN2C]
XcbLPFVJW^feM/5;&[;:=?5=MbUBI)f6#_d,CU)O+NTL]V3.HH)YXfbB\:e?MQ-W
B\U&5Q?-8a_c7@Q941-1H](\CRMTO37_+Y/&4\.JCDS>J:7QBK322SVDc]B?=6(G
>+V:eAe.A-MJ[VMQD>6Z=>M1R]MDGG>^eg44M:6+T;8b&PJASZ)I+H7D.;KaTV[3
?,05(XQ:LB7--D[,.::C.8DWK+W_3?1bM+A]&aMB1Pc])W]\8/PTdM]dY5H;eK.[
1ZN=K&MNYQ7+ZE/3_81[N4IVaBNVcT1)A[Q:Y;19I5:Bda&O,@?65?[..9/GV=(@
;\<I34;_1I56aAXf_/J[E)0_/;NY-g=-^H_;=?(,f&?-+^K[>>B2&@Gcf67IO(.3
dc[X;PSBRAY0@UaaET]7<B9dW==LTBKODKXB3c8WK.V6aB/gC#.Q[&CA0Ec0]VV6
69PB1,LG_(/Z(F&9HS^<,8>f19Tc3]a3ZT<R7VF=eW_O9F]4GL):Y(GVVOKS8J_L
bZP3Pe]N2N?g_SXIK@b?@CDO\.B?ASRR69N_1/^F18+a[=b0G+5D\gZa[[g<L#T[
9(89[:3f5_]8]cB<e^b-/5ITX]dHd.4WUH3[7WP8.;K9:S@54_YeON:(:A+5W7.W
1YHPN:c7c/SA@2/7f]7Bb6V<+/OZ)=AQg^aPE3<+X>b=LPX-HP^HdA.g(^CU2L&?
@b4WE#_fZ36OZI&LF65#Y&GLdRe2U70)Xg\U0#KP(=].3S].(@(g(.1@:eYD4.Y3
.0GV(9#MM4U#@-1eQ46.AEY)QM@W7GCJ9:S5@[8-f>I,E:4#c)=UH@O:M6_AY(d^
EV,7c+4f,+S)CWABH2Z4CV_.YZ4+-U2=/Te-/E8A/+V:]>TIT1N(dW\=_RZH48gW
AB@(=;/EP#?74?C2]MJ^J\e3+T9H06T2[(#U[T-c;TQ7PERDeZWXaXE^<J<JQe_g
fd0dT_VJDG3g8RZ#UFdV;D=^gN<a/LgKD6V;.ED#LVJYH[aT:DI^LIT-711N-^Oa
<;Hd4>GXH=[^fe#:SW[X18]L3_F682gC<4J9&c?#;G?/W1/aTK?94ge8>6ZO0:e+
EXea\INH#3NL1EG<6P.4,7@cPL(AK.UUO6gT+>(24FY6F(gD1AQTCINOT-32HB-A
(?D))Q.J8WN@a]dU];dM?NO4(=W&#ZP8R?@0e+D;I]a@/\-4==(B;-Lg^L8(c@S>
<+K[-XD=5LAc2eQ[R(#ET-KDUW<]OK,fX>T?:UUf.6]:9,Z-1M?GNdU9D4-#<REX
C8W2.,\eDd>_aFST#)_Y+5>3Y8P#d)IM#7FX\@;L@JO346=/U.B>)ZbPR(f9=88@
/fUT#-FB(SJ4S8L#E[;:R7LFWdN2K^9)Z2]GdJ2cKNS-E&CYNKFPU)JXc[cE;d_U
cAX)U1&#SfTFIMI;+3L?1A250E+VaaE21RV24UZXcHfU)6M>b-+1.AJe3_(VAXKK
b//Q+Q0/?+HFG#YUY>>CM?C92D>/5@2\Eb(YQ0W?BK\4@R?643>?cg;6O_R@DSU6
g76W4X#B\UTO[Ag>1E0-TG<b=^=SM)3)bXR#/>YS7U,Q;^]g<)A98@&RDKP(HN)K
Qf]<R@61DZ6d_52PCTfHYWIB:71(Ge+#Fc6FX4e@eg:^gSLMVd\,9365<H>S74#V
A:9ZL[)71SLB:@U[]=,Q67D>>+<Sa<:SAI=L#_Kc=_LbU1/cXGd&=Z:6SJ?&,9].
AdQa+b0eMa@A=_[Bd)]20Vfga:X?Y(XX-:S^J_)eZLOb/bZ\?GSc;2.,HPIJUJ+C
==F^0b6=<K.JJ6]eZ6.5KgeEb)&:-S9NWP>/;&MNW?GaW8Hed,<cQYK+>gV;Z.L2
Ag6JU@G&aJFb/\62\a8aIQ6NK]59X<0,<[1g2_)\KGU+WfSR]TOOOE>DV6[OaY_;
I1_+@QI;1B9\fbfFD5VW,(MGX7C0eBbG5^V=7=2&<W0523WU/RA@+,A6/#Uf=;;L
dW4,CC(;I1BUE),=8gQ=SXSQA@a#ZSdK#=2M28+I@NWO2.DDIG,/01..U+P849;)
8(XBdWP2=>5K++)CF\^/)YKI?Pe:N=G_>W.-BgQM(PaT+F&JREM7ReFJ>DAC5RHA
7[RdI(IG.117,_A-;J[@-TFK4M.;f/10UN9VL6(8,Ze>3&L,6(;c+a9TP<ccM3X[
N=+;Sg\(53T@?;a^DF-I9O54DC37R53W<E<79[aM6=RT]5NP)ga32G&D^^QH9,[,
W=/XF;K#NaJ<Sd@OSBMRJ@S]IV>LZZ#)CecMP24e?X^(INMC\e>(:HRc744P3E].
b=7M:Y>C_#<GYQUGNd<M?RYEVd1VQG+AJ4]OFUBG@V>3_6fIVg0aaOZGaUH&L[QG
==;P-O-S5F90g2)eREdEQ;>U(/]c]KgS#e)J>a/6NGL[DJ8XU@N_+Z+E_(8UI9KS
T=Jc.?YELBdePU5TO:?;NMW[V0(:&)JK[KA&7@.PDEA[cP-;5)V/YR[L#9A=a<PO
1CgeW/[.I;OTF9D4@@1?6EMVZZ](Y:2CgK^&:07<J1/[?(CbT&BWP)B+OQ6P_eID
@I>\R2_g8G#H&a6)(([g#/6;]Y^gT1>?=CH2O+44cVM[(R7?1Q3QfR?QE8a;aJ?b
\:cC:;ZNOdGW-V//N42+d&cJT=1bOO6d4a[NgF4Z<Z^^8[P_PQa;/;9;PTLT&ESa
M^VG]g[A,b978]D:ZA.O<_>N@E2WN_&URGf,:EXgaF8gH)D^^[ET^9Tf[\@(4L5g
,3.+CH8DSAW\;2-g57#d1@g:CKVC8aK+;C=L,,Pa-<((QD.W+=[gC.&_;S<c.aK?
3E/17BIYb?,E2>AL\/bJV=aLUD_,IAf+Hfa33:ZOTSLaQ8T(HOB[O6N@-B^H\YZd
&J5HT>e@Y87P?GgVW[Z[M&G3@N9\PIe#&ESZ(6;[,190=Q[GN(AA>=1-c)Tc4>+c
6\MHD0U,:4<#VFfSVea\+YU&50FRe6e(<)a3/fK^<6K@&@7DLXY^)ba\,::HdWN9
9:YI4IN#J4]39=P+?DDgSf^aB>6eQ(5&^fG+JR.-H8FJb(AGQg2D>PXI7471EIN:
g0_LQf#\JaG=c>D<BYV=.X.&;d3O=#c4-[#,e]LV>+I20B5Hd0^CEJA64-3bC\:^
X_7X:KY24NHbG-N]g?YBg]@,?:6fcJ](>a&9=KSS@YQ+@Y1KL9+]5f)DbJ4N5>Nc
cgQ39OGa:LaJ\>c.R(\dRO5PAfS+Z85-N#.dJT7X[bP):H.&=W3Y7_]IL>VK<9MQ
)T_97=[XXYXYe=/I?D]+_/ULW@cQUX=g?[MU+#DP(bG>TeKB8#+a]_Z=NF)K.=&_
AFX2EL(.<.(D)d/+;]Y]X1L<NfX>6LPT;=,-DT2PbA&&6e<.=ZH3/<dU)g_FDEFH
>ND8,L;[3fGY5?3>=BGGDIF9D^eJT/B+g8a2TWU=N,O>3,X[6TF<U:2K9]BB63GS
V84J_-O0a)1=PRe/c2+;D-H,gYc-Ed^JG@OgY5(AG]<H9;_gIOJGY9b:3S_Yc<(g
bY.&:Q3,O4]8NNfa_>J7M9G5>\P+^I0g#]7AK]@C3BM#cNaM]H2O;Aa3c1TO^,cf
g_9SN^[;[gg)5Te(-/_f1KB=&M[D1U4FaK8Sd5@R035I^da=aa?WW(d1Y?D75&-]
0U<B#-276;-f_6aVN[A9B6+R1GH_W](Z6:K5.LO-W<+,C7ae_D\@V7V=;?BQeg#P
fYQK6gf=TWH>VJHD&)^eaC41U.\?E[g//80dJKI&8\5QA9d.R6Q=T;e<bV(OP\93
TagBA5R:ILb(C,g^@:3AdIPc8^2=@ISSKEBYX+JRAKT)a:K:]4L]S48^>_S=eY3a
f+<7(,\8a/a(2M(FI8WH.9<R:/GL=MeaO>e)64B&<)]cOKd5]^=e37.^Q#3XC65+
Z;Y.P;,)<M:I.YZ8,L;J8-UHG&PYfa1DXW>W_8NfJ&MBH](.ZKWe,WL&U3ScEH/5
M+XR1&OSVVA^Q-0AW9VOD#R.d(9_3#a&g5/c^1(Rc+2f/2XbKc#HIH=-@6Y;V.3W
9Z84,O93R(c)/Y@c(1AOdEUEMeR;0cQCVUSR//^7\9R3#9SAWZdBa^5Y6:^@3TN&
0NK#?C4D;G(,\95[Q+4:2FT7A\^fZ9c1Z4;W8[Q52g0]XfgA(V8@(Qe=LFaH\M/1
;[(MIbK4e=_Gb+=Z36g37W+8)E&)?6C5N6A0IHaO0+BP;&58+Ac+GY:=+gN3=/eU
fK(g\Ee=1^a=HZGR>^<52+S.L^Z_UdOPc]44LB7N0a+IEE1-XL5)HF_X,+H\3466
Q,R4CV9+8\1A:NY?#HM7gMeU7(bM=&Zf0Kb[eY@9896Y2D1)C/HEL8V8<[Lfag1=
60W.-f0PaP72T7;c@<Z)&@&L.SdSN2@=c6GeO&BDN[5f-55g6MTY_WDKE<F)AV8g
^F_@01&@4,)_HV7UAC>3W^V^XZe<KTgdC>QUR:]/79=96.R,FaHH.5ADM;V9CXLL
0IS,1/F[F&b5SP@dSD6g;Ad>d^W[@?>9A97YcE-0YJ+EX:;8EGZ)D(A3RGPLY^>T
]7/5a;^91;S3;N)=b^00+?^1<Ff^gR(R?[,:TUV:#W[b/SG+/@Adc3:;c.:Gag7L
/gE=CecED5(>@56a;V,=6._g><S)adX,G-H_8XZgMY6?5^@FCX&aPV;[[fd)RgJ\
@>1[bI1Fb[7\/GMcYI;X45@0Kag4P&2E-\eB&=TV7INVg+C6d9MfWbd(-5X5W2=I
5WI0gUbMM>+2ST(6:KIY?]SKD5]d1&N\6GEC=b<,XTO+9,f^[F[)O5+4E8B\8[\,
GOIP:JE/2#]BH\-e(a#E1=K?9HBV-2T,-\0T[NQX_&5Q9g8T4B/N<L:U8c#G.)[A
4TA5eE2MWJ4ND;^47+dI\RU#\6Q&.V10bL;Z]=N9.]L[dg6BAPe<9G^\YQ^Z)SOD
fF9X/:UW7INWQC5ABNCNNK]WAGZSD:4[EH;_/@aUK<]4]#K_44H0<X7FBE9K]0RT
)IVRR2UJ?]eL.2Tc9dcP)...7-))JdYdJ<->AI9bLZF&QEcc3.PU)QaB7>g/&J7E
C+/N#a\J]2X>f8X)cGHVS>:)L,=>47U?22:GXT;+F2O<Q&Df[HZ[OQ\3+\\[#ce(
(eBKd-6=4VJ:FeXAfd\Zf69E<a3XH47#:T&c+RXZg6S7c?S-UGfPQU#X#/;cc6@K
0HV\1I3;bY,2=,]3&BYJBCg]>g=#-7+QAHQ)1:MO,6?>9I4Yg8&9d0;K_H)9WHV5
X@CL9[0_gXb4L7a(\0(V(BY1,A^JBL+?O;?_Z1#89dF?FI^0/?9?05:L1/W[M.e[
>)KJ7VcP_>0)BMSdRP5J@LFG_&d;+/&B12cD&Y+WULa98=[ZCKV23P11G,bR/@>?
4\/IHKX/BCgGS?<^WTJVJgT?>a2I?J1NX8V[MI9DJY)J&RM,0S6#-V>EOQ)9V=O7
[)W5JQ9OA.XK1<F//HFXU86:WZF>@+Q4KN+;R60d_F9[;5T<8BM8eOB=77_L18b5
+\S:7.d2O/^7(1NEM6-54eSJa+<SJERVeL<7@;TJV9K(9NE7)&Ze;6fRHTEX=C-X
H<bd9]=Lc8Zf4[@8VD#Og_?:e5H[0<3(e^.BKT,F7GD9RM5(;Q8S-\Y>U\ZB;cSG
358cXEV^@R2VdcF@f;fQG\=.3#,9@R;K5L8_,K06UU_H;dZR4XUB,,=E:=VD2UA-
6=I>Z.;WD#WU12>5?NBDM=I^@0dcGC:T-Zf3f1\Me\YSEI[GM]Pa;?VC1fT6G_(K
S0HX-CQ)9SU,<-g\DX44gQCH)8IU<.7W;D_3ST[W7]^a37(UXc.eZATICI_3JHg<
/5;5N1+O^NVRN1,e>@#;e>C#G<Bb;0<(4GO:Jd4Q#/Y(6e9g,TWBMg<7)++WQ8F1
=SLU,O78K4FgfQP09Q=<WVB]8]]DP=DF/Q_Rbc-76UcGf+,YM2Zc7?0(d_-\#d1M
&;N;\;TK0R=#D)5Ff<>B+(fPdAI@?Q+>==Vc/gRQb?ZT@3NZNBS\7.R78QcaJ(W<
Z?F]&#OM[@f,\eG[.Q)QAcPYPJA;Gg1IJ=59KLY?2BPX3>6GZH-]&J:[\fBP:LUB
dHc+gMX@8=b8+\&3RLEE_K0fOF43)9I.YPLN-)b-N6;8V;H?VM<W(9NKg\E:8C.e
OABYZ^M@7GHHF-F>.8T;2@532V=dA=c;Z&4,R[?J417[:N#V,T??_T/[10?O@/,G
I\-09A@VV=KA\?6:IPNK,C;>AL(c?7?MFT,</XeKfO48)J:d;L_IgUM/E;K>N<5/
LKJ4G2;5;U.aUNd78(d;M97[.QF];(dg[,F6@a#VaecPQ\UL/0IW(E[gE.>e4d:-
FeCT8DF\>OKE=1K,#621C/-@)5G.):gQD)_-EP.^DFZ9>QSQ7TFQ7(R,E+RdE]9/
=DPW>f\0:?P76CgE-V73M6XX@eLU?MeP0,4CUR46/:7Ce?N7^7#N3MO],>O<&a1S
70MLc4WUY;3EL#;(^7Pd_]].feW][OJHREP-CUIc.AC767.Fc]^3/Ad5WP(;O+db
e&T5W&[dcXE[)IcgS>W0VB]Z2a9>CZNR6#Z:1Q+.=E2OgQ(2#NSL^<CaW76\:56-
#B&W#/3fOTJAE&LEcRa(8<)&GPZ1LK9U(H[W4[(T2VTZ\^HJQX)E;E]4GD?M.N6G
]Fe9VL3K\_3/1Ec=O68NL:_L3-Z^N<N]g-C4(CA.P@MT&cgNLWRRK1\N:c0+Y)&:
Z#5f]53E>0[\)76G5L@b/N1Of2E4.W0/UAPa_B;S>:CJ52=1.2.G<a;IHRRT#b1^
.e\fbODTR1^-:B,^-cUSQV<M[F@F^aE\@A#LLVL3gM=.O;O.7OU+F.DH[aE8I8<B
=#IGR4\20,G&U>bb^F=V7#JdZ<cSG>P^-Md#cLS_P;7bD..dZM1AD]F9:T[P4@?E
Y/H6V00f=A-3,gB:?<b2^:_AV2EQGVL(0FR9SU@HM4^0PDT.ZNQ_?\-UQ;EZXQ/^
:G5A5;O:;0U?FgXc/R>?C/:[/Yb3N-70f[Ygc]HV5(6]gN_]5U-a-34Ga]FX>FH\
C2CGRb.I#5OaIFCg9OE.\FaMCQ6S=YJ5.]TC&_:0Db7L4d^&>1LZADe0J/AGH2X<
FV3K+QOg^?IFL)RIX(_MVVO&b5L&Q/ZQ_daC[G#A6\,[b#LHC=6T;),RaD=FBcQ@
XA:[KPc8:__.7-5gQKfS75.NScaH.QOJOaUV3P>US#X.WQKA6B:3.O@.DW,fHgBR
85-[IWCUV_gC3g@YP34L4Rb56d=Ud(PfagcKJ&<<f^JFgcEM^SbL1^RX/J4GZfYX
/)F5ZI#[R-^:#dY8#KOW;=T2a;:S(QD)Q3V-H&PHCa):Z\6:>f&0^c)TXNO41=6R
D14+S:[[aH>N\][<V,3Q.a(Q&WH()C(>/_FbMR[Gd]G&:d)e2ND\WE:#H^E>cM5M
93\?b?6>0TDQANM@fELLL,11^<X@A0Z8RQ99f137HG>I?b/Q&YI+-LAAGRf^5F-6
YW_Y)4&a/C18^,R,VO3^PeAaJ\QdTQ-VSQNQ>[be-8]C-HP&c+^T4F=YM&^ARS4=
g50Z3Z)4+/&C0DA(PRe4YWD6;Z#W^<3-MFIV2CLL-?V^:+01_D?b^C6VG(D@-R9J
TZ;;9N)1LJNB>Q^MEZ6&g4aO<#]0Q]<8Y,YK]R/:DKVO5&,M90XA<2)>HYW9:6?/
ZXgRDMf5.=QJf_OS<0L?N2HDg>PLYU[KQ@bLd0WO]?YE^Z#S9,@W]M-Q7Z1VK\a^
=<@SM\^@eAaY(=+1TD^AZD(AL]eOTEXd]=&(V#-W4HLX_KH,^0He\TJ@<:08(@>]
\X0&P-eAc^7/RRKCL+C^2b@<7^KWWD@&OI\aT\CV3f_&ggN>[&4Z#U/fB3L2Eg8M
/JU))-U_IH[MfQ4<ZQG;U?MW/_US.PCaM1P8G/IBA#Abg3)VULK1)G77eTd?68O2
-De0Z]1;#^b)9Kb&=929c>FdcAKg-?PR0d:21A)fXU;M2d+WLEA@X#P7Z=269bVd
W7fQ,M#[gLc]&HJ=GJK_9B0V^9Q^5>c0N(?#5_H6QQV>#;3f51\S8QTa><.&X8DG
&<8=LUR<A22adLR:80/RRZe6:\_7a:2F.W]_bD;5LF@)LVBW7-<d5P_F8E5[gfN7
LB08UOO,[6_UGW2c_4OA#,f?GA4RW6QbEe#8XH?.RGd>-3V;0^Q91M@;+Ea/H\8O
3Re=1F#af/6Z)_QH\cd]B&e9H0HX,01_8H.cJ:9<(YSK8&.&O87<DIK?3C/3T0Z@
18N,/&Td30AP,9)DA0QeO]OcCG8+2,)VVdc[Ed_f.TaN9E+]J1Eff5A&<Q:5CB_e
_/+Z.@YIKJ&Tca,f9FRZ]6M=@U#@6b,f13eWGW]Z:BaKJJA-ba<IV3J@d_(UF)HW
8:P.@,_V,K7]5PK;KIf<DILQQ1g.X;SO&7@=J7>?43XRG.Ta5N<?X@.OcYFTD+\F
^TeO)<,5^ed3DPPY07\PGGBG4ZVFf.T/[]_X>4E/1fT>)(](T[@\(f]435eLDd-N
#@9#M<;DQ^bb=c5R]_((Je@a].g\SRbBFRQ@F6AB0F/G=Fd/5YOJ4J-L/ENaD2H4
&,Y_NNX,99;;V7Ac?+DVbDaWA53O<^eC;4WU?TTb;T=)&\:6RUG3^edE[ALPXJ1<
,[f916OL1.[JCZ3NOHXC-H1B//]T]+Xd^B^N=E\K6^E)5d[XT5d1PSS?c2.-UE;X
WSSQ@3AF0WLBCc54H1BR7f1+,ae=DDXJMd.)CWMSMVZT8S<#0R)FGLRI&S<;MQDN
dHg\@<&a;#B+05?J3PY<)6c7fK#gUec2JD]COW7T5;<;CXO7AT#gUVH/WUAL+K,4
]-U&1CFX;KL4ONO>,9M[.BGVP>NNb3aGL(@5](=UCeMY6Q-R,<D;5S\g7#cW4c)a
\5O;ad9900I[^Bf6f&M0FfDNH7(#5(;GK51XBbWJ7e/]UNcB+>O_#A5Ag(/FCKdO
:1cH7gZbQ.I(9e=8->.AE]B/FS0I<=>#K[=P)N[@EJ#>XW?@H2B\g@L?2D3X(B/_
?=&6Y8+R1LA2[\])F<gO?7D#Bg;VJV6[#.U8L<IHBA_c/>7A69,;I;)-;9EU1IRK
S1?5EQ5RK<_fC9.4M0O0=Dga__TS]-:X=L&BG;d1RZ:U+29C(VF;S52,RV:L^TJ5
#@86Y<ee4WM4-2)E4I9BX5+J(Rb>_<TY:GCU=Yd^&@U#94e\BM_0PKJZ5;G&Y5Rg
/6ZYdNXE/BBHfKGVZ&+0?Dd=QX6G;LE;Re>_(,6e)Y6:8-X)^(>:WDWH,/&(B[R<
EcJRf(I/WU:KD^P5VYGTdH>-=^(XW;VcS4S&[.KN9>]99]QY?cI3E:_(H_1>P#8H
]QFKN2/K.=\,_0a]OQ7(MBB:D,699fI,^=dB<#a/T^VT,_DL8C0d<C@dH=;4dS##
]b<=W#2;FR]K]&97ZR(S3H&dHC@C.M@9GQC<<0W-I?M\:=C>G,0N;^_eA?O(T<][
4,,N;C:\7K6-4\8[37L2fL4Y70^+H;(cd9E6HfCPOH@Zd6.LMA]3eVQU:T[\?_82
.O=,=O2eI-e].7@,7;8PZ4=).N[Q?05a-2ZHYQ;H]J\B_8f+D,>ZDTOS.#M1>2ag
2O>?TMHX+:-WO3H8BS1?/Yf\H@e6SDM)@#TeWAgfY/VU90:&91D=]Wg=MM;]Q0BK
._/9D,4T^e:\ET#eI7G>LP;3IB)CNV1/9_[\PdQU)0W[Q&Z_]2T4L/4M.[_B_cE-
B]8S73G2/6<VbVKJ&+2TR?bcY1^HGE@I=77OJZDQXWH#:/P9,?DO[C8;A4,I/F,O
KF4PAEX_gNgE4>]=NO69:XUfH;g#G\<OANHH#1Z^+=;:E1Z@&L6\&:&f\&GbV4=(S$
`endprotected


`endif // GUARD_SVT_AXI_SYSTEM_ENV_SV
