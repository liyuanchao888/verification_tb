
`ifndef GUARD_SVT_AXI_MASTER_CALLBACK_SV
`define GUARD_SVT_AXI_MASTER_CALLBACK_SV

/**
  *  Master callback class contains the callback methods called by the master component.
  */
`ifdef SVT_UVM_TECHNOLOGY
class svt_axi_master_callback extends svt_uvm_callback;
`elsif SVT_OVM_TECHNOLOGY
class svt_axi_master_callback extends svt_ovm_callback;
`else
class svt_axi_master_callback extends svt_xactor_callbacks;
`endif

  //----------------------------------------------------------------------------
  /** CONSTUCTOR: Create a new callback instance */
`ifndef SVT_VMM_TECHNOLOGY
  extern function new(string name = "svt_axi_master_callback");
`else
  extern function new();
`endif

  //----------------------------------------------------------------------------
  //vcs_vip_protect
  `protected
GgbfYYec78&1)0/Z;N1?T=[^8D)2EF3K:D#ceI>Xf0]_5a)d6d<T)(>5WXb=S080
;KCe\+Ydb&6D#Xga:YM>L@A<K?f72CUdP)?AL<aU9gF;C<]Xe&:M5,-Zb(cX+_()
1OeE:][Ic1_a,F>fR<UNC:G)1,7DeHX6HeS4I?L-0QbE->SBZ&X86Wb8#IO5X#d3
OWID1e1)Y\9RA>PFX5NdG/)^S.^OOSWeF^E#8eGQ5cS:::?F1K3N\WI3?=CV1><1
E2]dDbbL.T4=&KTZRK=YYF3EgEW+J5Z@=/bE:3/7Ga-=9;@,d,SVg0UXOY&]@AEV
^bDN==_cZ/CHC-A3XCc><B7@G6]+@@D:@WI?I3.V6R5g76C](TgIeUFZ^]S1_YNg
6V^#d7e-N0b9/fR0&VF.gCb9SXcdS+)dIA24LH^K2bT9\WXEfT0KMQDI+]#;W@?_
=3cWTH5D9E8Vd-\M9OVR;#2&<C,AJf6>AD:;QH0_Z:L5[[4.2U\fbXKFR#9I818e
HX[=ScMEB#2-N2H\005UGC:#E:AU,V-HTHDS8V0,B_+(CS+.^[GWM>B/\U.3&&J#
B#QL\/00..1?eOI9>.U9[)8d9e>=X&.5f9X/T\AS>E_9X1a#/BK[E81\e]CP/B7F
F9ABS8#K-(:B6[cDO5_S62d;JUQH/I2+THW@ILHWaS_SaT0Z,Q1=[&42/(IMHQON
/>+K:P2CUgVfVd^f-49WR(aeP,OM+=Z(Zd7ID\cD[10.-=F0SDYa:5,NY([N?cKD
8T:_^]9&<3?#fAaFO;Mf90?=Q1[CJJ18::I#aQ<;PE4V4RL:b?X:bcZ3^ZdTf<;#
V@0,I\>1)/GF(RIZ=a4&?0]M(fM<-c,8\aLHVQd:/ZNYZ(F6O<4]][XT_(C_dJ-a
3QFDSME@8,)([Z5NLVe)S4.SdQZ6-NQDJ<g4(d.MfAW_/5E3F\.PU7C;VUND4K1]
OZP0g:5<)e>Nb/-#VHab,8=_L]V7>)RaO5<b,G6\T0f.F_#-(F&#^YIRUS/)X.fA
RL8M,J=fBA6N(a0LQ:UZ?9aE+9JG2Vf2?8#02U2:5B<2)\-DKF#9,&9)YBVLaT..
AL=_9;T/;bBV[J?D22TFeOV^>JZSJ@;(PLNXC^/MY>@BI.T0NO6QOTUX/M#[<\dK
L0bOb4-L)/d0GXL7D2dA-4B(5W(BI:f+5?ae(#^KOZ[d);PaBI2He#(+HVf;MS;D
]-._bffK\J9Y;U0._S3eS_&DaYHNF7ffE@/8^+>-W,C)OFIdM_+[=UaG\2Q6Gc+_
DGB&N<9?]<-=JXG)_UX4GM_GRgc#.@LCSKgXQ68]WQZOK0#Pd+2N)E&XT,J>XSIG
@WN1NMPMb=fE<T?e,dL&:X>1VR#\f/a3[1W#X(KM>5QNZVF[\Cf>(?GAK(4LWdK^
:L^].#b4#aWS/PR)])DF9A9UC6H+_O&?ZQPBUcAcT5c.&+\R2^H++Rd(0gC6KH+I
C+[c<QM_C\50\V[+_RIOPXeS9KXWP5N16?c#&fJ9bE7g@@X.:b)8F&3X0-VLeXQK
LVQ9<-H65;7aNbA4WT;78?WfR#fX<3-Y(KG]-ee343fO?B4FLL4d0Y8f6PU^NdI^
R;^ePeKLBZMVf8GCMPYO=:6Y;O-XYfSXd,TM(#500>6UL-<34Sf7Z?_b#@32H^,#
JQF5cdb,_JNXf+e:/gQKeaQDR0gQIPc&[FD=^-GRC#Z68]eAbYW,:3<#;H@RN\(_
U/K43X(B&4DZI2[RYA8X>K&[EN6T)F2(U>\H3dH;MW<<bX.3PGE(Y7,C1.-L=#Z.
bA8/AS_B&LfA@/:bOG?->bFAPG=&5^IP0IaJ6WWCd43UH(D7cOe5LZZ55?=X8W<^
FF-F<\eHeAFebW<8^Ad.UZ@b=FY3WTgcHG.a]2M3-TP3^4HSY<-MU\WeL8=E@MP2
3eWK<&C2+YL-U;-c&R7beX#>],S^S@D.]?eGb<-92d556ZP/1Ne.<@O>f30?<1S2
@bF;gNK]0H\aVA79>H\U&8e[CT;:f1K5\D>_1]TDdV)-8;b,NA8OJC0=1;FLS3RC
/Q44)0??fbR)#c]IQ[E:B]aTHK1);]ZgRGPc]).-10VRM#>4cd.E3)>R&OEW#F@:
^0XLR\6D27]36K:8#3+eNPFTY4;46NgLL;TN[W+RX<WU<FJ1CB.78\(^1:eHBY4>
(RPg3,DM=F)VLX@C;]28d,X/;H=2-2S@5_23X:DaQe;-(:1d##^PH,;ON+3dLVFg
eS?:P6[U6]DK9C,EFC8],830Y1N9,.@7@E:cGL?ZSVeJ>?AX[?-dENFVCL#2/KS1
O4:XQZWd4UH#W6f\YE(]:KJ.H?C3RQ9]U;QJ<F]U1<UAG/=YE5<MbXH\Z,P/-D(9
-d443UGUegPGURXRXQ.)BS95+8Q_F\PI(4@)KO=N/CFGTc#f#LJ3OHeeNO?EG_,O
+,2B=4=^N,<5MDgCcAUM/c=,ceb;.b0cIGQ67LdP)B/)cNOT/.X/<P+-XbF)JE/N
dP1.504X\KB@Eg\3;I\^Y6S3]JC9J<N?dWE>Xe7/O^eOOL)?A3MU6)XNG5H0Ke[:
gX&dE&0/aGE&g_,&72US^;._E\7>0f;CM/K+b9SKZ8^//,2ASUBE#K<DI&/<.ggX
JEH?1McFRaQ>.C>K;R8,[HPRA,.e.dL)bNe\(=7Bg(=3N6(_X-M(_PQe-c&F&&]G
,7J5,3ZY9@g(dD>R=/e\UEV(WF@N)-24TIeXVIFN@a6bV=;L^PK-<(RW1AEAXL_>
/0:a@W5b\c51;>.?#C.LIJR?)R_ZP,0]BE\+?GgG><^PYG6=MS;4@FU#WSVYF^DQ
Q3Md_d\,WH9/X0/F<UXEf<ZKUUCD/&F=IWCZSS3f4KU#^IeB.W[g?F.b2Ic),916
fAZ0)IY3J]f4+Y0E<#^UT[PMNW/:41-72H84OB)FgCaXJ<#Sg2B.(D5ULOR356>g
0V3>8R1;4B6Sa6Q+WZab-/B+\g-3HaC&1M6UZWVBA&\50G<<eG9/38_Fd_S,4X<W
.bZQfA\/C4J;E;6G8AbN.N?Ref[cLSM4,Af@7ZOH[<?dd&>>R2@SO1HK[HdCa723
dbKWE#M#U9&2XW>@>25bX(dU/8QaMQb=AEMEJMG,[_[56:;@/M&YUWX_\6B779]]
QH]D?:,2BeKXELfW@R++H4Z&,6DLO8@dg6QXb;\9KIY\._&J+_)67+E.HLAC.<Oa
7DdNRbO)OHfC3V&JB26E<[a^ZYf2g#DCd:9EL0;+9]9d#.3[&..UI[25=IaXN>R)
7<gE;)fBZTN#G;^U(QC58[XKF2KIgGAK\,A#<([SaB;^\fSIT+I(T8a)6_&Q:R>(
\P2TD<>eDV@K5R8M>C;3,2M)JYg@]e-Z12bJcZXfM>QW@RD)?SUR(-6#5fEK0.NN
gW]O6PfU:?+,L.Ud4<Jg1;655;YZI9[.HN@AZH[=d</GbM>KA/S8ONNQ-Y5ZaXVP
9+N9,T9.2&6G<#VU#VKeLYY7gY=5b&Y4D<6+Rb9c1?N19VcX\gYaX0;5EKRBfAdQ
@F-IS1;A[,1XRC?.NEO8[Ee:A.W=XN\WZHQ3:T3TZ1@d&.]V8:YH>Td#4#9A&5]C
SRI5KC?Q_YY8DL/TaP/3Z07_M&JY07=2Xe7FK@(cB0A.(YVda,L>A_GA<K\>Wg9=
Ce&(JPB5UOQ@X+=+39WKAZ8=DF_3FKF6eH2U)H-T;]DD;ZY=@+L<XKX5HKXMHBK^
J9WVX=CB401\Y)NB2L6:)I]G<NQgBWZT]/RW&Oc_ggDRP\XT,&a^d2IAAGB?gF+Z
KIM#B6O#>2g_DME)2Pc[^KDT&UgVHNe.LaQF+4V-Qg5@;+^c0+>CbgS8L67:A//_
D5U188\WS1Vfc8>&L>]f\H]dYQ776@0&2,7eCb;=#5Y3YFN_P+MJ^(TPI)A4cOgS
+O0_:FR3\_26LT=aL(PU3T-P?R24]dN>EUAY0/Sa__gJc53--ZKcgL1d.,>FN:#(
5gVY.@R2+f72JS<2\32e<EL4<&9A?_7O1A#IKJ&/:]aY7Dg8gT]KfbA34RJ,U=04
W_(GEP_4b#\#)MCRM@&PWZ03\1S6F]2-@^b;W3OOM@;DO?1-B,(g]TGELL.-+VS[
&,-8#]bPTD^@d(J)5?;@Rde6^43_(^d_Q[VYaFT4a30.[L[UB;a>XP=0L^2M#-H(
#]R]gOZQ1\ID\_-gc,H_=RU(??_3be_]fVaeFI#bVT#UUg<9U9a4PZLf+Qd[0RVV
<M6bJ>@d;J#1B#2SURP(bc3ceP55f^0Pg??41E@Y12N2SfJL\^d29<OVIF&IGX<T
T1K?.HD9d=()<HGD@7^Q-<dQ,bf(@1U)QYP:\.,CUEZ+6V39c,CZDX._S=f&E5I_
^W1LCZ([9V?8)72Z0QbT_QOVUMfb_N7UO,=#3H]a?DN^43(OOK^E)a\V;Wdbe,Q\
@_5P^g0VN\3U65d4HZg7.EW6B>/ZH>6^)++,N6(VUc+HSH&B\7>W3P/&d>]<;gZB
9G.8bJUG@XACHa9TPF4VGaVf:#Wf8Pc1O]UJ]^1W^Hf893#E#&9X>]E]L)1)PSS;
C5W6?@Def/@@,G>0AZ<H>Z2<-\f2DJHXDbM-&7BY.DdF/?OBP84D(5,gUL[TKZ41
##Y>D;:?J1SdSLCC,,]S?\N)<VH\NM[/d-C\9;80GNS.->9AM7T,8TS.d,c/=/J4
\gf&?-gbQ\N)\.Ce]c[JKcOO==0^gd@RKa]4:1Z_0KGQF,03f>Z-;=SNH;P@X:Y8
KQAZF4EU4DAC-#dSN)ZC;J.TNV7b_AGY+eUWD,V_-bE=a/1^:?6GM<aR+),#OCS^
1aK-?DO:=>.#W0KcPMOD1=X5_@_D/:;9>FU9\b>PF.B#Q36)C:\?(dP>W?Gc2-:3
0?7ADLM@>^T6@O16XRNaH_Q8B?E(?Zd0GbScM(A8L1UXeK+6d-0]f4=?;VaG)6.E
+YWVMOG=FCK7N(RMC:(YZSWa#fT_bW=_b;886;]LX-(HR;cUNd+Q?Q4JH?#gaI=S
0[B9-0&,4UdfP0EBE0bUO9]@UTgHZ[]L([6A=aDAJL@gQ;):C;K/H\;5<I8\2T@8
DUH)BG472ECgEaAbe:FM5A6UHQ3V.d?@70:@,c+SH[aXgb_VFC#:+#C5D0,G[\V\
&VE+4X.6gED=WRdc)S9B-;E;FSXF&6M/e#F?-RW8d-D1U3B(.+KHG&Pd^/Y.T<DN
5@.<;W0,[1Vg1.OcaHBf(7:Z2&PV0fOL_F.=dXO6Tf6RBD&ERg#7R,T3A1K8Q]GI
FDW(#N^]N/c@T7=+FO2K<<<URLdVX<.gKKgC,(F5:+C@44[KL=^G^#7OB)g1_>O[
a;/C90TI4g77SA2MgfgN+C4[DWVNVP;/P79<d>b[XF5BCDE=cc(1Q.VKBQM<?&L^
gd0+0:@/OW/TLbf)B6TF4;-XW(5?7>AYaJJW)/cO7Ce>6[T8QQ\fPbT\;.e0-FW6
Xa8J.VRD9[7D]:df&^L\D2VRc1SHe>0cEMGT>:NK#,&cG&\NTIRAD=g>#-f]RI\?
N2^^_Za#+_?Q]JfB7<RDB,<_GfRN^@H9]5EL.6&WO?<I5feC(\X&>D@C14IN^Ce>
E.RCL_R)BffWDg(NS5N^^PbJe,MWJ39BXNE2\8XAL^RZ#C#;6L1-IX^JQ0TMTCYM
@Wb&(L#&MW6WKG,#]dTR9,+TPNNYC:_d-^_5/#>:+WW2P/4IONH?EbD)fB,630K.
UET1\[@eWaVU#<Qg2bS#/ZE3^Z:Na,\BV1U;[DXJ+MIBf_+W+G-2@C&((P2Ha,8N
47AZaKV)5b9)2?aY_cI3f-C-,L,WZ/N_MOb(7HJ,S1O>e</2V[1QAL.)6b&eLFK]
U?;8Ma0(LE.\ebW^+8V:7JFCQUI0\+,LO3a#b+eMN7Jc^T,9Jb:.3;N4X(?@(:G<
Og]7?SKXOS&31#KY\:XG&Td(WBHA>bb1>01<RAD(D4d&/A=V3>Kg1gQEY?&+@d&F
^4>=1JZ-B[R@5SJB,)dJ.&[Y;^#TV5-We/Wf88aQPEKWC(IGU)EFBBFE\C&>]b53
M_g=&IX][#Gg@G2J6fEGI6A5fU7AQUgXUNF@BO&ML&N5(UI?V<T)GRY]Z\;KE-#G
;^CTKD5E\LVQ0IC.d&QO:=J#U9JA__;7K2fD,e_UU]/\>c05,2)/<fE-\,7@B?JB
0:U+(^SI\g_ce<_Tf-J=@Xc?(aM2)Qg;cTA<;P59R1.,.gD)0=89)F\G,g,B1L#e
bdHAb4,?DTbF&bWFM9d8aTI@G#A.LDG>&Z3&:+>>:7U5N<>&63bTXGKBHfMfY\?Y
0_-R)-Cc98M0RQ.IG4(E8=.:URJ9LQ_)+)^7O6=32/+6G-F:8NFM<=I;,R9EWI5@
bbA4N@eQBIX:;X(HgOb##VRa_J)ISIO)N]XB8:c^;TU_NUO7T(VGEB>)[Q_FNG4V
RVX&@B^T0.2SSDf>Z52KZ4TC<fIW1.d9.f?dG0TOQ@abM]-&S9_6X0b@g_4B[DX/
TUQ[.b3]R+@V?X[S[A2>:W=;=0EW,Z)+]XR)cV&VEeWJHR)\H0b-1SHAEX?<X\LT
W^CU[LT_M5VXU2902gAS?bGT/d-ePJKWO(HK>+afc8ab=7A-PS8#>F=5U<3[RS2Y
G@;,_OO-NR\XX/ZJSNJ4@^\4Z)=;=(C?Za)255&Q,;cLS/WR5+f1.d##E&EO^,K4
\aP<(4R2ZQFSJI<U(RD5b59UGSCA\=U,4.U@0DaDE45;cTL.Z4_CY?Q)^b)G/:AT
TE]ZNTa<bR3ND-;HD^(A:LE&M?UCM:g//0#@K-:H)bDG,-&\TLH\\FDQT52f7R7)
@S>:eF2\)0g4YT4,WbRUdQ-:=T,+K67_eE_fM_0U>DQEY9cf7>UTD<3_=[;7CCY<
GdFg5_I@F2,7a,3(a#Gf,Y+aU6M=^S-a6Z:>ER=95M=/8F(OB3]&_c?O5]_IA^de
)Kb4V)cL4I=X1VCAGQ4Mf3?Y?@1:b2c8Z/cb@B)VANI&)W9/..0TVVgDIK+EHbVN
BZX7#f9;>bPR;>K7/)Tg+6#0L;X)EZ+;18RX><H\e5G>/AEP7P6,GG;?5^VX_D?V
F>T7R@3\A76]Bb?A8#_f19EM.;C9(;IB8^UKb@BY7[?AX))L#Hb<([/U#DgUL(;?
Ud>VDA-^c16ZeSC.cLOGAX_-B#M^>0T-X0d#>(X(fd&f#/3V.=87^=TWFa#BU1?.
>5H-<H?6@Qc9@^#S@HJ,YK&f_Ce<Q:L05:.SYH?\e]_TbbP,.g#@@[/WPO@7=V;]
(aXf<KdG-_NdVTaZ.(FZQ4T#bWQZ-CYZ:\6X@,-TXQ0,Zg.1P)Q86/>439I[e_?U
-XEUX]KS4V:,_A=-44[UF.c54dF(&UN<E\H&_B@WWOf(Pe>>M_VTSSJ9RL3+;^cQ
&e1L>0=9?G=PZRUW3d9f)QD;,]ZRSGL?QW0O&Me3<DC;UT_(\2>J12C7QON&V(#U
f)#U#/Q1H96g5T2-41E2=R13eI>M&?95#H^/N<,E>\ZGWg3&TG#Z^a>#aAAZ?&,F
^<(WI]a/B[E\1?8IGSK70gX,+5=8UEeO^V_;K[/7>#7dgM(ZL;f&4)A#TO2Q31Q.
Pg?c?0g=<-3Z1BJWEgGWAd^H49Cf8D[9Pe#U&cX,\ME^AU5dZ._>?FMbBAH3c)]d
f[=)b>7UM[d6C;dY13UP:#L(3A^6)0f-4J4YOCE:U@?4^N#g,_^].8IfZ8F\R,=a
3dB=T8I.c5&N-64F\FG1J=@P:H@Gg7-4-:QPLBQ6^=_5Z;&I5=R&?3(PV,M??^S8
KJR@aQQZX^QcLGDTT@/=N,3L?\BMVL11g,.G6dgAM)c;6g?aRFNAGF614R<\9WQ5
MgS><:TIVE-UeRT>HG5O&+J6)U3UQB2=1@8MXHdcP8dF?SK0a(<UKTHfe:J2#E)T
Wa8J-NWaB0O?\&[ZAE37S/g.>3@C;[QKKbW=>b]1DA_DAVfGBf_;H\XdYD8-35g^
B&3OKR9=8V&ZcfVc=dFQ(NReN4O,,:U/9,KG#,a8[AS+(Q@bFa2MWVLOZZc92HVT
S1/MTeDCbe=177)F46M>\S^HLT@=L](YC]S#=B:bdMSe61;C7V[2,??<4HK/W?[-
>_T)d)bVbD76_MV7V,IPbP:cAeb^/KI[@HNeSUb)PC\^9GA_4S\4([.89-F46B7/
XS@D\4^<<FZS7\\\5Y?A2M)B81HR=L#<f\eKfWf\&fWUcXQgN6TVT2F9=_f[XXT<
T:0<0/+QL.RS1]S#YSPb^UYY@4L67IdWFM^T\T1ZJ<A>,R4bA/E=EBSPdN1>b/5O
6=:CJ[>HCBM.2HJOXaPD2MYdQ56;])@USMeS?<Z,DaaZ,3aVF)=O+Cd[(NA3Vd#d
&AT-?3HDId\E<1]CG8/(^2gB8CSE(>^Ie?.B69SGZ:P7.LW:VU^e#(EANE;C:@bL
49f)eH+3==_/-a9>X^>VAD3]V/eJf>>,VZ+IJ\ZNb1:d_1?D/DPOF\C89dREC;ZD
EX+Q^AgOUc<:5A-2W#a7;=,OY[bX/Jg@H&\Ne>G#L3>35=](L.RX9&dJ@@_FbZ>E
@]H.HY7H;5Rc\>W&+<P^gaBTT5-[<S2RV=)_E\Z>J>9_DW^5^[eVCabNGG(SJ]2Y
VO[M,+a(3L?5U\?F[LS[EZZ;_72,G6Z,C@Y0\=F(YHIT.>U2_2,=Z79,?-M2=:XJ
JXIeX(FW&2B_0+:SU.Ye??Eg.&bS(9#816_#81?/aF2?#3\=#c=@78?c6+C\6B;_
#K=GS,3?e#W,?<VVCb&_(1[cV0)G=#N2+Bc]L;RD3N.IO/f,0,5XSP_eZS@MGIMX
61XEgKO?R]N.][M6WOKH_P;LD]5G^8<aQ9KccD_59CG5/c?fQ[TAN86>)DXd8JXc
HGOL+^ZGVaY9]Yc1B4@GaZA3=[GQ_>F;cQ5=LdHUXfRb1DDJ)d;#ULM.^I<#VJcJ
J9,&UV=N-4BJ0+M,X?=UG.EQ#Pfe[#0?W2bXFX#XY-JcP(FJKOc>:@2Sg(#g4J8V
?g9HVEI,U:Y-f1BB2cX#/VTf/Y\@_53=9aQY>5.S]2eZVBL]4-9RXTIW?WLP7d,3
7L#R,-F-g>KDQ,CRU6FO5P[;Q8PcV\Gd6I1L&9)f>B@+B0<cOG\_#gJ+#JXgEWfR
+T7?O-;U6,3)aM]Z_eE@(8eDI(543+IW]CfKba1?-OHW0eA&QEf#B?&]+^Uf4/&K
:0ZcTa<[=:DSR(Q0H-CDE.F^>g]SU>bT?,])/[B@A<3BD3[La\ED=c,2=-1>EN8_
C0X<+)>ABeUB23<2b5,cZMZ=;g(3:C&:5Y4XI[CL),-g_]/_Kb@Q\<7dW,d9]3:3
B0B#CRQRYP==a7?^MGW24WHU8aGGUNL&bfYbH\PedV[S-;??\G#O0[DgXW1I?W20
^TB#9BG?>[+cP-)YEcUFZA<YHNMU4f?@4:GZ<AW6S8:E4H_/P@49U<G]X)X1Q&=,
KD\=[^_V,eCLDCDQ:6[O#QUIV;Je^dU94J:Z8g6;#a,G=>DAIC5E;GRY5[OW\C7B
#Y.fSM2BecY0D_CK=;8RZ)]60eAL3PN^V^9.fYGHK6NZ[E@RN7_(0EM)@d6F)cbI
AJ\I2CF@F:T^D(4^a<gegEB:>S7<^d_b24IF24P]QZ+gV55,f30/g?AJc692_^I.
)I8N96DX-JZJ:K+AcE#)C4K<5=QMe.TPG@S&[XCdZXPdb<8/2G7BL)H-?.g4/ILN
)I3O([[g^ZQ_2\.WV5>OL1C=cRFg8EH_:Je^EM(SFYa=XFbAG30XA5Ue+NCJJM,?
-DRI+RdOWMG)<baP+JA3Rg+<If-f4#<?3d&&+b/[@V_#VQX7g@4ZQ/34K9M0IGK@
\LSX@d#)/VUZ1c;;GTW1SXSZ6Z[I&DXYQ<T[6T)0P6]E?Y?_A\O/]>UPaeHeP)VV
HW]I<F90;7M=NI#<<H99cS5HBCBdf7aT-Z^=AKWe?CC8e=IbbSaS9FD\I?F^<J)W
]aX>SUWIYWV?PbGT@;c]@BH#YRITS4JT7.1e9Jg@W9+Y\3^^dE2;U1/XeQ]JDAg2
EJW>DSK,PKF6#&18POcJ0/2W\+M5P#1;;L_(9IBK8E1C#9BNM[G?\?@ZGOMecO[D
VI094B?;EM0:LMKYU[BHJ07-f8A25:RRQTaXb<52;Q=b3)e.;XS@A+Nd@bd(fI\X
:Uef.=M^U@76A.1F:J[F-A#/K;2NL21UVVEQ-eAfAT,@G;U(Z17B(X^3d/EW.^La
F=+ZBQ^K#Xga>f@V=CB9_?)<,(HX@=Wc/]93b5U3S8&I2>KX,-b\.3NA1XD;ZObR
4JQKT+&LKLFDaP1+7]>Y69O7HR(T>e/EA#68LaI6X6-J5Q0K+[P)P7VW643ccU3?
SSXD=;Q<HG=(.MTUMWT=:TJTc_N5#089]5b58TO>6NZd1X=<<I;3LQd)e,KF4WAL
3ZX5V2\W<fX+c@\UJ#;[QBO&S7FCG>>CNV/(5J)E&S3J7)1aCY)cJWFKEgS<dT2Z
]@aDUXA^L>S]Mcf+P&>9_F1(94R\9:IZUE&3\\=_agE_P5]RK)[Kgf<5GQ31X1g=
QeWPA:R,+JIV]GF\QH<-\ABRPTf0&9MNEaadd0/NAKXP#AIe#_M@IM;(H>?8RL<&
I]S3T^P#D9gTeAf=Q^M6R#LEX0<04Y0eUZF;4ML7ZC^W@L@3>?B4)fWOTcH/4DcR
e5]FM)4)T2=#d(FCaER7L65+>-,X#>4HN(E1b,<(02DY]4FbXI.DK>E9CUIA0<@f
NEU>K]+:P:D]#P<YUOZPN:gMXcL.++SS/-Qd@)f8]/H[,&J7bJf#8;;C0>9;?2YO
Z5^FJT0J2J28P\OOcL.g2?K=LCP)8gNPeDf2(^NA13T20f8XES0:4a2,,H,3?T+Y
J@A(9F:_c7M,5fIgRQ?NQT3>6HTJO4g#J2F#DNHb;I6YTC(,d6XH(L9@a1MaWZeH
7A>I[JKEEJRA/fgbY;.,62ZH<>e_H:&)X)UVOda-gP31X5_-DH#+R&3@E+F75_KY
]AIV_P,[LH(.ZU=.S#6W?>?TBE3cdS(6,T:2X\Q-UAHUWQ5[QbY\3)f_dW>S/B]C
ecK2R.2Pa,X+8]CM3Ud+M4WVYLI.T3Q((&,:VGF__V-D+SRVWJ\4)535PfKb)&]g
?G>P)GCH85,VY07LH;B[P0&ARPB&b<5-RU(_c#1<&a@1IWSb9K-8Q,5c^^fI-ZY]
7b^2HR-4R>,-:Me7TMV;eV4?#2d9cLZZBPOIQ8O?CZ6PM/)31QK<AG/8YBSKS<FW
ZC@C?9.4VYWZIL@;g:#7dHGg;fTL?V>H;9;^C2FO2IQ40[P./S>(d0eL^FBE^;D5
VT]E@9<W&(3U&&A98U_K>T1OVdBbIdc1^-/T/7;deN3DV?+4,^.GfPDH?M#OKH#g
W#d4+L7N=ed0]U9c6H@g]MW<DRBH=,S[?_8BcJ3Q=@(@g;;@T85dG77c0f3FOIY\
6Q,3eTR5PO-UY3]#FeV72bMFAOAOE_QJQQE@A:NTY]W.7Z:F+J,[N/]S=8XgOK<Q
#]24H4)M#g+7Y+#M>cK+XI]P,ffeJ^:I4+bNE47.+M))SUXJebP2+G/ObHbBgZd@
9g)FeOB5KL7=b?ce-PENYF>.IfT5#R4f[=3V1DLgXdIT)0>da&;-H.K&3aDbQ>JT
dKb38RSV=)4T.DC)g/Ia^;=S-N+Y[E/9/54:@;1YWd^T1V<A/^&8<ebS\),M^RS4
Z2/@a;2[.6806df(RK/HP1/N40P6g&F+Ee.LO^<#>Q3_W8&:FG_6;B@MWc\c[3[O
3PG/]A76c]#>X&Z@#-]85G2R3]M96:4U4cf_>4;N<U;^_Sg2(&,.D_)19=V?#AES
_64\Dg8PKLUd4:a.;/H#.+&CMFgEF#TNG@LAcVF?RM>?I]RH+J44L[.8TK)?L>DM
,#PdBfbB>F^fGJ?(/ML0T[ABc+_Y5\/Y_BQ)=D63YW.d.LK@;4\-U;O)g;X9.JAN
DCUT:=J5-.B,<CTb9,#?_5&@/fW#e;O,dZXW(C?_9+S;RX_A>LB>./@KJAC4)gf_
b>RWN/7;OH,EPD#dOMgRII6FPFFU_O6DT\E?V&;W5(\,35REBM,g<a>J>b.E+YQZ
391\#4#E^BR6U?96=,O,UJ>@SfcV)N1>>$
`endprotected

endclass

`protected
NW@@Sf/eaJG4ZK/I_;7c8X.OV@c\YFb15SR,/)Z;Y0a@;I=H#g6W2))[.:<&N5,0
O7#SLQV2\ZdCD810\(MWV&+_ZZLVgL#UDY^XB1@YH3d<K)M/2g75;5/+5J).2dHe
4fHJZ>]X0Jd,E_+,HLSIFgBOTcR[EP-JeXL[bQE&Ga7b7Yc2IfJ<LRJF2XS:g=NX
P^?U=?TNbILJ3aV^g2<ZS#Y4e,?[(KF@S97,6WHZT&NC71_VO@F)0:VQQ(=[P25g
/R<L0QV<DfV)JP2R+fY,<c\=7>+#Q1K/K-D3(:OQE@_a0KJQY?7D),GP63<XXU?W
a9eZK;-24YMF&O69KXKSG;g.1[=#B+QV?$
`endprotected


`ifndef SVT_AXI_MULTI_SIM_OVERLAP_ADDR_ISSUE
/**
  *  Master callback class contains the callback methods called by the master component.
  */
class svt_axi_master_overlapping_addr_check_callback extends svt_axi_master_callback;

  /** Port configuration of this port */
  svt_axi_port_configuration cfg;

`ifdef SVT_UVM_TECHNOLOGY
  uvm_tlm_fifo#(`SVT_AXI_MASTER_TRANSACTION_TYPE)  axi_overlap_addr_access_control_fifo;
`elsif SVT_OVM_TECHNOLOGY
  tlm_fifo#(`SVT_AXI_MASTER_TRANSACTION_TYPE)  axi_overlap_addr_access_control_fifo;
`else
  vmm_log log;
`ifdef SVT_AXI_SVC_USE_MODEL
  svt_axi_transaction_channel     axi_overlap_addr_access_control_fifo;
`else
  svt_axi_master_transaction_channel     axi_overlap_addr_access_control_fifo;
`endif
`endif

`protected
V27ZN3/>6/)NF\L@[/T.0/ec-7J@-d;A^WLUGYYXE#I/6WaS(TC>1)W5=]_aTbd_
IV-9dR2Y.0)S+Qe?)fb]-0KQ<.;03aT<[W=/CFbKC0KY]9/FD<BMENV9VZ&c1R7g
Pg:.C@T1S4(2#=<FFL3.1^[fC4\,H]7])3H>ee]D.I<.fbXF0Q?Qga&P376@(#\8
.]VMBEc#+Q)WKP>:dIFKEVF(9H(-MLD?46V=S75]Q2SgZ5XDMWa@>d@.]^K7,ORf
TRU=gA@HQ8-<O2FT]6Z0^.Sg,M[=a8^C\;5;:57TD&Z:PaIPD&/:;f6HNC8DVdU8
1Z8/e6[DI23^3RX_HP[X)6MHALBb&]]JIQPK+@c)465?c2BJ8EOH80[_J)=K;3Wb
CdX1dR83S<>BZPG2OgM=66J&X).K^WE&cRL9BT/D_gc0TfM#c]S)eFP=[(I/ITB3
\f]R)]Xg>)E&/HL/b8PZT]:>IXU-]aF:E)3Q(5#IS#52)c@Jd^-6I:6HC2e@9I,N
@(bZ=ZgBc>)&MFD/3:aaF-[[JA4/YLAc,c_K72f\,::/QcPFCE@KF<93_+52OV-9
3KER>)4(,4TgVIb>e,T72Z(fI?eR(,cd,X&W/@[gCSLP[00/,5e7?PV<4XGE-ACP
7eNEJCIESP4F1Sa32B^O([/&5Z5^4@/;>$
`endprotected


//vcs_vip_protect
`protected
VO),E@K1I6.7::OgY)FK+6AUL;7Q9dT@[1H6E&B3c#TW#^4Q<(1#1(:_N0<=DRIU
@=AS5?R<_K.1<\fYPV(:dNC>GX/gG?=R@L5c-VV)&DY;]b._F=(<KQ[AIE=Zd]e>
GI42)de0@=fXSEF^C,4A<(H_VV4RWJIVNW0RZ_IAN(0?Ud;]3=D3YEff&BdZ.S+2
,S1aX+UP]MK]]aA<BTI]92c<T+KA<L@ZBX0\&,0GcN_F)/UDMH3XY0V9-)0.PPfb
Y-<T7-/aDQ3L0g_[:7V)^;W^3M&&T5dQfBM+ZeJaNKDQ54PEBUSZM^<#M\UJ(-I6
587<FO5Q(1&[FT=WUKE+aJB.+H(:F#>WJV>R/-Rf3I;BTbI:KeQX;G/1@;>:_@6,
S.FB68H1K52Q])H_)\&W/PA5E(f==[accL;WX6U85&U)M5e0;G[QS/0\6a2M27Ua
[f],BHb,X)]U^B@g8&F1\?cSd\1UCP/JO?Cc&_1TecYD]>LGTHEO4/XG-#T)-\9S
VP.PFg7:IHbfVW+U3-&7\L.YE+=3FT)YW3R/WGX=-F[,7cI)].Te;8AMEYAU&)D&
[bPL]2dBTf9IaJc[Dca/M(/PH=F_=GD4TB][Z4d[GA??);6I[.\:BZ]8#11?PM8J
A(-=aQLLfYeS0ea@Q,S=J&5H;7CdaTLOR^)+9N1?W(SPeI?Mee>O@acJC[Y,RbI[
6X3230X:H\8#f-EbG[[fCde,VCKG]0f##@e@g(aZ-eJgCVD#D9JP/0W+)VBWMG(C
V]c?)1d.Xa_M^+S,ZL;KR/g=7(46,8+)-eX>2Xb(#L;Q>+;Ed?T(ACDHPPUVGI1f
=4W#,8PA4?6<PWK4VKEV76UaD7X5V>&e\>YR#^#HSUYdB&MV2(gbVS)UG65a8)\J
M>U(R/^U+L\B4g66VQ2<0Uf,D^TNG:7@3]e^Y8#ca=8RRK1bF-Z8BKIIF6SWCY;B
:UN7?=(6_f#_?WfY]M<68S^PUC9BM=;eg&WMPcDL,M+KZ3<\]C>dJ+0J]4?-@NL@
B,GN,QW0?=H#O_/3R:Y1_?XR58I>)CBXK6)ac3#b?1&;02Pc5D:\Of<.&]UFbZB_
^g/G;0bJC+260C>\;Ha,8-3M413.<WMe8INcZbe(RXYYP+1:;eQ)#U?dP=]dEN3-
&=0MUd>>:F\,.I.Bg^R:<Xe>L#ZQ]gPBPH#TFS4W37a4(,dQ[3V.EVR@V?_&_+U+
GFMKK-:3U3R,D>4?4BN;U1(g/.TOKEK@AE0Fg>Q?WMc/EA88:J?aR&9>:H[?R:CX
OC3SOg&NWM0G,Q^b)?@[G3edL43J1?/QN126PBG\d2VHMA^AWO@<?3CQg=/SRV;<
ZJg9X]9-_,F=6)ZX51O),HJ.eLE[c:U6BdVE-TN#FEK?J@<8O:SB.dJTWG,0CP6?
cO:>Z\TH+36BD=-^L]JA9:0Rg]AL_30[:\TKab,&&7OL#[<5+RMb?XgSM^8a/Y5H
R@E;+2LSAg,2?+UG0-FME4<D7gL=C@8]D2H1QV.T3FfCVI9<2\Zg_]O17&([[?.N
Ye_ZgLfP&^DP321LLW3GV8B:&_QKP@N9MGIa+T@<9/SKB47#Heg3BGa\MA>7DLAI
F/d?_.9^TbBf:d\-eb6:A;)A<-V]:4DH\dLR790^&BR1KRJ@\93d9^QR4J))ZXd9
T6W4dgK1TRHfKT1a7#>1Z98+Z(,c.L8&X>6CPJQ8TPIH#0XOCOWBa@W9XT/3eP_1
-;X1;THXWVfUJ/X5THS_(Y+(F7<7+4&RO1HB1GDEJXfdFD@YJ=E(18_D\e/dXPZ1
;e>8[Q6Q2:#FFV/U\NITK^6GPY.E+/_]a8ZJ5WMBX]+NJfC4;X7+0,eH_..3?Z-_
+V?EP+)[/K.,7;VR5eEJ>7N3)7)HAKYF1XEW1BI/<EQ9OE+>IXZ3&?33T#abXe;g
I4efW3T&BYeE>U=K@KTA)12VL4E<;/L)[M8/g&54KcBWL>-aXI4TASI5.a0VG+ge
F\cU:\?_[Y@DT1f#?@QZ/\2.[)MZ([V0[J9,=CC&YPDY5d@_b_RBT\AWRa+@B+AA
c_\Z1_2L_<LgQ_(IWKg-<fBeeO;:<+cA3()3XVYF7\Fd04&0L@\MZbD9d8,=5Ed0
^CXZ,1_eVCI;AM4DY^<_bIMKgIQSb]f24C104C-,/=>E4=KC8L4T@=BC9^W1VDf9
c-ZcdJ^c#5b8dT@NeK>aS^M2UcT_^Y8&4+_=9:c;:-OFf8Yac)TI0KZIDOIZ9N/U
E0=[Y5W73PP;]T_SO:&064UQ.LR2KML=I2>3-Z2JY8-N=I/1NKGS]TJ3XA(PcddH
EXKI,7bVOV:P?^edDD3OD\DQ(E4TZ;f&7SdP.cd+-YLI31c0@YQc];@@D;d)gNMP
1#=-a?b+CW[XS@CL.F,2g&,3KS4C73QM=g-9)[J])Y0V(0<9.dCaZ;F<KW6Sd8[\
>+57;V#^cL];OMB(X3cAID657(H;gg;b3d/KBH5V_ZL=e8QcZB=#@I5WK54SZKe2
J:J;LdMT[)0;VZJ8ASOWD,f\IBF#c7H@05,V?&YIX8U;-J=-X;<^Zb<0_Y+EZM,3
D@NIPD?-F8[0a3^.G1QS=_<fb1K(40c,cR)_,d7,EGHI5R7^Sde8ZcQWHHXL/;N>
e1A<9T.J#5CLZ)GRM]<78/FGSZDZ:eFA2DKeU)U3g&1de.dFRc)Y\?E(UZ@320IS
P;A^8T>8X0B8@I.XeD<MGN1M^[L&LKO_+@,.MUGeM5bR66fK(+-2bV.QA<&Q]F#b
5fBJZKXVga?0)V#a<S@Z8c2ASR=T7TfC0D?B6b6X8,b[6B6+U6@Fbg72c+[c2dZN
0]:ed6DX=:f3g5M+EWPM]D6[(H<PRHPXRc\.A6))#FRN97.?K24V890EB>g;)I67
dIHXB5fSE34bdAeHd621(S&_@(2DAbP5>#2].+5Sfb38.aP)FIQN-SG<ZR=bFEB>
0O8H/B=]:-H#c(ALd4:J1URC1V;/ND6]O9^\D]\8CP=a,adc?adLWV8@]2e/ZRY3
L(NCF=;6,OSU3DKcIL6P5PcL33BSGZGH.7,M#)5GQG@@5RMbSc5M7<fOAFS9N&SB
<P;8.d#TeTa8LCg.U]97RSK8?<@,dPa4LIgQ3J7]L7XG/+,#NBT<OJ<;ZC:F^Da3
>JWFP(F#K/R7=_.MO]d:=?WJO(:ISW[T/@/NVCZHVfWRdLK5)L61ZAR+.1IWWTgE
:)Mc2P-0[D;C6c9IU<-3cSVQ<GOIbGLBfDUO/.Xe<,V+?gWV//U#7ZdY]NdTZ<bD
(PGg5b2NZXCdFM+c8PM[LBG17M2<E[J;gN4#V]b&\e?eL26TA3<bP7XdE,)Vg^Z,
FTZV8K9A^eU7Qd243T#=Z#?e-Y^[^J3a:F5feBESIIS.6LY2J,W,2QYg2M9I<__5
8,d&/f4#LEM7-c]H&2J:7)NMRC09+?G9)A5VT);5H(cW9gLQg)XB9fJ;95?=MVHTS$
`endprotected

endclass
`endif // SVT_AXI_MULTI_SIM_OVERLAP_ADDR_ISSUE

`endif // GUARD_SVT_AXI_MASTER_CALLBACK_UVM_SV
