
`ifndef GUARD_SVT_AXI_SLAVE_CONFIGURATION_SV
`define GUARD_SVT_AXI_SLAVE_CONFIGURATION_SV

/**
  * This class contains configuration details for the slave.
  */
class svt_axi_slave_configuration extends svt_axi_port_configuration;

  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------
  /** 
    * Default value of AWREADY signal. 
    * <b>type:</b> Dynamic
    */
  rand bit default_awready = 1;

  /** 
    * Default value of WREADY signal. 
    * <b>type:</b> Dynamic
    */
  rand bit default_wready = 1; 

  /** 
    * Default value of ARREADY signal. 
    * <b>type:</b> Dynamic
    */
  rand bit default_arready = 1;

  /** When the VALID signal of the write response channel is low, all other 
    *signals (except the READY signal) in that channel will take this value. 
    * <b>type:</b> Dynamic
   */
  rand idle_val_enum write_resp_chan_idle_val = INACTIVE_CHAN_LOW_VAL;

  /** When the VALID signal of the read data channel is low, all other signals 
    * (except the READY signal) in that channel will take this value. 
    * <b>type:</b> Dynamic
    */
  rand idle_val_enum read_data_chan_idle_val = INACTIVE_CHAN_LOW_VAL;

  /** 
    * The number of addresses pending in the slave that can be 
    * reordered. A slave that processes all transactions in  
    * order has a read ordering depth of one.
    * <b>min val:</b> 1
    * <b>max val:</b> \`SVT_AXI_MAX_READ_DATA_REORDERING_DEPTH
    * <b>type:</b> Static 
    */
  rand int read_data_reordering_depth = 1;

  /**
    * Specifies the number of beats of read data that must stay 
    * together before it can be interleaved with read data from a
    * different transaction.
    * When set to 0, interleaving is not allowed.
    * When set to 1, there is no restriction on interleaving.
    * <b>min val:</b> 0
    * <b>max val:</b> \`SVT_AXI_MAX_READ_DATA_INTERLEAVE_SIZE 
    * <b>type:</b> Static 
    */
  rand int read_data_interleave_size = 0;

  /** 
    * The AXI3 protocol requires that the write response for write 
    * transactions must not be given until the clock cycle 
    * after the acceptance of the last data transfer.
    * In addition, the AXI4 protocol requires that the write response for
    * write transactions must not be given until the clock
    * cycle after address acceptance. Setting this
    * parameter to 1, enforces this second condition in AXI3
    * based systems as well. It is illegal to set this parameter to 0
    * in an AXI4 based system.
    * <b>type:</b> Static 
    */
  rand bit write_resp_wait_for_addr_accept = 1;

  /** 
    * Enables the internal memory of the slave.
    * Write data is written into the internal memory and read
    * data is driven based on the contents of the memory.
    * <b>type:</b> Static 
    */
  bit enable_mem = 1;

//vcs_vip_protect
`protected
QgL<L)4K]G1gbS>G=7eF#)a_E;U^M15B]+[P1eX;]>A.;1ecQ=e_-(Pc[J_#F)_Z
ga>AL0-cB13Y3B-G><3IK3a6GZU0>7B8.:>QU2T:aHH=(G5X]4\U.6SX0WRDAOSb
KR(UDEMJ&&=IMGIV8G9J,(NL1PO.efUJ^QC+#QJX\3Hfc(P67:S@HRA.?>U1J7<J
UO;b6N[Q?(R-dg<M5Y:HMKD+R4[PNPVK.JJT\V14=##WYT);fO-aB7(Y6ReY\\1R
34L^C<DQ&,eR99HHK<W7@VO9\O9ZPCUY.YS6QZ,GTb/<ObI+4aM@C;dJ\/fJfMAa
E2].N\NZ?;PgJ1?TEaE_,MC-Ve52cEPf>M_0(Z(RA-FTV?W6dI@AgG4SJILaY0]e
fURX5&@D#J3\Z4KAL_3I1#[=^_dg8b(YTZTFbSe3Q+?SF80T0XJ);?Oc#7+JWLU#
HZWR-FIQ;^85b)@VM9aWF80>JgORRA@Z81^UI.X59[6C&N>aZT0W+1f<A38EJTK^
V(CBV=DEDB-e@+86<C5PBUL,503cF=\c7-ZDPa8]Ue=W03-V/FIY.V@45/OSHCH&
gY2;;fWTF(Hc;1?5BV,9&,=d1I8NM/&XdVE84E/\Z#H1Z9ZDOA(0/g?a/S&IXb&8
a?-[Y:.>=:PPU8aPeaU74.C,ce,K15bUF3K<E(:;=2_LI?J20fHWINY^[M#Z\fW1
^<\)FYbD])+O#A2GTJ=Y>M.fb(fOS&9EZY@#bB2UA4BH0^=F,VZ4D4#>A/aJB-S?
H+e(XL-1F1(5D@Gb_f-@;FX^gcL;+7?_I&VN\(EEG9FYUC83fWc(GCWAKT5c_W<Z
eE8cHL_+D_<XcfZ,aZ&7C<[WY-dJ@C:38HeQYL52aD-EQV8+MHW6E0T(^;W3?e/=
e[#d/XBacbI?@HU^.URFaIa,Ze\[a#fSV<JWE55-^GW4f2:7#,NZCABB(E\fLFZ7
+BY0=&0X[D^fdfJ#YM4RZ#RRGRCMI+R<YG7/c:b.&P^Q]g#.SLPeZZVM^3:\(E9M
_];.8.1>7DZW\I;DS8,J;dRKf9f:L6P0,/c)[OT6EIBN@E=&,DDbCLMXG^Ga-64(
NM?gHf6P-V/PD:HC2/Me)@3A1Td089:bBNDe0)1MT1(Z9<U>RNUCCd:NSdQN>aCA
687N:---dY,:\IZaO5?[2_C8SETF/NF:M\]/DG8(e\[3cLSge@LVU^/[O\T)TL,<
/Z:A8J;56gXA=3U1(]#.b>_:-TO]J=d5P>3CW7dJ3)fKOX\J_eP6U+76K-SJQ^]+
H7gK^P4?3J.386(fgQ<]KgQ,(<P+](HI_.^@IV(,57U]B8NTZ7b21ICC36=-39G0
<[GCQ9^,B8LBTa_>bCa^@J-A792f)-\cQ>aN<\e7D.F<bfYQ[;S0D?/[OSBHUf9U
[+J]#KB+2#Aa<5KcgRC6MY9c7OJ/R\\]PI19L<YW_8^3)&Q>L/9@(UK^I.X10:)7
=0S\,J9ePSeEW;(J9KX\/0d4G->P\/WA/9+>2e;b?+?L-=;><Hg^5>S3c>E3H?&g
HR+fX:?(>)I,befOK8&6Gb<dd_)5@C[JNK3WZ3ac9)d<N(g-H382a]H0:^Y=QX2]
WI_^fPZQc=Sf&]gNX/LJMN#(7PTJM^D90FWNaJeAQX?I\R/APUa4#T;ZX43TZ=G\
UAB8AeQ(VOQV?#]S1M<LWRF,-WN)KQUd:=7?9LBUWG9\^Rb/VCP4M9J.V\TT-@(?
XfDCbgS_HD2S7DQ];0U+T9TFG^c]:IeeHC,[FVf[,R.HY1V@(C:>23\[c6HW2cRK
K)^V[,VeU=XR0FL5[g=cN]QA8_/.aDd=P8aC<JY<Q98^eXRUE-A/G+0M2&0D+#CB
E7WS_S0d3CRC]A6S&c-TY^bC0S[dAQ+.b^4gG].Yf-C3A,M:A/M-])+<b3CaP>)R
aV9;<AXQfHcA+@3;bFGNFL;7)\\B1?3:/C9<]S(&1M9W<QF<MeO<J@WKS=bbLG?e
Ec.WI09;0Z=B:[R?B]\392T1(Cca>L)Q\+OMBG[#g7dVZ@.YBD(FD#^A;VS47G0Z
d0a1^Zg)-1<[]:W>21Y1Fg<4>^UWUHO]2Gd>T);F7;MTT?3&NS0NP:CIB7M.GO6c
@]\d@+d,HDELgA7B[<6[XD9XEb/ZI,=0LX:W8/G9N7I,/N+;W;UV9OP@NW\YB/UD
1L67+Y3\8,ATU(0G5SSb[,)9W7H1R.+N4A.T?E.OSe(DPFR/WdV1H^JG3#](5VYJ
K8b1\&YTZB9VNC[N:K7cWRJ/Ae#cMT0;g@2d9_?PUL,LUMGVKFY-AK0WM^JN(&CA
E2aS:L>6V_,;T]cT\9XMf4a<@=g[=(_eYI/M];d9D^UKSQP2XO[:C\\6>a-KFQ)P
9=a[7DbL3;\>/F__OYB+C.-68Z:0AN==/YD58EMYBA=4Q\LJ<gHLF5+X.-D<K/FY
.TGVJ=Y3EP/0TK<fT)ECSD:8eb:QE.S5+7,LD,NbHMVYJ/UK1,O35?bS38ED64/:
cATX?0FMe;TRY=I=#KT=]L^O:/gND(=U3dGMVC2PD2O081CMJ87YNY8R;LV<;K?Z
5S->=#K3\3G?V+B4WB3+5]2]Q.Gb-R9gW8^PF4CNR?JWQ1ZgKNe0gJ.E[<XOAU>>
DW<#A?EB+XT>be^\-_G-]A+dI>97baFe5<Kg:QEA_CMAJMgT+G[YRK\e_R@:9TF+
<#>,8a^gCLd:[WfLNDA_#)]b;U()HTc.4.1.-I\[e^3I4G:S7H^2.R)(334VI?G2
?#UDW5W#3T<5[C3bO&JaKgd=WW7M-GQLWL#M]3[3/]5VXD+M4A?VL:(I3aAeY[MQ
Ifb++#DI/DC5K4>3=-SJ(J6=,F<[88<?,N3gGcd<a3[\FH)\^#II91CB(VZ/fc6[
HRIYVESZ@X^TS](b6&C0RS-JPM+&VX9]fW0APT_LR(<:X?BTF&E)30.C5eP-:&./
<Tc:\cM),9X;43BU__3abN0#:DT^TXO;(30cbg]]d^R3H(]F:5Nf1,P9BRW:1E,=
+O@J@,GE\Rd#/^CEMb=\;[8FRQ9KD.U;#SNW#/P;O31R4U3:;S2V391g2974SL[/
4>>NVGI+;E6@AX;.+1.GK-2>M3eYY]UBI0Z:Z@>/4HX70B_4,H_FW.LUVH>]aOB;
R,>fdSf>X)FeA?Rg[(J^DX:F?2_?Q+JJY7MKP#I/-.G5H_(RRY\X@&3X2N[S\5#(
(^KS[N=:^HMF=MKLH-G5UeeY>&f46(cWXc5FL12X097Y[862aE6RZ(fDP[UOPT]D
?AE@6<I#B-1DGcK/eBE@1GJ5U-UG+VT31WcFd90J>fZ6I6KWN.Y]-D@eNAe>@&,g
+Z>H/\<:61\NA80bY8>.;N<OOX=Yea7CGNF(^S7B].EB-48(3(PI,cdH(fO54=ge
<]^#ggHPVgFDFWTFZ8[L.9_]@I3G<L+&_NC7Q&KN6IG^Y1SgR<70ZHQ3T^R010,H
/)A36[)B&cKV,^ZJBZ_g-(B2E/3UQMRQ_:+/_TBMXE7T=7+48)+@2=#\TCQ\-&)F
Q/9Z]VM4J2-Q9\[?(HO:>,P3H>OEbK:)aWB_F96QMM#OJ.4>a;,>FS(W/6Q)LU6b
88,,^P5F#cL1Ra46APdQ<e0.CPE>-2?b.]5/^b_5@UX1bO2K9X44K&OP]QOZ:[N-
3bP(JK0b]7=&XDgU@=)#F/6KQ.J_#+]d@U-IBRUSa(N5Db,KaH9aV0DB/eMEaSG]
Cf&)b57NDg@BR6QJZ5=bKNe:(_+/0C)-HS0ADU&dVa:\bKeR??E]17&U_MDO>\eb
A:(^ZDKac+@;b..9+S02eA)M0eTY]&.UJAKbIeMBJ<.f-O3MbBFG#W^E&1VB2D4<
=W\BIW2-:HaFF(M7Y&9W+AN#=.;]HBTIUM66(7TNSW#-Gb;/7O6JYCRP;bMWA]bd
GIMZfcWJY6YSO;=[W+H_W/#+YgGYYfM+2]2Q=0)/^.X4e-9-,Y)^J55RD5(KOMM2
3Rb&^ND(_g6JY13]#:F/&VgAXG+R99L4eKM[#aH.Z3:WU7>+:e6U+E&]).gEIcZW
>E]GY0LNQccPL/b>f;#87W0JZ9H-NP@UeIPgIQW_\O8Q&M@3>bfS2C<M?THU>LcW
]HQM(.F[JL^W&O;[ecK:eR=3A&(NR&H2KSA@\8>E\R=a59PU3J<bHde:Q76490Y(
O>[)[8LcW1]#W=VdIeAHOfE5=8Y@0c7LZQN#CUg9.gG8L-D=S2&4\6[._N3O5T^P
BeI[>]6H=^fJIaQ;C7RW)9?76aA,K(S:];:4e0FCR\XQAg^,1C?3\U&IKN6FKU3I
)>B/eTVX8dJ,F5<#I];)O<UUgdV3(+,,ZW]b_2/N8EVTE5<H\)0aFD_4gMfCb<V9
g5[7_;>f:WD;ENY:=g63J41;ZLOYg1e0a[1H\._FX=-[Ag+;c8b=Ve_4K$
`endprotected


`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
  extern function new (string name = "svt_axi_slave_configuration");
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
  extern function new (string name = "svt_axi_slave_configuration");
`else
`svt_vmm_data_new(svt_axi_slave_configuration)
  extern function new (vmm_log log = null);
`endif

  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************

 `svt_data_member_begin(svt_axi_slave_configuration)

 `svt_data_member_end(svt_axi_slave_configuration)
 
 //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();

`ifdef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind. 
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.
    * @param diff String indicating the differences between this and to.
    * @param kind This int indicates the type of compare to be attempted. Only 
    * supported kind value is svt_data::COMPLETE, which results in comparisons 
    * of the non-static configuration members. All other kind values result in 
    * a return value of 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);
  // ---------------------------------------------------------------------------
  /**
    * Returns the size(in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack ( ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );
  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);

`endif
  //--------------------------------------------------------------------------
  /** Used to turn static config param randomization on/off as a block. */
  extern virtual function int static_rand_mode ( bit on_off );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );
    //--------------------------------------------------------------------------
  /**
    * Method to turn reasonable constraints on/off as a block.
    */
  extern virtual function int reasonable_constraint_mode ( bit on_off );
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>read</i> access to public configuration members of
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  //----------------------------------------------------------------------------
  /** Used to do a basic validation of this configuration object. */
  extern function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);

  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern do_allocate_pattern();

endclass

// -----------------------------------------------------------------------------
/**
Definition of the svt_axi_slave_configuration class constructor ;
*/


`protected
5fd,fNA+-)&FLW;7(&Q-N>I7X(O4WLR[,H5R2A5I;2+WQga.5#QT4)NM?(P5d+fV
(J;?C[XD4BA8&cF^\J1+]_.1Q^WVB41X7#XS0H^B=@[81N]KW?5<7L,TJQ(82A^7
#aH_Rf,bO^KU)X2Q?RH@)aJUG-=a]HXU]>@b.UH7D]W,[P1NVe\+G[cX(QP]V4<Q
1DW@1SJ7ec0>K+<^QfV2/&J4L+P[c&VHNK&Gde25K82c0b9+M:c,OQK&-<P/Z@G;
GfaWWQ\S1@LUMbF(_Kd6CA=XU&Kf]0(Z<^Y[9P\6<\2d8[@F^=C_\Y+7TVe0N6?_
fCWGD19?[Af+Pg3:GNADcADSXC;++RR<f\K<1-3/eMK>59<cX=T_dQ+IZ5FO(KQ1
2@&L^bEE1J05^CI]:_39>_P9J]+I@JW,72B/C@a3^(R@WVTLOCd-^^4ZAQ6_[XR3
T:f&G=\-A^-B@Nd9,B/#64+M]E5P61GVIIFTGYS5A<LMOZg#(2-9<MKg6&5Ea;<Y
76DD9A##d3ZM66H4YX];Pf><6G;?Z]aA<MVD:ddN;K4^U+MIf8]aC8_HJC#L-gLd
#=>YEcI.K^3L+9D@eabD&e#V#MG,H(WW@^4#S\G)Z9ZYbbD0Ta[563\FO0R\]Q-1
8&:SLVW&[7PQQf7-<,;L,).M:G\_A\P/&F3=0BEOf@LYF$
`endprotected


//vcs_vip_protect
`protected
[:EUL[2PN;61baB>LBKB.-329(F&.:6PH^69.+860XHZcA4Q1BAF7(01fEJT__N^
<4Y^a)+R+Q_OV9^2Z>]MD,)(D_:X/649F\<PZSRd5gcUg&Kg07gaO>QDQX&(X//c
d5B/,A]MSMWG+Z-2::NAbg/FR-YN89T?Y,\aV+VP=S,(K/ae9BL0VgQ;&GA?>;;7
KJ?HQ_Z034EGFAKG8c^Ka36JR-&<>##ZPMa_U]0a<H4-47<eTVZWaG0EfF4LLR=N
&L>.f0_-fA_P5(],G2V=S55ZUEF5(f<PB8H>;N7bY9>cHQ\7BgSc(f-e[Y?EP79K
]5A]Ge@@gCgGJU6Z=1Df]0A073C@2);WKSM#SP<=>>@KSa=2P6).DXM-YNQ5,U8[
3/LJ@O+@-5@g4U,5,T+?c\6(;O-J<a:UW;M2b51U:[U0?ZJeC:C,.S7NU?#ca=5H
;SJ3G5bfTZ^,eb_WHbZX9-GEDe@<Q_G<1M0??;^E+ce4=#_]RSd44HFA8SDSa3F:
QMb>G32c\O2?T)Me4[[?XUQ\_E3NA&\,6)E)e3\?N>\>IT5Xag&258WZ.,]_?gA&
?2#+>CGP[^=LORZ6M0VPCPI?KBM?>S0,5<H2I(5HeFI9BAAd&eMcE>O>M7<VP@3[
V#0Y:,He(@C@<-DU5:TG0-->S-YD;,F)FC/?Y4ddZ10_=DB_]\GZB\S,JQB[3Z3N
N]X,AZ;G^K^5dG-e8.NZH-HH>.N]R(R<MIf3c#1^&C4GU60a4G0W._/2^0MKdIc9
C8PT57.T))@FbaY9E3:&fVIUgUc,X^3HV1:fC(THG,ZT:E4:d>R^[5Nc;=e-=HP_
,?Y^/cD:1f?B=TY_G?(H0_M?&>U&QW+E#0:HW53J9BXT62?aZfDAg6/H7F-7V1c.
7.?dU)>B@#]WW2D/6L.J(DHZg)R#,YKHeI0fd:GMK32f^0eV/I79b^SD<T-KBg9@
ebZIE3WFJ.[M#^8;RdS&R&&-_:d6K^J;Y<,,<R^K)_g>OXAb:WY=6&F<OW]CU52;
&^CdCW^HNa)IJf;M#CWHQ:5^_R7GLE<B.Ja]8FMYT.f^R.(Bb3Jf^NbT)UaH3&2X
adD4I;,B^-cO(=]M4BQA,KZ&0D+XQIS@b,_d-D1Y0CGVB3c8>[-?@fWQDRT^9C(5
\2NX<6,/=^C_^eJQ/>_K41(:743Q#?B1AN4;Z?=R#I^(AgO316L\X14Z(db9,0XO
U[Zd:-L;I0A,#UPO9Gc9;<I<cPQ0CK,#>)-RgUSE7Q)7<\A.39S:d<CL3JGcW,W#
]b__e[d3e?Pc>\;.SCOH+F41ZG#Kf_2BB(<)TO#0_54[SA^P)gbP.SCKRUKA\bDd
RF5Y\CR>+229]088JUA:Q94->X\#/,aD)aJSE_&M,=;E3F4JFTS,8T<?;fS/F_4R
S_Q6b0A:g#_b?gCW>Lb=&28D\R].<[P,DH#-XHb.V#g#7<2SbACDfBK9@8;=c.1a
1BddCM?N/5Hc,/ZVV\YD5\TM2;@,6f^K_W13+S\<FM4?=gDf7)dI[0K0XW8G\N<F
CfbJV;M^ZZWZZ935[c12>c@-J@>U?QPK.ZR3EY6E/570&Wd#0(,Y5.+3-2NeH-ND
VHB[,P8BG&,_Z7&AUd6:^ePL-B4.7X:_M2^+DQTTH(6NgUK,1[Pd=7Q251872F7S
d>7F]P0#X@)56OY?Qc(588dCJ6a2RPU?XJI2)GCa94Je@[J;]4GFbFD;1b:1G8Uf
]g-_OD7FBb]UJN5Z/7IA9<1bDb8M@b)>XNRBHLI)K<+F2Z<WU;>&&]5E=7ZSFa^S
+\,IW#Kg:Hc<;LGY#:2Kb;a+RJ30_.fZGSRX4A;3UaFF3<TQbd<4bbbc=^4B30FC
D0;F/V?[91_\QIQ5V0T&E9LJ/U4.+W3IW385YIHbV^[O+URZ1aNSe88[\K?CT7EO
aT67=DaS;e@eQK@eW6Y#2Y+S-;^8Ha)fK-(H<&Ma0:N[U\9;b>P.2,HM+K5_6DNe
.ad2<?LRfMI^]_:Ld,N^d7LXM:P2/b,[WZ5AFG0DZ>c93]XWEc8g<0>?.8]KU;Y6
0CH3CIN(UUKQJK\618&@Y50:LQ[5&d655RQA_1dL5?6\d<5Re0D;FC=PaC=BNHE7
X),><7Z8<:8Kb\-528A0d>?I\=2Tg_WU(F+SAe-A[A/\H-9>><@8@g&8#+gQ=YY)
<.(4,<MHF98S59L^MHBgD^)^[,&cEA=g?c?LFFS1.37+1QA+,AUM>C#>?,G4W=68
1D?(4FYZGa]eUGW_9bH[5I.NTGR\d.[CPXfF=1g=)41KO[A+c_@,TRNe:OBXJ?#,
5G7@;>-?>KES<I.g\+d1@Y<Pb_0_V>V:Z<#<+YbDRD/JR5FO5Y]bJUX?G:NO9<0,
_/?EZV@Z?(]\K=#K2\S1O?1ScRT1PZ#@]K)bT2@5P5CYF1Y&B1eE:+X-93&GN,58
?@,WcC-.#55D/f7T6)bOFF4gH:,bTOP59Q^IC=bW4gC9D86;)_:4Mc<(]6e,3;/8
XU>.1?<5[MNH9.1OGRCWI@3N.OOd1W6,3Ya0PP9@<I8JQ(eF1D&^dH4JZ^W[_.@H
UX;.E_;T9)R>O@(^&T=&@6RAJ][W<7(?14<Xe#<HCd]X#b-K.eUL@63CT-W@?eZY
B58_f(:B(V&T8PF_LH#B+/JH[I\](7^GOQbRHe[WHG<6YVgKOe[N>U76_RE54[eb
B-Y=B\W23Ae:X6[bB.9:BEY>W\QZT)fB#U_TNFL8+VO@ca?6,b.6@5>J\1>C/_@K
<c=7EWO[7\YP;-]a-?geaECD2[6)&RcL3I)Q7C3<?gGgY+[N7f/6QFBE\FMI5dG1
OS\;(fcNVE0=(O^>HH5.\KRdef._f0>@IgaY(f[U52T,)[AH<,7)1\-63S?e/Q4H
g-[<.FNg=F0][[([_40Od375\03#QIdAPdC5.D>5K0FAI]cf?S:_3WW8XK3.Y[Vg
(@4,78P:_7T1-F.=&f^gb).Ig[&YL>[.RZ5eW4EZeNdba(eT04P@d[CIWPS[>PWU
3VUdSXbH@1&[:-)@7OXN&aGU44Q&c(WXO5LD8bF?..CYG>CT[4.(a)\:]#<.\(b,
W3d&IgP=.4V5PfaJQ.(PDGR+4&RU/?P#2V(<,4;>NFcJ13L\SYe.9M+[T]f@S3=3
a.eJ>R1U\VbG=35=I9B:5;^T@/]G:DBZ,6R>:+R#3(]4Kc@+RFYb>)WP4_MXG2N+
#6&IZ/A8(ZXGdV86@Ya:\2Jd#cC2dHVIL[cM1Z__Ff=7U8R.Z,b41J.A_L0-e1Af
ZO1g)-D>GaWTf8_gg3POO49(YG\:&]2ZN[T//I3e&_OIF/.,PN/VWWFB&M0I:EWM
c4^>M5GOW,YK-Sc.+/#A96:DPD?8JA18=9,0e-0Z8bF((^-8a:]-5;=b2WGP]f[g
@[gZJACYZ/B<IAME=cA02d(PF^L_cKDdQ?2YL=geH4Yf2gF-JLTgR>?K.=9EO?\,
TQFeGH3Q6f;CT5MU5;58^G^.Jc=KR+VRDLS\QW9T/>-4>9G&F#]8Q18>K6:\CHcT
GOaOdO5.G.(Z1GB/F/ZL-@cEb)[O5ZT@WT,5.L=;0G5e(2aIR9Y[Y>;\4T]B=OM7
V5eWK/<B[D?-+=0)C=>L2GD0PPKI[a:<O(V[H\XHU.WGSRW54GgJCgK9a)XFBYVR
EO3[U8]VL=8A7Z]?A6W/_4,HF_TWMH#NU81[,AN]cKNeX1U]\W.6VUTT:eN?/9eP
eP_1\gWKe3NaWE?1)GaXN],U]W>a)HG4TD&GRBDT)<?8gL2:eKce1]Gg38>cDfe&
<A(A>&a.=fD;K]O>SN2S]R-6V8Mg?ITC8.be(bE;KAJJ(FK0[3>^41d&dNJ1b?a2
9Ac_[Pb#-==^=D-.,]e]>1bWV=f)gG;KbE]#<TQ7b=GZ^2_6/T7NYQ]:O1K=]AWR
P;6AC)7T=fgLEEEUEKLQgSHPJ]OgWP-c\AMga&AeQ7fQK^f=)a:S<A0BLTDW@#QK
c>D\]gQ3#f8V2:?+49:beVHb9I5=8:&PJY,B<J9GWVPgeDK@JEK.>O5A(]YK@,RZ
^N&HfQd^K-6\Q]gBS62O,^S7=(4,EaFd_g?X_GRfg@-FE),=IQ&@9Xgd0];J&C6)
>Yc@6<ZfM&_;Dg#b(d/6/25I#T:)=Lg0B.UK&M\APg#-0&SCRO70eP6LV:d&7gfR
^-[I@NNRSLW11@g\23ZBGJb#F<F,;?gRc7.A;F#[C-9e3L1S\GEI8Z;2<MK,LUTB
BJ@:gf8[R=Pge]Ve6bdC[_V2W6GQ,=4NOXYF1_:,>-a7LTXIG2UNQ,EGLI;PWT-W
))HVfNe,M^dC@P[=dL+T+]E,L:NPDTHHFJG8N5>E<L\C??a3<)4)a6bFZHHf@Q5c
b9T_>f-G91PE.eVT7FPEcPS1[-G1PcCK(#H:@GDHbd8FM.R)f9E\^aL^1^:L8:4A
TRUQc^)D8C++9FI&/)4[AgAN4\68OF]<g#DNd0BEeaJ3dWcXAVO<SUWe:,B=TD\>
OH4[AQEX[PM^d,B[?DUQR=-1=AL6>eD\J5J/(H.1#3#0#HXI_MC??HYL7?GYePR1
>Lf[:&S>9NMN3X=+EGWR,ZDL>Rd]1,@6eY._72f646,Q?=,IUf5aM2cfdKZ(>XdH
F&5&6(;\4F]a&b#OZ2K9//VG)L;.<a.LUA9:Y_ZITa=;aZ)-C7e\KB@?AZ3R>L.2
V<?Ea\Z\>?,8I0=4a1OFCdTF487-U=a62M1LH_[SP68g.R5=G+/,EU>O&E@fR-g)
,ZB\Q/6/^7OU6(C6=fd-TG4eQFYf(=ScW@_\ZH#L-J2F0Y@c[^-;LZ./f0B,QG@#
Kc8U0.GP:>f#B5-,N_R@c0H=.YB3&U[>SP.1aMeWSOJ+f6,JTV7F2\+2OB,26P6F
.@K6YcMLDP]2GJ+VcEF+@TEK-QW]TQ?CPLL23XBIDe&J.::L+)_?)APDS[;A\GT^
\X^#VL0V>f6(RAH]XCfGV/BR-475,>KFH^gOZ5\A4_9M/F7#=2J,)B5W<)5937K/
GbaJKOU9];#IEgaU;@YJC8&T-TOHS5Ub<@N#SXcQWVe&M8^H-AWV70SVD5-AFT&)
ea[TO)XgUC<CI28A[9Sg0R<8_YCCM^Y/-=g:09&VC7-^dM112:MICU+.cUQ1@@S:
\4e&CYb7[-#,5729JZXa4X+76dKZ#ga:Y.6[Y&X3d[Pc>U/QON\V6SaV_RH5>-H6
(R_dW(73_Cd06@HLEK8+];TC[-ZVHKe=>]?GO9?LAgAN\5E(;KK);T#S#1GGR4>P
MB-&,(W2cD3IdC_T=J5;cXOTW96/].YAM;48A]1<RI]-gS0^J6>R<2G]68M,c>L&
/&)1]GR^WSSOJJWfGG>(4fWZb81D[^L2WTMBe1:..3U]JFP(7Q/\8_N^VY>MG6a5
d]Z>1MK0FCBC7KRY8.f];P3ACLBa?8N/=DPb8>YX>]<[NH>4H^96^Mb,_A^82@2_
&Ua:7@,U<)b]=U15,DH@gW#IedJ8\1E]aJP)Yc5FCB(C_^g0X^c\V4]\=25BBbX9
YJ:7HH57.04YX7S_dCVg;5+EMPQ)a\a;cR[#O+GL5#C#=EG73PPF\Q:(_<Q/GSHT
BQRISB?D)O2FM1+Gc8Y2^KCg4fA.P4<YcU,IS3G\+(08XXURGM0ebdd868P+;_ND
SD2(cB?:c&L>;7;:X>>AY^>f4RT_&^^^e1@D.XDKgX2gOI+V?9,-8A@a&6C^YOfQ
R8/VN#GA&gDI_4O_F4[MKN0P2C@_f]GdA5S:E,>^(7FVd@I?QabRE4=f(5H39CNZ
W/9F^((1-5Z1E9Y^&]?.(#agE[TSFU<<)H6cb+dd,cOQ>/G++?N2_XDe@bUP&bZJ
OZ>WYIASY=^CR4<:#YeENM-gG?=ZO+UeV&N-2e^\RI3K1/8(1VWaY38@;GRTW89W
V;]IGS0,:cBZE\PL]c1Ne1;[\S[/Va)c7)OMV?Q6ZNK5\-F_N7>>Qf<HSe3M)K_M
Bd(GG-F+JdX_JY3cI224gIAD/Uc[BHFIaWHP#NY3(6#JPE_LN1YM+RQ19WFAHVQ]
T4Wa#Y?GVebX??BWQZ9#dH]9ADXXgbId_-I)3\[8bdX,S3bQf<)XJ20J-;&D0GX#
[.T,VfJCV/#g5OS[)W1X9\GfUN(/CYJgC6NAAQcM#NfAWPH2Q;(QUA6<,e\J[]eF
I6g29/6V6=6PfYc(Ne2@V^O8PQ9Jg\bgNO:.=QKCA:cVORAIL?5UNG2VYcO1T@V\
VXSEcAQ8.C26e0=+_&8T/e0H08d2&V(?LIN>GT@(_M@RSAHa1#?fGH.A-c<9&SIC
cVPcd3R.R<Y-<M-K68-,7)@E=9Z+UA)&>;Z9(Y@7bPHbX3@+S,BWG#X8&OYXXY)P
aQDPQQ6,<N#K)M5FW:aUA+b3H0#@^]77RaW7\.4:8a9]DH+O+)8E@dA4(d^>24;]
P^:.TE)<PVO(eD_,,14;<VdRa9gRL@+HMe:/3,F:RG)?bL8g,+,<AR<?,D.U]COe
)@-ECZ:>5>:-3,&=3P641V04dL;_4&2RNIZ^;^gGI5C\E7JN5).S_@6II?7I3a]?
]_MW)KTWgN#WVYUaD5[&+R@GFLC:\^Q_]gg6f=_bg.\.GfJb3K5B@Q/,-H&A8f#F
^gfXJ]BDYc?g-56Q<JZ5UG/.D[+LXaRN#eU@9;+cC>6Tg#IeYb?3;;Kd?:>97Ued
X3X=PZ:U,19VT=KNE?<MfAZ,+X(R8;E7M1_J6:(Ae]G[]\Y-Y&8gNQ8O=Z8L4RF.
1W>d136[TV38#Gf+QBg)U((L\0##=3F#&1<8][]0U0#+C@7G:-?aU@GQY]X-H[A2
(UN&NZU]_[&U>_,S=bJ,(.E3Y-g7RN4cI.XO:4DO2fF_1B43\eJ^N+C;87YA)F<H
1A6LDB72aOL/[H)U+e[a.@UM1(4<(LV30aOPI>_.(G04XIc+^@C+OGYEeaBDXBUR
U]F0882XH0bM9S,XY4[gEfZH(FAeaAHC^J0<76d<fTL)U.e05c#^M@F#6VaZd?8I
I+D_V@/XA&+EgC2ES=#9O\K>3WW4B^.6-4_]fYJ.e=(C61PBS0G9Ra^?(M#9/#Oe
8^7H4E3ZGP(^FQVXOdSNZ68?+WCQY\QV<;]^gN&1FK;W0M+1d>@<OV6341\9F_0.
73C[U.)#BGPJGgMO&E=2AMPN+^7S:+UFI_-&QdE8@1827KcQ#bPWW(/1LD05_05@
0d(-U2SQfJ</9B^V>KIHJ1dW5ZP8=P[HY_W=LJ03Y@Z2M&7/d-X;3)EaR^M#B^&:
<ce^fW1?c@Z;-RdS/M&-bFS9A]WG,b5K)Df=W6c8;9)+#G.I46EKX61^OO25D=]]
bFAf_LL#c[EKS4[aNKf5\=,)T:eKQ:X\6Y4@#6RDOe:4P(,9N?Z>8g,XQ[KGZ8&C
GW)WDJ+-MQ=2I6CB@=gaB+2S-](>4Wd</c.=@9fGK6G61R/J(@OP(]K_ASEdgI6=
B[33Z4PGTSEGX=OL/TYLb5JJc//\g6=0WTYJ4-15AO2B79d&45AV_AUQ,SKUH/Ac
RP?_cM4UF^Sf(,:[AM9B=IEHU\e^?_\aBM2J\L2KSHKe-a;/c41VY3c[Z]CJ2a6L
Q:YfWHb@e7+6R(9690d#8QDg\Z5@QYWZ\BD6QTU,Y+U3+^+7K&/6a-QIO@^e(dD?
3WVZAK,7Ba4)dKdbJdTYBUP+-JDU(A8K4,\-YKf:b?BcF-R^c<bZ(/15DHKSB+@.
GN8cX4IH=UQFF?>\/M8YE?)\TOLQOa6\YB/MKB)2SP+YDAHPZ?K\79F0;LTCe;gJ
K;[XTA,2^g-O)>GG>[(=V+<II^\EK\eFccFR^g4&K4:RE5V>eJ\#Rc>2]2@4A:C0
GNLX5d61U4e4HOWdPC5#(QM1^&&VNU+BHIW0X<N1ZV:O;N5eB2?(:D@NZc+R2+[T
<P)PdP.2^WDMe_+CU5(]dQ39M-I5,2Z7Z(R5&#_,-YgU#5YYI[,f\(+Z^X.GbVU=
:=\@/ZU-[8f,C>8?3P;OKF_2\3QP66e9J@=eRCR7.O80R([fS+H6ZH-=Xd/6G+Pd
+;G74>Z(?5GPR[(2JKfaEKMSdXVH/X7aSUA&_K.9YO0J2=<f9^(4<H3VBZ7dEeM=
&IG#([86<=FeGIZ_V[C&]=\7gMGYXGa(5P-9RNb^A/Q0N0aeOS<U3/Rdc@0M]L9/
V<\dK81>#LO9B97HTBI+6Naa1L==LDTNde&f;eU/HMbIFB/b()/+Y;Pd7WUTN0OI
,(1/aM4X@-&9H:VT@J-KDb]2U1@YF#88D0KBXcCf.a/VB:b3U+:XFC,PdFLQX?\b
[9@e02VQY?&.XW^cb[Z109L<.dSAcBIFc,Sd45=<#\,/>[T,Obg\8ROW+.60\(<M
MXUBVERF&NH^U(U0F.@X_00\XN>[3F3#8gZ3V:,Lg:,HfGJH5F#Ie1XR@9^D-#I@
ba7<8bU&,3<Aff0DN48(aZQZD?fM>\CRa&IgfMW\UBHTbbT^WN]II5))cX:3d.+D
F^8d&+:,IHO<]2]B6=EbZ@VdEZgKR&OX=5Yc_O^&G<3QZW;;I5UELEXM(CM<Jd]&
OX^]eMY_-N,##a56B&_fHYR_dPP7LR:##0DZKQ^)]&105J<JI;AgTR5N_AX3AGKE
A4#RPCCY&a+9#2KL(DZ#I>7_59>T#O;6&T?a4-#+F4)3=[[-:(,TbOD37QY/,J4\
Ta))Y1IF&&JEaPB>^50;J4UVQ?.O>beYgPV<4a@A<JFd>^=)cgV;QE^N<LG147:<
5.@9ZXL^_gJ_fS9G_PPF3)>:#CgdE9#S)0H=0GL_b(eg/J(\KR0(5@[Q:<[(>V&8
^Q]4J5)ZRU77-8aS&eW>>M)[,;N&NM2X_ED8L[C\d5<++,TQUZT+4IPc>cR@A_7R
f2ba:6C\>7<\NG<7,g4?0U?WAa4UbPc]05FF@]P3&PGSJZJXDHMVP)=fV6/945Wd
Y#O&/V73KQ02L?/fF#U4e+2G:(P-&_K;GBB662N9FK.0H2@XY^3Qb&7&[7MH]b^2
fBAH]S((.8==?&I(HQ,/7[D?TU=/#_g2X&;BB7/+<:\ZBCRX],)XEY\JB<MG8eVM
PNC:OGY:]BR6aGWY[D/WOYMRB>8<g0-,OQCE?Fcg8I#O4BJ4Q3#9K-(bd8^Nc@NR
3E=C2I<c#.R<DI/7:ZgN<^(42SLCaP5W8\cO.7\VHF2V>.Yg73-fDIA=J,Bbe@J1
Acf.UK<-XN=^1\0&ggJ]@dY\6_^W6#:B6/])<A0:>KYK<0Y7IaZ<9/2+&deO\T)E
N>f[Obe=Y/d7_3A)#KF^)2X=U=#:B)fK6NX@,+0K^Z[(AX[AfEJ5-f(M<:=JFV:6
&JWIX]>f/?3(FLS3EH8Ca4;_6P04&7aPHHW^#]QGDP<5EV>L;7Vc\1:dWP<YC>3,
V#PQH,Ye>1_YKX8:Ud,?+ea?)e7CJIP:b^5X?EP70^faKccWBIFF7b^bc-\7_GH2
7H^;+852KbaaK8,7.C+bR0C^>R9IVcQ]M0.(Q,;I/_E2dWM-8-T@Z2I_Kf^2g7TK
<&1+2=)9O&O#3W=/^XV)e+H0_f^AE9cBdJ#UdQSS8?&7Wb<[/20K@+aFS1\X^GGC
@EUTL(.3YAW<;WMUcLI-S4YZZL]C\&)SZU-YM>@c?_6M79OfUIGY5(7YRS6a.fQ_
K?,<L++C3((PT#ebdd,SdZdI_M<P8bZdZ3#A..=ND;afZZHb.V-Z?Z?)]HD-64HL
Db\Z(QN5N&I\]9d-T)cZ25PX(58TMGHA&^CKVW^\B0YYO=WgY.(M.]WWaBE\R_1<
5#8UNK6d7IX5I30_U#3KePPT);[c(+T:[^3c?eSL,\K)9_=<A>XBS02L6<DWVeFb
>:QU&VGO3BGC:S,+P+)?XFHcdQ_(,([NJ+FJT6a@QUR?5./6FHTVg2=,=#e^.^f@
2&@B[MA#07cJFTS8cb:-f?fW[&@:Ic4a#QI(aMO6a&SS:RAC>[()A,/Z8=.-P@Q/
QCbU.4(WQRV_VJ3bV8eLCgM=O4<88SE=f8S?V3#TVCM/WcBLed26:I#3&>_I1URV
d23FI:fbO0FPI[(W;538Q#5T0ZLZ6E1Q8AI.YR&V[-HU[LMQJe6Ce^fEaR+eDR@3
MMT??OR(cKY21ZcEDUf2GBd\8]?6M6Jg?3XN5/_(g:ZQKbRR4fB4Ya<12X.Z>^e^
DQ9;b##]NGfL.92d8W);8@edUWJgJd#7Te4ID@KW\^5NS23<7@e?E@fMe1Q8\b>[
E9SH8O8QL)&V>/b.;^VI,6U48H@cH,E\[>)4Ic+eOP_XIg\A_)NF\X2b3=UWJ/Ic
fK,-b,VPIZ^93LfbKKU(]]@WP/\dEg_.5-]PU3F-^g0@=UVKb3BJDdfJFJfKF79S
Na\;EgZUGINPadY4C5fdf:7/8+,TFBPW_JZ6_O]C9NB9f,1IM692Q0D-UZ;g>KG6
I>N&F8=Ag?<2<IBLg\=\dG57SHMO?/LC-G>fXb\VEC@]/^8fI_#U>acA2b5EQ8>a
-beM^>T]3#9_ADY#\3UX(+MGA1(cJgIc^1dD5a,7C-R)b3TcGf>=a19R1]KJ]ccC
WJ0IM/-D)2M=:RaI?ReKXS((?G9#T:K;fNQVX@^-Y.DDO3XQE-05,#eU#\/6L7Qg
>XfX1F2MSTD:3-C(WM/6#B:EARS(2TY^A>SZZ6N\9d.?Q]#T6.?E;ARXE-(XQfb<
8[a?V+5bV=.7ag,WELMgH&@113])V^4BYdENbQWD:.HQT>R5?#KbM0<cJe4K[6XM
+e9QY2b?_H_?XNW)Udg^R#&&d4?7B96>a<=H@La>/9Jfge(]:8;H&H5Ec(E.J[YU
_#TE:N.KPgR.TK9,G=f;A/KA]KS##2OG^@adAH>X^:YY+;3@35_Q:GUeP.]LbPEg
5f:]Mb;D<\8?)+7/e)M_TW7EU#AaHM&1;POU\M^3FE(50NFZ(8OXXER#<675f,Nc
dABUW6MN,;2:EV&/ATH,#FM)Wf6A;_eD4)0L-Lfe?0d_W]g^fMUG9>dAK9^?-3P_
89I3,CTFNVNE#K(gELPc:PK]:J5YGXJUUbIg#ZUB0T1?98+=YB<a_XZ;^V4(Q6G4
KX5O4U^2H:RA@>,=1_,EY_;dFe4OU,+IIP-5dLTa/9GA>/W6+N8c,XK&A-KRBII?
FHOP8U^(;V06Ta1:[7]^<=QgI4G?PY^)(ae\d9=]f@KBGH<JF4>]R99UD6ZU)g@G
f#G;L=>>S46>2Y^\BPY-_0gDAPbG^e)[<#<_Q,P52:(H\G9\3bB-A&;C9aM/f@1^
9+[8YOc4];1?KV3Rc3,N,L^?</fDa)IAWd#bRD4V/+g8YdY3:HDX_]FMH4EVRZZD
6^gP+J,2aCF?&:4<e7OGKZ+[?A=(-/R]<BHJ3g3PS@6P[758/[=]:?V?Q-X\acY(
3f?_&I\5.aDMb[X9-X4?d,ZUPd.SY(AT&R(Ef(Tg@fB<ET,BeGLLY<_SKVT)J^58
N\bM>@bK[3:ba#+[cD5VUC9>6-1c^BdbV&0f)?3UV[^TW57+E3+J6+1&3I@-ZB2&
c)@6/RV7FJ?1;V>&Mf=5=1MH0;H#b3J(B)SG=BbQ_Ac1JYW95YNI2;SVf9V1U,HD
&V[\CbH#BG6&U=R9M,]<)+/X2[9QI\]De0^gL0L:UV6_P^B+FWOgAZd6A9+,5-/Z
HTD1a0eO<26E=eC2BLF;gUR8L>BB<53c&MYWZ92NA:X;[:6HV[\=K21V#^+0)2DT
:BCc413(?g:eg;CXLaXPCUSTce?RfO[-MANDUQ=2Q:Y7ZMP[ZTc;/<GW(C#_W^0/
HO^Q84E-1^<TW[Lf;FX;I+^T2Q0_@;DTHU>gRNRIC(A&&G5/PLad9IgC[0a9(_#W
[_+c1]#f014<?K+G:0-c/:@_3/>4?O6F?XU(JFM-gV;.R9T3[CP;@P>Y7,BL-bec
BacSCg+\^g5G?X5E(:NMS[O10448:0XSSAJ1>AAU&?O<ICb]>=\G0)<25-e+2\8V
eZR2=,V8TJDS4d\EPS?0L;9<c[R@gW/=Df=7>CK9LCUCEPFeQDTPPE^9A[&&31VD
O9ZaXV8?[0H/;aUF.7/(=NYFd(])@B1Y?:bdDD1C)0OS0[=Q5:5dF9AJ=4?^[H[a
E?PJNE9IL)c1-<dc&9F40JI_T-QNE=R@d1^29WC@()KQW]-4MAV&cZce:+VecAQG
E5.]0UI.D^f>a#:5/_)5ZGf1#d7:BOA^#Mc\+^Va/^3Z,TAUI,AQFIb=-dYU?LB)
<BN^:<a>.WG2-B4d8INGRA+c<a9NAC4GUa#YV3GU#If/[LOI]E8NPGgJ3R6+L-YP
D^M\X9&-7WbS(.UK\=\93;S.A^\;(HALf7C6aeaDUGCG3YKI6d4Q5MHgdFFX/\PD
XIfBVde1[/H4L,QM+Jf\4_4VQJa7MSZY3]DDMT-0]7[HAfF@<<O&eHcgW61^b;80
R&7HOd>@1@V63Z-)0T25=g[C4Hg=W,fU->FA(cXeZSXK3]GXYD5>\Db1BNe.&6Q1
T1gB^d//fU60)CJK))\DTH-6bP68EJa#I>Ye,J85V3+Z/:]AH##dede\d&[-ASRQ
9HHfFbOBT^Q3O:)&_U8C3T/Pb<M-I;(2Dde[beI,_dR(X=&-LS79F;9V,S8VU>Tg
+ba=C5:JO>DAT_ZTWCTDE)E6,___?:JXZ;Q8dC\gK_RbB7/7FXDY:8aeKg^2ZJSR
D7O82CU2eH7TAPEY#O/N^U^^,FK&9VIE2f/^EF47K+Y).;aYI/HEF7]9YQAXW;b?
X;[;1/V.5aJ@)3<_H<caL1/@KW1cd+(H_9[\6RXA7RNS6b_QFH-aRTLe#W)(;=_#
T?E-0&AA7F\S5Q(,50Db)S&168P0;9P#G]K&S@a;ST>6-/9eY#^T8aDT3RZD2dO3
4Of[/[-+06?aK7OW>+A8^7?D2I,bJgI(ccLO13-6J,B\LRK1R#O-48g]7V@M&,2.
M.&Y;KXSTV,\\X,?e1HfgTb3NA/cd?NNAbW;W+0M>URH4570FWU-Jf(:U(c&M:TA
eT7P2<.Y@T8PdWOYJX/NK5dZVB&.#._-:A7K-A(;=TO.99-X-BY:WEYEGeYP7b>R
<DH5:Ze3GIG>FgVHE6/Cc?=_>?5H)>;=O#OZ-^b.LT+6NO=A2T?b<OC5FZa^+YN(
;1Z6&9&,#\&(d#CE-K#6:\7HH:GX;+5L@ANOUf).AV?Hd&gX&AdOZSKSW7IPOWQ.
JCP&[B(@1J1;2AYE:C:2C(ZJQT@5Z4L^KE?aQWZe/-bd#c?\X&:MJ.;V&+R>V(VQ
bPWOVRAU^4RR;)\A=WBfF+6Dd5O;H(db\DV,H/&LBXCMa7)7[)C-KCZ4X1ST70-/
3dg,fAa=(.5)5=,;Y;6/9^1JH;WCBTC<D^bJVS=]?@#^Z#_X([YAM#_cP8FL(NI\
,K+OcfB2_Z?3ZX^I0L7SQS>e+A[WQ:ZD@:6AOI,&AN])0XR(aOGB:[_ITW_<4NGD
R,YU(,QEfM6RJ)?@8:NOO]^4Q_^<3?CB;B+2B4R@Zg5d^)fO1U+QE(7--V2cc1?:
0cY3&3.X);HQBYAYe)B2@T)=TX8@FFPb3H]Q6KL&]RB>Hc22.f@C1@6HfR_UW=87
M.WE:5B+?@[PFS21>b#L^X03,8Qa_(PY34A]6)Q_L8WL(W\:5ZNMGK4J=cL\4gcd
0>dY+^f37aW^_S7_&c/WR0@8cY).XX>^UO&g]^dKQOLXBeBX08c&I@UX#N&g?c9^
aD/L\\IW1e&Gf1;9G-6,Q:,0OG/W/OTNO9J@d9&d--,a2I6M@)8V6@WS=-OCO,/M
Z2_)ba41efCb]ce1M[;eA@L&_)NECN]aQ>=LM(39aQdB<Ke>/5=][+a?4b<Y.P_J
.)PDE>(.<eg/e@J8Lg,Z^2Z&KP6c0M?cg(Ubb4LR/=LafWc<8e+,KP8=/-a(3TYA
66Bef[VRRdb);HNe\W2=396Ha4:5H#[DM\=e\&)](<1f09A(0XNY2+:]WU:&V<g&
bO(?c0/ZQ@+6f>PJeOB8f0QEKD&AXQ#\I,&:1&CbQFE\eX^TeS10]\J.G^KZPb(#
?=_Qg;-VJ>2BDON2\bgWH,d@;>-db\73OVcXCX85<O(?_5DV=M9bPcR+<:Y;\+aR
JgY/S[=fOPbRb&9UW=D)(Q_<aEd==TG;VDfV],db--R3Z]GT][W]86fDFEJ,dZ3S
0^&Wbb6;I;2MJ]([#GSR)4WXcBUPg1/];1KJdI[>2=CdfGf7@E_WbF<#[+Ed<.;Z
IF;F)^MOe_cP82/VSeLV0D+12AXdU?05]5MH9f?8)M)Sa^G:9A,(Z_&g<&#G?2WJ
ZQTJ>gS<Sg?;9VU1[(VAG]HM;-4A:f2HTL1P&:K74W;:[,C:+B(3G0aHD(LR>MJV
_=85?#]TT?=93]+PZeH,E1BaA_KZA[^ZO^ORAT(ZF4JZTS#[I@eG:]3S=>J_\>H(
@G<608=c+/@T(T4[6T2(#?f1f[1JDcJ7O6e([@E\O3)F@g8&JP81[1Ee/+;OeEH;
=\WcC8=Pd_M@XK\8]_T44DbH6c,.cC)9[;(;IBF+A@RA]FaI73S1Sb3]+cb5=8P^
\U#^-O]-P(Ic,;6_C=Mb=5U8EdOMb7ML<H-agI3V<TC;>GFZeN)8M[N:FJB^/_C5
HO23IKLK=OH8TH\]D+PUH@G?E7RC6]1WdCPIAKeJ(\+=g_N-U:+G-)A\I0f-#49T
WVb4g@:&5N)<82-:+-;<Z_b&(\Uf-1:#1:;:=aWg9P5.,Ma;DLUP48.,27ZH5;Dg
7R22\E5+GQGJdX_geX,aO(7f&..;-+IQ3)RfMT#SN&;YYI^I81O78^QVBb>2JA._
ZQ;.LGAV2BL4CC;N.]e#@A=/.F:>95X.V6-QMYW?C>+-M9\[/)U:9I41BJ,D?#E@
@D-1fe6O&RQHRUFTaPQ-XQY]d+MA4+4dK(>H=>B[RU+F8Ve^gA\Ea6]aI^_&AK<U
Ee=G(N6ZCbL[4?QAPWaB-XZ9D?]V0:T._ZaZ9[M9U@IF28Q57cJ>.],H#18IN41L
;f]0FC?.g[I7K)^H1Y1c&O@SQ>Z1&+JJ4_2)b/0\8?FOg&Z/RP,X?9JbK^dH=bHP
Wc2R/:2\Y[&U4+165BU^I6,M4)+L@DBE\J4.c]M)QC;K29-AKTU\b(g;+Y#f05S\
J/b>N+OR#II:2U7e./;Aa<3.ZA;X@1ZW=P_GM0^bR,S@[F0TX[(M3Ka&W9C,Y[F]
,gPcCM8>LFH8#4.9aB,PbPgB.b@BE8V7E3L1A(]Y^^HWAE/9fQ74H62HV6.(^-RG
+e8Xb8KHN1FcQP0]20R:FeB[4A7O?;gfAJ#PfCZ9;/]ge&OQP:Q,7V7SRY_g#K[6
8X+MT7FAQE.6a=T-EA^VeQ01aE+FecXUDD#4T\<A=PSe4LL?JUePM0f:/VTX14:Z
BD784]_g6>CFP^RK[5.4<;CJ(5eC>3FeeaXRaIIO^BU\cKQPMeRdULcMHc&A]YJU
6<3H9JW:MXITEd;:I9_]Sg[L;OQf/;1GH2\H&)GZf\YWR0.)6O\2PB,0[N.GZ;T?
MXG9))9:;8+KA7M2PdBET)S&MMM3JR8aO_=6FTXB)NI:)FXOc9P)O&Z8eA<7bXMW
<@&S[J9I-bY?BDWYgYF;=gf=bbaBXP6H6N2Je)+/2,(EDI7TQeMN-Ac\XDfM\K7<
TaLW5HW-?1&L+1JdQd.A(3d;I]F3N,J8GHdJXOE2A(b<.DKMJgc/-W.VFQZ;G,-G
(eN)@.RgYQ-4D7=T&)NG#I7:HPHC2OaAd07-6RI(Ae5->c]\+G?7+,A4KANK_G+&
#MP(<.169&>Y-Mg&ePQQ@PQ@BL?[4(C/1]I^(G;TETYc^QXM&cce4gc..RGH15Xd
/CNXWW_S;?JIVd#B(_O4@[Y8R/Ug.>H<<a+<BK3D@GD@?9L?399_)d_<XDWJV^Xf
[KG(U,=?QdQ1T[J>W^LLY27Tg?d>-7Q)c]X5P0J#1?-==X@^+g.XAL>@&Af1Zg0V
&\72])\I8]S>77_/N.aZB2=ENY]c^)),7X^HG;bdYQ1<>(9\;#-DVe>,;-D66UF(
J8.VFJM9;;2b2,<NQDDO)U.-3\g8,5BEI[SC,fePK;,^(3@OL+,\:C5)VB3J1Vb4
2HE7^ZBN=8=,2(Md96_FHNeQ)42]+/I.9_;.BfW>Z)Aa>,=03GW]c2=34\#7S>_]
g:-:EY>/6<L;QJ[68A:Y-))8f,>-F9-b&B\__88N1BaHV&GUeDN-,1(Ra:E38eNF
da,CDWbE12-X6f1D#&NdBL=/8.9#[7T#Yba8ccEY19=7TJQU[MT4;&6Abc?KY;_W
,QWB?/7S@d.DAaW8Jd11N[@NJY=5c]E3P/(&C>2D(\1a=FC4,8g5Q0_Tba<7_Q>C
Hd7V7DA;fUNcPK,=3+&B;L/8T7Q]V4K^^S3J?FY,a9fXGO#d1MU13SV3b6,,gTZ<
@I]5c,8g5Y?&^T6eUV[^,=XK>)RAU\#Ra8b:6QZ@0HaA9NKgGE?W<5.e-<7aRT5+
AZdWP5NB?[@#J]ZUT7-gA7/^T9@;6R59DO?0L)9M+E=I>2b+A5K9IA]^S/11V;Xe
f0\NI+dMg=R9YaB)6+e62(WY2c2XBRSg@O@\)b8XQI:BPEWOG5.@a(>@6H[=^B(E
FG=4G\]KG:ddC[]HQD][aX#JKC#NdT,TcXVeaCJ=J:0ALOUD^[]DSHU4\[gJYV[0
=5=)U+Q(eHS5T@e\&GZD_H?&GOFL-2C>X,LXOPd)K9cUQ^A9.9F#\b-I^[S7\IHU
2FRcPg\_cH,a_cC0/a>:L,W\a5S37T7cZUQc/+PT8#\[dRe1&3IIf)OR7KX=).MA
bU\76dXH6[>6)PBMHQA3L]]B#=M4bEB@Q+eA9<A>3P<3PDa\eP<FEKfY37U1X1LY
;EV&bW&57,[_PWcOXZ=C8fY]L<V;/U6D&<8Ydd^+C<YWc=]O?51SC6H+Hg5,HOJL
XcQ\:&0\FGdTX+[g@FVTM39_J<S;d<8AZ:QOA?7TfL.NB/A+H#E>>W6&,=H@f1MX
6>f>5\2XZ@;>e,Kc:[]8YY4Od^7\C&/OCcZbT^]dQVWc&\/Mb@7JFc[>K.bZCA)1
MZ0:3GgOTHF?@#_-(#8L5;I9M0Gf,AZ/gLVHIOe6VVU+_FMYE1MbTSV:V[b-,:?/
.P1G0:<\MTc]EXLW3;2;d4+Q]O)V+CI<H3GE,780<V]Y+)-#JRA53Kd[E^5/5]:B
K2[?H5934Q<aWM+Ya5O](?LS?QQ_8?TW\8;OY1>7^S4<.]H5e)^&HX<;37IM=0Ib
SB0d,89_21DgdF]P6A>4>1G3bWf?TMD6+;/60TTf6a0XD?4GJV5Z\(,D^b8KY)Jc
,T]KT3,/=3Ef8+&.YZKF+deR;65MC5D3[K#80RZ-=S,4c4[]cZSg,X9-??\FQW4-
7<\1_Dc1UZVQbLT_@N;Cd?WNDEQ5[J2#+GCb[9S5C7<_\bb/XV^-HIAS8>XU,U):
=^,;=cH+MLK.DOQL&9V?S8[PR]bXR8UEL@?>8:25QeTP#,0GR1T:4)ZH^2]N-/-6
MJJ[H6MA39XK@.U<a@6Ie2)[S=Z]=+C2+b__?g^UIV>KQgSBMA/-&\DMS.U&acf>
MS8AG8.PG=ZI@GOd]b?G=MbC<#;^-2(OH5e=]FJ<,g65.CB\@L1SDX5>ZR#V-E)#
C>gd-+SYT/#.H0PFAS&]UZ]3@cPM6K]PU6W+?C6MOdc.[A-.6\6a/T,e,_T.>LED
IFbDC0^U[M1b[KfE6#+[J3--#0DYc3,8A7R/Z[::]L7\X&MZ;G,_Y1>VH-XAe2_)
5]^W[TM/H=SK-2b0eH[ECS/@YP:96eGfJgZL+abd]9Xf9JUJ#K7D60Wa2H5P(V^Z
gS&UbM9[=f\B:V+bf\X>8<LdSLKgg,YO(@7Z?;c6=SE-[2eM9O&IRH..Y/PJeY#.
6V5HNEa]VWB<URegHZ)dE(U>Ic(M>6Db,=^T8#P[bN(B<0-I/-A&0d3MPgLWVS9#
5I>b6>[_^K3]EF^ZS9A>)./;,U24X1IPO?<BL-QZ::&ZLK<=C4I3E>/K5d29?I42
=Y\D^OA(O?L)])eL=0^(D1<d.7P4f0;C<7Q<5bOeJXA)/bX<=W:C^.[?UdK5VeWJ
UU,JA[fLLJE1E-VS@JK>g#O2E5:6bBd/C24c^6YFC#^fdOX>NA8T\SZ/C1&.0cWW
&1W@JCIR2<7F;7(?RI&)]cQEaYYVGg;#3;@2=-dZR#c=9G^6+OK>R/KI,GdRBN^P
5^1bVK]6JgIOO>,&ZJ:YdV]Ge(VPJO]^AVQL:T1;/dZJ^@D]L^=#+bF7)RO>1/Nc
U,:DKG#N4.5U+S&V]AQ4>b(4AIC>Wb(9AU[U:,Be_N00JCJg]UK<YCAg?#0/D;a.
;LN3N,=P_5?T<161S3dBE4V>O>.^b-+5WHN,bV_#T(EAQcU>ePQFMgA(K886B,DF
G5eY19INT_N+K(;G&C;T7MP\7OT]Y+P/DW?7,^K6gH:K#Aab/VO43/<.:BK?/1f(
@V>ZCI&-K8C>)98C-/Ub@N#,g;#K<[,[M/.>gO,HAM3+]/)+LT;_W&H3+:05AI7H
1a@T>1>9B0ZQbX,@B1&[]NJUbLE)OVHaYHOGWLU2E<#M>&3,4N/L>-;?HX_^8HP@
,B7KKN+S(0MNQ+<Z,&8>Q]X:</d_<I-??I(R&HTJ#]7YZI)\C_E85SF9&=RI@DNf
+YB&JW9SGMO\.<?a<2BMHXX6TdF0NR/3fFI-FX.bPg5IS^L(^DXOT]WI(VcMN17<
=0_4e+0g1BF=-)gK-1]VMf9_M<:gO++(CVeHe4_7f4S5(X^@H07U@daBH#WM8XaH
Y+5.Z7\=-C_S^(fJ>S8K#@S0)H&EK1+VbZg--DA6O\&SLK#228XbDFF6H#FP8/(+
g-819#AdNb\[6:cPR)U]45f/A]RDH/CXGc&_J4d9S(0TE</]1c:JE>JGCd.:A1a[
.SE_M0bB0>U(5=0-;Bd90&L&V5M:Z4<(9+GTTRXX2A6>JVVc1Udf\a<E0g6K.;+1
Ec=RC71T)YY:]+O<9-RUX/L<<SVKP\AU&Dbbe\@gQE:RL4TGTSP]141T.a@f;bJA
M;OO1;420E:Jd-UX;=G[A>N&WYd^gfa]R?O1Y(2SY)5EH-K:[&Z04eEe]g96LW5A
fED8(eY64Cf5]PW;90SMJ6D@[cCK#>MR_&<\H6fTe>WUU8R)&)<KWNZK^GQU\4Oe
R/f4a2C_+&/CHY9=X>\HQ@b]XI^fK9Gec]W(0U7N-67744CRLA[aGf\(K>?Cd<LF
0:+HE-TfO:BbD87IM&@F3./f]ZF&ADRadC(&T@-Z;#cc:J20&gB9f?+X^=K?5X><
N61]Se/.,fQ&[E124>][3821#_O7:dCH^)T4T=/6F7g-]2GdRbJ7RF&U-9HJGP<G
G/#WJX1N.-&.YU11ISZ=#I[[\(+(Fb.>0O2Q<g3Y9V>\#&IJCcEVg8Q+&<[RRY1+
.2Ucd/0=[T5(A&5JUOa6ZHPH[[Wd3-UEX6H089VeNEdfZ1^cXP+,2-,^ZFcG-W8K
H\_##=3VeE7LPf/K]gCZSW>5afICFbY-,]G_46>IgBPBWUS59Pg,?JadF2_Jb[P2
>6?2UROKRFEKT#SZ7.QR+XMBKJa\)Ja.OEdN)989.\F;FgZ,-Ge#(#ZR,KO6(5@0
@1aF^^gMADCQ.^@^SU.+Y5(&W3\gWIUV<\][IbUVF4/Fb?E0B)3GBJSe+2?gT>)N
:]7)Rd=3R(]>V?R)@dT\7?fQ4JeH7VF(Va/a/W.J\]A044M[Pb28X8VPJa\4d?b.
E:cbXPZGAQab3<KW^-TG7GOP838dI+0e(<,CF/EA&7\&;S#bP)B<b9MQ;T9?<K9\
@997>/-),;OQK9cL3H/>N[QcOd_>H;7UKSZf81e;RU&gPAU:02gf9=cfCId@eX==
7QX,(N=:<>D&TY:F.DD(Mg-Q5e]?DS3<V@D?6E.EI&O,U>?J<#D<JMg,XegDGMfN
GT:Y].bNAHf^ODEWbG[B=_9[#R@E@#+-aLg=&&I=aY=+2#c9If54,/J7.Jed9B2b
BA3GeH8bSg=7bC]0WGB:#>..7Q^cb&;UNaDWCS&;-g088-N.[D:G:I7.1L<3^9WY
P=(bXCW&AQ[bbHR>1?4g3g<WR0C8&CNGcb2ITHT^<3I2U=C=W#[2JCFUL4Z#Pde+
4DXK.3R,G>C2&8;ZfZO,UJ.F_,D=857.1aOB[:)I,KGA,0;UN[6V8(Z5DO?R^)7]
#gOX,;=Z[7_A21T/_Ufc7^c[5W14[(=;@AgCGB-PYP.JB[BNgMQ6(&d_IEO;EK09
YNJ6AM[&8B>Z8T/)@M(JK)cQ>060CDgTBTQD#BWZ<0?7),eJ.V(d5;eK8RBM[gf^
]cZ^J0;a.Ja7PfJ7:LJ@TdgL2VSf5cT^&EQ7?/3>Ra4)fI=GK[L(F+7-+bTXC(+=
c^Z8;?DKGGRYYcT+c29K</L5[.[D[9aIZN3ebB)H<F0f1X/6_AE:AK>cd42E0/5X
,37\ZE3\EdVQ6I^R_-[U-<W?P>.IK9?MRbYGO/N@N/]>B^d)M1GIZg.ePUQ[<\SJ
W=fgFDTY6d2.<#^SS>a>[>^A>L#.)<ZW<7PF/^MOA_Tf7)F?J^6d&5ERDeLdZ4_V
202=bbEO_)VLRM2cLY4CZ:SdVL9(/D)B+TBGE2;fc0UX\1\A/0NE^YFHeH>E0\BN
<_3XS:S#Dddd,d+&(K&Dg89)Og+?9Rc00E&f4G-=)[H.:?FR<1.ZYQ]652)RI/e3
d1D@DZGF\[=TfIALW+XA^Baa,?BLI&RT.&1O)B3Ee?RKN9PI&##CQ&?SY1cRGXKT
YZ6U[+Uba/YVUP-\Y5994@3a-RH5@XS@Lf3bXSHU.4H348KQ.+.>^.+Q.E+K;\(0
J;?b@P&1gT,ZLOO.LG/RW1NN/>[OU+?JOK70SF[TR:(G\VF:cKQ=Sg9F&>GUUR/B
4:AR-H(g-2ZO8Y.?XcgEM)09>Zd3<#<2c1EQHFF2E/VBO_ZLONN;<3LL;SV4U;G5
8XA?:C]T#Q>IdM:>DVS?:d[OMTF0g,[#@eb+;-DVZ-(bTeENCOV32dbP3F&]7ac:
Q\282d\1/+&J0bdc=.&?=_D(K?H,TS4K4?5Z7T.Z+ZX=WfVSBA[F-I24N5>H5?Q4
//?CRCdT[fFGBXY:eC,gAE9#RcG-S2L&N7BH/:?Q>@]M6D-IYe>Ef[0f?)/R>Hb=
g#B#HZA2eRdB7?GNFG+7f#a\?8fJeddAb7.NU]MaS^::FF>7HZ^>Y4;a-<dcI)Te
/:LZD:g;;_Zd&.gK(@U#[#W<.+R-RNJO-I<\YSBM\CE5?f(W8[/Bf_O;eV(1;a^S
?Q>YfZdc@_f-,b\3KW^4VN;Y8;:A84@62E>(8Rc?=J>.NdeCF#&3N-?#8XcK;KET
4=D?Z.WNG7]L<MR1bb.DgOKadRH>)db3]dO\f.43PBg:Ya(<EWP^;L:,D-YA5=dM
S2OBH3<3ZC<1#OPO_7\11\/&[D^bXgSB_5S=/),\6U4_eZ6GTBe>F(d^[70#G]][
XP.9UGOB^B8?cG0MYM[RAQ-aN./X8_g1cb;3dSLR<P@I9)X7@><U&LWg,V3<&ON6
\De=K^>XQA)\WNBXYB+>.DS3=Kb3g[&=KG@6=(WObdc;N3GP=)@QM[8KJ(3_CeUa
gR^[9@B17I2W@BJ3?8M=.+,ee(S:[TQIT[F4\1^.^_OY5<220dXY.(fSBSbXaSG(
_1Ua5_+.])B?7BggT[DN]5Ve&4(6,(d)INgb-_0FE+>T82,4@,^&21[ZPcJL8B.D
IQ;.NA9/ebDA2(HZN5U[RWNV.K[P^^][K45??B.]7/5]4<=[@?E&bAS/8Q\&=AV@
NDL/V)L6>O(6QQc@\HHXMeb1b]?MB+<MPcDeD8(QY=Z>IPVJSAWT])I].OVgA5:]
5A1]&f5bC&[&EGF0)GC)FF\=[)-S6#48ZI]5^JM9Kg8g-1N(\TPVWMbED=ENgTXC
?I6_a>D#T/ZbQXX6UIMV(04cD<[),[8d^OA&C)O.-CW.X@(f<DaU@@S.f)USTXJf
dT]DNO_Ad#XOIQFB^AGeDEZ03#B,01&OQggYXH/RXW^U#JX-b3+3+>W,SS_0Zf9X
MI0Y:)9^aWd_@=F9_cd\;T06@3PIENMR2GdM?A2D?;6LRa(N@:Y38W].UIB\=S7?
:fDW<B_+1K9L?-<E8OHBeb/4c;@Rf_c(NT45736&a87I2B)680\75#gD@e^V?#gP
b.c21_<O+,<7Y&^?+a<Mdfb8c-\#FaQ:IS)93//(6?AQMaTY3W>H/TBeUb80Heb4
P:?;WG;J=Hf.Oe)T1H?BT(\?CMM(C3JQb-&2>D8])^[:;QeZCBI=.UcZK]Y,O?IQ
2DHVc0@)HeR)U6M<@d4_C?bV:fg<5GD<C17]-TS)&.]<5RH_;L8PYISMN,Qg/cP,
7DB@HJWe&4U@(U9_EU>K3F?^D)bQ:KQL0SE4GF,S^=LPW)#S+R+K7c5.g_0f2T^)
..Z?>D8^V)F\CcWH_WLJf/&SX9+VBI.Q1@+]646].QFZQI2]#J,c1GU:[4_^[\-#
?e2JPPWDQEL@TUW9<D.;_8=gDB9R5])K8FPKCVWfUKH6(6QR&U&aCI4)ULbR<a]S
bA-,2e8KD3d0=0H7UbIOb8SD\e&5Fe5TA#57a+R:G&#YbcU\:C1OJ^6/[?f8BALB
8f0c0:9-g3b[)W06Ed?:D??V8K?K+RZ:>DK[:MG\+,+4c5UZ)]^(S&e&d,D(]V#6
>U2]&U,A:e[PC8(WbQVNYR9DHBWZL>JK?&g\MfBP;PFQ:3CP7P9;REe]a48\K8MD
\?>1G9_-g_@[8C0Je@)H^.d1Z-DVKYX.&[BM=+c[>C,8UU>U-VBT(6(,RR=,f@_O
RRNO.f^Sd&QEU\=GHB740+F0cQ,MJKEGPE605R1=\U,EHK(Je3CK:T<cfd8;Cf[7
\;)=3+JY<E.4E.EceMY>1)]+1Q;gcdRS=HU,CgORfH+)0\d6M>5>MScVF+]/BJR1
bIO(<[V_,;]Ad23BD@U3/eXI/#OK[DfD)TVNFc;D.E5[W01L6dc5P)6#-;:FQ9U2
L2?+^SO?+Z]S:B:d1<K09;G+G2(J\/QdI\KE(^N\De+-X4F;5+W^:bWd#1T\1>9b
\&N9>6bHL3.QCL+<(L)E]GU2)=1C^]IcaB9OAGEFOK=0GH>;39W#??fLYORAF5MD
_=G?IKWebHV^C4\=//TDU)1J;fWA/;6B2)]M9;-KdSJ@7X1WI7g(^YBc-<6.#fLX
&&#I?1Z?P;gK3e<3]b=eL+R\@I\1&/BD@8DF;X@:@P#=@7_RMI6(L9AD\/Q3BadF
>_g(g4&4M3&4MLOREg0^>I9#LE[.f35DZ_&8EeaW#_CPNMd@FKT:6[23:94>XIG_
DdCc+g=d96K7b(U+Y-9f]\C+.6=c_^f+e#;0Md_ACR1eA-#9K[>ITWQB70)2N1-/
#Qg\0G\:LcC?.2XHa1_g3@1d[64.+\@#R=QKc:VIa\J2_>\?>R@F_cDS?3YPCCUd
4XRe.E,<D\T5NN8XS_01(U\)#/.9_7L@R>NT--g:[6AgKF2OX+D8<35cbM(V-,PB
X#[fZCaY5@5->_/#J;JQHNTN&A3(<+LULH-+X,,H+?P-23YR2_U8NcDfE598bdVM
YL+.LHQ]1+8g7V>-GJW#d.Z[[0YZfUQ_=H#;X1N)#HT6PbaO[T3WV>eV4D:/]R_3
(H7BU>-X&=Y&NW4+V8F(7Z=+_3JSV;V(H5PF8A676UFSSdc92-247dW>I@4SZ5a4
9V),_AI,Td.RW;9,8&?,CTJdg_II-7MAe<dT.F[bEH3+7O_S-IYE^FWQR=2AW^f/
-H@^8VBD.I63E5Xe,LcQRJgL@#ZIf:4\VdEX<7HcPSE@SOBK=)WUV87#:MVDP1,@
[1MG:<52=/-S27;PSgM\TSf7;7Q/gC/fF]7b<9?QUg&04\US7H4Fa:8-Xg283PbW
f=c-;<JC2:72<[AP/MeY=L/]).PM:XFQ0\H,S.+9L<;17bM)4OGQFN4EX3#_ZSbg
gL7YHK9KH;23WAQM_>T2B<,WKTA?NWX&>\0(gZXR_[+Eb&G,EcRaQO;aCS=VAX2?
_6>U2Uf/aZIN;5BdQ#+T4XXc;<=]dE]T_S<O(eWWMXA)P1&T)[e6ScG6ee,R6Oc3
g-.UJ2RHcVYNB=@7OP.90T[bU49SdbAd9$
`endprotected


`endif
