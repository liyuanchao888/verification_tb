
`ifndef GUARD_SVT_AHB_SLAVE_PASSIVE_COMMON_SV
`define GUARD_SVT_AHB_SLAVE_PASSIVE_COMMON_SV

/** @cond PRIVATE */
/**
 * Defines the AHB slave active common code, implemented as a shell assistant
 * which basically just converts requests into VIP Model requests.
 */
class svt_ahb_slave_passive_common#(type MONITOR_MP = virtual svt_ahb_slave_if.svt_ahb_monitor_modport,
                                    type DEBUG_MP = virtual svt_ahb_slave_if.svt_ahb_debug_modport)
  extends svt_ahb_slave_common#(MONITOR_MP, DEBUG_MP);

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************
  //vcs_lic_vip_protect
    `protected
6&^-W;_:BSf:I9NU,;_K,2LD^03[eGb)Cg1&-2LKD&]KSD:ZZQER7(51E?H(daQK
beG,\4(58O):FMKLG8,C=9Q+<c5V1]3-;LaXS/&C.F+D)5?<?4XU;2eF]\\G]ce[
@#_-J<>0U,c&J6-R>S;gaV)A(LC9&DNMUFTcOa-+L,Y1-.[XQaQ)?)W2F0YKb(X3
\X509E9e)(WPS)_TKb+7b7,A:P/W(I^[W[.eWF7@Z)F9I:e&JRLV>[0;)Z&[>_KZ
>ZgcFG@=3TM;KEg5e,9H-:f[O/QdUAFIO),K1HT5>-B9E$
`endprotected

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // protected Data Properties
  // ****************************************************************************
  
  // ****************************************************************************
  // EVENTS 
  // ****************************************************************************

  /** Event that is triggered after every sample. Other processes synchronize with
    * this event to ensure that all signals are sampled. Note that if a reset is in
    * progress, the reset_received event is triggered prior to this event. This will
    * ensure that processes that are synchronized with this event will be terminated
    * at reset.
    */
  protected event is_sampled;

  // ****************************************************************************
  // SEMAPHORES
  // ****************************************************************************


  
  // ****************************************************************************
  // TIMERS 
  // ****************************************************************************


  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param monitor transactor instance
   */
  extern function new (svt_ahb_slave_configuration cfg, svt_ahb_slave_monitor monitor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (svt_ahb_slave_configuration cfg, `SVT_XVM(report_object) reporter);
`endif
 
  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the signals which the slave drives to complete a request */
  extern virtual task sample_passive_common_phase_signals();

  /** This method runs forever to check that an active transaction with trans_type
   *  IDLE/BUSY receives zero wait cycle okay response.
   */
  extern virtual task perform_zero_wait_cycle_okay_check();

  /** This method runs forever and performs hsplit related checks.
   */
  extern virtual task perform_hsplit_related_checks();
  
  /** Update the component when reset is applied. */
  extern virtual task update_on_reset();  
  // ****************************************************************************
  // Configuration Methods
  // ****************************************************************************
     
  //----------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);
  
endclass
/** @endcond */
//----------------------------------------------------------------------------

`protected
-Q:4N8PT]/>Z;1@>WTAPHH.e?WEaO://8CEO2C=7/f6=E@[,1cK\3)g_eCS9A,4>
L1@E6^9UM0P)fLM-cG>4_JCWNDa6e-EK\c_LVgOg^BZZ?7RaBYbTTS83:[eC[49Z
+?BA<:2A_QbOJcEeI9PGHBO@_E=V6a(Rd8)48Re8L(;V2b&2BfS0D0T?\N1GLbU4
<>18+.aCT)&HMWQ:@A[))db_TAA]34gCJCG@J>AfL#:SgL_(0Z@2(+,BJDLAEEEG
54b?^F+M+T034M[?=M9bK;g>HgAf)HY;/C8De[LY=?29gRFg74Y7f,NaW##V76EP
WU9d)ZYPIGN+cLb2G&ULA@WbYec0U_Ue:g1O7dMe.6_]8:QI_/1+GZ>?FSOYLf?/
#HKRM-AAA,1MeH^)<=]WeTf4cBB15NLNbH@&L.cfF5JZa85W-[88[:[e7UdDQ_X2
4L1CY+D>OaUK)1eL+d9).d,S=F=[&QOAG#.F/OSXWF4P@54X]9+KHV&/F5#LCHeY
J95SLC6XLX^^AMGBRSA6T05VNT=S/EM)2[/.6BF:#^]QWFa=G>b7N_c6ZD:85GOY
OfPI\Ad2R,8TC[_<Q_6X+N(:PL?_Y2=(=<,Y<O+WaC=(\R7R_f?#d,/4O4D/Q5He
,#PE,X1#&2FN@d9KAaHT_GNUaPH7UULD7/2,=.<K+4@Q7f4S_N^QV#b3U4?5]?_I
L>KIHN/aG^HO8Z&3(PW[gF,5FUe2@\9&X#bK:B?=T7cAVJ4]A;?FTLQ#?P0IULbK
gV\C85AMScg5-[Bb_?IgCg^abW/&.].)LH/d#^R)=+4DBd2UOX\3bJ/-gR25.&QG
1Hab]Nd(=8W.eA[S19\F.YYBF5P6IS8aUW19/5)\a=LU>:SW^E/7C+T6N>Ge0LE6
gTb]a\(a]0O+Yd+@6TEWT0M,G37E.W=\:$
`endprotected
  

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
Z?P9,eI@b[B<XM)QC\f95]Q)N-e_CM&^gDEI1VHU.,3F;9_>ecg:3(cAXQX?7bLg
4HZe6#>g2[a5-7b:Q>\dJ+.RB)_TGP&.<U65G:3)#_;[2:NN&8EVb_VM5=IXK(12
V4J#e-)LKO5^PQde:g,F@,M]L#O:C&,+Mg<BLFTL5\C=L]BJ&KLPafIN^g(A9C/;
LI,XaZA9d^,4[E;B^DJ-fQ.M65UeSV<R4_:I8G0LI(<ca\UA:XOL[=^?_fY]5IWU
HKRAGN0R.g18X9/^b\>D0W&5fd98[7g87[UJXbIf_L#?aCeEJ34)I<0]1gb0U\PA
AM>UG/YCC^fAA1NTc7=fF[_;@ZH,fR^V=GP=#F_Be15R?[9U1+K(G_RbAFVbG=S,
,1&a(/Ge7BXeRVDHKS<4d#d14dWcgF^O&BCd6MF1\cbHGR@\AF9KbY@WIVV\(bU\
D8#VJ]fU-cTNDQY9a^UH0aNEcN9?LH(fO@@>#)G4-KJ#]6U=Ad</N#0(e<>;c)Zf
<cQ0^e?/@&4S8))ZBHJ,?=42.g2aGS>+T24dNZ+9WDEYI9TWcc6]/PTaND&;9BL3
gM_J2P_@C]:/0CHB\g+2]:@.fOO8[H#eSKLKS153b0OSJ,/MU]WB6Ob-A^NRQB8b
>7NR2dU]7O&X@)EQ#UgGa0f>>b8(W<-M7.[b^M<^_2f=c1O)/gb;aO8,fOO9d/#:
J.V7b_gD0[7dWbAOaS>IT?Qf(1=HG?e#H/dQ:N3=&E?O;8S4/_NIV?<=JN^97EGc
&SR=M[D_^<.aU]dW;a6P8Tf/E?f,\X,aX?ZU[]N)^NG0,D;e9BK[a@]4RVI0E?H2
a@67?Z[;N[V0B_.\gB2N4O06:#5)0)B1OJ_N-Q(JW]WO>>7.CB,S\+8C@B[OP0DX
af>KDU-)FeGC7RW:e.]c>L3[)MQ3WLb;fBLf2E?E_UA\V86+aO]<^E4/_J?M>0(P
B]@8:W9?3+@:/_<7cgL],=DgMZ4(/?Z^4U?VF>W[eadV=dOZf<RfDgc(+d]\M-1M
SQB=_J&H1/V5KJO3V]UZ9dB92_FG8DSSKD:IFc3H]0GNRBCCeP&;[&=[[)A_E<8/
VaXfKX>Z&=C@KQ(=B87fX,X)Vd:^05>&NV56>R8,Z3&8+0LYXHA-FQ(==abK->4^
V\EIAN8KRBdb9WK0[?=F^d]C/A;-^0G/2:cR(g?)7Y\CB4A8T99@+?X_#4>U(:,[
.FGH,O[6,;cYHU-bG@^f1d]B+DIcaP5NKB?JZ+gf<J?96-\JC=Ed_7[WD0CP&-@J
@.<XGQ8c56,]JJ1N19PDLfJGFELLZDK.7&0K81^/5.QR8C+Uc7?K:VY_\1P^Z8A0
]V@3T5V]]FK._]35IaRKDG)N/:+N7)9U;aSJ2c5,e#/DIJEE7K&=57?Q6.L4&J&G
4NV-6\>H>#WU\LGI8H.@-Z64HV1J5J3-&\1,D@[c1O_:\4g:.]0?6X5_JTX_22cN
4;QaY&aHZY;ccf6<fGd7?D=XZ0F4;M2#Yg6):<)@ENSKUg,YR/GIVLEJ]07[4af1
6.Q.=EMA]\M@H^M?Bed?dIfT>UEf9@5eH:@ZM4:8V6?H@f_dgU<)D?7VE)^F>?>P
>6#LZ-S@FAECM:eA-bfH(1(/,I#[WF,WC9Q^4)RI]AO2K]IY#-<_RKS\YW=X;N._
2I2:d15Nd<:NJ0VeZB\]PfD_):KBCH#FT#.MJSg4&3,3Z;U,+DfP@;FfGK=&_B)(
EaP9NGG#@W;YM<;5RJCb.>8WZSG&cbHZ#_,dMIT43_R>Gf^91#\5g2-c>X<6=gW;
BR#?IdgZ^&CV;+T.?CJcWYaQ2/ZP2T<MZHT.1B9ff_S?/DL8Z[=DE?TEUS7aaAPg
1&B:+\N0&g_Q\cB9\-JZXIb5dZ2-ZEQ4DOPdA/K6cNIYJc0(+babE?D-&.V85dK?
5Ae+BKC2LB=Gd0bI/HXCRf7R10Hc,LULW.@de2e[BG_YX9+a#;3eB0WA>@Wb>+P?
+/X@=;J@:M27<QH4[GVSYgW^&3G1=M:>3K@3fE[WPFD_CN?K;cIZ7/^\FE[VV9C6
&33e128ZGU,eZ6/BKP6OC/P9>M5eF7:W8[Z^\W<f9=;:G6Q5:)CK6?ZQ6ZQFf8X^
FH/BD^&RR1]SBY(WN>CK1V+PTO<a7D_\4abBHc8aMc\:A$
`endprotected

`protected
aKPKc>IB/:#B-1Ac\]DCZD9Zb6f0UOf,_gPZ3?J>I=NWa_]L#5^M.)e:eKZV=f7g
/51)Z9G<8&cZ@S+OTY<.#LNV[E9)X4PPJ]Fa:,Z)DZVP0,9eJ3+C0_AdFWLG?+VN
IZUROT3,YTfV5YX2<Q7[9#JJF32d+B8XYY1>3/1_W<V()bPCFIM4aCH10=4(.J97
,)TKf6G?UJAZYDLXD(45<J,MEG3H7^PL/T9Re1NdCGH(A$
`endprotected
        
//vcs_lic_vip_protect
  `protected
#+Rf]]:)FOPJ=UA,_+VH.+gT0:5Id2]F<EA8=2?Fg1>ad^/8>C6V+(LBMMN0--Q.
LBBCE<L-AVSP#3>#T(T21XaMZgFM2]?-ad;McRa68/eYL>KPQ@:)f57TEY)58+-?
&;H@4=53\_6W801FEB;T>[bZeWQC\@&7BA#G=8M1F\Y25OY(K??2_;6>#6;?#@SC
:/?W0PO]3e[=X[^\D\8_FZ5<Q9c)_f(:<7GE,G,Rc+FC.Te-G)WBcQIY7g<?c-QQ
G4@=8/IG+_6M:^+^[_=1c,+]2XS=8L.:8/^@CQ5BeS@#I>VVC(e?MDgQSN=VGZf>
=00]98fHL.G?^9=S^Zg14RW@X,)fKXUT7.O=<)R94C-QX?@FU)K1>,dc1#de;9J_
8U8LL(;(8Fea,0Zg4=S=,XM1G;dL>P=JTWLAU2-<(;=]&66338LgV/,3?9QdM<<g
B0]L\=5Y[UTQ;](cFCbE8.1Q,.EgB))E@aMUH_WJ-V\N54N]J+5a--CF),J^0>?I
D_#g0@,8]cg@C#X97^7R;(Y:];Ha2:5fK2d1?XLA4[L\I/H@X\GXC#YHFU-J?+d:
2KYZ\YbJV80/aOTJ>.S?Z75VdbSdH58B<D71FeedHBD/##faRW.HIHagfNX:/8.T
We,X-?M9CLW]O_.J71B(Q=8&PJg144BQ5e3#R7-R/5cM,FeBQE.Y?G+L>XT9XSPK
;3^&^b<??CX6fH7U:@[AH#RdW)LJ5D0PC&AOS8:d3M>Hf]^><fU/Nd2CVA(bBc7B
A_6abI:=3?[#fHRF7f:?GO0627Xg-47F4>ZD:7>0b._R58J8693+VPJc=Z(WIc0_
ARc]IXXR;Tc+W&V6(ZePC6=7WA^3KQC@P3E,-&#VIU3Y)<-Q#VAO5H1#AAY.\&GU
?S/ACCB@1&&A3Y9aff4].b16LP[^UFOM@TIPPMa0A:<AH9^d2b(.cNOK3e1D]X[G
#7I3JJ1)9DJYNW/58NC5;VK-bA2Dega6a6eX\Y5a2\@F,N<6H8fF.e?c<Z7I:DTc
9DPA>=\^e^@^NOPG?0S_5Pg,1eSMT=>R<IN?S]=Y;;/H0]+^@aOQ0&,[Vc)Of&T?
,V#:-YO-+e_4S>&&:A](<=,.N31gBb5WeRf1a,4H)+\?O\C[,POLH([XVX1]+B.a
XV4DZDOVWQ&&]R65SGQLSDbX9VAILT)ID&8@M[4Z<(&PO.QWK.d5NAAMGgcE.I:=
.:#]3e:33()^QZ=CH#LM@)()YEc,=e=FTL9@;MV\aCOPWdQHD1)0\<X:Q>[MAA\S
T5?Ae;,79^T0(VgFB,gI;PQAR[R7cY,/HLH8R8_8@K_1@OFN)&?/D,KAX?g-:1J>
1EcdTH]?A#V5>+IY39^@-1<5.&FZG=9DG?WDBJ]GF;#_OfQ][K=.\S/eHW/<3gR3
PQ=X>B_b@cK.BAY33H.9X+G#e&[WcO@C5\7CYe>^F9#F@33M7P^#7f_bAS<?72>[
X:E4_#-:d&KNYKB^Qd4CEaf02I^)>;GeYZI8KU8;)&/]M<-C7UEcXcJdgQ3HQU?c
YIWeQF\ZfV8f]_P9bfK-8eWAXW6Q)O-]]A/?L2,+-.Z6>AU=IG1D/cg2c-,cZS\Q
/+QXK3)Ne8Y(We@_.@4Pc8&C2\(dX>V#JFEN>RNNfY@eU9DP&W&3c^\QO2O2N<>X
8F2;CXae?UKb@(E0B1T-A+](V(64<WFaO^-WcG\X7MX<4EG:S8R9Lf?6W82@.HOU
f^9Q_Zb=;DHD-d<)g7FHFfN(A5)YZ->54A_5[AIA41f9N@4D(fH#9P-LG,;^3/W1
[-T,L_EfdVGZ3V3J=HH&^?APS7T=7b,:,=8=+:YcN7\BV_/<HMP5(FgTR3U>-II:
bNW(75aU[U^6dM9K;<aKKP_\J2;gG6U7^&CLQ:>QR@>^+1PDcfU^S2.1fWBJAAYO
08&+6^AdIAA@X2B3^;2GF5:4)A@(XQ>ME?#OV>)W>S3R_XeB,SZWeK<T\JS.(4;R
63L:Y)JTMD]96c0P&[f;gHEaTAO^[&dUQN[B?9#\ZNL@YU8#4eWY_UUYV[0_R9b5
4C68CJLc<3^[_7R8@]S+a&Y)Y70Z,W4:&:(aH.ZH:ALA(TX:8^4>g]^[)]0.G_P+
JFW^P4NA[e8;I@_<3ZDPN7-[Qe6cK/3@COP-EIO9aBA#9#G;?TK6)W,d[/g;Ie/6
43E.65L;JTIaBHV,QUY18CKE0_T4[5If6NC:^.\M1LPaZ.=)8c+eN4:V>+B7[<ad
.[/[-K>1+2g)MEDZf4RNYZ]<I,L(ad0-HQ8?@ee0ZCd4VOA:SZ#9Q5e]O9ff>@A@
><E>\\ZJ>-J&R^L]&-T(I,?E7DE-VL0Q7?GDH8(-RbU=A,HMaDG?95R2;H&C;@25
@RE9e-ecU.Y3]MTHI_gH4I<)8Wa^7KL+8E)ZR[LPAE+fP(_7=>GKI29R+?\c3(7e
_C5N==LU4d/97X71R0.TUSP9@e.\SL9KNGT>^VV&4U/TGX/E+@;]8RadZb2d]YCT
GA=JC-Uf7a#<4g7-D?EAO\5S-bJ[a.Jd5Me>a1b=\SXM?+A#OSCd-?X(2F\^.?:7
+S#DD0SR9PCJfA6H,L6&>dE_5Z9Cd.)IGa<9McEAB@3eNXE,2Z]@]/EH076\E9Pf
=f;SWZRbXJ6OKa22>JXBN9A6d[0E-S7+HXLZ[(/NXc20daG,-O,cZGM6.YNHf2b@
UD(Xc^^aY1KD>D/]BGgP/:1A2f3Ld.ddHFNcA)Vd4#1d9#Bg&V4[;XRVN-:RZ-&2
fb[U2+I^=FD)T^BG5S@#8D5I:6-SEI?P0><DJCeA&If/eTH@T,gMV?Qe2?VT=F&V
_MK<b+SS1d-fW9D]^SMbBS&]?([T#HbQ0PL/QT3./Q@c1I+8B\XL#FOYO8ZULT+D
[G_Ic3)[]a<Y_dQXRg1e0Ac4(bL.K91SLXHLIY&FD(d1WI<SE:=W6M#JUA2aAVVT
QCKJfgAc56HW;3Z3<Q@UU^d#7e0QIETU_D=SLK+N/I]Lc89-J#_92_IU:;+RWTV>
)3.K(;5.0OgLf\1DGQ&G=P)L9cbaTP3e5=.SG[:=>d:<:f3+M#+1.S[1LG>)\?a>
[:b\Q)FB2/TU+Y:/+1Ea@]4X[XHF.K/H.2\K[OW-FSfZcOXDUD#LaKGfQW_&C<SZ
L1-e;JdD^a+,<#-dWZWU\d^+-6YF#a@:9K)f[=aaNaF\Z@ea^F/N)0a]>c?Rb>AY
.J:W^T+&H,]4U9>/QAG<K,f8GV#6?CVCT>7+6(A_>/Z_4a8Z;?,dR_4RObRJRdFT
3(3b2LDb8#->G+@W;5OR78,FGKc>@MO.bE3==XPM<SL@/1K.gf&78X1:_QRB#_X_
eO?R^G624^XXJ_)XM@GQ_8:5>N@\--6OL1:AE)dODg=g81NZ(Z5Hc[H5;(ac;HNI
dC<dJefXXPS^a8WTJ#c^cdf:W&\O+,AYG>#4VF.4+\@NI>Ve+S.=fgCb-RB9?;cP
XNS<@)W[/L0IRc?MBa\.GWQ3<^g6-P?B=DE1+Ie7,QW9^D;>8L_6+W-EY0;61]NI
/?&PU[WG96.#48I?&a+[\1E<b_/MdX3ZC>W3-b4K)\X^2^V.QS9^OH)U:SF(KB;@
DS/HCE-E]<P(W-R]\Vf)L^LRI13_4\_P/NLS_cLX9R07=e>B3-O@Z9:4-ONM10:F
=ML#>=RF7_>cITMVJc#FK>)<;a>3feJWYV+HNbZJH:D-gdR;YW5H_\F;0MeTC3>T
8T&C\JYI1OTaS[V]O5-7UFa#U&LMF?2P8bZX:245E^8OM<L5aZM<5Lf)M1=]KF6Z
[C:\+.P5E+S)PZVFaeV3FfY=Y6\P=G1A#).AEM_]X-_VUFQ)D[M+QH9W^B>=081E
TgC=IT?;0b5I8EQ_F7-55HUG[a.Yf)>0dA^+,_dcE:\2bCKa1T;:/T9G[M1.Q4F+
0L#[Y]-D/bW=ME[,A665JeD^aE__S]#V,g,8^51U.dfIDULHc1]+K-[L>U]96-(d
Gf>5RA/RKP\1GeH\f-87]TT_);4c#27.Y/-S2D^A-,6;474<V(5JCXT5g+MSJdB,
HXPUL_)/P+5(gQQd>B4PY6Y@5/U2ZDMb>4:5F_9L4R.16XKMH(]OIdP^J/<\,Xd:
#2MDZ)+F/AeOa^UG,_aJM?beU;9QDHBZRG#0==R+7-77)W]:.VEb_EcN20V([@eD
[g9+4UG/>X.AKfW)NJ^B?Q@N#+L+1RcD7-PQ.OF(d\;R=9,DWYOVX3/@MGPb5ADM
-\H2U_Z#R9D((0F4UAVFdfLKH+.(WFH).WS6N56Bec6;8Rc;F\gLUb;/HB.XQ9Ta
gfX.XUX,HHY<BJF..#?&REbgCD8bg=(ZH\<5NPbO>38^OQKDV>PJPdOd9IT]KTg@
#XQDL[ZVO5eaH[6RBY)e&ReMPg,V4X@=N+0HA#Q(H/e8TJ-99V@5WCf].)#b5]_(
SJD)T=7IY2T/G)]@NME[V+?REK-.FQEFH&0SK<W:Raef2^_IM.-7NT8XfT>7+G/L
+0G-#,UAB]R/JM8G>/(b@C5LX&Q\DLYBB_P;6b9da=L/g34V+,g^P&Z#42V/VX2+
R.4UD,B@AZ-A1eF#]W)9]g2+4VJFL<^c,B._;>-c1C>c@BgcQ8[Z7g8CR-gM87]D
7-X]ee#g1S]B(.2J-E^KOc7KBO+VQg,Q.PBP,fW]&a,b3/a6H/4E^ISHR.+4+bH7
[cU^a7d/2dU[T9Y@&5E?fISI,Ic-]TS@M53D,Nd\f0\QN([8e<V0I)R8FI.K/:O?
^T:dQ-6+6)fL-2QT26+@5PHZ0?8PdFT<g@S&^@V)5QdU_f@<&Jb/\-0.WB9REB1#
bWG5)\D+,3EWWU1dH#+S3^GM]/=L4e+dAX+?ON&&7WQc.9BIcV]g#8#Ve&1XC/VP
-.H;--a^L3:DA9KBW>8UR9P2Y#DE3e5.@G>FccC6@>X@#(ec+,^Qd(&G1MXEe@G.
GQ1Z_=W^^dFMY2,;C^ASA+F?OK:7D9#G1<ECPGFN;:P35f^+>X[,#MHT^D1.SUS<
YC7&(1R9TJHU\<eCL063>SJ:E4O\RbN+?EM2U(+fWb0H5V0A>AWCe3_dg)6DB[da
ABHgA(8>RG5d678CJAK>U;JHGCI:2&LA2/D)^8CDbO;@=,f20><Y#Ub69RSS/YHZ
N>=VVKEGB\+Y3eAO0FTKR(E<f\6_Z7Z6Bd1]/2dS>0FJ06E(,eeZdU#=^311?a,E
JRaH,B^8?LeNb4C@W&P+A?BG,NXYLC1Y:E]NJ7XVdDPFec@eY)eBT-3N\6gJ7C6X
EBVF(&,#I5&#fWTAFG5a\+I6(O/XXVFIb)C]JDVEC4I\\70aM#I/O,_W2B,-S=,+
]/\^.0\II3A,?Md=eMf]E^[B74.bU60\Y]?Z2Hg6_aNS;Z8Z^@O#6;CWH3;>BRP[
e_R<R?8[#XW93S7WQOB&8/Kea=^K&eYDC<VFD=@\(QcPB<4)bAIR2D#[-IKL?_2:
[QXP\0[3W23,bOF/,#WAWO>C(?]gBcC][E443.NG5(5J>KQ1P^84MJ+L0=Jb5c?^
L6(f&\K/+@5f(b.X]+BU#9QBIc^C_PLA>RS+P>9.4T3JI;-S[A8&CWS>7SYc-Eg@
N&?ZG=S:3EZQ0\&c161;R,I^#58#1Y=I9cf,_8e5A(XIQI<;:??]aKW4d2[=YIf9
IZZgS1\Z@N2IK7ES&D;X(BF>UGW@O0<8P<N:3OV.-BeaPa18)0-\]\VL@G[K6JAc
P_0>G6QFASeMK#9?;6\5CK:3/2d+2CX5\;d]/IX]LQ#R>2V6QD86K56KUGbMJ]2P
@ZIRd_\a4]1.<C<IVWf8#HT7LTGQ,^eGHI4&LZ1d_DMcUc\8PLcJ,O5+TC@\XQSD
7;=P(2VAN=C3aa=DO83PMcAKSG+&V?8\Lc44&RNQJ1/-2)P1SFf_:QZgbDP1TA/+
TL,K;Q-QBXaZS2_fM72U\f&QCX8AeF3IJ@+^P)e:_HA38c_[Z^5/e?OE<.=B@]V/
Z8<O0@_N9E<SNP&^,K56IgV94SAOPa@9ORd8Ae51=L=_7b\SZDTN.A-204KcREF_
R4=f_c)6#;FWg;6)B,CT.U8S)K<4P,?2[#0^)-#CTDP=fZ4f:T_Rbg\L?&2,Q)Ab
Ag3065[E=+S9A(I<SKFN3_25@70&[FT1[+8ZK1T&<J+gWS9PQLW7Q]1LF5fR1#bb
[/c;c(a41KT-F#cZ)\;K)]Q:=dKMV3d(M3eG?MeX=?2CB7W/AHe(MTEcQG?RIODE
NcGLJ:RdIMF&;G@ID6HX9COa)#.eFF>T60_;F84L:HX&U13N,-^G4R@CA4;V1KIJ
U@LaJ4EbQJUY@e/++NZ]#)aX/,[8W,KL[eAXE:XYFRC&E$
`endprotected

`protected
&E_e93.eL5eJ?eS_CC[eZ=#aO<_X4>@=EWeb)_+K9dD_JV&@IE(G.)WQOV2D(SH<
@M3._GE?<V2J/$
`endprotected
  
  
//vcs_lic_vip_protect
  `protected
]&K(XJ:;S#FG=KVId-R<JIa?^)71I(._KQ[)M.FHTAVU\<=9./W>6(I)[,NRd?/K
Y2E27:)6e3-NYVbRV9-VP_LN+_6,.2<70Tc]@,TW8TZ2Zb_;9Ga(J]V/\a#^^cg;
M;</L=UDHBgS>=eb7M;S\I[[9\VQ8/\7)cL#/SIWI>+P4Z,^2CJfNb_K#Y7)/\F(
XZ@M1;)/<aM.f[_S&=JdB9Lb;I=eVNgUCTX7f0SP#0d4ZTUNVNCcF<?^R[^6e+K@
CA57)aC#Yg#)D:+^TB<RV7I]ZYQH<0Y0]/bRfI@SUe/O96^^1(JdG+.;]8eD6W,a
)^d4_PAA[ZH?bJ_-E(;>(J@5Fd34gG]WHJP+IMN[0]OV5De7TB/Y^@g_<EAgS\P_
Q8Icbf24G/VcED?L,O=e@)7]:R59A8FUTM3BE+H-XQFN<88Sf]+d30A;7^gC^C4;
\DF?P_,+VYgaD57E5SA([GRf2O.1fSV-(VgdIf0JLX)HO6-0bbK[4[K=c/A_K@/(
XfZ6GdHJJF;1D=0:.b[5A0X\b>@]1NXEC=X3R@,NT_5SL66;64::KU>@I&<bOR?-
^4-PfSg(DQfQ]QV-1T_X_fM@=T-:C0V;4A8+70=?PE6XG@M#c_cdW-Fa6AA9FL-V
2/QN,][_FGZT:@LCe_[7/dX^K+.+YaScMWBX[DD)8VAG.90:.]),&4+?fNK.2bK2
(YQ>/:);Q]<9TcGeZ;F&7d-/QTH:_IC02)VN7-/Ye2=3?B^ISd54FdIG.TN?O8Pe
_eH0B(5fA6DU1QVf.3+N2=dIV@9a8K(+WYg=HE,OML\^GRZ^QGAV@BBAU>-7><U8
.WRA,S)D@0FPe\6EgVKHW.>,@;R1Z+eL^0+,:.KXI2]VW..#?_/+^XFAA9=9Md=G
1)\K,+<c>17CVA),)e]+7g?M1aN0X7bRP>A-g;_W+G=PSK1_IHdbBRQ4DRT((5GM
]XL/gcB#7V5&7Fbf>FT,BadF=5ag:4R]9@&:J5.e7/ZID@4O>>g9U_Xc\.&e&C&.
2.6;VVYN,A,GbcZ19KU:U/4LHCa?WFa,U&(Ng3VAQ]9X9CNG3TD8&aLF>;L#</Yb
>R:EgTXOCWfK/A/P=8Q>Df:4OGUY8ZOV4K35MH3S>J6ZB&GEE02^gQJ.6=;5,ebN
9^#aKH3:M^WSYZ856N9U3.Eg_,GZGDKQW?VRBOUZ-1<^N;[>;HATSP308JfF)@Bf
)d)-PSCXbPEHaF(49X^7O(KK(GA1OL)(UB8QLBSG:HR@9-f&df3C[K2Ue/XbPZf6
@e]P=32Y0D4eg?=Va0gGX(&_MXQ@g:(4UPR<]+MAWPSHLZ+?7fW7SY=K>J3C>F^#
V,>1)RcDP.=eE8e@LSF5e#/\<O<+K450L/83I&,14K++..C(<68+aE9R:#J7G=X0
[IgQ.b\PJAOUMZa@VR#JM99ZN^03ENGYV86B_#JaCEOW=?Y+N8C-f-e^fJ7,a>1#
>;MIf^f)ATTe;Q]43aFR>X)>:QWM)]A-;]FUB(VM89O1Ig3L)I8[85V_:2ZUf_ZX
^+b=)5&J;>Y9e00X)FO8N,g53P+]2ON]^-;IR=)ULQT_[,eI3LTQg;@6.(F@5g>>
-(:XSN1B5-;4]ABCL.d[6XB9)M43M@,J<J,c^GgBFe#-N\^R#7QYKaN39PO_UO,H
.+U0TO0);Ne3^0PbJ#TQUg/\:<d:E3.a-\GU:Y[2HFVX+AaZ-^XHFAA&;E2)RX8V
1N5SPg^O(d0UQ7WR2@+:bY\UQCfJPPX=K9Q/01>39MR38X_cfJM9_Ua)2XJN&dAK
);5FPFKQWP@f0QXTG1T7=(2\>gaEZ_X/Ig]-BgAP+f6PWbC6[Z:W6EODeDFMBH:\
KFdWZ\a_3]=T+9b<\[(J1[Y&MdS&.J5+3K#\0K;:LSb.:6]5Gb(5V84cLT:7^/TF
?gAXZV&0MB0QS:NY?2&GNSXZ];+QK84SFVT&Y\_cJ;6Aa32/2E.^]EM<FJ(RMG/F
42P,G2Y2(aT9KN5TX-c6-\&5<5.HfNU+IeF4AZ#,XC_CK_fCL;X?eSL)0aKd/gGU
_]MOA6]GV<^]C8-V=?N1ABXRTUU0TYWM,EXXCHV3V5fLE18@<7CE:Nf^A.dXSg\:
CVOG5:?eX[>_P#PBK)Y4O1I0Je&VXd\V7Jg@]D7P8/cgLeL.C6+Ma1)VU?/I(NZ?
O--Z2[?<COQD^T>e6P#&EI#T7Ca2CbY^+4\b(d0P/HG1:e?_;@>=XBT-S8852^-B
6SQc@VA6?OE3@H.3S8YQ07V81BYY<>#7&gU?FP>[7>_I7EN&4NM15@b\Oce_EHY;
1OT3_B3L0Og;K^g-VOf+OG\FBe5GSJIeC83<;N-#3P08g2[/B);S]ZGKME])#T,<
(MUJ,ZaUC3.]SH,7[g:I5]L^9>#N7TgR/5K]g3A7c@I<b,IXYX3C#SH,1f\>PXDM
R&&(<>M4e1D3JNaZ@#Z8a/(4PWc3^;OA?be&282Z-E&Y-,[O&\HM:<;86VA3X>=\
+Fa[@R^;P4E,YJ]:+ea/@8+1/Q-[8g5:L&UHQcX^e#],+KYQB+3AX]Q+GWee\:^Y
2]X3LLeB_IM=SY,\5PYgW>Yg8LKYb/M1H95UQP0JL95e\ZK<:dY5OZgTYD/5HP,=
1J;F-cIA2_F@)1QP6X-O&^@;XG:P<-K4e/)J2Q),H9J5A9eS(W>;aK63d89#)..8
ddQ8[LW@:45CK),?>4G^?#Q(N.>3[9/.+8]P^6aN;_;?NQ-8fCSEC5B.]f<P<;8[
UZ.:42f<5S^K\SNIZe]8\FD4)OC<3F)^/PA(._726=66G\dU2BAf#DGC<e--OVV]
G#b/WfT)B3LZc9QbYJg.#5ZA7=0P-VSfQ<4f079Y\)Ba^&0_76;I.)2E7=e:HXHg
[^C:<de=XV?Z?/@#-XN93PHgcc/Z8H)(>Nb=53,I4aB7\XDJd),,;_Q1-5=.&OCK
bP86&_MT@d?\@2dEFC2[8>HR.2#87MZTX3K]0f4,d)Pa?fIKNEeaYG?E[a,2M67\
N-\4G=ec8^cSXb6\E-\^f(=ae<KR32R]3YOS5Q2&6YDG-4VNe:b,F2CA00/(?@bO
I-gP\,[ZC_]4>Gc8BCIE.;5M4^+N99Zg1,=-d5g,QC3GeZX9RZ?M+OV:)DW6N)2P
,NL5CZeCbQOCe:4QIEJI>HN<+&@c(e:Xb7ff,GCD]HFWe6^TQRM&f+G;H\cER\6Q
;g^&Se\:dM<O_7JJcFBMJF(c>CUBCJ_fNC41C0I5<RY)4.G02(>B4JML62UZe?6U
=JUSg#:EN&/P:)&E6RbUN4BYbWL\TJ#d942B_C1>IPI[]NI73SfJTD?LQ/E366:]
9Z&L_-F-)RRGX^Y]ZFdY74Y+C<.TB[U,E?60=;(2TP99&DJ)QUA+PE3_^B701ED-
GcUWRPPE3AK(4I9YLKM69FS,W#QWN@)@#9[eKAd7eZNd&/W<ObX]aQ/BFMa7Q(MK
J];C93][0ab.a[<WTHPfbLWW^319NY[-NK:UU?Va&WdQN>SUL&7BgV6.&-;@(EE9
G:L]PUg5Pc5B0BS,ecE\bM(-&Gg/@gZU:/(cdb7-ZAEJJTNaOLT(fY8S1=ICH:5B
c)MP[ES6G:WXe(:O&^J2JU&fCe+&8+c(f>a-)5^3#)2&0E9K0&I6.a0Q2-/5M9MR
(K_D/+]HcgU-O[H>K#_2NMVFAf1g<KZ71EaLCf[UddRaL8X2.#5GHGGFJ&@PT085
f]O:<-+T,DBL?eSM;(U5WW7fgH4.2)2Ce:.U#LR^#E9J0fb<RBfRT><Y&1/<XKc4
5Q(35/CMf<CNcLT2&[cV1,R,G:?Q,EWC)gd)=1DH4@AME))<:VVH00,bLEMIOJQ]
d9D_O)5f\eCRKR;FHTS\.:?8@@2>K8JYfV5f)WeYM.FdEXW2ASedC(F5d5^K(72A
LgI]b;?/MHcIY<_>3RMUP>DO[XWA?A55WDVR>MS[Yf.NU#EaLWR5<U8?9aOZD-,N
9dYW>_2C[F.:(;]G0ff_cbf/gC<Q=YMS_,VW1ACV\97IJ5H&bEW8_1-Z4IGFTOW>
9FKKf6:Kb<gA.]ZC3b)bP[JZ8:_;gL/>U5bRS]d).7D(@/HVO7V,Kb8VX2EQ3U=F
7Z\Q77Pd^1DMZDTL^3?dRF0SJ,3K?agcTCI8DL?I^YXQQHM0QbLDJP:1D^eDY>MI
Gg_c?e8X^_8RJU(=c+9Ib0PF1e;g_:T??HU/_dLR/6+4:-E2g4I@ID;1XJ>]A9SW
ZgU<UZ:0_-49MXUKJ)]QR^df(f^KQI)+M6JX@=g@R(KV_T6>bYfRf^K6[fMV5\A;
-O8CZM-cJ/[W:0UXJ4E-&STeE?)_6@>9O#M?3Q^##g6/TK^:-VRE^VOFdHSMgA_0
5(MX/S_,X=b6WVF<#[;fCLKg?d?)9.:X;O]O&#fX-H+K_]7@Wg(g+2gBH=Cd+W\T
[4/=FVSEK)Rb0X@EJ&>/<X#YbFICIC\&.eQJQg+Gg5(HEL:+@fb(bBKA8M88AZO7
WS\R7NW0R;<1O4-F4Tag7VSZZ@63]@+JO,NLE2DH)++@?7LaDO\XeAQC1\6W,a^V
Qc:M0D5M3.WR8T[OeZ&PO3-bf9]NP\3/UW@6g9X8A(OV8c/SG1DOTA[GU1T4M0aM
))3[03Y+;?Yf&/)M@O9E]#0E#X/?E:OM21Y7,d(V7I+)PFR>E1?V@YZ_B63[;JU-
J/Wfd,gB[d0b407\3JbWZ4S-]H/7WM2>X/7e?<@,f408IKgQ4(Ug9E42<.<BYe<F
.\QD-IZ6SMV_I-V8X&CGWF/./#WdGJNMg[SL1FP,aQcHA#:?YF<I0:.M\,U6_+U@
Q.Se_U<6+:X0+[X,2R;H5Dd25M6LRV<ef6RJA>baXbF5FHN]Ic(/NKb/H1&dC0<Z
N8PO(=@CR.N+.=I9A1C<NMe(RTegM,W7O23#DK.0;8^,QS4ecU)MN@=HI>B8;0=_
be4BM2M6_FO]>-KANRa,>a@-TA#/.5H)7URDX/[F)g4),I7Q9)2-HKf/8cDCcACS
E6X^AXCO+TA_B&TNB;MH@?dUcdV<J[7#eH+L&MbdVMd:]GA/L.K7(d-/ZOaI+)4N
8:;Bf&V0=KOe/:a<M]Yec[?KL<(UB[:QNGH0UTe1J\^#&3a8^XK@C=X-&590XFR.
65]>^[#b<GM>4;\<30eZO0g29FIN-JJHPdG?R6&eUB<CU@C9;Pd,:+DgG(^G:a?O
/XB:/8CN-DEG)20>-cCX3BS<\YY_Y1S#P5(L<Q7YE]4^,H6aD+1G/&8+<?MbRWZB
@I7X1[J6:+H;\X:@\Y]E-0P_JKX)9RSE,XVBLSZ]8#53]M8Q5D7_=-J]QG^&F_]E
CCY;;gS4UA[QTSBIXN(V;5E?MY#MU@Fb6G6\6?A4/>(BPH0.MAV>_]QW7XC;:&0I
CX,.EPb;Tge<VJYZJ.OSWbZd(/UK?aN>9(G8@)^;?Bag[D\>]73?=#?H07[0_3G,
+->5bTcV3.P,I57Odb[Ka#2]0275[OLAbE/BeM?,Cb?U4&=Z\Z=1(4&MQB85H=.g
&J4P]YMbH>8HE?d,.Z^&SC6#Z,U9-#UQgI@dTVeg<Ga.PF@)VgC/C#K6eE(E8IG(
&gUEN>F1Nb+?^Z^QEacCc;HPDSf>FfGBE.cD/)4_V[7dN7I01Ae]7M7@.GDX^<:P
LJJ>4#d^.?F#g1G5^&#cX_^R<1gCa>C]KV33OA:84^He,MY;^Z+S7Vb\\@\:YQb&
BG;d,?J.(:D]bP7SQINb@E<1c]37+5:Ua&J03TVc+QOR[5?3KHF0_Z\Z9Q?-XKH@
bZ6GMF4#;>)W+KXZ3A56^HWg]S1HPK>[_1L+FK+[JJ0RaP);a;VEX8,[]91QY+&^
=FbZL.O8I^8GEO^+MdbDa\B6]3&Z^>5aeD,7GB?NC#+T_-A]Sg;QZJ98XV8R/0/T
S7UXdd/_>U<S@YP,Sb\4N^b4fa]XU]/Mf[(;/DC57WP+,DF3.cJ\?e2E^/CHPS[Q
IZ;-((KV^-B:,D7^.F]+e-O8HCUOBf@KQ)R+M64JJ7I8-OZgWbJb#IO]9:Re]QX/
WVE])YWEM\[]]dO)+;=6EFK=F:)ZS4)>[-ID>,(^XH+5D>^(\W#b@b?MbO]4=[87
_-<W<=YFE.M>/G:M=O?E9G+K=D=CcC.Ia15MS5Bf_QQeI<4:Rd+PV>/-:#T_IaAM
/_T71K0S.E6SZ9d7R9:fe6fdI\b;<G+d?K]0c.TZUdH)@8O[1MM/7/24HBI;=4&4
O.^Kd9H<(a#6GB7R)1Mf+PG<bK6^30Q8UE.+)-g@6@/WYD(R7.QdJ1U>0@60c\,;
ed+WS;5aXMLa)4X2\YH4gH06&R.DG-G\Jb5f:-=J>/W_L)@B6@HH?YM<>OY<W<;M
cWF575YR>U9HN]1L_B.9AECDA>P:_e3>R4Oe1;5.VMX5^2I(:gXDP96--=WV7LC7
MNV^_E=O^0.D>Vd;=HW<3KQU34^<[#^2a]ZD9dJ4>Ka[/GeDQ@[JgF?4d=5R-CJ/
<Y<Zfb-2b(3LaX@7YW<Lg&cQV<P-YA&HE.D1>f3+95;X:&C;Y6H<6QbOI>1]<;eH
O#N-+:0ESK=d@+5RGbX+3>CE=,J9dc/RFC:@E0S9E\&1.]V>GQZ<7WAP_)>]/Ra?
YD+N=Wg:V(:1KJ+1aO99;AP\0+gC1:2[<DHcOcReB1(M5K:8-9KFD2>/@:Dd(0?X
O+()1,>ANbWGO8W-^)gb(X3_eU\=@L3];&3U#1U=8G=Y1OXe20HBJH)e=]_3X9?V
]dH)G.>Cc(O2>@c)>11TXIW\]L:^Q<WOg#GB)SgH34X_4::g=N?GSH@F37LM=M15
]&[(2#S[NBQZb\g\A[d9_b?/+]1AXKBYb@K/VYF7b31aW>5\ZKA+H4c)QGNDL96W
<Ac(NQR4DZE^0D?b:OZEP)><SJCKb+8bEa@D=WQJ;]3Te5c+Ig]V6)OYc<E-cJMN
(K/&MIO\J^W)-+(JOEcS.7L<#(9\S(cNdVOY/<2D[UggAR4g\1&[CbXg_6a7LK9P
]<,REcc2,:gd[Vd\g/4[H(G0b^S@8_WZV7WBIF-,)_#G;BcTYBg2\MZaOOZ#CUT3
e;-FSY>HaP_4<5aNEeJ<IV>D7&aa[^[O?:f^CaQ0E\ZV\WDR/N2N[U7TB51C8CIA
@OV<Q82aBOBd>TI,11gI5/ZAO12R&[Y7^L5^I7E<8U4d\b?E<Q8G5R-K6)d/9E<^
(HcdMJX8C59VW1UA1T-CZ[=^L4Q4ND:>C@IZ8=4A@8D\,Kaea/FL.36F)g/Eg9HW
H):g>H4XW++[DMZNE5UHX(C8PaWY<)1UX+H4BKYG:KW#,6C]F)YMT.JJ];YP.MT4
G)D@908CUb_K1>:)X-d(ZDbf2XXB/HQP_0),?55G68EM8X?NKO]N+3^e-)#FEA3+
BJ76O<#K6MSR.c(]]W<c;dA(=9_U23[J12DCI??AGKWBdf5O[)NdGJ4MLZ1Y5H/J
RLb4\,7RL;IOa\_VZEH5S:^KQ>329@QM16BABcSY3D@OFgQ6c:I(fRKQ63gF>TO6
7)0L;1APWaRdHZNaG5>D\E349L\S4gVCd9V?+E(@-L-SDU0L:Y0T+CJR,PSFAA+\
Ff?<#<DCX7CLS,<M=)9J#MG)Y69M\AI-3]2;<^GZJ)&+@JaEAP#AV3RWG&XF4JPb
0#S/EYRX5cE5+TN,D(QV=YLB@;@a/SAT44/W5ebT)7[L]cYX4+8/=-<CC&9([fFD
L.JdH/DVK5KU9YYK>77QCJQD6/2L&8d@P>K>WJ58?beV;^STLYY7OdN9NBUKBWL0
HFN,g&131-bbRIg5+dXfJ:7QdAE2P6C:E=)dX8CB70\,9EZR5LLXK-8-[3RLgP0d
1)C^0f_:E^UE5&?A/78,6DCDZH]MU>a[4V-6^M=HWHB+bd#7F<1>G&1.7=B26TQ[
01SP-faI-[;Oef7;F6fJDXSZKK[>?-+&.9>XR^;gF_RUO3BcA:d@YNaAHE<(JI?a
-D0_HD#2a#P[DG.E:9dR//.(3Z8b9d)G_7<[?]Sa)+,B9](1JcO)YVLGYBEWXDL?
c2VaEE:=V_3WAD[U=6^VZ9X\RZ@3)g,K\C]:Z#D)NJ=L5IX:A7NVFF7C/97\+MdY
DK#gVf9A,U.HLa<YdSLgEbJ:M?F8UD4E<FVO45A5MaT;U,@Q3AN/Ff70(9,ZO:.>
Z3F^ESb87\S3[f]FK-<L(9/OfLI>gJ5b-)U4TJ1.RG3&CbZa@W9)EH@#Wa@IAK)?
/_Eb.)Ub)5F3<[=af1K#VZ9aJ\K8VOG+FUH<)([=5B@YXW^Rg_ILaK#..f=S)1@8
9\H&1VH2ISPRc62/#f\Oc4BHK0Y)R_Y7dXYC/\+>0dOI2e/b=(5L9Dg5#eR:<Hgd
F0)Bc-S4c+VfQa)NWABJB6D)PgAFO-;(NTd54fXg/4^)R-FeCf3WV_VdWY)L#KM8
c;MFbABKGgT/G>]Y^9/R\WYT=9(eE,-AVFTU8-VdaR.B>[36Q8gedMET/e_;IIW_
.JCe4OG:XBX9@aTC6H+@BIce6,g//e)ZJ;2cB(bCf1e.JD(UX0WeAM(fUE(e#E+?
YU(_HUEg4WA+T10cB_=2b+?.)_F]^1)e,Qe>ePN09B5,Kd+043W5=P@,,A=[BRI@
7P72EL1;6d8J>4(=:GOO7ZB1AK?-F;91O;gdI_I@Wd?d#R\8-ABWNB\O?\2UQGU9
#bL.(N+#N4b[[TA<IQGgbM/&>WOT_,BO,>c2fFKg=g#-B+dU+G<,d<6BTEER]=2Z
/?)Y.2O(ZFPc>I92b=ZBUL?OaP;Y+.GZ4)K2BM6(Z?C8F[dYO+Z4:gN#CN.IBF;f
-)NSCb=IUY2a#2#A[G;J>SI]8WH><J]J4F?T^T91gae_0DNC@:X;RR&8O>Y<]agM
edD=@UFf+049&eR?302POYQ85\6U6Zd?3eca[:LZZ<0VC7RIVD@KCQ7UJYLYC-YX
[;8#-K8GP?0^Q;2[ZN^RWgf-UA-c1cg(L)ZINQ4[WJM0RV]DW<PC8MGRN[6>GXR,
[/UBPLHM^;(&1VUR-XeI?CXCbP)_O;Ue50\gaHH=WJS_R9E<=?gd#>=1L/ABe2.N
g28cc<+(@=JaI/I[TX;70F(EZ4c5[<RQbX_-cK>d9ZL>dF&&8L:Zd1X?La=>ZPPF
;>:<X3<XSS=-06F=+^6RRg<NR2+/(g0X9,.UJ1E0/4V;B5#_fg6>[<W]MLN;g0TT
4ZPF:YI-RSFac:=0C8<-:?a5,UJY,2]ZHVAN9E>[;?B#bRU;:T/D^8c/J4BDMVZZ
Wf)gT5LJ7gH.Q2cI8.;=XgdWUe99.96RK>-.9Ug;\)CS[PTVSZa4baV9.W7I2ZS[
,UI<4P-5e364\&^e+=T+ANOE06)376a[;Jg7&?;>GRUWIX-^a&Nc1)=?_B].=EBW
Z9=Y08V\cZeTA=bfRfEdV?Id^#W,0XDBA\JA\-YU[0^8bW5DQ9+dIKZ5[TN3&G@G
XI2/DP,g_(<+5eNc,\;G:-H;^V^KIa&ed[)XY&5AcUE9SXTC&+F:J14P0FPd__g_
E=Y()0/[(_e0I5[K8-RCX^;,J=U\\/9b07[BE5B#[(M_U3<PK=E+dJPYLO2Jb3A8
>3UZ3HIX<-<+PWBV?>19025<K_L&8RF&d-KMP=d>bZ:.&AdT;4LAAW(^S(TW?=K=
3(VM]8ObA5]<-Z0bbe,g]d^1L79/(T&3>>2_CGLb=4Z^/.\R,F1J+<gL7JXQYML&
7dIcJ&[ffZBMR-FdA;a]9[f#CdeT#fH#\\CN<D@1GKL]F:=0:c,6d;,TV(D+#K[]
&GR2W\-DW=GN@FV<4,a,;V>]DO#WWT.a1<S5X=02EfUae]>(_6&_8NBPV.H@YFM7
QZQLc/[[&LWf8=8:+M482H<;HOc)3f.YZ96J[-.U];=DR?D)5@Uf4<d_DD[.RE-b
C>=bFP&-Ne-IWFZ74LJXc)1]G)/T-99(A6d]0G+-JSW?)cUS5_<:9I-fRK+V_;8L
2/LdWY5-W<PYV+gKf(gTQ0cJJaa7bZ3dB@CM?IL9)(JNFM^Uae#UB)PAfS8N9-8#
&D,e\P0Z&JBXSYK>F31W7B:T?40^W-W3&3\]__KCI@b@7QI^CTV@>MG#S3ITFM;?
N5LJ-aOQVeBgUCgeW5R0g5g_Z=:>25-^/UU=,gBATXHWd,(PJ(Q@T0>-Ld)cb@71
fYC=S4Lg/KG=-03T[DO;5d;=f7<9RHeMJ135:PEKPg1C7c\#=2B,V@NdNH+BCg9M
,5-:d.#5,e/e+/7+f_9a)1M[:1[fY9Vde^5JE)A5\3-;10d4][UWSCJO\:R]>2@#
H?446RL,[6.>K_BL=:Z:/Me3e^=Z4WR<\[240bEgTEZ0M,(Nc7:(7H)M(OD(I2bX
HEX]ODaBCadd)UCVXYS9RZQTKE38OJVH>/2YafLKX4K2&RSe@gCXJ)/2,3fZ&P@T
W,JE&5)X#76=3LF6I,]a-\]=<@f0AYRXd;DB]d^;e9SJ3=SFQ@7&IG;^];2LBfVT
AWbbMZ1M4g125g6b<5a?eJM,,I-&LL+fb>>-9^WDcGe]:.MUA;MUg2,S?KJKC-I4
H=?0#U[(69WT?]V5-X76:SD:-BcC3#7I?QX9=AD-KeCc-JNIM0S1SLH6(I;dW#XW
CD?C7T,.R/SGOZB=&<NRYD,;L9=;U7e9e2/-5cNIVFfJ#c]MX=/Q3Y71>FQF7<X?
<Y,9c#^.0J1\0B5M;PeKcQH0G9>AcQ,E[FZ:g-3[)K8e:6L3Ac<#9c(CeDPA4\P6
V_Oa:IdQ(^BJRD/KXa[EEMA;Nd:DW9W30O:@&>e&BQ,O+@1^KX)=3Y?+&/^\J?Q[
Jb4?SCOZ+?W#)TXMSaINgS@589DX<:4c&V(#23U7&F#S1KW4=a15KY=Fb8QMf@f1
Ga?=bI/f&gHa95H]H@HI0&BOY(L5ge[g6F9g?8-cS5(E(;;G^(QId-?@L]W6YRY8
7WGaHfXD6-Y<E\6X/:RUKU-RP_UFQ__Ig_?\A[Y:HXbII;#R3AIEC6\52YRL+gg,
6GU2a2PKTW4?=gPKJb#EOeJ&OZ+aK<COP?VMGBOSS(ga33Hg#8L65,BBVX/D?^8=
-A:,X[4SUMXHT&5@.B?^5CX-CS_SSV+-.SRE,d2Ka._-Y=cS><_;b2L-3c\6<-FV
[=&Y8SNDH9.PSL3aY9-765cAbB)S[@5H(/@Z?=^V]\9Y.e[BaCf-M=8:H6=4K?+U
.W-L6#>c[QM_Xe.;Gf,@[Y)OEaTC@D;&(S[4BM<;LUX0IOGXQe4UbMeMBg-S7J_:
T&7//([I)&#^Oae;?>XF<+#3V&Ad@^L#5.K[f)N6eP7cFE2d&;=S/U8V==KBKa]@
5O5]A?>3AbGVd6IR[LWd:+ZICXg<]>5Ce:O852@K=[K3IgHHF0EQDX9Nb(>[+1D+
H=.a8A#cSReTB4\c:GJQ9Sfg=I&V0:RD,2gHg91[gZVZ,aAMO4](./O361&NP(gZ
aHMg]H_ORQ/<B__[W(cKG#[FBdB,@_\</50I;=CFE&53)D)gf>-W]\_:9<P#2MaS
T03fZT[HYXAE=,=:a01=_ae36U<A&534/=RFIV8+V)-7S-6X-SE8@E.[e^&g:gP2
.Aa78U<_L5YcY/B5Q5:?g7TRgc3W(ENPQB&e-RUDY:V8&#I^Ja(2D\bRGg-D/Y^S
(WAG/N8.-XX<II<(aR@cXY5IW7+WYXPIeQdDfT[S/8;38SUW5PWD3]@C_\(,a@3<
#C75>?.6(YSV<fg,+];3C<KXB#,WVP3KZ#BTN2PE7e<N_S_D)T[NbE=PFSKd(:1M
O.JcO^NJ5FMZ4MK[e-Y+6f->RAYM/Uec8QB[BNEV7YJDN7[SgLOE^>XC135\NWAb
f)LDbT?)KW71#N]N7.e-e57/<e@0SR)AL9>1X2=7AfTO\(HW=;.03(c6[2DRB3[<
S/1eSO[a?D=^NT>VB&]LcG^(0ZRJeNbg-A6fSHgJ5e/],#bc];g0)R,c5QC9<@4+
-eP\dDABHM-I\NGGO1HE4IS)d[5J?ccN20#W3&A2:7WG:)#>+A\F(1.gX/(XY1BH
J73^AI5c)V(,KWQCQZEeCF8Ie<WF#^#Q\9LJ8fQQUI#Q>UI3W8S7(Bag@E2Tg#3Q
2aS?S?L8_]I,Y)8[O[66--61bfbBN8:g0c+GYOV]B-b2B_C;483L;,7&#0JK@YCB
VM4<fb@_K\TeE1C@gd>Q^M5E&Q@NRNNM,X97dO+EH<<U&OYe1=N853;aVHVATMT<
G(5/\V/TAc_]]fG-USX\R?0W1f=_7c>e:.<T@J7>#R9&3-g,<X\O)2B[B.W456)2
B9E4_)038A_?-U,g5PT17>+8P8@EdeN)?HLL5DRVDc&+O=\e8d(1H9@\^Z(7.)59
2P)R5A]<M-\J2UXTYTO[HOb)SW)b9EfK+g&),=Ge.SeL86V8#P/I>2H((Y8#2b[-
1)/1AC\JW]94dD8Gc=-[#@cQ]4H95:=H#?0A^-S\5a:BGV=O5Q1JgZ0L.H2H^3.9
O0Y;+R9B8IbJ:[C&3TAU:\PcN-?UAI_-#@eVUfR/;MZMG_]<H5G<:3\ffd4\e]ec
#\&GXA1XAUQA[AIJ=:ISP,1Hb77K1M7\7HOO8XKW)11Vd+,X+WMQK:H((3QGRaJ5
KX+CNcD15?RG]d#&C]1-RbR_;b]/18ZJ)\a\],[MgdW,3.5X8a_NW6<[01&\@HJ3
3J(WH2&<-KA+,D=ITdL3Y1dX_/_U&HYH[2D\d3<&]MgF]X^4A&D-_=G,;c4DY(b<
6,VP4#136L.=#NUWb\bf:H=J6<agR-PF)#cHf=]>CcG5cG\/C;19^_R]C2UeVe[;
e^@,](QOS71]<^^VIGK3261MP1NBXT<7RFY(FLC?D8Z^eU?#),8NVN7-N/[=9f1N
XRcM=:O)@SgG4[+C?#O2WF\X-d.\]7_Ra#fcSDKK(HUO7<@&UafNSALE[V<=\&1f
(H^@722^(6G5LHD2VU5f4V::,#b5FH#(Z8J9Rd^,L:&2UG_VO?bGb(-_Mg&g.SM/
XdF2OdME^ZTXAZ)X[/\=/;c(5-8_J;7dLH^66=5C_eFSN]06TF]UdQ@JCgeFdSK1
dgRG-#5fc1IM(eI_#ITNdR2-5Ebe2<Y5,)W9=@_[E,MBG@B\MCVJX_VM#DCd6^,,
.[4R;7A/7J3T::-T;JP&IQLe78I_DT3b_bcKZ55)<IMWO=.TJa3DdJ_.N3-[53V[
P?EBYD7F:_SV_f5YHTW:R.4bdd=N>[=aeKO<?e;CBL[+I\W;(RAOH\-B;Rg>\Tg6
b#LY(Y6]Z[5+f1(#.a2)4e?6Y45+\^0S=9IfBb.[Y8a]@,E@<)6TaEO7.V1T#DEA
PEbf+J:H_Q5RBLP-#B^[b&_\W,PR76-Lg-?0TcQU9\6<+8[3XX[fHe[\5CP)>I=@
S/@[be7BG&UJ<E]&0(9L+1Td9Q+g^E_][6)EIVIeg4/QS;_,>2#TT0FO#c6=DAEC
)B>H99X][R6RBW7<Z=\D^E_#\eT[<F5;J<H=;5)@A:P1MCKJ=6[#JGW8G?(Y.)D2
c:)_S?G#2]HB_/E0?4-=)G><B_6ICQ_b5R0T=6V3SAC^QFIJ7@7^9RPdFEBL:[DM
&J=<MMB8ca&GF,^-S#G2M2Z#g6MW24afMYJb8RV+6WUAXB[e;EQe8PUX][(BMbY/
E+>)P^GA;-^=.9^RZ:Y&dNEF12\FV1NfF[YW:bQEbgBK?)QRDd9-W#-\MZeJR0Hg
UGM+:M9#I?U>#JZTaGP8\,YO8OOO;=JL+0X.7+Y2X+7&?#I30KaM,_FgN)If^V5+
_RNR7PUbCEXHKHCGHL][>E-J,MYZA-0:B/)Y=5,Y]HW#=-R&W)g.\;B=HObP^#D5
W<59AIE43)CPEL.BH_f)AGYK.#YSJ31I<Y(X,g4R-SQ9_U222AC82,&[_IO@^X:\
6\JX(.0Y5^N#P,+bNY7gd:JH]6HVJJUS.MB/)>)2?aUR0NX[IBK8C/]QNN]ReC[=
b>4C8:.X/&1];bP5?d[:A6WFR^(H[@IIN0QY>6G&8(0VP?-4KDDF)0]C77aH[AZ9
PL]KINH9T@I>N6R7XG(HVbH(BK?,bD2Y_V,RV_7<P9D88b6d-V2G4N9C2PH;bZJ;
cEKRa5#<>6;.&W>.L\+F7[C>fd9C:e:N]4^,CWL)ZT_?M5Tb20IU.7HaAHVX0ZO3
fK3K/7XYg0Ma-<:ZdSF+d8g:WW(F4cN1^=?_SdJIO\@]7gf;W^.L&_&O67Bb00a/
O,Q^]I]&aP#9&>UF,2K:?8PIK7ab8O2X6cFHZPA=XFG4JDgNbO23[;>6HKH#f1.]
S5/a)TQKIdPJ3/eGU#U#F1_(E_#^>FbNIF+VU=7CF9?ca_JOG&aU4K8O=G1(QG0K
RR>:CU5GMG:f;/RLP?7M,2DbWB7FXJ:g-dEf>[GE(A:PM0,JQ])T?dSN8_E/@PEQ
FDg[4UM>ZE+5^c,-2KcJ0Z@MEP3Tcb]C]SeTCGDPY1TNaK.5VXDfGBKAV0C..I8&
USJH.S=C1@A]Y63/>\I7B/Ze\Y6FC1ZM=^C)/P<#1eDC74cO9EgTV)Z[K#8;YFWO
JWK>-^F;KOX?\HM&?5U7-O=M:FT=S=:B)02AY>P]]I\\1F4UT=g;bDd4abDX5/PN
1cU.EB7E>1#C5gNR&Fc4MOF:&Oc]9<bC2KCM\YF8&JZ1;d6PG7Sf=&;AC:A_Q7K,
[-JAV)0X&MMVRP/+,M1TCJJ9e&Q3@fEY5^-IK<3H\Re<5c,OV_BOPFX;Cb9TffV\
JU7c+]U3P>NSZ50&HN46>(9K-\A;GIH:_7NU:R50.>VB2egZ\O^6Z)<NFMf/bSID
RV3WH)L6D).2>;7-+3#cN>d_8[c6?ON2U7/1NR(SQ-CgO2:Y4V1_ae=7FGG@eU38
L\ZY>f^=Sa>g,TT?=_H7<H?^b0/bA:^S/DVCV/JK&VgB5+PdJL<B2_V]:CNa.CWF
)JW&DRDL#E(7F8A3WPbPSU5V_.U:7I2d1JB735+eUX16#d:A&_DL\NYd+[PPA)=5
_^I5.7-9/0Q[-[FR(T.:1g)-2;/EW@a5;bcBAeL7e4e1EX=[7QcCP/GDeJ?V@[8U
M&Z8_&8-NJ9,L^GZf9f]G=,G9N+?_ET4e+-R.W6^a7K\)<<6+aN\5N4e?D0cA_a-
\_QK/85YW6B1U]4B,W=4/TZSfAVW5NE3a>-\N(4RG1QH2P##F?)?<ROO45Nd+>+\
HMADO]KN@\9,5_)@\1UFDM?^F5?dTY5M7TLb,35]aI,G>ZHS1DA_5O/S93/+1b51
IZc.W0EG<e;+gH[JSM;(KCY^4VVWX\F&TKN[M?IM@]KK>T]eW6^a#c(MHYV(cFaQ
9;:0b6((TO^JV>)<)DO&C]Z@/Yf1f.CGL(8ZIcU;5Y[7AH<=d;[]-3>EN-/cV5#?
M5N=W]P2NWUU(^C@@ZPAMBAOV3_0P?#I.D86C0H/_8H9LGSU36)(EY63#&V4d1YV
1Kg(H1G?OKe<TbBTaIf\bL_(=+]BE/2Y=9>&Lc/)>7VFS^Q\0:D#5&e8_1AG2cd5
UJb3#I#=IbBY>/0Tc:)IQ&0_[CJ/3\&Xd9?2.Z)_@<)RNEYG?6;H:.)Ud2.X&917
A+/MaP0(Adf+f.0A22KH52#La5XOaK;@CR=Vcg=4_e\d9L&>+G-PaB5&CJ71WV_:
f:(P#d&Dd8#c/A60?bTA[Dc_UNbe@c4K,R&BbXS/Na:@2]>AZ-)C;\1LfLg_&,.?
4KZOBTA50JYB?#@U1:ObHDSGOgI,XJHZ\Q/XIG<)ICAMea(V,E,UXV4bM_-A<<[;
EHR.F\OAMVP#C3[EY;1+bO5K7ZL5W6.[[b_4O.51N,Q-DG;>>[Bb[AW_:]1.H_Z9
09g?<PDdTGZ5_0aDb\-,,b&(_[QT8-[(EA(gQRPT4Sg;QfE2JH@&1\]T[>[KR<UT
Eg\b^=e.,=-3Ya0HC:)dV_W?T?.?XXGGNdHK2e>+>]\E<L:Va7DdU\4\S4W04;,Z
6eL?L5]6@JMFZg=B6RXdFXASYgGf>GFI8Id8UUVV]d@3THg6\@9A7X2]a.7>CQ)A
[ge_WcSeL\0/MX11=3BVHO7We+J;9UVd>\4&=X/1Q@bHa_>&Yg?(IL25,+6E,)EV
MC4NE.SbfaO.99I8<0F;XL18NYX8ePN;_\MYYV4VB;#/WDMgbMET2>GG6AN[ZZ58
=7-DXXX)IVL<(&G4SIgMA)aJM1RP]CC7I=@AL@>]9FZI:AGJ50ILN5F]K?_a;.TJ
6d;UG=IC]41aLWW-)[BC6LU@^]d3a2UZA1#\C<ZT7,Z<USbaPOgD[.;G\BDJQ03d
J</;<Q7AW2Q8>?6W9R5a7Dg8Q@C+:++/6^+d6bH-,A0V.0AR7d82<@eCRU8T#>Kd
.=UE<fY<O[<M<Q4,Xe?cV)LNQ_+FKT,&0_II&T8O&L;M5V(GDBWE:#&GMcG4_@==
;ES<642B63>KKK[,IdQEU,J?8?8XMJT4Ed_e7O[2\Q=J#77]GOIaaJQfO^E#<aF@
fY@&JI#VaA_VC&2ELZ]IdX[gC#T:EH^<_<F_eOdU55_bNSc<Y5N)G9==#RZ8?HT3
^fJ>@<2+V.c:U?gZFP\[aGgOLD&S=C@WL&7W:f&2cb@4<X0Y./Of^d=7H=&a^<KJ
#g&X^G,J78.O1e]P7:CWX.I18<bI:C_6A/,[FK05N_:FE=>,bO(<#77YOOT??F2F
+K=_ZaI=V,[(LaE[TZM7<A?X<US(d+c:9/D+^YJP9,LJaSC6QYS/7^/c7Q:Z9:C7
X=&NVRZ1\g+cFQ4.VQ@[3]d>NR5H9[aCae6/.8MJR)5ReZT+)O9V0;,f?eVV;VZR
@e&K-ROc;;gZ]/SZSFO0+ID:dC6J<7.+=5gB<,eGRG(D3UE,dA(9,P1<)19\f^P8
f,N#_XRUb;]R740T3RI7U^gHeEP9#0>2Q]>bac/(-VJ43?@E5g(_12CJ,_-cKYI7
Z([>:6)U63PSLbb]T(3MZdZ>f<4=?D&Ec)9&KIJ9#U.R@(KTVP\e?9Z;e3C._UYC
A#KO;6)S8VL(3R5NZYRORVX:U@&]KAAY#TR+O9=XS=?;=@MM4O&->4(+9KdJHMD0
]-E4>BGIV)e(AB35//ag0[)cFT0bC@2:]cG:NLbZ18CXSdfI5B0#>YSaTU]>(=@2
CX5M-.JAD2PdgET-F#_=FH>C&K&;31?dQa4JH5.WW,1e@._4.YH+.g/ZY?S22QNd
C@Ob2KX1SW>Ua2P-?A0^R#.Q5<L9IR2Ca7#;d4#/#-89LDC-cC-b#0&\BK#32AO7
57UXeVB]<>c4f2N\=<=])K#BZFZd=aVWK^558A&FG&^K)-2ZP).+_9@DO7=0>]^-
?B=ZEF?9S;If>d26H0IF5<gB/Bb\8OcCPdK&4>@cAd#>W,-D+]HQ0(^D[5aY]9S-
Y]C(Y-,IeHB:9MC^CF+IR3^4FIM9,MN:[JCC[dSa)]T_V@:8J#EZLO/+F<\)V&(U
7Na6::=,G7\.ZBTOb0;0D1Xf9+6HKe#[27V]M#/WTR8g1TcA=-XEc5IY?X40^E6-
)b^fSXOROAJS/..Q<)^AKKTI+R]#E6T)c_GP4YW2Q@^&U&>cd79(XA(6HN_-P&R(
@bUAN)HM?;^B[L1T;Yg.D8O,6(#)g6=M<QS-AaRc8GQB^bfP-DZ79<5?g3-Y-TFZ
g]L;@J3AWX/eU#1HVO9T4T0N,&@VZGIaS569A76<3f3_^K?(Ff0H(JV?LVCO5WO?
HAg;IZFc<3H?EVUAFYP;HYdA(EIgN^30We>O)+cEP_0ML^/4e6M/HUZSU10<JSDV
)Q-KJ+4^c[=_IC5+6(KCFfR<I<)L<XTcT5N;^J&eH5?cObH&eB#c1Pd2](5aLWI1
NBa5?d3Y1/K8@G]F3ZfcL<P\W^7@7P]fBB6(3aG:ST7=\[&V3-V78I7B12:)-F73
X:QX+4[0\F+OUHY7f1G:<P6@bbC=;+)V)P90^?WK,MC-<-795XLfSY&cS];T-EL[
D-#)]1=b5>1ES&1a[.M70M]Egg^RKD]46,CWf@4[fXE-:IJEfL<#YIK35,-4E13e
c25ZG+DaRHVKc()QAA0SU#,aO320;SG;>9@0faQ(TIfWF=CN3fD_4CQcg5R?-&J\
.)Y_\UXfI1DbJa_5T0I&@M2a+J?/-,ZQ20_@eSfB?g]_<E^I.XLH:.6f]=\<H?/a
S:eQOQX/VW]N;b\1Z0>W3JHKVCD_SQ_ca8E6O49[K?P&I4Pe.bI]Y;/G=>T)K)EX
gP7bAaD03QA.#04QP7@CN7-e9CA&DN^+g\Qb,.O&0e3A.#fC1;[YGcPW86(ILOE:
0a/Z3G+[&&_<a37J+VV_7.Zcd@@&^786L,R-_;W/7^M^#=EDK#>(;IT_FIeJ<__J
Ed-f6MITT,0@_We+[P)3Wc/#UHcf6)X:3.)3AVe]gLQ)Ef>Gd07?I)f2P(4eB9M3
RO3.8FH>N]-=--3F)D6)IZW1B&?P?ZOXP_UVE8ZK\ee]J_W2&-]D<UL0YC[CG-HZ
[+)Y+9EI7PbJBUETC?A4g@900EUZg0/S-Q/M+RE6cV[;b@6\EA]LBJ2956INPM#2
@E5[VUd0Ua3cVc]SPH3]CdEXUeGDc8SVe<71::71GE&/+8ZaSU=b-7a&#HK2c(<f
]7Rc^@J3HI.gUA>=I^JdTOH1AM/EO.4Q7^BV6S<QH/f__9GScI@/NDCUcfJ54/9\
)3,@]CbE.TWTORB_R1TI>93QG1FXXf/\&:?RAEg@f=^BBFe5AS:\Z?MJ77<;+4U:
<7_L=5V.>EYW+).-2+AG2&-W0aLUcXQ1(]bXfTcf?-U)G(S]:RR0(H8CX0N??^5Q
._0=V+O:MAS+_6\<g@2P)Q:agbRa<&3]eE@Z/cL6KQg,(&d>H?Ndb/EY@+Ad]1;]
<]/>/>7=]cX.7KY,,Y]AE.e5>1I[:P^.C;SA\d4][077C4dTPg80XKA7?XF?gXIW
3)Q-/D6YH43PTS=EZ<a#_C-HU^F0K8\N+C??#T/-b9^F^E4..?G,-ZZ[>N3cO?1E
YRP2T256I(+F_UD/U@?@A1;D#TM7HDcHI7QP[2\&bOBKL/NGd:#0?e>a2d-E/:PY
=DfX[&A\RSTcDC&gIDYTfC3=,fC/G#@Fd9e<CYDRI^RDNDHM<>HFEE(fZIfQVO#(
J.;ZE:#ID+[B;?LS=VXKg/K>B8:Tc5W7A?O:B/]9..71@,+1QXL#Y&6\6<\(AMSG
f[c0Q9YZLJf2G27_>IL2C>b2(ag_Ya1KG8)8Y3?ObPEYCd>0dNR5W=6f2DAUE>P7
(dENGT,Jb4D[;;fO.QdXB[L=1/-^;KSeZ7FS-?7PNM1CF,32F)S?d[DCK(6+Q__Z
V2Q2=)K@6(ZPV6TdV2TPaZ6>PL+V[I5M29SYGc^?#g&FH1Y3U[UG:\)GY8(;GNZX
_58B7_85:6W_1de;>Kg-OaAb9:#Kce(OR[dJYK@3:/R:\:YfO]XQ4^;Y_C;4f)CG
>NN\d9]U=I:3/>CH4?OeTQ]#+;d)C-RS9CBT#P>IbKVfeB5eMA6.<>S\U=KK2N\^
D^dV(ZSH@e#3Nf&0b^LASB^fLa#b)K6@^=W-Q3cI&5LVBD?0W@3250@dK_7Q+.;&
^TdP#(?NV]gZ66:LYBB):)P_;^Vf=U2BRVPVA77;9c^+<_-L.^V-(aCS<b]28)>5
R0#W7LG.:S_9N[[YGC,B#9#D/MK1NUN_3RBKH#Ma<_F]@eZ.XQ^e-WTC51PS;WF>
,I93\21dW/fV3)6^1+[,)XC.&Y?Q=bFODU,.JgGHS5e-2&dBSb]b^_:CgXMS:P31
eDI]K=5;O-XW+DX02F?<e3@TJO:bfC-Gdg)d,S2=>d]4J/S41&C@C.Xb.\+=g=Xf
86^Q[WUPOBU,/5dSMS/O]&5;NP\a_.I9:_[)2DJ0CR=M3S0RJ=7#W&Ie2?^@@G6(
9?_Tc2KS&QN1@FgaCT2)BU1cD^1T4XZ2Y0)C:DYd7HI<&LQMURF_^Ra\N#5WcPJK
J)E2QQ9Wc=[IXPW<3E@NOV?,3JSO^2;(>.(f:2J@XO).G>gQT0L=SF&8Q6E^Q]2Y
?5;KQ+Z&N&SWZ2?af>PDN8][AH#NZPWd:UZB;7_7D:_REAcP[^B(;YKL7(.0SRGF
BI/3g>TES,M5aXJReQ;5XY8fT1gM=T_27MVL.TdP=951c[+OJ3PX+:<MQ:P9)TTY
B9?b-]-:?-]K4+c>GKe2/NIab&/IC^&USIaaJ<>GXf-e,GKSU70SC0.94RgG>P#>
KK^^Q(Y53(OZ3Z8ITd4FCAge/=V994V5@#aG##=0bDX6-\.8/@b(bVGOI/.48^La
>N?_eb?c)^A2(<WU3C5C65Fa8SVK,a<2@cWA[I-#71HC08JK54C._#^AV4IU3;Qg
R+3#<RV:Q3^)##TFLc(LEN_V?8H9,AH+eb)GVSK8=<Z0/B_M#TI^S7JT(b(;]HK;
+F3,=#;[ZKLWY1=26>@6f.T/P8&_0/4TU2E.760^#eN9)A4QV9_6^QWA;/B+&AE&
C6ILf<<PL^(@C&>O-UN>fME]X5a899?<]D&RfH_=E9cgEG(1IS@S[8AQ2H>G7?=P
VLGKV.Y1Z5G\0?F4SJ3/H&3H)W1#\IQ7JKF<TaY-26cP7H@XJG=_;JDbOc4T#E/g
F=?J,IfB/e&KfI?b\7?d3gH@gd?&#NbQ:H-8c_F\PBT1bC(/cH1((DA,IN9#=\e>
NN2X/,3E;/&V-1X::D)-;0ON:Y=.+bG=eZ;1KP-bUL<,^S)MHbb0eD-+PBR_++TR
\,,TU#P[c7fHOg,DHb24+9e&R:00=R1@cT)S>ZcF:Ta26TNPC4fa-]1gc-EIa228
b70W4@F9:?1\VgaH&eT.6;1.Q,c4X#ca:+-caHNY4RZI3\YBX2+[2^4484c5(:a.
JAEAH(U@HI42+OWdg:B,L#dM-CX\1gbJNTA31MWI6LWB,G8>@Pb]PEO3[-Z2/0+@
4JY??R<TSR&&-c8ANKS;=P1(POd(:O+<GW3PPNQ[M>PR2,.11;D^G:&g3T7:ZO&T
L@]I:/d4639]<+L:B9Xd,bOC0JO2ZaTcc>8Y2c&24]>P9gI=JVNJ<,PP+?)DGTKf
M@=b0]8Ye+;9(4N>\TE-J,XT6UA1RY;T0HR>_>cEBbLd:&94RWHaP+F)G2<XL\/d
<V_6[OC_JP(Lb:U7X8:DBaJ3[PC/S<_<B\,gICAI)b,?4e01c7b\3#?PN&#/-7e@
C_DA1c3;A((VdRXY_CRG5VCQ5<0?,YB]L45WC\[R_>a@OC0HPfPf@LNDAX]H##J@
;5:HO;S</U?Q(/KV4ec3<Ob;8D<)1Jb=Y@J@OVMU:Pde4:OY[?VTOIC(-F#&eJH@
bZ8FELT-3J3PSUM(+L2SbUQ78#B/[SPCA(EN>AZJXQIV=,U)__?^6-MX^:dQa7#-
A-5gUK6a<B8>1-=R-:6^;ea1;O+7HO1&EOZ@c&I87C.e_#@H67g8XaZ&:5&&SKE[
e.GVWIF<aA?2[<,U^;\^=_SQP+&45(&QF&K@gUGG@>2O(d(X+G>^S:&Hd(C:@c\G
Ob_FXVNSC]G0aJ?DS-&Nb?GL/,R\5)FFS0feeQ7)#@C_6M,+0TJ>1b+TEVde/&GD
NIHJG8;f&0a[f1[U^>\.N<IN]PJe5V)0c::\97DMG@We[<AgZd>(1_52IJfK5-.0
Z;)P4^[RQ^M^,-76CgB[TaHBLD2V3b^B?J7?cOKCGCS(SU__g:-\PM9A\FZ&?Q1b
gJAA\d:H4ZaO(7OHe6MYPfL=\?Q-^^);]7b+AXgC[^TJTM-5[_&@\0T:V:Z;HF?O
SWA.?P<D92,:3JIDMV>]N.a[1.G=/05LgeL@fKX&W/VX@Z+cL#U0MN-FR34JGg.Q
;\7&fa/3]EOE]eA=852fZ+86]71T8A.b&JdHS2ZS9ELb>#,@eTcUV((G]^U9-(96
1TZ._ZX\4Oba1[:bP_3cXI-PO7@@-695&M:,#=BAadW2+XENO-4=GYZ=RY=LC3#S
J?5e0B2_K+#5#cD9WF3-?:PWHVMYC4>I9RP@O<4FQg.5)U@N>N7)?)&(D+8ZH8N6
IVJGP\L)/97NR5/\^e;@OOSa31X4@PN]_DS0NK@9U;OLGG5XgNT2CB0DN]f\EGVL
XAA6HEIY,N8aE4XKRcB2>;dga1C#C546.J^^]N>2^TK9C[?ZVY<J^T?f:RG\MZWY
MUDO[P9X2X]KV\U3+=/fDNGFM,CTQW_JBd3YLEE]4f(R@e+D_:ZHHag;TRX,BVW^
VfbD(E#_=AaD9YJg#VHEM6[E4#aKG,\^E(>B5&&Z+2eX92VM(&)bH8cRE4OB,4>P
LJ#4a\;IQ/?U3W5P?cBS,>e5/Te]K]A@?RO-NN^_;U0_Z^P\H23a1<,=(LJM_SQ&
67Se[PbSY#bIDE6C/P3)S/X<&;,:+(d6,<S8]T#d)3.S9>DAA7P.PI<(Z8FP69:3
/N?I;9E@6Mb4O?H@#RIP.KE8@KKY+TH8/IC5/A]OT^N.O3&/V4Sb-#(T=78YSMHC
ZVJ4Pd5dWQQ5E\]\aN6&/V0NE\c]/+#>N+^IPbM69J4(eg297Hc?FTfN(04EE3#8
CI1NX:[@/WFG:O/V;87gZTEbZ0ST0-;+P1WaW(OK(D(AZSOXb-S@/\JX@+SM-3S(
^&M63OB2<3SB=]<bJYaY;[+)RX7L6S9<:1#2S56bT;DGWH3),8dY3WTWF1a3-.,Y
N#=OZdaSULSH@U)N9IN68:0#\.WFH16/T.BdR-+a,G;CF+b^Z3C9=HP3\E.=fMcQ
f]3R\KQS]WD:Sb?FO4=Uf;\JEJSC=I(eaJZ(@@L9-e^eW+Ke-ad(2L^-]9ca1L?Q
:b_X09fG@;+O..Y.IE9^Y[g@;Jd9+<NDL?ET#M4VT4O/+eK7eYKO)[1&8:gbX(fO
gLfYGJfb5c&&,=/D.<-VF4^GL&>_D\e?/W7T:A[L]g4Q.6<>7c;V]T;QN9QDFJ@F
gTZBEO\E]U5@=O:N\(/7Z_+-.bK&S-K6-U1HJRDf.Te;>RY&@^>4MN3,?34I5[6g
6dE6NB)R=SHPdRSNKHVW+JM)^@LRN::)^U<NV&cFA?eSG@>5TL2EU=?__G+.d;\f
&9E3X.[R9[]DS8P)X4=/07TK/Y?7C(PbM;e;)8?6E9DK3.9J>JQfRBf8:Zb(U+E5
DfO#Z8F3b88X<P+7GRB(=DDGR&U1WCS[8Z34)9WNO)R2c,9&^8ER[OQ^N/42>aO>
(W=<^;=(\gXg&]D=#R\P6UP?T?,<ZO@-,cQg&.We(W@#K;;Q98d1HRG.@cD1_F(U
A=Q:b@24G(a_R7D]YF9-)-9Ca,9bbQHTMO:C3\F/VcbX&eUWU+<a/LaC@d6LKK6/
)f=b0G-F6;LJ#O+#Y:7JQW(A1C<J9aR6#]=R9S/MS+H,1WXN:NAd?Q55gVf8PFFA
O8F47X+K#\48M=Ke4PP@TK6EQGH5-9f:I_5Meg6]6;fX5a7WMPD(P[DUgS>g)5V>
+_5-g2@H10R\U8GbH6=;^HTI_eY0_(74/DI9RF,C,cH?T]EM[a1L95A7MK.[I]Tc
_e--+B8VD[Gf)OV5\N3DPA/RIb9=#dG(S\fPaNV550X?Z:=>TfJ@9.#B1DL-]:\\
WS8#c<_\D66QT:X[(UUV1c#]Y>]^HR)P;@7IM5/J,FOMYbC:)HV1GM@;P4[6O#>Y
T_AFNbdXK2AY8dS,UONO)Z/SeQHF=A?V9:HYA87VPT(?[[P&gIT-?]Uf>,G=KU:T
G42LHQ1[f1OC,_DDJIU0)78IQM@Q#N(3>CXC58fU[Ieb3W[GJ<IE\.SN0#XD6gL(
I70)T3VI8)5_bU6TX5cUb_E18B-KL5>Nb&FaA.])@:cH?BX=QE#7FI#O7e7U,^8g
5cS2Y0C[[+ZQ\cENDRG.0<--C+L<fXW92P;GT7aFQa1/,P5JRKO6dUL/Q5IYe-Sa
RHK[;JHSNB/da-2W\<&0MJ<?1Uf6OKQAe;MBP[L@7^H0f^TGTK5XdTe((^]CZ9\J
<+1HH@a,50OS;_?[7PE1@3Rd/6+2B]-TT-.#6]UJ0N+F/SE\ZD=:C@<XW;05<,NO
&LP2I1?7#J+fO9DXd/.A_><S;..7U+E3)CN8[=;SB?OMB-BL]SV<Kf,<HaGLNAVQ
89LU5<)0E(M8UK0HHf1BYLb3J_M?.Zf:TE<5?SCQ31/R#GVZ5<^(f<[Z@[&e]E[?
G,?XbE]DSQ+ac;O,WfX)cWV38.6Gg4LLS4X&H.g<>X3&4J85V/QZ@cWVX4<9Y[+,
JZM\M/:^US7]dZQb:0HEd6LUBAID7@,1T0b#WI+Hf>OPIXGB3E@c>?W/EDb)30W4
:-0?_7G])33DYB?>;52_KG-0#AO2\E82^\fG6>eI3=EB&-g\c/b\O\fJVLSf,/)c
&]FK@^SG2M3eTUIa[RaaZ_6^R]9cN^:[gUMeLV>dN5-ZK[0/T<Dg##C&U@G.&M1J
2VLR3;F7gY,CM;>G^G=Jb#X@#c.^/QJ0GL)\66MP5WI46IbGC[\Z\9?SA0M2&U=D
?=Q-A9U,VJU4f_YU52QO+R=X6IK:?7URTC=KF=MAd>Pe#Dg9CD],Sb>Kf.R[dRV[
M9OYP8g/D)\@VPUG4Y@E[W>R=O2#+F+FOfT04S.f@GPREM/4.UZ?3@cGVOg@7PRB
c:TD(VL(E&DBVGS2G5L=f:._\3;=^Q_XGTBaKE91bY7Q9&7bb^B3;@IBAe0#@2O#
Xa1FHf1O)V]TS.Q@.?XH:7F?ZORbJ)f#/1<R[49b(Be0_\c1N1631IC^]4>QR,-C
ZXDc-7OV&C@,W&5Z6N^=W:Z2-=__KX4Pb(>Y:H5>_g4W++We,1ff^M#YNDQA-L=b
RVbI4QH4TICSQ[W6/dYa-a<OfeTW)Q6-&2dAe9NRT5LD4M1Wd/_<X3Rc3-cNLbG4
FfDS6HS(0Q<:)15&a>Y9:Ie@_0fBKO5N>8PZZR=06+(E+PO@21cPQb#G)(VcHPIM
[bLA5)8(Y7HNT]=/];D1Y;=d@VYA79L#40EGB+/F,6[Ad9(CaCI[(Sd:8-HJ2.MD
,NUKA8614_Q2;XY<gD1N2TaS_C7)LS4<a(S^15779fe.c_)bCa/Mb\D=L\M+^dK)
S:7bJgTVb-N(#]9N]^9bFg^aT90FXBRKeR6)7GH44YOCO0MAA7_gY3NKHYgMZ77I
:5D&?a&&K6U4E)(+MGG8;g9_Z_#c.../4^A#A.6:@/X0eeE^7K=d]-_[SJMYYP,:
[Y5C3+KW]MR3AaRBY\YcbLe/a+P#1f5T)9RB_+,6JbI#ZAZ;W]JU=O)MGHH;,28J
XX;6UaQ4gO9^AG_=WJCX:?SgN)H&W:T[WM])H7ID;\bU9MX#OM3ON1,==d2<<QV4
B[^GeCTU;g)EE+B08_Y?H,g5g#>fe&9d--.8@N@0ecI9_BDNfZA>F:O9dOZ]S.07
W,>7)K5Vf8F^<Ye8.ZRY.ebY?VN,&R\>.2FOL7/KG<HH21>H2JaT9PP1>E0<BYR:
K#@W>B2V<5C\JFc:FCB(\N48cPfIbGEKWd1LI:0bBL+=@]\VCfN5_Z\ScL[R23GG
]g&b?X/IC/c2B0YRWQU9b:6G\V&?R-1I.1D>VTB(+0dEgD^4P6:fK2BQD[4P[@12
\T^Ed[4_f0Y@:H>@5ZT<8@C2G?eR4)8#:WWa93FH<XOg0&b3DG;:3\ea,&Q_XS2)
LD:TBJJXF:[?:.LL=:,bLZ?R/4W=01LU_;I>LIUC,gJIP8XNWXCJ;:[VWZBLR&,1
fgAf+Y87<CSPH<9dO4]be?W3VJ,@_3U>g2W.0NaXN12b2T9Xg-J]G6@]>J.7F,_>
?WFfTcQ<-T7+f+[ICINSF\R=6IR80/CEaMLI=a)Bffc9<M?G;O[]<6O[R1&ZRXK.
\N)Yc(e==><N&_J@F,XM0DT];2(4]XCFQBVGNCAPJIfVGKK-QEE8LGPQB>]5\?8V
?2A.L=gM+aB3c7[2cPM<?;VfF</\)[YS1&S1<[^MXE/,Z&67-,Ug?>@_\-ffdD.#
LVOE@d?YM]8?[ba[2cFTE2YP\T8#^7?5+MRXA_ES9I1/TBLRJBTY^Ic>@J37CD0?
@,&T85WP.,RXRLD\,XE,-U13c600S7B:-NAOZC1dW;10RH.>C^L,3QY;M8><.+GS
K/VZc&0.=ae24P\RcL)TE=V9[\<H)?a_6,3MZ:H/@>eO0F_fGLI2QDZSBRZ.F4/7
BAE@+JN7a:H9\S]4/]3HO=ddb<fdYIFT2WBM0EYFcf=Lbf1bdebM1D&NRdD25A)_
3X@R&]K[Tb\PML:__8T3?,->N\)+.H2N\&;N5f;N?>=2?0BV];C1#22e.&,K/)35
2eeT(<+=6H&UJQT18P=).Z@BU[6d?1W/EFg@6<c,deMB7-V=,J8c(DNV,XLG,H8M
QQ_SA>HL.Q,1PO9VW)D:F:\\^JSg[I@BAKc?IFO&=eg1N&a?OED,\8M_5B\1I4;B
NR;G+0)S2Z>bbDJ3aLFfWZfQaN&S?@=>P&K5IK8^\.JE[g9HB0-d9AAD31_SDU=3
-7I[29GO\2/Y.MCT;f:8AR\FRU]dKMJ)8d1+bO71/2XU9UP#?RW>-Z#,5QK0RO<9
]C\d(DcdVBKYGE;P((S7I#8&<9;YZNH:8<H7(c[[<KP9)3Z^dL>>DZ601eMdb,3:
F-5LD)#V1dVPO)>96C38OcA?c[#EH=,8B(8g5;8,L41P8E=H)1aeCIY8)DJX-d].
LP+G=T2=,A3M2;#:BXa94]d^(XCeM/Nd7:,DIeXgGS43:T-Z#+[;\b?7fJ+DX<CM
8QDCfVdGJ\V.RC+9]/QA3ab-4e6>TT:O2XgAAO:O1MD&S>ZTW_.S0E?ZOVF0bG8g
.30HJ/EQNF0:^KF90_7E<MU<LE&)XF?;O/0AM7b1OX:2\?.GG,F&/+7GS6W^&B<]
G30IN7OBWTVE:##4_83KfHEL5C:Z2E@^Fd]+b[YagEP)OO#BU6R<;R;E)^-A.\&,
ES\0>]bgE,)LAB0=NDS>acAV^bD@D1SH-dE/9,3;0A7FI@:7NDQ1YGd0G-A,D&VY
THPB5X&D,bV9EPT(K&C)TC@CQ7cWObR@=DRLeXcDXG[g3M^+W_FFEFWYA:VP\:e,
<;Tf+V1/H^H9WDJLP-cJL?VE,MM/d.GOHbE#94EU\FX4CQVCN/CL9e@]FH3N)RJ7
+V4&QWMJQ>/XH4f6ebGbW,_\e^S7T#dF<W.\A0^/B)\H96]e7bN?DTZ-dN.V9Z&8
6:KEE:-eRf@\;L?&UZ8:4D:fA)J]PdVR4^R8L]a[?/LMa&V;HKYe]2<_I&E:&@6O
S\)_Z7AN\BJ#VJFEU>9]1K&EH_;_IL-62E.bN94:FDCG/1]^G(FJ#2RB3&cJ0<(+
9Ce>.UM]Q>,&F0W=c8[^7]N,F>1ELV+bZ5:?:a-IFI^f,&PHOXU0R&_PAM-g-KH.
#A_)X]9]a<,/T;8I1XZ),F5gJgg/@HI.UU6R7fW/Sb+NTRR)EAb+W1Ma./=X36-1
NQ1_=aDW:<2Q(#SX:JeEf5>#N6[A3[D,DbHM+JGUTW6McM6_dLMb3+c3Q/SbBR0#
fMbO4N0eGV?7[Q,3G^DF[V166fO0AV(,EYAV?Mc/gVUg&VE^Z[bREC2EU#1)#@]W
7/QMJ/cT+<6-QVM9KHV0_G?,0QOg&EV>OK21UBOaJ[ZIN-&EF7MUe,7Qda1eQWN#
OG-egLKUMZOH91#FI,C46RS5dD+bH.FZP^S/^/PagM(0;c\.\@;^_I^Yf,P5\VE2
:bFf)E;DMK@(8=UP\DTLRP[<cM-I.UF;VK)fL#KA+>3LO6@\0Y3+<@Q,YCf;[GS4
e@V5.7PU94TT2^3b6;(1-?FCJVT.dAV8Ac.F14d_H<1OfKF9LM2J\B/,V(GQ@I2f
c\BCLb;^F[IWf^LI@&-J21AWE1=J3aGW1dJC.c&JDfVBXVc6aU4^;QbAPPA.[Bfe
FIFQ[3@+@:]8BD:52IA#7)NH7ZO-6T=4NfHX.XNLR#?V4;I&^@Z]H[4BBd-XW1V?
F9EOX=c#21d)YI1aP/T-@GE3f:ED8^>6e-?1JDf:+;RK:a(Ka@TW>\cQf37/BD>c
W47^5+.:adOC=[7[0RB7,2BILMfa7N8^\7#3g(DX4,c?CF1.F((JH37?5?gAK_D+
#D@I\Q7UPa[85839eS/NA.:4HM#APd6gV6-BcOIN+:W/;(ZMQ;-:A2>&UXG](F@3
/64R6V)KBcXe@:[d;_=84^e=<a?6NF0ATG4]+K\d(R-G4;3<HKg/-6?2eL>>C110
g]]KM<<7JAU=\:+>F<BX3+LGbRUWeYf+-Y.B^R@(C/FJMg6R:&W8,(L^5eL,eGL1
Z#P1N8QJE6Q:HG^-Ya]Y/AAZ1e_N,1ZdU97^]>VE]^06,F_FJ;Ma6WP1#X1W]?Cg
+?ac?1f3;8WagZ51Ke]ab3RGKb5-g7N?)FM/EX:SKf3&Q60324gT2BcVNaE4R/4c
OcC>SL<eQOIf_-aM5ILV&E6:H^J3.H6F7g?_YQV-O>1+7UJ=U\9g=TF(DVBdbRgT
d3dFOWP<.&)g7A@CRD-d./3D#]W/87G]0>BdOE#\2S)W_B7Q7;VNY#5KOW.J[3G9
DaZEHdYS(TZ@Pf6-BQY).D^Z7^T8F^L&O.;3Z4K<H-dPJRN)3BL6-ZPSZZAXM2(+
+=3^BA.^12EURCITKbEb5=LQ[g1+.Q9(MZ<H\?e=-_3/6(GFP0&=d]@BP+:XQ0@@
-QaUR1]@1]UFF28b;;@cd_BVR,K75BC@NbY22P9.D>QRILLMN@_5?U5;Oc0UQ]bQ
eUNZ1OPWALRH8G13K#HOI@e=6c;e^DKMOE^Z@KDcP8RI;5]7gI+BL/YJ7PJO3(JX
D+O9UID9@&1[.4/-8LX&F_+VE/5,M-L^YJeW@QPP\=DO]=#1B?B9b_ADPMS:)41e
V6eAM\3HH.K\UM:0d)3#WITX.DED#<?.WbX&.c]_,\UC)2UU^(D)8LBAX<3aB0g^
-8VT[Z=RfbA==+gVTO(FF.)LX\M)A/29-31-9fC2ceB_)\GN3/cMZBQ8a739aff/
:UKgWB^_:HEV0gIQfY0<g_<FZ].RddT;C8]\:6J752&SCNg4ZJO>C5_d/Pe-[YW9
P@7cO.1Z7g,35B_AdG^QH2d;&E_);QYMSEB?ZD_R13+Z\F[]FP36A\g,>HD;\XVX
_MKMV5L5[#:McGNBaJR-K=4D9eU,D-I93RH/6S\9E<>]>fM&]&OA(>@&,\dIU55<
;]eOSCM=M7(AcL6_TOJRZ@5;AC++CCg2559;>Ne18FO#YW,-65HG2D>AeHOAF4HU
(<8>FaZ+K\e@cMe[S-.UAE[P^c[gI^E8P?A35U5E3LFfc;f(>?8D5e7S2cE8B^TM
Q[0E^D+geT??O8a5>Vg\<8KH9+=,#7]PU2d1-F?-^gY7+?fN(=UG6LPVTdc(8g@e
F96aCU^Mc\0>[YP]H96+:_g@8:[3\Da52KH1;#6[7&E[:HD6X_-W\+0(NN99LG>)
SXd0\Z+(cS,0>MIfD+??_YW1X#a@Yb8GPbf;CYW=a,JAJ01BJ]M.^V1:>-T(3fZ-
=2bUO?R5,6O0#W>]D?FMT6g:H]&bFLR[c=_VIY_=4T8@OSTO5gTPfBLB_MO05A5U
#ZIC?R0OA3H7/^YGEJb?Y_L]RNI5+9H<3=O2K\YG8f,X8HK_NF1LE3bfX:^2f[E;
6O0/e_L:5c2LZHN,&RFF_JMc(-KN:@<Y]7W?R5gT?(R34=Sd#J_E[1[Hf[&)M2f\
G8T3@dQ@fG_(bMK6e3C?ITG7P6(&CZ@KN_]V58))7A&>d&))A9g;I?#GAB4+5>1]
^^(=><75B.Gb-&Wc^XA(P<1aVa[[QB+ULP#75IS<&#\M)Q&?#7+#@8_Eb)U<^&=X
6bQE-<b92]>&/fG8gUL+H)5e1O#OC:cOA1,7[0V:SB4@RAcQ=>CJcW&Pb;V[XfJ1
XOC99RQb/g>1dM8e(0DZAgUMTGdfG1g0K(0J^-+OOZT3)J=Zc_bI:@UV]eLFS5a(
PGZSV3e0+3Bg:7+<7fI9J5\f?<&gJ_YfcKD/^1a&VD^T>fD6[F@e>4aUJI,7FO;2
.E__;(:;&631\6U4Yf0?LLCAKEX^D^UB(F))Hd_@1F38&,8-S(A@0F6be1D_b19S
Tc,aX]:GfDWD\+92;+<R&e66\/d56=FBKcK_c^ML#g>,OP38Ra3B7a/[K?7SbXLJ
;NT(e-+\97;JB#8_[UL--,S@^6><0]H?bI>(-HUQ23BA,9T^7-XRb9DXAJ)QS#:D
C=]?GJJQVJP)5R6T#6d1g_F>QS1AVLAG=-26]9E&-4W;GU<7)CgL)bU]<Q9b-VN;
c9fNHI>CZ?6,@b4#WQ7&_PPCZ<_M17eWO/C9HCL20IAH9FK8V2d-f29ZBGDeeQAW
[PDO:f)bV3a)(3&G=)PO7c5;dAMd=R+T\GdTNZ<G\0)7#WQ(C9\##L]=?4^LdJ@+
B[()[\/QHfXg8-EV;O#gfRgR^fF9LP,#J_6<Y;#2TPKg><:?ab(c]Y>==5&.(>\&
W]K[OWSFCI?.R=d8#=;&IM<7VSP>P/d@)R,3R,ZB/)#\IKD6e;3T.8MEXYBHBM.U
N_I1[R/3NL#^YdQ&YFLHMO8WL1,[2g^Ae\8]JL7\(Fd36,>^(Y@cYA@Q7]R_FdcT
0e@).c<K(3C\Z6#]Y^S)7PN#=e?_6A4e9bD1,AQW]/,2L0b((AFg2)>9EP_,0DJf
.2&U]+>]XU]+8-[#B:]>057=g-E-A;A8.cAA7M-(=)9;4L5>?.8e,g7[4cUb=(6Z
E9,\f-<IK2dW=R])dY1\(HXV0]ZTOB?8Ha@1VAS>2::.Zg;#EB-4Qe-]8MQQA2LS
AAa(N(7b>Y]:M<R5\POd1I[SfKJ8Y74PeM)HN-V=#&GJ1QKXa69);L:P\JKRQ(R7
9a+e6R55?1K=^BbY)9&:WNe7f[SEAA_gG6Q.=1aSUZ0=XUcDD+DNPSTNDZY@()#R
RZF&.DOM6/9_HUAFQCF&>A>OI/+:^IIYEVA_I)Ff.\\7bSM^f1dCEA;;SEPB97-H
)_PS:=.UCPEaY7;E3,:2NI6b@JP3&/<b:MZQ>+\)Y\QU6^(/cN4YEUM2\#]edg(I
#>#=X9E(96V1S@[<A)5^/f]T,f9PX>-C8N]SON3#dcD_Q=bC5L\D^:IJFYgCUU^@
?DIg0c0N9#5I3P65-^57UZ^&.S&O32U-D5#G-)(a@XQZ/2+gS\:LQI7#SETEf2VL
Icf0C)#P--#=70f7>/ba2HaLTV:RI]6/a-M#,f13/50cLS.C0Ie4gNO#@=XSC5(I
QZY:N7E\fF0:eUeb=[M#4OW3W,a[THN:E&c:DL;3ZGTe,)](8\Wf5BYA2H(4?C/B
e_/PV5>)GbUcNXB[0U01V^2bM.JLa+,^[5Z8eE#T]c(H7WfP<M6?fcKPCL?FgVQ?
/A7MSFOdgGfBBg8^@+T7Q,He]/;O//3PIV.C13]2@_]))Q@V2Md]UJU?4fUc@/C4
ORGNG0LF1V29BOf._N6PHR-H3\<[^/a_FX4Q_5GH2+FNNM0G[=G#Q<P[Z:-,_>#0
ed-HVQPIeHOS^PUD4UQ<P\e/WJ1dcLf8dL+&5#fRg:D5G01V5&83OfBCLUGF>/T5
,2de69FM3L4g]RQ18;/cf,Tf[[EME8R@3.<)9/L6S8S8<2VAUD#^^K@,We3W0=2#
J/V8NIO)2,d-b/EZ)Q6?-?-fJ3E+T[VWX<=&AQ:)JG>?b@P+M0JUBJ\<A<Fc6a-V
WW^e,SA_LF[VG_5R5_B_F[^W(;&L4<U-&+(RO)QZ2^MZ5Na=P7E8ZMG0V0Y#1&1f
]f0&Z4Q?=6e0XFb.PH4T<?=_He9CB5.^c[)Ng,?TCXWUOV?LGc?^1gXZ]2PLR]N0
<TdVD?P&a;cc[d;N&gU@0c=(WHDf8N2+][X\:J&:I(IV8[[1J.UaJ3_F(RT=@@D>
\@WY3@K-9NYQB6HN?-O9UB@),A+#(O5QT2MOf6OY,aU(\A<2_IL7&THRP/7bWaW5
fYEJU&[?1:X+14]PUM25H?<R:RM8_+^,&W^O#A7N4@&QRV?#@Te>YN+JO_#WW(]P
FCJfC9:?_-J9B]4)-a<:>B-7B,N-))OI\?3P<gQOT9;:QDC<[LaI8-^-RW16;EIU
X_GS?XBH0@?+?,9?/&]P[;7/7O44L,97b9@SV(a91e-Rgg@&DCQ,e8cgd5E7AZT4
.Hd0dURXM16EW+R&1H@Yg?Wd-0Q4]a63gg.#V,@c;;c5_3]K5Ea)2MGBH;JR-&6>
Y-,b4\@\Y8H-D0,<)4N@..[5KbY,;]gBKK/?Fce(fI8)@c9e?Uc(+W9CVG9_W)M7
bEG.8V]4M7F3O4>VI:4IAe[GT(+.Xe6;4K]T>M:D)cIGZ7I;H2]?^^^DBFA/+33X
WKLYI-]P04W^^6@==fL>C_13&3@Q)\QB@YfSIQ>US+UH<C<b3W@(e@>A,+9=d;#g
?;,bDM/c/1=EE7Y6:#FKX#(LR<WPYU]cF8@gMG2#EgRCDD53X(f.6c+&.5LKI;]\
I_(QaTcM0@JP0D24>.eU:EB<R]J66(0Ka12R)^)ATTefGb0<U^LZWc=HJ1-a)f^W
f.<D&:G(FWEX.Y54,X>e5QR34A08JbL//27+016g29;4E2:]2FRCeSC6=M:bO]5B
IacWYOI.<[fXRJE=G;Va+@F,fF_7dWOdfV9KJ0c13OMZ-2.?dYI:8O)8Ib_f=)E;
Sc.9]7,/.gfcCCD8?5&FIQ;0#B&[ScFUNN2Q)Y#1b-aO-S#S^A).bd+ZJ4J\bHI_
GM.1,UbQ-R0:29D@?7Va#_KV3)U#-YPV:A<,\&c?=MU3)\-.35<e-e?#^E^=;G/X
S#1@F);VW]29&#(Z3?KaN#UJ;TGU+2U;4[TS1,b21D976,6FK(2g=QC3VYYPNU^6
O&6SK+Z(ee0-]IV4-MC9Y8,RX)S-^C+[3S^_&7#/I^A[0Mg+0e-)c(^6#>#:OAM8
G)DP;J[QRNSD6b_^:=gefRW<>e;dc]YJ^<:2(Ec#@Oa);?4TT9_L37R?^4BN4Z_W
16H@5.(cM+cf;)+eMB[/I[IY^6)#3dQ7.0gc@^K@=ETP)WF<P@\]3--O3g7P\6/4
:?&S(I.g=d4#6c55UNfQ^=A@1]9C_<GAef-g\c^\3aGQFaK>0Oc16JRDWP8dN<Y;
-AI)6=Y>0^<41.:8b<&4_+VZ94fQ+>3?S:7APB=1ZN8a4F<:A2=aNW8eI:8I(K,B
VH.YPf0Tbe37TS_/9b^2dBMRC5L3P_69U?_\.<VO^[\OWc_Q>O>#JPd0eDP7Rd\F
+9TZ_;@7V4S++e)ZHBf,L.gS:YEE#;H1Q2Ff1YXeCLg#MX6,^)XcG=?5#2gZ+I),
M;89N\.efa1VR1FXB/K83=C6.7Fb;@NUgS&K]LW6_S=dG]]^4<68150+c=d&SC]F
b53F8LI[/9UA:d59?PGA]2S8@fd4DKd:@#W05B_8HP)J^6BG7b)?5Xe?&-U,N,ER
#ST+F?#Qc[:6WUXA9fU9dB.(BOF./,K7J25gPRX_3^ZdS_Ig34/H[[&ZgfU?#JF[
ZJ,4/XGX),0W^9]#_QJC\)NdA7@_a#[&BD6HC=9T-+WI/dHND?fLBON&@#f<\K/?
bX-;]2EL&#ZC&__\N.NI0KNV?;Cd_HDP2OG(L)HX_cTK88/fHM96XI&f8fK,^A(g
E8/O3U+\K8+WT94:W@1TcW_H]N2U_\9SMb:J5;?;8Od_]f5>/X\PSaTO_cZYC_F1
[J_G\,dK#&+SY(T_XS^R&54PWG8/3LJ>N_Y51B9.0O4Ig^Z>d0QVFOXLDJ922_O-
O&NfeHUO#b:L>1BA1GI3?UAHC4,L[@If?bCC:B:\T2U#/(0X6?J&=/+@;4<R-IP)
#MF(L6U>#XZF7LS:]-ED0d93NG?c-c-@+b@DM+-ERE@>c@X<QDIE6HSd^G[2QS71
S)ZEDI3/GJ4PSA]bDGQ@;[8K[WM9^,;57D]^b17,IA7B1.V&O\EVYKbJHYJ?CS(G
Jfgd4f0GEY8D1ZJ6>_G8gY5d1_,fdg^T_->)=\,E&1>A00K_N^2D-b(MC@Wf+2DU
g4^)OVW.]PGg]=Sff_<.93(F9D/5Kf3N^g&S.)?]Y>L=X4+4.e=f\T/SX>\[Q<<8
]YDPVaR&H^;FUaBOb24RV#2>+RWb7T-e8-YA8Z53@?\\Og;&]6W,&E32EMDC3Y53
8+64];fW)0\ZU7(DUc/YNLbJS6#Kd()T.VZRAI4XCBCH\,3:K,#A#?6V_^eAfZ?d
\VFF:eJ@]&6Sf(YG5^=^]J?WeLQP]4.F3T6TNQM18.D&g3F+K/69a.VEH[2.FbNL
gUFbYgNdUMX/=S\ScQbM<:SEDIIfT(MB_<5YgTU<GN],:-N/.:@6#66>-5MLNGV+
@N>028N\6=8&\FWIAc>RTDX[cM.F=Y[F+7cKe^WUS4CKAe9;E^.),^eCd73;Q<?I
[C7\1T+Dd>ZQf4A9,IRVUGD0PO@UJ]^F\bT\d6?U>@2R]Ue#47?V[TbWg1AZN.YC
#6FN2g1cGOK2dESJOO.S#6#RO71O5,g_4@GYL./eeN\<;NS#A/5#=:_VWVZ?Z?,W
;VP]^PKLH0a9J,_N9YN:5?b_FB]6ad?X[RW6N5e5(@S/F(g26?MYf<Z7Ld2dUB.2
PEQE.28H_9Y4_bXYQ>JdI#6UAdPK#b@)WCT^gA0\^DL<cR,OVKV:6X93]:O83/?,
.PHb?1a4d[B_+>6S3-D<FT[?QQ=<0<E5-N;6^9\K^PW\:FX_B&d).Td9^Q6bJXFD
dEBWg5/;b#1Y8WQ0>3[ZX2LCaZMDbA;QS@)cLE43_;SH.a46+DO[4M_K3FV2UHIc
L8]bS9?\^dB>P1TI+5DE]+J6MY=_<(9^PZM;FY^QU+Gc<EV6EJb_LEYXfWGG9;Qg
#.U[-Rc;R/d6LJW+M[@[U1\.DC;2JcUT+[^UDA(\-a(98+.d:S>eFY)8b)L/+YB/
??;0e8H[)B0)gJ_\K#KY/T\Q[Ta;C3X1J9#dN/Z8G3A7(af.8:N#0>JbT)?&(-+Y
STLOCK)3eO/IJCUWZ<B?67aM6[fF?FL@_6#fO4D5U)JERDCcHT)@G(_:_FQT\d(3
X[T^SdW.N7+QDUN1>94][cHbG<Z47(&f]#I&0C_]WJ877V79912RO?W<@<J5bS:<
)<SR;fG]Of?97281>C,^2,b=7g.)7-F#_-R2P2-6gJ70;S>7YLUbA.J0&486Tc-V
@fKE4X(WWf0/]fF&V9\,E1Nd5,N<_LT^399SA_^X5f+9&(JGC,)R\>U)<e8@BbEB
=4U(d&<:??Hf9[X\B?XL.g3#I4KIWCXg:\;()U=-BHDQB-OJ=DdV&_X>C_ES&E,@
fZ^F_F.E2<gMVWWgX2F[._27Y@UJUT8H]<#D^-U#<SWW2I#b@Z7,G,\^aN0-HWTW
>aS:Q5beCYc0.\IJW[2edVL_6b^.:1A1a4J@QE3a]g4;;W@>SAW\TBVFNS#+R\<&
^.7P8TX\3I/FBIC_2+@AcGMYPQQbAMW3Q2&3(T8_K7=9/SC\0.BEc))R8&B8N:41
&E?/R76PQ:](@J&b\gcD,Z(e5)DYPJfc\]WaQ#L_>BYPFI(dH9=@NX?0UENRZ88e
N.<65cW_4H-Mc1,2+CW&=XR1=LVSOWUZWcf/e8DGC[W)MN-O]7Z.:)]OU/_7_QZ;
LP34=.]]3I)P?38399A2U.K_K^cB\.65C;>S>J2NIACeC=7[eG5+<P,&M^2;/5RC
X1A=^f4?1&G+P?GSVRF]35Be(H4QW^TY6I\.QH@&:,@Pf(f)c=[)1&;O2bZA8<Yd
Oe8g?OG_I<M.>B/78D33X99eQ2D-NGTeL,OS955?]>g=d1&_dZ<#9(O@PR#/&9&H
S:NGN4f6V>Z0c+ZdTG1c9cI:-7US(+^fA]FB\HT\cY^#=DKN1HeDd-_Q8O=,+P[W
NC:]VK.G(+]^7>GSTKQYd@ZXdWg,fWZO>)FHHD(M=IC0M:AM8A\QdQNA8N7RZNUJ
ADS7Q8OZ(OR)XGKR#.O\93a#]1^T-IT+6(?G;0BS+QPU&:NBVQ0JA2AfY&H31O3Y
8XC/A)6:21)bdgP;4EG4=eDdW+P,ACQT@T-/5f[)(2<NPOPb/G>054MO6?(]S^+B
3gR_&NJRL5K..Mb->C<LXJ5c+7GHZC14_.4))8[&9;91YKO0b)I1A_W<WQ_J\dUP
KT]_1ZY1:DaE9gWQd>2-3HD^UDN[H-IfPH+\6&O\cT8;@4eH\L;NY:)W^[]S&&:A
fIeJLb@0BXO7X>]_)?YS+FTPIKX74-c8Y4GB[Q&WZPJa]bB1DC+dNgb.e3<\R2/#
UI#R_d\OQ2G:(?>)J]=[<JJJ>_=;<OfOD@=dbN#&YO;?2#-_N3J;/ObS3PK/QTW6
Se#+[P#P,<LAHU=4gY&\_=>AC=XeYW7]6W.?A(Kg+Hg7&E+8#GSgE<PdgS90V/#Y
[:7a2]H,1VCS^77aH@DA?5CXB(M&45YX(&3gS/QD^)6Z\HCKRc&7.WNK^0MDHMD.
5NSHUR;ZTW)CH<[aR7MKf-eXKQI]M(=Ie6U9>4J\6Y;M9d_1EVSA,QPgQcP,R6+G
5W/JK^c(OI.c-fdZ7Y+&KLG2+cH-K=2GNHOK5LD2BA8O/DC>\+gQ-IAW(MUA.TJe
V>X28T):7UF=VO\+3-3)@FTe(S+)Cc6(V<+RM5CO?A+ZIg-TNC+GEOLA981ZIBW7
T48HFI6Q,a^^=\[b=)F1Y=V3>5eMbY4<]L<0U-)c-].BHZI)I=VU3G]3Hb:5HC/P
8,@].SEFT.30bWTZ_@>^QB8a6PLWPL^N6+]4eG)4PD3EO=g.fB+a=@4F2@]MbIDZ
_)3]E+Bd=^2ET6]U#0-5YI[a@Q[Z-_QU-=J)0-TM[=,45SR_)JEaK52&FDNTfXEC
dGI.NC2af\62CDS[B[gMX>.ACI;H_A#QERWZ=XNTXH+af4B9C_3;:.:;4BI0c][+
Y#;?0d79ZZ<.+=f@8K)c^cS?0[OCfb5d^F(XKaedYcQfFD]+.BDg#NVM9DTZO&J/
g+D]YY#.,Q/5X&5.JMN-a,dGX#CWPd[1&Q@ZZ/1@XET=_8SW-YHPS;(dJP.GcTB#
M)HXHFE3F<F2;@LcaAM)ZOQUNCT6Ce:<[9,5^gDI92NC.CgDCJCO0P(=&S(F29d1
cJWEQ]HSVg]F8g/Aa_AM9]NFS#(#@]FYZK@QJ_:D8_fFHd+AL2\R/S+^a,;H8[>#
+gOXC<a?1UI-1a2/&@2C,;J2gabg_[HUX_DJ6HTK-ca6c[Ff(L\&L<f&US(Yac1O
If,M2:aAe#PR@L#9Z0Zd.\&\,,7(TbF>NXO.Mg<gV@aXJ@5XcfE/U8@c>?(@2cOc
GQ2S_Rgb_6M77ESPG7b]M&VY_OMXa6<^=YRN_P956&CRMd3b/aHc8:H:MIV?;QE1
>Nf\cecAU.#,K_<3QIf,165,H[-fVZNIUS-J91^ZZAYMU,BEB0cLISSI+MBH;DQ^
/gIF]T^9M1<B0YL)QEF#Ja/Of)+E2=)GJ3c&?VKS#Oa_bZ(;f(QSc[E64O)6+C<)
^-WHU,XN8QAGHb[3f.f/TA0;3G9J+EHQf0Q,ZH[[PKOg<<+:+I4A(@&[)AB,eOPK
>=SbA.1\B9=&#_FU/.M=9B5J02&N0Y35@33B?_J)Cd\N37&QE3dB3#?.VZSKA2V5
[@D+W\J^TL>d+1dZ=PRWB)ea^>U?W7HRf(J/>2PV:g3BT.3c<0/DLLC+e=)dJ86#
-AL]YGJDD396XdVdb;>C0.ZT1cK/6HQYQ26RVDOS+-J(3NF894Bb>]3_g;5<)N71
/,BP3_4#=/c3QB=A]Y-\GE/6CC<I^gde?&#f;4QW]62^=GAU5/W\?)0c>gBXNHQG
;8Z7Y9ETJ&KMH2?@J]JHB<I;c57;:;N,WAP7V=18DA]KBN2AL-O/gJ^N#dcSJ\gP
ZE>Z-KQ42O7-ZD@B-2H9e;c]7K-,3K;;0<?f6B4N8fV5#LWPGXW;e(B@=;b9^ffO
M03Q_G6E.+YRI&6Q\-\;#A.BfQ_.TK7R0Pc]VbQE1BdR@F0[5]KHOe-e5=#aF+2T
K0C,@-Z2R43^a0[RK0+a?N4U@:WLXH_D/\W>f7W;dBfJ-Id_@]626G7^J@:gDf6;
7\f&SJD@4J_HcO2&)ACG^@60X/_b+40eHPC3A:V6U:2;2g821NS812-23.1+\[==
cM8?]e9:_dD#=:^IOb1[2D?(SgP;)UED/-ZMZ<L@UM-WMOML\DIeQ\=E1C7&J\IL
?=gaI6+9dS>O=gH[KQP[CeVCb9?=V=5(6;dO8#IO#6H18G/1?CP:T#6IYU/UY)N,
=,:A/.6[Bgc]246a[Pa;S-K7<=\YfeLL3BH#H90K)#0;DQ#2YeWJ+?ENQBE,T[<T
VZ@F^)OMeY.4H4/O8X]c9=Q^641/<P(ALU2B>B>-\@^3/S?c1N]T7;#9-eA9V0+,
b9NVF163]A;4Cb2^1+M+FSeIFg.@&e(GZ.db(=1LZZ@O3.-[_/:M-OL@eJO2c?P4
d.NH\:,9+,R[NNSDR?dKN->3V[eEEFGG0A,ZOYca\><+(6GAaQ=Q.<gK#+-_0-;5
fQ^>0c7/P7Q\W@=g;84T:d&a.B[=MCGBJR5JKS0)EN,ZCV?LV;9AZTB+<@8We<6.
4N4<U#A)WL;D-7PdO0S7VFTB-M&<bId[GHQP+[IA\,S=6W#ZKA=dB<a/MHAAZ)UJ
.E)&I4BR=)=VgbF2L8K@,-AR..\()OHK?;]<^M=aS.EOVOSXI<55HY.>-a5-SWS?
IQLc/R(XPB.IM9E:NH#MCJAM1.c8cO9[Ab0ILfb&ZW.#<UHKCF(/=4EY(@bc0LIe
N4>3AP1W>@<+;VfGLd>/CVW83.QcYY50<=#6UVY0c0M,c5cU#+:Yf@IeU97-<G]d
B5QCU@5@d,X2b5faU7W76M7g&\=@72]SNQ>)\H+EUE:1E?]G.Nc/FE5g8]<JC]&^
]Db:QH\T_Hf)eL#4ZJ:ea;B6]>::c/PK1C>CQ]</A8b_Q3H+/&U)]UU)P9&dMbC#
O,5S1YRAQYc=]5#@Y@<8R>/54O@:KF3VEbWT^9aA)[Z(XTf,NP.[O?6VY1Tc1MK9
87M(64d@gT)5Eg:ceD2IMgPC>L?)5_c@,8KXC=RR6f12cXDS&M7^TK6]Q7\Y15YC
FZ7^:NJ<^O1:8?1/3fEO\^14EU2g[eLd0fOJA_FGO-B((]@@EP[ZYBBKP5EAG#VG
+,a(;V_?S:=MG\d+=MW__H1ANIQP[OJcS0?&A<?Kd49R.UC0T2gAPFXX^Xg3+fWT
P7dJD&-dY(S=-00?T??UP3Bf?=Qc?(5-8K6&^[&,-#ZSYIb0.>>(2_,WM_[OH)R>
Z)?@ULT?B@cB#2EY.CV92LSXBb:d<cZGAIc^#I+I2fG6eGTF1dVcMEa)B4)P>;?6
=6G=)8,VWeLPg&MdcYP/WCE&Ba+_Y9f&TM9;D[AR.L_OMG-ADMT5b+U)UXG1@WQU
+V2BK>g&Qcc4I<0NTDe?WcBQQQCYJ(1XMd\8LC,W9\M?EC=Rg/bVbHN7f.;>F5?C
EUG4R>B\,e8LcS=#=F0c\O<OX<+H+8WQ2Lb=M7aZG9NVK=\E\,_0D]WfU)J]NF=S
9UK<cKL[>S]72&A295]AB;\fPUQf()X;Q=X8.BJQX2@RAe_G1HZO35DP)TVR3[:L
A])>ZWeIL-+PcA08JF#UO+W^G6.KZG);><QGO,eO<FO&.e]5@]X.C/;H>Ef-#WC\
D+4,,b2)A/N/EU-YU9..DCgMAJKd\7I(8Y8.5BE_/_W4(:9cP.Dg;3<2K1+b\Q(V
eCdTQLB&91P=E7-CTBJbcB>VCDP@>EER45g@OHMLYb6B0A@C\H56CGSZ\0F6^_2I
H9D<XUEQVZ\W5SM[H&_YeT_FQ7)&f=WB<QVVgaE))?>=Z2:K9e,[e?(JQCI+DN3@
,XY/1LJZgGCO5fYb57:+Fc>IM/RC3E0:G-g@PJPT(3VJE?=B0P?.&e0]4V-I9->a
eG(4?CLg^ALFA>aF^JI_O_DKDO+[3-9_C\Te/7V>RXR,&;S,F=#V1\P)A\-]FWef
d&=bDL_W0;9bc9A+_)\dM86]14T+I:eSeAS/RX,aTZc,QP,HFcVQ,YFNJe)c87.\
ICg:ZOK;M:U;]LEMS6@6WQU7H:3MNa-.;Eed00BAX43).2f_VSNe/\Ld#<@J+-&?
Z,]8O;;:-._e?=);-6_Q2>SBF52d@DeL,Z#^V=^B->5.dW^:5.B4BSE[eMMSW]H8
:PH<@a@gXIP3>7aZb6-NF9/SZWCGR<PILK3DDD(/gF=Y&U<^LK=+<914Rbg1DI_O
?Q6b/+]<CDGTbSTGP_I@SU#X=Ob2<I\1_SGV&&G)&)g]Rb#dD&8@[_TIHOCBd35Q
G)4.2CMfXG_a9LaH,+&0ZgOF4Hf)Lb\T4^,B9#Dd@H/80?PZ.5E8DD-cdQC(?R6c
Z5TH2=Ta9R]DG:2(MQ0L]4BEVD\-==<@@dGa5SbY#NdO7a(N,g]7LYLE<(/[#@EK
.d_Q.WZ2FB@1Q]J0_81-C=<aUH.\/9&@_FfJCG1McK[W8SKTO_@R-d0(FLD0<aW@
.L3:?J8I1H5K,UP>b11BP4;Zc3X5H,U&>I_CINdHeUJK]LgGe\-7KA.BGN=-eAV#
+VJ:P/@HOB0&\aOfQZ72,FW8bVGT]LYf3OA3HL\[7QM6CEXP)YSB?:CGHC&X2D/S
IE0/^;0M-4[0F4DJTcE,A0aD<g=X_VPd8H\e\EE;LNS@UIeZZZPA>XV3>D>=;4.&
(/+Lc72GfC[:?L^e5&KOM63aW@M6-MM0G(bF\RP><-/<(4<g>1D7B8FEBVg_<E6E
RS-4Ld3N)OWD+gMe[C/]1:0+4=1bJ:]c<Q_&((f4&f/cNgg#0=G9YBE<S.;3/Cb1
+bOFUEWKGB1?XEQAeA4.Qa&2aQ[SE-:gP#.>QBABM6X2=_D7_e.IbZ+^8QRgL?8>
:YWGV)6R4OO^A2[^?eSI#MUfbKL?;>7S9T?G=0LPZ=f7YIAcbd\P;G=(C9=c/>Q^
#D,A99LV2??9HF>8JU/?BB5)f8OS8&54-eHe&QKdBA<Of3+WSX19D@4L8dFNKE_W
B;.;R^Zg7GW.6(9B?ZHJA#_M<g0Y,@YNYNVDAcABa@Me5&O)ZAHJX-H(CD.34M),
b^Q:J@JOV>40JX^IeAf[9-2N/22PIAOBA3<G/@MggLR#_Q[XVVI@LDR0UTM+N>Re
H6SJFeYX#UEB0K>2VCT(f^\-<?#<C.UH6]1/]NYcWcPP(.D3>Ib])E;7VZd3(DPR
8/-#8HU_&dD3\R/285d<SIGa8^W=aA(77fUM)G>#D=#7-5aLWI^:/WgXTXTXI_7P
5OKQJb5VGc-I\.7g5cDGLA3>69B:EGKHHBE0]MIMEAB,_&[d&7,TQLg8+Ie?=/b_
YU=)/:O]MUF7Y?5#O)-eYU;FQ#T;QA8_:YL820dE7D3?ggJLCH/>9\>\5Y.b<:[[
)PQK_E<gS9;7S+:XADe/gEJ_1FRTG6.1H8O2(dXX/VgeXcE2#gd)I58I6g<_0VN?
-50&Mg?T,<UH8(#/E6,<(S0YY6db4;+C?cf3(Ee4G@e_4=U:A5_]<,/&[.,a.>)J
b0SM2<f3M1=J:^+3\cYH-9-P7\Y+:&&eESIbNKI>K3NK@g-.Z@OZXBR[M)9cU.5c
f=J+VgJ8&.f/.AY)JJ,9Lg0@PK/S2f@M-WSYg,0M0>&#YU?PY@BSaKX8OP9;ZCNb
SMN0<?0I4aL0YfC71H:?]cR>G?.\39P\(-]6HYJ;X693@McHLY+KOGN7W:RR@)\M
44ZNK7I<9;/L9MZPK)T]<:/HedYReKLgSNULL;e,9eAa5P5).[f@_a5@dE4E=GGb
2Ff.231O=.6E6^AES>bX&T?()PJQ4?_7319>D/AC0664AF^6PV&K+TM416,(6X78
M^b5g2GW/7;>HaN:7e(+c86DH=,N\)GBS(787S4ZV#0@^F-_Ad+^7?9I\QPQ=</.
?N2^2#J@VYafd,]_8\TK?9()O1c8UcR)Q4:MJUYa]F,IGR1/\F5(7:8#4/,<R-#f
gV6FZ8eY44.PF>)<TWP6T?IfZ-PdT<>T6<S(S35JU>2X8EDb<;/P_-1W+7eNE.d_
35NB2NM<]WNeR?Y93c/@EcJOeZdfH4eF^b#+I@7ScfUd4#SSI[&_MO&&7#gAa_BE
6H0DJ\R/GGKO[f81-JWeeU^7XWA7,II,)2_]CQD#R.c@gPZ63X_IJDYI-OUGR8MM
4#UGgKfL#/4b?1?&<Gf>aMbCM2:F3Z(Y^[)-,7IN_:gb;_U7_=+3>UU.VQB@A64G
eMB<6P(@<BL-^3Lg3C:QPc,\?@;4(EG^9Cd&4#<YB-#5:gIQ/TgR_O)#?BdV:1,R
H458;[2-39&J1S:61YRC\_W.CQJ<GM.bLOIDG?FO:Oc;D;aZF:RIbFO0>,WT(2;8
=I\_0A9aT.9<?a9KHD3TQ<U4:f?C&2dKUR8;f10+:YA?[GI:A,+25ZU55@/RF;L_
3a.>-5:=Kc;K.F1^^;N@57QWN3-^K1fXeS-EQ0)1]-bgSA(IgIYETJc2(69E6b@[
7=E1/+bc6F928a:2(e<>/BCEC\>a0OYb+)U:,&a,G#?)3fR[TLQOAb_7X_LR(_d2
;13Gc^)YR7I26ZJ5D1A^7eeQ@AUIKBbB&;GSRE,bS]R>-+Vc^U;_X2@8f=\R?UQB
VPbE7-A]:C,X-(dUW65:<[QcN)CJ_]K3+)\#eUb:E2g2SIZ8-.QY#5O3F([-6A98
,gU&/=+O,B)-DA5=&b4RS-T/^,aeJ8IQe46RW2H[HgeDACYTMZQ:1S+E75cgGdU\
.\G4YGC>e?eg&[XYY/^+I1J88B>FcB&OY&cE]3U&M;>F/VP4(B.1)Z3R5gN>^OK/
<2P]dRU94J.9[=W@:f4R:ec37QYc.92W^XT8<Y?g>RQR:c<797X>>;([18E?1N]W
g>7a)(VRVXW;Q50Q1;+7YfQUJ\^I&aU>C7\@AX3H9Se=fX;94GD56M?Q=YAJ@Z+>
GIE#T8g&YagXTG:4#J[1)]U)OZ_09-0eW,X1LZe=dR9g=OK1H--LI#Z-B@<NO-A<
V-/e,XfJV.c<Cc#6KUfM<(AcPf@QYB=;U/O6[73]V&>.ITW_cAH(f=?GWE1b=J[E
M4)^e4P33K>c-O^E8d?#?L6Y9@Q\P2-5M-.9BgR?gZ]Z;_e#&b>XF)@aZ:fGCR\W
2&M0WVFG36d;+,_II&bY8Ze^LBS50RI9W:HaBR\eS]?c9K_R.R@2KeWAF573_7O@
6EM[/[B<)\GBd9Y7Y4)?_J3JI4]eK+K<4Ze@2S1LGYgQ9&A_YObK^ZY6+Q<cPYe1
O(XW:=e#7ZN\X_Jd1bUgE01E&D(^2e>\U>92K;)LHMVEd0.7GECLa]O0<=B?4Lb8
?TD&6?fEa&\;QIQY/D_g969=Kf5R__aaZfWLKV&I;(_0#6GL.B2=F+H=K@eG:CB0
OC09O>OWM&I<>^,EHeA1;GF@\?MSaVD03XG8CLP\],EPUN#YXM^c^g)MT.ZIV^_#
B:Y90P>gQbQFc]SM^-4((e6?Qb=.2BX/Z,g9.TY@+>\P8Yc2>b)](eV:;6Q7:)]f
5BA=IJaJ&N&F4_gM#[_(CgSY[6W-dF/2&QCS1ff>CU[L;81R#f3MADB.5FD7UG1_
/d.b&f,F]QC&S,HWLLPVd8C1R3IRaJCecZ&.cQ6GG?(I^<R[_HX.0:gWJ1FAZ.gJ
)F,c,@7MI_(HR4@KEB]-S72^bU[2LNL)<PL[6aAIVB2/R-.:?S#VM.aFeO=.APd6
?J2TR+;SZ3TTABbUWU.eVAfANN:eSM,\KHFT+I-ZD>HSgN_XJMg@=Y]NGC,fBRBU
X.9&ffI=g?RS(L,Q@]dL8;e+#[1MGC)MN8d<RT1CBE:[7&.+N@2?(>PSI=U=?>,P
P5g;5TYA4eH\_EQ0?(,)]4)QC],.A<]GJ4W.4O3]<:-dECe/8)VF5OMD<_g.TSVV
UNWY?2NP/AZ<D/]PPX#)M41SPCYP@L1_Kc#31gL2X_fGLMZV+\9>AB#9daO:b])H
>(1S=3CIH,.1BIA_N1JSA9<0#gO/(ULE-c6Sg2OgM<)-I7FU_gY_-H\7X>E:9^1,
HX?P?X?2.eN6H5Beg-?8,aP^VT:(1G[b8)XK)4P6BQGQ#HB&:3<.+L[Nc@b=#(=G
:3#.^aH[I_2.33.((XRV@H5B@7;VXb^&ZFPF9E[#&ZPR5@A+K(@;d,<<=CTHXWC(
O;61cFZ+g(Ec>^aA<)&@SINNfc9S2_9a@(]B#7.6\:8cB1T/QV^eAM6aOJ@I;?@c
&cP_gEe&23cBJg7PS-Sd/FSTE0S.9e38]<Xf:TH5c_7VPQ[=M]3XR5?9@9]=5eYU
GT&J6ee/SN9_&e^Y9]T#D@>^QDd,L>XL)<9(D+?TgPPC#&]UG58d_T@RPIJO+:X>
Ob[2?.UZ>Y4IP3@;-G#I+VY:b(3Q;(aU7_IXDV&&?683M.S)+D7[BaVUD.E7U.=a
8HO;E^ZLPLK&E,LQO95_K5PPT5MXMBL-N><G#-cD(a#P([XU_AN;P8a<27+(-]ZX
#IUfg3)bTNATS/?6;K0>VS)cL.aNF#/3.@.WR#=e_cNE(J[@HeC9gW]C[IKc473B
+NQ=>#L/>JWLgH^c_d-@<<B6F.TX^MND?:T:2&I)\]g7/TBF78\=\;#7^Cd/P)c=
3C;PC;LFY,S0T^=dNZAL7Yf(5Y.IYN8)_Z_@U&T5I37b2/&K\Nf2GB+V_K_6OTQ.
M/6eM[+N7-0JI1de=OQP0c_+N437N]J/@X^<6cP)UU;/Z=K/1eS5YX>Y;B]F;R6^
Hac;H@(](?VCO>fbWY9N[HE4+Q(,^@)TCXdc>_L#4R<eUdU/N&UC@9?BHKWKb&&@
.Qf]Y6#ZWdSQ6+F6RR[PR#Y^:??;A.V.Ud+d7&;4?62E;]U:[9LPOIASgC>3b>K<
I&fR2QQM?6MY7)0NON(.0?EfIIb]M^(YZ5WgIF6)FHA?7S\V8)Z6^38.#SKa2QZI
E5M<c/:IP<(/V/]P+#JYDJ8:aKDH\KUaCdRgKD[)b8-0dHVeCP8:)JCgAE0CBbIT
I)L3UN)LP9;bOTKPAXd8ITcdO5:e5X+M#e-8?09G3-a9RdCD[E?d6>N=[JHY@X>A
^2^BNM60Y@2N(/>T-,1^4d\Dc#0]TDcD-4EfRC>QBIZ<7V#LD0@X#W])N8EK/-IK
<Hc@)ZZG_YO:E[]a02=Mb7J1d\CeVYJf:I?][a2GQ_Y&L9,X=d^HIGC=dL^Wf#7.
ffN<;EQVS[Pd<Sb6O#)=RfOZ\/JZ>,ga#OcB-ZR6;f1g.K7L7^_6ZMM^+Y8+L2EW
U42c90_J2VNLD7P2K.dKc[EVRYUNTVC#;@#O[Z=,?CL6RC6\85dVOZQL7E>^D#S4
IEb\19<S?:VV=N[P-1+&K:f#Ug,RO4_)UJG8E>0MUHBKdJDUK27N5UdK-FBN?E+5
ZCe9AaQ(3FW+cU7N_I1bEeD+#@G-RH(.cQB3:e(M<5+AAY&22&a[O+(^8g.TWO5)
N+Wg2c6;4SdFFe&_+CQe(CaA2^+6Lc85Qb>QOMJ_\N\0YOOGMSV:U6b#KVa66GY0
7H2L#6@R]8UG,EUVN-Hg.PIe(T(bFR2(/4.>]2_^=J(FPG0f_O#;IbUF5/cSCV<N
.4MN>5:3fF4bUdABCb<;:\#G=IVHQ9450YD=K+MEGD)LW,J(:SZ51LVJJ&\+\?SZ
M8b)Je)J.a^+7]W?NbQ.?SB#)c9)5:(+6,;V/d[J2P)U]1_A?,I]HIH0+f(CbR8?
^gL@#>g?ZG>3OR^2R16-V]21\1c67IGKY#D,5K7Mc00Pcf,X0gP<;GZ88dI=ZbMD
1\E&e1,^I@R9g6e9/a)-dQ)H=2g@QEdJT+9H^DW:[gc)2I,.>fX)Hd(?\YIT(B,7
W(FD=\#70M3^E)\VBM#e4dXJ?DC+<7#eN^DaPYHT/a)X9?eYR4A[<97_/5WDJP06
6YDN]3K)KLT.#XdY=3_)YVB)<03gR;g=HXW5T6CSPa(Bd.9I2Qa_R7+eJ-;KG:V(
6]+WAD)&AT<A\0Q=(Od:;VG8R^eR0C&=gU;EHI0U<Vd:W\e-H#N@2(B^g:B\,HL<
NBLZ^KGdS;IA(&8ID/(X#LK)DF83DZ;fTa(?<<A41^RN5,]=B=Kbf5bGJ/3VDX,^
+YMS7/,85:fU6aF0LQP?G,-J?ODZ6Ne#gA&,0^OVOCR5^M;(<;>)\O\=bX4U;N7S
(B\2aA\e\g2>LHUNSQ)AV6e563L=2]Y=R:KK,NM39T\g(fab(cUA3W2e]1>g>;K/
>@UYc3^E?W/8_aS^.cNg[;,-@Z12<^S@a?#5T(d,]I]4g5/>9W_f,c+4WN=#9bb9
[;MI4Wd/bc,)0Sbc)&@VSY#;0dLBF/b2-9<(_f?\OOD^<:S\Q78eFC?UCV1^bgJc
Q&1W;IPFW7fESa8Y2[Z>A@&1N>-2O>&6+._U=b#ES.^FLBC/U^F00,.<W1FZL:)Q
#825ZH9)5-D31WSGJ,40RPE8EQW:104YIYNaLSd_P^T;>Q+M^2cg66CV0\)UXNRY
FY,;P+cbZabd@K3HQ?.0UIU9e.bIRPPHTb36UKTTbcQ,4@&b,SOTICU;W@WX>NC5
JZPF>ZLKD=+=:C_(UYe,)-0B##I6C9#8#_NRIWe:+9UggIbMN,b458b(d\ORf[T@
\2)T5C/8+WeKY=8:XDEK(a::L]NLL61?a&M](4-6MXMOD.IX02O-2e1#P&MTF03#
C40S53=R@UAK(9FMf78-?9.EU,[f/MM7;,F1NWLVBdNUN#8B#gYX(Q^[5&&Zd5Y]
WX-)Z-)K\cfOacJaY7<A-MO?B8,D;X&a<V]MS(a&0M^4[9dNXHbTM43e;)-=-5,#
dA&=PcLVO]c8ZEgWWMPXN1CCB79PRbI2,/EA?9Kd:X;CT#??8Vec59KF+Z&I2HJI
C;Mc7a74c.@YQY\A).;N2X0T\Wf3f^(#EEO/YI(2V):eP4PNMKS+BJ@><;MWfTH2
QGSCfK.Q/:+S4RJF<M/,G>SQ)1AGL_6G4@_A[.?3P7T@5KE_GI;;^=42C\SG,T#.
]4LP[BPc\<6DM1P?N_W7e>E0.NcF5(:+7]>N0_308,MQ4<<I,Z7[F.2C^.JUG7K?
:-><2H?)f;9Qf7?;ESSa?=WX,=VEZ5+>]7,QB:A([U>27&e#\b&M=Y67cPKBW4WO
XPJ5+)ACDP;S<c,6,(9b&X@D5Sd=BSDeRESKcRa2P:1A0;KPGU8?(@&aEEW]C>44
UPDb,\CLV[KO0SbIJ?(dOe9Qf-0FZ>BJHD>GGZDcT7,7F^C@E)(JYOWC_AXM/AAc
UZ,]7<N442dVD\^0^-D=,_[9IHDgZ.HdSXI+X:5D:0=#JPg7H>J=c4J7]L/^/-],
\B@76H_)1FcMT+2Q-YIMf/A7IVeOR+M&e_I_@MdFLaSKgY7C<^SDL8C[8]_>C.37
J^6V>()]WXbL&G@L30;WZNc>Z5M^N/9W@;#:TEJ]gA#PbPbI^aLHN3Y>PD_AdF6Z
P3OVM?g48HP3g.bO_7#],b&fI+VNU]PIEa6A6UW7H?1&GNEZWO1V@OPTHIfVgXe+
2TSK)ZRZ#>-\BG##7]+YX5DL>=bWY++8YBbO)0E]P/&R>\)S^d9]1Z]K]8R>7L\:
/(69:\Zc:QJ^@.cR#7ZYOT#E8<PC6OMN;Z_e[J<NJYPe70f2\.G6ecU<(9AQV;[9
92\IF;5<))e<6MR5@Y=;SP4RJ.V<_K@&]5]M;<]2<[NXDIQA5/V7A;R68^E@Gb(1
T+PWGC1,0P#&H^U2B9?.AJ,/(F3/9fD6<RSXd=fKW,X\6:C-E+I[[AHCbcS@5B1T
Z3g+#Q-NE7V_e#c^61./e;Z],&cAK&SZgX]DVA[)3dT(5D77f#gDFCR?&])SJAIK
LXY]KADb7./_f4fd1C6GF^7d\+BH[.4,N<(aGAb7/+C&XUdTUXbVD3/DS0&^-UWg
:+H/])bF2Oee7)#BA>]GT=4B2ReOB^bWK&O:?NSF8.Qe;5;3H4QOPKXJKDM^8T.8
QSI=1]LT@2IN&[WMBX2d=0bW0a(/b>VUbF=Z1:aXOOd=L>/;4D6Uc?WKSaVH(.Yc
BA>[_AK35P]]UAf2?AG_ONGOb3AX]9I8\Y875eH=3J<I;HD&Ke2?VRJd#YA8(-4+
8O#-\.O45d.Qa2-Ic.[A@@Z#X#^5JGNde/A6^6TH@6.#J9F7O)-O20aa8_0FHVeW
GZ?[ObL^g)./T3N+Q<02,[NICADCEXPNII8H6<HYQL,[fFU:1VYd4,<?X?8IJ[cL
CME#?<9[]cRJ9[36NWP(6FUO4cG#D4V_00^QD>U/=0OMT\Z;a.2&(1BYWKUF5@fE
&VOGWa=3SQ7DR+F^M.&944?gF:,d2)b&8=MW6cY,L]<V_5af+HVf+7:.&[G]9V^>
NbXV,<1+[J@,\\@)T8eD+^K9^&.DM>JBeBVGA5\.gNe67-W&/AZE8Z87I6eSG2=_
ZHB4JVD?H<Bb[_5f3&+aWCTW2NM@D^YP8NM;D5]AaSS<F(D(0Y4CFDDMEX6X.II]
UD1KFP@\IJ^;d4>N+Y?CV7+g[RL_DM][SP5_UEBC\]Kc.QS#]BJ;T_BN=LbE5P3]
D1^RY;fR(cY,C]3FfGK7VR5>^H7T,FU5>FZ9T7IPWA)\F\X,#f9GJ=4QTa054.UQ
74CZN_W0MGb==;B;^1?V3]8I;3PRAU1V\^>NE3e7gd/RIEcODLa._aZgP(MPK8(&
R0@cB(RF;9dY)+Ib>B2(c?&LH^01d?&e#@f.b&C9HXMeS&J2D+SE#,,#5,>GF_SB
g+-&KB/8V-LaKWL#0@9,=^^>5A^A)R^,@M;>A_;VU2YV20S<c)\LC@-L4K=3[bS6
=C#MQG>aN.D>:T#2>Y&J1<EYF?=GSA)2cPM(:b#Z@])-GCfZ(c7aG&bE,8LB;/_Z
^MGF>N<5.;\K10YR[:[[Xg#^L=C&]NSX,MHHeNdBJ0N]7M9+bWDU2EPeV#L;KUJU
b:_)Od;F)G9#eU;+g3:9VHcU=R5??LF42>aIcc,^FQ8fC8<=#F7W>D?d7a;^2Z#,
?]L3_#5?Q;[5GgU863LJ2W[2/6A=>Wcb70TfM&b0_,&4aaJGbQgM6DE]NP<9;&/3
//fTP#^:@7Ce8LG+7G;V-1e4+N-GKN2g]0P6GXW/I[VNES1A=f(@;DcJ_Je;HQQ4
:]D=AKF07U8J+,P/?20F2Y\Z1])/ZGNZCHF/YDL9@614>G-G<1DBAL[)TWPK^/fE
S-:V7V9ZRP,ZTL7+M5\^FHJ?X)7][&1dH,8F7=UM:<DN9]#])[]#aZ\^H22gaUJR
2V55V3\)J^OR)YJI69:;1)SJUQUYQ;de?J):g:)?^8:LcaDZOS>Z_f>-eD?bY+,J
13#e?UW,G<Sg^4WEEDN79Z5K5f?Yg1W=C&?JN^abd<;5@(2T8?gXS<>VQ_ZY)76F
<d>)_Q6O];?JT)aac&NR<;VP<d\>YA3?&R^51])=C6f=B>JRA4/Kd[EC.f\RU6eF
LG?J4V@3FdWK5K?_SON3.gFDQ=d@Va)&Z7RSXUDGCAB4+(VRW/R1T#cACYcL>LG>
QSCUa0MT2^F9OHWX+9P[K3a[#8dH7;TMg>Z8HIB#AME,U?.1aGQ#cJZ7WbaT_]17
]152P?QJ[D]>17UGR]U@B<J\#GZ06C#aV9[U0YBI#:O-+b^_>8H7:XH14=MX7&?Z
;dH4)C3+]Q0)-+=;#IUW,eePa2#>[_+0V^E&K0_.aBMZS9SPS\?LDFXJK/@KR00g
dbGW_8&[)LbX;M)>>[;KP@BXJIJ7&13S;KX8HP3(YU&W+&eXc?D284Lf46=7a3(M
7Kd/4T(;++_D,/2W6LCCV_^A4BXZ?Z63&,S=JGO,RU2T9/,bC6)V>2ZUQ[g+8\c-
c0d)fQH:G)HEGU5TK@?QZ)4][33]3BLH@,06K0-6<\]:82\MGO;UL>H/NIK,_=,\
#V@b?)LJEY8AcAE&+eZU1c-L^FR872Qgg:ce[49\N>Y#Gb[F8=TDC8V=dc+g/:VF
[+13M;ZDR8,.YS9.Z6B;WIT_EF?#Egc,PM5(F@F[;#Q/[0WgTC1+5D=J0QRL[bW4
_f6?6_TZH-@QfVeg.:#4I+&Q@?W6&J<]65W1AP&aH_Y=T(]M\T6VNe]>NG8ABK(Y
F33N+E)>L-6QEaXX(&F_/<.6dI<Q9J>G2.-a=,0[;F43.P(#HfW]8B<&d=]B,NMb
A1]7OLH=R<L@QX,0BY_=BRI]He)1K(R1XOc-c_Q3e?@^X,4.,L6YAY4bGX1>3O2S
:QF27:dBKPLZcDdL?IbK9_BBCJ-8[6:E&RUgH<0(I8W#5#)M8NbF(AVP4>069>F?
KR4B3,^(@]D,+PeKG\0:d[KeVXa#RWg/U27;a&c]3BWV\75Uc<[&)=9[V3I5X(@g
3(0e>8:9].];FKMN5QS<0)4Y;+=3_A+gIN=Z6HQ>NKcOT9:YRIb6XM+d/W47eQaa
)(>I,4g)dLP2=QNC@QQeb[6,9LM/_3L?TDLZFg2c]HfbYa9@T8ZKM8BA4_LdK:7I
GJ=f7C\C?Fe-/:MRK_7YB+5b=fdOHXA+Td(\JGN-R(2e;UNO5;O7@@][2B-8d.-9
X0A/_=Q^O049UX]&-HW9&cafd;D9L/8/2@9\^>dF6L-&@B2YLf7>aJ0@.H7=/7[A
6K]b\WDb,9H;e5d9AfD.C@)DO#7ZVW=?gE-gNM:[5MEH>D<I?gZ--W(S)9XO,F<B
aEMSR.TGeBeB4?C7NUH;&Y27@Td]2_^1N@A4C5;gN(41R7]3<)7Z/]9QLINdSbd@
WI;LN03edcJef?3eJDH&.D1F<IgeSaDS+RI5C@a;3FL.gd0-Q92Hd4Q+ffe^=^RC
_IY0Q5T2a9&_^L5\XA^8QgFCMcF^B0VHYZ<&8J@^@+]KdL.>+QT2BA;R40P,+L1S
GaG;W1EQQc7=dKL@C5M7TQM#[-@2-IOL0H81N+)8G1gK[?>+MbdVG9N?-3=)DR:D
]Q841YGD9LXfR<P@E8cM[]O8H18)9;__KPD3J<IW)T?4Yb([H=2V2NNB5WU&NO\4
G[K@L9U??1bXRR&aV.,3Y=EV[Gg[=aG<JC7ILN1OFDJXO/_-Y(ALQ-=5C@M[5738
2K\/<]8:IMbOV;,AI9SJ##I0_ZF7H,EUO[(60E=<d4<N1=5=<YO@J/P,/1+ZKXFb
U5;[:CBdJ^B_;QE@5>)1+0W3I6;eL2CCgF_OUWbS\)PYbfbKGaG>]X(Y5:X4d_.:
HV)P3UE-2P./@M\)N)RKY>cQ]^V3X8WE)CQFD30)cO?74,?>VX<_ODQINaDP/H:g
QC=#.(H706a>;E]?J[4(/KcMb]N/+H]e)fB0I4:CRZF/YROb3_W(f.(,]-gEZA5)
5(C37gcC:c\_18FDHU44T]UD7[:a3Yc,_5fFaLH(7XYbB)N&6Qc<4,IR?4VGR(C2
2W=>ef4QLaDAX0ZSe4/Da9H\XP:fT^g^FY?GZN[HAW3ec9^KS:U<0XfUd/]1_7>F
O9P)dOD&?Y1+MG+S6I,.gQ2Ja-J#P?a[HU257ae)]<CS5dR-TOO?-+#b[_f?RSa?
53,7]WWA-7EeVAR7dZR(Md,)5eG,\e4W8.d=:Z<AE=S^=5=_c2GD<D7ZRLE+IS0,
5L(+UF8<.SIS_E_[#cNeZFH)P,00H(WBUTRL)[:S5VcM<bSO/c1.,2R_70NaENc=
7fD04OJf7Q(I^>#DF7GC_[c<I6H\E^9EU)F#K4A)+57.EYHJE9@a[MI/dPR/V=W;
F;+KdUdKd#1>fQ_H@;<:F;>E3Fd<S)9b)2H,:eM4?1=;GS<A.:2<Y/R-Y<AfZ8bQ
1^[JIdd/aO>b(a6D=RQ-+9.VAUC-^I^P+#4R5VGN+V_Y<]Bg]4OdNfPZf_>]0eeO
APV-HAYX[FOM(;U8Z5ff1-?g;.-g#^F=X7HA]]YV>gKC6JQ2R+39NI0W?>&^6e7g
[98BX0JWMUU[6<RZ?JU^K/WB1CP)RZg,-8-M#X96K<]-0A[^30FDI2Nf.G?Q;acA
]#@?>64a8;RH@WB<F?<f:7be3GX1NJ8X>@MN3;G)C)4@\05(;(4PH@gF\=Q,A9NM
QM&7BZbTKLACAOP?a1HW#?UgN[;3>eSdOM/#GJ_?d(<X00eC/O6(#[)VH-8b7^WO
)5_U07V:dGG2._>eDcC:@^;fg8-:#<+>9GK)V?]QJ[SB2;QIB90A[aR\5H@15^O3
>)W9]Y00.?I.7?FX+\KMC(aMgR^,.R,&OUbK-E7W<E)K;6M:QFA;.5NR#-3]d@8d
U:5F>eaQ0b2Nbb<:fbf0FR-8]<EGcLTMH0XRcC_]I0TJ;f>H2+@=OFGa;GZ+L0g>
_JH\NL?eC<2g)K,TeCHJ7ZBg_Bf.3BV(=E/ZQa4c/;6;(0QW:>MVKaS^HY47>[N[
YDH3JTHa=FbSQfBH)EeJ8XG)0&Da\XG;[U/2a88NWd8O(B7V.@gOgM_VJHD>MX1?
04,8C&-:6>AN/V/C=97Jd2-13=EZHHMfFg)(MM36#&RY5<3f^AJJF>^eGG/HS^Oc
:7cP#]S,7)I_Q&JC9e#N1#/38@#V;K\9>J,[DRDb6<MO^FMZ/)(>7)_)GRO[V1d@
H^O0N7[e-M.([SNYf+N=8Y^T\d68++5CE+HAE@OTM)#_PD5TR01;aIXFF>4O8DcK
2NKE)\Qd7Ra5gUE+aSPV:@H8RK85#_UT:TF8[RK+HeY_c]:Y_#LE3I.CM,/LC0F&
?SH55U4+>@b^3TG@4Y6fWMML0=\WfOM80A,Fd)c)0^6H.9b>La@W]1AMT/)VfH3Y
J[YM-9R874_\EbXF&SBe^X_FVc/+/\J;GDbOX=X5=TD+GRTP=QB5U7DMTZQ+L?5E
CS@GPXIaDg2UB.gJ0GO0^L+:)PWYgJ6XFNg95g.d.9YL290G2^@df#GAYGB2^]]M
3=WCF?F=O()CFd=J&/S90.;Q+W?AX2V]\AV0IF6HNKR[+(F?gMHGPS-M7PQ.3e)5
:/0ab#QgF1HT;_^CW+GW<7B\RG6_77.3;IW/9TRVS/4gGYVI[I-2Sf5)6(QI0&YR
]R8U^8S(495_I?KG#HF9FT5T<dTdD97HAdLE\)ABP-#7C:PJf3T2_HUCT]H=9TFV
&.fZb14XG>,8SYeGL7<(bUHI:1.8DX;RM[#^;[<5ZLM:dcHeQ>2gE1Q;#D^5A20W
ce^YFD]]?ba7XH1I06^ZJ1BPS5EOCHUfcE]PJLba5;?AHZ(3RSD9#_S6d:P3@.NF
-:QE,=(OV(^-7dTeQ)0.ZcW\2^5He,&BfGQHg82F?@)^aVY,63D:?HKC)P+8U:,]
2V.]YD=,GA>2<FWa<RI5Z]T-/_]Ie4WMR/F.e\A#]#G^]>_2H\6ESf]TF=206YBc
-K,GU&aWf+QcPe9QgYR=Lb@fV&bM21=P\M+EJ1T:0c7/e:N-RZ(UZO>.K=[18gN(
b5=gP-HOH5b0H7W<)CYd3#@M9>T+Tg5&_0@F[@#YQeV[CT\PO\J:]31PHAJ/P+EI
4V4,VX;M\O//\dcbb@gCeDG.P\L)SYGD\MX\\=G:P\7>K@S2#cOP[9b;.R]3DXD5
3TDB0-RW7eVE6#J#[?5S=U.6bPa33NN)b(U0H_bGfB7[/U=5O\2#I<H;WU011g;F
.OQ>79CW3UFB]\RWQBDE5Z0R1X#eGBG-1B/NNZPX11IgaF-^e2>O1.LQ]IdO,I6(
QUT\M2;N,eg2F>OZMY,E;_+CFY[f6;d--b-H?E7dD>RBOM6=N_TR<NDPOKO_[ZfN
XONH&a6.#8UD;-@PJNZW&:>3P1G3@TS[P]KJa2B8W0(M,^PNe)cgNPbNV+Q#=,dW
0e(;D^dFg;L7++4M)NM-e2/4HQT&M&HNGGTJSK?I6]AUD:)HB<;Wb&2I,843I-\-
7ebQIa0,#[/+Z8]:e?BY:?]?^GYC0]RRd61MNBFEe1CeQ(eVD8+/YGg>?1UG+)Z<
bf16bOSHAZK-;RX.3&,Ug-^T&I-gOTQ_ZFe:01=C;7UA0BE68F/6G:eNT..bfNc&
NfUIGaY#HOF/<aFGG3BIA&eX^R#7F@GN&TY.G8AJ\eOGFQ:A3X(Vd1/Y#1U>Q+_E
;]85FH\bG1;6>bZV^&<F9,+I3I4_]]Y&78G-JVVCZ7Jg=</:\XfI4/CA90?\83Tg
dI87-1<EV<9RF[0:.X3Y4WV,C3EA=>H2<A4=@f51Z5+^>f-HSY(H=ZS/Xg_>Ae,5
NJ^&3NQG-V^J(ZINBf.#0?V>B:Y(a]H8\d.H<<JeC+G/_.WfV^gF<&fJMRg@]Y8A
&(&6JWVFGe.9;>(S#^7JZgHZ)A.[8H;3A^3V:d@c>ARHIE2RJgd]+;7S0-4+VTQL
EB\.E@dWcB<\Od7=P7+AN?S-#KZBF04G3A/gDE>If?Q8(]HcY:+9H.3Z3-00,D@Z
[-5e8V(F/G/,\:Y-H&[#[;SbL(#fWWc=@149[GLcU1X0.)N6cYa7+EFIGIO.f^fe
8+1K0/OWa-G8=LNL_1>B8&C+D[50MPF<T_DV)Z?.+8Kcg+R\,O?J8[c9\K:H_e-(
2/aLR&+:K>8[H^eC4:0d:AKg54\@SX@L0f).F&36fGW]^24O4DW>:=Q]B;V^5M,W
12O7:Q@NOD8J/=?ga8>=-Y-4I?WUVgUDbf=[:M5_=647-1QST?]@feZFG#)483EF
,>&g4\Lf-(OdX4Ve=P65T9X.V6<SN0gUNJT+Eg_C6^dKX2eA0ReE5]Za2+RUSAEF
9FDYB5+-.NA)ZYG1)Pa@\MEVCQ;;g/D5Eba+TF8)7PcGNK@=UQ[c3];<Q0]C1P;4
bW0U?aRd,;:V79cHRDQ_b7eX)LPMNQ@JTfd\<<U:[1bdG5eK/gV+HDF?3g#-gA9N
K75ba\T<WO=NOID334^E-9c4/=2a1EJ7V6ZNJFbedPME+#_U6E\>8VTcA1&OfOCC
B#dDN+L(P6(?YeNe@/dJ-1)^c1MYS4c,LE]c@+Q??R,,[,CQPAK./c<f.QBc4RF1
J>ac>VOe.9>TR^X;NLPF:M&?9;FN(ZQTF&,E=(=/\>UR_JV+@B-\ab<^U:b67-cW
_?I\d&)=Be_a#=ST+UV=)[HI.+S7.fA?PH7PM7OB^8a6BdC&e&U[UZ6\NdJO-85G
L0)9#OGHUaK]]a6]RJ\92-@K1P5LJGKfdGO0Nb=BP,R=_7@J2NV7?Ra,M?55e#^X
+#PLZSLXfKGc,[-aK>3=(/[:9_NeYNM6Ve;IXYG>BGY<c/00(&\IJaC\F>/Pg_:>
::\2HOKH>UdV.C5K((\G(/@aS/K@Z=^2R>-/&0R>AKKNTXRQ4Ta&A#HJOU[_aKG2
1,dT.a#P.5(.;H(47XZR\42XS:OMF<[3JGOBO3ebZ<ZB]ZV@dH^82Pe<00=4[CJg
9BS]&J1acbB<4+FW[NaH7:SQVTD_3J]GD3P3[5-C^:F2+I9]0CZ2_g276W+5Z<PN
7bHY8O8D^b\LL&Y7E,g:aM;NAPF6.d/Z2g47@b-H/1WDbV?T;.gJBc??&H#G8,3M
\]e656?-F<1WP&N(Y(V35Lg3&+Jf;SMI270gCWO[eedOT#ZA_OMf-c4+/2Nbf/[f
:]+<2JW2,FZ1dZ0KX;\:C-dRa\D?K(63e_:6]=Z#1K#KDcIKBHZ6cGc60bT))=I^
1LXF5JWYM/84QA;aDL1c[&6W5X[eM]KY44\a7@f]C0,YXMb-#VD]//;9#>^\)AN^
fPKP7^Yb=]Q97eQ@-D;B/;MZbH[8W/_16/39Q7_9MC,]P3Z=NQ&fYg+,7L]6)\/.
<=Ebc5<91.b#-bc_>Q5_C58/DD12dTTD_8##?2,&L^Jf5E4c0:a-23d)7YCM&1ea
bG^HN^9[L)d&cR>I7U],QEZ2ROQ?bD6>GFQ]/aU8HG?)//&#5DCBT(?3424V+d/\
J]M>U_gCG\GTRP7]B]QTY0f[7/DB9dRXP#fJc??L2Z>fU1;JJGI7(D(Rd]W>?+6(
aecBJH_^X];^D=03.15@A#5a1\UVW4/HfO9a\&N64+)Y0C+QBPW&6O1WH;E+KZBS
Z3#Y:bc+SZ<eUVTJ4LRH,5^6KSDg?dcd9#EK_OL1#PR.67B.BF998dJ\7VS=5I9@
OD_C)DWO#0].+O??O?2V:XD42W_+]XM^4V2FAH<RMaFAV=4g.=_&M>6QYX-?)0-a
0g244.BEEd4R]IQ5<f)L;4BNKDR3,Z<Wf2[)Z&c;O95PeAJ(80DMQCe9,-UbV4-b
NX^N>HL?>P>F_cH^/-BIBfRdEE+CWB2gZ#,gf()C,.V;fD60d_<EFRf-+U;,+Q71
L>+Xe[6)ZP+M^<V>U2VWg0Y4IfS<d1b+E=>:@T78C6HP_.L[SZJ+0ZUd@)CA[aT7
W6:DI6>-6S;7J__TTQ]SNB.9^C\W\:5:Q3.K4N9)G7[f[.^eB_V^;S/G[:4.ZbVK
B+B&&4LZG&<ddgba>39,+^dDc[_+L7FTc6#&BVI;H@/I4CX>&L&,D;a9d.[AMQN(
B;Vf/T<[BRYd=<;W&d3QA>)>5e)4V8(ff8@g);4]Ef>T\8UQ#g/;)IV5L_UBY>EC
PL2eK._@1QZZE/@U^:0&H<A/cZ\H^_-:80JR6,IXJb6;Jd.X-Z0_-d7-BS9RAU-J
K_-Gc1-3aKBe_fg8.XWC\EDPb,52=U659:G8ZBDLGGSZ/WT4XVDW7?O:C>A)@We;
#0JDOBM27)#RL^E#96DG>44:aVC_a.gda,6R.Zb9]0W6C8C7KND\XR^M-)7EO#C[
7EYSZSeg#5d1.&(]bIN=6D>PX#:4AALNG3g^-]Z0LcY\_#4>/]G#ba]?TefX^N0e
NE[@EU^6ZMF\]4KI>TE.gAg=;XSeH_P0N4&O:YdD2T7ag4](5aLXBQBGAM,BV3,Q
;O91UK:DG)JXU?dLL]M1cT:Y;8&4?=F,e=Ge>@O4VKPU(4cdI46@ZX((&B[I=+E[
PJ7:E-V]#WYDVV<7Ib<=J@>4,SYf4KHIZa[1@^7g/6L[>eD@.:YBbJAP&\HS:4G/
RA6QK#LPFBSBJ@V[&DI2\JYPgZ]+#?G;5E08]ga8d4;@J0KOT=c;#LW>ZFW+/[GG
G(ZB41Y5;.,-/LE-N?6+?c6FO0N7.fJcSZ4V40@H#GEQN/gUef:CI:RU#+/eEM].
8eZS]\64,]g6gZL.8((68TXcKW2Qb1-C2Hb2Q,:VX4>adVbWYKVO9[S,bS?)(g6W
c7><fV;&?X:MEa\T]WJdL,-Eddb2f(V)6>]c4-/<1JC1f_X2);W<]H3[M1g-NA,U
YF,Ma=M9_YeUMO7Y]CAW_K6/)Rb9#S3:6/]D=UNGEaRc#C+?V^.GXWS1\5B]&K?4
UQec08.-,.#EWaZOPN)V.d@B&O+(90N@EF+;9__U+Y_=WVQ>S.D+;Ad#2b0b?LQC
b/IEIIUS<XBE)$
`endprotected


`endif

