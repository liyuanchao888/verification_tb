
`ifndef GUARD_SVT_AHB_DECODER_UVM_SV
`define GUARD_SVT_AHB_DECODER_UVM_SV

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
WP82BPaitpr9NizqH3Pqym2LCRZyCFLrkQ/GesYeJJJygFxu82FWQOJd9bKjlwYe
q6SNttgKk0cFfIQFKBQeAhx1fcFlKB6dydlO7V41nhY/GIy91mxfOsKfh4pgB0Mu
1mpdmMzhIqQu6OFmbxDivF5J/UEzkE1e/vmZESZhGzN33x6guPTcgA==
//pragma protect end_key_block
//pragma protect digest_block
zlgZs/eg47tLQeOoqvxGWslCiKA=
//pragma protect end_digest_block
//pragma protect data_block
iNYNfEeTb6r3uZB1WrF00zOXOQrF7FbeNMKBl6SMj/p1PFTiv8Uz3JYFgLEJJANS
wkhXIK4dmeBwdmB0MGwoFsL41h6xAjPemCtDHEzDKI2T1xxTFCwK5HXqHwTvEz2+
dtQcEFMwAlAKLbu2eQZ6CEQKZWHgdJ676MhAalj/RY1AL3IIBkafCfrGbJRF82v9
+Qxq2PvBgavwTVaDDfYRmBroqvIR+51qAphMjy4cJ7G3iIdpdthZXd2Sf7WOSZlj
BpozaY2J8Tpd+AKHzMUc5t0dHsgisGAudVswbMFqfrHbKsLUq6RsiUIHocYMC2Oy
6h2UawUXrdGmn9VUyCsDxt2oUniSMJy8JisjgRaKav/pJFaMoK+aIc54j2FsWwrX
1+RWf617ZEaThbFq5ti8nobTnvnRiANW0Vgzt2wT0mNTeLYcB+leK9na0hBwWWVA
72DE4ck/DwKjqhiY87iyskduRxfLAPegrwIpRoK6cetRZcwXe+VumEYm3/qho3ll
BaRVfu/GB6ww8yLTwX6FCd8w1ar4/y3XGkDq0S9Kb/AS7MJcGcUwIhl+qwUTg0TP
bGDyQroLr3JAgC21iuuVv/qGwYp40KhAhGAJrsIUmZ6zXNF+eAHEDTMt/u0eAuhb
fPGFOF2Uy+yhwP22pKm8GbZL9GqmVqaNVAwfp7AGPBffMYVauy9zKd9+TfjjT5fw
Lt2GCtG9Eq2k8IdqhyTvbhId7PeLAflZ5zHJ1pZ7b64=
//pragma protect end_data_block
//pragma protect digest_block
vbsiT172sbfKfHu1pcclZUHkNSs=
//pragma protect end_digest_block
//pragma protect end_protected

// =============================================================================
/** This class implements an AHB DECODER component. */
class svt_ahb_decoder extends svt_component;

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
TByHmShFz4GLrlfzSU35rldhLeK+vQh8S916v9wTmDu/EWVCKIcWjTi6n1Zr83zw
dou/dz8nialPcMPCHHeenM/+VJjnjMesyXlHSNwfDQeUfwULnDJkRhcirfbyX38q
hgtJ45JLb9mugyiBFqlV4b9xQQ6zGP2EY0+Sy9w8gViGr9rdsG7Izw==
//pragma protect end_key_block
//pragma protect digest_block
2dQhwuF5pvJfD+udjtwMT8WWE3Q=
//pragma protect end_digest_block
//pragma protect data_block
FaPKm3ronXrk5Yjpfh14Tajer6wI4d9RKKjJtspTser1E2RHB/n4G19jbAjfTd9/
DBf+BPXbttqT2GBUJ4FzMHPnD3uAfqj0REzJdJQSZtt/4ISiMTF+/NMkA2A911R4
kHy5LymI2hfQNe/QqWxNfEmAygCj0K61dmZ/XUpVm/ibeEwbclgYyQ7jBu0ItLKn
bRLJ6vu7tchROd0Nr3A7gLjkxxPKjew8TnG8nM3E3QriU+io7PHG8eqq7gMulxVb
kmXN5JLaZACnEY120MsHgJN+cGH4duTRfVAsUsFOSa324Du7j4TYd6gESQ6Le07Y
c7Zub8xVyCqeYY3KbChlSiRcX69LoRSwsOjaD+ZxxTzc5ZxRzszhIku+DBxCzwiu
1COKr/Y4gTxbjvIUSSNeYpeIf0bqjPUQ8wBNJLIbTkXgLszU0FhNZaqNcxn2to7Q
T9tktqOEJzSy8CvpfPmJOTnpi9UHwrZtFxyYMdIjnSNDSxVNIV9flBKxY3cbJAGN

//pragma protect end_data_block
//pragma protect digest_block
e9sRAGRkVfCLSsSwkeWGIjA18j0=
//pragma protect end_digest_block
//pragma protect end_protected

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************


  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  
  /** @cond PRIVATE */
  /** Common features of DECODER components */
  protected svt_ahb_decoder_common common;

  /** Configuration object copy to be used in set/get operations. */
  protected svt_ahb_bus_configuration cfg_snapshot;
  /** @endcond */

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /** Configuration object for this transactor. */
  local svt_ahb_bus_configuration cfg;

  /** Transaction counter */
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Gx8ZpRCQ4Y1SpJw0mM3mB+spkc8ALFMXSaTourpGd7OGS+fxg/lqU0mwBDORdbmI
pyUwvfMi1Y5C1D5kpr+UmQMPpXhZIi9kVUW1lE/yQF62slMFIRXvaezyBPofwyxR
wHzdzVUR46KEEsB1fzGr7RWcIBR4qJoGf8xeRV/QJxfOziYPUfoyeA==
//pragma protect end_key_block
//pragma protect digest_block
e8TA4tyzwz5gDXQWAeJxh9BO52Q=
//pragma protect end_digest_block
//pragma protect data_block
U29ZAY6imuiqdR2Gm4UBOwB3X5iI5U2imKFAVZYbGMTDsHzqQrHd2h36pTfSUeVO
qyFcCIMBDBq4Y7Syv1HROQ+T6M7F0qcZpELkCRuMmTRohEnhrWTaJFMGixSJxq/S
aAq2UW0eT3uVYWb8UEPutFoze679fO0Xs7Ab3EaghhgvuycqxuhDiqIGo3+5xaZQ
ETtEdQFzPQrmMXENLYWGc30fKTCK/cfMkiM2ihzVypmsBUYtx6PTIQIElj20AcLB
EBLY3/OWxhWErfMTm9GXRzoBHTTa7EEoAfpf1uYSex//1N09vuQgqw08v0jeWaxW
xY5VGPDL4RJ37GfDUDYVjE/huAHQdhgtGZ7TxSPZCi+4rtbC5VEwvtbgb3XiDi7R
w0FOFDYPm8CTAWbc4gTdH6e9/zRbkMkxOmIaVZXgPnhYKLs+/3u5XDYXifWUEVcK

//pragma protect end_data_block
//pragma protect digest_block
mkDdGBeAemX/xd8gKXzZvuj8KLE=
//pragma protect end_digest_block
//pragma protect end_protected
  local int xact_count = 0;

  // ****************************************************************************
  // Field Macros
  // ****************************************************************************
  `svt_xvm_component_utils_begin(svt_ahb_decoder)
    `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE)
  `svt_xvm_component_utils_end


  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new driver instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, `SVT_XVM(component) parent);

  // ---------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the common class
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual function void build();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Run phase
   * Starts persistent threads 
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif
  
/** @cond PRIVATE */
  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  //----------------------------------------------------------------------------
  /** PRIVATE METHODS */
  // ---------------------------------------------------------------------------


  // ---------------------------------------------------------------------------
  /** Method to set common */
  extern function void set_common(svt_ahb_decoder_common common);

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
c8DUWe27t4OnlR0vMhu0q9iakqaX63KqPWDidwkHawnVEDpuUoVcFn7RHqMoH7f7
D0OYVQd9k+Iqwf0NtIbk1Y+d7LaacV6glNXhTkrecBOmuB/SCv3uS38YtGhKJlZ8
oLOMKGKUXHt3+onhHAVEFNQtaRNaREdPheqZGVgakWpdwgeMqets8g==
//pragma protect end_key_block
//pragma protect digest_block
lC9XGenoXYJAiIpBQ75oiwCA+hw=
//pragma protect end_digest_block
//pragma protect data_block
8P4+L7kNjX6u2bzR2CfWuf+SZeJe1oBVNl9VSo/9tLTi1NHVH08/9j0PVREJjUfi
7sPoIS8BEXQ+j0Lr3ioP4LtdvdnzIMlrL21b91IjSJXrTb6M3WdBtPbz+JblE02b
ok5Y3GrSAtz4nYjJ3ZWuB3dsi+lUsCRzhPjIhEt/VgP8xBSV3Rf3SPKn/hflud+W
wxAiEOYA0j1zSaHxAcElvhx/X4T3Eg3k2o/4MpLNp4Nc/p1wbYXNzKDr8UbCHdpC
1uqiaKjGowahg/lmfzbTTmUWSSNxLz4lYxEDwgWFXdMmuOLcxgduPjodEf7/iLYK
rp3aPd6UmiPD1sxMxKVxNIqC12j2Ot3dbyjQBD1Y7RYt2u2XsrtWTbflIwbO5xb4

//pragma protect end_data_block
//pragma protect digest_block
LqEHybs7dvAojkTmLrzkfFO8Jkw=
//pragma protect end_digest_block
//pragma protect end_protected

/** @endcond */

endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ZlzGdGUaXj5Z5iDVuiBAMyZ2ZUV0Lj30Hh6yphYe17QA+k3kkTrj++oZyUk/0OVH
aI8nTGwnp1fhnPhXJXWcVK4v3tJ9ycQ3DGXACI4/dr+i/DoXgsXK6QStOd3NYleB
rTIdGodF1GNUEys2GIzaV8OMuc8zLRN0PGDLTbNHyG0KkdlXnoXEqw==
//pragma protect end_key_block
//pragma protect digest_block
2Osk5mHBW8vUGqdYhPzGUI+fuzU=
//pragma protect end_digest_block
//pragma protect data_block
1gZybwOsiGICbLSXlZ1/2wAQMwxRA/teVoxU0Fs8EEpc0ZW1kKQM0oqQREXnPpxA
CJY02zTpM3sibdy5sQ2OxKVlbpmLcLYvAMfpXF8pRs33d6sxIf/Pz48ST/RM2fvi
+7gp+SunRHOXRzgkKgTuxgME62UIK41wXP9I6i+UylalHpUjqghulzbvtCGIFwAf
/YxNNke+QhN3wA3V9XvkROr/6S0U0kgAagCqNfZC9nMGKD38jeGFRUr+D5Li8yzE
pyWmHeTf672sicxlt/TJNRe8k7YC+eqQovc4/XHKDl8ypwc44LPaZ2VyBJg7Bq0G
fQPC7QNBurcX/GP4qpDAcUBZs/6ykyl0iSWpzGRVi2iGTJQJPqm68GNp/h1Zt4je
slt6AJ23Yt4NxzTO0RnZJ+yiTg6sXrURQhzkaAmUZYLE5niy/Ic6wBgZ/EQ0WzHr
S+4Xk35aGFnOA8vhh9kf9v+zFEuiHQodJ0fdaDa0eGBaCfmj9S9vn77/yPuncYtq
CL4r8tduFJGvdZEvqJiB5GjUrbVyj7/d2YAkiTO4lVjRdGk8HrN6r26Un7uxdIg1
ZTt9dWlLzoQF/XT4T/eDIjFf0F6WKSqjXa8/YArE0wYCPP2jFtDNsruR1Viw0q9y
XALSL8bexgn99QEwzxDtfmhIC4lqqtjcWkr4rXHcrXr4b9PSwf2cMNYwwTnHMCWR
hzZdZnMF/AzBeDjhOdMKZfH0Qf/yb/J7y1crVy6vqelbCGvFv03K4+DBtvCHIKGJ
0L+LRNt2RSsMR197jwRDkrNlT+Oyh0XuTCj60beJU2FFLn8mg3idYLOTtilcgOOg
wSHyfBt8f8sSUpIEKcHsUg==
//pragma protect end_data_block
//pragma protect digest_block
NJ9u3C+3X279TI6UsEPPXqA4f6c=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
34J4QyhVKqrYsPYS2P9iDtHiF+uABzSRBaXWTltgKQqfQRhEVR7EefDqnXTuUMIF
uS/+Xp+R5kUTamHLSrJi7qfr1hO7KtL8COLvXAy5jko9tYJxNfb2h56mNYGMz6Ki
bqr2yJRrcoaB0a4GrXhXSozHUzWwZgAKEbH0QxaBecg2AlE9h0YY7w==
//pragma protect end_key_block
//pragma protect digest_block
XypbdT5/Hher7b2fEa+2SbsZdW8=
//pragma protect end_digest_block
//pragma protect data_block
enXJ0TEqiuaIFktUWWekopTc2KGDO3xed4gJY3jdUZXhqePThOOxvIPg8xKLbG/V
8IzJWSNxt6OxWGBchcGQ7rj3VRGNXAVWu09O6n2V1vlvm4pfKtgVXG+nJvacdfO8
ooUJESHG5pCjYR6LLsCzEriXpNpOakTpZc3F/gFMpHEDGQ3iJK+p8y8Bs1yR7k54
CIlFYXGR6lTm6RmGJEP5RQ3vZyESJEdAgU2mtVNJRv9rWZENbiKWDCeIUCr93MMr
q1CAjsIggeztckDe+mMU1ILcoU9f03CqY52XxO/6+HQEwLuhOFKpVnvuTxyn9V94
SGltXZq34Bugj2esBDuKpLO2Vy+nHLpOc7Vc13K62IgCTswH5VSptHdXKars88e/
w3pckJXQ+CqIYSXlMJyyqmMf6D7o/1I6txiVuTRTePpJQN1wiiDflYwGplMsAH5X
EQ1lgISmu61JyhJ+cDkZkTpvriCfGfBXeUE9W64rG48MJda/wxPHY1zfsibQSKgi
THi0bs+muIVAQ3/3fALWw3A1LqRYeSMabF24r8WXWQweJF8+x4sM4EmyVFKnvD9P
Iz+BTt7E6Cmv2kq6EMQ0fodw0KuXcMoEBMkjyEpxs6OaraMXBKr06+uBivVySkLt
kl7MdtHJarcZsfDpqC5WsBRo84ThFf6MOaa66gzWqQIaModGN4p4sZmXeF+IOJrc
q+sqtJpjGGrEXoOU28oxn3aP2uVxuaWCl+iIpOWtw74GVUa2mfnzyY61LW/s4CDV
RSXM9Bt0+CaKqT91yG90YPi8FdrY1xilKtVKRZj0/ezes+/2eZJzpAJiytvznk3u
NoUEzB+UdajXiXJkuBzE74MwPqeH8DONPS1nQY1MuoQgiSqhZhc8v0bmXGCACUa2
tq2v2ksvqqV602eKyqaJ/gBPGy1aeCu7yWV1tnGh4S0ko2U/mtvOiv4Mt3zT5ZMR
glfM+YfU4Tbk83dzrWEQe31UzkBfzfIpDfxWwLCmRaSGJH97C8AEwvDuc1Z4tHcN
A2tC2z/e69XdRo3YxsRb1i5Y7G3u5pmlKL0hWZ0wxldkhL6hGCXDdf3Mbel3xleb
aKyX/T+NscDj8tpNq/HAqj5okjoUmhh5lyXJCWfXvxDSZ6KH79Q++t6jJS0qfJAT
xVxNhcP/wS8Stg3DcPaeaZPO6kwF6Yk4jdEx37/09JWWnM9yUJuHAV+737tytIry
FWYIciV3XAsH3ue54x1BzA1fbcdsTwIq/44DF5Aq/m/N4TiicOI7VqfoXIl+7m03
oJO/+bJ0t3Oi3mWq/M4A7hlDDxxJuadO8TghCpt0gXNcgGZxmAI4EtXrV+zcIkvB
5HFwkYzTX0g9ceXSeX84yXWZYqV72T/zpjdf4wTu53AC0jd44dh+wBpjBMMBugk+
7yr8o2+4qUxetojwnv8vqrqKNB9bEOPuZAf70VGt33URuVPXM337Br56kI+E6spS
HK58eWP0958typ0JopzIgHAoH9x5EPn3GQYHEbFa4TZo+GuW7ydFfDcZ3nNCQ1+V
kwEAGYbMGGbuQuyOcUyV4HoZkzsSfmh8Uc/iP3mWlG9/ra1KNRoNyemgRUdTMllH
77iKzKvFwS2Lg4Rap+Y4KkklnAdtmirWqUBfOmdWwy/EYyBvvzrsOq311g4Z8gvx
uWEFVycPNHweeynVpI1aq0t/5zrzJqmM3JmYvT3vKwmi1U6G7CA9V5BQV3AJ8yvI
vdSbUfuMDsEVgN/IiLDdNr7+gQvnDVMkdiwM5dRAFkfdRzrhnnCaMmcdNaEZZBeP
CDc5NWAuPBs2VTGemS8YRTC8feyzXa5H/dMRrunU0Tw3/rlWyhJHgBkazOFI56DG
+EqgOJlw/zz4LAqUlkGMCNdxEf9lRPjSBkTu7MK971l1SEySKMSbPqQvNIPcSSn3
mhXxXYnMhJZrfa8uDSqb2ZT79J3a/pG9XXnUk8i8avQPzjAxVs2oKvvwIZMk7ZJy
v7xoR+cUxkwZCfEou3+nIVgqXwmv9UkQDibXfZGaRwdoFOoRZKZmw7JTCKcD1ELB
NgLS1tS3CDFNBrUaBA9RIQSXx2LK2OjXFmJA0acbpG4inkHt7+rdI7ihy/IqtC+q
tdH/pPip1v5TK236d8IoxAo19bPzjXEA68LEH5KZfuczqegCsBvvtlkXvknT6Z4R
/7xUz8Qu5Cna8QBN9oVitbQzpg/d2a73H0REk/QOHyTt6FLzE/mx5BBJ7LHv2RKl
dLqhVP7ZpiZXLX/WORzydNxIbjNYhGKNVV2DseRFK/DgRzttiKtJUv+wO5Oh/ynv
3JBLRU9DZEFkAHB4r1i8/1cY/jACcSn7ltgSQRNMXNwi4lDR5M545EIC3axCPtWr
A6hvxSkKjhEsV5oX5mBgPsWCDReNh2A8jXl30b++PdLugJdmg+q0c6iCGOQr30vo
NhZVXquWwmcHPc8z3EuMnykqXbd8dX1kTD/umNf7KS/wBiLuxMOzqv4V1bM4OE/r
LudETKPrRHSYgCN8fV0hBmgs7zqGKDIVZMHb5jPbNBKzJGw2KLOWmGoQNGOp/nIo
GR6u9QX4Hzcq2iHe2W1DRFJ0X8EY/JBDUlLmEFPIl90PXePGjy5PDXsOcO2nfkv6
BNFw25qH+f/4NR2XaCRDBThCIe9vU8Wmialsdq7xWu19UPk3LJ9jRHC6f8g4ZE9t
NaAMdGzGS5wtOGgu+hkSR7R9A+lI8qZ5D+qYExFtKO7zSsnmfi+MwWf7IdyMdzl7
Ngq/gKYNnaeKUYO0GE13V9TeDZZQ71MAWYH41i6YubU=
//pragma protect end_data_block
//pragma protect digest_block
bqT7e5T0T37webdUNrmkbuqOiC4=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
CexwURQQ0iw6aOu00ZhUhSiqdL1+ZjxlSsF8Zjaso0ycSUlmqMpOqXxBseJu1Fwo
qZdGOh06ujUscLPymQN1tvFFf47/ls1EwdCWm6xyvNUrLfoL4Lzi9H9zQDYp3JtP
+9+X/jGfqYM7etlRVLoKVDKTl9ICDjxYEHtU1hjRR6yqCxtLgSXKjA==
//pragma protect end_key_block
//pragma protect digest_block
O8gIEgMpThbFE+997bKiDiDZwDI=
//pragma protect end_digest_block
//pragma protect data_block
2WSItIEt9ZyiqWgAX4h7+q/oDSyLe5KQYlUzcliBizFu7uXU5NhgBf7YkofBp9JC
C95P/BrStlUUmkPqNvDUgEcJnNOw1q2vuixxZDQwR9aT7auuxEjc6ghJMTIXZA+6
OSrJmUoNb8MzQU+ON9WKHiwW9G64w8hyNH0WywB9Mx+LUQOu4yO2AoOy5fAvBGfG
rSOGScUdQfHzqxgZedUCu01P2dUOcpyhmURBKOvsW85n1pOswPPUVLOQhJHKgru2
XG/iYWfeI3W+IRkMXJ9uCjrxhbFAmRt5QEf6OhkArwlMr4ePrhet5eoDpPpSO5ar
y1kmY317tm40uaxdpFTZ73sT5d0oDj0YwqG4ZBS1LcK6e8NbAFyNlWRMYUEWlQL2
dtoXtFFWyhGSsK4qgK9t8A==
//pragma protect end_data_block
//pragma protect digest_block
FBHwpufMjA7QBGlawwvSIez4xsY=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
WeX7457h06/NfIWlNT/5zx57EnmwLzlejiNm9oAzGi1Q51VBVdYa3mIgzowi9E5U
BOaJ1R22AaBvCCetDQ1azeS1iH2YDnrhRPrBOgB7KUzgPb+y5sIr0E9HZd4KmIow
JXa4M++ohM1Ynu5dVOy3DQZpK5Ycyl6VZ9tsV8eowc1UhXa0JNJhrA==
//pragma protect end_key_block
//pragma protect digest_block
ws6Znq3Hbe9ykMxmiqbhGZfI2Ic=
//pragma protect end_digest_block
//pragma protect data_block
q8cxm+zb05UhCevR1zx73JQKBgaGib21WG+nYMA6tl9yi2n7B9LId+yr4+793qrh
pmBsUdHJilQKAnVqX8Zs/tkG5FXuD1AxlZWul2+l/SYlOvjLDNAWAWD5wgXwXn+l
1tWZlRrmU9nXr6DIix9+33UcCj8cR4oUSNJslj//cheIvqVLje8hAqNx+Zgxm685
6V+DGcwy/ysUC2gEKa2fWPQscwfWYiY3zu0pBeYQbCJk2L2idMTH9f+5Pi74izz6
Eeh66wsuvWPAcqsc602Euu4gUnBHmieuoj6LdH3M9G1gYm05ddlSLu6Jvmb03rw2
XkjnFH8gKl5qSip9J9325If0J3jeNzBgj53LBcn+QusdgHEyPodrGVh2/Bj2IDmJ
VirPLFQJAVZZ+vc+Nvu/3mOEWXohC07PLyb1jMmrfBjK1xOxVXCpwMPY67wuQCgj
bhwzzES+K9AmPc0IF2ZJoPcfMTW45iulku3/k8xbMDFyYPuxVbzDp8m8PgLI59yp
W5hznykE+RMt6kD9+VgXRlSgRKR0BLwJn2IFNXqwOUwpmufdmtipXaDuG/PB4qGs
mfM3AdrS4RcgBsmwZSf7O94h3aZHO4f6LuMiVyqLF0zpmiSGu6RtkYacEejcd1kZ
hISH5cUgKxhd53pkWuZqmDQrFEb7Nc3SNHiVoYQsq/FuzqIVKrQHPKIjN9O0UDv/
rv9NzzEziHmfdbPLqM3ImAum8dDX7/yr18qLspQnpbeuGYjibiO467Tol6wEFzhZ
XO8wYQW/4LNSqpghkg5aIHxIYYpAfSr8e47HRy/ggcipnK+eGqG4gs1z4SrbDpLd
g6Q/ogwEWkapSdhRKykPiCHeDnuWTAGJCn63no9ealZ+Vue3s2O8C68RNGP0hYW9
vZ/F8RCYsbRpVEV//mjI2xuSZxQyYfjTQ+HdOhvMIIMmx0x61PsRExSGHeLyA0fr
AJgn0IwoLHljdCvpq5KyDsQaPNgWrEyE5wEo/9mM7h9I+WWbTeKrB4O4CQ6PY/ni
DSoyoYV5YwXSTrgHvx92ipKXpaqU/VvsttjScnNTa/IvAIbOin0mbWyMc3egil0y
Y0O+9axHS51uKJnlPUSRVxU7NkNCydH0ePkwDBuOIzErK+uKZuFmkKETLW/CEO5a
7doB60fSrYzHGFm5mS4t1gwbiFNlsOc5rAWuVq1kA6YkUEeBr2f70BHclAw1Wf1u
IfyXJ6gyT5x1mzmZHB6/VGDJFRnyxt3Ry/Wa8+YRXOh92VGI5WPmdmAamOCDQYud
ELz5PR2MMIlIAysuPZ4btVt6VejmfZYBxhb7p8tdeCA6i+x9PVPtRCoDGXaDeY0J
hIv4DT7yne+IhQxOTLZDS2sA5La3kNMqw2obYjqD8/mOE+4lnpNHz+oyJdNSjb21
JTCh4+xla0fMuB4qpt0h5GoOHXl/ZB7KOysJkbyez4nOyhpCXzrjS36w6xBfjiPR
mZ290zbvEnQW1h8tnyOG0KaCZl4t1W68V82P9VW+gdVP3x7c69cPrrfPVPuSX/PL
8Nf9FwWlpAIZri4TG4Q0kgGoFwDNFuRn4yugxDmTpnmdVJ9jMHK/+j+BpzQJ20jD
UHYJED8hkWlZHmUPo3HSeHOBK3GHPcYKEzhkg5DBM7b38G8+7z7+amh9bUaevOKY
ZXx0pm+yJ361iTO4LkB5B9FA3T634ZFGUWg1BOoNekUznR26FW4o4ZsiZ2bi7BKi
Ob5n/kLg3WFRpxlg7TMjpsdP1oIUUP97s6PZY6SV3yqDHhYNHYyGArM3PeeetCOt
vBzoniQm8G1xIw6UxgezwSkazvDchOx67VOrA5XwPrLHjEx+i+wvUc9VvqA3WT62
XP9b1UnPGBJOSUsrjse56PybH07LPYrV49WIOm0mMMQgoSR/y+aYWlSWC9cLAGTU
LUlIR+jmvXIq3XTRRJwsiN6+IQbeotrgXwh40z2Fk8yH6y6Bxd4ekOsNorq5cP6j
Nuqct1A/i50OczLrvqfVJfq3zeQl3gXdBMQbqQJfjuOyST43lWJDJ2ol5DfyaVUK
gtyed1vpzw5r1wH9tgkrMIhC2wRMRZOBs3uW6OcHI5LWqOUR0F0AC6331oIRHu2i
nItLvNffEVXhO49rW4kpKnBPZxDPDk4TvI8tsPGIBcYKa50BvLzC+EHksfd1oych
txhHAtBnBE6zHgo+8caaMyrfCuA9BGOhGCySmBFNNOpq+3iv7mCvX3mjc94V9/Vw
Kyd1t1/4wPQUcpO90P0XQe3/txcCNb824jD0q+lNaPTMTXac4qCF5XF8WVannXNF
JrLs47MU4st14Xz/wVcyMkF+AUp3ubGX5D31dlikHzecS8ttYBW4vffT3mC40Ttq
HKYWWWZKHaiKRGGFD3NUA3bbaCrZ8L5zxmX6fPwOfL2ShrNv3TSgjvAENNtKtmlH
IuvXbjHZ17Wx4E52/8vCDiskLTAeQilv20BE826gcyHRh3blrWYmhmbv/2s4dRTT
bm/aQ9lxKCTNmXAQcC5LbHbnCInHZUQPCKNKnSJK3hjWgn8iPwqvsmBZkURcwN7C
nS+jqaYfXt+fHlDTggFU3DAHYpwspN3N0Q3gVHMC0yaikCUzk+HJWZT6GBNX0QUI
rv0B5/ySq6LL3pSBnj33EqgRX/wxkeJpCXLwp203UV5a6V/PJEb7f1Jdmm8+ndsA
6tRpmAwLmNBGSsbNv76lNBpETf7mY5e9mm8mQox8iTdGH6/Z4rS3iVhYesf7wtgK
o/zgh/dJjztWU59YuDxetfZsqZdOuHlLXif+L679GAlGDJ9M/PQG0MSqC3e9Ix1S
4eIC2z5hM87yRWjnPdCTDSCNoIyd5u6Ctr7nBn4mhCNwNURZQy8B7Y/ZsmcH6mn8
EYYMOK1MAymK78nzhvm6FMF3ZgMZlrds2UtDrfF0qvlqu6ujC/ws3/IM29uoAtQT
DGW0+7XIRssm1MTJh4T3jjh62OSevQ12orDRJWBEEVZUsXWvzrnQ1n1hQ9R/w2by
xoGH13euT6M0vaClWrqZ7ollN8ov/AGXsbPDjfEQMtUAHjpSEoHK/40fhZtX/weT
6VUH0DFRxP6YCs73V0YDZh9rOH+G8mBSO0GOS1S0zCMA1HROu4N+m2ECEvvtvCGM
B5h0aJdsCFSj2x/cLBwJViND17Vd1xsHZ7bfTCxR5kmtbWuYuSdWUUziXrnqJYKE

//pragma protect end_data_block
//pragma protect digest_block
B74KvbMTKWXvSVAHn1x/tdC9f24=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
zNbK6F2P5JhU0pfcfATj3fzdBF/z5SEqfuQ4OYMayS5FxibNzB0h1Byn1cG0pSO/
O9YHTM4RZb8dFEJmtph+ZWJpWzw2RfOPKYdH41wW70g9zLzTB3Y6DAcdzs5Htu3o
88JDflKT0csej7zJhqk3Av08Bwnh3le0wLEqnyJdm0bn54+jIgBL2Q==
//pragma protect end_key_block
//pragma protect digest_block
aPgSA9qgrXlWKRuZeoLnu6R0cIU=
//pragma protect end_digest_block
//pragma protect data_block
dx0b9WxsxBLm5XLGWPb7iBplML1nLHAz+zlPkuNhCbyE4MfblhFzLuXfed4CfYPR
jdjcXE+wzOCNLkV0yW2c58755lFjQgl+Jxb5tnXPFR+JMxgX88klmfxyMQ7I5cxL
v2zisITQ0zmhjHZQuJY+i90xTjQdxPbF34Vf4UsPvxz7Cz7NJf9g9WaB03kizlnu
8P8VxEY0BC99DjenGXBv37N54LwKLurFvma5K6JAP9D25O5Hde+1W31p6lMXyMKi
prRB/rvZTkDMRYn2VOTmhQL7B5PgHJugzJLVGYnZr9RGSmJ+RBmzNYwZIwcdY9MB
zRCuTq6VeEt0EjVpVvHCRnv7+dUY4hJhurVRAzla8gCKKCbvmFleczWGLBR3PsHi
QEw95DdmXkJVmbAjRF45fQ==
//pragma protect end_data_block
//pragma protect digest_block
dodvcpPcyKPkqH6cRZKhtH0hf4A=
//pragma protect end_digest_block
//pragma protect end_protected



// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
VbzWBUajfQ0LDjH1ifioz06Xjk9PnAbKblz8Z78kP2NFKiQ/bB/vLR1OU1LJaEaH
OPbmGFMHPSMn3udeMe0AnKi3UjxLU4vDxDl9VcdMFng7Gv7Csa5zcz+4QmVAP3h+
phgV08W1SYbfVkREYG1gCCHzZv/FWDRDMYJyMsQhTVUaKH7jRhErDw==
//pragma protect end_key_block
//pragma protect digest_block
pkCnr3Z2cy5wA5PVioOFX9qqOMk=
//pragma protect end_digest_block
//pragma protect data_block
fv9bzKpswOaMcoQeV1ULDwmAU7Y3oyM46vr400szKElKY3+U78MXsQk7ZhTacun2
HanZIVzcXiQZBT+GmqswN7rlIQvQ4AbGMdFtz7Bbj+AEJucOkmb7bQ8W/JTIZncz
fE1u+U+9f7mTNr6Vcej8RFz3he7nHSPiCvGO9QEZiF3+0g2dY3inYJVZqKzqQZHU
qTGHYISdeIaLdCyiRArdEMukWs3I/fs6atVfIGb13NMAAlZKZiMLaDFgL6AmhqFz
3aymHhVfusyUC0tKLjMD8aIsn2WrTiyeITYdsbhtUkizeYmajP4GGirYFKHeWUw5
2Ph857CtRzHJDRnXsN9TuA7+z2GrnImxPdbrwiim8FLPqCv0MxM9a9shTbyuSnRq
560TM6JrnMKMN5CJODrz1c0hQA2PyOEBNTFlcqaqD3dlVWEGjdZ/ATi9ETGdiuBJ
YiIj5L007p/7Nt+s4k0IxRW5ZhhAQ6PL8xc5VwXBp28W5QMCV3yj9ZZsYoaPesiq
JG4bWQixFQMvXt3yo+RQ6Q==
//pragma protect end_data_block
//pragma protect digest_block
VypwXxQAzb9xwmKaAF5hvUH1rGI=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3sSLT58cQt5cPGaHULyLqIvmMO4OCjsSxOMQ/N7w7MBLEw1wrnQFyU1oxDvkQqId
XVIDFgRQuYhfv/4wI9eXbwsQwsKhVlSVxDwbsKNskdebqG4tJqqFe+3+7Ry9W86E
gztIS34N7WUhmRcG+QXbVemk8WsxILW2amNhBdFwZj1AbRmY1d4+wg==
//pragma protect end_key_block
//pragma protect digest_block
b7x/sCE2MZFDhvBQTjiNotJ85jw=
//pragma protect end_digest_block
//pragma protect data_block
1wiphiDdKzevFpJXkmV8y9bZI4bw0klUFKV3DKzR7VZJFjLNzzPoI2l+57GvqDbW
shK6vxuqhrPzwygxn5R84HElGmWpFg36TvpFFugEhcNcPsKTlcdnihqZfdU25MJ4
hodp5lY/gVL7uLg94c2K9/7oTAgRso6jbsLercfyN7jspSVEm8beKpq6KQZ4fAtj
JmkWVUAnCnT+cw5fHSjGe5HvMG6ra+84+FCrZRDrXpuJm/yra8h71SYfUVsyvO+v
eog+6VAQbywD1r7EN++tdu/PNCkQu4ejFlo2trD3eXejcsAw5yzKFkjTRMwzW9nb
5O1qPg3ybAAh7gHPuVjhp4zaDw1JvV6eDVh25RwUTt667EySNjnZicaCdMnHeAza
LO6O9YUqOfzkDVyFPm4xJg==
//pragma protect end_data_block
//pragma protect digest_block
x5UkgvKinU38sjCWb1DLoL01DkU=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
uXN7N2WFEY2in32MSfbRT/cbbQ9HgTw0qjVzy/X7TAXhPP+hlfIErI2lHQCi0Dhr
k28o0QCM5U8e6CEnoaCeaYBEqTSwzKfpMdcJ1JGqoX70Db6eM/WcWm7AGWZhlxg8
ted0aKkWLQvTPpr5+z5n8PUTgFPIqfjbRadJxiWs34xVuPpZNzlR3Q==
//pragma protect end_key_block
//pragma protect digest_block
uP/atWOpsKHxFwF55Ai8/L41XPI=
//pragma protect end_digest_block
//pragma protect data_block
/vOJucyUYEiQ2KWRk+94SoeWcAT16wcyTVPHnSaqDcFxPRj020h72+DsUfO5tvRE
Nt2VImmo/6OFQWy0f2FRHmUkrBrQ69CjUbOyHfyhv0hMmTKq2P8fnfg5dx03d4kh
Ugt/xIwzFarp4CZ9PLFW4c9xmO9MwQ3tRjTKb0RfKnMftDAOPVUUZ8pIGi7TF2II
2FuB+gILu0rFOegFj5m09mLihw61BzKVtkAnmKih5zaSNCP0VVSVuxyRlZAiwJGR
twxCzz+9MgSmfmNeleictQuNVUPlMaIa57tn2ris6lOaey4mZnWTfEVQ4Y3bCMYj
mbl+33h7mOHPI1oHkCZQWqSExzenQxUfLQRvLAn3Pe3h0cKsU70pUC0WIxgBGmdn
MVaij3gQtfiF10krPfuXTQ==
//pragma protect end_data_block
//pragma protect digest_block
/QBRbzrBtqovEkV7P46qGq47nfQ=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
2XPGM4asFgeULilqslz3UArlBzyiWHrlcMP5ImV39PRHCHMB2x9E2LgfG0KFfLP4
aWs4PSDSEx+LKQ+Ht/73uzu99zkXN7SvpBh40YsJsBTMOo46e8dVLkWpeNsUgVL/
194l2L4SQVClP2i11qGR6WXtzPj3Ava51mq+z5epvHnNjQmMT1csFw==
//pragma protect end_key_block
//pragma protect digest_block
3l3idk7YgxFAMDNSj3mxdSImaPg=
//pragma protect end_digest_block
//pragma protect data_block
D+7z8xpKulrdVlc2XQDRlOazVVQ93on1DTtCQZNwxxBjq2WK/CGMoUUyaC0ggS2z
a1IGW5vw0RbMEf7Op63LSdKIHgagGxWzWlsBfVNXZYFM3sIlCRytnwCLceVxbHWE
nRjs/pZPpMMrWkutSg0VYFj/ngwxh8Le5D/1Ss/wZwaWLCR87oE26r7m6gaKkj3+
JmbXIaTZOQtztnrY8NCa9e+pQpyKg/2mMNw+WERHwshEd5snroH+ivPFPGhm4EJS
UofqQ44urkqu+qwmp8X35U72h9RXnUn53xCbEum2YLoQ+PlOtxt6f6qCjoTEAp4L
CfmBTtj+5aV/HJdd8PiKE5G9j9163OSNiyOdQR1NUXXRn8H7naf//MjkKsJB+v0L

//pragma protect end_data_block
//pragma protect digest_block
KWp0XTdVai07OxRfreGA1lDY1bw=
//pragma protect end_digest_block
//pragma protect end_protected

`endif // GUARD_SVT_AHB_DECODER_UVM_SV





