
`ifndef GUARD_SVT_AHB_COMMON_SV
`define GUARD_SVT_AHB_COMMON_SV

`include "svt_ahb_defines.svi"
typedef class svt_ahb_checker;
  
/** @cond PRIVATE */
// Note:
// This macro returns the width of data bus that needs to be driven.
`define SVT_AHB_COMMON_SHRINK_WIDTH_FOR_MAX(width) \
  ((`SVT_AHB_MAX_DATA_WIDTH > width) ? width : `SVT_AHB_MAX_DATA_WIDTH)

class svt_ahb_common;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  // The Analysis port for VMM are declared in the ahb_master_common, ahb_slave_common
  // respectively, which needs to be parameterized to the Initiators ahb_master_monitor,
  // ahb_slave_monitor respectively.
`ifndef SVT_VMM_TECHNOLOGY
   /** Analysis port makes observed tranactions available to the user */
  `SVT_XVM(analysis_port)#(svt_ahb_transaction) item_observed_port;
  svt_event_pool event_pool;
`endif
  
  /** Report/log object */
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_log log;
`else
  protected `SVT_XVM(report_object) reporter; 
`endif

 /** Handle to the checker class */
 svt_ahb_checker checks;

 /** Sticky flag that indicates whether the monitor has entered run phase */
 bit is_running = 0;


 // ****************************************************************************
 // Protected Data Properties
 // ****************************************************************************

 /** VMM Notify Object passed from the driver */ 
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_notify notify;
`endif

  /**
   * Flag updated by the active or passive common file which indicats that the
   * address phase is active.
   */
  protected bit address_phase_active = 0;

  /**
   * Flag updated by the active or passive common file which indicats that the
   * data phase is active.
   */
  protected bit data_phase_active;

  /** Event that is triggered when the reset event is detected */
  protected event reset_asserted;
  
  /** Event that is triggered when the posedge of hclk is detected */
  protected event clock_edge_detected;

  /** Flag that indicates that a reset condition is currently asserted. */
  protected bit reset_active = 1;

  /** Flag that indicates that at least one reset event has been observed. */
   bit first_reset_observed = 0;

  /** Flags that is set when a 0->1 transition of reset is observed */
  bit reset_transition_observed = 0;

  /** Sampled value of reset */
  logic observed_reset = 0;
 
  /** Event that indicates that current_data_beat_num is updated. */
  protected event updated_current_data_beat_num;
  /**
    * The configuration that will be used for the current time interval
    */
  svt_ahb_configuration curr_perf_config;

  /*
   * These are objects of previous transactions for tracking the active time to calculate 
   * throughput when perf_exclude_inactive_periods_for_throughput is set, and perf_inactivity_algorithm_type=EXCLUDE_ALL
   */ 
  svt_ahb_transaction prev_write_max, prev_write_min, prev_read_max, prev_read_min; 

  /**
    * New configuration submitted by user which may have updated performance
    * constraints and which need to be used at the next time interval
    */
  svt_ahb_configuration new_perf_config;
  
  /** Timer used for performance intervals */
  svt_timer perf_interval_timer;


  svt_amba_perf_rec_base  perf_rec_queue[$];

  bit stop_perf_timers = 0;

  svt_amba_perf_calc_base perf_max_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_min_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_max_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_min_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_max_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_min_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_max_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_min_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_max_write_throughput_calc;

  svt_amba_perf_calc_base perf_min_write_throughput_calc;

  svt_amba_perf_calc_base perf_max_read_throughput_calc;

  svt_amba_perf_calc_base perf_min_read_throughput_calc;


 // ****************************************************************************
 // Local Data Properties
 // ****************************************************************************

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_xactor xactor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param reporter report object used for messaging
   */
  extern function new (`SVT_XVM(report_object) reporter);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Samples the reset signal */
  extern virtual task sample_reset();

  /**Performs checks related to reset and update variables*/
  extern virtual task process_initial_reset();

  /** Detects initial reset */
  extern virtual function void detect_initial_reset();

  /**
   * Method that is called when reset is detected to allow components to clean up
   * internal flags.
   */
  extern virtual task update_on_reset();

  /** Initializes signals to default values*/
  extern virtual task initialize_signals();
  
  /** Triggers an event when the clock edge is detected */
  extern virtual task synchronize_to_hclk();

  /** Returns the expected data value for a particular beat based upon address, 
   *  datawidth and endianess.
   *  This is invoked for Write transaction by Master agent and for Read transaction by Slave agent
   */
`ifdef SVT_AHB_SLAVE_DRIVE_X_IF_MEMDATA_X  
  extern virtual function logic[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] generate_beat_data(int beat_num, logic[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] beat_data, svt_ahb_transaction xact);
`else  
  extern virtual function logic[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] generate_beat_data(int beat_num, bit[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] beat_data, svt_ahb_transaction xact);
`endif
 
  /** Method that is called to get information regarding the data/bytes for a transfer.
   * Currently tested and applicable for AHB_v6 incase of unaligned transfer.
   */
  extern virtual function void bytes_information_for_a_burst(int beat_num, logic [(`SVT_AHB_MAX_ADDR_WIDTH-1):0] beat_addr, svt_ahb_transaction xact, output int num_bytes_to_be_transferred,output int bytes_already_transferred,  output int num_bytes_remaining, output int num_bytes_for_curr_beat); 
  
  /** Returns the expected address value for a particular beat based upon address,
   *  datawidth and endianess */
  extern virtual function logic[(`SVT_AHB_MAX_ADDR_WIDTH - 1):0] generate_beat_address(int beat_num, svt_ahb_transaction xact);

  /** Returns the data value read from the port for a particular beat based upon address, 
   *  datawidth and endianess 
   *  This is invoked for Read transaction by Master agent and for Write transaction by Slave agent
   */
  extern virtual function bit[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] extract_beat_data(logic[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] data, int beat_num,svt_ahb_transaction xact, logic [`SVT_AHB_HBSTRB_PORT_WIDTH-1 :0] beat_bstrb);

`ifndef SVT_VMM_TECHNOLOGY  
  /** Returns a handle to the local event pool */
  extern function svt_event_pool get_event_pool();
`endif

  /** Creates the wait state timer */
  extern virtual function svt_timer create_wait_state_timer();

  /** Tracks wait state */
  extern virtual task track_wait_state_timeout();


    //-------------------------------------------------------------------
  //                       PERFORMANCE ANALYSIS
  //------------------------------------------------------------------
  /** Main task that tracks performance parameters */
  extern task track_performance_parameters();

  /** Updates performance parameters when a transaction ends */
  extern function void update_xact_performance_parameters(svt_ahb_transaction xact);

  /** Updates performance configuration parameters based on a new configuration*/
  extern function void update_performance_config_parameters();

  /** Collects performance statistics when an interval ends */
  extern function void collect_perf_stats();

  /** Creates all the performance classes used for calculation of each metric */
  extern function void create_perf_calc_base(svt_ahb_configuration cfg);

  /** Gets the performance report as a string */
  extern function string get_performance_report();

  /** Stops all performance monitoring and kills the thread that is tracking performance */
  extern function void stop_performance_monitoring();

  /** Enables/disables performance monitoring of each metric based on configuration*/
  extern function void check_performance_monitors(svt_ahb_configuration cfg);

  /** Enables/disables of all performance monitors based on the argument */
  extern function void set_performance_monitoring(bit enable_monitoring = 1);

  /** Prints performance analysis summary report. */
  extern function string get_summary_report(svt_amba_perf_rec_base perf_rec);

  /** Returns is_reset_active value. */
  extern function bit is_reset_active();

  /** Perform signal level checks during reste*/
  extern virtual function void perform_signal_level_checks_during_reset (
                                                                         bit                                         is_common_reset_mode,
                                                                         bit                                         is_ahb_lite,
                                                                         bit                                         is_master,
                                                                         bit                                         is_active,
                                                                         bit                                         checks_enable,
                                                                         logic [(`SVT_AHB_MAX_ADDR_WIDTH- 1):0]      observed_haddr,
                                                                         `ifdef SVT_AHB_V6_ENABLE
                                                                         logic[(`SVT_AHB_HBSTRB_PORT_WIDTH-1) :0]    observed_hbstrb,
                                                                         logic                                       observed_hunalign,
                                                                         `endif
                                                                         logic                                       observed_hwrite,
                                                                         logic [(`SVT_AHB_HTRANS_PORT_WIDTH- 1):0]   observed_htrans,
                                                                         logic [(`SVT_AHB_HSIZE_PORT_WIDTH- 1):0]    observed_hsize,
                                                                         logic [(`SVT_AHB_HBURST_PORT_WIDTH- 1):0]   observed_hburst,
                                                                         logic [(`SVT_AHB_HPROT_PORT_WIDTH- 1):0]    observed_hprot,
                                                                         logic                                       observed_hnonsec,
                                                                         logic                                       observed_hlock, //hmastlock for slave
                                                                         logic                                       observed_hbusreq,
                                                                         logic                                       observed_hgrant,
                                                                         logic [(`SVT_AHB_MAX_HSEL_WIDTH- 1):0]      observed_hsel,
                                                                         logic [(`SVT_AHB_HMASTER_PORT_WIDTH - 1):0] observed_hmaster,
                                                                         logic                                       observed_hready_in,
                                                                         logic                                       observed_hready
                                                                         );
  
endclass
/** @endcond */

//----------------------------------------------------------------------------

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
l/d9zBFrLL9HFYdqB9As3EuP+eXV9sEMq9NUyv8H2n448tiz81vc/2fVudypFEXE
lEb1zlKkmVD/pIHdDiNSF51XAjgZYLzbckaztTbO9UErOxWKWGl98czmtiZ5z6il
D4pn4p6ISVSNRfNXqTOnpQbTNdu5oggt6pkPNU+xNLE0d8i5PEYY4w==
//pragma protect end_key_block
//pragma protect digest_block
nsuuC9CfdGtemXAVIjgLMWwejrU=
//pragma protect end_digest_block
//pragma protect data_block
Oxt9QnsB6YAKpEJiV+4fwO4urPVtcJaxJW1xFeWCSstbTRLsLm80vwnE0kc+pbDG
UsRKkCTiUcT+rmi+JP3bNI/qIFBPprrdiYPwJ4YSZ1HgTEL5KkTk/Agf0HVJ5pYg
2uYbcFXZ+m4TDCVqEd60Dms6pT+znEQxF1mQz3NzeaMMX2bpDyQTwhDBqTNnhyqf
mDuXTMgitB+yp807s6Cn+LNITKLxfrDvjPW5rs27NvW4tblnDvLe30LoXB+N/xXV
nIYU8jbOBMYB6myWBvTGaO166k63JwI96uc6c3Hzv1IxYLePgUY+YN518u0QEbCj
CGA/rgmtCUbZFV76IJBIXNJkHiITS1AMbqW/4S0V1zkpCFCe4bZFoK4b+llXVtwz
IaUBXf8drGsOCljn6S33b4QehLrh3JWe4l+q2LBojamjguFfsVhViTCiAMjnRQ3m
Qo2elHwp7iUhGCx5LdXl7vJRwOsbUELSnvQEGdJCqUd9CfhB70daMLXYRgWJbrqu
EgseeAKV2hdpvZVuWFzE/CGKlxbzQbPFVgTYorgKa66eYtIPohhUfkiWVVSX3RXK
70JmXy+LtR7Bh04AezDG9MHk9awnLFpEB+T3Wr2cKOTEAjZ7IUfNE7Cex1KO/Grk
6heXvh1eAtH4fDXO+qRpE0tJZLxCB/n1XlmMhnZLA+o=
//pragma protect end_data_block
//pragma protect digest_block
zHwnOO8BQqvthjI8iISk1dgJZ5M=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Cc5tcxfAaABPwRcK8ObiJlmYRC2L2KKcEsp85l6SvwQCjMd9c+9b6n9E1pXdJrlj
Aup3F97mcoulS+b8EbAoZ3Yjy0aLj1FprGnfVf7Z0jUGVkbcvehSSwAPh5H242BT
U1gg0qe8Veg3eTN2eWGDvC8lgdQDI5VlikcB8wvRht69gMY+LFe/Ig==
//pragma protect end_key_block
//pragma protect digest_block
eGZcx0UM6SG3oW3Unyh762uGYNc=
//pragma protect end_digest_block
//pragma protect data_block
ZTI0gsoCpeYT+EkelG/vva6wIedXtqu7V1kecxq55yHwnw+C/MiLMT7/XZHwMCWe
iVWcxvv1Kz6U+YiZ1PL9Oaeq2cVpZ6A2ugvoxlgsV2/mU/obsmgbEW4JcDUggKjI
Pm+AZWpwTdM3h0+8o7IcZbJ5r1ojpiqYTydSfbYWb70zs5fTe63S46VHtXBRrLTv
UC1WaFkQCyB0wPmrjk716NKBAEik/8DIAbMn3k+lguWD081PxLX52ciEo8/F8a+2
iFfA4C0528Qqaf5dtHswNeoZ4wol2uVcimFY2UjWTzBKVabmnL/YUASbEQD60Yb5
r4+EKOKArC/5hS4TiJsLyfCvSfSirzt9Le7zzHvSCrkfwU6zjcSVJw5nr/YpajNU
J6dKH3sMDpImz1pV6aXo4BPwkp6Rj0abZFBv30mrRR/RkmPZqwAzjfsCGuqE0UkS
rcrD3Ln/wn9mhX5nrBtfCBfGyth15JB754RYiTNc6jiJvd+QaywfeB8rM7BtfrAR
xRKi2sTo6ZGQXoMlKbsK2eXjlm3c1m21mFYnkBlqeo2X3cYw4lu/xFhcbf96gw8G
nniPWjLTc33cjhN0TP4aVSMT9SJXNYuUn9rdIlFP+ZDJSRZ82Hr46qjXNsTD8i6b
v3hzJka3eUoGg9Kgtgz2C9GDaG14MqhUgMKVYYKOamf2bUirw7OzpckKuDG1FXBH
f7oXYcmYnAdvrEH5BTrRbNknheeH8sOw6wvDZxDm+p9sIggH8TuDe3cw5AcZEyGy
pPmq/9kgV76tawTF32k0GA1qBcaMZx0ADEEff6TqW8rV3dLRWUaoAeNwjQwNzgtq
ueNZu8TM4SPusRQUwdn4oYABGJlqbci9NkAK4otkd+IQjgBDnVx1jKBCGcpWJ9vX
LG1s+bXjsxFS+CWcRq6ioyapJQzEE66WNvvzIUMry5y1Yg3zu7sOHAkoKOm6giag
TPnjP1kkAbgTfcOCVjRNpgEjuUxDXa9RLVilyO5TeAOYdQNLeGZ9Q5HC+eyZd0EG
XrHtw0woALgitzyw6RRMVIUDYuF22Za1YzHK2m7OH3uxRNcbTONKhwCmkuKypnfH
NRWcSmivlakgXYGJ4lDK4Jqk9w/pRyzwL9o+GFonN4BncNHu10MFIBDHRcPlFQ0n
gEBcZQobGhpzFNVIeY8A6+r09+Zd0L1lYOvGAeF8yf8xBcf7nUSXBfiBYq7oOsEd
kLpvnOFYbS3W/QQqnRwtUAtsedoQi+/dDtPPzizpTueK20hHDoZJIfKIWxxohTQt
bb7WFXqkQ3kmtZCIGEWQbFMwiqFeqGXlJtCEkaw/SVik+0/7ZxJ5L1iNPNrmd5hu
TonVzyQxXR1o5wEiGfyhsu+Ocbi8fpLPDRW9oIEfdDNghzfCMggh0nzb7DPjBCh0
dp7ej+4LD6HG1yJHvyuXuAwR98fjaSZg24feG6Ir/U4CiKabB6ptLOZdtKOdzf9B
OxY18AaNwgrC8gEjDR+OCGhcHioOIkhFrDvSm4Z54dZR1TXcN+em7GEe84rKLOnl
QUFRP6w/tGs4FdDO3QMn9pj3lqZ8d4OzF4TOuMtexMhWhUcdFwaX5BEMTaAJUVym
L1moujJyohTWnwZJeMH30Yep3BmDhw3FMSINuJvgZP4D6IZcrrQLnjnRVkeMSVej
e5d+ZtkG8ew2Eb2rQKoRtqozQxW962yheM+efP5udYEe/bABKpmeT2RkvAprOMEw
wp0BOsHzn+wn8Yl/yV2fxxZa2JIYwJQiuXCkY52tnkiXu08GJWx9/OM48HyMBtid
rTDBKJzqCwHGppNYiRYXc+omRi87rlwilinhplgkWaCdAlhDLZwsXXSyiODf1k8D
Ejo2IkzRESH5XPY6iC7A/Nm5AMS8yXIjVfdmsIKIWB9BxQuZl+P9EbEBMWMvEd2b
IvAstMDu+Ju3FBH8nRCddqHX3IyV4IKb8riRBnvPvvUdOdAw5ROW84zClOsz11L9
yuOzLSQpSZs1qmX4erlR3Wm36CiSp1vmexwRdjxtCqsWDA4QldgskRk9x7UJjG65
OyWvTEMXI2tZkL/1Qo69bfUiHv/ZaXcCLJ2ric/eAAXsEJLRsmy2YN1khaTW+7QY
7SK9vCgoK2A0bv2HMbLSO6vo9f1P3lLw2+P/fZZoIa17+7AGG1ZO4WgmQke15Zns
2v+rPszKF2xGp/oDK9+MBxB8dN33LDn2O8pIRwxUAFDelR7RO/Im/OuK4ZG6A4RB
ujNL8V9c9EmtXlPvyuvLo7WpsZCpUnagJFWXnoNtMF0I6bgL2prhnXpko/4O34m7
gZodEcYdS3cwtFf07Dv5FmhB4nSB19PpduoPIVW9Tetyb6oT0XXNEbag63fwn2vK
mOItk9VyI2lBnNK9BNAzNiePnc99aSAFzxiqUV+oedfFsqPgVY8CHypOqnIhusU3
XEgRtLSnFaiieLk9Abn2Og2QdudTGWkQNbW3DxnANSvsOTQR4XPYXrNzVqzpCcyB
dhFXrbNeuk1WTYcAnv9KeKw1YXZNf6IID2IZroz8ahtElX7g+NJGZ8nND7d6GsMt
BqXZoNbUSgpSyIbRbleSLXI8N8m97/JSXLpdohAWqg93vGmUyBOEngNC6ayfdfPg
4MG32zKXxKbD9FoGDHBRVGvXl75WltX/eFyUL+Li4kws7lh4eVLMYlSilI4ulOte
AnitYe5ka+5ssQFtXQc/TEekCC9ZMHVxQ3qwM6La2lcRJqALRgCfrO2qxsMpJunp
8vA+vu7y795wXj+AHwKbm3VUbA7UIeVBVDBxLfWpzCVoo4zj2h16P/DQvrxT+Sij
WVhA1PV1im9cHTwerB/uSzjetmZ+RjHbv3PwjwtmGInWGvCMcQYaox83wBZyoncL
1fnWyryZ5J0SJIcn4q1oSwAXJbBzmaNuKx01khZt/t0JI0Qs77RiyVxOytcYXmb+
YIgLFVKGYb7dhx4OZ6ihANn5/nKazY0OCfcmIsmuDVZyfufNVJtkStb2Ww6bwHVK
rOPB/duDwN12tNvs09zAsEdkZiUyz/nB0SzZ7gxGhkoSz72ixGxC/GsBJDgPPAyW
h+Atz5iHDzR/nVndvmFTmcYGcLJniflg5LJ8Nqfo9Tm06OBWKjBX9cbqdlvweJDV
iqljbOY0vFFphQz/+Ub3Yc3BgGjPu2xqGwRa6Vg3iOpWODTvAKiZjjLn8DhnfM9b
eMZFNH70r/WO94+dUQveVKYbV7cwdVVXYetEX9BWySXIT+qLQvn9Dq8dd5oRUmgD
HlMkA5BATJZhpw9AGQHm0t2EGPxsv7djcvKzcL2Ud543kw7DASOD6paoND8ljyN6
ospoERp7AeljJACRBTqngLQoH6xc/AxkdvGCg61UTY+PbNlLYVtJaLnEQtfFyQ2k
CsaK7sFsNG6kClUPs02z/0HD9nfTDqqqfnGoVMTH8Oqeiu1mXy8enY4FBvpaLCmP
rjkqKKk2yBzwjszR20fK5WvfNbtnAcc13hRJHZR4qlJWYhF1s38zPmrrESRQM3bG
TKOyWgZ54INuyC2g3AfGgWYkLq32+rMt+m2csXgXJUqJ7RE4FI/80Cz0MEhDfRi8
uVNV3M7zpNqFgnPy4g9EvGNq17wXGRaOpXf+sWobNevUvk1V/iVtGUtunvOkPlrM
Baccux2MZgEMC+3rgZbiLolnPvEeC4TJRser/2JVJvOoViix7WJmu1QZPCr9imOq
70zzM1U2vThQr48LIwGjD5sB95lU1lM5dE1M+kstfZ/sIf4gXGp9kAEF/czXqBzR
Fs6hq1EPEZ5xdFuBzMuY0uLx2Vm0bTqFtA+5OEhpV/v7eQnim/W7uiF5L6tMnrSg
ZhEb6nkse5l8M+51zCCLM/WtKeZldxEMz/vyMFfA6MQ7QBLk+XuJHg8qEKm8CjKz
BrRTfYYOtvqkLQFKCB5gWigUfDq9pUkOfjfdW6CEjFhiWednsjZaOzTts4OBoDEM
3n5yJykrdbnUsPjMwIvYRJmlCqGw//imZbsDON43a5tm2kJrPOs00YsE9lHuqIvU
nCRkgZgwYo6uyf5GWchB22Bv93QyMGVM8/LYTh+3D8SBN4VVzHBPj2gbuCdph1hT
mUQbWehkcZbI6+b/TBQhlpsvLNH0SNKPCQUGzfKkaUirSpbMF40UyB9skrn2jr6N
7K6nTrXQR9DNaACfKlALL5Zk3xL0oPm4fbB7OiD6tk8qmWktZxgj8JFt5YeqroQM
E40VcC+bENQBe6X2vqFV1vNPPFN9tQUEeDOrX6i9e15PzZeSB1/TaKybtnRwVyH6
LKSkQ2YTf40YskrqpvcUckfW5s8tYbltuFTgNY2k4EQcIx6vTClQn5TRIbU1XxQw
ScFQsI2eGtXVoNFNT+0px3tJvzbHzOk2f8A6i9Eo05qjBtu62Cz0VRISUJifYqa4
D9NaOyASc7gLcSxm6C8FkRLkzEQj5MR4E5VNGc1DatAC4yt2RUlHlHyNCVsTWuVH
Lnklq7n3GhXU8D/0AIMXE/lMF8q785z/WqO937l9u9bH6g0iIQyUs5GOEez/nnfX
kV5n/NKT7L61CZ46iOHOy3zYgQYAD3QbXA2m1MnqQ9gkoX2HJ+Dv8p011AlWk/+K
uDFGJe5FO+ByFOqS+CglyP2Zqpb5QcVWmYPA4OsAB7ob9277c7IShctderT1BkEH
URQRd3fkNxLa3qeWujnvSEBtKQwN2NoXNw/PxqG4APknSDJ4UfKACiwn9uP/c4kJ
3t10cSjtftYOyOM1VEOl3xscmWM2DxQK7qRXM9CtsApUJlX3OfGnGInSPIgtmKzw
ZSiaDkeqHobHHUHhQKXKo1hK4C/xMF6nW/lrl9MYc+p2zhz+HfIE7ZfSyB0l2/01
YqvcTRZYRtoo5qftsoxxemrLSottfiLsqw6YjwgLCAkMBc4OZNPnSq1j3FhWoFrA
/6eE7zwVzXZYuBFPaGidAcRPrSyrpHpJIebI6QCptoZQVVaYaEu8rYsHhNcgYvix
yEZB17nDKSYhfJzZ1iuI9r/0nZuc39fxjVnsWg8gH+xQHzkg6mGXLXR+9sDXD9Iu
kVA5ouyHhGSY5IWmITZ+lSqm7kJ0YQNb2zN5hwb4pe6PLgdqRvaxWl9izdZcfKJx
7MBJbw0odujLmtLQ25zvuqYpJjY5RzWCvdsfLICrSR8ss9elxx+JGa+/UmWADNn6
WNGiyAc6Zt+xI+BQFIkEKcCVpLH2z867CsOZmOvqJI3MAdtXFI1FD6ExyxF+L6fp
VjtUYbyTFfZHfeZn/YCuzoxMlWCSwkW683Chi4yxxaNqc5P3m6JqGJxyu47vLfKb
8GN8rmeey7YI4UyqAje//lV0uH/rKMJFJaexwaUiYMgh5CxF+SbhThMnhhCH9gxm
jwbXCVslwbF4rof1GbES7QqY9csKPTUq6Ua7eXCMvlkUwO6mQ8HgtHPYbmNUqt7Q
yA9IpR+FQXfrpt9Y+4LdSzSaYgQpucg93Nu+As8sIjY66PGn68CIlICPLinKUBZG
I1/xRgQgQzd9T/IEjJwcGZCkHm4qsNCj6Z+5HGz547V6QlVHcxk4CBLLfvbNxK7e
Sr/Y9Jr2z5V1WY9SbhNoNW0TsEyRppmr6VpUOrYaAOosk8ISitQuvn4aT0DcP4XJ
/tSTsomDpipFHUxqNLVsW9u5Ccn+xlDfA2r9bAlnM/e2L70dPg7YGi03locit3k4
cK5CtQBe5/lJixTmBUXMkQckytrB3le8eMDkhbqM/4Qt6l6IcRlRVp9jZPW+OjM7
UtMGPKYCgJITV+71EdLbhr1K3S6UGwsHsH+Js9cY/I01fo5xhOHmiFgmqjwaKyiK
GoOjER/GCxX+5YLcAECxKCWtxXCV+XhOeAp8r3MPWvW4ROpS7T8w+nuEhLCwTtaM
rXKfLvvvHiraZzJo+oP1RjAHoecA9bfhRTIIJAa0M7lFNbPQjsgmraNoWneddAF/
CJ7EFl3lkPRoHGctldaE4Xp8Let7QeutXD98SH17Y1lvSwvpPUF4V9UyzNT3Hx/A
ZtcCLQca2x+qb6vVV+hAzssZZ8AuDSugfxx3TNAj4zXSMruwWM3DX2o62VUH67Z8
hYm1JdNt9DMnHYtL3n+FI4shZVfgCTKW4lVYSfq+DNzW4aKXKGYRh4jDbimjrXe8
IAdQZLRk3TzEEluhGkmhBtOSnXwMIvpVGk0pTkzsKij5sJx5g8ZcBW1F5JiLlo95
ZWshfkFW3xb0pA5tKu4tbE6ttNfOz/6WY37Sx+1FlLjPImspW02hxt5kGpLb++8s
9dnU26KghTp8JEXQU0obIu1wYMICiL5JJlyrS3eJnMU0MRMC9ZNuJHeoYDbThYQR
At9HZII7SQ/+VuUAVlZj//ofHgo12Kxr/15OWAek62atJ0Rj40SP3rvyq8igCQTH
YNpKMcaz8TEicnEcsTGwoqsODATaVKsONQIsqVjQjxLoCxUpEDG4Xd4GVMn36A39
zJucW9D3RDn0BvUU5H+2YSPsJ4gT68b0KFaAgRmnr8NI4zx5JMXcEQZW0pCrqLRb
Le8fQ0ai46lBe9y+nGsZ4xK1Din550K5Vpz62EWDfUEjcvZ1Egn6oQ7KBj3FKuaD
/c7CuzB1OXySMVyYIBJZtFWpMLplhZS63bhwOjeS+ZDCtE58bV+Ajz1vKQQPb7bv
ZHhnadgtHctLOIBz6NTvzQox9qjVfMsyd9GWKHXFiCqgfPWS+hZIt3GtiF3Aqit/
tHsHG655YBjx/cUHrgI7Hc3rDU0XITAXfW//M8w5Ab8WOS/GNaXJu2JSdgDiK/A1
J+1Yd+g4RGdvSuORcbCKz1YOhrQKi+q21GSl9ZS862vwt+RFEA2ZgENAXaGV6xwP
6ylO8ef3nBkzE1eLRZFL/vq/47xy952Enc6rolIlvCmr1jSA90jwlkXVU3Sfmd/w
7I9lFxOgDGoduAyRJHwv8BPtILz/2xEwWqtahPJQj/U4gZQ+OrD0ZpaM4+nrmAdQ
I1bxX0szLZbRGJcAUGHDlMHDuJTd7sXzLuzRY3s8xHn0yqcsAkqvz4OSyut3dznn
jKsHoGv5yRfy0yHlf8ygAkcrNnGL6Z/39BjRf2jrzE6yxIbTfUuirv9xxrpIpDvJ
ja27iWNkHnJ8KbFRDDwHJaaKg0dTL/EXm8VGRsXwIpZT5j/E1jfe+ZJhyDLY4EqI
ot9FpbzSWgHxPbdA7GFvF+o4RcBC/Z/+VimTOeBqYn3bKmxWw4Xp7T3lh/u1HlO9
nbXLMzvp81LbyV19NyIxcj31RX8o8/BVDZB8Pq3Mcc6Y4xfjxq1GIUOK/VSVGrWe
aT49U42v6COyytGUuadRazNK5XcNjPNguHxUPLgBoVREob7f71HArj8RQK2wcz2I
22GI4NrgyHcELODWP2IS8A1tOdzdvnYNyMQvoB5RbNXbDzsH5lLtCd0UrDTqA1QK
qr9Xjnf5Ln1mISGC+G+VCN3xJewzc8Hyrc81TNhLcuRuyCkU+hOJfSGMAkaq5IoW
brFXWEQPrIbbJZZTpeyUARKgKhI2ZR53UF70nnRyrae9TzjSj+4RXZbOSzCuMZpm
NRTTeYXzzeUkNaUwa0arwJWCnCbLTVxHA7Uw4+skhLVLVpXcW9sa8ztW5mAR5zMs
edjWUTn2w6dcsrn1Sh11k3cSgkYrS+7QuHiWpBb5trNaXNj4UrEy8QjkCtRN0P/F
PtBdlxJOm/Y2JAcIBfshw2Lw8Z9dbNTWX4SCxDy+wrHJJWOKI7RousSRspYe6sry
IHFgHuhaD/3pj0B5Vb1d1izUyzprVHson3vgkZMCz7nIzY458LiCR7O8o6r66148
aNwBLcGYvfmlNBcFcaNjUuGqLZV4WZB++KLqfp8Yiqm1kpICn9Ug5ljkndzJWdBI
xBLmOo8pNwZerM8YpLKAbFDcwgI//6KSMorg+E8iKgPtAlyR+cCUbOWhH7+ATyeX
A2yr7SeywRabmML3KsM1lZ50p4ahnq4SOR2bMfM0gJmaZTDpv5KD2dwCn8pL7S9H
RGrmazAlgceIabXbmAdex8GyPSQI1vpTAkJVV4Bp7nNsetmMYS3uHG7Szk8aboIn
BfAFX3gFHsaOYCX/QoWrxJLvF+6+/BE6pMzLYI1BEZdy0cqExAhmKM7/FsbsLZXa
qeubgwJEnImXCpdAzycuOnu6ZcibrWB3tRk3bnwfDVE53YMueB2wLs2PdUbn3xJh
qYMYz2Tfj3BIfVeZF1IQOhO2vYI6+5LvvMBRgeyAlZWolgYjWYBY6OONPRJ28bgG
xUtw5wOM9xlRc7oyDGIt4BIjetUAvDzzZHL8r4EoHbTLXT8xbt5KKH+dAn8Fk2Wv
xpAtIF3rsA+dSMgQKPICle+blUUUuXJUd0qFI/E0hYGF9NaAXTHfGzlHn0N8jQWB
M6bCOj1cp6pfgZoIvu2Z3QscBM/2K+MNiVWW3cyjfDsVb67eA2gI2+Gnd+jePO3Q
gexiwqK+wU86L4LPZ8737SlnNkrAKA175iUTOE4KQF3wqMztdhpEE8YlqnVGdCDY
9rSqRX8qdtguk7AXCXAaznMYbroFfgtocvykt6lkBr98kKg0Tb7W+ETSytiP2xVN
C2saBMv3tKaaw7ktl067Tau1WI4iZgdUz5esSaiz4XbriLuhyhdJFwZc97HUGWpS
2TincWVxxBpMM0mzFcc8awot+109T6QkGxfPcnLoPuYDabtLiCOq/uH+e0EuLdlo
nGoUF0gzjMjGnIzVTmr2DehLLnHEgcFAYm7EO9YDvqG88s7p3ap80K6fgG1Ue2jK
waBtAmzFyMT7v9bc43bCc55G02CXkQm4tFc0PxC/aoATaklIfH8fz6VGcRglFgg/
uI9R8HSY8Ukx38H5CK5pqswYKsQS7GywTm2Vb9W6Wj5Dd6M3tdaGQycVLWMBd9ot
gbKvXI75McGC30/700xexm5K4FyX4ygv7z357Sxff1tyAY+jro9+FZKAKqBJTfXQ
YR3xtM52l70gzt3BYxtUET49dpxlarHScfu9VduIoIFMrsJg4xnVOtUwytf5urpE
cKTpot7IML4bFYVPVyub3V+OZZeAZwBI2TYN2qE2eZtA/khqO3uJMANvfLxey07e
mXXXClbSrqEAZfYqcAjTBRqP48RI050U/7EcCYs9jaK5p6b+Xr0vnhcnSYrFuRE/
n7lMJXt7eCpnDozbSRrxxgT3k8sd1bEcsDcqKSrTDSK6AAd7GeA5zr5UAI89nsdm
aG+Ck6bPewPIneqYBt/eJfPHPhppWcB5NkfunPOQJ6w0y5yPMIHDhU6aZFI52IoM
nJ6QmK5dspsEd+hAOevIBiune/AJn0VjEUYhhOJ2MPvU05bx81O7Ivu8KUa5Ek09
1ZhRDI7H/X1CKERRriUMNXZb/aI6NLa6Qb40U1euDfHSr8U1kOnse87rq8ZT6V+V
/Naui7UdcDW7g7o5d8oMMmf44mq3UI0Fd1W+ZrbUq8fwfeuSV6WvSs4HdRc790iQ
xph33SA2QXVCy5Xb6PEFTlB0rmTLkUA7y8aIipfxAQ+QePfyI8ar5dnKDgjM9TFJ
sxV88dGqmOnzMUUhDfFBaGLXVZN1l+9sS4Wlccz5DCeY+4j6h+f+1nE0xSL4JzPv
eOFKrOuUG1fwj/9CjV2koEeuQZvEYQym4fI/2QAnDHgZOoFV7agqaVLigKWWvvJQ
Y5s8wogzAoFnYelFOzpo4XQQBqxnvaYTOFsLffkvI9gW0YB7kCx6YdelMGr5CiXM
hGRa0fzTnyMlISGY8m3+WfRllM3cmS++canmUDDKeYz2Rh2Vw8BEMZKbDVW7OqPK
VFbi+2Qz8/fNQAB1qsM82H5IF+5WV6l+cfVV2JJ+aNiJzfwmq7lV85JNTb6+VG3C
HOMQZRq0cx7lq/I2IVLUXvL6yOSHqCFhDylrqZESvVZUCzJ+IoKowDhSYjfp/1vk
ndphobig1aQtN720HbQ7CyLACFasodY9Fl3e+QjdYX2VVT0nq3Ucg/xf9f8uMh2a
uOg5eD62lrEpgkD/kFSQHhEMByaVIA4J+TtZHLC5z15l/nxhj0JqT6wIcmqqyV9d
59oE2u1GN/5KAMWTr4g87DYCH3Hb8dxz9I8RxW8XN/1MrhwMSbz41tjOF3K7urv+
0Yt50vzykfK90qo75Q9r4lpXvyZwGxAb8ChkBSj+4ycnrzFZ6oiuTJBKfT+G0/2y
KW47M5mRB01AVLXqebNwYnnbSi+O5qYXXVQTmMlCYLb3IClxImQjV/zz9QMfIK8Z
saAdioTt9QDlwsHQSZ3oEoUWA5B5ZPBjBUo18rfOWf0AXLOa9OU9r7utQhF1o1Ao
ggm6eRyQsxQ81EioBTZtuonYMsMMwQQ/ocHjSQ3yHH+/GDiBppU99bEYH3htY9Ru
SSoJ30fY1wzTyPCGhZstbq+yXZM5s0nWMKXqAJIYz27OrVsdVof65UaEFvX/tSFj
vulmEauEEs0Kn+WMbIvn4nZZ5pXJWN46moc9HlFuUtAhDDPgcQxrBVGyAG6RI1Ht
phu/MNoUnsq16K9cZNlm7tTieEb7bo07XazJlb0DmjNmg/yJ7uRQmySPctcMldw7
k1j0zXeDUvg8jJt3Rkso1/mlKF7AYxizP0j9g/DWIxEoN61g04mGMEF+s+UkJQxx
gP1OW3DVDwX41Mhqr2oa8WX9b7t6MSwc+NAaebQfR7iOx94Djjvu0V0FaziYu1Ui
ESX5DCzZFF1PrqTw32UY0krehCQf+P8OZbJSE6bfYTDVlovUeJrdPLEecOz+608s
irYCTh0ganP0iJskfxNZfJ0nBTL1UOTHko8u0ubHaNTZtqNJRRmz+8VAnTHGbpZN
4/sL2r5epZMeFhe7XZg5cdc2RfOevTdT7wMb/iLO9fZWFcBmcLPhxkY0WEsnBZ9+
wkVx1pXO5DAYiEamGFC+jm1jCPuWPl1lVMgiGnxaebrpCViHomRIUxoUD5AbbSci
3fSLPTVpHsXT1mqbO/2YQWqAo29vMAglOuA0GFyqQwKtuw6hsEy41WViBrxMM3H3
ebIvZ+jisqepplL1rUigCUA6ieDqHnFH5PcmeqLcXDZdrguXVMYIWrwrNr66JNPK
gexFVcY+Bv1xe/bHFISXlG8W9DLTLbmFiLXJhbCYszAtdQBN/4VH/cT+4Chk7slp
sY/lwlhwkduQu8VWz0g3Pa0t7+vUFXe1EhdfEw+j/kM5JUw4LgF/+Z8RVRsM0yY9
hrMDvnyNvn4kKZLgIOez+QK2f1vdPiq+xVHLNqk2Wc8fgmvjnxBhrp2OUdREuUmc
i6O00IhKySgU+Kg9ZB3NUbKJ63t9bRgo9pCjBi0x4jS2U04J+NHYyO9CH5HAuSKq
XmKrg3DOaSlxzgyLdNlQNlu6ApTOBseQtUrBiv1Tue5wXsMVy+6t8tYc4qB6gQKc
0/G7DVzvPqxqfa9X6fPY0zmjfLDUHHBQxYeXYDjBK3lz3hn0+o/RqMusr9/00Znz
w8wT3C+wJzteMA6o69QepIyMnMRXdTkUmd3flW1Yx3s88X+QH9c2nNjJHBroOi57
EsRP0xYSj/gGNjYNN/FE1ymbnoO2evQF2JUFymWdfD+CM42Nhhz9Fnd8EuPcWx9x
4C6utY75FnAFY7ukvVq+Wq43NIFPcaSQzxB+FTMcHfPK4/nVUjWJjRP+oV9Qjkwg
v/hLGksE2E/E6po97R0H+ibgvHYFx3V1G0iV7/JYkTBJdCFRMv6vSpPM9KY93QcF
cQCMcGsErpFRbxUIArDwkzcosTuszSgOR/7aB55SML+C73b9qZcVjX7/6QmMvbTN
VrV5gLgfkBmEoaFfrXQYLUC/DQraGZ7DKJY/Duh5yQIt2LWLNJI6Va0k105Y6TP3
W6d/oKQ2Q0xcGY1f+9b8xEYXNfUE+MX9dTfZrKfwY1Eb3UAO5nE+qUYg3/Gd35JX
XwEL4dPoNPHlzBzQTCF/AfpsO+r9/KfqC+Ror7ERjYPXP7b2T4tF8CFDF7Fsp+ZZ
GSef1BFBvJv3mnzQyZBRm9rgY0OPsU5oClhVPTD1f9tHq+QD2MU/rO5hQpzDq/nm
jma2IdqBCKmGnDUv+1oUSHFYN8wcO3a3EXwEfh9yf1ahwpTL59OYpBLM4U/29cOd
v66FoEXletzg+IhomUV1GLFzm9Vzamn3LQmd7quVKaZ24OXzojq7TQ4zzZiCWT3L
aQoC3adLPwpjZ/uC9oZHcAiPL6Ovuuxc8yxkTVBsrJt+wS+rXh5D1wHcIsZjsuZI
O/zaG/kyc6n6WlsyFiFM16+qAkbikTczkC6LASGeMWNWx8nQ5hH3XtqwOWAFt7GG
Bjio2sT1k8jpL8kxJ17qZdrxSXrE0io+m9hC2CJWPTYoXGMJCafd32Do10h50HXZ
jjK0Gr/gMlM9XRHv2IX1nYFiiOzB2PAOfECAsjIkiUdCa+dIFbvcCLsYjdSSywqO
ngJSYOSDDQyhZONyPpQCHmsqVEuqFAmNpNQX1MKkx0aySAO2BMG31socMVBsddY9
LzxTzSrJCL9at5i1W6zBEa2YPCrgY4HWPSjlm646vaGMEwRPQ5UBIQnegxE40Tt+
Xh6u60oc2jksPHtxTYoMbLeb/ICgg4XWcxv/L7hmrcvovUAnC/OeLRLtfKa7QnBH
wIKlBCcdevdi9fnkMj5NMdssh7ifN3NS0pERgcVKKAjsNJ+z7cjLXOJy0FgJc8Xj
5GeB0BGUlg6bNsiGcT2pnKIckRo6VDROMMbZTfjUxUShrewBf3wWq8cPt2k9Uyfg
HlzMUndlHjAhETonf6YeLkbyeGemYRgkHkFd6k3nsSd1N/HQ1dFF88oKzhFlHCpo
UGvtZaw9yk8jQKuBilPCbc6K0BdaqdB1oZdbIwkDxdC/vTcWMQkLCnGJ/U8GSbo+
D8rZrmpUbG3KR8Zk5rtW15hLAnZ28LLnyg08IEnuSKJYVmTPSGR4zbjuQzKeiThF
XAv29aDno6I2asGzBkzQKh0Zxnd1Ey3BxAbjx7LEdS3k8Rocx/JEPxtqlMjRvdht
NCLoNCVj49H+mItKzxlMh/z3WH0et0iSZyQJINIKYf5s1lD86tRGpmaV5nDuEYXc
u89UFq9y+KhFeglzQkmTDoquoxpHrYlRJwkV4MPeJNHH/fFxBTH7GwazTSr0+55A
KMNHzPitr1XG3nrpiFMJn8zvj1qA5L+EpmBTWYdLEemSgXOdkLWRDzsAKWrgs82b
d+oVgnarlmBtzxesd9OB4qa/XRKdro5H3lFONlwBApujTFUgelHvR/mFMiB/8C1C
pHeSAQIeqny2TXSUd4bClajAPrLyOPrHDSk9CwzimjCGjgxRHGtacV7eihbzlCTR
aGDmxFt/zDVtuIX+J84b8fk3vNseer8KoVxlgSdwPO5hES9momTqvoOXv/51Gkfu
55V4921+LJMQA8UZbxXaoxFGYRXapebGTd5zCG/S04cjZp4mzu2MmO84v7ibDrcJ
XSbwJs+IMpq7HiMrL4VjHE3nS30mNddzBRm9/Xh4p9Udy30iByM/gB2ZhTcI1Rpz
38edQ+J8crQ18qDkd4NlKkNvoARiGSqjZpFDHCckwMIQ6VDkLLE0Pv5wHwZLZsEV
WknyJLa00Tl9Y9fElpQtg/3gtfY8/6YxqTWjGYS+eY3gA6o/bCYOAsk8/XHsnRCM
EwJvTwFmcYRWIsi6T3a6y8BAOrT0emaTK37A0MEOWQQGZ9CHqdGn3DcREUzROnIP
arQ3P5LCbMzHTvRD31E/KAqng3VZvGtj7Psc2b6XhAqQL2DNNei9fnsDoZN0Ngd+
9K4XQg1sqRrw+5yGZyRrhwaiRRt2+EdXJ2NcdrWtIIh5sgt4P38tk7yYKfzzLt7v
ymzaSnaC8Seo3h4nlCuzis/Z22OvYo2C2E5cC4vWLp7ur7tsT+wX7Og9orCKCxIm
per4MBJCMWCG5/DOVbM0B1S9W4k/Gn+ZP0Ko+2wIFIYwtRhwlO3TTwtJHFbWHNpP
k7+eap3tvrCMhFnz/p0u0tLo6vqFJSYJZt2sGv/E7fR+gVcwcK2HyS41Hl7eudTw
B+pVCfJr2uMjIu9Ac7+DqNLyZPYYhTK4up4EmCZmd+ojN38GaaJpSllRehTaHyYw
91ou+QDDg9zVjx6jxdf0wBZhwUF7QTAaXn/xZITHW9Jr4TjvKK+8BmCN/mHt3n5Y
r9srjoqzYdCKIXMhxHJh6/ifBj1V+sQL9KXk2W9Q51CX7NrT7I7jdFFyt7MU8F/2
PMvP5TquCXNcw774Fw5HQeoY6oQ9dMU6GR1Xe1fFo/fzlWfCqnVnDHo7C/JDB0xY
WmCJM2pdi5TUaU206WN9xBklQOrtGZaDm9yPAKXd/bq1TORIEsJ+YTm7t/h6SjtD
vCbdNdkaa09+pNTXWQpsRr79oqjo6CWWE0HXxamwIf0gwO0ak78YEFfh1/yzU0o/
LqO4naK9vbcuOaH1fkMYaWrB2ze940Nq/t3puYqhiFDukD3xBrm7G4p2yN61aUSs
5dMUGiipRIt/KCvymglWDAwToD04WOUT/NS+S60v+hw/vXXhhYOD6Cq4rU7F99Ww
Qbg/w8Cki3oY8JEuVlMTQi+qvSmvuIo3qIB9e0aPmhBZYGkEuHqeCehL0Z8NGApk
cMunAey7DgssM2ijuWuJa7WAQVmluFduTcS6hxtv9OSNjE8pceIlIrM4eG5Z2cdn
lp544SeWTtW8wSlHhQtAIh7a+ttNiQfD40PgTejesuxsM1jkMFgRPPvTciT2mbw6
CBiELoWBMgr/ZDzMJfiBdGWhpI1v+HwhQQKlERX/z/TN9ltH/g6ySxXZphhvZF99
wJrjgfsCobMEj7qYlzXyvCkUcxUMf6aBaiQWoWNrIy5NtNlou+dA2Q8HOWo+sRaZ
DZM6+6NapnJYDJ+rqQDdH4QeQWYXfBcdo5GvXBJB5SyniBZdIg2mxJ2rTaXoSgpr
2vE8GW52GZzy+GXPuP91PYOnly/66s8yWBbZm3iIec0iK4j2auI3GNqOsb1bvxdH
DtYloEz4NDaa3DVKPQRURIV1qzYOmcsG3YBRQ8U+UNutGbv73pX1bJnFN34JrQxW
L8FWA8glugXAsTAhLiKMf4/7MfNo5AwOAuOsdwbelxKolDBEeAF4W/DkNpGP9TtZ
7ykkU6LNs91jOxIsb9uXKGJJQIW/D9l36Ho3ze0gxIbUxEj/yZDfTcpzFfv1IpGo
WobOgcgiKVGemJ0AcGV9SMDq4OVSLvmh/7DvXtjuxZgeTDZpe6AT7+t7E2zQw6Zm
h9gaX3cd6DWR93mBLLKZ2BLo42UyCoWY6ahdlIk0egj+WBVTnLiauQT6b7bia/0D
IzjArahv3ulAIWxg2MGeHa8a9wV3ApiCXDpv4xh/H5BaBy+kSuj11Q9Z45iHxQmt
JMdxwmA1MXmno8CHxpfkW4cIguBy8oGTphtT2h10ornS372/ZHEz7fORbVd2JmZu
RiBdD0p+izoBzQMWd1+dTm0YFxXUzIwTGIQNIb09m/+ZvWZnygUs+L1vs+cQD4KD
gofIgIwOQjTR8/NrwtkaBNkw47wLPqxbfNdXC6zrNQ+c5ppk/Ysdib0gRp80DFQ/
UCqTt6fYE6lJmS4W67QLzliwQ5y+priGs+qdCCh3I/lcJBvim0A1mAHwNw5RmJZj
Jewxs8XbUELuFWCTZgEiBFTZ7/i9iuH4D3KATJd3J8PLRcflZuwGtsa7LN9VCGdH
Op7Ce5Q746+p7cWQInrcdbQMncu1wbzm/h0V+KsDcUNhC+EJSQMvhUzxqUwdOuWK
FhLbFbaZTn0lIe0BGZ0UcgdJQOo3I31lbKbboCj68ZizilFUF7C9hBAUQljAANjH
0VZ2b35u84fDKUy7uU+J1vufsWHZGyciRktaXQr/a3aWHkF2vKuua6UxSEQnCb1L
qB4gnUc9AJNp0U39DkPaoaG+JpKldR31BNs17+0WPew7gUuoH2ySBZRFiPu69jOP
TIogkNE2iRxRJGJKiGdgV7an5BrhznUoq/baQgtLnEvMHWdXFQo3jtw5K7KxRZxZ
FoiDSHeSAYheMlAINz74sNnLRj/S8P4vXBheyT4Lu96zkkqJj0kfoPljbSUwDu/7
9uevBUt0/oxsTktsYbRgM3OHiazrZXK09bntXgbu1JXI/ahR8tPzbWcxswLR65o3
eyhMOb+Fdsut0SU+/C7YS40SQIPQWmo4aOZBx395pVJfgQt4j6Hcqh/+kOAC+lp2
d1tKtLEHbpqQoMshpC0p1voWez796M1S301zVzUSXQ3cPiRZ/E9NU9iah/6JpqGV
H30ctTjmpWhPXCYxagZNlh1HaZwQgUBt2DlJF3AH4F/peOFMhttD1E1ZzMhwcjpp
K9vO720+eVu+D4AuDRQuDppRdlzQpdoRMPdoUUIodmDWoVHjfipWns3dewlG85zW
l1YXL4h5nVzUVeGdmK/8lwSxdhyyvW+2aEhWYykWne/id7i1oj5LfO0iJDi92JMO
mJeYswMgnMMvbJxZwscQoK84vEUhViZJuDua1/HKSoaQ8zRItU/Rt7GDPVGd0nfO
dpVrdt9ML/09vFBCOuY0KMxzH/rFrD2wZunRkukmUhtfxrOXmab3aCkWl2WAtCtp
LoMZgoiykDtamR9hiwiwoBCtUkCtAwZQBypsmyfhXAdT5ukjxmeu3wUvpRQMUTs3
WV0ERwW6hRVY88Mx2GER2ar+2VyycIheAdEMxZN16JugD4Z23SRKsYjx/IUQbpjs
20u+zsSkAQ5papLSgHGv9T0mdajZrzPViePWwUgSKvCQHm84khkYXsbvNL+mPF2T
pNofMIf/DV1cy55X51orx2gfjwQuXY55uQHL7+4HnMFb8JcDTxnsr7GT5Ldstw0l
3lLfrx9GeTdIjgz203vlDwipy5kT8xMbHnMm7Ip6uphtxxPAWBdgf4fQxUyKkgVz
ntXaKJgvLEjY6tOII7eIPnkHXVOWe4fr6m+nKcC/q5tdm4BJ0UpghrKq1ALfDSdH
/6dkxyB9h7md3GMFg3FFkaMrhMtZT5VEJY5FYOWyvt5F7jW8lzSLQVBPTjemZUqj
oXjrNCOFyUqUFnXyECbL9efLFBDd/H2D+6gt1yo7JkMqFesxBIDTFIJHgFpDSIjB
ZRJ8QCTyMAckOwrAIWaOYQkTXf83dBvA9A15g0ysXmOEnFA+NoxS6hnL3pp4CSd6
Y+L/uUel9ilcJ95xlRFDJG1v3OqpocQTIeDEku8oZq20hoSBItD9Ri3wQ2grLjQE
/kduqBv7jarFrFbL+M5iCsNrkZLSMwTVJv8DcCTrRjA0IF+BmIU+FU6usGoLl49h
ANCP33QkS7aMqsYH09lGEMem5T7mqova1+chKFfcxNX8ZinmwX64rLjTc5I3BPXU
ZQUFWDsEVOEHeWeA3dFlQF98hj8Xa2fa+VwTCOcgwIhoKut6K6KUVv8G4b5a8GC8
Z/mCxaT7eYGSI0fFJYzFgDvWdarYAnBgtBB+eEcspY4Hmb1JS+gbbS9VDy1pCDwC
YoDlkpOmI29qG+eRKxMHdt1mWCX3VFXDveqWo24vu9RZEcRMExs13dcoCKhFvSWq
nbWK3cCdCQscOUR0GdMd0EmmrttCWkGOG61ysEcVyycrD1/htFHQI1tmO1lU8M5y
7tRWHK+w2FHSTD58QM5ntvSOTL+Z9orvFxap91a6i+D+LMtSsyjf6D2CEQQdHJ0B
LaiE1x6rNwJ3c/tBoKAy68l95xAjCAoZJeNfjQ8joLCHmOuorszyJEyzcPhPEpyu
AOfQuHloYbkuIMP5588+W5tdVZVT8WjtQkYHnWaBpNEgepXK/naYW80e138NHRAa
oNQzJaTweUUbg/QrGBhMh5JJhAS94uVBE3kXQnf6d9t8Xq3WQ4i8XqNHUM8+L3pw
wTiHrdH3u/G2nzXsg/6qIqu2pDcNYgJzjMwBy13r6leBYmuUCqNqSvpY39tsgTK4
56DmcgQr3tav1lkf+lAr1RgPdzouqQi+BslDw1h7LwZtY3NwZywlEMGNmLfjetR3
uQYxTr97c9b9memTe60U8dI5qh0ENoTqt2U1BEL2+ub6eMNji+70EAt1lPR5RnKm
wZtgrZTNX4A8MndMFvNxRRdMXrk7jy8zWQD4WPMQoLAVYWu3KW1q3/UgC+Twb+Hr
BJsdBHvLQAHDNyiO4kLjSBj0kMGKQ2Q8uOUImuh5LEK820ZhAkkhVhKSQEoc16wB
jhP+wmx+XbqkZi2RBc1WDFB8VzHQTqGSYHWocIFTj83SEom/efGGUB2D1JC3qvWs
gPKL/AD3sXW0bCQDIFTpbFbU6Exdwav0p+kV8YxWYlSbZYs39kTygtUewyr/1xtz
Sitr2KjI+PwWjFzLuGQfRgWLx5qsp70rELXjNZ5wHhvctTIQ1XhEcTXq5aXc6nU0
jynL0lk5oaknNEBGlWW2BY4aaClnXBgFYaP2wpool6+2OVw7athCNYGFvaC51Dat
jGZtKbRz4z8GqUdOOccnku0jv6LKqi921bwM+LK/t8BVEnc6/4E1lPT5uf/5DEzd
W9xr9VVmDfdtcpTjPj+OK83R1CfbKoJjQLUU6Ay08WAGuAbQSrM1dq2WFakpFE5n
DIVKu5XYANzLYtECJ7RcAq34ODtyMujkrSZD6dtgSHOivQPb57XtXv9OJg39BEAK
WLNm8ASY2OzdfPgPLf74Mk+7fm7p+sNP2HTkQZ/cgg3fJDds/XJLggbaz7RoYVBE
zW02CfcCI9yDTTqgx5tsWZ6T+EAqNJbLluRZnskLpFlMXDt9ZdYeQ9k+H7P/sN7e
8Y4Iz+Rw6OBgTgKrHsOfAUpg/F6JtKCwVitN/gPgiMCwPwoz1JBU4YnyR8NQZOvT
MEPSIYOcklVauxbEJSst9neJ4yKo8k63GL50j3r5FVluZHX8gyC+5cGM4STG3FQd
JhA6b2n34Sq//13eV5Q9hxShGcGJWURRnwsfqrXOeMr3F4H5Pts9l8WCQXnDhYh6
VpSez9MrcouowRc3YHqd/F23Ei5HZ6slbX1iudNuzfmDxB4WlaetoT445fM8ALKs
ekqtFjnBTtLB0piCVUa0EvSUAoBG92RAtCSD/22vvmOzSGFaVLjZErGrq55/cI1g
OgXOG/JFBh86FVrizOszGoPbHgI8dRixJNccE48oXyPOR4yNdPIfv3yhOgFFKWVQ
1uxnlxmMgV+AtglNf5p4iF11NfCwCR2DPzfwYik5KV3D42vPITeBkSWMJsHkwDmW
jRIOsD04gaBYTDVoppMLTundZiB6uSiAwnSPlCM25md1IJN5ROtjq5mKseTwPDha
kzNJwV7774wqsRJf+U8HYTxS8v9cYczXs4n2RF5H+sqO+LRGZPj+8l5KflrpKjmo
fWSSpiLn2QYNoht1pdVP+VQhpiYQIrnqyL/W8VMLU1T24AUo/dc9bYzbL+CiPITr
8PLpMk3zwD6P5y1r6t9zR/yOYJA/qZGDzq3XaDLLtlpqsjMVhS755Z8YxmviEw5z
A+P4oA26LhKCxDr1mLoXSGoka8BOqzd/Puw/LQF6R8rlPQjp7Q9sg7TbMRwkc+Ie
vF4pZIS3jAun5tpwXHMiTtu/IKHybz0PdfkaXulh/uGl98KBzj/Bbg9eFNVpIa2u
noVCDxYsgOcTio0gSqEKur7nkjnc/9C1gson4QpaDAnReo6S6G/2wBkCAF73qXng
sYAQ1VBjm9xz/kvAM5iwbsyDEI5/v8G2E1/zFRAIIhoYvwO1sh0SUnyKZEsGrHYD
/uTLPlLzr/KqYF1oHtVT0/P8MFVhS3MGbVsMQCI6jLT8GvxFml5XvW7hCvwRvlQW
h3w5C82q3mRoEnRHUSEsF4Vs0brkZn8TPM7Um2gT1FYL9k2tAQQfLXPgpMP24KO+
yJJ16Jj4BRZArtapDkeJblvCTPurHbg9qmRVvIbmuad7Tt6WRTpixVWow1kyNu+p
txLg3whYqwqNGomWjR/t78HO0sXMaYmcdMt+tvtQNiSU+nS3Emfp3YzRyts2Uokh
pnlgitxR3VTOlq9va9aCUneHWHksYk9ybOezGbHPvulYe4yytxwbEahFAmcdSro/
rW34YGL1h99bRfazHXf6kH60Wmo1qloGlfLdK7rHX/F8O0xfhl1OGmNwkttECmG2
PLt6YDMKUcHnonWy39MKOZMi6SYuKHtdpu7acOIt2gfQSbNN4PWL7MTvj38jXFmx
eYj7goQk9NqJ4ufZ35BDRWjP1mLOlVtqw/hstXpPY3lA/YGBY9mEBLnBBe2/OPlF
GDLKWpKZDCo+4ZvSQ28Q9WzX+09Huusf8OCJEXzdoyvXVwURQBaqY6wwRPis3TxO
ZuhJYyYQU/t1MebEbeTYnaQhhCWlYaClqJ5iHRZAw4ihjXn8IzM7uOnfBDF1iY06
fHe+y8A++haZd8gpU1F8lxw06rB6NNEG185QezzkQfumugXBy3BgzrAO+axfFyZ6
R1wtnjzXPYPU2n4JOaJfCuMvsaROZCJ3INpvBA4X/7O8sv0IvJCtZu6HmYNf7VLb
Z/WaKcEwHSukNnnFk4Jx9nP6ZoRX/bpO5bJODW9fLC1oM7GVgnCvoEOBXSgbsmiC
kBiRLWQD2FZ2DCymX8BQo7mE/lOnppaTkqRffLhyJyPfRLJYoIbHmyiln0XbQlF8
cawgD9Io3YwbHqq0nS0GwAKl7XeOS5F+bes9VhBKlYrABJtmGaxmrcBJlXLQMmpG
N12GGp60eVCrOiuNhupwcXk4BJ2Zp4vfKLrLvrvrWkbvMn/Jgop/dSZLJkm/Tixs
LMIMYeeYFNqSaNwfLazNKwVcosS57QBARaqv5gy78D0mKfuY94P+OmzNBycy1WIH
oYloS4IydTfPdzxWa+mWgBcbxE1ZtjaURnxezENnR5H3ceNtgSg/Abe5KHh54bf+
RWxbyzFfaQjJOg/12YSShkwuxhCqiqPAtBEEuNp4He97jN6MJYjAdPT8V3g9O1kr
hfKFsgpod2vNuthi/Ydkrdt0XZ34xqQuwtKOUEJ9GQ2BgdByD/M177QQZNEz95xO
18saXd+3sseqO5YFE42qQ7OzFar88blo6SZHrPK9EGAr9s1oKvK3Y8Ftgt3uafua
bnqRct1/vzODgNUOga5APekUNEtmdjtk8Er3H2FgVCDpPwFGcOHBTmskdtDgsECE
NWYQhmSY7kEutzXq6zY+By0zr6qSyE1+C+6/JK56uqe69sC9EUI9tXesPFx7rV66
SgynSh4kz6wfNSdlI/h63eJp2d8qxQifqZUsRex2uopPhww52lmN2lrpDXzi4tiN
ER5rpR96pm/c0BeTZjFGDzl08fMDreqPv2dB2TmUJ7Ms5kZE4WMuzhmESOdZui0d
dH7yU2B9A247STmx+31Aa78wOnCucmksTnyXvdA5XObxq1CK+1/q3ORohkY/5hq9
RU0xFC+5ZxJeiEopYuPIN+yjUUDEJwXHw9qXh01RFABQoSNf/4a3T//GAZDooJI4
hR6tkfUMiDxgKPZlRZLSP632QTc9zWsVWhed9hsZ5KbKMkL47suPCUOP6fitl/4+
8u13f9qlcbArhw5aQD1butVYcPVMfIKihO7izuS+5XlbmXtI+fGj8d5D1GHjAzHh
jJnHIWsak9y72MkI+WIL7W5z19vGgyyKKY3S845Dalv3cCbn9SY12BFOtkqUKda/
KYYWYYJMFD0+T3cFiUgppi9Kxj4NMUIKS5xL/6VunBJE+ALN4E0lsG/R999LY7pB
5eJ34C3gKBjv2Yoc/WWH5MG2tcWxumc0JFjcZrze1A/1mnm8WMNKpjJDZ7EsBMSL
RzYTC4J3QVpWdsNXxZ0q3y8A+5OSxvA61ipGeJuZgfY2nnG021RnJIbLMR2NZ65s
fw+hwKo5bPbvpkX8DwpiZ/kUWety6IOouQPeLg9XA41thFZaSWaQ4XhrEkMmmLV7
MCr+y+XuePONSGuv55rH4uktg/vIrTInMiRIwa/r6Eo/0dHkiNOAB9P1EDFoZjY5
vI5pngyb7anhRfrqH33LUpLfUClwtztz/XNMfOre6E5sEZIGra/Qk8PV7SZNvwSJ
N7JV36b7UAN01vTpaQSmf66QKzlBNRHxAg0pSaOfqvBCshQfB/RAickouJhCKy2u
/PEyWmT5ZHz/7p0Ia4pcCwkdVCwXvSKyHRZnTfEvbQ7plnF8vBPliXvI9a6TZibp
HZzpkj6UmaPJ0iYWsa2pfzP0hyoH5MTVymgSBbL/sCc9rCKqNkf/b5TkCwTaPSeF
Lx5hTcPBOKDqOkLw3G5hm3Vql9DUjMLlsuz9wIInTufdnXwcK3VMFqnPJVbHk2im
JUy7KzVwPrbWo2etT6QMB+0o1RKgnZS1EqyCdVMobP3n3630clhDpFP+1PHgpd1G
d3gxbBFR9pDrfGVKmi1MFIujLuOT+EC/DtTPjVIhPKtjmc3j8Hp2CLC+xYyEVrnj
Dl1POF9VREzFPt5uFn9MNsdPSawhyGRglctH0zNdlg1fh4DqG9sjuNdMIWyqac2L
HD6rCMyYu8oRHpLT6wQ4amHgrCFStqhckCUqw0akSdmUc8yL/S6BG7Qe1OxUZD0r
QbuLRVc2tL84YS6upXkoq1KA3AyfLDRWIOuVrEcMDxbRzvsTm/xPzXDgP6vtAxXx
CdDtBSANSIJAdW2CQTjIX0XuzhklDXVrGAaVj8WtP3M0ujC6MKIiGAVmWHrMOy6y
/KRKUv2WlfvxkpuMlnMZlHwlKrqwBHkAMSh2Kb0C+8eK7ggvbL+jAZ8XOjOAdkWe
w5y2yyxUU7GCpAYjhJ3zTYxsKC8sqHbFgPMdNFwjSl384NJZQ9JqRY/ntuVGVJYA
6SdJV6ngq+6xix1BCgm3aN+6MLGfRi9mFEGYocVisED6rSN5g7ov6fTssYYcgzW6
0ApUVcysClZMOKB09S7BPgTF0snWPPdhJtFsExXZLlc2zOwqSx+L1v5y/VtIygyK
+51WL60/Fd6V+FyFEqkUJgXV2G7+5/kjpyKDafAZE8LhscVww0q8NKPmb+EiWfly
ND0Iabt9Tn4DetMFARVWeSWmcott7862e54mm/ULMTSahGgUcsWr98IqBjUtpLDc
O2j7PPnB8FrruLFeDYJqXrWY2LvCYhREdfBIKyk/eGnoCL7krM20wLis5qTCfMlN
vx8y8hJgSxOWoWKLwjVjMOhrJTWyh/1Niyzr+nUJvW07nvZucvrIYKzrzz2ssWlV
dBpN637BC165nCk7sUHEWThCNBAyBYpRNqTuoXbTPae8ScOVN8G8btpp/AKNqzUA
1+CN+d1QxIw1eEJ6tM7CCLKkJK2ZLCCfITVG5WtTTNluh2vD33lnNakZHXTUBsSO
pNG7YspMHXeQCxzGkWVTeUHKh7KCX3PfL4G9aIUlLdW9gZ0sVbt1kRbSVf4FOsLU
GyP/Kk3rdxLWgidTJTLsnnylQNPQFXlkdOyM562mOChzlzDYxFnMrQ4cDUANk1yT
x+nbcu2E/8V6pG8BWfnfHWefRYdEcbE30wZ+cr1mN6Hoc2V/ZPqjinSOP3Spe4gp
he/HcEWFEWX9IDH5IuTzsxATzSmTVqrYUQeVH3z2Zrman3PL29dyYH0zQ+46Q88C
QH2Yrk5LgH2BZrtqXW9fSlYwPl4aLevvsk/SWIsgbZnlu8KN7DyFOXoXuxp+5Qjn
Bm8O2JZXZmCFL1eClB7qoUExDbhwIO4kUrrnO36ApdcOshgE+HJHasbP5nLdJ1tg
IQlwZAnXTHX6KtgYFpTMOS7Tch/tx8GYtZVtEBgZ+LjFHgvM50gTGaNqxpAvsiTO
W1J10IFTWt0ABvLiTVLiDrpoK79uxe5cVLZvh9tjKiaPh9qAPjI+AH5ggHqsaV5A
cHwnQUfuR5ZyIC3qHvF5rTognGSmIGfmp6R/FsBQsiHl241O1c/ojTKhJ4R5rkJV
eKrGt0N3haZUkbBJulUis5wDUcsEwEdiCqJlkjjX7ZLlhWYh1dP7Sadn/tU7IfZH
leiwnHF6I978Ie6Ydon0Z3J/L0K9b/61zK+buHapkP2gkod7XWTs0NB/s/3LKqtG
lcw4Vo9MePeq/fcFR38LFAx/Vco1E+4QNZFV4DshNGJLK5VNDRlKCtImpruttGt+
nZJdQj6PEdQQWWTxltJ66OEYgIAGJQJkB+sHXZwNrK8IsYrWA1jnDs2LmAU4uxcn
AIoUIpA7xZEskbo6hSWgnfMiuhHKM2iznuDeBDCXtoKRXikrc3rCyIkQbpAgx/VF
4xVRqgFhK9pvNu1Ad8EblB675IoeFdeVwCB162kWtlgwb6xA6R2cNUwDjLmBhPOG
WCjltiv4YDhfEI9sWQgaDo1yeSdcfYZm7RVc0p5cQpxuFFGItZLryZJAtafoDiaW
GTRXkZMcHwiJ0+f2KvXaCIrvoYZ+ExdFHespN3L8Gi5wIi9V6JU7yIW33xg/gkOC
/y1LbPTCTUzF0PODxoYyDxtM6gF60XjBWyHMtjStYwHhpry0Vnue50BRU5jUtXKi
dRL9ppmnGIGXdQZDlvkyIKrnDy17FO1gLW2FWL4EMYOtHm689mkPhBqmnQ7SMbn1
trKD2MGyolf3DpfpMhpotSRVlMi6BbS9hImX8kBFq8UrI9g/sd/MvxClX/+p++X5
YNIYyoIcPxesZcg8RsScAem1R1mhr5t8M6WQBqzFRZRWXXZvBZJcgJisZFal6IzS
EPmr8Isank4eeX3Kvpt0xSJmvSSsZ83tdAcZim36nXDZitdlwlaQBCn6c4E7O3Gn
njDJXI2KsCU1cPVC/yRrxOVJuBkCMd04uNXn4neYuAsSxovyLezK1PReTTYMNOzk
FNUjLAQ8uYywfJskUcEXNhMVbdS7ktFR6C0DN6ejA6X+Rh+2mdlrrXNE0YHFYMDA
3k652QcOtyY2wUqcW7ylsr3Shd2tV4L7OrI6TrfnTiIutDCUIbQytNzuck6TRWS0
lab25SDcV/W+rhpwfTKtrOu+5IqPqy7+nhhMYl75gKSj/yuDOyMcT7rbrwHN7UsH
bnJ/YyADkejSLL4y6NlbW6J1DsHRW1behIp0j/84J34xyB1ATZhW/pQHr1tGWfQy
nM+LL+bFQIT/21fQkvXsPLSn0PHIZ1QDwNSJ65BENgNRaAwrOhvq49ZIDmE4lhJ6
D6EL+klk2C7dwIy7GaMzxlw6fOUfEg7feMK9Q3/beKv+F0c0xw/MqeEXuI7LctxO
3md9fG/XxLkS5BRegiskBncQClpDQvVLVI3MZXfivrG44GlLU2zMRbimIAoYDr4j
+GvKx7AUClplTLIyjYtKquY1GGprl/h6qSnbsRth6Nd8FbwXEhz+scxsI3xLt856
B9jgv3EdY+5g0amzuGmepQZt74wRY98O/SBxl1M+TtXcIvanIfmPdpS2hgbw6088
e0lW8vRV/ITExHrh3OM6TpBQ4W31mA7Te01/ea49/oMmZiOD16MLyfD+v1RJJgsN
Ddtfgm+YD3sa57YXAGtmwdlyHfwVFdlQQg7ZAX6/NGq/uhmTsmET3ZEq+ZZcsoFG
j9QOkW4uChYtXmwLXnM7E3OLCAIqkDJu3BhCTnMJfqh33HMSnEAS0N75UGDW5Gdq
MV0TZYkml6MPhQJrnPrn0PY+MgQdyH+2UYQTaA3CZtpOYY81MYtrZ0xW8ufQURr1
MkIsoZXhtOmBp2Xgu+wgQilTqOpEcafWy+RFdFuDNdANO2d7KSbzFue2MkkjVmk8
hzDQeAoL5uD/RLTemjU9vr0TJ0HlO+AEC+NdCsqmwXXEF5MGWbQWmnwKfYAcbkAG
u5i28kE4xbaZBI0jyHuc6H2iFiHtMUn8IqXVPOYw7fXoRqe/47tCIn+854yPResX
F5S5BaKVHglnEbojhPWeJWMs5sZMCKsd1VXKXsEOrn5qJm6BiIK0+uvOgSGBbwIg
/AcZRqLY9Z710FGHWBKsMiECtbP4CuGUqkdbDDCUpw9qUCvjfEpgfzpqz5hPwAvl
BBiEoCvBYoP+I4+HzhXsKqgtDj0eS5dRL9iLYY/xfmg/fUHJi9h+n04+EJ23HCIL
v9UXy78nQinr8qh8ED5MncVX+6Di0lr0psc2s/NwK6emFgbWv3xRH5zr0PxPf8Vl
Ndf1ZNtLPbXGXECA9stmOUJ8c2Ge7UBVqxCmch8lwc/LFWLj4S/gAmQGaDt2Go38
3me+Q53uOC/t2nD/bE5vxjSDtR1mFZfJWKdJIg7E6AmmALDfzujbF0VrYKgibuyu
n8EVRAM51+5TVcdH9zBmTfaTxRpQ5V7OdArncgVBJGsNhsM0YAsOwRKdnCJOy1Vb
uiJDG33Ew9UGKO8GE9iIiWhCMrLrpdCNv0ElybpTDpT8YFTyh6wHYCgA7Ww/XI6Q
hFXrdkcxlhhR6flBk3gq+/HTra+j5EFFUfuXow3Fbxes0DFpQ/7Vi2QS8/w5q9oT
+gr74sAneZAJsSGlHx5tJWJsHpvm7FcUiNFChoXhdk8AaulC4jgIIVpfK4imgf3s
IxQyDGWHQMDbxC73AVEQoYQX9vnEUQUwGkQeqFVxb24SwtDuhypAz3DH6gnUvWfy
p41FEC4fxyTQVUm1LBFUGlqb7hHHy1M3COuhWya3idrcYxARv5/wuuC1BwVU/QGr
JsXSDYnHR32Uutn29BThOTkbviyg32y+J5V7PO720+sMQEun/LvmBqkvkm1bblCW
CvQogIS73R4vgq54gVl78cXSwhMebr8Xyt3sbwKE6tAri8SHk4K3KHdeVfCGy9KE
LBfP0Hy4GL0+hlL1XziqOGoYBB7m54YrMgREZ9H88CA/gaVC3YPXvVWK20MJqNEi
3eSt3TUP2v7AYQGZ19+tpomXrq3rBf7Ny3l4CG3gfhQp2mrhjQUPvWioI2uNbu0H
ZChMhWtNtpzBqEPzetXJjIrCOZsnF40LZ7eege1QeEdKdHsFV8LRidlpE5rcotrR
stRda7Trs/pITB2UiqL+vAf6AUujSUW3eq89vClJSwCpSehAifRUnCrtSsuKwATT
rZiUFZ+WLR3yZd8svRFQWbQkGGO98LMZBbCcYxAarhXcgpZFRyi/igN3JuX4a+13
3Y99iFUbDmAxU61L8ZewGf5lzTLYjqjDZcWlc/1tXUuKUS+d1/QbjhjIUdHnQ8Xk
IWBGjbF5OZZoogW5X14357W7VGB8lsPCJgWEvicZn68BOdxd41bLWB22WI8nFmt0
NSWELUvGWrqnXOjFFKO1Ikvw+pjgzh8O5qxrpQkKzaG8kxMPzSLtnyndfb/C9Nhl
RGV+e00zYOdRKKmEETYMlYqu8NxSXoo3OQP5GKcdk6KDmdlmNflhW3Yj4L/fLcab
ihyZ8pZNzGN0uMIQmRLcgq1RCXKZv2+hpTtBp1F9i/oHqRCsHrVgZwC7hVjbFQYA
iW8JToAdZjo5o8uhnpVx1kySnzypF4pym+n+SOxzQdkcbGEM6AjHaV2Hp4msWKfM
fJGlrHTYYGZ/83KLs6lt5jsdtYHV34aiu9RoAH9Pk8E1gOLFPF7KakE/Kreo70IZ
RlIxz+O2i620r0bbYIunHugQtL7ynoM/eCzxEqp4ufbve4CBlqI49UroCYEMUSV+
85ZoTKz/OnDP3PFqXNV/AO4fS9+me6AJLbsdAFNIsJnaqIFzIqGDqSsYxKfvTJYP
KcqhSF80UIXy+67gGIQFKHJ3zoL/Znp2tqPxeOVpiSMO5ogliHwRKO8vcmJT642r
O1DKatwD2tu3TeM1TNFBEQ5AilxfNhUJoktTSPxncqg/8Bgb3J2rkVkrWF6QmcQA
loko2IuiBAoWqf29bjlIcxs/GhhHAk365naAGZA7ZZ/Z6Txt9Jf16MMAAE0HscW7
t62ssaiEA8bF7aKmwp7uxiZkIe/ECHY0iS2KAL/IoJ1RoG9hlTsuZpNcUj75iB7Y
8X2eqYb43twX2ekvneWcm8+GPBNnlzaI+zWm+WTUnsSlwgwCxWuSLAL2DJiR/CGG
KxoU/+uac6qKCoe9hl2bsb5WveMWGCYFWODgfzWeiF6dRYGteoKu1gcBcyjaPthZ
9DUoIcUFLDdNxCPLp/79xMtzxNyHqiiKoZwlrvKGLo8CWwdn1oO4ZDQaSWYQeVc3
WHcExKXLQfHmRIc7Vi/z7YZ3zBCc2VPMbQcGNURFDdo3+lmJzznmaTzm9k4yC5M/
dnDMaG5DfEM5Rx0/lE03YZBOwLsGe0FJ4rjAdwBKBhjMJSKsBoQQt7uCPlQb7tvR
me2hho2Z14oSOaAJDF95tlKR2gkkgQHl6t2W+CTzi2+URIx8MdAH3JX/I1nJspsb
cy7jR22ymrQiEB8M82ZyQ0COIjb5HzsI2eLV2Is6rDmbSpziOpoX6suzTDoQSttZ
Nya1NOmz00Covo0sIKS/KcGZWwRf3OzDl4krPpVg/XsothpcTzgvmmR1cE6PvWK7
DF3xJF2k/jg46Agw7chX78nQgZba9Xx/CmHFwkUaMKqiBuZ5x63TB7FYD9qRRK78
gFtZoyrKtBXWOKWCpEPAUoO/eulGiPfUMuy/8ehJSC83qQ3IAPhGS/YTJt8Tjwjp
Sckhh0u741zvApQMcto+VQvGhMVfQlQi5XZx1mcnYUDvyBkw/mnLk8EUyWxmj2u+
/OnMH+LTn7IXJq0Xj4zWaTSlOLZ97dDo2pL3csCAu32XNE3Ifo4Cci4IMxRm3uY+
2HWTPbmByQzs9UQKdP0LljQl2tWAutTnIXsniTZIg1wyzteYDQFalQPetMeGpVH4
z9S1uwz4bazIH8+DDG3AJla849etvtS4EjFaglSO2Dc9SGykqy5x0uvWOHG1I6Ca
6tCLd1GBDX0O2LCGZCdT4QMqd2FuDqKnVVEnrV+ad5DttnTary2KtdF4OzToe2c9
7NBDL9PXUiOcVoSEUPP+FFWwdaGQBtDX0dAKCmYUJG4M1fiUScqTiGZh+ZWjLVu7
luPxebitNbEbSt+nUJBOW2uVVuRDwkuc0Aw8HJZBqNK9Me7m6+9o97uAN2Bpwu+D
+kHHNbCh2Qnn0W2Ir9PeUXIfCV9VmwcPwO6RpoplhE4txvcFd2RbQbpNQBNFynqs
N6YUPHUJC8ysdku7RGORKfzCIfuyr+2D/NJ/S7nfazzhxZZ9G3liPXrRYUNjr56q
Lu4Y1o+T3zN7O7Wgu5t4Q8heZ3B9N9BQsDInBwUBMazBqFGGN9OOJbVhIQOFmoiY
fTyI6LHyWOX/8FwwtqC8tD03MKIkavbypbosmToTwxSj9aWEgjUiydLGGbOxCbdA
607uCqSCluOqMTRv1N9PzAoTmeNLmk/Re088i8qwJgbD79I03SEbmY5auPGvLi3s
n+CZ+Zcza6Bhycp59wksYlVpz//tEX5gW922kIlIk3aqas1w9NUaekCJnzOjMBk5
MzZiHEPtHBO4CsLDWfKm+C21+l4jBouxdnNfgjX8xCyQZS70+PKUEWWYR3jRX6VW
S5HR6SxFUG4Bhc9Zj79n7QYYoitDT5s3sOzR6R+7Wnd2Y+OdmhxGhoVdTDwMiXRp
SPM7G/IkGGNLqNQqhLnpk9iqxfsPRvn4zyDGkZiA6At9MWB0LRWVatP7Q/ngo0cc
3W+Kx8tMMiAQg82J+vPQMIXh4FN8qxgJSP7wF9lM4b9V1m/jBpOSMZFosd5+AAaM
4w2MfB5LGLlfmjhcZg0lWi9ZA1GMyFaEOx0P8tOK+PieyBBO1gS9hbutP4nPSurU
GKTOWKPzEQDPbsMPKQcfuLCTr7E5Ymg4eRw+O/RrDwYAU6Ps/ZMhwvFV1cFiSnfx
jLYRF+2QdDvgCTfQbvjG+K09VQegBStUWpBTXSaaiInmLbtfh/5ruk59YFahbf4Q
Xn9rQyqLhhIP82wa31pQGa6sk+wSzVZiaqs0fHFuiCK2t2rlF1UX4hz6xLq1hQvk
wZz/VaIntal2x52O+oUK8ykk5+2s0wEoyUrs1035FXAjq2ZyBH5JC2pLP22g0FA1
S5Qx6tkXXU8fKv6hcWol0Mxfo20pTn8Q3A5gwGBixlLq1zSybm/g9fZOsWrgFsJt
Nb6kLy0pj+os7QRfEyPEeX9yxaRaJfMcUuwdqd8d3ScQwXKipdBY0DzDX5qmDQhI
cKqfdUIQvWw4q8a3hwYy+wYwx6Ij4lpV7KRkdF0owVL9vEQs+QFHftiErs57ws+b
JI8lVNDzsh7V5Gyf9S4K1Ib+hXTCM+rmoMR2uVX+4kP449wklJ1nxVHrLIp4i4g0
13GKtvKhHPHrSCPXyPaYd/dWVF0MnQ6knw1Q4CUTjZ06Ql62iy9jNUXf9emMOjRg
kGINT+HRp0HES+eu+gM0fgpgPIdeqil056LBQfpcaujOglaeYEPjYe7lCfTHbhls
/L6IauTGn+AjdTVOk9Zph5mznBOjmBVxVIdzIaCJFCnNKTYiBNQ3KCYtRJTkJzds
KpqFeWgxE+FlumGcNA/i6j+VC18VtlDSPzif8WcKXa6aFYUYqfGOiz1hDt6tk3uR
wS1y2wsFuetN02MLpjeQF9/O2yqmSTK3+anIojMJZSRMnSWMQIN93Oi2dwB64/sN
GthaomchaBc1MxZNUwjWXFAYhpteGgNYoTj9xgz3KEWniM2oZGOa6UCLc+LiCO4h
wB2btKL5SVSj9lo9/cWsQztPL55WBwkKJvOI19EygvWr1JCpYQm/dgtjVD5i9j8I
ntJUtiUAmOyYSN+AH8XDMM1USjoiayugLtBYUrlYSikLP2HwAj4W/toYcLIeEz24
Nhz9v4vw1K6Wq42OGN/njvv+xelHcdKsrD2mxeoBKpJxDWQmtSlPScy1Z8UMrQZw
jA3l0yYELk0Vr1An0ZJs80sps6a5o/TfCxPQ/xulVVo/vDN4J0FuPGwumqkH/RRw
/YNn0RFgbnpJmiz2u6z9ha545zSgrh4qOpXY4Xvg140zRxtkCFkcClLIyzrObC+5
xYjcXTdpQd2J9LGgmi6GBS+h81ILID7V1lajs0kXHnp5SKW9LAUdhcJsgGDEMwBq
OxZ+k3dM1Uiwhoya4AzjfZfGskXVN/KzjuTWFOWYpy9nrOgDl0Yhg1XWjIrKB0Qc
XF5Wpapvm6zCfh7HnTTENgdCDSxho6P5MeASSCuOzACX4b5kNCg+BOGw+RhOn2Ed
FjlPCn+4cF9baWu1uur4fdFqQUJRr1TMKn2CJ/+Ez8/QAW1mv7D0shjYw1W79JXw
O47njo7wTCClzEaPjL5RxU42aAP3hsQT1oRSjFDMuPPMM5s9oTD6mO+fY250ayWZ
QGSRj0lp4TnR3NXOLK8xLGdUZldhFiy9kIvXIGakiHR8NvMvTeYPmaIiB60uyfFx
FN9wWxBydE7j6dWmcdQfF1O5Ild39E54UY8q2xh+fT8ldHyC6FXPI9KIbdexgu0o
RBP8bB3uBcHkLMZ04Ri7bQ/f7taB8ma5THujPUcvR+Wabcc8wZDNGKATLvh+rCqS
+apbwynstYWziLx/Nw5O1V7GMOcbvWgdUpJ3dNNuYfvcbvALy+JQrbYGCwftYXWs
Qh/UjjJBXwz0If7Uz/DANxJKuT5vGEBxMAJ6TvZRHzJ1mZtH55wmJe+xHHJaYRkc
JiUcVI2dLXtOPvBCKybiXy+xiV0Zh7szzngu6ASCQOYHpXZnnFDhr9fHzqWXsWSb
FFG+gjMWQmWV6/Q0/Xk2Kefw/n8H+mS72ettoujH8fEuc+Cwu2AIB8+xjR+kiOfp
TsfNuE+t9KM0CZRkHRqNoQ+bj8Hv/9wUXGx99DpXDK5SJEZUPIIHdAD5vKQGwwag
GOfJiirUaqut9UW8ugQce59LjoQab3O7/RukDwrSJk5yifTYVEWVVXemC0o95UVR
tu2H9d8urWcOayZ8nISDhouY0MInxbwOJilOjknhMgVZlL2T1bFQiJb4pUfgRTBw
qTZKTJoAL4kJ3KKfWBZz32dfRbNQkj/fvEdWqTVcBK0oO/Xeob4NOc8Gr+J8tctm
ehlVT5H3fvnkl8njcsqfB1ezlO/3HaATLwxwy04c94nHBeAZPE/bvs45YCosaffo
kGwb57uxlkw9R2e5k9b0demWIHk6ITX2zx8lKPNMeIPhpAQ6z5dxIzlGnCj++ag4
it2JQaQcRnP5NgB2R6x9KD4dXSTXaABIfBGewTLhGPqvkhJ5nbP8VVyTN0nozsW/
MbH/OGFULdJsQRBJJAPTLxd/eX27U8T3McRql/8z6wLKVInqekjehnv6ctkURt03
Lq6gZ0e0YjX1Zr2WsJuocU0LeM0UnGBbpRev8foLzwiDAzCQGob4y83iTkEuyRKS
HHmOCfFnJvpK/zbGVyw/DcroezDlCg3PcT9VBWv9XDTHRM5SE3KuD4U0c02YPMyW
P8pOoF3YJ5+ZoOIy1xgVqFunGs72Co2J1c1mZRmPYxKqXhknFMIhhc/Jcz0wcFRL
F7LzEkWZOCtQv7Rlj/5yc3Y6MTPAOJi5tCSwzlaaxvTy4997fLOZC/bBJBFaYffL
5TEvuXFtJpp+G5/Gn0SWKOzxV/DnPw7fDcY7pz5fwr+1pl5eA45O9ZkUUmRE4c8M
5h2WQrKpD4c8N73a++VmW9sBkBPzH77nLABRIPjVe3vfVWZqEOwyLDk7j1Zii9ed
awMaG1A5Q0urnEIAEYEV7aEU4NtBTK1R31NZO9cz2zTQRKTGupR//EFO0fBGshy2
AxjjK9/Ae1i3vjf42d4bnPu5q9/0scabros8mW/lYdlD40jxh1e0tOLJE4B72lo0
93vcjXgBmkYguBorh+UQr1Gt3K1QWphLm/4cRsuK8w/W9sp4GOVTz3fZOnCGrjm3
XTKxu9iExwffjxKn7zvUs5NgXeNMsT9tC/077uiT8FdJGlVAxpgyrRmsnJULz7Hq
2yCG7+QrK6XK+m02mFREgpGzbbEK21TXbxthHcKPA5VNjM3AffOtRGtqUyrk9f+N
gxOg4frDNfFyT8ewSaEV5ls8OHSnt2Vr9WmEYIWW1Jgv9aPkBcAnGInhXhVAti1Z
+3Tktb9zTv7AJh+0dIhqTQw5IzwdCoxMtrlviJDKdsCqhNufjOdn6Hm45H0md7w9
6HA7VZBhl68zwueb/rETrD+vGgNZgPJiTV6qkizFcz2kYqpo9yWPWuGO5WzOERlK
mS5KN/eq59lE9K9ke4ucgn+beF0r5t1YxFIrfrn/CeWZEbnSb9TjTGDRQtMJQeYJ
ygxeKhpp2HGcQNTNbsqyWVZqJM20MPYATOPx0HonGroht6F9xUlmzDUZ5OclPqDi
eGal8gACwg+o8GAdPH/FgVLm+MzWVX9gnjxwkJ65uORYWS6yEf7TQu2f363UhQvO
wn3/PsYA7SaTFfLGgSLewI0eNLXIsbOQ1Ul2sHvFAqgdjqah2KgOCLT4TUf2I12e
/gO+ol+oR3sYbqy7zOjLX9wePYulJkrcQINbKKTa92IdR7ULb+4FOG2ysa+aqcVW
tAdMs2CBgYi0W4gJVTv5ulDR6u3UA80KE9FQQlkd+q+i0FIoPpVCh0IgwutrP3Os
lm1Ef5bboZpLU5r6eeJfYRgq1m7rT6QmNVagpZrU3dB3vkbOCXPuKYcU7QzKNn6I
dzF1DmBxQcb9Q1zOMsU/HKQPGjOm9FIlDGXqvaBYXFgpfBDfiXNeQVXih0kDjThq
i0jb1OpsaLSBLMN/wKTXzDwaH3Gaoigby7RCi2UAvWuvB7Rp0gGc/W+NRybGBJu+
UvAwfz5/ZVfBiOPHMW377IghUyl+GqN9xqDd6paBH7W+Gi6t8F1g5WNmor1q4Ezf
RfrKn6AUl8a7ylYis1y+EJasXIlQAgLXaZUI2jf98q5daMctYGmCp8evqF8PreLq
9mvEmN/7fpstUlAD0/G5osvT5aamIgcHAo0MuuAGo9oEnBC8KLCyuGPG8Hxyclr3
Mld6XBAaAiu+Bb1Ic+jxOQsECHYE0Iddpv+6QQABupyv9dmFft+GWshzBhrxil6y
1kSm2+hU5M7QjboCk3AntRh038IG+Lje1dt0JM3RXe7w8fw+6pdiZw2I+ieh0zuj
5AZrgOXSXyQREo9Kjp7jtMLDRzEhtbpjN3yhqfEMOPHtQs1FR2eXuZXB3neArmTr
X+my3HuHEnX+L5Vhzk2f30TV3H1D4pOO4YNjrcOMlRgK1u8aNH1itHo1CDqy9mOD
T/cv92rx7PAvPyjJ54/3zJFudFsnNsIsnbK/PDxD1KKgcRbQEgdux8HflGXT/zbK
OJD7KQqAR2XTSqJiKp3O71ypMZDABsst89baSzfvljaOpiYGzfgvFi2zHEoJgCjb
yoRVVfHj7FlBAYuM9HMSS/458bF+SEQ3HZgtw3CNLQwQxj0Dejp94ZtBD8MF7CL7
NGo9ZNlWBDbaKd9ueGmTT4EyarDOOjvA3S6ELOAYwz4hIX5hpbCoYIoouVo7fDqG
zPsnTSn7wnBNde72V2vDGg/WqDAfD1WBXI7iNV+16t+CHUSEnvk4AHFkWLaBGuHS
f52IZlBQ7zkFzS8GM9eKKArgB1Qs0oPcf+7QyAI0K3WM+IS9Wet4a4Rgx5CgCHH8
P73TgfQ+KiFVOaNTHK5lyG54HyELOaFpAjFDxawUH/gerGUFmIjSgI70ze6YfiBe
Z8QPByPVzcItS+ON2SZtYC0WYLrl2F401tnef5s0fMpANDztIvzbc03dlIyMeXI+
0JY2yQCNYdflM0fun7+tbmb2rCheNE7xrO2hrA0BtyzSQNQXW15GDOopm1ojuAVm
ru/PNi2vyP2sB+D16q2bgaSpbTuWjDBdyjzOGdylIrbxEg8/oSydJxPzHZiCHY5n
4OEL6VWyc2FqzWn829SB7/FdOAlv9yJ1xd8XwsnWMcckrL3LC5hJLKdwCProwygm
HtX+Gzg4WsJlhoWRIpnnPs5zz+qmnbLp5WCGD91T45RtShZKdTs75OSaaaTCKnZk
FP24XIh7bzjJkK21EyUCGjBORp9kS5iOnxvghGil1hbGkyY8C+xjRu0Fg95MaHJM
2UZwR+wUlldh6k1lPLEO7QbPoA232A0HJyPbribW6WdF6cz2UmMx7fVs++o+G7YL
9dtd7h/rQJlc85YSOwPUZxLmwwFWFsGr2ll8mNQgF1Apslf2A6dMauj5U8xQLM2e
5p2JNvEU7/vKIrFdebHYl9ZjA4rbUHVGLevZmTMePm51AJ+gLkXyv72JT7bTI3Ph
D6m54hgLd3X7JINWWLvlcwCduk6HwDMTy0r0vFx3ENAJ33vf2MybKdZiiQA+/+0l
qXNvAljbbgaEf0VtFvmVfDCOIvkb+aNoJ//VEe7zUSIITkyXXcbn9mByirP5pp1O
7I0v50SPONCPwXpF0ogXU6c5Adp9BkI5PtYauO/nnZOurq9hUsO1aABUqkLVmbTK
ntRYIdmsA8Rtbo7WDEe0fomOD0hQ8z0vCqBU5MiOwSBmYg6ZE9X7tO1RxhxITTIR
WVDAbYUKrSPkOg60tM2qZD43mT2lisn+rSSZRTQ+RzhuAFUYqq1h8BKmHLyfFEXt
bN6h9Gu/MGmVhJI92ulANUD9tnM4H/KXdmxs3OZddgfWGGJuDIPaSmjhUGSjjyLC
8d+6bDOKWcXwRi8Wo1uz3Pq9T/mW8oypuyUaLbKz+h8alV5XbPOGXUZ3o1svK4VY
7kz7ahHVDMIR07o2DTkwwkQJhMPD3GLKAnsC6sZUb3M/5lzE9BEqad/De804/U2M
QtPfHXEbWE1b9NPsZW+rYH2VGPGyMAgMYOvDFwCjLR/b/q9mbiIc0J/Fs/aPEAM6
NTC0/YzR19vThOCZGp18T6eiLLfHKr5NbshrKlmfrZt4L3eNTsXElHeH1ITL7ZYk
CJD6H8So7cVRcm86R6+eGi2sGJdd30Qq5AGmawJJ9mI+0/XGVjoUV+VF8apUeQN1
NpjIClBhCTotf5XUl9WypjCSuz1Z6h4oloB629loOvPl9z2zj3Lb9aUBErNqRzmp
eqszaphoAL1An/IrK2K/NnVrMrC1iMFxLMRU5wviopcRi1T0fExpJNoVI/wwYvGr
ycV1IyCz3aiu3n5JANv1WHr6CuEQHivAlYNCcfItSyhf2Y70j7AVf4VFHi0DMLjw
/8ItNiSkyDzz9b0VjZ91CIBf0lcUCdB3rCwb1FVNYND+jV1/wcb4qOnWbt4bAkgt
/1/1iIt/gQgVGOJiy06EHKuWhRAEwpR0S3saXNBifDL6bjtb+dQM44izEzgE/5s7
N9jL0MEmNsIAwnhhg8OAtSxyzMWPqu5Er3viM+lBlyGeUbGAC9ZNllJOFxphz1Qp
ZAJ1MtQ58ET3EhlxraQtQLYNUXr2EXjQmDArRYSGaQmYHIHrPAdhrVQk5JaHedJq
EKy4YpJXio1Jaojt1koG54ViJPzoQlLe/cjKy2zBvuUyPvrM7uI8as+FwHF+L9ri
xE2FKJpeTQME2WhceWNKql6XnFzCYm/06r1BTcnruO9e+y1z3n9RKZbNCJP1/1LL
7tBKSCBzZ7rfMw1W/xNeGO79nwkNaSJWw+sCOjFePGIjIcVnilxzQrikE1ZmWzbf
eQPXd+/UU3Fwd20nATtXAPWVRHn0x5UEM5t9g+G/Vuk/KToidisk+7ExiM5wvT0a
t5WArm+SIdD3aWNaWZ20CfhzY1rmtsz5PyvuD/lRvFdVeosCgLOQSFwJT+QzVopc
BjxaxKiyNghii4fVYIODyVr7r//0Rj+AKyimmEpDSlMYSlEr0ClxknOTwTCsTsUs
xhXl2hGG7dGMpAJhz2XjN9xWIRBUm2ju1Hy+KOscUGLE2rfB8sOXMmQSxC2efZxF
Yj3eJB31tNbC7eK7rBm4Uq/uuNYts16RBIkpXENXLektY0pLPxWcwTOAngTOCsuO
1nL77TqFw5uLMy5qs8yFaWxxLsy13/9CNzKml6sIFZNZTZd3IVG0JWVl0LXx3PDA
Upt13QJpBTTN1k0VJAVvywiBomum+plrFY/BgWAR6Kw2vzC0ApV2s5lbQshkBQAY
zGya+EQ48NSb2OXpKCS6RLvj3UDQYG9XQrPlgQs8ymdbZJd34okDi/g8l9BTol7P
uER019U2Ajf375JiI8qCGRuZhvb1KjjInw3YDTMpjL6n++8ZLw0YzjJMSUX609yQ
TRk5c6JY3HLsVnjq0QhCkbxH31Jwnmwffu+BOZLSvHKwRv8qMGfYNhRY5aPEQW5c
J+M0zR1AJJ01DViJdwaKOhQQqGdt/yWGGJFy2mOgSASZSL/hUhq1pn3tLrufadwz
6134jPHazT2yATzrPWj680Q7DnqsRhDIaMBwPg/tlDYwNzzOxmLkkP7MpEyM5xX6
HrlC1rUOCbnDSHV9tI3IFj52TtlymGSnpQh1eZHYO+5x812fwmLE87yuNoVws8nP
zvJGcppgM2+GGAWOQP101ysUuXbkSApVqLju5rau0pGRH7UiLzBUEs2gAb4IrSws
PIyPtmRi1M8TAxcc2bdgQKflo9zlnpkx3U1r/W51w1AnW6hC3LvbXeqZbNDV1zx9
8pJjyd1e4lNsfaq7YSjictSYnv2DANbW/SuEcZdmeQDo054kNmBwfedydrHoTMyH
jd2OnKGIhyk2b56kwbxDlykIHzyFRX9E7nAONVrfmgQQIo6abm+5pijTJjDvVP9b
E6EJKl6upRBxvlsEoAQJkvEtZcyI98spo1a3bSp5Zg5NiIXVTrtMomqRPXWxvDow
s/uMdOYUN0Q0pW99AVHr/pwECOSeBv3/CJk/tzrW/1WRMzNYu0Kth0slJb7cIu9I
62Uf56nIc0rlBy9XTNJ82LuM1JxGUoee6+U/CTZpp80=
//pragma protect end_data_block
//pragma protect digest_block
ftXnVGHOYLMbFTbsBCrHvj9Plxw=
//pragma protect end_digest_block
//pragma protect end_protected
  
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ZEfxZ5Lz1I6RVnZFPg8QhhdoQaYkzaA/NxMLWLF6M+3hLViZ9V9IypfqJkryQ+TH
agXq9QpwdYj7MvXDldSr+KJBh7fpi6yraOFrryGJGo68nS6sANY12YaVp04+sLh9
j9B6O5BwPmECHZlZUYLEzTa6VYsL1LWGF83OCZnGwheCg2aY3GO4+A==
//pragma protect end_key_block
//pragma protect digest_block
CZ724colXf27XxjysdaBYbh/eZo=
//pragma protect end_digest_block
//pragma protect data_block
9yWK/U6ByLNK5qGOD5T7D928LP+C/Qzeh02q7baHAFG1aCVuTRXoGeK4K5lAWc8E
+MJh/UuBgopO/xNPI4hC/C5zVOsdMdnBaNPCg1cIPt3xwJpH/uhWZV2HuBSKVYSA
AH5VXcIhBiBy2qJGkLa7pvAvn3Z/IJvkCBJPujTHkHS6Sv9ohJ9mnjWe9riWrBQv
uB5gBF1DuR1/r2CHPFGCPMrcGGvOLYxt7P6UOMfa1juO77kWgvD+90Nscx8N7fuU
QZD33PcvMY14DIFTNNAnPvX97C6oi4lT3seY79fcaarK2yoBfnKNJD5tWJ6kzybV
buDYL8s3ZBfKnq+wPqhObXM+vydzJuzGM+NWi1KMEldjPpX74GXe3vBfDhSBROhA
OTTl2fq7iCxIelUA0lU7flAQSXit2lMisT4hhpLKXOvif4A6pSdKKoNg+3Pkvf/c
5efgwTnnpyiDTRXVVntexYHBvxA2jMe2jxfVxpKGyXJVoXc9bfIkoXgEuU0L58GQ
0VOsFrxylcE8asxAYn6iugV5KujtMbU9X7wATzmxD3CoO3uPNdWMhgeXc/iGOazy
UHKDzc3yhbDzQZYF2M62flHiYn+QzL20opshkwWq2vqRryvBtQ8TAaQApASLp9uf
tgWK5/cAPLj7p00H4IS4bL5lPatbse0X8hLWe3mAXyYQ2Lg2HdNG2/JGXp88vMOA
XvpyuzB/QMqO+Ao+a8SxN9pmICP1RXLolojYFEKI6m5OoPw6AYmHiNvZPNYBvVcJ
UC4D5ewqmqjD/AFvGZfzKmGvRuBxSbM6PSQjzTcg8yKoMdU1h9TdYuq1Pz/iOODY
eFaujUN9FcWdXeUZWRCpYOa0Xlcc+vXtnadczXc5FnTI5C17TFRWm7YcqPPp2HqB
AhiSZHZSRbsrMGBi/7WsGX4EkqiKg/DoKWGM7MBGeg08UVphZRveYUQpWgouR2B3
scmlXoNNEC1BQG3BTEOe8Xv+e2mvBETC7YZMJKnIFUXcweckM+uxGZcWz5K0Yqv3
lfVgsRlQBrUdu8Nl8pBLyMwUGniT0n+KLveD4yySbzDRPdiDfVPFa8wAzzQgm8mY
lD74DJXRTJtQ5gY91lfOmfvsFN/HtpIXZDOZNLtI660zbTvTC5MUu92rZtCF8I/v
n2vZU8eg3W6yYR4zBHF7fH2aqSSJ1L0XXW4dygUmXRGPjb18fT9FC56+1bM9lKTC
Qjnx/WzgF0ADVuwFmpB9YFhjK7E4en6+0dYSNUlENu+B3Llqt19hnucztbRAgpJw
1xoN6wbfam7EOOpMGAJx+WDN1gslA/SD1tKTPM/GmyFmTpTg/h+vtFiGgaALRAXx
xPOS4GSF54zlRJMBeE8f+S5cJKPWC1SAwromby/hm5/CzvDutb/IV2Iih8EtdU9h
sfrnB7vQ8d1idAGpxZUiaqqTFiJwJbclprlAKqwEl6dpZMZFabi26MBMtldd3ae/
HKJYIL9q1EVfmm2J9pI5j/MIEM3e3942Y44JD/bi0PrH/ysfxwO4Ak6sfwZS1gB6
TbPljjiyw2Q/CLmijfZAQI1JSPUJrqTn+p9wlQnH+x+hdrzZg9YyoQgy21kyoNwM
ZQWqPW5C2K9PuBctLKDCLMldh2CUbmkzsMeD3iWmpopYkpI7qQ8W/QsILQ34zmQg
15AJA7XGXfcqWkRX3YJOjZvaTQ4v7W0zYCJDzlBPMlEUvomJ6w0ywNHHV16iFv3k
AkKBCVgR1Z597Zehx05QM0F5YjdNm7W/IkH/tHDy6K5COVavRrhW1rOu2YZjjD7G
CH6ZC6opdFiCnJQePwMp/axVqXJnhf/Tng+Dlk4SYRvSEmNh1JI1gTUPjooTIGr0
fpOqfSyfAkLWR5DeP+OyPGDp2GpW29uB7OcsaTS0C4ZS0SqFBMWGfI59zter91PG
mcgpWp4Dfs5Nhl8/yJVmWIKT8U0juX5AR9oHkWuI0Kvg0wJXKsIsLe45dEoeVS52
G/BBot7US8//5R8F0B2W/uMqhDUdicCBi0fQKFj60pZsc5AMInbgyxDE0yvz+o8I
13jhDar7eYvNPMYxRtqMCojWGKPZTgwVhP9m//6b9XsffDVTQSbqzSnUlKP2lynI
okC1c8fFXwtMA233WRKargG9sG93l1JfF7JU6PNFGU/HMCz4fTGOw3WPMW3wkANj
eQbE2QN//VzgkOTm+fCDolTBmdusnnkqzvGhRPE+MoHioWKM/NYK10vaDGy5Kaw+
FHYKQQWnA600fhR1tXv2cg0OuCr03QWLYBf9RnW3qJmA3iKl41KN/KRP0rlHTx8/
qrM/CZek+d6YqanlDgZ0NP8QjF9WOHCpZv04fKPoOaKiy9MNqNfxODAP6xcXhYCZ
Wywo+ibD+j8/2YF0ZqBPVySDsHa1s22zyeyYctkoDmk=
//pragma protect end_data_block
//pragma protect digest_block
7WokiHWoj+TkhbOYoB+yxDiqdT4=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
G1nRPBUzxk8BRddHyXasBs29dVGJ47xxeZr29PnVWJE+FyQweTlWL7Ub1UBSplDC
YTze+MVu3IBsmaf38HtQ2yxZJXdD4PDvU72GB/IBXhVfmRvwSe6eoa8rF8/aLtzh
iaMbVBF2C4OAXTe2CR2zz5q0cVD/vdRqsofSGqlSeasZGjW8NOhf9g==
//pragma protect end_key_block
//pragma protect digest_block
fCf1cNBs6ywBMd2yNmqVIsdnX3Q=
//pragma protect end_digest_block
//pragma protect data_block
/uERWc0eV0/m7gt/n9E3Ur2in9kWrhixmDxC+76OyA/cMYhuS4APGF/cKMa250FH
Vg+6c5qTXBVQUnaGCcHTQGxLrsB+RhFf8fqGWRFQrs63YdSG2JM0NRxpvNJxENoA
7SGD+3NfSEkflCDL8oQPNIugs4hLXWoC0EyUqJCjTZma6ORKiAnGJCTDDIoXiPy7
NgbjUBQJOxeK3DgWNoRCJOgBd8Oy8x4L6G1mBTiKiy+RkMZWd4VIcfUDa913p4qk
it7z8ap40tvQ1Vu5vVxir972+UtkjetdePLUECdMSKk5rf6hsYhV3IGEpC91QVtg
uc9hBfKOqjDvrE0GVoverND36K0tGht0LKEBb0TRdZuin+A1YhfThAbPnFQklNBy
QjuolMeWoS70tROnvzjmXKODnDmy+IuyvimHtvOXs7y9p/qSZEsR8Qmnt7qrei5z
ZZfDMRyU6N0XxBWwqbM6SwiS7dsQ0TaYH3HwFtO0rW2Yq2dh0ZHf6nDttnCbcC/e
vG7KHxk6El7hBwv/Yy5EvCCW62I5gWhA259pi+s9Ybl7c+hD4JfGsBTR9Zd22DWc
tzmAqDDZhymN6IbH1iExI0IhYbbTu5jS0AZAmjvicGhmZHFigqyelmwyoNP+P4ae
7cdXtpp04TUvJvJsp6Y3reanHa+9I9KpcucfBEA5exGTBo9qh9ueDUGD3VrYmmyb
OhZiawPOG6uuXi7X0eliAF0vUaJLyCx/r9J/xcKB9SsE4adFcBJL9o+CVX76CIUQ
lnMy91c1mYN7aAPk7QoQSoaRU3aCYX0Tlr0DFeZ2ZADlUCNBO/P1EsUIGCU2ksph
A/oZwAWh3MbgtDwKbU9m5M+BJKRrFXJnY5Vfxlz4tXqxYU02+ZnWvbkXuXwsrMuE
PxjWJJFWu8rDEFYXZcNlkUF4lGs60vcehrtups7mmPOTTIIgr+if7ZGWVQ8f489q
c6h2VAfnGuDyUb0W73U8yEc0zy2HEe+HifPThnpXfBkOy6PPUcX5Ki4GuG57n2hH
oh1Sx2DTA9lrcl3Tm767UM88rOoXoZmaIoz7ga6n2NfEKjfxBp8Dr9UwUX69g2Yl
zaT8+LwWnluYOEgJKBMozmIukUWKxLk8kiBXWrzReKzzHV9En1RzDEKe+qTzmQCk
hM3i/b+9VtoeJd47dAR8TI93xrzYgrbq/sCvH9h1ACL6Dl5OXzieBQgzhiBxDSXq
Ex+3rndaTistI2tvXJq2bmT+UPiR3SjAOJXAyEruHykHZSuZq0Qo5+tY/5tkx53H
dDL9XxsRi+M2bcpF1rLgHnD+2yepBVY1vJnMzBsAahafRMfUpcuAfNQZh4a9zHCk
LF5HYso2ufZBGdtPQzncDRsnAXJBZPbkknsrGlwK3UXeLhN65qfFmoL/H1fs4EEP
bepFJsnQxt0PekCB05TGlize1CuWM1B5LxMlDnexNIGbnXucMTLjXkITX/xLl3a1
feSGBn9p+p85fyMiA0h3NSHsDsNOni/sCnJ8MC/t080fqAPaFG2HiO3NvHxHQNQ0
zk4Kp0dLdX3j2WwrRLZ8MPpHS2E9Men9ZLwM6U2c+mCWVFnhnDz7tlaX66P4K8bT
lyzE6h6BO/Gqgu8TbIaZ7pGX5LQSGlgtdRF8qu+eeu6RtsM6LsoOM87j09rCbHx8
OaE5oLRKx8/Kpe4n7EfXYGA8jV/TmHJoE2bpe5P7zrDwir3BVqoZ+oPjQR7V3Szo
uU+BtZpoSPWKmfhkKSvxZy7BWLPhd53pRN2ejVaMT0E6FPsTbh1h/rn5Wt3zhhU4
MkS02HvsFdv2eVyvmNjyt5FAytT8dKBko4/JJkoj1VYvAv8loe/jBU8GmXJr2b5L
XVCH6eIwHGxYH10jKn40axoaWvCPyPzut2ymh8j9vNNL4qaj5J8HVcgnpwqfuGq8
DRFpssmps3JyEWhXUowZIHL6gF4tB0jgiUb9vroisDs2xXdA0UnjnnLw89udJdn+
w9FSTpBWWI0/QmHdtNywirHE0g/dzJy+MoXXFqn6z15/omOEkp8ADdBOU/imBy6u
lQvclix1KrgzvwYesRn2xNPjvFz5COKZ/2VttMUOjlqjKq3/wU2JMoaqQhv+swUX
fL4xKaNc2+yuf126fe+AMXmEHmdLAyFquLCsF3I0g5Pat8VNuEKTLYLnE/jH5hf6
h+VMOIK/qBwVy8EAEgXQGBF4Dn5sHe0mqeyhN6LWvayUfliTPdcxkdfROYkR4yP5
VyEkLSNB5XH9RlJapeeSERd5sLT0XY4TVsYfeIHX9o8gQIH5RFGCvK8WebJWOz5q
ctW3aXtal457k185tLul/Tv0mkqf5QUBsspU87g2Bfi1nuqyaZxz+Nadw/QJqqBg
kTupwwO/w+x7KadvMq/FILEX9vpyj8l9drLFJBXX/fBHjpreRKmPJAzJT3iUtwmQ
y8DY+Cd76V4VsEJ7Dtgtuf/BDV/lxeqfZLC1dXoUJpjbHcWMLVjwy61ljccRy+4G
NbFVRL+QcAA0PLwTWTf2lMeEPoxHUQBrIHgd+TcRq+gmjXXEc6SS8VRHURROv9tM
MKLS/loABVPL4OY+Qbhsa3K3OqJCUGYgWEHboQnZO/n3eQcTOzlZQi46NmbV6IUs
s62WgatFnRJ4fnAiCkMvQ3Eh0QFYC4opKFLTqsjxcPKca+4RcNhTPPy5iKc93WL5
5uzF8Vo2DIxoPVfDpD2/qLABK6ldRp6E5NqGmBvON4wIAt2RFQBteengyAACS1lA
2GgRRZR0M5Sk4f841GajUtesKRqPehjJLHUnaVTlPplwBqoS7jqSf3oc0vu1Ah7j
eJbs2b1jbU/iWt5soQRCIuhK+2b1NnSPbm/szmcq42BY+ZQ8kAHlZL6owbKdJMOw
RmVEHykIVborifK9n3rOW6O2Jmxjg2WQbdl5UbQZmxUmvPiMo4ZxcAltd17Hn5e3
ckOPYG3wo1KhRQcJb8wQfgdGp4L2FxWCH0XcANf/dmvYuApFXrGz6ie+ICUDF6WN
c2LWUBK8CY5/a49fxSy2vJRRKS8WQDGkHq0rlfilO7wVQMot+gaKftWAT3Xj/9Nj
vrIka5s9JbLOtgFYdFiP4i37uPEN+ppqGsHom5qQbOdye3qAz+1Rg5sh3GitfJ74
gzkSC2Ykk9x1/3G9Kdde77947Thasy2bAKireaJ0FlKNCWwkc/QxMV6JNkZjuUEh
fZaFaUqbsrdxPnhfVolCDhzCaEm3p8x6bUji9LTpWG0xtMslSjsLbpz77AHXJ+zy
cifHn3sNILnud7nlx5vDChzlHPrkfQtF/DvFCfjdsn7VwpxOltq3zWKSJBVHyKBd
kXTcLM/wYtHtmWiIQEkyuwca6+oBr1zOAMeikwZ5LmSD9skh+i80Vt6zfVc/d4Vn
UPQK3CU0220mHJ4D+2L/1+VzllxG5Qz0/FDIlMcueUXv38fg/XKDmSedqNA4BvJ4
wA/F0hVqqqtKgR7YDeU+vLtSid+utvj6ZucrHgzdkiO6JUo6FUPzlVQhRTe1I6Fp
V1rD+rxHsgTzxKaSp6wxDPzxLjpjsTu50tDTFKte3dq3RUMz0Rs01u9OcJ4ryWhc
0poMO1cJftDRZvZ9A+the42NfOVh351loehAoH6Mc/pqRStr8IsjefRAlUpKyJRL
w2J+NwBGGxMaBYDIgIlTpft53qC4V1fdPi0eDLusYo/uRHGFd8XhRLhMWh1rkaJv
bp51UUbxUPBlrvkOEBh1KhjKiTBBgFLImSsssKC2/jDOOpUHczpSfcyveN1HtNX0
KPj6qY0deStOI4hJLiGsmy/Z/xPKQSozHdjivdHZ1KfeHLfSss0NvC4oZTj5jaII
pZwbqd3oUsqIczJ4r7Bt9ILzypzQbpTJrct5RrN+MVTlXjTujMKhT0byJG+NqdBF
pDrMQCiBEOU0exgCnzLZufYEynalt1oZuMN7LU8Rc6uQ9Ivw/mPHLcwJkai/ZdQW
cdda5T5TKjGqWs2YzpmwyXANd66jaRulKikVyuErRW1nTc0Px+qvwUfEtY1smWAk
qHmXW9Jb8xt8USXAd/Vjk5qkE1eqGP8KEz+ibbMImIRBSf+TbBKRn6lEonm3yS3Q
MX6LFZDClJPdq484DkoF/qeSjtuMIXZxtdonFXT+lKK92FYoGmtwE/APGw1tU78i
pEYsecyz+P565QjCJcSGor0rj4BIovx1/ErYmeiTy+yzPaX5tqQjMarIfzJuXlqq
0w6in7i8BTOBnrFW/rZdJgSBImm1FAJuLhbGJCS9niCdmiua/AucKBn7RuGA2X2g
71sV2q/jnR2QE4FLvEhwbgPZ0SBNdLjHCTWWJwUaovi3TRAsfiG2xVD/0yt5TFfp
Wz6NDsDqGLztj7belPJOnI3mAOhpnJBpvdovf9a+Huv3+lx5nQ/mUFbN1oxE1IyX
jhAmRF1AqDcVnW1Sqe8wePPgbLRNU8c2NGfyaTDVcQPgFjeVxS+nVGb6pfB+dcSn
zNipV+7eTzqWhFBsOfUWdnnHewJKXiEXvHMHArRf2K1DVfvZMSl3syPotNncIYLT
eWnVv+Fkui6Z3EKGQ5u4azyc2sVHtyhN5/85KIC/B6Y=
//pragma protect end_data_block
//pragma protect digest_block
CbFlCgb1sMOc/r1eCfPCFOJsQbI=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
xRPzr5VF7R+T2r0qHyOCn20YYecgRPoYFnZPKWt9u3/lKIf5fSraWF/5srIoa6oi
r0F3f4I2Gid09ED8z+4HJq/m+XcxN3cmTwaLrCMAPfX6ektjiWuds6cGkR4d0XK6
kQcJ/CBRoS5zBxB0TQx1NDyJJCl0tlwKf1ErfriJmX+6/i3dgq0pHg==
//pragma protect end_key_block
//pragma protect digest_block
UoON7oGJfV+H+bPi3yT0An1Gtdc=
//pragma protect end_digest_block
//pragma protect data_block
GEcL/LF3PTcq/12VciCxb+hECCPf2kT6EFUnAhLVCmaEF+Ns6RHGEaKyPRSUQeE7
cd3KiKtF6Dj03TPSRFlt2U5egvlbCGTIhylX7MH2iwLClMZa0HrIHnj3pldU6gdu
A3Jnu/h15LMoBMzxZL16V4lwWxqUm3qdxYxADpomHnCKN08NuM5mOm9AyZU2lxk3
ztbXLag+XOAk3u5cmwHnJKiIOcVd1zOyUasAVKTnn0jYm/cpUWtlPDRXJaVyZy1j
rEL/rAK0fQj9sx9iFPSI5yUqfdVUfSvwZlebweQY1B0F1cGuoWsV7VsAUwfHR8gk
NXx4qeu1s7r9Xxypnz5+08/k/suKKZ9VJQlfg0TB9IHiHKdjYePnwYScB6AFzZ+y
XwJyqlUv8HT29RLdRvGiGIUU5zcqzGIFT9gJ/RHpwDWmmHepySitJDASxgA+5BXq

//pragma protect end_data_block
//pragma protect digest_block
8GSFNhkZ1nm8Yf0nD3P2Mq0wOhE=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3m48Dl1gAscwg523lmeYRd4i0sTXZPqfgMCCXKDeANXGuRQr4vdaqWKkhr9h7M45
F286X6Bg83ZnicZ1lMQxnHiYEYw6/snJnVFaLVHEvYbPkr9VytC1ew3Qld/YC/Yf
8uNBH/sGWUZToo6zBwJY7BYPKJKUlxs3HChJqKFX4dqYcRlycysddw==
//pragma protect end_key_block
//pragma protect digest_block
cW6x35ff2udJe8LUWCILzAWxh7I=
//pragma protect end_digest_block
//pragma protect data_block
okZkzh93djTrVzbYfSrAemR719+iqOzwdtiqy9hxh43n0KWY6HUbcV9RsquX2rn/
dTHoSrWpqAZpQoCzNoUR7x4+HKWh5/GhJz3KegIzieUtC4YbtIiii7qnW4cmEt1x
Zhddry4hDgJJqfGeoBuLC/8oJOeNocVuD5lNrk2mTbKuJh8uGe3UASPNm/JB5r2K
G5jEWrhkr9eb0THNGfcxxsn2oRWLCN78kveS0ofVn2FwrJQrG7eTcxY/pAeIETFO
Wggb7WITqwa6RK2Kv8cYs73NRQUdsD+bUcCS4hgLgtOZTPNu7f+5msZUpVILsmYe
/vrbNdlEesDjuq4Je7vRVpc1x/mGjj6xzhpKIb5Ns50YYHZj5Brjw8oz0pFCfq9j
jt6V+UPNWaKpuY78kyYVmR5aNAMQn1YpPxT78a9G8MGaY9bSVwbS1Mcqw6OVLt3v
B3MPA0Nnc5xACLxS1J+1NzDV2PgT08mUgal/fDJzB7F4Z8Rgkaskccs4F11kBJNG
XYm6YoCWXJCyXjuqWvIIyx/9689SH3F4ytGj0AgLM+ZF93JSvqN54kVIyZYQ6qBh
HcgG7zyEaH5oJMXEI88aK+gS1/0hZDbUAb65XMlGE/A4zyQliTS9Ffmnyj9EdnKX
w9hGghSIfgbSFV9wpPmOrzSf1WsUyRn5MAX4neXrVYYWGxU9FRlA4P4acqWmNbfW
E7BHdZ0BBDE5+MGFfuOJ1zyH6kxkiveuAO4WPpD+MLtlxtFi3e32XlYLOwiFAGBG
nS8bq4bFuypXFSG7Aksz6HEwuSPdHmhQq6zpL4uNOjndTZ1vb1RRb31IZSh4yezq
88IUYBW24UrPdHSkwm7L7NKiGA6d3XmnzNyKY4uWB0t4WYqt9QwaZ4P6YmWqOSjs
/1RixMcCNMoYzsRVvrUrSZrN5o2uipiD2KURfTKZ2yH4MnItP5r3g6KHpQqaejrV
wp8XFTbYnO89DN02hYfKFKT6hdGrBIs+BxybZFQfEilI8soz57DZR0LZ+wLda3jA
RE56p6hI3bOD/1twwpYiQhAwiYJd3L0kZr3azsDQQ6TWmYTOcGRbk9h+VdPhDuyE
cpRgWhlnSUwKyyKFYF1nk2uesoQabAYQc79c5eTPqv6RJ2lP1gcRqYAeGMVXFn0V
hTCtG3cNQxgebg0/gc/4TUYav8ip9hXTzK5orvlb26Kf6i3pS1syfpMeHiHc9Iw1
OW/Dsv03Qe2Elp8pVTVXiNa0/FJzXqo80kIkWAW2oJTc4liOCQvJxz0Aq/OPqgQ+
PhKwkNmpljTR97eLa7EwJh+0p3h/z+oyGfYojQU+psmouq1sg41Uo3Xu6VkJqmpY
tsAukzoNK1PV5exwSqL6miHdrxCtvGu79E74Ilcsx6BCvCVMA3Msv5OK33sqkWmM
yXQAEvLqbPOrqR4Yxoxd+IRPyV+a0PoJB+iHunnZbMwLWGpw9pyPbHSAKdKp+nbC
V+bPaRmBJL0Ri6umpqVx70j78MMgTyte9Fy+XQp6wpikutZ9+OM0n7GAE668NKBA
jaY7LcFD3WmjVCd6BFzc+DL+SQux01AAnk1bDSr4/8aEtLBqdokXhn6iJ+Y4705L
w+kp9eOwEZTm4nF6ygwC1XbkAHBdpuX6WQ8lyGAgtGYrStPRWhv2fw8ePj92SKxJ
PLYnh9BjwH21AYe01hNPp83Tl48RiUZxxxlrJ2zY2Vvgu9yzbtv/po4OhSBA0MWE
Sidm/9UV+pWk9pg2rzooog8/+cmYYvSn5LyC96oGm9oa3kIMjVRVW0sUIlqf5ZZA
7xloSXcmZrEL7ITtSbajsuYUTJG1q7ShvEonjh+0VmHBsbeOeI00VWQvdv48kdxo
h1WUEjlOtcfZPvo8J2f/hLQMUZLQC7H9vS4okhKJHcqZVoZ9wT6thnPYL2XbwQVD
fPBDAv5aPrwW8daF8S0ki8l1pKAtuMu20D4Hw5VcdFfRP3XVhF41BXDPdeKiTlay
uZZwIITwZKXNW4v1KuFZUY9VtbShutJOzKw6bi08lOhVC//tOsKOcCTk3+zAn37V
aV+jhjiFOdFFQ+kmvmFY8r6ir0DiBASCLhDdpe1jSUJzzpmuyIN2WTjN7IgM+0X+
FJuSGrEER2Z1gktIFccFMCWewRXTLr/sX7EjNzhApfeL+3DuAUBn2zKtWizfnVjX
6bAPUc5zuupeS+cZ5ZapsFcDAvTIV6qzLupJukPPRU6Jg/ixFm3pQ/1mjwMIXW+Q
PBIaCSOOmRnWLO6i7oOYwXtMBeHUrx29/ge28dyGdp/7fsNcm3x/Ob/dk02FHbk/
jzYtlJJ28oyBdy4bcnTUj6Gvm278LFkvVVbDvhOu4a+UfU5QCR+8aCVH2DeTOBUu
RW2ajF2+sRBigEsX/iuv4z1zipgj4x8N7gzOsejtMXBoLkY101StwGvjDQlW8Gvx
3dAz2lxlbqL/R5Mnjn5VxsKC/Xmgc7jXaNk+eSUSqpMQ5x0yFb6NCtl+3sf5qrx/
Iz2m1xW7fU9fsEW6cCou8H88jz/fmgsSop3fJj1cyueYSz0sQJFTT4n0rJq6YwL0
g5Vw0b1vNRqThTX13RM+O/7+fBV01fdQdkWqLBc9TGzkOLuuBBtHgGmZGKMccXPw
jdR+yZqJsfERKmP5zO8zpa27tr0/F/p4ApaOexMb/xYa0a3blMFo8UEmll0ZFObi
0W9ti/MRKPUu2VgVUvW6f+6SuXFrMoOrOPSB0qamWcGS00KmDAIs43JQUYCvpMUc
JcTujpEwUiaEziTCGb0gNI9X14jbWy57Nc0UOVp45B1+zpNVxakzg8KfAClz20ba
FgMnaWq5aJ+pgWO6/YcU8rJHohkSVS+qwLnnmScQFwoJ/R8o9BJYLUZHmwJqQv7e
D1pHTg5XUgaZi8fX/OBScrCiZrhaIMKnxk9GRoJvgmadT1oGcR8kCW9z6DFIPSHt
JVrUmuCwjZ7dle4MTEexaswr91Bz72KLLk/xTFcTDLUbVgl28WBKDGna9Wiv6GRl
eK4yuobHElIqWmlkNEJNGR/LhJ5P8F4iz4paYWG2irGi5sft4sepNChT+Bwppjyd
PfBiUjG3o+gLYkCFeghUU0IuUYaBQLa6gabKionxmpvvvVbqOx8I0hEQ1UIihC81
4BbC6HkZUWOxrLkkQ+HDRGPb004AAtYtdAFQajfd3kFi+DZBB6Hv0ATAHFkDc3Vs
BdCw0a2dIWH5yhZiLbobLs5+Efn/J6LY+/5bVua2g0dhACnJpglLzF+j6ULvHs6/
+Jmu4MQnzJ9SiP0siRGl5UlkzjVn+4IVK41fcwnGCBZqVDlpEvYOR54bCMPGNlA8
YI3YnH7x1YwmPJy1MNC4Yu3rq5hC0Do4lznL5pVybvnxGthRqycLSek4NXgzmYBv
4+NOteTb2T0Q0sucVkOm20iPU82sJ+nBuTI07jaT4nMHcvhFwwGZxTCot9/UnMI9
SKWqhw76jZn0z8cRb8Ju6wnFgZatPNEPM7jqlEMRkx4yJfrkO/y9jRauaoKy1xjq
JLuwfFdwo6zrKxdlQV78qm7F2iuFd7U9ryAlsSyJVV9L8cU6ULfSYW0jSjEcpOxK
HNC29RmB9/Orio6gJ9ifkAgsm9T9Zk7vUp2C5sM5+LmT1fr91gqcIh4Gv11oJyOq
MU78pj1oVzpfXIFY+Yz4YxxzBEMsPN0Y3mbCmXywm+5gbmF62rtrT0ah6upxsGdy
zZ4c7LU37Hkw4GAj3yWKgE2i84/c3J8HB5eMV3WK5tDY8toNVd9n606UQqlOOOyO
5QhWY12ybajWHtdlavwhPuO3/eUZbDFy2GMqQBpuUDMuAMrP1z4JFazw4NcONeY0
gwXUyXkShb5x0qq3bRBQz4YF8yR+X7xmQyj6ArT6dVPcLO40qlo07qB0azWBYF6O
w/yyOBOfH8H3+j5MYe818s5au+6Yjtpps2cyPDWxb5EcFNhiN+tbEc42+4rp2Xy2
CvD3qYj+DMZZSuX8tOl3mcjXzf5wN+Yfi7XjIcGRE3sMIP1ZTIucTQGq6jsc8wxr
ZeQK74lDbD7R2Tf7PCaQJSBcwJFmtWoYsbRRMQjoohVO7nMjnO+Y/Kzy7fd6mm9g
fOXvdtVYEbRPO1s3CIK2rb0vbuPYXW/AuGUNdORVn3/Vl6J/TC5r/18T5WcRjm+9
nhcI4zC9uQT/oKR2fuASyUAfY/T1IZlsYR75boQY8iG+XEgiUWOGiMoqDpsXge7o
N29hnaCSqNh3MZf0Ughbd9NXUidmZqG9mNQWvFdGwCz9gCPeccSb48BNsWyzsOk0
B6YwNoX3Bj5LDG53+WvEbQkxHgD47Pgt0tSZZI29aqKF+1pazl6148G3GQjva885
JK2v0vX/AwESBDEiRO7rbqrLC36um5KGvnPU1GkJ0XxVapRABiSz6AZbPkhpxPJJ
V9tdZCNo4mPw6uR4fJd1NqmqIE6YCy0rBgmBmqghq0KETmxKYde9pZJsaqkTbU0r
aY6M0YAznL6cLiSHq2DfZhc9RrSgsz8+Bn82zVTMu1XPua5mHXC9J9TZar27hL58
RBbKPlZ7VlncJiZ28NS0cUyYAPjV+nnP2iTmZtV1zN4Z8lHVWwFZEKToNvS4/FOV
lnsKUqGv7amdwp+AF+qMRxpXs/Gv6aFMKvhsD0EIIoZhU6hpqKbn3lGuZgzrCwSp
OpoRDiuqZZ7dguNuABEeezk32GsRygIcEyunwxkH18zFI175Gh9V+XbkeRI24fTn
vK8X+EKLlp+YLY/n6QfxiO/naqwCZDM47t5YF2E7TKSKfAy4pxmi4Ra18XnEw/Qr
Iowuf3xk7/4CUJPMaX3hiigzKGEJ5WIYxclTbQvMZ5aTZbA41T+4r7hw9HaK3noP
2gtrHGHW+zB4LWjCKor/KbJrYn6KxiQe4enaWinadgr4+1FMtxrPv0OVRlo/rUwc
i7khmVaJSOBb2x5EK/bZ/vOlqbPN9YLPhOiTYRBGyiUdDb5thsvwapFxb4fpYfF2
Wf1tORCqQj8aNmtNapLE1FOzkYFQJ8YInV9JhBbCE9kqP2yrBYhRdJuZUecttw6Z
oiPuzUFhWQxwuAxVLJrSD5uZcPsEiS8eaWjsaH9zbwWKkolWESGKeqsg7Zus2J0F
LP5og8iXP9QYUW/1BVkYeIInro0EcWgr5ga3kRjeNXgGegK/9ERl2xSSMMRagL2F
cMYzFT7ukjZuyC577+xPOmgFmb6npH+sDNqWnMR67J7wqIrsSYK74yVaf6k2yuiE
jA0jceEkzaFp3k6T26aNJ/zv5RzpOQyymbp+37NJdN37w8tcXFj7ITZIuwwUhTaM
4+xpFqHQhw92NMZR1+MhJDf6e/0nfRGJZYBL5kaEKI4gDnAtfQwaSwGhI8OhVpVr
/g79icnoaIzPxei1lR4e1upgYEzN44gHpYAsHUgd4+//bAUpjse0B9LsMMImmlNo
rstrdIqxbZYjynTHyEl/3BSTdeALuoyZNy+DA+N/8oLAGeKv8Di4bNmy2pOUnTK2
0v23SGweIgERjYbto0K0jSRkySH+9A7+Jza8qolmu9jrCy+tpHGp8H5wQkwZ3s1K
zdGXK5RcJSEZuBQLIieU/S0TYSgwCiwss4tQE0/pzR9NVJ8J4s3cl77uwPP5ua1G
hIHYw41UWcYohtWfqgDIMGzL+8bdAyTLtOH/GewcQdDv2Ryo2DQVgUXJJMymwkUm
7oKuZ2pO1e0+wDou9qu73LMBmUC4vTMrd3iLTDV1m0/SZNOg1tWapEfohK5Vi1EY
Vob6k4zttvr2qoSvdtIszG3zXBcgnAIDsVhukyO/WhR0HIYbyh6QKn2HCJCsR+0t
I0nn22QtxMxpptqLw5I2Sax98PKYr3cuJdd3alNxknZK37TnBGybzldW4nX4/FYs
g5di2BmrsKY4nonKU49uLVEU3Nwwvxs5ce6jjpjhXvOpr+5/hQ1eVyZpAUBTgRmy
UGpyrLML3GNEgF5e0hAVVRUPNcO1AbXywOStMoAFOfSo7xxraRSHmHWlBLo6ZOo8
f3aMEtylQmxquQF9Q6U8VPHcyzM7mQrKspoVsTZxyV4pKVy3LOsB8jfYu04J4XA9
tQ808tuC3jHpLz+vv2cQ8/obgX4og6W13z/NOscZymXAmeBO+VDMDGCk/m6Wuq20
tL/CpeokXW8Dd/Ez/JFiu2Y/Nk2VeqGrQYvqP2NeczFxXw+L1mwwejAVm0bV7mtn
+CfFCMSSUykXnk+/lZsDB+MjfqdWIGLlS3yZeW6BRs01bMRRkKJvCGgKDwY72Fe/
nC8oXAVlDhMx55hH+iuEmW+wZ2qx7GvXc9BdtB6DeZBQ+MreegV//BwWeKVyGmah
cZyw9qOza7rV29l1Jg5VYl+kIcGVb/reSqchftb50V0AlJwYgBQTEk/tpAKbUUlc
8mHYe2JgTtctKfViOEmHi8EEwFtfH5A/uKET/0LU0VXlIegG0rVfKG6DWoK1HzAK
hAyWeHjUbkNtwB3C70cJExfQR2AmnCj26ZWzLtZkKuFz95p7StzGyMuqF0UEJT38
aYqZXeWA5cJMe+Fm8Y6iAP24yW+v5voUiFKDG0oBuRAz7VQhzbDhhcLAwk2wZdmS
904qbWmWDnysWnsqLoSRuYCmBBhZBYb00i0iDmLLbZxlyW6iY8klmm0MUrOA5mxp
BTGzb4lX/i9nCANPKHyD1THqBJAL9GxPNujLIyU/LCPqGVQqe7BTrLqQ7jx2ZQbS
IcaKVvQ3s/P+b3/Gj5GiM0FfghuEkaqKX9RZnqN/pe+ARNtck89REK9mPMjnzuRP
bwTAuN7Iw9Y3Zsfgs3wOnxLKZnz4qGm7/6SSXcgdWYxiwQ9fJNzqL4YeyTrLZo0/
t9AEl0yen55i2g9s/fmWmNiTZFzSVTrnizwa6T9qJQdHrfkxWMVxVBtCM+EAeeQO
PZfT4qG07Ln/IAjOHjVLtol0puj4VKJthq26pk1mKSsSnTHJHhJv37HA8lZep0Oi
j+WgKBPQQvY5PgrUsSAUVctP0pjc2CTfD8uM85yOc1pqshpkKOp4qY9ssHNo6gqP
6WmFsdbViniBdBpjajD5oYxhITuDMLnQbsk4AueQxRV42w836kwpVuN/uBGORj+C
b1AHfL9e54shbHsY9lTUqJwPPCnJXvHuQqVxmuhFt9ciASK5RBwphi09K1yhAWyf
IUly4RjpmI+4/hP9R2weLdFyp6YjHl4sjc5OKZ1iJVTIX7+1OB4JSdIBWevQoLqf
olhUCWqeIcnaGLggHbNKX4kZFzZPObx5+eY6f+fwtGJqGNCoOAjYpIqQBDU3D5N6
/yO6pka6bWyog926efBzNFhqHMBXMSQ3JbDG+pwvevDrizqclZwXnjBzf8w+y6TD
/dVNgYMYP6YR4uXaIfowenjGmf5kbpcGLze77on0aEh6HZx1Q1bCsLnK7ngZOL0E
Y/0/VMW32MwYGjKu6aNIyYXy7Xpz4xFxhUpdeYWFU65u3N19XL62ngyy6Slo0heQ
v+zorM6DszokKj0j2jLYEXh5FF3BkdyNmQoIPrxCEjxBioh9fymRKpjSrv4XVXBM
8iIZwQm9eZFv6AdagYaP/u4MDtoCaTXRnqFkCWXR+bFqmEc7dA0ZveHA67Z/PVxY
hWjJ2W2uEq2Y6uJh93V70wsdSwhO2xN/0VST7Q6U8naIhary/fr6Yx1QVoR0rIuY
6OTh2DlG6rppFKW3ChkA2zvg0N+VBUBYMk3BUt7A7OJX6wm0fGcifQOn3utu0oUZ
E2Hx0zNZzIlBWRwa/oIhP/k/PkS0KZJ+2Fr6Eyo1k6WCibmSXfB/xLRQRzuBdT1r
xSFqhs7nvVwuGw7eauI/rJtHx+zFAh2ekOy0p6/RgY1KLYaHq8fAgX0fPl5xW2Gn
4wGndXjCTqC8TPc3VIOiRHW1UZAkWwmlLmVpo9DsPyD6dEwthxZNwYJQWKZgot1S
wA8nRUAECXc8ZsTvtMX6krdZZE12953Pf1UlzhU5Rxn3odPNmr7OdwuSRuDdTsRC
1xgBsM7mbDTASA8RAKBqQLyj9reb2S+BWVKvFEmYahfeLelCDVTiOS0MdrInRvFm
Rb1KTg9XA8gsB3Kf0A2fOCSOi1CnDvtfAOT5QvYaCFAVbLzb4enaAqa5llhqr9Qn
1N9RGQbMTqBoIEK3wrD01PCJfp/N1s9NEqrMWrmuaLFmuAlzWaBpxEHarNn3SLiE
BgJQBWQIwox+SL2Q+kNOCrbfe8R2frW1igimomSOuZolb132zsGZyczn8Rw7MyOx
T72PRI/Zqv8sGVfAaReZYJZ2/dn2wqXYpJmzxHeoMMN29zqp/aUvzWxJ4XqYxwPM
KTfCllneymKXMQuhKbR7oor6vYRo/dzX7NbRIHm27AWf46111dSDEpDe6WzfY1IF
J6bGE6ET/6bh1j4WVQjQTlNoFCG6zaayB+kbA2xm+q4Fk8ISfYOr5THZ2OWc1jE8
4K/dEkbpcenEe45oHOpzZCxzjMOCIqpHzjMvm/KKYoj9FmuuXlOyxPF+aLvmIl+r
3Tm9tmqvMxBkZZz0iUYJ0+IiU7yc1ds2wVzAbcYDN7ahS7TvhNCwNBLV+hOXqGRi
U11bd2EfJ2F3R0x05DpXmt2xUyA2S8JxmNtQeVbOQNfNYSnkEHsOP3LVd6/yJta8
ihX3lm6CXQrfdfCu4zuaBIva99dOONrQCgqcCFfMVHsdM197R11E1VpQ8wrZEVW2
jAVGv5npDM6iHQFkdwgpBxyVnHKns2tcWrTowPb5rgBqZxl6NimJgzfraA0YC0qk
Chg+ytrnnbPWTWxX1pcwTnDLCEYrRMZCYNk593grRzabflz8BYKRmUaEhi5rqPEQ
zvP+avGIgaPJWqZ6JU9nq5LnwLws6oZQUbsVHdje29kpMvf1WMtroU4rz5t7xB7T
OXHTo/EyypZTqKk2SFeIyDVz30qDak/0kZFb3NPeIVi1fFl4At3INpVmXER9SC3K
Bu0T1BtmH6qrXRYglimVn5vCA8zbM4dGWhRbn3t0yCNA2nEikvNUfl/jt4Euk4d2
4zg4F9gi5JkCEy8wc7+Dx3+Q/5bPe1n8j3kem3LocjhP/WiTW0QioUpgMEHKjAHQ
wUuCw7gF1SdorImd1iJu2jyLcNE9FPtPqaai2iUE+wMn17V24Usojgm0vJ8Dua4w
wzJ9eypiyq3cTMIJMzjwseFwAL+KDvZJD/EMEEiXd6luq/+9JmJh/txXWqjWeHPg
L92K9UlgjUSAGdn35jCsZOhPWhBfGphTIcub4HkOhgzhbtDfMfMkn8djxSRiKJ7l
FixCcNUUUqenJsaOHgis2MjQ2pxEkLNr6YL6ywmtMPJBTPQrL10LVAZ5tI0/uQpd
yPCXOWxCElpEN7pVd1ozWnbKSm7kL+HBP26xW+cR7F9WIcQXhz/Nr1v1Gy6Z6u/J
PozuMgj5os1cleCI5cIJU6XIFoIa4Z0vY6HUwDM5yTbXZr3sWQo5ytqyECpDluCk
P5dTtnL6XHKA2zbFuZO00Ev4YLsK0x5QJ/PWeD4bLWQo+g8TwXqQO3GQ9iIko0wA
SAPJGWWt7rRNi3+bQxK/rPuLIQnhD5/vbLr0YwzrULYnpfr1G4DvlQzOchAV8OKM
ujsFgSylX9hfB+12gbGwouNTlWrBklggJVkTvoQ3Di7J7Mg7vuzRxhCgyg4O3971
H7Ey9LzmSW5LeyCfZ11khwxmY9Ze65O3zEBj4Lf4VwfqbNr9P3IMr0vA5hDFOg2A
LRuPTGrnaSA2g/qLHQwqZhVbFbp8pe38SQhTWqI7O37fW+3JUoqrs4GJlOPsojFA
6vJq1dG/j5AOflls5ix9wyHgPXZxv6z7WhvuEsb6XGVULDCsCSvx2mNldUN+EEqm
OPMcycyNqefTzLQluZsuYDi+IwPGil/Vfr3p/GIcjfZRN0bEdjUhnn7/QwEZBQKR
7yU1a1dnmY9e9IUearu9QwShmhA2zNlrtaG5KHZHEkjQSZddcZt+t/ChbgtzxKNM
CjLkP8xHpEK9yamZJc+GoQJa7klZdcwG5iE1dWp7h6FgHyCDQYBHM34ztdLpLSX5
QK02dOFjy9J96anEPUSnqQ36HMb9/B04OcuDAhxq1FOWNWzO1djzrdeJ33ej7YGt
L21LJGREM1X/MXsoQ4NW7HzABHkczeGwj3lt0o8HqBGB6NdhQLVNu2FWodGR0fsF
18kPSWpFUPChhN6TKQ7Z0pzjlT+IQ7cuJFpAN+lX7v55KEIH6JdSxznl+iMx3I2g
0I3rEh3zTI38ZDFqbnS0e+kePJdoDLFrjNAvGLRWZ7DQvAqKEb73gmIrEdNnzbbY
9LL3oVsaiGB+9XZy7C0gWqVc6julBCSp/bc6ErDu4IORDrr1dQ1t376ZO67sVRWm
k4A9eh8bluFOq4DDRHEnsU+FNxrWkJ9qQWgT4hVbPoieZQ2eiihj1XX68Pe9TNxt
8Kpycv1OGyLG1VsRrrR2Sx6Np6XtFOJhgRufyaTBgzMzMQjiCsXtDqhTY+dMN/mL
vUHN3iqDbBX32fhzubGxz1HhhOgzV47URS12SQuF8wAHBsbTS7MwFADujrSw+V7I
ob1mCxw38UEJxsswk5l2Q3HHmkFs7eI/sTjwLcZWJilgDq4hv227pJpeVR6UNUum
5znR/QEGR/8tBKSyDyA1efXD0EHCd5vO3+uiuOMxXvrSmf71eROX5EHf8Zn70fJb
RSCOKbTtNtpkoqua/vzrW3r7XyzaHKj9VVVyVID0NvvZtkVl1+SwUHbODJnMTkF6
RfW2AXokyO1HWCrp7136E+GLkwYV6rALMo4ETzfZAOpic9snd9Di0Cldr/NnIMPA
sFmnW37CUS8IZX6mI+1vkKHSYqQXjiUNLDCRbwjDBUWuUGNRJe2p8bAcmFlEAkQ6
CEQDJeO7yfNpGn1Jg0CsaA50LpMOJIpzTmYo+R68bR616gwTyRcCL+G8S89Vv9cW
GQ7UJ75WtYs0C95GRopD/lbQNcGyKnFJ84pyYdW7SnY2GP9PncECkVCFlrgRnKNo
D94xG1mJGIu8yqeE/jG5T46NSUpLwZ78r/ZLy0pc5MQvc59NdqsrB/8euCwIAJnj
/azawG0HYm26ZeLFD5bGhST4OqUmkHeKZf0FuR4IAFa/YBosLssUIp5zp4xUd27p
AIkq31h8o/GJreAYB28Mufbz3+Won+if2ziMmLhPAhscGEQfm211xfzW0CBS5Alh
wvO09+eiJog4dz2W85ix94mME05Js1cS821hDpZhDJXBQ0Yrjq7neqh0rUYmaz4b
e+p7OzICuxB8gEvB9riTPUFO+FfGhKhFEwlt/vBUAxPXs44pkRDKDeOkmCrRlOjX
P9HhHwSaoCACROHLxyujFcYqjXf9YX3m92UJ+dGPCdiS6Gr4y+tvgtJDBrUTcDe6
Ex6D2588g9CIonALL2wlUN5rpe3r4dR756nm0dB4OHjcx7ENJSiAEQxUo4KkRAOb
ZjW0PnmXtXx4fyGp/y1afDZZ+7aFUkgCS6kRaD5j653ZuuJzY7URhx8RFf8aoG3l
NXhSziny+AanVqR6vn3qWHjeu7ELNnMuf14p48Lg1lYf0NK/vBLKD8nSZF57SX0M
Ba5e6bITRVLnb4gvV2VMiQEpo6TARx62AJrWUJMLLBFXBqxBP9xdgj/7DStX33uP
PeMEOanW/KgSgpRimxEgXzJ0RCGsZRtYCVCNBscqHDmiaIF1y0swMWditMA+BWdp
/GMKOugRRkfbzLNvn4WMZAwJT6Rpiarh+SoE9YgQuNtvAoxfc79y+5FEuwvpG5BG
D1czz+9dKmPOLjUtTPzfvFoHtBEmfYB79pjr6JQkXYxat8sWmtVCUu3NySbLQ0ZL
DI5r+7Jvudrx97tM6w2fXfk7Z8pUlyRVow/JpMaefmGQElSJorrTLZfSJYNaB8Aa
MZyXTLqVr67ohCth3+DhuPG6xZvPC3p4Rj2f3J4FPH89hJaARvQoUBH7ST4HK73M
Kn5TJDuTQAjbc5WCOfOewblihwmOGtKR6zbQ/Gzj6xE9EMGB3VTovDAnHqEDXj68
6x/h08ty0iDgSAsAZusf4BmSwO/1nG7HL/roaD63tX6FZp139nVsoWaF0fYzqrFc
eIvEVXqmzFDqxsUUe22c6o6kSkoVkWV1nSnBpDybzNAoHEjRbZoeVKqPk04VA9wN
R5lg2igCVDvlDnRCyWI0hLzcJXVxQsoYmkw46ixycSADzQ4W3iFIGZZKR/zbgn/+
JIZ0HCUjuidlSpoTF0z0bBQ512b0fHfRSv3Z1hN7GKqdwOHZ0mTfneDciWSRv588
c4x7ZOPjG5SlVft4zSUg2K/YjmQzwOxik7gfLN2zckkikatJ3eDTCPt2uU0E7Bwf
XrpdcTZJMYKMa1BaSz2JPmMiDUbbmUznbz9vP56u6pn6taK3XQBKRkbMmEgDvks1
3X4Sdp2AyxE4QQNwMwqIqu0kaaBnU8pYDeLWGfJvl8xIEgdnL6ssX/Trz2PYcX28
i4Cdp5E9Eh2BEsX9dkKsNsqGEAg6T62rN6ICUBQXCbNR4BOzT2QpCHl3WADsfaPG
VW4mioExNmy4fw8sF3+ay9/V3URzr0S+WopCCt8I6n5JDYIV1w7MdINYWkImNmzN
E1V5NjNn8Vh1PreXkEMEpLn5eIhA7L3UbWBXMcs+gAC83sMbfRr7DhEpQ4lFzjPK
Sdvgw1wUhhadi0zNNUaIq3VHHhL+o6VXi7wYDYD3rDTW4exF5QdyVOfevru3kRsI
XmzETSlfSBXNI4MNKAu2RGI262oI4A0OOsxNL3+OdFCDyicvQ2lCmHdWlWtmAo+Z
KPKokyKqCq5bS4UEZL/QyYbtCGxucLquucYWKfmDZ5Gb6ziz49D69gtzoNYTKAvl
Sd1h5zWTwD76YnpCuvL7+MWQi1DWIwvjzIFL423heqV7w/ZLDqVMs0MFkQYJCjdp
e7VMkOSUFcN+wuShH+qmsJ7yiu2Jl7hlOwV9MFo2tRu8wLjEUlXyMZo/n7Hmt0LT
zPR5VHrJI7kv+mfadBzUyjKiOcNVc9KekvzdnK+jYi1HnyNG6O+dUFk4z8SXX/Mc
ZqZaDv2mlmSeqqpHHE9CYq4W5bK27xnbKye+46Mw+e61pLXZ8Js12OoAWj8P7Shj
fVmxfAvBEo9hBBZ9Hjiv4VhXUUS5gpXmDbxjtcV8kyGAtIC9WA9uHVebUPQ8fANB
jEzTADjO4OOazXayAHCB1utkp0NbSNwpTtlFDTgUNqnnqcvC0sebSAIMz9m0YhUz
7du4gNrkXqvTevSkIfxEFfRTeRqASDUirLHOlhriM1SSHQSY+lMrfsDSNM8ZyhLw
TmWIL0Sx8wvpP+0fQvCgTAneAfagvIgbDbMiEPj8sqlSiHqzFnLRLa3k3I3kes4g
WEV0vmR43bEL48VQptxZkwDZISw+0+E0iBtDQxUsxmNEpw7Y7lEDdk5/11BgGqC0
rr9o57Y5VNx76fPOdCHmJ5ZtJ/pSzuB1ulRCxiNwQrzKeygx4jsGVmOLhRNlm3Ez
yM7MRAz+6GoUiJj1xuQRJZS6IXkAdUGXrtu2GuvirN9gCNbiytwYgFbK5eSJW8PQ
+X1lVZQTDKvutoA/d+ki//eMqHvmWCAJP55w2HNUKl+5nXVB2EXEL7cgRat13W8w
5kUwLcK3qG2gCsPxpTeQeQiwMdhcFAXiZzsmAQkZXTePAQcRuVEnREn9owiPczTt
GUVni2dRLN3+twlsweQl0/3OE1MLD2OCis49r3/EVnFZzbHR1R+Ichw6kA6uLMck
k01jVBUtmbtm12qG83bmgE7HAeWMor9QN0EpLsIjoR0MirGsE8rahDPAj6fO7p+p
XMFkd/BPpeduW8EMrYDqLzzjlEc4A1xjlxZ/bnIv/ZBHCXIqNtgOPWm/wxX0HHS5
/HT5J8z63EFmJ7NkCMK+UkQusXv5W2sbUz+LmUkzpYP5uTBgUXPRUs9ATTXoe2Uk
fpZkdRwvDsy2FKkj2mWwmV3Oy6akItwKEjN49MM1RIiFXZw0Heq5B29cfBh+1+ed
7kfmtn/7tQN6rRY8te4khOkQqq51sGLMieU3IMvo0J8WMzuAH2oN13ZKTU3QyplR
ib7fRGBdM/bXwJ920JWAu4xACp9AJVuy6RAnVRbyEKzHmMYXX0rXqMnEz6jylaLM
Tg5FJTqLx4hJiB4B6npBGWf+/QJ+56wPBrisz5D6pei6QraNyj8pAuvobgfsoLkP
DM+k05PlLLDnprcmpw0difVvXn0ZQEMkuiULNHu9hCFYq1hs01AG6Jt4TzSO4Wzi
ISVIm8R6x8y46mzy7iL9EkvU74MxvsH8/6Y7rqMHu1TSNtEAitrhFFbBT4ZBNfyq
+5myj1GoiCCjYlVviTznt9JgEWtLYE3yyYFUxauRPWFu57FOFyNIvHFCxpA2ToXj
UDxcDEaQpVGXbLdsukyx1PlKW//Sb0gStLQizeMIZC1raUugt9UWzzd5Zb99V7js
bQq2bhd931F2g23Hx3Oz3a3xBdpGRm5qgsxWlTivV556EO2NvYkcrMcuub4Djl92
6jPCD3tpFA+3OpJAc5VYrmupPHTzTuLrRjIan3uaNlqvUccSudBo5Gk7g1w80n3F
pMKJtgr0Ysjc9vxeqjh+xsxVQgtonu8I1IXcc24u8qiTQlagmqOCHw3qswsiRV4O
BjIjNV8h7ActWauxVGX3cVaC+u6yzS21Vx6N6HO/inLFE0EdDQVchMBWw+NqMWqo
KDuwcAk0wG70u4EmnSRRl/AIjP8768IiJ5ULCS9mDau7DYD6MafEb74v0JgB2uGO
pI/IkPIBk3qP3QF97V4GKb5Dz7sYkHrvRL/rRbDwfwrEJbX7FXe76NQJ173cIx7U
skQoOL5ePbS+wFFGFZmCWnCttaaEUFoN21coHzpsQG4ppIqOOl+iM0eTk2Thfv/V
5jK4zRC3BTNWFcMOImnCWBCs1bbTB6y/p9IulUn56wFbnoNiMTJ9d/jptlWiHObQ
4sdF1bwaFdZYSD3dtWiFqYJGyr8sYWSWDFOq7RVuprPiYV5mKOucxKQsDPu3c1je
GzOkIywFRhFy6HeVVcx6308voTafUUc+G1e74lUIPfKUHxPczCfa/DiH7zoxkwAV
Dluk100lMQTGwpYxbHYeQ2RRZicEKId6NAsbxDESOxUQavrLM9uZF3Qs1tEIxzC9
WDpP52yNGUis7/CH1RAVGnSzmdZi5WK4bqRwidOOydvOkQgicp05XE4jSE4DkAxt
taqtM4TaZIR0XPkossCCx9ubDt7nV3q0EEkC6mUY+HM6H4CbEWi02+nrHztp6M8e
+1M3hV0OWs8QYwViNmOZaXjyVdbASuSsAz2pNfYbF1T3/6tJSo4AQjnO8pWrkOSb
mhsMczQfYnjqEyoBDIs93oQi7T9dSmh72MAWNeyQO4o2hRWjn4aUm5MQAZt66oKc
EtI5ldCTELQ7GG1bQc75z+SateG2v1tusnJcoD/FcE+EFeKeIWCvaIaQ4PKJPoQ+
1EQ9/9eJEaAaUsNzVLnFP4rKhE9nhKAEdXj0WSzn2fKtH/IdecveKy2J58O3LTWk
nvUV9okK0KkxIeqAJVxbA5wGh+wNn4eVgPEhNINfa+CyApU0mfkv90TR+XDbaeH8
mi4bmc6r6pdulfN9Ipiq/uEFHr3S2+tVslSHkUM/mBDScMi+wW+06kYIMlCZXbC+
+Ro7WhQ97U48shy5dXCnlWwyP996gPcEhdTbly6XLEOkduhQwMrVqiEsTLy9n4bf
s+M7SZhn8xpNvJK0cnNTF9ULmtRs66/vSsxHK1VrPaVzcfit/7Fd+3TOvZIuvDkq
aoaYVD0AEvkWyRD+CwdKPItUAA/taYrfX7/rtxGoQ9eAwQtMhTNIOb927Cn0xU11
yVShrrlHJ64iftn3p/bOdhPYLGejgBSVaAKL4C7bZa/2xU/5u5iwgpXTybv82075
2pDcl4OTlKi40dZTOz/gzgL3fUSoNd/33hqDpPurqNF8516s6lZxeCPG8S1hI8+k
0wawwqbqNoeFQmX1gnFJfK+wbzhLlo9ygeI9LF+XRtICGhuRe5utQsRHUTXPe7l+
8O/QCccgre5CpAM7j+piMEfaWxA0TKrVCc65DtUJIAp/5BFttQ+eX2bxMLNi+Cdi
g/j3J8U3Gv2D/PRAtEsiYLRfDY+u3HAuNt+PIaJ2pWDbm5EAP2tDpLs21mi9kjVu
VRPfTTwcfJrS1RvKaPw61I4XVmQm2h1+zkWH+lZhLru+vbAXKEuIj7TE+3Xdg7T8
4XMfL9qVFWZo73k83/xidkGG3A5a7SN0uV2MwaarqdoggF+T7wnzQ4ewdX7lx69G
xyDMPv8ApgOe5bW+a8mucHY0vJWvhM5yLGEcwmYmR5FQ6owXz3tjnKlWvI1jogGf
1SJ0r+2jE/FwGHSvoyYw3DOElHB2Br6Z1Hj6phZdj7N0K7egtUAbs8/1T0QhqBxz
a5KcV7pV2KaRRTn/J/rCmVMLtt1vijRLyGxV6OkvYSLWRusfr5oqyNfTWUAYdPbt
lachfA3kFBE+jdEDVj9XR/EezeZKDYfsnZ7XWLfJGOOhmRVQIMRWAcHmvbKbTcA1
0+WG8xxG6PLowS4sZVEU7c6ZjJujye+6fdswHW3PPcu/P0F86tX4NaWfxkYNIXeN
WgFcnmyXFYPBsp9/5eNXD6v0p9PzTVaLJGhimAEr/+7o5N6SEyudyzr3Tj4CW33M
2nxyOdSXxI9GYolHTXpw8HqXtFEmQy9mIgejz39DJQPhua4Mj0FLbHo8WOQf9Ieh
kpZQLLy18srMk/31kZKx3JWB2x+qiaFysCz85DdrckQIDckGxkxxujHK2cDvCHK6
2D8XEhzfxl9B9xDcVLlG4eZKCioKlRODlyt7lGi7cEyKytt1pYxmRZ2cvS3Zu4RB
CnfQh+aJ3G6z9LPwgJczY5788/SlWUcQAgrNM+f76Db2KDk9tN+D5fuZfrjgt/6a
Yxy9HHUeH2ZfrRtwpcK7SdwoHcVTuCe+DLFAKryVkHvFgNUlAPy3IZ2DVg4i6MtT
7r29qICVNTjoAECQYiR7qCFpdlmMS8cO6Pt+B7vfBKA/kv/RFwMlORsreOrK6jLi
KjgTGPsCFfC3Wp+gNiHEFfy8Qsuxs60xP/g/KaE/OVT8vzjKc1Xvv0abDHUd7wvh
5VC/8y7ur+6wKPm6K6SvrReaX5lyprjaTAVNXc2VBUstc6zLzuepPyMTjC0kw1oP
pu0VjrCOskNeHapVtLNf6J5k4vFdACPosxPMq72S0Xc/u9bDI/DjjcqCTRKup5cY
Fntb0VWaIu2d8VoGBkEFMh/vjuO+YmUF8z5ZZhUcDXm6BeK+jCre4LEtxFFj+nb5
LiunkSIlTSgM/W3A//SFax6j/x0jXEautZu0/ka8f3gjyfrTLcfrtISB2Yt4aWR8
JH0k84A8Cnzt11slRSwGRv7MpEotZYxkEAfeHVAhNaii/XGinO3oU8YefluaeEZN
DZfOhnXdMViUkIziUEz0GZaVOR1FKX2OB79clQBPDKeMmfMY9N0nq5r9WCECoxry
vcY9YszObjeLkXmGv+5cBqd+ezjQUSZWfGGCDsf7TyCERUgEn6jCysosEDIvaCjE
fxckzipZ9SUZTMbFwVZVHdGVJ4xuEqg0kiBpapFjhsGDBpxaCx/LockWzkQwZ1sX
G3Zy7wIoIPjrqlbkvx9znIbKU0NXeTyJwfZYjcxVJPA9LxVdhCADZXmagZAVsGY/
HidB7p8/Qx0KQPnHh5nJ09AaIMxHBAbYmfc1AKHD/JdMFQoagczXyTc/wNYuH9jL
rN+qIb5Dty1ZeriOqhoXVWSfq0N5VaEC0ser3x67hLz+Yp+KfLTZlCiTXl3tqolL
w6rVzyiyLUReHECndT5aRV104IcKVoBkdX8oRHkbAwSq83tU7VHoPEYD1c4EOGIB
7aJ/EE+MO910ASNtTTa0Tc8qZBY7eglQwqzVH7DMO9W+waQY8f1a4S4UkxZLpcXE
rLMcqc/O2h+9RCOno4WQl39/X6XdftESn/oQO6DdV/BcyoaXk5jc+ILFt6cjmhdp
UCmPkHPENoLeyZaE6qBKQ+A11iKAS+HmQtujKY+5oSSyfBxv0zYWgIXJK3VABVTE
E1mVh5+DPUeDBbClQm6sETp9oqaNzN/zfbAu0ZlLjykagANRd8Rz757Rx8d8/rtE
K+oamesg+hQed6k5moiKxuKTk6M2aks43AwFSwC2Prvgv28Bd2sUASZBH5kz2S7c
2C6WMiX1CSGQhZNN4OmHgzWz2GpbLsBuPdFw8F3USg7QbXgy46MBxa3bylgX4aaN
VyHrCFhbcSeQmU+X3lioSHQmi/EXjse3dFuNcBIty5VcAvBUxJnKD+vmLtic1F0P
U7eyOKNKsfCgKp9e1CeEcnatt3stWTkU2x/1pfCVp+eUchc4z3eN1f8dvcK8EtH5
WO7x50ZnhNbMZ0R/1mX2KWz90jmZjezm12bfDQrP+9Z8Zm/aEfFVeDObSGMKwG6a
/Z31bgzZllfCghywQijKBzoaLq2/FeCQWY4l5OW4CR+Cz+/Nvf/R9YE2rAvYqGss
tb8atTpBfHgjEUlsjAwjJ5CHI+0P5Z1nZsxFKlJr4ivrQzPJjHmJCV76A7oOCCfY
jQpzl/4Hf3vmqdRLkz3k2fHSzg5tmIwLu+e5jWHT/nDhrw7YqrWJs5Z/4OYB85EF
XCS62SFy5ExspAi5lFmqPkO/MPGe8vDtZRvz27cb2RdnBu6FhEsiOdRV7LKb2b8q
DQ5A6uUjOtDm59/NxN9AueypKoXxSM8/ghnT4ivIw7x3PNJDcEOp6PXv2SYz9BLp
miUt28aCi9xF7CUmv2Wo11unO9Wjgeh7EUUxVcDvLoiTZHJECR2Km7ETIRA7uHWr
jTXW1TnaR2A4kLZILsH3hJRiRQILrUM95UfVmXhVaLy/0NBQ/6OB5xVQWYAOmfpB
/6zic2OABlfBTlyS4d62q9Wo2a9FyFf7ucP9XgQIEshIamWBbocAXNJ3XSua+JFW
6OMY4Mdp3jt543UPMTWXz4IHEoLQoHukqm/4wbk12MaA9Uq/qeGIcyLd389qsqWR
f0qf1aIncn0XBekfqjvyKQG1sPF8hf6MKBlAZfmKbkUhJfd0rAs6kXzBHe4CHwQO
h6WldabNvbdpSuThxepxIYyRt4acAyOeaeNOT8pezVCGfh2DxZt+WdlHhDZx8GaO
EmVsyipRvAjbqRuDlAaidf7RTDmY9E2StqpSXeogX5a6H6yv6RNK1kUXhVZA5eds
duzfkodhbHVW/cNXlUXBUdYhMruu6vz8EvpgmJxYd7+99NzKmoD2QJj4z0wYlUpJ
75fGMRxh/SBrFFpJKWHIHPb7SVO2cWXRdR92ACYMz3V3Xth0g3TqXnmdZc70dGyZ
d6ETdVOnvj980kTU9XUEyuaFDaMC2jifVhtcGS1R/k0xd8BHaTrPmu6Rtx0HjRLA
B++IttgQDXpPnaZA87SCgKKYovtX3VWng81hvKCSTbBopZ+4zDKZ1JkhmQ3qInV+
TagB/N/WVpP1JFOMIdeKd6s/ONmmo+pDFKmc01pWaJSJOueD5VimkGQTRDnRHEfo
xfSdBVRuFDMT2ZwDSNQpKyFoq5i+ndrRZMUjm7KsTylToPEBv9+XlZ1HzB1Uim5D
PzLbA6nEX2iXIUE369mLD/gcMVdpLHqgR+oX/06TtsymbBntMnK4DtB74jfyA17o
ujvJqc6ow7uhWJl5U9HdZpphv130MXTuPER64PMUIgxOhVMuVwXDZsMLuWKNVbiL
iKdKS+uCPJo5Yj5GCUhM8lm1kEvoOdfMharjM7Enol6VdMeCEOWLWKEoNy8eRIqU
T1Qrx1HzE/d7NTcU+822mzWPb5ZeKhZV/MuVb5M9kcAbHJjyPfwYdy+YQu7RcyVj
prbHm50EBW3Iy/tSldBLb9mIuRcAG2XVaVTrIjwTU7Z3XWlz6ym8mnUrbmdhpvTs
TTlUkRVORbc2Ue5Yq+qFuXZPOeQ6Dp1kZPZ2M+eWONxO7s3g0QEnyv2wVSlgXbzG
7UtoWbVs354B7PR8AO8kuRZ4X4c+VAkKN8HpGkKDq6R0MfkpZMb0aM/JNVpbj2QU
hA3gFt8xiccQ+nyhPEsPNB7jnH76hBOIwqtCRWxQsgUA8NAMtQmilP8wEmfBVNxT
UvZOVFrHYIoJDL/Uh2j0qPVD0uHlRg9gNUodufJha6Ha+8Es7wGWaiSwkyliRefK
GU/KXlpi4SABQCu7j1TQYkV5FKBq28aGvz5dSVlBqx1Cz3mahW62mLD/tykAqMTe
nZf2NYUdPn4068gmMeuoMBVxeyu0Hfz0b9hEx1ctTy2yYS+GtiXslAh6LdyOp66o
MGXSvhJ6zy9Gv3zczLNcqPcaMViYxqjHurOfIZW42kPVnslfe02xbBL/dGoKo6pR
VLqjdf6kCzOAS/S48t3W7WwtaxXCy6EMajqTopTfZJcZ/zxY0M+5Wm+uO7mbDrpi
VKc2GXbma0F54uZZ5LHc6ZUav4YD5QbG88cfa45GDHef7DJjm2zJdcGxkQa/IQT5
oeg03TOX9iIj6pGNBpd/eysLxsHKIrcRwuud40dAYUDQv+DEbT6NrtPjWE3YB8vK
SiTL0hMDT4NuXhVdUNeg1pchBO6Bw4ZFOh7xJIUxXijEniwVQSZBTCdkgzLupK8A
f3/3QgpLYmsQ4M7YAEve396W6ha7nhPjPiHzjSVLRSPM/La8FmmUxSRLVqYmHys4
DUmh/VH8YpqOBQ8XLhPeLGdwsX7+uE/m7ePQjIxhRvhZtcvicycF+HNucnXdmrXk
9uwX6l6GGQWSDVnISXZ6vr3EJ12DlTYFe2f+JtoZe9/cLCI+fWG6Jnn+U3OkFCkg
ZX53q6VhvZBb5wlps1lXzU67uRuEIUuL18IcRcXKhSB2twGN+Kd+qA3hw7Rh+VML
d9rtS4ndzzSUHKVt75QZME7prBH+1PbRk4u+pMxEeHDraZ89QwKUvOf+QA3QOsXq
wluHtUKE9Xyn1zsmD5u+oT01cZQP5Z3kw7LtPkn1K4KtM6qLjMDLkCgXCpaSi/NB
fx7uF2Z1eXM7P/30OGDePHcaDnCGpjmWiALJuMVMtHkd0MhUmjhGYBYNlpt7KGdr
EHFmhaZ6JQvUMPNTEWXYppXmHpdGlLDnd6HIjDPOQDzoP4RF8cRRzPgm/D5O+59r
O0YHgR1zWQjaYHyEbxqDjz0IBiLWqX3suq1dez/lvVR+O4XaV9Ya2PQ8gWMEjiKL
HaMGKinRf7XOkv6lhPDQcKOrh4yI4LcwtBGf3Pfow/He+e9ovwLDzSrfC3R8voiE
tYeLNc0I8XfbvwqRyfVuJMGZMnmnPwLQFjqG7431k21KyYFg0RW92GNVIAP1DsVU
zD1g/R4xKcTkpZXln5ILcwbyI4RGPlI5ypCt/OJ7d3caGl8Zl1Y2VI3sAPhblLHZ
AFwhDa1tGaBFiRhfajDgdfTtIgDkdOCdend9tM2pNSJwirJeXIGq3wNqeNpKLos8
KHXG/hXQAL0oQY7IEXcR1e+lZCsEn/83KICLJvtiW8skD3VkA7b+DYaUTRtFbEbs
dlnqc8xpL3+C4kmAe7kPzXfI21TxdFu2NN/h+0Ih0QLvo/XSse5j6WhwitOFd90I
9Vmoy27+DUNKwhtRIPkfSWRHsYd1rnzlHgwamd5D7fYhlfHR10Dt4Rs3fpxFew5z
1EUfU7+j4kRaKticY67ikcuTGMYD78BPPx1q2Rl5ckjrslDEttjohwLBOpti3VXZ
E+9CU38CKxidy76gWQYFmN4/PIwgUTIxsF6vmPH1OtE/gjkeQ0ICf9FtwGZHEe8y
YKsLs5PYmha7Olv3EO3a6nXf5d3HUEJlggM46mbjX/luVEsfni3F3zbARSRKPzrR
M0BXHASkVNkvrk7KzYekjqEBs++hFgjveo/M2PEIBbAya6aNBGG014RPLPJNuuqD
IEFebNZYjj/t5PiRZdRO8/f0d14k0ghn51gSW+PD9VIKw3wBCu0LbQH/cxcLU6zH
Djy6hsDoqiNz9RzyKxE865rhohvC3IMS7o2ugharkIUgnsOu+YESBT2qJPI2IYTI
X9SJxMdl6rVv7cnpHjvvDZrKaBJMBrce+UITMSd0FlgVYggzH9E/vRloy9Hb/yiE
Ca7BoB+2v1MOf6RJM2fxsOW+C+ZQYD9twg0xtFP6hkDH9ibmY6WKlKy42mOk+Iev
XQx6XXIUCWN2WcNLAfQ93F6cU9VSo8ziwIK+m0iNPvVEU5Jw+nOGU4qRNywoY6ZL
HCihsr/akizwT6bCFJqvAal99Si4wT5oiIpgrUG5gghNsbW1+hGzA0hnE0/zgcOM
rTgqCKT4vJ5tnrrzMOzrbXyCiTdT0NsDW/UEOlM3iGl/jgpTEjl3EkTMQX+/Q7Af
+9BXg2xBLAe9Cx13t+q6c8sAqYSppIeydJH/pKzdRbrdRmXmRxULM1CoiH/3PK0Y
7PgsB/FSxcceTpfbeZmB5xE8jlB4WYGpeqCqBHwWfIFXO5jE+tYjR3Vye6+5Xhp1
Yjsddwy3crowDV6IFwsdnyphkQlIok6fbsMJ180lZReHYSDYtQeN5eZXuVWgPJbS
IPlsRadwaviOcoLKre4V2mdZn0PvGv0vzXP2D0XoFQoc2x6b6zPBzS5Tr/VYUCgP
XBJJ+cs1FeNOFGprIWpw3B3zbInWnu2U9kRWzSEuLNRg8H+yhAcsSxbXPAxsEEsr
1NsVos1yzyeSSMrWoSeNkcpvY5NAAai1yW0rAAlaQvMLBCPvHAzYfcS2lrHDZ9O2
YbQ+2ADrtAoIjSw8VKXGOsbHf9d9RyUHmGOz+2a/za4DNG5t1iEG9evy6Vib6Q0A
IqKPftv3r0mG0pOJySf6NTxLi3c5KJZpCP6MUdoTr9+AhlMqXtNHkP0eKUR8WMgW
vCcaPVBWOLcpPOAOOKQrZgOjmpWvBkgfkfWjEpaipez5JKqRKRMdmROCslGk1rUl
XlCKUIXYTGGexWGeCGS36yqAnvodTPbZahaLokr7rPcrDbK+ginzPTqD/tDVXmHL
za3700kxSPZKCREB6eiCoOZRo/e8nbZwC4Nzc6orT6qp00e6N4n1qqr1J4FTopwq
pAWp2JdeOuEg6JE+FV7eg9kdEt9LqpKVEd3bv+s9qHvmASOz2/fBFQoShBC77Z28
xaNq61yzOrNTYn5ukkq2gS6lpK0vj83NOkkBsCdQJyTfYueI7Z2l/HvE5peX5o8/
6Lc/lQ4hNHza+poiB0rOso1xEsOAjTJ83ZcD+axX3mserp+lvVEXqgld9X/ZMNCy
8Mo3trMCr+WmcpEtFlkF4ujPDu+5hgFTfRDQNHpzTCZecmGP2SGjDQd82WrYl52V
Uwuu0JSija8IrKjKg4iVCE/4zyHZSaPf3z978TPqRYnGglSL6oES41fgfpR9R/0p
dP0+kP2FnBUPY2tezpWWyeFwracn3bFFcigmjRFOX1xryXZgr2hRwEe7l6mPYNJ+
IdC2AVUhYPrP2QkGMVEeev/pBajqsUxdzdyq7Eh7n2wSRxoW7k6c+8jJ5UsaBQMo
maAXwMqMCR4dN+Qzzn+leckxXG222hxrc0WuWy12Bzd52PJu1o8P2cmtoQfPGgNG
QgO6p4MO0oSxn6u2hHwJNY4KSF2Ar0muqLdYbfDEwXY9edoHH7tHPPg9ABim/uMX
qqJQ9WT1wFfe3GULbTZMj0D2kg3ZQ+CVLWmceXPD7vFLQd1xjPe1egDiiDNJ6nJ0
YylHJTZ4wR59EJFZqrchT70m5V24UwNn/qo06638gU6t/JXS+L80Hf6JA9Imobm0
cs/A1aW/tbpx8FImMHHBSH7maGHLxUDRYstXqnDVFBSOD8NbhPSa4SMrpKTKepGq
J6QyaxL4NQQpMBp3WzKX7mYW5qoFvTpd7C+EcMDY5KC34lfEqA3ucuugead/SHC1
gHSJR+KeiFssjQfIAhXIqhTdFaVJIffWmPqN6yYyTTEeYiTa3P7f46Q7EZ3sjHN9
RdTd1KiD246y27Qhq9ycqvgXz+pq6aXOuuT27ePQ+7uXBrma7Uf0fdLMYXX7i1WE
8hPolP7vauCszMEbmOM4NGQTjV+VGYhrA2Qi7VdA9AXPId6o6SM96iqNzLvriV8G
TOEpVn0rvceKcSEmTt+BQlDKwPWn+TEZg++pLFaYudUIRvKpDWBfi5knbyFLeP7B
UMhcPL4RHPDZjeVDScviAdyvNFBlAvZ/eG87OYtEQM3SuA8PjacbnpMaxPwyYZqk
n4kN47uiDWi1MYMgnzodEa23TsCIM4EuI7P444ejmQG9ZEbL1YM9yNCYtH7ikxdw
8320vr1bNWhuBMuR6ElDw9lAnTJWSdEszyg+gApRVmqHyt5bK2bEmrrQHflRaegr
KKSIEPNWBjRnoo5HOjSVZ3meUEBGR8FLwU7L/O+zCBuUOJ2ta6qFutKKr69uRezU
n1+i9N5W3CjsQQz2dnYz82WoHK+zibx8Nj8gCbPpcdA2w0lAtnq6P/CH9CGWsYM6
5CP8RiRNcDfRfCYx3p0oryyLuSpk2135h9vhvMTgQo7OsWn/TOLYBg7O6vk001TE
U64joKisPYGDnuVuNZZrydhv6W7oagh18GYmozdx1/Jx6NI8SuCbaithI1SZt5aw
7HM+0RXPeW1/04XSLApUovsDX6FD6Uk17RMk3/IP68nWbbZQxFRmGCIbU5TbrxSf
E4OdCkwcfaTsX8X+sA5SfwNVMAqBM7JJLWXAaGT72SBws/p2uKvpE1ZWcGbPyzg9
I6KeAEe8XH2rSRQSLrWpxGAGQus/5iagl51W/1ZCRiiIlNTp5T5956dRwxCo7wub
NcNCPwCHtfBjXb9Y1yqOUB6I3PmizlWdCwxI/+87020gQMARuIhq26DRJuPuR85P
76oDd7Y0U8kIAgJN2zDZ/T3aQnNF8icP5EsQk9USwTX7I52GJ8LENheWNNFiuSzt
xyqY8BtG2+pw5aNMGl+oJHEw1ieuvJrg+LI4Bt8Ow8PbYD5yVX8irPe3dussfb0n
yrE9/t9lHjbFncnESvX1074QML3/bdxyyNKNDMOCcJgnUEspiKOSVgkKg9xqfuQD
6xe67f1ruUcaoq5n3lXyJmbkuRFYctUlpbXFDYNOlFWvYmeJ4hFspTwarDFph6hr
3GD98HFL5R0XgYmMrzf8zCQSs/AnZvyzGlG09GS8fZ++8x30ak0SAFS+o0PEesmW
9Gmx3TxFu9+BA9rDmsqNkwj+lrESR0mPiewb2OGmVZyP+/UHFeFw3BYQqU5d85CV
sq+O8zm8AwYYki8ZaUGCy9uNoaY6h/z9K8M8hmGLxuCtE2At1AkiL7A3moy91AVi
/i+yaDZdX/36w6gTqjrWmf0JT8d+89rO4wdySRyR4VvcqjzJWMJI7TSLodOth++9
JJ4B6VNV/OFOS2DreDwHTZSQlLawqmT0TKZqlL7ONh1Yx/xuylK3tAJp2zk1iyaS
3yYkzzGuo+EMeq7PZle278eUCLNWe17hm4GdNUE7JeoRs91TOfO1jpAgfPwP4lxb
6lERnPO0xKGzlICBZmKGt6eAPHKMDRSxgSwZG0VlqI3SvyWoOVXwaCVsHk0hMuyG
28k8ElxewnuaO0IDBYMUrAExSSipVMNorzyLCWYYFhuTcTCXpAXnKnRlwgSxbHoz
VYIcPtrMSlNznh2pwR96nVUTlUG3N1hIrJECp8cp9+TOhQn2dIO3gX9AneQyPICU
iYOuy3YrEQhu4jNG3QWeG8kYJWdxJPUPkFQgnQkM/o5sq1i/7zPynUdssvSQjzoK
YQse2JXZPiKfV0FlZeIkxUScc7tqhiCogYcNv71pjsUZ2/aytYixuBUrW3rsALYV
vuaAUnABpRoQ072wo/bGHlPOL6kL2irU7cNJtPkI+z8pN719NWIDULlvjpIkZekV
2JjKn8O+Nplb1YyaSCPsUATPzzFVpRR4MpThXfzVECtz1Dljqy+QKXRASi3Gymfz
sZEfuw3IABNLfTAKveW1XLtPoKNSuODqW1vc5J0+YoiIin3251L3kljE77QK0q6x
Of/eulQh/Ridr25aKaIMwYVudn3mEFDTSeTmu6htod0aay6lwv9jWdk3teYtPxSf
miBirNStQWEMSgO15fS8qmKwmP4w20gzkxb7gr5osqYwqW9EvvN3Ba/PX8Mvi1bs
XvC2X3HPBp4IS033BPDu8cX1x64Z1Svvhh2mHPsTxkU5p2bi5hiHCt04uL0Dg0qr
QKqJf0mPHxtnz7EUkQT//WLAOqvu7FEwJT1fXWEKLzZuLR64iRndGubZcr/gLFBi
pGiIXvspRJEle6NQ2IWm2caE6ibkTk0jb9ubUmGZDerHAtmlBWKjPKnPX3xGGxdT
aT+AcyMdz6PJuQcaml2sPpyM0M4FafICeXX2a+5cvf7coPV5sf8aJOBJxnm5FJpH
s5uJeB1h48MtGfiqsRQJyqSGmD1Mpwk1prck/0AgaQEMFct3zv9VIUa6yzdk3W8Y
923MKroVyreoJxRfKJabjAvtDXdfhBiYWk4n3gOM6FJ60NNgUaxhg1qDUD4qBuVL
kar9p18krmwmYYc+7GVfeSY87RWstg4iqH1Mizhs5y1ud+H7YpndOVaeRg434LJY
lF6Oq8Ip7H5Ort+Ewt9IRRf9AIqEo+51nOqwmoqXGtsuYrJ6NPu6X+AiwJc5fKq4
JRSlUdNVmEzjElh9UZL+PAgh79hckWdmRUW/BKErdiIjYrDWbrnkbd+ENICljyLK
BXpQ0MVWGDocuSijEuX670QjiMpJkRWhpUNuqM0qSCRt7WlisCgALXL45Q1rhRQ3
y8p15VhFf4rP7CHctST73Asjkx/7Vs2wAvWKjtBLJsEmfb7dkVwSAwKlK04ufoxL
aHdTb2MHAvOAVGkVCqLrtKCtLTnrxxlZ0Yb3O9ORWMBJGYfB8t8M6jt4pHUs1RG0
phYUu6qsK+g4+w1GVWfMo8xzMlx7ltKuIO+/b3zRX0m8s9ZbSjEhyAz06nFJ6Zb2
ef2kcpenmq5ZMGjdjZp92qjHQrD405ToWv+fprUUnfL55fljPQCWIfibVbLaBAgX
w7F5NPF1SpsgOpv5FzzuA9FsbzpasId2vinI28h+3WRgnxIHmPqPtt1doHPMnm6e
3441PAyj0LcqkMq0ObzqLW8bo23zEvK00c/BN3YC0Knm5LwpxKTowJF0sZlUR/kN
OawIa862tu7un3c3CMMeHr8TZBHDFIGMlGLAF0lTOj6r7G1O9EKQZ/lYui6eSTtJ
kNP2nX+uFK+Pb0+3BkSsH0uIUlmF2b6Nb+5nq2Pe5//aRaxp+Q18sdEXHCAX/YUP
wnPKCnpUb9JPdLoLLm4zho4x1VZ0LChJBhvZKp924UgYSxOoo2Ss2P1Qu6fr8ovM
j9oki/+aLwc61UYcYjQYqo7anmHUhu8OJdY85Z3f+ujeSEZZ7uXDiNhuSrOJ2Xr1
TH0PlJBG9lzep9venAh7ELmNWKNjACa8lOuMAtHShFFRBO8cZHDHOCjK4tIncc73
2fJz6i22AfZMRVXdyawY21TzdFBkH8hU7G0TNqSB7r86PIU6KwXHFc8U2K4jARoK
C4TwusrbmxFbCM7VQtmZCozyzULmCmnYUcB3NTNMsSNpwLb+UpvLkLyA5GwyzK8M
ZWzGPi2M5M+HZXOazDEMrn/NFdPUPfbRE6MSTCPtS3+xqzEZDU/lZ+hYAgos047g
kbcHhpp5YZxEQVibbumir1U24uZbAJtmNGL7xtaGdRJttwrAy2adtCsWzFEUIh5i
hyrxIqKIyHCtHMgqrHL1dyCV5qod0uDoyWrvvE7U106AuW4bD0/GyCPUEyj87QaU
si1VZ/G995C5M0DIMPapvLCmQSytbFW5U8I2/+UFr5Z1lmkgWPa2EVQGnqLt98jx
NnY4S29Yvwpbna4FAest4JTfgsZtmT1sHkMQl+RClQxR+Q8V5oR6yjjKPmMFEjIx
vNdIU8/Xda/Dz6RlVtzwQuyYHGJ55Q76J5Db81zixpPCWj9cuge0GSPYfFvkZsb3
NV0BcWgafcEE+rFaoNQKekiI7X74LsPS6NSgkMvJDDD0ReVES1rjitS1WklMYxM4
VRRsiCbHTirOeGXWf+LOWb7KxoaxP+fAcgfN16H3lWfKhlnydx2pbTzzL3y64Hrn
7+ZYd6t+VR/KxHrznEuMCC4qISIr8i1uIH7Mu1OC0+kW+r673wckB74pcMogAWyf
vZNXYDKFy+qoEXnJ7mt8efQ2m1MEFI9NKPGaMuouQLa0MzXdNV00npgd9BAytN7e
Eb2HdfIabOMhhHxp+k+Qe4K2y/nlalhIfZKQ491rLnSDFmXSBwYinokuz9n1sunI
P4hQeOR18gEW25Ck5rxTW23rrBlttVWjhqYKRNw3lgXmOGe/4CTEALnS/+Bshh9H
l3kCrTBpz2kCQtLeC4FA+g9VZZaMeDK/E1tFc9kM01k/zGOvGPKbZQY95XstGOLN
gfmdDU63M8lx9rGU87aTP/kpRbtuEbsSadLTY8V2dQOP2jcc9nH2x/8e7js1yB3A
X1IuE4gTIvUl6NjGefCUCo/UdvVylIvgaexWVYmdpPwvs9ObOIuuNUb1+aensken
umY0Jvv/AjuDSI3LiR1blVMzDksWm7N2p0EJVdUmCg6ujDDYHEmflcADUWi7gCpn
6Ect362SyA0Ylj1zhNICOJkqn+zLy5a1eR5sGtA1ELJYTqF7k67snsM5NjjDGb6c
XhZfnku4JTgpr2pwDxJ4Nn3X5bEagZZ/1Sbm8KVfhM7HhAy0ZM5EGGclwbMFBRQ3
gB+i3NePiEaGOpFWNMpH6UgLb7/5OLmXBYqyvgh4yao/9wtR7oQXHZBFSbGuuOxV
FbZ76fAbGIizlSQCSs1vXAVyhCUccYVPUNew/AkqlpWsN7BYRBNHm2uUzYH3Gnwb
C93Gi5MGldYzjQkYYIy6CVxsDCbcvDSslokX0IbBj+6L0sV8+KlHReQSDPghiM0G
MyPQsO2SNh1y+UzgNdokmM4fsgx7LJAmGfIxUUBSdvyf+ZAmUab7ki2mN5bFr5it
fb1EW5wtomguQDt+Ke98BXQV6RFuYCl1HfmqEwDQqe0nc2ZFgWY24k99y4ZfrJEr
6Fi8G/ho08AzX2jtMzlMNj/g4GxphBHh3EPtcs/EzUBcBECbkaObEW//3LQAb4Pc
3/Sm4oyYTqPKEMmyZ07L8gWPcWVLA6TtMFN0Ccj15nRbphqGAynuRq7PjMxDUK6W
90vt2IVQOdYtuUSO8jKhpHGhwXUvCQhspDoY4NxjqiTU/nnwh1YoWaTzumi2Lay6
6RxMyDJQ8Bl4/ilp8qXFAS16Ubo1onjcHuqFlpg3Ggr6jOb0pS70aRcO0isi4ACv
jBt1L2jhUv5whECiTlvVX3J9z1yFGaDqtROm9/KCbAHrGMgMLaEZ8BztjAcTmQ0d
mUWD2lrnPGWKklrc2ZTEkwm4n4mdek7GhgidvPkJXdPlS/GqcijkUEIiv10RCbdU
ViIRlufmM1DThuDLy6SNqB+S4uZZT2F4LDt7lR5p1qrAH2+AXzRkitgJwzmPXxsF
rIC9ELlc39gLi+tO/es7RK7JRWOsHxAS+QqC4w2qz+F4bFOAdosVUsspxLw9FsWL
4J5S1pdW056mc3O0ol032XIretjo30G0AZwuqMUPhT4SLb4XBbOPd6YC2BYldUWi
Kzd1h35OUuqXCEzhsGiXI5a63vWRKi1TshN8mIIRa1OzP9d2NFfIB7UYsqAqKXm6
SNLGfP1qZejdhdE5iedGw3ideAOg2mbrwg9QEdx4Oi87on7asHkoHYwb56qjVCro
Xl/fd/wxoyaFmX4JD3RVCK2ZMTEbdqfvlZiiXmOeR8TbJrsBBv2HBmnpN42gaPNd
2AGGArAtotJs8uLc2UwG0Hd+QerXThmsspOoZva3eJ6fgu9UJi7wL0oodc1xtL9M
yuO+pDOXx2ekHTVxNWkv2x3SCbmBTB06/qbsWa3QDJ5khZnWKeVJCUcjeCXK6TcN
D84HKumd9CaxldJzkTaJ1VcDoVfU7+/avmcSvuZDYuRzdl+tD4wsAcX988nVBAOX
Va14APh3CkOcJCdO4Tbpc/iG0RBU75ySAuS82WbLiZ1/doqdZjeKsm+Zf7jmVjiR
X1o5O6LvOItqQmv2kMuUIy7Bhufqj9eGiT19/X9pwbyzrA9t0lObzFYV7GDdU90l
/BV33dLcMQccyvQM8ebp253CTiSB6t8hew6Y8PrhJNgSAUd7Eixb+0YHAxyg/OW4
C8ZbSQtO6VRoy8q8KytgqpYthZqLH9F+7kHQIl6VP303PFNTStz5c9iSrpjjhssB
tnNMnsb0ys1Fu4tRiKSUVRGHWHiPTHyh7jUFE7DUL6L117ZqsK7rOwSMCQhk1zta
xTNjTFf5rGoYI5XO8RspIM3aJyWtzMxBcYeYGFNSqsycjLD+7CfNtHjXg9n8Hjpj
hVhC38osXczJiEEQtxLI3ySPMShJAcr4x6oTmb0nEy22OwPNTtPvPWXCdHBWmn/3
XvAvwN0JsmWboWpv5Y6Xf9zVQCu2eXkkZjrSXYrbSqgfzqLaDsYNa6ik8yhNYZ1C
c6QNO1o0944ajewvTDZuefATrm0c5To8trG6I+nQIgzkulol6cWv1XjnKb7hamce
X85xpVBU38CZrHuQfKrWLuTrqcLdib/I3/lIN6MC4LUYZN6uLqFGFedy+5kVnnOS
fx8oS7bwuvDBYFfCQyZYAglMun/eJRmLtNgSFXCAIH1bal1RYqD7iCuyDpTXKBpx
FdnliIEUXua2fLKsrd0nhLzY6YiJvVHXJHBYVdAkAb79bl2Uji6Yah56dXonmXYV
iu89SRJkOXFFuVKtaDr0M8JbMCvccUMyAdCrKselgImcuRVRLUfneBkMX42RTxQl
nPi/mAei1ToIzZF6EKLgvTMzDcgyyQkl3JJJg2bz0cyjY+ZF1KjxO5w0FFBle+jP
O02Dt4yol8APcy/p7AoM/dS9USD9UqkOC2iyFRwMycjqkk79Ok+3U4v7rJaUFAEp
X0P6ySmkgPTWJS88FAWM6eSnd6GgSoCf9p6v5DTi/+H4cM1mb5UJ4/rMjgrQrTye
Fyke8W4nR/YQYXT/2RUGP3Ep4/nONgOfvuTFRrq6atQ9UEtsEIqMKluQICPgnBDm
aQim4SIZEbV0Owo/VJFn7r9uSLAhHv5hH8YYmGWHhfoQ3SpnvURNEAMZZ0JwX3F1
HuC/AkbBAkD7kWfxiIIDZKG+WuQ3F/9F6qwoGZMCk4Jq2Tz1nOPW/QeJl0gPbEUj
LXyLIDpwo0pgYzeeOhlTAP0cG7jTHCa2PHQ1xWXjXpruCDpOEKDE0Oly8WAu+KYT
0QXI4wNc+VcuK8Drf9PuGkYXNTR7LIGO+g6tjhQ5RaXWP0OG+WT85xWDxvcEjSGH
/pbzSZCs78x0HzVpz+reHj24zn1h7j0hoYAbnMxuRTLGhRVLs0QdGInfDyerJWQA
eIbKz4bpnN0WhyJub5LF0ZO2nl5HYZrkfNMBLHamecK5356uL/NV7B/byn+7dBiN
NQ/Jzy5GJbpk9H3ZERkGclZlkuvfXckm5Mwu3F9pntEMbMNb/gMN9OPoYP/u78Xf
TevZ4kk9e00uWOr1EavPPmPcdgNklUVtIHjfxaKmghRwSTDQwq4h5o/E7uN8PRhH
FBrJPPBTusUqN39mGzGWTMPJaoqwVnmKS3WZ/T99R6Cr1zGnOnL6+pDDh7Sn2EcB
gipCfy0v+NySL30wOXbqP/BY5z/ZIaPXNibSVSgt5++5DyoMO/OcbB1NpzX3RYqs
VA1B3k4QfUsflV3OnvTYkoLsB4c44l3qxrR5QUJNOeHb/X6MajQ3vgzjxrbfMHow
47fLtDZVqeFQiCSiQw5/UCHpQqspbUs5Mevxp8XbzN+2LwX3Zj/kJxsYt2r11CfE
bKEKgADal+kA7RXP8hvqN7snWiyRc9c7kcHiBwUsrg8suWHA57W6nAK9BURBz+BH
7QnSohWZxLKiJQdh9uQ6kWaQs3Am+7L8iOd4yiRsPULXby3BJ5aPhv6ZbwRT/+tN
as1QTUkDylyYynD31nvzxNPk8OvWkNWIXen3oAR+DzY2PcZEZXDGojJlS94xIZnE
3Kw09h3+30QNfqM0uopO7cMJZG8M1dlWGqwOoocdoPbp0tSDVUYaHxeBYlPDZqPP
XvvGm5M491m3uq+9dtCZcOR+khs+JG6yCJ8XEdAqCxmxpYIkROOIxNy1w/YVQlUA
gl5kKewJKsLhWR0QmnFr1ElkfVPmucPUXl3V8NlAOHs8w3U0ZeXvr4h41lVemRus
+vAu5Pl9rRpvHejG0+RRElJ5nQ/N+YJh/qxJEX6f8U3nigOnRZVZUnEo9MP+IvGU
5kUOIRaq9NTvTzbQcQ2zwd5TF/QUeMMZrOEFdSpZdQ0AcJNacPguOcR4hb9JH8Wx
KpyhLC7nbKl4OuGhgOrPIi9gIYWOOw9+Pv6dg7XikSUOa/EvUf/rwgD7o1NcQr1u
gcBASH4Gaxd2bvts7vkb1II7bdLcMEdfH5iZ6kZPQHgL7WOR/S+A+ptXaFZzWRAG
QDJomn33vLi6WWXAo4cgdb4TdRaDPtuSm0nNQKu7P33WgkNpMhcxz97Q7LuXuTKE
t+gTTHdmGDJwFaQuEoNZ7lrlhZHXgB2MnBZk12R7/N3EBD8JgcwfGRo/8+N5HrM7
zUT7KEkdigG2RvC4XTathAROrwXcjhJaOHXBjsj1h62v/JbFepMAVU9G8sudtkC2
AeJ2v1ikchMgysJNztJIlcKOB+jHfqrwxyIWjhLQkFZkOo3t9jHiUbUfmbE5Vdo+
zxdbOUGQ1aqZVS5PQPZylA9DioI01iB4eul05FGqnpdQoxQIx97PYFFBztTZVELm
1jyL5f0zkEW9QCdrEmzoOazI3LBd9dYobV4EhR1Z29sXCJYRRwtv/tBm1MG6Iaqv
x2Deva4gPuKmAjbD7CimVFLGDawHZL72aAF5bqThotvT8rc2V/UpOmyaezvYbE5R
mf2TdbLxW7JikuF0/LndU58sn3resqMNsyMEYVQv/5aiA1gI2YkHMyHwqSb72z8S
ASva2B7oeLL/FPyTMZQk07e/FBVBu1cHaMWDRr7RCDXy5GqH9HC2Hjlv4KIRfFwz
nWu4BP2FOxjl82uPDmJ8SMSKsBOa4rHwmY2Dt+x2tLJlJIpmEAd2+TKtVddhsLHd
1bQRSK4DlNqfMpaCmAqWhUAym3pVSpWmpHL6NyGd+vuduznw+zsMzwXRdflHN+dm
7u6/aCe/fAEtWjB53iJpsHmVWcggHpjgT1FvgHmqhnvmalzs3YK0H7W0DBEr2b8b
SsaHEwmv5NRHbMTykv3x+7zldyeElk8w1hPZSEhOJJIDhN6Gfm3YeV12gDplG5L9
1+wkvdem841u0XFoBap9p9iyw9vvxyxarnFnc8p+Dp8FR8Upr+U/AciaIroMmPy4
Xd2FZtF6GD3jgI5Pr47DMyz10PB8quC+ztgls0b2mkMvor7ydSOmOit4Sfpf2es/
Iu6Oj5zSWjOTEmBhun4r1a+pM4gha1h2M9X350cYOdeur+mGYgs4TutcnEqoxNtb
+Yw4djF4ulWALvgGUV431qw8/xKZhiN8xRK0FBU/cNgw7EQKv4pr7DESy7ioTGmz
c9AkhBFOyVS19IsoHq/IW25RYRuTRnAUlak+teZbigMynvh9Gu/eNQZiplST2olj
PO3SiTOshPR3VOrm78E7EO7Rzpn+L1Z2KZjgbAXzq5ZRQ+NQ0/Laaptnlmp1uSWe
Sa86n+alRxpz18OWlkxW0zkBcOGxN4vfHCKDIoH9IJ0udL9wrI9glkAPIqw7Gd9N
mEyipeK8nCedbh/HZcyKkb9hLXt3WeRg+/VfPDYUM0tOrHVLqxwr0bVVF2tGNoaD
3IpKsRna20FkHD2g+/4TKudJ0ftAp5vIVyxHKPfvzmmrRuZlA574klhJUNUsohNH
UYLptqKR+NLixafAnbo1I7Zk0DnLmJv2yHsuo4ozmqZeHytJMgT5TcFK2PXIr1mv
L/DXHJgR0Zl14WxWrkF9ZqVJohATQgLC5wp0E9d1lW/VdKd7l6IpPM1tIcnFZiP1
syf92kFVNsMkqH4trbPecmEvEEkPQ0H2XnmYPEu25ygNVc1rQSuVlpRXEFUcydYI
uY+NcSMKY+Tvggu0vmIDflmDRC0BbZD1c78KDLMlfHD+10rp6RgfWv0NoWgDvxHb
kfpcmtBeGsDYZnOiVZE3UmisFFWlxNqDhR8FtLUbbbv0OD0rBrNqCNKnG1Z56ufQ
DeKaNhLgyyZHOAidX3Ixiyk35enOnMxLFc0+pldRY589WRr3HJd2l3FE42oBRNFv
K7AVtD4EK7XGBRxsxwOkN0XXSTBPQ1zhyG7h3Urq0faEkMO/DQWKuOKTWMUxf6Ta
BQVmvWrNBO6xVTxuReqfGo4rVoA3hZcnI2Qro0dsuu99T9SuSL/IMK5ImT8x9utq
LpM9G84aGHrCPl83gGXaLpryywkFC5gB0UxzI1mRPSl2Kj2F0IA2y8upyVNdCXTO
WfXcGgq2NNGwOMnokXN7w+BPHY7823oPwf3NsZzdrNKkGcvrrHjqQPdXcZEeiHpH
FXgHudEq5zq1LMLn9JPHZ9y6l04Rawpj9/qXwgLEWp7Zf+rVQ0wu4QqW+3hwayqP
qJI2YLr2lD9m8TSUiiQ1wc0DgxnDzpD4Q8Yohq96ULNyW0MX6pF8Rsf1Rmus5sGr
dEPikReCrrxYbNBG03GK/RFCdARuGHflG8eo/0ouXsdAI0707FcqRS2Kj9Fr0URk
BriCMEGINyVyBgT8oml5YITHvnRxHzHXt6+nvUjTodgrCDzTSpjqMQNtpR9Teva/
55+OyZCiyEdx+/t70TRc8yMnJrsg1if8Pv7QqcJOrOI8gqBdfagf71/mtW7juprt
GOciXj92bVhIv3ojMvUy5lqpNJbuh8o4n9a7U7O6JymQz4qHr6NeEeNAFKoTQnCj
hklegcXnhl5GND03TQCO5EJuqXLldIafExaLNc3Vljn/s+afDtFKNzNWEDV9uwdb
KqWUaZ36RCGX9HerSDWA7jv23ZLYyaH+yAOJTptLJVLKeV7+ODpo+Fa5TahxP8F0
X6I23LzseDNOhBgTk90iGral4E49n/f7Sggbwft2uou87EwbsIGOG46sCVoiAeIg
7x7Nky+OKS7rAJLAUtggpgGuTC0kEaeqAI4ek+t3oyYmpwTSwt2NXgPglge3Z5vV
7uW6R7/OVfLgE3yZAFoyV5sgbATMg6Exd2hh06hdzS8AojOSMHqnOXqPXN8MRXH8
efY5hFIVV4pYv6VIfOiUhVzRQGzrOJ3eUGpud72Lyjdu80LjGQhQEmwlJOqjPDHL
dxY6gKRw25e93k2hy2370/PEkzqviaUkxXuyfIYe99OIezWzFzq1MSyJYzEVAt8G
zXF7nHm1x9UOLSe0TIeQNJJ7EA3RA/C/6KccyFhwLsdNTjC+PFkge8BJKJ3RY1Vp
Y9frTYodLZ4wMsDJJBTJTFskhbZWT6Llm7NubvDQnlxLtASTnnWfBtLbABSE3mj5
E3CBDO0lHIeRjUho3K++z7FNMDEdSAJZ3zRf0wpNdmHB5CpuhaiOA0mAF2YOQDrN
bQMal1esHHb16VuSFG3vEw3CEFWZiH1xg5AvYllam8dk9C8MsD73LzuCZ3dGLUk2
M2W/IWYg7i9V4DVMnrymoce98V29a0gIdzfDnnLZhH6XZ1zMHCxjc/VF+MaYLKYY
pqV26BXRlc+91OcwKqm7tcTn9wtgSIsXBdEn56mYUUDWgkiXHTSiRtHuxkBLM1x7
uw0tKy2ZVW7SO0F4HbDUcwzMon5R/fsZ6z79tXjXal4g5jAfo1rz+vWIreueesSA
tUBkbEJIziJ6v6yI/SrOh/BQKXn5XKkcryuJShu+pH50qroZHESGosWLJCd3ZEa3
mHR4QLRT+XvTRmNqJM6X63X/Lzv3VFb5sUZWMTaYRNScviAS9hdcwdSnzPLKgBgP
tjxjzur5OviTMkWeD/fpGF2/ltM3ZXEmqURBwZw2mSnsvl9Kdn1r7lFURS4IlQoD
1PQBdhli2CRo1Y1JyG5gTsdMCd78DvKFDV5RjzKUSV5ank+NpHgXCk1MGlKHpF75
5Oa+aNnGX/ZjDOt6ODVBFpNPTdphh5iWz+cPxGwwibig56rfewtf9MBL7P9WLhAc
Gx/Bq7nI/Nwm8MwvOpoUj9mLCiYk/PENrwmHitXPh8YITROFliwR6PDwdts1RP8O
A5MIb3dEN9DL7aD3Or6KqUYr4JBJxT2pN5VcTw31pU1EqJ6ClnBVZInAmu1AR9Zz
u9d/acHfhSAe3bAhaC0nWFdLHhVFaHnx/vzwv6DXSGPBSZm1oAh6aBuktE9Mm89E
we86bMLhYqgRnsbBOfH9UjKdxquL+ZbCOJLyH8LH0pWbovv7ybkrIQ+DFUOi7iah
X+kDFsKIE9urjNBLcpwLYpVUjPay+yxbwhzFWrWDUpMwN+xWRgGserYguDc+6tFE
BgeQSJiv8qvMWQVoEwLojzfbKqsSiynmWWuNHKXN+FolgPu+xkrV6PoAd8gS0Jdk
0Ro1S53++bhbGdXlZtbMoVfLfFM9gSl835x47l6//y1eG/gOs5vkegxBvjtJ8ycU
afX/pd6sLlcfcmsbvsYjgAsvDTei+8X55iXCq8c0l6PIlrJf1Dbq7Ms7MV0zflMc
Sn3lDCwQAepRKF0uQc/PLFWa9B5JBgEwPSWWIXkXcC4ds0gWgOeL8vPasLzcMbjj
spMcK+EbdpRTBYmw9h+bS/0u7ezosSFx8/JdJtkY4SPSGCDg3FJ9WS8xI2tIwS9/
B639faqvHFqPxbjlMBP6QM2erAzKklW0IPO7S4RbGcfDQ3tJsT7EbXOwv4QEaxic
xdOTgFnSMXn+E/1AvflsGMdnpluAAJgfunN8hbm4gkNrJzuGpZv9Cr1lpmvW5ddm
a0y4OgabO8+ZdCPLikAjMhInsK06A4fKdI1DO9M0DbH2Jk1Ys6VzZ44K4R7fs5T7
e0bj1RptClWpmv4Isvo0KY970l0QpU/USdwzpeaRWDU6Yao+Y/3nLSVoCxdnT39H
9zjr7NyNQhwCiGFleeDBFYkhc/g0G1nx9SjbMMJ+FMmHUwe/9TrL8Dh6UZQp/BwS
fYi8ZPygj9ToCDFOkt+9ZIwndRMS+/Vcg1dT4HlXLEQ+LspHY0wxgzuFIlGqGo1i
Vz7tOp03klDxWWXE7clxwJP0ELra8ksYm4gLXLSMzIk+6+umsex/79CH0eIp9X8W
s55pKuYzrp55pxsnFamwBSBeJwaK/GGS4qohFTc04NhsXw92FLoadXuonYh4X++x
ZMombdBpP/2T+nj9XI6Hyr7SZ+y2KFEEQ1bFCh2cKbEUKFJ5rqz49jgpYNoiSrln
Xw0LTbDikX/gLVKUOgPW9Fz8o71a/TNZrOT8varBZ4VzfySl2xG/Y3Ue3x+/KhZS
ipQAqzBAFxDrqdA8rtgZGY4qrNyP0rbSnPh8bPxJ1q8O2FNSBnrLMqIN+0cZyGTl
kW25udnACVTFhbtk0br17YeMtpNo7M9c6rD3m2LUAoKZjsWQs7rU0p3kLrtVlwEN
6plVqkgJcPQv3X06vSNpwsP4pZVWPAgAXaJETnRLblV3jogeE68kn4L9SPDZncRP
wrg9BjzGNFJ/k0e1g68CQpGR30SFau/3mz6Ktv3RFuTMdQrbZtD9kKVer+cWDyYk
lCchfSlbypGr+pqmpGxUaWWOBjk6Gn/4RMroFSPlSoSRDp2Oo7tbQZLGz8e/eAza
iQ6cv4MdyRASRmorERroAEvdOCjnLs43XA2LcITBSL26/w09OcxcMfYJxawHsCZ8
VZnY8exuxZy6VMODEuzdHnM2je0YxlPYZf/rchiOgYTxUBL8OPo4JuVfVKheCnmR
jCs/2Lpqwc1zbfHW2FtG39fw4jKbY2t7mInNJ+g8zT5Ojk8cLJj/yTkOBErF6RTs
S6xhs3ocJYK/Ri/XuuszID0ZSgbBZpd+H1p3G7+Ve5BdtTpDK3ZfwByoFEHcUNxo
gO+ywAi5fw9Z7KZ6zVSSrn+kBNdjdX581TJHkQE8Kxz9093kdJwN7jUKfSDFQ0ED
hjLxN7Vr/xoSmih4ouJPM5bEsXW91dfsVuoYRNEiaWgRhS3fdIJU0yCJoQ68keD/
+afEnoeaeTGLdAvuWHg57q2T0q6tQg8HCuFhUw0lrmmgmqHWaN219bBIdwA22i4v
0qRzMXy0/8HV8I2z6Uo7GjUQqyAv4udi+VuWzMkY/MkAC8WPO8XURXi2BD5GG5fY
n5wrUfzazidw3y37XjJfk8Y9Gqr6ZbxuuyO/3p83W16K6yQYXfETZQ5perKBqQpO
e9zWRZ65DlZ01V0cY15awphYtf8klPBXR9FWgOOeLvkIsaABGtWkWrvENCCkF+xK
u5rz7bNGMtLvCqNkN4yNO/wY/YpwKq21H5v3poglQJ3DLnfDve3tFSEyiFW12V9u
jsCZXVPPFphzXnSmgM4ibM6HYAKAqnVabsc3aqRdI5EAtcE/o1esK+Uw3yQKUVar
NroPTZUtqjrn+oxfpnCRKVMDIumH/u3XrsZZvtki3MeLtgo8ZVP+rgh7me3CY0Wr
NO8/9ZsJc6Wn2v4XU8ZyA5sxXdh/olueIZkTlKX/zmbNUBoLqPTWPFF2AxeYYI7R
isjm7GC0cv5lBW3JKyeYvqF5pSV4FIIbJmh1GSUZN72Ydinksazzrxef/cOz2A5M
UyLERS5sFzspL+7GyuCBqCn7sKsFDXPDW+FaRoeNGnqZkSzLyKve4p4TnOmE9WAl
OUw5V0i2XhdBEhaVS8v0GDxCvrSvJysQKDzpRmoHCbgSVqm771c50R3I1iXCzCJE
kYUyCssxddEzIUuIl3G0WWdmrR2elKQF6nL+4Ae0fFJVt5K0T5bfiSFDD4jaJfmN
sscuu2NizsSrzxoymdz3uehB7aEctbdSszY2I2qwNYV7k69n7+sllXVOndVdVidr
tRX4Zazr2H8xmEvPLqCq1byB07YWmkG+ZM3MH30YqX6TX1a+pbi+rduGe6FLrGnU
Fsgqe4QwFOyjvJjNYOkty9C2Iph3OssEI4P0dmLkJDg1Bk4ZZ/BLMKaly7KdKk0i
TlGaH0PY823CiNiSXyPfU8xN6dctUPcKrVeHBlBUlIk2Tj/TTzw1kXsmvrKFyizO
5KXFY8UHCEBBvji1TBgkghqVVCKVl95/DUSFe8jfg834nvN7GMfTPpyjNdgNpi4w
0VkwGAL8K9hPdOKUmHBvR+5xysygV8WxqZOaztiNVCmDCdFPXSGLeHwDDsEKiq9H
oQ7V7tEoyAiM4C5fosJ6nVM8uf8LCQEupPovFnm8OryPpWSLpfKzejlZFf8pqB5w
3/5SvnrzXEYUBkvZNc0h9T5HKvC1As+SYrXW6W5cW/Wb5UPwQy0lMThuurdYPqWW
bwx3XhrjWEX0umF95XBaSKVOGmZsiKoehnGNC9+qj/Ed1FtxlPxyYdLKvHYwfUQp
Lmcrajp/mLjt6voifs67WFRUumuY9Kwyt7F9SiRaBaWLYrVSg2C9qLnXMD53Rhuf
sS4rqYI0c2sK2j6HUlevZ2bnI6J5Ptx+3Rux/BrrEUmlZoVMeQSqdViyJOW0jpUe
s6d5E6kTd4nxiFV3m0EXrX6eL9NnZSQppPCqiqnD0dCaedjfwkB3on7EE2/tROQr
WeSvlWxCJEtpzlciLhPAvxREn3sO4KF9Ta22UVEtz97isvh66el7FfFS9H5+bzGK
b4AtsO6mUnTOJzB3P0H8BUi3fq/qKSBLtkSmewjURWM+qC5EJx+snqppZUU+gg5w
lHY0VsOBFGqzquVwr/BozU0qe/G8X+2konpuhtACivTAmJPbQUx3RXBuHbA4tUtq
D4NEpnu/jDpU704vMj6d0MjTc4kmdwum5GZH8PNVtKxfdYDWOeYcSvJNZrnDidb6
5xigvHj4SJoF6xH48d1D7477HtT8a3XiJJsEd0Q0+2sukwdC+S88T2c4ki7X53vC
aIuHYaBYIlrt5uRR6CDhvcg2/hH7bKIUhkJgi6nFUEPXnvzmxN0hzXXnqthhkcG0
mlGUK5SKkQJj/JFZlcwlJISCJxCdLe+5pViXzYKj1YErfETkzLmosGVTdqA2501P
EbaPYMa56KgdkXqiju5B6HgpxyLzYd3uR5GSNEQjpI0JG5CTIrTUgdgI8LHplD1Y
LgeeOrC+5XlMxd//r0QULn42zE9REx5kGQ3/MLzeZdu44vAoeIaw+RIJfHN7QHHU
oJ6fbdsxYtu7u6AMe7WPfEOR270rWldjZ+y/quvXN6ZzVAJS4lYLzuzENk7RfvVf
eSmrm2ECW8OY+4n34cd6Ph+BBpLLigAAY2CUaY2LbAwGMNH8m09msLF7QlNdZ94y
fX96sWW2hODgcs/IyQWecvkzheGiG29eyNwm6esZnEy5C5RG1uDqmM7DharUC+l6
d/aYppy3Qauai2gX4+o3n9XznBxWdLZp3uyzs4GcbC0MTGR6W9bG9yFQB+QMs+LW
/qXc+OREYd3E3v49GICk39yaGZvFVRDCGNtxVxyvIiOsIn08KS6N9THvNSpnnnTb
IB4zRgKEZOuFgyox3BwUrXlOPz7O3+ksOk0KwGCM7MtPUGMCCruaAlsJH3H7Pfjf
s+wzUS14BJ3byQeWz8IGJYOZuYg9cAmfIRA/eGM576eaiL0mHKj1/yt6v6E3LUQf
19CR/kFN+Nk8sx0hpN67U+z2ptVxaA0D8ExLDozlw/NasybVDbVpcLR8aCrkgHoE
tbQyiILMcSiUSPLPRQGtpUXLvyZymLQrv/4XEWSbVKaihpO3zIQAbNDcYz6nUmeJ
7AlgJVSMV8CWPJdSV6Lcm/Zwf7co15pzDkMxDTrQ2SYRDYduzFnbSd2ne2Kq1JgB
fIspgW1VfCC/KueULmZ3r3eDoxP/UPn9oSqDt8dB2COo4HjMZiAw49c0iFAkFl0t
xgP4OfMEiTIan2kTMW1t1pWqDp70tRBmG3A8AFCaYbNmxxR5OEQWit8FyPRgkGRj
Fgm5CJU32O28vEVrGifpnr0GGwik855D3dmInVB7DJfmLaUlQRkqa63p2Pwj4q5j
eNjw+mDUqcJ5dj0shnN+N+MCt3MsHqdb7ZSEpd1VqWdqVLhilvrXRjRnaSV3h7Jj
0mtVIjZzpWpxN6g3CUFzt2B71uleV1zgWw+A5VBeSF9ErXZomDjYdjOc3BHYTzsK
pScjnrUefdVMaepcJU/Ww4mC15kSpzVgMiFFah+FCnhMCbW6HGlWnBfdRGQkmggy
xudqRYgdKTQUIu8xv4QBDcmsldhf5yDNW+kldANJvECJyqXU7qI+D+12GgxK5EqP
oio0ypnZ4eAw+6e/HMQWhuMnhYy+J/BgZCxR/lRhW1MGg95P8UdqasgS0NGZqUJk
Jtv148oxbqUmOyt+KPWT8wyTFArj81LP+ejkF0OJMfDeONyAiSqeo980F0Xn9CkQ
NqHZPdUrx1E4CTUdXESegsb040LYCQYppa33SIfsw86Sx3KpnR+cBZcMn/wI1zLW
LnpEIUKTgeW+O1uXzsTmctvaV+pRkh/sevSalYBHDztaPi3TX3uj/1snOWwqRSt3
8kw1x/tp3oDzWIo5o2FcjLZ3N0vGaOmRR4CfVM4MYDTZGTENL8Re/8znzdorr7ii
SV3JL3pPsfsxKP1xuoT8J/w09w0HhOlIdvfFN0E65jv4B9kGi3ugKRRJRnCINTt3
olBAm7mEIPG6gwZ3MoxCZzOu7iJYPk11Z+4vDiVWeov1KDP86a1sihK+ErnPUQjS
gehKFP+sSfFNwEgOX8EL2g+SCWgA8M2PV8sIC8f+Ai/SP4AQ1BBfCsDJkzdtJr3V
GWha+YJvYc/o0Rm6uYiYkp85cs0MLBXc9WSOnaaADLRBGQs+2qy8afNAewrus2ej
PWSGPV88y/jDOwPMT4rjXkm1RIM9hCcEnqj/spjWe1YtG03fn2Dofs4VRv7i1+if
80W9lE4FNT8rx7+9T5s8SpwoR2gBc9zUZA7PxUY/NaHJptTm28Q4AVwf3M2v7PHE
6sT6reDTXvfJaSlKgvAudecqW+rpoXqOPNZidtFDPQxiKtpnBl+7RAjXboXARKr+
Cr86EiT7RqpxkvujW9hHK223RgCX3A824r8tmmfzUU9g5NOswtdT81H5MfdJ3aW4
CbCsRkXxmxNwNb1SFxfYa4yCkvaAFIiLMgX2wg8myauhrH+ayFlGOgnwbHzFyfUe
RtIOqYKMvqiLTA9Zb7hcHVP3fuPR8Kbfp3dr9uxcHFRcMADm33VVmfp0I899c+dQ
fWwfqb2AivQ4MYN6woVmHwzCW2H+0kdIh7tGL6qJyHLgSU0yS6K8YH6CYRHx84p4
O+6MOS395QmOITtECtvPFbvA8WGG4FHgWzO69pu6leBCHsBwXA7JtRuLnWNB59qP
NEDhJQ+l3cQF60Np7IaCuJWpAQJ4Anl+04D/NCfIlc9X+aYwL/aPfelDv3ymp+5x
4FkWJZHlzLjSkhR/Dl2D/fXAjY+djCiGQhDWZu8J9Vh1C6/mmkfp4/isvNpqg1Xs
l41t+OWaHHre8BNSL23zi9R9/D4tp5GMfC3wLuBI6pU2BA7SlnA67gwOJSZw58qG
hP+5ukq5Iz+ZAR2EZZucHWM7nvJmG0Bmmwp2AXI5IHa7INh7Wbw7+vHZqEbmc2eZ
2YWHMPFlMTS4VYNTtOSl4lr1AIg0sjd4qtRjyjz7NCf3Kg08XzTaKIyh9hpA7kD5
pxrNhRf8x2ncAazT8KRIzqdQ+tKiSPfHeABCf7Pkp4fF/fhohn7cr8lSjoQjeYPf
/42Ylzyua3Zb8L3PCfW6Ab0np6yxLqutdccwsCPwPq4WqSDvfWKWUBNgdTkzKRNg
Wt6Ix46wW7TZ2ZcN35lpBoIqDIhu8T5gsBzYDbb7pQOAKhrXAwWJLQvJHsVLnq43
gG6i62DHxSg5mG2UGoJ9IU0IH6gUXpFfFIQ3/hZAD3rmBqGUHwBZOp4Lv3mVcczA
GQX7tKjikmrhfDLqlR7lI9qr2ZGA86xtYNNtDYYGQQgGXTJ4ldXqRpIgeybopdS3
hXq2slIou+I1H6zn2v6I8Fzo1Sw8/tiRcjHBkprWojL7gK0iCrcjj+e/AtVUMRpU
srDGko9CHVjjg/3Ie5fngGkD1MuT+LG43ND3AhdrizU8KniLul2PCeJfbuFE3by5
VzemgF70vlmUQ/RoH7rh4nR0u0yzuAsfx3GDqsI0IrM6rZLjwJwBQP1a5FZ9ksvL
mFfNkLZ1waORa1x+jotq1gTaR5g39v4gvTgEt1lIwWPK+q8yGIiMDlT4jd6zao7R
aqj0QcxGhpJrIXcfgpCNw8SpUrVth6qbzq/L0E32zoi1c9MVgjqxAwMjhQfw9lSs
zjurO6N+i+pYKEaOjqK1HHQ2RlpKWuI4lqzzarAlNdRby6g6RJR5mbWxMosVbG3N
rfejlZ2sgJjfAlB1Rr2b3CZHGChCbLtqCmol++vyAPk8p1z/cEs5ObsX331XJWFo
/dYbHQ3dvoRgJHWgz8Dw7hnuEIvGJcuHsjEH8+8vikFNukha2FoDpVhzfO4Cj6YF
ffkrYz6JJvI0yUFNySbO7byWzTzmj6f/szE5Qa6GSrrHg4WFDC9IpyseXzVYicbW
MwjF5q69aBVasIbDt/GNxcC9oEZ9flZF9b4ahFa3/fA3yTohFrtc4v6PfSwyZxGj
8gKA/2E3xsoiQn8ChWFzHAuU6RmGmkQLhqtLh3jJYGTK/emTeWgC1x+NAU0jh/Mb
gkzwXVKNBM2lz2PddzP99GqvX+4gQdanHOjT4Kw09tVe9rD/NZKC4juFjM2Y/Cvz
lhW0Ic42dqNpGPpu/z5pAmL1dxsUxTINKYOx+p/H0kcfh8IfhdN+DcTMCeC4lZy4
NyRuU61916SseQLfESHRxCWZRSaeo1ZZ3Qhca6wDgeQYo6JXkX0FhrdlFgobQM5B
YaNdPmmPTULDBmvhQiR1qCTfqlwOIJWE0YmjBbQj6p38gUT5DHINzg4Xp0yo+//1
govaxGV8r4sVXulw77e9l1CbzL1A3N4d+hfkP6oW5Z2bDq9uVG7jbQJUHNPrOevZ
TOu7BIFUecgIMA27vRJDpm4B9bNT3VM3nRfesfgdnfpQbTinZG3rkSZbw1BJWpTC
Bn+NsT3ipUsrcBqWsgSD6XXlrYHZnFLpXMHbRawhPANV5rhR3vsg5CJw/IYvh5gF
sCNETNDS6bStDetG58dgY30zXYT1P4HxMxyXbrkbgWc6Ux0QQntWAmUf7NktDMq5
iL1QWCBd8IOZ00PY4hJL6WJ/d5MjwBfqBT8Ao49aXUv1Ipd7Wu8OZMo3Yd8HQ9jD
pLKZ0INej/VclA8gdfh07I6g7VLpMFYndxesI0FhBoYG8Y51lPwW+Jh3EvzobmWG
vFdcHkBcN3Q+Bh5VxbQqqW0nvdfa2+faj0wB2BKAT9xhPh/fbN32i6mgnqNdZb6v
Qn49EShmegij+CyKzdUfRz6mtCoXv/jmZe/ib2muKBacGzbLyXAQolZwlvjmF4Gn
DiMChUIf+oikR6DDziodvvbsQIAN4IUl0hxWcEpu36oBntpD5z9+PALmH7Gb9Hf7
9X069QVPfeM5Rn67pAcTBrHDirhRnW6TbGhYkWlr9wxsm20RieXHnvjOCU2X4gwE
OxztidqjgeU/oq6jvmbZqhoyceKDwXsnqGf417S7uh60BjrEjFV+6a7egasn7cq+
1a8CF77Y+5DTnS5PCur88hocBwky1z92871/cRRx1bUydnXe3AgknLDiYXB5OmqB
o2SGBdvYgDyaNHgKQQp2jxCRZHu31bXOX9Hne43sqx4IH8DKvX47rwByE1HwPch5
UVnsnRwyZ0nxPjOl9D6Y2pwbOzGMKXEKvxSupOnBflwgHktDQ4qiKemELvFIllga
RixFwJo92bCxg466OkcOWL/BCCb5ElILlAiO9OD6gXCI5MFSXxUW87JGKr+KPAg1
b++6LQaKhMh4TTmkuC/O+03RCTQ7Oe/P69BSbm6OcEdZPMMZYA9jkUrhuJTGTG09
mTO+n3THiatjfxf6pkvsZBceAZYX4wNR69XlTOk1FcgRZPHcfz2IXO8zhphjEPii
SXy9ytR095oy981LQsOP2mKHchClejogV0QR7BiY6xA0hWXL1UKf3D7fpR+cVz2C
WJJoY1vHvAEJikHDEkwWSstjlqsFcrKBsZdJG1OCy2SIFLUZJ1K25OEpwip5e86r
fTPvz0GORG3F8ds/6AA++leSaeZPWqu3fn1cpkjSEudDJkeV2rfCYCPHDkkhdiGh
Ve0fEvntBpQqFgM4nbOqFaqaD7sY8FL6zW2ooZqyV/KioaZMNyETu2NhlQJaolHR
TPT5YpBcRcCiwSci3sfxl9ibjnelLWfhxNcbId3vlMfn3gPrgPUlWJK2QOX96X11
nHUSZNnatrxCgiRGqW5sh/mmZcREQ24IEsHZe4z0zk6YexXPwUVCud61ACz8HbkG
NvivC4Zp0uTDXUry5atx/Om73mjjf2MuvpwaHlijC4hvEqYuOJnoNHk+oPCKveKi
MQCKJ/k7vYbQ8b44T96IHYB+4SKfFZ/xFd0aAmYRZ9YjL2ZH0nD+DcAzGrRXBJOQ
b5zSDT0hiAe7vDJGYXwVTqe7qMM6FmZAf2KbG+k0+era+Vdxo22JLSTIae0D6Xox
Opyh0JUJxoJsLTCEbauWPf7puCkPtd/8evaLE6nD/DvRbeCRrPEADqhwuD344rQr
HXKjqqFY5VbAzBOJ2eKL4DdEq9V2Qadlkdd9ob6RSQdIODlA7l92Hy8hBJAxJxdA
SU5umN3iCNO9OBxd9GGPrNXiSImXEP1U82EZtZ2ZO7qIjhDofFLoIrdg9oN2rXYG
xwDH+vzU/+23zU6mgvBKVhaggOJ7k/h3aA77J+wFjriIRhe6Q1t52AlUfVumrX3/
7fIQD9fdLd5LYJ7pCNNKdjIceQ3pzv91hrd9gkkM+JuYDL9Rq3kMP+IcOVlSiB1z
7EpFQODBt5smUlBuRE/W/oBpi0RC3+cuGoybrwHlVXgQbi1gd6O2yfmAiW9Rgu+5
w8EZjtM12fY/oXS/9Y6Ysqt9oYW7bjaLE0m0EispHFR8dVwBJo5slS+NG8aXSKJC
qlIUH9EeP6m21FqJjdrTgRMEjwy5XHvJzzgDn+AILyhSdPz6A/STSElNhtl54bl4
hNM4dAsEYM+a8CDY8zGvFIZljeBm9HyJMA4rWxqLSc5uyn/hhJaslZhou9NQJNT+
c9vrb8C5c8fzSHSEUpCqqvYMB8efUaHuO1hEl7IH88WpSC7REmp8Ze50XO6L1WJY
jJ0uo0gj/cJTgbhrBNGM+NDgNI88r++dpE7t2/6zGMy/uDKTh5yTaOO4me9jWd1p
z2KvHHLlUXCZjYs7kO7+uwLlBYpio14ATRpYILlRhT4g/QSJvZChaxVwnz2yDRoj
D1E4OjVquLOc1vnAC1xfQPB0L8CNFrU92mza8zN/4+actrKnEW7345shSPJblRro
Rtwn1F/kjnYyZo5qntRzFobQphTkDl7fg31YlT6QEKf9wmjWc7M/GalaIQoIvG5f
dZ7WmtZolqLWAhjoYCXmyaAdyw0mKF8H9sAju39ijgOhm4p1N7m5tpvHQzGWQ0Uo
VMKpD5deJjH7tdgBMJSWdUXpVFF+vqbMyrYJFp0dMwIrZ2gsHOKgbVhkqyc7/Yek
C+eHu9KS62qOw7Zb6MmPbfBz8SyaDTbh6Q6cAO/7QReCSJQy/i13/uPwmEXLckZZ
Azp3UM4jBp2v9tbn1VTUBfRKj6ts4hwb+YYITL1M4vWeEHajmY1nfEdDBMszgJMI
3IdSjrSPjxaLbYLSabh7h4zT+ZEVLjB2lGvdsOxcjdhaFE7bNa9ydujbrSBgDPx3
+QUflRXBb8C7aMD3Huy8UVqFIQm0SKpBJk2N86EXcGwEdz4ApbGxi3FTEYQq/j75
dVSgdjWWaEG5ZdXON8fp+bEyQ5w5dq9drsFJsD4gYCu6mhy4FluPZ/els7BcfdgT
iraXZsc1ikAV0YCQhmd/GZiQuFrnrzUuG+awjaWGohRyjAPcpL0PUXM2kqt9SRXp
SKvxYv0fz3AcoOgJ2h4GKcph4ORXH55tdbFm5/4wxIpBC5GkAyWdumPlN4BGllSl
5smpwmSBng6coQI9rQZzSDKCIdSVoDiplcR9MohNUAuwLjDrBzcc26E267VX3ldZ
MZ5wof7O/Kbsr4gbpb0Qe14idrVZyAzjNv9np7jVqwdRZOjm0upM59rHWc/ykIKT
kWPPVSIAZ+ICxSTWeFhLqIhm3dpyuRx9d68S950O2o+nVq2Y9PPaiC8SHOFNO5dz
Z4UND5yPGLHH+hqjdRtGyUhJUcP1GSzqmeMZyPsDHxEREFcYoPTQSJ3ljeQUpX5j
8ozVj11T8TO9Fp9j3Ws9XXcnIB4wkzjNza+2+ks0TvbvxHGkZJ9xdZEAc0yLyao3
EiW+jphFbRd1r5IQ/a0XDC9YRsUvUro5xMxE4rOgHk/pVsXkYV8JGb18HgchEFhN
eNFDp39iJsaW7SSVdYqvusi+f5FZv2uVUFz7zCTpgpzRa8XTNfEVhAFvt0lKHlRD
KZsNcAQVcvf34pYwulf/TQD+53h1aR3E0xRhTV1ZIyGP/xcGMkqyWGgXDi6UWpJx
AHyXdANI74pKBE1lwDS26wxuqYnJMnohtKgmEoDZ5Sm6zdhH2wobhclrrN+6Qn2R
N6/Fco+lY6+c5NwPWTD/Qhgnra07a8u5OMgCkw5ZneJaUPg8m5BphGzvolTTPA7r
LAwpzH0TrCwQfFC4nTOYhVvn7zFSiXvn90k9a1sb90ctYQqztDRQ3abriIojGwkP
1h67Z10hiX+DwWAOlt7rwpDcOfhnz78/+a/Xmw9BGp25nAKvZjc63WJdMrarPHg5
SqvD0wTYOcTp31Jq4DLTE0+YR93WiGMsw6GSxY7s5nFCjFicoER7MbuiIbqZHmGF
WSMaqYpI3xtGAh3aWoOaP4AdtgO54QG+4wjhYqX6NTXaIMvQgnfoeR1qCMgNRZmS
IR40U3tktMGHuXo005YpELlbNxy3oSoufrUANyU922qfSMnJiqQV0aCASWsFKDbz
jQEnPWBp7ZpE3fse+vHcmQ74TvkLShXWBBSKjVxVZZE/K5EmniGzfWh3OoHVAoY3
bKW5c0B9ACL+3YQCaWfnbVbJrPJJqhVEM9Ay0ugzmDUZhcAcNd5kcW/MG1j6efMs
6qK5xYHzFFPTCk1AwA1q8o9vRuhe6fSIPATmQ4FvEuRfeC1vk3JaeLdQEzcfKuTL
aHjdFR/N4ft6fcuUMILrHTD+9Zuh6mf7CuI0Z8Xm5R9xL4NSjBkaCLXCPvR/qas5
pbxH2YKNCwhB1FOff0Qn2jeMqHsgN8puz1qq1PQWTObkuA1nSwTfgoZAfgruxq6D
k/T+aXUAoiqx9Lz/mi6cNhj94zvOC4elR40cTRkTPtcKqP7f5btlkuoGB2BOnuux
TdpCEsIa6Mawm431anLj9o25gZKOMC0eP5iGneR5p/EPypSqm8bACSE6aNtGjkgi
zDSynb3U2/WEcOYrpSGfxKa169e0cK4eV973IOMiod2SNvMwTOU1QScUxc+oHd3j
O4IJPhki65lj9iodjLpAEYTB+u9aXb1PNcOLOh7P1ww4smOi7lRNOHfUw9uCX0Lo
xI9to2G5yxc+gAiO6DWhJ9swNtcbxbhhNR+Axxuh09psa+jkQGtBIHBNDzy9buRj
YGAWMmMMC6jKSJVajOJ2sTNd1FNlXzRalngRQEAXDaOWxm5xUSClFWangMoMOWcD
ML6VBKI33ePTR6QQNqIQEPOKeh1zcwmxqabXvbkdLpI+ppMG8RtCMaIGq/kOsIb4
CKWkYVW+1wQg93pA9hTfX1fuGDtNzHvnp7R+K/Ye2RkbwZVi2hJN/YKm86PjPadM
GvW0eQGRuifaK1wdEA/6JRw9uW3MOV92m6EzcJI4307Ly3mO6GejyrKGZ60+sQ8Y
rwwNfBNFwEXWN6iqudkZalkvjZTD3QAWfjJcQjUB6iNabc5AItPYKbmJuDlRI0YS
vAky0cVEVW6IBnX2iUrOvyO2A11jskJV8WhnYHxwwlaocEMzbhpoyjXnnj0sxHIb
VPEfSyUnLcXhJQrXALhyYvoL4z5AqSx0ZxXSNvXJKwz8nkC8g6JQ+ZM0UCy+BRe6
sPLyi3zXWHsnuBPf/i5blsPHt/O3JeWjrT4iivmiFP8yMIxXE5+54j3USOURT1xg
4gMnR6k+A6PkwSt9Gw0YBYqVHY6An9Xjni6dtjhCZoutIkyaQOTge1zKafjq8tXd
Hdkh6qZZf8WipjdcrT7hnpTLWDNVzyvcfqgSYFeQ5f3msJajXIYNhoH2kZAZPvD9
ZBYDk+qmFgsSTASaj97/uW4GdB/MXfzs4PDoHRPqIlosVhASDhVgymXCWpYDcF75
5u/roiIitTu9NORpgGNiajerfhOnpdX+hRtbzrMENZi5SWzvWTJtP5gpcJhpd6NY
ed/YLtOyt23qFa/x6Z2xZoal9s2x5u0yxQckMgEZGcCF7YWtN8YL4sOJhWg7Y16f
jS2MXvRQbvRo0v6/vG7d3jocGWxcE8tdzqpohqUIN4v2OAdntywSbBubllZxSDxg
VyzV6e3x++RBD/y8OLnD6XPTNr0+o7tnykAudqjmCKcgxfHi3bhW3EA0Sr+OYW2n
39pY/+LV+7ywxzVMcSgNZq/ISBzNqEbapCeGw3xYYDmhxOkKjPkzEg3alo/AdIYq
n4vWEnuZx3RWrVG4a3hFmS+PImywI8CVS9S9HCwoB36BEeyr2Tjo86UqG8QMv04L
1oeGJJ8nlZS3bcdD4+uvO8HPaYapZjxY+2luLYX/0yDMqKHTn84OCn7bl4XxvN1H
QSX3g2QzFqTJ4TAbQ+RA+Rwrjpr10nOU3C+U43Ln5Y4Fn/KQ2O/NExasfuXKjhGk
UOSRa2995/SQWZH04b2aRpwTP7DW2KjBwfz82BclImY837gpFHN4gxhgy2yVjI6I
JQb5Dvp1xdX7jZ20PvCb3E0jTkULY11iaLqxH8Rkeh7EmgtApMe7onNr512uZeZq
sBlQVTpC+nqA8aGbIGLLbjC8lV03tGh9/YoRPgFOTRRBreWvZAQcSAnF4i+fwuxh
pxoKulSWgJB06VoT9lJUyk8XUZul3GCT+JTJX2F8VYoyyaCKcspN4LDektcqXoUn
OjM7X77O38tDXuivqWQEYR/QqRwOa8i3Q10b5ZKKn77oxkucYqPzyuxyAXKnO3ee
nHxQSxY/O6Y/c+7v7hgamjLRgAAhOY/NgObv7kB/5GhxpIPWKDIy2clXLvrgGnYy
Py6MOGnR8Vz4RirfzKwtVoOg6IeqseizmphVB8w5Jk19MYVGpZcc0OYGBwmdJEgq
C99ZlUNGz+C5dg37agfFdSx/w3xefCNsga5IdBnkwFapfDOYgn/nH+hs2Q1ueuow
iS62sZzmODvUl5xSA/uV3zIgr3n0apCbehxz0YTI5qF+HNxyLs1pnRmGcep7PxUz
CiEBlx/nOCA5xTrPWANVVEi1+EP4lkl9QfS2vSVTr5rCiln/w2amT90qpEZ6p+wY
FF1hBMGwjLVyyfDtuMByPzvlH/meSnZNFI0QcIE6LTsyyUWRRU5LDg7Iviprdm7Z
ARWP6/znIb3D5e/tIEgiDAx74qFGxxG3xBjXSaCUw4sG3bnOZjvqvvCqqC1pVFw5
ECXJWp5DWII94CCPbssMZ4+HtxUVP2QC8colNi2kvosV2pGlbWvjYNJw965aaZ0z
rxKyGz7XLn8DDl+sFWxqm7cOA+1ht8I3Xaf1d/uOkfKu/pQ4SH9A8ZEyRH18bJn0
+7RgP0XDr4f/QxR5S0qNRZvr7CAQfoYnR0ODxszITerR+pdJlSFT+ZJP/nqfn0ia
Y5o8NwpGwkHQTcgL2i9xQte8eNQkZIyOWGMzZ5tkat9HRTAKhRpD+qJMbWbqpWwc
KLh2lA+eYFavn24PL/gAjHpo+5BUpyHqWTW+0sO6aiZkMuHcNpl11Wm+86Si2+NF
NdpcMjT3J5EZBitc/mpVVTsxSI8WRVaNxodtnmKe6eo82CEHTWdcy+ko8TKtdm2P
6Vrdz2lTZLTJ+R32vx89DHVNRuXDVd3HTRqioAY0/eCXkO78+s94zb8u/21u2t2D
jR2n2yu1Ubu67n049kT9ZlB1WBJdPmEEE2K3pWgu8S3Gha/TLfOntTBjcKia0xDU
sjHoMLAb8K7MvgGT5w4zTYAkRsttFq2pSp+pd41DDTD0OE7nM0Qya+eThOyYbl0m
NHMJopMTH9oIztHutuC6wtlTWWUymFGlJF7YOw2/ARuURAvNT2Iqfg+X9B0MVPY5
YHs3oDLXdxjSdS6HO1KXXs2BXxn/uhVViz9no+pmgsVdBorqMYxgz3IIpUIfqUvS
ALDJTERiQVS7AQy8Hyj9WHhEeg1RTZXCXIJrxFunL6KVvhDNPDbB+JsnkdpPi2K4
1hfS0QwlpEAyxHGe77E4cqRjH7ZP5EXx1uIMXJGXtt84JM9KPeaFkAlrHp58+PQG
OaFPSWlCuXxSc2ckTmuNOUKoJl8gkUnvThUbKhptnoVY6S7FL5/7Xasmme7/LSuO
fL0aIAnMOv5AHkvIhBDx192xBHIKBvDghn7l9x1ghXzG4vZ1+h6TWG9/VraSG1BP
02OQW4j1urHLWqBJn43kRqoPc+QnERiz9pTLsOtmdfOvBFvLaryHl5vhmnlp4eXQ
1PK5htg9kGRhWP15I5997aZcpC8IYugwHPfK+w1TgQM88SutHw2DGQxfgnPtCP6o
AyyRdN2+Bzl38fCVnuI6kSsERb87Z0KrgRYv3jUBKRrztZK4yE+Pg81NoWCedIT4
u1OSyI2TPZIbIgBKl50F1YkXolzMUkiiSbq2GQq+s9///10Os1jilCoP4hTfsWT7
CvyFABiI1wlJvGkt1Wt5zhu9QOeQ9P08fp33me/ZVlVRLOyw/dyIOUAMFTcYmitT
0shFajqRaMwqiQ7zWJ9DK7/CZI46/jGgIasIPqVil/itDBN6apOBi+EpcXgToiH1
dEGdd0e9hCFwBgtyb2ajbQQlmvsZ1TnEI/rbMLTr8YsS5AX2Je0eOuRgJFNNvjUl
bsixFVEoKeAy8BYUTwLq2Epw8ctGXiMEdDFXzupSIoHurDiCG3RX3eNBJQSwFSE5
KCHnUFf93m16/+TS2N0VJwFP+BeIfVLwwssLQM83rsy0wntgT+QhIoqSOUn++3UR
sj/gOgxMF57V7nwI40rxBSpWdnJvMUB/VHO+fNqa2fSQ3q7L5q7jNQaM/zZk+hhz
uV75KWoyb/XTP02q8z0YCY/zCdZRS8NprIr44NL6zw0YCLRZOKHVt8oV7X6hr6iw
am16wwW0ilAbGSFAEh6y1c7qgdCep1G7Gi1OXgKZbb/ZRUEl6Qbyt6i8LQIVBOZq
JmbB9hpAGR+lmAFA9qtSU8pgnOucAokYLq2lquOQUO1XETdQjkaRGB24VXa5BsOl
QH3pKZKSkVWpELiAikheRgKmZnsf6/0frRyvg0Hpg7rU2zkIBKxt9GkvvWgpptHx
5Vg1lW8VFV0mw6F6ypYXYw0xk6aQzQlL0H0VfAgITbvMXT1wJK4udtYoEk/rgMY3
iHMm/kOSTZduqnOf7fA+H+5h4DZQjVJG9tb/JSEuAdz5OCbJ9jeNzvTpARLTBSuJ
AUtZnrH91nBSPKpAGXZNmMIGCbSZJV4XpTbrHV4pZmJS91M/kJ9EGXxEr6NCFTcJ
CT83uEqBOXfoz4zyhscCnffweLZmjbjfFZhi/4wQ4AEuF7pJ7sxJxpBR/y4yU10s
vXUfeAwOXd+mTC0XNyeUj3gdS6dPOEvN6kfPGhn46QEmOFtR2Tlvkz7AUPQYTTBe
sibbhm/6eCoMLHGq2Yaspbj+eg5ZnMAAQZvUumQ4PTj+yYGTfWpl2YtG0LHwtV44
V1FSGHnLC4B5G2JAnX81PSC0iaLUiL1HQDfMADKyuejiH/hXpEHoqFj7a6xBVwCm
GIeex0GS6du29CGzt1YIP6NVCSXH3NcF1zIXAwwTQK6e1TWvXHJTYzukj+Ld/6+X
h+GV/HcUWgUnt+GIk9zCbGIK5v8faZ8meCSoVD+ECxaMNfTaZPw+LbA2ggZ8ImSg
G447Bv2tyctFr9+vmASkygZ3tdZdvNT14CpiDPnxdfxx+7zedlc3EzheDZ07AXwE
j1waGAmSWkASN/G8900+sRiEbzDGMuxmSvWv1BoByK+u9iBcmJwhYCYiV05jjlDx
q54e6Df4Zup/bPrs+kPb+lnWJRUJ4Tfm1vIkWp7YrSDI0af17+OoaGvV48qNE4JF
cDyGUAzyMbmJ4ajbHphpnDcfISogIbuyvT3qK6gxODBtkuaQ7tY97TS/HJIJ1+Dw
o6p4g4ivbVmA2g5/D/NKW8zGHvaLLJ0YlyhQV9UAQY+IAK0nActAQTQTt2mzvpcX
nFsdGhwxAyywml+14KsMJSiPuYLkjvOt9tPvFWMTrGAHxXjc+/efc7kNj2Ay2+P9
9fs8dSlrvd2JkbZvm2vRN7PGp3/kGmUDNduOv8np/WHMFnQkxT8XgiSVKvcgBeMy
ChtQtHaAiYv00PBajYc0H/bif89tZZOmDwmvhBHOsWCQdTOOdy/0soTn4OMyAuGE
Vm8pmwU6f5kUJ5oy7jQphpzSUg63/nXsfArNCR1ekRFfJkrxAQAOaluLD5HEoK/r
FL/yBMXQ009SMhqSxOUcLuMLov4oZ1Cfd/rUIlVG3Ayuhbd8hD+sXiG2Xf2Hrg9a
KBWM6dwL1zaQwkIHoSevovGO5dSL9l8XTwKpf9TmmOnlU5JvygMHaDSgloq5bsXX
O44C70Xt6gSyFv8m6gR4bsSat5y1g+68SfBVw05cvbteDVAYhCD83Q4D2sTInpMh
4ex7Wpfqb4Gw3V5x2vcGe4VybVzUxNm5GKGb76FjlIMMX3ibcbWr9xTYgsUr3Hi6
iQT8uggytURTGvEQ05yEn4GcXoxenKJxJOD4iDtqwsMaUlEiYQd03Ah6k4nfw5Or
taJIgCbth2+HE46+aiHK7AubnPoBAgzMDS+WLe6yhFWIe07TLv2QqGWAejLwvfkt
L2WC5/foZcIKvu+lpyhro6m3RgjMNj+MQhG+7y8RxSKG73Rz9jFnU08IEzLPyDSn
rlNrhwWrxL6J7e7slcdCGih+knjsvwbHUPjXhCZONVh7Vc76ajYHA694Yrn9043t
CRqqJ/BY7ISmFL6dcBlerigw4IPXFSCLD0rEcwtvZoLoNLzGB6SnyCFeh40gKmp7
/StQHjGKOV4DSC4xhYVxpUuYs8JkPeFZOveEbRdyT8Bl1XkfzDyX4lVvc0mUAhnk
RBXlIGOQ6T7TZD8BsoLmOfHNg8zUF8LTNEoxG2koQttupMeThBljlsasIQ4YE1t7
fmcDDviQ10LMhQpeaxNCR60unVYU3U6YOoA2IfO/mTqaWstOaTLcGUoV74xzVJNa
Xe5IQEduJfK/yJ6hv0grMsd0RLBZalI1tRmiQ+X0aHFjoM/fIuIriAmf8gaHEpxN
sbTD6Pp/l5kf3FQepkTnAWK8nARxlYik6NdhRQHpqJvtIh+DR0gZInItKHKYQNpQ
aKSmrd5TDRMDn9orym0gj/l/zPK0XsPGq2XgwV9CKyG2cXWFB/Oa87QzP7cofUoG
mfDhtqHqofzGVZt7TC6FJnyD6CpLN/WKrtFBxqYXmZtKCVuZZOSDCGzqwJKxRdJj
eawouXKyb7JEnd6FOBZ3YT2CnnC1ZYRBnYvg3Bq0D7pxywoARAbovrlhbcKVmX2m
2WWvT6Tugh9/aGOOGqZqOAR/nAHQdCqM6zWumogshY5el69aASbMoGXFYP74T5U+
mLislcCj27+YkGKMvWVI8eVUq7M5qgsnGYHTH/lnEUE8WblVhuJ0rLfL/sprxNej
+2KtQZqAe+XVWWIMHhfRK7Xn9FDSRtkZlkGCT6N9ozzZ6aw27cPf6bk4lzjgrvrd
13SeVZxdoJt4iWWqVDSYMlkWBpQYKiOT6KFF5bZwRds4ij6hA0Sommk2MlDHwp2/
w4dBaqD0IO6WYbhCoK3/gaCrtArJxWmL8F2rBYv54gubxBv1PHSdkrIK1nIdPRIZ
LTSPxV39dOC35BDABACiBGEAvWFkBO41pz0AguYAcv89Uvy4gw2ODRUEAdCeLMG9
AFDCpywCVbchEEHWSI71UGlS1F6sZ3gyQwtS9094GysiMf7nQIA2Oyrc76HgFtja
E6gBC0mz2WnhQbP2OvUa647Us47pEC87AhvcQHH5AcyJL0JJY2OMytPYcJyAmvfD
lA5F/NgtNtjoGnVccpzL3JX7J5LGPT62HkhJZ8Ji9crOi+KOThc25o+ff7rj6lHp
tgdU6xx9ZcO/qJHiS+o6+B+0t2asb1FUDF5MpcuDiSBD4hvvk0kiZEKbxwhz0vOq
UOUM/DJjWTMliVK0oeI2VlixxPQ2mNymAp666tbA1Ir0GJx2oaX9Y5LkYk3RqycR
aj56689RGs4THuERMyPIfZMTOpg7fB6nfCYmaGykPJ1IUs0NdGAZbL3KPmzMMCCf
3ks/qQMN7muG/pdaxYh3M9o8D7+ps9+azOHvd09EnU9YVDr+IW7NLngkuDMhye4h
z4AYLg++VhMsYENBu7KJAXcuZshx0yMa6k6dhCa0v4lh0IX1GVNe+pEiCse48bJJ
+EBxqwr60q84ixo+YNmKzAPFGshpcNaRktEp6pzrR6TT8W02SqwqbeCpsFMT4Ry7
Yfm1gpvX8z7FnIgsDmvLvQYlF/+ipI0OXGyRJeTgJ3zCWX9fwEEP5fZsdtyABhKA
69gAKNYxslpER6zWz6g0R0Cc9CAsz7IwJIe7ryF6oos0ytMrrbkPVPeqF2RTOA5+
EQjR0cjgDeZ/LSfYDmPgU6iIM9KKlugTG9Tw/IMG5eGsPg4/0kwtd2uxXhioP357
7tkY7982ZGRLb+2LXWMpnD7rrjE6/6TRVDsmF7iT62MxyOJn3eLoxurgxcWV//xE
gAVTlEMDKbmV3FeyxFbC8DFj6v8ywFewj9c5jG6DX0m7UMfMEyizrQukCiP1OK8R
MYx7w4wD4d2i7Z6ZwW70yTqpXDwdnwHc74VWn249ebamqK+9z/qGOxgs7QUN5bGj
6zRbKPj7JESUdFcGiEpnXDrPEAuvkMahtY34u6elP+XvC/rzJZWfxvVZIpUaSuRm
BIv1mOyoP6H0Y3jTEXx1nlwi5yZ0YNq+s/j+K6K6qovJhD8PKcmxWbRPL465gmqd
hwWNBdS8J+ZdkrsMOZpXEbRgD6J70+1y1HjgNYJ+nzu5n5gBEc9cft0t9Cin6lNy
YUnoIQ6CMHJNz7QVGTZy6Mb7rbpt8CnW7f3dg26bN5WiLZ/Este5Vq0XbFN0TZUP
JyEkOGhbreBUfTbX6+wsNzTRMUvAyy9etwTENvfZoMsqgA7Tn/sDSNEDpnnYnXVf
R8eCJtDOO8/oFed0kxun1K+TzcVDTY+UxYA8HijjFheLsrUmMcq8IfCzRshuTXNj
nlowN73mUFzWaKGrCLfbt4INvxt0LtUVfHW3T3MGxpsOYtvP48kfkS/ubrK9EK0c
Kvf4xEm9ujS6CuyeHP0duz1ggX+cgM4WPVC6a9Qzi1LF+mYt3xzfZYQMpYKqauKY
hwFhP+QiiATXzD2PCzzf2VP5C9Nqb2wyc+BCqs9GKxhMnPTiPadSPZOnoP4GZ9zE
u675cDXlutj+cagQFd2gotApx94aDnKDgMLVZ35E74SsldW74EGqaxEfvDcS6Aar
OIuW56Aqy+FnOGF8JrudBCOZ7EDOfM5Py5T47DfaEgR9ZWTpdtqtHkoUBWrbbmAE
GTob7v8f1+alIy3KZsLoFODDi0dTP3TepFUg2vwk0SGYglkhzM5f2+4eIP2KOMqY
0N8B+W8ph1+JTUGZRYimw9NrpwUa3ICWPOtzOEmyjt/o1sBn/43luEcXtCJ29Bds
W6OF6Bf6r89a7zYy3xwOWNUiHoyRQahWW1eQbnc3O867G5Wvs3VXO8yVptAzLzH0
Y2CBZYBB8EjOM9UnfEt90JcTZRN8J/HhHqP4711yBw0ZNoOHxi/lbJrEaSsb5aGk
YT7RD1KSmUuz8sM/BUxzAK85tiv5hid4y79nlYolqMhhY114h+0h/z3EcGDCZNbm
iCWAfw4I6+k4YUyvDhws/z+YvwVDVmJku5GnQmskzeuSlBVE5889w0rZgOkLiTpU
YpIoo67yxHeUXDxzeDE7ec+V3K+r3rSU88dFZXRfTTF+fqt89TAhSzYswiblxpy/
t9FXFxjJQygGuJcOKDX6bkyb/xUUamuKqtIuXRpA/xzdb9fsUBJY4jmBICHT9Nm9
9umcyE2ik69sTs3be0S39iGLs//yuKymKbXsdE0wNl1/RMkH+FaijjRIk7R5IObW
625H86qRrr1ICxtoVnHNezogjdWo2S/wTr97ue9vb6OVsrDFZkIqKs3PHkCksKGY
LRYaRMX+kKZprUWQ9WU4HWEiwDqp8p1BHzmUJOg8jaWnNr1H/ol+rVVmNTXnpSqT
NCaPkb9J77UMifg6N8/l0AW3GoZVRoB8eIRG01hIi3NXGoHUcQxL8KNXPRbTqaGh
fo7V5bxERFIquSeKVU2wwxo9k8B7gakxZ5kdAbTeSUl8AkdavyqX9fTv3pFIBDlj
BQEJKvXjZTzQ6c7CzOUeYk9z/Uw0kOdYKizAer1hcYmSNWOlz3j8baY8PI21QtmQ
PF9FRtbyGXVrp7pCXnrxBhsE99VWxMx4kQRztfl9PRCVxbGH+5Qu2iehYQjFt6eU
w0dbYRtozKf8uPyGscG4vmw0asIDDzQGfYX3RcstYv2TH0vtuTXZi+qjLVKDTwJJ
3eLScD9gtOJEVXkTUnBQ7z8FveC+/qyrhmaAaqJM7g28Jy/fJCBlzgbaXx+yNIOn
eZRV1x8KRst+3qa1q3MDXmTfimJ73xokgr06fpe0up/tYGrYkadDVVfLVfCDVe+g
YakcU2ipB1DaEH5gW7JMngR6NCEp4OYln4k+0SxPpPlvvZPix0CvbpG3kZSVdO17
Cb6SIeuPrnxwiC2yKS75jOxYXV4pC18ZvNlv1PDl9RiyMxR3GMpyquQCz4Pc3jVa
kqGl2SSZaU4USUSbqktYJL/jQGk5lvogmAjocWneplADOyVmOHVBoPvPJRU1xARm
fwN/ElwXnU+Y6UEpxx1JhWaE1eSd02OYUPFHpvjKhAF05l/ZxNYuxqyjUo5Swb6G
KGj70xrEKj/0WkrjTf903ini7NPSDA0c4LadqyhPKmAwh1nw8/EZ2JUb5CyVm2Im
HzhKW5K2SqV4PUOEZd2aoccZth0bLUey1Bgf/TcDW2fV+3Xs2azetDgvBaxQXjIN
RzMbd1tu28yWbWWELt99k3aCjogUqCMztJXceKqTlzpdi/BoA2MsnWTKbiGgY6tB
aDpDmwtVBrI0Z3ZUxx+gVsbAK9P6pDV03iOHUs1cvecwlnJQuB/Y4kY+I5AEmea/
dUrhrO82uUVqn9SmdN7ubUSXz2Qc9pNIhp3kt5JZITBzPRm8MSKgBjs+fpmiHioU
Ez81bTWfYrdjAmbKD0Q4sNZhrR5tqPEcjqysuTD4l5UEQ1RHpkiBAshRzKypx2LN
v5Vc4j7OsicG8J4uJixI3kZEFVAME3Y0UAho4AmVLwMg4wT1ury3F+Bc2ju6ywZ2
wGyGJiHRq0ZTYn44SjPhkWI1dlhfHIPBFulmBMm3VDPI1TW8WimqbO8i83WYVC+v
T9hxucMaLSZTvzg8uot8K5yK0C88ucZesX8o1AvCvBeP61mlP7Pqpilwalh+ntwG
ktGSmGAatj9qYdhwcGr34z370V/FfNQ6nSvshi0sYqSujPq9G1E5+L56JeV+Jg5b
yfVoIRaW+Th4MiJJYxZDs/qbyeUX5UGeaxrRDlLp/8FZM2ap4QwfwLQia4T/l9vC
mfkyFQoELnde8wHs4h6Fl8h6jpla6ttx8z4vElR/ge3mN4Hi9YqBEWMoAfOo/Ckz
m95JOqfE4EH+nYEFefWX19QaIKjcTsw2KbgYMPwhqdZWSA4Sd5ROzrZXd6FLgGu0
vOGwx7MQ2ELyzu/VZZV3FyfSg9H0y0ykEs5nGZ/eO+8fgK3rOwqGPWDElBIDZu1I
m1udgPt7GmAQb6tOstg/metUEmQsnThvOdx0z8io13jcVXsAgwqLMShBNVzJeMh+
41733WKBGEZBVYWpJ7PFTdivxaDCna7TCiR2MJXIyyynlXshoTRT67GvxVsgM4TZ
u7RW1MeF+g3BUjQMdiFNsGFz1gN8N5tO0KjcSE1X/h+V0F4iQPtbyc/bBSWg+l7d
FBPsVcXJAGNROtbfrVxjH6s03FV5TZY3P5+z9E2AEqmyjleLXeY7uuY4QBuwVfzK
K4UhcDO1bbx9aHfefXfV9ezPmjLWI5TccHLy6AZs3TZvVMZvJ5TvwOYOrH8J/WHn
EbY7++jE3nKGI5qGQWZVRMKGLAOP/j6XVlQ88Pdq2eMP4llKA5brNFk1ZnX/pV7D
GEw3zdhm0ePSCItWhu3kFSBP6tu9//qIInx15zIAaWsV1V5fdUnk+SRVb4QwYj5a
OGRLV4fzvpS/n4B6VsdhiFYcVNCcj2AiuQIYdcp/aEK16gfMpC+gaZZwSNYBHLkY
SFEllEyDQJuh+I+iOjpznyzw3omUxXr0/nDPrjE6ZdFk1xI1YDdVUiruxiooUzfX
V6Y1KnDduPCgpi7Nh74rnnDdM4PVE5BW7xrjIbLMdhXiuByUXv3WwEEpUaziJgAA
GH8HItMeh5+XEheizLOEy+9y2WIo3ZwSM+RLeeL7J0z5MLQgUwimwAWAVna0yTfk
rGNPpgum+Nye27CQwRTeng9ENEkmujJuyj8TbiYvPSjStnkqCqKCV601wRmyYBh9
Hj+Lbfj5FgCYQTVOJzI9c8Mj48bm3APsIXvm7svBIfORVtUyAcMK3pViYLALXXqv
I4nl/kG3++NBvCOiEsYCKzk3NTJv41N7rP8TNTn3gFU9+jo8uYlo1ZBNcbIalOib
/8iDv0BzigGc/+rcgjz7rDGXbM+doMW1lT3oRLWm0s1L2/6DM8nLL1lADJSj8+t+
c0wibkXZznQlz9XyEgzSYsGFnzayQEly88CQyDJG09s6xDefMcjEBGNlz66Xstdp
4uxzOMRjCvL6jqLxvLyZU+OUGqsn0dcTHvRy58WMCU7z02xliBLr3DFc82Tw2vEV
XqVA41kZ+QX4h+c/Ndaime0hoYt60hQ9w284m/+p73te9Vp8/xW9A+tkZcWL1woS
S+UfFd8r6nQ0rBGBQMqInmzNEUqYorhCLdQmhLfsm1MD5lZz2MFOw0dDQXqlL51/
SDmEVs7rjexRg+XSc9X8rfhmzya4zQJIvizSPpV/sFE1oro84x/zZFiBup6EWhOr
0KszjfjAOSU9j2rIv6X5fmJ31FjNO4dvuP6SnDYmoxCvD5GJod4lIPCpfkO8u9zC
KF+3z5UdUNYPjvbWwgt5S8wUEGn7BOjE9vsUzihgjvgtmV5e+ob89p4QVdIyhpTs
TngaR0Aerxa21vJ9J1dPhvZBFtpTaEKZ4QTya+J3ubLMZutffsb/gYxfWvZbXdYe
IWEINjluTvJRLi5ZSXaCFo9C2P0NOkTtpyiqn70ujyf90uM7R81XfN6MLWN29WVV
o1KHfpXykzXiZWlBLYbj78yiu5T0K3mZtJsjLfWSIVigknX42c02YmC8/uVib0hU
va0oP3liCxoq3Db6W1LYa6NetgbQgR6daHuITv1a45NAoOpBqPDPBIGlysNZ8zOV
14BKnrFrwnl99AGXFmuF3wcc+ZU9A6nA8Ez9905VCHXhiS6cmQYxhE1PAhnZJz/e
AM5xD3vgGxnOO9N2JtHc/brn5RNU4ZicokhAtL6MRo7GVf0rmfruzXNAWJp91rNo
ifAwaLdi6omMsIssfLNYQMJ9ycLXerA42cyJoJ6vdTXvV50D6lUysC/9hvevvJKZ
P9aFNfonNaHW0lYJVb6JHLlbhv73WF7eXjgQ2MQmA16fvufmTT9+RDSlnOqJXjP5
ypt9cf3Jhx7WEFQb5N66fZg/LuYF+2uZ6DNcePC31EMXu/grkryzRxkm1Bbcnsxi
qEFnVxrZby2EV1mHLPbyGjAF04qs331mVMnwEOrUzT5IO0GMuwwKHdas+eXzEkXE
uK+pQZQuu7VJfXke3MFr7o04pRQoTukYOOF8JOswN/p3zlasObEev25zR4xZs3de
cLEonQQ1SeDlgRksNWaeqMFpaJ9N2xbGYE4ZHvunGc5O31wtJUa5pIKRYg7rNMJN
955Wqn0aA6AmmWFojaNjvJ1dJnL39p6aEVviaLeP9O7EsEzNcR/MUSnbLDTyibxQ
i3WVNt+k3Th5m1EBZ6HnOHGyC7O5k0hmd9lSfGM4FV1jYoYZgaiT8RJhGwP6EQa7
JP0P79WhTP82AUA1m7kgw8HEYagT7zNfU1WeMDIo1eXXAiU4OC28AegHKd8rvR8Y
2t67kh/un0wARyZ0uoi759bpz14G+neRYCb0mWWm92naBOpoRNbOChC2J5dky+Oo
V2ZT9uI/G2MyXJmh3hVXOjJNp9CcyJf9UbKWVev5eRLufTerafFGAXxkWm4Cga5D
2Ukc0ws9OA21wEuOmrHC8DeBCr/dhqO6Ae733eh54fsCWTBfpmRrK8PM3baKraPS
q8rg/dyKhKqBcqgAvDXqzb423NrZT4Ycay7PkwLX2zOppFQauWMp0bWVGobTTN+z
1cJErUdn7nk4ZKZQ5+2dlAY4ae5zucTnBiv/lMkIvaECgMZ4s7kFW1a+QodTmCQe
2A/hoZB6FZpTUxYtvKWCpW5LMRdz/HyoRt95U6g1MDYa/M07Oas5LYqqXIgUDszm
9O2vg5lqlqtnlBRTkY1XF0TkzonScbn4S2cJwKqsVDGgsbEggTBA4Fr0u9rE/d9Q
WjKITK4p2z4vRTAqK4+3LKLILs+tAc9uKMXyp5sOMO0WxzrTjKOnwFoyw9r5qpd4
HOFxoCqACAqeVShOWl8ja6NLzWqEBdYeXXLLtgyf+Itt+lH+5RROWA3lzBvGGlGO
SI2JgPqnZSgf4E9rAwHJF7o9r8YUIdSVSLu8TpAlwCFYUOGIgbmBbxb48IcfYwF/
js2G2lcD39FkyZzfvUFX0vbcwnN/84Yz75I5r/ilhjMLHFT5E5RAn5WvFtrLkfBQ
8AlaOKpxp8LeJIDFMRKHeEh+zzloZ63J4VfrNLOe7CUV2zgQB/3uZhgjQ/U2b1tv
xUIZPWhJYfVtBgnjVz47hlEAF8bUxrjT3V7ILX8hg5tl/uBnSWrOWUUoFbSE05Bw
iPjSJRrJAsWmucB2WfCZrUoIFYnrcicmTfSICyoPJ1UV29AbIg8/P/yz6lIKoaRK
YCAQ832H9pW8VYpdw67tKo3pLpmKtHwC8TNL/5kxKBe5nEsVAA/DzQ5H4JNSuQ0c
WSsj6m6gBy/Ut8K4kw/gYFMF6na2CzS5VBRg10qMkNSb58ZWIET70FaAWVKiwFNF
UeVtc/VUSXV5dpEIagHVizhouZBU8iJVtsNbpgfJbwyzOFxCBz5R4/lyIavUO3LR
+dEBHKS/PQhFt94Ub0cXVyejJ7X8CvRwe7348FZhDbdVHv2shdfv68xbdo2h5IQL
A/zlaYHlf7UORMNmZUhy0zW+cWG/+0ALJ+cQWl7PW2jSqrQK7w90iK+NGAXdcKC5
zB6Z+dh0YqRsCbv4wj5BRvBvRgWdo/Qm7+jxpQL49N+6k8Kfcapg+cfX27OJoIB/
2BOW2fxh0SI3Or5sB5B7dNJjCFm9QrvWix3G3/FLmEJrq2HkXs+GErGTlgOoBR25
/CASAoLJBPPzdfVjeKm8Giq9zzAOqgkIkoENfVbWtKK/uIzz++hab2rGjbCweJ9T
z1ZSeNLp4wBhC0f3TOmNz9V8EsQ+JzBG5JlSsVqUBpRlJPc3JFPomaLttUAY4FWF
pJClBJPFKrRDrNwRgCUQUitJWTR1Rvv+cue140phot+r7cEs6d03xh+ddgfqYpCe
LI9//e5djcPvJVFBwCRQx8W0+LmxArT7n2CN1NZg1ktcmbdH9l83AeBsBVhDokvL
gJY86M8hh/y13VnJrfMKuxLXjn+aO/+ewqncaMCz9YiPaunf4O8LOLvtoXf+Fd8D
Zh3sUpaSKPwSSLKvDbb3btsfBC4Jwnoitazan8mCMvrtMqp9q8+FFqlXWI7ta8bz
9xDJnDhBrooiIQ2duNhlSZ2ygwby5CkTFNd6PLDv26gOvpxm8v3J5G3rE7lxR1qO
xQVQ3lDshzCyvNNURH1cmcj8oXMvGz5f0flKm/YBYWDxyVkGrTGSoQrsS22Qf/Of
oPLw3v6XsUyJgC7xtzmg44QlAUxczsV01iDn9pjGl1+l5uivFD3jo03ABc6N9qXI
PwO7YQ/OyRazPyRCwmOCmQXTkhQt7WIVd1ersjQ1abHw/DBfH80VPOCgV57N1V1j
EbIrt8rS3btlQYj0U8C3j9keDRoxDNl534LWW+Re4c1fZTSGzzL6ksdof6LP8NO0
FLiFuOvYKALu1dlXdVemzx2SaofQ7rENfByPTpvJAXTyls4YjymldmX2AhRnDgbZ
/yWxQse4xKAutcxPK2VtUBAdgLN2xThBgrCxb1Tn5KhzneTykuevuszLc9DTbGEe
kJTnp/CCp42CzRQ/QwOgZ50yaz5xEjZo5Q2oydTPmwtEN5wJeMRb28tal/f1GMCx
C4ZGp3Yub4AVawZ0bLdCdBpSbwVGMAVKft6Bzh6g6UgfGV4xMxHerX3GrkcehtX6
cDRt7TNq7ADkaR65+OwvkMGAEmbeBcz+jWge4vk65r+pkckBcfkN1KFydGOTB6Zo
4wozFEsBqkrNbnkSpCg2Cq6wdPx92WGjfGev36N/aoXhYYmY4t6txZ7BdYFdU3wY
cXxHIs9Un7nELZHFDYOAW6/8TBBVyWfyltLd4D9f8gM+iI7c1bDcQ8/peMwf9R+d
cNC3WekNFlqD3ZdYqEWD9GJEbkF590jjBngyLhnAicbvIn9BZMGxzYuF+sK16L/a
LlfOUWBxwaUGuypwuWc5MwGgP0w4LRD+I1nQReeizu2mVbLpXuRtDmCGmOumJEUf
qCYMEVlBRWRqg7Pzz7qPHAhynWFdVxkbL0Lu9cfTBSh7nJzbHETF14nwd7Hg8NSI
1LEDDPpJSmXVsr+08PaMtm9F6Jj3pO08b9RhvLUgJP42bSFqSMQe4GDXcV0OfcCL
Prom12f2xbYhOSJf4vR1bQ7UGFdw4dIv6+tP1qKTG1Qzp3Iqj8zjZZ55rr8JALd1
cVeoZ8/jpLzSV8jrWESFSCA6GLyAsSMVKRs7gGcWF7mjAPlH4LD5fK/3Q3DtPICu
N6jY37CEzAxOK1mzupy/Cy4h9VXlBiRE/w/Fsqc0x1jmRjRWGkcKw8VPoiQp10Sw
opcrxd5QEsc/vC4iVbJVd0o6bIWU/6s2t3zYublic13hvDGLSmcNITMmGUX4H9My
4Xip2BaW7XRh9tHURux2QDCMvX8OrX2mRw9M/admAWTjH3S4KaoFT8lXQTCZIXe1
rwkKShflEt7l1cTNyY1Hjpljiglen5lrMNybHGvfL/aQ0h20NJbgA+Va8w+PjpmE
vfKsQ7YgQGDw2nW29nN1eRpp+YQxOyARNmV2QnPnYaCzJhYhBf6V7rnd+Vu7mJFY
4CD1vcG6DRoOmitcattIMuiALMgIs2lETEqpP7meIl9EQEHmuWpws2AO2F/GSftz
8u8OdrcOA9W91wKwJ8VSjeLES873wj4Nnwo5bcNl5a01Jy/t47aIHIrt15N1E9iq
lunmHpsKPjDRRsno6FXmic5GtFE0AIFtpnOJ6o8qGiOcKqMT9kaMMfXWe1smObuq
AL9zGlcdZubah+tcPSP1tfkik9xXLf/YIn+2xqa7c9gPoZWCNB51bmeRQEwYXAM5
ApinRWveUPSCzcejmaNR5KqmkZc1Wl7CzCOanGJrpMUQA8JhpHwy3P25l+9vlos8
fTETPD/ZLefvzXXn4T+jnJHP9gc1LZNcu93peVQrNLJIIdVDUKmKz1gj4KREqxpl
4gKeqqA9+jb2G+BLkX73tab202dcHmL9X1TxxLq0IzeNIKkko8v2/97G1L0iLU65
aGQYIAgQYtSiQXPiCdccN4FEUxFD7m3VqdMHJ1UtoT3JLLh9C+frK3rNyhcnG9eb
aYILGXBJhhS15EkmMOXkasP7iZDBHwscWgA+hWUwG/RDNsh5uldsXjr8oO1DfE1c
bhhC+iFveIhISvZCVMlXRdBNAPXKnvFdY+f6Fwbyk908hAeMs86WQfJU3lSh1PpS
KaNcmBJ/K5XwYJy6t1YIoRh5PMB3E2HrGjngraDgpTj+WT++2l2rSUZq5u3zrp+i
EXb7izkyjYkLCo/viq0TQZCxJeBQjxMiXZC0XKhlL2e75yhUOPycC5fDzrVjYl43
uzUpBOXf8NbLWg1j60DWaXO8w0LHerjkLu95uOVtZ9lSx6KPvWsURplnNHRNwXUw
TnlSdO4J0e+GR1xt9bxhPFuv5At5CDwDdmNEt+xtJHws41nMBrTFhjArnVamXr3d
CnjUu1StYYU27p+3e6mniRIsGbeqJXfPb/gkqBsOHYbW2l6VaG3VBZrVqET2Z+AZ
Gh3zZObk+Tckj+6skKPCggLALSAW95z7MBJ0zkJB7i0dmJBGwILgpe0u/26CRlLE
m+xJ+c+WvadhGkFyOJFqyCvTmzVmYqa2HUMWEdhrpOMA5UGnIL5ioP0mP/7mm+XM
m1qNXwZGFBIYVOh8F/wp+tYMsG1PklZqnu+PlnsVV3UXGdNh/yiniA0quO+/Sxts
mLH/DMd6cPOjfFw1sQcyBm8rWOeT1M2OCeRF8Mczul8vZ5JedZDUa6rOCcuAr4CA
WNQRIH8e8AjYkuyx/tczTJ1PjR2GvWp7pInjTTa+4KUZ33EhFat1uWKSDcTeY15L
DRLT+TtlI8OfjTx+YD9cf2tcX93uIIOPA3rXZQWOQhGcIPptctCIKhzDW5COahnn
WN3RvMdY9j4eoEYkeKFGXPZi6OICNjgq02duUCceKAefPILD6TWmv9OwnN6YV0nM
JxjV8fdbWcphSRYBJViWEiIdbp0jmAGbHLTq2NCBFM8zWqDFus80I9fLelMDD7ZC
dzeo3XN7tvJZIM1RYwU8UhWYHgLOdPkdVTXAmI+7i6nh5ZKn0/zGwdevvjEpLCXn
SgLlH3eVvYYqOQzGGqO1Ys1Yl+yM11sRLlA1yyELYuCUZseCTudMPi3PnShRpv4l
qTvQEHzZD7FBVg22f4xN5DNfeJL1K8qEkgL0okm5hLIurMfiWh3VOrK5LBy0ckL6
HiG+okOr32qD+f4ijKBLt+pY6LeVToiPllQRveYMx3kmBfTHfbO23rLyEMLGrm2G
GxZZJAQaPNtLIvFke9FswxFM/v8VqB/lNG/PMkbg6JY5mB4uyl/ATSbKj+rLLcSY
K1JVO23b63YL1+Nt/kvyT0r4da+zKPRJ6iu7eUG7u/W1bpNyl5mhX8CnrM9wtMY4
Y4bqkfXY1wMMCUOpWuUqdhR7O7EBoBmgxFW0DCJ3V39gyhec068Eq8n7PXLa2X9s
XF4ksYYjPLBYHvZ/7ozhSbnT/5Sf3u5M7LDHgkKjdds0NpwbCHWib2nC3kdMPV5I
dXrqPfmII/0HuZXNqDYPEBC1MioSYNcvGLUZfOIWV6q60K0TTdeUwP0MVuMxkbap
/B8Bdhid+kZ/IaD7OUqoQPNu9bZzyE+0LwCIyIv+3yLqqT9NNJAv+Bhnv6mU9MdL
xhfiV8foNkMG0f5kLSr8sekAE1gZXlDuvgDFRgNAg8jAYCr1ilNMgFtajkbzmtg7
zndg8bEYIQ09IYZmViiFYFf5v3wLpHVjbhNo45aUikXNFJptp913rEClkFTvfIJL
LMT21ZOJ1WP3gcJAGs9kSEhIti7E0D8RoR4ZJ/nWW2mivfHfSuI0P2HgL+SZlk3l
Q7AaCUuPUix2svl+drXfIKgpII/ITOvIk+sl8VAHLm6ip38OPDLWb5g8GDIBSnnB
u6S1s6FqgBd+fpcrON3m7D8/EABFm98/vIdrX41D4zgUL6XZ2euug7ImV9iFstxk
RwKo7fLFmFwHUsCBluII9LhXRtBBktBXfFzKR0r6ueOixAyYptuEHZgSAG7BgqaG
XY/ed3igGs1lo9zmRDjWSSFGDcKl3ntgDsukphwglGttEXenI7oRAmv63cq0+mSd
OgOgq3h9WR4JZODMxCEHYEPjWIKATggDWbqBnKXsa8fBMk2oNIUjAUwBr6nxa5FF
DKiarvewd0cjmvNEF+au0jxLIt9W7xC7+0YgZVFwZ9aJJA3S8MG1bQ3mPCfBrwsJ
VgMjCfx3BwdEW+evCoQ/m132c+3TItO7b6SnJkXCuUwQof60bmYw77L8u5YMJWqT
8qT7a9XYx/5bc+ao71dHqZuTVriVLRS7ft1i9jFxi5iqIxptg9wCH8sd0SaSfYWx
HOKhhF5EmqFjXubgTsYdrm1PwUmCDAj4ZxGOlsc0T/kAnk4gcKCCCz6NDjdb19Yr
E/4W0GSmU6ORmKTgAsDn7RkXJbNkiEJlZQu2PwnWWsNKoILHW3M0M2su2N+DkfVO
HijsOWU0QIyjwK5tJkjRpTdVb6G5nIyGis1Jk5a5BKNY7XVB5QKpcT89LSwgvE87
AzAUWlAUh/it1x4PEGe7PAbfNgXnaYzz6zcfMlynBQaNmtj5lM1bHPA5MJS7Ui1D
YeTix59tRexhe5BWzD10DvTws1n1kD/ufvUqVp+2x2SjOyodsrQiHXd/pP9Ufo7V
fYKqgk1oJSXbYwp8vIeDsrG+HE+I6+YNs2YH0yth16nzP50+zZFCRTITriZ0Tk51
WB/s3gt2NmvcFTusjvrb1gncG8UoMt8biYgpJzPsQ7R/3bPCF1rxF8N2z/PCR5rr
xDJpUgLP5msMqSqA0shu9LhRi171cQsIR01wd/JJqp/23YenLHOWrF0EwA0c+0fk
16A9livChkR6HNZSVL4teoXuVbAocxap38eP82plL+GPx9jH6nRYO5YJlaWK/NlD
YP0D0KiUgtK+2xe8TdPgyBnnVxODtMmW2dIiv6pTD37ZKcT4kpYhsoS82p8PSwXK
PpZFahXSAQpm72oIkxwSlNDyoJ2bTRdHpOB8Z5ryjoJ2KY/zKhMqNEm8zAyJku7p
vwz8cvkqvMOwVLEvEfinhRXMLIt/zTYfa4v3wKA9S5Uv4vrhtE89jYWSJtvJLCkR
7PMTDTiN8M6ZWQT2KSwwEM9NAT6GIeXTs8DXFKR9BEiyAoARnuGcq03Z5xJs8D1c
BxI9TcpoFRpBoTknsp1A9eAELAjU80f9R78QoW9Igywup/i7zJM8lx36DeXjoBcF
SXotEcmvM2Or7/AMlU/r+Pp/XMtEV7sJ4dWp1IWbQnce+AISQlflWSkmsYsqUJXc
WdntlaIoXeshN94MhgzJSKA4A4LmTt4PAIqyeKfMt52zs6aBcUnt4BJIU2wEbOPV
DGZNNGP1fYZtBFk/0t8aGFCLbVjAZcMM5DsdhmuSbiWyUpQxRWDawRZPN5TZVJf8
nxvN4cJ0Si582EwL+3X85H0fw77V9tjPjnabIf87e71EoxUi9F0CQNTrXifDmfg5
Bpca1zMhXdrB76YWmJ0QID4a92AdP9Y8tZMOyGDVBANhW4cxr5xVCsf1tw1D8qDc
yCdWWJnwv+GrNnmUFv9SRG8sZslNlkycHLY8u+aoh+cK60gvcIphs1Jftd2jMF75
fA/ZBSZJFhgStKNPWPeAfPsby3l3r0DytiqLBuuQIo+BdSw8WiuqdP29wxA9BsSM
SNFoPvxN9WYHgVLnf3tDZOrY4dTp8iRcUMTFmxaIEQRPJ19aFOmafg73MILHiJlJ
/QDNWhiDxhfyIQSVzBkSfjcSPpTxP9mAtNEK6VIS0O4rgZVZSdMnRFvkNWk6Imh3
4BXtDrTWtjRE8qIXzFSjXfFI2anbXzlIuReAHcn6qvoZ4uzusUMOVp0AdsrZlZOZ
KvYhXBGOGN74S0Yq9SZlgOsFDFrIWa7XCln45alLW1SvpqzedQG0m9RT4zKfBz0l
erzigU6do7ks48ynRRPrWQZLd8WEuNExslLo92wQwYJ09hIkeSZcqTDjh8jeDyHs
CZhrVTdmWKzmOR4jIoG8BUejm7e7VOZl0UQxJ5uw0R+4CMDaWqEADVjsigF02LiW
kBvSFOTihQyQGELIRxYEIUg2BevHTB8Pc7HRm7z3krDZ5+qra/3Ydce0Wb0KBs8G
pXL4KyIEvnAgzVIN94cVUG8JHVvE7jfpstR1mGwhGzPDTfuQtkFU4DF3vgLeaezK
4XK8lSZdbtaO8qp0JKg9jv5MCa/QE6JMi5tQ2YbWXfy//zNrqsGZ9isjgrpiMiog
i072cH43F3u4zb1sz4XJJxnFvRRjSbssXhGoj0ni57avgYfBMIbBgrLvzI/EpBqD
ZZkqWkoG/OgWvHaqo7A1USMmJauCkKCU+W5CEFwvWAsVmK3igk5qATC731k73AMd
Ewlf0DhPo0N1apYFAbVWf9cgBav2aUnsrBW/tejeylsffYfqr3XmqQOsu+a49seT
vEoiNhwUQelslyQ4JBY+tiSp3U4JPlugXAOKQUoFV7GrehkPbrd42v1WI6o41/fg
FT6BMv9hYUd7rDCJZAADRzRuhvJZ7rpyVzvBDfQbJDRi+SyimXny9MHh4bR4slWo
TdVts4xJfIse/OVWLLu2jUrlOqXy1HC96+74g1mcP3Ukweh0Qu3zZMB10kFPyaG+
EG8shSUoLOqLW6fl7JtUgi6fEHYT9eUUhKVoEITdOBncfW56XK0KaBPneX0wY9j8
B2sQgDSFR5SecZC9VVEhs4YBe9a/KKgUhQVyP1+ANERE3XEwg6OVIiP9mJJ7VxMp
2pfZKL57L47kv6UB26+w4pLrmX/Qjs+lVlY+wPfjJrYQGe/d+gJ/XPDdUUTqf2jU
5bP0pnP5NgVafX+Sx6BEuxNped/P35Ux91ipjBUU1xt7J8oMk10gPhZwwPWLtt4J
XCJf3v/U11Dz6SgEbfClwGrChyN8xRDy+WG/m6a/wQ74TESSvI/cxrf4U3vWkwoD
v+MuS7W5Y490CkgCNGit1FMBjmE9KZYuwqxcVonEsMK/MA+vL40aJEbwXrX2Alcu
Y7m5TveDCEJuj9Zti6S0x31SELhDCCE6TjG2sTZlVElplrdNlxFM90/W+hrUMygw
Qzu59IFlOe3iyS+n3lWuG1RQVjfUnyj/85br8ipMLE4PBjU5BCFtXPsvQUpBtL8J
8JRr7YbNfHLx/jCvSeHPnMcgX1uwkQsSY01m7fdZmkQBsd5AU3NsRH5Z9+/hLl88
hwoPx7o/3ouj3s7NqVuhnSguWYnhaj+dhCJoEQGE9Nw+COwK8FnD6VSTLn5I5pGr
HurIwegkCWyUjEpjHsXb6tXHPkq4GmvdUYxH9fctxmzztFWU4L332TvjRTpN6jXi
JM6GvVyb3vRZ7XZnRvJ5vzYLk3tSKuHdhOyXNT95S6EUNr6fBxGsjScuNgX6AMc0
QIvfZ2/pOeDsGtqMz0S6mcqfrCX6MpEjvg7TXbwGsK+37RSifnphjvJDbav4+5Kc
5NYpXT38rcSAcELvxkTmJoFeNkEEKtuKlTYqbu/D9ybbvvyd0BfZdpSSNUourcaZ
6N4t97MBDUfYO6zU0JrFpHqvi0MksWBYm23XXfQIcQNRylj92ljmp4lVSrrvBc8l
TF9jmZFKmT7BBHQGz1NcO6/YecUBWqSt+JsWE6A9Eo+UbyaHN0a1/6gx/qYai8IE
xA73VH+3+PlShaCBnJj6B3DGAKmDuNt6LB41mcXG2m2E1bKUWx+AF0KGwa+i+BgN
6zukEe/sqDWueTBuhZ/SehccCPVGjNfDR3RtnBrm41jrP9cWg2k7Nb2VKHbrOgfP
TZpmcLQj8wPzDDfTDhPu+LUQBNF52Zn7GPAWzbBpHep5KN4a1ku+OdlW/JvOAwIa
qDkxWBpRfMi5t5L8g21y/EiVK/g3z0KMwuQNRxK2d93SThyHzQUZxUBTzhkSyyJ0
vWh4X1WTxgOyRqp/dj3KrDSggFzRjXzHclRaoElNu2xNZaj1fa3tFWTeoIb6CQ6Y
DiB0ui6HDBq7LIT4U9hE0Z64o6T+q7WagOPh4W+udczvMu4h6qNofPKFqjcmJEmm
dvXRXThAQS4OVr4RIZ8lXsCKquKOUNl+gtGVQyXC53WY4UFJ9jumZQKE6SJ6S2W5
LgENkm78XS2PAsCyf7Y82HYXA3Ad99K7N+XCYPx+rJJYQBdTX84JBLsxnEbOB4Hq
/J6LRGOW/BHuiSNVr6+4YO7MMSbMkXvlmbvRnp6/GWvRfPWdtD/0sVPSH07DtyEe
Z9bkuTZ6v6lnRdJZF4mQfQA4CCPUP70QLIoFafZsKwFk+zsZrH/aZ7+EjWYtHssA
/4kClscXZAzV0eIyEwnd39bMY2tBYi9F71Ykk4Q6KPXfRKLE9UKCoG/RtqyVG4Df
e1o/He8Y/VOVraOFK8iFIH1Mzq/ytsmKRzsNYG1/L9vMqVir9s+tJQys2OzSzPNa
GSZQymZMvwmp7q7183A04RF54P6Rff18YoO7Gxp+d1cARhJwQn3+uPKp2yPnjqVx
9F/GWPM9vfvxRWIwQRotOZeS4D39fZFISQufmliiU/ErpCjopzW55h+hIQ9eStcU
NHKDaf8XxdzFVRrInWQ1hkAmGPqN86PQWFVu+qWzZHmGdYCHKR0Lsj3UcoVXN/01
8wpTqihc5v8ID7QkVYHB0Jdy1tP+uVz6gxOvEVq9Q5yFnS85OTAp+jQ/Dlqog6tW
SwmcP4+M3UoTySR3xR0so+5CPO4KtSusskwaU0GpTnn2r4K9ne2GBazQpvaaXptw
uitqRXCCzKkwJFqfd6troxVM9qDQ6376LfghnBvIs79c1ix+zRmtYx/+jBc5HxJV
scgid9mUZVr8bAa/6WgOHlgLD+KlZtUnXbHd4QZvriAyqV039NIAjEwIBcZLMMCR
mE38qhX2t8X/eOdoL3Gs5oTN2dgSBQ1qBdNr+oj0m2oiiuHdG2LebUadUu6xApQ4
n/lL2Hd7xOrHn6gM+QwxdjHgFlnboK0usbe0UYE2OuuP1qT1GUL4/8i04X4mU7wz
Dj4PA1K1qzRcKiAAarHVgSMt9ccM0N58NIX78uTamFmALD307fwGLeTlp3TiAkdo
+qvdGK+aIklvGi0D74/Zp1vNyC/V+o5qZnHFMw3si4WHoXu6VjQtl8AEk5Y3CBy0
Ve7WJI0sN2Cortkf8mzQdYhiSU5eXNtAlmP1LjXFpvZReVQ2oNyRx9SvkmUDgTMW
jDnMcAliwHoc/gfOHpyKwa2LVk19LWIgvjr9Hq10WArwETPFNGNZ7l7qTY067tQT
5bHgSUCh6gySkgicQYySM885O5YP56XUfkRIjm2PJtwacO4MXfwqiYqCdyxK9OLH
9OsWYyVCU1xzRAOp5EfGSvgAw0EvLT+PTb/o2dUBd50JeBAPwpRkhhKk8a1IJS0i
w9fJiqyO52jiePcICNhyi1r6ip9pAFTG9osJJovCCdjDhe7pbsuKFDOnd3KCrmhx
OjwpLS6klIH5P97xDx4kd63xnGk+9+nqT6zU3RlDQXuwEKI6MeKxO9nC9gUytI5M
ctI7MhrPDeCKJn2OzPbCvD83Uv1/LaQwf/ahH2ICXqs+0lvxDVvP+2ECNJ8wMgUh
IXMngixCiqxPKUEFP+lPU9DVjJb3m7Z2d2XRfuPWt/eHdPsyHy1LxaWr9UaWWtPR
75ar1fBI2qD+iDxCmN/oQM4d6ccOb4Zg0uz0QHeOogTo7HR5zoLLrqh/eAERepIE
uJSCoblV5zDZ8chCXd3fYTTgsU0WtTBHjpgg/nkTWMG7hwJhLw8+TL95XDidjuxA
eSTSZIgf6uIRGSfRNqH3Pfy42XzBdmMy2O1lbivtQoKditVLpy/J1QgI3ZML1Ig9
ww9rrLBssC6uPtcnjKpebt2BrVJu+Y7auF7n0u1/Rb9iFMD41kPvT19RbFpl3cb3
IqrQmH/M14UZOEtQhct09TXDT4Km+rcFpXrf3NNccBgNs6JbrfdLU0sX/a+/7eLx
ptpG11xdZw8ZUKrGZ54TZ1Lhg97WXNkwhNz4Re043jg0t362JjU2Ia0Y9FBDHIJx
/ilNagoOVXQ6Gnx/B0kM/PRVupE5sqi9uuCWwCAjcZzHwW2fjs/ffkujZ8+YLyvl
2vOUwYQIhVZtNrFz2R2VkZAapn1mUprG800DLx/ZfkJuHPCy0y0LGMeN0DX70WRr
t7VsQqIr9kKEdhSMoDMh1J8VjHwFdjzE5er4iuq/Fuu6i6WdS9m2xTJOE4G+4JPa
8mTfNB28maSDmk2kSs7zTl2xFIQEABWi7IBYTvqfp4czMaWLmpdWQ/BOUWJDElxa
X3EJ8jAsQYwCMgdYrh5FSVmAkOI0BkD2UC5OP3NFIqWPU9oY4qht/aZObXhmJ5c2
DOJag/ErrrkpOCUh6xHyLURqFOp2O/In2zTY3OadhwRKbQBpwNp7qOesCQ9sB8rf
OYoKvOM1r0it+GY1w3MvIe1AdwMyuYna/33WtIGhumUksvMsEL374ZuJxyVPy1Ku
nbcwCrr5uSNoj+0ICJZYI0Ct7SZ33PYO9nR5EZ5xqvNtSnw5y5rczoOEznMrL8Pc
tALmDYmOY3l/HVWZF6S19Htg2GMSk4ciDUTbayLUmlLzV68bgKZq+9JlXHjGuj1c
7gli4JlC1ouhUjbjzSmN/QTLyShdbpwKpq2lmPabV5YdEIHR+11YSmMgWlX7kUpc
Agf3AMrXcDYJis5kLeLIZdGusmSTcPx0nk7LtZznbkGsxdVL4a+drFaZgNfFuZmA
SpYyHVZdjKWw2gGA9TouCAZ8/i1IceuAYodYLcXZU9fhWEteNUDey5Yh97AgCRnn
KkQY5xLpCQnjeUzy+F0VlRRxXMY071SAOTFwXP4CzB3/Z5/XRoBFv29z+BjBTRpy
JMK0wbNDQkjDxLm+rIXffzqGmB88WD2DE8pZrUIC6aodlYKsz9GXUOlwgxbB3Wcl
G3YIH3RNwqW7Y+iOfhF6oYS1dqG+CbaQlpJQl08GxUIGmJIJ0DsIvH+/zsZxAus/
rjtQy/NKaoniKAyzMNxxaFc0U++GbAberFYYqe48wMwE73zWqqe5wAHLGXum3zlH
rwCX/HZOlMrEk7nzgQjo2ezdwfq5q+7NinWGTwq5AkiY14mpGR8AxDhcvdP1im0N
ZIr3+/hIbXs3pBJaD1L5yieYJXRbuUa2VS8BcXL2UPs/eK4I2Luy/wdUDKrm27iM
2IfV4YUovctgYgv2U0PMSzbu6YdJxR74Yi8EfMsNygkXQ5vHvk5Jy2Plpn1dW5qg
URd6MWi8lS5i9Rok4dc3fbSwWmBM8SLBpfyUnJD/7UbEnbvQSfVxJSbve6vsFh9H
CGzncmmiGHbiqXBxHCpzLrEVZlyjl6o+C7RvMlq3vGM7w4dRT/NpnR6yHNbD4chd
uoEUS4Zw95sO+ixfiJH3RKnH+qXks3XaVe79eP/r8h3uZ/yzumXcscbcUbviPMED
EB7ZkFaBhs9w8GYP8HsH5BDiPGxzEuPB/GYofOpGUJONUUGzssmptzLaAgbI+XNX
SEptmyqMtXVSo84zTuB3PhFUV34CwNyP4beyQxSK/J+Kr9Rpsm1lxZA6gpnu5cLO
IYojioxjPBnWCLojd7shthlCrNKvziQvq1qOmI7RcPKJH1WKAbLE8cfTfui6XXom
SyqJDDM1DQieFjfHqMPcXmLrq1f5eWX4sIQXllgmvCXOsL/ilERX/Wd9u4b01o1H
lU6lNWqk4vMkOyzSF7USM+9vycW8KoJ04KmpU7F0kd65cZ/qNBJFXqmBbjfV5Ih8
InboMpWz6aBdSLxzG2CoKdAXBcyO2tkgBvLmlsSsHoXDK5s2hR/TuVncGxzHujbp
ixgpuuEdFL27STlBBNevny0ehDgMlr5ac+/bvINnwRf1kL1vGreLom2v+8sve6bM
SsZR+f55C/BSihOt6/1stfgnqckKZaDX62I1IsloB+WPE9ZHNEVRO/5xQ2jL2OqX
GN+xtZpVBrw/Ki+GpYw9Gl2cplQUYZSQhozOGjBSjXL/AKvSxg3lCUVYYbQCc13G
tqXApD1EYAeau1D8mhBv0hp0iqYpd6y3929+mMTs86qCOH2puaHkmiVj+u9FmXNU
YEzFazvUtYdMh7VFqDXWTJC3T5qpTmJ2OAW2Y5BXAyJVw+ei/XaDs8JKrf6ia8PL
zz/0sd5tZyOlVyoziekq64310l0+vNGpsg5iXO0ZqW73AwCyl7/ixNP+rOvGeW8x
M0WoOghgrsqHZfGLThU5Ynfss6PJWf0r4tD1lMF6c+QbjOHUgubqaQ9FXmEpSR8B
Y5SKbHMYjRlFWD3G+qpZf9Gl7oFn5m45Hca7+YBVyQS05mg6UVvfHtlPzCZvhLtN
0YpPRqg/g5q2y067NXczzF10Nojl+Ga2X9YprWw4DRjg5iZXLckbc0HPa28I/ZmO
qVxeVUhZJhDKYGZRDsPp2OrEC0uRfPhSAuVHdlQwHFZEDHFFwB43k6ZUlq3PA3YV
/R3l+/pYe/L7Ml/8i/TNjSvMB16LvmEBpQjhg7a0VgsdSmvOnGrXfP2kCxXdk/Op
n/mx5v0Cyburx+1PTftkCPqO1A79931mXBXq+IZr/btltm0+7Lb/WOUJU842QF/U
nJuOkSAy/SkugoZGvNdJHOkyK2js0cJKY0jwzzRdrUOuGwF3jdiyY79/cgjE1bvC
TdYLVsNOFx+l6XrYaGF1l7b7mC6lbxKfhi9VqkW3xAe6gKdEpQzqBSScZ6ew2aMk
RJrZh+QXnxXl6GiWX8mx7+z7T5nLGQIePaNp3nPGRTlh3AZToQoBBmlbywwegLHv
v7G0Yv4QKZ0jc7r/OqtdwMtOhzhnBxVVjWbxFPz58V1nS6A6WD/E5ZJdL5vKpsk2
qYbGcpVi0X8QgbLgCZJNNt0MgCF+iPE2TV2TCaZREqXU1ABCUbombDMe0b2vW+QI
2r9P5wk4lyy+0qVMb15+MSmY0IHIFxEaYe1BX1aDwJcTXWSobpmR7FuIYrv0QgEr
oZIgjFDSilTBXiymxoi8zUMJ3z2DT6IAXMdvH7HyRg+WO1kq7aZc6d0AgscUfh+v
bdqdZguV1IjzxmEsnjDl9cTAgDWt2Ho3DyH51UaMQd5pI1Hwj558iNSMBfrfbq00
IPq4WuSg1i+HMehfNwBget4/JZa8xXPgM5Hr4+zgNePIlF0GZyW33cEmoWzTXTOv
2+yDF//Xyup9pdo/8QYSygdXonBlOTgNXBBgWcNfQY1jpYt5SQqadpp8l+0aDNtc
WVxHOJUlHVKDaDSHGuE9T+92R56qjGfClgF2FC0j0R8gYJ47qB62EHQ3aytRlLLY
yvJwm/Eaifzc3fAObIn74ql/gqt4QJLgSqgklSjPlaIpG1dD12CpAwJAmH4uQ89T
Gsxlwsk4F/kMXl8nr2fh7jjtNfGLbzOda9cuPD2LktS710pKr6MEuBd0GKkniZZi
7u8ymK8UKfiBfyjHfGK8WOvPghAWm1hvCbpKtXG7vBFFKtZJH8Ninu+fsh4j8ACt
mog6meMrSqopivTpzP9Q320y2EloAZL6dLYprqDM1sjda3CbrHtq199d4iwf51XM
oqV5R/Ii5z3pMOL7TQwmpPiYSXzstjF5l4eIArRgXDMa4F3ph1K0LbIyHfe8AEnJ
487VCIJOKxpTkiGzhCZG8iYHpMsWSIy1unVBXxYBVzhFsamIi76ALv9C9jmscVY3
5Bi3x3dwKlyWimowDkuCLS4Xb1pEbMeglwrno8LAqnz9njQF+0EqTTHSfJNV/n1X
4qObfjX/gqusq7262r9cQREuAegHs3zB/cYjZ7K4nRGgoekL5O3phTwrW+wugmnL
4rGOgDwmp4K2s5VFr6NrGtSkkC20aWgTh05SAiwKfhPG6wlL9aCZLf3/ay2tpcWl
QvOU0Z4h3570omkb9LGvNI0AZOiDolTyYCpmR4JBYYO32HIn073EmNUY3lkcn/Dv
CIPTuit8AYoENh/j/xRh1XiXaEu1Z+Vsuh2h4qqM8zrCEW5NtQbNfaFbbZpYMW+q
qoSc13E7EJniIEetkY/Z277lZxRl6DAISyfNv49iSccW43wC8Twe5xqjSsLl0NeX
dBKJ5XWKGc5VyXJNHMKvIPW3VcX337FjOKp0Sy/ZsNSIvVll7arC10kVF/HzeuD3
fEO8//z2aA4mEyTznLOzevmWHI8pxAygPIIIvdsb5w3LfRxHJotvSNzKVbVvUgkn
HWx55cfynskg/PEaj27xVCu553C+6ZeeFkSCxKwbFICOcEu2IaFN7AjFoDV8tzCc
nBVpNDvIPMgAXngiwdJWkoa93waeAo15wcBt6rOzY6zyd1G3aNnZOdgI6duoecrp
2Xh47Pv3VvciNJtXSeRYaAN0qdEW4Zik6BtjEItLQUXfCuqQjDmvFxKBiBtSRNFV
eW0tXuSOvk6DaHalhY3LLzcRfHH5BJg5kqJDHa1EHJNwwKrSkU8HNPcXZnRfDSNZ
t0dgnjhuBV/Va5lNSYVjwcvVOB0fVC8ZM4nFZwBA9BKIhv3873crh7H6fSVvviXY
xlC2qjc7gFgqdoaHgiOxp5+Blz5lnSszaHwuiXfC3OiQGxDbprsUFFhdepi/8rIL
LzIf0BMyH9N6uQX9D3vs/yHvE42e1yjdFiRLDBDhwOdGsygw1swWGF3pZKzpR86H
9hUKiw4u7BW2j+cJd8ZtUloJa44bTCMp7zhSoFMtDLCpFIxJj18y88HBMSw4xVnN
y6BrfDc4YBLd5JW782VQoaqfNikT9HcK/FgppNnJmc1Ks/85arkmRf/YNBJVztI7
LAn1buNHOlgkEeTfVuXQskPtksyccjRA+tcB6eGFdggv4UHuoMx/4I1f0VM+xXJZ
p1W43jmi7Qn/TQPXjc+xXj5NVrECg2WgEjjk6EBPozNMzB0kM/P9a7BAG6LUUIUr
6G3cB4gc4Dk7DVmjI0rnYeR3VkVXDCPoRVtdq/dpygKEydNfsyWk5iwhDDH1BkGp
IWAJ5gfpMCicnVnhKXTp2eE6yjIcNUsf5+kmRcj4XckxIouHyUjZx71RVgnjRmcW
IAyXZ1jHlVCEgb53sRlkKp6RrWeVeZhcsLGvewpk9RdXhTpI/hVnzFHMDaBMPqYG
6vA/MsHr1s0xFL4Noka5gd/mLHQohzkElhJ9hFIHaWCrh6rO/YWbqfcvRRctz4qH
5QztjKZBkLW0NnIAlhWFtUBTp59Tv9039faZMSxMpvljqIeeN5DnIO26XZDYfoX6
YLAzXAgGdwx7hVg3BLT+cvmfsJ9N5uynmJ9EyS9/18Gu6tOwq07LhEPtksLF6oOf
8M+2MVhwjzExInX3LvGKg3tdyHEr6q9hqSekzDYmaemQmOCNDsu1pOppaTe6FBXJ
7kbdKot29R+hvRvC89IdBM1BT07CeaacyHGZLTInyU5JMufTJCyp4IZ4MSvNh9iM
XT6jPb3GO78F7HWtI+BC5JRjeB2+D4gect5uJYCnJkiP0WOas12M2jc7fFBWa/ce
IPdKBv2Y44Icyx/EPvzPWElRNQCDwVbRPbFsu2ub4cT4/wNafwjXO7WF0308vIvO
+p6m+REa69fk5E0MCfvIl3P13hFbjXBm6kD5Zm2wmxJGd9VkZNgQOdiooDlUXGC3
r+DYVXffNIcqOTBg41FKNa+F/o1mTCPXzh4/oWAj3Yh3C58+bw9YD4EM131E3u7y
RzcAJJB+Zbv36yaWRml6fAf7Vb716X391hBIJjU+lH4TPnZoCBO7WWYnj+UStmxI
e4AAeKG5NMo46MbVEj2kmzIEdEYtfGazmStvnfBATw10B7g37UdSRG9JmWL6EzmW
z7+UrQJZRM73oOZz4mPyTKAlPyGPZOXv/078c7ro2n74wP5n0hU2Ef8GnctdeLkN
HyQjNEI08ftyiyMfRPzZZ3zhQjyj1xauHTbdZ0BiqChNa0QKpWsXg6P8RK8LeGrd
iErIMJHMdGvjFFExCZFMNfBnRMpqMCD9lZjQjBygoOr01ZLXD1huzrJhfC1eLXPe
i+PJDNSH0MebDeuvAVI3Xvrg9VLUdeBfnCZDwZamNN37VL/7wAF1NtUbJsY61QWI
Q7VoRbFbDK5dCrJ34yLv586j6Fw7/Wp2rqr2Xs09EHTCfqVGx7bIhP88yj+TjtxJ
fLX4Zk47aoMVkw79ujTZtOOPm1hTlkvQuhAzdX8bZcAiC35ycSR/opt+G9wTNML0
O5V84r+M2QOy7Y3B9NpMlraeXIq3b3otVxuAkjrMhh7qVw6HVUvtGB/hu7He7eEF
7kOE5xbKQO/EWBRfdg44qH4CQboCFvSYKkrYAMaKUbPjrDREG4B2fL3xe7KEpseu
jJZml5JOGJUOGCUrKS5yujWMcgXAxXTCoSyNtOp5KiTa8Fow1Etnk1AAo+1ewp4G
BP/V7dj/pg7QpqEU4Wu3+d1ZpgjIFkWaXPPi2TuFilr7/bObFvL6n+LUKoHPHSyw
MnbI+bGlZBrpF1MqkMXnIbsNDDn6RKLbbjBPG1QTaGb9wZyNfe6e5BfRuVjFApAf
ebLPViDjoZpaHX/SCVcJnwiynkKriAvetkIEPfUY4cVtJPxdv+XBxCFn6JnsHu63
SDp2JWj5503CXbmcIoyJyySjskVzv2yXOCPZyk3OnMtJYM28whnJbx9mnusKh1Tr
7a2Q1HfgvDxsn4DBjAqWzz2pq7XeJDptxWF5m80EImqzP3u9YMXxtSeptdeBGyaR
2qeJjyhIp9+pFkC3BHf4HI+SHZXcnqM+/t1I6XzAkitijodBvMWYvm/vyoSWm19v
HGe5VXs3bDw1HrdlY0xjfNp7oGiy5Y6ROKJszl1Mjkc6inB5hT4uHlicgfGAARAY
+dAZsc+2lDf6eELbGjAYe3gp8Io2tUQbpe5Ai+G+eLJjWyhr/g3mQnm6x/kFB8gP
kNV0fgUozaNUMPih8JGIl3iJQMa5kfUaydCNkm5FVYuH+Q82FIaJpGQQ2FCI+xcy
FK+vw2aYx6ER86LfHzRF7HMhRbhcRI4pwYEzNLmzvCvG+VluhUEA8NuMxw99uZCE
YOvC/t1pyJ1h3ZqT+wfiqAqEiMuimOBr9oSfLZoPxX96T5HHxAsKqUg9VQ1ad4ib
g4tauJZxqXH4Lmi4/Ia8q/UuUiFCy65bpgIlAjYLtJ70jWq19hnSFMPjNm41r0cz
2ZibY3eR+5w6OEx/WSap6WpWRcPL+O4JCjQoCWFDWHk59qdUv6jKm6qLh8kFnI0U
xBNd50o+39QN4i+/tvFwDtuWua7idgkgUlUDrmAQNBuZoUMn2kBHBoGAhVS/bqaB
fWAIN4l438WPmSUIDhWYuo8DSVVyo8KVkkkEwgy6Whq1D5XFrvgn1UJF/6ePxsuX
0SpxDbqWnhTh2JWhEG86ypnc0gVbiModCZzFHRhih3M3oloOQw/ztejK7LL3YWyx
x8cQWBdsAMyhl2aXoBEQRyrdrgeLX3U0D5SJeEpNqB5ERJybyYOBYH5dMBeaJ81r
07XICu88I3pnt4V6Hx2RQywlXf1ft6ZjoC5KUpKz4/prLP0ZEfnW8ac5ETSa7eSI
ebQ2BSrRguek7RbI9u3pubiiLkYsz6cf5sfFUTNfe9BhDSDIYYwaJmndwmmUcpyo
CdYwuYyGJpLCiiSvCa8NK9s9nN9sBnThMO6fo2NKBlGHpzjh3rnau79LjOpNBTDV
PEVjxVNiD59O4eok7TIRRtXpKr46vBkaFuFghqPE9/pYBUQ04VCuVnl58rEWC7ts
RrASLU9wQY7CklZ1HM3yM/2IKM/Ryl5Wc1SAY1C2JHLh67+IoP8ej6jqyaxkWRVy
1zGmhXLhT2D6JbTZwk5SDtIuCmlwwoYIAu6HwUdPz1BAr/4yV7zYPDGjUB+r8JU4
U2kjaWkLKZxxn1jiiTwsc2WDbNrH3iyPmiCW44w5wX4usxKrZDnr83xQriPNs7XH
Hwfup2u+lsgxP6uSPMveIw0uY4Sj1Z8Oi7rjptC1W3qSK0a09dCgyZ8ab0MB0FzC
AbYqPKFQCDweIQev/ornKRPmFfaQ/1/IYwLhXW0Px6fM4B0af1eeUyF3JJQcZ+FM
vkrYmodmZ3Fv1Ntx2ShjxXoyiv8raUnXRuIpQg5hIk/xoDf6MFYPvQ85CAp1LjWf
RR02n4Mvo5iCwZqcZBSfI06mUNRgxEQtQMXgMFr1jXCQtnkTbChw/qdCDSd3ojkE
y8HKAVLFY64xuKnQDBMxt0umw79sHyMnVQ5YPRbOn+Ep2tcmfCysJCunqTkfOIOb
BObqiYkmodTd9+eJ3+toi+YZJtQy+BhpQ/yhU7hFf77AD5WIerW9x+ft/6uS3Hd6
dGnPnA/DI4x/VKN40Kd1niWof0JfA0eLli9BtNlJrW+P+y+ENsQxGZN196Vr2Z/N
nTMTdvJgfmHx9HyM+D+EJUwH+IdJYr9RB5QsW7FGuZpMp9v6APDFbqIDbAfT5gNQ
n12QU3E+aBQAZNA6Xf2auTy1UOPG6LxP8m7o3+wuxaI+jdi/Xyb7l1SL2Nmo4dz6
XEhtcYeT/EoxHlnyE6HLFmwg1zUegafiAwmDccPD3DULW4ZD8IXdsU6Mu1oz8d24
oq97IydCvz+7KFSu5bLJqOqrlcxv7Dpj2QVeHb4cjbpNn20fRbpifbQ2x9ti87yW
IW75vZJw6SU6qH9O3gHaHtcQnBBhTqZomMZZerZWl+Ker2PauhAU0e0jNqLQbV+l
T0uLNvn5x99DqExU/Ze7ZXoqk+uYC5A0XMe+SE7azjYc//97i99G5gOq6zMj0NkN
p/1NvdcVH3n8WF3rVsBYdGErcCIqHI2aESXITx/owk993AJ3Ga45Gzw8sJX0U5LQ
GLpi6SBCRrjyL1uyy6S7FAtFJT0if5Hnac6Y7MQjrLM4T9c+NzsauXlLvuXomLtc
fkNNcnFATYHmBjWX3pRauFwTbhcvsXGIXtZHjjhDUKzuvl5ZqQie20wsWQ4ZK/Pd
EGILZip+hrCRIfddVTriiRt+HEuu69Ey5pGlBE/QXUxzcMia2Nqb/m7Lp1NJZW1A
hYYMhY89sIQpsSUCsPI6Xe8QVe/Aqb9inZNJnjcvf5g=
//pragma protect end_data_block
//pragma protect digest_block
Rr7nYtT/imb+8ktQfa+gaLQlZEk=
//pragma protect end_digest_block
//pragma protect end_protected

`endif
