
`ifndef GUARD_SVT_AXI_PORT_MONITOR_DEF_COV_CALLBACK_SV
`define GUARD_SVT_AXI_PORT_MONITOR_DEF_COV_CALLBACK_SV

`include "svt_axi_defines.svi"
`ifndef SVT_AXI_EXCLUDE_AXI_PORT_COVERAGE
  `include `SVT_SOURCE_MAP_MODEL_SRC_SVI(amba_svt,axi_port_monitor_svt,R-2020.12,svt_axi_port_monitor_def_cov_util)
`endif // SVT_AXI_EXCLUDE_AXI_PORT_COVERAGE

// =============================================================================
/**
 * This class is extended from the coverage data callback class. This class
 * includes default cover groups. The constructor of this class gets
 * #svt_axi_port_configuration handle as an argument, which is used for shaping
 * the coverage.
 */

class svt_axi_port_monitor_def_cov_callback extends svt_axi_port_monitor_def_cov_data_callback;

/** Virtual interface to use */
virtual svt_axi_master_if.svt_axi_monitor_modport axi_monitor_mp;

`ifndef SVT_AXI_EXCLUDE_AXI_PORT_COVERAGE
  // ****************************************************************************
  // AXI4 Covergroups
  // ****************************************************************************

`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF  
  /**
    * Covergroup: trans_cross_axi_awburst_awqos
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - qos: Captures ranges of QOS values
    * .
    *
    * Cross coverpoints:
    *
    * - axi_awburst_awqos: Crosses cover points write_xact_type, burst_type and qos
    * .
    *
    */
  covergroup trans_cross_axi_awburst_awqos ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_QOS
    axi_awburst_awqos : cross write_xact_type, burst_type, qos {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

   /**
    * Covergroup: trans_cross_axi_arburst_arqos
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - qos: Captures ranges of QOS values
    * .
    *
    * Cross coverpoints:
    *
    * - axi_arburst_arqos: Crosses cover points read_xact_type, burst_type and qos
    * .
    *
    */
  //covergroup trans_cross_axi_arburst_arqos @(cov_read_sample_event);
  covergroup trans_cross_axi_arburst_arqos ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_QOS
    axi_arburst_arqos : cross read_xact_type, burst_type, qos {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi_awburst_awqos_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_QOS
    axi_awburst_awqos : cross write_xact_type, burst_type, qos {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awqos_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_QOS
    axi_awburst_awqos : cross write_xact_type, burst_type, qos {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup 

  covergroup trans_cross_axi_arburst_arqos_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_QOS
    axi_arburst_arqos : cross read_xact_type, burst_type, qos {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arqos_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_QOS
    axi_arburst_arqos : cross read_xact_type, burst_type, qos {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup  
  
`endif

 // ****************************************************************************
  // ACE5 Covergroups
  // ****************************************************************************

`ifdef SVT_ACE5_ENABLE
  /**
    * Covergroup: trans_cross_atomic_comp_awburst_awsize
    *
    * Coverpoints:
    *
    * - atomic_comp_xact_type:  Captures atomic compare transaction type
    * - atomic_comp_op_type: Captures atomic transaction operation type
    * - atomic_burst_type: Captures atomic transaction burst type
    * - atomic_comp_burst_size: Captures atomic compare transaction burst size
    * .
    *
    * Cross coverpoints:
    *
    * - atomic_comp_awburst_awsize: Crosses cover points atomic_comp_xact_type, atomic_comp_op_type,atomic_burst_type and atomic_comp_burst_size
    * .
    *
    */
  covergroup trans_cross_atomic_comp_awburst_awsize ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_COMP_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_COMP_OP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_COMP_BURST_SIZE
     atomic_comp_awburst_awsize : cross atomic_comp_xact_type, atomic_comp_op_type,atomic_burst_type,atomic_comp_burst_size{
     option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
   /**
    * Covergroup: trans_cross_atomic_noncomp_awburst_awsize
    *
     * Coverpoints:
    *
    * - atomic_noncomp_xact_type:  Captures atomic non compare transaction type
    * - atomic_noncomp_op_type: Captures atomic transaction operation type
    * - atomic_burst_type: Captures atomic transaction burst type
    * - atomic_noncomp_burst_size: Captures atomic non compare transaction burst size
    * .
    *
    * Cross coverpoints:
    *
    * - atomic_noncomp_awburst_awsize: Crosses cover points atomic_noncomp_xact_type, atomic_noncomp_op_type,atomic_burst_type
    *  and atomic_noncomp_burst_size
    * .
    */
 covergroup trans_cross_atomic_noncomp_awburst_awsize ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_NONCOMP_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_NONCOMP_OP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_NONCOMP_BURST_SIZE
    atomic_noncomp_awburst_awsize : cross atomic_noncomp_xact_type, atomic_noncomp_op_type,atomic_burst_type,atomic_non_comp_burst_size{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
    /**
    * Covergroup: trans_cross_atomic_comp_bresp_burst_length
    *
    * Coverpoints:
    *
    * - atomic_comp_xact_type:  Captures atomic compare transaction type
    * - atomic_comp_op_type: Captures atomic transaction operation type
    * - burst_length: Captures transaction burst length
    * - bresp: Captures transaction write response
    * .
    *
    * Cross coverpoints:
    *
    * - atomic_comp_bresp_burst_length: Crosses cover points atomic_comp_xact_type, atomic_comp_op_type,burst_length and bresp
    * .
    *
    */
covergroup trans_cross_atomic_comp_bresp_burst_length ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_COMP_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_COMP_OP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_BRESP_NO_EXCLUSIVE
    atomic_comp_type_bresp_burst_length : cross atomic_comp_xact_type, atomic_comp_op_type, bresp ,burst_length{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

    /**
    * Covergroup: trans_cross_atomic_noncomp_bresp_burst_length
    *
    * Coverpoints:
    *
    * - atomic_noncomp_xact_type:  Captures atomic noncompare transaction type
    * - atomic_noncomp_op_type: Captures atomic transaction operation type
    * - burst_length: Captures transaction burst length
    * - bresp: Captures transaction write response
    * .
    *
    * Cross coverpoints:
    *
    * - atomic_noncomp_bresp_burst_length: Crosses cover points atomic_noncomp_xact_type, atomic_comp_op_type,burst_length and bresp
    * .
    *
    */
covergroup trans_cross_atomic_noncomp_bresp_burst_length ;
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_NONCOMP_XACT_TYPE
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_NONCOMP_OP_TYPE
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_BRESP_NO_EXCLUSIVE
     atomic_noncomp_type_bresp_burst_length : cross atomic_noncomp_xact_type, atomic_noncomp_op_type, bresp ,burst_length{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

   /**
    * Covergroup: trans_cross_atomic_comp_rresp_burst_length
    *
    * Coverpoints:
    *
    * - atomic_comp_xact_type:  Captures atomic compare transaction type
    * - atomic_comp_op_type: Captures atomic transaction operation type
    * - burst_length: Captures transaction burst length
    * - rresp: Captures transaction rresp response
    * .
    * Cross coverpoints:
    *
    * - atomic_comp_rresp_burst_length: Crosses cover points atomic_comp_xact_type, atomic_comp_op_type,burst_length and rresp
    * .
    *
    */
 covergroup trans_cross_atomic_comp_rresp_burst_length ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_COMP_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_COMP_OP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_RRESP_NO_EXCLUSIVE
     atomic_comp_rresp_burst_length : cross atomic_comp_xact_type, atomic_comp_op_type, rresp ,burst_length{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
   /**
    * Covergroup: trans_cross_atomic_noncomp_rresp_burst_length
    *
    * Coverpoints:
    *
    * - atomic_noncomp_xact_type:  Captures atomic noncompare transaction type
    * - atomic_noncomp_op_type: Captures atomic transaction operation type
    * - burst_length: Captures transaction burst length
    * - rresp: Captures transaction read response
    * .
    *
    * Cross coverpoints:
    *
    * - atomic_noncomp_rresp_burst_length: Crosses cover points atomic_noncomp_xact_type, atomic_comp_op_type,burst_length and rresp
    * .
    *
    */
  covergroup trans_cross_atomic_noncomp_rresp_burst_length ;
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_NONCOMP_XACT_TYPE
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_RRESP_NO_EXCLUSIVE
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_NONCOMP_OP_TYPE
     atomic_noncomp_rresp_burst_length : cross atomic_noncomp_xact_type, atomic_noncomp_op_type, rresp ,burst_length{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
   /**
    * Covergroup: trans_cross_atomic_comp_endianness
    *
    * Coverpoints:
    *
    * - atomic_comp_xact_type:  Captures atomic compare transaction type
    * - atomic_xact_op_type: Captures atomic transaction operation type
    * - endian: Captures transaction endianness
    *
    * Cross coverpoints:
    *
    * - atomic_comp_endian: Crosses cover points atomic_comp_xact_type, atomic_comp_op_type and endianness
    * .
    *
    */
   covergroup trans_cross_atomic_comp_endianness ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_COMP_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_COMP_OP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ENDIAN_TYPE
   atomic_comp_endian : cross atomic_comp_xact_type,atomic_comp_op_type,endian_type{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

     /**
    * Covergroup: trans_cross_atomic_noncomp_endianness
    *
    * Coverpoints:
    *
    * - atomic_noncomp_xact_type:  Captures atomic non compare transaction type
    * - atomic_noncomp_op_type: Captures atomic transaction operation type
    * - endian: Captures transaction endianness
    *
    * Cross coverpoints:
    *
    * - atomic_noncomp_endian: Crosses cover points atomic_noncomp_xact_type, atomic_noncomp_op_type and endian
    * .
    *
    */
   covergroup trans_cross_atomic_noncomp_endianness ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_NONCOMP_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_NONCOMP_OP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ENDIAN_TYPE
    atomic_noncomp_endian : cross atomic_noncomp_xact_type,atomic_noncomp_op_type,endian_type{
     option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

   /**
    * Covergroup: trans_cross_write_xact_type_awmmusecsid_awmmusid
    *
    * Coverpoints:
    *
    * - coherent_write_xact_type:  Captures coherent write transaction type
    * - stream_id: Captures stream id 
    * - sec_or_non_sec_stream: Captures whether stream is secure or non secure
    * .
    *
    * Cross coverpoints:
    *
    * - write_xact_type_awmmusecsid_awmmusid: Crosses cover points coherent_write_xact_type, stream_id and sec_or_non_sec_stream
    * .
    *
    */
  covergroup trans_cross_write_xact_type_awmmusecsid_awmmusid;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_STREAM_ID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SEC_OR_NON_SEC_STREAM
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    write_xact_type_awmmusecsid_awmmusid : cross write_xact_type,stream_id,sec_or_non_sec_stream{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_cross_write_xact_type_awmmussidv_awmmussid
    *
    * Coverpoints:
    *
    * - coherent_write_xact_type:  Captures coherent write transaction type
    * - stream_id: Captures stream id 
    * - sec_or_non_sec_stream: Captures whether stream is secure or non secure
    * .
    *
    * Cross coverpoints:
    *
    * - write_xact_type_awmmussidv_awmmussid: Crosses cover points coherent_write_xact_type, sub_stream_id and sub_stream_id_valid
    * .
    *
    */
  covergroup trans_cross_write_xact_type_awmmussidv_awmmussid;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SUB_STREAM_ID_VALID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SUB_STREAM_ID
     write_xact_type_awmmussidv_awmmussid : cross write_xact_type,sub_stream_id,sub_stream_id_valid{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_cross_read_xact_type_armmusecsid_armmusid
    *
    * Coverpoints:
    *
    * - coherent_read_xact_type:  Captures coherent read transaction type
    * - stream_id: Captures stream id 
    * - sec_or_non_sec_stream: Captures whether stream is secure or non secure
    * .
    *
    * Cross coverpoints:
    *
    * - read_xact_type_awmmusecsid_awmmusid: Crosses cover points coherent_read_xact_type, stream_id and sec_or_non_sec_stream
    * .
    *
    */
   covergroup trans_cross_read_xact_type_armmusecsid_armmusid;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_STREAM_ID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SEC_OR_NON_SEC_STREAM
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    read_xact_type_armmusecsid_armmusid : cross read_xact_type,stream_id,sec_or_non_sec_stream{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
   /**
    * Covergroup: trans_cross_read_xact_type_armmussidv_armmussid
    *
    * Coverpoints:
    *
    * - coherent_read_xact_type:  Captures coherent read transaction type
    * - stream_id: Captures stream id 
    * - sec_or_non_sec_stream: Captures whether stream is secure or non secure
    * .
    *
    * Cross coverpoints:
    *
    * - read_xact_type_armmussidv_armmussid: Crosses cover points coherent_read_xact_type, sub_stream_id and sub_stream_id_valid
    * .
    *
    */
   covergroup trans_cross_read_xact_type_armmussidv_armmussid;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SUB_STREAM_ID_VALID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SUB_STREAM_ID
    read_xact_type_armmussidv_armmussid : cross read_xact_type,sub_stream_id,sub_stream_id_valid{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
   /**
    * Covergroup: trans_cross_stash_xact_type_stash_nid_stashnid_valid
    *
    * Coverpoints:
    *
    * - coherent_stash_xact_type:  Captures coherent stash transaction type
    * - stash_nid: Captures stash_nid
    * - stash_nid_valid: Captures whether stream_nid is valid or not
    * .
    *
    * Cross coverpoints:
    *
    * - coherent_stash_xact_type_stash_nid_stash_nid_valid: Crosses cover points coherent_stash_xact_type, stash_id and stash_nid_valid
    * .
    *
    */
  covergroup trans_cross_stash_xact_type_stash_nid_stashnid_valid;
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_STASH_XACT_TYPE
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_STASH_NID_VALID
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_STASH_NID
   coherent_stash_xact_type_stash_nid_stash_nid_valid : cross coherent_stash_xact_type,stash_nid,stash_nid_valid{
    option.weight = 1;
   }
   option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_cross_stash_xact_type_stash_lpid_stashlpid_valid
    *
    * Coverpoints:
    *
    * - coherent_stash_xact_type:  Captures coherent stash transaction type
    * - stash_lpid: Captures stash_lpid
    * - stash_lpid_valid: Captures whether stash_lpid is valid or not
    * .
    *
    * Cross coverpoints:
    *
    * - coherent_stash_xact_type_stash_lpid_stash_lpid_valid: Crosses cover points coherent_stash_xact_type, stash_lpid and stash_lpid_valid
    * .
    *
    */
 covergroup trans_cross_stash_xact_type_stash_lpid_stashlpid_valid;
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_STASH_XACT_TYPE
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_STASH_LPID_VALID
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_STASH_LPID
   coherent_stash_xact_type_stash_lpid_stash_lpid_valid : cross coherent_stash_xact_type,stash_lpid,stash_lpid_valid{
    option.weight = 1;
   }
   option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_cross_rchunk_xact_type_rchunkstrb_rchunknum_length
    *
    * Coverpoints:
    *
    * - chunk_burst_type:  Captures burst transaction type
    * - chunk_burst_size:  Captures burst size transaction type
    * - chunk_length:  Captures chunk_length 
    * - rchunkstrb:  Captures rchunkstrb values 
    * - rchunknum:  Captures rchunknum values 
    * .
    *
    * Cross coverpoints:
    *
    * - rdata_xact_chunk_burst_type_size: Crosses cover points chunk_burst_type, chunk_burst_size
    * .
    *
    */
 covergroup trans_cross_rchunk_xact_type_rchunkstrb_rchunknum_length;
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RDATA_CHUNK_BURST_TYPE
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RDATA_CHUNK_BURST_SIZE
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RCHUNK_LENGTH 
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RCHUNKSTRB
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RCHUNKNUM
   rdata_xact_chunk_burst_type_size: cross chunk_burst_type, chunk_burst_size {
    option.weight = 1;
   } 
 endgroup
`endif
  // ****************************************************************************
  // AXI3 Covergroups
  // ****************************************************************************

  /**
    * Covergroup: trans_cross_axi3_awburst_awlen
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_awburst_awlen: Crosses cover points write_xact_type, burst_type and burst_length
    * .
    *
    */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF       
  covergroup trans_cross_axi3_awburst_awlen ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    axi3_awburst_awlen : cross write_xact_type, burst_type, burst_length {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

/**
    * Covergroup: trans_cross_axi4_awburst_awlen
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_awburst_awlen: Crosses cover points write_xact_type, burst_type and burst_length
    * .
    *
    */
covergroup trans_cross_axi4_awburst_awlen ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
   axi4_awburst_awlen : cross write_xact_type, burst_type,  burst_length{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF       
  covergroup trans_cross_axi_awburst_awlen_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    axi_awburst_awlen : cross write_xact_type, burst_type, burst_length {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    axi_awburst_awlen : cross write_xact_type, burst_type, burst_length {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    axi_awburst_awlen : cross write_xact_type, burst_type, burst_length {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_axi4_lite ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    axi_awburst_awlen : cross write_xact_type, burst_type, burst_length {
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
// `endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  
  /**
    * Covergroup: trans_cross_axi3_awburst_awlen_awaddr
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - addr: Captures min, mid and max range of transaction address
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_awburst_awlen_awaddr: Crosses cover points write_xact_type, burst_type, burst_length, addr
    * .
    *
    */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF       
  covergroup trans_cross_axi3_awburst_awlen_awaddr ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR
    axi3_awburst_awlen_awaddr : cross write_xact_type, burst_type, burst_length, addr {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
/**
    * Covergroup: trans_cross_axi4_awburst_awlen_awaddr
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - addr: Captures min, mid and max range of transaction address
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_awburst_awlen_awaddr: Crosses cover points write_xact_type, burst_type, burst_length, addr
    * .
    *
    */
  covergroup trans_cross_axi4_awburst_awlen_awaddr ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR
    axi4_awburst_awlen_awaddr : cross write_xact_type, burst_type, burst_length, addr {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi_awburst_axi3_ace_awlen_axi3_awaddr_axi3_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4 
    axi_awburst_awlen_awaddr : cross write_xact_type, burst_type, burst_length, addr {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif     
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_axi3_ace_awlen_axi4_awaddr_axi3_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    axi_awburst_awlen_awaddr : cross write_xact_type, burst_type, burst_length, addr {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif     
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_axi_awburst_axi3_ace_awlen_ace_awaddr_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    axi_awburst_awlen_awaddr : cross write_xact_type, burst_type, burst_length, addr {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif     
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_axi_awburst_axi4_lite_awlen_axi4_lite_awaddr_axi3_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    axi_awburst_awlen_awaddr : cross write_xact_type, burst_type, burst_length, addr {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
 `endif
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};
`endif     
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  
  /**
    * Covergroup: trans_cross_axi3_awburst_awlen_bresp
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - bresp: Captures transaction response
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_awburst_awlen_bresp: Crosses cover points write_xact_type, burst_type, burst_length, bresp
    * .
    *
    */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF       
  covergroup trans_cross_axi3_awburst_awlen_bresp ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP
    axi3_awburst_awlen_bresp : cross write_xact_type, burst_type, burst_length, bresp {
      ignore_bins Ignore_invalid_excl_burst   =  binsof(bresp.exokay_resp) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
/**
    * Covergroup: trans_cross_axi4_awburst_awlen_bresp
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - bresp: Captures transaction response
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_awburst_awlen_bresp: Crosses cover points write_xact_type, burst_type, burst_length, bresp
    * .
    *
    */
  covergroup trans_cross_axi4_awburst_awlen_bresp ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP
    axi4_awburst_awlen_bresp : cross write_xact_type, burst_type, burst_length, bresp {
      ignore_bins Ignore_invalid_excl_burst   =  binsof(bresp.exokay_resp) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  covergroup trans_cross_axi_awburst_axi3_ace_awlen_axi3_bresp_no_exclusive ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_awburst_awlen_bresp : cross write_xact_type, burst_type, burst_length, bresp{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_awburst_axi3_ace_awlen_axi3_bresp_all ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_ALL
    axi_awburst_awlen_bresp : cross write_xact_type, burst_type, burst_length, bresp{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(bresp.exokay_resp) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_awburst_axi3_ace_awlen_axi4_bresp_no_exclusive ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_awburst_awlen_bresp : cross write_xact_type, burst_type, burst_length, bresp{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_axi3_ace_awlen_axi4_bresp_all ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_ALL
    axi_awburst_awlen_bresp : cross write_xact_type, burst_type, burst_length, bresp{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(bresp.exokay_resp) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_awburst_axi3_ace_awlen_ace_bresp_no_exclusive ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_awburst_awlen_bresp : cross write_xact_type, burst_type, burst_length, bresp{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_awburst_axi3_ace_awlen_ace_bresp_all ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_ALL
    axi_awburst_awlen_bresp : cross write_xact_type, burst_type, burst_length, bresp{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(bresp.exokay_resp) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_awburst_axi4_lite_awlen_axi4_lite_bresp_no_exclusive ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_awburst_awlen_bresp : cross write_xact_type, burst_type, burst_length, bresp{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
 `endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_awburst_axi4_lite_awlen_axi4_lite_bresp_all ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_ALL
    axi_awburst_awlen_bresp : cross write_xact_type, burst_type, burst_length, bresp{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(bresp.exokay_resp) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
 `endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup


`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  /**
    * Covergroup: trans_cross_axi_outstanding_xact
    *
    * Coverpoints:
    *
    * - total_outstanding_xact : Captures total number of outstanding(read/write) transactions
    * - outstanding_write_xact : Captures number of outstanding write transactions
    * - outstanding_read_xact : Captures number of outstanding read transactions
    * .
    *
    */
  covergroup trans_cross_axi_outstanding_xact (int num_outstanding_xacts, int num_write_outstanding_xacts, int num_read_outstanding_xacts) @(cov_outstanding_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TOTAL_OUTSTANDING_TRANSACTION
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OUTSTANDING_WRITE_TRANSACTION
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OUTSTANDING_READ_TRANSACTION
    option.per_instance = 1;
  endgroup


  /**
    * Covergroup: trans_cross_axi_write_interleaving_depth
    *
    * Coverpoints:
    *
    * - write_data_interleave : Captures write data interleave depth
    * .
    *
    */
  covergroup trans_cross_axi_write_interleaving_depth @(cov_interleave_depth_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_DATA_INTERLEAVE_DEPTH
    option.per_instance = 1;
  endgroup // trans_cross_axi_write_interleaving_depth


  /**
  *  Covergroup     : trans_cross_master_to_slave_path_access_ace
  *
  * Coverpoints:
  *
  * - all_slaves : Captures all participating path cov slaves
  * - slaves_excluding_register_space : Captures all non axi/ace register address space slaves
  * - coherent_read_xact_type:  Captures readonce coherent read transaction
  * - coherent_write_xact_type:  Captures coherent write transaction
  * .
  * Cross coverpoints:
  * - cross_read_xact_type_with_slave : Crosses cover points all_slaves and
  *   coherent_read_xact_type
  * - cross_write_xact_type_with_slave : Crosses cover points all_slaves and
  *   coherent_write_xact_type
  * .
  * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.1.6
  * .
  *
  */


  covergroup trans_cross_master_to_slave_path_access_ace@(cov_master_to_slave_access_event);
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE

     all_slaves : coverpoint path_cov_dest_names {
`ifdef VCS
    bins slvs_b[] = {[path_cov_dest_names.first() : path_cov_dest_names.last()]}with (ignore_slave_func(svt_amba_addr_mapper::path_cov_dest_names_enum'(item))) ;
`endif 
`ifndef VCS
    bins slvs_b[] = { [path_cov_dest_names.first():path_cov_dest_names.last()] };
    ignore_bins ig_bins[]  = ignore_slaves_list;
`endif
            }

     slaves_excluding_register_space : coverpoint path_cov_dest_names {
`ifdef VCS
      bins slvs_excluding_register_space[] = {   [path_cov_dest_names.first():path_cov_dest_names.last()]} with (ignore_slave_no_cfg_func(svt_amba_addr_mapper::path_cov_dest_names_enum'(item)));
`endif 
`ifndef VCS
      bins slvs_no_cfg_b[] = {     [path_cov_dest_names.first():path_cov_dest_names.last()] };
      ignore_bins ig_bins_no_cfg []  = ignore_cfg_slaves_list; 
`endif
      }

     cross_read_xact_type_with_slave  : cross all_slaves, coherent_read_xact_type ;
     cross_write_xact_type_with_slave : cross all_slaves, coherent_write_xact_type ;
     option.per_instance = 1;
  endgroup //trans_cross_master_to_slave_path_access_ace




  covergroup trans_cross_master_to_slave_path_access_axi3@(cov_master_to_slave_access_event);

     all_slaves : coverpoint path_cov_dest_names {
`ifdef VCS
    bins slvs_b[] = {[path_cov_dest_names.first() : path_cov_dest_names.last()]}with (ignore_slave_func(svt_amba_addr_mapper::path_cov_dest_names_enum'(item))) ;
`endif 
`ifndef VCS
    bins slvs_b[] = { [path_cov_dest_names.first():path_cov_dest_names.last()] };
    ignore_bins ig_bins[]  = ignore_slaves_list;
`endif
            }

     slaves_excluding_register_space : coverpoint path_cov_dest_names {
`ifdef VCS
      bins slvs_excluding_register_space[] = { [path_cov_dest_names.first():path_cov_dest_names.last()]} with (ignore_slave_no_cfg_func(svt_amba_addr_mapper::path_cov_dest_names_enum'(item)));
`endif 
`ifndef VCS
      bins slvs_no_cfg_b[] = { [path_cov_dest_names.first():path_cov_dest_names.last()] };
      ignore_bins ig_bins_no_cfg []  = ignore_cfg_slaves_list; 
`endif
      }
     
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
     
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_EXCLUSIVE_ATOMIC_TYPE_AXI3
    
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_AXI3_AXI4 
     
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE 

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_AXI3
 
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE
    
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LEN_AXI3 
     
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RESPONSE_TYPE_AXI3 
    
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ALIGNED_ADDR_AXI3
       
     axi_wstrb_beat_0  : coverpoint cov_item.wstrb[0] iff (cov_item.xact_type == svt_axi_transaction::WRITE) {
  
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PATH_COV_WSTRB_BINS
     }
  
     axi_wstrb_beat_1: coverpoint cov_item.wstrb[1] iff (cov_item.xact_type == svt_axi_transaction::WRITE && cov_item.burst_length>= 4'h1) {

       `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PATH_COV_WSTRB_BINS
     }

     axi_wstrb_beat_2: coverpoint cov_item.wstrb[2] iff (cov_item.xact_type == svt_axi_transaction::WRITE && cov_item.burst_length>= 4'h2) {
       `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PATH_COV_WSTRB_BINS
         
     }

     axi_wstrb_beat_3: coverpoint cov_item.wstrb[3] iff (cov_item.xact_type == svt_axi_transaction::WRITE && cov_item.burst_length>= 4'h3) {
       `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PATH_COV_WSTRB_BINS
       
     }

     axi_wstrb_beat_15: coverpoint cov_item.wstrb[15] iff (cov_item.xact_type == svt_axi_transaction::WRITE && cov_item.burst_length == 4'hf) {
       `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PATH_COV_WSTRB_BINS
     }

     //crosses the above coverpoints with all_slaves and slaves_excluding
     //register_space
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_LEN_1_ALL_OKAY

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_LEN_REDUCED_ALL_OKAY

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_LEN_REDUCED_IGNORE_RESPONSE

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_ALL_OKAY_FIXED
    
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_ALL_SLVERR_FIXED

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_IGNORE_RESP_FIXED

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_ALL_OKAY_FIXED_UNALIGNED

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_IGNORE_RESP_FIXED_UNALIGNED
 
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_ALL_OKAY

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_IGNORE_RESPONSE

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_DECERR_LEN_1

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_SLVERR_LEN_1

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_DECERR 

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_SLVERR
        
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_ALL_SLAVE_IGNORE_RESPONSE        

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_XACT_TYPE_LEN_1_WSTRB
     
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_XACT_TYPE_LEN_2_WSTRB
     
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_XACT_TYPE_LEN_3_WSTRB
     
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_XACT_TYPE_LEN_4_WSTRB
      
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_XACT_TYPE_LEN_16_WSTRB
      
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CROSS_ALIGNED_UNALIGNED_ADDR_ASIZE
     
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CROSS_ALIGNED_UNALIGNED_ADDR_ASIZE_IGNORE_RESP 
     
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_X_WR_OKAY_ADDR_ALIGN

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_X_WR_FAIL_ADDR_ALIGN
   
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_X_WR_DECERR

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_X_WR_SLVERR
    
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_X_WR_OKAY_WSTRB
       
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_X_WR_FAIL_WSTRB 
    
    option.per_instance = 1;
  endgroup//trans_cross_master_to_slave_path_access_axi3

covergroup trans_cross_master_to_slave_path_access_axi4@(cov_master_to_slave_access_event);

     all_slaves : coverpoint path_cov_dest_names {
`ifdef VCS
    bins slvs_b[] = {[path_cov_dest_names.first() : path_cov_dest_names.last()]}with (ignore_slave_func(svt_amba_addr_mapper::path_cov_dest_names_enum'(item))) ;
`endif 
`ifndef VCS
    bins slvs_b[] = { [path_cov_dest_names.first():path_cov_dest_names.last()] };
    ignore_bins ig_bins[]  = ignore_slaves_list;
`endif
            }

    slaves_excluding_register_space : coverpoint path_cov_dest_names {
`ifdef VCS
     bins slvs_excluding_register_space[] = { [path_cov_dest_names.first():path_cov_dest_names.last()]} with (ignore_slave_no_cfg_func(svt_amba_addr_mapper::path_cov_dest_names_enum'(item)));
`endif 
`ifndef VCS
     bins slvs_no_cfg_b[] = { [path_cov_dest_names.first():path_cov_dest_names.last()] };
     ignore_bins ig_bins_no_cfg []  = ignore_cfg_slaves_list; 
`endif
     }
    
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_EXCLUSIVE_ATOMIC_TYPE_AXI3
    
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_AXI3_AXI4
    
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE 

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_AXI3
        
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RESPONSE_TYPE_AXI3 
 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_AXI4
    
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LEN_AXI4 

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ALIGNED_ADDR_AXI3
    
    axi_wstrb_beat_0  : coverpoint cov_item.wstrb[0] iff (cov_item.xact_type == svt_axi_transaction::WRITE) {
  
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PATH_COV_WSTRB_BINS
    }

    axi_wstrb_beat_1: coverpoint cov_item.wstrb[1] iff (cov_item.xact_type == svt_axi_transaction::WRITE && cov_item.burst_length>= 4'h1) {

      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PATH_COV_WSTRB_BINS
    }

    axi_wstrb_beat_2: coverpoint cov_item.wstrb[2] iff (cov_item.xact_type == svt_axi_transaction::WRITE && cov_item.burst_length>= 4'h2) {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PATH_COV_WSTRB_BINS
        
    }

    axi_wstrb_beat_3: coverpoint cov_item.wstrb[3] iff (cov_item.xact_type == svt_axi_transaction::WRITE && cov_item.burst_length>= 4'h3) {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PATH_COV_WSTRB_BINS
      
    }

    axi_wstrb_beat_15: coverpoint cov_item.wstrb[15] iff (cov_item.xact_type == svt_axi_transaction::WRITE && cov_item.burst_length == 4'hf) {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PATH_COV_WSTRB_BINS
    }

    //crosses the above coverpoints with all_slaves and slaves_excluding
    //register_space
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_LEN_1_ALL_OKAY

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_LEN_REDUCED_ALL_OKAY

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_LEN_REDUCED_IGNORE_RESPONSE

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_ALL_OKAY_FIXED
    
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_ALL_SLVERR_FIXED

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_IGNORE_RESP_FIXED

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_ALL_OKAY_FIXED_UNALIGNED

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_IGNORE_RESP_FIXED_UNALIGNED
 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_ALL_OKAY

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_IGNORE_RESPONSE

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_DECERR_LEN_1

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_SLVERR_LEN_1

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_DECERR 

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_SLVERR
       
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_ALL_SLAVE_IGNORE_RESPONSE        

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_XACT_TYPE_LEN_1_WSTRB
    
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_XACT_TYPE_LEN_2_WSTRB
    
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_XACT_TYPE_LEN_3_WSTRB
    
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_XACT_TYPE_LEN_4_WSTRB
     
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_XACT_TYPE_LEN_16_WSTRB
     
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CROSS_ALIGNED_UNALIGNED_ADDR_ASIZE
    
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CROSS_ALIGNED_UNALIGNED_ADDR_ASIZE_IGNORE_RESP 
    
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_X_WR_OKAY_ADDR_ALIGN

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_X_WR_FAIL_ADDR_ALIGN
   
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_X_WR_DECERR

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_X_WR_SLVERR
    
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_X_WR_OKAY_WSTRB
      
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_MASTER_TO_SLAVE_X_WR_FAIL_WSTRB 
    
    option.per_instance = 1;
  endgroup//trans_cross_master_to_slave_path_access_axi4

  function bit ignore_slave_func (svt_amba_addr_mapper::path_cov_dest_names_enum myitem) ;
    ignore_slave_func = 1;
    for (int k=0 ; k < ignore_slaves_list.size(); k++) begin
      if (myitem == ignore_slaves_list [k]) begin
        ignore_slave_func = 0;
        break;
      end
    end
  endfunction
   
  function bit ignore_slave_no_cfg_func (svt_amba_addr_mapper::path_cov_dest_names_enum myitem) ;
    ignore_slave_no_cfg_func = 1;
    for (int k=0 ; k < ignore_cfg_slaves_list.size(); k++) begin
      if (myitem == ignore_cfg_slaves_list [k]) begin
        ignore_slave_no_cfg_func = 0;
        break;
      end
    end
  endfunction

  //  ACE DVM overlap case related covergroups for ACE and ACE-Lite Vips
  /**
    * Covergroup: trans_cross_dvm_overlap_arvalid_arready_cover_acvalid_acready_acsnoop
    *
    * This covergroup is cross coverage related to  DVM overlap case in ACE-lite and ACE-VIP and it cover acvalid=1,acready=1,
    * and acsnoop=dvm when ARVALID == 1 and ARREADY == 0.
    *
    * Coverpoints:
    *
    * - acvalid : Captures ACVALID ==1
    * - acready : Captures ACREADY == 1
    * - acsnnop : Captures ACSNOOP == DVM
    * .
    * Cross coverpoints:
    *
    * -overlap_case_dvm_arvalid_arready_acvalid_acready_acsnoop : Crosses coverpoints acvalid,acready,acsnoop
    * .
    */ 
   covergroup trans_cross_dvm_overlap_arvalid_arready_cover_acvalid_acready_acsnoop @(dvm_overlap_scenarios_snoop_addr_event);
   `SVT_ACE_SYS_MONITOR_DEF_COV_UTIL_ARVALID_1
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_ARREADY_0
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_ACVALID
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_ACREADY
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_ACSNOOP
    overlap_case_dvm_arvalid_arready_acvalid_acready_acsnoop : cross arvalid,arready_0,acvalid,acready,acsnoop{
    option.weight = 1; } 
    option.per_instance = 1;
    endgroup
    
  /**
    * Covergroup: trans_cross_dvm_overlap_awvalid_awready_cover_acvalid_acready_acsnoop
    *
    * This covergroup is cross coverage related to  DVM overlap case in ACE-lite and ACE-VIP and it cover acvalid=1,acready=1,
    * and acsnoop=dvm when AWVALID == 1 and AWREADY == 0.
    *
    * Coverpoints:
    *
    * - acvalid : Captures ACVALID ==1
    * - acready : Captures ACREADY == 1
    * - acsnnop : Captures ACSNOOP == DVM
    * .
    * Cross coverpoints:
    *
    * -overlap_case_dvm_awvalid_high_awready_low_acvalid_acready_acsnoop : Crosses coverpoints acvalid,acready,acsnoop
    * .
    */   
   covergroup trans_cross_dvm_overlap_awvalid_awready_cover_acvalid_acready_acsnoop @(dvm_overlap_scenarios_snoop_addr_event);
   `SVT_ACE_SYS_MONITOR_DEF_COV_UTIL_AWVALID_1
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_AWREADY_0
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_ACVALID
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_ACREADY
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_ACSNOOP
    overlap_case_dvm_awvalid_high_awready_low_acvalid_acready_acsnoop : cross awvalid,awready_0,acvalid,acready,acsnoop{
    option.weight = 1; } 
    option.per_instance = 1;
    endgroup

  /**
    * Covergroup: trans_cross_dvm_overlap_awvalid_awready_cover_acvalid_acready_acsnoop
    *
    * This covergroup is cross coverage related to  DVM overlap case in ACE-lite and ACE-VIP and it cover acvalid=1,acready=1,
    * and acsnoop=dvm when RVALID == 1 and RREADY == 0.
    *
    * Coverpoints:
    *
    * - acvalid : Captures  ACVALID ==1
    * - acready : Captures ACREADY == 1
    * - acsnnop : Captures ACSNOOP == DVM
    * .
    * Cross coverpoints:
    *
    * -overlap_case_dvm_rvalid_high_rready_low_acvalid_acready_acsnoop : Crosses coverpoints acvalid,acready,acsnoop
    * .
    */
    covergroup trans_cross_dvm_overlap_rvalid_rready_cover_acvalid_acready_acsnoop @(dvm_overlap_scenarios_snoop_addr_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_RVALID_1
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_RREADY_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_ACVALID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_ACREADY
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_ACSNOOP
    overlap_case_dvm_rvalid_high_rready_low_acvalid_acready_acsnoop : cross rvalid_1,rready_0,acvalid,acready,acsnoop{
    option.weight = 1; } 
    option.per_instance = 1;
    endgroup

   /**
    * Covergroup: trans_cross_dvm_overlap_awvalid_awready_cover_acvalid_acready_acsnoop
    *
    * This covergroup is cross coverage related to  DVM overlap case in ACE-lite and ACE-VIP and it cover acvalid=1,acready=1,
    * and acsnoop=dvm when BVALID == 1 and BREADY == 0.
    *
    * Coverpoints:
    *
    * - acvalid : Captures ACVALID ==1
    * - acready : Captures ACREADY == 1
    * - acsnnop : Captures ACSNOOP == DVM
    * .
    * Cross coverpoints:
    *
    * -overlap_case_dvm_bvalid_high_bready_low_acvalid_acready_acsnoop : Crosses coverpoints acvalid,acready,acsnoop
    * .
    */
    covergroup trans_cross_dvm_overlap_bvalid_bready_cover_acvalid_acready_acsnoop @(dvm_overlap_scenarios_snoop_addr_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_BVALID_1
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_BREADY_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_ACVALID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_ACREADY
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_ACSNOOP
    overlap_case_dvm_bvalid_high_bready_low_acvalid_acready_acsnoop : cross bvalid_1,bready_0,acvalid,acready,acsnoop{
    option.weight = 1; } 
    option.per_instance = 1;
    endgroup

   /**
    * Covergroup: trans_cross_dvm_overlap_awvalid_awready_cover_acvalid_acready_acsnoop
    *
    * This covergroup is cross coverage related to  DVM overlap case in ACE-lite and ACE-VIP and it cover crvalid=1 and crready=1
    *  when ARVALID == 1 and ARREADY == 0.
    *
    * Coverpoints:
    *
    * - crvalid : Captures  CRVALID ==1
    * - crready : Captures  CRREADY == 1
    * .
    * Cross coverpoints:
    *
    * -overlap_case_dvm_arvalid_high_arready_low_crvalid_crready : Crosses  coverpoints crvalid and crready 
    * .
    */
    covergroup trans_cross_dvm_overlap_arvalid_arready_cover_crvalid_crready @(dvm_overlap_scenarios_snoop_resp_event);
    `SVT_ACE_SYS_MONITOR_DEF_COV_UTIL_ARVALID_1
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_ARREADY_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_CRVALID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_CRREADY
    overlap_case_dvm_arvalid_high_arready_low_crvalid_crready : cross arvalid,arready_0,crvalid,crready{
    option.weight = 1; } 
    option.per_instance = 1;
    endgroup
   
   /**
    * Covergroup: trans_cross_dvm_overlap_awvalid_awready_cover_crvalid_crready
    *
    * This covergroup is cross coverage related to  DVM overlap case in ACE-lite and ACE-VIP and it cover crvalid=1 and crready=1
    *  when AWVALID == 1 and AWREADY == 0.
    *
    * Coverpoints:
    *
    * - crvalid : Captures  CRVALID ==1
    * - crready : Captures  CRREADY == 1
    * .
    * Cross coverpoints:
    *
    * -overlap_case_dvm_awvalid_high_awready_low_crvalid_crready : Crosses  coverpoints crvalid and crready 
    * .
    */
    covergroup trans_cross_dvm_overlap_awvalid_awready_cover_crvalid_crready @(dvm_overlap_scenarios_snoop_resp_event);
    `SVT_ACE_SYS_MONITOR_DEF_COV_UTIL_AWVALID_1
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_AWREADY_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_CRVALID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_CRREADY
    overlap_case_dvm_awvalid_high_awready_low_crvalid_crready : cross awvalid,awready_0,crvalid,crready{
    option.weight = 1; } 
    option.per_instance = 1;
    endgroup
  
   /**
    * Covergroup: trans_cross_dvm_overlap_rvalid_rready_cover_crvalid_crready
    *
    * This covergroup is cross coverage related to  DVM overlap case in ACE-lite and ACE-VIP and it cover crvalid=1 and crready=1
    *  when RVALID == 1 and RREADY == 0.
    *
    * Coverpoints:
    *
    * - crvalid : Captures  CRVALID ==1
    * - crready : Captures  CRREADY == 1
    * .
    * Cross coverpoints:
    *
    * -overlap_case_dvm_rvalid_high_rready_low_crvalid_crready : Crosses  coverpoints crvalid and crready 
    * .
    */
    covergroup trans_cross_dvm_overlap_rvalid_rready_cover_crvalid_crready @(dvm_overlap_scenarios_snoop_resp_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_RVALID_1
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_RREADY_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_CRVALID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_CRREADY
    overlap_case_dvm_rvalid_rready_crvalid_crready : cross rvalid_1,rready_0,crvalid,crready{
    option.weight = 1; } 
    option.per_instance = 1;
    endgroup
  
   /**
    * Covergroup: trans_cross_dvm_overlap_bvalid_bready_cover_crvalid_crready
    *
    * This covergroup is cross coverage related to  DVM overlap case in ACE-lite and ACE-VIP and it cover crvalid=1 and crready=1
    *  when BVALID == 1 and BREADY == 0.
    *
    * Coverpoints:
    *
    * - crvalid : Captures  CRVALID ==1
    * - crready : Captures  CRREADY == 1
    * .
    * Cross coverpoints:
    *
    * -overlap_case_dvm_bvalid_bready_crvalid_crready : Crosses  coverpoints crvalid and crready 
    * .
    */
    covergroup trans_cross_dvm_overlap_bvalid_bready_cover_crvalid_crready @(dvm_overlap_scenarios_snoop_resp_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_BVALID_1
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_BREADY_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_CRVALID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DVM_OVERLAP_COVER_CRREADY
    overlap_case_dvm_bvalid_bready_crvalid_crready : cross bvalid_1,bready_0,crvalid,crready{
    option.weight = 1; } 
    option.per_instance = 1;
    endgroup

`ifndef SVT_AXI_PORT_MONITOR_DEF_COV_VMID_UNSET
  /**
    * Covergroup: trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb47to16
    *
    * This covergroup is cross coverage of snoop DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_hypervisor_type : Captures OS type
    * - acdvm_security_type : Captures Security type
    * - acdvm_addr_mode_bits : Captures addr invalidate modes 
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_tlbinvl_modes_virtaddr_msb47to16 : Crosses coverpoints acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,
    *  acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb47to16;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB47TO32
    
     dvm_snoop_tlbinvl_modes_virtaddr_msb47to16 : cross acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart {
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_IGNORE_TLBINVL_MODES_VIRTADDR
    
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

   /**
    * Covergroup: trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb63to16
    *
    * This covergroup is cross coverage of snoop DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_hypervisor_type : Captures OS type
    * - acdvm_security_type : Captures Security type
    * - acdvm_addr_mode_bits : Captures addr invalidate modes 
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb63to32_firstpart : Captures firstpart of DVM Virtual address MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_tlbinvl_modes_virtaddr_msb63to16 : Crosses coverpoints acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,
    *  acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb63to16;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB63TO32

    dvm_snoop_tlbinvl_modes_virtaddr_msb63to16 : cross acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_IGNORE_TLBINVL_MODES_VIRTADDR
     
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb55to16
    *
    * This covergroup is cross coverage of snoop DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_hypervisor_type : Captures OS type
    * - acdvm_security_type : Captures Security type
    * - acdvm_addr_mode_bits : Captures addr invalidate modes 
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_tlbinvl_modes_virtaddr_msb55to16 : Crosses coverpoints acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,
    *  acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb55to16;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB55TO32

    dvm_snoop_tlbinvl_modes_virtaddr_msb55to16 : cross acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_IGNORE_TLBINVL_MODES_VIRTADDR
     
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb43to16
    *
    * This covergroup is cross coverage of snoop DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_hypervisor_type : Captures OS type
    * - acdvm_security_type : Captures Security type
    * - acdvm_addr_mode_bits : Captures addr invalidate modes 
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb43to32_firstpart : Captures firstpart of DVM Virtual address MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_tlbinvl_modes_virtaddr_msb43to16 : Crosses coverpoints acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,
    *  acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb43to16 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB43TO32

    dvm_snoop_tlbinvl_modes_virtaddr_msb43to16 : cross acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_IGNORE_TLBINVL_MODES_VIRTADDR
     
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb39to16
    *
    * This covergroup is cross coverage ofsnoop DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_hypervisor_type : Captures OS type
    * - acdvm_security_type : Captures Security type
    * - acdvm_addr_mode_bits : Captures addr invalidate modes 
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb39to32_firstpart: Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_tlbinvl_modes_virtaddr_msb39to16 : Crosses coverpoints acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,
    *  acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb39to16 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB39TO32

    dvm_snoop_tlbinvl_modes_virtaddr_msb39to16 : cross acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_IGNORE_TLBINVL_MODES_VIRTADDR
     
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

   /**
    * Covergroup: trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb63to16
    *
    * This covergroup is cross coverage of snoop DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * - snoop_dvm_message_phy_inst_cache_invl_bits : Captures physical instruction cache invalidate by pa etc
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_phy_inst_cache_invl_modes_virtaddr_msb63to16 : Crosses coverpoints acdvm_message_type,snoop_dvm_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb63to16;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB63TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_snoop_phy_inst_cache_invl_modes_virtaddr_msb63to16 : cross acdvm_message_type,snoop_dvm_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
   
    /**
    * Covergroup: trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb55to16
    *
    * This covergroup is cross coverage of snoop DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * - snoop_dvm_message_phy_inst_cache_invl_bits : Captures physical instruction cache invalidate by pa etc
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_phy_inst_cache_invl_modes_virtaddr_msb55to16 : Crosses coverpoints acdvm_message_type,snoop_dvm_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb55to16 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB55TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_snoop_phy_inst_cache_invl_modes_virtaddr_msb55to16 : cross acdvm_message_type,snoop_dvm_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb47to16
    *
    * This covergroup is cross coverage of snoop DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firstpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * - snoop_dvm_message_phy_inst_cache_invl_bits : Captures physical instruction cache invalidate by pa etc
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_phy_inst_cache_invl_modes_virtaddr_msb47to16 : Crosses coverpoints acdvm_message_type,snoop_dvm_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb47to16 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB47TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_snoop_phy_inst_cache_invl_modes_virtaddr_msb47to16 : cross acdvm_message_type,snoop_dvm_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb43to16
    *
    * This covergroup is cross coverage of snoop DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firstpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * - snoop_dvm_message_phy_inst_cache_invl_bits : Captures physical instruction cache invalidate by pa etc
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_phy_inst_cache_invl_modes_virtaddr_msb43to16 : Crosses coverpoints acdvm_message_type,snoop_dvm_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb43to16 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB43TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_snoop_phy_inst_cache_invl_modes_virtaddr_msb43to16 : cross acdvm_message_type,snoop_dvm_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb39to16
    *
    * This covergroup is cross coverage of snoop DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firstpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * - snoop_dvm_message_phy_inst_cache_invl_bits : Captures physical instruction cache invalidate by pa etc
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_phy_inst_cache_invl_modes_virtaddr_msb39to16 : Crosses coverpoints acdvm_message_type,dvm_snoop_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb39to16;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB39TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_snoop_phy_inst_cache_invl_modes_virtaddr_msb39to16 : cross acdvm_message_type,snoop_dvm_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb63to16
    *
    * This covergroup is cross coverage of snoop DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firstpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * - snoop_dvm_message_virt_inst_cache_invl_bits: Captures virtual instruction cache invalidate by pa etc
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_virt_inst_cache_invl_modes_virtaddr_msb63to16 : Crosses coverpoints acdvm_message_type,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb63to16;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB63TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS
    dvm_snoop_virt_inst_cache_invl_modes_virtaddr_msb63to16 : cross acdvm_message_type,snoop_dvm_message_virt_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb55to16
    *
    * This covergroup is cross coverage of snoop DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firstpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * - snoop_dvm_message_virt_inst_cache_invl_bits: Captures virtual instruction cache invalidate by pa etc
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_virt_inst_cache_invl_modes_virtaddr_msb55to16 : Crosses coverpoints acdvm_message_type,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb55to16 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB55TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS
    dvm_snoop_virt_inst_cache_invl_modes_virtaddr_msb55to16 : cross acdvm_message_type,snoop_dvm_message_virt_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb47to16
    *
    * This covergroup is cross coverage of snoop DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firstpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * - snoop_dvm_message_virt_inst_cache_invl_bits: Captures virtual instruction cache invalidate by pa etc
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_virt_inst_cache_invl_modes_virtaddr_msb47to16 : Crosses coverpoints acdvm_message_type,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb47to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB47TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS
    dvm_snoop_virt_inst_cache_invl_modes_virtaddr_msb47to16 : cross acdvm_message_type,snoop_dvm_message_virt_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb43to16
    *
    * This covergroup is cross coverage of snoop DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firstpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * - snoop_dvm_message_virt_inst_cache_invl_bits: Captures virtual instruction cache invalidate by pa etc
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_virt_inst_cache_invl_modes_virtaddr_msb43to16 : Crosses coverpoints acdvm_message_type,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb43to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB43TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS
    dvm_snoop_virt_inst_cache_invl_modes_virtaddr_msb43to16 : cross acdvm_message_type,snoop_dvm_message_virt_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb39to16
    *
    * This covergroup is cross coverage of snoop DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firstpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * - snoop_dvm_message_virt_inst_cache_invl_bits: Captures virtual instruction cache invalidate by pa etc
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_snoop_virt_inst_cache_invl_modes_virtaddr_msb39to16 : Crosses coverpoints acdvm_message_type,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb39to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB39TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS
    dvm_snoop_virt_inst_cache_invl_modes_virtaddr_msb39to16 : cross acdvm_message_type,snoop_dvm_message_virt_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_addr_range_msb63to16
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[63:32] and ARADDR[31:16].
    * The total Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_addr_range_msb63to16 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_addr_range_msb63to16;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB63TO32
    
    snoop_dvm_firstpart_addr_range_msb63to16 :cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_addr_range_msb55to16
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[55:32] and ARADDR[31:16].
    * The total Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_addr_range_msb63to16 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_addr_range_msb55to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB55TO32
    
    snoop_dvm_firstpart_addr_range_msb55to16 :cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_addr_range_msb47to16
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[47:32] and ARADDR[31:16].
    * The total Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_addr_range_msb47to16 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_addr_range_msb47to16 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB47TO32
    
    snoop_dvm_firstpart_addr_range_msb47to16 :cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_addr_range_msb43to16
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[43:32] and ARADDR[31:16].
    * The total Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_addr_range_msb43to16 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_addr_range_msb43to16 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB43TO32
    
    snoop_dvm_firstpart_addr_range_msb43to16 :cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_addr_range_msb39to16
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[39:32] and ARADDR[31:16].
    * The total Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_addr_range_msb39to16 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_addr_range_msb39to16 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB39TO32
    
    snoop_dvm_firstpart_addr_range_msb39to16 :cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_64
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[63:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[63:4]
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * - acaddr_dvm_secondpart_64 : Captures SecondPart of DVM of width64
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_secondpart_addr_range_64 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb63to32_firstpart2,acaddr_dvm_secondpart_64.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_64  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB63TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_SECONDPART_64
    
    snoop_dvm_firstpart_secondpart_addr_range_64: cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart,acaddr_dvm_secondpart_64 {
      
     ignore_bins   ignore_bins_dvm_acaddr_firstpart_range_3_dvm_acaddr_secondpart_range_2 = binsof(acaddr_dvm_msb63to32_firstpart.dvm_acaddr_firstpart_range_3) && binsof(acaddr_dvm_secondpart_64.dvm_acaddr_secondpart_range_2);
     ignore_bins   ignore_bins_dvm_acaddr_firstpart_range_3_dvm_acaddr_secondpart_range_1 = binsof(acaddr_dvm_msb63to32_firstpart.dvm_acaddr_firstpart_range_3) && binsof(acaddr_dvm_secondpart_64.dvm_acaddr_secondpart_range_1);
     ignore_bins   ignore_bins_dvm_acaddr_firstpart_range_2_dvm_acaddr_secondpart_range_4 = binsof(acaddr_dvm_msb63to32_firstpart.dvm_acaddr_firstpart_range_2) && binsof(acaddr_dvm_secondpart_64.dvm_acaddr_secondpart_range_4);   
     ignore_bins   ignore_bins_dvm_acaddr_firstpart_range_1_dvm_acaddr_secondpart_range_4 = binsof(acaddr_dvm_msb63to32_firstpart.dvm_acaddr_firstpart_range_1) && binsof(acaddr_dvm_secondpart_64.dvm_acaddr_secondpart_range_4);   
     ignore_bins   ignore_bins_dvm_acaddr_firstpart_range_1_dvm_acaddr_secondpart_range_3 = binsof(acaddr_dvm_msb63to32_firstpart.dvm_acaddr_firstpart_range_1) && binsof(acaddr_dvm_secondpart_64.dvm_acaddr_secondpart_range_3);   
     ignore_bins   ignore_bins_dvm_acaddr_firstpart_range_1_dvm_acaddr_secondpart_range_2 = binsof(acaddr_dvm_msb63to32_firstpart.dvm_acaddr_firstpart_range_1) && binsof(acaddr_dvm_secondpart_64.dvm_acaddr_secondpart_range_2);   
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

   /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_56
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[55:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[55:4]
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * - acaddr_dvm_secondpart_56 : Captures SecondPart of DVM of width56
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_secondpart_addr_range_56 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb55to32_firstpart,acaddr_dvm_secondpart_56.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_56  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB55TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_SECONDPART_56
    
    snoop_dvm_firstpart_secondpart_addr_range_56: cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart,acaddr_dvm_secondpart_56 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_48
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[47:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[47:4]
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * - acaddr_dvm_secondpart_48 : Captures SecondPart of DVM of width48
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_secondpart_addr_range_48 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart,acaddr_dvm_secondpart_48.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_48  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB47TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_SECONDPART_48
    
    snoop_dvm_firstpart_secondpart_addr_range_48: cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart,acaddr_dvm_secondpart_48 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup


    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_44
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[43:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[43:4]
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * - acaddr_dvm_secondpart_44 : Captures SecondPart of DVM of width44
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_secondpart_addr_range_44 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart,acaddr_dvm_secondpart_44.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_44  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB43TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_SECONDPART_44
    
    snoop_dvm_firstpart_secondpart_addr_range_44: cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart,acaddr_dvm_secondpart_44 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_40
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[39:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[39:4]
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * - acaddr_dvm_secondpart_40 : Captures SecondPart of DVM of width40
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_secondpart_addr_range_40 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart_acaddr_dvm_secondpart_40.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_40  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB39TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_SECONDPART_40
    
    snoop_dvm_firstpart_secondpart_addr_range_40: cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart,acaddr_dvm_secondpart_40 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

`else

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb63to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_hypervisor_type : Captures OS type
    * - acdvm_security_type : Captures Security type
    * - acdvm_addr_mode_bits : Captures addr invalidate modes 
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb63to32_firstpart : Captures firstpart of DVM Virtual address MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_tlbinvl_modes_virtaddr_msb63to16 : Crosses coverpoints acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,
    *  acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb63to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB63TO32
    
     snoop_dvm_tlbinvl_modes_virtaddr_msb63to16 : cross acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart {
   
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_IGNORE_TLBINVL_MODES_VIRTADDR

    option.weight=1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb55to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_hypervisor_type : Captures OS type
    * - acdvm_security_type : Captures Security type
    * - acdvm_addr_mode_bits : Captures addr invalidate modes 
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_tlbinvl_modes_virtaddr_msb55to16 : Crosses coverpoints acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,
    *  acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb55to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB55TO32
    
     snoop_dvm_tlbinvl_modes_virtaddr_msb55to16 : cross acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart {
       `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_IGNORE_TLBINVL_MODES_VIRTADDR
       option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
 
    /**
    * Covergroup: trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb47to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_hypervisor_type : Captures OS type
    * - acdvm_security_type : Captures Security type
    * - acdvm_addr_mode_bits : Captures addr invalidate modes 
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_tlbinvl_modes_virtaddr_msb47to16 : Crosses coverpoints acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,
    *  acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb47to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB47TO32
    
     snoop_dvm_tlbinvl_modes_virtaddr_msb47to16 : cross acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart {
       `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_IGNORE_TLBINVL_MODES_VIRTADDR
       option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb43to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_hypervisor_type : Captures OS type
    * - acdvm_security_type : Captures Security type
    * - acdvm_addr_mode_bits : Captures addr invalidate modes 
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_tlbinvl_modes_virtaddr_msb43to16 : Crosses coverpoints acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,
    *  acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb43to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB43TO32
    
     snoop_dvm_tlbinvl_modes_virtaddr_msb43to16 : cross acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart {
       `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_IGNORE_TLBINVL_MODES_VIRTADDR
       option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb39to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_hypervisor_type : Captures OS type
    * - acdvm_security_type : Captures Security type
    * - acdvm_addr_mode_bits : Captures addr invalidate modes 
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_tlbinvl_modes_virtaddr_msb39to16 : Crosses coverpoints acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,
    *  acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_tlbinvl_modes_virtaddr_msb39to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB39TO32
    
     snoop_dvm_tlbinvl_modes_virtaddr_msb39to16 : cross acdvm_message_type,acdvm_hypervisor_type,acdvm_security_type,acdvm_addr_mode_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart {
       `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_IGNORE_TLBINVL_MODES_VIRTADDR
       option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_branch_predictor_invl_modes_virtaddr_msb43to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_branch_predictor_modes_virtaddr_msb43to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_branch_predictor_invl_modes_virtaddr_msb43to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB43TO32
    
     snoop_dvm_branch_predictor_modes_virtaddr_msb43to16 : cross acdvm_message_type,acdvm_va,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_branch_predictor_invl_modes_virtaddr_msb63to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_branch_predictor_modes_virtaddr_msb63to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_branch_predictor_invl_modes_virtaddr_msb63to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB63TO32
    
     snoop_dvm_branch_predictor_modes_virtaddr_msb63to16 : cross acdvm_message_type,acdvm_va,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_branch_predictor_invl_modes_virtaddr_msb55to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_branch_predictor_modes_virtaddr_msb55to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_branch_predictor_invl_modes_virtaddr_msb55to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB55TO32
    
     snoop_dvm_branch_predictor_modes_virtaddr_msb55to16 : cross acdvm_message_type,acdvm_va,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_branch_predictor_invl_modes_virtaddr_msb47to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_branch_predictor_modes_virtaddr_msb47to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_branch_predictor_invl_modes_virtaddr_msb47to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB47TO32
    
     snoop_dvm_branch_predictor_modes_virtaddr_msb47to16 : cross acdvm_message_type,acdvm_va,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_branch_predictor_invl_modes_virtaddr_msb39to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_branch_predictor_modes_virtaddr_msb47to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_branch_predictor_invl_modes_virtaddr_msb39to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB39TO32
    
     snoop_dvm_branch_predictor_modes_virtaddr_msb39to16 : cross acdvm_message_type,acdvm_va,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb63to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_security_type : Captures Security Type
    * - acdvm_virtindex : Captures Virtual Index
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb63to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acdvm_security_type,acdvm_virtindex,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb63to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB63TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb63to16 : cross acdvm_message_type,snoop_dvm_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb55to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_security_type : Captures Security Type
    * - acdvm_virtindex : Captures Virtual Index
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb55to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acdvm_security_type,acdvm_virtindex,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb55to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB55TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb55to16 : cross acdvm_message_type,snoop_dvm_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb47to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_security_type : Captures Security Type
    * - acdvm_virtindex : Captures Virtual Index
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb47to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acdvm_security_type,acdvm_virtindex,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb47to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB47TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb47to16 : cross acdvm_message_type,snoop_dvm_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb43to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_security_type : Captures Security Type
    * - acdvm_virtindex : Captures Virtual Index
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb43to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acdvm_security_type,acdvm_virtindex,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb43to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB43TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb43to16 : cross acdvm_message_type,snoop_dvm_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb39to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_security_type : Captures Security Type
    * - acdvm_virtindex : Captures Virtual Index
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb39to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acdvm_security_type,acdvm_virtindex,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb39to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB39TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    snoop_dvm_phy_inst_cache_invl_modes_virtaddr_msb39to16 : cross acdvm_message_type,snoop_dvm_message_phy_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb63to16
    *
    * This covergroup is cross coverage of snoop DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_security_type : Captures Security Type
    * - acdvm_hypervisor_type : Captures OS TYPE
    * - acdvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb63to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acdvm_security_type,acdvm_hypervisor_type,acdvm_vmid_asid_or_virtindex,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb63to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB63TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS
    snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb63to16 : cross acdvm_message_type,snoop_dvm_message_virt_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb55to16
    *
    * This covergroup is cross coverage of snoop DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_security_type : Captures Security Type
    * - acdvm_hypervisor_type : Captures OS TYPE
    * - acdvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb55to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acdvm_security_type,acdvm_hypervisor_type,acdvm_vmid_asid_or_virtindex,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb55to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB55TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS
    snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb55to16 : cross acdvm_message_type,snoop_dvm_message_virt_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb47to16
    *
    * This covergroup is cross coverage of snoop DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_security_type : Captures Security Type
    * - acdvm_hypervisor_type : Captures OS TYPE
    * - acdvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb47to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acdvm_security_type,acdvm_hypervisor_type,acdvm_vmid_asid_or_virtindex,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb47to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB47TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS
    snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb47to16 : cross acdvm_message_type,snoop_dvm_message_virt_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb43to16
    *
    * This covergroup is cross coverage of snoop DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_security_type : Captures Security Type
    * - acdvm_hypervisor_type : Captures OS TYPE
    * - acdvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb43to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acdvm_security_type,acdvm_hypervisor_type,acdvm_vmid_asid_or_virtindex,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb43to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB43TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS
    snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb43to16 : cross acdvm_message_type,snoop_dvm_message_virt_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb39to16
    *
    * This covergroup is cross coverage of snoop DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - acdvm_message_type: Captures DVM Message Type
    * - acdvm_security_type : Captures Security Type
    * - acdvm_hypervisor_type : Captures OS TYPE
    * - acdvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - acdvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb39to16 : Crosses coverpoints acdvm_message_type,acdvm_va,acdvm_security_type,acdvm_hypervisor_type,acdvm_vmid_asid_or_virtindex,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb39to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB39TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS
    snoop_dvm_virt_inst_cache_invl_modes_virtaddr_msb39to16 : cross acdvm_message_type,snoop_dvm_message_virt_inst_cache_invl_bits,acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_addr_range_msb63to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[63:32] and ARADDR[31:16].
    * The total Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firstpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_addr_range_msb63to16 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_addr_range_msb63to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB63TO32
    
    snoop_dvm_firstpart_addr_range_msb63to16 :cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_addr_range_msb55to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[55:32] and ARADDR[31:16].
    * The total Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firstpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_addr_range_msb55to16 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_addr_range_msb55to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB55TO32
    
    snoop_dvm_firstpart_addr_range_msb55to16 :cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

     /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_addr_range_msb47to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[47:32] and ARADDR[31:16].
    * The total Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firstpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_addr_range_msb47to16 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_addr_range_msb47to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB47TO32
    
    snoop_dvm_firstpart_addr_range_msb47to16 :cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

   /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_addr_range_msb43to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[43:32] and ARADDR[31:16].
    * The total Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firstpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_addr_range_msb43to16 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_addr_range_msb43to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB43TO32
    
    snoop_dvm_firstpart_addr_range_msb43to16 :cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_addr_range_msb39to16_vmid_unset
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[39:32] and ARADDR[31:16].
    * The total Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firstpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_addr_range_msb39to16 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_addr_range_msb39to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB39TO32
    
    snoop_dvm_firstpart_addr_range_msb39to16 :cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_64_vmid_unset
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[63:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[63:4]
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * - acaddr_dvm_secondpart_64 : Captures SecondPart of DVM of width64
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_secondpart_addr_range_64 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firsrpart_va_or_asid,acaddr_dvm_msb63to32_firstpart2,acaddr_dvm_secondpart_64.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_64_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB63TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_SECONDPART_64
    
    snoop_dvm_firstpart_secondpart_addr_range_64: cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb63to32_firstpart,acaddr_dvm_secondpart_64 {
      
     ignore_bins   ignore_bins_dvm_acaddr_firstpart_range_3_dvm_acaddr_secondpart_range_2 = binsof(acaddr_dvm_msb63to32_firstpart.dvm_acaddr_firstpart_range_3) && binsof(acaddr_dvm_secondpart_64.dvm_acaddr_secondpart_range_2);
     ignore_bins   ignore_bins_dvm_acaddr_firstpart_range_3_dvm_acaddr_secondpart_range_1 = binsof(acaddr_dvm_msb63to32_firstpart.dvm_acaddr_firstpart_range_3) && binsof(acaddr_dvm_secondpart_64.dvm_acaddr_secondpart_range_1);
     ignore_bins   ignore_bins_dvm_acaddr_firstpart_range_2_dvm_acaddr_secondpart_range_4 = binsof(acaddr_dvm_msb63to32_firstpart.dvm_acaddr_firstpart_range_2) && binsof(acaddr_dvm_secondpart_64.dvm_acaddr_secondpart_range_4);   
     ignore_bins   ignore_bins_dvm_acaddr_firstpart_range_1_dvm_acaddr_secondpart_range_4 = binsof(acaddr_dvm_msb63to32_firstpart.dvm_acaddr_firstpart_range_1) && binsof(acaddr_dvm_secondpart_64.dvm_acaddr_secondpart_range_4);   
     ignore_bins   ignore_bins_dvm_acaddr_firstpart_range_1_dvm_acaddr_secondpart_range_3 = binsof(acaddr_dvm_msb63to32_firstpart.dvm_acaddr_firstpart_range_1) && binsof(acaddr_dvm_secondpart_64.dvm_acaddr_secondpart_range_3);   
     ignore_bins   ignore_bins_dvm_acaddr_firstpart_range_1_dvm_acaddr_secondpart_range_2 = binsof(acaddr_dvm_msb63to32_firstpart.dvm_acaddr_firstpart_range_1) && binsof(acaddr_dvm_secondpart_64.dvm_acaddr_secondpart_range_2);   
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_56_vmid_unset
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[55:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[55:4]
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * - acaddr_dvm_secondpart_56 : Captures SecondPart of DVM of width56
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_secondpart_addr_range_56 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart,acaddr_dvm_secondpart_56.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_56_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB55TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_SECONDPART_56
    
    snoop_dvm_firstpart_secondpart_addr_range_56: cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb55to32_firstpart,acaddr_dvm_secondpart_56 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_48_vmid_unset
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[47:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[47:4]
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * - acaddr_dvm_secondpart_48 : Captures SecondPart of DVM of width48
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_secondpart_addr_range_48 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart,acaddr_dvm_secondpart_48.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_48_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB47TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_SECONDPART_48
    
    snoop_dvm_firstpart_secondpart_addr_range_48: cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb47to32_firstpart,acaddr_dvm_secondpart_48 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_44_vmid_unset
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[43:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[43:4]
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * - acaddr_dvm_secondpart_44 : Captures SecondPart of DVM of width44
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_secondpart_addr_range_44 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart,acaddr_dvm_secondpart_44.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_44_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB43TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_SECONDPART_44
    
    snoop_dvm_firstpart_secondpart_addr_range_44: cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb43to32_firstpart,acaddr_dvm_secondpart_44 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_40_vmid_unset
    *
    * This covergroup is cross coverage of snoop FirstPart of DVM (Virtual Address) on ARADDR[39:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[39:4]
    *
    * Coverpoints:
    *
    * - acaddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - acaddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - acaddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * - acaddr_dvm_secondpart_40 : Captures SecondPart of DVM of width40
    * .
    *
    * Cross coverpoints:
    *
    * -snoop_dvm_firstpart_secondpart_addr_range_40 : Crosses coverpoints acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart,acaddr_dvm_secondpart_40.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_snoop_dvm_firstpart_secondpart_addr_range_40_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_FIRSTPART_MSB39TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_ARADDR_SECONDPART_40
    
    snoop_dvm_firstpart_secondpart_addr_range_40: cross acaddr_dvm_firstpart_va_or_vmid,acaddr_dvm_firstpart_va_or_asid,acaddr_dvm_msb39to32_firstpart,acaddr_dvm_secondpart_40 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
`endif 

`ifndef SVT_AXI_PORT_MONITOR_DEF_COV_VMID_UNSET
 
  // Added in 2.43a
    
    /**
    * Covergroup: trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb63to16
    *
    * This covergroup is cross coverage of DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_hypervisor_type : Captures OS type
    * - ardvm_security_type : Captures Security type
    * - ardvm_addr_mode_bits : Captures addr invalidate modes 
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb63to32_firstpart : Captures firstpart of DVM Virtual address MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_tlbinvl_modes_virtaddr_msb63to16 : Crosses coverpoints ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,
    *  ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb63to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB63TO32
    
     dvm_tlbinvl_modes_virtaddr_msb63to16 : cross ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart {
   `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_IGNORE_TLBINVL_MODES_VIRTADDR 
    option.weight=1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb55to16
    *
    * This covergroup is cross coverage of DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_hypervisor_type : Captures OS type
    * - ardvm_security_type : Captures Security type
    * - ardvm_addr_mode_bits : Captures addr invalidate modes 
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_tlbinvl_modes_virtaddr_msb55to16 : Crosses coverpoints ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,
    *  ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb55to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB55TO32
    
     dvm_tlbinvl_modes_virtaddr_msb55to16 : cross ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart {
       `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_IGNORE_TLBINVL_MODES_VIRTADDR
       option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
  
    /**
    * Covergroup: trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb47to16
    *
    * This covergroup is cross coverage of DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_hypervisor_type : Captures OS type
    * - ardvm_security_type : Captures Security type
    * - ardvm_addr_mode_bits : Captures addr invalidate modes 
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_tlbinvl_modes_virtaddr_msb47to16 : Crosses coverpoints ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,
    *  ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb47to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB47TO32
    
     dvm_tlbinvl_modes_virtaddr_msb47to16 : cross ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart {
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_IGNORE_TLBINVL_MODES_VIRTADDR
     option.weight = 1;
    }
    option.per_instance = 1;
    endgroup


    /**
    * Covergroup: trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb43to16
    *
    * This covergroup is cross coverage of DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_hypervisor_type : Captures OS type
    * - ardvm_security_type : Captures Security type
    * - ardvm_addr_mode_bits : Captures addr invalidate modes 
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb43to32_firstpart : Captures firstpart of DVM Virtual address MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_tlbinvl_modes_virtaddr_msb43to16 : Crosses coverpoints ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,
    *  ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb43to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB43TO32
    
     dvm_tlbinvl_modes_virtaddr_msb43to16 : cross ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart {  
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_IGNORE_TLBINVL_MODES_VIRTADDR  
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
   
   /**
    * Covergroup: trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb39to16
    *
    * This covergroup is cross coverage of DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_hypervisor_type : Captures OS type
    * - ardvm_security_type : Captures Security type
    * - ardvm_addr_mode_bits : Captures addr invalidate modes 
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb39to32_firstpart: Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_tlbinvl_modes_virtaddr_msb39to16 : Crosses coverpoints ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,
    *  ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb39to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB39TO32
    
     dvm_tlbinvl_modes_virtaddr_msb39to16 : cross ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_IGNORE_TLBINVL_MODES_VIRTADDR
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb43to16
    *
    * This covergroup is cross coverage of DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_branch_predictor_modes_virtaddr_msb43to16 : Crosses coverpoints ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb43to16   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB43TO32
    
     dvm_branch_predictor_modes_virtaddr_msb43to16 : cross ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb63to16
    *
    * This covergroup is cross coverage of DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_branch_predictor_modes_virtaddr_msb63to16 : Crosses coverpoints ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb63to16   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB63TO32
    
     dvm_branch_predictor_modes_virtaddr_msb63to16 : cross ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb55to16
    *
    * This covergroup is cross coverage of DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_branch_predictor_modes_virtaddr_msb55to16 : Crosses coverpoints ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb55to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB55TO32
    
     dvm_branch_predictor_modes_virtaddr_msb55to16 : cross ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb47to16
    *
    * This covergroup is cross coverage of DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_branch_predictor_modes_virtaddr_msb47to16 : Crosses coverpoints ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb47to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB47TO32
    
     dvm_branch_predictor_modes_virtaddr_msb47to16 : cross ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb39to16
    *
    * This covergroup is cross coverage of DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_branch_predictor_modes_virtaddr_msb39to16 : Crosses coverpoints ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb39to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB39TO32
    
     dvm_branch_predictor_modes_virtaddr_msb39to16 : cross ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb63to16
    *
    * This covergroup is cross coverage of DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_virtindex : Captures Virtual Index
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_phy_inst_cache_invl_modes_virtaddr_msb63to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb63to16 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB63TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_phy_inst_cache_invl_modes_virtaddr_msb63to16 : cross ardvm_message_type,dvm_message_phy_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb55to16
    *
    * This covergroup is cross coverage of DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_virtindex : Captures Virtual Index
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_phy_inst_cache_invl_modes_virtaddr_msb55to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb55to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB55TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_phy_inst_cache_invl_modes_virtaddr_msb55to16 : cross ardvm_message_type,dvm_message_phy_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb47to16
    *
    * This covergroup is cross coverage of DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_virtindex : Captures Virtual Index
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_phy_inst_cache_invl_modes_virtaddr_msb47to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb47to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB47TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_phy_inst_cache_invl_modes_virtaddr_msb47to16 : cross ardvm_message_type,dvm_message_phy_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb43to16
    *
    * This covergroup is cross coverage of DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - dvm_message_phy_inst_cache_invl_bits : Captures types of physical instruction cache invalidation
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_phy_inst_cache_invl_modes_virtaddr_msb43to16 : Crosses coverpoints ardvm_message_type,dvm_message_phy_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb43to16 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB43TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_phy_inst_cache_invl_modes_virtaddr_msb43to16 : cross ardvm_message_type,dvm_message_phy_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb39to16
    *
    * This covergroup is cross coverage of DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_virtindex : Captures Virtual Index
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msbto3932_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_phy_inst_cache_invl_modes_virtaddr_msb39to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb39to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB39TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_phy_inst_cache_invl_modes_virtaddr_msb39to16 : cross ardvm_message_type,dvm_message_phy_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

   /**
    * Covergroup: trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb63to16
    *
    * This covergroup is cross coverage of DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_hypervisor_type : Captures OS TYPE
    * - ardvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_virt_inst_cache_invl_modes_virtaddr_msb63to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_hypervisor_type,ardvm_vmid_asid_or_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb63to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB63TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS
    dvm_virt_inst_cache_invl_modes_virtaddr_msb63to16 : cross ardvm_message_type,dvm_message_virt_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb55to16
    *
    * This covergroup is cross coverage of DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_hypervisor_type : Captures OS TYPE
    * - ardvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_virt_inst_cache_invl_modes_virtaddr_msb55to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_hypervisor_type,ardvm_vmid_asid_or_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb55to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB55TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS

    dvm_virt_inst_cache_invl_modes_virtaddr_msb55to16 : cross ardvm_message_type,dvm_message_virt_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb47to16
    *
    * This covergroup is cross coverage of DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_hypervisor_type : Captures OS TYPE
    * - ardvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_virt_inst_cache_invl_modes_virtaddr_msb47to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_hypervisor_type,ardvm_vmid_asid_or_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb47to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB47TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS


    dvm_virt_inst_cache_invl_modes_virtaddr_msb47to16 : cross ardvm_message_type,dvm_message_virt_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart {
   
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb43to16
    *
    * This covergroup is cross coverage of DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_hypervisor_type : Captures OS TYPE
    * - ardvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_virt_inst_cache_invl_modes_virtaddr_msb43to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_hypervisor_type,ardvm_vmid_asid_or_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb43to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB43TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS

    dvm_virt_inst_cache_invl_modes_virtaddr_msb43to16 : cross ardvm_message_type,dvm_message_virt_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart {
     option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
   
    /**
    * Covergroup: trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb39to16
    *
    * This covergroup is cross coverage of DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_hypervisor_type : Captures OS TYPE
    * - ardvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_virt_inst_cache_invl_modes_virtaddr_msb39to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_hypervisor_type,ardvm_vmid_asid_or_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb39to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB39TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS
    
     dvm_virt_inst_cache_invl_modes_virtaddr_msb39to16 : cross ardvm_message_type,dvm_message_virt_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart {
     option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_addr_range_msb63to16
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[63:32] and ARADDR[31:16].
    * The total Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_addr_range_msb63to16 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_addr_range_msb63to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB63TO32
    
    dvm_firstpart_addr_range_msb63to16 :cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_addr_range_msb55to16
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[55:32] and ARADDR[31:16].
    * The total Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_addr_range_msb55to16 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_addr_range_msb55to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB55TO32
    
    dvm_firstpart_addr_range_msb55to16 : cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_addr_range_msb47to16
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[47:32] and ARADDR[31:16].
    * The total Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_addr_range_msb47to16 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_addr_range_msb47to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB47TO32
    
    dvm_firstpart_addr_range_msb47to16 : cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
   
    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_addr_range_msb43to16
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[43:32] and ARADDR[31:16].
    * The total Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_addr_range_msb43to16 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_addr_range_msb43to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB43TO32
    
    dvm_firstpart_addr_range_msb43to16 :cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_addr_range_msb39to16
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[39:32] and ARADDR[31:16].
    * The total Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_addr_range_msb39to16 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_addr_range_msb39to16  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB39TO32
    
    dvm_firstpart_addr_range_msb39to16 : cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_secondpart_addr_range_64
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[63:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[63:4]
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * - araddr_dvm_secondpart_64 : Captures SecondPart of DVM of width64
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_secondpart_addr_range_64 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart2,araddr_dvm_secondpart_64.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_secondpart_addr_range_64  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB63TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_SECONDPART_64
    
    dvm_firstpart_secondpart_addr_range_64: cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart,araddr_dvm_secondpart_64 {
      
     ignore_bins   ignore_bins_dvm_araddr_firstpart_range_3_dvm_araddr_secondpart_range_2 = binsof(araddr_dvm_msb63to32_firstpart.dvm_araddr_firstpart_range_3) && binsof(araddr_dvm_secondpart_64.dvm_araddr_secondpart_range_2);
     ignore_bins   ignore_bins_dvm_araddr_firstpart_range_3_dvm_araddr_secondpart_range_1 = binsof(araddr_dvm_msb63to32_firstpart.dvm_araddr_firstpart_range_3) && binsof(araddr_dvm_secondpart_64.dvm_araddr_secondpart_range_1);
     ignore_bins   ignore_bins_dvm_araddr_firstpart_range_2_dvm_araddr_secondpart_range_4 = binsof(araddr_dvm_msb63to32_firstpart.dvm_araddr_firstpart_range_2) && binsof(araddr_dvm_secondpart_64.dvm_araddr_secondpart_range_4);   
     ignore_bins   ignore_bins_dvm_araddr_firstpart_range_1_dvm_araddr_secondpart_range_4 = binsof(araddr_dvm_msb63to32_firstpart.dvm_araddr_firstpart_range_1) && binsof(araddr_dvm_secondpart_64.dvm_araddr_secondpart_range_4);   
     ignore_bins   ignore_bins_dvm_araddr_firstpart_range_1_dvm_araddr_secondpart_range_3 = binsof(araddr_dvm_msb63to32_firstpart.dvm_araddr_firstpart_range_1) && binsof(araddr_dvm_secondpart_64.dvm_araddr_secondpart_range_3);   
     ignore_bins   ignore_bins_dvm_araddr_firstpart_range_1_dvm_araddr_secondpart_range_2 = binsof(araddr_dvm_msb63to32_firstpart.dvm_araddr_firstpart_range_1) && binsof(araddr_dvm_secondpart_64.dvm_araddr_secondpart_range_2);   
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_secondpart_addr_range_56
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[55:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[55:4]
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * - araddr_dvm_secondpart_56 : Captures SecondPart of DVM of width56
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_secondpart_addr_range_56 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart,araddr_dvm_secondpart_56.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_secondpart_addr_range_56  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB55TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_SECONDPART_56
    
    dvm_firstpart_secondpart_addr_range_56: cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart,araddr_dvm_secondpart_56 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_secondpart_addr_range_48
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[47:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[47:4]
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * - araddr_dvm_secondpart_48 : Captures SecondPart of DVM of width48
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_secondpart_addr_range_48 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart,araddr_dvm_secondpart_48.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_secondpart_addr_range_48  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB47TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_SECONDPART_48
    
    dvm_firstpart_secondpart_addr_range_48: cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart,araddr_dvm_secondpart_48 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_secondpart_addr_range_44
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[43:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[43:4]
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * - araddr_dvm_secondpart_44 : Captures SecondPart of DVM of width44
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_secondpart_addr_range_44 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart,araddr_dvm_secondpart_44.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_secondpart_addr_range_44  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB43TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_SECONDPART_44
    
    dvm_firstpart_secondpart_addr_range_44: cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart,araddr_dvm_secondpart_44 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_secondpart_addr_range_40
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[39:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[39:4]
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * - araddr_dvm_secondpart_40 : Captures SecondPart of DVM of width40
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_secondpart_addr_range_40 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart_araddr_dvm_secondpart_40.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_secondpart_addr_range_40  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB39TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_SECONDPART_40
    
    dvm_firstpart_secondpart_addr_range_40: cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart,araddr_dvm_secondpart_40 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
   
    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_secondpart_addr_range_32
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[39:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[39:4]
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_secondpart_40 : Captures SecondPart of DVM of width40
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_secondpart_addr_range_32 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_secondpart_32.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_secondpart_addr_range_32  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_SECONDPART_32
    
    dvm_firstpart_secondpart_addr_range_32: cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_secondpart_32 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
`else
  // Added in 2.43a
    
    /**
    * Covergroup: trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb63to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_hypervisor_type : Captures OS type
    * - ardvm_security_type : Captures Security type
    * - ardvm_addr_mode_bits : Captures addr invalidate modes 
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb63to32_firstpart : Captures firstpart of DVM Virtual address MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_tlbinvl_modes_virtaddr_msb63to16 : Crosses coverpoints ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,
    *  ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb63to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB63TO32
    
     dvm_tlbinvl_modes_virtaddr_msb63to16 : cross ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart {
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_IGNORE_TLBINVL_MODES_VIRTADDR 
    option.weight=1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb55to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_hypervisor_type : Captures OS type
    * - ardvm_security_type : Captures Security type
    * - ardvm_addr_mode_bits : Captures addr invalidate modes 
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_tlbinvl_modes_virtaddr_msb55to16 : Crosses coverpoints ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,
    *  ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb55to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB55TO32
    
     dvm_tlbinvl_modes_virtaddr_msb55to16 : cross ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart {
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_IGNORE_TLBINVL_MODES_VIRTADDR
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
  
    /**
    * Covergroup: trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb47to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_hypervisor_type : Captures OS type
    * - ardvm_security_type : Captures Security type
    * - ardvm_addr_mode_bits : Captures addr invalidate modes 
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_tlbinvl_modes_virtaddr_msb47to16 : Crosses coverpoints ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,
    *  ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb47to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB47TO32
    
     dvm_tlbinvl_modes_virtaddr_msb47to16 : cross ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart {
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_IGNORE_TLBINVL_MODES_VIRTADDR 
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

   
    /**
    * Covergroup: trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb43to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_hypervisor_type : Captures OS type
    * - ardvm_security_type : Captures Security type
    * - ardvm_addr_mode_bits : Captures addr invalidate modes 
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb43to32_firstpart : Captures firstpart of DVM Virtual address MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_tlbinvl_modes_virtaddr_msb43to16 : Crosses coverpoints ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,
    *  ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb43to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB43TO32
    
     dvm_tlbinvl_modes_virtaddr_msb43to16 : cross ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart {
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_IGNORE_TLBINVL_MODES_VIRTADDR 
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
   
   /**
    * Covergroup: trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb39to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM TLB Invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_hypervisor_type : Captures OS type
    * - ardvm_security_type : Captures Security type
    * - ardvm_addr_mode_bits : Captures addr invalidate modes 
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb39to32_firstpart: Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_tlbinvl_modes_virtaddr_msb39to16 : Crosses coverpoints ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,
    *  ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_tlbinvl_modes_virtaddr_msb39to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_TLB_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_HYPERVISOR_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_SECURITY_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ADDR_MODE_BITS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB39TO32
    
     dvm_tlbinvl_modes_virtaddr_msb39to16 : cross ardvm_message_type,ardvm_hypervisor_type,ardvm_security_type,ardvm_addr_mode_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart {
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_IGNORE_TLBINVL_MODES_VIRTADDR
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb43to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_branch_predictor_modes_virtaddr_msb43to16 : Crosses coverpoints ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb43to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB43TO32
    
     dvm_branch_predictor_modes_virtaddr_msb43to16 : cross ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb63to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_branch_predictor_modes_virtaddr_msb63to16 : Crosses coverpoints ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb63to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB63TO32
    
     dvm_branch_predictor_modes_virtaddr_msb63to16 : cross ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb55to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_branch_predictor_modes_virtaddr_msb55to16 : Crosses coverpoints ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb55to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB55TO32
    
     dvm_branch_predictor_modes_virtaddr_msb55to16 : cross ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb47to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_branch_predictor_modes_virtaddr_msb47to16 : Crosses coverpoints ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb47to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB47TO32
    
     dvm_branch_predictor_modes_virtaddr_msb47to16 : cross ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb39to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM Branch Predictor invalidate message type,invalidate address modes and virtual address range
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_branch_predictor_modes_virtaddr_msb39to16 : Crosses coverpoints ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_msb39to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_BP_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_VA
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB39TO32
    
     dvm_branch_predictor_modes_virtaddr_msb39to16 : cross ardvm_message_type,ardvm_va,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb63to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_virtindex : Captures Virtual Index
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_phy_inst_cache_invl_modes_virtaddr_msb63to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb63to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB63TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_phy_inst_cache_invl_modes_virtaddr_msb63to16 : cross ardvm_message_type,dvm_message_phy_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb55to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_virtindex : Captures Virtual Index
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_phy_inst_cache_invl_modes_virtaddr_msb55to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb55to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB55TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_phy_inst_cache_invl_modes_virtaddr_msb55to16 : cross ardvm_message_type,dvm_message_phy_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb47to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_virtindex : Captures Virtual Index
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_phy_inst_cache_invl_modes_virtaddr_msb47to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb47to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB47TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_phy_inst_cache_invl_modes_virtaddr_msb47to16 : cross ardvm_message_type,dvm_message_phy_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb43to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - dvm_message_phy_inst_cache_invl_bits : Captures types of physical instruction cache invalidation
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_phy_inst_cache_invl_modes_virtaddr_msb43to16 : Crosses coverpoints ardvm_message_type,dvm_message_phy_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb43to16_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB43TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_phy_inst_cache_invl_modes_virtaddr_msb43to16 : cross ardvm_message_type,dvm_message_phy_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb39to16
    *
    * This covergroup is cross coverage of DVM Physical Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_virtindex : Captures Virtual Index
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msbto3932_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_phy_inst_cache_invl_modes_virtaddr_msb39to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_msb39to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_PHY_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB39TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_PHY_INST_CACHE_INVL_BITS
    dvm_phy_inst_cache_invl_modes_virtaddr_msb39to16 : cross ardvm_message_type,dvm_message_phy_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

   /**
    * Covergroup: trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb63to16
    *
    * This covergroup is cross coverage of DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_hypervisor_type : Captures OS TYPE
    * - ardvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_virt_inst_cache_invl_modes_virtaddr_msb63to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_hypervisor_type,ardvm_vmid_asid_or_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb63to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB63TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS
    dvm_virt_inst_cache_invl_modes_virtaddr_msb63to16 : cross ardvm_message_type,dvm_message_virt_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart {
      option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb55to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_hypervisor_type : Captures OS TYPE
    * - ardvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_virt_inst_cache_invl_modes_virtaddr_msb55to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_hypervisor_type,ardvm_vmid_asid_or_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb55to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB55TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS

    dvm_virt_inst_cache_invl_modes_virtaddr_msb55to16 : cross ardvm_message_type,dvm_message_virt_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart {
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb47to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 32 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_hypervisor_type : Captures OS TYPE
    * - ardvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_virt_inst_cache_invl_modes_virtaddr_msb47to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_hypervisor_type,ardvm_vmid_asid_or_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb47to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB47TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS


    dvm_virt_inst_cache_invl_modes_virtaddr_msb47to16 : cross ardvm_message_type,dvm_message_virt_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart {
   
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb43to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_hypervisor_type : Captures OS TYPE
    * - ardvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_virt_inst_cache_invl_modes_virtaddr_msb43to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_hypervisor_type,ardvm_vmid_asid_or_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb43to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB43TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS

    dvm_virt_inst_cache_invl_modes_virtaddr_msb43to16 : cross ardvm_message_type,dvm_message_virt_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart {
     option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
   
    /**
    * Covergroup: trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb39to16_vmid_unset
    *
    * This covergroup is cross coverage of DVM Virtual Instruction Cache invalidate message type,
    * invalidate address modes and virtual address range.
    * The Virtual address width is 24 bits.
    *
    *
    * Coverpoints:
    *
    * - ardvm_message_type: Captures DVM Message Type
    * - ardvm_security_type : Captures Security Type
    * - ardvm_hypervisor_type : Captures OS TYPE
    * - ardvm_vmid_asid_or_virtindex : Captures VMID and ASID
    * - ardvm_va : Captures ARADDR[0] which implies invalidate by VA or invalidate All
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_virt_inst_cache_invl_modes_virtaddr_msb39to16 : Crosses coverpoints ardvm_message_type,ardvm_va,ardvm_security_type,ardvm_hypervisor_type,ardvm_vmid_asid_or_virtindex,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_msb39to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE_VIR_INST_INVL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB39TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_MESSAGE_VIRT_INST_CACHE_INVL_BITS
    
     dvm_virt_inst_cache_invl_modes_virtaddr_msb39to16 : cross ardvm_message_type,dvm_message_virt_inst_cache_invl_bits,araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart {
     option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_addr_range_msb63to16_vmid_unset
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[63:32] and ARADDR[31:16].
    * The total Virtual address width is 48 bits.
    *
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_addr_range_msb63to16 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_addr_range_msb63to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB63TO32
    
    dvm_firstpart_addr_range_msb63to16 :cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_addr_range_msb55to16_vmid_unset
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[55:32] and ARADDR[31:16].
    * The total Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_addr_range_msb55to16 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_addr_range_msb55to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB55TO32
    
    dvm_firstpart_addr_range_msb55to16 : cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_addr_range_msb47to16_vmid_unset
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[47:32] and ARADDR[31:16].
    * The total Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_addr_range_msb47to16 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_addr_range_msb47to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB47TO32
    
    dvm_firstpart_addr_range_msb47to16 : cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
   
    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_addr_range_msb43to16_vmid_unset
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[43:32] and ARADDR[31:16].
    * The total Virtual address width is 28 bits.
    *
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_addr_range_msb43to16 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_addr_range_msb43to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB43TO32
    
    dvm_firstpart_addr_range_msb43to16 :cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_addr_range_msb39to16_vmid_unset
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[39:32] and ARADDR[31:16].
    * The total Virtual address width is 40 bits.
    *
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_addr_range_msb39to16 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_addr_range_msb39to16_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB39TO32
    
    dvm_firstpart_addr_range_msb39to16 : cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_secondpart_addr_range_64_vmid_unset
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[63:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[63:4]
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb63to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width32
    * - araddr_dvm_secondpart_64 : Captures SecondPart of DVM of width64
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_secondpart_addr_range_64 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart2,araddr_dvm_secondpart_64.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_secondpart_addr_range_64_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB63TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_SECONDPART_64
    
    dvm_firstpart_secondpart_addr_range_64: cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb63to32_firstpart,araddr_dvm_secondpart_64 {
      
     ignore_bins   ignore_bins_dvm_araddr_firstpart_range_3_dvm_araddr_secondpart_range_2 = binsof(araddr_dvm_msb63to32_firstpart.dvm_araddr_firstpart_range_3) && binsof(araddr_dvm_secondpart_64.dvm_araddr_secondpart_range_2);
     ignore_bins   ignore_bins_dvm_araddr_firstpart_range_3_dvm_araddr_secondpart_range_1 = binsof(araddr_dvm_msb63to32_firstpart.dvm_araddr_firstpart_range_3) && binsof(araddr_dvm_secondpart_64.dvm_araddr_secondpart_range_1);
     ignore_bins   ignore_bins_dvm_araddr_firstpart_range_2_dvm_araddr_secondpart_range_4 = binsof(araddr_dvm_msb63to32_firstpart.dvm_araddr_firstpart_range_2) && binsof(araddr_dvm_secondpart_64.dvm_araddr_secondpart_range_4);   
     ignore_bins   ignore_bins_dvm_araddr_firstpart_range_1_dvm_araddr_secondpart_range_4 = binsof(araddr_dvm_msb63to32_firstpart.dvm_araddr_firstpart_range_1) && binsof(araddr_dvm_secondpart_64.dvm_araddr_secondpart_range_4);   
     ignore_bins   ignore_bins_dvm_araddr_firstpart_range_1_dvm_araddr_secondpart_range_3 = binsof(araddr_dvm_msb63to32_firstpart.dvm_araddr_firstpart_range_1) && binsof(araddr_dvm_secondpart_64.dvm_araddr_secondpart_range_3);   
     ignore_bins   ignore_bins_dvm_araddr_firstpart_range_1_dvm_araddr_secondpart_range_2 = binsof(araddr_dvm_msb63to32_firstpart.dvm_araddr_firstpart_range_1) && binsof(araddr_dvm_secondpart_64.dvm_araddr_secondpart_range_2);   
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_secondpart_addr_range_56_vmid_unset
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[55:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[55:4]
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb55to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width24
    * - araddr_dvm_secondpart_56 : Captures SecondPart of DVM of width56
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_secondpart_addr_range_56 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart,araddr_dvm_secondpart_56.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_secondpart_addr_range_56_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB55TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_SECONDPART_56
    
    dvm_firstpart_secondpart_addr_range_56: cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb55to32_firstpart,araddr_dvm_secondpart_56 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_secondpart_addr_range_48_vmid_unset
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[47:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[47:4]
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb47to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width16
    * - araddr_dvm_secondpart_48 : Captures SecondPart of DVM of width48
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_secondpart_addr_range_48 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart,araddr_dvm_secondpart_48.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_secondpart_addr_range_48_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB47TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_SECONDPART_48
    
    dvm_firstpart_secondpart_addr_range_48: cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb47to32_firstpart,araddr_dvm_secondpart_48 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_secondpart_addr_range_44_vmid_unset
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[43:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[43:4]
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb43to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width12
    * - araddr_dvm_secondpart_44 : Captures SecondPart of DVM of width44
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_secondpart_addr_range_44 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart,araddr_dvm_secondpart_44.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_secondpart_addr_range_44_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB43TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_SECONDPART_44
    
    dvm_firstpart_secondpart_addr_range_44: cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb43to32_firstpart,araddr_dvm_secondpart_44 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
    
    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_secondpart_addr_range_40_vmid_unset
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[39:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[39:4]
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_msb39to32_firstpart : Captures firstpart of DVM VA MSB to 32 of width8
    * - araddr_dvm_secondpart_40 : Captures SecondPart of DVM of width40
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_secondpart_addr_range_40 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart_araddr_dvm_secondpart_40.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_secondpart_addr_range_40_vmid_unset  ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_MSB39TO32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_SECONDPART_40
    
    dvm_firstpart_secondpart_addr_range_40: cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_msb39to32_firstpart,araddr_dvm_secondpart_40 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup
   
    /**
    * Covergroup: trans_cross_ace_dvm_firstpart_secondpart_addr_range_3_vmid_unset2
    *
    * This covergroup is cross coverage of FirstPart of DVM (Virtual Address) on ARADDR[39:32],ARADDR[31:16] and SecondPart of DVM on ARADDR[39:4]
    *
    * Coverpoints:
    *
    * - araddr_dvm_firstpart_va_or_vmid: Captures firstpart of DVM Virtual address or VMID
    * - araddr_dvm_firsrpart_va_or_asid: Captures firstpart of DVM Virtual address or ASID
    * - araddr_dvm_secondpart_40 : Captures SecondPart of DVM of width40
    * .
    *
    * Cross coverpoints:
    *
    * -dvm_firstpart_secondpart_addr_range_32 : Crosses coverpoints araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_secondpart_32.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
    * .
    *
    */
    covergroup trans_cross_ace_dvm_firstpart_secondpart_addr_range_32_vmid_unset   ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_VMID_6_BIT_0
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_FIRSTPART_VA_OR_ASID
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_ARADDR_SECONDPART_32
    
    dvm_firstpart_secondpart_addr_range_32: cross araddr_dvm_firstpart_va_or_vmid,araddr_dvm_firsrpart_va_or_asid,araddr_dvm_secondpart_32 {
        
    option.weight = 1;
    }
    option.per_instance = 1;
    endgroup

`endif

`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF


   /**
    * Covergroup: trans_cross_axi_atomictype_exclusive_arcache
    *
    * This covergroup is cross coverage of READ Exclusive Access with all legel ARCache values.
    * The legal ARCACHE values for exclusive read access are
    * -Device Non-bufferable
    * -Device bufferable
    * -Normal Non-cacheable Non-bufferable
    * -Normal Non-cacheable Bufferable
    *
    * The protocol permits using the bufferable versions of ARCACHE during exclusive accesses,
    * but the system designer must ensure buffered exclusive accesses are still monitored by the slave i.e a more sensible design would be one where the 
    * buffer looks at the value of AxLOCK, and after seeing that the access is exclusive, decides to not return an early response.
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - atomic_type: Captures transaction atomic type
    * - cache_type: Captures transaction cache type
    * .
    *
    * Cross coverpoints:
    *
    * - axi_atomictype_exclusive_arcache: Crosses cover points read_xact_type, atomic_type,cache_type.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A7.2.4
    * .
    *
    */
  covergroup trans_cross_axi_atomictype_exclusive_arcache_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS_AXI3
    axi_atomictype_exclusive_arcache : cross read_xact_type, atomic_type,cache_type{
    ignore_bins   ignore_other_than_excl_read = (!binsof(atomic_type) intersect 
                                           {svt_axi_transaction::EXCLUSIVE}); 

    option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_exclusive_arcache_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS
    axi_atomictype_exclusive_arcache : cross read_xact_type, atomic_type,cache_type{
    ignore_bins   ignore_other_than_excl_read = (!binsof(atomic_type) intersect 
                                           {svt_axi_transaction::EXCLUSIVE}); 

    option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
 covergroup trans_cross_axi_atomictype_exclusive_arcache_locked_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_LOCKED_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS
    axi_atomictype_exclusive_arcache : cross read_xact_type, atomic_type,cache_type{
       option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_exclusive_arcache_normal_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_LOCKED_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS
    axi_atomictype_exclusive_arcache : cross read_xact_type, atomic_type,cache_type{
    option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_exclusive_arcache_locked_exclusive_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS
    axi_atomictype_exclusive_arcache : cross read_xact_type, atomic_type,cache_type{
    option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_exclusive_arcache_exclusive_axi3_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_NOT_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS
    axi_atomictype_exclusive_arcache : cross read_xact_type, atomic_type,cache_type{
    option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_atomictype_exclusive_arcache_normal_ace;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_LOCKED_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS
    axi_atomictype_exclusive_arcache : cross read_xact_type, atomic_type,cache_type{
       option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_exclusive_arcache_exclusive_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_NOT_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS
    axi_atomictype_exclusive_arcache : cross read_xact_type, atomic_type,cache_type{
    option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

   /**
    * Covergroup: trans_cross_axi_atomictype_exclusive_awcache
    *
    * This covergroup is cross coverage of WRITE Exclusive Access with all legel AWCache values.
    * The legal AWCACHE values for exclusive write access are
    * -Device bufferable
    * -Device Non-bufferable
    * -Normal Non-cacheable Non-bufferable
    * -Normal Non-cacheable Bufferable
    *
    * The protocol permits using the bufferable versions of AWCACHE during exclusive accesses,
    * but the system designer must ensure buffered exclusive accesses are still monitored by the slave i.e a more sensible design would be one where the 
    * buffer looks at the value of AxLOCK, and after seeing that the access is exclusive, decides to not return an early response.
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - atomic_type: Captures transaction atomic type
    * - cache_type: Captures transaction cache type
    * .
    *
    * Cross coverpoints:
    *
    * - axi_atomictype_exclusive_awcache: Crosses cover points write_xact_type, atomic_type,cache_type.
    * .
    * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; A7.2.4
    * .
    *
    */
  covergroup trans_cross_axi_atomictype_exclusive_awcache_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS_AXI3
    axi_atomictype_exclusive_awcache : cross write_xact_type, atomic_type,cache_type{
    ignore_bins   ignore_other_than_excl_write = (!binsof(atomic_type) intersect 
                                           {svt_axi_transaction::EXCLUSIVE}); 

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_exclusive_awcache_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS
    axi_atomictype_exclusive_awcache : cross write_xact_type, atomic_type,cache_type{
    ignore_bins   ignore_other_than_excl_write = (!binsof(atomic_type) intersect 
                                           {svt_axi_transaction::EXCLUSIVE}); 

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
covergroup trans_cross_axi_atomictype_exclusive_awcache_locked_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_LOCKED_AXI3  
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS
     axi_atomictype_exclusive_awcache : cross write_xact_type, atomic_type,cache_type{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_exclusive_awcache_locked_exclusive_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_AXI3  
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS
     axi_atomictype_exclusive_awcache : cross write_xact_type, atomic_type,cache_type{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_atomictype_exclusive_awcache_normal_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_LOCKED_AXI3  
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS
     axi_atomictype_exclusive_awcache : cross write_xact_type, atomic_type,cache_type{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_atomictype_exclusive_awcache_exclusive_axi3_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_NOT_AXI3  
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS
     axi_atomictype_exclusive_awcache : cross write_xact_type, atomic_type,cache_type{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_exclusive_awcache_normal_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_LOCKED_AXI3  
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS
     axi_atomictype_exclusive_awcache : cross write_xact_type, atomic_type,cache_type{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_atomictype_exclusive_awcache_exclusive_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_NOT_AXI3  
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_EXCLUSIVE_ACCESS
     axi_atomictype_exclusive_awcache : cross write_xact_type, atomic_type,cache_type{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF



  /**
  *  Covergroup     : trans_cross_ace_writeunique_awdomain_awprot
  *
  * Coverpoints:
  *
  * - coherent_write_xact_type:  Captures writeunique coherent write transaction
  * - domain_type : Captures domain type
  * - prot_type : Captures transaction protection type
  * .
  * Cross coverpoints:
  * - writeunique_awdomain_awprot : Crosses cover points
  *    coherent_write_xact_type and domain_type and prot_type
  * .
  * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.1.6
  * .
  *
  */

  covergroup trans_cross_ace_writeunique_awdomain_awprot ;
    //`SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    coherent_write_xact_type : coverpoint cov_item.coherent_xact_type iff(cov_coherent_xact_type_flag){
      bins coherent_writeunique_xact = {svt_axi_transaction::WRITEUNIQUE};
      option.weight = 1;
    }
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE

    writeunique_awdomain_awprot : cross coherent_write_xact_type, domain_type, prot_type {


      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                    {svt_axi_transaction::WRITEUNIQUE}) &&
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_not_write_unique = (!binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITEUNIQUE});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /**
  *  Covergroup     : trans_cross_ace_readonce_ardomain_arprot
  *
  * Coverpoints:
  *
  * - coherent_read_xact_type:  Captures readonce coherent read transaction
  * - domain_type : Captures domain type
  * - prot_type : Captures transaction protection type
  * .
  * Cross coverpoints:
  * - readonce_ardomain_arprot : Crosses cover points
  *    coherent_read_xact_type and domain_type and prot_type
  * .
  * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.1.6
  * .
  *
  */

  covergroup trans_cross_ace_readonce_ardomain_arprot ;
    //`SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    coherent_read_xact_type : coverpoint cov_item.coherent_xact_type iff(cov_coherent_xact_type_flag){
      bins coherent_readonce_xact = {svt_axi_transaction::READONCE};
      option.weight = 1;
    }
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE

    readonce_ardomain_arprot : cross coherent_read_xact_type, domain_type, prot_type {


      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                    {svt_axi_transaction::READONCE}) &&
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_not_readonce = (!binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::READONCE});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup


  /**
  * Covergroup     : trans_cross_ace_awprot_awbarrier_memory_sync
  *
  * Coverpoints:
  *
  * - coherent_write_xact_type:  Captures coherent write transaction
  * - barrier_type : Captures write barrier
  * - prot_type : Captures transaction protection type
  * .
  * Cross coverpoints:
  * - awprot_awbarrier_memory_sync: Crosses cover points
  *   write transaction of barrier_type MEMORY_BARRIER & SYNC_BARRIER with awprot
  * .
  * The following bins are ignored:
  * -bins that interset NORMAL_ACCESS_RESPECT_BARRIER and NORMAL_ACCESS_IGNORE_BARRIER
  * -bins that intersect transaction types other than WRITEBARRIER
  * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.1.6
  * .
  *
  */

  covergroup trans_cross_ace_awprot_awbarrier_memory_sync ;
    //`SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    coherent_write_xact_type : coverpoint cov_item.coherent_xact_type iff(cov_coherent_xact_type_flag){
      bins coherent_writebarrier_xact = {svt_axi_transaction::WRITEBARRIER};
      option.weight = 1;
    }
    // Only MEMORY_BARRIER and SYNC_BARRIER are being covered, so we need to use only the BARRIER_SET macro
    //`SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_TYPE 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE
    awprot_awbarrier_memory_sync : cross coherent_write_xact_type, barrier_type, prot_type {

      ignore_bins ignore_normal = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});
      ignore_bins ignore_non_write_barrier = (!binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup


  /**
  * Covergroup     : trans_cross_ace_arprot_arbarrier_memory_sync
  *
  * Coverpoints:
  *
  * - coherent_read_xact_type:  Captures coherent read transaction
  * - barrier_type : Captures read barrier
  * - prot_type : Captures transaction protection type
  * .
  * Cross coverpoints:
  * - arprot_arbarrier_memory_sync: Crosses cover points
  *   read transaction of barrier_type MEMORY_BARRIER & SYNC_BARRIER with arprot
  * .
  * The following bins are ignored:
  * -bins that interset NORMAL_ACCESS_RESPECT_BARRIER and NORMAL_ACCESS_IGNORE_BARRIER
  * -bins that intersect transaction types other than READBARRIER
  * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.1.6
  * .
  *
  */

  covergroup trans_cross_ace_arprot_arbarrier_memory_sync ;
    //`SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    coherent_read_xact_type : coverpoint cov_item.coherent_xact_type iff(cov_coherent_xact_type_flag){
      bins coherent_readbarrier_xact = {svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    // Only MEMORY_BARRIER and SYNC_BARRIER are being covered, so we need to use only the BARRIER_SET macro
    //`SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_TYPE 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE

    arprot_arbarrier_memory_sync : cross coherent_read_xact_type, barrier_type, prot_type {

      ignore_bins ignore_normal = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});

      ignore_bins ignore_non_read_barrier = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
   
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  /**
  * Covergroup:trans_axi_read_outstanding_xact_same_arid_cache_modifiable_bit 
  *
  * Coverpoints:read_outstanding_xact_same_arid_cache_modifiable_bit
  *
  * - This coverpoint covers the scenario in which master can issue multiple outstanding READ transactions
  * with same ARID,taking ARCACHE Modifiable bit into consideration.
  *.
  *
  * Bins are interpreted as follows:
  * - cache_modifiable_followed_by_modifiable: Bin is hit when an outstanding transaction with ARCACHE[1]=1 is followed by another transaction with ARCACHE[1]=1.
  * - cache_modifiable_followed_by_nonmodifiable: Bin is hit when an outstanding transaction with ARCACHE[1]=1 is followed by another transaction with ARCACHE[1]=0.
  * - cache_nonmodifiable_followed_by_modifiable: Bin is hit when an outstanding transaction with ARCACHE[1]=0 is followed by another transaction with ARCACHE[1]=1.
  * - cache_nonmodifiable_followed_by_nonmodifiable: Bin is hit when an outstanding transaction with ARCACHE[1]=0 is followed by another transaction with ARCACHE[1]=0.
  * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613 ; section A5.1
  * .
  *
  */
  covergroup trans_axi_read_outstanding_xact_same_arid_cache_modifiable_bit;
  read_outstanding_xact_same_arid_cache_modifiable_bit : coverpoint read_outstanding_xact_same_arid_cache_modifiable_bit{
  bins cache_nonmodifiable_followed_by_nonmodifiable   = {0};
  bins cache_nonmodifiable_followed_by_modifiable      = {1};
  bins cache_modifiable_followed_by_nonmodifiable      = {2};
  bins cache_modifiable_followed_by_modifiable         = {3};
  option.weight = 1;
  }              
  option.per_instance = 1;
  endgroup

  /**
  * Covergroup:trans_axi_read_outstanding_xact_diff_arid_cache_modifiable_bit
  *
  * Coverpoints:read_outstanding_xact_diff_arid_cache_modifiable_bit
  *
  * - This coverpoint covers the scenario in which master can issue multiple outstanding READ transactions
  * with different ARID,taking ARCACHE Modifiable bit into consideration.
  *.
  *
  * Bins are interpreted as follows:
  * - cache_modifiable_followed_by_modifiable: Bin is hit when an outstanding transaction with ARCACHE[0]=1 is followed by another transaction with ARCACHE[0]=1.
  * - cache_modifiable_followed_by_nonmodifiable: Bin is hit when an outstanding transaction with ARCACHE[0]=1 is followed by another transaction with ARCACHE[0]=0.
  * - cache_nonmodifiable_followed_by_modifiable: Bin is hit when an outstanding transaction with ARCACHE[0]=0 is followed by another transaction with ARCACHE[0]=1.
  * - cache_nonmodifiable_followed_by_nonmodifiable: Bin is hit when an outstanding transaction with ARCACHE[0]=0 is followed by another transaction with ARCACHE[0]=0.
  * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613 ; section A5.1
  * .
  *
  */
  covergroup trans_axi_read_outstanding_xact_diff_arid_cache_modifiable_bit;
  read_outstanding_xact_diff_arid_cache_modifiable_bit : coverpoint read_outstanding_xact_diff_arid_cache_modifiable_bit{
  bins cache_nonmodifiable_followed_by_nonmodifiable   = {0};
  bins cache_nonmodifiable_followed_by_modifiable      = {1};
  bins cache_modifiable_followed_by_nonmodifiable      = {2};
  bins cache_modifiable_followed_by_modifiable         = {3};
  option.weight = 1;
  }              
  option.per_instance = 1;
  endgroup

  /**
  * Covergroup:trans_axi_read_outstanding_xact_diff_arid_device_cacheable_bit
  *
  * Coverpoints:read_outstanding_xact_diff_arid_device_cacheable_bit
  *
  * - This coverpoint covers the scenario in which master can issue multiple outstanding READ transactions
  * with different ARID,taking memory types by ARCACHE[3:0] into consideration.
  *.
  *
  * Bins are interpreted as follows:
  * - device_nonbufferable_followed_by_device_nonbufferable: Bin is hit when an outstanding transaction with ARCACHE[3:0]= 4'b0000 is followed by another transaction with ARCACHE[3:0]= 4'b0000.
  * - device_nonbufferable_followed_by_device_bufferable: Bin is hit when an outstanding transaction with ARCACHE[3:0]= 4'b0000 is followed by another transaction with ARCACHE[3:0]= 4'b0001.
  * - device_bufferable_followed_by_device_nonbufferable: Bin is hit when an outstanding transaction with ARCACHE[3:0]= 4'b0001 is followed by another transaction with ARCACHE[3:0]= 4'b0000.
  * - device_bufferable_followed_by_device_bufferable: Bin is hit when an outstanding transaction with ARCACHE[3:0]= 4'b0001 is followed by another transaction with ARCACHE[3:0]= 4'b0001.
  *
  * - normal_noncacheable_nonbufferable_followed_by_noncacheable_nonbufferable: Bin is hit when an outstanding transaction with ARCACHE[3:0]= 4'b0010 is followed by another transaction with ARCACHE[3:0]= 4'b0010.
  * - normal_noncacheable_nonbufferable_followed_by_noncacheable_bufferable: Bin is hit when an outstanding transaction with ARCACHE[3:0]= 4'b0010 is followed by another transaction with ARCACHE[3:0]= 4'b0011.
  * - normal_noncacheable_bufferable_followed_by_noncacheable_nonbufferable: Bin is hit when an outstanding transaction with ARCACHE[3:0]= 4'b0011 is followed by another transaction with ARCACHE[3:0]= 4'b0010.
  * - normal_noncacheable_bufferable_followed_by_noncacheable_bufferable: Bin is hit when an outstanding transaction with ARCACHE[3:0]= 4'b0011 is followed by another transaction with ARCACHE[3:0]= 4'b0011.
  * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613 ; section A4.4
  * .
  *
  */
  covergroup trans_axi_read_outstanding_xact_diff_arid_device_cacheable_bit;
  read_outstanding_xact_diff_arid_device_cacheable_bit : coverpoint read_outstanding_xact_diff_arid_device_cacheable_bit{
  bins device_nonbufferable_followed_by_device_nonbufferable                      = {0};
  bins device_nonbufferable_followed_by_device_bufferable                         = {1};
  bins device_bufferable_followed_by_device_nonbufferable                         = {2};
  bins device_bufferable_followed_by_device_bufferable                            = {3};
  bins normal_noncacheable_nonbufferable_followed_by_noncacheable_nonbufferable   = {4};
  bins normal_noncacheable_nonbufferable_followed_by_noncacheable_bufferable      = {5};
  bins normal_noncacheable_bufferable_followed_by_noncacheable_nonbufferable      = {6};
  bins normal_noncacheable_bufferable_followed_by_noncacheable_bufferable         = {7};
  option.weight = 1;
  }              
  option.per_instance = 1;
  endgroup

  /**
  * Covergroup:trans_axi_write_outstanding_xact_diff_awid_device_cacheable_bit
  *
  * Coverpoints:write_outstanding_xact_diff_awid_device_cacheable_bit
  *
  * - This coverpoint covers the scenario in which master can issue multiple outstanding WRITE transactions
  * with different AWID,taking memory types by AWCACHE[3:0] into consideration.
  *.
  *
  * Bins are interpreted as follows:
  * - device_nonbufferable_followed_by_device_nonbufferable: Bin is hit when an outstanding transaction with AWCACHE[3:0]= 4'b0000 is followed by another transaction with AWCACHE[3:0]= 4'b0000.
  * - device_nonbufferable_followed_by_device_bufferable: Bin is hit when an outstanding transaction with AWCACHE[3:0]= 4'b0000 is followed by another transaction with AWCACHE[3:0]= 4'b0001.
  * - device_bufferable_followed_by_device_nonbufferable: Bin is hit when an outstanding transaction with AWCACHE[3:0]= 4'b0001 is followed by another transaction with AWCACHE[3:0]= 4'b0000.
  * - device_bufferable_followed_by_device_bufferable: Bin is hit when an outstanding transaction with AWCACHE[3:0]= 4'b0001 is followed by another transaction with AWCACHE[3:0]= 4'b0001.
  *
  * - normal_noncacheable_nonbufferable_followed_by_noncacheable_nonbufferable: Bin is hit when an outstanding transaction with AWCACHE[3:0]= 4'b0010 is followed by another transaction with AWCACHE[3:0]= 4'b0010.
  * - normal_noncacheable_nonbufferable_followed_by_noncacheable_bufferable: Bin is hit when an outstanding transaction with AWCACHE[3:0]= 4'b0010 is followed by another transaction with AWCACHE[3:0]= 4'b0011.
  * - normal_noncacheable_bufferable_followed_by_noncacheable_nonbufferable: Bin is hit when an outstanding transaction with AWCACHE[3:0]= 4'b0011 is followed by another transaction with AWCACHE[3:0]= 4'b0010.
  * - normal_noncacheable_bufferable_followed_by_noncacheable_bufferable: Bin is hit when an outstanding transaction with AWCACHE[3:0]= 4'b0011 is followed by another transaction with AWCACHE[3:0]= 4'b0011.
  * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613 ; section A4.4
  * .
  *
  */
  covergroup trans_axi_write_outstanding_xact_diff_awid_device_cacheable_bit;
  write_outstanding_xact_diff_awid_device_cacheable_bit : coverpoint write_outstanding_xact_diff_awid_device_cacheable_bit{
  bins device_nonbufferable_followed_by_device_nonbufferable                      = {0};
  bins device_nonbufferable_followed_by_device_bufferable                         = {1};
  bins device_bufferable_followed_by_device_nonbufferable                         = {2};
  bins device_bufferable_followed_by_device_bufferable                            = {3};
  bins normal_noncacheable_nonbufferable_followed_by_noncacheable_nonbufferable   = {4};
  bins normal_noncacheable_nonbufferable_followed_by_noncacheable_bufferable      = {5};
  bins normal_noncacheable_bufferable_followed_by_noncacheable_nonbufferable      = {6};
  bins normal_noncacheable_bufferable_followed_by_noncacheable_bufferable         = {7};
  option.weight = 1;
  }              
  option.per_instance = 1;
  endgroup

  /**
  * Covergroup:trans_axi_write_outstanding_xact_same_awid_cache_modifiable_bit
  *
  * Coverpoints:write_outstanding_xact_same_awid_cache_modifiable_bit
  *
  * - This coverpoint covers the scenario in which master can issue multiple outstanding WRITE transactions
  * with same AWID's,taking AWCACHE Modifiable bit into consideration.
  *.
  *
  * Bins are interpreted as follows:
  * - cache_modifiable_followed_by_modifiable: Bin is hit when an outstanding transaction with AWCACHE[1]=1 is followed by another transaction with AWCACHE[1]=1.
  * - cache_modifiable_followed_by_nonmodifiable: Bin is hit when an outstanding transaction with AWCACHE[1]=1 is followed by another transaction with AWCACHE[1]=0.
  * - cache_nonmodifiable_followed_by_modifiable: Bin is hit when an outstanding transaction with AWCACHE[1]=0 is followed by another transaction with AWCACHE[1]=1.
  * - cache_nonmodifiable_followed_by_nonmodifiable: Bin is hit when an outstanding transaction with AWCACHE[1]=0 is followed by another transaction with AWCACHE[1]=0.
  * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613 ; section A5.1
  * .
  *
  */
  covergroup trans_axi_write_outstanding_xact_same_awid_cache_modifiable_bit;
  write_outstanding_xact_same_awid_cache_modifiable_bit : coverpoint write_outstanding_xact_same_awid_cache_modifiable_bit{
  bins cache_nonmodifiable_followed_by_nonmodifiable   = {0};
  bins cache_nonmodifiable_followed_by_modifiable      = {1};
  bins cache_modifiable_followed_by_nonmodifiable      = {2};
  bins cache_modifiable_followed_by_modifiable         = {3};
  option.weight = 1;
  }              
  option.per_instance = 1;
  endgroup

  /**
  * Covergroup:trans_axi_write_outstanding_xact_diff_awid_cache_modifiable_bit
  *
  * Coverpoints:write_outstanding_xact_diff_awid_cache_modifiable_bit
  *
  * - This coverpoint covers the scenario in which master can issue multiple outstanding WRITE transactions
  * with diff AWID's,taking AWCACHE Modifiable bit into consideration.
  *.
  *
  * Bins are interpreted as follows:
  * - cache_modifiable_followed_by_modifiable: Bin is hit when an outstanding transaction with AWCACHE[0]=1 is followed by another transaction with AWCACHE[0]=1.
  * - cache_modifiable_followed_by_nonmodifiable: Bin is hit when an outstanding transaction with AWCACHE[0]=1 is followed by another transaction with AWCACHE[0]=0.
  * - cache_nonmodifiable_followed_by_modifiable: Bin is hit when an outstanding transaction with AWCACHE[0]=0 is followed by another transaction with AWCACHE[0]=1.
  * - cache_nonmodifiable_followed_by_nonmodifiable: Bin is hit when an outstanding transaction with AWCACHE[0]=0 is followed by another transaction with AWCACHE[0]=0.
  * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613 ; section A5.1
  * .
  *
  */
  covergroup trans_axi_write_outstanding_xact_diff_awid_cache_modifiable_bit;
  write_outstanding_xact_diff_awid_cache_modifiable_bit : coverpoint write_outstanding_xact_diff_awid_cache_modifiable_bit{
  bins cache_nonmodifiable_followed_by_nonmodifiable   = {0};
  bins cache_nonmodifiable_followed_by_modifiable      = {1};
  bins cache_modifiable_followed_by_nonmodifiable      = {2};
  bins cache_modifiable_followed_by_modifiable         = {3};
  option.weight = 1;
  }              
  option.per_instance = 1;
  endgroup

   /** 
   *  Covergroup:  axi_wstrb_to_signal_unaligned_start_address
   *  
   * - This cover group covers the scenario in which a master can provide an aligned address to a write transaction, and use the write strobes to indicate unaligned start address.
   * - Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A:3.4.3 
   * .
   *
   */

  covergroup axi_wstrb_to_signal_unaligned_start_address @(wstrb_to_signal_unaligned_start_address_event);
    type_option.comment = "Coverage for WSTRB to signal UNALIGNED START ADDRESS";
    option.per_instance = 1;
    wstrb_to_signal_unaligned_start_address : coverpoint this.wstrb_to_signal_unaligned_start_address {
      bins wstrb_to_signal_unaligned_start_addr = {`SVT_AXI_WSTRB_UNALIGNED_START_ADDR};
    }
  endgroup
`endif // SVT_AXI_MON_CFG_BASED_COV_GRP_DEF


`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

    /**
    * Covergroup: trans_cross_axi3_arcache_modifiable_bit_read_unaligned_transfer
    * This cover group crosses bit ARCACHE[1] with unaligned read transfers.
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - addr_offset: Captures transaction address offset information
    * - transfer_size: Captures transaction burst size
    * - burst_length: Captures transaction burst length
    * - cache_type_modifiable_bit: Captures ARCACHE[1]
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_read_arcache_modifiable_bit_unaligned_transfer: Crosses cover points read_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A:4:4:2
    */
  covergroup trans_cross_axi3_arcache_modifiable_bit_read_unaligned_transfer ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi3_arcache_modifiable_bit_read_unaligned_transfer : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_cross_axi4_arcache_modifiable_bit_read_unaligned_transfer
    * This cover group crosses bit ARCACHE[1] with unaligned read transfers.
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - addr_offset: Captures transaction address offset information
    * - transfer_size: Captures transaction burst size
    * - burst_length: Captures transaction burst length
    * - cache_type_modifiable_bit: Captures ARCACHE[1]
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_read_arcache_modifiable_bit_unaligned_transfer: Crosses cover points read_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A:4:4:2
    */
  covergroup trans_cross_axi4_arcache_modifiable_bit_read_unaligned_transfer ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi4_arcache_modifiable_bit_read_unaligned_transfer : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit  {
    ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
    ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else // SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
    covergroup trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_axi3_dweq_32bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_arcache_modifiable_bit_read_unaligned_transfer_axi3_dweq_32bit : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_axi3_dweq_64bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_arcache_modifiable_bit_read_unaligned_transfer_axi3_dweq_64bit : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_axi3_dweq_128bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_arcache_modifiable_bit_read_unaligned_transfer_axi3_dweq_128bit : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

 covergroup trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_axi4_dweq_32bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_arcache_modifiable_bit_read_unaligned_transfer_axi4_dweq_32bit : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_axi4_dweq_64bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_arcache_modifiable_bit_read_unaligned_transfer_axi4_dweq_64bit : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_axi4_dweq_128bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_arcache_modifiable_bit_read_unaligned_transfer_axi4_dweq_128bit : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

 covergroup trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_ace_dweq_32bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_arcache_modifiable_bit_read_unaligned_transfer_ace_dweq_32bit : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_ace_dweq_64bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_arcache_modifiable_bit_read_unaligned_transfer_ace_dweq_64bit : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_ace_dweq_128bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_arcache_modifiable_bit_read_unaligned_transfer_ace_dweq_128bit : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`endif

`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  /**
    * Covergroup: trans_cross_axi3_awcache_modifiable_bit_write_unaligned_transfer
    * This cover group crosses bit AWCACHE[1] with unaligned write transfers.
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - addr_offset: Captures transaction address offset information
    * - transfer_size: Captures transaction burst size
    * - burst_length: Captures transaction burst length
    * - cache_type_modifiable_bit: Captures AWCACHE[1]
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_awcache_modifiable_bit_write_unaligned_transfer: Crosses cover points write_xact_type, burst_type, addr_offset, transfer_size, burst_length cache_type_modifiable_bit
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A:4:4:2
    */
  covergroup trans_cross_axi3_awcache_modifiable_bit_write_unaligned_transfer ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi3_awcache_modifiable_bit_write_unaligned_transfer : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_cross_axi4_awcache_modifiable_bit_write_unaligned_transfer
    * This cover group crosses bit AWCACHE[1] with unaligned write transfers.
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - addr_offset: Captures transaction address offset information
    * - transfer_size: Captures transaction burst size
    * - burst_length: Captures transaction burst length
    * - cache_type_modifiable_bit: Captures AWCACHE[1]
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_awcache_modifiable_bit_write_unaligned_transfer: Crosses cover points write_xact_type, burst_type, addr_offset, transfer_size, burst_length cache_type_modifiable_bit
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A:4:4:2
    */
  covergroup trans_cross_axi4_awcache_modifiable_bit_write_unaligned_transfer ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi4_awcache_modifiable_bit_write_unaligned_transfer : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {
    ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
    ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else // SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer_axi3_dweq_32bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_awcache_modifiable_bit_write_unaligned_transfer_axi3_dweq_32bit : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer_axi3_dweq_64bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_awcache_modifiable_bit_write_unaligned_transfer_axi3_dweq_64bit : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer_axi3_dweq_128bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_awcache_modifiable_bit_write_unaligned_transfer_axi3_dweq_128bit : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

 covergroup trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer_axi4_dweq_32bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_awcache_modifiable_bit_write_unaligned_transfer_axi4_dweq_32bit : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer_axi4_dweq_64bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_awcache_modifiable_bit_write_unaligned_transfer_axi4_dweq_64bit : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer_axi4_dweq_128bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_awcache_modifiable_bit_write_unaligned_transfer_axi4_dweq_128bit : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

 covergroup trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer_ace_dweq_32bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_awcache_modifiable_bit_write_unaligned_transfer_ace_dweq_32bit : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer_ace_dweq_64bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_awcache_modifiable_bit_write_unaligned_transfer_ace_dweq_64bit : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer_ace_dweq_128bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE_MODIFIABLE_BIT
    axi_awcache_modifiable_bit_write_unaligned_transfer_ace_dweq_128bit : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length, cache_type_modifiable_bit {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`endif // SVT_AXI_MON_CFG_BASED_COV_GRP_DEF


`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  /**
    * Covergroup: trans_cross_axi_fixed_burst_wstrb
    * This cover group crosses AXI Fixed burst type with write strobe
    *
    * Covers the cross of  fixed burst type, & WSTRB 
    * Coverpoints:
    *
    * - burst_type: Captures transaction burst type
    * - wstrb: Captures write strobe values
    * 
    *
    * Cross coverpoints:
    *
    * - axi_fixed_burst_wstrb : Crosses cover points burst_type,wstrb 
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A:3.4.1
    */

    covergroup trans_cross_axi_fixed_burst_wstrb;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WSTRB
     axi_fixed_burst_wstrb : cross burst_type,wstrb {
      ignore_bins   ignore_burst_type_other_than_fixed_burst =  !binsof(burst_type.fixed_burst);
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup 

   /** 
   * Covergroup:  axi_four_excl_normal_sequence
   *
   * This cover group covers specific combinations of exclusive and normal
   * transactions, for a sequence of four transactions. For eg.
   * Excl-Normal-Excl-Normal,Normal-Normal-Excl-Normal etc. 
   * <br>
   * Following sequences are supported:
   *   -  NR_NR_NR_EX
   *   -  NR_NR_EX_NR
   *   -  NR_NR_EX_EX
   *   -  NR_EX_NR_NR
   *   -  NR_EX_NR_EX
   *   -  NR_EX_EX_NR
   *   -  NR_EX_EX_EX
   *   -  EX_NR_NR_NR
   *   -  EX_NR_NR_EX
   *   -  EX_NR_EX_NR
   *   -  EX_NR_EX_EX
   *   -  EX_EX_NR_NR
   *   -  EX_EX_NR_EX
   *   -  EX_EX_EX_NR
   *   .
   */ 

  covergroup axi_four_excl_normal_sequence @(four_excl_normal_seq_event);
    type_option.comment = "Coverage for Four Exclusive/Normal transactions,for Ex:NR_EX_NR_EX,EX_NR_NR_EX";
    option.per_instance = 1;
     four_excl_normal_sequence: coverpoint this.four_excl_normal_sequence {
      bins bin_NR_NR_NR_EX_SEQ =  {`SVT_AXI_NR_NR_NR_EX_SEQ};
      bins bin_NR_NR_EX_NR_SEQ =  {`SVT_AXI_NR_NR_EX_NR_SEQ};
      bins bin_NR_NR_EX_EX_SEQ =  {`SVT_AXI_NR_NR_EX_EX_SEQ};
      bins bin_NR_EX_NR_NR_SEQ =  {`SVT_AXI_NR_EX_NR_NR_SEQ};
      bins bin_NR_EX_NR_EX_SEQ =  {`SVT_AXI_NR_EX_NR_EX_SEQ};
      bins bin_NR_EX_EX_NR_SEQ =  {`SVT_AXI_NR_EX_EX_NR_SEQ};
      bins bin_NR_EX_EX_EX_SEQ =  {`SVT_AXI_NR_EX_EX_EX_SEQ};
      bins bin_EX_NR_NR_NR_SEQ =  {`SVT_AXI_EX_NR_NR_NR_SEQ};
      bins bin_EX_NR_NR_EX_SEQ =  {`SVT_AXI_EX_NR_NR_EX_SEQ};
      bins bin_EX_NR_EX_NR_SEQ =  {`SVT_AXI_EX_NR_EX_NR_SEQ};
      bins bin_EX_NR_EX_EX_SEQ =  {`SVT_AXI_EX_NR_EX_EX_SEQ};
      bins bin_EX_EX_NR_NR_SEQ =  {`SVT_AXI_EX_EX_NR_NR_SEQ};
      bins bin_EX_EX_NR_EX_SEQ =  {`SVT_AXI_EX_EX_NR_EX_SEQ};
      bins bin_EX_EX_EX_NR_SEQ =  {`SVT_AXI_EX_EX_EX_NR_SEQ};
    }
  endgroup
  
  /** 
   * Covergroup:  axi_four_state_rd_wr_burst_sequence
   *
   * This cover group covers specific combinations of read and write
   * transactions, for a sequence of four transactions. For eg.
   * Write-Write-Write-Write or Write-Read-Write-Read, etc. This covergroup is
   * hit when address phase completion of four transactions are observed in a
   * specific combination as described above. When address phases of READ and
   * WRITE transactions get completed at same time, it is not deterministic
   * whether it is a read-write or write-read scenario. In such situation,
   * either sequence containing read-write or write-read may get hit.
   * <br>
   * Following sequences are currently supported:
   *   -  WR_WR_WR_WR
   *   -  WR_RD_WR_RD
   *   -  WR_WR_RD_RD
   *   -  RD_RD_WR_WR
   *   -  RD_RD_RD_RD
   *   -  WR_WR_WR_RD
   *   -  RD_WR_RD_WR
   *   -  RD_RD_RD_WR
   *   .
   * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A:3.4.1
   */ 

  covergroup axi_four_state_rd_wr_burst_sequence @(four_state_rd_wr_event);
    type_option.comment = "Coverage for Four State READ/WRITE BURST,for Ex:WR-WR-RD-RD, RD-WR-RD-WR, RD-RD-RD-WR etc";
    option.per_instance = 1;
     four_state_rd_wr_burst_sequence: coverpoint this.four_state_rd_wr_burst_sequence {
      bins bin_WR_WR_WR_WR_SEQ =  {`SVT_AXI_WR_WR_WR_WR_SEQ};
      bins bin_WR_RD_WR_RD_SEQ =  {`SVT_AXI_WR_RD_WR_RD_SEQ};
      bins bin_RD_WR_RD_WR_SEQ =  {`SVT_AXI_RD_WR_RD_WR_SEQ};
      bins bin_WR_WR_RD_RD_SEQ =  {`SVT_AXI_WR_WR_RD_RD_SEQ};
      bins bin_RD_RD_WR_WR_SEQ =  {`SVT_AXI_RD_RD_WR_WR_SEQ};
      bins bin_RD_RD_RD_RD_SEQ =  {`SVT_AXI_RD_RD_RD_RD_SEQ};
      bins bin_RD_RD_RD_WR_SEQ =  {`SVT_AXI_RD_RD_RD_WR_SEQ};
      bins bin_WR_WR_WR_RD_SEQ =  {`SVT_AXI_WR_WR_WR_RD_SEQ};
    }
  endgroup

  /** 
   * Coverage group for covering Back To Back READ BURST. 
   * This covergroup is triggered when address phase of first READ xact has completed and
   * immediately next clock address phase of second READ xact has started
   */
  covergroup axi_back_to_back_read_burst_sequence @(back_to_back_read_burst_event);
    type_option.comment = "Coverage for Back to Back Read Burst READ -> READ";
    option.per_instance = 1;
    back_to_back_read_burst_sequence : coverpoint this.back_to_back_read_burst_sequence {
      bins back_to_back_read_burst_seq = {`SVT_AXI_BACK_TO_BACK_READ_BURST_SEQ};
    }
  endgroup
  
  /** 
   * Coverage group for covering Back To Back WRITE BURST. 
   * This covergroup is triggered when address phase of first WRITE xact has completed and
   * immediately next clock address phase of second  WRITE xact has started
   */
  covergroup axi_back_to_back_write_burst_sequence @(back_to_back_write_burst_event);
    type_option.comment = "Coverage for Back to Back Write Burst WRITE -> WRITE";
    option.per_instance = 1;
    back_to_back_write_burst_sequence : coverpoint this.back_to_back_write_burst_sequence {
      bins back_to_back_write_burst_seq = {`SVT_AXI_BACK_TO_BACK_WRITE_BURST_SEQ};
    }
  endgroup


   /** 
   * Coverage group for covering Read/Write Completed out of order with ARID != AWID
   */

 covergroup axi_write_read_diff_id_completed_out_of_order@(cover_arid_awid_diff_out_of_order_event);
    type_option.comment = "Coverage for OOO completion of READ and WRITE transactions with ARID!=AWID";
    option.per_instance = 1;
    write_completed_out_of_order : coverpoint this.write_completed_out_of_order {
      bins write_completed_OOO = {`SVT_AXI_WRITE_OOO};}

    read_completed_out_of_order : coverpoint this.read_completed_out_of_order {
      bins read_completed_OOO = {`SVT_AXI_READ_OOO};}
 endgroup

 /** 
   * Coverage group for covering Read/Write Completed out of order with ARID==AWID
   */

  covergroup axi_write_read_same_id_completed_out_of_order@(cover_arid_awid_equal_out_of_order_event);
    type_option.comment = "Coverage for OOO completion of READ and WRITE transactions with ARID==AWID";
    option.per_instance = 1;
    write_completed_out_of_order_same_id_as_read : coverpoint this.write_completed_out_of_order_same_id_as_read {
      bins write_completed_OOO_same_id_as_read = {`SVT_AXI_WRITE_OOO_SAME_ID_AS_READ};
    }

    read_completed_out_of_order_same_id_as_write : coverpoint this.read_completed_out_of_order_same_id_as_write {
      bins read_completed_OOO_same_id_as_write = {`SVT_AXI_READ_OOO_SAME_ID_AS_WRITE};
    }
  endgroup

 /** 
   * Covergroup : trans_cross_axi_out_of_order_write_resp_count
   *
   * This Covergroup is for covering write_resp out_of_order count.
   *
   * Coverpoint:
   * axi_write_resp_OOO_count : Captures write_resp out_of_order count
   *.
   */
  covergroup trans_cross_axi_out_of_order_write_resp_count @(cov_out_of_order_write_response_depth_event);
   axi_write_resp_OOO_count: coverpoint this.axi_write_resp_OOO_count  { 
      bins write_rsp_ooo_count = {1};
      option.weight = 1;
   }
    option.per_instance = 1;
  endgroup

 /** 
   * Covergroup : trans_cross_axi_out_of_order_read_resp_count
   *
   * This Covergroup is for covering read_resp out_of_order count.
   *
   * Coverpoint :
   * axi_read_resp_OOO_count : Captures read_resp out_of_order count
   * .
   */
  covergroup trans_cross_axi_out_of_order_read_resp_count @(cov_out_of_order_read_response_depth_event);
   axi_read_resp_OOO_count: coverpoint this.axi_read_resp_OOO_count  { 
       bins read_rsp_ooo_count = {1};
       option.weight = 1;
   }
  option.per_instance = 1;
  endgroup
`endif //  `ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
 /**
    * Covergroup: trans_cross_axi_atomictype_rresp
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - atomic_type: Captures transaction atomic type
    * - rresp: Captures transaction response
    * .
    *
    * Cross coverpoints:
    *
    * - axi_atomictype_rresp: Crosses cover points read_xact_type, atomic_type,rresp.
    * This covergroup is triggered when an exclusive READ transaction with rresp of exokay is observed 
    * .
    *
    */
  covergroup trans_cross_axi_atomictype_rresp ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP
    axi_atomictype_rresp : cross read_xact_type, atomic_type,rresp{
    ignore_bins   ignore_excl_read_other_than_exokay_resp =  !binsof(rresp.exokay_resp) || !binsof(atomic_type.exclusive) || !binsof(read_xact_type.read_xact);
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else
 covergroup trans_cross_axi_atomictype_rresp_locked_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_LOCKED_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_atomictype_rresp : cross read_xact_type, atomic_type,rresp{
         option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_rresp_normal_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_LOCKED_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_atomictype_rresp : cross read_xact_type, atomic_type,rresp{
          option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_rresp_locked_exclusive_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_ALL
    axi_atomictype_rresp : cross read_xact_type, atomic_type,rresp{
    ignore_bins   ignore_excl_read_other_than_exokay_resp =  !binsof(rresp.exokay_resp) || !binsof(atomic_type.exclusive) || !binsof(read_xact_type.read_xact);
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_rresp_exclusive_axi3_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_NOT_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_ALL
     axi_atomictype_rresp : cross read_xact_type, atomic_type,rresp{
     option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_rresp_exclusive_axi4lite ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_LOCKED_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_NO_EXCLUSIVE_AXI4_LITE
     axi_atomictype_rresp : cross read_xact_type, atomic_type,rresp{
          option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_atomictype_rresp_normal_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_LOCKED_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_atomictype_rresp : cross read_xact_type, atomic_type,rresp{
         option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_atomictype_rresp_exclusive_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_NOT_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_ALL
    axi_atomictype_rresp : cross read_xact_type, atomic_type,rresp{
          option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 
`endif
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  /**
    * Covergroup: trans_cross_axi_atomictype_bresp
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - atomic_type: Captures transaction atomic type
    * - bresp: Captures transaction response
    * 
    *
    * Cross coverpoints:
    *
    * - axi_atomictype_bresp: Crosses cover points write_xact_type, atomic_type,bresp.
    * This covergroup is triggered when an exclusive Write transaction with bresp of okay/exokay is observed 
    * .
    *
    */
  covergroup trans_cross_axi_atomictype_bresp ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP
    axi_atomictype_bresp : cross write_xact_type, atomic_type,bresp{
      ignore_bins   ignore_excl_write_slverr_resp =  binsof(bresp.slverr_resp) || !binsof(atomic_type.exclusive) || !binsof(write_xact_type.write_xact);

      ignore_bins   ignore_excl_write_decerr_resp =    binsof(bresp.decerr_resp) || !binsof(atomic_type.exclusive) || !binsof(write_xact_type.write_xact);

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else 
 covergroup trans_cross_axi_atomictype_bresp_locked_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_LOCKED_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_atomictype_bresp : cross write_xact_type, atomic_type,bresp{
           option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_bresp_normal_axi3;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_LOCKED_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_atomictype_bresp : cross write_xact_type, atomic_type,bresp{
          option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_bresp_locked_exclusive_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_ALL
    axi_atomictype_bresp : cross write_xact_type, atomic_type,bresp{
           option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_bresp_exclusive_axi3_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_NOT_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_ALL
    axi_atomictype_bresp : cross write_xact_type, atomic_type,bresp{
           option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 covergroup trans_cross_axi_atomictype_bresp_exclusive_axi4lite ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_LOCKED_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_atomictype_bresp : cross write_xact_type, atomic_type,bresp{
          option.weight = 1;
    }
    option.per_instance = 1;
      endgroup
  covergroup trans_cross_axi_atomictype_bresp_normal_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_LOCKED_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_atomictype_bresp : cross write_xact_type, atomic_type,bresp{
         option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_atomictype_bresp_exclusive_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_NOT_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_ALL
    axi_atomictype_bresp : cross write_xact_type, atomic_type,bresp{
         option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`endif //  `ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

 /**
    * Covergroup: trans_cross_axi_read_interleaving_depth
    *
    * Coverpoints:
    *
    * - read_data_interleave : Captures read data interleave depth
    * .
    *
    */

   covergroup trans_cross_axi_read_interleaving_depth @(cov_interleave_depth_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_DATA_INTERLEAVE_DEPTH

    option.per_instance = 1;
  endgroup

 /**
    * Covergroup: trans_cross_axi4_stream_interleaving_depth
    *
    * Coverpoints:
    *
    * - axi4_stream_interleave : Captures axi4 stream data interleave depth
    * .
    *
    */

   covergroup trans_cross_axi4_stream_interleaving_depth @(cov_stream_interleave_depth_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_STREAM_DATA_INTERLEAVE_DEPTH

    option.per_instance = 1;
  endgroup
  /**
    * Covergroup: trans_cross_axi_ooo_read_response_depth
    *
    * Coverpoints:
    *
    * - ooo_read_response       : Captures out-of-order read response
    * - ooo_read_response_depth : Captures out-of-order read response depth
    *   - out-of-order response depth is determined by the position of the 
    *     transaction in outstanding queue for which response is being returned.
    *     Ex: if outstanding queue has 5 entries and response is received for 
    *         4th transaction (i.e. entry[3]) then depth will be determined as "3"
    *         because, response for the first or head-of-ooo-queue transaction is
    *         not considered as out-of-order.
    *   - User has option to modify each coverpoints through following defines.
    *     - VIP Built-in IGNORE_BIN define: VIP provides following "define" macro
    *       <b> `IGNORE_BINS_CG_trans_cross_axi_ooo_read_response_depth_CP_ooo_read_response </b> <br>
    *       <b> `IGNORE_BINS_CG_trans_cross_axi_ooo_read_response_depth_CP_ooo_read_response_depth </b> <br>
    *       _CG_ provides covergroup name and _CP_ provides coverpoint name. By default these are defined empty.
    *       User can just define above macros to ignore certain bin values or ignore all bins and
    *       define entirely customized set of bins.
    *       NOTE: ignore bin name is completely user defined, VIP doesn't have any restriction fo this.
    *     - user can override the covergroup by extending the callback class and re-defining this covergroup
    *     - user can disable this covergroup and define their own covergroup extending this coverage callback class
    *     .
    *   .
    * .
    *
    */
  covergroup trans_cross_axi_ooo_read_response_depth @(cov_out_of_order_read_response_depth_event);
   ooo_read_response: coverpoint out_of_order_read_response_depth iff(out_of_order_read_response_depth_flag){ 
      bins ooo_depth = {[0:((cfg.num_outstanding_xact == -1)?cfg.num_read_outstanding_xact-1:cfg.num_outstanding_xact-1)]}; 
      `IGNORE_BINS_CG_trans_cross_axi_ooo_read_response_depth_CP_ooo_read_response
      option.weight = 1; 
    }
    ooo_read_response_depth : coverpoint out_of_order_read_response_depth iff(out_of_order_read_response_depth_flag){ 
      bins ooo_depth[] = {[0:((cfg.num_outstanding_xact == -1)?cfg.num_read_outstanding_xact-1:cfg.num_outstanding_xact-1)]}; 
      `IGNORE_BINS_CG_trans_cross_axi_ooo_read_response_depth_CP_ooo_read_response_depth
      option.weight = 1; 
    }
    option.per_instance = 1; 
  endgroup


  /**
    * Covergroup: trans_cross_axi_ooo_write_response_depth
    *
    * Coverpoints:
    *
    * - ooo_write_response       : Captures out-of-order write response
    * - ooo_write_response_depth : Captures out-of-order write response depth
    *   - out-of-order response depth is determined by the position of the 
    *     transaction in outstanding queue for which response is being returned.
    *     Ex: if outstanding queue has 5 entries and response is received for 
    *         4th transaction (i.e. entry[3]) then depth will be determined as "3"
    *         because, response for the first or head-of-ooo-queue transaction is
    *         not considered as out-of-order.
    *   - User has option to modify each coverpoints through following defines.
    *     - VIP Built-in IGNORE_BIN define: VIP provides following "define" macro
    *       <b> `IGNORE_BINS_CG_trans_cross_axi_ooo_write_response_depth_CP_ooo_write_response </b> <br>
    *       <b> `IGNORE_BINS_CG_trans_cross_axi_ooo_write_response_depth_CP_ooo_write_response_depth </b> <br>
    *       _CG_ provides covergroup name and _CP_ provides coverpoint name. By default these are defined empty.
    *       User can just define above macros to ignore certain bin values or ignore all bins and
    *       define entirely customized set of bins.
    *       NOTE: ignore bin name is completely user defined, VIP doesn't have any restriction fo this.
    *     - user can override the covergroup by extending the callback class and re-defining this covergroup
    *     - user can disable this covergroup and define their own covergroup extending this coverage callback class
    *     .
    *   .
    * .
    *
    */
  covergroup trans_cross_axi_ooo_write_response_depth @(cov_out_of_order_write_response_depth_event);
   ooo_write_response: coverpoint out_of_order_write_response_depth iff(out_of_order_write_response_depth_flag){ 
      bins ooo_depth = {[0:((cfg.num_outstanding_xact == -1)?cfg.num_write_outstanding_xact-1:cfg.num_outstanding_xact-1)]}; 
      `IGNORE_BINS_CG_trans_cross_axi_ooo_write_response_depth_CP_ooo_write_response
      option.weight = 1; 
    }
    ooo_write_response_depth : coverpoint out_of_order_write_response_depth iff(out_of_order_write_response_depth_flag){ 
      bins ooo_depth[] = {[0:((cfg.num_outstanding_xact == -1)?cfg.num_write_outstanding_xact-1:cfg.num_outstanding_xact-1)]}; 
      `IGNORE_BINS_CG_trans_cross_axi_ooo_write_response_depth_CP_ooo_write_response_depth
      option.weight = 1; 
    }
    option.per_instance = 1; 
  endgroup

  /**
    * Covergroup: trans_cross_axi3_awburst_awlen_awsize
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - burst_size: Captures transaction burst size
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_awburst_awlen_awsize: Crosses cover points write_xact_type, burst_type, burst_length, burst_size
    * .
    *
    */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi3_awburst_awlen_awsize ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE
    axi3_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
   /**
    * Covergroup: trans_cross_axi4_awburst_awlen_awsize
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - burst_size: Captures transaction burst size
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_awburst_awlen_awsize: Crosses cover points write_xact_type, burst_type, burst_length, burst_size
    * .
    *
    */
  covergroup trans_cross_axi4_awburst_awlen_awsize ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE
    axi4_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi_awburst_awlen_awsize_axi3_dwlt_16bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi3_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi3_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi3_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi3_dwlt_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi3_dwlt_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi3_dwlt_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi3_dweq_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_dwlt_16bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_dwlt_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_dwlt_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_dwlt_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_dweq_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_ace_dwlt_16bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_ace_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_ace_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_ace_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_ace_dwlt_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_ace_dwlt_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_ace_dwlt_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_ace_dweq_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_lite_dwlt_16bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_lite_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_lite_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_lite_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_lite_dwlt_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_lite_dwlt_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_lite_dwlt_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awsize_axi4_lite_dweq_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    axi_awburst_awlen_awsize : cross write_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  
  /**
    * Covergroup: trans_cross_axi3_awburst_awlen_awlock
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - atomic_type: Captures transaction atomic type
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_awburst_awlen_awsize: Crosses cover points write_xact_type, burst_type, burst_length, atomic_type
    * .
    *
    */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF       
  covergroup trans_cross_axi3_awburst_awlen_awlock ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE
    axi3_awburst_awlen_awlock : cross write_xact_type, burst_type, burst_length, atomic_type {
      ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  /**
    * Covergroup: trans_cross_axi4_awburst_awlen_awlock
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - atomic_type: Captures transaction atomic type
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_awburst_awlen_awsize: Crosses cover points write_xact_type, burst_type, burst_length, atomic_type
    * .
    *
    */
  covergroup trans_cross_axi4_awburst_awlen_awlock ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE
    axi4_awburst_awlen_awlock : cross write_xact_type, burst_type, burst_length, atomic_type {
      ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

 `else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi_awburst_axi3_ace_awlen_axi3_awlock_locked_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_LOCKED_AXI3
    axi_awburst_awlen_arwock : cross write_xact_type, burst_type, burst_length, atomic_type{
      //ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

   covergroup trans_cross_axi_awburst_axi3_ace_awlen_axi3_awlock_no_locked_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_LOCKED_AXI3
    axi_awburst_awlen_arwock : cross write_xact_type, burst_type, burst_length, atomic_type{
      //ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_axi3_ace_awlen_axi3_awlock_exclusive_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_AXI3
    axi_awburst_awlen_arwock : cross write_xact_type, burst_type, burst_length, atomic_type{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_axi3_ace_awlen_axi3_awlock_no_exclusive_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_EXCLUSIVE_AXI3
    axi_awburst_awlen_awlock : cross write_xact_type, burst_type, burst_length, atomic_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_axi3_ace_awlen_axi4_awlock_exlusive_not_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_NOT_AXI3
    axi_awburst_awlen_awlock : cross write_xact_type, burst_type, burst_length, atomic_type{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_axi3_ace_awlen_axi4_awlock_no_exclusive_not_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_EXCLUSIVE_NOT_AXI3
    axi_awburst_awlen_awlock : cross write_xact_type, burst_type, burst_length, atomic_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_axi3_ace_awlen_ace_awlock_exclusive_not_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_NOT_AXI3
    axi_awburst_awlen_awlock : cross write_xact_type, burst_type, burst_length, atomic_type{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_axi3_ace_awlen_ace_awlock_no_exclusive_not_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_EXCLUSIVE_NOT_AXI3
    axi_awburst_awlen_awlock : cross write_xact_type, burst_type, burst_length, atomic_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_axi4_lite_awlen_axi4_lite_awlock_exclusive_not_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_NOT_AXI3
    axi_awburst_awlen_awlock : cross write_xact_type, burst_type, burst_length, atomic_type{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
 `endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_axi4_lite_awlen_axi4_lite_awlock_no_exclusive_not_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_EXCLUSIVE_NOT_AXI3
    axi_awburst_awlen_awlock : cross write_xact_type, burst_type, burst_length, atomic_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
 `endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
 
  /**
    * Covergroup: trans_cross_axi3_awburst_awlen_awaddr_awsize
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - addr: Captures min, mid and max range of transaction address
    * - burst_size: Captures transaction burst size
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_awburst_awlen_awaddr_awsize: Crosses cover points write_xact_type, burst_type, burst_length, addr, burst_size
    * .
    *
    */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF       
  covergroup trans_cross_axi3_awburst_awlen_awaddr_awsize ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE
    axi3_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 /**
    * Covergroup: trans_cross_axi4_awburst_awlen_awaddr_awsize
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - addr: Captures min, mid and max range of transaction address
    * - burst_size: Captures transaction burst size
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_awburst_awlen_awaddr_awsize: Crosses cover points write_xact_type, burst_type, burst_length, addr, burst_size
    * .
    *
    */
  covergroup trans_cross_axi4_awburst_awlen_awaddr_awsize ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE
    axi4_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
 
`else
  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi3_dwlt_16bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi3_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi3_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi3_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi3_dwlt_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi3_dwlt_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi3_dwlt_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi3_dweq_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi4_dwlt_16bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi4_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi4_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi4_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi4_dwlt_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi4_dwlt_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi4_dwlt_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi4_dweq_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_ace_dwlt_16bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_ace_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_ace_dwlt_64bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_ace_dwlt_128bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_ace_dwlt_256bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup  

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_ace_dwlt_512bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_ace_dwlt_1024bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_ace_dweq_1024bit;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1} ; 
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst); 
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif
  
  /**
    * Covergroup: trans_cross_axi3_awburst_awlen_awcache
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - cache_type: Captures transaction cache type
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_awburst_awlen_awcache: Crosses cover points write_xact_type, burst_type, burst_length, cache_type
    * .
    *
    */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi3_awburst_awlen_awcache ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE
    axi3_awburst_awlen_awcache : cross write_xact_type, burst_type, burst_length, cache_type {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
    /**
    * Covergroup: trans_cross_axi4_awburst_awlen_awcache
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - cache_type: Captures transaction cache type
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_awburst_awlen_awcache: Crosses cover points write_xact_type, burst_type, burst_length, cache_type
    * .
    *
    */
  covergroup trans_cross_axi4_awburst_awlen_awcache ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE
    axi4_awburst_awlen_awcache : cross write_xact_type, burst_type, burst_length, cache_type {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi_awburst_awlen_awcache_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE
    axi_awburst_awlen_awcache : cross write_xact_type, burst_type, burst_length, cache_type {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awcache_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4
    axi_awburst_awlen_awcache : cross write_xact_type, burst_type, burst_length, cache_type {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awcache_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4
    axi_awburst_awlen_awcache : cross write_xact_type, burst_type, burst_length, cache_type {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awcache_axi4_lite ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4
    axi_awburst_awlen_awcache : cross write_xact_type, burst_type, burst_length, cache_type {
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  
  /**
    * Covergroup: trans_cross_axi3_awburst_awlen_awprot
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - prot_type: Captures transaction protection type
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_awburst_awlen_awprot: Crosses cover points write_xact_type, burst_type, burst_length, prot_type
    * .
    *
    */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi3_awburst_awlen_awprot ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE
    axi3_awburst_awlen_awprot : cross write_xact_type, burst_type, burst_length, prot_type {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  /**
    * Covergroup: trans_cross_axi4_awburst_awlen_awprot
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - prot_type: Captures transaction protection type
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_awburst_awlen_awprot: Crosses cover points write_xact_type, burst_type, burst_length, prot_type
    * .
    *
    */
  covergroup trans_cross_axi4_awburst_awlen_awprot ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE
    axi4_awburst_awlen_awprot : cross write_xact_type, burst_type, burst_length, prot_type {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else

  covergroup trans_cross_axi_awburst_awlen_awprot_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE
    axi_awburst_awlen_awprot : cross write_xact_type, burst_type, burst_length, prot_type {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_awburst_awlen_awprot_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE
    axi_awburst_awlen_awprot : cross write_xact_type, burst_type, burst_length, prot_type {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_awburst_awlen_awprot_axi4_lite ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE
    axi_awburst_awlen_awprot : cross write_xact_type, burst_type, burst_length, prot_type {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_awburst_awlen_awprot_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE
    axi_awburst_awlen_awprot : cross write_xact_type, burst_type, burst_length, prot_type {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  `endif


  /**
    * Covergroup: trans_cross_axi_write_strobes
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - wstrb: Captures write strobe values
    * .
    *
    * Cross coverpoints:
    *
    * - axi_write_strobes: Crosses cover points write_xact_type,wstrb
    * .
    *
    */ 
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF       
  covergroup trans_cross_axi_write_strobes ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WSTRB

    axi_write_strobes : cross write_xact_type,wstrb {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi_write_strobes_dwlt_32 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WSTRB_DWLT_32

    axi_write_strobes : cross write_xact_type,wstrb {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_strobes_dwlt_64 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WSTRB_DWLT_64

    axi_write_strobes : cross write_xact_type,wstrb {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_strobes_dwlt_128 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WSTRB_DWLT_128

    axi_write_strobes : cross write_xact_type,wstrb {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_strobes_dwlt_256 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WSTRB_DWLT_256

    axi_write_strobes : cross write_xact_type,wstrb {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_strobes_dwlt_512 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WSTRB_DWLT_512

    axi_write_strobes : cross write_xact_type,wstrb {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_strobes_dwlt_1024 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WSTRB_DWLT_1024

    axi_write_strobes : cross write_xact_type,wstrb {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_strobes_dweq_1024 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WSTRB_DWEQ_1024

    axi_write_strobes : cross write_xact_type,wstrb {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  /**
    * Covergroup: trans_cross_axi_write_narrow_transfer_awlen_awaddr
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - transfer_size: Captures transaction burst size
    * - addr_offset: Captures transaction address offset information
    * .
    *
    * Cross coverpoints:
    *
    * - axi_write_narrow_transfer_awlen_awaddr: Crosses cover points write_xact_type,transfer_size,addr_offset
    * .
    *
    */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF       
  covergroup trans_cross_axi_write_narrow_transfer_awlen_awaddr ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET
    

    axi_write_narrow_transfer_awlen_awaddr : cross write_xact_type,transfer_size,addr_offset {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_0_TO_F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_10_TO_1F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_20_TO_2F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_30_TO_3F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_40_TO_4F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_50_TO_5F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_60_TO_6F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_70_TO_7F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COMMON_IGNORE_BINS
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else // SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi_write_narrow_transfer_awlen_awaddr_axi3_dweq_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    axi_write_narrow_transfer_awlen_awaddr_axi3_dweq_32bit : cross write_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup 

  covergroup trans_cross_axi_write_narrow_transfer_awlen_awaddr_axi3_dweq_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    axi_write_narrow_transfer_awlen_awaddr_axi3_dweq_64bit : cross write_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_narrow_transfer_awlen_awaddr_axi3_dweq_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    axi_write_narrow_transfer_awlen_awaddr_axi3_dweq_128bit : cross write_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_narrow_transfer_awlen_awaddr_axi3_dweq_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_512
    axi_write_narrow_transfer_awlen_awaddr_axi3_dweq_256bit : cross write_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_narrow_transfer_awlen_awaddr_axi3_dweq_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_512
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_1024
    axi_write_narrow_transfer_awlen_awaddr_axi3_dweq_512bit : cross write_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_narrow_transfer_awlen_awaddr_axi4_dweq_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    axi_write_narrow_transfer_awlen_awaddr_axi4_dweq_32bit : cross write_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup 

  covergroup trans_cross_axi_write_narrow_transfer_awlen_awaddr_axi4_dweq_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    axi_write_narrow_transfer_awlen_awaddr_axi4_dweq_64bit : cross write_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_narrow_transfer_awlen_awaddr_axi4_dweq_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    axi_write_narrow_transfer_awlen_awaddr_axi4_dweq_128bit : cross write_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_narrow_transfer_awlen_awaddr_ace_dweq_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    axi_write_narrow_transfer_awlen_awaddr_ace_dweq_32bit : cross write_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup 

  covergroup trans_cross_axi_write_narrow_transfer_awlen_awaddr_ace_dweq_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    axi_write_narrow_transfer_awlen_awaddr_ace_dweq_64bit : cross write_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_narrow_transfer_awlen_awaddr_ace_dweq_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    axi_write_narrow_transfer_awlen_awaddr_ace_dweq_128bit : cross write_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_narrow_transfer_awlen_awaddr_ace_dweq_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_512
    axi_write_narrow_transfer_awlen_awaddr_ace_dweq_256bit : cross write_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_write_narrow_transfer_awlen_awaddr_ace_dweq_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_512
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_1024
    axi_write_narrow_transfer_awlen_awaddr_ace_dweq_512bit : cross write_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`endif // SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  /**
    * Covergroup: trans_cross_axi_write_unaligned_transfer
    *
    * Coverpoints:
    *
    * - write_xact_type:  Captures write transaction
    * - burst_type: Captures transaction burst type
    * - addr_offset: Captures transaction address offset information
    * - transfer_size: Captures transaction burst size
    * - burst_length: Captures transaction burst length
    * .
    *
    * Cross coverpoints:
    *
    * - axi_write_unaligned_transfer: Crosses cover points write_xact_type, burst_type, addr_offset, transfer_size, burst_length
    * .
    *
    */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF       
  covergroup trans_cross_axi_write_unaligned_transfer ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH 

    axi_write_unaligned_transfer : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
covergroup trans_cross_axi_write_unaligned_transfer_axi3_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3

    axi_write_unaligned_transfer : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_write_unaligned_transfer_axi3_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3

    axi_write_unaligned_transfer : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_write_unaligned_transfer_axi3_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3

    axi_write_unaligned_transfer : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_write_unaligned_transfer_axi4_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4

    axi_write_unaligned_transfer : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_write_unaligned_transfer_axi4_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4

    axi_write_unaligned_transfer : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_write_unaligned_transfer_axi4_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4

    axi_write_unaligned_transfer : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

covergroup trans_cross_axi_write_unaligned_transfer_ace_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE

    axi_write_unaligned_transfer : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

covergroup trans_cross_axi_write_unaligned_transfer_ace_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE

    axi_write_unaligned_transfer : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_write_unaligned_transfer_ace_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE

    axi_write_unaligned_transfer : cross write_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  
  /**
    * Covergroup: trans_cross_axi3_arburst_arlen
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_arburst_arlen: Crosses cover points read_xact_type, burst_type and burst_length
    * .
    *
    */
  //covergroup trans_cross_axi_arburst_arlen @(cov_read_sample_event);
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF       
  covergroup trans_cross_axi3_arburst_arlen ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    axi3_arburst_arlen : cross read_xact_type, burst_type, burst_length {
    `ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
    `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
/**
    * Covergroup: trans_cross_axi4_arburst_arlen
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_arburst_arlen: Crosses cover points read_xact_type, burst_type and burst_length
    * .
    *
    */
  covergroup trans_cross_axi4_arburst_arlen ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
    axi4_arburst_arlen : cross read_xact_type, burst_type, burst_length {
    `ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
    `endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else
  covergroup trans_cross_axi_arburst_arlen_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    axi_arburst_arlen : cross read_xact_type, burst_type, burst_length {
    `ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
    `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    axi_arburst_arlen : cross read_xact_type, burst_type, burst_length {
    `ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
    `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_axi4_lite ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    axi_arburst_arlen : cross read_xact_type, burst_type, burst_length {
    //`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
    //  ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
    //`endif
    //  ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    axi_arburst_arlen : cross read_xact_type, burst_type, burst_length {
    `ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
    `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`endif

  /**
    * Covergroup: trans_cross_axi3_arburst_arlen_araddr
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - addr: Captures min, mid and max range of transaction address
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_arburst_arlen_araddr: Crosses cover points read_xact_type, burst_type, burst_length, addr
    * .
    *
    */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF       
  //covergroup trans_cross_axi3_arburst_arlen_araddr @(cov_read_sample_event);
  covergroup trans_cross_axi3_arburst_arlen_araddr ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR
    axi3_arburst_arlen_araddr : cross read_xact_type, burst_type, burst_length, addr {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif     
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  /**
    * Covergroup: trans_cross_axi4_arburst_arlen_araddr
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - addr: Captures min, mid and max range of transaction address
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_arburst_arlen_araddr: Crosses cover points read_xact_type, burst_type, burst_length, addr
    * .
    *
    */
  //covergroup trans_cross_axi4_arburst_arlen_araddr @(cov_read_sample_event);
  covergroup trans_cross_axi4_arburst_arlen_araddr ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR
    axi4_arburst_arlen_araddr : cross read_xact_type, burst_type, burst_length, addr {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif     
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  covergroup trans_cross_axi_arburst_axi3_ace_arlen_axi3_araddr_axi3_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4 
    axi_arburst_arlen_araddr : cross read_xact_type, burst_type, burst_length, addr {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif     
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_axi3_ace_arlen_axi4_araddr_axi3_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    axi_arburst_arlen_araddr : cross read_xact_type, burst_type, burst_length, addr {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif     
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_axi_arburst_axi3_ace_arlen_ace_araddr_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    axi_arburst_arlen_araddr : cross read_xact_type, burst_type, burst_length, addr {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif     
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_axi_arburst_axi4_lite_arlen_axi4_lite_araddr_axi3_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    axi_arburst_arlen_araddr : cross read_xact_type, burst_type, burst_length, addr {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
 `endif
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};
`endif     
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF 
    
  /**
    * Covergroup: trans_cross_axi3_arburst_arlen_rresp
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - rresp: Captures transaction response
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_arburst_arlen_rresp: Crosses cover points read_xact_type, burst_type, burst_length, rresp
    * .
    *
    */
  //covergroup trans_cross_axi3_arburst_arlen_rresp @(cov_read_sample_event);
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF   
  covergroup trans_cross_axi3_arburst_arlen_rresp ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP
    axi3_arburst_arlen_rresp : cross read_xact_type, burst_type, burst_length, rresp{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(rresp.exokay_resp) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
/**
    * Covergroup: trans_cross_axi4_arburst_arlen_rresp
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - rresp: Captures transaction response
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_arburst_arlen_rresp: Crosses cover points read_xact_type, burst_type, burst_length, rresp
    * .
    *
    */
  //covergroup trans_cross_axi4_arburst_arlen_rresp @(cov_read_sample_event);
  covergroup trans_cross_axi4_arburst_arlen_rresp ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP
    axi4_arburst_arlen_rresp : cross read_xact_type, burst_type, burst_length, rresp{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(rresp.exokay_resp) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  covergroup trans_cross_axi_arburst_axi3_ace_arlen_axi3_rresp_no_exclusive ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_arburst_arlen_rresp : cross read_xact_type, burst_type, burst_length, rresp{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_arburst_axi3_ace_arlen_axi3_rresp_all ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_ALL
    axi_arburst_arlen_rresp : cross read_xact_type, burst_type, burst_length, rresp{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(rresp.exokay_resp) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_arburst_axi3_ace_arlen_axi4_rresp_no_exclusive ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_arburst_arlen_rresp : cross read_xact_type, burst_type, burst_length, rresp{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_axi3_ace_arlen_axi4_rresp_all ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_ALL
    axi_arburst_arlen_rresp : cross read_xact_type, burst_type, burst_length, rresp{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(rresp.exokay_resp) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_arburst_axi3_ace_arlen_ace_rresp_no_exclusive ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_arburst_arlen_rresp : cross read_xact_type, burst_type, burst_length, rresp{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_arburst_axi3_ace_arlen_ace_rresp_all ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_ALL
    axi_arburst_arlen_rresp : cross read_xact_type, burst_type, burst_length, rresp{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(rresp.exokay_resp) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_arburst_axi4_lite_arlen_axi4_lite_rresp_no_exclusive ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_NO_EXCLUSIVE_AXI4_LITE
    axi_arburst_arlen_rresp : cross read_xact_type, burst_type, burst_length, rresp{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
 `endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_arburst_axi4_lite_arlen_axi4_lite_rresp_all ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_RRESP_ALL
    axi_arburst_arlen_rresp : cross read_xact_type, burst_type, burst_length, rresp{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(rresp.exokay_resp) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
 `endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  
  /**
    * Covergroup: trans_cross_axi3_arburst_arlen_arsize
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - burst_size: Captures transaction burst size
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_arburst_arlen_arsize: Crosses cover points read_xact_type, burst_type, burst_length, burst_size
    * .
    *
    */
  //covergroup trans_cross_axi3_arburst_arlen_arsize @(cov_read_sample_event);
  `ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi3_arburst_arlen_arsize ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE
    axi3_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
/**
    * Covergroup: trans_cross_axi4_arburst_arlen_arsize
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - burst_size: Captures transaction burst size
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_arburst_arlen_arsize: Crosses cover points read_xact_type, burst_type, burst_length, burst_size
    * .
    *
    */
  //covergroup trans_cross_axi4_arburst_arlen_arsize @(cov_read_sample_event);
   covergroup trans_cross_axi4_arburst_arlen_arsize ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE
    axi4_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  `else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi_arburst_arlen_arsize_axi3_dwlt_16bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi3_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi3_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi3_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi3_dwlt_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi3_dwlt_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi3_dwlt_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi3_dweq_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_dwlt_16bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_dwlt_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_dwlt_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_dwlt_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_dweq_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_ace_dwlt_16bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_ace_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_ace_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_ace_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_ace_dwlt_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_ace_dwlt_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_ace_dwlt_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_ace_dweq_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_lite_dwlt_16bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_lite_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_lite_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_lite_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_lite_dwlt_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_lite_dwlt_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_lite_dwlt_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arsize_axi4_lite_dweq_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    axi_arburst_arlen_arsize : cross read_xact_type, burst_type, burst_length, burst_size{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  `endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
    
  /**
    * Covergroup: trans_cross_axi3_arburst_arlen_araddr_arsize
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - addr: Captures min, mid and max range of transaction address
    * - burst_size: Captures transaction burst size
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_arburst_arlen_araddr_arsize: Crosses cover points read_xact_type, burst_type, burst_length, addr, burst_size
    * .
    *
    */
  //covergroup trans_cross_axi3_arburst_arlen_araddr_arsize @(cov_read_sample_event);
  `ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi3_arburst_arlen_araddr_arsize ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE
    axi3_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  /**
    * Covergroup: trans_cross_axi4_arburst_arlen_araddr_arsize
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - addr: Captures min, mid and max range of transaction address
    * - burst_size: Captures transaction burst size
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_arburst_arlen_araddr_arsize: Crosses cover points read_xact_type, burst_type, burst_length, addr, burst_size
    * .
    *
    */
  //covergroup trans_cross_axi4_arburst_arlen_araddr_arsize @(cov_read_sample_event);
  covergroup trans_cross_axi4_arburst_arlen_araddr_arsize ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE
    axi4_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  `else
  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi3_dwlt_16bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi3_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi3_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi3_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup  

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi3_dwlt_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

    covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi3_dwlt_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

    covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi3_dwlt_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

    covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi3_dweq_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi4_dwlt_16bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi4_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi4_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi4_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi4_dwlt_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi4_dwlt_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi4_dwlt_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi4_dweq_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_ace_dwlt_16bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_ace_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_ace_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_ace_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_ace_dwlt_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_ace_dwlt_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_ace_dwlt_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_ace_dweq_1024bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
`ifdef SVT_MULTI_SIM_COVPOINT_GREATER_THAN_32_BITS
      // Need to compe up with an alternative
`else
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      ignore_bins Ignore_invalid_max_addr_wrap_burst = binsof(addr.addr_range_max) && binsof(burst_type.wrap_burst);
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif

  /**
    * Covergroup: trans_cross_axi_arburst_arlen_araddr_arsize_axi4_lite
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - addr: Captures min, mid and max range of transaction address
    * - burst_size: Captures transaction burst size
    * .
    *
    * Cross coverpoints:
    *
    * - axi_arburst_arlen_araddr_arsize: Crosses cover points read_xact_type, burst_type, burst_length, addr, burst_size
    * .
    *
    */
`ifdef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi4_lite_dweq_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_32BIT_AXI4_LITE
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_araddr_arsize_axi4_lite_dweq_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_64BIT_AXI4_LITE
    axi_arburst_arlen_araddr_arsize : cross read_xact_type, burst_type, burst_length, addr, burst_size {
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup


  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi4_lite_dweq_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_32BIT_AXI4_LITE
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_awburst_awlen_awaddr_awsize_axi4_lite_dweq_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WRITE_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_AXI3_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_64BIT_AXI4_LITE
    axi_awburst_awlen_awaddr_awsize : cross write_xact_type, burst_type, burst_length, addr, burst_size {
      ignore_bins Ignore_invalid_max_addr_incr_burst_length = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_length) intersect {1};  
      ignore_bins Ignore_invalid_max_addr_incr_burst_size = binsof(addr.addr_range_max) && binsof(burst_type.incr_burst) && !binsof(burst_size) intersect {`SVT_AXI_TRANSACTION_BURST_SIZE_8}; 
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup


`endif

  
  /**
    * Covergroup: trans_cross_axi3_arburst_arlen_arlock
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - atomic_type: Captures transaction atomic type
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_arburst_arlen_arlock: Crosses cover points read_xact_type, burst_type, burst_length, atomic_type
    * .
    *
    */
  //covergroup trans_cross_axi3_arburst_arlen_arlock @(cov_read_sample_event);

`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF   
  covergroup trans_cross_axi3_arburst_arlen_arlock ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE
    axi3_arburst_arlen_arlock : cross read_xact_type, burst_type, burst_length, atomic_type{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  /**
    * Covergroup: trans_cross_axi4_arburst_arlen_arlock
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - atomic_type: Captures transaction atomic type
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_arburst_arlen_arlock: Crosses cover points read_xact_type, burst_type, burst_length, atomic_type
    * .
    *
    */
  //covergroup trans_cross_axi4_arburst_arlen_arlock @(cov_read_sample_event);

  covergroup trans_cross_axi4_arburst_arlen_arlock ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE
    axi4_arburst_arlen_arlock : cross read_xact_type, burst_type, burst_length, atomic_type{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi_arburst_axi3_ace_arlen_axi3_arlock_locked_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_LOCKED_AXI3
    axi_arburst_arlen_arlock : cross read_xact_type, burst_type, burst_length, atomic_type{
    //  ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_axi_arburst_axi3_ace_arlen_axi3_arlock_no_locked_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_LOCKED_AXI3
    axi_arburst_arlen_arlock : cross read_xact_type, burst_type, burst_length, atomic_type{
    //  ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};   
 `ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_axi3_ace_arlen_axi3_arlock_exclusive_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_AXI3
    axi_arburst_arlen_arlock : cross read_xact_type, burst_type, burst_length, atomic_type{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_axi3_ace_arlen_axi3_arlock_no_exclusive_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_EXCLUSIVE_AXI3
    axi_arburst_arlen_arlock : cross read_xact_type, burst_type, burst_length, atomic_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_axi3_ace_arlen_axi4_arlock_exlusive_not_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_NOT_AXI3
    axi_arburst_arlen_arlock : cross read_xact_type, burst_type, burst_length, atomic_type{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_axi3_ace_arlen_axi4_arlock_no_exclusive_not_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_EXCLUSIVE_NOT_AXI3
    axi_arburst_arlen_arlock : cross read_xact_type, burst_type, burst_length, atomic_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_axi3_ace_arlen_ace_arlock_exclusive_not_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_NOT_AXI3
    axi_arburst_arlen_arlock : cross read_xact_type, burst_type, burst_length, atomic_type{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_axi3_ace_arlen_ace_arlock_no_exclusive_not_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_EXCLUSIVE_NOT_AXI3
    axi_arburst_arlen_arlock : cross read_xact_type, burst_type, burst_length, atomic_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_axi4_lite_arlen_axi4_lite_arlock_exclusive_not_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_EXCLUSIVE_NOT_AXI3
    axi_arburst_arlen_arlock : cross read_xact_type, burst_type, burst_length, atomic_type{
      ignore_bins Ignore_invalid_excl_burst   =  binsof(atomic_type.exclusive) && !binsof(burst_length) intersect {1,`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
 `endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_axi4_lite_arlen_axi4_lite_arlock_no_exclusive_not_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ATOMIC_TYPE_NO_EXCLUSIVE_NOT_AXI3
    axi_arburst_arlen_arlock : cross read_xact_type, burst_type, burst_length, atomic_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
 `endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
    
  /**
    * Covergroup: trans_cross_axi_arburst_arlen_arcache
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - cache_type: Captures transaction cache type
    * .
    *
    * Cross coverpoints:
    *
    * - axi_arburst_arlen_arcache: Crosses cover points read_xact_type, burst_type, burst_length, cache_type
    * .
    *
    */
  //covergroup trans_cross_axi_arburst_arlen_arcache @(cov_read_sample_event);
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF       
  covergroup trans_cross_axi_arburst_arlen_arcache ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE
    axi_arburst_arlen_arcache : cross read_xact_type, burst_type, burst_length, cache_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi_arburst_arlen_arcache_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_CACHE_TYPE
    axi_arburst_arlen_arcache : cross read_xact_type, burst_type, burst_length, cache_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arcache_axi4 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4
    axi_arburst_arlen_arcache : cross read_xact_type, burst_type, burst_length, cache_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arcache_axi4_lite ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4
    axi_arburst_arlen_arcache : cross read_xact_type, burst_type, burst_length, cache_type{
//`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
//      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
//`endif
//      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arcache_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4
    axi_arburst_arlen_arcache : cross read_xact_type, burst_type, burst_length, cache_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
    
  /**
    * Covergroup: trans_cross_axi3_arburst_arlen_arprot
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - prot_type: Captures transaction protection type
    * .
    *
    * Cross coverpoints:
    *
    * - axi3_arburst_arlen_arprot: Crosses cover points read_xact_type, burst_type, burst_length, prot_type
    * .
    *
    */
  //covergroup trans_cross_axi3_arburst_arlen_arprot @(cov_read_sample_event);
  `ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  
  covergroup trans_cross_axi3_arburst_arlen_arprot ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI3_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE
    axi3_arburst_arlen_arprot : cross read_xact_type, burst_type, burst_length, prot_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
/**
    * Covergroup: trans_cross_axi4_arburst_arlen_arprot
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - burst_length: Captures transaction burst length
    * - prot_type: Captures transaction protection type
    * .
    *
    * Cross coverpoints:
    *
    * - axi4_arburst_arlen_arprot: Crosses cover points read_xact_type, burst_type, burst_length, prot_type
    * .
    *
    */
  //covergroup trans_cross_axi4_arburst_arlen_arprot @(cov_read_sample_event);
   
  covergroup trans_cross_axi4_arburst_arlen_arprot ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AXI4_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE
    axi4_arburst_arlen_arprot : cross read_xact_type, burst_type, burst_length, prot_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_wrap_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::WRAP} &&  !binsof(burst_length) intersect {[1:16]};
      ignore_bins Ignore_invalid_fixed_burst_type  =  binsof(burst_type) intersect {svt_axi_transaction::FIXED} && !binsof(burst_length) intersect {[1:16]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else

  covergroup trans_cross_axi_arburst_arlen_arprot_axi3 ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE
    axi_arburst_arlen_arprot : cross read_xact_type, burst_type, burst_length, prot_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arprot_axi4;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE
    axi_arburst_arlen_arprot : cross read_xact_type, burst_type, burst_length, prot_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_axi_arburst_arlen_arprot_axi4_lite ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE
    axi_arburst_arlen_arprot : cross read_xact_type, burst_type, burst_length, prot_type{
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_arburst_arlen_arprot_ace ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_PROT_TYPE
    axi_arburst_arlen_arprot : cross read_xact_type, burst_type, burst_length, prot_type{
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) && !binsof(burst_length) intersect {`SVT_AXI_WRAP_BURST_LENGTH_RANGE};
 `endif
      ignore_bins Ignore_invalid_fixed  =  binsof(burst_type.fixed_burst) && binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif

  /**
    * Covergroup: trans_cross_axi_read_narrow_transfer_arlen_araddr
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - transfer_size: Captures transaction burst size
    * - addr_offset: Captures transaction address offset information
    * .
    *
    * Cross coverpoints:
    *
    * - axi_read_narrow_transfer_arlen_araddr: Crosses cover points read_xact_type,transfer_size,addr_offset
    * .
    *
    */
  //covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr @(cov_read_sample_event);
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF       
  covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET 

    axi_read_narrow_transfer_arlen_araddr : cross read_xact_type,transfer_size,addr_offset  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_0_TO_F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_10_TO_1F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_20_TO_2F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_30_TO_3F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_40_TO_4F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_50_TO_5F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_60_TO_6F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_OFFSET_70_TO_7F_IGNORE_BINS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COMMON_IGNORE_BINS
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else // SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr_axi3_dweq_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    axi_read_narrow_transfer_arlen_araddr_axi3_dweq_32bit : cross read_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup 

  covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr_axi3_dweq_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    axi_read_narrow_transfer_arlen_araddr_axi3_dweq_64bit : cross read_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr_axi3_dweq_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    axi_read_narrow_transfer_arlen_araddr_axi3_dweq_128bit : cross read_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr_axi3_dweq_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_512
    axi_read_narrow_transfer_arlen_araddr_axi3_dweq_256bit : cross read_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr_axi3_dweq_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_512
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_1024
    axi_read_narrow_transfer_arlen_araddr_axi3_dweq_512bit : cross read_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr_axi4_dweq_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    axi_read_narrow_transfer_arlen_araddr_axi4_dweq_32bit : cross read_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup 

  covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr_axi4_dweq_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    axi_read_narrow_transfer_arlen_araddr_axi4_dweq_64bit : cross read_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr_axi4_dweq_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    axi_read_narrow_transfer_arlen_araddr_axi4_dweq_128bit : cross read_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr_ace_dweq_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    axi_read_narrow_transfer_arlen_araddr_ace_dweq_32bit : cross read_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup 

  covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr_ace_dweq_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    axi_read_narrow_transfer_arlen_araddr_ace_dweq_64bit : cross read_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr_ace_dweq_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    axi_read_narrow_transfer_arlen_araddr_ace_dweq_128bit : cross read_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr_ace_dweq_256bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_512
    axi_read_narrow_transfer_arlen_araddr_ace_dweq_256bit : cross read_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_axi_read_narrow_transfer_arlen_araddr_ace_dweq_512bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_512
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_1024
    axi_read_narrow_transfer_arlen_araddr_ace_dweq_512bit : cross read_xact_type,transfer_size,addr_offset {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`endif // SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  /**
    * Covergroup: trans_cross_axi_read_unaligned_transfer
    *
    * Coverpoints:
    *
    * - read_xact_type:  Captures read transaction
    * - burst_type: Captures transaction burst type
    * - addr_offset: Captures transaction address offset information
    * - transfer_size: Captures transaction burst size
    * - burst_length: Captures transaction burst length
    * .
    *
    * Cross coverpoints:
    *
    * - axi_read_unaligned_transfer: Crosses cover points read_xact_type, burst_type, addr_offset, transfer_size, burst_length
    * .
    *
    */
  //covergroup trans_cross_axi_read_unaligned_transfer @(cov_read_sample_event);
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF   
  covergroup trans_cross_axi_read_unaligned_transfer ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH 

    axi_read_unaligned_transfer : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else // SVT_AXI_MON_CFG_BASED_COV_GRP_DEF 
//this is resulting in 280 new CGs, so need to check for an alternative
covergroup trans_cross_axi_read_unaligned_transfer_axi3_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3

    axi_read_unaligned_transfer : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_read_unaligned_transfer_axi3_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3

    axi_read_unaligned_transfer : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_read_unaligned_transfer_axi3_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI3

    axi_read_unaligned_transfer : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_read_unaligned_transfer_axi4_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4

    axi_read_unaligned_transfer : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_read_unaligned_transfer_axi4_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4

    axi_read_unaligned_transfer : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_read_unaligned_transfer_axi4_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_AXI3
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_AXI4

    axi_read_unaligned_transfer : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

covergroup trans_cross_axi_read_unaligned_transfer_ace_dwlt_32bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_32 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_64
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE

    axi_read_unaligned_transfer : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

covergroup trans_cross_axi_read_unaligned_transfer_ace_dwlt_64bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_64 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE

    axi_read_unaligned_transfer : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
covergroup trans_cross_axi_read_unaligned_transfer_ace_dwlt_128bit ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_READ_XACT_TYPE_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_OFFSET_DWEQ_128
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_TRANSFER_SIZE_DWLT_256
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE

    axi_read_unaligned_transfer : cross read_xact_type, burst_type, addr_offset, transfer_size, burst_length  {

    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_INVALID_UNALIGNED_TRANSFER_CROSS_DW_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_4KB_BOUNDARY_CROSS

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif // SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  // ****************************************************************************
  // Delay Covergroups
  // ****************************************************************************

  /**
    *  Covergroup: trans_meta_axi_write
    *
    *  Coverpoints:
    *  - AWVALID_to_AWREADY_Delay: Captures min, mid and max range of delays between signals awvalid and awready
    *  - WVALID_to_WREADY_Delay: Captures min, mid and max range of delays between signals wvalid and wready
    *  - BVALID_to_BWREADY_Delay: Captures min, mid and max range of delays between signals bvalid and bready
    *  - AWVALID_to_prev_AWVALID_Delay: Captures min, mid and max range of delays between current and previous awvalid signals
    *  - WVALID_to_prev_WVALID_Delay: Captures min, mid and max range of delays between current and previous wvalid signals
    *  - AWVALID_to_first_WVALID_Delay: Captures min, mid and max range of delays between awvalid and first wvalid signals
    *  - last_wdata_handshake_to_BVALID_Delay: Captures min, mid and max range of delays between last write data handshake to bvalid signals
    *  - AWVALID_before_AWREADY: Captures if AWVALID signal comes before AWREADY signal 
    *  - AWREADY_before_AWVALID: Captures if AWREADY signal comes before AWVALID signal
    *  - BVALID_before_BREADY: Captures if BVALID signal comes before BREADY signal 
    *  - BREADY_before_BVALID: Captures if BREADY signal comes before BVALID signal
    *  - WVALID_before_WREADY: Captures if WVALID signal comes before WREADY signal 
    *  - WREADY_before_WVALID: Captures if WREADY signal comes before WVALID signal or WREADY,WVALID signals are comes at same time
    *  - AWVALID_before_WREADY: Captures if AWVALID signal comes before WREADY signal 
    *  - WREADY_before_AWVALID: Captures if WREADY signal comes before AWVALID signal
    *  - AWREADY_before_WVALID: Captures if AWREADY signal comes before WVALID signal 
    *  - WVALID_before_AWREADY: Captures if WVALID signal comes before AWREADY signal
    *  - AWVALID_before_WVALID: Captures if AWVALID signal comes before WVALID signal 
    *  - WVALID_before_AWVALID: Captures if WVALID signal comes before AWVALID signal
    *  .
    */  
  covergroup trans_meta_axi_write ;
    option.per_instance = 1;
    AWVALID_to_AWREADY_Delay : coverpoint cov_AWVALID_to_AWREADY_Delay {
      bins awvalid_to_awready_delay_min = {0};
      bins awvalid_to_awready_delay_mid = {[1:(`SVT_AXI_MAX_ADDR_DELAY/2)]};
      bins awvalid_to_awready_delay_max = {[(`SVT_AXI_MAX_ADDR_DELAY/2)+1:$]};
      option.at_least = `SVT_AXI_trans_meta_axi_write_AWVALID_to_AWREADY_Delay_COV_OPTION_AT_LEAST_VAL;
    }
    WVALID_to_WREADY_Delay : coverpoint cov_WVALID_to_WREADY_Delay {
      bins wvalid_to_wready_delay_min = {0};
      bins wvalid_to_wready_delay_mid = {[1:(`SVT_AXI_MAX_WREADY_DELAY/2)]};
      bins wvalid_to_wready_delay_max = {[(`SVT_AXI_MAX_WREADY_DELAY/2)+1:$]};
      option.at_least = `SVT_AXI_trans_meta_axi_write_WVALID_to_WREADY_Delay_COV_OPTION_AT_LEAST_VAL;
    }
    BVALID_to_BREADY_Delay : coverpoint cov_BVALID_to_BREADY_Delay {
      bins bvalid_to_bready_delay_min = {0};
      bins bvalid_to_bready_delay_mid = {[1:(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)]};
      bins bvalid_to_bready_delay_max = {[(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)+1:$]};
      option.at_least = `SVT_AXI_trans_meta_axi_write_BVALID_to_BREADY_Delay_COV_OPTION_AT_LEAST_VAL;
    }
    AWVALID_to_prev_AWVALID_Delay : coverpoint cov_AWVALID_to_prev_AWVALID_Delay {
      bins awvalid_to_prev_awvalid_delay_min = {1};
      bins awvalid_to_prev_awvalid_delay_mid = {[2:((`SVT_AXI_MAX_ADDR_VALID_DELAY + `SVT_AXI_MAX_ADDR_DELAY)/2)]};
      bins awvalid_to_prev_awvalid_delay_max = {[((`SVT_AXI_MAX_ADDR_VALID_DELAY + `SVT_AXI_MAX_ADDR_DELAY)/2)+1:$]};
      option.at_least = `SVT_AXI_trans_meta_axi_write_AWVALID_to_prev_AWVALID_Delay_COV_OPTION_AT_LEAST_VAL;
    } 
    WVALID_to_prev_WVALID_Delay : coverpoint cov_WVALID_to_prev_WVALID_Delay {
      bins wvalid_to_prev_wvalid_delay_min = {1};
      bins wvalid_to_prev_wvalid_delay_mid = {[2:((`SVT_AXI_MAX_WVALID_DELAY + `SVT_AXI_MAX_WREADY_DELAY)/2)]};
      bins wvalid_to_prev_wvalid_delay_max = {[((`SVT_AXI_MAX_WVALID_DELAY +  `SVT_AXI_MAX_WREADY_DELAY)/2)+1:$]};
      option.at_least = `SVT_AXI_trans_meta_axi_write_WVALID_to_prev_WVALID_Delay_COV_OPTION_AT_LEAST_VAL;
    } 
    AWVALID_to_first_WVALID_Delay : coverpoint cov_AWVALID_to_first_WVALID_Delay {
      bins awvalid_to_first_wvalid_delay_min = {0}; 
      bins awvalid_to_first_wvalid_delay_mid = {[1:((`SVT_AXI_MAX_ADDR_DELAY + `SVT_AXI_MAX_WVALID_DELAY)/2)]};
      bins awvalid_to_first_wvalid_delay_max = {[((`SVT_AXI_MAX_ADDR_DELAY + `SVT_AXI_MAX_WVALID_DELAY)/2)+1:$]}; 
      option.at_least = `SVT_AXI_trans_meta_axi_write_AWVALID_to_first_WVALID_Delay_COV_OPTION_AT_LEAST_VAL;
    } 
    last_wdata_handshake_to_BVALID_Delay : coverpoint cov_last_wdata_handshake_to_BVALID_Delay {
      bins last_wdata_handshake_to_bvalid_delay_min = {1};
      bins last_wdata_handshake_to_bvalid_delay_mid = {[2:(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)]};
      bins last_wdata_handshake_to_bvalid_delay_max = {[(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)+1:$]};
      option.at_least = `SVT_AXI_trans_meta_axi_write_last_wdata_handshake_to_BVALID_Delay_COV_OPTION_AT_LEAST_VAL;
    }
    AWVALID_before_AWREADY :coverpoint cov_AWVALID_before_AWREADY {
      bins awvalid_before_awready = {1};
      option.at_least = `SVT_AXI_trans_meta_axi_write_AWVALID_before_AWREADY_COV_OPTION_AT_LEAST_VAL;
    }
    AWREADY_before_AWVALID :coverpoint cov_AWREADY_before_AWVALID {
      bins awready_before_awvalid = {1};
      option.at_least = `SVT_AXI_trans_meta_axi_write_AWREADY_before_AWVALID_COV_OPTION_AT_LEAST_VAL;
    }        
    BVALID_before_BREADY   :coverpoint cov_BVALID_before_BREADY {
      bins bvalid_before_bready = {1};
      option.at_least = `SVT_AXI_trans_meta_axi_write_BVALID_before_BREADY_COV_OPTION_AT_LEAST_VAL;
    }
    BREADY_before_BVALID   :coverpoint cov_BREADY_before_BVALID {
      bins bready_before_bvalid = {1};
      option.at_least = `SVT_AXI_trans_meta_axi_write_BREADY_before_BVALID_COV_OPTION_AT_LEAST_VAL;
    }        
    WVALID_before_WREADY  : coverpoint cov_WVALID_before_WREADY {  
      bins wvalid_before_wready = {1};
      option.at_least = `SVT_AXI_trans_meta_axi_write_WVALID_before_WREADY_COV_OPTION_AT_LEAST_VAL;
    }
    WREADY_before_WVALID  : coverpoint cov_WREADY_before_WVALID {   
      bins wready_before_wvalid = {1};
      option.at_least = `SVT_AXI_trans_meta_axi_write_WREADY_before_WVALID_COV_OPTION_AT_LEAST_VAL;
    }        
    AWVALID_before_WREADY : coverpoint cov_AWVALID_before_WREADY{
      bins awvalid_before_wready = {1};
      option.at_least = `SVT_AXI_trans_meta_axi_write_AWVALID_before_WREADY_COV_OPTION_AT_LEAST_VAL;
    }
    WREADY_before_AWVALID : coverpoint cov_WREADY_before_AWVALID{
      bins wready_before_awvalid = {1};
      option.at_least = `SVT_AXI_trans_meta_axi_write_WREADY_before_AWVALID_COV_OPTION_AT_LEAST_VAL;
    }        
    AWREADY_before_WVALID : coverpoint cov_AWREADY_before_WVALID{
      bins awready_before_wvalid = {1};
      option.at_least = `SVT_AXI_trans_meta_axi_write_AWREADY_before_WVALID_COV_OPTION_AT_LEAST_VAL;
    }        
    WVALID_before_AWREADY : coverpoint cov_WVALID_before_AWREADY{
      bins wvalid_before_awready = {1};
      option.at_least = `SVT_AXI_trans_meta_axi_write_WVALID_before_AWREADY_COV_OPTION_AT_LEAST_VAL;
    }
    AWVALID_before_WVALID : coverpoint cov_AWVALID_before_WVALID{
      bins awvalid_before_wvalid = {1};
      option.at_least = `SVT_AXI_trans_meta_axi_write_AWVALID_before_WVALID_COV_OPTION_AT_LEAST_VAL;
    }        
    WVALID_before_AWVALID : coverpoint cov_WVALID_before_AWVALID{
      bins wvalid_before_awvalid = {1};
      option.at_least = `SVT_AXI_trans_meta_axi_write_WVALID_before_AWVALID_COV_OPTION_AT_LEAST_VAL;
    }
  endgroup

  
  /**
    *  Covergroup: trans_meta_axi_read
    *
    *  Coverpoints:
    *  - ARVALID_to_ARREADY_Delay: Captures min, mid and max range of delays between signals arvalid and arready
    *  - RVALID_to_RREADY_Delay: Captures min, mid and max range of delays between signals rvalid and rready
    *  - ARVALID_to_prev_ARVALID_Delay: Captures min, mid and max range of delays between current and previous arvalid signals
    *  - RVALID_to_prev_RVALID_Delay: Captures min, mid and max range of delays between current and previous rvalid signals
    *  - ARVALID_to_first_RVALID_Delay: Captures min, mid and max range of delays between arvalid and first rvalid signals
    *  - ARVALID_before_ARREADY: Captures if ARVALID signal comes before ARREADY signal 
    *  - ARREADY_before_ARVALID: Captures if ARREADY signal comes before ARVALID signal
    *  - RVALID_before_RREADY: Captures if RVALID signal comes before RREADY signal 
    *  - RREADY_before_RVALID: Captures if RREADY signal comes before RVALID signal
    *  .
    */
  //covergroup trans_meta_axi_read @(cov_read_sample_event);
  covergroup trans_meta_axi_read ;
    option.per_instance = 1;
    ARVALID_to_ARREADY_Delay : coverpoint cov_ARVALID_to_ARREADY_Delay {
      bins arvalid_to_arready_delay_min = {0};
      bins arvalid_to_arready_delay_mid = {[1:(`SVT_AXI_MAX_ADDR_DELAY/2)]};
      bins arvalid_to_arready_delay_max = {[(`SVT_AXI_MAX_ADDR_DELAY/2)+1:$]};
    }
    RVALID_to_RREADY_Delay : coverpoint cov_RVALID_to_RREADY_Delay {
      bins rvalid_to_rready_delay_min = {0};
      bins rvalid_to_rready_delay_mid = {[1:(`SVT_AXI_MAX_RREADY_DELAY/2)]};
      bins rvalid_to_rready_delay_max = {[(`SVT_AXI_MAX_RREADY_DELAY/2)+1:$]};
    }
    ARVALID_to_prev_ARVALID_Delay : coverpoint cov_ARVALID_to_prev_ARVALID_Delay {
      bins arvalid_to_prev_arvalid_delay_min = {1};
      bins arvalid_to_prev_arvalid_delay_mid = {[2:((`SVT_AXI_MAX_ADDR_VALID_DELAY + `SVT_AXI_MAX_ADDR_DELAY)/2)]};
      bins arvalid_to_prev_arvalid_delay_max = {[((`SVT_AXI_MAX_ADDR_VALID_DELAY + `SVT_AXI_MAX_ADDR_DELAY)/2)+1:$]};
    } 
    RVALID_to_prev_RVALID_Delay : coverpoint cov_RVALID_to_prev_RVALID_Delay {
      bins rvalid_to_prev_rvalid_delay_min = {1};
      bins rvalid_to_prev_rvalid_delay_mid = {[2:((`SVT_AXI_MAX_RVALID_DELAY + `SVT_AXI_MAX_RREADY_DELAY)/2)]};
      bins rvalid_to_prev_rvalid_delay_max = {[((`SVT_AXI_MAX_RVALID_DELAY + `SVT_AXI_MAX_RREADY_DELAY)/2)+1:$]};
    } 
    ARVALID_to_first_RVALID_Delay : coverpoint cov_ARVALID_to_first_RVALID_Delay {
      bins arvalid_to_first_rvalid_delay_min = {[0:1]}; 
      bins arvalid_to_first_rvalid_delay_mid = {[2:(( `SVT_AXI_MAX_ADDR_DELAY + `SVT_AXI_MAX_RVALID_DELAY)/2)]};
      bins arvalid_to_first_rvalid_delay_max = {[((`SVT_AXI_MAX_ADDR_DELAY + `SVT_AXI_MAX_RVALID_DELAY)/2)+1:$]};
    }
    ARVALID_before_ARREADY: coverpoint cov_ARVALID_before_ARREADY {
      bins arvalid_before_arready = {1};
    }
    ARREADY_before_ARVALID: coverpoint cov_ARREADY_before_ARVALID {
      bins arready_before_arvalid = {1};
    }
    RVALID_before_RREADY: coverpoint cov_RVALID_before_RREADY {
      bins rvalid_before_rready = {1};
    }
    RREADY_before_RVALID: coverpoint cov_RREADY_before_RVALID {
      bins rready_before_rvalid = {1};
    }
  endgroup

    /**
    *  Covergroup: trans_axi4_stream_delay
    *
    *  Coverpoints:
    *  - TVALID_Delay: Captures min, mid and max range of delay signal tvalid
    *  - TREADY_Delay: Captures min, mid and max range of delay signal tready
    *  .
    */  
  covergroup trans_axi4_stream_delay ;
    option.per_instance = 1;
    TVALID_Delay : coverpoint cov_TVALID_Delay {
      bins tvalid_delay_min = {0};
      bins tvalid_delay_mid = {[1:(`SVT_AXI_MAX_TVALID_DELAY/2)]};
      bins tvalid_delay_max = {[(`SVT_AXI_MAX_TVALID_DELAY/2)+1:$]};
    } 
    TREADY_Delay : coverpoint cov_TREADY_Delay {
      bins tready_delay_min = {0};
      bins tready_delay_mid = {[1:(`SVT_AXI_MAX_TREADY_DELAY/2)]};
      bins tready_delay_max = {[(`SVT_AXI_MAX_TREADY_DELAY/2)+1:$]};
    }      
  endgroup

    /**
    *  Covergroup: trans_meta_axi4_stream
    *
    *  Coverpoints:
    *  - TVALID_to_TREADY_Delay: Captures min, mid and max range of delays between signals tvalid and tready
    *  - TVALID_to_prev_TVALID_Delay: Captures min, mid and max range of delays between current and previous tvalid signals
    *  - TVALID_before_TREADY: Captures if TVALID signal comes before TREADY signal 
    *  - TREADY_before_TVALID: Captures if TREADY signal comes before TVALID signal 
    *  .
    */  
  covergroup trans_meta_axi4_stream ;
    option.per_instance = 1;
    TVALID_to_TREADY_Delay : coverpoint cov_TVALID_to_TREADY_Delay {
      bins tvalid_to_tready_delay_min = {0};
      bins tvalid_to_tready_delay_mid = {[1:(`SVT_AXI_MAX_TREADY_DELAY/2)]};
      bins tvalid_to_tready_delay_max = {[(`SVT_AXI_MAX_TREADY_DELAY/2)+1:$]};
      option.at_least = `SVT_AXI4_STREAM_trans_TVALID_to_TREADY_Delay_COV_OPTION_AT_LEAST_VAL;
    } 
    TVALID_to_prev_TVALID_Delay : coverpoint cov_TVALID_to_prev_TVALID_Delay {
      bins tvalid_to_prev_tvalid_delay_min = {1};
      bins tvalid_to_prev_tvalid_delay_mid = {[2:((`SVT_AXI_MAX_TVALID_DELAY + `SVT_AXI_MAX_TREADY_DELAY)/2)]};
      bins tvalid_to_prev_tvalid_delay_max = {[((`SVT_AXI_MAX_TVALID_DELAY +  `SVT_AXI_MAX_TREADY_DELAY)/2)+1:$]};
      option.at_least = `SVT_AXI4_STREAM_trans_TVALID_to_prev_TVALID_Delay_COV_OPTION_AT_LEAST_VAL;
    }        
    TVALID_before_TREADY  : coverpoint cov_TVALID_before_TREADY {  
      bins tvalid_before_tready = {1};
      option.at_least = `SVT_AXI4_STREAM_trans_TVALID_before_TREADY_COV_OPTION_AT_LEAST_VAL;
    }
    TREADY_before_TVALID  : coverpoint cov_TREADY_before_TVALID {   
      bins tready_before_tvalid = {1};
      option.at_least = `SVT_AXI4_STREAM_trans_TREADY_before_TVALID_COV_OPTION_AT_LEAST_VAL;
    }        
  endgroup

  /**
    *  Covergroup: trans_axi_write_handshake_delay
    *
    *  Coverpoints:
    *  - last_AWVALID_AWREADY_handshake_to_next_AWVALID_AWREADY_handshake_Delay:Captures min, mid and max range of delays between last awvalid_awready handshake to the next awvalid_awready handshake 
    *  - last_AWVALID_AWREADY_handshake_to_next_AWVALID_Delay: Captures min,mid and max range of delays between last awvalid_awready handshake to the next awvalid
    *  - last_AWVALID_AWREADY_handshake_to_next_AWREADY_Delay: Captures min,mid and max range of delays between last awvalid_awready handshake to the next awready
    *  - last_AWREADY_to_next_AWVALID_AWREADY_handshake_Delay: Captures min,mid and max range of delays between last awready to the next awvalid_awready handshake  
    *  - last_WVALID_WREADY_handshake_to_next_WVALID_WREADY_handshake_Delay: Captures min, mid and max range of delays between last wvalid_wready handshake to the next wvalid_wready handshake 
    *  - last_WVALID_WREADY_data_beat_handshake_to_next_WVALID_WREADY_first_data_beat_handshake_Delay: Captures min, mid and max range of delays between last wvalid_wready data beat handshake to the next wvalid_wready data beat handshake 
    *  - last_WVALID_WREADY_handshake_to_next_WVALID_Delay: Captures min, mid and max range of delays between last wvalid_wready handshake to the next wvalid 
    *  - last_WVALID_WREADY_handshake_to_next_WREADY_Delay: Captures min, mid and max range of delays between last wvalid_wready handshake to the next wready
    *  - last_WREADY_to_next_WVALID_WREADY_handshake_Delay: Captures min,mid and max range of delays between last wready to the next wvalid_wready handshake  
    *  - last_BVALID_BREADY_handshake_to_next_BVALID_BREADY_handshake_Delay:Captures min, mid and max range of delays between last bvalid_bready handshake to the next bvalid_bready handshake 
    *  - last_BVALID_BREADY_handshake_to_next_BVALID_Delay: Captures min, mid and max range of delays between last bvalid_bready handshake to the next bvalid 
    *  - last_BVALID_BREADY_handshake_to_next_BREADY_Delay: Captures min, mid and max range of delays between last bvalid_bready handshake to the next bready
    *  - last_BVALID_to_next_BVALID_Delay: Captures min, mid and max range of delays between last bvalid to the next bvalid
    *  - last_BREADY_to_next_BREADY_Delay: Captures min, mid and max range of delays between last bready to the next bready 
    *  - last_BREADY_to_next_BVALID_BREADY_handshake_Delay: Captures min, mid and max range of delays between last bready to the next bvalid_bready handshake   
    *  .
    */
  covergroup trans_axi_write_handshake_delay;
    option.per_instance = 1;
    last_AWVALID_AWREADY_handshake_to_next_AWVALID_AWREADY_handshake_Delay : coverpoint cov_last_AWVALID_AWREADY_handshake_to_next_AWVALID_AWREADY_handshake_Delay {
      bins last_awvalid_awready_handshake_to_next_awvalid_awready_handshake_delay_min = {1};
      bins last_awvalid_awready_handshake_to_next_awvalid_awready_handshake_delay_mid = {[2:(`SVT_AXI_MAX_ADDR_DELAY/2)]};
      bins last_awvalid_awready_handshake_to_next_awvalid_awready_handshake_delay_max = {[(`SVT_AXI_MAX_ADDR_DELAY/2)+1:$]};
    } 
    last_AWVALID_AWREADY_handshake_to_next_AWVALID_Delay : coverpoint cov_prev_handshake_AWVALID_Delay {
      bins last_awvalid_awready_handshake_to_next_awvalid_delay_min = {1};
      bins last_awvalid_awready_handshake_to_next_awvalid_delay_mid = {[2:(`SVT_AXI_MAX_ADDR_DELAY/2)]};
      bins last_awvalid_awready_handshake_to_next_awvalid_delay_max = {[(`SVT_AXI_MAX_ADDR_DELAY/2)+1:$]};
    }   
    last_AWVALID_AWREADY_handshake_to_next_AWREADY_Delay : coverpoint cov_prev_handshake_AWREADY_Delay {
      bins last_awvalid_awready_handshake_to_next_awready_delay_min = {1};
      bins last_awvalid_awready_handshake_to_next_awready_delay_mid = {[2:(`SVT_AXI_MAX_ADDR_DELAY/2)]};
      bins last_awvalid_awready_handshake_to_next_awready_delay_max = {[(`SVT_AXI_MAX_ADDR_DELAY/2)+1:$]};
    }
    last_AWREADY_to_next_AWVALID_AWREADY_handshake_Delay : coverpoint cov_prev_AWREADY_to_handshake_Delay {
      bins last_awready_to_next_awvalid_awready_handshake_delay_min = {1};
      bins last_awready_to_next_awvalid_awready_handshake_delay_mid = {[2:(`SVT_AXI_MAX_ADDR_DELAY/2)]};
      bins last_awready_to_next_awvalid_awready_handshake_delay_max = {[(`SVT_AXI_MAX_ADDR_DELAY/2)+1:$]};
    }
    last_WVALID_WREADY_handshake_to_next_WVALID_WREADY_handshake_Delay : coverpoint cov_last_WVALID_WREADY_handshake_to_next_WVALID_WREADY_handshake_Delay {
      bins last_wvalid_wready_handshake_to_next_wvalid_wready_handshake_delay_min = {1};
      bins last_wvalid_wready_handshake_to_next_wvalid_wready_handshake_delay_mid = {[2:((`SVT_AXI_MAX_WVALID_DELAY + `SVT_AXI_MAX_WREADY_DELAY)/2)]};
      bins last_wvalid_wready_handshake_to_next_wvalid_wready_handshake_delay_max = {[((`SVT_AXI_MAX_WVALID_DELAY +  `SVT_AXI_MAX_WREADY_DELAY)/2)+1:$]};
    }
    last_WVALID_WREADY_data_beat_handshake_to_next_WVALID_WREADY_first_data_beat_handshake_Delay : coverpoint cov_last_WVALID_WREADY_data_beat_handshake_to_next_WVALID_WREADY_first_data_beat_handshake_Delay {
      bins last_WVALID_WREADY_data_beat_handshake_to_next_WVALID_WREADY_first_data_beat_handshake_delay_min = {1};
      bins last_WVALID_WREADY_data_beat_handshake_to_next_WVALID_WREADY_first_data_beat_handshake_delay_mid = {[2:((`SVT_AXI_MAX_WVALID_DELAY + `SVT_AXI_MAX_WREADY_DELAY)/2)]};
      bins last_WVALID_WREADY_data_beat_handshake_to_next_WVALID_WREADY_first_data_beat_handshake_delay_max = {[((`SVT_AXI_MAX_WVALID_DELAY +  `SVT_AXI_MAX_WREADY_DELAY)/2)+1:$]};
    }
    last_WVALID_WREADY_handshake_to_next_WVALID_Delay : coverpoint cov_last_WVALID_WREADY_handshake_to_next_WVALID_Delay {
      bins last_wvalid_wready_handshake_to_next_wvalid_delay_min = {1};
      bins last_wvalid_wready_handshake_to_next_wvalid_delay_mid = {[2:(`SVT_AXI_MAX_WVALID_DELAY/2)]};
      bins last_wvalid_wready_handshake_to_next_wvalid_delay_max = {[(`SVT_AXI_MAX_WVALID_DELAY/2)+1:$]};
    }
    last_WVALID_WREADY_handshake_to_next_WREADY_Delay : coverpoint cov_last_WVALID_WREADY_handshake_to_next_WREADY_Delay {
      bins last_wvalid_wready_handshake_to_next_wready_delay_min = {1};
      bins last_wvalid_wready_handshake_to_next_wready_delay_mid = {[2:(`SVT_AXI_MAX_WREADY_DELAY/2)]};
      bins last_wvalid_wready_handshake_to_next_wready_delay_max = {[(`SVT_AXI_MAX_WREADY_DELAY/2)+1:$]};
    }
    last_WREADY_to_next_WVALID_WREADY_handshake_Delay : coverpoint cov_last_WREADY_to_next_WVALID_WREADY_handshake_Delay {
      bins last_wready_to_next_wvalid_wready_handshake_delay_min = {1};
      bins last_wready_to_next_wvalid_wready_handshake_delay_mid = {[2:((`SVT_AXI_MAX_WVALID_DELAY + `SVT_AXI_MAX_WREADY_DELAY)/2)]};
      bins last_wready_to_next_wvalid_wready_handshake_delay_max = {[((`SVT_AXI_MAX_WVALID_DELAY +  `SVT_AXI_MAX_WREADY_DELAY)/2)+1:$]};
    }
    last_BVALID_BREADY_handshake_to_next_BVALID_BREADY_handshake_Delay : coverpoint cov_last_BVALID_BREADY_handshake_to_next_BVALID_BREADY_handshake_Delay {
      bins last_bvalid_bready_handshake_to_next_bvalid_bready_handshake_delay_min = {1};
      bins last_bvalid_bready_handshake_to_next_bvalid_bready_handshake_delay_mid = {[2:(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)]};
      bins last_bvalid_bready_handshake_to_next_bvalid_bready_handshake_delay_max = {[(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)+1:$]};
    }
    last_BVALID_BREADY_handshake_to_next_BVALID_Delay : coverpoint cov_last_BVALID_BREADY_handshake_to_next_BVALID_Delay {
      bins last_bvalid_bready_handshake_to_next_bvalid_delay_min = {1};
      bins last_bvalid_bready_handshake_to_next_bvalid_delay_mid = {[2:(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)]};
      bins last_bvalid_bready_handshake_to_next_bvalid_delay_max = {[(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)+1:$]};
    }
    last_BVALID_BREADY_handshake_to_next_BREADY_Delay : coverpoint cov_last_BVALID_BREADY_handshake_to_next_BREADY_Delay {
      bins last_bvalid_bready_handshake_to_next_bready_delay_min = {1};
      bins last_bvalid_bready_handshake_to_next_bready_delay_mid = {[2:(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)]};
      bins last_bvalid_bready_handshake_to_next_bready_delay_max = {[(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)+1:$]};
    }
    last_BVALID_to_next_BVALID_Delay : coverpoint cov_BVALID_to_next_BVALID_Delay {
      bins last_BVALID_to_next_BVALID_delay_min = {1};
      bins last_BVALID_to_next_BVALID_delay_mid = {[2:(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)]};
      bins last_BVALID_to_next_BVALID_delay_max = {[(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)+1:$]};
    }
    last_BREADY_to_next_BREADY_Delay : coverpoint cov_last_BREADY_to_next_BREADY_Delay {
      bins last_BREADY_to_next_BREADY_delay_min = {1};
      bins last_BREADY_to_next_BREADY_delay_mid = {[2:(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)]};
      bins last_BREADY_to_next_BREADY_delay_max = {[(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)+1:$]};
    }
    last_BREADY_to_next_BVALID_BREADY_handshake_Delay : coverpoint cov_last_BREADY_to_next_BVALID_BREADY_handshake_Delay {
      bins last_bready_to_next_bvalid_bready_handshake_delay_min = {1};
      bins last_bready_to_next_bvalid_bready_handshake_delay_mid = {[2:(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)]};
      bins last_bready_to_next_bvalid_bready_handshake_delay_max = {[(`SVT_AXI_MAX_WRITE_RESP_DELAY/2)+1:$]};
    }
  endgroup

  /** 
    *  Covergroup: trans_axi_read_handshake_delay
    *
    *  Coverpoints:
    *  - last_ARVALID_ARREADY_handshake_to_next_ARVALID_ARREADY_handshake_Delay:Captures min, mid and max range of delays between last arvalid_arready handshake to the next arvalid_arready handshake 
    *  - last_ARVALID_ARREADY_handshake_to_next_ARVALID_Delay: Captures min,mid and max range of delays between last arvalid_arready handshake to the next arvalid
    *  - last_ARVALID_ARREADY_handshake_to_next_ARREADY_Delay: Captures min,mid and max range of delays between last arvalid_arready handshake to the next arready
    *  - last_ARREADY_to_next_ARVALID_ARREADY_handshake_Delay: Captures min,mid and max range of delays between last arready to the next arvalid_arready handshake  
    *  - last_RVALID_RREADY_handshake_to_next_RVALID_RREADY_handshake_Delay:Captures min, mid and max range of delays between last rvalid_rready handshake to the next rvalid_rready handshake 
    *  - last_RVALID_RREADY_handshake_to_next_RVALID_Delay: Captures min,mid and max range of delays between last rvalid_rready handshake to the next rvalid
    *  - last_RVALID_RREADY_handshake_to_next_RREADY_Delay: Captures min,mid and max range of delays between last rvalid_rready handshake to the next rready
    *  - last_RREADY_to_next_RVALID_RREADY_handshake_Delay: Captures min,mid and max range of delays between last rready to the next rvalid_rready handshake 
    *  - last_RVALID_RREADY_data_beat_handshake_to_next_RVALID_RREADY_first_data_beat_handshake_Delay: Captures min, mid and max range of delays between last rvalid_rready data beat handshake to the next rvalid_rready data beat handshake 
    *  .
    */
  covergroup trans_axi_read_handshake_delay;
    option.per_instance = 1;
    last_ARVALID_ARREADY_handshake_to_next_ARVALID_ARREADY_handshake_Delay : coverpoint cov_last_ARVALID_ARREADY_handshake_to_next_ARVALID_ARREADY_handshake_Delay {
      bins last_arvalid_arready_handshake_to_next_arvalid_arready_handshake_delay_min = {1};
      bins last_arvalid_arready_handshake_to_next_arvalid_arready_handshake_delay_mid = {[2:(`SVT_AXI_MAX_ADDR_DELAY/2)]};
      bins last_arvalid_arready_handshake_to_next_arvalid_arready_handshake_delay_max = {[(`SVT_AXI_MAX_ADDR_DELAY/2)+1:$]};
    }
    last_ARVALID_ARREADY_handshake_to_next_ARVALID_Delay : coverpoint cov_prev_handshake_ARVALID_Delay {
      bins last_arvalid_arready_handshake_to_next_arvalid_delay_min = {1};
      bins last_arvalid_arready_handshake_to_next_arvalid_delay_mid = {[2:(`SVT_AXI_MAX_ADDR_DELAY/2)]};
      bins last_arvalid_arready_handshake_to_next_arvalid_delay_max = {[(`SVT_AXI_MAX_ADDR_DELAY/2)+1:$]};
    }
    last_ARVALID_ARREADY_handshake_to_next_ARREADY_Delay : coverpoint cov_prev_handshake_ARREADY_Delay {
      bins last_arvalid_arready_handshake_to_next_arready_delay_min = {1};
      bins last_arvalid_arready_handshake_to_next_arready_delay_mid = {[2:(`SVT_AXI_MAX_ADDR_DELAY/2)]};
      bins last_arvalid_arready_handshake_to_next_arready_delay_max = {[(`SVT_AXI_MAX_ADDR_DELAY/2)+1:$]};
    }
    last_ARREADY_to_next_ARVALID_ARREADY_handshake_Delay : coverpoint cov_prev_ARREADY_to_handshake_Delay {
      bins last_arready_to_next_arvalid_arready_handshake_delay_min = {1};
      bins last_arready_to_next_arvalid_arready_handshake_delay_mid = {[2:(`SVT_AXI_MAX_ADDR_DELAY/2)]};
      bins last_arready_to_next_arvalid_arready_handshake_delay_max = {[(`SVT_AXI_MAX_ADDR_DELAY/2)+1:$]};
    }
    last_RVALID_RREADY_handshake_to_next_RVALID_RREADY_handshake_Delay : coverpoint cov_last_RVALID_RREADY_handshake_to_next_RVALID_RREADY_handshake_Delay {
      bins last_rvalid_rready_handshake_to_next_rvalid_rready_handshake_delay_min = {1};
      bins last_rvalid_rready_handshake_to_next_rvalid_rready_handshake_delay_mid = {[2:((`SVT_AXI_MAX_RVALID_DELAY + `SVT_AXI_MAX_RREADY_DELAY)/2)]};
      bins last_rvalid_rready_handshake_to_next_rvalid_rready_handshake_delay_max = {[((`SVT_AXI_MAX_RVALID_DELAY + `SVT_AXI_MAX_RREADY_DELAY)/2)+1:$]};
    }
    last_RVALID_RREADY_handshake_to_next_RVALID_Delay : coverpoint cov_last_RVALID_RREADY_handshake_to_next_RVALID_Delay {
      bins last_rvalid_rready_handshake_to_next_rvalid_delay_min = {1};
      bins last_rvalid_rready_handshake_to_next_rvalid_delay_mid = {[2:(`SVT_AXI_MAX_RVALID_DELAY/2)]};
      bins last_rvalid_rready_handshake_to_next_rvalid_delay_max = {[(`SVT_AXI_MAX_RVALID_DELAY/2)+1:$]};
    }
    last_RVALID_RREADY_handshake_to_next_RREADY_Delay : coverpoint cov_last_RVALID_RREADY_handshake_to_next_RREADY_Delay {
      bins last_rvalid_rready_handshake_to_next_rready_delay_min = {1};
      bins last_rvalid_rready_handshake_to_next_rready_delay_mid = {[2:(`SVT_AXI_MAX_RREADY_DELAY/2)]};
      bins last_rvalid_rready_handshake_to_next_rready_delay_max = {[(`SVT_AXI_MAX_RREADY_DELAY/2)+1:$]};
    }
    last_RREADY_to_next_RVALID_RREADY_handshake_Delay : coverpoint cov_last_RREADY_to_next_RVALID_RREADY_handshake_Delay {
      bins last_rready_to_next_rvalid_rready_handshake_delay_min = {1};
      bins last_rready_to_next_rvalid_rready_handshake_delay_mid = {[2:((`SVT_AXI_MAX_RVALID_DELAY + `SVT_AXI_MAX_RREADY_DELAY)/2)]};
      bins last_rready_to_next_rvalid_rready_handshake_delay_max = {[((`SVT_AXI_MAX_RVALID_DELAY +  `SVT_AXI_MAX_RREADY_DELAY)/2)+1:$]};
    }
    last_RVALID_RREADY_data_beat_handshake_to_next_RVALID_RREADY_first_data_beat_handshake_Delay : coverpoint cov_last_RVALID_RREADY_data_beat_handshake_to_next_RVALID_RREADY_first_data_beat_handshake_Delay {
      bins last_RVALID_RREADY_data_beat_handshake_to_next_RVALID_RREADY_first_data_beat_handshake_delay_min = {1};
      bins last_RVALID_RREADY_data_beat_handshake_to_next_RVALID_RREADY_first_data_beat_handshake_delay_mid = {[2:((`SVT_AXI_MAX_WVALID_DELAY + `SVT_AXI_MAX_WREADY_DELAY)/2)]};
      bins last_RVALID_RREADY_data_beat_handshake_to_next_RVALID_RREADY_first_data_beat_handshake_delay_max = {[((`SVT_AXI_MAX_WVALID_DELAY +  `SVT_AXI_MAX_WREADY_DELAY)/2)+1:$]};
    }
  endgroup

 
  // ****************************************************************************
  // ACE Covergroups
  // ****************************************************************************

 /**
  *
  * Covergroup     : trans_cross_ace_acsnoop_acaddr
  * 
  * Coverpoints:
  *
  * - snoop_xact_type:  Captures Snoop transaction
  * - snoop_addr:      Captures Snoop address
  * .
  *
  * Cross coverpoints:
  * - acsnoop_acaddr : Crosses cover points snoop_xact_type and snoop_addr
  * .
  *
  */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_acsnoop_acaddr @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_ADDR

    acsnoop_acaddr : cross snoop_xact_type, snoop_addr {

      ignore_bins Ignore_invalid_addr = binsof(snoop_xact_type) intersect {
                                        svt_axi_snoop_transaction::DVMMESSAGE,svt_axi_snoop_transaction::DVMCOMPLETE} iff(cfg.dvm_enable == 1'b0);

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  /** 
   * This covergroup will be created when there is only one ACE-master and
   * minimum one or more than one ACE_LITE master in the system. 
   */
  covergroup trans_cross_ace_acsnoop_acaddr_one_ace_acelite @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_ONE_ACE_ACELITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_ADDR

    acsnoop_acaddr : cross snoop_xact_type, snoop_addr {

      ignore_bins Ignore_invalid_addr = binsof(snoop_xact_type) intersect {
                                        svt_axi_snoop_transaction::DVMMESSAGE,svt_axi_snoop_transaction::DVMCOMPLETE} iff(cfg.dvm_enable == 1'b0);

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else
  covergroup trans_cross_ace_acsnoop_acaddr_dvm_unset @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_ADDR

    acsnoop_acaddr : cross snoop_xact_type, snoop_addr {


      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /** 
   * This covergroup will be created when there is only one ACE-master and
   * minimum one or more than one ACE_LITE master in the system. 
   */
  covergroup trans_cross_ace_acsnoop_acaddr_dvm_unset_one_ace_acelite @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_UNSET_ONE_ACE_ACELITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_ADDR

    acsnoop_acaddr : cross snoop_xact_type, snoop_addr {


      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_ace_acsnoop_acaddr_dvm_set @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_ADDR

    acsnoop_acaddr : cross snoop_xact_type, snoop_addr {

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  /** 
   * This covergroup will be created when there is only one ACE-master and
   * minimum one or more than one ACE_LITE master in the system. 
   */
  covergroup trans_cross_ace_acsnoop_acaddr_dvm_set_one_ace_acelite @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_SET_ONE_ACE_ACELITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_ADDR

    acsnoop_acaddr : cross snoop_xact_type, snoop_addr {

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`endif

  /**
    * Covergroup: trans_ace_concurrent_overlapping_arsnoop_acsnoop
    * This covergroups 
    * Coverpoints:
    * snoop_xact_type:Coverpoint of svt_axi_snoop_transaction::snoop_xact_type for all snoop transactions recieved on master port . This excludes DVMMESSAGE,DVMCOMPLETE transactions
    * coherent_read_xact_type:Coverpoint of svt_axi_transaction::coherent_xact_type for all coherent transactions initiated on read channel of master . This excludes READNOSNOOP,DVMMESSAGE,DVMCOMPLETE,READBARRIER 
    * transactions
    * The bins in this covergroup will be hit when a coherent transaction  is outstanding while a snoop transaction is outstanding on same port with overlapping address
    * Two  ACE  masters needed for this covergroup
    * 
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.6.2
    *
    */
  covergroup trans_ace_concurrent_overlapping_arsnoop_acsnoop;
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_NO_DVM_NO_BARRIER_NO_READNOSNOOP
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_NO_DVM
       ace_concurrent_overlap_snoop_xact : cross snoop_xact_type,coherent_read_xact_type{
       option.weight=1;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_ace_concurrent_overlapping_arsnoop_acsnoop_one_ace_acelite
    * This covergroup will be created when there is only one ACE-master and
    * minimum one or more than one ACE_LITE master in the system.
    * Coverpoints:
    * snoop_xact_type:Coverpoint of svt_axi_snoop_transaction::snoop_xact_type for READONCE,CLEANSHARED,CLEANINVALID and MAKEINVALID snoop transactions recieved on master port . This excludes READSHARED,READCLEAN,READNOTSHAREDDIRTY,READUNIQUE,DVMMESSAGE,DVMCOMPLETE transactions
    * coherent_read_xact_type:Coverpoint of svt_axi_transaction::coherent_xact_type for all coherent transactions initiated on read channel of master . This excludes READNOSNOOP,DVMMESSAGE,DVMCOMPLETE,READBARRIER transactions
    * The bins in this covergroup will be hit when a coherent transaction is outstanding while a snoop transaction is outstanding on same port with overlapping address
    * Atleast one ACE and one ACE_LITE master needed for this covergroup
    * 
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.6.2
    *
    */
  covergroup trans_ace_concurrent_overlapping_arsnoop_acsnoop_one_ace_acelite;
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_NO_DVM_NO_BARRIER_NO_READNOSNOOP
       
       snoop_xact_type : coverpoint master_snoop_xact_type { 
       bins snoop_readonce_xact   = {svt_axi_snoop_transaction::READONCE}; 
       bins snoop_cleanshared_xact   = {svt_axi_snoop_transaction::CLEANSHARED}; 
       bins snoop_cleaninvalid_xact   = {svt_axi_snoop_transaction::CLEANINVALID}; 
       bins snoop_makeinvalid_xact   = {svt_axi_snoop_transaction::MAKEINVALID}; 
       option.weight = 1; 
    } 
       ace_concurrent_overlap_snoop_xact : cross snoop_xact_type,coherent_read_xact_type{
       option.weight=1;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_enabled
    * The bins in covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_enabled will be hit when a coherent transaction  is outstanding while a snoop transaction is outstanding on same port with overlapping address
    * The covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_enabled is applicable only for ACE Masters .The covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_enabled needs at least two ACE masters in the system .
    * Coverpoints:
    * snoop_xact_type:Coverpoint of svt_axi_snoop_transaction::snoop_xact_type for all snoop transactions recieved on master port . This excludes DVMMESSAGE,DVMCOMPLETE transactions
    * coherent_write_xact_type_generate_snoop:Coverpoint of svt_axi_transaction::coherent_xact_type for all coherent transactions initiated on write channel of master .This coverpoint includes only those transactions that     * generate snoop.This includes WRITEUNIQUE and WRITELINEUNIQUE transactions  
    * snoop_crresp_on_ace_port :
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.6.2
    *
    */
  covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_enabled;
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_WRITEEVICT_SNOOP_GENERATE
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_NO_DVM
       
       snoop_crresp_on_ace_port: coverpoint snoop_resp_ace_master[3:0] {
       bins cresp_0000 = {4'b0000};
       bins cresp_1000 = {4'b1000};
       bins cresp_0001 = {4'b0001};
       bins cresp_1001 = {4'b1001};
       bins cresp_0101 = {4'b0101};
       bins cresp_1101 = {4'b1101};    
       option.weight = 1;
    }
       snoop_crresp_wu : coverpoint snoop_resp_ace_master[4] {
         bins cresp_wasunique = {1'b1};
         bins cresp_wasnotunique = {1'b0};
         option.weight = 1;
    }    

       ace_concurrent_overlap_snoop_xact : cross snoop_xact_type,coherent_write_xact_type_gen_snoop,snoop_crresp_on_ace_port,snoop_crresp_wu{
       // Ignoring snoop_responses where is_shared is asserted and where data_transfer is asserted as recommended behaviour for MAKEINVALID is not tot transfer data 
       ignore_bins Ignore_invalid_rresp_ud_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::MAKEINVALID} &&
                                                 !binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b0000 };
      // Ignoring snoop_responses where is_shared bit is asserted or where data_transfer is asserted and pass_dirty is deasserted as CLEANINVALID will transfer data only when pass_dirty is asserted 
       ignore_bins ignore_invalid_rresp_ud_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::CLEANINVALID} &&
                                                 !binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b0000,4'b0101,4'b0001};
      // ignoring snoop_responses where is_shared bit is asserted for READUNIQUE transactions 
      ignore_bins Ignore_invalid_rresp_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::READUNIQUE} &&
                                                 binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b1101,4'b1000,4'b1001};
     // Ignoring the below ignore_bins for writeback and writeclean  transactions as mastercan invalidate the snoop responses 
     /* ignore_bins ignore_invalid_snoop_crresp_writeback = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITEBACK} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0001,4'b1000,4'b1001,4'b0000,4'b1101};
      ignore_bins ignore_invalid_snoop_crresp_writeclean = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITECLEAN} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0001,4'b1000,4'b1001,4'b0000};*/
      ignore_bins ignore_invalid_snoop_crresp_writeunique = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITEUNIQUE} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1101};
      ignore_bins ignore_invalid_snoop_crresp_writelineunique = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITELINEUNIQUE} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1101};
      ignore_bins ignore_invalid_snoop_crresp_evict = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::EVICT} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1001,4'b1101,4'b1000};

      option.weight=1;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite_writeevict_enabled
    * This covergroup will be created when there is only one ACE-master and
    * minimum one or more than one ACE_LITE master in the system.
    * The bins in covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite_writeevict_enabled will be hit when a coherent transaction is outstanding while a snoop transaction is outstanding on same port with overlapping address
    * The covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite_writeevict_enabled is applicable only for ACE Masters. The covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite_writeevict_enabled needs atleast one ACE and one ACE_LITE master in the system.
    * Coverpoints:
    * snoop_xact_type:Coverpoint of svt_axi_snoop_transaction::snoop_xact_type for READONCE,CLEANSHARED,CLEANINVALID and MAKEINVALID snoop transactions recieved on master port . This excludes READSHARED,READCLEAN,READNOTSHAREDDIRTY,READUNIQUE,DVMMESSAGE,DVMCOMPLETE transactions
    * coherent_write_xact_type_generate_snoop:Coverpoint of svt_axi_transaction::coherent_xact_type for all coherent transactions initiated on write channel of master. This coverpoint includes only those transactions that     
    * generate snoop.This includes WRITEUNIQUE and WRITELINEUNIQUE transactions  
    * snoop_crresp_on_ace_port : Coverpoint of cresp.
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.6.2
    *
    */
  covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite_writeevict_enabled;
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_WRITEEVICT_SNOOP_GENERATE
       
       snoop_xact_type : coverpoint master_snoop_xact_type { 
       bins snoop_readonce_xact   = {svt_axi_snoop_transaction::READONCE}; 
       bins snoop_cleanshared_xact   = {svt_axi_snoop_transaction::CLEANSHARED}; 
       bins snoop_cleaninvalid_xact   = {svt_axi_snoop_transaction::CLEANINVALID}; 
       bins snoop_makeinvalid_xact   = {svt_axi_snoop_transaction::MAKEINVALID}; 
       option.weight = 1; 
    }
       
       snoop_crresp_on_ace_port: coverpoint snoop_resp_ace_master[3:0] {
       bins cresp_0000 = {4'b0000};
       bins cresp_1000 = {4'b1000};
       bins cresp_0001 = {4'b0001};
       bins cresp_1001 = {4'b1001};
       bins cresp_0101 = {4'b0101};
       bins cresp_1101 = {4'b1101};    
       option.weight = 1;
    }
       snoop_crresp_wu : coverpoint snoop_resp_ace_master[4] {
         bins cresp_wasunique = {1'b1};
         bins cresp_wasnotunique = {1'b0};
         option.weight = 1;
    }    

       ace_concurrent_overlap_snoop_xact : cross snoop_xact_type,coherent_write_xact_type_gen_snoop,snoop_crresp_on_ace_port,snoop_crresp_wu{
       // Ignoring snoop_responses where is_shared is asserted and where data_transfer is asserted as recommended behaviour for MAKEINVALID is not tot transfer data 
       ignore_bins Ignore_invalid_rresp_ud_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::MAKEINVALID} &&
                                                 !binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b0000 };
      // Ignoring snoop_responses where is_shared bit is asserted or where data_transfer is asserted and pass_dirty is deasserted as CLEANINVALID will transfer data only when pass_dirty is asserted 
       ignore_bins ignore_invalid_rresp_ud_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::CLEANINVALID} &&
                                                 !binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b0000,4'b0101,4'b0001};

      ignore_bins ignore_invalid_snoop_crresp_writeunique = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITEUNIQUE} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1101};
      ignore_bins ignore_invalid_snoop_crresp_writelineunique = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITELINEUNIQUE} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1101};
      ignore_bins ignore_invalid_snoop_crresp_evict = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::EVICT} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1001,4'b1101,4'b1000};

      option.weight=1;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_disabled
    * The bins in covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_disabled will be hit when a coherent transaction  is outstanding while a snoop transaction is outstanding on same port with overlapping address
    * The covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_disabled is applicable only for ACE Masters .The covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_disabled needs at least two ACE masters in the system .
    * Coverpoints:
    * snoop_xact_type:Coverpoint of svt_axi_snoop_transaction::snoop_xact_type for all snoop transactions recieved on master port . This excludes DVMMESSAGE,DVMCOMPLETE transactions
    * coherent_write_xact_type_generate_snoop:Coverpoint of svt_axi_transaction::coherent_xact_type for all coherent transactions initiated on write channel of master .This coverpoint includes only those transactions that     * generate snoop.This includes WRITEUNIQUE and WRITELINEUNIQUE transactions  
    * snoop_crresp_on_ace_port :
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.6.2
    *
    */

  covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_disabled;
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NO_WRITEEVICT_SNOOP_GENERATE
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_NO_DVM
       
       snoop_crresp_on_ace_port: coverpoint snoop_resp_ace_master[3:0] {
       bins cresp_0000 = {4'b0000};
       bins cresp_1000 = {4'b1000};
       bins cresp_0001 = {4'b0001};
       bins cresp_1001 = {4'b1001};
       bins cresp_0101 = {4'b0101};
       bins cresp_1101 = {4'b1101};    
       option.weight = 1;
    }
       snoop_crresp_wu : coverpoint snoop_resp_ace_master[4] {
         bins cresp_wasunique = {1'b1};
         bins cresp_wasnotunique = {1'b0};
         option.weight = 1;
    }    

       ace_concurrent_overlap_snoop_xact : cross snoop_xact_type,coherent_write_xact_type_gen_snoop,snoop_crresp_on_ace_port,snoop_crresp_wu{
       // Ignoring snoop_responses where is_shared is asserted and where data_transfer is asserted as recommended behaviour for MAKEINVALID is not tot transfer data 
       ignore_bins Ignore_invalid_rresp_ud_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::MAKEINVALID} &&
                                                 !binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b0000 };
      // Ignoring snoop_responses where is_shared bit is asserted or where data_transfer is asserted and pass_dirty is deasserted as CLEANINVALID will transfer data only when pass_dirty is asserted 
       ignore_bins ignore_invalid_rresp_ud_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::CLEANINVALID} &&
                                                 !binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b0000,4'b0101,4'b0001};
      // ignoring snoop_responses where is_shared bit is asserted for READUNIQUE transactions 
      ignore_bins Ignore_invalid_rresp_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::READUNIQUE} &&
                                                 binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b1101,4'b1000,4'b1001};
     // Ignoring the below ignore_bins for writeback and writeclean  transactions as mastercan invalidate the snoop responses 
     /* ignore_bins ignore_invalid_snoop_crresp_writeback = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITEBACK} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0001,4'b1000,4'b1001,4'b0000,4'b1101};
      ignore_bins ignore_invalid_snoop_crresp_writeclean = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITECLEAN} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0001,4'b1000,4'b1001,4'b0000};*/
      ignore_bins ignore_invalid_snoop_crresp_writeunique = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITEUNIQUE} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1101};
      ignore_bins ignore_invalid_snoop_crresp_writelineunique = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITELINEUNIQUE} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1101};
      ignore_bins ignore_invalid_snoop_crresp_evict = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::EVICT} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1001,4'b1101,4'b1000};


      option.weight=1;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite_writeevict_disabled
    * This covergroup will be created when there is only one ACE-master and
    * minimum one or more than one ACE_LITE master in the system.
    * The bins in covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite_writeevict_disabled will be hit when a coherent transaction  is outstanding while a snoop transaction is outstanding on same port with overlapping address
    * The covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite_writeevict_disabled is applicable only for ACE Masters.The covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite_writeevict_disabled needs at least one ACE and one ACE_LITE master in the system.
    * Coverpoints:
    * snoop_xact_type:Coverpoint of svt_axi_snoop_transaction::snoop_xact_type for READONCE,CLEANSHARED,CLEANINVALID and MAKEINVALID snoop transactions recieved on master port . This excludes READSHARED,READCLEAN,READNOTSHAREDDIRTY,READUNIQUE,DVMMESSAGE,DVMCOMPLETE transactions
    * coherent_write_xact_type_generate_snoop:Coverpoint of svt_axi_transaction::coherent_xact_type for all coherent transactions initiated on write channel of master .This coverpoint includes only those transactions that     
    * generate snoop.This includes WRITEUNIQUE and WRITELINEUNIQUE transactions  
    * snoop_crresp_on_ace_port : coverpoint of cresp.
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.6.2
    *
    */

  covergroup trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite_writeevict_disabled;
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NO_WRITEEVICT_SNOOP_GENERATE
      snoop_xact_type : coverpoint master_snoop_xact_type { 
        bins snoop_readonce_xact   = {svt_axi_snoop_transaction::READONCE}; 
        bins snoop_cleanshared_xact   = {svt_axi_snoop_transaction::CLEANSHARED}; 
        bins snoop_cleaninvalid_xact   = {svt_axi_snoop_transaction::CLEANINVALID}; 
        bins snoop_makeinvalid_xact   = {svt_axi_snoop_transaction::MAKEINVALID}; 
        option.weight = 1; 
      }
       
       snoop_crresp_on_ace_port: coverpoint snoop_resp_ace_master[3:0] {
       bins cresp_0000 = {4'b0000};
       bins cresp_1000 = {4'b1000};
       bins cresp_0001 = {4'b0001};
       bins cresp_1001 = {4'b1001};
       bins cresp_0101 = {4'b0101};
       bins cresp_1101 = {4'b1101};    
       option.weight = 1;
    }
       snoop_crresp_wu : coverpoint snoop_resp_ace_master[4] {
         bins cresp_wasunique = {1'b1};
         bins cresp_wasnotunique = {1'b0};
         option.weight = 1;
    }    

       ace_concurrent_overlap_snoop_xact : cross snoop_xact_type,coherent_write_xact_type_gen_snoop,snoop_crresp_on_ace_port,snoop_crresp_wu{
       // Ignoring snoop_responses where is_shared is asserted and where data_transfer is asserted as recommended behaviour for MAKEINVALID is not tot transfer data 
       ignore_bins Ignore_invalid_rresp_ud_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::MAKEINVALID} &&
                                                 !binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b0000 };
      // Ignoring snoop_responses where is_shared bit is asserted or where data_transfer is asserted and pass_dirty is deasserted as CLEANINVALID will transfer data only when pass_dirty is asserted 
       ignore_bins ignore_invalid_rresp_ud_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::CLEANINVALID} &&
                                                 !binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b0000,4'b0101,4'b0001};

      ignore_bins ignore_invalid_snoop_crresp_writeunique = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITEUNIQUE} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1101};
      ignore_bins ignore_invalid_snoop_crresp_writelineunique = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITELINEUNIQUE} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1101};
      ignore_bins ignore_invalid_snoop_crresp_evict = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::EVICT} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1001,4'b1101,4'b1000};

      option.weight=1;
    }
    option.per_instance = 1;
  endgroup

/**
    * Covergroup: trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp
    * The bins in covergroup trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp will be hit when a coherent transaction  is outstanding while a snoop transaction is outstanding on same port with overlapping address
    * The covergroup trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp is applicable only for ACE Masters .The covergroup trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp needs at least two ACE masters in the system .
    * Coverpoints:
    * snoop_xact_type:Coverpoint of svt_axi_snoop_transaction::snoop_xact_type for all snoop transactions recieved on master port . This excludes DVMMESSAGE,DVMCOMPLETE transactions
    * coherent_write_xact_type_generate_snoop:Coverpoint of svt_axi_transaction::coherent_xact_type for all coherent transactions initiated on write channel of master .This coverpoint includes only those transactions that     * generate snoop.This includes WRITEUNIQUE and WRITELINEUNIQUE transactions  
    * snoop_crresp_on_ace_port :
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.6.2
    *
    */

 covergroup trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp;
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_SNOOP_GENERATE
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_NO_DVM
       
       snoop_crresp_on_ace_port: coverpoint snoop_resp_ace_master[3:0] {
       bins cresp_0000 = {4'b0000};
       bins cresp_1000 = {4'b1000};
       bins cresp_0001 = {4'b0001};
       bins cresp_1001 = {4'b1001};
       bins cresp_0101 = {4'b0101};
       bins cresp_1101 = {4'b1101};    
       option.weight = 1;
    }
       snoop_crresp_wu : coverpoint snoop_resp_ace_master[4] {
         bins cresp_wasunique = {1'b1};
         bins cresp_wasnotunique = {1'b0};
         option.weight = 1;
    }    

       ace_concurrent_overlap_snoop_xact : cross snoop_xact_type,coherent_write_xact_type_gen_snoop,snoop_crresp_on_ace_port,snoop_crresp_wu{
       // Ignoring snoop_responses where is_shared is asserted and where data_transfer is asserted as recommended behaviour for MAKEINVALID is not tot transfer data 
       ignore_bins Ignore_invalid_rresp_ud_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::MAKEINVALID} &&
                                                 !binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b0000 };
      // Ignoring snoop_responses where is_shared bit is asserted or where data_transfer is asserted and pass_dirty is deasserted as CLEANINVALID will transfer data only when pass_dirty is asserted 
       ignore_bins ignore_invalid_rresp_ud_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::CLEANINVALID} &&
                                                 !binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b0000,4'b0101};
      // ignoring snoop_responses where is_shared bit is asserted for READUNIQUE transactions 
      ignore_bins Ignore_invalid_rresp_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::READUNIQUE} &&
                                                 binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b1101,4'b1000,4'b1001};
      ignore_bins ignore_invalid_snoop_crresp_writeunique = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITEUNIQUE} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1101};
      ignore_bins ignore_invalid_snoop_crresp_writelineunique = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITELINEUNIQUE} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1101};
      option.weight=1;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite
    * This covergroup will be created when there is only one ACE-master and
    * minimum one or more than one ACE_LITE master in the system.
    * The bins in covergroup trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite will be hit when a coherent transaction  is outstanding while a snoop transaction is outstanding on same port with non overlapping address
    * The covergroup trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite is applicable only for ACE Masters .The covergroup trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite needs at least one ACE and one ACE_LITE master in the system.
    * Coverpoints:
    * snoop_xact_type:Coverpoint of svt_axi_snoop_transaction::snoop_xact_type for READONCE,CLEANSHARED,CLEANINVALID and MAKEINVALID snoop transactions recieved on master port . This excludes READSHARED,READCLEAN,READNOTSHAREDDIRTY,READUNIQUE,DVMMESSAGE,DVMCOMPLETE transactions
    * coherent_write_xact_type_generate_snoop:Coverpoint of svt_axi_transaction::coherent_xact_type for all coherent transactions initiated on write channel of master .This coverpoint includes only those transactions that     
    * generate snoop.This includes WRITEUNIQUE and WRITELINEUNIQUE transactions  
    * snoop_crresp_on_ace_port : Coverpoint of cresp.
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.6.2
    *
    */

  covergroup trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite;
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_SNOOP_GENERATE

       snoop_xact_type : coverpoint master_snoop_xact_type { 
       bins snoop_readonce_xact   = {svt_axi_snoop_transaction::READONCE}; 
       bins snoop_cleanshared_xact   = {svt_axi_snoop_transaction::CLEANSHARED}; 
       bins snoop_cleaninvalid_xact   = {svt_axi_snoop_transaction::CLEANINVALID}; 
       bins snoop_makeinvalid_xact   = {svt_axi_snoop_transaction::MAKEINVALID}; 
       option.weight = 1; 
    }
       
       snoop_crresp_on_ace_port: coverpoint snoop_resp_ace_master[3:0] {
       bins cresp_0000 = {4'b0000};
       bins cresp_1000 = {4'b1000};
       bins cresp_0001 = {4'b0001};
       bins cresp_1001 = {4'b1001};
       bins cresp_0101 = {4'b0101};
       bins cresp_1101 = {4'b1101};    
       option.weight = 1;
    }
       snoop_crresp_wu : coverpoint snoop_resp_ace_master[4] {
         bins cresp_wasunique = {1'b1};
         bins cresp_wasnotunique = {1'b0};
         option.weight = 1;
    }    

       ace_concurrent_overlap_snoop_xact : cross snoop_xact_type,coherent_write_xact_type_gen_snoop,snoop_crresp_on_ace_port,snoop_crresp_wu{
       // Ignoring snoop_responses where is_shared is asserted and where data_transfer is asserted as recommended behaviour for MAKEINVALID is not tot transfer data 
       ignore_bins Ignore_invalid_rresp_ud_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::MAKEINVALID} &&
                                                 !binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b0000 };
      // Ignoring snoop_responses where is_shared bit is asserted or where data_transfer is asserted and pass_dirty is deasserted as CLEANINVALID will transfer data only when pass_dirty is asserted 
       ignore_bins ignore_invalid_rresp_ud_sc_sd = binsof(snoop_xact_type) intersect {
                                                   svt_axi_snoop_transaction::CLEANINVALID} &&
                                                 !binsof(snoop_crresp_on_ace_port) intersect {
                                                   4'b0000,4'b0101};

      ignore_bins ignore_invalid_snoop_crresp_writeunique = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITEUNIQUE} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1101};
      ignore_bins ignore_invalid_snoop_crresp_writelineunique = binsof(coherent_write_xact_type_gen_snoop) intersect {svt_axi_transaction::WRITELINEUNIQUE} &&
                                                           binsof(snoop_crresp_on_ace_port) intersect {
                                                           4'b0101,4'b1101};
      option.weight=1;
    }
    option.per_instance = 1;
  endgroup

  /**
  *
  * Covergroup     : trans_cross_ace_acsnoop_acprot
  * 
  * Coverpoints:
  *
  * - snoop_xact_type:  Captures Snoop transaction
  * - snoop_prot:      Captures Snoop protection type
  * .
  *
  * Cross coverpoints:
  * - acsnoop_acprot : Crosses cover points
  *    snoop_xact_type and snoop_prot
  * .
  */

`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_acsnoop_acprot @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_PROT_TYPE

    acsnoop_acprot : cross snoop_xact_type, snoop_prot {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  /** 
   * This covergroup will be created when there is only one ACE-master and
   * minimum one or more than one ACE_LITE master in the system. 
   */
  covergroup trans_cross_ace_acsnoop_acprot_one_ace_acelite @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_ONE_ACE_ACELITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_PROT_TYPE

    acsnoop_acprot : cross snoop_xact_type, snoop_prot {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else

  covergroup trans_cross_ace_acsnoop_acprot_dvm_set @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_PROT_TYPE

    acsnoop_acprot : cross snoop_xact_type, snoop_prot {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /** 
   * This covergroup will be created when there is only one ACE-master and
   * minimum one or more than one ACE_LITE master in the system. 
   */
  covergroup trans_cross_ace_acsnoop_acprot_dvm_set_one_ace_acelite @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_SET_ONE_ACE_ACELITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_PROT_TYPE

    acsnoop_acprot : cross snoop_xact_type, snoop_prot {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_acsnoop_acprot_dvm_unset @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_PROT_TYPE

    acsnoop_acprot : cross snoop_xact_type, snoop_prot {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  /** 
   * This covergroup will be created when there is only one ACE-master and
   * minimum one or more than one ACE_LITE master in the system. 
   */
  covergroup trans_cross_ace_acsnoop_acprot_dvm_unset_one_ace_acelite @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_UNSET_ONE_ACE_ACELITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_PROT_TYPE

    acsnoop_acprot : cross snoop_xact_type, snoop_prot {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`endif

  /**
    *  Covergroup: trans_axi_snoop
    *
    *  Coverpoints:
    *  - ACVALID_to_ACREADY_Delay: Captures min, mid and max range of delays between signals acvalid and acready
    *  - ACVALID_to_CRVALID_Delay: Captures min, mid and max range of delays between signals acvalid and crvalid
    *  - CRVALID_to_CRREADY_Delay: Captures min, mid and max range of delays between signals crvalid and crready
    *  - ACVALID_to_prev_ACVALID_Delay: Captures min, mid and max range of delays between current and previous acvalid signals
    *  - ACVALID_before_ACREADY: Captures if ACVALID signal comes before ACREADY signal 
    *  - ACREADY_before_ACVALID: Captures if ACREADY signal comes before ACVALID signal
    *  - CRVALID_before_CRREADY: Captures if CRVALID signal comes before CRREADY signal 
    *  - CRREADY_before_CRVALID: Captures if CRREADY signal comes before CRVALID signal
    *  .
    */
  covergroup trans_axi_snoop @(cov_snoop_sample_event);
    option.per_instance = 1;
    ACVALID_to_ACREADY_Delay : coverpoint cov_ACVALID_to_ACREADY_Delay {
      bins acvalid_to_acready_delay_min = {0};
      bins acvalid_to_acready_delay_mid = {[1:(`SVT_AXI_MAX_ACREADY_DELAY/2)]};
      bins acvalid_to_acready_delay_max = {[(`SVT_AXI_MAX_ACREADY_DELAY/2)+1:$]};
      option.at_least = `SVT_AXI_trans_axi_snoop_ACVALID_to_ACREADY_Delay_COV_OPTION_AT_LEAST_VAL;
    }
    ACVALID_to_CRVALID_Delay : coverpoint cov_ACVALID_to_CRVALID_Delay { 
      bins acvalid_to_crvalid_delay_min = {[1:`MIN_UPPER_BOUND]};
      bins acvalid_to_crvalid_delay_mid = {[(`MIN_UPPER_BOUND+1):(`SVT_AXI_MAX_ACVALID_TO_CRVALID_DELAY/2)]};
      bins acvalid_to_crvalid_delay_max = {[(`SVT_AXI_MAX_ACVALID_TO_CRVALID_DELAY/2)+1:$]};
      option.at_least = `SVT_AXI_trans_axi_snoop_ACVALID_to_CRVALID_Delay_COV_OPTION_AT_LEAST_VAL;
    }
    CRVALID_to_CRREADY_Delay : coverpoint cov_CRVALID_to_CRREADY_Delay {
      bins crvalid_to_crready_delay_min = {0};
      bins crvalid_to_crready_delay_mid = {[1:(`SVT_AXI_MAX_CRREADY_DELAY/2)]};
      bins crvalid_to_crready_delay_max = {[(`SVT_AXI_MAX_CRREADY_DELAY/2)+1:$]};
      option.at_least = `SVT_AXI_trans_axi_snoop_CRVALID_to_CRREADY_Delay_COV_OPTION_AT_LEAST_VAL;
    }
    ACVALID_to_prev_ACVALID_Delay : coverpoint cov_ACVALID_to_prev_ACVALID_Delay {
      bins acvalid_to_prev_acvalid_delay_min = {1};
      bins acvalid_to_prev_acvalid_delay_mid = {[2:((`SVT_AXI_MAX_ACVALID_DELAY + `SVT_AXI_MAX_ACREADY_DELAY)/2)]};
      bins acvalid_to_prev_acvalid_delay_max = {[((`SVT_AXI_MAX_ACVALID_DELAY + `SVT_AXI_MAX_ACREADY_DELAY)/2)+1:$]};
      option.at_least = `SVT_AXI_trans_axi_snoop_ACVALID_to_prev_ACVALID_Delay_COV_OPTION_AT_LEAST_VAL;
    }
    /*CRVALID_to_prev_CRVALID_Delay : coverpoint cov_CRVALID_to_prev_CRVALID_Delay {
      bins crvalid_to_prev_crvalid_delay_min = {1};
      bins crvalid_to_prev_crvalid_mid = {[2:((`SVT_AXI_MAX_CRVALID_DELAY + `SVT_AXI_MAX_CRREADY_DELAY)/2)]};
      bins crvalid_to_prev_crvalid_max = {[((`SVT_AXI_MAX_CRVALID_DELAY + `SVT_AXI_MAX_CRREADY_DELAY)/2)+1:$]};
      option.at_least = `SVT_AXI_trans_axi_snoop_CRVALID_to_prev_CRVALID_Delay_COV_OPTION_AT_LEAST_VAL;
    }*/
    ACVALID_before_ACREADY: coverpoint cov_ACVALID_before_ACREADY {
      bins acvalid_before_acready = {1};
      option.at_least = `SVT_AXI_trans_axi_snoop_ACVALID_before_ACREADY_COV_OPTION_AT_LEAST_VAL;
    }
    ACREADY_before_ACVALID: coverpoint cov_ACREADY_before_ACVALID {
      bins acready_before_acvalid = {1};
      option.at_least = `SVT_AXI_trans_axi_snoop_ACREADY_before_ACVALID_COV_OPTION_AT_LEAST_VAL;
    }
    CRVALID_before_CRREADY: coverpoint cov_CRVALID_before_CRREADY {
      bins crvalid_before_crready = {1};
      option.at_least = `SVT_AXI_trans_axi_snoop_CRVALID_before_CRREADY_COV_OPTION_AT_LEAST_VAL;
    }
    CRREADY_before_CRVALID: coverpoint cov_CRREADY_before_CRVALID {
      bins crready_before_crvalid = {1};
      option.at_least = `SVT_AXI_trans_axi_snoop_CRREADY_before_CRVALID_COV_OPTION_AT_LEAST_VAL;
    }
  endgroup

/**
    *  Covergroup: trans_axi_snoop
    *
    *  Coverpoints:
    *  - ACWAKEUP_before_ACVALID_Delay: Captures min, mid and max range of delays between signals acwakeup to acvalid
    *  - ACWAKEUP_after_ACVALID_Delay: Captures min, mid and max range of delays between signals acvalid to acwakeup
    *  - ACWAKEUP_ACVALID_same_time: Captures delays of signals acwakeup and acvalid assertion same time
    *  - ACWAKEUP_to_prev_ACWAKEUP_Delay: Captures min, mid and max range of delays between signals acwakeup to previous acwakeup
    *  .
    */
  covergroup trans_axi_snoop_with_acwakeup @(cov_snoop_sample_event);
    option.per_instance = 1;
    ACWAKEUP_before_ACVALID_Delay : coverpoint cov_ACWAKEUP_before_ACVALID_Delay {
      bins acwakeup_before_acvalid_min = {`SVT_AXI_MIN_ACWAKEUP_ASSERT_DELAY};
      bins acwakeup_before_acvalid_mid = {[`SVT_AXI_MIN_ACWAKEUP_ASSERT_DELAY+1:(`SVT_AXI_MAX_ACWAKEUP_ASSERT_DELAY/2)]};
      bins acwakeup_before_acvalid_max = {[(`SVT_AXI_MAX_ACWAKEUP_ASSERT_DELAY/2)+1:`SVT_AXI_MAX_ACWAKEUP_ASSERT_DELAY]};
    }
    ACWAKEUP_after_ACVALID_Delay : coverpoint cov_ACWAKEUP_after_ACVALID_Delay {
      bins acwakeup_after_acvalid_min = {`SVT_AXI_MIN_ACWAKEUP_ASSERT_DELAY};
      bins acwakeup_after_acvalid_mid = {[`SVT_AXI_MIN_ACWAKEUP_ASSERT_DELAY+1:(`SVT_AXI_MAX_ACWAKEUP_ASSERT_DELAY/2)]};
      bins acwakeup_after_acvalid_max = {[(`SVT_AXI_MAX_ACWAKEUP_ASSERT_DELAY/2)+1:`SVT_AXI_MAX_ACWAKEUP_ASSERT_DELAY]};
    }
    ACWAKEUP_ACVALID_same_time : coverpoint cov_ACWAKEUP_ACVALID_same_time {
      bins acwakeup_acvalid_same_time = {0};
    }
     ACWAKEUP_to_prev_ACWAKEUP_Delay : coverpoint cov_ACWAKEUP_to_prev_ACWAKEUP_Delay {
      bins acwakeup_to_prev_acwakeup_delay_min = {2};
      bins acwakeup_to_prev_acwakeup_delay_mid = {[3:((`SVT_AXI_MAX_ACVALID_DELAY + `SVT_AXI_MAX_ACREADY_DELAY + `SVT_AXI_MAX_ACWAKEUP_ASSERT_DELAY)/3)]};
      bins acwakeup_to_prev_acwakeup_delay_max = {[((`SVT_AXI_MAX_ACVALID_DELAY + `SVT_AXI_MAX_ACREADY_DELAY + `SVT_AXI_MAX_ACWAKEUP_ASSERT_DELAY)/3)+1:$]};
     }
  endgroup

/**
    *  Covergroup: trans_axi_snoop
    *
    *  Coverpoints:
    *  - ACWAKEUP_toggle_Delay_idle_snoop_chan: Captures min, mid and max range of acwakeup toggle delay
    *  during idle period of snoop channel
    *  .
    */
  covergroup trans_axi_snoop_idle_chan_with_acwakeup @(cov_snoop_sample_event_for_idle_snoop_chan);
    ACWAKEUP_toggle_Delay_idle_snoop_chan : coverpoint cov_ACWAKEUP_toggle_Delay_idle_snoop_chan {
      bins acwakeup_after_acvalid_min = {cfg.acwakeup_toggle_min_delay_during_idle};
      bins acwakeup_after_acvalid_mid = {[(cfg.acwakeup_toggle_min_delay_during_idle+1):(cfg.acwakeup_toggle_max_delay_during_idle)/2]};
      bins acwakeup_after_acvalid_max = {[(cfg.acwakeup_toggle_max_delay_during_idle/2)+1:cfg.acwakeup_toggle_max_delay_during_idle]};
    }
  endgroup
  
/**
    *  Covergroup: trans_axi_snoop
    *
    *  Coverpoints:
    *  - AWAKEUP_before_ARVALID_Delay: Captures min, mid and max range of delays between signals awakeup to arvalid
    *  - AWAKEUP_after_ARVALID_Delay: Captures min, mid and max range of delays between signals arvalid to awakeup
    *  - AWAKEUP_ARVALID_same_time: Captures delays of signals awakeup and arvalid assertion same time
    *  - AWAKEUP_to_prev_AWAKEUP_Delay: Captures min, mid and max range of delays between signals awakeup to previous awakeup
    *  .
    */
 ////////////////////////////////

 covergroup trans_axi_awakeup @(cov_awakeup_sample_event); 
    option.per_instance = 1;
    AWAKEUP_before_ARVALID_Delay : coverpoint cov_AWAKEUP_before_ARVALID_Delay {
      bins awakeup_before_arvalid_min = {`SVT_AXI_MIN_AWAKEUP_ASSERT_DELAY};
      bins awakeup_before_arvalid_mid = {[`SVT_AXI_MIN_AWAKEUP_ASSERT_DELAY+1:(`SVT_AXI_MAX_AWAKEUP_ASSERT_DELAY/2)]};
      bins awakeup_before_arvalid_max = {[(`SVT_AXI_MAX_AWAKEUP_ASSERT_DELAY/2)+1:`SVT_AXI_MAX_AWAKEUP_ASSERT_DELAY]};
    }
    AWAKEUP_after_ARVALID_Delay : coverpoint cov_AWAKEUP_after_ARVALID_Delay {
      bins awakeup_after_arvalid_min = {`SVT_AXI_MIN_AWAKEUP_ASSERT_DELAY};
      bins awakeup_after_arvalid_mid = {[`SVT_AXI_MIN_AWAKEUP_ASSERT_DELAY+1:(`SVT_AXI_MAX_AWAKEUP_ASSERT_DELAY/2)]};
      bins awakeup_after_arvalid_max = {[(`SVT_AXI_MAX_AWAKEUP_ASSERT_DELAY/2)+1:`SVT_AXI_MAX_AWAKEUP_ASSERT_DELAY]};
    }
    AWAKEUP_ARVALID_same_time : coverpoint cov_AWAKEUP_ARVALID_same_time {
      bins awakeup_arvalid_same_time = {0};
    }
     AWAKEUP_to_prev_AWAKEUP_Delay : coverpoint cov_AWAKEUP_to_prev_AWAKEUP_Delay {
      bins awakeup_to_prev_awakeup_delay_min = {2};
   //   bins awakeup_to_prev_awakeup_delay_mid = {[3:((`SVT_AXI_MAX_ARVALID_DELAY + `SVT_AXI_MAX_ARREADY_DELAY + `SVT_AXI_MAX_AWAKEUP_ASSERT_DELAY)/3)]};
   //   bins awakeup_to_prev_awakeup_delay_max = {[((`SVT_AXI_MAX_ARVALID_DELAY + `SVT_AXI_MAX_ARREADY_DELAY + `SVT_AXI_MAX_AWAKEUP_ASSERT_DELAY)/3)+1:$]};
     }
  endgroup

/**
    *  Covergroup: trans_axi_snoop
    *
    *  Coverpoints:
    *  - AWAKEUP_toggle_Delay_idle_snoop_chan: Captures min, mid and max range of awakeup toggle delay
    *  during idle period of snoop channel
    *  .
    */
    covergroup trans_axi_snoop_idle_chan_with_awakeup
    @(cov_snoop_sample_event_for_awakeup_idle_snoop_chan);
    option.per_instance = 1;

      AWAKEUP_toggle_Delay_idle_snoop_chan : coverpoint cov_AWAKEUP_toggle_Delay_idle_snoop_chan {
        bins awakeup_after_arvalid_min = {cfg.awakeup_toggle_min_delay_during_idle};
        bins awakeup_after_arvalid_mid = {[(cfg.awakeup_toggle_min_delay_during_idle+1):(cfg.awakeup_toggle_max_delay_during_idle)/2]};
        bins awakeup_after_arvalid_max = {[(cfg.awakeup_toggle_max_delay_during_idle/2)+1:cfg.awakeup_toggle_max_delay_during_idle]};
      }
    endgroup

  /**
    *  Covergroup: signal_master_valid_ready_dependency
    *  The bins will get hit if signals are deassarted for N clock cycle mentioned by the user using port configuration parameter. 
    *  For Eg: The signal AWVALID has to remain deasserted for N clocks (user
    *  input) after wvalid is deasserted, then coverpoint AWVALID_WVALID_Dependency will get hit.
    *  In this case N value will be svt_axi_port_configuration::cov_num_clks_awvalid_wvalid_dependency.
    *          
    *  Coverpoints:
    *  - AWVALID_WVALID_Dependency: Will get hit if AWVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_awvalid_wvalid_dependency) after WVALID is deasserted.
    *  - AWVALID_RREADY_Dependency: Will get hit if AWVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_awvalid_rready_dependency) after RREADY is deasserted.
    *  - AWVALID_BREADY_Dependency: Will get hit if AWVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_awvalid_bready_dependency) after BREADY is deasserted.
    *  - WVALID_AWVALID_Dependency: Will get hit if WVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_wvalid_awvalid_dependency) after AWVALID is deasserted.
    *  - WVALID_RREADY_Dependency: Will get hit if WVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_wvalid_rready_dependency) after RREADY is deasserted.
    *  - WVALID_BREADY_Dependency: Will get hit if WVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_wvalid_bready_dependency) after BREADY is deasserted.
    *  - RREADY_AWVALID_Dependency: Will get hit if RREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_rready_awvalid_dependency) after AWVALID is deasserted.
    *  - RREADY_WVALID_Dependency: Will get hit if RREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_rready_wvalid_dependency) after WVALID is deasserted.
    *  - RREADY_BREADY_Dependency: Will get hit if RREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_rready_bready_dependency) after BREADY is deasserted.
    *  - BREADY_AWVALID_Dependency: Will get hit if BREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_bready_awvalid_dependency) after AWVALID is deasserted.
    *  - BREADY_WVALID_Dependency: Will get hit if BREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_bready_wvalid_dependency) after WVALID is deasserted.
    *  - BREADY_RREADY_Dependency: Will get hit if BREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_bready_rready_dependency) after RREADY is deasserted.
    *  .
    */
  covergroup signal_master_valid_ready_dependency @(cov_signal_dependency_event);
    AWVALID_WVALID_Dependency : coverpoint cov_awvalid_wvalid {
      bins AWVALID_and_WVALID = {1};
      option.at_least = 1;
    }
    AWVALID_RREADY_Dependency : coverpoint cov_awvalid_rready {
      bins AWVALID_and_RREADY = {1};
      option.at_least = 1;
    }
    AWVALID_BREADY_Dependency : coverpoint cov_awvalid_bready {
      bins AWVALID_and_BREADY = {1};
      option.at_least = 1;
    }
    WVALID_AWVALID_Dependency : coverpoint cov_wvalid_awvalid {
      bins WVALID_and_AWVALID = {1};
      option.at_least = 1;
    }
    WVALID_RREADY_Dependency : coverpoint cov_wvalid_rready {
      bins AWVALID_and_RREADY = {1};
      option.at_least = 1;
    }
    WVALID_BREADY_Dependency : coverpoint cov_wvalid_bready {
      bins WVALID_and_BREADY = {1};
      option.at_least = 1;
    }
    RREADY_AWVALID_Dependency : coverpoint cov_rready_awvalid {
      bins RREADY_and_AWVALID = {1};
      option.at_least = 1;
    }
    RREADY_WVALID_Dependency : coverpoint cov_rready_wvalid {
      bins RREADY_and_WVALID = {1};
      option.at_least = 1;
    }
    RREADY_BREADY_Dependency : coverpoint cov_rready_bready {
      bins RREADY_and_BREADY = {1};
      option.at_least = 1;
    }
    BREADY_AWVALID_Dependency : coverpoint cov_bready_awvalid {
      bins BREADY_and_AWVALID = {1};
      option.at_least = 1;
    }
    BREADY_WVALID_Dependency : coverpoint cov_bready_wvalid {
      bins BREADY_and_WVALID = {1};
      option.at_least = 1;
    }
    BREADY_RREADY_Dependency : coverpoint cov_bready_rready {
      bins BREADY_and_RREADY = {1};
      option.at_least = 1;
    }
    option.per_instance = 1;
  endgroup

  /**
    *  Covergroup: signal_slave_valid_ready_dependency
    *  The bins will get hit if signals are deassarted for N clock cycle mentioned by the user using port configuration parameter. 
    *  For Eg: The signal WREADY has to remain deasserted for N clocks (user
    *  input) after arready is deasserted, then coverpoint WREADY_ARREADY_Dependency will get hit.
    *  In this case N value will be svt_axi_port_configuration::cov_num_clks_wready_arready_dependency.
    *          
    *  Coverpoints:
    *  - WREADY_ARREADY_Dependency : Will get hit if WREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_wready_arready_dependency) after ARREADY is deasserted.
    *  - WREADY_RVALID_Dependency : Will get hit if WREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_wready_rvalid_dependency) after RVALID is deasserted.
    *  - WREADY_BVALID_Dependency : Will get hit if WREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_wready_bvalid_dependency) after BVALID is deasserted.
    *  - ARREADY_WREADY_Dependency : Will get hit if ARREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_arready_wready_dependency) after WREADY is deasserted.
    *  - ARREADY_RVALID_Dependency : Will get hit if ARREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_arready_rvalid_dependency) after RVALID is deasserted.
    *  - ARREADY_BVALID_Dependency : Will get hit if ARREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_arready_bvalid_dependency) after BVALID is deasserted.
    *  - RVALID_ARREADY_Dependency : Will get hit if RVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_rvalid_arready_dependency) after ARREADY is deasserted.
    *  - RVALID_WREADY_Dependency : Will get hit if RVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_rvalid_wready_dependency) after WREADY is deasserted.
    *  - RVALID_BVALID_Dependency : Will get hit if RVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_rvalid_bvalid_dependency) after BVALID is deasserted.
    *  - BVALID_ARREADY_Dependency : Will get hit if BVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_bvalid_arready_dependency) after ARREADY is deasserted.
    *  - BVALID_WREADY_Dependency : Will get hit if BVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_bvalid_wready_dependency) after WREADY is deasserted.
    *  - BVALID_RVALID_Dependency : Will get hit if BVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_bvalid_rvalid_dependency) after RVALID is deasserted.
    *  .
    */

  covergroup signal_slave_valid_ready_dependency @(cov_signal_slave_dependency_event);

    WREADY_ARREADY_Dependency : coverpoint cov_wready_arready {
      bins WREADY_and_ARREADY = {1};
      option.at_least = 1;
    }
    WREADY_RVALID_Dependency : coverpoint cov_wready_rvalid {
      bins WREADY_and_RVALID = {1};
      option.at_least = 1;
    }
    WREADY_BVALID_Dependency : coverpoint cov_wready_bvalid {
      bins WREADY_and_BVALID = {1};
      option.at_least = 1;
    }
    ARREADY_WREADY_Dependency : coverpoint cov_arready_wready {
      bins ARREADY_and_WREADY = {1};
      option.at_least = 1;
    }
    ARREADY_RVALID_Dependency : coverpoint cov_arready_rvalid{
      bins ARREADY_and_RVALID = {1};
      option.at_least = 1;
    }
    ARREADY_BVALID_Dependency : coverpoint cov_arready_bvalid {
      bins ARREADY_and_BVALID = {1};
      option.at_least = 1;
    }
    RVALID_ARREADY_Dependency : coverpoint cov_rvalid_arready {
      bins RVALID_and_ARREADY = {1};
      option.at_least = 1;
    }
    RVALID_WREADY_Dependency : coverpoint cov_rvalid_wready {
      bins RVALID_and_WREADY = {1};
      option.at_least = 1;
    }
    RVALID_BVALID_Dependency : coverpoint cov_rvalid_bvalid {
      bins RVALID_and_BVALID = {1};
      option.at_least = 1;
    }
    BVALID_ARREADY_Dependency : coverpoint cov_bvalid_arready {
      bins BVALID_and_ARREADY = {1};
      option.at_least = 1;
    }
    BVALID_WREADY_Dependency : coverpoint cov_bvalid_wready {
      bins BVALID_and_WREADY = {1};
      option.at_least = 1;
    }
    BVALID_RVALID_Dependency : coverpoint cov_bvalid_rvalid {
      bins BVALID_and_RVALID = {1};
      option.at_least = 1;
    }
    
    option.per_instance = 1;
  endgroup

  /**
    *  Covergroup: signal_master_slave_valid_ready_dependency
    *  The bins will get hit if signals are deassarted for N clock cycle mentioned by the user using port configuration parameter. 
    *  For Eg: The signal AWVALID has to remain deasserted for N clocks (user
    *  input) after AWREADY is deasserted, then coverpoint AWVALID_AWREADY_Dependency will get hit.
    *  In this case N value will be svt_axi_port_configuration::cov_num_clks_awvalid_awready_dependency.
    *          
    *  Coverpoints:
    *  - AWVALID_AWREADY_Dependency : Will get hit if AWVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_awvalid_awready_dependency) after AWREADY is deasserted.
    *  - AWVALID_WREADY_Dependency : Will get hit if AWVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_awvalid_wready_dependency) after WREADY is deasserted.
    *  - AWVALID_RVALID_Dependency : Will get hit if AWVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_awvalid_rvalid_dependency) after RVALID is deasserted.
    *  - AWVALID_BVALID_Dependency : Will get hit if AWVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_awvalid_bvalid_dependency) after BVALID is deasserted.
    *  - WVALID_AWREADY_Dependency : Will get hit if WVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_wvalid_awready_dependency) after AWREADY is deasserted.
    *  - WVALID_WREADY_Dependency : Will get hit if WVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_wvalid_wready_dependency) after WREADY is deasserted.
    *  - WVALID_RVALID_Dependency : Will get hit if WVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_wvalid_rvalid_dependency) after RVALID is deasserted.
    *  - WVALID_BVALID_Dependency : Will get hit if WVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_wvalid_bvalid_dependency) after BVALID is deasserted.
    *  - RREADY_AWREADY_Dependency : Will get hit if RREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_rready_awready_dependency) after AWREADY is deasserted.
    *  - RREADY_WREADY_Dependency : Will get hit if RREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_rready_wready_dependency) after WREADY is deasserted.
    *  - RREADY_RVALID_Dependency : Will get hit if RREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_rready_rvalid_dependency) after RVALID is deasserted.
    *  - RREADY_BVALID_Dependency : Will get hit if RREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_rready_bvalid_dependency) after BVALID is deasserted.
    *  - BREADY_AWREADY_Dependency : Will get hit if BREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_bready_awready_dependency) after AWREADY is deasserted.
    *  - BREADY_WREADY_Dependency : Will get hit if BREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_bready_wready_dependency) after WREADY is deasserted.
    *  - BREADY_RVALID_Dependency : Will get hit if BREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_bready_rvalid_dependency) after RVALID is deasserted.
    *  - BREADY_BVALID_Dependency : Will get hit if BREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_bready_bvalid_dependency) after BVALID is deasserted.
    *  .
    */
  covergroup signal_master_slave_valid_ready_dependency @(cov_signal_master_slave_dependency_event);

    AWVALID_AWREADY_Dependency : coverpoint cov_awvalid_awready {
      bins AWVALID_and_AWREADY = {1};
      option.at_least = 1;
    }
    AWVALID_WREADY_Dependency : coverpoint cov_awvalid_wready {
      bins AWVALID_and_WREADY = {1};
      option.at_least = 1;
    }
    AWVALID_RVALID_Dependency : coverpoint cov_awvalid_rvalid {
      bins AWVALID_and_RVALID = {1};
      option.at_least = 1;
    }
    AWVALID_BVALID_Dependency : coverpoint cov_awvalid_bvalid {
      bins AWVALID_and_BVALID = {1};
      option.at_least = 1;
    }
    WVALID_AWREADY_Dependency : coverpoint cov_wvalid_awready {
      bins WVALID_and_AWREADY = {1};
      option.at_least = 1;
    }
    WVALID_WREADY_Dependency : coverpoint cov_wvalid_wready {
      bins WVALID_and_WREADY = {1};
      option.at_least = 1;
    }
    WVALID_RVALID_Dependency : coverpoint cov_wvalid_rvalid {
      bins WVALID_and_RVALID = {1};
      option.at_least = 1;
    }
    WVALID_BVALID_Dependency : coverpoint cov_wvalid_bvalid {
      bins WVALID_and_BVALID = {1};
      option.at_least = 1;
    }

    RREADY_AWREADY_Dependency : coverpoint cov_rready_awready {
      bins RREADY_and_AWREADY = {1};
      option.at_least = 1;
    }
    RREADY_WREADY_Dependency : coverpoint cov_rready_wready {
      bins RREADY_and_WREADY = {1};
      option.at_least = 1;
    }
    RREADY_RVALID_Dependency : coverpoint cov_rready_rvalid {
      bins RREADY_and_RVALID = {1};
      option.at_least = 1;
    }
    RREADY_BVALID_Dependency : coverpoint cov_rready_bvalid {
      bins RREADY_and_BVALID = {1};
      option.at_least = 1;
    }
    BREADY_AWREADY_Dependency : coverpoint cov_bready_awready {
      bins BREADY_and_AWREADY = {1};
      option.at_least = 1;
    }
    BREADY_WREADY_Dependency : coverpoint cov_bready_wready {
      bins BREADY_and_WREADY = {1};
      option.at_least = 1;
    }
    BREADY_RVALID_Dependency : coverpoint cov_bready_rvalid {
      bins BREADY_and_RVALID = {1};
      option.at_least = 1;
    }
    BREADY_BVALID_Dependency : coverpoint cov_bready_bvalid {
      bins BREADY_and_BVALID = {1};
      option.at_least = 1;
    }
    option.per_instance = 1;
  endgroup

  /**
    *  Covergroup: signal_slave_master_valid_ready_dependency
    *  The bins will get hit if signals are deassarted for N clock cycle mentioned by the user using port configuration parameter. 
    *  For Eg: The signal AWREADY has to remain deasserted for N clocks (user
    *  input) after AWVALID is deasserted, then coverpoint AWREADY_AWVALID_Dependency will get hit.
    *  In this case N value will be svt_axi_port_configuration::cov_num_clks_awvalid_awready_dependency.
    *          
    *  Coverpoints:
    *  - AWREADY_AWVALID_Dependency : Will get hit if AWREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_awready_and_awvalid_dependency) after AWVALIDis deasserted.
    *  - AWREADY_WVALID_Dependency  : Will get hit if AWREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_awready_and_wvalid_dependency) after WVALID is deasserted.
    *  - AWREADY_RVALID_Dependency  : Will get hit if AWREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_awready_and_rvalid_dependency) after RVALID is deasserted.
    *  - AWREADY_BVALID_Dependency  : Will get hit if AWREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_awready_and_bvalid_dependency) after BVALID is deasserted.
    *  - WREADY_AWVALID_Dependency  : Will get hit if WREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_wready_and_awvalid_dependency) after AWVALID is deasserted.
    *  - WREADY_WVALID_Dependency   : Will get hit if WREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_wready_and_wvalid_dependency) after WVALID is deasserted.
    *  - WREADY_RREADY_Dependency   : Will get hit if WREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_wready_and_rready_dependency) after RREADY is deasserted.
    *  - WREADY_BREADY_Dependency   : Will get hit if WREADY remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_wready_and_bready_dependency) after BREADY is deasserted.
    *  - RVALID_AWREADY_Dependency  : Will get hit if RVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_rvalid_and_awready_dependency) after AWREADY is deasserted.
    *  - RVALID_WREADY_Dependency   : Will get hit if RVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_rvalid_and_wready_dependency) after WREADY is deasserted.
    *  - RVALID_RREADY_Dependency   : Will get hit if RVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_rvalid_and_rready_dependency) after RREADY is deasserted.
    *  - RVALID_BREADY_Dependency   : Will get hit if RVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_rvalid_and_bready_dependency) after BREADY is deasserted.
    *  - BVALID_AWREADY_Dependency  : Will get hit if BVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_bvalid_and_awready_dependency) afterAWREADY is deasserted.
    *  - BVALID_WREADY_Dependency   : Will get hit if BVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_bvalid_and_wready_dependency) after WREADY is deasserted.
    *  - BVALID_RREADY_Dependency   : Will get hit if BVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_bvalid_and_rready_dependency) after RREADY is deasserted.
    *  - BVALID_BREADY_Dependency   : Will get hit if BVALID remains deasserted for N clock cycles(N = svt_axi_port_configuration::cov_num_clks_bvalid_and_bready_dependency) after BREADY is deasserted.
    *  .
    */
  covergroup signal_slave_master_valid_ready_dependency @(cov_signal_slave_master_dependency_event);

    AWREADY_AWVALID_Dependency : coverpoint cov_awready_and_awvalid {
      bins AWREADY_and_AWVALID = {1};
      option.at_least = 1;
    }
    AWREADY_WVALID_Dependency : coverpoint cov_awready_and_wvalid {
      bins AWREADY_and_WVALID = {1};
      option.at_least = 1;
    }
    AWREADY_RVALID_Dependency : coverpoint cov_awready_and_rvalid {
      bins AWREADY_and_RVALID = {1};
      option.at_least = 1;
    }
    AWREADY_BVALID_Dependency : coverpoint cov_awready_and_bvalid {
      bins AWREADY_and_BVALID = {1};
      option.at_least = 1;
    }
    WREADY_AWVALID_Dependency : coverpoint cov_wready_and_awvalid {
      bins WREADY_and_AWVALID = {1};
      option.at_least = 1;
    }
    WREADY_WVALID_Dependency  : coverpoint cov_wready_and_wvalid  {
      bins WREADY_and_WVALID = {1};
      option.at_least = 1;
    }
    WREADY_RREADY_Dependency  : coverpoint cov_wready_and_rready  {
      bins WREADY_and_RREADY = {1};
      option.at_least = 1;
    }
    WREADY_BREADY_Dependency  : coverpoint cov_wready_and_bready  {
      bins WREADY_and_BREADY = {1};
      option.at_least = 1;
    }

    RVALID_AWREADY_Dependency : coverpoint cov_rvalid_and_awready {
      bins RVALID_and_AWREADY = {1};
      option.at_least = 1;
    }
    RVALID_WREADY_Dependency  : coverpoint cov_rvalid_and_wready  {
      bins RVALID_and_WREADY = {1};
      option.at_least = 1;
    }
    RVALID_RREADY_Dependency  : coverpoint cov_rvalid_and_rready  {
      bins RVALID_and_RREADY = {1};
      option.at_least = 1;
    }
    RVALID_BREADY_Dependency  : coverpoint cov_rvalid_and_bready  {
      bins RVALID_and_BREADY = {1};
      option.at_least = 1;
    }
    BVALID_AWREADY_Dependency : coverpoint cov_bvalid_and_awready {
      bins BVALID_and_AWREADY = {1};
      option.at_least = 1;
    }
    BVALID_WREADY_Dependency  : coverpoint cov_bvalid_and_wready  {
      bins BVALID_and_WREADY = {1};
      option.at_least = 1;
    }
    BVALID_RREADY_Dependency  : coverpoint cov_bvalid_and_rready  {
      bins BVALID_and_RREADY = {1};
      option.at_least = 1;
    }
    BVALID_BREADY_Dependency  : coverpoint cov_bvalid_and_bready  {
      bins BVALID_and_BREADY = {1};
      option.at_least = 1;
    }
    option.per_instance = 1;
  endgroup

  /**
    *  Covergroup: trans_axi_snoop_data_phase
    *
    *  Coverpoints:
    *  - CDVALID_to_prev_CDVALID_Delay
    *  - CDVALID_to_CDREADY_Delay
    *  - CDVALID_before_CDREADY: Captures if CDVALID signal comes before CDREADY signal 
    *  - CDREADY_before_CDVALID: Captures if CDREADY signal comes before CDVALID signal
    *  .
    */
  covergroup trans_axi_snoop_data_phase @(cov_snoop_per_beat_sample_event);
    option.per_instance = 1;
    CDVALID_to_prev_CDVALID_Delay : coverpoint cov_CDVALID_to_prev_CDVALID_Delay {
      bins cdvalid_to_prev_cdvalid_delay_min = {1};
      bins cdvalid_to_prev_cdvalid_delay_mid = {[2:((`SVT_AXI_MAX_CDVALID_DELAY + `SVT_AXI_MAX_CDREADY_DELAY)/2)]};
      bins cdvalid_to_prev_cdvalid_delay_max = {[((`SVT_AXI_MAX_CDVALID_DELAY + `SVT_AXI_MAX_CDREADY_DELAY)/2)+1:$]};
      option.at_least = `SVT_AXI_trans_axi_snoop_CDVALID_to_prev_CDVALID_Delay_COV_OPTION_AT_LEAST_VAL;
    }
    CDVALID_to_CDREADY_Delay : coverpoint cov_CDVALID_to_CDREADY_Delay {
      bins cdvalid_to_cdready_delay_min = {0};
      bins cdvalid_to_cdready_delay_mid = {[1:(`SVT_AXI_MAX_CDREADY_DELAY/2)]};
      bins cdvalid_to_cdready_delay_max = {[(`SVT_AXI_MAX_CDREADY_DELAY/2)+1:$]};
      option.at_least = `SVT_AXI_trans_axi_snoop_CDVALID_to_CDREADY_Delay_COV_OPTION_AT_LEAST_VAL;
    }
    CDVALID_before_CDREADY: coverpoint cov_CDVALID_before_CDREADY {
      bins cdvalid_before_cdready = {1};
      option.at_least = `SVT_AXI_trans_axi_snoop_CDVALID_before_CDREADY_COV_OPTION_AT_LEAST_VAL;
    }
    CDREADY_before_CDVALID: coverpoint cov_CDREADY_before_CDVALID {
      bins cdready_before_cdvalid = {1};
      option.at_least = `SVT_AXI_trans_axi_snoop_CDREADY_before_CDVALID_COV_OPTION_AT_LEAST_VAL;
    }
  endgroup

  /**
  *
  * Covergroup     : trans_cross_ace_acsnoop_crresp
  * 
  * Coverpoints:
  *
  * - snoop_xact_type:  Captures Snoop transaction
  * - snoop_crresp:      Captures Snoop response type
  * .
  *
  * Cross coverpoints:
  * - acsnoop_crresp : Crosses cover points
  *    snoop_xact_type and snoop_crresp
  * .
  *
  */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_acsnoop_crresp @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_RRESP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WASUNIQUE_SNOOP_RRESP_TYPE

    acsnoop_crresp : cross snoop_xact_type, snoop_crresp {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_IGNORE_BINS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CRRESP_IGNORE_BINS
    }

    acsnoop_crresp_wasunique : cross snoop_xact_type, snoop_crresp_wu {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_IGNORE_BINS
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /** 
   * This covergroup will be created when there is only one ACE-master and
   * minimum one or more than one ACE_LITE master in the system. 
   */
  covergroup trans_cross_ace_acsnoop_crresp_one_ace_acelite @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_ONE_ACE_ACELITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_RRESP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WASUNIQUE_SNOOP_RRESP_TYPE

    acsnoop_crresp : cross snoop_xact_type, snoop_crresp {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_IGNORE_BINS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CRRESP_IGNORE_BINS
    }

    acsnoop_crresp_wasunique : cross snoop_xact_type, snoop_crresp_wu {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_IGNORE_BINS
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else
  covergroup trans_cross_ace_acsnoop_crresp_dvm_unset @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_RRESP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WASUNIQUE_SNOOP_RRESP_TYPE

    acsnoop_crresp : cross snoop_xact_type, snoop_crresp {
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CRRESP_IGNORE_BINS 
    }

    acsnoop_crresp_wasunique : cross snoop_xact_type, snoop_crresp_wu {
    }
    option.per_instance = 1;
  endgroup

  /** 
   * This covergroup will be created when there is only one ACE-master and
   * minimum one or more than one ACE_LITE master in the system. 
   */
  covergroup trans_cross_ace_acsnoop_crresp_dvm_unset_one_ace_acelite @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_UNSET_ONE_ACE_ACELITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_RRESP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WASUNIQUE_SNOOP_RRESP_TYPE

    acsnoop_crresp : cross snoop_xact_type, snoop_crresp {
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CRRESP_IGNORE_BINS 
    }

    acsnoop_crresp_wasunique : cross snoop_xact_type, snoop_crresp_wu {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup


  covergroup trans_cross_ace_acsnoop_crresp_dvm_set @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_RRESP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WASUNIQUE_SNOOP_RRESP_TYPE

    acsnoop_crresp : cross snoop_xact_type, snoop_crresp {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CRRESP_IGNORE_BINS
    }

    acsnoop_crresp_wasunique : cross snoop_xact_type, snoop_crresp_wu {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /** 
   * This covergroup will be created when there is only one ACE-master and
   * minimum one or more than one ACE_LITE master in the system. 
   */
  covergroup trans_cross_ace_acsnoop_crresp_dvm_set_one_ace_acelite @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_SET_ONE_ACE_ACELITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_RRESP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WASUNIQUE_SNOOP_RRESP_TYPE

    acsnoop_crresp : cross snoop_xact_type, snoop_crresp {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CRRESP_IGNORE_BINS
    }

    acsnoop_crresp_wasunique : cross snoop_xact_type, snoop_crresp_wu {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif
 /**
  *
  * Covergroup     : trans_cross_ace_acdvmmessage_acdvmresp
  * 
  * Coverpoints:
  *
  * - acdvm_message_type : Captures DVM message on acaddr[14:12]
  *
  * - acdvm_resp : Capture DVM response on crresp,
  *                accept = 5'b00000 and reject = 5'b00010
  * .
  *
  * Cross coverpoints:
  * - acdvmmessage_acdvmresp  : Crosses cover points acdvm_message_type and acdvm_resp
  * .
  */

  covergroup trans_cross_ace_acdvmmessage_acdvmresp @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVMMESSAGE_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_DVM_RESPONSE_TYPE
     acdvmmessage_acdvmresp : cross acdvm_message_type ,acdvm_resp {
        ignore_bins Ignore_dvm_hint_msg_resp = (binsof (acdvm_message_type) intersect {3'b110}) &&
                                               (binsof (acdvm_resp) intersect {5'b00010});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup


  /**
  * 
  * Covergroup     : trans_cross_ace_awsnoop_awburst
  * 
  * Coverpoints:
  *
  * - coherent_write_xact_type:  Captures coherent write transaction
  * - burst_type: Captures transaction burst type
  * .
  * Cross coverpoints:
  * - awsnoop_awburst_awlen : Crosses cover points
  *    coherent_write_xact_type and burst_type
  * .
  */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF 
  covergroup trans_cross_ace_awsnoop_awburst (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awburst : cross coherent_write_xact_type, burst_type, slave_port_id {

      ignore_bins Ignore_invalid_fixed   =  binsof(burst_type.fixed_burst) &&
                                                binsof(coherent_write_xact_type) intersect {
                                                svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,
                                                svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) &&
                                                (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER});
 `endif

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_awsnoop_not_ace_lite_no_barrier_no_writeevict_awburst_axi3_ace (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    awsnoop_awburst : cross coherent_write_xact_type, burst_type , slave_port_id{

      ignore_bins Ignore_invalid_fixed   =  binsof(burst_type.fixed_burst) &&
                                                binsof(coherent_write_xact_type) intersect {
                                                svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,
                                                svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) &&
                                                (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER});
 `endif

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_ace_awsnoop_not_ace_lite_no_barrier_writeevict_awburst_axi3_ace(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    awsnoop_awburst : cross coherent_write_xact_type, burst_type , slave_port_id{

      ignore_bins Ignore_invalid_fixed   =  binsof(burst_type.fixed_burst) &&
                                                binsof(coherent_write_xact_type) intersect {
                                                svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,
                                                svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) &&
                                                (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER});
 `endif

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_ace_awsnoop_not_ace_lite_barrier_no_writeevict_awburst_axi3_ace(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    awsnoop_awburst : cross coherent_write_xact_type, burst_type , slave_port_id{

      ignore_bins Ignore_invalid_fixed   =  binsof(burst_type.fixed_burst) &&
                                                binsof(coherent_write_xact_type) intersect {
                                                svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,
                                                svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) &&
                                                (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER});
 `endif

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_ace_awsnoop_not_ace_lite_barrier_writeevict_awburst_axi3_ace(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    awsnoop_awburst : cross coherent_write_xact_type, burst_type , slave_port_id{

      ignore_bins Ignore_invalid_fixed   =  binsof(burst_type.fixed_burst) &&
                                                binsof(coherent_write_xact_type) intersect {
                                                svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,
                                                svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) &&
                                                (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER});
 `endif

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_ace_awsnoop_ace_lite_no_barrier_awburst_axi3_ace(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    awsnoop_awburst : cross coherent_write_xact_type, burst_type , slave_port_id{

      ignore_bins Ignore_invalid_fixed   =  binsof(burst_type.fixed_burst) &&
                                                binsof(coherent_write_xact_type) intersect {
                                                svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,
                                                svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) &&
                                                (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER});
 `endif

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_ace_awsnoop_ace_lite_barrier_awburst_axi3_ace(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    awsnoop_awburst : cross coherent_write_xact_type, burst_type , slave_port_id{

      ignore_bins Ignore_invalid_fixed   =  binsof(burst_type.fixed_burst) &&
                                                binsof(coherent_write_xact_type) intersect {
                                                svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,
                                                svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT};
`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) &&
                                                (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER});
 `endif

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  /**
  *  Covergroup     : trans_cross_ace_awsnoop_awlen
  *
  * Coverpoints:
  *
  * - coherent_write_xact_type:  Captures coherent write transaction
  * - burst_length: Captures transaction burst length
  * .
  * Cross coverpoints:
  * - awsnoop_awlen : Crosses cover points
  *    coherent_write_xact_type and burst_length
  * .
  */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF 

  covergroup trans_cross_ace_awsnoop_awlen (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awlen : cross coherent_write_xact_type, burst_length, slave_port_id {

      ignore_bins Ignore_invalid_length_all   =  binsof(burst_length) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT};
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ignore_non_power_of_2_length when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3],[5:7]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`else
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3],[5:7],[9:15]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`endif
      ignore_bins Ignore_invalid_length_above_16   =  binsof(coherent_write_xact_type) intersect {
                                                        svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK} &&
                                                        binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};                                             
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF 
  covergroup trans_cross_ace_awsnoop_not_ace_lite_no_barrier_no_writeevict_awlen_ace (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    awsnoop_awlen : cross coherent_write_xact_type, burst_length , slave_port_id{

      ignore_bins Ignore_invalid_length_all   =  binsof(burst_length) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT};
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ignore_non_power_of_2_length when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3],[5:7]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`else
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3],[5:7],[9:15]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`endif
      ignore_bins Ignore_invalid_length_above_16   =  binsof(coherent_write_xact_type) intersect {
                                                        svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK} &&
                                                        binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};                                             
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_no_barrier_writeevict_awlen_ace (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    awsnoop_awlen : cross coherent_write_xact_type, burst_length , slave_port_id{

      ignore_bins Ignore_invalid_length_all   =  binsof(burst_length) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT};
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ignore_non_power_of_2_length when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3],[5:7]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`else
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3],[5:7],[9:15]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`endif
      ignore_bins Ignore_invalid_length_above_16   =  binsof(coherent_write_xact_type) intersect {
                                                        svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK} &&
                                                        binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};                                             
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_barrier_no_writeevict_awlen_ace (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    awsnoop_awlen : cross coherent_write_xact_type, burst_length , slave_port_id{

      ignore_bins Ignore_invalid_length_all   =  binsof(burst_length) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT};
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ignore_non_power_of_2_length when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3],[5:7]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`else
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3],[5:7],[9:15]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`endif
      ignore_bins Ignore_invalid_length_above_16   =  binsof(coherent_write_xact_type) intersect {
                                                        svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK} &&
                                                        binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};                                             
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_barrier_writeevict_awlen_ace (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    awsnoop_awlen : cross coherent_write_xact_type, burst_length , slave_port_id{

      ignore_bins Ignore_invalid_length_all   =  binsof(burst_length) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT};
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ignore_non_power_of_2_length when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3],[5:7]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`else
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3],[5:7],[9:15]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`endif
      ignore_bins Ignore_invalid_length_above_16   =  binsof(coherent_write_xact_type) intersect {
                                                        svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK} &&
                                                        binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};                                             
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_ace_lite_no_barrier_awlen_ace (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    awsnoop_awlen : cross coherent_write_xact_type, burst_length , slave_port_id{

      ignore_bins Ignore_invalid_length_all   =  binsof(burst_length) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT};
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ignore_non_power_of_2_length when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3],[5:7]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`else
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3],[5:7],[9:15]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`endif
      ignore_bins Ignore_invalid_length_above_16   =  binsof(coherent_write_xact_type) intersect {
                                                        svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK} &&
                                                        binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};                                             
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_ace_lite_barrier_awlen_ace (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    awsnoop_awlen : cross coherent_write_xact_type, burst_length , slave_port_id{

      ignore_bins Ignore_invalid_length_all   =  binsof(burst_length) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT};
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ignore_non_power_of_2_length when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3],[5:7]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`else
      ignore_bins Ignore_non_power_of_2_length = binsof(burst_length) intersect {[2:3],[5:7],[9:15]} &&
                                                 binsof(coherent_write_xact_type) intersect 
                                                      {svt_axi_transaction::WRITEEVICT};
`endif
      ignore_bins Ignore_invalid_length_above_16   =  binsof(coherent_write_xact_type) intersect {
                                                        svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK} &&
                                                        binsof(burst_length) intersect {[`SVT_AXI_FIXED_IGNORE_MIN_VALUE:`SVT_AXI_FIXED_IGNORE_MAX_VALUE]};                                             
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF 
  /**
  *  Covergroup     : trans_cross_ace_awsnoop_awsize
  *
  * Coverpoints:
  *
  * - coherent_write_xact_type:  Captures coherent write transaction
  * - burst_size: Captures transaction burst sizes
  * .
  * Cross coverpoints:
  * - awsnoop_awsize : Crosses cover points
  *    coherent_write_xact_type and burst_size
  * .
  */

`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_awsnoop_awsize (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {

      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_no_writeevict_dwlt_16 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_no_writeevict_dwlt_32 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_no_writeevict_dwlt_64 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_no_writeevict_dwlt_128 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_no_writeevict_dwlt_256 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_no_writeevict_dwlt_512 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_no_writeevict_dwlt_1024 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_no_writeevict_dweq_1024 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_writeevict_dwlt_16 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_writeevict_dwlt_32 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_writeevict_dwlt_64 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_writeevict_dwlt_128 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_writeevict_dwlt_256 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_writeevict_dwlt_512 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_writeevict_dwlt_1024 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_no_barrier_writeevict_dweq_1024 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_no_writeevict_dwlt_16 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_no_writeevict_dwlt_32 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_no_writeevict_dwlt_64 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_no_writeevict_dwlt_128 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_no_writeevict_dwlt_256 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_no_writeevict_dwlt_512 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_no_writeevict_dwlt_1024 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_no_writeevict_dweq_1024  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_writeevict_dwlt_16 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_writeevict_dwlt_32  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_writeevict_dwlt_64 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_writeevict_dwlt_128 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_writeevict_dwlt_256  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_writeevict_dwlt_512  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_writeevict_dwlt_1024 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_not_ace_lite_barrier_writeevict_dweq_1024 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_no_barrier_dwlt_16 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_no_barrier_dwlt_32  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_no_barrier_dwlt_64 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_no_barrier_dwlt_128 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_no_barrier_dwlt_256  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_no_barrier_dwlt_512 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_no_barrier_dwlt_1024 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_no_barrier_dweq_1024 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_barrier_dwlt_16 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_barrier_dwlt_32 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_barrier_dwlt_64  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_barrier_dwlt_128 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_barrier_dwlt_256  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_barrier_dwlt_512 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_barrier_dwlt_1024 (int num_slaves) ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awsize_ace_lite_barrier_dweq_1024  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awsize : cross coherent_write_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size_all   =    binsof(burst_size) && 
                                                 binsof(coherent_write_xact_type) intersect {
                                                 svt_axi_transaction::WRITELINEUNIQUE,svt_axi_transaction::WRITEBARRIER,
                                                 svt_axi_transaction::EVICT,svt_axi_transaction::WRITEEVICT };
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  /**
  *  Covergroup     : trans_cross_ace_awsnoop_awaddr
  *
  * Coverpoints:
  *
  * - coherent_write_xact_type:  Captures coherent write transaction
  * - addr : Captures transaction write address
  * .
  * Cross coverpoints:
  * - awsnoop_awaddr : Crosses cover points
  *    coherent_write_xact_type and addr
  * .
  */

`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_awsnoop_awaddr ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR
    awsnoop_awaddr : cross coherent_write_xact_type, addr {
      ignore_bins Ignore_invalid_addr = binsof(coherent_write_xact_type.coherent_writebarrier_xact) && binsof(addr);
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_awsnoop_awaddr_not_ace_lite_no_barrier_no_writeevict ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    awsnoop_awaddr : cross coherent_write_xact_type, addr {
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awaddr_not_ace_lite_no_barrier_writeevict ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    awsnoop_awaddr : cross coherent_write_xact_type, addr {
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awaddr_not_ace_lite_barrier_no_writeevict ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    awsnoop_awaddr : cross coherent_write_xact_type, addr {
      ignore_bins Ignore_invalid_addr = binsof(coherent_write_xact_type.coherent_writebarrier_xact) && binsof(addr);
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awaddr_not_ace_lite_barrier_writeevict ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    awsnoop_awaddr : cross coherent_write_xact_type, addr {
      ignore_bins Ignore_invalid_addr = binsof(coherent_write_xact_type.coherent_writebarrier_xact) && binsof(addr);
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awaddr_ace_lite_no_barrier ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    awsnoop_awaddr : cross coherent_write_xact_type, addr {
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awaddr_ace_lite_barrier ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    awsnoop_awaddr : cross coherent_write_xact_type, addr {
      ignore_bins Ignore_invalid_addr = binsof(coherent_write_xact_type.coherent_writebarrier_xact) && binsof(addr);
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

 /**
  *  Covergroup     : trans_cross_ace_awsnoop_awcache
  *
  * Coverpoints:
  *
  * - coherent_write_xact_type:  Captures coherent write transaction
  * - cache_type : Captures cache type
  * .
  * Cross coverpoints:
  * - awsnoop_awcache : Crosses cover points
  *    coherent_write_xact_type and cache_type
  * .
  */

`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_awsnoop_awcache (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awcache : cross coherent_write_xact_type, cache_type, slave_port_id {

      ignore_bins Ignore_invalid_cache_barrier = binsof(coherent_write_xact_type.coherent_writebarrier_xact) && 
                                                 !binsof(cache_type) intersect {4'b0010};

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});
      ignore_bins Ig_device_nonshare_cache = binsof(coherent_write_xact_type.coherent_writenosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_awsnoop_awcache_not_ace_lite_no_barrier_no_writeevict (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awcache : cross coherent_write_xact_type, cache_type , slave_port_id{

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});
      ignore_bins Ig_device_nonshare_cache = binsof(coherent_write_xact_type.coherent_writenosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awcache_not_ace_lite_no_barrier_writeevict (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awcache : cross coherent_write_xact_type, cache_type , slave_port_id{

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});
      ignore_bins Ig_device_nonshare_cache = binsof(coherent_write_xact_type.coherent_writenosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awcache_not_ace_lite_barrier_no_writeevict (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awcache : cross coherent_write_xact_type, cache_type , slave_port_id{

      ignore_bins Ignore_invalid_cache_barrier = binsof(coherent_write_xact_type.coherent_writebarrier_xact) && 
                                                 !binsof(cache_type) intersect {4'b0010};

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});
      ignore_bins Ig_device_nonshare_cache = binsof(coherent_write_xact_type.coherent_writenosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awcache_not_ace_lite_barrier_writeevict (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awcache : cross coherent_write_xact_type, cache_type , slave_port_id{

      ignore_bins Ignore_invalid_cache_barrier = binsof(coherent_write_xact_type.coherent_writebarrier_xact) && 
                                                 !binsof(cache_type) intersect {4'b0010};

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});
      ignore_bins Ig_device_nonshare_cache = binsof(coherent_write_xact_type.coherent_writenosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awcache_ace_lite_no_barrier (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awcache : cross coherent_write_xact_type, cache_type , slave_port_id{

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});
      ignore_bins Ig_device_nonshare_cache = binsof(coherent_write_xact_type.coherent_writenosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awcache_ace_lite_barrier (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    awsnoop_awcache : cross coherent_write_xact_type, cache_type , slave_port_id{
    
      ignore_bins Ignore_invalid_cache_barrier = binsof(coherent_write_xact_type.coherent_writebarrier_xact) && 
                                                 !binsof(cache_type) intersect {4'b0010};

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});
      ignore_bins Ig_device_nonshare_cache = binsof(coherent_write_xact_type.coherent_writenosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

 /**
  * Covergroup     : trans_cross_ace_awsnoop_bresp
  *
  * Coverpoints:
  *
  * - coherent_write_xact_type:  Captures coherent write transaction
  * - bresp : Captures write response
  * .
  * Cross coverpoints:
  * - awsnoop_bresp : Crosses cover points
  *    coherent_write_xact_type and bresp
  * .
  */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_awsnoop_bresp (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_bresp : cross coherent_write_xact_type, bresp, slave_port_id {
      ignore_bins Ignore_invalid_bresp = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                          binsof(bresp.exokay_resp);

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  covergroup trans_cross_ace_awsnoop_not_ace_lite_no_barrier_no_writeevict_bresp_no_exclusive (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_NO_EXCLUSIVE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_bresp : cross coherent_write_xact_type, bresp, slave_port_id {

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_no_barrier_no_writeevict_bresp_all(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_ALL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_bresp : cross coherent_write_xact_type, bresp, slave_port_id {
      ignore_bins Ignore_invalid_bresp = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                          binsof(bresp.exokay_resp);

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_no_barrier_writeevict_bresp_no_exclusive(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_NO_EXCLUSIVE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_bresp : cross coherent_write_xact_type, bresp, slave_port_id {

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_no_barrier_writeevict_bresp_all(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_ALL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_bresp : cross coherent_write_xact_type, bresp, slave_port_id {
      ignore_bins Ignore_invalid_bresp = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                          binsof(bresp.exokay_resp);

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_barrier_no_writeevict_bresp_no_exclusive(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_NO_EXCLUSIVE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_bresp : cross coherent_write_xact_type, bresp, slave_port_id {

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_barrier_no_writeevict_bresp_all(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_ALL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_bresp : cross coherent_write_xact_type, bresp, slave_port_id {
      ignore_bins Ignore_invalid_bresp = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                          binsof(bresp.exokay_resp);

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_barrier_writeevict_bresp_no_exclusive(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_NO_EXCLUSIVE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_bresp : cross coherent_write_xact_type, bresp, slave_port_id {

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_barrier_writeevict_bresp_all(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_ALL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_bresp : cross coherent_write_xact_type, bresp, slave_port_id {
      ignore_bins Ignore_invalid_bresp = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                          binsof(bresp.exokay_resp);

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_ace_lite_no_barrier_bresp_no_exclusive(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_NO_EXCLUSIVE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_bresp : cross coherent_write_xact_type, bresp, slave_port_id {

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_ace_lite_no_barrier_bresp_all(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_ALL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_bresp : cross coherent_write_xact_type, bresp, slave_port_id {
      ignore_bins Ignore_invalid_bresp = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                          binsof(bresp.exokay_resp);

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_ace_lite_barrier_bresp_no_exclusive(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_NO_EXCLUSIVE_AXI4_LITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_bresp : cross coherent_write_xact_type, bresp, slave_port_id {

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_ace_lite_barrier_bresp_all(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP_ALL
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_bresp : cross coherent_write_xact_type, bresp, slave_port_id {
      ignore_bins Ignore_invalid_bresp = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                          binsof(bresp.exokay_resp);

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

 /**
  *  Covergroup     : trans_cross_ace_awsnoop_awdomain
  *
  * Coverpoints:
  *
  * - coherent_write_xact_type:  Captures coherent write transaction
  * - domain_type : Captures domain type
  * .
  * Cross coverpoints:
  * - awsnoop_awdomain : Crosses cover points
  *    coherent_write_xact_type and domain_type
  * .
  */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  covergroup trans_cross_ace_awsnoop_awdomain (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    
    awsnoop_awdomain : cross coherent_write_xact_type, domain_type, slave_port_id {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_awsnoop_not_ace_lite_no_barrier_no_writeevict_awdomain (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awdomain : cross coherent_write_xact_type, domain_type , slave_port_id{

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_no_barrier_writeevict_awdomain(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awdomain : cross coherent_write_xact_type, domain_type , slave_port_id{

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_barrier_no_writeevict_awdomain(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awdomain : cross coherent_write_xact_type, domain_type , slave_port_id{

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_barrier_writeevict_awdomain(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awdomain : cross coherent_write_xact_type, domain_type , slave_port_id{

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_ace_lite_no_barrier_awdomain(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awdomain : cross coherent_write_xact_type, domain_type , slave_port_id{

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_ace_lite_barrier_awdomain(int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    awsnoop_awdomain : cross coherent_write_xact_type, domain_type , slave_port_id{

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

/**
  *  Covergroup     : trans_cross_ace_awsnoop_awdomain_awcache
  *
  * Coverpoints:
  *
  * - coherent_write_xact_type:  Captures coherent write transaction
  * - domain_type : Captures domain type
  * - cache_type  : Captures cache type 
  * .
  * Cross coverpoints:
  * - awsnoop_awdomain_awcache : Crosses cover points
  *    coherent_write_xact_type and domain_type and cache_type
  * .
  */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  covergroup trans_cross_ace_awsnoop_awdomain_awcache ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4
    

    awsnoop_awdomain_awcache : cross coherent_write_xact_type, domain_type, cache_type {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
                                            
      ignore_bins Ignore_invalid_cache_barrier = binsof(coherent_write_xact_type.coherent_writebarrier_xact) && 
                                                 !binsof(cache_type) intersect {4'b0010};

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});
      
      ignore_bins Ig_device_nonshare_cache = binsof(coherent_write_xact_type.coherent_writenosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001}); 
      
      ignore_bins Ig_device_non_system_shareable = (binsof(cache_type) intersect {4'b0000,4'b0001}) &&
                                                   (!binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE}); 

      ignore_bins Ig_cacheable_system_shareable = (binsof(cache_type) intersect {4'b0110,4'b0111,
                                                                                 4'b1010,4'b1011,4'b1110,4'b1111}) &&
                                                  (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      
      
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_awsnoop_awdomain_awcache_not_ace_lite_no_barrier_no_writeevict ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4

    awsnoop_awdomain_awcache : cross coherent_write_xact_type, domain_type, cache_type {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_write_xact_type.coherent_writenosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001}); 

      ignore_bins Ig_device_non_system_shareable = (binsof(cache_type) intersect {4'b0000,4'b0001}) &&
                                                   (!binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE}); 

      ignore_bins Ig_cacheable_system_shareable = (binsof(cache_type) intersect {4'b0110,4'b0111,
                                                                                 4'b1010,4'b1011,4'b1110,4'b1111}) &&
                                                  (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      
      
      
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awdomain_awcache_not_ace_lite_no_barrier_writeevict;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4
    awsnoop_awdomain_awcache : cross coherent_write_xact_type, domain_type, cache_type {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_write_xact_type.coherent_writenosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});  

      ignore_bins Ig_device_non_system_shareable = (binsof(cache_type) intersect {4'b0000,4'b0001}) &&
                                                   (!binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE}); 

      ignore_bins Ig_cacheable_system_shareable = (binsof(cache_type) intersect {4'b0110,4'b0111,
                                                                                 4'b1010,4'b1011,4'b1110,4'b1111}) &&
                                                  (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      
      
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awdomain_awcache_not_ace_lite_barrier_no_writeevict;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4

    awsnoop_awdomain_awcache : cross coherent_write_xact_type, domain_type, cache_type {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_invalid_cache_barrier = binsof(coherent_write_xact_type.coherent_writebarrier_xact) && 
                                                 !binsof(cache_type) intersect {4'b0010};

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_write_xact_type.coherent_writenosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});  

      ignore_bins Ig_device_non_system_shareable = (binsof(cache_type) intersect {4'b0000,4'b0001}) &&
                                                   (!binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE}); 

      ignore_bins Ig_cacheable_system_shareable = (binsof(cache_type) intersect {4'b0110,4'b0111,
                                                                                 4'b1010,4'b1011,4'b1110,4'b1111}) &&
                                                  (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      
      
      
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awdomain_awcache_not_ace_lite_barrier_writeevict;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4

    awsnoop_awdomain_awcache : cross coherent_write_xact_type, domain_type, cache_type {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_invalid_cache_barrier = binsof(coherent_write_xact_type.coherent_writebarrier_xact) && 
                                                 !binsof(cache_type) intersect {4'b0010};

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_write_xact_type.coherent_writenosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001}); 

      ignore_bins Ig_device_non_system_shareable = (binsof(cache_type) intersect {4'b0000,4'b0001}) &&
                                                   (!binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE}); 

      ignore_bins Ig_cacheable_system_shareable = (binsof(cache_type) intersect {4'b0110,4'b0111,
                                                                                 4'b1010,4'b1011,4'b1110,4'b1111}) &&
                                                  (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      
      
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awdomain_awcache_ace_lite_no_barrier;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4
    
    awsnoop_awdomain_awcache : cross coherent_write_xact_type, domain_type, cache_type {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_write_xact_type.coherent_writenosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});

      ignore_bins Ig_device_non_system_shareable = (binsof(cache_type) intersect {4'b0000,4'b0001}) &&
                                                   (!binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE}); 

      ignore_bins Ig_cacheable_system_shareable = (binsof(cache_type) intersect {4'b0110,4'b0111,
                                                                                 4'b1010,4'b1011,4'b1110,4'b1111}) &&
                                                  (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      
      
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_awdomain_awcache_ace_lite_barrier;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_AWCACHE_TYPE_AXI4

    awsnoop_awdomain_awcache : cross coherent_write_xact_type, domain_type, cache_type {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_invalid_cache_barrier = binsof(coherent_write_xact_type.coherent_writebarrier_xact) && 
                                                 !binsof(cache_type) intersect {4'b0010};

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_write_xact_type.coherent_writenosnoop_xact)) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});
      ignore_bins Ig_device_nonshare_cache = binsof(coherent_write_xact_type.coherent_writenosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});  

      ignore_bins Ig_device_non_system_shareable = (binsof(cache_type) intersect {4'b0000,4'b0001}) &&
                                                   (!binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE}); 

      ignore_bins Ig_cacheable_system_shareable = (binsof(cache_type) intersect {4'b0110,4'b0111,
                                                                                 4'b1010,4'b1011,4'b1110,4'b1111}) &&
                                                  (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF


 /**
  * Covergroup     : trans_cross_ace_awsnoop_awbar
  *
  * Coverpoints:
  *
  * - coherent_write_xact_type:  Captures coherent write transaction
  * - barrier_type : Captures write barrier
  * .
  * Cross coverpoints:
  * - awsnoop_awbar : Crosses cover points
  *    coherent_write_xact_type and barrier_type
  * .
  */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF 
  covergroup trans_cross_ace_awsnoop_awbar ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_TYPE

    awsnoop_awbar : cross coherent_write_xact_type, barrier_type {

      ignore_bins Ignore_normal = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});

      ignore_bins Ignore_barrier = (!binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                   (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  covergroup trans_cross_ace_awsnoop_not_ace_lite_no_barrier_no_writeevict_awbar_unset ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_UNSET

    awsnoop_awbar : cross coherent_write_xact_type, barrier_type {

      ignore_bins Ignore_normal = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_no_barrier_writeevict_awbar_unset ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_UNSET

    awsnoop_awbar : cross coherent_write_xact_type, barrier_type {

      ignore_bins Ignore_normal = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_ace_awsnoop_not_ace_lite_barrier_no_writeevict_awbar_set;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_SET

    awsnoop_awbar : cross coherent_write_xact_type, barrier_type {

      ignore_bins Ignore_normal = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});

      ignore_bins Ignore_barrier = (!binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                   (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_ace_awsnoop_not_ace_lite_barrier_writeevict_awbar_set;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_SET

    awsnoop_awbar : cross coherent_write_xact_type, barrier_type {

      ignore_bins Ignore_normal = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});

      ignore_bins Ignore_barrier = (!binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                   (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_ace_awsnoop_ace_lite_no_barrier_awbar_unset;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_UNSET

    awsnoop_awbar : cross coherent_write_xact_type, barrier_type {

      ignore_bins Ignore_normal = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  
  covergroup trans_cross_ace_awsnoop_ace_lite_barrier_awbar_set;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_SET

    awsnoop_awbar : cross coherent_write_xact_type, barrier_type {

      ignore_bins Ignore_normal = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});

      ignore_bins Ignore_barrier = (!binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                   (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  // Added in 2.43a
//`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF  

  /**
  * Covergroup     : trans_cross_ace_awdomain_awbarrier_memory_sync
  *
  * Coverpoints:
  *
  * - coherent_write_xact_type:  Captures coherent write transaction
  * - barrier_type : Captures write barrier
  * - domain_type : Captures domain type
  * .
  * Cross coverpoints:
  * - awbarrier_awdomain : Crosses cover points
  *   write transaction of certain barrier_type MEMORY_BARRIER & SYNC_BARRIER with awdomain
  * .
  * As barrier types are memory & sync therefore, ignoring bins intersect with NORMAL_ACCESS_RESPECT_BARRIER & NORMAL_ACCESS_IGNORE_BARRIER
  * and ignoring all other non-writebarrier bins.
  */

  covergroup trans_cross_ace_awdomain_awbarrier_memory_sync ;
    //`SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    coherent_write_xact_type : coverpoint cov_item.coherent_xact_type iff(cov_coherent_xact_type_flag){
      bins coherent_writebarrier_xact = {svt_axi_transaction::WRITEBARRIER};
      option.weight = 0;
    }
    // Only MEMORY_BARRIER and SYNC_BARRIER are being covered, so we need to use only the BARRIER_SET macro
    //`SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_TYPE 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE

    awdomain_awbarrier_memory_sync : cross coherent_write_xact_type, barrier_type, domain_type {

      ignore_bins ignore_normal = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});

      ignore_bins ignore_non_write_barrier = (!binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /**
  * Covergroup     : trans_cross_ace_awdomain_awbarrier_respect_ignore
  *
  * Coverpoints:
  *
  * - coherent_write_xact_type:  Captures coherent write transaction
  * - barrier_type : Captures non write barrier (all other coherent transactions) as its normal access with respect or ignore barrier
  * - domain_type : Captures domain type
  * .
  * Cross coverpoints:
  * - awbarrier_awdomain : Crosses cover points
  *   write transaction of certain barrier_type NORMAL_ACCESS_RESPECT_BARRIER and NORMAL_ACCESS_IGNORE_BARRIER with awdomain
  * .
  * As barrier type with respect & ignore barriers are normal coherent access therefore, ignoring bins are WRITEBARRIER with Memory & Sync
  */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_awdomain_awbarrier_respect_ignore ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE

    awdomain_awbarrier_respect_ignore  : cross coherent_write_xact_type, barrier_type, domain_type {

      ignore_bins  ignore_memory_sync_barrier = (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});
      ignore_bins ignore_write_barrier = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER});
      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
   
`else
  covergroup trans_cross_ace_awdomain_awbarrier_respect_ignore_not_ace_lite_no_writeevict ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE

    awdomain_awbarrier_respect_ignore  : cross coherent_write_xact_type, barrier_type, domain_type {

      ignore_bins  ignore_memory_sync_barrier = (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});
      ignore_bins ignore_write_barrier = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER});
      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awdomain_awbarrier_respect_ignore_not_ace_lite_writeevict ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE

    awdomain_awbarrier_respect_ignore  : cross coherent_write_xact_type, barrier_type, domain_type {

      ignore_bins  ignore_memory_sync_barrier = (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});
      ignore_bins ignore_write_barrier = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER});
      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                           {svt_axi_transaction::WRITECLEAN,svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITEEVICT}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awdomain_awbarrier_respect_ignore_ace_lite;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_ACE_LITE_NO_BARRIER
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE

    awdomain_awbarrier_respect_ignore  : cross coherent_write_xact_type, barrier_type, domain_type {

      ignore_bins  ignore_memory_sync_barrier = (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});
      ignore_bins ignore_write_barrier = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER});
      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITENOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_write_xact_type) intersect 
                                                   {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE,
                                                    svt_axi_transaction::EVICT}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
   
`endif

/**
  * Covergroup     : trans_cross_ace_ardomain_arbarrier_memory_sync
  *
  * Coverpoints:
  *
  * - coherent_read_xact_type:  Captures coherent read transaction
  * - barrier_type : Captures read barrier
  * - domain_type : Captures domain type
  * .
  * Cross coverpoints:
  * - arbarrier_ardomain : Crosses cover points
  *   read transaction of certain barrier_type MEMORY_BARRIER & SYNC_BARRIER with ardomain
  * As barrier types are memory & sync therefore, ignoring bins intersect with NORMAL_ACCESS_RESPECT_BARRIER & NORMAL_ACCESS_IGNORE_BARRIER
  * and ignoring all other non-readbarrier bins.
  * .
  */

  covergroup trans_cross_ace_ardomain_arbarrier_memory_sync ;
    //`SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    coherent_read_xact_type : coverpoint cov_item.coherent_xact_type iff(cov_coherent_xact_type_flag){
      bins coherent_readbarrier_xact = {svt_axi_transaction::READBARRIER};
      option.weight = 0;
    }
    // Only MEMORY_BARRIER and SYNC_BARRIER are being covered, so we need to use only the BARRIER_SET macro
    //`SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_TYPE 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE

    ardomain_arbarrier_memory_sync : cross coherent_read_xact_type, barrier_type, domain_type {

      ignore_bins ignore_normal = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});

      ignore_bins ignore_non_read_barrier = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /**
  * Covergroup     : trans_cross_ace_ardomain_arbarrier_respect_ignore
  *
  * Coverpoints:
  *
  * - coherent_read_xact_type:  Captures coherent read transaction
  * - barrier_type : Captures non read barrier (all other coherent transactions) as its normal access with respect or ignore barrier
  * - domain_type : Captures domain type
  * .
  * Cross coverpoints:
  * - arbarrier_ardomain : Crosses cover points
  *   read transaction of certain barrier_type NORMAL_ACCESS_RESPECT_BARRIER and NORMAL_ACCESS_IGNORE_BARRIER with ardomain
  * .
  * As barrier type with respect & ignore barriers are normal coherent access therefore, ignoring bins are READBARRIER with Memory & Sync
  */

`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF 
  covergroup trans_cross_ace_ardomain_arbarrier_respect_ignore ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE

    ardomain_arbarrier_respect_ignore  : cross coherent_read_xact_type, barrier_type, domain_type {

      ignore_bins  ignore_memory_sync_barrier = (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});

      ignore_bins ignore_read_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER});
      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});
`ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else 
       ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  `else
  covergroup trans_cross_ace_ardomain_arbarrier_respect_ignore_dvm_set;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    ardomain_arbarrier_respect_ignore  : cross coherent_read_xact_type, barrier_type, domain_type {

      ignore_bins  ignore_memory_sync_barrier = (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});

      ignore_bins ignore_read_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER});
      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                               svt_axi_transaction::SYSTEMSHAREABLE});

`ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else 
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif

      option.weight = 1;
    }
    option.per_instance = 1;

  endgroup

  covergroup trans_cross_ace_ardomain_arbarrier_respect_ignore_dvm_unset;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    ardomain_arbarrier_respect_ignore  : cross coherent_read_xact_type, barrier_type, domain_type {

      ignore_bins  ignore_memory_sync_barrier = (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});

      ignore_bins ignore_read_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER});
      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});
 `ifdef SVT_ACE5_ENABLE 
    ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
 `else
    ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
 `endif 

      option.weight = 1;
    }
    option.per_instance = 1;

  endgroup

  covergroup trans_cross_ace_ardomain_arbarrier_respect_ignore_ace_lite_dvm_set;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    ardomain_arbarrier_respect_ignore  : cross coherent_read_xact_type, barrier_type, domain_type {

      ignore_bins  ignore_memory_sync_barrier = (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});

      ignore_bins ignore_read_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER});
      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE, svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});
 `ifdef SVT_ACE5_ENABLE 
    ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
 `else
    ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
 `endif 
      option.weight = 1;
    }
    option.per_instance = 1;

  endgroup

  covergroup trans_cross_ace_ardomain_arbarrier_respect_ignore_ace_lite_dvm_unset;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    ardomain_arbarrier_respect_ignore  : cross coherent_read_xact_type, barrier_type, domain_type {

      ignore_bins  ignore_memory_sync_barrier = (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});

      ignore_bins ignore_read_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER});
      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});
 `ifdef SVT_ACE5_ENABLE 
    ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
 `else
    ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
 `endif 

        option.weight = 1;
    }
    option.per_instance = 1;

  endgroup

  `endif

    
  /**
  * Covergroup     : trans_cross_ace_awsnoop_awdomain_bresp
  *
  * Coverpoints:
  *
  * - coherent_write_xact_type:  Captures coherent writenosnoop transaction
  * - bresp : Captures exokay write response
  * - domain_type : Captures NONSHAREABLE & SYSTEMSHAREABLE domain types
  * .
  * Cross coverpoints:
  * - awsnoop_awdomain_bresp : Crosses cover points
  *    coherent_write_xact_type, domain_type and bresp
  * .
  * The EXOKAY response is permitted for WriteNoSnoop with domain innershareable & outershareable. Rest all other bins are ignored.
  */

  covergroup trans_cross_ace_awsnoop_awdomain_bresp ;
    // Only WRITENOSNOOP is covered by this group. So cover only that
    //`SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    coherent_write_xact_type : coverpoint cov_item.coherent_xact_type iff(cov_coherent_xact_type_flag){ 
      bins coherent_writenosnoop_xact   = {svt_axi_transaction::WRITENOSNOOP}; 
    }
    // Only EXOKAY response is being covered by this; so create covergroup only for that
    //`SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP
    bresp : coverpoint cov_item.bresp iff(cov_bresp_flag){ 
      bins exokay_resp  = {svt_axi_transaction::EXOKAY}; 
    }
    domain_type : coverpoint cov_item.domain_type iff(cov_domain_type_flag){ 
      bins domain_non_shareable           = {svt_axi_transaction::NONSHAREABLE}; 
      bins domain_system_shareable        = {svt_axi_transaction::SYSTEMSHAREABLE}; 
      option.weight = 1; 
    }

    awsnoop_awdomain_bresp : cross coherent_write_xact_type, bresp, domain_type {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
//`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  /**
  *  Covergroup     : trans_cross_ace_arsnoop_arburst
  *
  * Coverpoints:
  *
  * - coherent_read_xact_type:  Captures coherent read transaction
  * - burst_type: Captures transaction burst type
  * .
  * Cross coverpoints:
  * - arsnoop_arburst : Crosses cover points
  *    coherent_read_xact_type and burst_type
  * .
  */

  //covergroup trans_cross_ace_arsnoop_arburst @(cov_read_sample_event);
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF  
  covergroup trans_cross_ace_arsnoop_arburst (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_arburst : cross coherent_read_xact_type, burst_type, slave_port_id {

      ignore_bins Ignore_invalid_fixed   =  binsof(burst_type.fixed_burst) &&
                                                (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP});

`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) &&
                                                (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                            svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE});
 `endif
      // DVM, BARRIER :: alen == 0x00
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::DVMCOMPLETE, 
                                                                                        svt_axi_transaction::DVMMESSAGE, 
                                                                                        svt_axi_transaction::READBARRIER};

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else
  covergroup trans_cross_ace_arsnoop_arburst_def (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

             arsnoop_arburst : cross coherent_read_xact_type, burst_type , slave_port_id{

      ignore_bins Ignore_invalid_fixed   =  binsof(burst_type.fixed_burst) &&
                                                (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP});

`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) &&
                                                (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                            svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE});
 `endif
      // DVM, BARRIER :: alen == 0x00
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::DVMCOMPLETE, 
                                                                                        svt_axi_transaction::DVMMESSAGE, 
                                                                                        svt_axi_transaction::READBARRIER};

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arburst_dvm_unset_barrier_set (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

            arsnoop_arburst : cross coherent_read_xact_type, burst_type , slave_port_id{

      ignore_bins Ignore_invalid_fixed   =  binsof(burst_type.fixed_burst) &&
                                                (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP});

`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) &&
                                                (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                            svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE});
 `endif
      // DVM, BARRIER :: alen == 0x00
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::DVMCOMPLETE, 
                                                                                        svt_axi_transaction::DVMMESSAGE, 
                                                                                        svt_axi_transaction::READBARRIER};

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arburst_dvm_set_barrier_unset (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_arburst : cross coherent_read_xact_type, burst_type , slave_port_id{

      ignore_bins Ignore_invalid_fixed   =  binsof(burst_type.fixed_burst) &&
                                                (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP});

`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) &&
                                                (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                            svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE});
 `endif
      // DVM, BARRIER :: alen == 0x00
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::DVMCOMPLETE, 
                                                                                        svt_axi_transaction::DVMMESSAGE, 
                                                                                        svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arburst_dvm_set_barrier_set (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_arburst : cross coherent_read_xact_type, burst_type , slave_port_id{

      ignore_bins Ignore_invalid_fixed   =  binsof(burst_type.fixed_burst) &&
                                                (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP});

`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) &&
                                                (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                            svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE});
 `endif
      // DVM, BARRIER :: alen == 0x00
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::DVMCOMPLETE, 
                                                                                        svt_axi_transaction::DVMMESSAGE, 
                                                                                        svt_axi_transaction::READBARRIER};

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arburst_ace_lite_barrier_set (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_arburst : cross coherent_read_xact_type, burst_type , slave_port_id{

      ignore_bins Ignore_invalid_fixed   =  binsof(burst_type.fixed_burst) &&
                                                (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP});

`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) &&
                                                (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                            svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE});
 `endif
      // DVM, BARRIER :: alen == 0x00
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::DVMCOMPLETE, 
                                                                                        svt_axi_transaction::DVMMESSAGE, 
                                                                                        svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup 

  covergroup trans_cross_ace_arsnoop_arburst_ace_lite_barrier_unset (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE_AXI3_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arburst : cross coherent_read_xact_type, burst_type , slave_port_id{

      ignore_bins Ignore_invalid_fixed   =  binsof(burst_type.fixed_burst) &&
                                                (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP});

`ifndef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
      ignore_bins Ignore_invalid_wrap   =  binsof(burst_type.wrap_burst) &&
                                                (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                            svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE});
 `endif
      // DVM, BARRIER :: alen == 0x00
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::DVMCOMPLETE, 
                                                                                        svt_axi_transaction::DVMMESSAGE, 
                                                                                        svt_axi_transaction::READBARRIER};

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif
  /**
  *  Covergroup     : trans_cross_ace_arsnoop_arlen
  *
  * Coverpoints:
  *
  * - coherent_read_xact_type:  Captures coherent read transaction
  * - burst_length: Captures transaction burst length
  * .
  * Cross coverpoints:
  * - arsnoop_arlen : Crosses cover points
  *    coherent_read_xact_type and burst_length
  * .
  */

  //covergroup trans_cross_ace_arsnoop_arlen @(cov_read_sample_event);

`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_arsnoop_arlen (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_arlen : cross coherent_read_xact_type, burst_length, slave_port_id {

      ignore_bins Ignore_invalid_length   = binsof(burst_length) &&
                                                   (!binsof(coherent_read_xact_type) 
                                                     intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
`ifdef SVT_ACE5_ENABLE 
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ig_len_for_CLsize_coh_txn when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`else
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7],[9:15]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`endif
`else 
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ig_len_for_CLsize_coh_txn when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`else
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7],[9:15]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`endif
`endif

      ignore_bins Ig_len_for_evict_dvm_barrier = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::EVICT, 
                                                   svt_axi_transaction::DVMCOMPLETE, svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else
  covergroup trans_cross_ace_arsnoop_arlen_def  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arlen : cross coherent_read_xact_type, burst_length , slave_port_id{

      ignore_bins Ignore_invalid_length   = binsof(burst_length) &&
                                                   (!binsof(coherent_read_xact_type) 
                                                     intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
`ifdef SVT_ACE5_ENABLE 
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ig_len_for_CLsize_coh_txn when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`else
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7],[9:15]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`endif
`else 
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ig_len_for_CLsize_coh_txn when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`else
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7],[9:15]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`endif
`endif
      ignore_bins Ig_len_for_evict_dvm_barrier = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::EVICT, 
                                                   svt_axi_transaction::DVMCOMPLETE, svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arlen_dvm_unset_barrier_set (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arlen : cross coherent_read_xact_type, burst_length , slave_port_id{

      ignore_bins Ignore_invalid_length   = binsof(burst_length) &&
                                                   (!binsof(coherent_read_xact_type) 
                                                     intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
`ifdef SVT_ACE5_ENABLE 
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ig_len_for_CLsize_coh_txn when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`else
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7],[9:15]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`endif
`else 
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ig_len_for_CLsize_coh_txn when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`else
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7],[9:15]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`endif
`endif
      ignore_bins Ig_len_for_evict_dvm_barrier = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::EVICT, 
                                                   svt_axi_transaction::DVMCOMPLETE, svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arlen_dvm_set_barrier_unset (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arlen : cross coherent_read_xact_type, burst_length , slave_port_id{

      ignore_bins Ignore_invalid_length   = binsof(burst_length) &&
                                                   (!binsof(coherent_read_xact_type) 
                                                     intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
`ifdef SVT_ACE5_ENABLE 
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ig_len_for_CLsize_coh_txn when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`else
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7],[9:15]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`endif
`else 
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ig_len_for_CLsize_coh_txn when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`else
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7],[9:15]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`endif
`endif
      ignore_bins Ig_len_for_evict_dvm_barrier = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::EVICT, 
                                                   svt_axi_transaction::DVMCOMPLETE, svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arlen_dvm_set_barrier_set (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arlen : cross coherent_read_xact_type, burst_length , slave_port_id{

      ignore_bins Ignore_invalid_length   = binsof(burst_length) &&
                                                   (!binsof(coherent_read_xact_type) 
                                                     intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
`ifdef SVT_ACE5_ENABLE 
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ig_len_for_CLsize_coh_txn when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`else
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7],[9:15]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`endif
`else 
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ig_len_for_CLsize_coh_txn when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`else
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7],[9:15]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`endif
`endif
      ignore_bins Ig_len_for_evict_dvm_barrier = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::EVICT, 
                                                   svt_axi_transaction::DVMCOMPLETE, svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arlen_ace_lite_barrier_unset (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arlen : cross coherent_read_xact_type, burst_length , slave_port_id{

      ignore_bins Ignore_invalid_length   = binsof(burst_length) &&
                                                   (!binsof(coherent_read_xact_type) 
                                                     intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
`ifdef SVT_ACE5_ENABLE 
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ig_len_for_CLsize_coh_txn when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`else
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7],[9:15]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`endif
`else 
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ig_len_for_CLsize_coh_txn when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`else
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7],[9:15]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`endif
`endif
      ignore_bins Ig_len_for_evict_dvm_barrier = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::EVICT, 
                                                   svt_axi_transaction::DVMCOMPLETE, svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arlen_ace_lite_barrier_set (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH_ACE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arlen : cross coherent_read_xact_type, burst_length , slave_port_id{

      ignore_bins Ignore_invalid_length   = binsof(burst_length) &&
                                                   (!binsof(coherent_read_xact_type) 
                                                     intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
`ifdef SVT_ACE5_ENABLE 
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ig_len_for_CLsize_coh_txn when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`else
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7],[9:15]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`endif
`else 
`ifdef SVT_AXI_MAX_BURST_LENGTH_WIDTH_1
     // no need to ignore Ig_len_for_CLsize_coh_txn when burst length width is 1
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_2
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`elsif SVT_AXI_MAX_BURST_LENGTH_WIDTH_3
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`else
      ignore_bins Ig_len_for_CLsize_coh_txn = (binsof(burst_length) intersect {[2:3],[5:7],[9:15]}) &&
                                              (binsof(coherent_read_xact_type) intersect 
                                                 {svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                  svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE,
                                                  svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANUNIQUE,
                                                  svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID,
                                                  svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}
                                              );
`endif
`endif
      ignore_bins Ig_len_for_evict_dvm_barrier = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::EVICT, 
                                                   svt_axi_transaction::DVMCOMPLETE, svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup


`endif
  /**
  *  Covergroup     : trans_cross_ace_arsnoop_arsize
  *
  * Coverpoints:
  *
  * - coherent_read_xact_type:  Captures coherent read transaction
  * - burst_size: Captures transaction burst size
  * .
  * Cross coverpoints:
  * - arsnoop_arsize : Crosses cover points
  *    coherent_read_xact_type and burst_size
  * .
  */

  //covergroup trans_cross_ace_arsnoop_arsize @(cov_read_sample_event);
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_arsnoop_arsize (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  covergroup trans_cross_ace_arsnoop_arsize_def_dwlt_16  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size , slave_port_id{
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_def_dwlt_32  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_def_dwlt_64  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_def_dwlt_128  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_def_dwlt_256  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_def_dwlt_512  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_def_dwlt_1024  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_def_dweq_1024  (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_unset_barrier_set_dwlt_16 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_unset_barrier_set_dwlt_32 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_unset_barrier_set_dwlt_64 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_unset_barrier_set_dwlt_128 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_unset_barrier_set_dwlt_256 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_unset_barrier_set_dwlt_512 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_unset_barrier_set_dwlt_1024 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_unset_barrier_set_dweq_1024 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_unset_dwlt_16 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_unset_dwlt_32 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_unset_dwlt_64 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_unset_dwlt_128 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_unset_dwlt_256 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_unset_dwlt_512 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_unset_dwlt_1024 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_unset_dweq_1024 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_set_dwlt_16 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_set_dwlt_32 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_set_dwlt_64 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_set_dwlt_128 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_set_dwlt_256 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_set_dwlt_512 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_set_dwlt_1024 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_dvm_set_barrier_set_dweq_1024 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_set_dwlt_16 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_set_dwlt_32 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_set_dwlt_64 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_set_dwlt_128 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_set_dwlt_256 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_set_dwlt_512 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_set_dwlt_1024 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_set_dweq_1024 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_unset_dwlt_16 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_16BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_unset_dwlt_32 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_32BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_unset_dwlt_64 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_64BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_unset_dwlt_128 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_128BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_unset_dwlt_256 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_256BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_unset_dwlt_512 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_512BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_unset_dwlt_1024 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_LT_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arsize_ace_lite_barrier_unset_dweq_1024 (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_SIZE_EQ_1024BIT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID
    arsnoop_arsize : cross coherent_read_xact_type, burst_size, slave_port_id {
          
      ignore_bins Ignore_invalid_size   = binsof(burst_size) &&
                                          (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE});
      ignore_bins Ig_burst_for_dvm_barrier = binsof(coherent_read_xact_type) intersect { svt_axi_transaction::DVMCOMPLETE, 
                                                        svt_axi_transaction::DVMMESSAGE, svt_axi_transaction::READBARRIER};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  /**
  *  Covergroup     : trans_cross_ace_arsnoop_araddr
  *
  * Coverpoints:
  *
  * - coherent_read_xact_type:  Captures coherent read transaction
  * - addr : Captures transaction read address
  * .
  * Cross coverpoints:
  * - arsnoop_araddr : Crosses cover points
  *    coherent_read_xact_type and addr
  * .
  */

  //covergroup trans_cross_ace_arsnoop_araddr @(cov_read_sample_event);
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_arsnoop_araddr ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR
    arsnoop_araddr : cross coherent_read_xact_type, addr {
      ignore_bins Ignore_invalid_addr = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                         svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else

  covergroup trans_cross_ace_arsnoop_araddr_def ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    arsnoop_araddr : cross coherent_read_xact_type, addr {
      ignore_bins Ignore_invalid_addr = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                         svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_araddr_dvm_unset_barrier_set ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    arsnoop_araddr : cross coherent_read_xact_type, addr {
      ignore_bins Ignore_invalid_addr = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                         svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_araddr_dvm_set_barrier_unset ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    arsnoop_araddr : cross coherent_read_xact_type, addr {
      ignore_bins Ignore_invalid_addr = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                         svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_araddr_dvm_set_barrier_set ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    arsnoop_araddr : cross coherent_read_xact_type, addr {
      ignore_bins Ignore_invalid_addr = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                         svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_araddr_ace_lite_barrier_set ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    arsnoop_araddr : cross coherent_read_xact_type, addr {
      ignore_bins Ignore_invalid_addr = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                         svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_araddr_ace_lite_barrier_unset ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR_ACE
    arsnoop_araddr : cross coherent_read_xact_type, addr {
      ignore_bins Ignore_invalid_addr = binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                         svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE};
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif

 /**
  *  Covergroup     : trans_cross_ace_arsnoop_arcache
  *
  * Coverpoints:
  *
  * - coherent_read_xact_type:  Captures coherent read transaction
  * - cache_type : Captures transaction cache type
  * .
  * Cross coverpoints:
  * - arsnoop_arcache : Crosses cover points
  *    coherent_read_xact_type and cache_type
  * .
  */

  //covergroup trans_cross_ace_arsnoop_arcache @(cov_read_sample_event);
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF  
  covergroup trans_cross_ace_arsnoop_arcache (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_arcache : cross coherent_read_xact_type, cache_type, slave_port_id {

      ignore_bins Ignore_invalid_cache_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                  svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                  (!binsof(cache_type) intersect {4'b0010});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_read_xact_type.coherent_readnosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_arsnoop_arcache_def (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_arcache : cross coherent_read_xact_type, cache_type , slave_port_id{

      ignore_bins Ignore_invalid_cache_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                  svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                  (!binsof(cache_type) intersect {4'b0010});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_read_xact_type.coherent_readnosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arcache_dvm_unset_barrier_set (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_arcache : cross coherent_read_xact_type, cache_type , slave_port_id{

      ignore_bins Ignore_invalid_cache_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                  svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                  (!binsof(cache_type) intersect {4'b0010});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_read_xact_type.coherent_readnosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arcache_dvm_set_barrier_unset (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_arcache : cross coherent_read_xact_type, cache_type , slave_port_id{

      ignore_bins Ignore_invalid_cache_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                  svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                  (!binsof(cache_type) intersect {4'b0010});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_read_xact_type.coherent_readnosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arcache_dvm_set_barrier_set (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_arcache : cross coherent_read_xact_type, cache_type , slave_port_id{

      ignore_bins Ignore_invalid_cache_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                  svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                  (!binsof(cache_type) intersect {4'b0010});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_read_xact_type.coherent_readnosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arcache_ace_lite_barrier_unset (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_arcache : cross coherent_read_xact_type, cache_type , slave_port_id{

      ignore_bins Ignore_invalid_cache_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                  svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                  (!binsof(cache_type) intersect {4'b0010});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_read_xact_type.coherent_readnosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arcache_ace_lite_barrier_set (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_arcache : cross coherent_read_xact_type, cache_type , slave_port_id{

      ignore_bins Ignore_invalid_cache_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                  svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                  (!binsof(cache_type) intersect {4'b0010});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_read_xact_type.coherent_readnosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
/**
  *  Covergroup     : trans_cross_ace_arsnoop_ardomain
  *
  * Coverpoints:
  *
  * - coherent_read_xact_type:  Captures coherent read transaction
  * - domain_type : Captures domain type
  * .
  * Cross coverpoints:
  * - arsnoop_ardomain : Crosses cover points
  *    coherent_read_xact_type and domain_type
  * .
  */

  //covergroup trans_cross_ace_arsnoop_ardomain @(cov_read_sample_event);
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF  
  covergroup trans_cross_ace_arsnoop_ardomain (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_ardomain : cross coherent_read_xact_type, domain_type, slave_port_id {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

`ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else
     ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else
  covergroup trans_cross_ace_arsnoop_ardomain_def (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_ardomain : cross coherent_read_xact_type, domain_type , slave_port_id{

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

`ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else
     ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_ardomain_dvm_unset_barrier_set (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_ardomain : cross coherent_read_xact_type, domain_type , slave_port_id{

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

`ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else
     ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_ardomain_dvm_set_barrier_unset (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_ardomain : cross coherent_read_xact_type, domain_type , slave_port_id{

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

     `ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else
     ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif
 option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_ardomain_dvm_set_barrier_set (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_ardomain : cross coherent_read_xact_type, domain_type , slave_port_id{

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

 `ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else
     ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_ardomain_ace_lite_barrier_unset (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_ardomain : cross coherent_read_xact_type, domain_type , slave_port_id{

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

  `ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else
     ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif
     option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_ardomain_ace_lite_barrier_set (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_ardomain : cross coherent_read_xact_type, domain_type , slave_port_id{

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

    `ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else
     ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif
  option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif

/**
  *  Covergroup     : trans_cross_ace_arsnoop_ardomain_arcache
  *
  * Coverpoints:
  *
  * - coherent_read_xact_type:  Captures coherent read transaction
  * - domain_type : Captures domain type
  * - cache_type : Captures cache_type
  * .
  * Cross coverpoints:
  * - arsnoop_ardomain_arcache : Crosses cover points
  *   coherent_read_xact_type and domain_type and cache_type
  * .
  */

  //covergroup trans_cross_ace_arsnoop_ardomain @(cov_read_sample_event);
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF  
  covergroup trans_cross_ace_arsnoop_ardomain_arcache ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4

    arsnoop_ardomain_arcache : cross coherent_read_xact_type, domain_type, cache_type {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_invalid_cache_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                  svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                  (!binsof(cache_type) intersect {4'b0010});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_read_xact_type.coherent_readnosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});

      ignore_bins Ig_device_non_system_shareable = (binsof(cache_type) intersect {4'b0000,4'b0001}) &&
                                                   (!binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE}); 

      ignore_bins Ig_cacheable_system_shareable = (binsof(cache_type) intersect {4'b0110,4'b0111,
                                                                                 4'b1010,4'b1011,4'b1110,4'b1111}) &&
                                                  (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      
      
`ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else
     ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`else
  covergroup trans_cross_ace_arsnoop_ardomain_arcache_def ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4
    
    arsnoop_ardomain_arcache : cross coherent_read_xact_type, domain_type, cache_type {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

 
      ignore_bins Ignore_invalid_cache_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                  svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                  (!binsof(cache_type) intersect {4'b0010});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_read_xact_type.coherent_readnosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});
      
      ignore_bins Ig_device_non_system_shareable = (binsof(cache_type) intersect {4'b0000,4'b0001}) &&
                                                   (!binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE}); 

      ignore_bins Ig_cacheable_system_shareable = (binsof(cache_type) intersect {4'b0110,4'b0111,
                                                                                 4'b1010,4'b1011,4'b1110,4'b1111}) &&
                                                  (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      
      
`ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else
     ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_ardomain_arcache_dvm_unset_barrier_set ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4

    arsnoop_ardomain_arcache : cross coherent_read_xact_type, domain_type, cache_type {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

    
      ignore_bins Ignore_invalid_cache_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                  svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                  (!binsof(cache_type) intersect {4'b0010});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_read_xact_type.coherent_readnosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});

      ignore_bins Ig_device_non_system_shareable = (binsof(cache_type) intersect {4'b0000,4'b0001}) &&
                                                   (!binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE}); 

      ignore_bins Ig_cacheable_system_shareable = (binsof(cache_type) intersect {4'b0110,4'b0111,
                                                                                 4'b1010,4'b1011,4'b1110,4'b1111}) &&
                                                  (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      

      
`ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else
     ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_ardomain_arcache_dvm_set_barrier_unset ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4

    arsnoop_ardomain_arcache : cross coherent_read_xact_type, domain_type, cache_type {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});


      ignore_bins Ignore_invalid_cache_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                  svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                  (!binsof(cache_type) intersect {4'b0010});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_read_xact_type.coherent_readnosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});

      ignore_bins Ig_device_non_system_shareable = (binsof(cache_type) intersect {4'b0000,4'b0001}) &&
                                                   (!binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE}); 

      ignore_bins Ig_cacheable_system_shareable = (binsof(cache_type) intersect {4'b0110,4'b0111,
                                                                                 4'b1010,4'b1011,4'b1110,4'b1111}) &&
                                                  (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      
      
      
`ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else
     ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_ardomain_arcache_dvm_set_barrier_set ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4

    arsnoop_ardomain_arcache : cross coherent_read_xact_type, domain_type, cache_type {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

       ignore_bins Ignore_invalid_cache_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                  svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                  (!binsof(cache_type) intersect {4'b0010});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_read_xact_type.coherent_readnosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});

      ignore_bins Ig_device_non_system_shareable = (binsof(cache_type) intersect {4'b0000,4'b0001}) &&
                                                   (!binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE}); 

      ignore_bins Ig_cacheable_system_shareable = (binsof(cache_type) intersect {4'b0110,4'b0111,
                                                                                 4'b1010,4'b1011,4'b1110,4'b1111}) &&
                                                  (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      
      
      
  `ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else
     ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif
    option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_ardomain_arcache_ace_lite_barrier_unset ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4

    arsnoop_ardomain_arcache : cross coherent_read_xact_type, domain_type, cache_type {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});

      ignore_bins Ignore_invalid_cache_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                  svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                  (!binsof(cache_type) intersect {4'b0010});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_read_xact_type.coherent_readnosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});

      ignore_bins Ig_device_non_system_shareable = (binsof(cache_type) intersect {4'b0000,4'b0001}) &&
                                                   (!binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE}); 

      ignore_bins Ig_cacheable_system_shareable = (binsof(cache_type) intersect {4'b0110,4'b0111,
                                                                                 4'b1010,4'b1011,4'b1110,4'b1111}) &&
                                                  (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      
      
      
  `ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else
     ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif
    option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_ardomain_arcache_ace_lite_barrier_set ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_ACE_LITE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_DOMAIN_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ARCACHE_TYPE_AXI4

    arsnoop_ardomain_arcache : cross coherent_read_xact_type, domain_type, cache_type {

      ignore_bins Ignore_inner_outer_sharable = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                                (binsof(domain_type) intersect {svt_axi_transaction::INNERSHAREABLE,
                                                                                svt_axi_transaction::OUTERSHAREABLE});

      ignore_bins Ignore_non_and_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                                   {svt_axi_transaction::READONCE,svt_axi_transaction::READSHARED,
                                                    svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                    svt_axi_transaction::READUNIQUE,svt_axi_transaction::CLEANUNIQUE,
                                                    svt_axi_transaction::MAKEUNIQUE,svt_axi_transaction::DVMCOMPLETE,
                                                    svt_axi_transaction::DVMMESSAGE}) && 
                                                   (binsof(domain_type) intersect {svt_axi_transaction::NONSHAREABLE,
                                                                                   svt_axi_transaction::SYSTEMSHAREABLE});
      ignore_bins Ignore_invalid_cache_barrier = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER,
                                                  svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE}) && 
                                                  (!binsof(cache_type) intersect {4'b0010});

      ignore_bins Ignore_invalid_cache = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOSNOOP}) && 
                                         (!binsof(cache_type) intersect {4'b0010,4'b0011,4'b0110,4'b0111,
                                                                         4'b1010,4'b1011,4'b1110,4'b1111});

      ignore_bins Ig_device_nonshare_cache = binsof(coherent_read_xact_type.coherent_readnosnoop_xact) && 
                                            (binsof(cache_type) intersect {4'b0000,4'b0001});

      ignore_bins Ig_device_non_system_shareable = (binsof(cache_type) intersect {4'b0000,4'b0001}) &&
                                                   (!binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE}); 

      ignore_bins Ig_cacheable_system_shareable = (binsof(cache_type) intersect {4'b0110,4'b0111,
                                                                                 4'b1010,4'b1011,4'b1110,4'b1111}) &&
                                                  (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
      
      
`ifdef SVT_ACE5_ENABLE
      ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID,svt_axi_transaction::CLEANSHAREDPERSIST}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`else
     ignore_bins Ignore_system_sharable = (binsof(coherent_read_xact_type) intersect 
                                           {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANINVALID,
                                            svt_axi_transaction::MAKEINVALID}) && 
                                            (binsof(domain_type) intersect {svt_axi_transaction::SYSTEMSHAREABLE});
`endif

      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif

 /**
  * Covergroup     : trans_cross_ace_arsnoop_arbar
  *
  * Coverpoints:
  *
  * - coherent_read_xact_type:  Captures coherent read transaction
  * - barrier_type : Captures read barrier
  * .
  * Cross coverpoints:
  * - arsnoop_arbar : Crosses cover points
  *    coherent_read_xact_type and barrier_type
  * .
  */

  //covergroup trans_cross_ace_arsnoop_arbar @(cov_read_sample_event);

  `ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_ace_arsnoop_arbar ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_TYPE

    arsnoop_arbar : cross coherent_read_xact_type, barrier_type {

      ignore_bins Ignore_normal = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});

      ignore_bins Ignore_barrier = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER}) && 
                                   (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                    svt_axi_transaction::SYNC_BARRIER});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  `else
  covergroup trans_cross_ace_arsnoop_arbar_dvm_unset ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_SET

    arsnoop_arbar : cross coherent_read_xact_type, barrier_type {

      ignore_bins Ignore_normal = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});

      ignore_bins Ignore_barrier = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER}) && 
                                   (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                    svt_axi_transaction::SYNC_BARRIER});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_arbar_dvm_set ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_SET

    arsnoop_arbar : cross coherent_read_xact_type, barrier_type {

      ignore_bins Ignore_normal = (binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});

      ignore_bins Ignore_barrier = (!binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READBARRIER}) && 
                                   (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                    svt_axi_transaction::SYNC_BARRIER});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  `endif

 /**
  *  Covergroup     : trans_cross_ace_arsnoop_coh_rresp
  *
  * Coverpoints:
  *
  * - coherent_read_xact_type:  Captures coherent read transaction
  * - coh_rresp : Captures read coherent response
  * .
  * Cross coverpoints:
  * - arsnoop_arburst_coh_rresp : Crosses cover points
  *    coherent_read_xact_type and coh_rresp
  * .
  */

  //covergroup trans_cross_ace_arsnoop_coh_rresp @(cov_read_sample_event);
  
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF  
  covergroup trans_cross_ace_arsnoop_coh_rresp (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_RRESP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_coh_rresp : cross coherent_read_xact_type, coh_rresp, slave_port_id {
      ignore_bins Ignore_invalid_rresp_ud_sc_sd = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READNOSNOOP,
                                                   svt_axi_transaction::CLEANUNIQUE,svt_axi_transaction::MAKEUNIQUE,
                                                   svt_axi_transaction::MAKEINVALID,svt_axi_transaction::READBARRIER,
                                                   svt_axi_transaction::CLEANINVALID} &&
                                                 !binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_CLEAN };

      ignore_bins Ignore_invalid_rresp_sc_sd = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READUNIQUE} &&
                                                 binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::SHARED_CLEAN,svt_axi_transaction::SHARED_DIRTY};

`ifdef SVT_ACE5_ENABLE 
      ignore_bins Ignore_invalid_rresp_ud_sd   = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READONCE,svt_axi_transaction::CLEANSHAREDPERSIST,
                                                   svt_axi_transaction::READCLEAN,svt_axi_transaction::CLEANSHARED} &&
                                                 binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_DIRTY,svt_axi_transaction::SHARED_DIRTY};
`else 
      ignore_bins Ignore_invalid_rresp_ud_sd   = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READONCE,
                                                   svt_axi_transaction::READCLEAN,svt_axi_transaction::CLEANSHARED} &&
                                                 binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_DIRTY,svt_axi_transaction::SHARED_DIRTY};
`endif 

      ignore_bins Ignore_invalid_rresp_sd   =   binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOTSHAREDDIRTY} &&
                                                  binsof(coh_rresp) intersect {svt_axi_transaction::SHARED_DIRTY};

      ignore_bins Ignore_dvm_xact_type      =   binsof(coherent_read_xact_type) intersect {
                                                 svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE};
                                   
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else
  covergroup trans_cross_ace_arsnoop_coh_rresp_def (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_RRESP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_coh_rresp : cross coherent_read_xact_type, coh_rresp , slave_port_id{
      ignore_bins Ignore_invalid_rresp_ud_sc_sd = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READNOSNOOP,
                                                   svt_axi_transaction::CLEANUNIQUE,svt_axi_transaction::MAKEUNIQUE,
                                                   svt_axi_transaction::MAKEINVALID,svt_axi_transaction::READBARRIER,
                                                   svt_axi_transaction::CLEANINVALID} &&
                                                 !binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_CLEAN };

      ignore_bins Ignore_invalid_rresp_sc_sd = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READUNIQUE} &&
                                                 binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::SHARED_CLEAN,svt_axi_transaction::SHARED_DIRTY};


      ignore_bins Ignore_invalid_rresp_sd   =   binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOTSHAREDDIRTY} &&
                                                  binsof(coh_rresp) intersect {svt_axi_transaction::SHARED_DIRTY};

      ignore_bins Ignore_dvm_xact_type      =   binsof(coherent_read_xact_type) intersect {
                                                 svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE};
                                   
`ifdef SVT_ACE5_ENABLE 
      ignore_bins Ignore_invalid_rresp_ud_sd   = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READONCE,svt_axi_transaction::CLEANSHAREDPERSIST,
                                                   svt_axi_transaction::READCLEAN,svt_axi_transaction::CLEANSHARED} &&
                                                 binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_DIRTY,svt_axi_transaction::SHARED_DIRTY};
`else 
      ignore_bins Ignore_invalid_rresp_ud_sd   = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READONCE,
                                                   svt_axi_transaction::READCLEAN,svt_axi_transaction::CLEANSHARED} &&
                                                 binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_DIRTY,svt_axi_transaction::SHARED_DIRTY};
`endif 
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_coh_rresp_dvm_unset_barrier_set (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_RRESP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_coh_rresp : cross coherent_read_xact_type, coh_rresp , slave_port_id{
      ignore_bins Ignore_invalid_rresp_ud_sc_sd = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READNOSNOOP,
                                                   svt_axi_transaction::CLEANUNIQUE,svt_axi_transaction::MAKEUNIQUE,
                                                   svt_axi_transaction::MAKEINVALID,svt_axi_transaction::READBARRIER,
                                                   svt_axi_transaction::CLEANINVALID} &&
                                                 !binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_CLEAN };

      ignore_bins Ignore_invalid_rresp_sc_sd = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READUNIQUE} &&
                                                 binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::SHARED_CLEAN,svt_axi_transaction::SHARED_DIRTY};


      ignore_bins Ignore_invalid_rresp_sd   =   binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOTSHAREDDIRTY} &&
                                                  binsof(coh_rresp) intersect {svt_axi_transaction::SHARED_DIRTY};

      ignore_bins Ignore_dvm_xact_type      =   binsof(coherent_read_xact_type) intersect {
                                                 svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE};
                                   
`ifdef SVT_ACE5_ENABLE 
      ignore_bins Ignore_invalid_rresp_ud_sd   = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READONCE,svt_axi_transaction::CLEANSHAREDPERSIST,
                                                   svt_axi_transaction::READCLEAN,svt_axi_transaction::CLEANSHARED} &&
                                                 binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_DIRTY,svt_axi_transaction::SHARED_DIRTY};
`else 
      ignore_bins Ignore_invalid_rresp_ud_sd   = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READONCE,
                                                   svt_axi_transaction::READCLEAN,svt_axi_transaction::CLEANSHARED} &&
                                                 binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_DIRTY,svt_axi_transaction::SHARED_DIRTY};
`endif 
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_coh_rresp_dvm_set_barrier_unset (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_RRESP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_coh_rresp : cross coherent_read_xact_type, coh_rresp , slave_port_id{
      ignore_bins Ignore_invalid_rresp_ud_sc_sd = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READNOSNOOP,
                                                   svt_axi_transaction::CLEANUNIQUE,svt_axi_transaction::MAKEUNIQUE,
                                                   svt_axi_transaction::MAKEINVALID,svt_axi_transaction::READBARRIER,
                                                   svt_axi_transaction::CLEANINVALID} &&
                                                 !binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_CLEAN };

      ignore_bins Ignore_invalid_rresp_sc_sd = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READUNIQUE} &&
                                                  binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::SHARED_CLEAN,svt_axi_transaction::SHARED_DIRTY};

  
      ignore_bins Ignore_invalid_rresp_sd   =   binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOTSHAREDDIRTY} &&
                                                  binsof(coh_rresp) intersect {svt_axi_transaction::SHARED_DIRTY};

      ignore_bins Ignore_dvm_xact_type      =   binsof(coherent_read_xact_type) intersect {
                                                 svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE};
                                   
`ifdef SVT_ACE5_ENABLE 
      ignore_bins Ignore_invalid_rresp_ud_sd   = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READONCE,svt_axi_transaction::CLEANSHAREDPERSIST,
                                                   svt_axi_transaction::READCLEAN,svt_axi_transaction::CLEANSHARED} &&
                                                 binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_DIRTY,svt_axi_transaction::SHARED_DIRTY};
`else 
      ignore_bins Ignore_invalid_rresp_ud_sd   = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READONCE,
                                                   svt_axi_transaction::READCLEAN,svt_axi_transaction::CLEANSHARED} &&
                                                 binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_DIRTY,svt_axi_transaction::SHARED_DIRTY};
`endif 
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_coh_rresp_dvm_set_barrier_set (int num_slaves);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_RRESP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SLAVE_PORT_ID

    arsnoop_coh_rresp : cross coherent_read_xact_type, coh_rresp , slave_port_id{
      ignore_bins Ignore_invalid_rresp_ud_sc_sd = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READNOSNOOP,
                                                   svt_axi_transaction::CLEANUNIQUE,svt_axi_transaction::MAKEUNIQUE,
                                                   svt_axi_transaction::MAKEINVALID,svt_axi_transaction::READBARRIER,
                                                   svt_axi_transaction::CLEANINVALID} &&
                                                 !binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_CLEAN };

      ignore_bins Ignore_invalid_rresp_sc_sd = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READUNIQUE} &&
                                                  binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::SHARED_CLEAN,svt_axi_transaction::SHARED_DIRTY};

      ignore_bins Ignore_invalid_rresp_sd   =   binsof(coherent_read_xact_type) intersect {svt_axi_transaction::READNOTSHAREDDIRTY} &&
                                                  binsof(coh_rresp) intersect {svt_axi_transaction::SHARED_DIRTY};

      ignore_bins Ignore_dvm_xact_type      =   binsof(coherent_read_xact_type) intersect {
                                                 svt_axi_transaction::DVMMESSAGE,svt_axi_transaction::DVMCOMPLETE};
                                   
 `ifdef SVT_ACE5_ENABLE 
      ignore_bins Ignore_invalid_rresp_ud_sd   = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READONCE,svt_axi_transaction::CLEANSHAREDPERSIST,
                                                   svt_axi_transaction::READCLEAN,svt_axi_transaction::CLEANSHARED} &&
                                                 binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_DIRTY,svt_axi_transaction::SHARED_DIRTY};
`else 
      ignore_bins Ignore_invalid_rresp_ud_sd   = binsof(coherent_read_xact_type) intersect {
                                                   svt_axi_transaction::READONCE,
                                                   svt_axi_transaction::READCLEAN,svt_axi_transaction::CLEANSHARED} &&
                                                 binsof(coh_rresp) intersect {
                                                   svt_axi_transaction::UNIQUE_DIRTY,svt_axi_transaction::SHARED_DIRTY};
`endif 
     option.weight = 1;
    }
    option.per_instance = 1;
  endgroup  

`endif
 /**
  *
  * Covergroup     : trans_cross_ace_ardvmmessage_ardvmresp
  * 
  * Coverpoints:
  *
  * - ardvm_message_type : Captures DVM message on araddr[14:12]
  *
  * - ardvm_resp       : Capture DVM response on rresp [4:0],
  *                        accept = 4'b0000 and reject = 4'b0010 
  * .
  *
  * Cross coverpoints:
  * - ardvmmessage_ardvmresp  : Crosses cover points ardvm_message_type and ardvm_resp
  * .
  *
  */

  //covergroup trans_cross_ace_ardvmmessage_ardvmresp @(cov_read_sample_event);
  covergroup trans_cross_ace_ardvmmessage_ardvmresp ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVMMESSAGE_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_DVM_RESPONSE_TYPE
     ardvmmessage_ardvmresp : cross ardvm_message_type, ardvm_resp {

        ignore_bins Ignore_dvm_hint_msg_resp = (binsof(ardvm_message_type) intersect {3'b110, 3'b100}) &&
                                               (binsof(ardvm_resp) intersect {4'b0010});
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

 /**
  *  Covergroup     : trans_cross_ace_arsnoop_cacheinitialstate_cachefinalstate
  *
  * Coverpoints:
  *
  * - coherent_read_xact_type  :  Captures coherent read transaction
  * - initial_cache_line_state : Captures initial cache line state
  * - final_cache_line_state   : Capture final cache line state
  * .
  * Cross coverpoints:
  * - arsnoop_cacheinitialstate_cachefinalstate : Crosses cover points
  *    coherent_read_xact_type initial_cache_line_state and final_cache_line_state
  * .
  */

  //covergroup trans_cross_ace_arsnoop_cacheinitialstate_cachefinalstate @(cov_read_sample_event);
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF  
  covergroup trans_cross_ace_arsnoop_cacheinitialstate_cachefinalstate ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_FINAL_CACHE_LINE_STATE

      arsnoop_cacheinitialstate_cachefinalstate : cross coherent_read_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {

     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_READ_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_READONCE_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_READCLEAN_XACT_TYPE_CROSS  
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_READNOTSHAREDDIRTY_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_READSHARED_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_READUNIQUE_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_CLEANUNIQUE_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_MAKEUNIQUE_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_CLEANSHARED_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_CLEANINVALID_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_MAKEINVALID_XACT_TYPE_CROSS 

    ignore_bins Ignore_speculative_initial_states  = ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE,
                                                       svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                       svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID}))||
                                                     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANUNIQUE}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY})) ||
                                                    ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::MAKEUNIQUE}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY}));
`ifdef SVT_ACE5_ENABLE 
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID}));
`else 
   ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID}));
`endif
 
    ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READBARRIER,svt_axi_transaction::DVMCOMPLETE,
                                                       svt_axi_transaction::DVMMESSAGE};


      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_update_cache_cacheinitialstate_cachefinalstate ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_FINAL_CACHE_LINE_STATE

      arsnoop_update_cache_cacheinitialstate_cachefinalstate : cross coherent_read_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_UPDATE_CACHE_COHERENT_READ_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_READONCE_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_READCLEAN_XACT_TYPE_CROSS  
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_READNOTSHAREDDIRTY_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_READSHARED_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_READUNIQUE_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_CLEANUNIQUE_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_MAKEUNIQUE_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_CLEANSHARED_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_CLEANINVALID_XACT_TYPE_CROSS
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_MAKEINVALID_XACT_TYPE_CROSS
    

    ignore_bins Ignore_speculative_initial_states  = ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE,
                                                       svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                       svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID}))||
                                                     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANUNIQUE}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY})) ||
                                                    ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::MAKEUNIQUE}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY}));

    ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READBARRIER,svt_axi_transaction::DVMCOMPLETE,
                                                       svt_axi_transaction::DVMMESSAGE};


`ifdef SVT_ACE5_ENABLE 
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID}));
`else 
   ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID}));
`endif
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else

  covergroup trans_cross_ace_arsnoop_cacheinitialstate_cachefinalstate_def ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_FINAL_CACHE_LINE_STATE

      arsnoop_cacheinitialstate_cachefinalstate : cross coherent_read_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {

      ignore_bins Ignore_readnosnoop_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUECLEAN})); 

      ignore_bins Ignore_readonce_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})); 

      ignore_bins Ignore_readclean_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN})); 

      ignore_bins Ignore_readnotshareddirty_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY,
                                                    svt_axi_transaction::SHAREDCLEAN})); 

      ignore_bins Ignore_readshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY,
                                                    svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY}));

      ignore_bins Ignore_readunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY}));

      ignore_bins Ignore_cleanunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ;

     ignore_bins Ignore_makeunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN,
                                                     svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ;
`ifdef SVT_ACE5_ENABLE 
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED, svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`else
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`endif

    ignore_bins Ignore_cleaninvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_makeinvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_speculative_initial_states  = ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE,
                                                       svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                       svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID}))||
                                                     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANUNIQUE}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY})) ||
                                                    ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::MAKEUNIQUE}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY}));

    ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READBARRIER,svt_axi_transaction::DVMCOMPLETE,
                                                       svt_axi_transaction::DVMMESSAGE};


      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_cacheinitialstate_cachefinalstate_def_speculative_read_enable ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DEF
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_FINAL_CACHE_LINE_STATE

      arsnoop_cacheinitialstate_cachefinalstate : cross coherent_read_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {
    ignore_bins Ignore_readnosnoop_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUECLEAN})) || 
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})));

      ignore_bins Ignore_readonce_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                              ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))); 
                
       ignore_bins Ignore_readclean_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))); 

       ignore_bins Ignore_readnotshareddirty_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::UNIQUEDIRTY})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})));
 
        ignore_bins Ignore_readshared_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))); 

      ignore_bins Ignore_readunique_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}))); 



      ignore_bins Ignore_cleanunique_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY,svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}))) ;
                                               

     ignore_bins Ignore_makeunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN,
                                                     svt_axi_transaction::SHAREDDIRTY,svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ;
    ignore_bins Ignore_cleaninvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_makeinvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READBARRIER,svt_axi_transaction::DVMCOMPLETE,
                                                       svt_axi_transaction::DVMMESSAGE};

  `ifdef SVT_ACE5_ENABLE 
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED, svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`else
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`endif
    option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_cacheinitialstate_cachefinalstate_dvm_unset_barrier_set ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_FINAL_CACHE_LINE_STATE

      arsnoop_cacheinitialstate_cachefinalstate : cross coherent_read_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {

      ignore_bins Ignore_readnosnoop_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUECLEAN})); 

      ignore_bins Ignore_readonce_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})); 

      ignore_bins Ignore_readclean_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN})); 

      ignore_bins Ignore_readnotshareddirty_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY,
                                                    svt_axi_transaction::SHAREDCLEAN})); 

      ignore_bins Ignore_readshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY,
                                                    svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY}));

      ignore_bins Ignore_readunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY}));

      ignore_bins Ignore_cleanunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ;

     ignore_bins Ignore_makeunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN,
                                                     svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ;


    ignore_bins Ignore_cleaninvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_makeinvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_speculative_initial_states  = ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE,
                                                       svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                       svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID}))||
                                                     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANUNIQUE}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY})) ||
                                                    ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::MAKEUNIQUE}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY}));

     ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READBARRIER,svt_axi_transaction::DVMCOMPLETE,
                                                       svt_axi_transaction::DVMMESSAGE};


  `ifdef SVT_ACE5_ENABLE 
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED, svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`else
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`endif
    option.weight = 1;
    }
    option.per_instance = 1;
  endgroup  
  covergroup trans_cross_ace_arsnoop_cacheinitialstate_cachefinalstate_dvm_unset_barrier_set_speculative_read_enable ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_UNSET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_FINAL_CACHE_LINE_STATE

      arsnoop_cacheinitialstate_cachefinalstate : cross coherent_read_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {

    ignore_bins Ignore_readnosnoop_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUECLEAN})) || 
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})));

      ignore_bins Ignore_readonce_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                              ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))); 
                
       ignore_bins Ignore_readclean_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))); 

       ignore_bins Ignore_readnotshareddirty_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::UNIQUEDIRTY})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})));
 
        ignore_bins Ignore_readshared_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))); 

      ignore_bins Ignore_readunique_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}))); 



      ignore_bins Ignore_cleanunique_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY,svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}))) ;
                                               

     ignore_bins Ignore_makeunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN,
                                                     svt_axi_transaction::SHAREDDIRTY,svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ;


    ignore_bins Ignore_cleaninvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_makeinvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READBARRIER,svt_axi_transaction::DVMCOMPLETE,
                                                       svt_axi_transaction::DVMMESSAGE};

   `ifdef SVT_ACE5_ENABLE 
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED, svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`else
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`endif
   option.weight = 1;
    }
    option.per_instance = 1;
  endgroup  


  covergroup trans_cross_ace_arsnoop_cacheinitialstate_cachefinalstate_dvm_set_barrier_unset ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_FINAL_CACHE_LINE_STATE

      arsnoop_cacheinitialstate_cachefinalstate : cross coherent_read_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {

      ignore_bins Ignore_readnosnoop_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUECLEAN})); 

      ignore_bins Ignore_readonce_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})); 

      ignore_bins Ignore_readclean_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN})); 

      ignore_bins Ignore_readnotshareddirty_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY,
                                                    svt_axi_transaction::SHAREDCLEAN})); 

      ignore_bins Ignore_readshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY,
                                                    svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY}));

      ignore_bins Ignore_readunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY}));

      ignore_bins Ignore_cleanunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ;

     ignore_bins Ignore_makeunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN,
                                                     svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ;

 
    ignore_bins Ignore_cleaninvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_makeinvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_speculative_initial_states  = ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE,
                                                       svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                       svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID}))||
                                                     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANUNIQUE}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY})) ||
                                                    ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::MAKEUNIQUE}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY}));

    ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READBARRIER,svt_axi_transaction::DVMCOMPLETE,
                                                       svt_axi_transaction::DVMMESSAGE};


`ifdef SVT_ACE5_ENABLE 
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED, svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`else
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`endif
      option.weight = 1;
    }
    option.per_instance = 0;
  endgroup
  covergroup trans_cross_ace_arsnoop_cacheinitialstate_cachefinalstate_dvm_set_barrier_unset_speculative_read_enable ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_FINAL_CACHE_LINE_STATE

      arsnoop_cacheinitialstate_cachefinalstate : cross coherent_read_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {

    ignore_bins Ignore_readnosnoop_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUECLEAN})) || 
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})));

      ignore_bins Ignore_readonce_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                              ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))); 
                
       ignore_bins Ignore_readclean_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))); 

       ignore_bins Ignore_readnotshareddirty_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::UNIQUEDIRTY})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})));
 
        ignore_bins Ignore_readshared_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))); 

      ignore_bins Ignore_readunique_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}))); 



      ignore_bins Ignore_cleanunique_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY,svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}))) ;
                                               

     ignore_bins Ignore_makeunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN,
                                                     svt_axi_transaction::SHAREDDIRTY,svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ;

      ignore_bins Ignore_cleaninvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_makeinvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READBARRIER,svt_axi_transaction::DVMCOMPLETE,
                                                       svt_axi_transaction::DVMMESSAGE};


 `ifdef SVT_ACE5_ENABLE 
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED, svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`else
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`endif
     option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_arsnoop_cacheinitialstate_cachefinalstate_dvm_set_barrier_set ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_FINAL_CACHE_LINE_STATE

      arsnoop_cacheinitialstate_cachefinalstate : cross coherent_read_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {

      ignore_bins Ignore_readnosnoop_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUECLEAN})); 

      ignore_bins Ignore_readonce_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})); 

      ignore_bins Ignore_readclean_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN})); 

      ignore_bins Ignore_readnotshareddirty_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY,
                                                    svt_axi_transaction::SHAREDCLEAN})); 

      ignore_bins Ignore_readshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY,
                                                    svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY}));

      ignore_bins Ignore_readunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY}));

      ignore_bins Ignore_cleanunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ;

     ignore_bins Ignore_makeunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN,
                                                     svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ;


    ignore_bins Ignore_cleaninvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_makeinvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_speculative_initial_states  = ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READNOSNOOP,svt_axi_transaction::READONCE,
                                                       svt_axi_transaction::READCLEAN,svt_axi_transaction::READNOTSHAREDDIRTY,
                                                       svt_axi_transaction::READSHARED,svt_axi_transaction::READUNIQUE}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID}))||
                                                     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANUNIQUE}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY})) ||
                                                    ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::MAKEUNIQUE}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY}));

    ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READBARRIER,svt_axi_transaction::DVMCOMPLETE,
                                                       svt_axi_transaction::DVMMESSAGE};


 `ifdef SVT_ACE5_ENABLE 
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED, svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`else
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`endif
     option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
  covergroup trans_cross_ace_arsnoop_cacheinitialstate_cachefinalstate_dvm_set_barrier_set_speculative_read_enable ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_READ_XACT_TYPE_DVM_SET_BARRIER_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_FINAL_CACHE_LINE_STATE

      arsnoop_cacheinitialstate_cachefinalstate : cross coherent_read_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {

      ignore_bins Ignore_readnosnoop_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUECLEAN})) || 
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})));

      ignore_bins Ignore_readonce_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                              ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READONCE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))); 
                
       ignore_bins Ignore_readclean_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READCLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))); 

       ignore_bins Ignore_readnotshareddirty_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::UNIQUEDIRTY})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READNOTSHAREDDIRTY}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})));
 
        ignore_bins Ignore_readshared_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))); 

      ignore_bins Ignore_readunique_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY})) || 
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                             ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                                ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::READUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}))); 



      ignore_bins Ignore_cleanunique_states = (((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY,svt_axi_transaction::UNIQUEDIRTY}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}))) ;
                                               

     ignore_bins Ignore_makeunique_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN,
                                                     svt_axi_transaction::SHAREDDIRTY,svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY})) ;

        ignore_bins Ignore_cleaninvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

    ignore_bins Ignore_makeinvalid_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::MAKEINVALID}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ;

     ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::READBARRIER,svt_axi_transaction::DVMCOMPLETE,
                                                       svt_axi_transaction::DVMMESSAGE};


  `ifdef SVT_ACE5_ENABLE 
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED, svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED,svt_axi_transaction::CLEANSHAREDPERSIST}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`else
      ignore_bins Ignore_cleanshared_states = ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||  
                                               ((binsof(coherent_read_xact_type) intersect
                                                    {svt_axi_transaction::CLEANSHARED}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}));
    ignore_bins Ignore_invalid_initial_state   =     ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANSHARED}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY})) ||                                                      
                                                      ((binsof(coherent_read_xact_type) intersect
                                                      {svt_axi_transaction::CLEANINVALID,svt_axi_transaction::MAKEINVALID}) &&
                                                      (!binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID})); 

`endif
    option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif

 /**
  *  Covergroup     : trans_cross_ace_awsnoop_cacheinitialstate_cachefinalstate
  *
  * Coverpoints:
  *
  * - coherent_write_xact_type  :  Captures coherent Write transaction
  * - initial_cache_line_state : Captures initial cache line state
  * - final_cache_line_state   : Capture final cache line state
  *                              INVALID,UNIQUECLEAN,SHAREDCLEAN are the possible final states
  * .
  * Cross coverpoints:
  * - awsnoop_cacheinitialstate_cachefinalstate : Crosses cover points
  *    coherent_write_xact_type initial_cache_line_state and final_cache_line_state
  * .
  */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF 
  covergroup trans_cross_ace_awsnoop_cacheinitialstate_cachefinalstate ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE

    final_cache_line_state : coverpoint cov_item.final_cache_line_state iff (cov_final_cache_line_state_flag) { 
      bins final_state_invalid          = {svt_axi_transaction::INVALID};
      bins final_state_uniqueclean      = {svt_axi_transaction::UNIQUECLEAN};
      bins final_state_sharedclean      = {svt_axi_transaction::SHAREDCLEAN};
      option.weight = 1 ;
    }

    awsnoop_cacheinitialstate_cachefinalstate : cross coherent_write_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {
                                                          
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_WRITE_XACT_TYPE_CROSS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_WRITEUNIQUEORLINE_XACT_TYPE_CROSS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_WRITEBACK_XACT_TYPE_CROSS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_WRITEEVICT_XACT_TYPE_CROSS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_WRITECLEAN_XACT_TYPE_CROSS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_EVICT_XACT_TYPE_CROSS 

       ignore_bins Ignore_invalid_initial_state   =  ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITENOSNOOP}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY}))||                                                      ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))||
                                                     ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITECLEAN}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN,
                                                       svt_axi_transaction::UNIQUECLEAN})) ||
                                                     ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::EVICT}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUEDIRTY,
                                                       svt_axi_transaction::SHAREDDIRTY})); 


        ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEBARRIER};          
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_update_cache_cacheinitialstate_cachefinalstate;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE

    final_cache_line_state : coverpoint cov_item.final_cache_line_state iff (cov_final_cache_line_state_flag) { 
      bins final_state_invalid          = {svt_axi_transaction::INVALID};
      bins final_state_uniqueclean      = {svt_axi_transaction::UNIQUECLEAN};
      bins final_state_sharedclean      = {svt_axi_transaction::SHAREDCLEAN};
      option.weight = 1 ;
    }

    awsnoop_update_cache_cacheinitialstate_cachefinalstate : cross coherent_write_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {
                                                         
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_UPDATE_CACHE_COHERENT_WRITE_XACT_TYPE_CROSS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_WRITEUNIQUEORLINE_XACT_TYPE_CROSS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_WRITEBACK_XACT_TYPE_CROSS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_WRITEEVICT_XACT_TYPE_CROSS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_WRITECLEAN_XACT_TYPE_CROSS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_IGNORE_COHERENT_EVICT_XACT_TYPE_CROSS

       ignore_bins Ignore_invalid_initial_state   =  ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITENOSNOOP}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY}))||                                                      ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))||
                                                     ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITECLEAN}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN,
                                                       svt_axi_transaction::UNIQUECLEAN})) ||
                                                     ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::EVICT}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUEDIRTY,
                                                       svt_axi_transaction::SHAREDDIRTY})); 


        ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEBARRIER};          
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  covergroup trans_cross_ace_awsnoop_not_ace_lite_no_barrier_no_writeevict_cacheinitialstate_cachefinalstate ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_FINAL_CACHE_LINE_STATE

    awsnoop_cacheinitialstate_cachefinalstate : cross coherent_write_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {
      
       ignore_bins Ignore_writenosnoop_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITENOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITENOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY}) &&                                                  (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}));

       ignore_bins Ignore_writeuniqueorline_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEUNIQUE,
                                                    svt_axi_transaction::WRITELINEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEUNIQUE,
                                                    svt_axi_transaction::WRITELINEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}) &&                                                  (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}));

       ignore_bins Ignore_writeback_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEBACK}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}));

        ignore_bins Ignore_writeevict_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEEVICT}) &&
                                               (!binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) ) ||
                                                ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEEVICT}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}));

       ignore_bins Ignore_writeclean_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITECLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                               ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITECLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}));

       ignore_bins evict_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::EVICT}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}));

       ignore_bins Ignore_invalid_initial_state   =  ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITENOSNOOP}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY}))||                                                      ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))||
                                                     ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITECLEAN}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN,
                                                       svt_axi_transaction::UNIQUECLEAN})) ||
                                                     ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::EVICT}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUEDIRTY,
                                                       svt_axi_transaction::SHAREDDIRTY})); 


        ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEBARRIER};          
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_no_barrier_writeevict_cacheinitialstate_cachefinalstate ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE
    
    // For write type transactions such as WRITENOSNOOP, WRITEUNIQUE,
    // WRITELINEUNIQUE, WRITECLEAN, WRITEBACK, EVICT and WRITEEVICT, the possible
    // final states are INVALID, UNIQUECLEAN and SHAREDCLEAN. So Dirty states
    // are not included.
    final_cache_line_state : coverpoint cov_item.final_cache_line_state iff (cov_final_cache_line_state_flag) { 
      bins final_state_invalid          = {svt_axi_transaction::INVALID}; 
      bins final_state_uniqueclean      = {svt_axi_transaction::UNIQUECLEAN}; 
      bins final_state_sharedclean      = {svt_axi_transaction::SHAREDCLEAN}; 
      option.weight = 1 ; 
    }
    
    awsnoop_cacheinitialstate_cachefinalstate : cross coherent_write_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {
      
       ignore_bins Ignore_writenosnoop_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITENOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITENOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY}) &&                                                  (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}));

       ignore_bins Ignore_writeuniqueorline_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEUNIQUE,
                                                    svt_axi_transaction::WRITELINEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEUNIQUE,
                                                    svt_axi_transaction::WRITELINEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}) &&                                                  (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}));

       ignore_bins Ignore_writeback_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEBACK}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}));

       ignore_bins Ignore_writeevict_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEEVICT}) &&
                                               (!binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) ) ||
                                                ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEEVICT}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}));

       ignore_bins Ignore_writeclean_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITECLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                               ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITECLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}));

       ignore_bins evict_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::EVICT}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}));

       ignore_bins Ignore_invalid_initial_state   =  ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITENOSNOOP}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY}))||                                                      ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))||
                                                     ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITECLEAN}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN,
                                                       svt_axi_transaction::UNIQUECLEAN})) ||
                                                     ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::EVICT}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUEDIRTY,
                                                       svt_axi_transaction::SHAREDDIRTY})); 


        ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEBARRIER};          
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_barrier_no_writeevict_cacheinitialstate_cachefinalstate ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_FINAL_CACHE_LINE_STATE

    awsnoop_cacheinitialstate_cachefinalstate : cross coherent_write_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {
      
       ignore_bins Ignore_writenosnoop_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITENOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITENOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY}) &&                                                  (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}));

       ignore_bins Ignore_writeuniqueorline_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEUNIQUE,
                                                    svt_axi_transaction::WRITELINEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEUNIQUE,
                                                    svt_axi_transaction::WRITELINEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}) &&                                                  (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}));

       ignore_bins Ignore_writeback_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEBACK}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}));

       ignore_bins Ignore_writeevict_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEEVICT}) &&
                                               (!binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) ) ||
                                                ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEEVICT}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}));

       ignore_bins Ignore_writeclean_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITECLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                               ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITECLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}));

       ignore_bins evict_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::EVICT}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}));

       ignore_bins Ignore_invalid_initial_state   =  ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITENOSNOOP}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY}))||                                                      ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))||
                                                     ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITECLEAN}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN,
                                                       svt_axi_transaction::UNIQUECLEAN})) ||
                                                     ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::EVICT}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUEDIRTY,
                                                       svt_axi_transaction::SHAREDDIRTY})); 


        ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEBARRIER};          
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_awsnoop_not_ace_lite_barrier_writeevict_cacheinitialstate_cachefinalstate ;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_FINAL_CACHE_LINE_STATE

    awsnoop_cacheinitialstate_cachefinalstate : cross coherent_write_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {
      
       ignore_bins Ignore_writenosnoop_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITENOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITENOSNOOP}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::UNIQUEDIRTY}) &&                                                  (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}));

       ignore_bins Ignore_writeuniqueorline_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEUNIQUE,
                                                    svt_axi_transaction::WRITELINEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}) &&     
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID})) ||
                                               ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEUNIQUE,
                                                    svt_axi_transaction::WRITELINEUNIQUE}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}) &&                                                  (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}));

       ignore_bins Ignore_writeback_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEBACK}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}));

       ignore_bins Ignore_writeevict_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEEVICT}) &&
                                               (!binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                                ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITEEVICT}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}));


       ignore_bins Ignore_writeclean_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITECLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUEDIRTY}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN})) ||
                                               ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::WRITECLEAN}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDDIRTY}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::SHAREDCLEAN}));

       ignore_bins evict_states = ((binsof(coherent_write_xact_type) intersect
                                                    {svt_axi_transaction::EVICT}) &&
                                               (binsof(initial_cache_line_state) intersect 
                                                    {svt_axi_transaction::UNIQUECLEAN,svt_axi_transaction::SHAREDCLEAN}) &&  
                                               (!binsof(final_cache_line_state) intersect 
                                                    {svt_axi_transaction::INVALID}));

       ignore_bins Ignore_invalid_initial_state   =  ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITENOSNOOP}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::SHAREDCLEAN,svt_axi_transaction::SHAREDDIRTY}))||                                                      ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::WRITELINEUNIQUE}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::UNIQUEDIRTY,svt_axi_transaction::SHAREDDIRTY}))||
                                                     ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEBACK,svt_axi_transaction::WRITECLEAN}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID,svt_axi_transaction::SHAREDCLEAN,
                                                       svt_axi_transaction::UNIQUECLEAN})) ||
                                                     ((binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::EVICT}) &&
                                                      (binsof(initial_cache_line_state) intersect 
                                                      {svt_axi_transaction::INVALID,svt_axi_transaction::UNIQUEDIRTY,
                                                       svt_axi_transaction::SHAREDDIRTY})); 


        ignore_bins Ignore_invalid_xact_types      =     binsof(coherent_write_xact_type) intersect
                                                      {svt_axi_transaction::WRITEBARRIER};          
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

 /**
  *  Covergroup     : trans_cross_ace_acsnoop_cacheinitialstate_cachefinalstate
  *
  * Coverpoints:
  *
  * - snoop_xact_type  :  Captures Snoop transaction
  * - initial_cache_line_state : Captures initial cache line state
  * - final_cache_line_state   : Capture final cache line state
  * .
  * Cross coverpoints:
  * - acsnoop_cacheinitialstate_cachefinalstate : Crosses cover points
  *    snoop_xact_type initial_cache_line_state and final_cache_line_state
  * .
  */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF

  covergroup trans_cross_ace_acsnoop_cacheinitialstate_cachefinalstate @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_FINAL_CACHE_LINE_STATE

    acsnoop_cacheinitialstate_cachefinalstate : cross snoop_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CACHE_STATE_IGNORE_BINS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CACHE_STATE_ONE_ACE_ACELITE_IGNORE_BINS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_IGNORE_BINS
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /** 
   * This covergroup will be created when there is only one ACE-master and
   * minimum one or more than one ACE_LITE master in the system. 
   */
  covergroup trans_cross_ace_acsnoop_cacheinitialstate_cachefinalstate_one_ace_acelite @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_ONE_ACE_ACELITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_FINAL_CACHE_LINE_STATE

    acsnoop_cacheinitialstate_cachefinalstate : cross snoop_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CACHE_STATE_ONE_ACE_ACELITE_IGNORE_BINS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_IGNORE_BINS
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

`else //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF 
  covergroup trans_cross_ace_acsnoop_dvm_unset_cacheinitialstate_cachefinalstate @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_UNSET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_FINAL_CACHE_LINE_STATE

    acsnoop_cacheinitialstate_cachefinalstate : cross snoop_xact_type, initial_cache_line_state ,
                                                      final_cache_line_state {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CACHE_STATE_IGNORE_BINS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CACHE_STATE_ONE_ACE_ACELITE_IGNORE_BINS
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /** 
   * This covergroup will be created when there is only one ACE-master and
   * minimum one or more than one ACE_LITE master in the system. 
   */
  covergroup trans_cross_ace_acsnoop_dvm_unset_cacheinitialstate_cachefinalstate_one_ace_acelite @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_UNSET_ONE_ACE_ACELITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_FINAL_CACHE_LINE_STATE

    acsnoop_cacheinitialstate_cachefinalstate : cross snoop_xact_type, initial_cache_line_state ,
                                                      final_cache_line_state {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CACHE_STATE_ONE_ACE_ACELITE_IGNORE_BINS
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_ace_acsnoop_dvm_set_cacheinitialstate_cachefinalstate @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_SET
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_FINAL_CACHE_LINE_STATE

    acsnoop_cacheinitialstate_cachefinalstate : cross snoop_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CACHE_STATE_IGNORE_BINS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CACHE_STATE_ONE_ACE_ACELITE_IGNORE_BINS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_IGNORE_BINS
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /** 
   * This covergroup will be created when there is only one ACE-master and
   * minimum one or more than one ACE_LITE master in the system. 
   */
  covergroup trans_cross_ace_acsnoop_dvm_set_cacheinitialstate_cachefinalstate_one_ace_acelite @(cov_snoop_sample_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_XACT_TYPE_DVM_SET_ONE_ACE_ACELITE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_INITIAL_CACHE_LINE_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_FINAL_CACHE_LINE_STATE

    acsnoop_cacheinitialstate_cachefinalstate : cross snoop_xact_type, initial_cache_line_state ,
                                                        final_cache_line_state {
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_CACHE_STATE_ONE_ACE_ACELITE_IGNORE_BINS
      `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACSNOOP_DVM_IGNORE_BINS
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup
`endif //SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  
 /**
  *
  * Covergroup     : trans_cross_stream_xact_type_tid_tdest
  * 
  * Coverpoints:
  *
  * - stream_xact_type: Captures the type of stream 
  *
  * - stream_tid: Captures the value of TID 
  *
  * - stream_tdest: Captures the value of TDEST
  * .
  *
  * Cross coverpoints:
  * - trans_cross_stream_xact_type_tid_tdest: Crosses cover points
  * stream_xact_type, stream_tid and stream_tdest
  * .
  *
  */

  covergroup trans_cross_stream_xact_type_tid_tdest @(cov_stream_sample_event);
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_STREAM_XACT_TYPE
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_STREAM_TID
     `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_STREAM_TDEST
     trans_cross_stream_xact_type_tid: cross stream_xact_type, stream_tid {
       option.weight = 1;
     }
     trans_cross_stream_xact_type_tdest: cross stream_xact_type, stream_tdest {
       option.weight = 1;
     }
     trans_cross_stream_xact_type_tid_tdest: cross stream_xact_type, stream_tid, stream_tdest {
      option.weight = 1;
     }
    option.per_instance = 1;
  endgroup

  // ****************************************************************************
  // Exception Covergroups
  // ****************************************************************************

  /**
  *  ----------------------------------------------------------------------------
  *  Covergroup     : trans_cross_axi_awburst_awlen_awaddr_exceptions
  *  ----------------------------------------------------------------------------
  */  
  //covergroup trans_cross_axi_awburst_awlen_awaddr_exceptions ;
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_XACT_TYPE
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR
  //  //`SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_EXCEPTIONS
  //  axi_awburst_awlen_awaddr_exceptions : cross xact_type, burst_type, burst_length, addr, axi_exceptions {
  //    ignore_bins ign_read_xact = !binsof(xact_type.write_xact);
  //    option.weight = 1;
  //  }
  //  option.per_instance = 1;
  //endgroup

  /**
  *  ----------------------------------------------------------------------------
  *  Covergroup     : trans_cross_axi_awburst_awlen_bresp_exceptions
  *  ----------------------------------------------------------------------------
  */  
  //covergroup trans_cross_axi_awburst_awlen_bresp_exceptions ;
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_XACT_TYPE
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP
  //  //`SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_EXCEPTIONS
  //  axi_awburst_awlen_bresp_exceptions : cross xact_type, burst_type, burst_length, bresp, axi_exceptions {
  //    ignore_bins ign_read_xact = !binsof(xact_type.write_xact);
  //    option.weight = 1;
  //  }
  //  option.per_instance = 1;
  //endgroup

  /**
  *  ----------------------------------------------------------------------------
  *  Covergroup     : trans_cross_axi_arburst_arlen_araddr_exceptions
  *  ----------------------------------------------------------------------------
  */  
  //covergroup trans_cross_axi_arburst_arlen_araddr_exceptions @(cov_read_sample_event);
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_XACT_TYPE
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ADDR
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_EXCEPTIONS
  //  axi_arburst_arlen_araddr_exceptions : cross xact_type, burst_type, burst_length, addr, axi_exceptions {
  //    ignore_bins ign_write_xact = !binsof(xact_type.read_xact);
  //    option.weight = 1;
  //  }
  //  option.per_instance = 1;
  //endgroup
  /**
  *  ----------------------------------------------------------------------------
  *  Covergroup     : trans_cross_axi_arburst_arlen_rresp_exceptions
  *  ----------------------------------------------------------------------------
  */  
  //covergroup trans_cross_axi_arburst_arlen_rresp_exceptions @(cov_read_sample_event);
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_XACT_TYPE
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_TYPE
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BURST_LENGTH
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BRESP
  //  `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_EXCEPTIONS
  //  axi_arburst_arlen_bresp_exceptions : cross xact_type, burst_type, burst_length, bresp, axi_exceptions {
  //    ignore_bins ign_write_xact = !binsof(xact_type.read_xact);
  //    option.weight = 1;
  //  }
  //  option.per_instance = 1;
  //endgroup

 /**
  *  Covergroup     : trans_outstanding_read_with_same_id_to_different_slaves
  *
  * Coverpoints:
  *
  * - axi_outstanding_read_with_same_id_to_different_slaves: This is covered when:
  *   - A master issues two outstanding read transactions with the same ID 
  *   - These read transactions are targeted to two different slaves
  *   .
  * .
  * Note that this covergroup is constructed for all master interface types.<br>
  * Also note that this covergroup is constructed only if the number of slaves
  * in the system (svt_axi_system_configuration::num_slaves) is greater than 1.<br>
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613
  */
  covergroup trans_outstanding_read_with_same_id_to_different_slaves @(cov_outstanding_read_with_same_id_to_different_slaves_sample_event);
    axi_outstanding_read_with_same_id_to_different_slaves: coverpoint outstanding_read_with_same_id_to_different_slaves {
      bins outstanding_with_same_id_to_different_slaves = {1};
    }
    option.per_instance = 1;
  endgroup // trans_outstanding_read_with_same_id_to_different_slaves

 /**
  *  Covergroup     : trans_outstanding_write_with_same_id_to_different_slaves
  *
  * Coverpoints:
  *
  * - axi_outstanding_write_with_same_id_to_different_slaves: This is covered when:
  *   - A master issues two outstanding write transactions with the same ID 
  *   - These write transactions are targeted to two different slaves
  *   .
  * .
  * Note that this covergroup is constructed for all master interface types.<br>
  * Also note that this covergroup is constructed only if the number of slaves
  * in the system (svt_axi_system_configuration::num_slaves) is greater than 1.<br>  
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613
  */
  covergroup trans_outstanding_write_with_same_id_to_different_slaves @(cov_outstanding_write_with_same_id_to_different_slaves_sample_event);
    axi_outstanding_write_with_same_id_to_different_slaves: coverpoint outstanding_write_with_same_id_to_different_slaves {
      bins outstanding_with_same_id_to_different_slaves = {1};
    }
    option.per_instance = 1;
  endgroup // trans_outstanding_write_with_same_id_to_different_slaves

 /**
  *  Covergroup     : trans_ar_aw_stalled_for_ac_channel
  *
  * Coverpoints:
  *
  * - axi_ar_aw_stalled_for_ac_channel: This is covered when read transaction on AR channel 
  *   OR WriteUnique/WriteLineUnique transactions on AW channel from a master are stalled 
  *   by interconnect, while waiting for the snoop response from the same master.
  * .
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C6.6.1
  */
  covergroup trans_ar_aw_stalled_for_ac_channel @(cov_ar_aw_stalled_for_ac_channel_sample_event);
    axi_ar_aw_stalled_for_ac_channel: coverpoint ar_aw_stalled_for_ac_channel {
      bins readonce_stalled_for_snoop = {1};
      bins readshared_stalled_for_snoop = {2};
      bins readclean_stalled_for_snoop = {3};
      bins readnotshareddirty_stalled_for_snoop = {4};
      bins readunique_stalled_for_snoop = {5};
      bins cleanunique_stalled_for_snoop = {6};
      bins makeunique_stalled_for_snoop = {7};
      bins cleanshared_stalled_for_snoop = {8};
      bins cleaninvalid_stalled_for_snoop = {9};
      bins makeinvalid_stalled_for_snoop = {10};
`ifdef SVT_ACE5_ENABLE 
      bins cleansharedpersist_stalled_for_snoop = {14};
`endif
      bins writeunique_stalled_for_snoop = {15};
      bins writelineunique_stalled_for_snoop = {16};
    }
    option.per_instance = 1;
  endgroup // trans_ar_aw_stalled_for_ac_channel

 /**
  *  Covergroup     : trans_xact_domain_after_nonshareable_barrier
  *
  * Coverpoints:
  *
  * - axi_xact_domain_after_nonshareable_barrier: This is covered when:
  *   - Master initiates non-shareable transaction followed by non-shareable read/write barrier pairs
  *   - Before the barrier completes, the same master initiates any other coherent transactions with 
  *     inner/outer/system domains
  *   .
  * .
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C8.2.2
  */
  covergroup trans_xact_domain_after_nonshareable_barrier @(cov_xact_domain_after_nonshareable_barrier_sample_event);
    axi_xact_domain_after_nonshareable_barrier: coverpoint xact_domain_after_nonshareable_barrier {
      bins nonshareable_read_barrier_followed_by_innershareable_read_xact = {1};
      bins nonshareable_read_barrier_followed_by_outershareable_read_xact = {2};
      bins nonshareable_read_barrier_followed_by_systemshareable_read_xact = {3};
      bins nonshareable_write_barrier_followed_by_innershareable_write_xact = {5};
      bins nonshareable_write_barrier_followed_by_outershareable_write_xact = {6};
      bins nonshareable_write_barrier_followed_by_systemshareable_write_xact = {7};
    }
    option.per_instance = 1;
  endgroup

 /**
  *  Covergroup     : trans_xact_domain_after_innershareable_barrier
  *
  * Coverpoints:
  *
  * - axi_xact_domain_after_innershareable_barrier: This is covered when:
  *   - Master initiates inner-shareable transaction followed by inner-shareable read/write barrier pairs
  *   - Before the barrier completes, the same master initiates any other coherent transactions with 
  *     none/outer/system domains
  *   .  
  * .
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C8.2.2
  */
  covergroup trans_xact_domain_after_innershareable_barrier @(cov_xact_domain_after_innershareable_barrier_sample_event);
    axi_xact_domain_after_innershareable_barrier: coverpoint xact_domain_after_innershareable_barrier {
      bins innershareable_read_barrier_followed_by_nonshareable_read_xact = {0};
      bins innershareable_read_barrier_followed_by_outershareable_read_xact = {2};
      bins innershareable_read_barrier_followed_by_systemshareable_read_xact = {3};
      bins innershareable_write_barrier_followed_by_nonshareable_write_xact = {4};
      bins innershareable_write_barrier_followed_by_outershareable_write_xact = {6};
      bins innershareable_write_barrier_followed_by_systemshareable_write_xact = {7};
    }
    option.per_instance = 1;
  endgroup

 /**
  *  Covergroup     : trans_xact_domain_after_outershareable_barrier
  *
  * Coverpoints:
  *
  * - axi_xact_domain_after_outershareable_barrier: This is covered when:
  *   - Master initiates outer-shareable transaction followed by outer-shareable read/write barrier pairs
  *   - Before the barrier completes, the same master initiates any other coherent transactions with 
  *     none/inner/system domains
  *   .   
  * .
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C8.2.2
  */
  covergroup trans_xact_domain_after_outershareable_barrier @(cov_xact_domain_after_outershareable_barrier_sample_event);
    axi_xact_domain_after_outershareable_barrier: coverpoint xact_domain_after_outershareable_barrier {
      bins outershareable_read_barrier_followed_by_nonshareable_read_xact = {0};
      bins outershareable_read_barrier_followed_by_innershareable_read_xact = {1};
      bins outershareable_read_barrier_followed_by_systemshareable_read_xact = {3};
      bins outershareable_write_barrier_followed_by_nonshareable_write_xact = {4};
      bins outershareable_write_barrier_followed_by_innershareable_write_xact = {5};
      bins outershareable_write_barrier_followed_by_systemshareable_write_xact = {7};
    }
    option.per_instance = 1;
  endgroup

 /**
  *  Covergroup     : trans_xact_domain_after_systemshareable_barrier
  *
  * Coverpoints:
  *
  * - axi_xact_domain_after_systemshareable_barrier:  This is covered when:
  *   - Master initiates system-shareable transaction followed by system-shareable read/write barrier pairs
  *   - Before the barrier completes, the same master initiates any other coherent transactions with 
  *     inner/outer/systemnone domains
  *   .    
  * .
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C8.2.2
  */
  covergroup trans_xact_domain_after_systemshareable_barrier @(cov_xact_domain_after_systemshareable_barrier_sample_event);
    axi_xact_domain_after_systemshareable_barrier: coverpoint xact_domain_after_systemshareable_barrier {
      bins systemshareable_read_barrier_followed_by_nonshareable_read_xact = {0};
      bins systemshareable_read_barrier_followed_by_innershareable_read_xact = {1};
      bins systemshareable_read_barrier_followed_by_outershareable_read_xact = {2};
      bins systemshareable_write_barrier_followed_by_nonshareable_write_xact = {4};
      bins systemshareable_write_barrier_followed_by_innershareable_write_xact = {5};
      bins systemshareable_write_barrier_followed_by_outershareable_write_xact = {6};
    }
    option.per_instance = 1;
  endgroup

 /**
  *  Covergroup     : trans_xact_ordering_after_barrier
  *
  * Coverpoints:
  *
  * - axi_xact_ordering_after_barrier: This is covered when a master issues transactions 
  *   between issuing a barrier transaction on the address channel and receiving the read 
  *   and write barrier responses. 
  *   - Such transactions have no ordering guarantee with respect to the barrier. On the address 
  *     channel, these transactions are permitted to remain after the barrier transaction or they 
  *     are permitted to overtake the barrier transaction.
  *   .
  * .
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C8.4.1
  */
  covergroup trans_xact_ordering_after_barrier @(cov_xact_ordering_after_barrier_sample_event);
    axi_xact_ordering_after_barrier: coverpoint xact_ordering_after_barrier {
      bins read_xact_overtake_barrier_response = {0};
      bins read_xact_fallbehind_barrier_response = {1};
      bins write_xact_overtake_barrier_response = {2};
      bins write_xact_fallbehind_barrier_response = {3};
    }
    option.per_instance = 1;
  endgroup
  
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
 /**
  * Covergroup: trans_ace_barrier_outstanding_xact<br>
  * Coverpoints:<br>
  * barrier_outstanding_xact : Captures total number of read and write barrier outstanding
  * transactions. When svt_axi_port_configuration::axi_interface_type is configured as
  * AXI_ACE maximum number of 256 outstanding transactions is tracked. When
  * svt_axi_port_configuration::axi_interface_type is configured as ACE_LITE, outstanding
  * transactions greater than 256 are also tracked. 
  * This is as per section C8.4.1 of AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613" 
  */
  covergroup trans_ace_barrier_outstanding_xact @(cov_barrier_outstanding_event);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_OUTSTANDING_TRANSACTION
    option.per_instance = 1;
  endgroup

`else
/**
  * Covergroup: trans_ace_barrier_outstanding_xact_ace<br>
  * Coverpoints:<br>
  * barrier_outstanding_xact : Captures total number of read and write barrier outstanding
  * transactions. When svt_axi_port_configuration::axi_interface_type is configured as
  * AXI_ACE maximum number of 256 outstanding transactions is tracked. When
  * svt_axi_port_configuration::axi_interface_type is configured as ACE_LITE, outstanding
  * transactions greater than 256 are also tracked. 
  * This is as per section C8.4.1 of AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613" 
  */
  covergroup trans_ace_barrier_outstanding_xact_ace @(cov_barrier_outstanding_event_ace);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_OUTSTANDING_TRANSACTION_ACE
    option.per_instance = 1;
  endgroup
 /**
  * Covergroup: trans_ace_barrier_outstanding_xact_acelite<br>
  * Coverpoints:<br>
  * barrier_outstanding_xact : Captures total number of read and write barrier outstanding
  * transactions. When svt_axi_port_configuration::axi_interface_type is configured as
  * AXI_ACE maximum number of 256 outstanding transactions is tracked. When
  * svt_axi_port_configuration::axi_interface_type is configured as ACE_LITE, outstanding
  * transactions greater than 256 are also tracked. 
  * This is as per section C8.4.1 of AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613" 
  */
  covergroup trans_ace_barrier_outstanding_xact_acelite @(cov_barrier_outstanding_event_acelite);
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_OUTSTANDING_TRANSACTION_ACELITE
    option.per_instance = 1;
  endgroup
`endif
  /**
  * Covergroup: trans_non_barrier_xact_after_256_outstanding_barrier_xact<br>
  * Coverpoints:<br>
  * -non_barrier_after_256_outstanding_barrier_xact: Captures if active transactions on write channel occur
  * after 256 barrier outstanding transactions are accepted by slave component
  * .
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C8.4.2
  */
  covergroup trans_non_barrier_xact_after_256_outstanding_barrier_xact @(cov_non_barrier_after_256_outstanding_barrier_sample_event);
    non_barrier_after_256_outstanding_barrier_xact : coverpoint non_barrier_after_256_outstanding_barrier{
      bins write_xact_after_256_outstanding_barrier_xact = {1};
    }
    option.per_instance = 1;
  endgroup

  /**
  * Covergroup: trans_master_back_to_back_write_ordering <br>
  * Coverpoints:<br>
  * -xact_back_to_back_write_ordering: Captures if back-to-back write transactions with the same id
  * is observed
  * .
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C1.3.4
  */
  covergroup trans_master_back_to_back_write_ordering @(cov_master_back_to_back_write_ordering_event);
    xact_back_to_back_write_ordering: coverpoint back_to_back_write_ordering {
      bins back_to_back_write_with_same_id = {0};
    }
    option.per_instance = 1;
  endgroup

  /**
  * Covergroup: trans_master_write_after_read_ordering <br>
  * Coverpoints:<br>
  * -xact_back_to_back_write_ordering: Captures the order of completion of a write transaction issued after
  * a read 
  * .
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C1.3.4
  */
  covergroup trans_master_write_after_read_ordering @(cov_master_write_after_read_ordering_event);
    xact_write_after_read_ordering : coverpoint write_after_read_ordering {
      bins write_after_read_with_write_completing_first = {0};
      bins write_after_read_with_read_completing_first = {1};
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_master_snoop_to_same_address_as_read_xact <br>
    *
    * Coverpoints:<br>
    * -read_xact_to_same_address_as_snoop: Captures read transactions to the same address as a snoop to the master. 
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C5.2.5
    */
  covergroup trans_master_snoop_to_same_address_as_read_xact;
    read_xact_to_same_address_as_snoop: coverpoint read_xact_to_same_address_as_snoop {
      bins coherent_readnosnoop_xact   = {0}; 
      bins coherent_readonce_xact   = {1}; 
      bins coherent_readshared_xact   = {2}; 
      bins coherent_readclean_xact   = {3}; 
      bins coherent_readnotshareddirty_xact   = {4}; 
      bins coherent_readunique_xact   = {5}; 
      bins coherent_cleanunique_xact   = {6}; 
      bins coherent_makeunique_xact   = {7}; 
      bins coherent_cleanshared_xact   = {8}; 
      bins coherent_cleaninvalid_xact   = {9}; 
      bins coherent_makeinvalid_xact   = {10};
`ifdef SVT_ACE5_ENABLE
      bins coherent_cleansharedpersist_xact = {11};
`endif
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_master_snoop_to_same_addr_as_memory_update_exclude_writeevict <br>
    *
    * Coverpoints:<br>
    * -memory_update_excluding_writeevict: Captures
    * WRITEBACK,WRITECLEAN,EVICT,WRITEUNIQUE and WRITELINEUNIQUE transactions
    * to the same address as a snoop. WRITENOSNOOP transactions to non
    * overlapping addresses are captured because WRITENOSNOOP is issued to
    * non-shareable region and another master may not access the same address
    * as that of a WRITENOSNOOP through a snoop. 
    * -snoop_xact_type: Captures snoop transactions other than DVM transactions
    * - trans_cross_memory_update_snoop_xact_to_same_address: Crosses memory_update_excluding_writeevict and snoop_xact_type 
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C6.6.1
    */
   covergroup trans_master_snoop_to_same_addr_as_memory_update_exclude_writeevict; 
    `SVT_AXI_PORT_MONITOR_DEV_COV_UTIL_MEMORY_UPDATE_EXCLUDING_WRITEEVICT_CP
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_ADDR_PHASE_XACT_TYPE_DVM_UNSET
    trans_cross_memory_update_snoop_xact_to_same_address : cross memory_update_excluding_writeevict, snoop_xact_type {
      option.weight = 1;
    }
    option.per_instance = 1;

  endgroup

    /**
    * Covergroup: trans_master_snoop_to_same_addr_as_memory_update_exclude_writeevict_one_ace_acelite <br>
    * This covergroup will be created when there is only one ACE-master and
    * minimum one or more than one ACE_LITE master in the system.
    * Coverpoints:<br>
    * -memory_update_excluding_writeevict: Captures
    * WRITEBACK,WRITECLEAN,EVICT,WRITEUNIQUE and WRITELINEUNIQUE transactions
    * to the same address as a snoop. WRITENOSNOOP transactions to non
    * overlapping addresses are captured because WRITENOSNOOP is issued to
    * non-shareable region and another master may not access the same address
    * as that of a WRITENOSNOOP through a snoop. 
    * -snoop_xact_type:Coverpoint of svt_axi_snoop_transaction::snoop_xact_type for READONCE,CLEANSHARED,CLEANINVALID and MAKEINVALID snoop transactions recieved on master port . This excludes READSHARED,READCLEAN,READNOTSHAREDDIRTY,READUNIQUE,DVMMESSAGE,DVMCOMPLETE transactions
    * - trans_cross_memory_update_snoop_xact_to_same_address: Crosses memory_update_excluding_writeevict and snoop_xact_type 
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C6.6.1
    */
   covergroup trans_master_snoop_to_same_addr_as_memory_update_exclude_writeevict_one_ace_acelite; 
    `SVT_AXI_PORT_MONITOR_DEV_COV_UTIL_MEMORY_UPDATE_EXCLUDING_WRITEEVICT_CP
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_ADDR_PHASE_XACT_TYPE_DVM_UNSET_ONE_ACE_ACELITE
    trans_cross_memory_update_snoop_xact_to_same_address : cross memory_update_excluding_writeevict, snoop_xact_type {
      option.weight = 1;
    }
    option.per_instance = 1;

  endgroup

  /**
    * Covergroup: trans_master_snoop_to_same_addr_as_writeevict<br>
    *
    * Coverpoints:<br>
    * -write_evict_xact: Captures WRITEEVICT transactions to the same address
    * as a snoop.  
    * -snoop_xact_type: Captures snoop transactions other than DVM transactions
    * - trans_cross_writeevict_snoop_xact_to_same_address: Crosses write_evict_xact and snoop_xact_type 
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C6.6.1
    */
  covergroup trans_master_snoop_to_same_addr_as_writeevict;
    write_evict_xact: coverpoint write_xact_type_to_same_addr_as_snoop {
      bins coherent_writeevict_xact = {6};
    }
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_ADDR_PHASE_XACT_TYPE_DVM_UNSET
    trans_cross_writeevict_snoop_xact_to_same_address : cross write_evict_xact, snoop_xact_type {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_master_snoop_to_same_addr_as_writeevict_one_ace_acelite<br>
    * This covergroup will be created when there is only one ACE-master and
    * minimum one or more than one ACE_LITE master in the system.
    * Coverpoints:<br>
    * -write_evict_xact: Captures WRITEEVICT transactions to the same address
    * as a snoop.  
    * -snoop_xact_type:Coverpoint of svt_axi_snoop_transaction::snoop_xact_type for READONCE,CLEANSHARED,CLEANINVALID and MAKEINVALID snoop transactions recieved on master port . This excludes READSHARED,READCLEAN,READNOTSHAREDDIRTY,READUNIQUE,DVMMESSAGE,DVMCOMPLETE transactions
    * - trans_cross_writeevict_snoop_xact_to_same_address: Crosses write_evict_xact and snoop_xact_type 
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C6.6.1
    */
  covergroup trans_master_snoop_to_same_addr_as_writeevict_one_ace_acelite;
    write_evict_xact: coverpoint write_xact_type_to_same_addr_as_snoop {
      bins coherent_writeevict_xact = {6};
    }
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_ADDR_PHASE_XACT_TYPE_DVM_UNSET_ONE_ACE_ACELITE
    trans_cross_writeevict_snoop_xact_to_same_address : cross write_evict_xact, snoop_xact_type {
      option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_master_snoop_data_transfer_during_wu_wlu_to_same_addr <br>
    * Captures snoop responses with data transfer when a WRITEUNIQUE or WRITELINEUNIQUE to the same address
    * is in progress
    * Coverpoints: <br>
    * -snoop_xact_type: Captures snoop transactions other than DVM transactions and MAKEINVALID. MAKEINVALID transactions are not captured because it is recommended that MAKEINVALID does not transfer data.
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C5.2.5
    */
  covergroup trans_master_snoop_data_transfer_during_wu_wlu_to_same_addr;
   snoop_xact_type : coverpoint cov_snoop_item.snoop_xact_type iff(cov_snoop_xact_type_flag){ 
     bins snoop_readonce_xact   = {svt_axi_snoop_transaction::READONCE}; 
     bins snoop_readshared_xact   = {svt_axi_snoop_transaction::READSHARED}; 
     bins snoop_readclean_xact   = {svt_axi_snoop_transaction::READCLEAN}; 
     bins snoop_readnotshareddirty_xact   = {svt_axi_snoop_transaction::READNOTSHAREDDIRTY}; 
     bins snoop_readunique_xact   = {svt_axi_snoop_transaction::READUNIQUE}; 
     bins snoop_cleanshared_xact   = {svt_axi_snoop_transaction::CLEANSHARED}; 
     bins snoop_cleaninvalid_xact   = {svt_axi_snoop_transaction::CLEANINVALID}; 
     option.weight = 0; 
   }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_master_snoop_data_transfer_during_wu_wlu_to_same_addr_one_ace_acelite <br>
    * Captures snoop responses with data transfer when a WRITEUNIQUE or WRITELINEUNIQUE to the same address
    * is in progress, when only one ACE master and one or more ACE_LITE masters present in the system.
    * Coverpoints: <br>
    * -snoop_xact_type: Captures snoop transactions READONCE,CLEANSHARED,CLEANINVALID. Other transactions are not captured because ACE_LITE master cant fire READSHARED,READCLEAN,READNOTSHAREDDIRTY,READUNIQUE.
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C5.2.5
    */
  covergroup trans_master_snoop_data_transfer_during_wu_wlu_to_same_addr_one_ace_acelite;
   snoop_xact_type : coverpoint cov_snoop_item.snoop_xact_type iff(cov_snoop_xact_type_flag){ 
     bins snoop_readonce_xact   = {svt_axi_snoop_transaction::READONCE}; 
     bins snoop_cleanshared_xact   = {svt_axi_snoop_transaction::CLEANSHARED}; 
     bins snoop_cleaninvalid_xact   = {svt_axi_snoop_transaction::CLEANINVALID}; 
     option.weight = 0; 
   }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_master_readunique_snoop_resp_datatransfer_with_clean_cacheline<br>
    * Coverpoints: <br>
    * -snoop_resp_datatransfer_with_clean_cacheline: Captures whether data was
    * transferred for READUNIQUE snoop when the cache was in a clean state.
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C5.3.3
    */
  covergroup trans_master_readunique_snoop_resp_datatransfer_with_clean_cacheline @(cov_readunique_snoop_resp_datatransfer_with_clean_cacheline_event);
    snoop_resp_datatransfer_with_clean_cacheline: coverpoint cov_snoop_item.snoop_resp_datatransfer {
      bins snoop_no_datatransfer = {0};
      bins snoop_with_datatransfer = {1};
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_cross_awunique_awsnoop_awbar <br>
    * Coverpoints: <br>
    * - coherent_write_xact_type: Captures write transction type. Includes
    * WRITENOSNOOP, WRITEUNIQUE, WRITELINEUNIQUE, WRITECLEAN, WRITEBACK, EVICT,
    * WRITEBARRIER and WRITEEVICT
    * - awunique_val: Captures the value of signal AWUNIQUE in above transactions
    * - barrier_type: Captures the value of barrier type (AWBAR), in above transactions
    * - awunique_awsnoop_awbar: Cross of coherent_write_xact_type, awunique_val and barrier_type
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.1.4
    */
`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  covergroup trans_cross_awunique_awsnoop_awbar;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE
    awunique_val: coverpoint cov_item.is_unique iff (cov_coherent_xact_type_flag) {
      bins is_not_unique = {0};
      bins is_unique = {1}; 
    }
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_TYPE
    awunique_awsnoop_awbar : cross  coherent_write_xact_type, awunique_val, barrier_type {
      ignore_bins ignore_writeevict = binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEEVICT} && binsof(awunique_val) intersect {0};
      ignore_bins ignore_writeclean = binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITECLEAN} && binsof(awunique_val) intersect {1};
      // Ignore NORMAL_ACCESS_RESPECT_BARRIER and NORMAL_ACCESS_IGNORE_BARRIER for barrier transaction
      ignore_bins ignore_normal = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});
      // Ignore MEMORY_BARRIER and SYNC_BARRIER for non-barrier transaction
      ignore_bins ignore_barrier = (!binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});
    }
    option.per_instance = 1;
  endgroup
`else
  covergroup trans_cross_awunique_awsnoop_awbar_without_barrier;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_NO_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_TYPE
     awunique_val: coverpoint cov_item.is_unique {
      bins is_not_unique = {0};
      bins is_unique = {1}; 
     }
     awunique_awsnoop_awbar : cross  coherent_write_xact_type, awunique_val, barrier_type {
      ignore_bins ignore_writeevict = binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEEVICT} && binsof(awunique_val) intersect {0};
      ignore_bins ignore_writeclean = binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITECLEAN} && binsof(awunique_val) intersect {1};
    }
    option.per_instance = 1;
  endgroup

  covergroup trans_cross_awunique_awsnoop_awbar_with_barrier;
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_COHERENT_WRITE_XACT_TYPE_NOT_ACE_LITE_BARRIER_NO_WRITEEVICT
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_BARRIER_TYPE 
     awunique_val: coverpoint cov_item.is_unique {
      bins is_not_unique = {0};
      bins is_unique = {1}; 
     }
     awunique_awsnoop_awbar : cross  coherent_write_xact_type, awunique_val, barrier_type {
      ignore_bins ignore_writeevict = binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEEVICT} && binsof(awunique_val) intersect {0};
      ignore_bins ignore_writeclean = binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITECLEAN} && binsof(awunique_val) intersect {1};
      // Ignore NORMAL_ACCESS_RESPECT_BARRIER and NORMAL_ACCESS_IGNORE_BARRIER for barrier transaction
      ignore_bins ignore_normal = (binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,
                                                                   svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER});
      // Ignore MEMORY_BARRIER and SYNC_BARRIER for non-barrier transaction
      ignore_bins ignore_barrier = (!binsof(coherent_write_xact_type) intersect {svt_axi_transaction::WRITEBARRIER}) && 
                                  (binsof(barrier_type) intersect {svt_axi_transaction::MEMORY_BARRIER,
                                                                   svt_axi_transaction::SYNC_BARRIER});
    }
    option.per_instance = 1;
  endgroup
`endif

  /**
    * Covergroup: trans_master_snoop_resp_during_wu_wlu_to_same_addr<br>
    * Coverpoints: <br>
    * - snoop_crresp: Captures snoop response values 
    * - snoop_crresp_wu: Captures value of WasUnique bit in snoop response
    * - awunique_val: Captures the value of signal AWUNIQUE for WRITEUNIQUE and WRITELINEUNIQUE transactions
    * - snoop_resp_awunique: Cross of snoop_crresp, snoop_crresp_wu and awunique_val 
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C3.1.4
    */
  covergroup trans_master_snoop_resp_during_wu_wlu_to_same_addr;
    snoop_crresp : coverpoint cov_crresp[3:0] iff(cov_snoop_resp_flag){ 
      bins cresp_x0000 = {4'b0000}; 
      bins cresp_x1000 = {4'b1000}; 
      bins cresp_x0001 = {4'b0001}; 
      bins cresp_x1001 = {4'b1001}; 
      wildcard ignore_bins ig_invalid_cresp1 = {5'b??1?0};
      // WRITEUNIQUE, WRITELINEUNIQUE can be sent only when cache is in clean state
      ignore_bins ignore_pass_dirty = {4'b0101,4'b1101};
      option.weight = 0;
    }
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WASUNIQUE_SNOOP_RRESP_TYPE
     awunique_val: coverpoint write_xact_to_same_addr_as_snoop.is_unique {
      bins is_not_unique = {0};
      bins is_unique = {1}; 
     }
     // When AWUNIQUE is asserted a response that would allow another copy of the cacheline
     // to be created must not be given. So snoop_resp_datatransfer must be low when AWUNIQUE is high
     // So ignore bins that fulfill that condition
     // So ignore bins that fulfill that condition
     //when AWUNIQUE  is asserted snooped cache will not be able to retain its copy and will go in shared state .So Snoop
     // response is_shared bit must be driven low 
     snoop_resp_awunique : cross snoop_crresp, awunique_val  
     {
       ignore_bins ignore_snoop_data_transfer = binsof(snoop_crresp) intersect {4'b1001,4'b0001,4'b1000} && binsof(awunique_val) intersect {1};
     }
    option.per_instance = 1;
  endgroup

`ifndef SVT_AXI_MON_CFG_BASED_COV_GRP_DEF
  /**
    * Covergroup: trans_master_num_outstanding_dvm_syncs<br>
    * Coverpoints: <br>
    * - num_outstanding_dvm_sync_xacts: Captures number of outstanding dvm sync
    * snoop transactions. Note that a master is allowed to send only one
    * outstanding DVM sync transaction (ie, a DVM sync transaction to which a 
    * DVM complete is not yet received). Therefore a maximum of 256 outstanding
    * DVM sync snoop transactions is possible only in a system with atleast 257
    * masters capable of sending DVM transactions.
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C12.2
    */
  covergroup trans_master_num_outstanding_dvm_syncs @(cov_snoop_dvm_sync_event);
    num_outstanding_dvm_sync_xacts : coverpoint num_outstanding_dvm_syncs {
      bins outstanding_dvm_syncs_less_than_256 = {[1:255]};
      bins outstanding_dvm_syncs_equals_256 = {256}; 
      ignore_bins ignore_dvm_syncs_equal_256 = {256} iff (num_dvm_enabled_masters <= 256);
    }
    option.per_instance = 1;
  endgroup

`else 
 /**
    * Covergroup: trans_master_num_outstanding_dvm_syncs_num_dvm_enabled_masters_less_256<br>
    * Coverpoints: <br>
    * - num_outstanding_dvm_sync_xacts: Captures number of outstanding dvm sync
    * snoop transactions. Note that a master is allowed to send only one
    * outstanding DVM sync transaction (ie, a DVM sync transaction to which a 
    * DVM complete is not yet received). Therefore a maximum of 255 outstanding
    * DVM sync snoop transactions is possible only in a system with atleast 256
    * masters capable of sending DVM transactions.
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C12.2
    */
  covergroup trans_master_num_outstanding_dvm_syncs_num_dvm_enabled_masters_less_256 @(cov_snoop_dvm_sync_event);
    num_outstanding_dvm_sync_xacts : coverpoint num_outstanding_dvm_syncs {
      bins outstanding_dvm_syncs_less_than_256 = {[1:255]};
    }
    option.per_instance = 1;
  endgroup
/**
    * Covergroup:trans_master_num_outstanding_dvm_syncs_num_dvm_enbaled_master_256<br>
    * Coverpoints: <br>
    * - num_outstanding_dvm_sync_xacts: Captures number of outstanding dvm sync
    * snoop transactions. Note that a master is allowed to send only one
    * outstanding DVM sync transaction (ie, a DVM sync transaction to which a 
    * DVM complete is not yet received). Therefore a maximum of 256 outstanding
    * DVM sync snoop transactions is possible only in a system with atleast 257
    * masters capable of sending DVM transactions.
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C12.2
    */
  covergroup trans_master_num_outstanding_dvm_syncs_num_dvm_enbaled_master_256 @(cov_snoop_dvm_sync_event);
    num_outstanding_dvm_sync_xacts : coverpoint num_outstanding_dvm_syncs {
      bins outstanding_dvm_syncs_less_than_256 = {[1:255]};
      bins outstanding_dvm_syncs_equals_256 = {256}; 
    }
    option.per_instance = 1;
  endgroup
`endif

  /**
    * Covergroup: trans_master_concurrent_coherent_exclusive_access<br>
    * Coverpoints: <br>
    * - num_coherent_exl_access: Number of concurrent coherent exclusive accesses on different IDs
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C9.6
    */
  covergroup trans_master_concurrent_coherent_exclusive_access @ (cov_coherent_exclusive_read_access_event);
    num_coherent_exl_access : coverpoint num_coherent_excl_access_threads {
      bins one_thread = {1};
      bins more_than_one_thread = {[1:$]};
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_master_coherent_unmatched_excl_access<br>
    * Coverpoints: <br>
    * - unmatched_excl_access: Captures exclusive load accesses which did not
    * have a corresponding exclusive store access and exclusive store accesses
    * which did not have a corresponding exclusive load access. The
    * unmatched_excl_load_access is hit when a second exclusive load access to
    * the same ID is received before an exclusive store to that ID. The
    * unmatched_excl_store_access is hit when there is no prior exclusive load
    * to an exclusive store (CLEANUNIQUE) transaction. 
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C9.6
    */
  covergroup trans_master_coherent_unmatched_excl_access @(cov_coherent_unmatched_excl_access_event);
    unmatched_excl_access : coverpoint coherent_unmatched_excl_access_type {
      bins unmatched_excl_store_access = {0};
      bins unmatched_excl_load_access = {1};
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_master_barrier_id_reuse_for_non_barrier<br>
    * Coverpoints: <br>
    * - num_barrier_id_reuse_for_non_barrier: Captures the number of times that
    * the ID used for barrier transaction is reused for a normal transaction
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C8.4
    */
  covergroup trans_master_barrier_id_reuse_for_non_barrier @(cov_barrier_id_reuse_for_non_barrier_event);
    num_barrier_id_reuse_for_non_barrier : coverpoint num_barrier_id_reuse {
      bins barrier_id_reuse = {[1:$]};  
    }
    option.per_instance = 1;
  endgroup

    /** 
    * Covergroup: system_ace_coherent_and_snoop_association_recommended_ace 
    * 
    * Coverpoints: 
    * 
    * - ace_coh_and_snp_association:  This is covered when the interconnect issues recommended 
    *   snoop transaction to the snooped masters, in response to the coherent  
    *   transaction received from the initiating master.  
    * . 
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Table C6-1 
    * 
    */ 
  covergroup trans_master_ace_coherent_and_snoop_association_recommended_ace; 
    ace_coh_and_snp_association: coverpoint coh_and_snp_association { 
      bins readonce_coherent_to_readonce_snoop = {16'h01_00}; 
      bins readclean_coherent_to_readclean_snoop = {16'h03_02};  
      bins readnotshareddirty_coherent_to_readnotshareddirty_snoop = {16'h04_03}; 
      bins readshared_coherent_to_readshared_snoop = {16'h02_01}; 
      bins readunique_coherent_to_readunique_snoop = {16'h05_07}; 
      bins cleanunique_coherent_to_cleaninvalid_snoop = {16'h06_09}; 
      bins makeunique_coherent_to_makeinvalid_snoop = {16'h07_0d}; 
      bins cleanshared_coherent_to_cleanshared_snoop = {16'h08_08};
`ifdef SVT_ACE5_ENABLE
      bins cleansharedpersist_coherent_to_cleanshared_snoop = {16'h10_08};
`endif
      bins cleaninvalid_coherent_to_cleaninvalid_snoop = {16'h09_09}; 
      bins makeinvalid_coherent_to_makeinvalid_snoop = {16'h0a_0d}; 
      bins writeunique_coherent_to_cleaninvalid_snoop = {16'h0f_09}; 
      bins writelineunique_coherent_to_makeinvalid_snoop = {16'h10_0d}; 
    } 
    option.per_instance = 1; 
  endgroup 

  /** 
  * Covergroup: system_ace_coherent_and_snoop_association_recommended_ace_lite 
  * 
  * Coverpoints: 
  * 
  * - ace_coh_and_snp_association:  This is covered when the interconnect issues recommended 
  *   snoop transaction to the snooped masters, in response to the coherent  
  *   transaction received from the initiating master.  
  * . 
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Table C6-1 
  * 
  */ 
  covergroup trans_master_ace_coherent_and_snoop_association_recommended_ace_lite; 
    ace_coh_and_snp_association: coverpoint coh_and_snp_association { 
      bins readonce_coherent_to_readonce_snoop = {16'h01_00}; 
      bins cleanshared_coherent_to_cleanshared_snoop = {16'h08_08}; 
`ifdef SVT_ACE5_ENABLE
      bins cleansharedpersist_coherent_to_cleanshared_snoop = {16'h10_08};
`endif
      bins cleaninvalid_coherent_to_cleaninvalid_snoop = {16'h09_09}; 
      bins makeinvalid_coherent_to_makeinvalid_snoop = {16'h0a_0d}; 
      bins writeunique_coherent_to_cleaninvalid_snoop = {16'h0f_09}; 
      bins writelineunique_coherent_to_makeinvalid_snoop = {16'h10_0d}; 
    } 
    option.per_instance = 1; 
  endgroup

  /**
    * Covergroup: trans_master_ace_concurrent_readunique_cleanunique
    *
    * Coverpoints:
    *
    * - ace_concurrent_readunique_cleanunique:  This is covered when multiple ACE masters
    *   concurrently(that are simultaneously active) initiate ReadUnique or CleanUnique transactions.
    *
    * Two or more ACE masters needed for this covergroup
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C1.3.4 
    *
    */
  covergroup trans_master_ace_concurrent_readunique_cleanunique; 
    ace_concurrent_readunique_cleanunique: coverpoint concurrent_readunique_cleanunique {
      bins readunique_readunique = {16'h05_05};
      bins readunique_cleanunique = {16'h05_09,16'h09_05};
      bins cleanunique_cleannique = {16'h09_09};
    }
    option.per_instance = 1;
  endgroup

  /**
     * Covergroup: trans_master_ace_concurrent_overlapping_coherent_xacts
     * The covergroup trans_master_ace_concurrent_overlapping_coherent_xacts covers coherent transactions initiated from different ACE masters concurrently on the same address.
     * The covergroup needs atlease two ACE masters to be present in the system.
     * Coverpoints:
     *
     * - coherent_xact_on_ace_master_port:  This coverpoint covers svt_axi_transaction::coherent_xact_type transaction . All coherent transactions capable of generating snoop are bins of this coverpoint .
     * - coherent_xact_on_other_ace_master_port_in_system : This coverpoint covers svt_axi_transaction::coherent_xact_type transactions . All coherent transactions capable of generating snoop are bins of this coverpoint .
     * .
     *  Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; 
     */
  covergroup trans_master_ace_concurrent_overlapping_coherent_xacts ;
    coherent_xact_on_ace_master_port: coverpoint coherent_xact_on_port1{
      bins coherent_readonce_xact            = {svt_axi_transaction::READONCE} ;
      bins coherent_readshared_xact          = {svt_axi_transaction::READSHARED};
      bins coherent_readclean_xact           = {svt_axi_transaction::READCLEAN};
      bins coherent_readnotshareddirty_xact  = {svt_axi_transaction::READNOTSHAREDDIRTY};
      bins coherent_readunique_xact          = {svt_axi_transaction::READUNIQUE};
      bins coherent_cleanunique_xact         = {svt_axi_transaction::CLEANUNIQUE};
      bins coherent_makeunique_xact          = {svt_axi_transaction::MAKEUNIQUE};
      bins coherent_cleanshared_xact         = {svt_axi_transaction::CLEANSHARED};
`ifdef SVT_ACE5_ENABLE
      bins coherent_cleansharedpersist_xact = {svt_axi_transaction::CLEANSHAREDPERSIST};
`endif
      bins coherent_cleaninvalid_xact        = {svt_axi_transaction::CLEANINVALID};
      bins coherent_makeinvalid_xact         = {svt_axi_transaction::MAKEINVALID};
      bins coherent_writeunique_xact         = {svt_axi_transaction::WRITEUNIQUE};
      bins coherent_writelineunique_xact     = {svt_axi_transaction::WRITELINEUNIQUE};
    }
    
    coherent_xact_on_other_ace_master_port_in_system : coverpoint coherent_xact_on_port2{
      bins coherent_readonce_xact            = {svt_axi_transaction::READONCE} ;
      bins coherent_readshared_xact          = {svt_axi_transaction::READSHARED};
      bins coherent_readclean_xact           = {svt_axi_transaction::READCLEAN};
      bins coherent_readnotshareddirty_xact  = {svt_axi_transaction::READNOTSHAREDDIRTY};
      bins coherent_readunique_xact          = {svt_axi_transaction::READUNIQUE};
      bins coherent_cleanunique_xact         = {svt_axi_transaction::CLEANUNIQUE};
      bins coherent_makeunique_xact          = {svt_axi_transaction::MAKEUNIQUE};
      bins coherent_cleanshared_xact         = {svt_axi_transaction::CLEANSHARED};
`ifdef SVT_ACE5_ENABLE
      bins coherent_cleansharedpersist_xact = {svt_axi_transaction::CLEANSHAREDPERSIST};
`endif
      bins coherent_cleaninvalid_xact        = {svt_axi_transaction::CLEANINVALID};
      bins coherent_makeinvalid_xact         = {svt_axi_transaction::MAKEINVALID};
      bins coherent_writeunique_xact         = {svt_axi_transaction::WRITEUNIQUE};
      bins coherent_writelineunique_xact     = {svt_axi_transaction::WRITELINEUNIQUE};
    }
    
    ace_concurrent_overlapping: cross coherent_xact_on_ace_master_port ,coherent_xact_on_other_ace_master_port_in_system  {
      option.weight = 1;
    }
    option.per_instance = 1;
   endgroup
  
  /**
    * Covergroup: trans_master_ace_dirty_data_write
    * This is a system-level covergroup which works by enabling sys_cfg field system_ace_dirty_data_write_enable.
    * Coverpoints:
    *
    * - master_xact_of_ic_dirty_data_write:  This is covered when the interconnect issues a write
    * to the slave because dirty data was returned by one of the snoop responses and that
    * dirty data could not be returned to the master that initiated the original transaction 
    *
    * Two or more ACE masters needed for this covergroup
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; C 13.4 
    *
    */

  covergroup trans_master_ace_dirty_data_write;
    ace_dirty_data_write: coverpoint master_xact_of_ic_dirty_data_write.coherent_xact_type {
      bins readonce_dirty_data_write = {svt_axi_transaction::READONCE};
      bins readclean_dirty_data_write = {svt_axi_transaction::READCLEAN};
      bins readnotshreaddirty_dirty_data_write = {svt_axi_transaction::READNOTSHAREDDIRTY};
      bins cleaninvalid_dirty_data_write = {svt_axi_transaction::CLEANINVALID};
      bins cleanshared_dirty_data_write = {svt_axi_transaction::CLEANSHARED};
`ifdef SVT_ACE5_ENABLE
      bins cleansharedpersist_dirty_data_write = {svt_axi_transaction::CLEANSHAREDPERSIST};
`endif
      bins cleanunique_dirty_data_write = {svt_axi_transaction::CLEANUNIQUE};
      bins writeunique_dirty_data_write = {svt_axi_transaction::WRITEUNIQUE};
    }
    option.per_instance = 1;
  endgroup
  
  /**
    * Covergroup: trans_master_ace_dirty_data_write_one_ace_acelite
    * This is a system-level covergroup which works by enabling sys_cfg field system_ace_dirty_data_write_enable.
    * Coverpoints:
    *
    * - master_xact_of_ic_dirty_data_write:  This is covered when the interconnect issues a write
    * to the slave because dirty data was returned by one of the snoop responses and that
    * dirty data could not be returned to the master that initiated the original transaction 
    *
    * One ACE and one or more ACE_LITE masters needed for this covergroup
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; C 13.4 
    *
    */  
  covergroup trans_master_ace_dirty_data_write_one_ace_acelite;
    ace_dirty_data_write: coverpoint master_xact_of_ic_dirty_data_write.coherent_xact_type {
      bins readonce_dirty_data_write = {svt_axi_transaction::READONCE};
      bins cleaninvalid_dirty_data_write = {svt_axi_transaction::CLEANINVALID};
      bins cleanshared_dirty_data_write = {svt_axi_transaction::CLEANSHARED};
      bins writeunique_dirty_data_write = {svt_axi_transaction::WRITEUNIQUE};
    }
    option.per_instance = 1;
  endgroup

    /**
    * Covergroup: trans_master_ace_cross_cache_line_dirty_data_write
    *
    * Coverpoints:
    *
    * - ace_cross_cache_line_dirty_data_write:  This is covered under the following
    * conditions:
    *  - The interconnect may need to snoop multiple cachelines for a
    *  WRITEUNIQUE or READONCE transaction because it spans multiple cache
    *  lines
    *  - Atleast two of these snoop transactions return dirty data
    *  - The interconnect writes the dirty data of the snoop transactions to slave
    *
    * One or more ACE masters needed for this covergroup
    *  .
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; C 13.4 
    *
    */
  covergroup trans_master_ace_cross_cache_line_dirty_data_write; 
    ace_cross_cache_line_dirty_data_write: coverpoint master_xact_of_ic_dirty_data_write.coherent_xact_type {
      bins readonce_cross_cache_line_dirty_data_write = {svt_axi_transaction::READONCE};        
      bins writeunique_cross_cache_line_dirty_data_write = {svt_axi_transaction::WRITEUNIQUE};        
    }
    option.per_instance = 1;
  endgroup
   
  /**
    * Covergroup: trans_master_ace_snoop_and_memory_returns_data
    *
    * Coverpoints:
    *
    * - ace_snoop_and_memory_read_timing:  This cover point covers possible
    * relative timings of snoop generation by the interconnect with respect to
    * receiving speculative read data by the interconnect and bin snoop_returns_data_and_memory_not_returns_data 
    * covers if a transaction is found with snoop data transfer and without associated slave transaction. The 
    * various timings covered are:
    *  - snoop issued before the first read data beat is received through speculative read transaction
    *  - snoop issued after the last beat of read data is received through speculative read transaction
    *  - snoop issued while the read data is being received through speculative read transaction
    *  .
    * - ace_snoop_and_memory_returns_data_xact_type: Covers the various coherent
    * transaction types for which speculative read was issued. The transaction
    * types covered are READONCE, READCLEAN READNOSHAREDDIRTY, READUNIQUE and
    * READSHARED transactions
    *
    * At least two ACE masters needed for this covergroup
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; C 6.5.1 
    *
    */
  covergroup trans_master_ace_snoop_and_memory_returns_data;
    ace_snoop_and_memory_data_timing: coverpoint snoop_and_memory_read_timing {
      bins snoop_data_before_memory_data = {SNOOP_BEFORE_MEMORY_READ};
      bins snoop_data_along_with_memory_data = {SNOOP_ALONG_WITH_MEMORY_READ};
      bins snoop_data_after_memory_data = {SNOOP_AFTER_MEMORY_READ};
      bins snoop_returns_data_and_memory_not_returns_data = {SNOOP_RETURNS_DATA_AND_MEMORY_NOT_RETURNS_DATA};
    }

    ace_snoop_and_memory_returns_data_xact_type: coverpoint fully_correlated_master_xact.coherent_xact_type {
      bins readonce_snoop_and_memory_returns_data = {svt_axi_transaction::READONCE};
      bins readclean_snoop_and_memory_returns_data = {svt_axi_transaction::READCLEAN};
      bins readnotshreaddirty_snoop_and_memory_returns_data = {svt_axi_transaction::READNOTSHAREDDIRTY};
      bins readunique_snoop_and_memory_returns_data  = {svt_axi_transaction::READUNIQUE};
      bins readshared_snoop_and_memory_returns_data  = {svt_axi_transaction::READSHARED};
    }
    snoop_memory_timing_and_xact_cross : cross ace_snoop_and_memory_data_timing, ace_snoop_and_memory_returns_data_xact_type;
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_master_ace_write_during_speculative_fetch
    *
    * Coverpoints:
    *
    * - ace_write_during_speculative_fetch:  This cover point covers the following condition: 
    * A master issues a read transaction. This results in interconnect
    * generating snoop transactions towards other masters within the domain.
    * The interconnect also generates speculative read transaction for this
    * location. Speculative transaction returns data while the snoop
    * transactions do not return data. The snoop transactions may not return
    * data, either because there is no entry in the snooped masters' caches or
    * a WRITEBACK/WRITECLEAN of dirty data is in progress. The interconnect now
    * detects that a write transaction (the WRITEBACK/WRITECLEAN which is in
    * progress) is received for the same address for which it did a speculative
    * fetch. In such situation, interconnect performs another read from main
    * memory, as originally received data from speculative read is now stale
    *
    * At least One ACE master needed for this covergroup
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; C 6.5.1
    *
    */
  covergroup trans_master_ace_write_during_speculative_fetch;
    ace_write_during_speculative_fetch:
    coverpoint fully_correlated_master_xact.coherent_xact_type {
      bins overlapping_write_during_readonce = {svt_axi_transaction::READONCE};
      bins overlapping_write_during_readclean = {svt_axi_transaction::READCLEAN};
      bins overlapping_write_during_readnotshareddirty = {svt_axi_transaction::READNOTSHAREDDIRTY};
      bins overlapping_write_during_readunique = {svt_axi_transaction::READUNIQUE};
      bins overlapping_write_during_readshared = {svt_axi_transaction::READSHARED};
    }
    option.per_instance = 1;
  endgroup
  
  /**
    * Covergroup: trans_master_ace_xacts_with_high_priority_from_other_master_during_barrier
    *
    * Coverpoints:
    * - ace_xacts_with_high_priority_from_other_master_during_barrier:  
    * This cover point covers the following condition: When the interconnect
    * receives barrier from a master, then all other transactions launched by
    * other masters in that domain may be stalled. This cover point covers
    * condition where master issues transactions with non-zero QOS value. Then
    * another master issues a barrier transaction within the same domain.
    *
    * Two or more ACE/ACE_LITE masters needed for this covergroup
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; C 8.1 
    *
    */
  covergroup trans_master_ace_xacts_with_high_priority_from_other_master_during_barrier;
    ace_xacts_with_high_priority_from_other_master_during_barrier: coverpoint is_xacts_from_other_master_during_barrier_covered {
      bins xacts_from_other_master_during_barrier = {1};
    }
    option.per_instance = 1;
  endgroup
  
  /**
    * Covergroup: trans_master_ace_barrier_response_with_outstanding_xacts
    *
    * Coverpoints:
    * - ace_completed_barrier_type: This is covered when there are outstanding
    * transactions in the queue of a master when the response to a barrier is
    * received. There are multiple ways in which an interconnect can handle
    * barriers. Some interconnects may send response to a barrier only after
    * all outstanding transactions are complete. Others may forward
    * the barrier downstream and wait for the response of the downstream
    * barrier before responding to the original barrier. In such a case there
    * could be outstanding transactions in the queue of the master when a
    * barrier response is received. This coverpoint covers the latter behaviour.
    *
    * One or more ACE/ACE_LITE masters needed for this covergroup
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; C 8.3 
    */
  covergroup trans_master_ace_barrier_response_with_outstanding_xacts;
    ace_completed_barrier_type : 
    coverpoint completed_barrier_xact.barrier_type {
      bins outstanding_xacts_during_memory_barrier = {svt_axi_transaction::MEMORY_BARRIER};
      bins outstanding_xacts_during_sync_barrier = {svt_axi_transaction::SYNC_BARRIER};
      ignore_bins ignore_barrier_type = {svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER,svt_axi_transaction::NORMAL_ACCESS_IGNORE_BARRIER};
    }
    option.per_instance = 1;
  endgroup
  
  /**
    * Covergroup: trans_master_ace_store_overlapping_coherent_xact
    *
    * Coverpoints:
    *
    * - store_overlap_coh_xact:  This cover point has follwoing bins<br>
    *   overlap_readunique_readunique: This bin gets hit when two or more masters issue readunique coherent transactions to overlapping cacheline simultaneously.<br>
    *   overlap_cleanunique_cleanunique: This bin gets hit when two or more masters issue cleanunique coherent transactions to overlapping cacheline simultaneously.<br>
    *   overlap_makeunique_makeunique: This bin gets hit when two or more masters issue makeunique coherent transactions to overlapping cacheline simultaneously.<br>
    *
    * Two or more ACE masters needed for this covergroup
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C4.10
    *
    */
  covergroup trans_master_ace_store_overlapping_coherent_xact;
    ace_store_overlap_coh_xact: coverpoint store_overlap_coh_xact {
      bins overlap_readunique_readunique = {16'h05_05};
      bins overlap_cleanunique_cleanunique = {16'h06_06};
      bins overlap_makeunique_makeunique = {16'h07_07};
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_master_ace_no_cached_copy_overlapping_coherent_xact
    *
    * Coverpoints:
    *
    * - no_cached_copy_overlap_coh_xact:  This coverpoint has following bins<br>
    *   overlap_readonce_readonce: This bin gets hit when two or more masters issue readonce coherent transactions to overlapping cacheline simultaneously.<br>
    *   overlap_writeunique_writeunique: This bin gets hit when two or more masters issue writeunique coherent transactions to overlapping cacheline simultaneously.<br>
    *   overlap_writelineunique_writelineunique: This bin gets hit when two or more masters issue writelineunique coherent transactions to overlapping cacheline simultaneously.<br>
    *
    * Two or more ACE / ACE_LITE masters needed for this covergroup
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C1.3.4
    *
    */
  covergroup trans_master_ace_no_cached_copy_overlapping_coherent_xact;
    ace_no_cached_copy_overlap_coh_xact: coverpoint no_cached_copy_overlap_coh_xact {
      bins overlap_readonce_readonce = {16'h01_01};
      bins overlap_writeunique_writeunique = {16'h15_15};
      bins overlap_writelineunique_writelineunique = {16'h16_16};
    }
    option.per_instance = 1;
  endgroup

  /** 
  * Covergroup: trans_master_ace_lite_coherent_and_ace_snoop_response_association 
  *
  * Covergroup for all coherent transactions generated from ACE-Lite master and
  * the correponding Snoop response from ACE-Masters for these coherent transactions.
  * This will be a Port Level Covergroup and will be applicable for all
  * ACE-Masters and will only be created when there is atleast one ACE-Lite master
  * in the system. 
  *
  * Coverpoints: 
  * 
  * - coh_xact_from_ace_lite: This coverpoint has bins corresponding to each of the valid coherent
  * transactions from an ACE-Lite Master
  *
  * - snp_resp_from_ace: This coverpoint has bins for all possible values of CRRESP[3:0] (Snoop response)
  * that an ACE Master can send for each of the coherent transaction issued from ACE-Lite Master.
  * Since this CG is applicable for only ACE master, it is required to check whether any coherent 
  * transaction from ACE-Lite master resulted in this snoop response and subsequently hit bins of
  * coverpoint cmds_from_ace_lite. System Monitor provides this information to
  * Port Monitor.
  *  
  * - associate_snoop_xact_for_coh_xact_from_acelite_master: This coverpoint has bins corresponding to valid snoop transactions issued to ACE master for coherent xacts from ACE-Lite Master
  * - snoop_crresp_wu: This coverpoint has bins for all possible values of CRRESP[4] (WasUnique)
  *
  * - ace_init_cache_state: This coverpoint has bins for valid initial cache states corresponding to
  * snoops generated by ACE-Master.
  *
  * - ace_final_cache_state: This coverpoint has bins for valid final cache states corresponding to
  * snoops generated by ACE-Master.
  *
  * - coh_xact_ace_lite_snp_resp_ace_init_final_cache_state: This is the
  *   cross-coverage between coh_xact_from_ace_lite,associate_snoop_xact_for_coh_xact_from_acelite_master, snp_resp_from_ace, snoop_crresp_wu, ace_init_cache_state
  *   and ace_final_cache_state.
  * . 
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Table C6-1 
  * 
  */ 
  covergroup trans_master_ace_lite_coherent_and_ace_snoop_response_association; 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACELITE_COHERENT_XACT_TYPE 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACE_CRRESP
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WASUNIQUE_SNOOP_CRRESP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_INITIAL_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_FINAL_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACE_SNOOP_XACT_TYPE_FROM_ACELITE
    coh_xact_ace_lite_snp_resp_ace_init_final_cache_state : cross coh_xact_from_ace_lite, associate_snoop_xact_for_coh_xact_from_acelite_master,snoop_crresp_from_ace, snoop_crresp_wu, ace_init_cache_state, ace_final_cache_state {
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACELITE_SNOOP_ASSOCIATION_IGNORE_BINS
    }
    option.per_instance = 1; 
  endgroup

  /** 
  * Covergroup: trans_master_ace_lite_coherent_and_ace_snoop_response_association_specific_id
  *
  * Covergroup for all coherent transactions generated from ACE-Lite master and
  * the correponding Snoop response from ACE-Masters for these coherent transactions.
  * This will be sampled only when transaction is having configured specific id.
  * This will be a Port Level Covergroup and will be applicable for all
  * ACE-Masters and will only be created when there is atleast one ACE-Lite master
  * in the system. 
  *
  * Coverpoints: 
  * 
  * - coh_xact_from_ace_lite: This coverpoint has bins corresponding to each of the valid coherent
  * transactions from an ACE-Lite Master
  *
  * - snp_resp_from_ace: This coverpoint has bins for all possible values of CRRESP[3:0] (Snoop response)
  * that an ACE Master can send for each of the coherent transaction issued from ACE-Lite Master.
  * Since this CG is applicable for only ACE master, it is required to check whether any coherent 
  * transaction from ACE-Lite master resulted in this snoop response and subsequently hit bins of
  * coverpoint cmds_from_ace_lite. System Monitor provides this information to
  * Port Monitor.
  * 
  * - snoop_crresp_wu: This coverpoint has bins for all possible values of CRRESP[4] (WasUnique)
  *
  * - ace_init_cache_state: This coverpoint has bins for valid initial cache states corresponding to
  * snoops generated by ACE-Master.
  *
  * - ace_final_cache_state: This coverpoint has bins for valid final cache states corresponding to
  * snoops generated by ACE-Master.
  *
  * - coh_xact_ace_lite_snp_resp_ace_init_final_cache_state: This is the
  *   cross-coverage between coh_xact_from_ace_lite, snp_resp_from_ace, snoop_crresp_wu, ace_init_cache_state
  *   and ace_final_cache_state.
  * . 
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Table C6-1 
  * 
  */ 
  covergroup trans_master_ace_lite_coherent_and_ace_snoop_response_association_specific_id; 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACELITE_COHERENT_XACT_TYPE 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACE_CRRESP
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WASUNIQUE_SNOOP_CRRESP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_INITIAL_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_FINAL_STATE

    coh_xact_ace_lite_snp_resp_ace_init_final_cache_state : cross coh_xact_from_ace_lite, snoop_crresp_from_ace, snoop_crresp_wu, ace_init_cache_state, ace_final_cache_state {
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_ASSOCIATION_IGNORE_BINS
    }
    option.per_instance = 1; 
  endgroup

  /** 
  * Covergroup: trans_master_ace_lite_coherent_and_ace_snoop_response_association_back_to_back_xact_with_specific_id 
  *
  * Covergroup for back to back combination of CLEANINVALID and MAKEINVALID coherent 
  * transactions generated from ACE-Lite master and
  * the correponding Snoop response from ACE-Masters for these coherent transactions.
  * This will be a Port Level Covergroup and will be applicable for all
  * ACE-Masters and will only be created when there is atleast one ACE-Lite master
  * in the system. 
  *
  * Coverpoints: 
  * 
  * - coh_xact_t1_ace_lite: This coverpoint has bins corresponding to first
  *   transaction of a back to back transactions from an ACE-Lite Master
  * - coh_xact_t2_ace_lite: This coverpoint has bins corresponding to second
  *   transaction of a back to back transactions from an ACE-Lite Master
  *
  * - snoop_crresp_0_t1 & snoop_crresp_0_t2: This coverpoint has bins for all 
  * possible values of CRRESP[0] (Snoop response) that an ACE Master can send for each of the 
  * coherent transaction issued from ACE-Lite Master.
  * 
  * - coh_xact_ace_lite_xacts_ace_snp_resp_specific_id: This is the
  *   cross-coverage between coh_xact_t1_ace_lite, snoop_crresp_0_t1, coh_xact_t2_ace_lite, snoop_crresp_0_t2, coh_xact_id.
  * .
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Table C6-1 
  * 
  */ 
  covergroup trans_master_ace_lite_coherent_and_ace_snoop_response_association_back_to_back_xact_with_specific_id(int specific_id); 
    
    coh_xact_t1_ace_lite: coverpoint ace_lite_coh_xact_t1_type {
      bins writeunique_coherent = {svt_axi_transaction::WRITEUNIQUE}; 
      bins writelineunique_coherent = {svt_axi_transaction::WRITELINEUNIQUE}; 
      option.weight = 1;
    }

    coh_xact_t2_ace_lite: coverpoint ace_lite_coh_xact_t2_type {
      bins writeunique_coherent = {svt_axi_transaction::WRITEUNIQUE}; 
      bins writelineunique_coherent = {svt_axi_transaction::WRITELINEUNIQUE}; 
      option.weight = 1;
    }

    snoop_crresp_0_t1: coverpoint snoop_resp_t1_from_ace_master[0] {
      bins cresp_0 = {1'b0};
      bins cresp_1 = {1'b1};
      option.weight = 1;
    }

    snoop_crresp_0_t2: coverpoint snoop_resp_t2_from_ace_master[0] {
      bins cresp_0 = {1'b0};
      bins cresp_1 = {1'b1};
      option.weight = 1;
    }

    coh_xact_id : coverpoint ace_lite_coh_xact_id {
      bins ace_lite_xact_id[] = {specific_id};
      option.weight = 1;
    }

    coh_xact_ace_lite_xacts_ace_snp_resp_specific_id : cross coh_xact_t1_ace_lite, snoop_crresp_0_t1, coh_xact_t2_ace_lite, snoop_crresp_0_t2, coh_xact_id {
      option.weight = 1;
    }
    option.per_instance = 1; 
  endgroup
/** 
  * Covergroup: trans_master_ace_coherent_and_ace_snoop_response_association 
  *
  * Covergroup for all coherent transactions generated from ACE master and
  * the correponding Snoop transactions on ACE-Masters and snoop response from ACE-Masters for these snoop transactions.
  * This will be a Port Level Covergroup and will be applicable for all
  * ACE-Masters and will only be created when there are two ACE masters 
  * in the system. 
  *
  * Coverpoints: 
  * 
  * - coh_xact_from_ace: This coverpoint has bins corresponding to each of the valid coherent
  * transactions from an ACE Master
  *
  * - snp_resp_from_ace: This coverpoint has bins for all possible values of CRRESP[3:0] (Snoop response)
  * that an ACE Master can send for each of the coherent transaction issued from ACE Master.
  * Since this CG is applicable for only ACE master, it is required to check whether any coherent 
  * transaction from ACE master resulted in this snoop transaction and snoop response and subsequently hit bins of
  * coverpoint cmds_from_ace. System Monitor provides this information to
  * Port Monitor.
  *  
  * - snoop_xact_on_ace_master: This coverpoint has bins corresponding to each of the valid snoop transaction type
  *  on ACE master 
  * - snoop_crresp_wu: This coverpoint has bins for all possible values of CRRESP[4] (WasUnique)
  *
  * - ace_init_cache_state: This coverpoint has bins for valid initial cache states corresponding to
  * snoops generated by ACE-Master.
  *
  * - ace_final_cache_state: This coverpoint has bins for valid final cache states corresponding to
  * snoops generated by ACE-Master.
  *
  * - coh_xact_ace_snp_resp_ace_init_final_cache_state: This is the
  *   cross-coverage between coh_xact_from_ace, snoop_xact_on_ace_master,snp_crresp_from_ace, snoop_crresp_wu, ace_init_cache_state
  *   and ace_final_cache_state.
  * . 
  * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Table C6-1 
  * 
  */ 
  covergroup trans_master_ace_coherent_and_ace_snoop_response_association; 
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACE_COHERENT_XACT_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACE_CRRESP
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_WASUNIQUE_SNOOP_CRRESP_TYPE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_INITIAL_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_SNOOP_FINAL_STATE
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACE_SNOOP_XACT_TYPE_FROM_ACE
    coh_xact_ace_snp_resp_ace_init_final_cache_state : cross coh_xact_from_ace, snoop_xact_on_ace_master,snoop_crresp_from_ace, snoop_crresp_wu, ace_init_cache_state, ace_final_cache_state {
    `SVT_AXI_PORT_MONITOR_DEF_COV_UTIL_ACE_SNOOP_ASSOCIATION_IGNORE_BINS
    }
    option.per_instance = 1; 
  endgroup

  /** 
    * Covergroup: system_ace_coherent_and_snoop_association_recommended_and_optional_ace 
    * 
    * Coverpoints: 
    * 
    * - ace_coh_and_snp_association:  This is covered when the interconnect issues recommended 
    *   and optional snoop transaction to the snooped masters, in response to the coherent  
    *   transaction received from the initiating master.  
    * . 
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Table C6-1 
    * 
    */ 
  //covergroup trans_master_ace_coherent_and_snoop_association_recommended_and_optional @(cov_sys_coh_and_snp_association_sample_event); 
  covergroup trans_master_ace_coherent_and_snoop_association_recommended_and_optional_ace;
    ace_coh_and_snp_association: coverpoint coh_and_snp_association { 
      bins readonce_coherent_to_readonce_snoop = {16'h01_00}; 
      bins readonce_coherent_to_readclean_snoop = {16'h01_02};  
      bins readonce_coherent_to_readnotshareddirty_snoop = {16'h01_03}; 
      bins readonce_coherent_to_readshared_snoop = {16'h01_01}; 
      bins readonce_coherent_to_readunique_snoop = {16'h01_07}; 
      bins readonce_coherent_to_cleaninvalid_snoop = {16'h01_09}; 
      bins readonce_coherent_to_cleanshared_snoop = {16'h01_08}; 
       
      bins readclean_coherent_to_readclean_snoop = {16'h03_02};  

      bins readclean_coherent_to_readnotshareddirty_snoop = {16'h03_03}; 
      bins readclean_coherent_to_readshared_snoop = {16'h03_01}; 
      bins readclean_coherent_to_readunique_snoop = {16'h03_07}; 
      bins readclean_coherent_to_cleaninvalid_snoop = {16'h03_09}; 
  
      bins readnotshareddirty_coherent_to_readclean_snoop = {16'h04_02}; 
      bins readnotshareddirty_coherent_to_readnotshareddirty_snoop = {16'h04_03}; 
      bins readnotshareddirty_coherent_to_readshared_snoop = {16'h04_01}; 
      bins readnotshareddirty_coherent_to_readunique_snoop = {16'h04_07}; 
      bins readnotshareddirty_coherent_to_cleaninvalid_snoop = {16'h04_09}; 
  
      bins readshared_coherent_to_readclean_snoop = {16'h02_02};  
      bins readshared_coherent_to_readnotshareddirty_snoop = {16'h02_03}; 
      bins readshared_coherent_to_readshared_snoop = {16'h02_01}; 
      bins readshared_coherent_to_readunique_snoop = {16'h02_07}; 
      bins readshared_coherent_to_cleaninvalid_snoop = {16'h02_09}; 
  
      bins readunique_coherent_to_readunique_snoop = {16'h05_07}; 
      bins readunique_coherent_to_cleaninvalid_snoop = {16'h05_09}; 
  
      bins cleanunique_coherent_to_readunique_snoop = {16'h06_07}; 
      bins cleanunique_coherent_to_cleaninvalid_snoop = {16'h06_09}; 
  
      bins makeunique_coherent_to_readunique_snoop = {16'h07_07}; 
      bins makeunique_coherent_to_cleaninvalid_snoop = {16'h07_09}; 

      bins makeunique_coherent_to_makeinvalid_snoop = {16'h07_0d}; 
  
      bins cleanshared_coherent_to_readunique_snoop = {16'h08_07}; 
      bins cleanshared_coherent_to_cleaninvalid_snoop = {16'h08_09}; 
      bins cleanshared_coherent_to_cleanshared_snoop = {16'h08_08}; 
`ifdef SVT_ACE5_ENABLE
      bins cleansharedpersist_coherent_to_readunique_snoop = {16'h10_07}; 
      bins cleansharedpersist_coherent_to_cleaninvalid_snoop = {16'h10_09}; 
      bins cleansharedpersist_coherent_to_cleanshared_snoop = {16'h10_08}; 
`endif
      bins cleaninvalid_coherent_to_readunique_snoop = {16'h09_07}; 
      bins cleaninvalid_coherent_to_cleaninvalid_snoop = {16'h09_09}; 
  
      bins makeinvalid_coherent_to_readunique_snoop = {16'h0a_07}; 
      bins makeinvalid_coherent_to_cleaninvalid_snoop = {16'h0a_09}; 
      bins makeinvalid_coherent_to_makeinvalid_snoop = {16'h0a_0d}; 
  
      bins writeunique_coherent_to_readunique_snoop = {16'h0f_07}; 
      bins writeunique_coherent_to_cleaninvalid_snoop = {16'h0f_09}; 
  
      bins writelineunique_coherent_to_readunique_snoop = {16'h10_07}; 
      bins writelineunique_coherent_to_cleaninvalid_snoop = {16'h10_09}; 
      bins writelineunique_coherent_to_makeinvalid_snoop = {16'h10_0d}; 
    } 
    option.per_instance = 1; 
  endgroup 

  /** 
    * Covergroup: system_ace_coherent_and_snoop_association_recommended_and_optional_ace_lite 
    * 
    * Coverpoints: 
    * 
    * - ace_coh_and_snp_association:  This is covered when the interconnect issues recommended 
    *   and optional snoop transaction to the snooped masters, in response to the coherent  
    *   transaction received from the initiating master.  
    * . 
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Table C6-1 
    * 
    */ 
  //covergroup trans_master_ace_coherent_and_snoop_association_recommended_and_optional @(cov_sys_coh_and_snp_association_sample_event); 
  covergroup trans_master_ace_coherent_and_snoop_association_recommended_and_optional_ace_lite;
    ace_coh_and_snp_association: coverpoint coh_and_snp_association { 
      bins readonce_coherent_to_readonce_snoop = {16'h01_00}; 
      bins readonce_coherent_to_readclean_snoop = {16'h01_02};  
      bins readonce_coherent_to_readnotshareddirty_snoop = {16'h01_03}; 
      bins readonce_coherent_to_readshared_snoop = {16'h01_01}; 
      bins readonce_coherent_to_readunique_snoop = {16'h01_07}; 
      bins readonce_coherent_to_cleaninvalid_snoop = {16'h01_09}; 
      bins readonce_coherent_to_cleanshared_snoop = {16'h01_08}; 
       
      bins cleanshared_coherent_to_readunique_snoop = {16'h08_07}; 
      bins cleanshared_coherent_to_cleaninvalid_snoop = {16'h08_09}; 
      bins cleanshared_coherent_to_cleanshared_snoop = {16'h08_08}; 
`ifdef SVT_ACE5_ENABLE
      bins cleansharedpersist_coherent_to_readunique_snoop = {16'h10_07}; 
      bins cleansharedpersist_coherent_to_cleaninvalid_snoop = {16'h10_09}; 
      bins cleansharedpersist_coherent_to_cleanshared_snoop = {16'h10_08}; 
`endif
      bins cleaninvalid_coherent_to_readunique_snoop = {16'h09_07}; 
      bins cleaninvalid_coherent_to_cleaninvalid_snoop = {16'h09_09}; 
  
      bins makeinvalid_coherent_to_readunique_snoop = {16'h0a_07}; 
      bins makeinvalid_coherent_to_cleaninvalid_snoop = {16'h0a_09}; 
      bins makeinvalid_coherent_to_makeinvalid_snoop = {16'h0a_0d}; 
  
      bins writeunique_coherent_to_readunique_snoop = {16'h0f_07}; 
      bins writeunique_coherent_to_cleaninvalid_snoop = {16'h0f_09}; 
  
      bins writelineunique_coherent_to_readunique_snoop = {16'h10_07}; 
      bins writelineunique_coherent_to_cleaninvalid_snoop = {16'h10_09}; 
      bins writelineunique_coherent_to_makeinvalid_snoop = {16'h10_0d}; 

    } 
    option.per_instance = 1; 
  endgroup 

  /**
    * Covergroup: trans_axi_num_outstanding_xacts_with_same_arid<br>
    * Coverpoints: <br>
    * - read_outstanding_xacts_with_same_arid: Captures the number of
    *   outstanding read transactions with a matching ARID value to the one
    *   programmed in
    *   svt_axi_port_configuration::cov_same_id_in_outstanding_xacts.
    *   
    *   The number of bins for this coverpoint is controlled by
    *   svt_axi_port_configuration::cov_bins_num_outstanding_xacts, the
    *   default value of which is 64.
    *   Configured value of svt_axi_port_configuration::cov_bins_num_outstanding_xacts
    *   should be less than or equal to configured value of 
    *   svt_axi_port_configuration::num_outstanding_xact or 
    *   svt_axi_port_configuration::num_write_outstanding_xact if 
    *   svt_axi_port_configuration::num_outstanding_xact is set to -1 which
    *   indicates the number of outstanding transactions VIP can support.
    *   
    *   Example:
    *   If outstanding transactions have the following IDs: ARID1 ARID1 ARID3 ARID1 ARID3 ARID2
    *   and svt_axi_port_configuration::cov_same_id_in_outstanding_xacts is
    *   programmed to ARID1.
    *   The bins hit will be 1,2 and 3 as there are 3 outstanding transactions
    *   matching with ARID1. 
    *   
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A5.2
    */
  covergroup trans_axi_num_outstanding_xacts_with_same_arid (int num_outstanding_xact);
    read_outstanding_xacts_with_same_arid: coverpoint read_outstanding_xacts_with_same_arid{
      bins read_outstanding_xacts_with_same_arid[] = {[1:num_outstanding_xact]} ;
    }
    option.per_instance = 1;
  endgroup
  
  /**
    * Covergroup: trans_axi_num_outstanding_xacts_with_multiple_same_arid<br>
    *  This covergroup captures the number of outstanding read transactions
    *  with same ARID values which is in progress, if master is programmed
    *  with multiple same ids. For Example : If a master is programmed with
    *  svt_axi_port_configuration::cov_multi_same_ids = new[3], then the
    *  master will have three different ids ARID1, ARID2 and ARID3.This
    *  covergroup will cross all the 3 ids with
    *  svt_axi_port_configuration::num_outstanding_xact. If number of
    *  outstanding transactions are 50 with ARID1,then bins read_same_arid_1,
    *  read_outstanding_xacts_with_same_arid_1 to read_outstanding_xacts_with_same_arid_50 will get hit.
    * Coverpoints: <br>
    * - read_outstanding_same_id: Captures the same id values programmed in svt_axi_port_configuration::cov_multi_same_ids
    * - num_outstanding_read : Captures number of outstanding read
    *   transactions with a matching ARID values to the one
    *   programmed in svt_axi_port_configuration::cov_multi_same_ids.
    *   
    *   The number of bins for this coverpoint is controlled by
    *   svt_axi_port_configuration::cov_bins_num_outstanding_xacts, the
    *   default value of which is 64.
    *   Configured value of svt_axi_port_configuration::cov_bins_num_outstanding_xacts
    *   should be less than or equal to configured value of 
    *   svt_axi_port_configuration::num_outstanding_xact or 
    *   svt_axi_port_configuration::num_write_outstanding_xact if 
    *   svt_axi_port_configuration::num_outstanding_xact is set to -1 which
    *   indicates the number of outstanding transactions VIP can support.
    *   
    *   Example:
    *   If a master is programmed with svt_axi_port_configuration::cov_multi_same_ids = new[3],
    *   cov_multi_same_ids[0] = ARID1, cov_multi_same_ids[1] = ARID2,
    *   cov_multi_same_ids[1] = ARID3 and outstanding transactions have the
    *   following IDs: ARID1 ARID2 ARID1 ARID4 ARID3 ARID1 ARID3 ARID5 ARID2.
    *   The bins of read_outstanding_same_id hit will be read_same_arid_1,read_same_arid_2 and
    *   read_same_arid_3, bins of cross_same_id_with_num_outstanding_xacts hit will
    *   be read_same_arid_1 with read_outstanding_xacts_3,read_same_arid_2
    *   with read_outstanding_xacts_2, read_same_arid_3 with
    *   read_outstanding_xacts_1 as there are 3 outstanding transactions
    *   matching with ARID1, 2 outstanding transactions with ARID2 and 1
    *   outstanding transaction with ARID3. 
    *   
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A5.2
    */
  covergroup trans_axi_num_outstanding_xacts_with_multiple_same_arid (int num_same_ids, int num_outstanding_xact);
    
    read_outstanding_same_id : coverpoint cov_read_same_id {
      bins read_same_arid[] = {[1:num_same_ids]};
      option.weight = 1;
    }
    num_outstanding_read : coverpoint cov_num_read_outstanding_same_arid{
      bins read_outstanding_xacts[] = {[1:num_outstanding_xact]};
      option.weight = 1;
    }
    
    cross_same_id_with_num_outstanding_xacts : cross read_outstanding_same_id, num_outstanding_read { 
     option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_axi_num_outstanding_xacts_with_diff_arid<br>
    * Coverpoints: <br>
    * - read_outstanding_xacts_with_diff_arid: Captures the number of
    *   outstanding read transactions with different ARID value.
    *   The number of bins will be equal to the programmed value of User-defined macro
    *   SVT_AXI_NUM_BINS_FOR_ID_WIDTH_GREATER_THAN_EIGHT which has a default value of 256. 
    *   So, if user does not override this macro then this covergroup will create 256 bins for ARID width greater than 8

    *   If svt_axi_port_configuration::use_separate_rd_wr_chan_id_width is 
    *   programmed to 1 then svt_axi_port_configuration::read_chan_id_width is
    *   considered for creation of bins. 
    *   If svt_axi_port_configuration::use_separate_rd_wr_chan_id_width is 
    *   programmed to 0 then svt_axi_port_configuration::id_width is
    *   considered for creation of bins. 
    *   
    *   Example:
    *   If outstanding transactions have the following IDs: ARID1 ARID1 ARID2
    *   ARID3 ARID4 ARID5.
    *   The bins hit will be 1,2,3,4,5 (for outstanding transactions with ARID1,ARID2
    *   ARID3 ARID4 ARID5)
    *   The coverage is a continuous logic. If there is only one outstanding 
    *   transaction in the queue with unique ARID value, the bin 1 will get hit.
    *   Subsequently as and when new outstanding transactions comes with unique
    *   ARID values further bins will keep getting hit.
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A5.2
    */
  covergroup trans_axi_num_outstanding_xacts_with_diff_arid (int num_outstanding_xact);
    read_outstanding_xacts_with_diff_arid: coverpoint read_outstanding_xacts_with_diff_arid{
      bins read_outstanding_xacts_with_diff_arid[] = {[1:num_outstanding_xact]} ;
    }
    option.per_instance = 1;
  endgroup
/**
    * Covergroup: trans_axi_num_outstanding_xacts_with_diff_arid_range<br>
    * Coverpoints: <br>
    * - read_outstanding_xacts_with_diff_arid: Captures the number of
    *   outstanding read transactions with different ARID value.
    *   The number of bins will be equal to the programmed value of User-defined macro
    *  SVT_AXI_NUM_BINS_FOR_ID_WIDTH_GREATER_THAN_EIGHT which has a default value of 256. 
    *   So, if user does not override this macro then this covergroup will create 256 bins for ARID width greater than 8

    *   If svt_axi_port_configuration::use_separate_rd_wr_chan_id_width is 
    *   programmed to 1 then svt_axi_port_configuration::read_chan_id_width is
    *   considered for creation of bins. 
    *   If svt_axi_port_configuration::use_separate_rd_wr_chan_id_width is 
    *   programmed to 0 then svt_axi_port_configuration::id_width is
    *   considered for creation of bins. 
    *   
    *   Example:
    *   If outstanding transactions have the following IDs: ARID1 ARID1 ARID2
    *   ARID3 ARID4 ARID5.
    *   The bins hit will be 1,2,3,4,5 (for outstanding transactions with ARID1,ARID2
    *   ARID3 ARID4 ARID5)
    *   The coverage is a continuous logic. If there is only one outstanding 
    *   transaction in the queue with unique ARID value, the bin 1 will get hit.
    *   Subsequently as and when new outstanding transactions comes with unique
    *   ARID values further bins will keep getting hit.
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A5.2
    */
  covergroup trans_axi_num_outstanding_xacts_with_diff_arid_range (int num_outstanding_xact);
    read_outstanding_xacts_with_diff_arid: coverpoint read_outstanding_xacts_with_diff_arid{
      bins read_outstanding_xacts_with_diff_arid_range_0 = {[1:num_outstanding_xact]};
      bins read_outstanding_xacts_with_diff_arid_range_1 = {[(num_outstanding_xact+1):(2*num_outstanding_xact)]};   
      bins read_outstanding_xacts_with_diff_arid_range_2 = {[(2*num_outstanding_xact+1):(3*num_outstanding_xact)]};
      bins read_outstanding_xacts_with_diff_arid_range_3 = {[(3*num_outstanding_xact+1):(4*num_outstanding_xact)]};
      bins read_outstanding_xacts_with_diff_arid_range_4 = {[(4*num_outstanding_xact+1):(5*num_outstanding_xact)]};
      bins read_outstanding_xacts_with_diff_arid_range_5 = {[(5*num_outstanding_xact+1):(6*num_outstanding_xact)]};
      bins read_outstanding_xacts_with_diff_arid_range_6 = {[(6*num_outstanding_xact+1):(7*num_outstanding_xact)]};
      bins read_outstanding_xacts_with_diff_arid_range_7 = {[(7*num_outstanding_xact+1):(8*num_outstanding_xact)]};
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_axi_num_outstanding_xacts_with_same_awid<br>
    * Coverpoints: <br>
    * - write_outstanding_xacts_with_same_awid: Captures the number of
    *   outstanding write transactions with a matching AWID value to the one
    *   programmed in
    *   svt_axi_port_configuration::cov_same_id_in_outstanding_xacts.
    *   
    *   The number of bins for this coverpoint is controlled by
    *   svt_axi_port_configuration::cov_bins_num_outstanding_xacts, the
    *   default value of which is 64.
    *   Configured value of svt_axi_port_configuration::cov_bins_num_outstanding_xacts
    *   should be less than or equal to configured value of 
    *   svt_axi_port_configuration::num_outstanding_xact or 
    *   svt_axi_port_configuration::num_write_outstanding_xact if 
    *   svt_axi_port_configuration::num_outstanding_xact is set to -1 which
    *   indicates the number of outstanding transactions VIP can support.
    *   
    *   Example:
    *   If outstanding transactions have the following IDs: AWID1 AWID1 AWID3 AWID1 AWID3  
    *   AWID2 and svt_axi_port_configuration::cov_same_id_in_outstanding_xacts is
    *   programmed to AWID1.
    *   The bins hit will be 1, 2 and 3 as there are 3 outstanding transactions
    *   matching with AWID1. 
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A5.2
    */
  covergroup trans_axi_num_outstanding_xacts_with_same_awid (int num_outstanding_xact);
    write_outstanding_xacts_with_same_awid: coverpoint write_outstanding_xacts_with_same_awid{
      bins write_outstanding_xacts_with_same_awid[] = {[1:num_outstanding_xact]} ;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_axi_num_outstanding_xacts_with_multiple_same_awid<br>
    *  This covergroup captures the number of outstanding write transactions
    *  with same AWID values which is in progress, if master is programmed
    *  with multiple same ids. For Example : If a master is programmed with
    *  svt_axi_port_configuration::cov_multi_same_ids = new[3], then the
    *  master will have three different ids AWID1, AWID2 and AWID3.This
    *  covergroup will cross all the 3 ids with
    *  svt_axi_port_configuration::num_outstanding_xact. If number of
    *  outstanding transactions are 50 with AWID1,then bins write_same_awid_1,
    *  write_outstanding_xacts_with_same_awid_1 to write_outstanding_xacts_with_same_awid_50 will get hit.
    * Coverpoints: <br>
    * - write_outstanding_same_id: Captures the same id values programmed in svt_axi_port_configuration::cov_multi_same_ids
    * - num_outstanding_write : Captures number of outstanding write
    *   transactions with a matching AWID values to the one
    *   programmed in svt_axi_port_configuration::cov_multi_same_ids.
    *   
    *   The number of bins for this coverpoint is controlled by
    *   svt_axi_port_configuration::cov_bins_num_outstanding_xacts, the
    *   default value of which is 64.
    *   Configured value of svt_axi_port_configuration::cov_bins_num_outstanding_xacts
    *   should be less than or equal to configured value of 
    *   svt_axi_port_configuration::num_outstanding_xact or 
    *   svt_axi_port_configuration::num_write_outstanding_xact if 
    *   svt_axi_port_configuration::num_outstanding_xact is set to -1 which
    *   indicates the number of outstanding transactions VIP can support.
    *   
    *   Example:
    *   If a master is programmed with svt_axi_port_configuration::cov_multi_same_ids = new[3],
    *   cov_multi_same_ids[0] = AWID1, cov_multi_same_ids[1] = AWID2,
    *   cov_multi_same_ids[1] = AWID3 and outstanding transactions have the
    *   following IDs: AWID1 AWID2 AWID1 AWID4 AWID3 AWID1 AWID3 AWID5 AWID2.
    *   The bins of write_outstanding_same_id hit will be write_same_awid_1,write_same_awid_2 and
    *   write_same_awid_3, bins of cross_same_id_with_num_outstanding_xacts hit will
    *   be write_same_awid_1 with write_outstanding_xacts_3,write_same_awid_2
    *   with write_outstanding_xacts_2, write_same_awid_3 with
    *   write_outstanding_xacts_1 as there are 3 outstanding transactions
    *   matching with AWID1, 2 outstanding transactions with AWID2 and 1
    *   outstanding transaction with AWID3. 
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A5.2
    */
  covergroup trans_axi_num_outstanding_xacts_with_multiple_same_awid (int num_same_ids, int num_outstanding_xact);
    
    write_outstanding_same_id : coverpoint cov_write_same_id {
      bins write_same_awid[] = {[1:num_same_ids]};
      option.weight = 1;
    }
    num_outstanding_write : coverpoint cov_num_write_outstanding_same_awid{
      bins write_outstanding_xacts[] = {[1:num_outstanding_xact]};
      option.weight = 1;
    }
    
    cross_same_id_with_num_outstanding_xacts : cross write_outstanding_same_id, num_outstanding_write { 
     option.weight = 1;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_axi_num_outstanding_xacts_with_diff_awid<br>
    * Coverpoints: <br>
    * - write_outstanding_xacts_with_diff_awid: Captures the number of
    *   outstanding write transactions with different AWID.
    *   The number of bins will be equal to the programmed value of User-defined macro 
    *   SVT_AXI_NUM_BINS_FOR_ID_WIDTH_GREATER_THAN_EIGHT which has a default value of 256. 
    *   So, if user does not override this macro then this covergroup will create 256 bins for AWID width greater than 8

    *   If svt_axi_port_configuration::use_separate_rd_wr_chan_id_width is 
    *   programmed to 1 then svt_axi_port_configuration::write_chan_id_width is
    *   considered for creation of bins. 
    *   If svt_axi_port_configuration::use_separate_rd_wr_chan_id_width is 
    *   programmed to 0 then svt_axi_port_configuration::id_width is
    *   considered for creation of bins. 
    *
    *   Example:
    *
    *   If outstanding transactions have the following IDs: AWID1 AWID1 AWID2
    *   AWID3 AWID4 AWID5.
    *   The bins hit will be 1,2,3,4,5 (for outstanding transactions with AWID1,AWID2
    *   AWID3 AWID4 AWID5) 
    *   The coverage is a continuous logic. If there is only one outstanding 
    *   transaction in the queue with unique AWID value, the bin 1 will get hit.
    *   Subsequently as and when new outstanding transactions comes with unique
    *   AWID values further bins will keep getting hit.
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A5.2
    */
  covergroup trans_axi_num_outstanding_xacts_with_diff_awid (int num_outstanding_xact);
    write_outstanding_xacts_with_diff_awid: coverpoint write_outstanding_xacts_with_diff_awid{
      bins write_outstanding_xacts_with_diff_awid[] = {[1:num_outstanding_xact]} ;
    }
    option.per_instance = 1;
  endgroup

 /**
    * Covergroup: trans_axi_num_outstanding_xacts_with_diff_awid_range<br>
    * Coverpoints: <br>
    * - write_outstanding_xacts_with_diff_awid: Captures the number of
    *   outstanding write transactions with different AWID.
    *   The number of bins will be equal to the programmed value of User-defined macro 
    *   SVT_AXI_NUM_BINS_FOR_ID_WIDTH_GREATER_THAN_EIGHT which has a default value of 256. 
    *   So, if user does not override this macro then this covergroup will create 256 bins for AWID width greater than 8

    *   If svt_axi_port_configuration::use_separate_rd_wr_chan_id_width is 
    *   programmed to 1 then svt_axi_port_configuration::write_chan_id_width is
    *   considered for creation of bins. 
    *   If svt_axi_port_configuration::use_separate_rd_wr_chan_id_width is 
    *   programmed to 0 then svt_axi_port_configuration::id_width is
    *   considered for creation of bins. 
    *
    *   Example:
    *
    *   If outstanding transactions have the following IDs: AWID1 AWID1 AWID2
    *   AWID3 AWID4 AWID5.
    *   The bins hit will be 1,2,3,4,5 (for outstanding transactions with AWID1,AWID2
    *   AWID3 AWID4 AWID5) 
    *   The coverage is a continuous logic. If there is only one outstanding 
    *   transaction in the queue with unique AWID value, the bin 1 will get hit.
    *   Subsequently as and when new outstanding transactions comes with unique
    *   AWID values further bins will keep getting hit.
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section A5.2
    */
  covergroup trans_axi_num_outstanding_xacts_with_diff_awid_range (int num_outstanding_xact);
    write_outstanding_xacts_with_diff_awid: coverpoint write_outstanding_xacts_with_diff_awid{
      bins write_outstanding_xacts_with_diff_awid_range_0 = {[1:num_outstanding_xact]};
      bins write_outstanding_xacts_with_diff_awid_range_1 = {[(num_outstanding_xact+1):(2*num_outstanding_xact)]};   
      bins write_outstanding_xacts_with_diff_awid_range_2 = {[(2*num_outstanding_xact+1):(3*num_outstanding_xact)]};
      bins write_outstanding_xacts_with_diff_awid_range_3 = {[(3*num_outstanding_xact+1):(4*num_outstanding_xact)]};
      bins write_outstanding_xacts_with_diff_awid_range_4 = {[(4*num_outstanding_xact+1):(5*num_outstanding_xact)]};
      bins write_outstanding_xacts_with_diff_awid_range_5 = {[(5*num_outstanding_xact+1):(6*num_outstanding_xact)]};
      bins write_outstanding_xacts_with_diff_awid_range_6 = {[(6*num_outstanding_xact+1):(7*num_outstanding_xact)]};
      bins write_outstanding_xacts_with_diff_awid_range_7 = {[(7*num_outstanding_xact+1):(8*num_outstanding_xact)]};
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_ace_num_outstanding_snoop_xacts<br>
    * Coverpoints: <br>
    * -num_outstanding_snoop_xacts: Captures the number of outstanding snoop 
    *  transactions.The number of bins for this coverpoint is controlled by
    *  svt_axi_port_configuration::cov_bins_num_outstanding_snoop_xacts, the
    *  default value of which is 64. 
    *  Configured value of svt_axi_port_configuration::cov_bins_num_outstanding_snoop_xacts
    *  should be less than or equal to configured value of   
    *  svt_axi_port_configuration::num_outstanding_snoop_xact which
    *  indicates the number of outstanding snoop transactions VIP can support.
    *   
    *  Applicable only for master and when svt_axi_port_configuration::axi_interface_type is ACE.
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C5 
    */
  covergroup trans_ace_num_outstanding_snoop_xacts (int num_outstanding_xact);
    num_outstanding_snoop_xacts: coverpoint num_outstanding_snoop_xacts{
      bins num_outstanding_snoop_xacts[] = {[1:num_outstanding_xact]} ;
    }
    option.per_instance = 1;
  endgroup  

  /**
    * Covergroup:
      * trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid<br>
    * Coverpoints: <br>
    * - num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid: Captures the number
    *   of outstanding transactions with DVM TLBI requests with a matching ARID value
    *   to the one programmed in
    *   svt_axi_port_configuration::cov_same_id_in_dvm_tlbi_outstanding_xacts.
    *   
    *   The number of bins for this coverpoint is controlled by
    *   svt_axi_port_configuration::cov_bins_dvm_tlbi_num_outstanding_xacts, the
    *   default value of which is 64.
    *   Configured value of svt_axi_port_configuration::cov_bins_dvm_tlbi_num_outstanding_xacts
    *   should be less than or equal to configured value of 
    *   svt_axi_port_configuration::num_outstanding_xact or 
    *   svt_axi_port_configuration::num_read_outstanding_xact if 
    *   svt_axi_port_configuration::num_outstanding_xact is set to -1 which
    *   indicates the number of outstanding transactions VIP can support.
    *   
    *   Example:
    *   If outstanding DVM TLBI transactions have the following IDs: ARID1 ARID1 ARID3 ARID1 ARID3 ARID2
    *   and svt_axi_port_configuration::cov_same_id_in_dvm_tlbi_outstanding_xacts is
    *   programmed to ARID1.
    *   The bins hit will be 1,2 and 3 as there are 3 outstanding DVM TLBI transactions
    *   matching with ARID1.  
    *
    * Applicable only when svt_axi_port_configuration::axi_interface_type is ACE or ACE_LITE.
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C5 
    */
  covergroup trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid(int num_outstanding_xact);
    num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid: coverpoint num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid{
      bins num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid[] = {[1:num_outstanding_xact]} ;
    }
    option.per_instance = 1;
  endgroup

  /**
    * Covergroup: trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid<br>
    * Coverpoints: <br>
    * - num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid: Captures the number of outstanding 
    *   transactions with DVM TLBI requests with different ARID.
    *   The number of bins will be equal to the programmed value of User-defined macro
    *   SVT_AXI_NUM_BINS_FOR_ID_WIDTH_GREATER_THAN_EIGHT which has a default value of 256. 
    *   So, if user does not override this macro then this covergroup will create 256 bins for ARID width greater than 8

    *   If svt_axi_port_configuration::use_separate_rd_wr_chan_id_width is 
    *   programmed to 1 then svt_axi_port_configuration::read_chan_id_width is
    *   considered for creation of bins. 
    *   If svt_axi_port_configuration::use_separate_rd_wr_chan_id_width is 
    *   programmed to 0 then svt_axi_port_configuration::id_width is
    *   considered for creation of bins.
    *
    *   Example:
    *   If outstanding DVM TLBI transactions have the following IDs:
    *   ARID1 ARID1 ARID2 ARID3 ARID4 ARID5.
    *   The bins hit will be 1,2,3,4,5 (for outstanding transactions with ARID1,ARID2
    *   ARID3 ARID4 ARID5)
    *   The coverage is a continuous logic. If there is only one outstanding 
    *   transaction in the queue with unique ARID value, the bin 1 will get hit.
    *   Subsequently as and when new outstanding transactions comes with unique
    *   ARID values further bins will keep getting hit.
    *
    * Applicable only when svt_axi_port_configuration::axi_interface_type is ACE or ACE_LITE.
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C5 
    */
  covergroup trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid(int num_outstanding_xact);
    num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid: coverpoint num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid{
      bins num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid[] = {[1:num_outstanding_xact]} ;
       
    }
    option.per_instance = 1;
  endgroup  

  /**
    * Covergroup: trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range<br>
    * Coverpoints: <br>
    * - num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid: Captures the number of outstanding 
    *   transactions with DVM TLBI requests with different ARID.
    *   The number of bins will be equal to the programmed value of User-defined macro
    *   SVT_AXI_NUM_BINS_FOR_ID_WIDTH_GREATER_THAN_EIGHT which has a default value of 256. 
    *   So, if user does not override this macro then this covergroup will create 256 bins for ARID width greater than 8

    *   If svt_axi_port_configuration::use_separate_rd_wr_chan_id_width is 
    *   programmed to 1 then svt_axi_port_configuration::read_chan_id_width is
    *   considered for creation of bins. 
    *   If svt_axi_port_configuration::use_separate_rd_wr_chan_id_width is 
    *   programmed to 0 then svt_axi_port_configuration::id_width is
    *   considered for creation of bins.
    *
    *   Example:
    *   If outstanding DVM TLBI transactions have the following IDs:
    *   ARID1 ARID1 ARID2 ARID3 ARID4 ARID5.
    *   The bins hit will be 1,2,3,4,5 (for outstanding transactions with ARID1,ARID2
    *   ARID3 ARID4 ARID5)
    *   The coverage is a continuous logic. If there is only one outstanding 
    *   transaction in the queue with unique ARID value, the bin 1 will get hit.
    *   Subsequently as and when new outstanding transactions comes with unique
    *   ARID values further bins will keep getting hit.
    *
    * Applicable only when svt_axi_port_configuration::axi_interface_type is ACE or ACE_LITE.
    * .
    * Reference: AMBA AXI and ACE Protocol Specification: ARM IHI 0022E ID022613; Section C5 
    */
  covergroup trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range(int num_outstanding_xact);
    num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid: coverpoint num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid{
      bins num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range_0 = {[1:num_outstanding_xact]};
      bins num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range_1 = {[(num_outstanding_xact+1):(2*num_outstanding_xact)]};   
      bins num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range_2 = {[(2*num_outstanding_xact+1):(3*num_outstanding_xact)]};
      bins num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range_3 = {[(3*num_outstanding_xact+1):(4*num_outstanding_xact)]};
      bins num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range_4 = {[(4*num_outstanding_xact+1):(5*num_outstanding_xact)]};
      bins num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range_5 = {[(5*num_outstanding_xact+1):(6*num_outstanding_xact)]};
      bins num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range_6 = {[(6*num_outstanding_xact+1):(7*num_outstanding_xact)]};
      bins num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range_7 = {[(7*num_outstanding_xact+1):(8*num_outstanding_xact)]};
    }
    option.per_instance = 1;
  endgroup  



//----------------------------------------------------------------------------
  /**
   * Coverage sample event function.
   */
//
  extern virtual function void cov_sample_read_xact_parameters();
//----------------------------------------------------------------------------
  /**
   * Coverage sample event function.
   */
//
  extern virtual function void cov_sample_write_xact_parameters();
//----------------------------------------------------------------------------
  /**
   * Coverage sample event function.
   */
//
  extern virtual function void cov_sample_axi4_stream_xact_parameters(); 

//To collect covergae of dvm multipart covergroups
 extern virtual function void cov_sample_dvm_multipart_xact_covergroups();

//To collect coverage of snoop dvm multipart covergroups
 extern virtual function void cov_sample_snoop_dvm_multipart_xact_covergroups();

//----------------------------------------------------------------------------
  /**
   * Coverage sample event function.
   *
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for covergoup read_outstanding_xact_same_arid_cache_modifiable_bit
   * and read_outstanding_xact_diff_arid_cache_modifiable_bit
   */
//
 extern virtual function void cov_sample_read_outstanding_xact_cache_modifiable_bit();

//----------------------------------------------------------------------------
  /**
   * Coverage sample event function.
   *
   * Calls built-in sample function for corresponding covergroup
   * in order to collect coverage for covergoup read_outstanding_xact_same_arid_device_cacheable_bit
   */
//
 extern virtual function void cov_sample_read_outstanding_xact_device_cacheable_bit();

//----------------------------------------------------------------------------
  /**
   * Coverage sample event function.
   *
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for covergoup write_outstanding_xact_same_arid_cache_modifiable_bit
   * and write_outstanding_xact_diff_arid_cache_modifiable_bit
   */
//
extern virtual function void cov_sample_write_outstanding_xact_cache_modifiable_bit();

//----------------------------------------------------------------------------
  /**
   * Coverage sample event function.
   *
   * Calls built-in sample function for corresponding covergroup
   * in order to collect coverage for covergoup write_outstanding_xact_same_awid_device_cacheable_bit
   */
//
extern virtual function void cov_sample_write_outstanding_xact_device_cacheable_bit();

//----------------------------------------------------------------------------
  /**
   * Coverage sample event function.
   *
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for covergoup trans_axi_num_outstanding_xacts_with_same_arid 
   * and trans_axi_num_outstanding_xacts_with_diff_arid 
   */
//
 extern virtual function void cov_sample_read_outstanding_xact();
//----------------------------------------------------------------------------
  /**
   * Coverage sample event function.
   *
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for covergoups 
   * trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid and
   * trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid 
   */
//
 extern virtual function void cov_sample_dvm_tlb_invalidate_outstanding_xact();
//----------------------------------------------------------------------------
  /**
   * Coverage sample event function.
   *
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for covergoup trans_ace_num_outstanding_snoop_xacts 
   */
//
 extern virtual function void cov_sample_snoop_outstanding_xact(); 

//----------------------------------------------------------------------------
  /**
   * Coverage sample event functions.
   *
   * Following functions triggers sample event in order to collect coverage for covergroup signal_master_valid_ready_dependency.
   */
//
 extern virtual function void cov_sample_awvalid_wvalid_dependency(); 
 extern virtual function void cov_sample_awvalid_rready_dependency(); 
 extern virtual function void cov_sample_awvalid_bready_dependency(); 
 extern virtual function void cov_sample_wvalid_awvalid_dependency(); 
 extern virtual function void cov_sample_wvalid_rready_dependency(); 
 extern virtual function void cov_sample_wvalid_bready_dependency(); 
 extern virtual function void cov_sample_rready_awvalid_dependency(); 
 extern virtual function void cov_sample_rready_wvalid_dependency(); 
 extern virtual function void cov_sample_rready_bready_dependency(); 
 extern virtual function void cov_sample_bready_awvalid_dependency(); 
 extern virtual function void cov_sample_bready_wvalid_dependency(); 
 extern virtual function void cov_sample_bready_rready_dependency(); 
//----------------------------------------------------------------------------
  /**
   * Coverage sample event functions.
   *
   * Following functions triggers sample event in order to collect coverage for covergroup signal_slave_valid_ready_dependency.
   */
//
 extern virtual function void cov_sample_wready_arready_dependency(); 
 extern virtual function void cov_sample_wready_rvalid_dependency(); 
 extern virtual function void cov_sample_wready_bvalid_dependency(); 
 extern virtual function void cov_sample_arready_wready_dependency(); 
 extern virtual function void cov_sample_arready_rvalid_dependency(); 
 extern virtual function void cov_sample_arready_bvalid_dependency(); 
 extern virtual function void cov_sample_rvalid_arready_dependency(); 
 extern virtual function void cov_sample_rvalid_wready_dependency(); 
 extern virtual function void cov_sample_rvalid_bvalid_dependency(); 
 extern virtual function void cov_sample_bvalid_arready_dependency(); 
 extern virtual function void cov_sample_bvalid_wready_dependency(); 
 extern virtual function void cov_sample_bvalid_rvalid_dependency(); 
//----------------------------------------------------------------------------
  /**
   * Coverage sample event functions.
   *
   * Following functions triggers sample event in order to collect coverage for covergroup signal_master_slave_valid_ready_dependency.
   */
//
  extern virtual function void cov_sample_awvalid_awready_dependency(); 
  extern virtual function void cov_sample_awvalid_wready_dependency(); 
  extern virtual function void cov_sample_awvalid_rvalid_dependency(); 
  extern virtual function void cov_sample_awvalid_bvalid_dependency(); 
  extern virtual function void cov_sample_wvalid_awready_dependency(); 
  extern virtual function void cov_sample_wvalid_wready_dependency(); 
  extern virtual function void cov_sample_wvalid_rvalid_dependency(); 
  extern virtual function void cov_sample_wvalid_bvalid_dependency(); 
  extern virtual function void cov_sample_rready_awready_dependency(); 
  extern virtual function void cov_sample_rready_wready_dependency(); 
  extern virtual function void cov_sample_rready_rvalid_dependency(); 
  extern virtual function void cov_sample_rready_bvalid_dependency(); 
  extern virtual function void cov_sample_bready_awready_dependency(); 
  extern virtual function void cov_sample_bready_wready_dependency(); 
  extern virtual function void cov_sample_bready_rvalid_dependency(); 
  extern virtual function void cov_sample_bready_bvalid_dependency();
//----------------------------------------------------------------------------
  /**
   * Coverage sample event functions.
   *
   * Following functions triggers sample event in order to collect coverage for covergroup signal_slave_master_valid_ready_dependency.
   */
//
 extern virtual function void cov_sample_awready_and_awvalid_dependency(); 
 extern virtual function void cov_sample_awready_and_wvalid_dependency(); 
 extern virtual function void cov_sample_awready_and_rvalid_dependency(); 
 extern virtual function void cov_sample_awready_and_bvalid_dependency(); 
 extern virtual function void cov_sample_wready_and_awvalid_dependency(); 
 extern virtual function void cov_sample_wready_and_wvalid_dependency(); 
 extern virtual function void cov_sample_wready_and_rready_dependency(); 
 extern virtual function void cov_sample_wready_and_bready_dependency(); 
 extern virtual function void cov_sample_rvalid_and_awready_dependency(); 
 extern virtual function void cov_sample_rvalid_and_wready_dependency(); 
 extern virtual function void cov_sample_rvalid_and_rready_dependency(); 
 extern virtual function void cov_sample_rvalid_and_bready_dependency(); 
 extern virtual function void cov_sample_bvalid_and_awready_dependency(); 
 extern virtual function void cov_sample_bvalid_and_wready_dependency(); 
 extern virtual function void cov_sample_bvalid_and_rready_dependency(); 
 extern virtual function void cov_sample_bvalid_and_bready_dependency(); 
//----------------------------------------------------------------------------
  /**
   * Coverage sample event function.
   *
   * Calls built-in sample function for each corresponding covergroups
   * in order to collect coverage for covergoup trans_axi_num_outstanding_xacts_with_same_awid 
   * and trans_axi_num_outstanding_xacts_with_diff_awid 
   */
//
 extern virtual function void cov_sample_write_outstanding_xact();
//----------------------------------------------------------------------------
  /**
    * Called to evaluate if there is a snoop transaction to the same address as a read transaction
    */
  extern virtual function void evaluate_snoop_to_same_address_as_read_xact(svt_axi_snoop_transaction snoop_xact);

  /**
    * Called to evaluate if there is a snoop transaction to the same address as a write transaction
    */
  extern virtual function void evaluate_snoop_to_same_address_as_write_xact(svt_axi_snoop_transaction snoop_xact, bit is_at_snoop_addr_phase = 0);

  /** Samples the trans_master_ace_lite_coherent_and_ace_snoop_response_association covergroups */
  extern function void ace_lite_coherent_and_ace_snoop_response_association_cov_sample(svt_axi_transaction coherent_xact,svt_axi_snoop_transaction snoop_xacts[$]);

 /** Samples the trans_master_ace_coherent_and_ace_snoop_response_association covergroups */
  extern function void ace_coherent_and_ace_snoop_response_association_cov_sample(svt_axi_transaction coherent_xact,svt_axi_snoop_transaction snoop_xacts[$]);

  /** Samples the trans_master_ace_lite_coherent_and_ace_snoop_response_association_back_to_back_xact_with_specific_id covergroups */
  extern function void ace_lite_coherent_and_ace_snoop_response_association_with_specific_id(svt_axi_system_transaction coherent_t1, svt_axi_system_transaction coherent_t2);

  /** Samples the trans_ace_concurrent_overlapping_arsnoop_acsnoop covergroups */
  extern virtual function void trans_ace_concurrent_overlapping_arsnoop_acsnoop_cov_sample();

  /** Samples the trans_ace_concurrent_overlapping_arsnoop_acsnoop_one_ace_acelite covergroups */
  extern virtual function void trans_ace_concurrent_overlapping_arsnoop_acsnoop_one_ace_acelite_cov_sample();

  /** Samples the trans_ace_concurrent_non_overlapping_awsnoop_acsnoop covergroups */
  extern virtual function void trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp_cov_sample();

  /** Samples the trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite covergroups */
  extern virtual function void trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite_cov_sample();

  /** Samples the trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp covergroups */
  extern virtual function void trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_cov_sample();
 
  /** Samples the trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite covergroups */
  extern virtual function void trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite_cov_sample();

  /** Samples the trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_one_ace_acelite covergroups */
  extern virtual function void cov_sample_snoop_dvm_xact_covergroups(); 

`endif // SVT_AXI_EXCLUDE_AXI_PORT_COVERAGE

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * CONSTUCTOR: Create a new default coverage class instance
   *
   * @param cfg A refernce to the AXI Port Configuration instance.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function new(svt_axi_port_configuration cfg,  string name = "svt_axi_port_monitor_def_cov_callback");
`elsif SVT_OVM_TECHNOLOGY
  extern function new(svt_axi_port_configuration cfg, string name = "svt_axi_port_monitor_def_cov_callback");
`else
  extern function new(svt_axi_port_configuration cfg );
`endif
endclass

`protected
.1LY2LUf1Uc0eL<_cJK9=A#:#3E;[5KR5:M4CASIfY3=1J=H3PP07)C13/fT9??L
Y41EH/LJ@TXKLZcN:E3b/2;U>716&A4]F67Wb&9aPA,@9DX?Kg,Y5=,-&TP[=<UU
B4.2J&B7\0-V/T&G)T7e,V]J2f2V0P9\#bM),K\=:bX<PLKCN(P]FTdAKd<)_.?-
]XHbcZ,e[A?Q/B??]Z_0&&,1\P25Pb[UdDg1+gA:bF4ILVcQLCdMGVT70/@PcP8[
9Q8+9\+Sb+(;f6EY<_1X\KNL,@cK74d@G5P<QgJT]N;952W#FW;B;#B<,)U[ALYE
@>05TS/2W<L6BKQWS0XR\Q31\&eXTX5JIE^#^+NN-96]<-BK+ZfbV\)>C,/Z0KK;
\X)1a]B(IU5XU:5K)(PS\:Ng8A<]B>SI9VU#V)7.HNJKNB63a#::JC(.dbPYcEAD
[BZMgB?01cJ@@7TYe/8Q^VV>Vb\P0)gT:=Ag#.#@[^U3_]T#N#ZF1/6:L<2)(aG?
U#QI.-&#93M.7D\^18&(A:)M3-1]51?DBS:AH?24>VF]gC2bC6eT)6(A_I.\F:RN
+gE:ZQ#;Q(Z]ePbdPbNSB#]V&&45O?LR.<R]ZMOTDe40K])B1KTF>B(2K&1M@289
fGc,a[H[OaA+df[LY>&LOCQe<#S=-<]I3/UMcL9S,A3^GMP:3H)f\eF:@&@f4-I&
6>fFM-S,S\>C[VYLaA2/8^&_;SCAWaLPF0Ka5;V:-Gf1<5<3JLB[]#K/R?9GQ8f[
4]]]gEKO<^A);P/[?Z.8e.&gTL];31L?[aL_gN<@C)>-f2W+5F>8aI<P_E@PI@JJ
7a+5d;K^\P4f/[#OM0F-R6T4HLT(1[A+UfP,EI?LaP#COJWSU=AS9HA_/g>VW6RS
EG8Xc5IU3EQ+(;DY2c)e9K]d@6=(&H+X6^6GNA/>85&CJJYI4R:F-^gc?,7gN^)@
/e<M&V5O-004]A?-.FH</C]AMe[S53U7>cf_^Id4;WPJ\F:[Z(T4(:BV5JZ0K\@M
_+,N0O6+ULH@=IEWXK;b#NCY4gE&]M@Z4?AQCRg1;MfYG4<NYY8)\T6@ZGEa,^dR
NH48(UB#BLaX,P[\=::f^(3UgZ65d/((R,BYB(-<9I=#Of\EGcZT[=P?XXNBO8X)
b8.5bK;^gf4&M<5I79<)#_7E.,T<[/gd3G797M?8=^#0\f\a\<=0^Q\826W8<Wc.
ZVY&?BXAN<1dQAF7e0:#/gJB[[N?)a2G</,2H>08.:5O.)TT=KLa4:BF3gI3YZ7[
DNLc.PG[gY/)Y_#>4gc3^Pg=,2>=?[FFFd9MHS;.VQK:#;>>4,G5?A7XD2&<V/fb
O,L:8]Lb,=JP(:NOCKUJK/C5\\DW86HU68[R?.d=1]L<:2Xg],faE+)>fZaR_:6K
@4(=b5Z^Y\76AL).TH5C3:U;D5?aRTQY(.;1GNICA<a(b[V:dg14fH?)SbMGXOPg
?ZJYJ.0RZ97gT30eBTUY_GR#cPe?I;DMA:7UQVRP(L<X<d?LaUJG:#ZI7eMQLD.-
7<DZ&M<7_MTdVV5B=D+]VE^IHF]b=]O^ZS<Sf4_CL9Og[0BeeCXZH51MV/c^8;ON
(V10,186c=3KZC8Re(?MT:NaQ>edaX^\&L15C2)NMR,2f?CTW3(^-5dT[:QEQQb@
>\7(IMG+_K.eS;8W7f&7;BS7I=3eS+GS9U+1bFVf>/5Z\aC]fHUYP<P7gXZS>&LA
UX/=&0+?AXd@0XZ+c)#(WV;B/I(+_:.X0G:cQ&Q[_]((VK0H(>I4=I#<A6WHLUOD
HDO_eP;_[9H@\H6XaIfRMA<;++W,9D+])eZFZY6^ASI,4A,aV40_gHCV2B#/&H#<
aX/b]1(@\]g/;/eW(V]4E9X:Q)>5PJf?B_RW]X4T-6&U.KMW<7Zd2?3^D4];^O8.
[+D-?ZbRPgO70<]Of>B-4:LDbR;JJQIb>OB-:T:^[c4,E971D,2M.]M5]WQRb?N-
B&M,fMF]7b+XNIF0V)/)Nc:?F^24H[JK,.XDB3dCD3aF<MMR+A5L,,W[HV5Eg=A@
N-6O?&^QPQG:55^O\]ZL,7[a[V57gBQS+_:/PJRe-g.FP>=K2<UL1K&+T;D2_4WL
^]-6>C-Q2].ZfF[d3BX:GeKB/6F]\c:(S^:+a9Hf4[Q6:-+P=A^H^JS,79O=XN,)
5eJ9(O/--/.fbJB86a@2;IX3EYL_RLCg3P[)-#c+GGD1GXZdcSHR@@]QgcV6LQc>
7HQNGPa3Z_d?4.#f7TJQ3dOD^)c<MBF_9=(9GW3d@SSXPdSQI1&\9YP#+5WQ3+B>
LF[FT=,?-CdKBXdTPd\5/Ycb)6_)/8Q<A-fE0=DDLE;^T<>:S?33bMJXbOa,=D:E
N-W4K3O?BC7R,Z.[C,HEP)K3/aRYC/Z<C>/]#Y\N.<g9<+U9MfGQPN[/B-J5ZV&M
b:@&DB=-4H93A[TII&;-:2WBP9:[HR0P7[a5/c6@<1>#:eQ6D7R=eR^:>3F2O(S;
H;NYVIR-R,C.dO;bS(E[dBC7#6:N5JNNeTA&aJ_#Yeg&GC50723K10(S3L.a[RdO
9H65T(IJ3MHY.^NE\I;dM30/@7@1(/[60@8D?#+&Y3a6SfZ2,^8)104L12@fL4);
&=ONK\O?WEME_cd4FSY;dE8J/@6VD_K+fbIXXc.[g@&MK=NN;7fcSU4^#O5+I9a/
>J\fdV0/aU4AO?Ed2HP0BZFg<G)2&bS.;\^QIH99f+eG_Qc-Z2e6OQEPBfW[F6Q3
+(,OZKEa;2\RXa<40K:DZU]T?8ZPY]/f#OORaEeFg.a#V9AdX?fOZNce02B+W3J]
3:.a]OZ=[]O8BS4,B64TFNV_ELA#^LA6XWBZTR<&R1F@/9[:DVB7GMJ_Y@3/]<_E
61D@1>d\#ce8,\S30g9HJ/\Q)T&-ZI/FGOX<8G6;U:Q0P^.U;1UaV]HS71Y5_2(d
4FZ-d[?-Zc]O;QJ3DP>D&+#^TM:K1&&;Y6eE59>,cI43S6OFHecJZ>NG+Pa7LB?R
).[QfKde(JOPZEZFTQ]2<<Y=UD&;65)8aV\N3+?8RE?G,]2g(.[GSLb(:6]30D6M
/84C(,>4MEBNDS,R5;F+>@R5F2,aPOCWE>5fN.,)([SET]aP3Fd.A\F30?=KW#d)
SS?FM-,W8>27<0NG<[]O>HE4?dNag(ZgaC4.>M8^c&eQ+gU[6XN-B-?Q@6]9fBI?
fg2YNJRPE[?>)ZI_:2NHT6YU.3DR^4eT<&^]V6JOH,G5;/8A_\L4VX&GG]09Ja7C
@B(4>8:LJNQf4;Ve)E5S^fW6V1MTAbH/Gc]Q4Y,DGR9O1S4Vd.YZgcBT:fT@T\A#
S\KF[2QL),XcYRAaY@34#E<01GDGHTJIN0547dW(AYQS(XYUdAJR>D#DEaIGF6SW
;JAD2&^+O@N5Aa[e;KF4QZ/b3;df:f],QDegNIB&+61O1[XG=c51.+-E3Q2gVe^F
)[B)LDA6bGJSMNY9YA#B+;:]P+2>DO.K2IDSA3(5:-W\H=5399NIJD,9;F.G9.5]
V[WW<d:)-GJd6ZF8;)ALM(XP@G=7V[/ZVK5GOA9V<?->)cPYaX/DNFgW)K^C21_g
M&E?PEOEW[HeH<:_.JGV8e&F&eX;25d9?&bBggMY;Hd68/[P<,^gS,0&Z1gD?B.I
d)Q^B[0@)M6/?H]8K78@A[@M+9W+ULOC;2d2+Z2GG(I:5AaYZgS9Y1WPd2-aA@b_
VH/D8gG)GS^UN]DUg]7,4eJ_6QHfHgIVELR7&?c63FaGOT^1N]EW=TC3_?89Tf8A
OdVcE8X4\?1N?+#N9J=5AM]GY.@^A>/,MXM;301/3-V9G.Qcg,_2:-M>8XNY\^10
;AedJI6f7b9J93aA]#;QQG22a0T9K6]FUed7e?Y=8;@^@fAA7;<4^NF[JgAG55I0
-9.#5)\I+M@6b37QbT9]-1IRa<TEQ<(8..#R^.25K@CG@91T=(.dRTMe\Q^]J.AD
R#LdQf(6&^MR+H+8Z]D;.RTS.G;Bdc))0K&2]g8SA>XSbSN\LOL]QL?-^C[Z2+9D
JAQaK7Z\O9U;S@KP5GbN5O0/A;,RK.\#bNROCWO0_KP=ZV]J5=I^<ddY5FHALT(L
BBfb8P^1FF8<+:&Y45>c([+]3gA>L.HMC7K6GLb3c5T>6HI^NQT_J6BST-7#KfK>
DbHV./S6AYS.WGf:[3J9]Ke:aCeS@acD)[aX1f2f\U&:1@O40P3J_&D-6=QM&=Le
WZ/:^PHVNWHc;0^Q6dVMgCE0CKUd.9UPM(cLS<Zg79KX.09L#9L7>#96DF0]6)SO
A_(#>QA3,/\__K[2R,KE-K/e8Mg>XH7OZ7>2CVO,[&?TX&(@Z5SQAd@(CX&E,8<<
FND1HCPK-/,CM0]]]?X7f9ZKX>IY9Ig>O.-8Y-\BUb.R8RX5BUF2E2e9f8@5S;c6
&]&=Ug;51f(QbJg-BA+H@A5a&&Z9,Y2/)7EY)DU2//T2P@0JTB<&)_O[>3Z.5^,0
ALM_#\-Q17[7].XSEKWTGTUC)b@agD(EfQ=C],^,AcVR)S5^W@+dD>,\RCP?PI@@
f^F_<2RO5UOD;Me@KB3b#bDL\B\+W30dFd)Y\O5\U\#J51K<.ZM[W0LL_4\cIB+&
gJ.Neg0G+IJKNFCRA[4B^S6(9RPV/G5/I\:#TQ-<g7Y8^eQYRSVd+&8N(SC^H;]1
[->2\Bc4d/gRY+1Gb)CJ2E:)>ae7(O_M)JOd&dO@/<;QZWK877S#[MUWH2OcD516
E9Q^BJ6;bRUbb8PN]_EW7,MTH^D,P2-a:X^G7]#gGa,+>N+;JY#H\:;Q>9:)D]DQ
e@d2KcGP-F0[@V>aG:H8_W?]_?LO,4CdS5.S@6(3=U7.:G5c,2/T/7WV\<C71^>C
L-YE50=G6M<McfD0/T?>0WF55[c4B;MZW79[<6Z-EeT5[S1[0VWF?=]D5L;BRB[U
6_(\,JaT,EC)e_7b(.G53[29bc&A]KK?)C8F4S@S[O<0+=cfNKdZd60:?eC,.S13
^2de\;#21]D9/M<5_KC\_X\0UdGA#DJ+IYX#1)Y5:M8R=\[#;Se^4cJ>-?ae]>^#
,gfX&9ED@7=W19E1.+JS]4gF?Q9FPX8#U4KXGYB1Ige1T]4e6TQQ#-<WM-SY:IJE
d.5[NFI?0\,0CPKNWA8)XeP^N85Y7T+cD_SJNP:OVaJD[Hb3d=5RR[XXZE=-WA=]
;D^LTDa(>FC^?#T+0D]2TP7/eH,LJ;K6L)3V\P?fB@4O&(gdG@/-@+^\g[,N3<IQ
c.XG_QJYgVI+<g:5VSH71>SRa.E1-AKVZ[CO?>-8K--bX0@J0X,P;NIbWQ4I6g..
I80G<a(V(6]2B/N=(FLWTSD+6Z;e.;f8DcD-/LIDWd/H35L<Kg&PKKX[I&^/:8@Q
_MV>XdN5<&N-\D9DV@.6;/5f7AI0I.-#[#&C^^N5[?XK[<WR2M68^,G4C10g_#+)
S9W\843Ng1.c>;bgg^KM,C)JZ=8f_X9S3.g##5T75QK@gJ9&#7A^]0U]LaMRHN<a
F]XX)47KaQU_]EA2T4?g&>1HfSN?>N3P8dARg3c/BC>&(FTK_CfN21<\#d:SJ\ZU
8_6XbZe9)ZL6?DM;UR])bA#732aZ:L@DK=&ECL/4HYK\]I8+Icb,&4;048:27N<-
cHUYBZU?<>3HP0)K8L_/?VXc1:6MUQ#HQZ3UYS=f85BY51:()-(,LO?Q:Za?D+>&
-Y?CLR^e8V.90:D^;c[CK^OLM91.b\Q:,M,A:039GT8LO>JD1daIBL,4<Z]E>P3R
1=.5AHE0+[dc?1^CV;+F.M_9)C5;aMT?54bVOgU_XCX?Z/[+?g&61+^AN+G(GV_f
4GM,Y/D:S#Ye8M>FTJS2]X&:fWYF;HD;Z5P;/YfM4Kd)/Lg88>Le()>ZVMWf1Q1]
>#+?92J\Qc&3]:32U,KBNGd6-Le=1,8;;#DZ0b:28[KQ[5f]V<Y82YWc;OD1:E_f
]&gLXc.1[D)-:JSZ?)C\NY/>dc9+C2NK5#c]8>4W=e85BAF?8?#FYFcd:XK(\(Kd
N/9.W]A,K;)e.Gg1S_T+31+[9;EOD9[T2M)]#QVaNeGQJ?-FYdNJJ:E?IVb8+ZSS
6C5E\^5@,NDFFR[S8g(cIdY@YPDO8QREZ-9IA+IP10L<5S1d.97Je:e?X_<Q;d(@
F52N#S]G#>((P),H:e(9:d[U4>eXY@ae3-9W=(=FQ(Ye(ZO]9,V&:\,R\EAD_0Z;
fVPQ)O>0c[/1aCB)=UV:,>#A?F-(2396AecJJCe,,:26J^^Q;AP2,CW1[fTW+17;
Sg66MJ6YHKeHRBB59G/-WD>[1?d=8Fc5ZZ15G=)fVa9COA@Ce+QA^A7CFa;N_,CS
K=9dR)I,I(@4A0WaEJ?JREeEJ^0BT.E22(.H#8OcV,U8Cb-WXTdLMYa@>.H^6.8/
QN1B#^417EM5U4J9cR@45?V,eQW<,Z]b#7f]Fd-bHSZEZ@JAB,PfPJBd#fa[d>SB
7CO?++KUNOB.McGK;RA:?TF-4#S747V\F)D/d;DFNM.B:f,@-URbVDN(QY8XMdT5
N/)/dZ9\0N]<>W]W9AZ5\DCdbKD=^;;0MX7CER4FUP5.O2[4/fB;WNGF\MM#g3\3
>_Q&DO&G7JI7_I_R3FDW-4;)6#:T^KGSRQ\>O:/0(MU<6.26UIC[<DDF#)=)FR0S
dU3fUFFgS@]KFEagT6EE0),X6&G8[/=bO8/T)@R1HS8,38UPeeZ3GK\TN)=E([_a
@,.c=PJ?8\EBO8g7;]V2RI?9B6cN5GFD:URM;7B&bJFDG?e13<4O.KXEFK(PgDa[
Y[WfTbDL7CT(b;eX6<1:;XOg/(=J:2&DCJP\[aT-NVL:H,&253D#,3+OaW<[DAX9
NO#_6+0KfTL+[_2MJW4J.VIdIP/\5_:fTa;.,Wcde+26NN(J4#8&D[AcWR_OdT6B
/8PZ7_AbZbM)Qc<QHf4DN\D,dGM)W@=c)B,^4Y7IO5>[0&Yf6ETL@9XUNAfOFd4(
eac5>83W4&^]6,S9=<J4;32DBg-R)ZQ7V5W#M;]#+QU[BaE>-0(aYOH2MT7/aa]C
Q+=HTGBN)_)4ES/-#AS.22=>\>C9:0R))N1GR#4g]&g66#3PRR7BLQMac@R:=ZRF
Q8(1N@O/QM<-K?ILZY,T\SGN153E7Je8#+ae0S9UTYdMHVX^B8@6bcRMb[MH]2[M
VWBSAfHgTUV[1>CdVV=9NGEU0;A?7612+;C/P8U3cJ=e381[L_6EdT7(G)ZAfDL<
VCY=46TH)A)@6ZeLB4&Zf6H=MIAc7?K,S,#H1B+9:3PK0@VK,)^@ZXL),eR06.++
0CJQ8\JX0]@3T;X>CIO^f7&-<2PNRO6Ka:)<6>be5C@\.Y;+49gNBY@X?EdJB_,d
M.7:)O1QV:g)4C/Z7;(<W#7MQO,GL,/C#^(2S=ac-;8_T8N8T11J1e(2aKU&+H<T
YbS3c?@XNZcK:?LG0\,bB@@#\&F=[g,9fSU+a<8[0JY1:U3_.1/-:-QQGCO5]_aN
MFGL#\FMOETP^]B7]APO-80(\WF2V>-/[-bc4357=D0+a]8G5E_83<]GT(,,DF0H
XE@BHCYSSQ-VEA7A/R?XGA;^,cCC7.W[I,)A7[B+E+f7f)S+\=NKW-&Y<D,V.LBe
U@N][<e&IM.W,V(,:bWTC5,4V7a_QO=W0]N3.G(E(72Y7O,:UZSN<BJac(c_cA:O
b8BH4.Q+/:@M-,FE)+f#b=ZFK<HF.N@.DL-f?AY&Oc4f[a3a),[(G?7_<LIOG/#<
I&AH;0P=9fG-1#6NRWSV)OJa0Q=5(H[MM^R(59_>d:FTT8LC>:),eQdRWBF^G]E>
Q+12/-G&0DZ:B4B_74+,6_(&&[eF>T>6aYgdE,C^d&IFRf#)LAd.@O])P/KI@c\=
Cfgc?A[bbEYAB#fX(XYJ#NI\^:01\D\I51YSK</F/eL+a1cTKF0d?H7IN4NN(c=F
)1:-W8NfaRL;).\;)BXc:&Q)O@?Va]e@L#7c5F]Z)+?UNJdUV@FC[L[+D-O.WZ^<
M^?2+eT@+D#)KFD4#5)-@PL>M7Ed#G.CIT0;&6[^05N>8QfcRL@/(X6:.5=3-c9T
>[\?,0P18##>-5[<]XO^]VO^.G/06O6B#;=bKRCdZF?df)I)7</3=d&?Q]M90T3,
(?N-gc;7eBEGHB?@@C;<af4=2Re2DP6+^R?DaO^<U)b,MB8/8\K@9>MdYT&3&P[/
J>K2>L9B#B4<B]JH4F7)2DKU7,bE/WUQc2&2NA.Y[OYM<A7Qb5fKOgg>DM7TY4aJ
3>=e]=8@52e0R/GEO0ZPb\gT1(@H5BBSOZR+fH-\g)IObJ3Y>8S#)2;G5[\UV]+^
>>a&c:;5?2e[A_G7W,N:J?V8f<#+^^L.XI2O^ZB@FA@+36NcUL?G/7?MD>0-0..?
(c6?c(U.S_&Xcb)R+,7V.4:K/@^L(&J(Y&g]RBA,U5@.Y4S^-bFa^53:RIFEI(>^
M5J.K+a2,a?Lfb^^+6BOS,bAFVeF>a0gBFFCgA0>Oe,PfP0/G8?VdQ._J@g3AAgX
8@=#/E/1FJN&BXg;F/OM0(<gHZHTe&4gA3TWP;7YXIRH6BLb)N<ffb+5Bg>)D[d)
EgfVdM4=K<FPDJgE:LXAM0K<Ng2aec)4E@CeN.KC][IKN6d#MI0^>1E\HU5M35QS
EG=&#\5ARe&9ROF:H(6L8>,<Yc8?1_<E\67e^,)GF^&6W+c:#bGa)<\<;g6,YB\6
@P]2ES?I8<9--.\IDg8(N(/2f-C>Ob_E/c,bV14J1-J49^Qd>]B+8#MNLXTK0K00
gP7KRbNAd5UJ53TF\BXB@LdP5JBZBMNJCJCG-O]J+cB^^M#ZbdHYLAgNN3<-U^1C
]aMMYN(#D,aYd+6Od]]U__9?KA^CU0D@L+2V#QQM=8LYPPRf7<?UC<begbF==P,=
@?Zd/:P=3?YS;_b1Ie^/L6V<<=011CV)AYQJMf9g#)aH]Hc[7c70;UE,\Y^Y1gXY
B^0SgM:;C8,2C=M4:4-[=:;]94CX#^c_Ga[a@GY(d=W;&LS9280N^gKc@XIUa#XH
&#\\WX<cJVfMH@O,f4N=7B.NL3EJ&]&.7.+QAU9]UL#]:?>fd-HI&G6V:K,(_eWa
ega/N?AH05N@E_(U@@8HYOU=R,8eD\C5J91)#PcJX?-(Y56#:<KV8+\51:P4C:(=
6dAD.8[WSYSb(G4Q\WH6TP:fZ6Of#2c6I#]2=06fE>GB\/)T8C<N^F?N_LT>6VV]
4JJZdG,5^;S5U9-+?YJ=&OH-Y<J,0[(7C?WQ>Z95fU)]@PKa+\S7>=[8:eXVKQ3<
KdZCRLE7,//EKF:?C&g9GPM1T720K:YgN3e4E.=6C32+M.]I^#GR(A3,V7b)@IQK
D?/9:Sd72.@C3B/^AX[9C1S[P8c29KDS2.?K79;G?FR^[5U;VbNYHb<CA-R=cGND
DNee&-S1XCH<7Q=(L6]:2e>8e(#KbcL2a(RQdC(KI0DaA<I&Da?@S<X.3(?LUK)3
HL1(=2^C+?W15b0e?JMV\0D&1.9c(9)L1.OP4;09OBGa#0-gaQSb<T#1E\R],32e
P4gcb@K,I.Bc/ZET3(3&\c7T:K+P11.17/X#/JEX@HYg55,<?\,1>f.X0-XQURMI
K7A19-bbS1Bg5G,@I#9-IM,Zf/T+RA)+JQe2J#TYLe+egfC_&+Ra4c1<b,SANVF2
4]8e=;E>I\/@UF(86d),F[>2(EVgb3O;-=W5-e5>\CK>B\=UDK?+FO<LbBC7M\fG
@RAAQ3,YXK1LB59I?2;2d:NbY;=3:D\YPMMM32PV.@XXWDbT;N.=;-=fSYa6da76
^f0><+8H8TeGRd[M+5@6,]PGD\D;@^4eT3:U9(,b+KQM574Z8U-DSCBV)fI?]PLc
;/Te7E?Sf/A?;5b)TbKI3RGE/)ccSS?/02EGOH)RP#<T]>>dGeNVUMgXVR)P:.7N
^=7OYJOOLM?.33d^AH3OYA40U6\d62RZcDP82?LCG1e+&ZLWaWA/Tf3N7aH0NX@J
S^d;T.>Fc7UeR=N0)Xd5BP\KZ[LFJ_S=QU?C\@9f=DIL(EF4T5O0V?0\;),:4^Y[
VAf3UMagUM#;F.IaKC)fV9B5c;R&\&(G:H>,\N:]W4P13c?-/=8J6V]7E\YR<?b)
<+T)Z,<Nc#=#&47Y?//T=7_63[H+@\T\_E,=&@[=3D9aaWAHe>bIIM[9836VXMJ2
g=eB>g@UeXFNc.8,7CM3_3U0A,Y3YETP8VZ4N/?AcP-987P1Y-[Mb@9E82M##L+(
g.Y-e0SAA<?[O5]Y_)-b+,@C;-9#O=]^dN9JMf@/TI&&Y+85-[D=eM\AR.VDT+1U
f>A&+O1LGCP1XdX2bI]>6R(gIf3,E/3HY2<>0_NEG&13\WA-@478O22gN+-I&Y8V
4:G(1U=P.AK?f_DdTf5,/4Q+TW^M.-e0I@K(>#g#U>B^](Ld]DZ4SBI8F=DeT1#Q
0286OPR=9LRXR<F^+8#36gG^cIMK&]9E(?@R:f09EW3ZQEXF6F?]9[2=\=,/]YMA
fe2J?;YS1?\\-fYF_W1Y4REE&K<Db4G9-L@N+,JY+](McSKT:N9>M]CC7#:CS?(F
#V]QRX_ZG8fc8YH@>.[=+IEH#=+g.V&U)fS(OW_eOXX,3\=M:WVSFc(\?b@+KV.\
ZDZ<8bK)aG@1@MSQ8JTL22[VPX5C;gSYQ+HOP_1736L:E3]HJ-F#NOf=,0T.VO;.
g,@X>E/[-478S)&3QSG(88Ma<adTb?VU9=\:<@;<0Y5,XbFV]cg\/bY#T([+\DdX
W\BL(/YS:8#c:;3R=b7Z?,cRL>_,aTYcX:S-INLg2H#1])?aP-C=R_6S=c&HNBa)
-dKY9XE>#]X>cXNMRD0b@,g0FVcOeO0XKef;J(:DcL=^FU>3@SF-MAfeENO9:-Ha
QU7OAdF,g>[cJ-?D&Q0(^1V6=DQ-24:]4A^(R=1Af7]Z\Q.G>D@Z4OQP0g=W4)W\
-DOS3<d##RGbH1,-UgT_H4C)4WRgMBdXgC.-XIcMH&8a\5CH;H0Tf4I&;.U7cRFa
bH>L0XQ#VbbW3Z#LN]TB.,#[TANCYK4WH8ST0O.cTbMdMfLO;Y78I7TF-^?.YbZ@
J7RLW^R5.K6A12CC-5&[gXL.>U(1T;NCf@#)L&9D1DKK^db+4(ZY,RLe+F\K#<6V
]P)3a+CXQZI8b&M#Qf#YW8JdXNW<?R\QG8;8]C.VQ7TR@7,RYE3J3-RD?L+GQb\@
NeL-844C&=OeC;NAN62?d+](Q;9ISbRgS>UYU9K4+gD+\/]8WF,7^G^@#0#Q1cGA
\]a[.=a=EUZ>@.I=7L01JcXbPNbf4>W\dH=X4-c^KI:79Cc7BC71>YFFF9.VaZ,g
N=@Kd]M^8&TOC+C6J;@-T,F&PHe]EIGLQ_K-33#&ITQ625YZ4aVQH6#_@__#(BH/
Mf0[^c)S@\H]ReE17b^YJXITH\-I_KA;;Y>GHX/.L.R]gFd.14W8R.(VPFeLS/L\
B,K&,L>.FC#-SIVK,aMO?)0^0A7EYIY-8+9GXH:C>_5-S7G0f\(.ECd^&35d1gH_
=Y^0>C50<(gc,(RV9#);4N-F<2S])\f)R7@-7=B6BD&_\4Q/ZK=^Cc<:+J/HCI9=
D<]S<F94^M#I<](b-:).]]e-XaLAS]MgYO/8[d,6\VbWfKTZ/:\]J9K4?;=GaDYL
#2ZbUaf85;W2a/)e?\bX+O\U.)0-USU[;W?I^P9f7MAb\D?FSEY?;)MLgYa+gf(e
9La^8&N[W/BA:4#7N-@gFPL1BHOCNBKD>c4JM@)e.V2)O@YB;gV1^5PL?9==X3Q6
<Q@MaHA9fR7PeZSTB#@e\6HaFWHROG9=Y7+X<IZL/\MLMX+b4A5<eGY+4Y@=5(+E
#c9Z7YZa?>\]OX@V;EL^H7_;FM9P8Y<;@V?YgaYTc,.;47B?FQ^0@W08#aX5f<ZM
B6Y.X+HX_KcMF:4)23IEeb]_Ae]&DI#2G[/X1^G1L5+#Y^[M:26.+T(<Q.RZ.L,U
cBN>33\/)NTXHQ(3.NM@6>0SU##W(]PQa@F6L8TIMX:#\>E8d>4(,@A9f@[&)M9>
/HWb#fG9b)Sbf^F69^O\1eB<#80Mbf3PE/H,_@HgfeAAP[JK]c449WRDMYKFRUA-
-;.;?D._/(0D3.E[+.VNYFKNgI?EO7g[6>LPP-=F:X4:Xg;;.JOSK@UD&-XXc<=N
8J,YL.bdfg[/aB,@\EI+2G]PSc3/Z#AcdS774K<G-Q_L,?Lc04c<_2@aCGY:QOe;
&76@YA+/TYb9<I7H8T#RJO@H5.Hc@ReaN3>1?;XU[=;O&\e;G<R&2Z26QG;HZ)=6
cf0R=VB:,AbG]@&)_XYP;^3D;L/O@gJB]Uf1D&W4[-G9g&;4L5DI2B7/Za(03KO&
@C18P:EIF@+5fD/U\/E+QaV0R.MO1^SUXFN@dLHe(@1///;0d5KgL7T6aPI^2)_D
;KWEAI)S:U]>1.\B&HdOH<BN]E+J8;;Y+P642<M<)g16f54CJKPHd/RXAg;W=V44
#&8U(<.d;\-D)DC<C-e[+;D8.9O8O>eX8(0W0^STeZEF<E8F@3WN=QbL]a:MfUDO
\ZKFUDWYaaR0Xc^6]eNT=0I9AMUbbXNL<;#\@:Qgad;,YUB0.-\0G3UO5I-^K1LF
HDD85VT5O=L#\e//b^O4-&2[U.Vgg<M730-J2c[c?]M<R;L_2ZO+(H1C[(:+VCc^
f=+E7c_.P,d7>dT)KNIWH&:f(=cMRK[9RHEGVP#-0Z6]c+?&06@=-;1YcdBA;H,U
R93KO@,aNa:MRM>@4L<]V&W96WP_d;#Ze[WU3e6=WTbIcNcNFFWbce])5_RdZ-.T
a&b39W_5G65^ZNG/;aX,LJ=AEAYK7N#/(6QCE>BBa]:#4(JE9BI8eI)WPS5[Z)3,
Y^&HA5f(^F^gW/Z@S_ERD.Q@+)1(Y-_TRKUF]X@4fL8WQ.ENUMSR?:?L17bg/64=
NNR^ROY<JVP2Y=GMU[Q/ccb5R+2:YG>UTe>J/\fU#B[.=GW?Bg/X#bQd_NUK4V,=
L:LYH=YG@dg/:E(gd4Ee8.IXD@VF0M1[C#f@_)IT]8c,a@L?(fU#N\e]XCX,Z3AK
K+_CH\9:W7T\fKSR[+_6EFPBeX-^a./TcDcSaMbF&Xf4&B6<<M@00g:de2LaU/C&
^&c:[:N)HaEBMWCBD8TX1-^S75AL,=3_UeYWZ3<_^)#^#0FbI/,XDT^S2>eV:6LC
^;a@Pb@6A+@.D3aM0NYee:JI0X3[/?R^.gMP^gHC^4//OcR82LZV:+=^L)P4[e\,
#d>M5:KdN<L>dO\Y=SGD3W>F8_(.?aD[dg(_T(NMLY>]fU/gK[[3a].Ra>RIb3R,
/=[/d-S)P\[_X8I_XUH<+&.AJI54(]P@E]DK]6?+&\H6N_3WVV_AQgfW._YC8TD@
UK8F<AA81TWKUTO?>ea2M<K4+H@I;c]\SMO[XV6K[gP6[NbIBaT@5cL3O&\1#?HO
_I<gLC/B\/=IAGf(X\NU+^eTWRJZgA_2C7>YbLBLK#=@)<0E?fWYYQX>5:fD@5QP
62MAEdTU@]dO7IQ0]Oe@2(^:<.0HHB72Z\e2TfN65_H]F/2Ua2S&TO@SM0L=ON]@
.6-^F<VVNGZb8:g][OWDe:@+ZA2=Y^fI-97;8HCab)12a#Xcf^gf,CZE9XHXTZ^/
V4a=8-,^K[]P>-gfMbS2I)V245K=aYD>EDLDcO8AFAC60K[I.Z1GZ:#=^GIT?26J
]AH+SNgELHZBfW.<KXD+&]#3E7X#[0:+6Z.9W:X^V3(&DGRac/-T5)\ADT8YdJWY
>9_If>O.B94O/e+?I>NG3I)agZLL,W#86FT+5U_QEK6[;eTGIOTVHTROL_;UAV^?
[<^+@:J]94C-O#[Y]M(:-Z&f,1R2IT..F4V3#@]@4Y?1E:_5ba=\V[Y7[E82ce@e
:5^YZC53GSd?cHaY\XcFB.EP6<B0(b)(S=F>S7=GH5,YF8=OX:a]\6B8@e:g2I[C
>+3d^#&[A&PaWafbS=CQJ#02^bg<Z?IE06_EY2?QS&VX+;KCdDIb(2DC-YcFg3DK
5IAJZgO[KLQ[c5aXQ4G[74@FC+Lf+</_,;4cYO6.<E,N@eR1-9]BeOI]7\2[)Qg@
eF]J81.a1Ib^(fW5=FeCQ(&XPd+Ye:g4S7@,/#<M7Sf/dS1#(.4HD@b7UZ,1PL-:
fC]5:4>ZJ<JR[K>Pg7ITHN^,&.(2I5,CKf3BM_A/(ag;0)],D)EQZNL@_=6JF\Hc
G[M<MSSf8C]d#EOd<AEe6OQTaTF<1,(bP;C?6,.3DJd0CCTHX-J1.a69aD67XJCe
O69RB>B?]eLH\<M=gY&_^ZTN4WOI.gT5J6>9Qa##;d:1\XIc)9<^::^aTf<Y8XT3
/21Ma_,J9\d[g2gEMPHd/?dBHS90X._9=G4bC^0C\(;9V/B0^P,;Fe(DDc@Y5Z@I
d@Fc+^d-ANTZ\=AJL>AZA2cB?TSK)UYgMX)X+LUL+E82>#MR[b&,V#313K8@TMe-
Y]TC<^V5bU\a?DF?RXb<897+7O+)beKPfO++1;YT_d[6?XL(bM24M5F84\2Xd5;d
bgR9NM?gJ34YO,QW0X&Z9UMPJ11VM3^5J1.;bCL?APYMO0<7D6Z,#.0<RTTf.e^]
1HZT_UI<MbK<@Wc5^TV3Bb]6,^ADQPH3-4+NXM+3^e_Z63Pe;+233_3<9]EV3aa4
OE8GRQ_V_MMPXE_^TUWa@U,]9>DP<5EKfEPO=4X#J3Z1fP+gO+5B1:eebdGD9cEI
R.&QTd)RA@OI-,N_GI\g=8&L+5U)f71Y>Y)[.-cQ6FHU4Qg6(&37;31VFF?_ff>g
=G+0#[6ZA._H>.K;3QB(9f[e_1MV[,70I1fb]0UARRH_)(ZB?gB+?NKfKGSM<2gV
^JF:^UFC<D:[IN&NK/.g,JO?(0gSAb?3IZ<Q[\Q^:6#?O/1A=96^@(D,>c-#7289
]HE<SLH)5c>))&LVGe=Xc5E(FQQ0@eDJ\D=:d9d5VX>VIV?>U3#Od+6Z3]U4\E+1
[:a;3?a@/FMED,e/YJc4H,RdHX_#GD.I&3O9F+a-S,?)V+#Y(6bB^IGC1C[,S<[X
G<#ICS5VJDFC5:7=B2MS--F=c47\<_OIN=TEHHKJY9,#GA=K;cJ.Ic#X?g71>c#.
Z2c#SNZ-R\^:d4e\]8XX9GH?3+Y6?&:T1R00OX@KDM+6>CdC-R+XE?JBD+A\38Y6
f#T37bZ5<7N\d;FHRD..VM:UZIWVKU-gfSdK,f/74E3P=f)>R]/9V899-Nb6??eY
TA+SE=1H.;S0D/AS^X5N_P\_WO:ACM[4-V1T@KF4a:-]dMYE_IS_;A5Z3ce7A8d0
8PL2DQG5.Q/c3+7TM(VD/(,L6PM-8bQ&3fV<2;<QTFA1GaPc7.f@.Y[Q(KNc#G_)
2#9#@G;/b44CcHcN;_eG,a,KJ3R;PW5f9AZWc1L[Nb>(;OCA6YEL@N?fE.X-G6/X
Y08_I&6]H)U#Ug4J@Qd-9.:8AX>^8bH[dNJ,O[0ZS505M^B;1>Y[UK>X2)baME>4
HSG2B>7>(0_[[7aXB.;FY4TQ75Cc0S)F)BX_YX(9QB:TKW/]4REfPZK5CZ31f5,;
]#4f:,&dUMX3B.UN<\KI[^#(KUR/\/?@>)\[K\4dHdC5&5P1)R1)2Q?.3\5U..IU
O@(9&[-X)&:=eL8.e1^(_3\4>;Y79Gb7,557?J<R#V;?6E?M/f@)gF;&cV#a3f8K
^@(M&7WJYA6Q5[?X@6A,Y55/M<aE.-GKR/aV6ID[HTe<<2]WL8SF5X(S8c=?4dJ0
QH;=.IIT\:F7L,MIb[,H4BVURE5gU7K&ORcFJE4W;^_HR<Sa0RQ),L0O@85B,cfY
UELJH>NG]V3W8/ES^Q#P+]fL3[X=cOa1O0+MB]7,O<Wa0BcM]^EHY7&/T\)f]3Ff
/GfE):J2W,cN]Pa[(TdLFK6?=.1NC^+]G?RW=]1=/+8,dTf),^8ESL1O6B)g5W=(
_L@U1U>C;UfXJ@33Z6=W;;-PSWE3KY#HcGcEWYF1dR,P#J:70#?Ng+CKT@:-egWD
-_cGLD:Y4<XSVHSL\>e3QdG1^+85+,-8VPRF=GgY;1>>\LO&).R2dfI0agS]cGK2
07]<</&9+IGUB--F?e0_NcNC+XP1^4&/O[CJ,P7,]c1BBX5aL4REeXZWQg>MEU8^
QHGV?+:Y9G_f?GE2=7GU:X/CYQB-3bC1?-)_QR#5+1)Q2]VBVc\d:660[((_L2_9
J&85AF1FEbaSU;gE?PMA,>=HS3&J9]K03FN1g1J13\>>G0^I9MG)L>G4NFW0CEe3
,)NAPT#M[>;25YPYOO/C37089I,0;IC3>3,HS]YZ4LP0Y[.UT1e:<_)?a,eTB8M5
:D1B(.]6?CY&I796<XT/HUa7CM__X^;#_KZ]WaM0:bCeGPUQKQ9>K@c-]f4Z.M?Z
W7DQG\0O7_TUP]+L/;eCA7;X0]&]dN2AEZHaG?HNEUD;FWVUTbWcTSd6bS5XRH/E
,A>ZLH;>S#92(@_5R<H-D/:S[70dQJf@.QA/VdSS1aXM>UO0FZH8/FG2L+gce3&f
]MJ=-154MZ]E.@3eaa>77<::gJ;/C>[]<BCBd,g2JWb2KI#7IHa@+WYG-HL>N,]T
dPL_U;B,JH(V\3?YIY3SN(M/aFV;[UF5]M_80EKCBO#>=FUc<MN]8BUSA2PE#GS(
AII?<TO?3g_]7+=202gR?>G#QEG_XFU5X3IHAQG\/:PgABY4YX#@-QZe&W[W/f9C
IRGW6S/P_[TC>BHD]9G+Z5#DL^-WJD@]DKIQDW+W7GOMSSAI//FLIc&AD_^=FW7a
R.NW)D8[d.=U3)&:3Z^JO?FL0X>79^#D9/Mc[YXgeNWN-\BA_O[YR>);e8=<JC[>
dUGabeONC)8:26N,OG^;^WbRF7FX05-:7ZW(RX7ZD)H]TW5XFV2O;,HKQX;]UAWW
@J#Ee^C&Z+0Z60fIa@J=(TMgWe8MF1c@d#\\NOU;@=XHWCNAIgE)-dX\>L&YGGgH
NW0Q6fI<C&]4f=PNNU0c#_=,aQ0<J1d+S^=/4YCR4\MQE3=V0bD4;_SV9;?>gM\f
&PR0;M#K9K#Vg@UOg85@><C0A=C0N[>[gY/WbfG@,-90N2a/d9c2_B_.45SBDO34
;L#<7)CQ)7/PCT?fC04VII#Ee]eX./aS?P[9_A,-(O7UE=X0QL77PK\eAEY-YN69
Zd/8dX3X7XIK)\/.2[#RJZ>L\8)ERf3M=cfWR6\V8S>WDJ<F_GKCBc81LHMO,IP.
RJ9Z3./5==4NRgEMU&U/#XT^HQIKIC8C)GRB2Kd\4==E.d_QSHe(RdC,=BaCK1FC
]Z1R\@D52(gIOd]YJP1e-AS_OTBe5H0&U-\TVO@4@>)RL8B_Eb70CU2e-D.P.V2e
TS(X9]eA?5CAUB3WQ(.]a)3?+W>,21WMDga.F>O57.5565d@OFcETCg0,3a-f?0?
E?]@CE<4HZ)cL>GS(c1a-Ta?3TV[D[TC5QN->6IFfbXXF(W(Jf4Q#g\09Y846=\Y
BS@7G2<5#bOT]+;M5XND1Oc8):7]F\X4.46P<HU\0FTU-0^DSb+&80g)8N#_1YYW
QZAU+d/42/eD0D-CBSCLggYb3G8,;@.f>(-;<T;2Q0L+d8=eHY+J&fba,XF>JUc+
QfZ;TTH8I3++:(;#S8#cH7ELGS_ESB4&((X:CB.+f&?5OHQJLQ1ae?5#.P8M[B]0
\JX9O53^DdD19=[HaFb]f+0F/M+5d@,&&2KXMH;V<;.?.cG7#0/RLV<XF(>,b<-C
_<+(9K&,41JZWa]fM+QR(/NE4XRYf-TO\E9gE_VT]Pc;g,Y9&3016-:3g+2Vf10K
D0aPgb]MK68A.T-ZW?,?V9UCUd9a2(,=:gI>Tc8W6]cBG=2_>SKgL-)M[)bX>E>V
[#TH83@@P8N)9^dC<(&/99T)<R-Hd);Yade;10(LF:#7A>.WKQC9<+AA+U\<C;Z_
/=/KX,\H,a#5L^^89^g4BVK/&@E_EY[S@K5.K]-e9ATfbe@5Bb5N6P])bC2T&FLP
ccf1T)3:=&R.COW>.[XMG#-YFfY.VXIBP@_Q8D\I1@5YQFOc+C6H@>#+g9(Z(P>R
E87D1(EA:4U19-1K@M1O/VA#RT6:)DT4H<]?N2YG-Y1>P0)MH./R7ITB[(Oe[cG]
QDBE_\d;XU>F[>D[8^eV=f,b.Q#+f(PX(gZB14QR[AOUa=H/0HTD]a::H77a6R5\
+(gFaE55WRMP&f+BR<M\>+#1(^_;.:/Q]=gA1L1(9FKQ@\@R.9-:^[EbZCYO+2#,
/__>/2&.<XfMCL2V<Hb:X7YT5ce,ULcH,TYC<4/aV9=a)R#fD1f,TB+R64-.IfL[
5\e4>\&QP&Q63#dbWZ8>@>g.=^c)^C&ZI,B6G)b]4OVC[W+=9Gcg58PgQ+d1>Q(A
IJ/1]5+]Og^LcS_E88N0]c#1^J]HdLA?cdH2<aI^UL46gHSTAH5f1W(L]Vg=P[&D
R0F7[VcOE5<IJAMS_;BY&O882G,-OK,,\PEDbe2?XS_eQ,?\N[LGbY3agB4I[;>@
)#eZadKUZL;,#H+38fKE8,_<LK:F\e+E7fWEGR\TF&e[YUS(OFHMF,d/LSX<,J^E
#5NY<N:^#9D?58<&g1S1]dR?5G<32bE5W:A:&0-+UIW#-K):HPT6--.0,,M1Dc)M
T@QBMT8Y9eVOMA2EDA9?^TeBW+HVP0T.K0>3O8cE>/_1:_7<5UP>\42VNE[4gC(L
ON/H];)c]\V<;c3:JC01eJ<,PQ;fPbFHY/6aGOBS]/eR@DECgM6V.]888Vc.dRBB
ZMQP6c9I[]\M3>51G0/ZSRTN45.DN@[7(3UbUgFQadS45OJE?)>a#.d7eF6:G=gb
&6Qff==Q;AUb7.^V?6cf:90H6e=AFJ9HXSW1g_E2YS:D&=UNO>U;f,Ua7<J;ICP6
SAW8XHLK[^3#c)-WYA0)M.Me9d3PF8NgIO3U&]4^-VAa+;dF<\15VU2A8LA:0;D\
9W7M8B?+e8:eCY(,KRCUE=0=N1a#YQ1Q]Z-5@>I\CfV^[SQ)A)UGcK.N#]5C#)Oa
A#gb-a,=H5((<XbPa96D&TN2=M./IEK-Ae.=PHc6MBTR>])OC7f8&\F-7H^O7OJ2
C<3X>BV9dc-Y(:g8ASe=++>cMYCe\eH-U?0VI;TA1aZ4T6N7_1#5.U41Rc+)L\.8
2Y.FB_76NN^02d(dGDF\7#T6^YB+EfPXS4=@G2HUATV:[;b7#;6fA&YDG#YGG.,S
cRgBVWKEdC8S+N\Y]cH)9>d2T8fU=EfPLDRF3HHb;D[+JMRYbO9(&7I];=Z7d4,g
;&:R]2:1_FR^&(B);&^96-e;VWCL;D\XUTV.aBU^?2,_e-d1fN\=34^E3C9DRZB6
<(+H8[==(@@@e5>S#LP\gKd7,JL_#^UN,V+gJDYDcc5@Z2gQB4R^]J7&dRR:U[V+
ab96L<T@N\6Fd(aCN)J/._@J1@HN)D0=PKUZf9,GR#KDQf?QWEg-_OEb0TR;6Kd5
YHQ9X=8e/_LV3Q1N,L7EbgO-Je+C=PdeE\M<O,_=9^CEO8#a54M9-CE-C]<^?9=;
\a97)7^3Z//?0E1UB0Mf2#>)Q2+80)A/8[#X.R7E\9;]<2QWO6ZQWF9f/d0/#4W]
c&?DQ9E#b/U[UAV?8eEK57LG5N+\<N)XL7P:a1,?I2\H5)H6^BfP0<Q_Y[9T7ZKJ
]QV@M(JDRb0-7@/EC2VOZYAY+=8e7bQ6?&BJ,P^JR78BZU_R38:3dGbQ/\^V+9\-
A4#I#XWR(]OFeY31U92=\D[V&,e)NHCc&MDMN^SdEI[Q0Da\F<3HN;&cS-3FBP+a
:P+D9,ePR5+cO@48AA_a@gZ0ZBSCUNegH^K<XeSEJI6020)@cdCXZ&^+WVK\ML</
S.bG27D&bT,U/4-THZae\?JA.^#&J_Xcb680UP\GF49GP@:V:U]XZY.1Q1/d<6AP
+d9N,g&ZAXIBf,aTIIf6e5?\7+&OFf5TSC)UTEY@D4&W)XZ_2KK@I5CB<>ET0V+a
HVg\78e?d\)e23L]dT(RfIBE>@6b0EDcNDSX;a9>QUUJ?VM[WWgbdLFMLX.-ZdSK
.XKaX7BS-7AP749H,g1AOID,a<PM7S6<fNK8++6O9:QeFK6(6+BC)f&[=73R/g6O
\(.P6WJ6HRDQ_?>NN_FCQe3aF/e#\6PgdAg7^fU^5dMS@3)#VPP&aHb>._,UI;Z4
9#eMG^A,-5.\)c0f7&(Ded^#YV)K[Z3/A7PgC<.e@M88(CHba<9KL]a]WQ7UR6Z(
,XG<@C?YH3TF<-=2.ZK<^S#3dEgN[+BI.RaB-ZS561Y>;+4RID.:E:FeXU#f<302
T]VHa=@U&eX>9I^-E>2F;-/K;9TD.5O#[LUSFRP7bB]LUUL&#KO\P?\7:DNfFc,#
]^8CCe9U@:=dS^IJ_>WLE&c[VB^1HZ4^)2;e=g=gEN]FL>aT,9EG4a71Ac8)J#eG
YP(+B)b]dLYXG/(1@9Q+W7/\&M^UEb6DIW-T:]__eg4bF:=0N\[K6IH\D4_3fKe^
FZdC[68;0X1SN^2]=/f+M^<[OV=R[[E-+,^^O>:?bT\bA0S5gE)MGe<D+ef3AGcg
\UPW^8PGXST_6TJ^LR9=Zgb5O?3/M;W,,7cQM^IB1)dRL\E@T?OP9\&@Y,F+#P^_
CP@)WSfG^(W[Y8X@0KL>U\-E]=&=GDN73IVYYgBZJ7H&2TeCMA:b99>R-^?WVBHg
VXU71^Ac#RRL7P]VMHC-VPWAP8O5F3H,2<Jc9-<dT#2f5@E^\3T/[N#6+4L=dWGR
63R9^T@SE@(V5/^?EgX1UAQL3)5d;&]f?S6MWX<fg6,4Q)(Q#6_D:<4)\W40D&:.
QcMNYRZ\@UM-3^@;5-eG6&SU[HPU0=S9MMT<NP3&c8)-?GR?1CCI>V/Y.NJE3,ZU
[FHR2cJfA,b#,:gc)C716>b_Ofg4^I-E(;@E]b-D&gQfgDOCgOCf;[ceOVUc1S_M
9R+eVX8dLXY:;]+0Y=>)IREgV3D5ZRM\.N9,^;@a8\KbL@EQ<V1Xc;D1I0d3XW2=
3K&2<_]c#@[4]0415VB)<:[.]\VA5XEF(<IZEU?\;L>LH)61OC#N(fX2Gfe:02=<
P@)G_S>PNKOS73AQ_:BKUGgR3C6]G29F2GGT?K#?F^G7C6@R\C2]:Me_()B\Q4QB
#2GE;LHS+9LT;W7SW=+/E)0^b#LG99d)fXbY2+EFXXb+)2RI?X30HSBIP-U&7VKT
&ecYYF;B6R5ZcESXH5SKIQW0b9UP(a5Y=<WDW1X8))]7.336U#>Z?3AV4+g&G4&=
M_2WM@AIV4bL0PS490@c3LM>MaY;gcD<?IO2_\.[?X&Tfa_5CB9;A@/.9\XJBW]M
U:4K<BaG<P02agGTf7BZ.76^-ZaYd-5f[bG6W?JX^;ZTC9T5ZFc,aD;=-MS)Q#.=
>:-(caR273a16Xee.:X1&4(YCVQ:2#/KEJ[dK4Ng+]9-5FUgBb4[U2b<aN6>)\\D
;1ECabWWbCbMH13.NV-gT<#T?c93+VWV2#CY>V.6S-^4C1_DGO_S]/J3G>/-J1Uf
a=bWCFg&P1Zc=bV<G0LA_=5(B@)0eR08)5J=b[,O\5fF>M\A66=,X0\L&:>d<II)
H7HgE+F^,9E1\>6/MfEaeAgZU(\P;)cg&_&V5.J>2^<57?=eD#<,Y@9JYP99RSWZ
(F&T[;/J5E/0EY(=)I^:?g5>CZ<^SOZKNWB<+HSZO2N>0LE0E6O9A:gc>&R2gcTU
dLY^D<+37fR494Yb9Y[],8+-,R&M>(\e#,YVa#fVC82\e\F4M_2M7D//-@^GU-9a
LF4-87UV?D&MfeFA?J/Z?W4(D)F1-1Q9@VfJ(-B1b.J_=>^9\=O3O+T(gC?c[KLe
IUHZLGO,AfG\K3Z)B1^>],B]FL+)/QaG#Hc.9\ZW)1@#+Q:#;6O@e13?]X4+VF_>
;PW?F:>#&Y4)Ic-G?Ka[;8K+C#<>bD1NJ[6L3U#[IcV:(RM7cCPcN5L75@1dA-0;
@0+bfC),(XJ4E6VgFL+/2G?f4_KHV().IIEG+Wf@#D675Ze+Abga],,LBOP=XMC0
FDaUS5OI3P1fGA-KTT=YPXOE4>[3<C)\8)IO1UY)V6f83g()IcXY,9U7/,&KT,gO
T2P)9c/)\-M[\1e=QLPg]NcafS.8F8PE2.?FfT<Hecd.@21:7IfS?/E3g/OdNc>P
b?X>dG8HJXZ1<P5(PKG]Y9fcB<J_P0Ag0e<KRQJfD)R.TL@;TX)::=N8F+a7;6ON
e(CCK_270(K.Ug+^2^&S#)4K_9@d.WcD?-e09JdER-2WK97^]F2=]5U&b4KD&@1G
Te3:cD0(\;<6TId^cf&(?&[#WGS4g23_D#>g^d)V@28<UA-?DPS=a.XPCVCKI:[-
9UZ>HP_I4IPMc(Jb6ES0\>A8-KA76DKZb6/]c4U#ABL)c3-F)ecVVQ)Z]/#I2Kd[
R[+a^52YA/1O:)D)(_#,>Q:cPQN_R1S4_EgB774>c6V;6NJH0dQFE-3e:_2P)8-<
He>.:eE)^+]a^?M=2:?5;0cGVVVObRBUA6)PZgZ\OMG:48Ja>B4FTU5@+S#ZdcM4
CAdHX@E/[]H8R?Qd5Zd35U\R\N:_e-MdfREe1)eNEE),8g]3PJag[NTN862g]Q+e
>AGfeQ^[N_3818OVA[++G=U]RbIg..(RA)/&]?\22;T/M=f=L?UN?2D5fCKCNL=)
d\R#HO<g&.<#AB@BNPQ1fFJN#a_A>?/^+R:K-]7T8U5C+V5:U->>F2G.TNg9/@FC
(9e5VeDZ_L@]44FX&2[SE?OdO3#d:\]eD5IKU?MG5?e4P,_gRIMaPQ#TfC6)-GMa
VfZNQ,P_5F@)\.SdE?RE/I:ECDI,(C]S<#8N)@9R+<KPPJEXb3#3.JRa>7Q.)Q_4
:SG=QXN==#H8cJe;)21G^L>K<[aF_IPBJQ;KEOfR;D1>H_U+LgDHH9@_0;MXJ]4-
07NR;J5K^e9&fT)3P5GEaLF@W?6NJRdf\:><#OR^N-bT)EJE3@QD?;YHc^6O?R39
4fe^]6Q?\A_C=9N2Bf19DKI>#fcK^+NZ.B-;V+<Zda87cTO[QF;JSRQ>8f>^f_G-
K<QdWRLXVLba7TANY#6cTQ;g8bfe^a>>6:3]a/:+WP3&8L1);FMQdEc7:)L)1XeH
L/()@?Fc0>5Dc9E2X5aHc-D24X61@849ac6;gD=N57,.+eVRV+-D6fY=.gH0=Y7?
@FL>0_\X+[V-8PS<<Z4J^)\gK324QV<LQ#WJU>ge#77;8\K.B&X>d(YfD-5:C/?5
R;;<7L2--0Q^TZ:GcgH7B:6KaBX3/#Q\]#N7+DCZ?_,]gcLR&4bO=JT6ZbM(]A)Z
N?1EBd;+^-2)92)BFA=96UICfWE1NY6[MQ:19\C]O2ZZ]K>d(;QUbU((=(\e@GNP
J-)UE1042K-,STR1VN/I5]F]7bRG9]:8M;6aagH>IWFI).M\&=7_@\@>67QFg4BO
\&<]H&>/-9DPE4aXb<EDY(S&KU\ZbDRQ<eI?<<M#eKH&+X,Wb3,\T20eB+I5=)AE
JF78_<I1b&3&QG^PFe+Z/M^:AC;]F;T@X?-aMY?CYaLe\KT\Vdf2#,EF0AR<-aDe
E;-eK^Xdb=3fYM[.=]f\]g+KT5,T0-W]fTDORM)+:XeRME2Z--^8.4fRY3D8>\Fb
H2N994(])g53U>)F609GOdb(V&-bTT5FPCAQFC-4,fIV(OEO;__f?.,2&I+L[G)#
6.V(<?&f:(0U#^Xc#;G@+F??MEIUba>f\f/.ECQXFg8@eV9-UQc@^+.aTL=PSCIf
0d^UP?H_?].ON-K-<RIMaK6ZXf+/QMGOMOUPX.[;QAJE]6K[LQ3WE?g?4]?7F?@S
PN6aT23GWIK^N\EYJT1-?5GS;4XYQ;Yf?Tg5GC>A0)D(93;1U+QD&57ORX#,&BK,
]>7cb09>@Hd+9MHf([/V/FKUWQFMYBCY\36M[eXGEF.8#:Z;);J<N6LSV8_X#3:1
f,/]-7T1T_MN(3ITeS0&WQ1=H;EG_Ia105=#YO\H2WP;>RJ:.gF3V@?5f4UZ+K84
@F)S@938;(Nf>R?:X1d(Y\T-^S.-<7:c7cN1IJ-=0S88J-?T0(g<12gH(WA8;Y/7
c>?+,(&W.KcM&-^E2ZS^Ia/4Y8BSXW5<7807IF>8cM)\O<Y#J#)@OKR>6TI6F0&U
FOA6V2PB6?_)THg3/O7O_)KLB?2=cbA<ZT,0P\cX/X+)()L0GERLBQe#7gH/D:?c
>N3(DMU:4T-V>ZHH[\^,JG.QI)E6:^gFFBHT>5(]13ACe&)5S3FFLdZ:918.Qg@(
BF^9BT&Bf-DY>:c9ZL#9@QUKcBMM5KN#MET,WIAcW7BO1F\,P,QUUA?BP4>EfDe5
(b=cH=QYC<GVQa.Y,?^<HKJHB;&Dd@3&X]fTYUY5TEBC3R<^V6M9ee)ef2Q11_ZN
7&J/B:Z9=I0;^>O^8fD,C);H5\Q76GUZ<#)EJTQc6R:EP0CXEM?gM&dSE<MJgTJ7
IE.?e^?AUfbaTM-THedJG:-TGIG\KFXVc4(b.MJ,,QWZARgP5Z,2-.;/IK-\-0[F
6NBCE;05c_E+U^CXWVHN;>L2D#2KLY;d1,>_]L.O+6,@/GcOd#XG>JWMLLQ_-aXc
Nf4&f-UIfL[9faXOK7A2.e8N@N?T6KR(/FB2/cP3SP4&KS,dQP_ZBbIcV)CN5]0B
?6B4Qa.<LX##Q6DdS6=fQ&b^[BLP=Cb=)e<P8YY##e(0X8AWMR?##O]6GLL8ZgI^
=6?WV-BLc\a.]@bd=[##DBeKU],NDH8&)5F6D(ID9QcU,.1.I08U=JR>QM:JD04-
eeF)6faZ>Y+fg[5,.#QHHL/(BaN.LEgW>RL[_>)Hc#FB;d0/9R&8Pb/@:0V1;--H
YG23FXL\I;+SZa)K#)A&(SgYP&</2TVNT7TT_LF,KKbE4SL[5]_PE1g,]LTD?>F[
LF4aF^<V:VSGX;FOZRG]cJ+M]>2^CC.CaDC-(P2a^_Q;S1^/af#DRZBPQQ<4O(Hg
])@@Y]QEA3/,g?Sf7PBEdS_U,/+gcD_<&--QA9Ac.@M.dL__J2[&0b@TdJ2LP?5W
53[f(P&,ZY5UF<8:C4?+[;=&2IfX2aWU8X#AUYZ4;P<C,M^87c.a1J_cXZ]UK?YE
d2#:+B=<1??aD\IV1_AXB[^S?c(1Zg,/e/(KWf)ETPUJ53PX74UEE#\:@,:g/SFA
NDf[dO)K^fZ9501HL549<]M/P5-7)N1M4U;&,F<=KE5UM^7@>RUeUIRcV+=6J)2D
7gKb?ZF4SaA0[3NEIRSD+O)6,O=(6K6YZaS_g8TC?LJR\G@^(Q]Q0-+LfCE3&KWb
[U7).f:7B&8R]RIbI[0^bP,PGU^@,(9/ffB#I#Sd;>0Jc<CWTdX(Ma)-KbL1=RY#
Dd1KF7@aU6(+Qd]SUR7<1G>0=+c@<8H1#d2/c(AE+;->,-T#Vb.fMd3JU(4#7Y_W
Z.2;=b83;126X.#6I/2@/CD>+BEe8=E7C7VF,<=IKEVO0I]BD+]XUc[f265OA8?D
(aPUM.^/0+(e<R.Ec2Y4SZ0:A9aCRZBd&B^GP1C8V9DC1PSQ_?UbD[#CT/X=Zg4c
HVYD+f,^B[ENdZ0>V^CT27RKKZ8bK0L>UKKF82(bNF?bA^)dbK3W(NRD[:@Ka,Lg
_GERIL)OXL.U<P(U^+f\^@^:V^&24)[^9^\PI86NS)2)1f[]X0)Oc@=5GY;:gCa&
bFX8Bf.GP/RE&bdG<ZbWAY=<2?c5NS.[<eS/\)\f8aJTA4P8faA5Hd36N5V#[L>6
RT4M)CJFJL9Q^H>1YH0M,CSHgfL]Y+V;1FbG+f]EO7D(/e-W<;E=)_:S.:T]M?#:
TKcB.:))9B]Q<D5P^TU2:72(1EIe3(\J\OXDDGe5D?+P.Q^ZZI(716?9)(]\\JWY
/.8-DAKCK_fFOcdQXA?I-cX+11V_7.Q46VL?NK[45L?;P\,.a:>dT,8H_.5A;EVD
\G0QYc&@edIER<cUC6S1a5W3:7aa>F7=#<\Yd2:8K=.RRXG^A+gNJC-8aT#,S_Y<
+a3,e>EGSaJF?N.()>dX_Z_)=DdBPb/75BN,J0,.E]c;g0_92CF:1D:/ET@e[d]Q
SOc1CHZg+\I6W]QG09V=_;J\PVaH0QBD[;/H(HYU>8H55VMcNbS0)L67?E7f1cSY
4E@D3SO&2f0&M<CIF:_8=d.Zd<If=3VR4R>@]-aGF/NYbRT)2.(UQ6>):4W922;)
QA4BSdA)AI]()Y3cSWH9_>aPL1ER3<#M=V((ASZ?AZAIY?UJ&<>F-+>a5+Rdd2H+
dP.W_=+cI<Q0-H)(9[#W[=66eDd8LOW,+R0+&5#]1d1Xb4ZDb)C1bD]J4G?YeJ75
I^0,dgQRIc5PFYHgHJ./U-Rc-gX4C#RX+?E0]PLgNQ4)I.C:0SW;E5f?:LYaTTd7
7=FO?ZAd5<Vf_3PQ=8FHI)_dS/VM>d3)?__H\N&:_f_H6/LRB#a)3;3,e1df3A<P
O48-SVAgQ4TSXd58V2TH/0Z4.Oa-]U;T<HE<9Z++?NT)V.)\[3cg-/AINX0Ca>f7
K.0E9-eL4?]LDfH:A9OfEW;J5g]<7f>,7UGVO\VADd@<\6BBCX^70>.9]e#<A+5)
QbaRNJ[AT.5TGfG#?/JIJ@3YVSf=H3(R;bR]N42I>[SO;U2M\5fTM3(5&^UH7a(&
B9?:B1=_<@g9:^@@U]be3/dK[#V#fabHG\L86Jd5H2g>Y62CPL(WV;C,?IB6E-W7
YgL7KLX?@8V&Y)JARME@AH=UK#UP4a-a/7.6_?3OWLP>DA\9Z6=>H1/-Z,LK8NZ2
E#0V4HPb8DM^OL1ENJH/SG?DdQY61Rae2I=T4JJH]C:)He&.aC-^A&]SUAW0+Gd@
U8MaC?cT?MIL7;_0K+e(M^S=WTZF7E]C>IRfc.bO44=6XPQ<=Ob]?79M82F<>+cM
)/\I,&e&G8>d--(J#_FTg;A(:W>DVBV?NL7L_\,Q-L<N1=<d[<NfI35Mf1#GYK+_
PK)QR,d45cA5NgeT4@SB\/J#XD,PX?U3QMB6\-LKX(XJBP^4GL1A?,?+be4J:&N&
[UL7cE<B([b\>0JTWc.8f[[_&8V=Za9I(1aFLOX?/J#TR)70F:F?DI&=E7_^WM-5
#VR#[bSG:NAXC18YeME]L\]8&G3T6MN.bV3V,_GdEB;E]TXZ0GJ]T\W(a.4X7+8>
)17//g+=,J,TSZWVKJ(1KKE(W,K@-MDAHD;^7.1]g;U/S0-@gX(5gb0M=#F9Lb2V
9K:Z<4KY5(cE<V0P&SL6O(?B50bK@Z3&W<BB46e^WV1\E<J?T[g=X?VG@+BR.V]D
Kb^C16S(ELeQT6F?453d94OF.E,NCW4a1J194/]JXCP/KfFAS>Ae=bEcQW(CW-a(
6e@e3]-5T)6,E<9)CgA_Z4E?Q4_cMH:I4CcEV+YB&]2377a;P)DJ_O(W<E(EVUe:
Y+72LUZ^]<63,UC8W20+VKE<Q2+^3L_V^3cf]P?;]4-1.Ua7#8;5=F?EA-4QV-,L
EL8-;N&C#KeX3Q;MT0(G.^TF,XU)(?NZfI@MES6L-06BQR[d__7?4;5&/6SKY1)T
^R>ERQga:3I-X,#T>4K=Y16G;(IeP=+M#-O8O67R7)]6;U39g<34OYXZC.&c49N1
C&]>gT/f?2]8>bZe28EY1G(_aU>d(RdSYY,D;a6.Y[&d9[P66#[Q6^SO<WL0eR1Q
Z5;SA>K(<c?JXU.gRQ@P/XdNL(JIL:T9+O8;>E&d?8YE6eWF/42MBMVF(:ddM9QH
;S,J@#R@La2=J1>+TH+3\@]e.RbAYRdN/)U(.[NW&BCXf:c;5\OS;(f;]RbJa[P7
0X4]6+c]93S@#\-SLgYGEbc>]TA:Yf\BDPE3#6MF1?TU)>d^2H7J2aUfdM(VD@a:
NdAX:VeCB649^-,XfM:R:3L+Dc2)8[f1?[R[O.FaRZWF0#9/=4W8AX./XZCZJ05=
/Kb8^H/aXNPWb[-g^&2C>VIZbc+>UcQ-WEUP(;Y02I8COQ>C?a,DX&0QOKXVZJ,K
]C^f)badJfCHS_fGZHT#UFS^#EMc;SSQ6eEU>g/#3OWKNA(:_>-@SLNAa^2VEMS(
A@?O.<Jbc@NN27C=5#/dUa:/S0Eee#J&DG68V0=G:Y(1S0IP,Y:@DWLCD.\A@(MO
:>\J[]1<[6#ZgZK_6caN>UQY-^:X:cVM-P.Bd&)RN\UAC[9<1CMSIVT<5=e?e]W)
3&(QdPd:O=M>+AOb/)acEQO1#ZIUc)aFBV/J?6g)X#<&+^F:>Y2e#1]\aY-G_-X2
E5..0S9H>H_6P@0PLRHZI-&MU8M,_\=\U&.,5U0#A[X7V6AS),34D=UV7U&S1&<[
US_]OO&WPg;#aG.51cBH,A.cc1>)N))B,G0E<KS:HCaFSMDD8<U=??TN5S[.(gA=
)A)L?.@5WgUI)?M_Cd347S+89c6JKLFE5(>)J_WC1g1Z5GN9Fa>:7XRTAFaI-=A-
N<Y4XSXKQWL_^@NLI)b/cMdbPRNV;)[AZ4S5g>1MX@<VR@GW#Y5<V\7cB]>NG1<E
RN9b[F;THN()GC\UB@3:3&>X?+KB4S)71c??_STd8g>CVCV_BMZJREVS&JG@>VEG
@[225LN[^CCPU4JF2\4Bfb:[J=AbZ]]\LQF8/OQ\OT(_FN^VKd7>K@=#.J8NJD^e
.LW7@b-_[M-9\dJ:effJ>;^DK^XOC^=a(>Mf^?<PMIf7&Cb3;AV[[A5JCcf#&gOT
H_IPH=T2dba2U,(XCVBUO:A;?7ZQRZE3WML[<FfP+4YF26[A[>6b[Z#fC2]GZ55Z
1EJ(^;76H7B,VRYc.7,?QSVJXYMJCG.>GbM8+S+\BC??;5ZgQS92N6BY6\-8C27/
8@7_UY;YI82;]aZWBPO[=<,_XP>^@6-U_(75[Id^[_#KT+_;@WV^>FaKD<ZR5[,#
@N7;,b9MWT2FS0V.YAM\JUf(dE_5a.MMeDd2fdd75=2FY<J,<62+S2/b]9TQU::_
Dd,OEV8-0Fa]ZePfH1-K\FP5X=O?E,]8/,J=H5JFb)>#cA.7AeH+fO@+3,eJ+->O
1J(/066fP#5A:ON/Y7<NN\F-HF07H^.P&.\N6Z(+06;HQ?IEe&f9CB4NO?[25Oe;
gI##JY#b.7//J1S:NZ_\CK1,SZ6&603DT2SaB9A69gO&?[PP?:4/#?D/=2PVA#J(
aY?7T>;\GfX-0.;7SD#=^3T3]MQI=D@WB]3B(HUIc3C-W(1,F4;bVb(DS>b,G/Q9
c_gG+gNd&dTR5CbDAK)e;Xa1>6-^XN^8dP]_&]D25Z5VXfC\fR)-.[fD-f,IYN58
cC][>EZZ<>42Y690[#]cc1BJbbQFaNAN]LE(GFRgQJZT.E@?^QJ_Sa?-RTCc6?_A
T:WM8Z&^W#K-]8#?D743)7K0\S5<K&C2;-<AK@fNbaJQWa@e_O)527,PSQ4&OMJC
P3RCTe&E4]d27NMc=9c8\&Jd-J^3@,)V@&G6Z)W\T1A<-Xf9MZR6QEA:_^c;DY[6
8QA27^^Y,KY]J;Abg),7[:AcX/>C>X44@EbPQG;[]O6bdBXO[,@4N29Q[#<&XH\X
V^(6Wd2bB3f>.DJX\CF0SR1G;3=g7D2dLJ;BFGKL@890H3680EB^;#V[MEAT_e7>
&)3N2gD+>&=]20KaMd+^Wbd).E)=d@IcL]ILU,A=;BbX4KG]SHH@Ef4PZ/.:AZ/>
@_4a[EAE\7OV8,f4QA6VGA-cd_D4-HFMe?-PB2_H^:-D//W@MFg.&<-7LB/Z71MX
=Q#CT6QWT=g/RZa--7@O,A3R_Z],PR/B<KW0aY][GZG]]SD@NVW?5&?TJTKOWM7#
DY#Xc2b/,eCBP7P9,A;:fF;^B[<EFRT05U89>LJG@Rd>;\7:RXD(9MbN,L:TURXb
LeaZ\XT]H8WYWI)FV\7AY[BaZ/SMOY=c#dJ[b1?J[?<_S5;NZ&&E/G1-E58H5I;2
D8IJP8Q1U31E&eSf/.(@OXO@((YNM_a/\VM[IH/?;;SE2](7XOB3MD+]fc93[T@1
dVI>4LY::RR.-R.RZ-R\F5Gb6YYN^ce1eaca+#GeI?(A9SHe:0G8?/PM0VJDU3d+
IL(0=ZbH]K-<I[BTA=2#^V\MLg)^]AW8?25RO+1.=@QHWbFeZgKD/+60T/,gTDAB
7^c7_CAVbDVVF6ZSb;PZKS7T1fgRC:\A:&&&-H.[7>gQQ;BW,(73T4>9FL&\AGAD
R7=;=<T77Ya:PXPU-\QDM(U+_\Lb_-4)YEF=BXO7A#2&dA&CZH:)88d86+O<OF>,
<aJP@,.;7G(U@Ba_EM;C]cbP<([0H&WeHRW<5V0\G2^<ARME6@8\@P7BR;T<?a84
.JbE=YUY?Ze<)#M+DPBXP9FRF8VJNF,F6?AWXW#Kdd4aAD]VN_]B:^ND+2QM9,RU
/2GXG[_NKg#O.-,^DG(]7^1#[N02Fc_SdfcJ4PTd&1C(;cAc#P:fJTG-V?[b28\&
b4AJ.D);9MHaG0^Ee2,C>1f/-P;AW5bdKgaXBLJ97P@69GRZ-J92MKM>)-&YMdH#
gLU)d6Rc;ZL:d_W;][:2:I.HUWXAXN-4a;1(3UTW:eIb?=LH+;T9GI=2Ga@:/_H#
UJ_Y?K325^;2Q5;d=7PU=4#?d\X8X(VO/4(AF_\Y9[T@(R=]M/4K#ZK[#cASUb;c
\Fg<b-fe&JQ<fUNU>b9IUM>?c>Ee3)d(-b0g84EVBY_gbcA63V(1;5#N07P^bISP
+dLT=75dRX)3Ta[5_JW:gd==N2IR3_b3WH&cV3)61Y_FT7\QC;,S[NSW,ObG0-5-
A:R#Q<(.aQgP#WW+8LeA9.O@0f22PI9-3O._EEAJ(NC8;.ZWE6-+AJ#+);bO-71)
.SOY;?FfRJa)_72+2YWF/8[O6O89D7N#QQ55]U]?LdS^6D>NHGQOe>[SGRP[BFK^
S;_0[L<5NL#C:4QJ>I:4[);^XXF&:PD5>6WQTXDd:Abc#&QHdS?L&]:EL6;a^_Zd
I:T:V+FCWZ)cf1X^NKZ@21;d8H<+Vb&S;\2R6PJM[Q;-:e>Hb,(FFe)1@Gg)0@fN
V(T7AX-bb:gJ)UU#W[)A;;.6WfM(\IM6:C5Sg[<8fBTJ^K]gJM9PO2IDITgJNS8T
;ad,AMGP0^T;F?CZMIC=bd)_aFO8K5f>#fLH[P,#bS4V^QM\L08^ZWLHXCC@Ic<E
Y/6+Y;d)Z@.]c9dG73bDV^BUH_^X=JNBZRS?2XC-8P18RK3:Z1fgH9g5Uc-^4W\_
fF\)/5D^-0.e16?17P-\I1UAgYUS/O(GW>1U6#6cfZTI>3e[\P\S4IHBVB-dI@_?
b#_HcVEO=&Q(95WN/_XK].TT(9[H_#D?1VD#>EIcNHbA6IH<f17GWKM6HMX6CT):
83L?bNVBG=39T3?UBXQ_0fX5_GSUMaG[c2[@AV0#@.gPEWU:;\Ie6<TVS[@LB@_H
=;?W=OV];=EAKJQ^g:CfK9b\\HWZDP+@WGC<Q),fLDX+G?RSRJY7?4.eIAXBFJ]:
1;[Z3LPL@H+WG5TcE0P\R8Ag:fKQ>:55&eLZ9NWF)J/EgEW+W0Ef/ZAEagcT;4-I
\[<;7RYfGZ]EM#CJZbFJ+dF7^,V+V4:3&3O?g;GT^SfS>#679<C5c?15L1_O7c7^
db.7-OKcKX.HCXRIC#1W@MSM/\#N-W[<fcE1]#L6).Ne2+gGWDcH-a]PQ]cA_U&/
MK@>=ZTQF-8D9A-(2ZeVK<1-B(46KFHD2=O?SI3:7>3P5[-_<K>&eW\aXa(2/b_U
T?E2KW8P8f-6bF7Ke(>TV9CZG]I//M_,0J;N&RSQfK)O7F1\UgQ5QG02gM3]DWS<
AG2VKH-5<O4T0T4,X.WEfH><UUMee2^OcCV(TVN/,4)N001?4-MR7WPMD3/>U/^d
>,H]<15A1LNHC&V_0#>:R)0L6)Y>&RGZ777(P?=]:H\Y6HG</SY^&GW)QCZ4/6#A
]KWF,F<bDFSOE]eY6bTA=VgZMGP_,UK4=7M1SKFV1[U0U81:.ad65ND8FTWO\?#D
@T=b1c0_<PJ#DPde=/VRd^SfEJ<1,[D5T<Q?84=9&&e2ND8TbeX<OQ?Ue#RFQ7c)
\bI^017FO:OQ12F2>(_Q;b6.[D#0GEag?IQe>+VcWSRJDeb,\U]-.7AC+#2WF29#
:g&e;^YR4fIG?H,KPBGYXVDQ+O?c3;a#6PI0#9AF^4P+;3<;YC\bC>+e\5CH_J;;
0bKNDe&IRVI2c^2?Bc6d>FHN\FF(GN,2BER\WVQXOe3Qc^)VNJP8NHGO_1^W026=
AgT60d,<e&.e\G@Fg)>-MWBgP0ab^Y>2fW_/@Wd;cN5[2W2aP[:PEg#(-KH-R\N\
GegBQ67=+X[a(Wg#IQ<0PESSEZ(?aD[B/4XN1J2[aCD7#]Q.X1HERT=^FIHg+](0
7P2bd)Z?L_@:3PHTLK8b9[@6WP5TV.b]?b.3>;8;<0BdBST>>S=0E3E=5fT]K)T6
X(CIXQ\IO^DBEe7Q-ZP0W=1U#I?[a(LG665A7d07G6\T:D?IaAY&8JDMH&X4f+G4
-<Y=5P&e5a_1D4KgO#V\8N]S_QHb_?M:6.A\BQcO>&R3O_?PBNSIZ5a-D^E+LK:L
BZ3C,A\/+^=QbM+2,=a3#>MXcC/Q6]Ga3;3^7d:K&[O.PQ3OX.D=f2VZdI(=KOY=
A24/)]#-D[9gaS@V;7#H.>>:N=3aYEOVgUX?]/;e2&#9_Cc,G5bIY9VC]84BfSOW
<):\;J[<17;SQ:/_gX8:1[:26EdI1G=5eX+H#/e-M@N_#UZ-#^5aMXce,H+;7^d<
P(B-:R/5OXE#;DG4JV+Q+e21bP+I5:5DX-gY)g6^6bZEeJ;?21-45?R#=1>PMUL#
D8EMT-?Pbg]Y0)=Zf05FAG#P99cL2BDKEZ3J.HAB#9TZ/8a=[S,C1&[edY5URJVE
AP;-BEVE:K1=?IPZf:&VV10W0?DF\VPI6T,7Q3]/]e-f6U4OZXgD7Xa:>9T&K#Y5
8A^\X#\+a6@KI?_J<LRA,H/)<8=ZSf^d6ZcZ.#8cR@2^VVP8PXU0ES\IUSbD6C/d
^\XPgW+dC,5FTJRG=ZZ83DPbJZcKc3Od<_T>15B/_gM#/MDGL4\A7<J=QReD^SFV
^W77IHOc7INGFO+@>FV9PZJT5gB(^b.^b+3&=&#e2N^.),eO>b^3TD8Cb4?@ca61
9/HPQ2TW(Eb^80GD3QWaBfCH;-Y#,D8OD^Z]@>#@7N3D-+YSP0-:.PgCUO[2aDE1
88]J<8Y49\OBS,RMbAO^<a(e]:P8H8#Y]fbQ9<dLY8OUN2+Ub@IQJ\QGgfa_^DB/
5M:K0ZFCD(,[LXDb&R@X.NF0QKHS1Ib;/MVC<==X9DJ>4G5X9(5Kf;;QPVY9.M(?
9BL6caNG,cF)&GfX8d<(2e-N5(\;&?\QX=2;8WORSVe]F03.XYSI-YK>dbFIM&K0
4bMg&B<SMO2GK4\ASZ,XM;aRb>PA3)P?DIAbFB2H1\^e\WG;+.g7)4\-@;1#b3&,
-fYIOW<,(41\#>C:?3\O@KOPH8K-YPf=MN@Q+T;#_0cBR>>dT&+1d>0UQ9)=54+g
3cC=,e.abBb=^0([CV,-+^J2PPCW\@^IJW,H(>H_KU]:JQ]E@F(&5+8[X^^(K;Ma
8&N2]X4(O=T1M+b=_<DM1\Z[B]3E7Y(^b(aD5A5Z#gB-Kd]XNKO;a\_\LEa..J<D
<9?8bZ@XL8]=e58)V:>d/e;L@7E&64J,+f;RG;A(<0[EOJDZSZWc6;[fF.X^=1>g
9[+BVMXQPLBa9RFI#KZD>bEOFEOO^-fM8E8/VV+<eOL)e0A;(4Z42aS#3;_U@2C_
+.gU\+WQDGS9.E>&g?#39.Gef.0RYY.SYD9Fd\.]M>VUcX(75,XQJTHO7R+=POe<
TZ&4D<2aNO+><VS:S+1)P\SGND9eRe5ZJS@EcQ2:8PEK-L.RgaL(bC\-[J6Z>GTM
I3e?\[I:K&F(X@,.IFb;XUd#I^L>T].IS4/EcZ;U;&?K<P98N[G))_P<D5HUDdde
C:@S&&=P;M@XcHO<M0NP[(X4.ERaT1f1@)d?cX[=]Z.NEK,=B8_c2E]IOFIAF3T<
GRe7LZDPTFVf#OJBaU6),[H7d.7d;aXd/I&RXdF:X+/Zf?0?=L,RSKY+A[IbIJ+>
&J\.[__[R.X/+YS]d-]D^bUa9,3HLT9T(LLa?8>]94NGe,#J[aNB_L#DKK&X7YNM
dH209D.4c.<cO(Xd7)L<C@,g749e63e,9He,TTg?>>edJ64&5ac&-(^GIg]C_Pa?
[_=_4+RIdAB\,bKdY?9&N;HZH71GafJ\<E#:gIK8&L&Vdf26-8(^fO;VRF=C3YG/
HH;+dfGN0JT-4(&54_;[(8D+^0g26e+1.YM?[3.ELX@3bU@e/^G-AY\W^K^O9Q.E
0<9TgJ8MYNYPO9Mc9=PHC,Xa/P8]_0J8H0J34ZP:FN<+&NY+eR826GU,B)+0<7US
3NT[5C4-8(QD=(.XTaX#C1R)2b5@aD,(e50>>O\\?.7L_8UGDO)GdaHgGH\<(QaL
A@FK9,#TZK+:OBEeXfY-^d8A3.E\(Dfg-g;GF\61@OMFY\O6b=6D741WaJe:\JF(
bLZUeXcF()6DNQ[G-OI#.Q9@U3?9PVNQP<9>e8Jb0Sc+ML^SXgU)dYK7^e:8<)R0
+H]Cb9Kg2?I(9C13A,G,8ag7CSR,XeeR?^&^\GK(<?JgV;b?14T5@A4IL+J2<0b?
YNA51H_X1G(PJH\IdG[bAI;NIcVX:DT:#)Y+;C439<e1b?MgVPKRCHYH.HM@a;RM
8aYTI>/O<eKWVBPFPB]A;@57e]:O<\[d91BY\O>@JJB],&6ZNJ;H5TaA@9&1(,)+
D[6H\^EB#Od0=:Rc\C]#XRU3)77:T0cH#Rf;ACYVa;[K7Uedfg]S1(-VG7XT:.b<
[43YTJ9e#9EPE5f^SE#;KG#@_8@VK3FBHP:\e@0fFEW.X@06BcN?\@CN4+NgPBCP
O.L@TS5C2IJ,=ae(WG[:K[9:Z0#6ZbQ=WDUER0@G>2eX=#[;^X_@S\OW,Hf[VC6U
Qa8N,43DNFb6P;MFJ4.K#e,Aa3CP:0^WcF\;3?])Tg,Y\>1XR>)Z.PaXU.gC7:&g
>UD[a:Gd:NgFGL/A+SbcS^K>:@-L#,#R;02&4X44V9aPdW9W)L&1(]8NQ-1(-b;O
?JOV+e.KggE(@9g;aJR0Ra)0b2TNg-N+Rg@I27DZf-WSaUa]N=aDe_c9N6E:)@[E
?G<2[2WQ^TE7c[WB<B07eT:9Ie1D46H?bd,#XGBf&WfF:+;:aT/7J,f9b@;>N7Qf
?HXO-6d044YOSZ.Z32_N>G0?&:3-[AVc8H0XFX8PaD<eE\>KL1<1N97cJ#e,I/N0
Ce?ZZ3]T^>[&8CQ=(/J&5;,OJ=f+HBCQ1M;G)@^Y^SOb99PH010-D=OF7;8SND2M
;43E\WVGRK2e1:5N2YZXQS<^Q59Q13RO].>aC<957>@T4gf^OZ1&JL,UYd@0OWTS
c.G[]6[_(A:1=eC#B&B[V7Wd=OgG;[2/[E#K1XSNPVEGTILC8.S.@/9TK<[.<JX<
9XL.2&JC\S9GEGAW5Fg?&83KYXZR-NaMOV@RM61O:#&CB7SGbK41IFBYNL(7:P:O
cI]d>bXT@AV74_gH+]FH?W7IDC4<g0HWX03bgc.fWZa(+IJ//?Q^e.C^4^B11JCQ
9&;#d#a##EI\Y?eYg^Be,DR/15IYL34ZZ71)2#d6S(+4?YM:[1R9.(1J5cAcY@MG
b72;+,HW&\5QadaIAZ:FSKT+;U#a286D<(PO&?5/-G>c>;K_>F5dgB;0,_SEA>O@
#0.Na3TgHL[RXa^TMd[8/)0+HVeMY-[N9?8JTE0U3E:2<6R:a36E.N&_SaQ:+]82
J_dfA56?4#VWd)GUaJcW[Ma29+dfQ@<Yb=:]IFJFE<&AD)S]BZ@8eb2I12N-]UN^
7>+dYN[F;6cB2(ZEE:Be[LR)0BBX^_c/VNIdL1(<DZS0X@g1JHc@K)c?e\eGbf78
?(([&S82\-=SJgYY(@PU#baB5C,R1GAg3S5GHV/]ODfA.^66eI/]:I2.:D2aOSX4
F3HW^1XAF-_9T1\G(?,a2ELd.EP#_><dZ+c]eFH/)Cb&2[9QbDG=^=e-4L&MRK<d
K#G?<#D/;Q]_WWEc<^O0P/-]\OSB7FgJZ;dRPR8^,G7IHg;5>:KK?DfQ(W:6]0>)
G3B8I_HX,[?eDJZ:VX+>RaUb.CW0.VTP+Ef5Oa9>(G/E/e7C\WF0B&aEDB.FcfNJ
/F[HF-<ML])?@ML,UV+;U2)W(c1Y/WU-L/QN9F,C1],(?]A&GJfGO+@HU?O-.\=d
M<Z^=9A4-1,UdI;Xe/M,4IKBULNV91[<F#]9K=(1Q41_A(B73FJ3ac=FA,e\H-:-
YHV^G7\H>2>#YVWM6@31Y=?M4;UEK3FE_.0/dX<(^)JG.f-@[8#W^V^?D]WP[2S?
C.05(aA>^JHJe54PAO(aRfe@&,?2W3AFd7babI-Q6([8<3FL-BNQ34>?UA5I8]e1
TYdCUU5@I@Kd:de@7Ze>=JXf@>32f:R.2UTeWWfJ5<-CJ+_UGA3a#gL98M1Ka43G
_DD64Df1YgG,RebbfK(c<g+=V3cC9PQ[Z+AbHG+K9^++AV>CF)P3c>#94:UV2M,^
5^B[]JC4dP<LA94CSIVJFTMd=\2F]aN:0gP^fST=752E0-6b:P<Md43,_\9-;F=V
4D03_1c3QcJU0b]Y)HfW_U0695&?IWM(BW[@5LFHQ[QTF@/R/;B[;3B7,EQ+>S@<
9WBeVCRbHF78+V#S&E0)>E(>0gXf=JFfe6@.-+^cZXSE]g;?>5RXZQB_)-=S]A<)
g4W\M4N4b]Jc)PQ8UQ2?U?_1GO>TG_#BB2M];M2dFU23<N@NFDM^AOE>+dG?aRPQ
#)41RN7S140_^@,6_KA24K+0PR.HVO;Hg)e[404NSA0HG(d05FE_#M.W+,b[KUcW
RTc(>VL;C0^OE)OXIX)G#BKJP@3#_:#b=_d5DJI)\W=[c78&X--D/I4I&H&aSFQ_
L.H.Ib<=HW3FAD)[b8R2H?D8L6L#e<a0CQ)A=:7.1O(8^+[#M-4\CTG9dGBJ?LA0
OOUf:T[\702@ZK>5EbPfN#8f&P)68Mf1-3ga19NQ)cXC_c+-=T=ZI<f.\^P3@.H?
A5b_V]P@6]1B>VGH-M[J_bM^AE7V1]X5&8&#TW<e9\=[(DcA@+Xg&WQ#JR0LEC0I
7LQ5:dc9^&,1R_P>,KL>?M28J-@._<O5ON85DK)f5fZO=AUd;bfe^7BOQKgD1EfQ
8OU,Qg_D;gecI;4?gVPSgcB&#FT^]PUE+\JH5g2QUTD@KE7H(A]/BNF#J8-NO6H&
ZGT2M8BLIZX<UFC@O?I-_^KZVN>5I=DK@5.<3&>,1R@TO\7D^R29FV<D.CaPHVC[
-J+)D&2]V,a=/)dd9D1/ND\WWB_8U=@@</^(B/8<-488:P\]&JV@K(QVTS?>=BT)
Mb^=?XT)I.5C_M]0JRO.98F7d)#&IU(<6-^YE97;6VZ@ff:?gZ8Y-_,JNLMc+#\W
3SV2b:b7C?IH5cRNJHP#5&UIfI5S@>\,DI&WQ32:OJ:WdcJ&1)1XE:EaNB8?)cTf
BN05b4>gWP;[S5_JCRV@\?M/->:-J^O#M2W;3ZQPWXGH\I;8/2Q<VfJGMZW:GF#H
H;d]U@3(8[M6/0JIB2:/WZ&d6AI8&(J49N8&I,2Me?6V>cc\_5HL^a>[XQTMK3>+
<aJ?ZPRYc\PJ_CWS_M>:7.TD6KLTKLFQMR#(bRL=C8O28H_@GAC9:&L]_OEd85O?
@J=g;05e6gY-+K9]-7G/SX,FGRU+.3W,H(ML2L-[/CFJ@c[H_b_PcEA2P<6MC2Z5
V:?^0YB(E4I:d-)ZT@a56A1:HeH/KIc:(V?\\aJ<e9V7+Zc/U]UL>+.TDIC^;<GH
4DNV;VQA#b5aUJcIK0]:^H+U,:L0;6GBTMDK(b;\O->e/EE]B@CMSLeQKZG_cTdN
[RgO0EU=\(H[)bU8;Q05)&V.#P4^-4HLBHM-gaY9:3W(7NFA2C@KZ>>EFa\XPbET
Z(WUe5R89[N]:&LYaNe^O,:@_JZg&C6NL2,2fE4#b#9e_GUCXJ[CBOVK9fAPc=cD
S.c-@0S=SfC&3^^Z>1R2MP&88)gf>ZJQU\bTOY480?,<:EIdI\T>\/^T:7LAN=TM
X;aSE<8S,V\XUC4A8UZG6.MDHBX3JV+64XSW>&Q(936\6fKVNJBWZ3(_8@ba8deb
6f<RVG9[MZb;cPSK2.)bId0Qe/2U1?0WgL\-c,8WUYS&I@0e>a+DITB)O@?/b[-)
(VV=N1W_P2bI8Q(Fc+\F<)N3)^;EEHDH;7[&.:3FB2XOR=?L4g/MZ4d&8E9(YL+\
X6>;H@WL_FJHDSIEFa?J2f6O7f?e8BcNLJ(8I,aO:cZ;g(cA9cBY@QIX?gR7ZI;B
AAMRW,f?+W]W2LJ#5D_d?8?ddI:L8=P53YOF^f9[5bUdFF:3;-[^GY1HF[H-<8^&
L2H^dFc\=7.4&ce_XYa7J+N(W&)_e.EQ1EX:f64)J54NOYe7?-WT[H)VQ)/.L7?Z
g>>RG;Y7#V]eW_bT0Ja>K^AEK(D+2KIaN&XPSU8A(bd5@HI[@\dA8TQ+dX+b-b^7
JTILHDO:XN@6[S/R&U)b-(HaH4IE@_#MNIg?(bS].?N_(UQP\)SM)X2(McV4fV2e
K6R\I8O,NH.YLVbFOH8/R-JY;Pb;ZC<[/)10N#7\BH-[_^):./XN6M4UP2JY86J:
a(ed_,MV]H[,\YV\<[.d,dBU/e10N9J9]3]E0^^.e)PB;3gWO8Tf)HAOPQ_O]5J>
.FL:=]B:3?A0KDMbg6O]6f>=.=Rc:CZ[#H+HQUV-NQ<KDdY+X6AM@U@6-#/=-R<8
[0d>\6bJS9?a,X.#JeI>Lf6eL7[Y9HWL.L+6JJCXbcF/cf5/CK5c#eOf-Y3I:a94
SEN,6?5UJSUb-X4-\-b_<c_g+X14AA:b]F=R5R=F+,?OU:NVc;7N9UC],)ObWd7=
<a,[X=e9ELeG3PQZF@#ZVe)WDR3?e1@+bOY7BP>,+UC1;W@D-PSQb[DU+=RH5\df
TgeUD36QL]g-G_?f25bU5<#:bc,?0_7))c@2JJd[V57@8T0;+cd6D2V8=,d2^HLX
,WO^1#-?eB8G#6V3HedcO/S85QYe0(I0<68LNKY:#8)?(/.QI6,=9cTSe]I+ZfDM
45\W<_+#494ea9;BN0DI@,.F&5M9H&AUQU;P(C1^LI5@PLI8eO&GdQ)FH12<eYcB
TQJ/AXL2PQFYKcP:DZb4IJ]ec0):HCKBY,42[9+feEKKF\g<0DV[d57>:e^GJ3/U
<g[],/MBLL]75c<?PGS)=P9LI:9GD/^#.]/0NU^5T3B^<1C3PU(P=H+H_N>^OS92
3I-UaB0.7c976L<B[1R\4]g9\1?=+a1E7H64?P.GNP\U.QfA,^ODdWBP88F0]FMf
/RPE.@9\)7?YK9f9e.bNBKC]1G18.+>(1IRG?5Q;UfEQ<B4E.><_2;JAIgLSZGN0
6cJ1@&])L:6-;aII3UXEVKEGW7P]LWS/(gS&.+[c,/,;(,O4e,;bdNTTYV?G,[]a
ODUa<TaJN:/JXLF4]+;-2aJ?;?,988+A<M.#LY&F+_A]bgDOYJ>IQ-eX-U<58M<R
Rg6HKNP5ZfRYI8CbJg[f4f>&VdVU.XW3YKR]e1J1f;QY5R+XY)d^]@]Hd/:A\=VY
,#)e<U,TKI)M(2,8<EYIBd(ENV3:f];0._9JHP.EUFL+S:WaQ,5gf0T,3\&&]Y.,
JY,L5073B4fL@4K,/5E@W=-5[LKF9B>1HfTa//58>=[feK7C#CG4IG4525GcB&L2
V8+ACL@[3FN6KULd(\)O=bIFI1fHD)N==YSW[[JJ)GgY;=a<M[ed8S#M[D[^F]<O
bS@0c;36@-_\@6:MdAIKDd0Z[A,V35Nb3?gC7V3b4f:][bTaRddCRb_W8#MgW99_
^R2@K=DSLYbgcA&Ef.1cX&.8T&^SZ0+afR;@</XQLQ(X6)8aQ(-eD7D5BP8ELX<c
GgMg<[TB#3_>\LSX3/5daE0UW=YJMXYD_98ZBT;I[4U/V9LdOd-Q(5=7V^U13=(K
)R?U[a\ZG,&8K&HI;;33L\]/KJa2/OB#\a[&VUKMKY4dTNUU[;c_,9[H;08NeC,F
GLL?b?@EC;FeR@UA;Q=cVP,ZJ\aV()/Ve)_9DJ?2N@ZgUZ&@45S;#HIZ:@e32P6M
^S_BIA,b.YI.UeX>A@9EJU#2bM&Gd(PRf4EKBE4^.O)]#Wae?@LM:BOZGP^FZ4g5
?X,0&R3E;&d4,Id1.-Q,IEKRK:A6:G4IE,R-Hf@:5Z)gV:,J.7^ZcJ[LEBd4^X,.
<d>;[]<TRG]2ff@):(KeRI<;-)2RS/<UF<9FUb6AEV<_EWG=e.W;Z,6O.3\.H3(,
UU6BLP)BO36NA=]Y>]DOA/.+83.dK>YDVU[C_Y,&5G5GPDFMB\gJV,2A(.(S/>)1
HgYLIAd+36+VLI@.2Y,1:b0N-9=P2QM]R\E90&I)SN:24JKVG4=00[X@.LSOHD?2
)ZCW+CQNNNA?[#adI\Z)AXg)ZedLBU]O]/\EKb(e#UV1/MSde:,L;S=RNMeH)I@L
UE(K=4\)I/>@#9-[c>#ZKGeZ@6;7F<RBa(c)#eJ=bM@+U8^L]OceAY\dG#^H=SXJ
e5eW)T_&\[03BEFS#ZT\WU9K)1K>DV[T8eY&M7Ug-:dV4M.IHP[/fKTE1Q1<U@;9
RdZB,4&)+^6U_<L/>CWJ&HX7F-9J#f;VBe6/0O9K_P,]g(YVCO7Pb@SL@<^,5A1K
[=SUeK[(7W?5+RcQMQ#(D9=-<97XR5]d.FbC1_G-GO#4GF.C7TWRQaBE^0EKM>-7
84.7;&4fd4?eKPg/e\8M@Z#L(.8BFdK[:YE[#bbbPCN1.P:8)@0F.OVB6:;A4X>1
Hf2_2\:dVaUa]g&W=/a?WA4d28D.aTSc<J67eN;2C>b+C+b1DHZZEU?NZ=)_e4N;
VG0#QbEd\@BM]T,O)R.Sd0/aZ^F>-VL>D^:]4cTJ6FP=D#F^L.UYAM14aKbHLW<2
SU5PH&UdaG(+f_NUZc1.M?=Z38[[.:=K8@PH(TYAc0KY1>FMfNGDQ,/:,7MN50BQ
@X\TCP:YXI;V?c]VI/43L5&Ea878A<a[Lbce+-Z:ZfZc[D\JPG&cGYaRL+@PZL8R
@XM2#6:Xd2#4UUHWb8)a1WB\&?8]6,e4^#X)P8I\>7_AaVXC#eGO@Rf43JIL4Ne1
/f7:6c/8#WK>^]8S?_AI3F3UbYg&]SA9:FgB&Dd&=O-]N^Vf3KI<VB0_FafYKKe#
SAI(dZ9E8NL<U@-fN=NPGP2P8g[I6Z5QMBMOEJA#+0S+XK7O+\:-J/8S5OCOL]XQ
ASAS-:B(a#Z#TGZRcB[T-]J-Z-<Yf^_:1N)gU(g-#R?E--GX8V?5gGG3VCC=:/D6
GN9E+0N.aZQ#[S524e(K((<Wf&G@cF43?dE+0UDE7:#-#^0Qa5]dAJM]<]7f7,CJ
:X@F3&9HI(?8?@7EMS9Y5dEP9]:]P(B8BYU;-C0V+\PC<@GW4TWO^K[[@BHG6XA+
1,-M\[VgU(,9P+;G?[FE1\^bX&1LPH4RUSXg4:Hf(G8F_IV/gN:(R[WSPa]/X._G
W@f3XT]AWgOb)X)G86^YdXda,W9&P#670;WeER[fUH^RWR@A(FVb4VddV_UT/Cd0
P4XM0NOS)WFK1KZ0Fc?YU?[\-,gXJI&P,[d)e]J2KB=<KI)FGFK1G#S=:-_UF=cG
Lb9,0g#-YY(:,\f;TBeP7HUKVZCgXRCLB(##TCU<;9ga#X\g0d\VeVXGQJd?)JAV
4?_aX4U-8gAI<[(EI<g0W[LF&C6;/N_N]BcT/2EQBO1BR0)II&TK4=T=dGNI[gY)
@^_(7C\L_2?g-666a\g>#ge/9\N6KMC\9)GWaKG_7E;-9VJ/G]S<dgV+@J6:IL(C
^KQ#@\784-3>K#/0Gg6O1>FaOYgD1B(R+SJS=TK[A.9f&cI[WJYg/DfNRBYQM6?E
H+b/Z852B9<53[a/5;/44[9Z7Zc,Q)G-(/<5PFU]_d^-U4=C2)1PM;:YRR.:8-V5
DgJII)V(SUgL<;C.FTd=IZcD-ZN;<Db5-K[5@U8Y,TK;X@AJOf7(W^#7Vd76JSN7
0+M??0F#,.Ed4+c+R51,E/3+DJ0SKS:E8WQaV8ID1@a#aRQBIcE:HBUA@UB;>(1f
eZKE<dA+5_N)UZJaYA==Cc1gEUD>P5A1,3:]>g27gY\2UM>[6#N,)S0YY_G]95YI
[QOO5ER&>^8bQFAPU4JNb((=)5DH:\6GX]2dCPfEAV(6PIL-GPc81VI_4d@Y?=5f
7XYW+A2LJ>aR&=a_.7Va-eEF,(G158R)J<+aS5Y_P,[fc-^G@+X[F<.H4ZY(H^#:
1DT&+;g/BbGCbRNP>^agCIg-JQ4S0+.CaL6BVeRgQJ?&&FYT<FJ^c4L(Z;&MD?e7
+:6/IS4GROZcQ26_MISS@##=3_XK?>QQ:(#B^]3R8(7=9DHP#V;O-+1@=#X1]Q(=
,<b5TVWGRV7Y98,BOe/08ZA5EO(JN;b02]U>/2>;BY]YAG#->:B2>#dJ5RA8)T-:
72G;d>YM+_U-WF/_:95/P>23QTSHERIWd^S;?dQIKZW=fQUPWY:=BE_+IN-)gBJ-
O[c&BU&6<V5>=TQbQ@W]9.fP2]IW-98#3B@014;:35&X,=5cg<Y]5?_5,<@e6T#/
;\fdK_.Td_.ecXe6fcBN2#f&W\X3]:QVXN^\X0CT=&Y-,Z27IXAUU+F4F;2cO51?
G^F;=&B7:07->.,]53Q64M^Db4\TF<#A6P@S-V3LQ5B\fbVD&@D8/E5/[&(X1J^;
9b>#P&9(R#-@-Z7,4XY5Z?D0\GI4;)D#G>S1+f9,UEN6.V7=SS\1dcT[)2DY;abc
aGRVFIZW:ILIAbA?N8:f5@-fZ4RU4:?OT]OWGKTcgQQF>:Dbb6X,+1bggGW>dYZD
0Cd019<e#:;3<g4=8R4)c(7VVgY1Z-Y5c[&N,03@U]g>Xe=SG[D]Af?T51+6F-VM
@N-cJ+\2fIU(aB\XYbb69ONG4R.>/354@/9J)^_>.K=SK93/)MWT.#fQ\?9,/377
5D#.D1:A,IT])cIaac-9dMfGdDMc2SW@_M1K?IX3OfX6NM+D[+?QSQC-R8/Pge8&
HZQ7W3>DG8+,8/BQHP[f;d^QMCR>OWGD=?#fOd\3VH\Y.Tg@aCU2V5;Y@K5T,AFL
5(=G2(3W/<f[8W0;CDf@1J+:WJL4[-3I>M&aLgRQYZR7O&X&ZYe+f]dFH=g41<C.
^Y_])He2IL1YSITaS;.[6K0[AMF_MO#<9WB#4.[_,]7K2TB<_M;-Eg]&]VR#[J.F
1XQV&5ZSXNQ)QT7S8N5JM6U[Of19+JJBb(0B88-1<f),XbDMc^/6K4YRM@#D@(eZ
]:8DFG<(U4I\GU:=P1aecU]T0E/N>#,>a78\GDeR8G31<&SE(@/cJU4W6@1b)^,E
921KWSNDH[-1Z:C/+4Z=Y)XU-B/O7QTU14/C0f8(BC+)NOO&7,5F&Q8-HD=eL&29
+d?A:;P=)c1BSYW_.PdI?\2I8Z;7g_/2R95-)H4\>&P_J[^]V?:8J1C,g[8P6CEF
&\ECYbeAbAJe[SfPT]R754U6f=IU66IRHM-e1aJSO(8E1:3b?+_a;a.G1K=7-+-V
1_H4f>O]3+4M<]S>#;8]bdNT,G0W?.&^]1T=X\>g7-bV=>ZF)/U^[^NaBAPAg)9+
W>7H-QJd4NV0=XHg6#]=FH/Ha[-(.+G)-4I7_OdCO7.E05)0JH4e5JSM_8D+d\[e
,]&=P[;;g/;M-CFU6(;7fB\(2,G<=?I(Da/>aFI7MT]cQJ?ac@4C#:]@bd9.@VA\
Z;P7E2fJ/S[BE<P4a5=46@D/86@EPHBV.VD(T:ME@^C016N8c?^YgKO@&7J=RJI<
BGY&\78E0AbcKL97SOU<A7)Of)3fA7J/:AHY--BZGdCXPD.2(R^ZW>0@b^A4LVQ^
1G.5.IJ>CXHUY:;GV9JW=^KgNK(:;L(L1[bIQC8K:BebQ:,&dD,HO?DXd54[W7Fa
DG9#7V[CfDTT&.<M5TgWd1&X4gDe[2eb68T2;]eT9b9aWbO.:S3bf(Wd@[LDI#9#
HR=2(^W9?\a:9a3H2^:(;T_5[HKELHL@(M)_aW-85?Of0)U/XFQQ^K?.V-:4)=Pd
5F[VPg\UT\=YGHWJ5;aA9;>5:3c-2f_OF2J:TR<eJdPE&Z8a_H)RW196\O/[)\+Z
I280RBZTEA98(g[@Y/b)8F<2;#UHEI\N2&Z6&UPOJD8c8F;97[8,]RG)9WeP+.OW
B@P7/@<Ta-UFQ5c8ZX&X=26E9A;RcWMVQeVL10T_C]YS\NOC50:e]a?MgG?JX_cV
9K(N8IN^2e-4bC63N0UPS74J+LODR258d7<.,SA@K+R]U?(EW;O,@FPb_XGG>dMP
TTgD+_ERFFe)(NHSf9_5Qg/.R^SEgF>MZfC@,K4HR?cCW:-;(cJ/gTa,S8C_0#W]
PPgUI=HgY@W)#=KbW43SW+(XJ/V_LNcARE^.Y[UdM[=]2?<\##B(&I&P@0D1U^_T
g?M#/E18,D^deM5@,PN0Fb>aJ9+U&ZPW77.4<TJ3BH&_46GNPH:110d[MBXZ./_G
I6<=UWS0;CCSP9Z:ae#4OW9Z9e9G<BU9aZcbG\?MXJ7>,aaE2\^U-XDB):eHKRQ;
80g>W#2R1QRgdV:5[2c@J[=fCX6gHbS4L=OF=7d1ABQXbHa3PJ[9JZ2<d->4.N+2
7Ud,b[3-;0H:H1+W@K31J>4]5\N15?UGSF65f1[+;e[cT-WVY;EI(SR1.gC,E5(3
V2[-OCRfLUE6-f7DQF]@352T6gB)9S]?J?D+@CD&B4EJYMQ:c(,Y@=]5b4RDEM71
1QX5]\72\\2=0AIKLRO=3W(Z).e3JM&fReCES]?.U;M1C/d<3U..B;]5JWe5U8J9
WccB_9[X,fD(#/?PI[X1-.OTMNfJS24MLB^#eg)1/\LAbY+H?^3M^TLNN<;ZYaA0
F3;8I/D=RD[V#HF].I>4F^NaUOE,>BA#7,+/Q).Z;0SA\DUaOBM&LQ@,UG?E0?61
,f:8TL]Z<\a?g[Jc.HR^0-29=DAX;#:6b=QPd2W^XCPUf#g@2gYQS=&V-J-6(Mf.
V&a[KU4-&b9>LV(Z9PaG6],N&CR2&/9YJeLMa-DL#[:IOB&5K/)F8AKW(SDABdf9
bOY16ReG.S^a\5CcPQ&#/GW;M@Lf?H3(&P+]UR46LY8+eDP/f/)c6a01-b64:Y+?
Nf/YVUUe-DLe3SK-TMLHN#M47DUACVFTO)U[G]@5KP?=J@?;740L\#+:O?#>C8;S
6fV:&&Z-P(a3IO7+MLTDADf?L^\SJ6I<)&dac09(QNH\QaFPTR41+aR5J?[;?FFb
W&3@WF4;,;+#08G)ec,OO>VM1_:/_>ZP((&7^DG;<.N6a@K9Q=OL];ge_Q:=+VEf
G@=.W\2=_IY=91)ffUAG8U<X3P;;^,Z5_1ee-)7:ONaWTFXHUTKHe&F2+g/;+e<V
L);YA.c]VTI,XRX6T,[&83+3+0]cUd971<YK1B=bH4YS8bJ#d):RJ8)<dS7P.D1&
8c6_E4]8aYgcbY6,8L@?6R,H<+VMYE#+P5L//gb1:+6gT[g83/25F&g=LNTNVQdN
f/H1-3YE8(/1;cXX7,7;&N=R@3LGYf<>6/bBb8Q611.T+>@ZCG5cRMfF3R5JCL5@
1FF/W<]a90-7@R\U66DfFfBOM65.__]@[YBDBf>XWZ7WD@;dV=Z)8P1M-3:-a/54
E4[ccOIT^^6<-15T<Q1HAcA2a?[AEf<KMKGG?+])fJ0Z182@=-d<7d/S.@OV?L)Z
2-(0#@bK^c)XHI>0AX3:4DX_e(-EW>f.,ZV_<0B7MK)eKUMGI:E9LS>(>Q#K.,^A
cR&:J-(e:@2bCQcKK6FAUE^[C&_=VdF7cJ_NW2&Y>d7,28R7IK0VFScR3VLbQ0]#
9E2X:_4SXBNVPNHeG65Q;XKf-B(&:+;F_GO>B-Q&(.4DI@[@:(4\T^GB@[@TR)FC
INSS\bdU[\B8-8CfE6eE?6HWM(CV02E?&K_S-5=<OK(I&?XY\:ga7A;5AQ0gUX2#
9=>\.d:E_].c&@F#:a,IZ7>0N:&G->/_RIdd?Y&XWH#X0LG_WLd=1e/CTf.]>YfP
7BdO5aIAUYONSZOX@aO^V<-##:g5C,TYIQX]c_b\_aUO\<BINFaTS8W@9Z#A)GaU
OecK@W5ZWfA:fJW:FCQ3FW]0FV][F=A63OMZO[EgZ@N\JR#J<J73ccV/7>^Z1B7P
cg#c:2bLHMPZSg15S0T_\E11QJ.MJ<TWc;9J^WFAL8W&\<(/3<;c(LXB^@096-<Q
UEV,IV+7.M;&Lce&^ET>T8VR[YQIZLaS@7(AQ?N:H=OI1(bgJ_=X)/-(YC/T4\]H
(e9e^-9S=<FXaFJA7/.:Z2EPTFI6?ga5]a?)faBIH/V)\L5(@@,UbNDX+J4CE@E<
.H-8#a?@N2cZ>F?6Kf6,HU;=E6F>RL#&)J5g]&daIT[PP?3f4+&[M>aDS3McY/W+
O;][)6NLR)OBJH]9.627UbH138:0&^#-?a7XQWa<<QJ^\^.BLFI;Q)0eWF;-LU9.
>68OC_VH6B]KLdB/S(S;Z6N@)ac(98F6R.8T^2^Y1Ke:^3PAD&g&#-CC.V@&S]Z\
QMF\a:2^U#-/[H1[Z5XKRKH2Q5b)KG5EVZJFJ2g7C5:bV+3&Z.@PCCSb?-,,e?SV
b^Q)G4--)[dbgQRL^B<2dNW0g,H2W0XJ(>^&)g-NFNAF8G650SKE]MU7;HGM)R9^
8HZ49X+-2+Od-.OBWD_bLVg322]5)gNR;^N_6f>C+@f4+5[,KFd=e7X8^H.+JIJ]
T(bGKb9E)a^N257?:QNdeTbQ;(<:Ha)<5W323MAXK_We88U6([V<;C8(8D6:Id+B
dcU<I0GOg#)YQE9<W>C^<3QF]PBOWDVAL(XgC<R/a1?R4>2(>,+DUZ?]c)#Gb^=g
VG?9B\MeHaB[]HMa[-GK?&)eb/]3+Lb,R+NUa)9bO0BN<RQC@bb<gR4gL+)3UcY<
1c8_#1R^ULD1A5XE_3SL1:JN9f6H>/I.[P(_-;;AM865@CZ?;W2^Te:);BQfa?d6
&:MSc-680WOfP,8:(e--MQb[Z3?9a[]/_O+O<U2^MVSE9.0?gcJ@;07.@=Z+\SP:
^TG6/Sc=FR5N?,<]PZ3@Y<&]ZX=Y/3]D_FPNdE2\(;I6]LNd3/Bf&-gd4]+E,d)7
(gd2[(/AN74XXO8:YFXAGV:g3be1DZ=dYW9FH\,;K:BQ9e5<?7II#\W5I=e@FJJ>
^(QD,U>JK?^MUccLZU2#RA2)1M3c_]LcIO8#S./W6,7,N:#[IH-@aB/7c,)b+9FX
?EO\[U#O0+^,^,^e&&A\PM7f#U\:(3Q6M.EFBFV.,JYBZ:_,[(<>H^<c,G82AO2I
\#E5HOB]NU\KA<d0B62bO1#G;2HW,VK^D[ae[>5d_QVbUK=4aceKJS]0C&&1]CX6
IT#XDaaSQPFAP94INNTMA5Je-_b;/efU#4F>6NP/0f@1>O+)[0.Q\QdFAdA1#,=;
5Y-;f4M0/R_&A2+M=I_bX,NIaSI5L?7U(9CZ5MH<aW/5d_NAV6W4X4IgS5ZDAV.a
1)2G\-)NF^9GX&YT,c+]GYac7W-BDg(G-_Q=7Z605UVd.M\c:,_0HE;V][gPL^fF
+6\[982LbM3W)C=eR)cLcYdRE9>06ZPVA4c/8NK-+<,=95&f=NS4HENKb91V.MM+
.2,S4C6AXYDO;O.;/,Ag5-;12f^M#a,^ND/6M7),fZ,4<;Vgb<6MV\&b,=I36,2C
T)M4g6E/-K?KO0Y=FAC260:<Bb:EVY8L5H)W3VRG4S5UL+=5PZY);70GeG#J_6SR
R@/?fXU/HAAQH/P;QXQ&c==1@#ABa=OD+2)P8=^QC8<QC_NZXXI;MUcC+REDYV]X
^f_ZXGQW&HgSVK>J0N;RPOYM<8>]R4d\(V0K7+F@AV45FO754QZ)CD639,^11JHW
RD0->XMXLZ+eU-D9dR01#N(MASXG0D@6Vd)@P=)<+<+4]&2DGV[L2C#M)\f=RdH2
PaD1E<S4Tc=W</-c]S1\<N07-L<KQ2TQ??YbVe=WRL)7,+XYe\bK;>/]A.20D\S<
)OTDM:GGW#^aM\Z7#\gL2J+=<N\>)ZA5V/6;-1E\22H(c+WN3=/0J#+&0HOB0[C\
FfC:LS3V^g/4;@f7Kc#)7WX];O?\<Rc/S8H3J46Ab=H1>YA0(^=A)I55dCdbN4[<
AgF^QM>#2C_b0ZYZf&5X&W=Q-3UF+g-TbIBKJ.^/T&11DI)O=CET\B+A.M.(fO&@
Q/fTKf[aeRg/@>O0TM8NK-E3XK:IRd6HOIF8&+4_Y=DP:=EP:V7Z9cH@F&dAK&g+
G7aP\7W-[9.K^b+.CaKW[BH91);UNd+D1\Vcb]<2dA-_PC#.BQ6+.b1#BZ2#eS1M
D/Y.YHQZb+9.deA.5Y1;0N^W,JWG<R8,TNEG^Z#O8?^&02<EJIe\a74AOL#3(GLL
U[BI_NT?^V^BH2?/AV@caZK41&>3&>VTTJf<,cMMaBPHe.SR0USAO1Z>GDc:;a@9
LFNO(P@GHY-M4_XaaE[_(BA?W2Sdb>??;?BJJe5],VbT/11:]]-XPT[.Q_<@baHg
#XdX/\XSCFGG.PDCR>3FQ<[TWGOVOG_X9QGM6A^0KYa<:ORfX4,IU3P:Pa1US<ZX
a2_dUFd7fMbE[9_\20gcL7QR3(WC4F&)JU4gd0FKY@<g8=3A4g@51P)d19JJR287
@M2C]<7J/PbR((g?\)aHVTfG=fN_6HVP+,?c(__G5ZNDS?V=>BX=T6\ZQVA_[X]N
/@D1[SWNf)9W\<7eg^4FA]X;ZB+Ug_dIN;\&#-:4adSE=&SdB?P>P?;XVUWP@g21
<gHD&20_[HL_INK7J1N1eeY-5)>>-[3:SgS:SN;;DOMCZOS]UM640dVNR)8?L6]I
&\+9e6FE</bZM#MII4LcOcO1UN.Y84DgE1K]dSP>L<U>6KQ8TXaNV>S6:XgDdUE2
45C.Y&M8_M5aCfDGJ5dV)_6&ITB>1>QaG<Q&)>M#cc@ZQ?-+>_dWNEO@H)PHZD8W
+_Y)=I<f&T2PQW,P/65^>JY)f)b@MK.=fe>T+50#_H,0+S2d2(F)=BJ=LI;-SVc-
FF;4T0LAZLc9:,2<)a^]1aBAB)^\#dfL?9H_ZCb/Q[d-M9LXa)GE\6<\-@)Z[6>-
4IO=@V@B[EVVME?NP^A6dCX-32JO/NZHZPF&N5722./7+ZA[9S35>\3-4=V6&2C.
&3eCGW]P9LQLfE.MSB0>[UP=SUK;X?)T0bPJb5QHXWXfM[WXUBFZ\B0a:GeM&4?W
BD2^A,a+B/5YLE(P[Oa,RP^3&2+d+S+Ib8N89g:CS#U#ZH\d<W8>:bN&fHJf>W_H
O<Y^d<.5Q3KJL3&g\NXcdQPHg.88>N02IaF25US+E&\FXS2@_9Z[<=J:e8#>B@Cd
@?)<\g)N?BEdEHaB>XO(g4IBM9gG93XbGUQF#<.QT5:Dd-#VP]2.QH1^Yb9K=VL7
20O-+=;GK&\6_IJNA0/?6;M+B;VZCOgB<IFBX_E^S\d.;QN^?,;-K3Q6@c:D;4NP
_g:.54-eDbZ@RdI2ea.2QU1aY3<+DBM)L<2=7\eTD5LMT/=B=KR2A6QKI0-^fYQG
;ZS#AS##?N82;Va_+GP#c2Re/c4dF_EG-b](=I#.#,&G:LRXSedKDTLc[ONRU@M<
f/9IQ<2&17N0c)+Y-RaY-Ae0eIGVdb[cAY&VadgRQ/Q5Q3H&fE7)#R6>P>a-/NgZ
;V29+F+TN[5Ca69)=]V6@G(QA,UP]21Q8ZW<b@YJB71I09bZH;EeH\#cO(V]-^a)
/-9d22KRLN47W.>NZKZbPe=a\-e4&LNI\8DFb9^QW&feQ+GJGTE4#6aOAD)2X0)Z
[c=<^#dN/#;DPMJgbcMcXW;Ib=HF?W23e&;0/4EPc-E85cY@&>+B<E2KB:.<6UZ/
N<H&)M<.LG11\UgPOE<NJ-AM1Z3;C5Xg;8V8M7<<UP^AC)WVgYUX9IDP@+PH2g-F
Z(V2(D8_T>Pg]L?1;RYFPX6Jgg?\<-+c1Ka2TU/K?d5J?;R\TN?R&;bJc?_L6d^;
2<Q,e=Bf>^=Z1GB4@0,(1W>[W>6[?;)9P^I^29e<5?/JX(.5cN2)<&V=(N0T71-D
68DAPSL4WCRdT(IMa0#N<OQBg;BYZF:,5R^0\^XYO:dYLCcJO0aR0e(/..5eJ45F
BFDWM#gIRH\&]DP0_f,<<gXUT@V])#AG3J&]6(<QGHD\RgX(0^C?4J,B1+d>U?IG
B(^4B[(^<<&C>bQA+<H6^Y>10NAN_dM+A6XJ\W/[fJ@O\aa#Y\(KR:))J5-\O(-8
Ee7;Ha&XT;ZIOH><?.B)e-OI3>)MM/:(._b[C_@]05(\@f_\c)-8FI&QfQ+AOJS6
C+[a,(NN:1T3_D-N]eUdg,3g2Z=bPa3(B)46?C9CR2]LggRg1CL#O_2&P5M5),=;
CZG:^JNL+GZXZ.?AI6]JgVg\_,?WfBDf54eJ6_&,19B7L(Obafe;Q>1a?Wb:I0E\
,G7AD]35ZTR17/g^J/T@,Ob(aTD4]f5;]H;Z/]5CI>,8D8gKU:S/#^]5GD>IB8&W
QJeTcEa1<PbLBAR7NP-+DY<3PYTe3]H@eA+GJdA4ZSON8@;PQYd61e--41Zg2I3]
ZR(D>Q2WWQ\PQ8bSTcCIfO]Rc]\^FPG33GCH2B.+,#:0aZ>ZASgMRJ7@3S8INGK[
C3X4d>7QCbgX-,^2GW4-XV>cgNOE?/-;<D0V8H&2+A&G/DC&S]HZH[fX]_ML)M>(
()?bcUYY#1#df7RdBUKI;^bZX4VRA&/83K94:]<[\-62#37+WT=_TB&]bWDQLg:f
B+X+G<b\=0=5DC=Q^^Q(EJM15GcFM.,1QA0+8[1Q^Q\6:Nf#U7&OB\=,Y<HIUNdU
>e(,))_(_N_HFTN3cNT;?<I34QdSYO[)<APW(0W)\eY7548c&a]/T#&7L5a.\7ZH
VTZ/T=3]046XeY=+X4\L9OD3RA.D+@4;#8beJ;:/H9.G0,Y>C/&.J301WcPIf<>V
6+fe_</<KTRZd4(.T1aD]T]6G5cYLeLg[dE\=ge\4Ac,]S2;eO3<V7IAO.NX:816
R;P)\)2.W(:5//RNK+d/d5_3MD94<#N,3##+bDef=H.L7HJcY0]VW.;cW8c>GB68
ZXIRAKFf2Z_^+@FAY&F<8ZE+3(5->Kb-@73Oa]L:+gH0G,QMDSGJeCVB)1<#0I7/
2RZ#AU:NG5,EZA+I9Z^bGF)O;>baDS3Vd2:2BKcH(Nd\]UAfA<Ng3XcHNXHMY+9:
#c^IGT;T/aV6&]2LP4+#aR28&#5bO#OI+68ADR4dH]FcEFX>2e[VBYDRe<#[2[4Z
L:QVS7.>/VPS8Ec0YbfW1B]GXKSJ(L9]G:1aDg6&Z83B]+/?U^<#L+2N:g+-c(Jf
RR.>J;4+KUg4I-)WR]GbG7VLC^Q^BC,A#(QMG?ZFSLMQQRf26I[Q7LC51^,;2-[U
&dJER1923d6Sf4D<Z=_#@KM&3Z;:0HgUd1O.(UfWC+6+FC[BJc6-RM;Y43#Ra,@K
_a98:,8=1HLY@b-,Q6^^K0/aEP+8>bJV<K0LWNf<?CXS579.CKSQGH3C=QgLeOZ?
+MV1F#[9YL^JKcJe4N].EIa.[g7a8C>=TK50ZacP[1aAC0)5=S@2ZJb6bKJE3/fK
D3D3LTRAO_e94D+G3aaa//;\E?R7#]7fE=gCJ(b<&@<SYEgFAN2\Sgb<aH^HVNbP
W8INV3J=3.=7])V^Zf)-OD8/UbODPX20U:=X\T(gfWN6SKa4e#@K@KR-X,bS5cB/
I&)+:HHT79=WI<Y&@5>2),7)A;.0B[ga1;&R?=QMERBJ9CKD->W\a40PaL4/W:c/
6@@SMabPLLW^-aGHRfQX7I(=_R3e:(W#+CZBRNfG9OVJO&b[=<(_IJ213R365Kf1
_Z@XcZH&5YV\JB=+K+C^(eE2[VUH(GKD;0?&-g.T..\U#g5A>bc[S5D@Vg:Le#O:
Bg?XM4XSL\.g)H(:Fab<7d7d]NKGO?>gc.VUg>28e_B/H0^+NZASJ>XadVIT]+Y]
Z+<,UN=7:S8=BX80D/=9^EV_TA+V:M8@4O_0CFPJ+ZQNMI=dWe8UBb&=0]3&#g7L
W(482DB:8#D>ZPeGAfQDQ^3KeAXBORANX4-@:dc8-SQO+\XcJW5>]MMYM-=<1XGf
)g/F5Oe;34FBDY5\\8bb^E&>UR?K\F\dC;DdK1N[LJP(_&2#-;G<SEZC9STS?&QI
E]0A,g/[^I]UCeYG<<Mb)Y:S+3S-ZU&D8?R/cf^14<A<cDYB2+N4(ed7E9cA_RX7
N6Q4bPCOgXL)^LgT].MYdH#M1PO:)aUPE=g/^EKGZ:g9Re5>1Aa8J5>JH&TcdTWL
Z3.3<f=+30PZYAL<L).?NOK<_6QfIe^e)UBJf(d5A^f=#@C:SM8]/E1>6GggZ-Qe
:3(,FgEdE@0N(gTN&dJc<[BOAAWcH[1gdC5T4T9+M(W5&>//S=GTgVRTG9Y,&\7S
Eg\f8;]]_.fG#M6#[28&)1S@X-:S]DPGW^e[OR2K(a[[9^TTA=B[B)RRPc0TFD60
\KX6<_EKee:O&@@Je&G;OfK5L;TC5)M4[FE9<WYMXd&@9I/2N==4a+S57:^@7\Pd
<I]\9D;=6SMa,;8J@dB8YT9#A#c14_)bOdc);F211Q?9C&[W#EPB4S8KfYN]Z^NC
9YM5(M-9B<,NU6PZE(BNbA94(.?,N<b;/b9Jc0dfLgJO9MCFb,fJ1V178LYANMQT
7K.gB[-5bUB>HU,c1dU#0;6\,U\A&W>[7ZMX9=S@cC&@AbcC/VP]D=6^UQdB9Gg.
PHB+S?X,SO.)MNKP<(_9>IYDGQY_VO?bQ7.G4g(.W@;S0@^dA&)<ZP_aU9-U:YE=
-1T(Z2TXZd8La<L.3_Mb,+V+&-cce3?H?,G^#c(:FX1L[KI#,;TP.9NZF7=0AeH#
.XC2bVXYX_U<0ad5?@1EV4gg>K^d]1aa:d[4)aY9&+62fN;FF-KPeWZ>-(-[-g,H
Z-I3N&6M0<X>O1JP:@<8EbZMD8>NXXX-05#J;B@cK[I8A&/GQb?@X<ga;#aH@e<S
Uf1RQA;3O2S4TQ.&MSLL7[e]=2I)DR4Cc6fd-69I4&KUOY(#;W4016MIN+^+([2+
Oe8.Te=0&#9PRaFQbPb[bHT>2:LW:L+Q/bbL[QZC.S+aSVU]6>UWQ1?A=5KRP?5G
9gI(GG\<R\]DU[E&K0a6g32+IgZ>0>c0&fPK1CAC7;0bWKXZK8PbT+5;g11E,+AC
=ZfaLOAX^Z+f^9E8M@AZD+Wb;U6E=?eQ4@0\,/g3H^YLP^Wc@-OH+07]6/@A8N[;
cPF=CFegI5?/aR=ESeY#R6OVM)S;8g4K4^edE@(]WCKe#>(A;ZYZ^Y^\QZX6gML?
&a]42ICEHKK),1[Jc>^:\Z3))OQ;bJ[Q8YDI-&c;dF((7SeZce^+&Z[4KJcO;@14
,gI86RU?9+fR0(Q8G^T-5C0^f2&c.CG(gFg0f2JRW5T<<A:gW6Y)\,_]S^S6ZY[D
/Q&WNDbc=b9QHXENQN^eG]/g-6cE-<_:>P+a0UdQ2[cbR(?.^O(SN]aP,g:_1=>E
30[>RQR2Y_N\gGe.e)@=bD1+9\,J,WY12X&N@fcZaSXeAMYLJF,P(>^:CQ=OJcV+
+S#KI94/-ZBcO>Qg:</WK19S(F.BJ#d1I5.g9;S<RV\M+KSZ?6Ie[,->8Y8^,YXB
:ZK[L1?<(dEH5g<KT7c]GR4,4V@K;g1^[T\)0DO[<WE2C7:.--M6W+UagAL2_#@:
bZaa=N,&]PTbO62EbOV(F//<OVaYH/G-/2Rd3-T/d6QQ36Q:N6PDgDK3@<;4>aeJ
A9b;QZ9RgMR31KfC>21RBQaKGa_HbUL\-5XG/L_+-H[5.V,A^HGf7,YFR9W[:5f8
I1[IX\-OJH&3/M\Y[e;2X##5T6Z/<[baT:-f;0)QD1Of79RQYbAOAV.=A^4?>JLa
bD-GA-BO+&>SR42C83DgW_\bRQHD.J3S1FRQ/d1A;ZfA?X&b(2W-8M.^>CR&U^cc
B\]6X3^g+0cY;2HP6E&T6MbgTCJc9LFINB4&Ve_+O>9D2+,>6,7aF&_c<TTCGG7#
DN9QXW16KR:2<-8^CT0RM?bE:^OU^R;Dge5PD1?/cTYZ(\,^-<Y1=O:2?KIHcG6b
?36E;RDaa-N7II=\9g>UK-FdD5cegL/[:NW43LBQ#M,KCLA2:0H2<](D+.3.YGY;
&f9U_\U<IP6-UP>NE43SP47;5YI3.\.12UbR<?N+6RKfW[S=fg?T0M8_e.6Gg3.,
>eU8+9M#2#SV)2K;G[[5DHA.SQ,PBcAC>2;)9NHK;US01BOYIE#;K/bSd#)?A\bU
9)IT/AW5G-0JWNJ&SQUc;K_1=9&-IVD62O66c-_AK]#P28ZKVMb=db.Dg\^65]VL
)\Q_FWE=3_J>bVQM/DIMV&@;]a1<]<e_DQ72^G0fB/G0=.JBGJ/DMPUS4LP?XUFT
;]eGBd(-7KVJ[?0AFfZ#Q^)BR0X&W]LD.3R>R#GdP6b6;/M-0FacK@DeL0+8E\M0
.f1-#UAUG.#a[UgAF:<(/?a6I-P+J+_0eBB/>D9IbK=[)f)GAI\g[QKH]M.T#8Ig
C]K&][JYU,>&[X&K)DFO_=EVLeD<-A\UgfOC^KY&c[BO[WW)-YZ]9//D7TRVM[^f
^4a>J7&55Y[b&83e^.)]3<#e_6JE+V;T8TKYO)K5;UML?0ZK)IN73:D2C3+&O]W9
&4_KOQB9fPD&1D=cDIXgTTN8LM_JP=?2W]]KH6?+)P39-9Q1>))e=C&4@^\FRd6E
?C=B1E8INV=BS^_DJG/NNd4aB(,=TTM^:JAbBN@O:&I.R_bC47c9b3.Bc4D2F(-/
TZ6\fBY#a#XN1CGgK;2-:c(?aea=J#(ESQZ^K0<.MG&a&.,_J+WMcfe#<<(YNEKV
;BJ?^#U8</0MaPXR4fV20(6;b3gZ.b]?XF^L5E,L2;D?:c5?3f>#0eeV@X89O5GP
GDP2-SGY\4#W1MC:>EQ@66,VX7[RWIPNFJQ+G-]=73R]MI+B/.U.612<:fT3W]fQ
M\Z:8L2F[PJB;XP=b@7<(XL0<A.d[IOD/52V;c225ZW+d_A-F7^I+08R7G>HZ[F1
db=f#^323E-<1H/P//O2-U=4<QKI;b&M;]K(P9EPHJWdN(&[_R96?>TB)6<A(e\e
G1g&LYgWU2f0RYU2WWQb<2@++a:PV),=F+#5f\e+6#1C,@SIH1\4@1F@Pebc,WX=
.\Yag?fU]ROgO>+JM[(-eJQdHJZV/V?A7LISHI9/a8M,D9<NL[[OYWQ)=>-94e;A
0b82aW]>MB_Gd038g+d@QG99]@HT0YZ&4L>9MA1W_(M>B]X-K2]HJ>6&&J,AWUPB
P(_E]WNZQ)7S\@):\Da;7cZ?a2:8R5G<:X:E4(<1J1XMG4T/1H9.4E@,>UaICVA]
U/a<86(dG7G&?XFE=K0aafX4A70HDe(5CBAR]?MK1cAL06\@8\?A^G8/RaLEQ\gB
7:).X@B0:X).2>aB=76XUVCF6dLVF9V7^d)07<J@c+^+:VBY4ND^<Ub+e_;I[-SW
H&Ab#I1943<5#GNOcJK+HC7faK:,I2[._9=M1A^CZ@^I_+<D0T]K)PB2KBR:U>O)
+gDcFM\IC;S_PL4RHgP+HGfNA5#Ig:)\7J^)&FG5=&7)bE6BUd8@O2/D>/;7;LU(
NK^N0XSI22MDIDD0:84-:3S/V(7f_B98]P7.aZQ:<G-(44RKa4N]@^N<G&[40\1.
)b9<_220TD?KU.FfZI;@-dKDR;64JNR]5C_K0cNG^cedg\4;/-g)-MUR@1\2H4OB
D^.0^(A[6\]e\[B-8AN[2>Y)A<I?R8&c<Re)<?9\EW8)F<8TSUeG6S&[T#]H7UcH
]Q7Zf,=]P/8d^U4I?9[PS.>Se49]ISdR5(<)Z/S@=41;c)eLUOCK\O?JN)M,+PI-
gGW0#X;RIJ#DeZK+1K1UcFT\S(EW01P+IW/g45g8a-aN6JCNgD,806-gRd?/:5O0
8&Q&3X;U-:-QWf0?UO3N@B&-/a+Q2P1,0_g-39Y0?bH6U1K\,8.g3:-f01@_[12#
7J/,E#J^ff?=CFYBMR@deJLHKEE)LeVgWYGR0&CUWd9AdDAbP.CH1/N\77?1bUN5
OAF?DDYQZ?eER<,TXBS]#:??+,OT\X+W3V/QCYM<TUd&=S>1,(R]+MF<#];6X<E_
O+WBJCbJUdEbDHBgOfJg22.^f/K8&TPG\VC2M?+1(6=YceW]KL(fAg62N^5W<YEM
D=S@;;AS(CaP>0O^6?U5,R<42QBKL8@:ff<Z55bLV1<]Q<a&HO,B[NYZSb5UK/@@
>OQUC7[L5^<[cM@9c,.ePNeU::9C#T:;PH53^@#EgN@@W,6N1cHN\SdB;S/.CF@)
VF</:2F^UX34I4V@:PQaD)6625_//=g92+:f(@S1TRf?:N)G0@_<B15J\IU;,;ce
PE6eNJ/b3fJ;B:&[GA)HcGV\#]6ZD<RS..F.L,d:-->4-&=b#f;84&49=)>2gEA=
]SM)=6=fM-5>9?OQWG;Q_3QQ<;T,B>#>V>/J/1dX48JQ35=5@2L8[Xd=B-?;IQF4
7S#C;b?GB42f-TGJ#D?QbcOb.ULCU>T>T^+b\6-BO03aGfW&(?]cC#7[V>WeFJ>\
AgTUT[=D?02_\5>6T\;Gd805@)fB];R07NBJY>dWMJDS>F/8^R)A;.TJYA.+G?D)
WWGEPT,ADAgV8&cKC7K@:)WME70YK>&9;a1&?25Y0<[f1;O4M^\.QQ8(#f6@N1R6
KQ\N#Ib@c(2DEUM21OfTEW_)7+A+&)7>F)NdA[e<NfGK9W?a_=)_K)D0Q8]HNWVe
JN8DOc.TDBCJ50V<<QOHGGF8B7e@cXfdGXBV/X17c_SSbR?-NDHIKa[5;:]->YVX
&SESO^I<^FL>V^Q6C.YVU;T)N]^4e^eAGTCdCAa=9S(,M,JV4TN2aWJgd76Ue8Z[
T7gIRD@2ON/BDZHYRBRFa6N?b[bTc9/UV&PIGKCSS+dV.Ac=)PLP=3Q)Z&)g_U=d
Gc:b_^\-D8<55E7+47]]B:CA.Fa9MUHK)2C6TJL;#Dd^Ig=MaX.0X()_gU=#4OH@
cO]W?3eTe#-BX0,11S2N.NDS?.5^/P6g:^(C]7J8V#THFHEdV:(d28ZJOP_.2CD&
)M/e&4Za\/BG@GMG)H[I+[QU<>9NAf,->HO;g02bO6QREeWYcI.JO6BMR[KGJbXU
6U:P=P7OJ1/#.@0eGR0H^:VeAGUPGN&?cD60g:@:S&V]._(7GPZ=62.@#I7Ybe[/
CU]=K3G^+S9SHUC;.d&,-Y\(Uf7_]Y;+c99D7g+UU1=7#=]UQD-TGb)OP)HU4-FI
)f9B;A;I]U#,DY5G?b2JJQCNbT0,^XDf,bNYA>@PY#g49)QNHR85&Mc10a]7LU?#
+D5RG.24+N]8U,^;XP,XEW+fbS.N+g([eL17g\X9#;Cg/^Za.L[^_X59WDYK?.3a
Jc5P-e+D^&7\I2)B&;+A3)Ed>[S]?bJ2L?TD+_N?9d&I_N>_PAfgdS1/#:&5d):F
cc^1(9WW,N?:g\2X;-QL>ZDaaQW=V57&WA1TXR6A/W=+&FLIZ857Hd8U#.F;M/?+
F_Ia&F)+T;Fe=0IRa:8-&OTY&??OF#V:&LTUN2&d^\b?2@FY<7=368e0PWBAT?M.
;6ONHR].U8C]eA&K\.J>ZB5c[)_eMW7(1WNY/GTCITaU@BWfP7#2_QART],>=^M3
ZaD+bU&D^;EWIR+g-?XZKE_.)EX^8._<d9]:B[gTY<F_cJfG:]cAfEE?2A_ZTHKM
9,a2KDd<cZ?F>T>=(gG[C7?@)+Of/>_5/MA#D9Q[YO;4=[H+<J[=-,&8[)9e\4KK
QbY,9aB+J52E#,Y#HM5TTOXT.K;/)(9.,Y34(HI7>LTLH/g/(KZKaFA\)06Y/bJ]
3f<]U<_+YCG)A4d+cJMaZ)/DH-H@NDKJL\e7P4UM?cLXfP2<G1YbQ@W/Cf2>63c2
LIYXRTO.6K3Sfd3(BeD^g&Y=>/SDZePVA6TCd.=ba:bLHSZQ9?XD-D6A8XT9G:G/
^69C#X>I<7Wa=/LDY1e[,-5cN@ZZEP_<RG^F\II[Xc8=\f.^JP]3(4<[4X[H.V:K
EcKD/?f?1/?G-FA6Z6,9_LQR4,b8B/QA&TDS9bC;QaafX:E26//BB)E^;&?AFEeM
)LK/_5\S5P>Ggf]?Jbc=c>;KS0<<Y=)H12HCb_+&[]^_O:]VOR5^1PZY[O/E=K[\
@PR0G=&,M_4TA1fDE#-RfXe]S:f6aAV9;R#,-4XIU5G+?9e7_H8/,I],<LTP.MD<
12FYD?JYBR&=IWE+<DGS0>3-d=F^]A(S0;N3<g)P0HM=Q>W[@/]3O)N<b#R1Ke_Y
Pe0XS//DJ9+e/d)4(7DgeO&2g^MEHK<\74I&GW)>O4:8e8F<O_9#FfN=Kg@,(/#b
K&c&eQ2^<cfGgZ8)Dg64e&AREQ<GK^K2M0I+V:.U4_+\H#<RK[ZYMbc=?JEYDg9b
UbU_;L]IYU_H_<(6Y+ac:R7PPBL8:7&5Y)?:=f0C.I8cEWf,[2V-9a;.g#KD8FTE
Q2=C;dPKd<K[cR@PAY-MGWF1GPK)LZK@LX)#fD4@J,5V6M3b^,/-0U.aY-;_3X18
UK7dMO3KTQb/ca&^.(OVf5R)>U8,;3##KS>3Sg#G[>RHV[beJ2::O4II>L3e#f3.
^EG+c06-3.Q2CZeGge-03PZ=VU@2f;^KPM)3CI?N\(B/)2T<PdY;5Me#XL6OXX)c
#6cV:YAJYb=RN4474.Y=6=+I2Wd;O6OUcIc(0WOD8)R&TbUAKQH&DCRaKc<]eEUL
[R35b]FFD<NW,N5)EUID<Z#BBYK:FS^9=<JB..fJ&02/8+U,YY#RME3)??)Nb0[_
T5>QfQ7G8Wd+I-OI[eC77F2W^/2>=2?7/;a[fSPA;HfcYZ&d7G@O0>3\,[?Y<-WD
f/\VJ28M97Q?]N;_UbR9(7>aUMSP,XB95F+B\c0f(RRgb1MUT[CM[5R<OY?_YUH9
QC\6c,(:>3J&H-]C]E\=\fP0:/4F6YQUB#)<65-R)U1AQPFbI_D0<g,H/C3JI@9D
gdK^U1K9-B&?2<?K1I>@0@I]3X6V_b4W3/B-RW4B^@),2f0\J-)38,U<J_DGS\W/
02F<1_Ec4^3N7;QG.7HX?1@T[+IeTVOTF98X0L9fGQ;b^6ZE_.941O<g+>K6<J]#
GU;7aTK;/BDa>#N91G-FC4<gf0H_I?O=?e\AZ4IPXAB_e/Z5:HP\.17R_ee^b:+[
4:EXSbT0O6Z]_a^Rb>cEeWV8-W>ZSN>Sb8O_,CN@;XZ_1R?^O_M=8,Q#eW+DDWJa
gU)AXf=A\9f;/:X<3D=6>Hg_bHJ2-00B.+e(?IO,?VR5M[ObI^-)19->FccUJRSO
^:UPY5U]e+&0NW^)F7a(_S2_FI3QF04C:>FR4F]8(+X<X,U;U,?A6VU;KAd_<bAO
E&SQQgFdVF8YB0LIZ2674X,)I^Z^aA(a]MffT4cOFJI/AY]+ceQPf(;>#_F9[\4=
M\F4bZF?]Sg&XaZ)C[#)#]eY;Y^2Z.<,B/Z-AA]RIabM1<6KB510a^]f[eU-S^Rd
a(T+;Z]6W=R[[CLN2Z:HHX==DOcI+U<c9I8SY2VAO77CFFJQ_ZN<?Zc]ePDL-5)\
TJ[Z>d;5I57[BL-5FJT?+4fe5[RK:SEW_0a5+/6D8<^YMJQ]caGfd0]L1+)NL4RZ
[@.Y7QY:NF2Y_A>XR8d)U&,W:3&]-ZIIWVBHK)6OCP,XfSW-3EITQ[ZK&E)[;O;-
WO@MgZKDO(UD1]MEK8C>DPQ(?]aS2eAO-(Q-0O2eJ)W]:[C+RE=:[<5^[,27\P6-
HJ^D//><AC7BM.C1f-B1c\<VdJ?=Y4Za\2eDZ]<K_;F>((XOZLg8QQ,=YHL#>?-E
FX-37AS<JW9#<ef1X?QQNGO9SFO]>I32LU53aKaJ18XCd6NWQH/8.:&WLa2._F,0
Y,@[_A0QV_I=7/a.;J3X?La]8<fER3<#:/0WIE0./U2A^WRK+B4.]Z?L1Z#R@cAU
JCO1<I@C+[)eOLWa/HRV).W1Fd9<aH\Z8@P1]68<6<3^]=UH^C24CAK^GVR_Y?GY
^-H4cC_L<8YUU[1W;#1JebJM2V^LP&1QgU8FWB1O;1O8\S@NN[cA<b3C,T+[V@S:
]gYATPNT6XC<:X69&;Z/^Vc@<J45=;1<45=4@ZZ@\ag@XML@BQ@eg,]YbE<VF-?K
>,>\UMa:d2T:+CfU?ffJQT1BV26(7[1c^,2@4\TDUVMcVOJMc@Ba@A;PbK&,g.24
<OA:^Y:C4#0B>3SZ8P=52R15LaV,#VM2T0JY6H@4<TZ&_^VBV1d(LIRBO=<?3R13
1&A-R8>d3]BSZWA,]R++YFH5-JWcX66K\G+;MMV2ZF_^1I9WA-^fF[:P_..D7I\d
gLIH-&F-6C-W^M3e4I^RUY9N/4(0]77)[MY#P6:A1aUG1GgU)-aM]fP-@?C]BZD>
L>0TD\;K/3?_K7UYc.MSW#\T9PHG9;SL/I=,B8QM0GB./5aV(dE\VLH=V&DIH/0\
_TF)Ma#KO:>@.LU5EV[.&1K.Y4\L7_]A1-6:5L\e1U]DcU>KC=d-CU[RU8^G@bVU
O2^Z?72]?6>bd,Y#0AL#G#[>F&a1Z#[.R:bBQJ;_D([;69dc_b-TSdBYb>&<NaB(
0#0<a980eeFM_Ta9,IQb7;21.R^4M7PD]FdDKcN8=Q=LKMW3J1gBd;<Yd8XXVBYC
X\4\gMEYF<aP16C;FHJe85_1?C8X:C_1<A&ZHD)=BX^O28RK=K8/0..Mc#1MgHA^
EO;PP+FV0=2TZ[9GA4)bWH,NcR:feUP7[Kd\JTU[RR:NE;PV(EZaKVY3g[WUAD4E
2:307V:=+]/e@GJ:c/.7ZUMJC&RK@ME5@B>b:V(eTBb9b1UM5^GWBELbXPd-@GUP
A@0/[.S6<M\GWY<)aba1ceAAX.;YN&(4I3XWY4TO8/G2MH#ZaJe__S9Oa(Q45>_:
&)/(;[Y]eX8,T_Z3-.^53H4Y8abc4BDSI+:0W51D)5.gd86EZ@5Yb[=#S4M58L;;
]]EQAQd251,^0GD[2?L7b=SX+&JK28R_+GV,<<f@4Y;8HRF[TN8Qd[BF:\61Uag/
bU-RL@+eGUC[49D?KBMZ:7;;.;/SR2EUQ)IE]IT[,X-bTURJ-I#UA^BdeCgTc=4J
VDAY4;\0G8bV/==Wea]SB?M/7dON,MOD\cR)=@[]?gJG/J:&Z-J/Z;\Ngc#=QPG6
0=H::-FR=Q6;.RD-C9aMeS&g>EOW>((4aN>Cd=C@BZ\85F>Hd#Q5>:^a4ZP_(J+F
aQF#6N=6eD5N8C]\5[Y=W+VZMY8C7MJO9IRLGM?[(21cNHX-Ng?[da/;G\-P&g&K
Yf0b3a0_E)F+U?aHB^R/E\VD,WO6Ee.[Ld[IK^/FdZb\G.;WC6FaL+VJV+Xb_\8_
V.LLf5Y8P(TNZQP(;eI[MYMX[M+>ZJS6W=JQF7VGRX]&4CO_F?dY2^._Nf(:-&S.
YD76#P/cULT=YS5ZQfXA\bF]2e8UP7D81/PJ9AK(XT[=9f&X_NMYS7fS5+#a)IC;
NI4.gWUX2(N.N3P;_f93.2/Z4D//T,Q]gUU)MbIK1>X.aDU#T]^<^-,:GASGB2R)
TC)V3@Zba#L9[f?T,B/@WbV#+?]gYA5bA<,Z5AdGK;3K1@aNCa7&Mec6Iaf,eC;/
CN=RQ]QI+gg2-DSBL_?T;,DN.WZBP75^d(J2Le.&:M1F&<Kc7^D;\SM^g2]g#78F
75Gf^P/_2NA_:BD_\H==27Q/OcN/Vg]X?5Y(=)b8BZ2.19^0QV1bJ3+P58O7-F<3
Idg2+S3,UT,dHU4KEF:ELfc9[4ZF47XN5\.-DFaN3J:O1fN54?EUK\S@8/G8cg3-
RXO2YDBY,PPR,WZ<d/+0?8f=P6[+W/N63IR3OC#=.&E8C^:Ia#(L?OFYJ+d1?Y0-
USJUcZ+9=BJ<S(2HDO;.B(JGRfGIU&=E9&cF7M&L\>=WG@KG&#Bb0CZW1.7RP)/d
T0XP2fG10dTbEgX5;EV2L)KG0/X\1-Pc+Wa<1QA2eJ^V1QF=dX<L>eK8Y\?^/56C
G;)ZXLHE[H_)D#S6Q,;]&&J/1/V[O>1BCB>-NDX^T[W3IAQ3L2A8,?3e+6MGAQK7
UB/3a19\T6AN7LA0Q]gD&QAIYE0D:2cZTOP\RDNb3UID1._7bDeH/cC.AKR#RP/X
C&8Dff;D6K9FZZ5d,.Ig4aBF(>NV(+XWY+9gB6BWGfg5?QZS052.g@RT9&a@V6D3
DCGLe,@dK0>343&W[PdSC>LgZJ,&.aXB[1QN@W&-U4_E7.&T_NNVZA[+dXNXSY73
T+W4ZH3RaMIB:UB<2I3A1]1B8W1Y0/4E2dFU,3##cfdc2P\8#c#,?K2=b^a.&O@R
]+,eH(LC),O#RTI2f3_RQXS-M?@<3@AYOIB;+]VG1N6AOD\2>MCSQEFG-La71C3<
&CE)1EeL>O86Y2000AW^db<gVg1f#HbOPF-?\R+,[2DZ[LP5ARc-XU3W@bR&A7^Q
aX?4dTLIQOEQRUFCe@7<#cBV8_4S]8/d9b&?@fA#bFQF2J/[=EQPAIPNO61QXTgE
CXX3d[))^,5>.BNAEX.MT3J9X_eL[3O-[d?N+d9bfIKG-=D=\Q]4R51;D3\eY7I7
TAW=dK3>QMSM[PUPN4#7_4&D8b4?4Kf(W?]M3QC>12g3(BP<JTV1Y7:L-)?4JDW&
EI[@>?If-VX)c_cNf\C,Vc9(;4XDE,G7M))F<5@6cd-TZ2^?Ic<6Db]SCWUDXYMg
AZCKUT?P>XY]a\1S^9O)7R?D<6ZXRE@7)_3X34O\<+&JKG)N=5RYfUcALTS,R.OA
a<;GMB4W\Z_-Y9U]&E7>-28#42FEag11S6X7e#gM7).B&RY0H0E9a[F@U>0R.785
C.b/R&JbK.d+SE&fe\[?bBUC6KegdP6XB-F._dO7_/g7JXI25&N?F]0F84>8VT&c
VN)f\FF+94PI;(=5DMJ<:L9#38b,FD.?P_6ZS)e@KL-U9R=ae0Ff7]5R_M[>:>G2
_.ObT<@Rd=^F>9=Y&a<O=9+Fa.;97FDK=17DSV__aTfX&A>8],fJ,DV;f]YJV)^:
-598.+Y(&V\Z\90@6F&+YV<FD0KaJ_P,#;<;HY_,57WDa33<1N(6e[A,9b^d5Z0H
8_fH=.KG[>W_;9\dI)O;8G]CYe(AdN+<6;RMW/T-_ZR?M=)^cb:)dKbH()P^P_,S
B@7.L/X?g)3^N(?:HN6X_UYF<6K;AA14=bg<,FHF4<QL#R),M^b;79R?LPK)+SGc
Y3\NBF4/.(+g3(WLIY,HQ+@@IRGCc5\^1-JF)[XPPLJ3ND2g\X\B6f&;+J;ZN&9G
.UW>\RC3A0gBdQUH()BXCE]4UEbbU).VBL;bD6U#0C\4cIW^c#.XP_a>FBK5^B:]
-\@M+>6e3-b=KGS7BPJ_@@77KC/QN(+B]=R&9R;CZ>GGS(S@57cM9?Z4G0[3=2MB
U6EY2PIcD8FG^d3ZF69\F_:5&ISU7JCdE)]..-SdW>;@?4>HAbZ40V2S+(d]^1^3
U?.9HIT//E3G5Q_C3dEcF#S,[e(J+SP^8c#0WZP)7O5fAYOOC0&P_F62?AYe+NW5
@^[fASI4?A.f85Ea&Q,SQ/:KT_P[DZe;2:dd3R>MY&IZ^^T)fVWDJ(Oee&g@P5Jf
Qe:XYeeYJeH(]]J)Z[<>?Aa#Q5H_H.?c<,DPJ5,C@a#GX/B0H=#>->(A.2A_4/J;
(D2)<)UUZ:GMC(=4#9+CdKFVK;?9XOQ:HG#G/:V<W96ZU[M>SdaYK]B8;]ZCY=P#
A>4I+aLQY0F#CG(_ffM.ZQ-GP41\@7URU3,:Db>WAJ:EHAP66W7geZMR:VME+5MA
]S/8#fSK]J3?Yf^gE?a,g)CZ[Q)&dT<X(O.Q8G+,\2ZH]-JG43(Y1McD-G/]Gd>b
B5CF?@G.R#e@4/eE;N@?A..dbg7^3T3^&JeI:S,2aQ9_F+7-QX/;C(B_0,)0(R;-
?D:[X<LG=\#eC=..?-U,B:Y0c]f)9VE&.e?.@:^1TURC6&2:\47W;_)),E]UA5b_
Yd+9YOW+VW<,NcY\S<=R5UaHfcAFXfIW]+7++.5U0b34<\V[g&#S@1AQS+?9A]c&
<F;:5Z6^b[f\Xe4SP:CDcGc+9\+8&(\3F(BAL5Y?+5GUgB9V-<>0_4OGH@KDaU:a
>[D:OA:]\()G\?P?SOS^+4E7)-)D4XW4HN2U@B#Z-4=<;_O9I^H@H39_&aa6-+H6
ZSX&(U)O-IAV:QA)b10);R(3?O3QE?9EC6>HEaS(,Z(JP5F6;5;Xg(3E9A0BOO=&
Z>0A=A#H-E]ad5828VTKK/dWU64;;E]]]O]N4B=8LTD^93=9OTA92fMHc[d0\\L_
8DF,D[XJHH/1L/6fOb3-Z3X_Y(:<@@eg+R+8?BR6@e@Q(>ND>aHF]B0#GF_UL.;O
LVR@c1Z^I,BEG&S2a14M,NN5KC=J8);XIBQFdSZ1[?+gZDYJFCcBREg/QeUb1_[P
6GTcVa@ScPfT0gJ\a74\+H:c/?dI@6fC^5HEeA<X.C4#T:V9M\T>dY.Tfg+L)^H0
>d<+=:fJEQ8/S[LX5@YO3=J^];SD0.4M:I#4#0IE>0F?IR>)[P6@)7QT&IF-11#&
L2TXXeFD8S=)IRBBQT>SdaKJN)JC#+\N=SE<^T64fe0DADP<=GI1Gag1-;J]cFYH
N86<]&c+0S=XgcG^bd>C@I3]^e_DX(]f8P]@\Z^MB?86)A>DC,\)F.\501KL(&gO
[^9Kb@Bd][>a:fBA-N>(\J(OZ=(RbO3NLcdSH01RdJ4GT_R=C^X=g#gQ[E/9OXfH
26D^.,\<>@UcT>Ad)K&WSA6N01(Sf2)Q2YT51-DL(4-DE)8T1b#U0d75J#/Z[OIX
8N=7PO4a7cK1TZC-Df()JAA#8_ZegXROJ9_L6X._fBDRZ_^&[A/&_Ga]F82T3dL8
:AX\EB51=&8^L>;+]^DON3LNQ63a6+9IM9ZR[Y?X357bC,N5R?F,VQIF9=#_2d5Y
5aZFG7XTV5)2/CKFX6c(D[>Ba7WNDB#>c4/=Tab?f,T<^MbHPY8KgE7UXQgO@78<
_/9cEe)&SCEWOI39E8[I6;I9JcfE1dI417e7R/OHfRGQ@DFeDV?.,J_Q8;&_?aNL
Fb(9=E7]^==2<PC51FL5@WH7V.:3.fD6U0S6F#Z&]UB8dV72d[F?T-H?=f+Ye#T>
B^DYWQ3DKG+dQTGGZRPYC(-UOZZ@]4=P#bOZ(Peg#GV(6TP>1@4g>Te0R/,(:]8)
RA[P2_UD0HO5TU+DC>@,H07J>GKa0e2gf^9#>f6/Z,+cW.^UYN9P46P7Z\aALXEH
;BI;&F2QZbXIR\772HJB5R.F&3S&/;6WO#=X+&Q^O[3.Z&Z_C00>33[3b]#XA/G[
PBG5K/0#S9=;P;4CP<;(R7g#W^D)&\b:G,?E0UAN\d4YM.dW5,L9=BD+UUcO/ac5
O+X1M&X22/]ZQDW_cP(.Z.GEXKS_J]f(II/R-V3LE2\@F.KD/]/#(/3^;&O5EfdB
6Z&W^:9GJR\DF2+#5ff^916cHT(Qc\aceLWHdbfG9_5WbgJCcaHHV&&EI;,3gE@&
aEWC[U^D<=HfQY#EaR@GY/G_:)\5Z]#AL9V8I;V+AQ^V(]f/M64-(>(Q.I)-6d12
Je;8W(=P0C>]WTNNIMRd&HYT_6#K=?2<UGcfU(.,fR3GANP.^X=D+&9(YA+Qf6/_
&5aT+6J5:71[_RZ[H83/c[3LRURN;MEaHHQ&(N:OLGGc-7:f=>#7(ER]R#C=g<Te
1N&^T&6^X\SKHa@V9+4),2^LQ#C6NFfQ8?b(gOAVYfWa#VJ0CQ^CN4.Vf1aK/#e0
.Q;3;3_>G)(_fK8]P;@&?K7BRNS@?FKQ#\K3MBU,VD78S^eP2O&1gZ-V8:aCgGd)
+]O:>M3W;27^Q3C:=#RZgQg1:6\<_KF<ACX\]&]\>W,H?T2T5cW=X)cAEb2_=;WL
0.N3R8OCdM/Wa2>M\P/,K99N(KJNUR@d\[)POK-<]B<\T:R>\1H+3&fdCL@K2=0U
/GD/V^LB)WAGPg8YWI/1YLF=.71+BI-5+[?ZGE<_>HI:;b>PYY0N_YFb/Z=GcMU]
O9_C82Ye/QBD;+.GI2+NTR-E0dRUO7a:;@A,?>VJY]-g-1cc^R=bH/UP.g[#W0f_
K,W=D(A7+Y)ACf16U/.V>X-&GYJ2ER#/Ee?W_[]XC()I6.F=/Q_ZJ>C)&;UM/-2+
e>2T98=/63EA_?QSU&U^[ZRf=I;0d)V2UKK#/-SYgH[^)2e83Q\5L#(\.[=<AVPH
QG)2&&9PRF8+HP@L,2Q0cTS78CC4/[LBD>/fL#e\;1N3AI-7?@Ma8^08Z.4U<c>^
K8&YgA2g@Y&FBQCR_)Gaf+@fgH),M;e]\2Z9JMDCK&=6Tf.;]b;WUA1-01Oe\CQQ
@+X@8fIUF578#gZ4gZ5.H^cRJ>Z:PNc\9H).^6<Z407GE>^2Y9gVQcC/3(8R,P6;
I=JaI[e/bA+a3fRc+-_;?Y1FN6JU[fQ0NI3X+]V5=F+(70NF:7LWK#8I+CP^85I5
_^Z7M^Fa.ZEU<,?Ab9aADNQ1=DeBWQD=&I5a;GU,[@WYAdc3dWJ,fda0R-XS_+PS
]a@R)O#KV+g_-<DYNK281_>\Q;aSK4QF83);.MRQ.<^]QH8aURa2>SF97Y;.3W:^
2^.Id288&ZIJF#\eIQ/PDKdcM_9cN9G^GBJ4-7SQ&cS<YKfeSS#3[7Y&\SWWKI,,
W53O^\bDg>1?LTc.FX>eHJD)b\I(-17HWO5fg<(IK:)F3AW8N@P?Yd8f\c-O\)L3
R?(RI?7PUMIE/@S+A_P?JbM&&ULd)0D.?@0ge6+&NXf:AWC1=6UULG;AHT0DA;9d
&:;;LJ8ES[W0W+K3^&<4[2/0:;4>XLF,=WRG2L=^1#RTKLP=O8\aH&+0M(<7@;UL
P7XR,GaZ6-.X10+3:305H:U&1HY()cOCR1<gZ&,d_1_7g4TTa(RYA>9C79PR<YPS
P,4-:V;6./I(N,Z]>9eNOO#MDQe0<[SBRW)14SXgY=?]I&OS40J7AFGb4b<UQ7fU
PeGWSb/K<_PT,7?FPYOH@YfeKc)0UX=-beW<M\>XMP3JMYD4b.S-,d(MWV?E7>E\
FJ?H[PSHXU9dWg_cL)(OYO_>IYEW?HX@BW0=aF^D=OX@Z@JI)JYU]U<c5L,8XPWX
ggV+\>^8TC,+MMNL-/Lg(-R/:[Hfc=,N/#A/X9()D2cf&W(__LNI9;F)e@9?ZU\6
/]gLg44NOegGD22dJ(ILcK(X1GC4Z:KUX?W@F)QEd^??bBVSTC@+M2\fTg1.YeP-
f1Tg7_T1b\c03OACf\3O7HYeYK4W&N\E6=OD@H1)WR<^/D^:Fe+(MWYB0@X_JP(;
e#9^<ceL4X;F^S.XU@7]@G5;B7(Pb^]9e<Q?QH]THdb;;84E=b3)f42)\TS1K0M)
bCPd8L,?FU.de=c@T1gB/7#AX^\_76\a^P.#fOVC0ec(]^BMP1S)HD?ZRf(JPSWP
5>/60\B>J<HK.HgUV@fGc;E-2gT=,JEIYP]VcE@V]E_K1:](7Ma5Vd^.GdU42:#<
(@/W]]UBPdgDCL)7):4MRQSG.O=+fKgc-+[N&>Zf?e[XaAR<DMFN4QO556U:K<2G
2.7a30OX/KR5\[>-PG+F6Y?LA[-=g1;/4F_DX_;;NaANG]5,QaY4JUW.ebN(A;Z&
Z:M[AQH&GB_NW0OSI]2LfgA9VeJGU[^GD(-3J1I09;d[U[13dNZ?O>Wf.#2g;\[W
<5fEL)_\K?JN<8(2.B#7\a/G\O9bNPZUg;TL+OZ;+T>JM1aTc@RX6/dOfC],SXW&
DFM\<,VeR3+/EVIK2Waa7g9dLLYN22+c]Q:<[POdecddMQ>g:f;g_(1b5cJ6DdN8
2?TFA+K[\JO2@ed>:MYBX;dgePaC=VgMO^f6L;+:&,.3\_Y,4<cW55]98O#96[=U
)__VNZU:WXSO(WZZ>&-3BcWUT4TS5G5SMWA\W-0DE3[K]e+;@X@CG:;E-U4G+L(U
bZ>>K29.(,O/8.B>8E@^.:SIEcBEULO#@;Y6/QIebAJeVGTZ:#Ld#e/2H2YJfB0;
59[FcK]P7SgC#[:=LOW;\D\G9><aCSW]XDGSDe+C8MR>93HWeUW/4^7ac2/Z)]-g
A2&EgX>7VHK^73S03Z8[TBUYOP0de.X2<.7M.5._6\O[fYa]T[8P+36_7VT2Rd?O
C6::2LHe?;[8O,B9Z1:dWJ5XPL48Ee0\Rf9Z5R&OS^J8W(D8b4OOIV5N3;33/NeE
=0/0@g500RFfKJUBYCK0AfUE[_,e36^EZ#6Ya(G\.T^UCc]M[c.Rg=Zg+-Fg-#4A
cD9=P&bA^c/74-@ZLd/^QecY>==@RLfbL9Rbc0aMPHBGZ5eSGU8__\G3fV3);+PS
b@JG@\1AOIARM272A@IX0Aa.;K0K.E1>RD05S?A2Ba(5&4<PZ3fS+^c##0<B3.43
-]-TO,:VB.231XTLMVN/1XMMR7daJ:YF_2b[1@=OZ^Gg79;)B2^COdNc,@A#e@&H
Y]-;Fa\F&d7^LE=K75ZeWAGB\XF)R]Z[b4J#>WHN&QND2?c7g<_=DO@QACX8DV4]
_K@ZbP]^;K,C+KWTC7aW8G[S5XF@5=/=25L6)C#/,GLM8]]P^cPH=Q]+/[Ag;3:d
D:5dfCf0R1>#,[P\\&DLN=\Y[1AS-6Z+VRPL>^BDe1>L&\cP<O:R0d4FR2/1/9a,
3Kd,g4ST.)^?g[085U\[#=CO@6/OS_T2a,9I2IfB./Y(X]<OHQ4[[WM9]+H^FZUQ
4.FSUY0>UU;OQ_Y_B<X-,(-N=2:NcB@RKEe_4B7[JX#R]V.R>f68D)8A>CMCL>XO
\WEUSfH#_La\75[Gd6,J)\@57._NGdg3:CTdF_0<fB0L8)bKe9d3-+aP)O<?K48K
U&=@TbUOSKbSF@g4X#:EYEFeZY]dN<V)^CAZ:=&DSXF>>5FPgVS4^KLNU[__DX>?
^Ee1YU:;(bT1Q3;GdJ+]S,6c#Kb,B8dN_FU1aDeeV1W8QTS7e\49cFCWH9UE#R2S
AKT;#HOX<?2C4U+Lf;Ze-_,g+#&<AML]a)>)d1QWYA#XR+6SV5WeAT)?&-&3GdN[
IFU1KN[A/SETL#15=@KF2ZZP-C.(GGa:(E4GQY=7JIQg[a>BP3>\M[If4Hf&9@La
;C8d4aLM)OBgW:Q,Ig9)2-7g;MQM6d3dB,0=#C^YIFa7@8eD\f,X/RG[28F,OF._
eWH3]O4Q/S3IKGR8cJ,]2Q=TXGeXB4EI0]9/=#Ab>^UgXG9,BXYLdXKH89M,E_I,
/M:-5d8aLZEQ@d9479X+<MA8d]9VPL3L6=69+:LcKe<[PQUaO-)/)_gWB^cf6aFE
g3Y6\=I1P]5Y9/:^RJ>?/>S_6DWX(\.@:JHCL4g^g#cgaGT]4;>#>/93,3NbY]+g
OMDW7a.M0?,=J<W-]1Db]D\<1J7Be[+TZLgbD=>Q;X9,R_egT^<L?.35)OX-N;GG
E8FUGccDbV)ePXM=cSa3a0ZG=>e899_@@W=-DVdH.6=MR_6LDUd.114Z5aI3S6E/
D#5@dOD.N+OLGD&AV4cMPc]aIBEV6)UC^WX-_72:&bM/;V+1Wb_IB7#aba##8SL8
K#3ae.)L]VCDF.4&/2T=O_gM2@ZCQNUCA;O^XQCEFHXa8P+>-72(YBZ>6>Wa70c0
V]ed(f+:AY\6DgE[3PN;-Ve74LgK^XY+a114]_YG@+Mc]dEDCU(KcC/GeRaB\d)G
X6DA@UeC0;:C_Vb?YFS<P877-F0<X06)O-\N=a<;a&fL=T@P9\dI;>\JX=E3[\/f
geP-g>FaLX;DX8d?^,Xb1.1M)5D?J)HP1#@]Fde[[Q)N37dgecCUT8J+eNQGLf<P
dMUcXg346dcWT\<bZ9gEY;1>375)1@JQGScD&4=,CV@]dYJZIaSSA?R:9RD1HROV
a2]Y6ZM,4[<2_Y3O2_JAg45)R3)FML=>_O&G3ZV&E3LHC5-AI/bQ?1R[-WGDf,TO
./4B</K.;<6<)=Z(eg\:UgWIVMe=Cd]U4B;_[@^Z(8V\212,Y&@(R,1>CL)JZJ_2
:^#\HMT]b.__B&fO4INBZ]?Z+371S1F>XW+<5X&HgNR=X8-KQ@A?.=)U8DA(,O/V
2Kg2QLVHW3X>DP<D:+Cd2>_41Qc+WJb;f(X#TRg/V[J?>S6,-UL1Y2CUH+FX([HW
JX\5gML0E^I9\\JV87C24dJ5c8G@_]FB2)V]f;50XMICYDNfA?R8,Dd>agK-9]65
O)VX<cU/2S]e9YUKHF)a=d&P<fAZ^2Ga73PLA\#<92[FbI?<CeS/CXD]be4W\e_c
Z-:Q#GDgQ\=COU.<W=Y3fG^\2;Y)5\.^IG<(FfG:B1RLPJ@T8g2:Z^S2HVBP0PK1
9FEUS29W3/U&#C+Y^d68Ub-P0=-b6OF9<M0P>E4X--8L=6[A=2=ON+#JAI[d:[E8
.c<JX>JN1^X)0:<7:dI3;:EVQeAAAM34_L&NfB\0<4R_]KRZdcX6WS(BA/M@/<8\
/?;@a[9&14Ab&-FKLH^I5f./TZU(I],]bMY93EV+U&?:@.I2_/4Ibc2Rg-AWB:U@
;D1f,HZ-@Y:dR2A:)1E.[d9+7:c\59<1859cXZ;BUM0b77,8LHUf_P1EK):G61)O
QM?L)/04NKBXS(YC92:YZfD?&>/E;K#(DeK20W5Y)#3eUf@X>?VR2:NGLg42:U4F
LB]gZCS<D\LdJe>YA5GG2[M)\7^cfI^OB#K3OP1CZ+Y[ZYBJdO6?UOgSS07C-?MC
(aRKO+6JXB.IWIE@>)L258#BAB)ASDPZVFNOG25WBF(WN;M]Ybb3O\FJ9U#eO9&L
_774THQ35N+AW-YS2d<_5T=O)IX(]SI4N<O3aB_(I7N.ZK+.7F+O[6-=cFZe+UV[
e9:2<+0<Z.>F?#PSN_LILFT4P3Hd?S\SC2@7HH?d=\a@Fe]DNY=CF3HN@GfcQ4KV
4AFKeUg;BE^#/C1=/8#):OJ/d<5S&9HM]?QSSA>cWWa1;e3fQ>A#e4([HggeLL7^
(89=Xg&Mb\J8D[\dQZI?;P&^^7]]_I[9]<=KHUaRWGa156TPYS;)MF:62AF/Uc4R
G&,Og<:#DKGFYF&MZ7PK0+SLd]e;_#K19GJ^2@7R0A0+&16eGeB5NT,2:,8OZKSK
Ge>ad>OCXVF-<VUJJ7H\^eg+L;S\a\_/eH19BNC:a9[C[S+NR7V5A&8aVOYOCY-&
/eLfIJ2)9ebSa+GKDSd\98EYANg):^F3ZR/,TO<5S8P.<G_W:<&D9JdJ2(X);,25
A:F)40bGADAICQ>V\GX[OMf37@a4aAJ.A0FU#eL]OdGMNRN;OG?9G1HSBNacDebJ
,QI-\_6&KBU[[3P+;WeP]2QX;.2V)85.@]X/aZ&+T59RU,&<^LAW=#B;R;XH(UGZ
Dd]<5:1ZFbYR1\4=B?DfD7ZXAO6L0eAKf-4P^NFHNPBJ[@R/1ZYf>OSTfNf-BGQP
HIa_)\V7(-FWX]<94-[GV2X/C>[C?#ECVGfCa?NX4J44_1790UfA7RR6,#JI)9Q?
4Ec6fZ;S2GMXP^53G=8SEL)IaF_=M/Z=85I41caVdH60b\6K>0/]P/;VP<^Y?)&&
a[T3_1(;<b,=NXTeU@7W&+ZPgf<DG[Q-=[PL=eF1QQBWN8O\>1_\W4&8Y/EIS_8f
(D]OcVZcQVC6R0>2)0EI5LdB9H59a].6M=+b#DEeF:&I-G9(.0fW:GZ)K6ST[RW/
_,K=.M=7BHOAU;R:C2@\S)VAX)@9f=L]P65J2g^\ZE-=0Y#+[,f/O.eN][T[4JG.
gM,<#H^Kd19=IF^LG#@UR]6e;O-ON-]gVRW4NQZH;c<H]XC42c5N37X:4?GC@[8S
e=g@Da2^M:;N5#G7+R9e954B-<+1a8f^B7Ne@007@5(1F90db/a(Z0]Q6ge/Q;6d
Y>OCC=TAfO;148DVD#I\56305J?T/a7S1geLQ]L)6OQ]N1cd#NN)D4GF+YMgdV2-
X1KQ65\#ZM+@^\JS;PQX[IfE:g0W3N9?ea<6JQ\,NFT^;fCg,#P_)/9[)R8>,ROc
+fI(AA_S9.TIMHVC^(J0EMA7TSf7F_(d-WPG^N_(Qa0C3f4KDTG(+SB@]RLQ9,_B
SKUb&.Ab5+f;c.(7T]TT+92F3JgYSI_YC[\,)><.RD,2<XH?HNWFN^#:=NLB.4?W
&6Q<(.Q:RH;GVYTO,W\:(:BPb(-53L)e9^._BFM4@7a\bW,4O\dH#aLZ,^4<GN9c
=+K1c=5QOe\8,BXf0&NLZ,NZP>PA?0[/U=W3I]B4DH\):b]MC4Q8R>PCBcYKM5;A
)W<H(O[<]).B0F,YR(PBX_U;4L06e(K:O3fNL&:T=fOS+,B^+;+d]aB<K:_IVL+a
KTA8=O:#^&9]cUf1&3)dT=BKM+:<3_]76#Da,RC9BZ:Q__COP-<fYXe/0-70YKWW
4>T#_I82-+UVGffF)L&-Zg.8BG_6Y9)]]B=J1PB81>?V(G><.ZHPaUO)<?OeXON_
/?EBB81&@DeV<#-[L[dPRSe[\25(5c]ZPUbZcW)@5#<AUX0S^gVXZGR90<R7]&R@
aF4)5SO3Hb7d:)eTM7Y=TK9EcP7>Y0WE3Zd><Q33Q)SPbeEKTNLDMMdLcLJ+U<f@
F</a0aeZ-g(#DS?L;;<Kbc^,VWK/+JWQ@24JVYbf?0EEg:Vg<7^NP5++^4\\c_9C
ReDT=_b,]Zd&/)XfdJG)?K?<O-@/5ULU++((([4Q.&V^F2&f+[(b71>WJ3g=R[KQ
4MGaK[B>ed-RNNSM<A?0]77V(DgA]3KB/KV_6B6.UPT1NB:B2fQ&?E-P.S_c\Kg:
D=1HVb_S836U\XDe7Z.+8e0\(8M/YU.bV:FOgPN3R(+#@_KgUc93(:Gba&3,G&0^
7IL[3=)X^1JD<UH;7.4J#P<C1YFY<Zde(=?.J<UA=8DdIaX(_SCVe5Q6N\5fF,DT
32fKY,];0L1)E[K.f:3)-X>Z?LLb]Y2;=G3PW3A&[U5\dSKQLMXQ,FG7@>bSeePd
?eER;YY+[>gVd6<E[K_((\L#EIHfS=_76+^T^F7<RW0JN_/1KJO.H7^BMB62)>I>
)2=eJA?gZLC<6F<,gDDR\,6N>B&(GK4A&)Wb492U2b:dP35UX[HO<bgcf841Y7N[
Uf\-?NO(<;VKf<;Veb?M@[_c)F]BXF3P>CI5B1+d(96S-gHc1>AOYQZ:EBZe<N\2
/<KC=(BeX+;.\?Gd6IC&H;7Zf8D8Cd@L(HM5,3X;[ddC)DH7IXG8\-63bfR3fL+D
J(<D+Vb^.,c5Q54=\>=dS_U/YG3P/.;15#K2]gSbQT8\L5OJLMKK&H1)a0dAfFN(
E40EF0]L_UR7P3-4MYKD,AfXO3T.PU#U0EWGV+#<W:M?c9EMJ9)D&eYRP-Y1F?dL
b#gR<DVCJbH?L(FX3daG:HS_?X/-1)HU49_QQSIb?7b2FOdA.A8UTU)_:4MXfLI3
?BMYUH+F1NS1^gOda&a<>.S];POF[T\DCGMH;@Ug#IHR6G>MF=A5R+4IA^8da;S^
2=\EEK?Yb)MW8XbU0dH3.XL7Gdge@g85XQa8;-,^0f,AELLaW1X@R-@_1?g5?]ac
W]X\T^1ef=[CUH)UPM>TZOO8G+f>WfWV/@RAf7SL8A_A7CTI>2PDdR;N[4R.AN7Q
+J_cMP&OHf:gH\&S6-H1F_:B6NWAW_<aHZQI60Ob07<)EVZJJ<)L[3<8\aJ+V>GU
bR<4H#fa.gV0[5McX75<DH@(WaQ:.Z2;UaXQMeJ<-(9=RLU6@CQ?EOF[#W_0KWMJ
WEB25UPF#>.)^GH9&PTSFQ]_GPX<D?19CK>agHYcTN?&?>bcJ/OQ.bSWB?R[Z4_B
Y_GZ?c;UO\V1b<(A\H5(Z:&VZ@R.\8:,1Hcb]a7(RJH)/Q)B)7(>LR_?>4B1Kc)d
+N_?(f:?ES/BS5+<[aNN;2bTd6BK9Wa)>U&LR.(gLX6<I>#>A^MdU0g0<);P7=+S
M<D-,HXb:M@D:5Yc)V>gEc>f9H/1KO3E]_aHB+(CF1g6Wd[S\,_L0F^\?:<cMQfN
3KS4:_98[Ac/P,dR<WdGL[^FO/\dX&]=O5H76eedU]H4Wd5<ReD[dYIK;^#;-)fL
9)N3fJ@EUE4<b62[>YdWN7HLWV[/RO_9eEcQAdL;6WEKWY[<AN:LP]XX&#P^E:cV
#Y_JZ,CXABg\/:&)UF_1YN].@R-EJ7e#<812,:+=AWd/4HHJT^<ZS:HM=(-(S>F8
g67_H\f^b/.ZeG3U[Bb]OWXAO),]SXaDFHgYdA&\/24ZRc_[+M_()QaW>EUMHKB6
E_e]3fSc.00V>Q=/^5695/&3+.1N8MGV+63JW<d-c4?9e-=9UMb_DA=&Kb,:4N/O
FJcM=:#L<U43^X5=F:C(U1ZWL4>PQL-P=DJd(B))YZ@/PX_0D<,+F>G>/-;K0T[.
V2+7/S>ZdEC;_D[bQ9f63A)=EY(G,;.dLc/-fH(;Tc();F9[)QOQ8GH4egUZ^VZB
&>(SP2XIYSSBK0VN8D(eE7N,K5HUBW:B[TS&G)KX\2AL,[-aXTP[>gU:ab5KU7GJ
&2A9M42&PSXB_U[=]>bFg0M.#5?V.Y(A^5USPK+Aa)[E>1/7.<]ABVT8MbcJJ=W#
V](^?83R@M)BJ-8M06g1I:C[DG:D17[VX=T)b6#1,E\f&F#I+;P-I))+3:e[/9@E
L[ef7B25;PP9(T8d/>06HPX)46+EB^\0LJLQ+M<GC9a@Q8?V7.I_N[=,]:dRQ:??
77LA>gL:4#88[2V@a.52=,)71DSH7YR4Y&8-63RcBfHdIe,OYb5U+I-5[I)PV)\8
6XW9>W/S91@-SM4UW499_\OcUFZ3^J\XK>(c+;Od1DBRJ),@VF6QWZ;5V0:G./AS
J5a42AXaDAbLIVKQ/d?=]6+VAd-O>GW(#.V+K.7_Z-3AHTeU3)5.V)VGJ\A+^&XT
bK+WZ1Y1#M3XC&AVeaR7?/d^<QJ(MG+G@a5I:cDc5A3WEc?bg]RT@d2Gc?CTe9I&
9PZ/\BO_(d@@c8,.K?I..d6JXS8K]Hc-39BJ\?+<F09<\RN;CPRgOg4_S^/g&Z,X
TR<8BQM>g=#K=<E:N][P3[CX]X+_8Zf]Q4:2BOWN]L^87:bVY)-#>0f8[1BDDc3\
(,=28&a@C#E00Q9G;-g:D+Ve??0Mc,I>BGF82E3cH/WDXbU5db.L=U;^F-Ye<;gU
:UVa/WC3+;(Ic_EQA6c#CG[3O+&e2?[<:<B4,_4-Z[^\\-=WIGf:6,U,cI#-9?bb
&IXIdDN6@G6ZI9T(CKL)_&Z.944\7\U+E/3T;4Bf4::CY0([A;7D8MWL<a(fe26c
b[#Da<0;V/C\=WFcAY8Z3dFBXceLQdC.=<U-0MC;:b:A96/6#].05Ce>1>X25^46
0,B\[.YSI6&BB76(L8\M5SH?O+caF^[McXRE=M##>>@OE6GIB4&D<O=c:H-b\fHD
KN8[cF&gb]DI0HLDNOQK/ZZ#bA958ePYMBO(CZRJS?V=E4G+A_d1fLM4e@7b(JgD
V:a6a.B>X\dR))1Z#,9<(/E=/C7&c9RU?RVf9J.)4R6T@6V;IYZF48LITARMeXG7
EAALCD]D.M.0,VMe[O7=eBgPUYQ3SJCZ-BBPECCF7#eO[NfG&TNK[YX;@H8OIg<]
:A1JeLQD;g]_e#FY)[6=#6UOe&5c.9KAf-c#KZ5/ZgS<I4Q59.G\6]E>]8LK3>.U
?ga9SMf.=M3d_Uc-/.692_^68HQ0<SGIG,6_6V#AB>/&2&GFJEDA)XI1O3J<6RS.
Z@bEb<aQB^[C@MdB=E;^<5BH&_.SX?a/IC[WT\\=_WW;5cD,<4ISLNc-@9>E)ERP
ANc=#QVQSQNd]b:-gQ7U.8#@XBY_IEG+JL-@O[+B,6#Z(H7cQ@\W3M<PH3C4?PXf
-)C&bc#4.W-9I#=C-2#aMHJKa9<Y6S1]EI>H:+8VEH,TWWV#VgO?O7K\,_/T.<I;
2.4PI^<(=-+>/)W^MR6;,Tc),7fR_e[c-02<OFX@GCC;1JTA(1a0]]:EIfI?3:),
9.X3+<(aD-gE9?7bb:(PQ3R.SFU8;5#H+IUMX5>;GKH.;WV_7#S?J-I-/OA;ITcL
S16/gB7^L9H,5UTE#Q[LB&\(:?H4FELO[&J>N/>^4I,INXA183K,F>OW1\\<P\1Z
VPeZ\RW?&9]YaD:>ZMDPZLFI(.(UQ3Y)P--68N2E\/7_Ud8O\]9;8^2XOc7G3E24
,0NVXM?QG-.+>R6IS;)E&OIG]8/Kg(5]5;E<>fAa6cW&fE+8QIGb47JeLEdG70]#
(RZS,G[Gb6TQ@^c3>a0edCBGW^BCFT\YRScK=.fP,dU\]ECJ^2VDYCBNR6LHV1?:
F#M-c>XUf1.Jg)MMI?OV;eQ\/E1E3SFLUUNEWOD1\B<bf\U]:(</TH1_\.a>&7eY
F(CEW.bUJE-2>>\S.7G(DRQ]KL1AD)1d.<8CLT53XAXE:/:I=T8=RJ<=?8Cb;+D8
JTa9#cT>J:B1Fed;/:ZOO=\2EQBK;;36&7W..#DVM,KG.&1?C7969DJRdMYYd+:&
2[RLH,3QKaZKSQT&[C</I.eVc3\ZaALaD7],K_^W)<Ha]DFXO<S;b=JHFc1\>T9\
6FVB7V^(WB3GB]Z0@X>N@7C_L_<g91GP2,c\=FJY2b=/L:N;\,A.MR9=aA,;NJ]7
&OWK9==7VT6g\[@B]P+T9##]b1CC+WTNPT^,MEc;M3)b1+0fIFM3B(HT@>4UTRdC
I^N_?,&4I[,E;PV7L3P\eQ=9dJ?PgT@cea[0?5bfB1>PYRe^H,==W@Z[^G]VH0F1
S;W<.D0Je:g<FgN+=ge2<SX#O]-;@^<W?^>K6:?bS/O1&2^72\,Me.QJFBJU#UcK
Jb_IASgMaSA;=3M[71]&^T>R@aRR>>;S(#(K488G:cR,@2@;JeA,YgOGTT>,8&Q;
/BL:gFJ=Y=W45NM<G?bP]:[df/MD@/WYN5KCPM?15@P^5+F=.d?@-g)NX<f7M?>&
@MKHOV^N[RW_I,Ngg5Mcf9<-2TTY#15d@YfYIB>181IZ(#Y13#-)KHMXVAc\5P1:
[Z)/aL^AeeEGP?TBDFbX8+#WIZY<OcfGgZ^d.N6)gb3:((a5\0YfWRTb1EOW?6/g
)CH,3W\W3Df2L_?8UD[G3U,.M?9TK:#R^O3>7_V[T9]f8^(#.1,;]L1\:ICVa/,f
M+_X\8DDN9eC>Z,GOa,S179GVY2OEH9@MGI]a:M?[8W;/B95S^]HJ80_0ZVK(eH6
.OPXeMGH:U+@[(eZVc2?97F[^eU58UI[Tc3/Y8I96DRF&6OFVf7LNJI_dITWg+-,
B&P&TG((M=61.NWN-F;4[6L]C]07AEgS1(gXHY5=[HXRU(AL1L:-,#Ia[)eBF-A\
ZW)2_YSe)2/(&A0&)7U-XQg4PB#/F5g^B(VR;aJX9ccd?T6(&[C>R<Jc[fB7.O\U
HV391ZN0P5J_G#/ZRGf5@\R7LaHeG8?#(6/?U7+C_Y0LI&EdK,/XTCF7K]e\D=X6
8YNCcXT&7])Qg;\=QO0>VJASB3\f[3BEK-E5/4fG/-SB+@bf:^\U@U09>f5UdXg5
dQfLXb-<,aX;Q(aJ1d0MZ2=/QC88\-6@Wbf/7<1K&O85IdP&IT\6=]ZIe>@BNQd)
/E8I(CbE<UYHRFa:[:M@]K(7(]VAa=_4WK\FIXWOKN?ORD9?2A3D12).FD_;LIM[
>(3?RQQ,[?.H3ac)U/:3DgS/;^9\f3Q?5fDS>T#U-)100OXH4Td2U(c_Q5K7KNU)
#ZECH61IXgOVV6N.V6?d4@e95DdPH\D8H0AHB<N/>;g=I<N&YX3BIPAIZ>\&/;4,
3Rba\:Y9:9a+P,+N1[.=c1Pd+74eRUb.UL0J,9\#X]DCdTd72bM/c3PM5d-3^+8+
>/ZBV6gc/fCf\P[<,(70/Ze,=DNc(Rc[6;#X#ZN40#=B=SI#C2Z216X[R;1:5+\M
=63K^@dfOQ8S;Ab]d6cGBSgSY^?(#W[L,^BfaQ=V0X)<D0TLCP9/]Q(adN]<)AOZ
?XMK7Rfge5@P3IbGL2LcLR-V42O_D\L<IKJb3I=2M-0Q&bYd(42W/;Hb)O3@CJX5
Kb>U3HLHMSIb:5L\,bWU3.3Wce&X9IS)CY&\ZdJa>66;4Z5/Y?#VN-8ZaSb]fcc<
<2FbZVB=XRLL>F0/-?JP-Q@ceQPX6RVc6(2QN2<1HF.V1T_g24I,QPW8_T)FFSac
c_]\7GKLSF?c(Q9FFN;H+.a[Acc?.VA1P:Q:1WR]=GWO<P]^W9gHB8QH3019\TeL
ADYV\>7.HPbPDdS\MC>gS;,8M7IeRWW1/(0(9XV/JI1eS)K&f8]WWD\BBE:P\.)W
9PU]XEX&#0_TPG@?YW@V(A1L)R^8975a^9@AVF+T(0W3Y;O]=N=#9I,bbMB:Y]d.
6HPT<R5-95fH^?^DDLNN,AO.N9358/]5\QFANVX#aP499NFd4K:H=(02MQ]C<KQ.
Qb:WKUBg819a1:XL7QaB7g?RXNa^8&ZT+V[0\VJ_^&>D1@>IA1-f\<W:#7:bO4(d
IC@cKBG(7d_9DH6e&VY;]\c&UPadRT5cHI3Fb<@1&AVfT5e?8,1Y>H,A5F[bLZ#N
S>L/=#Oe(a7_8\_=?^+\BDJ)V=:B>-9I7E&@J)b/^C,S#Xe)3NZ#Y7GHMA60R4;H
fZ,g=6;#?cGES0c=7V9)Ge/4@HMZd&48YE1A;=78+_V:H(NDCAF[#.-@8ZY.2)dc
<TOd(8H1&=]5Y\0/B?bX)f=P,G)3#Z4eK:]C0<J@c4;C=3.:Vf+4WgA+dN,-[5dD
95(,(2]4_ODXP(?KE?86J1d09a-:&8<4G/\;P^eFT4eS0O(g9OB[\2:USCI9,<-(
?U[fL(JL1U&G74CUPA5<&T=6O2bVK78?gLe7WRSY:WPeJf\TBRV([KP6dWa.D<D_
XN8R1^Z,b9NE/./RB.+I@A_,;IHDO97.S#Y.8S7>R:g.43bSP]/USGEV<9BKO.V&
CF\a4O:[#VLg6Q),@;\<E?V,d[=gTg7Kf]3d95TTOE83FdK#D/;4DCZTZQ1=62T,
25MIV=&1(Q9.@/gM<GO0PH&.7#(+V[/=ObX+[:dX+/17MWb)4<3bcIYD7Y7\WZ[a
aA3dJ0gY#&]GgL:HDUQS7UFE0aW+E&?J=]JNW,M0DbHUX?U7U,]8dfc1OKC1Y/&8
Z:U9aSGBURVPE^\>DMTTHaA-L8:D#4<8,,;Q1/I0E[e44_f@fD7U@1VGRFYbG-bV
eJf@-?3E(O=G7;d^g@,b^/^R_[J[:BEdT7SPab.G^dU(_d3.MKd<1D6bK8&I-V+=
^ME2ZDR?H,Ad8].SgU1d^>-3/0ZNL-ZW#IeI3</+VE:]V#HU3@^6/dSU#9TS?W</
fCPPf&.V82VN20,Q#KJ&H;]1Mf>I07(Xff+^>[L;ML:7,)SRA_3YDLbQSNQLbb^^
11&Y(\IPT@RVc5T=(+BA=OOXKF(#6F4R4#QS]U;(H(?[(^Aa]dJdYMHU7/@79LE(
+(B;I>[+e7c6CHF2C=W4AJ2#.E5::fDG]],#3SI&K_d\<[[4,S.1:3<[\#gQ_]Ya
1=,&KcXf[Mf\+cB=(&MO#WPLbc#X718HG1S>Gc\+@=[E__5@^,7^Ab+(4WQBFc7;
<5N)87,SKad2;Wb2DZ19W4F=2,0AgOU01B2XDHAeHF.\V?XG54@D,6&Lcd5UKFWC
5D(>O,FIH=ebTUeeNKTeF:U8;Rd1DUU0D_O\/NB:)HC58]41R1N+E3ZH;D;2W>bR
.#<<F4a8=_C50badXeT).F;UQN@H,=F\(D\7AHY5I:BWaSf82Z3KQS<\<-IDJ@.0
JZ\Z=;AeS/Y.YG>WLVFX2)gEdeeCQQ;Sc/H?D&6&b.MCJJ/W-BBQN=Z^:G]c;Ma1
=EJA/IO<Wc[]bAW&X=+-egQBU4?2^0==XD/RNIO/bG]6:EAW&EBI#AH:[G-_E<g?
b0MUdQ,b_<,.S;4Z^S/DfYG]YJ>E4L^>&Q#51dK^OA;PKQME6.U<C\X)\KH43,BY
(39&@(:#_5KXO,L9N9W,U)\<\=RcUV9^+2-^9^<e4c<c]72AVA#?@dL,4\2K-&RC
NbFIA]=af1<V/>dELV2_bW>&MO3^PGO7IZ/d\R&6:^YbCDA+M2dM:Y^8QIZSN&eX
<114eB9;FAD5Y0O7DH_0;F]JPPe7YaUG<0g)11-H#PL_76/V)d+.0M#K;#DP>]>H
-a0\-WU@CgGO2g)DZI<f7?S_OV3W;)L.U1/WJH@Hg/#PWgRHU,OTNZDE?^HMAO)S
GQH):Jb6ZCW7I]_1e-<C=-LK7+cC[5A1H74J@C7A]4=a:NV8]KZ:&[54HS;Uf#Q:
)OPP_XKDeS,SM6)e#YO,bHM:D4a@NAbadZ@+8PCZd#CX6PcM&9N5D+[6\f1^H;L5
&38,UVd)ACCZMBQ/SD4[E;eHJ#N0KEF2]IG=aLTHQX@-UA+c6@=We4.VQ=MTDd<a
(3bBM9[I9MM[L^90UUIM9\bXAaFN7.RAdG/SYEWA[U:503:O^C1=:7,C1&YMIMWJ
R5ZU5<;77QAB&,1-::[T;/B<CM<0VGcO(_g-1ZGf8-Wf^c4KT1Y]?Fa\OHU<4X_4
QBDXSN4I0XDEdN^LZS+]+LN]CV.N7@J0T/Ybf>+-&Ya=[EKV80-BEdQVEA/83U8Y
C\7;F04IZH6WFF\+W;?1W:eDf,W.D,L_YI),b.[^I5@LW>QfE3<Jd5DI,fK\;_^2
BVQU\A+#;^gH+).]4;<7H/VZ4_[6KK.V\PE\c[RO\U)8\ZR-HQafR:Y:?/L_g+VL
OAL/<]B6UdL.B1-TOR.c4)N-Re<6F;],RWf:f_gSJ2[7_0R80+HS9)<0DY@.(d7e
2EgHgE_51KfHB@VYFPL&gAK/H(6]deB8]/#@b(VM+[803[0e2>P#MbZ(-5Y>aTC,
^VT\_YTWNa9,N>0CM=RC2T4U;Q1A@AA>QHGRQ&:(ZBCAY(]Z+0S2#O?41:WG:^0^
?aM?^e?;)P)M\,K4BZ\60@F^;)a2&>>Y5>KCeBf,29EJ0_4T55AQGHSOg#-Y\3>H
AT==<>\=#R)I=XB>dK]cB&5A787,a4Y:>+EgDS^,8N/dH)g_)Cf[Q,GS?4\+0OMC
<9RU]5-DAT3gL&gFWK8R-;_MO)F1C3LE()gGa^dEgZIU32KBNbWYNLE(HfPUaaOe
;G,71FgcJI.;R3#Q/OAS,1MPV,MGdcFGbFcXWT;E3\8U,@3DeQ.cd?C;31eR9,QM
MW8PKDWNKZY63H1Z-Y/APQ8P@R;_0?f@;75Df3NIcH07(//CGgefg:E-5YFR.a.:
954X8DHQ&SdHZQaO^:YZMLR:\4\^22Ia(gO[YT4)]b1?+Ke4UN9aMXQ&_F<EV\X+
0+SE@=X@=:N^P_4cS)I#U8D4:YAKWFSRIOH)BNU=C[[/Z+Y9V?_O7V;3ESJ,gY>,
d;R863=PGHF:40ec160^)0McL]c3=<@?_;0:db/ca7d&;.Z#2(e\O+AN8DV)3@Y-
F76LUKJ;-NM1W(SQ4AQHPV2?QENSU@6NUA-=7J99:T6I2g9N^TWUPRRL>N6I9gU>
Z5dKf):X9ZKHNE>GDWg3\YR(HA5]8JW(U&Pf>.2VaV:Q^6dMF1FgR7@)/V>d9>6(
QPX_L\bLWDN^JEFAG-Q/+OEe3TL#)^^78.UbbRO?NT&)4@Gb8b9MVQ=Y^]MWcNS<
d:LAF1eSLMYM[I(=1C=2+OHg-a,/dYBb]TfY#3:D483BHVY2\,C:=:eRUS&G>NZ7
41S1cG1SBL296(Z#+TB&Vc(MVNL@OT@FUd_c>V&f)AKZdZbO\?PD,X^f[<CVZE):
&1_JKg?aL^?+V#L#7-g#Z>43fSRZ;<;2H)BD2=V>\\Me.(-+X+R0+,D;cHY5>?1Q
AIfQg0GON,gM>f=VI7WJ@7Q6M8NRA5>N:W6Hd_+N[QReI[FXg^VIE89V\2WOUXLK
E,[.(&C&6Bece]1>LI_0D]T@.C^8_.SaGHJ<3NZW>^=)FPI8OO860a430_7KVU1;
9D.2=1P>5,?e88-)<CB,?TbVO=H/NW96DgS0+TRLQU4RdNVVUH)BM#NB1a+effRP
dc?4,]gCe(+.47.HgbN4VdVG0S_7e@]Y@6IVZU8_SP<0@EK3V1(PdLL1)1>:YVY)
e73NUEV)W)-/\C<2-I3]MB=Bg(5@:BDL=d.63?QODENN<B,^LM5gH18^g&+/[^>N
X\_-R?:E^12+:8Xd43Z^Z\eC56&JUMP1O]eU>S.R:H<G6VJ/]A9)L?PESF9&<#Ma
=40IggM4H#HGFg0:1dJO]A60aUY+@9+K]].TGU5>9+QQTSZN&JN19c0E^1Rc0V4S
[Y>X>.\,\>DZUQ/FJA,IQ1QDEgbRC2d;/G&TW3PA/;&SZ33g/&Ic-Y3ag,IcWdR?
L3(XF&eSEVM[e5?:&QUe(4/AOQVZ3Q^_6:F^3a7LWd:KM?:ddf]5D:+C\@=0J=:E
)RL#0XBR7X[T+X,IcR3<+VW:A02YX=\H9aVXH_T9a)W536]CZ-Z6=aIXCDRX1Z8^
UB<B&B3OA>AdQNQ#X#MG1g@P=bb6^LD+N+3UUI/(Y:XAb3:YYFH@9RZB/,HGgO?6
F2IcK-;&(ZXQ([@U3+YL@FSOeRZPOI@,_e+IT#K\F1L:PfbUZIg_FNMe^=\BVGHH
#&aY+OSFa(U(,K\J6+a@C_a#W6,5.c\]ZDYT,SW4.=OQ=4[J>W5VdT12#1.?E^WX
<G[LTNg[VXd&T@[;KIFXg85NcTULYQOOKPN3Ic/UGAP8C35g367SRfV8a@,:UM@^
,+Q1\BEJ:MQMH5[3;g4C;;cI3cJ<(CRIb=UTM>?(>T<BWFJKB0.G/R_f=8];C6\\
U[:3UA78Y^@Ud9J5\\)bXAYGJ7LP9-?>KQZ746FSUa4@Nb?d=>8fW]SN=TB]9=g/
:J\KU1LD#_FZ0PH^1[FX?F5<5HO\(fJWEb?-KWP_P]_#RJ?a>BEA[Z,8V=GZ,5EX
HIG(I(H&)1-dP3#5ISX\(U.);USVZf0d0JOC#+079#e_T+?39S=)/CMN]8;@?;0=
#[#Q&(_9SA3)X8ZLR]XU=V58[9bHCVS@efB6Ef#4F+)Z-b&^T=4F/VS&9U^5G=Qg
H5E&-F,OG4dGR]3QY=.g@TJ/-:7B+5SF:?Le)F^VBeY7^;]+:B;G\YZ,7T,LBH&=
B2:ZE,0PXC(VBFLIKaH>V)S-22D&&6]6Z?WV8&g0cQA)b9bb\6LbO(BXQ/A3QgOF
[;c598ee/FIe.C2eK,84)WP1/0K<;UEb?8JI=M6ecND&XD8c^ede>XgcNE;@d4aM
LGIN7DUZ&,M4-+cbC0LGT[&VQUFBT9U=Bfg<CRY_=Yc9\E,XDDGT)NFeHKH\QW[X
c#XA,J]X[CMH7S.8XDV6+GJZ#OW.>eSKb@<[QQ)Y[?W..a;K=T?&7)Z07>)g?:B-
+(8:RSMTYOD&VXSMa4\1;MUHO3>&KOS=gbDGM/:&.2/)3CW<_ZR)BQ@.>+\NcV;e
Z@IHD-J:[,NNU:8a^S3@D]+G9TXN3Z&\=_=Y2\]B6I8WdWK-;D#>aPSPN/fT/Y#(
U5?FVP_#=2^2M<0V[7IJU#VMTL6:SbKcOIF&43Q;_:#R1BA+@W1IOA#JZe8951f@
V@/aH1&4fE=^7UDVbgUNZaR9>44+)OG;J-T\.,,2N74>K\X&F5#EV_6M)-^(ZM)A
IbIePag9;dDHe+S.f:6dd2FY;79f=Y+/^I;&VLU:+c[XTgF=;N5A?615M_0cMVZC
K>8;3FUGS;d,Ef;-N?G&Y71.\4Q4=JfT#+3>Z-d)?U7\BZMC&MO4dQb29)JNPXFW
[]-#UCS?3T.Q<YA9XU8_S@D/:<e8Gb&@5==Z6RReG6EbHU4Y/Sa)R<Id=81;?:GM
=1TPbOATeOM)9Z0aRg>aUPHd8QGE9.I5:J-[<;:H+&NPJLU8<<.XegJ[89GO#HP/
.DC;>K<Z?WOKCVD5.<\0IX=A:B,AeA<U>Pb)@H>[VRNMJD+YB1-YC1b0@Da+3.-0
EV#@&V-TbW\B@[7OM0V:W+g25\(@DB4Y\8HYcGNK+^)g,f>S-d:+391V&JN6>JcA
RdB,Kd9X@XedR:,3g9755OS@)^;=59_?RN:NEA3R-QUPV-JWHWPJH(+(PL;X/>-f
eO#7XcbBY0Y5EbKIP7[?N-)&/K:8f)]f]\c@/f;-b7Pba/46U]B5U)>39aYN2DE+
W5GC_ZeG4P)_gI#BITK,4cW\f&Z]C4[gD7f-H1a=R(T?T,E/G\:Y<K?#FbOPLba>
aVc(8]I[<3>,ORe5R]LWCg_TJXXD8+<gJ61SAO9VIg&IK4#+7bI#)-H\83&?F(_a
M.08[91UE<_<ES(5?@85N-?DUa2g[F#I@,4X_\d(BZR4[Oe^?1WMKP4_WV-QW^Gf
#J#L.CaC_9[#0I@0dce=,,cf0>;aEZ_IJ-4F#KUb7Mc5^_7bCUZc7.L^GZDY0HGQ
4#;Y9KUXG>D=4A7CTZ7Hg09)5,DU#-W=@BWXYGBV7^/DU6/5.S1K36-Ab58&_&ZI
2??UPe4bKf?WSFg.3OT:N<ZOBC9BR22OG\<QGK;QXJH_a<024eG<_V\U.:-OE<[Q
e2G;;<GCLO7)^AgR221bbUFE2UE4=MTV1a#CR4]bN4Y2^AXV)A#.K;L)G3cbX5+C
KNaD,TFW7]B9QCU+R4LURHQ3>Y]2N9)2ZB6B(G6/J?Lb(cFbW):_\P4\LGN/FQ]6
b8NZSF>J07M?)Q.?+2J.2BK:eOU89\g&QAE4>JBe_07UZL1^Yf)FJU/):P:?6DKW
\U_dT=#3#7Lf1F&5b25M(<QUY\;gg[E4\Wf?\cB14OdM(+GL^Y]=[N3X:\bP?+EH
3dE-NXgVY3Z@aa,,4E=^L6B;8SZIc05+Z/L=OW37\<Ea#-3-[ARP70E[7YF2;eRa
6;HJ3gQDZ,<HN/92c->Mb:GPYf>^U/OWIGGQ#FR4QS^Z8T>fU#]d+SB<-gJ-^AJ-
Ja,H9?4/]bGW[GZAA9Fe.eC,KLP@b1CLRfTe[a6TJ6K5Cfc.AG8=S<?8/)+4IJ=e
SN-:+N.UZ/8\Q+ELbHd=WZaEPd;06GD_6Q+/ZZM)\3_F/1/NDF/F/[_PV/DXg@I;
#,&cMcH1W[(D47SeL?gPeBEEZ#8#:\-#/;><74g@Da61/EA-?/DUD_a6;0=(O7#A
LDO^:b.U9-gK&fD&KW<1C0fI16#_=WKZ]Q]Y@-FeQ;Sb(EIbKXgRICfU6H5dC1WV
4[WMJ1.2T+<5).N:QMC30_S:9Ne]#QTG5_W2SU]f#&[5O8>M+MBW>SLZPBRg/JDQ
IH2>4=\5P^;0I#=Q/8BS[FEP=B,IP&gYBc8-KET,g(1J9beHd^8>Ef9ACc[EVg1)
\JC<_a#7bJ8@HMId]]eX(OGbBFKCUE9^.CZB;M4_<;.aX1d+SZ9aP/^12FPNAQ]G
a0\N=0b879WNYV)6aIQ,2@W+9/)#+VI2#b+2F#I-/@WMU/&H_N)D]V&IAU8e0?RU
cd;XB[[N=O;BBX@+7IdP=CXWM[KL4g:@Be^LD,T##USgI0D)75>c,FFeLMNdbX[(
GMQ2UC#aP,A[\a5F5OAeA3-8<9UN?c]27Y&L^;b#TeA&/[JX1(XWLPS-@2Pb2QG?
@7QGED^51U?3g^,[//-W#baD\&<Y(4.SW,=XV8PDbBFYIUU[^EDJO=(?8GJL7#\F
H)-VD.SN.XgRMEfRYY6-V@dMXCcG#gCRT^JaWb6SEUC=cbU;-Tc8MLQ,c;,9Q>,5
gBK(dOg5d2?bF)FRQ4;a)SW^/fK.AY#0+1,AM7I+4OR\7;aX]BQIZ<1Td#JBdN:?
?A-QM\4=.->^MWFWBP[)&Ef7_eZ,JC@K,eYegW\I-MN35PB&@9d&Te?@B7fAf2_[
\UP3KC2BKXTbGI=LS#I?O-=+[E(F5LU\;POf].0R+PRA<E/[L[cIF37M91>FAB:,
2a83T(QP#[SW4bW_2g.@fAV[D:d\gBK^3J4a[RPX83ZJXe7\C.YJ7\7KHIJBZ:.=
&ZQG9RdX7gDG1B#YV#GZIW@OPY1??-P=a6AWI25>c-_b7SR5=JGDedYHAG0fD>.8
9/JTUQ);T]0-^5=9dJA_8FO0SaKMJ@WSgE\SKR#:N_=-VMP;gJ419W,[\)N#7@#g
M]RIg10WCM7SY9RT:#/KZb@gX0H,6W^dC\cK:<BW^PJD)8M^8Z1XgODb0UW6#OS2
CF&IGSb<+,cN7aSM(HSJOFH>BBbEe4SgaFYE5/b^]V2H(?JJ5F0g9ebcJ\cL7WUS
55g&AeV7X;Z;Y=P=LNM\L7_KT[I#-(VWR&69ZB@#U8TDgUQa6ZVX6?\_-[-1,_;B
FYETTXSFHU0[L?>f6PD=BW1J.#QL8gO=:R8_\\DQ/1]^2U:D/Q:dY#OU754A=g(d
TF^b&#+\QZ70@1F;<M&CNKUOM?M?JZ@3Y8d=1MKGL?gB/7P&#&@@,0R8Z3O?N3Rc
VJ_8_;<XBFff9gJeE\^H.\Y0cd(@IPR6ZL+eG==JKH9I.>O:KOO8=IaN<BX-#3/<
W0E[S,BNCad\=#A?H)#C.EIUf8U@]HLO0/NRcg;&\4.Hd7/^QP4W3+S6M)O_bf>#
SZ9\YC<&JU;@Fa[WK--M[[EWMR6N-;b^;b?05UEXV]T27?(NT11_C2eDXCMS&W5c
7^<1Da_H]C@[_#gEa70CPMeKCP;\cC+ZY,;W7DGJUGgJ^3Y6(X1SS@Q](cHbV)/e
4<73g]2(^1=29.Z=E[c)J5N;K^+,AAgd7/_1B93-@.2718E/dU?H.C=Y9c)G.aRc
ROUc).#AW_H2:]PG2E5^bB_Dc+db9a+gQL=)9)RF=[/W=8KYRC3bM?Q3(&ZQ^QYQ
)F@8MD@RIBNT-/Sf2?;YdMW)\,J+.CX,+4=T@eE/ZgI^<RedCB>^TB0R7,DggZgM
e1^fWQ-ZY=M))I^H\0:Q9B4?-QA;D2NcAIS9MMC81gK?.CY>;0]N@TbdZC=2OS8F
_L7<<F4bg0g]_1C8(dY4(9HXb51]17L?NSdK\RX8#_-@CfW:^b5C<LGT@49TT()Y
(bH&JDegf@^1D2e0..cc>/Fc+/6Hb(f7;:Y5#=Y/dbaMcVEY8e33gC_=:4UFAR75
LdT-f@[M/f4d9[MR@S2-4VLQF9M8ae#RX2+X_Z=+c\fTPF^FbH)KebMPK6>7QG2G
WL,[GfR9D76H0\-]:]8ZSI#UFMV,T7g.e0ILA1RXW6.+&F[a#Yg>@#1fKfCS0QP.
e::Je?Q7d8>IZB=D>Z+/S4f:JC<13++/M>(M@H>=Z8M1R3+ZQO<6;1;8GWHPVP:K
RGLZ2Zdd(X^If<Z1T9c^YUJ?86QT7_]9NY6\VN)@860P(\X?g8.WZTW_;^&&>e4-
A/g&;2]=c8C^^aG<AcD:GII5H#S&=/3KNd/0:5-:[(W,#[=g&5=F_f0E4-3?6P/N
fX?UBCcRC+B_YU5T/3G#SP.Wc3&K[DCeAI.82BGU<FWF>EV0GFf2@L;VM<5\@52U
<WA,L[M;V4+)XcXA).b]W9Zc/Og2KF=OSR9d^Z[?3M:FZ+2g@2@2g==P#cU[7>RR
L,BC&[S-:dLZcVTNDA_&;RY)WI+D5QIIeI:C@?:5O=#EEG0Q:W3QK>GR],T#E8ZJ
<:L#_S<S2Q-:WV,Z<SPPREY9?VPH0JBRe]>T#;@8HUa&9@0d677ZKVO?FK/.,9JE
ZG2IaZ0J..Y8<,-/E95d&1C=Ve#_2?Q7c7)&YPVDFd--?eN32\Y+fX5gadBJFWQ-
)E20_G0:SJ0NfeAfHF8C4g4edA(CDM/bSeM,X]geIP[CS&?V\LICV)Ubg\?af^[,
-U0@HNMBgUHMLbbONX4gFDHEC\c&]F<Y1PBV?G?L[NL3eJ55=c:JXR.&-F3N;@I,
:D18d^@:QGe#f^V3GIggQY+I/W+G(dS:0?Z(dBBSGVa+d6/HIVI<#c9c9^f]:S7U
;=N_(E\cTc2QS1dS\62=]5W[EV_PW-8;_H4MEBP59R3K_;/FB4I[DeHMK)]1>MOZ
-MW]R.d&R>9U>UWG):=5Ye@.#CM<;f2cgHbO+LA-dCE)ee_E.?6/6SI;E&<AFfBS
Vg?HaR\3,0aU#.#1A4bH@W1/.e7,fH\#DY20EcdI#3[c4&I@>7891eVA5Qf?X(^L
_V0,:N1R]f(DJXGM3].H<VUM\c?0Z09-3?fMfH9X1f#WJd4?I:FEfaPKfW_PUW0-
:D&b=R2gg?#M]Q0a/IHB#9?0;L#38KU6;dTZLXGQfO5@2<>cO_U6F9[Y?65AEY<X
BH&JXZ&0&eL\<b:(=bVVG/AZJb/43L04fC+_1dUK.?BS_C#[9W#R(X;W+Q,a7FTE
+:\gT<_&7P\;I]@:^CAUDeS&b_&^PPXE<G7OL(V;.cCG?(,:SbVVSbU#(7V2BD?Z
>FU1.^gS8X]X[@#<e&gTN^_A5R9G)>EMF\1NS2R9=(Zdc2dQD:QSQa=0EVXXf.dX
(B(/d.D[KN=f^QLa-:(3GaTL&G08&=(bK4C_#5@>.KFGOE/J)SXZ+-[ICH\BK>=&
0@e;E3TY9)HTF#@5XN;SVM]N=a@6?69&g0JC;53e8#.?VAa-DPWYZ7WI,KBR[P[X
+f-?Mb;fPVeH:^M#1]#e@=HG]8Zg6b1J7\@P3[gL/J?gPY9gSeSNO/4/Q.(^>(VX
e#1AdTP3HQS,DF3EIc22#,2K]c&M_\(-<Q?e[(&ZG1Y;bc-7da-<F[]Y/KfO]W26
dfKAECWV[cQ]_]?0YCAKbG@(GD9Be)0AeEYU\:HU)Q\(0I-cR,:[#MJUK2U(FH_]
4Z^YND9P_Z/fE_W=.cegFIT)0<A+49=449&6#IXDGVV>+3g.+3H3L<5-72&ZO=BC
b,:O,>)[?@M3H=3-FX;02PZ8-NVcf\<^2<UR3/X3ffV\I3HYD=-d.:D>&aUV/2-R
S(.ED:SH0f/<?&V(K;_0UO[R[,5P(262]FU0aC,G4gdR=KMSY?b+\7cJ+-7ObWB_
RfZEc>#Odd8@?Q4Y/)XJe#>I4]Yac\KFTLCM:.GY8=c)R<f-&I;F/1,P[]@B1N(U
HXCDb8[+ZZS_)@@/UIWR<E-e753>>:Q/RTRXJ967?_+92FNM\O[)7CeQ^3,6AaY1
(9YNU\cIa4R#3Z55>P/09a+(RF\U,]R/J8VJ.#d8GRN+HO[8LG)^^UM64/+&B_I&
5]&bc[VTaW5Y3<[R5<(>0B;VC@J68W(W)dHT?)LedHPH8Z#ge]>FbK=)bO+&VM,2
_2JEd51;1XUW<Z80E-@XM5U=SZ[4A9e\ZY.Z7A?<0G9ecJ9(UPX@)N&?a=\#9=?C
BM<V7O2L6UX4a>)^C#6&N>AQ#3dDBd>>:X\6=T=1:6e=Kg284Y,4M^TX.;Y+&cPY
MZ9O;W#=?J84<6/?,cfBE=a08@WEM/f-,V]LNJXL\GBYLHFS:[OIXdO7W3J4bRNb
SYVV9]PKX]UTLT=9VG:>BQJ8OV7MP01dZ)RB4+-CKZYL&L8U,U@GMeL4\HOK1-_C
QWK:6VW[4Aa-G-<I]f.]D6;O2M2GV+3SQCHfa&ASV1=4\/Z8-E-8g[/T))Ac\fe\
I2M#M?KPc.G2:XQM#O_9QFF5RS^NJW0)cQb3FWLEIUJag8^HIeJR96Z(<V/B?6@0
&8H,7[C<61b6G]?M,Y^X5MM.F/7=OEU(bdI<Lf,MKZ#WHe#43P#G;KcD6QJFL3P6
G&DD>O](WVV9J,Z8Aea>6^JQCVdB4_]=J23L=BacLaVZI1RNDOXD1O48)4B=Y8?H
2<0>-O<1Pb0R0gLf-CJU#a0NAPYJ3I20;;.X\R?&)PM@FI^bXQ7a+bJV?D?dZKHG
c/-2V7/,5WG#KgUc##&Q0NI?S.??V/T-3(2FVeMPHe07XC0D+=ZO3WAI[K>a9d<N
g[V9<91UA43L?b3a=g2Z>aV\(@VQ\JAdE+K+YI,.[6_)WJ0>6e@8A-;:S#2YL]a>
Pg#L]&g[aEeDW)ca7,ed^;-H.@OC9fY==55<KLe?eB)ASc1<X7-T^d_BfaR;L@S<
PINQ_Sbd:4+<O&SM@9_Nd=Q1=H,KE(Ag6M02>&@-XfV?(10+DE\=B<cR-G04R80H
C+Cc,17MdE5@:90HNAPdKfN<P@_Z/f.I\E,/JXEeS3Gb_8QF-4?D>P8GT>FV+1:Y
5HeC=V3;a3JB=>X?;WR#)CWY9cN:5HM1[C]3PS(HR>a.:V6C:^QB&\L9BY@[61A#
NAC+ET[G.Ac0CW04DG6NA<cE-f=2MZB&.;O,GF7Ge)f.ESOfHf(A23L(fF8]+O-L
[Fc5,7I?_;&N/OGEgXc=)K)40XGD[VEdV:eI^9O=J]SXeFN7S\LbKO.GI80?ZS,+
F@W-A\2D)_J0KOB-)JBKNN6W^4b>K53E/71eYL+I)XdHGSAZSCP[7K@&))fJ0>/6
RGYDW5g4J\J-HM)H8DRa,MWgL4>0GfISFN?DKWY=&]]01<:ADV/+d&a@^[6gV5G?
[U5U_L68+=f1/3.Ob(d@D&4g44IJF7(QIQ<aVLZE-(+79MY-AYaa]g=B<V:I)0=D
9QL\fR)RN0+W4O]?<\Y:+YN0N6U;@OfMU-V.(WdQ>AEY]3DfMK.4<T4YL8;f<B2F
BbT/]f75?R#HC(LS&2ZDF4bH7K@M]bO0I.).<DZXW;\4-(,]NeZM7cE-Qa3JMS,b
PNf=>(g[FffFaHYbM.<aEOf)ZR[\4</3P6=+;H&Qb[f_&JZU5)O30NN#^3EeeLaP
28)2bg3C,4O.>W:f+AI.T;(aE92EVJDMCe<Q2?13(?b-GCf5g,RETCd]=7O@>Z/>
W^OJbb)7J5U:7_+_>9,]E-1_Q\7ZN_dJgcEK?V[g@UHII2FH:-Jb@EL9I)I2>?O;
CR.UO.a_1DP;8?/N7D00U=9]BcZFINJOb=LA#6O#\SL@DK8W4@+]>MNAVTB13WC7
+:JIR;.Da7UYUeeS&?4PW+:aX)dNEc[CfANaYB=6EXcC@,675G9Q7g:Z9BEDU/8G
UEX-64M6>1-;:]93O[\c<dfSP<6JVDW#SRYAYB>:X?56(?ZGX4.B-^T@SV7P8ME9
588HD/VL<gP(,gY-c0HF[&a8U,/Wa3(cXB4F?]aW)2O[A8BfU3.+L?;cFYa6.WDg
8Nb;L+40<SE#AC&&GOULNJNX3cP#eF4X@CIZVFVTU&:&1(D1e^8UFJ57OW4;N&=7
.5LVPS/A4[[9D[.SI()SS/D>^8_/OH^Z0ZJ.G,3)PM,e][VEV/=U6>Q;R#gSM7JE
JJ2e:EP@E4<G+NIF-P+&\+RV@YN_TGWY?N45Ra@a>(fV(Y2#Q1^/PN-KcbF0<)6G
Q:,Ba0]VdEIC3ff]Yf]=E8975SAV4VCdZARZTAGD#0#fDWH-BWS@-]8=E&NX8JQ#
,\OK;/H([E8bN]PP.PRP5>d\LbPeC_/AUGLD(dZV;Q&1=8TSe=)(TH^g59gEQRWg
0ZNC^>TJAD8/Y_</&QJ7#]A,8+I&?D1Od+T2;M91T&+8UE>(PO#Y:af;2/-+Z&B+
KaYL/[?TMF:dK/,093EDdJX2BcW=TSe-Yf+g]OWK>>/<M(M?)OgMW[A_V/eBPQYb
db<LdK/A\8e;?XCSM#/=^e16+;;)PTB.+R5I3aXXO+[&9Y\_-<A=#g00_:X7B9?G
+QBUSe9(>K,>L8A;?EAXI>].4\eR2+:^<XHFVFD3DdO^3R2<7QYX-L#[9cXaTKVS
f8>SQW_ANHHG[Rg6e]J:51&2[KLR[IDFNH=#RZT=\4)KaY/CXIaDgTWS)@M^/R62
E)N-=f_?U?Z;EAW?c,8e]Q(,ZfXgX>gPe84CBB5X?N0/@B=]>4-:&>HLQN;OQ\<[
b4<LN0KaU6.CQ?+/P3BMV/N.d,5g\6Mbbe39edVY:/9@_Y(?N.J9[6QTF).@G:]X
:2QL<:=98b4b9(+PO82LMJQPW-<caf1ZE87Lg,^b56GC4&\OZdUa2eDc7H2R?1@P
fNN9H\(J8]KRMOIg;2ORGG44=dU?G9#8.E=A/:Q7IJ0O[^e5JDVGe(YL?IO7R<A@
OJ)LS0Vd>0D&c#g4KWKE0TC1PXd7_N&F\1+egNX#O+3;^:[2bGI8Q_M=Df[\NN28
Ma>GF+^.54?e@@\#]]PY:/2>83d;Ubab(/13@g5cHfBe\bC68O8e2g>IJMGf</(7
NNb_RgL9J+YOfbT4A[Y.:C&c)7bdaR=JRIDc<XgC-.\=GD#+LYRZ?E(.2J,LGDB5
1_GR<UB;,PF.Z<T(=_VBYV^YWcS]SJDYN@UNBLS\1A<Pf3RVbH3J8XXf@d-^B[gT
WM)QZR8K5NWP7CKMUW+g)36U<?_P(&aL=_=[.+&3/_ZgM;cPS7Bf:+S]d8K@?eD#
.YU5MAVS67X3I<U@FS.#KXFS^([/,-O0[R#J6M))>8_gOU@+.[2O(JZbSMT@O++1
GJ&YA7[Y^W#)\dTT6_24/]Af,;V::>0D7^[dKR(@-C:Y.,B@&LT@>K[\4^B\PASR
C?<P&S[2FCG4OQ,?b44Q[)6,.Z35gHQR2M0f-N&EB,W?7,)f?JO>ec5Vg:X7Hb(,
_ZV3=:4SP\I-^8,e[7K(e@g&JOLHO^:f)I#PXB1\2)OT^RbgF]ATUIB9TgLa2<L/
\b1(.,>d>>#:T+_=K\[Y0Re@0]-[S(,VHSP@c>SPWS(5\abE,gT#F\7OR/7V&GL1
ZT<ZKaQWd8YK\(/4@dAafN7GF[1UM;V2#D=#E+92-([2b92DCIJCg0]J2^A.CS>\
/C]0;VY0VIZ>D-T(7GdG./bL:J\cLA:FcA7#]]EBPFcIaQ2D8-FH1(>F#XRUU4LY
V,8NX</@T3_RQ:DDOY7bZZ43R4[e)7dC^]5\+W@@<7dBaDGN1QBBJK-aAJ\gPC&d
Q2(?SI-2T]TWG]64_]FXW\f=?7<(U7<2?K@LcD282@0LNM#>Rc,LWE#7>V5,_4>&
:(E^Cb8LI^RJAG)TBG8FI@INAY(0QSXC=:H2B[\32B20()W^R9^E#E@-:#+1RA.Y
aA^J2+@4U5egf;bO5g80EPcfebO^Mg9aBR=:DS)5;W3bME/E=69;BOJ1J+AH^X&L
._a7GJ#,J>caEVWXe;e]_?gO99.[3MPX9XSc1BHQE/>HRDfCB\#ac?IRNE9J=f2[
fac>\J=33WG?AB&L4ZK9E_Mf10G2CG,fA,Wd>+d\A9DQOZ#Y(#Hb97U=4S+Iace3
eMg15:&M\F=a_^2g_a4H4^727P-g9;EMb.UZWOIIcZ4e2V\^XK<SJ:,bS0&8.AAC
GOH:Kbf.CZg/[CWLDeZRbSX3A18XAHP8RaZXbPbF6H5P9,Y<g8OD3&bbWJBSE2\S
U7b0Rf5:_[NgadDI=F3:F],85ecT114C7\F13N)49@decP,WJI#LE#UBP2gJ]-.W
0CVXHTe=&[)bL-?dDW@Scg-\G138T,^/9/ReP?7R+<3L_eNY5F[W2Q<AN0A+7D7^
UL-OH@ZY\f0e9G-gNc)GU93?1>S=+SC.DI5U9MZe6<:b]]0EU\#8Y\aL.^VfS[_:
-;=.KL&+,>:DV-8WfbB6<Y3GJW>8D@QM&]?<H-^\T@+20g>.0KI_03)ZNa=O2f_,
-?XQ,B;XHSJVP(Z0E)A7CeJ.C?70XQ\,50V<V[T2VW01),0K^XfdHF<5UE(1Sb1S
Q-+Y&<fDOU[[(L\LKd>dMQ\.@:+48)CCPML_94e[V3D.4J5#Qe;)<:/CX=\F<?9P
>HR)^J.e40AZ<DXGA1QUbL2^??25-W<RF#ZB,f]c@.J;Bg6R>^[,776/ZFg6d6&_
f9Xa,T)3?>FDF[U3.&4D.XCdF[GDY)F#HN--EV:T3Z^^0,/K2W8.4Pg@Zd@708HG
=g1>]:[R^]R/48VC_]7]##0Y3Y/=\>3WS>OaPP6-E@Bg<6,D\NP@C_(2=.EARJTS
&.N_S(,NH6Q[(EAU11MS[T98XDT.6F(L>7=HV=@F(>RNQU4a\EF@R(A?@6Q;)@OT
=(^GWcA-cZA&MHY)#Z+QfU6]:XV5Hg(54TUQ9KO>HBXX&^[Eg)IR&;W+(R;IMaUA
BO&^5T0Y,H#V-LNId(O+5C=>_@S,]9_>c@Q:(fg;D5^GU)HMJW0\N+KD;JQL0.@U
Ngd8)X5gc9fZ&>H9WSf0RQ\A=EASHSI6XIKH4J.5UOY6?TMQ3W[.R2#E\0-YF4X&
bCC;dBD]LM05H3)DXWB7EU:E\4MB[&J\3P,[]X5#YN+?3<>::Z^UPB^HF;+-2D8;
D^2QPRPTe>Q\X#f>TLBR&-7?1\/:b/@Q3AaQae>WQaf_=:#QN@,@dDEY.Z#c>Z=>
DQ>_77I]gf:YO68<fR1PKHK\^a;,P6I]9;.bY#?:4(?(@\/deI;V=3)Sg_,b??<X
c2ffB]=6gH75eg1d87Qd(U4@SO;K@bgYQTP,OJ5]edQMgVXRD0JS3R6-Z]c/dDZ.
#?4bHg1BH]NNCF0Q&.JANZ#9fO)fP7bSW08<NV7dT20eGW#^I:W^-@YQ.]D]C\5B
HcV/7+((IG3LD/a\QDNM8W&5;G3)BU=)@gc-@&8c7D<TbX<&-UEWaC4J/W?UU2Wg
3#M<5=JR&-J&L(abIB\Pg=.M\+XgL/N<Y@;+)+VZOMcL7[1#a,]TA+,],5DcQ5P;
DcMXD:94Hb37^]SHBJ3XT\DV^ff3=[;L9#GRg7Jfc1g9>I3=1g(/YWM\e_OfOCc<
Cb#>CbCb9BUXfR[NJJ\[4=X(J\d]e.,7?.X0b?<f6OXcH#.Je+S+A-c(H2X^5AB<
U+b-b25V\L+;1?/QAWJ.T0[1NQeU<T8M2J5M=2PBgX25]U/?@-A0dJ@MN[K2E9KT
+?<aB<R9SO]QJ(aa22G)=L\d-U6T\C(&W8^8e0a<aRS5bd[^J81;FD?)C7Z,7X@P
64R^E@-=9:+4a5aC+fD5cE7D</LW@+73OVFIDI=2<)\7JSWRA4ZNg=>g3>Ef2N<8
5X+BZ5[#3-[#ET)8@>#Z+7/6@RPf+X6IU<;2]^78=/2@K(VIM-,8.IX3g?.@@@a5
^&e7^QKS]RJR-d^,cR3(2+7J1/>8FG]egXX)Ed2U.[<J1,cD[Y+B+0J,9.1-5JH7
=>OH+fMCUe;eK.59>OFHJ?V,M_6+d+8DK9&XgVK<8RS\61Z]Zf-S-aO0fA&-gH4;
CG9E[d31]CS]=Nbe][15)QBc9ba>J7C#](L[NKI-?PNICK8>9RT4Ec\W1?2:O_6L
J#0/X=J9_ATgA:be&V3Z?<d8G+Z33SJE=cPGQ)WH_M93WMRH>:4AF?eGaaHJ#D(,
XFL(R6YL/OQ/98UU3>[@-_(;0MT?Hb0MJIg;QLc:H_#ID34-W[@e65YV?Y02P91^
Y_d15++Xd<].WS0A<9G;e#3C.?F6UO_fJ(A<=L8EW(QUF2f[)=fV949X<G2^[[.C
6gUE]f,4EPB6#/e[2Q<;^_Y9JC;BIH@;db2bf:.;&WU]QJ[=#NQ;4:0d:^[6NI[,
ba2Xb23KRL>^VNIQ,UP#OIHNM3-_FRcU_1fQ.6>#b<D@VN6^N^9B2D2)cA.Z&C3\
S:7F=8B602c^;EKIANTf+.1<QSM:)?e[[QS+CS/BNQJ[4MJZ)(ZW_Z50CFYF0S(2
(4^H0Z/B?-E3/P<+GN\->4K))96LBJ#]&M_-)26J5PC,QIKM0L08aXUWNWE>EUUc
-?JY.>GfL)LAK+EPDR/.^2X(Z:5X^Y_0LeXU[JP.a[=L<BW;T0bfO7AKC@AH:AXI
2_K)]R<JG\c08LY1LgFeZ&Z+AWbT6\72DP2DW/OM\//./fLF467NENS[1)X09JbH
K+PP_eO6+F;2TS@ZD(G+S;.U&E(;2QB)CFSU_Y4aJG?,=gG.3#gV&E60\Q_3J>:K
I(,<fd[+1dc2K6]Z)1+./&JB+A>G>S,a63Q2aMfH>,1@C>KW&SDCKN3C>US@(JLV
__#bYM,1UY?RIb9aF(0G:@CJ^8_2,]dXEP_&\<:S.0_ePRSbRF0:BI=VM-[bD2C,
RU0;9dZ)_48F)>MeX5e84.GZ,@A4bY=a1_e>KZ9A,]]=@V04+4d,[c_79,:KJAbG
B9@)\Wf#]M?O^0]2e=SPa6DA_/]6.JeR,ON?RP2@0b[EBF(6g++N(G@AX]He8g1Y
5JLT5^NCeQc,AU1>U:U<2SPU#LT>L#GT>6Ae[98,.ER2#[/Z#P>:=ZMUQT+TO;LT
H<6^1K>\Z@d566_-CDR70P@BE5,g667E-6aK&9N9ELC:bYZEHU#:.;f6]J=[L4/N
8<6LVcFcW/)@faXPRML(D)^FQB,@,V)Rf>E^V2F&2NC(+2RPF,C:c>V^]L;2^?(G
&N^V4_<H+8D;2Q14c@^A=(-H[:KRE(&G4MA)9\]>ebHZK>#&27DTJT=@S\279\K8
NYL3JESUT4#P=4EAf-I)ZFaGDLHG:@2f:6Fd(SB^/\&WM4MXN/69Z.+A44K]5L8e
/JR[T;2R&(UMG+8T^HGL1QGd(5PgA[b&4.7T6^bO/gT)S(6ED)NeN.#:6[2Of_ed
X[):S^3LYL56&a;A./98?N1Q(KIbE^+&LAgf,LCT&X->_>5O+4=FL&B03cD^<d@?
@:UTHcOR.&)&^cHN)7J&X[>Oe1-D6]Te)Q-:Z+8EM0EcX?AF0/;E5P43RL0g41K0
\a4WZC=D<V>@aWLY2]64#EWM@MJ,T1fX7OG/:aQ&>GNK)^C+P;K9]W(<047;A.,?
#+>THd1>L/RZ^^@QM;d?NKE9]Z^2/7-=3REU#EV\(SRHVA2KF?Cg#.YVBV[9Mccc
76fA4Ub?[:f-^N7BGDKRZ\X0c)_,.PU3)Kc?];_>^H^>5A(?(88(QQ0R.;cVfP0c
=NdL4T^f;POGTaSUG-JZb4D96?.4(-[>,<N&0a_OdN0YJMYZ<AA36dP-]55-9H7Q
6\#;F4M]3H)DMC8J>8Pc/M[JQ]KL0Wf#16MNXJC2ZXWcJ#(U#CA\C<?fHE=:<Ndc
<FQHMX:c,W\e[XR_D)2ZKKJ^c@afE8FJ_4W1:3Cb&#&/8&#N61.SV[Z1SbG=7=^:
-gX\10G:.Qa0\EEMZ4)8Z0Q6QdYg;e6JeFZ0>34VH]]3O\6Z@>g:A=XAUR71Q_T8
Z6LW@==X==-LXbPg8d_a8T,/J20aSD(ZDe?eZ88[@0;,09F+b\,DU:J).[UIXa^N
+RC8GH_X8f^F2_eFfZV2]ab7JM55R^J#Z@LOFHG7CeZGM_V9gUHV:-PT]0(Q@M)=
#\M&7PS:dE93O(@W4J8X/FJHOR06\TcMPTX^-Q5?Cag4C.GfGY5N:U440M5T;I\V
D,U#4)7P6?,?^LBD(@)d<cc1V64S0N?fH#C\IZHY<8JK7_/PIG7YNPMc2eEK][J@
;79J/JC&eA)[+A<?\JG]NN06AN7&8?BNXTHG\:X4CS--2K3#.;N#ED^8F[g)=cO<
gQ#3KK..Y@WW&W?FB9\JK.G&RPM7H:_/fa?aS?bGaES/V;b040C.F>^B-R\?:T@3
AR]F6eK=RIXW55>E<[X@(G#\B\)KdX_;fJ/B5;2_;BX#R1Z^J5[GLIPEL4d,(R11
74OZ_^55b>0RN-cJTO-g<@ZJfBXR2LaeR=J#,UfQd9NHH+^[+eXTEXeLHTH?/Le3
<S]P6=?BW5FD],3c@<8MBK?5RB/GI0/1DRZL=4,;)M>+U1ELgPCQQNVR>T-(X.b-
SbMZ@5NNe+.?.P4=EYf3#3FcROb9W:.--=[7@R#SZg3UGACUN[bdR51DQMAP3,(+
F1C1G6AN]K\K18]=5TY[M]KN32]@f[V(P?5ABQ4MB1L;BT0F;E,NLU#UK4^?bJD-
)[bXCX(AJZ;SUDR/W0DA.5adUgS/WZ2a@Kb2\_C/ff7Y1F5,;6473BE;EP?PegX9
dGU^YEc^-.7R.,]8LW7U43HC\TV8<C7DB:4B1R:#&[_UI;WS5DBIQV1-[MYKF2+Z
L<1M@ININ/\].bCb[bAg@]1;K,;E3f/4WSH)O2aJFR8f5XS6aA(IG,V:&:ffe[CX
/,7X\0W/d=R6F-RX_cg1FOKe8I9GXZ7A-eZ/-)Y;dd\cQ6[DHGIgg(NFZ<4fOcTE
1gETIKOgBe3X3:D0Y6:_Q;HJIH)?9B:O]6b_R,dBL)BG-]4,1<T1C616TG2NPeZ7
6XM\UKW@D&FJ-QX;A,5H?YD)[T,6LeL16?VK9U+XS9NP6^O=.&8.A+]8]&T/93(^
B#X6?1BNWI3.MTEXJ3Ng+f6CT]##?MU[78A[VN(Y=eD&:3K4(VLP6I=5OXG1gO0N
MVL6TQ(5_C6QK&:B@/)L=5Tg5Y[COAS^KTL6a;)gZWTSU0bIM:VV;M^:.(M4XW<X
N^1KL<DQUOC#-N1G)P6a17OH8H5LYX]<OaQ,]c^S)caHAL=3++H1[9L4)7-2V(?J
?XbbXJ6GT0E;4PMX.\HQ+fYJaO=ddFG;,8CPK/.FGD^@GCK0J@)R<&1XLO+X>1+9
/+T+4fDU68JZ5aA_IDF[@67N77bfLVF2,\O+#:cECfY)5CXP)Hb?-G@+YE+T=@C1
LdDD03(K.G9?+P[NCd0Q>5UW58QYFNB&FKG[IL_,Mg#8&GZTNVcB:,a=C;5@c2,P
</GM)L]AY6[J>dG>/HPA<6fQGD<.4/-#PIRQY<9gHJ2SQ/_(6QaCA68L]+0Je;AF
BaR)GNW6X,._/I6ONF:22c]Ga#I51eb47)e@.@:QRM^/?44S]>IA9<fcAa^67V3S
2UVTNe>Z)f,5.X7/ID/gTdfZ0(d_)4^\R(eg.=&bg7g[TU_Ib=CcL1UGK>3BcNQJ
;@06:3@d&Q8M^;eVMRXWd4K-P.fLN2df@AMSG5N0]B^1R8:BX+=[#@ee[@Q,I<UW
75d.P9<&_Q&>Q)@e?>RV/c,QN\WYc5],La#((\#Kea[M]DT_N]HaC3^1-1gN:dG1
)@>2-U1<g/_Y+gOE<A@[gM:ZNcOdXOU_+VN:&eVE8H^HfK-RC9^Y6#:?M+U.PNEg
T/.FVGF,D(gbK#H)5bO\:+G:N1_U=[+V:X>>g?D:;Y0)Z3O65=X8P7^S7,M-_8U[
[?(3L4@CYQ1GTMC)#C\Vf1_D(aOS-(RXWF<4^D<LHVI,(9A-&_?/Eb/TAbW\V<XI
F.P(:g,;OLUS=98_<?XH#,3OWYW3c#HW@]^0gUDDb7WQJPAbVXL@+aQ[T[?(f-#K
:T6],[U_),MZN1L5Y6X=J9?G</aH3TZJ\Ze8Q7/@P=#2?R;fYGO[J[OV(A)XA0;G
<_:/Y2^><5H+bQQ4HO&VPJQe/YP8c#+Le/7aA(ffOYD@GMY3SD0J/QFWQ#2ZY8Z:
F&T7BC2XCSX;K]@/E-BGfPg=NT2_X0YNG8@ST(_gJ;.Z6+2C=E20R<g(dYaI?Z+f
d,eQ6AN)#0A@[)]Z:IYN6>49>G+^GHO_E?g_J)5@A>7EGB;3LTVG_,:Wa,@XXLf+
X)#X58VB8<R_c4bY9FO6G+_,[\gSd[IE]4P:K(NL+@OS02c#<<@5b9[Ua&d3^9Oa
[RV&fI(c(?f1&fMW@T--N=?+&?O;@S]e&X4VB=NC>c6-U3<D-TM]O7)P]-M@_3NR
E/\TGGFb/T_60G+\GAeG6R)2cV:JfSMM4M-)ITY&cOU.g](<GIFeENI^)PR.c_LN
D:GN[E(^dGMfG&A5/>CHE>1MOQ=[R@>#4]W(B4>JJ:_a@FO&a8[JJS;FNEUHT^HX
#_6V;f]]a?XUH@)@,,<cXB5>/X_c/47.:@Q+8:=JRM,@8A<],9CDS[J,GCLd=A>;
?V8+)]<W#=eX:+TC,c1#/7e:5<+GEbUGK8HI-=&/OF8#Id8Z>^C\:XE8^4#WZM=0
3b3ca2\IA_]E8fBVZ+M4HN?cg5:/H.2F?E-AG[B453?Y<YM>X]e/baI?52-CA:eR
;?c9Dd\/+MgOcF&b+NMNGYQ@g;@bfac]:&a_M9+g02g/cZC-dWBBFIGBXJ55(Q^a
e]Q4H_)]I([S/H1PE=PV_Q:3W\W@--YTZ8cN^@f<;78?4A-TM\SK:PJW12&29d3A
(==G&B&c8VW5_CPLUcUKTb^]GdMZ@VbOWM^I7cFT]7S?^=Hd(8P+0b[TNAe96XV-
YQR2YVU+IS6H_-MQ^UUb[VcEM\1(\Ia<N3P#?I/?Y1C3Fd8[]0Z5XgS9_#14I<]Z
XE3E2&GM&5B<&c((:KM^d/I;FgSVGD5aQH[C\GHX:_IMK-T:,aEWQ4239CD,J[,[
BDLC?5@1?&^T24fN<G+=3:3@P8_)/S),ggYBKC?@W(+AYM0Q_-K@GU<>UE)=Z[Y&
a]aLT<W+>5WTHLVRW-I4RTXfDIT]OKLV/5N=T+DX6Q]?3B,e]=<[;4WNN#/Z;MS8
UZ,NQ)LOa,.;BVBS/DfSE1=4SYLbU,:[&B4\QPZ5Df&A9QJQ(D.2+8SZ_&VJL.AT
7@X./aO>73YRaEg/Bg<PQH=gKe9F(R<^YL,0SZ[V.6IZ11^=7<BZ4?7^YbNccJ<W
>b[RU59d\#e1dG;G6MZg#QF5[e(Q]0=\^C/L+Z&]FfebE#6IbR<VN1:cQ4OT6bU[
VeXX7.G]fC7aUHUX.B35cZ;J>HeC-[BR7Df=7T\>OU+H[YYc2f4I+36BZ;)GMM#3
7B+fK<U^/bZTS>@LN1]5_=7YT:J@.::W,K[84C_11C+S/a<2L2:[f?A>eI#eEgE:
:90eJL,MeZaZcOPBPI2<aJET.b8^,[:AO[.WYV3C0Q2d+)_fB5/:e8eJ_,A/WK(3
F9_S21OP)[dJM\(dT0WE=LUV^6^0?(5FO4eAc^IJ79DYEcfQ9HW8f]OWX^dZ:0HM
83C\<4Y)>Z+UIZN>-W:9(&g^L[Og8/5G:d7R2+>O@:/<+cQgcV,:a([L#CI+f<EM
W)9@UXg=WCR)+H8^T?#&:FVK,e>@JfSL9eI];H05Pd=#]U5F<+/P)L?a#6_M^=Pc
>Rb+/P5K.;9<3<T[8\L:Ed5?8UIS,0d;Y/GU(^VcgTWNL<)1D)D#<T@R:,9)IDZY
(_H8[M6\;,WO8[5S,QOR,+E1J1^4/L.2>?.PTAV/<\.fD8;Q-Z#L3a,Y(PDRFc26
(?&H1/<)DNb7a4cN&?a18#ZDe<KS2<TCOGKEUA9,.LHc7-R++OCB\(+G4dE7PK5A
?fF3T?Y(8eU41>HOMZMRCX+\M-?Y=Y><U(QeHG_gD5K2&_HFac4#YRAf]TW+S&M]
<F.gN/dVU_ONC7]2CfBN?XLTW,U1LYWQU?d@38VW^8?W&Q7(I:R7d8C]AIWbdVL3
bL7V\NF,B9N;R^9TKGgD2,A7)MD6)f((MMe7ATT(/5NAB>JIK;\bbY[3KQUSVF^U
GIS&Y>g8?Cdf:XIIN?V3#_GUJ5c-M2Z/2:I]a(b6WFV],04Y>V6QJ_76(LVC[#@6
Xb8K7\6T5)C;==.,-DQL@EAJWEPVIaC@;D6Qc&+LY\F0B9X4RC?F3Cb8W0LP64?E
NQ,QL1R4WFD8=+XS:#Q;Y1;D0c/+O_gT#,-+IFd2FL.9IOBY2SR&@,:_I;ZDJcHZ
e:;Ne.ZQ11>&I?4#?cJO>R-b2f&3Z3gFB2);56&<f,_37T;g>W60c;@g)Le+_&a;
(_P+[P89,LC,d[^#c4<AFe6B2Q:c86E5A4:=^A:98S,A7PKdHY968>C7@]Ub).@?
.C:U1,H/-57-JQ(DOd-,/5:\),BY+Q0a^+6WBW+>VdMbZ#/RXPJ]ZE+c_f3RG\X<
2MP#3SCV[PW^K.4g9)T#W]5>:@L\gHM.f+C):\RP9E#G;e>;@d_]4XV8NN^OKI3W
D-HLKQBHNYYIgXEDOa#SMg^S9ebM+GW:7#JYF].e,?BbfRG(&14/Y:S-E,_M]>JF
L5C<P)#?ARdMW0A[,OD_X7L;WX,-B;S>PCE=:&AXDM\42P=K;P>CIW;L313PGY)>
HY<,Pa_0I5A:^(Y#A6T+E//0Pc)=eV5WLb&4@2,P#GYWE14R/Z?\65ZA+d?+MF&c
QM&QLgN+QaIV?[M8K7PB=8(1RJE\G;ZS4EH1Z(SC5Z^4U\Cd&<3+d7/RW,dJ#J=_
QD8;(U7.H>H2QIE,_JJc1bBOQY4)=ZX0.XG>Wgd<O#=HVLU0NNM6RC+V)(Z=c)cW
QQUO8EcM@&I-O\KBINdWVP3b)HY+4aF-KcZeF^a.YZ3H9:D&#aaTY>))?>=O#9Z,
b/:#QX>PO(^(X2^df3^JP(B,M54L_CRWg21bTd&=T.B\8e515^<-/R09SFSIf7K1
,/&b;XaOT?LEJ1DWFeTBaddf/9e&RH09D8O\9fCagS0bT;C=<?<e\5fEe+-MMA/U
5d3#WD+:-)H6NaDg3AU:;1@+T7BM[C_W1(\R;5E_2>;+HX2BX9eP:&:W>2,g2B[0
[?R<KE76CS66d??Rba?7MM#5<Ec)02WbX-&^-@UP/G8DC5H]2)>1Rg0D[[I(AIAa
1Aa(+U?]7<fJ,2&J/YSR@YLR:;#(AZ6Y_A47T#R8D\W.OHO;L33B/KfVb7Qf,G@(
;&Y2B\9J#2,,54)4]a/7:2/^T0/57DH)XV1^]d^U9[=d:&cPdCZ=_eOJ^(&IeC>J
>I]^?#HRe^JOgY&5E_dB#-2GIdCW(@/1QW&2Gc.fFV,JEE.^N-[VOQMe^.f,+cJX
KT3&B[\H4@YfV6cGbb1SH=C_B^Ta3AB_(?VO&)D.Ob&:g0HgBO=>a#(#,73A<ZdU
g-QbDH-aV<\@,(UYdb0cZ\?&TRBcgZ=+^C+\e?1IN3&\<fGOPD)Sb1STR8E[;/J;
=TJ(G&.bZW<=Mb)B<,T+0e/gL0\J+XXTNSXU;TB[\U63fM7?-L2e?UEHJ?+WaSR,
CIOKU1[=e/D^H7;f[>[BXbUP1\-4+HW31XK#ASQV^S-.^K(d(MdbdRDZ&;F_Wf=.
K?Q=)M?/;N#]98]9a3_G-;K2#d9C)cDV=XT.\.7()6eW2E1-eMXS;=dRLgQX3M@;
RN5XD?77[.S>;[UaLV2-6g0D:9VcC(f-eG3ZW0JC+T<G@1NIOb^>FUKXRR(##H\2
P546dT6QBC)UD^g<NLa2?,PGEB&FPG2+(ML\7S/;0CEBd4g05?ce)d2H-14dY7S&
)\U=2><H-b.[FR)?KMHQXZ\B^I:1UE+Wf]G-RD^::G0/g\Gg1]1[-V;&c^0YLHdX
Ac<JcF/S91&KFYU)&Y7@&40?6DWT)/4L3;5FCdP[?<#VSP:f:U,:&]J=7#(?+9(&
bASWZ1d8-c>FcYVN??_IJNf0b+D<C+@G6e(Q78,-JVIN,JE>+)VR<[H\3TLEY0,N
Y]438)6<FZ0cE.]/V[Z:e5_9(aTE;Ke&6P3gW=RZ@3bbB7&fL;c6-#dA7KB^E2aT
++e81a80@H;/6<D>bLg,HFKUM3MAW,9e2_##34(-_d_71M;#gPH;ROFFN#I/dMAg
_\3@4-SOI377TT##5PLY>dCQBcefD,SIDFd<^fEH>NB/@Rf-)7[Y5L,C2OJ2&=Z4
CHO4(bQ>Xbc2YS>M0X9Vcd^G:<T)?e=)A9?:<bNO#\TC.F<&;f07W]SN].=CW2E^
bDdR<E),[[E5U^N&Z&SbCWTadbTFB,X-(->]H4CgWc,X#U.S:8VGdcJ^]JIT&4QD
)adMf)MT<K^dM(_S5),7K8T)2Ec?X@S/a#3#NZ,eI\;>8a+ObLR><64dFcOD3&8/
QXaG4E]dG3M_EX4<XZgFc13IC8,A9eb7UY)82-_4&2AHO-RM@:7LW@dSGZ/J@f2[
V^5,[V<9f]^Y=<JP)X&QN<b7<FT>-7NS4W.E<>J3agG@OF37d7LR@f6YeW?]g:e1
M13UU=>6UO82Q5ZYO1&Y0^RT?I-8TQEEgP,XWb(\G/-J>47XD<^c1_[7W&N058gd
Ja.M,7Zbg)1HLUU@NWNYeR_CN<7fV+X[>LW(dU#,2bYbPeQ5:c6)e+5gA#cf#?CL
AQWUMQ9NTDN-@7E=9)ddce_)aCV.FabE5?9Y\32MKca]a<(GbA@]M>DG#2f]=_EK
]a3GX\<CPJd+^V3PD>>UJQ-W5WYT;)0,,374NTX3L=TL4IH_8C6HX_K1)4dX@3&c
.6X2US9.V]_<>c>0A:H9g?QF(JaT92df)3#d/@\BO+9Ng1BJTPHf2V8_DC3g3F\N
TK6W;838fBZ<gM,XHd;V.7R2JWR,J6PP4[D4CQ7=L[9FgGU5M4\/L[P[,8K^LX1V
K+HF.N/DJ&DN<<8\d]Z(fKa,8(K)C<TV&@2fBaVBeOJ)L>([OG]S_8-^+_.G@&DQ
5JL,/0#&bKWK]\9.90?2^ZVBVd7E<6IbY+=>M>aFg7+C&a_?\&KBOYOGZ+@[>[1T
4UH[LTHUa=D:YC>SHIIQBb_02Q<C_@+WV0(a^b:-#)FM22dVE&&JVE?/2VKeMV.2
E431O>^IJ\<Z0@/gdCaLd/:AfEa#.K0Jbb=e=>S:4)LK3]\K3C<YK3HdcY7GeId^
UYX)[5+A(1\B,8?LG3EN4@O<YVgTYM=N/b:NKAb))+9_,EGL(S(T:]B0;.Z8[+09
b:P?31B89VQ/WP&.)-1<Mg@ZDa=f^SZCI#_NT+DE]R(ZEE6BW/XO,=C=&J<01N)U
LIagK2YQV&8^M_fF&I6Rd92J7<D:#-U@egCC4QeKOH84H?S1L&bB2@.CM_1-^bU@
Z&]<XIG1N<P4OcE[2QWfRJ/0UL@9=K8/Q^S1PJOcC^>ZH:E;1T.BF>.EdSJaBfB7
@UDT#MMO\H[Lf_SBQ8]&>.F7ZGaQ9Nc6f8+H?&@Q-BYBE-XV\QB<X2T]R&7#@;J+
+d2B(Dg+(&Q_cMAc#+BM@)TO9b8+[,aL4ID6ZUP+bJ?41ZR\U:DDN:_8P=FZ66MW
AY[@I4_KXB>H)[3.DdJIbad58^Kg#DS]9G;/QM./,<>c?e@S90VC+83e+UUWI0(E
aMcL.]MK/N:(@)fcfD^Zf1\M488A1eYC2SXSa1T3a7Q-c^-6O^+)fH[Y#0;+)U7+
=-2f2):+6SF6UV0KdaKX.aEY]L#ES>KADYDf22J0&FX0.KF\a.NM_U0N&c@:b<NX
AXcK_HUGH<cOFHHg9eJe6cX1UXX_bO4F6Y:V(??#G2+IV0eW&.AM))5VY&cQM/T2
OHWCUVU#CSB_;908>fIU8)M9JFFX3=N[XdQ7;X4&LRS@1Q>9B<E+[;]_IG85@5^A
/&-f#gALgP_[^LcaB5Mc57gI@][DA#<beP^VX3_Y1OI/RA3XZ&TDS(C:&a37OX\c
2?/?7(HI0N0b/\W3>I.Q.0P0G@PAPB/f1CgL8O?&>M(1U&W.f38]<H]U?0V(GI;G
N-8/@_&R5Jg/H.DR]B2/R++#OJ)LdC[QMdc3B46JG3VP9D,JLODM6cWW7X9Z4O9O
aVI8@S=6.TN\8+N)(:>J(Ab4)B8>@G[(GW\D#[Xg)Ab,-YPMOV<ZWV]Q9LH_5^_6
VWF2XYDUO7UFA@\3(:?P,6>O5b-EXX,\KC@cUG,L]UW^[CB;.2<b7/_@9NDF>6=:
WB8bP<Y[O2@>X(U;7,g#Q(Yf5(WQJdOXX64[\9W1f&V?Q2Fcf<.0,YJ:J@BQ-E1(
RJd&(#/D,,>9DfF4GO/H=\1:#@]4DXSD8W9#Y_B)<R713.\]2;d\JEI#g&f2)ZC)
cEVa(8CDH_d(7XJ<+cfQObOYL#gE7bPU#,\?_O6Qd>,98B0?1C9H:IO#-YIWK5]P
R[^>BBX9[KI=36e3J8G3^W;SH[\0^7>0^N;WJ:3+eVUcbRPMIa_X5]R2GD<P5[d?
IAb-fY#/9C=O(cS)2g5LT)@gM_ZS1C&UA2Jfg=QJ-@aHF]D9ee4?&#79bXPWe.,9
bRORJ:07RE96.IAcMQ4QE([)O1&O#5JZ&2-DXP@/(F/\dLI\O1M;<V5d\(L?)g9@
?38S-E(-C#HY;U],7,;BS),4fI;bO#D(IOb.Ee^A9LH_7>,L7_0#QGNANF54fW&=
?FKgWM-+KJX[Zf=5YEc.Lc^DYb70\2RV\@]Pc2S.\=EY?5:5&29\6D\FVWN=Hb<.
7W:aJ<#WGMPd><8CcAfG0)I&,\K.NB,<X^/T\O(FH.8RNNQ/J-#V<3YW[<E^8/PK
0K3MDb;78Ce0bKRJ2Mc?ZQb5QVG8+)9YV<c#LfKNY;dM:1B///bb@@/>TVTZ=[6)
&GEa&Q=M]@aF)c1;O;a</F&>DJ<&d3M+/+,JLQV?)A]2?-Q4JcVT6aWXb>M?@>ON
^?0OC2H.dP)8^49-S@OAU;@c)eSXcBFcS;XObFR0;&?<R/;MD_X9da,fg8PCPB)d
3c(f-F2b(S)dPJ4Y4@EI_=B^A19A8+E?>XNF3Z0>cJb4ON5O+O-#2@c_(Fa>X\@<
,PQFdcfS09A_GNf+UFTO7)NMQB+A1aU:-],_,FI^H:@)VYXVgcd3b9O(GA-]S1.J
YAYID&[7H;H?8IH;=_TR3(:?##V?]a8&g8F4Fc[dIg)NeP5X1dDX4fGT+64+&A=(
Q8_+D5L(Y6_YD_/-K][U=CW#L(4BT(,C-MA0W@?:Eb]fO0..>VWKYe]H(5e,1IEd
,YD05((c\M]>[WK9>6\RO]\7&,EA+9N)>#V5J4M4ZKW0X0eDR#d/712,S928:?U=
g)4ffW#4AB&M_@YKC2>5D+>PHSIP?>@LJdYK+WJ>f>&B9g<\Y:)ZV-AJ]X>3CEQd
;FXeA0H[5cZCM-IE^ZV@[-?7R8K2[/?a1#4W.]BU#Q69WGb;9_(d,?^+NQI6<+0.
>]1Af3G?UGU>\0_[a,c?C?UXA/F,H0#MNVD9VbIM:Nc[(;ZNH:cHO43:95PId6.:
E21Ac+ZP?;?JA#398M5F^&e.(ZRI70PYVGQc/F>;,5>=BWC<S[(\.MfOQT_bCd3L
^E&0=Z[dLK&VT>M#FcK>eQ=S(MZX+Hggd@^Z^I&3J8((U/>E(Z,f+eUD-eTJeC9[
<2:YJT+\/HZ3Z4,TX/[d1/])ZP[\+NPa2]Hb\M0Vd&PZO>BQUP\WeW67aAg:c?LS
:7;,a)MfCd^W>I46?I2^MG1(0,^4+\(+N:e9_S?b-@EeE5-744@VQXFML\N73CX9
c&4=;<9YfOL]\@]_Lg:>PJ+d2g]ZJM:1.(_DLR.,6J0/U?BF+4EG?U)91XTI([4g
Y&>:6N(-=:)T41X:(aU7&@6A+7DJ=JZ5V-.3-B/7O#M(_KS8I=_-I5([7ERN+<DF
=2=Q,g,DK&6TQTGBcJ5C]^70N8gWAP=)Kg(I2Zg\eYgVWDSER:Y@<]KB0Tbc([[G
PI&)36eTSWYH<31<3f2HE6(U45M3GQ?]A8<_1C#^c9fb2Z6P[g;U,BB4L6H_BD#7
0ae)2Df,0YHH<Y-#2#TCQ7>T6&/QWb2\/3f-V2B39dO)Z-0b-23eeATP+->[[O+:
@(B7Q8+_>b=X.\^b2R;(2(]0=DS,DH)].)aTOB(5GH[[#HZR8@\],MP;a1M(?]D=
9XXS-I;D3#VUNWFaT7_?<R/CBMedB0U@>K+=)GDZQ^dD.CQ80:HVN(V[G.UQBTC.
X)#@O)?O+#TaPBd6A5:e7+QAfA5e^JdB)L7JZM),59Ndc]_OH];95(LTD2]NHWR,
<C<XE3f+K>?b27G8_V4_]bfW[g4W3A6?gZNA7^M6^ULB=e-fY1_QXR-><;W<.YQ.
0;K-L,c<:TdV2Sd96KRN8CB)T5Z@F^H,AS]H]_1A27a8gH.6N;YdU0-b91HZK7Hf
KP=fSNAa@^Sd5HcB5:AOQC=.\f.:<J:LTYMTG+OE=&89#b.=0NHIS:Me8)/U:,[2
R:=AWPDLcK7KT9PF>19.Z0]1N]]2]_?PB/18Q+SE2,T4;KTf,+C64VG-OH2B8g20
CG(:acQX3L<D;)=CAGX8\VJAOFZb@W^RLRUP/)UcCSdQ[^SN&:5a./Fd19S/T5_P
gL/5KIc63@e=4UNXWaR@@[@3Rc_Q8H,&ZB>E&8T#bHC\UN=(g;?Z1Te0:Z)\H/].
Bb0Y0VW8-:2-KcH.(PMU:-3,&:<6()6dUEQ5a/CfM+Zgc->(EFe65<.AT^UUX7:(
;R(8b8>+W//Z]4I<4DQ2BV4#e)>3e0e#HOE)GFG)SVR(&=:3<c29;8EB9XAC>V0S
[MSAT85@,gCS9EGKPJ);KaTG=MaT/4AfOGKE[-;C/4G:G=7QUaBg]?^39WO.a/.S
)MNOaJJTAgI8.g&4&C+\7e_[-\ZR8UOc?X21O5a5VR<QW)TWD5J7H6,TRFPJ)Jcc
8CEEIJb=g5#I);a-fJFW0I[-ZIX\6Dcf@K?7eXIIgQ\D>3#Q4LM+f5H,2cA6]\FB
JD.CW-aD#@RDCIQ_#,M4f_.(56S+b-OfF4;IA<0+85F+(A&8:XReNFTJ@8\W.^ZW
cCK&SBb&H/-@JM&UQM1XC-<gNJP[+;FJK[Ee75;?@[YaPTXfgAfTCb2[:.FbB,9=
M&H6I28C3g;b_+Q5AEQCMd>K.4af6;_5)R1JXW7[U;]gLW4_UEC4UfO>LQ.V/#dI
#b=B+CLGN\@0FAO\.Me3#/5^Ic?57Bb.(3D\Z+<^BO]J030WPBJ)&1a(&dIC&[2J
ENge>(,FgAAJ_d03.ZBdA65Q-(LB@DV>BGeKV=FNLgXL0&DN6eF.VC?5AUYEV,J3
?b?[F(Dg1#^N=GE>3PBU<Jcb/G56&D7B:U7WH<R2Y1A^?QBX<7MOE.<H?2)Pb8[.
DC7@AA3aUW>8PRX0.IJPI?0C4.bGY/57U@[O\WG81g8>V6Cc;=?=]\>N.X1S1_K4
NXb7L)(QLg0a2T0dH17OD81[ZMN1Z#8g.^IIJ;a.\U-<;\K^;&SNMK^e#SJ8TV@+
S[+f+(P@>?E:<C06gGUKECMLa=3P/3L7\H-7;W2O1DW(C@A+;c==7H:>].@aW4O4
X3<ecc>gOU[:]a,=8-P9(,MCAgFV/:_Z93FB7CD<\bL&V_WA7HW1P9]b49HHC#(;
e_J>4[cEJ^#CFe=D5O13B?-7;MF^9U.YBBR4&#Ggd@)H_(88Y&.>/XOAa@P\B^G:
;(S-W=[WaLU](D&DZ85-<?RU8[U2cTgA,.3>9>C<?,g[4Ic6a\YF.U;8-#d=A=N4
5&B@9a-1IcRHgdYf1Z=S?53#O^F+)72LVF>WAa:^H.YKUD[4/]6-](Q7+L?RL9B-
[TCV/H&L9RaY>U[[N&/&CW>Q_B4]0V2e[)M3b9dCOTNeQY3,NX@U9^^V)6B](AEX
Y\?RQ0HcgS.3W3.&>QDP_C3EQUK8H5A7BfY+-\fVd=Cc7fL+^_6]1?bSI#O3](=b
_R0]GHOJ)K7]&7K1WE(C3+UOVfW+?CF<GYABL)DMITV]b,?f+U7]D.@cPK/-YMcb
S3S,A<Y\MQJb78]6M>daA(P5WRD6bBLA:K;4Z9E(;D=6SR0]WfIdG<T48Y(]6b(1
g#&@+],Xc8DQ,^=a+#Og5:;eg53KL[M@UUbQVDZ;F6HgG4=)NM<O])ZMf(>aC-K3
dg\1#FAX4,+KD.=DV(5(HN7_=c3Z?:=Q9]R]YaB.C6Z#Y=<71@,64_E8Z<R)B&G:
(_AfO)Z,cG<^c6>&S3G9^6(+@#D2GTGJ7ZOW9Q[^T?UI;,;)2-7M@C?5YJTT;;AD
<a28<cTQ&D-:9[//G@)42/&FaF6\4d]GB]C9=7]#4(bH:F(4R;6=(-.KW<F<0VGU
YgG9Q[B8@(P[ZU3Q_)ETSBPBO-3Z]>SR#GE5Y09?JN6X@b[QZV55>OY:P^cdaaY:
Q/+[JBO2<<FD(cK5F9);)<^O)&BaDMWEFH1=@1^P<=V9VX,?_EVUESc=V]+IBL@V
UaP^[90E(F/(L>W3AF2M2HYSWXCXK1J[P4MS5L^:&B@Nb-;>6d,G&?5LL>;=/K.=
b/)8^)AHI3g0+5+E@]T>Ye04,b/PX>.;J^MOCN:XIe)#d4D_-5^JT-8[\5#AedeJ
CBNaR_7a/N[faF\G.HHZ-E@+?)(6=CQKcV]2<dR;g50;TUX_MJ;B:\RVGU]#c;S,
FJ@(G6-\;;_XdZ?G\K3UI6L)6RA/b/,+6]>\\WGIP@T9H0F5-ZU\P04W@>b(gS0D
QeIK+:^MUA+5&(1>=bH/UP-V>?3FS&-dTOV,-fIAbR,/(-Lg6/<#c1XSgHGJc;80
[\@d2JdRPN?2;>gQXDEcE?5Q0c_>.^e_B1L)R1Z_KKAV5&K#-]VbEJ@O,273[+??
YXE:\/LF^S@..JT@:EfEB;gL5b0ZJIB<H\S[^@+S2>7=f#.)39cFI,RMD<L#T]/7
gAEJ./5OYcKLT#O=.NbYSZ;W)(=&IWG9QM75aab=T&]e-1WD<XYG\AS6-d3a<,?f
&cc>/)c9DG->A=g#]O/+S2CNd85,#+DdWIH1\1EP49U#a^?:LM(bTd3>(5[8P;PE
FZ1_1a;CITZ22[.)OMK:5=2MYTK[UNJTJ<1EK=T(LLB]G]&JeD-D,2NPE,8J&P1.
A4(3[WbcVYcQXYMA.#)N4f+aBU]8&2FE\.A-J@a6[5RX6#(K@Qb6=.JXXVHK5))?
JO2]OL?<fWaV@25a:eW(ZN+aFf(;V^NaF3)A9c.F_G1QCcDZ>8MRBEFZ;G182\bG
?KaOZe:67RD&/T^<Q>1Bg9;/?CYJdUD_O=&3LXRYcT?cP;2ZIB-9O<fAM5/@?GJb
S&+Tf#_0M+g2K_139Z/,-<^B(UTe9FG5.M7c-&Ec(.-9SN?b+V1[U6D.&P)<6Y[L
L-A?9^^5Le.3+119a,N/aRa(IBXbZP0R.1<ZA0c)VBca[[];YE0H?D.E_JXP^4)M
CMWN1+\(7#JVE5ebN,2&b0:(TCPeJ9G#M?>@/N@(N/9.[XO#]:;Qef=SV3;XV+LK
U>Q\Q#3f6/#ZWDR?V4R(P\W-4.b4RaAW\g&(aK.1I#HeJA;#ZB-YOJA:E-V@NbX]
=+#6]d0<a7O>X+X;d#K0<7M^Re?H:K(G)aWLBWMEA_[(_b,N(T@)KOa@^)K1RC\Z
/B7OLPO20M=:=M)G:Y:L-Bb9(/M;e(a_fBRF6)f<8Pb,7N8(QVK.79^64W1\41&D
76?Rf&FYTU&OYAcGAP>M62L7M?N0DbKBL3fP?aK9-[WFY=JCJ=W\[QB6S+9OXS>J
cd<LFGa29IgMS#G1ePO#>DgS]\Z))96MUW=OT6CKC1L)Hbc209aKJa8IT06#_FM#
VZT\3UU(KU:Tgg9TaABVX6O/T,>URfeA(#HA?9c6HS.8Da16TUf3PB>V.S:G:6ZZ
EIP9O[Z)1&B.c7.+Q>_TN8ETR+;;&R1]Q/bT-NZ(AI#4B<P;Ne_3/E?QAR0<8^E1
K15/>0fWc@gH^.&@\d(^dRg^AC,UN^N.;YLI:2\MV)BJ@:D&d1gDf_#7UT.#9JS)
75KSLBO3Da0;4OO+BaFN:Q+KeJTDR7U0M+<__N80<dV_I)I3[12>^N=@G&)e7dPA
N545b.C0d=H<R\^(c6dBdfc.=We?<1Vd+7.B-,8cOG0O&59@M+;>B]8IE(PY8OG[
4GA+D[YCD_?2e>S-,b_4^_4,3QY-IBE@,D(/;F0:GT?+)\C<P+W.03dN.4/L6C/U
GM>EAWMf,EB?SCg4ed/T0deW)6O>^dMA/-IfPOYDU[SS(12B7Rad7fG(d2E;e&FQ
25[gZ@IQYMP,N9G=@?JQG=?LBY(W,++e\NZCX3+J/O&NDA7,9bS_P]d@bBcOeZ(N
D0#d&.M]gWP_^/6+O1V1K[c/6[A(EX257.<N7fe96cD[J6WF\R=VZ=;>RQFNCRZF
N9NdEWPfADC\=S+OU/Y7-2WQ;=GWg71CWccX<X/g^5&Y[.Ld5d:N/_C8N+P6L1+D
DQSR);Z)9[Z8eg8M\PaI29/[[=1gDEJ]Pe/CGG&/3a9;d?UD8=Sc#LFY\)VSW0X[
_f:8?SCdaD[IbQ&N;/5ZSQP;XW4@T@Y:#]aIR4STa2NQSI\9Z_2_H]25-,P:+]#3
4]4BW(f[?e(@<V1BG<VW6T?)9>UF\5J@Z\adYZ[VBdA@9YNBdDg=ZO(Y>gCK3AVO
L6?GI+9@,fK6S(/+d.\a].gIK)eW9,L>+B:2B^6#GYN6ZC,W/&d1,DY6[)J3<&0#
6Q6+FDaR^XgLO8/TT16ae-[B[Sd0Y\/d2_&EF3[,R+bX,4g-&5(GGC9b=Z:AW\+X
T9-fGKO:Z(EF.LKV>Vfgg[Hb?&8]b.OgR5/9_??)#P<bF@K2,cND:QR];LC-PI9R
I\_MZb#a/WNL@O_>:T];8]F[./T9;#Q1bY[HEbEK^KJ&(Pc5>C;E3YMa#_Z4X9g&
;OO0P_/??AXZ[:4\P7e[JC6__c0bDf@3BO1#Wa6[QLfeaA0ZHFg0BH0gEM>K;)G,
K,(bU9D/3ORGML#&U--J:0\c-,c0#3[.</8\e[_@81eMMdDR&L/[(K>;PeVVQePZ
NfA,E<8/e==S3bb6^He1c@[d:gGdF+I^I8]@W;HJ,aD=5g2Y_B=GR@,UH;FOTFB:
.aCEeD>1;,/6\gPdMFOTCe>9b7S83]Me_&)fB)eQ.WO+&e/T,4(eG#4)<IU\HQfb
f)0RP.AgN3O&ecW<gJ8f)1;8=e(/]CZK483<7cWW)7WI>&f6X]A/3(R@b>&fB)_?
TPD7XeEYZ=P-6^eSeC3F+T:SbG,b[BC/)&[/9H><NF>E/PbI>JB7N</<F<[EbR2a
dZ]HA2c\I(VOOAT.gcCUMDW]BA0._Jdc6K>:+GR,[RA2<b5N3WREE\ae23&TKd;7
^K.4IFTJT3IAR(H6-GJ?4d9NK.K9bLU&1J][ba>,;@LW\7]B?)\N][49@fO16cBI
PPFF+Z\e<.VOCTe3Q\)WVfCK6K4G+(d<+<DQ9]TbZV_;c]efeg(@=FM&>N?-CedM
L;?F_C_3d4>fR(CV)\2RVT;;\F?0T59?^&OP/[JEU]8P:4)=BW9dX+/M+..ae)JJ
X+[#.,2@Rc32>MBFD]3c6fbc@^DF-9HGB,45&F[&MQV_HeWETUAB@7)Og=P<SWQ7
Ve[_>SOQ(I&\_Q&MQ#;>e:?YCabe=O_BWV14E6YEG+LKdDD;8g#+De3;]b9:S3G]
_b88L_1P6gYVb/FD+P9[M>(7CJ)#W9\:d3\a<Ud#]SIM90FfWG3Ha,0@9=5e3)[;
ffXE9=dDAR:-68IdC2GNL<3<L1b]?0I9U_2?#Q=RRC+<e[bZ=W;<34IS;07cQd_Y
9<g;(E)V)9_K_c\1cRO^T&YAS5PJ4J<7+1f?CI5cU<g&T81F/@&QN,U)5:^90gYC
\7ED]Z;.<T[BN.[e:,>LSM6XPT:2)EC:]QcQ)4;QbP4Ge\E#L<A33><T?GP6<AQb
6_^MF&Re+/8C4H5+bU/?KTJA#FMff3,XC0+eMdU\1UFQ4X(F?DZ=7^^8I85T7ad=
@6C.JYA/_&FYA?\J9d9>9IYIL^6JUFaa+#>N>\[H)8SM=d\75+eJ)HH&N#Z<Z>X4
7^D0,OT#2W_0Of]E>\4NZ_/:gIHX9G+dJ3F_VO\R/Y,N8DHHNT;a7X:_)9VUV9L2
-/9B@)Y2^-ZdZU0g\3=;4Y.7d=>D])9+_fZM@e2?#?\:GFF/B@LLO83BCbKa-&+X
TW/U^S:2,=&4(-E7CEG?f/4H44)Q+729CATU2e;1-CUCBBI>e[PSIJ_T_=A><DLO
fc,<6>7U#B-a>AJXQ8:<B.A>f18>MSQ;,/?e/YgG:fHIQ@1ZQc7ZeQPNQW_\Y02;
_DfNDU5/O,[/F.;M22Lb2&5;RZUN2R>gd5WXebSaa[(W[ZaUaO?AgPB^&<aSW9a:
I^P[YTNUGF_f<aO@\bC/eNR_>SS0V?3FASTD33Y/5H8Gd]TXNK/&R33:Q+AYe+O7
S?178_ELVJGf]FL8@5<;FX@@1-MXSH+BNA<&AD<4LAe9<TG&),E#5]PMF#<EL;g=
\T:/95HgB[L<GbH8^B38^?U<Z_EMH@/DLCLK.HC9bM#RUfN75)7@K=(#e2X?I/_A
O2Y,J0U2J]7\HbUT_72E]f&#:f>EDJF=9JD1V@R<U+=ce9]7KSb1,2GO\0XNg1#N
3#NA]H9MWbTPB[TQV+ZI,/P?Qg,8dLe6gd/-016<7(Q/[Q_XCe?:fNPd?8/M4O\4
?J4e_[E?,=3/L_IEJe,9+,SPW-JgL45ER2(?UU:6+Sa,Ba^VJH/DB(O3QK8DY&NX
6:@-5XTP&[6;G=VZ2425?18(=R_F+gW^[N#)XJ^8CL,X?B7(]/1C0.I)+A:LJ;5K
7_&O[g]3](#+=1g3Z#\=V-eD\DS&g[U#37gHN;fYC<b7?(CT3#NIRK<^a;Z_:0Qg
8&dX^O5b&ASPGdNV>Ke6]<CGdCCF=cBROB1/C=&6HeN@N\92X;gGg+G9Ia=TRG@G
b:a)YB9eFaZR50e?>EJZUW/L1+T?#I:&c_XgHAWcK97\@VACCB?3G1]0WP;R<UPR
0JdBeZSFNIJMD@UZ85d+\#ZEfe/L.,SfbO-#e]G?3P7/FYY+&79fLc-AN,e<IGBA
&G6Z9Y6e\&#,#9>5W=Z)d5R+943X1D5G5XYIgJ+9>5GHd>B+g#[HGCH\W5:JZZ[]
/:FRcT<I7N4Y6?VH>:^a)UX7FVbFTUIg(NP58<BS@HI-2g2;#Q&O5Q)VIfN(fJ2e
BWdLS1KJ(4LQDcE#:,-MQgK5:<P)B[QG2;_4EI0?DP_Eec<aW2gPb8WDX[F3I,)4
0ZAFEdMF[<BX(;V^GX<UWAaJ3(<dS[4F<QFNP]N)+;]_Xc82,2f[>05\[<&YM:^e
(dagZQ)cYJaCL42-]U_&OCP+JR3@PMM[B?.UfP1&0S/?[T@A][?_Z0AM4=I#JC[S
dU1FB)NVRd,@S/6Z7HL;4_KQJS1&Z-JTc?7R>@L(=OUc>N><(G?Jd?>H@O?>9B[a
S;L?2b.+Qe12=-dZ>d3#H=<VJR)@NCeYd1Bf2ESAN-&)V\;PYCT,6&#=W=&^9GFL
_4)PK&I0&H4,acS=R_Mg9DE7<MVB-,JFY0S(#):,@9)aICbgQ3LQY><&X1US330M
]_(UUa?2@T1>4SXe7Pe]G\<LZ..g+ORG@+<=O>:(7H-5]A(8dAZ3/MGeHZT)E<aM
Wfc]=aZL/5:UD1Y4#I-f3\Q4>a3_^U+4L(@#SAXPH8/K^TbHBTfBWQ^_AScOCFRU
\^KaA_[fQ[3=@3:0@J[VP(^?.9GWK[9b^SS5H[#_X]<JN+GM,Rd@BSZE.L+<IaYf
LNZa@X:a0>OZZ(:F?I1>@#?BR.N8@7cJVYK4fDC+=1Y8DZ@.\L4=4e=J@gC\\]/+
Y0A.C3WSfGU\Yd4Va0C-U4a8D=aL40)?QJXJaUE&7,bR5UP[+KQ=C,a\+(SA9O<>
>A?=+9:(b<JM-.3@P1C>::S_DR&A]eCK;LIcAS].Hb53H0^1&:=[J@1-fZ(LP4Sc
,#Qd[<+ZI5+f.KR\Qg-<@f^Kg--XTRD7SG1SR#>[=O9W:5:U:V:YGc.CCNB+:_,T
NUATfL>d9@1/.f>V.c)^]bOAg<5AB#H\J2;dcJ.O2J[[]7SE_Y6ONCYYR333ONdP
9Cg2HI-98+?2SDBV5g@)QK+J/OcLC<X-JP>eGUbF:YbCCY:(RTZK(NZ#gM5GGaJ#
X<;+/LT-DP^f98,e0Jc1ME?N(c3)M1ICB8E_cF@4N2\VS+>-ZT=IPI>7;8MXeI.e
&b7-g5K\#>I+-T6KVe3gTU6bg6T=fB\VK;^g22f7L_S(aTX.]LIQcZ7=&ed6C4O4
a:LKP-#-/[g4AMS2GCEN2VSK?g2/E8dP7f6-_V(e@.2&^X=Ba^#(?V(Z/,R=[a_W
.#D#7^<[BC[]_JYCEWIM<?dPBOe7]T^#_T;fb_Z]R_>80[2_4TERB=Q]6[(3PHHU
E8,d]G4SQLfQ#,cX]UX6A@U:R1Y#7DIL0@S8A8L3K<QIU;BPc,C)UYL)N.Q,W^J-
?U;B<Gb]f+2:<MRcR>+b,\OIMX:G]G30+M[>B<@V(f[G\Q7:P]<?PG&=-OUA@<ZX
EF?>@=eFMbU&M?3fBfG^^C+>\?U=Z,P/08D[-==1bC2-&Ea9fVXW/^^1XKTeAIbT
??g;.dX7:=^^[(/FcTO_TDT0)3#SEAK/0J2+@>GS7WB-=92SBd=SX===6\(L8-\_
d]cV.IBJUGJNME87@.R)F72.M1b8QL@28f+.W]gdXPgN4WbJ_cQ4077g>fFMR;W:
<6#&WD.37,-_93e#EKSQPeKF+@#C.O/IZ(bM5]=WV0./6;5P5b;B(B-8>fPH9H8H
U/:2[<+LV#DD:?9-bVaD.&-.?eX/WE)H1e2VF6ABF+0<X40+e[4?S&Te(921<G.A
RaI\3=.17(OK3ZP1BR_L>HU0^H5LfRZ>75cYK-SF[DF_c\B7U--&M93:J?Y?(PcY
<[.N#&eeFE0<<6B@_:2gGLE,:IFZ/?/>=?^81&D?W?8,/ce4JfY(XD+B^[;f<dQN
YgHZgHI>d(bKMW>a-36ge@RI=dP(ga>bM@AY321eM;63>75d-[7<IGP3cEFWEc(2
\eZOR+C.#9_c]Vg^(Z?VZ3&MAc4W-9X([-g?,9Rdffb9X4JZ+R_0@-LFET5c1aUM
UFL#;OB/a@^]8U9aDc(d5.N_)fT_G+3@(0.T-T>E[>E0(#-52DX2X=9EK&6I44_g
A4gWY[&@VIQ[#HbaFLKD2.HDE8/UB^[=@S)2CQJ7a:^I78;-29.@9Pe5RAOIQK,\
K7_^H)A_HK9>E]1?\.LM\[#D(.,2V+N(K#B8^Fc,//0.0FLAZGB(XCcR6La4GU)4
+EQ7N+I>>CYSH[FCZKP&Y.cQZ8/?RT2(fEga;/C,<QV86d9]>)5D#\[db0RR#I:G
--ZDJN5ITI28#>T0WR\@fdg&2O2NUUdROH,WZIMLA62^/?(.0g@:COUU\&cB,UWX
2P@YO\Y&<TIWY[H?aG3)MH6?d3E.4bJD(fg]F3(7=\GG.&eE9^)&JO5&[eK9[C>(
C\&b\_X?7GN[T;?_NZD_?_^S6/PJMMb8e[]XcC_#Z8Y3^E>:eI[6U9)B0?Wee30^
?LgE72T;S,.AKHI+000@7Df(C]:4?NYBH]-EXX^54VQeG?NgG:3,P3(6WI>./+.J
dXb;#.(QC=RUa>FUIG2_<U,->1NcT[]3D]-eW9DJ2OHDM)T@C+Y+X\)<DHRfYQX>
;HN9JKZ2]2:g/DdYdK=Z_DBGcc)1X;<GSJc.2T1W8?^3MJ8]9V)-R\3RfMJHeF/J
S0KI#A33&.c0[TP4ZQD&D?2&FV_X;0MNECgaEQ=:I?I3GeYBbHd?TSV^19<@(LXO
5a3=<=W+3A7HE^d-.^?#L3I#a9N5g]>R?2BQWcXb<6.+f-QNH]3M,(5#RBP^>2^<
S8E,CcG7VA@+:a+L\]QZB^K2)5J1e+GQ\7dR/)F@DbQL(#[2\&KN@g(1JBJM__UW
)Y97H:GB]OdAPg;7&ND&c:JAc^8PDURT_.U4R1e10#e\=,89=KD(eP)Fc3LQAO_V
O7ZZZC\,S?S:2G[9TSg7-BdHZaN]CK[#8WEBNVf:UfY1\V>OR+8:D<>DV]QM0<Y?
)KF#/E4517TEKGe^)E4+8OSH9G(d9OR\R\6EL/Tc3fS-3#FbcX7A5G45D8MR;CK/
?aFc.K->M^Hf^W&1c#_-6ILQL&^+3[\S&CaaMC\@+EG6gIWg9G&5;7?/IW@a#[NO
+#__J8?<QU&7;#?]NY3V?bWK]D#X]dAOUY.Q&-JBJe>J6P24XaK&cF.0dTZ:N]1b
U1\2DK&ON>>/KJ?-Y@-^@@7ed4Lb:_b/Q5JH?aAX(2QLMY08N8[31;Id8GPSfE&Z
JDP0[MH7VRcOS>5ga<M\@)(BcX#L4J@YBEZA7KE[YT#0_>-QPRSUERA]\Z4(GAUa
WB(d059c8>7KK[/Q-;I5JETdZC-O,Z<_Z^5JN#QVb(Y,VSYeW.1[=)3A.a[=4E-Z
QWN\/+W5FGO3)Mf,;[?QMBCA6DTf)T.8.1+9X^[,,:3H3I_5F=F?=<W&AH@IV7SG
8/\D>@cTc)S\OFQ[NM>V_0[/.1DOcH-J#eYWMOV94Ic7ZYG6LSfbS1>S@NMRa#aO
=Z?.9QYDSHQJ[-A?:)8]aKS6FK2#U#&,6fO5Q_O2B/;FA\9#F-MFdcI6AcP[SJT+
@->S#HX2#HHe]]^@AO7Te1A;R-HAU<g;\S/83169\(I7[R&H?CO\-S/8ba8942VH
-M[2g)\^Z)g1Q13EG31YD;XBC)O3?,SFAEVY#ReQ,:86XI7TZW.EDG_W#QAJEJMR
3U+bbc@-1d.aACNe5S#9S3HFJ=B]JVU&PAgL8c;Q)(fMSA\<\+U>.=W_K9P;@aF/
QSa/3cV\&7\,Kc41#UYPeV3UTHH@F0@5#NSgbK\=0,+G.,c_Q8H\4OSdB(G13;3g
EgM(bF.KB,8a>5).,(=+Y<9^6EH;&c(?YGQK)3Q1ETe1Ge.&.:gZ-RJWSgM02&,S
T1F;7GI7UNgRMY<EDJ91ORZ&0Tae87IB,a=^Vdd/c\BO2:Lb[]](e]<e2:W9,:dS
5OT;2S3Cf--Q2cL]L-7)8=)EFA\&[_BPd]01KO)O.HBUQSN;Sg,3#/dWVaNd2HQM
L0XMSdb>>:fdDA1AecLa8GP=#7?L8Z<ffb5STFM=24(C73fJU#ICHCaa?PHM^ZZ>
EF:F(RY:])gQ]CK[^&4C^W[Z<.<a^QOOE5N#R>FSZB3dTF56JA/9^Q[U^MdTMI2=
769.&5.#Ja.YQ4MT(XW9-f:_MG1HWGCWX?_1>dO7DYBN&I6T<^(L6CC0Af_?O\OH
5-56-1K(IgfH,X@SVXH?CW/&1PK)13^[QM\R,>4:\#.@AC6aXA<_6Y,>OH.@JGY,
HTHPWC\2)TaD0SD528N@VMI6ZQ,F/4##^GM6SE=;H;V]PJ[3Xb9JX>-Rec[:;Ja2
6S1fD(X:)5CR\>R?X26Hf#/;Kf;@(E]LX0-<aDa[B.?LA7>)fR[^D.=)E[bXZ>XP
&O6683F].3?aD;7?.QRJgVD-M1=YORS.23K.Q)7K(b5RT>(=F:JJ[dB&[1=40,@F
Ma@.A[#Vbc;c)LfW;9M].&W34@S61HX9d:gMCIE:;0PK7AAfBg0KS3J/]C+VW?3&
bG2\7gcE:EPYfe]FBS+D-Ja?>E>b,E(I?JX(7O@KSS]ZcC+ZA4SV,2;TK]D[J\@f
Y^13,8=2M:LgT0W#S8FQ2eGdcGf=HGc+(1\\-WT=PRUYQ@=\VG[cGTgBA3cOO[UP
H;cR+B93YR1e_VW.aQ9ZVa#CU.(\<5-/GU)?-U2=dX]^:N,b7)c=IGDN1U)Z482;
+M^f9HC\.;_7D+;X4W/A\G0;OE:))bOL&F6]^;[UJ00.PVM=+GWBD8\?L>9,e6DJ
AY2b^X:fF#=[__a;B3&8X:QF57?>-8DbTe?4E=^1Za,XYc94:X>=Z;U/E3_(DJ.]
6BS)HAYW@?A.\?#2Hc56@9UDJe79_)ULTK><15W:a8.UJ@-A_+@9Kd?fb-442Ad)
6NS^\P6(>2TB<NM2^W/I;T-7g\6bc>J^OKUAO_AY_Bb@H+SgR;@0:R^ABB@]I/Xd
<O(>>MB7f>(DMR(MEV@RV2@Q3N,\81Y.07<T_<64?Pdc^84+WT#8+d5K?e)YYGdI
OG)U&KXHD@APaYO+NSIf=_80a262&A0+R)[.NPNKYC;2C4Jbg@gZba.fe#..[Z:0
;0\,IEOG3S/HJSK-NF<AS_R9>_,T:RG&T8G1=AVC?EU?U4H_Q[_/+d15dbe0Hc(<
L0ZL6O?&^1._7,1+L)_9D3].9Nf[@K[\f=4J)K0?ONSMfF4cTe2DXcAbS4>6Q^(]
N=Y]BGbT+4a3bUPSI/ZB1[0PBe##YU,>bMD=DTF39f<O]df;EbG1Y/]5EeQE:[+g
E-cA\F2)\QY,^=A?NcC4b(X(BYF7AW&04d?TJF^EQ0:7YYG^1BRGJ_SRO-ZK/;EM
e/U_HI/8@H#G&#=JV(T/NFUJT+PT<fDV_6RT7;MX5e?@+:6RYF&7ACN:&UfAL]>)
d4ACEX-CA3W)+3ZBe1?R=DAVB.a(I^N.GI9:#10S\KLD=^4gP9U>b<Lf&<L\G-&S
)]<X>./>GT5XQ\d#dP8NM+T]P</H;O=8E4g;/YYE2IZd]I+>4F/1>CYV@Y=7T6M2
K4<+;X@]NPg1LQ>de8F4:/1-<5L6WX2&_B#(D1M7W1-cfPE:D.^&aW,EYK3D6,4[
<]8Dd\@9e4=V[]g5aZ8YUF_Ua9^9Fa^N+GJ:Ac\b4-DWO[1c87<NMNM[3ZBQ&9=W
g5E&A:fH\=1<TJR4fL[e3HSfJb.g+^/HMI,_0.+S6#YEBLZ4G>3GU>6#gL/S@BN\
bX@>)U-9=)(K09VOF<CR>0T\ef2PPc6YQ3H#LL,M9;=BG])?-0Q/PCWZ2SH09QEf
ALIM)3-H5LJ_H_>Y3c/STUK09K01+PP.QK]QHgC1Jb]R:6?4c99g=c&<:>64&HJJ
)Pg+XLE1_)=IM[>BeEWC=BI9/M_P0]CEU=F8IW\BR(LDV(-bW)OP\LV6\RR:fe@/
S)E0+4cPDW/]]STc21VH)TfXg-Mf#4?]@7Sf<Ud,.F@>RUG2,?\VffD:4G=L;DKU
]&-93>9C7@V.86;3?6Oa[fa>Y1?GR;5fJ)=,J0?D?D&C2.#RN@gHUfGGE#^MU&@E
EKS0069UI.FT#]V(0T2@Bg:/DcT68W,e1^4CL#B5RBDd?G..@A:Ha&Ub_Ga\50?J
.4a1(8/T-f9-9_Pb4]&E&)-3CVXb<RaPP+,>bf(H[4^4RA,V1+5d^e+<cFI/BHWX
+CA0UEG^,?RPFe0XXN5MROf0.7A7,bX<DS:&D5PZQ&#gD33U)9d3ES_10,.4H5/_
)B1W:.)=<eTZH23;MWM:W@Z37(3,>08A\P:]F@36=ED?Vd6bS(G5/e]g;<,)1&bH
#XHA.,I]7-#-[O?BS&H:][WF<QC=O3dV>NOAINF5#3R,5,d?V2V&3?N/TU]MZ6>=
SX\I/3/QRB[[gIU)caJK&)Tb7L-2GRQIIHFS.d3;<:/Le,Rd</EAFCbS<;.B5;6Z
a6fX,JBfDG=\c289(HZM&T87SK+7@9IU-feT?2_?(abT2@#->>V\AS)^:aY,F?\@
MEaXcb>>?UHg7<IV.PG=U1BMYY.FSYZea^gUcIISX;B7Vf+>PF#C?N6UR6\bc^#:
B(4;HHD&5M4/;W^Vf6fFFY<]>5^JF9CSG#JE5NfS7#>DB^6FYZ]e#90)\ZcGcSF4
]]1HDS&=.TQGZ#=<d1gS:K:&:DR/SbD>f#ZHL0T]F&,2c[Wb6Z](X]RAg&S#1>ee
eYS+F8I0(=MC<;eO\-H:]H#TWIe[=B+JcXfIbE6SYS<KT9A4&/4I5d^4=?I2.bU;
4W^_bgd7f&+U&C7ZTgX6)<c7SbF8+5GV&6H^W5_Q\J?e>LPA;WDe&YFYKa:40WV6
E[&QY^3:+feH66@M7XfSK=N\5ZSDM=0E+ba,JRR14eJWe0?aD]=]abb>Z@A;>IME
+T7_Ma3-cNf&;M.-B8@:L]4B3YIQ&7LT4(VNB3B&)<YFdR3Ff1ZP-R?&XMIg35fK
RP^e0\#eSfR.JK\X:N-8?XLZa>3ZY5OLVCCQafY/JDaT[)W]D?2g(Y,^7)U>>TKI
;EPNI>cJ&;2_OFF8aFfPJR:SGXZfEI,VZ2WYN:XIY0BHZ\#0f#TJSc52CQUB44DP
NY.IYaH:FJ)8;;F-cA<[]B,A0d5QcYf;VR[\D4Jc>?g1Z/G_&+Jg\B@(0?GP;=>S
;=3]48e46D;FT#-d+2^gHL>#_P(L0H70=PW1(R.dF@[d/,UHS5/VN=3]GP<VO&[6
Z#7dJWBc:MBQc/YV@RKLGIEe_Y\,A(EaW+Tb)OQf791aFV6__c,OV_<?2e@:7:RS
>;F_(6_ZNP.=]+=12_5\cD:-]ge2-IFUO_39;AF\F/+-Z>_-<Q(HcWW1;EHKOeL/
U0:Xg[\_I,0HbQcR&XF0J4]9TE.dD,O2A0f&ebgP<JUZ<9LD^7CEI,DA+c\.\+^9
e-HD&,J5dTNe?(T;?2QD+#F7Ia&]^I9O0UEJOV(0JM9S)?)&UK?)E^^XQLaLEAX0
QG__)@&?c,6gI_IV8]8AYZKH4;RZd5.0:D;QCK[Q2BfJWE6D+?WXY[MKYO>8[d1/
&(MSdLb:GCAfQ?EJS,OA1GN22gE@J].&9DWGG/cdEe:Q.XKA\K@gK=#+e+Q@J,O8
HM>C@SKLa:)=+8dg<XR:fTX^K#c25#,a7VK1+EAG@a\EV69Gbf5FQID1WH9fOI#0
fDX_0=^KgCHV+]&NOB4LIaT98?@S^HBC-)V)JFB(&+-)=:^cHNSEQJ#(bbE].g_,
@^8C:;^6)C1eGcJN]g<>T(EG+>)/+#WdX1HDX.50_->GSI27RVJ.<8V0Y1VO]dV4
^:OaC(HB(\Q1cUBD0)Ya__FC1]B0d,(AQO6)Vb=VG9BOZ5FaTD1QD?VN2d]PcH-P
[]@d]\ZY7SFdf.#1d(edPP:eGHd<7XX&Sg+#f:b8JUeQI?7RMPP62M:0DFeL(FHU
@gSFO-CCa9]5JeSW14@:=YUEWY=2,9VfGFG?cOR]QQMH7acI1AO^gaTEO^0\X3<D
.DB);T=[B:IY^4Jd=9b;4X-@MXH@]M5OQP;F,ESO6b-H28E5+0H&WX-Pd@<_/2A[
H[)VGbfY+O.[fgeQR]BC90FPdWLH[6W/TOBa#\=;?4\]109?HYe))X4Sbe&e-3)/
K0]XD>G[2e&2#)d##G^7G7cdd)G=.><Pg-CF1PRcVaTQK9J,P2?@T/G,0&00-GH\
]2NM:158([b3,=>^_T).W^f5L33J=N0^eHZ@?(-P>P5cID-D:<E5ZBOHRUI]6bAB
fT-=N2F7(/N&E&L:>gZ:/BK88PLCEYcV4?I@6g[4f5K#J<,>I(McYGO03A3.J#7+
H6cFLI3KGgg;Tc:Jg>HX&f.1G5=fLV0b;U48c=JJ03Z?#4F@)A-5<_:7gRdgC]EH
Ef)aPb-e;W#,3OAP>OOc?F#,KgDBXZOc9;H_(#I#^[1:&VEa0PEDBH>4]:CQXXJ.
+)6eVKO8=H1IU/NUBCe:AB.?SEgE(3fEU6e#\I-?;A:;3]9g-Gedb4@8IU,UE,XI
\WJbScI9[LfJadO1//,Ncg\O,6HPY#cX#bFg0@#_8-ANB;ZV4X0bF<WB4&aN(#]&
3&\>]K>\6+_>UbTF7XT^EB?57H21GKI_6/QK\2;Z.R2I#:HLU>R3?9DRV=J6:<P]
2(0^DSDPK_I=D[.74b=;XLA2L87@;<?Pa7cNUe^W4+A2^Qe4#W\TJ=dH4?[6^=<\
HYP0O)CdQQ0.U26+IB6E\(+/RUAMUeEAH<#DR3E1P4W(?&b33Z6/dCR2dK&BFcF)
AA@980Y?#P)0O6G6Pc41A?2^E5U\KG2.^R#AZM0;5)GZBW?L^&^5N/5J\CJ]+89I
e)-]Zd&NR,]_J:#I>e]VC?cLcYIP]aA,L,6/NeUJ7cg[f=V)MASJ;,Gg,D;)>[^F
@-ga>eBQA040#&L33?cd;)D5<.X,I.L+K:&X@-aMbC5gC0-,&XNRK(\e:_HE1#QT
_#YFDE^IQ=/7D=0(#gg#2.A_0f;6fL#[(^-I)NRXD?YE4^D:CJAZ/WP)JSdZa^S-
)U24N=K6@H(+_K_MB4=XR@)TcadR3:0+0VN8LEg2+\,U?1JGK_HIVN,4:.LD]cA-
AfE8,0(1a15NeR)];gQ;efY_?L-6g7A_F:LN31J4#\:,8OBba@.W^#d,Fe1gYS[0
ZW\)+1)bF\#gHe?SA]KJG-Qg<e_RSTN-&247]6-.MGMb7=MDRB?)4SefTID/f&:-
JOLed.VC<IOEeJ=YAD4001>Y)MZ\V^]TN(cQdAZKUN(:RMb<6Ng8X[e)8M48?<2)
34?..-g)D)#6/#/T,I4TW5UZDW;BSUN=GI#gI-&+ZR7^7O3I3_]<bI(Ub\L/7EeX
<V>3XZ>M76bE8<DLD9M7g3g>LE/^D3e<\/T>:S^X5Tb8L3E\&GT\]M&S:dOdKKf4
(FU89@?Y\:Jc]C@+MX3:M3C;Od-c,1S7.aHU7O/X9b,3+IHKUP@6bb,Q0.,R]a;E
+E9V,cY?:64YcM96=5HCX_V26AdaHe8E,B:.FC@c)a@CJ/UfE,]G9:OEZ99eS?6W
I26(M<:6WbLBU>_@XT)VH5QRL1GcH^6SNa<.I]C<H09,?#O+Hd?PWf^]Aa0P-6H9
))\VXO4C0[_J6.GQSK?e])TZ4/ZQ[?1SfFUJIK.=HNI6WHX8>?4b5>.\90G@(-2e
WTF[R>MYP<TYU0;L:D.FR@(,7=@(YeNF.TdTLP8^T6,\VcU#DU_OROEW<UAH]XfY
DcW.\bY<^;FQA=E]M?VHPEfaF^S&OX5,]<bM_e2G4g?8aN<Mg=;fX\Z.KY&BEJLE
I5P3QV:3Bd^JC2Bd4g?Y5#cUC=XFf.P+7-R@)/@<3b^W>_F2@TN@;Y&UdJ<)J)48
DF))D)Z7.K72E)/UTE,)a7M.(ZcU\Jf/P,@d)/cE-/Z9J]4NM_<Y#AVPDEBY.^K6
DK@6MCE+?+.U(WKJ28UH<6C)D3M1MD+>f@,b99:Ed/K,Cg9aY9cbZ>53&KTI6X<\
71I-5eUJ3TKHG2-Va+#/SBfW\_SZ_e.G8_222[f>139RRCY[=\?IC,T<+_Yf\XIR
KNW[^DTJ;B5g<;ZD&23KUHV-+[@7S<Sa/R17L](73\0+UM_-^Q><7\2.9;706c/e
Wd;AbFVO;VBJKAV@#FEG[]##(-N:@?Ng(?-N=EdT\f/JF]Fg<C56@C[BB7XYV?)9
<?-e#^4Wb\LB_GOE[8-3LD\LcW0GX5(ZH;JFdS30<[-a[I?J7@)\6.eCZH])?WC>
;>R<B+_RKe[f1NS517&S8LgbV[95F,cOAV_fSQ2BFUHd1_EOJW).0a6KT\(A+Q#H
@N9fJUdf>F_CVCZ:7R7L+]a+W3V&6Z7T[.5&Jcgg,Ia&XI^+dGG=Fd1E&:@KdW+G
C4dY2-(9,S@Fc,^.5AACA]>>c2LS1bdF2edHU5/3>KKdQ3<ZAKY6X_4FO+5T,Ag^
e>&3&6?4.^>9a>Y)AEILTg?_2<C1H3SJ\9#S?gE/HXcB6\;.e?(O,+1abD23GJB<
K?H/#f#M]gCE_D&.YE@X@A3T^/EY1IRSRf+O^C2#_7R7U#X>e6b?Ve@34>?_RcNN
4M5]AOR9cAPINa1?5S\eJWFIAKL7NS/6<1V[#e,)?c:&#UNbIHb87@UJ4O[F30Z8
<<:cJ];T4g5UV>.Kda4NFC7)d2+4F9P@J\be^3[N;\DCN?44O,J6\(b@0-S-I,LS
KJV070#=-9TaO+LYKWNXJ<)e(K/9e?+=BFW<g+\\3Z^77EbTaX.@g67WBb\5(.J/
d;5ZU47(W;cU=,Ke2\CO#cW</:8a>Y-gYPab=RZ_VbZO6XA\;)UP3?L-)+,[e]=#
9-COT,fQ\6R,,\4,BH)VLdY_K#HaX0e<JG?@A9AaZU1J\SV>JS&D?L.#O@;Q#40/
ETFM>#K(X7?:EQ;1?J9KD1PB,LUL7=2.0>d:#&NW_J,Od#a(E#>7AL7g,EE&3:&]
RQ-=\/22_)?a)3^UcGdY+5KYDK<RE#CYDLd]<Q+KN=.XAP>6,3XZ2YZA#cOWP84e
JC2<RHF));Ic?g+1X+_YNV&X#:TLe^e40JaLJ)3=:bNcdYf2MU6d&F6.I3#ZJ@EK
DNE[K_3JG?d.NC5bD>5VJ-HK/;Wg.dJ)EaD-F#<OOY\V?:76NN[SARM);]3^8<14
^U&dF+e4KO<9AgNSV:RM>bc;?J,UKH1@Y?;A?E\d-7XKCcGAGC3:Q]??\9#5_+M,
=Sb_,I8D:C\NU/0R=?VgZ_Y:8&F_e+V.DG<aWA0#,d&1[Z^Q?VGX(5,-8K65g]C=
cgRfFS1^DJdX@72P6ANf1\Q-#(-a8[fC)(6R2ZV,NG7bQQ)]eOWS@3Z?NcN^-G#/
96a>Ee^/-JY]BN+N>2b]-T276E/bW_7-^BG?CD2bWCO+b]9\J^MdeQPHa3U3E?-)
XN_Fa(+@I&WWZ53>PZ=:U1Cd=1^f_cY2,aD6d5&Y+IW+@I>JNKFUXB&c:=9I#VQ[
A8)>Q\LgRH0.3+HX#268=d@HdW@SgC[?M&4VB:4f?:S)BY^GE+8[2STPY1:(6)^G
.IB^7U\AIJ&CPQY&0FY>POO01^_3V?d@cI#N77CR487B&R2OIH&06P4_WI78BXa8
8S6bWdB/#E8>5,5de/AZ8R/ec7P;UcA-.Sc^#QS=T=:fOV8<B(GJ08bfE?9<[ERf
,:e;)Q&=\F2<HP1F+&())&K2EJ^I:N=g<_D#Q0-0SS.S)F5\W8\.4#QBMZ,P+P&D
+D(Z>aPAf(fE0KFXHC52KWH#eZHI]3;+#Q_S0W,a8BFI./<g)5).=]GF_2_[Z6d\
f9CaONTEKR5W1S]Z:DK79+<VM)&.UHS:9FfRJ-d>?<d#61&LJ.NEf?BF=HT3X/05
_;;].)N#ZM5&@U9)<#54GYD^^1Db8]4;JOVF.J5-VcS>Q38@]P9?TdK6LLM1df(1
FU6@1M8N07>631TC_4EP0JQ\agKG39-467Z0<B4@6ZZ8fYA1W-4[;#;#\W0c6.a#
6#Id[?/J?OTc;;QG&C[&M,-FT^:)4Tg)+aDaT?,(S[7TNV_YYJ7^>-]7P:QddX,Y
MVH_;^OZbE=H=SNMDa)ON\bPAd;F:)dP<?gB=BZ8Y#OGNNL)EIG1(g3L03BB4bN<
[G;R2,V,33PV.G8g#DNeb5&TWJeHSb_YGVD?+0@g@aR8?&GEcQ:OO?,MWAYTgUG;
#aP_5H.@9[U]0/VQ3]Y514JB(HQ2G/(IQ_bHW;Nc@f;^a(TfK>e5E,X&S+^7GL_2
-e\U[H=U])V)<E\AFWU22J]VXEWVYc#T\:AV)?^3;VHI9,YVdRE(X4T2W_HJ]/OH
cKF?<^H:\XW2HgG/>B7Y4JeSFA5M)f,5;Yc?dEg^YH99PaB;992ZAS-.YOO?CVTE
f3B&#S,TDgZA:WCW:5J9M\))/Cf5B3T@-6LU[D3_CR7NI?-D7ZI,Q@^S@;J8MfQ-
8ddK=\_aBD:;S@-I1=G90TULM10\49<4a0I,)1W3WKX+V[=5D,X<EL,/TdeP:a>f
b#O1CM047bT&V3>+VL#AOU^OJT[g,SbXCgaE6QXB:@?2D1F8[>B?Ae9D8EHZM=6-
\+H4/FARK_W:X)>?[Ve_(P,c./YQG937\.3+H\5-BEABcEceE&J69LIN.H^;IGcM
a<N>S.#DFHX14QWX7VYJO_F;GQ5Q8M+C)5;?967cTNF+^.PZf\C]#66eQ-\;dg^[
eVK\(bK8:-Rc?_8UIe4Z(EH\RE2M8>RI5CTe,W9GWGL;4a,bY7V4BSDHYO:I:H5P
P&7I&KYba-UDH/U@CD^R9J+9KP7:U&:aPdA8Ec;Z(OO.;e^VTf]DO?X0OXdaI+YH
)]E)8UH2JgD+BS]cM?aD-gf^11N\ab@HTPY(Z.B2BKa^,3F3/(I77GVQfQcI;Z.8
5STg94Z&)0/F_8Sb-g62,[+;(d=,gXO1)a9Z490KDdg@C:#+08]5NTFNL])>UH(>
d-,B@HHcYR)^&Q=,f[?]?P_fK(4?<(]=XG1COTA(BHVYEGa#=(c6b/f2+6dH7?GA
4I2;U:^E>d<DCbGLf>_B]bL[EJ5Q6,e?]N4^;5e3W-I&?>?ZW2<gDc-.-H>O^N+F
a-&T&)1;,8b6f#FV:dee^V.E./#COH5-Dg)YHX&&ZJ7BFW,c,_A5)]5dD2#^=dB>
^X[cVI?5L_BYO@cDY15I^LJ#)JV8:PAEDVFWWKg>Z(VG4Wg,+3WZI?HGbESR/<X8
#E:RLD5[CL;KP55\8=28Dce&CI^TcG(^AfA>YR@ZBgVS_R@ffC.\:d</<L0QOGHJ
+2UUG\_T\a2A2XdfO\F;NJV.CO4+#EB@A1;2gZQ(.NCWZAC)Y&W3WL8bTF=+FY_J
X)\B(>9_a]8[D&@.]b&E);X]>aCI,Ff1DG]Y6g<_X5@]Fe]GNP&dZWP8[YM]30Za
:M_V<_7HEWK)/d\_X9J+5061<,CG_U5KC</7.Y+HLZX^cJZS>W+f<AHHG7@eR/_&
._K8,XU?f7_Z<^8TGZ9+9;OVGbV3-c.g+L2Z@_NPgVB1_]DTFDIg=T2[GRG[e@,6
48NS8DQbTBEQ=/C?_4:HGg?4[(-4IBYeS>__QU0O7fVEf^EX,?1]@AHA2HH-,LbF
M63]SS[_ccQa9L?AGa_:LAd1^96NY<O8(SReUW,f7fVU3M<.+0b&-@0Od)=T+XKT
CD[.,X:I4:B3DZ5GYT3Q8g+a&Q,#gUdPgXT;<f0AVMa-B+=J)T8-EBb+AU)(W>GU
c/9WCPY]0E+J8=-0216>9#P00Vf;\YTONK>NVXX(4bFSFN6J_1QE,=gc,/T,.TWg
+\;DG?e1-\cK=SC[U_NC7X=;;?8)<JAXbDSEZ9V<ACZdD18S>[+,^0,3YM0Gd,;2
-)SY?)6J396:cSB;O?=Dd(+S-I)8)0O@^^W;/X_6S<dVf?SWW6OM__9a8<85[G,[
R//?1_&_#;=(3D(?N,C59U6B3-CHXd_g=\G=>Y))_)/60S#ABIBfI#ab)^GY3?5;
;4)C\N(G&1Q_16ZB4.Q+JOYZ[+fNFJ=&OaND,CX\CQ,2N3@;UR4#g[5@J#TNMH-0
JT@TeR2-L)[<Pea=-B-R2N<_[V.CLeMY7T-R4/30R?GKT;;S;B;];:H<a\X4Q,aE
5KeFSe/)XM6b[^[DO@;3Z8;7L&7,^XJTVR\P(O;K_U>e2CaIXEbK<=&-IS66,S>P
4#,=+@F;\0QL-,gOC_K^DN]G^&4)F52f3aU\Y7T43ZBE4CX<&FFWUH/LM9f&]5ZK
GT.HNWI8\@U+QTfP)J0)FT=1EN:gF@,GD)(F=L;7V/BSSQ/P&78D.g,X5XB:S)F[
+B_B=PdOJW&T2ZU;5+Y(9CUf+fFBL[eV&0O-QNb:@gM4<W2^:VF)Zc&@(T^3MF0(
]CUT22Q@,ED&9^L-0\6X0[c&fG2^<B7?M7+?V((OWFVPS+g&K76^XDdf^,9_:)PQ
@9GD<&KZV],FT2Y;bg-4(0CL)5d5EB-YP4XS:80/g5IZNaES4bZWJZA1GV@37&C7
8D_:9INBUK9+#LUTf#VEC2fPN4W^HbcJS3(>ag:.-^=cO:F4:)\:TAB\A[A3PAe^
G+/[a(E39,I&T&eGI?AV>(4cc\bfbQ02+>=c,L>9eIRN#.9WSJWB/25.89R[B(Cd
,<dEF=+:R9d#T8S1_=@)\DY<H\2H,aXA[ZKRfYL_bY=F#G:THg+Z2e5=BF;5AH7H
<ET4<N3&SLR<-)AK#]G-_SN.IfUYGR?E.0HIU#d[&N:Qad=eM[#(g@G>4.dDM3K8
09ZQ/-;daU7[XS,WBGV\bI2/;9HF.WYKYcM_G@-EY<O0&HT/HC-GQ,,/-SC<:=<b
TT?\=&78LOfQa#W8fdCL0gNO5VRfV<@45KZKABe:WCM5SaA0KD92b[1IQ,<BaQ23
)S6K42QZ)Ic-Q&D.-P/>7.V<>2(=<N[@N+JcHTKEJR<_OXW6W(K?-O5@?.c(N17P
3DPebQ,JOg5>R;>I)8\.cXg.]9.U=XPWQM./IBD2MfM;=-8ED2&R0<<W8?=]=-a4
<Hb=941PY:7:V<LYCS>_Z<]=1&:Xa;14?Vf2J)>8FW_4cRGZ>3.XSf;+1+>(F1[N
D@EX,ZcN[FGQ/LL_6B9/T;cD_U(5HOV]c6P@fV;QJJ?2gV3,&XZ_BX+#Z:D&ML;H
(84#Q2LQg-aLBfI]:8.:F0]T>[RMAQPY[WegROX^T3<Z-73,GA?7=[]Hc^W6#?eM
0)eF.#d#TFg]dc:AR8JbD>)#7Q8?&E<0FI6<98ZH)2]L1B^_,b5P_=_#J(QN<OI1
O>,eG5.D(B0)LU9#2cc-^dUCQWcab>_=9-8&f/6Ee4GDgW[#E5W7+c6WW/6ZM:c,
.0eNW,N1I(&TVK+^SJ<D<KdP=6UIV1F:Y0SfU/NJ/-U-.9X6EfI&T3><UcA.2[#b
7e)9Z=)[dc;&a#Ged1K,80e+F_=SS/5P^Vd@6X=^^-+gA+]7_a#-G];)YOe)MacP
J#NYJ+8Zf6gVMa0B+>0[RW\_&BTE-UV[FeQ#>C]I_A7aW+3)>FR\dI>8Rf+M)[Xf
FNVeP8[EM)@dHb..ZOQC]MJ:?H#4KXU+\0>^P#[=BGQ/ZFWU1R])#+PaCNDDa&Oe
J\5#\Q5;:MB=-A=TR.?JK]9[):>AT.7\d2WB^]AS5K<?c=^1KRHW2eAdcc,[T8L?
;IQ=UQ(]\KLc+dDEV6_LeB+BcX&U^S9#FD6,fLd.UA948\ELFRAcgS<9GP;L\^fc
(VO=&^[RRFAA+S=]Q^^Ca23U=YZX<MHbH<.Hg5b7\EG[a:dEZLPc.>6cA#AX1a#f
&+7FZ]_5^1\--&bYNU=]C=<3)D;Z&f4/7,,=R?B\]g==HKJ^)T)8/0;9,edIf[-I
eC#9SRf@)H+M-O]1\7AG:(6aAPgD;SRA7I0_b;K7G]D@DJ7=[NL/14Lf#<#H.5[<
(0>A[d8CQX9K9C2RGR6DV7;DQ&I@/_XGQ:PPGZU1/)(BF>U54TS-8&]EEWF#&E+0
V>P+d1.PN(>c:TcB&][c1[8Ld/A4/&W_7de2c[GR5BJZKL/X(U10+70NAgffdNgL
9:N#FN@FBI&QSb9PPOXA>.63dBQLS(8g#\]934M0-N6:@d9A^.9f?:9T\Rgfb5\g
_RA(P0=JFKG@5:\Q^7](JSGEB8aa,=M)e8_QQKXSg2Z[&ZPL,QN@#Rc+RQg[29T5
8PMLZIc]U^12,/(fadCR\R<+g5TF@CdcO]8O6:7d:a0K\bPe6IRC\CfECW,.@f+Z
BS7;K9#d,Z6dQE5-.f,f</C)O9#XC3GWN_.7QY+4\_XPdJZ91L;KNVBJfONBBJ]H
gd+bWO,D80/X4P>JG69\US,\acFU1H3e#fW5aS+8A,:,?EA7&TZE^W1AXcCc?bNS
/J[#7O6_)G-Rd@cA?Z763X-T5PQbg(&:XJ[c,PF(B8L,YT)PJQ8J&7Fc#/[e,(2g
.XA3a<gcBa+OaF^?0NB5PRMIRZEDW12][I#@Q^RK9QNB-a&R]<;f+aZfE2=EOE^\
-L@T_cf4P^U.J#IA9PFdcFMG)<EF+^f(J<dU0e?JIeGe=Oe3Z_BcAe#TT-(#^KCJ
=@\(03VeJ=]:N3c=GSNBQ=D5gdB[SW+39_=K9HK.]B/V@+6)\F/N)#VKRf--;4M-
Ra;&]2RK3Ga=/ANXZ4:,\R;#V#EH9dQS(V.[D6Ie)?Ka,O^_d(-[aXCKJ#@Q[?QH
ba)B5\0Z8FMSBJ-MP[M+fWQ#EHB.9=UDedJ;1IMg^)UV0IBQ;]bXG._&AgV/4T\U
c6ZZ1O=<[9X._3TLC?7=J@85IMD8L2NLBgGgg-KF@V,#V]6?fWMV7#+e[Gab?@[:
TG^_=\#^aC<C([(JMCK-<S04b0LXMFN--[egHf^a8NGgL)EFb>(BU)7#@KD+25K?
gHCG)g?53#I^I=d.ZbAP&F]7HbbE2Xe[afV@>XHA.U7U?g#e#>ZbOUZBJe+UaK[<
_7+TH1^ZbL9/a6[8C5]Hb#LMS5W:UHF#7^[L6BND/TK_)1eQ3O?ZF0\F@PONNAfQ
IWKWEG)]EN&C0<b:7)0]E.F)Vc9N_::I?&D/Pe<J((MBG&AGb)T1^UVN.(>)FXf.
)=Z0L9F8eSe+^WG>ZL@S5(D)b?b:]R#L4+)c4\7MXF3(Ff>SOI6S_g>b3B3Jc1Bc
ccMQVE;QQbLa8M,3IC&Tf.a^DeF5L+GI,081O<-XG<=1ZXY-I2B=+(2_+F-OWD<H
AF,J@H8TGdD(d@&G+XY?D3)R9F.)EW]KRZVL6>E2c^Y\D8Qf@3+6?9L.bgd)A:eB
R+4<#J204.8R=9K4@??B6HQacXADRY36E?PZ_<8],=8Ff5ZZ2WL#UQ9b+^]E6@9-
^>-5I\+1.@bb:+S6,SbdWc^?Ncg>6M4C9e)V/A(+[=ELVCK0=FLQ:=aY@>gg1^OJ
1B_e,E?MZGW:JO?K:3?#\3KDC]\-JKc;X2(0Fg#,&<4DJ9W36A,gM.^B)(Gc&P8O
>):Kb1@[b:MTe:a:3M3O-fOVafb78GTXOgg(e)X[@Q(aRa[0=((3:5RO/?PKJ\_<
5:aX^+02(KL>V77S#TLXQZeHV(03,]/VfEJ<81+B\])-#8D)aLDfI&HF&4)/4&WH
W=GRaQ#[>dC>?[PW7dGCWX/b??@BNgT3Z@Daf3.H4\Z>#2E[TV86=-e.H_F[P8g&
NOd)\WVKWcWR7F[_gFLXLOZ44D62LUYID\JOPBH)acYK9;EOX6McFRL3KOW9B4)K
^ZNa.NNef/fZg>[d;Mf5U8_VN3H6adG4>/9CP\0\GAT?07GLXMSBC\+cZIWYTe9M
>6^0.-a5P?]9GFfL=TB8g0TZaI;B\A0?gRH@FYJ=93[M6P5_),G17UY0aVLQ6SQ<
/ZMOY@Z972WM_&@K[(K@aBX)H-<6L0EQOEb14S)0)b0O[c=AaSJb4JgM)B0a_bfU
FD7GcPU_Q\&[A_.c@B5.M#(<FgZ9NT>_N.+5Jb_&QX^B0GK#X=,_NV+NP/#;K2B=
8.^bWWPSJR)JSZf[1^1]&U<;W9JS+AY.Vc(=J&b;V@CK;A.6\d7;f<)+Z<AV?WRS
4SZ0^4WLU:G>&;V#.&U07Pd#FP[CWW4;S8/-\@9Q.]Pa;,LH3-Y/3Mc0Nef<[#72
Oe:B\M/7@e\eKA,GaL7cM-KaCeNLecDE2^0+b.BPW<W+[)8THO?e\Z[SE)9;9gC9
_H-QYT4dJ2c^N./3[FK/RC:#+1F_I,@>&B1A>)AB6#I:2XS(X7QLQZKMg-+XB2=;
)2L:&g18cU5-/<IXQZa1CC(F8Fcd8E<KFF&Of\D(;)1P6bOSf8W?(bY=KJ@-#3)W
PgVXC/[;-H,NAIMMGaI38O2<,bYdKSOdLKCI]+Rab,6G0cQdF-IG#bd/5<],=7HT
<DB23=,/BSG1P6/_f&Fe^POHICZ/9c8Bcd4@BO4FL=JFYAR+8B+C<fJ=2B2K3f&e
=b>P;(;>:_F?GZaSHX;DcfVAX/:,,KB>,@&AZ[=MQS#_a86+PH;cU(H>[@_L&(J3
P)3&,N6[/:Y^W/^MB1fVL^@42-BB-(K6YX-3=9,-3/+_8F].8_R2IDdD&>Z&cA<Q
6Z4Ke<WNMS.dV8PJCcC@V/#WF,Q+T8R@=HL-bY12@CRU==7IS0S+6R@Y]K-/FU#U
c[PMSRVYJYCM)=+VdVX;,[,gVN.KX[\3Z/MXQ>@G&=@6Sb\+<691CaKE@M]QOGN5
N(TP.GbePRUg&FI45L?EdX<R@8(g5(Q\,.2AN#9RF^7#>Zd;\UD_35bg.T1,<U@0
<3L[[3=-X3(TeGMAd\YIV>e6G,e_1:ER^GHDd..XV=bNAR>Ee/V,7==c+OKPR/07
PMf(dPKJT;-I8US.T91O_K+J5;f&90X1B&K0H+e+QBXOQ+_RBQRDUQa^PC];GNeO
A(+;-D610QKe1=]3cZDJ=ROJV6Q<4D64TVQ]<E)3@^&Se,:+JF:\V#,K7dYd3XF;
HK:WfJDZ>W?:Uc6:N<CLDNQM[:1VE)&09a3.4KKXS=V]LSI=P#Gd/6/5?8QaP7^B
;+W\IOFR\Qe_Rb[6RMJ7;R<(BEBU1-8OeJEIF[_^Yd?)MSD:XbY&La;>)IDIaVS<
N\KSe&8ZY[J62A(KNSQH^gX/2c:eTb_Z(@Kf\,>PY7#:=HDB&/:7cd5+S:&;CJ4<
J&=Q=P(4fXc:@d,L;.RSVULKR269S^Y779D<1&&f4GQ3VE+gU#d<=cCTL.01#17,
?0E_c3VCE1VKAP^\ON;aRUU9L)BVUeO]&:dGOaI3)=J007NXW-+69bTOB;NgF]a\
UK>/0EXDBfHHP5RV)_dfNDEg]L/>J=UEV23OJ9M:\V(/Jf1F=>9[@F=IK&B;:4,g
V4GZcd5)+c=Y;#@+V4:@,dV#Y\KYR4Qg&4d3PEKNBf]S]\c-#E.DA9E3L^MM>ac.
CLV<FQU2Uf^&(Y9><90eFNb2=0Q<7[;WV&62,_P,HF+=+.7J,Eg:bTB5:gB1O,XO
-d3Y[0,4KYQD,MK4/fMG:WgZ5fFF#R1S)Z_IV@<HB;8WWR[Y6T=.MIHXgIXWL32P
f8&H;-55#bQB?SdK4Ae2gH4_B5^&Z&b:TE9cY.J)gUGQNa.9ZF84-_dIS[ZD3PJ&
,?TS?:Ad\&H9]Q\SK?Z;AK5Q02M:,1IIS:XU2e2,#:N[KRQB2/F_>Y=gb,:YfY@L
6\4_GI#TgXT+W[KJSNDTB:STO,Z:c@<YcDcLUV97U[\M^g_/54aC:g,S]&6F@,S/
KaX^-WXQaL1N7<Q&J#L:+&,7)MC=Y(+&#Xb]+a=DQ,/2_E34EHT3e5c_?:)?(@])
86Y@4P9S0;dT8U]F@QZ)>RT)NfV)2QP2&A^dZT.I^H<1DL,Dd:^eSLSR4>3>dd1S
bb/ULd9V6&MgY-57e5V9IAWMSD?EY6^SJC=?MRA3]E/;QG6dGZa_?OM(5GD/,\BZ
;)WYa+Y<d_CB5C2OPAAI\PH/)UeS.ZMCW\2&C#_NPY9VD(NaD-@dHZHGa:5-)P]6
PGQ&2cN&\Q&]1f)]_I4(?/]J^b=#J7/f\/SW>Z6abg4aS>RfE1_g]VYXDXAg)@)Z
L>T+VZ2XLTFX&La@TFc\(,f<G7^;:4Q:dQ-)VY[RC+GQ&(&.4YT#IP,(;&,>TeWE
.D5E(_:[@-BAJB)WG64Kb@V[V=)>Re\B;03&E\^XZ>JNg<<5b3><bdC6X#PDaDeW
Z/D<?FOIXK9#M81O&C<]8DLCc.9&?G^ZTTU:F5O@AI24YJQJeS3C[\-LA_DL6TW6
(D99.a7cMK0RD;f0X>[TB>\dM+DM0T__OLbQ;<;^76@I,AbGdRCWg<M<-bF^eeD>
\I1/_=f2VX,Z4?B&^949]8?K&,GH64H7^T0B2OWYBQfR82C8)3O/aVeZ4T=,CE6)
,N^09\EB5.d.,3((#4D4JKZ2S+gN/614&/#RX]ZGDCK9<I)_[YT05CF#LEUBMMFY
eJCKBU&-T+acW#99f3\H^.YPY<H8M+I8S64)67\7(2e:7I\[_A30^3HEJM11e.B>
gbMd)N&VBLY_O8[D4ZH_NVU0cVZGK1I^,+[P4e35EU+T;J2DT2GHH<eG1Z4DgBIV
a#7L\bY=F#:9Re1LX3TT@R1N1\FLA]@VZ2[1aQYI0P_B_KAO,9QQ8AMB8WN0OIR;
SX^3+@A<d-K#?0,+B5<;L_RXA8TH+_cba3JNQFcLL>K[bL^-4@Qf=_6:9bFT4EM2
2UC\5L27Y9EK2c9\7gT:2&d[L9)L0I<8#;?J=(/S8+X_BC+7P2D8B+QX8U-OK\Xa
<6\&W_Eg8c6H\0T^Z=Bea@\#e=005FTZB0[,8;G?acCXN&)\>ZLEa_1M/JCFDfZN
aZO+S&)C>_P0+B/.bAd1-J4#=[(#Q-SDYPH1[4e(eN#N.4R<XbW/.&Z6SI:BWa#3
2//^63X9@-JMaeI0V.06gb^2SJ49bHbDX-)M6dM?#2L/=3@H5>8EL6eaf3Ld5NBX
M<e?RD39:cX1fNb?C4?]K(I-c+BJ#G4W?N][@RQ(ZCX@eO&#f_=ZbBagOg=\b_,G
R9NUBOK#KKB_N?TYESW:.92?EB-3KC@G@\[3bU?6R@21C4I/OJT[OD8dH8)a#b5O
:S?OTIDWcST;=VJMd#<[WV>4N:KL[C)Ge[F:UOXI8XQQOC16&DP@6JNW[H=Y1;;Z
=;^T?a1&_F,7+f_AQfO/)C#8@Kg^8B:\;MA]B+:SPP@IP@&Z\2A251;f-2/6)TOe
a/>DU.Yb.V>FPIL6_X9K(V6LEW)Sa9fWfg9T.\PHZ>W]N/]=6ga)^U:EYeZ:7J?Z
c)UTJf3I\]K?2T2:0B+X>&&D,ZSAfb35HN?b&].P_c,X0_f_/B>J08?_;U#<;9dZ
74^.GNDA9cP<5YMKbYMfXaAY+gW@,M#@.&YVMVW)XXP_+SR_<bZP1(.(YOL0L5M/
(LA4HV8IB56A2M0,-_E]7?::.WA/[;CM+:C\6>PJJV=.(IPG83N^O+>)WKN_]5;A
XFfW4V1GIAKE3f&U<2JQHG?V/VJ-D)XC/bP@0G;I7B65CI\?))(UeC<,E&=GI3,b
6d4DH@M-@>L.0acc83=3E#e0?M0;:X:TOGOK6Be>3&M)6TdC?g2WYQR2]O,+H6#a
&#?JUg.4(R(.BQV94UdX.f;b.e283QGFD/M4D^B,K<0CTLC/Oca@PB+@P6.X.Qa3
<IX<NY(;T8]U-FV.R28+8U=e5#b^WTFa0^5]K0MQ^^T[(0(^ea6EST>QQ#_9EQ[3
SMc1NI.H6.RHD-#EeE(R;9a&BN;XO-BKW+?XAXU..Z[Q@C;SH_[5bVRd1W.(1Bb1
3^2Y@+M>PL)c\HW3:FPZ+7P?L:@YI&3H7dBT&V^:N37WfJ8RS7Q?LA.3]F,a;-bb
UC\TdU6Je<OS;JZS;V67;0bJD1WJTa\)Df/F2-B4;V_aHR1??7Na+H35:41F4BaA
[W1K5gBaR>C#8O@)>AFCKM-e9AUOF9D73Z4K9;M;Z)8PUX19>_Ng7TSa6L:QCRgO
f:T^G/;T<ELQHFfX/&>)12]3>#T@U&:&#VO:;(R)^-1N#gaTPY^&O\dYb_E1I7=R
96Kc&+R[_?c5J/^.H^+)1-1__3E[\9HR_.V,Ga&;_@8-NH8/]#)fcD.fX&AaJ8WW
2+[@SM,Vb=]F5KbMa#GTdG?JcA-5V,>U65HIHEF#ZaY=Ye3&+VA&12#;1e=+AACG
YBS5/O7?Xb-^Kc\@&:;31g>0[?FeSU4Q-MW/XHNBGOYSe4IHFNX1(>6:[Y5=58^4
#D_Pe(&X-S68_7EA8B(-=7J8)KB#e&.I=,^5.GX-Ae:8eI&NHSa4.aQ]-P>(c[P:
/PU#GHRB+=dbSPJb96K3CYBDLX\Y4e\6TQ19ZR-c?79T-9,\Ne;,2RQZdC),9KIQ
&/G9#F7V[.D(]O>0XZMSe.B4Q:?LI^0>[G:dbTP-5Oae)gJ_D5-(NP2?EKA(F:[9
\WOd1;K(eXD?D?AB_>=9bd@5G297dH>#OC)g?\PcU?1R?ONU5I8f->WZIIQC477W
a#^,.KHY=f/+U.3cRYg?)<B<Od9HV(eg^^CYX<AF@.\^AIT7GRQ\E8R9Eeg4[Q#d
Q[gI8#BcU?\MT1W&,A/fWMH>\Ag4-[\(,Gf=V8,MbM:ZU:^T5QGPbH+Fe94G]e5T
f/g/6dM?f(]@#LKQ/b+1:<A@\f+g493O#b/R9\4/AgRg9>:DW7NZI8e/ZQ9Td_]Z
<.\<-?.gUHefU^_HZXP.6.->N-(QDV+)Q?fLZ.W..K9Hf9A+Y9WBPY::Ya6YO#J2
eATE+PNO0DAL\fB:J46DXJB9g;M(gDDbU02XG4ZaYA+LFNWEM-3gNY9<DIH8L&9I
P@ORXEPLS;8FO]R[760dZNeQT-@K@<dHJ_MDg7>5?Z79a^P^_YFTP>]Pd1gI,Y0H
WRN+de7]OCMG)dHe(W0:S5QGe[QH:ReK7]G7;<A#\XD-4WZg=I5+U6=SW)HS9TKD
+DLRFZ\eHU<S6GI(BK7TD40VCSHe2N^2fN@>S>4]MQaP9\.B0e=TJJ:a#g;-\GVT
Y0LS]&aM(9gXAUPX<Ocb1_AfgSR84)GC_FY.6gff<E4NH2RO+>N?0C<FMK1_+U9;
WeG\T1GCY3/K(,7dX;8.X3+J-^Y,e5LU1PB9B0ZNB89fP1B(5:P3+O7&3(+&HgPf
e61a1=>TRO>C-N2L#DcB]CBd?c_Q^:GU0+bL/ZBA^c.8)>S4_\RF>Z_[\KV(_<E]
Q)b/K5=OY=E\ZQ<0VCZ6E\\K>GVNFU;3,SB=F0G1CB9T,f-7:D(N;7(N<VNQSBVA
A1,S0-80M9(@Z:A-+=b-YOS5:R;EM1D)MK(ITg1J)6FdXZ/8_Pb331R6/7)J[3T[
](0,@;PWFZ@8KgZ\M8,Z@D+A:,.^?ESg]LU1OLbE[J;??TcaCRE8XU3F&d<X8B)O
-+9<Pg6aBV@dfgR/:H&X6<WP5FFDC_3X[6KdL^,&G>[:eTR#B>YAaYSbVJ/[(FKX
b0.aU0@NbN0<e<(+=8F.:S9ZbNYg7?S&6B,5<+S2KPc:d6e=]+VT6FcP.PYYO\<b
\\KBX2^2QG/:?fH5fJUg.S]5BZCMG4^.FbPI;1QKSEAXSOYN:Bc<N<9;L\G.3fd9
f//EPSE[eed3I3UDc\a+\#Mee;.?+L+#T0,U0R5699PSa63;+K/K7egDdQMaC/T0
bN[Q(GN9JB<WRWcH7JC7,S\KU][E3(_.TWd571:^[?Z>;<C2B=DR3X/_#c5cA2f6
SJ)fRMY2H52&/U=aeWBb&G1+fFLO+.#0I0CAS<U[8F_TCCgKJaD3Lg+dcS9DQIf0
^]0;_Eb2Ja/Y^=4U6bG9CYIE0Kd75a=@eNIDfN;bV,DW3+19=a)#&Ga]cc2-&(2+
,71>8Xg]0U5J4<DXF1XIKMB90RfWN2@QSAeAD4=GeW\#Q@#,)R_GMdIJ?2@,8S-;
8da^C&F^W^,4#6]2AD<a//daL74VL6TgF/Kf)2_ab03]?/8dP351<Ya8^+U_VG@f
IJ>bc+Z@[E/-:b6/A/5Hc8=gf:f)g-98eL]G5A)a#c(I+JQcI5VY18RK0L.(MG:-
L4Nd1e;EA:HE@_V,YX+-7]DH#F9GH[?YF<cZ2QZZ1#F^&P[N6aX)aEcX1KA;,+_4
?L8g/?3.Z79EPX,&8QITBXDNTY[5I.SH?B)]32=a4A:I?X3^@\65(e8VXI(JQ&N8
CV7=8)d7#BR0bObAeOcM8PO4=CJMe,d>68@LX@KM2,H&2KVWW7U@VZ++Y[dGX5P#
=M0)CEU23[&#CF(]f/CMLK8CS<\/^]#/3N7K2UUC1#dKRaLV;Z?d4J/TL+]WUI/J
\16HQ^@\a2)SgIZOYXeb>WROQ<>3<XA/ZA02APbFa@79NC/#Y;2XRGH8?&(D9F8e
e>(Q\/1R[KF+<]aZRUX;[AVIF8H-;F,eG.Q\=FI5eW<,@R#^SP=Jd<QKWF.LB?YW
R-2LR_,#\I5&.S6IgR2OIF[:Xe:d+gUR</.dC#EACHPF<(bWN1XZV<>^Q&f4E39]
8c-V.\_QZ3WFAU?;O:a-Y@0^,&B78]^)>HfA>Z(?#e2>HSXP)E&XQcN@<<U\[TRd
2=:Hf>(;gUVP)Q7CZbfS7gF:QCg:+>M+N?P2MAWYV@5XIH2RU>B-:M@.9Nb6#=6+
=)AHU5,eeZIf0)R=9Wd??b^RbA(-P_fedC6\gKCM8#(GD]a4a/;I;DCf5F75TK/7
-Cb6BCU(5),H]-DGd1]e&O]cT=>@>Ze)[+=LM:b1b@,U6UR3D(X,(SHZFHEI>9Z0
a_@[9NT&/+VOW#A)XIg_dT\G/UBV[=J-Bab_RAeG5>4H,^<6DgU:Q_.-F^>:NNYC
L?&G0C39e-]a,fA^3T\a\a(<C;T:690c\7O=HEGBY]MT&?;LQ^1&V6I>UHM<].c.
&fF3[;<Cef]O3^.)Ge),Be6^1@KdbC,JS=^Ub=LQ,>3T@GfS.GU_dQS1YXB&6APC
5Z[+1I180dO7H]1HaMFb?c1BaBI#0Da0/Ga,O?dcge/#8@^CTc[N.6YZ@\]R80c)
SNQMWCSN9G\?]fZH=3eIcPDP.PYdAdHf+3=?_+.H.f@<+L7U;;cNaa8M;IO,7QCM
a?7ML1W>PW[b(G#XA[,T5DYBL&2]H=(9EXaN2f_S\#&\e.Ca\ZfeHV?Ug,F_bUfD
3Qf&MD^K.?8-df5[f5Ug:b=#1DIc>U>PBP8AWJ3E[WA7TX-([&eLKgZ[Ic;@9@UX
e_GB-ac_Ab_P(e+Z/eM9Z[Pe6LQM+aS6HMd]a0U.>8R?FTfN96dXFFI(1KK4,[4g
TU@A+GS=(&X./e\e3?;65NAMEa=[g9YFF6REVP]/ISW0cTC8HR=S_c4SF\R_>6__
c>TUX/d+NN3Y8)-C9H5D2B1K[<Q[-2B8;PSQ#\/FD^K?UFA-+:>^)<&eU<(>_F92
CAD>>]cY6d:&A8E9FOc:3^.#Oc]Pc0T>X2=0@V1.;E#0@4P_6+J0&TF3T<e/WO0O
N4fXfA-=M??JI<-XLdG;T^N;9Fd-=W6[HH;VN^@)F@IE3<K:AfY.P.HS0)Y(N/:T
f31g2dg(?2bLd1V-GI9,IBc5,24:(fGX[HCgU>#=(MQ3CJI&cCK1GX;^/)L^DD9W
7KSED53/I_[Ce#,:fZgbEb/FP3;[8cW41TLeYeCXV^VMdTUPB+QdP&2C6LG&RC3;
.8;-NQ_(76<E<8_@Yaa^6Na89/.<OcX=2-:>#Y-#>@dd1VeVS<#;-W1:Q7[)@]20
A9;3W6#?REFQBgJV>DG9SaC0,6aF[;VG3=D-NF^C/dbY5JJ1XIE&^HB(1;fgV7JV
.:P+/3O&08^W)10JE3H2.S/H609HZ7S/>PR7?bdK[RW]19>Ra[N;=X^:eYN,Ca2_
S6FW5GFR.]=cH8F,.<#.KVE2OeSd(OPdR+,Ue38RcMR?fXV&;1[DEaD\=MB[.d5]
/MAb5+d+T8DG3=gbGSd]-Z6TILDb?@G]gN<@A@JJWY@g28;(43;Tdbd&c]f:SNed
@]Y&?BK[<gGB7C1>2LbX_>MfYD6M7HI?=&SX&=RMI&g\Ke4P\/)I(_+G0U>ZJe=E
RSOKT)K53O6[,JQMgdYe[_L/YDd,4L6N)IR&](4Lc86/T+A2G?g-ARfAL\-H4AcI
TM]\2LRC?::e\^1OLM9Z#O]@0ZO(W+8bXd19_+b^Z/)N8F77[RbVgf6A.R_^Z=VQ
RVdM:EH_a)MT?.Sc[Ce@K6H>YOV2CLR<F;VZ(SX0Y4>,GTM)@\V58_90;0\P^De&
,E&FC:.dY5IbXGc]cXHe7I=I<aHOG8D43=3Jd+-gd@XZN[aVE+OZTFVM5:^^B,0K
?aZa>_9[TC=gCJKJ8;B/??O7N3Ae:/67;IPeFU),77DgK]]e_T&AJYO7/ZZW?XEG
,TcFf196ZeTDA\b[,g.?-7VLR:R;#N:<;bL/e^WHN1^DIN3cLL<Gg#ADaOKWd[4@
<bD&L[I62HB<\6-eD4M).a/_//M,1;E+.58=c7N?W]-NU=?@f4G_Xg4b\BaS,;P0
^.MVS\1Y3?.^d.7+\4R9NOd:\eP7.=-2NRAXL(a4H?];VL\ZJJb_^BXO>AVH)IIX
QIC:A0WP?g,=RLbc]@dF39&#6A.-/+26fML/@6G,ZA1g35H7N1H;+IYORgWGD7U?
AO[05;Ef+^gg50[<bG[RLCP^AV,bXge\@aUQ0\dS@UVc4C\].2U>ZRTDH]P781>b
50XVf1cD;<ccXS(Z\7E-P0:/4T:H#AQ?O1_>e9YSc.?RR0ZB6(09IU;OY6?c[]C7
Y5Z7Lg1RaR6YNXaa[9+O,=dS4IB1R2Z9:QG+HEMXF=T[b8fY.&a+J^KJ7)9\[_Z-
D1efb3E8TG(F93U&Ia-GL^33ATG5TXVKOeR@EA8Da0T8,9DL<@1eL+2PfC]aW6H2
Y(4cU42>3g#\/IaZ_U)_E_7PM3+A,cN^F.+PPRe<TQE\NMVK#91HBC9T^&b^^/b0
aWS@IR(1X)6]+#d_\4-H7C14M\.,T9ZIGA>cBLOOa?0#-=?J>K^RGY4Cf-:3HC&T
-364;RN:BGURa9?6M8O6N9Af17Q8^,,a0;U7]817Z?SG61QN=<VE=d51EfQ>=?MX
FU1;GHSe3XPa>HAWDDg&cDIB,G42+4R+F/;A5YMYb_V,\G,59a^8_+-d-\fI5Y<d
?O?KX:EfAHbeXe(9PK@OMZ-aH)Z,=[;a\+,f^MTaW++J&LG(H\0gDNQP5-IIR/XY
gQb]+ZbZDZNBD[GQ1JeXZER8(SK57NN^cG=eg5#=CUU.dF:D03R&9)98&^Ta60&=
;LE,D_:(O@MGJ^.TXK9eeRLC;S8TJ(_I]X7+0>R)gC)d#J7D2;U5LWIT@[;PG?;>
<(2W(SJCOALM]MDMHPG3MYCENZ_WX<R([>9NcG9FOKfE;d\bK?<2PgE1,NKY32W(
+91C74E<Y1HEO]a2IDC/W5.Z)5S&NU9JI0_^SJOeV1+7XRMf\U]4WNWJ).W.X)JK
.>A=P)0Q_]9=Abe_YS2adZD,P4V/S.@PYU8bOBE6Y2J_aI@<]PRd/SKR,.[VP\2N
>;IAY:AWI,8;L/]S#[OKc^cbV.IN_?g039<#UT>9Mg\e=CecJV3CL0+f1+UPPRcN
0=9\BIY\(/NO13U8LX7WA\ODWE_1dLa+aQQb5QN,f]7VYMIG)2R>YXKP]F8D0V\>
6F.>C(PY#N^ccNd?X+/DN):@7)38);(0&?5D/;SP6P/#[0M1SYL@#V6N3)PA:B[)
;e;f+LI67([CVJ\N77K)[Ie.Fe8<._7\dS<76_/7PX;DUf/UOV?8@WX+SB2VGd&5
F9cgZ.ee,(O=\EKH\1I.YF]>g\+R&UEc7Gf1+<,<BJDT-:0a]R>;aQeR-3#\T:KX
4N=?=W+[e?Rb=UU#g4dBXe;:263VX;7Yf@d@SL:VW0Eg8bQ,#7ESIaeegJ.HP]d.
T5&ENbee,]f:\1(6CdaPHMJSa#I(FC/+N3ZAEbe2BF,IXPCSKDFEV/\NbF7Vb9<N
g5;F].8<];<Z?;<FAe):B-&?0TD;B.QSNCAgd]1XXfLYY1[5FWHBJg>_I27^V?Rf
5)IR&gQ3H65b8HHU@SDA?UUP@aTF0b]+BT(AUYeGWA;#W/P78CGP:.[KJ4HFG]Bc
+dXS_;&PLW9J#AO;)B[PH1S)Y^7U#[JMJ;M#K)_2[\W2J_NVeRA)a8)8;H,>J4_L
M_3TL(4#@D^=V&D6W^2-0bS@4SHF-=6GT>I1;gS:NBKJHEScTJ]8VS>[0I\CKcKR
-.?/_CV7T3#T-_T-/WE-ID?>A.D/K>^6DJ,67fK:>Z]2:B_N-&15_:I56DH:L.f3
<W8LOQ?YBE1.,/a828PZ]=4>F<d<0;MSgNDB=T-.EV\._B>Pf;7?cU<GU:&Y(GDO
W@2-@X]2IOV,ZYgf3>R8DU)DHSI>S_UWC.I>US)94R3ZD?[1DE7(EFc76Qg]-Kf1
/2?#[\]FcAC=<H7M=b6997bc<H;)B-#U7aLXD4Qa\\#8;LD8aN0/4T15G5PQ2A5+
I+3H(+YQgA\8dW+G6dd_1f44C#F.7SJEBN_YXC?Q3+6cP@Z:f#>7e(DT5L2V;=2<
A=(Q0WG(FO\7-/Ud0Z2]7dR=U:HEDU62PVd4KDQPe@IC7K;=+KUAf]RSDJ\9Q6<M
@9dWf=JN]XQH_URB.-TE/bY=][T6:,4Y8D3B]@Ya,N&KCO]+DZZUY0XA7UdJG<9F
>Wag2<1P4<1]V-A:5PF[[H^H[4ga@c+b>c1I<d^Kb0Cag#5[J\#f1e#1a?d\><IM
\Q=F1(6[QaNIO?ADCT2eIQ?M>GEDNQ<<3BagN,>#X&1]O/#P.?5A++#Y-bG3KcSE
.5:ZTENG02##6#TS)]^#-D-[Kb0c;A2V1PEW2,:_8]:Q^^/g,\KV5WJb0J;F@&;N
4[6#I.C_c[G=MdP>.+.OYRP\+c2B?H^2KM-cJf7/F56DP<#CCVWSa/J-/cNbfU<X
PS9FQS9++c.dL-L=2-(a6B\[49:FP0O;/0+[&4,FRcB2e.<fFRM^@3H6Md&Z6f]\
Ja0,gV^:&g]VLR11/X18D6<.7A,]P^KceJT[POL4a=I9.5-2MGbAL#2eSJ^L\I/Y
TM]aFA).A6f:a]21(0MW0RS/:79-d&>(FDLGW#:U.297NO8WX>W]&PM:>:7U1H@5
4=B6f_>?(XQ+^J#aZWWf[d6b8^]OZ6V8a7RbOEM26YPMK\O6QXV>=R#5Z.TG]<1/
E,NU@0<U0b7TPM+d9OLQ/3<GVGEULFX#<Xd7:4@)\g&b&IW/L+g3J<ERWF-L971g
,,=?)(DAadM]>6a^7F>LVML;FdV\0BFOE\S_89O1&JDa3<ACbXMH>WHH&806J8E<
Xa\7<8dP^fQI#)SXAT/P^27=L#029XVVaFHM(?QIKOI_U,GX@QPY)17FOgK+d[V@
G)MU7@.7GCFG3?\3#/JdT-Q3+;_]a&D4R/H6K\5H:H#>5,=A(A4POfe6#JDSGK/f
e>5\L>OG&SXQ41M-RC[.Ne>d.AaFg5BR^?8U014W<TO9J7UHeKA=.)PMEL+dF7Fb
=^?7=/c]6R?=:^PYH71^W1aSXFJ[)O&0F9]9O?#bWO?4TaM+9(D271ANCN^dHBM6
R?fY8AUZG[X;JN2(\,JGM0<f32><ZV3L262(-f)4.QeTa)N=0RTH=Z[+A,>G:S9/
5Acd>IE4IBc&;1Q_#.JFMd5)TNa.UO.99>79IX+Z2RCXJaEacabWXEA,9Q@E<0ge
WYVTE3IRgY6#:(bMY;#F)M0gW?YLF/Q#)_)M&20b67-KTAJYTY.IK>]IRMPOO:>J
EV95GTaTc1e3+ADLYM1JL_1^<+5HHP9^:INV-TC7c-_gNH-:dbH:3N_FI28P>7Q_
2RYeg1a6B&ZGAeYW[[DV8/E2E?ScB^B]+LDIb8RF8c=g8Y&gAK>6YD7#(JdKT6E(
,.+fKbIH+A(GE]Q78U+WJQcBPZI.8W6:I(D?3b#Je&V>TQc.6BC.KcPg4)F3d[Sg
AOcE5,>/S?)PBE6fZ4N@e-d^dbIR#gKe<#XN5K/IV/\3KcF;(cF08A)[4I(\SMZ=
6R98.V+Q/7E(EY54ZF_O11)=4,)B1U;#_UM0B:0b-?,Y&\YJ2:1DaPfEP^Cafd8[
)0-aQ.SM:C\RYPaO[6_N5EFP^6(/+):H4+,f\<7DYKZP+JV])Jd9Jg<=g=AT#,AW
SMc\JR;aeO:5(HGVg(]KZ[;)X,KLG=??\(;G)/7L+ffVLRfES-Vg?eN5g:C-OF&R
?^UK+_K,@0AgcO:VdW\X--Ne81?9X\CQ[>Td2<gbb4eaM_@-J@;_EH9&Y1e.3C(#
S-BR/.R<L<U2C&?_/[eQL_6b#d]DHR>17=U+V#&]?#:7X1?H3M[6_F4VI0^-MV@M
F46JM:ZcbAT8]U-A[\F2([8IW:O_L?Ia:[IIG:bG+]MeEZI^LEV-U/J07:-LC7NA
.K]dNJ,UdJUJWDT@#f4[M.eF:B[48/__+\@gV+-5&HMAcZ_NW0=_We//KGAGg3VN
8FLRec.6f+1<4C63I3f->?-66(;@^VC1T\[dMP(WX_DU=d3@DdM4d6OdF(a&#X7Q
-9(O[d^7Cfc9MdKC50\-A/)9QQ7-cB\.URTd:5L#O@:OKS1TGM2,Z/QZ-TKeW)>T
,XXZLU2^<+JRBJ+N[HY\e.g8Xg7Z,#Z7]RA+aKPB6[E=FQDI6e>9FFV##1_b]FZ9
@)6.fG3e@^>,:9?-HX5OX0,8RQ;2:F6<;d(aORK#3^6GaHb-Td_AcB(L6:Og,&V.
X97cf6d3FML^IfO)H4#0F1Zc]DeY_,ML/TO(^/=ABbC)V#a\PWV?C@SccORR5TZ_
Xe;TWPBMc4@QUMRC19D]=2<Nc6UF.[X908>)09fD\<=&H[5,]Z_b&e>^?4QCSEC]
VQ;,RD&O7HRU@Ma+YEJ+@R_-I[a(bU_<1R\WEdZ9_LS7CKQD;DaC=+.:059@B19)
C\]7F4,0F?e1]CL)gN-&1SHF[_0RVUIg;f\0+BNfIb\U6>W?)T7@1Yf<;Q4)_=0N
LO;V_]0P8:1R2DIb-0@0LNf\-M6aRK.Z=./](7<3Qc,dHV<>6(Sb[9X11QC@@FV.
<HRJJI)K:>c4?U/ULRV)gI^.E..+/=@)K=/3Q+e_0(#8JP+#_PVN3JW+Ud\Fc^35
5(NRK9d\P&,b]/]PKR<3SP5WIW5Mg362L,&F75C(XY:/f<dE>aKFX5()>SXfe3A3
de8@R\cfg8L4<RTfaWg9e[(2^Q#Bd_.J1B:+Z<\RZAV0dT)[^^:gP0/-IT]-[(A=
RYXYVcaHIWH.[.RLS8b7S9)+PLD#TNX@L&F@[f8NP\IV;e3?I/AY_/68]e@EgNB_
AGV]_[P^D-Cg2[RTgFdDX(Vd1(SX36/Z>(XMBFE=\eL?R<1ZcDg(7TN[(>/>P/FJ
T7(_fd2K9/AAXb7M^c2_FYZ43XH/.gE9E+5RDf@HI27eDKW:N5]?5)N30]DP4IX(
f2_]?,S<\8D@D484FWH091;OIEHF1Q)2+C^a3ZH,85VU.TX,336ZJe#0B[SbLLO#
g]D9.8X3bYW,aT3Y?Q7V?80F(I&6]PY\ZIOW.#@GeLV(4^<4T;09+eJ2fSRH?0OK
V)-Z@P(V6+/TaV&bBH6Me#GBa5LL3JB/IB<aO_6<VZ46<P<e@K7B5Z]KS.gS5d40
IF893Ve;<,DPTFU)7/M4)2)UB)b\e1BP?_OIMXY;_CIV.4>G9[Ka4e_&g,@F#N/(
<RD8_Z._:KcAffUR8JW[2L.P8O.)?WE;O_5eF)G7UbGA&4eH4<_JAH.._J>YZbNe
\YF;5?cC;:1ZBJOP:[Xd6CH2X_<KT_I9c3_D_Ng]_=&C&f72QN1BIV<B9EENc5@@
GEDETd(@UT7FSUJPX:,E@6>.a:f1@)(AO6Y&b[dCd/b/RJP@QW<TI_C:63PM)2@[
EV6(BS4;I.#[,1A[[d):HPa=Z@E4MK]MF>Q8V(TfYIXU)FIWBR:802FT+I>)@UX&
G[JTA?;#BZ5?N/,XBLOAD+&N;/X4&4F?VQ&Ec[_^+33RB7:FP+K2P3;;K&9LUWE,
9J4c.>&g:@G/N]Q_6(ZF)MT/,+Yc#],;7:6R))LI4UUJ[(Q,AG5MGLNN=JYb#R^=
TYGC(7A]#))=+XcFa]C.19<H,f?\3R4/IX_HE5a+PW=:d@)W/7d[.ST@La9<<9d;
-\Y5e_6]K.89>;MC0<6,8dCQCCX4fO)=U3_+8OJ-<NGJd1K8cdN&>)S1.9I)J\24
[7T.>CCC,+_\N4)KQdTK;SNg4OE:c8?@IG<+H8^Y-L)JEa)@Jd=Pa4J0e]48YCO/
3>9T>O@4d8ERI0-cdP9\Y9HbH]4)#6C[N97PMMQdb1?EF</)S,g2?e[Ba0HD2<V;
5e\WgEa?UU80YMP?>N@LN^Wcd[;JWaDJ]cX+F-&0Y:gOG8IIffdZ<#2b\#]MaBR1
NUX#QZ13gRWF3)PD<R@3V9R_()g4b87J\?L4^DI]U><bg=_cKG8A?8;9bNHHFfUc
H?+O08D?B@K?X[[AKWYEeBFI&WgC6JC>X73>d/a0GSFY;2Hd5;]\H2/+XD]bb:[S
@+VGC/JW-2#A^7g3O#;2BUFg9KK^fJIN)QM2J:_f1ST@]_TJ\#BF(HWPYB>MK2V?
;bVK+V\1cH?3Q6-VR)BCW65+0Q].X>f1)P5G^1D0DGf+c&HKabMDPN[e;YO<HHNM
<]I<\6a./5[ZWC=@80OS&#,DU#R46FQ(8/W_d8\Q7NZA_3GLM_&XV01;GB3+MS6E
32[f/DdMAdTEAgN/G@PN)SA(@(P(8XLfbKCF8ZJ_#gKHZE]V]3YO0de/8g#ECKR:
)?c9d=W63-J+CaF296CgW?(:+I;^4H/:-G,aISaa6XIXF^dPR6<Y#7^A,>X3+gY/
[:[^]><M4_A8HgW[N6\[+b]1\3DF5P74W\?Z2e89b>7ZCT9^E(FfdZ70gO9>@d@X
+=F-^FWQb>44cCMKT(558>SLXQPdBBK>[+I]U^)/(78eA+-=3C)R0V5P>)XLBDWe
_YU/L42?((6V1770/>Qf9NL?QV),.CPV2;A@cY374\[ASb9P,4T2=^E]1+\_3/FY
a;=<bd<dQe32Q=<D2^A,E&PCA^Q8#SgQ</_;QYRQ,>Qd6^Y&ZLO^WXGQ/.f-L[>]
:Df#BbNUg1S00T/JM_f;HI3<X40T]=6Pe&H\]3>dNFHG@AY#>gVY+a/@GX>F/-TW
7OI,309f<eIgEL[9,bYP,,S8MY66TL>1+T,Q.<?#FSMSIQe.RRN+S-Z_McXTLa9Z
6-@+E8SS:)\1:b(ZRb+d(C89V1V]JY/>HK^.AUNPdUU@&=+eRAWUb=C-)[cc)GVa
1NdLH=B4MW+37ef\+bV0RZV:aUT12gc(IBB1F_\S9dc2+#2cTY8b:;PB-B73b4A2
)1PKLd9=LQ_,E-4/@c:RZE\?9[;V+^=\-7U->bX&/;AYe+41C8&H/;f33eVM/RX@
?+KZX4?I:aWL[a.GS\\Kf@P0_D0A()3OGCf6<X7Uda?A=bc@Ye^L.N<Qb[J&S&Yb
P)\;=b\[M@PQ?&^XZQ3/NIbE]5ORgS26c:F/H;d057LVgbaRQL5Wd&X<=dXVNIX9
3OH;/OTHGUaXb3]&)^-6e2/Rc,)1Qa+,0<??F34M8f,9J>[]<R>EUK)]9:A=DI1P
2)G:HP1S#g;H@HT7RPP_<>eBbcedV2;/g/P,.Z1H8@/W]N=]OUcINd7->(,J+,#N
@,&#UC/_L^c/Pc?1/^_:4@QLKeZ/PM/L84aJLO_]5-[a45SBA&8M?XGQf86O5,MS
DN#\.?\:B<?G4f46\/5[./>>BH;<E8<7&5bW_5E1e5J+OBX50H_-F<RL0=]fbF1R
]Va>+bS^\;f0UD2EMfRHANG:&W>+/7[GJ=De@I[KSMgR47^]U.;(fUA\#6aWNR?7
-4PK=E&:VaX\_Y,/HX?0FNVK>8BI)]gGWOL[]S=]9?T),RQG#0a07/8c>Z==4L7?
>99,L;2g_)E4>YgO/&Gfef552S+KG@;a,G@b]1_XS>XKN_5bGSPDF7>RKd&X^M))
/G5F\.FWLI;O9I1,fb05F#>7^Y2=L=>V&VC@-AHL.eUQdTOQ80)PK]P[9H^[24L>
0b@P10(=<6K@FO(G6D;VUKcJB@QdR4f<#@QQ-@1bBT)a#6V7/(4@/]aHGF7#W+AN
9[X?#.]/LBV>T6_)YgWe3ECH>ReH9-gN>SZKL^2(LFa<&WME5^C-_(.BW9C4CV8(
2F14Q-V-V_\CcRUL<G?0DO?-,^IIUdYZ#E5=50cE.^73[e6XR5D/JR&]\3d=e4=P
-3f[@=Z9#WZ&THcOD1cc@d6Y=df^?Ic6e&^1F6_DV/4VL&M5,[RMBDC7;3T1g3L(
W3eLbdf>4^QbdQ0[0)#NEFJ=M0PXXNc#,^X;M^GUDQMW7J(eJ2A+_(c3Vg?I)RAA
U5FB.>a1\NROD#AUH0Tc@A33EId9KZ<H;@97/5UI&E;&A8)cSZQD8b/FXXVG^DH_
R36(UMA)8;PHR)Y>FUd\C_#&6N7442U<TgY?0?e8WA]RgBDgCaZcVCC(=RLM&US-
LDb082@O,eIXO0OP>GAVV5QT?e(7A,1-?WeDgO(,Q<B7-DRL8CN[=4X8/KVeUa&W
6]a]PeM(JefAQZZ1H7(I7=LZaNT4:7B]OUTA+eIgQ]_Gg((6YFcJ_4[U0dM_fBEJ
S-c#gF7[SG/f5dT]>_aXFa4Y5L:_@T&-ZAV#c]^XgFV_S;^ND2<eVTH/<;MYT)\0
<XaHDTEeA=7X1A[]XJA1f\KSJ99B89&_AOL+52A/#U?c:^E#09-N,f.7<+/8@>?d
FJK-CRV9?-?5FG#OM2Sb)9-:LTFSAU1P,c[Q_:70(GQZ;[Jf@,I?b?g1<THaK&?H
BeRZ&6,^UeR7R,2K3:R)OAOb>WD.KBR^,]]S>PUTa)8IBb/acKRa33PAMYK6496U
&Z:>(5:F>G2+QA6W>93H==<1gBeCgSQX).4G]>K,Je_F0UNfS>Wc>#>bdcKXVZeG
J\2:D:<ba1R,D-6a.aIG#W7+1_#d(X)bdLaHU_NTYB0CYb;d><:gb/CXPR4EUXY)
J1+71F6J-HSU9=XdDc;gKR:#@aT.IF;WUI6;XM)NIF[cdGbT61^?)K=[L5Jg]L74
C/24(ZEOQ\R8d6B2^\;ZC,+RVY;([BZcS^-VafCNW3e9dc):RB))>H@b5e75PdL2
LQGO+gA2dD1?[Ob@QEC]AF+G2XRf.QW8SHO&PH?&U20W+G03(<(+51?XMP/7-N<f
&CLDG&Dde_Kc@F26]#09_PC_4TPA=?OG;UBD\8Ld-+S&SI:,@K\],G\3[77Y@B<6
7f5^:/fIBN2?,[;@b.D8V+Tg+H=ed9+C=[e&;@U)NJ@E0DE8.L;D>a=g?a/ZV8,F
VW?,E=\EbS1MCLO<.c]OSO8FDc@D]OEe\+4-C:.[K4=#;WdX_IPM+L0HaLg.-YP/
F9UYe0,?0W,6MJ+XA[F6@25Db-G7\CR=\R9>g34DE&&g-d(L)?5X)C+&gLb@eA)V
@M)V2LMY1;RQI^/^7ULTc_IF;@C47fbC/cG&HTXB/H@bEY1;Tcc:g.,22Pac9DQ[
5=)=1C4G:JY2feQ)@A>CYL^L4D?F4S(E(6>0CeG><K0BYKM&-E/Cg?;#23@X3A/b
ae0_6>ge)>3a@U2659PM-b+DdNBY-NR?[SL37Y?8LA5,SdG=Dg(A)AC]6@^:WR-B
2UT9-6)LKb,YF;b4^;/8S&2(?IT4f<E/A3Q11S]^<,<SP^3FZ;>1)9M3KSJC8J)A
cFOCAdd&7U,Q2fTF+C?8&\AX,01SHc?/HHa>SB698d#UPB\7SL^V9[XSJJ,N+00[
?:YSPB+T;YABCfNVHN(#38RC)VgbJYSWZGU_17aS&16+S2.#G_I,]&fJWge;X#:e
1#UCMaWDJ[)7]J9eL&R=2X,Yb\AKI>Tc-c&O^DT&TJJ.LUMT\6H:V:Q7_W=Me&6C
:T0V.-;OH5K<NHQ+EHJ?PFCTS.9Z9KY-;a?XRL-TO;gYC2cDg8Aag/1/#_YBQH87
dfN17e&]GgP+RL.+\OHH<Eg_+<@V9-^-,-^F371;Y7d0-1>AQa+:PQPXa^F<TEKL
H.38@:?HCMUXaJ6d]H\1PFUI[<33b(??ca(c?N]BaH(>2J\W.8abU+30\:\Zg<_T
FLZ>L2F#TGc05+be-F#?[\e9GdM)2+GE320V5+-UY/E8Ecb5N(0MJdJ\4aZUKY+f
I]XX,16)=<LUAaFPN2<OT51S2XLNeAP=K-#@OQge4O-Uf<fM?bK)-3C_.aD>TR5B
[Cg0A\QETE+=QGC^OE6W\5(UNFFDbNTR67PVI5#U4M0N6/X0-30#+HOVF&f2<XA7
@Pc4J4RU0(=Ked;ZW:64?YSH1)Te<[\00+EFd0M/\LZP5Y7KM1:7W<MMN.L?&ZT/
^S(KCMFZN]>1D/Y>K=J-];/9UeOd3M8f?;KMX2Hd>fO8_Y1gKR>G)5P2=G(R[KQ0
AQfNbG>=S(BCc\M-[T3[9+S\R=MbS,+LQ0QG@KGP:GdT84Z,X/OE\(##fG+G.B(b
1^&QAJ6e/BI&@&D.c]VS;(O:g)O)\gCSS(3aa9Q/8?=f#7Ig56(Z4GUbaIXNO])Q
U_NBLA4&U/-WV#cH-)JK_>PICA2Vf=,;:-f+g8HJ82C:RYQA<1(VXf:;BYb2aO6F
3F.2g5>U_X[J?YSaM/ZTB+>;S5dB]UPG=+ZRR(HV7P=_gD3?c=;WdO-:+,7C+#5-
c0N>A8Q:7F@0Zf)918M,[GbPRc?&T>=90B\YICM.=/4+Vf(._AAUM@RD3VdX7;ff
C=W=W.#51;PfF7(6SOEJ_c9&GHYG8@)@2ffWDbdO#J2R:(P1@6KY2TdeB7K7H90V
?bO+_2-YXFg(Q/:eY0A9<]IYROG99^IMSDMUE].R7M/&@B62X;^,V3L_Y_X;a/GI
EELHD3cGQN]JXIXaQecFO/3G((+XTD7H2_+]6b5<d04D]GJI87d\&^_479gN>5=c
4R(,/X00LJd[.(8Z/_I;NZ8)&Ta4fFDB@d?0@)QXDa8GPd,)44PYd88]IKXHg#WC
gUDZN(I8::GLG,4)-BBM/(?L@XZQP4c6N90J.Td90XYB:6M:C,CE+:(OSUAWQ(e6
DD_DI&0]F7F8K-;;bG.>#fHFf/fN_&JZ4fM#MISW^+[=fGYbS1/1.0/]7WY_>E.G
P(bI1#fNe&\L<#2JMF[?J\2\.YEd3d\3bNTc\9(>]]4/bZZ,14VPCQ[5(63e-@2[
Aa-9?LfB#S6=<<].c?(fgb)CJ:WNc(Q.)>._9OaNDB?GfO)#.M8V6dK1C<^d)a_F
&)^E\Le33&RNF2Wc_3eV\JCP8c6g3IV:D770Q19]aV+YD?]UO=AW=E=?a_K_)?.\
^e@VcK\.b8e5Uc\ODS9,NTcE(T1:eC/X=Y+96P_c&<[e(X8QGMQ__ebK1CY&egV]
RCQc]9.A/+\ZJ&f\[DfM7;[6R)bAXfgRO#@S+5=]5]@J2Q9b[/-9+5MC?NGL/I;V
1UZQ30gKf&F.Kg;Hbde&43=>7A:D?(VG1=00/5W5;-Q#c\-K8Z\6Dd-=AR>C_[^>
VH&8Ea&[&SKH;R(+]<2X9L6V2Ff+DbQE1>UJ<5Y<7M=BR+R#J5c0&ILCefM9/AG?
BAI4^G&3A=(VS:ZETN9gZe8bW,+-TP2(RVZgg7eF=0?OW<GJA&+RP@]f_AAEa5OC
>U96Yc1?,BZaR&LaK+87&AO9Z_:cC>c;8af/4ZKZZ&b3\fRBeNdab:gRd7eaDe)N
I9C-4E<e:4f[3&WdG:397GU,+4&M-#)?&>:gD;(fYR)@4;Ha0@K/\<(VS7Z/DdAR
;&CV0M3S7GW:MUbUS]^g-=0U-U0d8cNg948W[(I^V5(]L+J#T[UUBXQNLP3#g(@/
^gT#;C<8@/T2YWQ]1AF&QXH//FZ_(OUK_T@<FFHCfJD:@\OVaJg[IWGcfQIea31]
<Hf6F2G(>K5DFcQ1@8N_=D:I[ID5S[a&@bW=A\IXOJHYAGeObO&9M)>^PAB3dGV=
VfBS21?X74N>S_LYP[IcB@^.JVPf./B;_20?=\P:c=EAA7H_cI8<3>K2c[-VefcA
[IW_1f_4D=[X-L5_<ROOMC&DTNN@Ya>D<;95+^LNG3MI4JZNW#>;8AeD>(4&R)+?
TABd>,5d<ESVD2A\LS2793:.E9Q&&VQ-;_4cN\&SPSVCFP[>(b]T\0&9/Oa=eKU)
>FWN(AV^2(6_GC>_HIM.F4._b>B4c^9e,F[7_f_Q94RP:ZXAI8WBH4,3d6>4N<O=
V2(VV8K#M5,GB#-Z3&Y(<XacX4&7[8=Y#;a43b[N_:.8^#8^]IgH-ZM1>W;R0aAK
)A<8<,K)aZA\W_Q,<7N>Uc]Wc?/@71@F.<D1)2B+0Rgf\-/@d,V<CQH-:QTJ,=^b
U?K55X97<LWUU#+\T7P\?M3.;9@e75_eLW[&F9Q>Q-ac4ebZXbG5O32>+98c<II+
<..3.0H59ee_e:BR5V=G1W_JgTQF;9B@49bY7_/)K4JG@<;SSTBeA:3N#E2<)9_L
P<2L(XPDDF6<d]@cfVRH3\_3d\IdD4=\Z@_Ra&+;cR[cQ#EA8UM6F57Q4(ZfT5Z6
V8EH^d4=1&@.Y+7(5K]8<H8Y@0XB6a>SP5Z5C6R=0f,a2,7CN)Q/b8UUSB@X-;64
Z4E_Q1S5K,&_>=REcN^:48fK/?^[23PU)6)H^>+;)_\dYDGOFVcV;Y<RO=17A_&L
,(1fG>0S_E-<XaFe.<(MVDXA_Tg3\8/))M0A]KeF##37]U2#LONBNE>^LH)SDf_)
7C1B;+G;P3QCE2fU0-C),&a(3YGEQ6gN4\EFF2/H.eS\=H5TZ8fg-LC@W7b5a]7Y
4YT@7#)aL_9MET#^>T2B-IGgf_Uab39P:<N<C.Z5Q3VD1K#/DD;,Ed6W?)#06Zg=
@g?MGE>d,<LJ^2UIg2SW=9Mc[5ZMX_8D]?P25Z5cI#HKKL:2#4AOe1N&4:aaMCHZ
EP37dJ[.(;0BYUbH1\M8]=a;g2[OYH=IL\?T]#cW?K/VHe8J>@_T?8UPf1;<EE;G
EJH]:0cf;_-2_?J_[2]VK^RLVE6W:;@dW1)0DH52I,Y0#J&B>;403C5T,2?9;TeD
QgK#H\DWA1.]19:@F]eO?AXc:Z_f>^[IAVH?4\5SG/T;J<J)Z<Tg/OBU<9SHOL:4
b0H,I;Rg,GgUMXMRJSWG8M6NDa<f&IVH05fC:390ZQ=5,:cN88(7,P,]5MW9&7[;
/.MNJM0ZYE>/,&@EY;?(R8dM#8K7ZH2--?(]f80>GF?aCd+IS#f^4Z5[-gO-HW\J
\#OC:VM03>&[,IRMN(BbUA<VF)+:MYNP-Y2K\UaJ)fEFa&UBb/<W/TJM:0R@DR/)
bQ<(HeH8DV.EWXPa_AJM:Rde@G-&]Xb#-3F:SNeD7X+U(6IN4^0J@S[B.\f\c.5A
W=95I+;GQc7)Vf)S1(CWJ9H>HIX4cSA,R8;L5C]Ef0/5\#<8IWD^Z[JJ-Q&/];U9
,V1?I#C/880eVMV(69Wb>Bb[7gX](@4)\1.,D29VZUcGHO/HE#Ag1E&-HZ3N(Jdb
DDYACY/_NLcLDJb:9Q?FK+6I3K=<1J=(;Ndec,LP&/]M7d?eMAOcXbLV//?H-e7T
bP0O#(UVKEJ]JHQ(Mc\^OGSN4X5,Y6>>b)RJA\;#S/\e63D1ND.1PUD7:OJ8Q:K#
T@d8V\E_.A42<R+a8fJ_SHd?Q]=E#a0KWV&B-#WKRS<Q+Hg@g0:-?[d0+I:F9(->
0fCHGB\/6W[]^Q].TI&4JF_E\S[7U61CI_88bf2T+3NXV,1dfa_Z)EaR#VO&PbH7
DbTYO2bN)9;^4I)Of#OXHfV4;=eTW7K]:^=dO(5_Y0SA2gOLCP,Q@UM]O[W+)#dD
OP6(_gNB?6YQ#c>gZEY,N=?#9)d>3c?-06K5HSMb>aHH/L=QLVVRSI+M(]L5&)HH
(6MV5^dRP8QgQJR+JU1[:G.80#cbPbB;7C=.I9)K/-e]MC(BaJ<\JD0.^W1GUU;/
<-^M/0SH2&LHC;W,HW[^9EN(0ICOc2d\-deRKcOP+cB)(#@U-_KBW<I\Q,9+3NVC
6f98&W<a7:[E&;D0GG9gI83LNNZc+_2Y_fL[+1;FH8=+;\#,c^TQ8[TK&d;TP>>-
_KfW)WIU9GRZ]HcX+E:HE?C.#,D?T6c&=A=SQ:a<ZMR60bT89SFL3S]QT?\LcXN5
ZKI:KO0;XL]Cd55IZcT9;]JAEG3bK9?NUfUYLQWIO<]X+WJ>g_6g0ULHS-0DLO(_
LT(5[NaQ_A.;\LH;&=;T6OPR.AEVIVEfB@(eJ<7O]:dg6#E2L]>?[UeS&_FP1TNZ
V(SW#)_K+E(U&942+:e)K7Y+RHBD7D#D:=US(JRC,IWR8<Y7P.aGf3Q,-@..8-E7
Zf4d++FI]Q\((/f[^H6T]bV)&(f<6fd-JcD1Q,7+5+[@=/3e+6O5^?B=,Z]GKK-V
_?Tf5)fX/cb:33e)@W&T2DAS1c<>Y,TDKcY;)e;cN-OaT]70/.:6_M@9PFaPGYU^
>2@=OU1>UL&O@EQB]9KF,F)V1a9AbM])X:eNH>3]/@A_4&;@LS21-\dM6WCC7,AY
D5#L<D<EYNIgGPBWd=^E8UREHfF)=W/4\O_&eE,\&MJGJ?KZK?6:b<M?.dYb\I1=
>4)GAF#fHAP3A:TgR1J+F+6dWcR:J3+?RXg@KV3V85X,]:8I<IJTZJZ;b)[]6^4b
6Na?b/g;ca.e,ETP6GLO@8GQ0O5ZMd\/GNK_2<@W5EV=<N3?_=dQ.+;fF;9#)GZ^
eX7BQd:0(K+<)GC<:d_=#Jd>L2SLIaeR)#&K[0O>8?V4VD[R&KC6K^e(T0?=/MFE
_?cWRWK[/2:Z[^Ecg@2L9Kf=fM&N.P>M8XN(L_>SC)#gL>:AD6C/JN5OJb_-Vf@=
>ReC2/cg>/1GUWQG5c5Y[.0V&GL.bN.[A1@VM:#V0cF5>e5))W7fAB\7]a:@O]PL
J/+TJHd]SWF5U3,eKggQdE815#5<)/T>51JIA&P)@H0W^XN,aB1NL=_N&_cFXEZC
4=?MeN;-TfVSb2BegLP:)1LK7_Z9^KU4AFS.UC,OY9E(Z3aUI4LJEfG^;=>U?U>K
S?4fACF=.?fK..DJaCA1=ZZ--W5&SgD=OX+/0Z(M_=bN/Lg\H741(e#8/W9?V]#0
RP65JSP32Z7\H&J?[2)0>9DecZ(]A-\B-HBEGP[RJ&A#5@b;)>3\X(E@gREKC6RO
6AcTZ4_HEY6<g#/=8Y5<QZO[Q:U6>LO;:YRO)N2+LG4Wa][W5Y#eRTeZUg7,?19a
^2^=]G?>G8c7fZe2MBFfW]V9.d3gT9F[=D&@^0>TT\NUJ7NPE83(-3]AKVfQOW@>
c]JZK:=F3K20T#6_Aa@G#AEC6,+\P5:#D>-2(X50851RZ,?3AF2FPDY,<M+_CbCQ
>?B0GTAI[fI)d&F(6;VV7&S^[&BH=DV-<P>3Me<M,@LFMI1#<B2C+ZaG9##Y[2X]
#Vc[E8IOY91&9P4M6KL2ReJ3f0/\S5J<[gPI?YG;LJ3QAHKSGQ0]74.\N_UF2ELB
KMe1E(HCFV6,_7L?a6O4[8DW34,?RJ6dM9TgJC3KfHSd7D=)X0(KfIPa7^>Z2=a?
Wg14Q<_;L^ZTNEcWEeB.,bOV0,3c:>Y8,>.8T]W(H5YZ>,e[.W:b^CY#+4Wa8\e8
1N?#.K6BW-OT]F0)/D(O;>c4O,gP^/?P3_c(LLFFc]8I,PP>^ECdBA/4J]/(,]Zf
fU:)dS2[fGIWQ]=Q?5df_/_88ZIFg]<VU;O])g^J/]5QCW04dP#@+<dHeMFXE8^F
\>0TQW;H;U+HA\:9\?QW#Q&3Y2V]<Q3)ZDHf:7-3Q6/YReML291HGGdFR4ZK=aCN
a[V)61C9DL1d2T3)bcA^DHNEFZf-N4EV0P_eTPDM^g+1<c(.M5E[;)85a1Me0/4,
d5>;C9ZB1/-_X-d_Ne#D_X(DIg5+E:S4HAAS?e8eMgB@IK,\AA;[F[KQR[b?MgS_
WDG=20:?BgINGYVB3N;XCFYPX-6)]ABQ#]0A38>_N^>-+5C36(KV,N9GHU1e\b1O
W<_f@W]d#GK9;N\?0<aD-7YXURXN]LIbLN-g1J&ePa2+/+S;ST\/f5Z7+<gbC+=.
Cb164fIfIO[6O=)Db:<J,(LTKR])/+>?L\(.B=0fN+>F/G/6Ye:G?g?TG9Q6aJY7
R?J=,[.30:,.PcTY+T_S((@,7dY?fWPDF>OS;HeTZ>?GS3YQ?Ub\OU7Q,=UD?0.X
&aWY.;4c/JCVdcd4eO]gM;JGEgYJK2,J)b@/>]#+R#54Cg[Sg>^FV]1WEK>H@KT)
:fBE-?A^JHXB=aFa=5Q8bXU.QL6;F@?Z+,f7,O_1e+XV,c4Q;WNA6EQJYUN7L/UY
d\=+B7XB9FQ@_)_FU9WJQ.0?>Nf12XEE75=O;H_7-UM:A[/X4[Y>0Z+_bUGXII[I
RI4+8YeC\@XY09dd@S0IVf5Ia9?Z=5+bWI5T>DYQM7?P8-M_LL#+/XS<AJf_>4J]
CeLI#47HdV?cO,W(42b2G64Z80XOQ/)4L<4f\X9O]:8bK.Oa=D>Fdb25.)<GP8\Y
G03Z@3.]@J>W,:-Wc+[WG/1P2bW)(WMTGAgZ-D9=C8T2A66D=7_MEaWJ3GL9d)6K
aXf8e:.]KI#dU/9:PHg7CfQ0PIbASDTS3#>N7S2;ORIb\F1Ma[a4F;H:1.]46,U-
-#T+GL8(eF8bKF2[,RL6UfMJ;-9.G#@G8FLbI[Te[2)K4b?BSN5_Rb.>[C7,K\/W
3KL,PLe<2CZbZK03;+RgZ\cc\D6@EXS2RZ^,]RbTQ3GPQT[=?EOWN_A6O?SB-NGb
[3U0=dDbZe,TdPH&bOH2I?T#:/6c@X3a=><66W+PW-8;QSAbPKR3aP/XXS@DK)7^
eQO+N(dMJ#26Lc/DITBND_dQU&2?I:TPaI\_15SQF^5I9c/fV7f>Kd).CLCL<(@J
JFCY9XPRJfK6D:aD<_-51G7PL7/&#QgNS/T\+FB-.AXL4bee.T,HJMXZd:<1-+De
XG:aSL\L#F7T#FJ;bZ4e54#^S-C)N0Qd(,3J)L?G(4dNG#(#_J-88[COgR;>IGB8
Q6]2>27DPOFOA_PedF;+4TRYa#,E8.<>E;)0]8>H2+Og#A<+=-5_)Q2Gf13W+E.3
d_7Jc6#/78Z0fe/4Z4KfX)cQ4S+_Z\/0I<6X<[@0dfS0M,^#.C[B5F_G^CK;LWQg
70#DJ?cK@d@:A7^VfR,IJZ5RY>A&WdF2K\b4YML.E2((dB2-?_MD\?<)ESgAQ7(0
KAH4O065#C2fd6aG/gdL^01@-0<4X[+CZ3b.Tec#V_:6?+LV<]&[f&NZ@;2gG#3#
)G:(b_Tc#3Eda:DD=W-g#g56+EW\NcK=<f#_eWHK#XMaN#I:MLH9@F=#1SL8a5aP
gT<-V&,FJRa;K\LS.A(3I)Z?[aWWGVV^.cc3F3McCZU:)KD4/Oe\AKCGAKO]\\>1
DEOPAC=DH,74c#efTS<Z1M7M,+.Z[3LddVOGb-&+^)H7.;\7I<JK8RC^VT.J>228
B-GCMJ,+G(M\=>97BY/L=;G\)D60a64I?@3,TPYX,MaSON:g)_,eb.Ff&,8R#0Sa
XN6SJVPSMEC+.4P3]T1_9K]1Y=U]U1[3f.U&CeT<K//^GG9R=Idb8AQM&bS5T>>I
5e4O)@M(]eRSe]-;gCIQ#?/+SeFc8/87>C-O\M^[V5:&?-2D]@#f<1Bf^X\@[Ma/
VA<QaG@36Xe2GK),^VO6\e9c=RNeZSQYU)1[\\[46QH=_WJE7\)_[-M\P9Z6;fg.
>_<>8)]dOS0Q7<>2V)&OaQ8+,c0DU8A(\;eKaYB2R<VQ5MP;V=b4=-IX^?Va/.b^
C&(Z0I3.VR2XJc5-_\N-;YL3g?^02-RL)UCKD4H3Wga7U:]B:6RUJ+A(@D#O>B<C
:,;Uc.QXNbcKPS;D_cG=,37a^)3J=)gN3I0E+TTgHR38,DOPIA[T\IJF2/MAHXSg
6+e5=6[Q:ICBCDWMR:5XO0OB>MT+C#JZSbJ]CQ^N(1H\0F>TCDK#_Z5cILW&gXKF
<;R]UA?&ZJOUf-+g4<801)S.FN,((:D\^[5Q/B]PPD+)(c;FX2gg\Z@X//Pf8=]R
f7bg,JMZ.1W?c/Y5T9DWCS^+-b?ID&_0L_12N+ZD1&gG+JJ_].&)[c9^X;&C<bZ:
#H:G58d/(8Y<:@VRC_\#3>EaG:3\KffbY])A^X=>f:5-FX7(Y>J92K-O#RTJ<J@[
<R&4NNTGOL)gJ&IGR,98JVQ4H(O/&3cb^9GULdb>[&D[4:/;AD23:A+c>XK74d2<
CIP_SWBNYfRg1@PYGaG+^Hc/fMNX:<C9D>&=f\g)?f@U&g-)9/;eN8LQG6K\eb:T
#TR+1;.U7QZZWW;UHQ-V\=PW,e_E62ac_,<]STf/N0641Z@54TGd^cNSNC]J1HFP
gQ/N.EaGEV5gXQ9bbM1ca+PKf&<H(e5e-UTE;(0(f1^=#MAVBY5?f3O<^\G;9F\4
R.N7eBJ)dPaGLM5e=EV0+:J8aUc4<R?PRZY97:F_;YTf):1[^3<eD70FW(WA9S]#
<95TOX\9\8?W6W4,P#:#NSf>e[g(Af?-Td+KKDO.M^G]<P@H<EPH@Z/&\#g/b1SR
PQ5=T>0&-UWLC(I;@Wc(Wf;/YXMd<]2[J9,IRc?0?XE(=MI>g=6[d[<]=@ZSCT91
3\/P(=Tg9f9KR:^MgEW?WBNcRa=^;a[LaO[51@DPS@]XB]G:TJT//L4AEX\BZ6eY
:J5+g_7RF1.O:#U;#\MIEbbcUB2:gb;7Y:/SR<Q_SK5ITcD8VZge_)K<=gN7K(:B
:I7b>VR6(f[]c&^X;J\MOXH=TZU2>V]3DET.cKZZ&VKZ(OX-@>AAD+OQ.N47AeH/
HF]#.K4;#CUZ@8TaF0&f56YM:VRZ>-AbJBeNB<5O6#BW^AeORL#Oc4bFP8EO2<9e
,/K6G.RObGe25LEL]J<)JPBdVa(XK)/F>GLR[0KX)2IDc<RbO4[+WEa8._<L<KJ9
,V@S&&bSc942);43&4BH2b:H:\B:S.OX#JI09WS[?&_G:FRE+#2-OINI\Z4T1REO
DIQ8Q]>-c[#aN@>S5)0fD1BY@Y.:O?N1_=cL5/NS(_X]T:5@MVCHc\e>9/Vaeb<+
bJ(I2C[B:X,B)&QS\c);e6,@40dcHVO)U&_cEb8U2=YMV-8U4SY#HX?Kg)5@8TTX
CZ(ZOC.g=?31aUTKd^_A2[&J8#fC:,Fg[G>/&_N#2A]KD7#6))KUdaJDB_OU0V_0
OX(I;.&P;9\DLG)2B-9K]X:)?NT<Ng75e1B30RCbCJ9Xe7^PL[&>@Rb&.MMc]H#7
M5_UA.?VTAd\W/8,99\6I[D9R<?@6;aS1IbH&V=7-.PdX(&V>@aDA^W^M)N?\L>C
E,N[N=(30EaJKO4X2(K0c_=e=cNa:A<[_QIDY01QN8=e#+GN:7\8(48?MG6]X6[S
fC7?\,@e8F:Kb=&,A>/K8?Q:?,b=G7V,PEJ?\[6P)=I@T/Nf4+<AQ7]VXG8C#(PQ
4cC^XT/cOIU<ARcJD32YaB-EJO4H+.;()3,TF--F[766D9,E2M/\4__P=QQZI8/M
Q4fJZ#Ya?R9,XC08SP\78Z1dB4GR^62XdPRa.D=+4g#O3dC+X6INN@f4;YOAI:b1
>K]K/NI8HP8@6::ZY^]5bcA_LV#1STT8R4;#--U=c[5JMg47:009C81X0;V<H,(Y
,&M6.1b-#]ef\YgPED\XL0XRJZ,(OZ&@HEOX+?M)DOWQLX@_(Jc[TO<QR&03ESa1
NeZZ1QKNRW@NF?3<G^<T1E?N57WC]JH?UF4^L.EMbe.G=UJ(<d160X8\L-PP1P.&
0.dNCKeg76cb9f[14GAX1UC7DQ:b,Pc9AXacP(^Ia+\5A>6Tb,\ab;:9\W[HYe/Y
W,/UN#O2K\d98K_aeQcC2J4F^CNVESFCXVfC)Z8F/^-#1&F>,4TJ/<-&M6OLe,M<
G\JQ8b9[D)T7(;SP(V>[@TUMCUF#dZE\d200VU9)7OSZSUWQXYIWXX3F_NR71,_K
6ZO^I[,BZ6>L&1AN@Bb-.+1Y9[0],\OK[L5B8@#@76d&fLc\>ZXJ75ZY5<\OM=8D
bR^JId/=dIdWOI,8a&YJ:TY@D-.)O&\##&a.;&,D0M2a:(-d8@Oa(+a?2NGg>777
NU5_W6TMKIK7Ng4BCSV?ZP;ZbcSV(O#,?+^R66@P#3U^D\80&=)W\_K(#J8MDe..
cb2QS#>LP2T/]S&:)\5&?dOTeE6Bg.KF(W.\?KZAON9B]gR--bT#cCS;=BT,;b\>
OUN50F>5@/9EX8W^?.,75<K<Zd>@NOBRRd@d2\#PV3UFfV]C<\<]@N,?gKHB@>D(
7WR6eC+\:NCT>90?O4Bcb)\8b]&D-_03V8PVIZI32[E(C3L3JP78.0.^@F3?=1d9
A7gM)JaTLf,Y:4XN7JQV-]9ST&N/>g)=\7NM<Q(+RW@._C[XP8EaA.4P#_+6&^,/
Je-Hb_Y-APV<APC.M0TX=a+VdE,4=_6X[QDbT7.cGPI^V>EaDb(QE(5ZEAC#aB\V
=f3]17VG_a_8(#K[5E#+_<&/V-Y_FX&4+DZ;99X+gQCg]aYb^)OS,(1IPfZ2V\:3
;&,FC-X?aI;+_:H2D_/\#3-0B#-(=\Mf<P)Q)HV+ea+b>1Ud&a,b8=&aP3dMB\b+
8cYe;OJ=HcZS+Ng]:XH2VJ.WGVN7QR3HeFUZZSRMNA)]4RXB^\Kcf4Lc32L-51gS
HFRY).CQ;Y_dG:d1S26f./C2C1&eFP&S84XTbEdG#7GMCb?/O74,8;SgdCJPC]fD
7KYa@aG+_8:B3_7CE>Z&HC>5&1UQ+WJ0_+L_f-bP.Q8^(eg9V6A^(B<T4?;&8F:d
TTB4)&V)F.;F.QX4]7ONM2_.&@^cPS(7AW9?RW\#I#b+7BD;.8c\#JS1d5BSf6Rc
cIJWZHfgDSG5+54aHO+(DdT0;NCZdWD3/]NFBIE7SaA[._RXa>POBc]@@+9Hb)g,
YV:^eXL3[N=B4;X?g8YO7:F+YPS-O7Z^?@YVBH5DZ4CK4aU^)[OKe]-JXF9@HPML
S3KN8M8U@3a[IGG5,bB0R6PBLfOD49R<+HdP.3R#7@YG_)->+(DU#]?3e8R?g:gb
HcgbD/c#]\0DYJ[Xg\&X+>CGLUU37A(BLa9>P2=USB^?0RaQ?4@a_8:N52MW]LTR
^,Z>A^EFEX+9Vga:):dXAdOU_Tg:D>_C@SaD8;cE@UX,bbKPP[=9VE3-#JK[DFbE
#ac)XQ25fR#IER6)aMK6^9&Q5]b3XO;QD)aG9TT\)H0fH2:0+?YD?MC016)C@W1X
/S4J.B2J#Eec6JW?G:SZ2OW8,e@&UD-><A\AV(2R(-+d:G7:]<]H87#Jd\SO+4WH
E3O=SU,;DLG@^#?5V<)=\G@G)^bcA94:f;B7BH,O0=FH,6FXN<;LB1?DONC^_bOG
<+\,R_LB/BKaYJ5PIL+2@I(A,A4XdZe1QOLTU2&G:TU>ISUH:]7A)^RL;5+e1eC^
.+S[,WLA/[/77:Hd4T9I_e?JO>faCa9^J8F&/SX-?ZDUa-ESdMTP=+LaE0H5A\]_
ICbG2O6)Wb@L4:_Xg_45A^VG\KW=-Ug8@4#1UC(g-cCHB?,3Nfd,SD(]I?T6a9OX
Ue+\dOYX&PKQ3?46QK8Y1/8V#18[T;g_VW-)(2RLb0+GWW_ZYcU-<X?;fRYbJDfb
[dCc^fMGRYdL@4f8Kg@TZB5IBXCfd+GDa=Q)-C(:4eZE3Y\>g27=c8:_EdX^ccSd
:[N5ZMS@UNQ\X#Be8)>\0;+3P^Z?=X<;NGM?],P#d)FYYH#WX\S/L=QS\846S;JM
/fI8&-5=GE\RW@KZ:fS0d^D\K3#.Rd0a0f/C5D]>HW#+Q(FHU79<==FJQ^,H)OOe
ES&E=/UYG5055.Q3Kd@G5a9fgEeeW(.@;:?[\>b2(&-51J71>\-H\B8SdBc9Y)?a
I_//]X=OR.S4B4.?8=T486G_NE)S,g-0db:R?[4dCE1BG<U83\WJP)=26WGF#I-)
[b8P;XbaA+TU&RI=<R:YeYQV4cC8g=>SYNVgW[ZOBV+fJKB8G^f,SLJ/W6f^U,GP
J[?3#N-J65-0NfD4ZPD#V6FdIYXc]Vc.TYS6K=Q5G@BU:g;A50fDd^WN62+D?2B[
eB((YFRJ?T0^NO5@Ug3G.B+X2U5M(Xc)OcLbOHdJ27@2ZQ:dKLa]f0FOgV?-WI,0
GJ8&IJZ4FMEBTb0EA1=/c::g_\W,E)P=f6/+3SOR;8>Gb+<WMeC7H]-/WJKF;OO5
.WdCaWJK-)b;22,2MY;]-SaZ<:ac(#P_bWLU<=TXR/8e(=]#8F]CCN4YO\[cQ3SB
LP2-SMR33B)\ECP0FG:;7MXA_^R(M:&F4VZa=@B6EaPbg4B]E5T3:QWV4=\@2YK+
J(VU-/]8>;CLU>g:HPg>ba7F)^^@&0MK7J2:0?\JI;Af66(.0_X&;&](TbGe^ad8
ZR4=d^MI:e3GDC-U@6<U^]5GNQRe0?\MH-7RcB..&@WDWV25;(0.2U7)Q&M@=V&,
IFA.L8-:Af&IN8^#bC4Be9A<EeI^\=&LE/\Cb&F3(F-K3S.[HPWeW5QIN\#FB[G8
2SE=7I,,:OXN82Q.#8U=ADN5WB)=O16\?@H9?\Lf@R.)TY0,]FCSRP9S67+U&5.O
])B[I2]1+Z6d<b:NF+QQ51@-[B(=fBVYT<6=^GZS^U4V]B&eB/c=L\4A2ZV3;#Ub
AB#CR44.Y+^RQCH;3O]>U;+5&E^31O,7Pc9DIM1N2/P/QF>37A^Z3H:]<7^?QY4E
MaN+Z=)EC9Y9>@?#e;THIGN\#aN@-WFReV6<NNVNHP8:0a;<X8ITe=D)0XE>[VeQ
UZf5g^_2BQSQRc7V\)#9J_8]aGJ,,5BeEf()/Q.7R>JA81-#HU=Q(2fdQ.^2<HY(
X.F&P[eSKP/HT5\#.[6a.0bIbb+E2E@M9=-FeaKFZ@@20XFFM\g\#VWXD?DLM8D0
>.N)L(=?;VZP()&LD,@GCaaXX:7T#>+J,YRgB9CF>8_Z;/N(REX80JU>6_96HXW6
P5M@e@AgOPBa?GVL+#A/,VA;2^F_HJg]:KH?+.Oe6f.;;A4WVDLWU@:T;Db)0Bfg
&;K_1\LaaBY,^FJE9cO.K/MSG^Le?K&4M+5.Ma^^[S/6d1-bZTAdX(g7]F)f>KGO
CP+^(,a-dB:@DN>cKC,cB@=fIA3eOV<V2YeY\L?e.9bU.RU+W8V\\]\1W:LW.f94
SddgdG<LG3]\g4Y8B[f>Tg=MC6b:+fcb<3MWKJ4K1)eR+3Ef2@g<I>K<\[dTgbC)
2&JQ^5-0N[@M-J5H?Y#<;1Pg/VA1:0DaSV]SJ)\Se[dSQ,YJ0ONDT=B@/P;IdbU:
.4Nd&Kb+TCg:OOP1)]@RX1-U72Oc0I1LCA4&FSCP&AKD?)GSRLd4fJ053I5&_5ag
^-UFaO<K@g_C]K6,F>JZL_+PU.#;Mgg(fP]3M=dFN>I9\-9@5(<DJ/ET#-1a6ba[
b1?c@LF5,/c3X<+bP3]=J\Xb1PdcNQ5:MRB2:S^+:1R;M0)]9Q8TeO<afRB-76d\
&Y9gZ:F<O->35MQ\3La8VN5>(4P(g6=fA6Z3LFa\>0feF5^1/4Q7KC/L/T(W#_2]
[+RA(F3?A<ZLOMAQ9.MYAIN05bBJd?eN,Y;UO^a9aWB.Rb)fg]_e(f=4e&_<WZU=
\3PRR=B.MJ5:9Zc\;bZ5f@25Hf_PHA1],Nd30.aAfJJZ6Yc3ED0:OCO\F\;?O:6X
B3+T+a-g?\b+G]f3f-T&>1d[B>#PBd\9dT5:]?O^aR@ZUdM.#7/B<01-AUHaRPUa
E.8=K-0dD25/cUE6^VU(&RLaY23#JGM+A<@9J]N[HF&7]5\9WT^+7Q/1=Y^9QB9S
I-M1?G:NJX+48R6,/dTdEeEOJEMfd7,:/a=U];b+=L<M\KQB1\=Cg\?=H]]QN>Ic
]E)BE1],G,-_WHG0(dT3<X/HVSUeT)QS2QCX[NcbM>^BK7I08T7EA-,G3\Sf)=+0
aZ:]KC+\TaM@F(.XbD-U9L+@2^8)eZcc?HM5JZ8:G6DUe=2M-Z5X7=_2F7ETH196
/SY\[(ROUg,)6A<UMb?Y8d9D^5ceXgg.U=IV6T2AIJGg1BTWZ4EU(A)L=UR9#fN,
W-e-]KR9,50ZKT1WVaN-#CP7P#C=aSEN\3d1&&4.Le8@D26R7.gbS7XT29FYZWbg
L?WMHRZeSRQ\NTSYBgO/;4=\W5DB=Qc]&+Xe8#TUPANg1E9AD5]>8\dAI^fZa=M3
,MT/g?:N<bWP)4MRb4&&[E@PfObe@KDd^[MC,3:<N_7<3Z>=fT^ZB9bNNV-M7B3[
-I;f&TIGB[+-dWUBUIGEHccCKU>CU_+4f],aaeU>g0^6c>0@<[JdFM(HL1:=>)QP
8dg:G@TU>(T)Z0Vb^WbEc&IEUN(94@GIWb8Jf4YP:X,OR;26d=DYU1d\8M0#0(Y?
M078DdQBZ[aV[d9U[N_&]M+QE(0SES7N>77UN\Ia]>TY@THBd4U&(RZU:8FFLDEU
OFY7PD[J9>c)c;8@1EOc4V?8=/_;)M8^2I)J^3YgLUE.-Qfd)C;&\+]?/&;_-Y>V
>ARaO--RSZ8dN<7BJe-=#O#2T<7THW6P0g1^_G.&RA\:)cR3ed4L]-Z&4APBJ=UR
CTPSAF;UE,CD<AE\_;\NM0W>)8Td7H]-VE,6J(.Z(B@XWI1c(E22BN.5(Q_X;H-+
]=W/OUcPc4.&5V-&9OIQEH,Y5MFTS)PCR^LRE.9A7[>P][&F4KGQ5d:W4ACN=c;<
7a8Y_O540N\D;=?TaLM]/:Vf//S<^)N>.)Y1BgHc6;_=(f597fBdXHTO#>:0IdY<
<L?K4#T>_,(CB^:J1SB3U[8NPQ_#-DQ:cGL3TM;[LJ7Y&-=)C:3N\eY.R[@a1K+]
8FC=I90J-AcWKPe&fV^-U4\SC6M4[e6.bgE03eY;e3Y;FMaQV5+<F&62f#gbG59;
fQ\0<a-)5]D-SWf\Kd)c^?c?bKe1f6U0@9>?=A,Q@aD/V6fdfeRX<9MZ816AD45Q
B((S&Y^>RQ2]Q9DLX,VHIZ_H/_e.&1?<,2bc+Ab)8\e>OTRG^,Yf,7bUWa>NZ)db
4^^USV/&-+EII/CF0cQL,db4&;36V:+.Z^.VgN=^\aHAWIOB93>d.J/fFOSe=KVC
@;J2C,1_JKaIVA1D3,[U@S-#H7&aSQ=VQeN#)9F?UCQ>Z.He(+9WQ8#SY)O:TO[D
?bIf2TSRc21>QT.U4C__Yc3c2<&#/VMc;PGfV\A1(M=)EfB96KXSe==<J&NA\N3Q
G+NgUOg.VRWd?4@UcbH<e3FeQQ)CVW@/<?JN8&KEJQ(L3d+e2HH59RDF/a&g.5GJ
e8cJG<>&Y5c;N>0&B-[BYRY5d8;Z4/;O9Be7d4^C^g);ILf]F=)K)-XbC]OS>H+<
]7N.#@Q1-F&()/>O;4L)8P&/RQ,eb-&BW14.2\4a(,)H\T[YZb\I(<K/?<_M/@)3
CH<IC^=SDW:<W&FJ0Ob(AT&H229<Q?,<3Cd#bdc53a?f@RK]MRN[I[+fL/=ef[N9
d9c^(K3d6I4U3#D(C@baO.76]@,:2a3e1(++7LC]F[:\0g)=I+aWGW+Q[aWWCdF#
C=WYRDIGTI76:8]b52acg,?->6g=eAZe-JFDA[E;^P84BKM+7KFTgX[0<OGd&]d/
MX/V)2CeQLQ5d./];4b]Q5C9&4>_0YS1N,8(aRb+[]c0+C>_^](]WNCID,>;^cW(
S\1PGRA8:.&<6?b<dO3[-aSDaISPM8d@P@E[X6+9aEOD#EQ\,@a=-?VJ\GHCMR)]
C0b6]SbOaD53:3aaS^E,LSI&V4\3.B^bGU(3X#((KTc#S[#JF)OLF<EAKX[M1(RR
CJ:G0YP_f];9OTX<LF.D4/PYdW7d)#P3XaO3Bd9)9c@e)&<=Nd[C,(Q@D>-_D,[7
AUPHHC)Z8g;;,RLQb.N[JEaZ/U5E,FdV)V@8X-?4&6[7;L5?KfE5:UTP89bTI-6I
&[.;5gRWSF0cGN7LA:6#/5@bL.aDbA]?B((b[-a89C-5\A\PQc]X.[^1@9BBZ/3>
J@X9)N(QMP(-.ddEI.78V\;ULZ.,J,[63Q/07>XW@C/&:YP@:(M:)&-J<QgN+(3Z
_J;\^IbLH6-VPJ^5)Vbf5:<S1b[#4c0P7gKI]L-;V76,eB5H@5Q]UITZ5[2]J2AQ
:Df^=M(U1DX4Da]T#M>BH4443):K?bXaBSXXg0OYKB)GP/2R=1XY5SF>fM010,3?
AC5SD<0RV-a+@<:C#<Hc-U5LH.HP:<;2T^07_g,(F118:28UHgd.B)KQ0+T,2&_(
2APX-7@I)<W/2dB4O+A5KMX@CZM;a+\A+J:T<O#YTg<b2J50_<EW68P6cA^&JHf<
B/V]IFJK<O@[6I=&+?f>8GcD0Ie0V;9XW\&HD01fAKG&GD8b=N;g#P3MH5@-H\6B
QEHU0,6GED_3N^Q0L)Z3B_^gYR:5+1[>;-5J5U<V_bXSA?5);[Q&Z(NF\Y5B3MGO
@O.NUaRS=[>6G,\TaLFLB,L)CA0CLD)_]N3B()F1DM>[4D)(W9J\b^H?C(,VWgFg
SV#L)S@IW]R@[A-PfG,aR;7UX4;7A@:IUe@JRT_IO8FS3^-M9AZK-c78APNc?H52
b[72]KDS83P7Q2T@YP:K?M(aLfgPgVY,-:U]NBK#NOL9N8U^6;>09M8/aY(b9:P?
:J7L9NCMDR>-9>Qf2]AC&3JDg;GM>@;?@#S@aV]PRT76.[g:[C)&V(&fcVH\S5WJ
G:f8E[?DON?gMT&5\K=R1e6eCg;?eT&cI+XORZ3-MJ]],ETKR-Q76f&6&EE)#K0:
9-V_d#XP@6[YV7I0<WW,Gc:=_#W8:ST_0+Z#3FY]^PTYY&37G-#RST-dX;OX2Vaa
48LJ+eO3cD5<(JPP9@)80I5FYRIJZb&8eP<.?]S@C#9GKU2A27aT^ceWcIJ6JRTT
Vd1a6#U+0HH))J=Z.:[Af]#[K?YG;&b:[#b(1dJbceXB#2(eMTD/2(cU)G]g30@1
OPL,>QFKD/_f(T^P)0<2B_#E=WE?,JAJK5<REH0#10fTSKRY.,aAZ>3NETbFZ:UT
#R9gB]\,=7.?ad&ILbYP&)d7Z>(MPEL:YXdIO6^BFGADB3Q5K.3TCO]]@;BMV,FT
M<[F?I?A85)5eO]1VFCMW:5/1de<feX:XL1:/N4Y#=8@POMP9-N]95Rg,C5S4MVN
(MB,J+VT[B?;V\CU-F#9(&F)]/3_VM/Z)ASVLWBF0b5)LX@(ObPWC9K7?LLaM\0Y
Ne>&#NcZ;HREbbNV\^;A,E&B@KLE;-OV;9>0Y,\BcM\F;CRcM=>d72C]HNGS:PS6
G&9DFW##]c4)1F]XG?Qb@+L[aJS_?&&Sd95F@.gB?)+H.NO1geA\Y12>\T_C?[JV
CTHWPGV<>dCCQTCWW<bd=1K6M_\C0D[?<4+.cOV>9.0OW5c87CFO.Q:_[HO]3BO-
e3U0a8X;8_)0W)9K)CZ(V0F-[GDAX]TdF:[cL(N2Kf^Ab:b3eB6G5LcN@dT9dWe<
-UOTLD<_b1MJ-,LE+@)P909GfHbV-=&/JV^AQ37JU0_A^8]9=L,I+ZRHg2HP35Zc
^@I)Sg\\\.NTW/<1Q?3=FB\eDg4W53d,-N1JQ8:aJJD309;M<0C)aE73>>2d,d,F
<3P3dgXH[?GMcM/Z3S49/bW6:K:dYBb7VXV@9a91@=(>J<Qf^CQF._cQN+CT@?X@
BK21gV0f)b?WDVHUB-->B?[a#@Z-I^[^Z7]&280^IdLF5bFf\BL;Pf:-eXJU7I1#
^=S8T24-U=dV8E4W@H;WP5&D.gSWd-AIDG(aNc1>U/\-D\_<[Ac?7/_.2SIQSFF\
>65QOD(^dg2+;e0RVcOU@2PA-7U:?>L#b:c649(&E#9a,.FaOKH2fU#gNP&c@)YS
<BR+_99T1W(034PNG-b=?ZcMe?cg>+J>X;S:X-]=_##c+;L#WG[ZM/1R&V3&g,MB
^VbaG^d^-D?WT03K\Y_1@2(ZNKdS>H.Na+QH6(CGYJG7F111,+cE[>F2g1bA=Td/
f(2b_20(SH[TJFS&9JHD19-(>Hf^6?dN0E6_D^>8cNA@N[SY6b05MWOEMF)/dYGK
_D-EQTMbS7a>8fZdN.-9/@41X;e;#KJeVT:^M1^S(JXBV9X6\Wd7;ab46MRCVDZ1
H@FcXS3A2dXLdb8(UV\7G9J51@+9WX<NZBXc2GVW;5T;fTYV<YgJVTb)JPP6.]_#
([)AV5<,:GI\DS0GJ9O[cXQT+7-5:GPdV+S.:2P^Rf48[P96[1#J.US=fLF4-1QN
5aP=@W:/;O+S+U@Ce9_ebT+U;gegXE3&.A(_N>bT(_4gc.H+b52]JJO,3NP+?aWc
:YU^;;Jf#M<d@I:@5.F+:8g[C)O/G-KD3ZQHY7GGW<<>UAA\2&#E10c7gD#PHgf-
M4^aUSY2)3V_8.96AHK99d6=884f09R1=/?V,8DgSX0&A/</C_V:C\4;OfX(<VI4
#?/bC;Z.4@.D94_,99+0FYD^e/5=-3<[UICS>Q9)Y8-TYE&6NTUg(c\2MSDLDT9A
@(e@>VCb;b\Ke4K6(;LPd/#,G+bZV9OM6UQ5\A&TCMBNH2&RMT=,gH\8U-Ge2K7#
Y[#Hg?Qe3[U\?R_aDI@YHd[#D@G<7&NT.GO<F?I9@XUceXT8N\DUJ>eeX3e,SI5?
2P\3E/T^&E/)W(6&\b2C]O>?2IS0L&YEd(K_VJ4-;DbYF5G3#?837)/C73bM(:6e
EUO^e9O#J?IH5G;=4e;^2O>aJ>;0+NggJ0YJ3GT[@TBf_FgM#ABU2J&ZL@@6,[T)
14U-&a2.,Q/?:gJV5#ce6dR\O-XLHe:YUAF(L0dFR)BYNcC8J\#e#2B.ZQ6[2&,^
5b/F_9;^98QbB?3&[72b^f)&<\Qad]XJH+@\1&d4,Od1>C-N)WOKb1AcF??8EE#3
.>[Q#(@##\F:8eXTH&9T7G&3a?cA4+]MD15G]\bN_e,(4X+Z82?VE;.UAa1R_5YZ
?(X,&.+#MgT6[;_(B4DTTI9+F]7C(RVBaOJb(dA@G0_X5K.#/\b1&L;cD9LXb99f
(GOXG3W,7,a_H4bQVN_2TS)#&/KIJS0;/FU+O.AB50<4D-<W+LY=Z>2VGd8)&T,a
6&dKPL)O&UHC[-cdJ]bIZBWRNEH18\FY6&T[J:PB<K_C5MM;)4-HZ7MF-)(_-De&
SKX.TVI>L05:K2d^dNWH;1T<-M4d1J_TAF=Z(N]2R9>6BQL\O7A1=[:c==DE1a;Y
MPWFD>E@Y(]K-DV0F>)0D(JDFC(I79&XBI(&JSX+@,c:g]-I#K.NH9?4QU/AH/.?
5[-#;A186UI\Z_#IOId<[Y4GJ5>PMP3>;G4.aY9;_#5E\WEeU2[Z8X^]7d+9=AfW
9VK=&CD4S+TK44U(\#?3XB+)NW?V^\RR=N<GWRSVV#/U5:O&8+[1#HK0<87T&1,1
67bI>-cfcEa0g]P2I^0S@XZ8]?^T58++Y^d6\dKS4;4^>;:FWX?cTG1DZT1,8Gb_
ZEM1eLG<GAFAN/2&\KTT8C;@+GT_];Y3DJGMDM4P-97WS4&IBaF==.TO5DKB;Y[5
8JAb4=7=M.6E]DTPZJ)GP8#g.7#,+(T\:(RP)PcDS-HE<C6.^]@V#QVPU@EU+V>H
e:DT^CS;T1c]c1c_fSYG8&,&=(?eVOL,,M6&87Y<1+4CLTPW.,7CZ,WOZZ,+ZAIU
5T6VVL?DNd^^,DSYP&/c2R5PdRO_e2f=^1?N/^d^0NL/T#9&G.-_&ZG<CMNBHOH:
(fQF^e1[5@C/W2/4@?#dUO2H<-#MURadd4VcaP3V9I(N0T1,D>1U89)6\f:)EK&4
E+\Z^LbdF>EQSKH>2N&fRLTGe_XF[@P,=Y=^cYOR1=cg4BI1#_<6GHHWEDSRUW44
7PO5eAP5;AIaS3=48(SO7O4.e=Xc,8bFb7;L:&NYCS@,AV^07g/-Y2d(1<<2e\g-
X=>5CL:c81ILKZD1#X\Ie0QPEDLD_00UQ=@D1.5__HV4\47MZ)-(EPF,dDW6__>\
/3Y=.KZ\)I_IEHNO^OTUAa/<2[c@a[TQ2?++Nd6W3:_#_Gf2J)f92.a8=#GHHNGc
>U?T>JR3UE#KA,BJ=f89FD4=7F3Eb2Y\^QS3&eP1BXX<e)dFE^;,5X3>U,2&Ya0&
KY\R:M#bM^+>A]cM&Q^MB#PTfAH)K5LZD:E+ZLE+R[V?I;+<BG89McTY>;7)2\eD
O(5[\8HD?dY^=_5VP9Z(8@,]Fg@_YT88B(9@/Y>()f6B4X3K;6D4,8U1&aMCFZ+]
Ld8:)?YbQMA0Fb&KEIOM>G-KgGJ6T6g)?KB_UZWW_/GgC1FK_FQ2^M-]9>U#NJ1>
KF>.PU:9]dG)EAAbVJ_Q^2bRU;BAVOD+@@2VZKe3Y0JJL]W.>O^Feg1#_)ZfgTC7
T:<Z0VCReSU>@<K2N_g35HI.=a/>>b,,FP;BUDO:c[IfQL>KCG0QHW]1J/,[6,6K
8>Y+,#FD-&-c:TcFK4U+cYe<,)ec0/C-YP76=BR2,:_>#7V;(eIRQc&RBc5aHQN<
OM;CHFY[29d+bV.\#CX&+))J@S=gH\UIK<ZTfHNb9FK/;@Rd)ORPBN:aBd;#G#>a
M2_,+gE)7_1<H>+<AR/<?[W]?)KP(7V5/Ia8MG;#fF&3?VE]]>3PV4g1VD0K;[Kf
bF&@#a,US^<3Wb+CfGMb5>-eO5#RFgGR5+L.O=;G5U6R/XQDBP7]f?FX0VBO#Y8I
S/MI.^UJ(\Gab8a/VT).;ONE73\SA^fJA=ZL\g:E9:N3\#FdWeYVN;YGYN?7_.3O
ZbQAHH420-?/95>#37d<<f&DV)4O&P0A)B,=#FPd)U1]#8fOF/;BW9cS>Ha).d,V
Fgge=fdBf6^IgI[XL>d:CIc_Y5S]5^^SH,(Y3S-Yb<Gc+B_9c,1;#-IKIMAg82C:
3H:C)_5F.RJ7HK9SKMW)JY_6QaC^E1R-8eUfW,d6_,X(OfQg-V+A<(Z9D6;F:HGG
WKZcEOGZ=Z&NRH..GF<JC1^-00ZL_VZ()^C+=)NYe19)bZR-RR(O1QQeE3DUHW/a
,)2G^cS=gR<E.H)f[,B\SDe\1F(GOC[SHRT9I.]/B1C;#&P]>H(BCJUWH==,Z>8b
Y\dQZ3BI\gB@2U6YH#E;O8DgMU8/3AP77YMNWS]eI)<WIgFOV6b8H@E;.Z=bP\3.
2fJI)D5E5&/;)SU65ZM4G.fQUD@gIR5Q7XESZW),=\7LeQZUL9S_A[0S+3Rfd^eC
cVR4,V]X,@\SgU1#]H:ZgMQ6G^IYTNS)I<1Z)<P_179QEC&OV[CBgXV7QXB=F8V<
(K-JAIU6ZO2V8M@2c061&[P2[LDGO(S]U;:^P:g#@Q56?/aabQW&T?Z5feVF:9\e
>_,MRYZRd.W@KWgbF3O=(?Z\d+CH_RQMgbfP_D>_Qe[:3(#H.5<G>5QV_E9K=1SL
G;1LI1c]OZA^HC+c7dd^e,.QdLJ1F>GAM&UcY\)[4(I)B90b1UXI&B>a@U<5VX2<
DgV)A&/^P_MaQF?@_2S7-&H35aR&E_U(8U#VA.a#F)PATQ,>NL@1a@0(5b#&<gZf
PE\:O?X;d=d5f:_:OQ57=RYa;(aM(,dAX4_W_FY2KCc82.JIE\9MdO;aVMKC[]1O
TV8DJda&A),a[+-_,.:FJRZ&]=F+,Ha6:Y8;I&>SfBVR5Cg9M,(06g[CMF5HI<eZ
(PGH.c@+/D042f9UY+/EXXRCF)NT8V2CZO(&d9Sd@GaP[ca(]eFRQU1P\SO.1)XV
U+<().U8EUGH>d4H;Z3-3-&@5fe7.YQM9]KWYb[BO5L]/<-0R(ZX+?]SL[b:NC=f
c7BZc0eG3]K;9[59^GD<WR3#I9@8IXL?A\X#B23_\/0BYA5E720cA9RP_a=J0>5A
07E+g>+dDMLLfT1<.1I@;D=5)I<ETbC5O0b]64bM^0),_F(f\JAAV,bCE,EV0Z;W
AZ=_.4CK\>..dP3[57O3<SF=R1FA@&W#SXB(N[Zb>#YDVR(AQ#_:cId>7E>^C[N.
ET#S6Jc\JL9T<>3(de1K?fIT52U/7<dLM#3?6BZ=5JCD>b2^L,c_RBY(_6=&DdG>
83c[027O?UXQPM7GQ]3eC7[/:aL;cNI,+LRd^F=/C\UE9_06[YE\5OKVD=a<N(Kb
@_eNcXRMb5)^+/T:e=O1J8;[QcgPW-8AA??-DgF1fZJe.IFZH4#aT27I+3\0LC\#
-MS#;_RR6M_H^Nb,McTf+3/)8H<QS5>@IX1\<_PX.:bP<Ua;dBQ8gf]PW][KeHSM
[LOVIb)UgAWS&QW?=]aEJO<BE?E-DVMB(-MI@VZ=DNUG5.d@1FfQdf1^[eWL:CMg
c+U5>B@McEa4AMLUG5GGb3Z:6ReccE[31Z<>L97c<;4McQK]J6#K0WZ3g3V-YF](
O,ZA^>Q]S@88TE3K.39,@g\S;S,]:IaBNV<H.G@dcDX0/M\SgP:BTeG<JT>[GM2A
?54eY:T((6GM3=D5\H62Y9^GM/gJ#BSd#J@0P=RIF\.2YKX^H66Q+)<4/:QbI[=X
RMN-gQF=<Z.01C\QH[;.+Y;aD;d_V30#e;<@&O,Z0_H&V.gKO&&C5Sb_I<7KU?eF
UXC<_Cg<Y_b>?,>6Yg#,0R5MY@aATYB515M_<BC.P+;NfMa<VR7;+TM=a9Z9Vc07
Y7f4XGTZEBV?[V,#Z&EA+@I1cKZCeXRI@SF_RKYfaeD[G)dQNF9)]c<^K<(^V]S;
ddX]SWD+H67_B1b,6)U]2Z.4=K<ONX[I32)8b=:Q2UATE,(96_,V.[f=@D_I:PTb
<K@5d46<UOD?T]c^Z+VTKZD+Z\_6N8R2D\R43/\YEZgP]bXUK3]DMZJe(&3Ue^S0
2Y(T&X2WPQ)FaT8SG4\\>C0D(::a^H_C#S^MUBFE[E-+JWU\b\N:LKdWcWHC/gU:
P^9SbYE,42MGN0-TH2#NbH8[6b)2ALd4LK\+O<=c4.JQ[Of=Vc1(]#UBFMXF/)H)
ON[K9cdBTS[ZcI&)TSScK@P-,D22K:X@L6d@O?P+3?0D5-@WI_S?=:X39>X#J6;&
bIa;Uf2C]bRUcBJ>Sg#^3@g\.SB3V@KTY;2SAa[48(<.aAG<d;ANA7XYJ<6d&Q<^
:92Fgg-&)V1>-ZcB.HT+HggY.HNO5=J:I)A:e?#f5F)W0#01MaH#>F=XEU\?gQ(A
XBP2_a2+1:,S;(R)aLLU3.;e6(G9T0bggU3/MeX?KQ9>FP9X3gN7F4-_\[MX^E=-
O,2NZ+d=)[8=J&L;9+7(-/?N<?G>T;^L(5F<C7TUM)]C1+?^FY>[\8eO>DQS&T)+
1).8N0NV;&Oe-:_FEb<>QW=T2?>_[Yc\WQ\D[=_Z?TBb)7ff3Y@[(7ec7b]<1,g^
fNI(Y-.E;TBOd2DYZVUg3a^,YNg_]77R]A[3JJ8QYg^C1fg)Pd5fT4(cL>0IeO88
,8LBL6eA=P6//DNZEW2g9&,TQNT,QEU4>4D9>5)D[+8R,CJ9fB_B71ZgBSB#aU:C
].6.FOML_R=\@Y5U)ZOd(DKC2_8=S_86;)VU/M1D[&SE@KP(]QEQ[GV]LHf+.(:=
H=0PVXSRJdN9f6gY4CXVSUQP232GH1Sa\+NG&e&I\AP]fA^@YS#G\/IB6WZ@cNDb
1=QV)U+@e1XVS-AH#A(D)@bTUaA]/9L55O)KJJWE#E\64353EMAF4U)f1IAKP1V)
_99EdSV>]+5ND]T.R2L2B?[.J>cGLg=?KB]H>_FF=;-.a4d,Ee#FQg7.SIF5c:YK
gb?0B)5TR[a(d#GU&I(F^8(OV(Pb2TE:K8abC7SS9M1AgM,<cF>7\b9AV2..-JSa
[/HM^^0YfdA41LcE_ZAE7ZZX\7,Cc?59D.#B+J7+=fU?7GQ^B=O#9\R,G.;(.?Yg
-7L0XaeNM7S?Q[&06UW0^eaA(._^@>);P&NH42b[XYY[^J#/1]YDLZ_1g0EDP?T[
GKTa(0<?B&)aN+WFa\=,_^-Hf#?a;f]\S@(&,Q/eEBRV&LQ\BH\ICGM2cU^N.c:)
EcVU;.>,GOD(V>.#6E-.86X,:LcAdA=)(4\Ea+EPcfWDM#>B)g,?6;e.V>Z:NAE]
,T4EZfePPUQa/=F>IQSZgEB7HIO-d8_)c9N.3<2=6.8A>^9(2I.?17>K:R?U(H9(
79A\VCeWIb<><I3T2(ZeWFUZGAf[bf?E7-dc]_cB=bEUNIW4)NMS9c4/B-/OX@S0
Y?ZFW237G>Ae3AC9Bc3HM)Z(P-Q&.0CcL4ZabJ0f0=EW:^HHVFQ_g@4e3VC3Tf2#
RKP,cX0.)[9A?W4K^C:OH^9CX1#BHAZG;EVafCX67I),VJ69Y._gDGHCQg.)&E+N
O+A&]S4dNJ5Z\S+IW6@>NBQNPG/_H#Hd(D:_V\g6I<\ZXC(Ja/?4-].f8Nc7,@1?
^/[299gFbLSW0TH:OY=U.@(LEL/?1F+60d1R<\g<F_=>B@feb2[#9ONR[^I<E4\L
V)#MI_M-Zd??:<6G]]WL0O<0b1[ZE+9\gG3D+4C5N.&DV69ZSA+:[&d9+25EYD6S
KI?\A&#VcELMP3IZ6\MT^\)X1[3PSBZc8_f()a,JJ2?+)2FFLE\5b:XH,>&5Sg[E
?H(1c1-3LaA_H66VGb>d\(6Z<95@YPNV=f>#M<dW;U.4fB-9#P.]>NQPR:JI7:V.
-bS7B>E+)^b?^?X^@M8;+2dgA[L#3Z,7<;AbS5aQQHgX_#_#E3.VK>2ZBb;)Zbe8
:93_^FQg3?QGLK>2KH9_I)aEVV/eV7\3+8VYJTAP5b&-)fFIHBVD\]2SO#R#=18@
U42S?e@YC&8:+N:2Q;Vcc5YD(D&63FGRF?MLB<,+C=:ENS&XE>(d/K>3(#^>M<&K
+);CZ4Z\FFCQ++eeMJb]6V(4TM&2c)_J,H2O^E-5H_fMJDg8;gIN1//4g&G2d/Ug
cc>^O7K[P4K(S0CF#eJLf)/JIg1HA0)Q?[V2;d_MF?eP;E<4S+VW+2DPA=\b,Y>c
\/GGC;<aHPaFI.NG#;]&P9g&C[87BXbH,>&Y5C,/.:TMf^SO]=&-a[6cd-B4U&,=
7_QO^+TdV6TA:+A41]T]e62fI#XY(#@0(5JCZOEJ;(e;IT\,X5X1_JYf+_.:LHUU
.RKD39JaHNH<E]#G_M^@F(8\.6X.91V82&)Fd=J\+8_WLR2/Y^1Y/c62#H&IBQf[
a:Y=+OCd#B6a>Sb8YH)DT6S9=H(6S5eI0;MEf.G/MP?QATgI(/+KDN;\?IeE?.&9
;ZX3@9d8b&LZ.c)6?RHA^KIeC1?7bT>G\WGSJ^V;)GeJ@990#O0]G?&Y:MNQJaQ_
Y<0PWP:0+=1QfU7S2dET-.>eQ)Q8\:6aEdOg4fOM[9&/aYTJ-S-U7<#:DY4(c=Nf
6-SHRQJgb;OE1]M3-0JX[aZcO,\OI^?([E6T,RHW5FP@H]8P6\+#&JU5Lb>:TU<,
6A00)/),a8FK/d8;L#16+/FMg1592JHg@,^L-_=FPMQ#2g=MLL5T5=8D(-LFX9<_
/:SZ,H-f7.L;Mb)LK#0L0[(?Z^J8;7K7,PW)+[8@E.JU<B24?\I1V-aYM9JI>_Y6
^1&+.ICS/ec=^d(#3^T]E?MA^Q6:ObY,&[GVEL11U?OaHbTM_,e(Ff=@Me>gVff+
:Xc:],O2f&D)]WbE\@AS8NI-?Weg_cfH&HKD71]D,fNeD_ZaL]]@+M85)+2Pe>Ac
2+A:>[QbAUE1;N9>6,69KX\ZD3;/H58GX;-EbR2XTJ3G^GcS7M[9\-3_I9>3[YWa
WBdK(Q)]/?RDWBAB[)1UY=KF/.^19Z(SEUaEY]0,Hc?c1Q]/.,JC378Ub@<,HeMA
I@:cOaQb]B>GBXE58EZTS=A9g;FF9<cN9/<#f(Ed7HN<Ggf0SJTH?f]9E9JVT-5F
aP#]T07.C;ELe)F5/YN#5aX69+.9UF0D[BGBTTT5Ub]QV_J@:CY_FAAQXH3?I?<L
UH1PB5cWHbC7,4;8/OUQ&M;U0b@_.a+c_DP1E)<1EL98_3>)G/H8]01^O)H[Z6>Z
VZXLJ>U?(F.C#_,:b]AVTASM3<D;f\WS@<RD,Kg(F3-cb#<]RIeP\#;&5E#H.[5P
+P=_\#9+3cT@FUL;IS_cS@_E.c1Bd2L&+RWT9,cWH>SZD:\_9<PE@N;5JBCN6f0.
R[)/9/?8ag,\3K0H65P790^_aPa+8GL(_U^e9SW+T]UJ5QdO?BY1a;#B;W[ASDS7
+H(=2VcRI0ERSgC4+e##.f8=)B&E70JI(:RGbMU^J833AE0_?SB=>=eN+GDeC^5+
R?7HRgf<D:V0H_.:;2(YYMBTTG9RY:CQ7\+BdQ[a^e_K38^fee;JF)-G=GUDIS>E
d[>@,H4+80^C?EC2F?A_EM/Q1HHU28JXd>JRd:TA<R<5=[9<P[2MJM\gg,:<.;3a
fUU<??HK>TO25)VKDIO[_aVc.;54bfE>YGBdY5^=3;cfEI0IVFfGf,aS@)#\Z?II
A_+EM/>.JXF=dd;D,d;VcG>=5YdF9UbL<I#6P2FW2:@D4^d7>&O_@XBQ6DV]eTae
&Gge)C;O#[O2=G\L45+LD)4AHe7Y0,OcU)NKY.:D96.K6OW<C<F_=5]E>R?6>I.(
#7_IX:0gRf,3@aIS(^Y04MT7Z,fWVWd2::G6gc;J(;MAgb7&aFR#20FL501c5W#0
DTb#gd97&D-H]+/;a7DYePJT+AOe++,GMU+<5NPf.0X<-#H&aMNeK>?-W.aVH7OO
LBEg]UZ,@-1-_R6K5<P=VK@BKE-BU@OX8bKb1MNSe[#5?_&AU,6:YZCLM0=:19R8
NI@V_d<1C1Z4:W_M:H>97(/FE1?f;0#?75_\X2QZ3acMD@2K6=S.c)MWg@\GFOOS
6@NVCe(N[_?K9Sf@-ZV4b.N7ZJ?Yfd4OH9@aU&R2eTad@>G2[EL59HYGPRH3LZ&H
1WDX(XWA&98HZEKbJ+A^-D^Va?P.=1:HQEIJK()X.VYZ?#=d[8=2Z5PKBP6Q7ga)
/&61\bTEER3KF@/UTR]X-QcE-5V__3SXQFJ5#_\6cJB1,J>LJ8XCR0F=VK)9/8R.
A9fOEU,INXCT9U8SDE7X2D8M718E/JIg)2M\N\80A:[a;E,.dY2_UZI&eI1?XE&/
L]]?7+=IBfL(-d:FFROR@:Vc9QHIdG.I@0/(V?UZc.Vf[7YeOX.SUYH,L-bM+KZ-
VQ\)]64e6Q;WQOb@fI2P(C&=B?&O2UE(AdLGS(D96G5F94KXdb&b7,M2K[PUHAc=
b(b#2H:6ZO&FAL9X/Zc92[99&@NK:ZgTbR+/]8.&A0<UM(KV0&6/07YZJS(:&_YR
A030bS@BM^8HFN9+)(7Bfc&]\2aP2OMb#VeWOcZIbTJE-Ud,97<#KPdF-;Y@3<JS
33?4#BU+-&YP:2,TMFOSJ@C[UdF?f(Ic?@<H@SK)?\)d)cP\F.)L\:>HL0^Fg&_7
02[2gY@7<#eUS]OS9NI7YRMU:W0GQG6A,(>XU/a.@g@-V@ER(15ZR.K&\Z=e&62X
@L.KNQ<CO=e+cTLPQJ299;WcISOHXVT=,85=I0WAJOX&EW<XQ48S>8(ad+-7(4L^
g0/1H&.._\H&OI=\A(7^MJ8.F6^:<dBIF#8c[\B<+S4(cV,Wd1e5HBBU6[6V?BCP
X&LHB4>S:;?b8M)#g:F7M5EB+]b2HO92I)L98@5c9U;,CLM=Y=7a2K][^:&aCTd3
0/5e\69XfEWLF#,M;.1YZQ?XTdP2@X^0aE=K4(aRCF)4>SP>32[N(J[LN8V?RZH;
^g5]25I4E8_[M:Yd).=#f;^.QISJI?XELB=FF<:XKg[Be85d\Ib;LZ;)f6fD.?3=
5=(08ef?N=C4[&<bf?+I\)7+]XeI+IS?,5O@VVe;_8aVD.47F5K^FC9ZUT?OLD)c
fVUYVDQb@LV/<&)CMF)F/9HVZJZO3GQQ\[a)_R3@[d7J^>FC/WVS(Ggd2I1[XWCS
0-MD:XQgJDfI/IWYe>4dQ_bbNPIBEA8D@bLg45)e>Q)a+O2MQG,993?Z6/(NKaOf
\EOV6AD1e.ZbTCg_]K>HKd/DWa6D=(ERINX-Xc1C>481_SfX-5^3Q&/7a#ZUSGWg
6+0QCR\=@ge@ME4=3(SZGR^#b.,eW,XX<[=0GK_UEF\RaQWBe-4XUeZ[+\;eN&cd
W4B@89AWWR]g,)FK:BG@R;A7^d,-8+J6FagJ:JZ7FV0H;ZbSA_)MBR@NPG/2<D^)
83K1HGbQ_(..I49EK9GSGM.\f,J+aG?K+Y]_aK)ZeF(-]:OFZPV:+\&WcdI3KM^(
2fV/>S.MSa/cSdQ,MDR+cASKCd,#ffN(H\#g]1]52g#2PZ/&BDI_>2M(=R+Z8?=4
\E>@,C60Z:4#H\5WP&X))e.>[1D)5QZ)4<IOK9Bg7,=G9,^Z875IbeJJ;Z1M>-F&
[;3Wc]9UM?(G>OgGW+MER_:B0^N8W:DE2]<c,K.efEa\-?c,FWKK(Q4N)WS#:RH.
?G;5Y5JVNc5d:13YB(gM)2=_30gQ0Z026P&27Af8CB+93(RZYfd#U#G3==(g\\JE
:L)^A3\\UdLJ;1E?#eT>(6aDDUE)XF2.0&P/b:gNIM,,cLUfV6/1.^6?K/BU4d6,
K&5\#_XJHLZJ<@O7QK=SJ;L+MP]IWI5Dc(4&WV_,^ba&^2WH4Z90OP[cFG<[;cV@
gTZHcK,64T;(J)5Q)FPN@W7Lc^:=0_>4TJ?gf+H=/?AP08<8,QHgKL96#?c@MVUE
0Y/JV^Fc1[>Z4_9fR=+_T&TV8&3XOb6F?8ZJXS;F34GT&VRS)gW2,#F@HdTU\,-Q
QeZHNC8;-Gcc,[e3:AC__GCgNP:CKP[I3V:DIG;BXA@DHKZ_fdY6-Og@FR]?=-6,
V9)[>c6@]adYJTc@UP[GZ;.^N?:&29R>\.8S[ea(V@0.3GLCfbJ;H+W5Zc<GQcDH
<AAZ@6YI]86/4W(SIOHAf(3?f0MK^QS?99>=e\YXKe;^7?\#@1:Pb[^YE@UVVHO/
HK6E)JWBS07D@=K\^2M^UVRYQb(3T7V5.&?MBCNcXO9>^_>a(c@SM87Af\24@b1\
8MEc#XD<[#TCXC[3K)R[gcU3Q@P3\;<5QB9:AgHHNW)E3Q=QagBAW-.e\ZXJKa@D
^e:DOS/J@[2/>f#7PY..M1W-MI&BWP#.@U_1LdcNKbCRLS./[V8&L#9KOQV@YI57
8:VT9LeHaa7K4fS?)D-c8>-UGMYeXH/?WSH[4H9-ZaY?:P,4U+H/VL;EL>FS\9(V
<<,-SUK=GgS1;:4L]Ic?B0/a.=e&GAA1IcdHU&0^D9Y3,O-K#EAIcXa6MXN/GW+R
0&EL1MSf?:V1P6D=\_dFb>QJ,_#)[IIEZ/LD3QO18#M?<S<N<JRJ@#A\X_)fe?_K
P&7N/@YWce4aaOd]-YF+AA:9G@0IU_Q2R(1+(V/)QdI9ZOcA+)FHXY&)D50&.eU>
RFPX@(Y/R?J>3;-Y/)S.YgUOSN7WbJ,D)8FVJ:HedC)M>\^?AfUE_\P5b4cf@bN/
eIf_EgK7MUB41Ma;#X=L_KSMG10UODT7DH<V47AXg/)D[R\D#+GaQ&E,43^ccBST
;a@e=7dE.XE,JQ=OeOa<cQ9IJEAE8&3D^EM.8VFRR=<[9ab/=QM^TOK4EE^d\X8,
#YIGL?5c)_.L-:b])[[FBBT/F64d.NNBQV>eDa37&\_#=HRT1ZV0K)TNLSJFbOH9
5bcaV[@N525NQO0?NI3,5.DAVR-f+9;f3f;FY2V,P#e:I=^L@@T@QLR7JN&&S+&R
dBVV2;a4^JWg=[U-;9A_D]+LL2J42:+1RLV&I>W:<O6NE;KSe^KZ33acg(OCAgG.
59D8d:O164(:.&@bFDKLL]2./^gRD\@[?GKeM&5DgCC&_A1c]?.6?F/Kcg[>e\0\
:AC,Uc4Q5dcNTLC[+NaS@f?QfE5^R,IC/3BD?O_FGF9-+gE9U5#X^CDF&7c<faPU
G<)QKY/?>[8VdU?7_+E^L41_H\N/:<3KB,a-P.XDP+2HG>5F^PNI)+(GVE5d9ac-
@RdJ1?M\0bKfF-=dPG5Gb[)-g_\WKGMe(Ob]+Y(WO#N3&Gc?.(B^E&:QZ2_Da9\[
+#f2TXY[Od=[Oa;MD#^D/+9?P;UWM=[P?V1,X>b_YLc(6TP;U0P7Ka8Uf=X2E6aB
8.4aY5UcS8X20Fd2b8M\0>BHa:_(724AVf7RKJ9H8ACVCd_-KWDF7X7(JSMCKK59
g_W^4e82adJOQTV88Q4CE9GId;4GK^?S(6MUT-Z#U/FK.W4#KYe;?EYR&dAOL#;=
&PeL)V433Rg0KJ0CbEQQ_7MH)Yb>dEPZ;J(J7X9dV@GLaaH:O0-]N_<4gPZHS:+:
?)E,Pa8-^[&QRJCR>f[aRT[<0LJO+PEdU&GfC._3JHQ;VZB6TdS>1YHEg&CLJ&Ma
begd4TQ&@UZS2-ZG,6>3,ZTT]U1;eeC\VcScGU/+Zf#Hg[C(\C>_#DB[H59XAF8T
]:H;]\fDbag#d;=ALSAe3ISeTQA9f[/cC@=C8BUDVRPf5/;ZFJ1@3MddYD4<,\Y?
=R#b+8TI\g5M8DOR:B.-;C<9)ef[g^+5ZTc?][FH^/I^7ZIe6>79DC7/;Zg9\8?I
K.>Y/F>@FCg@(daKf0abC6H=E#(\1&#3e?\E5<I_A[9)OcdfN&>931@a<-ec0bS5
@4&#Z,g/Td(+[6?CE),J-gVY;RH??fB72;?W(,4g9Xg+#)aJ0H<+abb\b8G?D8EL
C.C5=7OHS>ZU^1Z6EYMS:1I<PGe[d3F70d1f>Sg=5:W<]JYUgQQ6DHWPL44fWFbM
C9X+?@)9&MVf)I68Y(G9AHd#WWA7Tf4AdOgY^/YK\U69-5JD]VKC7AN7>UPbT_a1
(S#T_7d;e+d;NHC4LIM(-]O8R0ZJ_fYIOL1@,cNgC\KG:O9=;e.NQbH,;U<fbOS4
_g_FTSU)U_AB/I(,gG>/M2J]C<SH]+PNNPd]fFf@\H,3PP-W7P4-^0J\1:d?2]Z)
7KHR>d74S=8X7)#ITY6=CLJK:=3T]?+D6WL),VK3egAb86A[#N=,T7I/,;_3SR;e
;\WYL&]^XAKC/6PQ?C[29E+YKCC7TKO:,Z<NE08EJ>#7dL:]0[=WSC_1H6#5HQOO
6U.T1IY0dOJ@WST8K&N2H[c3];\c:aP@be_J49D&#2;+6J&<_gbTKJfU[H#cJF]6
5P2DT+@d5;31DeL+VAH5N^+f@1c-G-7ggCN<<:;X,3d640FR]JM0,(T0W&/EYO3d
.R:dKI+[OU.8_Dbe5U+cV2G-BUcAeOKWRIOg231U-()I7<A[_P)/5SDC\QP)P9&e
d?,bV+-(_d;^R+f@I6BG1KZ\9X1f(+\e;6>=YP;Q)b77G5)HX^[^,.VZXW8@_Oc<
(S@Ve[aK@T3Qf1W^;-fG^6F[aP=g=+28f9GHOYC\)#+@g8CK3D:9=g^1WG.N)Pc5
T)1UNO6Of8ORaKE22-6:W2RHc#9]O6aD<^#@0RC94@HY,FX,T46PaU2:6T.g6A5)
d1:AWI-g+\8fc@>)8ZFM[B,QZT9.62e8VA\/33bU;,P/bHg,NeSI19O-1)M57<@O
IZLL^PA]EEL)9#MT9QY1;O60-48TI7V25M/LC_)TTX-Id;]TKc_8BV8CgA5HJZYO
/Ed^X+)AK:=Z<f:Z]0X^1aAS=JZ3=^>b&;;OU\50F#,><,FCXSf+EEfZ7\1=0IPb
H(5O2c(=H;]S9EF5aY1YJ:KNV\FFA6aFdX1/?Ee[=C/,H3Eb7aB-_c-H,Q#U->>3
cX>D4=ff>IHRUXZ5]QcgK1?dg67OU:6]22=D8PF+?PEH3,SE8Q6gF@#2J/LJ/7QP
F#UF+a/7b0W@)35;5B_B:Y0]<NND<DDFYY0,8g7;:Y:DgXFea9VPaa]/WB<VK#LI
BF6b05g;eU];&&88VJSQI+Nc9(XVO)YG/CVb80Ja@3f,:Zc7F::>_<6H:U6/9D5E
#OP3K.Z-V:I?3L/@RZ</\cD57Y5VCA3_(VL[cVY@O2A5gL/..0[^33(__gQ/A,/b
abFWd,;;I]I-:4Idfg/9F8W_>^6a6-F1MLHUGd]+M:1.\aXK[b3-,gBcI=ZADW[-
4a.UDcW/J\VM_OJKO;+.DW;_d_)[SV:8<B(N7^a<226JW9T[c;@@+bO>N)@-N/5@
([0]5]#-:cQ78(@-[2a81^]E-e6L>+eCTD&HZW()BG?WH/98;\+-KgaA8-DNUcC]
TNc?#+I^Gd5.@FC4&A^d0:0\;@L;faIg=GQg))c3eEI:e7X95/K9&?TADSV>fWA?
T<[cS0f5U8GA^:MLCW]g@8QL5PdDff<B5R&)D=ZBO)[g0dR7Q(CgP#DQefd88]Xe
_fJCb2\Ma1>(8XXD)AOXLWf(=eeF;ETgF54DLAc2BFSd([E=T0^A\OA,Q1?/CDKe
Q\-=fU5LaE?=54_-A5B)-LH:aQbOGVUg]T=].-7T>)8:R8P2VAPK[fAX^1\;f?DD
H(&CZOUP2\]Va-?G#8&X8G+NFf?6dH^/)0G:53UJ)?-OED<^HJ_8[KR6]()-(@gf
=.+Q4-D+d,c#,^7d()YD@QWcd+620AF^EUA<8-EIQF1V3MYZO,T<NXRL0dOIN3GW
1=/:4>E+dNYdARcY6TP)CE45aF[^Q;GaSC)NPSG4&4DV\gN+3VZBX2^).=^7Ff)\
3K\DL5(?PPDC^ZH@(@X/Xc\-&N\aUKbcIaNBL3]8PK5>(b;?,S:FD)6Q.)P]W2FQ
.B14eQb2@WgH=0R2g[P7@gVAUY2)JgNXI.56E&eTQ[GbF6BU#f_g\Lf:-)4c8]O4
d.CKKc).NVS=f.aZR6D_DK4NDPW+f4H>\7d0)If6g)V)1(WWXR5,?H?JIOM>fI,M
\Le/H\O##G=FcBLa[S;P0c_,&^7OfIXgTfFa0,TAM5S;V,U?eE<#.B;OgO6[Qf?g
C#Web,M-<^3<5Y47>ST7P8<^dZWG>[JaJ:)OH)aLK2@[T:8HY_L<;6g:HKaOe2Q^
]X6c/b@+IKOA<[L,B#-6X#2d53-#1_7=_XOe:U55I6CV)RJ6\@fDB>?N(B0e]./C
JC>.1M4=]?G\TOd<R^[H=34#4)F(+D4:451-QRXQ2N<[=);<A,+1<2-<d/Da[I;Q
>0&eG45_2b/&#1Sa?J^D:U@Oc6F<SNgP-Y(e&b?HAD[E[I<(6VZ4\_@+HaJ+YHHI
<5>+^GBM1>P-\.JG#f#]Id438J+2gf(abW2fJ.6655<P:G=Ha(P@6CfAOLf-.KaP
RN>F\fe]0+1:>_7GYHE6>[90dJ4&4PB.;9P]dN&2Y:-)Q/F/6F4,W\Oe@PZ7RL.C
^KVSR):)6<OfC+cA2H;COMfI>f;VE8becK2BK0T152(gW(A)cC3T:8<8[<c(IV3-
MVQW9/_Of#)-67^2GE2.Z/^(?4T0YJI/HH>M^#JTXMgVPNa5^E,2]cUN<0PW_:5L
CeG0Fg.HJ=H1V,P1:DgTXFN.1EM;AV-f)e<DB;d4F0VP7dMDgHO[S7J7B&TE2c=Q
,07fM?4-U[b8+<P_6+Q6Fg>^:2g=8;]_9ObN&1gf>KDL@U=^.#R7I>STBgR+(((B
5IBP1aOVLFR3P+EQ1b<=OTBbbN=O9GIR:Rf7,A^7g/^Rb.a.4[4,4ZO&OH.J]\>&
c2?J;d-@O8RVeE4LUa/[QPSN@+fSK5XV\(6SCO1+I\QNH)6JSM]1WFPE.#PQ.6IP
@3#-WcNObSL)^2NdV0FP/Ydg(VXIS+Ag0c]^KU]Q;F8e#0G.A:ID48]>>9NXCEJ_
UT7/&\bXfBU(gH3&@cQUg#UBE(Y/]4/5fgV2+H\@.9KfgW^RL<H&\gMcTbg0IIO(
#af;A\VRS]G=[<3,?K6d3g,9M(#W\5NcMY?OW<&M@1J_X^ggNg=G:[X]S6M+:SVD
>8-V;+KKP(Q?H3H[2V,[>/E.,OO+6]1@/MZa1W>\_9_NIDXJ,W0,QQX#6Ua7,LUC
g(VOZd_N59,-7#K?eRG=1H8DMC1690&E0g.G3a0_CJG@R:dQTCbX1?ZGPWFb?;-d
UW0I+>E@C0QQ,M6M3:Jb4?1,7RN7c)g[>BVdM^Rf8F8&C0H<<\K[^N4FCGQBXTH2
OHgV+.Z;8AOOeROO[38ID7/6Y:L.Y#E37F5bdRb8g\+fY3a:V=&L,>2)\c\G++^P
=^-^+?eLMebg?DU^[RCc&I^8U9g,B-_^X1R8W=FSD-&6\C0ZRKEf5ALRPf,a?KcH
>eSZPDQDXD&:0(]LM\g#2I=DZWWD<B?Z94+eS3,ZJ=BHOXN[UE)3aEK9-Z98^4?#
V5&O/NFe^3]g:>);OVI-^JJ(5(]NL.aW0C\[FQSSSTZ@_E_(Z>WbE/V+-OEHC(RX
IDRF)Ig4+M7MP9WXB]G)-H1OPA.^fKd6PU9;66a?QTG>SXT7VN2SX1]aDK<#\Z;G
IF]I--?HZAK021cT-cAeE.2Q/TX&4Gc-f\E+0a)^1RXL/]OO-f@K<(SO[=,Ygd60
_&W_6:388^7()/F]@LXLdJ_.g_S]gcS2_F\6NLBO^4/F]ffIM<_7<+O]NbBM82,f
Q_7:^25F^.S-U4+a6?LY^E^@NS+P]8XYY&U347=WW6Z[7K7b-ONJP#8@>[DHcL\O
EAAdP\E68:^:-?8fEZI^@f#]?[TG19:;)XgBT),F1@FAY@6]111YGGBED+H&O8(Q
>@ZfC>3UMV5,^Eac(YXYeY5:bg6[/[CS[@C031^JGQE>D4gKO>=:CgO0fbP3<=1J
b((42Z379\JR.5Ug[dB4L-ZgF;@\5>R))LKF/F#=\WAL-P?SHe</WB:>dSFKY_SX
&GFT3OC<=LXWfXL_eQV=&BD4LaT_5^+QO0E&J5-5-BA]0e9M^<OfX3;_YS?LS4>A
TEccYI11JK=<SHc+e-REO;?(-)Qb6[(b^8)G[4LS#::)b=P-QQJeFIRY)06B]PG[
NQJBI.FE;8)-3f3:a?XY-4[53bJbN_YGR92A<T3DJ^J;.g8g],_;N&-]JXPZL^N3
=V#=_?/Da=7@Q4]EV9VE3b.A4YV:AK<YWG\1C[FTd4N.+XD1AdF\5ABOc9@(\&L)
^KXTM4<ZZ=ESXFJ@QAXaNGU@[EeDH8F@a<^#)AJ&\:C]SA+,_Z8O3-&gBf:8ddXB
A@S-75bH193-JK,P#M9W#F2IU?);\#[IN/b^5Q>?I(2<a?eaCBVH5Y_/::F):Rdg
3U2-,32#X=U:\fUIZeJ(&0g[Yd+@+H(f[gL&XU(Kda3B?&J+W;DH=ffS:^D:N)W/
fRT@>#cD6A?&X1;7]5PdLS<-IB>[,SHXaI,6[Q+1ABL0A,@:bSDb;a7B0=T9FXc2
TLS2H@5f04;b5&A,WN+DcQS)N]9HB=5SO9LYR6B<.&B3,,,1HM^R==Z8H&J=.J,/
EWN#?dHSa?8PabXXaOJI,231JbV+DcPD5VD6,&#\[;B,c>9]Bd1-;]MZ96ZD\MP\
^>fN0g:++?]Z:GFcS6eB-VO_\1aYb+<@GdFK\L+S\=,=ADCVPXd<<IR#cG/4+b?(
YDc[5D;QG:8XZfgUfV[(Pc>:5/BH2ec<X.@1A:5&fO[7MEKB3SPF#[XF1/9[+X-U
&Da.MFS,8c0,@)(dbE]ZSMaaJd2<Y5U_D0/VfKOc]8FI9D)._5\K90Q51:.]IR]/
^e4:c6S/EN^VQ4<&I?M\9R:&#1,NS,CgA,OfLZ/LJgcD[W3a?0U&_P:E:BE(GTGc
?XUg]N&@:OSPdW[\3BVP]_ZSL8G_D4R9D@W-J4+O58#EU@W9R9E^D9Vg.HIH2ZD>
K+GY.<d-R+TB8bOU>-V8JMD/=1+6GIFLFZ+/W0HO9YWZTQ.[,F>6,-c+=UT5aA=N
58Y1I:(XB/I#Q3]?e<@MB36<J=:?]K7&^4V[PHN4E=V7V)5L7(^+gGg[(d1b/,#9
C)-eA8NL]QZN>PB(^c5TUU)S\4695JJVRdR<e6Y0O9P3W=9HXMd1A&Pf8GN4NTKg
C40/<7^M@+5T46/I82RPRPaNa-23-><D9S/L-2NK>#Y[E8Z/GY3@Xbb[dDb&,PeU
K5R?HEP;31-QC[fEEEEQOKCHMdNGb&<\FR^L48UD<7[Y]W?>#cW@6ARUeIPW?6YV
[_g>SWSRcRa[[<)a=YTB[U,-0IGTO--.]bB:O6HNTR846d&=;FeI>])>6Sa>)TbI
B3_(X(2CHZKO)JDK#=>G+^E-JZe(aVfCd2>.)6/JZV1LO)33(S7P[#RZF&0>H5>H
Cg:DXJ90&PH+.X(#NIY(W6SdYEcC_0@@VI@N;P+1A#+XJ5^DZ\&Ef@)Qd9<Ud4+c
fM=,G1>_=c_f\<gNRG3aag/MZ>[A;F_2X.)dPBNIX0.B;dJ&LaA5J.-G.T2g1D<@
FM(b^[)=?>O]aBH71R]>N0[PW5NS&Te&-?E?DPAU;2B4OO/7LEID^IHGY&f)US:J
;<Z1130I_L[KXUFNGBHH:Nd3]\9S6NF1Ya2KNA,8aX13(]<\KNV@XHVgX7[8(BWW
6-4VSM]=(OG)F9B].?JB?7G^NDF>d>Y(NdgKI+O@X>a;ccc>LP)=C#G1>9G.Fe11
H&T576R6HR=4R>eV:_3b5XYHO^#)R6/>^.R45]59Hc8;8fHUZ^cZM)1?aOT2QU;<
+FGIFc6Sb#]U[HNN&AOg;a<[.(,_0UeCWa+>\;PETe5ae-dd.Z>=P)ec^S#RA;?I
Zc,RZ@PMU=-HI7>R,DPb6R0ZQHPB;@AY7#<B.V2\+dAeA/2Vf0#b1QIfD^H9G76S
(Y&Qa^FJ<&dNW6@CeBM(\??A)6^<e+:U>&GZ=fKC:I\]R>Z?BeKS2-UFNS8J30Zd
=CeY+8&2^;D,a89R7(I&Fb\Ec7(&CRd8_S+@.?2deb08NRJ.[UC-J?_A@^^M-0Y[
.B>;5#6V:&2eMIa-4FT(L+>V9(f4=4:I9CI,f8Q96-5L\K8I&]T]QE=U1YQ:87<^
9@^GX;dP(R7#e)2X=SC.4Fe9[G9#_(UGPfZ=gNR/Qg5&3)Vd^O1/S#^KcHL7UL3=
FBe2(U0&:0@YP=eM@J=<(0c)+aA@7EAQ<I9.V6HX]X?XRG97B#Tf1M/;622cL&EM
c9M;P[T5/@Ug)N=WY:/0QS55.:_JgQ-<S+f&#5T[gH\^T4B<G6f7f)g6A?-.BNDK
4N^(D)#]a1U12D=UC@dDVW&WWdCPEPBZ\II+g;K?0f=CaB6c0=NZE@-<R9UAX+C#
@U3+RPV,#g-R5F741O2PR[7,#)Nb(:8NVY?W6VC0=SF1MHe]@<456UY7C.B-915:
#f1,[)M^?IKDfF[XeM[(E]LFQaRATf+500)YLML_1C.N#\V=;LT+3^[4G7#7Q_Y-
CH)XTDC#Tgc)MO&&EEBU3X#&]S(_d=:BP24,N^B4A2B<HH7+eJ9531V1>3\YV&&L
)=&dOX/<KbDS/R;N\[@P,A/2.b,V7IO(:Ga5F?J518B,]T&?0((39E+MJ2S8(JDa
B9bb>D>+f_g7,-M21Mb,87Bf3STZDLNEIIUU0\B?#He)JbP1DQK=+[XPGF-6#edH
TO5=7EGF,#65-VGMY-#2@L_/a.eOd3-V9OGHb&T<-9FM6b(f\IQ:+JC#RK@#7bg3
V]UgDHZZD>F70S.7XQ<056c==b1&X[NB4]Q98,gB<04A>>>0I/VgTR&4&:+M9,DL
RbQ2Zf3J@^egQCM5e6XN4,<c[415>/QE&@J_T-P]/1:_K)?6GC:O7fG8/MZX(?&/
1[<L2R-=)(MUI[:fe>D4J>DT7@VE8_/9DOG-A.MO/aN>Z:TG?P;T&Qe_(0Q3P,QG
J./#=7D&CbF^2NCN(KFR^1]eK:AadgE7UT/@=6-Q0#IKHP.b@T,ab#&RAS>bgDYP
U#2LKP+R,:U#(ef<U:LRa.KIYcMK]Me2DDX6fS@c,0/7(_MSVV.Zg-+_7U)D\6:A
.7d1f-eBHO9^+@#M-[^D^;CTE]X4B.Qe9P<g15SXI9@AeZ_VOC8gb)4gcg#]A0Y2
,-8)]6g#PM&_G06OCZ[e8UL,N][]>7&V96#H#TU_Z2/(A#aLM+SB1e0>f++BUYV?
45b4e<0:.:N^7EN,Q);WYBD84:3ET=Y+b1_b]C-R4M+T.M[DB4FM;4WW7TMPWfQM
fCdQHSHFeV;NLVI6EOX6.P<(=K@:1B<aScQSaI^OTHA9Sb<3b=@cGTfY.=Cf.d4]
UJg8LMa#GO>Fb+gC;+?#AY<@6&)6AAA43JS0UM.=U-=(=QPZN&:WQ<b@/4#,01cO
+I674.KU(2aI,\4HPCMJB9ECKT8(4^P?#bD94#PQ5N7=#6@BUZR#@_-Q2]S\:Rb)
>SdeB20TPX_4Nd=M)>3QS)J#LY/3K?WZJfD1=FA^gA=,(XQ/2_([:)4MAEGa/@)Q
bHO^112)ROZ;G?04#\#QWP7HIfJJ=D48SHL#BD>.,fcC?]HQ8[JDDS9.Y7;)g_?7
CH(\&g1cD[XD#:6Y<Y?W5#A?#MU;KN/PG8fUI)Z?E0Q&NSUR/^[^2SDbLQgWO\.@
QRNDBG7?X><UTB5<A#\bfGSWN?8420E:LD:[_:VdJ.Q/],Q<-Vc7YPU]_@?IJ0/+
SV#)fA+VW9DNZS,\#/;4c?]?BL<Y+VS\#_R<V_.:[R6(cJ9VXeV3K?OF9U<CAfJc
0@P4N\A^,=@fKV.Bg(HY>>BG)DC.c--.FbV<HOg6R#a0ULCYN/MZ)NNKK(H=Ua.Q
_c<?VE&XSLKQ-7EC?A0_?:0\KFKG?_4-c#X0BSEZOM5@BQ9EaMDf<fWL=ZR6&:0&
[RZXf:[D^H2P[JBf3SSY#^B?bW0cd\]Sc#/bE.XAMH5a3#+;FT<gHMY35FB9_]_,
C^e>_UdT7)E+P(^2Dd;73&>=6HWcW(DQJ_:)Pe#DRSKE<f\/e;^#PH7VBA,(@IT.
=0/e7O7OV9);0b37e_Sb@WAC&Ia?Z/,K>MG5DM]f53>c3ZK\/.+[#5AVXLT@>XDe
#73F3V]EEVEH1+de#Q\<@e:Sa[Z&GM-L]dW\.F7bgeD;^9G:CC:/H0].?5==(_Sg
g/fgZE(,bC&ecc?]MHPf252N+SS6YS&L@[4+1^3aJ4&^J#I@OXcf[KbZNVDKa8.6
=\#Ma9AS<-L/(,fRC?Q?3(I&BQCeD?=R;N:NbP:S@23DT1P5=-6fVC<(d#2fT,>I
VZ6d;51VRHOVf[Rb<>1RSY=9g3T1Y#cTbU?B_IQbE.WJU-&8I=+(VN.>MKA1^Ad\
=3Y5S9PH\H=2#KGeRC;\8&]/Ta3K[Y-6P^U5E],(7[WV#:?,e,J^LZf;-U3dOD)\
a9F4>ZcW/HF7WPM><eg]DH/SaRbMJeA.ZR8OWLYV&L&7<LE(Ib]^&J@I-3D&BPS?
7eQFEe1gK6F[fGA5CUWVgO),,G,IROf\/^U4-WZSTDd_Gf_U13Rc]UUfK?Id2<=D
@=99(&F/30X@/?HG?Tg#8a+O^J:/V033B()Wg4,g:f,X1Vc6T<QH6QP[ETBfG2LC
B(1HO]\ObE5?cR+;WP,P\SWAAS1A5+1AUD0@0S(gcP?O90SBMNd3&)MH[[/fX4@a
G;CE8YF/@gJ(-\-?\<&J(f1BFWbS?EdI-8e,GUP^#CRbeJB=b)[NVTS=8@fS23S5
KWcV^XIS/C/I9RX4MA;FBL.5B4@aQbASFV>0L(;4(2+)>9)W?2R:(L;cML;@^0F\
A1Ec31&7A)(U1X0RdO#@>MPOR9YGR<JB@:]cA02X=(&)R6:<Y0C2HO:ZX1>^LSGO
WX7C6QXC3L<IS&)QRbe0)fJ@e(,d4;OS>:R(bgZQG4QbLe-SD?ScHAEfa71@HKQC
I/Y]f2]8M9T=a;1dISWS/cGa1e++B;Ic(=9^e?>H\^1+A8?eEJD,4X_K=[UZ3&;<
gI7R[,3R(F]JRL;@f^VP?2Nd&2]3a5#WD);81CBUN42Y2cV.KRU2N0XDODIMc-9&
[1;RJYVKd3N[RcMP+:B1QWc;/\:DcY:K;IRac;E/:6@4-KP-:UcIXYH61C_>F_7-
fK3;8aS]54=HffLN07MM0>\f7837.)G(&=-2QTIa8VQ^K^T4;+;#?,CPMT_S[9[D
XWg_CQ+\YD[O;:6#PF#RH@0[_FEc.[BdJ)NNQWgNJW<2OT-f8-ULC&W5IC?B;YV6
f?M;V1?H5ASN2,(]#-afbII>+7Q8[ZJ\]B:G3J_5TT]eCYfSN2/8QUF5.<6P>E<K
[6gb80#[egAU<HVN#[0I.LVA3K.=cQWC8fO<22T\MA.ZXBE=1BG4YSFY:b41/EdY
:8Y2Y>gVLeQND6O,MCY_6b^,U.0Zg4N6[7JHRgQT_#_[?Z6P\5Q+)Se8bZ(-ST58
N-7X0(\,RfF@XT7:/6M\7Hc@G)DB++P++\aA#@B9;/K:)TfXI(2#@G/SBBa.VGNV
D:A]3g7L:IXQW>32GW_F]ed?X0P_7QUeLE-Aa\bUc-9b3e6Y,Y>;KKCJIZLMV=[d
.O63OWA<[g/XfBbH/5\PeN;#C)eO5^d8?NVU47^LKdCfN_Ag0,(8V/2L0d]F^M95
TR1RY<C0.^6]/Z4U[_V9S:VU.(IS&&^gZg(I=0HU,+^ebV:JIJHg0N^0>F,SOV2c
1&3.bOA)U;+TZ;;8cW5+>=-VQ6P3=W[V1f-C6H+UDdf<6Q:A2J9P0IK.^fT5(P]X
QN-bZ<?W.+V2ec[EWWd-92ea\<0eUPNgd.21J.2b.0:]#+&Q@HLX_=Hcc>_Ke;4B
AM<4;;9eNA5A3K)3:\OR]S3Fg&9GXD[A,0-HTU-9]P[aJ6?&_#c\I9F/V@5PVP[1
(+4RMTENf#V(6U?J+/O7R-UOW@(JD7BJb+I/H_&#E]#U&\H/g_3)bbESfM3eVW_b
[L<eR\Q<)&ABeC2AS_^PfFW(M5d[]<^+4-8aa@=0^6;Cf?#WQNL#13DS,Wd9_>T;
>6CX]d[F2)62@PR]ECf&_6N@V3-M2Nb)2(KHd55S&BH>_]A)Hb)7_Og,>K^-8UT@
CgO3KLHE9MXN+Qc]>_H=4FC3fR/XNYa@fJ6/Mb?46Ca\P@/&6FL9T_;_LZ/HNIM]
4Z/LF8&D:<0M@4E]:16)&GbUO,[.cTB(SE80FM6;da<9B^1_H-:6[^1eR?d6X7TP
d4?g88IXc:G[F:U)M4?H#U[APGBQ3E\6KG7N</08:U@27H[/@[W\F>/7#-gFX4]_
).#ULM)=MGK1BO-?B^4G7aY,XAREV37Xf])LfP;FQWfN4[4Q2[?+QR@H#]X?T_Qf
9,\QEfE<-LUad_^+UE4fb:XG+4e,=gXV0U2^d71;W6120HdW84c7<V>.P;G9Tc=f
9.OUeV;6UdDEH9g__-PK+628PNCSE46:ec0dZ2[)F3B8#[7P[O5^G44Y>OC)(e9D
:4:96&G?4&,U2V]\T80/(IM]<:=Q-Y2_\([7DPP_FLSLF90IQC^#&bBd_c=UgD:X
/(=FB.O2PG<,1DVXR\9)H95KJcNc<CUP0[P/RD:\/P3HGUY([d-Ja?G)AC#@2)Q6
QgU@S\IV>ec74#QNNA;;#G478ZVTERW3QMef0/A./ODG+dM>bPVL[UX6O[I5WS&B
I9?IA29DdU?-EZ_A[):AYG8;:)&Y8/SM+U@S7VZ=DJb7T@@&&E1@^,SB?-/D5C16
^T9(/MHg[;;FaY>K[?#R@H1\1<M6>^-24V8Y+<^\P\JT<4P=I>]ETa@&;d=g@_Cb
C\-P<V#.RcPe\N:3fMgGWF+H]R-2I@]7[bVZMY&(>(@9.DZ9e9R,fIT&FZ5X+]NZ
3@=]#eQAI\dNFVL4).Tbc8]F11@2)^Yf(_]XVA[O_CG-13C=gGBGZfa1&.g#-:C-
J]+aH#RHSf,M_XVTf#U.)WNaMYBYPI4YBZM;F4fe.GLe9=6+A5P[2B#XTT.XWc1+
2a-4-FM>@24LGdA)DTIMLaRbIO8H,CLD5g]9-XLaK.WYJE:;g??4\C/1.8dV+c]d
Y3RP2SeK1/S6<P]P@(-Z(1dd<-;GaV>9D_I^#?KH-cDRaDO/e[NTJ3Ia@RZWC]K^
2+eQA>7;:+;&FU-_gaK=.@OD_---dK?R(<Zc3]TYW=3C@Q;GVSXT]g5@\+Y=DQ]R
Y2#+8]&8.:PC.?]<c>M\95@YP)1@B8FC>8T<HSCfHE9]PAEe-G?FKR/H6NJdJ=<?
L4DL;KA0aIKX3GSEAX68OOXgAU::1Y@F]SQ#UX4A+e\&f[MULRNQGd60Z)T)8)@<
4)ZC&#TgTdXSf]=892?:O@,8&D?]5a;0Gb#CFII]YM<-Q)V<@YI#YOH2XfH8:#]3
fGBbd^7_19VV2@=<a4<a1(<W>YJ09/e^5WcM8&GHP=S@NAN)B<YX6J<+,P^d.I@[
C^C5fcTA37fWKF53<IJe+OPe#aKF4Id2Ae4Md]^NDH9O=2SRJ-V^XTN&_#(&][LV
c]M:<)XLD)>eK;?LM@\ZFf;c70J49/VW\Ge4.fH-[SZR3<->LXNQdP#LE_\,70c=
](0d<H(,(ZEe]XB9M&+V+YHT_5F,aYAUER\\EA9EY[.=2VW&6Ge/&S^2fg#+@N7\
bGTE<C8RP2_/=6_gA)N1XCS+D3_F[P0HYM/+_0ML-Z^]Y)cS]TcOZAAe(&VY5TI7
+\J_BY6B</MdPJJ,O7c;.A#QRDRd+e<R\Wde&OecOKb66Q#e[?KQHgS8#:RFE>:W
_IF\S]?(#=MHWdRE@>PGV=:-PE&S:QgRL4WI];=>1&V7N-N;555d+OX?gC<R-5BI
R.FWE.I&cO_WOcCTU<9OKSB>?2HI#?@d(;D<Y#7eZab<5:&/+D:1I8R;+8d^V;0-
cAdg+K_,\cRHF;Y(RQ5=J#GGda:6H)QG9^9Ad\O+RU)73&ZRM:FdG]UbQ[9]3B4f
/&R^R7WX/>fO@6]5E\]VBEH05We;XH-f@A,SS2U-.53N6<I3QV7RQ&YFNcG.+?Q9
2+AXSL@f;NfY,BC<ZM3<H5/)Zd+VY/.6)>:P&7ce#<Ab.cKGHO/,S.>R]I7O_:)Y
84-&6;JU@#V#38K;gL&C>a22dTHQ@2PNL=+]_]8N0Q\@XPAP9SUc3a6gEPJ5<\(_
[2NN,D\V^RHI.--65IQE;G<FX44#0J./OCDdC(5BdM9RZ4/dUL=e,,(1+\KOJFKR
2SA]U:Pa@OWG24?9&IF^ZZe1+,=3Y_Y(29V9:De^-&QV1C+^A;EaV(Id_;EWT?c,
+fd5@O,K-R]OS5A8^A\3X,Pa)4[+B^OPT8,MEOBRXHHWb9a:DWc3F/_A@GgM.A?=
J)W]1X1A1@4QG9[D,[6?R]AFXf5?,[He/\aEXAK3?8VCf:S+Q-WDC&,&4f:Hf^K^
KE,60bb9?/.42Y>#&7Y4YCP\1J2^F7HXbTe-c5:9d4>G]W(Q\P<?g6CH.::5H,(a
@)O_X+ef<Y>\aH@RH5O^.Q,&1MWX+88NW]9SLK5a/IaN6Tb&/JbE39_c[Uf,;XGc
]0[4Y<7EATd0;DC3Y:J\K41DFNL:7/cH.GK:8;0gXdaDa<ARP+Y7:O7^_KEB5RW,
6gJ/,#BeBe9;U#gT8_\N7XA,Zfe\V8L(f,.:6C@Z#_QdXF^?ZQ)J-2bIG3P=9)db
:O<;GVeGa/37;XBfOSb\YCUZ\QY\1F.WH9f4]^YOOKE</K,)5\J4U0R&5/PCF7<R
MY\9B&3=_FU)M=ZT2H[^^_\V+e?+L(&_2KU(80J2H:MJ._H+8:/R:G:,;(c9YCY?
(L-B@G\fI6I8_Ae023e-H)_V&X0UMU.#1Xe,Q,dOJIB(@BB0O8,=^(3=2]R6G+FM
C@H/I?ST]3&[U4,K[MRfO46be;6?=5RM].(-YU1Tdc7_+f)Q\VQ]F<>9.aQ8Z[.R
^PE=5VSB:gZ.;48dEa>=3QB.+cOWaCNGKaeSQQ07C6Y4XHZ4;6f]e@+7>2EfUYR^
Q&\G=e19,8DK?Fd04;QHZ#T[_CVZ(?)GeBe/W)X[T3eBL,D?-2KS3dgSfW[9MPEH
af/PTX,C=TgfbP.eDCVBCY0E^TBPTeE=_TPA_?:.5SOd7#F?RN>R47fG49NVXaab
3;>O2.@+,]gEF[TU+b[>ZU#,M//RLFW4(0&&CC+O/)5=^7We@+DS8Y[c?_4VB<bS
6;9YQ9GS@9D-gN@e+7B20GAGOZ_N4)&GSUQ712H(+RJ><UNe+ORMKW4.#ZHM>SPH
/D9;R#fEMA0a#5/P&/(BV:S33ZY4Bg6V9UY+0F0Q4^KSL+eb\9,1J;[A7YY]fe/_
cFAF61QYF=+\:W6,\KG4Mg:U3O@0V=f,=/&ddW\d/+OT#WB>PZ_^=,XYf77;YVUg
^8)-50B(\3DTCEbOdGQ@:?.P=\Of5dR?d3;,7OH83K=RI_4Nc&P<#LJbI;Q1BXF^
E]U.e^3B/<1;#OAPI1-BPJTgAHC[BIRMf0QI81f&eI]E60[#/TLJS&TW-bCS>8J3
@>&TZ@6b=PD[+R5V-KTFF3NGTBQ2VVBK0@gIFPBD7&1NL#APOZKaJJaS/2C:#U3Q
.D&F#e6[W+L(Kae<IDRgML:#7f.[Q?VHC\CF>]YWaMO]/>0_FCHg]5MX)Z90@NN9
?#3;&8BOUg+U&-f[A?7@PF[59)YZV>L;;^?68^(M,)<2Y8^T/PN&f+0)e(X-Z0JL
SPOY-H;3fa0;Q1\G6ORX@[_RF-M0P#:D9bNaOVTDd<e)=5I(CN&.BE2+LeL#JO^R
;S2E^=USX\1g[BbR,=NMB,R.PVHNFA0.gfXJO@1B6@T,T[W\VUL]UH4<#TOAcK\M
W6-7CI3]IVXJ?;F[#UFZ-ZHFba<WQP(fF-R86G&Zg9R(&#S;3=M>A3Rcgc]b-PdD
g&[R:FBGPa<abg/(gHIM/K;^]#Ued\V,J585/YV:dB(.RGNFcS_<L64QVDRS4Fg=
JU2:D73dd/5aG#aT7e],F^b6W(C,RAFc5;MNFRF([;#NGdV8#g]A(]#87T.c=#(E
\R[_fEX8-I>b=5CCIgB?I=BB,/O]?aEQD(f)6FCWO8\;DeR4^C?c8F9=2_@W-1PG
QJG18YCRJ14d#gROTO0)/]XOU6XP,(FQ9dV>?G2)W53)XQ+eGaWW4eWQQD#>(#SY
a80D1<cDKM#TIA0<fC6_EJ^e;9+45N-K)dH4:[;WdYK9#/WFU21eG?[EY5V10QL>
_QRHdEBO9+eBafa,U:QH?;C[#IWX;]Y1Z;YFD\#YZXg0Vd)3TM\RcW),f;J=;S(+
H\)4JW^Rb6J2d1[[OT8:YJ>JVS<Q1b+Y9=Z;Lg=dZ]fdMK7dcc.FBbCK28\IHMS2
VS@HA&;I,TE.G]6,bD6@M;NW(4+IFA3Ya_TIf=O.@^IULX42LWe,1g2(B-(4YS<W
M]<?gEa,C<_\54@.18R)Fd80Z68Z>ZCX6PQQH0134((;HHUP950#-FTH-+DYDC4B
@L&gGHD26OZ:4U=5FUAD>[C5TQM]PBHMVCCSR>]LM/5:AE/[-GATHa715;BD&e^,
fPM&g+I<7DZ/3^a#@8&Oe_DbH3c?T2++0dY,YL8^b9APNF2]FZV5EIH@cEP&.SF.
aO<<UV@=4PS(XJD#,\23]H)U-C#>D]PPZcE5[cR#A=].OD:9QJ)?3>]fD)4Yf@#V
(9DR/F##^f+A.BAJ#S#b@3S::#8e+,;<d6U<EZCD8;5R_/]?2N#V_EPd/8b<WW3a
8Q@72TVF42&?V)c6McV5,[(a?TQD^B^CSC;/W)MeHQ@7\R3/OcA7b/.])+gCBe,e
cVR?UZF,1a+W5/gdWIAL5HN20&O0R9).RZ28dVUQgIT8]3Y=bWRV16F9L@6d75//
8BBVO44/_.9c<KC_<67ZD4)3MEVGaYd=Q<81H]cRcTaD^H=D;J,H;K##<T2/9_JK
KgRUK)?@gGZV[cbJJ30T:.TQ(c6:7b;8,O3\^a2aYNB(OR2;:8\(B0b3PF09N^Ge
&T^AI6RZ8#;<.[-SM&>fKc;P)^e7SF.TN92-I==O;N33ARaZUZD4Ad2Hd&9V#X:#
K4dcb6b#^28ZBH.NPC^X;6Oc4?--E]c9LB)LTfFLM6:[(5^LE(34CffbYLC[a7+.
C5\gdB<)6O&OJ([P15gQ]5SHC.L&W^ENdHg8Z;8&ZR5\d/X<9IfbRF0DPCbB\:T\
O_d;aPVeHbMD-&IUE+X>].;#0b8;aWK_^f+^@MFZ/[K_f7(d^L(Rg_V<G(Yf/?PU
aS&IMB6ZT>4S6dM9:<@_.aAVL4\N.::\]D^IeaTeCQ(W1+deBOX?W4B(E@+E^cd(
3ca5;d=#LCW5\DTRK<J;:?3YKd&c4&F7Lf^JIf&4#->LXaD)M)7SaeK8KZPYbS7G
?0=GH55_MA16O?gY=0T_SBNN><]c?.T-MGWLTJSe(3XM3>\K(#@-9;6([SLVRYg?
HH5,+9c9Lgd^&0TB<;P[Z0^DSSWT==3?:_AeIDJ^7</g\[aPgb7P6@J+L9<LP;DA
OZ?UW]d94\G+SHXR]]_U##[=c;H(@88(:Ncg=@?&-6=Od(S>-7T[?6,[&f?^61N3
(,)9D+K<7RQ:_84GEG[I6_9FS106O8-V<1+1J\@XKW/K8#WP5A#JZ-/2P0.P2AGR
C5,@@Kc>fU\R_9=;[dPY/aJK7CDJQGVe@5IWSEWJdOG\K[[Bb^O\cK(daG/2(V7]
eF+Lb.RB<B@5UJ3=B?>1<?C+0M41;WYHV-_8OU9#d7>H<=13@Y2^.V-0d##&RL5g
[Q-DC/[SD(7V<d>;42H9Ua#g4;W?P6Sfe3W#OB<9MTgL&X^.>(+BJ&PBe:?BGe<e
[ERA.D8)GMXLI[BUCU)4;9EJ>3QKUc?]V2f]AXf_GebIg?MD;IKUL39GUDW#LbUX
V29aP]^BNd+ST/P\MQYYG\MBY=S4.6@0AYN6[X\VO[^(6+CbM@a?)MJ]YJU+#?3U
9X<FBB(DC8=N3)@@O\CEBP^4c6QK=SOU/W(9[^Qf31V1S1VRJX)S.bb]]b1]HLZ8
(bN:;S&]=5T1L;)>7ea;a6]/c0E?ZEXPP&<^_<^6,^)06.DT4O#9D6#,TT?5G6OF
V+=gDRN9:)K?+Q]QX:]/47FY9UKTOQ,-4^<:M04UHe?0[67@,Q9<:&KaU6c63GQ#
U]IZ.<O/S5_gWGEZF_+R+5GA(K^L?I;f-2GQUI7]PLRUPSR4HRf)Y9,7MD#>[9C1
B0;:-DQ@ZI+BHTBRDe+>7g@(@aXRM53N2J7/96IeJT=3>H]]P5]cSL/0W)1WR&++
WdD\K1.^F5GgGLX3E_F/?LT<I#4M/Cd&bTHD?RTKaEHg5YGcS?D(??c+f[d5<?/_
N(JbA&,3A0Q<_RHD3T+&GKICc]BHD/AS]+^].)0YMc<R-=Fg@F62(U+_>@:e<:9?
:d;c(6cY84_(d1@WX&Pa,aD/Sf?O#+<.N)D2^K;&JO-cgNX2_1JV(_FJ6ScKU6Z,
[LaX<[]EdMI.g=Df8c/JS\b3;XU_GL&NIf.f\KZ7X7W=g2938<gRE;D+d\O&cG(\
/b0S_c6(L<CMKRBDR]8FO#/JDOF[P(5F:1_F&M_58]Z7aCFW8L)G7&.dB9X2R,>3
B>CK/.WJ?)f>5?>Z[OAPL8DY9EM/fF+_bO4,YLJ<DDIYQI8&-85S^;Q0.&,<Ge(L
eb83XR.fTKCJ4DaU3a=,R[3J4@YIHM:OcFC(bXV82G3X(L8I8>AH/]I//[FeJWY?
K@DgNdB9DG])Y8;e]N_AFJ7gbUH+bR+=XMRd&0GT@)3Y@Gf\5ADO&G:N/R6=8#K-
WH<9MM(6/[]Y]_@7@B+VHZgb\-Jc[NX;24N0(Vb1g,@D6a5e\a&.@HBc23--#dO;
-aK6S].f;84PcGSG[&=K>T^OdHNS[I53+SZ@dQ.8Pg2M#T0C#UGTWLP8_WLE85&,
fIB#NU;-bL@U>R3PINO1-5S#.bO4c8dH5^>>)]=_e#W]FL_/L6,0cU=1RS]?d_DG
ZE&LM&-CWdAH,4VFM_dUHOHI[XE=UG;IJ-d^;7^S0-?BY#6@+WNgb(fQ^F.B14RJ
dD<XH;6+6LK;WJdSS9M&)_gL95\XWf./ZW9fCUdYbK.2PK<_)H7\>CDI1DMF;GDU
.(aKB>G5f:5c8Q7O?<T-cUW;LQ2DEbgX3K1e]R+HJ<=G^d<@Q\e,FHK\aL_>PZ6.
#f[FD+B4FG#)02,-=/HNLFZOD904:?WS=YV9Zf3?b0026L]I_3LHCd.40a_=UDT+
571VdJZ@M>MUa0Ra;@9JE^b7e33.D1CPJ1^Q,\X^K?FW9C2+HYNESU,0gGSNNeFW
8KcAV]C1<MG8(:335>5(^7g7B.Q?+5ZG2fCTQd_,D7,LD].-J8A^OZWFX(GR+;c?
_ZPV,F7GMN_3W+_:NF46I>Z,O&,JM8g?ZCQXAP<0/&1[5.NL9bW<M+M6I..G_F4&
g.?25E#.CH?8B[-/P9JG.)//F9?KAJSFR.W<e<(]ETL^[S32Ac46OIF^(>I&eePW
P5cVW<WABQM4MfLIeR8B4YK25.WV@T6@1/-#EP<a([&LA9+TKY,3P9-XR1fPV:N]
P=J.4UM.,9<Z<11[-/A>7,OKUGQNG\^\>=D0&GJEXYT8=EA#SN4cgQ5V9QED+dMa
0QCHQ2,@(VfFc35:=/&W7>VK:V\YH&c+-I2NX]c89^b7-^ad>^&e)]JM3TBN^MN-
5,S9?()dTLF37R/UOb)/f/_IJ6G?CH,)Jd4>.#HP2PI0J?89=5B>NF/,HPKG#P42
X>YLUeJ,E4M->]]9/9N,3-AG8d7QB.QZ<,L4USB]HbLcTGG]#LJ^F6/Y@5N/?#:B
>&8R-B)3D9]H5L+IA0ERcOO)W7D<L]FgU/Je<PU)SA[g^6Q[<+g0FP+d&:&YT2RQ
W#9\\,3_WD@#@4UeCURKK9aQ>)Pf5FFKf4K&MV8HS/AaJ]N/0P--T7I2CQ=c-gV+
(fS,NTU]#\NA:ZTB[BEU+KP@QQO-J?&,5fdeeE]P25@EXB?2NX@=S/412L1gUYL2
=A80-G^[c&K/_L:e5@3e@HPS:.^65d9>cFP(,L#,S5e2+BS.0NJcT1:F#IAK<=K-
)5(K_K+V8<g2IC;bQ@T7[//NdSV<ANU-[6F[Z966W_3J<YH60V&;G]bRXG^&JF/9
8J9B0_aJL5TG5@-c=<>DR4-,PgM)/RW7S/T595=ZP:_>1HAb?UWT3?[_CDZ2dOV@
0\<TX=R2fWA28_&70e&?+N4G[A[:99bHLI<C@[.EbEJfLMcPFBDNEE\IS055D>\c
]](6?NCR+NU##e<1_a/TW@aOP1N+=0J>86IH-#1.aL&g?c4R5Y76A/6@1<S54;/3
,JM5.6]&I(1SX3bQ;MY7G:HN&NLWC,?A[#_FNPa_^Hc/(E#.I#ONO1ICHfQVG+<Q
O#=;A-(ZY<IA;,O/\9#6_42:7LReMY@F91R7/?dfU<CV7#JRa@QQ58eN?W(\/1(0
UTPbI>QRKHR7[+>16?4:>0>SBgE@FGQ.5BY3UCYX=a=NTgXA6VD9FM1eB<5<765d
dFL0B]cDLF#eZAMfS.@_:T=Kb<>?J)ZXZJ6-=L0aOEXdbH,dHI6/<L-TF33:XBZ;
adG@KZM^YWCXF;L=@B?<]C4,.dT,.I)<+^9g;EX3gIc=J?BP3@IXY7\-6&6(>6;b
R[3ca=>eDc<DbCSZ/YbbU)L7#CY#)UaM@XQ:4TN.BU:K;EJP7X(e6Y9_:]CZ>56G
_)e^,X1I+bO^a]@XD9Qc5ZP34J:F;_+T/1C4@Q\e4B:@<Y](\>8BDN6Regc)V3&N
[-4Ac_?e7&O@5JU<BRHU?Z1O+aA^U>FA#ASK\[CR7Z-Z.7>/UAGC4OdI8bf2FJdC
>E]X95b9c?=N9(W)LC-18@\V>>6g[T?-,=eQ39^4?#a65#RVM],B[59]HQ>9dJ#^
+Fg\Dg-,c]BG[A(R3<SB.23@C?c+T9YT5.Of&XYH#C;C8,ONO[P)OF,Cb##P2K2f
,E+)5W7\QPTaJI,+N_5HS&g(]f9K3E_Td?6?35#?G-B8_A:9^_QC6-@Z8L4-A0&b
3)JTP4H#I5(7/DS=4bXQTB=@=QO1D<+@^(,a&YKdN/L=+bPVPR[G+aB-E4F1&L1J
&eM:#cRP(G^.:^bR<e/19:51C_@W8G+CeS_N\aDHN:F6L9-ONMR4#8)+O6f&+D;/
Ya\K)HW:/C\U:YaX(Z[&JVG(PAg#gE55.IGOJA,=T83\E0MJP(0=TZ.@;.=_1aI?
@dD3,OJX86BPKJH=GX5.F3_KdWZGgdLG3Z11:&0B^J#]RSC.B23JUC4O1bDYc?42
)(\^8H84SG_<?GT#\S^(R64A0RM+EAVM?ON0H117]f)X.H&BB^^.dSW#P3=7W^<P
\^VZM[SB+KRXEG=.7J&:)SC:DPZN>4I??=S1ME5G,6f3>KF2692A^c:W)YVXac#J
C3#-fQC\DUJ/]?7,\_;MO_Sb]7J;=QfM#3EScU(?@,/<L<=ZVV1=K)(?TgK[29(]
L+a^CS<;-9P[.T=VNH)cMM&f>EI&7),f.ZO;9OZPYg(BD8>4NDVN\D_68L78JAZ=
:#1.ZIadZXKW4d&=9a@S?=]8@&0,7Y+U,?FcN4<B1;X<9YEZ^;_1QOQQK)/cPYR[
-U8O=.+\V(PP?BEII9NH</JfdgaZ+bM9X4<A,@<f=6=X81dI\,VS^QCF1>,#1--C
G[GCf0[@CS/)Le>E#_TbSNf?,cD/Of@X=0[^\A^?;T>ae4\2051O=DF6##VX=Z,a
><,N=G=(cb/6^A1c.YRQW]46E+YQK28SQH9H23e0#LMM9=HV#BG@240bI\KFJA_a
M3=AO--6<C2:?Z\5e?/,]ZXUc+OPT:-X]VRe:H&)>8ZV-0COD.<b&ZCKQR\I90D)
-bcX^.(<O-e#[B5B0X\68;4AO3cA],Y)JGC4d7&<,@9X6C]K:8++LE67DIX/]RAg
HI,PgAH,JUV\38IVA[cX74VR5>KQ[J8#@GJX.NbSeK>eBXBY,4&<(82>7G(CYdKJ
UeR_Le;IKV#(AQRdfeK2^c6dD88-5:IcIY@c:,@ac/;P_0=9Y)RV;B()\d?L(E6I
DI:IZdPLe__U][XA&BZ2/9L(f5GBSLV@\;FQ:Ba0f(S?HM]cIE9E0M(I:YS#/bfB
5?fF7N](1^FV0QT4NIXYAbGHfD,2bVaFC57Q-?I+K8gHZ-.V_PHEKC2P.-YeS-,&
59O4R0)V5Sc36bI4;9-P8Q>8Pc9HT,V[\JZ]a_g_?&T.K5_14L4AUIcb^YXO\\+,
8b^MZ(,XWdcG-5KOQ=-],b#>/c-2e.QH-:X]>CL;KR)+1\U41C;NH_S);#2c?.^N
EZG;L0L:fJ,7GXg7.7G#3RMF;D[ZS]5A+/[T8e7&UVHa5-a.a+e[dcd>Jg6ZH,9X
6PG9#4.)>KGGO0EDQd\ee_I#5GgbO6N&I4^)g2R,LO^MPEC>_/T#PJBcD;&@O-@A
ZJ5(M\=O\(ZSL_^9?=L_YR>P?BUF^:eSG6J#T7dK4JZFBA<I^J/@V,MC6R;\FW;)
AJ>3a8G0N1,:.gSM.GgGbQT/:eC]=Y<>M8R)U2<\\.MJAO3G)ZMLbSP>fPNK<>8/
M;F4fEL[DgQG]P\V?BgZM-79]@JQP<aULEM2,I4KZ<@XcQFPDR6;>IU)VVMd]5a,
JTHbMF&8DH482UAK_0@DbI8^0W=9._U52K-e5Y.)Q6PK9O6/FVa;,K\M9ZT]M+0\
Q3>5V-/Y&S9(9R;0/eD3De\ZG#>CQBYZX@>6&L=EC>975@[CS;2N]V#cg68?#+[M
W]4KA=F=aBB&]#7#P(CBYX5G)Y,^C+<^8>fC8/f9dSgK2e=>CC1=Y0g\EWTA6XP)
@gABW&)1=(P4&\IY\#,A/5f<.:SfVOR76Jc_=?U>d]KMC7GO1:HC2<B@&>7Q<UVN
HOK7-6M^<889C\Q^9cF^C:O7dTe_--R]X0g4H-M#J7;eO;D1NA)&fR3;JKFD4UQK
GRg>eC^B3Aa8@JLB&#\2&eO8G+dNJ.AMX>cNHX2L]\eB5ec;Wf[>-3<]&I).,8Na
:RW0f]cfQa.?2H2Q=)(F5Z_P3Q,8)QP7<>4,_C+1cad3QU?N+LP9A_<<MFF?(DV^
)6>Y/&-5f.a]EG8>\<e78F97b&0)[/M6E>&PPe2&gAF)S)g4[;JfMJd@Z7O<0J2)
\KN7WGE(EgG9<OZ,9I]eMgTZ>O#g5:<CNXObQ_C2,>#8&^L:O0(3GQZ/1HBQKSbc
/&T3.8@PSA,L=SJ&U<[a]1Z+@=E6.Q:FTMDZZBN;R?TEPG#?g3bU?E]f:FM3:0=G
3V+K1+H[acO?T>03RANZ.1Mg]C,<I1P^N@^807][];gcST@ZN8a48?H3\1SN2K-2
0fI:+D0(#f_)@E].c0:HgMN6X^F3@3/3)UCV/:1DD2g/2a[aeJ&]_e@S/U,<8-dR
d)AWHg>[VM1g]I0/^(f2_,Y]-d(-ZM-;.EgMP[T^ffCCBXa&ED^;I1-5/_+0W\Tf
4AO49e.EFY]IaRV45CK/SC1bP1ZY.=g.ANG1UTG28cU[K8VLU8G7WeV0:6E1MKKI
+1V^6=2/ZeYfVNPTUZC>4)DJTJ#DMT-c@BA-\&O-&LW?\c>]1a,GBS_g\_V=S;(>
Y9d\+>;B-#+gg2<=>Bdd:5)cCX]T_4?1BW\LSX.SY&P:LIO]Ne_MNAB2]:^<(_67
NCP)W^I)O9>a\EMacgA(2/92671d=Lf<N5VJ]EWA+PC?Q1E5CY]GPSM-8);BJ4Z0
_g13bA22CIKX)KEJ8IFdU+16EPF_KW\.TJI8Q>2.JPBfF3#bZ?df;553\e#eAOG6
],R@T?F+#0NC-X840G=dFf<ed@Wg,A&XXcBeW.:[g6TP?K;f/^MK5-+eIFIC[Pg)
O6e;F_;WXe9[b[^d.aHc#g)DS.97SX+@a\W<?@\-S3bY:VV.0I-E9\R.I:J/J+a<
H-?AD@MMFA4+J<Q718+)=?LM=R-@TcP/e(?b;M.[S8&]+D:K>5OL?I:G/J@Y;1AB
5H;CKZ:If?@CE/HG/06cXHR)L-d#7cNW-#7R)ZgB?5ZLJL;aZ:7\1RRd9I3UDbc^
NM^TG)<A96MAb.^LN=faGK/V[G4FXR1+<RUN7+U=Wd3g1Z6?^eI9R&N&HZ35(MG\
PS&#F]BE;_KbDL0.7YeD(RZe.;?eXE+G#MU<A5g@)Vb56D2dc#J0=Z(,BQUSXe)<
B/5eE[P5@LV^SRcaO77GX-B5=LK,HgF\[g/YRSe6N+X=C5PHR6?:befFZd>LE[?F
3ddY=4+EJB00Mb:ZBW8V[#Y,\=Gd/VTM/HRD^Ke@Q\-V1AGD5YJC80a8.L[eDCB+
<3F1-\+;@\Sg9gR0Oa<Sb47F=>9J\1,#<>;gN8:Q3gV(<b(4=&/D0)_M+(K>-G-]
[bc/X-5AK,Z#9U1fX=F222_BG/0&=?<YOW_RGK2F=f]Ub[gRJPI]c0YD7TUO4DJZ
/?;\KY<SRZ=DHWSOg3IPMbW]PY/L^V;Ob8<S2_?JRK38K1>Cg(TWJ[Q5L.LfX;V^
[9e<B_N8IW\V;e(V.TD&d;L>>F>/COT3^_+dfOHC1Q?ZeY0&M5GH3B4=R)J626H-
KVA(dERE<DZV7=gMb-Y^O#A8OeLIbNBU;BK5\R&cZ1,IcRSCNSWD64WPNJN6VGJZ
0RI^F/+(OSe\f@T7+,KLE#7=,,RgR[LK]-Oae:MM1&GEaDQ.:?91,)f(<+b<^#F&
H1<R;R_3+^I\g=#MB>R]<2Q^_R#>B,,]JdR:Z1a0UFf^4ceS#S-)Z]T@D?+Z^,ag
B3E?f?CUD+^,^f@.Da1cQ1F[6DKJ6&Q&L?-=9Z3eY7TfX8U[2XM_R;R?dc@eV0cH
D&0J-#Y^8D_M5,=X4ee;RJJIH9T(35K<AXW2@Y+\F)3S-O1#H>O68SJEd.c;Z@0Y
e;YOO<V1/<e#KXNQ<1;0L@R\>PeJca;f-)<(YeXfacNRZMP+=1K.?2^<^5HG8;gH
#1>6YNKD4g6;HX;@)-?5/+O5J1d,U_5a9<-KH+N7CSBHQ5IYCBE6C1F5X?L<;]VF
<E?P-3PBZgRM7+T@/QY6#@/cC_fY40_XO?(P>K0F=U<K:3f?35/P&2>2\fM16JKe
-39.OeV^(EbY0WV[QAg,:[-JFP+;Y0VVTUQV5@2>g=Q5AM.YaaLK+:Z.XW02ZO[F
Ie]bFSE<cJ3XMY)7K]Ga?Q831(b+7B-3L).Sf4;[L?+eEb.)\XR-C1M(3=L.-\VP
JVB2[DJdDGKBcVG@3,Z9-Ue5F]]@2IZWZ)](fc]QUV,f<1X+a?AHI]YA?@];e\;1
4geXPY/ZV+OTF:L)@CP?&,>?^HLG52VACUR_=a#)F21[[agO.F9gNDELKc]QJ@aY
@GZbf)?N.M_g9K,3G(,G]C]9;5KB4J0=I5/)A?J;]C^g)^9+?O>R69KPFGR1>AFO
CY>\/gd)HQ?=RZ=J,>d.4KR\0C_FF1FS2K?(KV,-#C&PE]V_M]HML4Q3BJGFES=>
X1I,34@#U&?U1]7T1K>9+P#9-.Of@T.+6\-:fJZ6MB)(1NP0MKa@?;2WN0ZdWJHR
\[)/0^aV\PId:9WXe=K89TF3(+dA]IDG[WC+Y>6L&bVEW8,JXVb(8(BC0OfK(K);
PB8TLP9N&aW\8?bDF@S]2\WFdQ&TU)4Vd-\+6&Xg#,0eg+H?T2B.NU68&:S-^4LQ
a1[YW636<HK99@QKM:54@f\\E>C59/L,0eMcY\A]K8)[XEY8F]^KeLaT98+>=5a/
+Y(V9SZYRdCICM5J(L[:5e@,;HNXT#8_1U63^.1DKW]5cQKd.Q=TJ<OYS]&^?#5I
3<JXQGXNF:O[8f&9d(e;8e>H<5]<A4QE(2S2N_&/AHW]ecLaF/NG:c=NL);?]LJ,
N4Xd@L#HV&05]ODKB+3AJ(EH(>Q=,S?fA^,0F2a.N;QE/&.fIG)^>C_2,WX;TPd^
DIJ72#R3bCJAdc2?cSag5])TQ&&Zd=<g2N_^&RZK>13Z+fS/[c#UZLeVG;7DATZ[
\dZ-N]T\QdB\E2&\V(U5KL=LOMV4^(@RgBD</aKT7@=Rb6MUB:&RM]]+d.>Cae?T
^PHU))&FXdCKP),]:?)2Y89Y#9[^OW0VgMGHdL_c5<a1=8+OMPH8a2Q8Q)BIZ,8#
\]<\db3M>;HRX.H1/(Xg8E)eY#F\H6U;^Y>3BVWE-10fVN4Z5-WYBF;1\=:DJdM<
c[KK#&Nb3eY+8HbPT24/7PQJ2?)48]6UNVgbN]6c1HQG/LW^a>R-LNTeSNHdfPPg
ZQ.>(]LHe#JV16>_J+cQP:(C2RS4AK+B5dY^?fL9/&9<9GJg\^1I#^((3g8Nf>K3
0.<IF&b^S&C+3JA,(Z##?=8AJ.+AXEB@]WOL/295+WS(ZMZ\d],/E,OXb5PI]Q1L
IWZ5OL?P0H0>I97OH,aL.OIJP#df03]UUI1N;<de_;.CVW)6?f.4FT02UES,0Rc8
H2]#^I8R3ZVPXb/S7C35ALF3L0LQ2DZP?.g\(eYJ>4VaNY[:P8S>4W^9fBHM50YH
GTP0M7fM<J1TAYJ@7BY+B>5A?Mfb0A)ZXaAQMfR,Z/9M9:QC&#f,ZQ6M&Y:[9<ZS
??5=5UMTNQ6CW0RF0PF>?VaNJA>gU<ZFbafBJO=aBP_]JX76#-@[)?5-B.>V_<#D
B1UBQ3b#F)G(#P;g&ZVDGA27]ANc6[Z?7V\94#2AFVGD0DC@QgS,^)=<,ZZJ[Qb+
Yf(]IeH=7<2+@e/FNKA\KU_gC]E:WdYFW-6L@dQA=9cbCAT^21B&M3.?\Fc=1B2b
TK8#A,UP)(7=V0bWYCPf@-3+&.e3A^ZREd;5Q[X9fgde?STSQ]#KWPBG@G<IX.(/
M+O\(]aQNK3[E(1eT@;-Pa=,EM,+AJ>?-PG/PTIA(9<WO8O)XMd]dcAf6?P/;TR:
B</5cMUg)PXRM:H.(J/fNQ;f0/ZVBJF8U/gEWgZM&X,f&7a2WUaZ8T[ZL@5?Y=d:
7M?TMX-D[#4bbQcHa-M)+0-5-#:UB7MEE9@N>[0N>A)A:74Rc__LA?#0+,56IRZD
3<JI8Z95Q<Nd<F9315I21OgVVDBM(+KO^+;;?WFABYJ-NKI=WKP&G[HJ/YI(<@e]
K(^1#C8E)b>ZC0IEAYB-W;X,RT3+&-\ORe533FXNI^H8R.NP.WeL3d&LXQgGOXD_
;3A2>EJaKT4U#:YIA8#F@V)5R:Z+bb?S6bQ1:WF]GQA7;;aD<.-EB:..5LLbCMbW
@(.SXWT<2aL^P?_&_YS&/QNCZ>KII>H7b2[D65<ffH_PaK&I:/3.9gMG&fL[J#X8
=/E;HJbEB<T^AV=&F0GD,K?.P&PHU;KH#R/(3,M072;8ZM2)2D>2eO;5]aREJ0[A
>[F+FG2Q3Lc:3d>:HM?d[=.JW6/FN9]SISH3T63D#=5_NDKX=Z;D?U:-cK_+9MF+
V2+,7b87\.C=/c-2?EWVCW1=:#-bG4Z7EFHF0SZ.,BHN/c;&)7N4IEU)7K,bHQ\Y
A-RR,\PLBZbN7>/HaE2c@/_+&T7(NU_:[XF[680_@,e^#TT:Q-JGM^3(T0-2QFN4
(0A?BW\M_c>R4H0_b?U.N(6@\SLSU.,+62FNgc[b2/ML[AI\Q>W34HA,D.#ZO4J,
R9cCLJXN.G3a=-:b4VaR?Pag4X2RS(551Z^Y4gP2S;KHGSFL6./(D^8ZY:U37\,;
6e.Pc^d5F/;.:.^SMbAIE8X5+KJ&a[]E:X[V9<=f>AWGD<R3[U@E=8e2bcEcUFM6
=C]8KU64&RO,30R:4LRR9K;;a#RY:ZEYZag7^Q,XOd)LE)1OLYV#1HZ-R4]DT,QI
^Ee^VAV7Y3@XMRJ&3RO(LNKW7/NZJQY.CI<AG3REgPZ1IMfJ#Pb]ZG8N/]^3Mc2E
I,&9d=TW@e-=QL[+Y^)C@D(A)[K8@6:^Da2A/]G98U[LH##/aeMNE;9@[f?4V2&;
B^C>2#,a9YEf?E.6g^F9/Z#[Le&I=>Kb/_IH23J#_.C8D96Re&A>?#MW+7V4B<PU
2JBGc)[d9DdT,.VIM0EWO.c9,K;CLW2=2GeR(1J&K;QEDf&FR841L>8?KaN.IGWS
P_W0BZ40#)NWH/aLAH\,=X^4^EPL2.):M2P9a+WgH3\+6Wb#:?4E_=DgAB>QK\BL
26\<)E@8+4=gf>FEcN&J2[Pe1-8c_]B)BaE0G/g7bQcK:ZFI4MWC>RQ,R2C[U\B4
GHWV#UH5[cUYAHY\:=]cNB(2K?4DU-]Pae^A/,cOX^:H1I+(AKLBGga0YPb3fIVg
:.0>\@MV6U]G+C70Z1KMaB5Q(WeQ0E@=0CgGF.I^XSR0OK;fEHaY<^GC&6ZF[7LS
?eVFff9UVT9gXdF<+N4c8LIKH3N#JX[6bSMTLWc4QA^E/4e/R]?1/Eaa&bC<Y8S2
,7A[g3IBgb^S+UEKBCa:Jf]<6b/RPE3f<E+E8A-f0RXGD&,@Zb-^6<QHQ/7\FL65
.;@48Z5@#bHV+b66+PG-:>W\=5d;T&]SNAdY#(OK>^ce9,&SXEAWMX5[b#U<@/V_
],>G;@/V@479B;?(g+HIW8D9UMK;dMS09L7CN]RcGcc,V6FFB656052RW)Z(U1?O
1F.?c(<RKW=/2_7/7C.<T[?U<LVKB)(=,<H^1=]UZ41KB,OT0._9<OZHE(R4CDGV
D+8+O+W_)gON&;gXJ<V8\ZS3(2G)4J7;&IB#6/D2@X,e&GFH63Y2=R#PBEK]</3A
O1UaUR3<gL\d@W;LGe@QMH_.&D#LYN=T0Aa5MXAFGDb\Y/U9/Lb/1,01:dc,aI>D
F6UAJ+NOA8fO5:+?4N9N<IUHNE@e\=4DHOU,B#?YSRA[SBa_W8?64+bd+QVNP,6X
<]+>>ZF&N7d0WC,T6B7E>J?9++[gD,<>3/LKaQGY=Fg-Wf#CBA?AgA7b=,(F58VT
0;e?beYPPR52KT+5:3S]7Q,->>ACB?[f.L6S.7Z]FTg2+SNABDIE(DRRe10I7aU+
#Zb&(PI5:GX<D5^6a:V8_,WW?KA<3SP]0.aVE#dc,bO-3PE1]b17R<(\BaAHQd/4
d\,_;RHeW5S06(d^YK1Q&)YEE6Zg(#(/7J^DDeP@H1&fL1,cR]ScC34Jc1=K6KS(
?WN8g^bQ#]-d(d-c=Q9M&aeOR=PK[F80+?]Y;(9@;6E[_;\82Qe5_+1FQ3_C\2S:
Nc(@TebE_1CeYWDgF(eLaOf41,ZQgBV;d@bGH=W[4B#L]NJ@N85KS2@\R92FF2=V
5LDIME,BLL5IN9YC)_B8CA<1g0?8gbM(_H/aF(XEMABNI8^O[P>TNO#aQ6ILO\0J
8d+/f6?TO/-(^/#NE^TAa443aaNPfa^DA(B<Y-,8#T)H7W?g@_C&\LS=UFCZe9X@
MA<;&;2>Md8MEQH=GJ[=cf3(24E92(.HYTIKcF6(RHR[6\,^B02HGg6:D_)db(9;
XFZQ>RF7ZD:0:JTUO/N\_+]]1b)-H?+<e)O.5KZCZ?d0BVH:0&c<P,=+V/1D^?/0
/CZPeb96e3#[01CB,8_0\3B)69#/c>YKNWPOM1]Gdb)WJ)C6EZ;YT,>g88T7Z4+@
4H>dL4R-.4YW[O9<-f^?RQ8gDP8T.:O)8E_eJ;U8ZHN5=0:77bY.gI8V0XC65U2M
M#(@1fe7R4M<LF=]1(dX<Qg&aUSWb0EW\B0WO<IT:U=[AT:a^1-N>_M)GaH=bf.3
Ea6&]fUX^/;G&E]9-GL_+[\+XR=YY<S&H5<IbUHB_9E,0d,BAXMCJ/HAXNUE&cF(
3X^KH@-X3L6e,6DA4AG+H:6&[(C#P.dT4(R1>Qg[+K/ZGaT&)W(,=?8Xb#6[/T/:
cN&5VaU[]O(5;761;Pb?O[e\FZ8U?-8>J&(c;7O6EU;5.;12cSJ#99K1@c3RGL_#
W^7(dF^U:.SeXRNOLC0[2[1_Q@UI/9^D33PdFb&&d0(-D8-K#A#-/4NX?]7U:8SD
:<FL3&?.H1K6-2F,b69RNc=KE.#:PS<L=NeF[1,3O5DE6[[D^U6VXVeB:RSBR-?3
+.M)b8-gBEe/3XF2YD8W;d4?/Kf1(U)#;W5X)Pd29MB-A^0(,#K@Ie]H<R=?KSA2
,=;RDPge>3SG^1:bOfTaXE=XY9\5GJ,WA1@YfM5GV=+^#?<9^ZE-<YXDWWfD:L93
3.D;<QRG.RZ>5c]NW9P5&,[Gc:[@>8&4Z.VSdE8/\6J&/I1F2SRCZT0=UdOQ#5V2
ge6/SH9cD]D+dM4<Q4&AdK9)1UOOg&)cHHW6+4J2K-J@OL:OQR82A+>A84BTFAHU
@>TX=O0S\Z.>#Y]6H3K;&)7CfDfSSMAUZadW8QM;EaKGMDe;>@;9[4P?ceJ,cSKJ
>HX4:e=@^7Kc1Q@=03+e/WGc#89HG_)e8_G>V#ZgRf_^8N@_NP1Qa)3H[=4EA?d]
T>0TNZ\B;F(e#/gS@&E#W.R@).76N@Hc.ccF(Z^b,0.QDQJZgXSPdBIC66MX@ZH2
#\\#=BB^L_OKIPeU4ZD.R7OD0IEG?QXM24c&UI=_XI0NeP24EQbK2>87<PHRSNV)
DQC].,7;<)LaWeKW6Gdb@R4=8>1Na70<,5XPZD-M5M6I)26)f;HFA\RS(GM5P/TM
4;EU_^D,,B9UDT&\MNY<?D[UBF;:?Z8:-RLJ;\/C-d8UUB33G>2R+9\@5Q^e;&Sd
S;1(U)3#/M4>(9JY(aX,@N@G=8C]<V/?;S,UD>Ne7Q^M9;V;7#7;(bKN1J7TT?N,
21B?^.5/J;YQCXXY1#;0K1ZH).b0RYTVfW\;)BaR8Q9QY=#3:FA9;a32U\7J];7<
3NT3W<X?b5C6=aFg#RW-&\/DQTBSWY+NESWAF(IOTXC57QV(BQC[aOJ7-VTA#3#2
7(BR8dVcSTJW2b/BTN):#.\H?A64BSO.@UL17][A.MWZ\a=Y/QT=:I6_LZVb>O9N
Yg?1U+V>_5?X)B0B&/c,UfFH6SYCZN24YW^#E/baR&(8Q#8ZbR_Z-<)@b+3ME<Sa
N);>)6-EST3O.F2))P#20]XVRcgTR5J\<F?&<,HZ1KcXEB[_O<g\+bC-Mf@65+LR
#6fM&GXG&UXYFHfbdK5>fS346a5CS?#STYIO^6C]O<KK(>5>Q@9a4;Uce0R=E_N1
&NC[0#f9N,PJ\5aGI)-F94\-3G&L]B_J_7Pb-M=;J0;VFQ[-(b91JKXT(NPY]6H6
Lc)MX]T.[15Y_S.HJ@KTLa4Cf9d=FQS^Z6d4)Wg,J5R5g9:RKLITGP<cR_)@BN2#
Q^5gcdF._K32>Va0X1ODDS8#M]\&PNE5KZ\>A#?CT1E#J#?G+8+VR3TLX]2G7]&H
cY63TgO,T>;65-;&?Q+>dA8IR:2AD>I#D1K6(<La>>P;]eb_L:CccLEA&O:b;H/F
I.TSM)Bf7aJbKC\:D.66K.)dJKU?F0I2KDN>3SLL?3NHV=GE>KC]JE+62O],-#AM
E9EaE4a;aW1):G7Sf?DffMTO->WG.f]JCY5D^Q+)6GAE7@NHM&C=+0<d#877H=>T
8]HM(XSFGJW1HGGT<W/5@3U9b@8BCUASNHg@_NZf6O..Y6:X&7-@80<:P=-DR\<>
@,MO\QZG@<WOJV1./K9,#7(B>NH-(QCcdG=X#/H8@8G+).Je>aCP/T4&:K-Q+6/@
4KSF9>G++JQMM?c0;K[fQL:8eY9dd]T/XK^2SaHG7K&U[FI\a783P(AegTG.16&a
\BY3WE-5?9ASSL:38W>_R].a9A-dga2-#VGW2TE)4(cX39ON_(+4X\T7AB41B=XX
a:#a-e-EBI_AP+_6K;Hb4MPYWOUbf:a4PJc2gW1-:DI^;[a5aQ3@P[[K7G=;ZL\N
aHIAgKWF\?]UeTVK=4<D\A/7BDee8#DJF]0V>_K;b(]W/3QNa[K-JMgYRV1;]B<6
3LgNOV>SdIN&gO2E_g#CaG0aFY+eYDJgUF;Q-C#;LCNMcLJW]=X=<RX\.W,@CF&N
;Ddb[5-\,TY2(7FO);4^]&7\#_GYBMdL791d32-Y\a>@WVdBH=&RGJ-YEO.eI6,a
1I[]EY3SAQTP^C=A;U;9;H@[ba/;FG7c?V5)\X@f0d@?RNMNRJ7g1[F6]?ORPdC=
6PQKTZ;#6Y>(#\bNGf[9-P[]Q_X,X45^KK&3Z5b@UcND?IX<.Eg<PAaDcW)VJ\]X
;f-CRO5E^/Ya48e,>e#(9cJ1#;K;9Y]b9F5OR)8gd9/NWOZU5UOd2IEBe52H+B-U
QD_^0e;@cWDBe<L[>Rb)/-4Z89@BXD1,;=X@+O/a?AK67ND=REUPHULc\N>B3c>E
#B:FO6C.3,fL,PU4>1THF3HEL??UL_FL(Nca\L[>0QHNdECXQ/7R2/@TX+7.UGT-
KHVfA:fWbJUT@VK/Z(FMe09WX6GMW85Z^<4(/ebI[EeMM&MHK\YPNg]YCK/6HC.Q
B@X_IJ.ZKeU8@NT\#,e0_W]E8#G-)KK/e/c2&d6HX7PMfZ+23(M#JXN\KB=]=G-5
VQHd--E[=+6fAUT_BCX+)E>B]#6G4f;M]#999,7>YDbYb?WLbEE@0?RCQ[71CIaX
]@Q@F14@:#/MS11+[Kbf2FF,XD9HRQPT0?aF@>B:)]5SS),Y?JVR^G11QN?\c17a
d,LN.@+C4Sd6@f-.16,[\IG_]T[b4<IS6Y#_HN/f2A&Z&.)@bbc9_C[32Y,4G]UG
JaJgM./.IS?V:W1U)5@(.Y@eL+ZSb.E.F52F/9fN<Dg0]45((--5BdY>(2)S6DYL
3=\8<RLW64WTgQ&M6Ec(U0P6:+T-c6C<OMBGJT9^0<&ecB)8]BX],O5T9=3#=;EN
(,ESFSD;J+.?.#(&S0eRW@^7KCb=EGbV0LTNQ[QGAaKA8FNT3_/AP44H0MQHXFg:
=U\9CHJ<U<;XQK+LAT]L7;@:VSUU<bSG)FKM8GKY6D<&bOJB?XWL8_;>TP;;:C?W
^U8(#8)eK9L7T6-JcK2Gc0UFdZ?J[P72WZ1V\(L9.KJKC>&MJH:Z+MdX@;RG1&K?
6,.(=c^NYaS5FdeL]Q[@)G,+R1:33bTP-W(P4-1>g>./@\+LLJC3Q)>2:@d,DU[T
)Z/7_LEA7Wdfe3cQX:A>BX]NCD5[5V#^;Z3G+PGd)30^1#Td]?JH1He8c_EDP;2g
@=A4cb61(:LX-E70C]eA0GN[JcIc?_O]Le&O[LB@8YY1#3CTT962;+\4.P+X;#g7
@8W6gOHUBH4XBBJ-NMdMTb2X4VUN.5C>.\eZ9K,.497e2TQ[DS2gP)<[X6g4+CfP
T)Q7.A5#8L\S16[7+])Y_H7OgV.ZA8d+0J^==W9H#D,XdGLZgaD@54c(RPS8CLY\
;IZ#Y<CIc(@4VcN:D3?^C55/K,@K=HAV0I&B4_c],_\(0(BO]3V([d[c,c/G(>Q6
SZdGgE@XXYL@#S7Z@b9+eEa>S0;J)\=gZ.OX-NcHL,7/>_GFdUKLR3L0[O.ORNPC
Y=J[:TQL5480:_cM]839H^[V;B5H74TLI=f()LU3g5Qd(b]-g,Yg,Z2K3?_4KCLa
&YYd98+46_.Q]XYTX=S<ZXAMMY^^a])2)GM1RZV.W/d.B#G.JQde4@4K0f\Od1TF
;9R^Y0eQ^&,0GI-(5H,Zf&<@4U93N/1_=,WF6\#;LcO(Jf_gg.)f5SF9(-^_SN(I
dV&7BYT=)>0\7_+g511PaM24A#TR-C+&[\UB>aUf81-Uea^>IWb;K<g1Ld<EFMNP
GOc(S4fOI]aVAN3/Ye8d;8]cYYeE1]Zf]IQH1&F)a5BJ_.ZAPZ>7)JC@4LZ1/NU7
W-8X,0;VKgJL_Y:1+aZ)1<#T7&O13>QR(@=DQ03)SdBJU#aQ(W,<TB\_86X7)C@(
?fLF69B/_TXDG.#4_E7dbV>Ag2.aJXb5+W5,R0AF?#G@BDP\G?VdL(QULggX.02]
#d0#ef0Bc9M8Y:?Q4MS]8/g0T<NZcI>3bWdFUgM82VX3\RMCNUY[efI,U(S3K>>F
TV2@B8/[M(KEW41.FPL-8d=N[79b\5[V2K;70I7881BL4/9TPF#N4AW/1dR5I7-8
BPYE^JU[SCAR:b^dU]V1dA9Xd6E3AfSdd4JT/6O=,Z59fDG,\O<P/T3[;3aF(<dQ
6?O&9XPHQQ;ePMQ2H71/V.EfT5PdRFXQ-7,CCS37e>A4PM1QDVeZW6&S1L]b@P+-
-cU-/CPI[JIFL8XK;4YESY^7BAe9A4Z7J9ZNeFcS8-^N8JB1S8/S^NP7_=R^_g<X
GR(8a;d1,b)_8C9E-U[NcD<;H_5VY@U8I_Q]b=N]HD?Fg39Y2C,DKUUA+QLf+I(=
DL/GSdNaa)[LDY>.KcVQ-=J/.ER_d1gF\I7RYTK2NF8L&0fMd5I>(7DRV:6?0Q@W
61G(5a(c4W<)ecNaM2Sb?(g8-TG-/c5OOe1Gf=>9.T)0af0RY_A/aA3A##?+LLMV
6V/2>MUB.CVO^TObZPc@b/V?Y4P3@]D-M&;X.E1CW4K-a#B[[-bMK7[J])Y0X?/a
-[GQTfAf:-aZQUGc@2>-55.?IB774;EO\+EJ<6gW_SWEM-GX6>WGFCKT8KJV_)FI
#I9/DO4HK)Q96)W0-#OaF>VM@XJKX2MTe;OTT\A&JZN#7a@7MYf4VO2Z2-7N?QH6
GN)7d_P>e#(](P;(10XZZGB4e^GTJD0>c4ZF&S2W=XLLCV#UVIK#aO]1^OL&6?TT
F9-3LE1)MEIQQB3(:RCC-M8EIW4G.Q;-Zb&)3HD;+,GLT)-)W9QcW@4:aH]&S--:
MC:=HN&2S=BbLW#N=&1_HeB4M[1L@YH3_BcO8+6cZD+@8;_]GIS+S\]a)M^+P.YD
O7JggOc4KQ)-BBg:f\5[54@0e51B>:4AXU(_D:NUD9Sc7PPVT22;6cE\^C7Y^)e;
8QB.+BL\Z2EZ@F=>M]>YR6JULaU)IWfF<Q@=Rg?63M-QBEK<=QU7QQQ>O#+R(?1F
6e84(V823(J[R-EXUR0BV,5XF#S]I4RSOF\6f7FQ6I2ZE)d(>3]^-)\A@7(WE/Cf
e]3d,7&f1cP0HA;E^OVE?:Z)f)P\Fa+ZcR\74c/6X,=bO^C:(Jd^E^1a/S.3/NJT
DUWHDaf[0KP?<M2-2N)QL1-[,YZ4G^dNP4;;b)cS([WNg,#RG.UU_e=fC=[W@J[A
5\\A@>>dCaE]LJ7DdIN5e0M^V]4(:QH9F:9dA>?DA\_]?P=c8Q7G9E@+PgA:>L&#
36M:GZ)+<g#LJBb&TNL_&A<c<]VK6+T=#&FW1?Z1g7C[ABXaZQS;@a+IAWUK:S>:
1OTe-Q1aL^A@ba#9gDgd=Rc186_AUGKH4^5/V5b;f:_^]3WF=L8@E&GDCCTDEZ8<
52W9e>G(VIR):=MUMeEUZafQD1a_?6E3+YgN7N]0g&e\7Y06.K19^f+/;60,.12,
\]b4J<L<,BKD[#&>EZ::7Bg_51FIbCEXIZCZ],>Q&-K)Q7U6&DM8O]+VEO2OeX(g
Nf[5PcVO158U=PV1N2)Nf>=?J=Nc9J#B@Y4^_bWTAEJc380QR9aWeJHPVTZDEG#V
2DRS]f1W<]UU</H=J7GAX]c>_.eBTE\Z[G&d&gd[L+JW^S^eW^dJ9aaNYY#gLg&\
@I)8MC=RQ1SVH,)EQaag3=8&YOB5dM>B(_P1SbEf56DbIa55GP+]ZD(>,.&^[.CO
,#EE@a_6#B9#B559C15cP8=UHVbO\M?\T/MQKW_6<4R,:^MN2IGH=9F^c6fbI1S#
Eg6-E5^aaTg;LRS=J-Tc7J;dObE3Pcc,705ITZ@]_V94&2/GT>=N.A37+8--dB7Z
[6&RJ>CPYP1_9aL>21KI0[a:E?XJ_37^;^a)R\OJ=[#7I/&Y1S2[HUJ;9GZ7HZ.Q
KYU,\LFZSFVJ(>5>=dDGTZ7Rf5Zc0)@K2_fg/WUfgBXUaE10T=R>Zc=_E)X,A,9K
/:8&@Nb^-YV_gB_7JC3daK-A\B.A<MCOS-(BdRYe0.HBNBXTY.9#:V+^eFEC=,4?
D-(1-__f9/^@&/5K2beMQ\]A^d;(?YI?YZS>Q69U-\ZgP]2@-+AB.&,^M(PF\G?+
-dD.T[W;>BRD<JE4WF3OLH/P8a28TKJdQe#K@TCg8183-NOW630+?]1aa<Z;)K^3
S+/OgS/G>P,OT)8dF6P5=0bc+9+8EG1I-@0(=,V^?X4dET@AJg-&9b23gZ=S<F-7
MR\2\7.JFZ_7CG98;L+Q2BQ+Ha/;+D69603WA2EH_U\2(=C+9OF/A^#=E?G,S7J6
\?7:#]TIE<JPbfaCbTMJH,-d/RFaBRBS\b,\J,&YG2_9K:H@EObcKHUgEC]5+fbG
8a#gLDL+c1^+<EK\@f_5dd>62O<TSK.3XCWGCEdV[gV[C#KDXA@@T(=cMPZ;^Q8D
-5&^1_)M)-VH<QVa;6N3F?d-8(:^cegE>c>-N5A\E?9[W#:F1?ZN8>d72C_3V\]R
DVg;P@5RG4_>N57[?b(e=58@/gW[J8aVKK2+<>IgSM\>0)(;KA0Z.a/I>_K9Z2Y8
Oe^B(X/FZR.EZ->2;^Q&4/(ERHc55+4)Y#JM-_D,JOca[H7Q1O:a;5f;E/PLAAK>
_WaOb-@gb;=eLAT,=8d[QY#:UZgCEXB],QFg2&>7=,,(<Q:Z<2J>Y3:<a_>572/H
9K(_fcD\;_9D5@]3Y,C55[e=55aW)d,FW)HP_X)IQ7VMIOJcFC9L67C#_(7>.QJN
Y/PG5>J+JFgcDCPRWTOX,=@H_f38CZQAId9?VQL[2Ab?@5J.7fR2L:MeB5J<Ddc6
BRR.@T_C3E=9Q>VHVX;W+dUABC,7[8[b:6RDd9N&O3RD;7&98R2O56IHGgEDaF5V
?Ca85NK((9]I6]?gV<N9g1UJ=WIc:K96V\TLZ;(/C)4PfFVHV/Z=DF\EbEc1+Pa&
ECLNE1P641+Nf[-J\)93WGU/_-U2F5)bd2E?M16@:K+#c]W,?H=P2VQ91c#Z14.M
EVd]J28_U:C7^U,20g.]2T#IP+>TXR7,SVVJeY9c1G-d=?3HO-YIe3R@N8;<7KNV
?-b]HYad:BfRUN>C<O]:/Q-(=9Gb(6+OL7bbHN7YfO(f2[fN)GTJEUV\27^RCM>)
4J5S,\V+7+)5&?2U)aVb<gVFVCKQC)B8egQaJLKL8)?]=RGC1<850^19E,&D2Z7S
LMQ26H0G.(+W@ZBWGMg94(dOF,CIF&2_H:]R>5^X.[K/M4F.T^dY0L0(\Y[\VeW8
?.NYOV,b[2Q>].:L-QEagPAP;56WVYL6GQYZD].HVDd<)f,QZXOOG:]PRIY8,dCG
Z[TW(CQ(E>1PAMJ,e(X72AYY3F;H_E+\&CbBKNG>^J/R)J/,C.O90c+/GBb7&P4f
_MZOON#JM]M=#)g,@Y:fDc.TYPZ_Ma25PG:L\^L_4aLKKI0]dX<Gf6WXeOGL^fU1
[a^3Dc63=^,_KLSU>BV^WP:<0UFH^=)[Z1gR-/XRfXdC=99_-S3)9/](:\I+9E]b
?aaFYWVJ?e0MX)B^W->[Z#-X#=[<XgK(9geDc@C68YPW(FD2-2fdYMY7B_D[DaFc
,^E.(VLI:0U>PeYfE9Y7^F>NSS6>B15AFZa)RAJE[K\aO1[OG^L_65&X0de0F=2d
6H9&bc(PQTQ-/M[1gQ_M5_8EL707S;K_-Za_H0IE1\eN74Y?eHFQ9#5KG<81;61Z
B\3>29X)4d61?<9@<f>d@OS4K/VBU)GbS\YeNe@O5S..__;M(Q+8C+>b+aC]@HTZ
Z-4)b#_H9Z@463DV^QIZXO_;4^TC.=PBb8FLcQB&>DF:ZM4ZeH\_g)c.E&9dY&+.
P;[>2g&ZM@a\M5ZMd<:XCGe/\_C-aY\8UDEGLOf@QQK1CG-fU@UNV^V27HFSa>W+
6C]2c6/1<dbPC)1)9FVa7\QK,>V^]W1R0&B7U0WD>d))-XCeY1[()Yd,-[KL^HIJ
f&+EV1;6EI#fLaYL<0Z^#)K(1^=WFJ(B.OQJM>3gXE=]HfFb(>-F?Q_Td#X?JQI&
<f9LEM5#Q5S?-TC:IJ3eVEAg@4<_J27Cg_6=eBR\&M0eDXZN.d,;8?d5J]2YKe0<
dLMZ51>Y:ATYG2T23V-aHCE?L9J1geSG(M@0R^fVQ\@g-\)W6ACSC-S[[:(2>/VO
Q[feSRgcVbeG3P8#9O[LQ2G]\AHJ-<&/L#M#Q&\Md_MG57]#=bK0\g84A)N6_C81
3KLSG0<#08[,([1RO^Be(cT>>>bG[W?Y96NVQbKZQEQ9_M=/9UC+E@^4DW2DJ@c/
Z_2TQ._]d(bIG.C^gV>0#E9;>_^bLS;N?7YKg.RE8L/<VCI90cYU+Jad]_/M5T&b
e-^]],XR6\ABdM[(#?[#H)-TdC?#N.6N+IGXc0g9ENL^7d5T_H5L18R<Q3X#V7U=
+46&^R1d/cUAc;SN-REg^Zd9]b>QU>6R1M1Rd_\3GS?Xgg^@g@c?VBJ+HRM1I9eK
I+c,#])ec?E?A&5e^,5b(ZR;NQW+YL&=ZM=O0.f(f4EW-7C??3]-ff;O\R/GI5)J
)HbBB==bC,>54XDA2PI3Xc#eARU_&H;.TCG><d,7CV97e6/VAXD.V@\,Z5;e<157
<^eN9>1eGSbD<=FZM8-(d,T(@N;QZ4]EGDa1UZSH&f3=9K.5E9@,FA=dc+ZG;]H(
B[cG\UU&,24-a)U;I/Y,DUB11@[d1LXHZ8S[QK02YHH-I5MCddG]+PN>UT>:R?Sa
JX\7eM4:[=6^H-/5A1YV<JTHT)HQ(2F0Y-R\JT@_J4)g-#Dg4A[>SRPR_G32?RE^
<VR36#.Q[YO@^HQ-S].1a5-+5.f/BQIXc=0NK0P3K6[TN?fa85&_M_A1gf>,27I_
eM_?&B+HS-Vfe7.8>M[<XFa@-&e7CU[7aT2&^_+^e5F0JN?aG3MPgL7W.4B[Hb#1
]0b1BHcHE(.R3WaE:B06HeNFT]D1I#7#cKMb9>-Y\Ld<GW&^c31b,T7bBDGb1W.[
TL0CN.?Y040[]&<cBD(Y#)(/?AU9GUg9[P8_I31Y<I4?TE&2#+JIM7+1aHFUKe;;
g7)PC^+VP/T=ZbBBFg2Q#SfNA]cN?g@UH@P_bWF.g)BY4H>#3[JMbGf-NJG,220\
+Q5)<R0602])S^B1D8B:KNFLLQg&S/\..7Ng[QVY??^GO>0>5;A,EBGZDT0TYCX@
F6\L8cOUCJ.,5,5ANGP[0K1J&<e^HI;B2d].X#6I-)U1Bf@BSEB8I)-QI;eFMa;.
#5V[[<3^+FZNNGPJDK<<[ZS/IPUbG,^(dW:5W::O3@LG#C\]6Q([OS^E4(KR_:D9
[D=B(SD+Qg7#5&S8WX//Y5Y23cJZB2]M+4A=[P:>NE93O[O;^+EHZAJIHA1GV4-G
\?eDD+c,]7TP>J.d:3\Ff/4)LYG?\5N7UL_1#N0>B?QTafR1Nc(J=)+0CN5E5GN;
a+U<6HcF?S254#R_9?.XN_BIU#=R7)P/F<LPb1#M=GVag4/TaMO@<N2=3R[:A)95
Sg/L[-#JL+)bQS\CKPbY(B#3,IEfDA;\H^ZGgY)UR#P5D7L42C#\F4VS2e[:_EK+
@P8LZHJ];8gP?G@gY>[aWE2H^dg4gB(Y+OPc2@WP5C:FE7QA]_7dOf>=_[a<AR)(
Y?Q5E,=9AUU(MF<6V?E(5J_CT)_b9A@66=5eDKES;aN)R#4DSAVW1.G+;OV1Q7N,
ZM7e9+;D@BVM@G>;-.V(&BT,9S;VOR(9LAR3-8e-D>?cE1bfTf,4GU-XTf4Y<@Ue
L2.[S]-,<#GXOfec\6CP3]9[)3d<.Y<2)He,d-[D4:+:2JE0Ra1-7b,Bf=/g+V+5
[eE\^EMceHBX;KM#3HAM;/ZTAgdO[Ve8.a>1ff8@T<Z)61H:-,dT[5b_?IJWK5&F
3gFKV8=/9bO?7XcB;dXYOIU0G:_V1]2@33&AE&,>@&@Z^/F24J^<?K(MX-5,0b7f
WLML7&dKcM;7)Xc3FVJVBe7?H#gdJK>UYC_AeV.D:7SHQY.WVA@DQgZ0>^E5+9S;
9ED?^Ve]E6=X2e:-F@?7CCdP/T<_X//HV\YZY;@.:T-M2[HK?HQ4#&UC8a?ZU4cc
DVb5#Vd5PHe=M.gI7^TfL;RJ_b&/<ED^_Z+#=38DG]Eg4IBe:(.L-M<NX0G8\VCC
R,(9.f>S6X\b&.4-=R?89SD04M\2HBZbEg497\Q9DaP<_\I\(5Y:P(aJa3Wfa:VF
^[@C(P5Ne<+FN+]QA7UUX:Eg(JBOO>OS;-0HD0Q2\cE1H]gMD&V2Cc]H?MFXWV-C
S0JZK24O1J(WI+Q2L-JS()0T+\[N^cg\0VBZbXUDNeHfYEg9-\LSd,DfLS-O_b33
H7aNJWYUUL2V[LRXA7PYPW)gUJCD=(X+bUMH3aHaUMgGUNCG0ZV>\bQ[=.bHJF_,
8BVB-L+P+,>\SFT0(W0XJ+FeGB\)Y8#3^O)DMaDN)\A^P#IJ+I=0LA(c-a+W3Vc5
dMFZgcQ@ad6Q2_dJU1@5TRMfT_]&SAS6&_FXR=U,4SLcAN4Z+FGHY-R8Z\(93MPM
b(^=F\JZf?6cG_e+74M06V+/_:&44.I90A-?F1KKe>cGgJ5^4SX#-G5I;QR(C>8)
(U<:5e??(<7,GQ^d8_WRO8K^/T9]_&,AfeQY1I1#&IIUHX911PYD^f7G^cf[[3^C
TfH@3S+QEC9_Z8[PCe+5;b[\G]#G-,eK,B4+1Y72S1:KL^/Bf(F93H[-NHT^KU^2
0]ZW07&XcZcJHF.[\BY/FcLCHYL(^9&^P8SAda]RADPAY@\Z;#HZMd/&PX7+;F&<
9B>:EM39]6g6#&D.-6;>I?1PR/_dH7IC@A-#V@[bAK7G<]P<X@>D[5^YZ,A,9aJM
a6^(CAETbB7gMX\D0e=[&O1S<0SM@Y]JJ9b^7:#eGLXZ1dGdM^,Y3JA\Y0(7NW?4
b3eJOA[Z?,O]-P_=>edIJ]^=d=H]b_GA<:94H#&g@ObT)D/Z2=R/\ULVbS@&4.db
F-#\-TB<^9?cU?2CK.>1DXN\6bF(RU3Z[E,XY()D,<f9)6/fK&6fHRb8==ER4eRU
[_:@?6TIg1,?36_\-_(R9(P??YA+R<@d/dc&?@NVL42V<?I(,Ae](0g()M7+IFI.
YP3W8DV8WE6DR/U_=&cD<;])bVM6b,=B_V-.--3YP>ILa2KZGK0(aVS.[g#?4XZT
,700V,G&7FUIe4f,GfLZ9a<K0+D8Za/@P_d@252>XDZ^0QK7bP[@Y?2>/Y:fA^eR
.MDe#<MGP+&Uf&VXSM)OZ<MHX5@cWM=DaH(O83=K(-0.Dc.YFWJ:O/@[-^3AT\gU
Xd47_c<dfC>K9:CIDR@<^WAe3&3GF-c)aOO[R/]\/N;]MZ?)&R3VT,3EcL.9&+\F
XE3S26U&T/+ET9(LJ]Y[d;0&_S.Z.,YU/K)1D6cV>AdGN)#,X.)Y^)@KN_=C7^6\
_3#a[=H@XZbJ9f1Y2IM6;9O[H8HQ/:E@6]:cdWP=-U;R9UUg2/(M@#gY&JC^K4Y&
RBH-.6_@6Fd[0<bKIRcYD7E?)((1(ddNFb:Ge<TZLV;DGZ)_BKERMfdH/C)]b?AE
@bg2J-c]V[Q:6U@WE-\RVA,2::2K03+fW6af0C.QD=3IZ\Q\RP6-VaFccg+J[4=C
Z4Z9XE;#OfZ?[A?N=FD9,Y-T5:/^29XL(F6R)@T:VC:M0W@J^,2)[PUCAGKXOZ.Q
6bd.,><&g:cP/+NC26B/d96R5C-A&ee0-&M6Ic=\I-L^E27669&9_^,;9&#U3GI+
X^Ob<8Z4_48OAEV^-?C8^P\=OX(E1K8UTT2NNdJL0_5_\VORJ_I&8<efZ>AD1+Q5
V+Q];RcgdaI77E\d-^H<<M;/\U.-E+)CLa\<,+@K=_9Z,X7W6M&:\R/5E-TIUBJ^
#^9TIT_[CUCT<-f_>Pb].f=0I(\<+[[,5ZVS[3=Fd[DDNCUEdA_:7;,SY\K.YJ9a
b_BE)C&P#ZdIN.T40.3E&HD=R(Uf7^<e&4)O&JJ+&89-Bg^7e9/7D4&,Ya#&bG53
YNFX9VXN&^bV<54B5SY@HSQ_L.C>043Y^5N@(T22c7D?Vg08_WA&^>K;E+29CQ<a
/4+L=._R[<^R9M2OBMeaac\e\)G_)Na&>F79[a[G2d6833a88D[\0SLO?8IPaTX9
R973@QN:5^Z;89S;\DG9V,aOeGWUY1J[;Q>aaf[b<6<e2BS,6IT[B#T-G?M<@TMZ
&Ud3;0.Z<A031UXBVGL+Q52E.:KDQVXR[:_YT]L5H<O==]8P.=8)Md3ZOe-GFPKV
?NV<0V=CZeT3#0(A,bBDeX5da=9_NYAGX-#a>M8^VO][FZ?gGa)6BRS]F:ZV]5,^
YD<N\A(3Z#RRE[PYb\<51^J3f4WB3P7]V>fDB3Z&(c=P:(\1FK(DcM)PX,CPJ4_]
@)OBg4d5]#f@9SR.,7bAWU2./+9Z3.H3^D^S53Y.b(?\:8=-1Z@,Z2P6M8DC+P2:
)=IEdPQ;WGZJOE1>9OPaOHFN8Q55MJ;LD0@SE.2.5K-[8A5UbGOWVZB2\<.BOVJ4
-5/+:cY3YbRKEO9PAS78\Z#&dM4>dEN/A8.4FC8a9(GVb1S8[-TE7;K_QUPf]HEP
;9_6]@bPK<b@0JPL8M\D#;e,1FYG/<aIPV>@=JS?G=2@DgUL^OGef2C=d^:HB\2A
]L-HPMa_]HD>C?Q-T>?+&6S)O[TT:)_FK-WAZVU6F>3Z&H<C)_gI+V\c.g+G>,C6
bHU1dd-83R//G@S-,dJ/T+GDYa#ZAD-W)WL=C5SSUQVQ52#8L-<EF4JWS-V#/A:A
2H<bKR.g6XZOSgSd+aT,+fT18OI7KE1;BJ_LUV&7P:98HLEZ@._0J9bc#Kf7N4gQ
?0^WcO@O1(^Aa9f/+&V[P4X)5fPRCMMEed_fdUa??])?&^M?1[>H51.DO@?VTT=#
MV4Ma8J>KfZEc[@FLXL5MfS5B.4/ZI/d@Z]2&)Z<?CRg)LW(A:gf.#DS7OcXXIXK
H(U5,bXZ(.E\Y))@C9+A+ce=^9(U8cZ^V5X1ZWIQPH=V<@&8-ECXd]5A&?T6?Q,G
YG(;_#(gIRWT/>U0IFdUN,K7N:@Xd.CT;2QM/@OFW#Z]X@O;H==9_O7J<VEI<S+8
_C-bH:VMd=,4TL)b7RBT:bV]9NMW)eAc1\C28^&0B?8aM]?24<:<UD\e?faU/3_a
E7Y:PP<4@)?BANC<DH;#CDa>W9J(7<>J?(Z,]7+7OX#J3#Q31Qfe^W#01FeUe61U
,4<H@Y]Y6V+K^D)XXP08X/2(HXN-e12SH&/3;N(cW(0W12DIAJ]ZMM4cR\/)^SfK
G;;8-0NK,A7==1WSdT\DX<Z&Jace+D3;-B^+OD^,91\dM(43@+R<Y>GQ./aIZF)P
C1\<b0@T;3^f2Y@#E_G55LMSgOO6ANR]6.1?[F@,P#GVb@VTMc41LYUSQ)&Y]&02
?3UL)LadbLSEMGUKg26YV_/=UgdRe.)GE77D7>,/5;4T;BGMU/M:9=c.)E4@f76E
@fB#D>_;dAB3R>T?/=MQHT9,H?>Zbe::J4;.@b>OR=LQ)<gES^MN66K6a=:3I0(]
VLL<f-6IVABFY8ITJ#>0HUb+GJ63B(/]Rd86FGFYb)4)PBe2J3Z\3HXDKUFYAYM+
L6VL-b76V_Z_[I-c+7PVL8=9Y4FS(A)N-3/V@FW58DJAc]c@b&-aQ^4C#&#WZ[(G
B=8g5]9Z.WADTL[cT&UXNKaa,M\(49^6H8?0JHSfNX0\5>WXN.#bEGX53)O-,8gH
K=SF5O7CO^BT]_fA>VV//I_QY519@O&C4G)/C_HGB-SQS-._f4,R<WC2QZ0/J/&c
LRM>6^fQAWZ09P()e@CK-:RWDH7<::YIHb>+I/P3I21A4E7M\B(:FeU>:ES,S0V9
>SYHX0QLX)30[4M?dC1#3V/d)7M=NY&AN_X<1?]fFg4C.;\/MAN[S4F]ZH]CED#e
NgSA^g0T28+WK/77aIRYH4BbSVf,@_eS,YS)0\.bL4RJ6C0&a99g[c/Gc(V>H+_<
\;fN]PQI.I.<c>)@;[N(UgA<\9,ZNc<;+/HOcT#,:I]c5[I+;_Q?WD.OBT/X7M+4
f7_)c?6=-&7K]@_f9@AQc(Q2W46(O8Z)+PWJ>;@<FE-JSP+Y@+\N9_XXYOZDVa/,
28G2D>1@Q[Ad?NB6L59O/^IEF=UFPb#&S&][U9W;6f#Y?)#J&)T0AVB=+>7e5VTX
8MVgL=g\:58HW/S(K^ZV[RPcQS9;3G2Q)O4+I_X<9<]Ecb0@Y_3;g@Y]ES:_GE2[
FF=)Mb<W96UB;f6J;PF1_?NU=)[DBWF;P?ZJ9)U1THU73@J)-ZL05YYF./YO<KZC
XWASf71b(\O#\H6)CXJbCW;G6^bB/2K?4;D=aM@3XJ@H<b<401RQ/X8MLc^>7,TT
DCK^YFdcFQ94Af-Qa:fZF(<X)@O_5H1/fKCc24K;=F6Q0CKY)TIA[)Qa4?]2ae[#
1f2cG\8A8)6RB_+OWIgP:0ADa4&TA0L;AdL:[<U5YRg9Y67BK6NK@=]53<;HVaKI
KGd1?FgAWMHG?VXLO,IYQeMcKN_0BQTdMS34+4@eL8^_B5?#d,S,0,NTH(W7)JO?
A_&&IU8B3I9JV]&(2UX[@.;fFTRdKfVQfFV_)gN\UIXcde512[7a59abQ3gQZV17
Q:_GeG\D^>Y9IRde<<U]Q43(>NF?CE)AW=3P++GR&XM/@9Ef5Ld0dWG51V?b8(]8
UR@B057P]B2,GV+&]5E4U.(M[UTKQ.HDa&gCI3]Sg\NDH-D&81F+.3I:PQI97AW,
H\_c(MFW.5,P[D[bL@K\?a#\#<AfDE9BcKG9+7C(Q?&I6+5=GbUU)M6b&eGD_PKF
=5fRgN>\IO<?<1K_RW,ST_Q;U6^=@I+4T0V6^M(.[OW(&_7LJaSf8X^6R(.0/W4?
FVLaIGYeDLaK\fDI;BW1)\B:N;Be\TX/cCJFfTd9[K(b4+E9&)<)F@U_=(VX>BLB
SUZV;dP,cX5S_?N[F6\c?^Tadg;a-G3Z/#fG:HM8IY9>1>3+DS#+=PU+2POFO4[O
5,J@@.RIFBKI1]_0X=:aJDMKgc.DHT=08\2X9+J4DLZ:f?.[=:_bTRC(.aRR_[U-
>c]46B2)4IH]Z#E&CEB4BFYcR@+@_B&Kc3d,(K,2I,PWCYJ7\T+dA/7GdfU=B<L4
0-X&F(;@TgbS+H.(UMHWG2_G<8U&(B[V.MNP8>Ua4J1:3O]G:7^3SC/KAR1fLZcI
eKXU9Bfc8P_P<5;905;<CWNV4e&I)V:-0^G@9>fXc682DU:JXQ4V3TS7fN=R6^Qa
Ig;LLIQ9V\<7<XdaJJKCJ1GYb@VL#>UFNBGO(aQ&(aX(SDSbaZD.c9&aa4K.?RX&
e6g_5f9X(Z9>,O]eB++^<QdJRLHgQR:G?6>,XFBcRc-URG](>&4</7)@WbZ;5CeZ
X3@ag2B-)N,18dC70b;HQR16]/D]6/?eX_(]7)_D54^#L.^XP])K;2ZV7cE5XHg2
FAIL8aH_J[ES^Tb)O6V;3/?,5.FF9OWS,,JaNW;T,a\IZabX6<-WJ<_?61KK&:C.
83=?4T\,;_096P:9QD=^Z_34CVYUFCKL.aCP5WXVG+^b,^9#:RC(C3;]&4V=QQCM
Z8WAXS>0bT&IH392MC,NB8Q+K4RI2)^g>]I(&33.3\O;](3&J-<=3TJ5R[b3^8ff
OGR\0f,^+L(PJ:5]9>R;/\WWg;549)ZG[7?M<_RU5Y5[X[JTMf8aI,W78+KD(HJ[
QSgWS=DE3Fc^;[G:+X35^BN5Ug38eK4A20XI1De:cdQRLa6\LYO^H(Z?6MdKA-7;
Ua<;_e7@U23YD^dNK,/V-[EY/.SWD+UEUF)gaBMRO0E5O3N.)<YKX,T9U6cZ\Vg8
3492RPBT?gY]>eK0B/=0_-b/L:XF]^NM.MBH<(.-N@9YNIeb.R8P)4&VNX,G[e=b
YI5G5ZF.K_PN:&U4^fB=-a(cVYQ8929bU#7FQF67JZ=faJBf2Q#F_89<#a#R2JKe
c@A:CDd=A4>cB:;OL\L2^YR\\MP^KCJFOF-@&8:/GZf<OJC3(7LK,(7f^Ma(O38K
#dbE1^0AIS^IBYTZW)4O&-R-B4Q/g1R5SLV>D[-=KM@SGdI5-]/,2O8E-C-:M2dS
9+gHXWW;dA;@^HbI?->E]&f7&DF6/)-4LeWf6&);EDRaL(@5c>[&V]@(=Y.49KM]
F^3(XdP2U<C2:Og7H>)X?QD<?AaVd+D=WfX.3INN+6[SG(1<?N_7M[CB^&CEU4R1
dX@QKW+<<M<,#S\X.\+=/46ENN<>920E(@E]+)_[\U^L5\F>e]+RIeS:5f91B^NU
CZRA]9VGagVW9\Y=L7X5U,N4c08SIY2fY:(/<W_XI#Q9^,cW9b7]E@4U0PJOER/6
ReVTT?eE14b@3R2CYI>T.1ES>N--VRL&YBbcFXd_RNJX4-JF4=&5gaX+_DY1F3dG
5GF;eDJ+C\+g@([Q)W=W=K9E.E),3H+,J:<]g>EOXV@.a10,bgKJ7YZ=@\:5d.E;
a2,7UF)AH?42F3-,:YG#V7F&QgZ:W#1EX>LKOY>>A;Q@FJ9JU8PaW]5MPN@=WK\=
.AT&)I<^e=(eW]#5g<EGUOK7JLPDKfP#^835J(ST=OCBDQP2&1f/(53F7BAUOEgX
+Bf9G<ReQ[T_:,>5#X,)fR.ITf-#O-COb#9G^\W\=[g2]]\WQdgOSG,\gCNc4[Z/
G[+5A-BK38VW5EU1I4)3=F@8.6e&f6N:\^.N-&HMSg>Xa9)W_H)G@CN[\Z5OQRY@
e;Ve@gY6aZ=AfLDG_&63R6-/<M>;AYS1D;?cLIcA?TNVacL63#@XA^UXcS3NJ)+M
M)3Y6;YM@;B49OAJFJ:C=NIH&gHc(AILGDQefTQ1,@<E)J+JYT,e0FQ)@F?XQg9_
dO,SRAC2GOWZdRD,FRVGY^W5/@cUF&fJU]20Rd;DQ;3K\2?;DG>D?@X>8-;+WN;g
BYK7cTJH2\1&YDC?;_\EQNe0H6D9E4#QPP6D[.K[IN^.Y0K>Q0SZ+g&1gQNg2JUd
EZ+X+AT\BPZX)fV#S+/C/VQ4G=9g/)5K?6((_HI5ZX^1:VCc.QcP462M-+fA8&UP
)K2+CP&PdXO>^Ag#]XcJ)cG+/;c\LN>6)/2D37B_)D_O9e),LEG779:S=U.H5L&M
/TD]X0(3?7G,4]\Lc9_N)NgL)PaCT@I43K).(81_bLYHYS7LV3;J\=^Q8AHI[1Rc
2C+J?5N&]JJgQ3GS4YTU9E=4e_@f8d_3XS.G>R_:@5FIN(:F[8g^FcbDRQD/MaTW
c55D-e\e]HDaKF<f]G_9S3^AcU)M4HXO_F/[FX>7H54:g&fW2TF>VI1(7L4RC8V3
8S>D[M?C=4Z_X9D_BX:9?&M:\d?KTN(1S]@Y.AF7W<>Z>.KaC1[+-)Td2E8/Yc?B
[Pa+#,Q(P4cg]-)7[09M^Q)(F]-71ELYcA#?XG[](XgH9G-W-gE8]Z<[.VH2R&X(
.B(=^C__&fJIO/:\H0eVV(Wf>[;MMQ^K4UIG)c;BSEKER)6a@X;7M/\?aQKC.1ZJ
[L<;XMEQUI:FA8([J#/Ea,<g??eL=L:QW[SC;.C[0]L:@fBR7c_T.b5##UReQ137
^/<JDWP\41CBK6QagC>aU+8,Sddc[.>bGH2IeQg(ZL;O2K(e^5)KNgEAg4D3\Z?G
eQ.aDfRG5WaYOYb76F[a)P;>59JL9Q[CL5=DD-A9]bZ)W0249Ub7ENZ&gQV,SZZZ
LK)0F&@)6_-B.N;7Y>K7UX5X=(0Xb#C73UI2d8+B[V>HYA:g](1CHB=-dU.46RaU
28,L#N8R0][D-W[gM@TA\Z8>g.TXC-T1GIID5SKADX:gOK]f17ZC5PfP6U]@_d^V
@8X;R3c,&IEaG.aTSWBHK_\/R/cgd;8P/X4U)(aT;:.OALH2[=:X#;M&TQEDVM1O
b?e,SW+U5O_L>:[SK;\3RINcMX5[Zf9XAS.OAK6fI9NK04>:g&.DC<F<&>:>#Q#6
D3dX#>dbNOHQ3]1^;7fIRQ=<D92W#BGRI6>8fVN3g0^J^ga0\_K-0&>,\]T:&/eG
KH1aQe=>1]HgMLMaa&SZ\E;2\M)J;26NBA2KXM,W(77=ID;Y@\G_V54,K[.1=UE4
.0/8GK4cUZBZ9PM]W=f_)=[9MG,U1W#aA+RTXN.Q.KFcM&),0DI8CD6QC)[^XX9+
9,4>QcIZ6<&,+B(a(NU&9_<:/81M<8AN_IAf>.R_FL9YJa&4>d=XN.BOgcB,N4gI
AIL<3CJg?E5S3>ZG.),/+9N<59(O=)Z1H4LdXX@\C[7Zgc)e,(U<0:+a,X.0P&^@
F8<OCE(8MgO+E7.C9_Fa?cJ_ZWcL9NI5:V]L6N:5ZJOb8Z_502ZH&DFRG1+Ha/ee
(V)^S>NE&?,I.R6LWSG1/7H7=5KUOeQL>U41EdMS_Z=0<[S_T]OALF]?MOX\246K
=N_D.N?G\WWB&=I?Z[M)]M7QW7C=9+GV@2])6J?+g)RdK((RM\G/^VbDE@(KCM7f
Z;9[#.<=<=E.58aOC61OV2:B7e8RKO[Rd.EfTJB\)UVAN6#J5>LfGFcfAOfSQ[^]
[QCSZYLN<BCc3;Q)WNH_J-BTK1/CK9)]?09FTY<CI0HeYIW?QG^W?-RBA-0CJc@0
8Id=TN6/^-Eb&g()e]NB>_c=&4=N@\U=fe75)358b_,b)4<)>307V_4/YG\S\=^&
X+\PTgWM1e,S>LL]\:,W/Tf/F--P^ET)TJ&@0eO)KQ]H.C6AbYfNFN4Z[QD9I,<@
RU^_#f;.YZZ)I<E_<IaAHE@[2Wa;a@3TT5DfPbFKaP:G94BGN.a#(f>(+@-g>,D0
@MI4T&UcGPMQGUG_U])cDe(A4]AKK2Q#c58VA)c.B.LSK:R<A]7ULJKS//-WUcfP
CNg0Z:A8:QDb2d24^?00FS:1V9ZZ@WCC0#C7N^VCg[)[/&.L&>[G4HVO18]+V?,N
NF@)?QWeJ.g=U/Sgdd18E(-2\SN2_AA?)J:(5&5^K\?=eCYYTD.JP)\60J[FcXTP
]5D^C^7Y9BdQ6XY_B[G]:MaDP57MHgGY/;@,^W#3;HNfTBYbTQ)LbGb_5]4]J[MV
a8I@T.N?7.5+/=GM6060L2?T[369H^(87EMW0?1_U7@IJ@,4E7AEgF_34]2/2]/6
AN:#U720?7G=BK6XbPS_>+1:)5]4BZP[6,UG,CC@G7[(NT)KIBCIg+Vb0dd[D25X
1U7:e-UZO>/53gALY;?HFX.CCQ<TEL,>Q\;.MP.IW7^[>5#G2;VLL]&,UEJMS4Pd
#6]JFLE9AA_7P@>CIIFCM/4<c<K4.C9fJ0_284RY:G5e]VSPb@:19KS>&fX>EY8]
;81=@8C0E1Cd>;M@.WN[7g#N)DeD3S^7L9B_NdRMFDLCYAUQbb6d,P03De=:>#ZS
9DZ[Ea9,f)0TIRNc1Z)+>b;41[CAGIb<=EGD;d9g(_P&W0T7\gI6WU?cQS#N91@7
OE\CaKg#1#716QRd&&K)b)]J:IEQOR2V^c/M_dGc7KFAK2e@H4(D>E?I]369AQ7a
I&6S)3\66NRe4,\I.4-NZTAL13+S^fYMRV>MQ\)aO\Lf4cAJFOa0+,X;P,WJBVIM
:6ReIFPQ:B(4X+ZR0#\NC\V-d8(^5;.^9(8gf@Vc>=(BRc9XD.?)(g[G90MZF)A(
P)I&56:/+MZQ+0Y_=OdUKHFbJKZ2\3-TH6PU^E\&L9:=3,>#Se1&-_&^>fPb@Q3:
9Y;V1,PG:IJ-9>\,de2:1C3H)7,V)fM\??c,0+gDX&.a?/WS+)](<B\Z;A/<M-]9
2#[@,(XLPD_<<eL43A_7BKB&g4QM.&H:#2dUYeD3W8H+7Q3(]BIJ;\SS\.<OTFK-
;9F@QeF;c,\bNU@5[3CE[/HObYI11K)^HN?&DZYG&5Kaf)I_-,/525WN?[FPP&c=
&fO24HC/SDEZ1)HaGCgeI//.?aWS18RR88IF\3[62PSG/e.2^UTTLR##8gUQI\P)
:(TaSY>\FL@WM5I^<6Q_Wc8g3:/b^T>=_fQ(-ZIc.]&4CT[@>LWe\=\BYA[ag.NU
<S]d[AJDR,+2HbH0O06B=_]Y4579O0JTH-FTXEX?/@WA6;WC2B(?U_[#DAEBVVF(
>WC.-PTW]Lf0(PE6A57+gQQ=KJ/3TU+(#751<0\X+e@/d(;8OY<5XBTg^Y3H;4\@
/\Z[I^O_YB;K5I3g?g)ILY6^g\/LOL&1Od4.0C\X-\?bM]&R-3@99P<_SbOA(1\a
eNK_.\BREBa4>@D.5Fb?b_^1W>6XB&)PIR4&.C[I.X.aDP>P<4#EXB,E_H.OfTeH
4ZO467Z3YQ<X>)g-6F&T,1#94-M.H)PUa5\=6/CZMDX:4AI(QASdH?^F,/3_@TM3
JPB#+RYfa_&?W.[SdIS/4C4O-_agRC/F[AU#EQG#IcSD,UPDcA\Ha3.Dgb7fPT:^
D=A?^b:(UQJRAM-;_aNW#[,_@a?JSd#cgCQI#=W((HLC/_-SgE)=U2FJQ[Y>OB5L
ge=+S1EVM@#S.e2V(FY_(]M\KC7GY#7YBBK3Cb?1g@cSQa4_MF^f-JdCOA5ePKED
#94QN-a:U;[/W#9BCg1E(\L<5cP;MF2AXHW05gKX0HIc0@N1]XE-:QWc49D_eQ@6
8\6368Ig&QI&AVPf1_If#;-/4bG1UNZ23EED?/65/+81&Q3C-K8OA(PBV\OTf)W2
Vba4GYfCB>X?g3K\eZHdN4BW70LZL@#8V(PT=<O4P]^<,f/4ceA<f7,Q3@1Yf;:M
:M0ZU0B83I2,fJS2KW@Re8F;@DW(4(8^XEdJ-7[XL(8_H@(,W3^AZEf(aeVC<[P0
^A_1O5Q26X+LFVDA_R,@\Q[^SB>I/A<FL91^+T^Lgb[\NSN8II7=:aPKd3.Haf?a
2JKCZC:eAHR(B0(AVbL\cA[LPaaX0<N57RfQ27=4EIe<8TOR846NK0VDc_?4KeN<
8YZ,dD2K469K@5=3N\E4+HE;fQ8#Yg3W:C=Oa<CQf)O(Ze1NX9<N_\FZ6Weg[]F8
EcfT:L4DCC8LNB_C);X8(F/Y@DRPZ3L8\d;NE?3dRHP9bWE4fE2#eNTMY6E13c[L
I19W5cOJ1Eb&>EZFHO>^NXKa\[@G3^5?HFeOAJB(gZ[D8=F)]c\>e?;bb-XfR/W(
U;@FAa>_;fHDJ6R2Yf/S8^T][P#\NaN&JWROZ(CN/&0])EMdd)KXK;[\@b(F_LKA
:K&bYbad(c(dB5dJYFD;Af#VT,B?.4IKId33f9[/81NW?UaB2;PMEN4-e;FZ/GH0
WW-4>9;-KZR2[]BFbW[gI)4:/7_S8X_0Y=(C9+CJ#0eI.R)Cc8@[d]4W<7_O+VKb
:OC.gCV0fA(G[+Q\ZW<D6R(NUMU<_faBb#c.Z1caT6K8Pg.B43T6@.\]LL]QDZAP
Z1[&K]GJ,ZW\[)eLGeA1((IE=)e@]&a1Y_HaD\E\8QH[G5RXCf#A4&[E<@JG;>L<
C=c3@cd8M7;f#S9?.L(f8If72E7/#CVVQ&<Kca;N_>CIEQ(FNE[6(_<2eG/HQ8_<
gZSe3;T/O\+cG[-=Qg=_QZf@#[9MG7S#T0@b:8[1V7&B.G-[216Z0Q34/R?BHJ6B
dZ2;Wb48L-/DEB+7?J=bS4IO<F3C_I@(\Z:=@Igc()ZL(CD](?]L:f6R,Cg63EYI
R7:f9?^>)?=8UGV;M2)1Z>d4^T[86-1[D6JD[>/SM2QXT(.eM07VN=F4-)E:H<:Z
=P/ebRUTK=J5,T),94[?#U8KPcP<^+\[gEQ0f5?f\NMG3QG]9@HMQe/Z6.b\F0#S
ZLdRU>ec>D+XR,^/ZJ&G):M2>#(DL^gOcU++PIeU&6f=Bc)BZKVP7O.AM[?)DFf;
CKHL/T1Na,2^IVJQ4@ITLD)DWd3NXNF)U<?;:R6:\HPZ\.)16P&E56b[DV0=44HQ
WLTV8RV.JHL/3>GR8>GYS3d?5f87&??&QMREcKJDV<1&Wb2:_Dc-7E=f#P&KK2^D
(X5Y,-<PWH<A:O\[HfEXN4B7,\MU(b\cfZ49M(CMYMI0.+MG8;&eG<4-)#bEG8#B
G\GFRd3#1U-+@.E/Z187@[TV/.O_7ZF.R-406H9[=f3-E);N[38^>+b<EYIX.-3Y
ER3816WFQY7OgdWcLC,;#X]<?[=P+GeYZ)@EU&KTA;I&,V/3LYI\KCHbW7A<CEE]
(YM1_bT<cR6W87?GZMYEW\T2L:+cTX<,W;/Y.(gf^d7<RDU<GGRc>]NJd><2XU7c
1=3=7@:_4C)\S4#91SJP?YT^R,U9)^[fdFZ>MHJV>fSP9TefcZZQ5+@P7M7]MJ-.
Q;N(D0d4Hfeb0DJ;H)LaQ#K00Q&;4YB-W[;UJ(E7<S7:1;^DZNg9;CbL:<g4g=O)
K<@g[dF+fR@;^SPHEgdT8M48YK(dB3e_C5+9G^@I_CN(:9O>bOdWQG^)#KfJMDN[
&\>U,+#99T1AC^=L/K29#dXD_H>Z4;<OY>E/7dYe9592fWN\_(QLE2aIK,N5X1DF
.?]?;<UfOe@7/\V)X)MG:2dNHdf,AA,b/F???[=D&GH3P8IJKM9JcM3cfAZaP6MG
#P;U>/0)8#6Wa#f(YF9VZA-DLa\K6?W/>7?UPS/YP(df#[EO,=32F)=9+-BK9Q&<
D4F,<g5J90.Q(a^]P.73Q_\HAbZ0D^c@??7=-d^KcJ4IEY:e9VEF8YSBOcHaZ&=6
fg:@;C7Y7)>0gEET07C0PR_^7M0SRF:\BNU<9Y:^ARYJM0Ze&=;5IE7#LJ?b6@cS
9XJg2_5)CYefU88A:/T?N)L)YM>J0FN;&c1F1O=7>?a@XS<S&^(0RJIA3[UY]F21
X60EaM);J:cY@7cAUPS+Qe,AF>QAHUJ>M<->_XG>c7YNZbF[SL&BSOI#Z-?80QZb
B/I_dO1UaIBFKXcM[ARRdOgQG]g3=UH?PKcf(0]3&LN3):Te[G8T:#(_c(;,1HR8
^.2F9:4MODX,gS#972&?e@WMUB9Mg9.XM&).49]@MIE_,X=aZb0ND[6MS:_bM=eY
gdO,[BZ<;VBQ7[1^RIZ>]dYQ=J,S\#+cbBFOL4cFX>E8#f\QfeK#.XRHV<9UZ<=a
C@MS/N6\#6OJ;:A[1[(@]ODeB.G,AMM^#QZY?b7G=G7CFO@-&J-#M]8F^XPMNc1B
0L0:<?6&4g@;R,0(cQ&bc+^_1B.Z=28T8_^IG8>a17;7OX9Y/H+Hd:G[1g8\HO3Q
X.d@.\T+JOL_DY:#-40X_DR:e//cEH8gK?e=I]=0/1_LXPfZ^#PB]Gaf;=5,c[^/
C[1XFd6^UGI(6f@?XQ5Wa2>Dc^=eK6(eY:+04@,WXN)#bR629BXGP,>9]9RVP9^:
7TD5Dg,O9Q9[cAVFO+2QYK@J3/84<c^\+_[UPQ8cG?5Rf?)+F3)LMR=NB-e9^3\f
)dQ4\6&HJCD2,=RG_@^MF2\<@,]?,W()>LPBWa:QDMG.EE4Id;64ESP,+_L[X2N\
dGa5bHO)1/C?BfX7Pc);1QW35(+S>b[]V:\b=>A>-D[TV?\^?e:4414?E&S)1J#9
JW<I=:</5]J94T9-4J)8FQdeZ?Z)/517c:_)U<d;2U7Y@B_NX,-;EJY5E,/;(>0a
Q:C83Q4XR&(A6;ABS0Ba36+dAQeB[=[-Z0Y(@1d3\d2G^E7BT66/;)BWPNCP0gNO
M-cV&-c@11K<<QP-2[Zd<e7,1J;YRIQ)C0D^U+,N-f]YT_3/#B_S8?F^D[(4M-=;
1VN5gTZ,[DVPMZgbY6^d4)ZW7\Z8VTHX?Z(d5[DY3JQG@#6.fP/)\_EPg>EKcH?:
L3+c4fK_M,DAAWEVH1M+>JISUCQKVfD&M[#X]YV1,X\bE-NX99S;^C6,C5KgEJ1B
F2QKYD-_OU5/2R>dVa?7Lc\:G4=B4.K;JH<2H^:IY_:1&LQEBCNG)+OEQAUKZP,7
AW+X/KXX1PeG79J5JPA4SG-&Lf_9^5)gGV(gQF;LeECb=G<MNfY4LI<5_<R3BCKg
TNIV?<eZY)Wgd_LXFK6aRadZBg+;gd,-_g(8HSY2P?9A>M10>_ZS2N74Ta]XBPOU
?.d38e(+T(Z+#IT<:U[7+<.XLQ8)K,7#G2+S.\:C2/e5&,A=M5MZ<3eF:^)I=01-
(IA;HUYB;E^0EKD#/U9@&g,NIN;-CD(74R0)C=dZOe_7P-4Ja?0A\KWf@BSUcHNO
9>E53eI(6C4#,f8LNfA].;L+9Q>+E+&6<3YL9DcffU_OV6^7YbSdXW)?8.&DQJTa
;Bd4+DE\aU2gb:4ZK>DZ(ZDCe^#f34WCeA?Z)I+I-0@bQ+[/M3<=GedEAMg.Ig_9
.IID=N<3>4a\/NZa71)e0/P\9]^SM9QEBSaE6Rg+3/fD(Z/4dO?RL=fCG;bKQOfc
S[UA;6dJ1&0c,H43a3gWFW5PFH\8<U<SIL[SM/c+[R\E73.47#7(T..Z5]&U<+]:
LSdV5[c;>1g>-Y)J^AT.2B#0E0PHSR4[2Wf-,U-^C8f;6MPSg8;WVfQ9)0[8P>>\
afNN:&;)W.DP5X-;8&C[:K]EL->BO3D78Fd4UA\A^bEK)2<,VYeW::0)ZQ4)VLE2
GJbEa-;CAbNbeUc.H5VIf)aRY#5/WXJHHWR]3N^@(cU6<.IC35]?6]f^dc?_PCF+
C_,24V&/ZETGbZ(Bd1A7Rff(dUD;IY=a(F?7KXAe0f5/K/TAB]8f<F@Ige-3.;)B
GE4^Q2TffR5\FgTSe&F&2\MNG]Yc0JPSTSg347aZH;D?NG]Q93d<Q7IC;N_468_6
0W)SD1P-fO5<TJK90IdM#L)&b\[L6_U;@:),>77K(SaJJ29.]d98PM<:.L],:3W/
.5FB(3^e64Q0MZ:6?4_F3LL2X=X60>bYZ5NDP>]/@=C.,A3A95=WaMgC.bF;6<,7
+QWLRJL+@:5C1GHZd]bO0WN:?5ISW2aR<+Fd4d_)=F_4U0IJG?e;J04Y/;M>>9V)
YMDOX5(WZ=-?Z0NYWVZCM_@G9X+9?eN_?RQP\2(?(K>7S9Rf2?8MKL;cBR\Y2Z\K
,B]8BJ#Td.PVbG\0bdF;00TS^[(HfG3+M\:dV>d3L93Z:N[2L)5.#U?H<LdN\)eM
2;8OE1#gRg@e#J>_9D2d<?,g8RBQ.X,e4fBf[ObHVB,03#X3OI8g?Q;VJ>+]G9gP
-R&.7D&;+#:A03C@d5B-,&A[Uefe?@M\31c/aDd,/HbMfPU)>^K-1\&EUg8:e;W#
,c<b?79#UJ\(fT)MA<YN7:#\US#\KdS#ZL96R-]8@a.V\HFL]^KH1+-f^U(=^QB9
PbZ8B_P2f4.V=0aY=4bC2RVSDBN9RDAgRTK9O<b=bSRQH_Q?-a8J9\=G7_Z86aU[
0A=R&bIA#II,F:@[XdG2=BY0OH1HK/YAF\GH<DLJ4Gg8RaJM4daNf/YBHUPQ@[7,
MR7&^GF2dM(a[eARNAbPb?/7c;V_Rf6@\;^NU?0GC;[;<7,UD;dQQfV89+9[U2O+
NEI6OP<D>-8D;]QWQ?bEFK=\4)fMec6KX&;3AaPf(AX]@P\.X>1ETbO\FSG<P[U)
f-)2da9e>.9L_De77McHKb&eSUS6=BXD;>9+Gb0V+0O=1ZLdYD_]4)dT[X?G84bH
-,aG1NXN:5aD8^)f4#]a<;KCR-Aa8./SP,aQTYKPbY01Kc8CB7P0-3&<VWJR\3Y\
ePcXYMg?0[DHc/g6<(YgZM((]gTKI6L#F9)T6TZB\-Z9a_+6aOY;c5L@B:R:B;&Q
8UT6)D21@@TPddET^PD0G;+?8b#==@M1[XCYOJO<2Y^27\.YES717E.QeU4ITR2^
HAB=\PKALF9QP:bT2ccR0;P@]d_D]);CY]gT4FN9X;eR?2V>XdEO/M6:5JJ4#N6Q
@[3^ac\-E&DQ-U(KA0&.(BQe#]-6J:CeGCdICW;PaGN]<E:6<,?-FHQ95,PTKJaJ
&d.feD9\M,5N)AUR)3?B_AZ&#8bB5:(=b?,U5U.<&RQ?1;E5C4_6:Ce#2#+c+)B4
;<A;/=d)]&HE:Cfd:OD\)@J^,87<N#:KU(^UF)Jd,PeHb>#@/#R/9b\bNDLO1Y)B
c(75?3c;E^,EL+0W;I<N0YQ./O6Bf3N?)5.6(HaP+6dPL<#/F;b1UWcL2c&9fZDQ
-=AW67^+WO.&1fRI5M.:?1BEg9[KS+>+08VHQO./.O\<>3Z#OH/ZY@G^[LL=<e3d
IZfC]5YH.+_-8LVH9IQH^JYGR=W15A3eG]+H5@^SJNW8SS]ZV6VYL.JU\CHFAS=7
\NQ/>3[ZA;?)PI5N;_6BgM0(<X+-A9DKC2;RK6I&a<cB56P,MFF6DFS6EAMcQ#XX
?I/2(<#<aB<J,YK52[C@T-,&.)gJAF^=HcHQ>8KYYP#KW7RC3E6ZF5T[EbMDO&N#
WF7W+]DX2CJcff;_I,GRa^VTIF943Cf&>_@NbV7=BQI@ID?F2.gDOW<AE1);XeW]
(9?e111D32&>PgEH:YD<(g=]=95TA?<,^[Ca:E#8JB3/-BA9<#MLW(Z9Eb4Zf>&L
8\BGC;&\D@\=Hfd)L0Y5CLT>L3+#HLGdNQgF/,BM47b-fAJdb.dF1MJS)/3Z_\]g
b0C\MdRI<5VQOLA#K>,X?.)L>#0f(NU#H><_QQW9N9JH>Aa00Y^G-Y>dUXM++c2)
\CcMVPa28#B_&5d6b:_>D_+/VKAKB:,3[@GOY.e1TY-J4GG\dBeP4./9KC9X?+=c
QZXKOaZ/J7Tb76(X;4;VH>](KP_HWa[P[/SL9S-XCM#EDa1f-YVD#34P0U04(A,P
EP0P-TaaL6C0?ZYNMNQFdB9=4?OL6Q>KDL=b&&Z(A,H(U,;EV8COD\R_DF?E9-RK
Y(C(+D_OZC,+Y-=TaN&LH.O]Pg&f=\SO;(N;]S8P:bNP,e).<c12(gZL/e7R9bW8
_K<XWYQXF0WFP\^-Z2+F+JE7&F9UZG6&4QFP2>d:8<2=NS>4F\XY1M?f#Qg?HRH-
_RJU0AAZGL8]C5N97GGH_g49@P7<eW>;#N,232/X0eM.>K;6.aZ&L?E,3g1AW[&<
J]/afdM6[[G\O&,.TN-V2Y\BO8,+,:D5CDa>gPaNLGS)NXKL#:Y8EK.7NJ)A]XU)
Q&&FXgL>E\gE-^--6T<-2E#/HF0.^bK5G,O^ESW9)K-K:&QHYb4&7+G&_+E\4TXN
#CLZaM3=Y97GJa]BG_1Z@0g8S/HNa2bfA:P6UdGM.VGS@+e+dQ#0:2Zgf(Mb/X?B
#Ma+K?DRU)P,aP4&.2cCL\F/c3#G\^gdD]+,FHDEFOK4f5Ud^a=d=_f7c5Zb.6W4
S3R;X#9.c@fPFS82F;9@V0(-OZ)W(^D:H+:(@6NX/Z;&VF.[CPNe,)\29J6AM-X&
4]7&Z+fQ=@A09:[/1BfFP_e0)Y:29^[86g>VC03_U?<:FbdTE:9^b.+^3SV80#HN
)DUNGQa^IK/L?4M.aZ:g1I4ZHU8>B#[OQX?7>OVR?3A1ZHI&UBcDVXc2UQH-:+?O
e/e.-P^,WcV2^bSI-3V<a)Z_XH8JfWa.gLF=.8D._f=B=A5?TU4BA_:EHQSUK22G
-g9gCV1J3,@Y5R>4.C18I>=55):X3fdP^@I+X<[0F6CQQ8Jg6N4Q51Xd;]GS>YU_
R34E(geWXfMK#9>cF]^#N8cY63\&8(a6B=8=O]==cW75&UX+5c#OUR6O#EAc-W?G
a_8b1e/e0Q6S[TQ[;JCfZ\Dde\NW^KJ_bQKZ[+K;HT.Z-=WG&Da<:RGYfG6O7(HM
AcR>F[AJLWga[@-L]^55L..a5_8?HQ1XJXM:e_e#0@O^:WR7CJVI:B?2&E2)>U0-
>6TbX,B(\[73,=BEaY<H^Dde4gQ7VOU>=.2Hf6LLe2Z(C4a5ZDWH(+,V9P9^#S(8
5CPe3.6(_+]G3&028#=eN74?baE)&#^5f[D])VT&U^e\L#@Q/-T#O<5YP&N;.4FE
1S^S(CJN;5Q#fJZR45@8<^&/;CHW)JZ9WU,6>M8A^PI[BPW,;JU/7:JH=LQ4];U-
+B:d2/C>cCKFIOIB:QX[B]2\ObR-6c/=(S12#,L<[dN6QBc#XC.I^A)Mcf41Zf.4
d8[I^PC.TKMg/0JQJ4>OM+QY-00<:a@eCHS>:ZfQ+fQ76ZHWA/3)POa#+MD62WLb
EGCNIbVIe_&Y).1)gJ=;MYaTC<TN])[.We@P+QTXRKc1Xfac+8\-cM,L\R_/,gU4
+=OU+f@5_-3RH:I;,_58;J5U3J7HR,VS#TG_#9&X>D\\^/[SZ^QTae-HME)&6:fI
,GW,NeZXAa3_Q&&-990VTJ65NK#0@dT51HNZDJUOO][=B\C^^9V_QQcI,Y;K2ZUM
)LR6D3YC[.gBC03WUVW.VUPJ&K&[JCC&&Kc^_T7[L33c2&A#09)a-K8M>?\]aR3g
[=2^?_1?/4R7a+369bNEgedcJ4aA.>/gD[:M6\UTQZ5(M+_:3Pfd2M2\G:54/?\X
RXL@6>eYJLZAf?LVF9>1-@\\L]AE789NDQ86#UWeP:.?b@0ZCd?^Q^LEK_PA6Q@.
1MI?KdUd,UKa[G(O/7T;;_YW-4+EPM+-N7?C6]0E:OW)GWIbaV(Y:IdYg7fF30e@
-2/OC_PQ6X8AU\.D93+<_3<BgT1P(7N>Q#>+Z7=+V8JQ:1WTC>?>Xb.88SFf#<+/
GCb8&03AY0;I_CU\E3Y-,KPegCZfC(e1?GT/+233:7BK=QH=f/_MHDH(CJ)S3B:?
0VR//#Ebd5;#4TCULLQR-(4<ZG\>3X(:U^d:=<B@Y0_cD4H682ZLC[IO;9bR>>J[
3ULUQ9Md+FdU?2gWM1ID,UQ+dY0NGQ^6T-Q4N>aGS-)AUQ(J1faMK@]PE,G41fBM
HQ+D@OD3K4TVcVN\W<E?S[W3R3HN^XODU9QZNIcW0[HC;E+NB]1]eF.8Sa6O50UA
-7fLD)K98Q5[9IJ3@8B<PbN_)Qb]M5e1JGE(5+:aWRI5[b\de.G;dZeF28<bA]ZV
>2</.M&M8/aTG]Q\d7KH5e22\XJKX0+A^@^2P;X=B9:+?[URJ02@Cg34M>_>D)>@
(Q#7b::S#]a.;E\)__FHLd8Lf0.PBMXS(MTZ#)Yb3L_]aS^H+FH-NQOa&HV@ceb^
D0PRZKWL77fO21X,gbA?XKJ-.+O]17MX7d]3U9A-V>>LN9JBF[Z4YaG)BeQcW=HS
)LTId2+e20=K86;+=.?7_MP#bT\20KP<RbUCZ/&35HER\c5fX75.a_Tb#-LV9#BY
bKWB]CKHQ>Z;EG/A]+6ZU]UCI#.J/>ZIQ^&fd2+3I;QL4NXD6+9<.38AW95]__a[
]9XG8C\H#ZF)28ZZdJ(4P/.<[+M^B>OPXf@9_:.X;?DVXZ?bUQ=HFM&NUK8Oe@Ye
H1:QH;85U#;?31cAQ><edT_IGRWM&BT2X[)5I]-D1>WQ;e/bOaHJ9+6S004>933\
2=a7P4bGb0FF[?1F^B5Y:;7Y<cRE?EU5K\^.E#4636)QYP@4dQU13IG1J0XVDJVY
3TY])S4&Y3/+(=)K)\bMc^?@3X5U/@c(^0gWTSZ#^L-fd?;UF_Q)Bb-AP.IU3N_8
[3RTa&@:[@DaQ7?Z^IM^G0Z59^N<&C>?^#F]CTd2KP/^J@0;71ETe5(edG^ZUeBN
e_\1PM9?QOB@\?cJfWF5U7CHgR8L<&C:1@8cULQ0GOb<L_C=Y^Oe<2M8#,,OO&ZW
d:_bONT5^Ve@9Xb(.+P7+=NeWXG3fQ2EW)X>a(-CP0P4F3&^+;5^Z76RaA^7QeB:
F>8U.[dbcY@@8Y+WQAE7^G55?W2NM^-I#[LE,4E_6&0ZKf4[,5J_\\YFW)df28-1
>JC>+9@N3PIA#PPId4I-cg#]=a#HC2aZ/=>)cTRSJDeM^_e[APBeAJ<d12fYK[68
>&@_/Y]6869/Hb#9.#Zd9@\8\A2R:S,#SfbA.WUOeKZKS\G+f.WWF3NP62FH.6VS
+ITFR4PfG=d/Y1&OEa>&M>+L4_3ERBKV>A6X&&F]5]Y9gAd\X]Jca4,JA.ADNg9U
<A?TLMR:1<R50Z^=(:=VN/6e0H8:T?;7+c9MP]?0.Q,W)42TD18[9+VUQe74>-eg
J/aG.)6_@-PA]\9)MgD:R1ZK]/_?-X=aT&6=c)/Qd3FPg,&3bOgLNH6?:&ebH4V-
d-H@(ZeRNYbU/gCAdJFV);\cKK#/8<Q6QS<+T@Q5c:)HA>3N#cHF2M+]N^gZE:C=
]W,/?\J_EJ.3a3XPF[?]cZLgUJ1Q3U^M+gTS@,<7=;ZHS,_e3f5gaJ.HO]T,[U?M
WUG^1C3(2M:.[TZ1EHG+c0dH<3LO=-9?aIQ[J@-95SaS<FH2bY(PB1GcPSWYW?9d
e1aNc5MYd3Q#F/I700D1Ebgf-E_dK7fGB1:783CNK4\d;bUQDQ)DZ.aYP-_RG(D^
7If7Na7.]OX)EUF38U+1eP2\P?C_\KC22dCcX@(1J^L?5:@gaPbePYT&C/V+2P0+
2HFUI2#RB3^&E9S?5:F3[_Re6WSB8)2C0\[CS@8[-VgMfIa<RTX,_KLd0gJEaD#N
Z0Ja/TLM=4f;Y?IO)(WKMXH4,^.YKL6V11ZB6J.FD^&19Af9U7>PZ((b3:^R>eR+
E6OUGGAC&/TS6Y;a,EIFd-&//B3D^#L_Z1E/YM)TgV&c)H7gC]>S5A60>TEaY>Q-
9=Ua;_<NFaN-I--GUZ+V.[.<Q@.C[RG60_<#?MSVRA49<YBd;L#U2(d]F(<QR3NJ
Z0ACb&B>_<f_YfT_4L,4,AAVDf@Q_gF6F#,2RQ[7T5NAMK9LXUNa]4,SDK32U?Wc
a[T#Rb;WeB]^RR6D^bSd6A1Y1^N/I&fdMW<Z<d<eG8OL.L]O_LB8Y(FHI&XE5J_Y
CTWRUM+RZYH5R.(>-[c[B(dF(AI;D6+]>(P-^QPbFS#[JNdL^&#,O<eUNKF5LH(]
2RdfRN^Z:\egKHDH<3SST@M<3(_R?Ga6Z-M>QPCbG>.4gDEF_XAI+T#b1c?A)ZV)
^caU=[8M)J)U=R7D3a\D0UITgD.<S+^K>:9gT^WXaU<X/<C(JVT<UI2R/F<3;#P8
)\8AJW4bX[DYDZDd2gZVTN>OC4U>2c[P2.L0dYN#;V45R;dKLgX,V9UC:<Y;IZQe
-A5PC7Ne)N<:\)B:b/g,W(HAB4U)]AYb;g#_;BDZ=N^@e203M#+<5JEc5e_4(Z_)
<TUBOfJ\8SJgS;\HeKgR#_LDXB5Q@,YY\5+.M2>]P?EBT4d9>[XJ.;A6gCE^H?AO
3T4N--FcH=>@W&U&g()ZX=-1cVFbG0J=<,P@?KA\3X+HBY#g)WTb0??4V]eNN>@d
K+c)9gHU[e4e[@A)#]F<(f(>;YO^I5GIc2D;AK.bX;\;+fQJH/31]aQ]F(T86,Y.
RJOENLU&AfccT:F;6A.V=GY?2C:2^d[Z-\SX[Z#eBM.1>?TR7?(A0(Y)6,[6Ufda
F,R,>1.Y3g.E6WRE[4+-b7f,^Q_N-N^BYCG0TLC7M]6Z\?O8eR[.K8]E#Xd4,C1N
X(f.D2\Xa<U)bS4(M]=9,VVcbgN>C-\/a@,QG);AZQ:X10WS\BV08LDPd2?G:V.\
-EgOe?EGgB5aCP,MIGY-(:N2UN(V+/]a?A9+D.Gb+Wc]@_PJWfCM:<=L(X.3NHV<
\WFYY&WLL6[c:;fB3C?=:C<GE&#fD(K(ed_E^Fd?)BSIOM;RDe.<#H?IF470];bc
>H7eB:QRCf9QR+&B3O,LA4bV652JDQKE94\I@O7EOV(.IJ@R5^;PUTVYXR),V=a-
-IX9>-CMQ#@/.KgT1,.,&50-LLYQL>9T/O#7\#Mb3/8F<IF@Hf@e)LcX2Xg5^>M,
XN6C>W#)1S)XILfQVC:[/V_X<B,[d[E=c;FW3FE.CQ#;Y&Od0&.74PKKXF+RUU<T
+,<]B)?,=bOSb>;_dSFeX\4LCcE/b=9)f<?_^S]G,\;Y/K0^bQL).Afa9(c&WSc1
,75.F0I0Ee:deL()^&TONWUL3R_8Y5UZGQGeOXWb8)V_Z&BZ.c)Lc726S8MTUB@-
f69d)eY4.bfdGAGI@^+V8T\d__OX\.SBH[]\U;=<NCL+;1eD:5,E8NT_(-?WaJ1N
gQ9WERE+@5A6gGN>La95e(5AUcN;RU0KU\2Ag07=UAPRVS-Nd+54A3<H)FV&MEWU
>EX7fPIgWg::AGT;.6;2^#fTNcWRc>.(]UgFNC#._U&)PAgaHga2Wf9L3094DQ<,
Q\27McZ&;\P]^7Kc97RbKF9^.VALC25V+;X<G&PI3:JECO3e5>.(-A<bP8P0fQ+2
FEcFXV4g<Zf>O:8)e6NN=6</BFW@?MI@\-MJMU-dU94UcUN7+,4-;J7Z.dM3K549
cJIO@-X_6/0LcbMAN&T(N0QFXM4dX?G;QB?<6KK^Xd=SLPV1;2?\N&+@:OIE2W7[
S]b6M9<PE61-RZJPK>,aNgcYB#,)/0<0RR:4Cc;)];GF2T-L)H2#8eQK3\<Z^7[D
fBEPLG3ST?_J=.AYXR>\dSD)a0dKMVU@-b+670S^SJ^6#H3bT2W?,g)T8c[58#4R
_8J?)#&caMa>c/,f9RgC/H6[FOG#OJL@1,@4Q>07JX113>B091=EERH7Y)=W+6&W
df(2^TDPUB-Q(ebIAGXX;<O+]gXM>+Q>ZRT7BEM4V]58,I8MGJIdbD=fX3;BD3M>
FB.DUe<ZI==20)[CJ++c+T>9;;b,W:H@7T=G@,5.CS?9_(VTB^YU77:B&/(K8aCL
^Q\F5KE2=,EG\;DZeV1V&,9@\3TL3-01OHR?F>OWM[4Nb@LG/Bf\U@S:]4e13YB?
P6K<3fH/(2_\]/B8=L1dbW&A>\SCE<1.Q#DH4&1Ncf81@>7cKGgKCIW_1ac73TE7
\YW^Z1IFdBK#OAI(U;@1F@G8\GNY7X7[94@AJc88=<4#^8?20CN4NNRDJ@4VEF<M
XAJL^3W^aE,eC-S21FY=C+)IJ47[-W,_?+dR=QA<HHW(Y#K)IK^@a,58[JUS44gT
I_FaSf^#bT,^egLNP:A+2@YJ_cYGL(3e+DT@0[e?+72JdB^PVLMcJcN4QZX=5J?U
8<0(7dC40[75&03aGT<TX(1NNcC.8,4;3KeR?S,b1/MR:.B^S\b48H/_Zf\UKUB=
b+TL1^;=<#1O/H7Z&]<UN[TcGD)VOJ54848/bZA4[+JXP6U/dN))+TA3\2/J-\9P
?WFVAIPCK,&AUK<X=;9f2Ea/_N#SB.15[Tc2[,B.KQYGOHRDb;9R>6;U7a,HV7N:
-L3WA9d5X#_I-W2LS,cB.QJ=;a-F+?R3W+D8c2YQXD;-I?<2b8,aJf=MeJ/.1^VV
d?T4O4S(RX(Vf_SCN]J.RK4<P7W>PS0KCaf@M1V:1Hd0<)@9K.eDV71aIbD2Z#W4
;P2+8.,EW9Z_WLLD72LHf-L65Vd[6UOeM[?06.5](9WHQEE:3Me;5HX97d\@[=_e
W;c=[gR:MGHBf+4]+L8f_=L)B=F6WgP6IIM8JIJYK787ccf_M.[\#(N]1>NEJ8/+
]IK6-;ZYZJ7ADZ:b>13BCD>VO-2_b<aLb>[&(>3[7ZQSY>Sd9I(<LO)Zd\LVP3..
W=T-<^3_GN2H<H^^BBWI^c,fA[A4NOS148g\HNB9aX0UN=/XTCd1S_4@+d#g)YQ0
4D[2Be&R[#A[9S<7F+@9S9T86C[\LJfbeR0/+eQ@&F&61W+SRg/9I67T0@8(#^_4
#C_3+P6T]2.WV-/[R0(D00c_A#F.S&])H6X9GD<3#0WE52O?VP]5TB(Fcf]5HaUN
UPIdW+4.;]FVIS[G:R47EM0dNL&.,FODLLBF>fYG)KA^&@IL14;WRXYKa7[AK#R6
WU;,bS&,:L8#fd,)W3Md[X[FWQa[?aZLW(G6CVI?2^3Z/AYX<Vd)/<7?g?.f.Y.@
O.MB.R^6SG:1ZQ?_>S1[SN#=7([+G6G>^D_F[?CbgV<<\8#7YLR3fNI?]R[&H]CC
,N9.CLRL&I:A33TWC8/Zb=)_8Wf/=Gd,](2B>gNL[BN1fYCKR793ES7N2K<,:PE2
<\W-F]V,N]>+gdI:?H^@[Jc/B4H[Z):6F:C6[a]&We5>@LUQUfT)XL&L77Y]DV1d
9,:K8THbGZVU3G\E<>OEdGaa5?<SVTW83?X#+Q]IBd3RC4<?E0W>X.QNEc5JOD:5
8C+5)>ZNH.7XH0TH<?)-1fcfUD,aZ[E#/1:A21]a7QO[<EFf7VKE:BJ>g_=WA#\(
AIVG9d7/CEa@L>4#.^bG7F_FGH\M?>?K>^84.a)\=H_#a/#-&9<[;a(eB1Sgg)8G
36?,:5R6XLO?M:FNb,F5eOa<R\c.)_3#86DUQeIMY=6^8B3RgSeA//((;a^)XB6g
2((X0cI,Sg\_TKX5/74KO#DEU?P#/9gQ9RYRTRQBf-_PH-3_PRg5F)9:Aab&EV-&
58)BP>1R9#LSWAb3+#CA9.-CUE9#cF8YE(g#[7,Y9)&f-7-EOIa/I_FX]&PDf,K>
5(B?>_MY\a7<7;GH_MMH^c#Y95U2f_&YM0MAf/JA14C&Ba;-P2?U:S)-#7E3,7NP
]Z8<KO\YRXT:e,)ASZGHJU_21g\O)GaT16^BHA5c>@4[a)bCH0CQ&=K?e^c=4IV3
9]?O:NIPZI3DY:_4D@2b?EMD/a=c:YSZId:78T00c@IG(Y2SXVGFW(]3Jc=9RN\&
W)(db0bWNS-\K^>J@X;>EBX#.O6=A:Y3]H0G7PYHT6>:3GW-U0C0ca5?g8G.ddRZ
@c>#CM/^,bQMFBYCJ8f#WQ8(&,7cfe8R^g:f:#5-)1V>\5V3@?1RFKOZR,GY;8@>
Ca_Y\J_PeW>[Ze(NKIMUC_&8:#,\2_/?f;(HOA+#?<E(8f1C3?#b9,RTELB9_0A9
@37L/J?b7N/93^Oc\O3D#Ka=99+PQQ^MVL7:Qg+ff:]6#@f#ZQI.3]g/ZFQ&V(D2
TM1G)5SE,R))\U[,Cbg>>?/_.F1@UF&VC]J77Y3g?)NeX,/PEYgZdN?#1P:]\Db6
c\J.[P3O>VNR\bVb=;1&9S_:^FAX>;5?bOOL59:0XGOW1,9c-[1cRQ<.?4F9H&fG
C2VE/cb:d/2Y4T>D?ReC5;9Xd6L-aBF>DbgbV/X>+&NXe-9PSd;7P/LdCP#O4N>A
EJY@Z]5UG[:&<MT\NY^63cH(_D+O#fV>^0\_SJ]fS=->Y4H\Ta+dC1#E(L^3SMcM
JVAO,agVBEIK3C4)1<:]d+O_=b>^9=?Z8E??L&X:/dE?KKMQE:QC2[A5[75B:_b:
;&4EW;D_)I16QG#:;AgQV&HBM(S1)Q\CT??L#Dcc,beMb2J1]6HDIFZa0^37&C7C
cCOM7HUV)O9U4#5:BWR(\MXW]YZXI<c2XDY0E5O1J@;??b[Sd=QT_YY0FV[AQ70?
&01,.9+4.W]^?QH?#RYHQ@S8U,_0VXHZ-fN=(3()aYOgB:Hc\N-(I)(b>HU\(B1b
ZdG)Sg-.DBB.W7)=bFRWXU)NGR8M4aH@Fcd#HM<bK]KXMbU83@R+C8S,OH9Nce8I
dI5&T?QV&cE>@01QB;M(KZb56IO95TXdWY)AfOGDL[/KE;VPDP\YD+S]Q3FJPKBZ
W?/+5C8<QP#c0+9[2;2#A8d4SN_K_=X,[[?.aaR&KQN,Q+S97MIE@E;@gQ6Q4EBJ
1da^),JA5]FXP]f3:6#e)_-_^8Y#E2=6fU756Wa/23AcGOgB\2+?=8B,R/5+P4,B
8@;CcDU\[+_T.P77TLc??8_E/Gd_][b,,aR2,C:GM\Ug#JZQC;e0UWQAURU=LOZ3
UaVTKJF9D.L,TN=C?UCGV#DI)<>@]+G5(cg#RIT;/-;Y][@WgPD/9Y_Z0^E.V7.a
=Jb2AZ(?K8-@E/W^(339Y##845FHT-8YP;VB>ZVHTg<M@+f<&5A9#R@D_4)JN:2X
FRAQ4F]A>18O1dTBZGO8V[CaNAZH8aZW:>D::1;\[C#+f?M#N23Z7/][H4<(U+ZW
[WQJ:+II2WfHX:WEb4C-WJ4>6][J+UYRcfW)G/CAI<ZKb&_;^g,#(EH6#0aM?4+2
#9,1d>YBWV-4Y0<^fQ)G^BGVbAI1+0H77GK).Z]E?1)aYUXJ.5P=Ca#)Q(S=-3UB
MFD5_.T>[/(a\^DGGXRZD(f-OAeCbRbWFg,D[<W))d1(FIB#b;;XUQ3^]6&6>@g<
:C6(^ZTI#V4,c9a_/JS<@eM.aN:+Q,DA1JdH7W>KY7N\bTT+\agVNa<NO+V2.cFA
C.BK\FQ1M(S\A</#YAg#P\A7751-^FNMF1g<M818+;4ZKS,M83PN;?f0#R3PBVU?
)7GB]7#_G[dOCT<1UU4>IZE/W>II?6200#dd;R\.D=a#F,9/HNd04B.-?F[B-=/X
^KT(;Y/STKL4Q2VMEQ#IE6I#@?L,\<VE(Z2,e5IK9/@DS7-;OE_YRd]2^2X:4<a+
M;PZJTF@>g[f_bY-<e2/[JEggfabGaGFJdF()K)HH.4OJc7NZ;1.g69,dfP=#R-U
PJ^F9,aY_W<XO8/N>#=_\PUdQUBRAZ-fK>H@B+GP]3J+A;BM@R=Y91UcK5f4KK3.
0=V3RGYSeHEAb.9)8<\O1<SN?_Y94S9/959g_AWO8T>(U7<A;>A#K9(aL2;+BTcR
/]9;2^eA2P=XFFcd7U,.=IR(c,QQ2?F+<2#.Cd#gA86(H7[K?6_4SE]eF8JJ;72c
8-5#_QU#aE-Z;6VL;))@X<Ad?M,5<&LRG-:aB.29[@UG<-MPY8BA=G@NcAI4?c6G
C4IKCFM6I&EC9]fZ3@HcdV;472FE9Hc4S]<gb0#Y1]cN\MJ,:K_RIb=4X]#EX8aA
2F4_+0>T4La.O=D_;bg;>@G?XM/3V)=H@LIX6RW,[:O--1)bH6Ca(Xa.0d>^g7Ba
GMef7O1d]WIc)4NRF<\b-=783S@HH(WQS#EZE\aR;0_-0Mf.U47/L9:H?T4?6J28
8_R8EY]PS/S:(PLMe#e\&2W.?C3,g5d8(VYCII,e)M.a4?C6F=I]Sd16>P7bJ<2;
>D3#Y+.MI\Waab,.)W;<KNcY,Hb--],eI-<e_I]A3g>aU(&\;XWRG5WS0ZDafTNd
@0)GJ)25S;U+5/O.->R8;8Lb?\DQ+W;7@d^WP-9T(.DZ6Q,=G9,[[U(0A7T<VbY1
0NH9ME#4V.@@_DU,0IL(53../f3O8AP<ZC;8CX5IPWY>9G9DA[1HJV6P^@=Ke?J/
0TWS]1Tg,VW?130X+#PT4M@ZP/4C.B>8W9=&76T+:X+Z_]fN^NG7dIZT+=1&[)B1
a)L&/MFA<2UD=Q+I]6S-4[c8H2OKMD)28Uf]NVICS<H09BHWGU_7ZF_W+\7;5UL1
DHJF\[>W-0IYEdZ:_+9#&,QP6-#\gT8VR01_I0-c.MZ(77ZdgIYOV[a:gJ>GR:YB
,SX(O,08D+Q_NOd=41,=_d@Jb@C=YPK@I#:d)JNIRGEK25M6agSc^e/d<c>[PODW
gRS+LZT>\O1a6F4ARWL-1K2@aF_MWOMW=.-aWf.&7dS?ROf,.>?M\K=;+EAeKcTc
XR9L5/?&B9[39/-&YQM@cB+G=bQ&\?EJU[Zg7A6#5[e?9OJfQ3Q_9RZ./P0PNE3&
2+6cWNgBBZ#3DCSPIY(@J-BSdE0Dgb59-d#R(ZaP(W\@DW/6AQ.S>NI/C)E/gc2V
VT.&GOWdM-^?A<1:JW6RE8bgO\UVNe3<N639&BaBM0?47.U(cQAW;-1]A;/&.UO[
+I27+;6d72K6.X9X#;<)4a.]2;R=,Q[(JeV_9^[[#dQVc@?NL.@7?(#Z+_96^FB.
b#OfK\.KGWSVScN\1#^T;BRbD8?bN>gdAS,S/R\YdDdUVO@==RRI/1)F]GX+:.SW
I.UA]GZTE/H)86Q6JVP:bWZQU5\JR#62Z]]6.M0Kb30fVdPVf3^=b2W=Y;.b?Zb&
,/35R>^a0Q]Va?Y1_R=Z37>WC>>JISV)^^12#<1[)EJJ(Jd3Ebbc3OR<#/S3T7,4
26)?Pg?FO&L]BDF@E7HU\R2+,,GW,SR81J?GNf<AS4f\<M9)#Lg<O^(2U,SKSZ(I
BY<d5D&QK#)X>5CHOO>K2L:]/3ELY:ZQXK25\?3gP(,]O:cgO4bL#PY\OeQaCW(>
,_P0Z1<[b+9NSY+(5<41S[9]B8&Lg=a:\VIbU)1U1X-^6PNYd=ARRMQYC=BM[e(L
(Z:d9Wg-91)]d\72\:L#<Sc+)TMRcdg-/>3[-O@#eW-NZ451]R,Oe97.#Y;KO=KU
:]5DK1V#/O1c:\_]g3U1/,[RU(<g:?g-RCZN(V&7f8f:f-UA_STHCCT/Dcda;(C]
6,WP:RdDPeWR+CJAaX7/E&@LaPT45c2E2WbOE@)_N?AbC?Xbag.,^IKPAfeK\F)+
g+L24N/,J)W>\CI[Z4Ibb+(aTaQK[J&@\\d9U7@EE6JZ@d(7FXYA,OI?XGIYK_aY
MIV)L+@Y#5DKGE1b@)f5c/8N,_+\3FGQDHf3V:Z1KQ3f7?Ie]/YaM3a<A2Mc[-/f
21G-,)G7=V4+ZJ(KGJ(>e?C42_?YJCNZ24f1feW1)MXQHQ#./0N37\<[g<4K5JP@
39I(KMWM(CJ4O[A_I1ggQ-G5V[)LJ:=4F1[ZP]NM6=0gd85,Q8)G#9>2Z\,@(6BC
D]FFYcF36Y;:_(=CEAb9]ISVGb6d4P8#WQXN,gJA,ZPOdf@8?[Z7T0[])-Y_d:/(
gB@W2FGS+A10;e\5S8BK5P/^6e@OgKK8HD]G7JMU5JMDT&K\/OS@B:0,JR(5ab)K
=0=UXO+g+3IAVD2)LDfcA?E6R5LgI949&#SaM\.g[(JMP7XQa2U_0U\dH[<DgA(c
KJBfNG+3FS#OYA=@#agD[(cVCG@\Q?;DY#XNQD_20CcEU)dWCD5Sd(#Ba\9J7]7f
[EU7S#BJ3BBCHMW7>Aef:aXg/Z6T3/N0N-[)C1H#]\g[AB\^/Z27S4T@_c3dFQJH
fJKW2O,5AUS&dP_gK4ULOUYf6WOEV1d1M/N0^H=3Y9-8(X<2=;HFTDZFgL&f1@\]
W(34)fQaI<#W&a)a<SaIYED-NK-2VGU^#db_1)-NEUYKYJXLPW_,dM48JYP5^(S-
I^7g3:8RL<_Ob9SZDdf@VeO>QP>I&6+))7E^cMTaR;NGO>H>1.WCScZ9bFMOYdc=
3fa+,?COM[f0=MW^S_b)R(ND@TB)G=\3@1XP8H=ME_5Y@Qa&_79NUA@GFI6(QJEe
QWe>3\ZLJ1Oag244/RLd6ORg+fOIS:HKef#J+(5d9:JN;<.eSg7a&9TC2Q>_WW<O
)M>D.I=R3Tf2DH./Uc9Xbg2<e8LL1+-QL8Z2G9Wg>\[cb.bcJLLPR\c711N?A^?g
)6Qfb>BB.\B]&&&_P2EIP^a1(gO7dDQ?6Q6TKJc,.C\3GB8D3AaS&V>E)Gc-P+,.
P[f664IWC^#b,72J?1?cYN::EM)C3OH6d;M-?V,ML@/D:I+V+[PT-BZ]+^bV7G<M
cQ?^Q,EONDgBA(M>&aN#QE+I3P#7A?TV68EDSHbSWTbCWeQPBc@L<),)B+I;;E1]
\4e#-+fOcaRR<gX/.J+.ZWC-K3QMZ+RI\<&P,_H:UL4KOZ/^STL9Sb=+XOZ2V;?f
cba.#QGY6,Y(>SR18S:MERZI#&.:Z5]N=P1KRU3^_([a=efI=dR[<,GE+@b]>8)?
J)TR;CO^GF>W9b1X8dMaB2cc,2b\K(-/S5dC@BVEK-S1@JLGfZVeN5^>?X20=)fa
V>Yd#92Q2\&&9cXS0VJF[c#/.]Y_Y=NGf^=G/BP)UC?&0-VUS2GDJUc&@TgN,dP?
688OG&,We5@eBcPC8\90,EH-c=/[&NUE-7IP@=YJ>Jb<74)&)CGT=S8.b=N<@R^]
Pe&KCKNdBd:L\393#T1]a>5/=2UE7_ge9b^>/b))Z84)]KEF97NB.VAVM^-5+GQ@
e5fZd<DC)MZ&_&2[-T8.V29LQ]6f-;=RcJ(d:He:TfMA-R>#)HF9NP<#0#RP=@0<
I/MBRTPSN#:E::\e^,\XQH\2):3:41PL[EJ:3C=71-]\R7bd[M^>GGTF-0=(W)PH
>30MX^A-:J95?&SFH6BA[6aZ-\XWUH88.-P?OM3f1T496KVce7JC^BF8LW?Jd4O+
:)291?T7,O_=[&LG<YSaU;8?N&&GN/1;3Q1U?Z&dJW=_&B@_.[3+++#LS)74TP\g
]Jg7HO0C(@Z53F5g-;JB>)PI\ee15KLG&Q,BH#1=/6]1]_3[F/08F8(L-8CgZAI6
6>LHKQ7a)b-,9ID5)-]#e2\RH?,TBI1K;K:/;@\(J2&gQ2NSFaLU&bI6VF,VKWCF
+^MM<[e)^NFD&=G/D?(d)GB]#0d_OQ4;Zgg>.cT3V[\5D).BgZLOCCg?T6>NQKDR
QT7(.ZN<@:<,d&U8D^+E0_+dX[9?U48gU^IDJ_d_UVMaSM\?F]V^g5<RD-W6dP:C
W);J,TV6D:JFS-DbQ9(D9FKKC(2O5Ka^\bfM:QAS9Vfd37/J^E@fa\6+We<3:([S
JH<Lc#7U:ggf\_(2LQ-&\3.&N].f_7ZaR4OT/,,3K+P]?68+f,_#cU1=6=2-,L&.
A>[P4CK9YIX>-/24=0VC_X21GEWA&KgaTL71aFY)=2ZVeD3/PDI#8[ITIE;]R(Y>
;PPQ]]IIB>J.fP@W\4FRMGHcHM/?HL[d.2V\fUJ.N[@6a#9dKQ23EO>11&HAb)9H
HN05L[4:)S^Qc6MfD\BcA0gP6M&fTF24X9S)D7:UXPC>.f5]@V3OKRbM)\QIEZ-X
_F@G^gT4aR4F^;_V#_bT9GL>5B2g)cNH)E2@[=1;:F6/TCfeMZY5IO#bM/FU?3?+
OU+T3-G<HMeaA:BWZd1K4(5-RPf+@,Sg:9CeET;QHU5BaTI?R_bEPZ6Wb>#<#D,8
U9+C9-KWOf_,(][(c1_N_EC7/-gFKPNP2,UXNU3[b(fCZD>0-E>a(>aF)gUT(NX+
I<#a760S\@[X-I7<E0[D1Y6#gH;=DG06Ud^Gf)>#g\DbL+1GWKbFL-.WRe3+gb>#
B;?6-EXT1XBeVd?4>K4;D8I#3+:FIU6Q1eM_geE:_Q0]Tf-VaN_2@IP?A:3bd?69
,ZX(B-BUF8<W\-4OY^#PBM6O6c+USTNL(Bg25^EV.0/APVECf-CTP&NdIZ147:1V
9]1@f>7)3<f&#?(PI=g73;9\9>eLZ2GA1cT5#O(::VCM,Ug=\7)70;&W.:BHM(9_
1C?S4Kd/CBE5fWJAMeA62XA;HE5FYAZaAc[\a(_,Xc6AXb,;a[bL0FVZB3XJf7K4
5W.c;T81C#c#JE;D8e81ZHd(b)V8aH?N-&IO\5),Od();1b[<K8[d:R3Bc)(PM6^
Lc.6+-&g,O.90Z)OY=&=H#KL7d\#4-KH?E9?1^K)e?d#),RfgFX)?UEJ)3@_XF@)
4A;H8Z#LX+=#A3Y\CIRa1L<X#OS1,E8UTeC-DcGI:>A1]bO.).0L6WJQa,>>EBN)
,R^6APW1I+_Ug0L7)HZ.Z89+,5)&2]f&f)94#cNL]EWJB1)QIaeVKeV^W3EA+/:^
8b;#:,Qc:dI:f4]?A>A5V]9&8LfV5JUOX.?X[]02..0-DeBQ3(,\C#2KRNZc2\aA
&&,3\Db+AVaB=V/f^eZB&.MWg^b9c,J^:UDZN&:-FZNAVD=:dB(9Y3+>W+M0W2]N
41)OB97H&N6=;SQHZE)daR>YGJV;Q0^?e,e7PG^C5WcF3ecBQZ4JM0DV.b2ZQ>Q/
Z]NLDf^2PX=UdG(()=2-ccULgRT?SCQFAM\^dfBY,eaQ97I?,_e[<;IXC+#3VW]A
Q3+.25S>NAQN8?d+f7H5RM,aLY?\-B5:].G)J;UU5KW2++K]J;-2]U@c7e\Wf1Sg
#).96#A8^aB6gSdM.H>f09bf@X<@DLNCFWg:N/Ef^b.?_08<&&e;bfU1T,EIb.>Y
[gI3gD[LgSa-PR(:VeD4f&5Zf2Z:5@5g&J&^<-EDK,4T_E>U:,d=P#7Y[IJ/BO&O
E\\V+P_3EdB;@L;Y9eUAd;/?H?#+>WD5U-g=PcGC0XF_dPS8D/[EaGVJKN:Y\VQL
JE/BbMST_?;cWP^cbS&SeeTL9MRg@SBaZ0T?T[?aOgNIQ(#Bfc2eGJR0gg@J0@Vg
>NUG(2d(9[7CLW16_W,?]=X?3IQYA9BXdb)[=-C4fWY3aMI]IaCZJ#YDT=Ac0I:A
O@-DN=f_X):Z3;LZCWJC#8IbM?^2=DU<CTGaGe[bV]-8bS1c-gMg-B\+V5DYd(^6
(aVP2L?K+7#2S>JY_bRaO/FV=5.DgT3H?J7aOHJRJg(0Df<O#E98Mg1EV)HTD^-7
I,<K)72O-X#X7D0\a^F^/WPA;>?,U>?\<H1ZQO7DE28H905\cKX@U-00a^)Pc=(S
2D>Q0=Ug?AR:?2Cae1L\A24)@1;Zd=g1)(ZXB-)SgP=]W@@_X(?4A3Gf<-[+O^S1
V&78N8UY]S@6H(cI:HF8:#_8fcJ>?M17:\cS^736@?^F4D8gPKE&OLfYVbTLCGLF
:,[H(DF)^V11O2<F7.a]RA(6I#YP#d&DHM\A;ERNR1?N)_(=PF?,//0;d5+e.G7P
L:+g#&Y.KBgIgJTKZ24,?FB?=X>.8US5NgHaY,<V4KA[gN^MTLH@U:dJE>#f[Z>;
TZJ<_BA>KW#[Acf[>L<FAM&Uc(E(@ITY<&>-]g5-Pd#5)X6a215)UPFKYYe6YB#Z
-/G1f.3L=-.e7&4EUJ=HG\b7HGN_B15.7..OCFZ\_?73F.(P2X/]EY.c917@GVGP
A9&A>;f.U/)D7=Z>feG=<V>c3K[L+<^XJYYUK6Hb.D9(8>aAN3^L5#T#BU77[_eG
#9D?<;F^QEa^_EaRQ=;KY8-ebP28a3(&MEZRQ1aWV,Re6>7gQZG87K4QH6V=)/UO
+Y>-6ZPX?U_cIQ=G0904D:DXQgfC5VXH/E^N=]D4aOF.D.ERD.9+_eNP&6P@C\G3
Z7>L\Z:@cD,d>^&26C.DX@DJ]^SBO=@YDJ[?)ZQfJb(<:#]NB84W^1#;B+69.]B:
8WPg;,.#DDg(Y;:VS&I@EG:5JfF.94J6NgbN7#S6^.2X(fOHJG3,U59EN1c+e?g,
3,XHH=9VAeYc6#.QH:Y4@ZeN9,9=8^;.-AGJOHNHTQ/aaa<e^_NdF6FC8fHP(89S
1a3gD;/;)<(LX^5CZ,LceLP/A&GecBE/&cH1be^\8X<;OD\J5[_DY7d(ST#S+/H:
<XG2TD:^D-9^^F@g[VZ6gNT.WL1e/^5dR?Og>4[UTQ3:;^ND&;#Z0ONe8b;/:ScL
OZ^-U@:#4b++aG4Z&>ESEd\<)V(gUDfcR15<VITf++?H^YReS=B;Y_-Y:/>ZG/Qd
Wf1#^L^YfJEIEL<5JRTQAXB,1)-STJTN[8EObX0Ke3?->/U#a-0#&G=Q8CJA]8OH
230R6X4J24)b\JT&ND0LVO[M>+?HeK&M=:&W&IM8EeK[C>N(H7:Z\_?;5&O5;GUY
B<:OLSJDfZ9a@.;Db<#=/<5YfPOK\2]\-bXa?E:N:ICB\TKJ525RA,3L15e_.<fc
6_#3K0XO_W4\]K4Yc@=IRL.^AWcT73]]Z;b<+BMSF_/E1R4^fCCQd9d-E^SKNd?(
_;8<ZA0GI(C+:9#>AZK@?XC(4@VX\@aH,?G:L\VP?:<52&#I=_[bCNMM91NE;\7[
+,?Hg[Q.R(R4/AgHQ-;QeZ?B.#W.4SFL@a2058XZCS3X#_;T0;RO+^E&LYg1dC_?
Nd;N15SK@Z]H9F(,g;\2\HP68KA-R@76_RC8]:Y1SOY/_:+IV(<W=&+V#-KO6aQ[
KL^FXVLdM6(T:6/C?gIJRLA30(:L-PL.\>X.775^G7YeP;V/R3?G6&-5b\]KFdaB
>C\CLK2ME^)1&V-KQ?5+M@_4^=S>HD/XKFE-,YS\RbUC42Kg[V&R\QU^LHc3ZAFZ
^Ya0#;DI?N[#CH4.RD(;b;-DJ0#WBJ\TNW.)-cDGCW_4IWX==1[6XSW3[B(M:?KK
_L?cFb3.2NJ=^J:QKIJ>GeJ7ebBMbJ26<=LQ/@)Z79X7,VNc^:eWN2AU\X2TfDXA
cXgRVL.RKD:1+07Q1CB6I5#SQ^5#Fa+#/ed,QI5/>CR#b3T),D-N=6a,)ZRY5CGd
JEW9b&03HM(K\4,g58_BVFX>f(.E0REJ44>aF@\T<f=5LLJ-LGV93a-=V9U#bHMC
HXCX2-<>[YJX=25OM[TGLO^=P0&??1PEMI8I^(G5#.CP;_F&#Mc1NPLdJK<LQ71e
,#(X(DCE@e9K+B9L=c?E&F5:5c3HZF>Z#/KBDV&Id8V;KRFS1MWg#TVW/-+E?_E;
=(3gUgVZd-d\R6^W&U&=4QDd9BPEP3Qeg?ae5_=0^A&dG8LSB5/OKed3\+_UI]J_
(TC,DK)ZE0f5]ZO-AQJJ));:HgRUU-d:DC2+10#^P8W69LS2g20QB/2<&NNQ-KQ>
/MC@?UH[(M/#P4:+:X7Q.de2S1(]c9KXAWJ:<+>:V-L@@DKOGQ89)4BJb-82=)YP
8B0+:^=_=<dVR[8^f[fIe@N>baG6#^_:2HdD7:WXO^=R\Z25W=_=MFOE21?c)I-=
<R/0gEd#4]\&Y6T2F>DdOI;7#8J0cC&TXX8YXe7e?H>aKb+?HX+5)LaKMAM37d-a
dVVO&8UR8KAPMU1/;aD6fT=9+SKR3)f(.[J&:S)A3-^I7;Pf,VbIS0QM3-[\[@1H
bE[cgIbDKXH2;=>#7&F.R>9?;]]DJK<G8D?1X=cZ+KgG-NN4&c^M4G[^@(RN)UW@
cW8F]P@&5(J_d<RUd5ZZ\IGg>?C6=D;^AQ,c[&R_6GT,]cI=>\HUMfR9]BWGONLC
H_+78YZ@H#VeL9+[e3^abCLTeCfWP7d4_dD]K<J[APH\d++>37+>C((@b.#faFLV
TAPO9Z6]#>F:GDWVMM6Qe;VHZ(2Qf.,EC+[)461cE]+7O.E#[R,S9;3=(;J^aY[\
11V[CMf9+bA<-D6PTN[#4B&fY;HZS^IXZG^-g@gfMXXO4UD#WY#PPZ\gP9(WGY?-
ZC/c9YHWUeDE/VOOY/2cNF3/AFS^7KUCXMTd1/582SDbX^\^@@0W4&3\..2GWPRT
^=#K\TO\Bf1DRXS82M2O.eU]C8IHL(2<SV=.I40YWF5#X#g5IM=F]^GM,NbMH2;:
\(ce?M43=VeCO<E75MRc/]bd]+5;ebHJ7R4\P2J2W?W11^g5V[cI4[6:3RWYQ]@V
?a):#AC41.<[#4\4&SO[N<Yec.OfGNGQF;:IWH+BF8aC(6Ng][MVad/=/R?GY+W&
LS(<gJUD-9Q6.#[A_g#G(Q0c=a)[UWeN/@_aQ9_G(B)eZVJKSAQD@T5>:?gU(UY2
SG0c6(O<#AS=U57ASXF0T]ZN_/:MD#K8O./2b7PSeRXQ/I0&M:.;bXIX->fS\FEN
QO+XW0G,PHg_?2>[f+ddB&0(<HN/_SRHQe.:EIL,@4Lc.[OSLf#E5H2gd9?E(D@B
.G8#SK:X0_DPHLARcZaBLM3gKG>EaSSCbL6S7]IWWJAgS,;)G^EY>(?abYC\FS+_
@T8;6Z&g2\8IVGJ,H&GYeQR-DIF>IU3PM;7=0MA#d#/2<#+SfUA6UK/OPLU-b1gG
T9P=-_C]Tf\ZI.5[E13&8M;>0\[#>+2>ZHZIPNRf_4ET,#61;AEFHcNO>Pg9+GV>
0)_8@\R8@X.)#=VKZ^5N9)#AV^19@g]HCdE/5C,2]Ue;B9;&IUb7+a#(,DF3VK6F
Z=NGSMT,Fb-ZW8GG]N.Z#ZZ-)=32>fAN(H&M9#9E&be=;V>CTX5YA=:Yg6\@0?==
U=a2]BBVD.;0(1Pb;O<eARTWR^_UAXc6QTU_7X\?c(E@.LYb?EVcGdbOGZ;B[9#e
W>9dZ3C.fK63-@eX.aU&X2G@U:;UMF(DbY.1AUfZNXa#JG_Yg5;Q.2KZ[<]UWWb;
WKQ@,]R,S[]f,IaV@aHE,/d:fUN=,GcGF.fX&MV=[2/^cDJOY;YTV\\G-J)8/9\=
SYc1.F+?Y)Q,3R8<_KL8YT[W;.U8(P_6:.^,CA&ECZ-9)P.FQJ:+.)d3-cc)Na7B
JW9+T495[I)Z.T7,[g]WQJMWLNX9ML6Ngc[#JI0cdW:[YRHH]-7:D-,.fXYK(5g8
TX?S8_Y2DVee9X.A6,,XL.RQe:H==6^gY<3/4a<URI=7AULZS]a?12__cE(S=O[S
(X[@bM-M<+5(Q[A7=+a=?.OX/DQc3-c(4WZaXD>YN45@3fF?Q,>3<R2BZWJ;M)-:
NcJ0aBY8G27fea3WQWE15.-Og)g<.(/TO0Q@HJII&OCb=9KN+JK/NZO2>C3,a-&d
SZ)[8M(H]R)P4g\T)HJ^.Tc8XN3W;V(AOC975-NQMfB6N^AA,Z8Ae>JEO46>b,VH
?Y@.<?6E6:aEb/2\:ANGHA[\<(.LI98_>cRFbKYVORR\f2EeM0^1ZQM#=cb;S_/Q
/BJ3@Z(\@AWJSXDbQEC>f?KE2?_5eW.QRgWeR5e8HBK,MNgG95;4gZ_8>S@9AbOP
\6AYN4PCGG8()3_?C0:0MJ?+Tf^5G680NO9;+JGBB/7J7Wf]1P?44VSP.VE-KJKP
HPANP\_)U<<c[0J@PFI:;L_]aK,ROHD:VCf4:>:9>6&EQZ8@a#//?]UM]aM7eK^5
6\FVYf#B@7KQ9T=IH8C,VN;>,J76)F,aaJ59>RM/J[6+T9R[O;>9&ROB:2Z1A-_W
25I/;RaKSRE)@fRJN/.b:O7^>,,:&a4e#G^XXV@L5,J4M.Ae#;HCGf8:1]^L5O:6
VZQX)H24];0GXT_+[O]d@(#)Q/2,Q0<;B^<Pdce9?PN#KH<<9Ec3)WA7:,<aAQ:e
@8SeKYeF.X&4U)QJ#KA^ZP.Y&cBa>P-.?A_6.dg(&9V5WL0;+g:F9-0aQ3&-=QfH
<#N&MZ;G=J.c,OH7.-6N?+da;eAZ:1720UTf:,J_=a=@MR]\0U?d0.U3<LR)7TfR
C0-@e)KfAc?/Sa_X>#abFXbXfAZ\VCKHF.6@6RD&ZY?9=9E@gHLB-/G(+:BNCH?]
?&]X<?9GUXMQ.1-0RK=Ub6\F:f937S9@KLMKPW.JU9/.--K#@gaCBU6AW&Ic]BW0
e6a[F1O.Q#^KUD)C5,Q&KfID1+^H;>4a6\S1_KLVI1V7JMUH0eAXRS0)>A<I^294
9H1)WgMcE^QDQd?;HHC4IX263Y[c)DeJ)U(@9daD,70:c.UMbY<MEAQ(NZ=>R,X_
fL):c8R:DFC>ff4R]54<JF,R0YgEF-QfG3bd=VGNYM,c[1OM:3Id)V2GCQYVKVQb
I/deH^2^3KFDeGG;]A):L_L.7d)RS6GY5K9a=WbP2JDg1_,IAK1Q5)TWG1LaU&NO
C=U3W.AB#aC^S6TcX+,^c;S/B2-<T)2A#^SRR\K\@TG/AI53^#IObeOEE8?.A]&J
>-Z_VUEN#0Q,/?VTbDEP+A20QM^?)cU>FFP]0B#Dc,XOd8,MM]+J^aCCBJV&CIVH
.@R@8W:eZ#NR>cf.PAegUUKbL0;(9B2P.fMS;HR7F,2a>9.&W^FI7_#QD#[?5bb6
bg?Fd?Pa60X)8[W-J+<g>VgK5N?]@(c<U55?0^PFVP2_Z<ZS@c:U[H[HPR8//7aa
a3N6_@:@@S9KJQc.LB\&ZT]e[@aKH_ZL=;SM,]aFdHY-3]LAAgZ6KR:_?JdbRaV[
>@?KF@g>A>4;B,LeWHO]b>BFZCD9\LQ?CJC5c??7=\bERN4H6NO:3F6#K,)F>;X-
GB_5PK0^UBFObI+]\E(dYD:^e7C-05K15f_=8T(R4WSU;@/)d;>^0?86<]?_&&[6
Q]#4HI..<aNC#SaBI>EdU)7eLS6TL[0&>6Q-4S^MfJGC+=Ae^W7G86.Kf9.e?N^_
<b(R<^E<ga+d:>35L0C?CJ5ZH50^8_[7O1FJYc<eV6CE_3F\E8XH0c,HTFR@^:7T
BV?MBMLH-F0?7,)6,U.R-OP6BX:?c[QRg>D#WNJ,S0JX0H+XNfO00C1e1\+/9^QK
ZS^(:gG@MU00/[#YPF5/;(V84>D2)D1,/F-/EBT[()=,9&+KdG:QQ\?e3LM+27G:
[I7>+4/<&F/FaZ]IN#[Y+#RUY)S&Q/f[:?dGR)&77g9dWRBK7=5?dU_IU9-+Fecc
[8e)e&BW4[Oc/<SM_YP-d+YO?MNU:7&;:ZW@0U0+-9F28#P2d3Iab=JS4)=C#0O0
P@YB-@[)+1.,Z2,L9:-8/M8EU//#b\P^SgA9@g7;EN4@fS:=Q0Bga5NCW@SMgP-:
.5gQU)^A.1=&[gB<RN+1=]Faf&RO(dIXLL[E_Y72EH+@H-EFg-]WSUaSNfV?;BJd
Y3-R-OcX]L9\[_=G[(4Gb1KaB,)Vf0?d>:fa(4FXOa:/9V0VLAI_:UUPVK7U#,0<
\HY1R[=G;e)=-QSG^&#SaUdM3\[_4(=_:<Y_6c^\.9LJDaVCK6<D6T@bT(F75Y3[
f0aN?1Q)<:[cbB(FV,(-Oc1I5GE@d@B-c_0gF6U=371baD29JNV,>LRRK;N32MeC
NU2.?.-H,f=H>GELP<?8FD7TB20e#HUK9DdU_RM5X51AgP)(L6O0-NKC);e9<JX8
_=d/849Sg9?KU0e2b-J?c-b7\-K^b/Y)[ALcJ;F1P@J=)DN.L4/W9]T4SS@X2QZd
1BPBGd)6[@#4W>U5J-XRH[WbdUa9JGI.=COdY@f\28d:defeWO6CU4Ne)^7HV70K
JN;K)=O=N.9V+4R+G2@5)+--W)W?->:I_1HcJE\&PgQYCNVg^RR5>cIYQ2VUCL5[
;]_C:]c1.6dc.KJ,<UOU9^M]TdA,HBY#)Yfe^9Qd<5[@-3bKKI<ZO38&L@##-ReI
bHGeYZRL;-\,/_ca.M2;0ND[JJZ<,_R)YPOW>=9ReW+2)21QZPN2@V^S9L2I?>,\
f+NY=+YY/]K),1f1FXB1B4dT_fa3M2U9UL(0+U^/=_[P5aEL;c#f_KYZeGQ1#HGG
eAGTSa\3C/]9V&Fc6f,WK]+8\[@YT._QWcUd90_:F<([bZ[[MMW+0^Jg@:](8\6A
+bPHWG];3^Y#;WMLZQQAV4AS;:M-c=BJKQ2cX4N61[&UV2O3&;7][I@6:C6bM:/V
VbP3_?S,^W^d0ZR2^N-QNG+#g7G;9Jg>8ga+gB@SYeR1DR0M1<[=X>0aU8VQ#cYG
/:;.^f5?/Aec,TTg4f)-VcUD\#D8Y9VC9<f(]I&#\B[GBN\)NJR4/AAF4&)eeQRD
Be8V]K;+R8.ebL?U@(JOL;,L^/W\egK-]7X-.\AP-faM38f7P+bAI>fH(gQ//g54
a?L@XReZPF7>@SF?cRT^;-TYLTQbMMf/cMb9VCVVV7YHg]ZK6XO<QeC8LGB<-SU.
:O902caCgfU1>JL>RNGG>?b.dggUZbUCX92CPGRY(]Q0ORdMPYQWE98a-<[MM84.
cKFPE?ELGUVNMdIQ)7.&^?])E3a2-+#a/Z;^W?2BccA=OX^L9F-_S>?_QX9G)4-\
dH+_32RUDV5bdW4Ob-=5X8EQMd+,a<I\.P)5D8LJ,K6,R)?^8^<[DFU4/-4c]X1=
>d(&aMO_-H2];DF5#7)5M:F8&\[;N#(3-LJE@Z_AEWJ/JP:C2+49PE6#d7QM78XB
4,b2b=AUPC2ZP9DMV<&dOS^,(?=0S;57\>8V?)^^S-K?bMVD3E4?X;YDGc\b-UPW
;/Xb)R&Ba/Q=f3@dM?a1,#1#6L)EDP3NSP1STU]G.ggM+7BFYfb9&<MK2-0QeS;^
/@XM/LXF+S5V6?^,4.,^L+:#6G\[c(&W<7<GA73/3=6(g/^5OV[&M/(Q&D;)\=>(
UNVdcF(K0;87B;aRc]8/fR3EB/+J\V.\4]H,=E/MK#4PgS[7UIZEgT_.:fV.0S.M
9].C7W9;9N<QSMb=Z^\?_8W\H6TcP8IN[,@)2T0N:a/;Z&+aA+[-6VU7UG(M9=bB
8G9N,>17YT<E[H7K0O@N.dV;c\_=7@]bMQF9Fe#/I2,_XKb9b]:ZD<>PO?S7(WSF
S_Y_JH-/J]-KU&MN1-dDecHQbQf.c5@>KbNB-M5CJb\]R(TL<,RJN0,&RBJ(MVc#
26<68V7T+BKa-2;/4,Z]f)F[1Ue7,6+17(aa5e]cH?Ve5(DeU?L4C.YId8JNc6]b
TYVVYT</J=_4UGR:^FN=(<TYbYUE@Y[c^;aR@aO,WQ[;-PdK;-OFDJ&672O=7(J9
+0Z]/dA8[cDESNI]F5dHU_AIKg&NEG=L&THMU&#(4G_-]P\WF)I])MFYMC-T)6Tg
,M6Yc5-XIa0c&2/^W&_@eI?EJV;?(R\c0.A;fW\@7MJTM0dIKN<(TT&_<9Q8@1Y[
M[5QbgX[AXbb,5P69[W^LA/9XF;IcT8/;]=OZa3Bc)d0e]]IL2/KVA>J.b.(cSAO
M6WE4?ML?B9-CfGJNZ797B_2B.S&[\6T.5e-5M(T\Z,E,_1R,,^&)Pc7a2Y[_1\I
ZT[Q?c:5XTLPCc_0AJ:0AgX6Yc0,.F.3GAa-M<:7+MK?H<@_4=APEb6VB.RY?S;)
6WW/0\QQ>b]/SdTBDaIgJP]BB=>1ON6#BPHQ1==TZ3-RKa@\;1Cf[S@7b.UD6T0.
dMfITZ82[FH]AAWQZB2Mb-&MZfcD&dEP#WYZT[@O/MfJM6TgD/c)X_NA[F6X-)GW
PNBMb?H,aW0=9W[B[NA40P(:XW)@aXOKbP.?]Ue\6@KWW?TKVO_J15VYFL::9<cV
#N)0\GL-ZCT?H/A0U=4>C8C#.K^]1<#Y\Y>E^TLL_VUFLAa4UNO8:83gSGL1^B<J
eMdCB?_PC[]eIU4207NTBWe]M6BZOLWf2;X8UHDT[A/gM)#d1Q>;G#WeG7>&]K/6
C&BF&M.LWU=CLf80eAfUB\SJ3MC^EN9bQX8?DgG:GZ;R?=/6+\7eCCT();_&J32(
^:6K,E2GGF;OW],b[KNJ:cFKS=^a?FTCT+Gf<):C\81:MbH>]O)EO,]OPeG\KZ\F
O7E_EBc)+,W9gD0@37O?5JNQXS-gVc0HS[7fc?1O;+9^B&dK^J:X[R9)a0XfUE\G
F4CO_(A/8gVR2A@RB]GDV&[^b:K#V.20;4;-Ma[HWI\+FC,L=6DT1N-83c<SaUQ5
f[=gcF2UD;8^)W\B//D;46gGLJKA:eO.ARKWRA^LUH\Q_U9aV\+3d.:3Y\TSCX<b
TOPcD\8#Ne6]&8DSTUK[4WGb0;c\FZOFXS<SMVGR^QC-<a.7&JfLYbN=TeWceR5S
&_M>S&<Oac<L/A3FM.#3(BPR]S,<]DO+V\FX+WT>ES3bZI3[3;V3_B(aYPeRRVZU
?48FWc/,fU1=6FYW4W2>)7Gb9G_=5Q>6Df[6B\_&A];aPfOQB\OB,J<@e)X,AOH?
3+P+P5&5aFaZ2T^-4JfYSD?Q)cgO#?a5=)KHH^O\_]LA@0)85a-4;L-Ac#I?Y0N;
.DHGK(;EO41P-M>03NH(bB8Ca(,T(d1-8_aC+d1#7FT>&@K\NL4LYU#bMU7L167?
D.H\PE50+bO:P\,G:,.BH9^+JOd&C0,LUDP7W1GY@c&C_/U\_TRY47[X_MN/6=(T
>/RJZPE:X8adMSeZ2X<?L]<A5X#WH0R8QE&?9dPP#K76H&,7AH\A?<S+Y(2&=#Ib
SSe(J)bJ4.#C0/c1b=SD))23K0fP\SS#WC-.^;eQ0TQB,WGaBN-<SY^&fBH&B_VI
1;@/=I<XcCB636Rg^aVP#M+&EKI&CIK=-He&g&#0=722c8IeZ-Z6TSaL5Yd@_dNC
3J=2T??0MDgbXE1bR20^YA4H[.b\6QRUQ-1Q4,R/:W3PM;K<U<HP7>^W/=\Z_,6a
g](#g96FXYgWg/)4ENI,K\dMCU&;e6Y7:>)QN3&VW=(0BN6)2GB-d@aAZc?^BGc4
XWKML;TULD]FQL))8+f.46f=1@LW3Oa5<NK-(c2,W+M:?BW5c,bdTDaO0^&a2W=J
B&T)T5KA]3\GOGRb&YgDQD@?DG4@H\b^:6K=;0C&?:cMPa<H=f(ZG3>#GYf]+M9#
9-bUGK)6ZeOL@1:,&Ac^C(SPW4(FA#[5c4AHG11C6&=V9g(L1AS56;?UgQQaN>D4
S:7UR=;(W;BYA4N_#ETG:?.83bKA=5PQM=]D=OY9#-Q#_HYE<DAe0R_+WS/X9H1C
J9&FNLf.)T,Ad;)2DgA\L,>)GJ8OEP_>+-DO&\6MZa[b6?#d]/P+dc+f^6dIRg^(
[ENBFb=eEFN?3;A;_TCEN,E]H:&S?KK>BM9F,[X(4XOE#NBD)YVV/F1W?5@CP127
9:6A.^UHI7EIU6LAKG^KVB&/,f63HcgDY,b76+T#1A6PUZ2@8=RH[2^Ea>\(A81I
_7+(_XcGNLKCV0<>gDgEAR5=dO?6;YJ7f(XeGe>Xf[3B?44#);#X;c1:dGXX_:#T
_)A\R)g<Y#CE59OS#Df>>O]4DW+Ha:A1L6I.aX\1AY\Kg1Dd_8Q&/FD^b6MZ#\0N
L&#C?.9TP9G45;+P#MXZQW;XU_7FK-=#3Hd3_3O^_O/]]GM.O_d9\,E_&)C)HMTI
K0DI:):;&5H&96f))\fG3,)/Kf4dCT]^JV+V688(0>TY8J5C]/ZMFO-#:H,5Y,JM
,6@;MYCgdAe7a5SRSV8+3dD#,2(.?+64.5g_Y/Id)FA)]Fb;fOf#Y@@5C1dXd7I,
>Ic60[;8;_9C<6=E2P0C73R2fYUI[V\S&LKP/3C#d.#]2eDWL.a6LHY5NM:V@8.[
Db<5TLVFDBe#eJB;;7;8J3:U>,BgC?AH2-e^LQ@OPcG8TRG\e941TZdAUR/#@P9V
aR\A3]7LS/XIB:@8U<?Q3-6Q?:^7bRdP)ZcEf29a/Y6ZeEe^SV#4G)/\OSA&bfT.
RT8.;gd;ZZ6LAIT3Pb^_e+CVB)VTSBIWSGd>(&RMN5EZJZcXf</-_5^IMB=(GH_N
6TD/DA_IJ^B)0afJ2]Y^J85:8-;PdK#T=f7dfS@V=f4?K&OHY&6WV=(R#74\Kb[f
+dP/JV#2Q?N)(_P[+?.b&H323?-NBbNGb,)7+4=^_Z@6/2\;#)7ZO1_,a=@fS,@@
:7XNeMA-EIUa&\TN4WKaNRW2U,&+S8]/==_CY=9J^]77cd7g:WK,5QF]RNeAOQ\\
g(L[3>:>X0>cCbaUR;063I0_Z<#UYbU-N5d2@1TUcQdTH5cBG]e#;3Y+3BN2U39>
MKA+08;d>FT?X0\DaLK@)&F;7H+AJ/W:eQI;224/K/-IE&dFeL>T?JcJ&XNbZ2DU
?F_\+d5B>TY#f^aW7)P>.:JLDQMNf[KAECPEHS?A<5YF-3e8+^S26.Z@6CVHAbYE
[-;;0,_MSA.N1Ide@Y_9^9UF#B\f[Y[9/B>G->3[Z:/bf8d99>51EKUPQVEeV5c=
MaJL:LZH?7QeAXgPIW?(]RS@V6aTHTS?RQD=cW2E4XS,\_U]MDLE)BFZ#aKG)PFU
FFD[E@?aC9,?M)b/DH?K=VJ)T))0ZT)^IW[@-UON\_;J=cf=^ZKDa;>=DC]Q[gJG
L8ZdX;g7IRX:L([C80R5T[D_aC1=_#GWHO<.b04F32J#2e3#3A3Y\0Qc)30(#<g0
(dRA6X?I32CF<KP192_=aCT>>YBbfA_-;UB_>#^Y/QS)5.-4\_G4ZD^CSfZ/>a@6
#L^]H1F5@K@2FVJOOc)?9b>B_#cOg(==]?@&e11JWe@W8M[Q2^CIJ?1EX1eY6//4
.]62=c6IWBf57V2IZ_e@J26C[-_:)Ea\#:7T.:D].>X?()0H.QcJ+^83a6KPSEI5
0c?f-VO\HDZRTI6T^F3J3fR3E;W0HN5]NcfV^6?f:P9V4a7E7daUVL;\CZ:Ad5\O
Y#6c,IGP+WFK2Dc+/+-G^F7)\MDA2@U#8KH)X3Lb8V&R+G4-VZO(6\dTA0=JOF7W
IY;(CQ&TO+UK+0(A[R&)g/:33]fbA-7+e=IC@.9gSd0JO^,P=\5[=Z_E3C\BB2cf
8#J>c5AC,;+8DRZB:QaLR/W&F.MBS#gcQ/)_YR6GR503KCB]]T^^_M#4@D8:RdCV
NT(G9GX>3LKgdIXLSg<DH5QL;AQ.AbdD_afL&Y-9;IJP=?Jc+\_d:QPf4=DcG^D>
27KT@@#JU@f&2C(G(ZEXT#NBUN_N2(eMF1]fY_BE-8FVVXG:H.CJFMFLggZ-;Y7Z
4P(V&P?U<(1O@(G=IL7bEMHA-#:bTc4FPMIV42Zg3efW(+1@U^K^?HJ)V18PcGd0
EQ(>(]fJI,;/A5JF()JT531<RQ1H=6X2UQYW[A&>9&;-]^d_EK1fFY0)TFH:;Qb1
T)5-ggGPF@E,Nf#QT<H?c0ea>]MIb9ed)Q/,W0EcHfT9<KJHVU\Pd8>FZ6eL:Q>2
W2Ud\W+VO(Ne(.N/Q\QFXc>7[-+1&1>>XL[H#2C<HHZYB_T8A_?N)8fATR+E+731
.76;=gH2MCAL8WL/8N]OUOF;T8L@WE9]@B<]/LA-7Ha#Y[O2,2[MP+L8^AfR3]g<
dRH68aKD?d6X9&[XY>9ZD#0KY@:X-/2+0TXS\dR4Xd;TddeJEN<VT8P8XVY?Gd+f
CVIZdQ[G2Pb/D-\2af3C,^88NRCY&P-07@X5?Y70Yb3KWJ^/()NJRQAc9?)MW?Ke
7[&G>?e>7@6>d\V#]6.aL2\2TM]F-7g+,K)/)I>?+A6F^N@g)]+Ka#<N0>f@aW>^
2HHSPJOK;4ED)PD3P16dAMF=U:5-(XZ1?QCIUGbFS;&CC8T,BeW+-?VXf/:[YD1e
.2.:Y=b=aEH\\&cKAI0R)_IAB7SO1g&0GK,cX),SF&3GGR#9U:Y+1(X3&bdMbR0M
JY>9)3)9W)e<39)DNLK>@DNXLI(NJ31e+FD:E/d4c?HS:a]WOf6HbFYCA3+Q<^,M
2?gF7\c2B?V3@Q#YU]@O3<G2@KdP,g24S;<G2WZ>.gFTceL<P3eP)E1#Z)5JC:N@
F1.4O&(R\5]FAVL\Vga?f4606Z1KVRMfPA@N1XfJVP45=[=J9Ga/P<2TSbI2W(1>
1V,fa^cDcGI.P9f?)X:\FMD\_eM8DB&XTZM.S\(O:@9QG[ZBP-dc\e3IF&>-HO>5
BDYB?B6Ne6+?C7?^JdaD,8dR/IEXI&^K=@eBa68cS0Q&d1AX[RO40K;^@?+\.FDS
0B<AY>WO8\6-@(-H28?LZ_CU(e-,(9F0XT#(W:(<8[9_S<QY2RVNQN0J\2A96G0=
/WH1Xb177c_]8L1+81XFD6f:PJ58:Q=QSY>]IDf80SCg_M4JQ\.0^&M0SGPe5&)J
KeB8bGg;&V2.CF#_1U<M-AcK)C3UN:HK;PeL<8<]GVU=311JBeFf[+[aIL2;Sb>@
+f&@(YaK:Z;&F)g@7c^BWI#EIOM1@S.ZUcB?440/,+WN_=D_+3E9@P2S7VF[FdID
:b4K-gK6>D)Mg;P5GRKYABFNg#.]S5d6B-^2Ve;0g:0==P)Y-U[R1eY26)4R8f[A
dV?/^:[F4eNM5;a#AEEV92\:a+bTEFfZ/=<(6472]H8Z\cI)+<;VI2?J)3:e4ZKV
\e6I<EUSeGI4;^KOa&3B,V(XZUD0X<I[NG_f=XbRf5_aB=K+:WC-1=fe;f(Rf3(P
cO-5Q]F2L6#9H.c_E;4OG-3[?03CA+X]8UE4_8TKG6-SSdcG,e@70B-R3fNON0C+
O_X_MKeHI\[b-FXSOBKK,UQD?>Y@64]1A#DBS;eJNARXWb/S@Cg6UDQN/1XRKGeO
+_67)E4gKA&#1ZLHe9_9751-8Kb277O+#5A6d7G6#G\.#94Q/=b+LYG0#&E(FHa(
E^Q2D3&b?&D;6T=J)=W3KO#E;=eFUY9>].ZC7D#aKg_)W/85W0g45AZM9IVG;<U@
EY\7Q-0\eZa=EDf)_+EC>=<f=,[@VU^<QcB.A-f?2b-(@\Zc7P/d2_XRY2O:IOA^
#@c5\&6]Y<I-FFXV/Fa/e<23\4B]gbN)&B1DGW^gK1]^X.,GP79/g0M&1]:?I01:
X/\I3/TecfBQ3NFGg<1CT=J=]<D@VE>PT(5WAg^b<L6MbW,3]b6F</0,EL/62TK>
cc&^O2AUCZ)4g?(+_(/S]A>K[=@QO+XMMcD,JD<W9<3K4,M9D-DF\Q0<CTG/+(Y1
PH9\Y/F2d.D-D?DddRWY-C=ZPO@d#FK_[(c39JaMKPA(8>#7BZQI0P33,+MT+W+7
(3]4/AO:QMVA=/F#T0+0:dMd-Q4(Qc7_^X[ZN/.2S\+.GPS##d(-Bd2=4gT>b)8U
S65bfe3?aPV0bJ9OJD?BXO9d#(Hg2<Y&5E.==#E:[4R/DHOT>=:FLb;b<P4<A9_T
4:P[2b3_dDg=1L7LaC=W?,<3)#R94c(MPQK_dD412d&JT^I8N/<YVBQCCM2dM0_M
H[82LH&<._>VFW&+W]1YLG>N[B3+T]IF\:+U-W7Ef#BXQ2dQR4OB+?W@)c]\O]BL
9@,,g(;fEgW<e:dKN;E3ZCPGJQ39<X4IaM@a)YB<;Ka?F/f.TO&B/Vd7da7PTSWH
AcPNPB)-gL;?PZ=MT34#AgT2F=.P3R]XXTM5a=#Y;X/McYf),STd044QBI<I5(-<
AV>0g]7S9YaO.CFJb,HDBgM,O,2BP+B];ZB.ZKWbU)0FI37I[A[_B[2(gNg?54/H
eD.^,D_;RF5+V3URe\d@D/6+XEB4cLJ=IeX?/1RTJX;;.LU+cA<SRD=XC98?NJdV
S/c[W7-.XO].XQV6[a.>C:P=Lb,V4Kc/.-PS&X>67/\@T>B_L2A8-^D@:)MRW8g<
22MR&C0\HJL1]f;G.>6aT\83bNe_8N.-Ka)@&C5S(4G>Aa_869RObRZM<,>bLKda
=0U^RAP8SKL>MBZN(^O+Q:8H,:P^8R5)>LKG]^&MI^UB&dYXF@9+d#;EgC&J<K1]
Q2BEfQQ2L[gUSaE_OUSPbZd]G]L+DW@2OgJ7=^58_#)H5@dL=V59GZ4>^YW:d<P\
HTEb6bEPD-Bg=Wf(2VW[135c+MA0]5/L#?-KL:1/;;E[URQ+&g)3&]SP_QbW#KD)
1#Dc=26a6+BgNPD<gc-ag?:569N@^N2T]H6egZ]SF3#g4>ad7KE6)Z8@Q_KNB;OK
)1bHUe0c2g<]LM6N>2_&/fD/Ygb=-X,Y32.WO[PS]S[:>JD(1cNGJHZA=?11WWRH
_).W/C3M?9Of6g\ZgP2GH?)a]-@#[cPf05,abNN9MBA)3,fA/\F>A5^TG&-a3=f]
(dL1/1e;^OVOb),S7;.ITJV+6<1COX9.(8g.g80eaF:gP@fLZ.SA6D(OVQ+557Ec
/>\@^WYM^6_PB?WM#K+RObJV59)7\+[DG<\cD#G?KX:.V[V11f+?E#J=T,J^P?SF
HS[\)C==aD^A(g.a)R:ISS(JQ;,R\^&=U6+,2>Nf1>^8CVI>:-RO^?Q<g=T5:#XK
EO?Df4fJE41E+AcBZTa=;@)AZWCEW=dXS/(/>[XM.^=I8^L:=e1_S2eS,f_b3b^#
_B#_g&_&b94V.)O7QRN2PPf7(9)5N,4KF30Lc18Q5cf@./G0#VJ6S)(B0LE(L4C7
_-75GLfMVT)^1Z872>TWZZ:T2bD0_CTSf^O1:PH<ZbYR=-d,\JEEEbZaYZFNHL?6
F5;RQ0?d(dWd-B18BCAO?1,(@ST>(&=W4^,.Ba4+-aBb7&1Z_C-G&@a1NEb=_;>+
@N/dg8RGX8O:P+PI^4.WV18)DKA?8#P\a>8CG(aG?VS<12<&:WAG#V6-DFQVRNeJ
KbZ&\6AI,]QQe#AYV?cEU4)XG&bQ(<g^RUXEe^J#(+G><_Vb:O])f\E(<&_<A03W
__S^KS#fP,NfY2HX67cPP:.=_U)VXJ<QWU,Sa&]9BC0Va]>bK=C(a1RZ#3XCB:7Y
?2HFL?R:=&>5->9O&cM)T_]R6VEZ,NN<aA#,8O1S9LM+2O)<a,R@_J8]cB5IQ,8<
(3E;D+61D<^H;BE@K-18<_=FU8.,&3NSYPEJeZNS;K46D4Vddd3WN=DE=b0dFMcb
50+O=D1f#.+4<4.9MN+&I21f^T7UL9W202YM<7&J\X)]a#HS9gPFXDY\9U8-3W53
A6V7-,CY0?E=VAN=QGc,ZQ.g\e)=I+DQXMd]PU[fTV]G7J?6K=5<Od76,+Uc1VF;
[;a4+J(gbQf7M_5>d9-GC7JEeYb^(W#G.0^02K\bV50PFN0;1>8JbZ2RCcZ2XO<#
R+N_PM1J<Q[NY?Q7Q=VfF/GQ<TTD<QS]T4]RTSbE7FAB7IV@?g(8H-SIFdBHTC/7
3?+=#88]MFCaXT,,1V3I)NLW)QG2-+c:a;Tf,0Ib+<T]8/7:b[TGP8:27:5eTcfL
F-EUQ#DYe06YE;F<QWRM?RE//X6:@TI4FPDL)6Db\/PGO=F;Q^4fGEfQ3:NK5@2U
FFP9#?U3&9EO:D#44/2SF3:77G/g\R0@RHFJ537S-KVP[eDUM=4gNa\;)P?LSbb9
H5;e.[6NPXXK9L(^O]D;EQ[c&J#D/0HcP-;15R<eG1KYV:-MfP5H:U;<.f77_/[D
W(C0FA-4O0FIeSYX@J,3O_&.7Kd_3dMaBZ.RUHOT5=a(X2RFK3HGSEY->?^@EP)@
@<Af[C32>&>,PJ0)<U2N6FBM27+aGOe7_F(QSBI]1g#Q5+aYc0W79fff7@B?_(-d
48Y8C6^W,\[P?ZHb/TPLWW^#FXQKa[VTaRXZFBb/D=J<ed37:[I__aC(2J^NMf^>
IA#fEE03DG92WKF4P)#WaS_-(;e#3,3=]S#A-\bA)GD(:)Ta92M[cZ?YHOEZ&+(B
eX:gf0?OdZT=21/H0N:72OgU?TNUBZ0Zd#&bOUIQPBPK^]c2C:IO\=c4E5?V-[JQ
.<a<,A3>BEgYbd9Te+,g&RYNeE+_@+A\2ZDL?=ZX<LRRLfg4_^L62A95#R77>G]c
fZ]O0US+&VI]RXffZ<+/aYZ/:e^YE4AHIDg]Mg-4Af<EWQ;XKVQe4bE1YJfK/a)d
0>8N4A6]PIcD@C\7?)<GDH[f_SVH\4/RQFAXadY3bFE(Y)]-XJ2T<1)Uc[><]01T
JHVDZ1JdOGL1=:\gPM4WA&7K_5_c3A;Qb&]FYE&8cg95T#BJQUSP3FS5\EYQ3-S9
:=5)LJcZT/F/+R&#.]d?,UT<TAB4/gW8K9fa^O+JXPALKR^\VA0<H6774Ad3BQP;
DNGc4H.^;^_+IJDF:2dQ@U27GRV43f[DIZK@W]F=UgPc_WM=[T<gW7_:8K,J7;^@
>cI=[ZT1U3E1WYC64I=E7H\<:O@[4MCU,:7NO;TD6BZF0a:,+49UUD5R0QMVLcQZ
DVZ9F/5]38#b&ST)\?#=P0WVFdU8_08W&Zc)Q6aXJ5[>SP(]WBb8L.#=LHTE03VB
<O>OGP\/;TU8P8]<NM1]0ACZWD&0;(HaE1G(P>U[SYO9<.026T3F2US=+@L@4U0[
V7P34^WY?a?Zg8L?bRR@BMK4dFcV.41HY^^HS9W4_S.^V#0L,64H(3a5?eWG50XZ
FIA6>_e7?>AN=VQM:ZMZI&K3XY:3VPJ-g9a;ACBULS-aEEZ9B8c[72&\CYJ.[@JY
>.&#be?M4O=U3AaV4N>=4(DC.Z;<Yd4Y4MC9USE&(+=00[,7NAZXQ\/-@/YNTbKS
J=;8I^eGaHI)]+=-Q:WKI&dFf/Y7&@NZXVG2):)12#?#_F7?L?R#X2W8SZ21Y\E?
9aeFEXHHHV709gYaP]fbA09(Y@=GD-(&1<TMG0?D(\(+e4DNQS;Rc[#=0GY]^S/D
=J\YJJf[Dga;((U]5-IUQJY-AU&7U_bW4^=U=JG,AWB7f_D+URc\2X#JA3^E+YP>
0TaAag1VEd&:H-b5;EO9;eab3[,c:EPP1&CUGE:=3<I-8Y:E4&B?G/@f[1ae+?0)
5:cC4AV[f&2Cf=fGH3IL0+FVE1:9McB^I+0:<gJ:e.B=OK3g]IDb\J72N48(O;ZL
2PeP&6V/,:75[PYB+7)=9@16M2\[c\=L4d>6E@M/KD?#T+P1V+F/9W<98aVF#(_J
<Ke@AE2g2@A)O8#e@IfNRVQ\.NIb>D6?g)I8EZf?UJI.JcPQJ;WS?;1=QO243VF7
f=DCG?/2E9(WQ\&QIeW@cCXP?+8B,[CAPOW<Qd]CP=?CJS,UcB2/a&_Vf@B[.VV_
XF;Vea,eBeCVc[6GdM([C1BPWT:UB6_RgRDdOAU+=(QXL2SY][N5?X/^C1QdG&IF
?Q8&P_&90V;?5DXDH\LYZRSVGa[bE1Q@T52WdM(Z=1W5CX:)N8+E0B-V6_e?34_C
OA3R<IC+@)]N2@C:TcM.7I;UIa.8/9_]<Ye-A3dH^fB;A8S(#\7@)EbMM1B^8&KA
eK.JN5DBOEeX3;5F.W8Jb?6/B;RP2/+UF.fJBQMC2S[JG&OA#O0YQV.<#]_>.7/&
4LRD)dU=WT&L71Y5FU\/^g-#d@8W<BZYD9&C2]C]MA)Mbc4BE77(c.44=OFeC/g#
B^YJQ=?OV[42LFOKGd7Nc+B)&_6)TID#,,Kf0T@,2-F.9:NU.5?+bOO[4(Y.;BYS
GWH5F:]L(A/E^6RQ:&H786I<\5A#W;g]ffVYN?-))-MF;2W9],3a(4f,CP1A7,a5
=6a?/0>5_D,<f).,L&#?eD[dX&/J<:55g7BPOf9H6EfF(Ydd<5R:K7LFK6R.XU8^
&X=28AVI:7\\ZH.MVCC8URTVE9JC]K<-4];d8)60L3()6@0/4PDeHdWC[5D9c)#[
KG&Q4V[I/9[gV@=8>fb))a2N:QR?V\MJ]6X6+8QM03MXRZVJEKE]1HZST#b3ZSR[
AB]48D8Y8+0abEX#W<3dHMC7bZc]UKPGWZTAYHH+<,W_0\.R+ggCOHN0_bB9:KEF
&3+Ta:9<T@WfAeYL_B<N1(XB?YA6E+4Lf?(/:+_3P/H1Z=b:YVO86O3:f5UV;VN.
/EBF8:=/X?(UI>/4;gcaI3UHH/TV;g3?.XdR)dTG4b,4FZ(XZXK40_7?6^G16(72
Nc[&RO]A]#-2fBFYN]O+EH9X74K37OE?;HX1+CZ8S-(VGT2X_eO)L)LJ68A-[2XZ
ZUNA9ZL^>G<e:M0HVX;BC=5T,_6PP^cW7HIDICeNL_aDE(98RE7c(,3LQCS(e]#)
aGDFFXH)Q;-EBZZ9_0CbN:dUU_bAQPILT@DG[,O4;QdbaaV7>_Ga<]AW)IBIWa,9
<@(Bf9Be=E>7SCNg#4b5[/HZP^GZ.C.GBcdfJRVX0P39&+_ZJQ(]MN7<D+US_ceK
a(>eP9JN]-?UW&Q&MNFDC,MJb?=R\YD)<bc?TV:;^^RO;b63K7dcXVSe2,9DU@[X
5MEM]B)/d@X0,4,3(YgN\1?X@Sc//LT(.3eWa.];O^G8#HgI6/Ib]V5BY?RKM4RV
08d[FW7LK[_QJB>Qd(EC-/VO#USH0U>N:CNF;<-H]H(BA[W-_3N(B-L>8_I@0XJ=
[[W7D\?[8ARI+1W4eG_7?c:.GVCZ4TS<Wg+4G<#RC.dV(d2TgWVE&Q[2Jg+YQM=S
S=gbfc-QV(L.9-8.Y09&8I_]]E1fX2CV)YgT9]f6R(GVaY/,V22S.:_@.8E)7g-J
_1g<EL\cMCX<\T3_g;L+Jb[\A:&)8Ge.#0(9.<5HGJAWT033da/4&FeFYH(GHL]T
D.;HB5fEUF116,;Q5We_Y0GbN@7Y<^_^3MgDcH[9VH<&36-@F)SP=P,.0JacK.5D
^d]H3XG;Ed@[0;VYCTWca]).Jg0XY)XVOJ^7HZYF[_,AKed?f-DXg>P.W3?I)QZ1
VA;0.K1)K9?,#dIZ&_bM?2=G]J+2)dZM]b&gV8;IN0SBJH\Bgb6RGPV2\^52O5.S
g3dMGJRgVL^1]7SKTQNE2+=W#@W_#UIIT+\G95\5\PJNb3E@I3BfTB4[KWXA=55P
I]W@[f2M2SWU,ZDdC1V[F45Xe4/NVMB)7HN)SYIS0:\+K^bCB>A19&c=;I:LI+[_
dXQe=K?bO>0S&@A>D.H,1HA2JOL[9Y@b=P)?3)70+U;S;g-b.K#3Y8Rge+C@;:HN
X4a3GS8S@0<_b-FG-,>,\1D4)MfAc0g]f+PO93g+:^Q\3ZSf^XD<,3eMH/g#A_IM
VY??>dX;M7Nf1FH-25^gW=6CbUYR31-c(6Y03=e@d@@2_GWe>]:G<>6[Uf2EHM3G
(.[?ISS=2>c):0N?)<f\)X/ZV0,-0TdC3DRQ5OQaL&4=27Zg:_]#_Fb6RVU3\YS-
=6MT^4L1caa;06,dd05Y[>&2<UDLJLH.#D:JJF(Q\gbQZ7GG<,V.?TY_.Ec_?KX_
R=C@5#6,1Ag+3GMAfLD(YG&L3:\D)EU=,ecBLK55^A/BUQ?>[I6M13a5@&,,HSg:
]5b69W5V07Za3VA3VXH+6P<Ng3DJ@KK#B-f_F^WK=-S^1>fP45GTMbDHOg:-1UP=
gU>SJ/&+=N^E@8:H;.MW5f)@.UHC4KY)Qac48)-Y32,&?XC^dCM:cN._EWD8O?AL
@[E@#[UNdEC<Gc.@52,_YY26dc&O<681.^QeN@EG+6]Z,XXR/6/\aZa8S@^-N8Ua
\TP)QG:P36N<M7\3;95/WQK_;)VLC_1@BD1)?YQ,g@><K35g7b6O2]DJ)Ze4KKX4
2#B)>bCd3Z8(11LX3<^=8OFUCC6O\5R#gTe=4d<BY;6P_;V6P&dB(S4?\RAa3fZC
)>gDXRbIJ>/NB<QXP<MDEM9UMY]+]2./VM[dK&UXYFA8NXGYabNFb^Z<a8Lbc=TA
e\0L\RRKbd^TVK=.a1BaQP?,YS5&VUd(44W^SS43=4G<@-AHKJcTL2_G@4GT7W1_
?0CC8A[HC&QUaL0->+<bIeHf;959c5(cL;,,O=][81S;9cI_8>&O]aR?\Oca,AbX
c3,#+&(4K+&+]UY(NN\WOKKe2?,S9EaZ8T+4CcGVcVN[bb:T-1WU;_^HVdG^(.CF
7@dQ;T0C-E:L&XDU(d=F(Q_FT@gG2a3ce,PdAP-T+0<:@_)RMd:_DK96J?:OE^IA
2EF89N007RQU?W,?EE^WWAH[g0([e3a>WW]PIPS574?+^032T\CE.NgLTUf;]N^=
?;(,fAX:I(-3fT?VV>6@&[1f5Z\JLJaQUR^)K)0B1^MCa#U;LGTFO0T#a.DOI0@,
fFDCd?b_Gf,_90A&d3K>.LE[90+\Vc\#B3dOXJdMNFYDV):H5O<OZ3<]N(e:^;DK
g[2cOD4Yb#aG(UP[=d_gWO+F5G4,4#fe;d608JZedJ(ZIH@X,\]9c911[aAVU-VM
:XVB)4+7aZ659NLHWJ5bY7gMYBB1Kf(gLM;f>ZN&_K^KP>:F&63=c.HH,GCad_5\
Sf5cCR5N5WAY8bd&G/@:C0IX5F/QeZZAb,Z^>.N[bGL;2<C\E6TJUX/S:0\f=+3]
Q2K4#_6D=3=eIa]fI?/^HC_CE@-d#YR-aTLa0]^<<95B+\33;6R6:<Ae70KV?b;_
3=.F6G6G8D,^f;[T^.)/QY7Q08D9E5f&016#5<<DYQ,A8MWK_,b]BX=>H3[O8Ded
Le4P4eP1Q@_Df.+3V30<@YN._G4ZH+fT:Q@)ZLeM@4N:Q3DR>?GR9)S)a26S5ERC
Ndb+fU^Z^5:N;7O9[-JT);&22FRcYUPJ74UUH9=F.?Q7TDL,SIeBSM<0IgBa^=HS
[3N1J._KVaFaSQ8XRQ&-.;PIDEGVPV2G5@3>cCa/BDT7Ke^Wg9c#F_3O7^#GV3AE
_;+;&LDQ/RAE1>(1=#4QB_6Q_(AM[(1@O\-.BQMSQ(;47?&cIMW:-+H78<-]>>ML
(P_6.]Rb5[?H\Cd(cWN)3,=>DKI8[->U2=G2Pe<Y#(cN<=:aMfP\Oeb&QT^1Aa6O
[-DRCe2<FSW7g=\HaEA0ZK@8&6\O8)+Tf?[B)P?b@b0aP6N]9=B0:ZKV]e^fWFYd
0@&<SGIcbd\\^@@1T6bD1cVVE#+?^ZG9/JW?OccXJfa1^.3/.+ZGQBa5a[O>7NM=
+-L?DV0aF.2/G&2=2/@]<ZUYXbVT\NG;((^4@,;?95ED5HLa3gZ/IQaaZ2Z?]/6e
;]DWLQ,VJg.<F7\X-18c\AGI[02IC9eGL,[MY1I92QdFM+,8cCO\.?,76Ec]R4BP
?CM\eWIEM.Y-ZUEI8J3_L>W?3NK#V9c9Y)dG(PA-0VWE^V(3/6_eL@\=QNRG3#FH
@NQ1>=E:VUVZ+7dIOJNTHZ:aL/<&7fecX/2e#I]V+:7/RO+.T[T[>3^9fOb+^DX\
M?E8efIJT<RFKRS>OIKS8/)ZA-^+N\A=VY5<2^+BaT?/Y1-I(E1SK9N&8aJB10-P
\5MZV7ND^Y<@6S&XL7LJIO0J[MC:O.a:.Ia<FS>19:D(\^]&IC?a]NF=S?XRF4J[
a&.,+Pgc1372?P&3E]<(EaQ</0=bP4Va2TL#e4GCYa++5a4ZONQ97P@5Jf0(&.d4
VE[9-?M/c_B/[[4cJ?f;U_O[Ef0WY7Z@gbUWTHgeb@aPCZ\/M&#c#:IWF=WO#>5C
0RgS\U6\=\])HR/-[8aSO?5]4FdbE5=39I1VVeNg3;d),fOe2\cL14B+3GGCUeXA
Q^8dI3^[6^FL@B#BcUGWd8LT0KJ6bNebM#_=(Q9F;:RR4_dB4:T+EHX<^a+f9RWb
\J]CJ>SZ6Q)B0./PVVUQ6N1<7?MVE@,H2ROQ.Y=UYPC#gFc?C,E6FIOC9/f)C:3d
g3:))LG;/CWBP#=:;EaYb(W78:L136/9]Ob&/Z=8#OI]27X@7:7N9P.NPb&R+3YB
QAQ96]Na[)_AC,eagI.RBU_,@H2&XFKROG;S5TKVG.R#EP21K\:98=M8@Pbe\L4L
9\X-R>8F8#?N[BPRc[9:,VYWB>Q9,J-6IXf3VH,ReQ^f[/a/[WU4CP^Wc.3VJ4L3
PVYbb<3]DBAC#M#772b(V5Y0C9Y,ba7HRc@UYVbeMMbVM#X.>_(#EA1\8R0P9.#@
P3NWS/NTPJCfVD^d?Z]R-_=\XV<bFUT0A;PYLga(\J2[[#f4g6O.KMg);@b#Q:[K
G+C#FJM=HR[;7^5a^M80e<C<ag?6&?L;I)<]Q8#>VZLOU7E?54e;_1M.K<_&P0A#
LNLY0F<H^UJ:AIaaA,]5?)ag^PXL73]X3L:#cT7:+29OY^\<B[<bL56-bSed_6SK
<,:A^O@N@ITRGA.C[=\]9T>-91edfIDX@J>Tg#NK9bV)PZC[a(KFc2&gF3^MGRPa
J7fbN_VW_e7E&O7T<<d3ZD8Y+Ya^9B]^+&]-F8II-?0f[?HCGEdgb<HAQXQ/gY.a
HN+ccUg#VXZ17?=33c:?cRL1)fcbce;2-;3Gd:2d.V&g@QV&\;f21=7eE&6UF_g\
&.f.,?+,2BC&0.+aSbBCGKATd2aa6:4/<2#@,9FU47J_AS\F[I4I6CG./a1XTX]R
K,=_Jf9]=B(/62K5@X,M]eG.I/AQ<GQCFJ>UBKbTTRPW?<bO&6C,FFN?US)ZfE3X
?b(QW>Zd>J&07JBFPZ4EW_9<+K/fe/084P.7Q.e2J@^=4>MMe+[3TAP_,1#K.+OH
UH4G6W>?,9S.,agKR1gVVc:5926cB2<7S=26bX1:U3CbRJ8:dc+C_-/?KccR^0>X
F#EJd,,6-]dM@NAN;959c?S11Q2PFO362XME-[DQ8A&H7O;eH[(We&:/Q#IF>KI]
U<44+33(5<cQ2bfE^4,S)e5]4#U-)B/\=2+)Hd1JOYeIXWYc\FIXU^0>Qc8eVMSI
gRN(Qa1R0a<-W1S&fWP_9/]U=PC+]D=<&MPHc_eN[,P>Rc#NHdZc,XRJB@F,8DBZ
E1FKE0A+./Y;4842UP0@)Y(Q7O4B@1F8@-g+2:edWX?[][MWEag0(7I?U8#GdM.)
2LTLL>g&baK)0E56\d[MZA]^bO]=TgEgZc@#]:]Z_RH,D?6b2FdPR6?P)^e8g9.+
[+K:XP7>#4MKggKH6E[gG:LNH.4f-<<^5L3O/.+W(U+--4D(bb=-DFgNYL1dKY[+
\03&G)GGM^FA[/WX.#)f<<dIbPB;/BBK/_eg\e@UMUF/,NH0.gU5HQL2FXS2WG#O
JQ&,9b:I7@X>&L^76?@AOGc.b2ZN\)g)W]fM24:]/9Ic=f&=LMRB=bU_>]Z7/\^P
?;/4^(^b;fBY3-#bI-+HVGf0G3BM-7-[I:Kc7<gd2YcSZ(TSJESVNCTB&/KD&aKc
.YV9H?)<aeg@eQcL80d.:a1aP-#L+../]M\cV4W4LG(^(VE,Z\AdgcaM]FS9BFf3
IF=52Z:BY6?.,DTH;CD^J:5@^0AVIMce>RJCXWRW/dP[8K-9BF:HKS43<-:W3M0@
A>B8&:[NbTg^9P6Da+RaKXB)?bO/<3eA7.e?6X)?@6/6D;/CfX&5Q1Ke6BT99Q[8
WZ[Ea?HZ,F+OBZI()\[_E2NScB[&e-CI?YBAU=SUQd7P4KUR1?CPS+E7#O5N^T5L
4:U&SS3&DL,,P/^04,P5H0Z1O=?R6?OK&Y9_DLB=Bc0CTS]/g>D6UI)(S6//Z@g#
,aCPB,CN3#HHZ@JN8\63GgKXL,14dMF/<-J&d0.S.Q=6\](&048-?A?e]fgfT?/[
dB)9Y?=#E2gVKJSY0Q6,PM]N=5-:XMVJed:+.LE&#EV[>[d-<S=?=2;f.;gGL;KR
/.0NH0FT\1R;]--adLM,EHIVI,P0D&(_Ed_NGeFgNO\1;=[LNOSIY.b7H+T>(J;.
0d&:cU?-/IBP]3XHP)=(93TQY&b&\(PdCB2C8W@Mg,B&E#D-XF0)/1[[Dg6-OEfQ
H+]PZPDeVIQ@/MYTPZ)U&2-><ZL]OQ6UZ@B.((TGCcG164egTR1NSfb=QdD/B.3<
9X1K>@FcRUf5HV+9\(K[?>bFAFMS4Ea&2VO.+a5J(a4X@@O6Y?O/H@\Ig./[9A[S
LFHFE1SBE8^:..(#cM]]CP7Ue,;/81-TFc&/e()4&S0S)Z)D<3@eaXD.g?\dL(M[
]L[9TaBeNNZb;(a[^-gLEVfP/_?VQ(^,GEMW5DbCMg.9=67^G?2.TMF9W;=GZ6=X
KK#^(SH)dF5<[P@cR5e[&ST=C2a1d7TS)[AOG==:@#8M&8^Z@?7-4Hc4RBAe&_IO
dPDfL;5RWc))eDIfF?8-QW=@PH<JH#.@BZY&F=@WV1.1R6OUgaH]\]I20DaSMeBg
IMR678@WLC4ROP>;>?L^3&7TUQeGK=.^<?.2QU:MS]]>C,Cg)7DH0<f7@XZdNLW8
+QB+E+R6-3f(MPRKXX>#-8F48eFXeW(XBRdP#UBR).F2>Q^fO-IZ?VJ=UF=Y\:D6
;N><.W=9b>Q&<b(Ab?DFd&]gba7I7?+#[]#D\g=8GVE\-.63]LMDIdEJaZ4^:bVP
+fY8[8\4b.6?:=Z(EY^N&4^)bRae>3_(6\VIb&VQU,MdRG3EVKeV[LQe3/[]_H6J
3.\6QZ)eP4TFI/gR]/0ZZDYa@+A@1TW]Be@,=H@^AJ=#+G,,>N<c,gf7EMUSF):f
O:?Wd9,YLJ?3IbTR4BWOBWQGTf3#b^76BH?QF#DJZgF5;WX?eDbfT74gga6X5P_7
SW-0dP)ST)EX#IX9T5FfOD.(25Ne]IE_O2B._gZ.P2;T[REM?_#;(3(1&VWTM<c.
6#SXb>3.XIa?CBW6UK_]H2\/&=Gd.T4V<CX<,g[KLX?X0&@1U_TBEGgXYEJO?ec^
fc;WO^VA[9;dBYE@,#c2O2H-eaQUb#88][;G)>;dX:d&^/W4E\BPVJYBEL+efLQZ
5&79?A@3YRKIDWG,IbZ^ANJ^V//2H2.c<7f2EJ++EYTYPMX#,>HP0ffXPG;GV-A)
K5U0bM:D)^;C/QX7WZ+ALd,2V=QOYR.T+LR#BfGAG)?d-OKVBafbN,\AgcM7QIaZ
5SaK]3SLdXAAM,4LQ=WW9M1FX.QcY<J33FBXYX>Lg?VR7@W</d;ZO3U@ST@ReBTc
(ZAEBRI//ceO4C9gBO+.+V=DQQL^G8fe;6dKObD+[=9OO(]aJCK\Wg)OUH;2\)e5
+BaPgKK606^__;PW<Q^3KCX\eC/]Lef_#:/@4E[7^)+9A>)?P:EZM\b4QJCbB=[M
<HX]FDWN3,c]<\KS:a(Q7+B4=#^.R=dD/VR8DV]Y3[E:Wf]aXDVURCB_MA=(,K(.
79DaGFb>7)]FNJ,c&#QDAcG?Z1MO,@#/F<&/.3ULf,V_TE?5SW@aU7N.21LN6=OT
7YC(:5;[ICTXXZ[<\1;?X6g(K@F1V9=f]f_bgb6d(BMCX\dQ2)bZ8#(c0?IIFFaU
4Y,N_4F7L?TL_19=_Ocb4:;K=B&[dcYL0;ZG?HO2R^dL7.MKL]MR#)/U6/N5P<XG
2C3KWc7Pa/,RU=@_>Y651KV?gN)&bXN>D25(gDJ.1=2IQJ0g@4c96cbLRJ1T6/P:
2UWY>^/LLZS_]7ZO+_4NQ=)QD#VSeW:.PI-^(NJ2C2D<AW5gd@g^DRJ48AX]S39Q
43fefgN)Y7gcH0;8<BX:1-V1gT.VHDS2<V.;e<38gRD?MG3;B310AZGBVUOZF894
1dGU=&2cJ?+g<CGA1eB##Yb9(?d#acY_]Q19Z)V+b#_C0&C[00HEF58N:_/SNgYL
]fT=F:bNeOeT2X+71cBKRbFReAfIbE?BNS#W^)FQBc0f/B3;HBI17Z?A+#O>;0gG
NB/Qb/#.g>A@(6@A((F84NAS#[SfRE/)0gRQ]7\LNH=ad:M9SX(2c+f>X?HJO^YB
2I+BgVf&=N#6aPJ2ca9?OOFfeKZ[<-#>F)BCE]d=C8D>W>#]X+EF5?H=8_4=c^Z1
_-.SAYa9C6;8^VV&;C(f=2Q]gSKfQ#Cf?Je\6]9V=;OV=^F26D@]7:Ode\]Ra/=L
?2#T9b\)PNQUV8N4I-BD+V1>NER4#E4LL0<0YcHKVL2H:)CWHP8)[>0@THXYb#LV
RO?K?1&+6;B5N[POc:aO3+8H2[>\^,;C#I1(IVZD)YPgf?581d:3(/X>O^5Q:WM+
B5U>Je=4gV-gIeXLYcX:?)]+::FV&UOCTfF=(W#E[[=9-)U,9PC:Xc\LJ+a/>Nc5
gOZ/1OGE5#1e#[[PgbCC1AE\8[:R[)S<1_7CM/c.G8H;0[dTK57Q^1->6D2[dXIX
FI,CFHJK\[TUc2?=N.^RS5?H\2N-7W:#GTHf9?b[:P2TOb.cc1?_;d.=Pf>)\9O_
4I=)CD?B^W&DQbCIgJ8)M85RSJGBSMM6:B#:>OTV[E5S/B@>:N1G=O?MV;aL1?f[
9.Z5V9_/<N6>.O_&?N2B?(MJ:[NTG:8TgD.OTg#;N=ReB0(W1@^H>&3>;S:SGI.1
N<O;(ZSKK@:B_RT;dFg_MDVB(ST/=<]7<>[<DfOFHafXP5YCFGH/QVE+Sc.7c8(W
[/ND-E&(4d3OY1JW#Y0A_,2]CL,I<fR[&AXP@<B42;VD)JB5QCH<M\gIX)_L,;K.
L+@NfgaZ/NTE)M0U/#4A==1H3[+aJ\MbcXYTRVbOI#=\3bL)[U?H=+Q_^7K/)^5S
XG_+0d<T0fK<WN2BB:UHW=e?Qe7<&fLQ978,f;@_;:WJFA&HIO:9ACEbbc,a_9-7
=+F?TQdCPX^=TBF]^/9DVW.8#cNdH[W]LRf;GS_9=XB.4W6d_G1LZ#S[=P;Q+7KT
K:acEA06AN1.(D5#U_67)GX5YR#?SOXa1.4aJYFS:&Xe8#Zca;c@\?Pf)]PIYcRG
ZH(EBLLgR:(D?HSfK1H_<9H6PBE0A=a,IV]D&Cb=W&aOZ5L3\J9e:(\-+/V2]R7@
L,P[9P,JF@8VKCDe?E,7F9#OA+c6WZU<8LF+?L@U(cX>LK),M2(Q@Q?<L6..LM_;
>CBe+K^0CgD/?PXRP&_1cELT4A&IZB/;&_KU:aa:=DAB,0<Q?+AB+Mf97?G+bM]-
]DgQ+[=/6aMGGZ@@PAX\[7[P6J9Y-D+BD]SLa0>eP&RNSK]K4_XR],cX[Q25CB6)
)W16\&]>I0&-):;dEDb5O76>IKg48g,>HNXgAUZY,G0&IKE/F55TIX_2BCT]Qc#&
KZX2LSM4bedN(dRJ5HO-AVO(E7.=92C:?]fX>Xg-\:X#+;J2>I:3S>KWUAHBWa)0
H-Y4e7LO<D:#6\+2A<N0WN3F.3+f6>+,>[YKX9dSC+O?.ILR?+GYW0KYD@7GaBd@
<(GcV0U2@CH/34M1@B.0bAXNW8_4<2VB8K1:.Kf&?O,G=I-99FHRG483GW6.E8O9
^KFd>MAd9O.(a),^6P1dUO//QS/8g-LOV/4;XL]T.Z)P_59>0<Oe\URB@;X,T:1=
AOKXeUDTX,.JF=RX&PcABWTNaLK,DeJ60+^P^.1c9f2HM#g>CHF.?Nbf8&J^DZ##
Z;.(&&85;.8Q^Zd^#aP8>(+K-IB51a]E(W#]5D@S))><0\3X3f>-QYD+b]>M1<0K
M?DR,YIF7^RcWLBcGc\4ULIU\3OJ9MdWd@Z(:B5)XLf^M#J29GD.J3-eb3\N]K=B
@M4&\L13S/EA(S>>?^V_J[B<-1ANOc^/9Adfd14G9E=VS5P4.dFEEYCI&0DA)LCN
:&T;\e5MZ#68OMJ6N\\?>-)I_)1Aee3g6QW2]PRRZD?EBNC3\MW=K_V);P?U(2cQ
-5&Y:(fW&9L=M&A9=\ODPMK&gfffg]OKM^9MA?[58gg3>XCQ:U)/^=,SH3/JYB-[
>WObbVY=5;L8]/N83.?2ENYYM;E-.Fb:2L27C2]7M/[6G>,.Z,b&)0VH.U#eP5&c
W&JR]]FJQ(T-V?Z),L.&D_^f8<X6E=GHIX\LF/[I0a5S.H0XbEXc@EBX7<EE0G/1
&8XgV=0Y(8PfdHbbW>fQ^L3I@?UM]PEX7QCF&8F-^/WAIQbe?[SUC1&]1N]D-5]+
_3NPX&3#)OT98=51/KRNZD[dFFc4UF^D+_D6?f06W[ZH7^F,be0PIMQ8Z:Y)-?LD
^CIGG]PE\ZUGHM4E>/:dL?EK/(:_O/P#C4OJVHD9YCfQNATM/6:CB7J5a(0LQN>d
PFFMdQ[1)e+g?V[MA>4gC/_(PbF;).MPgZU6@5cgY/OY[_9&L+YJADH1>-#fNg7>
JKc#SXO#\_PTFZF4M7d@BaQ^FZ@1XGeRJeGVZF&e@>_P29cA2JYaa2S;BN><ZZ9]
W+3QY+NggU&64(&/.I>E2df:;H0-AG_5RZE.Y3_NF;@a1I09]D-,>LH+>J&c1O-d
DRTS8UTN)cc@?EP;cG(MYA8X>(GE99\]#FL#<Nb2RVD&;?:JA81-eEgX6:bN+<<A
@?N/:e.2>Q-D:]]@:#^3A8^<;3\g=;c;78/[bZW+827=ME0BaaE&9Hb;?=:MT3H_
TgAZ,VPX_/W[GB5deH?N09R7+.]E5d/PdL/2Y3]Fb0cRV77W3#<J=?3[JBA7HJ[;
=_IC[&(>?/bf=)2LN#=UK@KeD^>M.g/N7TfFGbacB/.F9dO2803fRM]e)d-@<.c.
1XEF5KMbdW0B3TXX(Y3EGPE+HBXZM+L/:2OC;6+#9]TZR>]A64/Y/S]R5;a><F).
YQ&Z02=dMWf@L2;<7_RL)0OW2/>)]\eKF-;3NLcc0@3+I(^5ZA916f=9)U4.7(US
X+@)EfJ&0^/RU#3^(?:?/QDPC>J@0:Lf4L1?aX90Hb:HUc7R3(:aCD\3Da7K>->O
<gWeddH@g9?VNf8=VK<,gA@aS:5b)_@.[0<fW_-<+4YFB.>JH6eZQ&b&M&&W69g+
0Z/94L0cK@Z>Ue5.<>A#eNO_D5BH,=Yc(Z[0KaE-&+SQ5<@1WL]S9P#M0LMY)&fH
5+)ZG.3@@44SG)BTAbTFU^4EdDOba1DX6_DO919=Y@FK68WCO5(f0+GQ(MZU^6[@
9J6V,G,=0W^4TN0#SBY6(GBWg7LL?()P_^1]U7+F^<P8cHY0b+FZ79(f-BTeEL\N
;.-G)+WT63H03^^N)SWO-VT;fENP^baDBb@V.D0<BD.(+d(BK>+)25@M&;)?7/L0
/5K=K37(Q53La_B>CKe\.T-a+dQ2,e7YXbCB?.0cYX7I-)\T#B8/+G0e+@30(MHQ
CD=a^;2,^B,2E^#VO^T0Yf+<73)Wba&4M+2TX@)];+.dgW5AW^Y#_eX=(]R\YA@+
Pb7DB9S#AA3WUR0IK8/GaUg9T^X9]?<ebaE@KHc;>^3SMY<RJaGa?9-<=gX+\c,U
aS^X]DOWTI/AY_.;^8,8,(FRB0#)CFBc=ZGa4-gD3cH]/247XGOA599YY=OP7T;A
cBLMRKEd#dA:b#O3ef6K,_<g4=KU4>]7UEADC#eeMJW0Y#c.g/?Q8#2E(WeH>5.>
>O_RBP/N?>0STWKUKU=^bD##gXdPB0I3a@L>fH:b=ORd\BUS[0V]IHDD5Q<IA2f9
[S@=J(BD(b^D^ACUD7K6g424F6Eeg6Q.9SPRC#(ZX=TN#7]+)51+[M0Pg/R/Za@b
e-#^N:U?8E]QE:Gdg[,@6BO(GAbFXV>F3<,2Sg<(\(8fUcU):GTB&>Z>JGGIF^A,
bQNV=^JO+O]XSLUF\]65-=2Hf(B:/6IGdS<T44WD0BOY&EYF6@JE(1LO?PIQ0#QY
+\<+/4Ie-3(SQX0c><LIMPQH_3Y]TNfKTUZ_CfSNeLaL?;[^_YYPV1)9I0Kg?](K
Ba_/Xc0I:b5FcNS7\5[A0GBT)\N<B?BHb6\.0RH7,0N/Oa<bcA>F.0TA-?^>&:bB
ff)\OPgL[0ad-13/VIb]E\R<<E+?(T&?1J&?L)^U/RfW>Z4NJS2&..C9>:1b61\Y
g3TD]\<5A+dAN:F=U1M15JTe:29RU)(<@3(Z:)B7U.-N9Zcf/V@GT?=#M,.;+5/,
1gE4#BQIHe,JV;fIg\::M(W<KHT:bMgK/W],EQ(M>D]6Rb\?b\IPW-a48=V_XV_N
&?e>:1?dF/eXG#Ua+E\&J)&<U40UJ;eH@=Z8cYFdTFIU@NUZI#<,E@-?)F1<O;2a
(GC;-FUZVOd0>eg7@>:+:SQ28MI-DG;FQ&H50.R@76/K/A\&Y[SX^Aa#?9<\@X?(
1G6]TIg)+A?T_,OQ\/FYXK):U-<J/[8GJX#7HV0&4]LF;g@><TRDQ:;Yg-d5gM]3
]/F5MM8#X,a_2?QWaFfRMO(>bI&51KGG9TW?W&H])2IWLH])/@c5,0V8OQ@6,<@<
Ga-J,APa@]GN5DdeE6:+4+O6e7NYRZTf<V5_FNG_S_VG/(7TY2c4N;^,,;,_&5J]
e@F;4R)JD(e#:fKW?GMI^UJSA7?,\BHN0bc>G09:GJRJ>3OXLJ6><^RUc_WV:FRN
O^Q9GS_)(/gQ]<IIS(XFGCN]QW[1AcfDQ8F><09dSbMU01;-3c?.2dB)(Y@EU)MA
H[JQ\/dbP<S^d==8<7]gU\8DegSSYHZ=YF1X&\+;?YX2O5[P5CfZ?dQLJX&N;/P/
WMD@Ke^\82B6eD^HWF_Q9Q8_0@XFV@BF7QSXc0:9K?)U:Wc^H6+7)OQ09QG>7=#^
Cf<[;ONICKDMfA:Q\T5gWIWE/gE2.aG)ag9;;4YW\19XJf<@gY3,GI?KZe(52>5d
LZgCLSeC)Q)A1V?-A1U3/N1H\-<X,N;<=5ga:5G/<26M(&=NK,YL/Bb&_G^f<[d[
9MK/9WP0G<4S\.JN&^#H=T6.7KRId1KNSMf:/2K;&MadLN-(B>SD?)AeK9H?HDVE
=EKfPVASXg]d31+B[TSOOa6&N6(;^A[AJ3&?RZR4I5Qe8S.-C+>NB(/3^W1<dBX[
+gTG-V>A02-Y;_CZP+BF+D#(#?&O)ccF1.SS6V4T::RA-HMN7gRO\Yd4+J>cOg\N
2<6DV/Y>THJbRZ70R.W>AKEP[:_F#PJJIO-WDU7[N6/(<A@#NM7a2d0O.M/7?3@>
061QNYE2[UN>RQ\I(-[Y4eWQDR-@)U=N&V[_O<#NK+>/_Le2@d4G8XPH,+DWe:\?
94\J&^/eac0cR<7;G>@[&F;d&4/bSYS(@e#@T)>Y@&0S-JG)F7g])1&<^]&^M-Y=
Q0X]MDRg+PC(QeG<\f,J:AN#NC7baGc]2X(8GFa4UT1R(2_H#&7b/5O<.cG\DJc^
9V^66Y5T57Xg(H:)7dcBeWReG,UgU<UT-B]3>Qe3C<D2[JPQcB:T_R,)a?+T6ZJG
\EP:S(HT&g5F<[I(Mg=,BCe3@\W_WLU0VHV&W6,_c]QSY3Q=BEH+L,DR4=e>;A#_
)b0.(2L6\6=;[=VA?MKB0I:g2;M=HHX[]HU<(F^;Z?X6K3aC[J(YK+^]@>&.R8Y]
C].YU[^2A&^J/)Y))HTeTQ/59N191MgfTaId/NO+Ae?I7g(;YD7R+973Md[?P@[@
#PVAE1>gS(11efYRU&X3\SNEY1a9G3T9I@@aXM.3eGMW^U&4<.LQBbT5V#0(4eYX
FQW;,RP.[T\DWL)QU/(-<]Pg=H^P#L^&7-cLFA9C=gG5CPcff5]Y+/#GQ7:Hf2>=
BUUG/d9+SG\Q7,^[4KDXVWg[K\=DY9D9f)XJ>1Q[-bFN-B2<CP?_E/Z4S#E:W9/]
fQGJ8RJ0;21]<_/_XQYV;5U5;A:MR\^E0M0;&)Y<,3dF=V\IPd1D8gbXg78LcBG:
ERd,^_T_eeXRI42X;S=:4EbSP4@BgFY&_C(&I[2K5L^,:R>_W)52&/=[<=&8(]/J
<RQ(8_9R#=Ub_N^bZD+]#OgFHVcZ\1+G7>=1MO0H<Qf(J9ff?7RUeY/QL]RL,R\1
ESK-A9daM+DZG>N1XA./Hb,CE\fWL:0Hc;UFC:Y5=UF#U0YdVR;]e&,b3BeUG-[)
?SZ(V_2O1O6dR21P=J99gbW)Ce[2cPgN^Q7Q4-D&9Dae^;X/==1.=AZP]0P.8I[L
G0PJWDU#(RW[b6((/cT:DD4&-;C3^c^H&IAWP96eX8@BM?#[395;X&/K(GOcSgWT
M<?07NA2Y9NbED9(@f[FJWO+IO:d;X-Y)D@]42H(TVE^Hb\/)7TOQUER5X\Fb,9W
C8Mg#KL]_6a&a.Qa0.3THH@)6P&[>HDgOQ>S-dLgER1[3G^F:24OH0N6E(/gR3d=
7E<C^_([]La;\J:=O=-RCUbSgM+H_eU0649G5eW^N;OZTIB@N?UV?I/NEe@6<RRT
&#J2L=^;@2PMDRPZQ?\XXU#QW=aHcW<.<=XM#If\DL>?e=O#1(22A.9WU6Q/TG@(
a:=JHf@^F:Q1&&&.aN<1[=@<ZXbYcWZ>R\VD&YFW=Z&Z7^6_(/W;^Y6U3G(+1P,L
B_GS((DUI0>a<7HEBK[A<5RT8cbZaEXL8g<;(/\>Z79SR<1;0bZV<S?JQGF1<;\R
4fbHWD\FX:)UIRGHcKC,^>)^F2#2ae_F)D?<PQ20g,BHeFW4b(OG^d)PJMFZZP@T
cBB/JMPQ=UH23W7YIb2VYL(&+4#b3C7#\bR0:dO2;.c0Y&bCV>Q3NQDD22/X.0;R
MI].Z&&D6B8WIa#WX,DGA/H3FWfa9MA??+;_-2b_&5.D&4&[L/aXdF[G+20=N9P8
)Q7N0<N_QTU[<RfPQEcX6H;dG8OS#.N;GZ.d^]KaLUY&A&dWN<[bPFB]ea4EP;8C
HY:QJFYe1T+MEf8/SQ4b5J2&4+UBOS-f]U#;^WM_4TJX+&LIUUD_ZDKENfbNA#56
B)\K,?PMP),VMN^,@d2c05[e9(0EMUECdbP>I4D_N[6.UJGH#L4Kb)RU(:Agd51>
Vb)PX&POYg.C.6^K4d<>9H;R[YA7d.2Be0AKdcP8(a;9Ag>89;B+2@gd</J;=eQK
;=+,>Z=2FeQ^ed>d]0/bUKR-V(?U]#6LNK6<5ZS-RZ=_4CbA?FJ[OY\Rb<NJSAHX
Bb<=W(UXN&10G;]WHgYT?F26)@Q:[7JJTA_U+/]S^)N<4a&6S&7=PNV/M(]YP.(,
082L.dc0D\61d2837RZ;+4RJRef7R9,^0@2WdgN;@+Y^EbHO\dC.PZ5X].<I)L)J
Q_^0P0JZDA.edE:5\Hb52,ZWPcZ5TV;4=Ld<eT\(XX.R.ZL-22V?+4.g7)J.S7TQ
06Y2.1R8<;3QZ6Bd?(-=cXGc9A_+-,6EFRI>KH:d+-(SH/BY87S]>#1<9;K3;K=1
=/DX\XZ(/)\L3N97S:^L;>K,QJg-e]/_W85@g?Tc[[29KARS778MeUCIgd-Y2;U0
@3#BU.PbaY[DIHE5^;+1EBB:T+/=V&8#Hb@)]NBA=bUP?DKF>S<QRP;XGD(\)&K7
E>L630[2C7S.^OESIR2SUKS4fSWMUK&2RbU+&<[eZ;CJ=FZg;5e6[[H<6)>G4c58
B@RFWVXZW:d=BOBOVYYMWB;J?N:H_ZP-#8=50f3M=N3AY17Rb1V(^YI9\[@VYZ@C
)H[39FAgDfHDL;YLePeDRKSfPgFW1bGVd>0EB^^C>-gF@WZ&I;F9@->#IULN\;9G
-_)_2K#Y6L0-S62U#ACF+.\f;^R):&9^/;_[ZMS-]1([f9)9@6TZeQQ;_=cMB+;U
LFe[XBNBM=cA@DY?]^.-PbDYBPQg<FbgP?=A,])DN<UZA7f(&V>Z0F[4;CH.B_QA
K+KRSICHVE+OKPLD;K)U0e#G,7@Yf)#A2/5#c^cP6CfQ=DPTDgX,,KbTfL&#<NRc
<)Wb(=#JV;-cXVA@A#8#@IPb[P@/@A167>a7X_W/_I\>PN+2a]e8#&0fgW#U@4QU
Q]5[\@Y(RLG)+O1@._.Ug&^GDYI&e\MNHgBC5ENMR0XYb@>YeARU/8e7edUZ)8]g
-82ZDXESNO2N))M>^68&CRY5:b-97G@aDdDX@W4]HK=8AQ<R(+2G7I<M5;fM:=C^
W(T<db#D3[DG=16]>cIV=+MC6NF>N[@f#RO1Jc^Z(VX,/2Q=<E,X2C39\HZZ7Z\O
^E-/5Za&;@GF(7MK6SdZ]U(Cgg]NW-(RA;-7d7_CfILZF/GbZV\DT3UL\._^2(86
GW4JHRQJ(Q2>NAP]S4//(Dbd=B20=13IN6#b7)1[#(VgGE<68QSB#[HQ1@H[ZCJR
;>V5a<g+UO7]11/E.JZda&MdS:=I<8IN5S&9^R/KE&N>DK5F<RE_2&B9D]e1#W@U
9Y/2>\4DQ_SZQ[bU&H6]f3NE2dVS+1V;A5L.Y.AJaG>2;PB3)>d##JV9a\U6171_
WeL3c&SF?1>Y@P36&N/I9]MMQK>C08cfAeWVKMKJ[7Y3WeOL=.&&P?]70,[P1)0(
T_cL#beBcE:WX=W4cScTO2JHFDY#;-I6M;.JaR(FHb\\PLF?:f31>\(86[@1^84F
8DE2&CgfD?<QG3?0c+42WXP+d^]+-5.#=,KVO<GL+)3,>U<T?EbX60Mec=+NE^ZL
FfBGM/N8D6Yb34LcXJNWeebcJCTg^+2)<FHgWU6?^U[)HLFI1Y]J9g;A)QG>W4TO
bWc-B83C1X069eI\#^A)EcZ0_OM2D>N^?SC_.U6GQc)..Ue,W&-T>@K3UOM?VR,K
g2fP)f\DW<=(W2RM8KLMON:#/^+bG:c/ea0XZKRCZY@TY,ec2S49X;#2TeKW_D0B
HRDd2FGWaH[SH0b]+O=8W/XEN6C17cHN?QJO4=QUZWO/JC:G\ETZcM5A.c=7BMbK
4I6:DI(2U]Z)CT?+UDP,T-[)BD\SUG2>YS=4K:a1\\->AAgC/LR4:JDAKQO\,2R/
+/^D2c5]@K/TC:1MU4[E7KBgJV-TETK[g+gdD/[a\/fe3.RYHO;):G5Z6?R@Oa=e
.aaB7g,CU.]HK]Db8<Yg2I8Xd@8H2DDCEgBGa4dSg66R9>P]<2]8Dc_/9GS\d)BI
NLT(XA#E-0@64M?>&3],XDO[>2c;P\&>^-7:\,6-97^,#W)9C3JOK\=c9)B;c_\O
W3FO98P(9PI@RE5=)3/^5d0JOAL.A4YO6e_ZMg?A/c8\EEa?(M4dK:fJ^8WH_YA#
U>cK0FC(IKI?^0O6#<=eL@^E\.F;/Fd(@:<<f;@QEA^](MB#,TU+CNKB]f44NW@K
)-ZdEC-8SB31UC_(^7c4@6+K1)W_ZPDe9e16<7&YZ=VaDR2DW>&LYYdb-DC4.X3R
Rf_R9ONQbNHNA)776JAWHG]d1.]f9/523O0HP4c9Q_O.[gWOS,PA_DY[J7HOGC3;
GN9NZHYOS5]2gcE(KANBM/BW<f301b>K-CNN-8F@1BcN+SFVN5gFfaB5HRYfgR(c
05[[<>cZZTB/YX&HX?--]\6f>-XXUaMCJCg6WWG[OP)SCfG56QKNZ3O-\DB=bcfH
CF@A0Q<,U]\TVAS)B[,:^P36];#B+.S3J?D(Z1BULP?KES)[&.N+HDAT]bF9\Uf<
@;VA[O8dI8>U^e1<VB/Lb7\a\T3\)(Y.:9L<Aa=UB;H^^5dV2HZTKN)3N4USRC4d
<YCLY8I5C4S9]J4]GN#+f5:IT.&b]HI;BbdT_+-DYJ2gJBQF-DFHa@6SJIU,B_<2
Y2<TW5<7WC)LK]U3Rcf]4RXQ>ILDAWbAOVPbLF=bgK(c1?HQP<UY,6TR[\#D/H03
Dg-T)?-.VO/bC/ae#:\:U.OeQ396MPg2]+.X]Z_&4Gd+#a@PHKL,U>IM?Ia,?<[Q
>V@DSKdN=#Q#G)9O?XeRYDCYYU^9X(b90eA2UB]6V6G_]]&?GT-(R4]7O&5ORHL6
b=de]VPdLJ[&Rd[0OfgR56WUD55W\d^9PN97V;<;T]FJ<Ke,NGGaG=2_8fDH3/M-
GdV@=8#2-WGFPJ7ZK<GXY:=a=5JV[0J?93//PB:]Q1PZ5G6ge(12>\8.R;<)<&7N
,?/,0SQZHgU)^++S#755GD?I3CV5cVSXXMQS\<Fg86#PX8)cEWX53f558dXCG(c/
Tf<0A6,g:&MAE/U4E9HJQ5c?3B<c()_OR?[DCZ<S<P^eVg.OBd_9@<YaCgeSU,(I
bAFXc1bf,T>#O0Mc>a02V(AC5<&\5Oc531XE6eG1=X?/f6TBL;4.8TVcH<DI;;W=
VU^<aH(&aYJ1Z_3J7]eJSC^L-S7]XX<D[C<:=.AYTK)Udc8GbF;EGF?OE,NXbK;X
/RVUO5ZcNLT@ER_>7ENW@R.H:OO9]XecKMH08)FR/LQ4]W91FabNcDC@,\d\:)J&
>A;e/7^(IQ<8eGS)_Y2F<7\B#84+5(F^9e]QV^eF5YY7(^=&@45SR]SLLN+3f7L<
N9:FWeMdDN[:#E9@3URb/.H@X>#^\V3XU_]\9]Q[S&5XeXKWYO+6I)fKIVJMJ&7#
9H/^?@:eZMNDBVMaY?Ia;[N&-\1BcB19[?/Hf^LK[SPY\BU-X+EbeGTD>OOIUL#3
:W691J724C8@AA@-c(XZ+Y_c5/#N,Nb>^abeU2H&dG#;^:3Z)JB.-N=Ic#FFc)1?
g8T5G6@XL8.3@I]d,4GO2M;RKU<D].O3X0@#J)-N_Y3)A1:TS_)(I9BJ4<)b#N@.
S03Ze,N2H5-^-/P_:[.MSBQ&EQS;+7Kab,0UAa)YY9),dDc([a+,g[.\^#d:Z3)W
GD/[\(BS,<G.\=/N9ISU?2RMAA282H9YSNa/#cH/VODFAaVSL5c#NdMQEVeN#.PG
]?Dd0[LFMIDe[P?;I,V138O5OUHYFJ-_HO21V0]MYJeFVZ[4Mf(UaM43J,G@)^<3
#bA:Y7g3.f<6PL8VMc(/]9(g_.g2LUME?PPb#)S;1c,1fF+Z3c[=0+RVNLEKP:AJ
RD?185S\Y8OL/39DR8KL>--2P.@dCWU46^A:?b1ENg==7_]VJP^6=L;F6aJ\&:8L
a1&G(7g1]@c1P#BU,_>aa2R,Lc(;+DfO(d=3WY0fJ/4#]SgX0X6OAa2(>&Q5G-W<
<9.c+#X9JcPDDMR?W4W&cR5J#581[W4P@GXGML-ZgLaSZ5XfI/>]N7@2(_/.+#M>
N^PgSW<gS#ST:9>^3;<Y\-K[O5P+<9.P\4XO9WM0^7g^MU08FS=TJ6C>P@DPF]_)
cbOV;)\)7cDGAD-Gc;8(?\;(V:]5+BCcU0=H&[5H5VZZ4.CY+><:-<:gNXCZSb;a
gMHg-H[9)1P6EI2@9C;/4W4RX8@G_7gZb<T);&^M&L#9g\BFdFXFPB.,@,BGHP)J
SZP&0,9374WN?XH=P2720.c]1cB9SA\&<,\#P^XD:<B>8#FQQ?UG1dBLPdGC9+5:
g7F7a56_E46E4UV)agX[C?QZVQ5OU;H6A82^)F:@F]J[>082-Tba9?L<A4@,(4c_
+P<3485Q1])83aVB2.TU^b4UKPWbB2XaAI);^AW-O/d48#A\[ee(YaGb8;WC-7Z7
643@=f:A_^23EKO(e+b;_WM;)YWOGdW#IESegdL4SC@-AC_74[5:VOIW7)DE;(8X
eD\K/f,>80Z^QMJAAcF(>=<@]f8YH6IOdZK\gSBQB&QL62X\^AH-Q>E^[P)Ob1,H
BXH?B.;JDf4CK=@#0N[6BRH^/a^a[\U+@Yf+F(Y>c[_/&LL\/5LZW^[HccCV6aW3
Hfg1B0;+&^FEMJC29H.7I[L5BUUG?dCJXWWa62[519_N^]2;2\AP0Q09@C<_]Z=?
;L24[_V&#U^Z-Y@>81c;I6eYUV@R2f>ZW5C5JeW1IL=AL&R=\UXJJ\FLZKW#Qg;=
XJ^/GNP#\e#WM^P++.#A31X<6<Z6NgEJ236f00QIQ=6)0;eSG/3J7c]d):865OQ,
=J>(V99_FWDGVcdNA(b&;EP;H[E-7)V8J(<Da@.1M9GY^S)[PQR7HZSS4+.,Z6dc
/ZcK-0\aE7WKR?=NJEABQR])]?/d;Wa[;64;B7bG>)8.9>.dcL>P],KI7K&8J30)
+.HI9T&.T/:B@1:+XC-6.NZ(/aeAgS4W#:WIS&0,MHC@Pg#_,\0R3A8=NQJH97d=
C>^4XA0VT1bagfNF71HYUEV4&G29^4]fKDfd_N#^7FOGYd,9QKeWa:DaFAWTB//e
C_MDRXP#F>X<TW6#=(\<)?g7:745L0VMP69Pa7Y2-]dYDagE>Ff880##?4>(O\/7
1>7.f-]LeOUc>P:+I[[?G4cB\HH+6(5?2fU<bK&JaAHba[M,^E)bU^/G7BGL_(GH
SW[OV2D>^N-NDN]VfDGZaMcV2^:,,Q(B/:H4R1L(O7A3J/WDN_8#?O<KG59Z6f?L
H4a2[Ug7197;M]?A]7VC..DZ1MBQUZPN;DIH7I6OW7W-@HNLE@#^:@HLJ8CD=S>=
R.]?5-J3@M\S\.B^J#bZ=DSE@<H4e79+UZd[QHN:=U@5.8>;:T>W_FC97T_7a8RR
4QOdT&WgKU]=N=Cd-A]8=GQ@0W?DDC?)Q0KNX;^F:PL.>T[+356H_f]b^?gAQ7):
?I6&9e[b6&cLUdY9N+>/X([VGI&.N1H7(RP]JV)I\K#71f,c:(S.V#;M8a&J\Z4_
M&_A9?S<F(X2@f^_R&Q?2M?)5>?:gK7Lad0#)FR^2H#]N,13T(7XQT;bE(c2g=7I
fYHc6TP&/dWKI4OZ2F2BO]9aP26-I/\KTAT?-+OP7aI1RD3O)MEYN\2,QDS0FWM4
B:FB3E1a5)^TLI#3fd+-aOW<1c369FCJHGR/Z-D-:[(BK>+7K<=QR2E0?>DQQF@3
[^4(ZU-RL3GaCId7]@N/g)Wg)5g90U^?TN9P4Sf4.6Q2LI2-BeAT8PNJ1c5dMK6\
G_0RBR;dg@bZSeMLO4D93>]0Z8S]#bB4+Q^5TaZAT#V)RQfN>VV);ga;eNZWcgde
15]C+P:]?I\:)Yg.a/.0]4-0Z4V2W?14<+BSf\XQI9)\?D@bFOEc@]E0#KRLWbW=
C&(f2NI,-V/+13S9T2UKQfg&gYH>(\?5.2QIdY5=>dB>W.9CH[X2H(Nef=#8ae4O
;+Og1S4(Zb[7X&FI;]G(.0HSE<IX/_&+64Y][QGE/dZP+NAR\[88X^E287?e=e&\
_M>/CZ\5g=ZVR?&FP\[0<+N@52e?<[2&PSEXG9F,#dBa??K>V,SKaW5bb9d_AQYA
P>4T?)_VHT50UfYQKI)WXDFCPJ@7THb(_eW5aO9X2^4-BK]U4V,77CU1Z&d@<_/=
MZJb6,=6?8C.UY+/ZAGSQ#@.Z[W[L3#\#M0=A/,IgPL6,G,0[O__E)+4fGgF3c\f
IKM@+X2+f0G:MU/Z)?PX/;27<f9#C-K-Y^)?X:@4^/1<.N]e9gR-H816FSI0LFf1
WZ:X2dTW&#H7VgWYVcPJgC:Gd3@C8+B#08GIc4dgU5K_6OF\?N-GHe+WgY.T-K\g
cZFA5fHFLGH1_T9+4)UJ?K3=G>:T5.]a7EW[Z-62.;C=:;578#O6VX:d[PIQ6UcO
GaSPPe.aQ1+[E<ebZ/40G#JVP]YTFJL0Oef=gBQ9c5O)?G0:9.QE[+DG6G)ebQOf
Bf0V4F?;abL;F4,(9g[+aF7]LHE.^6LS7P:P,:g[E5Ad,8Q&BJaUD,QY:V2X#)&8
&(]Rc,[>G>6<Sa2.1Q=@I?HN2f.@HE/ScIaFPU-YD@>C>SKK(Qe:L1?e&K66.(^/
6LI]+XOWS_:dc3>ebYVe)@9WEEID5A9M.cXaFDG9OW^&57@I+d;WX4.YEY2HGV9W
:5+Ya\=+2YU?^A=+(GX)5,d&D_^8?05KU,FHJ1\WfYIP0Odg=F_;a,#\Og9?]O;4
B_T[V@D7;8:^fc7CYHG:RTO;E=0X[TKGJcf,\:X#>GA9fNMM#<KATa_?3\cTc+JG
3EcaVg,]Ia4bK48.g:>E6XR+1P,RCGP)-<3@9cDQZb,KcOC<6cWd]g\_C[PZf,,7
4Ma#0\g.\Xb@[J6N(D?J)7/0:98D+QEO@(DdQHBU,)V?[8>;_JF.94O^^[L932e+
gg&C9LGJf3/HY4<BP9UVJD9I)(,=&.1/IcQ)H#?PaB.1_\eT-&-IPNK2D.AQ:NFR
[2:=)XJ\DQ0TXI;\9^:K.+2P:afZRY=&;.0Z@#K:3#V4^</<CEK61DT#b,M3KN=(
ITVRR?OX=DAZFN57&E0cK2fCb9HR6:6YI0?7EVF2@;54^X4(eBO4,B)aW>V4JK0J
\).S8^;JUS+,G&L;T,G/dDW&G8[&H]gS\\B88c9,DBOfQcFQG3L:gS.7>V(LR11)
<E;cGFf^XEKN02^:/924cY_4EAIE7CFKS+?C;5S2QON[SU^Z3E\HB;g8F=M.X[T_
NXD4ZVRf=537/+A<^V2PQFI-/b7XVS;L[<E,+.EFAPH,<(_?MJ3Ud>>&fE,_9^c^
&Y,_FAI.B-R]IfS,F-^5eB;:3??9IIIBe4Ib\&1W2_LQ@8.B1:M3=?U#3=8a\S-[
4:/ae^)g-f54&9OQ=6N1F(e9Xd0S?,QR0QG@:)gNB+6:B>;Wa_^^1)SW_D@01F@_
]a6#X\QcgCa&+NVX]H>R+1:[MV7U1[?&5?U\=5VeY_cYcV6b0ISYA[?C5:\&<-\_
0KM;3ZY6S62[1=g>c/5UI<I9:D\.Da/K3_4FRP22GET(6?1JT<GI:O:2OVO[(=NN
A/C(-H/.PF3QCKeZ8J<N+(EL>XYIABC?,I^G-8GCP/]R.Y+-^0b00<D&1TQYYYX8
fO_3JHY]8F1L-#,,WNC_QCdQN]^E-LMCP)75M5UB9cU>G/V)=;(U#Z]8..1eK;X8
d81+X<Q-3<[a-K.-U-g>:f=>3LQK8\7&ML/54W2CNSM+a>YQ3:PSE7]C\I.T30g(
cH?F6FX4Q_GS^,V18?-.RA?d_GNT5QAOE[X3<Q:MPbQ>C06)MF2=fR(/?V0Z2a07
C]#BcPA1_;2MRgHN;LY;/<bHH@LfL3813\_JaF#f<+aSXMS-,YAc\GMN<TIE-Hc5
4b(I./W[9OZ39;O(/.O5(aR7<U[^HR5]#S_Q23/?3Q6FDCaI2GdI0#R1?E@1_TNX
A:8_1Q+fQ\Wc1>#He)_\@0GNSUP#SF+4-@REL,/OOR6Q+N/a;;MJaXAW_N-28d^=
TM-0g5YX2d,P\S\._TQ#1:)d]Hb99#2SZCADe#VATb@6XH+2g+Uge-^5dN\EA\MX
C>9S,PY7P=5bDQ1^#VLWQLee:L94=YQU_6ND\ENg?U#CS>MZ^7f_SWDT^TKTO686
g:4.\T[<CP=bTQQS?N^f-?D+.4ANTD7ONf+FE-Q?6/KWBN](Fab&]PR_e8g)3Ub4
+MHa58QYM?Y>JH>,5^KVN059BgC@#Y5-fS5TXT.aQ8:\Z>,a#)4Wg_cBUIDPVCKe
V(X\,,ed5D;W&5M9^1F5XLRY84KY:<A-,^+>.LgC1:]f0Bb5GOgFgS?XUe096]T2
9X7US.<T3T0)+g.[,W.7ZQLCg[W>9;6,;2K6.UG8b,WZE5Y;V(E6F^W:YSJ;OW]<
_KNKd^FII1]bJIV8+IP8HGR0??EWDBe1/4?9@HC]IaA=SX49[#5GC)],=fF^WQAD
^WU5>A9@1^8V5A^-@ZXE3R:E2YVP-\eee+=Q;J:/(UaKQeL_XYO#804B@TI_(eJ#
MQHMPR\CY6EDNH)1eG1>H#GG4@>&:MH1Y[F)0FIH5J[4M=7A.]OTY<I(L_&TUfg4
O)e3;:V,.8(CS1&I&?IB+&YE,b(W8<X8,-7OMZ^X=BM44-6M73?NdD,VV&S+:\I2
YO&:e8&c&NB=FXgaYc:P14/LA=b4ZM8]HG#VS04;6]-EA[<XS6C].gFdId)[D[-[
,NWPW\^@)&Yec2Z82d_-RBB(@E<\T410<1HN/N(.^f(Yf]&MZ:a(YaS1)+9_XLLB
.-A[Z3Yec2DNK<>/K3GDE+.ffGZ]5:dQf5.M<SRZ_/.S2L.ZQCg&OO9(\:b>P[#0
<Y(CAM-1Q<8^ReP5NHgTbP56U.3+bKZ0J3b_&E:KWg5FJPDUXZH81a5CHB?Kc/U3
b)a:I#g35&<A(cV&)d4_)AVM+\aa#PR4a74f+VUc8=)J:cc=U;CCWV=3&H6=)8e7
=TZ]g@#(U]0&8>Lggf?PcggXHcUHUHe-]g#^@7WK4;<0_RQ<XbGM1^HI;f9HNaf/
Z,4f(K0K-dS[O2N?^25WC<ga_?1:[e^,IAE+GAg(7CL?]Fa2(H(f&&A<TE1X8U:/
NK,f/Qb9^#6I-KDgIf9Cf/,3U3e=da6A(.(a:g-[&GZEK;f8<1(Q^-Y>7U0G3Q:W
_SQ&W&YZ16&P.^_]Gd4>=\,YQU;^>LDSRe2NWcR36KP=COP=>7)O8Cf_Q&Sf<PaM
b#gW]-\7EO50X8HaI&<5<UVd@G(eG+YS(7-F]#+e?NXV>H\;GFQgSH?Q:[A<=6&8
I)@F\FX);1-/QKJJH_dK(.d1dQY_R3^AXGJK0[R)J?P7-.85c6^6N3TcCd/DaUPJ
GB@MS)2/;gOK3]O4?Pbe)Y2E@I;[0\;]>X=0dG:##^ga@IZ?Zg6dHaSV5Q^V/?1M
[c@975f)=[7ScV/beQ6KR>+a0?,OTZT7G5L(g@0M77A/:05ZH02[61BO-S8)ZL56
3;Fd3-;2J/@20T^?O_@E_2cA;LNIU8FeM#MXSUT;PA/1@MaL>gf/TB6X+:T^ER,3
Q];J7PW,eV5@+GRQGd0;\#826)Xf,P:]F^dSZK[D5:T77gcB\G)&DAYYQd=K[A]a
/-:))=8.+PJ(]TL3Be[D;=eb1&E(#Q35S<3AEVc?VA;]>HC,IVNCYXS[V+Y<.1BB
5IgSYGE&?VT0Bf8656@)4ZD]G<46S<LebLW7CO&+ZS@]UPB4O/c6e)J8VZE2OgV=
H9F#@LYXEE,<F&=CEWeEOT;H9/4@W9>?.MWM8JEBW^<P.fc[.D7CWe=Cg/c&S6:S
HQO@?aHE(1&<?gcZ__Y=Y79K=d&02_@VXG)6V-VfXce]W<P;Ed8+e,Z@&UcS3+M[
;)F-PgNTe5?_3SK#(.S)TLXcR\.1F>b7;-O)]D,d].5@36AV7K-K9c@fBAPf^4N:
bMKV/Eb2cQ20Q1O(45+52Q(ecSN[/afa&>XIZ7R>+OZ&##_1+P(R@HO/ELN5QJ+R
e-MBRE7](S_OPKVCUG>;5>2H93Z)0N-\BKeT[CTP1E6+#:f.W#CW8\F5:47E1GKV
<g-bA4^^R6f0b1F5fNWI>Gc1<MG/ZE<2cN,U<8AbCK(QEW=RL59@7.\X=)QP_JG?
D@DC8AC8F(HO]ZWDO^X4^Ld8]<,a&W&N5VKA?V=E9E.]?8ZFI=2BMJ9F_46[/[)I
IVa]8bNWO8D;P_A-EB3M7#OD7HGG6]>R[\acWTZL0LE8ER@[7U0&Y:2Wd+,\\b+^
0X0YR)Tc;F#RL<+c7X5Q38FEKS:4aKX9-&0Sg[KI/@A8Z\c)Bg2K778NZ]Cff.WY
f=1.?AE5K^[4XM??b#GQfM,ZRST(S<bFE^F9A7&/LX7a^+V6c9GYf/ePQQVfQYTf
.,<&4@a4aW)deE=gUR[>>><9/NHM\U^52>>.C]]<-WHSe@<;Z[F9Q@;=<K_OAcWJ
M^XO5+9HRRK\f@408e,,C>B;?ROC-EW+?6e57/0gPUB:L2I[6M?-d;_CO:a&_S[V
A,&^P\JCgF7#c+W-f.A2.LD>F)NI3Y[S^Eb1,0&E4Xb@,>3Z3eb/E7fMbeeK]_)e
[\F@<KV[JF/RAUb.>0]_HAOH,Da[GB_c)];b3P523^IY[/<@#]1\g0A]0]2VXe8#
#R<SJEKZXR&XU<\N8S1E,+g]PFaTJgNZSDEWM@f_=M.4bGEZc/]T3#W.\K2fMZJ7
B?DcG_@+X@W7ROOYT.E:[Z(6OO@^I+T4=#B<\61QKXU:3&Vc.CGe981BDfD-]ASU
3\XE0:VDcEGO?<H2C>(R2dZ?_7A;<+=AB:Og=1PZ5PCNb93;f70373JP<K1,TeOX
,>]b5.C--P?ae#5f1^g]WR)T[C]&P(AO>\/]9;7IM=UUMJ#G64GLBOI&T4E))3[C
.YCD9DM/^(@4P0HI]7]fF,.GSAc44QHAZ4+4QU#@T\5-0>NF=JE&f,Z+&bF92Z3V
E;A6K&b&=R1?FFYc5gB]1&,LYV.W-OTeS1-6.;R9F+AfPQTAUdNgMX=,=O+31dF8
\TMQ(L?N@RK=I?d<eZPS5A5P9ZJ,P(&EWB:3CcZ?@VOL)(WY\2+CA1e@WGZ]2H]Q
B(@VgMS0_QaT6\gR(I)KWW)Ve=TM8^K&/@^M=>/5\(WNgW,;,:JD6&46H>A^S#6[
+2S-=&BE)=TZWYDPS8A,ccG;Tb\;b)2XD9&gEL?aE7FGZ>T)fW[.1.8efdBbM?7,
:JJ^R1(RC/g]C<8VJ/ed?27L1,Zc;<8T[6P)[bG/8KD6&QM25B>-K&OU478L;AL8
HaJ<eV+-.8F&H5L.A#MLMYTVd](DU<6\/NGCX,IX^1<9BLF/VP<T.-XDELQfdOM0
ENc,?3RFK,<+#34&6K.-QHERZ1QBdGNf&BN62>@0?8-GL#T?eX_5Z.AU]8M1bTKS
-WD2)7:>gK?KH6cMS/L;=LZ23:J8H.FSX7R/W-(^NE3e[W+eX?+QUA=fMFeGKK&?
[6ZLXH>9dd5c5NP[^0JeYSEdJ=W>IU9EWNZBF[?5bd11VGZ<F8U04?&RYU/bbXMK
_3bNY(Q\P#Q_Z+)2M6QJPV2aQZF)/#5G3d1YAOc^E(_[AXaXESJ4S[09fd_Fb<?0
,,C:@BCJ]^.C/[YM[4O:]9&A,V7R5D7[T?dX.>HgY#X1K\IFZg(SHPYG_9VHB<]_
R<9Y2P2GF3B^d]T7X:\-(#J1ASVO=ZX&INSYYV;BAN:<\&W==LdJ9D]XD>KMW:Q8
Md:,-_ca1\[OY3dC)g-R&a9_.D4:a^Q?R\[9\X7<L_1+_c+N4RWVY&<@728@_?:&
edL#\BZUfcc5W24Y:61/^Q\C7e#SNL.?--UCR;9F^<DK<eE4,UcKG,(Z#INH-6,8
?f6gQ;AW,A>a/;R-XLB1U:8=>fgT8]c9?F]66c\E-4IC^J#880=\L1T(ZXBFR0HC
_+;\bF:PXV3E6e7EEIM3F.6)+H6BB@8TA3bIf/I:ZH[GB;,M??g)S.T(TeC\MdAQ
Ya/[R[gWQc^YDO/=ERg2,d32):\R0T2G?^LBNFQ;(ae]I\JQ)c(:;U.\MX_Kc<3+
:IAb=cB)7+93+#eWJ8gR;\,Gd7GgAQ;&A=b#\DZKe+HOaT-a-F92QD.&&]V+Aa-@
gd5_4a@IV;aUQH;,a\bd/2NaI>HMeQO,UPTgNbN7Z>-A,PF,WJ-V:E._?R2e,c_:
Sg]N1f9eNcUWL)d<Q\EM(\8eK+FB(]_;T=/LM@ccEN]9VB6]<24LgDDIOAUgT.2Q
R(69XZV&\WM2X-@]DO]\->.T0-d^K:#K8IJ/Ha2F(8Lb6.PK,cG2C+H6;Ec>-8)2
gQ+9)\1aB#Q8,fP,eE,f]N5GUQZ[[U_W>ed@VN6,66:]YDSKeX6QFc/)WX4I>WCP
5EaD?Fe8Fc[,;7Sd8;cK8,@UG6Wa(=1),4ZfN6f^&Y7gbg#d.JO2U.RQN)UKE#;>
>K\P:DS4?_8:S+-)3SWXA[b>V3SR\/c^)I9Xa-^L4H13ON(;0fgM@E^G+eU&:Pg.
4\e4_D-[+B3AOL/E46>=VT)G(2E/=d7U_f?XGJD6R4_I#;5^2fC-&5_K0Q,LWSTf
>SPHM/:f>^&A4JBT>XfR)=]E[]Q5GBeH5G:+>=(GU/K(c>dQG-2NC/E^4FN\b[e,
3EbW1V3J&e_YK)Ef?ad-]>>QDKB>_e<..#BYOc-eWD;B;eRB\6?I?Xf^X(NO4EKW
@.OVGJg#b-f<CV2U;/((gcDID-1_NBKeJPPbCGF[-ZM_;7\1XSE9CLVMbD]YFP&@
b]b0];:DS[VBM&T4<WL\;bP[C7EGM8)XSUDS+?C;7SKZC8BYdSD942GNcN@JLNb@
#XMDB><1bN[DREKKP-M]V;cA(S2;OLK2K+@-Z;=520JeAJU9<9c?,K,0V3V6;216
#4Z\CI-21?E0WZF00FgRUE&G_+X/)a6ZN4M]6XZ=eHCA:J2)/QY?(KX=N#d#bER9
bK]<VUbU>F+WU)A83L.]\C5A8-9T?+0]?<^@_RE9gYTfBQIdQ?L4TffSD30dR-M5
(]:ZO4F.>.2[S21NNY=ZNPGIY^KcDAQ^R?0(62;UIa)&H[5TgSMa02gU+XJdYG#\
J40AM#U]OWTN2VZJ,]a/8@RF>>IDC@VW072ag(8J#D7XORX,.<Xb9XZNPae0_[P7
(J?SZA36FP(F<DJ1ZQ>#OfVBXBKK(^YM_@J.J6aNF[4?L7PP3G<YObE77@g@IS58
X=<aePLZ@S#_1\XgV+TE6=[ZW;<-Y5/-g2R/bD254@,4;]JLMH[SM:1?<d:)H\Yf
K,g&B,I:^L+<T2JR\E_]S\&1UP^eK+cEdEPaGIUZ@^3P_M?/IXU),8,J22XS75C3
&VC9?]JL)[@U+Q\D;&/?/@aW&2:Vc4B/WBWZc[O\PTZZf+(7eRDL5O<<M[F/596L
ZJd@O\FY,@Z)4-GQ?W>/K-#Bfa=Q6c+>J(O9Da<6&K,^W_5ITC781+b\4;/)(5Ne
SEX^a6c.:?WTH]ac]K)RFPc@+\]HC3gCO<B/032I?^T[Kgf[gJVF?(ZH#B=(Bb&g
O_P=2?9J77>:>]8(UNPDcTBN:Ba0WOFT49F)F0=+<(KgV0-0aHAa=TfNX^O=IE2]
+;C:DLRcbWR5^MCO(aWWY1D3?_;//.U\LXG/.R)1,cW[gecZL@&7aEOO],AKKU^O
b32@b-@CGD.4NDebU=T6MEO<?)K:H#52UCBAH4R8N=PLW_,&=O<C<3aA2&9O^WO-
)44.^NZ7YQ/N.PD2f/>Tb3;SCL^b5ES<g69#CX6a+:Tdd,gZD(\b7M#_C/-NIB)7
\^N(^_KJG(VU95YNQQDg,^;b(@=.c-BQ2C8T9<#;+VFV=\/O^]PfSUFDOQ;G855)
da]7cFJ_Hf+3KYKb/V;+A=DPOUdc4,gb\A+^9_7,,(,GOba9=;Jab,Tg>B]cLZ3<
&][L8#cacOSb<6H=3G,aA0f_[7bg7C\aUH)?&B(--&.)SNJ]-OI4^5#3PTYIe.#J
Z6F=a0(JHe\Z_B.:/225F8)P.99<_X&9>E1D^+<fF:3KdP[a(-7J-5fG\b@VK9[0
7)<_XC=OagSZ6;(\@7LPDU#=3(;0#J>FOP,=<dTOb.OPfGZfVK,@IB[^J5K4HFZ6
RQc@EU<^D0>Tc</R\&T=6>N\:5_7PPGN&Q>IY^RP<ReSV9HLJJIbcQGK__?ARB@H
Aa-<,/0TM+NN8+S\3e3Z+062A6eBT]2RS/5]CJ)GECIP3X?2N&IeP?B^^2E8W]Pg
AJ<<SKR9YC9CGF0&<3M@gV;70.@1U/2&E.]Y]9BW2MDdL;4W[.+K\IUJKDF-+.4W
BQGQ(O1ZBaLOI=5R15Sef/aTYM>285BWJQQ_MJDC7;QBRe5?V-\+/bNUWVAYF^P/
KI)+VJLd5D;f^DKR+PPP1ba_DRe&T;S;<TbV+X9Y4Z[\X.<,;/McAYZCIgKGBgGd
FOd,La[<<.bg32AYE;>M4]M>9H_f55YILe<TU@CTaa2585B<dV++YTG\)8WZ]U;6
b63\d\NR,Y-DT(M;U30-@)gT.2YP7aE>YgZI)DJ@@]cgT#2VA2PMJ4<S=gZf&21A
FX^NX0aNBN,,;eW-/ZO7WWU,3<##cQQHH6HE6DcTI==ECR?cg00#\MbQ1M//TLfO
e6[UVdR#:.B8Tg;E6LJ&YDWIY1#cI7@M\,=PIc3P0.+X4I\^VVYI.\S?WUY(PQ>)
=U2OT,+DEK2X[1@SPI5Ub>_aP.aB\@@3H#0dWQg/cX@O5J:UK-dTV/D&X]\<,YUY
4RK]^:?9;3(X:26f69W/,^BJ#)?Ad-.]6&L7LXc2P-,X+Ha^=IdeEbLgX-c5<8OM
50,HF7?LZfI+A0B27>68HQ2gfWfFN7/E.G0(a\T@f.AZ&41/8B?Rd5P<:,>HQ<HA
c:0>a)O&K9KU;9U:./_SO8&Y.5)2WT?#PV3HdA\@e;00;>2=5C/RXJVAdT#VMRf2
_^\TG\1,G_6181)N57N1?UH6J/U/7JWJ/>D6FZV8:cF@VfT>XMBc87?0UIXT-O2S
\AXVg07@#N-XIAT7MR9&1N2AC65^0LfXZU/C=P,P89OO+aF3X_4582Ga@BU@75e3
F+MT6&P/PVB2#X2G6MY/g/^LR7]+c=C4EV]2K4B78W0?0L&LQN/BF:>B1.;,bc+\
Q@Yfed\(6E;c06O]39@@JKVc2aEJP(6f8g0Q7IO4.OI@(:Bg@N2H06Q)NFcY:42X
T1PU7W6+6?=6FWIcBPL#>FE][\KdH&[L.a+c+;RZX]K@JO3NHV?>dRSLgPJPW4VI
g2a9HDEV9)\._Ff,TVN0>:c#57I=9#d7.;\UUf)).\D5/(U>79&3-@X_B[N61C<,
>aH4;DCc/6]=GLDc[f:;,SFHT&X^<^<63bB_UOUe3J;R7aIH/CPbg7Y4e/9eg=+#
0HU4M?1Z)?VEEBRC3.R\#/TI-^2caZ.XN_fV.X7^,5g74g^9(([GIAVJ)P:0P\#f
P&;[(8d#6dQBP+L#B^+Fd?ZQccOLc+^75<>0Z?@)<.La76B,cUF5R)F-<C3c\BS<
]/;dOT39T=YZS\(O-=?(QZFRGI?;?#/GgF/)U#539+I7)9PcYgJR5eEP5<X)X8X-
-CF5U\;1a,(S1[=6de<CCAd4NCLW;@S/NPS4bAD/XGJDRI@\cZ]Eg7aYL>ZXQG.E
<&CNgDT,Lg9TPg9d2=3MUa125DE_d8D3UT1b@:+F73VD0YfZ4aIG^M8]MW<E2YV5
.a:M]AUYWC4_OaB6bC3V7GPFI6T9/f7gcdcU?7Y?E0\d&WBeA?8fAfM3.V9:Z5Z(
EBfG3TGTF8?_QC#@O03=IC5,FBS3[TJF;(e1R+1&:>C(:\I;+ZK<]bWT6(7a##J1
+=:6e3:O@7NJI#LIHR1fDfXN#D2#D4CcTXW/\b2_)5fg6U)(_)-7/5>d\4bNA4YF
Y\B=G/)_>)9T/Q-;I+f#Y>^N2DB(.U2&]@0F14V_bQ;KZC@d_ZHED@_:G>96=:3,
#;M]+>f:8:G^9;=KJ8NIPVNG\]B.](ac\b-]S4#-#/BFW660;SU,8aCb7ZaH4G3Z
57NM,Y>Ne69V/LV_/gIX/4dI]FJ]Z+:HZE1XA\S>N./0;#+X.,A\YA;eJbLXZX:J
,T2QN?S#R(FL[\e@B5V/^VRKe;1[=\#Ub.>#,?HNa>KaZXbEY9ZS6Y,geWdFJXWK
4F>7fR,L?G/)g:&F]^ZB/\OP3E;>BQ(UM]D([5:7TYUYAFU:C6CT#dGaO_dY01,Z
()C^1a#^7U/e)/<^&DVN+WAV>5M03?&aJ<WU\2J]]ESC=3P_e:U.bX.X:,W<:;V9
<-6Ge1TcT)DYH-2S/JCY07#:&TAF,R,C;NI5acOE]1=dN8^:AW;,/XTT\7BUe?2K
S9B)H=eYR:PMK+[L5S.1C]Fd=/=[Ba0QYMX?3<EFQ_b.2CMdK,Z1[/c7ECf&)FbN
=RT3^VE^c#IDaE>cH343GCgMPb-f/7ZXV8bXS+S\cR@_Q5bTJMO+Y^Le_Mfb7[b-
d.#eb0Gad>V:Ge1c8J>BgB2RYKcT@9^DQ,eQR=JYf-J^g1M&d5SCaV(TfOA8-Z1d
TQ[E>Zb,FXQ.00+1S93b>F:K_LgfH;GgR/@T8B.G(7/R9U9JG(B]+SWG5C6S3TY/
C;P@H6AbO.dNR2MN]3d4OPJDScNPNX(f5EJ@97]]0(QJeVQSLLS:[9-^MH(6F8+E
=)REVIHXGWE]1[CB_ee\?;f9G9#S_;E=&N(P;2/ffgV)e_O(<=Ab#1/B1T?B+\((
dR)8;gdcPX9Qd7C;g)#-\f<@9RLa@IBKHZ&X-1_F^Xf#@S[]_3#?gF;X+bAdXRU6
/^D14F6+0g&[g7NDTW-53&cc4:Kf@3L;[/BEf64)C^;UZ2)PbIM84V0M=fNbKD6N
R.78Y,AZ)G\/4DLP+WP-.4/]>J2.<_AfJ762LfV-eE7g/;43[09R(2JQ+Le&\-KH
>&)V&ECA5MIg]^.gZ.ZU^W^C\;YX^>M@S;b>^C[,17A:7VMVC>@++[9Fg^c8188#
&_-)PH(3]bGO=[1,23R7G,JSR,UR^:N[b^NSF-eOJdK0=FfA:B2FXV?C\]?G_OL]
d8JSW_N8CU4.D-;,?)LHC5MVb@#=_<_G5<a+OXPEM_T9bHEQ,66IQZBB1>A=L)DJ
Q7?#\5-8f.0JI6WBBC0_G6YHd(DVgE\+NT,G_9)?K5DR@K64PEfcJYcG6aWQR8W,
)f32SWSE1^e5.RVA4+]DE-K8/C4];V0PU7dc>Rb+bSDRMR/[([42IbDX5T<f)+O2
bN@-](6]GDIcZFWg8gOgV)-N>&bY>8)7fR:Wd77<B:BT,J7;O@,J]>YZE<8gVM:/
B;ZYVNSZLeXQEGE:3B8PCAgQPdc?68;\_YA]IfNBZTdR^4Xd&5c-YXeR)D/VBHZ/
7c1_05aPf5)bbOXeO99;G^5gK#ZB\e,)^RLAL_)/3.N1VL@+>:I+-?ACQf;9IcgF
=UI:5B9F)#\,:QIE,b1AR5&_<RF6gY73M#RTV#3c[?J].a3M^+e>LCTc3]Ta@)Zd
^V1XD=K9cJ2A4(,Nb6VDC9SLffRR68-e6^Y/Zc9C;M?WabK-S_57^7,aa\/SH(^R
4U4E?92/TgJg3=0-[BL.8gP43D]RQ.EAKd.H/NO7L389[Y\Y9D=)A>16U=+CP@SA
;B;Ug4WS:6>FFRgNd(b@<Te4/?(MO39-+N4:7Odc7^YgI(G+DHS_.E:cWPQ3>TQ6
@STO@d,PL4^-)96:Jc[8f-IT^0DWCHTG>g^O)/0A:3WF1^P+WeI;:9g?\WgM\CbJ
a^/M]Te6T4QO5B->#SFU>HT@P>X@UOdK14)I:Y_8/7g+;5535_dG;:7WeNA0H43R
CE7D+>9@,P40f]8.@?FYPL.g^_QS:d/=cYB)5#20VTg]<cG/636+bR:2V7Cg?fab
JD5JU^98EZb&gZ>LK>&)GCA#(3+>L0bN(bS^Mc^ebJ>dUPK5E7MU@7F#SXNZZ+JR
VX7PJITU.^W;;S]9:fHCM-]O4QX@JdGLf/-2F_eMRaa_<dJ6<88;EVZ)>VQAZ,E]
T3e&@G(?_fU-@\-.YQ?U)gBecH1X99&+,F(XUZ)A.T]AGU;1G=<;\S8d;6AUSHEN
bVE,PaAc3EQT)\a/R>JW7fC7Ua&2d+1PeZbX@+O#,NDgLff\MV4.Sb/24P7JPg65
48,Q8KNHV5bL((Y2Cc6=9G:;KHH[E.JXKJ0&=?,&=Dd2/7#b1V=7=O]RSb:[e9JW
N(GB\LB)9=B(10<I+aXD:aICA,9g9;+IRLRLFeARHc,H-.aYO3(aB6\[#FOC44]2
FaEO#TUQY;Fb)R=-[]8E;HeO5#L)H5)gK/B>[AFNc-\XgJ?=YbNc86Q@K\UdKd2U
];=MHR8XaG^_@dY3,bSNCFF#&PG5.gH\&GaE.(STAG=TJ)9##d_^N/cKL4)Ea_V2
H)G.2O0<eU.6d9(AA\]23@^VAPNcVCU==@DO\b/E#8&R6<cd6N21eeJ-HZX,21S@
HO5)\<.60X9PN,2Sa45OUCAg1D@(]/+-W]gUY6++IGPaYXK(<5JZ#:1CN63&099=
SFNXFV]:OcSBNBaLNB@f6[U50C&,#D:OXA[1LIg[+S,OCJ0GRW2Ef;-)c,@RC?1\
8/3,@Z;AIgMFBN>CK(.=RB9JMAOWP?G4Bf,27.+dD)C#\U<U;@bA)>eP#,KALT]=
&SY>a4cC<.IBbg7<MgVKFJ8[6(_MWF&g]T_N&7RKFb.;R0,MRH-ZX;HJg2SS0+HG
(dU-2T>C=PT>1?Ne.H2<a>8>L+[b15(JgL)A03<\eWR4M7gG7HN^YBFL+?K-\]-e
,Q]^EQVTf+Z[#-19_8d0IOZ<>I4-a\BGVM#HK&=fGb]XG2O?QGTDB@ATVPQ#N:-V
G]H<CK;Z;ZMgCcMP/A#MEJdT<T@b+4KbTQ(2>:^2J^Hc&C3V:0A]09<Y^YGfcc,c
NQZ4e9YJZSfPMVH8::K1.T(;fG\@A;L4Kb+.8:3ZNM2cIG9NM1[J<[+\5b1.U/Ic
):16O/c8G4X.dg@7d^?-2F810XLe?.bV7-,]PO?L/VP]RM<Zd[7_MS#8G>YX<Va9
\,GHCGQYJ,@-)12RU>5@6;-,2BE#0HI&)ZWd/ER,X<)6&ec)ZDBTgA9;BO:dA(^H
]?=5LF_Ee[&g9S+8#fT5g-?bBeP_QY/-LFeH41D)0MW#\U-LGe1MP:8^5db]-?8e
&G1dAJ&gVCfKJ;TX-[EXQL9?HGF]MFg1_V/d<5<JYWNWSKJGE_,E)ba)Ob&f=bgU
8T+L0bc\?SV(cRVVGa#)X0)HY[g]F6dRNW?G#ANLcPCZUfQ5?YMdB/>;.#9D<)HP
6=;\=BE5=RSARJeMgcAbG<eF1a@:))/:IKTc8&]eM0T#M;Of;QV43UTL7G3d4WgH
C5B,B-^[?B&^&ME<#KH5d;e:;FO@:W,=FP;3Y._6WIQ5HO:>US+:&_ScG9]UXb)>
+4a#b2)-I^1R,<4TC@Ea/e)@GM(U3N@_Q1X/&5Y;+fae(IC5d&Y0:@?,OYW?U=C_
RBcP<UI]G5SC4g2@+H0(^4,4QJMKa:g85ba58BMA42#.Q2g/G6M&Occea5KW;d6H
]Z,5G#N?Y8X..>M.e2WBJ2PF)F=Ka[M_4D1F._X_8MI0:bDV,=VaK;(&?fU+/Y-H
a\6[0+;Z3QKCgCG1E6DYX>TBKFK6e&F7fPNbI\W]&W2dd83C#:\I@4B.GCJcXKO8
^5aHBZ5Bb-Pc2d1VDZIYJ]45+JKY_cK]+6>5?TA5g[=1Jg(]/IQECE^VX2@;2#>V
Z7eIWTWE2,+@37;V:fG:Y/R=\P&;122Ab9@8c^)_E[-V;T:@PRKKD1b7HUU/2JFe
J[V824,ACe5fU-IMXE1P^Vg2E&5<M#YXeW^)=aVb,4U<bP_J1Sf=/D+5YH@5&NXE
:1-C<\T,=;GRe;S[a>_bcE0@B)0S2SAgNdYgNSDCF7G1+e0&g6]VA]Z,eIM.BN(0
6P5EJa]V2O(C7L?f.A7O44.;-.4SJYRfNDGd+=,T7<e)N&D6#Z(2\EZ(+1JW13#=
C3\Fg+=U<[^;A,QIK+@7<RER>VLM<\V5BeQYbJ-?:ZUT0@KN./f<eO(\eU1cXZ8)
M.)R\UZ=Xg0faYVW/F.BbL&IR,\dPL7AQbE6UQg1(0QKW2ANaM(JaMT(;#MO9M.+
\FK;6-)6b&/e(6+Na#J?g9Te&?5[U3aK9b-V-fCZO;F_X/TG\TBQ1GUJL2dTbcM>
_L((\..eF=-YQAOeKabP66K9@_3BK?gH/gO^P9c0<-d49XP,7;-)Jd#M<SY8,2XV
&cfMJ[Kf_U;O1Z6^66J0&[\@FEb#5bO3RgVR:-?)?ZR)ac8+F#fE,(><=\#5\N/9
Md:ZK/L@IFJG\dDV7YMKdD=1<G=WdUYf3a,9P;I5bScB:7^4W[6>_PP>0<0[]0;K
J+K31U+##DLB2bXG##D2+NIXBg/?gG?V+7L#)F&K,(BLB^;GGea5a@>Ka:FP/N[a
?>.E3.37e_Aga)13/ga6S6W=C?/.;1<@XHW(F1R=<H0Sc7TPB<-d&]ddPaX2.JJN
TCf(BE(Gg^Y)H&:0^GF/\W/KUdGW^GT2^RA#@3AE95AE-11f<VZIfQ=GU/Qc)Q_g
R<LMV]Hf2&R&@a&0gZTVe.3SEM9;P_Q_-5CGNPg>B+;ER<DW:<>9#9:0bI363P,Y
a#.IE2;&?6eLX_4)[/=JI],)Ig5AUe21#(:PM7:B9FK=^\9M;86\JX1>[(d_fX<f
TB8:R->4X,/:RT^<GV:D^C8+g63S?.C3/40P:5c3(AeJBD+A0UfB-cY^5c#Ma9aG
EM18TY?1+@@NGVT4K&8A_HQU-e=^JOC?1/g:]S\DRNOe5@gI,W>:QP^<0fYTO0PN
cU2BV5?[Ua)T^\e=XK8a#OXaH=;V6+SY3.:PES\>&b?Xgf[F\#[Q+P9gf4f^/S&+
QQX#9DBCFX3U=M\bBWeM2JbQ[)W,(_F4]EZ5<B1_QR^<9ZFR6;c,X:M5Jda35W/E
Z1K]AYK0aDJLC_GCAKTQKU[VD9@SDIJb,0U/F:dZ6R+@NZ]6\?YK7GCI0I@8U3Qb
0?4W[@=M&02,M=b6:#5ZHJ(-W2gXAN,Ia_5)U@RZ2/RJY^DD-dH@MdSXaHO6.6G_
]D&fD9>@)JTM>#g3RI/H3)Y0D8_WVUER78[?6fLg;6a87T.<;/aJ9)98YH:];>,b
=YYb#5QcaVKBIJ81W_.QY5_PF.+&,ST<M)X79#QH7HR<0J:7)<?N4#<WY/f)Q6b:
R?)ID><TCJMP#C&.633BbddYTA;B&A+C&O\JgUWe&JFCM[0P?<g?PX?^-+f0Y,gR
[dXZ0F#ORBHA6RK72OU73@X1>dOTV]U:,CbX35Sc]a6a?26M418O-&DUea7>&Z2@
+OQ-8F?VAK&5SH<GbReTT^+&Aa+9F@4=be:0Q<DdgH8Z8RG/Z28FS&@TM[AW783P
>bK#&IZ@;&+0_-EDe+#>Ra]FcdI(VXZ@3IX^Y-UFVD_??L[-X7fe=N()/^L)L:>Y
E_;)f\ANGJ&B+5/dA7SU9C46=W&c6&M,@MB,<5G0Z2&f1FT4Q,:]0L/LgBK#Z2WQ
8@VcJR.0DK@X=g5d>+A3IVYYG@aZ:\W,V;ZgP8L72PGFe8?A939<,(O2,(a^-7TS
=_+Y7e:dQV6O/Le,gN)WCI7O9\8S7e=71RP9F.Q0#OFRFQ1CSD#F,L>@+NM.(g1M
MD0H6_N<AJ/#1eM;6ggW3X4d[D^U-_07SA^:]I89Q><<6G^)GR1RJ>KgAO]B4#HI
Ad_2V)e<g&6>NI1N]eVJ[=5DdcO_#L=^@d9ceDc9#1:Ea4BReJ.+3LR62B)6dc]d
]HUNLW+.U=M-g;D^Z_UHgR]Nca?3?VZf#bePT&JWY73ZS29^,\R33Z?:XAYIRH;&
Ra,Q:79?c(LRS&7abE36<2@@9];aS^W9K48V+5-#.0<MGe/8#YCX/6-Bc.,2,B+A
\2=(MI1PW-[11]GRZ&^LcS]]>Y1>4U6N/P8\Y-=[,)g1dUSE-35bG<7/Y9#-]H9J
?G,OT@2XBUYSH9XFWc;DX1ORFNfS<&Q0gKcaLHG/Uc\NZB<6C>.)H)#FQ>SaOS^S
U8LL#ZeJ,^9<T2-eRO+&KLYAO54-bWe7]QbWHA)]^L1/Df-I#++4A>.6PAU2X[A4
FLM7_4?1@HBWMUJ_PZ1UB_;70^(E^AU2fP_Cc]-<[YbIgS5L:]OXH(<:169dA0B#
;b)\D[&AF8df5GD)+7(E1),Rc]Q0@-[M^U>2PG^RWc,0Jb.cB#D888SG&4HfHM@Q
.Z\^9cQDH98J2?d\4S6+URGD;MMZ/1(^eQKH\AAN[/9GM>7?:WO3VdKbF^M#<.K9
O1V7@RSM0=<EG).b,F(Fb1L5Z8QSdE=9>bV(P,#[\_U>bN]g^3K,&X<(RJWg_5=0
f3W#1KgS7Y9,-TJ5)M.e<A^JC:gB\E(&XMGa68OBMXBG^0C;+5K2\,Y)^49OIO4T
IEFbIf;Qf,Q;&JHE-78VEJ[2434ZWf02c-e:G,2fW:]LF/gdWLg9M09+aHE9>)15
S@)C&I9KZW3BRK]6OUXA?;&+Zb3LQY49TB5090@^)YAJIQ_O-HP4L6L,GDcPORcA
S5?)/52Gg6H6,_ETeWQUK#F3Dc)eQ^517@39&YT8OHSWF2PL;SZ2U/E:[/(GU(5W
[@a6gB]H<@[5BAW-BC<Q6b0JQ8Lcd:JJd^H+ME@Y8ZNR,H)D#8LVcRGY=,7ZP4+;
9;b._5C/;Q6TE35WV^g_S;_e8,NZVW#M\EKJLSOGBD-Y8S@aCQP)fDXfQ8;@>+CD
LM/T\YH^97A0814)V>W[ZfK([U^aEO^)F3bE&>cGOE>gdY5)?[]-cE1N>YgT3D&Z
?CY8K0/J&d5DbNT<SV4>..[SFZ,ETZ,g6KB&Y/2?CO_:/&8-aGL2f^C3EGgS.d^b
:CQDG\3@ZQT#/cf+_J3=_;IE6QU=BL2H:F=8O19>J_?CZ_Ce(I.Q#Z<D0F(;(^>>
_M+M;F-B,+<=6;.?2:SeI8X+:;MgQF+OVT1ICDb0a6R2Jf9_1WULCFM7bd#OV1[/
Pc,<XM.67@/N>W<3X<a&5fBX43MF&V1DBL65A>@HP44HIN)gBK,J].b=BCF+(d)K
[QR6_gJTI3MPLV81;e#gdE-@aKICCI;V]YQUG[NH1PQ_63b1)>5H(_?X9DgaL)>M
#VDOcP;BM8FOD4M24_B?E/JSRV:,F(D2bYBeUB4TMIGFT5W2P7D,FBS:V+@CJ^P#
MQ3L=R\ALdbQ/Tf=W86(Y0e35b9TXZ[89J^?;Zc2Y)Cg^7Mg;A<FGIaMTKM.,aX,
?C9)H1J0e]7eY<Y7LOg_2;_&b?C>a@?6\AU=O,##+QRNX33I^cJdPU9cX&gGeX=Y
GQQ7]SRT__SQM9T0<,3E_,.CZ@^OC6OTC[20&FE+G[53HFeRc;ZY3gd:HWOB1&?K
e\;U4FF#c^6_:Q3[9;36=)2O];U_d&_:9YB\19PJ4,T(d15=25,J/PdHI0D>;I^^
0CH3)Ea>R?9bS3X_(F;BFaZ\,/\FII[7V&09;b)2A;8A)WcD[f&@b4(2eFa2NV9V
gGd;-S<[^/DW.MK(-4DHR8-7Q)<E(BTH/G^SIQ6J@c98UGYPU01EY.ZS)I<:RA;.
N)?SPbg7f:SBgg^g7/&_EBZBg)/U7#;188\/daT[BO?bb,:HH+C4dNWGgfV#eR0O
][Q&\QK@8ca<#OGNK5HeCd?>/IJ]6MgeWI4d-?CP_B[]c,?F7-dOQ#5g5c(@A?QB
dPgS>2_.G_4-I_BNb4>/HPIIcf7+S-CGe/,46277D)G]=;<I+7Q)eed^fIPM43,I
6&CeD<X(/1Qd&VZeW15],C\;=eVOU5ECTUE7/<N8-+3^PLAR9+cQg)Q8a8[9-P_f
OH[5>WPRL[ZY6^5#9SVT1)?EX;fC-[]Z<&Y.bOR_@A(9e=(6LCZg7LKeMPC06O04
(P9HT4>LTbF.30GN3ZVfQK?8ZKZW1#K-#X8,8A00/-d/1RJdF1:S1FJN[.]\\TE(
RI5QdPM<1:6.B.?MBg2.9HY_.c9?=<]Fg@5(0eRIAC2)U_6C[eJYD69g&b74C[=Z
\_dC54\0D1GO(g?,\)[MDe5BV3;cdJ8&VQ>.MV6;gFTVJ75=a8Ad]WCHS(/SZ6:.
YdUKD@@D_>He9,Ub<J\Xd.@:2d)]>NR()^VDP=HCJ[Z@DHd4:.b-e>O[cN]A&c/6
Rb1eFgPZcV[7Pc^.T/&]&GT?+b.4T86G3/DH.>/5c=Z&2R]LT\CeKU7E3-4N5F5e
aVJXF0XC(#XcM58H:@0U5>P&<?GM(M=FJR2J[W1AK48A-W68[Dfe[OWDb,EHFK@6
11<d\?^dSDNZ:,P:5/K(19ADS4-NaYNHffXcB)3IV3IY___AP8?TCQ2/#-0_4/ZN
aX#+Lg(</@#,KS?5RP6)GHV\,(?Xg/Z<-[E;4CNIS2C8PZb<K6^Mbc=V_\V)(@b+
J&9+92\@WZ-gV1eW5QWBeF(Ub^&JE,@H]FBEG6ae/@@A7A81B4GO++/:UBTL0[<A
UC\\\BOMD4>]gQUH7QEUGAeW][H,;&]>A@-78CJ,1?VBEH^QKgO\C4C1^\2S(f=L
.@1<A.3-A,P&]fX[ZV]<-Y,5[?XQ&X>EL<S+3TeXEO)WJAX0WJ@KU>L@G0B1bK^>
,Jc)<X+SCdQ,;@P@e)7KW861+\aS].]B_=3f<,M20_gDNd<T2X?0F_4+ZgY7TF/e
F5E,9B498b]^-?50I@#DZC?[dEa7AU])6g&<W.1B58E0GcM2#-@>J(;;IAWS>-VY
Jd@#5V22[_W9PcQX0,LTT+I42?=/XILfE^CZ&R_cCQNAgF]<c,)=ST06BG/8@d=M
P.W]C]F(A1<XE=SY\+K._d=)OJ^4:053BgQd(<&>T_PJ]1WJL4Y?U+gLKKbQ-(dd
b4CHf6X8XD6.IO&bBG)QA5EgOdD2e(V8g>b&#(UFT@SGA[643\K_<,JEdOGBOM:Q
P2ZJcESW^Bcc:<?D5JQ1Z)V2XM>]Z#SJ(=Nd;+6R2Se]93aE5[-4eK4LZ>5B1>,]
6<S.^->=>29].-YM8)U6aAeK(?AF+aXd7()D6#Ba_HJ>X^7H+@)^.eV?AI^WI,#]
/c\\5/I(IG1)T;)gVJ]GG:d&c[X21P#[GKK(<VC#O1_fgG]\>GOF[U8]30BXGW(6
TPQ]//f#O,GdEQ@U,AZ/WCQE:?;[AY?5c[#E_&RM)1&11.P)g;K@a[G<NIf#WU>B
HU9#IT:Y=-O80E0&(Y/AcM]7V0H)77/EFHW82LG^R]5+UUTVM-e:],&d-bK/d.g.
A96P/.HJ^CZ\I/X@U]=8g;K;dOf=R.SV[9U;4eS0S&FYaVdgXNUCYZV@6QC)^\:4
\\bLWg2#P(.EH4PQXK8.=K)?\@;RN5/F(ZG&7H,/J+H^eT4R^a3\?EJ3+G?UYC9C
+5#_PTdHM-g0<)O(D]&KVB3QVK3#.Y2MZb\V/Y4T\<a^Fc#B?0a7CYG?a(B?b>\I
GNG&^+MbE^3R\_=H)(,OYf-;A34BB#4,Y:<@6C@1VI;(3C.T25(U[8afB.VBV-FU
8W^4@,SHDLX/:eW2JP#aY[Z2OLg_#[Og^VY;JFIELKKBE<QMfR16d]8A\TH+91>[
@6dOg&A3P(S[/LFOHR]LHHUg+(D,,88;3<>R/;B?FH[cW?d\D+d3@D&6F,>0L>/,
UGFX7b6ZBV+VcJF59(XL2d6DI?S/FX;8Bf/LW,25;(XG;/.M36J2bC993Q6X_7-Y
9SVfB+@QL?&40)<OfZ_DWC:CM63I:7LK5cPU?B,W=]<K=4a)U)3e>M,+R\:G+_2[
c-5<cERbVN^0bIL@AT&(>7BL#E?(\ELb^<O)?NY7egBD8d.OgXB8X\W#?4&6,dZ[
LBX=;YRWII4]9D-7GH0G\a?Q?+WE:CcWZ6RPD_]^P0/5GG\VTg,g^8d,TLQ;3P6X
2fLKd>GM&D#^;\@Z<JPb+gI:1b9-@<4dV#)L:cB/X/LJ<^<W>[;.gUS0YA]\HIG\
<Q^(R@B9/4=YKbT1<T;0])3\^03Ka3Q:3+bB+G31/b/4N+-KgZ,>g(&T?VQ?;)Od
<GJG<Vd.=H9VCW6X&[&H#fe7e@)PNK;fC@Hf;eYP:YOa=#f?/6aI[OM45A+V/2C<
HfMN92688Z)?DdF&5QKC@>_;-85JN)-E8EQ+<2DbJNV.cPJF<[E/J^Y4afXR@<bM
7b,a03/S&0=VTdI,FFTK##+gHBb(=9+ZB;ZYZbY>Q@HW1Ef8QLH8Z>+b-(;T-7:3
eJN-C:_JK([6_E[YeFM(-R?3fdR8)eSD5.,7TbKBHZ.c+RH4cVN?G7.-\(#SN7V[
M0TgbU1a.4=@_e^:W0M6LaR]BD#d3,/NM9H2WEWT77HD4/XE7#;ZI8))Pb@e])3)
Bc1#Q\^U\SBH:4_=5?AbS(H>F7GGVO_RW@<.A\OUB&?-WZR.fb5;eM,-I<Y:Ea<7
_a/)(aH,)#[5;FSX2e)Q3R&@dW1A,[L9JH&8:39O?_O_:U4<C(36<HgFDZg48(6]
R>8&6@/&:[T#2FXV+aZe[95HY-+G3\H?L>-B,A5d)K[U(_Z6V[f9ReQB5MS=LI:?
]<=YbWKd4SME=4g0McZ\eS_bLS9WfVVT(@R+G3..@7Peg9W6<=S^e[?SZ;S91gYa
-Cb)0D(H^WCOd;M-WMF9J,bDcS(Xf[GWPZf;&,;843S55-K)Q72O_f,ea>..)5P.
3dPWQD5OF&_5HJ^H<P,K[BD7#4I9>E9[V/FH[GQF/@Z[1PF@.D&6V+/JWV4+P1HT
MX^SS^e:cR[EV-L4c2gND3TF#cT+1S_=L<WWG8=9D7Q;/BYV779cZ?JSQ4+CQRHE
7AR<>\0?WAM)&7F@1dG&dOW5C/a2V_@>V[K2+P@V/-S#cW<D09NQRWX0WT1B\GK+
)eNY6c8-c1WOFE2aJIbCIgdVRdMW<W1I?[VT8R,]=]X.EMUVS3QM^&&&BGSa+c9[
&Q(NPdcK\&B[\6#28O(17&W<a5\_eAT2NRTXP;V)26<,I4V;(<J->Pd^cT-YO@/J
GKHEC0D(AJeVb#L>eU>R5bKYMbL+B3fZ^QD];#,ED[#)61VL[;?YQQOZ-_<&f75)
G[;U_F).HHQd^GAR)-;5=.UB<O:^_F@^.5,F_G[a2W,d,_gIC[NLG@PdBgcOE9a#
(F3W]a/+0WHEbgJ[D<6cUR>9/?LaH^OebA7R.9BgE^>9B)H2>+c&D0+:3C&)3ZCQ
cQ\>4dW;BOI2B[LREB=I#LLU]YcQH3KgdBIab5:d[W^DN14c,:\gSYVFMbQ#,O81
BA5a14O&YTXL^K+2Od:cNOPcFce+I<#NCJd.eV3<>ECE;#(\B]Q-Rfd8B_1TGLEN
dX?WUTIP>VDVb(d7]I-=bIVSY>8AZK,,V48E@?.:c)VZ@H@&)=2LV0^KX37#EC::
FFBSeIV7M9>aO<EARYY+[cX.:c/HZZNf1#<H,QGH])D#+>2aL+g<,<=DVN+8g2Uf
ZW^73/07#15=5PWdC[UKA1?,LCOCa4.&28Xg=4P.U=#W#(:2@YV4dY&[;:,.(K8\
gUZ<W1@&2>TA[1FFTYN36DK[ED8[C>8O-Q9Ga>56K08RB0cX>80S(cPFURVcWG\O
BS<^8Ze\Tfa:EeCO-AfFUZ[I6Z+1[G2HE>GY3M_ZZ_NA7AD2+<<UD,(YPd.c^MHZ
cZf\P)^@U<;NL]W51e?aSd;gBgYa:eBZfL?L:-agH&JCXYA?Ig:^:JGN+2.(0.L[
WUGD1G?):Kb^Y:?-d,&;FGY>>GP+C<4#M8bA:.If;UU[S=#(7W7&L1Ob,SXcdZ[-
,C.-QPC8V[EH0._)YX^SW&;E_9>@;MTc=10M]5I(KQA0[1f2KaMMe4_W)FL/F?/U
W5S;BOdc]f-fMX1_,5:bLd[M/gXf6,/-==4CF1Tg^W.3ZS&dB&:STD\:/K]/V#\O
72AFE7)d4>.4EV=-b.A-VN]bC<JH=OCCFBRC/BVK6Gc9V)LU7RIQ(+dH=44NU&G7
;<O@0.PY^L#;Z&gX]<:G8GN-Z(_7+Zd;9<Y2RJA_c>J:N]bA=/XW<[geN^,IQ)fO
+^8PV?c]dQ;?H3BHA/@]<ETaW;X^eVVNg)CUP\+@T;W<C8Y:(J5PQ++\(8I,)81d
EZ?<C1MPG)NCa?]3Z/PD;8(<eU=d;(S9M]L[d3YSNAU_S5R:&UafbJI34MQI0/,9
WR]RT5GO6_9_e#4d/ge=>9>Hg+YBO.N?2K^-&<_#VRF^78H^baB)=Q.eS/8e,S<G
C5D^LREPDC>V+Va4RT:0Q7-Z-cL3]5:McW(H)C9DN50_AF4MD2&dD07WI8[4HQcg
3_BLO-QN6ZBQ@_99P\aD.84=NQD[3;N-_Za8:7;&QGY6^NFgUREG&@G;.-MIDF]U
Bf_EO[C=0OE/\RW851aG?_?6O@cTC3;aQ#A\_BIHB(D?M8?9>ENPW?:=5]S8YKQZ
6Bfg^DYgTN:0?,N14dCONTMZIY<BNT+]P/Y+)2_1GCT3H;,eG80c&V#<E@/HFe4,
\,C9/7H=]Y[aPd^A\Lbb9@45=faI4(57:&^M.F:EaICcSa&IfSY#5W;:]SOg63b9
/L#_T@]_7(XR41<1/Y[]Oa#NWJ.bE?S-g@+^\@^Z<5N:8TbO+<PI5RFFVA@>g?V-
^S0PVf=8+Ud/GSVb2HY=f0ATL]\2/V4RP/FN.63?T\a?Ad)+JC+:K[;PWFNK8LEB
.[MU^Mc?DWU>;WbP(,<_C]#GA6H62KPfS@9XVB0(S>-P1P65K7<,->#7(.S&I^0;
26X8cUQ5N\N<(LO5P?]8F8Y_b,cJ^31+2,&=)NKNT_XK^?S?\PCNb.O+gTE(3S0I
?:6Q_CS)8M4#e3&)=G27)d)JIK^(WUZD/BIZ2TO(X0;IJ<+e,&?:SMIJ)/=AI8TL
W7f08L24M521S9P_3g/ZJ>&W#14^5&4FMG30=M/J/FYa(d9a.U[cSTFGHO5RCILb
:7.,eOZ?C[4;e?SeRH(QMI_+aC,VM+>A1Z5-<#)VGY8BR/^^O3=U85SEe7Y2WD;Q
Bg4bbZRHIe,Ld)DSf(Yc^XNcHWI<8HB)_@W()<e4/LG4JVQU)HK@C?RNQ0<FE;Ge
&;:I6O):E#?Xd^6C#7&3cS7=Z1RQeG3_T,N)2,_OEK]bTT=+=J,?G8aAPNA\)G@/
JW<XD>0DGOX9T;Ve\+ACdHHQ-L9T@OGB2Kb]Ag/3#IZHYHVVJQZV]f85_g0RQ<PB
b:GS,1+AY7MO[Zf(fe2>c9&c81Q@L^MFA:+;1e7LJ\H;BeAS67UgaN[/T:#71&>e
.=GA,250@[5:#0L3?d)>1)>d5^)SPa]d\OAX(0,W;5CW9TI\W(<1O_ZVFN^b.OV(
)a)Og:Eg\E]&F;F.#J6N]#:IJ[+[)Q,U4#8]]9c-CTA-&L82-+DUUX9e)1GIfGR)
B/\4](fJ5@-<@C4gWU:5?T.WJQ;6&\db0OeYKcfW-=SV6#_5B7L=1(YYO/:[LNa:
I2Ib71g#@I5)B,G;N#OX.>YXDDb-+WcF(/3BYVFY8S8K=<<P#gS9I=cWgK3Z,a1+
C-))Y:eL=faO-=5@#.NLMDfEe3Z(,3[bVY&R@a,Q(.9ceS=X[dM[([)PV2(E]3[\
.N7be.YgFRPA49[VNMEQ3+.CO#@Wf),#(U/EQUN_E8^DdG#\3?8;f,JD\E.HX?O1
/^3)/W/@UcH8[LfB+e2<MMLSMUJ+<Cd0L^\ZeN]6Ee\Z[g;?4Lb&B-;1+TI)26CK
+QU#]P3_E5(#OfV4\FT#cWHf0^X>)<BeXIZWP(NEF7UcV#eSb?Qa2gbMQ@1B8Q2[
9H_-.[QJFc(G1:<+7RNTSB/5G(3YPVTIEE-<32Q#DC[_,cFU^GS3F<J(N3)WS,Q9
UCWA(HIOgLN]Y9I0d5QIY=[bgaFTL=SJYKaXX-M14-II30S2?d8N.R@VF0=_gG&6
08f6FdRK;e#cTe=O7;OM2]<XEDUAXRJ6Y.-;CB+bF>f3T@N80C6_WN6Y#0DMJO(#
=<+XaO&dAJ09)OQ1WQB;ZP#>IEO8efFL6MZ/Q0SBWD?R:-8C+?MHB#EDMY:g?Sb<
6HZg@9VE._\G6B?>H=)SCIda8JK<=)g5NbdN=f^)YHa43OBKUCZGFgI6;@>]E\9[
6bHG-0R@W)J_6XMQ_b&+.&g96^,?3E9F-#P7P0@4gMCf2BLX.8gJ7SgQ6e6O0?5U
,=WFdZ[I010=H)e(=<C@:8XP,/XgLU-dIXeR@Z(,^<[HNHI].[G2:<:N_gU184c3
ZOg>RML<\J&PYT.71JfIUM9V8ZO#/PS___JWWUO(G)\Id<XTX19X_Affe:bN:UA:
AIETb=C62IaEES/3FD)143CP]PR1g[c:@LE/&e\d+c3ESedH.gZ74#GfXQGDI:Z(
/LWBQKL./.c0S:Da/2C+7,6VCbS(C#DU,dN#,V+S576d;]cVXTRL8I+QI7[)[GZS
Dg_WU<0d69>a-X9J;&CH,:&KUGOd\T9T&=#1?=.\_Y9<a@\A+0fP.P8Z4Va?A2aA
<FFKO_?5Sg\M-(.87X?Hb]gV5[f+YOI@SI#bN#ML^6Z2TA_Db2BFK2gCB>f=.C<c
QeL.V,VGBGKWI=fO(,:Wd,14D9K]O4b:25ED;Q>BG+W,?PY\0/30-<PQ^S.WeP1<
)G63-QF\0O.b&-PA;Qa>ECGGF4eX.HK+,JS?8/?)9)B&PW\IG]9TaKaGF/D)c6^c
<?ZdL=/[WAB70KZ/gE8;>&:f@6;3N\:Q/3KD:U?[JM(S0_7??J6=OJb\=AfP4=+\
:G-ZS73aTg7Y<97E^82[X?TDOQd)X/9cC+2WaA,W@<[^=Y@B]cO4XbAT2KND6+cP
3(.,G7T^C2-&d=/PJg2Ja.TT@R3XVe>?TM]FBKAAPR9e^U6ANU0MVaR-(9fRXLO0
7N8P(K>76@7eb]V?QZ4#+)?@M?K:4FAUQ=^A5EGCGSfRVEeJX.a&MSac0fQZgE14
b]KeAd6C>&/PeG/>;8Y08+e(G\1cfTQ_8Ea2>9:F?+Xg73-JZAFC/C@O/V9UX_5N
MTW81.QAEJ,1UDRHJTI/UNW+V7H@bEaQHHZ:)gH3,ME^.Kg8JdNC^9Xf>#D,(WK)
^F:Jb56V9-_>&(a#>-GQ:[>?#PF^a=Y8996N168b32IQ6(JR&H,>d1G?[STOf2Y@
\2:E1PJ,ZIBK3@e3/G^^(4a1<P=KMI]6fA_2><6?<@e2/<;(5L&SGQBWZFI+UYOS
D&<Y<b94\c-YBZ;V1FaG/=./QLCIT/4>##X2,\Eb9-4V>_>OMY,3;NYRS1(5=O_A
&DS).EYb9JBU@E,RM<)[E9=[;N=;0N@Oeb>Da<YPN5e^J8.MGDZ0b^98=K4=.(5d
cT#<):><D7Y&ecY<5)Sg<YF#E,ZcXcfK?,9ML@+AY@6;EVB-5QUNV7WGX6(0H5=]
IU^[QDDFPF\_.=O4]O6^d8K<d75R<;_-L<7?CJV-#O^UG8&Y\C->Pf&ZEC&<Uge^
7B_BU_&?JQH^5(RZ1Pf=f.?-)3]B:N9TKNX&GG^Ff3AA\<NW&[65+aJd3b4+^Yc>
c?6Sd@>V_Og0L3N[/L_;2JE@I,9)bPC-N>:XZYH5S<O\QYR:&_DPJT895;3c<8dT
F?=U:f\5/..c]XJY[6Z]62M8de2\8.\S.<733-AP.P?[&?VR?W.<^G,/1R#WQ^<_
=_3Id;]=Q#OUfa>OUSX;EVV)X/]MM+F1&1H\>?V9L-\OAUWA<3Q03cH^Q.fM1)d4
/)>g?>Ke<&7)LY=E)dTF32LE.YPHX]?LL7]>+,VfN5OW_\:]Mg=/R]b9+5S>>;fI
Y>R1-S;LI[Y-ea9_5B4+-=Q)6T_gM4#3YQg6dMHQGbS6:;6RS<T;@>bVA(MG0LJZ
df0\;8bZV_SUZG,NWV[.=c\D&B#=R?ab7f[:>HWS,6EV89A5QR,+@f[e8-ddRBYH
HK[WCgNS\.15-+[&^Y]1><Z_\^bFfE2^fc>0J&9-1@KG3HgWc&GS23H^#A8>A9T=
GBJC12+JHXUT?(>L(+Y(T0>),,(8?c5;cII>OR3[O:SC]IaH:/@/dC,I9SLS5O]2
NLaSe<OONTJ:07FId-RP(XaQ@OU.AKK>XMP]MGA^A20N=3IP\=.B)P?^d+HB7N8)
9HIB1GC6]2_1+d=J_d1N#1bSF/LJGeMd(2JWIO[KL>BN&3R1FB(VYNO,B)-3&W31
5D,/</T,:]X.@(Z=KX/0.QUe;-]4eB2[3cF1Y^dK2>[NgU<W+9c,,L#NJ?RL(_=#
K7AZ,(KNL#KB1O=Z7(W(#6,(51;[#YXCW3>c?^f1Y\g:a7BHHQR.2)N.=@K9c^1)
X<E(#&N>REg3^<0J;W^BM]T_P\I9Y1[D+F.VC4:8/_T550RB=R8fX,H2R1IF\\+d
f0A4ff1T)2MI&]\WC6/@<f+g3]MTObO:5CYdId4T-=LB>[gR]V&(X)S#:JM#a;:C
@>XS^P=eRKL,M)^3/Mgd/PPP1NObSZEB3MQ=.gNd5;191Q_@73cY\EN-2;I-b8f2
MOd<0=865+7b-1;O4+RS5U+=9\:c\+K,KEKV67Z@#J:/GUTCfN[7X:-fQK-LN[0]
f,>,WI=Z3V5?Dg1gK3-D7AOGW4I?,+ZTaeP[\JBWTLKMFbQ#\CNYZF6/L-I)EYAc
KW7-)4+bbG66>II906_PNQ5A?b1>DX#H:NS14=SeaX^PGHX:>a/L6G>de>/AW1[8
.==&0]UECXe_GV1AWIN8EG4&L4#J(S6Y36WUXM9;FN\/E[;A/=[NTF9,^PR-dY6_
:&Iaa+7I[^NB502Y_5G?eQUg\d)d]MfE+=:1d\\9>2L-8T&dMJa,.G7&;c(N):U=
QYJEU9];QPAHH]=2)K[aT1NM3=(g)(_<b>X7+ZQ5E7OY-eWI^,8K7\..VfB>b+;\
&1T:IC;8c2.1d&FIB@>#=0L#N^c5<#F+RHc=NN;6Y>^eMUdICfV:^:gWYY/-MHag
7f5\20Cc7,-8ED]dX]gN4g5PL#B_,/1/.]W^DZd)W1afdd@(,=,B+81_/NWYgO\X
H-0Zb&/SdMV4>]+-.Z7&^KVBN-)6[6Ua@EJ62?[2dLUeBC#eeeSFMaD@9[Hg<\,/
(E.0Ic#/]P-_S(>^1gIM5A?EXYf2Z,[)gRbG^-df)QHPZYH(LS\Z5fCK[>26C3/]
BTKT+/K]6;)d_\NHV5C7bQAbVDB]79VT.-R=DEM2c[=IXC)VIeAR7[6e^[9/f+(W
?_6Be[+d\YXfE?fd105TF#fa@@F1TS8F.a(E;b3eY>4X:)HK#LHPaJdCCZA8,+2P
;UY>H9NAc5(+EE((gPgLOENP#CCD4a:(fe++:P]9@CDFJeDSFEcfP/R4_;(RC]+J
H/bP1KX&O?)_;QL7P)ES:;R3NfHVO9LJN:H:a/6(0Eb:PH?#S/5,,SOQ[T,_U=dH
^:,F\VaI(D@YZ6<<a7?T3.UIWSfG@,&PfcCBC=R+EC>b,g/@R#4/d8S3e#dQ&gSb
_gb@C8+FEc[/g/c7LG9WcHV+DC3OWe^Jd]M<@V_cV?dCQ;6]PT+g.3?RN?1T0g1T
E@e,8P:dTT>LNO81)R.&_-8HZ4N.eZG#63DVB0LP>&=F2N-^OQ9N)8gaK12&(gTZ
+M&6gLbfO#<SG/:4_F(SGJb;)^>:P8I.CMKc9S(KRaOfJAc=FC4ZMQJc\g>7,SP,
FLG-Z?MZQB)YPJH5FJdb?>3JX)7-]-LFK=c5P-8:B76QBY\b1JXRcF7J2WI_L])A
fZIJ]ac?aLO[_P3Y;/?OV/;([dYZ3de]e^cWK)TE>9,>Q1e#1L+S7.E^GOV;bfJ(
_G9Y6eB/4&[HZgN^J4MSc:3eKO;]^,:#,g5(N&RT,Q71>CO8B5X[?g\-gZF[UR1]
\VXLbg&3P7AWSaWJb\d-Q6f#.R<@UMVOVg]>^,[fYLM@TWQ]=>I\,<X0dGRIU@7M
4/M8>DWe/eV+E\QO#]EZ9a[cB//@R/>B],D/[P<A[:WP5B=(gI53OXSK;Df^9Re8
71Q:c8VY5M@U(RfBW,].Ke><^X?7aUBIXMO6)<QJS4VJ4)(2\\;f:b-1bCPX,.W4
PV7([(C8)JebDTRE8>CP2H/)5Z&e4DR5F:9a>KbKFRRS-,>JOUD+VN9+OO,;g3GQ
(ZJ>]JHdV^2-3P<ICPSe/L8Ha2VZ&>;c1,YW-JO)J6A\RX5[cZTOSMUGGL2L&V(<
R>CTdaJ<XO9^4C0^G9_eXOV3DMK5\JG9A=&+A:QG(.:XMV[@7^d\5)/C+IV[&d1&
-9IEX6V<45]@JA^e1?N_#KB.2-,/fYC;af-9]Ma>9&YS;0,GA4eY(DYMF.L7.[2F
>+<\eY;DP+X7\WYA3cJ@XJPS38JVQ>Bb48WdCK-1S/aTOYZ_Q/aTQ8+eTPI<N\;W
N&&B]=#dFXN&Ud#_G_7>@Sa\e5-L<:egZ7\97AD&[5GKZFV8#Ad,dFMKECF9;IAZ
C5[]-d#6eXcFe/Y,7@IA/47af-^gUff].c;3Hb\Bc;cB?E8:3U+1&TO=&f;25N-+
NO&3RQbf0./=DHeGA__D1O^;BCcRYPDbS1@4/E_-@E&/Q,,;cP0BSZ#ETBRZ<D]T
OB-:PAKA]&QX1Mf\@UGA1FJ-CE2A3aIb-4>Y,.dY=DQVO#[@;YY2L/)a4c,:Y58V
Ed<MDV;HH,TD5[GW7D.TZ(&0eLE7QF]f_UT3O.A(X5b4S<G74beWFXdFX1:-a)PA
1W1_E[>LbV3Y(eS<8deQ(HG\f-A3H]3NYVV&AYg]ZJN:D;\)O-A^;L>=dRM&GbY@
cA9UY^AT/=;PGXS;5TaBaMgYTI&f=a?\?AH-78aUWN#a)bMW8[OT+DG8fZ/9:1Ze
b/]CBd-,V\94NT+;6BRFZ6K\cN9,fWGNYG>J2Zf/dcAegJHMF>f3+LGS_.^bFZ#f
b:XQ^FU9U(-;L.Zf5,#ARU314/H6NZA<AcBb(PF[PM;#4;Xc@#ELJRV;9<&2TR[9
.=I3W83+gc=FH<=IK,6L/(f_6XC,.SNK-JIPWC&+(H,6YN9;LcA,P;3WHVOK^SW=
>SDBBUVBIf(.4,0G.dQ;3bUY9M^0_EX0E(/^2T@?IaB7eWOcNP.B41SaT7-(e(LZ
1LQY6):RT]Z+>ALe(gSXVaOF4E^GLcHfRQ(<GLV9TTeE0U,(DKY8AcN4]MYAQWd1
]?#EEW6>M4e<S328AFe4Kc_+U92R]>Q;)bERc;e_HO]CO4Yeg=^OZE]8\S?VCYL(
GMJ\8;-M(C/PI=:PH8MHNSee30+C]2#PbH:,I[[R]MK-Za=L@G?3VKO+SN-L+[1&
2<UE:D@Y>-^>?T]PeM)-GT>6,NHK7B?M<JQ2A97/?7#74g(fQ94N@T8)HVMVf]TQ
Q,NfVH@D:DU=6<7&1>:(6gC[fS]]f:)::fd^=TP#=:FFe)4#.J66-A+H3dPTK:bO
,UM#)H&7YYYQ.K]D0TeZ-)]<c-<AQO(&TV@S2+BEegDHQ-ad9VN>gDG])WE55:6V
H@AGPYQ.JBcL+a[<C#:[4UdBDE-d8HdQOUHggC@E.;40>O=V8RMDHC9O<BcHbJ/U
;Ab<=^T&g/?WM(<0Mg2UB^#]e/dD_feP8(>CbcgOYSVRWZ<YQS6U\R40bET_C1VF
aS?&GK0L4<XgG@F+\:A6>C,PFcJ35RH[<XVE33&AW[PAZVSc.D,1/8FU-T4BAaQY
cCG#8ecISKBRIKCKK36=_>)W;X]dI)AB^:/?+77PPG[T5,aY2]NEN3/DOG:d1#@C
Y&U9>C_[GdbY9e.GMX92A&;EKdgQG[/1_#fb8&\7Fg=E2)W@?eF+O&=5X_R6U&J6
>R2=LMRF0@/W3&@=7<RfVKc5@I<#P<N9]b_5Q#3;0)EF6Z;P<M6+WQCb^>Z00JdX
,+2(<H:b=]OQ^ER>SJd-8F4N+O1\a[?M>,]K=Wa3.B=@N:+Q9Z/=,P5+6(R^JWL]
IGLP5TUOP?L-\)a8XU0V&(LSBCF/ZA#+FU8I7VUFIGTeG7b/131BK&V32Vg@c+?+
OTb([T/MRe[(6JH1)YF[K,T:[gSY>HXSR2S>KdI^ScP)/FJe];X(5R_)UD4\7YWe
5I?#S:gB6f]C+Ee9SUR9VCKUPI??HV:8ONcEb02>MTHN\CBK+2bgCGf5DB-)aTUA
X4G)aO?VO1@E0[9)NEg=2VH@/SF)ZMc]](bB0OCM-3;J8;TPFSTZ^g?_JXKYBG5#
&-cO7&0<[=eSZ3&1:+Og>6B,Qa3;\,f94dQ,H9UK7C(&UQ/+Y;f&XcBcB)Z25Qb+
&R/1M@c(Y8aOdC;;6:V1)\CGJLM6<P\+\0\#JQ-10\fHb:CDRJ#9d2DS./8>CLD9
YagI:=c&;Fd+J,IX]M7-2BeJWBY2.@C4?/AJ#^&1e/.2C_L5:5_W,W18A^f608OJ
e4_,ZV9\C]gI9I[;]T(aI\Q)XO+X5SV^eWM]>:.8bOLbTH(ffIaO=.Q(M:IDB>8a
VG]G?Z@]S,&F=H4gXKVHXMVA\VWBB<4_ZNJeY-b34W1PRaIN5=2W/+P4<e_(9X)2
GG18?QNY/fV]7F96A].GEHZ5KQe3Ld5R-EYZ6[Q6-aWN^F##JF:FZ1;40aT<)1(=
F7)_KWH6e94EWe/@&Q6KJMe;GDEb9I#C4:cbFL:)=fdeJ3U8C;7De.96<#f=]45Y
2fVKCgge2f=_VU<_)\,.V\L?H-?a_.=W#&PAD(&D:cgTXGg(QMN?7=7WE>FZ\).=
V<84+=3D7aK(?>bJ:0X2+Zb:HaNWdUJ>9):cAI?8@TPEfW)9TL,GdWJ[>0O)<cH9
]HbdUA,I5AP124Yc8,cGE_1&I4)R)IZLbH0K:C@]6MQbK\?1&eW8)==A0#Af_1f?
]MRZ]QSf_72RN??^L>]A=5dK)I[6cg30WCAP0ST;[Y9SB1I,]FA3dW@BF=00SI(@
A(@2a/P9Dc@F1BJ)^V<+#6>OfbL^b2?<@KCgXXfW-G/N1&BO/6LV>TWaUJDGW>W#
OQ,/0#RM3W6I86YORD\bV@L87OeW;>X:-C<2,2R(RLS1Y.IBN>(gQ<cE/P1(+O31
-gZ)D1;I\>;XS0(a5OGc@;:X<&EC_I??NGf]KON-2YL08FfYb1_.]1_a+S<X)_BD
L09?/S,;&??>.I)bS;NQ_8WTJWNOBa^M9Fb#,09=\7#g+Z8Y9<#X:Z^(R(D8PM9(
C:aYfZ6Z<085C-8\Q^+)T(?(9T:/b>J<S-Z3Va[)V(Aa1fXR-Q1-2[d<-T(I27eR
1AT7Q=EC4D9/EZ06C;S&;QPCc5\G6)8fR=(I6f9Y<.6>:\UH-Ca1SD5Wb814Ke&8
V2JPdV5-+\P&F6BK(>0B>2N4[dMWgY=-+4K>L]D\Je/DWfN@>SS(/V/6gW@[&9\)
<0C9M1cWXZfBT(9U;ad?SVAA&c37=5PZ\4eTLe<W^7/2DFM-0;b#BUf8W;Z:97,/
,GQK6WNU/2Jb^D1>:1Q(T<1d9G<BMMGUXKf?=ORcJJPEIXSOKgJQ1X^NCX(Y+A?\
M_fdT44GJ_@0#e>f\2)=N-)DB,NbGNd91>G0g@gDF4F_N[(_9b)UAcX4fB;G5<Q/
^J?66[@=4#]P\gV:VdQgFCXgF62We^)=,[G1Y5QHgV0HMAe#VNaONS6XJ4gSSW?H
T(\BJ49D(;T?]<c1/CgT0Yf]75>SF/-O[-Padg(BN?-c>.8Wd;W++TR<g)-UMR>+
P(-X?BfKAF:T)9/Q,-_\RU^NWQ.+3#fH)E<EG#=109gXAXLW&J#RZf>K;T,/[;P#
W37D(#&M0>A_F=\XC2MI9,TL;IK7@]D_fDY@d=ZWdcUa#OG&J;=KAA9:\8,eRfDK
5S[b4/F_-OV9DF6Z)d)RW_7D(6OdO^[gEH7dLL,-:NYTXA@@UUSUDc&DR[)V;(:?
VH0=Z99I_@CHaCAf0Y:C79ad>G^.E:,\LWVGA6C]/D:J.KU88=&aaV2XD>OMPZO-
+/]Q]DdARMEdIX[KAD&+5)#cJd#ZG8AC[_;7CTT0_:g8(-DPaA9Y@SeDCbQRB2e\
a0a]KXN+HZ#AXMMcgDUAK7>IPQ#Y/[O/(.X]&<#SXYWP/)aZMV+?+E1LN-HPQHB\
6Y@8_H-R\;:]X#;>#N6Wb?A4Cg:Z>)bg34A//L.;3C]B)dAL;MH_;SCA2dO6.AP>
5eTcd:^RK_fgMJ+EbL50;WbC]CU/6EEN(Y[c3\,_:U;>L_JZ&IGdP8A21c=P6JWS
N42Z-#3MJdO,HGBIV.B21g6O2aEYIGP4B#9KZ?JF?0P^M/8N2a2=TLD5Y9J&XeKT
B5G?c(^7=YURFLWbdI^@P-P&PD7R>4:<J2>]1b1#;R<_8AII13g6(-.\AMgEa\&6
NWbOdX#ITHZaQA1O4>98^,5Z7+aac17(-T/;8D]HPJWW7ZT@+(Z]8YSC^]N6(T3>
LC8,S0R7TG4eNRBT(AY;5GWd6c1[#BbY07\0=e36fRMP>0DfIdgdU9W+8&UA[bEA
GME6H94#[WEe5^C9&MZ2-I(CY0X5=H\Q4<>CWDDXMA7d)_TEI>)N06IF^_QEYIc.
T(\>c>40S)eZ);c,LH1PW6b,ff,693N:Ga>Jdf@XGL=7Af_@2#@GK3_IZ93I=KM]
Tf+FY4BcY9f/M0dX7HT9EFCTZNJICO/.#O(Y9^J;?CSBQ)5/?Dg@,)12-OB,R;1^
.>A+dRW@EJ+@]LU_8#_NQ5T/C^/PMEg4fG0d@#R8[2#69B7Y^7/)MYX3b?81G@^H
@HdFYYYN[@H;YIS7;\21WP_(XG#d1>Q\;P@[?g\>U]J@CG51B&=DA;>(89^C5KXV
.5.Q6^XH.e4Q=[HcU7+8eDRVG+EVLf+,e\aEc?AZ(d7&X)d.]HEVWO_-&;N9ZgD=
OV]ZPLUa0Rf7B9=[:d0/cQc\UF@)0#K?DWH8_?D(JZUe#O+9Zb=E(,E-If?S&Pda
2J?-g-2<V7<K._UbG6<cCE6Ob6X0,VS(5S\J>OS/Gb6,HJdO9X/Q#6<?)HaUV#?+
A/D94M:0K&QbQC(cE15/b@a#7C_fZaf34Q++9-_309H>[F-f._G3TMO,eP@HdW.W
6;34I=.)8+\I>d7?(+P2I(>CKKT4:ZdCH5>NaVMGAN60ce_S:>>N<-QgZIaP7FVQ
DP7M,,KG@X,+JRB<dD\e4WSgVP&8@T]Qce1U5<41J[?)//NC+QZ&EBY^^4GOCE.D
GeBHC,?(N(Y\Eb,ES)2)G0(-UIWPN<6S[/a7#X@/)Hd52,/ETfUfb-N_H1]f7P9e
>7DB>GWRbEbCgbEU:8;D(F_>f&LUS9LT\=63_2b2?U.-\)BJ_FBK#+V20D.dS]f3
UAX36KMf_^GbN11-+Ug:Ia33?-\R:aa00X&K0R.)M2#eB<EW4Sc7Gg2^)[,F?],P
BB2-PTO:+dRW+T_IX+D1J#AL_O,.?-44.&V;[#DU/.UB0@P[,Y#O2+R;#2(d\f3N
7+87[:+VVcQfHdTc2@E^R7\Ua:QWZ^O_OL95QM(1.HE7H-E:c1X:K([:J5\TEP0P
Qf#XU[DJ_DS<d\(H\<=X[/L1+JJ+-R[G.[.Y7CH)2YY^2dZJ]Ug7eb[7ON3(HgId
FfP?f@g^Q?&1]?dNf&c19Z=Q5d1_6eGZR=[JTc(KA=SWd)eG8f8SCG8b?BQ?c7Ba
M0Cd]d6V9_[,JVXW-U&fH/^K=W7HO:53)6Q0[T0=JK16;WfE\^\2@L_Z3&0bH2a?
@H2:CF-88e&K2]ADN]ZLCPAO<P)JQ#Bg/,C+:@PNf,YQ/:C,F4V]gQ7O-(+@;gC2
7:d3;VO/.L?D>+;J0KI28)#>e)9[@YXPI[bWe?S3cC^7VS\99[Q^g7MUOL5[bR+:
&^&Hf-3[bT-,]9)A/;YT9MKJ(2gcP@#P/\/YYAKWEW/=A6(]_^M[#\6<6C;a@I8<
CIR0:11(@#(?c0QJ>E<Y3UZb38)+43621@MO-JS=H8X_a.YZ#S5:7-@.:JcLH;dd
:&E/N^AbYWc/E1LgY@CgDLY_44YT]X[&c1EFfC,.df5D\/CdBY[bV&QE2&ag#XJ8
?.[gJOQdJB^<[-dW7-^UcH2c^#;:WcZSSMYWPZ6e-BWZ..5-0EIFT=P,UKP_#K<2
:V@P@)^5?=_G@<ggP)6Kd(K-W@FPDMSFY.@<=J?/5KF&4:cS-IR]4O3=JQ.4Z,:+
RMM1WK=7EKM+g&BHFO>/b>ML57MXSg(<@3R2YQ+]I90R6[;03cgPdT3CST]:@BF_
C03Zg\<DVW[X-;?\S9Q&)2N0.b[#U=E2YEYc2YR7C/<4-Y0LdX+Q6/7]_dTbe3ZX
9F/H0Z,;-#VE(AQKfJ.)C,PbUfIR5(g,;U@>C[ccZVY2HOV=ORAJR3Ae)3QRQa;X
b1DO>^PO)BH8AV[V4-]b?=-]&OQDK@gD;:gR1[(KF[Se[L4/B03[L2geO&REC/aA
98fEB.G,/aEZR7OVFg7AX(M(eX5WZE^XLcC7O&CR?8<fdVd0_PDYYdNc>e,P22\1
#G.O#9&c(CO2a37X8gFBY\WAHW3ba\>\Y2[M6>0[J_<ZfA+?X>ACO?K:H)dECG@1
CRM]61K>e2=dM-<FbPSNE5RCaSLb[g4&5+M3WU,0R;2UAW[A@>T_D5:g77)+XEae
Y1#e,&fPc3QRHKSAMQ7Ae+]L@J#\4>B/X<^+L[N0)AcRgD:-FJA)M[]FL<&+@E7J
db[9Z\BJ6U\Ya/ROVNN;^R&-Fa+&]BHfMASHH\aFW.g9;O)37:&Tab:L6A;;O=f.
]6_:&J39D+fD#]MB.5.;HffR?W3_31B]T_3XK)KSL&,<:W)=L@KTBSI+deDA5<T#
IKTfIO40ea8F,PCQ-dUP5K-b1JP+VbA9UdRV_7:aD;E=D+dX-\.:HC6I6:9K;KgU
IG>eB?UP\3<0+\<BPW]O1KcL?VOJfV\5g.8;;C[IOf\IK<9@K95VH0M[Ub[>#5L(
UGN_XbJ(A.O1LELgZNc2EPfe^8:f5NTMbJOI=.Vg)>9[(^:-IQg\+a)7ddf;CFaT
gS#I[@=R8B6.\>5bFUH^5Z9T:PGH^\3L[aW)9_8-8SNV/.0YJW)[5A]eCJDR6V(-
b;1]6I#5MRc]9&:U4_7QQd[_ggEKRE<_T?b6b;&Z0Y#G_._MIdDUSA_>WRK_]_6W
>Jc^C<>c8.8+_LHTWQbR:68<,V#QEfPDMK<>0VTKe;XHN5gNQZ7PcLC\^-8_DP45
G/4OfIVHGLM/=)fKd:?EH3_g6(GODf/H_CY_5dJ#,J[0<?F0QgcE\WUQP8Z[57/:
QDM#e^Q+F#b9gZ+YdY+0J5T_T_g1e5>dE8?R).D_=GK=6dFf?@>Q\1ZKD&;<T2<6
IYb<L;K3dEQN[?I.62-H^-.BS\))1?Ub+1NVJ3>Ke0&ASZHgfF)F#;JXYCOR;V0T
c3[=\RA2>S3B2G_&([-;cA0cOdC:^0c&/eUHZ^J=bI>.cA..be0Ab=e63GX_#PF8
>D:,#:M68;C:R)eNc+I?X]BFSN]=U4LD3RNLUY[3bS;T.3.1((6(@RMd4Z4eN^U>
eW^QQ;17_/FFQDU&^K6E^4fZ;01_HH)#IFS\,QEM><TP81A:<-<K\\AdHGY4>C/R
QSZ8&N6T6+Q=Y.B4[L@P1I3GYF:0YIG@<-M5F)XPTe]g,B7IN4?LX[d^#MO@:g?X
V:F;e.G-MedH1a:&8dOP:BAVHRZG3?L+?@@PXI:F9\04(9X-H:cGI7(7)I?:H<J\
@f0dE=SA&EfXc2MI?R-ONX=Kd#cK9#,UDD-eUECe\6T7ITYa+53BS9J@[PT_eKf-
BDef_[0adf(b3,-6E&2b2)_5(?_b]3245eILd<Sf+KQaZ&TQ=_U-0AWZd#\72f48
BGe:^HLDBC(d\<0D38d#6TBJF#)N<I4OSL2/4_I3>gQKK2aK\O(\dM,);S97cO7N
#\2+<JQb1C(a=Y]0Na>/56;Ya<YOW-eTeJ\233;JP1=X?Y]^KeeJ/T5U:&<X5I=I
:DA2\G=IS0/7:V4BEJ;H?5E/T/RAS-52JD._fZ?FUK5=8UfN(Kc18F(=(#NM,AAC
X<GSW]0UN_YP5GN(36WC.;&QS,7c1DVRYTcXU6_^\>eO?WBS;\Id-d1QMRERYE=?
:LSa9Ga55S[04?gX,-#T8/)EdL9X>dJg=V;]?];/@I]CJCOKg\<K0Obf&D:.;Dd-
+4D,6a=>:9I<PIEV+EQZJL(I^.b3gMIUWURe1K?UZL\PGd[1/(Qf(@[<[)4:S^Ma
#BMNM7gNRe5>X@PE[LA^X<T,)fU]J/ad:W+.&DX6gI9\8?Z\RR;;99M^[:aTc98;
NAdJM#8T#I7FV761NY-2+KfgBI.W3MO35M+S8Z+XC2WgAHSbg02J>]KG3dT)M,_[
]54&b:3<2[c#.cVR3C;B_Web)G9=7&)U]8U35.-AGa&a7FO_J13M6Lc/.7QP(BFS
E?=M@&fg\R:?bCVccH=8ES=fV3P]/SA\@Yg&/K?cfe(Za7-Sf[KFcd1O+?>^b3e4
S^&(Nc(W\QG27ef6CbWL;R=ZU]S22(dFaMQ;@3HQeZH[7IYQ[<24=GGB55IaCA+#
]-ANW^710129169TdeGbN0e+@OF,UXGNOUdA:\NF\U;93&(ZK=(R,M8U+:g\.NN^
+bW=+A[X^OW:/#=eeDfM8N(2,\0:W[eTfTEEfRTZ0(])4&B0^^Fb-04B>#WWdad8
45GZ,G,ZXO01]FGE5852GB+>U2a6XXYO.MbU0eN@52PXa?84/_bJ;248dU0RH)WA
Sbb;<W),fd4,DB&;.E&b6b_YA,-TWKVGHEWAe1^KG_5)bQ+ZYH_;N\ff3[Kfd+MU
Z(.S\bCR.Cf>XZ[4YR3N=gPd0-H]#S6aM8G?a6E4M6HH-;NQNU_3M/Nc8ML_\4Q)
Nd74I:;]fC(FTBT02:25c2Ub7:5:eXSF,TH2)QKF>N3FR7@-FaS=1&eDfXCIY5#e
W..PZd7L22J(dUg)U1_M#P-^1.-M0DVfCC84^@Nba?X5b13#BU+Rd<:L86bJJJ3\
W>6Rg2[ZLgB;bbRLJ.-<G__)JReGg]c@Z1_/N;;>D2JFB&F2D,D]>@a2debEVU/O
#>A5N;BPZH)aUO7G3C6W4V)QIBP#aKH.E5.>N/-3&cU\EbF?_e:[S;T[<BTGJ?2)
4:7aA4+2G<9&5958.ZV<E1Y9eY#Z76BfS&^>JCUBONL1>[T#S+8)YV6b;+76GR,S
WdIO<C)Y@255LVJHdUS;=5U8;SI;[-4b?D:71F4X4-XNgc4Z:FZ6YbPE4c[aEGVI
X..c?(gBC5YZ56KZET@HF;E-I6IaD^gV5eeH+PS5HLFFXbH7<bOZP2IKOELSI_;I
WF(X6GNXFdC-8Mf3928d;IT^_;1NM-K6XbZeGA6<XT?g&1)N+@F<?1DV5aR_>80J
56IE.[OZ;Y/A^#K+b/A>N3Ce;ME4I3\(fO=1LU^.bHNU0C2.ETLJgGAJN1#N\TXQ
UaWc-)L(4<>(YKfH7U@[9NKXP<>RZ#]]SJ<:bD5]^TP=QWgBT]V0AF@RI2.22ECX
[[XCANfRB=;4#eVEIbLPcY7,9C0)[Ug^TX]/XKP8II@dM\/eSLA=b\gFYAYMdfcT
X<#A^LY[?Z6D5Z/P&YTcPTC3)[B/UC&2T;\Bc]0<XD_[VE>KT7YRQ04b2-W##&D1
;[4-:eQMB91;MN)TaXX63)7X45S2P<CZ;d14_3Q3J2).,^=5EEeQLc2c<_5[d;GE
>M]0OJ[f11bca?2XK]9H^7])-/E#=8,<8EYK&5Y=\S.\L=8VCP3RL).(PGaYcN@g
#.WI@cCQQC1X7?,+F.U^;RWKLU],DXK[LK8_gC&.VAXEf#_ZFd&_Y,-E5=SMUf39
#4,.57##/HW-?B50N\\W;3//dF-D;PHY-OXA=EZ37]>5U:g9;Jb^1V)#8W#&eZgC
P2N=@&ge6/Y5a2&Z>KbUQK&=CRXCYB(4U4g\42WP?fW1d+cR[;R;;UXNMI=N@;B_
7LT+/]aG^UK?aJf<(PULWZ@O6;XC@bCCb0AGS#d\2KVAd/MN>V7gF3UO[/K5X?O(
A[<ID/cX9:BB.IQ/>aKOE48(=4T?A&Ab#V-BIPe;F\M/a(-d#8UUOMJ<KGU.P,F2
.LYZ&d9MM3#=NU,4VB\:FO32&L[AOU.+dacU/)g/@MF4-=?eb92FL(,CEL<6S81c
NT./:I6O,58X=FH9E/a79)XEaIITPB=TS9FS[([29/>-PLS]bOG,FKXG^/K4#RK8
JA^26e576A^IOK9;P#@#Y0-U8d1(OINaZ)^1TDCg+Kg@bT@g4Y5.R(>1J3:=AR87
4#.@[4L@9Pa_C)J-64c++,RPQ3f5,Ja=QXE5.YUR24/9LK#)X?5E9<F&QRfUA(KO
b@Id)5NWAT@8dUL.4aN.(RHXWBK\4_5\R05&^TB=2+>_O+YRa.b-W7;]8;C^,5O[
OeM>FV>ESN]g=22_.??Mb^R&#G5b@\4DK4Z/<YJSb7a9EIDdaU&[8CA.fOKKFA8X
@I?##ZL;4XZ<eX<A4a00_HF@6=3/e-]JDN&-DST]b89(Rgg0Q/fIO;1Hg2)Z>A\8
=VN#K&4Hf_9<(<a/bZI);K/4.2,a@\2Ig0\-.G5PQOAS(CZ86OHEa:fP&17)Y]K@
S2?2YB:(=6]bPC[PAd#g[P]+[aUZIF><cLR43KV?Y\8#KYV@.cXb^\++RT?fbHEK
a/HO.&eY+0?e4;LRd<#.XDYV<TY6AaY(eda8BO0QbAQSZ&CG.>4=A@AC>+VdEc5J
)=P2T.SZUeAG:O47.0CY,G2/??U(8)@Z+/;b(3\9Se8VL+D4CN&\3NgNL>1\/T-_
L7D/Ed20@)gFZIUa].;.:R)\bI8B<:(JKbd.6]L#1g)O?J/eLHOAX;@dEN76F20^
-F9UZN[:NR<f,BIQJV;ML.4ICWS72HeNT))O/f^.#,>BSB@.@#a[+35?;b>N.B^P
E[<<LZL.KfJc-B.J2:XdR/_^AN]HP/a\B/:+N##NOOW^G>AQ/C(_U8J9@:<J-FX4
(:>BTVR)Z<<8_Z0MUT7X2dPJX#[FS(>7C@D_C(\,eRB=VX)CAFJ&S5IE]U?]dL::
]A&1]&dIE2FY3WB5<4[2M\PS:RcMV]XXJH04M?KZM#_,[>H(abKM/:AC-c\:QK-A
7g[S=;-X;.^_(OWP5-ADQKJf#KSObVaG<QIFH:-][T)K9R;5;1aC[WCZH&:/Of?(
L_83d5L0HXbH[SE(&,TA]\+<;8aDgNQ7^NV@7c>ZJ;3cb,TL&]4(FR#0C<,@X<0)
N5cGUS>\2OX42ZdHWc.M_Q4SR;_>C35YZ^Q(S6DX3bA^\_Q81ZLBLbD)cYfT5Pb;
@fWM4FI?AKV3Q&d8K<TM^U-J6NedWTPbg5ITa)ce,BXUIKZ9LPK4;1R2cG9T=^0+
M.?bSJ&D5,EWI:W.P\XM.,\OQaYP<Z1:T8bTZG0:gN&,6MXS1R=(1_UZUYXO=_)4
2ARF3ae]>3B[fLT87fN7/PAXL9E80Mg+Z8gV/M2R^-/VS3+Y.)#&(.\T3E\S<D[Q
BfVR>M,<5P/+dFWKdcN?02:fK(:UUJ(-7^G[)BV+<2b0Q@2]MLCE47e38--9:MDe
F?<QW_<2XN/J(c0\<:bL43EP;#\=\?=]DA]_:\)76.@efC&c1JAg/9^;;8SR>?A5
K4(6:)JA4+&g0F:XON;_FFI]<^bZ(F(f:OOXRU)<JHf2.g9/7CR9YXEf[9CEZS9=
4dbTC\#6:ZW+UJC=523Ja@<)G?CM721MadY:C(YI5UfZ5V_[WN5-G87WbbL^\GaV
.^82=CX-/4MOT_Wb9XE,S+BTd3bY,F&4AG?Z<DD(bS[##(1Sb.T>>WQ7f,d3Xd#1
:f]<+BO5JMS3eG3c]fL7:Wfe7=TDCU3]c@]GX67IFFT(X0-YQPCH4KT7ZT5X18#e
2>RMTE?X2?>9(W,6;bDNDA,#0<b>eHZBYRUS:P#=QfWGUAcXGJGJ[RDP0&X8^9U,
d9U:Vc3)0#BeV[:1L#<Y\A8WG>W#R&[c,=a_;(7I?@bBU([-^_1a_IXT1L8MD1Yf
f(2C_K+UEPeGE]QK5>=UILJPIJYFcLbV-Lf_,Lf)7f15Nc4(69XZ255Zd_L8gH0X
]dOF_LYPUVEA,U_eP-dW./Zc0@3-./g.UNM2I^W2?>=PQB07W0IXC5-Z60K3DBPT
:9;FfW)cKdPFH3YO5BNgELcM.Y41[<.0b3G.GHT9AV96<11D<db_=Oce;S3HU=_f
FW9EAW#C_=B^LI,UMR(>]0]]+.=DF^FICZ2LXHa;WO](#P[+0..);I5+YLZP97J_
GHMIg>MMUG3X?fcP.bD]=>BD@/D=EgP_ATGDU[47\E)4F..(4@82DeEd3;IZ3CL4
:1_\49T)H)V96:Lc(?_KPQ&de[62=B886#.K,-Q^3(8^(YPH8gR(YPJINL\,+_\,
1:S&(Z>P6?<#Qc[K3K#CGQUP5<F4EWRL6,_0#^O0O@;ITT+KSMI1W.[#65fbg^Z9
GG=ObeaXbAY]V9:Q3f0O>?.3NFGBV,0dP#[FaIP&-JPEdNF^HNJ/dY6#L+FICDaZ
K:,F?]=P9\(0.^@M]0+79<E^+A&4/AM.#XV<#;(A]W(897Ucb/97N-8b;Z]=1WL6
G5E6;;2?Z?O@40[Pa]eaHJ3,2QFW6NI(8XO;#EV7D,VTX<aN-f0=5KPE+X.ID.gE
O3D=aZO30VFXQ+Z&RD(>3f3MA(cG4T51PaA?A+H>P4,KE;F0WB&,5TIH+Y(UcXcI
,0KM7TNL#SZVG6D.A/A;+d35Fc.TNRWUbM6D(0O46JXSUV0^QSE[..<@0^,)9-=H
dV;aC:5]&[J(7YN#LbTfAHYEbX^RRg7_7O/N)T=AK/G(63G-Hc\aZR&LX/;=X;e.
&:dcZ&[GgBK+0AUb0I&JDW&4T9Ibd75J6)J2VU-1;1--9HPFb0DM<[<:c9:Y,G:#
1@Aa8PI]/Na4:\8F070?GKE=?TCU;]P\fOSZ=[P.ad^.-)+1(5R/63->SK?VH.,U
)OS:TY(9(bR78bUc)Y:UXZ@,L@^1VL0S@VA@4If5cYW=Wf(c.(\]Gb.15EZc=XaV
2Z_JJKC^JNFP^YUL+O4U6:G,TXB=JZ>L?-Y=NJ/c[Ig-J1UNHd+HN,f8&MRAJ,gI
T>0&:;b7/+,#dOZR&/-<E]<9D:O066.eY,/BdP]3Fd=1e8PU=(X>,&/O:_B3IO75
EI/?IgPEa1Ha,0Z^@=[b19+Z^(7^_>JGY;_g[Le,2PTaFGbc9U/5eO77@-0dFB-8
8NC0/>R,?dg:>>MO_]^A1F[SP/9JS(WGW(T]_QW>>e.>O?[b(,0CDdb\:#N\YAgP
?)EHSV5&IS-7b(XW-b#HSU?WQ4#PG@c_>:?U6;25Qc/_2<H2]+\05GCB/3gQBVVb
;I.N;gTWBSOCMBEeY\&.FJ:][WYfXS^0W2TVf+Xe7gL:TV:.L#OBfg(ZF8c3@_@+
DN6PGNX4JGI^N#/P<J&LTf)Z(Yg^.J;gYbe\Y/&O7d<B/]g^RBaG@>?T(ga96-5Z
HP5ZZMAe0T,:N8/JBDZa^N+F<7&S?D\C@92bf12cQOHT(7^[DT0M6+K(4_DH?.Z;
eYUd\Y56XI@F6D6#IM+4M4>K5M(M=geA-Q>6.+M\B_Y1#+fDOgeQ^^Y,?IM90N72
OKH:8/\[#:FEfB_R;TRV<8A,D;Se#-gf=GO1B-EMfd/a-5O0=N)NCCR[Kg9AVS[a
D82QUbEU69Q6/+YdG\M:fL4P;G6_9@0P+Q]8U18^,(@USZWL&=(W3SW7,=S2M:Kc
+c@T5)QT5b/4GANb8;C:X,23H7-c\e2U[\COfGO\:K=XRF9+b]?A;aUBK^2<IP.E
GJQ:.32YX,D@._1BL<WN82KZLUGDTBFJ5(6,cRIbgLe^BX^FO4686fMJ^Y\fF]a^
?dWZH@NU6-&L4Y<STKDD/-(X0+(0aagHJFbZ,7^HBVWD]@@eUG(K/<1fb?F5g9,T
2H5c+M.a@V7>/?D[LVX4SYbE>+/H[_>,#:)S<:W?5[4B/31XaFV^:;#[);N]aeEN
#=IS02Hg^Y@4?G,^_0cb.aVb6A0Q(3(Mg/g5=GA:+QdP/TE/96Y3)\<eA,2](6GW
?&KcWdX(<IDHde9[e&O^=1H>T&WIBNe1Rf3;Cb;VN?7@>K#.-JVNf<DM2Q^.SD,A
SQTd3\1<7VPf^VPX3H\>HFU:TB(Q]EGIL?7Ie2Z5<F[8O8UB_adF<[7>J1a&ZLIU
bS-9Jb06V)UW)@4:b((g;S;8Q69TfV\cBU&GS-CZZdN?#>&[@e_H()[&O#B6D?;]
QCW#/?g&e,06-PN)_-SNP35P9b-1W7TTO#3.b&F<cI&/2#+8C>=Z+H[[ZNZTL9BO
Y:cM9T>PUOY,KO)bE7LAIQ-M6e=(fd#A:fM<18Y[IQ-4VK-a##OHIP6A1J=[W3N?
(SM6bW1Z?7GDV5.@K64Y/,0,8@-A[<F#5:VN4Hf5NMT&8b.\5@@E=1L(7WeXHb#Y
4e18JQ3-G7N#7QO7b0:VF#B?\_KKb(N]<Z=,65]?G_b&Qb,FRJ[Z&\\H;T_^&?BM
Fd-6;I]5SRAc8c(8TD;Q&f)44b(GNG7c/3S#ZSOJU7_==LNUU7f,XWF\b3f^W@b<
RNC645.Q7]-P[LCF?M(OPBWVVD[V#<6I\6[00,>]Z^BA?M[N7a]a=DH,2)L0>7Kd
2:?8M2?OEWD>_1?HC847,CIY:Q)0SVIGJ5Yf1XMN#.OgAcQ?3^34d:PR:SdEJQA-
R.4ZFX\8T,N.0Lg7GfV2CJ3R<7GC(G<5#]RW1Mc[4()OGUZGQb#3_/D2V#dbR5=X
#54RM94H2:(cLKJ4CU4d7UbB.T;I50,8.a7>[ec1/0VJ.\Hg=]X\5gHH6++.O>)C
B;d+B/^G_G96Ygeg<ZQaWKZ_6Z\#;QFTXTGa+c>HJ^aPT;-JROXZ4K_Q?]AL(VE[
+<0X(ZC&[;f,ZEcg?8,D6d;NL\II.U@b7dLg,e0)W4VadFS^Xd9_H_ce:G<)=:LM
R0O_L.--?BaZE849B9N)fg7+>FfaUC>FBDZPY;O+-cKVH?0]FJZ@LHeb7W#>+V-^
G(G66[BL\Y<M),gG_NXJ4,^)Y9T=dd[>P&A+R<;248KQ(MDG8&GBC?fI=>9HeCZ:
7GcU+M_22HQ>R<P+V>3D]6[MX\;\1]@d5+&.KTd-6X?;,6DEJ0/MHBYOM93A9?fO
I.ZTZ;,&e02)<C[fCZ)3/77c9I]#W66G-G\>>O/R3Uc/.@U2LbNA:&H98BH;c3@Y
&6^OA:4EX>,O2\cXH>&AFb:B+.RZ91bR4ed/#>GJYQF>Rd](VMAa[YL.UFZf0de<
/<92gWD#.4?].+?1d8ZTd6],F@B6/+3-GP54V#V.aE)44@8_<,XM/7J;FD?HSH5Q
c33fLJ:=]@b@[L935/-9,UVc;KT#G+JVSRWF=d_d_+_g.O];W.:a,DZ-J[<MS,P(
.[<N>DV#LL6-Vf]C.aMHbL((Q&PWUL:RVdB3R=C)7NZAML]>?HQA82@I(QX0BQ7N
gaUDM(O^b.H/L1dH^5WN7f_X+3#64H.B8JK<L0-F:-/<_g<eIH[AG:T6:\df@KV3
c@fEd1A;A/:8.ZP?eB(-Q#X9SG8?P9Cd[L(8]RMC9BT8^:[>MEe7RU(c@f9X/^MC
<#A8RVNf@F@_Q8P\4B[:XR3-/YK&.@]713D:A1(JITS..:+FPfSS4R?f8#1/d91I
b8MA.@JM;MH3CK[aa[Of)g;8LTK&.Z3Ve14)C?&0^URKZ7fcaga>Q5</4>c,I.E?
EfG0SNc0(6/QM8:E-&<&Z>N61.P(B-[,f__#.Q36A:WEYe]DAOL)Zc7>-I-6DSI(
-E9FM6://T;&LGG(5ZB44cAPLH4@.CU0D9YB/&:b[T9C8;D\e_@f<Xe.6GF-[66[
:D_<@X/d.P3#>cbZ@V0b;e]JfW(I<9e.]Ucg[;@R0BYUF_fc/DF@c1(T&64EV&V=
I-37CM<6_C5LTPJSA6]?a6F+(7>f/[N++Q.E:FSW>_/8&ZQ[XQFFJBA5#WX<2fb_
gRADRJE#fe4YEc6VgDK&KY9)d&@?.&Sd[+[RB/-CcM3N<.UeRI[H\=]Y<5e_/I.B
+PQ?Z3YN81f+f,.>7FLQ(4-NSWVL(YOOccSJSFEI1b=g_NS/DCa5U00cN@GbXb6A
\[6QFRBafdYAe@3-b1GY>G5dV6&9,&.)/=+:JAUf:;0&]9\7.XZ^)#0POJe/H7W8
P=R.RKa(U7@B+;88g^-P<OPS&Z@FGE630dddDC#AAbTf5ENE>ZGO&,#&869Be35#
+9KM&]bP/Y,X.2S+eXM,/6WURK&G7=#:K?d/)cIC(cER>@)R;([R7G,LNa600C_0
QU@6-MJSI\>>:P#8U8^IH#CPADcO7fFZd_++1:+HRdM[WD?K1>SDVG8PDJ5RS;_C
X:<J(.6N?Hb?.;A,44bf)Ud83T>AE9[6E8II,,2).5]/]F1/])XC9\XWa?<SZ3TY
/Mb3@)8#RDG##gDa+.O/F2Xg11.Z\f>F@IQFVWDVL:9X<0E/P)=O:F]g9[Pb+DBY
0:f8SX5D;a1KbPNZS\9bDg>YF>HUME?<.R#V]\QCL86P_L30^NLF<AHgJ(@W,<D]
WB(]WfW5T>J?D7OE#^dcZKXK>,TR#().,6b[N4MVbHbdIa&[,)ADfEg8JYcg-fA.
cb83[)eb<MDAgLRUeS,^MDBUC?1MV-A8cEf^L<CeCB4N/)@5:A1.c)be1+bM?2b^
WZcI)JJL_Y#Hg[;/AR5].@/>Q?+eLG2?&>?#K;7g\aS8^SFR^58JA2C)?<fBg.c3
96Ng5HH:J>YR[(IGRb9S?e0CHdQ-Ea6N..<(f4\I)^>WZ64\63^,W_VOCdS-)HTb
O>@0V5E)+1/I3..+3f9#f:2AE^f@6(bRQ?W)7PCAU6SARXWXK/_?BX0,[14GRVIQ
J<Jd)TXL_E<R_2]bbT=9@1TKHBB,,gaP5RL7/,=.FH4@Y(Y-:.\X^AC7UP2,EIT?
UH0G9)K_:He+C&)OZff9^N&\(C>M8T1\a4Zd]6K@XJ-4AOZ,K8/11+a?eP/@dT\-
=DT;6.DHLOZTQ<^,c&82P)2MEMX6)b27-@RH9^cX(^Vb9/f=[J6ecfeKJIS;Mca3
>>K[1LgXUH5GQEaOX[-B0/A(^Y<#):9_[_6]>(,VYfMW2A7RcA)7V.O(A90#Y4]M
_VC5<2B[.(.dH#6#QDQ=->g_MA[Zcc961]\QEf\LU.;?E+LV=45,<5/\FN.N8ED=
@;28?5]@d4K.U3H.;.9HOG,ad99/1+^;06L.dO[::fYUZ,d8+FOV>\IENAMEU8/e
+\.2\f>+&ORQ>\aU_N,0H3?)PF^ffPeF[H5b_&K^5=J)^ND1=>2g2Y6L5@CU4Cg0
^[IB05cQ.Uc5?XXMeL>R2T+^KZ/Fe46G_Q@O\:SWRgF&E[_6^7b--44Sc9AaN0S9
_KAd?&YO#HfKG)Vg0Y=8[B;D<[..-O\a?&#1R?2^QbXcE1XAIF#FB9GC+18+@e5?
2.VZ1&:K7FM-.11We/Z0G?YgFae#;UGYR,b[ZSQMc0\^KF,Pc:ZCUgL&(BC6cPMC
:\B=7TeL?F_4)6&SG,dbR(2KW\b<Z88@8G0N.>5J0Z2Y7XPIK6YGA6H:&&M^@.MI
dQPa&G+4#^RCQeVS=5g-0XWH\=H<eM[_;)SJ?O@C[dSgfFBH)2g&2Z:g.TQ4f9A@
We[VC5W&S64dgeTVNF.F,OY=4N;g17)BOG>R&RG85U>:OSV72#GVEb9.]I_P+;BD
7FHY.J;9>5F[<-FKe>)cdWdR<]/8&&ADK+P8V.UcT4-8[Uc=B5<d^)-/(I+MJ^AF
QBEPc--QBBDJ=:(@e+V8QZA)O.DUdc=Ia:_>0ZQ_LH,]YG2)d619ID[G[?a(DA62
\>b<T?]()H.<LeSf/RPMg\(:N9+_@DACL<L/+US_RE?IN=NU+JE?.1?EKDa]UL&:
&<Kd&KK:0bHF2Ff9:C(<b\-:KHF;OOfFE<Q,Xac.XC-_2e-F:f8TDL<4]GTT,GE4
F3dUEBO45+13?:1e5<E5;X2@]EYJYEKR096df>OgXLZ0^A:NUD9XRb]Zae7+9<D>
/(_QKECK:]+Nf1N,@O40TE]BH0:GH8#)P;ID61ER8><+[ROEF)>CAJU@J+ZP/EH[
;\E+J3RIDV_SF0LD,L9Y<1gIcN;\b#WU?1I&;M+LT3=L=SZ0=g1LVX_(NM_(AHQ&
6-g4d+Mg@=72FQE/g,_F.BbaJWF[,A)QI>Zf=T78?bSWF&P\2Mc2T6?_UU9M-V9(
C3b^^<(NVb(&X,Ifdd)VO^8,VXU[d9;(0=)\?BOPXf>96L5@LKBF(:T:bNP)-316
>75GTB#:\=/13dJ;B=IVAd(W^/L#P1c2U8M6&a@cK?V(/MCIHF8L(XBM6,?99OS9
Y[JQZS6OQ61bRK;J>A0ABG.c,9.5)_-HaPd+d^4Q2\?11:_T0R_S75&(SB.6=M\(
cX#L_6([07#)aON0EO:5V[HQF_S4KO?14,;6LIMDS((D+bL/WbWRPb.AJ0K0ca#X
OKC#B5?bW9FX)[/=@9,^KgP.XdXL<:Wf@\K9A;PUFc9MaLJ-;/^PK?AB7W0JO(9K
fBYe;CZ((B&JSAf,H]=d/EMa2fGQJOXPSRc2^_GE@V_g<a05X4UcTU/S([T+Q>67
6]K./e3<1=g[V;L(\^,fF0-_DTB6fH<Hc<?^2&5G-5O#8)U(4LH3^JU&a=,]gZ2W
,Pfg[5NSD/LO1L-N>+Q1-0e3QK2@.J8>U&(J;3gWd[21&3[DaANfU2;U9^/fFcJ7
b>D_@IDWa\>7#KR#72G<<Zf4_dRA:S4>.H@,PL=IVMTA[AaY97X_5^A@9/J+QXCY
/.^&NY9Q-L7EWU&a(87L,8..-65)WJ@:c7G#OUWN2&YSGcV^T=WDPN+J;^Q1>[^e
.2J1(G.\AFd\@:e1KZ&0(Y/aL+5c.II-KMHeW3B1ZM6TE-ScM0/2DIF/JD(\]g&W
,Ka=S;D1/&0MQbO(Xfg11XXL^Q\/8](NA,f)fdEGKPA&+I265/9L;fNE4.@?#OcZ
dV6YS8F:?^2Cc/4;#2THI7?\eeJ1=DYe&M-1XM7[(Ta8YbW/)G?U8S;1=:?8aHE=
9V,A-YKPN+]2Tde]5+TX;0\4ScYAHG^.]6_9-M:ZJ&K]JVM-8(41Bf0LQMdKES\a
;JEO\=NU+GL#e7BN-&H.PgCfW9fPbW&JA?B<@a&C8A3./,U@RV,bVdO#XD@]R;.f
fc7YD?(5XZ/IM6^CVX3[Q;[97W3fMe-D)g?5Q84HW;YgLc4MF3I+.+5aRBO,=H81
.1G,/8W)3)cJZ</@3f02b]a^_ag?<^4_7(JSKeOUG9_6=M]N,EW59-;C95>\_3IN
=4(<dZDO))_HP[_V&ESD6a(4&075@e;E=KZ-+cS3GUEb3@-;3_/&3=O5W-/])BJF
/OaR1^F6FGE,&FT71A:aHCUI[GL/LaDd(6UJ@#L:IZ^AV2Z1g+<NU)[W(5U)b9QR
-M-)g2X3N/9M7I_a[S,&,D[Ad0GW&d>dNg+2Md?DaP/,d[=CR&^QIRZR568X(A2J
>D;+GJ.,PXeK:KXA(L+-:X-?R1-QA;S[^P&>a9D4Ud=YNEK_[G/G?\ZaTY(J35HH
V=OMcbFYMX.@eA42C<7?ITc#+8e)bF\46&B](6XS)b?4&JHVL]Xeb@^9C\LLZH,G
,I)7=AR^X^15DI1-c15Y\P3#cT1GCa(A)E?<L(RZF3]dI^C4W8L].0-LJ5)Q+,KW
ZBE80H&c9?1eE@G];6_(+J?MRT\2C:a::3M<6#5>c6Z5ScG0P4UOUU:RVER:]+7F
>&&?5:L//HOR_eUR@&=A@)?/,,7,1HIRd_EAG3+a>@fX]A+073Z/T^5Cc)2XR;S&
9WIbFEC@J:S/0IZR5Da3\?X]W\ELNgWESZE7NgfXgOaQKZ?d.N)4-U\QBYQVd0.H
KJ&+Z2gKJK2@43]DL1^S65M3O/^Y+IO4IaT)Q#g2C)cg_=,Y+YPG7e@Y0JV-b=-F
)ccYDKK,-IU3W7NC,B6JP:3VJ2]PE0KNSbZM0F3Q7Ka6KL]30F\G9/Gaa@2EH(IH
GOSV(C.:YEcR\-gV6]D:T7JT=d&9-=(WJ(8ICTaPU=F7HYc-)+F^]-J>BZ.-<#3C
-DHcOV7F>JeEXN<^8\Fd)MK-73dMUfgF.bH/Z8O1Hg&_e3[e7Ac:3g+9//XPO35<
C]F]RAA11^3?)d(W3.Z1,?/:#eKbTJ>;/ITLIK7,I&:=VJ_ZD..(5TdBP.]3YVWC
a+UQ=;;77_<I+.6/#5A<J#B[?&=V.&G9&9>f2:MZ;@gMH,?Rf@[^IXbHR309begg
L5A#&_2RYQ3,<G1B5d5^GJFSfVE)SF@<(S[B=FZOAJ9K=P[a19JOe\8(LMVF?S6/
eS0FKg):Q,f2f>^PX>^UI4>C?(:DN7;LT#].[Ef2fLLSMa9#9a]-I98DZQOO@O7T
)BT@8gAIX>)RIH(XADa69\&?d;H@5E;DfIY<L;56\=0P(;<:]1X?FTZ]@-I[=<-1
M^D;OV&Je/RN2A=NU_RJU=JgVNDRE;LcJ=U,Q60-O]A?KD9fV<IIgK^fDA,_AaX[
2?#;Hf\FGS8:U-[7KTJ&6_=Ca34^cXb?HL27@d?K40AQP#+SC8:SAYPZ4Q[/31#b
WFeE1.[-G?0f\.#O:1E&LgI<VUII>[EA#>#U(18#7dME/^2Z5D\ca;3XXV=.,W;A
,P]P/TTT@Z444TDUYFT+]L94g7T7-P.FIe3ONM7f;gbb\9fWO\IXM-?(cZSJbg_9
_P.g6V_I,JJ050LbP6E=F7-MCLZO&.H^D+RNQKO^E]:_Fb^D8,)IA[@)H_JS0.-&
dV[.QOK\OUTaFF<VPScK4M==a1Pf^XQ_T;#e+M-NOSG#9@5\6+_bL&RS=\dfUK=+
ZN.fQeT<d:US_[9:/PaRXF>[UL;A?C93F+^C@LF]S+&QY^2e^CI[f\,4aeL+Qa21
[.2^d#,NU9)>D<ObGYR/GP9P=;P9>99YBUN>CADB+4<FI+gL:=])fb^>3-NUW\OX
SYgGBYD[3Y89BH./@.<8KF46&4-I76G/<5U6F3IagU:=U]OA:;\3]PDU(g4GLS;9
PScU7WNSSA-2:F;]#KKTM:0.@Z2[X=fEZPF7-H3BbIe,,9Qd]/9.+P(9STQ1FQ,c
A_]X/-K=aQCb5W&e?\M&+d;R]37L2f_B29a+IKb?PRLO+?\RC;a?Z1+bLQY_5H^5
@YMZ:_ZBQ0,BC5I]IJLQ+YJ24IQWD)9.43CX[L=8JJGE6)Mb5bB0PMTa].Ma>R6B
&G<SZg5I1=(QCU9)<)39MTH:OXLAaG[T)#GIY2e<YXHSg_NZD)g:KNY4X#5BV#9G
[:\=^I:e@2Lf;^I@.:P.O<_LPKKK)dNMQIa53_16B,;A)AZfTcQ)Q8gSGQW>@eQU
b\g<)(/<aE(I_FSNRNSZ>84bO-41D7d;A[b;=CC5?VZVG^2CY6PbbA1GVJ/L3WI&
#-aIY[4<a4(ZB:.:9B]<;W:;+EgHacA-JLS+dY^]7&;fFS\f&#6>9#<A+14,ecNE
@=EbS:C[X[T)F:1&^L5Q=EEU/I1#VMQ^N;<=_EWU:2N.6V7egLS3MU2G:#V.U5=c
RE=8A9V:8<FEBQN=S.VF/H=0J)\4HN,5:BTTEFF6K5>8)T]KE,fc]TN3W]+AX<3+
+0.?]KS/<T\IC>P&@+d-P=7ATKTc]=8W23R+b-@A8=/?+)65(60O=&3Kd3YXI\C+
XDLNP5DR92_I-TT&XRHPU##/CW(#6)b_J-+dC(YPbV]P[TH+dcW_\f)HE2ObHJ#N
>)V_R3<W??d?U4YG+gK42SUd&NMfc:76@D;dWOba=73,<9+K.=K&.CP[.?\Ub)6A
8O@g:<U:^DFfVLHe?029bC(,J,b)\ee^/?Pa+U6XdF3g5,_fb(WEdHI_&b+L@?Kf
3L:=L6J,YMYJNFF@F((.:Wa3I/=5@c/&b0=&J7Jc5OLNe2OMG(?/cc./#^5,HA62
.K[Mc_)F;>>+O^f@H2JTN9M]bM5GWg8@dc,(Zg@:bQ<2cee5\c4,Y.X4HW1Ng2C.
#+gA6SB<e+\e-13M(90+^(];48ML75J[e,Q3-WKaWK4Eff)6LRWgXA\Z[SZ1d#_+
+[aK9(&SKH6/THS8[)@Odf5X1F:P3=^AII7DI90W;T=U<9)\9Xc2^(/EEY2_2>DP
^)B.D.cNTb<]Re,IP4b-D[2/9;2D0=Q#7MY&=JRbLf/H9/R[ZE[YW#VS2J<Rf6;?
D;:^PJ[YfeE<O);NNQ5KgZd[=+Y5TT+LB/5<I54CC7;W(YD6dA1N&FD6@-FVQ+:9
B5.9f0P=dQ60Z<dG6O</L-6ZXYWc,0A#,B1c;R:=TN=c@WH9CSX&VZ<:GA,A_&),
#]=8_S=44HK0);@^d517596#f=\62WH3H[EBeY37MFc/Y09N6[((_9()>,T5/@fF
)TB>A6cL<c<I1Q\J5NOWdM\:Y7@3,IaD\;-;7TMW;/#R5C3d+P7Y0IcXP^bC-_f,
-G3W:c?MD9Hg-Z7bg-bE@ff)FXQeL)0FN6R182X#89=(D,2N)5;VKG,N+ZM0J25-
0Z1e@&U@E-aV++H+GD]gXWJW-S79_@]OK:G14,7#574>G(A:41L5EMVYfHa)S.Sc
\JD,TT<#Ne(AGCNA^Q.JW\4J#3UM]C39\I78\2Hc3W\[N876\;f.A+5D4^;-U-:=
3b)CbU8ZC8\,,JC<L2/[1KF6_G&F+^<)Qa&c4W=QT[Rc4@9EbgMW.3GW^U,BK;@E
ITQQS/R#T/];Z8b#R?JRL91?eRR/<A]UQc]dgTVEMKU#4Z3&O@,Y]-U3-GVb3GEO
.5L/\+DEW2O]GK\]IX<bX4cTI5VU>\3Q(P\\R1J;D+0a8JH>Y3CZK8eYgZ6g9FY)
V[H1<)bO@O8eP9PcIE-VK@1I<DMXaLQbH4CX<dJ\N23ZV5,(C5C@b?^DK.>6HZ;8
P2>-f@L;N#Z;2@2\YN9^C[-/+;#^<KNX6X9_[_)7W5eH/1J\X+c0C-&S;G#^]=b9
d)KbdH+RNQ(@8R80D?DbQSFR(FUP0?BMC_T/]]3I^EX;X-7:ZQVg:8T/69JRcdXc
?9c,Qgb4E;QC-;5ON6>=Z_Y1?\/LKT@UUHWI:;0/aB5^]c(/[);Z;9c3c3.Y+gWQ
)RR;/)d=XccM;(7)PQ,>E,)@EM+#,(L4D/F]K)+HPP9&D=UVQ>(fV\0-:gG?^c9/
CFe:P7<ZPfEX=c9VP,8R?RXJMPA:],>bV(d&0J[Uf@4gNM/f>5YEAZ.FFd[cb2ME
<^:@2IMML)CQ31EB(3-gI?)NZRPA8Eb2B[)/gd0(b5O[WB[MMG<=2#fdN9\VT^,9
b_D<ZVTECKYW9c?R7O:4T,I;D\?b8UfA]WS39c/.]PRD.91N&PA?A@&^9QUM1&Gg
78)-6?\?=8OccS\4^:<\L@X/@^Of[<?:7>1[(P&.R_SB7eZD)]#@412RO^V?(&YU
c2e-[MJH^)^2Hg#7,\ZD;aD-eaY,<8>bZ6eZb5&dS[FSfd[SSR_STd>PN5SXd?Oe
Sg;^7HG?T42Zb/^.J&T/9-KOTc8#NMB59CC2Kadg2L<>d^d?EKHMPL1<ZY@9GUO5
8S(0=e3R3YG?-;2_G:T61YMVRJEgK(2+eg23IED#>W0b8dK>2N_/d=cefRC-TFcU
b9QANTag2de<cF6/#Q=I^feX?[bD6PU0Pb1QR]VB&V0(TMW&1f8T0d\RJ2?4S;LU
SNS2A1c(>cIB:,6LM.>(O<DB:32e<BP>XY@3P3[N4<K;H8a+^g8B?^]g=D6BTIO2
Pg_U)DKYNMKT1?8\HAV6BFO>gY?5V,HOG\1Bg_\Sc<-U-JgGDCE/-^JaQ0VXG(,,
\Q>PEe\I]JS;\3:NcNT#QW6)Y3(AP[174FA-IaW>8&C<H?R7d<2V(OIc#Z2R2<Y3
6,DTA^8D,-R92PND9Q4feC7Y>)\ZEWJ]RK&_dLJ(]8gUXH>>96]Rg)JUA\UcEAbX
/M8^]fN/WI#A9J=(b9R#QS@@L5a0CM&J84+-[BP^=@dDHgB/Y^2G)/Wd=HN9d[4d
.SWOJ_@8KLf\>gggBc4\/?U^<\UD0)M<VQFL0UfI2da(=S+\U]&1[bA2T6R^J/&+
aW[0;_G:.f4]220W4\^Z\F.,S/,D>S555<(WCH.@PY:L7/<X^A43-3NJ(4:K.2eD
:GN-PBJQP,<0:#QdO9-R^Qd67Na6;a;JaP20^1VGBH\70#EZY,+@&:g].I#(,(T@
9XJ\X=K2H,[&J:f?8O&aS+c@3)Gb(+12;)5d7K<7FBLY?LT:^.DDGf_6d@I?K;JM
/:N3[\A(;+9@J&Y6c-_[6e:VBecVKgC4W-,)YR3@8]E6gJ6d>JGT&].-C:U^a22&
;:\/<II75EV80BgK:b;,1Ad\g\Tg.ea,e?6_O/C2:DT-ePSK_;M\abXF)CR=4,5I
-TO,ZYa/gCN+bQEO6<X#RV=\Qg\#IYJaMXP;.6UVKL)bZ&Z;W3?e)TTee\OQP0MN
1Y?=O8Ag#Te.,[>(D=_Q?<C#3-VD]&-0LQa]_=_A,;d_#6^D+MO@g&2CdL]e1C>Z
Jc#5.@S@#3dX:HQP)aKO=-QO6?VE]4[P[2-;bVRPWZ;PMB7Kdg-?O4K6:;.@#;F3
Mc&JRPGVQ68S37<aYDL)c,OcBWYJF+:)#9TDMHGIeE?3]N60;-&,BB)YFTTe,Z1a
6LQUPeXg@ZGfEZPW)^UV4/^(E@+_]KE(W68//3b^IR>)fT?U2]-bP59]6#QCSR3+
7VCe?H2.5MgDESCA92dagL<A(5/IWNO-_<@-V.;g<974<M0T2H./^N\b7fdN(DAA
+@T2<JgX\R@8#-SJKA:PaD5C^T44I^Q<:24d=:.C9W-S+]4#7@UK]<#PTa;f2CNR
-^8G>J0_MCdQ=EZJ_EM^:,EO<L4;^;BHYHTCcG7F@d&)XKSDFP,<@+HI29TT0ZWT
b/,Ke([[eEg-O5G5_Q/OP7^J[;O:XC3)Zf[QN,T/d9e5^X8b[Lbb^07FcMKB0-)G
2MKH>K61UZ]-4eID7C5C?d@Y&<7]V@ED\LJHZ2LL&46C?>QY8=3D4X-4GbJ,XDNE
=R.14AY=R)CM7DZU9Od7Z0cF10aE;+,0eNDQ=g2b?]AZT@ZQX3<F3\YgGKU;R+5T
?\]J49&H96<Y83EVLNP;5OP]9cSY+YH3=8=RcV[#HC0&1,;VKWJf>g0>OfMK@#A4
(65a+QZB^a\22U-b#CG@(d4Zd<9eWI;][]J4_[U(>KK?CY@#f1\3aMD?J</aYK13
CB,EK[^Ad[+&,.JG,.?UIDO:0&fPK&7Z(3)a4FF?^S=5>Z#C:[7-H[XYZ@D@./M<
L)O?OG6I@afA1\HTQIC3DRZC\Q=:?Y_)1O4)B1V/R_b[:OUd,VOF[-4@=>A702I/
\-=DB529RT:]XV(7)Ddac43OG3-SJ\a9762]8LXSG@4:)YN4[3(Xe?d8:]bOIFW-
=>U@9WK/1N-:PFFEC_#W:]LF1.]+;ReVGJ+f;.SbKYG;RZb@\<C&-46#U?,7IP7@
f8T1GDX6(LW_R7B1=e@gCeD[YE\\J_C/UT-a:(;SKa\S=)N0#eEHHXOJRbB8.9)6
fFb:+fB4?7=L[fAJB0HR0H3XV->X?YJfdedRaUWQ<9\<\+dXVJaY=[MbW@^_Y&2c
c+:?\K-OW;<G_DEGZ2IN&[#-15(K2f3F#B17JR76C@?917VA\^^bFaRW1VW9_>?B
gI@aF#L&_1]U<@WX,M,TR@):GA-Eb-:7G/H:\,.;EdT)g-6H@CZ7=I7I_26dd,LD
Y2ZO/017K7WVS;=Ob9GRCK=W#@d_NK;)-;EI-Z(P3=Ebf__Ra)7eT?.A[[OU-=]H
/;IO9adQ_cX\1-D^624>#K5NRI\c)3INCM)L28->3D9aK;AYg-QP+L#G4F^#cJc\
cU93MZcGPSZ+K@^2WV)e@7JW^?)ROPH&AXG5J&DE1AF\[++Z@_D]_;\FVW8]g8dO
_C<RT7SQGUa-3ZGa[,,/.dJ5Jc==O<=9@c-;[K0_0TD:E7MF1(+,\d17gAP(DZ+b
D1E(CJ05)L8ASFIC1&fI?--3gTf?YB/J0dE8IJ_MB&HH+HUGVYZ@?ET&QB.4B=D.
)P?d/?4KL5BJ1fBe=e]BDbId4(\Yf5:da?/Oe3f+:[056U#KaZd7UB;YR-Z^Pa7Y
,5-EZb6O</-cCMZ?g/,f-N)KfYZVd(MHLR<BRO_S+I?,E(c?0+8]c==04:>K2cAD
(d+>BW//[HGJUBU(VO<7Z5TNC(\K/&#,+^RE@WROe&OCY9.TE5<Lf.QR+JPd9Q?N
,I/_D1,cPFGMc(7PJ.WZFgY;-110>2[E(9.Q^;L>2AM9EHT;B5\=15V]LFU\Gg+T
4T>0CYU7:dEHEe<OAU(&[)9dR=758cF7/63dBJAH<7BKJb^B,eD04X#?V/AC+@9f
YH@P8aB7&Ef+ULbA<]IWM..E:KgWK0)7=I[W-2+M[9ZMS67UVH8])6&3&DPYAO9c
8SebRaG<LI\b@SScT3EcUVb\>.#Ka\:_eCQ;Ig2?K@VL;BX_Z/:S;Z[fAQN[e5JN
aNcI7aXU^Ze8WI9PUSY]JF^-A?RB(2f6cU_64JaOV]g([JX1>5GO]OZ/#^fKBAP)
)0]4WB<)-#JZ@&3[@b(DGcMdD=Z.bJC:Q#M^Vg)YT-f3RYDWE=#P?-HV5/ge7cbg
8;Z\0A45>95,a[PgXEIa.1g#?:)+R360aK4N[>YbY8f0fTFQ1BZD[gWc)WBF76O/
.(DH(<QIPLOfE5-BW+TFNWM<5Q&,@0Of7:Rfb,7a<R6K0\SS&-NU?4E&Z3:aB:gA
JT2E7(dWXKdE-<9:U#1.+.?W)&]:f=X\^QW=X9=T4B72]X9Y8NCKee&UF9H/WMTf
D@\4A#fAQ;9dF6SYDeAK8WG2SH]:B[40IIR/5]_UC20TE=+7>2fL:,e+9YT]UZSO
L/5c_4&N)THGbRF?:T=1#GH#2W04K_(N=4TZG7:?NNe1A,QQf54G>-)Q.(e0Z+TZ
@Y?cPW4=<IL[GWDBP@>Wa+);P[4XE/9R[4dZ.?N]Jc(SP<V6aG>#N4S-?DfHGSN-
P.e.9Q,WKV:\=TEa)V:FFHbc]1E.NdV87Ug-\Y0<bf=+gIB:CRQ]f=GGZBE;cM59
12;1QT2Vg//4MM_JSFO+V6?N./+?C=Rde-OMgQ-TXP(IO_=17)f#/dQV:VY)T/28
]LS.33YK:(a@[=/BDPf4>0F]bDU?@FB<:Z?(-KA/R7NfM;.a9Hc.E51W<WW#M]bV
;Had9f1C?A(V\5D97CQI1U=fM_>;<=)VCP\:7-_g:0K]NCe1)+>MHT8=_.Ud40eF
+bUS5fSJ5EcA:+>HafTL=J,-g&cY[)(LXV7\ITT(91H8.3MV^CX,U.cBC&=GL>W0
879R,7\]<72PG[PPDU7@0@1,@>_/&-F9-/13DG[^2]R5/@.^V04[ZRLbABD<CZ]=
EO4JfRfEHMZ2/D&I4;V;cc\2=b1ER04DMOZEeK^8W=BP,130\P@1)g(;c2F\ZPbC
AM67XEA_3BT9/Pb&SW@CS.4\\dg1829VM/PG2N,g_/BQEWT1L@:((M[29YVMH1@?
2_:D6:#C.C@ba:209KSE[B3e/M.cf3V:bV<MHISeKD9ZAI\IC(.Q^0&NT7?,)5D/
a2P2=R_HIXd),YES9]^e6T66072HIFE0G7;Pbf+YaMR:V@3g?^DJ@8NIc\L-e8fF
_>dQQ#7A3144IBIQV=bFe?/A#Id/@SFKOHX7]J-166(LC68dQ<RDS\4ZRQ6)R6;:
/,+,@4V&c:]OBf.ASa?T3E/>eR#A^?WeGN&8Q<K8PK(HbRc4e2)3K5+Leaf9&]-K
I)RV]:HN(I(:S\68d;ad@d/6S[d^XGK\J2g_gRF#WQF^ABT589a;9B\I\&gRCDCT
T5(PZ8c6O(IEHW(3b67Z3/X(CP+UTKc:X25aK,_98W:6a=_3<J6a>9QWB;6?g@^W
B,3@=\0U-cd2&+_K^g80F0KdZ?I9[]LX;EF7M0>/6&^W96.M2X^T]Z>?TaX-ag2X
ILL]HR#b0^c[=VV?JTEI[H;H8#N?+Wf3ET:LKDP,^K-8)<L=#^XEWEXEQWN1=\WV
a+NG>DOQ573\5?.f,ATRXXJ@8>US]4?P:Gca(3WL;.N;9:IgR;&@QCAVa<.Z2_#J
7_bH6B_O9QVLK13GP,VMM/1YONdFY,,)cIDP6)2)T:P#8XR@?.=(N)FXW89^c@/0
]GIRJI-:XHT&K(GBd=XQ[;P^706J8aG[5^dVCZ4b/N912\4U,fVSX#aR6-+e2baL
gSaUZ6FK0XLcLMHPW\g<L&,)c@XT^/]9U?A1ZG?I#OgV/1MGT,,OZLN\8M>9HWW0
L/[<X#?aa;S_RQM^\cLZ4PCa?C1HeS3:@5(]@ERa/V:<M4WGD<K.=.R27;7^.=Da
O2<CaY<Y<X9E_(BHF5,7Z3&e043gW58B_-f9WFcU.P2J_8d[]TfI^CLM?0GLeYVU
f9HW2GP4\,;,WB,4gdT.AWY[?<6bgI-RK8\-;D\>E9AbH.ONb^Z6W)c)>+,[=H=C
N4NI=P3]U4T@C+a:b9g[HV0dS0-^V;;LVQf\?_b510gN.>[0E;+=bNNW1DYA>2\G
KNR-PEV>(S97b<S)I3Q7_Rg-Oe<U:9VX#HaWF834,C___7=S;bM8MD2/+HU??YRb
cQK1OR0T24;JcH4F42[BP83CG-61gFK&c-BD-0Q[V=/3_X9@&K.#ae?ag+>>cOH3
O7:f,@U6=5],<W@XQ@4<RF:;08d,Y]JgAfW2e8>0A&[VAJdf6E8^c?6=_dI&[1T2
1e3H[4WVgQ7gS.4I&VO..X9T^.2Ha)?3R8)DY#F(B[OZ04@_#I\e[@[/#gUPYMe^
))\Z+O^;B0CYW<_7XC4c?U#+6L11HDTR+_d4MU=9W799^O5HAW\M1Cf[cW,-4O&4
/+,OLVVF@RO0=?H@#J.>@EAZ3Ka2<QBJaObg>H=,2M_(GDOX+@DGHC^c_S.2(1N]
a-&d#:/UFcO):A>EUGa0@&9=5UG:9M;<VYcH2Y+8B(gdI+X2&d8WS+_5TXLVV[Ag
HAUB-GfN)=;MU<LMJ-Z8QZ<WC4#,9Ae;Sg1=@N[YTTQ<&HFR9M\g,A(c>4J23&3A
^BG#&(NRV[F?WIQSVL/Vb@IY0LWZ./3?V?1:1QWFY5#FMHR3Q2,:@?f]2Vd5DABU
X2=;,B=-[(ed].)fW7?Q]5a86ZE\D#_RA9]@FORD50P]^[;D/I-^WDTQfg9OSgH.
2\G2<OM/Z#NQ(GIcUgK<e)OC4A9L;1O(Z8?PE-IZd_TWCH\RX44@/D\M793OQM<g
R#>C-a[9Fe9Ee:L;3F.4g_J;JSa(Z/?_bd.;g+C]K_bG(GBN9cNV>4Pf<95W^1&P
GdB&&G3-^08-/C7F,W+c25S8C6<7d,VPRb]E1]C85.9D8^7a^7Ied^W1d1=R3M1X
[3S5.@E<8PRIZgEBG,cA6L,HS:R].@DEbX>;+TBDH#Cc+SaTgF#Vd0_7<GL064gA
L98977eC4.+YTJM_d]\HT#&3L]1O3>_W3>Z+N\DF@;#I2WVOGZD]a\Ud)6K8(_EY
0e=8OODMXcbTEdb=O)OO^--(7/YR5]eZ-Y7OSbY^BZ:O?G=61+/:I>dL<9HdFE:?
NP.G0Na@E+dEB]#1HIJ2:W>R8+L-L=0[;LKXZ5NLLRaZ=9=]8+<O;]SV+fY_N:UW
>5?H_2(Ag9B&I+T#0Y2J&C#44R)Z++aF.ANc?XOPL0a&)1R\\F,a9R3I&Xe0]D3B
UY>E-0:(gTPc&EH]9b=D2+<4RL?:+:P@Y=#>3TZKHP=.Q?INLL/=W\7N7A5PCW+/
>df)SH=]Mg\6740U&KL_+:S2GP-IZGTK1#]>Q5H[/S4&QTHf7[_9g\KgXeeeN+Hc
UEB-8EY+DXA+;]JK^,OQSX-b5?-H/GJ2:5ETT.AGMJNHcKJ+1)+90EYGNY./gO?a
T^IRc7c1(g)6^\FH[FBXgOKd>@G>Q+/2ZQ/I7G,?A@LfaQ.ZG7:D4C8@fRPS:Dg8
L8b&(]R?-/@>BPYc5FB@8YBZJE/_\\QKeQBd.4]<dCfNL9LZU\P(YDBFU>;;1Ad:
cYQ]M2FdU6_IV6Z:8=AQ^A-:#XMC4E\,<ILHbX5&fg;=f+;]5U](9TLfB,Ua/H9:
992:OZfV\,]D#1?b@Y)X+E4#FYMa1<S)UJfOcF8WV.c^6&Y1.ecF/_[d:D.X1<f.
+:/4.aV#+e&?C@,DR\E@5#OM^+)\61/<@+>)a)XAAU1_-4VG/;H9\fY:_N(CZ8W@
T=Kd/2X\bBYR@g?[.<AI;33H;a^;f-8(fcGH^?-IcGU^KJAY6.O)c;I]9UI.Q:O-
Ye;g4GNZLdH59gFL8T?NZFVV77\JX#G;\2&<W0N\XbQZEJ/1gA3TL&]3BVfF)fYb
QYEB_8KdB//#,5R4U:Nc9YZ_YGe,WZ&QK6.>?U5?0f2c+CfI)X2+[OJ(]cI>N^Xd
M]54H:;X_77Y086d=HZe<&:LQCW-_TUMBI0YCg[bIDWf8aS>PH5E#C#_HbLU/66Q
(aa5WJ90,GZ4J0XK&=OX[DB(XX22[e5[Q;ET8IV>TJPJOYfS@;cCH^L82Ba](55@
X_)cQX+SKHd.62,)ZZHRH<e/=Df<5B@V:J/EL1ccG_LAU&-[[GS?6WP(K@+.;K:R
CC(cP1]f(O7HWNW&1/A4LOGD6/#d^(3Y(LFPEOU.Ga\((^4dTV[Ua8/+3F@-62f=
DIK[?C[2>aB1;NL@U/#CfQfP\IacWcH\BFdM,)J6_91Qf^UdYG9fe&e3F(<CA.D1
-E_RfE.CUd-^e+=4F#WHJ3)c^\;^6XVd8)0^8Tdb[^EIU2-8ZI0A(&4]8f(7BTd7
D6Hf3.4,8@Dg;;R1\4M/5.N+F=Y=65b3JL1F8A2WEQg&[U/:6E\&KT5dXQPS-b0F
1&L_MG#c_O[ffaIC-(MQ[_98241:T44XCRU<XMJRgbfM3\;LK6K13.TQg+<K-/a_
DCQNCU]JeAa(\5MJH4>YK^-L;9R:FKY6P<F^eF&>&#e=C,]dWCR_QTAI)dRLI;X0
LW5eQCNfR@4BIR)RW;HBA^R62K1)V58_R_d#6AH9\6@N,Xd@\\7e&].C6&e?8D&,
DT-gWH1-M6J+0ENG(eX8V#3V,&14NS0:49HE+9VA;A1DR@cBQRC=S=O09_CQRZY,
3@F07O:<DN[:VS6665W>\-K)f/P=;8Y[/a]ZQa)K@KHVdfKL(73W=aFb9gJ6_CX8
A#4=4N0<FRM:NCMUTb0.]L<8e36(T&>3gR)#SU6a7:W9X/<)4&#aVeD&R3dW11/(
T.][L?BRY1[61RC:b)&RRS?Je@+PcP1NcPV&V.D)X#NZ#/?EYCdK.AZ+?5(/g+BI
e83W)<O(?=#f-Ig),<U?:E\fV@:WQZ5U:C(1.BM-J37FJKb0-dNB^XcaZc[FEa_/
CXPEUR(44.?XEcf/Ta@(/KBWdE>:J94a(:HFZH1]E89.@fS^>R;O0D8<Q^VBAdJ6
6[;=3T)+R.\=8CXQ7_7cIIKf-E&B4@Ed0N1ZcVa(=\L:L?GYS;_/)K.SDQ6OUMUY
A,H+@2<KGd,Q4Z,I2EAX&[eX@(-0b^4Y58?MMSO@0.C5G1=4YW^;53_=]+a6b#7?
G[Me@G>&dMF\9\7PQ7OVIEMPb\UAEP:1Q_CIOBdAFF>MO+-bK?INJ.L)_@_VH-AQ
O[Nb2g).,7?T=WVWF5_-66E,<OAT(5SUL_\g>OI@<>NQUDKBC7-JM_C_J/K\KH/X
Qe;<0&B.XTbf_)>-LKK?+[FWIRKD59I:7<Z;J18W#;HR@^[_7#Jgf[-@7d2I]NcP
J/6,aa:UdU[T\8FX/GM>c=X^7Z_[SU^LJIKf<SWIQV#TL?R#3-LI08,E\P;cAIC>
S2FAg#\NNB)+O-LATG103d#[,8b6PGOcIf8aVWVb-3LRVK^M^@P?1XZ<O;0,d#Qg
&RD^TZ03K(Z5_W&ZJg\3T?.W3>8,Eb3LI9bC.bXbb@3@6&ZOVI5+=-<:F_M,S^Y3
NIa:Y:aa<I&ecR-^KTPVVg5^V+/=92g)PTF)[D.^.HV2L]@\e)?MZ;Q>L]V;=d)-
A^-b;5efa(^XF14DaVJ##V&TdNa?.V?=Y0I#U?FF(9<E=6A2J9><VSV(O7D3654L
6I89e^dN)_ZVDE^_.--1:Y+@U2_/A,f^U>JB\Z\(0S46A27RR[bf7g:62:K@]F-(
NX])2HLa]^6]8L/N#-6?>)c6<3=IS9>@>AH[DdQfH3T)(QDgM]86[Jc;\VHNW0.E
H+J,?F0AbALZ+C@K91RC:X?>e.AH@F56dQMTcRBP&WJ3eB=&\Y@Zd]+(_:>I]:0(
Z(+[GWNSWUY:8MIe1(^LO8&Hf+]:c_O?_PC<-784AY-53U&Pb.WN<;TX0W#RO[L\
3@DG8@U2QN@YFKD85N^YT55.DfDJN@e03@eN]fDWY?(0VP6ZFCNBIFX=a(H]&@#D
ZXFCO[86_JO6/=Wc)IBc3VW,f1b07LSaVg#gHY>24N+RV#b.0,K9)#773]0ZY2JA
aN5Pe\d0aX6^@T6I+<VK&.N4WZ<(BUQWAdW1NS5=:94W)QU1(SD69a+N[7e7FIT;
5C6c)XG+8HCEN(Qb)cFf81<gBH_H(>[[9O^dO_M]\(:+0P8AVd_=](<^YP)5.@&(
7P=,8Z^G_E,7BN@BeG&=9e\Za.5b[/-_?C28AZ2P?_CcPRT>UAM7FZ..(?EX,E4:
4I;;Dd;AN4WHOaACB\0(4aS<@,e:.;MDd5<Ub0:NB?X.VRSDNS#4V>@TA8#C=,6_
a;)44#D=LPK0A@8F5#@#I-.=396N_G-U4(\JV[)ID?^P#55HV&)Z<#)e;.S1V^BP
cYHSYYFec6?cJ0.@M(?@^5QOcL3YYOMecW#)H+,PSII[bEY\,-+(T#SDE#XYD9A@
.,UL8S3V&U6QKgT?[eRW-gXT9f1^7cS=R<U260M=ZCX514C=G_<XS.+G8]+5d?BZ
@L@H.e9b\TG9>S7;CB,HfL3W^21]9(PI??_4>B-<;Ef\-5McK^[?E0X^A7.Z\=#/
ZL+[-YA5Y8Ac[f/K/a:^H+=FZ)7HH&LQ0[Qcd=K&])AVAWb2D)eA7(^3@=8b4f;>
MI8V8]Va(]?T#b[ML^Yd/_>dDgd]6=eQCF;AGYJ^9KEDL1HY9+Y,ce[2#)U1_ea2
ESJ]G&PA0^GBGX9&U/8#G4-fNRCa5QQNI6e_f;C^61.(^N:HPc@B1&)F&fBZgGN1
==?0ER0AgJgIHG54LBCCVDDBT_5=b\>L.6IKA@BO.Z<,FL81\cb==(?Df-L2CWD(
C2Ba,b079GNP2.E#YMWaM5Q/T&=O^ZCLW:aLHdN>W>fD1cXJK<O?(QbD#PDJO9=/
7Kc?DaUKE-d]6PN@-fBe2=U#)Z(f(IU,,]#-@f(CTT<US;HZ@Dg-Ud.3O7+;;/=W
M73/#Uc>aZK6^UL&C6J.\M48_P/Wf8bRIf)N3-0Ue]:_JKb^F/8PY_V_NCe#8#C^
OM16c6:CbbgcT:9?);]=g_][<fO>a3b8[3>cH=NOZ3Y&[(SadX+<Ub+YSY-P.PHJ
H=OV&H#TCF+H5I24[GQ/OfALO?)H#W<DHf7F.:Le]dB=RD3YV(^)/eT\?P<>?D;>
=N,N:7,;#;2[29@S#\/VL)Pf#R-1[<N1OZSZgR]ed]Z+;SQW?]BULWVE/4b_<b]?
WcfG48NGd)1MNJVI;4IJ??2dcU#gVCMU=gKT)S[g)WSaf4a:;UX^]TIOf\Ed#N2X
Sf]:^N2\U=A3d6?M5/a],>0LGJME+0?5ZAM\5&F0KZ:Z^L24-adUXc@(f0GK^g9,
eW?e^77>T#8H3M-e(99PFg)FZYVR;:TKZe5dGV\2CBKZ.KPf7]T3W#?WOC[;(<WB
UQ/4;60,7;^KM(JL0-7R@>.e>H:ZH\a(c.+@IeP_1T3-1W.WOS4E4a#de5A;HQMc
GHI.a#/PNf,G^?(W)(^JcUXR;#JNLQ.(Z5.DeQ[eKW+eaGD8CYFKE+W@&I=&G7.8
/JCOQ^]))e7#2HFafXH-G5;AE?d^XFIMEL#ce.K;W\V@>-U5a<>V,.N#K/@\YRI>
SK-(LV&?(O:M(>O?AD-#ZDIRcJZRV^9GAUFD\)6F-SM4+DIR&L]LU8f)-=_XB0KM
GBC>7X.5b?^QW-H-,8ZL)eVI60D@C@F/1B@NNQ.>PWcQ.4)NO@.&3VcZNNSFUR#S
)UP#M3(=7.E>7\6OG=Z0Q>W[FfM][W>]D>_&/5fVND2:,:R=)9eC^Z@T5e]^P@:9
0OEg,AVPM99_FVPYCP6RD^95N0GAY@?1Y]a0f(<-G^Ad+N,A]c:7ZN:DP4DB+FS(
?]M&;-Dg4b(Z>5G/OLW;8(40eaQ(V32HG@M=Yb^I#WLY6./EC7Hf]<U,e@-H,>Q?
?e.=9)O<=)bX&D=5;+W)^S[.&,+_@_>4SBY<g/=4bJY4bb/6=5JM-NeJ)RI95].H
0D8:?FJYI<W]/>_f;-0JcN=G+.HP<+-[fE(XHc1g@G6TBK\Fb&S1e0?+fQ(H52A2
@[2O,9a._-1?D3K;(Eb^]GdVgR+NB8^g5_d4<?7bAUVL](DR>PWJNd50@D\A+?gU
NWe&G1Gf(gOCL(D^OgT@5:a8JT>-W([@BR1F7^X-+(267baL?LXa7SL95@R/M0B_
&.4b+=Scb\C(U)I4UN\O.NRb-#GHIX1V)P7:@Jbf2VILREMZA.9JR;?ZE(gfgfNA
>YE+Y1T+XdYI]JQYHX:7D,1=XcX-<.GSUb^<GVM3>1LA4H9bO>f4UA1^BY?[8gN&
G+A0d+]L.LBO-Pc-a.XN2_5/2cAUZ39fMG]>G;UYI,8K/;dg/C[Dc=3gXSbfHB<;
RJ+H1M9b;12+7@U6?)7f^17Ea);4?4Jg7=H>YPE(0b7A7O@)S0#3Kd4S4\GQ@92A
@+SN7JX8KQ_)5M/KE;JYgF363Z.>]]a,3,f@.T&P;NTU.S2XgEOCeX\]3.-2Y;T)
QRfJ3_g(R8W]SWHMUBC&1XWL4VQf\aa;?Yd+WURU:\,#-_eW(V-Z72+-[TZg-/I6
+Tc])374b4aTJE8O@T#9B0UM0@NE\FPb&Z0XJ51RVV7IM;-b;[22eE,.KOH;<DFU
+@XZ#bW[I+#>SBXS,&1.CW)+U#0>g\21J=P@6NQ>U@U56<6D\L;EU>Lcf[dC##3\
I_[(g=dIKRP0)c)3Y+JgFMW>aS]0L\ITWWS23WP?Rd2[R=_S6;R(+MB)?TGV/(Y\
>PCKU&XS_GB^O5?Xc(fNI5?=W+(?^-ReG0.6XK@#fSA+GOL(?VE431.#IT@;Y=[O
3(2aG-9SfT/+Z&&1QbH/+W8XA<8=QQXZ8^FDEB=1R?9((U9faGUR#VEK+Z?SH9HB
NF]=fd)-M6AIXfX+]/0OM>/#VeG-QD^>Ha5/.Fe:YZ2G/DLT93+)OE-/ICNFV\0+
cD0&LWMZ\2a@Pe_IF6d7M[.<JK>-0</7),3(G_^d(H(1QA&16348Uf8<FPM#T6DY
(I-1J8ORWJXWfdL:^I6ffW/))abW,;g9GR@+)_XagYI(@R,=aQMb,M-E9b4TPeT8
[cU(CW.#2^/<#a>>388N&#N1<(ACVT+T_DVV.:ENHHI]>Sd30S-9M(Tac5aS<0AY
U(-dbQ^.#SVUZfd7S(]Q-.Z<ee)I[SA/1@&(71GAX8#H&I=<R#7\[&XfN1:FB1HS
d-458-_(L\(a@P.Y#CLO7G(W??[33df_-_L@e3GWE6EV+I\O+4G-=)3[>d?,5[2e
HQZ@47FSE49Ab#]4Zc&>BSgRd#QReP8<H3Q&?NMK0GRLaW>/Zb#D^N(?PU,?&6E:
V=\G7R7_H3,T^L;HZRd4[F1>d5N+e</>>(CH8Mb)bZ);=0fa]=<^bLg1HJ=^95(d
CT?.Y5Ag08eS-]WN4a3^R(Y=9#Yg_6Q;62a+JN)ab0Y?Z)M@782X-WYbCc_N\I3_
\UH&@.,KLZ0gQ^UG^6-MU8#<4<(/^RE0?K=X6]E#(7f=KUT&&>8RX?TgcXbRTI\]
^e]=\1Y5fXHOOab8b^HXG7gb0AUF&#HE](.-?a=8E]GQZ<Xd.<]A;?]:c398U+_H
N=(Fg\,5WZ0X3>F9)c\KQ>B.2dC#OG7bWF;e[/+UEA>&FK^a138Z^I>bB02(K.-e
aJ1.87?@edXV5]XB[=O996D;D)IEPVK[?,EBd3]P(6S1ac0Z&FJ+e]c8_FZ:>[b8
7>;c1N;D=]5d5B25_^?=NHZ1Vb1R]d[C[?LQ+#Rd5J6C?YOT/3@K]g-bfXX1RR4.
U4U?+d4@O?PJCRXbP<e5+D/KZC)ZMIR,_LM.FW;S4ZPWD5-0@QQ@HT)1aI0D9Nc[
Nac6HMT)HL+DZc-cP\Z;NL>#6bS/>7/^X0g6E49)J(Y/1Q:.77+N]e:2Pa2X[Wa9
VLNb3&><gE:g:O[F^ebB^cN:<Y1,Cgc1YQ5@af;[0^G1I/;NDQV?d/F?HFaZTEdI
QVS]V-ZbO,8Z(eg-MQ4Ab)XcVGb&FYT(JM?6YATR0E0DJ#TPXRU+5G.aGQYEOS^/
CY7\<SDC2PLSYWYD:Y\.5-.4R7+U]H;+Z7dQ^/Ia&aIV[R@E2&VH>I&H9UW1RacX
E9H4DZ\-T;GEA7?O(>Ia_VbUdeRC;9f&R>XDFZF?(>1F[Zb.,+XY?bV9d4Z6-GN)
XO)HYV=V14>B]EG.S@LW9-WedQ-6B[/fOGY\PZ]0EZ/CIFeKKQP9[ZK8JfdC+=MS
ND8/c_@JG7I7cYC),XYb@+^OJg,R?42TQYF#YID8-KLE52Yfd+];>I-_9DLB:2Na
RfHZ+2FZbcI^?RI)]3FVRA8+#I4a65G3[VeERX9K9XN_O@ONecLX04+>dF6^V57L
g,)4/&9b:E=55Z19-^9f5GL06?SW?3X?ZTTf:0(NN[/\:68&FM:OSD<^dWe&.<)6
2R29gZ,S:L8I3LSES&0@Q=J]4@@aG#KdJ0TGX4c3+@a-JdJ8a\dGN)P8C=cc:g:+
)^f95I^JUZ+9-UP^J2b\3W6-CRf8LV1A;&[M0^+CK<)OJ#e,Bg\0];OPSFK?YK-S
D\C-=@NRCUG6bBac?Q5&-D>ZT@81MUT8IJ.&==0E8S>PF/UV,DfLM7Q<,HP@P@EY
UH7E5b37A_G5#<OU4&<KCLRK5CU-RB0U)UFfdfR9f78B:\\dRJO4a7DbL.(NgJ5N
+PY67d+AD<]SA4+3T.?/_Se#4D#06aD0W&C\)DQHcY3DTfe<@OFfW=C^?)GQ0=_9
T:0=+^)WVZE^ZI=079c&O73L>Vf?]0RUVQW=>e0:&Ab9LD8NAaHR&@;C]0>de9XE
?)=]ZNJX)3C/2O4-#?-ge);.b2])&0N5OFEE5<-e3gaZ>?OO^FG[J(f]G4(b8B2_
QfQS.\]VI\UJK:.3cV88(6\=O8HCcGAMP.eKFOTbCS:KXGe0afHD2E30,GL2LN(4
T9N]T=:_M3>UL\[^P,8Xg\>B?g_^0Pf>RObS8]cE5FUP(@F]<B+]fT>QZF6e1C29
Y2_:]N<cY<98#bE#9CV)#XSTH&a-E3DK8BQ@/Cf#3Gd(S:Ec)g#.&f6>OS<^#X9P
B/1fU[?._K;[QeMW-^-fAFFCF=F&4=+2f3?X8TD=R-H9\?T^R]I9B6J#+MEWAA,X
ba#3CZH4W;@gFTbYD2MZ?_.?Ya4_>^9K:QgB;GO3Q\N;KFS^H)G--6a[4INW]R5=
?)e#5e)##X9K^7+[=1;b^.OX5CE54FLaWgS3B^<>^^C(]238eQa(bW4Zb7Z-=FSJ
6T)XZ>;C4ZX?EBf\fbgL_\,K:.CfSFR+N4.Z>0NEQ,E\>O)(.7QU)PS14HW]M^,T
)B&ARb,8JU^X8I@P>3N5TN3(G,6:C/Q/_;Qa]<8;]c#-<g8Bd_/U8#>B0)O(+DQc
>bGe;BA5ffX\0A78MQ.F?=@96f/[8\6Pa]J+JT)#VT>K9H)&0JWEWG,[SMWS:WC_
Ag7VgK0(#d;g-EYF8POT7aOBc-,9T&M-)03<TKI.b06^=Q\C1:F1fW=1MO((@1H9
&(_:2(;AM&JPMIgfK9JIgaO7/S-.4C7JM(\@-OG\:2QaKE.;dP#+OOB=5cQ;5-TB
K2[YCW^S=)]5N0BD:)?B,GL^YRH=),1:C),@E2bTB;RcFL^cdU)R-6Rc7ZQFX]eU
JR6SdLCYB.7Z;>@gPb[,GNK=PWCPc8>beQV)LB_c4b<a&_6d9bZW^[]Pf7-X<2db
F?LP)0eST,8DJGGcXZ2L?GHXLDXIE,0]?.DcMWN,SRK3,:#+-W96bK[,N11\A7[g
6\I^QGY+Zb<&TYHb]_+K/c,P\^g70N+eE#?R7cJ^#M)^(/?\L[da=<C)TM54ccaT
AQXVgcKB1OCT=>R\E&cPFA:X&=Q_@]6LG>?10,?O:PO)--DA8b(2Agea@_-9Naed
OMdUHaO/+;9U75H@67Z(<CY/ZOR^d-gfJfF:9S,>/<C;Be0+]+@O/9^g1f6V<\1#
bCK>_1J&)]=VW44#GDaMU188JK^ET;E:82E1([M]G)_G9L/#@>M&(^M\GAA^2:7R
>4,Tf:3,R#]Q[HQTS>LGV_fRVI>;O:W-XY-cP)FaUM?U#W]WVI_C=7#@6^7CAY<V
97RW/)&CA&0&N&SK5,)9R:=3T:#K.L/O;Y+7/#YZdgDKAY8>0fW6@P:b>GP<Zc1V
JWgY0[AA29UR<5F&e]be:dD7HG-C@,e)g[&K,1,GKI,JUKT3>JPc;UJb<>(H^P.(
.G3Wc#OPB_JT54a#-G(&g-9B9_8_)0?)4>N#H(+YfJ/H=@=2eZVS3+[+9M(/DD5S
206V=).8.6QIOX#KZX6J[QZGT3D-N2d./2[/LWc,0#MK9+NA,^f3SK87gRdVF8cW
>^a,Cc?3O7[(9\K;MQW;=g\)DCTRI?AD/+IHEe_SSWSNFRPaZM3Ea>b+cd2)WDY3
G)C])RR7KJX_^FL4PJG^O3\e335=_@Wc49O&Kc+\GH3a^4\>fA]T#TZF_8=E8L>L
WT/W<c0XA9\6Q5:F12FWCQ7.M5Y&P:19DVNO1<488Mgebc9GO@0TYJ4I2gM6JIdQ
E_XFg9]:d3E6B/9+d10UfUdPX.f#4XX<;)-b_KPLd(:3&c7WU_M6IH;U_6gY?[0A
ZM;9R9g2C/67+V@@G4Y(@,[>HC[&[91_DQTOU9a(+EbYd[6dY7;X;C/A>PZ]-_JN
cbFXC.]V@Qf8M^Xc_P&6+6(Cg:FNE24e]5Q-=DgLF4,6fa&,Z1LBET-;DAY9gY5D
KTK[K)eQ5?[QS]+cX=S1Y,CdP:f7_4K--Ta(-WZa5(J7E^:<YGAV1;6IdOS75EC[
CVaYPS^Be0]D+I84)P0E([5^;O#fSV##LUc;BE&d#[YIQ46XZ>=Fd4?b9230]JPI
f0G(;#K(eG34D[2fJ7,(OE2))RO2U7?b(.=/6]IgR\@)IJ3bfX5[4;5g0DI+QGB5
3]A4#H_:c^LX(<+LE;C[=ZGQL43)3BZ7E,Y9X_BNS/DF5b&KXN6TJXHYe>cE;P01
>1c&_1LL&+<AAIG?bYDILf#Ce8Z<HTX>=V;MH(3;65RRSDaf;+S<_O4QXEK8_9,Y
K1aOb4f&-gH=P(YB5)?P5U<eE9+f[QXa4=G+QYT/ATX9&C&3gIU?_&A\QM0eNgc+
,Y+5WQ:.37b;Jg.W=bd<@UF#T5<#?DP:SD=+G91#/+4FbVTEDe5R[BNJ:S84W(b:
#@;H[ND7.YQU?R3OLcdTJ:JBQXVV]>\I:;gW)>#2+DU0.eV9]YD&#aa)5PYEQ,K\
-0/Zg-EbU4cD>cO-e6@..TdHc<OQ9IY0(/5X55M3?F(NX9aHVE]c\[;9J,4=c#)F
R^6L.?0K:;K\R#ON,VRUDQ]_\SY:+,HKI-OP7J8R5@7^_9e=:Q#JRRV[)Z(VG<-,
F5e.fEI<d+4YLK#CZ:eB23=MDWR=HA(3e+QO3D3f(EDQ9^N.HgefeYB/b[P:CcP;
]SPB/b_c.aW2W@LX:\=eP(/E9=6EG<-EfAG3R1GCe;-L(fHN:K9650&gaFUC:(CH
_E[ae5DP_1V7+IP//>++SB]>Y5(MGFKgZUX0IC1^V&c#^#OQDa-/Af=A)RQ_,cX-
@#Db7[fP\Y980O@_+5e;^:C\;+:T#O=9#9Z8KC>?\W&([?+LN/+#XKCG4g8)9\&F
,8>VLCZ[](9:LHb5Y0d\/&Z\Y\V]54VZE2;YG-dUPcI3XZ&cVG#g/]VNdY(@@151
CAC@_0G3Y]FR0^I#B69DIbV:1dM/<ILgUgM]ggB7Md3ES(A3?1+=RAJ;4[A6CWW1
_GXYOR2HDPPa9Ib.>TK^4.XB5g18YdDY-3LcH2O+Z)Nd2529;A_^=J;WK/>cHDa^
Fa)]+,MAVPI=a[cLFM7JA5D/+/Le;(/JAMQd9FMQ+]74S5bD<&#BGI;WJOg(3TD5
A:H@4@Z,eK@/T([@9(8RFRCQc6AN5c#a(6f@?eEUfDRfe<LO8MHQ^4#1:<RKT-d#
7aUaIBcc,PR6]Og:[239+0&&T.</>(AV#&9&QC2]5f+P7E^S@-L(F4BE6,-IEFdM
DN@Q73M5=3B_ZKY-5VSSRF]R4)f]&N\W95+VfPg4FZfdACWfU29UgI=L4FHRH1U9
CIE=&;W>4IZ(KY:DI1#3\f6:\aeTD316_,G_(<[[M-,U^&>;V0J#^SV+)aH5&KMW
HNA7Z68])g]4NO&Y,V6dP8KdWPNLe&D3GfY\483X;4T,c.Tc4M(ZfbK(Z#IFG&DM
5@Q@#M9DGa96RX]&LKBb2O]F^V-E@=b6D]2FeND?gc,(.6NO7fZJTNe/[@b>UE><
M0UJNc3S]NI#H)[3W9MgN>)+A>B;JZ^@[[&c?2(11_V\]LdSQLJ-.SPIcbT4-H>g
O_XL:N:C8cG5/CMO2g[eGL?Y0[e#d1b)EIVT<K1Z.7(.O;)X:-[IMDGXF7b#<f<.
0?)J5:8>LKG\IU-5+^e0(_bK/X8(QS#,2=WQCF[#Te6L@XZc9<M>TBdF(I7.4[CA
<Y,/Qc:8:]J5.G6CG-?5e0MPQ4a8gQ4gg1L#9?;4+GQ2?<#S1a>XKLDJ-\1R3]SP
B^[,Dg)(7W8V#R>]0B6=H+_eg@O119A>,D./83R\^X\8?M]#8H+KDQMYCMcMg86a
+NZ4cG=D]=8Q6Ea^Ye9\/Z]ZAW\OFLV<b:SIE.7>C,X4Yf=R8JF/]79:GV#G?3)d
,-db+d>JMBK[IBc9<g_[3AR>X:/C5ET1MFcTT&.gQ;d.]>&O/D/eR=<b+-+eW[,A
QGQe1/?/<e(fEZ@=XL?Ve?,5@4:)B4F@Q)MFG=4+Gd2(c.W?N65Q^GWJ#EQ/OPCE
SI@]NQN]K6/<M6Vd/aX<B0dU0H9[(5/Z9_PcaI]4]cd>82Y-H=WdbSL?c,]KfD6L
TFM@98UE?IVaXgY;-.0QKG\NJWU3O#H9;;_[,-1^B9+a:gZ:#(,]XO2&&Q_P\N,c
23L?.bD9MgUC93I4^)Jb#JPO#gN38b5;EEW;@[LHYCIV5@TN#Z^4E2g,J?)@Yb>)
c/H[?F]#&?3e7@U[[@:\49^YdQOB1#6LQ9WCE=Y+Gd_F,>NZ37bJH3NGN44TePAV
XI=\HASSCU_;I807dIEe8PcQ^_1eQ_/DM,42SQfCV:0O[G[.Dc//\8+;U<5.]ON>
3Q1V\8\FF6F1\D+8KBJ#8]Y(FCcD[H;dOA[-T8/<AMeDa@EB.7,I:1d)W<V_Rf61
_<CHSIP).3H^2E]\8;Y7Q3bI/.a+=QfUC?PJ(^476QE@V&cX6BZ0)9Z8CTA8ULM4
FI<O]P3(]80L&38W<f#TE6LGFaFF&C:3I.Z[,N#SF2_c,NNR(:9,LV?H5RIEI(0a
H]X,2W(52/W8&9\:2^Q2]+\4gf0#(c,6E8d6HUf4Z;cbQ<[NOTN<T0Ld<e+7K+.g
Q6_ZCH<:NY,LR>LL]:?,J[_AIW4]K^fJGD:CJY7JdN8;7KOHJB7B(PZ8Tc1OcQX2
[@,+R(5&([]DYDX)\-5DaLOf^f(62;PB->+VT=(MG58(9&fTYX]8TD(K]DeeQ9aR
/(cVK;WcYUVMKg//a3UXY#YX^08_fA#ScT@Ed;KaUL58S0,305GW7Cg12\S#dSbg
])(Q(aRAATFUNG#X+e:/2ggb:-\d&@&6.X1K065+6[L]CT(8,98_f&AJF9HO:DQ,
I;Z_1WR&d4A<0J._>/,/ACJI_[cGeSA93;2C6a3Oc.?4J(5.2-9QHRdCcgCW7)?.
:&9aL>6+R9fUe?ed6NZ37(:L)g]E6cT>4[T@6e0gT+.V.IN-:TE3GIgY&5f]b<-X
-)b[1;]\2;;N?A6[b34^a\g4?@OI:0g3M+gTgd5/0OV?P?AG20Rg3VBbbRFacLE4
<I;;XSE,-g4YXa:1,e,6=L9d)Z@@\<TQYJ@:I24)O7F)]adPNXbK#D?T;+=0:?]:
27_&TC#AdX]<=-MJRDM5CB3ADE3Z&]fUU9b2B9eR7<I30/8.ZOVH\P467D3B>59E
NaR6S;/@fg+dA6NEP]d1f12KYgXD1=(?9d#FDRd7QJP9?0N=3Dg3[@VWO^:0(O#;
SYQ](2T821</+9\JKTBFFb>f?)K7bLNd6,5<W:\@+ZWb(Xe22,X<Y):MSX:fQXHc
Qe>5@]<.S&\VH+38VJB72NB&+8Ibae.Ka7L+U0<:R\.INQ+=NJ/RT+>O-b/f:0MC
FKG-b,4Ld/1BYc(UG\bdK-g6/PdaTTA^d9V+Ie<dg,/fVeb0KV<T]@1B=L,gM<-1
&>#S#4THc4&A.9S&_Ad>\=<XAXCGO/WVZ)\K]HCIL79Qf83H0CPd/1Y^+X>Y0R1B
9N.UcI6P75YO6:)/GT8/?@aA_\Jf87[<4;30^W=V=_A^.=YR37J3Kg>\P&E)_<VV
F;Rf(&0]fUWOIDE,)f4_eQb1QA:]-PXgF;=?f(#PAZQJUKK\b4X4ecdPb,IFS9=E
_KH#JVB:>>=[AdW;F2>W/Ee2/8UP8?AZ@\4I]b[>RbZH,WEH:>OFb0\:X#G/>V>R
LfQ#[Q>3feT#PYZeUH\05H.L6acETBSKa^AV2#:@eKef]B?P[C2@:LV#8Y:+2W9K
E#IX#?dC-R,dCRN(O,&fa29H542RN@9:d;O[VeYgS[YF8,A^2a+>1=.8b?UUKg_5
6fFNHgfP;<,.dDO@5LLWO13H0D9-E61B.A3IQe,6=IMRN;b:)F16:1V?)bg)4JTM
16;539dI7TUeJX?:eIN=f+;&N5c&Pc28Y^^FVHL]@20eVdbQZ6C?4@IP\bE/(^J,
E>5JXb5ON4LZH/1T)5[=6BVNZYQ09(KVQ2FCDB^A/ef4A;e6fA\WKBDO]F3bX[)9
NT;?_N]gdQFA^F)3AC9,\;@:KN2L>gL@(Z(:=<Z3bN68X;AOD],V-75:5UWT7SbJ
7<U9)-L,g4+0<)aMF?a6F:=_fP#gA&3;VH^8K>,=>7-T=b[d/K86eV&#^a)]20JV
6c>QLBLM;1]0W<a-&b4Ze#??LM[_KGO_d;-X:)5(2G<U&f_U8_@fWAC+I>OSVU-0
PK<I)\_U7N63@LA9XKB1\X1P1#@(K<::>[=A;>d3YU7/FC1ZD]&]2>PcD3HI-LcT
aH=ZWWX(QWEa3A^_^,e+V\)(RBEZ:=LJS,?#.^Ae.LJSFX>CN(,T:gSV5][K,S?[
aX]P]M9<)OW>NQ8--27AKW-T(UCgJMUAeCc=9^;CC.MN8J5JHH(<BE#F.6Jfg:1W
Kbf)RQZ]N<C8>cN<LLRBcbDfM/&LG/F97X<K_HAT-5g/X3->K9LaH6EC[GPadea@
YCP;E\(;12\MAa4-N.YQ<cRPI[_;]25@5O-TP0<]5=ZR\L&Q?]G\-\Y(V>PB@:(a
a-LR68WLaHOQ]<ODJ;cE/85M00BbG&U(c#a]54c+2.0S[XN])MH=;,L:ZU)Z9FLA
^Y^2)L3A,8M<W^COfX#g+Gg(\;.H5;M1E6g?[]FdMYU#NMUKE?ZVA]@+dI_DF>BV
-7FZ(/(IQa9_?B?^>&ITD<Z6T\=7(-SeHeAN:e#.4M?K?T[)(Ac#=4),I2B<(8B+
Z(6fMST#I5I=UB]N?^NS,VS,8R^7=L@@?4A#)X_+YQP76?M0&LWRcDYX/>fHTYQf
LH2(]^#FX(B0FPU\G36K,Y39S>\6NYf^Z7_S;9&=<J)+9-QPAE5XUaaa[?ZD[Pa/
1KG#b\BY/DE..d^V.WC(;O[Bba)M+Y1T1#0B>c-?F>99T;fCNH=BIdT[+^5aVMP<
]Ze03)P16TPQcW^Sad/S4MHH:1_^cJJEV>a3&UUIKK^7EE6_Qg@?fF7P]L&^30H4
X<<L[(^RH\fB\3c)R:[)L049=L.f<]FR.J(Fde<:<@RLJDL.DU0gKVMcX>C+IL>0
K2,,[R>)1N<.\8bD8?Q6_H3@WH-_^ecHJA^;B7\Q.XU<\:716Y?B0Oa@A>EF,RBD
gS2<7.]#aOQ54?XXR?BZ(\-gb2a-B4IIa^#dLCHIbeDTY62[/=/RA1-BfE&-0L1^
W(J1R81&dcXM;S&VRF=5@+daI;Qdb86TKYN0BO_2-e0/)Ja@QA?AS/TS3C13L8a[
Y9c8ae?;TX&&\\N-TE;WQXbO]+^0A2D[COd>G@M7]9-?5SMIRf@B)DZ-V6?CWH6(
)=FU5=O[5TZ<.#@dPS0XQN-5XF^fFD6F2]BMd30GD<N/G4YBFR>>:/4T=g[G/e/3
<]IB4f;BWWgg[CM:1BXUO^Cb&4H;/EfB=4eWWC96<;R/IXRE2@/4-/+g/^fFL#2X
K.,U]N;9<;X;UFNAVN[Y82N-UMNNOR6^61Y5Ybe>KP.-7H,IfO+1b#Y8dGD/,6bV
Wd[bg1aIL>OBRA?d#+IgVO[4_6XcPBZ/D;/Scc?0E\cf.6bQ#bcfGCHaUf?=L.Yc
HC7&U5<D59&N?02[8\6_[XB[5U^JAO3E@ZA1eBWWTSQ>76a.(5<F&+B40,Z=5Ac)
3OSM#HQ3Y>/S[2E\e>?]Vg)M]c&9WB0a-:]ZHfYRL>D:P,OM0gcR)DB0G/+?A);<
M>_GDe#8?7RWF.T6C6=?E,cV(0U]_J(0LYK<;FTG=C1W2SE[A_d5db3b@+JX<.HW
EWHL_)#a6A<S_@?S<eVD5,_FK;=5K7D=:N/&>eF42;D^E4+JRF^AAG6CR7LEad[A
TZb:@8+g=))Y=8^a_-JY9L:aO[SGJ-e/TPCK+,Hc4,R]<C?T.8>8WK62f7(Bc9W,
N2X)IIH-ZaV4P=RY<);a=.Kc=YY2#YgL7+B:8N-YKG/BdF[<:9T34FXH:OY^[dD.
<Lb/O&FGO\+(NLHPb9Z3?4g(.G.&WW.TU6G)T6L5eag2&D4?0C42?XL]TZ3GE/S&
]?;=_J9/0F37+1G/S#&M5e2.^OLVgV;#)Y,_/S@9_7.TMLFZc-;=[.YBB^\26b-P
5SOH,O=:I_SNgdQ5I5==EeAQ(SbF#g,d]JF-S9S<A8(;U^.ZDUSE,UPEMW8R=d.<
AXN18B?JXVM:>0&?>HX#^)=PDS_\ee7I\?QE@4WR44.R2UbD_ZCg)YFG.UB/9L/6
gYV2:09;=e#4e2e&-/D0Ja?[R-V+6Rb_&C&a96JHU;-80SVW:OgH02+ebK2?^2cU
^.EZUaY,A1K?e=eP(4aITT^IJ4CN7^ZbKD?SJTb)gXd-#Y<2L-/DTR8.7f-R>K8,
HH3Y?94_a@fN=YH:9P..(bB@RW>6DFdFU=2ALT@.d#FQ^?C7U&e=(]QOXc;CR.GD
A/Lf)4Y[2@T#X7XZ4W[b&UcSIGFL8;I<(]Y0V2OOedO\0LeaK>2:4T5]J<^]#)b)
\C@9E7/DPW4/B\^<E1\IPAAQ>@GK\DJV:CIMO1UP?KT\:;554LZ1[@ZHV)@3R@8G
fTHIH]YA^,:8&5RCB&&K>9V5P]4PH#]IK4gM7?36A1d8WX/_)>[@YK1VO:PLTB#6
,@N\6,WCSKDeJPMG>(LCNIZ7;;WYG>+26MN,XXCPP,Td)_g[4C,X^SVY++L=Y8:+
GJ+]1[<)AbL;K:J@0&&2C2GKO9.2VaCF)7gQ\G:eed75>(2L3-S/egPG30H<[6eX
X6W3<96B1gJd4F>P6XQ#(KT:[GZVHg[e>OC5.5(@/?]:[#FU9(c4J]:#L/0Kc>6?
TRED(RW,&ZII)X7Y\?FP_WNV:1DQ^_^-g]X8HfX:_D.HXCcAV07>)W@4SC@RR:4J
VR0;>f/J-=_TGL:G)F3cN<,S.^D>7LeH.Sf?&,bEP@4W,dg8.#V(V@P?JS(>83Y_
PIG:K,V2V^/SNbgL/<P=CM_B,?F=.(-/;5cPCL-F;XZB]ZCWMDB9eH@]+2+cAM<&
D+/_c+#;U3KPWEZ\/I8\6C:V10WeDa2Baaf0B;3Z0A&VU7S/?EM[D-SC;JMa1R=7
E6)R@V?LVJGJJN:+R9DJ\]E^4TC^KI36a8QN\KY8LHD+cMQ(f,X;R1RdCb7#G641
b</a2E0GDa^U4IFIB)O3)SEYX&T8Z:3J/8=-6@<3YZga-aa_A>I/agU;bE?+f>OR
^#F,af6adI^.C2#_?UDG27#[4Mb)UITd4HP0b_Y,S-09WGaSU,ec1cCg=(a(&,T+
,2:FPNZ78R.0N2Y(AVb,\H(e/CIVTB?ee7.g#PI@KMRZT0/g>C,4+X#PdDZWD>J3
a6DSIegT,BY<Da<751be^X\@[<=M3NWQ3ec/A/7aFH@>c9PaUI_8EP22^HEKK=#6
0ReMcZFI7(V,Ed^&?Me,3^a66JG@.b>RQ\S/fPUBgFM?b6E_XUQTI>eTOg^^9?E=
_[Cc;Ua^;9Yeg\>1=/A+1GbVS/PS\I-S_a<6HH6[(ba#QUE@R<7&Y[HJA^]_L^J9
eC?E_&RFT99W&QeHMdP>bC-cLLPGQ-,7Ce@H29@(A@5SO)T-@Bg>LAJV\7Q^^d[@
??2M=R.+A?8CSeDZXC;W=)4J;;SQK6HS67QW0g]79[BNNG5S>UObW,)P)cR[?+Zb
6<TfggIXAWE3A5QD+.XcSDB3;VFe:-A]98WQ4eI//dEW8(@.@VC5KKe/.;E8I;;5
B[ZG+BN#,??2VY1aMHEUN8K>NID\Z6=Y+7GdSHNMQ>\@:aR5&:FQ(UN[_-A(ZU&E
GQA1QU.M(N2QC;SGNfeY@N/J+Ga.(da=MI?A;.AXeR@VSMBQQ16,7:B;\0.cG;O9
G@0I_GS-4?FB/VOg:HRA?E289(\?_+bfU]0#H2_E;GO]I_<UP(GL<6H^:A&C<<VN
D<IDH@[V-XAQR.M:f[@<?Q6VU#e61L\RU:LW5I=-2[.B-3G7F;;f?.\._00=<:aF
G&43J9?SLPTU@S)YL<+P_;^TD-Mae[&E0>N?+Q:>LdMY^I>@Y,DA/OGO3VS@R.E4
-_/8^JO&USMS4cBafK>dU-8,TG06GX<(@a4KO7ZH.M>S:.)8C/LOKLcFW<bVX=W.
0?R,Lg0N^c#9H=_3aG=<\4VTc,K]7Bc.D.PHEMH@8eRKE[&+Z0D(K8)/D&g+J:BI
X(H#GPfRcJdd[,R@/+OF2L(b1bc<C4EO(bQQ@09f[I.cUCbF)H]K4[,=,1Z,[-RL
F]&5C)_)3&\Dd@=>E&<N4I6T;a-ZgPQTf)QK(]Jf_5/a-#NE129T6gJ9RJ(f<(-7
>I^Xc1;B166#34:N<X#Ab[\<Pc@#_-Z=0+e;Z#9.Rdd#FQ9L(C\[NH4&#dKT[/WC
AGU&W(9KZH5aU;75?4,BO([=/D/g<VF^3<cb][Y0_&5?=;,<Z.2^P)7IE8@LWDD+
WY^1ac,GD2gVF8:.7J604&F#JO4Q#S3)QB=4\L^0(eY7PZ[5eLXB^0BR.Wa1)H<1
K1c[&e:K2D?_?LVB:F(025Q_6K)H+X.VV];#]gVcE_G5D:e<#/G@IA2&/T0H)g:F
-./L>&=4NGXaZE66<Yb=)ZMHc&99eeQ#UQUa=@H^g(:V?1g\]#W+H8GcXBHb,.+6
5KI,2;.5S(\VV:MH+<c=^IM,3W==.)IYD+TJOKAZ_OH=-D0:EUUZ1(U_>X?=MH<_
K.g^N0G1gT]/4:68614b=<#FU)BIQGG6@),U3J;S>d6[eI27#HXbZ=RG^^)D8aRF
79,#Qb\/:GENef4Wg=_4ZH/40.L(DF9KdPB;-;D0(b;1=_<VNdW-3@0E01BHeZK&
MGH^3]NQEd-Bg3AeHJ7=W[PYRRQK<8FRg_HZ4;@/a,9,d(?3\^UOc1((K=;]@<&Q
+G)[bf=PM9f6ePWL8MVNN3RB>^M)5F[AQKMG;\0Sb_6[;B2OL29&cSc^=fY?MJWd
+gF:<DI<^P_)&&Y\_2STFW@b@Q((M^35;7ZN1AD^cAba-VeQM&J2D^4_WEO9b>;7
7e1),Q<a7NC)=J-R#5[:YRF4T2?)BROg3/XO.6:a?_fHfT_A?8^F>bBB,EONKZH_
-V)ZX5&cD;ZGIS?eB,&&eIAbg#9Q/KC.HJ\Ga=J.eSJ6S^AT6.:F]5D^(S90@/I?
OHNC@J6KYPSB?2TgIbN,R@M<f56>^\R1V_,<XbJCD5E8deU;W5/eTdE8+GW_Wd7D
eJX.G/f+YMED.5::G]_^V]9BQ^UQ?TWQY>,DM(/B_:V?84=e=H/VL&5MX-/Mfb+F
[ZR=f?f:6I[MLJ4+Ae>7X0:O:/b77H/#3)cV2;(A.bI>BKUO\L-U,+9#(]S7R7E)
6gF9N.@3D;T]C[R(IX<e6UK-)Re7T3.R9,V05#Le#E7^<3Egd=)>>cf&T@b0,AO1
7X3;5ce@4D<JJ;F@Y#fYCa@(>ecL:_cPbY[)MB-L3<F5\EIX[_S&0<QWCTUUS@5.
)?XNe\O@L/Nf^Q4G4eZ.PFJ12S&Q(g=1(2;447&@cXYG+C>UDEeD39B]CJ)LU\1C
F>]a3=#1IF]+H#dOIf,;^+C\^,<<cA8+9cD&Kd8)UA.<5[B7R2J[_/MB,WR/cbTM
^>c>W.3LJ0D1-H<e-D5M-QaH.[CFOH^,SC)4(_JD;=FE?I8UKf-=?c8B(_DT]a.?
c/G^1@N=,6_:dMWX?d58+RJ),d4M41FU0:NG_)C14a28c=L&d>UJ&G>F>8XP)GIZ
ISE_/Hfa<AcD/H[)ENFKTg)a=M_Y<#<W_a;QF.OP>V7DF@OUDO;8eVLA3RQ19[\;
AA#BbDKD&<J-RO\3&;cC-4TbMCU2ASg8,cO1@LbdU;I94IC[AAX>A&43W\^\6OaX
T[#3(cJR9WG-V5H6N^a1DSc-gJ#.62?,GV<<2AB1_HaV\#+AG\.YL-WQe?84Y6V4
W\SX#@M\1G;+F-I#IE=^b/-]T0WcP34F[O.8[ZMW2^:_IL6bWaE&^,-5[G&B5L<1
^0+N)\)Fd(93CF0Z5]V]L8\4/56WK)@_]KY=[Q[.DT41VEgV,DPL++Q_<..IE;)f
>&S?0?0)=e=d;JTHH]U?XgC_;DKUN^<5>)+f#H@fFS\_[_1@RZ7EEPWK.>C&DRKH
;cd/(>?,F57&?U@C9K8_&=]]gd_Q:LBOH/I,ZI&VMMDd1WMIO=X>BG]1&2F9]-.:
-5W_UFL1?;KHGDM5@d5(7@T_(UYAY;d5X]cVI#&\1W085]]BB,P@eB[(=;bZ]1Lc
[.I;aY#\;Jc:W3d-dN7F?XF,-^X>1W?MEH9WeJ,P=MO(UXb:;)8^DF(OKJ<TV&UU
LBHP&=3YWV]=4)M2a8](\U,][_Df=YZd_HVg\LAH27WUcb6&^P3c+SFUeX,68PXb
#5_>cgfM4RdEW:(FgPbVd]T5LYG+I&bBd-KBAYXHeG0eALJI@H9((dDTNf@JPC1Y
J6>BGD9MZTOV/XdS\Y?KN[0M;ZZOU.[,,UXZIVGM--WTQ<7VY=.)H\GB/NRO2#Z^
U3a..IOac.T^+0-T>T=Y]V9>.BS+B[_ZSXBW8[Q?gK/=8)AM?CgR)7YTg#WaMa0G
1aNN]R02^>B:5K0f<1>g(<S96GH1;H&OBL(dM@:E_)Sd)Y-/FbPJQFXOK.E)8RJJ
BgL4M4XeH?HI.Ld?b)(E@IXJ#RJ]SB6d2T4QA0g#LAe?7(C<(HZCc+>4I.SE#]0b
YccF._6J/T;KXbCD+R?I-3_-(<40Nb;N54)5b;ID5@RAR)=7EZ6/NS.IO?URUCbZ
O@1Ig9=S2(#7BMA5H/2Bf961\FE^(7NM?AGQE;&X6)Rf#>If]LN6X5J-OX8QEL@+
HR>\UK)QP,QfNZX_Y=U(-PcR;9SEAM8T2JL1&/Kd@G3#3-9M-F4>>5L1NP#A(OHM
58@,Z(5C50V8.V82N),J^a9SUc#DH9&M740X8GYcYT\@BA#fVOWW#^f=?7(;;[S&
&0:[:D>Y@2RD<V0/(^ZYM^:V2+..8T]2Q>5DJ-1aGE>NA398#W6Wb6493Kd?Y8L0
Q8P_:0Hf/Q)VC=H)MJ2B>-..dG>8Z/N7Gd.c<C_4-^bO2I20-bENF^)R?<E2GLJO
3QPE\X0U-XDc()1\(;_U6D[fC@GBWQ-OXQU6H(NQc[M&EbOW53VTN8Q@MKR?4[&3
U[+7Q_cAK7.1_20I/G=4fGN2UTTgeZ1d&gOSf.V0H\15ZB)a]IbSMEAbdH@NW(84
)I<ZX&9/e7=[WGOUf(JXRg45ASeMHWV&AE3E#].MQ;=O&NNC#MLZ;/7K5ZMc8OGB
CaJ6JSNbSH?09G+^<_07L(<Y528>F)-I5Yf/-Og:#XDSa9POa:W64<3.&c>[b[5M
MX,A3NO9=[2B#8E;C0^_Fc0]FJE7X>2IK1<)@@?:?_,8a_e=CO5,EE[eL<b3Z3M,
5Be[47d-)V8AYN_=Y9Y?IF[V&60cP^5<_PR9gO&^?Y_E.XP]4H+7D9O(T7WUg70:
e5Q:7Z?f^]d<\He-@9UN#cJ7^TIK[gL3K9e[,\Yb,R>V6V83<#5d<)-;WZ770^-b
JP2#=T/8:[\bP+PHEFFME6?DEF1ba+1d4ZJ7\RVIHUb]VOf_R96\dJ6.&ZOB1:PI
(\MNJ=.&H::IEbF>+gPA3/_>A<g/XDCS)@LNDM_Q2I,TbRgeg2J&8_8BH_#]5)BS
K4ME)TD-1^W1OM?Q:9f&1+U#CLaVMf.g?Q)W7M/80,a:>^Qb=:V;XF&UP86De:^(
KBLVSCSe\T?8TSJg53g)7/)-RBZK/5LcfXI8#<8M;>J>G94H/ON&I\62FfKQ+Y+Q
YK\N.R\2/DcLM@Z=DN4&^]W6:RDXa_-XZ(,,;)V&INdT0)N<a#S[IF1D6&\f60&\
O8bebLd^;=M-PD8Ted\P?E7.OSM6&15bP1f4TVcEa5c^#5NV>C?V1)_FR=C^MJ08
MXJ20G;3W)L-:-/P9QP?8L>QM+4UeTeQ8ISIKBb+I^6B?WI,K3;<6BNJZ\>]Z>\E
OcHIU?=g][UNS=PcWD45I3[EEB&&#b_.Q7(IGO#:NRZ_&:OX<]dX[VYa/-EcE2Dg
LAR+5;<5PYc.DKXFI;JT<X&A,[?B<Q&1^1MPFe;bCT@N=KNF9(9LW(Y]WY/8:1d6
7a]L?VK\26VU]<gRd-Dg3F))4XeS_SZ1D[d#PJVZDB4bD]d(ePg2DQBJ\e<Td:]J
E;.HAI8>6\5:L[S^8EFP1\&)IHAHMPPH8B7c[X^NFa.7b;M&C;1E&1;DRYA_Ac^C
/baC4M=X@aO=_(UNB#f=M.8(7B,a,53BQ8gBFXGD+1&S;;P>RHM?dbFYgJeTPI8.
6ZQS<GGE3[De.]<&3:3C+0=R4VX196YNG;U&5+>^gSYNDEcQ/PBGH_0eLOW;79OK
:G,\V01gPa5&X4&@F.cM1H_HbJ7C?I8DP2?N4Q&\GYGS#cE13V\#W^F1UO1E)ZR0
8e-Feg[5WGO5Y)T_a7a?cBVK(9KAQN7FNL3M_=@LcLC7NTg29]A+.e.YH?0g.5:e
/@O[JXLJeB1Qg4CR^PXDTAMS8,X?[U4TA\7.cCgK:?AC&,DY2R^AKa=YQF4F&,dV
,3^H=>45I-68Vg?(NX#7NW:De@Ta&H6YM6YgG4,M_?6HA=&KW?>8DbEZb)^9YCT7
0G53/DA;d;<Od#RMS[^85H_R-_//3c.=5f;(U&^1I@NG9]@0\<GL.d9T\:DTJ\,[
6,dMBO0b/J_?<aGcJAKOXWAS\JB737\^&=LM+eI:3-6H+]^806aV;+VI_80ZN5;S
/9Ia\\<F?M:(7-(2Dg/[MfALg4b37XUTf1WPR2]@3-;0AT[ZgNCU\fNWAG/<ARZQ
->1[GFRDdLOGB5eVCIZKUX1[RGXN(_VI^+D3K+gL9:QfW_cB82=&b,cE9<:AGINT
QC=)X&SE7X7_VDV491dbcD>gM)a#fa/3,dgY19RB9+?54FE<S<b,]P#+U]K_X#U;
PET61dIN\LCaA#:P15B3Kd9IA^\V?;a]=2B>5;K?;ER1.G\.^CHL0Wb^96C?6W;?
KFB=gO7;R>VOX(dEO]X5eSVAP+fbAQMW&eQ2LR@9U\TR7;-9.8]+W@=I\Bd3[:Ye
[6YQ#<M)RND)WR:7eN^=&+]IW<f#I<g_G[G,R?6S]NB#7T#X,=4C(&)QF\(Rg;[@
>[)&)VVIg,,?65da1_9G<>X:XDM.=I2YMSDb&DOWZ3]g#c[X<53>d]S^_49E8D=I
<[N#T,;K]OK)acgP/+,@F_gegWUcL<O18aZ/9fUD>dcO0E(aV.VS5c60@3D7Pb@2
ZE&AK,[V>TAI2.I+5<g=KJAGY[VR3>FJ<9F7-+;7U\^FF16QK]b=:7//g.LTU?0c
;H1:OA]2ECBB]0ZE.770f;P9Z.gbG=^1WO_.S>F@8RBYP[,=1]O>DVa[7NDCDKg?
dY;:GKe(NU?&W&B8/<L-b\GUC6f,d7B-L_PNT)YA,5>NX#+ba&<I6CFQWMP0LZWO
bW:/BG2[MdGWAVJ96U[]=,V4#?a=4Nc]LA?>5AWeR<@?\NgF5d?b\IBI9:F_G/7M
Y6;9(0@SCV9YX^LR6N)5M_0QPBGVOIO0H0Cg.HWY)G#81(OZUSUg5]Hc2.3d@cJ@
9E(N[a:f>S/#,T#U9??Id:c(Q(-3I)H)&BcBBNg8bNMLK8S5<,CP9YDO51VK2D?7
7#GAQb]T_VQW)B96CeST]]=(6967M0D/^9a37X2dF])c7Sc,R\2G_4B,3IJ1@e3&
N.S-27JGb:bT)2];/DaHgSLD-(Je,:C3RT(aYNSX\b/\PWbIT,C1-RCGGgaK)(.2
g7@O.J0M5NJM>]HCD]dSZ2aKG?<TI#YabI]d^e2F<5Qg#\J<90]Q=A3&IJ&&9(0-
P2SZ?,,b:Fd3]b4XFHJUH09R^b6/6HcG5e+K1#F-.NTF4^J(dMbf_6B3H:He384K
PN\FD:FJUgAc;FJa4CVT/gZ?/SVU1[(b>V2OaC5]ECZQ9.S_/MB0R-W(^77Z/?>9
(DbKR&c+I&71V\UMFS_gTg.Ae:35)Z,B:URa,\=>0@DcLVT4N39#:5N+R0KA/?6U
cJ>@LP670CVR88(RgIW;@b.I?^IWQXHH;aT]XR@J53#98KbWV@LdGQ8C5SQ=9;FG
WHf;5VAN#3[AY8BP@F_#<=98QXE(LG>)@YBO&569CZ1AF]SQ=,D/76(;25#^<,04
S60OK=/5fDW,K>0T=@LFb)6M(g]SG<&+660aI+23MfXA2J3/TG@N.AAWNY>;AB6X
=&(Z1=YH0(9@SeQA\&=Q3=>L=OKH[:S^=DW?P5M;F(dg0>LENO(_9W,@EDT77Gf?
VPe,FU]3_)X2732d[bJ640G4(Z6;<SP.BTP0;7b^>\#1UGOSL_#LTaKWKg^7:f_f
^+?1N?bWa[66eD8c1aF?M?FZ;SdXUf]C1PJV?;e]CJTgIBXCX4>1HaJJ&67X;VU3
RTaBZCTYBABe<528bI8\_SN^e:KOZ4#R6.QQ_PN6J>M:55LO)?FT6#=3P&ZM0I(8
<S0<)edXHA#->5](TQHT4U_PZOf_P))2&E+R3;W5XgNW#RQFJK7&2Ya+_;ZZ#RL<
04d4\#_)+66V_Rg+>_e@.6b8<:Qb-E(dE>Eb8+gGPdC]0_F+=0R^W#JH2^QUXINU
)0UMS:]Q\g)XDd>a5P&9BYf0:dV#S&N9a1NWPKS;SY-+5cZ1-PNQP9ZJ1V/2ZTVP
c/bAX))>LNeFZ7a)V;/MG#KC)V])B6I.@&V[(ZRTa<M1BCO>b:@(QgV70:/>LZ9_
9E?#.C@c.:HPEe@0,;f40C7U&,UZ/N@S82\>gPQQAC>Wd_8,G9^#6S6FM23U)NQV
-R,XH6bd2Y(PFU1:4]D/8BJNbYWHc2G]#WQ@1fcL]5?N4750DD>ZIHc;Y,[D@<6Z
]9+K1T.;;aW+E.?\;BM.T<N1\A/0fU=#XY@\J_DPNOdU;@P>X-2ga0MY1(+K6_Z=
>2e_S-62e2]2(a=DF#<cRA/Pc8BDPPPN:UOU9S<;9L3<HK>1W;ceBcQ^@ZNa@5HB
;8]e7J>/IX>TG_NXe.+M>f2JE4bc^@#d=)ZQ+O9K&D.J3249e9=ZYO6)>a6AB\2[
AK-3DBTgK#Be7b1Z7D_8a(,@&74FT#]N:#RB9CeHc[9^)+cBIg/>7A4M;,gX1P6a
1.Hcf><#;)XT>))<Y7@f7I3<40HSD#NF^^5E0g.fHWcWOg>>8ecT.,4:9cQeX_;N
BaYa/0&0R;52#0W>(D;VHIXR7>Ugb[d8PRPA:N:MgS.07YUQ0/&8M7=P@gZ@=^Z)
9TC-?LM8S[9gK4C[Y#6fY<XRCQ6&^YdMeOFBO4\]?4-8M9CF^MO\<EB.V,+28[0T
Ee&S,>Wg>E7\G[JJ2IHF#GX_RWe5-<c&=-Uc^\F9RCN^-c6[QA]@@Z#X&@;(;[FD
8=d<b:7GQ&81<JIHIg?=?aYZYgK^&H(G@P2.VIWX=NI[AI,_E&T\Oc2#-:TKa-/0
>HVC.9?+8IfI6<g>d5bW8D=LSH;1M_SVf<d,3e3[[Q[I68G_PIIcdT:fKc=@X@<A
B6_(INF#7.6+a;.aRTV3]DQ::1?fQA6R/]-V]S+8\4M3B[fagT@Z.S6<&DA?X2JO
D82?O):]548NB8BDV(Ug&4Lb_aIHQad6[_ZW3^;YfRA+X5T\/^+#V-:3H.eGM\P#
fZ/@OSULC=]]0Z^7;]-@,95SN8BUPJUgY:PFEXUBWWWFB?A#NORG.,U)Hd/+1C9<
,&2UT^QBS#M1CFXC9Z4V@Te]EXZ\]+f_^PJ[D4IXSM/:WTgRX>KHX@RZB]gJ&;(a
1FZZB6D23/=;J2.ZdPeN3d^V#+f7bUK[G<=&G4MY;F6(EGfIJ^8ZR\g6O;P>H+Z\
-A_Y[Y)?f<W@O(N5Pc4A:9XH:Z>e0e>SFBMd8NQ=OJBBAf^&)S)3-P_XYN3J^S@1
T[29?L0BdQ(.-YN[U(9;[@&U&&cBPZB<QY<]^L=X<]-S.b(.@?5<G.SBFY<NJR7a
fDe:Bg,Z4K(/=0bQA/Q)U#?R6MTY]1)F_HNL7W3dUfKMYa9f/G,9H?a6S>&4&-?Q
BLV86d45@)EbA6FEI?[.O\41=<8)Mf+HU?2FUH\#5->Y>A7>G30SG\6DHa:=&PC#
Pd>B7e1J33Z&-^_XX3IJM8S@2/ZbPb4>\L&=[f;FNYF4(W5JfF-d.U,d@2a9WM[H
[?X[GJ.JgH^VUc-((;1]GGgU7BcL]d[2MI4,g/D:4e)GZaC=HAa,JDO]JG_EV?e6
^9-76/\9D7\8HDRQEV6I-2bW<^94K[3FT]_UZ>,VR[&^Md.:IP>_A0ZD=(/]7>\3
6>>DSWONO@1Hb-M/bANRSE]c@_67Y@SQ.<K:K]J<;-?UTUHDC3).dZ5:RQ7HEeL7
\25JR9MdKbR3FXWVW2:,EU\LK=LafO?HJ&_R?U]a)M?K7/DKefT,-D8;,cBDdZ8I
;0_5],Z;[:K^>g[X;9A,V9@LS^\g.U&X)2ce,gV/F/,9O;Wc>]>M.:W@=K2Y0(3:
-SOOaO4F,7VXce)c^e53D7R2bMZ)5^ZST]--UVf#(NB2PeHIY=+QQ@MY1g&Z@.CI
TA3+LO832BDS,(?:S4Z^BGg]GN@=MTgd=1]4/VOPb+;048)X;D4XM+=2eS[&AO,(
^Q;XaT=R.^YeS-1D?Xf=.?^P?+RLO5./bb0_GfL..A^W.#^_+F2ebN5^[Q[I=7fO
D30AC(De._Wc,1O.Jd/]&J.#H+LbJ#KC.bf21<W2,O=AR:O,R#J_@g1BCUM#RQ4L
+@&B5ZV[CEPPK=e/SLHG:_0;(\SY:=>?&R:2fbB85K]E3/,X,Q9:dR;HI)e_.cTf
LPDd8\6gU>dT94CA0)S=d^0?>T5(U<3E-]e]c:0NFTR6H>;f36,&;8/LUV)=M4+6
.(B>>M@;JN[U[g]&H@HRaS)IUa8SA&JMMV=Ta=^/2SZ@1D2&COZ]S0gQ6BD.LO\=
PYZP@>+LZHE1N2R\d@BW7QQLW(R.H5eYg;I2>QbK3PGSC(TTdKE>>V&+7NA,<fRZ
>HG##774PI7cb6b9TSb=Db[_EHH76+[:4eTO;Ha-;O)KLP8,)cI_#XQ&7d+d,)0G
A\f=ePcgNU6Z/10VeE9ZL+7JNJW^=EGM:L]c4U4ENaB>1W7=R\CPN#GZJ.H]2BA_
&)EE1Y,edLbRM07M8_dW#Ng9_eOD4^<+EALR.@2KW6(KXI^DaBdNTGU,0+IRXM8>
P>#_NeEX9Og(PeGO?4b,V0O(aLBO?H;Db.8R=>CEQM[-b,F,cWE1-?c\g@)X,0F(
P[H74BVgfHA;#A1N,C2c/B;e8,0HZO[0EeI](bZX=V4.PTe@WX-)_M[;1Z83W&ag
eg.RYJ_E,N^2B<YL5M(K=8]a/<09P8Y27cI@D>,Z8eT2;B(CgeYN5;JCDDA\M7P?
(fZO^Lg=3)<UH=<H(a&LR+Y8H1b6fZ=3@#=3K_Z5(RY(Ng9a3)GcG:)-)YJ;e(?G
cc&U[Z,Z_U>UZG]7]bd80LV=V)N?@]GM8W883V)?5@^^dLJ8+@^;V,8W+HKL^S26
9S:;@=@_c5SI@48\OF=+5g7[O>g(I;^2B^IY]9./UWUcM/ZZb28YV[>(Z?E2CH[d
,)/55+#,PAbNVY?>I_+GeIXbL-M<==D<e\M6Bg7@U;T@1S@R/JC]T:?<gT;P^]QY
9;g8Ga2Q/U#f#O-5;[Q+^/:#=B^NEH,EYX[DQ]Oe-?Q?T>P,<]J\0NB9,A]>&X8:
<2:A[JNB5F+;7Q<_9ZaZ81WS)]5Z(,KE3=.dUJ.>:YFMI09:>BH&?Y@ZW;]R2fFR
OL(LQ#@P4g-c@?.VHCNAL/N95[g+P54,B.JK()M-W^,ULI<<PI7F^#2),>H9WNXG
\3>W02?5QT;UX#,UVW<601[^6fN;LIa9802]=cPJYV1>gRCG<I=[XU0)-L@>#0Z>
Q#@?7=\+/)d;MGQ97Z/30P;cLb.W66K_cJ]WW(b#\X0#CYHD);_AQ#(bA:1f##\V
1WII3?@DTWFgf2gC#dVA>M5)H4QBUXFA8K1LFb71^81>E<dY.T=A6f,)B1Y;WMQ1
OK#-TCJHd&fHa&8(ZY,;Q[J>@A9SBMb=I<TVMJ3#9gd[7Id0bGJa]AeH#FbA6R<B
Y3gCb\@<NVMN@\.MTB6A6DeANEe5-VB-V8H@e\MA.8#_Mb>?;Q8B]gJ)c5=\M/c#
Af,3OAbRZE-6fP4JS9ZAW[0KdHA]ZR:VBPGa4Pga,ID\<[OEL,6]+K.H;cUgTPX7
R7BF^aCe#eC>aU;/39IW6)Kc9BeNRCW=BDeOGea=DVEQ((:CP9QHT4FYLGg.PI#[
](L-I7X,GEg2E1PC>#RYMWBFee_@/d^;aK2Bf^W?PJ(3Se=e47WZ8\c--8J@S?,^
Fg;IG[P#[<14^_bNd>6LI87S6N><?M5ZA&/,WI6M:EF8E7+(UC;3-X]^GN@e?17N
KSG8aW+&@QcA^Vf4\F]291UU,O.5501;WE:F-KJ;c-T_<2,dL&8bCEP-<R.gJda=
QCd^b>F?_[)CfW\JAaa[.97JEBc9cHO\\=VH=egAF=2>g]8;#agG-[X]/VTZ_Aa0
\\:IT^>XZPfI?JGLb(Y[3O]F=La9_SG^FV_#ce+-.2cdB2R9\)6VR+8a7&-PI+>S
0=M9JdW?_)-=L#&0/]3f^fA2#;1T&\1IEE=8G9-Bb,)eCM;2KfY5[5/;\^XNeJ2P
Yg@^fT>9c:AV7(]cM5VV^\f?c?Z5AS;;08a+9Nd);JaB_#V_0I?UHF/db53&Xge@
P&^5KOXCL0HPddAcU:4g6_PC]L?5C/P?/@f[WT#e_>M0GPE1bZ@FEKD0@#N4^(@b
);.A#T\T1BRdg4MO3)Q_>cc2HJK#NOOfED6)_[C1WS^+JCH4(\MT@@Z7cR7FMMA8
eY;1308K)7J#HADV1DI]=IEDf_JZ3(E3^/].bB^S:2Q7K)/5E4E7]T^Vg<O,/b-.
CZG<<;,R7(I86Ef@Rg0Xfc?LV4Bb&NbIeZ1K>K^^FIGcUcKQ78L)9HO4_0JBd6g;
dGeV#QTWZ)_4&VfZb]DHa7?77\KR<:]6:F+ebYC#[\.>1,_]NH4UL5:OAQWG&;:a
.&?/8/-?ZAA@aE(:H)R??KHHQ>,d\R7I(Zc5+T=LJMIGFeZ,-_067bUb(@dE7/ND
\6[+c@YIS+G:QH2cZX;NSS<EIg)E[?fX2(dUaEU=0EBZ&>S.L77aHf(83V\OZ;d4
\PQ[CKA1DG/II(G]#PI#eM0He(2c37>bR(XGb;@T8C=:HHcY(agJG\[G8;aMb^#<
@;B=gf[U=R]Y5@_ESH@>HQV8d84OBOH^A;-26UFDe\S0\2Ba9gT@XVGaIRB=(E[V
>X25/8EEMFN)WA5[b.W<-GeOA4-66/>(E1gH_9OQPHg(]-R=2dA-UJ_=JF.P^/Le
.:<X?.W69&e=+TRV.#:55(ZV\eV+>Na3+#3O/Y#,C[d7=79Z=S4B4&D#IN\_EJ@J
G<4Q;7T2gU,\J#^[^O#&+G[M1>^)Q\@HY_YW_<b72b(,&]7bGBaY\AZB7dSK<U(O
b#UAL88g=cX_M+0NNDaB6+QQJ:=QccM0(-]Kf+37-c9Gb4G?GMa[G)YDLMST[HB#
9g5GK>JUb;O+9DB>IVWNe5P6S?U.41>0&e8>AEU&OA,V9AE05NXS@)>5O?5\b50-
TKf#U(N-[e.Y4D;ZG(AZK)DVVX.?5cPO)-e+/\;^Y@QX0f3BF&IJ<K+AJ-fege,P
b2LQ1B18ffQ#a=4OXJP:+G/8TQCPI,1\P>c6>)8](5+f1#^[7D3U??4[)FN;\3S>
8(J>bDgPWTC),VZDY<N.4aSK5J/[Z@K-/G_;IDLNfP;?KC+=gKX6[0?6YVcg/3A0
1I\bJ^eD,9f:<[PaJULQQ[P)eHO9#8RF(L[9>#@=4aeSTScXWUPO7M^aLfH(Q37T
=;L8g2UO.aB2_1ab>H+-PGHTK)[F^aNbd@G)T9162a>D&b@&JWK.X/HP_8IDd4d9
)RcF?K+[#g9>E2R)YUD&IHOA&aSa^U?DRJ:+-T=?]\^]#>1^;bXS\dZHVS/:]D@T
)9\I<SA=1F>IEXQ:]IYE,78MN[SF++\f#-O:VN2Ma2P]XP>SY:gN_IVF>G\-ME[6
K_c@RH[cDX/FADZWcQX-->,J^1KOZHPN#>NZ@V_g;0+Cd<CB4E9D22XS+5MNQa<3
XO<ZNf9>VTQ4G-?e.ac83:K2e^)c=e[(YM-gVC95[K&)GKV&9D1;;0WL;13Xg_Sc
d=WUYd/2U@^(9Id?51N@66Q5^6E2f&dHD-UTB73A]NB?D\<U>YBK2LE;26PQ(O/.
,Q:DGO&T1?R<9?M;Sfd81;BO]gIg-W\?8JPO7H1I@MYJJ6A^8P]/LKR4FR#710He
F]>6J:)cXX/;&f,C=GQP9_S;>\48eMFYfN^M\7^7]]:\gU&AcQ=D@L7]MK4>FX(H
)W2(0Y(8@(1.(:;CY[LDOYS):AK[Tacg.A#e1-J@O(0f+AJMJW91\DXa#X9CE/NE
;b@H]QT6.IgP3G-+@F&I6b+-P\U6OfN44^HL3cTZeSMa4W8>2)TFR5>F/5fUS7/E
fX&Ff<LL4_:P;/8AR)QdI?eB0J-dSTW[[3,gJ.E1H^I#FbLg_1]F/b=?Z@c5TU5@
_XZ24/[PB6MY\]368P7E<YYGFP[5Q>,MBfc8/TMHb7#J3b2LeL6(-0A5AS9BVX#E
4)&OF?dC:Ea;LC1YSS^9H-II55F.]d;Ye>,D&Z:L5g#+IH@(OZ\.I8=Q]9021WY)
WXTVa?CQdNe,6=#(Y+#8W>V>,AGX=&A3.RY\_CZQIMR>T]3X1;_>5fC](6TGc#3O
S=fPfe:1bC2<Nde25/eEVgN2^B4WDgZP4AB1FW-.=\^([0R9CP9#fMWLC&aBX6,V
\)e<69;W9:\8:@FD.b.+[HK=BPZKg6)<_/XgS#W037X517[OCS.?NU)AaB?d\5L?
25T-5X.G1&a#NMY^O(LGQN(c->.BY4MR)VcK(fS@2H\4\)5B&Cd+a5[E>+29@SXS
;()1?VLKEPU>cFY6Z]/Ke#d5MURX1[:B.^5^O2IK78&OBUYC:V7GXT+&Ze#XWSQ[
?UNE15BH7VQFBB\3SP0BHT=KK3=XfH>\QK_Rd?,7QFL1H3#PE39VaX/BMTSM.2?6
0EN9VbO/(8J2cQJO/(@ERF-PR#X8R^K=g0=e[,1V7+<2-g_P#=#ePBIR;SJA[Z<=
YVN/.V\46-5&:)f\_JC3AP1F#C8F356_BX.HC;McJYEX:>KN)A]T2IKHW_.Wf<[W
=e;\W0)F1@_a,3f>XHQP8QGOa=b+W&)QOX2cLf=F;V5RdH=TQT7HV8Q)ZP4QW@EF
DXQ?IZ7<:V0-QQD&6g9TBNLOf6_W?AZbC=D4WV17ZMZR\[be0>/R5&KSO2LPf1-(
7E;c/[W,LA3Qf0#(d.Z\?)?ScRAJ5:/YaV8(Q8@5WNJ47O@09\EI;-EU9AK_O16)
H=5XSg>/?.0:aT^8<ZbXf:)GU+\[aI):g^6NV:G<SQCfTbd?EI6[DaMX-V[^0d.H
H8X^)QOO8-A.MY.^JC[AQW9CK,6,:CP2R_7A+?JZ)AKP0a49BB(TU7Va/\-?6(&&
[3?BBdWKRV8].7+ZU(<S>TeKHM:+@[ZS<-GNN_BP,&Aa\105c9.JbH=].GM+\;8.
LE[IPd-&6#5Td]_KEDeG,ZHU<Q>+>S;Af.#:2PK,2F9&<L^NMII?Cd(10<YA0:a2
Y2cDADEUCgG(^WX_24;gac>bK4ME-Feg.+2b1#HC=,9(CN(+?=;aXfL@ERCI4P3.
DZ2U2.MD\eNW844L;EE9V@\[@MJT_6+R8H/?GDBDd(ff.<>fb[W^,O;B&6TNOQ\W
[QF<5==4I@ddMY[+\=PbG#6))\<DE+Tb>):Mc?]<5/>F6d,<>TPOFDOcZ6,;(?>:
+CfL-8Z-:6CA]c_Ee\]F:B0P5D6ITPITJJW]D[ZUaA><?LT9acNU>Z>SJ^66I:8Q
WNB7UBJH^fa?^HA+=3+W7G<&7aL_=_9^#(;1=H4]ZTL\d=d<Q74RZ4bG(VW6U8f4
)-SVMa05&_C;XSJ/,ART-#WE;]LXJK-.3=AfaTU#:3VBAX-2fbSXPLI=Sb\ITgJ0
&aMS2-]eWCZY^UL&:\GVb-ROM,,P:^Hg[CP0.K1A\=F0Z)e.I.OgAL3T<K:\C5,M
DBTT1LA0UW7S#g1Y?H(K9/<BB<7:VMMcb.NM;##S22SY<8fU2<5d07\)eRaZ94_E
[.QDA?UYS]^A^O8:_#6S6BcR+7V>-4CVTGUNXRI&M#S:0g^NQIa,:39&7<O+?,,Y
#>,D<1gP))UMB<+/U/-CZEM\L<JR9/IH=XcCS_[b1KgV)),EVH.VXV^&JJVED/V(
0R\DbVJYXZG_ZS.][MJMYdO^O5)<a#DT\X?N3fN1a?4be63JQ/d]LV[OVZ[>OD[S
DafPG3B:;_K2HZ;_P@_>HXJ#T/aX7_R-17>5<ZM^QYKCFJK2>--Wf90]Qa:b9f_Q
I6e;1W&Y8a@B,MS\F,Ec_&P16E.C8QA,5\94G/;ba,0eV<#aaG]JWRV@HbB6I)f;
&[9?0K;_QfQUK[^g-LZ=8/9,X=X-4Sb2Ue906G^)Y=.S,C+B4_M54WU<</L#I9-Y
K,?@d(K:.=4D<UBg-FN9SX)+&aZ)K/e)/[RNFG1N8Wa)D3&eM+P1DMQ_OYOAA1JV
+,ETU/,df7#fJ.:Z&8^TUTI.E;9HBM2/9^2Q(07_2)IJZD6f6C+#AfX#9]K7IX>f
J;CONNXS#K>8F.bB_W866CH:JSfd\[MQV<M^<U])8Z.^)GY-BXKEBIVP-N0S;df)
<@W15,PEaNYEWf4ILT5MN^I#E0TTU(V0QGGN@^.Q&<12:gEGH2UF9R3B6F8MG\:T
80I]-8744U:&5-DBSdc(9,6-fUV;YgG8U9/5P0Z:eFbB7607cCQ60O<.#XU&9gKX
;050#BS>I7a^06/gO/08@dI9W&Fc)8PS>S]((Q&@J,Lc88J+a]\CI=NZ9aCe\4_Q
R+<7[W&LG?>cEN)^4^R0dHI8SZb=6(?(Z=#(LUR6KS8-g2,T@F^964c4.Yb]BF[G
[6Q4f0MVPC4>K?<1e3>,WcVR&I=#OPH6=R;1WV5ABV9G3>8VGaGAIICL@8Mb@cT4
.1ECUB^M\9c,[=68]gT+#3D:VK0Fd^2R2,?7@G<B#5g;6A96,2>IO72FVD5TS^@D
#YUTf-_5)RCCWKd;V_J;4H\LFB59JK@R+2^\VE<e0B<+_?7?@@8>+3cc&#.;7YFF
DO^+GTdZBG@dEG.E535^<[cYH)B&GQBSWU,@8-:NUN#)Ya1-Q?SON)>f\6c-0P[c
]\)^5<edKFa)gaUZKZ#OZ9AHd&3G[b#<-C]@M3UMHH6X9Cdb2(T;W_O9-;]F\fc#
4W=+>&6@_Wc@,aL22UX2:C-#>C6f8eOBeGZM?:dAC8.)4dI&6^82^#FBVZ0MIAJ,
Id)11]]7X<c9_gJ;4?KG^^.<#6^9B,RUK^L:T,O8a>@HcN]R4\AH=:S#GCEP;bAO
?#O&HcE8Rcc,FE4T1&K_K]d3/4gQ_b\NW>YV9#D\RF;+SJ_Q&>aJ,VTD7@IbZ8@4
YZ<D-U?1H8a6:_AcM5CL:E&2>XEH/fN89U+Me8,J8=4Z/GS46>?L/^?ACA_OHS=e
5IGZ=5]<a0P[A9f203AMG7G9dDC./A[f_.=d-A-Y4?aK@ga?,[W9)TA]ea]9FAcW
+K=^a^SGKObA6OY,G\/&c)]aZYJ()eS;Q?2JC;+TO;=4^W,&#3F)K(W#XDSfE^df
^9Kb)<D;7[7gM./,G-5[W?L;J;]5a[N/UM.7UGQ.8+8ZB#/LHV.W^C;S?&HR.P)g
5]Z_-dSbUOXOSe>4d^O:=+Bf:@f^9=K<X^Je]GF/[QJ776S[?)^J]GG0bW>?>;V/
<b]<HR_;X8Re;5[^@6@@KJ-1G^1Y&X+:@:7BB,H@5<W32@R;O0D=,#D:-bYHAeEe
82e<cY\Y0FHTfDe7E/=:&T0I[0H9-fU;HK3V.TM,B9^52X::(^-N3.ON0C-d33Kf
3>T7g0IT&S;Sb@NPe-+bC;Ef6g\U3DcM=@c^<#Z2/L]U43gBBFL,1#@7>N)eb.E4
a9_M<EJ]-\,7K8b-(ZOB@7C21GQF>W\OPTQE?M.6OGI?U9>)TB]4V+B78Z6cBYBX
-]9,:bKYaXWa5dWYFC2^XY,/2]d89KAa+DW[e@\\1]SLCb<T:?_/LfTDL;J\/<^e
(Q:_(_.I,7H\A@DHWO=F\a0Xd-VZ\8-)B&>1J8LC/Q0JJZZK+F-XR5,D[,&a+S.b
RPT^AVO(_d2]F<eA4SfOIVQD89T(LAR\DdbC<P<AYV8\&H]17e<-M@KQC,Z(a<?^
X]-R]E2?eZY5_RY44=)]dHfH3^U;c=:0FE.FIV2d/.ULc>Pb80[HM?6g&T?B<8(f
BK_=Y)5:91RT,RX=]6&dXSedB[HfTP1>Y=N<;Pff]Xeg5KaC&K\e0):TIg1?;::K
4;,.I=E?K<>=dT1De_RY]&Gf@RFAXVKa1)a+f5RO,[<@[;\DD9_<X0)Kd_4V)9H2
47WC,]I)U[F#aY>WUAFZQQBQ@8??:N&/fX?4VW<_-8[_S7D^?#bO2@.M2aMJfXK6
:Y;PCGR+ZZ&S-@e5aDda<A=NS<6+_a+Q(666Df[VaMeRffd_KU<S&5G3D8P/;.)a
+L+\&Pb#B8>VL<g:<(V&6QU/Rb,]H8DCHN0GV.bI0+0O<]d6#9X75<N>0:[P.UXS
W]WQA5\]9X2:\=Gb#L.8HA#0+I;I<gQ:5X#A.dB)1R:K++gWTQNGG4WFe^4(+LS>
3>U;U2[K+Ne0PdSH-)8fWc&NI?.?3X;T:>^JV#D:P)4dI]ZM5)N;g@U^N29O3eS.
U]7H&;>aH9\);(R&3OWO.WK4f\PK;K&W,ZB9-AA-;baC3FR3ZB9)SgN^3;5T7.3H
E/#(03A&=W/P^<D2(R=M_UT2@C<3ZQCG+<Xd.>@2bVgYQB=/-\E+H&/9?MQUJV2I
TSHO--BY)39VF9;#99#E,>d3)TY6<L9S\/gI=_Y<BAUX8RN7=McKUPX.7]5\K)=:
IA4YF33EZW-:XAHN-7&:TO.YX+ZgA.B,DU5&0^9E8W0,b_-<ORMM_QEH>502UE+Y
3)V,A&9VT^8Zbc=UK?<JWB[HRNJ>I9DPVU6K9RJT+4/>e&BdPN,Zg]g-R@,J<ORG
56J=F-5=Na5,[J(Z)O<GXe-H&f?6ZIX+LOIAB@JbZX<LG:.3#KNZ.M2-:c/eJH\)
8((PE=2M6cAA]5#\AMgLROF:3E#>4:[e86S?RY]:e0Id[0H@OS6+W7c8:JDc31?/
9b(bR<0d84[ZY:WIbH1R&S-L2a:S\^?Mg(C4[A&R&@]>BK+A+Y1(=1T_CcG(f>L4
:K2KARK,H,E<eb4V:B9.TP69&D:H?/QC3A;QAg/O)+ag?(5973:(;Lb-9VFcf(HI
;g2BKR2?U^YCCT5E4-CgFZ7SabQ[WW>0RZ/UHU1=\Z:\0]1K),\]569[e<&QGL(_
IV(W)eN(b^D:HP6S1BCHRA])db&?W&G?Hg/S(MT[/<3<&-;]EH2C3MINHPcC#^ee
_[5//WB[FaG>,+26?38:?6]71cSE9F0M49GA4W5KVMCb8.<[c[g4@^W_^[&gWEW)
&aFaUd8/E9CK+DHSP:U[7LZ4_210e<fYAVE72Eg1dcV3]KYV-/bI-SC2:9Kc4aXW
]7KbSH<]gf?O\cYI@dMJ<AY91?/4();)UM3JPX[5.MdXSJc33aCd/g-M,Z]?WFI2
CS8/cQf<.JHW1\dZTC4HV5)>?1f_+2-,].A]^DeC9aWH<_B^)&+9Z^_/.H-Ie(81
U^XYPf+LNHYC.GV+E_)M;fPM:/Z&V5Q7dSMVQN\@fZL>Y_Y9<cTgKLPHgLISE53X
BFLDb=\WLM;0bKEE[J&Y.N2.@1NE3;WZI[.;d<4+:<&8?9[)HW)T/WbB)\D7fDg9
+,.(K9T(=8)YAX-M(Y\41K1aEF@P4=4:ST-QCQD=E.<5X1:/)(RU-]I+QV&JD^3Z
(Ee@?Rb#cW#T-2[HW6Z+9IRVaHXgK=K?e/b?-e)(@JD>S4Ug@LZ^?WIbg&/_0.S(
/:[2B(_WMCWI#4-BN+YMNd?^LR;:]]?_YQ:KTQDf50)SW#\43G6;#9KV]O]Lb>V/
Of\XKPDPM#27NB)B:EZKfY\2?3O/=KEI1-U0W&S#P?W3E.&>c63]1Y?aEL@H&Nd9
EO7W=\[(>S>GE[M0dcN(@1#@TD?O,H^@TSaK;4^L#WG@VJ;]IG0<]-K4JD<c1?L:
8J6=fgRUd1\eG8I;@@-?#>C9>GJD.ggb_0:Q0MY@B7U;Ab&9?afGL><5.;>]6E/H
@X)g@;[U8A0L>7J_[)T#c)P6]MOPRV))/F-gSC:gSW7();VC4&O=_ME80@6BIV.b
4-bQQe]a&9/XJO85&3^T[NL4g^5-/YBB;3CAbA:A1>+X\@NQ4GK4YFY?5^TC55d/
KWDRDXeYK82e?2aMH@0d42V4<bDQ>aUSbR@/RZ<a_d<e\X?F.W>O&Pde],bCQD;e
.2>U8<g)#T,TMUYVDN;XN319U+bJRb128ST4&cL?a+g++\UBI?:WU8POK4[R)7(1
,E,X#)+?:HB.6DCGF\f^0Q-a\A<9@A(8#YO468>5G1#ABc7]-?[G5>):&J#=?I,R
HQdf_9M<NXSAC,#cgQNP>1D0#fL][NGUEM]Y[0;=R72+QQaFENP&4VVd4N;W,dH)
d&>^N0(&Z#A<b5?(<(:0Z;0?N)]L)@HY;@LP^K[1EOB6b:[SVA)@?1][)?96O;1.
YDAU59L43LH9U.)8Gb-\T:ZP2Z<=;AJ=1SPC26OB=@g\7Kf_\@L5>0J2,NI6D]FK
S]@A_[-fVT#,4[OMK)HMg#+\gBa[0S(6?>[(FQHC=P@1MHF2PIFI&AbMc,T-_e^F
FNA)F=Y28V\CTZ7<g\?B/<L7#O9H5H\VPe[(ZBBc\;RXAI3W4Wff_XHA</1[(Kf2
>OJOA=MJ_YM#?),1[COH>VU@=6M<V+\FG]T\fObSS<d94X9a&AJa0YeCOaMK:/QG
XK1WaT9ZP9^.<:E4Z)-&)\\IE8d=bY,Ag8O\VH<\cS23C[3=L(9=XW=DJD2M5GC2
SCc1@GF7Z?f<9ESg&XbI[-KSX&\).B0I85AaE#.4\EDVWC8^HGF(=<EP&9bCB?/3
[B=]&FR=V(,fQOIR8>G&6=_4&.8=CcbNW4W;E(6;[3#_5N]>(&7U<d9:,A,.IMe+
eSTC>@><\U)U-e\5-_U:adX(->9):\,a2(3&BCKg##@+IVM9O/8+/J-b:?\-I.U/
E9-9YKS,Y_f0X+VGgF#D9XVCG\a#YeIF?Vc]Q_+^^V(S78D6:IJ+^c_G^..]-T;_
\eeNC-6a[PSHFXccIX418<@PE3]b<[<&:)6U552.KWTMaT8UA<4LPQ,2TW#J7Rf<
CAc=V7?_3,+8OX&cOL@KWJ#5d2\#a;D2Ld;6I&;?g]U38-]UGB.OCQ)D)XCM[=E6
([fT?7AU2d6)Q,P+gP9K)@g>-cfRI:^=:e2].DeJG?3.)[a+gIFY;5A.8A]X),<^
?_AWU9941?)+FM-YUZ.@)cL=P-VD&4cg#T,G=R]OK1W>-dYA>JX6,e>#IdL]\KQA
1943^).LKO3Na-10#V6<U3+]GN>CYVBRWHO;4TMge4YIf.#2#PHVB=O2.^&L_N=^
b/../H<)?#<Z-0(3e_M=7@H2=0fKg&?EYY<WAcWK5;]Ob6GM#;DKdH>BOETL&U=3
cJ]&E500NRUV@UOCOSAO0=0H#_EOZQ0Tf,QXef?A)89(<@c79KO<Y&5LY]QAF]PW
c8d9#/aG[-BF?UTHg8dWAMV(.A6P7[W_]6+1_9G;3^e:?6ge#F7>KdDD/ebUAE]e
=:fA+UeWO2J7Z?8.Z/6f&=C-K31VF&U;?&Eb&UO&F/NF7F\[E(AdbI:NDBU_]],L
I3&2GYU7=<O]7=CN7&L7+gK3O5K1G[;S<4]G5gQb&feX@I1E5U;]PJFgY#P=1<a+
-=,=#4L+5@aXNX+a(0E&=-M?=Z\a]FI8:^^4SdgYXC:R])TR7#9])KK_#CH8fOM&
d/B6W#=;6<4&O0;e6>7WdI3L3^C5BZK6Q&[UJ=6S[OF(;#a0T7ZHXb)aJ3UX]\29
7;]67/B.^:)R^^T[\7)PW(IL(\+)^V8d3>]15#+\.Jc&MG?AfSXOGAC<_H.F([Z+
_I0;9M2.>,D#<EL\Q>Xc)5X6];_;O;;XOf6C4K(P6=?d<b:?4)K4&4[043J1.\SQ
@V71_aK^_\E131Bda@,L1B)^T&+T>R11A.KO7<:OU/cZQ^Z?TLZ)6<]C;936a^W4
HS\;VKA/6&LVB^WH,&I>P_TO9)<F,>)M&R_:9@AB-f-Y.a>KC+[)?J2PN5ac_#M2
cW@ZfcOD<;YJOCP<SX2GX,DN1;[J/E=@B>Sf@aCE4[NQTDQMUK.Ef#0aOL1(>bg.
&FC;\@B82<.Q@/XA.d?-R.0C7^[GZ&cY0-KRMPD[Dae/X8]06g.S\Lc<VT>P>g9-
,VYdN^+HIc8^B:dV0]Q1>6XW[d/1)ST7A6.E\:2R6QdZDZG^gVX;@FDMV4Oa5)?I
\0?._ES#/E5VGVaLU--/Y2OdU94:_=OA.=;;PbYdQT9FRc13Y6K=@ce0QIP).[M#
S_/OH<<N(+2]=6#[\VUHK77?).O,PCUYWIdCT2?:UQTC1#1.P(aJE[Q=eSI]6_AP
\b7,_cPL1]D(TYMT<=8&V:dG^cFJ+.COA]dOVaG5Pa5&VV,J/-C5b#5.Ub^,EDCf
e.?5.O5#D+_XWJU;>5=U2:dc194;.[-XR5ZIRaM^f95JSEd<L.>^X3--LSDC?J^d
X)\_GF;I]A&O/Y0;(-]_g+;F76)PAL6L3WI,I#.=c]06ZFAQ;W^5I(DAaS_LE91G
beK0G29f&0c161^fd]6@0A>?+G8?@&&Y\1M147ZR7gBZB[.7T?F4NB8LZ^,K]g#D
4.OF27EdPHJ]AbY(_dbV+W(PSXY/dO(XU:J-EWe_C46U]O(+V>U&M/N4c;J<]KeD
g?CC:-+NO9YX8S&d9L.7MIRS.dJUQ0>UEOf364&;b<Bd;_1_YVHUQRI:TdceLAKX
Y6#00JBQbHY;0JcG<(TGAG^&T7fPaOQ(X6O:7&6A_F]E9.&6[OT7UCX4e@;c,]^]
Y7@ND?8V2QWHV>H8@Y\/Y+9>cETdA<KUPf+^VCHEL9-DaH4C-^K[?TS4DSNCd@1&
_(^P2)#GfF0P4)<^MOXA<(;0BGdBK_f,=:FG,3fB58?)JPP54&?^[4)ebFRLFWN<
c+_N7?LUJ:3Z)8MEAGE[LSgR(;)C[7Z<6>be]G:P1;H<_Ea,5T/N;&FL:7EZZ,\<
>UO(=g4WPEO1bc6E0_C:c_bg4/F4AQac9Q6Za3V=.9eY@_CaQ)T(;<=@WF2P[-;Z
B\SLCV/f1IQQB.0dfe4AF.K?5GB^9UTHGda7FT9\W<4aU.A=&e\7CQ>fLI>R:99?
fJA2.BBJ]A@bG&dNGOSW#>Z1U:\CW65JNX6&^9;cG^YOD3Bd-@KEQTTDCFd-Zc,g
FG5<AGSA0CaZg)c0.^7Q6\N/>8a6LbD/@N9<K>[8DR\4RN-L3a:/9Y/A)1K1QP@5
EQbb22[BDZVI5(E/HY-=b)Y\8>M[c_QG;H2J=4_;91Y@(g^9>\G?9&CAYK^900eK
2TT[+7<c[aB-9a+,c?bXM=RXQJIIHa@L,>206-9=1Y\#[cS7>O+16cHE[-/8QdW^
#9&2Q.b]Z2,8^#3=[7QT9&&>-BDF9GQ0J.QTG?#>JVT16Q^#L\eFdZG#]Z5AO+fF
AIE4B3g32,=a7F>Z;;-2\^2L[5BF^&eHAU+#f5bLCQU2]YPDV@cZTJD]&AGR?Y0I
UceEUc&V\24Y++F_[eU9XM#C5:;?#8,d<X#]g^;.</#H4KTbE&:Z(dP(OT;_6c^2
@PfBaHOL?eIT#Lc33<@TC5>-L+eF8eN^H?XB.7AO;-&RK&=<_RV)L\_)9b5CPSS-
#71J_9QG_\L7C9A-0N.N#>E<W+d3b6W=C]6MB&Z9YHD7dX3Je5.>[G.LRBa_gH[4
QBM9FZO>:a>+(?/f[2Pg(5+DJ0K&#L8f\Y]1#F\817M?G(.-g@(?8#^/3?M\2ZK5
WS)2-eIa3PL>?fY#O([S);Pa:?g/PBS7g/IS;WIc^4AD]7SB)G_6[(_QLE?6)V>R
feH]d+JUcXgD4Q:dB>;ZJG/MeL2QXa.K@6&1+)[3RWA)7BFXJIVDL;AD>).DS)DG
C22_U7KfdBG802BE00S?]\.[KUEE5R^RdcSZ744UDA@gKHQ]7?fG0=F?fGBF;X#\
WgU#15GcAPWXNK^;N6O#]e?.M_,5ZFX)9eA;;/F?P?ETIH5[YD9JZdV5E?W+a(NG
PXQBQd=94b[-M>_2+?g?M\4FND:Bf3YD3\(R4G90&_J2,F+UAM5Z+AOU4@\TI3OP
26<-UG20G&9]+GQ8IZ)@a#P;+AIBYE7McY>GdM=MN6<[]f^H)ZLEg]2-66>Lgd=)
TWH)3VMPQ\:G=H)9fGFZOU=C9J^94ZM:J36;eQ_0H;Q?#<E_B\L\=BKTJ),0@[&)
GQ;&ZcJ[=[S0(W+]c0FHb=)2HP=X3g18f0C#&D/I-2&_CcLRLL86O\4&^Y;KH2B-
B[XS0E?fQE&D.(,5Z[)bC/>BMXNF;NHG4Y8XC)RFZXG41EU8F+J<^;g87WR\g.FE
K;A<\W3L^JHQ<(&E_-=FM).g73)>Fa]A9O>4EE^0@STW^-EcbC>L/Q&D:Tf/cYB5
M1[X12OV:7M^]2<a#MS:;0QQDY>8>6/D&\T;NYe9dO0J2@IN2ZBR1>8GDZ/a:/N5
.Z_#XO\L2X3/[bIFd4\)4#?J=9&<7N^DX5@FF8aMG.KL@[.d=f&?CXc(W-cga\ed
@2=13CN4-13_L2]S+.>28/<#G]^dVU[R^^&:(CgPIb3&4S10JRX;cV:?WQW,b?UT
9.[fde14NDPTgAA<_QIE:</NbI#D-:9<?P?.N\I1K;d?53T)&-M0Cc6FJ9>NSPMT
QXMaH;&g+L[>A-3Z7QTJIa&[(L\T,>SJXd(FJN._K4>Ob)^7+],dO,P<g=R+fb,K
\E:d6#35#\QH8T]-f5?Q,c,WVXF3[JBAR-#;#Q>faf\ag)-bR]W2a?cJ&JO.&ZZE
FZ]EJ95Cdd+.3?DV3/APbS();S97ZIH6[,R;,305=?M+CCb.RXD+<DAe:_.FP>EP
OU_0@2AVJ&d/R/<P?5f_I9Ug]_2SZM#3+1Y9c&)LEO4^ZReRSWAQ)M.I7TE8aXBE
d5L]Y_cTWg(c>gdUDUHN)67YJE,#I8?+KO,PT_:#LMKV+2W@.@Y^RQB8g;ad:BZZ
)a_TE.H]]7B:E&IH]fM-D0E^,CRZ14YIWD]B?ETHeK@FI/-DM#.&+3QgHM;O@\MW
G#@3Ad+UY2fWCS[>YGK#)X6D;d-#E)6IC9/DM6?5\cU^9bB[=;ZTR=a2.XB_=+H,
5/#V7W0(e_>@/T1N[2_.dZEe=Z9(5(>OWXcb<RDX9S)+Ld+-M__2EOVF8WR-ZZ\G
8?DJDS^Z?0-IEI+g=\ST(O=&A6TX[3^:O0RZ(dT4=<X;9FdM#?JAHTF5QU,8D(2.
W<Lc,;23I6a397?^e>7LWT4]0aM51=\O6:c0dHfS<SFFbf=H>dRgWZ.)9(853eAf
3Q/)/2Pa<:@+0Q[f^.BHMUJG(,U@@HJDPg<BAJU4_]4X=Y8K<RJ2IY+UM1?3d<MV
G;2DE;Z=85KQ6>D[)2S]SL#2]J-dG?XgR7FUC]<ZF(@Z<WVSb7b&X\_5cU.D_C__
CH>abHSM\7];6?UVY[^&SJDM=3?CgX,>RXU]OOP&/fa69GRODNBaI\X[LO3QDSA7
5_Gc_&:S;5Dd,Y.4GFLHZ\JC.,a0->^M(YT.LN[<K)\4^dKMNZ_.0_[B486I=6Q_
[Se8M(<\QILX5adI3V_&_]U,7LQ-Qgf)afFNGG?3<>H3Q(-/XSG[+O[c1GC-A,Z4
_9-_Mb.^OCZaa:PM]#c:9MYF<[]<ff5DB1M)9FX;\FECcO7ZIf7ZL+J#1Me?.6=N
ZESB\>&\TT[7>eS9/42.Tc\IB[Dd;He2<=>XNUG0Q0c^HCO<bD,)35L#>J0T6GdF
g9@=V[)3?JbN4<,TU+M\e,[b/-MC;_D7[._-EcK@cJ-V7c=8RU0[d[&-T^60[/9)
6J5>.QR.#f9@aSWXR0b^c(7W]_-XT3-R?JN&<(I/+OSObN)#P8>1C@b4_Q4/d6?A
.-cR_JJ@V<V#VH-VGgG,S[gReQ+I8_9Z_CMF+EWf:OH5X.CJ.T&3XH>e6Q6IbCC3
TYZ\g&\GX;-?1^(K_TXQ_72/5FDT91X-_8gOD<e)S6D^(T]8Pg8D5?KBEEb9+Rc[
PF7I>IXGgPg,^a-&HMPbDg6W\<3-E?)>@K[3QcQfVUM)<\D-,N@\9EM[30e7<^:4
@PgRN,REg:JPYd)?0#3-AQaMZ1M>g4\PZbd@I<\?aFc5#5XSU4DeRA.&8dFSH35e
Y7&c[DX2@;;P__MA7FfV/&BZB6(PYC#bfF+,O\WgE/&GBa33(ac/;eEVRQ0#cY3L
>gSM:L0TfTN@efK,,c7L=O.F9DZSE^0U?;\TT.V:-\.<WHO+aQG4KCD_31<-F_+d
cE:2TC1./CE#:E:T;:2/6.O.RX?Cg>X-B>[YaY+_bX,Qe9S1T/8DQ9OK)JcV/F1b
=[7E1LHg)cD@9WbQ;/aBQUT\R)e[4;9]aVaMbV)VG(]ZJP7cX&:eQPe.W21c_OG/
-Mf+S211N]>cN\eKZHWSG@b-/.^\,UW,5AD3V1>@cKM&/CR/N_T^W6.1=<..Z074
E85-NQ#J\ZK]F\d7>L:L@@VJ6P.47@0ecCe)AK[Ng6&+1X5G.WW9-5O74\(1G6MR
N9Ig4?;0.[,+MEeT&4(NEQ4AXf]CFUb25X[>W\c\P5YMWA5Z\6()G(8\8[fDT-=H
\#)5FTR2UBC2<WF0]-1_>HB[ZNU]7\B5/5TOJJ:4_H[eSO1Iae.&]NcHeK]?0J#W
.6R8XBB;UB6<5Y.1c0Q<,HCL]A7a6?N<5(L-8=#V[dSa?:3;_WfU4gAg#/-6Xa^-
f#FK+BAO0fTPT+E.Z<NP#1O/P&TELe;\;FJ)eRXSXNf[H7&:,ESc^QMCVB4W_7C1
&4eZZ5#.99B7[S[8@40_E(IFJ<]EG+#+N/4SY]AZ2c_0D_K>P-7XQa,DD]#fESDA
QA=;c:I8M[&(0&/<5eRW6-IHRL,J3-U6JLecWJ:N9C2F(DcC54K6QBNW(<EX.ML_
eEH6(C>MdCg:@e6f3Z=)]BWP9dcT).MQ]?,KZcJJ=:OM4f=SY@5,@7_306UeU2,b
1-P;gDQ56/L&05\CMYeAQ4]E^,Qc,8K^H)&IQD[_e7@W.8C=4I8MEQUaO3T7F]7M
F;FRg3)1GG>b.7f@@NF)ZbAWN.a.SD<a6_.R[4HS9[6;S^X9X^Wb(EbK>7I+ZR^+
;CACK8.?_/Q&UdV53-(ZR(_dA+5-BZ^L).CT5UBJ1F_Wg4Z:IfR<B[EZB<:6DV;.
U^HJP-I;6(253EWT8@S2LE?D3T8^7_>L:Y;.6[HPbQH.AE?)),7/@,UJR9/6NA>+
6fD2.U(bZg;S;[&[(\ND^=_=He.4.-ILU9.LT\EM(-(Df1ZUe@,.3)(5gWcaAR.J
eY-4?YdQE_eB8Qd[&SY4c5?&8S;&VUY_3T.O2/8<f]CIK>2O_33/7#=@9)8.I?G9
<B]fRARE4D8<cB.9,A+6;L3I67<XP<>#UD##602_1QCF[[?4>,H@W?.X.2L7:=M4
(_R-J;1K\0dL+GJAN[JWb89B.:#P3J,:BdcP3Tb.-9ZNYLA@>(RM/MP;1?cEdQ7@
J(7H.H\L@Gd.WcCMJ@MRd>4&Y)d6V=#PGY[,Hf7)A5T@I@[9#Xe<[4578gaX&9I@
V2DMPL@F38=MX#@BIbg[eGM.(2Z=\6=QP#3F#Md[0U@3MXH2-DN:1TfI=]ORQG-&
U4[X9#S:DeC4>ZU0@XK/]V<f(>^OZ>KcYBOV;d6DdH<8eO^B+0JK-a4Q22JgNQ5\
ba])#QLfG4:e3\0SIg-QW_67-U6.Y8@(1S.5eZG::2;S0,I?B5,PCD#+R@/(_Z,R
.@Cd&O8:#=_ZH:/.E?PG8>.-)]Ugg0BMK+O_B:0MD9.X:53AG5,K4SbUeI9<C\RR
<1bJS5KN7bC:KU2g,3,S[-RKP3H^Q9f]f6RD_-;&<FEUO\;+^He[>UNJ)W4cE>Sc
@>/\=BBaC@RX8J4:[f[E6]VcE[c91.5F@-7^5O4@bg?I-8-]F?(Ga#)=>(fIGWZQ
6_X6eBIM6W>1?D&#cM<J.g]e77f=Za<22a@MM:5]g^&H/A]bHIJ>:1XI_B)-EgYH
d-6>4Y5-O.KR(UR8DRca;3)d&8bcU_0<EY+aC))IC9cZ)G[+PD6LKTBLfFcV+3^[
aCO#]8ROYM4Ae.EEN#K)-I\5\6X+]Qg04@B,aOPa-)N6F=++617+ScEg2YL<J)T6
f?gFa63W3,f9L6gg.1Z:CFE;Q+P.J:V:g2.-?.4aBRTf8=TKLf]G)E6?(?O:CZCV
I#UAO0@_4c^L-6_f[/CVf<;&1Q6WET-e+g7H2b&SHI[RVV)aY0#;_(=.3E3K17gL
:b6L-.+H)5HU?(AN+RXZ(2b#4WW@M6.O^bYX@NL/TU5U4SX2Y5Z(^8ddT=CS;M5T
VA2&4<E1PVQNPD#DObU-V\?-H&1bXS\X#,@aK0GNE167VL\^FZ1-]0QA1\gPd/\J
HFWK08FE8O/6&/gfYWgO+Z]S6]e@:/eZCC1WG9^[7=28D9OKF0K.=-K>;K&G9UT+
FN]:gA,;-1_EY[:a(?HT3&IA7.:AHXNC0g2KVRd(SFfYe6T0ObLV]:c\C(NPf8#/
Ge73#2UdKB6/\NQNFW7dMggL:+A-[g&P?1d4Ja:O<&4SOf/8+OBW.-+a,18>Rc@0
c5M&cK0-J0c/G:B+9J.AV(P&,J2CR=8J]E?B)TA:N77+L+(N(US?E#?b/GCXL4L3
7g6E3@cYf(eGXbB?b<ePA(I-AV.Qb.D@NC7,;))D6L:F-99L)AQQ@2[+8&.Mb)Jb
2cF7\H\5g@B]O9<-80MNQA7H1.3[g048),NeJ1P[E(c[CLBVH2U)NPAgc^[(A)N[
L3-cK3?MQELE/&QK#CLH(6TI5@V=QB=6WMLLWg35cM.;6EO)eFY.)\FUcRQ:B8cO
ORO8^&D]f>@A\H(RR#/9\NOPH:f)L>>VH_FB[8e<=17YUE;JV61:/ef&<\=UI@R0
]K).2-&B+g1gZ3c,H,d5F(@=2X>D9#@A)0==ZKTC]IY)L3^(4ROgR0@:4B/Z<;0R
BeBC=6(^CIb68a:BCW3^0BU4#<3gCE\C(R@O-3ZME4Z_<[a4@;LbCfLRaMYO;U#D
K)cPY?2gFV3E>^9/55+a+?b:_FX#MY:gCL6Q3YK,e>>#<,5G2D\4D#,\9-DQ@Z&E
5MeK,#e<89S3AXL8a8c)O9A0fICT(@_B\B_03\4O#VOC:]_Y5(G4EGYgHAJFg.PJ
/P<SLZF14A7B?P\T-MGMPTRD0-<^]7FC+0VH+dBJC:>Z6H1e\9KKO>:#TCSb\XP6
9MVK>KMN_L7XGU7KWKcTf(KYc/[37A3MD]g=?>H+gBMAd?FD?;g,VXVYL\0gTRP9
A9^#<SK1_Q]#^][<:ae(3P(6Hg>Gc-_MD&d,)]PEB&2]XNB6@dCB5BRJ)UXbECFF
S1V+8=c>1AHQJ\ND&M)+=XWS3e.=IN8VA1.\bPb\.[e=MOg-VT^5=YUR7:a8bcV9
SITUd@T<ee-8Qd#G0Q\QAO#)GE>B.UZ-916;-CT@f)NVE/g5B-aMVcR0.-=,J\Xf
S\>M++YO#fO+-I6-,eMV7&e#->7D)+Nb2;RcMg/4M3;?+ZN=8SY(9Zg(F8AQ(PE3
b(K_I<HH@+3]Q\(c1&3^(a]CHL@f,<K]#P:HM=D\L#<M98L,Pa:5H+XW]VQWL5\B
_C-NYA1g<C@0)0/JW_)d02=3cQ=N[H[M/86d5XT<P_e>0a#?0QVDc)@fG9;M:#/:
/&ECXMgWG<G;0c:JU47V5]V9.X1DVdQBY_UP8LEC9\Y_XZ)(J5Z2Y8@]K8@^:[TX
\NA.gb)+2\H5A?@V-:NLIa0ED28_^__Jf<(D-KMaRb^C)gH]3JGFeL^fNF#Q/3Jc
G5(VXc^FJ.<gVNYS/cDJ;&Fe=B9PP-ec8Z/CB_+/6JTQ<=E[[@g4-FD4)3[NNZ7b
c7K@,8.YW(#Z\5JL/:JO_;>VF+>1+8-Wc:J[/g.eNa;c7cYgND8+>_J]=dRc0@cT
N0IRQ=1<.<#eIca=9V;Q:(XTdR68LTTga.U5T+=.IT5I2S;YG@6KYaGfR(M^/FN[
Yf^;&Nf5;7eBRVL[0JDRaJYH3JSV15-&WI#0A8+#K4/Z#GgHBFKQE#&M5/NSLQO\
<d@Hf.]2AXfK?g]A]-26&SE2fd20ZJ+6Z,5JJ7R9R2?36,G+-.;_1.e(=3cGA\_#
)]13U9Z6U4gd\Le@WFg2REfQ-QT>Lb/GMbg#J6,#B^+1/SaAgTIQ^8fd^RPNK0Ec
;>V;\I?SK^4/Y,MX1KUbded?NAW3Ie4/eK2bN;?>1>eA2@;SI)Y^,P1UH7046Re8
N..?cB=(>]X?+bb(Je(WJ8V2SDE0<QG0O2K=KI/fFQbb-A5@:?-Y^gQ=LT:G\M^/
aKQ\;Z8fNHa>H[KEF+AaT:\Z:1Y=2(fU92YeJ4\P/1M=e\g8_?#VW=6-QJ;(_.2/
,:W0D4[QdbbHE;18&-S932M3H4<6d^OJF7VTL<aJJ2&735,P=a=QOJ5SAaWGEAFN
:FHIKG0BA_O^ZMc.IR:7KOg+bFNbVFFU;^8cBWG+V-=AWL5)?LfT^G78W,\EW.c8
;c/[>QDZ-WD/,\_]O-DK+UgY(2X/^f3Tf,2/-2_]RTYN:,d3?^FCdP.F;SZZ8Q>T
Vd[?E]HcM>)[HKNXEK+fE;7=8@Cced1cP;^BP_Wg):;(Rf1:2)H7=LG]RYJ_d,]_
_d0a6/FfB[HD<RP-AOL]\cZaITaM@&](NU+CK,\:4]6HHeF0dM3RDH\,@D:d3Y69
?0+(;gE4)AAXKKd2WYd@?Q;=Vf_O92GE03WO=E=W,\@^X9EC?f]FQ8PP@#91Q+cd
;Q,F6;RFSXU<Y.1FY.3M.ga=F?3@?-<M.JX2SA3BPSVCIgR^_CZc4ZSc.W/&(^26
:(?EXC-7#BX8=dU(IK&0:?UNOC&W94^6G_=+N6_]c8[K#=ZePa:>P\-?b]\GQX\@
;3Qe:9bTLUCOg<,KQN7_5NDQdIB\.e-GQ0>O\Y#OS?-NDgMQG4Q_c,>=):ZVNL\8
g.a53:6[?S.dbIC+(edT(Q,1?2Rc:G=),V5fefTc&UJMF.D6aff\1;H-PSVJW?56
9]S8<f,HGMRg7<VJD71&V3e)g:R@d^^9Q5MZE##6_F5V.-ET4+LQ=TdDTQKWKNa-
R9aLV=-9<,Q<d-RCLfWC2G[/@NI+c5Y;@B2SIL7AO-OIE5[K0OgFHN8KMD#LQfTf
MDeW2Gc8B3(>-LAV&XFH6LB^U7<1S@2c1_9G-RHg?VTMVX:f129U\ggg68>[S+:Y
<^)]<@D1.a,G#@\D=]0-gBe8;;=\^La8;NIKfaCQ=1];F6],FHMP_;22<L2)HBKL
4I:?X2\V7;>1QKH]KM9g6Ve;=I@/egUd=9UCa;0K13>3&KE5MWVBH1T9-^K@&<EJ
_P0Z#Ea#M\f:IQZNBFYME(aLD#bGafQFOXBQc9+D4A.QE?AK[;,U--2\F&CDc?\b
K2(/]c]W\.B+1X32O.aG2\QUNZO9T;=g.<W>=B-A#;<&AL^5SB4bV(;e8cd(AVC#
b>IZ^@\]bg^MGVORYaG.;;g&]1?fB1DAAIUg0d,S#WIUBJKQO(::/R]Eb-OH8a@.
;<dI\WT3)00##=DbGZ#:1e60L5VdV4B;)1[Ob8XUA/G55@DYYVRA>O6;TcUS/7SK
9?5Y:AY+-6_gN#GY<V9),;5DK(=<>Lg/14=Q/,1d+M@P_/U<BFMJ:#X@NE[WH(,G
IB-J.<Ia+aO@aO)5?YEQ5SH[:&/T6b/0G#bfSQbH3L:REX;ORF-BP5_UcF_;0S<>
M/>EAU&08O,KVc\1Ue>&&eDcJZVeeQ(IH4#].4=#0B8.DbQe\H>F\,g7-M#>KB]/
5JGdfcJ>7WD/WD[B;_\&1W(_LbI_YHR;UefJ+X735Y.XZMFMBa0+Waf/GdFcP5:S
9K#e1P#,8Y>JJA:S\[YO,XCgUW,<3Me6IOIF1_S76U)PNZMB@6-F7KE@e17V;^<Q
U<)7a+6(L4&c?^=(X@Jc]T><T7aWIT&f7d(f,HZL>,cQa0]SSf<NGZ&A/:,.#S2)
E35fgTB?_b71DK_^ZT#;]H9O1]=58;TLcd1WV[NQ:),c(:)NT2,P:_a1LMH<AV7g
QBEgf)6Y(8UG0QOQ29Kb+aVT=bUeF[Vf:2G6K(>gX?Ng(eD=2c-:BLC.6=HVG8+g
#e\(S;C,5Xe1W\:<(?9OR&E&Q0a2+MV^@<=4MKS,0b:=a^];G_NSe,M-80+(G7(6
4Pa^[HU_^6?K2GfR&:Rc0QMK@VHT/:b&KL.CO(5G=CfObR5@^AQW]b2(GIaWFQX.
;B?Pbc79JDCO@Y)b7W)N(TX3O,^8_)X#G+YT.:(b.6>CWT-_66-DT27gPTZc?e_a
\C+bKVd0;2W9=CKYOV1=aHR22c?QRTDC^8b2.dXIAXg\D-.+Q^Z\d5EBTdRB3F>;
0IWJbe2PF.VEPM5cBIO_\_0WB_;F0#(AUE_H_MU#>X]+SWH?CLB7?6#+<K22Z@=P
;9;5NY3&74O,.2JP<7=)?>e7++1=I2.e&b[D538U0<JW&/eIC@A/a?WE.).TU<VN
a8RPBCAIOFMHa:V-X7)S<0RS_>/EeT#PbU87R4+(127/QU6_)5P:+\-D>YUIV7Ef
ID5524@9J0VKM=ZS7[;Xeg@-Pa?K)4_2aUL=e67d;g/4I@Fe<]^77#,A:?C?S#NK
[4]@/6fL2;+>a(+]0?Eb)O@@X<76O5MEdHK;PT\J0W2MA>YaOO?YGB>=VL0dPU6M
.2B1Z3),#E2c/C:Q;33]@9EffN-(5O:L<Ka:;8S,._T7-Z&>9H.)b-4H=dAgTR1W
.2^X-P4#1/&8d)g_+EC9@4-SM4B&KVC(:(gXX8=T\5WM7,Ua)f;>[bN[KCW/:dO<
bc0.YL1)^b-#SHQ:A[Ae[/)Hdg6O/+34[-\RWM=_CZH+g#9_)[FSaCV5Ka.I7SK-
gNZ7^[1^2RGBdC8-7K]4+FSef()e^P8/O?f(XdU]43BF?Wd#@W8@d-#,=,@9:Ge2
V(M^034I7HcO-JKC@Z5aV8.-eQf)S@O@.dOJ0@P[8egK5[7dQ)[CD.[@,BPUX??X
W@f^d..;Y+C>Aa1/I<>W.\B8S7d]5^&/ec(<33J-fA[AbB6RAF#6#QZf(cJEK?V_
PMH=N<1]7_c?cgFQ7YK8KY]b5,?LR5DCT8-MIGQ9Nc/CKbFGR\FG\Yg0(?9>d]NZ
INdV=Q[3ER\<Y\<4^_A#&RQ/\\IWc>H@]J2<gcfE4MKGW,VCO3VK,RdY96B/HF-N
K+;cN>67JHeDe2;gN7;f?PI3;Sa+QJDXR+WVW0JaF=96&DUe@:gB-&A/NWPWOH0[
I83NJd^MW7PY;;@2OWN9KBJH&S0;4]_C7P6V&XZPJJ=g\K19WbY<O+?VZ3W.f,eQ
]Cg]U(e8be(ZM9XdXH/LBd+]3e5-BF80Xb2aYKc0W=W\aW/)-.[T?+De,LXb<>Qc
Y6AV=BAf;V,Z>gV/:X./+6D^:f?DX[PcgNO4=?\c?Y\T0TL:FdYPXc;H:_3E,Q/:
DY3_.J^Bc6[#Z/_/N0aQ_:f14G-Vb@QX5HZDLJ9AL=9+GW<]aWAKZK,^>:\HFIY[
6.IWH35CJI=\W/I)f4B<-W-VGG34e,d6S)<_Z6]O2/C2P>&dVd:?QRQ@)V,LAdK)
RfIM5-]NYIcePG_a21--dgE?CIGgM?0V=f3SdN@(TaN^c&;c.U#ILIe2b<c3P=?f
5MVF/ZRL:]&C)AWD=,[d>H?>eg45M2JH-Bf.M0/4N,-74RWUJGGIWLY44M49E]:A
6XI9b.R\6aS4_,BNI&bf0UQ5CY1cF_0CWTPY_K\-\PYU[LI@,.1X_UE2JTN\E.Re
gVSC^BFPN_C<]-CGBQ-\4N7],EEGFC=->]eV4+>1Fb3V[WZdI=:)d1c8TZ-.YfK9
_JM@K2[J^L-)1@L_4V,?edNYMa.N0PU1EeT097DQLB?53+5Hg4^?BKS1a(JZ6)e#
L;ZN#HWE3JBGAfN=@:Q1ISR<AEHDO0AcQ8)\;=aT)d-#1BL&aG^B[.,)C&gJJS&F
2#6bKSeRA,9,2\;f[E>GS(OBDJcWMeS@9;YMF9</_FO-#a=-c1+;SBK>(0Z:4VYE
Se6?KN^I&RGN\@QPIAa:FVCY4=3b[c^AA1fWWQ6OD:;T\gbgDGLEaLBFIONU3[6K
c#&Maf2B2])A:IYg,HaI<aYe]LED:JMI//eVE-Ge=(@+Ia1)9#3&XA0aWRMJAC=#
X8)HRC=PfDD.P=P(\Z;7d]eDZ^>bR<KUb2P:@Z(d,=,&G;-J&VAZ2>2V[6_,RF--
807F(d_0MS63QHa(9)_Mc^EVXKC)W\.JVTWaA1GW]AR4P[dT.=NT7.eN5#T#/Y3?
YEI[N@[f5Oe66Wb1=,JDV6g-3bd2F/D__I/U:CF21/\^7V/Z.]V6:9:SH(#&@Of#
L+a1&RJ_UB?:Z1/7VVf8+>K>\-..9f.7>4d)?T#1\\eEWP>BOU722+F.bG_H5OLC
g@:&@@L,YAQL)7,d6[SPK5CT@F9@8;3XM+O,@NYaaPZ::T]Scd,3XE6XbVe[T0OQ
B^)(C&U2X8Q\U08]fNI8>WCe6HDV/Q:#V.<6<eTgM^O7]2EbI0]8+<Z[,CBR[XLX
DW;M(.D4RVE)b]0fBRX2K[O8_8=a\T6[)(7:]DP66>D@K9FDO_e^B^_ZJ7,+FK/6
MRIC\Z]g,@S=]V^7WTC+T[(KR/.AXf+#>Y1dOOA_[O8[c(17TAD)6=;CRBgK#A(J
>6DYUBLH<DAK[2TMW<_<P+T]Z?aA->/;;VY6G4P1J.&)UE20?4]GY-R\P7TOC6bI
H/09H2bCVV:_d<X/P[;23LQgVCRJ^^B6P?F)L@)HXCBH\DC>S9XAB92\FGR,K5LL
E8E?B<19\\-H:LBd4-,NS/FaZ]3[_S-TXTY6-OWeZ1NMO:?I[@ZZ;5O3/UR2.YPP
bVLC\KfO-Cf_aX<RcIGB>VYVa<g7<f=1K/UAD+/:SOI=SV:aE+?K7,dRdHHd#\U3
@YG]S#:\b=J_/=7X5B+Vf<D.4#:G33#MRS_)L-g<HWH6cTGM/996F<?R[A5\fPU5
[3cCP]&7\W[OX^163-E1D2PE9YNTNUb(UM?\g7NN3X^;GF0YY>RY^MPT)bAP:b1(
BLCbg#732KVNdeCGVRb5(d[N@(:V2U7S>gTaBT#\M(EY.J45YB:3eR&XbbP5QOW,
TNI2;/.6-^YJ15LZINZ1OK98IY/10W;c3D_;QZL<^IB#&Ga-0FL[_K0/./BV:+K5
SdKY:&efH#^QC+0b:4EcN^D4N)<X27=?d\T4?^2/d,gb;NA@Y_BQ(@.2eWQWB:c=
6>0/TE?S]WFY.E&W7:-&7;9&,K_T[;=UKYaW9-:DdUXVKgfAX.8:<P=IRJHNU9?(
7c0ST:R>L,^U^^E=,aD^/9bKAd+LX^(+2NLg9B,7G@5?B0U[[+(-PK<BVO9C#PWg
U81#)&XD,^5L:0RVIc=P=a=#2gMUM=0<8K4Mf<\\^+D[.,IJVWOPY>8P>DOgVZc6
GQR;\Q@2L<F:.A/C5^a[:GCWH:257PJ-J2cgK_Z:L:]1eOT9bMB5IEQ0AKV:eYZd
:)g;34PA&a)b\e(AdV7-CPII1K))cTQWcCCe=\1[;[D?=F@4-C@UYIOIHEAQ-dKW
5IPN3H,C-E/S3Vb6,UYF@[YbSEO=1H@fe@<QC[?SA8T,3MYeR16E647FIT2?Z0:W
D[/U]2)#Cbd1QJ_F(Y@NA5b7fJEfQ0ZX1)2fKE_b:WZR1^=27A.Y,6(HY^Te#Q#G
QR/UMOORSQDaW/DOA6f5QQU]30\GJ#C(:0=JTX5G_E7ZJI_3c_YI8#,&VLA1d@/4
>Z^4L69M60(<HT_[;dP5-gBONNK6.Q(fX13=IB]T?UO._(SR-aT+.bA5R1G:cae<
>94?43D>T^\.GE()C=]50(:=7^4a,c>QJFbK-HC@XMH#_P32(6VQWX2M2.?Y976/
Ve15UQ0GL-+GY[>QBH/M^?2OZGL?5&J9U5dJS?BIC:^a8:CN1U^RT+R89aCc-3:D
R?YQT,?(9f3RNO#5aP0>YM8/2;gJPL1R=L2d3CM5/<0_BI(GK5.^QAKJ8TQ(aS1@
QD6b2&IJDTYI^.I9B5[P]4[g22.T\_8:>T=A_JNb4Pf?:I<8c+0/NW]=.[VM#dBA
1bTT.]_=;OWB2Y,X8gH@We7eQ@O5]dEN,^\PdX[B9gL[=Rd+_,(.EZ2_O8,0-d^=
.DU963V?DBR:N<#UaM-OE.MbAR:^X^?G30)aN.LNKV#X=O+R1A\;#BMA_Y\(F72,
e=0;4:E.ES?.P=Q.c<6JH19K/6B6/3.?O=S@[3=/0(c-B^_U:K+05d[SeEVJ2.f3
a_P=8_I?N4M\2,WYG8NXc,Jg<g7PBa)eI@QK&)SdJc#+\2P8,4Kg6_R=-T&;=:?R
Cg/+T??c86RK;WT,&G-;;RZR2e5aU#>K=H^Q3UJX[MJ8-,1-+I0E4@d>:V_Z;0a0
D+QDD?UUG.eBYVRZ31]ZKW;+1dIFXc,8AL(8=L:]]CC?(9[cK\bc+<:d<]FX:JB?
FO>E1@=2TFL1-?=K&CA?_3JA8N:BXM=Y34L[da&f.VDQ9@<=+3OT7b9TG@B;:^Y7
#fc67;MWS3[eP1N,e5_T_@KT6W99P)Y&<_&0GY?;99+WH\gKeL/GQ:Z_0gcG(@Fa
7;IFfVK@1V^f6_\5\56YYPZ2L&e^;48](A22/c6Xb+]/Ea+G6U=RE++M)+N1SVJS
VeKB<6gZ0C<5cWC/:UZ48;(O9/9Y:KPK387?^M2&e[2HT9@1aQA0R;SZLYeG+SR)
?H#QIWB.A:De=Bd=0<SIWAB>aa[Je4O\b4fb3+NLUQfP/QYQOOd7FYSG_D<SDee;
8Ia1HQ8QR&;4gg?HP5>](?M8?4eaZ=J;-;Jab+5,^17+)3?cfP9:c>E))6Jff_-5
R^bd9.4-#7\eVZ]@S=9Y@VaJbSCU3-c7GBXK8B=gXY)B79^)/)76g-ag&F^R8[4-
K>Y=P6<d=Fe^&JT[\cDf\BGW9]/TQMS4aAC?\YDdBQ?FWOJZAPOVV8_N:=L<SL(K
fOS>-IU9B)M402TZU+_-P.V3e&:c/UL,Z9VM&e#[CPcO797I#7^O6,?Eced\.6.9
DN+BD>K3=7aHDA\M]].M[g=TG2HF_;RV>CDC6.7G^,YTMT]S5#IXa.)H-ZQ>b:eE
8[7fUgYdJKEMC\]7AYAOf-E#_28JQK0M&O3[?bPY4F+?-:-I<3X8^W]SdZ:;4<TY
LY,eT1V:V?GO5@SXN8A3_C&(5V@Z2GGWe?EOK9<K;>-55HObS;5KcYP3UNF6O;8H
2<\S=\Z+Ya1b\?+0M(ZKUU9g.OFL[CHS:fNB7.93AR],,2TGb?T.XaEW-<1]RLVb
)a]Ed:T.WeE=Za#JI\[E(0/CgfV&&O#5?.#?]_e9>X\WKE?-W]U3+CfCc;32,f/N
-P]823O_<E.G^=4#-2U8VOFMO6V3d[L,FW>gDXZM>eZcP]PS8VM0?Ce2_K8eTJK@
#]E-:e)dPcYC61JGIBF\ZR60Q?DOH+gM#eaI&(D01EaM67:eJ_R=H+W@W3dFUW(F
[_PC0Q/;g#PCFbggV+dRKU#,-UIOa5gJ[e_e)G#Ug?aCGH4->N<<=a\eN@.[E?gO
F8(B<LPP=@8R9ReOO65]E6EX6HY[VL)acH)DQLKTKgg/<CJPDX>Pg/8<N8IQ#TGO
RAdQH&))#Y.&D8#dZK,8AORV\SC;_^Sc>7IZF@UcMQIdT.9e2ND6#.&BS?_S9FWR
d?cTU(#:\U88^1AV<E/?7=OgbeA73?Q,H+0WK1_PG,3U_8Q_[^K4=_UZHUSV7@?d
81\gH6MC14\]W@@L@/=EIB[XDDUXd4+UH+5]=M7-X]C.?O_?=ILDa+>@ML(]]O[H
XQO2.UK;=F]?TB6MCQd&3@Mf[TDDU))XTO\<P3@(/O/L<6F_,]>R+Sf&Ae:DAXfF
LOaJF@ZZacK+X:(8P1F2&T?..SFE>V(DL?8^HDW57OQ.3.(>P=N]GCONbJQ2YX<N
EaCe3VFGA@8ED+Q7N#?/LaK;AUd<?Zgg]B=,[5WA-A7A&])#\cK1Ff-(>Y-QHe^\
.>eIIFa87cR7)ODaUIE^DI[M>ZH)QTN,W6.IgC3Y8^29N09fee-YDUT7ZaSWA2+f
^?#P_+><Qab,8S8<J=D3\Y=;AR7Nf^^@&aeNT30Kfab[De3#@+.AA28_R-L=TD3]
QMR:7X#cUZ1FSIJ&B?<H;e#,K6XaVLR>\IPPgY^C@@JN#ER0a70Ra#4e1HIC<IUA
HDW+Xd3^CS.[MBR@S]SFU@/7@Dg@\2)MQeBfdG#3YGA3AOXU-YgAY)4]fHQ]cT7,
V5G>YG((5GcUTT>(8]N4<NDV=GaD&6Z2CIc\Ra\0da@V=HQN(VUGKU5\S6Q/_+/?
2Ge#50RPVHb=Q=M/(VVX_\3<R=g<_+4[;GaG64/&SG^&cKG,I9H-L8WO\)D8)L^\
gWG2)SIeEF94;CY8a,Pf4(:da2V-4(O#CXeMT(T<]-=(JQIa=2-3f9C1?e<Y^?Fc
8F;Y[&X]998UU;cHC5-dJ+F8#E_>8e2U3b(YI:L)KXGGXeI9_Z5PYA_TZD-.4N_\
gR#NG?dQ9e\UAXaW,PRA8eGdH[9>.A#<,WK1#6I-I7YfNX](L:4GX0fW5JW<+OaJ
3Ce[Z#34A7+;M0HM_RX@Y6cR<7,Yea1M&EO__U30^=6,(2>+fM:9[S;]N,=D)DH#
/@V8J;<85X\J2=QBP1FQd?/M-P6O7NGb-.ce-=R8?<#ITSNJa1C8Oc52-5C4.1TT
]+EZ80ZTgI0>GM]2>4(B,-bFfWPDW#+cLI4Q5]>28<DK@dS11><[-#&<UZ^U8+OQ
G9YL-&M7M4gOV;+a4K&7@fDgZS.=L;+L,7F7DbOIbeDISa#[8[F0OFGdMP7A.8M3
EUNT;[HBdC[WJY<JGcZ7@[@3MUR_2[EaAU@8RLFgLK&+[;&^a,[\H>-8M&9+_[J]
QLZ:Eb(.Bd&0QCdUFQe@P4=f+Ac]Q6-4WM7W2,b(SaRN,.-S-EQbfQP4X@F6c518
PXIK\eHH\,L8L>3JgVI9bLN_(?+f2[UWF1#\4C)A@SH:46f8bgI;VC1@#D30&:YE
WWK2^(8ccdZE#)AK/.5EWW,?/G4#I-&=aDUI8&JcF)g>M<YERU?X7+IbR?QH_Q3c
DbH+/^g@^G9/Z;C=eOW>+IPPNTSG>aNMG9M-/DI]9&J,6389bPDB[Ud<ZH;AKeG9
ELW&9.#K0C>CIA))EdL1XSg99W6bI&e_N3FL,RSd1XMW?T4AZd,)\3K/V@c6)JC>
=c5KEQ,)gUJ9)#BE57##IFVC,YL0>Cd0Y>,9+AN1P;^:UUPD(P[RW?HAS63dJXGC
BTFU?W+XXg@G1<:Qb;&:X1V<:_0.LXd&+W[7\?+Y0,,eWGbfPPDQ&2Jb4F-6d.;f
;MLR]95U0M;g.Y1a9/BTO-Wc]UdfFLP<97[B=e^GIT7H0B,:D&2e2A35T@?LL+Tb
gQ4>8Q2&BF7PGROLJ]H&X6N9VJa1?#Q&d&5U8]d9^09B0>PK6,S-NG2-OYDMc8MS
VIDMPKAG3&Ve,@.X@?1VbE4D)DIM]YE/4,:2HL+f0M=U36Kd.>JT^W:1YH8&,K+X
RWQeR)7=J.E(gB,L.gY_9AG10-;fcFW>bEE=L+7/U0SLa8YJO#Z2PQHG6dLB4^C[
X3[1(RE<-5#++8:U2T12+/M^5]].&(VfYDd6aJI3OIZ<e>3FePE_08&+(==]6W_>
.=0,Vcc1075Y^Db[Z,95Wf]f7D[56);Z=D)e4b0;J:H#;eT1Va6A3KT/@URYNP.O
-[(^)M,D0LePM>/?OO@]e(EUZ4P5J7;(J_A9a@JAdKA1FGZ>fDFIOP3fDG+EAQ<Q
SAB_C/a;@F[Y9W/)&6+RDF]D2McW@Aa^b]>;&7g^?B<H,4e&0BYADa6a<\3Z^2D3
^:RO=.&+9FbVd4NBc0<T[gYJA:@/Cf=L,->:AN@@0@0,\(gNRXN^N1.14c:g.U,T
:[:e<)43JD-b7-aa]OQ/ZRCgW9\\CC:Z,)#7_\Dad3A]2F3XNU]9;[69<4@(5@NE
8faQ^YKeY<RNcg.>cLOD-Y/NQgXGLUICC/02<8(N0\HA-W0ROR7Cf=(SG1]6[G;,
DM1&1ZGI.BMSF2&@1U]aOCEUJg)9B_^:W?>#U:?aTE,[Tc-O3XA@Of3;6D5^JRc^
B6LE=SJEBadOKd<Yaee;E/#E<0(JBeP?#]EZW\SfgDR1VZDK-c2Ceca32(,:fbac
gJ29621\?H7f&K>]R/28a#+GO(]3[6CUfIRHTC2NOTOL5;fL5VB>IPEeG/8YcG,[
;/8?M-ECb;JYJT=9N-3_FdaAK=M.--R;2cd(S;@X(B[:YQV(b@^f6_dU^#U7J\de
Gg(aL+,S&UQS,U5,@K1QAKT/8<61(J@A12VeR2Zda#,eaY\DE,S4JNX;,?E.4_\U
;>TX4GaXJHbg1Fd?DA&e;X^AJFXB@B/L-9V04egLLIKY8/-VG35Ea6TPa&JK>B;/
eec]XHgKSQ60AgMg.=E/KRTHg>OM2:P6.^#YW_7cZeF;I\#MC9X6H84=IQMR7gSg
\[S.>@YcaJY/D+TI08g9RX:^/7R,gf>6O_BH>CK,KG-47=C)5S.T.X5Y&F=9FAV_
#?e7gHbXJ9E3?BTg(:A:&eT)KIK-cZ?\P>2Mc<D>]-cJ#DEZE4cHSB/?b9e.cEP(
66c8HZ^7b214GcBYP9Y17#.XKEd4cV_TM#VLP/^RQUK9QQ118:YZOS?)#PH9GKD3
)aI=Q^618WGO8=KcWXZ+<6BX_(4-ODY^7VRVET-^44ag1L.9XHY5/3?NW\T=/C3)
&)SU<CX?[T)8LT<39AB8BIcO3(DaQ/=#_N+KGgfJW[R].^&b1<274DfPAgP4gE@2
fPQI:)cbE+c_JPcdY&:a#,ZWOUP-Z\Z[M^]e0bUM7^Ne)H,g=:H7D;VUN=7fPdC.
B.1;e8^JAHG2P(P:,e8;f[8<5U5+Q^#XMcK))T)+XVW1;J_TDAW:d5+BYZ)&)O.J
7@b8@;-HVc),]GbgPT4]=6G<U;755J2U0KW7NRR=RICIK(0@I;YdeBR<<:_YUe;1
<M)S,.O68?d+,<9#Y9e[H<d,I3W[&=0D?A,;G)UQEQP/\,,O[OG3e9Z1:,K-dSR#
70^[a.QL6GQ,2DYI]bA[Xd)GEYH:?5V&YY(DSPe@JMe4<C,^IS5f59;KI@-.IRc]
10@b6bG4B#Q+#VUMEEDXQ;eIA;R8-OX<F7gDM:R4]bNGQ#MJf7ZGK-NNLf7AS;C\
=C^B3O-7ZU^X9((=2LgC^b#5fCWZ)A#Rc>NC/\7ZVJ5J.]caH,+4B#Sb.;JUa/TX
S8?O+?E;+NDRB_RI\B(.7CYBT,H3#@YM>3d\,gT.R.VdUCYB>)Tg6PU4T=eGK^21
9@#F2IH8H3\E7Z5=C/6g-_=7ML?fI__O6/.Y/PE+/K5=Yea^5,2@4_c2c>CVAI^:
)50&]@#P>6[YSJ,]#<A89eSJEgV;?=TMK5>fSL#^84de9JG&(e]H?c_P;(9c9_Ab
:7?2?;d^@a6.-Tb53)K(L+F89[/^C76bTF)WQfX]KW#BK]21.J/[d::Z=>UX^<^D
(/2FH6f2YU778W4R;/14fKHGX,VG6L2G>=/PS/5g;0ePD#EB/[\..ZUI.]0@),Z7
V2KQaLfe&dEg7AV/-AN16D--)c(b-Q#7S[80137<,;50V41OT1BTRU<_8N.5Ua9N
F<:EbWc<1_+ZAc?,^;N+HaR84:<5Df09QE+D=_Rb/<eHDU6SZD#Y4cY(44&1?-U8
D]ZbUCK9#bIY6S\Fd:G+\2+E9\_]Vac@6@AS)FZ<)@cFDJ\Na7E,UL>>dTM7d:Y^
J/&#I_BZFFL8D]dI?OcfYXSf^?bFC5SW]:A\c>T_bPReM9GK>XV+.4EbR54;W(+T
0[1+eK_?5U;V_MfMde.\(?VS6.MWNcM)6J]KYaCR^V;ZVA+b#4Mef>.TTT^&2Hb8
XJ2X@Z.0;T+E(Q4Q2,\^-\]1NLQ9:COQ==SONe;VF#.Ga#Jc.:2&.@^(PaK\M1?8
(CKEgVg@IRV+8aW],+=e]=S>8,KXXFR<E)#0N]1-T([)_K7TSgDaG)6R.4+2GAda
P[Ic,16XdM&NC(eRQ(D5cCJ#MG9BVOJ:B<fM>/bHTD)#e>HHCIJW_cL,553UCF6S
ZQ5<X@Qee\9<3?;NF)7=A?^YG6+D#ebEGV2gPHS4(YMH_61](1CCGJB,9NR2/9?-
JNfD:?0>#ebgPaI(ed>B7]\0H9NVgE\JC):YN?ePe]dA?N:DH>CR>aEd[b;g0^OI
QKOf1H7?.H&Ie6c9E\eVCAP5A=\f^,8YN(^Jb8KV>aLO8^L5Tb]727E[,^_3+N?X
8CBSDYR[3-[04<EB;R2=UJ,;+d-P\[a[Y<BJ#:BC[C]/_03&8T0-]C.D>2N>SVV]
5JT62?a/[g#//D?C1&YG_WR[Re:J_Y<fEa,I.L6)PQEe&c#XWO6[:BIZdLTVdSSd
2<V+_JQD_]A/WI812V&0,9K+8]/,,EJ&YJ_/bOL,F087I?;T<HD6/34E4E.V]bf[
RbG9[EAYYa7Q-D]YT-QcW8;U=W\UTMNc>M1M7gbcQ^dcTT5VFIJ0Cf-eBSgARF,S
2IU0/]GANf1aZ48a8^.WM&/.4cM=[^PQ&]</=I_N8696UHb9E+RWMO?_bCH(E]Sc
>VaPN(7-T^G3/<OR[8VN^D8ADB?MZS7g(@IE@_PY4NCO&&6F;:PRBd@:5UEd:bK:
AN/;@)-;>G.\[8[0SeRZ&905_J#W/Q<LR)\gPLRM/UGF<eDf)SO)D3QF+QK&WAKU
3dKI&AX=3CU3bYSg8GP2_gB;>#8_e=5F:cK#1P5.IL4Y.#,#M9BE]3IY>3a/N]-Q
(4bGJb;5DNI&/18(X_^J[&A)YD+g#UgfcVWZ_@Y<46:37X8>IU0AS/bOI=XZ-EK5
(dR:DE(-Ed^/^ZS4TVQ(D/]S7^IX/]4AOFMK^EDNN(?L-CC(5JF;[b567DA#=HfC
#R+Z11\2<^9;=.JDAD2GB[L&)\]7?O=\YR-e9@Pc#.-6T/EAJ/6(.C=FAdY<;Z+N
c9B9XcARG05W:^YOP=5,S#MDAB3QG<0>?2YOXPDF=_H)K8bE@fQ042e<J,)P8g[#
d)RF,;A@MAgKcI,6#\aPa90?R26EYV:/<bO2T.V/PZRN&S?d2KeZB0c2PYLP]LO+
:[U>?d>e..cTAcQ9E.KIFTQ_L2J4\6V?U/F2F?;BO>AN9B2-WX@KI=Ua-;&\9./V
cE=Ug=6@g-))+>LGK26JF?09JCV#G,6D=a]_/-cJG#91WI7d,1(eH&6CP4]^[Q;.
ET9]K<L3RXY19\H/_2E9-V7H+FBMY(([,T_P9eIJ6f:QMN1ZT[?W;Hb/K.KI03FQ
)2E(>WT5S:8.=Z]N_f94XT+ALG[?5(5ZX]@<O+MCH_H4-][gORM>b9#55;OeSf3(
CLdX(F)5N:YC-SW<[KGR4:FFKRSd-_IWRfCW9-130O-H+gcJ_T,Z?DLa2Bb)_#eL
e.D>YS<+)8U1/Baf#DUT#S:V+PLP4>NVF:DQZ=-?R(e4^TXI[O[OLHI?8Z9]A_[#
\bK@6E;R7U9-G[J/fd7OAL?.R<USC3O79B72.E3N4\6Y3GRC.<fL4e(>bf]U[U;L
L[KQK[?GXgK+[70#3IQJ,e4<QA(PLP<>.-4B41KBZ)^g8@5bO/4A3c&XYPEF-^V9
NSJDVc/PV2P2N/KJ83^J2#gF64#5W=;>FPdH3-+K]-PYfY./]7AL.AR,MK/^Sf+I
:SE+.UGf_D\4;D;ZBa.AV,:9@R@8F8:;7FR9>^Xg#N_V0DGWOIg.-5Y+\8+\:@//
\(74+20@C\6;RgWab=&S27dF)69I;I4+a4:;_g5_#QP]8B.V^G=[fZ^LEHSYOe.\
:W/V.RZSGP;b=3b6PZ2UDB2PS8BUbRIR=3Ug\POR?OG>SNJAR.LB3[4b]bMR\GC3
48eR[KF9fe]e/MZJ)_gXeWL[UR/]-]Ngd=H>=45VQK5_,Gd;:G63_dF?QC0.YZ?]
U:;ZI>.Oa1_2BXJL79Gg0TT(CA5<5C;5=.B7XG2IJ8OER9?]ZEF1HIFO0-ZeCHD1
6-d2/07Ng+/-R<S,T5UdSA/DfW^,]RUKIIJ6&Ma@g6BY8Z)C]M-.6NA;;:S:]Ga]
WOf01<,8)X[JCZG1g7\;&:.KGI2T[7>c5LWH94SLRbfT=;JEBa<>)S2aBIg<#H1;
-R/LaQMf4[4K\ccF9Q3@XZN6B[8BK:FGQbdR=cdSKGDd_I3b;df)88d+_,<@15+9
Y]E6JgD19UB#&e&XT0Q]fF<1MI.?4bMK[G:8<64W9;_,M)-O9=[B.?cR:TLLV&C>
?FF_8d6baY_OJ?54CHA<<^3(>f)Nc(CR0\[1J<,@aMVP.e/dS=1M@U:Xf9WR\[AP
2UV;?]gXUZEL/c>4c7P31N7[SSZN<JI5Ke1a_C#H5@U:)A3I&AGQP5Q2)WHf_4^E
fb\?#XC87^+K&JU#1?E()c<B(3/MM#6:0AV0/2=<HKFJVA1?TK@aZ)]0K3YCS)JW
FMM<b;-Nf9-P#<.5>.cH)L_G?LVcE+,3U0\U<?eNKUe//TMTD.I8Ice:(6Q41E2G
+XP5S60adCQ^d(9a/8Mge)5KFeg<&0Y8#FVfOU,QB8J7_bM8TQ=AAcR@ORAV;4.[
b+c9C:[;[Ce\_;4UW<_97\ODfVF76dZG]KKJ63RP?V8@STS16<MdPN_(JSEG?GWb
K13dDWF2GDgLD(CI_4&<D=3SNS#Fd^A=L0AUDO&c4EN/^4e1D]]O-U1#AKGdM[e3
ZPYO00\9[P(54?WY,WaCF&RG(RPEAL+QK^\?]6^E9O[JFN#1ce9GJ=-1]->,5aLA
?EH)f\DV]&<5g><4+QY3ALI@T8G?T-:Sb<6WXI4WV:R^Na]CO1-^(9aE1IH-)OI\
7<^_eB(>Tf,-7UYYVb]6[7_^(C>S)f2ST.K/E2Y8G62gNdS):^NL=d3,M1NUdK5#
G1SOTWI,0&(E;WHacSRH]O1:QT=\PWVLJge\(BHBO3,97X8OB[J7AGH2E#P&1W#8
&f[ZX@\=9Lg07&=FHEeKM([V4^P2T^#9AcM?gPC=H961cVa@]O:c5[Q#/6F?9Id_
>4L#=5L-@.@#<fFJ.cU5a6:Q:[[E82)(>S;=LM&1ge[BF27FL?QY9I_8LJV=PUeA
XT6_c5.MV3S&&EP_=DLNT]I)eT::NV4Y,SXb<XHY?^cK[ab+>cFAN2b(U@-)(XW3
dZ6(2&DY(\?J1J?PBJ9/>.,C)V0,6\e_&#5J:#BHG5c2T\2UQ^,0:PX8/3&G0MF_
aNT@<f/DZaBPVS,SJfLYP0W,1:aDS;;ST2,_7U74ICMX@?ZP,1QEGOR>@3DF3FSX
59d82]QG]@B523>Y43.(?-;Re,Fd-Q#DFUP7D+PFNde<_f97@Cd8gff_[ag,:(a]
-8,8T/fgP\\K;I=JWVWgbJIJ+=E^XT+>0=?:++.E(A@/;[K61NI3d_M:Qb]fYU.R
B\G/>@@GO^(NY5(ES7,L&1W;X)F9-&TI_U<S2U@M28>_dc4PDP?DYNaIV-RdU6UM
]&#-f3b++1>Z_G:<6;c+11+R8eS\7MM@3&U:fCI+#Af0)]c5V.C\C(f=AU&gUfE&
N;>QU=IWe-5NNX0&1<@aV&?IbR-)YK-fIS7#VdX>6a6_8fACENZ7GQ^.G7OdX[)f
T_A>:TL>f.WW_1D?1\ab1EL2#Z7:2)81C8F_(Ae\aSc5aNMb#49V&Z@=G00ZW[_d
d\>P#-;O,49Z78Z(<Oe]+e\)V;HEL#XFBBG/H#FLZ]KZG@c7X^<RaNW^P0+8N[BR
BQ(Sag3NKU>GTWC3[04JE+O5YeFA1JKZW+[P-7P42;OY2L+_ZI>WdJW5N5S4Xe@g
E/VPDbH;bN2032P-8N3Z@WJeU1J.6+57.U\,GUeXBE075b0_\4G+7fK<)J,eMd2Z
E&f@]344E11_+TZJRV?f)G#RKg:+UUN@A8???@Z?J]/fA14#:d]J<c8[^,a^dVf:
@P/Xa14^BW,>+??O5((M;QO041+L9K,R9d:7e0K6d[:Q]#2a1<QF>+4I3C@UJUQ-
bK#6HEY:+B1P?_^N;60=FL,SWRO^\@,,.D7^^2ReS,-EgEYZME;9DEL@9HE4=G;c
NE^;SRQPXHGgF=K>KS+<gOXXGIC8N]d3=b[[f//-\E>a/)g#[\JYTJE;F^;ed_/2
adA;6GJSKO+8gMfF\;Z8(?<a=4YdR(L-P.-M&Ea9c=5R]b_>E)?PceOVZN>Tc//-
X>C/(2=\AXSbHY<C.g/+e(?a3f.S+L6>MBKM-D^G7F]QAbI(/2d,@]K>fGYgQ&\7
EcE);G?@d1)Zb/<d)EVPVeWXJ[3&-)Za#6-(E&bCJ22:V.NPP<<Y.1PJJ<L_I:8)
J3b\HB)Z^a.5+>fMcOV&?^?Y=e)6fg/TZWZdW0e2LA\MDW-2OJ58BfBNJF:>78?^
)=MTR^N7SI2PHPA?7dFGD_CXW]?8-M[e=B+I^9G+&V:HdF);^_\)=e=RGT1<)&^J
60JXdfPZIE4Z;\9Cg48cYJ920JT9[dYP_\/0c)4Y7]NWDD@ZS.Bd24V8B1NR(446
1AB..L]YRL&-W736;ZZ+fSXa5@[^(g5g-b0+]:1UaH6:;eYW314Z^dC#NWGeJWF:
6HUTZeA/CM?WEFVec?,IdE>I[31/=:^NF)1Jg&=/Of=U09N[O_+5ZeV9LS=J]@IW
;5f\TZO)LLHB2f/:/1Mb[)?2ZCH-5OF+UeX_LZegYXEJ2X3c2?_G.2Z</H@H3A\3
Y]RE5g\O^37\[9DX/e#?VYN/V4Ff>#@S;RcI:.fb-_e@>^a51\#Y4D1g:CdbJJ.O
KO6fLeWMH7TfdI9dfP]]MD7WIC+b[.U-LE.>]AXETH(P2JM8UCUe^TJWgWXAeIGE
L\N>?ce8=-P[Lf]UCA8\Ubfe)0)J54N#dC(XJBN[=K?SC)Ua+ef25C0^dAW2U@M8
V,OQOX&-OFV,^@>KJWAH+DP2L]HR6\EU:3UA,DP:?\(gd@B@_S<a,IYP;(5Gb1+Y
U@S=3+cV:@(8(_)1DIOQYW^GFL(&O?J,W9g8gJcP[23U_P&KVADG8J6J]YW4T(O4
DSY2]>X8V?D?)^J#80/8>)7+M0.HIH#H]:BZ0a@WHT47TK#6&=F>&+)8ZC(c8+KD
<##D9,EWA7P[:@eYG&JCW[PLUMQFUeT]6SD@V-?2g/aG;=eRb2#8A>V8R2A9&a<R
Ha@a9CIH(8F[V/BLTfL09Z^bL?[()R:?RWVYLDGa;8G0)E?K65TF&Ha]#Y#N=CTM
_@VR6>UDG;TPbUJ+?3DWcbAC..I^BO,DR^6\THZgNOKg<6aBMRG33-=3;B5_HZ+Q
D#[LDYcVA]R^RYV?(:&J:-X7Vd,&20.LX#QJ+&+e7I-d#0@/[@F#C,P33J=ZUgLa
VM:beXPZML[1M)[9A=PZ9(RF.GQN)Ad@LUA#R0:>R@DF^Z0BJ.a0cZD0E[FM4F))
b?a28fU\)=Fd=?a?f#Z<ZM)6:1?gM=XYN7SFE^aCV(EVZ@?@+&g[CJM^0REKPJ=K
2We,f&NZN4:d&0]V:1<92<QRY\(a683H8>#_g^:PN/@@QDAZE8[]S)E?YAa)7d8#
0fIT7^)TJK#_;Z:b?:CZcO=ZCI+4G/=9cXP/47D@cIMR[HLO(0<&(SgKYON?f#TW
g51QKL=7G+f.A7=#EOQ#82,X(@TgS8]@a/J=S:g)]QQLLc1TCCI?)RLZL.#Y/bGO
gX4IB.,f>@_4+I9+NaOU]Wc?GCNLMb/Q,EbHG&ObPfUUN,KdaA/=MA#J.;5F/12g
>L-/-^2>P:f409E,:<\6GUc?E5J+4]>AYe>VN9aLc-8UZ&EN:]#9I8,>?[H:ceG1
MK=2J9HXWWTB8+-<ZYC_8Y\RWQ-M9EWW4TG+4IS5+72QSfFT2JacXgW9QX&9ILFI
\)_,Qg3XC4J-NJ#4H;4RB3)_gU,?8<d\X8WX&[Sb[/d7@d>G6>4LNII(\,fEHJ3=
?K[0;8&8TR8dFUc&6O=FOc7UgN[O.g_=aZ4LT5BK[26VGY:]NSTYH_GYDF9DegSQ
WUGX9:.&O5;g/bOON0KP;0S;=V8)GJ8U>0-W4ZQ+CG?&1e?bON15&6VZ#Y([C]gg
[>fHDZ/)S#12S1(,L[/6.;P_XXbdTV.g(aeH\eYW)2COCcPTZ^<_CHcHDN44deH/
aM\GX+dHUITL/Xd(V(]6E-Ea(56+\,bBJG058O_NDF-NTeA7V17.dLFIC2;<CAfK
7eLPF5O]?LNMMcb9+SRLa[YZ@H^J1bB0a1RTC@4D-\:]=FPZO99XW\H\3I_9_X:+
IP6HH\aS-fHDY65fE3K_&21cGQ^:0XZ]Z1MV\dFK+?2+SY6#SZ9=OB-3dT-bfY\.
PAg^&N:7AV/#IW:5&dJ=&1M>)^MB6TBGXZ4Ob>f6@,KI,>S3(F&GcEAXa(bg=47R
16L&gfVYJ)5V5+C]^@4UP_F^e5]gG[cY6T;(#.HZBYQ+B,g+F3^Y0JQ(,Xe;c\(V
\L:&>:^P<5d2\_>KVT[AYfWdS,[WKMcKH[U<?cc/9(YS9]1.Q^U1-6H+EW;M_FWC
+V7(]<N_P<BLTP,(cP0CV+WRZ;bbU6G26>]YWU7IKA@RJD;#5>94Z<P,1EAY3UIB
?L>C:\3NeZYE?&;^M8=B?]>f\1)5f3;Q^\XSaJGTH:Aa?X/gWM>@7-LG>b/FTYBe
/DUMC/5S5V,CAMe6R+JgI6Ie(_)CKS3-g6.84P;dTcDU>-,E5gg66HUa7H_egb5O
>@fUaL=gKIQFW37?If=XaJGCPQKO)H9VA#C]=fbUR@,T:K[HY^Za2C_NX=R;X:-c
^(9^#5JbX9_Ef-+Cg.OZ;;P5VWL=Z?K\V,)1I6L4/F\g[OB/?X4HX5I3&Oe@#WeU
)<_@#6F4#VdRCUDM1WbC[-\Q_5^DD).N[N1G.OS[2J=:+2@FLDgLZaRDBS=F@<@\
dPC1H6CYIg+5O1;7UeIdD2LJKeMLBS5P0dE=?^ReKBJWXX0#I@Q&Sd@(cHPY-8bY
/N;W(]SQP,@E@gGW2,Ca-361HG:,Ddf]Z]fbObT^I<SS:5G^Zg843IM/2Z>RP7cP
U]D[d),6NX2UN(4(2QR(Ja^dR;Q^b^=5H<?2bIZ5b6aHYDcX0NBKEg-gRSSC^gg]
MS/f&YFNLFO+dG8+^@DQe]a\794KDPN/+NT54b;2S:ZHN)KXcbg:bFMHC4R&A=Pb
A(Xe>ECCJJe2Jc>,+bg)7G#8F@/@<UU[F_,5RYM^J/d@<Ud?CBg@_3IZ9QT0=2@M
Ec&((>6YJ:9A;+#>)&4R3U#FW#dLN<5U1PAb<BACf@A5UD&K&fRC8_EPeGI]\-.\
YI/9@HU7A(>&@YP.9\Q2SdZe/R\ba6Z&cJM:<O#W.Wc5C:L/OgKT\_QM@P:dB7FW
38#a;af:#K]4>LPP:/B:-e-9a.d]R8F-(.SQ8C].2,P+[Xg)E[^3)P^W,F0\0;a(
O\BQG://ReJH:<E^_8[;Ua0NQ<fF@XGV20^(M/P>XLMHGe8HRJ^BIHc:cf2gIX,[
ZfS(@F_FYMfS4KaeB<g+eFAdS<>_K=Y_4HR0Tc)8^:bWFM)U(AZK^#;f(E>I4>,4
H&NHDGfaMIZ\H3fEC7.Vd=:badTNA\UcgUP\gJX^O,7EC+9W28e3CZ[@&U,3ZZ)L
HSJMG:VgaKOB4V[.5dJTPgB+L=JPLg>XZQ7fe2P;Gb<@ZX5XK5K(7DCd&fG8]FRV
9)H3UHDA@NAgg-3#OC2,W_Z08[0VdEM+KZ_FM_BdHK\5I#RS=P>E:fCG95:eHdHL
=E>LH;>aWgGQObWHgC.Vc_)B53:.FR7OH=_7O\/QSAa.NG=+45Q^4(=14&+Q2:K,
cd@3?N8YGP(eG6FeNC&->-7U?JY+3>1@/&&C<cP,ED(gH<Q1S\HF)[J;[+R+E/.M
(g?e0U5+\1_M^<aYZ<faC-^BKU?]8R)P;:.gELQ176\:PO#55V5+GD1LB?4K6AKX
\=fKH+6._J0NTX)BfAPZQ1&6eY,gfG9f4O0e6Y/cKDR5\0A?(VB8C3\8T6C7U6MO
)4KJK6&7fITaDYJ1WcZ?))Zd[@M@=MELTfK\6:4.?E36g6eTN[I97&)\J>)KAY@D
8E3YZD<3ZI\@GOBK4A>P<\=#dGG#4bY,_6EgOO1aJ8]/5T(MGBbJ)S3?1YA)6-D5
/O]R83+9WG-X3[0F1\I785@QMfK]EL?aHEXV);82gc.cZO9a]SG0_0)^7FZU+bDZ
\KCKU)PWg_DRYJUVU13436:93-[gc;H,O(1D#1/TT.SAAdI^,#@BXXI4XUeaT__)
,6JJLHZS/A/A?d_=6M5O7bgNP;2]YPR0P]0=1<-60,/H2,A+J)S>(_9c,-/(,J5b
]S5FX)@fc#9]5KWDU^L(OX@M\3S>@_9B<:.@PPW;g)8fWT/:c10<<MW_+T81M@_^
bQS7af5dHZ:XL.:[.Z5.]N]1W>H:V9dedf^NL:Dd;,X3W0DH2C#dP\J9?;S;3P3B
=eQL=VS@3:5NG1IgJ\RM_RU3L>3g1eb6cNKKaedBA0I3QJRWE-dW#1T-3@gXKgae
6&8S:OL>.RKT&P1/[?bHV)C39HG@a29I0Ub1JJaQf,KN8Mg#X;/UTXM:g2\HH\,<
Rd;8WJMbMJgV)&A#E)]+7=Q]&.WK3U9J7ZC>:8,/7N\ORLN,.36:bb3X<1VHUYUc
+eB<(]451e;0#K_CK4.^NSc/F<\;@bB>APIU)X>J)+S\GB\M-SZYcc/(>RTa:V70
WI/^+@TI1C=#28VJ6<_X-@HAUe<Z]LWCB^dQ/NVOH-H7YY.1<#/SB]:IKK8#]B#B
02=b;9X&X;MX7,1DdRI>J?A2)EIN])-7b6ZR07<74Q5][BH/1XF?AA/R^]/bS&8Q
73)d(>\=Q^/;f+D)SZ,B]UX\d\4@:bDS08]-#f8b03V/^S(c,&O-1:^R/^(XDGVM
&46>a&+[7,gSa[;@LUNGW#0^VGK4B@(1DS:^.17U)M9/f]2KQ+5bK?R_d_/ggab:
/;L<1b1<cOe58@[9I)P7=c7eXP#DG(56XQ=V7F=.:>&69JSe>G7DI#FOY1/e8K-.
ea1)YNG&^-L15:BXK6=2Xa_X?&KD@d#\CK[A;e9VUd9;NQ0_BNgD,)236J4AAWKC
YE&=gKcc+K@LLCLRXJUUd9PQF\+)fFQTI)dS1N[08>58/>e#-AU?P;@&,<a0#O&d
0=GM-WV7#M6Lb05-4d&eYTVAXG)6e2[.SNO\[/L\O@&Sd>a;OgAd_]=Za)cKBELS
1<MgIec]N_V)#X4&Y2_Ze?R#:UI;&N<IQB:N9Gg&)G69C06<7B;7e;J-G6(,SDWK
]_P]J+FKVb<KFc6QO)K)RBYJ.PCgc.WZY-(7@Qe+QA5EECF]2I5+S91=R7A&6R&L
dY&W[,DIddH>#DZ[:?BIaJ_8F@gSNX;LS,cQNa(G(9I-H@PfG.?BN:cB+=PVQg?B
NZeGQ0VSXNDDNSFQ<02/CXUKfgCA\4)Eb27OaKZ0TCa0@FLPTN&&BW&6A/aJ6KBG
LA6B22C>D[FV8.[,gJT=MH=\CS^S#cYb:S,6_QOL@aBM1BBWVDH[E4T^MVQ+Y.>b
UaAc64\>c24D:3[LMOX3cC,Z_e3C>D,U<8gfT\R.f^>6DdP>U[f&\B7V7-a2\3eA
@R^_U:BL<^(M/fc0XTd+RJTEU&5)JD1J73GU>JQS1_TA-;U.20->12I8U#)0\9>R
]99a,6CPV]D,-&/#MFYP..Y.LfdbVG@EW.H.YFLgV-bC=2L>R]&MB+:6Q9J-.4Y8
29MB1PK1g:E]QB[ca+AdeT<ga0c4?SdH<7DF@NH]eKAH0YgFRBRD<#\f50>E;8F#
.2+AGMFR1T[@IJO#O01f+[BQ8-b#+eXH7Md@e2&+<WI479UKfWK>OEEF6GUJbZ^J
bP&1XeZ4FS26:@c1PZK7fF)2,4JYdWLU=<NQUcFf+Ka2BNORNA#646M[[4.TF\K>
g)ZP(5MQG#X_1(C:OFfcLV140ffSLXKQR8dAKe5/8c6/M;/K07@.5OVFUfO==D^3
4Y:L4:EM>X<DZ-5#@eXU@[J5++><O7;?F<83+gYdcg(45_@)OG7_9IfZ^cbB18gC
K.T&_KdH+YQ91&()BTD#W#6#H0J_DN0O93RC&OH@67:[H/6BXcIA>MgZ9HfdI8N0
M8.EV:Ef_f]NFY);+=TF(B2(98^:fa71\cXGSe4QQK^C>R>a:@K_P(W_KIX//I0#
-Y4RBLaa7#;d7Z4VY/eC1(NQ,S-4C@(W37Q^X8RXY/[(5\U:4Ncg).eXRE-^0(_-
\#Z@QMGQ@Y2Me12T;5#B[B(\QPHUb/#2;P8HI:MNK0,X=5NL11L^?g1UVQ4SQ@EG
2PZf_EW+[..<>PQ\N0L0AU4[I(&@PV8/[Z5]#2\A-]@@8=]P@N?HI-_ACfaVDPd@
R;CBILHFH-(+0:77a;(5TM,/T+<+#<M[2]=+Jf_^\BP8[7@CfJ)ZZDH:=gc2]I;>
F0XB/RBb58Jc1?A3GYI<fDPET>8MJ]A\g](S91O/X/LN+?PDFB4GJ9,DKc[Lc7@I
[9a\&IP\^d\6D>JP3]0V[0I58A)CVAT[.Qb:CY?@L+A5EdODUDL>bJ3HR@Y)#0M)
]Xa1VV.)74^_4;]U>LD4BM>Q&Jb+,6LgT6[G^,dB5G4\\H3(:^Z]H4_Pc.B(5CdY
G0bI)_^[J[YMIA72&^&Ye:SE1L.UTc860OML5<./DK^)-g8EIa4<8a[SYd:JBO67
6>eO9BR(g8AD=[>L[3MOC-dZ4?.5UUQ->Q]ORFe64@.Z0<efU7>7;e&8SDGKOZ5Z
e7bJCU_387JF0_LIV0bR+6J^@PG[#9cSI4B39#1W22XA[CT=cVFOP#f=5=I;H?C&
eFP/<0:GI)Na8FaS+-9>HNQ,K[,43b.66cgZ^,7ED&dEXNOLK.>S&^U;EPG2agAQ
Qc0;dKUX/V2UNa788EaG@-Pd8<=R8U=_dB@O?I24&AN<WB?SQc9>[;VfUF^\>Bd6
09UBVY)2M#U@N1aN3(?=K;2[Ge7,OQ1daUL/0fB)#@9[&cC7X8RUg0]-#R/f9>XX
d&L=c)PVcAD7J5OPcP:c9FF3]MGcePAJBC1gf-bU]E,RSG?\dX0G/XbPL>MYQ2CP
13C(cUG(V^A;EWgdCbXD)<HQRcF=MQ(\+U&92.#F:5_,[_MY2R#F<1=7]H;BL:b:
R[YV<MCcXJ8/\e?.FeF=b7Y\2J+4a\A(2T(3.YN3.)-WaUc>@A9@J453#YbQUAa[
81DY>[J7[Pe]:HZV@.f&3K=CMXN6=fC,H]0Ff4_7>a\fZZ3IA^?PLIT[:?SVHM]g
3_CS@K<dD9321_6N_R5.6NPG0Ga&TM)\38FZGD-.9]O&4f,RYM^ME_FE&#F0^]/&
;?>?[6:2XHWIQ1.C^bMfMZ0U;fAP>RO<OW92FP,b8UUF4b=BK2.XZ-M0fD_Sd#3Z
V[E6EW&\.-CB/MCeSJEDER),>_Q-E/&DSDA-I+=I3T]<(&-N,RGcGb##X<RF-EY/
9>dEfJ+NBeI9@JJdR9cTM.:gRZ5bAENGgP\[5;E=JbK92H1dP8S?OcRXZDeMa=M8
2LHP(5SG+)9f_\6&\4B-T9BU=U^eUcIQ)Lgf>HOJJ].U^4(0fePD]DA22A\A+JFg
YVW4Ig7I77>Q3_I9VA[>\,(15M-=V)DGZXWRU]5X/Fc741]VJMb#:WF+XY^:4Ocb
e#2d2&#<-?dFA8Z4C3NTF(Fg7][T\K<>&=Y-7V:Med^&f^fe66SDb2KJ)gI>bDZR
NaO>G<5;DR<K^Y.K1+,X-7W:>&[(M+Hc\eg5fKgW;(VDMB3K]Lf:J5:VZ3G&UQK4
?^\37=<:+Z51J7S,Y0[3#\IQTEVBL6b1AcA-,E/#GbE23&M:XaaQ?E>-F(ZfO81F
0IHK66:O,K7YJ@XaXc77#UfB>L=a6^H7XfLQ33\.XS-PaO<f>Q1==J_PFL,PL&EA
3]+Yg@1Z(AI&KPW_SeBVaF,(I=@,]#aQROaW_;-N.7Z7;+(@\7==NRE)+FCM36[b
HbJ?8/2:[aU?W31ZEaPZ#8@],3N#8F4S-94;8a<&O:HAOYH2B0BK+WD\&Y#+HPG]
Ke1?HV95[,;@GgeUR_K13_TT/a?A^f[Hf2@;L8c1@-)93]Pba[_8C4\(J_&ULG?H
1-dY-RS:Tg?PKeW-VL5H0)&T38>NBDI.9D(7W3ZPcE)U+\g)02a?8/LBYU0BI7H)
De@gA#<>5/;6XFR>Ba+NV1,V&4W#40.D72[@SC591/Q_HW,1S_8R-<Z&.Y5=)-Ef
>dDDZ2gY-W_:,d,YC-M7JL&OV^;P0^NBJfGMSLW7M09fM6AU<c?2CWCWRcK<ga+.
K5CL8KE:&.2N_C=^dBHS-WB;f15NT;)UMQ?(5;HHgDGGN-:.AdT<b&8_#bS&c.e2
)OCD]g?Rc?;^g0_8a,+A8dKaK+<];(S(FPINQSQ7&R>eEU#ND4g,d9a0Q=<dSf62
:C1E>>3Zd<Cd:I[g]G6[^dAJaCd#DA1;F&(ZGZSf<2MJVWIXI4^8F3G8(M[V\2HZ
Z>LdXB_eXWCNZAQcUZ]\R),fEU@RR1-](.WXe+KQ1:Wg@I8G3@KQ&[4_8OP[ZTD.
?-OPQ77+BLP716.X8Rc/G#CXS&FOe5,R6Z:(;c1FS;HBDYIf?3VUTTT_&V2AT(1d
]I9+4YJ1&JPf,IL-,^@a]G/We4:8ZbHYa.:A+aNb]EF9=Ka+_1H;I1_3R[^]g^;Y
T=F@Q([[:A>=e0,FEGeW@dQALAXI[H/OWb6D:@bb,ETE)W23P7a)S0YX..G6&E#D
UeOe3@_MJd25^:)V,MJIC/-1L5Of@^I@4cQ]/b9(R9<,b9,2?8#DMV92TM]^0D@U
HBYP+]?Ke)6T&d7E&\/gK?VZc1X0Fc.JbE9:K47))Z#0H^RS,C\BWe@P/1@:gdV7
4a-:PT1J+BE7W/fZcf;,6JLeV(P&-1TVfV1c6TT\]<NAg&#QA&>B@=>Y7<#X>UW7
/XJWH\TNf_@ZOYM#4d3JF:@UK&bG>N-\1)B.@IP;^^FFZC6S)E(Qg+Qg?HKT.:6-
aRT,Q&W?R)WBF3\H]Ze6LYNJa@d2BLGZH+,[S@2W#.e\S(JMS)X=PMa5O\3(faa&
A<GGI@?=L#ffFGT&)g0>+6?KG0@EMN;,ILO>@R;AYOA\X^Y,51M\A@94X@-F^N06
=TS@:DV#2S&M9A7^;eP\ffFVP:GF^7JQdT17gJ,)Ba3UDUcA;ETCIQ0D#Z[8_UE<
dMI1Y]dcX:[(HF>e=YXfY?4a5,faKJD6.3)e#;Rdb.-K()8=G=3;;1F2-_^,>K2I
@DE-BGUG\EU_?EE@Bb2DZg(3_d:O+8>1C82ZOP[,)]5Ra\D7Xe]@8P[0R#)7]H>G
&[/cJf8].#;\FTa7\7-_-&&^D[=^9b@;:&\dE&D(fQ/M#50_:NUN+8JQC=B^Z,Zf
-Mf(e53WIdJI75NEa\;^92QICA37(@WSaR]D(#7;,@G]QQ>RR8CI?3DU5CI>T7#Y
@eLW,4[1A+b555J2:IM=fU_>;WTU]QD)B6?c)\&9cBX:&Y<DH;HYV2B2:I:dW<6K
5>1YaS..6Te+3;bE[E&QQ+-?CDPXDH;Tc,6.VNMg.1.dRE9/WT--Fb]e>I(6O+0<
YcbN4+0Y8[Q[ZB=VA;41EP(UT>FXg[fKR8F@W43551;NM.88\U\g>]?FYAL;WHN-
-:LM2;)#I3gIGOC@<:gJbS3I??2]([bcUT96)3e_[-a@#-<.3V3\BSS_MQ@LBCSg
VE8SR)\&gf7Mc-g+IPN4TSD@Ga;KD-)LIK1WPFD-1];08[[94@Z0<@f/_+]O][U)
b/FW:@G.:<O=UP^#@@QT/:N(^8[2V_N(HJ-P_M4P_cIN<5fY?KQ^bP11?FgT11W)
7Re[IXfXCM_YSa6-N)T#FT&&A[2fC^;Ac(K.T>X&#K;9)[FBZA8]+cXPC-APf8+<
2VP6I83RG-JF_^F@[DMZ17[R?6#_VePR^_5/I?6@XGNP62]5J5EW8AU[H7E::7I[
cf8MeM9:7F3[ECB@W(IZP/?c^)]4cA0=cM1+--^fO?C-<Q9=.QUIWU1FN]eU@GAR
)HIXV_I9#O&6;9e5X?77.bSMaa\6UZR:HG)?36833&>9+bC0:T8:YVKW.&-]-]/&
VAf3B+DK]T4C7=NDM;:4]^S?33bKGNRgJBZED\\NAWKC.Mf&0[P;J=,(K4G:LG27
&eBQJ9:[[Ra/O<a.AS83:F+7,K_-IcL3MJR<^62UGM\VB>GS&[:QGbJB8CL7]-/I
e<3K<DM5\+4-7]W4]-4RVA=WaXC_OYQJF2@_e7Z8G5E,g<JN7>R;WS@^EMf>B;+N
??^XZ-RB#0bXYgRMTeRg50c7bD0I?PGFIU,^GZ?5J)/L0<GD/=&TI]-)K=[175g>
F:PJ8/Wc(JQ2Q0/e?cbZRK=I-3\G/89.?@gWP?Z/cB]N?T3@\<0EHZ_23D)28A(3
/IQ,Nb@?2YB<,2?YFYYS5VQg&3GVJ?dae-29,\[>Z+R]>GEV/C=--UI3+@/Pf_^M
Z7+5fCF^Ka49T1#_99@OWd4NW.a.4G]2-[R+g0K;.cRX?#B&Y&A@J;YS5:?Q23b0
&YQa0cYY6?7gd4W6IU&/),VVW509gB-6IY(V8-C;8H1=9I-=]gJW+GE8eaSL6Y77
Y_/@bPZ,b^]#WD5IeQRG.L^O-FT&JN+0U1AF+)O<YH6++53+W?;KM:@fKSVf89QX
56\YU9R[OWQ^PRe4_X@WVK#1LK>Na;>Z[;Se?H:9>6S0TObaO:7WI4d&39SK+Y#g
Ba6SfN/1WS=_)XfZPUae71C^,#gFaHE@K>X11J&f767UaVg1G[#DW@Ve&-CUd8dN
P70Rf&.YO)MO40e:g]9b0aXA<QTF><AHZ<a.E&VW&XC9X.+LZ]AH>8J)@_9)f/Xg
0[?GJ(&K\;7+_P9SDd/C.HK=&/eHG&ffD+L[L9Q_F]IaUCC=/FTgB3R=;3a?>7@B
Y7>1=]31c=IFQ#5(@@LH/4SZ;gP3G>49#I39N/OQ6^;7Ke;e2#OMVI.MBf#bZ2@=
X9PS0Q@0GSKB^ZA(KL4L=Z1D6#[+cdUD:X._KK6eXDRT@FPXCC-O-,XV:)Pf4\Y,
/Jg\=3[O8P45]C<GU:XQcGN@WM#DbS5TXfOWT8/da3+e<VcS\Xg,B)GEDG1eW2>(
ZH1gK@KN[[c+A#QIXbQ?&)^He^)L=fBX<++03]NCN\9#^AK_>ffPe;JUVb3d5\C,
DD[R_K-Dc1\Ia7D5FOM+0&94;Qf+Z-+-/.@M^(Ib#<&,<DO:-ZTe(]#@_FD^@RJ=
f3e@CO8>2C-bLKF_GRf=/?H7b3^I[b8[K8,;+<4DR,AT-R<K##MM&Wb@YIf5;;Ve
5,UM;0ZL87,78]OZ^AY][]MGfc=?=TX;MC1N0BYZ?&cK&-:O]4X4f7](M;0X5+O0
PC\e<VEN.#0_GT@M&.38\A3WIAA7J,1?TO)<Xf.7L#Ygf_C[-(E@a@CLF(9[36M7
Ld)#69b6:>-@I304GbgbO@@I:cZ-Oa_0H2.UA1b&/WEI^&=]VVAb4K,>H^M6N(\O
c0&)-4I06\,.R]2T)B)WXN.I&6O.B9(HKaJ=+,=^)&N1,-P/+KIQ(2cQ_aU8WG#f
US)>RaZXT)13XQP3ec9aCPXDBD;.GDZ9c?0/T^c&@<FPPFW1#XD4[_5.W<K3CO/>
1ZD#2DL3X?dHCB=#AIWIX[[:g/EP&T3Z6FI1YI=VfJ4(e?/SFGG4&9;=;^Ae)OZ\
f=RY\_)\=^D]>7;QE]gKRUT&Qg-Y9;8(B=Q&J6c_Q(H[6fS6++6VN@U9D9PM/HbU
]<=c7+gM:]\BE/JJ@RZL-]&#c@3cQ,@>1,SHYB@5#C&d\BcQSU>C-C<]MKBa;D98
92L/RBXf\.UAY];Z=0G52+1Q70-9?O),T1Lfe6Y;[,&:@(;MEPUJ];.4P1R3[gWL
Mc]b4)g+()2dd[^SX#;HHEMdHH<Z>&F-BCYe8.-3c=0,Ug>9FVZ+Q?5aEFHCg8a;
0g]RS?#S<V;V?&-W4bDTUTAVG]_fN]=J.(WZP?]KDRa2(G9=7;1^dF?]ecN4<+3V
M._+3MK[.U:5,?Z)EF_C2;W>\<.Pg7BcIT8=P)[#[Sa\?ZJg1,[<@b205H,VfQ(9
+]LF=-Pf:17:DYAC]dfb1+EQZ7R4-XZ2>U.5;bFX(Ad/M[S7:H\5FJ74#V?ZNGY(
-BeM43VBBO9UdIJ3eS)-)b,[Z5/eJT,GUB07CLD,\F_R)_MKTO=FS@TB&FSQM?LJ
C4cL/8g@LQ<9SScB2AWgWHFJ?I,5]77UP64]9(eT8cS,6V[RM8MTR_Z:J6B89=+a
\@H(5F=(>N.B<]eYZ1TFJV90gS8SIfN488QJ0JI]F;g6e#A?KZZ_cRd+LV0EPT:)
XcJVd/G1X6HQCgAc<_f8R4eW0gY9H:fV:EQ,V,P#O8?AHQ[9V+V,/b+OPPc+3?N#
dTdYf+/E9/,=CfC6)9eZ3S_5A+G)/fC__D.;MOe;IEO;S0#(EPZ/CTa:R0dP1K@\
Y)fB(?a9ZKabCDB=/UB#K]=6WFC6R-d.^^Y##W+,@WU],4E^bE+8<PHE3ScKM&+[
RNgLGd?^=E)M7f=KO1Nb@/K)VJ^F2Gf9(S9.JD;XYK=]7MJ0Q3PR.F7aN:..b,^@
@W3>.6(\\YB5F0]HPOdR?3+++VDJ<365#0C^K1+d6TKHe<M&N6?CA[MRfD++[W\8
]]fe&Wbc0BOLPa#?1T@SEWJE\IH@IR6OR=cK)J5;;9](WgJ<f+M)XA((5PMT=07Y
^?RY7I&X<G9LB?JE@N#GNXLcBSEV[<UO[ENgE0]91gG.4:LDN1DYL]7D,]&0A2U.
@#U)]Yc1dPTZKc&QI@gUJ2[4T^MX1X38TOM1aKP/6[CG[Z,_Kagg7MfFR;390G0W
K)QSKCB/A6HC_ZXRCb9M@6,J7,#cgfF^C><(.4NU>-bg-N(S:GG3NB#+2)AB8Ee<
(19OffK?fa>+Z75_5[3V_K__(+8DF<,QI]8J21F9/F85L?K2V<OSgJ>cgHKb8KdI
=QQ3d7K=gD3/8FXe;3U;SMYH:9<)^NdWV\&=1d,=/SYAdDXR38@[I6U/;2B-gN[1
,G2SYZDP6D(Y70ZOaa-IaLCTc2;=8<BeY#:DT&4aCVY01:MIQD2>)</)e7.AAKH3
]+(gb-gQ#5>Z=3TY>g.&)_UE,]85Kdf7N4(/,0F77WH#;],?f-#ABD?PBH,NO=TY
HZFef_HY=48ZAF+_YbW[9g@_X9DW/0?RR&&9I750PO+R0R:Y5DeaM2)?R0C02PY5
G=B,#V&ORTE2=/>:G-:GSEJc+8W#:&__)g;c+W3P>3[8fR57V?cO^QgcS?6]I?+E
YbFY.QdXG\e&2F61F-YP>G2>/0:Y3]gef2.;1O?^d/OY3]<7a:EC&T-ZL-.9<aD;
SY5d/gd<QK19Tb=,gJKMV=#7V.8e;-HPMG^0TT(:&,XN0(:0Ib6.([/PP4/9C]DB
^3dI+F0P-:DQ+XNEUP021S=ZeMcVU;.,UQFg5EB?S+30@4-+_Xg@HgfYdRe-ZI_/
_,KLA>c?#+9TB3ABK8a?KBF0Y8Y[;L)N8<bgdWYA.:eeY?D<S7a>cCUW0#W(eC=8
KK?f+I0X:H)-eTfQ3\B:]4&DGZ\3L7[cIe3XFPZ.e.RZS8-4\A<>:^-CXPARZEPC
ba:OI2=0ZUWXN\G)OHJ7GF\b+=W=YM.e+d_a@\eSM\I2=_WA>D,QK0YKF[67/R_P
;AWI1NE1Jf8;JWXCc.R65A7(?^P2HQ&T08bE;fQ1U7M/)0(#aBK)D>e2g]K[(0I\
D;Q6b/4=HKQN?^^D64(YdQ)5<=Wf.D<?LTF_]+Fc,SR-5cJP&R.I+O>@8FH-X[@C
)[Af]^a>SJ@FDL5(H-6/-)f]ePGL0BAcOYW.).0DD#P5((2:BN\I0HXV/3==,VD6
0>>5^7--ecC&\W?dR&?CV;[=4FH5NbXY;;^K22YDA8DD?@XBSd2,@++&18dTPA/R
QfD42@U-2:>X5/L>L>L&9;6dV1#S9d-R[1WZ7>4b1F[/K5<^=b5Xa(WY/f5-K5O_
c,_U\T/XUA11YdMLce5.:J9QZ(J=d1:\fQJ-=W;:>G1R=E7=7F<[-Q8_Ta:J>MbM
&Y.U?aTJI3V_U6\V[B.8N[VO5Z)5<;AEc&8?[@#EPXaLU_T=QffG2E:&Y?:C(ZX<
D=1P@f.EK8W))7IF0B;#^6Y9>D:,RdEP(VDWP-;Q8>1<R7YCOILHH]F,fc)^LK).
WgddH>fFA@FfL)8gY=^QZ9TLUbg-YC&TJf_Qe[U-^D?AZV_T)EJeG5KN5d>+V(c3
Od<5P(.PE?+MII<RW9W#S:&W>/P/T[G\B&GRL6YCV<14RN?c)6gb(03V5db=6__e
dYfD3cRY\6=F2OW)P2179TFZ/OB2WUKV9.=6Kf.HcV@Q.:?L4ETI/d;8;]Ff-g]B
^aUG]Sc#H7Z)3Wg(Geg?38cY^41KMb_Jaf--K+LCIL,4_1d3LFaC,:e8SEUW?X=G
OA0-#:VeRg0JU84OIZ3#],D8bL0bPNG>;4JXe.27HM]5H5d-,:C.?T(5C#gbVS?]
@293Dd:?]PM+NMSO0?VQ1@DIMPS4(>?738)CM4BQZQ,1^c3O0?a?7EAZ_GO.?XdG
?0UW5A?B#?;W;4DBNe>QZYN#[ae/FHT>XG55X23AGG_[T2GB[JA.B&>0)#g97#b^
<9UPIXLF]7<;U53;>066.-@3VG4,G09?C^RPU&^5ZDef1Q.;MQ3ba.)Mg+,,g>eE
FW?f:>F#-QWe#65PA928^f;I&5,P+F-g0K(AX-)8X#93>Ld<OfD;3K1C#>G;[eU@
&SG+/O#V?WYBAOd6M^S2:Uc[1/KLU0E341_g\M&3g<N-QJHbMUFR7@aL5#YX9Eb<
KfYbBG9^QC;)+UCYgIC3UAe0[B]fXD@B;GX-cR78_:c4<ODWIC+X>QZ&1.3])TW.
EB##7LN=:;06151Of><^.^NTCCT#957>&?KS1E;IOg?12D@BU<XbM)>J<g65cV)2
G&N?;&\)X08J6Q&A#@G[2CQGNZRWXO6;,I.L-D6W\&Ug.H\8<VRQ@?fFH>B0I)\6
WcM:/:D2]C)D=JK:D&eIU6e</2f3<H1_\^PVP8YH:=88(N2S<>e?PJ)\cI)c[4PB
LVTTCXB@4Ne@6NA]K56K](#7Q<J&A0O2If]+9/OKbGcDL1_/Ub[WA_>_C(NAO41-
WUWOY&6E^3GUdNUMB98G7fRH>J^d:?MYb]MDEgTN_L/KRB/Q_>]0D/20<++XHQV#
T)f:DS9d#F&(.J61P#@9DMa,W)a/QHF-Jd=;DU(92(IG_RXN]&-f)^>eMG>2dAKP
@6e_V9Lb=e^f8B5#8#J1?Tc<DCU=F=,Y0CAF=NOH67G:O58g-WTP#?H>2g;MW+W;
b\#VQBP^>dg_W9=ZbPPX8MI5(AI29Cd+LY)^/]YeGV^6B+DT](]S_A7ebf/NSc.4
[@2Eb+\#S:)BS)03^:DXCE5a#>]d&1)3MKQLRHE3@.bRcgB#fa,&=e9O4BN>d[:c
KM+<Q<c@E,EGZ7\[>Y?&IeJaEGX>0L>20??(P:_TAS#c=/RKbW/0[Dgc)V:0O_^K
<[2V(RTF?#[88I<\4Y9R2IPCP2XG.D=S)=4V2<@WEU,#OF6c=1GXD[gM@.BE<UGG
3&a.>ZT[c8NZ(.:KPUG-M>QUV=O^F36eMN/F1_7[Uag#OKd#XE^bQ_9,JHHgG?SG
X_#C&//3LMfSDA.KMMUMc.D]Ea_af@T[^:B^735FA/&g:g9CaL[7D[6O(N4H^9/<
Y3<&?(&#W](1;?ObB?@(QQ#K/4?#ECH>QL.?-SaO;>4NWW,?_#6CNfJLN^K>eb&E
Q60\6PdOg;PVUQGYRMUb<,2<A+:P&f[L-C^T-eP[TV2]<+@S0T.4P_3Ia,)D^0@0
T303OYT2A->?Ng;LKB^=^<:NEdYX&@fQKC,D5MZ[:>V^cT):F@EJE#RbE@91DAbB
7_YMSN#]faN,IA@dTKJB_N3NXR\8/N8^(7P^Ob=>2L^Fc5,L?Fd,_=)#UV8+bWM7
1IZ_8/4g6=G,P=a_:U0^^1[#:D)EM;X8)3DV)G^S>K&YQZY(a]AS86=f.J?/(?1)
2X4-f)/HdO1K4UY6^G7Df4AWR\SEgQFUHTPe<OZ:cBc&VJ?G,Jb28X?2.PU\W8,e
,JaCdGF10U37^BKQ@.F</4,U):/3]N6@X>ZI-Ic2UNSF<<[gA<:S74gFLI,L4,gO
1?9:V(.+LLOV/KQ#(&YLbKaQb?YV#5F])0/HSR#/-,0#<6H@\JX92U6eDWSZ:=(c
,S-V+;3SG&#5?WP3U=bY[BQ_85fYJ\?bg/Ag^UPB]e42L4(K1afg/N9XLab9,HMe
1SU=N]@,#S-0cLL[\JL/0QO.@&WfIS8Zc9_V@Zf38SfQ>?,?V2.=-GE]O0gZfHID
E0gQ,;^)IA]Ofb=d95:G8_Z,E(?>,EQdXZ@=UWB\Z-/A-Bd62Fc&DUW54cE=O1\J
PUE9JSZeAHgOB5HK=HP?MT49(V>3AVC:8S:g?S-OeMMe0XIg#>(^/3IbO/R^\BdJ
><1Lb/b)]6e\^0eS61SS2\PZ-A/:.L)AZG?WLB,FH+)ca,;+FDff^(?AeSQJ(T^Y
a@,;Yc^:dJS=C\0M,_+72W5UVM-^bC.F.dFV-bGReWE9?VT)4?L\R//&cJ9IWL-7
6_X]NQ=ASJ;b8[Y0P/&TX)fE&OEU\.=SJG#T7W\U4+GALQ7/Jb[I8UF.X/6WdR._
UR5PUIe4P58<T:5&15?K^39\PaFcc[6X4YO:,X=NVK\[#U48cA\K-a(YFFHR17AT
M_g3W<YX].6>R#6B20QS.gX.0d@XPeOB:0RA<bTNEe5@&JZW?C<I[Q3JgV.OS]DI
#4eB</f9TbfedP2f#/(>V>:EYLWM0^=K/2^8PPa)HVL&7)4@=STJf<9FgZA.:E94
f?POfeCO1OY^FK<e#<g#fcI4V@J@DHN+bYLXLQ+@/4cUD<TKe5XLgK6cVEVIR;26
M.SZ0C8]0.gF=\H(HPCg\,0@O3N(2Z=#OR?g,BWRV7U(+WMHOT+8?Z;G];5-J/]c
/NU/1USVLGe+:X=YDS1@],BU=e75<]0J.4BJf\7_#BZg)NW61E_S^67O5[fNeD4<
D_YIf^[L6KI>/YL\_/HL5,Z6_86<AaKX8)B9.F)2Z2]\Ic]JH1=XDP)_eDS:)UPW
K]+TFb5P24&S6/LcL5A5&f#.HB)bY>D>&b[M_3gd9(YL7:<W20/1/3LDCQT#4D#S
W^5Af(J;QRB.cA9B?b2@Cfgg8=Y/:,I3E3PVFc_5,gXeR?S/3N]aRP6JK2F/0Ab/
Fc=9@e><5aP4)^JSE+^[0,DL=/Z2JD<&CJL1f:.d5RO90F?(^F^;E\dfUV(F_Kge
2SI?@1?BeDf,^9N,?/@8^B(6fA[LK+;?E_@XS.fc]Oc\gCUKKG;N9C&W6[)b\=I3
Y6;-4EPdcI+U@QHU1^3a709=QBE7(P[V>WeYR#JJga/7R;1g@AB]]X-c(>\I:f+;
RS3HfVCeVOTgD#D_MW3X29a0](L@^KQ0I9R)?<I[142BD_ed724&\Gc[@a@STc(;
PG&ab5f8],SgNAfAgA6)+RT#f_/IH_Z?d/&N]8/;W@afS&M[RO@S/-a[-@U/OJD=
7>cW)TX@FM^EP9fU&1?W[L:9[9:2:<=V-d4a(=EH?SE>eC-;EX-YPAXQ(^G2LUOT
T2eR+CEEW.L3=FKFDE6BX(_/K:UQB+Z#TFG00Z)^0IL(>GZ2KESE/^<FAMGR,6X#
QZ:2)0[b_B\-@>/gIFZZU<+FKf>C])WAa,M:0[M[;c#L2EgNIf@79bW/FHe]C1)I
+8M(3]VQ_>=_6I(OTF;V[>RW;>[eO>T1cAbF=XK(.GT)=[bEXJX[7J/\@dDA@QPV
<9]GY_aa_HAPbSS,5_Tdf@EJXQa/dB)1=#@=5&WMNMMJN;3HR<:/VHHSS4+9PFU,
&S]ABAa@8OU>d=<@@Ea[[&(QO)@83^43XO7.0E5]Lc4858d2I==6OXT1HTW4N[)4
U9(UHSAVV2+Sf).S)b5WY48BJLX-DXGP_D)Ia4GC@+b5gQB(4e\<M4CC:HR)eT;U
[KN>\)2<cXW://:_J#Qb_c;&/;.2-PN_^HTK#R_XeC&?Wc8ZI3^5>2DL[@d5P2P-
(BSAT^[8]P6cO)f5@Z.?3D]@J1;f/II_I5Ug-(#Ga3]CI5cC5RS0Ig1G[3aJ])-^
DAWL2^-GF;>0@SSWL^L<L,7dMIAJ8INUN)g=Ud?6/aR>Hb.(_\^6O9Z@ER&BVE4\
g=LdcN:WVQ@-GbB&DQ)\RI/VO<Y=..L9ec<:S?-UU[J>e]O9S<O>bMKO>EC#?c#H
TY\1+W)R,N?OMP(ZKKZ)F>9E:1IUTF5ZVS9gX2,&B8fB(L1R_g,<.&)8PCP/3D+d
dDD6=CSKJ<=LUSH=Y0>]4BW81UC&b-Q/f9d[Q3.BgE3+\;2R2TC6)S_JB-Ob#EaO
Y+B\^O9f<\AGPZ8,TdE6KE7^5AYU1g3P]TX.DHSHCg9)709c&@:E7-A)GV7.D&K1
:Oad9-Ide.,dM?>;bSb^O,b[\Rb^2.6W_QRg<I8]#PKCEE#PWGTZ>8,a,4\O-(M3
)0JLM2YE-c\)W;F>83c1CZY@OC_T5MIK@=G>-?38B)6C/.:.(4J@cYKQVYC41QM1
_cNbOJE_U,_E7]-^[\4Bb<eJQFcgEWVP#E;];[TK#4d@fNZ8UH3;CR)>gXM9@2H2
g=G3Z?PR)+TO-7>a7SE^\ZDA01U+,d=9R9)?OW>>HDY\W4QfI)8S#,]X^0D@V(8<
JHM6,F)e/F;O4D9SD+b=7XPT8K4]b6[A3<;2F\(39S#O+@8=44/4c8/bVCAPXPEB
OfN?TQ+EPMBC[?KHdU]P04TDYD(KfYSFJd\T^1PO>UPTF1GS<4ID-VII:97aB0eg
3<.fO,U]&621.Y]D]=,3NdfHA520@J-C48Q[3]<W0==@D+E-7_SEcf?BD_5Z5Z/S
FF[0.]0=24_/@AYDO@??0L#H+>38O>C2AO2.:9If>H/H;57(48[-Y7,8Y5/LD:1+
-R+e5ffVdYNe@/X?FTLEBJEWWOGE6VYc#?Z-;=K0.d#1+WNQ#?^QT[[R&bS_GQ\G
//g:>VHHZ8][Z8U-H)COFZBeQ^=>/QLI8-\TDY]\P+00WSY2?>^TWdA7A5:2C40A
4LGf]5LG,;ETJ#&[[#7BIcC-:0d)6RMgQ2.E=f=KG0ELEMG7dB&c346B/Oa;DcPD
g(1KZX5]G7<?3#@8gQRe<-UR\36SaeV=/Q@0[7:Ug5d@2Ke:.K@Q51)=>M9FTFV<
9G0GbQc.JL6U]GYI4+dcHa(L@P#]1E,,>YKZQe?G2TQ:Ed01DU_aLR)@WDN3H.GH
Y8&TdIWdHJHP85fT,H:O6gB4?\;@@8aGJ9.FUZ_NEID0H35(P<191+F<Q1I]1VCA
B?-TV_NN#QX\8N8V=_+[Z+7LcLP,BWEWWWM\^^(gBC5EM\99_T)_/H9H3f_[IP.8
<IS:Y[E=UHEc__+aJg97)cTFU(3+b@06WcOP&L)=Fb:O=_<1ULc_TcfM)?94D3,G
a^C]4cD:5cNd0RRJMPN&4:ZCIB?F:F#>W+[SMfO64.O<+-<=UJLa[6WOT<b.4S8\
L4Y+#(aI0?eL9]5BR3,Q5baW^DA[D8)cL&5g_0A.e@;1NNeB,Wf:/SHK1?_=b,HX
>fI)&MaaH6>H6]17\a\@DaZ.,8VTO?7.YXH\EeQ6[2^FBR#[&9AHb<;e6Y/I&S)6
CH<U]2>V>X8=;#YQV5>4R:629._D)8+TMfacF>N&9eeQ_:>1PFaJ/,Z07KH0@f+<
EQ0N5bX6;O8IVE@Q+a\R_:;O-UK,HNS=&14O,</bI.H;KKFEO3:G/M/YO58ZU^(f
AA59a:gTDGe>[Ze-WN3ZW?Fgf:D=gBS-Kf#f,+9c5YN?YD1BJ;W?Q-@C9XY/cYc2
U#4RL)H+<,&(R@b([H,cDH5BECZ[AU14QY&V#Q&3+-0A+QU@c9OUe>,gE_GCH&E=
BEcU+ZR-Sfg>W^gc3cSD^-FPE(ZXR+/gKg#D&<\=+),=VN9CJL7-4<-0OUS:b;<<
>6P6>0AH;W5ScRG6GE0UPe8g,GQS1WOW51&3G/(JANdCL8_M?b>9)31-H=Z=,:/C
;2/FT?dR[F\+W(a;5-/3@T[7a4AXDT+)f:8d(,4>\TXSV9aCUR;,KT^9b9<:,\fT
J]d9AaER\YO1/4]d^eZEUA)]N,/R>AbRCEDKJ?NWe^&_DC-F7CVI/Rf-cEKDaL69
ISZ4,Ue-N?Q#d3?-8,U=Y\)A5+Ce,cOO<E6^GTTDHg#[&c[,XH09;4Te/\26bGO7
5LM#dF#),a]I2K:^GcAg<TIVe,bWd8):@+A2K.D+.4EIEL2C&Y;,=3ENZ&U-DM7_
Fbc#Q(#:KH9J7R#9bd9LLI_QcI/N(A&PFACWRT4F)C8a,<=:=?M<E(Q>D\0,b3gK
:Uc.G/I=/7>=WVAX@W2SOA74b8-[(N4;g\;;\QHc-aTgX+C58\=J,;e^]UARdT:b
6>=Odb6Y:H?9G)WL?aE,1_J,M6=,93bV?V(+&Gf5((f??g46>EK\K(ET&:VXHd/:
I+6I3f8ePS1G33d9?8T7>7R+D3JZ>24W(NT^fP(Cc]>Q5JA47(1I85(>+;9NJ0Nf
72POBIdR_P7FRLH4-62e8fMTKGI[HGDMbR+3S>,#)KT??^72fL&Y&g-8KGFaLZOE
Ue0T#>Z^CS3d9Z-3=IU^I:bPW_^\V.R(9MDI]WI1#Mg<O?9^<QcfL?M/8S]2\B;D
D6.fW/e6Adb)G2JdgeGH]8ICdIZ]42/XIc@,OC0#)VL?I><HGZXgTD4?e^;5Kag6
E<>:4H9?;LTdD:EU+,2;I[ffA&0^M_aeXBfKFZ1L0.(?L)cb>fR4]E:Q?c+JI+).
0>N,dAefgKY\ea@?SBg-KcUK=(M6:,EUP+Q)2bU<Z6A30dS?92PT2ZIXEY)P]>Z,
5WP&2HASW9;>4FV8eXA?O&A8FK:VJL74-[bBf<.>&(YJ+Y2#P<GE0cS<A6>\/TE0
F??BR[X).]OX8D-N]J:TNQ&]A9#9X_QKW-(S6^dU6J(CSJG0fM.8J44g^]/]1BN<
F,+?6-<T\Ad,bfZUeH&VAZF-PEIRY:,I&)QD>\RM]7LTC^aLg7ON<M@8K>6U1Q(0
b8NO/@c&9DVT^3(PI2<0O1Y]..[fY3,S7UDf86<1G:3EKGEZKe,TY)cB=6RO[Z+.
\d)cM#DJ6:-P.:>cMcC-YGc#PZW)^0+HCS65a7&Ree=DTRGgX^\bH3GE6bGedFQ&
:Bg5DRHd6X4Vea.3QEB=11=5\I@5?W4^9<2<a6><VMT@.Y<I?1dfe+.AY:5F(cT9
S_CfIDc:4NcI-.P=75B_Q1<Ff>YA8:T5_-(M/5.c\dP;U=4Q([OH7V:#fN?@?4dM
I3(O^+)&5e];H(Ub<&TG:XN@Td<AHcOYZ#L8D-:PKW;MVR>&g.FC)DAM3>5GGdHB
WFb&FLB=L9O@Af6J>_;(Sgb@^YGE+DYI-4F0IVS6CNF,C@<Y1KJ,gPH=W-<g&SS0
K:_X;VEZEBd):=TJX2M5_QN=ZG7#Cc.F81YF_D5(_gV<1R3C)XgDS/HT](&@S6e4
c&PW9OH@0c9.eaRI>]CA#=<4J9UE??+a(J)U&bA@;L4IGWc_W6J0&W,A.(d;_,b,
7ED1OeacQV1&cg>ge>\fQ.4@ENO&0\<>dF_D)f_UAXC[UG4Raa+8FIKg_K4O)URb
[SZKY:.LB?ELDb>KHN5b0LPQg@ZS8S5+D:4UO&7;gL[L+3CUOSG4#Ad^2aPQOJCa
FDS,D4C0#+g_Z&#)[)g3]Yc+JU8bE@RS@R)f_M988-74T2E\LE&R0=Y-Bfbg.?(<
]MWb7;RO]4SIL)bdS]O&\TgCBUB;/==CQASf-c6#\G^QE;L1A?U-fDQPfZN.>\Q+
YU,6=fd)g<8\_7_5PP?CF\NGFS4=)O:Xa=DH+3>24]+2?78/#O=?WP7_<;fX+KYX
FG4DJRY]V?\N/f<,TENb(7T:6c6@=S;EZTU:g;5O0Z-S2/IH76N3S-)MY2<^0O4I
9MGU#V1B4[BVN@.5b8;R9WM9D=<Z[B:\>7W&(eO+8&G4,O[^^(PF7:MI;XZ_3[C[
P->]-defK8I8P(QCfdCKR\H0dEAbDT[]1)@)+H6=[&>.,IUAXH1:0V:HNaXeR#,[
EHAHM7T(ZJQU_UAV7V)(IBaI(@EB,6Z:DX2C>^=ZE(SE:M(e(@K6SF7@>2L.EK]-
XDMM1=QI:^)R44(UI3M#?5FWbUN;J3ZK3#5CMS+8/2K]GAIUM2XKeXd#/<I0G<#W
<5CSICN&V2D(-1;+G:@3eIeEfOcW8_dMLgV6G)>gM?PWF.fP;<NG:/)B/0)X+8YB
WK08#;?XZYEHPI-Y]8>#JHE#BPF<JDg_&[2,UD??A4Y.<.HVd+^7:WEE5/:_I)2(
e,#&EeO;VVgg0TG)Y.#22;V178:T9.\BVJG&5C:1S+23]1f^<KVeL?g1CG2J_>,)
TT3LU./0;>ccXH<FeZffAK\)GA&<g<N4I&eE#Q(+P\f3W?<TM3^TW&>e3NIZP?@9
-Q6_.VF>.@3B6O_HV]Z+/DV7RY3.:CLgXeKZK&I0&+U7\P,R0Ra2+M>7c9>+D-,\
\VQd\Oa.a&LfG6JPFCUHY\-GN9M6CBb<A>OZ^RG[UeaVCH;e=K,KNI)K_>1SDHVg
G.EfUcABa6X2ICf.PCVK9f@DD(I8CZ?K:]HJgFT?D-WHNIgeRaM7\I9b>&HNd.cZ
S\GeUfL7X0e+:HM4,(8eIB,d5]#AI8,[\U1fH^T9c>IbVX^]4X>Qd,OO[M>/,K@W
CZYD]8YQ+WQcbP-PMH[g46<BHQ]@715OOTF+X]@#.?)@5C+d:,90Be1NX.KKfP(T
4(ED\76#60MJULQ]QNSc/M1Y@]1dg_U+cT>Hc^PD3I#,aPW0+9g8gYfQI\f+_PBT
^2,edXFXPf^Ocaa68^N3VbH^7dD5:3H,4PIB2Q/VfX,=<7)=TURHaG#(:>W#7Z@N
&J(Y<b3=3:6<833adYd#,7ES@DZ179:3F/=P>N)bK0^E;BNV#HI.dIM6W5O=E/4T
.BT1R-5[cf2,,e58U?:WFQO.eHG41@S5K?3[8R49WMC^ZTX3DH]=Ag4fIG]a:BM=
O9XJZ?BC+BCM<Z\c3E85^^[b4B_9VE7E?KA,GDVNTbDG+BM]SC5b_^G4^Ma>/W;0
7@b7X?&7;:4<baSBe:H^(>P=M+?[\0]+(g67.\53B1M+GL72+]\bBd+R@U1R#U0M
2XC4NZPE9XXTdY+9(NPW]FV<2S+^RW>NAS75/SLHSCfBW+)dR]c.Od.Rdea>#3f0
/+7QH^PPHM;5?6CYSMY;-GT,B;ERG)K(8e0#&H3Lg4&Y\I/?;:6F=QT]d7PZNR\[
0NCG@_6TAM2eCN7L7=Teg]TOPFa/Q&5NHe,U[Ef+S&PYf0(+>K1#)?aZ(W5:10=C
<A@E.=c(R;?@SZYLJ)2L4A<NL@(G@<7#DSc1BJS@BTD8H4e0A\?//cg2M<53f\5\
R?YPb8\@7D0P#g.#R\VXg#cOO<QTZ[F[D=0DJGZJ(/DDJa&Sg8FF:MB378+?7<)[
;)>=e:9<KVc&-F>EY.+>Z?1[>LaM)(::?267QWA4-[Q<.T?A@@GKc[G^HAT^0A^@
<bE>g#^BLAPI/M,:W:dBFf6,VC8Cfb]+>T]=T#^AHg(;K:aWMR5;>\QTVA8;:H[,
,]>0e7&W+H6T&;RB,O\1E2CMV8Uf\J0:C(R-QJ;69.,(ba<;8YcHHA0&UTN><Sb#
d/)D;Z></Ha[Q0IH@5baPU/N,A33[]])f,L&L<AG3.F=O:33[JY>7ZMKd;\YT3I[
#<X.4(Yb_?A>\V8S9ga)>X#T<NJDG-K335d8gBE?B9ecR;]]1=M3ZcN9ffM)7Q4<
UY2=.&H:0eN@Z1(0.&MK&A#EG_V3D/C-J1@fIJO^\eS;[+8DOCbIPag+bB(E+NI1
46.1=J2)/)WQ<63^b9^)BUOUR&0T<?#?7<W?7\=]+Q4dOXUUO;c[[<MVN[,>C/.,
.Z4B_?F[0f..?:MUWg,&X)0=3X4bHG1IUf0F]DOI=YMUVB)WV((1V:/JS=P&E5=_
aUeQ;2R>AdH5HW&..T3-e-22S1,b^?Y+R4@[Ob_.N<I_M:1K9fK5B4PPS_MY.2Z#
NHQ7Q1eP&9(1KRZ9@)EWC6?.]C4caNN86.[@YB3UD2[K51HE:5f[[O&]([6\0)VM
B<UA\@G0;ZY]T,=.?52BN4-CG[@E915BgfZ4A>TN0LEbe[ZVDN8SV14E3aFIIa)3
f:F4Ae:Y1J^?&CS[6W:21SXSe2ZG#DAX&[SNNYH?a#WNX,8U^;<[V,PG?</e:/L[
Eb_cK3[#;Y?I(_1LM#X(+<(\b_b9M@JJH<+;(fVD]J><eW.O6DTX?2/),:L#3+H?
0S-KH9C8Z(SR6-:_K6+d.P_V7#P?5Q5?+6Yd#N<>d:LL(7c#=\<gA9B4IJa(BX1_
,1-;0:8EK@f_-3N0PIG/ea]8AMW.-;/O[Xgd^P3R>LC&>aC:KgU_49HK;&BN:\RY
I5MXX.FK7S0ac1=YEDPFK>Q4WF+e+],(@5dI&P)V3?2;U50?UMS6M>R02cdEBAU+
,R+?&Y^KAQUV+EbSHY4:Y4]C<D>U:_<TVRL+?)T_LA#50:A@>V0X&LMXCCGNMf6]
YRW>U:eYYB7J6DM,,+?POEIJ&E/,>Mc3FS4Y/e&Ea#4[;[5#gX^gE>>3A67[d0GQ
E0bbS+8;MQVYV\C-=_^G3&.X;W0=Y?(9.V5+S#O^C/Ub_IOLA^N/LG1^HZ5bH#B6
cJBb9\<QXCS._^K/#99&1Z0\E(D?ffP@bfb+B=NB_d=9=(HKfgF1?#faYE+Ce&E8
2OJ8f2I0B;YLJ>cgSMB5\a4&)^PbY621C2BP?Z9&?19a)TBE.ZeH\Z_ZPNcI<=^2
PH0.GMIV/OBaMTG.g475;gZbO@O#S@J?56(=7QZ]YZNE4aI_9Pc>R<UZ:U(F4.F[
89(IU;;HTT57M->V)=S:>bR&+<b)Qg+Kd&b.GQ7+GEQ559][)P[NKgQ-DR,C3Rg1
MHeTK3eVA,g7(N&XgY7=AION-;C0K+O9Qg8b3]1f+1d.HQE5=db<Iab,W+29ZgfB
P.Ab,2HS5Tc+P;XLSbf^QU3LN6C8(G.@&:TH601IJdF.YYU#Ag8H?.3_@D38,D6Z
2(;[La?f20Pf<2eAc]dC<L@Gc)8D2+#F]-K5T=FH,F)DS9(]@&E2eJA]K5\-K(:+
U@Vd8Q<Z.@)dCKHgG[BP26.PEW]FE\P873X:=/bKaOI32/J1Db;Ya9N_Za2@K+=+
QU0I-YE6@TW1V#]OIc.;(T>2Gaa+EM]eSD<>5bC.O?a>-3GR/O6g^^:egB;g]EZ5
VG+a0Cc-?FUP_AXJR^+SIS4-:Q3EO:?Va^&L[EBg-T?D-=>I-;+28WOFFYWG0NW1
]<M>77PgH0T-&+NXCDb34Df#fN1b4@V6bJPaBeROJ&2M,R?@6:Q29WH?afPf^Ygf
Sc[5-3QC+a4-^ER/2/G+f=(B.N91.eR)BV#9U0;31K1=4^E^]bV\OGS9NZ>JG@DX
3fRN6+B/Kg?f0Ea]VQa@;#@L_aIaD@)#T45>A<e<W>.2ecWEf#85#D_S=N\7^=/4
1/c?cO&4DK7g=c=L8_XcgN#7Ig0^6#JA&[]UbNX5ZPW;:7EZ?8>c]IE&Ee&UdfD<
#PM^30:eC+.-:O;78(KOf:I=N^NRf;QS<KPg)]W._dL^@FR9UOYbB)-A&J>Y-^S>
;E..5bQ^^K0UFX]\g=@JE<Y6Bb#ZC3H)MD,[HeH8@T^R;cPPN97aB#L.:<fQ6W,]
32a\VI6/8-O+&?A-2)F14e2X1Me3ab,OD@,BV/O?D6VD-H247UYc<R2\KGL(#6B:
Aa/NA)Q+R058#1#WK_;<feROafbKGeE@,K/77cT3ILX8L-LU:01EN.HF8&M<CJ.X
c7G^]0#YN5];8.2:\.9@]:/UfLU(,=GfVRK]4/<Z#)OKPPLTW>9#EXJI6I0Zf]@:
.EKF(D.Y<J]3_AZB+8La_H3@LF)1DCRa21(e2fdV/=2S9G\I8E650_K&E./^Lg^.
CeW0DI7fE24]+aU8+R]3bA:=#2-^ST\Od=#5)-aLB9e4@P#:^F-6_4KeH7a^@,<:
&XO#7[VbQ).@EfEM6DA[f+#N+7-O>,J6RCU[3E#O&8eM1B8b1[P7^44Q^@fPDY3d
cWT@C-[492H61@A:80e#:3,B[e:QM]UD_.=#ffJK\-Z>,WAXLR?A#7DH&7>HF+e@
7A6-5@_Rg:WL_C^,_S#]FeLE/9EO\dBaLN5I+[@Y0N;+9g&/)MF3,WGO,?@86Xbd
^HcL_Ia=?4eSNbg)JM04BVI6b(EgMPR4XVe@OVXU(T^Hg7-Q#73NP3f^MY(F/dYC
/@-^[4;#HG_-W&45H2<Q,D9d2V5&aX>eQ>9f14GX;cfZP<QKJCCVD9@7d&4^SC0@
:,ZOaI)&D&J0YZaD-BAL(;S3Q2L-XZ)UcWN8G<dB-LGGT8b@I4fIG4dCJH)-1V[6
IAEN=\,.Q10HV1d\F4[;Y=a(OT,0;U.+;>B8/LX,9O8\1?_;)G32P/g+44&__<cS
gZ/5]7cfb@5)6H1C1;B_A,eeR:])FWfcE>b1d5,1F)-(<)EW\^b?^4&e,-/P+_HZ
&B8)^H>Y4Y3Bf2]Af>#EaN^#eZ;^cQ1[QQ@ZaM<BOI]]FU1JA7>a2O0R#5MJT(M2
#HCS1f+?;849aJ?P0Mb<#335\e.-GZ])8]/PPX\X&dXc8aV?f&3S((_RSM</Ide[
WE^8b>Y6&13=GX=4^LL7VWbXQ_>f&82FXc:cf5Z6/&#W/[92W[d/7C:UG0W(LC+L
X^3?#I=9\2M>@g;NTVF(,NI65SM\DZW:O;#J&6gTB#0S+_a4;I,,feJLJJ=M3;^M
ZN1&bU6Q_0;.CW20SL2:.XS)H<]KN.L(B@L.XFO.[gDf=<#[)B/W5f7fF+085E[[
XcD+K)aY&QBdSDYI-\]&f3#C41cQJCC37e?<Y^]6ee,@,-3FWY([g=6T]\]JI&FU
9=)2#A>+gTO^9Z8]&D(gDA@K8<E-1P8H9\90S\@A:_\b1R9cR5APNb]Gae/2DQ&a
bTL2&>F/G\W)Sff;PPM\-g2ETLF+UC:7GW2cMQgb/I6_L2e60F?_^aV\;P:e1PAC
b4T]49U2LdS3^A0=QI[\P>1/<:eVH83:EH7<&)#A.F3J(bVecS?WG?EIJ&E\XP.?
AR7[4.F6:#27UK.=G_bdZc)F8bY](V_^6CVD7\f[JZV2;.@a9X8C91QKM+eTK-.0
eC;+I4M8PfYLJ__,c;VQ]eA2]F@YIPg@)]V8BGI,Y0b\M36.@[X3Q#fS,;HX]&GC
C?Y6^bQ\6NS3/=NFYXN>A_)@:]2_;g@S2L]\L4DNK1)^f\I9IXBD3#8S?)Y=CW72
IA6+20e_Rga9gOYKG>=15_WI>PA7F?RC#MTaK5cC(V.d.TKX>L]82RP:X=0PA]AG
dbV8]6[OdO+PI@EEW1\4W2K?8_&Td8aXLgc1CeQ0Z<B-_FY4DRB@>NF37?PUY(b7
\,;QI#9F1aMZI#^gf1../QF9ZfFL,E5c2S8f]?Q\@aFF\K4]e-0K(THAKP-.CIR\
<2>P^T_SIBK@;ZafIfeHMAJ15RIFg]?6)CZ)Z:Db//VD=SJ/D[dH5;N7db>L\9&9
e,;?CHTeSGHXAA:HA7S6(8G)DJIbX1AfXQTa7PPEHI:.[YSfJW@61L_&L1+3/7;8
E_6_WbFD.R]VX<RAN#Z#eOdG8G(&W)I0gUdT,+1\J_Fb?dE^@482e[P#N@;MA#8#
9.3bgK5C=GYUAc^<HV58&D)ZJF3XBPXAL1;UJ\7[X?R-@cI344G^Mc3W+=Q8[D7S
d/FP)6AF1)NaA.bI#&a0K2)8^b@g\fcNadUVbaaTFOG9I=O47.\31<VV4YL\6aV^
_V);Kd+/7?=W3DQ_e#6-]6VMS6POAJXUFL\4-/(6g622KEe3D0a,(:&@_\eZUS+S
/1Mcd\(6Y(>I0?7&E7.(U(gQF0DEaCTd4?7M:CX\,)7@7JgfI]FXe8I/A1dQ&^&>
DGTH_XgT\I+P7/3O::LHeC)aE]Je4cgPZCBCQXEe6g@01]XTcbW>b93DD]BDE@@f
f5ce_KFA4eH2T#bV(M(7M[I30NgO+#\6&=Sb^?&KKN[T7J86>gEP4E#-0;-3\4=0
+QaKN8af\@V@Y6ANX[S-=WJPKJ<cP0[_#[fNV;N.Z2PcU4aA-F_+VWd)GIeOZFK#
W@?M=<^<RgdC_X/)Rbe0;E<\_9EPN3?>96Ob>VK;V.H@#ZNGPK4b)1EKV/Zb.YDG
SY_CA1VY1COda5HA<#;E0;?.F/-5LD_=.[=e.g<ZKWQPW71fD>94FCK&(=.0ZE:T
7gML;N;;+]SP,>Y,#9EXL.e>d@8?;I[Gc9(@eE<9(c5@T7)7)\[I8H6M3UKT7g^Y
^;WfP?B?ggc^YF63T)Sd==4(4e.Z@3PgWCSVeYT5MTU7J:[A;H4WP3:QG5A]Ba4F
dK7Q-;1XX:IGF8/]G\VTV&A_.(eW?2fQN0)eDaEMXAG\cUW[U(W\;>.M-@XK.gD,
I(]b>7[-(2H9_>SW5@VVO+]F(#/VUY2/;HR_Q5G#/:VNHgUD;[C<Pd(f<b^7(GZM
7MKULH,?72BXS2[3)8W.+(0RaB&[]8_^d&1UWd3WH)dP@D[ga-#d,].cH?GO:SWJ
XaXJgB,T>?23M+Tg6#5K.NcWdK=[3W]S#VOSV6DA=C[G::LPb_^@@Rfa/I=+4Bg:
V9,41X2SG/e(XT@SY,8JRG<1=@3.W[X=9C\@J+;^WN8S(7T&(+@3,&U5(:J>R4/>
0>.^58)&54aEL<LA)@IFXa]&I=J7?Jc6.edGDY7@S169@B@dIc4#173QX7baA([J
AC(YM?3,YHDX])G8D[D.,eHP?7WRdXVT.ODd^BaNNKAaO6b>a-<;Y([F+B/GL)DF
\4UY[M_gC,Q]\b_E=c\+7#LR2R5a8[ed#;91<Kf8NZJ9\@(L,PZG#&W\(6CH.+X3
V+12g<NQ,KI@C@(WEAP&Cb3IF(^?)-d>-,LO3QAJe8QLLNI9O7;;4Z?YDB])a(N9
R2)QKJe-EW_J38I)Nd)K@ZW\D71f.GI/;?5,AdM:__X_E9A4WgS:.=.=gJ(9egVZ
?SeHJ<OHF8_5DP)aJM73>T)CCV-RP,SYb/D/2@]RY<U]TM661aLZUU])?cCL4Kg[
ZVW>XX+EX?]^5N64c_eJa-EbM?=?@\XC6F1M5;:QF#/b.BFe19AAa5HRQ7BbR_87
J<S9RH_]gD/N7[<c[gIFc8]LX5(03TUIW\[^3b>=[=7^@2:.Q>V^JGN)ZcI^JID6
_OacU+(TI1+\]b\)>T,0aC-^FB=;BR^BPKRL9M8Ec1@?=2=TRV9fE(3U;g=gR2)f
MAe=(>Z_9,^8O[e1MYP7W],e4[A-M)^;e)79&UE1g9T.Z9E0\9eSMVJ1&^S4DU<9
O.#1N9H1a3N/+^PA2K:0\;H^#,/^e1(\9ZT9(K9T1NNY]<UV8:@F&5^;Nf&2>8Z?
cRRLZFW)V[<6,6,I2&W(a<D4JO=]##d^4Q13a7XUWXD,f.=DfF5_gRZO&#(SG9B(
3S[PeHE11A;J^/[W^#-+8W.d\6P3K9\-N@NeNN\KgXQ2@c0\Q8[TSaVO-abQeH(5
/-CG2NacQO:PUaaGSLC\VOXX>\gb3[5COG\7K8_^2LHUJ_\94W:]ZI94dTTf<T:)
QZ:7@T6=3T+USLaE\2KMcOaYETAN@855UJ5&6[D)(=11VfF0E:JK3:Z?DaAD.#<-
52gb8@_,C]K[eBH3W8PVPF;=IM=7#Me/^b5KY&^JC3I_[WSLU^-O-P6RZMe@9)QC
fO<RDRIMRfG^5CG]1<Cb+UaII);532b>8H<X/FFg+TT2eVcf7<4]YA-c^#P#_R=;
eY;BUb:(G):a\6=f13;VI<[(:KLJF^6)#;TaJGQD?_S=K#eCHGV?HGd,)52G(/_E
V:QaA3^O[CGgVKg@>HBMd6fQS[5K>d?FM0T.-(8.(0&@+HA?/LZU,TO]@-K1TbZ_
Y;0X4?N,0IHe>/N/>WOc;^RXgUcS>NPY[Y8:6W:E-V3X5bX?V@;\J;77fb>THc>+
Ybf(OHOU#c22,O+?0>@O?71J(P6I8ZA6KFb1QRLGc2NHWN9V-0@+)F-&O2TT?b8=
E]JLef@WS6A_@<FZ,_BI9KHJ)>-#Da1O&5ag>PUcX?)#3_/_EF:1X@YE8IOW.H4J
b9)g#)aVEE8)?KZ-SPZ8:eAbF]CJA2YZ)B5?d=)=Qe(;)f[6X?6YD5=R?RCW@&]5
2]Rc^;VPVZ.2D9MH_)828I_W:R,2e=cN^gd;+,PM0)cZef,:H5@G@RdfTJI\e4Kg
Z<,U&H]_dWgB&YW0T7,F9SL8Tf8c/JKPX#UQG)8>(:THMNN#^L3:QMU-_(3Pe&0]
(+8DI+2JcJ44NS.eE_9A#EA#MDH/gN46K&8Ga5@QZc>V,NT?OJ0.G#0^]?]2Qe(1
L1@?D,cId;W,d#cT.6P4Y[6bI&JOag35?0FG\7X_(IMBIW/@?gP>Y7W8]S0(FH(d
)FSPbbH<U2,(YJBc6CCOJe;DYQf9+969U\.SP-JV.;.\#[4-/5P.[7.9VgV=J-0U
4GaRIb))5,f[\f0#[2I7A83Kf-I4KP5IZ(V#V:H[QKI0f;,W_)NXG790d3S();XZ
gG&e>JL/1Na/#5G[dgD8&a^Z3B87>P\S)JVXb.\/A_a7gE>/OX[?L)=U0RFH(e8g
4d11;&76&N<(Y^@_D^74fUQVd&O15S=YRO2=I/OR4#O)YI@\A\1.cM=0DC?Q#7XS
DIW6W&?JATQ-CZ996^[N2WJA6V/Ce?Kg@P<(?[GZcRNS]])<,UDV::8A:/?7DXVL
7LEYT?-/\aKL@@[gKRe-^G>\N^+8@_8#,a:JW3aPN1?gcCJ4P_7TdMW0MP-?Ud(/
52O4Z0R#_6I?Xa.6MOPY1HI)9WeC5=9LG;T9#=AN9.O;VUPd1.c>Z06H9cFe6OP3
d?OEW3IAT^?P?^@\B^B=<Q8fVLZLegMSfU[)V-.TB66WGJ.E@\Yd(7&_>N:7&OFf
;ZQZ)M59C^#Q-+8#?\W\C2PABXEM_+#8EF=6B8_MOPUW>S+:W8Y&9UJ?CA5A24d4
Na5BgbRSUFd-7.V7[PAUQSR@8\Zba+D4S1JaA@@7LQ?;31agY+#K7JK6QMJ-.&SY
Zd;.(S)#0[-Ze_:F\YfAH<UZGXc45Be.9VLE,>c;WO/1SVO>bD>GbGE;/N?dP+:d
A.fDdUgdGXg>-X,5<LETPSca:/=,LPMEGYU_X(R#I7?X+bEKRN@UR_LOQ^P&]@L&
^a^5UVKBQ9-aGL6=EUO:T/aL9MC#f2US>BFg1D^5C0Qd?Xb_2<S]=d;5D/&GKXcM
S,G21HT8g2&]&Q_]aR0;3VU-Gg2.9:gTK40f?aJ@_8DA]>Ig,ZHQDE#/5I.MX]+/
--HfeXU&3/<&EMQP5G0b+-A+R5ZeR53F:EC>=9V/,KY?#D+KS\J?E\/1-.I_-4R2
G/M]DPEbKS[#779+)LWX(3T1c[5OT:6.X_,X0WRG&+@.U?,Vc8?,Ja1RgFL,\SO[
][7_EO=N^<\0_;AJIbEX5@G,T]@&J\&;9U/WBC]\R(GHc,H#Ve/#-O;<g0ECL7/P
]EZ5=Kf1d&eK+.M-ee7Cf[Kb7<a.(bE:@SQ3W0,WE245312.^?M1HeW2V_CUTHbZ
Z/^b#KM?RT;:eb,EO-2ZQ<^aC(bcV]f^YQB^&D6Oa]+0206Z4,A.PWO75+)gPW#]
[G\HHX2J;6-?.)7B;?,ddU979_2-3@@K(^AP;CWC^Ja2&5;FYeDU?GV-_V0=G+X=
910.>D;TEL=FN(X]\TB1WJ63=X@LEQ.U38IT:@d\:d4EfUNa+7UB4]U9^dUHB\K>
SBHEN6L/+GQ:)U9NEQ\KON<c9]NH.cKfQ4K15\3]@>?IOTg0J8KD>MGa.cU.G^[G
3bdRVX_W+@aU:\L3IB-U=NC<AB-PC]B0I[=(Hf[[S1-/>\cd(KQ#/MG-V[VH,;O(
U#RJ>dO4@HO1>;WaLPg,d:F_Md9C(3U2-DX<aR8?c5K.Q<XeUe\:;\8a?Cc@P?)(
>;:_.Y<,[RE=2]D29/-&Y-//_ZWgOY<27Y9;A-#3?cCbE?+7+^PQFe_TK3BG7c<F
d2U^5(W7_d>+H/A6G&(]Wf-]^SWZL<:\[[B\-M]8RNA1HCZ+[[(1\/@;Yg]X37#Z
Ycd]Ee=[1J_8C0?0R)9#?CW&33c]]M@GNdae6-X@GAc3F=CK52bZ<cC5S2OC8C9c
,_.-^+d+#FZ.,7H>F?f([]BWXV#:.9,7b6A.)g5?aXO3.)JVfYTOc/[30E8(TJM_
d3&b<U7=fII]SQ9PPD,GNeO1]0IK>7D#5UDVZ^c,?SKFPBc->3aW>eU#K0##40@+
dNUa#BW07#58L2[=K&/E^JQM?R<R_UTU]:b&7Eg2\F+HCF-&^3?RggSN;fSU14b:
<a:=IM+CaG5<2+.R@@.X)9K7F6IQ+1A/f6AAOME8M]fX+]H7BafNEb@X3OBEDN8\
X8A>bR_g1\/U1ZO/P\E?;<L,78QA_X<8QO7TS)K&fWR5BIgbL0+d>2[\fF5KGR]<
AC#V9+-32&N]3<)I?D_d;,R0HGCO_<HIX]YY/5@eM^50H,CE.24XIPfFC[MY[Q&Y
3=QAD@Ncaf57\[5D5,(LCYaR4DbBTHT(1:1b)B6:Oe&KR7(2LG:2F(c6:O9O7F2g
H:Q-/b_S+VfW#(4BU[,,Na72:b[)1-DD[U8G@YKVUHI<3fb[:Q&@d.MF6979-7&Z
(Jf8(+G^5@d.NMX=1V.UI-88TbJ-cU6Pa6)V)SL?=7/1];D58G<+dEI_D5g67e2@
PV.;FCH].SZ54?3cJR/aYL/F4,2gX7U:&QEKLaT9UcYZ[IVTMSWWe5>KE+Ib9NVN
_5BZ(=C-]e@BPB\\47M5LZ:?C(fBP.60VI^=4,BQNK::WQ<Pb]H^.NF4e((K,SFf
YAY+OB5e0A(XH^EBdVLVM1-6Df(-&[4JdWC33[Z83EgCbXIM.Qf^_H1N#S]6&f=Z
P,?QfDX.7XKMV>5-\eFS_[Sf(157#6\B,f\QS^Y7R^L0a7X7,Y\<J,67f#RWJ2/)
=eT8Z#@[b#W04cCf/],b6Cc^dI\c+fcd9d1:S8:YE8QP[<+\@\WJM\8_^e/[.S)E
\,.TG])OGZ=A]T7TYB1DR2L^TXF(4Oe@D)7EIU=3)+GRIWU#+]YF]Z-e6.LGgSP(
3UD[Ud94R-b32<^(,E);24IWGEP3S:cI-]Cb-:[XR4@</XX,YJ^=N5;=;9KXg[0#
>H3[(1X-@U+^T4e4=CBPNTI\fF_aEQ3>MV.Ca(RG6gL?8<HME=L_M<AX.MaD#@#d
S=Y8KOG4)U7CMOR..>9eHf8EN_E&@TBg^g0bJ[H-M#RB5eD<PIBF7?eb=FGY:,AL
9Lb&NU,[Y+0\=>aPG\\N9MGfGN>K5>WQ6bF_1:.\(]BJ<M#AGJ7#GGB#LTU;gK)<
+g)dD#<PM05267e@faT:6fR<UG.2fMTUEe)dcAY>Z@C##/a30-1J[[P:]H>PFLK4
fT4RTd#gIRJdLfWP3TJ<F4I^8S/1eCbNfbSI]O+=]RT;a5)/_[]Te&ca)5D/PR_C
13]9^?:7Z]A7=_0dH5,OXDWUc><(NSXFMFZ_M9>2c1B,&e>Eb;UfLT2J6JIC&>I4
Q9e2J,&^:aI_f1IP5=DX3Qa)QbP3]./U8/#48CIQ#H1L(V42cT)Jg4BBc];@7e4R
C&9DOY?3ECFL&?CR\+fWGF2O=b<]ReL#e-U-[:.E\ae[UeTf16T@07[aX50TPPJ(
0.V9HJaE82]+edP>PW9]75IQYL[87V;BC&aF;8;S/2Ta+,D-H;JWe,FPK/cSIa75
F6FH.;HX&(=bCgdS1,R).A()L.LUX>Q:4-+eV.62A1LP9MW+IJ>.GI?@(<4\V..c
cT9GQ4dV]EVOGa,I2.VUOe;\BI8NEd7a=DCIG#1GI3]3.+b+?V2D2DEA^6]c;W-5
Wc^A#8PTB>>e2H<YS1]I-HEYc9R>6I=22<(db:A=<R9MORVRL1;__=3G&N:eI6C9
agd&,(d/\ENHN_HD2Mg[BA8>CH];S0T>VaaJ0RQ;.9<+1f=<FM:S,3=<4AAd3K;^
4\bEQ#+F850+R+83^?)1G[20&0bQ8D[>8g0@Q>3O<FJ_5_;=e0QSg3K0fN+2TYXP
7aQ-G;T/2_F(;#e),BfH53]G/CE6f5#AY9]9XNFSD0:f.&F@R5<=ZEF1F94bTZ<(
(XPg0YD])1:A&-ZZ(KZ@eV4gA;&DS1bI885/K?U<HQBcR.U#:3Lcb1O<UQ9O^2+9
WQ)fTT+1YHebb6P1\7MTKJ1@&JA_WRU?K(#,]M0c?2c]bN)\M55_W<Q@7g\PP@8C
+@W1SYD_aJ/RFd59#eE6TQ+D-[bZBTcce;_L<JR#TR6/&,[:A1;3-28<)I_Jbca7
)P6d=R;NYKd66O.a^J]:49Q,-+/W,^H@X])UX(D8=(=eQ;SRJdMc)SU)<<IY5b/e
CJ[Z_31U,A<Mb)KQ:?gM-:B/?+-[^<0\+F3H-1;H?:cU5MBf1+VM^S7AF1JL/D.;
7^_ODJ2DQ]Z@/a.:-Z;db9S&REFEbP&;@]EIC)HIaec#=4+8beCaL+UQ+645C9cG
^5#<6eR4+Z2;La(c:MH1acJ[=^-PL#Pb(..KIfc@Jf\56cOXae+70MH>O5I4.IQP
;3:b)WXEE8;cQP/>[MYP==E;KaKc-6L0g)DJLQ?M0I[(K9)>-BYKc,SM<P/2,OXL
[cEe#6^M2]MJKHMGA2DXbO&5.PHECK3K+R8SOY(2RW[d&SM5SD/^(.]IWD#)[DKd
#UFE#g9^:R.MT.<_=T(PZe[(<\)?J3Y<JWEJQg#8gZ1^(6_67F_KePS)CWMG@dK9
=Q\2R2EcAEZBJ-J8H>IGe3D4K/4Ud1+#M<L/OgZ/f6eJRMR3.gHG<-=^K/\fX^03
:..(aO-4[)3C:QH6K7[UD,I&R@QD+\]Z-cUVO<S^=^T@bNgM(ae:#\cP]--7GJC7
(EfU.;bY=+7L]5611MbgNO>XS2V(Q^a/&eC1]K[5cJ[]A]?H\UIP)7\Kc2L(5HW:
^=@KTfY.917G9C8M=CJ]@A><K>]?=b\&U<<I,YJZga+O#d+(B:G]FKSJ3c<+APUT
(KO@J_I>XQb+aOE)#,?SIR6.ge;\A5]VMA5ODTF5A(.L45<#:ZZL?eT1V@XQfKeI
_#:WNS+;K4BT/@5.U&RH#fT\J[9[_IQc\X);77:VSM+TT1MR=3#_FG2<62\G6@]3
Uf:VW26VJSX(Q8f3)f&HW/(9@\3:-XN9:bZIB8AC4cXG8Ge#\22A+B-bY]_9^/&g
B,Y^RRAdNW<dN@f7e6T=?[=D8HgMR:E\cC:HQPXADgPM@^VV8RSY/,K1L:LD@.X2
CFQ_QcJD#260Bd;eV+;6&KWPASP5@[f1/15:6G?RHCTU:1LM>g./3IPbg&b98#3T
bT954<0[eRLLa.8a<M^#H(G[X5OSY:Egg\V-V71S)D?Q.RcPNDLD?=/5T83IORK0
?S;f;?11I=eD]9d0f+?F@MHX>@\GEPad(@eQHIfSgU:BUWPV46^V7@2[4/f:K0+0
T&N+d5&9#<\&=)cL72ZA)cKR\fA5F65S&EU.R)D9d?C-TGEXa\d,^gP&=I:NaQRI
_[]^.-+TQMSK:=b[>KM?173RX-#ZI9FD=P,[D42EG4gBC)?F^[._=\((PGE)3PO8
&TG0VgT?]S[OP7cZC8gVBH3=Fa7db_^XPfVI,^OY<[b+]RIa=5EVJ(7PaW>3,T3W
&K_K;_W#-=UU5ZG&b+V]G/?:f3VT5bR;/24S[a&I:0.:YZE@2R)?9Ff0]^6R-988
_FYJ7:GBNTLUB2#f0@LM1#H;L;La4C+H#.f1#GeE-GJ/c?I^9fg&?;LDef_//<f;
@4M,-cg^E/<I:5LFZH+F?61QA#+CdP8:=WL1F;H\H^E,^fK^KMe7TDE6,XeQL5\R
ZF(;]CKK8R^P^07]Ue\2T#J-;C7L;CI5WXE[&6D05_>XXX_+^S)eD3@EP)JK2/M(
e)&)]2>dcA8fQOJ8QY^6,.>8H6-UC(;>H99,]6bS&@d_M4IRgHND/TGC:bba:7MI
cRbKdF[5K(fN+S>B9@5:eNL5#JW;G02BT>]XMcf?[a)T__ST?>.L)/HT6T?.gX/Y
9QLd0P<LMMbKBA\AMY5@6UI-g[Y8L\bXD8gO/K--ON-R#0JCGZ-d5a&:4VX#^<C)
HQ)G8HO))CWIF\ZMKJSR&GGV/P@YTNaGWPR&3>VVBP7]MYPQ@.SII/LYY.M]W>4-
2NOFXON(<2-=Df\T6ZXY_f&<c0Q4APe2J>96]=24IGL):)Nfd\0^8KPC4+BJH^DL
Ca=H3f/OI/;[D&RFeRF>0LQ:QQK>e^#F60:.aY.]1,)aGF>SWE>:8Ia5F3+gD,@]
E7)#_M[Oc#Fb1?;8&b665=\@[YY_]LY7Z?HVaM7cRfMcRAeL-_[G+[Y\Z>#0C&&9
QY@W.JU_S39(A1>YHKIdcG8L<6-5\YafE9KPZD[;_1NE_SN,dIM<3gR,X(U-f,#^
JHP:^+\IS\=8G:(g(6UD\Dg[ACPGccF36AD4J;S(@B8.AO+5aOf=b34C6FN)X)QY
:<cfS81&b3+g2-FNV1:CW44Y:9NL^)TEXcLP3C:I?(b?,Jc&S],)_N?\&(PV^-5(
TV[S]\Sc27O1Nf_#Z=/[Pd2KWF/#dFQ;AN11<])#XUR94=c&DL_-MFF93AHED)?O
S)#f3:X.WIWFH6PV:a\@\H/C,M)A1STBV=ea3EO+GYY)+=)EYaZXSV?,=-_<>L^\
TY:R53M2X-=THFBS<+H:),@SR<1F@5:@,EQ-3Pgbe@];CgP_N28+-f+#\_9fC?LU
Sc=4EMVT3CNgB8Y3U434D9;e8UA]/-(K(6XAbbUg+:(<OO=^BUWR;@SQY:.\\P^,
8Y7.+6.5&Q6^T-=3TUQ5D^E,([_N)Re]15fFGU4ALLZeDMF]_W^NBH[E,eXU86GT
:6[ZUK#7?3\47V&Wa_91FBX>1WQCd1H.DM34/XU,#PEA4?abgQ:TV4)85ZWX6FU(
0U4a]SH68FPL@[;&M1Nbd6,g])HQOLHAM)].cce646@#M@8FDSIaV6/:[6?RH@gL
b6[P0FM4]467V2T:-(+b^<<ZUWR7+SN(#N7bbV^Dd\3#N@48,9LgE)Dfa;1eAJ2Q
5X&[RTc.ZfD3;/;WZ7(+[1@aIQQ#gKLNW(\^8&9f_]J2)FA?TZ()dfWU5Pa8F<3E
@&329LSFFSN2dIR1<CXQf-&RS7M6JSF#Wca#<VXY6FcHQBY3a.[[EW>M1b>NC78c
Z2G++RPM[be#JCeTFO#SeK;B0.:<VP9>EY+1fODb1FXg<UMVXY<4B[LdHJ:PB&bB
5FMf[^+;#JZ/6Y.1CMQOD]0Z__Y-5Va2M@QJa]RO15HGD+_2e55^6B)LfdA^6M4^
>;]JM0P;E);ODHGg.O^NMdb20-+#6@\_EdYG.Q^U<.gO7Y3NX4I:dac3>DH/_Z9Z
GXXf@<7,5=7#B)W:Z30f/#@9J18^4ZH^DT_Kg2)+:?DfNO?ACL(M&ccR@b<2ACfe
(\4UT)IUb.YDC==b(7M@22FDHFA4./(YP#8fCSeT5-9D>V)V1;(N6a7W9NeZ<R0e
/1QKAGL4JQI8a3PaJ7QR@JGXR(b-\OCZ#7dDOf950@c;_Ie##AN@++)QfG2+I.JK
M(M.Y@B?R?.e9-DD7JdB0FT2a0K6GaXgB80Z::@/faI0Z:N;8@>MYKH(_fKV(K>R
>b9H(J-?Nd#<=c(J,c;M7G9BN3)5LLQE.HUGPZ6G:cO4Pb6gUM1V3YR)B?D8#>FD
Yf/VdA@aFK/9d,8A@-R^JIc<O1P:,f<;eS#IQ&@c4F^#9f20/_&c#(RdFC_I.eQ<
\D<9OK31849Q]33DBP=D54Xd8(JQQ<#@Cf6YBZ=A9[3?DI3?FR@P2GD:JJMMR@/_
QYV78,?L5.HOc];3K1>1-ZI\N>e.2-?E]>P2YOaF<+9J5/G=Pb8f\#J)^MS93e=&
a2H_WXB/X2]C<]cA2,7E2=Z_\#S1+TKKA,+Kd?\J0>Se/?Q4Af>RB#;CH&J=@bgg
P6ZOg1Q1GM9/7E;N(L[V_AIXJ;1]@Mf#6a065&(-F#JO#QeJAXX3c+bCX,);B7_Q
Z@Y)L[Z1G3Qd,4)<V-?#5MB9ZF^)gbC4\,[,F5=e(-U4\WC9fR[&Z:3#g833./R2
e5.Z&>b2Z8MV]a(J\=IOHdX^6^T110X3#S3\Z9We50497M7FB)+cKKTW8/0@2XJP
bbNHS,;9,.6IL:YE(/<?8H:IbL0J.TR[e)>[YM/7:9.N5,(Zc8c4DLdTMO(2<0;E
\^=Cf9W36fbL#1(.[84bMb.GgJ_QX5VNa-88[Z&GXT>&Z8,BHg_29Fc/^,S^@AgR
)^E=QHHPJ47K@FN<+T-V?6c@?VXTfEXLM4+d?7e-W?ce_GXZ0.](^[.0JRfaA,XD
5;\dAgL](PEcMG_Q?9IB1?8GT@647F+][\Hd^5@.)KKV#beO5&dM88X+.30S)M0c
#7(.\?DV9JOH1TA[&K-BQ@)\?Ld&QGaPc^O.53@&:-1,Z_:Y.9/2Y1G]\^SCH,>e
HXV+A._]N;C.I4K(;GF<6F1:C;?-/VJH9J\JX-W8,BTQYgZ,K<?4\Oa,]_S+c?ZN
^-Vd@U\_6C599&30FXH@)2fK[4D=]FfG0dRRGIG\3cI85db.aLN<[3YM9T].\f,<
e_d2@I58/Q2Y:,e5aAJU,:0<4]15K0UeV69K[Db?9IG2LP17D07;8-BQXDAC<.IF
cM2c:f80aPZ)FF1+6Z(NN\](J7Ob,RQ^Z?f,9S?:Y,AdKPU=aE15,RI/?];&IHYA
3E)FA.G,a#fFZU=a5F49QP?D#G8/0VG1OK-^&T?RID8DULP[9/D2<5@:#0R[.bL3
X-M(+;(<#VAM--d<>4-HW6XQbYDE496<f]\<b;Bb(ZHa2(K8E_H@NGgdZASU+Ib/
8dFU7J#+>D@P(OHg]UABSHAa7Z6NN\-QF(GMQ?H,^GV_LZ+(.1RN]EU1J7&OYJ5E
I#fIb?R@?IT=4K>6<1DdWKL2UVSU9Sc1Of-9fQ0+;Ld3D[D,>P<DBe=bg7&C^U,-
V)B4)(f\F>DL5X;Q;TJ5aBHEW/KAL[.VPL#L<3JeT#HWG;/.GUI?T:,[O9E[ZITH
1SPeAT0&&?J,4++/<^R(Y8fXF0@J>)?7G7JF\KRdH;/a5@B)JCA-IRDE?7fVFV_?
G+&TaQ+g>.Y9(>eGNXW812<)VFe(IY]\OUXS&>X^WNI>ga9HW6I,]JR^#I1GedPY
Cd_#B3OT#?4/?@3\1QQSH1FTdfdfR2:P)+S5FLYeR-dB;f?B_HZ]VLQ)7<#]O[;9
WETC2@>[.L#R\\U@QWRX^7\CN4=Z?@IV.8MJ@BD\#AIP,PC.R]DRGM:>QRf]C&7<
Bg3PQX\(0]QXK)W(b@OK#PK4\E\)>)bV.,ZY_Kce?Z9RTNNZM2:220;G>.\5bU&<
+Q5ABERW9ON1KO9B=CUUJ4,(ZXK,OR<NDK9F8f@32VJLc)G:7O>+M;22-Ud=a]0J
02\&ZY5+_c?8gLK;-Ta#UC,PF\9Pd00GcZ:ZGF)0fY<9L;cd8I7CYUaa>I^.WJ(>
BZF;IgC<>DbO#F3FZLD)(I:g+#J^?_U9U@TTeY5+9>b]c7NGOVA&7<Qc=HY.2Y-0
,[GSGZ.BE6,9]T0E4bRYP\SSH3N]3J42[E&)&WG@N+19UDVK/PKPLK+SD,-XU,W=
@Yga58aS<@bbB)[-OO3G4(^L08P<;X+-X60,JGe=fgYY_W1_D@-0]RdP23@(VVdG
OT05Z6.B?<,B)I=._IaQJ]_N94J[V1;]YY9T7=Kd,B]1eb7S@-@2fCAQE6Y5X<?0
OOFHNQb4R,c+8.:CeI,WH6X^a:0)277^KFYF_3eVSb0Z=G1;O#JFCOMa@7)UYZ.Q
RA@>=8LR_/5GQe1#R[fD>ZOE?]J9ePJY(>-:V@;=91c+8e6_8V98A>@D/9MT7;UL
7Ua49P(dAf)[=X+=KBP.H(QNO,[:1[X]RTWTAIV&NP/7SML0YP7YbfJAeV&db&,7
_Ua6Q>bTJd]X.)>;WR8J);/>.:e+P39gKT3+,D#^3E3=;\]2]T]608/+AN^^F(IE
F)<a6La-&=R9]Lb2>f8<cSM<4fbY-T>8FEZU2O^0B>>LZZU\WNC9.\NX\e36XeQa
MZ54:I31Y[K=T5F6U9D2Aa4K5;0CEBfK#^@K5<;\Y&WHRg>6c5eVfJ#IV>S->UdS
F?O>;/^U/NSGbZbAW,WbFP/M<(WV_GPD@@],dGb&fVD=B(L0O1]N#8)RR\XZS>4b
GB;S1G?b=0(TG&TI[PQEc65V8W9(Od@Q3Q^Jb7aED^GRD1BN[35P5R8S.c,CE=M1
J&PM))MgNOATC(T#_V#)2)LFRL&XV9aK_gBH;WK/:S[GWK.,U\-gA_TAc\R#[XZZ
YWEP3UbYGC+bB]/&E)@R-Za&;O[9g;&EJ9F69FJ@&CObL-+GJg3G/]V-=ZALMdAc
(_)7)6,SPcdOCNG;HD^VPI<S,@ISA,4+IT;B/B@f(eMAM2gZ:LXA+dfNYGZ;A>Kg
.4b#b@]>21gGf1Z0c;Z05gLHHYJN9,:E3C2//08U4VTUe[2Q_2?80H?TW\YNaPCH
;B-BP&2dW(V,JT=,+#Y&E_d44>R/?B]30-FNNUH=c8bdYY<??4\IJL\-,N\]62J,
3DDdg/>K_/L.A+1>aVF0=6bX473+cD?/5acPZ1H_Vcd[8Ub)d9#W]eUCWAG@.U+7
73RI\]^.15]._\F^C_\08P6.BH\UDCJIIc&_3;Tf:=9BU)aM1,GLgI2RaCHUP8F9
#KQN9=ge9Z<3<;GL_]G_,T,Y,gEc?LSZP(0F:,PccUUa/U,H47BPS2JNOa]\e?(V
79\B/KLWWA/=b]bK@d_K6)[<7BW9U\P0FI/6e[3&X6Y4c^H)De&YUc<)HUC:#(KI
O4SU9VR[HCUP:Y<(f,e>O0PZUAG]05[^#ZAc\I/DE<Bd>Xf:Z9M04H+^67CX:YC,
-<WQ56.bWDJ.9g+[D^e/-3&BgD8XX4SCa>#aeSMB,4bA.G)G\5(7Q4#7Z:<aQ7Z]
6bS/3N8#27aIV-b?9e9(0U(14;,B9Ff,3K^0V[>^(eeIF)]g8\:W^K;1S6\+?3>]
Ig#+bU(fH<A4,bG+8[U/KUM#;1.)-HcQWB0O4-_>5CP0_O(HC(@CL@J7^TV6e,_E
MTP<9[B0__;C7+-b.N<aagJQZI01Gba+)/T:&X&#.15?d>J@SIfZ109H[8GPOFSM
e5bT<fBHg.c^JR)9?gZNSIbbYeG77;5I[IRHIY/:PFaHGQ_BZe[SZ>43d9E>d3ce
7TeJCII44SNU__WVHGHX5H+:?EZ>?c@N^^+b\[KW#efW:M_Q_H:]g-I\G?c)]]KR
Z2ABZQ4LU,b<e.8ZM5)]168cRZ#dfIaN5JHK.GIR42VJ#EX6([1>R2;-J+<OGLC]
00MN;-FYZaP@(JB^LG;]C&/.&EH1g;UYY].F1RXD4?JA(1.5A7:BWJ/Z4UG\Lc[3
KBZXHTQ[7X7?[T289W>O(5CG)1c<W;P9W;FE0eS@De6<&1fdI6EA#N70ZM7VNc0B
&JcWEJ:0FXQIASIg;&g?MYM#7Udg()fP-B3(PA;g<_9\332<0D=5_HPeS\.W1KS5
7b;3?E-[]ac.&g/U^Q@C_UdR=\Z@aa[YNc<b1;2E=\YP04EeKO[L+_UUb[bD]gH.
T.Q8<:GF>bMTZM^=::5Z\C0AYUGPKF^.X@<&IA?R28+f0;Wg#@aGYM]F16J6=-F8
W&WYW+/467/.\DJAbUC>5ZW3-;0U8H[DNW2WTNe+-WYPMTIJba<9)@cU/3#]&eOa
@&@2;T;Q5UFaRRPB6C?QD<@BEc^N1R^-#O4E93&-2OSd]AM>4N=W?P/[0OFV;85R
TD?H-1XcO?d&4Me53.[e@HI:F23YSW.TXI2<I=>O)ffIN.[570[\a0C5d.]L3D29
&2T)UQCD:)fKJ@)#gM8./&KJ<)A4_,4:-=Z=gBJ,QD<4c=_ET?B?5@.-WHKB-<J?
=L:__7e6^f2^K3E(.Z&QdEg\dWZgb=;2FVD]29#)=./)5[^P3dD0P&9Q\/5?&Z65
f:2TPXO<5H:+&MXSeLB64bI12G[g/(C&-BFH/U\0fU\L\R@;G;F+83,^]fa,8_(M
^AE#baU;cbT5([dAT19(5+ENS+I_R5GF7gVP4N#b]fKT\G\68Z<LKYcdSV067@.6
g0Ib3CZJI3TH.RRf:ed+^dHME.LO:Jade;3TU;ARLXX(BK31G,:7YFP-)K>JfAd[
6>RgKBXc5,#B0b>];6f@PU13+:EEVT-c2N=Z-4WcR_BG(YP\6#KR]]=+#FL/Id^;
eEfJc(,?cO=gg;\K7^_9DYAc&DgKE<4:QS(We;Rg7/aX==DgSUa)7;>>bW-^bV5H
3&:U#Q.)0H0MPRB,5@GaDeQB:BFM3G8:c<GI[M9P26H>gR7C,I99=\_dP[JHF80f
@^.5W]-OUGSd[),^\BN_T-89e0IU;PGG^#_0;)<WVQ]G<(QQY3EL)/K;44SXS)(8
Fe1(M;)KA,bde_4[-=0-S?I5C_.FFY&YU)c;H@UEFB;bDM<]W2O-9#@gTY\Y.K;L
g26b^[H?[Q[)<U8<<YV8&UUVP1=SWd0=7LK-,+&V?NBNHU?f>NT>#\FH05H7;X.T
8:IL[O]6R?R^?IS#]G:Y+EH0De;gB(UWOFI5JgPC(,S)C5>?IDDA1(L_W4UE.D./
f&.#,(@D[S04_)Vc>0UWYDUG5)G+YA_OGW4.H4dPe5UMdJB(>_H=<1M/B2c#>IGU
?e_I3<K(]R:+e7ZT((8I67O?:/.GfAPR[M=gP9S;HW2D&cXSY_:2a>f9c]?gL22d
_1fQcRgSN?W\.b_Uba#PE^bR&YbF39a)aT(YA2<5_U3#b)Meg\ZP&;YKT#J@?KG.
0LdM\0++[>9M_Mg,CGT@,C/4(FTFF\P>NGF=EMM^TEZXFB(TI(UL9+RO)95G5SeD
cL[?6e?c]Pc<2e6K1DR+5IgM(7-b\\()\<,<NR+XOg@S)GY6M(MGTf&][Y22d(\W
K_;HX0OH9ZQV/0?QdDVX3\1)OVO1^(JWDOS:\^B9[@cVT1R(.H.KcZ\d+9YY@8EV
?MQ/9V#5g]?QY_6eVfL6:IE0SA&[#W.2g2V1A+1#;[_6dI=)H+59c6ADN)AFPf5;
8GXWT0:OgM753Rb<?=FU1gbSH3#UXM.>3_J>af_gbLL-9c1-Q)N3G03b?e464N;,
2ddMeU7+U<=dB,PE7b#71Xcf,T@(Kc\3d.U[;@8V87CEdH5)O@+5TSW_^WYXd,,)
GD8bV;L7CAJH&C_HJEJGOU\,b/aUI#:>S+/N.85<XYc7\/fUCAG/#N[96N.-F>RZ
&Hf)PYA.P,(c(?6Df-W.\H;L,Vd=MR0F63_8)/0eW>0P:.Y_>E/Za@AJHeDeQHMg
G.\TR4TER3TSX(Be^9IPO@3M/,(-e#P1]W=gW>NK]IOI/[;,G_^g(4BBE;ZB-:-,
#2e&KdZAYY,cfU9O#dNM1GOJL543UX7c?TA@E5AAA2+gHM,45UcPCCc[AB^T?EK9
[+,5?FSDUK[H]L[\O.#6B1/(eg-F,E1ff+L=+[98OEB#?=SR40,WgHU/:d@Y#@c4
?a,8dX3,L1QCB@3G]92E7ONG:H@+/W/N)d.8Za3FA9K?)_D?7Qg\(^2U=M,^Y_:@
Yf)G>B7cX&4K:[J0L/:.]/ffAdP9J&J3@DBMG?,51)]7Y[-(4(J&>cX,U#EO>G-]
3DHKO=&aIaX-,N18>8_\d<CNAWOZ5e.<3YJJAf@DNOFdCEEXPf_<Q.MYYc?EQRO-
B^cG0NXScZ,HQ@g&C9J2:[:75eAdJdII+;B2R-MSSb#f.cC^?I8b6d]6QDX<7C1P
4?,;ZgIPE8f@BGJ]/.4,_]2b6J5R,0g;SAO,CBg_5A9#N3H+AZ2-8A5PJ#Y0IeL-
cNFRS/WDH_57CU:2J1>&]E1QQ=G4.[Dd0SEHg3Q_C/V1Qa<QL5U):_<TNGLQL9XH
=6?H63,MfO&=JFSW?9e+Cae(<:8O9LIb\3.,4POgLPW7b/=aSa+.M7T>04SBSYA_
]D1ef&gM)?J/^?1DVE5AM<:ceTVG79#ZF2.GF?3.84QfMET<I_MN^(&Q01>:;QDc
S>aM]@M?-B7J^1Y&?J0]8P<1PZSX9&;6Q7LJXIKD[952K><R2+F183X8TX\?@(ON
RI3TR0G<=C-3e/Bf/4/?&VU(;3Q6e)A1Qb:(V3EEfJXT&:1^90?GRA9\,91L3ZDb
?3bS6fAB,0XdRY;>a[,SAf.PG,)+3XMb0HA:Q(]5=b&M4\4OAdIBDTI>-gZ4EL-.
6QBW)7)4\U+12bGW6X.Tc_LOMBY=,QS/>J8KR]1aaW2f_d9S7&6>GMfdKN,)(S?5
M,O@N)F7=^JGPbRGX,eBgB]\gLHIADJ1D@(P3M/L/.IbE4[5K50&O#UfbMb)5?f8
/H(Ue@Qf492g1[6B:Y(9ZD;B8JRdBCC_5O8[NM7[@Sd:O_BPaPE;8d@@LV^;3fdJ
d#8NLf+M<(03P,\A#/(P7+c:VRFWR<G#/3I((DMQK-E;cb,<Pd6#3VF^.HGI\<:g
fP7b8]4d5W55N@eS<JKgYO<S6T6f8G:(Xf#_2R;.BL.POASJ:8PUNaX+]cHLCU/,
YF-_>LDI@9#LOC6X-UXX3F>,=TCS-D]IgA_6&@-_f@c&[JbS+VY&]4.[766D2f8.
efKM,\\#<Gb0_1@bLO>7[=?RD5F.bcgWPL15&Y0d6Xg^Zde>0OZ;F4(626^?UGD.
#Q[R?GA/::S(SQ#6H>,@4,8Q3OA,#CJcc8b_CDdA7RF)B.TA2f3:9NNeac_<W[f_
>7])<H?/=f;0W?VW[fUBU+(P49F5,NB/36ZV._XHd=b9AH5_CN+MZc;c2^9U9_Cg
;(_c65FPQffJ=e/B56dBT>eJ^V^L#UIfMCd8/e2e_4X<FNQGfeVfM;B[E?X1UL)C
;[CSIJ/VV,9HIN1GV2L_31(6T5\=-@TFYXM+^OUT(IK06;gLYFVKeHBHMf3(,K(9
g/B(V&O\>gXeTR77LbAHU#&_JGHM[1:S&;NPa,I2&D<:bY#(M/gcKQJ8R;6@HVAH
#>?64]PFYX,d[;=ZTUg92;\d++-+V,6cXQc>OV0_RA9+A<EQ0+E[g&BcRSGTU)AI
SG7aU7UZ2L7L]f7<;fgP11gbD5L57?J1U1UIf&9KF#0EL1D(]Q-9K#Ec=ON[8IJB
,U9VY5+66H3GO++Jad3g#=.CDGAO[^U:VV)GFQH5CK7/:4@P;@Z(<^?+5@2#PUT:
V;D,1:JYLb>XP(M_)Z<M<&Ra1FPP[+QF&GO0_]?;GLI0-eeOSe)Og?(ZP_03\D9V
^RJ>ORd6g3Tb5&D5ce[#477?KgBC.BM58fVDBE9]H<)[5X\H<75\^NUW06U=1IN^
77#12R4G6>,4QJ_\6aPN<ZMe8fIGP_BM@PL<f<K<.TQ:QSg.R#7Q(AN)TDF0fM_4
./FI<K->.K[KJURDSYg-a/\0Q#=]+3fMg_?9VJZ7S[fJDTZbb&+8Z,cXYQaD0H7S
^)0H=f9g3K3ICF,QeO6e(:-MGL_F8RW+W<)#HR47:13dda;BQd[cI2gZ4G#>;KJ<
P,a]Ha,TH]5IT.>DW_Q5/H&AX7);ZVSM^.)9fa+=_\,;54HI-++]/=<V1MEQP7E)
_O\8ZCYde8I6DMU1MGMJV@13.K@G:??/\Ng9@QbLWT;O/efBWgH@&?L]bU.Z+bgE
7+<.J?\We1b66GEG_R[98F/)\3&LID@@Z(IQ,I8eA:U,Z5J=3QVL3f)gBdA.=OcB
/b?RE^4U(GG0c12HZUf?T&J.WC57J3F#VXE>4)T:];L5-gA5/5#?WE0)]bDCQa=(
_6S+<OT@3)2Z2^ae^5A5_KfA[[-M9UDJ=,<U-+1,62:JEVPdIcDB88c4JBX=EcJP
YC\T@.W9DT.\a89cQNa1P:<C2+G>^9g@MG[;d94<Vc-N^8A.gUc#T8-/<&A,1d5b
OSCD-fRc3>P[=(QeUG_9DRF;WOTLSgD:P]G[4B9gENH.T<6eTIHZ5Gc31&70^P+)
.L0V/dgDJ7B&a)_eb?_S6EFLDR^H\f=^VPee:ObC\FEXcEMb.T2L0D</.f9=M(Y\
=BER6D^4fJ,TdH?-@N(PGJ.UP58<e#>V,+N/9::SK0ZHA;P;Nb)^-Z-a^O<GL[,C
/HBaO1KB\NaBfe;.25Y:1N_Ifa.2(?/B7ILZ+QKbgXQD8YL5;Y4>Ac>J;cEcPUYb
>)B)^LOa7CSW1P&6MY\#A9UMT>V_S[HFcKDFSK/O0:U/[ZCa@0@#f@>@._c(A=20
U9VeI86KSO9,W4BWd)O#eFS&L4adBEDUdgPf/55@T5MA@GTJ75:V6.^5bgDbcH(d
a0=+U]Yg&#?a[XeW-gG^;77JDR263++^LDE1@E=G9,DWb>06>(aGG1c-V>&O424B
P,P+F=1VeYKH7KY&19>^A15D2+>3A<3dB;9+#4))[ZETK<H=:;7=FG1XQ-3f5KT]
(eJ3K+U[dO9#W^-R[#B_\C7f-ae#L,Q[L&]OaP8bGX^9aEdUSLR4Z-^],K+TBT:N
?J+AE7>,;<=.,,</2NM;0V]=T\#8EZN938Ree(42ATaC_W.;YafBW?\.FL-9HbQ/
RU)RIHF:\[>G<(ZGB<Q[W3TN;JVRf;dI;L.(;@S78<d(4_GMdS<-EB8#L)M\eXC+
07I^OV=J2R_3J7f-ROSMA2/d8N@.O[D?)+B\+MQ4(<g:R>K1YFACK\V7JY^I5VaC
<W5<YL0I/K.f)#V^\_7<ZfSM\NV6bP=]9SKXOO6DB)gdTMa1b^CgeB>U&Y(?&5\\
<J:\9/-bA1U-JU@[[D&5cR74bKVYG?a#:V]+\&@LaOO#PS9O<@L7O<_TA[EdMJ;U
J=@&Z8:HSH@9fTK8<Y[+/Jb:L2f<#,cFg@SU@0DN7ddgb?8S+d</=Je[V:G6=g@<
XWP<Y?a>O&:)JGJWf)K8V0KbN+&+8GbRG15e1^\.\N^Z;>>W>QJ&_FG<I+SFZK,;
gf<_bSCQbZ_B0@M-b\L_T)058>PQDfIM)?V01IL]NeEc4E,R)L<GKb:2]B\f1efG
V(VQQ;Z0,:6ETZ)4P^5+I>&?1R_=<W49U,E&Q6E0)\X(bI<C@/c6TDJ09T8YCb_@
HXEH7Q<E:Z\:)\[KDSg8-7g[:#7R,d06c5.eYDBU)+\V21.F)>f]-,PRC;,#(AJa
^DD]9VX>?5UEB>2>QdN6/N^/S2T_XcBM]Mb[/;XIV>eB1&Fd)f>8_YE:JD0bfAfN
FH.&[A9WU/L^06SZZ+ZSO^,>X/<\?gG[:K3K>\ED?a(3R;Q<5GdaK#-B3+b\g]G(
]YHa3XOCDa[aV,V3=-TR)GK:;2+fW[Wc(XX-)^\H9L3:CE^604&Z@8[&#E>-8Q+A
7/L=dM.M.5\R@XU,SH/PJ8_3^Z.KY&BY:+/D7N:_Q)f&9<>XX9D@XM6C.Y4)M8KY
Q^fS)[6?.OHI;d/K5fF5<d_?#>M>]4U0((EV/11[H]_[QL25)TGPX&H.0L?H#F<K
YAZJ0FO7e4M.CLK_](\bX1<<P&V\fM)=]NMO[L>8Q&61#NMH8O8;6NX-P3e)V&<B
_M:<4_^efP341fCegRd[DWC0cYS0>E7>?#J&8:=?&Y-[/1/N3>cfDWaFSOM.LS)N
-gIIb@a--Y:R/#,B:#W\7]c@e0-DQK(WG[6AC;]K0)d7+-6LUT9IC/Y[Cf&VaB/A
+g0@Y;D9[NLAW@f#AS]Mg6VaT+4M0RXM]Q[,J&@f7eS_)_cS0.E0__#4?UK/<@2Y
Gd.J8JN^0c<K1]FG3(D?GJNJ8Z-PV)I<-_adF&_-3NBQ.F]5=^E6RRV@@F^a9\Rd
/USc+L6ARQU3H9Z6a?@L52ZS9];Y>+DT:JS.N<]Ta)E^<,FZ1M@32P^#Z(^g)UOE
B1K]-X.RA:BE.3Oad\+aW/8+M.K/7T^F[CX2N4IJRT9\M8.Og./6:?c9;&YC=P_B
]9e@+C:EZcT?.)B^\-36Nc.9K5fbDN)]Ia0cJZ?1WaBId8W@/:[D(+:<NNR.0)A+
f@0YC_<SegMTN4/YW]#8,#17.,e_=:;>IcERffH98ZdZ>1bdX#a@g[+Y,,SWZ^F_
JXISY(g].dI?H])8MHC1+RS(H1bV?+f-5B?I1BDO6\U#GF9)\N5D&X2PP586Nc,R
+V&O71K=P-DF]K:eM4-NK8dFVGG4,CH34c;(DLD3/H>Pa=5b,bC3fQ[cHX;M_?7[
_Je@gKAa.S9c1;ICH.<cCQ</#L7J,[(RB[_T&_;VCES</UAN605OUOdO8H,&#8)Q
dg#EY_,HH@9.JX?@,N_(3A<.dd8XFUBC&O/,4E#]4^6\C)???g9B#-]\2]+b-DYE
):74NJ6BEZcQE@2L:g7(eeMaLFP_K<J;7A3?gG]LMg)#PX5P0dU3<S-c^Zac<)R8
#.gC]=:V#EJ3D\0e_0E]e5d&YI#CXa@3a)P01B<&2I)OJGF=.7T0Z/QfHBXVN-=_
9W6<>:BUeF1IE]E9LJA?B2#Y7Ee<I)&3B8:CN(R-gK@N[K4KN2Y1PW:8SabG4R-\
/Td>@:VGGT;fb,G3X8?5:a&eKaUQfRYXeQ<HCEN5,F;.@DJF.Wcb+171>]fD-R/e
6c^g78CQY9,g0B_g;<V.<8)aEPSX^EC6^>[<-Nc^PG5]]E\IT&>J28eM)X]T.:e+
,>M<?P6OBYPS_Z-++3^b>feGUbD^_Vb1@b?,_dIQS&X;X@S^LEb;8dW[B\N\:UF[
M&MedK]-?.#[>bW\Y^<@MPZ3K0+V(+?.c2Ng:gG&#]4I>&(4XR<0PcPgMPScAGGV
JPW&g@gJ3VQU+^Bgd9_^aM@R^B/HM;C8<.Ja)DWQc]2AS,b[+8<aGTd#+,TY]4M.
?DWfC36Z-X#\TV.=.5bA@bFcK:V^.:BJLMbFE:.K=F&YR#F0W.N.F\F0T<=5/WK-
Q]/JU4a5dX3f+H27QC#OADd)>Aa_^SKP?)WafP6<<4/>_.E9=UVJ&Rag=1?efN2/
03S/G]0+Z)-^PaJV>2;>)@^dYUe[[QH\10OWGeML_-Ce55N+-LbRKEUEBgVcKRca
MGTM5,AAZN4?1EXQYBCQ0-eH&@-[M_BYNQQ6;H7D_07f+C>Q/2[]#Z,17)/6IFPQ
COI;[Y[S,^ac,-ZaK0^>.Te]JWR)T>KB\D^?/\8/#L)aS.b.+.B+a/@Z7GGF?V>3
VTS9RO3@^LEPeJSY[KXOCQ\beLWF9g7c[7LY(&N)K13_?KJGHg97:PV2Z8D+g1gd
/<^?=#X;a^#\CA;[[<@ZU7ETN)1dfXa49^ATYAQW,X>NUF>^-UEaJK5#RAJH)Z7S
>;8W]SLXd4VX9>#?;/+g@XJ?=YNXVG:[?f58V:014SE2B=g3g+KeIYE,E2B?UFa[
I\.DRITSXN#g,Vg.eP6Ed)\(d\>Q@f#bMJOVG1-O>0W\Z,7g00U>+PVBBVFDMSe&
4B(=ZMUH1+.,)O6)NdDG^aggA&,0+B?Z=-&\R[0,bYO<BBSIY6N2?f7F945_&/4_
2?1G3^\J;8N9@#@SRUCTUdQ#dK,NGQDQI5>V5/a89&(=,+5+,G49]8#4@CEJ9L@O
A4NKP2dZ4cgF2?Wb@RC79G=d1W_e-3>#TNBO(cgPGNBa:4L]gO8M_QH6f5\A-\;3
;./[LNL^;S39eYCB?U;f^#LFe(MZ:Ved7d0P7+/UMTJU,(E.JYWV7C3M]I->VQfe
e>DZO?Sab@8\@@b?dGb8._:g88R1Z.X2K(YLRUONOb/?V^<Rff\69,XQ7@&?DTPT
Q[<:X\,)RF9&44<+<7+K(8)>T9ZV2U3^9+?VLVfB+HP6gC;?\)&.MSTI)])58N/F
V.=#E/g]fS2>M^EB6-:0(J9#(a+0B#OBG;861g6?#EU)d/OEb.P/;P=<>\2U&bV0
f?#=Og);a-ZZ_S_@YU]^g/^LT6e;Pa\Ra0bX24@QeOPc7AGdIg9Md>YCQ2CH=;fW
\:X:VH)8O-:RZM9@G7SO5+Pe-T&;,Y+ag.B-\-QIUGZ4Q5>-aUbO@2M@MK5H=aC8
a_7NQ7R\]aI;U<.Z>TD-bP=N)85^#NELQDH3/)Zf&_#U2Ua7)QU6eR10Bd;Z)/FA
D.S[1\8aEIDUIAX/\Z31IJ\BN,/aP1L>0Kgd44TW-^QW;3U^<aDT6X8dTX0@&PT+
?]=9bNDG;5?J.MYf_.;@<.T>+)f(9##)6(/Y-;TQJA&.=C]E+;/45:B.1L/-1:,U
+1#eR<Bg27,6T;:WcN2O[G,16VB8D76=RNaWPQ]P_,EWe:X^Y:D8@bUXg:Z2?R#f
2Q/cZCWT(L\RNN=<@O2;HZ5-g1fF;@A5HPL/7E[HGV7K2[Y5).bd8NC)9A^93cY[
cKP?5]gD/DY1TQNcF+4G^LEE@E40gg6a[Y#1,0(3bIAdEfa,>4g>Q@,?B1BE>K)&
,b;cO/NEI?[:3J#9?3=-[S2=A56URK1&2JgNb?g[SJZ,c]+gHE+(W8HL?:8QAKf/
9B_^fOD0PZcgb:aRH^^QQ5]gSC9U<9cddbH;=T/8Ze,:HE.c20L41IBTL@)UCZF2
U4M8^^\J7bc<RM8S/cEgeTT.dX(_V5N?(+H66[[FZ]QZQ&c7^3E)2=NO:6KV0\=Z
bWGTc0]32(/GJ@EaVL:N:I7e#7KddJ2^Q79,FS]deEJ#H(^g<<^0-P<>V9AK>(5b
\AU3Eg\WbBOKBW#Z9OPN;7=W-OU:U>E<S&C(KS(ZYO6S+?V3A\,\gNB/d_6?Z.67
[IWFST:],cfJTG=Z8+UKA@JI&IK(5g-^e0e93aZIJMLUeOP^?@+2>HVRN+F0.L=b
0\&:\4WQ>SC-_KL&FH<R_&-(2D)SLA]=WU_#M[X\bS5@;=E>XRZ#>e&Q:&&OJaV=
=@&Y)b38PR<4JK0.J^B/NGRROTH1NU,.CS@KX&S2O3+a/H)&K4eCKP.LQVJ)g;=1
N6UT<a.0cOU>2K\#9SFMX4/#f^efR(;[3/D4R2:S-VeHX9K=O9EXL&?<]N7/D)29
-QV78F9d:R2g.><QC;@eY^/9ddSZ9E,((P.eW,MH4f0H\>e7[#dFJKE5#dPeRF7a
RDbF^[fX_\0D#@3f;@82N^WX<U7W3_\NF#9CEGNKL2Aa+A8WX(?2)SRR&JUQW#7^
B@#fB&0&B^:;9US^Y992W)(RX[&<X+E&:1QTGFH]?HG^eQJe:1]P@X:/+)V4Zb0e
e&J?,>fE+eP^0#/C)AE+YM)^K__&cNSHZCIL@+fUF_I@eDd+?KC?O\&c#&Y>Dd0U
OFN(D[dASa9NdVV@Y7)B/A:4S,I6Q>6;JOa<V[&E&Z/CW9SGg,Y]GXQB,4HgUd6B
.c25S[;RZYUZH\E.3.WIQ.A]XJ,>]A^U944KSI]X_FQND8:N#G;cXK,@8NDaVM6g
?D1QbAJY-5A8PTEB1G6L#84Qf6>-RE0;ZcVUKITQY6=/O&dHaQC-:F)S6FYgO)R_
A>60;R>=6^4.+,.:A/8,Q]T:]ZbgQ&N0OUIB)c#3GVb?O,Ve&V8&L\@J+7>@bGB_
4#(7?@I5R;C=d)@Y(ZB9T1.R.bH<c)[OZWRJBLDdHQ>;]JO\BTB8^54>_G=[O(?+
W]ea^.#,];>ga4>#[6(S2-H0Tg0VdWU)9C)][/5T=DFMOQbW-1bGVGGH_dV^9\7S
LB-:[AITdF84;EB1D@R60+612(=34;CXX[TF#&:G@+3USFZfHYQO+3-PZ#>\Z:LT
9JYE+)@g8@:S+=9K=7&RP#Zf4P=.\\6.)7B\;XM4_H(aQ+K5VSRQG9(:eW38c_DR
2RW;<6=;@@H0A_3g,PXGN<2M6-5:54<aNV@-HAT^/C<]YKHBU:37(&7AXbKXQOI_
B+(1X;?=G90U+D[\0+DMMHN9&[9UTaY@+^[33eIRbB8/YE5LfPMAFK&/.JbNN#1P
5X376LWZJTZc).UH+M;1L^H&fC+SN]gfP;gIQ,AQ.11+XV/geDVA\_X84]g-UHcW
G5)^@SJTOdfM0gP4=\c?>>N;aO&46TF.FBJ4^ZEI#I?4YO,NET+@DeY4b0PKHSeV
:A53ceeT5:&Y3F>+A3P_@J]NC;]e</)]S+,MAC\RJ=]@VJ^B_bd]DZVS:Z:O\(9S
5IA?64Z5Z,:g3MK#KLN8)>J:,5DAFbDY:6D7?@<(F=BYNa9Pc=LR>G#f[,FZSL<f
/^:^76G,7g-&.]0U@J8VE972ZccHK1)YRJ-;#:FQE#)8B_J@<8K4O1;B>2OI4\@c
FA)_(C[SJ8>,,]9R(M/X^cS6HM:>];:]=W&WU@:Sd&d[c\PLX2+TeCLL_+)g0]C8
M--MP[Db&VJJ9@YffO^0-^8:5N?0UA#SX<<N/8EcJDAF_B;+VfX9Mf0-E:>Md7@A
]Pb87+O@:\^JA9aY.4_eQLIS_8,:&O]88c&d6O9U-KSP;+,S[2e01GD&dNP&fKfX
&=EOUDD6Eb_>Q:Q#W2-=b^EHFN8O7+6V9D]]Yc#KCQf(Q:?@14aICL;89<Y>;6=W
g)d@6Q]2))L(OT;C7NaEQZg)Y&W.&CDffRCH/ZDZ[[#-\:FfH6RP8;b;]6Q=U([a
2-#,6KF]d3R;S0B(/#g8Y9I1J5<fKQMHVSB6JLLI?VccO.RA1(B]bK&FMEC)>QSc
Y<K,-dK-.\F#e-2>M#P]Nf<<>R7:J+/,.bEOW[2I/=A46D/.[HP,dT.SP>&.5:]V
97_fP4^OHC-(&Z:6Y:/QGZX2\?dG9+^3gWR7_Z03L0Td2.d]4OE/0e,&aJdVEGF4
/5&JKdT)0()+S29,4FS<[1^D^4NgESM2\=S-D7JeVQ#=6+SaUPF@U(AZDM\^^RFg
=D:QA,KDPLG?VUZQ:N8)^??0d>1c)[.BAQGW0_^5L3TX)JB)U1?4d/PcFWag;S/A
2@fG[S;[HJ-@D3U7#5)2&.0I>b?4Oda#VX//ZdaRfU2B:U-JVK(M,gId4N/AS#/P
gC,)3dJ_FM62]4TDEcaO16=Ef721UdKHN4F^,60ENa0aD0+T1R[&PX^:FF_-OT&C
@BF8-gOW:T6V.P/D7OBUB@cDE?-+K3W7.bXJRCL#O\BQfXH]]VOTX10-@Q9JN7b&
30ZM9UYdaU(#_)Of@>fJ]=+UA\ZW#KW]g93RN3JF31>T7T.6dAZ+NY?VdAg:1<31
4CB.P\)>]Yad1OW4Xe;+3WbP09&1L.:cJH<b?39X;R=0Z36dc,HC]&4-,bU:[b5d
ZNK<;>B:7S6O&6\-MNRYZ38:dWLff>-c9Ng;e9\:)),I2:Q2@+XE.ee[XG6QPIGf
W>[T6VdBX(#HP(N32Y,M>>W;:eW#71bWZf&0eO1BE5=H_TAcHPG>\8SYFbX5I]=U
P[;P+c<=7c+Eb-@+eBN2,cR@GN7QS)YgO#25#,L&YKE_4V55(9(I#\(:+UIR6c+)
1(AWF/(Y[HR\41&>4Q5P[@26,8IFF3UAA/6dG?=>W)H=g6efJE6EQ:bVU/Y9VAD1
T?FE93S=IEeXI,C\):F&0Q-31#X+HC^[1@&UU\J9R[S0L<4U78TZ5OUf(77X4K+]
bG?910UX_NB4,ZbdGKI9eIP<^>;SM,AG<O]^0U\B^I?P2g,7CUCc<e1GBDH>a6>S
g,3(\^3?f;T=@F>M[(]KAfWOZR=((82C/b29[2e081&a7V:eCe6[]+XE@R7/2;)O
&g>@VG=01C_P)+gggWBP&[63e=>XB@2G&P;#b>LJCBPbg7J/8UcN8ME]C^&N?eGV
:4V9bM_OPUf#SMA#J\=ZI-(0>64>QODbfXV2]9=7F2_TH8<VXZgW-NG\a[&8,NUP
/XIDO69UGO)5^#MBIE+A6:)07\10&HS1@YIZ48TR1^DE.fEMc[+A1<@#H<3:11-F
0GQX9CEYf;X&&+TYeIS+NG0M?IR:g9HQ:DFJ44f0V?O#XZa-6VO[cf+1.=<2/(U:
KAC;)J-Q\7cM;?0IMg=;>#=SfMW>b;8g=N-f+[b6_DfR_ZU-7,:FYS2]dd0a[Ke4
?<@f6e.TJ=8LLL:a&d#g^>c7QR>OI:fEbD_QC#55H=.V]bVB0_PF<YAc#d_f1gU/
??-d7JSF.V86R@Y#XR6)bVTT/0@c7H-+(;VdG<G(__745:N2UfHBLL-W]9IB_C1^
Ad6-21gRA#;3V1JSQ9f3(,gTRIF.B-G]\HY#>ZV46@<1eZ170eOLZ-f#@8GdAOMd
^OGXO@eDZGN#\5X6CBI6(/3f.8SITcb?PO\O>f;A217&J)S#41._8.g6B)/2,AHg
4)2&cEdfdg6-^&7->W8eN+2Zf,-V:@NPJ;R;/[@>8c.\X+TEW;R)gc=VXELUL6Q(
M6QI&#>A_O9MDE.Je+GDV+]MQDO<]gCT:S+e)D=@eZ@Q=.;G\YB303.>c&B#YL>a
bgO]K7L_8NCHMTIda:4EH5FSXB\4dX);=TG#8dR&,e^bRNO\b,XA4PV)^\=_;RHK
G#<bCNWP09:IWJO\f@.3DW)Z?;9XV&]/TJV+5\D<[Sc(,PBR-MRHDQ3bWg90>?=a
V2YJ2e4c_@CJ&/FY_3^:AGHI\@+M?9GW8;H(YM:8CZDD@TC]13=1EA#O;@,5<W.M
aaCATFXF0Dd3,X5a_(/?1MHgc<(;RNV:#B_eY]G598(:L2)T.(#:;YdM,&Z/gF/G
Z]8PQ_He<LN;)=0;&GEONS3gT:2Q8AFY#:P/G,@0C>?BQR>=Uf;4;13AW#7/=BGI
CYA&M)[V@B]Y[LBb>e^=O^8>VV?a35D+HcHVJDX6,)V<_0K#X+]79MP@L].JL)R=
:X_^[c[=K@1#F+c8Z0X97:=4:ZAF1LGC+5cbfC0Z>gH0]dE_7@B7OS&-5R06g<I.
g.D?A@(e)bPF_/gad>=U6&+97.N#VT0A=?9G]K)R&K13536A2ALJcAECB5dAY@O:
PT8eV1B^]97#G^Nb:1)aPQG5&@:NEAgYNU\QX5d/Qa<\TB=&.:Q.5?R)QSJR\c2P
7\YF\WD74#0eOE=V0cR8++4@\5WX[O2O,LPW8EGWV^<HW<>1H,A;ZCH6Q]]:Ge4\
bZc]6=WN]P_&5.)2N<gN(^./GT,9,;Id)C(FMKSA-#MLe>,AMALQF6>7MY6)SMIY
CM49DF9/Lc2[\XeJ@eEX,85:bHMQPW-H^XHOLE\5@#>XA\Mgc)_U8[YC_3@KfT,B
bdAdN)@d[(6420)IS]e5cZBR3#1)NgLgR54Y=9^G=U,YC2a@:PC_(5_0f4HWV]:I
UK+&.G8#,_EWfA;#b7FV7Zd(JDcJYZJ/a2_8G]#5#;>MYD0JMgGSdaQ<PSLIcSC3
W+(IL&_(/VM^^C,AHQ/db^GBA13]#]39\L^N,[F<#5Y0cUI-HP[A^XM4H&98YdTF
6c.gF9L5K./W8JCB>)<KCdO>.#\cZ[3(QTb4K:3^:<A:bKcHC)g#U37)>e2W;_=>
,7Z8e-#9=AM?1HCX#S:X;+Q^2C]48CaM8\0V;Ib8eg[&e)Kc08dDFQ[)F<#GHJeX
7c6)9#Ha\(4GS]+-3P9YL<b#aH[a),XSLJ3?R]L;9WI6(O+GdNHA0,F=.X?Y\eLO
L@b?a(1OOMKY&GF7gT6b>4:Z)e^]g2LgV4XC5/U\G#9UUI[eKe=TeNL1[a_<(Fd3
,6=Z_R>#UWNFMdF4X38YfSggI+aBW>TJVWA3/Q:BL/eC8DQC<2Pe;S^U#\FMbFRM
Q45;;MJ>6[^a:<HV?1-3Q0RAeSS;3YZJgY6\KL88UfS-@#72AIQC.:V+M>>QS)b7
UY^3YaQd?E^WQ7;]WCQ>CTB>H4LC,?CbWHI_5PaU:X/AFP<AYJJc>CIUBUM&=Wa(
I]>=NK/^<DTg61A6O214KEG;d2.fI52c\ScZOYB>V^(D(J+&4b(UWgfBS3U)JK\3
C?TVL?a@L7Z/8Y-)OO@N;_F@b+BW=<>NeF>3J.[L\MW8fON/=TMKc-V:bX_-I/:Q
<Q?FDf9gU?-8cXY1D]&@Ke,3\Y[4N1gZ8(O1_7EE#c12,LTA3:>ZK<^^WJac;^:=
(cQ8<;=DW.CQ7HZ5VN@YR^[IbZ44OBF9)<;RWC&=>F^9R]LR.&33GIUCbM(KgCe,
bX14ff6AZHd@/&?MH=,D/3@7918PC?8TEFOR_L?67PX2AaN>W#dG6aTMUME9Of=a
>BE>-=:(H+baG9:(,MNV:aUXBaCXDf.K_\D?6);U&>X6>B48F>bd0/\<R6YV,g^)
W:K<:\[?S^KAC(E(0D=f)L\F&PGLd:?.ML-FaVRFN93>/B/V3]4P0Bc.8<[BaA[1
ZRf/F;=]L.2IV-eAX3BS9<7e65V&N^_H5eH<fRUN31d/<@L9=Kc\K/.#7Z(OAL/:
7eSC3D(gcL87bPOAcX]U?e<K=P0)642IIESCL:J4+4c)AIbG9EOE/XUX)Zd>[\0<
Cg^BZ.R@;^&6N8HMPA&J/TQPFUPX4F:6e0WE(\:H6e#7\,=P:<&S1(.1S7c=I2]Y
#/-MZV&T@.-5^WPBGE:T3ON@JR#AEOW=P[[dY94C\[<UI;KAEC<RT\;5/bQ+[B<5
NK4CRdQ320?Y(0OEC)Y8cMM3Y3AZ^.T)>#f9EQ^&9EKdX-C_b\e[_#36[[LQ\V1:
f4ANK;[__+150[I(1(/V?FPPTZe-(g+<L(?3PM_3c/J/G=f).SY;1;&8)f\SgI71
;[FBHRU)?>1F75IeIL+A@D1#Q&]bP.RZY9FIeANMXGBYA\#c6I)QW:4aPPWN[Cg6
d;JQ[X47MGT=D#04SYWRK;TWcYI)TLGMA8N.:V;0Wf([#CN8&+BMS94<W_/</IW5
]1\SEJN?.2BC_Fg,2X[M;G-0B]I&ZdM#^c0f?F5Re9(^]=/@1XfCL&^V?#eOX@[#
2eXFP=/GI3\.+KbU#H+aX73R/)V(PZMad+<>#>?4]75Y<@.^@B;QFM#AHJcMbbJd
4a-[S==c2F=T=^:>HPc4/+J:Q_a3+Fc&FNH39)G=45+SRcE=2AM>:T3aeBZ/)LQ3
9E1_DC\2&AU@SNH8ZT1)+F0.D(Z67CH=U>/;5?6YY8@;\44T+FHC0\R7->dL:D@R
RCV\B)NM?M/TQIf&R0N9&VfT.\R7HQOdGDS01<]Gg0)6C7a@[;.2+JA^KMPc#/T#
></Bd0^EW5#[OP1?,Rb-eBYB(;7#J^O_XWa4gS=MNZ/]Z?#:RBRRA]XddD8(8)f1
I]48d,0aaR3\ADbFX#=cSLZ[cD9TV5&UIa2R/,.cdKbCASNNg2DGF7K_<LR(VP.1
OQIHG/^a,+eg]+GNaG1AZ0_5TLT4U#VLPP/N^KLG7VV#.G:_(9<(?c7U7gJg_>L]
7&6D^4E,A.TRaC8\61e\I5[Ia:66g)BMZW[G.+.9O82)QIJ8Gb@EK9I128V+Vf^(
?I-LWHd;@R+d.>/Og506@#SIb0\aGV.b0b7O00WZf7EHK_.eCO7>K896^Z87ZRO;
SI5D;RHF6#<RggEV+I.;9(Z(1DW<ZC\40.KB#Y&\W6J1D_[^5,2DW]BAca3WD?PY
I]NV[&@UCc4^1:e^U=_4gZ7Zda6Xa,P<3aM:d3dH8Q^:)4HV7gX@9M0OZe7aZQA=
T?AD.QLTPf)/fE?\a]_+CZV-Z@G-IbY/3@MM_AcEOXS6Q,5+-R0M/]3-cM]A?O-K
4/db[:C7E_/ZKI76JeN\7WDFc#?0@:6Y(BD,O3gUe-G8GYVOB_L7>g+6EAC=e/d/
>L9&>C14#3).?d1TH3/(\#<1AFVX,G]C75I?#.NPL3_<ca\#5SUO&JBZa1_UF^cA
g^.aCUP^AY@313[eK@3]ZQXCLR8NV[;=#@A\-ScSbIFV49.NgR3]_O9D=UHX9fO[
WI,H(Wf0JB4C<6TO[fR:2JZJT=&g4Hg\g<aHb@1AO6BJE^<>O3X5:S&eJ6\B.^&L
.3>U1>),L[&Q-[WZBK,/2SXE.(R5QX999,T6aS]=)LBAH41bGP0+N)7VP4b+F1cK
2Yf]K.F;MB+J:e6e&@[PWRU9)\:Oc-cEC6J0#/QLO,4<f1J(gE7^(VP^f[AAH[0P
gfAd4IGS(R-.BUS+,KN]^cG^d:AI<>e9#4E101D/;WLNf8-<6VQXJ4ef^\2_eAR]
E)HYE8A93g[GF^C5HS+FVA@U)D]NWfKaDfLSJBQ1[&ZZLbO(0XQFX?-;J:0.C[C;
K)/RC23[BT)g[7e).NM-TcHdEeK<A]UPSaGIKQ-Z[48)##NNM>7Pa2KIa]8(QP.9
L_eR8c02XSE<YOAA+[&50Sf_TND,\]\MJ(<(ec\a2Xg#ZbZZ8/BZ#R:&F_OGd[O&
:?dO<195NP@UOTDb2bJH/UOL/,M)Id>IGe,B4OP#cQ3d\6J-G=P?4Q70YGN#f?G)
8K<RB;)^=f05UObX__PW:S9=aH\BaE:A.\eB5Z62,ZEe21,cMgV3H(>7;\bggD#F
1+X&&N#KOQ-E?#I(W/LQf0WK+4=F,S4Z23/.5@7;G5@.e/ITed9(IBFRg>a\bN4E
?[g\N<U/5&b+a0@?@J?MeCLWaWWPQ3&E[JCICGKXA04d9L(c;@AS9K1Mb8AEEDQI
=Va71KRS0<.#HTL9bF0(C.F&&>>?&Z5^KZWE>15bDQHX-D1]+/RXN@TBQFKXc(.+
S>Ac?[QH[?>&+-RG0#_H6fVOXNDc;bQ&P6+4#aabNa(VZfQ\=6J]UI9f=OaBDRH=
adN0#]ZZZK6XV#Q>Z.R.1Ye)7Wcc+15KC[>>ATP+OJdeQJ&.=O47.f;0@6?U:OT6
FY/E_bJS]X8\gXb&OFcbg79)^X5@51\\JO2DH?>4BRgM-M/6H.6e=b7AZA1-PK[4
21DL,>4JB[R:X5bHbFJ9Q<[eGGLJ@4=6=>9^@_VI;fC4?WY/(\+XXN-<]L<;#.LM
e^]gZPeML/)>[2J/e1O<G+HS6PC/5<(ac_J_f=Zd&O+T]<KceN)Ye+LB[(A,RLWM
H4FDcN,ecgU.(Q4T,].KW?)4?ZV[ad\7HQ2++5A?bF,#88B5X:/-ZVg96dW688]H
Nd&#GNJ)+0Gab4d:0-JcX4K7IK#;#7_5K@SRDZ))Hg_D6R<UQH3c\=\_&V6_S&9Q
VJ2VPWg:1[;V@AZOI,fQK,d@BV8CH+BY7^YUD=67&,f:+(Y)-(;7UIK3E;e69M,B
I>d.EQW>FG@d7[.c+?UEd,7S0]bW342Fc,;;3JINE6UFBSgMa.M/?YScS#c49a(\
dDg<fA7E;<9[=)a79MJHa288NT^YH?S)SNVd,MMM3Qd/PDO]EJ?@_aYEIR-0M:ZQ
J-Q.=N^WBHOHCV7>AA[>#0)BeQ:c@YCRK\W4KUT)3GX#R_Rg60/Sg5bQJA7B90+O
5U)eOVag9U2S\;-2L_6#6aP24@(0a04(FJ9g]<?Ogc8736W)DNOPQ30@4LAK#CE1
M&-REZKK:6DNEcITQ;X1R=A6WKBFE,;K/::-WI-S#L[)?Fd]DWT@KRFU-;,K2^#)
85=L97;gfRBO1+9FC5&@5HMf>A9ZT3:J[/c<g,?Qa_e:Y4W/=I>#5fW5\:N-L8#?
E::5CdI,\6aEWAAgUSZBOIDfJ:0#YA&+BZP=:LST\SEKB&Ke@c=FC3QU7>eK+PV]
bH3GV2d_/B-DY0Yfa8VcB]bGN=e#<2&-HI&L:3IMN(Xe4Ha9.FKX,JG#(JOa.<D3
d&0SR&?&.TP;B:6IA8MOR[NF8@::8QIL1@AdfB:JK30F,b4bH8<gUc]S7.g-)W_Q
^(F;fO93eb23,aB1W9eeV)UW0^5JCgQNE.H\J>LfcP0UTdIJ#Z56NA=_++X;=Da5
XHf[;fBSc)W]]a5L&Q:L--bHSKL#9ZK@NfNc+#(,]0(/U>9)A0LWQ;eTD2O;]c]Y
e]?gG0c]6dgHJC(3+;GR3@Y(&A2=YJODNGTE<9KDXg)Rb1<_55c7)L,gGRGcNG7P
]GY=GI9VP?f1:Kc5a9S;CP:9B0-XV91HeP+#1C>.8?Qg.#P_42IKF[ccf]@&d)18
fB&QGe3-AcED=7A,Y)VK_DZYR:>][KWO;P;-C[c#C)BKC@C&d5_X><6:5,223C8d
FHU:F6Y2C.eKM-USf:_E37S<I1341F/.90+<O5+TTgW[Ne=^NHe#5IL_&+f8X&6:
XcZ4]KA93?J0-[8HL:OE7gRgW>I8E-@F-,c>0/CX=CWKH4?eYc:;dWKWN7QGUMHH
^P^ENgHZS@[GT9CV)I)4#L^\Ad)eYT41^56HUJR&)4J5Y\>LUDc5\<@]-9@\6@I,
KR(=Y1&0AbC&.VB49CdLc3&7W7I6<OU66H]OIWT-W(g6#;4OHL=Q?OONDH+aC(B]
6BUWc_UC6_Af(X9@K8;S)J[/Rg^6C?g[IIKJ0/>W2H.5F-;)Ac^N(T##E(T9a1CV
1TYMQKTc5SG;+6WIc2)BAVc;UD?d=I;a4N7>+<e2Gf)QF<gX&aeJVBU;UB;bR0P1
)SRT6Ze+>Y+V+SP]_:9Od0f6NZEZ/R:+=#TF1\RZVV62)PZ2-d3EIL<P(LTa#-C2
H1P>aU=<ZMdd56@gSM4e/IFbJ>]OC@KU<1If_D^PaLaW<A<IF^3;>8<c^7TP)cb2
(3<eU+;aPfGFQP#Q,08_d[VVZ[#RNZ^::(5YX7+Yf_c46A3.b:[5,14JROd+NbK2
4g2/C_dN:@-8.O])fSO<OHXZHg),S\BYI5f3-]::LJL&,_O&60gX@f&b4#f;KfZc
c+Z0@dE30JfFBX;\-Z@gX/]<9[>2_&Ag<[f@QfPCcfJCd422f-0YBMP7P4^8H9AJ
b=RcTb2e&@\144e:aSFYFaBegJ<e<,#2)&MbBR47NXSS0:S=DASg[/<eI>?a-F,d
?FMWCcY(IB1T0>EDX36@Q\,?@CN2)8GA\ZTe;5UKL4)RZKS9R1V6\[VWI7T_=cV6
_H5D)0X=\+EG3&1f?(>)d0I<NR^O]ZIf_D7;K&CQ(BZ?]F4_DWY\RM8J5^#b;[L&
#eT4>c/44_@.H3,1KLA7/4K&QG4:#D5F[J8ODWZ/KZAgJYZW1?V@N9P.<NX[9&HW
/TeY+YM(,?RB6C\PbRK@&/e5EgeG&D]5=/0/c<L5_JZ\1TJ6d_TSYA,)eM1g_5MS
P=QKfT\K6>OOCAK=I<-@,V^-/D:[6=QNK@eTe?Jf^DQ&;SLg4/9KHP+Xb:7,9LH6
W5,Q4eEg^(fFV52Gf\C1ULLGC@/3NP^J?B=))@P\WA>b&T/=UD@_._UFQK6(,734
OV2=)#,3#[VU-c>-N52E)P=We/T7_QF/E)J+@b8M.+gW&@;/R61RN_AS/Re@CObA
QEfPU&YbR[SY^b9+8bg)=T_bDfY#W1?LL.A)](CYC8?/#6BO7M(&H^]-5M__Ef[Z
&?bc;FJ4V<0;fWON7XHLIN3FI8b=G=D=ZeQ#3R.20_59\ND:8)b?9U,3\(FP_(B)
d6g?_1U(_]15=\Ab><M@JQFJRa[\FbGFKKFNK5WT,N/LGF:AIO3bJ\fZBP;E[=5[
/37eIaOIZ+Y1R;>5T\^<N&Z]3_(WDMW1XM(XHBg<\7800^#6)d2]+V(eE0(0E=QF
9T#d,L1LBL43:HT-@RU8A@UU,MI6\3F,e3FHHd7E>.\URO/-;+^2OZ0RbUR=T_-V
TFcSBVDZG&(OYFOM+Qc26dC7H?WNOOH]F_?[B#egJ3[?g:]3;P@4,DEFe+0U=O-D
RB0CNeF+/=JNJG2W]+\1)@1\2Jb^&452,1QT@[(DKUDXFWISG3U;9a3[f#eXWUDZ
5bKS-Z\&Y=7R@Y;<1UZQ8f2SK&DUM4Z^3WW_B+^A--Y@=DC5I)XAF?5<ReHIAP,L
?#@>e]_dQG-.GY>B>#:Td[5_=\&G-:f=@0^C)L8d9(0==geY>?;YXCFVEDHRBS#G
e@0V=/R5&@faZX?F85a=UN<bgdO3#LdJ8I>-:@fWAX5&-ZU>d34FS#<_.#-0[Y:P
\5[1&99b=d2:1d7[M<3D@[AK3_S#7??D2/8,T.Z^7H4ZRMLBWPZ=D@/A=\_#USG;
2CL8GK/ZC_eYG9GQ@Fe\fMFYQ)<<5cDCCb&81Fb)-8K,-4IG@[3(K_BIeY.14,4H
1,6K@^1.@9P])eE@_S@Q4dPdU;AE.:#5;;Z@B]OSBN,_1dUUEc[,9XeM(GI+OSK.
X/T:47DgN[]a_=d/AAbPN14&;)dfN)]bV[9,4J0b3g9;9+N,EDYJ6Te&O;M<\.@Y
5W8JQaHJNW4@Sf4[UFN/eQO(&7P7_Q#e,MNVW.J,N:b2_XO[H=Q[e1PV;aX2A_5-
/B]7&>IV4X9-cG2LDCH7:@9MC)]FgE,fRM1A]9F&;UL+_V^YE5Z7OAPXe=(@[\QG
R(W818DQcE+EK#4g;ED)<H7T2,VKRg@#V40L&A]:1aF/^Z#5I<&&T3,UD0=^<F_6
^[HTWU<BGZ-3^TJP#,>5P>Vaf7)+bC,HP^=Hf,9WIS?Z3eLcUN0IPN<QcU02DP7^
>3EL(=V^6Zd:f0bR3dP\VPb6DOc_VM\-c1Y+UUK&7S9[1P4>=@9L[RVE#.bO3R>P
5,9.:B.2CRd_FLP4(#E;M93?E4]dg511Yff/JN@?/(4<f.[).H5FR7e,15CLe2[_
-J4L[(:aQ\74/5b?C-BWPF=SgB36UZF1Y8]>7]PT949gK&5-Dac,#fO(NO-e:bB/
a2Q_E=:+=<:+-V93/>f/PG/JC#<ZDP&8CMM8DL:.XR?M&\947dfBM#W3V94>^ROF
:,0O>)^d^2ZFYJ[T),8J8Z[;IVWUS2K=^dY2J0+d:X1X7+S8&@M;\(_F0g^eb#Ef
>7HH,>=D)&g^g/,UNMe.LbH/[ee1KD38/1QBK#KC1BGVg/^G+Q+32@5F]d9SR@FW
Sf[_9:0e[D_SdN+B.[2(XF))a41T5Y+g;KaB1FCH/C31g6<R6-E6K1dF0,J6#(6J
cSWbM(YZ9B?QY]:.9OY&QJdKDZ1<=V7^]E<#6GESUG@Xf5<>R\U-bY::38L#e:L=
&H?8TbIJGD1UGOXRUa=SL3BD[4PF5I43UJC6g?V0AH9)45):)c8LRW[B[UD;X-F0
(e@?&-.LaBfMLSH>Y1,V](@P(1=7R?1X/&^L-GBe72TKM,/J<NZBd+W^]Q6S>DEb
[96+@<U\1NaQN;SEP,+Z,IG8&O1T-2dde^-/&+,GQXHg&K([7U3U@Q>+4IK&)b7]
/IFVH9A[N9<9T>2&>[+W10#QK)EVMbXZ35[933Z#_CYT)eQ-b.2SY9><ORM4==dE
/G3OIGMV0A#RY;OGKO?N>A>9.]\+0U@01=GS,ge278QQA@TGUfDTcXTb:7X0CLb:
9(O.>?G26I0258fL3OO,Q]N/IR.Q.Td\,K7CLKd3>LbcE#d3R98>@f839FT^T(2@
J>fQAWMA8Q8W?6D_F>R2IZSWMcP,7>6:?f_BQb:(Q2/U+IMWS3S];R;[V5EU(V77
G/&,c(XK,<UFK(gNHC<R<]b;6<FS/=f#3JAe\93P74QMfIdU_VO4_6[/=SSD4D-)
;ENE7eVDE?.JF#cM,BFI1fGdd9YPQ//V4.b6=&:^AJf_PHaB/N0[3.)8\YDZ?@0U
LYP,J6H8HOCXIFg+a9:=5eTZ:I.f#JG@2/2P5BZU]g5#:(Y(SIQ@=F,UT#[1I#7(
+5eKM=U6?X+gDW&BWIX<>U2AP^a@2Z\[YWA,6IRe_W+JT@NEX)H3bI3WfGdJJO;d
Y6IR/::]>?;cDD-UR=KfV;GM(UaG<I>-;]P[4&XbZA@=5U4N21BY+Cb#7-NWFX2W
B[>_bfVWH@N=UTJ?8L3#5=f\^/XNW<b2XF5Y(=XASaKL3U,\4.H9NOcc7,VR(,93
4JRBeBPXI4E\)e.\T@^]L2II:#2DAX;8ZK,0QOUD@+Uc/6e:L7NaN#,Mg=4/2+6Y
W?>&;e;R_.AeEWRK9/-1He<Ed#g/RQb;PA5&M9FBT9.&7>#I9R0?Sd\&?//eFa9^
R.>?M^UU08SDX4D3Z:3DTD0U,<7a/MC@8c.c8=YM6KWd+dCX._2]\/\4;SL?W:U+
O_>([XdXb,&8cIbC#gg2XDUW7V;X]]:RG.?_RO3MQG>952Nf_fWd^X9Z=MXA^g&N
\R#[I3T-+YLI-.&7EW&gB3#\0+^+:Af\(X;:L1GBFNJXTGJ>QBPX&\;H9?@HXYMb
R9@;.#FINFY#NSOW54/32ZSP#4MLP1\JMN&Sb&,HMSB_d^^@Q@A2#&+LSDJUP=<6
/3B+C7_0&5-0J;A;U#@A@WM>K<7f9,F:^9_GYNXCc4)=;N0);eDMR:eKZf+OPX8\
\84J;.(]90HU^5\8]->M?8V:;3Y_f7I:N#d,.cTGWH:-C=]1;=T;AI=CPHfF@@fF
@_-:TI]I1X7;CTX.^S._J.:CgbXV9A2a7Y)4Sc]IU0WZR8gG]&00]O8W.IL3gcc&
MBS<G8)?N;T5(VQT(BMD&^I9^J#=3CB^K)87^=;Q9/C/DeK,A=G5;9+bf=UJ>+A#
f-8WCc=&^Q:E(;d/Z+d:V&FLP67R(@a>/&Ba[F_TdG,\BeQW@cMJJdA,=4cJ-Oe5
&(,]Md6#F7,aJYDI39-2W5UaQ?F.dSMeG[[_)&+]ML)ee:ARg.Ke\F\,:[(c91WV
eeQ4D4Q[0#XfbdZ&I]W5:5W]ga00RG7@g<M6<C1JGCP\AVEPA]-1\U-/5=2C6XEG
4E1ATa#7d2c^Y4+W?RcQWB(B7+e8+#4M?eab@:f14,U&W:5T+2S_V3<M5McYIY:<
&3eAM\+65;U.:)X4Z^J^OaF&9&M74.K]8\UBc0&Mg(;[85VHMa(dUUI5ZA_^YX\-
L@YPTf#\JUS)4),DfRKGC?-Q5JS+02B:CJ+X&>IO:bcDHB^cF.4+J<C[]CA\R+(g
X-OWVYP3QGFXdS5cNFY_T:,C5eZ=82KN9MP+I#SUFJZEHM[VG/NO<5>O4aOa5TX1
dg@MXQ=[g4Dd-9GRRg9RX>T9d,[VXW+-\+f2;GSM@>U?a=[K6QWgYDO:DF#O\8/E
_fH]MN-PO/Tg5A6=+afK-T.Z&-e?397/gMP\=^Cd54P5:<\\J/VI>F09R^,<>)&A
T@g07fBcCcbF8FI^DKJ(g@6-\&?g6:):gfKX,9C<KI_S(OM?.IEEA^,,ONSPV5QV
-144-9/C]9,.D_=b4=XSY8@e5LCSDeDH;.\HU5XN5\dE?<Kd^__=E56P+Lde<0ad
J:GJ+F5;YUbOTI],aOdP>Tc+Z&>c9(a,@-Tf3GG]NI9V?W,=a9LMdEBEQDAU+&3)
N14Nb0K+/3OZQ#aJdg6<;68A>f[=WUCNN?U_?T_2c2-aY@Bc60B?UE6geM;K+4V4
UEFHd485/aI5Nf)PCK8P7S1f9dQOAeeDIU2(0?eFGSJ577cc[WcGC287+_BZ)/@S
6Z?0]:4[P.Tg.MLI6-,]=9OA+.O0Yf9Z+(bN8#/>([8XTd(O?5:aSA05C4CAV\ed
PGF6UF&30W./f&Of=>=U,MPK\3Pa(R/c[KXM9]Q[=:#[_e;VCf+FF@IG:ZOc<O+T
(F/fI+P:@XBW+G]c;?Ka-+T4^Z8&B_L^C)IFMQ-b@+A^(.UT3+:XNOR+8>0DU4>>
_Mb<bc3SC/B,-_XDJQSZc#^AM4#64#FT1U7<dY:5Z\#_2>?6+7b?4+NJ))bT;1;Q
4f50&G<0W7d.Y<CRD+RWeK\_A=1]<bc+WGID9TCTB1&[)W7@IAT)9b7ZHFTOQHOF
/-?.+4P1d031O&eb1eE-B]JE@DYTDd([cZUGKC.-7TZEACEE#KE.O9N@0=La)RO@
9LO#JOY5=:\(V<Sa5Pd&1Xd.d2c&W6_(EI>+&aQdf#B69UP@KKEVADM45b:919Sg
^M<F+Te271+g^-,5Bf,:I7&&Ye\e4<>A67HbLdXgQ56J_47B:aI1;)f0(5NLd<F\
=QY8KYQZTM59^P3T.H,J19L4,U.L<3HbB-?483#AfAJ8(\J=\]8/c_TB9GDPOH4>
B9.22bW.Q6B)XDd-^U];9EeNAOCKXg8UHc,be7=VGGPQ/8_CQXBO(d)2,d_Be:D:
4?=?)#DYJL[T-Fc+A+WT?XN:Q0aBXS;L(YMCSXJ81\Q7YVWaNB#GBD4dL;LdYTCB
#J6cSDb_;X;5fT1^2^2ZP.-[^76e\U0_0c/2AF.6Y=6UTTRFf&-7S;J_KE[ff;O=
8==8Y#2?V\Xf+a>c_BB3&;T__Db_A1N6,_SUH-8NX(K]ILE<DY+G8#6=Y9HQ3IM#
JDXL<LWb^^_2-Y3\H^bQaT=I+cT.<L+?L(bARgL#&#8:+,g0]92gJBJ-,1.VcF2c
9L+Bge96\,3I>R/;D6KOWQ84H>[gPQ@O?9?1-J-bOcZgJe(7QD75.BHg1HB9OI_:
g7//EAET7)\_T)FBb=Oc2G.V=<cH@+AJ\029))7>>TWX;J0:671XX3PPL5eU:W:6
XT37M.N2MX;;-bY]NT:#g<(.H<I5QZM;0gSa3?DF=U(;7@G78#^U^P@RS=)dGKDE
@D<GEg]a)?7TeR4__YZ+&JM<>A-AM2(=?]\<2?:OC0(WeI1g]374f2^AQ&O/.AF\
D2/cONG20:]]BI]OfRa)/P2>U_a^Z\Q:EW?T29XY[JHREA]S\?,g1\ZRaR+L&^VV
b_=K(NBQ@6e.B;ZaO-@2E+,OHg9EE]Z8\(Xb:^bVd\#SIX-e92>S/-,X,U===:^>
739V;bEZ&,O^T_Z88P+;)R/?Z&K-A9f]+[=),]4OJ,\I-]OX:?9ecB>SOe^Jf5f;
bX78\=Zb7&g#LeF#a5#3A>5O;^>LEfQH&dCL1&2D.gIS,(.=-C.W>;/X(Dd69KC<
9-]Pda]O@@Fgc>0M#A6K4LeeKH?QMLg\/L_D,AR[M<JM9FeDI0X.:KWSHX6KL&CA
I-a6-#?(3.;I;?)eaYg/\K_a@]WKX9KFe=3<PcXVYHL=D&Ncda2A0>L#X0S47^VX
U[FW]_>M5,#AN3;BXcdc?>]]A):HK]0WYF-.+L7U5\)Xg7]8cAMZT\N(XM>&STSd
V8DN5aT3X>cJ@<=W?CUPDDV^)AcgfcG:;[46X/c4H0Ba9JGZEKWOU9;=X[,QOB77
8?#N4BRL(>15JB<d__RHO?+TO]/fgMG][-(D[<Xd3)3BeGXMU&cOC\IK_84cBa_<
TJM;<ae^0<JRXO1WEbG0/EV-T7U=LQ2@:9/,[4WIcK[NJA\>9:2<Y_dbMfG,[H=N
F22)@Y5Lb[O46Ng4)\bdM+NES9DN/RCcKQ3D+CME/]B.f>c(HJMfTW\>39@X;P>V
?QaK<-b.8HU#,2<+VSC788X;@F#ABYT4X/\:>VIf,bWVI<gNC.3H?;I;X66[Y[dI
JP)4S&U?6de.[+gP-,IQbfbg+S32:8O#PQCY0c=+KHGFQW#@FB9<73U-]gdFa+4;
7YGAgQY+N[NP5dQJT]#2&\Vb+^2Q:1R1d<(KbQ;6\MRK6-+G+9266[2^#WGf7-A>
NVK;V.C05GT->^2eHPb(L(51>Y]ScMTP\2=^QMG]32cVQFBDd/)aa7HbYX7+55;L
HX.3e,FQ9XBH0#f2>/74BX\-VTVK:=C9AE,c@S:6D/_XLW:91DUKE;=GgM>+RT1V
JO;,JU(#I_Ad/.=ZC)&Qg[G.50+?\8Q^O^Dg]Z9e(0-C7=D.7J-aF?eYQ]N1Y18@
ORX5ZEPL)&<XBXeO>[F5KZCZ5)3=Y)Xd/QeH(Q[;<QI2<KQ-Q&)V?19Q#,?W2D.]
+T,35[AcYf_DL]Q7I?YcSX-=H@Zb=12c)a2&/E-^R>d644&a7fb:6)H=N\@?RHMZ
M>KK1fKH^03[\K[R_1=NJdGY-;YIF6?&P-LTeGHfbTb;G0:bTW9MgG6&dND]NM#?
G?-VXKKLQ[&<#2N4-<Q/_GT?@QKf)J26_=G(cLCOJCfPO2Y5gGf99H,_c:NC>P[1
TaG0-=6OO+[)1Pdc<93,&JeO\P3-8C<I/R0>3_TTE]/Xca\#bE@fQTKg07BdCT?a
UV]#O:E@?_\AJHEQ?I8,c-Q&e0&]LF@XMICHWb<9+C/61J1=,)UXU+)_>../=-IH
L6;YE+8S2W:Z6]Rda#M8K9U;#9fOZGJHCI15J)/G-14P)9R#=JE)F.Z;P4Db)Qbc
56U+)N,cHD8bC,/SIQDR8NN_bW]X?P9@<PCR-;;>bFT8C2J0[G+8eZ4?eHXgMGQB
LYT8S8V^@+C#SCM;D7<(KKC;4UPH@Kg=PMD]5G5eVCf.^F6S?bS2:S^c8RK;_6P^
X+A5Y6+/Z1CXL;<&+;ZKeX5??DF/)P]959Cf<O?T6ZH#B]?1<VWHKK3#7;X<g>a(
M#8<V&_A87[f7=N^?RNLRZcaX5T:Jb/;.P]SgYAfPf,[1\2+SY@I52+0^-KIF]gf
AA&^Bg8TT][?,bGDbbRCDP]\M_3,D]f5)?PQ[^JZ.ME[[L;\;dP>Y#_IG9MD3</)
b2M(OE+4DI,FDd0e7__;X^P)N]R0c.9YH:cQPTHOQ3.WfM+gP\9bSfDUM)?P64W,
]:L]HT,Za018e&MccIHCF2&T,<-U?KJH8R5-9bDb>0W>1&+.6[/XD\g&R+^S;cBg
U)BGJAZc;RQ?459HAC\.<c2:5>]X+_.eM2.T_<^Te;F,]HUe^YGI8Jd1DaF5O4A8
0HM9RC;T&@#)=.O3e&PBW@R?XH>@4^=YXUK7O=/8)M,[8gVJ[]8\Y74GRTO/2#8a
KM#UCTO^+)dAFEN[XMCOe/#7+\ZOVc0&Z7UcB1?E0OK>YJ4]C;#f5CGX2Q(]2JL_
QG>?OMC)7+c]#--]59>aOI7#Lf&73F@(JZ;fG];-0dMX-.-0e9gNK?DZKdaa&-R:
AP92:OcE+4CX_bX6.3B[;I:MX<8&4bUGGH=IYg/@CNR7C:^<:aNRSc)#06)#+?AN
f[1J_#J8]F;Q@:I)P2&LSD50TR/[D3(B7.@N0TIXI@+JbOMR=K&KI:T\)#OC+99T
VO?AOH46TEO7=.Jee;XWM8Q5C-9fUAQG.I]-bDE^Qb=/?\8N6LTDUC77#EVgfH\e
:=>]::O_AZE8d(gB/3X#8&?7NXgL9PC&O9MT^H(X,7]>Gd-@[PUAMf+cC[^N+gS4
ZZ[ZBXYAU]W&>N;FQSPJ@)XLg^]+H/J/=M.ebW^gHFON)^&(J<_N-?58OaWXcCS5
1;Yg@2LTM:^4PM>/QJ]Ne60=Tb728eK0&FXKRG>K9+4L[fg-]I#TVcc_7&[)_)F0
K-U_V^Y0:^HIPY]AZf-.=KC?VUDMc7Pbd[;TafVdK95^BJBdQK.[/]M.GTQ+/f2V
GYLPYL6NaS1Gcf^+3b^,X37VA&f0.FDVZ:8EKC[_]\^BcGB)#E58E>.O]P?2Y5KP
_Y2/<:fP@^87Q?e8fULL0;94/LaS8N4S7V31F\C0EZUK+,<Q+92K;3bY?1LU6PGJ
RTML7T_LF9SI_:NB1fUDSLdd3V/KJQB97:1b[c5L,fSU.a.f_B.>T/c2c&+^K#OX
@3aSJ[b<0a3e_NBR-cDZVP8]NgPN)HBW<>:C,:,[D4_E>CW?=YaU,,e:)?&^3ReA
\-6bK_(L31c9-#-=T]H0=dC@(L7^g,^@Ld6-/XXE5XS[CF>b,XW3VCXHL1?,2T<a
><TJNe2+JP,WCA)JVBg.@2VcT5e-[)PFO8+g>9J1/S@W.(_U/@22O0Y5<UYFZ:AH
aH5Z\L7D2X82:39dQTQM=/B(::31@3)J?Y1Nc-32<LN_Sa0b>@#Q/S2R5N]b18A0
=fT?9TZ/M>]0,JIIe8=Wc,KH[T<^\2<4UX@X/dP==(2=N_:#g<3&5RbN96\3e#dY
N[CR@I[S:e(b[S^B37O@9>a[\G9YH8,SS/FLEX(<NC;MWYfKICG1+RW6:&#P<<0_
gW/G&J3g.L4dPaY=S7_?19^O#VLZSdL7YTJI^U>Q_0<.<6NQ.c5><DR/0L&DAg:W
;ccY#RGg8:)FXIb-53A1/1(e+>D1ZY]g/-0d0dM_+ZY-LAWMVD&.[?P#6=SV@7IM
b33FVN1Z(&M=HB,D):9d4H>Xd)&&RW>EKIe[[O5>087)N-(\:,8/Wf(G,921C:<]
E+6<H8>);1cEY#]?L1GYUg6T[^Y/JPB;A8P@10C5MaU=T/R_g;18Q:<7_^9\PL>>
K]Qag-#FEGR9YRHcV1\#,>1afe2F<<2&ZW?9c)(<c)?51DK<@Gcg[K:[G\dG4SV=
24.<]X4LN,]NK=]#4]=E);d0<I&)QZ_JF([=&[@7(TO9/1XTOb.#,(AJ3TcFEJ0:
V@\B;>+#YPSQIHZ+BM[:]bI::8AaEQD\b64>N>-?Led,J=]6\25U3;+4edc^1ab4
W&T/1[1KeaR(JSJ?ML_BTgSDYZg@8R?Ia[.P7:;V:;dCN\.HN)CK9a05HS9\\+#E
)R;UPYFTAEII-DW-K:@S8.#-^-1/#?#>YO(Y>0fcQ,[X<Q0JD0D>4,a.g,a#49a_
e0_)O^>@<4EQ2]RF#^J_9>\ESd47GVUMB9cA\8F233+=)cG4N#[8YN^/P]SDPb0Y
f3]E+B:>@\E_EXdd+3Y;]+fVaZ0S;TcW:ILK&7=YHA-bJOg4BTCdVK_[7L?0Y1TB
(OJ-?I>1f.@S5:JKB@b^AEFa9TEJ,5P17/+0SQ_P//a74_N[_)&?ZHe?,c8bg0OE
>O9_@9,)GV?O0WfQT:FY\0aU-6;.@0S>S0cYQ:368b34FaT6f3FH&.U_#eP>5Ee<
/02((LK^.-FNG,#Yg@1Ra.T0?5I<A.,e,Bc&Ncg-,VHG,4?abHDX\Y2fYI2)9-/Q
^fWCPVB9Lg\DTRPG.+XR_+)Oa6a7;:\]AA?DQ[:Ra=Rd(8+Ka7N_e9Q^<M8:\6DG
2J)TB/12QW_f<+L(^<b5C@]R(b]:)SbS1+ec&#aF:79dMR5J?>Qg5,U]^0?E3.>G
Z-5OG.MK8FN(g@E.dNgg7aO;eGMW,[>:a6:I3Y]X.b\<FPO:8TF6>SWcE&.D>^&A
?6eVU\G;1MH6abACbKX?,gS&G=aNac@XBL0>2U[gE0]#Md@C>BGQX:b@>(Y]T9O^
OgC1[)84fVaI@#b;dBB96.<Q&^FW[cNJ1-,FH9a;0.Q36;g?O)ZSM-A43O-<MH44
,)[OQ&AUB-QU.(-6@/O50R)=/4P=>\W/QW\8(MY2X-MdB24.IV=bS;)O?B2cDSMV
,6c/W2e.:a6O@]IdG<9UP[Z)R]Q:4NDM:\7?3XE>-Q,9UUQ?F3<K,6/P<MfFS0CH
CbT)c5U1V=A)D8WLKA.[N0S8A<dVg[&4I3cP/f8W(FYRVGJEb:#UQEL+1^5@7d_O
F?V-?#QIe6M[0be//\YeEGW4V6]9+V[BCE-05/fH0Ze>G<_4d[J,@&GSPZ#3WT#7
<Fb)\2Z?T2-cDM?SWbdC@J:bH@B(?//3H:.9C=^0e0J@=63X&>[E;bGD>ZeM<WU.
H<DeQ,;)2bbQ\gB/Nbe5[dc3R<YB9aI]<aW8S&#S<ZgQWE7CHSTaOX3)d-W\B950
?e_gKI1X#ceOW;c)[:CMa89b_K-[QSMP:T9I6N(6_=_5[)26Y=>6>D+5a.F7BBb2
SP9Nda3?R,W5C:eAbH;GX(=E2F1Q9MSV&aZ<C1QOX/C:HO:Z-9FZ-bV??->c^TGX
Q87=2][&gCH3:738.,LNg^MW[JO::2ecY4;LW3a]b8WKMf?e,b]K=8gDV[V@QKH@
1L<JJA[&TaUfgK_WAOGa?#AC#JJ3L<aTOXEA[g0Q.GI-4]P]>9WMZKUN2NN3ET,6
.LN6I8ZXa?2+:0FF_.((3)LNFG<;:UUQc.GOI;=DBPA@GOA281K;YQG.gSLTTNPY
V]dWT>Y[:.-HL8DV9.MAYIVL+2XfT]KHZ_BgPQ-V]_]+Z0A5=;XJBW6)1]L&MR.R
T;_U6S7=9R_8W2Z=Y++Zf6Oa4_.8?9d1Ca1>B96ef3bc(N.Vc7BW+.O.D)P?YGTO
>LOX=AdF/4@U3=3./H_4<39M7@VIIaD5SIP&bV(ObH+L79(4d._WNODS5Ta?T^WK
+017V)3QVQ_MY+T>/-[(fCbU@)IdJ[[AMK<[OGFFK^@WBSacV.fb/&O:A<aX25EU
CK.[_d+UGB@\d\WZL((G17V,JO&]-38IB_I@8&@X?ISbW_?aDX=\)Ze=4GKND]DE
@GA^\EOKMgMP]15(\[K2?(ee8?01H+RTVW/\5CB7)>QVXO)f4N[IKR96.)&df&FG
a<8Je?1,0@?[0eDCG&.DZNMCd#3RY8cFJQ;.:+CT^DHBT-VE\@NP&+O;0B4XA=7\
IbcQP_29GKR.:[P>bAb.41S5KZf[c5G8YQ/Q4/F/KO_aWC/R695YOAc\JNe(egC(
(d;GR-IBbER[Wd(d=F.QQ]H/_9dQ3bGSf.GaR?>eDABEJH(gTL.^_ELf&=F]Nb?;
0cVO^]2RDV.G)7;D9#]:9#:R-\=ALP]PCV>17bF3@JW8QMCG.9ROSN,&IYL[bRf(
9IHe0c7,fDHYeLV<U:OWb&cUGE]cb]KCIf-?Ha-T1](Q87]N:4.]SY)Yf&Dca\YJ
L9d,KL:ZFU6-#a(:g5OCeVaBG0Y>07<@5<)Z[T-R5_H:L4LMFW](X\V(U4>SW(]c
-]+:&1DIb>WK8DK4KbHUR?78WH_-Z@U8R^5-Z/I7\bSc#RJ^_]1NHN0G&1B1BW<J
K@eH9?J-JB47I[HUN\Wb#=#NZJDU,V/90ADc:&KJO+,BG\3Q?e4FTW\TfFaANFWV
IUX/WV?@(3bEge<b<OQ+=J6R(DC[4<RDGUB_TBe,/5()F+YEg.T\VDB,[A=W5?5D
bCHe,4#d.=2_2G0?WMU1MJY\ea,:0/#L@&\U/>B6O;O7B<&]::]>3TR)2P9#=Z1;
P8+Q2+?^--0T[#LK9C#FYP#[5eAaZ(DDe##EL,-,QCH0Q3V@]F.ea,,Z+CS@TXAU
A.,#2G9DGY>gVR,#S1Y3K94aOPYKWT5;W5Q2OH],KWACVf@+@@K)9=+99A3GT>Ra
AUaZ7J8):[/YIQ,J(X>TKYbXVNA4_;c0[>LKO0XWOd8R-Y?61g;cLL[@5Ga7F9?K
&C(_-K]]Y>-L&3G:95RBO9_N)6JCF9c+NUcG1]6BMK,:8)VK6U>TY5EXWVBP-D]^
]b&\WO78NDK\9bQU6S]6Sd1M[4Z\,4W[J&G+I,F?93gVb?<b(P[c?WD7Q9=ZNOS;
;H#K&d2=f,QOKgbZJ=NI63BD9=+_-PCF@#QDK.XR,&=AARVaDa?#A+GFFMXgA/\2
7eXQV+1\I,ea=I:P]Q\;aT8&PGI4.2aQJB.\(f+&:U9IIY9[:V_/Q&PE[7aaF3R=
MZ/^8CFdA/9-Y,4P;>EMD1:]&1;6ADH3OI9,,O2WW<;QS@B5HT[&-6)+=4XD[/@I
;9d:@gH5Wc#OQ#9/.Z1:gX^8Uf3#b)/&<eU]a1FRL?6WC9U[0#:W8[EZF_4Z;==9
G:<T&K(SXYM2M5b/,C;/0dJ]P)SbCK=D>eAN[RW^]IFH<@HN5Cad9SQCHSG:XR>H
&L?>PM)[1\C_Z=3_&7gWC-TLe:\]#c-\e]NE(&(K??O7)V@5M_6OQK6U\:I1P?]<
EMK\3bVW#AcBR^D[9_T00?Y#WF]K:W:-Qa1XBC01f&Ga+V8RUPESP5PD1)]LT\;A
U6C_O,N3@Z[L]KG?>7F7F^/1=<8(I;F-ESP]7FXVgILNP@+&g/_Xf_^^>EW8N1eJ
PTK7KcA2Ze]/VgA0N+^gdGX(.T,[8&ecd9bMSWQ,OA(ODcI+,69g>D<4ZfRc@aFA
&=d<MS5COW<OO\PYNIdI^G:&)7\gP<=JRUS5[QJR>E<X](-8ZWBQSN(1gT5+G/gX
C>59U37)&@ICfH#N3@TH:^Cf15OAN_bc<d/6HaY1?8eF9L88^CL1eAKMSb,R1A##
g60,>2AXE7GKSXbd]+RgA:8.)_LS,7bRBL6g^LZHHLVS@\A<Ig7XA[>B1(@.6:Sf
-GGA/Q;=DV@7cWZB2NUTSDgVS0E9e>49bF#@ZPSD==6L[R])1&#+;#8Y[[N4_AXd
c68]K1H9\:1^)1NW.c+UfU;&DNT#5]E(RE&;R,RXW([eD9X?#eD<TaWZG6YX_P(9
TLdC)K(^1Q2X_9[JEUJ,=(e_)S=\X7S;C=-+):.4V2,+Ue7&NK33NO;/N>CTT/[U
MG3JG[IAQeXKBb_TS0JG>8LLX[g:8SfR_XED2GK(UA29b\1L<\X>?A_\^Q0bK034
K+.eeEHW3XIdJ=Pb:]<H7O/L5QV[_Qe[MC_3JQF7=.]00-Y:EdR]]+V1=&ZMACM3
_W)ZWN(YVa1cWE(+(WTB;+CM;WbI,XLWaQ<.b=a6&OcJdT<,O<CEQcgWe7R^)BId
CCUf\g6CY:b=QfPWg<[^D7DcR7)[ReS(.Tg>D[@cSU^eD+<DD<#P5cd57:;bef8V
.?9Le,a1BMA^:+=_ec73@Ag769/\X>;(87XV66L;RTKOSCd1<+Baa,;f0EU()V/5
c@G=&XIA>Pe1R\P+)Z549d,Z2DJXcH@QTQ/C_UgY[0^IBMc#6DF6^&ZbDW8begQR
>G88d\eJa7/TOcC;a(B4XI3bWV7[KNM2PQ.)=BL=c2/FKZ>b_74f^5c.>NTaRcL<
(B.,Z<\fD=H[G-E0a(H>+D&&9TMC,0)#UN]4=GGdIBR\_@T]?UDHOC4G<#P38],#
,TcNYVfRU2UDe=@9ZFJbgODE#67L6?ZT)Z\VZ&.[,N_J6#N_+eK4.#ABHK95dFKE
g9W;R_VO0b6gG-a^)QZg#0+b5aBaB/=_2=(SDADLcaZBfQL@A&2]H1ZBT<Zf>a<(
M-3\HQ1WR643[87LPQP6&[N](+[G=8V>(WQTg1>F=cT?ISN\>;8=MP?0JEQ[YP7b
L^J8FK3VQ3VZgVAgUc/F>PF,.>S>aYRCe=R#/[[UccI:JCWGC##3/E-98X>+(&;a
)a5g1B.a+H56S8XLUNK)M9#DN0AYK6g-06)N4--2DdAH7Q]CPG-dT(WXLGWVIONN
OWfG:aLH+8bNXQVC4L8\[M]W6MT8a13ab2Sb703PP>HVYA]/D.b:\A-gS):0K^)5
#Rd]2YC@Y\5fbAT=N1Pc-27FU_\:1#11Q=F0a7YPO3g\J#6-b/9&^,@^27ZcTHXO
4c3;#\5L1XJa&BNdaD<C5G\QI2(S[eX[)S+&46G]=^LB@#JIF7d_84^aX.:GK>^,
_4U\8;?3S1ZF^9X8EVV(F-@]+^2;FHVgSeaBDH/=F?P<WJ<7G^d@OE[W(,@S:\<J
bf36_:A&:e_DA_Gf1A9RTIL5(_,),2>HM+]I2D\<VZ4USKGJ#0QT8[JNM?F;.>J3
#MQ\gYPO[)7W]Z\fY+gJVCfccK.+XfUD/3B;#WKF6<R\,eC:Pe\S/Md_PD@cN15,
)3>)<fF;5C&a9g?L=V?Q0D]^4g+5YFKRUB_aORLSf#d9]:9_U/cL\X5OBM7f#bW2
)3KHY&R?2Q@#MI1eM<d>+/U3+A^MM-3[g33R?^6#O\JR,())?gd&H^[3EI4f5Z5c
&+KC[CO[BfbP)CRf((;gg6;Y0RSOPgP]6GL2])K7UeV/?IO.M-:RKY^[-I3FcIHc
G[>HO&:Ob]9C12g8R4W\6Y<cK_60=TR.K6)&.X)0N=27;?4G2bX[P4O0&+&J[O00
gN85:[/dIEX^4+=OXO;WLQ.J-U+\LG4gc9TD/RZ],1Yc8dDD/X0/1:U/H^^AZe7J
8RdN(AaQB,X0P-J(<IS-<.Wd_eO5M&DRS=S(PPF@>aNSK;2<;XFYa[e7P&,7AXED
Y-.14LeC>,,dPA(7W)^=NC3B9Z#Z/<M]SKBZ>G2GF1KNd+e-8G\VL9_gDB\QPVWZ
NX027HDXc;+d?#/S:Q1(a]_#+XMBLR-@>^5D#=a[=1RTU_[^&ERN\_Z33O&Rb+cN
bUSW::+ZbAe.\#\(=CX7eYAU?YTbD)ZM.GEe3Hg>_V&4S.gd4:;5G^KUc04T41HX
(^\RJdZeRg#>9>1TZXAOG2BJ?E5=5)E<+V51O,A5&c6&:O#=IHT>a[LV_<9MP2ed
)E[[K@?F90-a(-IEECOZQ,a]R/@Ag-(2DLI,f8A&+G):ZT7U?EAe3;-g[8-P5:#<
)[R5WZ;<9gOX\3E\D@\c67e>c(J-:ELDOK2&LES/&?gaA#[OdRa+R&eQ+XOJ(7)=
K>A=QXBS?eUA=C,&I5RUT]0;[708]Pc?1-4gYXND5L=A&1#=O]SYB<&cANWDcOH3
:[GAS8XW[0,+5CcV&TbQ_NVX+P[TBRO2cA;3?08(U.6W]/W4/OE#^<,=O998\YcI
Y:M5>QGb[4J?143Z8Q@GSLMHIe@SIU^B.?+gCgMfFO]YSGW>[c;6]SM?NHB<Bc<8
e,HJ,EV(^T>;&;:2;b62I4c&#Z:F3PdGef9]NgT9d0#IIR6;S;)dR>+FCa-aPbQ4
#]_Sba][,A1HBQP1T4V;eZg:[KG4Y13.(&P-P03^DEL3)d_0LT@2P1&YEZA5OMR(
dQ+\CMDIGYA<GbKdPLQM_b-^X@\gf=a,02E=:X\KBL2+LK&eQDTU,>>-;7a<A0-e
\5BKF>W<<?EeTK4X(&]J_6WESggdWeV)4>_U@>I[OGQ7,4]U^ED?DPd]6dBg>U3f
W]Bb<eL3_?RgGR^)W8>KBKacO7<a+&Vg9T+gC:80^4GZ3IFce33>:&MYVW3YG_55
.FBFCJaG92UVBeD<_Z1-]KXfKB^eSUgF\GOITJ;[bc@<,<]_5V>Yg86fB57\5YQ0
F#efTYYLYPXQD34C.SVF#HTcL:V)QFgQIJI@a[=c99M76/^IeXTdfJXL<96BEG?L
Y>+c#^TSdFdA_3-7RZ510D8W5:\=XC0P>GUeT^SgGbO(]6bCXG;f@=<<G2P6MJD;
X_E46PU;WO-&3FR+a@]-LYMG]YcO/3=(d:3YgSR8W^8C#Wc3L>(WAeJU_6:629OA
S4<O<#Z1-]T+B(8&c<W6O4cB>.e/E/e@>=e4:ZI5Sf?^<,f&Na_.GOV41RY)1;aR
M,X4FBB]A9L-(3[VgB#=cT;VH)U^A+,JU2K2STQ(C[0H?f2-,DU1/D;5[S7<9Y(V
50@B2A4M\UX@+effQdR)DI-@QUZ+3X.@[V[AKJ/Pce&_D0XJLd<4U),FH3>/Q^D:
]2JI-@>#ZD[&)+)^=6E2LA6^^QE0+UgVf8,NeZ1;Tf&10;DBU;.+AUCbgPOa<^/^
(D^0P<ZP=/XcgPSd#/YRVC1+e:53cL0OI_Xb@:]]R]2RbEFVKG7AE?bXY5gBH/&H
2a5LN#b,BYZKT-YVLX5S[&J)0Q7NNI.FcQCHe-,9;(#1<gI;>bGHE3aF]38gAD^D
;=2=,_;S:+dEM8FTA3APX7N8?Q,G4WWJ[bH4f2=\-(cX9<O78Tb8I.Qe-UH+85d)
NUTHg0R_A9MGcQQeSR>G#V5;E568(Q(<b91KBCAe-F?PWgVG1092<\=M7FeTeSL6
8DUCb>ECWTB);+D=9O.YVXG/N#_=]WPCZbE=[X&E9CG?Td1(ZgFEWe9J-<f_dKdf
#FY6SPB@UCL(97B9/cI5gVUeJIB.PCTE:8H:#cF2<Sb\5),\12PLL4(TYR4T&8c\
]@Z:-eYPO4HL0&(C92g+fOJ4B,&e^[Y/@E0^a&D-1Q_:1_SULJ+89;X@1DUK^DIg
3G+;-/WR30SYXG;.6cDL__-?G]:]D2g4[Y#KIc]b,EUCCadELDB&4dHUQ@<S@^WN
.S1XQS1^Rd3\XY85=3IcEe3VKGHC#C:99adB:?V)Y>URF^U117T5[#Na#HV2H[P#
+\EJM@PHN#:fW:?DL,\Rf/>C1YK(D<(@Mcc==(+JO2D8Z#Y;.FJG7g[6#FOIYc-V
1=:)C^YFbHe5(c0G[HQWADXZ@)c_><KR7-6T^=:VVJa:@aJ)(P:-2DXd.[^4&A9U
:DI9@gOeWF/@,^EFQ._ZYZ8S@GHSQBaVR#1JN=F+:Ng6:Q889D8__&E0f&>@,(17
-:0YM+C(/.R(<CO]ScB^B<)D7,(CW2aeL1CX,A8D?&L>K2[WTaM56NG;&^,#DdA)
2][gQ.3AD-+FC:E]?8(b1EV\9]/(52^YQ\ARB-^J:O-A;(KW5e.B5K52.AD6-PM,
aL30UeT0GX<8];9SIDIbC,JTR.?V<C7eH]cH=)C?0WUER-L-g2bP=67K/AU+F+1L
?P4X93G/[9BX\U/\?dETUU7_R3;HA_=#>8/\8bSGH0H6?C3Ef5Q7.e@LJ018Q>,M
??/)G#/IFJC5a8QVT,I7NfRSE34O4[8LeAB&?2LF3UPUM/@&f8Q5H>8FQJA38cQQ
;G6WTJ&:)/GY;CE?,-QV[].(YSaAbD<CF.5cHJ,L+c]S7T&6]g[X+7Ga4e\>AfZa
2;D##cTbYd^3,_?0D=]O_Z@D[:[0]17:]7TffgLH2&1bd^fQFS;ZRN1;dNd<L6XT
bAXHd(O?4\EH)aI;aYUCS76GV_H1a[gFKAFGa8:Qf6=?,NH<S,/^D:9E=gW+ZcW;
g+M@SCEKLR2=We\<T=\JC2.;Hgbf-PMV)JXJ;7@X)a[C90;0^0Da(FNIBIQ,PaY_
O12&(P:3dJVN6C.2K[O@5.HI>2Db@dBF0GFgXFNF]X:>Ka3;;_]V[01#&:0DU-]0
VS.]2bI449>F0>]fWUN.O5^Qb>NB@B]95;9EDGXOKP+-eQ;1[eJ&^OLV4#+K/)#-
@cgZ&)E&/3V]_9&/7L=A;:)<A8MI09]@.QG.&3;4Z:(+3g2fPMS7M(CZX.)eO+&g
E&bLg@?eEAXBK[Z(-//<[CIFgN.;fcacMf@a(?AaOcE-(QMc-P@<6<W.VH&1c4cN
D=;KE6ec].11/#H[+P=M<V]T#;^gKORVaA:4H-<)D=XWXR(O?B.g=1d/b]EZ:faY
)]f34BK)6S11,]T9F5<Q,3P?eGY>(HR6d,d_PPP[3g+#N>c#/2:aDTSVK(1&bFOd
.5c-(:)H#08@K_<84=T)M-O-+K/B:g&VV[KeRLdFBW@VP\HF.QT6a&70A9.+M?,L
/a2)+=STf2NFWNY^+,VaFd(E^eQ>gK1EKEf[1(NYEd#M3&^PN_OWZW+/Z(CVPO+G
CP>W\[:GFC+O(R9c6I/<W4f(^J6O)Wc9(fYQ.7:L1/GfM<=K;Le^Ua^3ZbBb_,]V
F7,/V[M#]]D27b6c3,P@H.-KF6;197BQ1A@(+fAN6EC=Zd,[GZ8\2b48gDRCMY+=
>7XE?-U2PP]NCRN3YQE=@<]N1#[D3-c<7K(QS^@/AW&RR<J8K<35A5FFb+&:FA\4
e+g9c<1,SO\_SeU<b\?JQHV)-6R^/.SGHbNKQ-5UEMMN6=ANOMMTG2JdIQY<,I5M
UCBcG9BW=PRKF9(ee>>d+\YL<0b=.?@NU/FN;NX3_AR<H<W+H9]UdN3b&cg65T^:
+?NC/AV2#GQ+CY07AeT59?33cQT2>O=TB5C@(XL2&?22R:M(I?9ESJ]WV[cTGVI\
^MDLK(KM>&0=@3,81e./QA1W4?NU+f1;\7?GMd,9e#4;3dO]fRC#7)KIe4_KVa,[
Ma2bMP):=E#?NfAWRSC>(JX;Q?A(3/T(J,<:=Z.fa::L42RgAd1UHOYVYd<A:cKE
BCTaA1P=M6TQWZ+,K?MPN]b>Dc4gEAVgG/W/MC>2EBP#6R^N#A(3N@(;TAS?D3V5
E#93XI()PH0,BgN:N[]Y2g1[/edgWLD^ZDWf)VeSLZML:&Ug2e1VN,IW(ZReBMMV
0@@NJSgR2S2TJ@\?::2\8WcZ3Td>cXYB-N7ad6K6NY#C3XL&aJ?]a#6IBTKHWK;S
FX)B:1.bWKaK9>caTH^>Yf@KS(-BFg\06eD/d(KB;Q]]^D/eAF1X=1ZXZL/=9JI+
,GNGVOU+81IVd[KAafUFW]AABbfgQfRNHW7a412J3G4:CZ+<E68)C+Gf,OTXJGc<
(^]NHW;/)YW/?\1R&]/4)5=&.?+/;XeNY4;,adg\Bf8[1OVO;V\f&Q\8QJB-f=&0
/_NDW0@TDLLSaSY1GdS7aSK=S@W;TMC)FG10:M@T)V&RW1f@A]72__Z1C(L3C>ZB
3YcI9I-TGc2R#4-/aTA0U<90S@3&f02Z@NAFHd[<(YeY=f,07@\C]_BRPff0HMY8
8-E//I0V(J/C969-<<YX&=/_g]E?RE>B<^X\IWKKK>IW0OC>Ma\fD:gb^<S].ag:
O^^0/+>=1dG<U,0OREUKV:V[CGN<N\f40.FedO1NSB[?g)RAQMX,R6^+G>I;>3\F
2E54T#cAZ)FI^6=&=9b9)T-09Xb@9UK\gV1#V=+##/&aTK)L)CU7-U4Pb)LS4RCd
0@N.^^ZI;,2(dZ];T;VR72C)QOE7]N?ZYHJdb7V]e+)/MFEWCE[L?CF]34H?I5YZ
SSD<WZ:0?7e[Dba(#TcEgU?-U8P?bfF/8FWE+D@O\E@1D+HV:2[HDBCY:g_EO??R
.:(D65\cBQ.^+I-A/ENMc_+-^JO>70)WP:cK2\W?YM:fW[6/)O]XcTUc-_@+H0BU
42aFU1QT=#9_9e(\NQJaUHDM\F9Mg3@UDEP\B[&W<)9OOY=bT8)3L]Z47+N+XdS<
f8+V,&;C7eb@9ZV;@c&O-=>G\;5QK9S8=K5)HDFAad@FGS81&E&Z\L;JX/<?BT/B
FbO<8.2C&_EABcH(&XdK?4I.MdI\.HLM8[:D_N)&=X#+]^<D0<c/=U]JHS+LA7&F
<f:QTP#O#7G^g)&dJ>]DVZ_^NU[LIY1WOVHL-V2J64..LS)E#._[(L;UAH#J0M.2
>c-.I(G8QRZI./)R(^<W,MP<_C>1.b1e>HRbafG8?&QfeRS.]JO6?WDcSY&+1)+)
g2E3@cg4deAN?10U_a>-)CR5(6&WBHfD80Y0Hf)UH5D9V4E;FB9.cf[e=VZ9EcJC
6>K?a2CfaJ<(@0]7;<;X8:_(28T..I/0N>c[D_(D\IKH3[E7TQ@.NdV),>(M.?.7
+CbQ\&eQI;aYUDKPf^>DTLgJ0XC2_^\S6U:J-?IgKO^=?S8g,Z&+N/(-C,Xb,]cQ
7b^Z>UYRQ.3SRPJ9,O&RQSNA^0^b4S0R[A16J+PYO)FD0,L3=LXV&_C0MR2QG6=@
:-EYAOCVOCL_6P4f]/\3fN#6-0R-Rd82Z,]&3;5C7UQ:K-KL[J,W_/ER9#6GLea#
],M2K5T)4.0M48NP3B96A--YB]P8]cV#H&,gAC(2eR=PDI\&-39Y&SEf,R1N-6D<
VK#LWY<I^&4^dWc+g]0f2d6O?D5&RL]E/=VF@C7H37.ECV+4^^3f?)-,aJ<Lf^CU
C5F=DO\TWN^-475IR<+;,[I#cPMFXH0eI-(CDDa8\e9UK+M3c#e0d6\)ZR;BA3Q3
KebKB8R>X/(T:)[:+B>3d,M<(FB@G0ecC7OZ[[3KN>7V.2;QG8&81PbJH3ZIV@#^
+LTE_a>,I-W7O=#4-EfFDbgMHR?DV6419G;?9VgQAVSO//f=g9?-P#a3/=]XQTcY
?]9>b:RU\E@T/WCD^cKOY;/,B?e;3&O=e:2ReY:;AD&=<^<M6&_O,-L_+^+EM^5K
B.#4d.c@4=OS@<0:U_.8ST0ZZF)Zb\0gBd_I;7_LTLf=FaQSV?>5A>K]=X,T?K(O
&a/V5bWc[1G9I<E=>B(J7g+W\3WA)04143>OZQ;WAM-,3b>U[K7-QGbU:\2g,N:Z
QBOZ)D@HU=e@8?1_]DT\K4XUQcPafT,eI4DZ\-:0f00^VKFa1d3:9R::a^5D>1S0
K93>;cc+EGK^Q/&Y&\2(T/5Z[X08ReN)R^U/1F1.;W[EK;eES+1PC2\4]H53OV/2
b\:gM0]K)\->0I,H,ZS9747LX?cWgD>fPLGMQ)68I.eDUPfeD3#S-D;:,bV1=d:#
aDD<Y:CVMFG3bG)^Fd66\+ZV:F;5-bT\\2/GIA-;_^W:/CggKGg;85_51-.a/?Qd
WfEEN_gL(VWf.:e+dQ6N^7+VfeDEa@bB_2L?bcZG?.F>H&efaSPLFEHK1Qg,K-Q<
8fS/KcCSBW3V#,@g43=BL.A3FI1-APT7&f=I:\G+cM-c6OFV\0bG&9AdN^)K0Pe1
LKV>Zb:>8aEf;59WSffY]P#1&)MC6/PGZVI@IXNTO75C?W&)AT1E<ZT>[AE@--?<
e&;e,\2c_OY+S&QTOA/GP0ePM:Nb<M^YECU:1/]#J#LF0TSFA:33)A(\Z6eV>7E(
a\(^eD.RJ\G(SKbL./]e.,6XT,@=eNBXK-f0@?-dD/?#PKb#Faa4/X-WRc6MOgO4
I?AI_<;5d#06Y;F\S(MZTEU+VO@8cD9FC[S_&:1=RM3MHRX6K@U(aACA8a6I4BBK
I\-LIA0&/L,>Q9^H-(adY]-JW;)DUQab+6#1V&[UA7;J+<8J<WY_I25M>ELM@,T#
&XZVIAW4C+;4]PUJMB#bKaB/:Ub([4e;G+I=JfU:7,D)\X+-eYf37Sbb:7<3\ETW
@aJ@,@8fO@[[-9-CfP^7]-8(F^2R25b(N)@N]A]G_3F#_>&NV^0QW=g8Z;/)OND#
7VXFSDST1,<<#N5dRZVJIZ:Z>G8Y(c,1/1S4@_CbZ8#Gd:bYKDQY1U?L6+Y6M-;X
>&R(5UB;A=/#J;M/V77J7I3<f0&)T8-2>5&T]H6G.YS&ZcA58LF9++U1C<5DS=,S
:T^AH4e5)H:]SE9=IW\A.?5/170USW>)S4[gK(<(6WWO4WgLN9:<N@(+X?V\RIXH
d/cSMA8VQ3D+HU^#YE(_<MDFJS=[RHIF]-C7.b^gQbXZ7F@IfD@e)#P7Ce9ZcR21
?PA[5T3^.C+gUW+RgMUd_LY-b=E)J.YLYRV\TJ\)dIZ&XDdPKN93XQHQ.AX&N]#^
:7S/A=g9&+X?A#2?,3N/C>SQ;1<@bGZMY>:W(b2-_<L5H?AfaW:UgXS]Ag#Q2ZBG
Q)(CK909?0Y:M#4:8DA39c5(ARBd=NZNc:+C]ZLcT.c:CT#2;?WcCHYV+^0_,@W_
PQ5PB:6ZB:bL[WU2CgU+3Ia7;X_]\>;3TJ[CHNJ&EEB+gB.M1L^YE24>>MV0ZYSE
:>0ZX1fF81B[G82^PW8ME7_PAX_?S]H0gI2e5/d@W5@G7TMG#ZacaJ#5+dVQ0M<I
<M2I<BZgaVA1AUDL?][-e7B59BQX3N[&_:QXRCYN;08P2Pe)-WN;c9:_&FUKV,,R
=,I+e[ZMX=H:EC7>2:O)c2ffO.E0JH\-1+,DV<C&\9gIU<g<6I<[2JL#fO:)N78N
#)J8,IbfCX79V9N_EKV/:/3fgQ&Ugf?bQc0Z?W-0X:XKO0?)-[)?_BM+NW)dPIa&
3C-G4T00ZSD4cSa;>8f(@?^RFYU]/@<M@A?=,N<.XH/,PYH)KY\&_ED.MX(g@H8e
c3+DTbT9\[1fgcHCH.JU/DF:QQO9geQCAeaFPaQ]J[g1-d8RB\Vd)fVV&BI@Z\]_
d3^&EO2^)RD\E/GMIO6SKP?QX)WR&De^OBW.F&YA6&9V;9^YP;/BE\?9:=eT4N92
.gEB;5cd[H+a8O?[12[/+<>SV,(Z]UFI.e&#f,2GNg&5dVafZd#4R)S+WY-ZgA+[
6Ag64E\?((L=JT^_a/@Ce#_Yc&MIPVNMY.9@3A1fRVNYW2cO_eaWOG92W=-VHdN]
VLVIceFGZIL:SDCQK)#9+E)GIU(2LdS.CdD)Y_?KC<&B4D+VJ9A1IX-S\FD-0.IQ
7gc>O^4#0U-K\U1]/RP0(:,d]OPg/JV];bM@Da=02G(9&_/Jb+:B8(QbYZc,G7..
EK,5TV,0M:gQf9VEP=Qb<IGGcU-K8X5d=5/dII)FX\dDDFT,[NQN;;X<DA>Hd(_D
ISESR^8f#YRYPR/._.IM=aGcbT+I&.B]R.Pf?\^PQIY0PYZbXT]4C,\[?PLM&21C
V_9MTZU)6MD;Q:8#Od&H_24<&FfSFK7>YI91d?C]VUD,6<SRK9cZWY\G@@A-E>3N
VLb3K_gG5H8cQ=O^94H@\2NO^TBKcbeM8Y>@^f4dA0->7,Y+KI5Nc3ZHF]V[BF,B
,H_N):Ff<1)R:ZNF#b7(X3G&#\Y:aPC[?a#=+Ac>HGJ5-6,I;+CZ.KXY+SFRfK\[
&8T.F\.HF.4+@0N[W&<Rb;[EIcX]GU[(+CH.L26,WaHV&UO@CbUH&T8>S[GJUC1_
HJD&#Rc&USQY8[-@HQaDLX=(7Q[Y)+J.,31D:f80=.Bb)[Hf;^44ecE>/RI/1212
H-NGHM7#&E=UX6Dg/=&He^.GPfPg0^(N(9aO;W4\g8I2>HAbGQ+6MZC=4PM\?E(;
5F81Ia/eW7E^W5:-cE-M=8Y-b8AP41CBFf#9g+-/S+aa2TDK:#(DP63dF+;;D^+6
d2_dB_\=2dO<.bR<444<N@T,WK5F]UO7Z0X.>:bNK+EN>W#9YTV@^f0E-F,LYUY4
1P=6B?,T[_3&HV)PX(NdR;cX=UV<BD/1DdP31<B8CGSR7X0)LRS:DJ,:?TE3NeHR
Ca?\Y0F^U9<.PBfUS(=+:+b7G[I9EGPeA:e5IdO>;Z-=]-YbXd-+eO,RU^;]A:_,
Be+H6#5V0TaPM]dU=4E;TR?Tc25<=T2efe7b)WdbSJ;XS5^QZ/=76+:]X:(<4;]c
2Q?T?16YS+E5VRPf\?:f.U(;/cbHb)\X7T8H#9e)97fR+)[E&549TH0E:0[261g8
b8:6MCbO(;a;I^_c\eSfceAZaP67?Eg/<_@-/J47f\<GWNLE0a[e.Cf.=O5:S1d8
&L_a/\^.13_KSY/W)Q7G=\@afV^c_DO&)1E^TX8-,4N.E>8AK<.ODJ9NKPH/]BWU
I9[WaEIBJdM>(gf:#B:8^<NA)3H?1O9XLN+V[2#JETBc^+PAI&PB<7SZ)NS75aX8
K]\d&R.]XeQY>X9@O9&\?NSR;SfDe][^IK-K&F-,9^7D^21\@KQW?D[CBLKCSaM&
R3<M;gI_Z/0:]GbAH82DdLP.)I73D0e66e+KT2_FYE:;H@,HPO[(-6\Qg&.BNWLF
NWMLOC@Ze:E&_[..2d6c]8>]&?Qa@S4a9afC@R8D@RRAYOR(RL.=/,3gAIW[PaX8
I:2P?EIUT100-LF_,QUHcX;D=a[V@O\SWdMMLd?_P)1EB.4AEa#4TbLgaD9?9S/U
LaF&gJ)NY<WF_@:fMGD=e7I&##81V.?1P59XBU.gL.6;USA_MB7A\B[c6a@+G=g]
68>^gE;;e:-/OE<Z<?B;G&H+FN3SX+T[>6^2CVId@P.D>V)K:Z&J3<^N?,0[PL)/
b#XA9Ub980cbffQV@aZZ0dW/0g.=XdY)3]_1EI4.BVCHBO+Qe(112X8[O1?[c(/O
;f1>;G=<L4Sf&<&?.L2V9a[870BHU]eMY)=71=a+IIU69>(#OP->K[GZGZ5N-Z;B
)a]>GX.;ANB;[Wc;T.cAK<2Kg2CVJJ^:R&I?QT-0Y<\90]8Ycc3MaI:\GE@2,C)U
L@D8S6:P)S]eIEId-/bW<(DJY;BKWPLF5gd9-<?Ze/?4U?Ad:f+&QCM6TC0WBdY/
4O[&@R76QT@\])(ZCQ>YPafRAYSO@_O@)TDPed,U/68OL>Xg:/)1^4^[gB7VIgRA
JAf^YM)YA[,9ESMK]J3b-6R9R)#ZCI.+RRE&)>.d2HD@)fF5^=<gbII.DKCdSUPR
VQ2g)^CcO5Qd-M-8QTSD0(_E8Wd_4c\FVD_[]cUP?IU@Z;42[J0U0D)82UGA.F::
D.^,Kg(E+(TL9IITXcG^^[E(8:A[)T=Kb\QGA6&=(5eWB1Ud8<\:6ZNUX<\f0<WD
E,#8UN>;4QN;,)?IH&E/9WeRCN9OWJ0Rg\I^.2E..CB#LCO<:<I&WUZbR#W/F[E9
&J?RS09N[&aXRe[VCY.;b\TdV5R^<N6Q78>>Ida;/Y:C#;K)9dVKF;&I#J2D2Rb&
:(K(;&2H(YF(H,aI51/CKM=A;aRBB5?#[#@_./FbO24#fAO.T02&O/?WDdQfBT4a
(&(5FaJ;ZID90LA\QA/bQcG46fIV;0COKXIE[#NAW/[FTAEERR:M?NZad.I)FfA>
=7F7B0gg0<BK_&^.1^e0Y:AH>IaZ.3XE3PGB<d0]dRFQ8]WP^UQ45+dY.?H]KTCJ
gCHGA;MdO&FSf>HA_23O7D>Yd<S3:GZBG96WUGe9XX^dAKVXKDY,g]fe6FFB#Jg+
R:/4.[=6KB3V3#f^M7BcE)1CZDL557ff?MI\AN8eA-H0F3U?d,.GMgOZ<KJ.]XL&
U;5f<DI#?EK3g?G=GEYIg?NF2e7e]8a+ZXO62&VH?+PX:IEeRLSBeS@BFLZPYW?3
H5d5+XBMUR=@aUSMTMe?/(^>#BF/]e#VL:.HZ\7G3c:F.4:/-(9?BSRGF(;#/S^0
Yb.F;J^RR1SdY-KENE:D2>HJf+K(<TDC?FE]7Z;_3K1ZRHW&R.B#9.&5+R[V5#a;
?[((c:T#1W=1PYAeUE^7.;7P+2L3K([&O979^)9dQ>++J+eIUW,<8CI,0#GEG?1[
#N5S.FBX.@1OaAJ)BMKRHZ33.7VOD2B]Tg\DJC:-FB#234F+eF2TS7AAbe4>P^OY
D:cZ^b>/AURW#FPQ+/J.,bXXgPRXe&b<81g+)^JK,Q117ebXAWQ@E23UUNL:U#4X
YWGMaX1CW_^XQVR\B])ZA+AXMbHbBN./U^5B,6BEbb7ET^f0/[06gHY5Vb@T0G-F
X@0ZKYGNc)UOBc-<L\0aHY5\^f;#d78D2:12:?1ZB9FO+3E/.TD18()1,Oea8)1L
#)5+C,<B(45SHeg4=FaSG,N/)=E#Ve_HObW1\BPHULVEUF_FJ,:8^)KCL9NQU]KO
0G_aM/#8U#S>S4edeXQ7//daQ9,Vg9R+A.K4>Q::43GS1VK&^/E<6:8\>E\(JTJC
SCZN:T&&MO.WP2GWX:?^JEG4G/g/_>7)(RGFF4<:S.FT:__WNC4D&3CM7WGI>VS+
/.M?]2EGg6C#X2ITB9fQ:fYG?RFU]Ie/RfJ\09EY\3R#ZY^G;;(#ZJ#KBJ<,gVdG
SXI+O;M>=>WPHHDTQ840Y,c-IB,[)I#(?LBHKc4@H)MEKZ876D34aU46-g9b;@5R
1UJTL:RE_d#>R\3+>)C<fC^CG3G6/-T4T_48-f)Y2gT#,&#I+3^_;S)]Efc\)W-I
21+M&)1d&@CDg@Y,F&8g(9aV<##)8b#,20&54La&=cPK.RB7-<BU11H/[)M(bN7B
2U1O325<PE(V[\GgHXVKW1-eHJE9/X?=NJ9[fM(?65.CVOKQL48JQfSMeU6E07>#
B&L->L=&T]ca[d><AS[?5R(MPI07]:>],&\\J)?(/.Nd1-e-fLY^SS,G(H,\bNSE
,]METf@],?d-2f&.Ia<F0\&)Y4ZGSTC3f\#6(VUaK3QC,E4AaRg#c])cZaf8_fU(
J;7L>\gQ6+DOe2^EO;Eb>]<R@^D1Ka[3Gae[>4^cI8U7#0:aWHbBONDY>-/S5RPG
S.IJ^E?;LDTeIYO<L@(K5R,=e91#Kf.MG:X)2HVF-NI:K;gNMHEd&AS6MQ]2M>=e
(T/XKJfMH9H-OMY@=IQMSH0E<45\VAJf\C6bJ[fa+@U<8268)YYa]9ASIHYL,1O+
F9REaATO\d<a66Q>YJ@ZVW/.4A.d_0@G-I;e/b=3ffW-]AFg0Mfec7ML]cMFXb_X
1:Z.VG2>BUEX/<YE+E?LXRNZA(,g-L+1#:38SBKPc1g&-Cg;SLDAJHO[+7-5HET#
6f]d4aBWL0C,43[5WeRS716<JETf9N)S1-F=QgbOD5Ka?6]3C=8/6WF@5S2XLEVL
D@AA/dR(-61QD<c<FU[1=V/^R\WA9[?8c,^e4,e^WV()Z.^6OEJM#EUPDA^Q.Z^d
LKgKc_0?IffM16KUbf+(32c&b54X_Oe90>]]+KZ^S(@.<\CQ_M^:9SC_>^0JJ,KC
5H^d-ST]+TYIJd/^)GbcO9WX.a][LY#YTL@YQ59Wg._[DdD2<H>C;@U\M8JA;\-X
9=E@gQ+]HJ?2YaE]H-&OH\>M/T[(49RHL1/,7>T=4P&^[cJdIcQW@^=eG@U^<P.c
Y#EE&@6-g#Wa\\C@W5Q<TE&A<d\WJeG<)TFfB>4MgFPCCK8\\@/0ZRK,b8?a2A/D
(V;_70J#gR6?S)a9LUd3dW:3\D]Y.\I]e.O;AIR_8.(WKQ)L981\,c4AdAM^WKab
ZRc]2+.2H:aJGH09Y(dR@?(PZ)E?:4\2\NI8A#;[JXF_#R7PQcIVUQ]V#SI3B_);
(T4QU91FB&K)eABHR>bAIP?62K>(a04?c\5TQS^YRbM7dLW+,b(3;#3K#PJ,0/V_
2EKQNOd>MNPJe&VX046JX2a1V?G)T^G&2EI;e,E9D1QZ4<P0,O??1N+KJMReG9cX
a?_Y[S4X2Lb8aYC8/6V?g^@aFS46F6/=3->_00-2T[UL1Y>YW@2@2^M,UIO-8f=6
U)3+-+8#=[d;fga^FcY3(g&UC@+3eJRHId0_H=^V745F_WJcdH-d+V<CDNb_ABR:
>>BODDBF,dfM4)OE83])@WJ.Ja=XG_\FbbNP-A&6512TF9:OD4C<:T465L?CXO95
8U5LcaI9Ug3?^,Bf-/4L3][++C6<(4<4G^;)4UT0.8JBU[.I?#V4gY5a0Q+>4G:)
.E_XKg2QdV\=AX#+)[3@+I47-?PS<&JR3S3CV&[[BfYHb-)Ra1Tg5CJXT(=Z+&DD
bbNWIcFYQe1a))9C]51#AdMD7-8.?+#6bb8CW,8=d-)G39U5L#?([WFG@8)EI<)O
T)S5R(76#Z[+_XW@bBPHff39.@N[#B-[&#,Y^JM;=+a?_HH>a5YMEDW]F;BG_F./
LCO]aUOeT(#LgVR-Kbb@R#/S0ZF25^4LDdFD_>PWL>?)AG706.T@I2D:C/g5S,&3
+-a8G+PdOFd/YFR/0,7Z#JV,):EXUaZJ=bARe.2@PUE,cK=>GB;2#JYYW7C,\W(U
(VO/Z15Af#><H3385=XZ:+)_TPC[gFaBIZ[6\=^3DL6[7AcXB^X@fG4I7?96EFW&
>#?7OA4FPA[Z?U>.K_I@K/&Z-ebI)YD25IAQ_ZV3.^_AE9U1(U.d,3O;/_.eZ/dg
V>.ZH1=KBMK?03-UF+?Y.(c)c03_V\XUS&OI,^V07Z@6S\,c[4aL5VIg^S.@)^<9
O8OPSDO0P&]6RaTaY:aP=_\)17-d_+T(D1(OWbFW8IB2^>;X;TCV\g]O+5#6+=>>
6YYDJ?,1Z6G=Q3RfT\&KU]7f;CP@NHAed[H_I,3VD,DFUD+NR0DLS)Jb0-JXJg7d
fOSe;=D@:eSd8(8_7;SGJc3PT[b93cc[)V+=aH2>ELU^VR):D#F2Ng]#:OQW/VCa
W/;]76\(/A4BOdU2NYCPdd#,?e@T/KO0UfQGW76L^<K:IeI2/[g^0AN1;@YbI6O)
;^?b(8.AR\>K&X^e_SA7S1-d&=IdG,WO:T;eIW@?)?bB[JRD43?:[16+7cAH1eEN
&P5BQ/S&fQA=LcL]ga9RG^)GTfC\&>N#R?^.GC^XU\HU;9P84I[A3FXIS/5G6&4/
K6\Mb6)LP:_#F4FA?)XYKa[^2)H4ZKJ@X=\DK80\,#;AXBI^#@9(0(_4^9E5PNSU
JO2CLD?Oc0CO.8f2<ZX1,eYMfI)_JXAdF,f:+Cd0;DC]SC2ZK7I7I1>&c<+[X;KO
A_SKM^3C++T/1FW#K,\\PMSXC#)cIS5]:XW3@&XD_7(B.UeL]RC5c83.fFRbgV@g
[TY[e6@\?30@O[S,MVB+e.;FTCZZ2Meg/\Nd-IHC44ae9gHD8=&>6KQ6BbX#6X2e
0P18?3:T_=6g>X6AR=:67Q[>\EY,\]B0J5NO(GH[(?9_&KHNbN;Y6WJTG8-G+aZ(
E_TLGT>G1ZfQNOR/=W)<65DEd?P/MCd)UB6GCV+d2IUMeF:K48U?_]IG)#^#3&1Z
)=fP1WK,066Vb.XA2\+\:NBP3H4[c@E;=7VdK+OAHPBaI8Z66cO;cHNb&[RR2gSg
WEN<[?3Z,N_FC4REWIfCNO#@Gd;?+E\N:ZPc9N]<@D]aV?;aT8)?C7[<.;MT1LEO
K:[^2(C(+U?fZKWML8#D4B&g5Z9Fb9+.25,7KGLd774908ACW+1J4]&g.?Q9&\\R
&Of@[EB5)L^]0G0CAIS;O+@[<KA=PAY5T^+Z,@,P:adOPfV\Z_:^;V@JF)[c>#:]
=fGFF<H==\EBEKN01;.ZJ.We>=gFT:Gbc7>9_\ZX[WZC(,TE;.^(<EO<NI^-3?7f
-:;4E>;1A2Y&<18IgP3/32^J<_UXH40SIEdFe\0LV^a3-d>Fe0bJ=@-L>eJG:Y]H
K@,1#H.7CU8K8cP=+Q4]-7a?]#fUPDZHU+-)ESEa4<86.(B8LcIQBc_1TCXOP[Y&
2][=]E46(P^\6IM?6NV^JKN?[2+P3@/-UKOYHc/P?6U)I=DXdJ0>bfT7Y7I0_OBO
c7NBZaJ_(CC3+UWAa,E<\@4PgD0/O+e[GIa1:J0IPQ557NY=#+B#8e?H(aBTIR\9
]0UZ;?&YTY)3aa8.KC?[g_DL5@5S7/NNC]QCN+209S</Ufb,F0O@Xd<^a1_:Z9WQ
J[+21fZWaYeZ<0ef3+Q7X^-FT^EEGB(H=?P9F+,A8OPHSGW-eB2[K#?&(/0?K6<g
N,M/]L@AS0;Og+HZJUJ\9)-F3,[&6AL,\QWc;97XS73R46ZGIVGR[M4#,W\@.[d[
?OL?R[B_1VG?>HH<:^6c]T_+5(Fb.>ZfERTH36CH7LV?I3e=C09LJ?2ZbXe^.OBe
.1#OJ_R>V[S#WJ)2eAZ_9#.:+\-aAQcE+ECY>QD3ZNZZ:<V-[_#@=/K,Ed=<e_W&
0@;-<6DUN^6B,\&7V))e_.;CNUa,+YEE1R;G>LZ#ZgRUR-#J4dV8ZH);CEB.\J?f
=ZN4d5X;GeYNC,ZCYa8-.>[6fbBNJGMF9Q,c5W69<3I;H#b?1?HO_YcQ-?2N^-4=
AOSA/@8G0,+A/A@:LJ:bJ\YRdYe)c;DY93_S:T^&(7R+[)&Y:12Kf&,FdTGB:K76
>AHN_LU02VW[c?7#8b/SS1;G#+MW;\VgEAW&X72=f:UT]C?ZQW&WWA4W1<EJcB^(
6DV5<?BVHY?.efOXXe[W+UCM[)-V>32YM=aM]Ya9D-9G-@UBFFZ@HZd#4+>N:B7E
J8[X_&6Z5XHPgNJgGC=L>#@gIQOT3(@#J#HF=SY;I]6ZXAOMU0((667J^;RO^\2>
7fV&LE&VC8-RIDA+A__\+\UU?QJ.<FJ5ag6_-cE;>310S[^1M\8,P[5;TUIb=(ON
V&a#GKGSSd,6P1BO/X&+Q7LfPeRg[;?ROFS2,+c>Kf3(Cf9#G2;AHVM5:M_AJ#I@
Y167):2L.0EZPS<8>GaYDg]I&YIE/YILKL(A@Beg?UYFe_?2g6DVeRI+3=:gKXgG
#GX+BMf21,M_[d[_J8Z;J;PBLX_I4)[ZbI9?]#7/TE?f0(#CeIY?P)/Ed=M-H^A=
=#6&d,,CLS3UfW4B:YUeK,K[)f_3N>M6=#RTP9UC)&HMFAQ-dP<QL#B-fHJ/4\(@
a]PO17Z75HD2(3WIU06?+4^FNfgSfPYBIDg63LNKI+\]RYJ?L/c8NR@)Q:>>H[96
aCM\-P[8Q#^c68AF1^=S)aDK+:3gQ3X^B<c7@H<?bJRBB7Bc8O]Ca@(+<[>M(A=c
-+=D7.1CC0g)>;UN\C<]MMT.0H@TdDOBA[,I^-2b>XR?13(>:ZLgO^(A0[If4/<G
a\=]L5NeH[cNJ;K10Fc(0D#c#C@#E-]+-R-&;EDWc.,RPcc3-X33VY4Vb=OX]/?C
YXY[4T]MP,_?:X&/J/dS\d^>g[)<fa-#TKX@W8cAJ@F<MR23>)4Z?+FF./L:I+;(
DeJ/<NMXb=V-5K>d]D&gRYR._K?M);X,d)[Lg3<9,8RgAaKX&.XQE))/JELbd[Q?
()=bQ7OR70(JIEW\RAH)[E:UEWBd3gbQX&7BF7WbFFY4YFK@T038fS;G-FM9d,#(
\V&&@]J8@Q6@IQL49<RV6GN_)6P7a>XLLK1K?e@R#]A]P_267VPLNS4R^-c&e-W5
]9V./3SEO84H8718ZUSb_W?af^7W)AcXP.)RK\R/JRfQ@[/])M928gd[+85:P[OT
V^7W9X#<ga>,1P:>UXOP<D2Q31ZXFCgOg>;2FLF^\I;3#+>e?T^Y,Z>67[L2_]gX
0/G<PZX1UV[]EN7WIb;J/XKB+#J:83^>P;2H/5[U=YD;dQ[bO6S;R]F?dY=7LNNO
:gH_RQKUaV8=[GV\NDMIZcNA-QQ]Z3RND=>AT8bIAKa=I[7>J:G1+L:MPCZ+HG?G
@FNc=aRfX),(Ng=CIUI]9M@d/Q^^Se[K\XTPO=.]<:I+:HW-3K]<XIRQ6_YG@Tcd
TIJ^S-]J@WFBXA)B>fV@E8(;B:H)GF]@R(/)PDTKY<+67TR6(L_eC>>E=-CR#1e1
WGDOA;;@>;L;c^7\c([U7NS/FW9#<SQKL6IY:N+E9NBDX_VF2<=7>f7AFNFa(e]<
,6YY_#bb9R0Q#@<]3H/74Te?a-bCHH:D;SBG>-aJ84QXN#R/E;4:YX#O]AUNK3MX
XTSV03/]WSJOQ.Y7@5-C0<-C^-KQ\d^GXF:>]_U81ZgG<\bWY43K89]M_ZGWg>,C
e]FfCSS&2W_0)PL&GU0#dKX.LV^d1ZdLJN3c7,\UZ7PA[VEEI/;59#BJ7aL.P8Pb
IaAK(7LLSAF3bSC5#(-C]&_[acZb-H637UF>Q7(CI1B^=f/ST0BYTQ8\?M:(S8RG
[_NfHgG#b5LRM3JGd7gOSI\g7=V3TB+Pg)V_&&T0\M;#>E5Ng0GER?5_=KQD7EWA
M.3<1@D5]590O;DNg&5cFPReZ^9+/&&?1@BR+MYa8/eHU,9N(^g==O?)/JCbD/g1
;bZK_MLP]\0]FfF41RYf2Mca=Q>#=-e=BG.67_a1GLI8Z]5\F\KG4=FI.8A+B_ES
RHK)-g5#I<5fP.ed(#XJ-_@c]KdKB^W8cD>-]@g;\WD&Ed#KV_;[4:CJ,.e6P+9Q
J@-G.KWS#K<@OM@W-aXf1Ec2JA(g=3E7,#gR/aR-Oc>c&#A@9IJQ+SdV2A0gbaW?
BR((,.8JIS6eT3b6\PS-T8Q#H@3^Wd.1S4:Q8W_JA>A7N.P]aS]O(44Y[^Wg?KR9
R?-#3dM0/08>>EWe9-624/a(GF(KR3>30P@&gb\@ARPTW2fa#]@4L).fNYJU4I.a
fegI4_0Y:gaZ7Va2aA8<U&H)2S@5eEO([WO1D^:TEdG>2QQ7AWdF-5+:B>a=IL4Y
,.aFJC>SE)R#Z0A22.<_f7B(KL)0+SJMdG5cGE,bAgbQbX?F:)D8Gc3X)#BV+@DZ
dIA#D2b3>-\.&^W-&R)3:2@cM8eQbZ#(BdDJP356)a;)UZS8_-fJ/-B/N5KT8BE[
E+\]0<=VS+-.Q.8<\BAR-Ff&=g7#E)4(CYR9T>8R=LZ6)I83\UT<c7aID[WJQ^(Y
6PfH#&>9/,#RcAMQ_-F9Z042b5c;g\f^H=7JBg==#LUeNFC^Og4?0B>@B4Y56Q5.
RCL>6BXPd?<BM3/1\=?;,5_3I+4VMBEB,UK9[7FgdT1N2G\d(afgZ2B_R4?4:(P^
.DNGYU3+[7f,K)&Q7Gg5[CP+(L#QSB+Q-M;Ag=H2PX?U++TC9aMN_f)MA^U>5K@M
TZ[VETaY)<M@Y+]TDUW&CK7W0[X&+J[4ANACD-2TJP7RG_DE,I7>d7,J],1c0KNH
K0S,F>_/AEQ5_/J>YAX.I_&;E>C^M>:ASAHg3QW@UB4<H_?6_dPU(2S5BW^UGd17
>A-G;.LcJLQW^=XT,Eb9c2fdZNRM+118:+S/;@\Q4f<\aBb<0_aBDB?GLL_EGS;O
R_0eY_=8Ha#W:&-eEK7\gWYDP?<_Tc6XB6(FXRg(Q4gW\L4M^M3<;+g+;AKNG4UH
.P>XPY;&M_.=Y<-GMHe[E[60D5/SHDTfST:=KE?H\d/^<P&We0>/G24@2a&9&_\R
.5f[K8)0A>0@bd5)Y5SJ.^+?ML3B4S3I>PFZT)8W<0N:KPg\N/HO16BL6](XN[U7
62U92+5K.NPTLK_)W^;bH87ddS#YfcSK=&X;#\_L5,_Wb;L07-/--+8:JJgZ/F8e
T_Y1d<XUceZ#7a1<FIaef=f<+?f[R20XT;38]@DC5aK49==8:0^g=c]@SQ,<4RaC
PY#<2[F@;RYPRCCODX6f)]9TB>fSR/=7E:d59aQQU<E2:0f?M4\K[B_G)2W<c/G1
M1U=\&7C;XP&E/Q,QS@.,(S#+B5&TNS::]^#61+KJ(Cd=,K_J--59SXH\Gc0e?+N
D]F\,;gea6;Wb(8&gCOLA(cUFEE2X_&2_&D@<\]bATU+b;S_8U<5QDY++=@fQ5XR
D^GgI]G8)B2:M@5R5O84d8B4E]6O[.73/P/cUN&V@4S\@,LJ^H]NV&(B3(X?MB99
H6b?M)Af<LU#8;)L5D]3)[g<85LSL5F55=:@Ke#_-5-+.XUHRW.=4T9C+c8?T.,T
FM,<UOL&49/?@bQ7,OV,>)O/7>MaYYSD2,;L]+cG.Rf[N2Me9:<.,.D&Q>Bg>XJT
-;]M^gU.;4S9C+HI,/4.bF<P.W_g,Q1:\-F8>ZRgQ2f]g/&G)@59(#SNX_(5[#7L
?IUNZQSa]d&_Ic;V;I:(1c(QGBN\9GLK_7:R745N#6YMg1W#\;/f?9K\=H=aLE8#
;(:^OLbB000VF#c)_[-R)#,]K/ZdUFVI@.T4_^O?5ZQf-[YEF)T/O\OK_\3,g:.c
X[2BP^9/T+4d^Pa6QQA.YeVEDg\Z+>K#BE7F^8L-G,Q,ROW]@<Ga/VCJP3&2EX-_
.\?8KX9M]NNcg(+GEUe#VG=ME\NfV=ScPK_.>,>+L?P,SMCV3dEXO5O=+GA50X]<
?0&KG1C)H_PB>3&O0FN<9&.1XDCR^LDA:4Oa=Yf;Q>22XHYRWB[57MCJ@N3W(5DE
F<3H+#[fZU<3&g8V?]VX4D/R/64;T^FF70F:,X5Hf+)6:_(gM:&PZe;F4TfQ+?]I
K>E.P@)2e..N&WMK&N)Z]Z08XN>;T#=KVQE=(e0P9578FXdS19]HGCBS(71-c]6[
94P6e^&;=L=U4FD]2J@=8D16fF>f_TMFGF_C6f4A3/c2_\Y0D)QR\dKe2-X[RT_d
X]3H(]_d#@[J11>d1,ZN-THBJ24.aVI^)PaLfEY>1gc-,AUeBOXQ>7bQgR-YDaeY
B:&+&TY.bSJW1_dV,S,UFL_1d]fI-G3MQ22+=A2]&M7N33#00K5\4+.9?.b;\S9]
1^N-:e8#OVDY-BX-/@O+.+#XQZgTY:H8[&F6)Y3CXYPa^f6gG&0P9U5TA[PQ==FS
e?S081=381;[Tag)5aE[^g:[@b>4b/_b=JN_<5AWSc9;dQLIL4YL9:QTgb5#Z9=&
;eJ5_BPQB:+\US.89+11A\7fJ+.E4OARCS_OE1GZ[9[]3\gW=.I<](D?[EO8cF3A
8#:WE7CR_d[5EO66/W2R?McH3RaEIRNMC-8,:\-e+4BNf^I0(KHN#TY19)cUL:2H
Ge<D0?(b,(F-.?/^cMC??;O1/9H(+9&GY>9O+A5Y?bc&3L\JT\6[L\TPMRa[>Z/7
XAHT;N\HDeDD4VUgZSZb=K/a5H5T6e[WP7BN@]V5b7V<Fd5?LgdcH\C#<^EagQL^
.7fUU_JRg0ZT3V7;SJf:Nd1D)g[fA:F.Pe6#8S1FF8Lg[<Y7NOE5[L@>DWe:GKX9
JGf&^SZ#&UXLUgB0;)\-T/ZKLI9Jg=VWfC?d^1^aA1FbEZ/8/T>,0=\LGYE<1W7J
9?=-1ZN(@(1(,##cR.P6&,?P;0CX.4CW))K+Z6<BK.R/VH+J\^-R.YJ__X<54bVS
/aE+c&]+N\5E1_J6d#A>,9#c\(g,XMNY:G[L.;d,/1fU3Gf?Q(2])Y1>61Lf2Hf^
&_ZXf(d&Fb74/Z&U@7Jg5@UYE:HXNIPK3)V975G0Y[f=4\QLcJa9=fPWc&gDVXQ8
W\@^Vac9652Bc]\)(WX+#VdYMNXJgJMI8P-F+<G0f&WZ#b[<_OH4EOM:^OOb>I1)
47W][1bD^G&E\NR;QJPP>^eJA6Db-4T).CB+?58Z4?^NM5I3BbMe/573DK)\>7KW
cX-53]MSWHH;^e.4#caR7(Hd40O3Va,-bY>\HdWM-[NdM+JB+5_VM]USN1cNdgAT
U/F>,eM\N@+,bb)6g9LMDG)7KM?,W9(D2IJcR8NV5LQ#UM.R4CAZ\]dZL86NNdK6
]W^-F90D0&N,9#U909MXX?aOQV#].9XVCSK.&BBKNANUWL:^G_BbU(X5DAI#S@DH
DG69cgcc./68VMUQ#E8A(36;c@WZL0AbJC:9SP(da71HZ8(BK70@^Qc4.U(e:>FS
V/MNRH8LY:K6g)^g.BIP,e#3GbT^;3J-(@[V\VHI@@+5UTV[(ILd@22&CGP^cK#a
>R)V-X<(48Z0P=U_YU(Q]dJ5GK>EG\X\T^\:b<8SCLL@?7)08-EH#6J9Xf_#ZGG>
fZ^,J)V@F[+#&@FB:P,076\+/R4]Lg.3Q3&D22N)6H^BEM7=>HE2@(9D&2)Q3IVG
8/>5R]=+&99gZY+:67bg]\X6F/3F>H0FK))\_fgTd^-Pe[-^_CF5MBBZRKXa&QaP
XPdfZ&Gb0+)SRP-@75G6ZMd2WB4]P(6M=YeJ+bPB#&LcX&;eaF02fC4N6.97)142
b4P@P?.B5MfO);3UXJB^;6#ARb6c0C.VB++FOZCA7e8X_J21M+;&&R:PBc8,fA7G
,gVW@6)2NbQ99;),,gF-9XNIdRR1Yc]5WGgP8RgK[K2\A5HJCf;d05PHa36K9Xa9
XC,,X@(A&V<N;F9e3&DLR[9RXSX9fc0GgL)/W\A9K@;)2N\9]fE(@Y?c+C/WY(:B
6X[6H7AD5]OY,7H.O1NR>TB;\N)JL9KS[CARG0)]_Y;eSdX-;]SML)Ec];17T1X1
HI9)Ua&Y_NE@8_A+#A.:c5)AE,MLZK4:F0Y-J>)?FWD4G@gg?;b1&,cdFHTL_8ET
fMY6,R]?^fH/A2#e6_176-cE&/&/B#Y;J]-)9FHb3fUe/,+MJK8]Q;GW)T_I7cES
F/G7d=0QYe&9)abFbTPVdbfZD6I5A--#->NO\fB#U8,fV9(QX+0Z)WE.dc[X?=+9
L&Pa+4BWVF^;3>/W,ea-8a+51MBG/^&KLLEfg30=g;NW<K]XPbd27S,eeKI,([(,
6_M37IUB<e@<>ARE?a+:N(A\8L]Y,Z]T3L(U.=ZR-IPZQ7CWOP1OKM[dTS:[,Y8J
W_B(EWWCB[e3DeZK=U-fUcM^C+C(A+F_dBUCF1N\39,ID#(K#HT<:]-EJ]4-EJe4
GX]8WDaJfC;#/+AE\7?K?CgB/[^e,5J;LbW/K[0CFQ^MFET:M//bE@IY:0.M,JGd
cHR@@&QdfF9Y2V0/59aEUDa?;B5gYF^R<TPcRR]a\GA\RO@UW23MaZ3(gMM;<Bfb
&#.6?,3aTeS.AF:eKT/\/=gV7-QRM7^BE;GD_UD@VB89.L.,Bd+>^=D&:I_g8(V.
5XaONW-(;ae:XO<VQb@YA@UYAL0_1K-6^AOdRA<fG0PSBcgHD9FB4b-P-;T4GPOT
2>K-:H,A@3G_c]MT?8a:U.?CQ;E9:(\EZgPKU]<K0?/.EO^@]-gK3a#FTbMSC<HM
?OM5c+g(O.CK>E4ZQVed7ZN9[C,DP=M?6Nffc+ICaf=??35^6,1]TCA)OF+7^]fL
.<ZU^J#BeBFY->a4cD9,#5/>fNa0C\0+X/cJM4d>0cN41gRCd36/UEEKV)BK]LD7
c9Z(6H(([3XD8b7b2e._D[9:HA73CL077,bFN@#G(L+>._fZS5.FFQMdL?U\,SWA
g9([fLbC5a+:.PdE[@?R5N@73<Sa3QKFK7\9eMe:c?&.e3bg;?]VG_R\7LaJAM@c
TXHILO(G&5LKXV5I-Mg/NTQ^K?3@e,B0K0ZNOI1=8/,^[eL4WI6=,d6Zf89N,\F<
VRVW2b[2bPd7IZO#KC7U^c^MWHFW7E,SNfWY1ANB37g;WV??bMRaE<3-deIH;E^9
5Z:+-X,g9,UOX5(P&=VU+WL>?P1T<;5dYBX^012Te2gT6e#3cV98-1+-=gT\Zb_d
f6[OX0^K&K8,R,:=7c[Q(88,_].9PG=_T)Gd3R52LP9\Kb^Oefb/&ZHUNX1O7V>&
c+fe+D,EZ0:&>(6d##>8ZJ>b/_ZGSW&Sb>W-F+I^DX@MbWYcHF-JYUP/B1397&CN
8=UX#JC[EC;]71B.<5HBDXec;Z0Z;HWQU9fZGQ)cNM@cWEdGccB\O&Q:+[M=GaT[
8b,P=6-a,^Pg+HQ5-EWN\CO1+VO+S_C1XYP)\MNQ[/acSB7=fERR.TQaRISgUJ_S
Q/f@1CZeDQE3bVW?gDWG/agI3XOXLf7;L8J&.278[#=1.1.?G_dI\_4g3Ye20JY\
W&XZ^ZZ5L\efCEVO4D:0e0X]Y[O2W(U1O\V/(bgMaKZ.<-9fTN^)/MJdY3.C1Y5R
CV9X)TQGe^W.?aTgD_3/#S&L.XS8Q97f4?G?dB0[\(+.4/:/XVSU+@KVb#R5S=Y3
AN=2\T]Rg_8^Ra^86J-#gE=GK4G2d;4N8;?3;?LIeQTI4/ggVV2cV]TfDF8Y<.N1
aL/eLG[I@Id&U1T&,-3YD?58JOHX[\#I>A50LL/RBA&1dP7C3XKX\NPIU]eAQa9,
a)GECKC:K^F^7Z7]b-,6ZCPRO:N/0S=OA<X9+A[gT,D9TgE/:WPd^07,BG@9L9_O
ZV2ESI]<e,:_D.K+G@J<-Y0#=CA_A\eN;=J?BH=8RbA4WcI^?ND?<R,8QEN8+,?-
P<CfAH3G2S7R^E4bTDG8gP\Gd@@@AOG/Jb?LQ&,:I-,KO3X0U2#REVCK)8TRO5M=
;4[YHf1T/7O(;6;3,f&8TOf^cMMVN-<a<JEd-WNYFcVTg;NN&OQCVPMW]ZSO3f5F
\J9JN+P=N8W=/KOQ8<aTg_>PdBNfJ]=WO5GP:A\XA?1=;H\8?VZ:VUBAINg-_gZa
YD1@LMOZ)(RBGJ7QdS[LS]N5:\QODOKW80:C4+#IV;=e)IO7WXJB<dI\)191L3RZ
,^SNZSK7Db+(b7QZER3L/5EYIYD.Z^CaR1B1CLQ@f55&Xe/fFDJcJ.2/79TFL,U\
OP>5W0OG2N3W]C=RU(.0_HOX:_U[HaWbMd9V8NJR72F2RMXb0:-JN(36R3YERdcZ
/G-fMPRI5[)H&?.T9=#W(d]&@LO0VVUAJ=g/NLfbCe8M=3@,X+bS?gI.S0M\@@O=
)-(a;((6fJ[\F,[c[#QM;(UbP;^76HR_,8>V=I6/f+aU6TD34#aK4]142SL4G<3^
0V6I9MTUV_F1WgG:B(GJdJ9A#KUAC6.PRCJ?FYBHLL;g:L[4cA7BY32C=<gefQe8
_@+1H_c+)7^acgLR</IT5B@beA9VgUBg/0Oc:^/1LIaQP_(0c3HbP<:d#PXBIf;L
WbIMfHeFKbJaI0W78+<BM6fA:;dFRfU<=XTU,bV@SUNW-Y3.S;6C(A0#;Q;SHPVV
V:cV6fMM\48AeBJQgRR7E?^C[M@=dBUc4eV<H\-@KC3MgJHX#b-&K2:O)B4V4:CC
K<@d:C<O_\3/P#)agQ(#&7?2@-^Og6)O96(S=;;-P;+-MHJ:[55B\5@;=G9B59aM
K.9/427=7UVZMYH3bQMU?>_bZ4_^/G.<[;4B-TP9CH3Ce:E39Re)b;D5A.52L=EC
Y4=7cV+X(2L@NLF#7c+N2C7-;Z/XO=#]4U5DQ6[PL^WYd8X3H</d-4TC]f6BMY-3
_7dMPL0/F[TJ8B;]IeAY)K52T62/S_Id)Z@e,?DdSM&QY2QTE7>Y<C&RE@FL&YQa
=c3@-LI/<5.DeQ9.1S)#K\<PRU6:&5bPJ0W@@;]CH-&NCa<g#deZ-;6G4gg-MG&6
d<9(H/VOHKAWP?G0O94S;bUAM0#U?a&8Tf&Wb6MTc\cK\XbXaK#>?FYFg_^@;\;U
>aKP__1+)(#V5IbIb<0ZdQS.<P/630H?F1Y@A078@Z<7<EJ@_7;F;KQ>#7,egfFS
&Lg@:@bHQ0GX=-^PAW@KeAbd],]Z->.,ced>=S1O1dP_Z[Zb<#DX=Q06g>>fJPI^
=/&BXVb9<]C2a3PQV;W(gW3Pc-Z?2POPGM5J58^f7(^g3<)80\LG?;B<Jb+bH8R1
/4AXC&bWIc@1LF#@G27A<F:XA_A:8W3+AVM0RE9FI593A>dB@G4K.ZR_U9XdGgcD
89JZgc,:.a\-+F:_@C.e)d+5B;:_I,ON/;<b#_L>Y-^)@/#43dT#DPfXP&#<VLY2
AV[=.4Ye@\BITA:FP[L/SIOf.I84K\-9K6)<,3FBeYJFc5acWW,A],M_VKg]7b^1
&E</)P7a-bS1?<Y<Q)0\_\N<FGX[SICMH9SCf7[]TIdC[/?[&])Q;Q/6F#?]7_4+
cU>=,7S7)LSM:KQN+be)Z_=,.1e-SF3ZbJ[^L2=PB=XE>LWaQ>eIe9:e<,g\@^KT
DM>64Je5^LMZG+O:T)9X[L++;7K?A:G@BV^Z41S]-?C\R1R<(YW?F]_<O50K8?63
O>d@f3>?.S[XP^UId?VHOLg^5W3RP[V1;Y-^4),/8L[CfWWZD[YE7^+&<POOM2VC
D(I9^@Ma>eZ<a[X\_5E:4/B]/2J>708_g)?2::CZSBPO/M5@OY\f42#7c@P=F>fW
eYZ.c_G=D6&614DK6W=/X.Y5>SV-D9<W)1.=bZ+<:d_JE+4SS@LT<-TJZHb#@/8-
U?,cER4Ga<&BTMgd>SN&2JH,QU:#0XU?3NGXAJ5RCd?[0==P.Cb^DXU\,d0;Q.4V
BS22+GHJa^^U:[&V2&FG\;]?W_AP5AXa)PO+=Vc[NbE^_]\R-[agdf1R^I3P,a6g
__475N<7)PJ(TJbg]I[#O6fDg8bN1Y:\3C.=efC]([7EK5eDfcBg0Z08WLU7CFB_
2(VSG5?K;gO]Yg4&=FT<^6-#MR;U7A_f-AX-Xb()2DO;W[aQXLOf<AN6OMW>.CUd
.LZ&WJ<#2S93K0Y8VD3\8C^#d@[=I33]1a3V,\^A]d=]4XSP;>W8S.L2PHJLF0;^
fdY:V)BSFW4/-a];KA]Q&(UL/0DG+9S>-f&;(Q8RC1=ONfCG7d=-D^O:2M-0IeM\
T]\44;)LB[aR>L+_5JAQd,8^T>87[>+HD1b2_9):_46<V64AQBGX6LICTC[#P;;\
;/EZg^[+64/aU:AO[d<^]-WEREPTX4FI4F;UJc>fPPJOf3_=a:@#5;b1)TCP35H5
,2&3)1R57=GZ8/]gRc9^0>:QOfWY9=B7X-@9QQJWF_C_F3Gg?TPWZBT[V&a(cS_,
CQ3S0V\QcC59c)55bKFg:5K7Y>K_aZZBeWVG@/L@J_\(^Pb@7G6ad8(&ZK.S9eS0
L#^?<S>.TK3FW4@4ff^Hd)AS?H/L^;\.baJBD5b9aP\9^Z>(@GT=,&D@R?LFD\E^
8056]6(ID<?Md)9MfOG40;Z_GWVb())V\ZX1NET:IJVC5G<;<LD5M<7+^#eUgZ8-
3Y#2Rb1e/?/JfQ;BfRS/aC6G@M/RLIA1M#aG((,=PD[CEV7a-ce9KReeV_X,-N34
)XUJM7eB5dS7WT5P1Q<b]5=[GNC8^:1?&QVQc)(I7&DD6)?_(TfWcXe9AX(Z>=e[
_gTHZB\28SX9V;<>OUcP^#fBQgM9Y@3#DZ2].&;,Q=XOb;HAYTY)EH\/R^Y(d?P6
@_Mg;EZ>PaeH.8_O/]d:@[cO4B9E0.R<gBQ8_FQO>]J1>Y<ASNP/-V9+(2FN)dJZ
_4=PTX5Y/DNc246+IAT@-I0:,=a41,_HDPDaQa;_>>35TM47DR<#B2^J(_5=R#dB
.&==4)YZ-@D_Q-A57gEX)JTVb-_6gM/(-A2-B;+3\W0I<WaBI]M\A^fZ+BZ?[M,C
F:.Z@I@[-c?SYO+S5J]eF\;&L)>\N<-9)OOg2gIGea^(;O5K[#)SJAgEL9P(8bCQ
#g&O_F</<T6DDDde7,=/RT4\+[\2[[TS+,>]UWd7B+M1NZXDb&&JggF32f>>C.d_
cXF=b8ge5E\HO+YFHNdJZY>4C=)G2;?P.,/F:4ML/FMHP<[G8A2T[Xg#JC.UY4G,
_#5L32;K7UL&A.@20U?4+,)d>XA,6B>W3./CNA)/\?Q5@9X(=40YRRdG=8?45b+0
#DN0YPM8#O74MVCZJ)<fYN]Pf@4[XH&b1.\&d.C^fB?DX>dH4O2/aA5Ff/8E0CYd
;eR?dV2gRK3GF.G-:(_eSU)(O\8[66=I@[E70;@69?2d<5DL.6Q9G:Kc/Fe4R62U
45AJG=.\7XK=3YRa#(6dL#7(f4V&1aBME[S9S:8V9Q9,:+9dU<\Ud9G?I+.D.]c(
)7;<bFeX[-5bCCVYG45]G,17NJKWg691X@P5RIJ+QL]Q@4TG.C6S+c[>YEU2C69c
fKSeR).b2c#M7?MB<5GYD>?2e.=.Mf-(D=UJ[A,c?\HR[VS[D9KB\8KHZD7/Z?dV
U.FJ_eTA^Ifg_]^LMKB;3c#>L0QgaQ-6J:aFfgVZ&/.E[,W3^^CJ)Y23@;^WCMJ_
QdP5)05.dVJdS?W3+ER]c=c-K^/#G)2W)M-8Td0HG#_3->RZ_)BV(fcd7_&fCg3J
TKC/[)IB.c>Q3fg>VJL0BVA6c#TQ&?f]Z3T?,;@TaGAeZ#;19-&]ZIM9Gbf2K[>9
)[fA=EIL-;.^6J?JGE>:Gg@::]3.1M8<\1BC61&5_K3g:[L\[+@N,ZOIc+S>WA6M
(M<g6\]19_272/LJ&K9,F9;-&O-R[GD4OQYUT2.?[=?60EKRJIZ&YZZ4&=HFAV33
^(CU:QCOf4)@R#c8<1YbMNZQ/\IF9#b:9\5gU]PcHKMDX\MM85>-H?J)=SCZVf/f
0>IT)D<GIY06=8X=fZ\FHK4;/[dWK1(aQWd(1]a48ZAW068^S-&(=cYb(c3\YHHI
4]V8+N^J;K;#\D<9/40C<)S+#U?ONCD:U9D)9I6Z1N2EWSQB0F7-FTN<S\g.gfSB
QB+7Q09AVCL@DAJSB?V>+<PE5+WdS0>KDBLBB3MH6U\<+ED?[J10346:1N<MDYEd
(>f#]1dTM[Y88[5N<A>Z+X]-J4>638^(1VP,fYY8SNTcXDGSd(O,<;5AZ;RCdbb\
2+I&5KeF]IE@>-5EgY6=]gS^Na1g?(Qe&&?DOe9aEeJWBY<ca-?^D4Nc[a=-)\(R
X)C+I5ZH2RMC_e<S-2S2?g4DV\4S\91a90KD4^\fCFgcOTYGD;]UdCNAP/R[GPZF
ZHGd\A[5)g-bSGH5a&E>_<]GNf16fObaS/G^@;#T3+1[(b0,@X[B^:N?>]80]);T
5\X9HUV8@H3^0c^YO:f5-MFLY,_.a:6[U&BG-XJ&7Q6+dDARHfEaG?Sf9N&9g#QA
#A.[-NaJFJfDKU&4AO4+DM2(;.cU)5FS/BJ<WfSR(U_/M>OU8V37;OfI.A8:c[IQ
:I9O??]d<_&RVW[P,SWA/FW:KBI1B4@4NI<XcH.>ZKDJMYQQ@R7\:0.9<<Ae@,YX
?>D7)Z9<RZd@gHT9N>)].X3\dFe2AcEbgQ0W5[2,G::C>FC]F64GbE[e=RF>P[XE
F-/=LF]J7O(=N)@fH7aXXM60@L(S-9_8KPM#@:B?3B:WEeE[R_KDR<KfP\5c8<)2
4<7?KN4+[G3K@3N923-.A>1T0J/\.;B(&&Bc09eQ4>I(E+6ZQ>@5@K1&I&[/:E&L
;WaE-ef?(5:b([MPVPAV.4K/Ie?ZW&S[T4&YX=Dg/K4B_C6WZ(@OZ;65TgS&RTE:
63LPKZa-)+:N#RW>J,#=M+K>Y::2F-#._aEQg;YA&_[(F,PPL)URQ&@g:dYCS1<T
BISLaB5^6USX@XIdaO,+dXOU5W_S9c26D1+J5X>LQ]A(4fWE\Z-+LDA>gAYDd1b/
9J:DWZ4^ENI_DT@=&Oa)T,/I6R:ec>c_OGNC(Y2(=1L+g6M6Y^RV+F/ccgDfCG&Q
?afGF\bJHN)bM8IY9<bVK&WWLV.ZGTE=Gb39&>;ILQT;a^g1=[T39Og8?4FMZF+:
PR,PC\bD?>HZPE#Q,d?e_;TWfABGa?gHI?Y7;[UTFO3T2KF(Q0ZNb6]4>R=)=f.Q
X;IA<b@dK^E@^e?#BQg;#+@LOJ>Hf)=D0^+Zg=IBd/P-ESdP+Nb,:0-?\99S6TcS
0#39H-ReMD<<^V@I0EB2J3^ZM=X#688&V,947fO/c)-)FF6FU1WOM3TF-M:06RBL
]BDBX;N+U(2/aDegLe=ZZ2(V@fVJGZL8GF)7dJ#^@:^F\ZEKOA.c#8EU(AW/>g?Z
44C?]S1_JYSa(b&(ab]WeXOGH[eJUL46ZMfccL^4J?3FF0N#:O@+AEG\+FC>AF3:
Y^=:A(4EE;[4N,KVP84>Vc;:6A#QZ@#=Gg#:FFY8(DDLfN?+RY/GBB;5cGW3C7HC
K;023<PYa]5TB<S56-HW]LbI63fU=0=fG_H1/0;B2KRdH/7DD10\=;S4Z#<A8X)T
>T+5F-aEP1+<XR)9^be26TaZKR:FQ)T)bNKLR93IINQ@+.8_1T:cW8U;:^)8I:HO
W:\PW2I3_.02G;5C;EE&Q6>UI)aS?,(HAO@7]+I[IGQD]\B21cgDbGI64<G[N2J2
D3UZ==)81K.RJW3?\1dg3d2MeQJ///=g><0FAS+)f(DBG,C7&#D3B=S>ZdSW+gUX
W.fK,H)LL1:@0-b(MFHgUL&R,?a)Ie\eBY)TMF22CC;TG[=V@])#<-U0;0e-5d>I
@,MM)DBaME._KPfgKbLAb_R4TX.76UQ_ZM:DJ)1;TLEM?0c,15PL&;[TD6-5B#XM
D5,eRQZ.M+4H:1O7?a^5GY<3S7=.\gCO(bPSSCOR1L^I3SF+5UTcA/4fJH0:]C3(
](\7SK6?XZHZLPV?IAUWX5g31Ea3=9+d?1bd_JC^TR8-DL+VH;XM[8U>^A&F;KEa
)(S]Z]CA:0@].?(4c>Rd[:ANR)G9).C[eI,c]_;;YfLH5X9/U5JY5MTGA<3UbfY.
VU]+GD+T?]cJ^0;OSgE)cgZY)-?2&Q+Ze^_4]V)_5[KDOE;a40P67Of?5g+Y_=9L
aJ;Z@;]2][J6B;gc+<8:?G>]_f<VK5Q.M6=T@de)HJ[K;A<AO.0^@W\N^Z);T7Tg
c[BHIFcR1JSaLR7/-#Z]H[0?XQAOIDJ+)46GDNNX86NTZ@(^X@O+LG]+/U>,0Y-+
M]Xf:JE_DUX?=4-bX_O=&58TS<a&c2<PVHXBTcf/=UY4/9+7=3Zd.GgG+ZVHOZ7[
P<8,.^;IP<CW3W^A8TL&<RC9W3[N#80?@?Ha1/V6I7A?Z&L>9JO-2.W^U6NJ6H4>
M.&676^W5;8SSZ8^-c,OZJ50HbSCU8@9[Z_:#XEbE;P6CBdJTc@-;(7M>JRQ.?)O
EfK,:H:\ZO-4Q/__:C+A)b9]0DL01I]_LO]Q,=0[_T?4<;2FG>M[Wb<>9dO()Pe9
[480Z0c4O?0YD8H;:fWO+,c#D@0P?ReP3e.0R]CHS8)>90IOZ@/<caDK?g[Jg<Q/
>SY2LVAT=5\2S/^2-RNH&)K:P,[A74>3ULY2L]]87?=H-]K5eX3Y[Q6UAa_Kb5:M
-:HVVKR1W5:e/U,CO9PgOB:NCc@[OZ3K-^4d)TF@A3cc+eU-?H3J&+L7\;d81)\[
<@f1>HUZ]Z@D1=]9eN\cC-BZR4>4CWUe=;W)J2ZKA/?U]B2\,2#D0Q/4N(\H0D5:
3WEW:c6WGa#^+@4]M90RU1_Lf[&1Ud\XJTRH2OQJ\GU6Q+G\W9_(5g5eXaSYPXbN
,aG)P81;@^Y<+<C):)aN3RI/-\81e?_\T5\6ZWV2K#G/df8dA&^#M2,NC8</.GU3
f+a9/LTFWK8^1E&4=L,5MIQ_M4)c,5#YW/VO@[RTOMD3#UO3__L^0Pf6?)?8YCac
C<VP\8JTc_6.aX0C]:C6;FT75)f&:?XL^bL&N7F3I<P7H+MO4K=1G(YAeR0a9I]]
OEL0Y3C,a&LX<5LD/,>@_2BeN84c=RN.;4a&4S0d@W5549VB:VC#O^=/0W5JNB;+
GGe)dd:WZFOMA3+Y+,4=[a41KVD:KA+Oe_QM7)DP]JW^Cb@9Y\HOTf&[/_dC3@4^
B2^3H^4g,2e1GOG;KES+KIN9@VRWeS\[Q1)IF[cMg6:^3TKMe(<DL0PNdcZ+>OP]
\?[;3.25Uc[J(+ON>9[U3<Pf+U@M.7-KBL--0N8J/+#2=SS9e2TVX/b98/#H6_MH
92>5S5RG-c4D?@K.#C0S=E:Acb0a)F9@06(gJ2Pa<)Ld0VV)4[H]d8Qd=a.:,N_J
P=E_GaV>GYC,R1(;G(#PD]5g>#dR[KfgQ+GJUUf@G/cLb.6)HCT-0)6O0];Y\]c3
GE3;_^,<(-Xg29KaWH.RJ5,2ZI66_ZHKDDP)K/1DgB/C7?R#B[cCEe3]S<C>2&XC
P>]2+b1a]ZMT(H4\5^14LWL#6b=(\Q=^@@7I;@;[1Y.,8:9c2LL?ZSaJ^M^1],KH
GDPZP#[gR^WEg+LMKKO9T_AXfSddA2R;?^GNFP/+3\f/3^ZBeF,eTZ;EX>ZY2+0&
OdQ@DM,6HR7N,#ZQS,>]\\I]Q1\2@b>?R@f2U1eKM@V8U7IUM)8/64f0\@+,O,AY
^OcNPL)Rd3bbfc;g]b5@-CL;;+4?-@DRc<EV<(a6[L1K.]HANCGU-HV88>>HWde,
OdLYZ+3,d(60146d<gOA&_YS,CbQeT1;-d8,#Pd(2S8AQW&dc6Pf5Yb=8N^T3d[b
VXa:XWI1T3ZSZ^+9N_[:S;B1N20BAGKIWCEQW9(&@DJ/6X>_IVU&?WX<1bUT/WS[
QN:HAVVf;e/=X=4dQ:[ggOU2YR-&a_E^=\L_e(E.I;I^<GCJ4;6@M3T+@Af(]G)=
^\[TG6O3G?/:Qb&8J2(+@AUV&M87^G6Ma>;LA&97QH8+=.P>I7^>bKXgb4^I]<A+
R5M4VB/Z7](M&W?VT4T-ce:0(8)D_;,(b+V4CUeTE)HUTTF=?(DO4GeY#Fg/ZX(H
LI;;:G&G2=L/[0484@gM\.EXZ:7E2=4<UCBCg+VeB;02XHRU&L,GCcGEV3KSO>RO
d<^8XB-L5TB-W?E\e7.I7P341MCDQHWNL_(#J0EM[VU4;F6G5QCfYJ5Ub;L,:FZR
I>)0GYg.U633g7@Q\GTAQE;BMF;ENNEPa,1DD/TZ-d.bW?[JK@3]S-2&-BT)d\8+
#VKF#/QU9aX/BRM(.Z-3AW]bKSMP([Jg-,/Dd6KI3dD0QSW;#L469KP<4<0fUcIQ
2D;+,&W6ZL3??F)M/>(;IPe..Y.4M36S5BU/CNW_<&,^I57f?A1H2aEZ-8SQ>,c[
)^HVJZ:-#g#^Uc:fAb\Q^=V,2SE1[QE^HM#EC4XSD2Y<gfYa8:_7&Z[cB1-Gd3@Y
UI51)ZED#C?K<+b3RV,0JD^CTE2I]-?\B&_K1eMVATAD-,FBRUR@DP]UAZU97f7,
QXP_7Ee,[KS->AVU<@(c:<A8^;?Yb=a#PBce?PcX=SCEM5AggECYTO&)4,<@PH<6
&NS)DCPg4Aa/Y6T@Z9Y5K[&]63c(0?.RINIC4TR#_bQb:\&R?agX)gV@]N6^bZJE
X-G8X@N.\:L7>G,KR[=88a_A(d8F4I)>J27-F#b_eEQ^GUfBCgc;QbRXFF93?G^;
N_dU0LW<V,O()EJ0,&DW[DIM6Z]EJL<K9Z],]faH.^Zgd]O6>H7(5ZEa3JCD9f3Z
4VWVQW9AFd;CJC4&NTU4SJLDQYa.R5A&bJJ@R^S.](-?[_#cTb46Q=KQ@D35?-Zb
f6IR0O6?T->?O^;a^ZY4ISAc-GM9H]0&4^./HfXDFNNPD_[,\KNb-NXJDS@\Fad_
TV(J5PJRTX3]A[@R)]gV(CT3E^RK&a):f60B-UeH3/6_BE)b0(L_CbI.KaOAYL7;
?T]6V<S1d#Se\D=c-N/+QPKZb/NegX<a#C;T)@\c[dJ_<C7_5HND]L-\\16V@1(P
BI6/S&O3[H38PQfKa1##O0b.faN21/,gPG_@+&ZRD(<LDIOg9C6S(PZNbDeFHA9-
]DAeCQ?3^fE:V.F+WFaSJ[6IYF]D5U^&FGKf.]6Hd2cQ+g;J+5DTUAXIS=LAbM\V
A-#Me^/9YG9+A4f_9gd)/#:W;8TAKGK2QAV2M)JS5]4M#OC,>TY7>X@R\Y5W-E\Q
:UVE]gUI7##2Bd]b#d1V0dA1V78gS/HI&L1BX?<);&-OZL=K\.I9MZ3b0a:4I3>e
\(\HXLGCTB?.J8Lg2-0^X=HQA50>Qe@e36Od@]F94aCBP9Dg>7LV4(<0c^-ed5^@
1[5We+Ub3R@^V02PM=Y#gbe:d,bD]3;>IAGPDWdT=50PK)3-K4-,g+1P_?OSS2ec
eK[XH9S?_VB.e8+(Q@c.563EUBGO2c8Hb,=ZN651d50XFc)X3(OeER4EL7La9X<C
:e?Wa#55g1Z>:8dcN;ZJe>,b_&GDLa@@07+^db:M^:=P@a#TW7fHTH3RH:ES83CF
eV5J[/>bGR[P=AFfB5<,LQ>1HbX(gZ<TYG:bP&E2AIA</6)fA4c=289<62VWF_6b
?0]d7\D7TS-1].S340C.]TC@]OYN4K1/LV960.LYPTYTCT7?ZT31S2<96g[.7SC]
R3NS6+Gc<)VP:,M(+F;/+&JZF+&8N^=&<_Kd]64\=?H-Ub/0X67@NO2c4a0TO(gC
c3a,gCHYg#(a/2W[_]MB_gAaRN<[J(40?OHE-_I?7\D#J#01T<U:gC/M@2f5d,]5
D7?7SKD.Mg>ec1:0b@Sa9)661E6D[+95?cNKJ]bS=HZ9LPZR^8@P&(2@eY[GCF[V
G1=,LQ-^X?3O]AaY,P,#_CgPUN7P/80D#^H+fSf+U8E8G=&N>5>P]e>?N-(fA_af
-QE3Ea10#CJ7CV[=PXIMDI6OO\7UN5UQ1G,+\JeD]53ee38Y[Xc,:;<-L73+/S/E
3c)8,-5H#Z_]\0a;\M>4D(B/cLCX,1?:GEV1ad8)DF4ZJY8-LN]]X39;;.E\1[_X
#+BfS>;GPgBfZSH[2f,L:R^X-:+:EFU3X<7f86e@M)C189e1dHW+M_bVP22AKOb(
@[ZD;)_gg@4JfYf>QL<</aG0H?1:\=A9gH8UbLO+B\.d4NQ::#K@NC@)2\_5Z9ME
#P28UJY()[J_Z:/.2C(;8KgfIg1/(Oe7_7UGKUcX;^f>N//WZfYE5K.UM2@:LXX2
RW>L^&EWb@;,Q-<A0L;aN_H1(HE3dYW^HS;9Dg,\,03eVX8K0(\HU04)C@gH8UA]
&^a09IX__/V]O34ECY>&X4.E2a7597DE@,fH<,GL[@6SK_^fDO4F--gX,P,KPF8/
>P/+.0dS(UXD=-\&[2^=8U?,5.Z0gW30+<LPOVF\eOW]9(0Z_PO\^Y6NAQV&Gg2V
1Ge<G?-V^9L2O5:T2<#KWS4X_F(JWCc(_HL[;d8;;P3H+<.,2LZ_4.=:&Q?-(:MT
S#KQCfP1P)--LH^2N_E(<W9;+6Ef;a./5b,)1<cQ&?,.XfINRVB-#S4F+BK:Tb70
/SM1=I)?UDe]\F])aX+[T(O06&91AaR[M4/^JO1e-dP^I,B6A4V<4:S9V8YOfRF(
<UNb0L/-NTMF^<^f3)DRSfIBU=@BSX],/RMBf^e(Sd&gZXT?7P@4Q><3&@U7J,:.
9^;OdG?V+b&gEgL;dc-IP6[&T>_N\:B;Ea84)54K7AJ@67::>IIA=8@>C+Cg/,#K
/eIQdE@+JYHf+?8OfZ-UPg2bfKYBEH-AD@f:?+\7H--46^P?;I,\XX;M4/@P,6_f
c?C^IFL:HGSG;B>T0MCBK--GY3Vfe]ZDGY=.XeVG2))/Z9^TdbA,G,#@8a)1/+O>
bBM/S@gKa?^N[WU6gEWHM,U<5EX=M@C0+Q,5fP/JbV<aB.X)-=QB+C8J(#>BRA=-
O5RGG5<aV]DKO(_[6bXa8OSDIX617F_2XeR?eO68bW<FDK\0XTC;>P\QdJCK\R.T
20R=M22aHg?eK9M6d2J<+gD_1L9TL[g6F8gA)+C>6D)dDXbYBdRWcY_eH49?PG97
=;^K200CM#Fb8G\?]KH4<FV>KH/D-1#M=]Y:[],>)>-L=4Wd/c7PbQ+B)IPA?0b;
E&N(IBcC\I#;3=44OEH]V<cFe54DR#^gcaa3BW)g2]@K#+;;EZ7=478?D1LUL@;Q
>d&b?+I+QS+V=)1bNB=M?IN[7G./(#8T2R-AcE0\\TUZU7Z0(8Bg6BMOZb)PB,6#
))+YPP[SI5QdVDC3)b4ZBY2-VVV?.b#]L^@f9TaXFYca>&^./GD>9Ac)QMPecf^S
,/U(\D(92-g4=@SW<H(g:DV.VE?U3[[d_3^))RO+HYA<9fc^9OURLe+P?^aCP\\b
(OM-cYD\@a6^DE09cRHV.2N=L]ZY0-d^X85/&/0368UgAYeM8B?>R&IDKES:\TfS
U53DXede)LRW2O^CM1LWI3I_8FdHU6B(eI51^#<dDVIS]>\cC]7ENA(L^YC9XLR[
3,XSLG/YNOf@F#>[gTeL/O.g42Ea]H/\O,1&44E4Z>VS4Y:A70O)U5<YKUfC?3@O
Q1DX0I-NTS6L<UO-<^XTD)Y]cMA/)d(68Rd6@F>3\)PD4U,2?]CZfGSR]B=:eIB.
,.A/^Y3V83>J.^I5Xe\7EJFZK:@]-];Td&,A/.>:bHe7.7aPMCBaY^EDdI9AW5ca
1IWDQ7U<2<B9XDJV1D0D>U55V:VM@\WU6Tg_C>]EQaJg>TY9R;&CZdKZG.Gde/Ag
]<6_b\W^G&.[5Y)ZAcH@Q@+@b&KKSBIMG5IPbZYOfKH^6MVQ]/O?V)I)-9gN8OXE
f3N>#7]3O#O6HAcZ0eWS@T:&6McJRH#Y-;G]9)KS:P0>36YCC[T<I[EW>T3JWM:<
WfF+/<L0;K(VW9HJV<a3S:B;?9)fF;A23dK1]<F0KdUM@4Z65Pb[[>W[]eX)?)dX
VNCK(.6U2/I6eX9aecf08//RF0f+<CJ:dN5/R;e#5KV>0P?3YCC:DM]/P4SZD/&\
Q<bOU)YRFN=J>b_&SMQN(I/BYJ@;Z[=cc>[N:fS=J78X)RZ,65QgC-;f+EKb+[WX
CN)XAM7\Yg[T;ZYHVOVYg7-U0BZQ))2bP-KQS#;e,>@X#9R;]Z+HP.E3)T:W9=D/
\_XKQ;NM4Q]/_LP=eAR@3Pf(8IB:QdK4_Y/AKGM8S-X@a98[Z@RS1B321\g@KeTd
gaRgB-DZ\9W]<,Va.]AA<a@P;3X-FS&dUMBH4(WGc[)=dS)X10I,.gRQF2CgLW>R
94<2E&NE,e2f1>Fe[01g&<Y?:e]YYT=fEUI&A\&.M[Z6FR0]4dC0CPFa:9U4#J/;
DH&>gN8HEU0@YLKQNY&\Q?H3cTY[Xd)[TLISHB.6XC)2>:=(;W[([6Y>5^7#f9/>
G7b4UKR^C(@/>A-g(/^7_cg8?e9gKd-5cc18/=VK>.02>f)=N]E1,cMbGeX?VDe+
>b_K>8&69V4If_E66^6VN81S/c#Y4A<>8WgA-+dIO42gBM(DWK7aSS:)aQ4,+<FO
QNc:2eUGLF_ZV^@X)=L9QF@2;HIF;+L-[AgQb]8>RFQ9=@Ma@9)=7Q7.ZXEIPAb4
@;cJA0fM<][b/E8Gd^I=6)f#H^-8>84]aaR?R;RE0BKAbIUT@2aac>(=I/OR&NEU
9#&d>X[P.FQd6CJaUQb6c^LB^9CKJ&WRYDFcH&V.DVG^OW?0VAPGLBK(Z[IFC;UZ
>0T]9.K-NfFRa;C1)J=+RK>,g<M)P3C;?8[AQM,bE6CGK<)aKN9)dMHZ5?)dHWFN
=I7?7\R6>X=cDJ2SC2/_R,0#;[1^9g].c;I\OaSY0cW8Pd60ET+?=f+ZERTVZUPf
Z.]Y=EPSOBMBV?U(a6Ze\W.QRRHKKeE<Q3b>L/6[aSSU]N7DZ;4;SI)U5X2F,3JJ
BEgPT?&Wa9Pe&P\/C<CWcALJ+g\HZ0)2R.XF.-]ae?3#>0D0PQUPM\E<1NAW7JHG
e&H3[4<aV;=U62ed80EQ5].dX@IY]BAL_NW,S_HJ[/23=WAdT-:A^GfPa.=Pfa73
W<[d73ZBAD3ZVP,/YTe9?WP5P@4/(O[?E&AYQg[E\)OCF/U_5-]8[XT7VIK)Fb\]
1(J=6&=S7dHGf(K\+=YbVTCQ:DMM0WZMC0IU+TFEIG,<S_+&dOSGMY6\QKFDJ]_X
6<H;KH0M78/3FE@b.d+I5<?J=eT+EAcCIdQCH(@[WF-5]3K(\bV12b]1J7C+3-fE
:\=Y0#^:]?=eY3CKB7;D/A1(E\(bG)U0V_H4HaX67d\@C6(&2Ff9>:gfWg_b@@M(
X2)@7)98+^>0]V3F,a#6TeN.Bf5R_[.6a9&UVZ&6P.6bMGgC<@0Cg/OP+PY\#g2;
\P9/K\D0^=S\b8_[Bc/ea\4;O1GfY.dWMf_?#:cJW\SB#=\SAM5G8a(W&g::N2ZA
3LV>G^05\5aZ0Kf3GW[;CeaG@\SXCOS1><&VVc(5MJBUa)3Jc5I=XU0S.I71GF8V
3\.XGZWQP7K)EFfAVdB8UV.;SY]9/=#+WJQ-/G3(1?/)QW;<V?D_g?Bf(gEJ<,R?
B[US1_K^&3/9^T,92MggXCGTJVeLQ+HIHCSN2=T;-bfF2:@I=F,T_CX^NXF;MQN]
XJM+R7OC(<SeQ4.^bGA)M973MP2AV5&:>:8)RbdS]E8QS6gL+QCcfN2F^S2:#&C#
\)N(+@=YX6EF:B@/=QJ/N0a4HC/;RNLV7/A35-,cVTT==Wcd<[^YNQ2W.SCQ5)+^
4FgJ\R-X0IFgQ31ZO6WWM^[&:H13UJ#T^UDN]9=c2(:WOG7fUG[D1MW^[18HAAY?
?2IMT0LT)2<2a&4B.B,SUU7e;.3+-aK&:,gbXcB&46U7Sd<F:2DALff=a^-Z?_?D
HA8I@H>N=Z.V[N?W#3cBbN#GEDS>M]8Be)#Ya+:XD8K(,YA)XF/N;_>0_]9F;5UB
RCA6eE>I.L9(V-T2Y]-,b[_J(TT#VD=/c(ENV1,)dF92C3)+O)Kg(;)?_EAG3=IO
B6GQPHS0\[OJ8A5P1J?784H9H79LYG,MJ3FH61(C&V&6W^\\7@-b.d,D)[I3JDQa
+G&OX9X:I,.8<:25[L_XKZ<PY=?^/ddF(K3,X4Hd.K4f=H]7e&4Y(d6.JTL<,)@Q
(A(&YdTG94E4aK@5gT&;Y@aP0Z_G.?Pa;ZM4W-UG=7F0J\QXU=YJMdNV)1,Z=6aT
[/PQG6C&ZGC#3@EfdMecNJ#2Y2&g:&>-DH-?JY;CI;<2Q?-J.bYC]A20(Na_Z>Pd
;cMOY>IVK(#)67T/EB^M/-Z@N51>I^cDSBRc]]BcPC0P&;LW\)1gINB+OZCM28c;
d=LBfc#_:R/>\(T+(8\aQKKYSM7NNA73^e.<NeSVW<eT..+_1.T(IaT1GgP(+CB&
T-L<Ca6WGG?35cNbY9W24Zf57gUFB[+D(Wc0^;]//gIff^<_2SC<T=2BaYI6<#TI
:X6>^QIKSN7gdC3)f[AECVVO6R?ZJ04I1MZ6aLQVVV6J>6fD+7X8R&X[ff<20G].
>TV+B3PW:>^BS1@S7LHK1d6.9=[88[.89HT\L1Y?Wc)Gce:fB?Z2DD[N,dBeL_T\
-ODf-GAG:@AJ]Y]J840]3:,5M;40gfNO.4Y\2IMR].2[5.^5gY,^L\-BeAbX=)UN
_4L&U?(-MYS^a3deL).d.OZ()]:-bJ[=3cG5)FG@Pf.aIgA&M>0Fad6:/;:.4?TN
1^L_HfVNOZ@U9:2Q5K9+TYeb.0XMYG-\0c5Q98F:8782P,_9VgV\S-L3-,6L>-:K
>WTR.IEXR]5@S\3KbY5LLd@\UQe^D..LMST]7IU&8SI(4Sd95SF,H3D2#5]Ra-P)
;[>cBH-:^6.?NBP9+g-1G?Gg^K@98gG9/7,=..2_:aBZ/Lb:YTHfY5J?(J[.OK[c
TSbCgF;(H1ITARDDWgRW6+(X8#+0V(@d:ZAVX_@W<E9[8;3F2E:4fb7R)2Xd(N/_
QXaRg_Z,55PR8>Jdc<U]LAIM96^#.\#-NNC@S5;,#<I>cU5U]2THcfdM@6WEBXP]
@/5d?<774)a79DPUe6,^W\0K_bDL)\DBf[9O,TR[aPVP@EO=UU7/_K3J5=(C^^6<
5>KFYLdF8Cc^gG6FY#UeKC5+Me4W;=&9,T.AAL)#IWD^LEY_T#&T?R\D^#PbFMGN
QY_=LZ;1;Y:#4?V&?dMH<=EbJCDfb,NB3T2^>ZC2Nf9#]VTWgP^b[@K2F=eR\N78
[><I9gGG1aOP,BLcSZV-3eC2D90SB#P27&><.eZ/B:5TC(Agc]SFY\G8;Wc^&b6\
Pe6&ANZY?[7bG;TcRS[I5KBcP?N):\B=P9>&VT:_^<-FL1D5WE/>b9O;JaALB:14
/\=>bb=TEP,[=HA7QY4UVHYQ@^@[,H\Yf<PFJAcJ(/bFdQS;dSg/XQd91ZTG^NE1
BCGF,W=3-44)g+<&X]/SJ]K7Mf0(gHMC/1\/#:.TS0,)cDR&@BNg1,Y-A-SA0F^g
d9+ceDGL5A9>Dc0X+;:4/-@Q#WKGJQTFQUNIQ.8;NFG/N8?+c?:AZ(-VGN0LcaQX
Ag/5DXKGZ5ca=6M9S3Q;,?b+ZRVQPQ#<GM=.e.18-@D(S?LF7QK:;/IGYOC.:OKX
CY9;3b2-/WLQ;9gMJA/9O?+5J^7.ENa/R_c=JWC>bC\;RDFZZRJd.N[51J@fY[AC
=Oa\-<9Q?1A\L=\&R(;S+6D,/EAB<6f.F)TQ)4)I,)8)8CA&.;Y5>F\5SNFHYPTA
1(0-cWG0O+:NSTE@2:#>]KXW@WP&:/P8_IXV\&Ua]HMaWFdegYS50L-,-2QHIc\Y
WFP_b.]G#IH>R/He9&cE#MMeV-Z^GJLB]^UT:?e,/ZG=J[aPMSC6XK;1UMfGVN<7
8TeX/1F+Z<M/]RVR:C,UQ2QLYK7dBYaff_(#(1A+P&#8SHdOGY).7?K\O2Vc3W-_
W2HZU1\NY)+;Y8FSP3&._f=IdfRc/3GFf5g;W\HN[[7J#f[5I)G2aRB3;&,LJ-)D
:1F6K-E@]1)\?^QS4:F-25;RL:WF(QReL^e7IX/eS,?V&dCP2-O^D/-dMGN#]V#9
1K7BH2I>+gN0;aTVC3g@=GJ5ODGPQ.:X4.&Xb:J9E4XY4^ZW(?^_@N()+/eX;W>#
f](->N&0Q9],55M#(&c_35]?SMUf:S(fXf]IDAgJ=<=2[=RSU:/<I>cX?6TJ;9aS
4e5\?f_98W;71gV\S>_HWgATPLfIWGbeXM=O5_4U88HFQO-2bc+;d2P\R)?a6O,Z
_4?bTKd(RJ/2I>,RfHCM(e/?NS9HJRISJ&#/(MXHaWKDYP\N1QdF&EVd\WNG&G\L
bWV_GMXZEP&9;a@:X,@K80/G&eDSZ8R;U.DgL#4TSEEL8W3N\)ga:-8[f:9YE).<
a7.>XR8;bP>.;@,+GJ9UC[Sg2E<^[c./+g>-Y9FPa(]S20;MT^(XEU,1<7S=M9CO
)F?1YF=55/1_\2eJKBe^YeX-f(dVP+W5T)(@E=;</cX.LJB8631Z[QMV6_c)#4d#
D3_b_OL(-0)WP(ANCW<d,))].[M0SO1^BHEN\d>fFI)Z:ZF/4bgg&=OTKKYbe1ZF
aL)BFd>J[)d-Y[E-CBQdPBQ2JROJ#C8))IKe?I4dScCR,C,=(I_f3I9@#2;d?d6>
IQ\WSM^E):eI)N&AY>?I9R3ZW:4,3(6F:bcd#MJII3daK[K)5SR4g(3E]c;+6<Dg
N6d;:/8[O1CCU6;M[MAG0=\Nca^Pf7;YW<cGa&-.a]c:3NM7?4=\:U=DMY:X8J1C
CY2XEMbe(MdUO_=ZPTJ,W:#=P[(bRg2LDIMX897>&O:ZY2J_6\a0.#INTMUG2YFH
I#7=#JL+^SD-ZV;[EY1E,V]D8XQ8B06&(C?I3N&/(Y/V]\B9&0XbZ:,(@\L]FG31
E##Hb=bCb/Q>.9IM1@C34]>WM+)G-C_ZJ#gD)d+PA^JMVT6?c3XUCQdZC/4IC265
ff@e9)gf1^,3a8NB=NAOdYTHMH-#cD(5?2bEaf/36[;;07#0K)>DgX3#F>@XT_aH
__=JLY26U@bP?9?MDG=#)DM]^FC1T,e^6#C)0O=[e)bT=&=Y>3CC3Y+@6[LUMA8L
bP\ZCHU>[=F/(eSN>NC(:FO:9eSPcSC)ZDAeT/V[?//PRK1QCSSbAEZHB-b#;#b@
?-FUSC+2_LMV1.EcBQET:@=aPf3VW3Q#_1LVOQW7e,=UR)?[@I<0?Y9&45/H=\9T
0KLd+\DARI(eP7W[,[5ddTJM]HL72FP:76D_1W,:.gOb/&+[]GM;R4C+<M>_/WW6
c&cVIR/d94RLM,JXT+LM>5_/[G_[?^J;Ic[4,7]^HF5dI?,7O;_0G;/XU6)ZT/12
72[aW>KJYe>_@PCLU[e/7A:W8VM\9C+JO;0&K0B3FLN3aZEK+8=2R<[MMcf-:,[U
Y/?J,U_=\ZI@V4e27=U8+^J2:876WPA;H^=:T<a1W=Z3-7&J]WB>12AOAMK0<d\Z
QWd3NUeEO?+JW<.\\N?FTB/B52Q4KEgBHG@9D@.L-Y9:F;:/L9TWKC_(_>EC3gC[
.4Pe.O@J-WKXA(E+BA;1b4J3F+1:)&9?]8@?Y?-Q#:XS]HHgbKL&\?QE<)2=[\(7
=5KE,WM#I7;3+-AI38PJ3&KY1RgW0JWb,dJIYAWdd8)89[W=5VX<BFLObaJ>c5a7
FA6dYAJP[/MMS)L_J?(K?fge36JcD-,fXbD104H]d0df8155>\.&D^M+R:PB1A,,
8)+6[e_I6Y7][&23VEH9@GD,(N5/3F-)&=aW2YQB,^A.-,?9,IP+[;A4/\4J^A,N
Y-@_Fd33.J)c.BA-&2A<+;c&&\#e_H6A@&82RScDYQE<b&/bc4a@NX09CbEf\dLJ
bU:MgM;]W3e2/&^F2EfNHSYJ7?d^:4Q@/<K@;B?L1YBEI78U/J+6R#fW908)_g=+
CTG7eXP-AgGB@I^5+MPbA1R:17:9W>-F]@7:LAeg[K23;Q)T^A>[#.9V5E/_KcX\
TNZ/Z,&TegF8fI<G\++LMKCWBEYH9.P>We[-?EfFd/Sd\FV2^4/&(-XC9[G<cWg&
dPBUUC+cIbcgA50VeJHgbOXYMBXg0:aB8WQ6C]9F>fS_\ebD6:+0EQb_DF/J>c6W
&SeSd\baWU34:\:eE7bcbN-24@=R5:[]31aU(b5-R[ZL?4aeb[?TF0AF_c:^6-d7
d:)f&cK6&LF07G<DeR6aX:</[fH2_,K1MR5B&UJ-B;G3BCJEMWdAJ8bQPeH0L@E=
6S(0AFVJb8W<WP.:8_3=K/M<Ag(S&<H,&K>Q7DA-6X;&/?<FZ6Ed:TI[2QLb/1T8
=&ME^SXeVY8GGR(KQ7M7b4E#?5T@F3EY0-daCfN3<_KJM8-C]4-,T[C;:\H,Z(+_
BW\2,VP:V+2gRV8(f]0,F>]&@M;U;]208W<g:O:bPYdVbV\5Y1=[-KH(I[124-O(
3^fBDg\B)TR;4\4BAIYb=XPB\LEPNaYSO/4e1Q1.+07683@V6=JT,+ZP7UE?RMdB
cdgW#8LQ/^AC8;.d@^B+()T@^/SLCYB/TdU:SAYP]V@LIN/PN@H9Oe6CQOQ(0cWc
O0<VICV1FZ[#Z/gI]9/C9VL\Ye=dbIRA)Q+?0R#ZZQZ[H+R+d7QB,7R^:<EVdN=a
H,0;BIc2e4D_@.MfHJD35OG;EBSd7W4McAQZT#QJ>^\=dM;M-b>LHUG0gU:\589Z
)2#@7TANKFG8B4=&R<7R=e@M30AC&\HKG\@U8b:\Vg@9DZd9I8[PK[^&#OY[[HKf
1f7&/[HX+&5<[6.XB2.Zfca0[&e8SC3-eTJ)V(SU_8M6PQa,62A1#bU^8NbN:fG4
T5=4@A-IQCb_,/9P>UgEe/K:8O3X#1+d]LV5MIXC),M@[^aG[KMRb@b[ccRggEA,
^g[M])D(VcK#P4:b(P>_/<[W9:bBH9NS_3+b;//;gfcO6VOL&BT_7aH9D>N/Ge@;
G+VFMRSURR2ac.Ld\U7/KTcOY/Y2^SdPBE6/7.6FFFX^E>\<0KMS+FEC0D4gW9A=
5JMWcbe4e4V+]>fJ/EN#14Y?=Y0_PO/<+aKeEeM-L)6XV^FUHW6;Y:eP^BTCZ,]+
XRH@X.3-L4Rba^>.YR1Y\;;51dCe(gFY=3]LIc+T5RH5,d@\g_UY7dMY@FWC&b5?
HW+2-IUX6A<8bY90NEWb5W,>E.@+V(Z<.0c?ee5LeQ0-:EWLL^IPTBQ=+)OO7-\5
L@6)R0TX27PN#_a--9Y\g1>ZAYW#<:CZg+(\2&H8Qg:51VHCM8^(ZgJeNF@8O=1T
Ea^&.D>.@)a9L\OKUafT4(cR4HVfR2(L1dN0B=)9EY#:IRcFbQ^;IFI/@b)d5fP,
;FE^_=U>-\bK7Z1e#YTQc<2-J(H&W8:?T&67>V477=>6[4_/QA\^2+VP\78g5GZU
FT)@T7P[4X2OgPMC3UU?E4L[A_MUR@;DNWDT/7>5[e5fJO-XFRW04ROcLVNBHII0
/-K#d2E5/Yd.7RX>GZ_Q)JDCG66<_L7ATUTeT#>X_3HMB,Kb(U0H5LKU0CW-c0C5
M?,E5.F;V3&c5U/_<feM5.57d&AM:0RT-\G3,SO\G;]V-\X,[A?fa=K&/:.#JAHZ
BTA7bg-B>J5H@.g)HKN&fH>Vg4QA@7R&YH0ESC^THMRQ@b0Sg7#C0;QWWdFDCKCO
Y]^f0S.0E\(4e]3&EV0BBN<0[e;(CX;DHY&_C^#bG-I.4dTF9N3W)XIR2+[),63C
RB;&-OUP2dZ\bK0\3+6E6UCLN]]VCUd)V4<Y[<c]6\3>UZB#/K9[1T(_+b;Z8B^6
U;BV4:&M4c:(,gTGc_73I2FYO)g6XfOYURY?X]aFZVTc8#S;4\_-&#A9=2b]bS:K
W&,d(XGcCdf0)S_2V631d-Rb4KOVb][69\4BKO92X:+[G<83(_GaE3AN?Gb;WYf9
C7#W17-U6>;UMf8Z>0QaQS=&fHWBe_VD2ge<KQM@f:FW^O/M<-aNd5UgB)Z<N>Oc
5Y?/db5>KFX=9;=JQ/9C&#7@Q2C3W)R9.1(_/N.UR=d4S6J0MZ8L[\cC^]+g>XRK
=B)N35K?FDa]?Ia7\ISc)&&Q9g-IGU&UVH69e6PSEXgSQa@\P+NW\Q>+__:[_Pd_
bQ2bN#5RMEMS<Y].N4NOYc;7deC.TaJMDT+)O+.KD6Sf:)\=]HTN/Z@W>66g3MRL
]-#T_2Sg?XOcdL5Z4_e6DM4&P-?8I0OZ.#8cV>E\_UF&6+P:Q-O;0g6,3e;eP.<N
1R\>VR37B><AQe\+SeN([9XM6?EXaD:XAIF_@_K+IFZD7^6S#Q(He0E@/SQ/S(0I
FSJIA9>Z9#&ILLfJG>A:K/a^^Pe/.\RAfB?HI=+G9/EDbbT]0SRZf(>#AdXOcb_,
.L0g+NA/[Vb/.dHPPPL:g\Yc/JP?0LY6,20Kf3M:ZKU_.W4e,Oe#OAPV.H>8NWZH
I#96JPJVg=,GE,KWTC8+8BWWY3WYZ@3F_dWY1:PLAW;:M<76V>)?H@&QT&);O#b3
PPf@,#c\:?9g>cNAeZ>T4DaD]>\+>WI1?aB7__?F-(EF4R)IR7eRfcO9B3KEZ\H/
X[Va;N-0>5RN5Y4DY;H?;NCfgQ=P\=?P=5SW[C1^[@@eb>@>5__X-d:aRT/(cKC,
[+\_+&K@]..[8AD26[2VGVVJ?9d0CBe5+17_<&1C9P1Q(KY)gB7M.DXc#8Q=H3:/
E=YLPQC[=<K>)L4-,J3@,S(BF?S2_C-7OK5]SULQbOX-JZAdF=]F?/?DW;UKB&JS
W92NdUb]^>;5-_Fa55cLMe:M8=dJL\(+PR6?JP4gHTa\+ZM]H1WgH>K=Db@#?_3:
[0I>QAADT:0KFCN4X3.;]<MNOR]9>_6IDMB?HMEXUBIB=[\V1B>b#]0_U;CQ8-3_
4)\2S6&+B>G(T<Y)?]4Qg9AV]Ae0D(?AS,Ke?\gN\O:WN^)H)&N\MDDK^E;cGFJ6
:L(U1,GMD53>)F;f[ZHTa.C^gC>XM=ee\/,NbU>C_fg4YaT<7<g_gS]d^<>L1,O@
aCBg[GPGNaIA-;dcU[+;f6.<fR(/GbIL2aAE@f8IF>D1,RH6;CL.7V6UY@1(RG)Z
HN[F\AEF7W,<YD)b>)fZ;/d=?PB=1C,>/3[3bOC8:K9K9=G@7<AUa?Bd8\-6BI++
fYXQ53#(<K&F5R_dG/^N>(IC]UF6B5U/cd2-(@14\.E6dS+KM]2>HT0^X&@7G9<V
?WQ&:aXMg?UPWdX/I#JB>WRHc@X=ZQ(1N8J>/cC4]Z4Og0@_8Vg9DLHV12IN?#\_
Ze<;A1NF,N\ae9HJX1<>3L.>4,Yc_Z\B<.@7]d_POH>WT5P-R@,L&fYIbCAgEK&9
A\Nc9O(;1+]7;f,+.8gE814FUeIB27ZgML/G(.-M=SJ([&KK#&Y95?VA<R=GJ@cC
NFJA#I/]/]f-6NF.WC\=+2W+?d;8,;UUO#2K/TQ0<DT9IC&X)W8>.IJB<c-&TE/#
g,GI3ZHNLb9\TX3=;JC-W&U;Y)e:e<KYQ:WD#EUdW+-&L+9@IUedYf@4C5]E:d0D
=+2X4f@S@c7-MQc^&cGU>fP?=9,5dLXEC+eN#7O9P_gaL)UfLSOE18KAXUbFeb[)
M,^77J_^]\?da#DW?B_#K8F91gVXc1I1/P5-.LEa2OJ,aN>P_SO#F7eA8Adb6AHW
,H#B-:bEG<36+K;aV5T9cUD45CCVJ)bRdN-f@c6@.0]?5V3//<M2PN?-_MKC?0ff
:1)5=GeG[I#O<:gXU0\1AC9PCddJCP1-UQ7WgBLY3G&\ZB7e7T9(ZH.XY2P^J@7F
1&gGAZ4EaK&XLeF]K#2GL8@<gc\_(>^,RgcW#^D7B3^K)aeUTR>@@6KXdQfcW[XD
Z7HNYWf&[<S;d)[Vb3A,-\^LC>YT]ObI[Mg6a,=^W5SeDID[_-,&A^9U-(\,8f?M
-W63b(;,E#5D\&/VX<5RH)IRcDeBWKC)NR8ec5;DZWNQ]=N8EY@JJS#V6a5Ub]OH
=SB\(/Gf(=+EGAZ;@QHI)eWSZ3c4aO]:dfF)9;4G0a4K_IV#7cUI4E;V@gNK\X3-
aH\A,#d8LL>NB:L#a^.fH=JbAJ^1>GfW66]TTf)L8Ya-aTV7PbPI_YOXV/:fGWN]
=Y&WK.XJH#75g#GS:__79.7WF9<ARe8e9d@cE2PJNW-S5SROB0cO6YHR_gLgTF1X
&:4LX;,-@>-ZVU[42c3_.8G2>\[T^NJ4[[I91J[339G(;[B7L4+O2f=.BTB8#?N3
dUfFA(RH#4MPb0]c7>U2Z1Y/BHZ&ZVb30CN5>7XDKKK&A><,d<eHg);WUF2H.@Y?
\8:b<Y()Tc+)C2D-KY6Qb@[GA-?beN33KI-LSF(XVJ2[?X)[GKF0(AI)=W]5fH-d
C&H1Y[1V8dUZ,b-PL\6b00QeKD@4:P+]XJY8HJ0-I)<#H-SLDJda9\30FP6a_FCJ
g?HDFAVeFBb.SR1aZ02IOOd=EOP-K+Y(U#22R3LN<U<=+DbJ@;b5d2B4LgYETf/O
]E4H(\MYN,WM(9eH;M-.a9c-^f=:]Ta3BOT[)VMRQX.GKB86Y(Oe=8N/DGQYD;.;
+9O_\47](M^4g=CR5b8IeP0YD#/3@ZbY_(>RW-d#I_FQDd#4AW[VT.J2JWW50A^S
?IX+[Q/e0C@DX?#1T_.b?V9A8f,+ED]M?._2D=E+3>3;^XNF9ZSbLOY6Q^^,da&T
SW]P\D+@e/ZMS^/H&eCdUU3JFbI+ZOMGW8<b))V1NLR1N&-3CPKO5I2c9KY(UcU^
HC[H@[V//V_AE(2(C8N4?HXfZLI7.JX5B8M=E.^([/0:8SE=?18@QR_C]S7,,EV,
Q:1F@H:/AO5Q..,)98fJUH(Vg.,XGDX4aU?C\e;@EVPdV:S?31PZ4VW+7>/Z#7Eg
dZ22IB+-8M#IUQR4dBgHFf,@_VVVabbK^02T4(T6;c]Na[L8#QF&5:OYKFG91^WC
QODOa@^][6-T.8\P8.W+K5gV+D8AU6aMUDSVJX8L1aGV?/4(2EVa^gdK_.+SCH?W
Pf:8:,2K9P,S18#1QaKH?\gLgHBdK0:3;C:<?W7=I6/0_>#[2)R&-J(Kb4&T&,g8
7+TcM/S]4+/GT+bQ5\.^)?W7f.UC.;QOe?M/gFBV\]SI._5]IE+)a+ZcT=&05cf[
M&MDOe#N2GP=?XM??d^]DG#K?&7,L4d]X1dNT@[W5\&R/[.Y7ce-85RaBBK5(,3J
FAX#U&:LOVf>,JNHK4WC=PM&-4-fQC<\\.S:f79^N.;[SfQT.K>B8(X])eDZL>e[
,)KAJ^0d8G([=5SRLW^9ZJ,C<g@(HH:MYL\O(3[B--8\,a&V1^S[\5K&aQ?(ZVH7
5T=J)He3SdKS7)@-8&H&cT[,_S_X+,\_a18)gJC.[3?YNcZ?4<L8HHTVDeg?gG.Y
U:99?N2\+0@?]-1UM^UGNKD#^&>+RTC<_UC&b12O)dH0USQ6H+N([YMb]?E1D8V7
9X<fee9HGR4=OE8#aX^DK_ec#fbE;6fNAE.WZJ[@-\PD//LWCa(GE1J>=D[/2_J>
@-](PZNaT-I^YF>1N]eY2bB7W74\^+U[)-^0R_]D\XHCG6R+\_-T0T2T&<Y:],>F
OaCY#LMA108TbV,@/3K[a^BFOc^5B/UdIZ9)K]EYAK@8&[^)=X-VC9JeF<QI\40P
HLN-=A4X88>AMGCB1)7<eQPAa9Sd^C9gE0Y?&c9_7(A;?YDUA_5WMI9;IJ@/F<[;
A=I]66;CYeU#B3UIQ_<dYLV&dW.#F]4?+I(,I4Lb+8eV;aE2C/Cf/cJ:&OER2&J1
PH?fG,2>U_#W,F-+Zd2dYVVDb-5dCWN.1DeR&fR8:b5T5?]^,?VXG-B1)1K:G#7F
GX,PTI)?F([P-8beCX].Bb@aK5Y7fQPNV5ENKeL3HdU#Cf^;S+cdgWZ4dG4e<3Mf
SALX@Q4+gafV/_+MHKA<IC^d7<+M0CEKO.9VDE2?B^(H>2Y8]QGFN2LM,)8TRC;b
U,/OVJZ@6;dA#g2IA78FM(c_a[+]A79=(G5_56B<Y_]_aG9^,CPUS8V;c[R?&bQ]
?.g)46>X+I]QL4X1fOSdT6P;D?](e;V_f?OVWL[Z4bLR0BU=D;0M.,M+=[B,.6b@
_Z.N&LV7PYL,PPFVcIZTU;_Q/J\@24K:7-ZZM,#<RG^(d4N872,DOLQ?2U?D([@e
\4<M6&;\W6;S;G)aF1A86T9G^78J=7W)4TQ4ff:0^OL/8/CCNW80a/4/->9ad@8?
OfONLB(<2N==(K.0@/J=?9JTU&e4=,R?Y)0=2HgE(^1F24:]U52AGN;&^JN1[DU#
Z_/NWcb9,eNA-f#CA=D](-UJ-+I.ZH73OI(+0(J::bL]S3E9MU+9WWR1]f]K6G3+
Vcdc6TLLM8]O\</^-/=S#KD0O:_4G;7:](:SVa#)QE2C5eIBc-_-P]-T;#caXgFc
EH,1F@SX@gHIc/f/II2ae3J(US)O#ZKg&^OF_H^Z@[70?F=H_S0Q2A&.,VK/_HB#
_S;.d21=1=BaT+@HQ:Q,,8FL_0;TdB6J3Y=7WFY<dQ]2JW#I\;bN]2+gUg[?)+;:
0MDXRWQ4a]e)>\6U:2AP@;gd/N8HFGC5g[=)Q6.G.-+eND0::YW#QYWG?EFN@Y.e
gZB?+W]a9L_Mg?A5gS59e\]HFUQY8K,;O^]<DD-=HF@EI1(JM+/8R-SL+=^>_&V5
G9X2GFA:DM\4032)X<[+,L_0?/VN6:acOJ&>a()_SDU.#P;C+RS5a,;9SM8(31c0
fdfUV:(P11[BR3:<MMe._d_HQ08WP8[G)^f#SG8171116(LFegeW^fA1)(X)60;I
Y0YK:]OL5RA9K[=a^<:5B1\\(4VO^<-5=K^;>7Z@Z:N_fCUCf&eY\g<e:5aTc1dD
B^aCCe)?R6\.TL>d1/b^C985-DZS8@(WV?0>d4cgDL6S3.-,]?O-3(b?5bWGcgK]
8D:QagR912d-JG8-V?[@#J\+Je?:/ZcZT8@?gecc\?1VKVMY3e+8U=eTg]TE:XTJ
A9.FI](+7R.]9Z7^7U0Y2f[XKf([REJ-1S+GUYLK8X:<#T)c.24(P[+C-Q)74@]F
d#[S+#JXG,1TE(44cP)YCU-V<FPRA.M5>S&Oe^E:SXED1.V+M#)4c@Le>EXN^[_[
3RI[0L)&0Z]6U6(#g0&CBK9S+CMKSfOQeU=Qd3VT>8dJD8]+XUC(:;GNLd:,d,FX
8F7E<[HVBA)c]V,fMeGQfL&RgYV-B,fJFU+EZZ0&Sgd,:N9A3>bV?REV[0Vg=<S@
a]=RR,gJD7X]KD/a_)YQ#920N/\/12MB2ZZE0aIU:HW)]6\XaW6(B)F24X8G[7<9
c^B21(FcEW:g6IKMJcET.GHb&^#\#adONLSMLX](eW[d>XOW#&I\MM#G66U>GZ]R
:L?QdI^aS:c24@54+E=\P(g3C?0e-KS__]2(SP9<[96F46@K[18F(O@-;(ADf2J/
ZCL<[_Wf,AR)Bed?QC=C)2&W+6T&^58C1+a;(&bN/(V7Z\^]H<]_B[Z(D:KS#<&_
4:T+0+YX7c.L6YXVb,G.2<3?IJ24<XFHTJf5<E4;TL/B1XDbf+HJK&2]G=Z3PG3C
)ES0e-D_;QZIL:P=TEEU^?&Z?2X)EPScUI8Q)0XZG#Q\JI7gH/7FS-EAQ&)bVId(
Q\<<@Z+LNa&/aXUGKd?VV+b>GOI0;5T/gPKc73N8g&]VF+4F3OdXVG9H83#WegDO
15^UAb@R]0>MNca(41/,NE0<:&T_G)BT.UP0H;b:[Z[S,X6M<e)fV9b\HbT[bVFU
,KJ4X:ffJ)&A/ceAWWgOECR6G/;\IEaWFQ7/)[ECAY:eP.ab>[(_&D7J88F0MB0_
X+MTM7>F;bN,bL?@+_WPYA#Y\]c9O#DY4gT[DG@2D-\ZHgUDS6:=P5-=XdDY1]WD
[M438(<>G?/gKPdP:,3#bHfKEX1J=7FEEXBH\e3L:]BL,ADU:6dA-b,]ECNGHM.,
<X7/DBJbS/?3Ffe59E_X9a#2665f(EU[85fQ98;/7PMTEH/VgUb+.@]WO8T-F(:Q
V>A50+53B(ZN+[>;HfETW;XUR_.A9f@LCG[0IRgZF[D/F=fTD@^::RAK<ZbA(QL<
,FN0b1L3AV>LP/g1QK0)Z<.6]:M_9EO:M5;bA;@MDJ<I5>>Z4/b=O++Vf&;aOXO2
15Hb<DM:>RZc(T4[Rc^<a6f6;<&DacC7&SQ]^AV5-,FIVaZMSdEN1gTPeB>6+)Z)
9>(BL#X08[_R0=[SP5G^d..HB1W,A)U\AXJ.<d,7)0W_=/&L7I+7JHZZ8_[O=<O0
HJb?/S,3&P405.Kd&,^7:S\MZ3RLddX^FQ(91F>-8SF.b/<>JaJ^)M.\BI&LWE0(
bQ3II.,\@+AY@@b,_-P-36]32#SA;f27e>3J]C+@6PJX^bQg/8Of6M-f<e(V69J7
CdP3.AKPV-H:4],=.H:JXSI6G,+SSH1K8If]9bN8T\4F(aFd+MfU]FG\6Ic^]:&B
DD+F1RKM(d&cb0RI+&U)YZ-_fGaT9OB7OSFa&@GSO@BQYdI=FXK@e?e)CbMRF<Va
(SFQL>?SX[-RZR(>f#G:06,Q@N^F[d=6\RFF#QfTfB26+2XIZJ>M@6WI.SU-&QG>
A[5/Pe)_fM5#2O^]D3aD9,b;g;c1V<-7]YRc6#=#Ja=R[6=7J&K#2GADIBP)g3-V
>8D+:YKJQ8/>d->_Q4F6O.K47dAHBIbD(81P001@V\J;/8<?c[(\9T>.PGND7ZHR
9SXRbRSYfBJR<e]5ZSQ-C(>=G^.QP:1PUY_(1dLJ<:8K3U]Q@OXQ?5SAa8LV94e1
;eD3aUE=_TH@8]=GIG\@?f:(,_ZX7K.+;L+??R1a78YYZ0<)DMJN_Q8)X&53X\c6
A=_5^5G#,OKg&<E[ADXaLD&/P)R7BVR1cGVb/(9GS@cQGG.@49_>B;XS/d+JX4G)
K26<_WFTWS:C^Z(OTD<,\g7J7>f:R\0O_W;KJKKD/Nf]8+JG&?X^d>;3TCN274.:
3P)U-8-\SW=\^B^O=X7D=adPX(I[&3XARI,4^G4e<2F-,Q7OYW#&/P72?B(-U37@
OGNN]W5CgZg^XSNDSd/&C0^V]c9UY.WH-=[UdcOLC>3Y=fCf8-..2Zf8IRAL,I;\
0=[^[WbgK7P,1QRbgEC8V:1=^8^GRO;2\G^<_+cc@N4RWWOEcMAIW.\=&QM\80Y;
5&7gT2e1[3>^F5,()(7.b[XX4_=(@HFfS?AYGSYeTGV\&?cV(7#cQ10fVDgG3Z\K
F<^KAPNZc?]?0\^1S#D5f/,<^)9QX+44UC<Af?U:f0&DG]:JC.<##XN16PW0,UJM
Zcd6.fKa4R_c>-#[PCH:O-eKYWF\Xe14^9^g?UQDcfQK3+I5DFT1C1c+BR?gdFcf
2HDB+OTbb=FMXWDR2&#\DP-EAcfN[K,;71K+LV3G[<C4gK8MG2:<W0=]^LcGPXN+
g^P_Agd6)[ZB(\ZCOU_Y\4H,0T-21S3e0Hga>9+/VX2Y,K1<0F1?>ZTP[EM4#[V,
_A(_ODc;fY&Jf/_J6,F8c4SP<4G1fU7TSe(RfK5-ac6AR^4OBY@1e23gg;E#+@DU
+0KBLM?^\X47GWIA+75(/\(]RFYYY)HJ9KFC?Vc,CJ+JT[aJa;PQ=/##N@,F\MWG
6K1(7E=#dUN/.M8L)D3KbMV#g;),/cK.-Q9>^H\80Ed^F8abd0F<C]eX.cVLDcA,
bfg12/(c,,.9_WF+6#B0Q^gXEFZ^ee&0.0J7>bJ=-b+LR@PPNZ:YGeXb=H3SOHS.
R;RQREb3M^.OL89,)d(5??_2I?Q(CM0K)Pg0@CPZ3ZG31^]P0X88?3JO8O?,MC&P
NX@Z9V[7cFg=PX52@2USOI9DVP7,YQ[(A;]LGXU7<b;KDbZBQE6=JWMN8^;Q?1C3
eH:-+T_XNOU6;f1NE2QQJbPKX/MC3EKb#O[g1,=G6gIVE<R&3_Lg8R],R034dZMJ
]>N1IVVcK?(FbTP)0N]ROaKCZ#ZGY.R[VBRDe^e>5W9_.ARcB>O=gR=_<&U#ALR-
C<>1V?V1N/C1-()_WSd@0GD9b2R4=EEZf,c=Pe@S84I;Vf5WZWeOf2)UHB:IE3dQ
3RQ1[eH?SJQ12-^Q,DQ0S4(P=eX86BL.f6;YUZ@A=\R?O@J5.e2G0.H3FK>8WbL_
\W8K9_\/We]:+Ne@-\SK5Q[aQW=DS(#gM1b4FNWGd7<QZ-e,SFZYb2^BJ0+0H1S6
XXUfU(5f,aHFFDRYG7#;]5LQ02KNU9#6:HF,[=)UOJS-B6TG\LgdT@1Z(1CAG&:D
TNDDKBRJ38d\9I9gO=5P(VTVK>3;G.(baR8>aGQ;;=G/Q5dYZ/L2].[_+D7QBRa<
B1+(8J>MJc(7JWc,630cY\BX3G[R\:dNWE_VeRCY0\V=\^TeCEG-77;Z;N)PK,Ta
+HC>,[OK5g>c6&G>gG:M[=1H?\JMBA39-4TB(^SW?@99GZ<;=[9H>+Y5J>=W9g:V
]FN&GF:O9@c0=Z_<V^gS-AI-0a\8C2JRP[)fD6M@Q-+;-5LETBR:>06IQ&f@YY7g
F\E,E95Q?@2(gNE#^IB-Q:SDYXCdFY:(=GUU\FD^B>8U=,M1CO2[KZE,NL:a3#76
6H[.?9\L:-fgdW.^>f\_6O_S:RO5WgI>_KNYD_7_Ma.S0O+;849c.FJcBV98a(YV
d)QRQ?B+@MX<8&)9QTSTO\?.VGfb@0c[]FW4N:f]SLTX1PK4D,BB#89436V#I;_@
LJBCb4a_/WZ?XJMa,R3f-+8GF/FVGC8d8PU,bF11#YU5AB=^/C7_F=U_]2C6TPZM
9VEbR;8VN49A329-&f:/+6U[F<7VEdBFA@8JI?8D-D&@<ddXN.fZU53^RgX9E/LW
S?[eOXcI:NcETAFC0O(8a)IO1_(/4ZM[=LX]b_@;d3\E(5PcSIU<)b=P)([+aZ6>
B0/aU?<U8PG+NA,BUT?62YGY7C1UNF&><0HOXe6CQZ3GP9S@+:LGUI:+DZ;eYTcT
>=DPRb1dQ+@.2@5A+e<A8f.#e_C&ZC-aPNNF9:(]B<QC6SB3J\aBa-@..>#92X6B
)-.HTbVH9G[3_C<b;MBeP,,1?\,a#,<&6ef&S8]]ZXE3[Ua662IPP]40VZFL<>Q)
&B6B1:S\RSLP&37a,.5E;0+IIf\gU96_.+)/746+7Tf7W9T+XV-fMT9R/21:SR(c
f37K,e@f0g^TgcRgTP-:Y_f<8QGFLZ.#NU/Z=.Z+W\OT/):g7OdSBHT,FaZ6UL@O
ZSET.?,c.UB)[G:35U:2CU<>A3cE@W:/JMM.:@AaHET(KPCQQ/52@3.bRCTF6]CX
V=c&WW3-9Q:\^Ec@KER9XO:P0A<NW])A_=1f1,SR58EX6[MD3_9_Y]A#1FG_UJ[J
K]Q5a(T5K8ONQSN\;V\X/;Q9gbHZSQO]SDg71c_\2c@g&_KB5G.U@d[W[-eaC=K]
_[/f7&KME\e90If@.09cI0/88O\XK2e+1c5(EL1PBB:cXCM.P30g6(f;WY?G;\MT
R1#Zg&UX=HLIBG5AfSTZeZV]OTCFYUCPf9H2(77ADPEYeC]X+64R2QM3C[2UOd<Z
T1g4e][\SMQT[-d:T(FLX,M^2Y0]g7R7J1YEI8/:8+7\]0Tg6cH//+<NZSRfT.V0
JIRZa3,D6Q+gb)<3g(IadWZfOcOY@AY;/7XU:TMD@QJ<d/E]J(eUaG_H>3=b&9cH
#UN#5[L;BKJRU;W/;(9W0X1E=U?bG)VCC>2]3W_S-RNLWJO5M@J)TOF.2BE&RE1&
dc\+)beJ6&Bb\S(B0cW_VA0fFQ(H(=M_^;F?5I+8TZQ:>;MAN/+1OHSQYVFH+F/X
D12LXXS7J:P9:=/R[/YAaR=<0Q7BIFX-^#1I6U-^]#X>IdTR8U4&[E?VRLH7W[ZU
58+^d^K[AN^GJ=RMT-:;KFXTfCG?Qb2D6)K.P\Gb79EF<Ib6@H^+YQU?/N[7N.eB
&51I+KOM6cbNaF\XGR<V8T@3e:/1894B2]]7VB3(_72^4/e>d3,/ZTG,4F6f8PQ_
=WNe;/H2DC.fR@C_<GKb2e&4T<IBO)HPe0[/D,+gR(V1?V#-&(B?^H?\LccAFT6B
)T:]:LZ5EC3#M^1K,_?L=OaV6\K(g=1eFQUc<e@O?72(U5(F@a.PHDFB>cB/RYSG
8[319d#+aQV29,5[.X7+TG6T?TcbWLSg\:(-RBX)NP5[?VO2+8WW^,aR8A,]Z7(9
U-Pc;4Tg??>>DSXS<H+SW]YB2Eb()BI)@PMCCJ]SZEX/W-(/(72P;2\U;7Ia>##D
Nfd=5]<08A&SAX7AF79?([Q+,3bJ^&)5QXT7S\FaYJXH.4L^M-\bG0F+c</+B=PJ
B-cMD??VeAQ96@b,COD_c=f\)d_G7f\8GRdGBY3F_N2S1KT+.g6[8^9b.\EK08\G
<.1X?/.PA,E6A;:&31;,CN-^cG-\EP2#]f+ZAd?8/9ONPPYcc_YDXe=a4>2NK1J8
VMK=Z=\P[NT1E2H]HH]&+Z82F)TXPadU8a\M.D8B.3C413g&[YAT-7+B[7V^;0OR
:YBFTaFNXaO/<O:)ga?CLe4H8FaG?9.Xc79GKKLT9P<]M@T5J0R1P@@#Q+]FN>55
\e[8)-GUCP8<]L/8fLTXC(cWe]J@M[B[0X/;;(F)E5S0TD8\UeGWZLO@H#_:gXI+
53F)KX_-R,abbJ6BLDY6,@AQ4I6MAbe8T.2><L(,)RB<4[3WH(V\Q3@[HUO9dM9]
L[C-D;8Y84;YWC+b-PAH1?+((734&29,b=RT8Ia>AS/@O<W6-??M+@(@D6E_(R^<
e4VEWdX,9#GU3bLMQ(;QX;W[f7>28M?@9+YC6TM_2I_OKLdCIMaI?@Y\8JSg)IE_
6EGT8WEgIY7_53C@UF,BCEGW8H]MTV&X8e&_&4Y,-VdJC4U5^e[+5P&BW9X@-NgB
@g(O\A2-\)IdY4fTQ^IeYU_(KGb#GLRVKB79L;6WH1X_R>.RD-=N5d9XT8ZfC2)P
N@F-QHFMd9Tc1JN>e8U,g-H?)VM#LCQ)a/PJX#G(R>T2YXg8S56(a:BFc[6>9B[?
,aJE8ET-Y3QOPD][8.eT&<QI]ID,3KN</f_>2@^1E^X\D;))T11)Q>VH(O,U32M>
_FI@DB#f.+VO[EJ[(OI]BHeMHEAB0:1L:7BSWZ;:WQ5@2.]A+4B<HfD<&Z//WNAJ
:CIY=?\V)/6S4.D1d+O:=,/E[P^O;:^4BSFM]XM2VZB4-0Y[;1(ObQ<C_O>f?Q\S
M;MJgd^G+NMaH2M/U>0.M8_=QODAe(36\f6)A1:de<3-;0UIWFM,d+,GG>4Q\=g2
(@Zd1HO<aRDNG&ScOa_1]S]VQ]E8AW/Uc0+PZ7V,#0EWeE/5G#\;IC[YVg6bG<GZ
08PF[fW-0@#)C>f7;\[^?W\0OIPR24Y7+)2_Y.,<Q9_7(=[-]><60\7DTP?<J-_4
5JE/Ng7EHL_\9M4E&?3VN)Q-HYX1Og)c;IB08,9R_/<.ZM;_9fa/43SZZN1);\g9
TMO_.PK+ZY+3C.761/@UF#c;=9_HR?.5CS=)OMf=M?Ha+<_-eGS7R3Wed3B0XcTe
3E6=IF/SNEJIE1J@,E.^PcHP(/0LZJ#00ZgN:0PfZ-CFI2>dUCacfdNCd16Ve1cE
S&83(C:dS.QX-:PCR#eb_CRK,gRPIZX_I6KeG,ST&Ue;=Wfg(&96\4+G5e_(bc2)
.e>+^HE&8:@5T_BPFeeRVR4Yafe5IARa^E\9(RW&+Y>7Q]-_(TCc\J[,,3cS7=<(
P)4DIg#&RG42c63Aee,C=363GWEBXJ5ee.AJd3_Ac\UZ+7;(:7XGX0ZJ^\Jea/1U
?9?X5(/<bFAO4]bI/57P=_]/cMMK2N#.TET3\Y?WBXGT0>_RU0I(K6H8gQLf-I@T
_M;HY7=)<^aWNETCcS#[P+08&NcgY&<c],7YRcd_94N6@V)f.;D/;8\.IPQ>WNQ=
^5gf0[gVP0aAcQ&B&I;c^A?RD_RCQc6ET(gZ6ME@Q(4KMVB\JA0@OVV:=)L<]F+<
K6?)EPdS&#74I7/f?f]27FcHU1/I:b]P:Y(RE1FNA#6C(M@3WUJ0J_82&MSC\;IP
:&3-P<)3O)7VJdT9#e4dI^1N.2e(fG(-XFY:cSY#<N0BGW\b\7.fSa;[<>YKZJ&]
6TJC/BaU2+#(<84\C[5@+g9d;+A6E3Y)Mag5@:N3V9P=7W9a2T61X+H[N5P^>5?:
)B@aR+WdG3#?d\J(XE/f1Y\BOC(P4Q7<C1(:Q&LaJ&&1_GQ5YL;O[H5ae/=8?FL)
@B<X,..WY._AgaR0bVR-J35=FRNf@0-Eg3<3g\[OC;@e>A45_M-@#,UE3XQ-1,&\
(TG@V@U)R:,?@gOWV<Ha+0)_b:1EEQ.?b]:Z0ba2HQ]:,/&,6_;f=35[Y.^S4MXP
#IIfG:S<IN\K<g/8TXbI8AVB)>J5RAg[77+;],&@TE(ODH>>87)Q@cQ;(T#4M<+I
eTc52e9F<&1Wfb@KVB\8_d@1S8K/J>FfD[cD[AAf.2H7X99B3KHW)S]S33;_e#Eg
KSKI[^CXTDe#R3PAVcYFFDG1]2#1;e@ZeT65UV.4+18]a_?g8>a/g>;0R5:)]<)A
.:4@C39;C)+g0B+G?:(4#\([KT.KfISUb2I&b;+TOY0)0M9[O0GJZYR8QA(LZ&c@
L?fOJ9_M-3DF0&8AVV;V/A]C+MA(SQFKe,Me.SAD;B3H:=ZE:F.J4Q8&C<VVE7XR
ETIJSeV?]eHP]A^S@VP&&7[X0/6JLK@OKD78G063XY@fQ96b<-)H#:\a0+fg=]?A
F.feI_0].Q1OHP34deaNO8J3B8gC2U5N+H#3N6VGc@0Z[5)7E1a/Fe13V(f[:c:V
-5S[P4Z20R?b3M6WJ[D[Z&0._0OES4f#E<W3J#W2^0G@KBFOMbTDB>J4WI?YEEJ\
&9Y)_;4[[.g1K)=JH]^g<B6cA)+TCeFBc1Y>96\+7gMWY9J7,f6:R]51#^B483G&
)@dZH,\I_1ceC1TNK?S/bCe,>e?3^9b7#A4g^:R)UMC3?XOW//<=(Wgd7[fZ4=G[
]<?@Ye;=51-d;Ve@D9>DT&K9I);N#]eZ+EbHZA2T[V>_.UF:,X\R_YPfR_#;QbEV
d@&W+_CH/?S\6Jf99@-S5::QeHY;S?8[JI?dL)#[ETR8_#SIEJUP,G?+@^&_:DG,
E6=?Jc>VNQ&XNW5c+HdC2G[^)L)B^ZB><,_O23/O2,]SG9LXSf^A4,6P2/O(]Oa-
?LSA@OZdVU,AR<I=Q4M-c_5PJPSM?:@H-@WegcXUYL97RfeR_5@ORUf_QG5^-[d^
g=cSX,0XY-T7@X8J\A.C(H+-XQL,5;ZN+Nf>\SF#RH?JeZZb&RG5U2>,;6&Ke(L-
:7\b0J\P5P0YLc?.[D[c-=>S6PeC53CY#UM9DI;_.?^/aYFa12-faNFST=[b9?3X
NZC6X-7E[SUG#3<fI4D&VKC=S/X2&S1_Q-P0ggY)-Y2EVHO9M-EXc-IWV4QG.0a9
IeFKF8\(]#4AEdS@7cDd.^7.:2L2.N>IYR-D5+0e+Z5@2>(64X[>ZSZ@Jg?4K=Y-
IdA)QPQ46=QGbN&BYd=.K.5WD<R)4fVG4;#3NbHZ7F25JZ.)ZPf&C?[fB_(;Z,D5
+VXSbQ6efOQT7Q2Mc846)FO,NKC9;Q\IL+^=>E:>?DV,gDI2BC_RFQ+VEWOQMG.,
V&8F?^c_I>0DD:)O6.XW+^D<P?X=fH9O9D<Jc;X--SC0OU;@:UKC;(2C@ZV2^/A@
HW]d1Fgce?bT)+EcQ5</)eTC#7fE6;;S0Oa1J@f;#]^JG^#:BL;V\WBbY?^#]dUK
>]6ag#/3K@/gFTZ,,[?ODY7[W8Sd\f(>@[GNB?OF[^3SI=D&1-+ARJYM1,M/^;=-
2A<4:dS)95C5^9)KZM,042eNEWG9FY\/][d8&+Z[#,0>UA7I7@&I\?6LJ?>^7[O,
PA8?:6GYV3+(Qc-1/aZY9IW8eG^M/gX2[M6T-K_d\>\19\5bN-cX?H^g6:PUKZM3
g0P4e7_ZU<TY-ZK-YBd0\HF\0EJ^gDO43BF81J8g.gfbK_&0_&f\P>45,F#&EQW^
?1I4;92O(e+VcgSBPO:D/)(OXPW^?6Ed.7Y?4I/>Lg87K7Z?g(VZVTeaWRHa^#O)
?P(EM3+X]Yed7QHAT90#FV4BDDFXF07\dH4@05b>Ua)bTPP7Q@PKD_QC)WXKUQ#4
Xe-dfDDZOcAOA]c6b8^X>cd_;V0EX[VeQX9?b[>c,74^\^RCY_=eD^I.EF.8(bKA
LF@KSUMTYa-eY8g,#SZ3SH&ZG[>DHR#1^OT_5)^?9.2)M38<[O:a1CCd.4[1]\7<
9Haf#PSc;dbPHH9?R4dgRW;=+[W6DP)Ke0Jc2bAb2:)_^b;Z7bC\_D?50D@]cJLP
A9-gV_Ef&<_-:>POgD]OF5ce.]#KKdYgBa?M)cZWP-1)YXg_gUX-62d>94B8:N>a
L&1:B?ab^N50#TM\AL>^<Tc;P/V,ZG_dJ.eNeT[8LeNfZ[KN8_5P2ZQXIPH9TZef
\@gYH7<-Ra0R&]0UDD>g(\-[(e)M<(140C.CVVTAe2AA_JPcPZA15XUUa5=BP<OL
2H]07YENM\?;;Uf+>\@)TS&MI;CacL#;GR7X5.<X8A,cHVGK/<?aHN6/F_C0AeMc
VL]RRC6Y06c8UNY16[B-7MTDN<D/3</DEW)&)Q:NY;6FL.J0eO\b<;,a]9>QWc5d
4M1]\_GZag+IUT,=b^.]e7.d]-ZDI?(;,I/d1RUeJ;BN(X2N>>7FeEKLc#9.[9>+
#.B,-TN192/42^F94CJ\QFa&0Y2/?g=;I7_[df.@B+A,_5FY/bUeM=]3]RTAV@KD
F86Y&&<\GN4AO=T[(WdEZR.N^:ISR/KX?VZ_;[g:Y)EEgB3_gf6cR+<.C?TL,\8A
)V?VG(2CdYV8&;2H.g.(4Yb<HfS71?(K,HW=fH5fA8gQ0QE;YHDCA)RFY8+W9)gX
WcM.f73>^5T:@9]Q#:T6UMG&&W,Aa#3=Y)R4,BQ58M93LU#.LRK5Y?JY_4)05C7/
6-)Z03<XU9(5e,KW)=<\cdX@N61=Of;[,&T@B>-\_E#M?bY<3SH01_7D4>IGW:NA
:=V[9(cfKN3T8GL@Q(>YA_M505FRFC>P/;8<.\IB,-+?40&+G[1R05S?0I#-WD&0
<@I^-U<]+N9VTOP#^e/68UX^<R5->GEGS()KEMRFZRJ&.ND##M7fIb2061G4(<dD
fRA[ZU9d_d=bS0UW)E_Q)DY#]O2/P\dU.@P]IG>07X(-((He?E)XYe#5dW6LBAdA
68bQOKf?Z,DA6D0d(V&V=R-]TAL(MINFNX97&&+W\MQ?C^6L]3Y^Y^\DN(<NSS@X
-Td&B?VDQZB+BXc?=[a#_I/-YSNSW52C#:;IOD.O4OfA;<)3T@&T@NYS[a-.7R1.
?^/,Q5g7IR0@6F1MXcVFAO\X;=L&?=aHD-24:V,_\TI8=d/?3A2+M<K>(?HQ?,C(
&I-b>1YH:/II9+BeDd)Ud.NF.H)#(S8/IIdHfFGBB(6SK-f>ba;<Y_JN0FbZ>ZIQ
aLTGO3Ee\,Q8cXES/E4FV;)W3f=._74)>R.P;^GN[&3dKR5a<]Q5MVKIb#4FIYb5
)@_S5SP.N^J9Vd+:F6gVL:5<PP(ZL6_SB+7<_/+[8S5EE6Af+c;PIO)O?bP_=4BW
1Q43JX).F(?2T82,bNNKEgCcS34dc;9?;,Y=@7#)J:9c/B<7H,Ub&K@M\GGa^ZC?
:).E)J^QL(T2KG9#Q94aO-[T4fI_GaHE=?Xc1Z(D+=31&F[MRW2LbEd+e0ET2E4[
^G_OB<\OWcE.K8.3fd-NYXDC4A&LMI&U2@._>4AC&X+dPQ/ZIM.;1YG6Y-)EZ_>W
)fPe-C;cDP\=7:-41E,8bgQ01@=3OIC^W/fN2\XA8=.&9.\&^QM4I9fg-V.@]D8=
dREFZVBX.OP[-3HLR#MVM)D=/9OUa_6YY4(R)19[R^CS^MK(dVaYdR).9?eW,L6>
Xb;_@gNY6<FcD</(XIM]:,3WC\b>+MH>Y=V503I2^_<g0LcI@?8A8BLK#<N6Md<^
NRaB5agWZ8Y#E38CY\Y+;gS(]K5VS;fD&/60G;\(.-B\-9[8Q^@IV)@dVB_b0LgY
(I98^7gg1gRUVJ@]A-1JC0aWBZ8622\(?69RIJB2^MRfd-A-E@W6R8AXWg2D\CQI
8G+P50L2TTZ76g6]F9EG,VR6K,a/eARe^/.?baFL.6FEd#4Be\+M>1(U3YKN^9@5
[aN.CO1OVbI1GB37WDT]^d^.^MZYdG229^2<.e/97@S4b0b9K5KD.=4VN@@ZS=Jb
+BTQ@3_BWOR@c0EWI>U5;TQ\eg0.TR(+=UL0763.AJ>[9XZga]2L4<[JK(bb;\>.
)ZX6IDYQG9^]QNH5;=8/2KM9Q1/WZ0b^Z,YfY=-=;OR+\WO<1Q<)AIVRZ\.fF??)
^F8fC=X9XSNG(K]K+?8aH[X4Q.,3BPaD;2gfe2HFYZ)YWJI@cc3C@A:UeU0,)T=a
Y7K9C90Y2G2(@4S7Y\fWdNdXXW&_P-.Af:]]]Y@8>)VT7KP]7HJFA<c#>IdT#W=R
()&4cgSH^Eb8fd9:_R_JU3-aCLH3ES,=:93c,&:bRD^(J@DH7BCGI;((VeQ&;<VR
OO?@][9<R4@fV+fZ5SAdf7d<D8bYMFg\?@#H@ZdQ-d>;TC]CG/?0+P&W)eHZf,C#
CJYd8]ZRNd52#^,\]&]LNc@QO;)&?]EPE?/D,A01_-B[)5U15KD.D4eX)>Y>Cbab
[.(F2\,G/9C#&.@^fA+(.>S7W+2cH.d+@IBMC8Cd#^4DU5GK5#&-M3PG7Ma+Y),G
5-S8)S^_U\7BFWVB.2BZRWWXR<3Uf?H@G1/ES_e@S>(FbO?,IgK?Y[.\FRg/@.,,
4(67DbM,F,OYTB9BYFN@(a#&P0]8WD(e_6+3,;E#9YV)4&38^_[b\=5&XQ5^C_bD
>]df=c8f8/cb+^G4]RF)+/,Q9Ag4^J+=a?>.e8VKdVZYGaH>X-+07K0Se6:W2B(0
&31c9VFT\G/X(:8NAQf5V1+TRMH]Ca^235WC<\Y8J&1-Fae&_2CfKUKD1Q&./)O)
_>@+M/Le<:0T_N]&^[)dL.<V#<FIZ.58X0_b2T8-cH=]5Z4I8g>+aY)/BKTKFW<_
OKd923UR^T1gd26F)8DLD0(RQ2Y^TgT^J_d\WQCWNSA>#6QTF@>W,W>?C,P^[CQ)
)LG+@,1FNe.\]=cTMQXeC1B82PMPR498:5Y4N>KaNCY)5.G^?F^&O:P;YKEc5_ba
C_Ae+)Yg,G.XRXge:CM17[@=_L:M(B@7]d.YIG=/KGUa+SG]&<D=?H>[CXfOb//;
T/^,c9,9QfER7ZTDK)7X:KC4AQ59T:;Q5PF#@2)L12See,DSKS(b)/VGY)@\=R:Z
eZK@Kf-4cEfSA+>R@@ba+_2McD#7XU9)?e)4?)G3TM/)#PfBXbBcfSANMF:c&-2(
E5ZPC=[;M9T7f3ZE6V@MDJ?ENW(PS:LFORC67H&R0F]=,DOc7O0:/73gP:Fb^UT+
3T/97[fH/(HZ2N5_/[g[Z8]-G_&:T7V1?(K9<9/HWC/7=CRE79A/JU>F(#6#e21g
@PGX.UFLV)2L+#,9DH3H_C8/J^-R<1ScQ>QXbQ+KOI/A5P8=PC^N,\8O[4,_G6[H
/cEgg5I(ELT=;=Y@eI1&J=cY8Efd^Lf,2U_CX=g3C-I6PL6KggZbD-d7\_MXfA8_
[#EA?;TJNdVL,6/UHA-:,_I#K8<0Fg/4,T^/()))2/P^)Fg,bF\89CMgE9ZR&AW=
e@JP@0DV1K.Q@H/MScaZV&bUA5eWZZ^M/3IK1]R:BO.=\2_fIU\/3(I\0-E]ZFA;
g_3b+4WL.PKdWf.^9(S+Jf,@J+][W#[b4WaH\g66AO6:B[9Z+CO6:N;/4V[\PZ,4
D+gQUQ56ECAD;RGdg6BQB&V_cN@6?2F0517.9\.P,64dC@RCC+H_T/G\P#>09(W3
5&^LZWUB.Y;6RE4)Ie#0^A6KD?A=CC;S<;Tc&H+C>dFBfIUN6cUP41aTWUdA[M58
UMa(+H>ARPA8KY^^I<6_K11ZSWGA/C;:Tf<VS0e/Z]7S((Bca&Fa0DX-_P+I^?6@
H1E)HRKZG(U4JI314dO^N:Fg/<I,_B.9_ecQR19Kd@Z85.CU+9<3_(G;,<;T[L/g
LA4EC>^W0g\KE:DKPBR_NY046Z.S)/JB^FJ:FH7^O>@))SQ_fX;#ba-^25;ZJC:W
6Ld8Q6F6@R4\_>eC9P:\6WBMOf.K)L8W7<KX=].^f8&6OGH)?5f<KM,ONe345;gd
?CO5;V))NDJYg0@Je6XBL3+16GI)1cC4<.fT6AHYJW.M\Z-Z:4+@R8fKP??RR\&Y
.=e)UA-YYR+V90\_3\SfQ5W6X+\eW[)Qf).(M\d_NH(H5+e<)DO9&F-K:/0@;(OB
=Z:9F^>;7E3RDP)&@V@FQ,II?e&PRNWR@FQ@[MCFE#7[a?CXENMVf]RF7fUQ1LaX
IJfEH6:2EK9@\O=Yd7/bBgP@f32V0ab^U<g_UMW+1-A=Vf8-Reg?+#c:c:/NRK\[
d#;Q-bEDYTQHYLC&/XJ/+BX#c_31H9@A2N72Ng9\:&\BaIb>E[UbR0#W[D?7WWgY
f0ARE+_>#MGD4UAWI/^U=45^F_P&&]#(P1BQY=1451OFY>/4Z]9_?eGANG/,GVA;
09(?0S7+K,FcIZ@(F3-@CW^_&U+J7-;d.d;/,P#3G.J8H_,BL74-06UZ]Ac0XQOL
RH>?E4(9>,M]P<\;&+ES9^XL7446CB9.G&EKTILcG.H<L0HJ4PA7A&Qb+J?F2NZ[
cN6_YfZYTEPe4<M?UfR.c\,313#UfbA?a/R856cX6f+4#-QEU6^4X5BH7c32e<#P
J0b(g=\FTHYY]0?bG8V4+Ed)&1GC47LTGG8V29NM2Y)-O9?R#YD)(?/M_a#@^WHN
RY^W/03FNOCU6U3eEf4(a.5e?NNJET@1462g_4_#[gUK,HX<>[MfML])P[X+eJ)A
;L@/L<=&0L>-++Q];I)-6H/F(ZD2.#\&[\L:=g&@FKNa)F3fVaY.7R1,JZHfdQNR
E]dC7V6eHF\A4QJISP](GC\H,?SaEXGJd?9O/8+M>J)b/_U]M[8S28AC5Ze+UK(#
)Ecc@:#S&PQ,W9?65(N2bNHS9_K7ZH&5?/5+G7X9GaBZ)I&=XG_[;0:a\<3?9NKB
GJZK1e__eI/(F?2BTXQ1HST\&@DDJd_d[AVc[:VWZ6>Z5>R<=cZBDY:&KR?,c4_2
C_R=f#b?HaLN&G8WX<ZS^9gORCRO?RD9U=d7W[6Iec_\)K\KZ&=eJH:)NdS)I^cU
AXB)c_A7,)U;[dPURPA7JXO\&1&0D\@bg(8Ua^dUXHe1N8V:]RREKIGB4cL787:V
YdY8>fgXT=KeBDQ_:KERUL,DZ75-P3R:L?K35Q2OAUaE:UBHg^1<.a^JUZadH,K)
R,8=EJc6GN>QK0;JYZ<+PfB<36M?,O-47dSJB6+FF;H19MWG+cL\)^@N/.NTZ4<Z
#?+7@a?U<5#560,S?^:XfSb\GQ?.(YQ.fI):_BRcHT>cL^^Eb/(_19d6)0_9PKI9
NM?4DHc3gAg-&2[84LM-._a&eTLM>V)-]D4]gKA7;F6cATB:IgT.TWN2E5;&#8=P
ZV&+)VBK@cF6K0XS#(2+LUC?1@?SW;/Q6H0;=5F6PQB+92OW^0C.NSUZ?b>4FO&O
U^gW]Id8+fe1@-MM/X:\]ef-3JD8E/bAEbfee<9??7FdX(B3D8W6Y+e#)@?LOR&N
>-<7>]+OeWfB>267B)YTW4Q,Y]27768aX.^PZ#>#F7&LK5g1]H??HFUF<Aag:)H1
S=P1+K8I#]Rf48^S9fA8LTWW8,M<E+6_K],M.9\<4I#g8&b[UC.R@f1OMFd[:?>#
#0XW.,fP:A4V)B@OgdIgd\gBNG1Z2.ggb1_HY72)@\2UL:^bBI&TGC5],RS49:B(
^Y=U5G_VL+>.CJ//>^>7P7\/97[)4<\@F2ca^J<Fd&R18f@0CATD+/aSfYGd=J=Q
AV4aB:F8_3VPe[8+eFM-HT#=9QcPU,3DR;+PW<aRJ?A?9/[FdCJH0<DGJ[-O(?c\
cKQP-+YeT#KNGD/;UEKP5W](gDVT]?RPT-Q/F]-\R?Ob=R^92,9D2^>8P;55IV.,
84R;cDJ.c2^QT_)>aB:?0>1:=Q6eg=Kd;TA?GNDfSTA/>>8g>SF2d=_.fEaBS53S
R:8cN-K2<L]6aW&Jd,0Sb?QK0MI/RJ+e5(V1\591A>G3RfC>O\a(DHPRQ6SS5I&&
ac(\H>3A7fbc,IEHW5>eK6:EbUa;4Ka\HQB+2Mb6O7aM7c?X/3K[(,&a3A2K^ZaI
Mec]b8d797P<>+d]Zf\BPI_5+ALFN/WUH,64Y\];gX.g(-f/f5ERR68Kc39A,Z8d
Pb(dC#COCM:NP^-,D_9Q=E;bS)[.:UF=N]bKU=8<SfV7d,C,7-PQB:H]C4]9d<\7
,>L\fCU0.e=aU=86\?NHB#F[/E^#\+V)@2@2Z_(C9VAVd3B95/ZF<]X>>KBO5@XE
+?@<A7JH89G9/MY?_L-PC]^c2L-Q5\dA\\P1HQ=I7B)07_BF36NV.Rd9+7X5A[&R
2=E&\=V0a)H.=8BD?F(6TIO#0cae4cZH:adg=X6BA_KT(2M5A?].8EffEgMY+^/d
-VLNL&7V[@=(U^HMgf)\TH5BHe)2]TF&(:JQ4+@2F)T?KK793XWTDVY7aeA.+T-e
N->=64b@CKbCb0?MbGfDRG]9I4H5>R:?g25KEE,V?9GLAB&Of/4UE2G-cd=,DXKT
[WLJ^B\:.H7fYKd(6ZE0L2VgBb7?;UQ6=54d<Ic131,V1aC9.RQXJF#DA;=OeE+<
#-8.GT\+@6=RLLEc5C[/5.DADK_84>]K4+QXZ1-e=dU^84GB+W>WecH)/KFFT_-#
G>[(]?U_7[2H@Q?9cR1S_c9@/4?aaCC>GE+GV(&O+cGMI:G5YY60LQe;^d]IS3EK
\9[B-:HW&M^CIH0EP\VfC=[1Y_\B-]S&AB61&GZYV3\a<?:&SP;S#E58X4+I>\6>
#@)-K1&764GW@,9B&T6T_FFBJV&F/VgJAeRE74Q1b9Z23M17EL?fLf2E[;8A2W#R
&X9JO-_3CC5&UR>=T=:RJc6WTa89DJ1\=AYK]gLP&4gbNXIS4S:.B)N0?>2M>Q.S
K):BNW/FCIDb.)>WF\N44?d3_QV>VQ:YO#^]YU8H>:+/fHY0QCJ8/+^D2K5M0+>[
ZJMZH(<[BDVJE6:5KBC>f_)I?^;;/<A=EFJ<Q.Q\^<EC-&A?E8\9<QI+&b>/U2T;
?g+D+/5)N8R6gf4(_IfNTUe(f[39&/FZ@:@Yd>df^/IM68D_?8Xb.T[SY>I#LeX8
@KT2[,\.8M1)?/W+bM=>?&NBQS-c_L0M=FR5=P\T)K=<5EeCS^CR<VO4L:PVR8\.
C;Q97)Nf//dR/f?)<FNZ^g[0>-2P46/WA2ZX9=PE:3FLe87NDCXVO39KT2.3/QEK
@eDYSZ<C?be57>-P1fLQBU9+=3JY9^?K(>0K;UfC4_>LZX1ZM1JaXG1E,..Sf](e
US/<&;JDRD-=Ke)+:XQf0SQ62S2YOB_Kb[PHXTI?YegMX8P&_8:)M#CQ.:?M_[IZ
dK,:#_F7)>LM?GHZI<K?Z?adAba1LH5M8cFA1N<dJ<d.T)@\IeP+A8B5:ObBL,WW
]d&B#eBc4N,HWM=U?0FSTaRaeCdMM2XdV0RWW9X)=LZ0I)3c-;[^SdNVgfLV^J]W
,:f\Q&.;97C9+S71QL\2R@2PZKR,a+gLFQNQUFc/??&GO33Z\2[I+@&9KdO-VR-L
D0KS)\4W1U8:U#aAMZ);ZA:3:8R>?5<WUXA(73H42^cWS=UGfSAf1(.D#N)P7Ne9
_W[AT?Ud=bFW1J<Q?L?Q+WAWGe?&&9C:O[74[?12c9BKKPF)bY-+R-,L9)6d11Z/
3B.L8[WBT?df;]\@dF+G_@T_-Sa)M.->_IWKD\cM:d:]?OaW/PdFPc4(,Y?6^Kab
0FgGL\bZ;CIaJVX[RL9S)4Y@aR-UEcfS=P)3.AU9.2KGKW)?04EXUKN6O@[Ufca\
g@D=9Y6cDVJ&b63G88OQe/[TfLZ4)B;^JXZZ\4V4@[ecV@R&&3S-J)V\&\;JH63T
ZXO<1a[\g,-Y+aPgW+,b4=JZ[+-GgU#@<efcDe90B&dZCDZ@Yc?G..(D4KMb.dTG
+DEK8L2]3.gAO7OJ@Ab)RLY#26+ZL&=Pd1YH>Ea33[,B_9K<d1LTH^?^?],d2.X@
S&Z5g(326CK0>0YL_;79IPcMW:\&_@0==]KUXWYN@;720fV63E/RM.0eNc;^E4>Y
_=a>g?0_:3].[G#:SLH;F?:D]2;\@C?3B=0JDQ)X(_Y_D9=OQf6/#9aETG#f+K,3
cM<HC.J.gPW4.5]d7/feJJ<b4d8;_L0N1NSgUa<6SENN>4d2KY@>S3-+N;DHX+T0
QSP+.44#&&A0FNO[f6Tbb37:#(U))?=4]Q;F>(_CUE/R-82:&I3^Q5e0c1B>LRUf
L@=JO4?2\3K\-/0Hgd?6K&_bCMY:cP4JIN>7Zc/d9c2BHH0E3C<=QW_6[9d7;S0-
/:PZf&bfPCJ1=1e]7/7,cgNY.L9YQJ/ZZ3)OZ<7S9;+VOf:JP2]>#QO8He_7c\1]
[M?-(T/7&<#I[FEO+]:7)9@<f;c]&?E1KI+/+HOa\L/-QD(S7aUFRM6Pf:5@T<f9
.G5]NBCB=XZVPD#;)&<[UPD6KO-fA1BcZ;=Z2QC#,4]3Q.E_M_,/Y]BV6>DUG9<1
gC+>#)2XG-W9U)X1;#+K.0B^6,T2^TQM&^8Yf4,U:3<K>g.=6V9+g5b_7Ag0]\/T
aCX/QMXHM#-KT)_KJd4VCC\<WE)2G8OES#BTRe&((AQga9,\afM:LS0R6eE&L;;I
X\0a^S1GY7\#=^DHZ=;AU_eWG76=fc;2W>D,&+XB0MA&.FLe,We9>A[4,YYU0;I6
-Ra0BD3)NB5=<aGVaR)Kb@7E6V5G?&VS6d@1&G>Y=;,?OKUFC8>\>3Rc2>[@H(&O
.D,JD0NL0#La\56CX6^&A)^--@T>I-TWEDU+c?:TOd/W<YfO6T8MY#0:2=4,_X&0
V??+D];ZQ-\RG,IEODA@6McBJQR6M/5>W@^LBFVJbP(.1QVAD.A9U5/fG_W25gJ_
DV\M;OLD@(_QHG::6^2N+E@WCDQ,UV0fXcBRM)E6?_NbS^><_e<)7Ie=C[YC365T
P(WKPR]M8]e<IRc+BJYXXI)&2/PcBecC5Z)0E6^2<1WUSF,J?:8\VHSM0a\<[G//
;17,HJ&?+,=;?JK@]^M&C5O0&MaAP9\&dNaN[&BFWP^_LM+b7B+^_D;1?=>PP;K?
MJ_K^RS9)=7,/V?T_>@F)/-V=L_?H\9E)T_E]8BdYW-6\D3>cNf3;e1?C]@C;HE;
.1)>]e>^8e0GVf>8D]BbPGGN9&f>JL1e7CZ-6GPPbY#HZB_e2c]TA(Z[Qa4UPFTR
.KTg5d;H9D:,Y]b8?]&9OaBVEKEf@E]X608a3QBCQH78#9K_\ZRa6C>&.,2MC0X?
+)T:d#Z4]@4D9W6Y)JY(Z:,-@&K96_XP_f79#5\)+9d4Oe5e]C>]M4d0gb3DBAZ\
4)&BJ0cV@L?gH(&I-,/.>gO>Ee4:XQ]@Q0/MQJ]IO,dg&fe<DZ.^49T-I#fbNJ0/
&.b5LYFa0P/N/3V?49)D1>4/_1_N#LRNAX#9a<Gg&<IC8AE4L8SI)1];<HX2ODP[
ZRYPJ+JI+8D,)VI]+0R,=[T_+G#cV2[)a,5g3Ee@:G1=ZXfLT0QM(JG@_g9aLcU4
AdgX8S+EJdTQFdK([=Gc>_^7FEcb:W^GBQZg7e2d0C1[3HF:=d1;D5++S5)NMKI\
JCT-T3a?OA58X,Y#2\PK?^+VCZV[-K2<>8&>[]-ABV@5ILd[McOe3A3]CBMc@-F\
Z&YU;C5#J[dOWCaY^.3;QKGS7G^S0(@bNXM5X@^&63.+E=1Mga(DHa#dY^L=Q.64
V]>5PdM62KSDXd<[D0W80QA9JY_:U7BGE[H3PL\eOI,VX[=QMMI)3<HNS?/SEEV4
YT1aA5Q=)(LE.P,9IC+7)dJHC5T;O[V>1H>I,UI=c\]E<\N4PG=3AAdU>7CeaSC,
Vg.]FZ,\0-Ga=a#HN?AW25F[BgW3()J?8SO:5M;MX2]4?X>X3SQ4D+eVZY7e7>?6
RVBKC\K;0L^WbRKPHWN<Le,,;IP/6?FM<X4/#?[I&L&+M>75AcbIHeMGO#5JN:Rc
@a-,A)4<8T]&cU5-ZPW\D+A2K;8.,FQ6/\73C0:).2,[X75aESeIL+[L4@6BFLOA
UQZgZ_BUG.Z/_8-<:PE.d.\/(8(AV<31gG>[\U,/3K>2K1J0Ldg(OOd4P>X)2DM=
=^RQKTB;]d@+Ac=@G^ZD6A_P?U_Gc@Z,.NJ+#3aTQIfFDc<6N?6B_c#\Z;=E5HC8
5dZ..C<+>3)85Ee,1cG(@X+4c<A?A\AE[/^4Dg#-MMUB<YWMJ4/]?L2AdbS_P?>3
(0We5dLG9G\2ROO,[A[SS\_R3S2]G:;6eI+Cea,=aQ0B;AePI&-&X@G1YSb]:ZWV
b;7SZ3>OW0^)+HefaAY;YHHDQDHDC6:Ga:8:d:,B:BOVV/E<Mf#KDa+,PI))O-J.
TD)CY1-Jaa)REfSgO6M#9U@c#S>C]W>\?&+02PII+8<5\b&UNL4J.#eSa4MMS,1H
d8@:,eNK#FG@cg(Jg:-F4b=H[D>dYS@I\<PW+HLAHK-S+2#H#DX0TRRI58b987e9
+g.a)K3I<6^/V-.THBf&0[X(?F+R>I)(\/BP)G#8c5c(?#^K.bWTAE#?]fRUS3/Y
>[6aYLDS43(ag06FOI^/-CaVE:9NP#]ZEfR1[WWc/>)7^gNcG2\B+=fd9W);d:P+
DIPe8fKbXKJB)EMEK4)OY)F@C9LGe(T1ZOG\dRC)MJ2,.(0DHYISQa)E/f5Wg-K?
],@]<@4D<)@&eDH-_?>YEDd-BTVA0734ZO@ZcE@Oc,[G.GB/7g[a>L2.,(.S0G3D
fJGE\2aDK;dUD1eO^d,+2=<FbVbdZZZTgZ.3350CVF:6UXBe_K9+DI>dZd,fEbC&
^#fJL04Xe^6TZc9e2\e38c2dbM]?<f:C,3fOZbg00UT,LQ5QQ=-Y+?(5&fV8SQZQ
9T>/C]<;e?T:?\;-QASR1DBJ?@@;T3(6aG]H<1D]S+Q8DA=8UBJ3//X5)I:EIAHI
K_(a4@\#\0WCW&WO=S0Rf8X/K9K7B9E^T-DA1DNgM9\S.eaE8TJK=2V00/e]cg:J
AXJP<PQd?>S.\ORP,:9+_eV+R0/@V=7dAaO)&6=Q5?E(I9Z?=BXI^Q^-:T7T^<J0
.B/V[)]SV&.D9;.gMfB[7PB]U,(KV30bcP;_CaU[gURW;W7IN3Q&aB@a@:J>NN/;
W[6\6-3MMT:?@=0_IUSPNS=<S[SP9(dLR:D#AE^>_GP&A5G:bY4^I78V1/LXS8O0
<;@_#CaDLUYD5;)4gNMXLB=8ea:MAb1dS&G/WI_RIf)H<J\C>E#W6^]6U9LWV[J&
2FJ0/\TWQ&3eAU?R9QI(.A5Ag?/a\2;@7LP;)BQ1?UgHd-UJ7Zc.#Se2)]@S@U2C
^eaGEH96gWb6=JcH3I9I+TLU;JbgK(Q<8M-P,1U.7E7>ZTX,;1\IB4TC-4UD?7.\
F<>f^XQ1HSJS<dDATFbKI6+Z5GX6?f6=G@M>;V.PYa@K6T.PJV))BP<5?61X4##b
3S8H.FIF[;F66>P[]<CV6:#WL._[AaK/e-2_L-V8>^_0?8;/1<g[.):>4,/;WfAJ
]CYEI.J_.L<P:+b;XX0]=>a:?9B4T@TK_F<Q]c,I3fg]<N[Pg2LX^EXKU-I^cIJW
:E+&&(T8U&)GHe[b5e7H_BRe[9_^O^?0b1G+QNF.R\+[eR;G-2_)aC\E5\W&Dg-G
E\6<(EIAZfHGWU17I+Fb8bQH0aN@,WAD/C&<R47OI7LA.<3&LF>9B3]968bf2=1G
2Ja+^2EKe6.d:G\]b^3N3W]QG1_@O0<<R8A@O)TL+L>50cQ[X<3<OUE1b,/OOCW1
N79EJI-(OH:)gP[UgG:e,_\+.Ag@JPU7JF>C/XgI\aP<P8W]^ZV6d3D5^^9#/C>C
7^:^M#\8fV6U]eHSY(J()Y&FWVULg/eU\L.?2C_]7bEE29R;LRY.CXc:1&.)OBa4
:d0Z=+8\C1UA^a5^X.@#&1HNFJR&SIJ]+@K[HT@aGIEIZE8GJf&cM3]^#UI\__CN
MSdHMH2)e&635I7S0e>R>Z##D544-D1QVHA-50R\32Y_Z_U;>)A+E#.JfBA?:RPf
[@RdL9W/=:A>?_(;H)>VIV;KaIB^NgFZZ+H15Q3b+J(fJYdL&^5a4e];gLMVK3YP
I0EHO.6B#S01K-Tb/a?-SRd;#T(L?UN_2()XTZLHgT6+<(TW@>-Vg>T<Q)L).V5W
ZRO\>^G.R3&SS2/#,=XKR&&b_-7W;SD<#g2dgF\T-Q)H86+E2RM(KK:8>c=(SBNB
g3S,]/MY0E3a4.Q75=;<4L9B5-(-gY0O4?N3cb4JBVB(K#^VIV60[&CB6^YZ;WNO
Fd&W9Z]/1Z/W<OPfCU+K[V=cR8=R1fK<c[KMebGPR=+3gKC,/S=45>85C-+IecDM
9=;DVZ)^C2<?KCD6;^5]_EW,DQ.J^S?ED=)-1Od^.ZK=c326(cb?f-7)#dM+g)_M
Mc>]C9G,a[)YX(T-VcN/3=;TBCEFF-MRM<PN/7)6K2R.BOW+a6,@J3?>&K\NaQ+9
4KQ1[(-+?6IRI_f>@A^A0,<^MS6-WaS/=[RVK#P_R8I68N6;8/QP\-5ENKNQ28YA
f_J>=>17@)TN^8Z2@>[c_1M+MPBa8[>ACbVG5_bD[fR</UV&QNIPQda85IAX7a&=
.,O_I2Xa.(eU#=fVN1,QeYUQ33V[HD49OAMN2>gfRYT(RIbac5Y;SUW/[;TLB^[C
U4GJ3O1[YZ&P2@@91/C@2f-0)Sd.\+_@^=D.]3_46Z=XD_6T2[V.N6@EO([Z.SXe
d^\Ncca;[;[#]Nd;e@5P\Z5CGgD=2D?EE@Xd4_Vf@Yg)9+-?(X7DGY7Y28Y0(/>;
:Y,g&Tf]2Y-OO--;(JFf]=5>Q[2e(4<B6X8Ta9YSY1D=b<,Fgb,R:OMMb_G+9ILO
>28-#./-b^VDL5(4:Z[W^<PEN#8a,65F&,QLId+a;5Ca::41#QLW2TL3C+^Yc\Da
F1@BYLPNQ5G,d#:T-X6KQD[(]]G^d0SRO@95,f-WY.=D1\RFDJ@[U.LA8CeRE3S1
I?_N275)?b=16D<&d03LaId<<=a_]N]DRVWMTe_a1J7?AH\,1-ac@=[TC\:H_GI]
Fc.MU-;;T.>J9K@7NP8>TE6YPcQRaHP8=8HBXL(g_cLX/?E,76d.X8a6eSU3E[c-
7QEL.Vd=[dS()KSFX&4N]N#^Mb>JdBRgb@ffZDb)1[YV7bGYL(/DBDE,f-&eL+/R
F8S3EHfPROOe1KJMEADMJPf?2[6K+^#fNH=PQ6eJ#.EJ-)f;/RDM7WJ7+BV??X[5
@2KQSD(ZfVTPKF1G<T&<U#;&W>HN8FX_JG;U1V4N;1abH0fVONE65.5A#<(?_dHf
?IH&6U>8=>BFeJJ+DLD:M2LUf-EY,4I]O09+XN,#[X9(_CB)f5+(/g9UCP1-ef.+
67W@E5ER1SW.^J>g4U+;@aZ<MJJE0&@Nd+]L7>\KcLE;DH^NPIg9IU\@I67DND<E
VWL085Cc\\->afBXId0a04eLZH)D-3X@]NdXKXEYVKM&\bX@;=R&/+?1W2TY?H9F
6E<Ned]Fb9P2@27e2C7KQc2T((a8A2^aL7?LdL32Vd6>-FC8cOg?FHIYd26a<M#+
<d;?TWJ:O8WJ@^_[G^-7T1eA5QX.9<=1MN5OJ[Z[(L/:)(,AI[e[(;1CPO/O(0C/
a/+<XWge5REMR7#;9AN&)I+MH+E=P_A#:1/W&2G-7^C>(#QW[?KVUT@SHUc?HcOR
Qg,2S56cJb,B_/S93Z2X\<N7egT0#ZaYT\1::#]YRI(.7c8K6Z-<bL(CY)R\K1\f
(7B6>59CRJY8EYRQN9\[Q;:Sa;0?M5U&JF@4L/#9EFDPbc)?bMcc-a2G]X9W]=a@
L(SU_HIaa=FM&5C,g)FPCRO^LaWdXP&JQ5LI<F/H=^>/Q)9>:@+?7^O\?LG.E7EL
2;cR8aW\(2?/DHUF)fPU(YC;.7fHG,D)4DMgGDQK1L<^QA\dL:Ec7e54<UICN\B>
X5,XD4-Z5_?]CXgV(_8OaFW#a0DgSgfOb)I0;>V&3WJf<Z7ga.AF6&#;S#)?O<LL
.;?#fIKe4JSCX(gg-B8^<a39?TfM6UfJ^W4<515ZK5aSV]:Tg5\[FSe-ZW87669P
:>Mb@]c2\?dUI?R-,M:N1()K1KF/;^0SEZ2]7Fd;^HO?MA/_<WHTgX9U6]b;DU1=
&X,\:YHN(.XRR>4SEbA3J00\dFF/b\Sf,I4g7GdDWf+FYLV27[M?6C5CeFe8-D29
YW895P/SCb0YP.+PUOVTa.^Qe_U4?VEUc2[5SU=>.#L^YVf=J3)_C_JW[+.MU,5<
+1:;?D3(\X<OL6@We4>Ta6?f;466a<3,]baV_5^P-BfP.((9IN+[O9_11Dc]9?.B
3OP>O(+#[-N0[V.,:/].gG/,Je?YOVeKG_DC/<0GCVU(WK5C)(3/B=H9;XRY)c5[
59D+(U<:#@d_a,AU(KF5,eMZN^Y+G()5OK@ea>+VVN/5^U=b\GR3MEC9S(Z;GX?=
J]MVH\5?RM2H,UI;RM8@J@c1U3U\LV3,=N(5QDEE))QDI2UI?OA;Q-<5@:;cAG@_
R(b^T_Q7cVS^GW5B)YH880:QP3LQGPa&Ra);1JBFdG(HO4e]R/BX[V[e7BFM0(C?
D41D],Od\9FF-JL6WAT^D+L97/2/Td6)+CEIg@B9ZXdOZNY:XC(&bZ:YcR&P]@](
cFK^\7ZH4O:X16@ED#Ff(SN?2VL6KKTMGf<O>G\RTP(+Qeg^IM7]4C&WA47AIEIa
BgA5d/Fe[e3ICYgf10#SKBH7,F3[+.E@+\g;J&aI7V#g>g^3]F3e[@d+)d:M)8#&
,=B5C\^\^@g,d5L6JagK1Lb+UU+f/.?0@T+6_ZV(91(/&S86Ce_8gXY5<f8PcJG>
+gGMb,aD,NGII8K[-_bVN9]BD>Y5eI:80#]U61SZ-Z/FQ8WZM,#_A=)M<;8MA2.9
F74Y=;de-])/MdE=HXI@RR&6eZ.=I+AY6GP1]C#P-][N:b\JLMDfSN[)Z\8HOH:E
-b880V9(2H8<4a]R,c862KKf+@.#gJ;g7D0D=(-5&Ybb2EBF;QEOcdE8K#9Ba&RP
3URC@522(-PdS8VE5@\+)]N0P3J+dLFQ\RLPP&2.=>9+2fc+K6Y,Q_)Pb357WVBO
bE=B_fcN=Q+d;(792WF2;N<C?\\?O7dJBg/b(<=f.+T79<;:?32(7MF8TAT;Ga>]
7-:,NOHS@H&+Ob:[&X\=6YQfg6B26:QCXINYESb4CB\gX5KQF.60K^^:I+gGf48:
5Y]JGF[bI;-?0V1+U2>(TH<AcJ.-6[)707[3ZA&@]R]&YTH_1G_-]fP(BOX;30B6
UZFeCeC^fZMR/NO#FK@GWR1W8Tc]e<ba@I/O.O+3K,5>_LUVgbWB;=(?GO@60c/G
A(ZYBd;B:;XRZ&I/1KNHRKSI3bC\+XKLBZ47=EcU=WV?a[4;:c6bUdRQM<d:O-\H
X:R1QIFEH_e9<IH,b.0P]&0.S;#)?2B#N2e+Q&5(:&;/a,VK^a,ef&SB?C<3dTf<
J\#->XHD_))NPeBP(XX;JV#Q3<c]9BH#.34T(17V5YK:a+8d60JJOC)XW6:HQ626
)&_8G5SQD0=)\PEC3AFU()N-a.ON0F&N,&&P:3CKMgdaNVcI/0<.>TRXcRG5C5PG
4\:UN.TgQdH,Zd,cM94;Bec#\,9FL4+JU]<\O[J7BB\:;B+d3?2:[0N=SQ\GGP?=
&3WcW[-bc[2VO0B=RZJ2(((Fa3Y=CSO176O@DIe,g3CcGYGXg+^J,]XZOVL1;)6e
)C6KJZ-:@7W0.P7D(4D/a4V+8G(d<=Lb=[aI/b^6\@?(BcX.BDU#-3?25\OKG>]M
@aOd5VQe)\UZEF\3]J;N;OB]OD-/VZ87>N=Z=M,QUcI6J@d#./(2c/2gf&H24O]X
HSC7_6<(N-,EMTb^E)C67_eL^A^M#X?Me3cB[bOZBd+NKT=&N=G4[4g64C2LV2f]
>8;9,@A#b1+G<d)&6^5RG,cTFHOeP8]\?TO#BRMBQ3V5D5QIf7:^2=[S]TTWU=I_
Z/:8DW>35#e3eGQ4H(=#]SG\W)Y,.4[FVPL.@FXE[X\f(T,Xg)52Z_CE]/])faTg
QXb\[RW.#e>:IZfXXZK<A?.A[D@<@<&F#Z+(59(+E4YV#OcTH(]ZB4D[ZM+=\HUY
K29L?CEAP:K57#MHI^8?[<50&&KK\@Z^N\;)3(]/WbacSdECVagXY2^:5)XXFZf8
cNHYBaR_3>^W2)#JMNG6=d4W].)<D=^-d)I70>RY-#55G?-#c9;@69KC21-956#a
O29BU]QL._5cg(W[=+WYS?4H=/RC#L=AY\]ab?6(FP590XL7DH0.@;1AK3ZffFX?
85.V/,T&X.A<.aIP8F:,[&[P#&IRS76Q6<XH3?#b3VQ0#Wc-ae+LRA^1:PJe>RWC
@]P,Z7U)=gYdQbVES)R/B3Oc;XKFM,1/VG,VNFVO0@8#)SGFMIWZ)Zf(ee8@[Gg,
9[078aX9\bWR<FVO?&=?1EEQbNW0>d-dV]Q+TAc,R,0KV9L(,=1GBW_cPO+PQ6E>
=3N3\CVc/NNXVN)77A=6>a7(]#YU6^(S;_-N1)59UF5J9gN4TG8L8;GfXaON&Wb(
VB_3V[H37PAG4]EW]a?D]L5V1NR32DD5e,NdN7Yg:N^L+WW8G-4@A-)FgCL&H.6Z
81f(4[>1,E\\3ZTYA/^TbV-McX3eJX&)=f8G7=W]TG(adT4F#,eJc]Gc?X;ATBdO
agO)0=\M5dU_^_)XGQ)3A:B/=ZCYd@YSZ@BZ3NWA9PR71^WSJWNMXG;]N>B^1>a9
TQGgYa^CK6U2Xf5b3=SaBWO6H9/IFReHe(J9N>f\If?1P(X_0-b=\L(H=0Y=O1U:
=7PF8Q:(LKG44ZceD;+))1(\PU>W(Q.4_?TW8c+OWPU_GL8J-T.9b-[8>?H1/X@S
MNCICgST5e@a^@\P&TJ[^]D)1]Y8M;8+\a?_UNT6[JcaPL>OIVTOZNEIQNge-UGI
>P(D[#2TFePZ/5&-aDdK)d1E4\N#/\AIIc[M]]8<LUG0_J+1,-@Sg(Rb&3&L7VOa
MG#ANUO8?P5<J<&c8]&01M+9]0^P/.b)RJA#7.6NZFF:cG0PaK]SO.5-QX+BaUAI
/3=R-L_DW&A+<@gNZb)=?d2>gbB\)1_WeRPcNXXfI),bT]9_YH<CDf^+\#g-46?4
^E#:d4\\,If.[8HTfRccUU9UK.X.0N<L4Y#GTSd\b_NN=/]gA9KfLP)=J[A)H2,g
8ZSU]^@DCR@\9KHOV^XMG1:<8^HOf[5b7GYcCF\SB?3_-3\CF+&LeOdZb\d?E=FR
N\FRcd2DdE?A9]7/43f,N<4RcHVHFgTVY;@H#?HN-(RMfOc,SJ\?+KW,2=geHC.O
R<dY?c7=:6DH_?D>UMD^-bKe<\R(FRA\RH__KWX9^,JcbPV7QZQ5^F_3fIJ51SGP
6#eZ=2?V3+YM4a1T,S4<Z+_D^=:Z;BL\4Y//H[?CMObMb,95XfV^a)KVT3QDg#,/
0,gJ5)]=#eag\TFUB\SQ9K@[I?<@,F347O\aZ(<7dgCa>S]R^;gQ34R&5GaF:KN3
_9FUf(9Q8LY5+b[.VZX-2>#f/^[]Nc5O37/I\AP0Q3,D8:MC_K/Z.PUINXc2fP7Z
PBUL<1ZQA<KTHDdbM)M_PfP4T+A66E>G/J2WXVH>T7UD<]ca7.QZILW?EV@::6=#
;>:Gc8fS_P9UG+<^@Y9RG6XLN-KBf,9^\LP]gADQ4#8>a[^1:/;5SdIEY,E;Kb#0
EdbH1M^\cLY6GcE\0]LYDZ).,[W@feL;U3R27-7)B;JWSMLgJ+[,\(:F8/g<LdJM
]-AQc:[fGc#CN,->2MP;^&TF6eB8SYSIe6fd,GY2M<_^W4@Wd+[@Jf#b_X>BY[O9
Q3U.dWM6-<&XB?5AdE=Y<M3gV?0@]b>B)A^)]U1<;U=4DFIW78e&4X2cJBQ5cE-d
HaU2:Z8)3eQVJ7M>9L_2B/;@BT/&Q\eV]ffCEe29ES/1TC-6(IJ8LF/73Rc/O_+)
G4_DCgdVO8JP67fK,-fbE2e)RDa,3AN+46ZGW]\>3H<LdVc9Jb?;3\VJ-f7EETfR
62=^dHcHa.L:O+D7[0,@A8d]#1F]KedS+^XYNJ[F?:5?L#.2ORV^V<0\,#7T<ABB
UOPO/RZeFB(DCKRJA1>Yg/(MN9PI1e-Fa[_0N(J@H?.DC3f.M-3XUXadAA7<c]A>
YZ-B\A?//\5eE-^>?dYA>8[(+01aQMXH_^K=(LE5F3f&/b?VcSF^eTUP9g6,g?6,
bO27\G_(9)A9fN&UKa[/ZB2;Be=#[_0B=ObE[eY7<eS-NeIW_KOMMAEOXc?@>F.P
f,.83gZ@dQ)UH\=5<c160\O+&65F3<Q[:/BF3ZZ^M>;[LV9Te#+/DC;0c>1dCWW.
FD>8e<E+d1U?L[:g:5P]H-/e<11P/4SDg-H,>]b03U#P^@4cbG5_]^T2/4+:KWH1
Ce9H5#:(YB_]1/8d\=(<7fQ8b8Le(D34SDW#E=e3cI&Q9?.I&5\GZa/#1G3F>@T(
A<=6=.1a8LV/:6UF.HBGRKS,;dcD9EKJ=fD2[D]<[FaP_X@Af,(,MM\OO&e?4eY7
=\-Y2^8IKJ+=b1(WA:,I8D0f6W;@X\b;H:EB1gTU>/C6I9Ve2f)/R8QP[BZA]OUO
eF45(<-dZ:&VE.d/KX?&UMa>:V.\Zf50)8M8[@@MP@?([BP\,IFBKUBMe_5<8/[P
J>[\6cLCS=,,JGeFC[d\GL.0M6JLC)T6-N8LOM;]]La)SH[#A(7X/(?CYZ+D?[5;
7g/FScbc&K;.M4YaEcAd0LF5ZNJT-@XfE?&;Z\:.G]RY05_]1X;&5cA)#,_f^YAG
P>aYC0P:#>N5EE/4fe0&WL>56_\^=L@bC:1XIaVTgVR&IN\YA8/DNVE:=0/N_d_U
Zeg[ZOS9I2f1+YCO>)=O9B69@_\A@^&QQVd>5<P-#KeT-]]A+FY)\8_6I#O[0R8/
J)761&Ed6eJ[5&>8MEU)1R#H4Ef@)=785]@PRPR8F5@bPKPBC/OQ/7=I=N-#6U=T
#,J<;^1VN7UM^2Ad_XXC#,+[-;U;-YKD:8R=K\=[_RG[c,QD7-\5g_5?SMZDc</J
A.e?9H3?^(gUbNXP>HgS4C:P]7\_Jf/LF^:4XG3/gIOHO5_</;AA[+K+2KISGJ_L
3.(T2()I&NFa3<6^JE9V&1eL&48::E)_eM#9MQ.-Z-9EeGCa0a=7GEd?F<8N:bGV
>+f:+1-XU;>=N(/RCdL6@BKEcSUGf0=?^WBXSa<X<7PE+/?/&.#F(CE@K7SP4]@F
_V>=WJG&QfU+cd_3:OODST7?_DBG,F_<1U1SgO1?c14//g]R=&J4QJ,6(_.G;]<2
Od:2R-.bF[X5U:&UENPS#acB1+P-+E.<;?O&NM5;D9<W.O5<\ZSg@cVe6a7+MXc;
BW;\1]Q;+fJd#U7F.=1BVQIQOg_GT:MZG>+^&LGHH3M7-U#d,_J^26=39/QeXTYE
?X\IDK4P=DZI8:MT&8A9-,NA3&)MWe]+09I<c<FBE0e,98.DE>@;U_NRXB0&#.O#
9W]fL-,@DFcXN+T4]Nge.fe.]1^?>].#6\eAcI/YG;@;5AA>A5VV9N7g_._V,=+Y
WKR?9P\#:B=1:#GX-U2]^)P<EH&0FW:0[WU4IZ_<.eVECHOQc8f8=G5)#_CQ,._+
^<(.5N0=CaUeX,aTD0OR>FT3.-+5PPB,Xb??BSL5gb9&8ETedaG8N>;L.LC1459G
C&92QCLcO]cWP=9IBPU^-cPa)>D^:>[1934f)[/NTPCDM2;]2JE>a81Y15/P-?6D
S8#RS+RCX0IPZ4NX85>a.T(2+.>baLP\X<@K/S+U1?#J;MQAEe8.e+#@KV/J68+8
d(;]8c084E(f=>TW=(=d]bYfTdXA)DXI&VMK0a,DCBN7,=b(gL5-M6H_473KJ&^Q
1VFGFVT)92aF-,;<d]_L_I&CcH:=e:VQ3Zb@?b<HL)9XOZ9N]ETeY8S3U+T565?<
1BSV[D/E17]J#:F6MQE/;.5D^Vf<@-/TJ:GdP3dV-_83>I2<X2V2-^b(RS/CXU2-
@VObK/2^^NB-?c=S)NPBRFD0F6XgMICT&-A6aMV+g?Z<U4-WK]-O4FQ#XPU>^<XG
BH:1d&ZL+eCF<7.b.YL#dL[>6R71C-<MeJ<Lag_7e6,DEJ1:\+&>DN89-E0f[I=Y
0ZGA^5E5[fF6#IXMb3:&[DO]F^bJ6_VEDJKOL2Pc>LEN<DG9L:O0>NF4=XfNN&EP
(,fc0>D9G?H4Yc8IUFLUMF2Y:fOS4+/7g+:@/deBD+;aXS<:5\XKcWG55&Z+)YHD
\c>c6?R4WcIKOY90g<dQR.ZPB+NEP#)]F9/g6\^300f1H[a3AR(.#F/-)I/fV#F6
607Qb0GIQ<RCHI#L3Y#K,F<PIO1[gdB@IMYZGNZNS8&=L)c=K15SgK8W2,K9G)@d
DUR>Y7[4I@6>\NT@R4d92;a:S_RgWFG(bNE9?Pa2J<GNU,:17e0])\:M&-HC#NR9
)H6,JN[USST)WeX-YPY_&SW\I6\K8B]6<PAXb.CGUR?XBUgY>#P\;RQ=;2Z.XLHL
(0b>Qg@I8MY3CCc2C9.O(BI][ddB:c,9@a_9bORcH4D4LJRV7KELL_Q3\c#866V=
9=aUIV0VF6(UN:KcXFQ)&,B+@/DO)Y1c)])R<4,8GQFLd/g.K@PVM)e]B].W_FKZ
2M]bD^G9<//5LE>W.2ED@D(+6DF[GS3UDFggg=g^1/3d;/.U+OR+XbeUAF]-ZFf)
UQY9cXQZbgd:-UVUf5a.HX-+e=3=>@B1(TQLT+^D>J-SJ+.BN4,cf7F?RHHX30H<
^91d&+XS_H[:PT3B:^6/PYe>EX^:eJOZ:e@DFe)VK=5cO5]&S9.S/cXP]Ya;bOS^
7,].O28NL:4C-c<D;D#Q)SDZ8W4)Ud8]Q6Id<;1PP4+E6THP23-ZM4H-7-JEUE:;
LZDc0_P[^(TH=<777Ff\@J;Y<3=W@GGA@8(:J#BLNJ)<ZKZG,-2\_fe:\/dO]5DP
?XT.0_,KZLgZS7OVacH)<IKT2Sgd;Z\-^1eMc+51c8H=f(^2)]12BL5Z2\AW^RF_
L[Z&M1a7#9-?E032\3\1-,=(&ggYF#V(Z;DDQ_KQ]V,XXbH=_9:3BdU8N>PQ@[/[
PaTbWd1ZZ(F]@=efLW#dNB3@-cFA<#>F92TAef8SX?HCNW&Y5&g)H6Nfb-TcF]=d
HO0/IF7,^9P&K#ZR_>?)I2<OD)>+#9f>UH]J>]RSfUT1>95QaJ#:D>NW)3&@6H#^
#8B.#d_PW^OLcfVd<d=^acIE^B-Mc?0_.TC>e\1]4Y8(AeH?A\9:;7@O6XM4SVab
A;63?0F2)&WW(Bc.f9\g/6WdMR)C/:V>I<^M=2YS]gdN-41UVCQ>SAI:E)U)Y7W=
8eC]-ROY?\.)@0OQ0BK0H8QONX@E:CSge2[,[G03/8cBFH.S)ef)Z@dOUIgGe)De
<P:OP.KP3YE4K>,76D5@/(E(;7FaK:QR><##N#VB(2&?OOd_HDH&,HgbY,WBJVLE
E<Bf;0J<]bHPPFO.TXQfH0,G(/M-&.T;GeDU@MTA(ZH<G)G3B??,7F.WL1G3MB@C
7S=(-M8C:E/5d9Sg()XVM/.DE94N>JMD-cH0RQESb08)P=[=^cJ;XNG@#@<Q/P(3
Q^Qa_@X6:OCLL[,bC1O<Sc]J_2ZP<IIGYa1aS7E-H5^GI4fE8>6,2#XOKXE9#>;@
7Wd]7D(XZ&e5F1.c?KTZ;M\I5PU(QGf0Va6:NA=->3DA-V81V(4DJ[WX^>N2:5<M
H5+.EH)?+0_.f@Y>3/&I0b@\H1L&gXEIdJQA(61?8>ga-I[SK\EdC@]XN,?,NO_D
Kg0D9GW8T-.Y4ORC2ML,Q=8H:SW=b_OT21]+NF[<bOVcK1:-UJVcASH>[-&IXH]+
LgF\F0T&+D^(b0Z:Y.[.W?\:+1fOHcBQ6U@UFM,)8#\(Y5B@:<B>HcEU#Re?5?P/
]_/ScX6S7E6e@Q]f(?KV5\e1-]YLU49N9;_@<8,\B4bWXSWKgREY^bV-#&@=&BJ_
#&Hb7)@AW>SP8_OXMOXU<,c7]U+#c9UZ.g#@1>,][fd0L9>WXQ4YRb-,Z44R5;AI
5PRC#g&-;DC8>R2G.D=O5[^=M8:gLZb.3Q^^>Td3R.:.>BVIN7_:71@?\ZMP.f-B
MWDc=C25-+QGdbYBK)2-)[H7VJ>BQg+5E/9^8&^4E,1+2Ba(9.W09):YWZ,P^M7\
<a&C:QJ=P\,^PB7O>2Na+<f_UDI5H-UMU2.CVE8.bN@f:<;:gM(XbE8N\RO7TdF<
EC^;6GT73_Y9LcFAD]cf-c5c=:)3)<VE)C<F#9);I5Q^+ZGf;IY4O2BJ;FP=R=W6
NM&P<Ua?8:faFK5[<c<.L.;8-1B^,Mf;4O0HUUdV<9bP=GZ]Ue?IM74]W)0YcgaJ
(N6b^,=U@;I/E-#5IaBO@2gSKa3O)KX0d#U;(0fb;3STL/8K>QW1-J@eLU63QNQN
J>2A^TNBf6a0H4\MI9Z@:6L?Yb(G([NaIR[+(_E6HW2_83E4II0RP(@-1ZXTCMgT
FV[1;G&>D9>^a,6[:AT#QY33a<_VG9B-V+K6Z--X80Ce&W/1E_@KY65SGESL6+>b
6&PEV/a?.g;X64_][2Z&E1R4241AV?UJ>(cQ:33Na0[Gd72>Ug+-RWF./:UZ4WXX
<cR-9)\-_6EUHTM46APHd#,L]5g-;V]9XO^[ed=Pg&0@Nb6gUT\KA;.U,,((1S2+
O>[,DZgINJ3\6S^[S5/XEfcf&K<1d,D/?WE/0KM4P>eW57a\STI<>9gGOY?_M:_4
]\&(Z-6eR\73DdT?&\(D8dfBbX_N8\I_5[IYKEE.A#)aP1\IK]#M@bC6@;@MPCBB
U7)DKV9D.S6gQF-X<gQRcV\C)_:G>BA--,CJQ4]bdYe\.K0dDg591<PfX1ZB=O1Y
E,UC2I[MN,Xa<VbPf5T:+BNT^R?FJ(<HE85/>BBCSe0Q+->[fJR\FJeZL4d.W-/Y
O=^]\RM&YK]N5@&@6+6J6>cfNJID2CJFUZ>Mc9&ReI@FJP<VY)/H93VKTH_39EEd
.]<D\,S<dSDcZ3@:V;]R?6X78:&abP+Ib#b4=GB_a2UQGQ>562QH3=LeTE/6Q/NX
0N>d/VF&g5bRE>HZ_18L]c9R&dS5C49[>G4/9X@>6C0Xg=+LV+DX2EH/,)d,BG?4
SS(NP?AB&-XY<IEQ;+UH]4[1B:,caKQ6W@5FR9A37G.[BD=F+JaSYeXdJD<FFd^&
T6W[:GE2X)7FMaGBdAggQJ::f7NFUa5J+I1EXXGbHbY=XG>Y\R)fP>5Y<S>=UM:V
^X4G=GY#><cf)2V@\?2SW&DcI_ELa\X)gM82&@\[13(8F2.D<-gMBA/<B5a\?-(K
ZDSYSQBFHM4P8cI2M[>L\W03,dS2MaFRXW]#RA<;Xb)^.3L&2QKYX<-RXd0H/EO/
Y0N[+\)@FZ@6I?##;PHP(AQDBX6N5ff47=:_GfaQ5JD2#QSXHVNJAbP1abK<]9O.
24@33OK6cg_4eSKc=97]\3Z>@@T]Bdf0#Kf^-1Xe-A)\TDAWR=];^ZE?P]L0g+]P
<1JF35(5;0Tdg+Kc1?1&Wf5W=fe4(f?d2(P.QXIZW(,<YAI4(HGLQd=0;.B,-:;N
fD_[C(:[]IZ18P)1^;>ER0:6e(9D3C<+0KQN?RKFJ_DC\2XU,0CFQ&E9[d,,RJSJ
KQf&32-AGXJV&X0@aC4BL^F4[>43^W/Fe4XJ_NQP/NOI-1YcPH=1W5QR\,H3U>6/
L=IbK4PT3af5-,-g=L-H3HA6cYCZNP()I4Ub#VJ3]FX10Ked8\6fCc4>N@SZHKI[
2[7PB//FG8^:Y&RT;@9bUA(S0bGPL/5L_GS6B;M+bM20P^g8P9;G=;;I(<;)dbdN
+9cLHIAIB8NV=W?E1E)NLJ+DfLFWHMV7E4@B@7N.\3AP]SYFB>VfL@b#AE[3a[6,
cU.\BB:NC)R2+3_[a.=FV)@@463K1F@(4:(T?^)ZUNH6fc7<1#3E,bef@,(8RHMT
8>^G6dTdO_SMZ=?E/BYfeH_FbfT7(H9;A3OHc((M=AFZ^J,6[#B[LEb=KWB@\BGe
RRMJLOE(6&+KbP>PC)MEC-OgOe.)1VVG?Vb&>Rbad@f3L-T?,U,=Y@)P6a6.F#AC
R2&2Q.KDS?dc=e5#+AMG0\1(g(cEb+@IaKS)7Ua5TBG;Y_6;=//@20=S?<ED@H@/
a2G6;eC2O6bGe^+M6UO47P4AeU/YJGd=,SE#?2>I]^),57eXWe^-X,72U,):+Jb(
0CXYDM8@QE,R=:H2B6JA>Wf;eON&=-1cb7CdUV6<GIMf3W^/+S8M)ADXAPC/?N2<
C<EL<7,63d[F4EG8/9e]XW-7W_?L[,DDZUa?<MD.P<JD>B_Y@-K?S@Z#(0dcDOc.
a/+Rg0B0KIK+Tae6^dB]4E)?Y#?D\cfe?_Eb6?-:EYM:H_[@a5MbS4_Fe@S)3<[3
I_^E#RKTQ;ET/G8V#M8<Q:\cF:WCcMC@47a3Z]^3EBS\G;/@<1\\XZA3QaB.=ERZ
bc=^a@6#](<5fAYF@a-<R&H[bgGg]Ba)YA64Z4G?FVa9JbI>2=K).gM;5S;[A[2F
1aLd&OXW2eY)06=,=[ILD2N6Gc8aA@KITZBWL4JE;Z@12BBLQ&JIJZ[=NORca20E
1J&K;B,9(R#RJZd#Kd?]1(NYQ8,3IV\5O8F]ZL&[_/dR2^dfeIPH2K6EGG-\(Me8
9::&ZQR2++Dd.#Q9++b5ZeDLN,4RRSd62Bf^@=(A)0+]dRA-O6M+G164>HS1a>;O
-08IG-Z01<\\^4^U9_E\B-))@Q9.F=F/6?5<8]L51S,=d+7/b?K6LQP4\dFAU.&9
:eGH3b]>Z1BfaJ1.PXd>;2c5>gJM]2O20Md<&K>:L2&b-8/^,>gB1CKN]]CD+MCM
f1+M=@@((<Ab#Pb]MT+eg0MC]?8=&_:<)[^_R[[&5cS\C)eVdBgOc;4CfT4K)>E)
7H\UWS<cbef+3;8TgXE(GP(]366035)BJ281Z#TG#PDQ@W=QYFgZ4#,eUP@#B(<Q
#>S6/1ME1P2Dd2f9M7g?H9e@Y^D8fKeBZcS]&fK6_^IWc4>TBKT(:R6QR3U5]<UV
\FURS]XJSS5#V5U#0W.b1X6N&/&dLZWMaF-e3La?S_;UW+_/8Xg]7K:\>([LQ0^J
E7NU,X7JO<PDddET3Qa5[FI;=M#)&,:=1DK,;AIN?EZ3=7X4PcA@T_/XY>bbIcXX
+L6JbJV+H;2KW<RBHOI,2EA<[;\5M2]E291dfH2S3c4+]:VVcY;;@aAM.V4#-D+H
d?^BXF><1-_WMRA1DB.#M@LG4CVEP(]HAB]QV?8Y2(^Q_H80\W[H2GGd6I=;+\XE
eaYC]GEe:O:45[WgEKU+[1MHL_U<H_LI)cU:P;8[7c1SFb4@95Mc,Lc2.gG0[I[8
\56aTMY@LO_0OI;+cVIJ((;Q.<dU7S8Oa<;a.BBV(fG[N:bY-eGQ(OWAQ]SV0//5
,GY<38;I@7]]X\-A>]8FLYVgT+]@>5],MJ)A7,Hg)&Se9Qg(3QF1/:Z0,?7D0<c-
=R3aGPD[g69ORT3^PgJW^#^/7\(Y3b;KH6GEa>T<>]7J?;d6[g0>KGTdWX#Ge6RH
KOX^fC=M93&SJ5d4?[@+(VQ>Ye?:GA\&[27a4.S2I/93T)_L6;YP/.5,+B8J.&3c
DQQIT/]+_[>RKWW3eY@_]FYO.R_P02#:3Ka;X+I1IC]L.9G8V/]b?XOV>OH6dC+X
3@JTDT6OK,E>KNJ5dNELX]6?-@)9-V.YR5VA82JD_a+8^PDV\a6W._:3##.8^>MB
W;NR)Q2(GF&gf03/DW1W=/(U1K]IGe]N\5\5T?/YVR_JMaTMWAGQ:D=DQ]5&T)1E
SA&dZVA/W2C4?P8-57A1?L>@Y6#dC@.L(D,]:Mf17cbME&[M^[S=5&UaHU#3UFWa
[,d2=TE+Kd4GL+L.USBZA;&3Eg8:>8SDODODLR7/F@DEeM0Q2CW?V((F:0egA)\Y
9@34M.aFSQR[^IKH]6@U6__T4bS)f1SM4bZ7c-?=ObcL(HH=1[CI5+dP+#I./;?]
>C7Q.P18NN#f,FT:XGP;^#\>W]g,>+Fc\)1e--7_,WEK+YJ@(GKdF/-fZ+,G36@&
b@J8S:@_/P)Ub[1_=Q7^Vg;].a&71#I>IAOQ:L1)6V4;-4CYL1L.#K(B?6g9BL&@
F[8>D_SO&03fD[=\Add?[Y3LB,^^?_+R>Kd(O[d&HD(BfYQc,#<UD=9GVO&@ECe4
&M[Q_EE:L_8=/^,SWAf_?(NM@\/G9HM^#KF0+fQ80;:A?RaTN&;<8)S.FB;/>PR<
H=Wg[+7B.\7g-V->U5bOU6KU0S1,OM4UDaQP8+JC9X@(,[^Tb;(eL3Oc]]O5]VKF
g]Pa]Cd5#Vfe>(LUF9Q,Q0Q)]>>gK,UUUE2V.g@1@M>?3BQ-eJd]Bb8R_:BDC]&2
J,Y.YWSV\QJ2YTa:DY0YXD>/?GP8?&:__/N_/_S/OLJ9AQK5APG0,,XRF,;<Nb&4
HdNaT=1<LZPHeEF54Q>L>Q:B.H;=_XUcSJD9;D1&[[g5ffG0,S4fM&0V9dM_H@&c
RM(RJe=&(GMU>#&/L/VV#A[L-(D;S\M+EX/+a8N5X3/DK#=M.6YFV/BFXEEa]G)Q
D8-&3&b:P1I=_0B:AD?FGIH?10-^R&-1S[GQA=NI\VB4[BA)7<^7Xb4X36^XTD5[
TF(6.b918TP>>JQ#N]V7,^ebJ34E)\235fTQWR3M8)CL#K0?F9IDWf((W3D_GO>+
e#OD.N.4Q_7H8OM;f1V8b/(Z@S>IOP@f&5R;BB<H^D@?QUWL9>AQ2]+JIYYELfNa
H#AcW-b6VPa(+;O_.GIGK9S(O[UI0ZKW@<IEG3g9Q<3Meg0&@WAA5?6PSE[#G9EJ
<TI;4bR#+&H_WT1ed_.0eVB^8.^?Y?^eb8g[WdH@<Mc8WcDa-#OKb9#c/;57^2a8
6J6VN^U&D-<0Jg[#KML:e5&C7=X;fJ@]e8IR7R?\4EO4<FP]I#XC#)0Z>YPQ&86Z
EX0Ra^7^KHP\K8g)VdKNdAfZD9W,D2ce4E[86S9#fQ)eKf::\>gCH])^^7KB81Qd
IUVQe5T&F?)C+(XJ2B,I6^WYTR++J-2_eK84?eKY#B8IOL(.eB3AZN[VEB31eVI@
db9fQOfBG[L]FU7J759Q6)Z0C71M.+V(YUPT_4]SaH]Y&d1#cTgZ=TJb802VPW82
aTH&,bU1:ANaa_CgBCX16c#1aaB3K2S@g:8_eB>eRF3>,2Xe43J;/N/<NcV.>V>K
;gVZXVSO9f1c]c^A6&>:Xd.f_JG=>-.)DJT(gP6GEHRDO2?+3,ASWR,a0>0V#+cd
<_\VLa?E+-fRg4H#2dJ[E+2:_L.IXVTU^]RO\)MfgO1^)QKQA,e.QP>E_)4[.X/9
64S@<L/8/B^?NIZ<c:c],<B)YUd3[VCX[(@-X8RgNMO++]A2:V]#R[?T2&Z)U?f]
d)#V;OgE]bK/<6X.WL3#;2?IP77)LR6JLMJ6a[A-@;LQ_Dd>O3VcLU4H9,BM^6U#
ZeK.9.Y8G:L(EM@U&Y^cO.?7UXV#g:P)N_QKQ/aIeSTFb\CNS-;)X,?E):RP0ZS8
>I-_4-8c1E-Z:NSce]M,ePU96+/;U,@K3(QfO]JUQXg6AT.<BMB)NEI>)L-&J[E\
2-[R6_[M>0RAe<_&C5H8,EQ+DS?C6Pae7d_\<AQMbVgUWIV[@#7&G4IA+/T>MC?J
1FC3B;UYDIUScEW(B-H8;..DP-efUca>P@G0Nd1/b83Ig[Ef5GWPHR(CGA/&#RV.
6I^=#S43_JUXN=\Pb1F0f0Gg9CgWKLBQ+a))d@>MHg#S6e]MT,:GV2/,aIS]HCMg
db]I[VW<.DQ\2]F,<^+J9V1e6I[3#VR/>F[g5\NV][N0-4Ug(DE-I-W-6P\BAdH>
;XI2,T1)TG:JOD;e@S(S(ZY9_Mb3f92)6=^]_\.?.,>gQD0_5E(<?@84dcdbOOSM
2EDSfN\O5@2E3b&I]60^85B,ZS4bA3\Fb-^c?7)AUf^HTEgSX\a#.^T8dXfO#URZ
-3:dBd.VN>-7&1#eQ7ROOeVLa:UPR[6UI;=1ea2R.9]47?]19#3bUFDeQf>AbK[W
fBXT)SGX)eH&E,#(:KQ_JJLT(@fS9#08FFf6C1/I6bXB[b3U9ERZA,FGOG7&>V6U
][915BcMbOTJI&3CQ,JKD:F:-?aY/0\a6Sc=[P#]Xcc/3]:[&95;&cdI0LOg]4/K
WQ6I4\/0G)+_dg>c\=YCDM[SaYOa_3D?TcD[0AB,J,cYY&P:B#J7B,7\^5G6aKcX
(I#,N)e=VO@1Z\8VbRI,dUCLb0B_AQ7(cYBJEA;I]/6/+-,c+79ZQ:AW@]0B?+0#
T];a[>9MO3R3TG.HSf.9^P+8-]T4&QaGP+69E1H@?A9Q)N,c_VT#)MLF9KJ0Q272
X([RPdCNY#gB4Ffb7ENg=eK9>-\H/aXcH:1A?)1I@PR/?Y[d:A^@b3G\229A2G;a
Rd2@JB-)&,aeHDG+RK+8:[cg2G_KBV3CV#1/+DJ-8PLLBO?8fMX9Q\S&RZ(37YK?
c1H@3=:J[WH@WOSZ:fE2CJ9A+5CaX@8IcM&_-6E<1=M0IDUIc^\@.IB4).JNC\Ga
G=CHdB6J2YZF&0UU[+(M(6+RBJV-F\^X5MXAQ&JgFA/_e23Zb8[5-]HNLI;bT+;S
ZHQ:SH5YU8/e6I5].AaeTB?2&EcIW:XC/JdKAbYO8(bFg9TA;];4EH;,8GEeXHA3
J8/LG;N3Fg:1B07bD]1WWCZc5K4QVPWH06>1c]/6[0(WMJ+=_.@S;A+D<K2-;R7@
SR<H3d+]S[aa&2Z.c_WH5(f-()N4Q?g.JB;WAR:Na.A\BdeU10?a:8eW@&KfAf&^
8((D)^7#AdF-6VU:c13200VH5f1f@[Y3BeV75([NO(adHDJ8^PNX:3<HX7<+/&I5
7LTS@O#Z9W-@PZgA+IF2K.QSE<]fe?30E/-]SfD+T[;>]HJUUGA_.aUJa#Z3W.gd
IWPA2VP.f4CFF)8[FB+f/aZc+]CJIP4@^-D[T8YaOCUYQ&L)MHRcMR1e9d(,X0e#
R2?UNIE8LA8]S&2HU;KK.7==)Fb/-fZcACR4>c(4I\2O?3Cg4ef;(?Z(+bJ_FJ>C
MVZ;)0eCPaRbZ])T0^O3F,O)3V#9>PD?^JGNBB7(f9>1=5eV58C&.aa]BfZ@+D/^
4#9;-bN?b<>D^GdRdHHXZc]VH@eT8?RJ5@9b7]O^[FB7IFX^6(N92cK/ANSYc+_g
\d(Qgga>G0c:1Q:Z(TS_CXO]EW5]8Ke(;-E/S8GA<\8\FaP7?#-)_&0M[YB3T@<U
d/#E?-3]VWMIT9Ea)??.3>)[\Sg>Za\Sb]O19V]Y]KJ/LW+S&dM;764(Y+6&.gT0
5/GL_I-M[6&<7Tg@#/QMFQ/=IMcEM_&X?M5AWeXTWN@R7@(&9205A=29/_CX,bQO
YbPa_YT9I2G,+C9.8f:g&BUWW(+4^0,eMB#U/\Q4A8+@.EOHTWWZE.C^553EK0T8
+S05\YPHWH?TV@IL;-20CP-/HS.A<5N5]-#]f.@E<CBP&1FDF.;_LT8(7NZYM@LD
:9089@50(;CM?B\:B,WV.D./K0][/E;-OLe_^Zd4OX#\UU-7GcC6\/G9eECHd<bA
I4KXDK3.Mf5]HN8b>GdE+2(5P#5I0d_XE.0=N&W794\<1N;\7:c9(>WXPcN6J/<(
3<a+4K??d6(8N>?OKVgL\C0MgP2NgICT=#O:BZ&&4.FCfY6L?VED.,T990,(NRaU
8(P<UKe?X+2b1La(4?.g>d2/SS[9>5,SV_aV?:B&)4B[,Q4d3SE&A6OJZ&:e7>3-
gL@R(DI9?_3N+QGM?@4\>:O>-U:]3=)FVXS.X0OCHN^QXbT^4D@<HF8fg1/_YQ)<
_D=INGIO6X&Fg>Y-UPDO>7Qd])\Y[\^HcU_&B5AG?VcbQL-^@0<,g3&,c/ZMa-<#
b-L,1NBE1K#/M5^REfU48G+VQ3NaC8VIK+[]/@VP0.NCJ8OCVT8SQf-N,V;aJc[_
O4;.J(-3C]SCBcUJ4FH=X#LBML-MW;WPPW8?E>Q15Z0U(^3Xe)gLdU4eOega4e]>
YF5RSHa<=1bM2QLIB034(F(:#?RgA^T=DXN1<5&XEN^0K&(TcS5>6_=LUZ,OQ./d
E;0/cR1E-S+;]+0:_ffGN/_50f2==RL?)VG^E^X#_D8=UH9@NFc&K:&1[M_]b/YG
-8TK5A2.0I1fL5BA-7[_JR)d4<#NGA+5N+#\CGA7:,;B>Sd3@Lc]<W(YL/A/UQ^I
NG_Y.EfW9HSX@G/.A4]D>.1EUP.NfXc-R8UEC2TMIT(<4<PJgYN:X6-6Y-Zb/-)A
:CQQ#2:CUH&\#LS-)1KN8PX#;e;gOb_d#U3M+QE53P/G?W9:+^U@/OGJ^YB3f:XD
MLDG@[eH]495RD;+UTI1_A6E5[.D;Sa]6DNT59:<O=4D5V:])0K9[L2dZ.I9c-@=
^V#N3/\8UKOKfW<H9H[9LV?TeQ(ODQ=dC3dd20aL#\d;=eY;&E5QTA@CSQBSE_af
fHY06ZP,O5.Q?]439F90^-LNcX3]M\,_.V(N3>=UXPYZ^4e9_#H_DR=^9HA=Q/UL
CT6ACJR;2T)VK,=@64c\A7YT&XdgJ;EM;Z:<QW4gfcFKNG>5bTM6dR?6R@O)X0LV
XW&/dEb;JNQ9-#2F^15>,_S[.(0e#,TZ_+,BL&L/>W[OBTGB>PZY:G)VIbBKC=ZB
[eT?J:2DWSS=a/Y0JcHd?^O;0OCDZB5D8e)Cg1_2MUV6S-M002H1[V09WS<CWDHB
0a_/+.@8L2]dP#Q(:;UHUUFK2.;X\WDaAF=Nc0g/(gQ+M6BNYS+=IP):b^F_E;CN
7Xe9G.F22#e.5bHdL/?.0SQAT8S69;faG]e(eI,?YQeb:,,<,WVf]+;W0;HDXD#J
>=TSPC-3e@H>9C_3N-W.0J]:PRA]f26E><2NOVC+Z<SB+8EAUDT/O[&MN?3?R2V+
]FF;#><T:fYR[)=?FRTMQK27(FY4<dIRLc=J5;5ZFS/P6Ybb(,)N6R0K<dVgdd6c
M1cE2M@C)D9WJFTWDF91C3Q19:H2F/R;.f-\.\02Zf9ZL[2776HcYAFQ_00f6\GT
ZY^+B_a2,4^cc;^?3\6IY&LFaHYV;\-GA;8R1Q;eLbJ0:QdOZ[:2+^N#4ZF7A(K=
LedQX8ZA>#dJ2[L(Ed86&=@a1]?^df15+WDdW\[DK0d-7ZX8NUR6/V2:dQe&eU<g
9X]d7L;4=^&#4I14.A6UH1+MRaHP#WRdNd?,9CP_#RQX&g;35+NCOLQYM?/GTBg+
1b.cbH[2^@YT?Fc(Z/?DZ96S/dZ@)&/4=G)->-=AcSY<Ve3R1]4P;\/e.;3)7C\Q
f/93e4U2aY0TRL&a;7F+Q=0d???>C9\XMQRWTKPO:_<?7f5VcB;Wd[b86U#1Z_0.
g/]4EV)6CB9+)e1dU5Ygdff&MB23eb,T?gY@+@BE&7&#]E__A]/5QBVZX5.8dV\]
MP;@OMI@Wc6OOB7Ze=W8fH49RbcUDM:BM\+EC4=/NMZ_>58Zcc-[6NU6YaRUCDaW
J7,<.d=DN6F,51(V.@=GN.XU/&[/^K=&7eZ/fb_IG\0MXLb4,[O2dZVcfMGSH5P+
#@GB.V(]N3TVQYB8)<KdO-a&2&0fR8FMPEJLJCM<@MNQHO]3aQ[ZPFd9,^55,/fR
<C]>Wa#Pb&84YOD]V2D]Wc(+Q>UM[T-+F#LQ4(8__<6Q0QH\]b61X?67.AB<TFP<
KD6Y4\CR?/(U#d+X06N>[c2ded3U,U(?;O_9d1/)\A?#@UaE7MO_A:M>@6:+]+Jb
@(O:[C?]3,+DN3@>=G-6[&=9b4BA=YAde,7R9LAIBXKEKUd+@]PZEQ\Bf>[fQPWE
G#P0Z56_:0eHNEbc#IW0>(6<R8bJWbP5AAcL:QYYQ7G.2Q-?<X[1fCf5ORcVL-1e
c):TT,P^)e^:X_3TaH28=A&Z@aVJ(C]]JYWb1A;PQDbU=-bS&SDN/N,GO5^c-:fB
XKJ,1Sb=bCe?Y2deJb9F2P</4F<NID_NF&b7AD&cUb1VM(9L@?MeL9bFVX^Qce67
MCK8AF?.dFQ?\A?N_Q_9(AL,+)cNJ@H@4e=@ZG6_+<J:<Kf^gRagYV\Pe[]-LSaY
U4M,AB,<eQ1&B)QGDc:Z=>J\I/J&F_KAAS1E]Sg>&^.K3S;=dKK][(>TC]9cM_@P
C?XC1dM^#D[7/JYW]S],G&A>7:?F;[eOK8,\\#;^PQ\J&&NKBY/aS=__FDRIf]\<
NX5<BD+G5?U2FX#MIM;N3a9^SKP5LB9S+P;?J9gV&3-Y@I<Qd.DM_g?NLD)9#4X:
Dg,JC.51PIgW-7Kb8@fb#=.IRD>NfV+)>0##<]g8LHTRR<.3.Q3=N;(Sdbda]045
J0+ZR)+/QEN>-0e^2K5bg2GIH?ded6VQ8+-T[/K?NX#H)8IAO(;cJELUa6d6[aM_
)+?D5S)0P^gQ(PR,?d<XY[G,:BRWaS.UX,/IUgE3g?T6GNW\?f2\GZIGV1_:RL49
_1ef2;#Had/8YP(T#Y4?XH^/FCW?/U8:WeXZ9Qd>edJ<-b099?,BX1dW0/7)H>2X
4[4G]J/JBW9C/-I<ITA#&[A+90f@cOE.0Y/VVG0gQ.ZWQ31A[CIA[;B-Z[KU\/=7
.+6aDA+W),XU#M9RBOd#TW4_/&UCUE/#cOcO9?2Q,R:S?,d3?QRTWBV_>DW/R4a1
TW:>bO.a+4Mc5Z3A(aWgL)(9O(_D7XM(F0=bENPe:EKCGW780&#<H9]]X&.ZCZ@S
C/QcQgSWT;V0(?_AM,c0<Wd5c^M[LAC\;7XWF8BK(3@Be:8FWA]U(\bb6[ca[9AR
60(@.aZBI&cO9,F[KRH8.(:#-MXDYHVH//&?KVICg,SEI.:3H1d?LB+O31]O>TC,
/@UF1)gDHB-NJHf]3:1/XGgUU=;W8OBVH,#bJNCBK[O^XJcg+C#bU]:F,&W#]+Z8
.;d.:EXN,26\6IF_-854:AKQ0W:FQAT-COZ;99=+3I;a/)&6G/)-_6cJ>DN/RSb]
3(E<Z;faX;_278AZKEK+<1,6#33K4^H-2-)#9<+Y^O;^>-4f36OG1[I]J<RfKfZ.
Zb,FWSN[R12EPF7+CM1&\A04M0f_C=3,#+N1L.3T34N8E[gG3bS)cV>.>NZ:-7YC
fCLa,,Q&LSVSH#\(AW8Pf,KEN013Z6)HG/(<2WcbffbD,<3OeB@(0)H?/7#[I3]a
A^4CC:Q&)C+L4<V:(fYFFWVT_+dO7Q36gX92Bd?>.KgI=1K&c4XJd2GVJ\9b(TL4
VLTbF>4cQf99KQQ([e\Z_O;@T.01T7\<Nd:AYON>C)48D2cM,)Ya]HTFVMW2^TI&
b5/UTOV,Id.E\D<c7UTO:c>0/TOfRFB)FD++_bP+9]:F;IQ46P:\f&>]cQFb=@FL
e##5-Mbdf-W<bXJTOZLRXD@cY^Q.@2V2F/?#<D[dLS/gL_.IW>+K(AUH\BD0c;9a
86WDG1-e.1=cA>;6<._T8(BRLcYf>.#I(A2]MR:8>a)&R_VN6>-6/[9WEZ(f4=)W
?NB#-dBAZQ/ZXGBcD].^,dS/2^a[_R3cYSSAF)3)cYMb@aM4KVS=#).(Y-fAeTW\
&[Zef>44TK)He)Vf-0Uf.1b04d03ZB4,8g3bV6_SQ[MXUc=45Z0\D@I:J?^BA2fS
C]]V20@D6>E>:G\IeMNZKU;E42F.fg>AK+PJcU#QHcMe)+Ba;>M:UQOPJ5QQ+W.0
K?/LV@<0PNOEDEg?9OP=Ca/Q.;OXHW@HS&1SNZUB6Qf0La\@HcdNI5#OIS7\d:Q:
XV.Y27)0G\#P]@f70[RHGVZ4Z.#9eKcVGZMMOd1V8,_Q\ZcIb8(;(-ef\<BN[I>&
)N5V+:CLB83?_<:3b\GGN@c@WXZ5.)>PSfS#a&cX<>@YHL<N@77OTb\4=e&7M<GQ
UK@/1[>>V5D(b-J1>T5fK(#/_P9b88LHYRVG.[?AC+EV,MDC/YaGA/DLP,:SENSY
AR><NN:gd5f;>F3f<,^Z\b\eg&K8O+\BKFWFE^YZPc^A;f1?KLS)END)@/#g0OF+
:MTNeJ^_MGgJD)]W/-(),GQB8&LJXOP/+WQ0LZe3FPNg/^).Q0O(49&(IZH@M+G:
a^^XQ\PQ.->CX]?TWH2dbJgH/^2U^1P+&0E5<U=RF1OH\QHC)G;+57@:I4R&N,2a
X)68LGUPIH5T13[]23WcYJ0f@DO]2:\f/>e[P4E>#>g=T&H3.gIC4KNS\@#IS>;,
<J(((g58AKWU5c#?4AFPCD1Eda&e(H2M]7_H?[^O=W;d8e#,RbM\Gc-DgD/H.7,;
:]/-;.96T_WBbC3K+DLRf5c1V>7LB_HJV=ff?gOKWOZK@=N/LNH9HN4=CM8#a5Db
2/W&Qg,ECX^-P6/YAf5Y]WK;5cdHb)^<Oa&(C/ebT0ZV=9Z+=cE><PfA:BP[b1K<
EI/#G2=DA.E)V:UI>0FJ(33@;N<F,5FWfcQ=H_f__ND>2_.15]cf:RANLML9D;RX
I2+fB,:6^5:;c.E,[g>7NEgL9V6W3c=3_5WO.SF<(QA:eK<Rg;R7S16N;?1#=Q5N
FG=2)D^I32KGR]X>Z>H;=TR;^c<:KKce[XeOZJI@c8daS#<1JRHIGK>3;Cc6->Q<
L6IgLW/b6AA<(Q3T>W7;S/FbN</NVV(U]2;Re/]O9\(0,=YV501.8=U?JA5PbJ\g
IMKK._4?4Af<+D&9+<bJ:B3Z@DQ<+\gW4fTg]R^g3F+KWa>9WVAb9/geC9YR.XGg
2^34ACb:2FB-Y=G9?@UR\71:#H..D6KD0P&)e-HRO+EH#4-Xd0STYO+e/:b8@.S-
GYOU++a]5\a:75(N>ggIP:-)c/cYFV>D1A\Z]g.(T@\&GR8;<9W88]1_4FK1=EJ\
PI6;S..c[##:B7@PJ[;[;1#_N\G8/=Q75IKSZVN1?P^^H+]&^.KGFRd8(W^8&C\H
1T,0[BGDI43@3MVKX?LNQW74FYDPQ:^GXAf.gc48UgPbQM3-(T3A4HG/=(&&^5\I
c/=e:f?O,1,]C<_OE@WE92DJTcIg0Z4ZB#Q2daa),&QTZa9^1gS5O:NG:]K\#N,I
DeNQBYdI_/4MK-[=MbRJaYaBXKJ50T.UC;4K.-#e]g:WML&UX2H4beg.7THD8[5+
.K0L^C2<NN@>280/\SN]-=@13)g-+5Z,__(1_e#R(^1A3PCKgD^ENf\S_=5KeF.-
-P9PC#AO0M^EY3.GW=cZ:d<&QL#Sc@0BAgg2S,6K?G32V;QY6HXHAJRPGa?e+HW+
J6c7XU^I#bee6M7[X7-=4c,KCYc[cM=&@Qg=:Xf\8>7]XdbZO>MS/NRW<:UaDcE-
#0B;g@0M9B2d7dJ+^3EBFf8eOLdD6PF0N+AQD7NBBQ+82MOH^Q9-DdOMc)gGW:9_
(5VW588d&dM9KeL50URa^H&@We^=gRgKgNX33ZT.\TD=J1&/>D.B(>([]\dgVbd/
P?>aVCc0(XX6@ELHHU].G>)62]4H1=g150;21GN@J4LE\4:]M,bL4-S0A>[7<_<?
HR@bFc_W//_22^:FfA;3L6gU9[-#gT.5X9A_\Y^[QYgY-7ege6J&97<Jg7-:>DC\
WPf&QGPe075AN[eb,VB,V(F;<M85:N)>UPI#A);-a10HI=Z^^A.7UPdgEG4]ccQ2
EU9_KANELWce#VeSC<d+/)FfW\F87SB7?NI@HR([RV\M>f5UM6&K.4POEN:INc@0
aZ_7^S[.#PUg:8fRHW_aO7Qa=SbT6.8]MFf;cD&a/7+1E4T6+_&[M2KS[>ZNKLTY
Lc=1MT19JXR,,98;0R8;d1d+C6dQW]?4(MdUJ);BE]?#2cPHPT_R#RQ9DMZcU7^]
5C:-K5/a0L1-2^4dJL/I,T8=YRD::T(=:YU.;TMJdVPZV)H,c<V\ZM^cRKIc2U,G
2Z47BZZ>gdfMHW5V5N,^BNI6@5g;B8&X[W11V6a1H3a1?\:fS#87[=:6YK.0UZ/Q
N;J\H>J)I,OIZKKWRQ3f</^dgFC5;5E55fJBd&a:((TQFGGBAC\_VZf-bfE]ZE:#
,4Q[U;fQ49(1d[3N^Ye[LVE1LQYN,6CN?BZCW9;@E09=>4g.Q+#Z5K\=)f&8a3>J
H4?Z(?e4T5<._974ZYF=8e)WZ9QRU@Kc0((Yfa:\3NPX<M.X,JXX8L)EO<V#a]I8
PG0=MT35a9Yd&T@_;>.6/dY:[5A=X>B5#MN/9)7Y9[d#J6Id_NFOO^N(#-3BW7-K
=-AU^Y2_Y3A,[CWJKD15;P>1KZ:>DZ7_XHTSF/8KQK4552KT);H,UC4e6L/e;_E)
>Yg0I6QQW]W45?L->Z;#F<;28:LA-89U1,NGSCMFU6?D6HM=]TKYRML<I0@=@JYf
NMG&8XWaA/BV25PXLO;O[1#W;G;#dZ)3X7F]7UI156@-,HH+-Y5e(,^=@T<XU5HO
QT,ZG>2VG-J1V=O5<b(3bN;a<:]EUFIQ(K0BN,I./5/A9;11HMIdP<[eRZDBF9>G
/@b+K.G,Ob^+CQ42+_MF.(]VaUbDdc?EKOVPG+Y3T#+afPI4\NF(8GL[P7H]9.1g
NTU6F:eTY\L2K9b[NQ]W1E<@0d_[Qf0=035_b@SIc=2X4P06Off7.5@1B]&Gg]7K
HJ=e]7SPB4YG+=fIeYC=U_SZa+BF)EV::HAd[@-Ra-DA0L)b=e\:SO94^fGPa,;L
ec#,PgYN0IVE)][WeP_TZ^?_5]ZUK<e]?V)174&WR(JSPL4NSP?C-792#SA\>9UQ
?V\47Z/Sb1MIJO]CBB<UI9FN2TE>)AHB_3TGK@bW_=U#3L_=GN3@=E\1Q.RLK/BR
HMT1.<FH@J5c7E9W.(MEaV0D)c_B^#5EeIT0D<A>#?NbC\^.^18EFL]QE)fFUM8:
5D=/>-g&\0+;eYQ(:[(XXHT\/60(ZS[2.dVAMIAORCT+FL9,3c_-L)C87K[Y7Y8b
5+d4a=T]O)RW3(@_;;3(GS^>fP]N/]YJ9/)N+;PFESV-WE(8]#>HYIN[91g+.+W1
#QUc@b]I>bO_0fQ]EEBTRg#DRXE3,Fc3:#O9:AX3PYT34P,Y)?15D7a0.#1M1-Je
OBKBNN:LYS?Q\@.4YCc;SLBJ3#]^^Q?P^&<G-?#\D\\L2<\&S36WK97HC9?GaVL]
FEc,C_<>_O4Y]fE<Q(WSZf6+c]68C4&ZgdbV\XcOW8GU0FbY#;=<3.3W]](BZ671
IP@e;9S[/^e.b3#_f?f30;LUZcA\G&IK\\g>3?;f<W..^58X]:OYf#GgCF[X;^V^
aJgPb[JI3>WgbD5D.UAK-0Og1#?d<<H.Vg,S88<MU/2c1MDR1,FBaK(,AK>A7YX3
S+;QFPS]:0NW9:>C?798)/DMa_PT[A3/O>@Qe)J8A[=1?)Y5/JVR79XQ;TM6-L&6
U6576(FY==(;3.ZbJHf[X(H8FL3\b\(=.C>Pa]2XH<@:GA<G31?H<67F,844<7Ra
/M)g&;e9)V8fM/YMF5R0:eI5GIC_B>:JMATDIIb(J,XTQSE>=\>)c6R7I=7@\6E.
U1?B,Y;MSSKgO#J.Sa>BD_;GEe.[^RU/)@),(P:POb?:e1NdCf1Ac6VBT&>G@I(-
DGL9/(WPH-75@1BLV[P-.(4fAIXV]U,<)CDHRgV?L,d@Y+SO7c_/[93^K6G.C+=V
Ae[1I_Z_?=eeT.EG<.\:9;\6T77Ac5(D1ON-JH5I<UF^9V(-Y&BbM#&&D0B)M5Y,
0O#KD(IgT/Zd(N)JIcZ41I:WI?WS:4c6(7OHU8G3XRDAD..48ZW0).L5.^-@Z7GE
,Dc56G1ePIEU+Udf_=L)PX&g4KS2Y]Z&g6&ag4KAV\B=KP/(3WC3V4H?7_Y397_R
?;7QgGB&Ic#.IRK7dO&G<X,G\?PEgY1N,aMf:7.9_YdQ-e?&V-OSM+>;_8(D34A=
IXFSeAL;F(Yb]g#)\d>\8C6fZ1?T97Vc#Ba8+0P95KZYK#<=>HCPH=+a-c9](L00
8/I#,a)_6cC7^dgH;dJQQ>CF540.0+=L&7-d\]Ua2fLSS#dJC,KK#1Y]Bb<6e;/6
FF:6UBbTSP)P(TbB_><fZg8eg8SAYbZZ>DE/Y,GN,NA(3VO=VKX8#GM3CCZ,]3_X
MS=S+DLI#8&)(YT)4^8N83_FK,^8HG8C;KSS;;:_)4O_8>A6gAW5K)?YG:/^N0?8
JIV2a:1e5#\4c8geH)^X<3g.9,/@06I(&G#\V#7PLdNS]NW.N@-RJ420A4<SaA67
cQPb9>)?RM0KbQ9A3WXDeTIQ.O+.E=P\_6L5NB1d9;ZLd/>\J-VT42EB5C_(I/WC
E+7V&3/b:JW=\&a\OcA6&IA29b=-C_N.cONdbcg-OX98<7WD_[Yb]6&+9f/?e2K]
2gALBV?L,&#1@ge(XEWcMdA,d#\Qb1?=KJL,#J0C]<;K]S5b,OKGd<>M8W\56#a4
3=_.X?&Z]NTIC+]7EQGUATGOA^ZVQXUB8[YNV#)(L=IfT;FBIDZX86(I8F:9H;2c
d<g-@(P;VE9=C(@-U<O8WM[V2SG=J4K=)K.?4=<VYV9f1[cE:;CD@MM#JIS8CN6[
W^+]4_Y5\D87)R)49BF^QFGW\+A.9HT4+fC-MNG<g;8bgLF^+T+&YDeW#cVJ<B3)
K4/3=_:TZ7<P+5GdSAd3&JC<VS<]F50a>P-DS<fJ_.\&L/gL@8W347I?KUCG.(=J
-NMU3X2L\X=UV^fCYd@-HM8/5;P8L7e;fC7&<Rc:d8L.#gCeIHQ;MfFf+X>KXfc9
[Z7)K>d.HJaKg6f),8B>YG5)<[4VP[LaRW>P[0H1P381AdCNN<._GdTQc(-7X\/<
E:+^C3bf>]2(b:3g2SITga>]L@Y=A#I&YcB5N#7=NK+^2VH+<Se>3BMbCHg.]+_?
@e?+dLd69),H-<4:Vb^Z4N6:,d#bP-1AHMF3^W+Ebgd,38CJRgNe4b8Y3+F^a8^A
[;f4-&=381#\4d2^Y3HdQ1_U4<\XXVB\_CJ/,19&LIa,36<>N4.)a:],ZL:M<0PW
dJZ/;FI2eE]@<)J_XY?Df;\V+&+Ae<D4P(I64W>>#Sd4;.3\?.0NFCS\U&Y8H6_W
:,f<87;L9_DR5A0g+;0@3V&62@LQ<W<Ie2<Z)7T&CZT\1=&[88C3F#VS.g,GWMd_
=3D;VUY9J16^D^dN;E#=.3?^2)CAAN\b[RO.4.GX6Cc:4&8H7Q8?Ge\f_]C>[\Ad
B>+-O#++-#W_Q\3NT@F:9,27a\B62+=-/C()UH7.F?FSNDBf6Q^b-P>_CF5-@:/C
2@cHLJ9-U1bEO^)5J,9\]2P3@>dSa)@=^gce>W9C=d2@RRgJ;fNTVAdD6E)2U^>/
@Y9e[ORL<P5/^3LK/U4N?L?CNB30?/Ed;DM#<]BSBTKM254K3b^L:/e-?b7S0b39
(;JEQE/MO_9[JD,:61A<8@SeH>aV8>=L?M(1-@D50HB_F,IW@5MB,<9fBg^1T?4[
S5B=?Y#N5?-eRESY[f0_TV&#TKF]Oc/;Ud<4JQQT9J[&=^d1IR34N<<BH^S@&B-M
1T\:?e0))cc,d#AO/aFfeK2DWJZEE5^F]Fg4GQDTP5dAI8S6+U6FO<FZ_8@\).R4
?\YAYcYD<L6/,b?SdZ#Z2QK^e:OS;68b]CU](S6+d3cQ[.[:>ESYZ.&N9BTUEV0\
2I>D?&@OA)WM)T=,=0C=eM<0T#)VB8dg6@>?OZ9C98#U57;@0c#T/QSCD1KA@@/[
<<G)^C#\PL004;g9O@Y@ATb3Q9X]Z9.1d6@@F&3\V&Y+(<:N-?A,aa>?EZ0K3IC6
;WIfe-bILXTQ<>1;+-QV,bVJSN(K_739RMTX@EE]c?aVT8gB8(^a3E&G[JG+7E1.
#f&dM/aM@:gT)46D1,OF?gVFPKX@8+>@Qe6EB_UgNbSIA;.ZZ+W,Zb)+>OWb)H#9
NZ2+\2K(6E3cG[TPTI/geb_0P[Wc+P#F[38R02&_R_?YD(V[&Q@1<6Ic+\?-R7gP
KGAM\5R^@70RTU;PR3B,e#bN4D5g<F6WRBQOcC\P<0NWZ>g.WV&XED_&&DDS)gY:
VDVN82^07Y&8GT@0)ABX([-:,eKN04IKNgU5-60cC=,gNJ4]=KScLOUKKRH]H<ed
Z4Q/GAIG<.Z?B7&9-7?GXP:R0AF-XC#T[T\^(^0PBPS1YVW11GS;WV_M\;)5KP3#
I>PaA^C_D?DZ5:)6e#eI:TR-,260IOZ^??LN0NL]5b3F.b.e;AM)6G>eZb=DB@YR
<J2N[.@6#EUWRMUY6>DXA6W6\eGN.4V?G.V]Z?I?]E7c(5GT(E\@I_XRR7[@BZMa
:Z#:\N]T.0e)L.R\JUBRfL3>[fFc?OaE;Ab?@KGH7SFdA9UU-)cQHRG,E/>O__O.
L?U5(5T8Q;aMX5eG#:]MYPSWDT([R\U=AO[Qe+/AWHUG&cU<J^W8;;PcJ5Ud7-2a
g7S5.e#R8>9R3K43b<UTRT<\aTT7I][U[d;f1P3J;XVDA+P-]B7T,4(,4]+R4.-J
ETEcaDH5B3/7Q-/0:F[,VZeON+TFIPI?O+>CE\HQb1)&BD&5T(XLS28S?]E=<J?Y
3./dAdD?:1;U8DA.(Y#P5H+Z;<0<Yc&:19FWc#J2E7&#A.gDQ#g.5b,dISOS34d1
G3@0Af2=@dG\<b,<\2C8F5(;54?Q+(S+O9N2aSa-ARHgGEU([QT/,9Nd,B3_N&@B
:_:S4K&Qf:P8#YgP=T)P\WKD9,(L,M=b+50C&OB?-eYU/gNE:M.1\F?cWQfKHZA+
#9C_9V9;]?YD8bKVAKE?;[2W+:4]Q0=MBOb?0HXB)18X&=P[K@-&D13?M>1#K?27
,]VfUU[[WfGA6X9g]?J4(MMX=QdJ=>(-Q3f3bON,ONKBC6?XJ[((K0>1HdUB4V=P
)FeceT0JYI8^dT@RRI\F^XeL,NK67_H]/c:f14Cb.][CE(Q,[d0KO&RAeFO:O1J,
9:0VC+IQ\g=?Q4;_0K67e_HgBR3f3[(aVU9<dCA6)^@6YBSeRJOM^aF9(BI->)0]
DYX&Ief6RX(5T&951P:1YW]YUD/JP9=JSe?7LG>?@AUA#,2V:W7CFcX.g9BE9RR3
d?S2.b,COPISAeRZeVb7VM;QR>Fd(NDHW@M=3#C+M36PVI2e7cQ&LN<I1ZP8ZXY4
V+_,GFM1fdZXReb0.J6N+M/f<@?@@MX?e3A+Qc/FPFdD<@0F^QTQP-Q6P1ceKDLZ
Y:<g2ba<(2TaL&4K8BQ141K==X#,<(G0R@>=Rg18U5?>Ie3?H0GHSYd=PU37JB5-
dVJ;bB@^XgJWfF-<;Z23)X5R&QaQ^bHUTIgN=fZFSGe\=bfL-Bf,@YI_348#;XPd
c5M>\T8#EG)6<3>LK[e>8@2V;N5C<F+I=GKeca8-GC-12])L/gbP1C>[4eBS.21c
&V076XG:W+0\#DCGQWR.fY=@fB#G)a=2dKU3R7;D(3JG+13O5(BY<4;gE?0#.=;R
D@OOaf\<)481C0(OZ<+1Cc;eQ??K/4AOg_E6OFH=>:(M=\?K1Sg-a92Eg[R1KcHQ
G6c7J@PBa\VAbbRR,3J+OA>8CcI3^8[7Xa,]:>)W&KEg1PNNa#]]JI6K&O#+K6?<
URC^.;/:K1_/)6@^7\?(;a?61:ZS<GUN(_<Wa2KGB2@1CI<O&YfC3=&W\QIE2@f9
([M58I-PPZ)/+fQRe7N6LeV(V^2f>Hg\JZBZ>)VgQZP#;P^d243]2&,L#M^TEY&(
=20TMBZY;<[,Q?@_a=3J#YfL:I@=8G_>KW<Q]4(,dLfOG#^IKa=Y(&.@RDWGQ^gG
a<QCRR)JZ^Ug_dEQbV\)5<BbIB0-M>T(EVGBTEeI/<-U>O9b23(MVLOJ:]gRXATL
1>W?aV-I)&B(Q72?6DW6ZD(#f(GUJQIB[,8?OG]:S9VB-[0fgHc>A0Xe-?.cgc#B
Z:4S]dP:A)]BH0)-H]N]]N;7Cg9G8W<B#VKH3=EXD0feANYRga@=Z@/#;#VM+9^9
2f5Q@0d/MC_8V=/CQ&?c+;5,U)@[>./A^UU_YR9^<>GMe34MBS(3;BMeeUe:>F,b
B=T5#;d>=X[LCW>4,6\7,&.JI<b53Bg)4TI0c\6C:;&dVb4JJM_ZU4.MBJM6&B.^
V6I=^6RV/Y[-5N+34;d8eMIW1Sb,K/MbV:\FAF[G(MfR@8e]]0J-FS;XHD5-/9Q-
JEJ_/M649QAGWJA-^:OB&1_OC,.DR=8OFCcT])LYgX7aGQTVYWCCL;]6O<2C/2+-
<H(&d8?GLDO]II0;_eTNg#^V#Q&YSW:b0]Qg6gP0HJ#X?(<^.=L\ET^bf^G@LPbd
9:HaZAA-&eaEN<UQBNd?TH4#27Y);\F,Pd>^?CbV<6OV_TF8gYaFOWQOR8M7:#[]
bF2f;FTRId28\>&O_+<PHK.<E&T.;#)1^O\,ZS.A-RfSc1fL=^O_:;WM=Q=(cDA_
RTYb?0Nd+FB]M-&5]0:-ROQJNHSP>cJ=40++_)(KO,7c@9JgL79G52^)8Sd3NVSR
J?4QAGe\\cMB([LVWeG)&_&V?DQ@S8[?&T6NPA2;@c^e<;[K-:XLI(64[IL\fT\^
L&bg2T5.S)O+NbN9E@E8da0:NB/G#9dY2ZVDGf;gZb1?EH<Z4V(LOEZJB]>WU]:,
NaP2-ILC_JcJEe&a@GI3ZTg;6WSLa=^VUK#&/]be;\>R-5Rg[<5MLU3Za#8T7X9D
G@PUD73_I.6W8;ZAZ4fK(\2C&B3DR\TZ:2^.<Va0G)^9@eIZ2N30B7a]Lc&1D<QM
<2CZU;8DbQTL=<>?=CLEa=CBI8IX,a.R6d=_<Z;#U]7e_Kfe5aXRaeB]E1G-4O1S
C[<B.TO:^F.e6O(SH,A(HI#VJD;EC-&)/SWD@/#RUcD)ZK?8,Z.ZFUV13ALW&/-R
;(B&:IH\>XJZG7N9M+gA=?Q9?^MAGV13JLUDK;=1K\CfZ+[:4]V6\.^[8K2XL1SP
6ecfggbaK[7Z(EK,T-I<9.L=TPMbJ.MSWB.]P,1X98_Nda8<JD=[/B&_:3b?Tc+R
L^B6NS9S8HPe(\RIZIb(B;GU-=d.JYa,P19@S:^a<\ZCCK>DLU&7SN0SZ;=Q8:L\
8O)K^+8:GB76OY6/AL]A_KK1)E]d43f+CcH4WAP_AFb1H5Fc7S4Ed0YddNV>L9Q=
]US-GeA0fY>gGB98PX2c,9?>T>e&?=U<#7PV.KO4)TH4#4ZEBM;=CW(WL-W-F8aC
2Y7f3d?P.d8OVP7b1K=K>8IC8N0@II[T@Z[K2MS&4X,0FfPIOf;IPd-7UD>K.98.
Ac4Y05JQOZ3@HJKR+,S9cdSI>P8\0Y0@=N]>,_?d4AH_0/4NXGd3Ug]6)8PZOMeL
T(<<D4J^YGYX67K,0#O#DZ.J9Q>X/SX#IaGT-?\1>ZB<\Vdf4f:KF,,:-,-<FR?Z
1TI7]LM\efT7gW[S-=Y??7DJ_1C?/_J/PRg<AQ[0H-EK&YKS1&E-7<1<JQS97#0;
7QcVP^6Q3)J?aIQ;G#IPLC/DLS?3ST(V(4e-TUU@e/aQ.e;1#[+3]#JA[Cd0(U/1
P[6T&@9DMW5D8ag@S8J[g(?^.f[BB9f^>3PV8XA<gXcSL/CJWNFegGEf[Vd^<6&/
Ac#I]5ac^V?O9:g3N]@_CCKWTTW;KJIeeX+6c(LbEW9:/6Y#-+?7<8)#fV2IY9OU
gcY,8GFE[VLaRYCVH>.#Y\N)g]3.AU^+-/:_PG7+Y1/P;DS7?g4a0R+U>]g=dQV1
&U&PHOLPRgcFA7@4RbF=C]H\_E6b3O9(-^;B3ZA@Dd>4WD:]A_=bFA)3XXJT@Qb)
VS?+(D:XKH.:C[]?H;0F\G66^-JDO@GV73Cd+>GD]/JF?6C?\L@&W@&U7a:=a:>H
1+Z;RGXbBTg](H1gG#=8:[2[XKYX_C-(e\P?g69Ag3S;:H=K;Pg7eb8+.4EcPT)X
]I#+W.T7CU>7cEgce6XW[d-,cd_JFELAg5HNQFZY+2:[\=L)9.2X2b1AA@C@BNC.
XCC#9[Dd0K]4Lb4KZ79<=.:6-L\\=WL:MZ_X-.4<?>M]RD;EE8K.=@+O.b,_)1/U
AOU00(0IC1M&>SGGgRZD+XQ=6&+_/D?+A\:A28O>CW_.NM>1N^KMOJ\(3gP@UZ3J
DW\L+5@UT-PBJ>TJN>.F.&,+:K=[)\+(@8b6@<#\;QgUH<gcK=T\VJ8D;^d<))bE
K3.:OVNXH=?WY@49228FaE>D3D:;F2G)]QAKRfH7D27<3C<@2_<POMg2cT4UU^<I
AFSPSQc:+Fe?F_/]&<4[WY\M?7VCST8?ce=g7]AL9C/(M6OOa8]7WKSc>VeN^^KV
CAdcNI^2XPZb#I/64]7;:H3F&F<g(2^R\AK&WY4A0Ya\;AT:?\,RKW8BM?Z/DP2)
DDc3Qd/PW#4S_EX9cf@d[[.dPa8d:4MFWb3fDg@4He0#5a^UA-eF+IDVN;\#;J1M
T@D/&Zcg<dTY;4Ub^8Q1V29cVd-<5Fb2ER5J]1^E[6?[.(e>9RVW/1?#N29:#3#,
XeYX-6ZQO;6FC+,9>dS<1AOG_QF5:+3><?-,R0JCHDZZ7YKfCV/U]J/+fJQHVAA\
Z@<?>1)(IXT)),gK:H7GB0e.b<N4\^_JIAV>1M<dOP)VdYY6aT]H]6,PaR@H1NRa
>BgE[_1\O(M>LP3PL1=]AAc--<8L^aeLa+7d0QNMW>HIP3E_J=Qa&gd42N0OHfD6
>53C&@_28W38;X6^c6M0NSV0U=G59<>TL35Nb&>1#C\Ld6LZcGTaQN(@OB34WG]6
JM_&-SKJHE./7a.+D.B>E_[MD?:K;Q&2e8&1>+PA1LF<0_2-CbLf+XE8/(bb0Ue6
J3/6cG?>5;De0W2@.>B>UGIL-d.8;(VEM8g\JGOO\3&V)ITC5GM]Ac/??5(O1e2V
;I0/8GHTT]c:=<HcQPHX>XE5fU>0V,ZCM/8_Ca>8O<S#a^F\MaZ;9R19+6KRT;<^
UMU:+aMN/-b7PMQQd5U_#-]<2MLNB0Cg/^RM=3(D_BY2b2>R=-PF9T::>68fXAL@
U<DWQ(K2(d=e?)@.P925[29Od7O6XX2,V<_S<LB<,.>@YG.C#EMO5Q?/EW(R#27)
&4&W7N&(W/).FZF4SL-H]=66.=L2:\G;_JNH8\gaAXY9HF.Q):6&@DLTC:]&B#g-
,OfR;1JXG15<R0R7<;gQ]_DT.]MVR+<0A>f_;9d9CA&d,1,RKXQ[8](^46+SZa^0
)T_B^>Q\F6[4].)3]G>ZF61.^gU/edWH1;#7Ee,\XIM9VDe718Y-I/>;&X#5]?/T
;FCS9AUSL3\0c2RN(M0EWBeFd4Y/3@f0<@4CT4B<_9?K=T3AcX>O)^.]S+/Ue\[e
.=M?CVe)+ETf<;GR575BD.b;L9P2[@,N<OP9/BYe=^\BUAXN9&;4X/I=g;(;^-7V
ReA;F?Q@cTaZ\N>2_3VV5\1W:_I/4=MUcXd&H21AY6:9RHG)MQ26(C4D-4ALQgK:
,?:28#dTTCRHFL;]+_/\S_#ZTS);)2\>4D>>?((<W7>3d]);=OaGT-,HbGd/7[;9
<fX595g8ZP5J?e@5]A[LYU37B,#[/2.T2CgJRGYUbB^IHNPgTQ3a;SYRS#gCK+L+
UA>LE;Y;_(YK35_=Z:)16af)\KQBOg&>2a6BG](Eb>6G8/:LUXgFAbC9](ZO5+(>
0EFV(R_)^;<97Z#M/_27[e&GB\]]\UfD^ObD4\NV>IE?^\.gZNIg.[H6MOagA(OR
U>3B#_;e6gMS/5ANaDL9K0>+3GLHCXI9K>5[gTgMH\7_V@1M[RDeS5HC<gB@0QW]
g<Q/6Xe0&YcFHGN:&EO[e7?U2D#bDR9c=/d4Y,_MM2d?a,919\)P3?L.2eQe:3L@
M0WV^#P[U[O3.#T>F__8EN&Ra/.@Fdf3\>X(39R?>.SRE=1W#[e:I7c.0LB7^-14
KA)USdK\F-7=,HCZ[=WYe7-S0Ic;N62\#6\aae(QO6gT_&c0,>bLL1b174^&G1EM
6g83>-O_3726T9ZORAD:67<0I1YbeNNG530S>FWX8-Uf37<J=>Q,UJ?CW=/5?V:2
e6f#&A+Q1H<C;3AZDG&)W9>28d(#M-aS>ZeKIUM),;36a<e=3g_=N6/Cdd5X<Zc<
K#3LbJ)f@7_(;S;<)JTW?&2C+ZD&^K<G#&S@SI/N&HNDP/F4TW+/\Y4)(fC@OCP<
PH7:<,dY#d39>)8a#N<GX[Df)=1@]/@2NKILLXNPcd7D<cLZ#dFgUIS7^>C3UX0P
?V<J.4Mg6UAHZ<Z&DSXML,GDZfDfcfg=Acd@_UPWId4bLY3ecb.BLT^42N08PO:d
ZQ-UL\@AAfRbf;I>?WCLVKM,P6V,E=XY@gAA.Gfg;Yg#b1L/AG,<d,8f&3U1A.>I
4JO&BAP3T5(H?H@(4)@Rc2-G,c;-I>0>6UH_1Z;3^I^faGW?bdI->Z9_N>5D1/<6
3GIT2MaH&-TM9M,eP[RWLf80<\[F?0@BZ<?1H</>[G[6)BZ?/JAKO37&/B,RMRBF
4GHg(XXcCM3M(#5C9_1XYd3fLF[)V4;c=&3;H=b:(@C1g\X/)FNR;4\5SV3@^\13
E^,;0+Q/578cM;bO,US\1F^-bJP,<;aP-==3,H1OE9fVB&dF6#;+]RN2E3Sa[a9L
NX,ZUAK9cCT;a9KA#EAF#5Da+eMgP7-Q;#PC+IR\LTW.UT5P-a,RLCA3f->/I,34
#feLC>)Jf<Z1cKMO/A+4TXVdVVG25?7B09L(.CcL5U&c(&=,R[Z+\?=Rf0_=bETK
SA.^.-HCOMGX:?cg2[<NaF@,]6DL4GQIZVH#dZA2.:F,(#OUW_OeCd[&ET)GD@N/
Q]cDD4[bJZZL-M?f[#TRO5/V0(F2:bSE?S8FSXa1#7KaH>DLGb3A-__A6@5GY_2Y
cb9B26Z;=0Md=I]NPa.gXV3IT(VA=Ef=;4A[Q2&[:F_Vf0GOM>I;R.gaXT6V&gI<
,g_V30-;M50bCA)7S^XKE+&d14TJc\_)+[:?0G#QI,(_J>X:ReRF;55[e>d@VBb5
DLF0[-bMTH+D+SPS>K/JEO?bf54ADE;K)R85Q;dG)a0Lg<O6+K3(;-C6.QS@IGf/
>+=&^,174][4dZ4H1^S#Ld#R#@GUJMO]Y(>VS[UOf[_McIEH[6^.ZRGE<SPY[J9-
DQU1<.d,8=CNX2.KH[T^(Y60(LSLK?N94\:Q=-BecJUV?-Y@cbB=gETd><;AX-ee
e2<GeZ[WM<T4033Eg(e/5[&@OY#/R(c9#cP6C].=b>SERI4\P.X>),CYd8EGH3ZW
Yg#<Ig2D&7e&4:-e9,YWHAH5[+S3E^,b,K&b\V4?8\>WS2G9BDPP0KR_U/B]:d1#
Q,Y?C>G^Y7A;B[d5S&X[@TT3:+NLMX\O;g0VBT5(fRMD3W]WD87RTA-CI.+/T(a;
;9J,+NM9\9MM^O@M\g]](<6O<VAg(a21D-&c(d-=6]FU3[R5D3Mf)bggS\8DH&X+
=AFA+]g:43(W:P?HT(,U[G1J,025_QOM,;9_.#MVT1F1Ke19>F-B^E<7#G^+bee,
<D4WVT;_[,R[Ke),XA\J6YTX:R9MIYJ>51^Z?Td=&fXEM<G.O#WWLa-/@@]JcVJH
[.G#5bc67ge8KGAST@MW07FJg@^&DB]6e[8g/O1K1ODE_S/#Wa:JOC)M&#DB.Uc,
7bAJ;K>?5R5.7ebe9QTb+O-KH5bY]FQV0=5L6D7^,LCaA.N/ZO:U^:Z_\ZU[&4[#
#e5,\J-F[NQ-bH]I32?C8Bc-X20+XW\^E,&>?JZVO;)PRdd_6:]C8/56R._:_/Q/
CLb+4T_1[)GO/^I:If1WBVB8^ML@F,cU[M)FL7e>K&186?YVDMG(K89S>RaaZ1LU
<1>dd88cLBgI-;RJ+0]_EgQXXX_UECGadd\7ecN0>7E4KPT^;\&>HPaRe-KD-ILg
.2e:C-[MEKD8J6GK61#BgXe=,3M3ScHHENM,#Y<._(E9\/M6/FbG#/L,NT5_HU-<
2FF.9V>b&5?ZgY3\,0,Df(DO#35G..(YFFb+,HSP2Ge)DfO@13>dAf#dWaAa-WZT
J;_KEQ@dXca=f4J#]7VR8PV3JG-/f_,XMFQaQ>T>GK^QL#D_>O8^Q0ZA1K\G0Y,c
[Z043NeM?T4[_9e[L.^@H1X4-;dC^ecY\.2fI0>7]ALSR\3eYR:O(HAL&J-,UGZ>
O<M)NE.SZ]/e6ER:](]G=S6[>g;K]MNa)S@=@57XggF-G(O9gGO[2SdN^2+=_3B;
g7<+e(QW6aO\c=UBWAIQB>1f#X92bc_?]D::d^c8#,\#;]V&EeD#WH<3fe\fb0M3
:5+F.XGM)UP7dA7bWX^PAa23<.RLIE@CaR&]Qd\Q26)Y5[XFZ.4=PLW^+WJ+TQ-V
BD,f)QQ-)M-=@->P&V,FDc/5OaHgAB?_B+Y1?Gf_76TX(?FH5&335Q#A9bJH@Fc\
A>(PF+dI3MSa#:<9<#D4=].D(Igc1MJ^Q)D][6;EKg&B/2d10?=JB8^X(BK6##>2
[fKA-VSQN&2=YOZBZOR(Y;YVNaZD??7<WLQ5L#UEF<CfaF6WQ,(0)56Q=CZ_6TOD
4R8.PU+I\GNCJdKO:R:0@aUd=MgCL[NZ[;[<-^];ZdgfFN19;8V9eT]W#H1(9BBb
eK:F2FE.GQN9cgN>MJ#M5YBX3EUAd4.)2LT^aN(PAF\QKKa2A97585BOP<JQggRQ
I6-cdd@S[:;^/5_#-D@3bMbB4-Ra0PUMHKIP-/Q,/)A+W8#P&3YLB^)Zc6,7cZAW
>O+4[S2,<9[AXf00ZQXAI@d+>gXMQ2P0AUPN?O[Yc_6>N]cRMeA.eHGTOUR(I-35
38E5T<=aNP,I[J3>__cMLR4)H&53A3^IFH03J_+?XY^),K50Lb:QM9S-3D3T1eB#
V&88XGW(B[B/GT9[I#<;AIYF^AgaBFg0MYB:?YBH4;+/V9=Ib?;N;F,Qg^f/&PVT
3Eea@Lb#CG/H[bOKgS__KY.S[K1_5=d[[_S3B>QAH@)LTFY7fQR)XM[f/B/(fMcc
eCH2XOT_R@JDg#N?;gTG&,eN^EaXEfZEX5dT^9@4UBE&-IOcQO?VKOg.N7gaQ\=4
H/FGBU=/+IJZGf8W)2/APPSVS.8Ac,NYCWQ81#UDE?>I)G0Y9?g6:ZIF/Te\AN42
c]=@&LUfQLG42defL-TU1E(K635V/3KF00WUgYQRQ?\>HRg0G3=SeRG,Jb]F)FAA
Kf/6-.P\ADc@aD^6KTRZb]]T:/M+^9EKY#T=9HT.=[.=U+H8F56:a:U.#9>9GJV+
1?g<Id:R;C8SJ8V3ea^,Od77,V?8LGgCI-N9N9?-?6:<fEF?4IXE,6eZ::#;1BV.
CAF/9^:f<@]<GU,eaU2^\[)b,H:RLBd&\dELIGIa:d\/E9V>[dS52T2NX?I:b--9
ED0V.Z+,B#Gd[4\QLDDFc/Z.VIFRcE,YN/5IO,?(M@NeRWAV<cR3D<Fae4OC5B(3
F[@BWA#?KGBdI-OC;J,?=H3FDgJ8NKg8g_f/-<<QVeK9P9Z2c#^?_O_e#Obg81[g
,<)_AQbFI=Z[9O.XS[Rg6@dQ0>\4YB8\._1=IO+fcgf@Qf,K@&]FCW3+4I)f@<M?
N=:WEQB2A^d96FI+Q/d4)<)>WD-I3ZbUf2:TP@4P:a>B[S;7Q-=QE=6gHODU>KZJ
Hc)48HBfa^.TB)d:e2,2Cc\,/8.Q^66<eL=a9JT?g\(M-HHYaN:7:.5C^\-5^WI&
PXcV#Zb]\LR@5Wc;a0_6PZ#7-VU]cV(:UZV+5MV.C.b32XEdPYUH19IY@F)X8\;+
D9+^fY9eSgR\OJ,:M&3+2=,6T6FNUb;^dKB;cS+NX/4<@IN<,I)BBZD<Ed#?.R>\
Wd-KMO?UW(c&<7fbH^gVW_.]1GR]^<X7^.(D7QUK58HN9UJWF-W9E=a#,TJ6;ga#
MMG_FF(GH8]XD)cSe-RV,]a>cP#/,6g1@8,K,9a]2/Nd+M/:d2::O,SS+U6L,a<R
AQ]a\7<8dC(KT8eA7J4g?Xb[TDb00>BK^c1[KJ\b@UD\eXI+WU(4E1g(UaU.B(07
0+=[>S/gDK.;YcL;?3TMMI3?]UF>c0T]7&7d+e:)JYXd_aPG/D;UXgD(3)CdT[(H
J0=AZ+b2&F7S9(^V9&U/]dbR/Cd<bPXV1V170bJ2f\&^H/>U_?B:#W#Y&R>@02T3
]b].-NVT3T5@3\dS=DU.b08L^?S\9d21?-C]G-K&@G7\2D0:Cg\dYZUe)b4==T&W
>=E<^\[G^5Z:HIZC-aIMB4[JUPTJVY0YC:3fC(8J-AS2ga0/Z[WGSgL/]a[J]>:e
;IM-e,L7CSb5ZZ+W?_4]>Y&A8V\W)WGW;525IJ&,..CcV4[B[X;c[8PRQP,)HR0b
=AWE,e2>Y>)_ME/2GK+>&D9CO_e]/,_A8;A0[?S6P+L\]RO5+4LMRO.U^S^<9c)[
/[SEQZWZ40WV8)5R@>FVYJOb[UW(B.HN]5W2[G4cd@-MWX^4=12+:Qb<RO@G>I\=
=K:TGKVM77=BEdEMd[0_c.P988SGQGIb6RC?b1Y<N+@+EEJWTR\9S7_PA^1.?KGB
J:=,XU9DN>?9+C&R6]>\(]R>9,AMNGW1E7bO19=A4;?@+<bB#4DcV5O<FD0:Xf[=
[cZ2b)X@+OUR\f6a:>e2TRQ6UM2M)+M[P<cZd14M]Z/U/8ALf&D[@3Ag-BU6VaHL
<0S:/[4+IW)@<SIR?;T\MI;XYEY99dIP^IE@;+;aV2@b)C;WN>.PN[_b^R4U[I3b
2fP\dYWS7U(:=TPR63a4bU+2^]8Q-IE[S4WQ-E-#9CFXeYDS]\G^6-0,g#A:H=YN
O1OA5N1M>baMIRRW#PBb@8-3.,8N[Td,a\d,C+?E.2//bfBB#O)R,EaY:>.[]a(b
Z&f.@>NUC+f0KV(Q0^BD7),_^7:N@T(\A0\0?fffb@/EVb?@?_+[ZM,Kb&:]E_dG
bc/PH_X>6ICJ37R/)4&WX?S\#),DI<GC&)d1R^33KfO2,O0O2BASHc]B48+fBa2c
=0e\T>bf),4e]g[@Z31=aH\4gUQACR8Q+>I(R9.2PQ@[&P.KAJ_#Mc+9;D4;UJFL
XP.9f879XIB&H#Y.eNC\4;-[\[2OSe,G7CN0@MO&L^&:QJP+PYWPB4Ee-N26b[/D
fD,I@BbJfb,2U?=@MAE5U=U,8J>OgBVH=@MK3X,H0::Oc?JZNNgRK<@[S;-#6J&R
\.<.J-2aEFa_<<@P1V\3FI=KE-YE0_b7=9C(M&AeAHZIE<J0EV[<K&FN8W/VV/2]
U5_KdDgHe)J7W<)dAf_Y8&:T\GNZZ9=\[=08/[I>6@+QPA_(BW+:4C3fa.HM0/PG
-HfURR&_^J>4US0F>ABWTdRf)_I1HX(D&51Yd95LY>.Od+:VZ6BIg#<Wf4OX;6I3
6-W0/DZ=],V+cARK;)JYA-]E31Qc=g:A[[R7D3.?1BGH(f]U(G5/\8[8AQ-MUJKa
D<WRZC8)Y1<HPD&OT[L0\E;S[QTXFgVO[^CfE@K/\[_+_g?=N+,bIb\-]<Sd@=RW
^;R5PE83_28_-F>:(BH;&2#K;R,C]XAe+gFJ;7GIFU-EM,7[^IXN]11[7H96Q5/>
ANeY/ZX(eT=V#U<;XWcDVRLgQS&K0M&Q@U@K^\\Y\A?cE3[AP0+(TOTZ8:/^.a8d
Ef\2[T7[aHcc#LT_bM2Dff4NJE6T-NI?XgJV)M:_<2OfH#ENK8?#OO-UT4M_BU>P
-IZAK;fJe<?4N125+.cCZB;2P:4efH/R4f0.TJ5>#O0TQ5KCXdM\[]bBe.QZ:4BR
bUW:Y(U>W,LLP_HYLd<&Y0HP#\\-L>3g1AAb5U1.b5UX\YPR6,TDbS7P;f(d-;K.
NAK=#YV0\1d#[Q06?N;9f)W)?LQ6P1MI]?d:?X8-IO@(,AU0^W+bK1N_dU-:Z7(&
-QYa74^HV.=>c;:/56e+_2(aK?\7#;SXM,=&eT-]X=T_e+=&]Y7DD\VM[E)9fRP&
M6dM73?\>83P?eU6TeKd@<3JR&:K+=fef5JL0#_=f18<,aKIBOEJAK0Z72)K0W&g
)0-33g[94@gO;Nf+MJ,/Ga,ZA;/=O+=FLU_Y(-T^4L1fXG@[9\=5J<>JY620d,_-
=B24ZE#@U2BFCAJH\>AI,=OT/-=#W<5=SF;f3d&ILF^0Cg81\=/YaC+dEU)6gBL4
-EM:e#^0CM/[F#FC;JWJcS.F-9OQVNLZf+&P_ef6S.^5XQ>X85GG\g-YW[1aZ][?
f7C>T-QGZ)LYIO60U9,R3_M.66Hg\>N;122U)_Q_?a1<+Y<C+?=P.H1g?:C&MUBA
T/><0PYV43fb:(XLWL9SgWP.e:BRL^OS42E(1U=@++Y.O^X2BJV@7@Ta>5gM85L/
b)5J]<W)e+/XgS+:AMNJ/W@RB^37=Q]Y)D3II8OH8V56N0N\FZ-D0NU,-:W0d8B\
R4^:5X-R56\g01B.KSWF5U?C5g1-=6Fg6YD-S+f:;S^X56DY_8CT,Q+F(K]QAZ^;
>bIJA7GRZ94YYG0^JKNPA+YIAB;4(Z+/<;L6AWWAQE;8P]QLbc@d\RP)0BgddO+W
AX653a2(c&0(Z]FgQ5]BI>N]IBHg(7fFOE?>QGZ:b0HV?Nb/_=8\E(Z,;\^9H.Sc
K:@b/KM\O-R)bc?_c0>#GA+C#_@c=\5_J<LHb5J;)S9W+W,?G?]\U]X8C:>@X-Bb
WN]?CNVNPYd,gYcJ<=^.-G,J:5/C0^6fKga=J-]:33(O@?ZPXQTY@.FY(D7fcO[2
[Ke@bE3^?=#DE[+88gB(bN02f^9U3aS@W)L<9.@:QN#P\NP=L2Z:/fUO&IXQ43e=
24DSFd0_6^/4L9><#3NBN8G=VQ[^f7[LW9g5a5eZgF@0XRLAV@S8(9OQR/SAYaK6
-;4#,PU).S##7D@AW7C0N0EE6-Q.0dOWd4&81NJ&B)EUMQ27=#&IN[?-cfJAQdNE
@A.J;[68bC][bUf[/\WF15O3.UXRS^F2ON@)d(O8f#H(UV+3M=Bf.:+bgdCGNNc1
2D]NS.+c>1]N@U8H@/DH0S+)I.#U@UeQ1<MN5ZO5\_8?G,KZ3aT(A+N]I+(,WJ8]
Xfd0:.49[J\)[a4a/AI.:#3YcWb^?7dcHa/OZC[WgAV44;N>JBZfL(J-KP^2TVY5
JK?-.^LLZ&OS.gR=f7S-XU+;:)R:CGGSXGeWNO<I(FJ/85M+\Q[]L=Sc:dSE#4.2
EKHQO#)B>;<TJP#86CD0P9bY68^P:fK483+9<Ic,:8b90G,?^+G#T)K>cC8Edb?<
ZJf.X9Ye=fQB_7#0XX2cM,1&?Z/ZT.\/8@c-E95_+/b5<Ya)=^OU9BYO^HO:AHb,
<43H31(ca3>N1;@9c+N)IN7?<B&0a/.H10W1+dW>>_H)Tbe-MK]UY>NXTUfN>597
X7D&2_XV;=(U[KS;f?C?SRWcZ?CKT5LJ@:#NKB1b6[1L[,MPO&XD(91ZGWQ^><Eb
RUfX<FdbNeZ,G67gJ@0S8^V\e[_O,fcda/SeKW63P.>I4B>2E4bL\P=>S_<Hc++=
d6;8\b.)EDbR7UK\8S34;IC2@b7^OH5A9CTFQPgB(N^VJGR5726W89^9^J^\=?VF
[Z.7,V<@6,C>_,<-I:F99AQ(02UY4E(8:)EJ2WPCC;;=F=ed=\)_,4:F7A=WPW<<
g[@9I2[.4HZ5.^Jfag30HQ5f])E?cbc/5W\>RMH)54d=0dQEBL:QG45KYbRSMEOO
bK3)>MX^EI(-\0+/5efC&C4?M3HR_PbJN7#<Sd\@M<Z]SQ2(3.Z3_#\<f1[,WfZ=
OR8/:3Q#;0TEa5;2D:)PMX]a3B@_-f^:7<6QF,_Qb<N+-a[7E?^fW5,Pe?9(5NJe
EE1GDGS(MKB+cL#>8\IV_.0K_:750VQB6Gg0]=_FQH0?)>)dgG94bP?5b1OATV9a
2(.Dbda455JZdJ76?UJ9ceG:)?IRXSeNOe&E<1[]Of7EYS6O3P-5@]-P>R<dHbf@
FSWZ_:LNXCHKM&:a4]4^(KX,QE./HL]A#?,H1_\8EK&8W_8-WfI\66C#:].Mb\cC
VD\;+X3PPN&[_B\J=NV6JZ+4.dCNe)=5,):(0c5c#MZYB9=O[?;V<b0O/BQ&5Nce
;EVMY.Q.WD(-:3K=a0)Q^NZ=QEPYC9WT[TL#<0>;[DV4RU<4RZTgW7B.0b))-AJ8
c:C8I?F=_6d&GF3g;dYg_W0Wf3E09B#4]H0Y.K,]V[a@[EWe7V(^D&2XDY2[UaSB
3IE46;B;B<GZ&>N?]Af06R9U/H0@Z[](CZ4-(1QK1.4Y0^Y9[1\<R:>SF,,^AWP>
0_1DY7K6-O46dL82E_DDKO(&ZBEa,U;7dEELND(4Ld<NL>-1I1-c_U8R@V1&04XJ
?b&.3gcKa.OMZH27fFd>TU\a#cc)_#:Xd4=J(7,7LR^;^ZXIgad?;.0T?/^?S5dW
]ecLWO^66_X&A_A.#9UHADWN-R1A6B:^HL];Nd)eD>7_I9+#\=2_H#c@UHICY=1g
.?[gW-?YfY])Z.Y(PD&K/(N58PfG5EH@Q?Zag<5;P\Q_cXa0\,6g#Q@Sc3WZ?VB]
L\4C+[0NH):=6M[PNESUd=([?@E6I]9aMRGC<c[+&>?b^5QR:&b_RK:+c,&Z1(4W
^?6L#/5ZF=QXE3YDX5g5c6OY_(S?]RGA=gUG313V1gCg;=]BQ)@C1SL4K)/D0F_9
e.#QNgD0U=WQRI>&Y\1A8F.dD_-U7Q&fSGGPg9#bf(\IFLVNO=<eW6fd/3a/_dF9
E/6:INeCLIB\<FF+c8?6JHGVN,&BC9^L87YEd0TQ](/g<7A3#SPc^Q>acX9L>Ve\
<AS&Dd:NTZ_GO5aX4(aY0cVP/=@&NLfZ5P5,&e7=^.+Efa\eY>_S[0P2:16&JY@3
-4AbJ?0;\@C)DGb]YH-cf>ee#F;ZRJa&RNeH8FEdW=HGZIg5>D)^>L#NE#3QT]ed
RJ_fe@Sb?3W>SCB?[A?25T4c44La9T&Cbd=3?J>W&MdA\Z(XIQ@V.[bV7bC26@dE
B1@Qg1I1P,;NWaT=04V082a#N&(<2469X@F^a+TRFfMaPY@GT6.V^N#K2\^Y6/f&
U(/ZA^3V9+=YOOARaKW]L=UC;7+;QV8c&(1I)e2c&^0_V_5)64bMB]\fA\\#R7cN
MF;CEN@R.b0(7^VV-J@K0]L[Sg2L;R3;U_Db[>U_U1K]<8=Rb[;C1:U3c\@/HN]d
1ReN(0:[7=)8;\X>Xb-a/0ZQGWXA.CW1a72O8,E?TX@B_4]^53<,6b>e4V\eMD#F
&f4fN9_DZ/8T:RG^STcAU9+W^[=U,e1QM4/db\[aD\RbWH1[KJNIR^+TE_XaH[X-
MDO8:0.X+AT#>B\ZP3<Yc&cc2]SfV@XVaN=1]b\5_@+]Y[Z4B5d<JE&CW@)NOBQ^
?8Kc,X\PR21YFY?15cSW3H].0gH[5,?@d@1DN6MJD15c^=JC25c#DX.&eUdX>=+#
A=28C>eE7?2+/\<]8<=.[MRNWOf^PGQ_@[>80.0L1IM\#M2A(bg^1bE1gQ1/]RPU
U3?GIJZ,B6P_;44;Tg.U=J623OK8I_VZATODD.LVKM>S]P3WO6;cf62I7^FOJ]/b
)M^7MI64D1\QI]Z/(>8=QG?>-USTc.NVU2#]OB:AFcZ[Fb1/PY.[^&(4QF)S54Ga
5P;:6=a&7bEHYb?:>)]RU,<C<8M\2]@Q1\+0P)/FJeWXG5<Ma85e^^RdKW2@Z<b.
_+RX=-39WCg\XdGNY9_.9^W[/?JQ-1:X1dfJ:+EF9-,T[3VR@JeIH7V6CVeg8D]c
aZ4Fd@.6XEBLdZN12B<RL(NfM^KE?WWL@^e7bJK-Y,UHQb,H#;?UGE@Fb7^7Z\,R
V@MAK\_/c:8\AK2QBE&BF2@cWG\FK#J@:<&=QIF^F/^9+A>3RR@^KaJKd@_BK6CV
RIN4>e3BN_^/2\@,[RFbL;:I#4SWL\Z:Y9#-DYA)\^91[20?9[3gF/DUS\?W0&,a
f#X5<89U1Ab_<[PC[<?.e+d#<HdMA[PT6g=B<?BF]\-57RF+,g0O?0gOHUVgI<@:
b&;P<FVR];T0DKR[c\7G.5TTNd>B6dB?,(#\57C9+BgMb8fQ_JE^T#=N8g?bB^);
TTIAC.O0JQ\eEM9.S_#eN9^DHD3MW@(D5^47A^=a<g?5ELN8\G94J,eR.PAJdCeH
.V-5_(4aSN?VRA(+d=5fDc@L\Z:a/NcO_EAYdS_HQ+_?(7&P^(-QQTI#E#DN66eX
/6E7d</LNM4bZX\RL=f(P.f9\>6BPQDW>:_UN@]+Q>Kc,GGYWDMGM_9#O@H2?&2T
I\X@M[5(1G#4LIS8S-OX_,+T^:8b=A968C;Te/H:a3N_HMeWa+D0Y]U/P>/;<]VN
X(7J)&A,CfD#&0,dCVNf.[K[CHaVS>1DX&O/JKX2F0VO?Q-]:.=^N\>AU7\D<A_G
>ZFedI[Z>7>>/\e1SH+M54E:47)X7^MCY8)-gGd<U[N&>NK:G@RFHC8VH6FNOYRP
,gVUeS8d50MTP:9C:MPA=[I093BISQQLK1B5906;X85C-NV/e;4D[YT4(d_?M?R0
U\)9^_d:QGcb.U3KQ-(3P>_V#4KFafdc=M#D3,FcF+/@)=TC]?&O@YeJ3)cH[=d\
3QBINfSW;Oa-bDIR(eV9[(bV44<5B4D6,)G]U_.g&1R3F0@=8cL[<ACOW&FYZY55
/SZ#]1:G+AOG2.V;3gAg:]2G7fL,\g3fEBX2H8#dK1W.(-<bfb#aH<gS2@8J)6V?
&C:YAIN+_E@B0gA8ZF/W-2)fHKQ)SFR,&J,Hg^fN]EgYU(:MO0H>cQa:&2M:89;R
e4gJ&][0RW47CXP;d+@?EB++R^;d70ad)/)e7&S^YLYBIdT4SKKGdA]TTc+7D:W<
E3[:,NF5?J:XUJTQ@)ZFO,:F9feY4\.W.N\K<8:4-;_-\1MeYD=,5++Q0E,E-4C3
)O.XO+De(c,\5f=O/#b7ZR5+A1+85a(M-Z(7523[ILTFL4V?Y@P2DH#7SYMK.TI\
@V&f23X@O=bgH@LV&/BD]EOU:egY1K.L.Qf]:@9QcA#RD4#X46/Y.I<8YCXI?T.B
G9OHgY79,J)41+,5:L^BgQ?/SSP<\BC9+JJ3gT0O&A=RMIWCT&;;AGTF-V?4N<LC
[6/^F[@5O(,H1MEF2,:gT[_YP8_</fcSg0YAH)-\S)^=QP:a_R68\BM)CbDRb6M[
K6\)3C/XCYbK5W]0X(OV,0XHP?]#[P^QYGR4O47REXAGbg;X3gLMWFR3Fg.)?0@^
&NZRI-,dg(M&3_RW.B(RV))c2274:NX8SA-][XAbH14]BCe8GAX;ab;U:9K?5JdI
OGE-IN7?>#=8MIf^((Z@P=YLE)d&E4<&>BQ:UA)R2g]:,\S2<>IcgefID];WR^d:
6)-Z[e77Ja-5SG>;<&W([\ECC,5ZOXJf4E]d4aX&eRW\IFQ?Ag4aWRD8AM>dF>OD
N;O4U\X#a&df9=3_WP9LE\978TH\9fXARJM9]DA6T9NP,MVIOPXC)H^9dQ0G8B9:
g+&3^E:cT^G2);&8eV^7fH?HZ<5XH@K7+3Ma)(747P>Y4>S<ENZQf+Q>60,-&YYZ
_Q?LQM82H+R,/-HB0e@:b4)1GVXGTRDDJf+B25DK\S_Pa,R22.X8?\JgZgK2LIQ@
Vfe9?A?9A?DB.1a77_d7c?G;g^JA;]K>)A))TV=b5N<UKG#Ze8-9LTTRL;M4;UFW
Y2_#[#-fI2]91MDT>NBPIUcDVFOH6?NUQ3^+<^9-:788-[aP0(]RPE2G?7,@VSEK
QRQDA9VH)U3]DgE/C@ZBRT/P34K8>>CI6(@1#9:ZOfT6E]cLg.a^/=bDJ2WL[:-+
-;/_#IAd#g)AM[?#K<G,4T=[7:4YWgQ8J4gW5F0d;H@,_2C<G?=70e^c6<B:[MdK
9@>CM2edJ;]T[-+[Da1d,D3/cY_6>J.cRZLJW)[Ie=2A&a6-HHFSEO19P-,],<>f
]GeUa1:aM>FQVg49XD-[5?##fFFK)XAK>1M/_3(7Xc/_MZdHeR^/<-\Ue3086863
eXZ.AQa8P?[C>e[fDW[QS89A\d+Z6PN_<X__,&&=)6SHA6+W+;Of1&\I,;cO#15W
e],0F<ZXB.+8>aaB@Fed(eg0W)T6:(^\80+eN43X><e]fU7gDVg]P#XWSOA)(c?E
:=a7G#FX[/6#IDF>A_Q3@<90DZ2WPROGf>-=&N1^@-R#B&=8.U+@#)Wd8JbS8#CP
B7Pc(JE/eWTS;\BKe;ZW1a/eO]L&,E+B4SLW79@B7:f@_LBGEA#W9B[R5KMDAY-<
<+9G5<4CPSaB+c5)C&NX@G/40P#_L;e/#VO;O,L)g]FbfZ6\aA;Y4QUc>WO+^7Ac
)RA[g3F6MS<Q(/9G))4E?N@<UVeA,TNEe^7=,fJD\-PeOKGM=YMY267aH.4R]gIF
_H_4MJMd:1eD4;.FeE=f-9]?P;OdPOAJ@RS^PRa)RWX<3EH=]R6G,-@DFFY?]=,V
WA8K^]GU[.+7UU;XY/C8D<R/;c;.,4eP7RF2>/AecMTdI1>e0@bGEe=WND-<_.R?
_c+b+dE1@eKDR794=QW)7Z,?SAbWTUGM)Y<+_+KJUCQbe2>Z7P9PR=6V#A&:^VO(
@7UM\ME=d/ULG;YZHLC.71@IE?E48YJ:aO8.CR#S7OW?AXD_bJUdg51Re7=)E,7e
)&8&>5Y1Ge>.UV77JP0GLf1&,QIYS:eg,H]\/Q\79@R&g80C([9Z&A\5f1Ed)];-
H1@=N91_P(EYI5NXE2-/8L)_ON3D+@ff>@CYKLJ1VLQQZ<P#;@a78[F3R_.M&J;T
3_):,A4@33W\]IF0:&<^LaH:^fKS2f2EB/c:dA-^5O(ZQd&IF@+9UD>^)+cDJ,ZL
[&)CYc4>7@ad)J3J,S28EV@C[#<4GU58,?NCGDcL,aU.)&Nf7cA/,)JNZcY]EN5d
MJ7f?(dA,<2;4G]]GH1(6VBZ9HL.ED6IQ1(5ZB6ULQ,D1?bT[-[SZP5UDB#[:.5,
Ue)Eg-U\K3\;<?-S6?YGQ<8W7dfIg1<H;(CF(X6/d1J]U4ggJFEYBC##PN#_@JG\
#d[7#=#G55geLGY8^H:Gg<KVd]&V@B/gSc-N5,8)QJ[71:0f>A@9S-Gb(<DOX;28
>GUN_KG0><_a^g.b6,0d&8bTT:6JI^D,]#dAH(645HO6SUSTJ-9+&.Rg>RE7LI&3
V5d,0KKOEe]B9@H@5bH1+abRJgB;:Zc31/=-/c.[VP?c9a#]d#&g;X&R\^5^D[DB
/^Re/g6\5T?aQ5T@(>JEgJO[L:70:_74Vae>[U14&GW[/F5I5)7e27,R#TEM-G/L
H<R<I<N&O)P-=(/_cb;L^,\13,5D3OJF1,,P:Z^;b=+g0,5dDb5U&NK[E\LdNcXM
5ID>Xe30PPde13B[VT5bYe-BLYTDcDbd&G)_CR+?7DLOSE#?)90)()_4E2(^E]HM
Q5cAYaZV]OG?GN&c6-=1M\gH0+)\F>gJbBH@MQ7=L[)Y]\4XKU&Z_TK?11fXaDKU
9Z0:[SFL2</M1Lg.9I(AB8V/_(5XW?/4Z2W##CQ>O\aJg9CDVV-@&:cOD>eMKFKa
4R=WR?J2._S^=:]gQ;#G3>UL=V=)TR5_eK9:326Ab2G4A53=HLH<DN(\>^^SVM:;
@=K@BQGYCGQ9EdKK#]NPcR>&#dLXb_2cZ)@/;G?PW-5(1WS?Z5cZYV=Hc?=[B_ZH
E;b,1.&21JXV5?Qc;IZ/<YcRU&JMSSf4M(_Z#-EHcTA.(QI-]JP.eFG-P.fR^<NK
Q=b@8GFZ:)6^\QPP>DRL,dTP^+]b[=P&W8V8Hb.AdI9)BH_I4#N<5bGYE<D)O]Z8
1-AS(UX0T7QK3\KT#PF.?:T>fN#e@7;Z[[;DUJ:[7L>9@IfV\]4cBY0&gJE-DY[+
V,-WXObdd6#VNFP;6[+X-:DObLGP17&a[C)e-,aG34<=:\SE1fE3FfG;-Rfgcb;c
]VWC=S=9,O\G/SWVB-(@8B4VAc4L^?(/_^.#YUCNTL89c2W45=A6f=\T1>@DVK#S
YW04NY7T:\P\Qa-dKG\++UMa:X;/3A[.?DdE->aA?ML/c8HJ4-a93(]9]bQ(A,]#
C>bSe\,M6]].F;b,_)VaNYI7dH^9>D^JaW>EN(\d&,RdJPR>V2BGMN.ZY1Q^O>O-
b96f-Ve7]:bB#&2@#)-f+JF8:)F=[L\-e??>eKB<=g,Y12X1;-ZQK3\bcf<7@U0@
BB0[5/aBS7B&BCa7MG&QFfN-I#IG17N0.N<6L<[=7C6GG@G#-)Z?Ed2>YeJ43Q:c
>D_[4]\&QNcIf]f1K#7RNKR;_EF[dN?A#_3^E:)=<8dE7YU7@380;Z<>bL4<YHB;
=0<Q^+<?NK+c]=?dIcg^4bb+.GI1564@S?dB#/]-.f3-8AXN5c6IaQ^_]G#bLYHZ
?K,=^MCEe3HN:7M^W^4^VdC:e)<?Q[_=(6JZA\85732]](PRBfTTEDRb89^G&2+O
XGV&Af;\e3ReRK\A&6bgCaFe+6J/C#38O0G/f694+WAU5JR_<B)[B]G?0<^8);=g
cIK2._d^Y00T73XJZJ#f9(e0IVTg2QO..(F]g8d74)OI]F#<>FE9MW9X15BCg+6J
d5>2;FK+>MAY@Lc[P#fX#QeGIeeHIb:0-Z?WFW=.D^_5[S6/4LOJKOQZQ9#T\-:V
L^^OG().ITb9^CZ4]J[Sf.^fK<H[4Q(ZW>+B4ff0=B=(D\5/UH9NV^c4PYGD7GBd
,NW[58GPfgR2CKSMGaI(,.<8D<b.ID[()W<,E,\E?JV^2;2AJ?YYb=dRIC2K6-5_
@\V?N;QQe,IRIE\CFU]4_Pa6I,?MSJ:Ne)<</0b.HH)fT]]g((T:EHQ>]RKQ[Sb.
9G_-6ea^_bGW4c[W6FQ=:PFfBcGO&4U1C+\,(-8,dfB5-c,Y;76A.=3#dWEcd5/P
N\0.,eE<Ya;EA]9Ef@WDRPa^P^ZNWX.>O.@)G#>9.+c2RZ^V1JG[_,E(M9;@NU_Y
cg+25/KQS/G=[8c^c]+G[@IYZ15[H@OY[6Gg7Sb@D?5EH#.<&WcSe)QL<LOJY^?7
EWFgbQ0Q.U@edWbFa[@38K7E1M27Z/dLAD-c-f:?:)\2I<LMDB&#Q24(+gX2dc^b
CMRD;<88X/@YX@6/@N@PGMeUB;JCgGOM4?)5QU2f?G=g9S<UXI,d7+fJU@ED\LTH
cFB?N)_Xg^GF4>=c@[AHdaXSb=\FG0Se4#&DDg9)cg46#d,LH),TgZVb)/H@LCZ;
D+Ua8OLa#2ECC\3&H?I]^=?F=FeTAHTGT[ZX;fV<5<H9S-fe(RVbB31<,S6(U0RN
4N_d<=6a^ZcEW-&:6T>7U=UH12G1ZCY3_Fe6-YZH-5@Zd-/4PX>.e^UZ>7>eG:)c
IRGdC@X)].c-C5-6&:5Y5K@<LF-\21g:=7XB&Ad1M2.E(fPf8aJ?_]D=0bW3N\06
e940);9K6?9:RJ\DAZUc=&D0+NgR.1dB\I>R)fMd0d6)D\WLTb<V0MF+[2gVeM)B
;OI,X:]@X8e+c[C@5L>C5M+Ya8GCO(BF2#Z75b#[)W7_M267fS+^.D:9EHVaOFeW
R9cE?7Ne=B.J67Ub64Wf.0.efd3VXC)@F)3[ZXdF8BUG^:)/>5Z64L(f3(:.-/<G
)KYd,SM^0ILFW^B,^L]#KGZ(:5Y&6ID5&8\KE8cZ4FF>@7XI)^bfY;bcH659P[DA
3R(\P-5SUK>b2DZ[6I<FD3#-[(U7ZcdJG:_YAQU6F0@\_BE#;S,UDFUI<aH]cA]5
T@_]cDaRGM1Z99/>:F2VgC2LR[7[DXHfS[U1G\TePMYH-FVHc#I=HPQ#]GL\J,d6
X@H[O#Y^JQae[CKg[_0bYgD0fFDTT;W^ceZ)TE&\EZ?[f3M4DXa0?^B[,?D/HXN&
G&CNQVgLMc>94IHN9]-@BK)&Ne[7)JMVKCA)B+2B41+:Z7b0Z[e;^2#P((TT2Ab2
V&<B7S.9Q-Rgg;Z<4ZO:&+:GR_LLXD4af_O>8N66PO]E@^;EWZgc.b(<RC#W._+X
3?2\J8LJbCO@/e<HAMFF<>aa]U\SU?0LK7Y]<W^.]F]bW?6^f:;Z;:L]TY:a9#d+
aH?5U3Y-D8]7ed1N3<927ZM92>0R;=N3;#eFMS)F[2YQ8EBW7S&EK-N3FE,9#(+7
\43GGNVUAFYCg5Ra4[e.-E2fFRM1/6ZO>6RPb0KAT:,:\[2D?E85Y8@2Nc>W4#;C
2c4<c[WT+M1(+^O3YBOf^/.0U(4IH13fb5#H2HbXIO/a\T3Z[P=b0=I4GPC)bX,7
TVKdV)?]9:)?[LD):X-]aTF#BBX@([Xf.:<Mac,[>EaBKbDeXCeZ.05OVMTT]0U+
U5P9e7[cV]cVIC8\INcZNBA_D:8K8F55G:MXK64cFF(#Q5E,]:&#([_<7&)6VbCC
5fKUD/2;;D/WP;WfAcV>MgK(+B8E;])+6S;R-B6,6NJ#6^XQ\Q9ET3=>_7RX/\b+
2F7+CgT8RM(#/H0gTJ&TZ<9XCOCH,<]?,Q)C]:MH0O<9TTZAZ-MP#,PW2VTbUSfV
RVD;Nb[,LCLGCV:)a))JYX97[RDD#[-f4G?.(]BG^#3>,2>F74PBRQEJa;VH1?;1
gH1f[E613HfL8@#ICb6(Eb?dZ9&M\Af<H6O<?M@#g+;Vc9:MT>1C#]QIDB)@B;(=
PT,cGK)eKSW+N1>0)H.X6?Y\A9Bg6e#,<(D4,\O;NZ=3HG]HM?&,Q+BDE:6ca_d&
::I>)Kg)NfA+AH-2JMg;b;=?3+LMT5bR5a=XF)7_6OGW#NM^7D0.9B>L^-P)0/bE
2bQ0W.afKG(Ff,2WEE82F95-K_JVE6LdE[5UL/O&,6e5QF^Y.UFLBZY9,3Y9@&._
/.]CA\(P6:+5cT4PCJAbT:WQ#7aPFC^eS4OK4QOc;b@ZE2)K,)c?,2OfSF()QcI(
&gU:G[>_1-;,Y4W2/[?U&X6a15A3@YOP>==:g41C+R9@A?Q9bQ&>a+KC8X<\EV/J
NB#:0S@f1)gbW3bQ2]F;C=])3_Z+HAc5(JT(,2bGF;Qb\KG-?-84R-TI\1OIK=Lc
(e7=#8D1VD6,1:A+F;TZK:1A/.?<V-(K0IY\HE<WWWNTC58XBMa(LbA]4eSX&&g=
VH8=[Xd++<g<A#/=>VVQOI@P:U&<M5377d[R,728ATIE71D8GH_+Jb6dN]AT=a=C
Qa^7@=Ha<5-#e&5AC(FO[QB^TB\J0fX@]KcK13V&A2>UPA_O7X4(]6FS0.BR.6P^
eL,6LF^aXF=cJATF[,e7;TR\LE#gCA/H:(S),R<GXgG[?E&^K[#V&_+L19YYZ[N^
\Yg;I36V;If//7KLB8?ZRf&c3AI-b24TFC1PZQf_X2KVQ=/aTZY0S#[B@03H_J32
(>#T8EPeR)D-(&(99J;7;e<8255[1e^Q5_J-GOA<81dOQZb>AACL.KdE=A=WgKc(
JJC5(2f:9+6;\G9.IR&^ABAP.6Z(?7K1KT8=DT(/5]R@/bJX9Dg4_B36PXBVF-]H
_1&)Z63NP@;R]0MC\KAYCg;YNN+831XV8,ga.+O=@KD_,Ug-b0Caa7Q2cf(a6^U9
VGYLQ1E9L,A=Q94;6##)\XG,4,@6=/^G3Q;cATR/+0eRaZUe4\3ZS?S:S5e#gfI-
Jd/1RYQSBF])/b<+<@XgH0\(/e0VQ)^8NZ@TAF0K:/a6Y.SN..-A=I4(8AL9K5H0
[XfYR\C;JEX?b;E_92U7D&8C<2-QTNBcWQ:@4XB3+cd]5\AB=VNeO5VG/1Cg<SK<
1T;N21;JMD1e,Ia)NB42LG5MdQEaITJ6TKIe:FLVKB@Dd?fKDLE/e8,=/^Y6#H[2
87gXEa2Y)W@Ea#\MVM&ONTR-DA9O:NY04+A6c_g-S&^C/bReYbE7)IX;)&\1X2cE
^X]/\)8F?,57Zf2C&POC\7<Y31TXcIJ0g[9W2?TgUf:NeLFMKG)<D-g&^-#^?&0e
^M9SI5=bDT:dbEaE:d._S;REX>=DW&&]O75[;)P3Q@>GEG,fH(A9OMMWa4P6>[0A
5c<e7<Z@J]K.<J>XbZ&91(f5Wb+8T_HJfJcK.L=gNJUT&U4^(\Y&1VHZ=-33g4TS
MG=YL+8^VZT4_>]@?PH+7fU(#LES:beEQNCLMCSNHQR).6O+VG:P<_2R87L+92)d
YeJaN)]KQOR[IIcC3&ga;OC)U^FBb2[XB<Bg31Y@Q0f>b1-\4]D(PEPJ;A^37IL(
F6aK-AH\AD/6..^4;,c5VUaIT;9JA[W6N+3aL70fXCL34F/aU37&:S2b562DWK-9
MW-MeT&&#;6fOM9_T#MGY+S9,aGF+1bC7>BDfZa]D&,Z#Ib:?SDgR154a:YAO@+?
AQ3AXM_6^6MRef<W-3HS&.e61TG+)E45SMf7DS)BcA)_2O,fXJ2WFE#_7A0-f/3(
C?b8fMGP,(?_\ATSQI3+7MaM68.<\cCUGMJQ[JGK(V:I_B+5_J#CL>Q\(B<4Q[>a
Ge3A[G&PbE+E?#VJT_d(>6X-CM]N59&aV+CUfLR4@T]^;aOCOTW+6bE<7]\RdB#I
IX_\54L60T)A#<_JCS)/FdOd_I?,eLBD-6>?#f)g=5N8:Z]:CB&BE#OdX5[INc-T
MCFWEGE-BQSCd/E?V2,:L-_GOXb7S\K\+)F58],/N0#D3:,;^=-453T8Jd]/df^&
eT<Yc55<X#42eXf\g0Z@K5WR(2\gE.adW&Le>HeN0S;cWM(53@_B\d4-gc\SJ@]8
024Q#5[[R0Q3=Mg[BZ^RYGTD(Q]P;G,S?GXY=BP>N\YUH1LX8JTD5,P-b^1908XQ
_JJC48W(L5C07c^WH++>)(c\YMdQ+9[1_He(/\BeY^gOZTV^d]16J>)baT7(7S;A
_Y@D<4f?2BbXc/(IPGC)FZ/N0Y3[)@([,Z57.e5+-+bC:^a1&51?8D(Af/7P#B2&
(T(62+.OZ7AJ@2Gd50d=_G=9W5?+WV]].-\gM1/I[d<c,U<;M^TYT3K4S/)LPM_>
R#(7WDEg5=9=4IdfP9FEA/N69RC-6b>ce18#_f2S,3VR=NF_V0WfQdC:L4\<G/26
<C4.&:8/cV#.ZQSXEg[[Y:<,9(d:=aWADFZX[FD,-#QbLMXI^SJ@M7C>LX7I?Y^G
=;CD?[;S>\G016><SE;TG20AN[W@EGJ2N=a=c:S>A\B<e\@H\RWb\-4Qb+#32Fb?
UUVcI/B2DeAP)(^^&V[ZGCH2S/>T(Se9aIMRT5::N@[6)1]RFb;:XWZGDQ]A>S&F
ZU#L\2X[:Z_KU/)JWF&d9F[5-@V4I0GL2288[&de^O:-e2WU9Sa6_YC5]^P+FQ0Y
+8GU(-C2GYae\MJ0]D#Ng]:V/EW<8N;g/_S804?UVH9)-41PTV1JDPDbb]?O0])9
d(J.R[C-F/,<3ZVV1];87T)bcaVgQEC5bA/becE;O-PfV@I[;L,CJ]VYEC;_EKGa
cP(aCS]Cb>4F8HZ2Z<Ac75c<B+B8bDaHQTg-2<AKaQW>##9F#HS0:C0U2Z?.aK/H
#E9F7fFJY68=Y.2V9/P6<XZ):34d3K2K>d9O<PB,d<7[V+G3:&X+&:I7eW^(;Q>Y
OGKa17-78;7TGT^II36Q],T4^a<P-Cd7N)NXg>B[RE851,Hc+a3b6^gF=\Qg0dE5
Y@:V>Q1.=@3fgV@W3bMML[\84OQ/@@9:;[F=6;@CWE0(=SS1G.29Z75-(YB1PdX)
X3\3LQ.^5Ff8.C\Z;J.E?)Y&bR+L-Y5F]OPW28P=C6RT.9b2+@ONJH)5J]5a5\WH
ZU/-X5A#ff#>#Pd82Sg:eeCg.9^;QH^f639f,L31ECG38Q^>0JFA21a4(Kd6@@,7
SYgH0H[&M.2.-<)GG3ZLIO5JQe3>\LU4:2)FUf5EeOC;cC\DLJA3R.S=DaPegW4R
3OR.(WD8:LKQ<Z\KX<>/)C9KbX_K@(cQ-#XDf1FN#fE)_cEX(a6)>/c],@^e&>(W
f1+OL+/T=d:\dC)0HdWJ/V=XEQE]Pc8Zg^[L9b;<[#HZ<M\BG7QZ]+D6?_\-LE#@
fC6P@bFa>BN\UVW>Ha,eKef5aGLgLdU@[XD)9,:<]ZgNS;b<N&V_Q74W3f?-H#P^
79E,?GTS]^#CcH]b6C@cZOHP&D_;e6[Y&(L:bUf/b<:H;K3TO/I2Ea34V:\2C4DZ
Y+]](_aLUd_]Q6+bJG5O(RR&A]0MKSX(-5ea/>-3VWI:EfB:5gQ0[4Z^&+e;g]5\
\,+X12dO>K<S/ZZ49b-9?HfSb\U;Z,,d?@S@USO\#IQOC>>K+J6cY16QG6//bHRC
-S<^K0G5R(?M-HN,bL7./789;GY-@@;c]V^81)TZTD3O;dIdcD3SeSN0d.Q-VY5+
X;D^eX/II&3H3b9>3G(P>Y@ST>cf+7&EJXA_c^UDGQfE80,-9(2eD8WRJR:>ACGZ
R5S,N).<dA&ENX))R]S8gI:#=#9b.:b<d\MI-.-0(aFdE<0KS&g+;gGLZW^X+GP=
O4#YGWQ4eA/K+R-6UD23:]F^b+:efYEU+GJ176gKS0+39N31Ag.+SBVLJBga=LNe
;)WG2[E\cTC2?A&EZ3Y4?Udb6c&J#.8+O(aWS^,\@3(f<J;IMP#C1LTV6<d/7eQP
#GV,1D3Q,YEUIZYQ^G0:47];\\U)3gO_d07cV]KH,A^=1(@L(7d_IS;B/6TUQC(_
H=J:R=P+0:S.@1cfPI2:I+XK.J[95c3deA4&X--\=F<K?(6RVPG)>\E:#J1[fK80
]@8Cb9,6Y[fEJa_aKB-cBPbYYO5J6A[ddB-/E/,?#;;4O<GTZT2>gEdKT<DJ:R[c
Sd?-EQNZG6Yc(Q+e#HAQ4G\dXCR7II]JOS?O/H7,D^)d@M8.J/<;d1e;A53g\;2M
N\Y[3Yg.Y98gX+UgfR7:T_>.=E4]2Q6Y+^;>JWT&JCfcP8+^IA/GVQ&.9/.JdJW_
Z.,6,<EUW=6d>PEWL--0#B;bZXDZSObQU\OXR5Q=a95N=OMCc)fJF-4c\aT/KRcO
TVaa+f4F](UY4<>cL:(^?0YTI+A_Oa<a0<PNK<ND<_<+@W/=@0PaGZcS+_3Q]<1O
(V9.Ga4N=/SQ;M;QI=I#^8X3Md/W<L@NW,Q&0VFJ&9ac9_:SH)<,((M1aY<.\+N-
B1UPWIZ.Hb:_cXHOScN6A.HM<fL]G7([F3,aDA4?K]2)J8/,1Z3S(E8e5aH(H9R0
M2Z-B;a\Y<HT;&a]eV>@N]Xa/=5I:dd]2T>SdP9[VS[BHdJQ6<b&5gIg(:g-ASd,
:9/#50)9)>@L5TGc1Y\4?QCL/=4E^K>AWACA@(];>E.\KIBMBd9>D:&5/2#B4PNG
7<,\a,/,:X&&adV&4X.^1g7H8/[ACI@9/UPG@A(Y07RO#M(545^V+gGV9MV>3YZX
.]FO44QGdRL-FPaRF9)ZE.Y]BXA0NJFLbOWI>1F/<8:LRG:R@UXQWRQQC1COJ.4a
+dI-3M<@\E01S&B&NcRVHNB(C]FHHeagb1g-C_c_.8?c)f0>&LeIRcU4(d7(+5@R
&3c.)UP-T<8J6Fc_LW9(1dg.[:[B0[;;eUc8Y#TG]AZ8?Td\VUY2DKWCfE@?[F/.
LNe\W]V+a;XA\J_GROe@I<(4]Wc8G34^V_D;DBZ+:6_bYS5V8-NM:M/ZT@CB]?7T
4&e^PRKZGfI0bd#^U?Y\Pa-[XR(\gR,3[TYSA&7+^R13WZ\T@+UEc>Ob8V>BEEA)
,8G+ebgPW&^Z.D@U\gbcd)8K_1^#,3]@&VB1F<fTOdB=YXYg:OA]V2g&YT7IA@.(
TS_()829K\1M\35]C;+ac0ICJ[S4BOSAIR@a]7]:VfX5P(e8GBQNYN]3SV]_4?=S
0FL^_E&OAZP]9AKCANH37I,)1e-Ua?TFG4L(g-VQ4e#J:E7>e6M9b>.:fVUUT5[Q
0+D@_,A_a)Ge\(?+XCOc6gK8d5\<,WO;\WBAR.e;0M.WJKGC;@WfcMWNW5\=1K>D
ebfZ&Zb>Cc0C^T[4QC?KKV3ccC4Y@KR)(:fGRDeLBJM--f.@Ka^-DPT]8^b3;N#2
T7.I4GBbF_IP?QAG&fGEcH0P^1dD_EbSY\_.UcT0NL2:a@\]aU^8AYZ=8]]17?2?
\ZP&)HXY?UOW:[>aWCf9IRJ)R\FbG8d.+5<e]b(d>VU@Z@6A=+d0(7<Y0M[Qd\X2
_b:&a8cfBZL]8cQ;3H5-ed3f75]5Ffb>VFe>.\0HE=5[]L1Q+.ST(B&FT]MBa<4W
NADNcC+b+[9K1?e&IN7B\MJU.V(fA\f5F+:WBTa<9N\>D+1E;:+^.7)Nc?/.W2e&
a;9;Y?c(eH5FUOXfN(e[4f9\G4-BF-F?fG^8])[c[Z6gBCPW(XSAWJ?5&NGf,L>C
^bCMF_W(a^=G.0AY@?4]<.784D-1^VUIEN9]__YdQ[G<M),2QF=CP,IXY\;TJ.Wc
:R+b;/+H<b[7>MIKgMV7c7K2TV)SNXCKcVU26X/RBQ4Mg5I/T_(M-dLfF0A]8MY=
-V_ggVTVc4-6NTF:9,d>U7](>c#N_H9c(HF.=R3ED\V_d.[,CUd-DdZaZO\8f)<:
ScA]:?5EAKaCBU&DEIJ)K,:+e9Pa)a5;BGcG;Z=>&X\F+?MS<32FNJSdE]I\K;fX
820RIJKGNNFD)P>g(K3<O]2.UKFQR_9=EcH16g7.P?U5:<0L<Sfgc/S-=TF;Sg+G
FcDQ)eNLO=R37^^;,N>ML@K&fPX&U5T6J8F3EOK^0G^G6GMMX6M/44343_6H][U3
D6UJ+>\Z:a1He9;NN59V62EWP>E7<gf.bYK#U&YOMGI7AZRJY4Of6aR^UZYFD=/L
\Q#4O050a-YV=]X:8>fZPZ52M]RAT,BCR4L9JGZ1EF3aFSXf)B]74JE>99QQQ:c[
&.#<P,@<A-fcD:WgKT8\D:=:4AaF+[RTY+K(d/.g7f9A[\Ue1N#-IB^Je>(e\D1U
B,C<3/a5TdbJL5dW6DZS<6>MF4I6Id>f=--DNF45_CBLMZ>0:-HF61)E:=7P6)TV
RaGQKD9MUY/V2JM^2?MPI#3D.OcL2JFAX&O2OY0OF&:\S5CD\U?S+1)FPKN0c8)Y
Nf/U6QP_KcL:A=AVT7)(M_GITKY-I1_#Z)G3:H4MR.65H15M.>/];#(F>]JS#NP<
7ecKaY@LGJKSf<C:2U]Y@>9XbI?6+/,;8gCEB1+L,04X6++UVfJ\F@b)eMd]ENg#
11CM/.ePDTDQAZMRJHa\RY_.Y^:1Lec:F-Jbe,O8W<U-R^-WE[[<C[gY^+?N^2&Y
G14R/U;f_2,4&^+BYfGWM>_@S[MB_H?)2F)FH8+Q?Ag-gKUa\737@\fHcNgXQ9\@
:#Le+e:/cB=QKTa8YQ8FDTRR+.5LP@aLW#Rde(cdQ0_GCL-[710O/c^bY@0PGN-W
NcL,O)&W-dT_8gZcZUS,6CS-bV[ZQRMdV.7M]\Q_[GZ\5P/>KVZgSMCUI]Uebc>\
/X)fR[91N5B2@HgQ=L)7V4XHD6AN.<Dc?+^[TD@gAE0ZgVN+Q:4d)0&Yg,&R7HOX
HCN-[4.3fQKRM.cC3c+c75-dW<ZWK4KO3aY@>^0CQ6^?C<b>_/C&^BQ?<F0;@H9R
B8(MDS0)dd?^O=aAFPMgQ)A42g:XK-bESK^ZWL/f2YCB6RYEMPRI#W>.S7F,#O,-
AI:gc=4^[SF-VFFeAMHGIa.D,?XA,QW&d+,@@,:RKO(SfSAcc_/P\;De@4Bb9U?D
PDHBXU)RNe=KOELC=-b7^8^fZ+#<VPFMb-a0)/0,+5@F#a6DY_-bDAIWD_eDaYJ:
5,(b5O2UG#OQNGX<KH&O8Y--NRKPX]F^&LQ6C6g>5SDZc[T[A.aQCP,_3M.R_YAR
=/63Se+1D73;c/:Qb+FEH11]DJL(c#KaJE3U4->9L<C#S&2Y\0J0W#If&^<Y+C&e
M_J_.+02FI2NQ1<NCPGC]A0IJX)6fASEO539[-FW&OZ+2C3De)Y^]KTY((/C8a(&
aNDPaSB@?/,;f?K-\:5//=9b?>N3CXTBWI065KW99f(VQW@>B_Q[J.X.Ab#T\OSQ
Cf\<.,a+UgRZ3=A3X:UW63dKVA573L_3@3M:,e:;egcMd<SOP7KMe))G45E>A&&0
<[JdA4>R6#XccG)#7^,]O4VK)?[W\@Ra45GQ6b?ePUP\2+N1AO.Y#3WVgI@@O+EF
U6+>P4M-E^?,T1KTF;WSG-48b7)<fcWZ+)7\.EYA3@[24A2E_-f&6@;U04N^M=DR
VAKF6;FcbZKR;Q<U;&CB]R[HILNV??d5f?TdTKD2\a^]e6BU@UMC=W_UE.:&I\KT
:Y.f9#6Y]>5VEGHRa#cfXFAdIELd>J,.c8<==+8CFf3e-C&5W@b2<:eD5_PD-Pf=
WId1@8Zbf;cV^LI\N0VEASJSYdfT0,V)/WAdYRa-ZX_b8JNH4c@g9,WYW9]V)SY^
gb7E2^=N01_?b_F2Z@&Gb8[(40Ca(4aF?-H(6_LdTe:^H?YT/dK/CPUGWDPXW2g&
5R:/2JRAXA>ZgeIC;S@3MGE:KUYOJ\FES>LK_1GLDgCX0LH(E/5.7GfH(AW(eG/5
ZSHGO::<0PQ97?=^FdPO>c>T]);_L@RX1HN253BU_B;NND8-AVP_\cY<JO>Ogcd.
XBZMY2IWR=d6O72QgaQ6R(Z)\OF3_E_?T[N]eJ+:4PJ^^16,D>?Z866H9YGC--ND
(U>DXfcU]2<FN=@#R/N@624f.6@)BX\]CCW<:HFC;?<dHTS]X,egdNVgLV2M62<<
OcReQaCcRD[?JQ=F5a=L@#;8]U\V=6XIR#U3PH]#,8]f9__[\\3WD;Y/#R\Z#[]M
96YT6fHP\<=X[a3>F?;E,DA.CF:Eb26EYLbNaUJL4XX)\NMY0X5GQ+/Q4d&51:-=
N,AM^d<VUFM0G,40+O0Hbb31?&4&_1I-aQD\RN31YL9XDJI1):d3578B0(Z:YJZZ
RcDG;gS=YSe@D,VZ##5d.IFA92[NH;#USdKNc^c\J\B@]TU[U1DFTH<cF6?^ec4=
F:HgEB/D4FY/gfPcbI_.\W\@\\MC7SLbVMM&]3?>)I5[=1Qf4.:OdIC]T161M8P>
X^FBK<bGZLdP.QY338ASKaAHR5EX\8Ib-fO]8B5Q(=9<<1e1S-Y_VcT^3NVL[2#U
S;/)3LbA(I7509HN6+c(9@4NQM_U9(L74/]EbJeILN26KJO-f_J8d7Q4MGcV;&_Q
K9f+N1;F#95G2?&G(75#8FgXW15(,BHU06^D_JFPSaf(69S?=TIL.b_@1I]a.Q<0
aaLP_A0;@<dQcE:S0P4WVZ?T;O/(Y5I5\Z&a,5OfQ.1852G;^F@LKGGMO2+L?bb>
=U)a8S9]/6GSC\Zd/bR9+ARW.#Zc7YN=?[RdUWd<YP)af6<2H0,Z_(6F7-eB<:Q/
Y;:4#/\?MYEM2V>bFM@VSVNPA4RUc9AF=.[:FR59&RA<OX+V_U9E#PS&SIOHG6gG
K)TE;K8AM1:LS]LbY:@ZgZZOB(EeQX(;D<S,5e3E1cbE-(/:+C).CWC^F&;;^5<<
O/B8O@+)D_3g857NB^;&(:,9+3Q#I^JP&2KaeLO74D_KGX4@]K+QaP_V5b<N5[I-
e^@J?Y7TNXK:I5CYK;7<)C:K89S6Q[F>RdONUfCgWMTK;^bR\)eF8E(P17CK;Se?
CE#Uf)Re(<Z#e2LDQ8X8E\2VE^?&N1f,@?D;)\@c\EQ8J/dZSB&]>Kg(;OK^>R26
-/?>4fG)g-X5SbR)P2K;:/Q)HXM5dSCM6<0[VeZW5NL.Q9[E,A[aTYQ@O5e;DY)\
6VA5#IXEO.f4X9.];J17,X;\c.c1IZ4&UQA2&(_IG;0A^UP)8H2DLdLS_G0e_\aT
#)&]0F0S;QVZMZeFWgBd,#/:?TZa_fCN[&?6I@N/?<6+B8W.([C:#TaVG.fHg13S
gegX2=A?b#L7bdY@3,N&VKK3)-+RV=95F9.W7>K?Xg45,>0L3\4@644@gZ9W2C5O
?8=Y@CE]BMJZV[VeJV8G_@fce?aSUdNQ-ZaR&H]+@dR(WD=-2&^;8MYXcW1[EITa
.Ma\(JWI-E+3a/0C#T3O0/0&WU&QHANQ=G[S[GN5Y>_=a-+R.ZOTGcHD<ZKGV,I^
U@,4-LD1fMV1[3aX)H5a_;JCETCUN(HbK#2G#Xefb>B^0AUQ9c:S1C57e+H8YN.;
_MfO:PVLD_U=0:_P(65@I+gF@O]WJX+9[.UPYQ]^1+\@+L^8cT:U26?]J6J/:]?7
fGRHSf^1-:?fH(2TeH,<<DQKP?WdFEb5M@D6<6g2][[>4=,(daQZ^aUSMT@.TN11
XQ=;YOOA#d)F\]/bXU/435BDa1cGE),7H(RN@Y9R9@:4U-CdW?9g9M)D)APMJ:/I
A7YBE-E?-3_R@09W=;<?Q0AC7_JeJBW^af0;)OHS\^JgNYf8#@DA^bOI)&9M^bVI
G6T5]5R(&C^)&7(0^BPT^<[;gR9D+&EG_ZW<RSIXB8F=C3eKITKgEB8OObSULBA=
UV4Q^8WK-[f03cYd+Xe>1I[MB0MXNUg&EU/5<>:1Wd1V[O+MT53P@J/AO1_3]d.,
@L9^GX.);BT-;B65_U:8d@.8>-&b(8>1F31U4>\CQ]8Y03aUN#@.e<C-T<3g^87[
fH(5(?X6d7<+II[_S-g\PS9KQRF>0cRURWK@]WHRTNWUAZ@\)^Q^-MOZTfTF^S+-
OaB@;RJ/=Q7I;-@ILY]LcefCFb[ZagRWQ[LD2\]C2IL>.]5M3@]OYPS^O\g@@/-1
H]M#gaOOF<4&NSN1<ZfU7bDM=4TH:()_Kb_RHZ]f/TP&2X+FgG7g=_Q17L());d^
U&?bUZaZaT(]8[6#<,U84_6(_J^.e3aJc&L6ZZ)YP]\8Sf+8a40D\5=U@d5+182/
BVa-LNJR<IOdSZ^Uf#9@ZS^]EV)ST?Uf_Sf96XIfEW[)Z)41:+PTHO@PETBa_4gN
WF,:-]L<O@:_+-/cL4Q_+OP+86Zgc)\TKQ@L]XMZ7.K>[.JQf2K7G>OKPSHM5fD,
7VGdfD5#d9:E\ZJCX7OM3\/TX,(c.fXK9eNJ_4TQ=@SJHGffe@P3\\7[QKeF(4V,
R.ZQd#R?D]8ZNS[a:]MWP8K<A)/T:FS7NBR9\I]4UYIF@+0\<IK3d4ZVSW#=M1VL
V\+YJKM,QPa;KP3GQ\_)V?#VeZWVUDa_&:&DNQagE8?eQ5Z3N+4dV:0VW@8e:__&
=M4?cA[I4^D,Z-Bf_D?UH-Ce5BNWWDYHF)fZ4#R-2Z^F>P,4c)DgLI6N)M#]3e5M
+.>J-4VLFS48Y@e_fcV=\QXPAgRBAHM#Y>T?97;6:6-b#HKUHGFU=]F6B^B.8MHS
>d--CFB+(O:?)^QE\Y[GWN]>4FbXMC(L,1L6ZDc-f//,7]>ZVS>-XdF79YcIc@R1
6e..NQeP_Y]N6>^/X1:GI7>b8H(>@a;VYLJ6U.<W1>DeZNNg6)a#BbXRQP)Cd:GT
X.(EQ?LJ.:288&&VEA#BAC-9X5G7LZWH:CHSKH]K)A#6-_X;/:cgGM)dKM;)LC2Z
6?Y@6H3gC0Y.)gbd[G>f<>@EI(\#7KAb)aBW4];f?gY9OL&fa0I3A/4^43+(&?P?
5)1Z#QSJU(PE156)NAYP(FG=^d15\7;:IEV9;gGAJ6,Y<4E;,FePD@a\@LOCD&[4
4Cbea&URAaE]_5ZD.4Y62OYA1HWIO9>LTB^MSfX/A_AcP=U^0(e\)cgRJ221(S?4
cF7\6O8Z\>+WeKQda7&)50J7=f=\\5bYF7_4TLUeCOHLH(_^V0G-4@E\gI.+@^\a
X5U\7KF-4K165INdF53.f9]8FHT?^DdM[=UAcWC1)<BN]TeBB\_M>L(-#.;)FMVS
7UcJNF^?3497fN^N#-cP9S]c+E;1O9T=1)M=E=:1I2a]STZZY1/@[.Q:Ie?K9;Q)
MQN8(?D]P=\Af?d[+?C>[9CfH4B^_7;7A#?IY_BWS.BP90bG[-E9)35HW/P^;LNR
Nd(.da4E0<F0I&Zb(C8V-b8<\)OGO?]KA=[M/(WBEN_P]bT9LPP^55bUOg-KS7<R
&@gR>d]+8NY+O<FQ\>A3?CTQ@@&X2XXDY\68IXPNRefE53f\4C,+M;TGd5^_-g:?
&d)[?YMOJgW_6G=-)M+(RQeA\BP2_,.G\/ROO;D+DS#V(^Gcg2DBSXY[eDX_PdJD
,T[,PdQC,?/S+06(8^>09#03e>#M5=]ZGcTIA2JM9>8@c0DCK+/a18/gG&FG>_(9
(5]K[A<AJA2A8#3XPB+Z@/1.+8gY=X2ISIGB=SNb2^Z@O)T7baa=_=0\3)KJA38]
^e.>LNL@_F:/S1@BDNVaWZY5FEZLgca-:_K\B:4QN\LUB[00(VfAS(&f]V/#_G/9
8,C#>F<VY656,bHP=HOI=HL6SA7E03aMW;(Y_Ga6&)3>VBAgY7DC==\,9:(TWQe(
1,ND^#<EDW_b;fUgR9UVdK#5:F>>)2aJ5M3OFa(XSS?G(I)eO--O=)52/aXX[3W]
;2Bc.X5PbKS+-#NEL[Q+\W[6>#a&93Y8/&T&4eb;3DGJfM7PIb^Y66J60=g0#<A@
8cL.C32SJ/[X51ZZPVJ2J(N/5RL2C3:>P[4:8EYb=,HLRF:??-A0cNQe_N4OE;1T
E/XDFH3W@4F&LCRVM9cdcb.4OC]9DaB(NT(TSQM9bPWTN,ZH07S5FR+]c9OLT/1M
9G>1@bLF\BULFeFgLMY,JXOBI4EQT/O7dJQ2P1YQD:]&6fZKK&^(c[_AC+]HUb?B
4b2:E(aEW6Q5?+0BKd#C-#^FM+Z<^E>IJZ/]LB3]Xa+PG^_/b^E8@8.@);/HY_3H
<]Ja=7E-EF19@IB9fDWJE(>9OR9&Y4NaPeWc;(fcd22?5AB-T?;LcfT]]g^X.E6Q
[;.C2Z:]cH94BLP0D6K\RDdd<KQ-Ja.,A6.P^C@90H1dS2;f>cK-YK[N=O@L4@;6
Y\5#eVT#25e^6;Q#6(dggTO5b2)\.@Ldda2gQE7&++.6:[9KJ4N+MfA;6Va^5N\A
PRfC(T)(:HK80)W:[TE97KB<+M6MDC)33S8.\S1V#2GX&_/_]R@KSU1d@DI;D6^&
6XOWSW18B]S2b^HL\6U:>9BX/b)A=K&OY6]W\f/c<2>eMP66R5ZAS43:5O<D/?OP
f<PLfS)g[##&b5EeL[DG<EB]AHI_+DG3VO:)@48VJ40D5a+^gO5T5MU8Z7)aJaTK
(XZ<?9.Q5Y;XADXJ0=)/6/>4RON&O>OL4ZKK#,@ILg<gOEM6PG.gN)V>.2IN(N-C
eJd9SNVDQHSV/<GGB#,XZL^&fbdYOHI;/T.GD;RFL6a:c;II6/<V0b>^DRAQ_02&
6UT0?bgI7)eOGHg6=AO7A5>Pe4aCSU6#OK>e<LY:O[Z_M4:6c_LOFg)<7BQI)L=V
=HZ<?UZTW<-fK,=AO9#?KNJEA4?Kd81^GOC,g=_\Xd1<Q0KdXY5-XW56ecGT+Cf2
)D9fX7(43W\O#B?BK,X97+@T_N0I<[IgQ9;//(d)531P0e7@?P@VfUBI[(d,L>[W
RgXU-367#/f15Y0>=5/X;6VdLNGE?F^C\3aTYZ9gfP2ASI\WggXM@<T5C>O2EDH\
GFC9549X,A+INff+YOOA]]H@,+TQJ0A=6Q0Y<?M]DJJ;/cZT[KW?G_;ASDC]^OB(
:UHc=.9TZ[&<)6Ac_f\.6<-Y^#0Z;,XS(0+EeQ#@HNd<dWX;V6_4)OH[FB+[ITH]
:EZ1Sa[eSC9(D2SNH6Z<[0&4L2e]DaF9QB,Y9><@0TFUEYc3TZ6M_^H,fS\1ET(@
dcTcAY.^3;T2CR,5=&3QCE7167E,\V\baJ:+,L9^MHVM@(C4_OcOcW1C3Rf<5JY0
D#.PbD6&363Rf-B2V9HV;AK0b>H#^D==>+2IH&,d6FD)60.IL2X:XQC/#YE_91RG
#0U:]:MSeYdJ/ZHVQ/G\SPUe5Vg,?OB/bW:>Z/D92=a.T9>>#5d2Fb1V,]8Ia9?B
3_/3E2ULVOVY:O-5-\^d-0Zb^g)-6@eQT>;I3IUUB;(]fG9\[NcQ+<J8@7K5X[BH
X,R:AgD<;Db)ELgV-YYD4cL0.QV&B(#Qg=3d\b3a\L.56[788RdXD6PXJ)TDcW1I
)M^aN7Z5#(A:V,.6\-9NLI/I)VYg+CDW:Md1G<cFP3d>bbb.SS&(KAMeH@S)&^R0
a.-bK.<])V#F/>BM[MZe<=XB,E@dYAccR193L3,,Z/Q.+HFKH=cMX_L1e<5N<2\I
X=[->b1B;8QMgI^E/JR9\5>-@OZ3.+,)YBaYP:R/V:5\D_H2(ISIZO&Gc9(20dVN
)Hd0BF,-(aceDYFX1/5aLTF-1?B/f(@?fCEQ+:D+KLeZ7d2dIXOW)f4R/+,]^]5W
_E84[6f69:0RNRSD,.30aI8Z?If<+^d5e<9^RRSH),eM8,??>R[b&80eXN5IF7.N
552;OH,_OB/Y_L0ZQD1<;&f63:3]I]d/N2D.Q<b:=GTP)M)HC3F?2(C@B?b;.G(X
?1W&afM^V/Z()]YZS;UK-]66X9aY9FV:<RL5>aQ)2#Kbb;^d5VS7ER6,E=a@Ga=D
29f\C5[.91RA1B7+fQTI/0,.?bG-.F@24:7ZEG^+S(DX:-L)_]:)P[SWAZK??[-_
A/>UO?U&Jb\DA&A3c8ETSK]>E_fNJ)_V?aJ>+ea@FcMOJ9XPAfO43GYZbA^TEA8f
^cOQ_PdXMF=Db3c@/8g;95-&O3OXWGW5LDV=#7R;-?[/d6.aJC(0.dLHG+\:AQ.T
03JI/-Q]8WDaEC?a;QJ4ZfQR]A#>BSFPE7(P=--.9#.DP/6#g<WYF5ML>db8BR-N
?0RK4^aZ;.<:Wf4+cf.d,1Z=Aa.6:]?27Jg^Y4VKKBSC6-(E)Z-LP/&91:=HQF\<
I+FC;F^RG49fggPdW;9EIZA1GX_0^86N@:_X&B52-M.Pa;MGAO2Z??Q5NGU.cb2U
LfTaVV2e?B]\cE(A=:.PgC23?K-/B,EV;Z\E81:@>Z;1^W8ZU]TS)d(;+\Id_1ZN
VD[.;6[3]6c(H:9AQcQdf.K]F(YL=H69J0@EDLA.5Wbb?X.O1ONIc&<CX\QeCT<W
K0ON/beH&;/P?BUE\E6aXXA9HMP+/b66(,7AVgR,bO,Q;YNb2Ff)YVCaY0[>WWPV
3UA_9Q&Je7A\N:-4K-29GP5:Tc7@CII+g=WE7S5,9BYQN[]IS>W50KF5L:U2aaUL
WRY>RF(f-C..GN+X2cC)L;@3[8R#,2d8]1H4^+LA-1WX0Gd4g9Aaf?2::S(A>\SN
eSORDSW1W7g>_@\W3#0X]Y#eT7&NYY&?2(L<719La&B3>UOWWV7cc1[V6]._N,@>
]E;P6:J#B1MUE2QIF(I0=TI6\GfPf1<@8WEJRAc?X6>O)NXSR4@D6F\:Jd3LV<=\
a>#,T?_+e]OX^JeJ?207_<K(AYT&=U/e8K>WN20f]:QN9fJ:825dM_/YWSKTDHJ3
aP^gGCN7?\g7A])07:2=@JLQ/VY30=Pb#bW),0.ZP4KJa>;bN3/a]NaeAR&Y-]]+
\Y3R07Z9F;(1L,UME3IS6IE[8eC7#Y]/c+Tg)c(>=Ve+]J#D1/KA^8-(J4-P6Ae6
4Ce;TG>^[I@eC1=J3/F6+_I]b2X<H:<gaRC?<Z4]Fd/N49RVgUgKZ@-SSca:+R:e
#3U0X,1\T1[Yf):Kf[/)f)Ye;:)7E5FIJEIZL-S4079A,;&<.+ca,?,:=5P7\DFX
<6:RH;FLXP8P4Z_65;WH&G1+31e.+a:b7GHY=c=D;BNQ.gLC6^>6:^f+Vg9ef5.K
Q;AERB=>1+9B^b?BYYKR,_\H4,[II_ggNc_f7DE&9N9PUOe:BW<;BMd-SQR3=G92
(FB,<M9.Q3KeKcBC9XN?8<f4BL.49M&9FD+Y1)L^ec&S(LKXE9X-/IA)Ff;3e41<
?;I6ME>9@ODGC[R9a5GR2=+MT9W7U+@TaU1c(4J@^0YbRDD7Y6MJ2Y?M/?;(.2Z8
XR6P^X-Lf,YDFR7+c6BaE^:Cc,E4^Tea4,I1ZAT+/?1L&??=V&ZLH9.#W2)QH0F@
0aef(Pf^)35)A[PY;=CN3>27B7DT3[/9ZF=)7L\.1(4#0c?@6(I&/6_YF&_J[3eR
;\Xd1V6ObFWObS=I3/D9.:f>N@&;LCQ<\&[8Q(8GBcYQfJ9U\-F7/#?EIXd:A?gY
be)Mf0]#(4,08=X4(8.L.ED2.2L#VY?)2+NXD9MP@f1J^#O?<W,ME8(]8@6&cU=+
<a)UX?C+e&g+b#a>-&Tb]+,eUE+e_V]V]T&3aM)<5,5.+\R[+aaO_TeY[U->;a/I
?cLFgKY7LK@93X\T^HV8d(PA^_81a]Y_8D-PEa?2B:8@4KT0A9>Hdg3?a=f8)WKJ
K3QRc/Ef?b4(GDaW,Q@9eGD,-aG3470;,LF<<>5^F0Vc/-<.3ROFY]:67(;b<@dG
geG5?cKZ5(CQ&Z@?5aG8\/_CZ9S_:XMbD0cRc.1[F1^5GD^A)dc;V9O;B4eLJ,1D
\WMP_Qb<AeDZJO8@&=_P91P=GZA2B?FRCC,##e:?P=VJ&]1GScAL&S,]L<D=<E[/
cb>>)aVAPO,Kb89(9ODYI4)63JDJ/8G?N7cf[UJ_O=\].cYaS33(&:I>,deY)J&Q
6&,,44fY1J<F@#EES+,<^1/\3U:Ia+=?&P#QWL,-7.)@K??ZYGP0]#F.^:^HU4>g
&HL>I1?)6U)L82Y4J])G=a5ESHZR@\D?aWT2V@?Pc>0P&6M5Ab&G.<&8e@W#dYEZ
cO@]MOX3_FD(SCR-N0YU>&K)f.c+B0-=^T(2gP>e=O7d6_Y(]6V]Z76>9(R/<][H
[^OaXM5S4UIK3MgYM>>;BQ2FZOQL].[H^DC2JSV@25_&N1Rf1LaAY:e,FQMLFRZ+
1;^-S0[A<<ES:4R?Nf>5LDMK&fa/e5WZLHa8RO_.JW/M\@(I1[Wc6UU\cG9X?f-M
I,.<]?Z6IWBTcZ[.SFb,5P97SL=:dcBT3PJ7I-^5b2W]67O[E.MAdA58BB[#B=_0
BWW]/_49?-d2d?UN:B^:0OQ(4D4&8JU8.gA=:gOFWfV++R,(,0?8XKUeC1/[Y,F#
F>6K=Ae:&E52XKX&)&75(CR17<RSK^<g#2);7:/GAHNgZIc0X&2UBS/<d7gH0PgH
.?.6:0YP]X6g0N]8476I5;X>aOFU=:8c:<BP/,+B;,Bc@@;N3=Z,S9UeJ=FL.Z=f
B5c5b[PU,TACJBB49,2=>@LSNdNLcDWOK,]([HWZ=3B,GeYDI=?\F)7AZLIRBNXb
dR-,cL,8,b[5-LEIfXW5Q9)LK,-,;dB.;ZQ[RT&ZFcNHGfVR@X8cTVMH?UC-.1WJ
&5]0+]PN>T_Q_2:Ia^SUBO2/^fLTFZ=(P/85&U]g/MGCA]R5&d2aPELAQD3B#&6?
?BTFfb\9>[Mf^D8LD)N:,O-<;=EFO,1@HF6^T=[L8^1a0X[7-)GP#JM];>HY.PE:
^.KG;;eL,QFHVTgL#C>Q(F?QP9]X;3<@?ZdR>KW4[HL;IDf[6.A.R?96+L5USXLc
Z7\[(JKOTU2MA\E>7L;G,BBdBO&:H;G(DZd7g0/c.;+c7bEO16=5TM5Z&:eIeJN:
P;&JF]W-ZcRFDX5]M.YC/L]aFJ<ERGMJc.TPD_eCIc];KdM^=Ug^dI<X&KK?C\3U
Q+RL@)ce@ZJ&^G(f6gY#,20C=GL0C3++;@,+eN&b+CO,EPF:MW2B:[F57@6g5CG3
Z6aST/HXJbH)SeQL@&^9TLg#R5dPfTE;@4[998Z:Z3gFK3URNaYAbbUe5A,G+_5+
+D8R_ZXFYQ0D,R:PI9;@V?#Z(25#+eDH(@.bH09S-Q@.[f.;ZH#D]S5SKE^)1J@G
+5Q=@[=(U)-/LZB]eI1De=C/cgdKXE.+VBaMcM^:b@69P,D.+5(YKC)<J#RdHJH=
A#SJ\3SBeOW^edg#)W#456e:C89Y;e^/,/<QUH]7(\@f+9-?W\/A&Q5>._(&3+W.
d>9^#B:L>=A4gMQAI58E<(73^^UD_9@G-#=:>7U8WO21.8Lgdc\2S3S7DDAd-EYQ
I</YgJe+2A_[(?/X:c1B6X3ES;cP^X7=(IgF=>g\\e1X=158dd(98F9g@2/?+.6H
5?S4@#f9C;?g8I-Ja]=E6:8d6I97;d^#MU\F)X0Q;Oc87N<?CKP_RV_CY+<OG//E
>OAH(<&_D:gYZ@VR][a#?-8L:fZJJIIHC6G83SHP:V0F/?:KNU]=a148KBYS[,IC
R?J+T,51L):4.<1d<U/+XaAR2,Q=DI1(^2R+5,HAD?<-H[<T>S/f,#eZW(LG#GZN
4G2_Fb>Jb?^GO(f\e7g@TR>[6]XdOKaR,a08S/IIa]>C\<UU[)fZRH-<0&UJZM5K
1>Q<Y2I3682>8WPV6DNd^cCEDfRTO/V@_HUdfKdQUJ;RfNGKb(<bO4IHDeC7]_@Y
0=NCB_]487fW7\f=5_D?YAaXaQNQROMFP:7U_g-Q8JQ=KRgT2X.NV(:=?WYT6Ed]
&N<[2:Yf9E9#=d41,SbZJg(B0@aOE=IN,<H1K?V^,^LKHM118:1aebYbM@aCZ7DO
a+5Y3g^_1@HRD=-WcY.PdX\HHXeD\6(I(Pe=:0[Vd&3@;7NLdHBBJI_c.<;82NE6
4H.E?7&Q\XFeFFD7JK86b\U]GR+.CYLb?GP9f662H-:;I=0A,T,3=_[C@R6eUX/a
V#M0PFBV>@_]C)S(E=Rg[L\.e-+G9?9KGRW=c7c:fbR3OcDMJE5I2=a7bQLc:G#:
;V7+V&4#3MLKBZ1(>2f0A-bFFEfGKbHAb:a_g/\+F9(cQ:962^ZQR6\Z;/OPY5MM
+^R3AfE]>N#?2LEMP,^O=D7>2cdFC^(#@,R4SEcE^1(EJH;XTIe<U@GdXcLbVRJO
1O#L#NcTLO6KB(HR(Q3[Xc]D]K4#1:Y34?X(#A4V=3dHQ4aU68/M5F/_YG7Rg8JS
D6DG]c2,\?@IQ;N:/J3VfV0G(69(IGG0TZdOND]1-(&:4L24Q-[C;.M6I9D4VZL:
_TcV?37M#UKYHB@IU[ab(?D8ZK99CT9YG<+HN+YE8^.f.BM=b9Td;?P/:B7:X_KK
=7Sc[QY4:9.GIOga^2M&-cUC2]C5^&I&gcegE<TS)IRX;CO(Mb-6UOJ>a(bYSe5=
L\8LE^?K6Q[0gBP,fC&HYHgC+_6FdHVcFbb^,6ML7_45=5g9@4g<AV+#dM\2C/BP
L/:gKRSK0a(-b)SfZKP/_2PPUS2bV?g4>UD?-(([)BL19P8W_f:[XD[gOgE-YaDe
#OE::c,JHR,e:d[+P[2LF:JCAeX9TadI@HTg[A@4Y(d^?M&[S?>R)Y>Q51F<9GK;
:MBJCbBX#d]CIO=0-/187>(5QP50JNYSIOcEJb&EF#L4Q6)6;^Y=C-a]9NVV-J6d
U8,OIXg>XL><:>(>#DX9AT+NgMXa0;+/3DPHg+)SeXBdHQAA0:..;FK\:C,_#&b_
f2UfG,cDMSW06<-)W6WK(4J.#)Dfa=[KcDI2ZF#,EM#:XY#>U)B0:&8UEgP;cR<0
4R85O4ZQcAV7\)DJSDN7//,M+L9A,aM@8MQ<D9BI=65K:#+5;5))XD72=H1TC9OA
8Id<PZRJa>5.DW7f(L8fUOdM)/_CHYOARK6]0Z^N?,dc^UM-f_:LDC^B3Ze-<YW6
8>9@5c:T^e)X17&#BB:XdJAZ#H-8/c#7EHOZa(+SHVI_V7ebc9XePD&)Z?dN)4#8
<HFfPY81^D(746YRP9FFN_E_1HH4UMSc\_E]K2_>EU2.N=I]F7^><HX5VB9YcDXb
U\R3/E4A=Y(2a.7+^]DVIA7L2I15c@7,[MZHWWP6(?R[cM,,:gY]O<,K/&[T9,71
1R^eZ>-R.Md(e6\Q5g/=1TS-Q5SX(4N97fJ>U7V&A>.?X\&,cf9(J)-17e-C;.<&
WSE]&B,ggfd6L7UOD_+(gbMA:dc[O.71#fFR;?:UeM<<5\Z]8/#6TY^\P<g]U+NK
0?<A\bDWE@T3ON4Y@7[2T]Gb\[e@ORU.NK)UFA\;=A9+BL72+@5Y8C/FdEC],bH;
>W_[_FSG5Y6;=?CNg=;cL?ffIf3WSdY+C=1+[XGB&D3IN;^)15+b6QIW:VH,a;NB
:0e1>MZ\;J-DY](R7C[=P&G<G+K.6)7K?L:@H>2O0c@30\@E]_A:LC.#TBNV/,PY
=\_9G5M6F-O3D@Ka_P<=+7..-(Y7=97J4c0g0Q>NEIY4X8MKIMbB9H\-.c&#[=.Q
Ra:(c>WS@I<K?bB-)8IJ7RQaEbW+()Ee<Q2=6.CC<@UY]AB79:2EfGK\2d]/N<@B
J&--/@XSEFU:ZfGO:XPF:0_L.ZD55#RdEXED?NcgN9c5>5?89-Q4H(]aSR/R07ZC
#^5XKdOG,Gd+LI73V>d;[4bXV1?=E#_gUAHg\3)93&;),&NDBH_(</9W:V6GZ[Ob
0_\&;EEHa4e9WE_7079M3/F_b_4;UHf8BEDb&XV3[XZ8+-Q?>/A^:2;dDeIa4EB-
^C8&OS(+^<CZ?/)^eYW>8>X2I7BVJ+LN:DNgML>^EE&^2e:A-9UV6I>8245+)e(F
g_\_eYY06L3-L(f-bVYeBgZ-9G#cQ#7RfP#c,3IN^N#8b0.6/>,7<e)Da9Q2+b,R
?8+-dTBO_3AAYd.YZVQ2O]4aHE<;(Q6;2,#+Y5]L=ES(FK-E;V734?TSO7TJEG7:
]24;T\,>EOP?Z18P4UaP/IE7B(E\IeRXU/,.<8S+L9YURE:5V@=gMMG?YZDT2+gB
fVFS5OM-#0]O0V9X@Y;J6<D@IeJBTP.Q9O9Cd&LTM\&O[:A]YR3.491^(XbfWTc[
bT+)[G;IS7\I;7S&e9SS504=9aCIIJ?,L.&5CBF>eP]TH&7:da#bF2D>1d+G9F^2
FMY\T[7U=[\M;#46Q(<^^HMM-@WGc8NWDeX8<-JHb956D]<8LXN2Uc[^5IT2VWU5
VE[aN#Q;G:2acXafRTA:J61RG_3Uc-WadJOH@QI2M9H+Da=>6ADQe(QcTJ+dH.].
Ra;2.)a\FTQJ#FdAdIXTXUHeUO>QfY_Z/a)F4[BLN=9&SY2TFQFDDBFH8D+]2(H#
KZB]a95H@P1B(2RZa=VK(cH^H,(C4^Q(5\U^8&T_)4X/4@ZG#ZI&>CQe](ITV=Ga
:;d)?0]O_b>ODU9ZBU.X@_a]S6\;YdL5f>36-?Fa&49IF.]LTARE<)U,9=,dC?)/
Q:U[E?D\49[>K+ead]7dJW@/S=16<^a,\MGY1e&<3K1\O9W9dS>cG9Z?)1XeM2BK
2H&fKW/^UVZK>E<J)8?f[V,>R>Sb^g\/bR]:02)aU,PUbEL8Y3?M-CU7Z4.Y^7_V
-O(ZQ4+BGfK0=?F\S>J=X=\V+#@H7=+RPTTN3.6:R)LIb(5VQY7,8L/HA.O?XgQ7
cUS+a)M:LA0)A84^RATYMUIdaN7[?a(]IgBZOP:Z(LcP4_C+PWV:5R-Q90=0C:Ra
b,/U1CO>IJfc:0)Z#OMd^=ZC:eE7Ef#?58_BQ>8EbGJ=QY3NT3DdGID@PF(.3LL)
OJ=YAQK&U4GGBZG66WGPLX[E:8g\C#WH@<KY)]J0EUTcL)bK)T-22CFEV.1]T:J_
M7<)fKJ:@H6W8W):7[IRefJC0M93Pg9;Je4,&R5C6X51Y)b]P;JT4Fa1GN9\W__7
f:LP9]d):02[MIdT.AKMU4RTP4:EWQG];@J4Lg/WZ^e.1-S0BYA32-O)AaZ9_=I0
e?RW#_dZ]eOgO#0WB]K_e/K62>6EDa,)D[RT\d8FW<[\d5+_-<+5Aff^bL@aNI/&
a-+dWSR9SbLdI9G@_d&GV4\]Me.4(@_DV7+g5<N=3ZWH^6R50JU^3d),2D)Y0Z9]
ed,#4A(Z^HASYR3L(K/<5X9D\R\WH,ga+SRC[E>M_Q(eDPDCGU\&EG?N8X\_Y9-.
/].;F0UP3_C.Kb0fB#X+1>3=-1W3Y01D9>d=,_.;HS3<9==C>FaId2b50=2]b]>A
0>&W@BB-U]UU]>3(=)dB(@cf^Tca87<Q6^5+,2]/dd#(d#gR3cL\??;^/5\36W^.
>:Bef0G,WP:R/8KBE7QU);T-b3SMI,E:RR@R3E]U-D-a6+eT.)8WYEb>#.4(LD@:
.OD&3W?EKP4gA@<:@TRVEFcD:@O33Ud:6RdV^Z@37I0@-JFEN]:@_/?SS)NN\(]>
[D]d_<7Z(N3<O#R]:C^2)6?P5Hcd28]#)1-LTXf(dQ=,QQW^7Sc()6:+VgU#1L:R
R6RLNg73D.-c=<+1bU9?IWeKMXJ[+#MH72&63,)6,6>a<>B..BUMAbSTf]]8K#97
<S//=+?N^:/#a:P#]M_TRFE\(QVOR?:[g3@@P8-V3V6#:8,YY[a:3,I[aDD5).C_
GLCXPR7XQaB+7H9bD[H1W/F5ZX7.H9&\3=?]1=3[/8(>)GYJLSK4(7\K=Sc:<@R(
TO)f9T]/@ddZaFL\0DgfE>FH+J@f-/_f[d65E:Kf/1^6-UIdG4Y;LR)e[H<,?294
8E^NMG3#RQ7>Q[Z)6S-eC&0SGDLVS_PQEE??Y>T(YS&_A/?OaABKU16f0/>I6M-d
ZL0O5,&29/JREBRb:e2A7#(PI52&(R>Pf>MQMLc8B9LJY[0.>Ya7:GN\)#]NQ:D>
c\M#DU^8G.dXK\fX@:&Q:;d7HSVU-^NFg/D0HD--U&N8+W,</7V1E:^g<KEM1<&]
^S-.LUZXOf54W\ePPfZP\&Yf0Q^?NL6+)M/0_QTd8(,-N,)gR^:Jc688,A7MgMXX
N;7/<3.-e,.CA<\7LJWeL:0RF1=1;0b[,Y_3W^fE]LBd@KM2Q43^f;&M9AH?O<aF
^ZC>>>#7^4:GD@64UM7Y/O?14B1=DAJb25fI^0.BA2TC2I3Z9BGV0HKK_,A/dKB9
.Q;2H7K=HR=K6E9H3SAI-N\<fJ^4G=L.YFIG@a@f9dR8?.X0HNPLLd/CdW\3ZLJ;
5GGY6L,SE5a)FK9^ee[_H45XW3EC@K+W&:)>VT-_A/=(N7(Zcd[g<b5OMY_&Q#4D
L-O-78WOg&UZ1)BAFBb^PcRge#FQ_f+a,9RF9[<WDK[-O4FOeLM<>Y:/H#3YbJ>3
=X=;BLXg=D_P>e8\BSFSN&A=-e/SNGa>gC5T,HbT<+DGAJDW6Cf-;^3Q.S/Jc)+<
[ZLX:DW>&@45-=fMA&(,G5:O0MM><V,EI,:?\_L5&H1<_JCW23>Z]@0[;F_1WMfB
F:GI+V@\-D4Ob^=WWUSVCU2_TDgPGO9HTfF.5eFfVEeg#D<S)NV];-S9CXES3e;P
67C=OH7bc^a>4BTYWK2gXZbYbR^C4LCSK.E^6]fR/0e.g^(7>9Xc_DNR^E-^_.Eg
R_+,F#R\_G,N\;d-H(R=T17-ZNOcK>/\1YKNV7gMYD^Ef>NB+WOPQ.a7ccK^UUDX
7DeP#cVX5GZ+Wd4+5\TFg_.H,;0/\;:H>7YQ4[EF39;OAXF78AP:)R.a<,Z?=caM
(@C-2R)dcM8HLF:TX&+BR&R&LI?5,:Q]9K@U=09e/QYA.+.c:HZX<S7V>7FF<^#I
YNeEHP_/PFZ<_^M9g&DP<>F-c:\OFO^gb.FP26b7<U+>:[?SGF8T0gO(ZNHVW62[
<K0CP<)\/e71=7Z-H=0?e+=-fPVWXX(08MFG#UN,,f17V]+.f8H)B]MF.H(d#?S^
ZU27M>XLWb;c7W\]+Z33T+R<J/NXFKRe&I4_<TD>+L+7E_FN5D37f.Xa_9[PGg/F
[^7_c]P,B@>cT)>C)ag3O0Eg5I1AdV3GbL24QX[dH?)A))F;;Y[<#0.\b2<1UZP4
eF3.6,47d3#(F7\&XUK>5UK3A<GLf&WD>F.7e@73\+Nd-d7/6b=&XS/-M^(E9Z^=
#Y@@O=YB^@-4=ZM#3UKBR1A_WRUcH,-AGEbRKbVde(Z8FQTVAVF3=0_(2CO\KA@0
]bPI1C#D,\d+5O6I]B_68<6Z89LT\Ieb2Y-FGJ6MU^B^OWc@_2Y_d[D>T4Z(L4eG
0?1X><-^&aY:9X3=Le@J2fBa8P=5(X#YG4;9K(HG7/4>[O?B<A74R:D2MKK;XF2d
29)6;0DTHP_Y)bX[a5M1F4Q.MHbY7?-2,=9dQAc])87Pe:IE/:,OC9H41T<8=(&J
M._OggSOODa()Lb.0.B9-&WQHFQ2[,TI]fAE4MX9Q8T1_G-f0KSEHW=Ue=SU#ce.
R.U1^B>FY9LTgV<g72cD65P?@S8/GH(QZ:E,H6aRTMb6Fgdd\PV@7RV,M=?SIAJ,
-8ON[TN>Vg&IG.VI5Nf_A=5+377XF55g+2P@9:OD_NQ7c)(C^&e/,S0@ca7FW[IM
He=VcPC=?AKTWeD\SVWBQ0X\JYJSLJ9B0[)W971&P4)cU(WWcI8[(HK&>+d+)Z.B
Q?gccNROIC151cgKXZ=-JCL/]&C/ML.^6MN=6VEQNgbI;eEEHQ3/dBX)_2^?9c>M
.LNa-(&/A<ePA@D8JVYHLDYK=;JWFYg\V\(]Of2b]6Af@N>08&H99e,K#Sg9DfaU
NJ9Kcc32C]e+K3T<?XDL0]GNX/L;K<-b?HgH<J3LBSV@FIK+^fVA[20#_#D>Z?O:
K[Yc,.]-4MP4e:68-KOLP9EP.B6]N)5),CRfPJWc@4></+18CA_4RF-X?8^#b3+3
Z83HNC,E14g1&P^?7,2:MD#DQU#aGOXOLVX3+01HU;+ZCI-<&Y&J4d]#;SEIUPdD
=Y#36_DPAQZ,Cc-NMSaC)Y?##RYH]8#FBg13a&T1(5;K5gWMQ=4?0Y>-#5],L^J?
;T7QAU(=PdfR8LEV,gB8QR>g\ZFHc,KgA+X82Z]AV^HM@[48-BD\,^46Nb+Y]7J>
1AIbNQZ2I>.aCK;TIU;_GOU=LYB[Re-TO4Y]&5QXd-a<>g7g\T^]IAa9&>3F@708
>L9\FX.bU2.>>f-H#VG(3SABN4We<\JfGNR9:YLL#&ES5G+/BGaX-T0\KfB[I)2]
2Y0g/+3A-8CK[]E8;ZN<P5acX>UQW_[?80,d6LgVc:9E9^;1F-.0&Pgb@_?J>Zd0
V/NRgNJJ_FHL-c8XKGFU)dP92<OJ7b;?JEBcX^F:CZ18([:_10_PbCZ9FD,Ud2J,
((GWa,aGV@D]6d>>@1QA&87:;>.7[KNAN+Ig>KbY]@?3T?T4ML+G)4N^N9A/Ug+;
@@4PcA@5^-B8Db,/SUUZ0>;WM@ZK_:MIEP>,)>QI,:UcJ\d#_U]:?+J7>UD<V;Gg
GE6R&3E2BQ+ER.=B#V6\XXOOEb1_&V+24@,J,e2QbKcNO;+\9(/5Y+(@g1KNg9X?
^]4IS5E<BbD8:\YVc&,ZWa/Z]g0,?W4Md,Z;f+KQ_UK)X/-X54CR5.2?XAB6L:>Z
a[AeESBW,a#BRS&D;1>3#>77[D9@:)^X#X8<K-AG5KeA6>c<@8W(R/441P+aQ1Xf
c-132b_W6gEVIO7A@=cHg2C;,e./L[;&7Wg?VCEb1J^[8_FG9^FP1Ye_(P8J>WTS
&]I@TK4gA#4g+7G@:bgX?EOO,]4#@E;Zf6?N</e=AWX?fAQeBD7<O&Ub6W\+L?+=
Obde6@^O)2&9a7A<)&&S/LJ.Yd=1/&0JGKOQ8L6CaR8V<R<,17:P-F0fgODVNKX-
VfT+YRDD<E#ff7S@e)7;Ua-ccX[S^V,dc8g]R)OS76(ZO;(7[bcQgUQE?Z/.DWPB
fW:+-V7+,]YGN#>L;>GI[OJbQU;.++f.?>F-UZab_f+E;#U0.HeSJR,^aGg)@50@
QN@VU=?++QVPNVf5-4:Q,BKB1J\LCJfOA--GM:6;I,_L#K@;M#BF#/9KK.b1g(5X
F<)SDO;J(SNNE?Y3NBZ8AT4&^::KJIP0-^[DY:P@XL40fVf9S<bRR(,3M)T:fZJ[
14C\-T1NI16>P5L>ZbJKBI2-1D@=YT\H7-B\_>(CFbL(Hd_5II])dV-V2I]Q>7HA
DDbKUA=33XME^e)Z_5_Z/B;,@W((SE:bGK3OWLP_ZY#Y?ZS<&+Y0HK#,PP39PW7W
eGbJ+MQPYCf@:6KAL[:R8eV4eW[RX#;1-?VQG8A=<5I^fJ-2f;N@-dQf[Ca#I3,7
POIT^/f,3g8CDO871&O.T>0@JTFEGM^D_2-3_C;K:U8>bF^b,2=_dAZI]^TTG>[g
SY?aT&J#C=@QXfIQ6^b#/[ATN\EW54#YNfF@;+T.a)eV3I.UBgZdTW]/A:V//DBc
gT#WgeUMPfW:B=3_O?CAY)DcQ6dg)H0#Ec+CNC/_g@gL8g2ACOB###]1:57U-B/H
C105#9F)>)0#bQ/GUYJ[UN9:M6HgKQEbA\S2e?M-KG7TERT+N;[JI=>4Z1Mc=AGW
YMR>\^aHdO8=&:2N;,eB7-We(1C9c(\RAR=]Qb&,4a+Eg?4^b-B1CSbd>+)M<RW:
XYG^&D[e+?7J+LBa=f=.J]KJ1+V[M5Yd[Va\OF?c#Jc.\^<6aZN8<;>G)@f8R_4<
]:gdc]^D.02S=JQ4>f8=[E:E1?)[W_>,\&P?I@&bVOg\,?P2Q8A?e88],<N[F#bN
TD(P+54#B=<7<DSaf;MF7(L&g[LTG7(cL3=HTD\(SfHZe1OZ9f,6-Q6/Q\;>5=AL
TYGP/@G8VMOLJ5?Ba]#RCJZgCMY^1S0+Xa-K[_AHceBT,eQ[\VX4:V2^9Z95D=R?
)ZQY)(b^N;N@[=#/MP0?5^eQ&/400Ze<>YUB9WRNf--BQ+5I5S7f69239;URa^b1
&VHG#(YM=8YZC8SY89-g09&@/&@gK(Kf1\M7A+EP)Ha63<B,ReCVWW3UWY4B]5:Y
[](MF.-g1c+cDT7.9#E;D0<9V#0YPAQB9/TS03X)8D+_\2Y9D1Wb^a[[69WE-?3)
cO>K[,-dRS^\g\6NSO4=>7<-Z;3<;8GP>EE\W3DP+Q8a47WL<WWQ-:FC,M:]//=Q
3bPcI8=F+S]@/X^JQ83,?#:VeE9eO;OK<.<B?\c=TI7VJf9be>^B#SAcRPDNLVI(
_>.bM5#.-\370DBYc2Kb>N1Zb3;3FF2H,4S^4M-c/O--76:PF0B50?g<J[IcPOMS
HH.72S<1K1Y\_2e0ZC]Bg0c>b6(fg_/_\=cO;#3DJD;[@,HBHYU+0:Q?0b<VRZXF
)gZ/Q,/>UE+X_B4)aX=c@\):f0cRE#?D;Z2:(,I46RZ#NWW:1JH6YW0>OL5U&-E@
+P@^,0],2UF?4Q_;EF,&9-LYW@@Da@9=4FEV91(\D><UA5GNKY62UW:A,6P@V<C7
IJ#fLNdO.>@KNB4gF#5.I:Q\,GIg8<R6A</6Q9#cVZB-29L:]8WG/B@AIg0AUUI@
CE-aC-^GHV#YFPRPX9T>F]D#20Z7PC/N0>A2V_LZ(-FJ)4\45ZG\d9U8b^fO9]O#
_G/LceIB^)IKF#6?M]-0Z?2\B1F[>f-Za=8_40]^\P=.8.;Ya&W[K:&8=UeD8SLb
/7?BdS@(<TH5L_[\+aYg_R-gP;2I_](JQ2@=f4cYL\HY]MNK(6):a[1/[&RYR[=Q
V5D]f=]@9_)8).L^g;VJX+=O9Z8GPU^VU&F;CY)23;2c4T.N<V?>A?]/7Lg[YIX7
2XJ266.KKDZ1&ae?D-a@;4/_/ZD5K4<8_C-.g8aOR28Y^,D[Y,9>:7T?/;d@TV<2
g5O-]VA;S]L3[HGN&:^#2G+aA?2g3I4EBa2c1+fCQeEWHG2G+N=DBJF;Z6IKS=X]
9TUM]TUC/C.3:8\IgTTd^QB7F&(/SIG;;HcFC1C/5gZO_Z:?-fCD^ASQ\b<Ca(.E
3?E,6D=:g-CR6\()6Ye?#Gf=HL&@+^1#@M0<]-MeUNeLX1E-=Q:Wd6(MI\egMLAb
:4_2c<SNeQ@->76f4S)Q/X2U-&F[??SH:..]]B]357D)5d)I8GR5A156HG6W&49^
4#]N/I,.M]1bL0Q1d[V(HNgN.9#dPPS_PcgZQ^9[b6cI1+Z]NDdabOIE4Uf:A9e&
bK79VI<UXJbTg7,079PFIO1VaNSSWC8R:#TgQ207+,Q,C<[N?d.e-aY&YLGMSdL5
)@EU/TgUe0cTB-KW,-SgWSEW6\#d&CTFO9Z)L49\Le_,D]X-;<DeI/=NJTTf?Ba0
1;EE.[^QbT#HCH\VV(JJ&c?70cPb2a[7e5a;=3PZV1dL@TQ\=>BLL7@gK)&#<cI6
:PAWK=?G#g0e2P26.EIH(/Q5\XQ;9^GVR;Qd35LfWAU63G[aG^--)1-([)TBJ;eR
J1HR#:FWN(WMEG?T<dbV288EFU=RHe)COaWT@-)NaaaD+XG[M4@V=]FC]_GPXKXW
1G;W@cBRKd&M.7#cHJTD^BR/\#+UKMP)JYCc.b[^8K22f#6T&LY;/9@g^T\fKD;]
dd,@,CNJFPeH+CYO_)=b49^Ue]57eR9LY>XOH+c-0(]a;G:=a]WD9L]F=]E^13g+
SB0N(,e0@E]&LcN,-M.(?EaIR3L_]3fV,\1GHOGZ/FD4eVKOJRK,2.1,H1GPNT09
f03(T]A2YF;cDJX[:bg/O.a>>d]AO4;DT)]+f5).]M0-,-Y8BIPOZI;1:eAeJ67U
58b<-GaT?;43W.YKD/gCbO8aR.PA@(I,TD8RbNPg@+Tb3:O<B#,d7feFYC0^=T<+
He.5f.If^fT&75[)H+I/[KB;\1f8<+@^dVW4_eG)[bL4d0We&TIJY;T\55IXRX&7
=TC\Q)J6<+MRQG^,+LH&PO[aT;(B7RD)fK6;:-<bCN2#=44GE780;#0b-E>;Wb=:
-_YNIR<GQJ87X>A9@PCESbGdf(TLaMe<P_)Q8EZH8CHR43,e6.[4O<A<C<[LZSL1
8RCF\I9+BXdg6_2<b10D8-,)gG5M#D[5PZ?D2W6aMaV^H[IH]5&ZLSZLF:O?@J:2
^?P0Z,U_;AQb#c?(TTdKe0;4M\de:GUJ.>JA(fOL>6^IHPTTgI5V+0>>-0]4@W<-
8edT\,]CRUC\BT>La6Xc06N1LQ89^N(>2AF20<,A_ZSN_Q8C3SB=F)UfGJ-YUPF:
2VO[GLXM#WUZ<>&^&W\U.+^G3)S(^BQ2D5VC-QW#;?Y=HH=:.#]D\FDb-@T#=B]E
AO8&A(:-<fIg\5IH\<-O&:Z.MAa=OO/eW]2HDXJ8RPBe.@bb8eFUC)R&9NEECe\0
[8\#-2NQ<4L6/@@MUE2T:TN##MRgL6/cd]FK;f195_DHOHXVf>MLE;IE&PI0SJ,J
?KN41N46)7?<B3H3e.J4(J>ADRV\(Yg2;3Cb\4f)7S37]g-WB6AFLNf[&cN2H=JW
+_EI;7TS3)[B387g6TU+JQPNd7Kdf>7B0:-)UE(S(cVJgNO50?8,@(AW@@O/eIH9
>]BcJ[OVHM9fRCgb9Z5@93F_:ca()<VT/9g-4Q&3JAfWW8YS<?],5g.G;;b0<FcH
,d]8YUg>=R9#Zc<fB:&@7BP\A:f5BVA-O5(.1IIUea#62QbZd]9e6R<eN&7S;TK+
.,BgAH5]7Kd@R0;_VQUXd?2c1X@9>FM)IbYa2MFO5S9Y^fdX,UVN?WK7gbJTP?)K
.(-&#/@8G5]WCOcK?](\A>,RB0EQ9dRO34IU+NH#DL(^=@06cTKgeIbI3Lg2;\-&
V?&T5CB#(g[SA_f]QBEG&_bE6-f&TL9W&SF[,B8+38NDF5e9-b@d#NcXU.\HD-&L
P;UX(UL>-g^@P@M?BM2-DR78GUZ>3bJaYTZ?FAET#Af@>6_09G1&_QZcHWgTMa7X
KF3,7eCLRKb#W.O_)&JNfJ6;fHH1#GF[+gc>eZEU^Uc)KRQ><W&KW.8QH])OQ00V
DdW)fN13<#MWJZ2IKFWHGR66AD9T(U?,(?ERJWI-EK.EB,-DSZ1a8P6^HA2EO6F5
G2=EUJK3HKD>aEAA5KZT1YF/<UfSZU?BBT#c@30_@TZ:-e3>HVGg+ZR\8QH0;b8W
.+]Qd=2V2FLZX<g.:X31bAMZOdOJVBad2UZC]CBM=E8.\[S<:15FKC2NL\gI8.?Q
@Be/e9&;T8-GdI&fEJOM]CKb1db=b_:[G.a4U1057E5:6,1B54[Ue5BeR1+:9\-0
\WJ/GFAb;6ZeO@0C3cf36[de5M5ZSPO1989dK@Vg>]c^>K+gPH&VaY;\,>Mb[F&Z
>=#_DY_2[X&]4.RNb(I,Y/]H=?>LLZS6g7O/LKH<[^YF6R,4\F,NBH#12bO@FIDH
eI3b8b,^+6\Y8(3EQ)^?gd&PEd\;RWCQGGgJ77\I\FX\;g7f>&bDae4Se^3>,Q&W
T3G6d#-90XbFYg171NWUgYScVY:2)/7bWN2EG4SZS-/<9F7E]EgS5cV_fZ-HJ=ZP
C+?S50FU/U,&a8^^<Xg.0O[(0:9VT==.?b?X[1&Y>G^eO5Q_P0&UbT_ND^:D0_2<
^.A]7]FMRUNf5T)g0(EBQV5)>a6SHeWHaRZ2WTD)cbVT#I4?&H1Wb9QVL9FM1=85
<P),UX)3V<;d:Pg>:\6O#fX,SDYP4aHD?^GY5TE(Y]S(WcdXM3e>;Q?7U0]S0V<(
-NJ/:U6b2<3<SOZeUN0_<Gf,J^>)#Vb?&Y:RV9c_,JVE?K)Z#4D;18-d8Cg\Z4Ec
D0OV</IE5=6]b[JYL6HRI9A,A=78F?XB\GHDXNW&:]7#T>H=e#eT#GED:dPO-/K3
_6@PV(E+3I(L/0]b5[V<GA;AK2eKQLZR63f_K<AB9U9N(e/Y8(,D\H;J4/^W5KGX
OXRC^-3X)IK?WLK<FY],)Nb2bX?c^)W\OG#??DU7RH&P8e/M;/-]Xbd2I-GH5:CA
,2]L+SS_#HK=5RY7P^##C4UAaNRf:^Q11Y3T,Va=2.T\cRNe)4H]4ed8^88NGN>X
/;dc]\PddEP.e0XTTe?Z^8UQY9RCA[P#@QY\IF0_HI=WD6CUe8;AO?2Y^M8T:7?g
B9+g\2[1LO]aRF;0C?M&U2#9@3^LUAB3Q3OdC<<D?&T\f^>5)@UMW<?48(4<Ac#U
P[f[d?VNYfYFeV\D^K\KJSW17SN(XF2a+AgcK+1FS_3,2RJW&;7dP(_VLcfJP=c>
e.@_UA#?8U/Qa1g_7f@K2VcMbGJSc<<@bUU<(.2]MD])SB?<2,JUD+/&7@Bg&aNZ
ff@^D)BSHU#38BH/Af[D6adUf2gg+VBRZO,D?[g[HYI=EcZO[-,AQ(K_C;[806BC
7c9,PD9R/CNC/DW9LU]:=bdE>>&dE[(NP,GNCa5^daN89BXTID_8A.<+1RMXT#M[
Y^L,J/?R-K+CFg0C;e>\<V19b?>T^@=S3>UB(T51/;8Q<N=/6DHHa]U4\9+d(Z7[
8eYfKN;(fdKITZ1J2gS1^J24HEeGIJRRJ:2.)9^<#B0Xd<P#D&F#g-]?+L2XV61H
3B=H9a2/H,,T8#D@:/_ST3D6A>V_C,@g[Z-Y_/1V=1IX[QZIIX03_FQQUd.0SQ+M
_<RQ=;_Q9_T+N0=S>V[:bO#A^F#\Nf?C?BE16#J.Oa_^KAVJG^;EZ_gf-G>DaDM@
cOT5;T>W;DTg.0]BVKQ3cO_=^BF/#WbQUBYXTK.G:E<d#]N#PXKGDfB\O[R-<#B>
W&+8A)\fYM?gU0#+(64S@GAX-=.992P.M7L5(YM(@HBIfSa2+^XT)Fb8dMN&2S\e
F-IPL>JW3C>QB(>;Qc5NBc0>/eRV74+SZM3NQ+/KK5a+[/PJ0P9:D]J8Y4=)=R=]
@&1L6>R?&I\4H8)7c/MS9MAagAK;.FMI#^X[E#O)Y26I[VOUM@:aN\W?e\db#Rf7
c@G@VL5=/FY:K+A+f[EXW1,g.7B8A.>M>(3&3:.#_5&GH3/;g]]_4CN\Z,3Y785[
X6WI@JXLe3?6_gGZ_JAQE&dZ98H>4/KcCBYf2)SddJ(a5JE:?=#/?6KVRE9+D_ZI
S;Y(\HQC&P;,Q0.:-4/Y7SWV[Cb;[fVHg^SG3DGcLebfXfcdVOc#/TO1:4YL\_IS
E^eDDE>#Q)@eR/aRFaV<C=KEg(J3CEJPbg--[cWeS1RFd7-Fc-g@&2b[XI#QTgg]
0)a)1VM/E-R>?Le+73eGD^SQDSUU3-]Y;UEN.EANfAC1V&:9SLNcH9e20CJHG7e.
8Q.[;J+G6CH/eNO42&Hb)(Ke^g=<_+c.eNaNc&H@@dNO)]I+0?OT#\6;@aA.3X;N
UJIdS-C4\+[AP7S+4)O0A_bU+0:M>K?;36;V9@0]D3Yc;P<T9S-__]f1A&fS9?[f
U^LSRb/8#KdO+>KC7?]Z:YZ7gA;?fANBN(X&(;-SSK@3a994HTY(,=T;4(^&?>1Z
>:P(#Q.-B>:cbg#If9W)XLg_\DH.=?_U<:SBgfLO:@)FW1fOVe_6D.FT.(SFQV8X
BLORe8DP-@UIDJ&,AgPeJ,]59ABB7//GV(5Z@&_>aPE/W(3JW6(TD50:=<F8K\3)
NYQ7/G_]4c:5@#OP06^fPGP&VS1<=->3J.V2ZOZV0Z\4d5K.GY7RE,aCZA@Xc,G;
7O/X_Z[O=>LTX:=3/Fa<<cW#)AZYSY6NWCT(_=B//RHcCK=Q>]C,E]9\@#W6>X8A
Y&FH=\=5H<RHT>-,8EID4(Xfcg2(.6d0YCPN5]de5;a1\[O,6GHA;Sg1/I(@(6=9
5V:Ig6&D.B-KEU]N7Z@Oc7XKX14W2b<F+B4,c2b0AL64d3+Sg(Q)796?5Sb\:+Ee
^b.[2JHe[GHg@K/XOEA\g-+g\_36I4+8:69cVeZTGK_F1(@^RZeINY<\K4eX1)e_
+[F[5IMKZOR,&[0HC4;(M>cfQQ9dNUV6Ec\dg,:,1ObIdUPEJf]/^J6d]a4AP^<d
Q@f0,GXED]43]7;Z:XL(^9\PXI>/#I15Tgac?2RO]dP+7OM#+G6O&(RV@CZa28RV
AZL:S3@Db-M=C><N_:O&dC+\#O?dXD)a<NY2KFd;dY=&7fE#^4=/-OU5R/3Y@fGR
1]TC^0B\@;S[NK13=J?:/XZ3:;d^KLAMd-1MA;D(GW9]@gTK><?JCAM+(EEW<JPg
,LS5:#TEE;4B>c.Rgd=4S5dM-T\B#)4+S,,bdAM-M8C0^GI9M6NAWb_BO87YO+F@
cccZTNB^+e5=+^C+>Ye<KY;EWM9RFgcLP&#Zgf[]d.fPe2][<]+EYbL6dV]\Hg/<
,^fcI7Y0S[61XY>G;8U\XN6?S-Qa>9TM&KE;+V9#<#=)6:^#eeSaRVSX@)]cRb6-
4DUD>#Q1ZaY?c;#S8#@2(PfXC6W1AYAJKR(=J\QU)ONERL:R[6<Me:P48SB1N^(U
(I9Z@HT[]7E]ZVT46/128?f9=]:PABO?Ed@MY0JP>#<N#fHda5bMX]M=H@9[C(KI
K6d.b=RM=C<_F2#7a2^_2Y1W02RId&]JQL_YV:N=MYO(U47Ub33@G=F?cQ4SE]AI
d):HC0=.,)Vf__]MT&e85-4D@FA#X[NKIMWa]([J_&P2c;^5(-gB&\2V63>X,0d^
+VJ7ZK][KAH[ag6[XCDW?AUU[?&#)2;A8.N3L<YM89g<&?<AGZCP?6T(0MfV,JR[
?4G(7[L4#1EWJ;?I4-@&gUWJ7,6.ZaEFP>[:GQ)\b7GGDI)O2Ae3L&NI41Ma;T_W
-RYYeO?KR,PAa)2&)V4]NMC]0B[a(3JE)P>BBg<I>.+NRG?Y_NdP[CdNNdPLZ(M,
Y3aE<89JJ\F0g=?^T7GHV?0eQU6Xaf:EFW>[gbbb51OS(02_5YaV?@YY/@3<K]:I
JQ-HHA,)fM@,MS.Y&g@-?Fc&FGU527]ZN4fBFE9:<N[\>X/.CMW^PHJG_@C@?=DZ
3&&=[f=9b5g+2-2=Z.\>AC\A.<1&M:(M)g2Dc<WQgZDN6#c[LA\dC)AVSOUPg;H3
8.U);VG^]U5SSN+M#GV(/fdUg;a[@Rf6e_.)A+>-U:[:APaI?/-S,_d6R^_&K[W4
0VYF&Ze(R[X#B0f+Ud:Td]<18#A0&>F18G#IRO;[E:d\8C>@bI2PPgE3Zc[eFHP1
-]0/?fF7b+9caI7-C&<N;WSSVf&H;]D&7b#9Z@HdCCIYc02F&YHOd60T_>;/6(K#
JPINCFca^c9>DV0]&CRWP6V7Bb1YEd@X167:ADfQN(Xd:_MP7KO.^3f7<NAO_gH7
52#=W,QF;<+S_@^-HLB3HVNU?C(OB6@)ASdM)IM0?5[fcHe<?_@0L89-;M_GM<+K
:A42g/],W+I61b5;^H20M?1X5J3IO.I_V7aFRd<ZYP9#GcK5,g]0ZO=&79UDKZ^I
K.LRaB0PYIQDBR((a1)6F]&=S=#FfJ;MY<R>8H=(f4bFH)L_(>J[R)1_TIeJT5PL
9FU50E(^(5cF?H,L1FDH2+PfXXUIY(^>?73cB>5d+(U1_dW3)=?U0,Z.@.2#>/MK
VT6W,Ke#-[P+&KE:??+e>G<bK6@TD;O;0D,A>]#P:/@Yd_)W(4-ZVFTOLU\?4-24
P+^D]YVS3C:L7&C^==-T0,:D.2aDE4TN@8RdHd.:^Z)0If65KN?a:(Y)H6;Sg)SE
^PRSN14))2M<J\VA_F.,288@W5aKEJR#fac5IWP;)1G9VFAFZg(0@MTH#LRd84+<
VW:?=\&;Y\P:O8<J@:I-3/FfU5a.eVQ.\FQg>SD5^Sd5S6OH(;T3,269V.[?W\/0
?]/@9,KDGBN5b,P<fLfSQV5OQSU3,7T6Y42H_=#[EM_43\b0?8P9@(gM6O80T81g
M2NM[)+<5J9f=cfNN5QT[&G_ddfV2LE0.+0CK/f+8;0[T6G,&D1#7MB@^C-2,=YS
_Q(c\E_9E+Z;]B-(dL#adBH(V@2==Y<d_ZI(<A1Yf7.417b>K.Z.EA<A<]A[-7VF
J9DfXdW:9/TgV]<>6TFDJ3)JQ>IX]J&dc5A\JHQ8,d<X9+>=OZacYGL_=F=)X@J.
fe:P)=_H^])-.TEc[)eO3FQNbS6@=>2K(R0U3a4C9H/&K&,8-D/+0N5PMM,J&I+D
3g;1NA9DYN+[&Y805gBE[e5#E^^X@K)Y#@87+8C8([E6F&2U<\AY-bZ1TA^C:GJJ
>K66)g660[7Lc4b<I2R6F\I6U:=./?4:Y?O,_O,c/T0JfI19a8GZaQb?\3EURf^:
V]Cc<K)S29()ME/=@2]02cF?&Hf=ce>V/48,7DWL/+-7V]1X.XXY<9HN;e2?V>I-
4:T4gK10-[+RXSB@I#@)L8#TK27MM9gD5gb0IX:(W9ZeZ0^-E6>d^b/bL9c]]0fd
?:JJRF&2g^WfQ>SV<7Sg(16]=ad/9&>8a4/3YHb0D5e@6JQ?IRZ92NeO:bKgE-;B
2XW5(V7^K2HS.BW4M:VG-<XbK,(b.]=_LR=&YM&[cQ>.&0U&>=FNZP-FG[d?ZGG2
)[b41#0MPELD=MM>PfS#Ia-1+RV)5&4aYLI6?;;S3AQQT#;4KA3]M]&+HKRL,PdL
\6D24:A5:-?NAODcc>Xb=T0B-=B2Lc7U8&4]25?@2Y-UM@B3IZe4NP:)99CHT#(X
f;-^bA\9&C?=e2_NX]15d5#/\^F^88(.+R3,C3>?DEHdUHN=,>1W\?/[W#(T#U/<
UeFEJ:F-XSZd:)8R@W2^N09/d<)dR6@<cVcGWbMP<>.Z1SP+\Fc_EC4A:e=9L7.A
KcgGXdV=;N2A1DX,=0F#@D69aYA2LF9<=WPS;TO@a/fX9g:c#_-&I.5\8Od+C2I3
^a:3+U_AWYXHL#CTX4E&SLO+R7B2d>e4Y6b8=2ZTIVNL\OQJ.B\&?Z2_XZ\(A4\P
#c:LVfg7>WVSGY?[Dc7@fP\9@GbfA?H=3e=TYPT5#a,P-R-=5]6#ZM\VPQ1adOQR
3V[&MN_;VJZ\KbD<>8f@1]3EG_IZg\@DUW&KS7SDIVaY&7-A[U63e<)/e;;&+<7Z
=ON>>4>XYF&B7T3RAEXO7NUO6cP@&cX5.\9:9#cRQVcRDdWH3)@=b22d5\f2O0]=
<0CF#]2@/9_4OI.KV9XSb^)fJ@3;DQ\2S\8=J2#UgV1<C_NK\De>U)3]V&K6,&J^
eU@eBZ;/g;b\c1T]86J1;RL<J?FY20B9S?_g\XYc(XTPf^AZ9G-S]HUd#a_I0(BV
1E=/S@cL1<XB=OHONfN/P0N8H5^7;1Uf)@SV66>f3/L51F?5[IM2)WG7+_K+DO4g
cQ\b2N]4X2&DebA3GcL+F8c]fFWde-<PP@6\LT);EUR?Nf4\;;)3&Q:?8gQ_OYEf
V2ea0BBfFVEC0<>OYfWY,J:^75<WQ>=_6]1C9K7#Bb<A+9IN0M(K]^5PE3?6JQUO
>8S5gDE@\^WM9L.fF&74MT+,NbENHXR4Ag?\FdB&7FdY0ZS-Uc=E^^DY4^UH8=ZY
PW3g5;HFM_4(;\D#<JI@:D(GYaJ/Z:a\D,V)M^d)Y+LK,#+B[L2QP^d4@RcJ;L3Q
gIB?f<#7UgH\@F,44V9(X>IHZ19^>:_30.J&OT04fUG9+[XeK4<,68,P@Vb1aK]S
#eEQGFB]=(C-W.8WWGS9;bag)[dS2Z?0WRFURM0Mc2cBdgN3GTP3\A^Q-.)^WQ(O
Q)J/3e3)Q]V<^L7=T6?V+C;2F[S8KF[b@faQV08-\SC^M=&^P:]@3KG.OP:B:8Gd
\)>=3DX>N9,G)4)Cg)+d9I+eQ+8K6LH??KNb:>D0+?Qa:XdX^)96+@afG975=Z0\
Oe1S,I:-)#_DIC)0X)c(O9c@JVN3\c<>ZT]F?E)^]32>g^T-D&O-Z\-UZ7RXC0H7
MaC14=5?[ME2f]=F3Sb(G;I^OLO,dTG:O]XLN;bGTd^5<RU,AX(P4VR)(7V7]dA9
?(_IVQ^=3D]1^JeZ2&KDRFP<HGfe9MMK88/-[9fG3AAM-YG?2B:+=-<:KNO=X4S=
MY84caF^CBM?dI#.Ib+YeZU0N0JfQ&daI?6R?]DTKde4S7F.18RAP<g06;<3\9L-
+N+K[g3M[<]YI1QXF\T+Z)M)IUT(K1O#c)R]WHd\aV\M<V:L=H.[@B12[X<edK))
gVT1c_^7ZQE6N2(<P_3N9&^CdC^e#=]5\2@@8)e2[FT;a0Jgb+.:].LH>FI1dTG9
DZbXB0S7]f,Fd,).#]1,W\W_:gPZbZ5>=4DPJ/Aa6=)SO,3Ae<K/>O9B:Y6<g968
)52e((\ef9I=ZC1]EKXH0_@X=R),gYL1a[OI\3g5D2(bIAOUBT4d/g?>HHG-dG,D
PR.gI2:.H2b(&8R6cO;7N?=C>F&#W]F62e>3LZ^a#U9;S1\N_AdBaQMVL3-HLY.L
cPTFEYgF+T1EJbQR=>+L9)4AU^G]Le)<&C>ER@PMJE^^8LS5M3KS1?JETEKBLg?B
g6@0]2gBX8aA/aGB1.G&Scg6dg36f&9Z,RTa[4A9UUM-8^>gN?->SR=e_Y,C#Y(\
^-JHTGG<9,0Vg:VB=cXB<gG/33_O[YS<8OgbG3?Y:O#IG]aG;gA,fEPQ<M,B4I)H
_g)LbfRa0XD.=[P]J9.TS:4_QTB.\YPF0g58HJ>(KYQMM3cFKEO2+Ua0HI:/&P^X
U^/E88WKFRI)M:aUY;RdUPT1EV@@6U#FZbPR>fQZQ4gZUfdN0QWC(Y,R6HXT@TPD
D@3MaMMOJc;+:=dUcXWZJ0A[T(BT/G2A+BN_\(CUg@(K.F5>>>NZ7Y>JJ&VcI;b-
U4aS#V;>MVX7+4]X=JYObBH,:Y/U.UL5^e]@,6IJOdg(+[AU].3D/?OcV1@2,\)[
d5/R-a_@aFTZ:aJEL2Kf37INK8>2a;?/?YP+L\<V:]-0L:;JTX9S36G#&3YRdbbJ
afFYg):3;)=\Q\6faa]70d0b:8O9>QU;Q^ga1bdM/eBW:/bR0g@GV++K37FG5L=X
A;FMCc)<(H_E0Ra@A>N&2X>fZ24XYbRDBKEd)^2>P:_c/T@:G,_K^/^)(S4.-<\3
Q]c2Pa]-J=WI>Bfa4A>eG#7PC\QL^[eOE.FHR84A@=b/F&W;WDCg10/MAZ?12^,]
NI<gE:11XP^#HYVF7a;5TT4T>+1PR75+A_5)XENAI7IIgQJR6W<L&LQ6e]VEbW\+
]JA@2H:/.[a(;SLB080)D1&2A:D-/&ZHH<KGB3ReQB\8H<[e<_<16;2eeP>-0OWG
7c(97D668V\9,8[=Q31J0HB3dV;C\43>3U.[1/_B3XL>gD)4Z7G;U7O6)AfIOC&c
A>W??5E=B>Ac+[_Mc4V2YV9[9P]E,QgYJ&Cd0DTT)XRTK^8XCCC/91K]4dYXJ+@M
-+U?c=+H#\T+P_<[FD,SV1KZKfEbV#c,+9g\JJ:?=Ec]9Q[YPKPZe<O/[?6;MSO^
A>T^._W0WG3@TE;U)(L(PNRD(b(/fef>R9g3G>ZOS-/:\0#2gS1M4I(RNQ[&(\S\
aJNS_e-H5IOOg7cfbb3+Z]/\[cY&SH[0Yf5=^G=,BI6b(H,W?.&+@6TI[65S&&e7
CP)[V7+&66gfNIV=Dfg,&1V_=(-f.APR&LV7#&7SSZ\U(O_8AY[bQ9>WHL/:HW1X
XJd:^:+4QLP4E1^YT_e<eD,6XOeH]):@L[D..=N9A0b8?YWO)PWXKZ>S:J9aNS<Z
fG^QEfB1<f<1aVc-=V>c<OfGH5XQI1IK>K75g@>0YH,#OZJ=^EW(a-5age[IHE.+
35Gb1O\-M0M>RdWF^b.E=J1D^-V>-[:X=X/4?e,ZbG^&DX[,/3MEQGV;)-X,5&S0
O>D(EO4a2H\72U<F6>^M<eDLO];:DS#&39V]CQY_)fKG@g60HMCBA.PF)eD:JV:@
IJ><@XJX&JL4C+)b+>[(ATgADJ=;FfaUBDF;P)]-fZ3T]Q,a-Me>>Qd4]/H0<b7@
H/eU+.?-_&NIPOL)af#S85I2a^-^+RNaK^)ZF)<<ZG2WZcd,XU.,#f.#7AV.]V2]
SSV2U?fec.BL@@&LLL6_Z0I+e7eZ[Y0]C@&G?F::2+e>9&g2>;_QELCA=GKfOAU9
a)fTGFg9=Y,-<#fH<A9X6Hd>?10NNF.LXcD:587MaEL[XCEO^XFJ#:1J=.)E3]S]
M_#Z>3Z_ZCN-O9a2>f3c87+T=9R/T&5Y-B6.;M>B1KMF3b+5#cHFJbY/a?-T@P_4
5NI-Mg9Y:c^^UgX-O_WK7_25G+/ZVVgYM>MC16#),4Q5^?LI<-8/2:)]<DLdQY&e
4gf9IK85A5DIRd0f)Q@2SdZ>1[PC6C(16,;W7>FM[^&S.=aSX_-4Hd6eNd=\2cWc
U=G)B91U9932X);AR+IUAI].G\U>^f>BDY#VD?:bY]9H87#UeW>9HKU++D9fKV4Q
ELbL>SgP&deP5E;MH2^9IV,3Eb+:8ILOcN@gJ,._SWA/gZAWUeG+><g+8&\:b#M:
)>(f-;=\e2;SI^&8,/[AT0b<JfUY9=NG3LY/Af>I)5fVc@)LN?J5684YB+U0H);)
D7PI69?<9YfY--Z(<G_3#O\;PQNT:YM)2.YPT@L:=0Q3CIgJB]5M9?,.&fD6eA9V
L)Z?-X_P)34]M4cU4Gd;L/Y;PK;L_LA?-)S#6,VWb82>#:3H[^f1G^DPP&,RgT&<
FSRF1cV?V#2QJCaK=NX>&R;()]\>c;.O-024M)3HFS)bY#[>=fO?P5JMBPdULJ.V
57B&]a[W:/J=VK/fN]LU3a/)5Qb#d/W)9(-DB#FWZ3U_Kf5F=B5D[XT[Vf[F<Q&)
9=A,?S:G4eJ\ZceUT1-S0\HXCBO\B2N]RR50IeI^/_c#I_bc5<b<-Xe.(#2ON5X8
]=0:QNU,+JT1V<=V(WdI(X^;M1Tg&\d;YX)T\f&JEDPK<9(;O:VACBPRQfEPAYEe
AX3)d)\E<U]R/<bO/[J:FS4Nd:^RI2+acHg]d4GBCIAKMHaIUR>9]O:[W=J#-G;;
+Scgaf9WKX#SE?29dC+1(X87^#cW@Lf#=]deQ3B^Y\7<ZT;AVbV;fcd;>U#JB8O;
O533+F_@7c.CW2e7LVEVD>L5TUMEMAIX&Q?)1,W2-Eg]XHK;H0f8-?)[JM0c[PbL
adaB:Z]4T@#e/5]:V]CBI5ST/=TD@H,P[)16U+F\Wf>R3+>1a:+N<;V3.O;O.(Ic
L=;D+:CK7=5YW2XA.\?4\#3:MU^^cKcH#4D68WNT&SNI+bF)#R_ZHL#e\L^NIY\a
:MB[&]SGfF\Z9(G8A(A4B4&/P0=-(Y_V&c/@SAMB;\QEL;RLEX;H4OJV92I3M?c-
VJWK@GXcNIA(#^0b;<C,f@?fC)<fU3U^=E;QS19=Cb\.^<4eBT^:=5^V98#Q(KY6
IGOTMMX]072U2QQVYZOP.VGf\NYIeU^<2HK8XN9^C,,?^FX<1@F5#@E#O\4W&e_O
7T+IVeK:4[M+OT;VZ7>#KG[&QN(0X568@L<]FM#ZS>__4:(W_DFgCR<dP2eBE/UH
RG\WBffVg9^&>?\881fD0NcL).>cf\f#)DMX=I]DbJC?d?.-P;EK][B:_1f0W@Qf
;EM)R[6Z[6)fcXe1;c8Hf?c/T=(2;\1)T);D,V/aC&e>S00\ZaTS3>&ZQ>HRMg75
DIM-,LT^<>(EaC5Y52&;H<0W=#TCM7VdZC,cfe:.da,d?_1Td#,f2Gbg,W3eNZ;=
\7)+[0G@fB2]<,VA(>a_W5M\2L0WLUA:b2K)BG[\_P^6)SP@2&d@DD5,3UF02<)M
FMZKFR=b[8:#X7I40f,d-=DX326R]Be5)_GNXKRRDG<ggR1c7#M;<K_-4:O#>-Od
.L)gGNW3g.&G4GZD2&O8ETKPBH-I#?,dRA_/a5g>EJdATU^JfZF5eEUW6+VS_c7Y
4edR9RMea5JSGNJPW=\=/D4cL/AP-gU/81S>#X)_>([a>R0Zf#V6-T4)0e+(H:T?
S9175F=-Y0_+O)&f^&5UAPZ).H&,-QQfR^SD#IHdO[(VBaIGZa&4J>:C+08E03C;
FK>1W4b-UbC\(eC>>#SF3A#@N9M0+d.FE=Q71QO+86a\K)NOYGb1=IBL-P9I#C&U
AEcR5QLK.DI432ZMVA]:,>,R;][af#.H(1[R_fWBY6.5\,+LR+17[UM.U-3H;F>M
O;WLfZO51eMZ\;Hgg.RK#L[,DgV.N5@(OaZ4cY;@aD1SYU&L?b4U^L6G#d@030WV
0K9H17B9FK;(RQGI@U_Q>_\1-eC<[;,\DIFEM\N/)@M4.UF6JD)),?OI2PcR/BUJ
0JRd.HK_DIgWPW-YHgK/F[^./5QSP=:4)_P.>c@Rc@a>#E9I-M:2ILWJK@M/TUFY
3OSedL@XdT^NYaNF1d(g9Sd8TLV;c<A?2cP:DH8g&<8BENSXR#I?&=<EaV04QV3?
X6TcXXGd^)+@M#)84+0aQVbZMDJ3Z(/=R1Q/E8[5TV)3g&a^8TZP)>eG^+H-61@N
-8<[[8ARGY;>&F6T+IB?eUNEOZ8I.G.EIN5@9=Z2Y8&Q>LF:?eR/W\+VWLa@QZX0
,Z-XD?WT+6G\4_dUcDb@Y>FW_:6R(PY6]76/(EG9fKCK^P=X,dM6)3bN5=7ZT=N>
A5#LCQe91I;:<J4YgL]=I/\d(2de_,H1a-0,L<B,B&ORY/Q#0Y<<ZDeK>9c(5)VV
EG(=GG@6gf7M=?++?K1]e9cHXIP8ZDH-?)T=G]X)]TCMC;>#6S.B+c-dEJ3f1;V[
/BVZTQ/C6MI8Y+9L[2-^O#:<;fS_&=A8T3HY&#X:bEZ->/0R..PPA@e372RV)IZT
[8S8M\@,33^fP1_@8e9<;:BaZ+]D9<dY>Q4/:cM4\]2N((JHS6_c)>]R;DR9g#X<
Q9)GEA+aH1KBUXYY>g5R]:U\P7b+3/2fd>?g5SQ5>J/A<@\5I5S5NN-QgFLRSX<Y
QcX0If50)1K[91QH0DIO0XD2DGW@aKZU^gPUSHCfO+FU2AWM@Q4LU,1C+V6D+0@c
//9&bLVde0U07)_OTCL7#>+AL<<P<1e:9K2?b:.MK2X[;/.##VYI@4[35e_Pc<1I
VCFE;>EdUF1[aQ8AJ(]d-I@2:I>T4JF+<K]O[AAC2-IgdUJADV/SO(BIU_AZ-E,W
?.OCUQ3F1>0&S8g.ALUS0CSbc;6ARX]I(Z2-30+P>&R8)5aNYT30.#(+;C7+T]69
0]\;=.d4cJ/08BDQL_7ZEF4A0E[gGcJ0U>2D=+7D26OINc5O=fS(H^K(&d@VJe>>
a34XY3SR#NN\[T^.,GbS/XQ3Qcc_UW<d<:PH8>[W#)Q00/Bc+E9USV.+3E)]9>F+
AYQZbHCB4P4E]6g3E/+S4I]JBgWSDS:0d3^9JXKc&5RM[eE>9,E7#(PU?V=U^\O&
M@RCgPKG0+Ed:@)V/f&P=CfK)8GOU&fH555D.VYd)&>afPb(<0>O&B8?:KS-1M#B
N/8JLATQ8(g;e:<7f:^,\>Q;YX92F_Y[Y=b]/C@+G>^Zg(QT_LfX_SeL\bSVWaX#
S<IYC37JGI_[4T0[INUT/1M@@N.Qc3IG[CRI2N)b&KSIS#Pd&LQ0,FC1Me[ZCe9L
3-dF[;eUc8P:S(AfFLeDYV:WZ+F(0=/9C_T)5;5J5446=&4L-Z/N/;\JP,,Mg\Y\
?0f)(+d7>>D6IO.7D-A[\Jg7&.BB[C-T1O2:AZ7=<00MOF8GTXLDFd52,.S8_SE(
>I]^-f?_(N^LafG3KL8L>O#?3JT7P7I\_<_M4Z0Ec?B5bSX?77-\I/Hc?e3I5;BQ
&J(YTH1JUZ6X?4XY,&PGLC92K2Lc[TL+[)YbUcWT3Kf;RDN-gF1Q(<79g6fg7B02
,f:B(&F5N@ZETBI#b24Q@MR>G4AJ+F,M(PGJ>MXJL^g3ObP7]KWMJLH&Z?>7McUc
G)4=b=gDGZMaOT?13-5J[SHFF;Q1GA[VH0)?4<F<I>EXL:^SKZE+;CAJ)_0T\_+M
8<E_2<D#b@?TH>>HGIIf:C>4>(4YGd#,62?UG,[P8_-_>CAXC7+9_SUSP:(Ie(?7
TQ4CSH3BRTUaM[ZG)W/R+^C&[P>SdBV4HA/bdNH3Zg4@[.IB5H)/3,:\Z99):5Q]
9-\>C7;=<O)1(V&X.FJ;4eOZK>05A)6H=X@L_TK6e6e)<&K((6IS#XC-V62/4]MW
ZE;-9O_U]LOGA>O.g?H(b#F-aR3D:6]eddH8:IXU36S;aT,WGR).6RCM-++O/:)_
:GFAZDU\<00de\(Mc4QV?+C7\e:Z6^M(@:AFDFCY^;BaM2APN0@??(ac,.72R0/S
<g]gC@PJ#\>)S_6^/>_<gBaPU.1N(5U@FS:3MI9I[DF69=;/g_-U7P^[B_M<U=)b
d4WEK]RV_3V6;<A@9?KS:8BQ6?eD=(EEDEAU7SIZNb:[efD3Z(aZD:N]dI/Y=+[Y
THRMX9T(.,JJ/I0B5YS+Sa@3faEOI56Y5VQ54Sf3#.JYZ97+[GU<20bCOCe/0E+g
)^<V\N^Xe4(IS6JGRf71V;DN#/\PXERA)WJW]\IWN6@KBK_e4<1=G3MZfN4dG<3C
QI9:=IEO<U5^?_SM@FPX,]T>WF,VQG_TSQ2GM&.E0X(TdaD]DG5Wf<KS<AH?3Xe)
fK(IPXP#[7?8,ZLaS:@c=:Z4J-aICg0Q2ZW[:.c?E,-eX\e#<]O;S<cS;12d5-#I
M2fH4cM6VXFFB6\3BEc5X<?ed]QaV1]5,U:U0,aS)JJOYf7.6)ef?b[^^5617+,M
eBYLe7@E8R,C<CFJ>(:2,^FbUW0YR<7@I?=TM\E8]YT0;UQSCTUf::^T][_eQ_^^
6):-;e1O:7Ye64QQE@(&aIPgZ)7;8J<d^TDAL43/=14_77J];LAO@?>e5)\D^^A0
)W8?3JV=:N,Q6K)I,0-&U2g;?IF)HO9+QZ1?1@-YUIeODdAJ6SUA#W3gTCM=1?F:
XS9M,\efA[CV>IX?Re+K8\O);)>G\_0;Nd[^<^.&0fXHF=f[6Ee(JN]IC3^4MJ6(
ING.UY[&[Da3]-RU^NRLTU]9LY<H+ObG3D8eBXE2&P[X]SGg-Y7=3T5Mf=NA#CWU
EA,B@eNBQSgP\cVMKL<Y@,MgYG_1)bD^P]8F^TN=g<4aU=,>5F1cSZGeT\[15CYS
e4DN\-2@FK35_;KB>DQ=_f6#;AWWc#aDZWORWV_TE?XLR^SFP=S<4C-L)2J^,,6C
?0SXFTET.P+77g\9&]#G6=Q7T)-#I?Y\gKG9Z_@[4HETT0Og5-3bL=20>Nb5.-I#
]e.VQNYL5]M;/&fDEA\[)5@3&\@,\:ERcLC4Rb>YbS>>2R8V@Eg]5ddA:528)+:\
S(RQ&fJ1&/ac<J@7E>#N.JGC>K_G\.=((P&NFT,[]U^T_Dc7+TSC:^_+&Wg[_5FW
F#[QaRWB22V8/b8+1HacVE&M6G#c#0F.&6^RBO@TXFe6\/H)PL/6I.LFUHee_UQV
RS\0D--B@)cZ()\Y<@LP&#d3CY@3\9&cfg&[DO,[,I5S#&PU3-\26RR1-eW8^=gP
dGCV;8ZJ4cTMb+F5</cLe;YR=IQS+<)H:S<Y=?A8E/IEUZJGZC^FfFZ6RZ,a+LYS
&c.5:JQVZX/\-/&>R/@a+0<b_BU3T.<O>(2VEK\cPbUfRdA1Q&\X<#QUf:PJYDeG
.#(79Y3J2FC^L3g<Gg=<IgU)+RcJR3Y=15?26X>)VffQQ71Z.P2[0)<C_OWAP.HM
(J5H:D<5\fMfI5^b5-f8YLE1F)0T@[#<R@O]#T8/KU?_9)8=+C[-de94Eb40@=LQ
<VP^<f8#?PH)+@+[].5N=A.1Fca_W^,YfS-c9TO>7LGKT-JKZUBHb].cIMfHRA\?
bNU;La_?5@PGE^A0-]3&]L_@QNL44846gMD;Z6_WM+K=EdDJfO44JT#9UU.@)D\a
6aRMZ:3R];X@E;U-gfFUIX2[_a[;9(314)BMfZfK3.[/@X:]S7(5YBEA@][fMWa8
//ScI=Ke(+PP7Fb_W[NE<C#=g#;aM(+d6S0+DA#08SOe(JQcTOU9:1F+1WC/4@@J
9dTg//c4.@TcLWC_a\V9S3bC_.:;4)IIN-38dOU/>=KD3P7#--=)aEQg+>c]c))f
2d<-_f>=A8RCGS=gB)f,O>:f+NO)U^5Df1>S?[d3g6_,P>bB9f(R&a]\5=4ELE-S
dfIdMDY,[PC&BdEKI?<>&#,S\RHHgW6)54_,gY6<+)PKG\B0@P3/BH1I1gF<OdF;
/bf7T0beF9PN?W79@(ZX/QYS^1dL)14I^D3M?O19O/](875B</_W80]0:(RgJ-2-
_I;&Z>Z]3=+?3^8JX8A()N0=T71TH4A_D7IF513B_dQ53]@I&X,-gF^RW2C7.c?2
/@ZY9DcY\T0);TZ^Zb^+g;=S2>+S9X\=XH,W\6V>d9<B@7a7-X)==gbIJD07)3I@
I(7bFbQQB;T20dcTa:NU?ESII#2^f=5M,5U35^&K5_:QfK/3d_SV#L/T1f<B7.FK
E,(/O3597D,N9NR6L+9H3Q4=?CCO.aME&-Q8+Q_W(3aZ0/]MH#c_9+W8788>F1WO
_RZ[3-K3cY1+SIJ^)1?;BDMS#-32g:a@V=VDM;G/#YRDTRd8.P-NBf/&.;99K7cT
AcMV@#;10W+4E&Y7/__W&PD4^KG:5a(>baZ?f20QGJ1BIDNgE)3cE_38]HG0YD,:
M3B7H#JBYKCBAV]\C<1aPS;(FeCWYNGE4ZdGP>Oc:7X81&P5EKV8+SYQP;RQSUd6
(>Kc>6]F,-AdTc1;Q5I<@>NDE<US@YOOc/Q<F&=e9)/CI,-]3R25Wdd+.YcDbPIf
=\a1=YX6<[KRcKAY.1ED&gE>=]SgNMT<:8[QFX,(bC-eA2E0OPDK^Bc_fYZMH[c2
_bf[_f]VH5YO[=3]b8Qd\Uff?8M,BR.8V#W2]GSK:F)\W/VD@PI9H.;O7F3W1(Rb
(\8PK]&L_UD0Dg)ZB^a_YfJ@4]3FYYGVL][EVEffCH9/H\33LW9/,[8V-?ZMgcVX
bdKABb(@Zc_cJdQb4)]5UHZbCZUBDR5dOe8FSY[a?NR<+JDD..6_b<DEb63)EMD4
BgA1S6@c:[>Bc2:?QR4=3RbW2-W,f[SQ^\@W[JIZ[b_Q1U8^>O[]X4]9g5626BXN
(&]d3STfI5TW8S<DC4.eaQAdfBF1cY75ESZ0_.O6&[(8(WDEFUI>WG-1/4H>-/BE
2UV]f\IPdGM-QICg.K34C25,Y\?]G0f-c+MZU+Q?(]FV5/MdF7a>(@:QHBBZ2Y3g
98S0]1,Z;+cNA;?L&a=8Ke&3.R-3(P1]E<^81T,9fNB6FO^7\9YM[TCa+-2gHaWB
/N@MKg_/LY#3S3>fUX=]gbLeK#6A,:MMNRC>?Z8WFC1@BVVG6cC+NNI.;^(DJ2H9
[6f6b7#[S)A:=YBJ7/)&CGI4O7KDL45;KCE-<g^V7W7Ac88\6_A/@DMRW-&W6#=:
eC&6QV+(>@a552gcACP+g@WbEJM&Y3CTaJ3>[cGB,HaD2a/:#fH^\SRN,:X0SJHT
e/ba]ZeUSOB4,B/P/]-J.?PgOD2DG[MDY+((NK]=:GUdK<OaG[4d@e;0Z-M?KBY4
3^Fa4_C[&)HKF[U;(CEB_[aN1@YT,DB8(/HKCXUV/2e(W?8E,D5KUM)GZ_aWCM.T
_=OR3J:IPY?[_>P&E-Ra[GHOefN/1@UQFR<ec9I>Z6W15Sa_#54VX46>6FVE5?cU
<H<^0bKePM>SYF\e:)/JGIW5J-F3.C2=I3FVKY(0Bd<=aVS8X@Da,C+Z3;TU(:e-
E\(VK]<4aECW=?bO2(K>W[N^X?]O^I<KXK8.SYSTX5=bGU6.;J/?+3EUHK>c+deN
:Qe>KFAd1JU0.OH8S.8&4#P<&8\4.cJN8f=2bLP9WGU;R&WVd6TG?O/L9O]8IABI
LDBgXC31B\)-F?3d8Z&N\#I9<?4Vg19&P,)US@AO2B#IX6]3W_^_6[@3VO#5[[L+
S1?/7>NfXd+JKCJ_+OR>K2Q>/0^\-e(ULe+=5<CK84EbN9@fVC@(JaO.W45J-?Rg
ZSY1HQ<Q8bb@1bg)E_8G[Y+RUaPQeR,FR1=5Wg(5_R(a]=<a2DQT]K<cZeU,92(c
>B4Y/<V#6B:YecGE/G;M[L?V-29IP84,\g5_AcB8M#F2LC<?-8a9=aNZMSQeOf1>
?Q)HAdG:O#)Og+f0#DP2L>IZf.O^NfJI4.V>)TK7.f#H<R1V\OSe<Z?Qc:YX+[N-
;T<MLMAD=Y&V:7^D;N(Q=0(ZR]4Je6/[>ZOB<NZ+?SZ-3@_231H8U@?_>S:4)/U\
dd5I<aGX(:?>\Z#Y=P#/PH2N66U\SQUHI0cX#F^7+Z9&JRc/[9-YI.A=64\DN]d[
)Y2FTD_333d<8>=-B7abT;A<DL-:B<>-@Q>D1WAM2LLJe9?E[]&_54[S3]^a20.?
OZ8)3gN\C,>,^dA.V((LZU7?BZ/?M57.&S5QB79[:MSfW+4AL+1VBB0OcXEE)LV)
V2A7;Z.J#@#c#Va:cV8g&8/@IKN&&6UXgO4KdHJ)G&&(a<^M5KKCO-bHe1[TY>1)
fQ;bM@C(DJg]Y,^O@PU9R/=VT8KAA^N6c&].AS9e\YBe/_(M:b8F(?f3JK6)YMA=
MTLd=+^?gO>Z3Y@=BUgHcS#U8e@(=2\V03b3Jg_2H.4ENM@C):.[aR\/.V\<e01E
bY5aQ)(9dDLKTNPG9f4&R/]OX,A^]5,Y[9daFcC[OG^^cbF_SW:#5eACbBY]R;,g
<.50:HP.gLGLcYL1Z7deC+NNY>-J\,KNR-ePA+H_3?BW_\V7O\OPL@?NgC0C(ZFU
6-d-OX@Gc-\^D^C[-5)&V3a8.)HI_f/2.a)@NKc1@0+?_(#O9B/N/MY=e7XH;KbD
\:+UX&650?BKV40_:^IP+EFFB:;0MN?Ug/L)\04Q=+Nga4SN++:cO>YBg20[cN4,
4D)K:TZA;;)F_#G0ER2FFIL#,..,=f.\ED([?d.K1C>WT@:Se9VD-g&;d.<DE(7M
?]Zf2CQLS1A]IM4d_314/MG@TcD<FX@SU0?^\S9RUCBE;4cH)Ye=d79AUJb+O-B2
aQGVQA^W=>G1dcBfX5;RN^d([(\87;D@5b\SEED<;SL/PXZ]9=&bd/gJ\@B(35J3
f78;(LZ-H5LUA3TW2DV5+)7WC.DC[I^MWA_,G5G=6I-#(OaU[LFdG2eFJJS5dSXC
SAHOg>99&]=(HK>UYQ[ccgaIGBM4C)#]UPI?K,[_b7f1TOUQ@0<-#(#fXRSb>aU7
a?JW&/1J)Q19NX,C-<PE8dLe)Q<Q;3L:;3a6PXQ8/291MD[U/J@[)_@;[VKML9(H
#DS@gUbOQ\Y6S7(7Cd&T\GH?YX2G-Mb]T6@Pg>9,[IF+O43XRE,([R4d)9Q),Zc&
\#Rf\]M\4@UG,@W1DBg@1Q56A2fB;a,d;SX_J;e/JL#UcF8b1#CIF/gW1#L/@583
\EO7L9O4>Y@+:8P?9g-2c-7#O8f7-\+YVR-EPC:N.7,RKC#9G_&;Z]U<fc:W-daH
,6+PgP1+F4Z-HL-8V8J^OC>NIfB9CW?EeY66[,3g8_+e6DY?NZfLBJJYZ?/)H-2K
=eL@3N01J^T_HMN2bMd0.27@DH<72C[-E8B2Z7=#23U36bEJ1&A?HM63##UH6.7T
I2@KE/E_KPS(M>LW]g(Z>NZW(,8R_g)aF&<K)O4JcgLT6^Z2\?^Y</V>E]gJ-9ON
g3cVX<d/@)]GCS3KADF96N-U.E&(LONP54eSRCdZCY)e[KT@OZ<Xc3QcMYQYY?N(
R)P](.+XU(4HXg?U;Hb69c)5=DKP?AJF3Rf93WV6^MRae+eOR;QX.&GDe.:+(#.T
8_0I.fYQPO(:3/,;dZJ=:GRf&VAC3C7><A:-DZ\K9K7;(EB#7>X10]XM;Y>]^)gE
#>VCY#a(.16<CKc4,0VCB==fJ1=dNPT\IY2ef=[#9g1(=7)FE=KZ@+56C^]e;_?e
/6[;<3+&&3X=9QL-59-OEX9LB&7E@^T5/1aHU;a;?U1.^^R=aVL8S?dZfT_WZ3F/
(M0->]g2OBe@MVL3KK+g](4(0Bc49@>Y&,aCML1ZN_2G4+]NT(@[#N2AX10-\^5M
VL6]#)f<T#>[fdTAP@[6f]]N0W;(C6?-1K5I2/S4/#@c&\2(R7\],d#8;.DWQ1_c
[]cWgfJ==]S(ELIe:EOa^cbL-8fJ1B483?^M.==SCONY^aB6FNV-8B?ZM,4V)^2B
C<a9)Fd6[>8A?/S8bIYTXZY:G3<9cO>KNDI>e3?A#;7I=?\3,R(cc-\#8E+UPJJO
PCC6Q=6OeXZ46HLaU2&dNbf^6/<]14X6AR(/+&[Wf:=N@DM-?[GD.BVHJS>UA+OW
&=ZQM8?(b@?HL\KC)#+8H+E;FC+8Y+X3[E.#IN3PZZNA74gV?,,)AcVBAEFK4YX,
(N<19J6J,&[^QBZDM:e1F__#)XXf:0;6I@cTDDfc4@N[<A;DcFCG2#d.5dF;KcEF
N#cDE\28=T&B#/6Cf4G?B][+0)g3EQ^,:g@ZPF_/K;-f5Pe)[BNNVEWK=97X]^]8
-3GFK9Q7@c=_-)=&5\]RDaD1.dP93#BDgYNFWAgdYS^d:+/(WNW:>^]g4c(AOB:^
WPBMOfFKT-SQW@Qg9^QL5Cff=&Rc>+GYB>&QcNMZ[dT5>3aDb8Tc=7-Sg2/O]I-W
ZJHSFRF^NL^=2#<>R#,N8d[[B_0Q52fISU+BV#\C]<)MYgQWDDe8[RFF,@fccdM1
92S&gVGDODL+IKC38WGIU+P2d(HTZSTLP:OJ9GW]W[XUR_ZXLPC(a#I/P-E9]S#L
/POC5R<0)9/+L_7XDOZ&#>@JXLF6U+&R(F#O59DG#^=+WP)>W00(-a^&7?eQD&/B
?41]DL,CPYLR9R^]#4aKI>EJaN#c\=Y9_@;6L4ZAPbK4AIC^;054.G?X?La]_OL-
RgV<Q/H[13/ZXM,/gM[5BZW.<P&3+f:EPS,<:RS3]AX6A7W3bBN:[[Xg4.S+-H(-
A&:7e0ML^D]RZ?@X=UC2XN:Y3+b?a54[a)c-C^[YI3\AHc2\W^YZZYd>N(K2)6c@
VTB@JdBY9Gd,ZAW>O&La6Ng7GW0W(Y7_fXWc7Z\5+cJ2+eFT9.;ZKTBg(Q/3H/YA
_7(,KRKbdUE^^[+Ib,.792<H]=XCcAa8@@I#.JW@37XX(b2g[ZMU:SO&^R=A#AH_
g<30d05e#645UgXH,[a[g)Z4&_PRX??XMO7H-4Pg6KA7W(J@\RL=d5dfRWIM@4b@
_45,?cGGWV#W[#.-4=W,C;?IKW-&_c@;cXTHO/c]Lc=4T8^.A.Q+:ab3eO;Dc]+e
>UUTgOC3T[/6?)A-YOf9?9XSW<Zb=C?6-^+.YF=+UCb<&OR3L;=[2EBfFeD3HD:6
:?HHbWU_&LHH2S\b09&R=:=/@ANW.1e<I[Hf,)ZV9Kc>fFBB,_IO\I33-HDNC^,9
:;2FNYKCIE1+BZ.=N/TK=YUe9^SR5Jg57YEVK\4CI:ca21@8S/a,28eE0-D]:2S\
<\,=3<Od?VB)N0gEM0;-:JQP6,]9WcYIF:P^)=]bKI^&_XOXMI,N9?-6CFZ1=W\8
a1L249f1B_?Y^@AG_917^R,4EcI-0W/Ma>e[;e9XOB()J<7S^=CYc/I(B@)U<@(A
+@:g,UVJ:J#H2V;:,UFAac4>8KcA7\ZC_EZ\L_(&3e(d2#P10bS3WL+P#aM/#^Xd
+S_Va7cVO+FJ.+e;O,WK,A2:dQY<GUI3G<&AX(B256_+\T-=6JQAKXHC:T,OC4Y5
fcM8U[851SQ><We;cYL^]F1=OX+I1.Ad1^GPYFB,EC]67D93E092U./Z9T:4@QP&
3BFXWRDAO]KJ8/>WA5ND^<:<7,VGTH_+RbOL<>\IW=64BI/4VE=&ITQ6[H)9]bag
-b]RE4+T@,70CC)ZPFgYW#/#8<-B01<-=Uf4YIWCATQ0/d0c8<cS<GRKHa@R-+^7
?258JEO.0.86f^O7B0PC86V=[#SU#;H,d(@/dJ\5BPKLba^?>BP;X8C_->e8>UNe
+@cA#BEc2MEV356DNWY\.?&6H-bOP6#RU(7@Lb7Y^]DJYZKf&a+8X_b-?:_;KO+J
UfUaH-#e600F/LQ&=]X-,+G5?cLANJ&e6^T4M4BE>1J;EJFB-.eMAD<bLG>;090f
-a;^MeaS99Y[/5;eK0OZcZ#<0dM@6,6bXNUU_:[DC@_b6_eFJ>3=K.YM-c)=E6[]
;WU4?^eRW,&&b:AK+:]fXHFIL(-NAaQ:HP&D#ORde=CK7O1VNH3?^)ZPgRR,5><e
12+-?Z<<cH-+@RE,7R[OL4.-7L\/@4Y?V(HN0INad47,YI]a>BS[EF\De7+f#&>(
#0H7OA3C>7YTDAE7>e^23dS^6dO,H5IN@Q0)H@B?YE;;6?XUgAa<GOb<;)a>H(W0
^HXY:Ge-2PTGQ77_FNg7aU\Bd#3PUcOYcPDe:9AVb[IA6)fDgeM,+8T&^eHO357b
E=g+dX&aX04J,]=99=?Vc<=.\2Q)PUV^(c(]&Q.0O4ENdXCSA<2)>ZOMQ:Q90I2C
/F&UeT8Q:MVEUS65-#,RX>^)2NSJE4d?f&e7)U<1N4LQO.LEC@@LY5Q993B0:JD7
0?=fK:^I3>-Z)\]JJR^)>+9\1-S7((-AB+_BU^K;(Q^Fa>354?7WA&J)IdE\8aKa
T34Y9)[A\FA-[0c+(RK6U)bLAKJ9>2[G[Df<e5;.Q:C(?MCRPM]Y[VY(\LPe_FfW
?;Y1&HR;^Z\DD[R&[:Eb8Xe/F0;=ON3XRK8D;I+QXSWS]U6XeVR)0bdE>J+);0WS
_I,dG4-K<V7,d4_<cG>,e899EF3:C]ReOL>E7TYH9Rg&)66dKK&BQdRL0Y-OO;/F
gBK3LG@4:Pa-^6B#V0(0IHd-:G>bOE2US4DPC2/aD[J0>e:Q];(:,W/#:FQVF+f&
c,]8;RPC@,X#)XgU]-e7a5eH7<eV56-G.V)(&DW.X_#=:>?NTXH&:/=O?HT@cUd4
\K6[62SeW;bP_FGNIV::>C^5/AH@KVOA5PNSN?WAL_2E^00OTE<@XR9/Q6]fI=<O
B6+.R=aC51bGcQS7d]P=-ULIX\IdGV:<+B05)@eGcAE8J>\S6^D^_2I7T[,@<X\D
JDK2?RX-^3d?945g,APCQRZPf[S@bAacM,6:+YR0fTbLMA8.Vag3[Q]T4e-13^SK
;)LEVWVBWOgK(bMA3MEc:Z@\Q>fFJP>G+#9&O66DDP]4<D[TA[9c<:S1?8PeAQZ_
dH1CP^_)c^:YEUM\,J9^2]I^)(DHDD8>#Y9L0agJ(JO>QSV^H=+3U\\-8&?@JSO0
W1K8Y1GWQ8^2e/@>U4aB=CGV:/)eP&_2/=G/31Gg#+XBIX7fW(UD@E,^)ZJ3c]<g
9<JJTg+_TA33?Q/G9)B4@)IWLA1fG+25d0)Q78/-BC31f7=F8@e\5@UH<58:6;9d
J6LU0:-[@2G12VJ/^5/&ALA=;cY_)C7[\7MA)KSZcQOEU5&?5@Jf6U4a-A,;AID6
)5S2bGQ9NTIVY:RW^AGDUGZY6KaB=fRDLC-3B#HUY8Jd:(,gFL&F4KgB4#=]C.&T
:-)b_[a\aWX+]<SW#ZabSL1e:)AJfIg_A[:)5Ha><^d-]\H.;HI[a?RU386@,[LW
\,P70ZeI4372X?P@(B@.b(]P_LUQSgK^C,;aSQ+7P3LX;A9VBKF7G2?GeVQEGT]g
MUNe1>F>(,W?9Y2;SZcQJO>=RaP0M2H/CI/U?J0J4VBB@&17)W41cPJH8;0P8BX(
4/4M3V+e;FV/bXOPdIM)(4KO93;(H1#_C(Qc]4XQ[F5;5g)O^_B@CMICZ;T:H4<C
#(<5DVZL;/BWM5RHK?(dU#HcV8^4.87V\]B\#G9RWGRI2(AfK;>V)&@8W8@2:Nc(
b@#(D,D0Q7O+#OTU8bg59ce+Z<O3</2/,>SW#1[@85O6.ZANc-\K?@A>C@7+7Rb#
R2@?&LD2#R4-0Ig5JZ17QML7A4\EZR;?A,_8_:=)dPJM>Z\]DGOBf63Z\=(K\8ee
VM2/d1#1:0V_OIgBO=Z)V6+2E@^6YIOIOd+bM)LW[61>O<YTQIDK:O<#<O?_Zb(+
JF3MPL97A/EdQ1ea>c]^^\W_FAg11#3&fCDD@K;ET6Wc?DeUg]&?EY-HWWaZ;8TS
)8g4T,MTEUM];6LQ]<AEC.9=N]T+-@cRGCc)RXHX+P(:P1dS&XfT.3C/4gRZ];QU
.bF\X-3J_.S)a1;,5(gMNV/YVXZ;-+ZK_cRUa?1IKTW1)&U@\&++VM2]YJN\RFDe
H8#Ia[+F6dYD,,F22LbYeL9^K,1fDA^+GeJ23D7-)LQ#NeDNcXD</?/KXe+2cF&7
DA4aXcFH+&?TZH+)T(,_6I;_JSB2f(IF[?b-2dGGSX=VLca0/9c+67U<2YVc[1>R
J9]dXKPJR<]@?A\^#SK?36B:[:NMFXaY-9TA7FWO7#//GTCOKRTYaJ>U--^MA<ZM
eDbCW2Y1U+<]JVS(:?,dVE5I_CVafg2/&]a:MW]PFQPTW.2)=f<1K\KTg_OHXH0[
M4bJ6V/V4ZNJ=W[LEZ=D##MbT:#1e(:.FR#b88[?LFT)T?8aU[?Q&MIM?FDd;ZX[
3CT-<GYVO-&=>UM/4BbNPNa3.P2#CK<b,WX41.a)]KHW<-;&fM-Y:4TWePU0dZW8
H?H7g34>\M9cVRYANHgXM\E&7JH:?,.S##;06F3<#NHME[=355[]84S=^fM:CV/U
?WNUOR,(Q76Y9IIYCCgO][Y6HBVdWAK60YZ+<BUW@eWb/_J,)XVL.OFR2V><R;_<
6_I<56MC0[(\F^?/T3egW8<]3L>).@4aWKHNa3Y2+9;6.PBL2)<X/#ZL7,5[<7b]
V+,-9KGS2B6V1ZV[\8?:E(dWI[-cV5;+aFY/K03ZFXA-D9VRC\a+G9?>6[#UTUgg
fQMePEZ2.L+8&:ZIKK05Qg049E&RW=Z7MfH7V\Z0]dd_\78]GWJd7V\0?B9@+b41
WMbU6,E(bY9>X?LXg1<<X>0N)aNBI.Wg&OUH&@e<Q10,W&[8XQWJ];^7U;PQ#Qa3
.(2J@=C-]@A/(1]U&a(QEVa7J#a9M-_)BO[/T<<.bH:U7,)XP)1,@+3F)V1Sa_CU
#<2P9Lc7M;JZ_>7c_,,Z5+J.GdLY)e#HVOE,Q84K-XEOI?0A?OKafP8+5b/6f2+L
ad#4GK#;X4A24<^/KLLd<d^cgfU[R^CQCJ,XJ:G-HbONa0NJM]aKe00VXI-fEIM=
PBM.8<]>E:IUGQQJKQ/U0W)b<[-QbINcb=dFQ(UW[fP83bF//#eGe;Y??O)8GF4_
R?#I+Z=dGBI^b\X5,>5,5_fZNV^_5OY6SBLdKD#ZHBH9,WU+&(^8AHUXKX[B^_8Y
gLgP4D=5caXP3f^(5I._>L]3;&0+bHN[TX/V,4)5HFdVACCRVC+U:eVM^^J;A-H3
T-&\/,1P=e84CB-\QMJ:+4H>3,4f)f]E3_6K1HT-[4bM,^dZI8;-ZE;0gNHS=^dC
=,<R>E=9f<WJ4gGX.1:(]X[+V[FFDZ:ZEdTc.S+3g/]]5L06f.D:&2;0J$
`endprotected

`endif // GUARD_SVT_AXI_PORT_MONITOR_DEF_COV_CALLBACK_SV

