
`ifdef CCI400_CHECKS_ENABLED

`ifndef GUARD_SVT_AXI_CCI400_VIP_CFG_SV
`define GUARD_SVT_AXI_CCI400_VIP_CFG_SV

//`include "svt_axi_defines.svi"
`include "svt_axi_cci400_vip_defines.svi"

/**
    System configuration class contains configuration information which is
    applicable across the entire AXI system. User can specify the system level
    configuration parameters through this class. User needs to provide the
    system configuration to the system subenv from the environment or the
    testcase. The system configuration mainly specifies: 
    - number of master & slave components in the system component
    - port configurations for master and slave components
    - virtual top level AXI interface 
    - address map 
    - timeout values
    .
 
  */
class svt_axi_cci400_vip_cfg extends svt_configuration;

`ifndef __SVDOC__
  typedef virtual svt_axi_cci400_config_if AXI_CCI400_CFG_IF;
`ifdef SVT_AXI_SVC_SINGLE_INTERFACE
  typedef virtual svt_axi_port_if        AXI_MASTER_IF;
  typedef virtual svt_axi_port_if        AXI_SLAVE_IF;
`else
  typedef virtual svt_axi_master_if        AXI_MASTER_IF;
  typedef virtual svt_axi_slave_if         AXI_SLAVE_IF;
`endif
`endif

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************


  // ****************************************************************************
  // Public Data
  // ****************************************************************************

   // Reset time Configuration Signals
   bit[4:0]   QOSOVERRIDE         ;// QOSOVERRIDE;
   bit[2:0]   BUFFERABLEOVERRIDE  ;// BUFFERABLEOVERRIDE;
   bit[2:0]   BARRIERTERMINATE    ;// BARRIERTERMINATE;
   bit[2:0]   BROADCASTCACHEMAINT ;// BROADCASTCACHEMAINT;
   bit[39:15] PERIPHBASE          ;// PERIPHBASE;
   bit[3:0]   ECOREVNUM           ;// ECOREVNUM;
   int        num_cycles_of_no_activity_after_reset = 3;

   // Common Control Registers
   bit[31:0] CCI400_REG_Control_Override	;
   bit[31:0] CCI400_REG_Speculation_Control	;
   bit[31:0] CCI400_REG_Secure_Access	        ;
   bit[31:0] CCI400_REG_Status       	        ;
   bit[31:0] CCI400_REG_Imprecise       	;
   bit[31:0] CCI400_REG_PerfMon_Control	        ;

   // Peripheral ID Registers;
   bit[31:0] CCI400_REG_Peripheral_ID0 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID1 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID2 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID3 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID4 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID5 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID6 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID7 	        ;

   // Component ID Registers;
   bit[31:0] CCI400_REG_Component_ID0 	        ;
   bit[31:0] CCI400_REG_Component_ID1 	        ;
   bit[31:0] CCI400_REG_Component_ID2 	        ;
   bit[31:0] CCI400_REG_Component_ID3 	        ;

   // Slave Interface 0 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s0	;
   bit[31:0] CCI400_REG_Shareable_Override_s0	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s0  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s0  ;
   bit[31:0] CCI400_REG_QoS_Control_s0          ;
   bit[31:0] CCI400_REG_Max_OT_s0               ;
   bit[31:0] CCI400_REG_Target_Latency_s0       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s0   ;
   bit[31:0] CCI400_REG_QoS_Range_s0            ;

   // Slave Interface 1 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s1	;
   bit[31:0] CCI400_REG_Shareable_Override_s1	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s1  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s1  ;
   bit[31:0] CCI400_REG_QoS_Control_s1          ;
   bit[31:0] CCI400_REG_Max_OT_s1               ;
   bit[31:0] CCI400_REG_Target_Latency_s1       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s1   ;
   bit[31:0] CCI400_REG_QoS_Range_s1            ;

   // Slave Interface 2 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s2	;
   bit[31:0] CCI400_REG_Shareable_Override_s2	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s2  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s2  ;
   bit[31:0] CCI400_REG_QoS_Control_s2          ;
   bit[31:0] CCI400_REG_Max_OT_s2               ;
   bit[31:0] CCI400_REG_Target_Latency_s2       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s2   ;
   bit[31:0] CCI400_REG_QoS_Range_s2            ;

   // Slave Interface 3 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s3	;
   bit[31:0] CCI400_REG_Shareable_Override_s3	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s3  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s3  ;
   bit[31:0] CCI400_REG_QoS_Control_s3          ;
   bit[31:0] CCI400_REG_Max_OT_s3               ;
   bit[31:0] CCI400_REG_Target_Latency_s3       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s3   ;
   bit[31:0] CCI400_REG_QoS_Range_s3            ;

   // Slave Interface 4 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s4	;
   bit[31:0] CCI400_REG_Shareable_Override_s4	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s4  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s4  ;
   bit[31:0] CCI400_REG_QoS_Control_s4          ;
   bit[31:0] CCI400_REG_Max_OT_s4               ;
   bit[31:0] CCI400_REG_Target_Latency_s4       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s4   ;
   bit[31:0] CCI400_REG_QoS_Range_s4            ;


   // Cycle Counters;
   bit[31:0] CCI400_REG_Cycle_Counter	        ;
   bit[31:0] CCI400_REG_Cycle_Control	        ;
   bit[31:0] CCI400_REG_Cycle_Overflow	        ;

   // Performance Counter Registers ;
   bit[31:0] CCI400_REG_Event_Sel_pc0	        ;
   bit[31:0] CCI400_REG_Event_Count_pc0	        ;
   bit[31:0] CCI400_REG_Event_Control_pc0	;
   bit[31:0] CCI400_REG_Event_Overflow_pc0	;
   bit[31:0] CCI400_REG_Event_Sel_pc1	        ;
   bit[31:0] CCI400_REG_Event_Count_pc1	        ;
   bit[31:0] CCI400_REG_Event_Control_pc1	;
   bit[31:0] CCI400_REG_Event_Overflow_pc1	;
   bit[31:0] CCI400_REG_Event_Sel_pc2	        ;
   bit[31:0] CCI400_REG_Event_Count_pc2	        ;
   bit[31:0] CCI400_REG_Event_Control_pc2	;
   bit[31:0] CCI400_REG_Event_Overflow_pc2	;
   bit[31:0] CCI400_REG_Event_Sel_pc3	        ;
   bit[31:0] CCI400_REG_Event_Count_pc3	        ;
   bit[31:0] CCI400_REG_Event_Control_pc3	;
   bit[31:0] CCI400_REG_Event_Overflow_pc3	;


  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
IYo6gAD3I+0z6bsfPlWraAVOIBlGsJQw/RA6nUbGqO4oT4ih0spQFKdSsSIPu5b1
QhZcgEikosgyVlfd5ZF2YcDWQddf55yfuL4O688eDviAUP0jkJVRb3SrLhxaYfPS
Gb7ntiK9rfUZWxxksj26ZslXEjNh7JkrvSy4nn1qzqU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 13434     )
VULzbDJqqiMfUHKwcm6qBMjoR2T2vshQtoG2/Na2vYTA1/lfaPR7U5EiVIL/dSNP
UUKyymNLZ3tfGt2/SSwfdMK+3ZOhEGjVPp2kKv2n8mSUKUt7Ug7WmeFwHAbcj9+Q
4KcS3W9jaSSCXhJWpUNND7wUz9IQc7S0m7hqwWsHA2Dch23PvGrjfSqbVM4w1bW6
jNlQ8p1ixO426HhWGfPVQEvzv5ssGFd8tNe9eTBKranR3SmcdTbdR5xDa7ZEhcBb
Xv1eVj0qRKZDpOB6oY1gElVjvzGIypERLhtWnr3RHz1TCpuVOo0iUeLgiYNKXNV+
2qIicDW5Q5Jp3LDb6wUxDdMlD6nVInrSSEYKB4jRZRKcN4n5d3PrHTvu97ezOX8o
pTaAANG5FkvDvVD0J1luoauwjHhBOI3J+19yvorXEfRFdH0OgoE0t5B5P+WtkFLx
NHFjpixN6J16x8eIBR07k++zp2QxhkA5ddIhm8GG5tvzQ6G1u0ZqhBtSnkS1Mi1b
t8HnRQA5aewi5HyCuzQ/ey6GFcFJYW1nq/A2vGFEj0RzjLLsM2SLhpblo6BlK5Qk
dmfT82s3GLaUv3w9VK8t3ZqseKkUd8kcEQsQYuHTNdKtFyOwSQwQsmJG+/ymxOim
fC83Ou0v6j8/fFdYrh9p35pQHtCAw7pZnL5bAJ4AxJ4WaP0/jIRz2BQErC7rFSNv
ADJKUwCRL8ZJCzccQmtWCd1bdnlZRWDie5xJMBTTCGFu9yE4Z4dr4exNYw7+2YMc
n4Co7ksyROBFP7/s2L3GuYmcNqEv96GhWelInPSgcIFdDT22mHmkCIjKyC7vT8vd
RQqP3a3WV+O+NdpdwyA9f0hS+rUgnTVbFWPN7FKQRzFA3F/lu25uSSLOjwVtfiX3
mre70tOmdmamZpcgGzT4kVSV1f3fTX8WLoITKhyhTIJLUfmkrTF5NuXP2TKHzwVj
pxqtVi/SymGTAR1rQzk4goaaKIbH8kB0p1BOMUaqExWKEiLockDksdx5jPr7WN49
horBIVsqxndyGXs/Fge1qnXZjExV19GamoibCEEhDYTeGCQOwu6qZqKHCMqbDW9r
CWrafnQPfM1NCzJ6VyZva1hLsNNs14jeMjgAMMsz2kMXaErdChQuNDs1WUGufxvZ
pIe7puZD7z7XIbHfWSzVt2feJWUn0AepDslfmHgg33vDsbObNL0OQIWV47RwT1bc
ZBVKanq4m3YHxQG8qBy8HNW/QyeX9NwhZ+geMR1zAknszK3Ov7pODKTS22RYC8E8
r7kgmEapkrGyw1iEZLa/ROmNdPxE029x5h9Bcc4aNoA+lGoWbrgBaai12lFc9yfo
9eqTgOTEFCFwCgfjLlIZeHAcqzO6JZE1IrUdoupZzJ7n0hbCUPy6KMGAqxw+j6/o
bLrf8c0Bv+YewLs1cLegjo9q5TIUzmvaD5YOXse3QstSy1xAbWoOXV+lTGkQCPKG
ZJ92kJf0VrNTOeZS0+eOr20Et9rJx1Ilow5zYf7gocBhGbBXlgw+N4PSWAhd92JI
r1c/rhhbGmwI1hwvt2HelBP/Bc2fvDSG4Z1Xoc8RstrEVPJBqni4Dj7DBe2mSAit
rI8lV+sp1lNSKveC9CxJscAlZ++vqKVCnh0G9j/v32RneKE4rD+gNLNB4keSSkhg
EqfM8HKbONWPB4p8qYmQ6mTFz5anSQMdwKfIso06pwcSYDMYLYNSODBSOFMi/BER
ffA46A7dkqAGnYhJTqxg4HpNche6LK6jeDmTUuJXHyi/l+q040XYPi6zVKRbCw9a
yhUnvT2x7ktoLQSDluT29vhxbKSKnCgE/+m6/CKXq1YtaoL7QZuclGDQMHINF6Gu
4/llgGBRpkQ+z9aTAt1y7SMs2MDUICzWVS5wB1u4TuyDpHzxSVO56EgOJfnq+TEL
zk2Kvh371IDC4ZXtpa196RzaQoxP0bvu7nd46XHU6yOqU/GlbYpISWaC0/suO9CY
iDyTNb8GT3ZnCTYUrnZc00/LlKUrfsi9ffRwMtCTRzujzfcdztJQ+MzlyasUVdMK
Jac5frTpf4p/hsEyK9DrQD0kdJ/Fe6+t2WBfaQRTpuK/aXj7U5rcaKTICiLCTvRh
eUxYzzUaWiPxmeFLw+YGPhDMfvKtnH4sXBrhYh1kCz6lDtXSkAb4vtz0/mExznv1
qav5pzxs3WCidNPp7UMGVoQWvtiRoTque1F2ja+Y/QeGP56sDiwBkNCpz4ps11yT
orKf+pQ8uWU7ItIBhPXqhlQLAypmKsNM062zZIwNzFZSOLtDy/huTRimi4hMHyF6
wZBm7OlARaBrb4gc9cYxF/cyvk2i6HpOPJlB0z7e6KFE8Mbk7p6Y3DHew+J88GqC
k4tGuQpS7pv+DG8w5WB199YIXCDBkb2SMdi5JuIT+mMFQkDGlIuJnQ/e0g8E/ND4
bzWSILEd2sW9BBsETWcOXtnbC+SMztJkNFJPgR3T6iphzVu8bo+1M/0NwPm3QuX+
5T9bvicWi62siQg1xclmr7EdkUVh5JykeRWZvdWi8BQSa4Y/w23zefbhWfjJamGA
4FlUoH82BzezM32yRaNYWWW6UiUUVqHqmTcMyTsIz2skPXrBhNnHwSt3bbhWHD3F
pqAyFiqJDP5YZxmB8RWNK1R4rs7pwGm9QLCoUIK6Y4XEFxmgxvFboak0tp4zSIaO
2hZKY/1hg4VIgMZZGLwdW0T3qzWRZThVUYg76En9tgCbXshZSQG6wfgy1Hl88aUa
dSUMfg3ESftMR+HasehmyKWrKn0FrT/d7F6x6QhKO30t0x/dh8UVwx9D+l/Lb1xh
gLWCX4CfAXr9WYlfyolvoybMJGvGNITUdUCAfZ3jfsUNWRlFW6J9I9dDKyqaxyDR
sn/5D+VAq/dkJU+DZVEuZrQwd0qQe9SahlfAS0529zeqqJh9AjbEbGhFvkbDYqEn
C5ppSF3+l2jWs43QpVjy3X1/IK5O7xVK3GzDTI2PaW4pq57C+Zf7zMElMhdFxhVd
7DFeBaae6tBF81AVpbiV/g4u8p9OWYFfKz20xCZYRqcoX5nyY8qosTCJ/2cNFEX8
24Mdoci4gHVajZI8fYjeaZdx7szRFeN6bnxN31Y9+PXzIcnLmExgdmL212GC5Py8
YDbItGVdP5R7kaWcrEL4Vsj2/YO6X/cgumy44TdScyEmk0lYRwuXbBLjKzK6v0yq
4Y11E3YroSyihTSPi74v4f2hfhBH58Rwx6n5yNDWvAoHZE1bc1kmXEcsgtILynwl
2niHxGDsbB6BPe73q78Ytd7Ls1obNjLNk95yD8DXZvz2Tj6N2KrlCxDexQJqOCSb
nHvH059v0d25Zsj7741XeXsY4BdN+68kbDJFcKAAaCDTMeLdAINCKafqzVjdjzTk
afVqxyOPu9QowRTti/R57keWy5Ur/O8/NZzGO6L57s4B5HgAT7YniGDurYTRZpqg
VJ00r9OUNm7hgr0ssuM2EtEd+gKu0XVJsvWDfI0N7JTFrF6sECeOgjv99Sy4YiHk
n9oZnZ++bCHAI/wAAp7RKp/5r4vQ6JrYW0fb2wEYGqwmp2aajmG0tjhgPohNcaOB
d/aiQ5d8uKWIOlNvITZqnbW2b/bevP5OvId1/xfg7kfJ+dUbSHTulAGzf9yHcnqM
Mx7DySZ4F597Ov6HS4V5GYANKusehRqnuc6mVWnxHp7eNQsvGjoG9EC3wZPDQ8vp
sbWWDFj3xSQJaefrhJnlZAY3ATn3dTPXrOGC2iYJKJI5EIWOjQgq3AWi3uMgDZfK
wUmVr/1ufl22dEW/SFMr3K1pRHcC7te37yR1IKcZWZOOHRYfO57EWBQ5WX6uKopY
SnwvHKtiOIFgUDs0G0lK/S6tsbHrFC1rjvmNKii7dIkVR3mamJL1WzYcLwSVemrW
/SpNJNgBvDU8zB6sw4+BJAGqmgtZhRW4rigvF+aOuUodSaBtSYOguq6OW59fbAbV
3VgxNBhm/d3MSPqPVA/H5yAOG0kxHgK5y8QgW0AuOgfhR7yk3K69AY9xVdkL+HcS
iaSKoqncEQDdaFkzBYltwD0juVC3SKXjZHEf37lnR4j/xzQizLrEC/ZPy+Oozp9q
EGL+8dBwJaEIAucU3sZkL1i3LCmhaTNYU0CLHYfrYDHJ+NmEQ6gcwCwcjBtGTxqU
2kDlMniBHFXf5ElmqKGdAs96Je8r/SrvJBEn8iuZdLdbd1hulyKYFSSlKYFHWxAd
LbRskQ2RnqMNDdrrzgiRAgLrnOaOJ6cIJTFb8Vu3WKgG0XIy6aRrtKQ8EEeSFJB7
LVVqrKrmvR5JiFY7VmElmmKEGccnCWU9OOCnpD0SFHI6cBE5duhT/wZdqlkYC8GZ
kq+W1FMkBhCLwvsAk5Qzg6sEl0+K3AiUveYMvNTf7QE+gtfgi2zC6ArX0Jd9bOw4
XQM/aesQH0e2YoDXM1H5cu4URI33jaAugT/6+3X1p6KdQklfoYvBIWJTsjTpc48e
DYiB5gdJ+Z38rCIImYIIRyO2zqXQC+eKR6l9NXfg8dkMQ1yxuwDl3sJ977Cep0S/
ViO2ftHhMD7RdxQkKO6r1K+NrWpZWlYOOImo45kIF/szwjB/ek8JLUsUEigRynmF
pQFxwtxj8lJx2Z1xNdQ4ppKlgJqVxckuaqz5Ufv8T1E9NY4NmRD/VyJZatXD8ml5
glSH1woM6FXDABRSvqodPmO1DY+jn+qIlj9tbNnFs0u86C7Aww0In6r+JQBn6jXy
a6iiRrcuOJiJswNam5EZqrxdQLqlBiMitGmnQ+AFFuEpp9jch/J/zK+wR6IsT0l2
l0Dkxc15vzSkzCwgjOu3ZBOER1L/n4FEKE3AZF6VuK/NmnEy8vzqBWDl/kNkdSCB
Z68ZCZi2vKLlbdL1HAEVm7gpejS6q0YmYgmbpGMVAZmiFjVqElXrXYyyq5A2sieF
Y4/H+sBwvOBrn1fcT3C/KjEpUOqAtHBkTCKe0BtReytEgchgQ1c7V8rDh/J0OzIG
G5cHDXGxQ5OvDoDl2WPJvoWUPuVaaQcGnNXLMDtPtwdlvrHHPA9JvR8zOUfm5j5l
kT/ALDPUdT5LFSKjfyg4gIfyAtUITXBp52ZpN9q5a5MWd9WTIbEf3Y74kRq6Rk91
YVJspQ0ach1rHmd6jPOaqLqWtLZgT4583zToP2EgMZyHSi6wI2qTj9dANmfzBOfc
poUMj97tCXp9Fc2nfs8cEWxCeDBI8grcNl0IeZfvKidd3GEyirrBqwBvRxmzCFuy
bx/376DYBdDq/8/03b322eco0BiZVDlGkVRbNQRnUOMgDxFbCAtG6bBxn7vwr/2B
MakWL6H8czbT0Lrvf0koFGSN8YbzvtetGGDHbxHHbvQ2Kxai+BTot8T6zZJ3/JPa
vQHKHz/BmxCfbTwUi7EWYaWFTZOncG1la/x7UgHGjIrcGp7aSwUvLUlT5jSlSZ0S
dtZG4QL+kricoHJFVx+ZN6vSLn+E60ng009bW0zcp+n2+p4Pj9RK4+LaO9X6DKv+
H0LaxWzPITWTvwycxorAc9FWW4+Cn8Y6JCJmTsApSv5BEjIh7/s/YIUSLKnn3TnX
LFV2JciguEYIa8RkPdA6yP3RO6hClf6t4e/s5j5lq8HneG8htBevAdT6Do9DHhMn
QNtnLXgLj7rQS6i0Fv0Wd0AibCeXAxstuPQ19TxlN6u08nRJbshdEam4N39fnqB9
Czj/I7O09Og2xxWm5cKNQLxm7Te5Wvh+bx71jAn+SVdIfrqw4T947FzkE2uQQ6iF
K/A5hrFKoL8wFDoSlk4C/pPMMqJeer3Li9+C0vchU+iZkt0KgoqaISw2Kb0WbN7s
31PY1EHj4tlOe9bVU+bhwo9cHbY/2rQq0HI1X/JNOaEmNhZeLpfXkeT6QoFUeKCX
OOF00G/fKI7SNepZbLuIB8t1FTIxGwbtpsPHpeCmpYqxAjVtNrLTNKec1jUsnyaD
zE+m7HsMzCZc9o2WDtQ3x55ZlvDO3WkV9CYU1EkjzBL+epaaV7TOsTj+/FFnFrUP
6jc2lDJPzDJMLuTnXue+vyStn6KRAp8Q/Q4DTnO4FlvK/oCfYIh2d+8uRdNiJhwn
olc9k+dBSSDnszVUaYj07qysVgFPfsixSz0rwta/9OrX8zFkeGMfA5iz8m6SCiYL
jBHxgJG2MQaMQ+SauSB7flphLf3KnaPF5a4BJqW4mi93MkzjCjCRchc2yiwK2pw+
VfiIdMymIXrwM34u6atYkggpk3mMHDECg217MRddW9/oiL4PrljNuxW5fBik4R0O
NbtFJ1G+PGmFpdKNca8aK5DfqH9ZOrA2o/8lDwwWT9pAFQXhcDey44sgz6Xc5She
b3IHH2AqE9kB9tNRMZ/xfMOrtgI2hW6S8UGJwtLYz8UIANtmNeSwLH9odZUsEs1q
akzgBcdJbumU4jx8Z23b34zrMyFkn4h2HA1cAsvQbFQ370S8VFwJKQaRV+awb22P
1J3ERH0nkyx8xAoKlZqX1kXUXJepko9MCo4JQY7N6+kHdNrHb9szqB/xGLsygETd
g43WqUEFOUDCV5bMWiRw7GmTIDrZHo1q7fAYEhrPgJDpqDr1uisOIJoHt3zpMpxB
r2uNUgSuokbipwSirObI6hOhTtRfiCAnLzHIUJj6NsxzeO2aFHcuV9atvdMa5j3Z
MtLc9CaQ8X44p95KQpjzToHZ3mqqmLpiQAECL0wbPylnhS2NC6QuRuXZwgMG9Mrc
GrzuZ+u6rIN6k+mmfbvGdO/ZMCnNkLJdeIOUtroi84HEbjT8odYOXqENvukDef+u
ts/hlwsjNLbITjg4GLXlpcoBQTiWDPMSwBRnDabVsSoW6mRxve42I8R0WZSIU0+j
uAf9gdXEcqeqRQuc7jO7deRyHoCjrUZr9XQ4HKxMLRJBZMAGQXvJIHm+Yk/R2o95
r4cjhP2vidm512zvc2hrtKu8Q3ZHcKEjWAtumkoRSdkRYzSqAUQ+vcZOMLRjVO7e
HJShnbCajL/LLkCH5cGPeYtdylh1n62QIMtSj8ZJ9OJRspmGCbY/58lnZN3Tyqbv
hSJjsHFZ+JDjNWlXu4n29PBLUhEJdf6mbTqKpeBO9hvuR+fklr3UmTyw5w//SG7h
HNy9/pJh6Glh7ei0ncf4kUhoEbLPQFHAyIr6DP6S/QPl0SXOAVe87ND2stZh9Rih
fVlDpHlFXc3BgBp5Kwj6baj/1VW3E0tEqGCL+zp84I+IGDx9RpbsI/TjL90wvQZT
j6jhCPrzCx7FBW0XxOEH9q9MDK6n2lKrUwcRb4dXxKY92XtNugNMgKXlusNmaTWg
4tvwwmktcgPEZBlwk9iXvHTIPJxfrhazRE2azmQ8WSzghtJnM90juwkMISXPLVE2
QTGFStjLENDE8JmI3QLLKgawnXyUvOOAHajepWf8uRUa4AdWpaVFnAkm6i94G8vg
b1WOlAh2roUHZoizOxTs/0mHY0GmcEGvVMGoDDetsEAuQJOjjodD0EDzG7vCYR0R
DrhY1I9oH3lm7n7Tzfo5Q+0PJMnlkNgfJnKFkVDezJy5cwPFLbZgqqXh0yl8Jr2a
keKvIG4y3TjyZRisNS0HO4aGTivAPa64EE9zANdihc577n2oRxPbKyz5QbYkiEGY
GNq3wIov5OaxUUkPTN/0qDYv2cACdaQpXkeiJdHPgrqTrBiGNCMqZcTxtwMflH5g
JvmCGpx8TuZveWJisRDYhFnnDiRdi+Efk5Wt872LVpFURwYylONCc9iap8SBCpHB
r8Wj0EVAnqzO6k8cv+nYKRq/BylNbOrMGWPqOwoO+GFY+4Zy53WyH5wAdBpLamHg
m74skmWh7p7CV7H5pOIFoY24hbZvTxCDWuKRgLPZYW0ldrWZ3iEuRfmGWm7eMuNo
6lOYV2VnVSDmZSCYQ4FxGtqEg7tJ7ATQ1Q7pWYpBPNzvtpgSPopoy98M10OE8iW+
8CkzNYEUG3HmSsektpr7cAMa5aqopjyDpqGXKtkEvcN/Zny/qNykr9CYGXUAc+vW
4MbmK5uZTiHa1UjMxgkC9J3shYNGUOj2nWx14wHrBpr3cSqNbpE6mN47D72DV3rc
1YwhTmDM/M9EWG+rjw4IgSJQWmrEAUf+MhfM2m3DUaNgu2jUtSeFRdgq6kuMSQ1C
wjgTM/vLfbyjd1uH7WQnQAXoujOOXKAOXYrVUO2kLi2Cw1NTsVxRiDkP8dKGvZWU
VX0oSwEOc3V6ogTKSERvOICQ6IR/7qDW7qGCJAsQvKgob5Jvd9iuYqJIdx2cUKj1
XKTXv3cIr7RMm3MOFgQvR3WzOOIlZKodE5DAi+/SUtPbzDUl0aoTzf4hz3LPPAQK
2PS/L6WIONqSFANKKJ70nT/6HtDUQdNr3jeb3o36bI11ecHv79F5KleNnoepLKVa
oyJcLeIFuuuLZqeGRTAKAQttlLWAtDpTSSkT0FmDAPUA+ndsfVC/thy30paXMhdr
+BnQH/uOU+zjxZqPMtiW+mn/iLrtdjVhjyFYpL/LY7hOiqiSfGFCgimk3LgtCQsP
9plKt/nsIoMpNWB0gQotdMkaNuuPiCRocyBOV4GyPen+uV606ZcsNnlZ9ayzd5uX
vb+/og0E8VsRrnlByICnaOP/S4G7/6iZ06g6kKZ029QoFT7X00m9BOW06261Mgwc
VbapZnL2oikmsKGd70TSbj1qJoTD3L+mIArN88O+E3y3Lc7xnUnwILba0sIDCDVZ
F+cSf8HxNxPwbK5NZ4sLnltgZDvS+DfvLQ+lUpvzxn1xppaZD3EReQwgUG65oNJc
ASwjVLxjBFTbbefutZ/yM4LQLG4Uh85XR8xg2eNdo5wWyq1Az6aHEyP19kuFy0d/
FYyxuI62zvGQyGPaRSvJuyPxhWdwLETTCDRgN/iPoGZt7f/dstP+fZl798rtupCn
sRGRl2/FxKv48ZH4n73u/K+EDQLnOkwjEbUqcBc3KX+w6yZnlmD146qgBblwS02E
OqnqJgShGzUSSR52sJSTWOUqcer95NnNVWxxkAimx0J3hzL/FKTSJmcoH58tr6Nc
pUjrXYMhJkRcz5ECiTTvM9JrOUnwLQNLOV+QLKpDX8h6zYy/HFpL39OPg1YacebQ
KO5WpcM1BcWm+KKZoD/zpWPwG/0UEUHwK0Z75xg3p+xWYlBA6201H7uhJ5xRsEa1
k5/LkaWgzghCXDxSSTmKhsjfpNrlY9a/nWw+EFWwTOMigtGkahraA3BuRLM4HmTO
Ti+yB3C6N/e1Vxj0VGN4ng24zvE8nBtc0KLT5IGYtKPixOBv4CsttAhDk0T9lzw5
soBfCZ7m6vypS2EQ+J/KeXQ3dcC+NjWyVQVQ+o0GAfzQNh/3VZAg/fiCDpu+hMvc
K9QBJYfCLcc+QE0wwMvRjOk4MgfwjzPY8vElpN0vMGtyh5+K8t/ew3uiC+3t3Gif
2Om4sVMpwxlaCeP7B2r6cECDJuSX9V+qyNolK/zeo3og0j7XdVkO/oRXTy/OEY+w
zXXvFIqW6TQUIZSsZnqtXMPovzZuSthvapQL+fUv4uzOuXp5XucLvpIyJycRhTsX
f+O0SveZS7gXIjwRLs5tOGM3tbn6ZrLJIpMCNk0UF5s3Qs1YSRbCFFylVazgyddO
B6ZGHhBDIPNYqt+7YTpwfuYpSQDVkR88gMpL9esZB1uHIASsIzVwSDmGuvx3h0uL
veVu+2GIJzpk7Xrq+1pmrN9CoWHoSiBgADVlMbtnrMVtRwWBHWbqvUv3IpYdHvDs
OybUDm85t8o6MZiFrdW1GHNNAH8A2A+30YnqZ81cHO9IRiEvxdIWd8L0CDGsDy6/
w/IyUGp0Pi+cieHA2AN/vl2cXOvwAwDBA3slFIUewpme7G9Uftx1IvjlBvM+cFcz
dAiOVaq81wqdMgMgAIC7C+YXw5TtrU8BiDq3rV9CbYxx53hrqC4jW015O6CPy4tN
SWYXjcv8Sz5Wd1otn0HTJEsINCEsBWPG82ERpNk3GhwlKdbliY+2aSAA+7KOuNhV
GwShULFmJLJCp79GC7dbZmMOSIq9DydC9MKOJMWvPvgeaGlHxYU25BIJx61PZJu7
8ECbgL4s6sR3YYzZfZ29WXLA36CIc2GEbyXNa44gRnxqgBWtqWS8OJhMggpdfhAc
QFtN5oLLdaMyeDeNh1BRkGHg1l/6O29UcMAPwIdDSN5Og8JI7O5wFLZBj+1ECgLb
6kr4tfMrBkGnU7AieM4HUFHDrXrfTvjkG3cOGmdla3pQXk4KWC/bMPKnY1OG6zmO
US+ZBvwsVmwVNdq2QhIvZ8f+ma+Bd2N6k1+4x4HpgY2CC8k36jt6UFyot8k+NA6B
6s1v6MH7AXGF55hGkepCZ0hfHs9sCoz+Wm7zKHKBldWEY+Aj3nmacF2p0rQ3/tez
Lt8MRYAx6uO+B4eclSCSNJ0LZfedQ8rmoUb2jRzK0aeIqVNr0Oe14HTSAYQM0wV1
dre5pzT6gmO2s5V4PUDK1J0fBX7F3OQyahvmHW6h5UOOgi1b78MKkds3angAnu2g
1kYDJYqOBBlEnVoV10dgEKV7gU6sCukm7YU6mRZ8SMtfxwYv1txCc6BJsfL0QUzW
AUlB6CVecxpEXd+PH4J9Qgd3sZH6O8eYXlTqv58bVLPpKKVmIr2Wbp8Mmu9xDDIr
YhQkLG+hW/PP1mQyYmHGHNqRPwfclmwaZ+dYenMdixB7hMOOtVuVqfJ9mdCeR1a1
b2QMIslEEKo5ByAUk2VALcMSODD0WOioyomo5o6z8K4k7HIcRi+iDXbYJfN5ggjY
HFXBcTmbLYE9gNSlAIdwC4gDD1mxUAb3juJ1rdwT0E6/eo8kikIM8JaGrpt9LZPf
qmXjNRtVI0yP/5xidZc5tN/zashb4O3tjvTM5KT2P1xuAa/TpNpqlf/B53imlUzS
1He255lfKWb7tO002gMqcTj028FiTbsqo6F9GoxdGwrPzy0e0tIt7FqekUyky27r
46fJWLcpJDXLXtPJyailWspZZoyv9oOMi1eKgx/lWgJbBNmW+cPUzSLYUpp07mP0
r+CA7bkucy6NlilZioyEIFV/kI23P7TZMzE4rZfrDi7YYLLMhdh3+YHy82vtIYSF
UUi6pplkFqsJ2Vq3MdTqX2/NgN1qgkiCM/sVw8h/f9Iot61rTxM/RGtKN2szYniM
kYe2d9eNDk5BvBYp7XAbAJY4FX7nA6BSEYdOqFl5PIPoBAaO6XduIdRvLI74FSOR
H2/lV9nNlbwYIQWMJwSUwfpQp6VKFNXhns58NafX9bMeoAu99vM9d5YjUwAJPYmb
qrlr3+WnSsDqrgt7K6bxYoaZwTMtAxPjAFXULBljGRjhlBm5wUoB1ZhtTskAeaR1
3krGZTi+42FQ7Mq7/ZBF4gnKQvIngJ5CeA0T/KHrDSr3ijUHVLk696jRqaZGRDF5
ZCU/EmJltTGMoq+AH4woGVKCb8wWX8fi5sEyRAsnzaKsIjt6OyBXv8dLYNY0xbHs
VA/7iybixdakS4co/Cv/QWXOCfkL1zjLHKmv/uPSjPiYs6pmK7ZMFuiJixNF7HOy
vVJm/HJSW104/G/V0I8Gwf1oIG+u0BsNCKX3UejUqIGIrDggz0f9VHXurzw7mrh4
8iqFm5UhvsZfP0ocxTD3UNdZemgx7Cd4WCeAdUE2IEY1XqqMJmJUaLtcpo3ZehCP
Aa1FU4a2i88VMgHjbS5f77NtrNsRjbF8B3fh/8s14XOYoyZfJ46JqZmW0cOzPHt2
jDKOrwn3EmV/SQyNAv/rF/JVmFDI2ZgDD6ZVL+yHEAGXgpcxNCqdCQV3uM9n1R1Z
s7F6ZbRBNg4Zoxc+exgX9rLNI1MNoFxvv+K93YklWozBeGXNZ4gUvPWpRdlM7BBJ
XnuIjtUyR2ioaPORysZKw9Tk+gMuoExWMo8k7nazf6OX9hr7488Bnz/0gM1byqJa
cGwA/0a9dJ/qbQm2ljYQzwaSHzS1UuaD9uFJuD8OF3e88+T1BxYNhjkJKcwGSpdG
PHYX0rcg44MNGzmK9oXipuVc71obHtdm9erDFPDMmZX+M5Mfhb0MqRWvYV4dS23I
n3NREkoxoVvQd4DVP3k2we0LDYXAI9LzxdaLuEGuvtCIwK5HkIGwtHU7L4g0L44K
HRO47QEJj2t6qQNHNLuAPyki2vO3nCOC2uYAP7qXJOz+VcbIcXTm9RiXJPibXd7l
AQQR8YNogdH22LB3j/UP2uWylGR2c81y0oSyZA4tx5ceyw295Qe+qKfEA5iIe8z1
A06Na/udRx9jl1fFfIfePpb1u8hj+yKxdUp5pwhoePMw9i0Dhb085pF1wp8IgEQA
5sMUQ4nvdCR26i6Xk6orXZrSmYPh3CqlBVrjQyq120JH+wXWoUff8moyiQkUCO3w
tD4u2xxtA1WlFZMTMG7Aq81gA2QgPZUP2HBeCUdb9Md4U1JhO5JFjxiBl3zcSwXM
V8br0wRaJFuAI/SUPCUGHGkHBaq483NcNUDQUp9VlT1K74bGDo38rXGHRdFZ81UY
gessS1+7xuB5JxUueNr9slEf9VhF/e+ERoApz5jO7vrY+XRqtwwMj1eLIAc2TUW+
82nYBNS/fB6GzfoBIolzxagqoeKDzQANuKiVPYWAa6EKqBtme92jL/p503kZBthn
9l+GXqnfS842oHlCiI7KxHBchDDQKQUnpBxjt/HERCzfEkR7SMpLfj2HOZqwl5qW
2i5/B5IgTb0v82v4Ngjw6Oam/9fTcRcV5ixmBmx4sit2/sO9WaHfWDHTwGZXVWOj
ru04Ag6u7fIB7vj1d7mCON3fmX7MyzJgVGz/NfF1lWWtu+Af7n/A+TL2k9Je6QF6
JFC1MrmW6Db32h3J5BpMdkkI7/9wZRk8sqpSqolnaj/FyrHJg3fZi4OcunApmimn
1ukyFzs1MB9vlbu86FpHKUesn6T1OyM0G+RoT5TJ4S7TtB2+Xy2DrvmpRr1OSODL
orlOdVYPjjK358nDxiQeMmvTFDIicQ9bqFiDld+m2tVyrOk+07bq+Je2ahfmsbm/
kByKA9VQt/bHyPnklDu1e9dEjCDFEonAeuVX4HZbWKLVdEB0Jib2iiJH+lm8rV+C
t6AzQS/7jAay0vQ6wDehzDc6t6mX2bRha1uiEaTByIbDk6LurUF37YOEINfjGrWf
8idNlAsMvk1MO/Y85ZLvccFt+PLssJaxBt0PEcVxB7rdIiWPqqpjbgT4qgYHlAp3
Hlze7aQPT/clBmZg14biz4x45MsX0lsPOFDRNhSD9t7joffTy67eP4H50WqnfGUP
uVj6EOEGMlSpUnf1nrEV3z7PBtys0CoYLrn7/5DTnkrHPHatLUa+vzX3iD05dU0E
UTtYOU/w2YIm7WKW2Cutl5GSib8LULoxdjQ+eoLWmL4BY3CnopPgXCcgujpu4/Yp
kRPzXLVOMg2lRAkwD27HGwnMyG0c/zBOf9LYY12tv8QzxO/Ul/4PYfiD/yBJAIwG
m4CDHq1txAfTbsJzFdrVkt/fh3psLfEz5repmFUvoKBnpHw0ydpP6ENNveWZ/CL5
rmp6t+rqJqaYV/g6Zk/ZOuQAF1dRsfyz+l7yFaXnPUV3aD3zJz60ky+qQVBRfno/
zB0SroOW7urGVn7/jUkco6k0RocMCVyr5OXBenJbZPNfkx0Tj2eqLAzy1Tui80g1
c3sfD8AaWcJi1vEZPg0HuQWWy1KDBwGx4r9HO6PgXzGsF6s1+YXuP4o26ccIrQxD
Ee+deryrg3cUN1QyoPASPQGp265bVKLSUCjkTdvLvwkA2WSmz+oWfAGyXT29U8O2
BrP+xOxup4RFLEPGHEa2IlFBZ8yikqLtQG5ZaeXGgZ2OW+wvlmahQ/wofSXBapih
NqBjV5G4wsGBrkrZXps0naNZ7O9B39x4KrfHUkMFWED7YNAXBb1P1KGQ3TkPppiQ
OF9rmiAOrjYPbcXBhswecMi+KiTnkTzgZo4+2eJEfdsB6CbyE0zrpzDhYelkl3v2
TRQ2mjPSYS3yHRqj1WbfxWVfE6O2JJeJFRh246mQvJa/r/ndRH/tYG/kYaJKpxVB
qdMQAFDKUA0qvamd3WxdRufuJ5hdtiunMpUUUC2jWVdIQOZT9NTVZF1SLHBRcw80
tFSUWW3tA+7lWwQ4ZiKvEUcZGo9bhl97WlemYlaF3u1/j8bwxHw0sK/lBN08Nngv
JkmNSyDjjCkcTcMRkqWqQeEnxrrUxrIsovzaks8PImzmKjnNLbKDtrswlpOW4cCy
04e2WjuYWcOahRShi6VNL0/6PSwYBlyTM3+2/1OIoUH+f7AyzJ7DuIUvgcQqFd25
imGpM6+ZhQfpczVWgzTz8m+ncM9muHr1E4po94xk+mpCd/a9MzVjSiUpCuRu5NPQ
mWLUSFCFBv7YgKjMLFbOxnYqt4nFx4xpFd2j5F77NQuQ0Jblrzziwc43BCxAR9mx
/nig0ERffpokekz8hjdBrH+4cs+0+Avp0AQ7Fpye8AkuG3HMoZnPUnoaB4V1CNdm
ETXkR1L3X202dpaN3TD9ID9TfbMUFuhXFfpFqjGSR+nkFDpfbsD/unn/vv3KZ46r
/tA0cWdCl0fKpeBwPrqjWO6o5g1WH51rxmMck5OeSETPxIweByCq0VQ//eMX+X0A
Z9QcmRH9E/YdKHZIhz3TczVSGu2biQJUU8CzUiZTC36pem/I4i2ATheMd4XKy9nA
r8UBMO/SkTHDeDuPlz6TsE1fX41r0PTBeKb7UirasXAcd4DFpeOQGX3DPcZgKtxe
zV+7vLq6THJxSt+MxTH7M8ay6fx0xgKrmaKT00/PGxuXwgp3nfIAwmIMu/1QFIHC
lE7b8JRl+aEAn6t+mOANuPlbRF7mhUtsedKwDG2zb4an3skuaMsf9VBCyp5AiYtG
j0SHvhUqcRKh6ya+ZZPUOB4sy3IQbS1dsYWPUCMpde+rcSK0NQCILPbs0TStGOm2
IVCfHMJTg1taliZ0l54lripTXSpjdTkWXk8cMrzFWFqGr2q7c41QU3XqenV1tnCL
53TEpX+Erw5cU3GG5x0/DmtW6FwW2mc2Pa3rA/KpapDTfOYeG7OqEjS1RoFKjxXX
63sFeCfU4487EqRJ2JTv6hFaF2YMmZWBaIfatr1VGu/zs35HNAPa5LLgcV8+key+
NkT0cFBC6Pbct9PJ+VWB58pFQJEkdbB0XTtqp0uIr4ytpuSLEKEjHoO+xq5/ErJT
dCmzbAQWzySfC/i5OzuOm/PqmVo2KW9KVIaY7LezmDWnz+tV0eNqvRruj/jb/inS
CdnevOUdaLBMwpAhh7il0HT7bbPD560+aVrVnKLbELeEDKt5jKzLWQ9B0u3iDGSY
xxIfEoDD9FvaA62C2/YKsD4TjZcd3PML1/u11Ywg+COjwf2DpeB7rKn4iP1iSBIw
QVNV5jEc/mkz6ylR/Al8Br4jFxKUhropV8PY8htWHhEXSYhk8l4/hEIqwik1rhCa
myHzrBVY8Sesk1ij6cCzwOCt4jtUxgV+IkB7Wg2UBaBgHJVxiajnnCfcO+cItl4y
sj2mplBFjLEA7R1sWFZUNcXFE5WYz90BV7V/nXbQKHrwbfE69u/x7Mb8AE63Iexb
bM0cVxEnEJZirauBaSRLCKyPbmLR0ug8oKm/OSu7q+zb4SsamNNbtbc+qsQ0Kxu9
OQLmfJD1/GNFecEGVt/iC8W3ZMAA6lTt5fq67mwrO6/0A+4tQa8lltS5kc0yedLf
v6CsOVADp6emur5q4GQJiVLvrWNXVyWvA/s8bVeTDU/FDtC5Zu+9s82vJF3QF9Ip
ArY0RtAx7pcFrSIPzT2p9+j2q0PGX7ejdBocfhVGEIiJyC3GzWS3wraSzGx8EgJ/
EKDSas9QBXKRXLF/NRq9Nh7XHXk0Eso0Eq+O9hQBtDcqoFdFondg+/5uDhnYhaD7
vmjUWMFhU8SzVNxPS4LURtSef6OPTfR930Eu0Br53G6YPM6JECkJtFF5I1a1lO1E
ak3OlV3o9nKm50gQt6GD0x4CkZ6/w/aX+P7ZspNKJ9w1Y9cD8o7SdLoPbw0cX1Ah
qku3RL0p8LApVE1HOO1fx1dIKZ8svmnxraN+ieB/ckLFsh9F2kq6GJIZaUrC8WFw
4NgoCvjwhHzxJtzFFHyWP2CtlYjyGujNTwTsVxMJGQ3OdQpMA6+JTbPlr+aOISmx
VGCRtDyJ2oSNPGD6ipm1Y4kkwrzTgIsFSyW7OjE+9fRP2jFwUYX6AaAjLlRhAisk
F0aXuoN7h/AabDZ1Z8tiar7RMIp+oWhD77GzFfSfF+73TKwm80C+ydbG9eCkNbrw
gN4AJLsEysRns81jbJceAHIldZ/IbC56Wly39WKVj8VPGa0oTK2OaYToXHcy/9lc
zbvIqXhToemOPjmoSBYgaXXnHcU4UAk44GktumgilvF2M4KRlVk1ldbJKejLDuc4
iXrEBmhvDtO/+LU4GGSJtxW4T82G9SATD49FPMHtAWnsfMW+iWqMO0GN1M19P1dr
hIqYQ1Dt7Qegrnt5UhEaV07ACeZVHw6+Tfxlnt6YIKrEen1liZ+qbYmNCJzmmMSK
gtgMhKKuyhDRBLBU6AVPibLn6dFWpTadjIs/Bp1mUcKXpGYJBglxztRL6KL+cC5r
yEgJITIAmGpKyXpkKMZgcMP3JmrvZRemQqLm5MvCePBsOcujjBTdwaqx1XPYTDI3
a9TU4feg/sG438azk+GWO0XS9LGtIaA0EzQZ9THQfJWK+ZuPHescU9J47FMPNZIG
lBPyRp85J1UXl/5vZm9+TuUeN0JNmelKTZ7zxCBm7/o9grmVsvhdF4O0DqO53xJe
wrFf66N9QpeWxJFlNyaGxDM05fjFHyFJND4KMe9zYeuOGYgg8EPqgThNR9RuyLwd
uZLoWr5IY9jTSh3gly8yNcsTyh2H16XCIwAIUjbUYdzfiZ+WoetsM7iGlLITf4g4
FtlqvzJjNVVbq9h4l9EeQ/nqy0PpqBjwGP2jfulz9P5HUPkDE6S/wEsWpC+8rmoZ
JmHI0SSFXhQAGkNVDa/sCC7Hcv2utW6f6R1Ut9Yd7K14gmnzaklX1Zd59jFNXmbO
7/GbOYl7JRdks7/9xq/7yMTYE+l2JpvpwLTjEK0o0NcRwgE6MFDzyqfeBWYOrtjI
sm+g5DBPbZwsnT7YoVeSyCtEHgo+rd4mhorZcpnl6/GaV4SM1e06YM+tmes4FXGR
inr0ypeYFJKi4oqmiQ/AMr/KtO2A8uYOe7vmFY33Bv07o+dD8nJa1s/EUR2j4OK1
APByhjJR2jdasx1/fDyFedUpx00qDwrqogkieEQyBIpCOw2FBmhGZo3nUrHeHdCz
bhSQlHX4IBs0MEB2thM8v3/4USOXcg3LU9RhxdmHPTdbaZh1P4HC3qUfv/KMlAmR
1imzJ7zWLCINo/V6WqnWIeHzgTtU8Voel3O0Ptzbpp0Q39M2bx/nX3Lj8+6j/H/6
L2J4rVhjc1nJhgye4Z82J04lKWHmiRYycZOaPpxVVzxx8cjOMZp9Yxk37fZWN4Bs
kXC/a5v/QeSOfQg6DrIRsUxfidVjqHmqXYflAc3+1tQwIvfBlpZEPGI9VCMI2yL6
YKZISK6Yqw/AVBvTWLEU8A+6r99tH+x+HIAo46xpVf1dVorHw7F0q5dp0pjjdPAO
cepZq9KU1HkV6nfCmVldox7ym59Mud+m2TcyEfrMv6SYlao5hpAInSQje/0ecMt4
z6PJd9zHX7Y3zoAP9Vg9sDaIRpyCftyFsW5L2WOfszSQ/DH5YcPCPS/NF3lt3PeI
x1s6WTNjy5YY5C4P9lz2omvmZq0mejxnIn2chneYKWSe9JVVETJcEGUdVtfby0gD
q9AkY6WUmWrTwXK5NN3cpDldwcM41pLK+jKKJ2DZAxpf8ZnuIoKBw9J0DLz0kTZg
9mL73UBYGwJFKahuH3GURkSQMNIIKEF4uBEZ8GdFI0ytfcIuVXQaAScnLdLWChgn
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ZVV8ktB1lbG3FaV8lw7jGl9KR9Tx3ZuRlVvxirMa3UV4Irj/dhgr5qOsImMWLt4N
zTrTSToZhzvwxFuU6cpOfMyovkD7E/ArAcpI4R8iyPEIsb/Wnr/fVak/7Gpf41C6
2okLw/cf0hM2L6AI1xVTDsOwkBC+4QEFGZGmpPQU0j0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 13931     )
aPhK5XtiDyvnq2WrDz1z+pfvqW5K0UAtXE/B3YhlLDBmQJQyL18rB3MR7tUbPv66
8lYtNFoK8dK6A7++3lMoO8Oz6eqyYD7TRbttIdOuCgghdUESlw0rmpSkCzHTE1+C
ZIZxGtBihdR6khUup+xQq1TAwE1VY2SZzEMVj9xpDT1K6Gq6ygDDs0YyiWzkCWKf
/qwhKQKCoEz71knLfC8/Fw0loZAToOvHoGLkD2rJpzgs/Vgz9hGIqmuzBdGUtroW
PXmBEZwZXxnH+EGT5iQgjRdkwhgXwPpqiFGrtNCOHkMzSXD8cEktEfS/gy+oCWJH
4xY0ajMcp2naf/Pt2lw4l53brioxaNszAT9JUEwr3bFGXCzlJJ0r2oqKEQx5hotF
e/sju7b5EtZ5EhA7gbRiquHkO6L0TJzudQTePtUHju6qrdTLP3vG+zmg3YiE0QPd
3sxnTTpoxvxUpEf6r3W9sPpmbQJHDDdXkgLSWTI53fQ6JOp+n8la9qVZt0xhRe1T
Ls/Xqd0HX9SKM57OdCevLwQlftsUL3GegmDxjeJI/30aPTAZA30tVRSlKiGiVJgm
VCFD5z+FMECCkBU4d2Y0pheLz4wrpDMOh0PJo8tlpgxCp9xsv5AZbP8btSmeotKK
h8CI49JOr0b4xxL08QIYTAIgtY9m9fC/Xa1OIlTC1nQ=
`pragma protect end_protected

//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
IyirNbQDFwxvO48Tbm5KMp9XAHvdA2+J2wQpQWinlf+nTarwVENYuQdsbQGzsqe9
jbsVuWTaPkH8OZ62AvUrNTD9+yJqVX606JmXMVAxLFobB+djC3oHr81KxR7PXI7w
WYwEDjwodedP9RT7fUYjOczQJXkVMaUQdapR+ZIn0zY=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 82355     )
HLWbFi1XxwwBmVTg4lDnenBf8ixYF8IaAYXpeEzdVc+9ANFvGrBTSGrM/RF6slSU
gWiaSh4tmTjP8k+dkJtwoHX+AF8bn4wmWu45R+3Bb7biLLfY4VFBSOl/5+RwTcAO
Dm7zIoMpzz8DaHC7lukQlUdPVp34y4v4WRGdvnLgiI4xPKngoNMBSG+Uwj+h+bWq
Va1Z3seht9S8tPup9oeD1iQNU/yMGbsqzt+YwnMMoo5j3TlvCs+D7LLNg8NtqFU2
8d4vzrKSlMzYAIQMVmG6anux31MaOM5CjBcjFUCNjXUyxmhZRufuAlzDJKe7s1fQ
2tP6d78va9/XH4/QPN0l+2Xw5Oi5fun63eBwRC2A973ZPQ/8nDYZcabunhtpDDYh
VRzqYBj1tNVyaTwI46o67A6ejOYlsaU4c2fARwmxQ0JRS63/zCQUEFSB8eIol55X
rjAKAewjuWg3Y7mNCqKSHLRfw7o56SExq62wuxI5giPCvg2/IwQ3XV52reJV24wj
CzBwCGo2A7fPVokKBHMAbXm/OeTOT+Oe1pHgoMTyCzR3f+31Ol0tij7C0RaNd5Cd
nn/taMcwUGa44Kc+P2/mBhvgWypksDsSomW3Azqhaaqjmry89JMRJDWzAIw9Qe9e
gUBQUTpFLeSopwi0uEfDPFnEtOIsvVP68LS0s6IotTNowRpR1vE8Mm+CfCWr4Sjh
RLHNxv+kA58e5pEsglaQ6QII7X+XP6WvAT+8v38U1ITqu+lXv2LhSuHrRJRUWDAQ
wz1C9JNq2CUDEMSzr2xV4H3n8vbTj9b3B2vhjPybRo77aIXxxwfKy9CUTekZ9GTe
aBggLNrXEfc6Qb/3OFHXqJlUNs3xnfVVopMMhQELKOuKTawQHQodlyx6ZmZoS9z2
bR/gPb7/SnG1iUhDLvXm0yeOs8ZuLQcDlu7DgVK2+hfzJVJ3IWrakfMv+3Ai+mDs
QBSrxv3NzgF8aK0YrLx6WS2ucJUUSAMLLylBSYN54gWmRxG0Qy6x2XQxwn18t28V
ztmBKL+0obu2fTa3OxLvoQodm8IMLhMlGKUAxK2NVRBw/Hk0dX8oqpoPVt/kbwji
mmp75xRxiGWTWHE1YcoN08c8RidS2zXv1XEi0J+xpNXoBakIgZCXLCj/paUJsPiD
b+lHJcbG45GEvY3YEzd8EycZu8rDpt7UifW3yfiJy1/BRO3S4LdaMyZQRrOPJNB+
uMbGpDIZ4+apiOMqblCWComejF50cor0+Gq8beLfAlJ86KOoNct/m6P9bKc+W/jI
Sh+Pf/ov0UEkkviSUQo9Y17Y7zVZx9jZ31fQbWEtOmh8AgkXY5DiwIiDMTdaNVll
pyfTWHrfS5p9pKgUC3DQf45pzN4ghCGBVopWwQfSCRAmLxlJV+RELzkb6DcLItaC
qinLM8EdgM8Cx5DGHyCp2Lj8hl+ez0KRr36EXsciYMBnPkKDmdNLtIiiuq9px1ll
qAGmyOTpYi9Wb+Q5G5hztYGW6Bbz6ltKMxd46Kwn5rt/tQGwyYpFt/DZ/Lc8Bp6T
or4bMDPFBP3uGo9sId4G6cD1IEnWEQNt2VXHaX0EqdMsNT17fXboyBFZG5jnKml4
3qtCDg/jdXrNav6A+HPNbOnpFbQC3XLY2LMjIy5GKi8bzFkBRNTaUQQbpMSuuJq5
Z1Gm3jK9hnW/1eHvRDUbdmy9vxjXVMFkDrKVVSNTn5Sv0bL5PdiFZhQldPr7epCn
4sWCi0cppBanM0jm9jV8E41w6/I2jyiB6YH+hXtfenrehKgdWwSbspexVjjcHEBh
ziaKCaLeZHN7T+OQgw2q2fy7pWfnO/FiI0Te26EmU6PLizSIoAnFNe4eUuzcj07F
AKmlTVPqOgcH917Q0w2Qbf8Q/uEXRukxbs7Kp3W3u8Efg4DUWIOi5ZkX631dcN8c
p9+CM0bbsoey7Db8Xc/n3fHEqoWG9oeSRpn4aGpFLHEbZ8IliSPVwH3sOM1EhjXO
hAiCFIV4QrG3F35uOnjRHrajyuHrcrOm3kzxBhSKIjOFg2roPFJelPTQ5hqljcL5
KddvtliJBEnex5bEhZdDEp8e9WSQKL9p9DVOeWMly58u+ya/tlY/PEUHiDQw4xsE
hr4JjdLP5lsXvSkm/eIAQyvr3oXvG/ZaVBONIvjZUVPajA/aJmvETXXKxPTRR2CG
ztwg7gNLnRSl1+SmzWIo3Zx87Wie8OY8byqcc42mcBlOk1RP7e+8jHSZGu5ZKSVr
jlaKfwxrMrXXBhXs/w9yvnrLJ951NQABgFFdZLU7IEn62GHIImCHtstTOhs+WDho
nJDByJb9erGatTiTH4Hfzs1EH6OLqvQ51W5mBey5IJL7hG63x6TGXrsZVcEe6rEk
rQf6pOvo1ZSvdYGxIEfazWdtvnn/u8Hjv9rdaeKpHMFQlYiFvapoBNdF+dKv2jvs
bgkSOSvdXCFjDCU4wYNyu59CU8v32CTa1+P12kcpmHaxHZ5UffRaTrE24AzRYzol
d9Q9W/EyEi50a3spnh4vlGCbjq7LuCIOkpFWhFKHDIcDMQfWgfxsJRXGs2okitXh
5AEgY3CjkVbq13dij+LC63OOPb7WPd5yxtYMv0BgrsD3jGWwad/pBEitMFNrk7ah
SDgggdNJQjbeLR0bGbK1nxuP7MfbHlk2Le+bWaIIuF+tm3/OQH41BkYfD1TArfZk
rG6DXiqRJIShI3mXrA5xrXQSTQ069KsVe707ImELykNUFPJtNJbxAPKuteb/lECl
Sd3SYfREWMUEQN2LjYGTASN5/yKSZ3/Gzkl7j35hlE1LpWb+ZPRQoXHAS4pyHdCr
pp/n3Nf6Gt/sMsXitNqA7idB9Vx9Zu0XnwRwuwzfD00IYyrCc4YUX+x5zJqiHq/R
gg8uJUKCp8TLsrh/BD/uDd5v9etVVyQOINuN2hcaJ5rQHioZsdrXRRBsRoyGqiYm
s56UwUaYRDabZTHxH0cSt8IuXYoElUahl6BDmRZpVguXTTeQVJVR03XtTAURzmkv
qKsTTve1r+8P20NQyUbTiEfKSIv7KTSOJwvIyOvicJMbbq7Yq5rHu26ZGm6B8Si7
aMNN1Zwg8ZarHu2NZIcImeDp4CGank4uGqIRk3cXANUyB7r2rMhdQe3EdnkxC88S
I9Sd6RZWIsOPeSvsrnP+7NDWgTRDus4enKWV+8QvKEZwOhX2jcKvXvKoGc6YzCMk
oJxdQwMHMICBXdL6rQRn4x6hMqR7crAp5X2gkEI8hW3T0WXk4Sl8dTmGDBzAXXJT
WPf9u+iD6/0vbu0LF0mTOkCwU7CsBlUklazGOEYIULhlinbVDxZ+Bx/gF13SPalS
zpoJHyoETXNtbpTe6tdrk4QQvLv0puTWzyDi8KYlc33Vba8jQFU7vjEhcCAjNOJ9
lo0a/DCAgGNdaaOMfQ//Dn5eCnWBZbSEnU92Mb1G1fu9XmyoZg2m1DuZK/HU+K8e
RBvi7I16tGnmnozeLZR73sqhRnwMQpEuxmYJTOgeo42vDeqCQlJvNI8mb4JkiSBJ
88WOiiaVGfghppvmhyWqwvV5efbUNiaVzIavOYPVZZwNW/0Q5zzaHja6qGd1/+tC
ieUmMzKQsSr1fuS7iK32qLWZe7udkwrPUAx8hq1HIJueqkEEczuq12Gz5pJCG3+M
K+2MvWsBKQzte2+/aJZuFr6/4jq3XSbmyjm32V/ts5cmTnQzNQdcSlLmdoGENK5c
u9y3DRsL0Uw/w0aVKI/ECeB3zm2le5mBZ5NSia/J6NYWNqHJSrZVfCBdh/6tqdwm
5MGlyA0cClamrxUvmGTy+eGzHuqY5wfW/QJcqlC3tj5mxDfd7Z34Jlho+1eJJbv2
sDEt6wAneGA2EJ5DwMhGGkpH1rS4Tg3toJfiPAt+gPi7aDa5ggfYh0y77G/vr+IP
/vapUgX0+DJfrgRfegb8DW156JvldP8ptfL1baBGh2BNIv6B+Vai0hQq0msV4LN2
R3n3ScjKoqhp+6hiUUDBpCfGHYQKrIdsAEtdv0XjDao9GIOitBjpQUaK9pbzrg3d
1XP62DtCd2Zr3f7lBOGA23WkePLwbfQ9WmwpvjHmjVov074+AcNtOaj2uOxX05ek
pDqIfQZ8snPihTr1puAdT8NJd19X4aT9Weq0f44Ilis63t9XITjrTzPMhZDuaExY
h11PpzaYZjsjBomsvF90hng7hNGJwu87zEY5aRa7Tb/zD6tSGWuLJHMGGHjn3rdu
pCcCT4T38NyoYNgNOXu6gk+gm1vvuLcGk7f3pjkXEaPyUGGINEMRgPzHAzgVeaiN
+77BFlwTk4PnUBFXf6M8kQZfD3ay4aasa7IlyHvkF2NcvTHtWF0ywO0JowFWTOQ+
Qf2V/n/tZoHZpbiAeSZqlYjIZH5gmJn7SuJYTblsb3NHeWYQ8vPTF4wq1caqH7zk
220Ab9QqWhpev4LMcFFxhkJfPJQttDdRJ78geCfz1Lded6+g7TzwkKeIKEr5z0WS
Y7TPo7f2SjPvPS1c91QLLD/p2hLzTvcAdagg1oOnBhRr8cZ5W4BWMcwLZcrI0Udo
3EsMZQ5SAvprFJgARnaU2FqGH+K+B4qV8fr+os7ybadpNETO1MH+kMIz8Usbe91X
lfP0QMTP+C+Alm5h1DgpZr9i4++jO7kJMdqaamQ1R+rMbAGxhHnCEBUANmNHvp0d
MYGfVnmNJVfsyhaKE4YKCO4RiSui7qaKnTV3U70MTUZG74rOqARcfb16o0Y3bKNW
9jDERa/MA9yEADShjIY7vxm8xxkskDJOamgk5higk+D2EbxqPvVQ8e8a3YJ6m79T
vjVaP8AiJgoXjU53o7C/lShs8N/H1KWWMPWRe9ivX4Xpw86EUUxV4W4ku5zfEmEb
HCl3HYw+R82GT4Bbu+/E195TdT5uV3EpHJbInU9Udv+4fq3pC2OpzBhJXvjONIdu
FYvHaS77KZ1z0HNP536Ko0ifMaq9fA82WI+FcAdEIUKCb8cNEABOYkvvUzss/3uj
D7i2wSF/nnn0CdvgYmyx1XpyEghcKS+clEjcz677vgNOD3AOSfbq2wTqpNo2AX45
j7dWBS3fx9lKFEFGsQrA1k/m6hQggYuYvxwfAv+jhQCVfneBNjVv6Bg6GBZZyzPC
YUOC8blhT1OichMP52PXUrrIxnH1RRvw56Ceo6F8pQbj3MfnY3JFh70mgZviqJJM
uubbMSIYg84nwZ0u2q3CBRfUfypFeRxJtGnU5xGB3lsZzfLcQ9BFM42i0jogKFYW
lwjqgG33XhzVxnmxYm33//p4Qg4dSUipjXompPYs3P5ZZ7lXs+jb9AfeeeCLPjSJ
zF1YRK5w2MmCHMGbnPtpegQpxFLg152IxawPmE0gPQ373ai9tA8kToFl2vWoknRf
y/yWtfYwZZAutE8Bkth0nAiJUh6tTdc2nD3nkDL+f1C2wp/aTKC9Nhl1foBRktSm
7JtP4XCCy5QI+UfN2kKsPt8NgjEnSmXa70axAcow1f40pNfPHoVxgeFkjX9Lk/JW
Dh2pVXS6r3BkbJHOeK537Y/CKI2T7soE7t98TBQnoAKuI7QzHjgPa54eFeR6V3SS
KcLOgEM4iQAKSeoiyNKs2kLy3n6YwhHiZDqA63EV5rARy4n87o8Ml01Ozdvuy+kN
4FG9HIxrJ2AKz4F3/GyQ3gsLnEM/+9+SlyfgtlnyKS/K6Pz8O5UYslApn4FY0BFH
HzumC/ZA4X/upQZHGvDD5OIVOtZEta/B9vg8O9hDPyXcrw64cdmGUWrSFzWhtAKw
k/Y3yaTDkHZOL4/qk9jU5QkC8bPY9xBqL0ENIQ8XZhq5AZabjUkEuDJd6SMjhf/D
Cb3DpyIp4dn2YcCEzAUhvHI4r00AUqW6XJwKbMD8rfVNuaL3Q6+U2+PAP46/hXWk
2uvfphBRqCQjgCPjvF+0fggw5FZO4evMxqxX9z2bYCIgqKwDBocI7Gfp4gRNrIhs
i6GtyUowFY3vvjLOvPzY1zeWJ6tQpbzs4rkPZZzfEkbM3RkydYmjcX4jL+i7r+uR
NecPzDcnGz4FwjlYFf9iztbbBHQmrFQdsgPAdlIa89GfFLtlfgae+fB/WX9Eox0E
2ptH2LkQJoWGokrmJzNFVsIeQ3/NP4f/e8hMkYMp3tjQvpe2LvhIMvQAonnOlNbI
skxt6TPuXFNQUlC7gfeE5zxHdV4XmF+X2J08nXij7oO6rq8yI3f7YTyeeG8R3Vvx
JeBh+vSNMbfykK+OY2zTdigUoEQ2KV137UoAID6OsvKd4H2/SUq+2E9ALA6sC56d
Yk5MEPIwjgRO5cxjBSc3PJG0NIXEmaYTfvvP4Q1vDz557eC2Yb1C57FEggAxnfxU
eweyZtSuHXaPkWb8Dkv6GR1CQS9Dp5AX8yBy/srdaKos1hdDdHkALkvLPOkMHr3L
G7d3yUqwHhC4jjcEzAXXjKxWpfCzanbPlBOEIh+1OTXbKMeOvFgvhCA4mc6yF3Kl
lxy3aan4giGoXOLUeiy4bf9XSxvPukcXIvplKoWuBVXf5k8Ptu7KfdCYxf2vW0Yo
I2MAMFy98HVi2lAHcKkI3S8zEIA4MdXzoPxeNELHCNI6HpZGVQfDHkck7Py+Jh9s
dYv6Kw6AyJJbw3AtFrxsKXvWvVvNN646c8t7mSPR2+KqDbJRgG04AzySXYXtLVhT
U2axRkZ9+OroT07p4e0z7dJZGqO3kzvb6MS7OrmIr0+LCqeym3IjQ6spNIK/jO3j
Lagb08ms+UNtDAawOSIBY2aV/mantcIw387JLK1bb2TUY3Bq7KYnCOq+mBdP2sze
DNqa0nQHkRPw5QOo10TJvr1s3CrwLowYUVbp7Y6sYQteIMt1k2885Jz0KZdtiCNK
H05I1mHauBYMrzfSUPAU+G27fBDRDuPr+6OKDlh+AgF5NuTIos436Qy4Ga1c7ZoM
yccNIwOTRsdLPDroRC+rm+Z+TvnBobTj7SM4V6/h+RubZSqrPWx1rpgh6DTrGPrx
AoVXC1/PQK4fTmZwOWg+4ZwFsopwEeMy9wcNd7K+rrBkt5/i4V0Im6xFu1re9HqJ
S8XaezkvaOnBd2tS1sc/+90GB5V6FBobPo/Mk3HpI+9fpQaNzDafDWevfLZb1d+1
4kB6Jj+XbNEfaBm03UtImoFrbh4hBnzVHd/HQsrdHeSfvAID9VPBBkxFr7T/MqrY
X7fAtwUZCjNApvC3rOC6VUoABkmVgrqGHc5Wk1dz7ilGSp1Qz2hnrCT+u+WJAv7b
7uZK827aLsiNjrvR+XynscjcjSdDE3h9FjZZ8UqVo4tdDld5hZbTRG8+1b85egM5
59OfCoIyJn6Z3KgwNRmCNgaRsHBl0lL+pWO88a//ch48vSkk3oPhIHzeD20kJnYl
SWh0mpWLDCnx21qbZ8GmgVjCKTPUrtSOELYo+n+oRaUJKlg298OrJMaHReQa39cN
LZec3urYQ6Bli7Q9Zp96Sg+ChdDez525fe70An/1zSJ7WWe0cfMdWGCkNS9UIhTg
t8tR9TR3Ed8lVr3v9dTAIN6mcLg64RLtJZPkxxKcrf7V3aqKUEfWIeHruZ//C8nK
1EPf+k+CcAwEWP11FuzAseXoG5gZmXwv1pGUntnbV9dzTc1NCCLyJ6zlsOeFnHx7
YurqreybAXMQAQvmdgBL9/nMGvH0rAHyp93KVFUiYLyM8tJ+qy24UB1dR7dXXOam
w8bmcTWl/iihq3xMkkmXjh4l6u5Y6ZM9rWaK28oK4cqTBRAjJXPSAL2nAVxDRwCd
UHgYJm1uCyt8KgL57VPFf0234qvdNy/OPNeDJJHlpylwJ+ZpJBosUCMJKOeF3gRW
rOxohZZ9z4azvT3827FDIOZe3Q3pCLUORGzqKBRJvWfDW3qcVDvDG2dp9cCMIO7S
Sd2/e13xTWXLpsJ/1d1gt5Gd6i2iT82EjXxUE3Eq70lvhfrKwN1m0wSIvMbPhMMR
LYDd3ZhEUHYSMXPkHeDgbYzIqArM6hRyEyfcS+NELcjwZi5bGwDWbhUt2MTDSimG
6r7wXl1c6j1ewgnfhKtxm7iDEpXPBdGZQ8lbBWb30TGDK6mP3cWCVFlVZ5INdrtK
1gWspu6FdpDuHHLX6wGUxgHbIyb2Pis+pjSd6H2/J7MCo2O+NF6gedJNXIHqB7FA
y8zMT2d0KSpC/ifwkswLyJBiLBdn5ICmduDkVoJIk4kwcigJREROh8YuGl9Rp9tu
CaTxVDzZ+gAR90Y8amO3gZTsqsqs/7frj6bLGUs9KxegtWZ5r8BZKVmpgM7WE4g6
bPvaxoOXiuW2y4/TKqoo/I1+Qse53R9XjbQHmQuME5rEJQxgVynxuJ1hpSveLQA+
cUTOBmVrptXply7cs0MYEKE632yiia4zHfp0NSU5XALxdHswOlRHanXIPv3rzG3u
xeNtjtgeewo91F3pG7UcjHPYpET9ej7ICXHwwHV/T4bmyuuVAJ71HnMXNcfMo0g6
jcp0m9HKeoOqUQkmrz/iBu8Z1MlRC8xY5jOVfWQ8Lu+at16j2h85Xl3kZxBaXsJh
7GLEOWUGdiH9zwZGZCRD4tp9sBsUodocRbWVPEzZzeLJOF5QJJ1KAVsnzjbGiM+4
6fpB+NqDm2rYSQm0BYiBGWu+VoxIMgCgRrhpq4gtaQV5GeBMLds1mJmQuc462Coz
DBROUqzzZVExY2C08EQnzQN5uNCQ1/dVyuhp7Yw0v3SW/Fz8pmjWjBYTF3VLzox9
hyAKFFCdEfdVEJ4AojN3clNxAcGbWigZyOEBWI80MMjxz9B9zx1d6FtEI9NRdTX2
TnqZL/FA/M2zRTl1h7CjDr8TsHvCGMrM5n0+N0rYJ/9SI+J4JYFHjFGq8EUzYl3t
+L+wLQm5+FnR9/sTuTFG1XPwfCMufSY0qp0VqXnpq4h/yaMTzPQQMX8ALbLSZKWD
r4+5Qd1Nafzvdg/nrMuYRttTgVNCG7+YcogKyLB+xai81F1bvHj8Osb/z8VkdlyG
fILI5br72PY+oclbRvad0qQEuGV8UqCZceERpj7WnKiaJ4mJN1yvBg/WC211WNih
Me89CLN+bz2d5VxVASXgJ/u3V+txrgL30+zyIiZdbP+i0ifwYCDzgm19Y3g6kcKC
sfCmTRz8DTztgCf3kCzL1QcIGWfMB5OA74aDF9qd9xxvc4vcq5bpDgBR5zWXuKiD
yc+ijrBF1sifKoLun4WNdS94Ufv0ce0DjVJKTLipjRYEOh5OhQENodfHUcJdfuag
VY2bNqGw5DPiLbdwasbqxNh7d0xdFtNkpkpl0GPp5W38rzu45RjXy8HxVp1Gf6sH
vAYpwrEWbw6hDId6PmzIO0sFPNrOYwyc4iItVZvFSgMeRkC5k6aMF+dgDK8YcHja
gbJnN0kM3VExGTwl3v3nlPEGuIY5brs0R+4RN4tY9LH73GY2k2yjGlBdvUJUWkaC
j3DyLWi+aY21QkmX01xc3oUab6dhl4+DepivolemgrTV1Cs9qTijspDeIjNnAfLy
ccCu+rfXo9qe9pnHlwppTJVCTp2uOHJmgcErvlyjW8PrGegbN3xWZ1j29GqLMBM9
ypXYmFHNTZKx8Sm35MBPw6gJGaX+zCYAl+Q1KeMcccWqNGhBJtIaFRvQnDznBdBq
m6wD+EENbvAKKlj0qrW5ldw0t/qBnblFll0SDLrnTQWMYvXqUgnpst03IyEk6VGy
Y2Q3N4RQVmGpMLA5p3bFQiAwMbgztNfrUJ/ZCS4WSPFVdw/BoYqevgiyxQKbB3DU
tGr1qrZrgjMC2sNmAPrZ4iyqx3JENs9Mwf1+0arUiX4sMN+AUNot/CBiFZSTUCEi
bYRSFwoGUhucdF5w2LclmHzIxkrdR+HXli6QzeajOMnf6psEcd2EMRThgF0h4oXp
nVWrb6wkOLbp6nvlZ3WhmT/s3ptxtLMR5Vh3HrpNSI0yqrHbwDvqdlwhmdhUS5d/
QAi54wAkavLFwIiNCHuCzHOuS+7alvDD2Jxa15KMDkgnZoypR5SNpNeQYWsAuufI
+f+V+PD4GCS+eiqVcIFW4POpLNQ+bGpjClzgzJDoH/b49yk5k87M2QmCB0nAXfmB
r72Ohq4rAduNoprflFnxJQFd07gkJnjbWsHFc2uuZmzV6quIezoKgrYarJTlss21
CzoJErTNBAMqCA3AHQnEdIhZ0zaxzBTHHNkaxMYUImP+BdbWA/GdDOyv1wR+ZBPf
6NBSQKOFY9dIfFOMgri4yRwb9Rds+3CFqTOdo0cGBd4s9ezCdaseuOP6eC1UqOJK
17HzFisysR336hlWcBVw8Rk/Ik0GEHoFtB1p3c6nZU05lUGqVCvesvsZq+WFPzxT
v3/AY3Ob5OdMQ1KuIQ14Zhq715odDsXKaXsKQYZbY75XEwZkNvrpYz0D2z75b4vz
z2Idvskey6Jlm/QeW1YY/U19ku65JRH1V3bDzpJCFzJlrBzCtAhRQZPwE7C8vfoa
HbrtpeDBhxHZ3IQR3uk8QNdbzawcxSEsOKHuf98lqEFEMmgKmosnIfnBV0Gd3AOR
FXRr+OxwoAJ5PpByx9cS7HgkwkGlpf/sxHt9DqhEXupDzuvrtnQcY9vSoM1790L3
gFMI7m5hx7DIu0Vw0cfv71ZUnCZtqggVBfREqNJFVJCBiPhU6nfplB71p+Qa3uiu
facVM+75zSi8Nkmcv0HS6Ib2ggvV7SXYLtLqZklPQcoWYkn64lNlxmkr1wmamSMG
XQKGsWfmlIusrt7M/pKlOxeUU1PbxSVXcAGE3miZD2fEtnWrDQf6Aq9knpy0ikbw
/cEavLCvmkZp2NO/AWG+2ftO2I4lmydiGb8gCQvo/lDYwaCWVr22SN/encwd7vUc
0ik+IYEplbsMekonOy4UNz2WeZMajRrkOCT0Elz3HO+3EaLDEjMVz91CFjH7bjBS
Iz5iTV/5W1qkCI92hCZoIn4rG6ngPOn6tNCCWLDd19p3j5EPR6F9h29/QZvrZxQt
4MupGGmKqm8IA/bDSW95jZEC6b7sR2vsQD455milHKrBGdhGqZAj9CrlhSPEeWYJ
M/Gj3XPXZMnH84sQKXg6yNjtYfn4wIZqiFtawh+L+M9OLLqPeKXbI9Qs3a07ym0x
BimXxEmJrnztfgn6fEPfyDdvr2hVBHkaS4UU7x9SOVrMEZSXOjw21EFZHF90Mljw
qahn7x0Pijfugb0i/5+xvn8/BkCrOKpCq78a0vMrp40lxzkprH4G4he7KvKS0YKq
j0hO5iK2/7+t4/BijDs3345sACjiyYe681CP7lvsfTyJD/+iazRWJQT7vwRIEOJl
ey69iHpQW0nJYQqlhPEDSR3Z8VBITOngSfXn0vZENOtjNl1ecOfZ56G7W8KfGWfq
U1m27bJA1u36ZJwPazTzROdzBtmCXsaMLgJ8QHpMRAUX6SMi99ccHxRl1GmtMSZJ
bbB0aFHk1SO1aWbHPO6DNVmrpSe7yfQm6wc1nQWAYYdTt8Omtt/3Orl8uHQocCDm
p86/ugYzkjCnwKptO8idaluQ5QE6hyeIAgqAXvPiajCBwcQo/cSp/eL1QfCvsnQM
WQ+490p7IUgZlUd2Jw+2baDheFfEXiHuc+14zJUi9QnPi9iQHLcgru3J3Apupigv
MeE4Nx86lR/hzSBi+HJTDocRSbeKsCPzbgz2McWWnzOlXRemmYdpKXanL7SyjsBc
i3Kj27V/L3we+pK9HiI0v9okpQtoR7BkosYSCEkTlbSyTBIN7GH/A8Ss+T8VY/xz
cFYq5nHzIcRmXbCZWMkSNXJGjja8OWcfOLxT1kcQto1VCgIs2wuQb1BTWlNsQo2R
RKTkHByfXcq21irWp4kVZ+3L7fcBkUDoQjvVMGvbAu8yS9HfbpIFIhTSQ32Jeg8N
4YUjzcFMeBuS3qB1rZTYirznTCLBltFLaNWEdC00JWiaGGI0vLEzULQexbRILQH7
gBP0Sj4qrOIYhmJBXSSVrz8UD0EWlZPG7LXbcOejdlEsibnKsGZselSzDcdU+AT1
5luwYUMsYunXGXZw7xpjAcIi4E7o3IWFKRvvDT3/Mzfom/zITHjTqvxrZSWZdZ2+
tBLyqT/VpIl4zmdLZLO/pc9o+8Dk6oTpLcgLWKCfx2KOH75IEb28C3c3iuXkQ2jf
zKh4+sxmO9/sL2q2n+eBFsmIbDlq6piBvx3ELK2j76pQXw1Y+9yk47M/e8mYxFTF
rPtXl8P2USnRv7VAGXtHkgIR0ZPNWIYFELP0rt260K7SIbT/lwvixM2l0sH7xMB0
1+772OnBib9YmF+GO+VCY+K2Ih4dFXGyxJJ9BrS/DjV+RxEsye65FsCd2VgAtKZQ
W+mthBIYQNhcUmouHD1CAeG1phdWv6RafFki3oXyIbDW7oylHxnkMq9pbyfZ/rmU
65GspaR4dPXum6U21yG3HViPGFzJIHBW5SYyBrHxKx+hCire3wOmSv8D8LidlGUu
ObU28ytJhBu5ceTUm1jfred2OLzeZQy0AmVFuNvztROSNRu6L1j3drEhz6azaWxU
D4lI2VNh+WSmXgY7SW+HViPxS1FOPpdWnGSVYjPwXkonesI03rYwZBYM4Guw2tV7
2OuqBcqoW4+uaarV9yc0xdhNxUfSJRRdwoeUbS4Pkhx5abOhgxKdLS/xaTeqeacB
NjsEHBzjrRVwR1xA+xsOXJhNnFQ2S6xJEfcYPyEte3RMtBCiIMvYcleXT31IT3Mi
IHXnzFQdX9tXhWIRTKgXTPKS0yI6a/BBd1qwICr9wHAg/Z4ep/Tmi7oq1EJaA4Vw
3mHvG+JCnWxaw0vpvzrbQUudZQm+fN8PBY8pTpDvp5M83PEk8DI4I6mlCkgohEQY
jAfvPxzoohxLYLWmQONz5zB9Q1cqSishzJGC5nECRogNNucgNRbvVzWVgUfFhgbK
cEQ6KF7FhmbZT07RB1sA2xuW2A2GaU9T1imx25k2M0fWyWVm0U4qr9xD8nS3+gX1
oirzjZQEFPp9BCsqYQvXRO/8YzkmEd/sg5A5N71puCobbWMlTluxFXmjs2PrYArp
bAe0bH0JbiZZosOjESoDjMCClKyh4w+CQqrqWD66W0gUCbZMXwwKpTGcoggvxmJr
nzoRE7n4yyURnnEWR0bgc1oCal4U7MJvFGLqqz1dDkd/wS/x92Bvf+hjwyJEYk+W
nVutgj/FwFpxZcqepCDS2ABSp2arCQtkrKTlNTD0O/eqiMacp5IU0kTb/JWJSUKr
EgSySKr4NF6ktmMpK2uzIfskw90+hAk5QxMgS2R4Kv9rRZg3PPj6bHhiEcwGtQAH
cx0fAB9MD6WGcvJ/470zi+3Veh+GLrXySGcg40u1b7PxHVMT7XKrJhmtXDAsgZ6y
BPG4+v5b2YlaXbIfXWK/NHOJMx19/4R1drhSUoQIS3IvgAoFDVEhPV0TYRuGooOs
rkqiiw2m/Imyo8hJzosTpc//bUsmXcFKySahAkO9sflJRhsqPiZCQUmr2udNqja6
GyfDZQdhAhm2C1MM/PkU69J2N9SGyhErLPTCNIfFnPZGe8Tn3I0N7VO6H+pWjlmL
WVCde5lINbI8Ubte+EEzt/n8AHpgn9JuUCh0lWiOH4bQtbQ1Re/QNaymwXn1i1eb
DG0CueqdftV/mkHTX1mG4FpXaDjWodJTrcDQkXMnz89uzeALOqlCFZNJ1TbH3OAs
7HlBdBmiPW8Gf6a3u4a1sXrY5HSkKlTMZPOtsk4qZ0ng5ot2zGLAQYRjX6GYXIzq
qbdEr8uiFDI0GzYnDNv9+i8cN4a8itJmrT0fYHtvDfFWVefBBQpHGYetYei14sxK
vXvTmG35NhGTOwZGwn39RmfB1aV0AcOe6f39oixJW+T50poM11axZydMOzx/NDys
ay7GVmYKiqxrD6Ek8PW74nO8TewZFTVz8174OXEX4ZMdXF4eOzZUZ/jEzzBxKYue
+OxIm2wTeRAcGt3i/rJDwUeZBBhV31/DD0vPVN31MYbdTIRnQIbGxo9lTA4y8UtG
m1bWN5cHdovo6XwtzampBPCoFZGxa3ZHYIEuW9SoMRMS8j+uMw6/Blme6wz7V0FZ
FoNEUCHS1mRRYbCt08cxlKN7lJ03QkObBmQyZnmjMNfPITPxeEuNINT7cHL2a+Cr
vpgMaadXJMApKIEHJ0WFuHD0KkNfv6FLKJhfw97o1JsM0RREwzEY8mxEZDQqla97
VzJEjKIb+8P1qVzVQU7Gfqd9xEENl42YXFr2dQkUVX3ah3S+BvMk+05cz/eEAJ70
IsZULJDa8YZ+rjpacYbNQgqyqZPZ6X8c9gZG4wr3jZDQ9awev47gL9o8EHzNkaoL
QXQmEBfJ/8++VdFlissOOAk/pncrxYghABfzKTLuoJRxT1iA4d+tRE6IXo2Zt726
Ehml8kqGy488Noq/FAI1pQwLtVis1IdpHOV4aWFiMNeteur+hJ3QEzyZGQGkZ3Z0
AeW3wse0nWsm4HnX/V+2ukuLHa9LN4SWkbM6WFVkUFvmu//XI9yYqt+BhEtSJDof
HVpcuqFtCDP3lEh6xGLshHFu53S88Idn/4ro0kA9Nh0mtXmNxfe59p9lWB3C3+cy
rudbT+9MdM3RbDLAhOhdmtn/w0hb7D45vXBpbZU7ubdueNkvoLWgdcEc4H7IlJ55
jucKRs+qqGb8wmq5b2WFOGtmWeIwx07GGBdaorpsRPPxoV3+gg3zrn8wS9xV+c5B
/mJZkK/b3atscPsgU7MkHblw/wKkG3VoFWMvsOjsOV76xKoym+6evjjnYwTDnHwM
3RmxmXoikkAsLBOzsMzPsgPkrVlJJjhh2X+KOv+4HFwKu4QFRKUJySuXfZytVvyr
WTSjGI3KpuhcQYyzUlhbgsJMLOFx+Al8mRMrtaansoBjo3LP9dQCyfeHBvAWDwMn
1jrD8pOT/Jlq+gW2PUI6slM5lMUOHQ5cMfTEeHnDc4/L8KN4UyU1ToFdj26JIafl
5CmAi523EHAOJw2+Em2v249vwrP7cZjPSMCd1xtOa+8cz+NuOQJOLnH4FQ47oc7J
A3RUsUCRVny/o7LbZ0PanWyVm2QPSEkRxfEyg1oPm0rfsmj0musH2WEn8R5hGfnc
DhUPbiO2ZeAt5cbOZ8YsFTMJN0MZiBfodu6W6X5PxXVGERX1MYlX0slHS1taMMjS
MMlFEsX263arWnavI+qNH1WZorapCaAg5Zd4eVHRjfIEgrWONbfHFzyj1CZDpFMi
ALJZKXHc6/1jeYWNQhY4e0mfy5bYKNGtuc7T5UWpj4/T8VJ4DRkSYgqvQ4XRfVDz
jovKZJY/tRyvi+set5YrIWVwsZLGCF+oRJtsCFFtOK4uRFRoWsgag4HyOteEa3cf
eaRYSJpdp/+EdQIOkMiT/gDLZ/SE4G2D56HUeni8sG2SqKnk+3t6/8ZDX3mTnXlc
VZrUDzFAz2bqAUmPKwlgXQm9Zg22xUcelLkXdlOBoWPPR9y0fGOiq53wAZxVjox9
jktYl9XY9ow8TBHGWEzlKrHDMC/2ey/NX91msxDCnzP2MT6nhWLiky31rMYmPKU3
a1J4Xmpp6FIqYDzfVjQ2ZfOexLQV0v4lYzQZEob/UgUl+zloy5xtr8WG+f9Vi24D
jKQUMwJAHmi8F15vFeQzGWKmMahtiwL3HutR2smzocZudtLIla97dhmP8Ic3HMNe
0Z/uToyejomWN81b4Vn12Bf7BJzxVX/CRcL0AqWv3bnoXdbaPZBu+jYIBrS4zrJH
8EafV/N0W2DnnnkBdTYWb46UWvsNZbbBNYK9JmFwxwPf/YrsBuy1fyKSwyVuBxfH
ff7qdx77XrT51Fo+FET0c/YjAfNb6Guyx2tF2vqG9G8uze+cmvKm9a3Ns8GmdWTw
WjKQg9HkdpFeBWVnBQu80QMV799aVSVaDTV/ddToYCKwHeHQl8WYnUc1ZNFTzOaR
mJ+9N1C7kM3/FwRx6uq7cN1z0X9fWyUK2ZuPTXCr2ZSkoUJl/t56pnRfiac3n/ph
amdqYCLGbbxaD8z0m2TzbHqv4wydJcH//arqpJ/Lh+gNRjt8mDzyWQP0pytvZhYm
TANKRDnnKriYlcY576Of9YToZsG9HB4u08I9sBRIUa9BvP4Y1y0r6AL8hIkeJAd7
g6oh05iscMzgzgkKdfEvF6k4dXJScKt+APj9HI3DiyN9fTEnmzp3VQBJUBJPtJuB
HNoAZxG5pskjuPDKOwWF3wVQ4ckBjjWhP+/ZlPmHryKGO8hpSfUvyqtpQJ2z8L1/
nkXytYbGWS3vVvKm8RqVMuqjB0Jk3rvJbw4ymMmF4uaTds9AmuEqAtvx/ipdXZ2p
7yMhcSQrVhOIg7RYYvYNImyveizllYCVAiReYEdolWE3fYFnV58lyVCFwmt8ksXF
bSUBEkvXxToD9u+5lDNK2xpjqU6taEnocxUkjEhFBehINWFIuCHikglmMDOUfAHs
hh747605ywP5/RkLMMbo3FvLHuO2Pm84DA4g6PgiF/FBnGj27nireiZH8ar/QkrD
gaKIvOgNQzvwAOqiYzRr82yt+KoVnnhSfo8Wuc4hK8lBIvgTAFZOfEBxIFt41/m/
xVzRCAaO9nxX4jZ8412fSBDe/unfMy8b7qdOdeRdP/+9G1XW1H3e2dksZ5nPzonM
7zVP2eb9l+bvzi/4P1mupGDH+YmR1piS9VqsSQ30D1Ct+rlI43LXb5qi1M4nBoWY
NIXIrnbZIfxp/swICK9C0s/bBRcN1705uUtMHnJloXSP7UgQdQocBmT4pH5fAgey
2ZGL1h/d1dfw0mnaOwE5xO5U8H7sXVelkTgGbKvRlHybjGh9jlDpSBD8d5bv/VDT
1XH2MCtAKKtujHETrMzoXsS6vERTdxRpLGDcbphjFWuY8aD704poVVn1v7YHA9IG
Cdihl9iZUMGvyZ5SCB9qGD9tvsbSiAB4gNarNiuPzb6QGA8JpROz/czfbTuzScEj
iRtvDBjJRgi+MB5hSl6M3rNzoSIiNFo1R8VGsu+PMfLQUysheefEy+laTaoxeUuY
FKU94SQcFER6y6XmbFVeyz5uUI0628YtsxvrqiOYTJdO48VJux6wnInmT7ZZwKOg
T7eh3TYWbbvKbiK/MI/Wl0IvhO+j8xS/fTgTvXnLf5SkK8flT5VGQI+naHzxOJQp
kboBaCLRwb2GAah3dA2TZ3m7m9MqVD6F+kZ7V9dgkCdqSAenq2SdWWjm53jkI6dr
e8roc4fOg3Qkq1439YICcY06VEFJsf7t+phszahYfAh5NSyR2g+AABvZcofu9+8a
EZQTn0YbDnSGFnOban/TOHWBHyKJYfGOHCCnnlCFeqhpjAesD41ckrmpTjen3bIw
MzGvGtWVprcjs2viMgKNJXrwsMlOyQXFFNUG73RjJXV5QtgcCfufKjmdlVPu627m
1/kq+LeELDYqxRF6sGjoFXCX7QyvDRGHMUQZqjZmpvl/wbkHSrwTgEEXLzjerKeB
FkaFhZ0zkEKT1s6xcrInwPGxKy6MhJ9K+xcwfrtt+40O98AkysVKHQ6dJXq7/KOz
RrqnkJOcG821h+LfwQhsmVz8rPjeCASgurlTkKzihjjtdm+3PIzDC8q71xlrVFTJ
mr+VHfSFG4d1N/VF+QW21ECp0bK8DAnH/Mn/s+PSYxE5jZ8s7molt6D1Bf6pQPr6
FzuCDWvoR/PrKnWjZX6zeS2pxChI6DgG4ooaqc0HN1MCi7wFIJDCySj6+3MZ6ljF
8DxpAfNKu7ZbM1ygPwzX437wzi5tICJKmbtcddu/q6xlzYZ+BCGfG9U0f07M0suj
XuZXsgQFcIZrnFdHG5yS4wdZk123PR6RqeWjnOs8qTZCTsvSGwAawwmeauPTDr1g
Av88llzHHYsCfAom5lBSIXgwBMMs+rmk/eYNFwJNGwxppj9OfL1P3wjiQInodtd2
LHkYHJI3JghCXJPoKRLmXkx+1P6aWITr29bwXpC2eUMO/0WJ3YEiPUJZrCD+qk11
Pbtk2SE2UQuNicN1tN07e+Y5CB6loelRg7BevnPxzTt2Nn0jhNzm6iYIUx1o37La
ck8/+z2T/r0NP2Odn3bjOR9nV31T5srrywTkYVTVKsfU45tnFCBeQLM4jqYLpVKR
1e2j7o0wGD7s5Y7j2iZQ2qqNIvnWo5DKAiqPLORXKLuuCeEU0gsaNWxdJeaur7BR
bSRQoLA+g6eJRSj2b4vEqZLr8BCBVTmmpJmpapZCex7ewluWZX5Mfh1AEHzammbk
wN9Dm5ffHfBfptNQZiCnAnXJYsNm3QwWzRleulGASUeoKFqBbYd9zsQyT5Yzc38b
0Vc1yqyHgp/dsE0AyKWYbusbaY02JRXIGPX21suwsJfjT8qLb1Pe7TxK1TCmnRIu
dxqYzNJbzMnui4l5HwWDZ9JO+7comiAoJ8xtVkCCEW66N+3Ary6hYDuujHM4ISzw
tEB5xLcf0y/7SEobROOgqHp7zj7bx+V0sspEQjX17/emu11Ai79daw9oecXQ2MWL
IDbKPhLrupHkgxidQWEpmNv9m99/mECRzgtwr27Ug1EF4fEGQ9QVoZlayThRl2F2
kGUdzQtvWRvUehnurNuqeYPkzHiMBVODSE5P2EXNT8Gf7PZqHsgklb4ye1FVVHQ/
h+WjTFQz7ROrDs6e5naFq1kuwAae+MRsik0EMY48sl29FYSfbEN0SrIkIaMtfpip
retsdkxSZAXXB00lSIWrLdLNMZpBnxDaE+VFf6bRFD8AYn8Rbp1/G2zeRSd7AYSa
DCCYhFCngzOSCr9pIYo6V3OMlOaKLvE4j1gSpA6wbOzL1fuEhXb1hympAEzDx3/0
t8971YWPZzBVVH6hjdvAYv0ZxV2f/m5HEJ355F8zK7ijkvlCTFSw2vbqVkxcP8oY
urB1q5d54LDgoInLzTSjUFJgg8ipzc7T/R3EkZIhZqJIKlRrVL0BVIYA8+DqHK3W
czdgU7btDs9qQqN5XRGB95kTjRs9UQEKcNPQ50pvblpBUfb4tOWVMhiqjtfV5hxD
Zoiobe7WklOhwHf/lFj2h8FJ3EbPiazDctHkSxtmgxmkVtQGOTiKPfGSi65WH4Jb
tmS2FTq19JIJC+Acs7ZACV/78KXbGdNJ46h17zIOjSVn156LDwKrta1yMQGzeWge
TZ87Nky83wkswA8pvZ0IlCMnw24mROiFAH+U5a7Lm9A1w4ODmBGzoQduU/fniR11
VLlxFxZw+hRUrt1RIMS/ah8RhPif/G2uJgaXYuXck/PpkeeVbYYhu8COqJNBCMT/
4DEWdRdYRKd8YiVOGQwVEXdfdz2X+0rUA7gH1QfmSJDUR0cML6alkshQnpICt1xL
P8Lz80fOQIqA1fsptUOLxJMtjQrl48DaaQYm7NX1fL5e+uvZnsf40aH926TrK30h
mwYDd5Qrc51qerUL70ZPyM7bvo7ZfbGPcnuHFaxcPgR6t3u9D1fh4TKAALs1Mwtm
wYDyCZlnu3TPVeZu0hfZVPiF1BdX98f69Gg4nWszPOXWhRl6XNUH6mPIOith9GTj
wlrYkdTDMzOoYscjp/tniPIGfhIT0aF84BXFvGsyEumZlwHGdF8nSYJIJJdjGp48
hHLnxhsLFCHRcf2quP26BN/wtwQiMZlR32yetDoOtV5UnrWA0y7ywwVqw2OeblnK
q4EYs9NvX8Wnh26TjZIJUlGrBeFAZ/sckLrrp9I2P6gpT8OVzL0EcSRQhPiEyIoS
l4S1aQVOWxK5wA9rhhyIX7c7J43rAMqOxWMGyt/3ibqzvaztdDmzTScTRq/OChT+
62cNl5vAoG1XDa5/n1SO+sM8h/ZE188+7K6Hs6qGNaHU0v7FLvKt/iocf5ikqXLF
MvvXBKNe2YTfG/kTYd/Xkgj3NmISTTqETDA6ilW45f/kh0gTspSVruo86/uMA60v
rd7c0RvZmdOywPKLZuYcmJA4sN45oyZdde+EHBflIV+KTymvO0biwPmFXhJQxb91
OoLbvW1hK1lOpR3I9pfb7bIerhj5wBjIa9y0TFFF3nOYi/kI4SUREJ/7NSiygkuy
VLF4KQ13lQEIzoi92JZm940Dp9l/IyfYmlz2CFJD6iM1jHeOr8PvGWnydzCP9zFK
rSmK610TD8nJtIjH0sVCw+LQWNiiJGkQc5FjMouDpce1gJnAjXxRXICTi3gj/Ses
2AQQs+EZkCIYvffY253DnTB1Y1+hptLpuQ4q7kBINEfbeZdq85OvhK9K2q8BOOvG
DNWpCGQ/wAyh+w6Ubo4DAZHi/od3nwMOVGgToSsEHxZuDCA9hsy85nlIjpUC0dpb
0z7U1vGbfZAxnE+zcKheJFtCQm33ODywnsVbS+hTlXnaUSKNsD00k3LnylxvH/7W
6xLMpeclvdiwisbltXZ6h8vwB7MHy/zzsTZL8shSXVS3aLqy5eDaTlABzE+eJTu2
oHEaaBEJUmZuPjRtWP40Vx6W+yTMc+j4aWuYLdA36cJZJa8r0dH2sPMqVJWs6Laj
fpKzbSOp8ZmEJP5rQTNgVtEIFCzrOuvUv0vnSHZm1xejotrUSOatYlpKWU/lU1Ph
2H+/LH1TVD1b9YqAma6fwMBWnehGmGPYTJRIn7Ra+o2lvHTGe9CkLpI1a6ufRG94
bdeq17kvBOiMEm23O/6cG9pmvy0crWiv146kM+BHbNtL1c0mIwbzJ8+ikK7gUw6G
JYuJDW4WMdxGEtXTc+z51IrcSi0mtv/bQJLCVtdiYtQBrH72hltLoZbQ10dIUU6M
paFh7UPrhUXQExWKgW2PjUK+x7OqZcyrtkL6npTmb4ndyP/0Awctz/PMRRYC4Y/s
0oDa9moY/B0xserc6VpIcEKFHNHdW5YUs3JY3+TQZ7oEZcBldKoWofwzGwwQJhAi
KIcTE0U36RgeTflrYvDg8J4bvsKqM5cjdw3MLxBwHcyUhk9rK339hSaez8Mfeffp
dcyELYjxx/CB54L9SurNYAkExwnFyUHPlyLUFJXtS8SSrEHRZHsGpmgXQsqv4rHz
LZF8x9mxR8WmfKs19N++isOQS2+DKCD5M2CssQC1qNp2+Ou2E1T+H/9U/QbkpZ6h
b5PDWhL16DW9MSRFGR4D1PAcqr65fWsAFNqEv9yhkUEnoCOEl6Id+iaT0wXzmSby
MMCTDt8OUmBNCo6Ti9U8YzJ9+EQ9KTX2JruLmpLGI6THWNVQ9U/ROkRzHd4TiX3v
SJJnd+WagtVtrVrzEfgEnpFcP/AAS5pRV6ojGeEW4jsLCWXvEnyUcHfQ7DnyrA7y
2NGegqnu7owCTA7nOMeR+leWhMNfpGOtepyE1zGA4Pj9fVr2BsQpo/8mPYhLDpXC
ujzUr7VPJcXsO+5bMTF7zGZCv/G74jl9KyMRaZciB6aidPJrWvXtLS0zV5tjcfhz
DbBijDML5h6/aIVV5q0lHfVv7fB0sshypW1iGM419VIWEPgsCMdVwlBXS849uP2v
+YKMdBHEcccZKaR5ls5NAzR6Xci4oO/vBWjm4tmmJJmadIfgnUonlaZ9lcAMfsbR
4i9zy7TjUIaaiLu29NIEd0aLiJN9hdSK2gsLRZNIPKKHD3S/ly0bYNNpuQxtcs6y
ILGmmGaVaje8EIEyC+DPYrGkoNhOOTUgUA6eEGb54q3935YMjSRjPmpT1Cq6s0B5
BZv4tDLuOy6RdFD9SfnEDYhWs3jgmB0Gb2xWzoGPlUbHtwn5Y3TU/K+N2ZjHDwiZ
+WgwBo+jEq/0FJYd7gq2es8PT+WkPVGevVXdwt3hVvB721NiRfyRoQotAl4HPv2o
+cV1Tj3uazmFSK+k8fHb8xVOxOKkN/adU/MRzM3ORx4zHVolYtSn1juqgOS1WYAg
24qqjKsHNd8EnJCboFekq9uywgo5u7/0Ezpyomi7jCcrPiBDpiRiKD/8+pcBY6wR
sBrQjVUTVMNo3DQ9ljUG7GF3dLxlkfw/g63nb1hocpZH8G0C/xqBN0e7VAEnQE4u
A67jV3Ha9fP4K/li86QnNspG6Nfs64drKO8FscmWxh9pz++HIpXtTRPIBa00QeoK
vGCca+QUerMg8nIXQBe3vZUGe8lcPJ0ranUHvWhWe0HKNLMXB2pzVgZoPkvCbJug
r8HWRJs5pkQ9Sgo9Vwoj9kxb8+eYXiDJrOsLG9yBAczbk6CsQ4dEAcBorPhwizBp
UiZDjQU4eLcQv/1tQf4y/dFDRIlmHt7a5Z7VK6yqqy2bSXhFoflids87Tx1CPbGF
RYWauGKV1Ps6EKXxtlueai1YHLwwr+aXHG7WVCRyI9RGeu+NJTWXMhKq69FE1Ctg
ZAEVUa2sWgcZArWEZe0lxwHhDUue+ZZrIsG2IhckFa1Ko4YFAltWWL29UGvayd0T
IBGKUecDfAPHUyfyLDo1tUEDhHSbEsnYeEaHJ7hwSDwV2WMe9gvoHaswduDuJdqr
ijjQrHxRzC/vJENODfnrXyhQNVuuI9I4vKNGugfINkicXKBehwXaoQmnRT8CMU9m
KIaCDJxdBA/HRbzF8m/hYXQ2FUHf7jnC7+gwka8kWMf0ThexkTDUkKoQ1wYpXASA
QyNj5x5JR5n53ZSuUFMrXR6ZjTcQI05uk9WW57LhN1UVECCApy6ESCgMd40v/TLH
tf44dl1LU43hnOStWAoI1SgJaU6qr878kixJqG0pRcYYas4u3FrPkr1eLrHAXRrd
JE2bJpt+8o6Ua9SZvb0pe0RAT9yttQSY6fA0Au0T8h01Fsth4UC0tgoVR/Vu0DGw
9WoWrzFvTcqLk6HUyvfLCNvRoLEkoyEoOneVfGdYgb+A/Go00nDeSP6tE/FqC3xC
qbyYxn0UVfhF6F6fujvNIEikFMk4zCyoMiSHcTAZo4RfVJhgJFlA3Xf+b7cdzQQF
E1CNrYnxsMPNdQBfXbvI9P8ycwScthj8JqC1skar/w77foFFhD0HDsWvpRAR5XdP
J6JT0GVdNMNaolrojutDpKSrjdhQVknToH0ncHUO4vFdg2X8EVqoQi8cbJuasQno
/O71c8UnAqGFGrqs5Bn8rVlMc+AuS6AiyL7enFkyRm83qpcTIdS5W1HZN5XJyn2v
L3ExhNjl0WkpScUAUsNTkbk2Qs9dM6bFu6P6TPqrUBDZNPCnPiwSlLD0aD87Qj6y
XSq53tvEXAHUujARvAmqjz2Jz2sAXmGQy2DUyaYxnzCI4KYkDhj8dZzpBQhre+94
/5FHflNuXhyw2voCQDOKmE6RZGN4skGSwMhFoL27d515y4TyNkyeDU7xGIiHGq14
fpYFLil8VjEXuVrbRJrTsOWnpLAdDh/kpmdk4zeqL8hWaQDgWW5d8qy18oUeHMev
3yzBgTIbVL/jZfIuilO8RM0xYG1l/0b5M4De2tyJANYJJf6crXhB9Ibq2A6X3IrH
sESdB+FkMrFHqD9K06L3Bpku6RivLlvMhB/AAoiDt1zgEHmka7Pi2HWS9ZvAKlTP
TuSWauF/Ly1XjuwupIMvChgcL8rQMfklbhtGfWKPBU4X+8e5NZ4C5KqJapmnajhe
+EAUZiVGo5ocYeQhXWAEB6CROGdHeEnvqAF5eh3t1zJbFHBmVLj+et14NVdjEJ43
A/vwSq4/wdxgBaArP8Pk8cdKqi+tWJfiDabBSGNK+4o9yZHjcqbtdgecPkcqFEJR
ByP46vJQuE181eFZUjSA/6sgxjqjqVqStKmyg0TFC8mbGJ8BYEPQ8ZV9RB+kP698
n8H/5dhaNr653fbZzL/cyJy6A0koEcT2pytAhYV4PKGvCmBYjozv2nNXQZVTFEd3
VByABi3KrrOdNovNvumLTpot9RdMFa9EWctwPtr9dLRqGfrcZC8cQ9eV1bxmOnQK
ShcNxzlUR0fi7k29NYQIuFJkW8v+j5sonVO1UHrbt7XXpXJyN02uNfBihriU/MQn
V2l0DfWyA5qtrZTDESaIJlQevRPW91kwvB0lixSJ5/qHxSPgAOAHUWC/1+1Ltah3
jZWxVAZdTORbBv9/AijanfE3mceP3bowzYE8U5w1wUU4igqFuipxIQW8SW8h6fsB
/wKqJ7saNJd/wzkdaGyAeUo/33+ssRu7hoePWJO19mcmEHm8Vlhkhlxwx05qcoIH
2aViAfM9jz9SPZbUBOXBvCeHVDAWExapPGunOyfgKQYqrJ2zoSQGUfZej92G2ASJ
wK14C1YYaoAHrP95+7BuEi5mXmcd5Qr1EdI1Vddu5W1kmYKoiJq9mTdu3xmFOkax
tBvMDFXrvy2eD9RMpYTWzT6bI00AHH4Y3mQE/zi6X1sNPHcu7CRWNGScSyJPApl6
83tMgRFk39ucm5QyKLuKvi/MxzRbLEeQ0BJ0285NeTV3ouZ129pNGp43rxPp9Rbt
CfEq0S7e1T40AVc7IkO5f1KdD7iLY3mHkQUyQ5xO5fyijm6irAAYeA+xHjE5oXK8
QCSsrLBqLcH5DgcNkHBUbAxs9Z9SnJesJlj9lFAwRWOomA2IHUXSKD4oYvLnztza
PvWweZRi4IhU61ReLeVddgrdMgj/hjs4AkkHXMLatQdoX+8yIEjPsQLAh3KRn1L6
GRke8/b6MnsCiMUb5N7YXvFM+TOLgZvaeGqWXR+8qMFodhl094dhgGa585uDCfwX
jJOIFBfNbKjvpVSUKjIMi2eboO15YY6ShJQzPXNDbVqpNcuMaNxN99dCSirHCvtq
vYYp9yqP5oiP3YLYkcANQvnpM+3WL2xHExkelim3kMbWEa3d+q8W8HbBkiqUxzgb
WQ7BFMXupdu/MET5gK0IVeUclPRJCWpCzJePdRHhQ3fplMdBHeB+eE4s/rsR1S4U
sJBdT2Q+psx6TnQJJ3zGO0vNdMUPQYj3QMfpdSOqOA5OLc+hpQBGZBcPMkJSWlNa
c5A2nTZLe8W1YLouo/2mIr9pGxXV6EK+YzF668v4LLZ9aDQRx8IsIbyxTsjNk5vp
ZEYv6hyvB3n4Tbplzp4OZYn7JO+efOQC7BU27/wPXbdMyNf8kOdoZDQdbRiR21ml
frkIY6rImY3kOwRJ2YLIGh6vTZhlOwlVxKXO9t4qGcKMyc3IBU5K3ydO/VvzoDqZ
w+iL2BzZ+YKmhQDdk041R9Ndt/LmTOgzUs7P3aD0SW++K6hbWaSNL5kc2FbVTsxT
p2b3QHm7hw2LWu5PFP4bnisZslyt8uyPAIVWXWS1EODSEawQzudQKOMNny1ubymL
e2+J8AzXBiDTuo+svj361S6caFthWyX7iezuyIX4o9GDrXyU9pjrSr+Jqzut78Xa
AMdedj5WI8DvEAI3MNAWSdb0jlFgUi9qTvxCzZBGlGGoD6JCXoQWp8jUTf/opFY6
9eNS7yC39yqYB9OqGLnu3FV+9H84PnniZ7PjvIkeCHIXdkb0sKSZ0vTG77oaPImb
j7az4oQocOo/gQv+REp+DMYxjD26EjvITE6xhDWHERmvtGWJx1WPejl8n3SDsg1P
E6aNTbxCQv2w1pUthgwelvigHoIaHE1+4GEwCABaRJ2zp3+qNy8XZa3b1HY1pP4z
oU9VX9S/ViBYV8BVszNzeu8MvkQectJHjjbtkYgtb1GGwjfTa/gYiABCS2BooOEy
Js8l0eqGL7+PaFCw3N1YvQjDgq1nGe3UdLePoOE75qZl66AKkr6OFFjYpFV1X8Vq
OifsbbkqJWpHSB1VH6Y8LneDUDk0maJD8QfFlnTdkRDw/jY0mNvW2IRPb1MbQW1E
54J2lVRQIOrnE2srH7p4/nf877dAkgqsSsYcEFahLZdCdHuEoeTZ1B6aZZtVdVtt
FYskjzbSfE5l7NqtQCcJuzFRqPxM59nyvVRpoSzHlkhrbKosWRdjuZhJSy4iJu17
kDFUYg5BcBXr7KGBLTy2VciNZCFEVo917BVs4quMpC8gS9oNu52a/o+5XauiNKvT
ZZ6GoFnGSMnV5PbGzvG2Df7XLnnfZksDThBdB7dIc1pd4INJtHRHm/mOb6uU/vdZ
91yrG2PmuDRIYweZ03oywjfb/mQH7ZAw0mHcYguNBBrEXUs5I1pixAJGsvZykdOC
Kvk7oMptATbRg2ot0ypNCxcxWqekz794A3loUY9rn+qHgd3WhYwUcHME1qffqzjk
GnOQV3KN2ATe627zJowD95pQWwy9DBK2k8FZwJxQTTHO5nJUqDZiDbctR4QMIOQz
K8HFD1DkpsALMhGSiccINRDVr1S2wz0VmUPdL2thi1dYmXK4cuQTa/Af3+snEy1s
j8s93cwJSnQGeenZRzlSiZM8Zl8sGtyRPpnIT/fq+B6DGO7HiBqIvd7IIoWE6pI6
+gLddD82bXag9U1AdgNrM27mvQnb+fEwhjgXubaF0xH9TUUZVMAbPi9Z5Gz5raCS
Lpiqz4w6temYtqU/V/A4ZJMEEZcpvVpwC7IVH7V28LfzlDCqovjvDwb75dyRX09p
LgYvjzcIu+PpxmN3q3Fzvkud9FT0mOXmVH13ymlblHKmAZHrnRx73GDAZasYizDC
jeVnxMteNWGlpT78X1SuBOhRxOTbJEGA7WnjSBXiZyUnO2ej6kQElK1p1tJM5Cyd
HK2onS9PrZi4EweEjARq9VJKnANc96YPVMWBi3hFSOv4Tr8f5ouYlx6wstXEYdgj
0l9MMrymEb4lkyN4Dlaml1iFtcI7+puDWHo7bE08gMc5UWuzk50nKNby4iZSZ2u9
zRkoO+aWLqjuCMo83pk0QnhuonOb/G9QPQhaUpN0GTjNmj3b2k9WW0AYSe9aqs4X
gzr8e2hhqo44Gne5qHDl74mavLerJ8PoxHdGMM3CyK1PANqmgyUX4FvjLkDD5D1/
eRuBHKrpPmf6uRqd+g5VN/qeSnQHJF2n4orokRgY4Su/g8oNOXM5LEULgvxjiDxE
fM6tiNsNwISAfsn/qaayDk48lvuIN+69ILljejGVSvWY9BZTMyqDpLtHg0Sa8djq
0ct3rqlcIHe2xWgGj3n0YDjsk/MQJSrW1n9cATj8Tu+x6/zeO5ZOpkuGQmjEIcNO
FWMJFCPRvVGuYMlIjSZNFWwhcbI3m7vczTl5r3batHuKKWggaBaaBFpS0p8lFJUz
b+u9cbxnRv45AKlUbIkyLQWep6F8P2KNG/m0omlu1TymVQ89vp3FyV372ubI6Q10
6Yx8jFi2jXGmmA3nHWzyi8uzVAvOt0xzJ5v1z4vOapzTIF+c/BJxmywRYSdHa7/H
yZXAfwZ0OpromhzRMMV4MC9RJmB2vCJk+waFOGeWp+B5ghjcuMki984cEO4vTLSX
vC7Jeq/rNpstcmdm7ywRw6r228Y1kM973iRAYUEj6MBMsc5SykaBq3M0AkUMl/6C
sl46pHiHlMPvaZE87UGEmwG4hNoJ7qegarGF8er0Si+AN6nCZ9a/XDJ/fhdIBx15
pPLYHZdfpRwZl9+PO2Cqotaqs1n8dZZ9sE5LGVblbOslJ8e3byfndrRyno0QGwy+
+rFOIi8+fPoYB86C9vFFJADNZBdR8Du4XG4NSTBFqB3z7bov2nvoYst2NV3+rvDk
vAGIf04dtPUeDI94RC8jfYs69gJrK8A/whUhy28DJBFShhBqoC/GyAVdgFJakgwt
Z5DMUYuEfUuucmorHSxbUJWF0tLzz1weUH83akESCnP1VxKuG/RIlGmnhAju/GVN
0Ewcdm6ZzDW4bUqm6Pc7gk5ZMKfvDun45/Y7XfjJ9N3Oa1UYKAPvY2ehiAxbyylj
CbgpE9x7rKYXIeVZT6FB2bzHUN6UNM07Z9nckjGsgdPsm3OqpEQDP8w/B6Er1Nt6
w3+hxtNYruu/bCKLosr/ZzRxUPqNIoZ/Cf3M9jWF02jLslo0dIIz3nt1g7UhMOKt
2oMN93CiwYPZmicirp5adQuWSTv9WdP1sfxtfCLqfNj7qtxL93c+gQm38nj3YeBY
307cXePfSnw2vZz9zQ+acOnsordayHfa+cQOpuHig023qHHUAzGfuL5XBKr6kDEG
kryywMyiXiERVwLrVZrp7Ouvk8bZbP2jI4lnh2WsxfzDTvNtV/kawPTZTpqiKCr4
UjI1u9YgcT7+xSmXNgT8kFlP8T90lZqTKk8wC1Qdd5tRLZKM/7CRsSIfi0g/KliL
y4LN5Wo4nH2OjRmbT+lYKVphmL+5YbvLDIyYyBFV1o/OSyXHhtYxPlLJFX4D0lEt
mJCXJEKhGUmpjLyBvz8GIWRYnB6rYdK+I7CfHxkQZKv+/Cr5VMwvjU2+4eJUu513
eXd8IJyK/Due0Fm6reaZvVH+tWAKMpk8xXsf+fa8i/MiOB7gU/48xUM3w3BRqVj/
jI33QOsdzhZZbI4O0M/32aXVCvd/1sRmSlWgec/FhtmwleihiPucAJauuOF2i1yf
jWWmbnCKyLBcDWOZdoF0zaBTtmfcpnz6nhOYldKwsHDNdP1sVlWOAK3v6UVZLwEP
rD3ntp1hcMc2QgibPGCKQP9NEtk5oAnoD/htWlAp9MJeoRKZEDsDOy5ahNEYh/U2
6wVrb+5ihU7eRFyX6/DZ6f/NJrS3Cf4CA8HuNbMr+MHUhNTZkkcKMeD83pB+7CZy
XNj7FvFDlBK4x57TM7OKDyFQUDeS4bOsQDHdrbVFYcNVamtn83hv64L10VAsFC82
dWn9BsLpU3fdhPpQhUXx26Y1DJrkP4YUCpUe2GO4tvz8zEYBhl8CW3pWqDXT2rVf
nAXC/t1eyqmAkMMnkuOVTb/URr3oSrQxyDp3Pk3GGilJRNIx+QbuT91nSBHt1Y8g
g79jCR5dWRKJWm1pmiSgfNK1L14vTRssIhFjh3s8xS/HN7FQxh2s48eO2DTnN6vN
MPYn2eWAurqWYG3damFYeM6CaHu8hJn/iax90fdJPHgLYQ+IvuQuRnZ5N1eYmxY7
XErhy5JIgmm8fOmK8mJXUyQEBwvQ/5q2cuz964mwmfyRi1T6iGwmTFFrqpwWOKeV
KK4cSRZPYRJwbgJOGOy06KcjsR4+nqE/QPjOhIbwgKtmRNi0iienRWfJGBu8KLsu
ebCsz0Pw+x6TrOBXXmNlt3KUp4Cx0j9xYVbPt4D+VtWWLONB2Wz6nHsfqbNSTbgQ
C1tUiF6jl5m+1BVsKUBBKzHIntCaNbTSi0/ZvsroLArbmTaLWKPkNEm2qHfS6m6z
Mg0dWTIZY7VOj2lGTaj2IDTOkRPwQz7o1RVpiqoRDMwB9P7ohZyho5SX3G5iMzem
fh20zoHMLHTYy6yV3u2lfb5DUY0o0vxGP6sd0iIdofG1Z7T+7zgNwwTqI53GcUnu
fuWrLcUZuw3ePiqvSbFUwIMOONhEL2d8Ewto0sF6S9SyKkA1OV7K6bX1QC1MBaIe
YfqNazTMMq+eciVxWmH3PgDnAgRgVo8Y7YNjCUGL+pe30Q+9/ksrO1dd5vhQl3iu
SPJSfArKRzBGXzQinISK0sk1TTGTrEgSuNsA7IlsaluRp5MT4a96fVO8bJ1qEDOk
GIxxmBnDognZh+8WFS7kJ9p8vrsE0i2IIFtu58rrfZ7x3N9LSqPTU1HWTwmm9TmK
TJLfWixIAYODb41FSfVAAkVxFRvyyERGtxGKFXFaxHYvSU02fl4ueh5L1fZYPzNS
q/9mY7TsFYpMLSGn+5MJ3e0a0jIlJvT0nRfcoKklZHZHvVSVLKTSw9dhmDccdEW3
nDlu5dtSHXMv375IC5fwGPm00tvDoVBOmGMxWwHnMKyrGz3bahvYdcqJpVz+kPA3
bMuXfpIvkqDqjF7lC9zE2ofrKkli2xgiPf6pxq+YeXyjf8OHbWwp3XrYmy6+Jsc1
AuHVfjsYzPpZjQU/lkRYQsHnQh6Uf3QNTuD8watosSO8LzLUMjBZlaLh2tazCK/y
Yq/8wIG5zA9ZyzJ02RcbI11xW7bYoyX+z7XnxDGcZVga4K3VkyrVCdWGXw4hGaq8
zXyYBFA9mGzyt2shbuvWWxcUOJ6MiVSqs3Bshy81cJE/rEagLuD7Vb2VzPCfR3bL
RZja+dbK+q+t6G48KwOicT+CRd6v/hwIEA9UwGRs8yWOwZqc4Mxh0tG3LKMyVgkP
98/B7BwYKDWki/R6WJxJjGY34Xx+G78AEyOiJkqAX+BeXb1y9CPmwFClfbPTzQSU
CtEKuYlPbNxvIji7dzOBbx14tsJlYb9a4G5BzCJQ13A5hKENY61Py6IHMW7QKNU7
4rO6JQRvQpRv8sb0dZjMWzppo1pYXPm6gkOq1Mhm750Tozns1V5cRjtPHXyuob4f
miIgSocRJsbH4kljXMIUb7jURj7ntRRlNz/00MkZgPPkN/GVZxTzlZjxj88JCsWa
jTH1kWkwHv889oJ4qXgCEqqjYmFzoenBIJYLNeoS/6wXU+v1/AP+/AWthy9dsbp2
tB7XE+StPTWnGRHiJRFmI6nKC8YqAOyiE5a4b7Q/8HTJwm3zEapgNfXe5wjfrHkt
ub+abo0tagT9g/I8KCDdJ7FpmkOxVGepfq7ScdkeKS627Q0nJhS7DxXU0j2Rq+vz
RPtF2PuNxB8YJsmEBS23w4FTsC/LNVJZoFB3b5kHC3PNjrxWsu5wE1Sr3nRYmE+9
pQafVG6CQGtDn4IXpe1xNaviKGqZDM5XZdLVePkY+z9Ly4ovJrY0gzafSxO5mgcG
nWvlXVB4gz8nYM3xQ9QMorDdCtlPJUqStbkIXwbzEmZeYcB9SLCa4qpbsuQz7jvY
ePHMPhnYfrZb3Y6v84euhTBQlI7m/ecmMC2Q4jXvBopAHn6ijcFbwgiaKUc5xT0y
TTpM4jMrmJs3lkIARagZzyqF6lua+Xctqchlg3hcubthantElxkiWVPJnCJX8yWF
LPhKA5WudjtjqOn2BOQDVI1f4LNgzXifQlcnC5ZS0bR5R97KP+wjWppokOEuqqrA
YO3LuLblwmfX+NZN2nAYeXIbwkt1NRnUfL4P03MQnPOY3HRc8RETZzfKJbjJHNY6
4lK7Ln12c4IAlBkFC8Om9wQ5o+0PK5nNSsKIia3TO796RaAdz9j2Dt3sKgYaggaI
ZeKu7j/4iZTCOoRvaUaky6/CK0Wm1sJvYEu37YbWCBHEmV4cJPfLk+8d5EQQlzFu
+Hnf2DJeuMOo6eb7cuwWNocuy1965NBtElANzlHSfbiohAxact5dWCWlEQJIgf2E
WHKJyfVEi4GUp0NXhPCXPto5KU04lEA21/wTtYQpxyAUEQTypxqbJ/eOIlyfuo8/
H/N+rxv+PIige76OfNJRi+vlub58fqIyxEsocoWgPCmU5i+bNL+qHX6RUe2LEwF1
WuqIAT24b2hQfE/3pCxqy8wWRkMCNKqPR748It5W4ARzkQVbQIz1XlUZDpqJ0Ngh
kkT5XsXvus7bly0dq9CepwA3qSix+HJqiKHmMur/JNte/tvJJihVqrVbQD6cSsfz
R5Utg/eQqDdEp+wlorWJLfS4G8l3n0A4+UEKyMbU3axf9ek0zrAMkV9xmlddUSsD
ifIVoHUPdmR3tvsUUHQA9XiY9dY4Fzkoi6vOISHfJn8D6AK9tnc22bWFmQl7BQrK
8WyE7kGJy+Ocw40ekgUvAhcAV9VtNGy26+ncot2bqsxadjxaf/Klc/tlODOM493B
Likd/Datu+M4QYKQkgoDvrgV39ovceLi/Q224GWkZfxi6UW2NlMPq9y3xHeQzbE6
IyVeLeeL87UeaFeUvn4kCcF4jb4frUHZYkFf01D7b28Kg6YsYfHvQx3Q6+KF6x47
pz3xBcTFSG3OaHwxjRRfU6qaOIyKDn9ABY4kZ005pcXzbWVG9vJKFErxjKAm2m5X
+cpwLQrUEbTKtdKh2gLhS2wTQxtYyW9x21UucJyAU8ZaJl/I01WR/FrQvRMK7sN3
+jWoRGyGp1Y0k1XdlQPV0cxp9FUkH0bV8iTb5NMWhbQ4DDDidqGPn67tBItZ3l0x
sk4fOkBYxrKczFMib5fyb95M2iHaejfFgMOcOJSqEG8/+cVfugcrdkW00LVInHLD
4cDWTWA78Nt5dVmEKqdy+UavhdFNvh0IhiZWTjTTV0c4POQx5a7Txe2v6qWZL0JC
MemFltQ9hISyAgIbCbXOSVy5TFx95mw5f8JFFzf2XhJEosl+H2qUjCWCvPWOhuYN
Pop06gti4TSCqTv7CLVPySW+VjY/Uov7SZoSFEKGWkF9ysGKwRR+REqaQBT3PwXv
ksTRbGfgvzFzuzbuBY7sv0pLo00Y8zOrYHedLXnjzh3K5esYYYAInntc4Iq6po4P
VvgMgm95CODu3gZDMBo5X8dVsoyZWQMRyT0I/eYY+BLio4CQlMf2qKo6hav004C6
/gf7Rs6zSmqdNhWTMaCvyP4RFRo6qJpHOjPQ4HgZZEKVu28hWPZzEI8C18HvYwdn
VKytBqU7N2c5UxMV10LOATEP/rFvYz4Owpy+oCqNdFce64kb7oPO5ym4STN+VDU4
bW/+lVatd03TSlARgC+/Jr4ccmp4BLHk3EugGHr9vtrRIZjVigvvg9bMnbkuHdeH
PjrfiUhEP88e5AV68oy1Dko0AMgMYkI2bZYdYXfQxs+MGGF2ewTuJpsDmb99gBBA
uquRaIS9XRspZcyRSQ2IJPvsvEM+yMzW04FoIVQ0h7j4ylYN0CmBQ+jV6q6btqYR
eABrM5nhgc+E0zUo7dOZK7RIt4rMjB0io6kg3YWXQ0Wa4TCVb/CFaLTkUZWLpVPO
OF4I1Dvb/nddqt/JnttJ5peYo0m4M5Okb685mYZYbSIZIAcp1b1X3Q2iIWAFZ8rb
Gl4/3JtkOqbsqYrvKo3v4CmZ6UsxRRcp6VIF8zyyE1bLnv7/OmscRGEvRXDA2KlY
0J+6nZ/EUcvbtSbCKnqwlknv2Ku5ZiEodBn+Ui7GJgnltXPW43lSy40zZDNUUkmG
9ujbaO0T9v62heXonHdeMXUSD/B2GnUPkHPWKSlX/Cr/paz5JgkO5Kszg9DG/zar
aN8pOzj0i93T1TJFherJhcfIn+KyK/baNeF6ac6ct53fO+r+aYKXA0HEiM8P01G9
Vqrmry84emUNgZlW3hHeQfSPJDnCi/WvNAUXb3RTK0wxBipE1o2ELYHWt89BU/c0
9yIex2PTsvK4OISEjZJyv92iTbHsErbzFBvtdlzHrGh542h5t8z10aCPSK/AdmlG
3NNgohB/pqN2eL4vDl9LD0YqRs+3i3oUiLO9TD1JF38Ah2dR3o+vcvx/EW8ncPa3
ywFkRyy7vva/UhhTeGioW7bMHuCuuaNKEEuetxeWjfPiIFTmVToWpPU/x9FltTgR
sF8gyVcDZuuYdRski4BsdJKKeCmEHjtISjCu5fpKnfsw7F6doUe3cW3PzkXR1p5v
d10cUDYnieSkZ+kozpAiTjQ1YY1DCQ64vq0K3sBBq8t2VVmIAz6gLt7b3xcqn2v4
3UG7o8CGUGPJCvQ4YZc7ABculTuPz0mlu8uE+3A6w6l2YC+o7ExiAR48eaIB4sgJ
wxAueodePABnQJT8qJ9n9fT/U8Hw5Xhkc0FvIFySeDBuPeuWeGTRDqJJMJNbhk5i
PHdsY55VgvBLUK7idu4BaEzJ7U9UQp/iQr03e+snojYnZcBsCQZNzlT/AzcZnqoe
5fxMyYYkGcQbIjHldihnD3kIoDc9No724tRLNhJ5JWkO0FjosPMM9XACUzhgxbTk
8FItVvP7ZVuFCyi7XHApl6ga0ioM4D0ICKQTSDm2teb4yRseHJe5VoOd6XDqywCG
cjx4CXpEqyw39VYeeZ3yxuacGfjevVPrO6IequUiz1TSFBBrDW7jtmG4qhYgRqf7
V/Ik8hsTImopqpV8m8ij+9Fbv16h8Du79+o3+Sbb19A74UVr7+hBs2Yj821kRbfZ
rwLaQfE9g0nWS5SQOSE/OPssGe8GfdTqQ2JtXFfhBAY5/wVNxUW+OF9kWU+dj2qF
A4E6PB6a1dB2BXsjxWC4oRsbmz5dGbvYjPDtPLKzZtbipls6hE+ImCa6mgr5FzOs
uaJ9AKu1NkP6zyCWK7fzxZA5zXnUooZCVPU6u/2OflQvaxMq9ekd07EzYEAh72sH
gYjUo7Ix1j8862Uh5QFL23pbT0F6bjkEcb/A2WbMpa5NxZ8Y1n/nqhEb7SsdsK16
GGJtk+x7LLXftePG87ckySu2giitfHdGR4FD0lX7+haCxC7hdfgqhuYXP485vmZ4
Wt85+dTLqOqiNzz3O+P7x1SLLOF6VIR6QChiNWQ+gkOhfo0HRMQG6gPRStXphk+a
nFZqeatVz0o1FaJ1n9yDTyAOBbtlOCFTNW76ec2LFA158PqGw00nVDRAIwVaParB
ky6SrkQo4fhnQDjoy48kTak+MKsGwKQ+x+jjQo+fOfhd0arvuQYuvCQ9OMKtqXax
326E52mZnPqvKwY4zKD2nGuuZ0/1C0SBieuTBT2DXC3agcf87uja0xYEL8NBRtb8
7dwJ1xrPL8h+s7+DwBuFCbMfSO02cip0F4Gi45+Qg7UnpvBBpGqgb1rMgb/tD//1
4ID9a2hHLfKN8fkbgy/ArS0OuYEP2KjzU0YZQ/xp58bM8u61aFFx7fs7nM6ifGC1
oVzA3i7aM3u3kYgiW5E6sURZHrircC+HH56aU/mLazJK4TN+5qXRAC0qe2ZPuGNq
qZuRTnQkhGBkb4i6YNdYsAXMez7E8v34oAbSetxe+FAKOx6Seo2Jci7ff1iueMH6
NUbauQQabJPZEzkB7XviDRowJEpKFJHU498lHKiMgR88XFZFtLgxrLKEWZMcvFns
PdeB+LO7GD0nZXjyIPzDZpNu9RE0amjYbwv9PCo1aI0oLSI4DcPN0VmEikKWhpK8
Z5kg8HUJ3VqxyIqx5boalQibavlbAqmJ17EWcnYeFXF532rMDEWbhp867iBCdTOL
HXEAum469u93oRY5VPQ2FaeISw90eFRgPe9Y8Jk+dfy98tmjezY+oSiyA/dvvFLr
hvbGUZD9s6k9OZjELnuKblCEsRnpeQoXJPPdeIwr/m1nEr5cfNqyQwE4M1IW+C21
tRO/lU6gLaEdhS7o09f5Q/UNahFFJ4GSRjssDTUsMkJX8JcNdj9+tQEdnPZvY0Xi
PNliMFsx6/FPEBpXPZVpzan9RPVfmNtKTwkKiPwDM7AeOVBgJPppduTlSh/aIkGC
PtS8GOEKjmCh+JqJshh1SBR1YrbgnADBbikSKFD0ee9cLVsml3/9q+wG/mZC+Qfr
j27f3Wqg3chUTV1i/S0xWMIpnO9I+ST4CkM4Mhtppe9+rbAggu2GUGyWOEFdWr4n
TgotVSpnCDnAoKlUkYxbjrRqWrBQVGAj+nO0wRUwplKfcro4nyfe2YkkQSXkrYPh
jI4DtaflsNYgGTxw5/PmUxUMlH7NdLLyUgDgbduqJD3Mwbw6VO3nQ6pfwcuj5QEZ
jlpbEfjQH5uZhkY0MyYDhz/6DKFQCE1swnSyfuFOAYUT1Wq1mSAui1+umHw8p0Yd
NTctsVRKBXiv/TbYXu3TJkVQCqlMvP27mKQF8HuUAw35IsB/b371SnNp6zjd3EMa
wLYmoK6ZtQlNgnvUQ7rTcbf1CM3iplcTUKFEYOpo1PPrQpQr3q/YlrH8xdjMruC4
bHvVdc6D3ve1awNZAcOMwd4jfrFK0EqEVkRvCzQ4PRiinn27jB3Uei7PLzxcE8xc
yvaoqokyiU0/ZVbrufjJ+7DLt9bL9M9/klDzkpj4hqO/AG/Vi2ZI3OM6Fm0Um7Hy
N7ScgCRDnyB1Fc/n4FMt9Wb3SaI8PubJ0d05mjRtVt5slBd70FItTYuiFZn5FiT0
ooAEjNjH63WZCiC/ye2WR1IpaccFJWRMvtx+h/oGxjxGYD0vSKuBCyFzTh58OAsr
s8auk7z2MaVreJBiqWqCSdx91S01uH5a9uWifwFgITcJLjluT4yc4RoXH5oxqw3T
vsZNfzuIOlO9sD+TyEBkoXoWFaq7naCkBXUxhQHEe/DMUYaAivtDcqcCUjFVLZd8
4r/chheIfRrQ9/6k3c2jcKZdmB86ODEVb6TdIM1pVjEzr0WMZ9AnyaWxPila7r4f
3K0N4O56xTbrvgCqPlrn4cUFIjeXGMUxRh3SwEsjvgGvkIfIk2vgdDV5J6D96VD0
BxLLe2vGeUTVnXxj5QlUAUdphc6joUdEFGtzMJcUyH0ez0rEZo0PfynnM7jRqwwY
+06JTMSv/AloKc+8yoDKEKklvtJeLpTQAAfPNvFb6BuV+X3nF6n7+0baPVbyyy3I
ZdBZ4uuNXFpC+ZHICWmn8weN8cLqCCmxgEQ52MWY7bKoOZOssijQVRoiQdqb7ni9
A5PH7EcHA/E1BYZ2mKBmE4GmGhJ2JmEoEmcDqDtXPQwi3RunfJDoTpau8WUaa+Up
VxRjMHLiL11SY+jCzNfWE1QJn62NFgRJNRP/DB+uyJiOTtNNsxZHeetV2IOZGHCE
Ks4eflAn7BN40r7A9th69hAjCIfnlfte8Z0AsiEfQDFxuJY0l1DpVWspwZSvVH7z
2WQsMIbIRr54FRvq4EuWzryGgfAZCT1tV98TCYjhzZ+I85JIRQP+bjjGsvqZp4AI
KIEOQhHS9jcPz+1uRMvRZiT5wqc/sJ+ivtly8j/qyj/fKcnGnESW5mbw3sF7dAmV
OwuuQAqrPVTkFJVzQzGWq4bot50YkvSuZ5YB+/i+LUD2xuQJp+bD0GFM+cC9T0bL
XnbuxZW+StaDF2zesZ3tt5EY7lw8Ac7ZbBq/JG3ba2RKR3JN9VkD5y5Ln79nlBH+
1a8qhW/6IKaPpWhDLcNXSoSYb9WC753pyeyxaywtxdnty5n/aC9UAvNzrSHrdSp3
O8UgfJtclrGLbsR9aSthA8QpxhYsW53LVjGf6ZUO43RYLihcNUoc1cr/6GfKpaJP
pJKMdTT/9MeGQgZo2X990ZADG3aYTOzaM0cYWZPbzuDT3a805Zt64PD5DMD6BZOB
yI2N8uyHqm9aFntNYibqs6X0czBmgqXOAgk+0GyWTZ0pHWF0mY8BnmV5xj9StpEL
diKjjz8/gkx4C/CsEeRndPz2LgEBbVLBR4UTYfdoPhGXFRWneTUKNwICloXSzbaV
qYPXN6Y/GCQaThGPUZNHAmakba0kaBHXtITfxwWsI0+K8F/JvqwHIGvYvJSXXSj0
jIa0kc1NQuK6zbhyLbPUv3UrrjPVYXPHq643ju2+dx0VrUVOQkoYJYOtt7M8/Mu3
mQ8gaWiHBh9oJaGLmWjN3kTNenVqmvv/M8OGTeHzVK6JSxzXmCn2ooMtMUSwWYZ0
Pq3iszGkyXwbX+FjI6p/ZlplKPSJGyGOFAXANTXfua8o5kLQgphhDDG8ACjU2IRG
eNnywMY7czogbaU6GsxFZ3Nf3J6emFgoP6npZnfYvNHmX4UGq3+Gy3TpbyDUfYk/
XQmd8P7ZPYCUVklsaJEOgF4JyFErWheW9vdL5+VB/OCWG3hJKUGNbbRyiVCKpyWJ
LMlm0POOi2AJxk5w1qQyPLLlb178jk2KcpivXenbWtMuNcWPri4Cz/BNBZsnObMR
LiSwcZ8L3Tv3tei5FuDVS/NTtdNsEf0uAXQpANNwGgak8ld5zKRKeaoI5Pq8+qY/
puNZyVudhjwoS4McLdKgJ4kRN7q/yCl4coN+SNrJs0+szlgnHh1ymiOzQV47QXFv
+q8uRH3RInFOwKyB3tvxSeFFFBAMDX7+qsbTXkniD0NX8kPp41N7eBV/YAFGwi5q
29SRQvEkeEtkgB8Nce/F1sunp9JRpQqbNF27Eb3hwXwH27uNNzIXJ+0pE6Bp3dbw
qLy/zFw1spDRoh5GkKFB9KGn515XX7Fxu0JgBdh4b5ukETBmXkWuK77pfx0MguFW
jQF4BcFm7A56GOkcBkGgHOp/ijJNwvyDlYl3dvxDpg4+ICT3TzVjXi+X2DC/lXh0
oWkenBu55eKycRx+a19w2AjiDP7t01cuXAgUHndVYNXO+NjQxSo7EKGlwRTGOA7m
tF4T8YOUYrmnmKggDy6NyNk3OLeTpw0jsswoIwQ22zZVHEaEtRP9mveDjmu12xGp
aTIyRBg5fDqe3FuHKZ1hg9FqrTeU7X4gHTO0IXSdnm/iU2O0o18hTNLwA0f670wu
l1rPkpAcMl+nF6yTevRjCtUUh+RanEOXUgj5hJSpv5N7sLAgzxSEb2aDXs09nqrC
TR/W6fN8KFlifJTRa4zB7glPnWh71oL9cLZtMXqoiLuWkvUWk4wY0Pj86LcGHI7c
DrnHKWHYk32bNgA1KgKzTiJzkTWJYE57WnAo05N51Th+xR/dmVx05JsyJjNwB6Mc
72KjjWEzetTUjyouo61QsOO9hmtF3HTSQCawGGoOTEPE/ALXjF6KMMrBacQc+YH/
hg7hVwVHTguLR1rgvR+ua1wpH/0g8juywVRXKeVoE2OfOaf4poz8hYk8WvVm2G0l
SqAWgUfNau2TKnjmLXQx9oytZ9hc3vG9xApLcYlgZhOvC4RkZR5tmWVf94rSePtr
jpp3v6sM7+7jVsD3E2WHslg+cpNBQsX2AS2yfUyXieL3CgduxrUjSvcnZajJqQBG
+sFxqtoMAhZDC2tb+M0IzLIBHDJAbKTIsfKGnaE/7QtG8tHdx3oMknTHPsf2nv8F
PAV3p/naVIjI8CaaqkqK2Ej6kOU5qYjUeggMyiEZKxNYN6Ge7qT6W/4Pxaf9mzyM
kIwgW6t7GegXVWO7Aq+y9YEBz+Qq11b6PJpOoM8qSOWsZvzlYR4fLNrW9nxFCU5e
yYSFsS/erwJKEn+aMC6d9fGdAk44oxyyk/vkVEVgwmN5MaYCEpaEAzAvC0UkjOCq
VxYD24jMZoIuxovB1aufE8DBepSBAaUTiqsXEXI8CZL+BzQZhLkyrYeJk2VB7+QO
4/kg4EZDylG4yLN/KMasxr0bO9u7Ua77nc1mdHpomw/B0wP9fGmrpJZEDvdgpF9i
Xu2m7RIuzpv7g9uHw0sB4KpOjEXdgOCDExw+67TbCiGF2WBpYxpe88Nd8YDE69dz
Kmze+h9SXa6EyYpV9av6J8yyMPdQu7ojzYBzJKVFi5nKcgh3BU+mSP/pwA95pMvO
VcWviFGpLUyUYAsBowrJChsVZM3Ns+Vvs5aYjMxRAVBhzRckK9d0Fy2kO2ZC2xRy
vtDfXOpNwLz/Z4V+XCL1X+okD8azeuq3hZOaeTfvWSihnCEZslWghOKJbgNihPWG
BMF1A2tBhOSZ8ZaXbr45cYy/NALUQSm2iUEg55a2J/n4k6PZIjWKLof57s757Kqd
XojrCQtNKKxmBYFWD/OL5xRAPHaM7j7lk1bhDn1/Xvv8AGOPtIaQ5Q0F0mxv5fYu
jX/KR+W7P65uT82Yv3rZaec/42AUwyOKesnKhZ3QBUwjMtk0r2gpOYQEnsSHGN5w
IoHqvkRfBx6gKdVch/sjspzGhgj0u9j7cEBKQiF17q89ccC7HnQkDE4DF2jbIVQD
276R3X7Yg3ojna03GrUpwiXK9pxvs7mpmWeSx0jpIEj7WTt4G/xDOHd2S7eQZIxG
QCJknf/n8vRfKs9XfTNMMsNO25TQ+cP+8mcaW8UYnhQFHKLqlM003NmZkMrZfTiJ
4PssrD8AfoIuZXFCblhc4I2rZrx3pUy6UkalXQA5n83buBo7mqLT3B7cJDRkEzCA
OCOS7V8XtfK20e7+OBsSmonReI3MICU0waXMWxlbGr9hYWvMWSnO3dyYWrrkjbPy
FtwqcOi3smo5RzWB+E3/orp7ZpJjkmAXXgnvlnVJcFFxxJCQiKbpANPY53r+YuDU
KizWj/yUxfK/etad07Dr+iC3KRHJzAJk3SNK7A3In7BCukcuGv79FGrWXnzCTqw8
M6InI5ORKEt+5tdRRaNxPVpXnyr/aPtI3f6an/WiVjusYgtX/j1soqQZp25tPco8
kdPbufbyj2WPrzTL7uVlbqWiq1XKsod0zp1BsQktv81FQECN1apRR2lYNZryJNZS
rb+LwIZ54yK4vTmLh7mT951Amt/hltm88K4BdBCuHkpZXyHsIDytuwkUZYpA5gho
R8tWXzLQ66UTTJZJxkmvdS8fhYkuLb7vXS+KDjynP3FY0QRiOW0ehalhabXHHK/5
O8AniHQFYGPHPkVfXMgC7y2SaHJEf2/UJ1HltpAMo2r4r3uZa6+Fx9u9RUq0qd1l
eBPD7eryzMlH2jwQ5BIxBN4YXscEYR7DR49UhpIivGoJsb+Iwzz8zMtmMIIayEqQ
LOMwUPuknVFuo9Uu6cEeZ6Tc787L7uMJMhWxKHTRRdE6sKD5r5HoBF3SxD8tBSEp
Pz6Ochz4cA9FDlWC8Oe7dJ751FO0uxU1soI8pgacFaDJFl5bZZZ+lhIwnd87XxZe
gAOWKDbpdgQgo8wX0u5yOQQA1hmUziMl1DDd4rwZI/eHJOVfhVLDVWR6YhRMT9cN
dqU/sj8hRZOj52v0kci15ugKHibHU85Pde3Fffq2HRyN6uxWsp41WxYeuu7NZPRR
0mDbrfutCmYlXFd2xlj6F7bXjPAJAce5LW977ZNUdKUP9vEv3lBp0QWCMIYtzfif
DjYv14L5WfqtiCLH6zaKQHxhC9rQAsqhXWIpSTxd311+no7qXyvX+/60zXKUC19E
sxkbQVfwR7K0G6xUP+3ZcR6djJQ9ebr8EsgqAtGuD1tBgrVJ0Z6IFEuwHdoiE8wa
+xEqNi8glLgtGcofTcp9BMowEbyvvdoyvohKsT//VTZCGQ639cn1cD/6odlsliER
uZ73X7pfKd2zs4nmAVUxcrL0Gm85kHJumq4sD+ufGrzAqK5TeKyZo4PoeTpUFNhh
mebgF4C14tNm/lAntmrecHeEIjBWCCjygEkAKHzQrCiESsR4QKuC2MHckL2p6iVD
RD8JVgeetwLGXHIMTBfkhqriNSqomTHgxmV+9I85ZEnCLlC4TY9lbP7MdxMEhzXF
StgI1Wg0AaLOGyMRGY7xIGvWv82QhDE76xW076KxzbT+8+gSk1jE1npS6uRN1g3G
vltx1j3sQ6R9rwuCysqX7cJTwEsAPCkelTcufH0BYi/kBpGiMXUrym1aJAEgOv/I
7GL+Pl6wWRlvkBQI21WtedPg8kTkUv+3M0nYTTWXcp0HTTwviWkVdCTjHW3TuRRm
GiB5K5rlloW6LCPhHIvM6x0vznS83f8OIRmDJAmPft3xXclmhOrbQr217W3cheSh
39orxa/W49IA8i/qoWAB7OWBGQ2sE1GfjLoLqT6jsHqYQr1SRdH6Lag2wPTlm303
wB07t9qaniQB0RsR02pMlQkBqnJcsTCry5LVBrGDwcmy8fsM9eKT2MtBjHI39X/p
BoFonf9XRWQBPQgHF7C3toWIaO2yR5vT+LE4ClruPGhspsMff2K44iQLe62bBgJI
gWJ19AHDNuH9TMqgPVg/qwLACa4vDQGG0oYFTzA2o0V2sje9y6dgGycQE324w1X7
JF9MlvNuHVYPKZyZUFBRDMu3NQxMeVdkUy+Vv2pIFeXa0dTGEo29mfsyM4amE75A
6CgZG86+27v66y9p2/0D744UAwQsqhAXba6tAcc8IHAf84ma121LqVx836tTTBYM
5SffI97CArHH4kzFAg5LuBAZGmWCx0izoqcJ3NR02YpOzBwFL+dLybGzcfZXibxH
bz7dVxPmErnhqIhk8RnsAarfizyDnDRyRVMBbUrarcHqgYrthNeoabsCB63WPsXV
pJZJMt5J3whdjyFyEglMNlXSb0ecekId4pe5wtWbisRa5HDuYCJgEjsn7h/jzRkC
wMABC2EtRZp8WdPiKh/gi07AGMNiPTVGH2gwU7NLfJjTB1A2OiK+3WPWln27CeRP
bB1Bz5SmNdYoKGmHxz38YRLD+Iip60Vsb4erYcuog1d7PVQyG4A9fPnNQYUELSoh
BUtlZrJZUAd/Saf9U3jP7UNY0cGhqBREvWzZZgMw6crGZczBYZl9OcpFkUEz8TAJ
pwgHQAQl/FCKaShnDAHD0Hjon49iY1Cx27hhCkNxB4IlE7CSpP57N0enFiK+qw1/
+B3xvwaLewB6AF/eYKIniGty/QfzCxe7NqqCgQxCJpEoCR6Kp+T4cUdOwZ2bU9wI
DBs3moNU+WteJjhfTgDC0Uy0HXcu5umNsXvzRHMHBRmp9StfaCPoLSKgxKlZ9oEf
MfEsh2OT5tNeNhYBEnHmjXfk8GQ0kSwFqzyUhayoxW2d8Z5S2idA0Abs7ESclO8P
mfecy+d5Ors+mAAylJqgjn18IoqCwtE5jnf6tJxlndVP3KFLKH1KbjK/5JIhMphF
j+cm9zXrW8s6a2j+vtOQilEFhgWZG6dyLJZKcwRXgQ+pFD7xZu6Fstz5Xsg4bmXu
Qi6G1ZElL9GFfLM+VM/51WjO/OMZlHhqeOiMWZppGyPcHhA1OmQiC+xdvtFFKcsn
Yiauf7NSbz2ILikwqTwKDIIlNaQc7Z1XpmwrKlakQlo1sW/S0Ustr+OzBrU52t4N
Dt1sSPE1QgVVZS2cfyTrRn6Qcj0KUTkeStSPkEWSmqCPSe7MpAod2joKUyDAgYtQ
la5QdF/5XBcDAd2vzmgvh5Ls997wdFFj6I7pbOw3KRSlhh+L8GB/aSB+1q6keYyO
SX8VmIexlGiYyVQSZx+xCrpMu0u9rva5QMb1IqAhVRkAATG9PVqTMQfdwAEgs9sh
Xs5eInuJJ/maYKvHxjYP7z67zml43SXIu4mekZob2mmbMRTb62+/TWrrWzYqrxcu
WfF3n3rC+9vCQG+/Fpu+lwRkdVqsPXZZNiqMeK7sl28ltY2g4Oy7n0YRnonSQJNA
5YwltbHaXGtMrEVSn+uIKspHLXPXiIIymBcs6pKrZHLBw+4rHl7IQ8rczMS3nNiO
Y8mxjg35TLNkUK4v1tY5iQuuBGMQBeZPfOyaibugBMUalkx20YrzNtgcccY5o0b3
A3KXHF5OKVH9mN8Gk1XE/KWn5Gk74LtFZfn3G2y6VAMnlsJUxCBNxo8Z4PMszDxt
tP4Q8kQ5fubw54jp7BlcgEYkSyrRw/DHzPNdZvHw8vuIsnEoKqdNVbrGHUMwF6QX
LP28b3UMEaGjYRdvMsotbon+11muir11sZpn2rtHpeOFRlLbRIkuHrzK6XbbvnOD
JuEE5IR+x2TL02+jUb2a59o8P/dS63Vc2DhOpxFg2oqLS+lVhi0tKIyhMtKxNrKg
rEmqTx5Wsq6MjcBmkDCpNwzLOzBhqD3ifvFRrPXKTus7ab5jnOd26uDMtVPxL+mt
lsbNJgSHAHB2ASOUl0I/W4a0JHD7CCIL6jqM1pGFKtZcaDzW8893lQOdbZV0D0BI
cCwaYYn/7ztz723T51SSIIcTYVQ8nWeISOS4TWHlxwMZf+PZYVovypAp2j+AYvd6
Vgr7oSTh5t1EFqxdznj1z+FCXrCgxlgni9NLnc/O6Lgt63wczsxz6G7HclB9v3MY
uFw0ZeoCfUItXdYh9Y0Arsx2lPnpmEsZ/Ob/mXzDEfJ83AJ3ceQCiCT82CnUPDeS
UyYan++en0qbSIRsfgDtqp3bs8N7vMdCfKSrclK0waCcMjk/YalgrttXZP/V7PQN
w/mU9NSY3uPyl2uxrZTae6hI2MAFbBD8SRevtXPyoggLxxx5/kvD0FxDLww8WSur
scqnYtHXUUT6jXTq0Y8RLSzV6c5LgThMlFfL4ENSpEIE4dpmW5kC/lwajBBDSs/f
Z866RIr014dhGoiphB04wSxiQJm37q+Pvlso5p0DOQvyWln0R6JXtAoNyhoNnJ5j
4q0T9noiyy+JtJbXYceFXIExoRpVrc4rHsoICLMVcI9MNslQC6uPbCrRVvcEWWVR
kJKePrwuO/BbE/S7ISMWKCdexvsy3gQsAfmQhhF7J0+fUHADZVxk6yFM9SVvp97R
USHoVpY6PfkY2sTm7fTmmhozDvM031/K1qMEAn2jAFrWM120M7E9gmb1yT24fW0G
zlfo8pPaHKxzZa1lM6lyvf8eFQYtcvXjA2QWgvaSa1dDcZjo/5eqWrHZSvUqTtMm
T76aHQemqhh+lnnoIom4GI6iK8aGrl084kNtMxYIkkGjOQeC3rU+EHfFG/M2PS/G
aFkws4Vk3jdAN/DAPN9lF7EWOfeugCWlRGMEmu4R7SLSZXzzn32co1b0r0/h7pbH
RhcC+pCBdM2YyNXjw1yxk0cPJLdD1kFQjVBUSdKTEs75zAfU18L6EguHV4riuu/N
sCF+AhqmK9uY8RA8+u04hYGdDpPvc+f3MI2oL3uCBqZXyUI4onkoDIbranexhKwv
hh6azE9KpMZLCYLI40L400iuMkLT0aaZFX1rc//cAGm7hEbaZ+uP22V5eKHJP0RQ
mTkTEJOeOs9rIfYpNK6QjvRKHmQMdUd913SGQ0HOPahmvPhWQDKBd4x2xoFN4etH
k8HJhqjHt+MJauX5mGQVNS00vuUXhGB1moasLtx9X/HGqdG/L9ZJqZwqzmelbCb3
40WGAkyoQVnPxMiba/sHVEYsjBtsY7o/tX1QhWOP3z+NG6vLdFYEX25ufP2v78YZ
75dIw1GXnJ+GJLS+Zeoo+/cXN4AAvnmkwQ+5JPD+j+b8KnJX/BB5Y5T/xLVbEXB0
ox+YwFjsuouyE5At+dLN0N+e1iNHbHLIVEmPvraFH6VNNVpxbX1mfVYAhJ0+k/Ud
w7TwoX5RD+bywUNTGJWb1yyNGdQoD5H8kJavwTc62rqqUtlZN092FNJ2aHHdjHeB
FAhLK4/WqIs9r8d8WLa0AXcFYELMQY8fnUD676L8rr3K2Nj3Bu6NTGFoTwYVqfcL
zi0NncDkpf9GAE73OULodZf0hWn1vNE0ZtPNgVbMYQOeBj6coXeCnbdvgArVtTIE
jBWbKhdO+pYtmhLBBqhbgwQywg+zh3FLx4AB+Q/v4CWb9c0KjzaYrRK69tmRmEng
SM8sYLw+iI82PED7t/3wxst2qLmr2/mSQKXuX2HofXTRIoKNbhnJTp63Hp7L1B61
TPPU/evqzX3jmffKggeHYNYIALZDOnutLH1eO691D7zHuc5Be0euKngS2BCCogi0
6DpBUfiiSMG7lwkpT++n7JZi3LK3AEN0fBUXFdwFwr3P01Cww/vJrQzZ3VkbbkGN
yyE1oEUdg8qj8xLILGzEmUSG3auZhZVhNyZzhmNOROo6ywIKAfhmSi7FdZRU8beT
MpD96moKreKwhy3ALpzu0uzMKsXe9Ei6eEWjCyYlwYGa1PHOd+4vDp7PcbFIDgNb
N5nQ2zcXa5cv5roypFAPAL7/VKZN1ejGuxCECsGoiqaUhZhVc/Tg/uSfI/oZ9jEX
G3fw8Ebct8Ut6SiTL9BYo7Bp8ZBFJMYNjndcLijYJ7SIfMjkeAx6Tpu8nhzJ9E/J
UL7sgfmeN+GJLn+BEYySOAS+5RLOr4av97+46CjB9HPAa88dySVtkSJvZR0mF2uA
bbFckjP141CGP/EvVh2mD0PTYRAGLvABLoj9LVhtKI/q8mkwlktf1F75pQJwRme+
qvkvGqVCRXhjDFjRWPEI0cnZTDVCEHzZA8KxzZSj1II/s8CvAhhrM1lvfgJoC+Fq
xrbDi7USobDowTIbqDqLsB8nmtvqGl6oJyQSbDkHfRhwgwieIRITIZ90uUr373C5
OE3cSxifo+A9JIdAT6I9ORzopOKE57miy11RmG9p6OrvdxaZfMIAKUWNn2I0+O/Q
VxNJOXWbZMyC4XDfxVAzUjdXZYI0przQ2AQxPva93SCFgUYSSRXNx7dqh+fRhoKv
3Cv4ZtnjE+5fvFxNd6MsYxFXtCHNRZqPruqmC5BXP8bOMBgRROt5ie817r9dZd9e
NJM0bK7BiUR5dTgyXPK2aKmBtbTbl3L8zOEs4QsyBmxfg9Ae/0aa1gFlgYUmazC1
I1cuva5eOeeYxnMsKQPFxJNB/WzkqphlTJjAv/Y+rgu8retv9zEwAXOGMP9yiymA
PKbd3XScNm5KzMj3ZF2kzXazglzoUmmpHlQCUor/3l1B/5l8O1nTManz7zWuMPpZ
H2K0c+xL8cwlXq1GChU3+9YCtBQzpXWulS1vWts8NP+LxiOJ12IyJuol+T4UMuHg
Z0q14BjwNhLodcCT59Cvyw2Vh/4zuGSD9iHYAGyH+2+uQc73Keax0jaqhdZp1crn
ehzjyXm1ah+3yoNW0vq7SYzdvRR1ned8/qFWUSuy0HWqcDl+XGRJndsB5KsjPReF
fq0skMHyp75sXl/z+ZvepgEkASWgB3cYPrVh/IYZUMo7PLQouHpN5HfKZhDdtIaH
ccgkKf0UJjJaVsA/v+unnSG1jNm3vS6LTut0UR48JYUtiNmTG0CrbatqQdhbUJDu
3lgpMcQGeXgeIGg3pNBXQPF1J9N7/JpvOpASrVP2qwmCCsvb8XvvYbGjOHI5nFMq
w0QG6f1mi+c3BwcktitSn3KB6v3MZKxnwoJxiIioea2h0aj4vk9qXkCIT+5mYTI4
v2iN/oVb8tNlKUT+QgBecwR8JGhp9ok9yONG407VeVp9/qQLPGXSvkRn2gyHhPEr
cUVfOpa7dLCAnuclYUgpb1FD2533cGkJOw9YFkhRDqPnec0ElzUBA3P1K2oTJ/SQ
2LmNvWc9k/fCkViIJ9Xr7v7X3nRRK+lQGoSFjUX3V5bFOH0Vd9pi9SfNAStf8cZJ
WlBVRoiIFkeixZForRdvrtTl1kx+2FZtdKPVnHt5GoMqd4zIBBPeFpl+nl4Il8mr
Q0l29smJjb0YaKAF47l9Fgv2sRcIYIDVftRkqGReOlokn+02J7F0eCK9Zd2UwYiC
cguTvAd7uMNnq+jggB+klF2AvCOu7sAMk5+S9GgFpS/1DcnpghBJUZcFW5xMWooo
xxyrTrXgAodeuGuIMZyREdX3/dMR0a2DOYDp+C1NtXuLAd0umHIsg5ipVzxQ0pGn
Zm93GFjXcsDGCpHBbwwN5rbkKu4b3wnnXjxZahLmYT3+r9d3vL8jEiaPZDblNhGf
IXCcgqpYWkJ/uNcWCMVZjf/7Fm0Tz6V4DE5x8Ds2Oq8xpcvqsk64WBkf3Cfk4a4T
EuWsvV0V6yTZDgrlXcW/sAeboJoWb7JvEQll8bTsTqnIPzAxmitQkjo5NnYFBmDA
l8y2/f1oeGXEi9QHKLvzFUGckj2OzI7oaRsCnowuHD+KG7oIfLDFZKkB9gEWdUne
FAcI1DOzavzEChepuacQo6vjM/67nN+5nne/02Ykr8g97n26io0OtOYItftjpPAv
12aA21h2+hKb5JwnhvnjAJ9lebdWBrQEWFmwtq+2k3fdT4mnmr6EBqvGk9OteVSX
ofjqFB7VW60SQqT004gJKo6IW0DpTL8h9vkxZkD8wDgtrMY5LlCzCDyacMC3cGUS
5BW63vUFXj0SslnRO9yKtyihTzV96pUE7+RZsvfUrGRQH1a7W3UukGAnKlXrveKQ
zILrP16x0zbb+JKeIXrjFGx6Ombqjn42Kql75rsossXSURkgGEaSPhvWaMa6LAKJ
bGnbRHbGpKyJWmBGyrXvv1vZ+fSJ/xQMnBom5+lFU8Hq7HymDK7T9IwJ3F3tAO78
NmDmUR1b3VzjiuZ8cwD94xdbUfZSXClS3v3maMYRtEmDpiTs8pDSuSqZsWNKvsAx
XKmnlGHiuCDO7zCp0fyCht3Ad9kcAXaB1Jy/COSdzBftsdXl0z4qiB9fuGFFOqN0
UuZ3JivkHUzzfCj1EhKGmULuBsEWmhRMSoYuvj7D72U+4NXWNu9/q2+HQqAVqXUw
DwUP8atJV8rW84MVYzZ1vSKdDu9kPkVlMWovranMr563BrzOFOTIFEAMbAFRNcC6
B3OIibA6HrDej1sgMOrtqQVwb4eIE+TWzv9+w9QRLz8ugQDywrIMcoIMgs+xqubu
c8Cam2qh8SpZGb2WlKJ+sM++n/lyXsKJYZQto65I9a4KvPAurke1orLAEd+VmXVm
ibplw5/Gb0QL1Gonex4aTL/92drtnyIq8N6pntB4hnE8ItSvP5k/Asw3ObE1+Oqw
7rVe/vfn0BfUBJFzAoEjUgbON/NtD4RWJA5BhnPLsuokvZpTk/p9BblQw/+yXDrD
1yhR+hHzz7bSK9/zcm7Klqw0NKaUFvZSXobusRcn2UPaePa2AcrM/umpZ4pxHIhO
MO0QxemC5zT1rqtx/i8jfA02+sRtJYHskx7Un5wp32K8Y1qQ+6c+acmynPX9ry+G
YCGLGDkUsiZeMxv0nKSLPsPTQDEx/uTaxbH2ZxvfbmDp4Utc0Voa5G5k/jpn+5kv
wHu5D149vAbLDlcT+9SvwwCzpyGbvcdTJ5kdTHZQ6NiLIX2sYe+jiCn8b66k3DQy
0YNAhrsj11/I7NanV8FrIz33vE1Bf2I80/kwdgUvRCYxV2pxkUUnawcrM46mLHBK
nvo1tTnSTycfFZ4rFrFSPj2GSFJ5644nMrJ4Kj9to076fy1JGiJSEnUUTxsSxJ19
AGkWIyjM6oNHLvPmIbtuYNdbamMvHgl+dSOOISgHHZ28pH+7+iQj7Q2DwMNJG4At
0QD5ew7YGrKCo+bM3mhPg9DwG9YvWy1t3SwjiFw6VivXyEM0sXQLS+4N/zWeLJSB
DcixkNewuoZQTTHF0I3K7kF12bGQog8ricoN/duwdqqIatorIzJnlL7f52Hj7MIM
HWjXBuL9I79jXgp09eZIJ+7wn+oJfeWe1RmQkSqVSc41oEj9VcCN1xiHzwd77too
ocg8hPlUpBmXy0sKqpKqfFM/QsQzAtEWgfiL2jEfv0e/3Q63WrtqJFuKxpfdWYQ8
PPMfhtsQzOpKNYr7h6/b5GjQcCSO/TJVELFhypWPgY92eMqgJDi80G4blNxx+7Dg
xOO9rObiekIxltsfmzCzepssCPK1pEGbsZMb4i76J38bIzc0QxXSzdfsKdp5f6pj
sec+RVT5vBhZnYkwM45EquTWtwpsl+HBGmbOXW9d4i+C29q9aM/pRaF6O7efLarT
Yp/Np8WKIo5lT1T9ehidgLPGGuzzfe4NmQtVJV93tRsczsw3Hr/RJYo44rI4Om9d
YTiSj4yNqAJcvONAuO1sWGVeyiCQgvFg+/JF/WWl7fJpkm0acb3GuWjajKtzQ3BB
VLo46h7982rw2cDSZU92kSQwUs5wVPKnEq4E01zQ4nadYddxLpxZdFj5EXrRJ+By
G/XIrzk9yNKhSD1WIh0OXCWeEYqoKeGwtpI31kAKM+KQxed6q+w3aHvhHIuc9l+e
mhykSLoCocFG7yWMUmKF53AJDcs0zm8YTQlCiybeeO3vOra0qaPwR0rVGj56QZx3
jtWpTB1wVa9NNn0agAL9LDP7jBTH9nIlXTX7i/KjhKR8OOqpxcqbHMX0TrtDJO7i
ts7hmKhJoQ/52NptZT3jki+ZfUuy+PGICuoMNsEON9b/oLPB630Glbc0qGC5vNv4
0LAXLlk52TVSw1I2gN5NPM3Pn4rWYMaK47Om+pktv+VH+LxTFPThTyOB3bI+hWbu
CBxpHLgKqfJ4JgbZSPJ+t2pkFChl914utxit29FXMPh543QqF3gWcp25S5x9yH78
B8QuEld1oHvPMVt8SUh03LJYfvShuz3EFyzDCRwasVSfak/iq9JkkVu5vl3ZfGv+
aTAWOQQUNWVs3jfJvOb3dSkA9WMtsbG/7XKGcNZcS7nObG+WXM/Z+n/tdF9kphBU
oU9vJtw/k8LvikXTtxMc+7RhyMOUAsWBGd3+LLvzrglks/G45lDkE2o/MNtf5Alx
528EdrWk6xXo9XGZzCpIrq3k6m3ILTijxsPUygwJpRtRCPDDYm5Y+I9QkkCyaci3
6GsEKwldoAXMhrCvI8USwK7rzpim6Z9viPrFMs3iw3JtsrdPu29Scpjr188nJ7yj
9sIA0SGerjzTWNbNsc+T+s5lL6zPY5qrm0wNhw9FVL1xbkGGQLS5G+XudbywfCn5
VGQH7Y5nSaMcSKqYnvp8FJ+Kwz8y5YnF+MxD9oE0gwEnzqS/tAw42anCOVxq2ZiJ
eTrQkjetdO3eYCrmdk0Je40WmjFNQNNgNLKd9jFJCwJ8hJ7mo53HWUlaVUGETwt6
HT3XKVA/zmr1YYDAHKTAEtto5mdAahhT3pC3h2MsvPFdDP0C2GvtjWR3rpBDWtD6
YnGD2luH+stpT089jJpSKRgQv3ttqPJMOSNxwU5l1AA86LCBDiEyp6cEwvXX5rDl
CJqnLWmUl38KVDlKHFppmsOHIxTEnSzfdl+Sr9Yb34D23Rnh9GlMnNt9toXwa93O
+1WFDoC35rXKm/FgAhcpwddNMv+ETKPNM8JPglsAx6K4bEidt/xnzSJpkjOMS6PQ
UkgJCs3uh3QrkNoZeXZ2lwTskY8zU0Yh7NlpFwsjhfEVN64G3xLUEFxLB5xRUq2j
/Z/zzCibWk3LWz2I1Ul40upAZsuJovf5ahht+7gXYozaEkJ0OTrE0Fp0cbc/PWWY
EkgxosmhA5qPq3dsDytzNPw497OJi4m+vWUi4gAi8sG09wv4MMj2g7z7gyFfEgMf
zSzTdHy5s2fXsPFiLo/+hkZ3SMCPP2g+PyFGn03C9Icwy6HZ88TqqqwKK5Z8Df7P
Dv1OZAADxWOITnJtza+P+kq0v55rQuRb7SA05jO+wZsyDdZHA0PXt97fX5m7fUPY
Nb2bqBSItweLVFRxHpaLVNxf/iVEJiSrvdc6u/TQ0aqmmklH+vp0JYnZsPVzRlcZ
j34PuXwkOIZUs/rBNd6L/5Z9NiudQM2kbp2qmBG8470JdX5SionLPToeEZ1whYIS
/6C32c5/F/ToyqCgZ1edbqZqgKbkSVZIbXkRMwQyOUicDMPSPM7fCb1l2Tz92s1q
pZRet7ff2a239v6nMfU3rvNGLLNGS+sX+ZAggykVmiUEkPGWjWgRErCTr4SLKcXu
1DZjrx6nAR3t25QtphasuGTg9yBp+HvbsC+r6KEEe6rN/f8e6ZXkEnQ5YzaREdf8
sV/8nmOX4KJasxGm9OfI6kZgnNuZ0dLa95M1ge7NyFMTiPgCachdYwZjNzKTUDEf
UYLmNUELSRzABguWT3VRpYp7b97AzhOVQJDNgLgODEZqVj21Kos4UhfGYbso0ueX
XY4ByaTC0bV26ls41HCG4MAFtbEcSODCze8KTRFM6Ou4Aikz3+dLQ8Q+2SE4reb+
zRuubD/X5HdbZyUFHGdAsVC/12u+zRHr2LGAHzjM4Yhx8QmDVzRiwzR5szPZIoBh
g2IHDWZRKk7+OOKPFy78nZ+1O3QeTFtpLZMZMlVydlXy0mNWZXdII90Tn3FfeHtR
dUjMAQc6p1v3fSYlEvpHXsGTu52ZeWWSfEbHQYQksm6aCzILXmK2gE2DtItWHXDN
t9NbiqHhzwwWmffJngbw0eE0ciqxUnlCCjn+2lP70Ln7IeGFOB5Zl9AV5HjhcCHT
GsEZbacWt/+6JJTZDJLXVtDv96iBcCqEkTgSQev03reUnWvzvLxpp/3cqN6f+3pY
igWwPp0KWbxa2cX6xX7FN+SXMCKKSTgIa5u6irFmZaY/TWdpMIZWHV1jxDCGCtg6
8APkATRCfyQUl5ONHvRD3N4Yvjyd+T10/E6CqfGJKJVcWVRRAlbQP+G40csr6ji+
O5OSIxsktawv+LGJ/9dvIeBO4D57gRaBTBXIvNaEcszbtd3dFPLarcV8xTfFb24j
slilvXZrDxWFvWp0DYeJTtLknzeXQXAQzkG9REepkC1THE4n2ZPnR8tulL8t9L7v
OrlgUt880yeLHkNQY01aTtHAtPhW3fxQX7wrlIO+pE2sgTpn2iqc4ewAD+iAESuh
/I5o1XxuvIPbahOZPJ7DbvWn8oZA79oqg9rt+Wf4skCrcQxaR6YDb+QfSJb7m+Pa
YPDnXRK7vHc3mZsZ9eWgduPxBc7CuTac6rQxU0eooVxnRiB0gB9ZiCbb99GuojZC
pjNZEyk0CAcjqI7uZjDNF/aFlQsbjxRHFG0hqjJXPRcgB7mYU7oChcUGEIHUz6g7
R9R6qoyKv6aQ6vo/PK+g9LaABx2+3I6NuRLVLlww/cWRkvfLaWX++vWYjyjeTM/q
XgUgSKhVEF+XXwnN+zL4sB4KEeBlhzKvOIxiTFoWagRpOiejRbZJNN6eXdH+O/mg
9JcfjV++X1kaWdf65sQXJIlaRu2uYIFCstYTQC6d97orrsXMWXSzG8tKvj70yo9p
OJAiZPEEpZEauLPJQ+57Gs0xLfQqm2Qp585wzhDV7FYaJyEs10GQE/PbIAtfKOz1
h5k0iJ4cYWJ7WFVjXtHfasiVvFzxzqDMTBVx4933H47TK7zmpmSZJukvJdLypv2o
SGGcebDV6m6c7RlN3Z/cKYXYrX2JCClVgqjQOIoM1KaPznNwX9OCKwZr1Pc/8Eau
8IQ5hCtKu4qwTMeH+kBp6M5yAIcj3VSRfBw7/L6WnOPt11EAU4VM3xY7pEN0X93U
H2qkg1GhBMrADypjLiBkjAo9Woq2WTP0QMmkd0u8hafqPptbLUmR8cpUCd/f+pHY
Lpy7j75q3aM6cUVY8QuObvIiHopE+GEtjZTdpKz1QicBvJtnhdF46hCWZ4SJ3JjZ
8Hhq3+BKJAFNXHn8Gocb71k/rJR8X9wNEM7gfaDcPtKLS/MbabACec5yw7TZdIRs
qgeNltyti5KwhlGxO+e7up31cZcA+M7NHFM0wrNzYMWJGzHVBhLH+y/bXmKXhFTz
RUszDjPgSyyiv+fgO1micz+8gkAFhacy5m0i3Tuz4wdcb7PtbO+xLk56HWxBrWz1
s+9xXTET3Vc8LzuW31bJfV40xb0lGafowBI1xij6C8MQ8LYywIHFsykHT5MBwn+3
L6GlIWJv6Q7Ha6U7x+UbpaR7zwr8heVvFfauUv41bPhXtBk4D4NzDg06pXavkCur
uyBUHuw9UwumdKXlxYefYNnEspr2yYF8roXoOMeZqQ1MOPf9xFx3THxt7Xl9h2Tn
sGZCzOXhGkdycpTApjipqpIPijTz6GsMKklVekHNm1+/+a5EVhdkJRnHvXcduT6d
GmhExZzembt4K2vd5Eh2JEh4aSGpyjacy8NxBk46zGH/RDLZ1vzy9PXU2z1F6Hcq
NOub2Csm1ebRcwGIimO+OU7I6rMll0ZZg1ZmyPKYEajl3aN2flE4sAnhzYv6medP
QPY7f21wy0w6O44XrEjde6PaX1EKdSwW6rqY48ZR2gsv+BW+pkBZKMCFFLmzpRhx
Hb6H6cTG/xcYZThs9/85AzRSkd0luhammNE83Y14dTGx1btYVz9Xg1/juvW6Zrn8
JDDmdDY6qK/uBBjDOAjmgza82ILyBLHRxsvD1KmSnQFBGSZtbYc52dHwOYFCHuzz
4VDJR31aO8fuuOHMTUKQXjgeUeczin0Kt5T/qVODJOPXCjNymgXL/kmfcDE8x7H5
l/cDFpnoFjkX9eS0jGzt8As2nnIUIv+QId0URnxzo5fWDkwyFDTbdko9So7k5Fxb
YDe96cd1snpCD4DNzVahhT6LyvwE+Wdp3J3dqiikA/JwLtf5kWC8N7BLdsh8irKR
79aq+8aPVU/4jmCqI+8CQjf+1Be707PCPABGgGp5xiaFto9KJkmsURkTutxO58hi
PUcLwEQlPtmCXldZxez3s0avtiC5jbuzOjcX2j60SoxV6EOqzIprUmj8WHiG7ojb
EgAiVZHZjb9kGJe4hxwPiq54vaJrKq8hpTvXZvlJnNTflXM0LHA3IUw0nZnqQvoR
l1K4CTCk8agq4eZA1flP8DY9YkmlfiuSNOTER+mpO5zZ9HPaT80fNR3Tb5TWRHV3
8NaQNsP5eh0+BB4Q13hN8rqwTChCRbvGPD8yOldqIZ2z48xYUKeHNGcd4f9Q8GGF
FGC2AnuAQQ50qxPxX23Z7asVvOA3k5gEYCApGmqN+amcXgeSgkJZYRgWcOGW0/qF
BcRuTdG7gJqeL6y4deATtDilozPTB3tunjwh8ldMIsFHsC9PVl+vl1SsA1BSmbrw
bXhbAzEnMs39Az4wqzVYA+z4ntemKg4tpLo7m/4MykIGTj0SbHusDhrZjcG/Iy6y
+B6L2QCxWJ47S2fRZ1ZDyVLP2Ei1vUPNTSVjW0RyADgnk4V6Y9sgkaWx1n9Sus1O
dwM1XjtqxAUMX5pWGdvZ19dw8YlamIvM5Dnm1dL8SnDR2pkVwX9gdiEHMnJCki5H
A4tuVfakM4NGVnxH/Vw2zlmIDcQjG1Ilt5UFZIt5JgfES58RQJAhlFGr5ZTIh9P9
ajtN0jzow6VJRfLPkaHLA4ysjGOjiWbnCV+q0cCb3+WAhz3SsiBofyDS0mR+d5OG
T7go7tRMm/Z9cMZJ7xWUlsCHgzJvo+QQDb8d7GEKKvTWS0vyX468LlDxyKiFOfw+
Q8UgrVoWjImv0qhyRuI+/T0iwDHVrwUC+8+y/bEgdzjZk3mNEgUjEpPwJh+jqrTe
ggn2SrILDEZWuaQWxMyYo7fth3tCxWFsBbLAmsZkksm+cZSApl68DlUwWSXbcgwc
48KdYq3jGYSsVz5ymQlSRq+Vgc60RZ3HN47h9qoRjlmbzCGC6pTXtFuV/8kWddi2
jhRjR1R6ayapGshNZr/8C5l/LhyLtlcfqlFlW/wo/f2fI8DFtygPArgduyAiBgKt
iufHN3Ubr+ddev9R/ZzIRwJm6ucWFRONlowJrPYZlc9fupJS8OUlUeIX8VJ2KmKT
H0EGj6dZR5p6R17wazVLWugIWgdxz8v+6tHPeamOZyPxrUEKGzgei6ddMOSJoES2
H9B+08/udvzcN4jFLHozBy7X2iiGihhjGXidHOy57eNDQNh+kYKJfAqw/qQjwIZp
x4m/1mvWs88VjgB8o/zvWCE3cRHY+2sKDhWH6/CPnJze+0zHO+4LI/USxB77dca/
G8LsQaVP2Lg73PnqrspfLT1hoFMY9q+3Z2JiHbBDnDqqHqn8Fu52jP09IUH4bwUG
vh2bMMc7pKwi4QNhteaMRfOCiNHUtIUNOoDldAvAThGnI6NN87A8IrXJSc7N1biW
8Qb9hBfPoOxwqrTNI18hHZWSS9cuZYlCBRhKFKNXwTvcJPqrOKXZM04cLPIyhcR7
42KsOgJ7VqJzOYkbqKt/Ps4oNEQuT4CrHZYK42JaN+nqbeUH/fH73I/AcvO7/p3/
3IDziCqUQK9lA0LyuBzNkC0YFtelTBx/YcwNXrQBqJ9hxN9R0Q5KMb5yKsaQ4jIo
srAPGtIonn/s10Y0kYe+aK5A4UorUFdJv5Jvf0TCWsk2+6ZqOu8EcnPHHL3wXZkn
31YcqnAsTR0HLziYBV8u4x4xgmfAmSBHuH7QyPPwYS99nytuJQ/kf9j1CCQoQF5E
NNpy0jE4Oy2ifiCOsj1BKrMJZt/FhUeZn54EqRQk5nne3CJOBUSaZKQQgNcCdwre
HMdkEhSaTwyHtATchFW2EzFQWjuX4w39jR2DQ5hpSMUgBCRJ1KlC0+/HVPIDr5xn
2XAqIm8QUYnysTktBxs2ki6h5EfxnpCMfvfpBGOgcWZjSQCgHRVV8LLR9t2NWVUv
7IcEgAlpIjJ5gT2vlkaANzmySc505mmBrXv2MZMopAy9kVBHPuPJ/AGaX4jHoz6r
NfwuddgrDM6BLp4L8/GmCBro5lSOlnPMUOeq34VQ0PDaVnE4w9j6Q8N9Fuoisamv
qUngFZiz1PCqt0yd249xtfrWyFPKVnfiuvNKCWOZhyjVU5R/yzumGfLgiUujtKLk
qKV7wx1nfeWpy8Xxr3nc0U3Y4p6770AayL51od0JDPTPDWzNZHxJcye7J5loUSWs
ep8kLHYYYJCASC1BBAok5rD+Cmx4S8m69FJtBbE0jVr+sLkZcJdfYoKt/LVYkmaD
dkDSpXGP/VLHlTPFZX89apU/CvQbnPhuQfylFHGK7eNJHJX3b8DfiIB7yUA2fsmA
CPSTA63zYQvdHyJitPdIGOGm/dt0EiAugvI0JJ9v6BebtSJOcR+AT94cYqk1VxaK
4AehJEIrOyjqDAQkbWUqcT4pg50mIcmGrMkM4eogLp/UO57L8KkjsOk2HPCti17B
RXmT4/Z+TWRK1izHpzuPEsac2mCucVgeeQdKtTcreJIFAOIvH3SH5OSXO4kpB6uE
New29s0JjuEAXkazwjbnkWA/y73Q6bh/ZTy3KrYX4ET79RxFcFtLlFUbjPgT1LZg
He+Ty74klJQh3EviskPOANJg4JOMR4FvyXCi7RyX6gVqQ2lgGuTXCaZx+Jp0RT5E
VvIvLPKUNkO+WZneG09y8C4y41P+MrbLjt7r7IkgCxTVTHbNA1ni03iKMv7932EA
8yCTdocXD3dNrbjxAOM/SCeZwAlwDa0b0dlLAvhqweSfKIDf8BDaixaFzS/k7SXx
ABLrL8B/lkiQzquoJN1/Bd/zIEGuL+cYYnjEpwb/v+DYhaJh3mCi/HZwxNh9hbnM
qIlVJMhx29/6kDvADZJBwwQdbO2cTDCU+8pKzBZtNrXQtu/Y3yi2GAmm7HBJMcYW
W1peVvvu1XR9Ee2GLs4wO/8rs5p8/MAUkbVkj2vl2EqFktHzVNvfocaI1G+4kYAy
HoJblfTbIJyz6jz4jtLxMOrLnoCw+AHPGxfUfFvT6ax1Hcinza86jN9n/d/1925r
Qt7HWOa1Tyi42PkwgwytYwV+/+IkqwDcaY3DvwEEHUvIDpyl+OYUNA6OupHJccwI
YfQd3WZKP5fkLnqyelw4eBqAk76UWWjBKQJjIB5qX9wt6cjqf1eEBtT1F6IL4K0p
M/JM6QYK5nmZO498rIQOgR/H2/jKILJG7A3a99CMbQpNTyOEJS1BgOpOxj9uJJHx
t9s5GhlDsLs2CU2kYF1PAwBkOCtopTjxz7Zm9bTXuBZ+h8/K/V1jhPn5EYImTPiK
674FrS6Y+l3RzKr9YtHnQ7Tx/GnjwS1+Yf4sIwpOnQkpivblLA/DXJc6Uz9HnscK
o9sa9+69HhSdW54WB4cpFXneeS+S1S0uozfv+YSbSg7wULL2icCm74JQewIDvuOB
ej1NZ7bN4MFv+Y2hPihZcBEDFMXpOGdV+5DcINmVzTTbfDnMPqa2/P0cNa/aKli3
Y/4oRcbsiNlWPr/362hfuKij/6s+8QqsWiMUkztqoZYUR2pGVDNt594igIYzg+B+
8wnSdyDmuPlucRDF/Giwz9cK+QLuIEG4x/9qorwVxc0jmmZd3KH9Rh65vcnXaqUz
+kWtKiS/bHOjHEu0PPDoM0bb9p+XHahD/d0Fh8kgTmfTcWdnPxybrYi1XdV+/Yv4
0K8MLqbUs8kZPzyOWrbom4Tigj+dxtaQvNvus8tVttpL/B+ldDJvXDx6CTpTJCcQ
ZHfnPdMTOdKI7MY9wlK9nX4kEOkrV+MbTjK0Rwop1+IU4SE1+nwtMEeB6OA2ckNJ
wQ45M5dHdlY0hpuSkqABws3irFnCOVUqV2FtwQlqyfL1eo9dKxUim0mMB1NCspKI
XTSvOtpwP8BYffJZAVdEE5bRyZrbDdOeB9GRGW5YR6XndNNlkTOD/EG1FtObnwXe
Hd0HAjQh0IYbVmqr9Uy2fou6dL403PkbxhUQgDx+TpW3VKHXDTh2qlRBMV/Pd4IN
hrJSFuxfLV9XVZAGcPsBtjnokrkV2JTmD9CVUs4QkB1eHuHuVQv0afeU78Zg+49c
ZtOX8g+2tA4NomBKI6v02/GiuVvXncdeqSrdAcPfmFl68cyZUGs/pXC47ltWQhJz
SZDfDvJA8+dI6aHoXgAnW4a05YrJxAPlsgf8bcnWziefolDZyqP0Osr9OBBX9iJe
/jcQoFME2LwNqvaRQXHf1jUBtBCWh29kkJ3lt7kDQDmLx1/I+o5L3mLPCzvnRxna
tn2six459ajOt3XBYKcK+d+XXpgWh5wWtspEKtC+El777KV6L/Vzesf6wNnQ+cN+
ZaRxM3nodQSAyhtbQUd7IwESpJ5LRKINN5QH1trNSQutOGxhH1VVpt5fez+DAgL6
no1CuCHiDcxIFQS3LZxB4prDzG5iuOUhzkujSepzj87FKObCjy4pZqxE5V/fqlQm
EU5Lar6YyMMhALzkzrlEbNl896Bzsyhejo+h6AAwP2P4o6ly888nM/pZQs/hP1Qw
iBBnrEWqF5CguUnv6qj36FF7cFCEEGAYnG7fYrZ0hZFC0AqsFjhdhxN8HShG4Xq5
WqypHolU6WQvYmCAMpYpAZv5fmiwSLT4mmojCHLorr3DBCgg3TcE5KpvbynnVYss
kbk7oGw22mUQQFyOgzCEOEgahf4kb76cbOJiu7USHC11HoKduc+VT0Ces0jThUDZ
wIBpP6LuHuLvgv2lpswRvunypNvGe1TwN3cTvgSN6wZam4GzHlcODke4aMpf6u3k
+KTma0eNqh5yyaXJpqeBTRnufiFT5CwT6Dk5veQ2ZZBrcIBjhSTxawz48lD/47/j
beBCc+Vq0B52+r21vovcCt544qYqMNgEqIs98YI7nHb1UXsNgrhBwqA3BZ3NvQN6
P3pHtRrFZOtkxTFQ3zwswmXscT3pyz7caKQATjFOfb4ab0+rQ/dzo7qnkuEExnGR
rwXAw3s95oo8b+bSL2G7gHW8lhfFCW8VT84wKRGJNfAH+SujBXcxmDVXjCId3AgX
+cPssK4/nJvIElNJ7Clae2bNqmlL9AtVs9z0kFf36Z+0vpcpVo/E4mckWtsl56Bc
oyV1JJmPiOGKS2jpUzTHipLNrtm+6/JmI6mG8WMrxf2CQHXlK6dsqlPnWEgglk+c
ZWo3sJzO9uH4SLChBOIG0HKb47hN5j22ZfQmUD1iz1q84WhtL/BRHFRrQH9UENjP
NDC+2jPNlnPb+vxQYkC6jjItoBt23vD/nrhBAY9HDiwDE9gxcFeabU214EKcmbKl
C+7n03c8kw3fnKNZhJ2Y8R5vgrSguS4j3fCoeaF3uWM5FMXw0I1+0yvd40TBMcec
Xw+ndPrf/gBzczSU5GxLp+g7wkpc77cNXcByUjXdcLMQ8JpEr7W82HyWnNPw3ecH
Px0enLJ+F2Q43ZzUjH/J55lvnkLVB+wq5cvkFEZDHzAPeaMl+cJ38pMKijIZypE8
jsiHPUQnakSUofC6tiGnhORZGEUlbiowpFyEsxlud5qOybpxpBZjjHPTP/poFyTc
7vSq1JG1M8C3yKjyC2QrrGcYmGH5Exe+lZu1w2qweZga+BgDhGcf0Mduf5pbszOO
u1Py2Ghc9QV6F6CxLdYRFRy39DSeRaKAnM91ZZAV+GHc2P83sAwEb5Nq3sb58uwe
qAIhmjPb45k2LXNhVQYSh/rC8RZKYYI1sHRv4J0k5nFjKP3tdWJ0Zj1PW0IX0dVn
hUy0CmrPsU9TtK4VeIxnOUpUVZoRskRSfxVQdlvbz86SlhBCBKC3Gmurxm4Gphz7
uipZDS36F1zx2aqr3BXVDNaQFho3pnWVcbP93zJQDtE2zGPjnoX+GV9kAh0BuDJM
NoxExr7cFRQvgH9Befsw+Q55HYDvR9uxdiCyXWOFtr19JJOHVlqMTONoQ9A/f5KY
AXrWkZkDSV07QRjvrmAb9FkAIPlRUs7FD5kwpsg0pMaWBjGfGrIgD2YeiXVf9OLa
C9KxknD6rh+M9ca9PgdslPyRw9MTGZsR60go5/TNiooFKg1Pu3Kv0ywaqzqreWCf
Ai4H8ZzZVuVU3eQzIQt1pfjHkYS8oXfpB9/sWW4+IxFNQWQIZQ5CvXRmfHuDA7XX
qux+s7Gdi8QQ+RSTWj+q/MNb+AzpQkDpIU1wjqK6WsXzobC0YOyoc7S0gWOQs8Qf
AHZdZVZg72gka96NF/+MrneMYi7tajH6UWI3VpLqGJnx8mgfVyIXAl0R7eskLjNv
nIi5SeSmMZvlz0S1UkRkkX7SMsx4oChQXeDG9DnBgahENwLMijsSFSBF8oHMfB+6
lZHHWZAHt05GQa6P0hjrO01eflQbiasw3tHHFhv1rJVhB3tjLjErH2aNbSTbhrrA
SWVu/fRLE1lDn8G2tEEGI/D7wtZdt+eCyLHSymP/JGju17guPj2+JPWiqsN4Rc7g
3AVaV5Bm9fJKhMvchoEBiQu4OVkJ1lgj3xVAEU0La4/mQcBIAzRuUWIE+z3i6aLU
q3uP3IAR10O+THbi+elvZYIhHx7uR6AEuLG1miSGVdrkab1UHjrQAcw5R2mS2nNu
Qx0t+AcWbUO+b1nT8+LKUYnYreJDjcIYV9qfxDjvjRu14zTDRwOgiCStsTPHn1Tx
tuw2YGyt1YvCSemlQuuDVLrkc0iQDdTy1mcOLjWjC4UCs0rZEHo7QhgXyzuAhv8I
8IT/vyS0X1JHHgSNNgmm33va/wzK6Ueq/OXPR+LP9naMUfl8kw5ScYYC6+hHzmCL
nc1X2ohK4tyyC7Zg1HsB2nNn65MPa8l5Vzwg+mV8/uoeW75arVWPJdfsrDZsD5KB
Sq7DL7+SU/EccFnkOiaNp6w3NJasRyZu/tM8GMFrwv95jVTmIgt1DjJBOSOIivzh
wFjmyBWRGKdx3+fYWfrAbA+aGptXXwBaIaQbqq3+ASghXHhrWj9YPSuueec7p+/W
dgCML7sA5GWOw7wRfL/t5RcFi326mO2PCA7nGCYY6LZT3e8eS4B0pLozAWUVzNji
seQlGo6Vb/91kiye2vCzPFRgwiixHWVpvAKgnRlUbPqYaXWC2cY8v3rDvgzOReo7
qDJNosmE2CFxQBqw+beB45uXzUiF3gMlNxf1ViqRkYf+ss/7Lu3aTUrTjdMVXr06
ttCHY+tTxqqECseG2ErwIze4d7/q1F5kusvKWOsFmv5spvMLEb4V2gtnlrhQVLXY
B5Lid2WMki7xpWPGXv5VnE6TJ7+w0EaWhMRrlp995RNYMbzualxncqH0w//d/eLa
yhN52trgrBXkrWE8zz3sKVP6v7ckNQb1Uj7r02EIHqh+FU/GZADRrm7yAgLFgTul
3F09a+aRR4HspgjCE/+bU9NZuPqXdLDQhlhzJSgohJ0rRkhSEbAwnYld6M+glwHj
9qolCcCbz+J6Z55UGuFfGbiP5ro17TuwCVNsxZTmwDj+kLWVt20oZS8yvM51mJPe
bWYv1gZiL4CLu7W6f+sHzOBJM3jd+S0Ncd26ieITgR/cj2MtqpIctPSkuDRFwQks
1wxvwDvbgmYQWVfvY5SKcRJd03eKpu/IGFPb5DhgVtmRTOTQTez56GYFHNMcIl0H
wHWf/3CAMKofJV/RMpl6XkIJrdsdXBSZVTw2tDazPzH+gl4SCwA9cTjpLlkVtR94
NQg+3gk+cBNgYCP5nRD1TppPQ9s4ivw1o9T5bheZDZZPMSaGqkzzRYLyIFoX6MPo
ryxythEXqJZriFl8NCGoHHAowixkKCInvDReaTs/1/a70KJ8tnVjTNtIWVpv6B5y
b7apix+2lJe1x+gYFlwnhcl4QwyK+ZrKl/EzCxKQyD9fT8qhfL4YbrXet6KK9eVQ
uX5zJMPNveFfVfKxZv4/FnmHmydKWOOzjOBpVbezwWI7+2L9LL7AraTUKfl5+tqm
1bWb8D6bvXMkzCt19sHl4lECgvZvvN36s9HA9j4ffpS5jwOBIp+T1YaDAgYM9BMM
KaVQadbWPWXAATLC4KY7GX8acvbIA8OAkoFtZxVriiM7DA2xOqp6XEFoOvHUsloG
6qzcZ2VmX+Q7gr1neGK7LyMnaXRw0x7mjULiNkds2ReQOG5wNjlJudXlmcK4iDvI
jiUcIAHdFyOHBv6wRxMGRQUlg6Yi289nppQ1dCcNtUgGtPcIS+Ul3QPdFxqi9W4O
lRVGv7UuojDi+UB+tsw5hdOgwRx8ANcsIinY6BORWLPXGI2U67PJBbLOFkOYySr1
bY8H7/i8hxgifWMJXXH3Px0pNaHgQKREe2JS75J6MCqnebyAJDaL8aVshRcgCIBc
FBRpVx7W9KCzJFdIHbHA317hlib4WNxnPZbVP22wQ3QEoO8ZERygvcPzuSLzdYXP
PKhePHksvIEN5PJMjOxeKD5tlM4rQ15ZtabIuABcQDh8TYf43wwwACFTQKbF3odC
SR7FVsibC1cvXcZdEafUJlR8+igJG6MThpUJUuhaZ6o5ApHWnR8PeJQfU2qM4Iax
c0GqZ+yv2QcskJjxCU5RL/UEspdGGrT4pDMYEk5BNaQNYp+pEhCObiuQwevrhGlr
y9cDYWhtIl5vl7RSjYGTQqPrE6zs82QECBc/PuP0dAEGnbp240jzs5DUEXQJ7fQr
MXc06nGBoI0Vq4v/veX/mjvtG3oT9Peu8ZHkelBZTdAFvttpmCeoeBss+ZOCxOc3
WVH7UVQyJE/5ia3iR+5kg7f9A+pmYJhNXVBC61Dr1xmyKDMjjXazwC/bKQcFq7/n
GoYnw8C4dEEjcCpjzAqw7t3S3p0FksFCBahXYnWzHh9UbfYPCsblHIKS6Xx/RQQb
wvb7/ssl8DxlxUKseKccDzIMQwlnz9L+7M8NkihZx/zUYiXv4HTre3xwJUBQzmaA
2Lt7dsJP3B6NitsPNrSTvDlsh7CmCDM+Ml7xwuE/jrk5cvMrz1fLm/ie0QK4nMhC
OXYAgOo76UBcvZvZzsszrBNK8or+oEHyljijipcg+Oai5pSI5NkjAYUjjC+p38bu
dtKZVyP0W7VgrOyrPYRjJPapexqdDdL98mAquE6bdhxcNgapD7kzCemCSc8+5pQM
BRsgdd6mITScc73OK1JlIqnt+MPx65bImJEfmVv+ZRP/ofJN+6H+UGOztmRDl2gj
UBOmaG/6GV8UKFZGUKu4GD9Z9KWR/CDZ1NexD70eULlBEckTupjjyPxpgtGz/zJl
QO9yCi6Bbg9JslY/AjK3WT4GtHZYUuYXH60ZxYe8dLlTGqFoKsbu0j2FpGGEVYL/
g7PzNg2k1XG8vc60xt7aRHEAFrKf2zQHiCUzfpfoSHYAGG74LExCOzwbJSHBXW7l
dc2G3awoIRsY23nY3PTfvzkQKF+e5jvs+JDoyk95TrMR8vsvKElrVY2JOVx6feV5
QVftE3AMCaLsB8kDVH/xbzTGYWnspzyiZuNJfM81Y7hFXj+pF0ulwQ6xuV2/xeaS
n1Y1IJqQw5s2vvAx4Vjh8OkJyUpN7++I87rUTi+Cnn/gP2lr0UocMCzYOHMV5s/p
IhL8N18t9b4Is0BoG9GQE/IZ3iSI0QDDpNtcq1A5shQFqvlMXWMXOPsGqTunPRmm
gn/N1bHGY91DRpzwIPXj3TtrcU6xR/1Bn2BUTBOd/WK2ADLkcAUTKZKDKH5Pcil+
5871I0uaQPmt2IcAVn7YKWEL52zUuh88zfQgmay7J/e5VO9X2jXhI6laIazHqjhz
lVxyO5oY2N5N+G+pbA1R3XsLsYpfX+No2Vxcoat0JbuQS2fWUbbB8nNFr7qx2Ro5
Cq89o62Yk2dMzo/hI5RE9xdxdcXb6CJ/kd+QrrJPWHIeOtRrcE1X9bUgih/q4Tws
4MBpixr+ogl70yH25359MLS9cLrP+QxnNuh9FMDQtcaFZcmGPKhYSu5CbV8D0Qb5
UVtkrh3duzuIiMKtvg1GmyEfRmfabFreVbvia0SkPaJv7UPQDYIiy+orIygy1iSY
D0RmM83IWpEcw3rcqhqz1qrQUSgb3yJSwQTVqeeR+U0FcKYj9x2mZlrq9IFHW9c3
4sTIPROveihcjTzH2pxrgoGJmiFc5ZLBF5gqJ2XuUg7XYkcdGtAn+6mO/bJMJkIu
L1myylEMOai1oDYnRC1LkY99UoPqHIVzdGfAjaWA2esB1sapH8rbgJ2EuUWuhovj
W9XaBQN6lt6VeRDfsaSuQVonUAxi8YEnB9efOAxKCjsfQJkioUihRPnItlnFESYY
KxtIEjVIT/TZd7PaQy+Az8BsIFKENLkLvC6rHn9XiG7W7t2QSgC3M8KboSxGkWwg
OtDUKRJoFgsdxgaIbT/JptG1JgLMYwaLRPS/ydcVReQNeAN9NBFZSTbjdE4eKsgD
kBl2cfw2e5oMxxYuOE5wj90StAsf8IijCviP1kR40gaFo5kULTBZXL0dtFRptRY/
7sxQJstm9dYqRRFgCzxmVp78AJLUwcw93xdLMVf/4P/yN6YAaKl/nML08j5MyKu3
P2r7WEce4lsJKZdMKf1Hkg2jdWJfOvIXbR/2xffs8lXw/ZJoU26JORZ3FLkQq//o
P8wfE01wuOX9LDkPQH2cFd+RepIdUw1fu80Rn9+3ADoO26Id5+WJtkZ4AL99OJWK
PTMkR4GOGkq6igaf1fYa4li99uptid1uBZHDt70acLOZGXttN052b/L/jssweO4x
ZDAIhajUHuUcNSIQ69eLoDpE6MbWDrqGRxYlbQjZMU+E07nnUcKSmwE+v5VBZRcN
rFelIPq/QyIa61L+5lNK21cMDn+uoyXCnTBKvRoV36ysXhOuHc6TYI9L6Bt72wwO
xZKQNgmna66wbY0OB8Xc2ryaYJDsRqpw/mfoYCmEbWzNKvU31O+x9K40tWVq4G0q
cHTroDkHp82TlGEDW5wOd7DpfTxm9MuYDbynAKogNhTmPh8RiUJaRRggrpLzCblw
lX3AhkW8nC5F8k4v7rtN2wSupqTKdfwzax72k2agmtFk5KsmvKohGmWm9R74V53B
hBvxfmU6E7WFE4VczZAiwh/IQQ1P3m5OV79u2zu5kklaxODHnJanF6d3HELNUcGJ
VIN5+tO6zda51mnf7+MWnOXJmN0FEwEwBdp+DU+PuQUC2D48HQQV86R4gNnqNyRR
Eu0LJkv9PBlHyiY60RpDtEvWc4lN/ndr+w58sNRske31gfuYAo5GVSGZ2hwHmpi3
TPj02X25FiYTL+kRMVWEdyUCp5QcUao3kRhTjJPjf41ScR6HOIM8WYYYzkPjqo8F
/34khquGTAiFTLkvR6ldGjIYpN5a9FRGxeIxumgjY9/mPyWpqrJVVzNci18Nt5j/
9w6sVXBliKyP2jWg5udITf7YkymnYePUWsoJh3HCrhxHfaffpp5gVs5yRRe94m1U
VNu9QY5WlhpflBYvm8A9RjkwKvTf44ZB93Ov1YBA/o3cpfD9jI433NkZV5YuDLut
gJfiqVhMFLbOJTt/nMsDto3f/JdP8CH8CPGzMy7MXaI6zX5JbUh7RAl1fzEOLwQH
4Qy4LlFZHQWN267PbnHOhCOYYzpti44GHS4TW147RVu1UCZUWkcCG5+Xbm5F1uDn
rZWnO/jDp9ldFJudHrkKnAg1T50D4fjYoRTtJEghe41ShdoSekhyyPEsA+OI3BGX
+UgGNlWrdmGeolPoy2NMLNriHJccWhvvyuTiq2sxB057HUWG3v30bwwl9vd99w64
IZ+sEtCPH6g1imKOuyaqBVUdOgG4VxEn+8xS7j8cSnI3XezLJRG9nsSq+Vml+oux
hXbt0OgyTQrsVtaOjMfiayDhmO6YUeAIXnQS0dXB+KK5JQBYfUAZJm3tnEzfCVVo
NfMQVhcAjjHWKbwHpIucf7za70l6PIGqPjEdXuImNuBp26jUCDVs213zhweuNW4a
fjZtXE3GZcYNLS+AxNnFixO82rDJOQt3azgfHEPXK5oqwAv2WU4V0Smv5hUsM00Y
8uIzMKHr0xL+3q87Kh2NmHBAm7U7VdVNcY0h87uK3nZmv3l6NN1bILgta6uqZ5G4
J4BVlCF1Ho+vYwKQNfmKYFbdsj1SF3q8E1ufoVuj9sPO48guwiSIxL4j0m/yjhwN
ochdb8hJl4Ue63vWnq4qrjlLWjHMwr08fnI+0llxKPQvDXFY1Jr3mUpTKsCFYx2Y
/oytaADpoO4+rinpZnccKOk6NeJL5XWxNL4r2rD41zEEKZD3bdRvrxi1nWS3y54r
hRbujglJBtuYaI8L0yQHc455PwowLFVEuRaBU1vlpIxJDh4AFEYavfFephp1pCrn
xOyQcdUPJdaWVpVcLUGWf1IpM8ZE8FPDj+gXaAeWKX0g9Jc4vmRu15QkJH29QfvW
cIy5X43r0E1TmNLOIv2V5JwWPAnW1FLzmaaEPD8kCyUC+TkO1oxVpYJ40XzZ71ye
neN/ExLKNGsRQFVZXwgekNQmaUpvOKbcKqzUqYg28ys2Cv/M9RuqzkleEjl0DmFa
CeaBxldeDVio+Wyv6GStri0vcpKdW+wRl7pJYXc+xcHUxyd6N5dVqL+MJJ5dRn4M
O+CKLMiCaYyaLLjqw0K/1Zs6AA1Ifd0Ow8wDwgdsR/vm1+Pt3lZXhks2wrW4Ce7V
wwzOplF4tlEhof1S1qZXz1IjcotKA/ujZbNRoEMvixlHfaJrR1CT/lLuHXe4qGra
J1eJhZMhLZcxwFKOZWpVb6stqqFOk5Mk08oEjjcm/xQuqjaf9QiE+OxlPUVw1/Ku
SwaKMs2QXSIja2nhWJJiNoOgBYGyTglWCEIR24C0zZ2yHIIfBrzpGQB3B8J9faUZ
RIThNBtS8lSH3oUPPYfxfRi8N9iliCqVgPUNHe+CSvSZuFtJZog+PvAY2XC8MQrE
8fpykb+Ct0XTQbIp/fiuDHkOBYs1EahguChn0jw74P0yWXoaUx7WdHXq0nAL59Ef
azjQd+3u67ZEeNKR+DmuOnSwMWCc3Tc8r0zL6OX6MrHMH/LRbc/B6yJzBM6dhwqG
EQqXz7F1bTXDauoDwnBz1o5JrHV2mexpJjAWuXneDweLlAS0Y0Q5f7v2qAE06mlW
ZQS4V7F1019P00KATe+OfRSlJC69tK5co7EDreg5aLarZHHtqxOJFKACF4pJenQl
PIkKA8/XARhgz8ofoyawIdct8pRE176qXjqTYD3m4XahdevK3e2+G8HI86Z9lzno
p2gFuw10XiAUg9+3mEj1KHSE1gV1FOoKrope3PknK+XGZp/Bx1A6VIAF+IPUBhfn
lHH+cLhxQBsTNuxDtbki7YhsV+mXlalr0PM0Tovv6qX1JjK5fntUKosxAsDjxOvo
W7Ti2bKwPgOgt5Dl4SUpVIv9qhzdr4e3rYbLzej23Rep47/TrdM3xdkxo17/q3k2
aqNWZHIpH9y5PaA+vZvL1C3PCQIcZPjOcmydK9BSjScwmM3LD9yFIYu0tBgbyGp6
Xeth/2lvvAYnyRj0lD478Q2mjFZ90GzvGNkNxIWEC8s4LN5CLTOCOv+PzWpoowzz
XXizTzDZ9Wa41E6v9IaGOpYpusCCReVXUu5x2aGQYhvNnOQ7ZAfjPQSFdKd2HfBV
9qNC3zuixNbUaRI+aFfQoF94bOViqlhaK+DUMpCJm6tyPoIDpzqbDpk8agU5u9cz
uvUkjOwNCYPyApN+ytfKLDBMsFIOu8zAmaTHjXicyQuRaS01OiRGQ6MppxASu1rc
qbMaC5LdVl0hWi8GgMTj1s+bkjgEcYL8VmVtwOK1OynwSClWZLRl12SuE7/r55L5
MOkJUxlIC4qTHMyyt7wdZZ0obg3Q4crHB0aNK3uCDoZF5kF6hIqHNysSurlbilk/
y0Kr5epmH5RWEEcg5I+47ceqq8+pnN4BSZh+XgbtV2wbIfF8FGrfUEaoOzytijxz
xC9ULldWhU2J+B8EzibiaeiYY6ro71DGJoCkW4Mp2OeoTY2nNG2Q3nBGtjiumlUg
fbvZ7y6TFAHhCTkqcYTLQ43C/hR2xLXFtfEFDPC14s/rpGQJl38UOCeyVxMd0d1r
4pJIfqzlVJBNdNEmEyhmDtlrYf7JYDGop5O9v5P+7phO8aJLLvmpEz0G+S3+LsaU
BGKpab2gbxK7fYr969DOgz3szpN3xkjYW2eZyvN5wxoFhNqLPiH9/u/z9YDf71mx
0ArI2q6Px+1n9be2XseOoZLITGOvZsn5IRc2LAgd+a2i6KNyjYnpzjRJm9+u/S9M
CnHv70w94BPkvGaUeQjWvaIaqZ2h+xN3zdiX3l+TueJQgVydqqjoNEqA7GAiEJeq
Db4m6kZkyGlzVys4Fsa6FuwnuXiN+7LV+EsA6O90S5k4L/cpwsIdCChFv8ooowmY
9jFzVGLltPCBTVQO40cBiOmEssZvKD+Iz9i9nNPfA7lDMBKHQe5GweFiVoQFwpnS
9vOxuiJd6QV/MOfpwQKbmMv8+pTRNuzVOv8Ng5QNyGzpbJGuv2jjKjEtfatNq0Mo
RmV0pEWeiSvhj4FAqtQUd7Y2lBgdSHISpAef+BDE3/cDA9x+08b8vlneWClr4R2H
LaIAHDPXTM3MYX5iBNv7pyfCNxNmnxRNYYG9zmbX074kyRui83KT8Xv+ncv8WxW7
YnYqLKDk23XDSNBgrAerHupQiB4POK5ovL1YTOWAG0TrzW/YAxDPxuNzIq2ui3Yd
EqzBTzZG0/AijsqORJLVAGwSK0h5pEnS2g4VcbbeKknsddg69OhEECIkd5/KYgL5
yL6nYlQhxezEHaadJd+CIQckkXvte6Mec4lGf2h0e9pbanuP5qlBPfH0x2a9xkWa
SvjuV3fAT4mvsXVsiERqseKEZRgJ6+BhixWDRp7vVBeXKZVhkHRGE6zGue/hAHu/
ukDKinAajGtQ2R1If/JzowpOvbvPzm6mcl4xLVmm5DhLZWgYLIL5EqRe++Ode4FH
Jnn4uBnI8FPd/BNY97r+mJxOiyQl3Vc9j+/MNGKrfzwoND+SihNXQGec4uxUNNnR
XJGThNWzuCbv6VDfdHFOR/qcKR0qJWnNYNzi/hERkc0qOQWt50nq+zDwPquoaPGR
qaloFDmeSE8tTBeqimQugZeyoxC335dETf/+2GyG1KFhLQCygMGEG9mESBCBDhH0
dAFgv9VQ+RsTmma7AN/d5pNtXNQaiviWSkJzKpqYI1IEUEMNOHoYPE9MFnwdLwvy
pTtsasKPdLzbb66zZkzIKfjRbr/xiI2/tEG1HWbSntBFmWOAT6DrklWarguHwHqN
uS7w8IQH8MRmtHll6oNDXYCyj2GFQ9jBPS7xU6GWjACbn1Zk7DliezQMuB/qKlB5
s0FljF61TgeJXzIc05IgP9huDLYDtC2atCqwRVtO7DdSMA+ymuUyL7fUvpXqV5cH
l/ny12z+CrNn7qLA3p3YDfDfSrW27qYkY2yz8P5iVZthJljlDrG024G+zggYERLe
3Ue5dvJ3+vAew7dDcdnjQTaocKATO6nU/11Td/xemegZFd1VBdW1iO54od0Gu9g1
Q4KQteM+54eryoWZTge+zj0dvH8Lmbbfuhe2VYxdQt6bbvFsd0zhFu8GXomS1law
LKKTk+PTkJDXSOIgAhLQ/ecadAE0oj7E+8lH08Aj6YTAEGYKUqepK4ElMjF9GZ9i
4w0M+ffg3FMnY9XdhpoRA+VRKYjU73UMOm1TTqHKsL32X551HAfoO2iZI4+CYa/7
yZwH6P+c+QLyB59cYpb+/99MplPHlN1Uiq0lkp5WpBrBtyll//aWak3tP/+fju5v
bDg59vmwkodZ5ZHuLA4s9sUKZzvTAWjq2g0zHv9PbDbsnlUSMWKn/nA7G7QpZy7Z
wywdmsS6bgI50o304oD5tS4IwjIfEAG30rmcBYg1km/fR6NPhLwUm4sYw+R/zffC
odPBkf9SlK1ZWuQjxLCNg7X6QNx2kmtWl0EFr3pOvGSY/83kgCzuaw4/l564ied0
tg4GAdXJujB9e4kNJKr/USv3qLuenez6UEzp+s9nStruHbennHGTwY/z2Zo+tCdO
kCvXetWWwV79iOlBgljh4zRWLgzYqT8Tl8hAUSHHzrB5wIay+3oMJTsLwFn14ill
AuUGXDl9mh2G99cAY+GtivE4kVtqlTnHvxrTpQYPzXVQZG+C8D4TiAonYapLh8SD
gTJfjdN+2myjD116N480uo+mO7H69S5VFqkwRbVl4o5Y7YwETWRwDX2dKj/lxyCv
WzmkGQ2Zhceop09TLibV+j5uUdhKflLwst2OI6qX7qEV0kqlkOXt90xlxwgP27XI
b9ujAEG9g5M8hD9LZ2FSsDLVaXZEOLdq2cmM3NiPPrtqojPcbeGzTHI1oK9DrHkI
UyybibADmpX2V8TVfzLcNf1913RQLHcgrEAAVGn0ni24whJ5n+subjJwItEUzDKZ
GDbTu87zvaBWb2H/PuL/tE/CiH0c/6vOxBLsAOzUX9FOni7yfEJFnW+svGUUe3tD
vyPd2EB9A66l0wo4WEcAbri/5TwL5d2I0R3+TEq5DFxzZlSSlVW1ZEKqHIdYAQz/
NFCgaMP0ItPtyOHaeBU5P6Jo23CLxpmSK+vy6NC+KWrwlDc1ovccyhILeseHttAM
sow/qMqzaQaE1d3KoYbMwBS78yA/r3ZDoGmv/Wczs/M93g/hTJV1UkvtoOL7Rigd
LlASjKVs2XlJAQakmVpw2JswwLaE9DsOpoSCnPdp3iqqOS72zThNDlQXlzvDpQMj
BQT79GMatH6IKN2WVjlscfSOXL++BOiYKP4X7tKbVFOJr0lv7IknbSWPcdmXlJvl
Es36R7fNuz6NX+icSoFnjBQQho7gm99uzm+S09JnJUYaFohie0gSZARCk/scVSBt
IQeS/DvXgEZgsbIqP1kUlZRRhymHT7mhrrA7jzRgqMK706zV6obkoAYUab9mKe4P
T0sGxPnsVVIjdnDDEqK9M1sW2oTWW1kmWg9h4EwQ5L4LHTdUakOm2N3hdtHzSoMD
07bcdVy9H/uWnuhfQFGxyCMw4ikHLbit0GdfwILDjFHxFE+HbRtKzPCWPcWZnPa9
5EYjXdrxsR6LRDR4wuJ+Lj+hk2UFG7K3eLa06T23+lo7tHDSL/BYxNw0XLpl/H+s
nJXq4F09ZhV77WgY2sxilH8JrDxZstdXGTJT/s71xfp6Pqicqh3V6Ow4+87VA8o2
NkSzHeZCilfe0raH5ViYn+iy+8KeqOTZSMWHTpAfIev49gXDUVF1GGhbrMGP/fvT
yZPUtAIzBbx2MfCEhGynhHh/KIRsUXVtS0bFA2FKyRPe4vZfbVh2M10MQ4fZnO1Q
uFJ6Pk4z0Nq72rpgf5zf7OBUFxzZwm7cL1js/EZpaRO3XDNfmZyxaDxqUF9s/J4S
hqCiYPdevJnuAI7wgD0A1HtGkeiOXQJIQ/uMm/4eQRU9cDjaey37DAkU5CzmssZP
qpWRaTXbqx1TwhUspJ5I1fNkTQKy2WSnzQIuedv3tUhvgspIZF6dbKdcE60EoX5d
mR2tTnT+ewv0RWw/xussZbd21lrlzVEsVpKrR8dX549VALd7IMMNS0x9y/KYs29Q
4L+3d65WwvNjld3xP2RQ0jFHhH3Um59GCTBMNCAsgpyhG4k6jd/ew1W5DEFEEaDP
e+KsEck/KjW7Pi4DpiAck4THhPayHybF1oV0Kdw5UN/FnhNq5WW1v+TIcKxwsEhf
4ObUhwHo6BBcDTPTRamBzbCNWDM2rTqbJ7uMMX2F+2MUBU4xo9fTMwakywuLMB58
VqjpHl+Fq4d7BPqqobGWFy6A0tHk0T6Wcnp5ZYrNfYTWLhQx/wsJbxB9C5tClXcJ
rfXC9hsg2paUMuptzUlFA16Jo9aImR2GMMMRNBYxWwRqQ8MENQOboAENTFq3dXgZ
Squ5OUrCtv1kWJBhKsfb2qfUEHwo9eFsyN/RTlYsCBcG7ofMg21sLkMcMr8Ot0yx
n7+wUegqd0Koo30GaOte3CuCwComQxerzCcJm/it5kCEwnUOMHlVayuRLfJ17kum
tu6JDXyzsntJnIRTkMCuQWNlI3XyJyZm9iYb1iByf1yejphWPOsshIi+KzaHyex0
9K2DZHnBgi9FJbkd1sJVoe0Isq2/S+CbyYNND1GP3JVrsckBIzypdmoUwYTDSc0d
LcE6pplNKqiL8DmOtkh/VXpBBQo0TinC+5juCEKR2VZFLb+Sldxidy15Uni5VzX+
BZnnAVDeDUhHfN1pyHhWvuKvo4BN6EWxl/GiuFIQdZHOV+0zQrrJAMsqrTDgs7fs
RFv3rOZpY+xwbMP298Kov3RM0KKUEFc0rQK39Nq6drld104h5i/9aCWkyRreGhj6
Lsvcb2hYKtv7t8xAPxw5xN8yFpHWuVmn2j3A4bs0Ca9+vm9i+/NW4lHSihy+wz7p
FNmgv/P6hCdIcdje6afuJJ91V5+hBg7rDCaQqn6uc/W4NlIW1Ih9k6dKClHwIoS8
KRi17gNyo3WRr9PwUeE+elcGfiKGusk/WxZQ3ohFzILwQaOmXZlPGet77sBhHW+k
tilGIu0LXpOosQPro4VIrO03oLQetw0gp7H5sbrPvU0zDS9M2ioK17fWgXznxg7E
InrngX36eeSMb5Q3EYnSI49U6bjMgyIn8VsaPLbp++jrrbbubhHBozmLKv+0P2sL
uD3uVOoJ5WrKhLprn/7et4QzJeBECey/fWuI//oBnFpR0hvSqYHVA+0E8d9iPwwD
l9D+nMR7tIxqFUR6qk7DpAZ68X1i1zUZcm0Mg1u/3kG9OXDXPAzh1z462N8VPgEH
KdKp88AcUZx/3bKt+H9Kg+WKuX0f5ama3ZsuwblGU9KLrE62ux5nDMi7gSDsYHuy
a5D440q/tbLTHArksTTk6kypiwbzYHeScuv0ek6AIvFf3pIADE3INVGR9W3gZKe9
QeMZUoq0id2hgm7Z6lheuol/SKxDk/0IeIJKvHXUTSGqOmNzOiGFkUUkZjXOBLr9
f++YGfHcV+6j1C6Fez734bLCnC5TekUcrMJP26OGUG0V92n/84P7Y6+uuP3VtcyD
6s80ww0A/cR0O2i8FHop1qTIZ4Zh5eNrwE5Bhy5naS99IFgq+vPiJDwzVdTi7V6q
WBVki1zKHFoHlaIyl/m/m7hc2i/nyoNteR5v7VTIUAjufVSfTkR4GbHmpqDPf5Kj
TZpfpOjAR4F3gBxUHFSCS1R+bH4fhYfMcUurAPuHK5QIeray4pcaufttbiRMKbfv
sQ1TJgr30dg7+5MDa8vwCqce4S9YUMtHl8WXh9glD5svouSuwXzGnd5RzrjpHN7g
Wxw/L6M65NriZFlN90z2IAcBKaqa2PUe2fw9jBvUcDpjp6B9xSfh0knhXkYTSQ0m
01UM/Amb3gCpQFAmQtmMWAqPojztAOCEKLXoGC52yKpeYqfCjjysgZtX7bcarQ+Z
dhxLR26FpsRuNUoaZZ5fQlNJSMaS/OT98IwsfqXQzGCDhWwpkWCjSJlCyhWpxWA+
oz/7Tk5GK4kAU3ee8QfVJ4V/OQyKeqe5XZ1nLBNJqXcUy7JB/OYClrvC5OzbYHR+
6doBTMswmBixZBNn/YDvyJxRWoVLdXVzfzcFUCvCWFPBRU33CCVR8Xkd7F+At8tV
BMIe+hqSW6lFfx3ELeuqiXk5642CPuG0KfHfQNypw/wNOvOW+VFCoXsLNh+/miRW
xUnUTb0d9rocgtzqAqaxK/YKhna2XcQbrq/shK/75AgJnl8Uzs6m+KW2fp9+S736
3zUhE0xnzleQF12KuQz4rICDviA7f5bm6MCKCrrE6Kb6C2m5Kxu2/iL+0/PHtzYM
2WKDVOQkMWhwoi3J6aYiBFOoTB+mHnpQ35UvZUvSxsGhesj5LA6I1arXklKWKxvA
lhdSRKVM9uftxTXNhfhazOCbWKxMfT3o7J7g58ZEPJJlA31O8m25xpJxL4R1zmJB
5DgfYc06+BjLvpDqX6Yy82IGwh2qEmHgXPgTphOznKTKbRComhhaw8C9jLg/R3VU
RT845HpBZouVNQgpKi2UcFAzwgzrm+K24czDNCrdlCqpBl4nYUJATxdHenXFQvti
iUfYivSxPnN3ogOK/EerGBvrDanjAW52wc0SnCbbiK7pMapz/pFH1kF5dyVgUJ3E
0T7E85ZvyTcjMeGV2x7DXyalB6tci+fsSBj1Z6UC2Kl52Oa7H8EultJQviMuWz0d
zdtfJL6hDKFe9FN3zU7nLK3v53aR+votwzUZPblsZrSCFxI+6PPCLdOVoEPGvO1+
K3GQBtQknS995Z7xeT9xP0K4SsnnYv5X/R5vUPiVB7MPOBlAveG5PWo5Kk3+m/Xr
58f4rbNUDl3jm60Gaq3lbx8YuLJ38M84DEFcx4C1Cb2BcOKr2gjVllSByW4YTTcA
wPY3lMTDucFB7Q5EHhcyx3fKHg88k64XzCuJo0GC7hxjwwo8ucquw/dKrBlDdDDb
z5QOWbOj9d/3lF+OmquzIE+RWGcFErToLfMfrkKjvkCzWrlTdtvfJaPeDWtJ+3ke
Dznniz3/JrJVLuyXgX8yTfBTC4K9+QQ8Z9nvMsW+fJQajh6gruhWC8EKHArRN9qR
vTnmEi7sRatTo5OU0Nq/AGwefkTq2Yg6TuuTjtQXgtCpNQRILJcFxVxWeEirhj7c
CZW08ZFO59OOWa0E+v2sCzQqu14NW8xc+ORMoTipklyRlumc839vQLxENyPwlyxL
HW6wQyAGPU2iOaOrWN+wusGtbOCYNWgwnniSFcGVU2jmxbt1TZ9q2GLBvizK1Vb3
SssgdVryLQWOEVrVfmV/x2BntKUJNG4O9gycZrr5+UyWJanhWoseIfXBAQGnjHxi
ingy9s4PQPVN5kvn8CMh7UigUMFcdMhBEfsYr7jFFgLm90NnEjxKlzufIgTt6H6d
xikcg4yj+GhRgoxqLaxpjzNzANoJW39DoheCYDJBdgCbrI5/J40SDuxV9YESGD6r
8VGaHjJUqwUW9eeHm+irQCG8N8U3brOmSMzT6bogylZBPegwTakXu+aTuO+eCyg5
hf9ZvUAmM3zjDPgTZM4jaiK5az2kdHr9AfaMg/Jv8wGALBW7T//fjLhGrLbIezvx
8kicd7n08D/hRNUWHuTRuQ4GEND94x+uZpORkEBItGapGj6f2E1t/RAjdNEtYZtk
7kJjVu8fJ96ntkGmbzGhZa5i1oJS0RMkr79RwX9IUM0SE2Qfuy1PgRWpWAB0kFiC
6pa9+YqLpSOzqg+i9g17Qilfl5y20U+DotwAwJ2dSkzH8Ezh6mnoK/HsMK+hW+B0
P61IFs2jdGZQgN+XLzpU1Kze2P24kVnHWXXIYhJ74SYrZ147dhU5O0ImzZrAUl8H
OjVUrDz186nHEqhlbTGII1ZJy9QWnkIhbVlSWq4fzyk5dm7oRrjaQWPIcOuNDSyR
qE9e1l710111ALyxSc1zB/udgQgbKyGfjScj6jp0HedCLk30+Wh1wmaPaVSpLCW6
4tmx3wb6wHuOCgLhMMRF20AyX3wKmZ3mT29HqbFGkX/VOU+7tx/Rve+dfAy35sFs
bUryxubi55xvWxCfEZqJ6AjxP/HbEDVw1kx/76UOVpfSjSNJjBgyknzrlbD5Dw7i
kpjYJGAPPnlcbkHm2RVbeDF1vUI2UzBglbopxsEF8DuFTLQHQLAOJgrwhdmUmRFR
524jyyUCc2FjfepiwakhQTJtt2Q5BriOzyeiPDV9je1kEQ2hxRV+RX/8eu7Qcca6
ZMAeLeuotelSHB5+zp5/CnRZ30V0q+n9zCxcsFOEbzH6ULoDxeuOPy4lBF6KKgBE
Xa27Z0fBDBQfM+zZB5tmXjgJtMuAk1+eUC+b/SkS0Q1YCjCVltQpXw/eHOLmgboX
x+5VhW3r0y4Lw8e+f1/M7Uj6vZIdEiNpdvRWsaXA6XGaGQ1+a4GVOLR0zwM7SpjX
lSFIddV4CVsWmxHcsDQ+oY4Cc+/OF0j6O4SbW5V6Zd/tsMc1p1ByTj/4M9+YhCdn
lDmAubIz/DcPRq/bSQ9dRr99qBGLEr0htEjI1E2E1csrYUQSqMH9J0y/0DIJbKXl
nh9qd0fe8LkxQAaMTDo8WXuFOSeL88z58mrR/SmgUUYXELw8c8e0Gq3mKrYGj+6p
50ueWBNlww1A6tlk/VYNU9oSLGyaK0hlI4US+khxz0AhCWq0jF6ViwTHPIYfA8bh
JSkgZM4pSEyG25RGVhS0q71U+8B+fru2i+lJF1xvFJej/KdlMPCW13DiGDIUEO+z
SA1GRPqSbiNPn2yRkuz6rYTki7C7C+xCTW3t/8KgD7kD1Dy8RLn69dL2qarAEM+z
VFxp7c3m/jmYoDxaOO88pDTc1TyFhvOAE6xdoTNfULcAm1s3RqiQ9+xhUIuELAl+
t7g8LS/NamC0yAKZourbNoHEhgvOppcUPel9YF2Hf2aJ48mz4/AG1LYJGkwHfP+n
gZjtGcRqUJcOMTNno2ICiBdJfEmhyBH28OHYJ9MSrqJn7Is3uwjfVYw6B5zJd9rI
1JGfiLG6mo9EjRDw1sjjpWIYGVMcCHE0sKAdDBm569+iRZ3unsIv8iWy/5mnGBQ3
/gd/SSXfjaBVbxiZ4Kz2FnJe0BzrjWSQ3eiObepyh3Eg4YPzYggNRTr+ODrcsCsO
4or0G0n3eA8m8TuftcIbjFdty66BwKzmvQD7w5hJBAfK38rqoSLCrGb+cl+FHYBY
wrK/85jVpCKM8SfNAol2jNQBI7Q4p0dZWurTwx0tc1wcSAzE2zsdmu8ZY8tl07sB
vdoFAdPfnEcYJdQnfMNAgCrrzxkk4gj6fLpV+AIfF82c2YvnPrq0xAsL6zu52f+b
R4vpuvY2g+3V3nvOoD1ZIF9AfqMObcPCx1/Mnk8NVGqdany96s/Qbk+DaEyFPsrm
vxBx6HIpPWSxdyU7blREsgZZOt05Zblgu1alD6HkZrDYewnqrWYIWAfvqoBArOoS
jwunF3H6j2pcRQRvUMP9LCw9oHum6+91zoSep3mMjSM5rHwRu6Kwv2PPhwglcUc4
lBhBgwgDlT5POJKFGtaNAN0Vdg61zs9/90OrpoiX69b9cujWy9cpjTI1T/5rgov8
Zy7yGsQeoecToCivMt9Vk62JLHU2RR8EbcE5JYbA07dIa2yAumHbQFr4WIl62N2d
y2JoEkD8c6Ap0ypyv/zDV9iYa4roRiMoaUwtu6mNb15qn43rXsAwUxYckUCovgS+
Nbqk1s0Q5d4yn4BRs3AdOCA7mAZvYbT4D7cEXJPhZ/ArXwgDWhQRlZPIYd/auRaZ
V71zb+sJctIDk595HRiy+hD5XquKPqfXLhyARxCI5nHFxgE29qVD2dH2d2waTbdg
lf3NQNgg+bBcW9HuCPEmvCPvU2ObZzjiM8qwZ77QTzhFF9f4vQ3qcEFJpkeDbhCD
U5+JL/QeI/S1JKjlGE/A5uKxhRGvNq0JCCaC3YtUJjiuU9bcKy9T7rUV7Mk6ITK+
bF06Eqe/cAipESyR8YDiOvmU2TmfcepzvaUcQfA0I8+k+uGJK/N9ZQ/Fa3MVKrbW
bjvqc8uC55T4qV0mHoRGRpGIKURx0o2yPsQfAsLPB5jgDolbokaGkGS9YTfY8W5A
0lSbVDJVlqXcAevvJSHXzBtXGNqlA5fkq36SNfbwdDQufbEabPCiJ0D3WSBsov8Q
g4Nj9U9KcUD+mJT29z76oSamhQ3fobM0kiA+BXwjGvi5aW4mqgnQN5yvCXs/Zk3K
T6Rih9zbv+AStmRKfcRnBSTzTGifgIV1DJODEiEJPJBLPLFz6rMoEE43boIR8Bos
fBi/BG0kivfb3P9gIqBvEiwKZmRxxNl8mm0N2hZmLKUy5rQgHi3EHHKRnYSC6McK
b8Ek6z30J3l7ACvj0MTI29rDXah4wobyoDRnndBhIAxApGF1jH7lskZEOR7jqqWF
VnB/f5DYMhPHrNQ0b4zDFWqoac9N5dwDAAi97O+2Z+odL8MVGWReXQwu9J8XGIRt
DpAkH5ezzoS7BUQa9KP6cxqu5lD4CfuBx9VkljevikWVkbBfxtW2l5O0cCeZHiBK
c97JCZU6d2HxIs2hHMtj95l+JxbFo69A88kp37tdnbNYqMURf33ReLlVXbnyAOCt
4XNUS3oPMbEYlzC6nfbYTwKtpx5jJDHJWs9iZOWdTsQzDru2f9z56Ac6At7TbriH
kUnmN4aJBgYFvltu+BRhFXIcYX19IRN3XW4ibeXD02FJm2fjpTIpVsGDCjLUIPce
6O/VYx3eFrRQ7KEwgYZhFRsBflo7lC/eLkHNq0u5m9SJM0A9IyXJCaaPmW30AU+g
MJIVKe5gJ9CS+SuE8K9tzatgBYVxGriTn3jFwTlhZzd8InB53oQ2sE90mUg9+mt2
TUMlmqkIwnzPakgww11g4zTUHlDt6OI3TfdQ/fmgCm68C8BEpQsZiJeK6X/lfuuc
0jlddihvDNSh+FxEPqaB/iRO13yqJOek/KnjSCjQIWIZYFiCcPWSjHiomFHQzQdi
O6F9hhmNqZA4IpAsDNijVoegzEt9JgWJcdI3vVBBvU84QAgadyuvF14mZq4UxR2p
MWp5andjPTMysORlDfpsgclevhG4YqzdCyRFjb5vgHtkhFDR5qU9JTIjNgXE8gtP
+ADy7EKhLhFmHLfmmgTKEU4cge0kS8EA3e1GcbjRNdRiy2xl4Ew6DPXjwXW9DFxo
MmC49zkWHoFq+W74PubQQBBsGRaRdAepWEBt+PU0DLJXMtE5/TqwSVUsmemfetPf
sZF3Z7/TMeFN2OJn4SjtFqiCSCf9mvOihccm3vKB1YV6bpaA+6qpoeasR7ClZA34
EtIVrBX1ATOtQtl5TjmOyWWGLTW9trEaNEERW/4LhvaQ5LoxFuESKRkM9Su3cZ7+
SAPivoY9azMVJW22w8suW024JysKs5n2ghgmcx8IZqA4btGQoex8tPfzx2ZEmcH+
d77mVcHwu2N7cEDLie4evb4TlJ+pNvQPGeIlZgqLI3bKwrbN0uypIDey/mKbhnN2
/chL5JFAws/2O74hFIBaRTem9FVrqMR33FK+MFVg0jddqZLthCKviakUHnezjP/A
g83mJShPJw8hxTB634nlZArOpGyeAP1RoMzJpg+YYr8VHVjxVb4f2ZMe8oe11JA1
uEVgsIZraKiFLrhXK1SxxfJmgaIj2buNmHa+jLYasRkwl0tCai9i5T7vcgSxpHuC
lsmUhi4XJGvaZdsrsuqs4Ihgl4iTg3Q4n+JmenywSA/kdgBNpx8NGvKEayxQuIpH
vvFu4FjusEFpTzM65tGsCoSyDgXuLR0QBa68Y5SX4MnPDOkr67cAr6gzrj3AxnZ5
ysUGul2o/y1ncFIzCoRC1YOKCXm9dCDt5NBMUTEIkzpjm87k9IOA+P83iR7pAst1
DG5wIGIe5BoV1Jmn1Hl188op9XJYwyKR7uiJXiiSpbQMrIclUUDn/xXocnuL/bNB
yBBd4bXvucacI/tCkJpKLmnnvp2e7zkSikBRdOmrmSx91a9PCSH3s+hFAw93xiyl
WqfB4+q8QhLvha1ivI9rT8t/5h51iG1kfYq/8hjMezhGAyN05VZiquNwt6X9rBCQ
Thzh+VIyPMBrNalQhiKmamacOq3Re5Ta7sCfJfPwd0UxXVq7VSoYcfUOHJ6VyVwW
qHyaZvuesWKNnwZrwrPYkUP2fY+35PzRn4SgMYBL/a8WPt/N+oPVmRDCO/hRsYLF
KYs0K1SXXvv0MfBxTkzfAlltzLlQrIbxw2IaANZgTnl3zrKog1f9jnwY4Xd1AtgT
mwqlFzgl+zYMtVZULQRXUBAEZA3InH/KRCOHoNPN2p8+xWm8Z9j2vrcuQ90ORY+5
S8tcq1vN91yHz5pQCI8s1ajKvyYaCxj4fU4RCET4AIPnk70TmuLXqtBPNGSF37eP
yUOz5l/qzQrx1NuiUdQ5OEn2EbJKsOZ5LaBNF2g4ls2DWYYYKGHjjAUX5RdhrKxe
Muckd9kN3LVtonDXky6dv4VTo5bozWThnJbGAah867cLn8iLvkdJHHb+fhhKcgEb
1JpCOfF1SlJK5cJ0u6bK61ffa6POn57UTdBecu5CX79HzI2C1EX/PSpDOFxkHHLi
a0cwzlrxnxhrnCPLmlnBmcF3m4vIWWv7sHOrdjNQNYJbfRcyL9BZW1Ud9NCP+nJK
xFnjgT1u+BZ84wCvylmphSuc8ojk4bKerzCOezq40c66Ap0rrJ1kqi7CrGgnSBXg
pFALtjRoJV6D8Zc5AKHZNXY4ZKWaWgD9DcUSjfui/T98SSHfImciBjNexYCFl8UJ
dS0rOpqbJGPvx9E8elN+f32RBPuIpDcqlyAlRVgGgYu5VCP9rcFBmoGFejourQQ/
MXd6S6z0KaApyW314WKHEcV8y5hG6L19RKbepYf/BA910bo+Dg4iQZtxMlQjZfiN
LwV0EUfBooq02sGqLz3jLQJXGaTAWTdw9ZgV7mi2Z3BRHBzpQ/ivAxMrv9H5Hl8t
tnupwSY6CaSzSuen9ZoqZxp6CyETIoemYvURf0gfpzXHqDwzd+YOWBA/SaAErNnu
fLMiV8qTYKH8U7hwZB/J64b2HQS7tI0k1Afmz5RedkE9oHKG1MaRx/lsvWj20oM6
kiCw+35P69Q1/zdNaLdVgeyGg5fvX1cekEBenaK9u6gAoKQj8v6K1uLOXGQb5yqJ
/Nvz1ABt6OLXd7K4KtUhH7whbiyKsO+jdUjGvRGIFtk5PwUWlv8w2jGPEi4r5y0f
DSio0uQBXcID/KajRMiNh5H4ahzNCte/V7np5S7NZJU4AnOqqdw5egAmj366aTDI
sbPjdgp1hd/bqDB5gEuurbxWm4/CWJ0BuwKQIv7SMLSHNmnmfiOGW2g+XX/CjL3U
YHlZrUQtyN4D668Htj0snga2+K3+OubhDvsIfVrCyXa0jPd+M9ohRACY2UePFBZq
YSTkWFdtZPCFrY2yFSCxayoCIGt9dqMicefYWAvsLhgtNGrHfSZzRKrwfgBP5rGi
g+fQduK7UumVNQFOtvrA4oR2crsAumE2Wo0k7ZmvAsnimbbcxnqkGO7E4oQTSfZC
Q8ayvFHZuSXW672OOIEDYepk5giGzX5swlCXWuVtjUX7a9mE//+Jh1mkYA2gVSwp
rhrNv5kkoUYe0o8XdDmOe6jqoh/8olM/WRkDETZxMHLY1QBBQ57t/mu8IiA5f6VW
IlZ/mLXfKQcUjl+2hziDY0ifZPTf+kmD8pQm7vMQg0m6gTYdgVy1kSYYqa8wjSlQ
PcDDEJIMqNvQFKNRZtPET2+CtTAqnfuppngFHvH+TP5tbO+a2XMMuOOXW72tTMrD
dP3DEkpRdA7SvIDiuG+8fSMhHij98qsMeFrmd5Fm2XUcMn6tXMuRLOzQLLvRf99R
wY2GU20I55NwZVfF5sWJ/vlD5jpxT6QO07X+1J7qdKgFgI15lFqUmzPRp+wZ/TmE
fO9CzStGMiBRVzNIkVmkGQw/RelJPAu8DI5fsIgNZGxjk09Voq+BEn67Peg4722K
vBnvefGX6mRZdvDLiVgvBUDYOT84sBCo0js0Ofzvwl+PQbc495jEhT7FanjSe2ud
W0nHYq/vv17Y7ZIbqEMXZTx8/W8IxDLGvzsuiiGVAoYNddeJYeTqtUdT8py1a3oS
akCukPHheQ1vFkSteqcu+DZmQA8cjnlW0i7GLLofFOwzGFyW37ZYJWnatM4yYA+M
AemoaA0Pq1AOkOPfyobT+wUpgxUStKIKzcNIaru8OO5eWf2JqFuxnpG9202ULO9U
5p7MRrN/caFXNMw7CgXrgwlir54GVXIxZcQVVtrOoviQMklyyxjA/3ptDprOqsP8
4eb5c26gocY03vO8DD2k25XgjR37h+mVTiQaBrbNTCpMDuTeqh84nkmzBAEc+4PL
NAD8TG6ZNStcBpq8aKhiRkxLIoEJZD6yxG3dURM8CdStj/n3mgGkmZMlNJokqXQE
U9iRzG/Tk7866rByTGKVJdK1eOCI3rDZSMaWH+jkEt84k2roEcMoDKiCl3UhnLoz
mfROvC7keWLuzBl+fYBTeJGpa4YnaqwLxaTZCm4ESN5HsvMqmjvdQ33w8HLecn1Q
4J1jG0KIf/yM8CR/ffPlQscyMjq9hVUkcToXrKi1S7MLjaYOPA4q18VEW2DIwSrI
DxPiVYA7YyECRadoIDdB7WETk/FdZcRrnR3j7uXTGrHKLjfDxeadDKeT1mYYQDox
7+b7i3gAexZCk6ja//PzYeDK3GF6LYsYlQapayjBMoSN8jU3PW90hM79Q3BkVIiG
YIE6TGw5plzpfjFfAIg0/SPbWKTRYn9u4byFQ58OUgt8wCR1kalpMOjlMkq/l/HB
731dHe9+CCS0jAAAecm46snqYgiiBcMc1pmIFMPICD3ZQNVKH/QmG92q9mOS7Pyh
KT+cxvQ0Nr43c8JjOSsCnzi2jbTVyOUUQvWRXPl+lfuWsCul7ALqgKPaNzzt2QEf
PWf5pVI7hObvDvqda5FOkZst6Sqndd2Y7KrYk36X24yuQD+VX71E9+RFFd3sx3s1
gCh0gsiMb4cl6dJgKdXihDUXgXCzdWMrMRpk6tCADWCxqB3CkrVZEmdNPuVdbeRF
bzXCD3CRS6KLN+QQvNiq49BgYO+wP2nTgYl/M0zn+UGyNsCNxZ1UhBkNGzTRDZXz
9mpye6PLFLYe2DBp5TnS4r7VKuFHjH3D0b67ofJsIl3PzRGCCUN79Ph6Zabgncur
Z/N5B7Jj5iihDbt+5jPsr6bBcHn4l3rlnbvCgLRDako9DBx39Sgxb6ZMy/yDp9fV
/NFyLE/1MWanALOZ3h915+pbCJBDpEOFnVgrUjVrNKNU0i6wtWmTAEb0m4mYXS8R
3tjya5a9EHAgqARFWPjvdbJ5NbmoBzvwgsjIvYftPAzMPiJDOVuGsxb2wYYwJ0Fb
+QoG0uR6II0/fYKlVEdBRX1PfUUL5kAHAZzvMRW7xU1FWZ0+o/d50OIvD5DG0Vzi
LShPJSKAB6kXniBQG7ITqXB7UjlWt3vyq7hYS5ZONBd3TprZdJ66gzAaXoYfCylz
ejhapKOHm92n66YiyacbDURMJ9d80QtzBzJCO60rbhAlkhQRYkS93RoMOBXWAuGh
CoBFwOdTs5GNDjtfxPopzR1UfzdCC6L3uHkLnI0JNOx0phP5Ci9Sg+2Qbgyprjzf
CIuK6o7qshFrh2+DFHnyzeVV19m46KRZfwBsW9KK2fMH2d34gUfFygaQev0JP7nF
DSFMlV59i4witSBDrg5ep6ynbWlYYNpBB2B9VMDNQBT+OaDcjzfjFUc2oOoCMd0j
e+aN6Bj8ySOwLChzxO9jYx/sdCOxy7LYejtx5nRjEoeGGueswYSfLxzeofuQ1N1g
i9E90ttKYGzoi2+Ag4U6Pp6eCPhFdngDaJw8UOZOV3leVuU7kj/B7Y85dSlCBifZ
bxgpFjJjLiuLU64aqF54hHMLuVeEGAxLssfhM99+2QHBNwhlxLg+nHAMo+Bx2fjX
snQ5FjVfiojnnnihlf4a8AHt0CZRxRhH80u93XsV51V5jtckOTITSyDSTOo3PacD
lhBeOHPRytwmmlkYskGxAUs2mosHO6UoJEtg40xVjLgOMtkCw6yfR1t2QkhI+Vt0
MYUJVyX83+5hSmbmi0G/2E9p7ZMzH7AEzgyFhBN6lH6pGxCNtAyJGKfDHJInM5Wr
YonlWyOnR08cTN9XxC6zeSy8/cxWU5tm4IDEzV/NpQuV8p+UWJAVFfPoEg7OO5bU
USVkLR1gRjSeiEw+jROis4cywtNYkUiOQQmnzD8LbqIGB9Yt2tuaR5sQsTc/JyU7
i3ZBstnMgH4XRtR/LxZe2rB8pdDNlSn26UztSShhcn+F8txY6lJFkxuM4NcGLRIv
eusbJSaE5fz5rAaeZkfv9ba40tpgoZwHfZ9H1djpqgYxkrqgK+MV4nhoSsOomeDa
ifFSiL4qMK/ZGJ9nOySVFq0dhfP/OQmzHC5tyBF8cULEcHmx/iSdP8T1XjIGEa0y
RelnK2pEB+xjM0p4Gh8uNP/RYnOhA2WYF5S3fuOuqsAoAHKgTl8TJfvPW07P2PBy
sT5a4r2TriOLZWAgBf7bK1y+9QcAWnrNC31h4kWlmS55h2QrNy7YrEAoXL//PIDm
peQkSVCXv7zfu05HCC7HiIf07FiAi52LB508/vD0tAQalxKJ+/98sF+zeF1VWAkW
BkCDVIP5lNeS1pvZr0PkyhqU/aQlSKaUChdZKcQm/t/z6oMCphQQWWeD4nJkslhV
E5Wzg2Nj4nOOZZ/IcAq+f+4b3SamwmCQ2DykbZZXTsdzlzvHIvrjzQ7ZFkjSXeYF
mpnIKk4JX6P/7vbmUlM8CiUu0nlyLsetTsul5xCOyzGo0oLYL9uvoI6/bcgCfC5c
FmIJ0AYOds5gP6in34XfbAmq/MwzzeMEB4ePOZZFCnY2w5HaY/nPvTQo6n7ra2mi
QC4hhGNEJ6Oeyem7KFkW4u7KxAgu1avIwcS6yLtISI/UJq39wCx47tap7KBXMYT6
JCW54EYc6Tfvyg6knUSbDVpCaouXn9gVPErjdc6gOjMPFyBwhn9JWZzTEa0a2vTM
c4ErxqvrQOWe05P94a44t6LtJ9VHCZCCThi2mHPhWwMCaKE585uAhH9TS/LXrk+K
T0HQod6MDMRDUWgvAN8VKdxfxvbfFOh2OUjwrv7YBLkEz7XxTmq4UZNlZa+SWUDg
seBGmzCWn/AzsfsZ0zcm0jSCVf9hCs5aTw59UwZcy8njriAy3qHR/oNyAmpMBxg1
e+2AdwBPlt0OfyzqGq60E/k+NDT8UDAJ6o8dCggPA5k2P5d/daXn6+iyH8fSLiNR
Ot3sqzVcJPCVlwMfnUEpC4WVJqvZgepjaE9bZ5U8mfa68B85HjoLFH4bLqpEXGXh
egBSg/XoH17aLPc62nAj1XTT2ZDzEpTtblWRWKLzXglvCIPxutGTzWfJJRNxzkTt
OBjcBUcMNPDvWnSybWRq8Je/LsOXw6mzv7tliGRHSEd8HgQny+amX+sQkuksvwTX
3B0TGENIFG+PUDQAzwDtU0MQcOvtXiI2B9NNaj6orzkQUMf008fHuik5i6H/C2L2
Q38o7p+gWasojVzk+C0r5XjPpmSSmegbUm6C3etA75gX9ZPJBpiWC07g/AlTnbEE
QjAVU6GnhANmL1LfhLtDvHGAmdu+uvqRpRdXrv6L7rgYhsNQjRdtoHrZ1j4BN/Qk
DooO/gBAOE4Bipl+U2cf/u//vdPcqexSRs8nUFhdq2E+fwvBNwqyKGmGlgioBDIO
zsPG9E+bBR7BC7+SEsLTgW7MPiTq+q2vAXG3x+SpbrJ3IJQQB3T9uQfYDynisbx9
cTSI4T9FIdmNz6nNjeMULQklMJQNGv72KPynWgv7ifk9DFslTkZL3fZRRyRxrFQz
MHiTzKifasoeEp+mS5dHVl6vjRiNHg5WCaeRQQKge9BPyD64rP/xKW4iV3JBi2o4
PAJpbTUbzOjatCstVjWF7wYjZhRo8FNRU5RYWt/+9fxYytVRzrKSMjdU7gqfpvfO
mex759N8JwLWna/2QXusRa/ak7Oaoza+lMx1kzCN9DJ0wiN4Q5of8QvEuoZlN04K
W99ONPJWU469hpGx30f+0hJ+pZuU/8lnKWyu0mC+9kyhVtMW4KgV5gsdK6q8mAwO
dBhJuIQNn+6Z8iKqNDPDrup95AoaFWxWMtfNeJdonW2WkGHurEUjkDVGTNNx8ncG
vOqtnz+ApGhocoYKjXXBMJrhcFQknqm1W+i2ZqpBACRTB6JJfHvQGzJfJdWbdI0F
220wq7xt+dWHwz5lHrEO/gGRZCe9ICbJBaUgPduDG0nL1fwMHNys+JDCgpwj2nbW
OqWcTO+qbsM2A4No1zKw/TFL6iIw1gVh4wdqV/9csm1mcZyi8kIT0qsVCwJa3L+U
JafyLBfnBna5BeleY538xvWg+pMt0jcJ7fznUjEFHr1nmGT0CM3JrhJjn2qNpe6j
W9l9ujRCMLTbXNmAwnK3zXznravPJzVILmwPYPYhVoL57nxt74A5lFDQhBnL+Vmq
M6DobMfZ/iztn5xmhKbF2SFYe3X3qUejFZCV7qcsNg2EW0ZcEW7HcgwWMkpGkJMh
t4nsdrd7WRMsqOdkxo8Faycc2DdnLTOeQKrdVWSLjv4h2NzDe6S/s3nTr7VsUpxr
bRxkJNdw+HBQ24CFcsqrXCdxt8nBgKG1qy1hpuKR/71+bWpArSjk7PC6ke04Kfic
dG4AE3+TuqoJKiMFDuEGIBbukIDe8JV+mnibRro8itDSruRb6Ext4ENiFHcja4+E
seq21wO+I4VwQBUxZ+1WYy0FjrF/P9aKq+ZVy9Ne5ce7zW0JmESKAuiNmzHdsEjD
elPnxB2F6KlE2GH6TUVNcBcEygUyUBKXgHt4/vBAD911sqofntRM52CWKOL37DYx
f1p7yM5SLaigGImudtkxumYfzGcmzOsp5TR52Mbl/hs1vsAvncLpg5ay6harTqKy
kQ77mvAOrkW+Apve7kwzZRTYwvHHzH3QbhF+QaNRLinmBzCirZCfLkaGmJwoPoUb
ZMKuApwGXlwiGfkT0UOdeXT8PMZrO9JyzguwTIJ+EVHukVwIkwapJ0OrpxtUId5u
rG4DngHmGmrTKLguLUp8NSHn91MyerkfZOWLakd5PKqAYHnD9S/QgyPwrRn2ZXt2
9Lkki7Axtp5rIQhHjdU5TXmYfnI+8xhGFyRRkd/f2+BZz8bZLgmLIgwMjFHKsj6L
CX6HJxmLm4M58y9lCxvIF6j962j15g2039yAFzsIF3qms3dE9EMDOZXN0Vs0TKaa
Ij8sRDJla1Iy3gfk1kY7w/6zJOL5pWAlwPiMatLJDUuqg48CUBLtSc+wBgXNTaGE
aGnGRei432VdgNxRS+tU1s9URKbzf+fCu/hq00q8/lXuxW8UG3CNnRP7gAc4UNXM
/Cajd/kRvZnpAeAhFIqqCyjTLzVo9vmRLac7+ZKoaF4jzF0VUGzYcTP7lM6AyIBy
YUe1vXUho3Gl0OWThWrLXQExeSyTlT2NNvW5+j2QkBhf0ebgwwQ0xdR1lb5tIPwo
8dr8Mrba6VK7pW+qJYJHdBVBYp4o91xp/7FTO3KtDoPFWlX080hJvHjDO4WnAQEB
zT3gjtr62pgqE/OHf0gupub/+iUJGvC7xEve3EV0a7hcLsju/50sg8goneIt8Cb6
hTyNObbcFoY48lHbojlybadRaOYj82fcjQPh7DRYVcriwD8rVBrcaSLBDRquOsez
K27YXlkyi5GH4M+C4twq9kdzDWvfjR6pX/jNPC+j2RkG4AHEmlR2j4SG4kuEogkY
defYDTeOSrnYrb0VP1hCrXRPVuKGZiUyNhBaV8ax57m/muD8nj8r3vNF5/VaTvaW
EeUYL4TUNDe8HNvIfuPdzFOwKUYRkoEByUeMplvtz/JSEkQX0EmBvrbSN5AI0DNP
Z4+mxqKeePtV9ugiOifTelMYGXwiMYaFPFSig0uUFcSlA3PFuEht/O9ty3L+5Lki
ORV0dMiP5BgFVDZMWME1wHQpBTI027JFNCFptpu/8PCdVPY2RTivvFCHCOGO97xh
eLPXD0xoJ1uPRGtwz6qPzbIWe9mkrdgW7AUqEA2hK8zLrU8NQ4NYpQDGa/elyOle
jUpuEIkSfmQexlzdcdUbUnt0GdF264xzVDvP0x1tz1pHiuLPOLL25XXtDlKAYGAw
93l28xqZSm6euGxcRgg79RGq6nlUtlHOC1gtXoYeCA8E8ndILH3s+Sd/HtzacFQR
aGBbifO6xXTGdfSWOEOUJ/osm6rIWaAtN0SobKUnGmis3MULrIB4zTqUhdb9rXzh
Ps8QuL15Dz+DzwHxjLR07nW28Udpmh1u4ChFSwG1jaA3P0GzBLDybReMyfl2xUdZ
phoRKvmrvQ55Uq13pFpEXNqyQJV0VE5osL6LqyCzTJuifRnCLrwvX+l5VzLIoPUZ
S6zyXCEUOxA+J92/ehwgMkTdTMBO34a+Y/u+VmckWWUUFMkWwgCzucey3YIbMclO
eODSXZgXzQRpWJN0mrwXEvOoUKsDz2T5P7zYRFKcgxwC3yPOmuleJ3SXoiVv/HbG
9+IO/xPqmkW1endSnrxJGBfFYdXxIU0DZuItcxzHUln4HR7TQuccAmqKgDSn9dRJ
YE+ozNGM87ENn4uXtYuSrK669AHGaIqup2HF00rY4Oqq+UpfpEtoGB0TeU6zdSaz
AO9LU3pffJcr1X4+VwpBA0Ine5AzX6hymsYBO4hHdd3s0h9ORY5KE/43xvHqKQpS
SmubD/f7fkVOPPGMMBEzf+d45/46KgNv/S/fXKHon1bCK5fsP6W9ga18h/HkR7L2
hzfTswn1kYDKDO0pMT4SszR8RUd8T+8hJn7QuAiHJbhrbrqIvOMvkM9wL4qwkHMb
7wmMU72vX9wPAvYiy5CCAniujk7VTsaat0EbdIEEu9KkHr85dZz7APWE04rWkIuS
Q7hAZNLnKLdPDuSS9lT5N8NfPhD9B3sZGFAUKL+k7qi1xrSfBJtHuTsrY3LQxe3e
fEAArG3TXP8KJvLX+S3T67IGg8A1tEaNqzSjw5ypueP3HAepweGcleseMtNkz2n4
W/h3nHbgqox4V/9TUsdGfHNorMocHSstoXVqsqpGMSWbFIE2r49v/MGSzRhS+LO6
4E5ha9XuIRLzZe1ZCPwcajPghAswmTvN9j+A2tTQW56fbpN0L9b+mTvAueKfNRxs
unoNGRE7Oj8vW25q6YiOJoZKSM7bOnsc6NiCFYVs6GitJHWrDn8A8p5x1G0p8ugL
OprCl37bN2qdXFloOmvODQZDDi8rusYpo3DbKl1LJFbzJnjrCjTxCMsrhl4ZSLTZ
/nKVoVnoIPRnAe+fwNujQQnBeckhzXXa6b0GysAXAifNSMkDcHTAJonFdC3e7noW
JTfIIa2tWMCKfv4ub1RXqFPwKgbQrI7YR/3I+lt2N5L4UoyB0XpyQwvXIJwNgLWN
cBE2LKFLwtqaBXmQVAk2Jzxav4lXOdEmiyXz0F9gzcsyG9JxbCE40UO6xvefCuVD
310+ukLNhxXpcOvJCanCeYCXfmiEm2kySA1YMhDfxbG7dLrqbPDs1rGHtcdTCjIv
k2XGeT1+xHsfEtA6gIG1PfeTCvmC0x5FpCV4wuM7ozWDy2cB5b7ZHfbbl8QUO8AF
T+jeU+lLiv4FT0GDdK9qm4SxBrEWqXtBodFa8ml2t4CerXyPQRmTqKUdFhk9UpE3
1nYO/ijn1vsQQTMHfDx0SLKaZZ0hpSIMIv5zp7I+PAn5iXgUnAdbG4XMxVoeAPnD
slmUva6qFcFg0eQXrbEgxf0vdgWHlKU9JvszAmN9+D+csZ3iz3Uz454q9NDXAAAM
h/qh674kKZTJUAisAq49y7qVYIyc4O4jeVV0Vu1VY1Hz5xAiMJvsWuaH/rrikrVZ
dyM/isB+y4Di+2ogbWm8ZNrIS2/0eweGPuSv44U/0s54AcF284nKhcq6b6VtvCgD
Fq+g+r5Y4vxS/4eM43l0J0OcLV964F+/2UVQWDLduetyT5nuQ/al5yRaFbuJZnAo
262g1c3O3yU9xhpAYLNV0pc/KgDMwjb+x5oCXYrYj4tYcQhpRgZRjTfhTSU/Mh26
c7cipcXvrSAXuwy9kChqu/68DibJAG5CgLvsnKaKTqzmLSzCTtB0at7LaIqN7yjb
aAskHtfPVvlXLgj6bjjioGLOvLQdglOjX+qipfCsM+gc+r+xXdI9vplurxaRVPr/
CicOk7JolFjHF5E9w61l8eKrzplVSrxQaHO5nHafUxwnYuXCfGwRbqvJ8sfghAWz
GhuvzCNCozszc30g4sKq+KOddQRC7R2NqK+WEdpwoVqOW7MTXtzhnAWFy0auMPAX
4jv/CKDVqhu90PPoSiBStOZxcgTazNstnH9gcVLOM9W/uZ9BfbcpM0PQn5mLgt0E
vyQ+eXIDYa0dbDsL4X8QFZXWDs+BspeHVoR794mWVwyiubbYrAZTHy6vDa0A/i0A
GfGRKUH8M4VcyK8crwWCsQUkHoiAGiHEXcgs342JqgWRBQYGmxlzLtyra4xNE8kG
h5y/TS18FraqrT60zLrMrq3wM3Hz1ws1kUaREP4aLGh+gEsXOKM6sje4wQJqfZfY
WfA3PxuKqjIJ7miLr3eA2KMR3yLxds8eovtk0R25yM0sdTTHlLMHQSLJ2Yf2uqJh
SFn6HyTtSBH+SykxdFgcy28vl6jyVz8QRhacKRBtGruIGrC6R2wC3aCi3ONuvtCM
8lqQkN1F64kkefYpWY9LLUCZdowrEqxDmA7PeSjgkraVnv2jWOvPYikrExfV+LBV
GitrYEMOdJfq4FtpA8K0dF35iPrCarXARZYs9Y1UX3D8ALFXMGdVOaKqFH8tPP6b
B2b2NQJqq3N5VjRbcIzrJaCWAeXyjPpEf6N8BYaGh6gs7hU8b4zGVAedSugqyGY6
LA2a1pCoyRIEhwgmlte36NCIlB5D3VDj0R0O+emSlS4Qo82vFLRFeTEkO93eku0I
Ehj9FJuZt3wttX1aMpsZSSy2BXxbxggl3iboTw2ZrYHLOc/UImPkbSckq9mKr6M+
eJy5YhpcGnxf/3XB+/sruBeXc0QeePo7nSY6cGOLTHv0Ep8ItCI0FB9tsSrBcifN
x+0sN2GEeSErU5ze5bo7pQpkj2N5cTES5mA7GLhOBs1EZnQF24Dq1kzS26De16SZ
vV+1m8PwuZIt4T06SPcJ3cimNDNUH6XAFWh1glfhsFz3vYuY7JGxslu1XH+MIuCt
Bs6d3UdftTuHxFD78PGN5RNET3BIqxRKMitjvpl6sZ0pExmNi1DoU6wbErt5CGV+
vbdLzsjqYO/ioGAF8aqohQv4Gq6vkSLA39UeKgNERpO92ltYXoEjJhk5k9/zUSt1
Kh1aXfA2oscLkx7y1s8OwP6rMTnc/4jAOMyJ1Tpt22MvHpH1pA9VPgmROEmerBI0
CUCrg87JMjwqJfysFBHi5s2Aei1plzqyZXwQNAtjzajF7c5PdrDFbTUKevXNbROL
cxAKofBmoXkXLMkjZaQnu+in+xGYsHIneqYGATEHzYRhlc2/oVkD2tP5Dd3aeqHq
qX2EOGHg7bGLyhNEh3k3osIObgvvyeJwyBfZHHCxYtbTYjMNn84ZygNu8tem6Y4u
3UkcsSbWGCJpQM4/xmB08PywfEo3PxmrgMDz2kS6UPip+jKi5DRGaF9o0/Oe2fYB
+zF4yXwLy20cQpzARa4fs1Xmu6P8lw7oP5J56ds4fW0/e5seQeA01N3BZuDNW1jD
K4PmFD3pfa1lCpmO0S7CHJ9QOpNY9PJp39Kb37XAHRjC2lw+wLH3DONrxR9tYkWe
ZWU4Tw2UnDN9ke2CbffBmfM2JVgyayY52meGMo1PAgzYUF7XnwgQGqDp44Dr5/h6
tC7dgxS2r9e/DsduaqgZt6bPEn+qx1EbJkcqTBg9EUetl5Aj43pnkoQfBsNaQdw/
y1wlKCcyDoXfCEGftN2qIAsfXPhh3Z7MsD1ihjswPIFV62Yf6LItRDwLnYzXJs0k
5Cy8Nee7AbmMVvgtdoGQWbPiE6tQJoIYmhw9uTtwhXn6oR+P8/nAfnCn/8EiDX+p
0dIQLTedHS/Zjhwmrp2ypffhxFHkI9miWEDXqWrhvrfqLfSg9R+KGKc8H+Huloml
uoLHZT/ExTnHyuq4Z4sRGncuQPgOSniC43trKfoKmNsLSFJ7sxBbwOoWJB/Jr1e1
XL2N2w4HtszrY6Tsn1T7zOMcyXvbnIbMQeQOHvQo+mmUHVQXw8ajVwSLPIzQgysI
uwT67q+hbR4EdnWNM4oPVT5Xlwh06xBUbm7Pesq/uhl8/EZQmywNT0cRVUNm+fjW
KfOKHc1vv54E5y2FiOR0fAcIvqY1KrB4w8dicMUHPNSXC8QjsQM9zT5/jmxS+XIu
MjIyn5PJR9WqZPJPiG39Mx3h2qAFHjUeAvVclv62VIPJSJZscFpfhmRE164C1jMK
IteV3AQLIMf0Fnldj51/RtP5XZdI4su7XwDH5zHJQSA=
`pragma protect end_protected

`endif

`endif   // GUARD CCI400_CHECKS_ENABLED
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
g1LAQRaov79lRFBvobPxz2N2Kd7jkuKqswC1fyDPEK2Z/hziQu9IXHGudhW4vPc9
10hCr0jsuHojH76j3HtQyRKYCfqrUBBPs64746qwx0OQBYyCIeB6oY28/2MRTMvX
R5FJNQpd/KZn9XddWtnHK1JnYho2z05K6Byp9Bm80+E=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 82438     )
adGygn8OVLdbR6cl6z1t5iC4BT7uZyfBJQcjwTz5i7V0OAsZNdEoM4vvXHZdaOth
Z325d6g+WmNYlLfZCS2bvjaB2lnAD/ewLYhtI1MjuIT2E+qtEnEOERgpJ+fSwm4D
`pragma protect end_protected
