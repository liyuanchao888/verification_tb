
`ifndef GUARD_SVT_AXI_COMMON_SV
`define GUARD_SVT_AXI_COMMON_SV

`include "svt_axi_defines.svi"
typedef class svt_axi_checker;
typedef class svt_axi_port_monitor;
`ifndef SVT_EXCLUDE_VCAP
typedef class svt_axi_fifo_rate_control;
`endif

 /** @cond PRIVATE */

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif

class svt_axi_common;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** Analysis port makes observed tranactions available to the user */
`ifdef SVT_UVM_TECHNOLOGY
  uvm_analysis_port#(svt_axi_transaction) item_started_port;
  uvm_analysis_port#(svt_axi_transaction) item_observed_port;
  uvm_analysis_port#(uvm_tlm_generic_payload) tlm_generic_payload_observed_port;
  uvm_analysis_port#(svt_axi_snoop_transaction) snoop_item_started_port;
  uvm_analysis_port#(svt_axi_snoop_transaction) snoop_item_observed_port;
  svt_event_pool event_pool;
`elsif SVT_OVM_TECHNOLOGY
  ovm_analysis_port#(svt_axi_transaction) item_started_port;
  ovm_analysis_port#(svt_axi_transaction) item_observed_port;
  ovm_analysis_port#(svt_axi_snoop_transaction) snoop_item_started_port;
  ovm_analysis_port#(svt_axi_snoop_transaction) snoop_item_observed_port;
  svt_event_pool event_pool;
`else
  vmm_tlm_analysis_port#(svt_axi_port_monitor, svt_axi_transaction) item_started_port;
  vmm_tlm_analysis_port#(svt_axi_port_monitor, svt_axi_transaction) item_observed_port;
  vmm_tlm_analysis_port#(svt_axi_port_monitor, svt_axi_snoop_transaction) snoop_item_started_port;
  vmm_tlm_analysis_port#(svt_axi_port_monitor, svt_axi_snoop_transaction) snoop_item_observed_port;
`endif

  /** Report/log object */
`ifdef SVT_UVM_TECHNOLOGY
  protected uvm_report_object reporter; 
`elsif SVT_OVM_TECHNOLOGY
  protected ovm_report_object reporter; 
`else
  protected vmm_log log;
`endif

 /** Handle to the checker class */
 svt_axi_checker axi_checker;

 /** Handle to the port monitor */
 svt_axi_port_monitor port_monitor;

`ifndef SVT_EXCLUDE_VCAP
 /** Handle to the FIFO rate control class for WRITE xacts */
 svt_axi_fifo_rate_control write_xact_fifo_rate_control;

 /** Handle to the FIFO rate control class for READ xacts*/
 svt_axi_fifo_rate_control read_xact_fifo_rate_control; 

 /** FIFO rate control configuration for READ xacts*/
 svt_fifo_rate_control_configuration read_xact_fifo_rate_control_config; 

 /** FIFO rate control configuration for WRITE xacts*/
 svt_fifo_rate_control_configuration write_xact_fifo_rate_control_config; 
 `endif

 /** Sticky flag that indicates whether the monitor has entred run phase */
 bit is_running = 0;

 /** Sticky flag that gets set when a reset is asserted */
 bit reset_flag = 0;

 /** Flags that is set when a 0->1 transition of reset is observed */
 bit reset_transition_observed = 0;

 /** Indicates if reset is in progress */
 bit is_reset = 1;

 /** Indicates if synchronized reset is in progress */
 bit is_reset_sync = 1;

 /** Sampled value of reset */
 logic observed_reset = 0;
 
 /** Variable that stores the exclusive write transaction count */
 int excl_access_cnt = 0;

 /** expected exclusive read response */
 svt_axi_transaction::resp_type_enum expected_excl_rresp[*];

 /** expected exclusive write response */
 svt_axi_transaction::resp_type_enum expected_excl_bresp[*];

 /** flag for received exclusive read transaction error */
 protected bit excl_read_error;

 /** flag for received exclusive read transaction error */
 protected bit excl_write_error;

`ifndef SVT_EXCLUDE_VCAP
  /** The current fill level of the READ FIFO */
  protected int global_read_fifo_curr_fill_level = 0;

  /** The current fill level of the WRITE FIFO */
  protected int global_write_fifo_curr_fill_level = 0;

  /** The total number of bytes of all active write transactions in the queue */
  protected int global_total_expected_write_fill_level = 0;

  /** The total number of bytes of all active read transactions in the queue */
  protected int global_total_expected_read_fill_level = 0;
`endif


 /** Internal queue to buffer the incomming exclusive read transactions */
 svt_axi_transaction exclusive_read_queue[$];

 /** Internal queue to buffer the current exclusive read due to reset of 
   * address by incoming exclusive read transactions */
 svt_axi_transaction exclusive_read_reset_queue[$];

 /** It sets ID to 1 if exclusive access at any monitored read location
   * is failed due to current normal write transaction to same address */
 protected bit excl_fail[bit[(`SVT_AXI_MAX_ADDR_WIDTH + `SVT_AXI_MAX_ID_WIDTH)-1 : 0]];

 /** * It sets ID to 1 when matching exclusive write transaction has been received */ 
 protected bit matching_excl_wr_id[*];

 /** Semaphore that controls access of exclusive_read_queue during read
  * operation. */
 protected semaphore exclusive_read_sema;

 /** Semaphore that controls access of exclusive_read_queue during write
  * operation. */
 protected semaphore exclusive_write_sema;
  
  
 /** Timer used to track exclusive write transaction followed by exclusive read */
 svt_timer excl_read_write_timer[*];

 /** Semaphore that controls access of perf_rec_queue during read and write
  * operation. */
 protected semaphore perf_rec_queue_sema;


 // ****************************************************************************
 // Protected Data Properties
 // ****************************************************************************
 /** 
   * Triggered when a reset is received 
   * If a reset in received, this event is triggered prior
   * to the is_sampled event to ensure that all threads are terminated 
   */
  protected event reset_received;
  
  /** Triggered when a new transaction is started */
  protected event new_transaction_started;
  
  /** Triggered when a new READ transaction is started */
  protected event new_read_transaction_started;
 
  /** Triggered when a new transaction is started */
  protected event new_write_transaction_started;
  
  /** Triggered when a READ element is deleted from active xact queue */
  protected event active_read_xact_queue_empty;
  /** Triggered when a WRITE element is deleted from active xact queue */
  protected event active_write_xact_queue_empty;

  /** port configuration */
  protected svt_axi_port_configuration cfg;

  /** clock period */ 
  protected real clock_period = -1;

  /** current cycle */
  protected longint curr_cycle = 0;

  /** current time */
  protected real curr_time;

  /** Async reset assertion time*/
   protected real reset_async_time;

  /** Stores the last sample time. Used for calculating clock period */
  protected real last_sample_time = -1;

  /** The cycle in which last arvalid was driven high*/
  protected int last_arvalid_cycle = 0;

  /** The cycle in which last arready was sampled high*/
  protected int last_arready_cycle = 0;

  /** The cycle in which last awvalid was driven high*/
  protected int last_awvalid_cycle = 0;

  /** The cycle in which last awready was sampled high*/
  protected int last_awready_cycle = 0;

  /** The cycle in which last wvalid was driven high*/
  protected int last_wvalid_cycle = 0;

  /** The cycle in which last wready was sampled high*/
  protected int last_wready_cycle = 0;

  /** The cycle in which last wlast, wvalid, wready was sampled high*/
  protected int last_wlast_wvalid_wready_cycle = 0;

  /** The cycle in which last rlast, rvalid, rready was sampled high*/
  protected int last_rlast_rvalid_rready_cycle = 0;

  /** The cycle in which last rvalid was sampled high*/
  protected int last_rvalid_cycle = 0;

  /** The cycle in which last rready was sampled high*/
  protected int last_rready_cycle = 0;

  /** The cycle in which last bvalid was sampled high*/
  protected int last_bvalid_cycle = 0;

  /** The cycle in which last bready was driven high*/
  protected int last_bready_cycle = 0;

  /** The cycle in which last acvalid was sampled high*/
  protected int last_acvalid_cycle = 0;

  /** The cycle in which last acready was driven high*/
  protected int last_acready_cycle = 0;

  /** The cycle in which last crvalid was sampled high*/
  protected int last_crvalid_cycle = 0;

  /** The cycle in which last crready was driven high*/
  protected int last_crready_cycle = 0;

  /** The cycle in which last cdvalid was sampled high*/
  protected int last_cdvalid_cycle = 0;

  /** The cycle in which last cdready was driven high*/
  protected int last_cdready_cycle = 0;

  /** The cycle in which last tvalid was sampled high*/
  protected int last_tvalid_cycle = 0;

  /** The cycle in which last tready was driven high*/
  protected int last_tready_cycle = 0;

  /** The cycle in which last arvalid was driven high - update is deferred by a clock*/
  protected int deferred_last_arvalid_cycle = 0;

  /** The cycle in which last arready was sampled high - update is deferred by a clock*/
  protected int deferred_last_arready_cycle = 0;

  /** The cycle in which last awvalid was driven high - update is deferred by a clock*/
  protected int deferred_last_awvalid_cycle = 0;

  /** The cycle in which last awready was sampled high - update is deferred by a clock*/
  protected int deferred_last_awready_cycle = 0;

  /** The cycle in which last wvalid was driven high - update is deferred by a clock*/
  protected int deferred_last_wvalid_cycle = 0;

  /** The cycle in which last wready was sampled high - update is deferred by a clock*/
  protected int deferred_last_wready_cycle = 0;

  /** The cycle in which last wlast, wvalid, and wready was sampled high - update is deferred by a clock*/
  protected int deferred_last_wlast_wvalid_wready_cycle = 0;

  /** The cycle in which last rlast, rvalid, and rready was sampled high - update is deferred by a clock*/
  protected int deferred_last_rlast_rvalid_rready_cycle = 0;

  /** The cycle in which last rvalid was sampled high - update is deferred by a clock*/ 
  protected int deferred_last_rvalid_cycle = 0;

  /** The cycle in which last rready was sampled high - update is deferred by a clock*/
  protected int deferred_last_rready_cycle = 0;

  /** The cycle in which last bvalid was sampled high - update is deferred by a clock*/
  protected int deferred_last_bvalid_cycle = 0;

  /** The cycle in which last bready was driven high - update is deferred by a clock*/
  protected int deferred_last_bready_cycle = 0;

  /** The cycle in which last acvalid was sampled high - update is deferred by a clock*/
  protected int deferred_last_acvalid_cycle = 0;

  /** The cycle in which last acready was driven high - update is deferred by a clock*/
  protected int deferred_last_acready_cycle = 0;

  /** The cycle in which last crvalid was sampled high - update is deferred by a clock*/
  protected int deferred_last_crvalid_cycle = 0;

  /** The cycle in which last crready was driven high - update is deferred by a clock*/
  protected int deferred_last_crready_cycle = 0;

  /** The cycle in which last cdvalid was sampled high - update is deferred by a clock*/
  protected int deferred_last_cdvalid_cycle = 0;

  /** The cycle in which last cdready was driven high - update is deferred by a clock*/
  protected int deferred_last_cdready_cycle = 0;

  /** The cycle in which last tvalid was driven high - update is deferred by a clock*/
  protected int deferred_last_tvalid_cycle = 0;

  /** The cycle in which last tready was sampled high - update is deferred by a clock*/
  protected int deferred_last_tready_cycle = 0;

  /**
    * The configuration that will be used for the current time interval
    */
  svt_axi_port_configuration curr_perf_config;

  /**
    * New configuration submitted by user which may have updated performance
    * constraints and which need to be used at the next time interval
    */
  svt_axi_port_configuration new_perf_config;
  
  /** Timer used for performance intervals */
  svt_timer perf_interval_timer;

  /** Timer to track periods of inactivity for READ on the interface */
  svt_timer perf_read_inactivity_timer;

  /** Timer to track periods of inactivity for WRITE on the interface */
  svt_timer perf_write_inactivity_timer;

  svt_amba_perf_rec_base  perf_rec_queue[$];

  bit stop_perf_timers = 0;

  svt_amba_perf_calc_base perf_max_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_min_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_max_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_min_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_max_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_min_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_max_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_min_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_max_write_throughput_calc;

  svt_amba_perf_calc_base perf_min_write_throughput_calc;

  svt_amba_perf_calc_base perf_max_read_throughput_calc;

  svt_amba_perf_calc_base perf_min_read_throughput_calc;

  svt_amba_perf_calc_base perf_max_write_bandwidth_calc;

  svt_amba_perf_calc_base perf_min_write_bandwidth_calc;

  svt_amba_perf_calc_base perf_max_read_bandwidth_calc;

  svt_amba_perf_calc_base perf_min_read_bandwidth_calc;

  //vcs_lic_vip_protect
    `protected
MSg5f>XeP_<OG\#bX]+U]RF1(=D@R_:\BXZRSc.3FRT4#VeVeb^?4(NXdMD[L:.9
)fFI,^GT#RA7OURBK8Jf]9G64Z;Q;PP;NeJKC\9&GXOVN5e[O].[@8SaAHW:&QM=
YPB_JB<3WYQd0+?^A;AG&dO+RG)@/de3:T#WA1_8bGYBQ+7CgGa([T((EU=\cURZ
WT9#F_&Yf0@;@a=LHX&T>6=_<3#E5;:[E8GDV8XfPbf_(LLE][O^ZK_HX3_XMIJ+
LBV:SGQ/1Q+#^=H]KWF1cOMSdc_f.0TF#T:Q1b]/+TYaY-bbH_=d?HGY@W(FGDb:
DQ#-NeL,<FL)ANY70c.Fa9_R5cQ>S,E<;_[=;)Y.8M7A/-3Qg@MVW6D24cD_RGMe
)MY28aZ8JZc<I7=MSTB5AL_R7$
`endprotected


 /** @cond PRIVATE */
 // ****************************************************************************
 // Local Data Properties
 // ****************************************************************************
 int report_new_clock_period = -1;
 /** VMM Notify Object passed from the driver */ 
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_notify notify;
`endif

  /** Variable that keeps count of number of DVM Syncs which are accepted and DVMCOMPLETEs
    * are yet to be added to the queue */
  int num_active_dvm_sync_xacts = 0;

    /**
    * Method that auto generates DVM complete transactions
    *
    * @ param snoop_xact Handle to the DVM SYNC transaction for which DVM complete must be generated
    * @ param phase UVM phase from which this task is called
    */
`ifdef SVT_VMM_TECHNOLOGY
  extern virtual task send_auto_gen_dvm_complete(svt_axi_master_snoop_transaction snoop_xact);
`else
  extern virtual task send_auto_gen_dvm_complete(svt_axi_master_snoop_transaction snoop_xact, svt_phase phase);
`endif

  /** Returns if all Snoop DVM COMPLETEs are received for coherent DVM Sync sent */
  extern virtual function bit is_dvm_snoop_sync_complete_done();

  /** Wait for conditions for DVM */
  extern virtual task check_and_wait_for_dvm_complete_conditions(svt_axi_transaction xact);



  /** @endcond */

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param reporter UVM report object used for messaging
   */
  extern function new (svt_axi_port_configuration cfg, uvm_report_object reporter);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param reporter OVM report object used for messaging
   */
  extern function new (svt_axi_port_configuration cfg, ovm_report_object reporter);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_axi_port_configuration cfg, svt_xactor xactor);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Samples the reset signal */
  extern virtual task sample_reset();

  /**Detects reset async */
   extern virtual task sample_reset_async();

  /**Performs checks related to reset and update variables*/
  extern virtual task process_initial_reset();

  /** Initializes master I/F output signals to 0 at 0 simulation time */
  extern virtual task async_init_signals();
  
  extern virtual task suspend_signal(string signal_name = "");
  
  extern virtual task resume_signal(string signal_name = "");

  /** Initializes master I/F output signals to 0 at 0 simulation time */
  extern virtual task default_signal_values_async_reset();
  
  /** Initializes master I/F output signals to 0 after waiting for a clock cycle delay */
  extern virtual task initialize_during_dynamic_reset();

  /** Initializes signals */
  extern virtual task initialize_signals();

  /**Aborts the transactions and writes to analysis port if reset is in progress. */
  extern virtual task process_reset_for_new_transaction(svt_axi_transaction xact);

  /** Sets the configuration */
  extern virtual function void set_cfg(svt_axi_port_configuration cfg);

  /** Waits for a any transaction to end. */
  extern virtual task wait_for_any_transaction_ended();

   /** Sets the clock period */
  extern function void set_clock_period();

   /** Returns clock period value*/
  extern virtual function real get_clock_period();

   /** Returns current clock cycle value*/
  extern virtual function longint get_current_clock_cycle();

   /** Returns current time measured as (current clock cycle * clock period) */
  extern virtual function real get_current_time();

  /** Creates timers used in the model */
  extern virtual function void create_timers();

  /**
   * Sets the delays in the transaction based on observed values.
   * Calls to this function must be made before "set_deferred_event_cycles" 
   * (which updates the "deferred_last_*" variables) is called to reflect the
   * corresponding values in "last_*" in variables of this cycle. 
   * In the case of bvalid_delay, bvalid can be sent before the address
   * is received or after the address is received. In either case, the 
   * burst_length information is required to calculate the bvalid_delay.
   * If bvalid is sent before the address, the call to this function to
   * update bvalid_delay must happen only when the address is received 
   * If bvalid is sent after the address, the call can be
   * made when bvalid is sampled (as in the case of other signals)
   */
  extern function void set_observed_transaction_delay(svt_axi_transaction xact, string delay_type);

  /**
    * Sets the "deferred_" variables to the values passed through this function.
    * The set_observed_transaction_delay function works based on the "deferred_"
    * values of event cycles. This function needs to be called after the 
    * set_observed_transaction_delay function is called, so that the current
    * cycle information is propogated to the corresponding "deferred_*" variables.
    */ 
  extern function void set_deferred_event_cycles();

  /** Checks if the handle given matches any of those of the active transactions. */
  extern virtual function void check_xact_handle(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

   /** Checks coherent transaction. If data is available in cache it is retreived */ 
  extern virtual task process_coherent_transaction(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Reserves an index in cache for allocation of this transaction */ 
  extern virtual task reserve_cache_allocation(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output `SVT_AXI_MASTER_TRANSACTION_TYPE lru_xact);

  /** Does the necessary processing to end a transaction */
  extern virtual task end_transaction(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, bit is_removed=0);

  /** 
    * Updates the cache based on snoop response assigned by user after 
    * receiving a snoop transaction from the input channel 
    */
  extern virtual task post_snoop_cache_update(svt_axi_master_snoop_transaction snoop_xact);

  /** Waits for post_snoop_cache_update() method to complete if any activity
    * is observed on the SNOOP channel */
  extern virtual task is_post_snoop_cache_update_done(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, bit check_outstanding_queue= 0);

  /** Adds a new snoop transaction to the queue */
  extern virtual task add_to_master_snoop_active(svt_axi_master_snoop_transaction xact);

  /** Adds a new snoop transaction to the queue */
  extern virtual task add_to_ic_snoop_active(svt_axi_ic_snoop_transaction xact);

  /** Drives the awakeup signal during idle time period of addr channel */
  extern virtual task toggle_awakeup_signals_during_idle_channel( );
  
  /** Drives the acwakeup signal during idle time period of addr channel */
  extern virtual task toggle_acwakeup_signals_during_idle_snoop_channel( );
  /** 
    * Adds the transaction to the internal queue. 
    * Blocks when the  number of outstanding transactions is
    * the configured max. value.
    */
  extern virtual task add_to_master_active(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
    * Notifies the slave that a new transaction is received from input port.
    */
  extern virtual task notify_slave_new_xact_received_from_input_port(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** 
    * Waits for a new snoop transaction. The monitor uses this task to get a 
    * handle to the new snoop transaction.
    */ 
  extern virtual task wait_for_acvalid(output svt_axi_master_snoop_transaction xact);

  /*
   * Returns the number of outstanding transactions
   */
  extern virtual function int get_number_of_outstanding_master_transactions(bit silent = 1, output `SVT_AXI_MASTER_TRANSACTION_TYPE actvQ[$]);

  /** Returns the number of outstanding transactions. */
  extern virtual function int get_number_of_outstanding_slave_transactions(bit silent = 1, output `SVT_AXI_SLAVE_TRANSACTION_TYPE actvQ[$]);

  /** Returns the number of auto-generated transactions. */
  extern virtual function int get_number_auto_generated_xacts();

  /** Returns the number of dropped coherent transactions. */
  extern virtual function int get_number_dropped_coherent_xacts();

  /** Advances clock by #num_clocks */
  extern virtual task advance_clock(int num_clocks);

  /** Steps one clock*/
  extern virtual task step_monitor_clock();

  /** Waits until a valid or handshake takes place on any channel*/
  extern virtual task wait_for_bus_activity();

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_arvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_awvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_first_data_before_addr_wvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Returns when specific events are detected pertaining to transaction processing */
  extern virtual task wait_for_slave_tvalid(output `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Drive the idle values after initial reset */
  extern virtual task drive_idle_val_initial_reset();

  /** 
    * Adds the transaction to the active queue. 
    * Blocks when the  number of outstanding transactions is
    * the configured max. value.
    */
  extern virtual task load_active_from_master_buffer ();

  /** 
    * Adds the transaction to read_xact_buffer or write_xact_buffer 
    * depending on whether its a read or write transaction. 
    */
  extern virtual task add_to_master_buffer(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);
  /** Detects initial reset */
  extern virtual function void detect_initial_reset();

  // -----------------------------------------------------------------------------
  //                                EXCLUSIVE PROCESSING BEGIN
  // -----------------------------------------------------------------------------
  /** It returns 1 if there are pending exclusive read transactions in
   * exclusive_read_queue for which matching exclusive write has not come
   * */
  extern virtual function bit pending_exclusive_access_transactions();

  /** It checks the transaction with the same ID stored in the queue */
  extern virtual function void check_exclusive_sameid(svt_axi_transaction xact);

    /** Pushes the transaction into exclusive read queue after all the data beats
    * of exclusive read transaction is received
    */
  extern virtual function void push_exclusive_read_transactions(svt_axi_transaction xact, string kind="");
 
 /**  Removes  the transaction from exclusive read queue if any of the data beats recieves a erroneous response
    * of exclusive read transaction is received
    */
  extern virtual function void remove_exclusive_read_transactions(svt_axi_transaction xact);

  /** function that compares the expected and configured RRESP for exclusive
   * read transactions */
  extern virtual function void perform_exclusive_read_resp_checks(svt_axi_transaction excl_resp_xact);

  /** It returns 1 if transaction with AWID = ARID exist in the exclusive_read_queue queue */
  extern virtual function bit get_exclusive_read_index(input logic [`SVT_AXI_MAX_ID_WIDTH - 1 : 0] awid, 
                                                       logic [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,
                                                       output int ex_rd_idx);
  

  /** It monitors memory location for exclusive access */
  extern virtual function void check_exclusive_memory(svt_axi_transaction current_xact);
  
  /** It monitors the response for exclusive write transaction */
  //extern virtual function void process_exclusive_write_response(svt_axi_transaction excl_resp_xact, input bit excl_write_error);
  extern virtual function void process_exclusive_write_response(svt_axi_transaction excl_resp_xact, input bit excl_write_error, string kind="");
  // -----------------------------------------------------------------------------


  extern virtual task wait_for_cache_update_post_curr_snoop(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output bit is_snoop_to_same_cache_line);

  extern virtual task add_to_master_current_queue(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual function bit add_xact_with_same_id_to_queue(`SVT_AXI_MASTER_TRANSACTION_TYPE xact,output bit[`SVT_AXI_MAX_ID_WIDTH-1:0]  unused_ids_by_active_master_transaction);

  extern virtual task update_current_snoop_xact_handle(svt_axi_master_snoop_transaction snoop_xact);

  /**
    * Creates the transaction inactivity timer
    */
  extern virtual function svt_timer create_xact_inactivity_timer();


  /** Tracks transaction inactivity */
  extern virtual task track_transaction_inactivity_timeout(svt_axi_transaction xact);

  /** Waits until the transaction ends */
  extern virtual task wait_for_transaction_ended(svt_axi_transaction xact);

  /**
    * Tracks suspended snoop xacts and triggers events when they are ready
    * to be added to the queue
    */
  extern virtual task track_suspended_snoop_xacts();

  /** Updates response parameters when supplied through delayed response port */
  extern virtual task update_delayed_response_parameters(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** returns a single unique number from xact ID and ADDRESS */
  extern function bit[(`SVT_AXI_MAX_ADDR_WIDTH + `SVT_AXI_MAX_ID_WIDTH)-1 : 0] get_uniq_num_from_id_addr(svt_axi_transaction xact);

  /* returns address part of the unique address-id combinatorial number */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH -1 : 0] get_addr_from_num(bit[(`SVT_AXI_MAX_ADDR_WIDTH + `SVT_AXI_MAX_ID_WIDTH)-1 : 0] num);

  /* returns id part of the unique address-id combinatorial number */
  extern function bit[`SVT_AXI_MAX_ID_WIDTH-1 : 0] get_id_from_num(bit[(`SVT_AXI_MAX_ADDR_WIDTH + `SVT_AXI_MAX_ID_WIDTH)-1 : 0] num);

  //-------------------------------------------------------------------
  //                       PERFORMANCE ANALYSIS
  //------------------------------------------------------------------
  /** Main task that tracks performance parameters */
  extern task track_performance_parameters();

  /** updates the READ inactivity time performance parameters */
  extern task track_inactivity_time_for_reads(int perf_rec_index);

  /** updates the WRITE inactivity time performance parameters */
  extern task  track_inactivity_time_for_writes(int perf_rec_index);
  
  /** Updates performance parameters when a transaction ends */
  extern function void update_xact_performance_parameters(svt_axi_transaction xact);

  /** Updates performance configuration parameters based on a new configuration*/
  extern function void update_performance_config_parameters();

  /** Collects performance statistics when an interval ends */
  extern function void collect_perf_stats();

  /** Creates all the performance classes used for calculation of each metric */
  extern function void create_perf_calc_base(svt_axi_port_configuration cfg);

  /** Gets the performance report as a string */
  extern function string get_performance_report();

  /**
   * When invoked, indicates if the performance monitoring is in progress or not.
   * - This is applicable only when the svt_axi_port_configuration::perf_recording_interval is set to -1.
   * - Returns 1 if performance monitoring is in progress when this method is invoked
   * - Returns 0 if performance monitoring is not in progress when this method is invoked
   * .
   */
  extern function bit is_performance_monitoring_in_progress();

  /** Reports end-of-simulation summary report, checks etc */
  extern virtual function void report();

  /** format report string */
  extern function string format_report_str(string exp_str, real exp_val, string act_str, real act_val, string unit_str);

  /** Gets summary report based on values in perf_rec */
  extern function string get_summary_report(svt_amba_perf_rec_base perf_rec);

  /** Stops all performance monitoring and kills the thread that is tracking performance */
  extern function void stop_performance_monitoring();

  /**
   * When invoked, performance monitoring will be stopped if already the monitoring is in progress.
   * - This is applicable only when the svt_axi_port_configuration::perf_recording_interval is set to -1.
   * - Returns 1 if performance monitoring is stopped as a result of this method invocation
   * - Returns 0 if performance monitoring is not stopped as a result of this method invocation
   * - If the performance monitoring is in progress, that is is_performance_monitoring_in_progress() returns 1,
   *   but the axi_port_perf_stop_performance_monitoring() is not invoked, the port monitor invokes stop_performance_monitoring
   *   method during extract phase.
   * .
   */
  extern function bit axi_port_perf_stop_performance_monitoring();

`ifdef SVT_AMBA_ENABLE_C_BASED_MEM
  /** Converts an AXI transaction to memory transaction */
  extern function bit convert_axi_to_mem_transaction(svt_axi_transaction xact, int mem_data_width, bit convert_read_data, output svt_mem_transaction mem_xact[$]);

  /** Populates data in memory transaction into the given AXI transaction */
  extern function bit populate_mem_data_to_axi_xact(svt_mem_transaction mem_xact[$], int mem_data_width, svt_axi_transaction xact);
`endif  

  /** Enables/disables performance monitoring of each metric based on configuration*/
  extern function void check_performance_monitors(svt_axi_port_configuration cfg);

  /** Enables/disables of all performance monitors based on the argument */
  extern function void set_performance_monitoring(bit enable_monitoring = 1);

`ifdef SVT_UVM_TECHNOLOGY
  extern task write_to_tlm_generic_payload_analysis_port(svt_axi_transaction xact);
`endif

  `ifdef SVT_AXI_QVN_ENABLE
  extern virtual task qvn_process_token_request();
  `endif

  /** Tracks the timeout for the signal argument provided with its timeout value given
    * w.r.t to the event or status provided in the argument list. 
    * Mode will be changed to enum type as seperate activity. 
    */
  extern task track_timeout(svt_axi_transaction xact, 
                            longint timeout_val,
                            string timer_name, 
                            int mode, 
                            bit status_equal,
                            svt_axi_transaction::status_enum sts_val,
                            event timeout_event,
                            string port_mon_name=""
                           );

  /** Tracks the snoop channel timeout for the signal argument provided with its timeout value given
    * w.r.t to the event or status provided in the argument list 
    * Mode will be changed to enum type as seperate activity. 
    */
  extern task track_snoop_timeout(svt_axi_snoop_transaction xact, 
                            longint timeout_val,
                            string timer_name, 
                            int mode, 
                            bit status_equal,
                            svt_axi_transaction::status_enum sts_val,
                            event timeout_event,
                            string port_mon_name=""
                           );			   

  /** pushes an exernal coherent transaction into port monitor */
  extern virtual task push_external_coherent_xact(svt_axi_transaction xact);
  /** pushes an exernal snoop transaction into port monitor */
  extern virtual task push_external_snoop_xact(svt_axi_snoop_transaction xact);

  /** 
  * Returns the number of READ transcations that have started  and in 
  * active queue
  */
  extern virtual function int get_num_started_read_xacts();
  /** 
  * Returns the number of WRITE transcations that have started  and in 
  * active queue
  */
  extern virtual function int get_num_started_write_xacts();

  /**
    * This method is used to get list of all IDs which are currently under use by outstanding transactions. However, user
    * can choose the type of outstanding transactions this method should consider while extracting ID of active transactions.
    * "mode" and "rw_type" arguments should be used for this purpose.
    *
    * It returns '1' if total number of unique IDs currently used by active transactions, is less than all possible ID that can
    * be used by an AXI transaction. This helps in determining whether randomizing ID field of a new transaction which should
    * not be part of the all the IDs currently in use, is possible or not.
    * 
    * @param mode Type of outstanding transactions this method should consider while extracting ID of active transactions.
    *             Currently it supports following modes (defined as string) ::
    *               - "non_dvm_non_barrier" => all transactions which are neither DVM nor Barrier  (default)
    *               - "non_dvm"             => all transactions which are not DVM 
    *               - "non_barrier"         => all transactions which are not Barrier 
    *               - "dvm"                 => all transactions which are of DVM type 
    *               - "barrier"             => all transactions which are of Barrier type
    *               - "dvm_barrier"         => all transactions which are either DVM or Barrier type
    *               - Note: if "rw_type" is set to '0' then only read channel transactions will be considered for non-dvm
    *                       and non-barrier type
    *               .
    * 
    * @param rw_type Indicates which channel id width should be considered.
    *               - ' 0 ' => only read channel id width and transactions should be used
    *               - ' 1 ' => only write channel id width and transactions should be used
    *               - '-1 ' => common or either of read or write channel id width and transactions are used
    *               .
    * 
    * @param use_min_width If set to '1', minimum of read and write channel id width should be used otherwise maximum.
    *               This is applicable only if "rw_type == -1" i.e. no particular channel id width is specified.
    * 
    * @param silent Suppresses debug messages from this method if set to '1'
    */
  extern virtual function bit get_ids_used_by_active_master_transactions(output bit[`SVT_AXI_MAX_ID_WIDTH-1:0] id_list[$], input string mode="non_dvm_non_barrier", input int rw_type=-1, input bit use_min_width=1, input bit silent=1);

 /**
   * Method that randomizes DVM complete transaction
   *
   * @return A handle to the randomized DVM complete transaction 
   */
  extern virtual function `SVT_AXI_MASTER_TRANSACTION_TYPE randomize_dvm_complete_xact();
  extern virtual function bit is_in_reset();
  extern virtual task         wait_for_sampled();

  /** Checks if a WU/WLU transaction is received from the sequencer while
    * there is activity on the snoop channel. This is checked only when
    * snoop_response_data_transfer_mode is set to SNOOP_RESP_DATA_TRANSFER_USING_WB_WC
    * Needs to be done so that the WL/WLU does not get ahead of an
    * auto-generated WRITEBACK/WRITECLEAN
    */
  extern virtual function bit is_wu_wlu_during_snoop_addr_activity(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /**
    * Waits for WRITEBACK/WRITECLEAN generated for snoops to be added
    * to queue. Applicable only when snoop_response_data_transfer_mode
    * is set to SNOOP_RESP_DATA_TRANSFER_USING_WB_WC
    */
  extern virtual task wait_for_pending_wb_wc_for_snoop();

  /** Gets the time at which an address was invalidated due to a MAKEINVALID coherent transaction */
  extern virtual function real get_makeinvalid_invalidate_time(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);
  /** waits for transaction which has been blocked by other transactions more than `SVT_AXI_NUM_BLOCKED_XACTS_ALLOWED number of times.
    * It wait for those blocked transaction to finish. This will avoid starvation of some type of transactions and will provide
    * more fair chance to all the transactions to proceed
    */
  extern virtual task wait_for_severly_blocked_transactions_to_make_progress(`SVT_AXI_MASTER_TRANSACTION_TYPE xact=null);

  /** waits until VIP is out of reset */
  extern virtual task wait_for_out_of_reset(int mode = 0);

  /** waits until VIP is in reset */
  extern virtual task wait_for_reset(int mode = 0);

  /** Wait for start event for performance monitoring */
  extern task wait_for_performance_monitoring_start_event();

  /** Wait for stop event for performance monitoring */
  extern task wait_for_performance_monitoring_stop_event();

 /** Perform master signal valid checks during reset*/
  extern virtual function void perform_master_signal_valid_checks_during_reset (
                                                                          logic  observed_awvalid,
                                                                          logic  observed_arvalid,
                                                                          logic  observed_wvalid);

/** Perform slave signal valid checks during reset*/
  extern virtual function void perform_slave_signal_valid_checks_during_reset (
                                                                          logic  observed_rvalid,
                                                                          logic  observed_bvalid);

endclass
  /** @endcond */

//----------------------------------------------------------------------------

`protected
5RC:@V_+3d/W[7d])BM@7Qc^ec(R1[S9XJ8US<IYPL1fgF3-PBdP,)I@>ZbdZ2J#
M7GX,f-2HPg)Q0FMR]H->Z\\P5gD>^<[c#X]SY3FJf0?Z^22[d8Igg-DIWd&FCRR
eE6]8]Y=RV_;ZKWMbdagJENHcY+YL@a2?Y/,Q[gUM(3V-JB:_8VDY.D)SdBO=EXX
<1d)/0JQM+BH>(2S4/(3XG29O5ZbaU?TOCe[?Z>b8QKPM.6Z<^WFQXCF[g0Og&>A
Y3#6Rb)-^eTA.c4B=_?2^:W:-&D&JPHW4-]1)5T32g-+E&^.-)<H@VJF@72).1;E
WT)aABN_9E[faWe0B.4=7@\ac#@U+0ecga/6^[Wc]F>g>cUALFK:H+NWYNERO-8d
(^&eV?0X8U.:3;M3W?4Zf>64S;1L\eR@7/PPTSHED:/V:SXS<GC\(0AOP75[\acg
[6H<4Y9:):T>KS/0#T;5SOC@#+A(@B@.V?TVF+Q-KccMQ4T9^AVW:B?#0_=YgU&L
SC/:UXEF5TVTaFG2@L)B4D6:HW,E>XTJ[7gS-A/D4Hg?/EY_7=Z>/[?6c-cg7]F9
d),E8\I6F,?WEZf8Da6:>YO.::D,ONH)[b(\H?30GXHLgF]R8BLO&;KD>7(XEd.8
PR_69UZNf(WaH20;eDVGE5ID(7AF:XG;>+2fZ3YI3>WGc[2gC>EB^=.FJKX)1E5A
]GSgO09+U#f;=-(/:+7e_CbPKcX-R39WH&O@KHfdb(/dD]Mc/\N_a5Q#W4MMd567
WO:&,C#1?I]E\Q;aLfb5Ke0CHD@I2O^Z/f7.+^R./gK+U[Q#@0eOGa,\OM0f@J2@
8Icf:#fSU/AU<?)R7;,^^F@IU0FbU_NN;/VI)H/^d4:b&T:-+(g>5?T]9-6g9J9B
1+a3?J=U[^)e.O9YI8SG_2c[c-7E?5)]5ZH.JSUeJc:+<>^Je]YD<U+cW.#f<_RD
2W<-+aRLVdg@@U70L+8)\d.EJC.afK#JSETgX4eEe#?c-25D,HeXS<V&@OE:X8-4
:LB]5TF5@.U5+KV4\[C&-2#40E4Q8988CQb_cfA:8]0)R?HS)LE=SMX)1f4BS6<L
RSARWY0gPcGD+&H./a1HL-6([2V;Uf1A(WE-(0Y2,VDR#L6;b9PIXcC<.X^]<)gb
BY0@BX0<+/)#;-gG1A)8gg9\IW.KgW]D=.R^M=JLD=B63]64@UXITc0D:.F0)^WW
9PD:+_K:&I5LWC:OJO_)6J^@(:Oa:PO+T&f0+L8-DZWFLcNXIdIKZ08Q0<NSa/Ic
OT-=\fa2&gO/181d2/X?B08.87dDMLI8fOcdI?J;YV7J>&,#Q5;c,:Eb,,@_VIgd
JQU(I,F@af4cRJ0)1f,2)UG<E-EIdBE]Pc^G&)>?-U&FNCKEMX3G)g?D2-B>D/Q-
A14-9HL\14PG3C#;(.K54b7NJ=e9KHTcMR/<0:#@+6?+:\8#BV,Z<KG;cC^BYA4Q
OM+>DB&0fcX.E=OW<CTVK^(1DXADR_4eZTQF/O>O_Xg3&)5T4+=^FJH?=8D]GeWU
80EZ.@H/J\g11\dU9\B5=HG5Q84O1S<X(P:[GeNcU/_&^:,Nb>88_;;D?<U6+gA.
XXKV#KH5X:.cV&cA8BZRAcIRA;C@UfaGHQNb3@Ug>JN.[,eS,9,[_.H-,>a6\5AH
3?4VXe\>XS-BcJA5)[3P]B?X4[^(YKf=aMER5.,XR[E,d=11Q-_9PZ:5E66Wc[2M
3+=J7A<e.0V-E7PQDe6;\PaYcVDc5;EAM[0-+c)gID)W;8LQLQV\11UFYD[bNRb@
f-aH,Veg1=.A;&/8+\TOZI=(Ef2I-b4-3-(=F._+4K4@>4NL/9M@]9^MMcbC;;Vb
&0KJcGEQESJIf;:M0NH]=d&KS^B>VeJ.)&6dE]EX>,Y,+2M(3JW0d>KL,8&c/ZDD
)eNaQ28^D=W3eXML=@[I#M:0eQdd81-BgC&DLfCA0-6#Te.>?L:TEB<P>,H1f1D<
TARc<CD)BS3L&</CZeH?9OVe]c2Y]H#T2cG,QFAPPeT5:BBI^6>QKJ5@ZGNJGEOB
C>L><;^]<U<JN4]9[EP6T?Y^7(D@dA?DJOaR]<1)S9G(#f/eeK0Q:[X\^#&&PZ\+
,.44U)@b1(FbA5f2>.>aK4+.c@?1c<R/eN@7IfWOg2N52@R;BL6Uccb[NdEf;17#
:G5I^L[CE_SQW0++8DNcF/Q\@-[S2ac7]PTaG0/:B?L6K^X<6Pgc[(U-<^Y6JaeE
A+;_)NL>MXIH&A_UDUVV(XcPGX+>a:S.B2_:DZ]HG:/IG9gW802DINB;C2C3RJXg
1)0KTdB]XB_XdW1cB470[9Wc6-&W\GE#7:HFY_gLFbVcG+QVOVH_7WXZN(ST82E(
gSJ.0@X:N-6ME_e/f91SU>RZ(DKXL&Z_,df(c-HB^dH&KA7P-PWZJ]Ca0;^+]P=f
M)Yb&e_@^.^)B6(<@a44BO.EI.H3]3@FJ[]A5H#@+2HZ7VR(7YQ#))>.RU=UeeMZ
H-ZeJ47<CgfNK<:56=?FS)?#Q-7@HW/4bf30[)UU0]H<O,:=/bAQG:V^V9@&\6L1
4aL,Uf-^V)\[QYDOXR@HXAI&N/E109g;&7PJ?G;N-NEe]XD5T=QH)B#\TI3=ISNP
]HWEA#Va,)+D\dCZ[faFJbHUB9W.DOD6Eg9E[]9QM_>2:R5b:2Ye>/+?AF6?RGR)
dT:Qf2,dF3D7b3e?f6;-4+bH_T0g>a5b:T\)4B.+ID&g?+3R_UQ(eSa:^a\/@)J/
3Tg/[,#OWF2@X6RH[7O=UfO:_79TJB4H2@bcN)+HW(Q/X[?<=6MdY#R;db>+fdFN
7aVd;@3;+>(E)OY&aXc,C#UF0OeJ8WZU1#L\+e-L)4FbcXM5RA-&&<g>++#H<XA#
0^Qa(M8-(W@3OM/L?KRTBN<Le5P?/Yd.CI=H\?T7\IPc#=WZ[<7F+\.W+=NV@59C
\K:4K6=LW/,]RQdAA\=9UD=0O4W3>\b.U_Z<Pc9G@IX#H=?2=@^GB3ZgV83.&1Z,
DWAe4IG>f8GdcI4XMd@SXE6a_Ra(cXBI[WR60XfdJNTeTcU3E9KL)b\ZOKYNZ(S?
<G?CH1f=[)Z+I=EZXKV4?L=b239;GPe,,DI_TPZdDg/]D3eOH)eNM)4C0--gIG\<
+bMYH0+K#OBECbgRbZ0S<JDeVAR>+PPL.T=S9(CGUOMEC=IBX_CR7W2M,<2Y8J3=
;fBI-0S\/^5e37,Q7IBJRR0/g>Y-,58K(JA^4EL&N0Pg23CY&M5P8aQT@<.V&,Rg
(_-\=65X36/;f563bdFd.@-^?bH43Wd]Z;RgU\W6+0&cXPc<3P=2V+5;EGgS[GGC
KgT8#?c#28b;M79T9d>Da8N8RGOK]gKN3]LVVRX]TTGBN5<:#Z5BHPT)\COCBD\A
I?A6d,#WBGd?#bQT.N[]Bf&O,6D_G\#\F@dcIJX-N:?R:VbHT\<^3>GeW6_@--^#
>U=V&R1;U?Q&\HQccbbI4K?b@XLGZ@Gc>,2)bK;8]_J+9<5cT?:T[9WPZEV\4Y47
H6cCLU>D(eMeF-IB6?g)B=UNX&Y2X<,SOcdC=(e9S,@RQ0D\C_;L8HbaSU)U[WM4
.ZM\[6R,[)C>+^F4C+Zd>>@fUb1\CIf?P6UJ/;bDaaPGgdcJ1C_cZ7\Q,AOc_,Re
IdCO],[-1VP7BHQB#B+Eed-7aIJICaC_/C93>@aI2NZ#aVD2F1AFS(:^CgO2CfWH
\G/HY+2-bd.?2(EH-,VVZE\CQ_;3AePLRa@9YO92Q;.>A9J=LcXDQ:<Y0W]dFT]b
(dUSBg?d:^R0]D5b(O:f>Xf7&=OMU-M+7RM-F,<)<2Ed1BB>Oea:KY[:.7Gf#aPW
>^K1J(bBS8cS>WXT?:0+[3[VC=8b9]0@2HZ(-eFe4M=@_H^36V\3(R.9e9G[O47R
1V9beV+cEYIG7N^KO5b8]_VN#@L;d&]ZL4-5gW)7bUNJ<5VQLY1?Qg?S[2WBLI74
&U&TTRU/1.>4bc9LbM1eLI/VX^U5AS6(R2&XJ7N-P:#CGK0P<eUHKM_8F:Da>]Y0
?=#F.cX&fBf=?A7#:9CX0gfScWf^FIU+KV??,H45aPNMeVJQ)4]^d.2Ua5aa_T57
@3,,\5J/3W8=3e4+Zd>R=/>0LBE-b^UX&(7J&0-GW2BYf;#bK]>_S;PC\fO2A2PX
_#;e+S=,PR[A<AO5Q(,BO&IFf8E[ADGIA.Q8IA\9ee[cTEO1;_,&PfYC_&?139JC
\0_ZE&:J[67S8^+gT;HGGg)>e6;6e+3CDADe.PON#c9_FZ?903>GaZ&N8DUd[dQ[
GH2V;,2QG+7[\?Bc<HW55e&>1SIEHV(3WPT<GVTX_K<7Wf6<eM:H]IN4QK=T^^a=
>P@)O2Xge01b[P^V43K)P3a=I<U(615YY5XVERV<BRZ,[^,KR45R9a_<O98Q,0IA
a>Oe,JZGP#[KBMOY\>Ef@G+LE..75:TEYGJ:e/GaGL>C,?[5SfG(E-KbLTJ&#f<3
HKKd;HK]Z+P:c4LN(=5E37Q5E^f4O9M:NA&C/Gb>=eZYZF&Mf5a;LWdZUeAR;IX7
6C2e3>I\=#9IW5d/0>)Kd<:e-1G\Zc)GJK/Wbg^SYfUHRgWF@10C\;dZM$
`endprotected


//vcs_lic_vip_protect
  `protected
FUMa,Eb((HUZ7O-;W@Q68LacOg.4TC)U([[OeWd1&PKM?bK.c,;^&(0RB.H;1=+4
((U@X65bK+,SHIRJ_591+>2(Ed5a6-@dXLOa/aBgI-J[]LC(5TC>_[)NJ->bBJd<
[+\gD@.I]#@XeEJL8QbN=d70?>N#=6X)9<56c<QV#e\e1N>1\IX=]=/2V^Y]GC>e
1Id9\G]YX?U,N8PNHN[93:G6+dB43/aWJ+<f,M/TR>]_5&e&#9\^#2;=]WQ(L)BQ
BU0?<?][)d3IZM0\Ya\?,d[Y.8FO=aG52J.942+T)WX.;bI1EF#F[KSRA=:b,W-S
ecG2QeB4U<abY&J9COf;(T5;X]Q>><3FE?Ec:D_+\WXZBfCg(T&RXTYg6D?SOH:F
S?B;NbJ<[C\;L]dc(TS/[I(53a^MS2UBdZ.DY6@6TBPSC>&)UNE]URHb.FY_/,0,
:^+S5f4eTfBO6,(YaC)A;N:P(9_5N6(H6TEe#T0]A.,&7I3M_,(aeQ8Z\_5#H+PJ
X[[9+8&5XB;Z)D6XEVbC^5;8]_cV=+1UB.KQd#HcXA12JDceINNXMK4\@GM;BH^Y
.+]UN1E:)(fb<EbRSK4+(4Y:S]5VFe?QX(#J>>ZHE-U3RDNV&SL3E.T4X->QA9@U
+G>f/WgA8.H<[T(@)bRe?PXPEP2,HIZIb5Paa8A8dQB89SIPbeWJ0>KfM)b=,5+&
A+EP&,)JB3T,ZfT[[JU_H8Q>_)\>d@K6-GLe]ba\)RA=:aR^@EE1W@VIYW34_>2/
G.f+^N;:=&fI95WNZ>g7DC&J1/YK@3NV0DOGVEZ62T.O?BEd4O86H>dFfbE\:W94
,63>J)6=J(X-f#)06Y.5J^8[.UR@3P^bNFNK::,ZfCMXbC[D_DUWVHT<U:H1^@f=
N^^/-6=;8B?ZN_&9[_L5/09L^DfK/,XO&4QI3db?SLMZ^KEEbb+DI)G&gV9Y>T+5
A/G-&J9c+M(?W8T3D<dG(.G\QJ>)0@DbG>&B;/We&V&-a?/P)e_UT##<(e83[P9=
#e_)<Y#1>E(8-69M:U?/V/#\dUC5NY3#BgU6N(#>=Dc;@]B\KFEFT)Df8G/Z>P>L
d#Fg1L[I,R2YCU4SYdB4JT#6F9-_DO7]VTcd\IS?9R;,[^M#66PM88RR9f-.DZIU
bA5IV_U9@;232<Y.f=7ZeCD[O+g4b.FeJL?4N5e32^OCM19,H0ER3\_WFSA;&3N^
;QPa:[KE:A08.TNLE_>^PSXYFb.PI7a5_4UH7.D(Y1W#TC6Vf_]Sd@Lc;U,GIW5]
N4a2#^cQbd/R]?KL\:[0@T,/P<FY/]JUR)PGc9<cH_WMZ2@M?-7#C(,1bJM^GdI:
667BbB?TZ;)D^CCUK<N\C,QBQO_IB(,aM/(S6<+/A+KY\PUf&+Z<@#FcF.MJG@TU
cAWEdWE#WR+O\>6KZYO4YVIS[_BX38LC<.N^NP?3U1#2RX8+(HdVAEBI&S1g\g:1
&4_8f]-b/31V:LKF/KP=aJQB3?TP,<6_-=HNK\:KWLaC_d#D?C=NfN4Y4d>^a7E^
)Pb]ZabLc7&OTJX&J.ZUU[OEP#6#=S(.F&UCB^d:e)UA2J::Xa=)[+]=M>](-,SC
A;2HJa[e)@W^L>/KVOcSGQD7ARfF9IDZK;4NP^c7H<+&1FgT/_9)Z37@+]d]655f
,Wc;DSICaBJFb:<036dF:GDUb=24#+4a54]8.+g5=S>.0F<4E=1J\dHCNAZ0g0Xa
5ebNFX9.2+I]CMcJ)P#87UEU?@9b1:U>e_WBa&.B59OVaHRb^12T:9,c###TJPFM
#gaFKDJE^7b;A8E34(A^D[H-Eb^H\E:6\^^X9-55(QLWQ6RQY(>?HL;JWbKTD\53
f8QXVS60KEZA+:+CQ6Q,@V1Ua7MC8LJ[6YHAbe5DCH@2N2]JIbDBV-#]:1\U2IGD
I]5FSb[@V&HC(QO:;fQ+-R-?F>RQ[GD>#\+dF-Q],4bA]#VTQ=fa.WJW=7Vf.D7D
-)S>;MI<PL\))D7f^)ST>W5(Q2HePMAc([X-Y^-/IAM9#UP8:FH#-3PSS^I2G30N
1#S6.R,eL:&.P/?->9/Z[5YaC:N#CZ_QS=>)8564LO?N[dT4,KO+]<I-W&\WBD]D
b]1BV0Z54@0@2,5=;(QM_)2QB2b_9HPC1E;BQ^X]YH[:8eZ@Ab<6G_M>]?>[#/@]
0:+I0d@QA+)\LHbAV_MVF.=X==W;6f;TKIecAB--RK(;#dA2@GgH9/15[dD=9L_:
P#;RS6a;FcCEMd[0LNdQdEWFdbeb6<(aFe\(Z#C2E#4-.b53[]ACf4]>R[_E2Pe;
=9&ZD+HEVbZQZPU():3_Z^/1D8dcK13eY<KU+RA.J/3:9a9LJFG<#B=KQV7/:+@L
Yb5ON,?[HG++\YMCXE+=M-Q\:3^+AETF3@/+2C,;:KI>SLSWJA4S)7//NH1)@^8e
dFf0&I32[?X+AB-CEG?9B[Z3UJ1>,X0O,=gE)PFGe7(:.:bR(U,4QQe.52Z&^(JW
WXU=?.dLSgP9J(cL/I.bF[4A]P\^J7fQT+,aQW04I06&[N&R+1-7bYe&&g/)1IYT
BdePV0U4P(R<+&4W7aJ;KF#U)?EG0A/</3&80NK7(8\KWUUF-accb-\AHcX#-,,4
HePaCW>C67KYfC8]4)G;-]KQW4-L;G\6M@]9_[A_/Bb.K-4[/U(3XBYeKO\]RgZS
,H=TA/Qb<ZLNSS93HegbV9_&)MdV1^:9H_>N;13gR6G3M,,EOURPDg4=AR0b0?b2
I,@:_=dWSGVRZ<c@?8BU4)D0LJQ#JX3U1BI<?(3Vcg?,,SFSeVf^_-#8+T:=,\PC
e]#?7&O,Z2;ZWVaQIa4J8d:0I(de)[13\B<-+9B?O7eRC)=6gZ#+O2ZRU8DT;IH:
^bC[X(NK16M8N89BF;0_1#ZF/WU^fH\K.V-Q48WMQ6\NTL:HEZO3O2U/7./09f<b
\H:2>#W_#W2b]GUaSY7:&-F4Q<V0Lc/JGVF1YA;a\@W/,#Mf^#_?F?6JAMaF-fT2
dWG0FL2X3Tb(Xc;E9e]WVQbaTQ8<aS,AU]-8)?)bM@D3R,HEX44&9ZAVNJaJ/E\-
A5Se^7MRO/e.b6f\;I146)ZTBbZ,[-dGNQP8K5Da<83/;?La72[N7TLf)&0.We9H
AR:.]&b0/^f=/]>OYH&O^O:&=C&U0D<Z\C.c6AU]Z(3O/?Q@2=2>D22/31I=;X6I
11)TL>AMH+bN<2YQ-Jcc0BJg(J+YVd5WW1.e[T84.4c[6IBR?4+2S0.1ce+;@d7f
=UCI<E)HG>6\Ce-PR7:6Y1UE:aGE;#P/J6#OWbP?L?P/+:@X1C3?Sc/PK<EI:;VP
ZYX2,dUG-9,\cYOVc@MV5/4Me>V&8).J?A&8(T-^3d.&/a^G-7gU+:-<R7/aO4.Z
,U[Q[>bE5#1&/=HU3.dQ5(Q4N;BXHX3/P+PF&6:bA0>;6_KYV1^T_8WN2Q6Y0&#&
D7K)DbKHg2.YXV;AXGF<b:g7-1B:f=JO(E4[[R]EFe[-4)05OZ.RIf\>4;g^:+>F
:9Dfcg2VHLOOc/(S/a^G6-U#DAeGd9W>1OR^gDg-\#6Z;[>[f?[UFHGbU&MI72P[
R3&A2BW=QC\f99SC+aE5Z97>d[eB1g.&SC1e:EJ72?WJ0HYVBN<dY8J_JWI<ANO2
KZa1KF)<aJ;>Q:J11R<fYVOA)R??0Y[N_0GH3:?Re>M>YGV?##cUMKRc_/3=,P[R
;:d\LG&U,LC<_SOQH3N#B;FQDDW:I#KU_W7#4B+SM5&56#H/?V2XK7P:2B.(=Te;
0PbgN4.1SNZb;=.S9ab4_4R+HQM;G]/41Xdb?FC_4R[6HTa@)LB=FgHUA+6,QCH3
DXOL=VR[(,[7V>9gWVGAW.;[U7;Ob6Y5VREH+f(/B8(3_0-FABg7WB6f=cJDW(B.
:<R<5&cPW_9=OQbVO-8AL-\RHaVQXFKJ(832/\A:SJUNAK>cD;2.K@M@-B-W>gZ4
VFg+F\0RX,5ePFS=&.4;&4_3Z&J8ZFF#)L6/eR8Ng;9_N2W3WCO1aPXbTBHE?\>P
CR&MVP\cY6WZa6NN.ATRf/.OQ1:4RXM=OLT],R<Ng1HWJD+^X,_LI+d666#>C)NY
-b4RTSEL9,NZ(:6-BX6K75(()_=6dY0/YVK_b.3<61Q<OLJ0cJ=1O&,YDAKUUUK^
NZC21(F#V@::F2E>&Ec(LX#]O=/=<(K47SDH1b[ZT.1b7/A^d0,;SK8EJ8#2Q(<N
&DJJdW6K\E_\9&b([4Xf.D/X1&C_G.LHZddc8]T5;^#Y7N)DG^EC\-L8/4@?31NO
T@9b7?f:-eSc&VgT]\P^#f)-LDY:geE)X[EP/F+2LWIdPKT1T=@eI),g]^YZ#)ZH
_ZT^+0HT=LY8aLHD-Q7[O72J-Q;RR381[U7?N8begM+D:B]Y+O6YF&_F9&a(>HN5
6VadQMJda[FQc<H)^L[97ZEAeaJ1,,^3,YUgK:<GdT-ag]T)W)6[=SSfXb2\B+Yg
G&4V9L8&YVONN[:@Xf=OV3EQN)O@E)+UY<5@0?5^;T[P#;6-c[(#M6DD=&I5L<VW
2XIZZB])?KUM<KZVN?2&77fSAd(Zg6XOegK<V7ZKgC]ZE\aY[DA&1JAIaN<>>GKP
SE];#HTLG5768<9))_V:#I5c25B=:)DTHELABWL1Rg3U(beU&VN102>YK=9^<UM@
+6VN76U:+IWY4aa=&1e#[)X1daGR7O0OP/1AH]aPI,SN_Q\/GGQg#&Q(G,YYf8-g
-HUK/232=(_7=Ng1f#EW5JIbB&bBFa&+,CD46)GJdL+6,6:S]]YS>UZLa=?0X..#
6HA/9,LZd?TABC:gV.YdKQ#]_,:[\g+X2)^;8_gXI>e&,gc&\L4fS]9FfS&KEHRK
=+CAEfe&9CcR,7LFD1QT-H7>/P\L]Sc-8.aGG-bLH6_7TeSA7L4)>O:aAG+;O:VG
RZd=,\JRdf)ZJ9N_eC=3VgSFL40>MID]1#_Lf0L<^Q0MT_b2a7./FTc#;YXXZ&2S
eCUZbaM;JR1]/&eg#/MaQ=Jb=5YHY,6\?DUMIDC8aW8e&JEC7HPHH5[(\a)K]JH5
_?RRA)<_C>gO:c5XX:ZYH>V[G-\HLe?5[&L1\\Z-5,NY/DPX0FHac_4Q6]49<9FA
SXD7CA,9gR?6+eNC#<d)D5E8,?II]bBI^BOd>2I4&dZ+bbK3WaXJF(d:2YUc+?H?
3bbW2BSFeXWN:1FfCc_?N)\S^bV=SA[20Z&FI93M-6)FQgNW)MV.N:RPUZXQFYJf
;QL13T];1_^CY3KUa03A#0:NVb[=A5cSePeVa>f070a6QZUK-ge2_cZU/OWVW&cT
YN)?Ab>(P_8H;\a(^ETG4P]KM:(1(05<dd6=eTb7P=Q7P+VXWBN=P&@DQcae^U,4
40cJP1;]?<e=<Rb5:+U45>3VB<bfU#fKZD,M1QP<+N@UX-)=)P&FMD&X/V2CUT[Q
I9)T,.SQ0]K#]]+@3CBV)E\2^29?EDDV7IQ60Q^M=OSNNKC54\Q7HY_.D&R-ZD\P
N7^.CUIgeXfQa/>\@LC3.MdWS5/0\=#<N,OQ)T7S2(a7eO_H[E\T?2JC3TRUZCXM
ZXU@=K:,;Y+5+#@ZgAK?[[3fdZ);]L@bF)C0EQ)5LM8W5=[5QC=^TN]Jg5X]1N5-
Q)-/PF[8D]ZU^8>=D0]KGEZW^4Rf2#^.>KYS-XA^(fVR5cfHPS/;PV)F4B:L_;96
N<6??DI96H#Q9543C.g/VPYffXO;&F36eEK->Y?RWeNJg@GJF\=.EE+_;01IS=g[
,&HL9:eLKS2YK(b-YYXI,EZb:1g:.8MGSbGV#g7DB>TI6^D[C-K[#d9G^)L^;@G^
A;J(<b,eD3AbQbEE,c@#I7+)E<UQECT)5?[f[b?7TT26^1@&+[a>I?R=]C9@YaNX
HFJKPeQ])a5TQP.[&Id&&0,beFLE4_acP+N,CgJHM?^GK5Q83H2W:J(^69J+ROD1
PNFB)Tb7bf2Z_3Z3JJ+0He?V&AEK\>IWLLG27KUF\\>H[UWG>Q\FZ.=1/AUWCT68
]DO&fN;-PIC(E5;/GX)5T4_\:+)ZIXOFO;ePAae@#9HWI3XdQN.,U:d0Z^<7U=9;
(6Pf?1\ZT814ZJG=F4#RMR[P+g0);3^[..Ye4IZSG5=S=2Ve:NfC>>(aAbb?/f_=
Sg)8VKVb3CSV3@S;f/=36JGVBFKHQ3DM>TV7TeZ_R,C.2SP5/8=\dXd/c(OQH-fb
D,?EROg:gf6WWe9>IYX67O-C7;LVGH4&b&&J\-ZH7_JG(@1=BgTd,(:[f3cD-77U
cdc&B9PePW2:4#Y?8:&V<(UFS4::P<]7/=&Cb;RWB?]7K\&=NDa<5c_)\/3G/;JD
/f80<O#_USYOdS+].#9@eDPc@gK__XV>:0faL_2)W3CB@McX6a<N-P:5ZNFG^0W1
0BL4e;G<_Z0Kdb?^SeV_ecH4LY0_UNGA&Tda##.ZG:?C199:Z4668;e\ICB2eJ.#
[@VT@2ef-C/BX]OG2B)M[O9aN<L3HF8Q^)a&b#;[[Bd>WbA7Q.OeEHM83f3#\c99
O,4SXWMWT-GN)KfYX/aI9TO_=>H3__NRWXHeNTRWC=3fM4>Q&b5@^X);+<QRD1.8
_V@#;7=g^6]HB_XXgTLfc83_CXRL7Z[/0+\>G5]D8T1UD^ef?\]#;aZ>)R)K4AAd
&[\dK0+(/RaWBMdZ+Eb+AJ#2?Ng-XU\L:aFKV[>/NNf/0c.2Db8f::FDPNc/bT>U
B0f[<&c)#;LBOH_:[6H78^^E_)19?GCc)Y2LRf8OSS1B]JF));;ZBVN6JH[2EA0J
K.HDV2DNX+8WUQS,V.VOfUb#M93>=WG(JMS&\(^Gg&PW>G6AY-fd.QUggg^d+#I-
M-=JR=P[e_ZLWScJL.WL(_1&WDXXZO-dL]IY]>HeU0K4+1Qc8SQY\5D&Sg[?26C3
^.D(Q&PH-_dCe0[GDR\@PB@SbADK<\6-ag)K7T;OND^ZB;5<.AU@=WNdRV(N58>4
08B#AVZ9d^VZBLB[bO\PKR;C4g#A+98J9EJ0Oc=H@Db4GZB)]5<:5:?Y@\Jd)09?
F3gD0ceTLe)57bTAg#658WI&PX/L0#I4FND9>/_7(M<5?Z(NJV29+QK,MXX9.&_-
P,PTJ_1<]^_@b6ec^DES@]CUOOI;HE4<7QK/7.-(WAM4[9MaYK;9@J:G9?R4\__U
Z]ZFQcT?43f#OOFb6A66bQdF1J0?XGbcBZf<5)3=KSg]HAQ\\A9(F?M])aZYG<gg
_AZLS@dRCAFWZNV+LX\;Z?C[TM8K8M?eIPQ:99@&^)N&2(JRP(KCJ4_+Ae>cJXJ8
fFC^.77;LS1E6P1A-3MOM:fdIGB/DbJFSg5Xa4B,0e#X2[>;F628e>-@)>(?:5:W
2DgE&[6A(33,FF^g#:@I_V8/IY_^D8TXYa#JTQZH8OQ(20[)@;d&.MdMFc/Q.bTK
QUEf/6+P7I7?-H8BRR(0F\a3KBZ(Gf.<a#PJGc8:.X&E(UZ2\V9(WZ:Q)_cK:7@C
M_^OIB)DM[FfAJL.CIOH6\T6<\&E?H#O)?:9)89W>eLP#<2@>35G2bBNMKTO<MQW
,97W/gK=.f(Ef=JO+fGJ+Y4c\;AV@+(HO0)&+Q=O9&AQE\U,,4>(1cgLcSZ.WZ24
)3G99=ZM/EXXcC7g&[52A>fV)Y_BA>F<M9244+IaF=OZGHdd<TKC1-e;@8Z3^T26
?8\X1ARI7+4>I_a<a#(0,H5-F=5aG;D0Te4/Z_M\Ob,eA-NGNYVGf;I)L.e8=,)M
81g[9M?0.C9/g?>O0VHS4f0,65g@Nb/FH@P\5PS+f2e89a/cfA2T:,eZ:UfQYIR9
=J/gWI8.:#Eb2bJR2Uc\.cOEA5L_&LND?_:D>P\dUYe:b\ZZ/eJT7eDa/E#R#+;M
O:V^cL_fAe;AbG4_T\MC)R-CI[PE+EWS(E.d>fEU<V9c^HQ9;U:&NbUK&FI/P5)g
1&bHTf;,N3GadG,0\170F&]>d1HdC27QO^]SFMPU#2fcO;:=/[^fK<W.=\0OKUDV
gP+e<c2e;MV-[)6-#VDS]G+16#dG?BDO)T.>Y]<7N7/D3/dF,:+\L<EG)9Q]W\+Y
P[.8-fW-/?P5=/<f3QIc155WMAWSIHYVP7dCAK,IBL&OMMI(]P&7;f>;g4OSP/>>
_7dR]Oc6H\e[3\+1H)3,d8D5[#c5/L^<8]]2=(P[[3N,KI7[U+eR<M]H<.McWTWI
#:,/GPOR/G]6RP?K-X<ST&CHM&O_,.I.7db1/[S-d\>++R\7CO?D5F4bc[UZ;e@T
[_bVXJEKOB84G0MdIb7;M:d2>b;<EgF:JXW)X_98V^4K7KIII<f;_D8#HWC;)WR&
f\e8?.#C1]#6_N=JT9)8_QaTH[Q?g=A17R,6G8=FOF2?d;6^KS?R/N15M&H.-H<Q
;7Rf)3RAfUY)I@#<J_W7YXLDJ]RR><:I-ZEC^:6>RBCHFPe+DK-B1b=\H.WG0XY#
,2[+<)5#:<&dT,?Q#2Y\>Q9;(U93a\KM\@SCGJ/DIP3<,4Bf2We<DWZ6Y22FV_5\
YdGgK>;CSLHf<;1:39eS177gIQ69C-TMH(K#UJ&OO[WS@3)KP<;T./.KB.XeJaeF
?W&&Jd=[-fS#E8ODQ]5KGTDf=g/=B7a9?+?HZH\<XSA9MGVIeVB9/O2<2]K3NTL?
gZEC>Kb;.KW;;F8Q#&PG)T4g47#(8;>+/?aQ^PSgf+:K?/R<>D63cZ#IO2N=5.-L
;5fE2UL9^DNd_PIK#?O:&O^eBbFML/T1SHa8dC1bG2V>VG]XZCIC6KN;>VbQ,?OC
9BZ&\gY/90W0,9?[?;>6S<G9Mg=^^JNF[XbGe(6,:6GYJg,;+=15&DfA-Q1W(Q2c
4:NM\b_0Z]>..4LE2@gXR+./=YPNV^&,]3).E+J==B/0:dOO<_L.CdB<4Wa;SBUd
^Yaa&^WKZ=0:;9Q1S).3]GOYcGA&I.P#3.>K1#AbbSa]gD[C@1,=G[(geBd>)_[L
8^W4)JTY/V+1/M1?NN23TU+7F(PA[:?4D5A]9#]6[J/./Y4AMeB@<:K^M_S?\PBG
K>2(=TLLTG0DVX58?7Pb.S_2M_&GBR&b&EJ<C)A6(c.fAe#K8XV>K#cHD@[ASe,M
.[9AY1U:(d=C<Hf/f.(0Q]U7]2IGHY@f?7NT<e5S6K9Y##WD_)bHa5Ca(DaU7e8Z
AcS9]7F)4@eVe=^37BBARH5)8Y3^>bB>G?0XTI6>M,dd>(;Y6dTSO7UT3>&/e&QX
V_GOJFgEb^(]@Fbc.PU+SMWFe8a(7;AFNe98\a)F;8HDHGc@]&\8W5_MV-^d/:XW
Sda0g<1a@\AQS)\BWLaB)0_?^(H0-<&;XZG9OcgRVbg]>>RB8D6(^A^OdF8cYc?b
8g\@3)4(:WG:9;4_0Q@IL&NQ-HU0<FK#:JJMJ:Gb=>a7OZ+Y],dHfbWF68<M=40c
:#&49N4>U:,:H9V?gg2RAXDS-6XZS/@CW0O+:T[LVF5UYeQ8<=2\L883,>4/10]B
<Y[I4SI(RRG(9b&[;,Q0K60dEV7?=Q)3L7UE<2Y1H@Y:3G<abA.M\>ZWe-<]>7_1
Yd[.9&(dGQNOF[E;8W(;a<F^/YIT]LBHAQ\3@>SCCgL(1-S\U6[[1Zc0c&Uc-cDZ
0_)a^S)ga;4AGJ3?f07P4?M/]U\Q_R87YgM2M.=M&H:(7-4J=gBa7+e&5Pb_f2?7
@HDYUeUggNBKF6cbRK&9/+)DSK=P:8,HdQT,9J155_cYCT.IXDfCCG;_8<F:g#\+
DG2ZI+S3/D7V+#X>>O7.&feS2f\:^/g#VSI4Q0dA)c)N6U0\XC0+R<=Tgb2PYY#I
+&QUQ-D3^\#(AC5b68K.FYS_Dag4V.M2E>Q@OI>X#Z=)<+a]TTbVDU5S^2\fVK/0
??a,]agUGFV9JV-F9RQEaN3_,T?b?fOc(?<:3X74E7(.4_5^8]2G^gX2JS6(/WK5
C(K[K:dfK#=>?B:NTge.Sd=E0[W#2P\P#bb:\+IR28X.PT9)Ofdac<P6-Q81#^CI
QWf/d1X3J0;IS/-)#;aPPG:@JVcbC-HPDWL^C)eL9ff2NP]?B:DC;WYMB,N/X+P:
>J9B5QX)N0KgB>TN^2V@e0YY8H8S2H2g:9EV@ZPeX..bAIS8f15F&Y)<VB0Q58A?
G]H^(,>PNX50H5P6@>]FY[20^eI#L;C4Ed#-I6^VOH^b5<@B.VOZbA0&]5gPFLg>
K#Oa0.f#ZKPUUc+f[7VR1(5g)11EfJN.][a+UY2>M4&g,R6LK+4K_-V^<SDGAQ9b
3bd]118^M7TPa(<COf#8P&C2C<d@V5R;4:#9=#^1:4I<Z6LV>C-G4)RYVSC-<bGC
B?.S9SET\W.V2e#D27c\8##@0&]ED02T,>1O#?D9afK,dLZ;R.G0]+C(dILNGX&.
&SCbJ0VI/Lc.b;.CcZ^SM=dfdf3Tbd;-(ea<:5Z2E20F^9,N=2-3\./cW,cQ>32Q
/]1A(;g^3KXN;d8D43[4g_c&R<ZRT]HX0+X/S8UFUM29V&G>\6?5]bS?(UHNW:]f
2OGga-Z_FdH7#,[CSBC+DKc-5NF2RRfZ,U_;<d>WK<H)#6JfYNZ7UbEbaTSX?)&G
_;K[NGeH;B2PFQ[O6=9?S/RLE-J3LgPc70]&,P-)KgIRZ4aJ67H\AX/.[+:bF+9W
GD[?Y#&c6g:ed8&(1dd)QSZP6K_:;VbaG5I(:3PV<D86PN?gT,_9)46WN#.#L:&Q
##-VOZW@RVb@9V=I]J_aVE4,Y?]Q/-F544UTL9N-SGG_I0J8WOL(,_,JCB5IYMaB
f:[T?KW]Q^(7A46^LR+>W2FCFK4MO6B;I:X2^+-&Z[C/K@5fGE\D;Y_B/^[bI#[V
A3HCH^]=5XTcB3[6KA[_@dS)49K:)9KZCO3g.e?@]T5^7BdY[c^b.-S<M\:.0L4C
48QC]\6U#V?GM^dg\+LR=L3VedL^&g]2H,9--U7DP40d9/]g4=<T&&FIL[0>5c&/
_DR7V0^U8]bNU/M0[]2D-@3V5$
`endprotected

`protected
PU1?.f6]2BA-\Ug&H^NfLD-M88..T]#6XFfUFZ9W&f+-<R)P@(75/)XEHMN+?K)/
IEN-+B+6F1--,$
`endprotected

//vcs_lic_vip_protect
  `protected
f@DJI-=8(#3+a.><?^;[@OIV6])WN;NFAX3,dYV-Sab?I?BO<P,W,(J</J@N0=f0
g0JQFc?aZ]CRT.T/[B;/4GD:)SN[d1LWV0H]C2R,GH=.e6_a[,-^0(,^AC6WJ=];
V:??]1Va4,^PB9X/_6F+\(0UJ4dfJ9dO@ZKI#FXd9S_@E45\CYbFf,b(;(_5dR9I
#&ZQD_98I-=1JG/HU=_+#Z24ccbT.&0;&/.#cV6?S\=)W;)YOEL)FZETLY^,7f#c
1Q=DL0C7g:ZP:OWQP13g.+-+YFK,9>,F2aL?(:2@H_>cP6@(>0#)GK74R8e=1H7/
<-1@M[I5^C)#beOQJ:<6)?cD+MRC>)TUcCg/OZ#=B4Xf+5R<LFUe\:_S95;-H<cg
V07HTION/J??#E08Cg<c)N6S)YG=cP8[_<YLEA7?SIJ37Agf7Y/0#;4<>[5T\TX)
WOL.(]@YGIBXLg(V?H(BUJ)(UUC1ddIDQd3):F00ELCEK-Z>IMQV]Xe,e,ORQM;0
,\1eI1AGTHI]c4W(KX&4@\.6/0TD<IQ-U-:QQG8KTX:deFKK<b0J>5d?OEUJC_5Z
:RO#d7UM6;5)4R:#+UST,2KFDfF_XCGGH3:.FSIL:<4JN_H5[:;bPU3P&W]4@a\#
Qf:gC&K;RSLTb,BWSEYcebF)N//=44SY>8B==97;1Ab@b^DO?aD]_PLd+9:g;J]=
4D/=XN^QF)7cNN=6+DgVUdOSa(02ba1P+M8X-(N:UO6HeP6&+/-+C0?C_ZG54.UL
V:2Xg557NNL0VT-fTS@A_ZAEdKaF&-STZ1.)59LC&L0Qg&6/+;gAa50YfTe0<K/L
Y[.d1=BPaRc\.<8&9I;\B7KNb9bI\Y?IU8Ra>b/DLb2@@;)D>=5XYDID[[47>CX7
e&Pg;J7>D+G+_gd)LD4+?M1[9B28/QQYD[61QI6Me==<g#LQND?\.UaSRfd).8VS
@KV]UaI.&U/27ZC.CP^8.7GDN5Xd=MbLCag6;,[?80M6T:9+RORKMN#\fA4ZPS+A
1VJdP@=)U/Oeddf;OMbD/@>fdNM=1L2A]:FI_OTFBD]20TOMO-UcN2D0S^69+]GO
#UP[;,KSU3^^7TI15#)B8c;>5+F6I\<^#\ge8Z/f.dZYHF1fMUfeDNF)HMbI(\DJ
,<JI^(5=?_Ae+\aSM\NQ0+5eNQ>c<0(V\WN/ZHME78@2/RQfGce/Z?A+#-R7\>V?
OZ^6Y8/RW^Ic.WJd7\PP9MI4)G+6DV5aSGR0H_76V=?C:[9H14YLDF:=/;I+)VN)
ZQI9;YG243/>H0;dg/16EDKB[?W-2N(B+9e<3I9>+,B0Bc4R04416:(NG;X4#NM[
dg(I\+9e:5/U)HgLKF:E5P9XS_]+&eDL9MBKT7YPUN.AHEE52:/_\0>HPfTJg+Za
XH<)C18\T?e>F]HBe)PefJB,.GLS2+)9@E4-Ha4NE3/U8-G00)e@f)Q4AS?GUe&?
,QYD0<^?/JBa)ZeKcaD_,__[)S+95ZU\G<)eH99EXa\.MS_G&XE083(CTbC]551A
N8@5UaV=2/5.YIG?W([T3L[KJ]D7KHZ6>d5]LK:DWTFB^<-EY>LHF\YI[)<2,AP.
G&1<8>Z#JV8aPY)(IP]2VcH<18OOR8.J@<9d.gL,]<\3bO5)#Dc;(AJP01<>Zb&[
ZZf&ca+cXD0OV2KOT9.9\3H&:,\.QB^?B/Q3L/ea[>U,REH<QH^Na.P)EYY6^&\#
)C?[A\S/DY4;B(:&^(9E.LXD];9^Ia[Pb[0KO2Q,H0TYT9+7HJWZB+AfG^M],8SQ
e+\Xc:3\Z92UT910A@+:,AQ]U_\M3K76F5ONPWBL6K>;#K43MY5[cGJJaT-1-1FD
18NNXZB))VTg1Ed--D@c,T8A[V0?WOZLNOa5E,YQ6?[BK<&6B62Y&QJ<gDMH=@@X
9A[NYL>Xg,X@^&=]>^/QBLX7.5Xf807)FLX1+/]Va[CFb#E?LL]#IXc9g6?KHM<b
52V6,5QSc6X4N\HP:^a/Cd+6^@TG<^655)L,J&&MeM.agU&7UOTJ2IDI>K1/JW<?
A#QX;F7ZTU]&FLVHAa[/P[FJM<@O,YF<Ad)WGXG18cUdgQ@5IOIaWFQXG]HDR^aS
g.F\dXfc@Va8R8+b/YE[gZQ>X,P4M@FQ^XccZ)X]5TZ]ZBE6WO?:U-OaaNR:?-bY
4KCS6XOFB7@X\:1A-26&Q9]Mg^^T;d/S32d5M8cGc4@Z,PMGSF<U?WP5b8]b=^;<
;e<-TN]_AgBNe()N0Pc_CeI\H.(36S8Eb[LBPYY[1S[OIU]3We1-BLObPOGF6=XZ
ZML9:6:&a.WPB#,QC8[;.N(9L6gZ.BgB6TSf=F:0C)1F.>T&c?8BA;OBB-T6(OES
G,0fO,D4\P_K<IB5)cP/+ETH+HSgR#NZ+@BC6O1[)51@d+IKAZ/8J7S4+?b,7,+P
PI51d9+;&(BAdH1aPF\.+b43M700f=WM]3[eSEC;VD@E[UTGe\R^=/ZT7MZQ?M10
4/7-;;#QSIM:)CI=KACb.=KbS3T6<cg++a]5CA3SNEJ&5<3ED#DKf.5,B,\=U,W#
B/>E97c_8edB;C3gTe]GfX)+2+28g19U4cUb.f(FB<Q=@]:63FaNd_bGbJ.RHT&0
D8??9#<MK82N=NRaY1U0-V+1:QZXO7ZI-GUg,Z)75(LUM@2cgMW_U1[3Y4La;.BQ
HJUg:N(TJ9U#A@?:>_7VINdTI<@EY#6085NSCBQ-EA+8<LPI?;UdA/(/V7dOIQQb
\O>QIE-=CDd6B,NPEDN0eX[^de]Ib+1b0=b08J8JFeaLKK^0+ZSGGB8J602S2OQE
YBB7>4U=PDX&@Z.SB9J4G>E(8X59LcQTU(HJHE?S^J@==/]:aDWabFaY@<R<NZ)<
/#8.2f]LgX1agE:;ZBCQJ5)bMAT/MVF&;4H&D\HHe+OWa[.?>NCAI=X42=O/(fDU
N777><8f8caW[7e<FJ_VIb_UZe4>M\@.Q^;YR6<T?9W:ZPO1JL[gMQ70R>eU_UB_
X_#=I5_NgM]6>6FZDW2aB3FFAAX[(7@;[_4:5.dE6Hea<T1]607)SG75JL=FH(g=
S\V7/]96)>X->>b)FZY5.]-ZL]T)@66]/YSI]NKbFAC0D6PWQIR1T3_aUVCa#0_a
dBS@YFCP^W[=b_XcZc&RVUFIC+8a<F>?F4-d#<P.:CD,Eg@W(3DR24=T?S(D6[WV
\:SP<WLZFgE]30:(D7#JNPWRb+a^8C6N5cc05HQBU)3R?OcGZ]C[IfO3J:4gXENL
ZBB3O#ELbAF&[(W9I@K=V<UbgTBZ8CR_OTc/NcaX8XLB);RQ/O,M/)16JX8g0TR^
dNXF#P>(QB7Y7+#M\DTZZ=6CI:dTV>g))WZ964dN\a]P32UMVXf9H[M3(C.3[Y[>
-Qa9AB9N6P=6g//161&YTL&^:B3a[NJAb4C/1N3\]FLW3>c,Ve;-e8_^[,KW++AO
S()PR5PQTIV_YAL?ZU1fcH\<5?DRA[ZM;:DH=#<fYHY;H>G84UAJMNMTDV1>J#-I
Q9C)5#K4?H<Q(cLB<&/:FWc=aeI;[+H@XbW8<gP:JO+I+;NAfcJ+S2KWdSR#OQB&
e,<S;:2>FWd0Na(?Fd)I>F&FgYI[E@P0\BbRENCCQ-@[FL?3B5CVIIb3Z_a9dMb9
-R2X^T1e&YU5ZDBQH;^CXZgN]T]gGgZ])Q+7I8aX/&]F7A_\D08>.B)6OTcOgVR?
EY#c[A-fLOY3GcI-[U1H@6PL#4>OdNFF;_,4SFd/0f]2@FT1BcR>1Z.f\N8/ZHW1
_cf2f[?1(0fGB#3V&.J]GI?OFZY5/4^K:;Q]\64SfVUL]37g:=4MI++F_+#(X.F+
ML[?E(UER@?BZ#>?b\9=Pea+Yg^>a>K3QQ?1\:G#T<^NRgW7A1fB]#f2]bY+.SFI
\L9A)&D/WU-7-=dcV/DU56A^RfJ].f2D<VK&1_TG&JW^HT\-a6EHG;[d;_R2E00N
)J9WG/2XgPeI6Yd.75)#W,40D^4,R[W^;XPL/4ZIZ6?QZ^?#L(F,3]KJZ/;:KY,f
bNN@WT&=Cb2H7PZ.#[YNNcgFbZ=J#A[;L:A:KN&ET+<:YSbSI#6[AE5VZeZ9\_Q:
,2\2]M9W1-=LNG_Q1\g#HZ141Bbd?+1\E<=#L?S_#O4+:5b(E[[&+0F9KRU^7)Q^
KFa0#2BV,^:LZ9>@d80G4E-5cQ_P8S4+X^,ONR2I4/3AEO22RQ?HJ:2FS85T=SXc
>6VRW=]]KP=A3&f1N=Y-^&\\K-?,a<Oc7A4V.PQ4AR;(BF<RJ?14V>NOgMa44/;[
BNA\1SZ(dS(<;.O#UfG&D7+d5F:JAT9\f0XY?X+-[R/>L<8-[#fQ.)>(Db(P/&7C
d7>eCUKBY2gdOWHEd\-&-6aObX7Ve][61(@PH)#AMKc^N=FcEBG\[SHe71M5W@(;
\L(_9Y14B0U::#R6V\#>-3=56V5]b/M9_GWB0&K(5,g)3F#He13D^)b&2XJ]DHH&
0F40+8)]2,X>?f^N.&/I;C>]D.G\2B8G4,CeK4]HcNRI0Gf]R??gX\L,N:e77G5<
UE^F.=b@?\1M1&(]/&]Bd+/MZCE/<Q>ONO>YB>G_@&QgLWGF.,@VT=D0U(SX#:H@
0(3]P.g=1SHTg^_2UbWM;:8@ON1?/4Ec8OHT1bg&;TD@QTM;B7V<N\8J4E/CA561
V4Yc5M3.V>JST(F\=@OUcC,^++baV(Q-],6VJN<2[^fc?g5UH=M617#(5&a316=g
>?IS7T.Kc^XBPWVDc7U:aUe;#]^,4V>Oe)JY@Y7&V3&9Sc1aU&&Z6Mf.7WPPKa;R
eUdQc<LPQ#J2>a/b8#e&A(L6+?W2W:2SN:6Z]8-7MWe8?9Nf]6)PgMea?c4MKKGE
::5])+3_(La+HP?bXGZSTbANMV<[N85_V#X4D3]OFLU;eO.De.OfX8G>8+1Sdd25
fW(6c:?cFO]F&:AHIGf5ZYQb8e0J=-gZ0fd>I5F6;aVYSXYea1P79N42H.+(_EAU
3DN3U0EV6@)MANK,DH(?HV++N5bP]/8K#fHUNYXLK6T(c94).T@DS?BBPBKe4bNJ
QK^(:DFQ=OeIa#@8f2#T=-CC+B=FTc@eU9]::A^C<Y@5.\Ugb[T_b#K[Fa-:0?Y/
]+RJ_=_^;Zc;UO;QK<V5@4gcXF=cGTIS&9ZN/5DT.@K)b25.HWNFL8^O,CDQCJbA
C<9>TN=P<I>J,[M<:EHPS[4>T.DPce=;<XX&T_L?-Qc4JMP=D^-LMebOX4CG9=-@
]_N0@.g^#VcaX6+b33&2RZWTEGWaU7EO/9ABE3?58;4QM?,UOJ:=DN;_UR&_a,;U
L\(5gP2_d=)(-A<0dWeMYaAVLMREB-+INV\)bC>6Kc=&>:(S,;RL<E?)L#,L>7A;
P=\8:/WDDOXYIA<I=01)-6E0XGLZ..c=9-f:W)g&2c--#U.Dg3?\:W1QbV+:ALA0
\D8(ODJ:I1FUe?D?N_d,d<(L)&U934_E9dT:K65O-TZ6US2EXO2M)CcPQUI\SH/1
V/&N623Na15U[&W(GOaZ9D0@SaL6./ES:#9&(ac=]fN+91a./EHaX>f,e[8[7ATH
1E78,)1TGUYXW2T3[RZ#=E\RV/24KE1R6^5.8:UcJA&\Bc16Oe#[Q.RB8R+_85.d
ORUVf.9[@4&;<>(RECS>:_&:SUP)Q?aU-V?TTA#H2(F-9PdG#-G_#L4TDW8>K)P8
e#/XV0S+P0^_3W(gKS;=f5V[:G-IZYC47_gD-.RdX/?cH:9V[<O=K#;T=7UH^,FM
fBV7@22]_8(NJMDDWXH^F(4Yg9DOW]e[c]U68.,3#b6e.F<M1L81?R\1^bDD#Ua(
WCE@9.I^7IK\/=ZP^/b;6^NE4b36QZ-Jg:6?Kf>d[#Oc\T\KHQ=#[TJP53/gR/Vc
JJUM)QCL-4OJ[9f4@0V#6(T&)6#RP=cb>>RO-4WD))/]cCKcP6W6R=XD,D0f@XEO
T35ZaGHgANA6X5YMEM/E&N)W7R6D:;5AM)M>?0TVWS(7OFM;_DdO<)=I@^R7g0@T
#:-+[M>1<@BbE1EcBC#JF>\bM(@F<^=@V&a4/<[VA[1g9#3d?>bXV09@_NUV&+70
2O9@3,]CUXS6(?^aF0]RNE@dW);S]fWgDHe6,OT]a2D2,1ASO)#Y&Y[L#g66PU0d
[9KOa];WB&YETHZb/D-Yd.5?FXO8>;V.5/W4IA]C)C_^B8fa1;CRd,HY\FS2YKC0
LQCdW/f8Q=[D4@55MR70>BTA)?]ZX)aKB;:EC;A58e5U\Z1;V.-L-9@adU^JDVDA
J&);gAA&ED7103V:OJ;cD:>_fTHI::[9;,TK\9>RJeA-TSdP2GOGB^@\2X^eKD<N
dT@<KH8_?27Z&ZS#a_6D^F.?MT.;AeT)7;F-+>d&b#W)ND=13Nb<3#&L6_[)8b12
Q<2QR;H8\eeY.K+YF^IH6.TF<FgE>71SGRPI+H(.IZQ/1b;.FJ#ef#O\_Bf\SG6.
.1:aT(E=;Y0S1.>ZXH,S(2^0DJ[R,-JRZ6c6#(aM/\9UU#,<(H1K02.:8>M&Va0H
UY4;(eKP[\>XIJ=\FWBW73-C2VaG&0[:C]XBLcVg<b2@2U1#FCP>8.OG6gD+#FFX
e)fTU/LNF3UD=8C7b]f&X3]2:G1-FW+[,Eb@)KS\<8?FC=G?8[H<_YL0G>TCIL1W
HYQ+(J:>NMG]UW17N,g7:R+B2Xec9c2X\#ggD;J3),]6??E98W,2H.U6Qc>917>5
/CS=Z4D)IX03L[Gade/2c)]gY>HbK-SeOANX66H;Xce\Dc7E<IMH&Z\fW_G0A?KU
=R0-2FMYV1&Iee^T(6H(8S)ab+<Yb2E6d^C04I=R/G54TD..SS5#Z@6F?4]WB1^1
&=O/]Z9eHD+a#:E?7>CPRU@C0QGc[QSgN4WFATQV8.?K=f:f+15PQ7a<+NgZc^R#
/YJ8FCRc(\LGZZdX0e(R5d2bCI,VBN1NU#3D-R:gY@@gd-(ce/Y1+1a64C&[U2Ze
:LA-P<8+ADGZKI6^MD)6#Z1MRG)&O/A:OC46\.4GYB,P:W;1^?1e354Y1>+,WRcB
afR6DafN4bPQMfU-P0./((-(5.T\#]D]e0NN;U6+=/XFLP\9(WUdHAD+O[:Y.@^,
UREXNEQVf\=FO#)NI7F>@(J2G0J+VZ,.T+dMc7a(I23_WNXC<DebLZU)^ZISVIZ)
2[YT=dBUKWKCf7957P?@2&66K4HfTHEVLafYA1IbT[<eDJQOfeffPQIeS.?SP[&M
g)Ra4fB_Y4_a1P.3,f>T#fZ@[WgJ2L?EYFNCWXS/RU]+U+cM>>@51KaA:SSBXf\[
.&);K-84\J2AL7HQX_gcD<V>@979970gQbdG6J?V,(-DF0Za+[J5.HT=1_>U(-^b
(CRgbX654gG=(YBL[E7#387d&DO0P#W0IO2b<@04H+PH5_L@>0X--(?\V^(W^U:J
(+_[ZLTbQI\._SJQ<OXR27#K/<JEa_9&S+RdfNZQM^U97OV)Y(5D]OaW[39O\G6b
g>JMHDIXPX;9f@TCBdH=@MK_L93Bf=c--55;;A[a3N:I7>O@\;JgZC(5WS8ZD7a1
B85X8B5BUdc(Bd@CaY-+N90A9\29+1e<WZ88]&/A:G>&+JNV<ec8CF3JUcDfRXb,
IW#B6Lc9LeX]DTc>H6;HdI0<Ua=->edE+Y&[QX]L-Rg>Y67_W?TL2;JNg24)W_7T
56SC<R]5:4B\V)d;W(EV:Q>A[gPHS)DaNe9B278.+?7R9AY3W&?QL#J\XPM6c,+O
g@S]a:=:E3OC-JeKb;LP[G+J+=Te+JZE5bI4..7g4)X.)N/b5c]3>&DGDd>K4-=(
Xa[M0?eZ7V4ZK(ET4caTb<.#Vf#3e,#+=I.XbS[f)UOUW1ZF1O)[Kg-e>T>/>>V+
?[-;[=1g(aP5[N8a59Sb8T0=:49:fGQ&E#&_6,31UR8=cH0NHIP4d^ccBNXQT>3T
@EaH9._<A[8LW1dS=85af6PE02GNB:/V?05[Sg,V+6d<CfQX6GHUe#aR46;CfY/1
9O03HeVY+9;Z(dSCG[FS2fIH7RW[bI3bV^@N1DUc6;#:>];@JL^,1Z>?IadIE;YG
UMKAP_9:aVTb2.6Q275@gIM&GAH7^;(4FSO>b\UBg>3D4/Ld<319<DVX(FGD,OPC
]=W=^27gX4T=#Xc9L000AEdF7O.^,+1Rg?B:]]Z3D<c=EEZ8[IgNP;b+3T8Fe7(R
^+L_OA9L<c]DMdf,8I(((4@^_/?gc4V&Z(PLE+f]aLB6U[C>Z/fXT8@H@0X^GP6Z
gLA4CS[eN./a;P8814)-F=S4;(5G_5)DGcPYd\<fFJ10NeA^Q:=\OGA6;N+_ABF(
.JX6GJ;5>;KELAEa:#5dLTePNdRV)53H>#ZG2Z+E6e[ZM::0=K1;=];?4T5]2QS]
e99[U>[#<@FZd@bF(d?Wc+L2PM17=O/eHg2M<ZJ/PWF7L29G:&6bY.6V]#7W4D?+
I6^<HSgI8#6U4O/S2;5HccG10-HUS.eDagUXG?F^18NOd]<2bMdX(GWOGHK12<EB
<c\fA^R,CGRX8aWH2GAN>;;Y[2A,38=-EJUZ.(D;+f,[Y1N/40^O_0I7U(8f_<<K
S&SK460gMQc67OD)c5MTL^#1VP,;/V#VUQb>8>+.&++d1abd645ae7UQMMdB;b<.
VXPEQbUDAB<NMZ]:cX:&S4A5]@KG3-bW,^dBg)O<fVgc&UMA3?QZ;HYfH-CHJJRA
)XK><4//bY/DB1Rd@9R3RWUN:(gSeP<J)4]8]RCH_AHYHBQW&ZaZF>QaTY2A]D_^
MfNQ?6W;Ve&?XDP2R)0(1JCbB;OeNJc:#3ZTFE<f-HN@6]#IN1+Xd7/;-FLe)cf6
_>P9Z)fa8P6O@QMY9O^(A3ebd3L^DL<7<^[8eZ\MTbb>DdBc5&T?_L/2W3\HNBX(
PX8b<^0D?+Ic=,1d&DZ/#3N;JIS,./>PG94BZd/;+4g0X_L5<UcKRY-Z]I#&-O5f
)JMDY);VFGUEX]T^]?Wbcd4XNNAEb/YT3\^[T/AX&=#?DeKHZG8DG,KaH;^L@dJ2
4<EP1:0eeX9fd9AORG3&+@FDHRY2PMN?Xe?YJW\PfJ/JTV<-9U((VD-O@-bV.E<=
;5d-4MXbKTd5@..YX:,5F8e,Hc[)@CaWF_#TY8+H0DJ?9)7/P]b>WbR6FT5_g1[E
PDF)bFE+Q7WQKTI5B:4;?Z#a2F.EZUUC3QN5(R/KS;cW\W:Vf8Y1c/VO3Q#[\/+I
PM>OP=#8B-OOTCaZdb0ARgP)FQB_)6-UBdY;AIV-@P2?TJH\P#e?A.?.O8MWVeO=
GAZ,O?4[LOI9KeV#:>H30LT[+,\]:OMM&f8PNCQVYQd9Y3.:ZUX0,V3<&0O-6+(7
5)b(DM,+c&S&8gGeOg>dE1dFW+CK<SFgVTN]0+bZS:3_N]<LK1XL>ZGZSZ[YEOLH
)c<\G:4O8cgD1b)I\W+]1+R#cBP=BH43E=/):bZQ[:(a.96&YKXY#8<QCf#[g\#g
C_DF5#=JIXHPM-CWI?X4]fW_[Z_.4d@7_P)Q[aS3.G0TGg_G8)3JY,]9WaY.c8R)
5OV;IB=9XAePR3CR83/<;QLS#GaI.EZ[BgUV():6R.2SU[\b0f#f(J:8c4ZQ5RCJ
>R]97cUd9D1>,OR5>@?PAc<_?0T?fd/@T^efZ)e.2=(EI]-(/TMU(;E1g^dPT#Q0
W>L-RZ[#Q1dLVSgS6dHSa[U:?7Q[HJL.])=;^E<XUBFZb#0-LZ6+<G/(>aJbHf#Q
KI3d+V;&NS?\;G@S7Hf4I^G<@@5[8;OY\6_UP^QYU0OKHES18HgZXWaQMPZAA6Bg
XKVF,M&dZT;EP,7O<;+cFSf687X)/5e9/F(/da6?GU)F6K7M#-;8a(34#3:gVO.3
4EK1JW>O/TCdS.U>c9_85UW:BeL6+DNKAg?d-bbZ]KaT=G-YY1NY0FNQ6WB]2E#N
fZQ3efDg?AfO8aJSZE/f+.VSZ@:0_FEf+>d3Y:YD.c^f#WL;NZA,:JZ-WRPYOe+(
7ceO?UP-EMFA<b@2ecZUgXFB,:].2LANI?dX.K#c2#3a4KSI.AU)b9+8\A]F8^[V
N?2-LH,[[d#1C7dVOS?FUdHXJ/SQ@_N/Ac<[Q_.F7?GG?,[#:DgL/()+CH:4<Fe]
3&(,^AE>SC?(99_6EVV_633#A==J[.<^4CQBeB>PcP=DfKgP2C6U/;ZA)A\/TMHA
Sg\0d5.X:eHUC.6A98,,XV2(.eTUJ.++6)1cbd7-#NDU(-E/Fc5NI(6e536A81:4
JOY8]De\#@CcbXN]IcOZP908)XHW?BL)b/@<W,=cHLP0..0/;4[2,D_/^5=R@1V3
_6dQM.6/fDU-fDb?EKOP:SfdOLXM76:GV]ea,YgG:g#aUU7F0,Ad6O)4(FacQ5HY
X[Vd9M^LZ1A_)c-2:E/5WMH\7<K?N;#Rd2g^07Y<@_E^&If@GKH,-Yf<]c+4)BY6
2ePUGW:#EZM_gABD@6K5DdTG?<Q[T9=6_8TRMfWQ@W]^&YC2]@F@Bc&0V&NJ/fTS
HZ7@]RI,KT^c9aVYc2D:+/X-EJJK)[c<WGbG7<46BN/89R<+cE?2K202^49P&T:M
KQG74=&;;J3]3?5]:_f4Tc:[YA4PD5/G.FLGS80CG4:SPaNfY<If;DgaK-F[U-;0
>P6AWSe[L>E3Kb\2feT=:3Rcf#T77O+XMJg^;abgY.f87,/6Fd=gL7KF/KXE:5Y6
MMY#)#/2]I8Y0YYDKP2db4&&8b=1676GO2aZDGP&-M?I(3,AXdE@8S4f>\3c4EZI
cVL?#Pc:93LGIWAON+&\X[@J8-FH=-g=VF;OMa\@_gZ/UOU1KR[b-d.UM8A5e?#S
5/?Z35MH4L&/M7SW5LU[;GbJVWQNFc1CD\484O5ad3JAfCf:OA,_a8&#4K&OO,)\
EXVFWdNaHI:88Z>DD2BS_]:<E3TG0b03Tf/6OX&+W.24-Q+GPTTa2IWc81YU1GdQ
&:4102/7ScV]=W#TGd8U&BA.?_9R3HGT6)6WR&NF)-3,K[9I;UA@S-&DM&d4)CIM
DZe[UG<g2K3EXd281^9I.C\+XOOeR>35XQ;a7IY4O>B)bBbIJcY>GK/P:BeYLbeb
]&@/)MV+0?NS?T;b)b><W+PIe+daGeX)HW2/:=N\LPAWdGaVS5P=0ZIL6aJR56=P
cZT]P(WLJ4,04B]];Xg^FQ_g4>agFD]V0J#1+]bDUZN(B>PY.7b;--;16YBcL?59
61^GBW0.c5Nc2K&_/\YOP8LKT@=?V\?P0ZC\c1IU/1:_[f;:,-GfdJ83^S\)/XZR
g>_dQ1g&e09Y43JU/f);[[7J^Q/56[3c).H_H34@IP6W;7HK8G]YEAC&DReYdMM/
N6NMUb0c?;CJJX(#803O=RJ,c06[>(3d+70XTYGAYH1WcPM511cJcOa^8Nf#eA+X
8/90GK)]4(U5/]<;VEd:0g7Tg62PC1XZ1F@WYBcR:YFDWGVe19VF.9+RSJE7H1R1
]NLT&W#)De/IODGAH8ZddeI7A(^/^=b</Q?H>T\6FH7ORKOQWNN?JHIMF?JEE[Of
;UKNBRA>aIgS[OO)O6RT6@4N>-Z@@QRb\\6\#f9#9N.EbUO/;H-c:0bTOYG@^648
J0SF7(C(LE6]YN5>9dN^1KUW^IBMTZ1,V3cY5Z71;>:FY)c@Zf\0,<U^A@66:WT\
I1U;K<)(g(d_BU01[)aF<_1(DKdYQ1<52Y8KUH7#1^f:?E>?a,3CGb]E.Egb&DD@
-/gB86FU[E62YYNJg)RC@Q2bAY8##?U#9fRRVP@1UJM/W[CZ/5-Q_Rc1S\Q+0;I?
,&A/^a;ITg90^]:9aE1>>BI(TX53DGYZ<>#08g84:5CFc1\BCdWO1OQ<R7IYH)9J
1T6QDE@7@e4+/1D@fb9L&)O)GR0@BF[CG/67X.cGCBH3=c;#C0Kf9aW4[4GUT0AC
gcJG167D]8-Qb/FAT2[_FYN4BUGVSK&V/PWFgR[Q/2:8@Vd5J;gJ>C>ZF?5&WbR(
Ab.aGW([2-RI\)b8\KVa9\aUWX(B^W0N._-^.>P;X]fTH1B=5Bc<]YD^)bS_Na-8
:gO=_GS4R:gQ:\1d0G@P>64K<#+7f1-2TJ.bDYD:_ZBgA1?XfI.A7L2@(&TJP:[T
^]D<D+A.0;WK_B?Q8W4AU53XQ=PPIZbFK,0(3Ba7I,d<b8,MTN;_2YQe(LD?6Y2g
d.Y)I#T#0gT(Xg]R#8?Z;1LFcd.BC_#O8#)-7ZVNZ8bOC8c2c2^:_M_+-H&D2cad
>WO50=QZV[.D46g\;/F7(,M6-<:^N#7?G30Zf?Ya_\6)FFS=RZ>C::5\;J\,Q=(M
=&gT41)9gR+,5151^;4]6OF[BSY6B/)Z(5NV?(RT=914E_+^VdW[MX]JBa1-I/c.
BS=UP>IKLF)4)1-,VQ]R;VP2Y=7UGf]E]PXA2\QPAVVKJb.)\7J]\)d@,ZcST3GE
V(FH#E?5b;\HSJB2KCC-8-(aV2DH^WI2OF;(<H4acT4?.FH]DVI0?JLcgaBXM7F[
T#&#e8FT6\,-;aeB:RO1#=de^XF#35M?(-6)[(TRO[AK,aFb\(,N6YULb+><]0,U
^?ab0(QY)WO(?,PN)Yc#G-T_A7W7I(g\gg2HUCegS#X_<cH]M),eZR+I#1P<UH,:
EB#Q^5^0a+EXR\C)afG13D7.cZ;Rf::ZS-W,?2M8M@9)WB?Ja1(OPNLRE77SPPE7
P3W]IXOI=Y222GbgM.b(J8FMd/KRPLdT88H-=K[51#-C90NgOX]D&_7\3;4,9T_]
f2F.BQJfZW6.MCRS#F(Q1D&GRL@ZZX:A:(IK6ZPVN1.-S#)]0f53<SZ5Rg_THB7(
2>_K-UD^WUd:e6gT#EKF&d4ALMFE(T]B9J.DQc>41b.2=eFcP-?,b#HH7T3gg.gO
E4\6)V)/1a>7@(VQ9+gT)3c632f\;R)4F7I_G^YL1#=H47,bV3I_HT\e?N)=<0F]
)?C3^XA6HS:c/R7XF\S[?++-b\@&/Ne6D^HIS56gd(gMLGVUc57[SBdEa+?CWe4U
/[[-c^WS-gTc=+fP]gEW\/8G+\K?CTG>R7#-D<#5)fG+6Zb#X@_/UUQVPY7OIe\3
2PIS9NW7)RIFIPdeI>2PYP4NF_Ued/Wc_g)&ULeRR.\P8@1NZI58a_MgP8Q+9&[7
PWOA9X_^L,=E28b3>YZYK=322T]C31cBJa+0McC9GAU@BZ9A^5XT6I:e3X_T:U,W
SP0?Mf)d2PMFA\cW7R7f#^bAg//4U[+b4UA8f,V70a_F<TO@Y9@V;;-GJ^f[JA83
,gF?U]@J25?CC-S#^N/L<AWDG)0XL;6+5SK4+C@gD0\a(6S+UaE^PafV)65)<P#=
ZC_b[@I=X4IbZ=X;^GU?@CWKZPfQ]f?D[F_U<B?P?c0b8BBXAN7F;dTZQUWRS6,A
EgW,?I/OcAFWW3920Z-V6GfgQ,2I.DCdNR^>^GceMB?4^,E.,SES6AZ7c:S)H3UR
BG,?B5N8/-[Adg^M/CYM/DfZ4,TY09);WNC>VZ:Q88I4ccLI@[[/EEB-c841UN/1
6LFTb>g8ZA&Ma\M@gPPP_]bWT?0CJ9N_&E3=dOGQT3K9]-4J<?;U>T0TBQSgaR<_
K;U8COGZAE5]>+EI+D=BHV.d:g,:9H\R\QfSfX.T^^B>CSc9]2PY].+L2X[G;CQf
9QM2/TH1Q^L\>&Y[S:>>AdL#>R)O/Ff+Q3T=:RR-YfJ+@WU?P5U#GEdOAEFN0bTe
8a-V/+4C.XQ6I5[U1)SaU:0)#.:Ue:=gS^<X)6<gCS6,b)\IBaeFV2eUQed>SLX>
dY8fTX&_58RT-4UQ;4S?V2YSJ.BWPH77]DAL_F>,Rg&:?1Z#-6Ycdc]22]Vd(F4L
X23]J:;ZU0bbOT)9Y6bRX4^&R/3MOS.VO;/YCaSaGSY4Pc7\+6_U<RMN6b;5W5.#
b1MN9BA9c44YNGUP#2@]Ld4[A\XY_TJae^GeX<YDKYB5cZ_MXY&Ye4Z>6T;36[)B
Sd-WE/Wa^=6-XS8UdE[@>6dIY)4eHO2@.99=/bZ0W&N\]SS,8.[L^@dLFeL1?;<-
2VWVgE)H.d7Y=N1?]^/_dDWV9DMBIG20U;J[]fIO/6VI^@&NPNFeH_RP+O)H3g?A
1Y1V3BDSAf4)EK@Aca;RcDQ@XTH<6V-3]>IV9)Q)WR;SOS+M8?;7;E)=7J_JR.UK
O5XcSGGSYM@\c4K[DdSX/FZdY?)eQ.g@5_X=g,.OY].2T&IB1&Y[VaXV1X^+S#HB
g;O3ZCO;,&LMc_(D)A,e\9ZD/C<(a7B/MY+.202)]C:B6?;@3,^)F+YDcRF0@0N=
L:Z-4AB^ec8K_Cd4Ta72aME=UQ=42D]YB-c1Re_N0^SZ<8)0U#;9UNa;;C+Ba6;0
bH0L#BDA\C[e)FZFM(#d,B2UF(15McNc9.K^E/N2X@d4Ua/5IJ4W26Z+1DW/V1E<
[G<\LP\-&PQ7R:>LDS,:PNHR=IOW4N:g9FOWgLc2_9G+g;Cd.:3Rc31WJa;L6_;?
Q:0PZ.4#6XXLWG7]gD^4#(^ABYVFHS/d?-:2BU:0gSGB&G7)S-8M65f9gW<dS=N)
MNI5V-<?b8/T2CT.eJ+8-TYO1T>@B?7WJSO/AG=a>[WNZ?U,Fb7_=dacNfU^JY0&
deL-JD]90OX+JSQO\1E@cZGM+7]_bcVG>WAQ<E#0#@GB)<#W(Z-+1]_^_RZY?11Z
N^]0KbZ1,Y1FH:+Zee4Rc/@YNP&XRTCY]I?XDW4K6OG@=-)PSNH]9)F7<)#Hc#g(
bK,e[_J^Y]54_Y,a4??\TT16?11bLP_?1@f_FX>-D?X0B</_^NDe@)<fa37eF??>
.<T>19cB+#8Yd3C2TP^V_4=H3b+DYQc[5==AF1@/d1?2G3f=SST2GR90Q<]^Oc-]
S?=Y>a(C43-0:JZ)8Re8MD+Z))b)S7HVBb-W\beQ013?WYJP6=N_F.;AW;V?=P/9
c>Ge.SK-\&G=XS+7GLRKKUJXN6<77A,a[ZBCO8UUZ?:@@HG[Y0;,Bf6.-\3:(QL.
VSg.&20JQ1LTZ5Y@TFWD-N1c=3H)JI&Q=6=EK-;V(Qa@X1<<2gWYfQ&#[-AVgO86
CB+_B3.e2RGALG439>IXB:V)9b6eg(MW]5=^eKD0<>X)O/O_0&F_Y\ZaaaG(SZ1T
N)11[U13/c>bOdGb<ZCG)VQ(N7QK((?cCSF^c9&Ob#HC/.K^E&P?RTYCI]MfcG&X
8T01-/^0+VgX3Y12a+B5Y,:b.g,BNRKIDAXb_[16QR4-CFe\KVCc;bHR]LRG<DG:
@Q2)g89K,)OF9YDf<(EE8Bg>;F(c5AZT+H:a\B9aJF7=2)\#QeI2=6-+V<MbQa)I
d18V,]SeJLbO-FSZU3<3[,GLXRQ(/ZL?+]<YJ.;eYf[I:+0ZMaQ56dO?_fXIc_:_
2+:=4JE]WL&;,SOL(L4-Q#HbdS0H#K^E#R?&J-X:3I=eL4GE^-CJL,HQIS1Y3c_e
=4^F?aDe29D\?A,.)C018^=;b9>E#&E5eJg2#dG[I,?=M8ZH)#V//>\P7O901O5&
7TLB2[Sf/cF1V#@Kec)?AU<+(60Ba4:0&@NBUQDQ_55Ye-ZTQ9S:I8MGbfP(G6/X
0KDb/W75FIOf9)#0VFI9<;&&[d-0TGe0Md<<:W6B+.8&O4eT.-MHBE<<6//ScWM.
.Xef:<_Bc?Ff0R&J3(<#)I&XWIZaW-C7bBY[A&&3=&QJ[:b;.fKY,[AD&cZ6Q9I>
cL?@JYJ496DCYB>80M@dgJH/g5_>9>]9XI]c7;L_B+]IPKAL,.g.EAM3BC1V8=<-
QW0FIMUD)FQ05&)&<d((-D&HC--/Y.Z:;9-fGEGZeW4(Q#QJ)fWP\12X1/HY-OAQ
)14JY3@K=)3=]U\)3H<Q6F/O3OPQ.4-5\fZY:RM193NZ\WbPe^L00^[O9d?78_W^
LEbJPb>HY]d&C\#/fd8.IBO7L1.<HQA(b&J8?<&.NZHGDJDV5LMb<,NWCZ/:NdQY
):#365<60dT;2I0830.?P0Q1Q;\ZI3Q70FG]\F[&&+:]&XTTY,(GTHXb#(V.dYUK
CM;3J4^W?E#f5(N:;+IS.I)GO0#I#&K)31]0(gQ?,LZ=e5Dg)^IO3-SR@Z.f87#R
(0^d9Z3J&ZX9ZCFPALV8@TWT=O_:D6V_P4XQF[SgVH1a2/GbGAEEd=YBZL^96@]U
[YZ>OO5HGSR(Y_Z8;=_8+M_)FN=H?]@,OUV?V<8_GG]0]cZZKaKg83/R_PAdGKA(
4Kf3R2AZUC]>I1SaX_W2&^>HA8\)J2PcV(>><)gH_c+Jf;84fDgMFM0<HN2UA7(.
JJ(ANcEV30.Wc_MAJP6&)<R(>X\-51ORAGAQ(9UOe#ZX1VJ>&D7.e0F>2,f:aNYc
X4&#ET6A@.JRP.GdJ_I?/3\cH-/OO5<T/>]H3CJ5Q:?YLKTB5,P64=1[UNP)JITK
dUFdQ7:76GSV91/AXT0>JPZN0B-_FH\DA7]/GDQ)6G7<<\DY5dPa)a?<VdaCC&+R
NQUX;F=4(L/?;QgVWE#,T\.1T,UZC-dDK[N5@OIQ+7cTMeNVLf8+-)2#JW\DLPUB
3K@KV)DadeL=JQU<1\.F,gY+LCD44XOcA:<b?G9AP3NF=\G58V6^W2@ZV3/QIa+N
<P#d]IZc+D2M>#ZJXfJ9;b-T/f_Z9=V\TUK;C,/7YR4:B:R8ZTcdgX=O^F<++KGf
UfcGH^0LLCfK2XEO:DKDOB5N9L[N5.G^MUSaSe8^=4H]=GbL;X&d0\\Cg?=&)=9L
e9f@#4C1Y_\QQIIM&[])TLdT2SdRU3e_X)LGFJ4Tb6>KQ&VO]:Q9QgOL_.QYFe0P
d<J[70-6)[/RL+UE7+T5J-J\Q9Hd#5D<A?e5:OCNecI9dUSN<=D#[fUFJ9QVE)S/
@=?ZN<(Z(VY;5f-.&W-N&V,0=a(-ZcbP-K)e0fZ>aU>a_8AeD#LAK7<O&F(=H2C_
J66C,+<[UdaGFOS=Z-7;T32dG@W(?EH2Og@bS7R=?J,H^CF<S,1cG4_gFFXDR&]V
c^bXR^XSFeC#VK@6[SU<c86<C+@g8J#ObCG98gKX(4.HK>.f5@V(.\f/6bPY9:.L
]fZHT(cceeeX;M0>ZC<Wee:BfP6@KY5^a6)O^AAb:Z+F@)KYB8FBVBEK]GEIZ<7N
X^Y]>VeHN20X=bU59b(:4B5U(.:N7W>&JB4QaF<1dg_S/V+W&G;?T3+0P&33LP(S
<dME89L6CCbee6aXWQ[7e\TeUD;L4.FVF4TQ_,D=[THTRP4->?eb^a<U:5JgR>,J
BQD-QfKFNE(@QYc8)>YX_La:5<a3Q&KA2J2G_PH029.[O/XdGX3eUH<YW13aBM)[
#&c)C?L9((_Be65@/QXW\0gc=YbP(SHgF#-&(;Ib^/BE=LPQ;P\b<d3fe5T@(\&B
5^8)G0@,e((OeNX+45-L:_R@]J<_b(]?TM6f0)8<fBH)&Q.T3B&(M034)XXL7EAU
We8V8_a9X#DQW]=32+]V)\UW(J7WdZI(ZU_=J-7eGfL=T8QT3Aa/UH:>3@F@&.VJ
UQH#581&WCeS1g0;8c-WPDc[R>8@HCbFgP<b3L[\]3LLeN+4[G-N5aWBB[G^=0C[
bFW<5GHPK<WeK3]JeH#G#20&>?e#-#@WfN1SJYVR5T;D[0BVbd1EFC6WT<S/M4SV
P.MMOVS5U13<&cJ1N1XPagc_XaeJZB7\ADe>UV+]W:7UC):R^=9QL1:c(.3g#FZ:
WaB8G9XX-,dUCAeQF&?1?^bgb,_),OBR,\:;[bIDT7XNagJ\&1A.\0OAEXB8CeY6
7LZRFG:P:\,b[a+,-e\FY^]I#28?WJ#]4STIIHdCHYE@9[#/X19)aA\:C&bOZNFS
>)910cQG+bK[<W>5/_CDG?/a<B&.RG.9@+S&^Z<[KfIR]02V\@VFF^>aR5\JM7.X
>EX<-YaH#VS2@MgXOOOfB/ge0,0NIFIb8U4CTQadH)Z4De&F76L3-;JNIAE@MREe
?J6a&L,^CZd@LVFE:cK0W#.gD1+:XB/@+):E@MG73@^KC2]Q-D=93<9):0\_JBM6
7dE/]DMN6F-G<6]H:,>f)8+NfY(=BZ6HSF0=\;7\aE#\^UIgB_0W@O?(B<TS)2@[
e1I)A5IA),L@X]c&372;-JXTQVN#3XDF1A6/=(\WdN[=CA,cWC5#;&d#3e-ZIZFc
T(.eYUM_F]0/[^<0:=6=e768WL)6Y=S^-T=LSe,NE_/X-EfIbI:0U^CG-A0Je7#5
A\9_P7(<4A;8Cf/^=JgVObVg9A[9W)4T(/7e?Ce/.2J]QE(QE,DTQbN?;ORXF.8/
DZP=,X0#\J-UHE<-M:^I2@gA&<U/&TN=Q=U=[9O?bLg?SSVN]SY5Q6-\Z=15F[<N
T3A;>4gf5L4PT[Z-Z<5ZHC0D/gM[V.37M;cd@e.16\.NDYVU[fddcIFfD\7(D]eJ
._POg6eI&-[K^&K+M/=GJ[<,(aO^:eadU6e8#,e(&cRc.:=fH,UeeW=XNdDKP9?J
),S69]A0ZD)g/.=D-:XX^a(U#MZK6NX=\G1Pe(_S2\Yd]RT:_C>fKJ<CCKIJML\A
PZKQRd##@L(]QGC83IS49XQI+PQ3OXI11C69\,7WP/+U2Ug_L4T_U.5\36(P9#W?
Y0adDIc<a.J^>,_4HVc15O4:3&RM&:A1YQeRK2-XM2K72+d2Ea0(>D?B?F[)]4J&
:D>ATXgeIL&DII3c,URf1NJW:2#1/(VR2d7]PeOR)ENX+g1df+TS\0AC8]04MC>Z
&>/4+5SLWATIE^6Kf1@.0@V]2A0T9J6F(R2[2.QK^_7R&BdJFUQD9&ZU<XN1-1B<
J:=G.ZgSK+Rb&V.KAAL<9:H_T(<+B+G>4Y3BCI,UbZA(a>Wb:IN+QbK#aagb.ZV,
/<KeG/U=45(KgbMG/O[CY@Y=A[-fg&1VY;0#:#I.(dN?NB/EeIK:\@8+/)a^7Bb2
#?,/2[<EZ47;THc[eE_;IIbEOWc?C8[#=9A0>Z<68:X3/(1)UB5;=P86;?f/CNCJ
S#Z-&(@I>;Sb[/_.LG.gA@5LR[XAZ+18?WL@CeS90EfGe88Qg9fVO16K09;8WZ2_
F&d:gF#=AGW31#JaYD(]D(H#((9<aMa;NU)X)KcI&\C6Tb_eF0baQM5[V)]9\4M2
OH9;c=6TXc13__GbGc&UaBCLIN:MHCKFRU@-REdAZb15-A9W]Z2d;I=3IZ<:5#KQ
Gea_0DU\AJ34>^::D/B&VVO<]VA1IU:.RL:?V(<[NRA)9I/(:8BHWQgb\@2I\=,O
N0?aHOC(c5E).H(;#E8#QH&4IK^9@EQAL+1#]C1^5\Z<2VQfCQ]d?cc4VgG4C<_9
:bF7Pfg/\ScF5[g(-D>^NF,^3fVF?[D=+B/POWK)V43B[aC(OK_Y5->aL7BVYCD3
a#cI=f8_5+G+BG\L[T?f>=A6BgO83J.245b&^/-_ScO9)4ZW/c;&>CE0^QH)2VN.
OX/c62M6KLSLZAO0L)L(H=Y(9#9S:0MfV@T:/TOENeO;:@a?7D@P7_-\Y/CT3+6e
74Db6I8@BCAMNdNLLY9=]F9VZO?#5H7CL1,^\4CYIDP_a0K8eAFHGLC<Xa&960;\
5QJ[g1_XI@3cT(RdQ)ea;<HH+(@EA0b=b8P)HZ-be_Pb12ePG&WgKBYD05ZfLeAF
^d\1L#J,_^Tf7_2YV49;H#g<YE:^.RPC26_a9^XT]^&-]=ZT.;dOZ8&X)N>LVLJS
E8f=0PX6==&P&^9#-g\S6]4Lc(S6.=g6d776C-a3&0=I_5ddM1TEWN4L&+=I@gUP
@Sa_=H8XVO;Z+bMH8(6<R#>F,+<5_:E66S+\RFcT35bb>(g\ELINB2b-XT?2_D00
Nf4PeZ,e?/EKgYY[.+dTN>7SO5fdT)1L?6OfGN-UggLR(?gVb7PI6QF,3[AO1b_J
Gc_6-c:MP;Z[<7X=dGB\A<+Ce.8cgYJ=<c_ZHa6<+2:\EQ@T7+4URF/HM8J5VW(^
/=0,[GT4&\b],TH=OCA9>6&8VH#2(N+gX)EOSY\9WP_1.F)8X@=@])_BU4TY7C4;
JMVD<N<RQ)8X/5SL,Y8cS64HU#9bM9]@95RF,I8VTV_TAS>::24+,T56R-:7T\f=
LC18;,YN4c[?I+[If3:86N+@8Tf^SM&?A-UEOKAA-+#FJ5KN4/3NXDXF-L)2.XM4
UbfJB&?)&KX2O1IWWB>SaISPgYK,;I]_G_GF9d:(#,U7g-O8?X691IPQH<0]EMP?
^EW@e+11.>P?O2&\:T?;KKM4bC^5MXSF=95\_XR]<&,:@S2P2(.=g2X.DIeG,PAZ
d]4^0C,-@a36;]H<B)VJ<[L#UaV^U4PUORgJUP30e7)2B&OJ,UE--a10)N_NCNHV
0=D8gF8#a6HM2ZEM6-EJfJ=.OQ7GPV37b0J(dF/(VaY865=BMB4ZVHd/R7B\e[;=
:;)J#&LSf]dHDFfd?Y?CJe2OE=aHb>;+@^Ad/RJ@<GC<PS<?9Ic\>APD(#^\85I7
Qe^HN@C(U\(2F+C]Q8B@1BW2>/H/I@,@R8F=UA]&Db<1;(/QdG[YB-RA:>?#]Id^
be6&.c4JM#8/EIT#]UQS4dEQ#Hg-gUMbGW:KC;+TLX/^?RH+8/:.]]Ue?d(aW@5O
)+ED</-D_g(6_.4V-(XHOVV;GcA<QL[8Aa0.#_W[/SGI5LM7;W5:G@>.O[fe/N@&
62KVLTdCM52B^7Y[4M?RMBH)UR5fO7AVIg]Z&+.TeN7Jd+G6RaHc,+33[/]9[P6B
-3eQQbU&&=0:H0_Nae-O28);7-fSEgNFP(2fZ9VaVY>B=^F+P.)Pbc^X&9B@100]
&Nc?W[A>SZO>QJ2J2aS8,RC,Z#Ia)[OEUM#0+^a9a@+FN/NE@F](QdFeK-.><X&M
-cgNUZ#X6/HPAMZ3e\S<SAY_^S<bCe&&a0IU9X,E,gZ=#L;0NaE-G,7HGRJ^UXX:
&L#I_G7fWYNc=M0(6Ngd_R0K)M9U?5+SYW&cHfF?=]\F]:fD402P3HFQO,b-acfE
BM790+V6W7N?4P1)#IZ(c?[<-fW<G7VB1&<dP[MH]L])E1dYgHT7YZ^0K@93#<ea
;AcYg;U)\M,a<CZ<(L]#e8I^/M&e3I#]+EZTWJY]7LP6@.71/HBU@g08/e,-@=:K
,DA_=N._0a)5#0>fA-PS6fF4(GQUZfdHa[Yc<XO4/KEPGR,>aM@:K_.101Sf67BS
NXQdUO_7b_TaJW[(gQXF\IL,@c]H3XT2Z&RZ\XcTNGcY6c+>Zb,a;1P+Y2T)-67F
#.)]DC,]aaQHAGL@HfT:aRQ^J0HDZ+<gHcb23@M/ecI+3G=[_PXW39BX;J6c,FEV
9OOTb9=K1Sbb8CIOUVM9UZ.QV4TVJYIWK4C@-d^CG^Gd?V+-3_PZK]?dMR=G7FFR
)5,0\4YC3\YH8Rd>O3)gJU/(BX?.eJbPcD<FY#f=-3FJPFB;K8@d&WU[.c_(S^&+
_cMB=]7F@)YE3BB5<C+YIa<b1&UB92_fD,X^/QX[:5^L]bcC);a>\WTXef&N_d+6
f^?NY:>85A]+)#-NQ5NY?.AB63P<I;d9f4LSJ0NENT#=/^8Y\@2OUBH5(@?8Af08
1aRF9W9_Mf_fP(,fITS+UVAT]ZDW-))[cb^PL)Z-I>g8.e<P48)fGUfa-fSK?E@+
PO(gP0JM@^-AZ]b#(8GWYUEIC@B,_fb.&INBY<ANU<I\Cb&]OW0]<+Y-J>632+V3
5:WE)WSIeb3c(RWe2g_M\[XY&+eYKT50UAS;a3d-eNMg8[Z7@BOL4S-@c6>2W[IF
3<Q^ADe9.(g98XL>:d^/bM\Gb_9Na;;fKD0Y0>:DZIJT+c,H?A7)2WBJ#;/3@2BG
UbY.V7Z3[cI7Q/+:+d[\4@(?UDF0;ZYcI/^O=47D(UJA@U7&?>]G^a&9cI&,9f\3
YaM>ZYF)GWHI#&J3X>2EY7.BYX+f[]dA]e:9W/bME,Yb,4>.IF/;\3MMQ:&,TJWX
.bGX^K(OEED-8g</70(/BXB_9@6\\8(B2Z3@\]Z017D\:\c?D8c;ELb><AdQV#MJ
/bbUREOHF3U1UW8PHFP.H0Y=E,AUb_LBX2)^aD<8?FH.B-B#?M/GHg;+HfU/2d\a
&:TX22be0)I_,=N3;2:66ff&6\-BTQUB.ZUD(F(^;aU,E+VY:1,.>7O>CIAKDFc\
38OAHc^P.;^KeIM7KOGMPWFU-eO(MTL6AcI+93)BAKZFe4J7gUP<TY6#bWdeBaB;
YQU4gdOJb(W88Ra,Vg;eV@+aVP&P,ZCf?]8<,;?eeZ[AT7];C[7+bJSA6W[\ID+7
3>33];P><ZB2g=TTcSa3^/0#O.4:@.>4>;1@gQ2Q6.D5B+ZYSDFRF]2HEda?GN-2
e@(;HPKQSO6TcE)Z1a2,Y[PJ.4D:00\Y?F1<-J0,)/31IFQT)eL2U;ZdWM;+0RI-
-I\@>Jg=CO-2AT1G2I6>fS]65H>T+::b7CA^7UTAa.1^=7I(Vg/@Y:4EFW56WWKD
FR@K:0VFGOI,2-I2^/d3\^NH25c=28JcY>:]KII[(B>7AL\d4]5VLG]NPJe]g^TS
)^YG^<_8X+((a5+.<VYK^?6BB[U5_CB0V#:/SV_Lc7bFc-SH1DHRE#IGYeGgTeE[
6:[#CUU@6B/3#M&(\HFL7R,M@C5HCOO^:XEW4K#=.(SDf2G\[L@MZVXO@V@aCV=R
[QGPg&#RfL)K>OV-g\[WUX^R-gK>)APH>?L7aP(]HCCSQ+;bcTUR7LPAEU52SIV=
@,DN]@df4+N(:I-M<M]<O05dO,B>1=4>X(+>C8OUcT]\H6Ng:[UPIW[^KUD59;,&
IgG@fA8KN7FDfaBf&&7U500W:J[4/?OP<7#][<W:ZKC1I]<UW4/?B[>25IZ+@?eV
[T9S))ecH[8Z>eP.cE\&Y(445KM[,IJTW#5WBM([3cG\Y11HUG0IK<EQ3TTH\+7c
Fb&^@D2\.fPa,:^</\:&&f\JfZJg6[>1<7DPcK5dbAXa+0K^gaLeg+:0+M\Y41P0
[817<&fcfPX=@>>IZd&<S&SV.Ha6gWSQ[GEK[B]IJ1/:E)b&18]cNP2e1g6A=[),
.CUUTaF>GAf_\LY/2F_1b3bD#B&/&e0\LW^>eKJTQ>Sd<RdY(7fL#=IOFA7ae(^f
HfcMHc@D@.ETb(1A@,KH:V00Ae>@AdMU)b^b?Kf.Z[C]VO8VKAXd#=fb;C]=e820
&09C<FK:(3\d((4Y)^AcT,?V,Y(_W#g(:FBIb]C-4P0K(g>3/;a49e2KV?d7,X6?
AF>\#-Wdda(J+SQ&b/aaIH[HPG8J6YK+R+(=T]1UANTX7:]+a_#OdY1/).eT<4&\
]U0.ZJ@&3G3,+e8EN3C?D,+YEY^-]F^3bZ-25(#\>ZODfeH4-)PO&(GQ3\f-I1X(
1I_1]K:PCI]H=S&e3GL::=2#ea46)^L##ba4FR@GR=4FZ+B/bM<BAacKP1O]+c=5
C7,1F0dL4e-(IWII),5)X8J?Mb[cd>[7W)8RT(CD6bN_.^]-X9>O/-?;,FMLLeaQ
^c2K(UWGS@&ENWCWf8efb:IA9SG8LF(4g8d5f)R@@e(B_aNYZ2]MfF/7WZ]:L5P#
c=@8Ydg-:L?7&V+?/&=eGSQD8f&M9#Q@.Y&2Y:CgZe4^e(1]c?ccZPa703T;F53\
6LR(&X6[Ff#1e:?8U>F-:.gK(L7U\WC@3aTg6->/?BEL]TQFCXgK]-N08cNa<MNb
HBGVNcS>4X/I(C[R&5;P/H1_QSd5+U@,=:#(=[1C>XG\2WF9gF>_1HII(Q;N/5A9
I,BR7^2IVIJ<bD@P77dOM.]=JO4,Q2YO/b^84.[E<I0eQg:KR5+)0f.N9+K>c<(.
A:e@\&C]R[<+/Qd05U8U?TEFe.HH@MDM7OQ.X)UQ?<G&IPO<.:.^?(aQW@,_3[.P
,?7f=d=J)+CL5+-AeZZU_G7HOKHWV@Bb\)AV),>-NM8#Y1]Z/.&=cGA6]X(5C2b.
02<e(\1.NFRMC]e(,R6W#G@XL(PB>2a]A#)SB87Y(^A/361CH>:=8fQeA:SDfL_0
[Zg7MgX7X?<B#RAEI?30._[MJ?R_@WRG@UOdIGFEDS62b3P.G&8B5YYHQ4SR07:?
?,G/>E(>0V7(fI#T\S::3#8NeY(4-GCS(cEH6F5E,e[#;Ra^f?KO+3J#d6)aOBaK
=B^\IC^N66;FXdSMecD@UGVR@8@gcKRaI-V?=L.;^AX?Fb=^@bV/g+(IZKLB_)Ad
Xa:E.fXDE/++,c&UW)P\J/0:W&XQC]N#[AUC5b6TCIVX-TP&Xd,Q#?^8gfH7\CN@
REV>g.I\?:/3MH\4]7B8F6Se-HCS)2-+WC/[/NcX+Q0W.J&>L8].;=eLg)>LRYFM
STZ:2,c+.1c^8K)2=#C_1g5/IW\MKHE46B43B)SFbR34Fg4_20B@+YgURZ?70GX#
X^;()0e?Qa3KdA8F&[I5P@g5,O>@7\.WWG0d0HF\)92/J?@9\:M8@<?>,;JU:g0U
BVA)&.1]eY-X\&ABWdOBV0H_-=,_QTKT6UGdLI_9gA,>(=UU_TSHT8D>@Y?6Hee)
AA\:6]Z2+dR?42P&XL6YcC)9fbd5]g,/>LbA/cNHSI,W-:eX;Ng=\6)dBH-7<NO9
3U>TWR2P-3/SJF.c8/>aZ-T70@YL@D;7UU7Yc1(b5d:Lc@KG=1QDKK_K[EQ)&A_.
e&\4E:N=;ZIf;O:N\XCI>HGU[O:#[>HG]@0I>MUc(S9O?._6]\E;5>XQ,=]dJ3HT
1&@94VK-(>9Q->^Wa2E4bITe?,5F42Rd3\^=+c,EPB(\I:,5XH<[KM)=_S2N)4aE
+4U>4]Tc)D^WZdH([@W_<Wc\F\-J-QCY<&PfZD2]9bB]L+J&T<ca2[D4.,@07QbG
7B+-O6.T7&E5L5ZZQZ>2-f5IXL@4&016V3Ia=Rfbf-OKW3B8IGE7S6X[\F8fJ_f#
CG_D3Dc8.BULbCe(@?Q^Aa9[If?==5B1^,P<W/Bf7cfK9U+M?]OFT.eQ5)gD31+e
fHL4OXO_e+J</Z98.X/+7=<8d98#E3fX@fCKVR<S^#]H5G_9PY^g[(9Z;##^38HC
(WK7AJK[FIF5N8acAKQLJX6<TLKA(2S69;S&<-]PA5eW7@Bfa.<&F+95L#3G_J[+
ccZNL;=I?(&,#a0.E:1<?LE8ZX,,PW[[C:U,.JO\FO3XWZDJZ?B)GUdZ>c(3XZM&
2(X;IARX^GFf?Y/BTCNPgR7adD.4NZXP7[;TL2U6WFH\G-YE8Y3MZ2#0I8H)U]4)
B2WKZ2gP-0aKFR9^=3.-8aNLLTW&M(e\,#I-DG+W#.8J8FD[MW/;UHVYb<a0V^eW
?PB0MVV2.)A2ILZ12;WH1A[(43WM>V9TY??;b;[T\O4&DcH@fNL?F1/@gFdH6Z<a
=X:)FC\[;LVO&Z[6Tg9L4SE\[?PA<JIPPA[KKf#=I/ME#@]@Fg\7-2Pc2RXN5FHV
)eRbS0.@EFJX6O;3?N#=UggcUT3UR+Zaee#17d58ZB-<[H2V3Lf:S[Da.8=)IF#f
;P(4KZA,T::2T<A104adQfDc-\:)EXT\.FOR/DU^/(Q3b)@eJU(I>M<AC_[;0_,_
+>9)J.e0cYGQFd).[.C\;U>FaQ(R;CE#QU@f<WZb<Y&V:-aF<cYb]Q+6RC0?T:@)
8+C2IcF_LO/0XS.H9NGdJWE&.AYAgYI8e-()0c72a8>,,R5+KDYC=A.3&V&AD,1^
1>LUMPIf<d4(e0,BK8;\Y^2G&?c>/Wf7eSgJ4>V/0Fd5&11a=g^f=(91\+2,+4=a
LMb;.@VfYF2ORFbMO1D;7\dM[GG<1ga/d-/&(>g)_Nb^5N^O@VVK]<Vc#?DfV3:S
9O&1R?E3Y?.C]E+=5:6Vf2<LbM>)<M9>SOH/LX2,TXUO7\FM9IEFTQBOdeeW\XE&
dMWA]>A[c]YQ2cZ\MDOG)2][V<9VX&g17@#[YT/U>_.@=P\N3)RF].5KLgd)\_]M
J_5/W0;XQ5?1/S)PA>I)>041Og@4V5c&?;1?TMMg1&H?#(F8M)Y7TCI1BH)>#KN?
@g[NN,M5b_Ng^c/O(Yf#&)AH-[3G=LF/ANR06)D1D;?X90L)[_Pd+#@R6R]]a.T;
&5D&Y8aC:Q>>W0eF1e&Z2&0UCc/QS(NS)1UNaEE9P:,WLHW&BF3;YffMPS49-5)G
fL<JVaMW:6+=cA2,8N_-H3?G7^S(9)(S^-O105CA#\]IB2<-2b#V/[::E6P7C2B;
80[-]2P)231/5MBC-VH@_^5G3g?e#e[cfb:<7f5W-WE=-PH+Q11Y&b1B7eAII1B_
MPB1a>VL(Z=6CHe0@g#E41D9Q7O^IbNH4&_:Y88P]2HOW;E.R#^B/dGC17PI64gL
Peb>@YUd#c-3\XQLQ:SP;X6ZBb1?dPB?bMF6M/3F_dFA#:dQQ92\WJ3EA/U1@X-A
R\V2b?BHK8/(eOKFCVW_[LN.D+-8./@KB:/XECDY6H#ZOZ8RCP_@+PQc.b<c_6_8
AH@HG/_;S>UUPfUDg543bN,6Kc)JSI3O1G/38G9\WaG7.SbbG?WZ>VB<LV-89S?M
f=#8):U(_[gO;Z?L&7X,CKLf3bN#.Df9_/XN9ZDf99]P]_A#Q#KNK]:^H^6W&JKK
.[[ePUF6[&La:@a.[_-=G#Bg972OQXEQ:P<^e4UHFMEeGPBbM>7ZbA>8O9K1B/N:
7L]D(HL409@9cK8\8,[6_,EY;<b4T/A0X+UB9BL&QM7XKOL@I/[.8&)_MUHKYHTD
G#)K(@4(2B2X([D6S:?-gRRcEXJaR=6()7f[9,6;K]53FCd;,d9D=/f/-E.AAKg(
(\d.KP?ZTY.+QF22O+.FaT48d^IXZOHP-+Zf;Wg7-dDDb?;@gJE;HR@>GLN&[3&3
;f=c&+X9X0C74^f<^4<[7aR=?6D61HMCH730]/M_K2FHOMEW]J3/=?6=5@FgEU:?
DY,L[VK^FJQEW#[Y#J=R.E0BQEf/8&<F?9(&b:e:0\4JUT?GK.+=X@&[Af,1E6E:
OHKb+d5=AE6ZU+;:O/H310K]\)F_JC^dKAd7E>D1#e\^aZU5W0Og)b2c1YF)M^64
3P(GbMabF(&]A_:,Be3\FC_7W?ZE)DZIG7NPK/g.G<Mg@:F9Rg6T:gH.0.g1d(Y&
4D<1T=;/2fZ@;IQ,YSIgG9/cISGI7_c1ZJMVJda-BeQ:TV8GP6@cW=6U]W#JBZ]K
C1&#H5LXFCND[IaPLRA1PW\4PaKN(:\((N2]@G?JLC_28TRb?8MU7MT/YDAXN--J
KGQg\-2T=c4OAOCbGYS<&D)WQWABB=4+@(6MV;gGO@?DO&\L.GZNO]cf;L:We[V4
;T<gXD=VF>?bT_QcbI(HKS1+[W:RWEUEQ8.PVS[0c7V>8-Zg:F.^a<C@W42Ha@1B
_dDY<FD>K@L:;9L^:X+fU5HQ9#3]@]K@QR,.9QAW.d&M<gP^C4<e#.Z)^FVKc9@^
/Wc73]?/0dIWL2]G#1N/X8[]=J-9g9bWF;Z9.a:W+#0>,F;/g8b:1P<F<D@U(P0?
[L2Q?^\4UFbOXeK1Zb+IV]/KG_fTH)a],6gd,+4b4?+K,b0)2C@6)G&MY(Tb#LJ2
S[5]84RgADA^]O.]J_dQJ:D70URB78^3AL9b]64P.4(d8fXAH]1)](>#M6XQTN_I
)/A@aO@X3dObJZ:5JD9JcUabcJ[+R362R^P/eFRZV.DYaPICM-0^]D8dRe=CLeKW
565N?VP0S6cZ81O#]+2d-g#e]TSF5aa_+fOK/gc(NJVb^8aU^GG#92b6#VH\c-;X
T,ePO\b6g5PF<(,\KJ\BNUGf?cGX#/])<g/Rg:G(3K>>M#Z6J4I+@<f/Y++LaZ&A
.B:M&MY&-B5P^I22fT(+L[G_H@ded;XaHS=-M?KE)K-T&c-BOfVW3I#D-62f7=16
Xa/)A99f))L]39RS^gaNaT2Z@/<1d:8#dM5;T,e1PM.CDT-e9O4E2f+d.c.4<6Z)
-)2-PTTd/-969PL,f?I[=.bDe?d-];8;@PbY&&20Tdd_::=Kb+d\gLKg<\eF>;GR
1L;Q(M@8U/1EYeSV&&;GD-MO8?I8OE1]^b>_406D,.1(d]Q0+DBCGba&AMK9fD@V
/)R&]aV^I_HXI4e,fV<>GQ]RCI^[?82I)WXTO/g.gbFJ[IF7(938>EgI11SM9T_N
Y)KTMeC<:8H;LN@G8DF=NMP/aMD:9W\95@0TOK8-;(FZC2^AAAZJGD&0K:])YPNZ
[9SYdE0^=JOF9cSW.PZAM:KD?Hg&FU1+P2QbeaEc\:4S_[Ad<8N(T;HG<-YS-B>0
96aE/<ZS__b;L<#-)6#D]eEeAUMGEf)P[=/C+])/UegP79_E>2?SA>H;S41egfOT
_8NXY[EN>_FS+&4O&0?5Lc:9:6E_AGI[a&O54Y[)AQFDd,1V?H0Uf?406gF__B>W
00C^PFX<#GPTO>LeFK(JI.BZ.MYC(fY32IO.dHf)3DD;PgB4>N;624[<N?8eaII^
@.:M..:Td6YWG@UBQ_>_L,6AT_I+:DM#TBdDbRXdU?FY(H=CGL-.KP2E;dUCWc<;
a-HR5dXQJ?0LIcNP_/VKEA:1LX)<H=;Ie,e<ND-8((U<GWZ=8^;g,2EC<\]2B6Q-
,g1(F@WFBc5JE6#-FXeFf9ZH4J+MO94e#491^Y>3<&2#F+M#^D.&_Dga,7@0O8UB
Yb36_[+Q2_Q>OXQeM9GWUeFP3FW:Pd6-Zc;f1P_aMI4(41AGZ4:f(G<JB+efOGB3
7OUF,;A;.0gRP19B5]-,LT&a/84UdWf)Xa/?F8,C&6;3SX7U)D=RR@d#RJ]SDR^]
?)5Ka.N(,LEg5f:aOEZ^@6-QD+NfLOPg3J.aNET^ZKQ3&KP=e:5B+5VZ2OQA3NZb
c5.D6T(B#F+@DaPIa_bFK(I32JUcO@@P\_#U8/<&2BAJT74DcA-9ZD/PS^4Af)EV
PST520ZXPYN#H31HT^X/;6[cdaZSg1HGQ3SRB4[;S+O9)/X\+4C[^U^>a3)AC^JB
P_Hd=^S@B.RH/52:@E=AZ785R,34Eg>BPPGH7.Xe8MSGNBMP<W/RK4b:,,(a(d,.
37M-O=N6YKPMGg#FXeVRX4B]3ee7]_>P;.3:?VLW:_Mc._YfN;,RH7+[6e.KA]7g
,>?X/J?.B^5Bbd(Rcc1[E&)L-bT.N?R[92G3T_9\\.Ce:&9PEb<S;-,5f<^3:USQ
GI;gSL8>7W5V^^?Y/de#8;_N6ASD5+>L@[PWKVgYMDCE9(GE9_\D[FR_fM[+0X;d
MARY9:CH,GS>5S0#1,K>Q&(;VGNP42fW@X118g5N4FLDZ\=L/YRMe6fTI?DD,_DN
0T?#NbDI.]81,B9C#;(2:HW:0T-Pa.XU\4.)2Lg:+)2TC3:a1bDPId01-.dHB-A/
?UJAFE2Q<bYARdOL\BK_4.:HXZeD/2,G)28CeCc?#3e-\,-4g[-V47b96.b-)9WF
J:,FC?GY#+e\/F6a:[V10#a=&X4Xgb]UY&S=[[;9:DWeCVZ-33,B+c3(g6-5>&.-
UYYD.)F1M-Pfg4=W7]VUU+NF+<4;&BTGHHZ9P:I2,<FK-YL6VcGUL<[-UJ8(;/S8
<-&+974O<Y_AI;N/XFc_2&RcNGWRLPJRb]^3?U\2AAY6d6>0ZH3C(Ta;AD1,)AQW
[2LYUW1^+&QS(]CQ6:-GD(N=Oa^[N_-KOS3#>09Of;6d>BbdaM/cUF^aDF.AIfa4
J56AB[QD(#>RS6_U>g=OHV90?C./9;g.f/OYY<5#bP.>KUT\RTGgI6f>_MVW<VgC
f&#INA4VQKKBTPM4T7CR&OH_79//XR46QH<O41B)\BP1<8MZ6S/B+AI:Og(:0/@U
;5:RAEbJIW?G9R^#&c2XY^R77,MT(-VFE;BgCA,7Ef5c@_T&L:ZJD_e8=e+BJ3AY
6Ze?Xdd6B/?C,Y,2<=)_6:c5U]g9>caaEFf6EYb#(F8G-&#[DI2fgHG,DX5\J5Ic
LPeM4^ZfE6^OAd//&Z\V[MDVQcD&.X3FF]1D^&SY)?d6_F^\NSN:X]L,e^Z?1/>S
<fe>F^,C5bY+\X_Jc1?9VAE_MX.b+gX7ND]@=]_;FS/W)5_+8X(f/RaYOK3H7/G.
S^c6V02N[Z_G2dF<eLRVKW.?G=124B&#e0&-FX&d1T[M0J==2Y>XM+g65ROH_NDO
bJ#U<7?g5MJZ[9):J3CT[G=^QZ>YXHbcHHUF&Qc#(FI/SeS==4[&7d2I@[&a>_5U
<^P[KcJ[6/@&O:R4][Bea;)+TdDIEU#/8DH>CX?B(C+<3R=G5Z^\AXYN#&[R/ETb
P02?C7bWDOK;(W.OQPOE@^<:2)B/SL0\^A-<6^4<Ic:OTcQG7UR5?O,>@B(]XYFB
=b\K48Q)SEfWKV/gg5M:_=\KMW4S[Y1(?EHX3BCZ0QaTPR9IG-R^TXb=9b-Jc-?7
G)(U^K9#>5>7VS,]0#N(YN^3(J],/>,S6[I^I#R@4/5@1:3^@/H&TUdG0N5I>b,4
T50:E5C[:TO@MGOC/]O/?&deDM+W]]]b>O>b;XcbdLS1,U/-/(<]WZ<fGXIJ32^D
,9Ob4bHC1ff;TN7.3-Q@V)LcJZUd9J39?E3/_HMAT>1QW/K[e[KM(ET&/OUeYK#2
@aUU\9]J2RTFcgR31G^2VF=,/ab_YQKeVU^R;6]S\D]Uce699.D3GL\WL293CA6C
[HSE3TCXdda=U7aA)\?c,6G96gM],,.77^,[V5If>3I&K=#-.ag)+GgP=-T6Tcc^
eEfR)TM>VfADD7Ud@E:,#<d=&M,9;<?W,X.V6bM>J]Y9POXf[E4>6VQH7LJB_3=,
;gc343P8\f5>/]I<X?@9dT-bS)>Lg[&6WE>._9gCS,IZTT9NP(394;B4b)a2[Z(M
eaD8FL9dL1CKa+6C&E4)ACagff1_X\L5:5;-bMT(H02a6De8CYeN?1GDO9\0fO9Q
Hd6b:4SAcfM&AK;T>G0G;H=FIa[P^.#XfJW1#9dc7GXd/c.d+<Q@_V9+b?5aMH3=
=J,3U)_IcH15)f0G,LN;Fc>A)T&FgLVcS&O8L;76,^R2/MNA</9S(fXXd\)>[+YZ
MfA)O?F-AT[2E4-a7f9;aPbb#@:<D/2R\YV@<Hc4M)#BOC]SLVUHP4a^?L/P00J&
ADL[O-OL,cAa]F48^6;Ad4[f?ccX1_]JRC3+9Q6RML+M=>/_]_2,=O]cUJT>VSWO
#)@PK^ag37D_+_.[Ma<R(8#\)OYeg?dWV7S>-CN#9=b>9N5_gPU=SCEdXU3T_-W[
+A+M3A<VgW<OA?/E/OL[8_62.d_=NAL)4ASg4d;aS+O,?(J7e9dc+X=86,f;HEI\
Mc_66A\-LV5?LTO\&F.2C3T2NU08C/B[/Z[QW;_9;OIQU+4&JEG6>C0G2@Z4dDG/
)>FKX-H@b:;._Q#g=<_C??)?#)\+a:\GaJ.PID/c./BJ;00Ba-5RT</+APR.D9@_
JG()+aL?IQ[cA?@=;_KSD-c8EC&>9D=S-L7ZYeE+\Q\D<JQd[+LF+HfA.7/e?N^7
#IO:?Y:S-M)S8SS(0bY&cT?SeL,?6GZ8f;Ff7e4/dX17V7X=@K.bQ2FadT.SV-Q:
NG[\a_YJNP-&9#<+WA)\Vd9CIFFXP<>_PSN6X2f-]K54J=?HR,:ce.D\L,C7=8U-
U@>ffV)UZZX/ReY35f<[T[<C.AScQRFHRNFf[a[;=.U;Q^9W#g8USX\93S&aR)O.
BX7,Wc,Kf@aQK_L6UgA_7YU:@:;A_.Q=C7LBNf(>>==1DPd?5K>(8RWR;<\T1C(@
VQ>+aJ9I]9H.[R#HYNP&</.,RLJ2dHUBCDI,FPS[MP62a7/IIU?ICSaFQ1e)&ELB
:0]:baHG&D\9_Q/JJN?[D5Jd\2H#P[\GT_K633[R#:,,Z3W//YIaJd3bZ48X?+XU
]fgH(DUBGbce/<C^J#3P.R#CX#-HE(TENA;I81\fBbV3ceP=E4aJbR4#I5\fU5E0
76H/D^?Y9)[);ZMW&\NO04U/GS:CN,WP)=H,Mg9R3PUaF37C8De06NQ[R40E6f]_
0KPLYW3cAW_A/[?g/S)GURM0IB?TEcL5>12=+KIFVX4,9d:.BT5Ea5L/D18BZ)]N
fZ2+Z(\f5I26d&_eA0SE7YP;[[G+UN<,E-ee_80@:K81_JDEP3G7BZ(SgI^gQI=^
]UB<3MX;WOgH>Q&4A/BH_^WY[A8NL@,b]CDI0X4G1JWYbMP:LD)6GgD\LM1,M^e?
[BeCAPU\dY8.IJEE6Q@C?A^/^U@O9F_<ASBJFec@9?(MBa76W9@S6+OgRQQHff\J
DFXO?J/a2XLa8I)_e8(G>F.Y1YP796DXeM2Y[HgVCIY,,LKYH_?ZOSVeX=1(V#V#
dC\0[^/IPJ[NN^;SV@1J:7B<NbS+,>ZTX@bU=4Pd3Y#GLS9Z^8>W:7R@>G)>0Z_B
e]OK[^ReW?OJXc@>@dV>O1YbX<):JPX8^_?HcYSH,29<DbYd/B1eL__ESDZQU-WI
\DAe4f^K7&/CRXQC>+U-2f;T.9gfRc7>/LX8BK(Pf01A^.56\_JD0XTCETDbYSLb
)IPA4JJ)B0W.,IdfQHA;P\b2(.@L_[RDW>6&J,7#O4-O.AcTHQA^@Z[TLO\IOc,[
]X[eB7-X\[Dad)?2N?#;RV<HQ+-E/4=VX,bM9dIPXccIB<TD9AE(W<721J8eQ)M8
d[?B)_ET+MLE@J=AbUHRFWd+G](6#R14=/R&_C(IA?.daddH(@)#00?\I.XJ0M-C
&HJf08;cHXeQ5R3)1OBIe;Tf)DWI+O2A3BWc<<5A\9MCP_HY.dQKBZ]Oc9Ab<5W7
5Ee82H\M)>HdMd5V;NJ/aN?gPdBAFe&QC=/D_[f?^-==:.>aMP^+N3:T0b[c27DL
CHBe1UTGF.D[=EFXW1Ie7<.@10O5G5]faB..fX.WW04b(T.a,bRbSXL9P8S/O0I6
+W:YDFXB>6/>1\IDNA7RX<N4<cGE32\g/=\QSgOAd>1Eg[#.gIQd62e(;>fEgN<R
W.OSN.+d,2=M29G5WP&Zbea^Q5BRP6]aI;[Q+J=e^S\C=73P8TG>O.UEG17<XHM5
<R;58C.S@LK\2>9PF)]EJ+/U(-C1-aWQ6U2b7X.acYcPW1KI+cP1#XY9bNI?C5-F
0WL.QBCP/&/DaGXE8dHfP)?UC#-IF94QF\NN_&SUY.GLFLEb4:,L7/V<.H1K-9)N
/QG5c@RO4VIM&R]b^^E1WQaZ^)R[G4c\V)\\YGE^bb82b\;E:UN?AC+a:G[N;8H7
+V^]ggFaRDZ\.W)K.WL,(6#V_&XO74UL8Vg:>gEJQNM)K/JM8U5dR\7-K3U)PDF.
7ed5^B3a4&=/A\<Lc[FNX_(64?^A&dH/I<aL@3b<XPc#1-LP2P2^Z:NADbA6Ca(@
JOO>bH8,G2fXIAJ,]7MO9>U97>@FffC:b6;>FgXX\,^-:;F<[2G]<dQ]W?,5#>LH
c7FgYVE8?a-5C>M3YTB4cc[X_.@\?7,5JNg#\3V&HYX>?1=f3JP5&7=])+D9d/=B
?]X6UNVB.)U;8VVBQfc(7VQ3ALUV5Td0eF.0QV]6bf>bNU7+6B]HY.8=]9Ff-EdN
Wa^OMN9<6+9[X7RU5;8cB6NFRQAI@EB/D288?@X>PVJWY]32E5YdFH4H,1cXX2.f
LO31FCK26/;F9^20JJM+]+#9A;+>^_FQDYKI&Ya;_A--T[>Z;4A@+O)Y\=4T7+Jb
33)1_RX0+dZ#1g=)B96>OQ;=aG1-(,K1#^g[US7FcPQUJY(#5411PC)<F7b0?#<\
12<>HGdWT)4DSHH680gEG#e/HRV)F=a@=B?O)<Y[(-RJ>)fIG]Q5X-.TAedYW;Lc
8cFe3=^/>^&E=)0/)?,d20)4PFEUe:/H^bcX:cSY_L?_F2JF\S&_O&2S<dT?6#g6
[2KgUGVP\R?A_@^4><TK@.X48UD2);V9RMILNI50US].8+&-AGf@4G<;b7e[e3E7
Ibd7;AU_.P7,)b0HfO7,.W7STUJJ@_:Z_HLKZ.H/cIAH8:_gG7-e7+V,@5P><IQD
4](QN\=<90(X2A[+gWID7.GeBg,[WKQ/6W#5A;K68bRc/O44X7:UQ+YI[f,(f304
d</KLNK/GdK_86.+AS1AIJ44;.:b0Q8X\94RPD^G<<<_Z@PF:47gRa@<5<ca(+YZ
K(;1)81=I#&B4?#&,:T&[3#>\dLX10e7/NXLNgH>?49c@W^7/3I++gW0:S[.?I]&
d(GDZbFCO?LTPHFG&)dHGL\FE,H?VGFV)AP1[YY?O&gdgA_(,EQ=1cPTXfV=RPPC
:@g[P0\AbP]&NK&SSO=Y_]G/eK218,PLfSdHDeB_[:X+9QObQ_IUJ?@N53?Jf_=1
@]e06+R68-=D4;&fd^69DP[T<S.><T3W+C2+&;)H4S@KWWV435UCOBVJHJf7Ge+Q
.;J8OEE+OV\&M+?1V?@FF,;JMgbFQfXFM8+-b2X=U1UgAP1FdPK(NaS=1R;LH#P)
0+B,AV+IgSF97g3R=X&bD&CH_FR@:;Wg83BUI,\D/@O@^d\:WE089@aPAZVDQec_
47+@3\IQcYBC@YCc2/(@X>CR^;-/E4-XefS?HQWU9+QU1ND_P7Y_0;+XV7S-_?M:
41E4XXSacId01WeY-XH+3#CH@26FCa9.47e1/R_QMdc<M9MbYD8K1W_@8U8@BGO(
)K=a8dTAI>?)B6[JN:(VD:caF4;R@JJ/NfdKO,W21IGS/RcY5cNC]BW@1@@/\dA=
(5LK6T>#N:d&e(Q<SB85HTD259XOI;AYCeVE52-)HUO<@<83N^^^Me:ZP9[6LaH:
N\LEFe1(\]##H@0Q#0,;IVg/V8Z<,_AQB&@B9HfZ?eP8Yb]dQ=NQ]gA?A0.0bF](
1U[C.CX[J#WdLV<DM&^=dSc2#\GL)QZa#DFabR5A&(e)\WM2AUGBFL3;>P.cHfY,
00J-dO?_08)>94APQGRL:b6>GP^25.EB<fR_C1)6RPd>-PR;7BNR:6(DYND-_BPE
V>>U)-d;#3.+:L\a)CE&@E]/B:TFV7#L940UF30:TN:VU5^>g0.Z_+5,eJU3?KQ2
EKV57STO7_DG.<bfWPCd.]PA>8,J.KOW3_G_5/CcM9V@8KA6_Z\#CA&3ORf=>&6E
@<RX_W.7?_M^9N0Ad9,91egTfdYd&&DZ^_GdWNX7a1,&b01C4]L&TZG.MBLJX80f
@=&3IY^ZMdWAc^F6_\(8DRgRJ2?;#YN=QFJC.G1<^[OFd0V33E/[g6dHeEZS122E
@fH#P+VAN9R1Yg1T>V.&D/^.K\;+)eL)_3;9R@L4_,R_GVG/c+5JfT@^G=5&DaK9
3bGTQ;)^ZJ.)]#^:@fLd:(Q<&B^fJ.RP1agZ8FP^=KC[]T31)3TTg@c^dM,K6e#1
)AfPIbJ4IdA8G8,KA25RUDS;_[cV?Laac+@=AA#f^[NKMSLWF4/?[HJVH/=a\(-:
-g]D@:c&)K^_-4Y>\1RJWbQ#2CWZ]0gFETQ1.G-+-7e5^J6FcH9KG9KNHfLAD_B3
@d64c_FU/=9+8(/>(B-e93X>A8A^PJDf[#c.1WS;-BGKP7f#K,@-C+KD;U(21B0;
R=e#,>,X#aTFUC?>g+(/@L.=XEVY&Ag/WIAR>RcOF;_+^4]8)E3QO:\_KO_?eTH5
8)Q)S8M+0gJP0#5daJ)P?ZcWNR3U2QfbV<.B6[B=LK6fZX(N;0f^0RfXgY2PeR)#
19R_0C?I)>YL6gXRO30e&#[,2<KLPN9\KCfXVA6:AX_I9a?/Q<Q\a9MTY(1;W1?#
YUDAf1_X</aWg+7-eF1>>8TJE3VL<JVe-CBHLDUOH_;aIU&(6U-Gac]HWLfZDXM[
HI@S.-)fJaKN]5K4SUYFJ4IR5[b^CI.FD](L).87^^g^fHRBK_M,7JR)e,]U]TGF
W)@?)&P]-QFCU2K\=:W0:WcaE(c@]<Q(]HW&]a/30Xa/OM?C@^gAFEWQT4?F&:/c
GD#+>E-N\]=,.O\LV.d2D136ICE,)1V1HN.5KGIF2AUJ.D+2Jgb]#Fb5XT0#B;D#
5CI4C__AE?MPKMIfVQ3;]bI(MUNN\c-FN<P:YK55?5=Lb7=P9<HSN6:8<bXcT4V3
Rb&\\YJdG&PIJJ=d:E9TE\;8^4?,;W:a>9g^X>b5HNQEe7X2=OKL:F_@26a57MZe
[[7c\?46N_]I6<;4GO)^._8dDWg=YXIH_J+P0[@FU:)<M1<VGY3^-aNVMfe54?-^
99e@@b+@EafR&ZFT3F<+;-&+W?-O;(>7^J&GG]#M<fJ7[_8<V^Q=QPCG)1,bK0e7
O3P6\YJ(-Fb+NgE2&8YTY>cg7[DZ;SEQ;Y[^f(89NMC5I2eabQ.M<\)ST+-BFAB(
CZ;@K\NSK3,UYcVVC@TP7BHHD8&3#;#&4a\dVa@7DgVeG9\CY/b?PWf0.GOQMT10
W]_5#,0N0-bFRK^f@470#@4;H;@-D1)VG;b4aE=U71W28ZV6@K,N(=)M2D@O>O[d
;6?g[(G_KVb:/OeWF,9GJdc@9^Q3Ne3#]GN1XZFe]g4BNY@W9M]NCS098/)A_)VT
.UFZHc7_Wea-SMY\5:W@T&DEJ:B>6d^g5K&Y4g<3L+1:+7]8FaPX^(Y&+#,CZ68Q
D\>_I1T2D]M6b>,H9\AC59LH:Y6HWgRT-PEeV<cM_?aUG]SCUd45bWR;^3_d=&CX
4;;Y^B\PNM8M@J?^<(Ib(SPFNIG3#.5&EB#DVGYU8_M3)=6eecMKL?G7AHaJ54(f
<;UA.:+[.e2;3dITd?L]BaM[8)34F)&NZ60b-7aPQU1<8Y6cH^;=>JJ,D\=5.?H7
Q;6[H9DR5RZW5OM/[6=)S]MSVG,A-BW0fV@da11>,4C:+dO<RMcDI2/@fMJ)L?Q6
V-YQX1VVf/CZ>[c,aEN6Y3P?&;U^?fKMF#6[T7?7M->L,R\@XdU+&S\c/J3b:_M.
:aWS_R[<5[6&Z+0Pd7f8=-J.,_3dD&LC;A:>O\K-=G6E-KH2VZcH-L>-YAb1\LOO
6T@4-.2>9=7Q5P9&)/Z#-PG&8BHB\.X(cCCI_4OL-JB95g:3QLWW,Za?.I_WA>KC
5W0PHc2J+;eF9</VRE9I^1e[D1S)0Z&I5EZSdA+X;6^M3=P>2,=.7fJ@SK,3,6F7
SC<VN2VKaCDX^R1#CM;aE[\Y]M4dO7_.XB,Y8AMdI][\b#/JFZaRUW^]]?(G+a84
W1XR.T[#K75C&?SJFX7_6a27e;[D#GEb/IR+c,3TdB5NGd1fKB/C[cFU7EOb2U0B
H9?HNNA37W54(N:fE/gI(]]+NL9IAa704C1=VH9<T(-2XU1K&>&VB-H)8-9VV_H]
?gZHA-6\8(.GSW[W03Y?9#D)UR3CfgKEPNL_:.ZF?PL.8W/T&H>P\A)#+/:0J0>8
4Tc&F70GQ[IJ)OT]CNg=0^@+b#3-4g;:O8QI-)7)6g;A6SP5+TdbG_\^WXaVVQ3,
-PAdUX-DS78(XaSH\(Z]D;<FJH0E\L544[7J9E\8967cO(c8#@Z.__bS)YFEUf8@
STS?5GVJLFV0?AJHCHce@\9KP,4H\49/6CI#59ZK)^K9Jf#8gLI4TMc8dP<F7TQ8
4XWDb&J&OD\3\/0WVS\LbFI<G(8,B(E^3G<5]Y(.Q8N7(_\E6A(:28Q<WVd<6IAa
SfC3_=KG^fV8C<E7=8O@aW2+RW8f6G@:=((0=N:WRfQ9eFbfT4DQ8^Q&d_C.9>,[
HGeF4SLZHY;e#W1UY876-3P+OSFQ6TY(.&?(]W0N/;9A)99XIc;PCV1@)+0CKKDc
#fC2[D=Z2[d+gf))<\721gPF#1:ZaWIMCdd>5X]=OL87:+QJUZa;Y^gED>1(/?93
b34_FX(?B62C8(U]-.^J)(e4A;]6>68I\:Idg8;V-06(ZI=HC[&)++0N#@3YC4))
,AB]c:DBfF;&<1+@gB)\^\15KE9]#UW<>:(g6&=INf<HHH\ODAH]f4c4]5]W&R[V
3ENVb>KQb9Q4K>Wb6b<YIcLZ?1[]NS@+6JYe]S<EITQg9cLT<AWP7SIROBTgTb.c
MSQ))[+BD+:5TO@fD60]69<GZPNE/^JS@MgcaYQ;f+4\gG>TR][;^S&Fe4/aLCKE
)@,181FZGe&-fQgZZETfZDcbFX\\_2<=4724>_QLgRE?VCQ@#.[JaKU&EEY(caWV
.J_,YUa:]VJ3e8SbB/:]A@E2bGISb+-YAED).EUDRU([d@8J<>_PU8JP.&W]6S.1
9WZ_K0a8V?2]9?d&Rd9dVM2N;A4[gLc?c,0EUWV#?PCa:&\f.HP<#M.?G_:[8^]a
P0c#_DCfGMXH3V.R:(50WC7.M,LWU+IV)>8A^+aN2[S5I0<M/MIf#Q34Bf(1^B0G
I9ga<KW0AM\>/RO_b,JEES?S[.R:QI##R/>Md]Td(CeP5,SG31B7GH8,531&)=1>
ZaW[cJWeELQBYd_E7^A3RLXWHN(4[5(H6N6\KIRdKQQWSa8\F2^FZUg^9XDG4KB;
T:5.#<W7;,1_c6dE/PJMBgL/7F/HeP;gW@J8.?#_965ebFKWI4TS\X7Mg)LGGQ+.
(K^I(^gg[8,4c^3&gS@FIOZ>JAgGPO/2RJ&&[bWY/3]<F6g37AYMC9D4L-@ATHB0
b3/59g,JH)+]E;_(&&U&6X>.UN1NNc<,V?c?U^2]MJg60=T77b0;#ead3RdgCF9,
2Gf[6DaU,-](VW57#)?BPedV+O3a;K?[17=2P-OBU8J(dO&J)eZ<\fGG1CP;Sc<F
RF=AVIOaR(^/7CXVRBA_^H0If3888MFAXQ.]>K#@2[f38EgS>KeF7@\cUN&02AXH
P>N:C<M1UB(H4b7N)J[)D#Da-SO>/C-Jgbb97V^>__K/QY.Q6#PX;b3;0P[M0]1_
ceaV(R5J2[aXBPCP=Egb=HOKSW[O7fPf(Ob^;]]3X-F?a0=5G=U,CHA-a]aPM8C3
54,Y_aUJbc[F^D\W:8)b^VLLeJZ&2DVW\7C;J7#8cf[<T&[^^>9TbGFW#d\XVHJK
RL^4g(&:6BQH)?0S1D=NW.&.(AW<_[0c)/T\]LSAJb\;a+d4;JM^M[3\:<dT+K5(
#>5_OB_<f[Y5HV/a]<[cBH#7D6CUVSfUCK,?RWD1)Efb?3<bLUV,]:Ue85N-M<O]
XG(]d:>T4_#_XB+-eN5D/RV.>=RJdML3B/K1B^ScES3R\,DE48N8+9[bY@6@Y3=1
Lc^dJ#F&1#IXMJCU/^abDc=5Z],5\B@X4N(B/f<&/;]EK<L;H_1W2cS&g^?+I26@
4?U8/(_#N,/)HQ4C3g0Q=[<;b^f7M:@VFP(..,--JMCLcW&:G88OgeG+PCC.JOO3
?V_:AeVY,D6XZgT52\JQ<#L0VDJ8^R48LbUI+ISU?ARL3JAe4I.0dK<IYd<,U5DJ
QV(2GK9@.X1)JCb].gC:KUMNL#b;NP1?Bde:BBJaA4PI:R<:=,Vc;)G_E;#>:adg
MW&gC2FNf7+I-QAM\\EDcb?TOZ6SWZ0>P:f<bH,#6=TG31H)d./;=QdR\I&RQScW
a<]UeO^3fAc&D#^#=Y>Rg-aH@93SfM1Of:aE:TG@Gd);PEOQ67EIO]KI]Ya:4ZHH
2XG8f^C:d8(.1UaM&e_KYJX<gZTH5M@L+5:06;OJW]=G@MU<7B_K/&<5;RB&c\ZT
YM17=<1HW)CRQ#IL<S6E-RTaA<ZC<A@EC9EA@U_d@QX8.(QAI\].>TDBObQ@(fS3
R,<bI560E-Kc2O&WR,@b#K8A>16DM#6)XLeWM=G\KUVXO1P&3[0:M_:c<,[8aX9T
Z<GgZ6g/F6FI,>eT2V]Nde<6HNdAV]ZFW_I&W:Ibf&:e?,ULCX70b\]0XDRS?TEJ
?.YIAMNfV\Y;J@7CHHKIMC70PVOA<PFQ=JTSN>WLV;B3</5)?VOMH3Z3LdS=Ff2F
@A[X\EPDSJ_?#\aaJfC1\ID+G1,-dC^&)329+6FF#X2]a]6=M76XR@4ANc),c)=Q
bA]82bQ.Md6+O/G>e,+a[[6ebR].?DJ:aK2ZQ9L;@<>MP,g_T/Xb4bQRdIg<XAJ4
8<[)SZSgK,dIHB.eT7Jcb@1@#_7\=QF[N-J6Q@EDE_V9YYOdCG;f_35,]I==:L>1
Jdef9Wd+a)fd73W<+&G2]Z(;D+3:B986&OSIF.;3N]B&2OK1GbFX3gG0PEY?DNC/
0RY6ZK^gB/Y6Zg32Q+5TP+N->V[O&[H.d#)U,fGc9QD]8#5,MH5?[)2PS>;?C.Qg
_Ted@=7T:R?#RdI:cDNY/E#.(MUMa[X/(dF\L\X0^U42Sa4?\+gRPI>>^_@c[-XC
[&Z3MG:#<YC1#L(#B06\-QeX^=ONY?O3TT77L-21XKb7d&fL_79D&ABDYWA.K38>
AR:gQd42PS\FbQJ8bUc;UFO>OKG5]-Eb#4ONK^Y>Q(S1AO5#O52M9>R2_E0PKbBE
T]cBNgf=B<W@g=&41eGCC33),Afb<+B7/S74NR0:\,>,_<FZ#J;H?6e8,NL/&g(P
fdZ)EMc-f-^]C;&=/W:8g;K/[H;JMM./LaF9?W<R^IX9WUPf?7[\G?TMCMX]ecJB
6)68P(Z8#4A#QF,eCADY@F<AfP<^G&KbICG^eGK=_De7UIfX6d8)+FD)gaX&)4,K
c02+]WQa\>VF:@E:S/A&0TN#/0:/e8^UKD2Zc?D<YKaQME>(J[RH#CUC\1>Z-6MM
[O@V#c&gIUGW7@O<G@(KcVMU0bEF+5dXXHU<ECIXF;,Sd&8,[+.M1G?[LcORVGJ5
MD\C[([?(+9^f+Q04_OJD,:2P0bII:/0ePG_@IK+4cWUXY?J;6TM-RZL9JLK\aXW
_12YT3+Q)Be.V3=/,FTP^c+J3/B8KAYN_WJSK]=3,]TKUQB=&M;0=EFI0g2R#47-
^\[O#?MHAY.]\AfY7\PD+fg36F=@A:95N2HdcT+QLd6K@deF7CffV;:3&6^XJ9\_
0<5XN+dCXH[;4dHc7@04_]?RScHEb?8<P^>PJD&;OTgeM-AU6+.U+)ZWa+C75UPf
HNA5^DIQ)XR7\6d#a:fKY_#3Q]_?)bfK,B>(U=Ia4TS>S/+S@SCeAXSPOE3,Ob-+
^J<b;e/D)fOB&+P(FOMC1F:JQc6S^cD,+0)e#SB?2=cV?L5N)U^[bQK22ZWZ#IK=
CL^4a=7LdKXOS6c]Y1LPe[Q1gc[PW_4<DA77(#f0:Ac<D6,N0HC^;K<acMHX\\P8
fF/\44[G4H_U._6,LOe\;LUKPS.<84FX[PULNXDJ9AN/YaP3HF>]8FX63JD-=5eI
[SUD1fSQDS/?D4a)QFA;>&VC#&U-Z3=XXZW2ZC//=[.O2aY1UO91MCL7[b@KG?3(
QT-2JRZ1RNf_Y/R#=5Z\PH_R/S.;5,=N=_HJ7HN876\H(c:_0gKS4EV=F/a\b]33
?^IUY-VeSP;KSX(XS5A@#<W+3dE2O0d.A8(5<C]6aSS;(HZ@G)8>NM?CfY3S_9_<
8Mab0EU&BK?>)BI_3:U\.\VXUTFO[EdUKV)L&K&_RA::J>fAF4#+STM;>JVR)^36
OdMOVWc-H_8E3(A,YWJMG5c&3F2TGKQT-.ATNN2QUZWN;eBL0?G#H(,FUed4bRB4
aE11Sdfc,\.\ZSfceZN-eU+<P3Fc[[9:T8fH-9)I)@+E0J_(_#FEYSCUH6c>Of-:
-=H\fNQZA9V0a3&NK?d0CB#fR2\>C(=U3)WJAdVDY6fD]GR)CeA&=)9KW\F>g8@-
RSD[NJc,/G#Z5ZI\B1LVL)#.?M4B.F38+)M?0V[1PBR;TM9,;]eK<8C</R#;)>Ra
LbS>4a6RNcQ:&>J,7;JPEYe&4F]\OGU?@+/NIT[d=WAD7.=D@,+J)>M0/\J@=V_G
PD>BeCf]A=?#a(WZE5[2NTSM>=c8/<ZI=Ve2ddV-DEK^a=#D/e=cgUJY@bY7H#C.
SI/aRT39DgF,TEP7a&A9,^P3\7W>,ZeYTF>#J(Z::N)SaZa2.bMB</D6EdI;4YNQ
H<R?+)AU_Hd2RI_2bAOGZQ^RF95A;3+?V)LUB_#L4Z?Q&)BBK^8CSB8>Y6c+e^cX
[UH;bMJ9RQ;#4@MX5=989&_4N-RQ\K69QKEZIM2-&1[T9F3fZ8Y72G[ZbJIW_Nb(
3&AXad<6+C\7LW]06QVdPKBGAeL&<3e^FFD+LVN<8FbP/K0dZaUWLBZ-04O-DM-P
3BD3)GHRKQf.\;c2ORCS]UKeRE?A2BNC:Sf4CMc^C2MF6HACgDHXa/J=<[&HYgda
Q@3]>R&]V[:47)TS6U36<5(OFD/BIec@JZZg<<X&e#/a]8/g<I06_YK5@VfSe1bd
F>bLC_TXCO)\DfbA,=aO7JR?+ddA[&(LOQJU/BB4TdH(CL;#&e9NI5C0Mg>egfE.
/CF]+U_P(Ja(9HTfcY9;.VJ,&d]bE<dA+T1(UeeWV>\>SBM:LeGD/[PEP3E5T^AW
8Z3XOZ2.]=G76).@:(]4>8N\Oa&RA?7P[b6_S3d@:I/&XGL+2a,:NL0+M2CG84@6
^3HJ6(HT=V2&UA[40M6&<WTId=M.P#AUKC=D>BQ7>+SY:TIJ+gL)\0JSd4ET)>Xd
#@AI76X(WVSKS1SaOBOf(,IBN_d,BO2]6YYd)XNTdT=L18S((EX3LbE<9O1,9B;4
cGV4?3CX3bW-CWd0]+9UZWg#b^2V=RAX+[=-c3TdNLXJddcaa(N[aU8K3474YV+X
[LQ.TGSbE6+^#OJV=XaVKZeK>MLEUe;]/&6S=)CG3:e7(eU;Q\G1K/+;YE.A59cd
6XJHI0&7g?8IF\,U-:9JVTQ74MAJ[g;3--<eC67ef=_a)1Ob\+(,B6VaF/>T]8P0
Q<IH3H&K\cU;1N>K#Vace:V?86.,2O<1?..24A2#//=3R7_/&Dba-2^+eMbdL_Qf
eL-RO&7Q\c&aN&HHDe5HV2KK?QTDJX9+N]O+Jf>]&F:RPUPCM-ARE8aY,_P<S0d9
S9KFCR\P6FeVVNL&^_DH/61=4]ba+]fMebSK1;e:XI3U8@A+L(YIf^aTKUf5e>WI
/&M+5M6I?P=LG6(dM3+[&49e)S2:c=05;>_.F<^a\Ld;983T#b@I7B4:U.98;#QK
>aHWR#&[>F^1_\GQNQaZ6A:T8;ZHf^DG-dGHYP=caKTS#cRS=V2B+OHB(];C_[6E
&E^e=1^g.VfO;K\7RdN(([SRYG\cI)HdSCbb.,+&K5+22O)/@L8^=fK[J.C(E#92
FEAXU#d_2CYZc#/?9EK\F1G?]3C3PNI4]IKCY/9T7fUVTSOG&;&=7[&DW\9BTfZ^
X(ZbDT,@LPS#1+BcFU?5RE9&LddPW4HK6C^0V584)4\2QAedA<Z59/c:G<OGGX=F
>3(1e&O+V:+X6bf1.0F<\V-NfS1T?EIF;aWRA+=I=RJeb-]H2K_SO,73.LH_20IG
1RAF]@D@\G2&3NJ8)[>TWe<cMNRLNZfZ:3\edQSJ.+#ecA:CKbQ(E56,F3^9MdZ4
>8JQ]a_8\PHE,U6]<IR8PdG-?=DB(,6&RQZ3/I:PMN_CT2d7,9G.\+]1P3U\2a#N
b?G3f^RGG#H9,AB)&\2UeFdFeE7RG-&:?-L-#.YJ-g52^+)\.[,cQ5>bc+;)F?,O
>Fe.1>>67:UbZ^fMDK_/L[P<XB7]G5aJIPVY/BK1[>9@]DYX_S4P5SQ3JQ62b:\<
HF1>S+GbZFAIDC<9A)KGe=O]\5ERf9/PfWDIWWB511:X]U(UGf6P_VH/DE6;#W?S
&8ZB,0CaN#eZZLDE0Z]&EA(d7YZ(OD.J<.VUR/1=H.)+OOd@=1WSbCe1E@?=V^#T
)FFUeI:;Sa-I/?.M<;:_,@<FE1.4N/fWW#.f[\RMFY6,VSP_0.WCaMgS]<[bEV(Y
#>M8#aX4ZA(AEAAWC(FE5XYf<H/6#Vd5?6d?f\7]OX/:d/_4;f19V0FBX[VXJ;.+
gdZ[0a8=Na(V_+GWR9&+H7EU:\HAc\TeHUGO2322@Ob,5;.[+6)62,I@SFMV.bZE
dSYJK47B3HY,VV>dMUc7a#YXfbNDU[<&5NMV_a?3KJKgGS#UZY6b0XfJ2^>f3F<=
eUPR&.<50#O/#GOS1A=\FM5,cJF_3CXdU?;Q\NG5F+K8c^);]7GF&#.>Gd76fTc_
0B+J[-LV5S^_<8f@_X1X=#MUMf.1CW+2@1&M?HTb?gTRZ=?2-[C8HC[2&DEWHKME
A7MgY)Je?fZ-ZE\A391KEAce/2bP/2Z?DN=#,5JTZQMT[AEe^.P-dg#)10c&=]Dg
CX6TB(]9g1_UG#K9+a>KY&@Qg1LJbcXT0QdN[2N.XWP14a(c-@,>@QI<D#0T&(F<
;1L#UV6J@4T)DB.:Z-MUEUI&4b9337,1E8c>=1&e[f646aG55F4SQR0F9^HY<FXS
;I-]=95RV]d,\;##^&.==@K.(0;3XCD6CeG3Q+:2R3ac.WaWX<TUA?TYV\I?6&-e
XgQ)2PJ5=.67L36Ne#R=S6B+3LbRH4)><2GKe):cc1bEe^:9aZBc.U_QQYKZ)1_Q
M5Q>4X<G9U)K&]b)_#;>.^;0UH5KHBO_W0\/S:SOdU8f[S;98B\QWSH&R9_ge;WA
21F&=PNH<@35YYNL>Z(/)CSJMDZY5_F-=aCXM6BFEG@Q4-^F)4\5?^,>U/P?67VH
M=;_\9\gXWgN[:3JAF[c:42HP/0QW7HHD^:6JT#PO(B2RY/e]Y9Ge/cL/>/\5M/Z
=SW^K;c#Rc\\&T_RQ)Z_85&J_^P/A7.Qb-O>(87.c2_T@S5MMK7UG3&Lg4X5YM(N
eadB]B5d#\?/UNYD]:M)?YG^W?XWQP(Z]:(9<WA-J9Q1b;N=d@Pe=gHJI&\P/AQ6
S-Bf(cL;Z@)>eVP;I9aV^>c4cVWaXJ#5TbDRGQ:XfNJBgc>ALVGJJ(A=P;U-?B3B
O;8(g<f-D6&cd/G_7dZId9NDCcK]Q[0I:XROf(8XeDfU\X76/e.YIf18N.KZ<[_I
F=ga5GD9:TUT_dL\,d7(=He\^Xg:HYd_7PCDAVD5aS?2&#+-E=YYHYdAN8/C6AY@
=6T?bCWWYIbbO7cd2/:Z3EeDQB0S1QQ(\VU<fUgQfYU2:-OVD=&a@c?;-]fFGD4Z
g2U:[8gcJ6-H6N&@6U:a.4e+#R<B;ZR&#W4++c7/a[3cS:@8BQeOGU3,PX2<2fT@
gUYL4U3]Q601BfPHK_^W_(&WJ=S99VBZ,7W=_bYK<L/;HYP,&L[,K_3FDT22(L[S
[UTdX3A)^_)9KN[QMab&(CD\f=8b9Ogb]^GVe#0A:YM21;c^Fb.(8#[+?D.Z,S:Y
P,PROa?6bZ_gIfP3TH_>3GU3G?E\:]._E4VE=d])X\?B/Z82dUSG]M]56F:29JN8
TKP3_1;P03cJ)VW^P]SS5W;.-\HeZQPgMXO<)]YOb\B8[B@,\W134X/e+^.WZ(G\
3@9@e#ed14,79dW\0-:?D)\H>CG[?Gf:6GbHOO/S+2G5FM[CQQ1(VKE=&\8/+JRV
>&gMPMGLCYfQ#70I^0e2L?V_,:B3^DWSE\F6De8\&a.\N2FWQ;b&CfFRZSG7>ccF
@GBM>e2;DI<2O2>].>M(U:R&F<XDg4GT/1\Z^eR7B==gW6_ZJ;;N6Mf;/K94MWOA
G[fLf+]=]e+D)B6&#6aI:NEI:H1KA?bM\T/Y)T3HBU\\-=S01/?=&SMW]1H00:#J
9YJ6NafYFf6^,b(K#9-:>MfC(HW>B2^;Y5>[JHY(=U?L1FS)fYEVBb>&37:#W6J3
WMARTI:7NG@\fBXTaCT\W_P0D:T4eX(0\eH#^5/cg=N[6Ng7VK1beLR^WU1Ibg7K
3V,M+5CE)MB2GLHWY=\&WLTE4E4:GPCUQ<a+KSc7J/cI:[4Z+b69,Y5#Zcf5g27>
a7SSQ_0.DNG52<UX4?-f[E;O]aaB3E?(@//,V6414T@^U3+TMf;7^L.GJe[UUY#C
L0Q,TLH.EUT8PaV@aB^dDgEITCW8+=T?cN7[I46=(CDa([-]DBYLE5Q)R[PU>b(7
W;B#3#T+2;S0^RN7]RP2c#<bTLO1[#bXZ#H/IfA6/8g.;SD8EBCCBGAcG2(f_=+;
)e2dBLg(:I87SA3H<&bV&X8_1@PZ@;1R?)Z^W(E,4OQ9N[K\d5KW7\KGOXILdb[Y
LT]>0=.BYa+b+b/M_6(=^[/[G>Z58=+?gK-+NW-O)Y7CaDDaK>[K:1,Y[(e7ERY,
++PLA_Z4^J.6+XKNQDS_YWM0?RNTPBC[W@<_1g889/I9AP-JG6aH.ca5U3OSMYWR
XQ[;)_?##TSOSFWK8-1#SMHZ+0T>QCb9X(291T85e]&<13B@1I@RZ,T65T?dT>]8
BA#.=dTG=Z3IS^;);Z2KVV-#V.X9K0GAKIBY?Y>1g#1O=5V>FE]@^Ea3V\-Q.,P(
,P@0=ZP[F8#GTQ3FcUdZ\F>f0=[dPfKJLZ2]\<KM<9BQR4&6>\b#W#8K2gX-V)HH
\>HA.UN594EF:d9[8aVB10gGQ04-fR:MdSA)^=Y;U/VST]g[]>>K?5\]VXfUV+=+
GAQE^/ORG6S5cJ:MHXNbaK+WZN?(1=Y_aCJ#-7G,Q/C52.bOM<I[e4M-X:g^:KA=
YWO+@)4JCN>@I6+53eL)?RGF1)9+:;I-cUE-[VRJ155g][#Y/\eC35[?G&Z-_,aI
<+UVXSeV3ILYc-4-4aB2OT\ON)K[?],f.QVLgWB&=1+:Q-W9+JULD][1/e@2(8-N
=_ZU014L_4K^/A>=1@?\M)<7_=g#<[6+Qg12,Y_d.0V),aZMFXd0)b2e+#?HAF<V
L9>BKa8=b?:SC?OO;0RDcB>&MKN@)-M5c,CDIU\d=:Jb95DY1/[-DA_^.,aLW-]Z
gF0LS6NaaXIS3Lg)aAWaO1MaS5a(6R2,@:<Va[cIf>03U;>62/2ML..[W:IVf7/X
-3T5L+,CU2>@?OWJEfYJ\b\f,HKeNR^]aa/7S:aA\(b+C=-Z18gK?A#dQU8bE7BU
6D7gKR6[CBRf:bJ>Ka3L6,X<ROeVd(6^cbTgIb_^<2@;f/J,@I2:A(^-7XJIZe]B
>?S2,U.4@<HHOP(58Q^[SSP5LQM4:5MGD7))79YfdVC(PFc_-&WXG+)J8<=W&UTS
/IGc1Q-M.f8\=FL]F;(AcJTd]#3L_6),NOX>3H_V<d]cJREXS6@?CMXA?a5KGJ.:
Q6#DXG54BSD<?]MD0M9926_?3)YYfNUZQ4S]4JVW_bI0CBCbCAZ8.#L](bdC5VCS
gVcYY4_-e)S8WVIg(AaYX362&g34I<g-Q,g8M11/c:)W@\HHW[?OO;)0U:ag7WXc
Bf&]6D[OPcE8;PF))H]K[6?SG_JTAP<S\^RJ(aaMBgP]S@>+.0\0a0L(+NQ;UbAY
SG2:RQ#I..I^G^?&.BaLF&KM_0<B6Oe_P])[Z:QcA>6-9J4.&U6OXbf.?IN)ZGHR
@/B[+Y]8V/5IWKDKdc:7I(MG@,)V+3)QEH^/QeWaKA>f5W[-E,H[L\E-&Z26Q/][
H?E+WRE>/3LL>?WIZYUCV/8YJ)VO/F2)/G?UcfEPf>Q>)e,8O;95./=B.M03SIE^
DB(LCgENZBS9O(Ve[K)#8+cQK.BF75<X=U/)5cBBI)?^PMJV(#ga+P3SUCV0]DJX
1YM_N_eMd(;V8H.T-1U,H>B.60K5VP=H)3F360=VMLXWdOI(58Jb#NO;EM\SO9fb
B([C;A0T@,BJ,#)&dQY&<;\],.(T5R[c/5MOLEJ@0=]EJRe;H]8YPZXCW7D364G+
DP->T7U,W/.3e.-dD#Sc[42[fGR\6dYbU^GMaN,Qf,XdQ]bWLTe]>YP/4RNGGPI7
O[SRTGF_L)QaM)b,C=Q=B\KcY??H45[5<b3W6DFETU/G93-4Je5D=5V;I^/X?^ZK
]acUU49>1gVBa^]Aa6/E/(X77L]PD3:,cT+5H+P)<Q#Ba^WD21G@L801MR77)F#R
LgVeX[d@dbH#17X,@U2PEG,+WMQWG-BYDR8<IL;NI=&3-=FCB#JAZF=LBe,b;4)H
<)=34_]1fUYYR(2>PdJC=bM[<TNV?YSDTb;a8JY2/:;)<:#3ZL.(81(.H]a>Y9T+
FCY46S)V^]PdOA39KHO)2J[KX=BQ,:Y=cM1E>&X3D1;b>7L9_AX.:^T=SYOHJAe?
g2fAH\95G]\e6?XH@ZI/@GcZeAS=+;FbTbO^3/EYEb3.7W/\HOcbTRMHNfWTeWe\
_^B]3U-ZNL,H00D;e2CI0^2J8THE.NLIeCAeeFJO4/BgbJbX?FaSa+MXTW\RT7ab
aK)?6F=Ba#H8IWX-1[8G5A+IJ/XQOKGb):6/CQD<KG<O;I/&I?2N>d#[C/5f\AOQ
F5+LQIE2_8fWB[(,>U.[Q3e)[PIN>XOf2.BA9G)G&.#dXKT>&QQO,4g;E5,CIYG;
7Q]E[W0:8G7>>GU]bY[U@9WA]c68^#eGKTDCPM^\:fITd-cM<U<MLA3S=4Vf;=(Z
1(Y)^9a[daNY^+>36\=T<?87?:SE,;]>M4?P5\70]NZ+@9a,QJ&4fONbE.[\N4e\
_FCLa+XO&eVHB#)Zb;3IP2J-Vd/SeSE-\RV/MI)?D5+#K_H6Y.1fS#+7;fg-RF+8
\_+ASXPa;/\UJSKFb&BZT@GUQGDg:Q(VZ[Z/YR&Z]>a5UaJ/g?H1\Dc?09dg7b&H
7]Q0F([:Fa6LGX,)TPV?0f>.P/8?b_QUK,^)L:_dd9;&f;Hb5UT>JaK+GVV^[=/1
N6GQ3:39GP7HHM^VP/(YD5Z8IPYNZWMGF:-+QZRJ/F]F_O9.O-I?U&-8e0<9O[gG
65UVBQZ[d^HQdC4I/JTBQMdA+#NHT7+]2>^g.<VZRR1;O^d]PMK,B))<\H(D1]a9
dLFM1-bPW;XA:RU.LA)Wbd#[KcNM_/2&3](PI=c)_)?fR1DGbO/SSLH19MS]UJc_
5a]N&B[eUf)S3\8]I\Hc;&LA8[:3T,#42/H<EY\)TdX>bR4]^MWD[;8C:3]RE6O:
b?Yed?,2(TZH/1:TcONLBUg8I:+&]M>R:db#YUHaUE.Pdb<4L0<dJ-V?0Y^L-BWP
V6c[(;-KCCUX<HLVWTeJIC[CAD@G(QAX<\,E+=NM:][A,E^W&P>13@)+^e+J^c87
#@dD?<04VDZ10>OA<a5_UD]V<Y>4[BQ8TY)6g6[6&dEHUdQI>FOKUS);@M;SGKC[
>)YH3?5TCcY-G5G2WQ@U,JR@J6_Y+/Tf6g<)CBNXQ_QLJD@Qc0&R@g]W+R(WS>>I
X3A\:M&6YDCf1ZfGXg)=fH9f.Z1#^XSIY-N?bKc813G3-<13^b<A9>?H<;A3XM[F
B?D6PXd)Ef@F;:1YWUOR-522:+KD814QL+[QJ;JA=KSNAS]8J5-Y0),g3bT&b?\f
+JC1b,)4B[PH?NJQCDC9)50L<-[ed8<<+aUI_#Z/#S1&?J._X[HI6LA/3U@_DRXY
DO_AR;K0SZ4X3G9U&0NUFg@EP6C;JA(#Z6E&R)1YQH)5NQ?GdS,Z0>de<TKT4bW]
>@g8,cXTT^_e8HADN/KBYCd#bY6-7M2W-XEY&W_JFXDQP&8K6AS5c[3/8ge,IID>
R26+DJc1@[EHT?89E8J3DL4P#?QK>7e2B.J,-.02O\T)S<E&Q/S(dgCVZOU,(QcJ
\C1=6CI)da_=@).WE9JW4JHaPcVZN4+N)H3]S><W/+SGO_XBHL+7[CD,SI=OaN<M
#+H.TQEW]H,0PI-M5?\Ce+63EUAVYWL(,6(RA#_?a,N1O;RO-YdE2W&8LgHH780[
FBT(Aa]3BT(JbV8/M4aBcSINed((=7W0-bf-Bb&4:9CWAX)-e&cKUbL)cLFHPa\X
M@6-\=XAHX:N\ONW<)YCcE&?VIZ;I@8M,AYLHPE#;^caefg,)(_\d81ZRf^HfZVS
aU=7R9MXa;KWTTO46X<X1IATJJFE7@g2X@fAQJDa6[Cc(E?.,\FdK.1Qe#3[Q:AI
7</I.Z)G[O,=a#K#=;:CWf&CGSBVX@ZRYA_[g1=S/OD))?K=e#QX3gW+PIZfbRF;
Y34M2e&&H\Q^ZR7;@<FAPP5UA98V?-@^MB;P4R=(a&DPP(3N7J\BbWHF[V1D9c^U
U6Ge,[MS1Bf@I5cAe#BgcA]1U&<B=)?.7UFZ4Qa0U>\A-XaT;4Uf1@RfO-_Hb49E
F5/ZfAPC+,^<\N=.CAI&GM8KXUVc^S12_a:D#)gb-YKSZU_W=Y?YPEAg^D.Z-O<T
F]L0@9N[#If^)(\]&9<Y2WKR5BAUQ-[(&5K(A7E/7E4K@PefWYHS=QDXZ]J[G(d8
\#IaT)d5-;8/8-R1Ob+UcM=7:\JSa#6Z1U2cJ:9O9)LBX-X9K>DMGF]0T_ACgc?[
F2T4+CE/KMXOTZ:8N9T6(I[Y_T@CEAVV(PQc=&JN/C=H.OaJ0Q4;5Z96:,H:^GTR
a_>LZaG_.]=H[DNO0R+9+Y\>G/I==eG.W]@1KcBC;.O2F5__BYA^..#WI#02Z:L7
:.7>a-8]9)Ce7Q/PU2\ACHfdL9?d7=C5-@bE]0Fcc#\0_6R&\U:\+SOZf>5Z1M/4
80.EOT;P^SQD;S1YWN7O_>YG[23_I6J12J:X/(9Z@RWM^gB;@RARF96,4Cdc)/M,
RE27AFIWHa.H8F].U-.1G]]D2@I+P#7C?M9b_S[Lc8ZF+ag:\(ZDbM)+/DReR@P/
TS6(;6=;Q,2@S>:6;gK]\=+=Z5LL242Le24C2[<adFGZU9Y9?ZPgcC)e5gZS6@ZT
6.g??3+K8?R4(<INGg9<SWSU<>^56BZ\cW>+.Z:^JYZ@4-H^>\)@W\W^8ASX6QZe
<N=RB^@>D8OQ3@(aCS(M236W>Vd&@1[9[9g8ZC:G8\XCNV,Q&ZF@#0X34]gXC3,e
[PW^PH2T/W0e^MX9O=WL[0/QBXTM1W]B8g=N/SA]2)AX/&DCQXg./+69PE.362\.
=Ud^?V/?M^.6URDf:?E>4WI\C.K(,I[RZb=)-0V7&a63[E[=GYG7RH(42YJ,AMG2
f[gY1WR7Y]Y2/IM(gddM@8F#SN1/D&^F?YY]O?GP#9=3[DANTH3W:Y/SF0\]>gG=
fgLcBYO[,P@>>=:SHM[&;^<0:^@8Qc)HSBg^eXT9_?.B=&]54QFA]SXc#8ecdO9K
UYDF/A^G0U4=@/02]9>A;H@b_3OV;GPDg(1V(29V<1O&4W?F7>=:-(ZKY@C(G@QX
Q&NURU:f(EQ0bZ2.>===F5bSH>dZ-VYDS(cYG<7MLR+[FF26&M/Fd;>.]4KNb<(O
WMR<DTW+++H/.d[6>RacP+5P.J/0\:WgA.;V(8V0dBPeF]VN-QMJfP5BS9P&2V^W
YTL#@WDWH=a+GCWCQ&EOH?cd032:?9T]DP#89+&AgN6^G]Pc4/3>2Je-YDD6?JZ0
c=KbV;bBD73G2TMZX,be8egC,;^L0)IYF&dJZKOLS]EJ,T(BOPDD1Qg\&[;A4<V[
XcW-U5LT\SEKB-X6d6aWCVeVSP,)Mc>(#ZfR2gN>_I#RfD^)N(.PM05((bJ75P64
A[^MP.O2X7^<[Gd@<d4T0^_V0>SIPPVJ8O[_.&>]#Z,O7a[a@U]RKf<Z73H=dGY6
[?Z&+65\^[QX1TF^NLUgX\+^a2H<fAJ5B^F6eE6KWV>JFH;0OZ@-Q]DaRFN8K,W0
IbHDLa7\22d+O51_,R_d#_g/B9TLHV#bN8X]^AAWg=G^?9OR\ca;RB4PdOa@JLP)
LV(_46cH7C=CfJT:NN()YI672/D3[3ae(,2=LG0UdLVad\U:;beZ3B9S=LO3:3bF
d:WeZ)cbDIGbPL?E2GfYJ;Cda-A,4@1U7M,^/eb1a-eSf>F3e^&@<PU9/9I=<&d\
EJIZC\?=S#\ca,64=[4#K>^fd5/EL/CF-81e^6:;S<2:#E#-LNF7_Ye<_6UW6SbX
HE&5Y;+gNYd?(=(Rf2J0WB6(S2/+E<GV_9g)(c#Q_8?<D(L+e4M(T@?EB(>&XG3[
?QOGW/B3:8>dY/FK09KX#XJF7V.T.cA-;8B8-CcP+Eb:e8DN.>6TF5.UM_a6-Pe@
;=<4IC]0X^^5Ud\A-Dd[C@7:A1afJ.#IW07?Ffc&C7\,S?b2cQ^50Hg=YWO.K3PJ
(a&M0<,H3(;aC?3YFG3.WP19EKZe-(16S2.<C:8YA_UaCM9/3/\TUPQV;TW#2=3;
U#-T0\R_WV:6#0?LPE.7J64UaJ-e=PC2]X3F=7=fGAeU2VU+8D::7RWTdAPH_[4P
)[A)ENbO0+ff?9U)XP_T>4V<b0W5L>,.B,E76-.8]c>&1VC3B_[LND-,9<.P,PNM
>R9,X.)(A7SO8B7)>0H,>.[S4+A]4=(]+^>MH/.\15S;\]4DT73EO)@G/2<>V8Cf
eFg(8-5)a7acJ?DO#d-\;O60HMd,Y;bNUd,6RIb24Sa&5S)Kd&c91R]/,(@YF_#a
4gFg/bc3fA9-a\3aWb+0ZUK<KEM_eUfCce3_H,^HV:HgOG@:0WeO,?bJ@<7>XPW?
I8WbDg@N1^9F#f:(cB)8+=^+PO91H=3Qd#e.GJSd0[e/_])RGKYV11f\==RO30OD
QW_M=WN^?1POcSGd8T1)1D?C&P=^)UH9E=gB[)VXB:=V\-A);C=U?JfSaL&<YZAC
)]9V5+\E9O&\3JI[@ERTQBSC/KFG+,(aA:#M,:F:0DQSG.H&2aR4I<f]]a8Q]UXG
B)b)Ma0?[#fS3VPI^D<^)F4SeY[BGX2fKEYR?ZA>?YDB,MT)QW##3.DIW-DW^?&1
,DOXJX:,=>[6GIN&IC>Xg)HIH7^O3\90QWHA#0[#5D0JHaN/;KV#_bS>]gF&>QR-
C2RU0#F?T2F[M.:e,F&&W9R#+JR1F(N4-T#1AAd_<O>XeV^J1S?\JL1M1RG&EY1>
KXV8aM&Z/ceR<22ZJ/&4]3>#)<cb8S=:E.GT6WJ>]1YE^KXbJ@X?F_L@W#0B2@cC
IH8[UgBd5TZE3\/.4a]&WC54QbbK9-)DKJNCPQcKG=3c:T0?QN@6T9[97/8=RQJZ
TgEK;6e=Q<?b=TKI=9[KE:#0^dP8SX^g:JEJ/3HU,,bW/G3g.\Zb7EFSc0LA/HBA
/f)@<LH]+JFMbBeg\PPLFQ2\RC#a\.([U1R5OO1W,).]MYfQZ)aAPS?aH&+C:Q-\
\@,VJ>3]_O2aG4/B:FN7Q38.,#?1PAeaY?f+T31:#[dZggbcK5W>U[S\)(?b]fY)
.WLBSCZ0cNH@Pee\-#TPaOgS2D1?TZNOB0BSX/9H=K35+A0F-Db@_IeSbW]@#UK\
_3>Pe,4DaD;[M)R;?-B9gR5K+&PL3;YN@.F:]F[L?B5&eIP<V=J-Fe+CJQ;5Ee72
DZ4HFaD)NOTDT5Rd7[K=J==6@+B2:0U]6:P&M,e5c@.+f[c=>3a.M+VNQ^I1,Sg0
;J457Y)+HP=Cd\EMfA_d9N#Z<9b/6JDJ;BK])^V((13C_XZfPbG3IX1>#D&<b8-W
VNPM=@TDN2gM/@58d[A>N:-_g#A.O-[P2?gd]1-0KKIL<<BZVJYO=dHfBK0.BfE]
XYPU.JSN[GT-cLZ#L2f^b770Z9]89=5S.OGCW/.7C2&TdGAc_>-J5O3=-=,e@N<\
fNbK7R;T08+V/c+&VP;,]:+KVN63#Y=6J=C\-B+G1KD68&86CAQc>13dHMS]H;[R
W79\cEVT^PcR:3P:R)LO8Vb=S-WLT:V,0\J;,FMEdO+cX[c4^OL.-]d.KRgE-LQ-
\\Y41/VXMZ7OZ.(]\3<PA?#W7_.e_]LMeZ9V/#-46Nc.MII9DNR+UV6^E5CVG[Bb
H\,)P.I+c@Ab4<Q5M5^830<MN(dP)DNX9X=e>L0bI?D6,&(eJ[@:;6A5P=(/O7gI
3/21UB[]^G60\5:B53Fba.Ze-,([>)K,6#EBSUTLT(3<egd29V0#W>Z5FB1FPJ(C
@3_EcS5B?C50b9c<gW0B/S(HI;CT9UcBYLP52bQ,MA-\2e8AQY=DXD/L_PYR&X/c
6DQSPUU54^?NZM7BY\U8bA7?3)<b^O][Q.LEL(#-PU0U&O)XHH:;VI,R:g8NK]e[
NA6bJ.9b5aTJ6PcTY+cR8@\</V@?-AP7OU(eOeSe6B)4N[KfSI6Cd\\T#NEL86U>
/C=K\04N,(V29E-CFG:/HS9Uc?J/A&_II.CWWB8V+XDE-=?XfAA]g\10&TR3@[;_
RZ/&NBJE-.1\4C]\\7[27C)/5JHM)<Q3A:4LZ,M9G(F.9=YF_D38N[5@\XA:FK2@
gb>XX@ACc^)CGLbgb&;Fg]\4#.OFVPa?c9X>X1Id>+Cc=ZVP3WSI46_9ea;OOFS>
:T1;3PZ7B/_S:c28NWgaB1fKL,#d1ga;W:U>H^,=C]fT[,LWg\bWBdQ>EAae+R,2
cZF8Y)M.U0IOTS9,QFA\C7de8U[dFVR:S^,;bNQbfT50)O(CSY(A(MRW4.K,eNY7
_OcH62T7H[SK07,@O+Bg;S98gZ.f-MHOD0^_CLXOS(#B4+X)^V_.Q5/_/D.\N-ED
aU;bEL3PSXDE,#6327(A-+:d>0G-,M?>A?:Ea0^FGaR:7VG^Ocd]XASf1H#2?\U4
O02::.XB1ICQA\0,?/GS+4VG=&2;;T9UDf-#VefD.K9gV129H6b?eMd0YG;FIES<
\F/[@]EWI_Z\[5;7]Y[]DMY&K:Pe6LIK/ZJDG5Q)F@F_=C^afd(aNYAHIH1M>&1/
1517[)PKF?/DX9;=V2AcI>_EO1A4<F<CGLCZKV+2D8+E&F<JWXM9;,>-)/4<XM<L
N3Z,&I=-e.eSKCU6=aF:<#)L9N,NE6/1<9.,ZgF3RQP.=8A66\_#LC4TT.[^fZgb
6Y(1HZ-^-LO+:5DX1NP\6Aa[Z5DC;2f43A8V1]SCc3J-SS@Y5A>N3L[0/<J;_S\/
a(W5&[85c&\TJ:&T/G&)^JEYAf#G#PJ?8V+7FC&(D>bdVdY]>I5248]g26B[5=@N
9]ZP@Y6^HeN@E=Y_S<8\>,bUN0T[P7.OV,U5>E(_EDR8-IS5<97bRd+@f2X[[04I
EaF_Gf0^U)X,3XW>E]6PBJ6X,g2A@-ZIfI:2P,IM&ObP[3L7/?T7&CM8:CMa90>I
T8,#H]39K3+T8SM:N9OabI+4:#L-NQY?EUX-TC64AOXK=D[I^RHFg)D8(KeSDM-]
A.CF;.B89K];L?C8;#OK0BE]/EDd#-b,?(E_XIM+EKLcW7-YAaQ78)g:HHO,G^<V
_&,-C>H1SWLZg.Z/b02VK4BdDOMD:bZO^LF#LAR<\\L72C3:>5g11_9K9BCZbIMH
@V/=7<SX02gAWWOfVU/A8=T;+e,]&Y?;/5TX@61#W1@5e)Td[VW/6/#WY]TE3G&E
R<b3gU3NWfAULKOTU[>XaAcJJ=+F4e1g(S(D&.AW/PfQIUAePE=ADOW\)C4(M@&d
GMJ<.3GfGF04(YDCPdC=/&&8Q=D8Q;)6?+/;DB?Pb1([bH7XVd5>YYX?\AfH2P_6
H@d/_I(IR9dg(a7)(RH3=(]-eC,889;IGdH3CC6DAcP-YEK^d#,\ag,81bT[<HN)
::N57b><e^FRN?:91Q=.CJ;Y6A00K;gA@KE21]A#D;/WcAOS=QZYCJd32E7SQI@0
#EY<;NRDg(T@7^fL4RMVOaRUT<EOUXb\<1A,\O0A9c3)A<QYOc>6?#S1J+8ZRB7a
7>,fg6-<0<@0#M6E(C?0/(.U^Y4fFH.b-C+HLJ(W\25PUIC8,>)V7>DMPJ-Y_>_F
f<I?9Ye6M]Rdc[E3aVbHdL-Hc5ZZfZ(<0UB?\9^UI5GL-VT&51:Z#WXSGF7H9WA#
0ZB:N]]b7?[A3K1L1HN53QI>KFU<:L,R]>^IE2]]&b4O\>_-+eWK#RLA1T.L6:S.
>Y]3\ONa>e,0[Sd]>/F/GB2_O0B^/fWf>F=/(II3Q4+M2B4=F_;,@#WdP#?/_UQC
^9aLLW-8W727Ne?dRM(5,5&W+(GA^=R#RK/^3+?3LA-aa:&WfYC(+Oc)2>V^XRTd
d[GB0.f@Ve<a2[A>EF:Re<X@FJ8XC524+ALE&TRN7dA;:4gRO62F:BF,6>D[eFX/
b:HSfE1^:EMZ?LFIF2U/c)UV#[:Q\7cKT^>fKX8#Jc:1VbQX-HTSV)K6PRNf>V#R
IF=KF?ca3Z9.ZM[3:0b(VYcU0X-SYK(4aHS0<@FZVN7eTW9ZY9Y4/L\>HE9L2b4)
@)[+RZ06\-]JFg,CDL1OZb4=+1E\@bHX7[Df3O7MU:Q6TY0[0N&0R54]Fd0;4-+Q
e>9Ec?3?^7KQH6MEEL^HOPP>5<#O-e^H7)-N0T_X76eeM9M?_D227?WFSa8BY=d^
X373TCY\+[FA7g(OL3Of;VD/Y153;TM^2C87ff)OVQZH2VZP=Hd.B0-?2,E-HBTH
-6U;=X17E+0KH3ZA\#3Jb?\<]NEHbKXX3CJRHTPbg^_&O?G4g4.7,,O+Ng],]J^,
=(E^C@T\UV(?P5E6)8Q;bXNJD=Jc&1;LGd>#FEA8OaJG11/_82WWe@(@K=,7N?_P
;0#/E(aV_c;<1IR9^5,(c(<W0?a3GHQ+LUOf>,)/a7We<8@T@4((2)P;Q=b)?edM
Y-8RS.P(]I+G>NcSB:UAZ[W&HbcdZaQI&ASLN@-:0\)\57>E@C@#^98>OL-6+AAV
M+/-GafOKLNZ2e=L#V8<X582R0?6Y&QY3VM^8-)LY+GDeL#fgOCS&2VUaK)L=X:<
8O8Q&=PLfF(A[&[DgA?@>Mf]NR7KDe:FRD-04+b>Fg&KcIe2[Q;3ION](1I)c60d
=(AZ#,6P4]ZH)9cHDZE/BK8Z=9e1e3Vf@DPcX<3F=&.@=+>ZA]@E.g>JX80/[+(e
a:O](.WNP4-\a<Be+;[^,-LV6FB8]_C&N9-C9gNQ0?T3/ER<L.B#9:]3P41;8MZ,
TYH_U<\Q@7]ISe-MdH\SLL#>\)b6J=1)/9[S:A\\./AT3MJLJ2gZICPMCB>#2eW7
?Pg)eH#0=M(Y[+g65V0#:6X#2KAFF21(.)WHV#,=88Z)#HLUF\>eeK?YC[JSSN?@
UD):#E[I/FW44f0^2H,NP?_;>aTd_9.agH)9-.Y7=Q(OC[2?Y>4NG]<SH^c?a/-.
+&)0[RfT^K_\(T_[U0HC6W8bU2KF_DbWVBW&>_2VCDKg@L^^;KNL:IfA_\@G7ICc
.&WL(aWU,<H^S0LGYLI_ZRCWgfA[fSG#PI)(HEABW-K<PSK<LG#:76.;B]\)F4eD
O)Y1g77GJcI<14GSIL@a@\W:1W\VP5TbB)N.DR6^@VD25BY;WM5e,PB[ZT@,_Y35
QGde0_<J:4(bI,O@FKfRW-,5C<L5[cWK(X7QT>c0,]:(6aD,)@c0/YbbVg7-17/1
cAX<1Y@:Se7X>a5bQQ>4A5&789)4QKdLeA9/1-e8^Bdf_AZ_+634b8I]H=_ES8<f
;Db_^eR6XAW1>D:\_TFRG6?c[#c1T_CK+O^6GLWgC<HO5C8KURSBLec#SP&H:3]e
g2<:T]49IBF,0OW.<GdM+=>0eR/c]+\^)/^-5K&^OP@1]4Qe(K8bFV(TeO0IJ^>Y
>.\aX^(;T;)5Of6KOFbda&FVTM99C&+?=,.V51d0^5HW+1=aZZW.CAcdd#<P4^I+
^gA^Fb=99Ta9X[c5SaH)>BX3A.KP#WGRJOWKSH]fBKVefc)M]8?4O[JJZL#I59d/
4+&f5_C726+ef;QEX(^aHdFTW)(-9EgBK:bD-KPPI;/72HTdON=(E[E:Ag]\R]2_
be4.O+X@cZLVR[A4_S??#?JfaT7MYfS./67ZSKaYOXZEJMRN7eJ^1,.);LTMP#Hg
&3264AV6]B5D/-W\8JRGbbI6JK>d+gQbZB#FQ6NJ9BdFI-9BV3O7LfU)=CZ=)7Ce
\8/_TPE[[L>G;a]S5S-N+1M?ee:&Z5+OETIf78:Fa>W)<3,fcf,1\X_-b#bT-_>>
O35-XgF:YR5f_E9D3FE[K=F5gK>](#1_)HT1K\])OO\P@:f(7f>,Q682g3QLGTY5
GSHX;dB5aU60X4EA+ATXTGaRO_aJK?]e,D;YJP?CY+;8=5+<L_(WHe[)0b(X(ZgG
MQS3b]+X(B/]&J?.-PRR^^A<193^W3)Mg+SO(/J,\(IH^:LgSUf2Q4[6[D\,&E?9
.MPKPKD8gW?=1QUaRW<#7[C/W0[eN<FQE9bS5S8U/KEcUGNF3:PJBLO9M23@F2]+
:CbA9G)dfL.Y0/Q5CA=X.BB2gHMM:89I/MZR:(NWDDW0@&,FHcP5b#Z/cQGGD(/>
B(+KY.SRS@T;d8#dbJ2GW5UH-_:CF_SM(1GE@RNN_R0a2K;U:ge=1OS_&,dJ1-\\
-\S+:/XLSQUWb87-LU[gVJ<cY\,dR##\)K3L3gLM+Fb9T9:O;H2RH@+@<WKYEa]\
5eQGc/O\H9Z=<ILDc<+URZ;H4G0O1DC_SB1[BD^CMJG62b-E8)+32Pa=,@eeR<.;
\3c&-SLH(P^BI#c;FgGQURZV@KJ8-9<AH@GfgTBaQbR>F(2a?]EPeK_RE_JYM7BT
NZSGL<dYKX&fO_C+BGGe\>4_[1FJK0.Qede2V9FW2D\73F7U5gF,&NE:(J#C74[.
UKA8^X7bg;UU\-fbT0MEWaSd_5b>Z3N<@6S.7)\c8\MfL[PcAfD5IS<G_U.GJZ5,
X@a^Z4^)TD?6#KN;DZ)@9\_42@B71LGK\@baE8UFd<D89I,R.5f4]T=I+/-S0)c;
Q=?COLH=#:P#5HI\\>C<<0Gd2,X)&Z)(Z=^K>dAD:=1XO.A:(bA;g+O095cKcF_Q
</\WCgf@dd.8[ZS/gLD&1P?>?@.S42P(?HedCcTY<@<PWRY/:BCE+/NSD89S^+A;
YJ1X2/>Ve;1@O#bGD4DfTO+<8A?.KfQf>c?6Q>E9PC.BH#<a^EZb7SPRa&6[e^^+
4,[WLGN#4UdVF(GV>ZK?EK>QTdH:E]+SA)ZG##4-.K)@dJB^97N\#?]NdGUWU#?F
6gd\9)g_-(^dY4DXQL@Z=YO@5Ebg^@11S2WKM<&(_;UN3DY,T6TUWYU5g9<0<V9g
Q^W7V9X16<QHND99]O(\dT,ZT>g:K(/)2;50]?ZH]aGH)LOBODYNY8SQc)PMJ9U:
]Z<K+G?^H0bW+>Y1SG2FO-:<6dA88P[88/\,T538WIGHS@-K;4]MIB2(O-,80_gO
FS59D)4AJA,SPeF7X2Td)GBV(a5Y1P:1#,:fXdFQ?fa8&@8SCA#2_\JW3;_2eE>J
F+05\gIY=AO05:?5[MM_b\1M,.QaR-SR9_]B\V^H)3W/=M+_EE>ZP:)e=O96OE+\
L64,)?7,W=U9WW2(:Y</#4Ig..a:/fH5R343-gJQ0G.:QL>b;YYTJ(4)f1W]GN9>
dWK-P#gJ[/Q.\g2L>=31bbU#g[R]@JZ+GZSKK_+Z[8e)S>=CD0M=9^_g@OJ@(4;T
f:g>4.;gT3DC.<;7;9TP(U?6-OVD.7^QO)]QU^_A^fbWWb#)<L/8e\P1X73]3=;]
fU=f,D2X,.9<-]D2cf9Yb&<;74U7f&O4?CLUa\b[UU2RH+6HEENO\?d^#g/[f/)Z
O#F+Kg#60VW4)/USS5?/6S8=6].6/_A@5R2E,\A<L1J<-FN8RCRdIZL41:);UYGG
g9Qe@b^VU;^KXFSQY4F@baeF?:7dGHMDbK;33(>B+af,SL>;9GXc0;V^RfMIVWIa
Z[CFM-&RHAB&[Z#TE-5R/1TGN8598S6JD?YV#A>.SWbA=_\3KVTM/g3a&^9YRe/4
47&<Q6H8R-.5_5]E&O/<3EDV<4&BTD=Q19G2:P;G\B,f.[<0aDEKa()JMe/<<@e5
)@<<eD,2=3]T>3fMU]bg&]LT?5D\8&FGL@P3EP,TE?HeKO(a+P)RKbc[7dfZ?1+6
KX:6Q<&8J0#b#76\P-+I&>BE47RG0bX_NC9QI/##-LN:F9&9Y0g#b)+_g@NGgAAV
G/D,4TJH.BO=94W?&Z29^fRP[<,@I.?a;P(>.]Y9^@4WZaMMdBL#S)T,0P6,O8R[
9ML<MK\6A@S=I>.eaI(GS8UCZfG^40>:8)Fd<NF6cA+]5Fg33G_+OA5218THc6/)
]HCaTW>YBf8)B>I_=TZKVBNW+ZI#N5G&,G8GS0I2=5,A\GI3)-,LC#23_Sfaf-\1
M:&#F+/dXPJP85XBbP1^Y&,Mf[Y7?4LVOV:X#J1>53-QY&?gcAJ1b?&)N+#HbOXG
d?UbHN=),/eR,d];(QT?^(fK@Dc#D=R6W4PIQ/\bRH@^X3C(ce15,6&5Q0e;6Me(
6ELO37F/Ia#GT@c&=-_Y(CCKAB/[4Y_K#5D:S+]0FY9(YH?11:43&1:VAFK3[4d+
C+6+>g.\9I2CT\EIIVR^D]PL:b4[Ec-[.@533]]OSW/a:L+,30,5@/<LaAN>W_Q(
0D.1<d:V\4AXI/7VVb/V1.8g3HdDJ]H;#8RXWUUJF4PT[.>e#4CM050\eY+BdM(6
NU77OU5<.06_G:=/5eH)=UfPdUF_&SEGHcg@U;NV),.APb+Q_/#bI8,&?+6IQPT)
?M^)eI:)O[\PE2.#-Uaf<Q6Y0[<#JX5BWI+V>##;NSKFJg?-N3=5(-I.Q(&7NZWb
.4>,:F_e6PGJ#>LSeE#]]&Q#.B6=S(+G?8b;965PBU5C1P7=+A-\F4>#/OTcF#AT
-=P+-FES:HVcBe_F64,CgA)\07B-g2^BLK?c+]P#BS697>+d(@.H3I4fU&,b.(KE
P][ETI9JbQG&EGZb]ff+T;&P@SR+@.aW?L+aZ#g<1UN<:EBZ3bbCP+ab/Yf??X3W
?U\HL049?aPHUU&.d=)+BgJAFgDa>_7@9R31NMB..F)#bUM^PNYbdZFL\IQ_5TEY
:MU@e.cN&T:><^\5YIITM_0ES>=:E?E=1T@MM&\TIbM.b(NIAZIO(aB,@7^,U/^C
\Ig4KZ5?S+d;[:LU&YA_Aa+.?<XI3[Q^=d9RMRc^02d7D2U\fM4Pg7-7O[QfJb#^
1OL^2AcV#GGWUFVO/?EJc>66MI@51FA]Z]>/8V)<D[-:(_bBE_dUHF)NGU\#2,0=
61&SD0UK_#1eR;;d7P@a);g^M@d2B,cCg9C[PX11c)>,ea#1E]OXLIKM(S/,_E\O
RaIV^0A?9&?6QGA=K-D67WdMgQ:#eM,]ca#4Q1F#(<L5]@-S9PX\/5R(3&dGHT4\
_A\&1dVF4?QfJ3/W5J5[/_F28?QNO_SgO.8Q]JTLV1VYZN\ZH?ePHZ4g_a^6CW#=
F&TDTdPaBM-Pc1SJ1=JS1;V71Z\@QJQAQO?Q#b58<)+<-V2\J9.\7fPF19c3ad&L
PU7:0A?8BcbA6.<Q4b0Kcg=AW--0_1c.gG-A8_W&b_7<9,<0ZXK\VY26Ba)CFT_]
IC)(Z9K(K?Ra9(7cX0f+@NZdRR&:c-6;W2KGecJLLe+4XHH,/DIdeVNfb-MZCPFD
D80:f\IA(.eBMJ8OOe<b[[?C/L4&XC3NFCWKLL9_/@\UK1bGI.fTY92F(7Vfd,I.
0WJ,W?4A<74ReTcG(+6/A+L:\);a&D0+-.,1Jc.<+cY+LcWP(QJ63/dbK[6MGFHU
d:eF-RA0?W2=\Ef=,eUf=@OW-e09I(-D2.9_bZ0.4NH#CSZ)F#V5S)Rf&[eT4cN>
H6Yg@<X0_=RdVc8e-OWOH?#TC>g;S1-&8eDGZOcPLWf8,G[ZV1K#L&e];^/;dC@4
,D_8M#__(L19g)Q]\Me3:WVJg.93-:3CaaG/OZbJJ:02A2GC300I)b81/EJ7<ED&
[ZgP+,R>+\:/:;1;?DDaNDTPaD-W0OJ4+3,777I]4FJ)/HcP:9ZX1gWf]\1cGH?5
eR3bOP>g:I_9\_OY<8EIfUR8a1Wc]9Q;?):18Z.8(^TQ@ba]1(:X(2)#VZH+U.WZ
+fRHYI3C.S?d)S.>6YF?DA0ICH>Ea+VG1_0HP4_[N5XG@SOXNA=RE#B(_JF@ZTb7
:Ce<)^[HOZN9g:5TSVPCC7N=(Nd++S6XA<&8KX^MP(>a_<?Xg[SMf51,=[e]f=T/
OcQ-5SFP8T;[Y7JF:MC\>6<(?ec\dU1QF2cYQ6a;3?cX[S^b,./Z3R82U3g1Y<fB
aGQ/-#)_F4d/[_^-YNVA9NRDGCa/bSF,S,F/L2]\L5QF5F5^?R9e?.7/1;&ZcQ;c
[#(]cg>M&gZ0g0EK(/CVMES>(RKZEcA068);,a:Hf/#]+D<[)gU,J0]IeHK4=IXK
]IB,S.W82R]5XC.gJeP3R+S.gPZBGL&^@=84d+,ES(HT@aPF5RA6,62,[,L1.V6/
fg+6&.eUVOH<_5QTG#/LZ[0V<VX>9.c3H0F,X^D.F5C,,c1_]-]?d36@T3KZM\V\
:3bA0^,Ec(&_8NMdZAM]:(Xf,0+#V6;baHH,<<<=##e:]<W<ZU5&P#c^LOQP:(4c
5)(<IGGf:J]+UeIgd>-SYe6ZZ1#MNeTCbOX<+&-@AY:US;Kd?1[7<CB_T@C;Y<US
Qa#L9TQ:KD5Md9F?^168)d9a6N>e+L.1F0W-87>#[_(S:4;eWB)R_XR<W7QXe48>
-+[8V3RI++<6-QX\D\c/8aY\HN45B20:&64M/,a.GSPW-\E?Hf087_>S@[7D13eS
EH93,?fVcF]dSg2;-e7FcX(--1L;L7X<PUf]37\15&ec?D^aE?L+L@WSZNW-90,-
=D^47TU]&EXf(D^J;\.)PMW(\4B&[7H.f(VS<e-gGIRS;)=g?P)+3RA1WLT\))A\
Gf4>BXO\RO9-]-ZY-.K9@L.)Ya;^>eQ+?\(&S.&aDNTF+_Mg_B(#eKgR5&@Z7Z6T
DAg@9bbg]T6Da6WD?_).#5Ra;4LP0ZV]9;.W(2],.4a>:(,SSW6^03:(^#<:(Waa
ea1R(IUCD43(&(^Jc8D810VKDUZc+gbc=0LU#<NCCaP0Z+e1UW8a0B3>?[59[eU3
54Geb?10183VKM^YgbVd3SZ.=WG_I0Eg5D/W1UWe;#Y=E1TJQg@e_T;;V5#dKGU<
LXMD)Kf2>Zb>-&_:6LL,?,AO@gS1S6UgFFA5.YOSX]dUGD:@(CG_,_V>;,?GU4e0
g#I)&d3d\1TIH1S7+g;=C7]5:JH:[O_S[WWFA8-:Z)d?1g&J-GaN^UF[@ZY>JGOa
fAXHYIDS@K##V>G2e#e/AN^L8#/fEXUET_]KcDR^/_Yf:&29S?&Y/=gI+/NO7G)R
/1fBB+W8OSY[K3U3#:=.J@S@9#QW]RYL-Kc5/OY?aaa391>cQMF+<bZV//0S)9@;
=[e-g@eb)S,:PH(85B9>/a0JdMP[?]&8G)>.#@;ML./\\JEAEBBYGN9=0\&(Of^R
-P2B@5YH+7[#13]KC9=9V0H>.[#4<65f]0c0+@VDNR7Y]4Z1Q3&#X8]DJ_31GJMO
AeM-+H-+;GNH(]ZUGX6KY+@(ERC)U0^G7().g#N5dNWDKAM]#18f#QG(7IbJ8JJO
\.8+II8@,(6,5_+747a)7:>?(8c#F+>g=BQH\^L[W21c?3@a:B)E+2M=,2U4N^J<
2ZS8adXEdaUDeIQTbXN_-C(]?f,)F9VCJ[0X(JQg?J:?5>V[.9JfL\@Q2ecFL).7
YEO&&S&1[Pe<Y:^,LIcaP#9KB7.&e1NP-,GJ6@12:M?fX+_]+BVO@Y9]eJ(;7B&-
3T[W^?Q:-<aBR:#WM:?Y5=c;5Z&Z\\,2XW,c3#a+#7P?+1,L/LaWSB[-AJa?B/e[
cNA,10T(>c4W(AfY[>B?9IB(g8]C_Q2I4:QMD:D=<+PXTC2?=(fT8deRLQ;c:\Y&
+LR(\+6<=,I/gb?/_?)&Y41HN;N9FE(ZZC?83YW>+c)9T7,D(f8>MJZXG73J@a@G
(.NXaNAF2&aM5=UFGMHLRC>23c?O#O,8=:R.#94c3aeA@,J@1R8:2W0=/ZR&@9V#
135IYXG6.f&0e2cc8EIa5cK8d6fEX;J3PHW616XL./VUFDeJOQLe?+\DB3#cSNG2
W=K6Wa=\@,Y(<.FG9UF.H0L5L8AcJ(,=ff44VLVT_VIDHNS+N5/cZ6(e30=<H;57
bM#=EE\9E2Sc;cRME<UfPJ;P9TaVROaL>XeD_&ZZVE&F0WPJ2Oc8^D1;5?a.&M,R
<=F02E\QX9\IQ-]R8F.;/R=bD?:^DC&2AVK9-X/+18^^:g_9Z+^E8Q.X[:M=b3&A
:O\SGVNc/]IYA_g++NK87\dO:geXTLXMdG]&R@f(2e9L\UfL,^[LX>.5/0Wd>VZ_
]VH+D(>[M90]8VV[bDQ2e:Fe97?fXaQ+KHB@#]Meg4(WNMBXbUF\BSHb7[cD83c5
^QFCWfJ[X;C)T2NBNDf:JR8=JUTI4XF_2RHQ>Oc<:D]eMU3eI0=5.#@3.)<NHUQ\
d#.6TgX4.bZCa,aWQRXI(IN^Xb5&cQG?;NK\:_:KfMOY:1]=CC,OBHE4\3aK>Z#e
DG_\0+Df-N#cG3gK4I.2ASOF>Ac-W4-UV>._U]O=DKD:cK2d#9YBdafCRZ2?):\b
f>BDTUS+@3^<X5Q)FY+g:40[cK9_S.c:dd@Y..T.,g5c;:bDI42-KI^L#/AWG)Ve
M6fd=/LX,ZTH=.dDD>EENeA<E.C_A:6JDWc,@0I=C-@+fOK&TABGfH>Z^dSZ-K0,
W^NCV0AZE6A85ZPCCB]NKIO3ZB_L3>-7,aUD^@;ECc:9O=_#_E=)SU>[aVXaG-I[
[=b):/N5GHOf9gYb]0Z=c9==8=,WFLNPK:5PUNebGGMg^M6I@B__@TA6,ECc8b?e
2OPOa.N/7Y==[=&D8\R42Ia9Qg-fWZ1dXf3R9GeROVHU1KGdSc(\[7>FGU139bZ6
7EGceJ+Y.I4;KHA(3f#L^Va>M5JG:[W<-]S/X)bW\LO>Ld5=WR5AaEgVO,ATOWQH
0:Y<)SRP6]91FUGR=?@Rg83_0#Q95IT/()b:2W42(P9[bJ+2O_-,91Q(eX?-ELAT
g-FX74@SfO;]f2c6,^f@\bHB=CX4J[P.6Z@C;2XfNXEYdVY?LMHU/D+X_(,,U^FQ
OA.a0A^OEe,_)Wc^-B21.>ONc#QID00Z38)E7+C\^=<JeX@e=g-eKDGc2_MV>YNA
WXfECaQ)/;<,T1M(=B7\(\Q5:@=TH9,0L)9S@3]a3\c02_cB(@/&S6g@b]T_bg,F
ELWS[e_[Gf>9d,J<-7eXJNQ7BRKRY+=6]Geg;S1#e):B5fD>=MG)];0L9#eDg+);
#1\44@.SVeS#64]7(C5MA&F,_FY@)++K3YU_^&A3Jeb6E;cGMS3;SNM-S6Q#2][a
0Z^)4CV.L?KC@#2gg]T^,Z50F@XU7>J;2\EK[(KPG=MG2MBH2;1[9(NMBS_8gZFK
20]6Q]3SdGG0D_/UYeAAR5FMSQ_&SaB7OOa<CSZabcLK&#,\gRD>[e/;<\aFRb,0
e5TfP7;W>5B[,4B5S2E6c.b,CbI;IBAA6N2YNd,8>=LCG+:SI1H3CA]]DG07?./+
6P-HI4f/[.^:HcBQ6,USKW.?E^B\D3G9-@0?Eb:BE2\8a4INA?&<M9SIQ>RTDMK.
T86@+ADD?]_AB62eGWC\=-PI3&@I9J4cf9TIFXK=.>>/:3-@<NFD=,MY.\&6JE#^
fB81<B=Jf_Zd&FFGUA:F:_C2NK+;24R61^VC5A<AT^</&@fH[29E7cT(E20DW\1B
GWcM?6T9FCQ(+)]Ya/\\\4_EH+\</ICRaaO^CePT8e9@DDSL,</CGSI;8<MN][XV
[KU-E[M9aSS:1GNBIP=A?72)DWPcHD_]B2fQX?T^BB5[_><cGRG-GO+W?G&)(5NI
>.M6LNL6J[[)8:?d^O^-c-DdB@J.>QZ@963HJL-9EAE8XfTEG9WT.D&S,_TJ2^KN
PBZJgFg+?d^/(/EbBUC525fXS)aUOJE>=9ULf?e,[28D6EeD&5K[)G]M,eE9Fg-F
0-VFeD.F=O:8,=A]7G?5g7MeCWIFc81]&2R#N1>MR@6H,B)SP1<N=:Ld-Pcb5_1D
(U6=POJXLNb)&e32MO#5Q0Q5FBBZ)Q2KJZH_#=:^H2P>3#KG7CRK[63DVC/JBb=>
K&F^P7P&2RE\9DHBM_FOC2P]>/Rc5D)Z;fZW]MdD[6CY^@RN;B>+3K+)/^4SaEN=
CH]W3+HUX@)4eb\W/?Le:IRV:I0UZa_7U>2Ac#[7c3_QIUF9dRNK-gc>Z80V:=9-
f<,_]GV^21/XcTLW(.(QFI^D[daWKJ##5&_&G&gAX3\b6-<Udd2GCdDEPa9W13]?
6/<(CK,.e8V_9[MITAfTTGcAJGY;8B6^H4HJZ-IU8>./,U+ST]gTHW5g]B<E@S10
\Y:Ce]241dB\?PI[4@)OFXaZQM8-?HAF1A4]>ENA,3.Z_-d5XV1N1BLfP<@:@\BN
G.A2&K.;HK6+M-G#b/3IAe&P4/LTK#^dT<+J@>8<[V>0f&^&A/cPd(9Qc+^OM7<[
?[I.fRF(ORAVFH1Qd2+KaR2[/P8MD2.W(\/&I+8I?_]W.fH20_T\7Agc^R@4P[RP
CXR(]PZUSN@9caWa]L76Z1OKYd3R;.]f2)-XOR[LRYB]1VMEY4CF>)eEI=A8g0K7
Ne9U]AME.8cU2V^&A+KFaWBG9<P/2V7C+XMDe/d]@S8B&.DM1<E5fb3C-P-DE5Mc
EP.S&?-]SQJe?+d\C/#D],+4R&_1[gPUa)0g_(]U/g>&C^\V3aLMJ_+\gH?NUD(5
]S7Pf2)6WGA]).WNf6>;P#]PB_A_\Jgb]+0;AI\gHA:6+N&e/=LSVEWZ:TY8Y?:?
Vd-(HbN>\5ANCX(:6[1FKU.4Ue1-6Cb=dMATHB)eAFaQ&a&XA,dDET(2[)F=<;VS
4614X6S=4aHa&Q7G\T[96?6^I6SWbN8C212c5#Wc5aDWYG>ER\VJ\d>&FOX<UM1U
F2D^:-<Z4Y54_ZL(T&ID.c-DYA.DDB0C8WC@?FHf40W9Y7T1C<3JVa2GWJ?L&aY&
C\A;02\VI+GBE^1N1O/M:>1YG.YNNgUSIB]U3\f;ZZ+M?79f+K6]Ab+(/0VeSM-/
N@3H#+Wb:aYGRbB]]O4@=(<F/6:X::7,#JRUJOJQP+\HN8ZXUZWH(F&Z0U2.GVJY
9P+NMRL>>BYgd+<KEGE:-&<Xb/S_@S[X@GMS#-XW\IKUbU<cH@)L,d@8G[]VUR]T
U)+f,;Y<WBI,>KRTXNd/]#fAP<TPO&TAEI&R7cY;I[(g,gcdf\N1I<K_P-+;Y/91
]L>ed<9-.A2O=bAXRR0H1Bf5\9_R3:g7X66@ESLB)>Q5D^KUR^fS>VcG)f-);O\;
0(DCU4@?=-_fF5&RFD@XQ4;;;/-GCMY+e@5W+/Vc[-ac-B-0JDFK&G:&\5G_(JEH
Y0M_=4@DEX]WWZKKdR3F[84(7QBA?#Q1;M(D>;I#>=fE3\YIQH[KaJdJHIJO:PeX
[=J?A)U?N:GgRJ::USZa/1[?4^24fR2D75ebZGW#\^QI>.]_gL#]+]dX4?8\F&[+
EETaV1<3_1QHXV\52XacL9D##HL1TVWcW[YX+DFEa;I[1G4cXZ=HH8S2J_?T0QSY
^X:01b3G)+@^[4T8f=K/_=794MKV<QbRMc61>e?_2H5QN1KK3M_RZEaC/<VI,\RY
bYOeg/\b(,4MMM:#>[bXA.JSU-d\E8K^P79Xa?f5WZMEH<EI6N6L/E-&^,EfWO;4
Y1;7Ye?_fgLL3?PLHC3b3>;^;7=AP<V#2:WVd[+;7YZL,=g-Ga/>R3->2(a3H)B]
Q.99YY/JNP]6+N@b9DA)O,QAd19_c@cLBQ\4[b^@(^37SS/gW<>BC-Dg-?fM?P+2
]+[-g4QM<.8P20.-,W7\/^>f:,A8I54d[W&U1b=SSg04W8O+--+X3M>/<(JLNLH6
[9#8A+(0gQT5g\@_8T@4MP[553MgY]2S97U)LG7S_8IN.cTQLBG/T0PUO]L6_Y?V
A:XM[Xd:2KEWe0R\O5\Y.cLa9Eg55K+EbagMb7dZI#d_+DFXQ(V44Z+K^9@NGLUW
VV];K,F^cO.)4XVcP3c-]\-c6C6Z\(d,WX)CUF+?U,4B>U[=NWC+d,EZB9,?X]E/
(6gaULMX)Y7K/;RO:QMg&>8,4;f2,N3VVY]fI#De/A/DdH;^V[;eF@Y<<@W<YF+g
3cO#IDKE;[CXD^+.HKF(TORBYLa/S=UZgK=NL@)@QSZc,=.FDabS+Q5IE7@+U>CX
K[>FaFT8;>dIM5@gK4)Jd7RXd?=GR9-R\YB-TG+0DEaU\-6,K\QXH3.?#V;H:D<S
eFQL4\1/D7H;Ze4#B>L(LQ1e42]6TQO1D)PUH7RAa]WdR/LH/0^5MWRV]SPTEXF0
YW@1?S2.cN)G-8S]PM[V#SS/+/PGS8+P;F,d\FPR]5XEX84]TGdAXAN;&,+a&De&
R.G^WfBPgZC^[T\_)b<;cI:36>bU\&G#KAARX>F#T-U9886Vf3ULDV&3Q45(^\5\
LfDfB<>gEEJ<B2PNW&d4[1U2J>QIUT/Xfd36bb[2/f,4^e&Q>f>Ag&W_Z63bG-b5
SR53=J6UcD9:(I.CTSQ,V=CWNT[TQ;gU;78FK11TID(FC,0XV427PAV([IN2K1WY
>GU_@8L?>I#aaIa-=c#9#H-P,:(7]58K15+E#Te-^\LD@.<9aea2AM[gg18B24EM
DXY0.[2C+,I0/_D(04,-V3GYMQP=Y[f@ALG^aQ82eT6#cN[C9Z+:)FFO?>b]6TB;
7FIE4YD@FD#X:^Q4?=[=R3DO@a<W?K)8W2H(&Dd]Z_=#5MfU0WAcdHb59OND1(Xg
:;aCW(Z\d31B#2^c&]2E3D]?]MU_R=O<BUUAO1L77>6G+&@SJS><FFIN]<[GYc?&
9C:=C^Uc?aQC;(>8GKV\b?d[#&L=aReZ;6aH?B3E#=BT=P]7NdMgDZZ75=[)XW24
TDN&NdKCG#E_.5@+AJPN1E4P7XQU:C,JP;_Y>2f2FITb/I/1J2&(Zf5TD&G-6XUE
:\D,,3VZ?@^?B=@+,?5HeYP@,]>YcV6)U+)a9TJa.4,&D2a5aB3O0M)^J/?cJZJ]
C4_W0\fSZA4C^RIDed<3M4:5GOb;aU5)YNELfPQA?TCdUH,\Ed84,a=9\<H[0I9/
)[UA(&VB^Z0\]V@>B0:.=-_0)Y[M99=F9(26\/gHM]4eA4OGc><@8)KR?2:3Ag,[
OCBLP3b3VCA#3\?;E[KMb01X2bCgT(ZJLWE(OWWe/11B6ZB+APeP+N7;b<=,E\X[
eS0TdDOO\-1/#Q4FE#<-F?#.<ZG15GWE.Ze2KC>T2U16fXKS8BI/?d2.WZOdUNM\
Tb#_06_T^#]cUE5@\=bT-2gFLgIKY=UFd_=V&+0EBK?[?@N;V]7/?<2[A;D]WeJF
K[0US^AR:LO-(a2O1+G<S)LeZ]<MN=S4c6A]+#SaBb;^X6B9V)c.;SMPZ_J[9;9D
D[J#WXFdR26I^&-E>^ZJEg>)&]I3VA#6ACHPQ54,PV\HC2P9X(EE-F?aW]Q(2@Z+
/?HJRA]R=6bZM@,7@g(R]/HB])#-gZD,EE3+,3))@6/eLV[S<A#:/P\#PC0&1IAE
X.V6cR37>BW)5\0=KKNN87g0\-+3\A(cFgLd&9:RcZ@-(TH47AGGDIB)K3b=aJKd
&N;@/\1U9K7X<-6TJPb1AFbR0@E.^#@4c)cb#b+[(?gZIAG]0F?^)U:<fL^a1=e<
X(W8A.,DVZSc^d+;5X6K#Zee4AQ#)6>W8^S<6\>fZG@;?7QP2B?MF^Ud./5OA0aZ
YPA<eT+QD2L1ZD+2O]PXTS6?&+e(5U(EL#=<UX)RTS))(X6aLc6\1^;Va@)1-+6d
eFb:d4]&>,<AM<?^0YL;5DUB_RecBHdad:K3@Y/D8MW1c:+]ecV<@JOZf]WK?U=V
2U],JMc@C\b=B,+_<\UQ(D^@>D9LT_Q9;:ZG2=S/6U3DT/18@d8Ve?07Fd8#aO,V
A5U>D#OFT=f_6R9(9[070fTP\[V(E6Q5?^/U(??>66^D:3HX(2E<?0QBK]W90=VB
^b88#G&\C<U((e^,<:F(eO\P-E&Nd^X9d0TRB8SKWb@C3-V430(?AOXR[LYQ0^c0
Va554QXZ8ABa@J35YI6KFSOH._d^2dTP&D(YVKA?+Q:3JQA=c(M=,f)J27e+FTGT
^4]98)@6AYBYR9BO6Ya(O3a1FZD)=\9NE82dFPJeQD2B;8?HKIQ>>,2):7#d6#H9
M8gYQ1I[>_aL3eOO:]c+)WG#4TY:M^&6[=^f^L[9S.bWe)<+TKLfC[J,BUbG;A<D
Z^Ra@B8WMY15IZY+G_M&dHZ/UJ?AZScE&814+JKH^6?IM@=[0VdXMOP1gdWG;JHb
J3)+H7/TNbQOV5/54IfgY,J4NT7K(.RIg:VEAIGLa[^4BM2EaQW)P5QS]=,-(C@Q
KGdWc^@1(2AKM^CO(35BVbE&+/6;O4^9I1@g40aaWA:)Pa=A8F)e:3^_CG(&?-^B
;XJTLcNV?0)90EYMN:+;+e5.IE2#TP]3>CJ8K]IE;gLL6+ObJ1>E\TVJaBA)g_f7
YD\<R1YfS)B6>4NFc1:=NC.S;]4(E\Fc]Z@DKb[C8)=.OP_NA82b[F8-3eUbB]RQ
fUKRU0X3[CM(7gLWD.IHe>2#G3?gPUY62Y^[M&RC\P@L+3Z,@XT;Q6>85)e([J#J
b.N\b&-K6(XMEYJ7bL.KDPQeR2;3O.)WY=OO4(cV0(/ZOIRe#;NK8f.ged)g^_.H
I+GW9e@-MVaXAa2<XTb0#<F21\E#Q(2gZb#:LT]BUBKJe)W19JCXIX00SDWf1H[(
cCD2=CQA?W0P8(8DP#,Z\Sc_W[]5/OL0W-6&](BA6#AO>98SYV_5BX9H&D\e=B)X
W5Z[W8&;SQ/E./bU6Y+E=ZAU\3W5c77,?KfTeCXfLaZ@1cO(4U>Bd0fc&4BP2^/<
L>bN(^=H-QYHQ+QA)KK@\LL#/D9HaY/9P&dOgZ2Z13L,PWaY)e_]=[2XgMMUJ5EE
LX+]a;/I7#We+S-UJ5ZI+RX.&HfT>Ye78U1),>gK/>O:aS).b-3BRX<Z:[XSF7f^
PBG#^<#UD)<J5R)&_VZ:)V[,-L-<.&^Q^E29I1a?;R81A)?W8_;D0\7_BcAN?TP6
C;_Sd>PW6C+5(D1<=LcB4+P56U0EO8^^RH,1Re1BXFYKWXf+DQ:gDUbX87aF.L)(
)^66\VK&NRYTS&<H(X6fE+?Tc)M]XC.:ZIJXJTbQ+/_&bfIR\&:U10OL[+KER7bV
K=I&1)7ZG#g7\3f?QF(Z-Y^_[d;WCgDJcL)a@WE6BA_f47?E..7gcLd_5>bVF46Z
J1b-XOKW(>LG?NcFb.WR@8g6Q<51E5GAHf7#VIIcSc1G\0N\]L.WN&bXNUNB33,N
)WZLO2T3;Od,J2UE)/S+K;2MGeVaYH1gXf;6OD>)0:KYB4e591FRI9I0deKSb+@7
H^>ADL7CCH/ES>B/Db5bKEfIG;]g<SVFR-4,Q)42GCH?Tfg0VCX09XG/+5AP>1NF
Zf_QFAZX6)\559.F)Ne]ZO;c1Y\WLbKA9)0B\EG0-cQF>&FWTA,&019N2cN04WX9
572?@@HM7AX3EN7]P,AVGFbHMHJ4Bb_f2fFSbU=d?c]B>=MFDMfW:@V\XTKCDAI^
dV&GMVIGdS=Z7[\-&5]C]:LJUL)?SE\6Ba;3Q.25KEYP2c3F-;_UGgZ7PINaGe.&
Yf&f.SF>AJ6IY&#[Je@L=<)W_/R9),@3RB?d,?TJR:bR^B@JJaPJ9&B:Z(+L8XS4
JQS;/>F3?VK@JOg,-T_e&\_bJ8T:X-F@DR=ceFIdWKMJ3])=^be#M[J#T:CF8W31
]-KO_TU@dADA:M/YDW\J9b7OVJ/DF6NFeC)@XY1B?\;;eN3TaOb<J.abOF0-.B5>
2<fB6JKFed+QUX>:43>Z.S[UfJ9C__48>Y)F:_)S#9O&;+UDfKWZ>gSfO]+bM6cR
fZgTE=KE>FaMgR=.2FJ+H)T1S80V_Y7JBQ,[/dK<D#HMS5ODP^:5072g,De<@NNY
WNN[I[U,fONG>IKE^OK@+(MLU1dYFC..?J@L>,]CHN\&:dMg_NPFf5RRU24KJYWR
7O=.V7D0RJL+ag)cEGQ?5A/OBOUO-]?gT;SeTGgWO4#gRNfb\I\#-XFe@8@XXLS(
I;+UaZ1f3MRbAKAG)Hd:\AW1Z=\\dSaBZg[DL^..WLNP/E;BP-gd)W_3KG\#_7Ge
QdMd_N/a0e;d<M2HYG3Gg3N>/I27-@aNZDD4JaZ,Hb\?U[HZ>N2f+[./9bg\QL;7
3E\\@(Z0+4@?3E:2_8<.IaZ]7K4RfM)b:&06eI#/3?@Cd7O6RJ&eD7f^S7Fc_55(
g40dFX@S:gKIIM1Z8+@TP/fd#?-fK9:VJ/5L+T]5Pe&PKFSOQT>Z^,]=FRYa)^S7
G;A23Le4+c[N+XUg7H;4D]V#]DPF9<<Wg=:>G\_8Ga7AVZBZ4/G8Y/:3[L7.)fHF
=DcCW7M)59(E2HDCC1][.XQTPAc=@J6X@IWH+7//38<33Oa4fC^Z9J6U+#BaFVN]
)AQ1A+[gF;NfIJ3K_.cGJUG)SW54W/QNP[eRY\89.-_0HKV6R]69I9/.dAL+Z.[:
\(6Y:IIC:(SXdS72RRa(7bI&L]H0,A3fM)3<bZU\+:U]@Q^<^d2d32Y,TI#Q#AD)
DS:aVKK?]7UYT_=2WIZI]MUAKWXCKfISO(\>W[;c&_]+8N/4?;B]=D^0N4.8W/N]
YffIJ>GYBTKG]AdIMA(OICbQK10RK>.?9+FN[LeC)SXKc:Q5c(NA)LN+S_+@aEX=
<:CS?a6J2>OJ9;DP<6gWbQ/3D9<EG?U9b\6G7dJ/I-f&(FQ8a5A.OaXY<Qc8b_9)
^XOFbSS8WVM319.2ZL#HU:-ecJf2(V[LIZ;C#R6CN2GKE/3N0_8RR5CCSI@_CHY1
eWDX?L97T)=/.97F)<Y,^^S/+,fHf;T.fa&H]I?#(_O82(UL]8[XA)^P-[69g?Zd
G?dd:L@BPWBB421.3fT7IJ;Ce9b[67A2Se7<)Hg_Y[:^ERDGCCL.D;^/^AI1<JA@
^O2P?(2KR9.#VAD(<8L[?54C-=I(ZK[U)6eH.=>C:65>H/.E^(=aO6bI8@QZT_fM
\(>]K/LSAQb6AKDK07N?ZEc_a0#9,QU(O+Qc?QN,?<<_@@V.2gEQ]US&3aP]A#P_
Jg_2^WQWGMW>SIKM\@#9<gKXd#+5LFE0^6870[,bH&HV@g+/MaI^BdRSYF#RH\\b
Pa2)69<ga^CQJZ?#bQ>YfMO8KJ4[=D[B(-QIW6d)_b#/X<(K3=TPU>N#8HO<U^.K
C_LI<A,_-GOJa;D_QA,2[6gL?9S],W9D[#0H/NbO7M_4GZ4g?N&5:MW_YP5c6dJ^
K>,+dQZCQ0NZ^dD(.(@)M#^gH\;^-G<R[Ug]T5&QX[=D?.WKU-Y.F]5-1cf2_=?P
c&R\=D+J&3;fHJKM>GZ9a==6NE\1GXLGSV-7@UR05Gc8UNBH]UH\bO-a^[Je=?VR
Hd7WIT#NY+_S2:A6KcGGG0G+SVW3^,OaOJ(^<V>XU(U-[4RS5.[@M1e/X[FS_Mab
O9<J__5A1I.OM:fQ-Y;g@<(OM2SA]04,P:PLC,?62T[K22UfOL]>5ZS/=3?MY&7_
LS?#+IL_\(?>;X@HD^Ec<,<;DT._2f_+VH/>-0Z4VS0=#/\X0d:BV^@YX]Q@PM<V
KGH1@-BZ.P?1.8+DJVQ504Bc5GB+U0aJ,TWROeDX^5D+SHIBTDZ5+Z]?YbEB@1R8
=e8J_J;:PZK6\A,aLL6_>3^<WO0Tc/[^>@BR)#=Z3I_.U0cB0.5N07\\JTb&TbK(
/]24=DEeGegRdY-.#_]cKHZWE_Mb#-6UP_(LIC<C)7,GcBVa\_\X.8V6V?_M(;\(
2E11/UPC6\9_S6[40W6#/&S76#K+f#HSUI6F(HZf[]>J\QCFaZ<LM)^ITJR]>:^#
gc<IVA#8&U)>,Lg7C@UD0KTH0102VA9>21L/V)(MEdVNb17?8HM0G&-<d-C1aBCV
/=G-DbYKPZeELgV)K\C0W<KSRSH7ZKU0_4Y^N=SPd>WdWP4Gc5L6ZC_K)U^:-B)\
M?PQM\=LYRVT/<b,G<;0X6bYcXaNCK&cL1#T&c51:\68eJRBV)6EP^&-_J3&:M]/
KgK-b(M6^gP[;g.b9d3Y)R7Ad7[ZV]S>_6T2@RYB\;DY=JO^YHYO@4GE<@)J>KBd
M[Fc9(d>9RZW(Tb)=f>I1<B9O+4AS].X\Y:]/C_>a3FM;G+YaX#,\0FZg]8GR;:R
@_292Yg:Z4AfE/4Od7_Z4/H)8K2;,@3HEP9>KPV+\FMeaDMgN,e80U4C)&5_EP_E
R)L)C&SQ=8X7TEdd^<?#9a2J#[+a1@9W.+FD3.^0,G\0#<+f8XMUYBZWWSEe>M/,
.gH0F0EX>=M5FB9Z[E>J>^G-#G8NR0.&@?^Z=Lg.UU[CEB7^&>fKcH-)X3YF@38R
GKdRUb&f6:OY8NM:c9[U@YV(U)Q-F2=]0A>K6aVeE<>P828ANfFMTfV9^20N@:V+
#C[K;+/ZR5K4</d9^Q3(RG-3dcKQ79JX9LGH<U&MAZ].aLf<=JK_Q#O9IY\K(MXL
>?98AJ2Y7TUG[3L#g9@U;>IPa7FC;1e/fRe[=F^/[#G8WVfaA-9AS?<]Q-\-&?SR
8.#5(#\.(H?Fc3E),3N_6GA_;U&OY2_0P23,F3(b\2CaKf<6I:cAacQgI2ZS[bd1
J@<K3Na[A?+GPGf;YZDW2\5M]E[NPT5;T4L1BbP^FB1RTa>.B^14fE\HNJ:/.B\G
-?CLF;Yg5[YAcF#/B,e886]SGFMR0F?Of46GOMQBGA^QYR@;fLO964G51;43C#3I
f0N\DS3,C@-++,JY?[NQe]fbVM+_MI:T\M)3\Ke,\TDX\<Vaf=EHZX-B<)S]1W?&
<NXEKHg43_7;g:=?J]?KRJ6Z.D+Z0)>ZM,S[daOb))0_@#7eS(TG6KFZRR:YPIT5
f/?(0\<4Q[KG_H2cMTba[G+@.C=b[DKPP0ebAB.^PQCP]W00Q(UGF/C25J-E[;2F
^6PcXB_/;MX:eX)ab;5bCB:S2[>=BP=JY(We7?0Y3e;=MH)YQN=E^[ObI0]6J?G6
Ra1D=.eL^,GT+B86c[405MW=OUP[)(DZ^Q5Y9.^5QHPE,AF[?0G92VQG[Nda_];e
;(3[b.<QK=QK[\/=JTbXbB[1T3^O9@/>663JFgcC09<]?ZB576ZTK/POWX2,W9S_
ZfX704QVQJEF8:;CY4-e4)/g,f^U&(1^HB?+JL-KO(K-<GRZPNK:[DX9(WOd9(<B
,Zc>IIB@(QU;58>d#],S7gc^J0&S3e97[G:dW#S@g[^=P-_,6KZ7;Rg>1UP+>ERc
=_V<.><=.ca6RJ&2?O,MdRAVOZ=8IF:IPCL8dGG.AV9?]/?(QRV9I6HYJ3;HZ<4e
Rg;M@>@P2>#-&c>QYa?73_[<]cSbGDVX6JCNe8E#J_]YR.>_@.Z>(>YRgFJ6R7Y@
?P2@SeXVFTZH5cIH:E;b:g:3XQQL=EfR1B(D+ZKZ&_Md[(8K/,;TeNT7U8#>\[]U
S(2;+bE\;.eb:=SUM/7R=D]fG6J:+d7#/gO:.C0ZHJGL[YSf,ZSQc^DfQ&,^Z_F)
WQf(c-gX[,Ta9a[[N.&HWgG=NI3G48T(P8(,eD.cc5Z51RM#PJ>cK-<DZcSB:&6>
HS@Jc:g8J^W,K6LRS3^c#:,?_4?L[\,@,6^ELJY\(QH899d4,EC(=MQG>CJE/]EW
7&&#0.^fZ@27g)XKY1d)BPWQ\&-b<Pa8DBWd^?&-L)^,CKHZM[Lg<0=K1/2BdFM(
\5B@&:0[f?,MfB#354HU;SQ9,.)-R7<_QR)T5-\4,WcI[1=:VZ(3323.Y9&\=4Oc
Bc.J,1]c9K@c<d_Q9aeA_XT>F)5V3O366BLfL4Oa:PH\]P[E,ZBB[_f5\G9d4&Z2
S-S:g3AYgE[gOCcbbX80=<U)]>RQGgCg[U,)3X90G[6@KY1IC9?C/;9a,H/N\8,c
)cVV=YU6IGgT6_MI8B)LZgbGW<;?GZ=^T]aH9?:6=,#UR)Q2Bb4.O2c4&+c5(UJ)
XS8,gQW[&+G=2Y06QFY9HYDa;RY2IL5JDXT-=9WF^_AZX)^=G&[c:bJ,?T^.7fA?
04^-=X?JZ_C#-?.,--1A/^_ZK,)4]58BBa23_I7W9^UR2.TgKYV+Oca)@_4W8Z:#
gWbCZ#AV0&N2KC)40RLYAa,RSGXZ7f]^QYMB3MLa/C)\fJPU.W(E@UgU]LAF93N3
ZVQ4[gVMMI7ee_<H6,G,[a@\UQXI&0?<[QT8?OMa>e#bTTg6Q+\4&T>6\^0\Y?]G
+:N,:>AAc7838]7MOE::EZ1Z=LA\RHIK]TSbZ5Z&1d/R]E@71Z5I_[<30&YP>__g
g=d-fXHH7EZHJL^-Da?e&X<7>FAGIA_B.?KQB:4)ddc-9#:cT,XC\1Q(SZd7#Xc(
(ZbG[D.)Yb3g1235bW+SdSMXM0XR__MNNa_2D.6V]C<c(@V94cF@5=)IK54OJ>&H
-f;eX/UGU.3^X=W0F^X8-g.1H:JRUNS0a(VLc1^KRP<,RW:CGK.AO@Cg9/Q>W^@6
>,\TGEWF;GGP@Z#+6R^UZDQ/bF#&_Ha<e83ce7ANBafSB#4[274=K((Q2f#P@N+)
2PE_TIcIN\K3M#e6F#.:_1\?fM9G28L2@G^M/ZBXM5\8T:;-9_+6O)\NGMI#77]7
K0+gU)Z]YA<[QY)#RR9E9<(^MeZe@8U\b+aC@/5_EL2GbPYEV:.;<=K<E(b]A3DI
&[\JDGFTHHTIJ&Cg3O-(92?@&OE8Q9aZb3dNa]W84Pc\OC-Ab)@fI_BMK3LR&ZF?
;A-=GD@^#acNd-:;aFNU0D;N2G6+M62cK6@WbRM00MJ^Zd+f]1J)XX9Id+3.d=Q[
&CVd/.,#G#e;^/C=-1a:=B=Xab0Y#Jdd_;c3\,T?_7;XF8OV_+B#_AD;RNQSBeV-
C]C7?LR4_4]CE1CggL:FaRAE+KHfdb2@I&?a9/+2faY=KD?YPS^:^4&@KCEQZF<+
.:PI8e6Q[S3XWeNYD)I&GQ@7?3BO1a?30DZYX0:@D<V^93H-e)JfdcIJ\afN?M,F
C,PUZVKS.5dAfTS(JT#fJM..V[aZLE?EN?UWaC4&cYa0LT,2eDGAFdHg^]]_I4L8
d;C6FOTTaQKEdCRN]W7YWP+0=A2XGKg5ZPLO[)RW&?WSX7UC^I?+c(K/03>17CYB
:aQ<#,DYDQ69K5VI#RJ6fdPM\N:g69MC/a;Q_BCA^OI6=)Z1<.Gf^KU9FEC(X\d<
103T5]S0#QV2MP^29J>Hf?>I0Y_KeQ;^,OUNUTS+K/HB1J=E&\G-+d^1EI;4Q#0a
<3.?N+(Nfc8ddC8d@4a7-O<=G7DaH7Y8]716IQ)8U(;?bCF<Ce&U7RU93eHS38IX
JY/UL2P/-SEAF?KWO=_C1-2;05WHL8PW+7Q1NN<FMF4UbKE>0N0I)#DJ3X4,B2E-
811X,?=eca4GJdW^\ce,:MJ=T>TbO3[)Q?0GdG\KA858B?9=OE0DegIYK3D09Yb<
d:4]6NA?:@ga_0OL#cQe8)2LN-S6:@QX9#M01C(-)O?RU(.e+;YV7#IZCO;.<+0c
GHGU>f>[][[8VSgFERDE;dFAd5R?B=<Z6#&>a,V.KgGUG#I=c8S]9c0Ka@N0R)d>
NUH0dBPdLF#-e&1>W3\YBEU:^0MAEg?bf&Egg0P>25VL.0/:)^,MBDgf?(.TTXBO
]8O#);2FG-@S,X1<7/<^L>59<]B&J#=3=9M14^C)@2;A7O#eREQI]2Z24#f3bU?4
OU:XP#,:_;/ae+6:-G-UdF2]NJD&NM0Zd+F5LKCbccERC-T)O[E94e?.#V)e8LQ0
B[TPa,[W6D+1A.M)[2-=IX)]CG@#.F4</2G[f=b5_IEHY2=b[+X9EW_W]I(]J=I+
8[#V9J,CO?8ZgIIA-/(MA66ZAU,L5<-A0-5b1YM(OL85ae?WUI)IPZH#0>-/8<ST
=+L&&@+bSf4=gXfg&/Y0Ze:RFXF:aCF=QM>8d8PWRHO9YYXQ\]>RVS=^XED(]WHP
Ba3LaV+c8FGBU:ea5N[Ye0HgQ-:;H3ZE1#VaY,dPQ/?R-,Jd1J_0:1\_/U(8Pa5e
LCM\8_=ALWCbNK5G+V7PRIZR+\49B&M51CI>FM>AHDPDR6c:38+E9d431;<aF.+A
(I;f#f<MZZ^+3D2?eW@;2g]dMZ+JYbHeD@=0=L&#TfIV?]d#<fU5JAJa>YJ7M:S(
f#3a7:@gSY2ZfO]UO:N+42eRE5U4XGPL4#BD)&RQEa6-Egb@?:c4OHLJP6V_ZZ<)
>M7QLRQ-@dNe:4LFE,:>gXaCc6JJ&/;88\ec9#eMRZbN=P)XRe+L?F@W^5TS7XN=
TT7G>S4:H#+S7P@711_QQGRg+CZ>TXCBfGM8ObLHLNZ<OgH3PLKO.VXJ3X.U)/JS
G9:U)BYZRbg1X+^>_34P6A2^D-_,&d/2\B;6PR7266eK1BJ=gR+d=,LZ,5WaZ\FM
:C6^-B;XS0@dSU9:J>,E3a66\N3_R..H=1E0T=YLUQVMKJ]W@9DCW[E<Rbb/,Q)X
+TA+WO(LLVcPU[CAb/I_@Z(4cK4N+^N&OW;g(O.L<,\Z=DT-H>/17/JR?W0BKF?-
M1WN.\X,9Sa26YBEA47@9.&LU<54FW]T?Gf=0HIfW^dH.A0057?YU_Od6S.3=OGT
<<QEcdMT_\8FMS;,34&;&ZZS37UJEA[PfS0O:_/2?;Q#X.LJ8d_4J,6:VJ^+Z02G
DFP7N.#K5FJ2aEYO<>]RLJVLP,F[\VP\^/GUY_(-4A,UDUKeB4JWb-/MQc@2?/IS
UR5<\9XHV8.ZMIH:fYbT[0O61HGDT_G\QdSD(Rc.1.JC7Mc2^YE?M8[6;@]+X9WO
FLY#Zd4X]7AC)?f?X[:#WRH=,F1ZLMY8bNS5.^?DaggdA-3\dN3PAUF3H78Hc@:M
JHR9E<?MeG@RVUF_,d3ABbD80a45A&b>IX/4\T2Q4+S<ZCZb9Ze<==&_eAb0-&N.
03>W93M4)e^dYd8\3?fYc#RF,_bU>SV-JCJ4g7g7H_LU/=_9RCYTF@)(1K4S=&3L
T3VBB?U8Z)RI]c\eM?YF<GO#]+b1J32+H[WLDNS59U4O?,G(I0>341DUO0F=#W<.
9,U@c;6FR&#TaZ7-J)/80N\9YfDa[UWT+AK2-WHR2[TE\YeV^L5GD_PbfPNQW8+)
LdaIbR2D<\S9a<)=E\[A<g_H02f4cI&#N)<M^NYDQ=(DRRVSQ\-&C=K9CR7M:RT/
UT[F87b-2C_.H/O3BaOQNaJ@C;e^;H92Ge<OPYZ_AT_JSFAE@WUQbN2\F>FM,bZ[
[G@=E4\\:fT)>,7IDI><YQda.^@X-5Q:(RAP6I6MfC8L>[2(]-Y3_d0,BeR6.0fB
IH^.3;?#PE5OH2^b27-??;,AR5GBMb&7TWG-AB>EGE+,-57TK)1+APCBGaQ+#fQH
K^4>#7H4:?(2DRC>6;SAUBY.B,BW1fMLHA#D=3OE5OHJ&IO8M4<YP7?;VQb:5d-0
d-DYQ_8c+Z;K^1XALWY)HgR_R3FX:0NO#3ZC:62_7Fb;K07SOQ#43F^[J2A28a8#
^039cUDIO@BGAQ8D)F?7_5)\W@,.\(9OHaV/MHeY\O3V>]D[8[OSQYWbL-Z,MU8T
&)XD]0Wba->CM.g.@.aB),7QNSL\,F.gZ\.?C9R9H8X,AO(N?_(J&R/>+:\#&WCV
RM95PJG9HA3GPRA.EL2N.E?&UWbd@cUQYd+b:9[_PGG;O3EYZ.R@Yd-CV(2e6f/<
eg7[G1e_C;F_U7f[^CW6)<<9Ae^C,c>#eHF7Q<NaJ]gdb=8O<<PI8Oad&,S&1c?5
Ia1ENEg>9I5STZ]SPJQ[?WE6)-3Y1>#Q>=BIdGYVHY+aWg./0L)DQV:2_HDXZ#0C
^&)ZS\e37(/QB,Se,e]&XEd^B3WWSMg#O@Ugg9:Md]H?2e4e.&J\0c16R,EN?;8^
e.H6@<D@]d14HUW&O-UNTB9:]QR9+XKW[\aUeSeS4cNaMab]@gG^TMg.9)L#T0(T
=-<R38P7D\<SN&=1:+Qa1@1Q=F[&Tf-RSG(J6V]PZL(aLB<Y:fH.:e9ffO#:OT2D
6F8_)b6\BLeeP#T.>-Q3W#VX9XI/MIge.785+I.e=F,=^cTa@b;\5YFe0QR3+:KV
Q>F(@E2^;3.e^.A.GgAVFECTSRaE<_AcCMN(\I:WYX@O1[6M0YSOGgEe_N4dHc#B
E6L2K@_I8LHF[3SY3B00H;_+gg,:B<_R<[=G=Y&;\42dX;,,\#G,19bE<Bd)[CQM
Gc#32,LUE)[F3_d@L=2dQ4NVMA4aFGcb/O.UE)E)^a&(e[AI:I+2P2^4VV+bI7T>
;MDU0#-9HUfQ=Rb/WJ.LQO(CI3(S&P?#-QVD30@0d;@NSgZL3;Ad5aVSI#Q^9Q4:
(\DZ1P)K5#7086DU/.G-#6)(gOK#@HaV6aX<Z6FSK[O]@&B27a77gVe\ANZGNU;g
3(EcV)#QQCOSZ;L:)bD^[8>?Lf+9[#MBgYIE=L[QA?E3<Y5LM.dY-GacC@dLg)MX
DO1JB5QKE4fU.61Fg56JK#.9:N:>EOM:)ZeAF89[N=#CfJSU@Had&[G=5c@A7Q2W
>d>_eVO6eBGX;G=eKW_Ig9Jb6G2;?I(1N&7:eE>9afE#6>GODc:EI0[YYCNCS;Kb
XN^GdcR\B@[,:@^F[_8COJ>[372/D;f0@I/03Y4?/<U(G7IO,>E4T@YUeIQ;K+3=
OUZMD?BHJIdV_=+]#23W_WN](40N5Q6gL170783Jc,77Ocd;1OMM1>4547^YE[56
F7HDg>Y>L7,b+?O8PL2aTIPQU19]Hd]D=_GPgXLe/;7bOLN3.BHRKH[Re2(6+VH6
J1B^+6(W,6&VVZ-75E3G3QG-<XC+8G.aeO^9JYKR@&#8V&J83.#W7-JZHKa=_SY1
fAaW7)0+LXLFaORfMP4UFXPW([^EC=P=IL0d)TZTL8G8:1T_,VfM\]FcTU\bfDMF
LQ;f495J1.SF]UeL5K3f#UF1TAeGK#?a/(:b4UFNYeY)-WPRQXIPC)-(G=5]XC:J
JXaG=HNIbVJ#a?^@.e96cgC9@DAdVB^3K\@YXSZ+;a#-#]8E)PgLZYKXL3ZMIEde
\@.^5@;5\A[fgP:VXF.HDP6,:,AP28T:1@D<XbV5f0>c([]&.O.-;3[K4a[0Z0f<
8:)b\E:f04V^+Pa4M<S-B9P35A@59AR]>S[(+CeO?[C@b9_#P+8Ub7aAA8]:S&/N
cGfY,^]1d>5(XdC\Xb(ZP7QME+KB6fCagLcab:(/)LLKP#S),JfZ4Q\@JD)e1f.X
b5TZgOb->)8d#L94C<KOf45.W)GOQ4cD,a;_SN3g5ALJPb+Z=6KQ3,4OdIQY])8)
f#VJ)=IGSaG45f-RQD.a\c:]CDcaE4FL##afA10.A<:0U^+2b[N_Gg0f(/P#/.ea
SNaM\#C2D#Q#M-?fa33NNO0.[+((W]Y1#_F\/O?e,3TZA=]8(5Aa&;1AVZeU+SFD
WARc5-(\NI=ZXI(8@be;4.FHCV5JPRc6d3_PRM3-,af7eZcM##C7dQW&=\.E\5S0
:83UPA1Q-#7IFbbSK82,.T]#ENZfF&KV.BHOFNX#TH1C57[#_V>Qa11#/ED4JAbR
cI2WV.dFYIY<JIb&De6^bdH-[WG.C;U#GgP&<7&:ZZe.e-9PKcHRF4f]JSO/=OTR
[f3#+[58\:b:D;LSTDc<W@#R8-++]PB7P9L[G\<c)NO^H;>7HY^]8D3Y[Q^S_)Y#
ZCF^,(DP(IJDe=e_3-[+Z#9G0e2R4BXgC.e=L:P=)e?/N]XD8(eT28D9HF2a(&E=
;aI_JCUTXU5OLQWC0T0C/D15=UU?>41^LX,.X1O59c3BbG9ddX:@KcWA]5Bgg8;3
eHSgOKNXIf&P?0dAQeI@:03(<,Ka5g8O@)4K#)+M]3fRAE1)CCO[-2#QcEQ\YQ-1
&ZWK1/6CFH_\XX-b@8\).S)WgS<R^7F56eIC\J12d^Y+J2)(VMKe1]fK9]:L#Z,L
H#14.WKRY.B&?-\N&DcKfb5\NgWWCA__O4EK&ES9TWA6,2--W_U;7d#,T(D#F-Y1
RJ/_Hc/PO0-7TKLf1:-##0JKOLU=7d#W(/JW&4+:)fXOK@gDL#aT[KbE#5?#@8e?
J>d1A.Q5VXA?[TZCIKfN#6Q4eVLNadZ,^TO-)_CG-KM=YS9@gI9H#Ra1Q5ebb18V
=NL8K=?I:6T0<ZB]5Y)O;LYZ#Z=fPFId,Xg8EbG#5+A1OD@#810@7)g:<,dK8Q_T
LXLdc67[OD1C7>[<A4_gQ5I9G3DK(UPa.B=KGC:YVed.dW?W\HN/1F:)FESFIJ)H
NFd_2->@TgY22e?S7#M8@O\Ed/22.-G&)FI,EXd@aHWXGZFf\b[=MfRC&6g7HJMY
+LOL1,O.(KWV06TL#3bZBaNCA67M?LAMW<cT2Gb9TFLfQOX<JBg\5A7^\#Ud_XZB
OGLQCWNF1[,&]fDd1QV62#L/G.5OC33(g0Nd=>Z&N0[6VYM<VVAXB44E-&R=_@Kd
Fd]^\WXM7/+RD:cD7OfN4OYO6^db2FKKE(^OgU<EZ]e8?WA1>9A@gYM89G9WBZ;#
7JII;J0eFa8S1>/2)G62@b5+<\C9KDaO_:;2Ie4W3/dE,(9Qb[Ac4N\LUZ6B;X27
C(BVO-3(I/WW7/Xb8#Wb45=+6gJ>AYCH]92KYAD([662E-U:3J=GP\7g+R1TRgD4
78IO[AY,3=0H0P]\?@L1RFMRC56>/gaE@8EBRP>99BQQ^2XTeLS8B/WN0bge:UR^
g+cORN>@\b;TC66I,#1^D3253.f@5_C@O;4#:1P-+>>b<1=d)L,BR.H;^AZ8/SW0
fQ5G4&YHUF;E0>VUH&_XHc5@K+5]KLf-V>aU30RBV47RD&^DE9N&H-WT9E[#U;LK
H.g2g6+:ULb9TVSUK7/a7-K5TXS7W,0RbWZ#d5:_T33XfX)IC4XWQK@5/6FY]#d:
YNE3\;A,3(Sb\Tc>XC3QE.&[HN,BHJ5:>BUQ?S<EL7HgOc],;b,>1QD60@3JP4YQ
8-?cL6QeeCL7eG0,4IYDNG)IO<[QA07F,<#++F,N\fW5TdD:0;23.->-PUFLYHY;
^=-cZ&^M=;94\.&c+;E[UD#S97[/:?12-#G]PN;b0gCb+]XA,]M8@JCD/3WB^I<R
,@Z(=CMF(e2@268N@a0J8@@;=S?Q?Bg:YX[^\9H]Ag9K9SW_aON.cD=T&,:5g15(
;<b1?A;aV[MYR[3WP-FI\N##TQ7FXgV6d5HBb&P5KgMeT]=6:dX:Sge19U?4_ICV
<YA-C(V#HZ]SAX24g9a>GK/(R0A;fIR0N[<<V;Y@5NS]E^XEQOG=Y_US>.e=g/e-
V4O.=W\^4[ECb)(aLg7@WK3#1X5\PU4><+B^Ie+g6HE)YG0PP))dLe_MUTMLa:=6
.b5BBUV]7<CIZY(4M&M?VM@SgD3E=>DZ]4B)@Pc6O1b@Y2I=gTHS>@)XI+(?KSBO
Y&M:X<&QIXD>(WOc,cK5^>Be-Q&LS>+VdCP&YGWPVMRH&9>UKcU)S_QJ/?,23?V3
VSUL8)P:P:9\;@@+W2@TbLTgeHAN1e7R]d+5#XSf:SKR?T]0XE::A(MGDdFeD>@g
QNX6+3):7NgbZQ64[aVM/OgICNDI,RDQ/OK@M>e6;#^?\NPe5B[<WTYe83c9M@bN
]U;O5_6g/P_4PK&7ZG7X?OW0OTaaRBZ(;;I2;,NM_M5e;Z.7I=QKfY0J>+?A&X(Z
OGF8;c]cBdR#/.(3S=eC/G4BC<7J<052=.,+fU((b@Q^=87\__3A,WFg6N>1<4,X
^Vg4=c_f?LD>)IW8Z0,<N9KRH;,3^-J[a,[f5^PBQ->X,7G>TaDET?8_]AX(9J;4
(QF(]FZf?EDc_1?R+6^(@3<5@BF@WX4Y<4JA?E93PD\73QTaO2Q4cW0^>ae2[36[
S@E[R_Te5_YT;J,6f]2bIP/e8<O#T?Mf,SN^738L=39bgL96?MN=d=[X]ae^#SD<
YV]\0]b#LFYMCL_09c\b30.d<b<:Wd:dRMMOJH&.0U])e61N,Y))SOTM-<D5b.7H
c]M28BO/SN]9I7JTeMJg9,B5+-3)/^&147@:@cYbPf_OBC_dVS[]=G4[4;deUKS8
-8C.FE./VZ5acc_8M>3EDMPFTUf3ZG?a=S5BFGDd25Ac1NH5],ZM>M2EV+5PKb?E
HG@?BQaK3)=WgUUU0Z.7HPb>DEKD@_HAI;2MB)_>#Zc;fZ?MegADcBSS>Ie^<B_&
E1f[SbMKL,0]L70[,W+QI2]0X99?V:7U^&-9YYTTaDME&G<25OdZ7^RMg#.@d:#>
LR>_[T:7H1cQ:-KD;@Y_W[>S4N#2F1@YaM.)_^,)RYWbQBF(Q+SCK##LR5VJ99C:
:,JdXg]D][\[1]82dW7Xf-CCFOa;Y+8b60K]2F?Z\1->cGY<=0D4),WKXU1-a)MI
/[c)C>AfE55TgLWM<1DW>^H3g:?BG]QGb^cBWR7M&aM]H;]XZ7C&5>?dEQZRV]RH
78AI]8\X\<Q)@#I.4;^:ZL=g7BCL<W7fBcU:)_QDO8I;C-f<LZa#\9O)a0f.:NOa
:F]/A4^(::#LT<SA6>L[aHfTOT68W/6N,Y@SWEfT20W8#O\).QbB7=-.=9@HC+CI
>Z]T^;4DE^K1IG4OdIb]>b^Q+3]#O8(fDP&CFa]?_1Ge=^5K@9bUOFQ\E<I,HW89
8:XV@E4=\eeWbRG=9G1FRIO>FR2P106?\K]RDIDPf.Yg]L_1(_98dSGM3DHB7,JQ
E1==41LB[&:1X58QI8.D=f?[]YM9V6G.[\\g?d)[^)SCA+@Xg)E=GE+0\cWfcR96
]JB.OOL9S?d9H<U9]afEW0+5I5U;;c\&+BTY7@c766K9]HWF@d)JZBH=b9^J_Vc<
(VJ#.)SL-HGVU&71]_LCfO>]3WKC0_YW(Y.)SDJGbWBXAFP1^ZAcEJZO3aVe_B2F
R8U7[::&N&-;Ze:=C<4:fE>O/+[3eDNFb]SG(S@E\ACW\(\GUeg#BP5]fDBP_BNA
UL_Y(_afa3Jg8>B1_P^8bQ8JdaJP.]+L]@b1faN#U+YgPY[Id/.)fUDF9M=bV#_S
:MGaGX]3/EOB1)((e79MDUb<\DX5WP@\aATg-,6[ZXR6c#ZR[dO0?_<N[e/?3#U(
DEU4Y]@_f>J1U17Z/a3AV1RX9DV,JFIe58K_J8BA,4A2dR#^DfE0&^7NW#:X-Q6:
9=P9^-S2=)aPVZCXRJY]E7B;>;7M3:XAcd4bg[<ZDPL\8ETUTAKS<?G/>=Z?Z-J8
I4:?eA_5=.g0C8=b]Y87.HP//.IEV,>#C._Z#=E=[Q;R5=C,ET\^?O^=[+.U0V7^
A;QIbJD(05JH\f2gTZ>gf?[PZ;?:bS=;B\-&>5E.5DbgdI,gKODUZgW[G0,<WZ#V
J#DP3<NWc^V-L<CbX\Kba.6gI9(fT#^4R[19&(T)e:0=c^1\_Q#>NHQBA#gEXMI^
-e_]MN6X;HCE-MRW@DO^\-^WY@C1GOV88Q,OW=Ba5MEAL70<aY5T6<[9>2M]0>Ke
==;V#4;e4^3Va0-N2a.8#/U9fD68AMT[e0GOTDE\[I,M3\VgICS#A<<P8(S#M7dB
;S/ODeS6[(>>#YZUDf-^DBXZ<Rg2+MV;aRR98I,FGS+Z3/<4Y^:9fTWcOPM9A1R+
04A[b_=/[),(35M)3f=@Ce)DDRHBf.6&0Z&8.J3;PL:&LdL,M0<E(;/EUVLcU((B
W<_\6M.Q2Qgb;VG//[eDb1)7?]KbS5FKD0C&_S7M_/\0-/\^VZ)O)DS],9/X[A&&
DIFgH@gTSMWY(@P_7ZQL-V0F-0eSBDI/]=1D+ZE/KBf<=OX+GX^Q1>^;[CNZ@<9K
64IG1#gK.A,3;b>MMCEaJ(IS^4HW&e^M+a2OYBeI2G26CJZd,1II3V4H_;U:S]UW
HDJC;@8)QFJHQS]&3\dLB5/CT30/41RA8b5U>Z:3eSWO5[/LPSX2^3Q_3^cK=W>>
I:7ScH8dG,Z=B7(<bRNUY0X7R5A8_S#;d#K+VF@3@OagK^E8[Ab^fDLO=QX\8?0E
BE>]//.M/8:WFaH@f8LU5-WA<?-7ESK0Y1>:3N<H>&BJY<I1.:EfM=?I8=^F[S0W
[PHZb[F)B,#2d;U;[C;@3YE:L[B_[1YU>RK.6[M(;P_E4<^F,#,0_D#.(FSC]4+2
d3Y)?+ED.CWcCV5A36M8>3W^T8-J<LZfGLX^[MbDUBEf&:W7dJ_O1C)aOD9c)&]M
&03=+?f\G@M:?bJYB2##MFO.X6e_JPQG_\\CV&OHEO-g=+_D)_ZKgJ0a,06=\;16
Fe?eZA.91cIH696Nb..)95JK5FZOE:M&+R322FVW4G\VWaUU-3#Wdc@H28G#=)0[
Ta6\eHTF4PI+&&e;+4_KO[?5C7^Q_7Zf2E0TQOTY8=d^GG:[W6+B?\1NN37#0VI,
VVeNJTOV[b90=C_<Q;Q.,GfV@MS=_T,2P__INU00.)W/L8)-^;Zd=Q2<JN5c.:EV
7//(\Q66.I2fHH7#N)ME<H/Y?5XH+7.LC>a](YR0Ya60Rc&8TKb:T33cE=X-O4<W
YI^.VE\SMOc;71cCBTc(5XTIX5D(dH#GIgb=BR67XHKgINbFbK46>;B>4YPOYaB]
Tb[9b^UP8W_2dEEGa4WLD-YIHN76\33gXga-,Aa.I]/5df#6:NK;N<0PB3d0DJV5
:6BQfW1[EO>7:>e9&=LGN\O2D4&CBUX4:/8>4_P&:ZFSL8TV>cc8f[VX1Tb:Fb))
cK=1<IF7M4DI0Nbe6^O)HO1_M_NW(Eb-6YUJ/76S@=(FJFFPb35SUeFAUS7KE-Ee
\@RVQ6NKFJ8\I6FWac,S[KO>/4bK;KOS3TLBAI)b)87/8]\??WF+M-#6RJ3=;XA-
PBFPDKN_gf\gW&6-5D_Ng4YP@Ee,/I(M)9S6TD;I<-Q+M44:AKO[F^/Y125.R33a
TT?5GU,52B]gG=8bDTG^a2RKNVDeb\aHKCc#SDI2LZ[5,<68<UZ>PZH/QEXcd7=F
WdY.8P-^a^[_T:#5(0_g,8WN)9&^^(abb_LL#VRI.WFY<8LM.0N@X]N@5A2_N)gE
NPd7B9&\da)VK=A/-BQbT<P,XO3^TD\NOa2f.YAVMd9,RJ=FQC:>&;dV9)0;JVIU
5DYEC-L,A=-J#33F>ggYO]C>cPFZ:W@;,4PE+;<g&cOS.e35[;^2:Qe9]3T;X..N
_U,>K/Z-@+a(9=ECL3,@Z/(B&+KH=]-?>d;1a53;UF_R?>[W6a,;=6=N_<I/d4+2
].6HDY&2d?1HD[&dFF8_:2A,Cd[<8E\2_,AWI_6SAb5\FDKY:E/728HC:K,75g];
/dBP#(U4E[d>Ma?Q6@Jb1P1XV]^W&D]?5bK56b29Y2;JYEQf]@8^K>PT3<UJ]&S3
7b>H.B4/?8:U+;U)PZIN#EWRV(49VJ1;/4BXMPXW[R-3f^,P&D1Ic\#S^;886DAZ
fM9QWcNSZ97JO85=+-C;M-OJR=>#Pd&-7)18M45),+:fdcVF1&+)OA125B^R-Q<P
-DaKZM)Tf].?IG.Q?.;@=OK.AY[4PH=52#a0.c4F8?IN01[8-,VTDE25dQU,W&VW
D]B_JMZJ;.D9;5[7d;<e#;B4QW4:WH>FI6B,2AeI92cdJa=0E.c,06cP)QONQ=(Y
Q/<(ZE1++CF@JD=038UL96f:a:/=bEH^>g4U.AOf:A1b(UAH]Dc:0@(/;XfGV@XI
BUg.<\Y2BUR^^C,:dQ3>aCMBB?#_29#(9KA4,]067eOM8+\JZd_7T=B^:b])Q\O]
F?E9_PLJcEd?Hgg#N;dE/_2M/AFdKK^K/0>-6(,2(+6XU^.D]c?;d^)N4&faMF2?
Z.MR)bdSU:FI106DbQ9TbNgYOGF.(#Q&6DV+W&<AX_,b-JC#RM5HN1/CECe_EK\[
[XLUGd,L>3Z0bC9?MKS9\D2@Q>XeBASU6BCIgI?VKf6I<.P#/A0>04I0]eN+D2X@
DZe^+aL;a+1GDUOWPI\9_4V[LaF+84>:fK_e/EAfY-NJa2(:[NT7&_UK5Y0C+KN.
g]ZXa^OO_H,Y)d;gIOfaAARNSY,B;]c/5b]>H5(LHM#OCXD[]-9F]TMB<U#cXgVN
80U&)GC5:2BeSJb,KY:-7H_0L&-:G\>b,Oef4bDWJG<L-GfXIU,OF/0+4UH7=H@Z
Q7)QcYFD-BG#O&6Hba12>EWf31W9?SH+HeN[Ogeg61HF)6b4ZYH/<_bR3]5OMU)X
Fa,RQ9Q80eCKP\CFSge=673P(03a]_#Z:I-Y\#&PBOZbc0X5.6Jb/dL(e;.0d(K(
\PZ#FPce:eJeMT7K\.),,a&4a@M)cO)UV].aA>W]:1FYQ+FI.TUJ/^C(If3,]<.?
#826C3>FR97fDa?NJHZ\@)QUP^47cTRFa5]S+_:?S;c.?]FdY@T;ZcUKIJ8&^&Ce
@0+AT\^(A)gNSI2JA>+UXcO6I5-SCT.SCIgWb8\J\+(B^HE-WaPY)<E(=g8+LH/^
6/IX;@#J<-3OZYfAQ0VAb\a@7X[.K#EDYE#YaTT>>?CPf)A3GKCDaG5X>#;(96FF
@4N,AUg:\C[g(?MO&RG?Z@HX6/<#@&+BQV7Y3g\U>+XXQ5_aM(V.XPW+f&;ODec>
9WfPD>KeQH/:LN27D-#VOP=\RK3WOZ_X1-;Ka/<X_:07R:B2HY_Y[,4]CK,Jf2K6
)&fIe@EE0.B<[_GCPU:6T7P=M-#S/&QQE?+;L7H>[X6eK;<F78c8K7,+&[R#_e^D
&36_FVb_PP[gH61?;J_dLdLgcaX(AO62(#QCR1=gUb;:4ega9M_1e5>2H;E?Edg-
\Ne_J+E783Z)9g7J>\/:ZagKKQW3a;?0(_A=TSAORg3g\JWf&Q@^(fKb-KA3PYD)
b.5d;,Ud,G;J/9N+H.O1/GI_07HVeJ6_V=O4@1.WUZ)J,,PH7NcB,f13g&5<WO15
_V>]IG-I5N:K?>XMYg=Y&RD3W88g(^>,1VR?_D]&8@T(:_VRF>>D>7F@(G<6aLMX
0@UD>K7;BL_]46(OP?U4;Pd:UFQ(,&5(O\N)4N(-UW,;2S^>gUEfVJTQ&Vf-b,\g
ID#25(He>7&=&&9I1Z8R^e>.&e1(b/J3XNXF;L,b15.X,UL/=1/6e&F6<5gY-b=>
E=VD0J-W<]8fUC259(V<>0IM=:(O5H^U4.:e<R_CLD1eYY/7-f5.L;XaV.,VI;bZ
^DG_A3AI_>Gd?]._a#fAF]=55;M4@>1:2QKR4e;PL5EL/?<9K8)QfDTT/e&<HPX2
_J#XOIVJ>bfc_I91ORFCW-.H18GJT./]S[g\.Ze<>+MIV(ON90IN;+-0LD<g\U,S
NaaA>S@GX(J1M)RI&K?);3d1,@R\T)B0SY_8KO=.<Y8-?VDMHG8^?.aV/Y-_E.c1
2BWW<7AIAQ:aXY])I\HZ(^C<]?/.<:X2F9cYNI/A&4(-=4cDU32MdV:9([L25A>f
f]H\1#[RTdZeLMK-gZH9&,LXB2[Q/9&L4O#51d::L.B(ID?NW-IbN.@XKI2dA?-6
X,3G(U-YSFHOQbS11HV(>^bLTEX[a;,>/3L>#-,NeQT_A@3,J&CF:,70J(DZf_:#
=LG]T-,da^-F\f1_S);?-KY/:@RBG6VPJWP^T54Q?6aJe?fK#JTbQ&U9<QGE\UEH
[_c1[Q#9U>aX;eA0PIMS2GfKgR3/C+J7/WN6;V_3])-<f1S>C:SSZ#<O72]V4P8a
.bbaB&Wa:31(DW0^2L#A\<Z?PLPeRF=[>7L=B84T5LIeELg721U&S/bI?K.3Bb7_
+)BaQI/QHTBKC]#:>6TCa-;;3<TM+IQ1CKC&YQ/e+3S.JL/5V4Qf66^Q=/-S2VGM
(gb&bS\71-f^ad3aXT5_]UK[CJE5D#9ff2@(_7:d2J);H@>)X+H2CQFW664V>7bB
R@Y1ZUX_\e;GG\+fJ?K]5Tf,59\C\GU>BW>]?93V(aAWMg(#fTaf8V6MeIV,cEA]
WPc7@TUXWBKYNZ#YTQQ<M1a9=.D52BbM_9FGU35W\\_DBB@dg-\]2>0):X#N\8FG
J&FJ1b,J0T#S/H5_&JeF<?&7GM58+Z2)BJOF8#4VNGCI+NEFT(N^7?0(B^/MSV3=
7^#\UTHL9Z@3>4P(MNFO:-=\E[_JWg#B(YI0?Ja)[)OU8JSUI1AeXKO#EPJ(P,+I
34B]#^\bBC\O#]=+,_;;1abUG?9O>USHa,2d6ZcGe(CV[Z#BQTBA1L02R2/>S.fU
a:ga_X7XT&1P2VfQDV>#S?(b9UXI<V0VZ33,:<UQQbVVG$
`endprotected
        

`protected
_JH@a(/BDDVa>:ONB>HC:SNEd,Ya@)fC];GZVa[Xg)>6).3YGe.+2).,4=CLUW-1
(_E-a>Z8/YXY_gFJA^=e3=ZO_ABa=#)(;$
`endprotected

//vcs_lic_vip_protect
  `protected
3Bd2(a[RY#g?7:>1Y&?gZMHL/6=?5R+EVV?#Y9/fVBV7[S;0DJ9+3(2+gR3BaQXa
F>;D><\A;TLK;:[PX(W_HO2(ID;;V;,+:SZ&cK<WUOOD]W(X\E\d/LB5Nd-:[[fP
#;/X__YTL3HQBC52\@SQ5,5]2D^DE92M+1dI@g(K;(Q#UE+^1@M9bDXTH8A_J-BS
VN;V41PWM3RZ=9U0VP<>X,YIcIOI^=MG^0EJ_37Q=ZKRbU>,KN9Ja5HH+KGg)ZK1
GdKeB]2;(15accBJdHES[JN6cQJd_dE^.#1456b;4Rf[2N(H]Ig;+G(C,Qba#KXC
8;FKaA:WCTX@K6_R=E)0LV5(.e>Z7.,CC^S3AbG9(W)#Ab4\)+BK;_>+Te/OYA^<
A#8&/_VQD@^Bad0X_6>dHPaD:N\S0MHVG<:]<;:HPDf_Q^<VH0V#=JS?P,PH6KQS
5,R8VJgE7E.f,UU[FXI@f+S+2[WN5@2G:O\A=Vca5P@P3:)->b?=IK.H75#DPP3M
d4J0I0..S0@<[-4?WX+/IVUSYa8g;EE]e[eZ:\+gH\F#bIe;1H]3RC#FZef(2d>V
+\(_d/6N#H@OG?;Kgg:B6Y.8\BfR-/@WfUA?5+3eY2#B(I4U?9Q#g-;,][CXCb8V
(C7YM[2[BP1?PQd<6B=[^OR9OJCOYV2]N;N3:Vd0(D_0BWVeO:/c(T.KG9D7QNEV
WQc:RAaRJ],H2]ALD2Ca\PFe/ZTYC?\(Z;-(GM<#_NgNO>4AMFIe@9b65GW1Be-H
:LXNI(,INOP=),J?GZO/H[,I75dQZ#e3=3^1Z3MA1]2d09;:Y@^4d[.G7HA^#Sdg
BY\aL1IL+eV77g=BZ#/e192NdM_9fA:]fb/8A?\#DAb+&6Q17X2)6LU1GLR]KO9X
b59SYM8+5.C(5)6J^Zbd=8)1cK:5S>-J-V(SZe2MSU2?@^Q.U9L;SGNUS@:&Z?FL
-+BC1_@3J7-I#5YCI1/C9?,aVZ3>0YVNF3dB_egL:=K2fT-NR^)KWYUWHY#d3^+E
/45ga#OCZN#g-B7F&K:@I7U8NSd72&eOHK(R&;LC63_UNTN/ETKO4ZeKH)?f<ICE
BfGS<>4P:EgSCLaMMC3V#E]XeXCQ-QTcaHD@3A[1NQ8@J^T.K&eG?L1PdF<g+._3
^,91YUNR^faaX.:N3-X#R9NJ/4N3+MW8X8/S\EG47@a2L4J\f-<,^3Vf6HI>^(MP
e8ZQW,^MAGGH9-X6KP=G;;\(44.J,6A8?/CbGJ>I0V;A;[31KA90G]BEL@67KA[E
f3WaM8BH62T7GD#)7AWdD;8\RA::J]bfWW_Lb+.T^5ae7NT/C/LOTVb[c4\SdR.>
4?=C)]_?T\WVYIKD+N5@gE([+;]W9cO6fAdAFeeg)[H\eI4a:@Z?<J+NT3.>=_PU
I;R@L.9;7;]b?4eG55)0;P?US^Y&ae9-@U[ZL<P^9aHYggRFHfe9XFQH<YLfRgL-
W_bXBQ-8c_C5DM4PeA?(++eVEC23:.SVcXD>;U<M10GcWe^+;@(]#\-+B0,(0a63
4e9]6D4OL^a8H^QZQB7/XedX_c;C\Q:^ETaYX,5@VYG^L56LAG3>+L=:Z);O@IE^
(;S:BBY3d@d1M;W3J.+K(K_.=&0#LK1Wea_9Q#XJD:\M8QFX&A1bAG8NaR/f>+<Q
SXaa@81T+RK1OSBY8EY(dC[7^#EOH7.-MICMIIH3f^#cU-M8BZKTLF#_(4XP<XDX
IA#OPA_@2.UDGS9@P7XU;+bWgFZNVA5B.GVRfWD-4Pa8[QN?.R&cG9GMTA9E.A[\
=eeY7dF3&/<cJTa>BFU0+G+XQ-40(;e_I&?RX>DNLZ/]INF5Ke5BXVWU=2@S339P
7..+-5RGPF-JC7T,)]a]]V@ED@ZIb.X(C&9>4K\9Z:cB_<TXS2O?^CdVIMFfaG2;
3+eG0I7P8\G+Ze;4-W-1WA)1@(12O,8cNCX,4eKO0G?DaK>bO)0N]G4T-#LKP1Ig
/Qe8D,3M4UJ+@/=g:>a9B\WU>J/_=d0)_0Ug51HJfE>Z6IPOE:S([IXV;G?1Od)Q
(S6^/,6-(HC?-#])VF\5K26^gC&4>D#HO=WG3>X)^M\8K<:OAJEK859=d,Q#(3_/
GAL9),Xbb8dOB<FDG)/:=(LZ6<a>9H[H<0#\P1DW:?fITS(9dRU-LDN6A\\PA[]D
H207eO_gBV+:[8PKAPYB>_K68V]TQM2G2@XC&,3U<-1]&Y(.P[-&Kf<GY:R1L/G&
_Xa2&@)QFVUYKYCCaN_>eVS3cMYQ5,bb9;)8LgSV>A3QVGV<7THQ6US3CAd2GFDW
ZQ-()]<A=Q[-LWM(,9Y8&T)T_=2b960CMJec]8/D>GT:^MD2_)U\-aS/fDKfb1\M
,ea@]Q7HMgADQ+J3UXHGTU(_A;+bS&FeK#gFEVE^>ICGQGZXEe6fZ8YEDFKVGb[3
SRHB[0E]a8>Cd<NL+4cBbA<00INE_cZ_X;YK[:e@?PNFI^WDN^P6KNdI.71cQ95O
=5MP)JFRdUED+e@6^3&P6(KZD:MA_+CdA/[G&d)5Q.HZTbZc81f)D[]]A?WA,6?d
;T:bC&)70)BXM2M@BM:g@4P(F9OA7/\;07MHQbHdKN-_4/\](PQ(+502,@P(?LBR
e?fTf>A5#DQM/2.;6K>Y(3.gd:ge:;8Kf@+)J;>)9I5BQYVbBCd&N5Jcb#\T32dQ
3g(?^?-S?+)?C5Y?XP.>cB\]@]db<cEI=b@b\4JE5Q](2?0fgf6\e+/+(&11-MaW
+>1H-SgC1F59\+1T+Q[@bK5U,We2Q>(,g+Ic7[a9d(S0P1Zf^f)5a#\&MV(OK\XN
(f3U3&b+W:+AfE:2;6c&aB]e6<)4f#@N,&,MNb0Pa_/C:QQMfbKHb8H/U00U-6KD
W1f>CYVE))@#_eW\H1H-)[NQF[GWX1S#R._IKHbKSMZdI\QHQ5XB:TOgDSMA#]]=
67T/K27dRWg=)fW=GFWOX)36.5/Z_W[BVZB?@=+_cI@X;(:F&RV1UOI6STR#A5QJ
J^.,ZacG?#5IN078+Sd3]N8=SQL&:gd68/P^,QADDBZ+=ZDWWfAD78A+H-<48352
O<4GYG.63CRRCIJcQ3_,g8>\2a@TTHO3G(=J@W\_Nb5:0K0T/cKN2&TdYfX5MRN1
I.J/[DbJFc-&\bI&^]^cPF.0\@[+PgDgdT)-;PH05N@3K6T9@[5d;<1U9K7L,53#
#<4c9.d\9cXH;]?W)ZC1F\UEbGDR&2g_VPAEXf36dY3DDOG)/T)7F]gO/4M@c+21
KZ]8L.MFD9aER/#[K4Q@c^>437Ba,AXJ\V=+Y^Xc1&I:@?98OJU_YI>&J>TO/P(J
G3GG;QF2Y5_F=BHZCd7.P)=ae_LY#NeHEN/Q]0[YbNYVYTI5]H5g[.:4R\Y#TBXQ
7?KIXgf<>_B_N1Xca6WU:5RQ-JPOEKK.:D=Od[]8)/AI00d.+YRP+7L;#@RQee^2
YRbSC26dZM<M^YWb0OLQ;]cP1/P?ZKX:CA_&>AY9<,;>LS:4<FWO9X1__L3?C9<>
eb?Q(,_MB:0A]3/GLcc,ZR?A?KUCL>)V1Y2MN>gID9?,V?4YQ<@V(@KH0#CI4U2)
.,X,VY0(Z(Z>+]1CAc^=]\FGA?,O;0baVG\c:\L6dcR]?-cB0WS1Q2EDSbC+^c#&
MGVQ0b7<Pe.;7L;1UcJ2R4[X.L63[7b_WJ#Fc>^.ZX:FCT+,?Q6gR@c?e3GBOZ<L
gSWb51]YH8W](D?F-OV1RB,OZ/NF8bcdX)U<[QG9LM+63/ZIR/d12e8?KSL)_OO;
.O@WUeO+DSY2/Kee>>++dG\<++R]ba+fN-HZ,O2ZE4^H;]FHAR:f8SZ9(0d06I-5
979GX]O+Bf/^I7S#<P5Y=EG[R9]G945b;KR)O(KP@RG#?7JC5HQ&T<5^H]ZC+.Q:
&8TS2KEPZE,I+.>cESXX2XHB;f.EMA9=N81dHX_O?1K0<)LCE30DeEbI=Xc;af#)
M;SKL(Rc-]]-:QD8F5)C[460M60@=bJZa8Y81I8LM56E=QL-#ad)85BUfE[<BFKZ
/NdCB;ARNG3-X]DO]:S\-6U0ERO[7=e.(5<;F8V+7[bGMKed(9<7&MMc#5P,40VY
X1)>?4>FaY^D^:=39->bDWVY^HQ3Q3]B=.O4J-8&I,^C3#I,Y[>5AGb<F\[).ff9
;=Ha2P.R?^\dAbRCHN5SQGDTa8U:E]D]IDW^&R?/:bO7=AcaSZ<b[b(P+XHME1ZH
>F]9H4E(.bG+DX)F19HORaFcEOMaBL#@0;C8B7B5g\)FUf.O,\6#>4d3dc:6WV5Y
W.02#2[G=LA8+Z+Oe1dWNJU7^:R,.E5GZf#/UH4@3TI]CZ#TP80>ETaa+/KPIL]e
=H,#/[-L^WD3F<_)H95EWRe42\+Y2R_V#QGQDA(8>4DEJSG4R0Q/OM))(VG<T9bX
MM:cYM<aE/1KR6LGJ62S,<#.:P:JQ1W)Q?CDJ3KDX>3J8C@[WM=?aM>R(3^H(E8.
d?D4HB:_UL:]8S3N=R1?#c-gC.JQXG+X>$
`endprotected

`protected
?[[;=8:X3VbP?cMWG#g&Dg:B:7F:2dfCAgQNBA:>@9]G[?/JfZWb0)g[00_Z:1^+
28W/T8<bV?e?QCGN@EDQ]]Z21[d([gN]>$
`endprotected
        
//vcs_lic_vip_protect
  `protected
QD(.\KZUJ7Q/#\?A62O_BC/bQ<]f<I6eU;<[:-FQe0G/c/L-(>SE-(]&fMeQVD@W
72T,^5b\E7/+:)>>RSK=946LU4f>/IPg=<bNB?_10([UeCLN;;<,1P-dIL;&:-5.
@Y5=MU<]ZS+JHEM:4W^fQDD6?U)=g5V7af]JDAUG#c?(Hd-fc\0ALZBPYdE3fVPG
,(Jbd)<43&NfWVEUNT:@^W2U[+aVGONI6U.,X6^YdNL2a4<JNL4(+-eFY8Gb6HE+
2?_\O]BVLTH__^MYCG#e&Z6X\FL5:0gJ)ba+J&[K>e.:;B8L<\Mb/&#2(;30RL0g
=U@FTZSMT?#g4U43e=VUF;B1^<MR9BbL0PVeTNQeOR<G(W7+8d&NMRP,gK-0>(_R
I8HPcJB5&f?4\;=aFB(d+=C:>PaW7d8JW7H@=c]a[.#LN]4N5SD6+#0+1T3fK-7/
9ELBCM47U]]a45-dR)A79A(9OcXT</=c;@Q4LEDPJI6:-,NG5K<)XaXN6ED088aO
U]6^^35C;eZ(+]\aCJE2g=/E]gF\dOAK7^2ggcYc5Z,Pf\N1Q#AQJVIRS2-L08W\
9,A:a9S]3X]4f_M\>d_?T6SSYGLO++A&9a(LID_U9Q@Z,E=9T>P^^XAI+B<&b:?]
Ec&:]WE5BZcg[gYa62@NY_,J:fMU]SU58@]a>V:Zf?GKGbBG:NZW@&(P^V_-(486
gMU#XJAIMFF>]F?-(#f2HCJ9@GZ9+F:cM<[KS@7T:T#76)+0>PS(f>-,e)HPQ(DL
>V&,KC>3DQ@&8MPTH[;?NE</;>CR;.6)&0S-JF62BQ;K#^EHgBaAI>TFK-gd7Q9f
^5GMYK\A\2aUDW^>M8Ac,S5Gg#,7C2,2)Yg.(FS,_-[eSL/:@[+MWf@Da^E#NKLU
^5AK@cIZH2O+IU8Z=C0^ZeZI?=b>QVJV<9558@-K&VBY@9,,[N=137f/(>_CV.-9
:TPgcO#Y)Z3>DJ,[fL]8J#f/[Z.(Xf&B\4>I48C254XWf]aJ/@[3G/Y._PLI=MOH
-U^HU#6&[1cc4A(a.1NPQE5P(778G7:cN\-8QD@V9B4LBNYcKefR1PUSeQ##Q+H(
=E5d,Y6Z=@bVGX>>3])SPE1=c:@86HO?TS>aDR2L6>1N\fG]gT<@Bbed=.3MdJM?
:F\[2Y4fcA^K]\+IbMVY)Q__C,PeY1V805-eAH,9HJ/_+_PUIRMggbW&W8eS8]3b
#U7)4T4;fCH>R=cG@GMR0,G45H^gg8AIFNdA92[W^L14I/->Pa^<-S0_S7\KN4g4
>PO;gERO24;bFFK.XM]1EW.I,PM,=&7E&0XZ<fcRJ)<=I[63H;e#:1&6?)\C6?X(
(IF?f083UQ@G^_a?^6LK\ce.R8Z];=+)LF5P.)ccbb5FHN)MgO=PN<9dRFb\,QF=
bfFK#T);G0,,Z:fP(D+8AKRKb6gG\B>FNd63Fd.1J/)3=QJ?ESC)_a8QAK0=c^H.
b)+L8IbY.2A?d#.7?4.X5HO?LA,/-_NH:d)88RC0U)b=<c22;2J@-5]A04D>EIO.
/R-2b#e(V)FN_=b4-c)-UgEUCR8TcMI3>Id0:FWE=g/.2HWY4Aa)3,]eS(9]+(ec
P>g9\Ne,Se@CX#P&]CIX;=@NcCA:;TC8f:Ka?@B=eUc>DUS[]eb0/#;QB_^7&0,c
H=G^X?8A;[gPaTcJNN0ZT(>7FW&G)L-CXeNNEBY+QO4Ta44<0d&UWNX\g\NYEYb>
>:0eDC\RYU>f<6A7;a]/1:]=5DL#\18?CZg<5J:&Fa#fUXP3=;[L052<C:Yf^b&M
,<X_<Ze=GbP44>ZcUN,O-M+3I73PeZ[<:_N.\NTQ?Se^^^0dR@4&QZ(-+31gBN7B
1Ya5(CUKM]dLBH\[_&M?\;b^aM6ZdGP02a>3Lbd(?8Ce4IO5<W?1E&J8SYLNE:>/
UA<4=L03JL^VQHG-Y.c?R:aWZQB>SAB->7#>6TI3)e?ZJ=e[XH5JP;KB5^HHD,gT
76HEgcT,IN2+<B3]/IgPHIg(JA<e[DZ03X2eE[[KdYDB79EL>H#N?_eYfK2WEaZJ
]U75)6BV3?P6J\W:DY-Rae]9S7?DKQJ@eM+Ga>O:H?+Z6.<?NIK]Gd;3+We:c1#@
0B(=D6)CVHYgL)XCRPGC5b,B</^K-CS:3MN2B7.B:MA9<8HLS@OVGH\Rf;3#).WB
-UYNUX4Z#FTd4&f+<\_T/T\#QVJ)g0aZMZUU&&K+Kc(bZ6S0(aBG/.X1dYOO-NZ:
dTOdTGHbZ-HXMZSNB[[Y/7gHcUOW:X50GgeL.WN7eX_V29Y_B+((.42THT=<O[.B
NWBQWf(OL\\.<R]Z:_KUY3?@YU?8BXB-WXI[QYUVQ\2.//-0A@ETeP=aP4^&b0De
,/Q?2)WO]AHS)N;X;b/Qc=)8J,DEZIK.L9=,AW@;]7:@eNeMU\d>3.>Q&#MA:eF8
6DAXU0VMK_TdH>XL7RT+/RAIW/@^//P_FRK8:5O0eHX05+T603.[./V#LAARV+,H
N+)Y^GG\W[QLf&fAOVJ0).P57/eM5I@9I07^T2WMaOJ\I/=R8A9_M^g>#O7E:e_^
3IE8#VEZ5B\EJ/9&0,b0&+&Xf2W)#(c5V]/WG_c8gZ4P(8#:&54XFbUYUcKWJ^DM
2PMLc9TD\;KGCQMGSH((eZd2Eef6JF)H#5-GaN:Y30,NVA380AM4E,ggWR=:dF60
EUe(IZHW<.WUKc/MZ;A\b(eO.N2LCHGMQ2RF@),6]^CJL:@(3;(?cN=T,1K8L^F[
AI/Ng_8Q^f?Q8GOJVZ?SK6Y(>><9XFI0P03)]D=fT[Z+L+&gW[28:4NIY,54+YgC
=IgI,G;2AZ?_)>U8]E7_F+38RGM?:WSIc:1_,f7NB?@A:J_],F#&UFcLQK<GdIUe
1>>&&d5,.Dd+J+b<XOaM49_?Rf:;cRQbU;)YLYacO351JOABd_,U1&-&EWE)(c;O
J?;@O.^GL0(eGOD>aXT+XWe-X7d8)BDCbNCa(1J<gfWRX:fPFQS-J#DfYe033P+L
[&\S^S9[E6-..,WZ>@(d05O^BHT?SGRaZYF7e?fUe-0L+8DD+=K.N2SM0,_KS5gP
Z7Tb&G(LMe8DJ+C.\536ECBEO/eYAYRULYA=e.V2MU47?g2+#JS-PH0>=8aaFYcZ
VC#,/5_a\,7VB)+f?QIWHa2PXW##0BS>JVQEP^/K4<1Y3U=\V0E@C#d=Q16963I.
PBDC#?N;^4[Re;&Z^>R8+adRQ:A<d=M_SE:ORUZX1@AHQ&8bQTE&]M4,+f.f?6fS
[_9+E5d0,IKZcC(&T<P)2P:,7,,]#d7,0=J6CdKWaFAT.+VZ7CgJ461FeES_BX]6
G9KJR=]&0g\OLJ<;_gdQ((2EVX>SMLQ&L(57c50d0cgF.=V+,<H2C,_I\+U.4&NF
T5a04Wb]PZ&.Nc#H:;-&WT4@WcET[&LZY+b+0S#c-[A7^LBKZ=[F7gNJW+&26DbD
<N^TV08/YIFHTO4a&BG[8YK-?SJZ+HRBT?&KLTNP-]R[\^?;0Be<:>b9<-f?deC=
.S6ID+P4K&@XT4@U5G34Fc3W&S>,U<7[>R13L5#C[=c++,e_6)FOZHIC95C:.dU5
ZbFG>4,75[E+9(U,WbA\([YfP&d9EE_KAGURef/,H=X6f<;2#e23>a.2AX,VT3dJ
ESXW/f^(9_1[X<;L7:@,#_3PNUFP<VA\OYgXcSW,#Q/6fDJ3[R]N:2D=#H@WSLN0
Fe9R?,:0JB.]V98OOYAE_8]4MXfdRe&KI1L5[YES5a?LME<J)^G(;/+)9eJ+TR\G
4?QC7-b5K>:PH(JJ\+RT5<,I@X260dFRf#d8H[G:.KAGJaFL:4DB-a/T/aY1HI?:
0a\gZK;1FNC7agO@3a(-^2[d))CW_YK6C,]/N]-9_(K-BQaMR6&\>=L8Q[#CEbA@
)HQ(C3@>X0OZERB?IeWJNY<:N<NQPI3PR^40=MRRa=CL#D8eTf#bAaG(dXg+L+5S
.T:WdWOC7,(03eQf@bM&[@g9R73g7e)]S#+gO.=#bURM=#c;WO,V4P1/<FHE:W?F
]H\gL?6&LK=,CU@C;7:Aad2=bX34aUc+M#L;aeT1[F/HY\B_HIC9(Dd4G@([;b8.
)K(59K97WD+SSMNSfKJ,Z)G/+V:W^1P@9K=QVCSaR<GbH#Y.1RXAI7,.G7Lg+_7#
&VfReH3c=d20gaY2f_>\@MNE<AVa^:Dge=DQ,2Q&JQ&9S6JR-OaVQB(#>C=Ya[0;
Y51B(X6fF5V</[;f1RSY+&&M;A67g-2+eg@1GZeCZE_X,3SC;Dd,R6+8cc7^F+A3
?X_\a1<8]5(J@EV/J>GU)KcLcf(G/D]N/:JT]+Mc?I)5.0fZg2W7V-@Qdb?[FT^e
OOIE0S1L;<_ba57TPb4HV3/^VKRg^+7dDJM0-(5CI03K)DfGFHU)-Y<f.D/V:0f@
_f7W&0L_RdFG,5(W<@)K_0V7/6=C0_=H]:e&\W5e4a#^\)U/-+f(T;c:,&B78+Q(
X2)Lb.N@e/]6Z5>6Qc&S-[77e#3=PVT+H&f.7FM^C-PI#5=\Z?UQPIGMEBaFU4E:
H8Q9;MQfE40V^(CNe4>(-25GUUP./^PPV9dU2E#/We^J/4SI(/A0R@U-/XM1#E85
IFW148W/4]YQ+@X0WO&bWN?c,\eF5/P@S9Kf2d5IL4g<V?R7_7R)ZSY59M#HW?.T
CaD:8RQ:ae?Y<c=/00D+bRG8?M=8_e+bU([&JZ0HIV2RA94_M.EZ<ZH6&>X@HMe@
gNcFSgDZ.0]31GQ:6TL[>9M?:/efE^/MYRK;[9-S,a]R+;HB.I_)U#-aLM0B(aX9
JT2<R]e[5N#.,,<=Hc9\H(&I7+d&f;X;G?DX;L3gHC?beEP.Ld9Lb>&>APN_T=D0
/5DD_CY-\;2Nf9X3_3+RT6\)BT<c8>];=O11AX6f3KOBYb::3Q:&)+f=A,N_ON-F
:>;7ZH33&NU<LM@#KH7D>?W5C[0=7&&aJDPXQZH6.<45WZ3.HYZ?,,Nc=NY:4Vc)
VQcJ#T5--]b0>Qc_C)E//3S<#-GGS6fYaSPU(6><,XOU(HY\)WUa\&&LUAcF1<D;
R;<7?M^GTIFHE#3O6UM;0JDO&.Q;OUWY=]L?P6H89KLUYRHVaLO3M.AEM_D#91^S
;,UPId=5RdH2f(:Ne(0KM)7S>8b6Q^BJJ&5(^[\]UW&>4T_HPJK#,/3B^YPR5TI9
\FX[#XaX?<?OfAQ,DE<5gF+-B8eK8S>FGC]DHJ;H:+fKA)XSX5\CG1O<7N/D_XD[
^CSX.:=AB6Y&?5eXNGfT,I7aY6UfRATN^)E1]RU?AZE0/28WVJ<dEU@g_K,<;X@g
<QJbEBQ6N=U(</A?55:ZLA;=ED@S<\@(#a<-_0?=4:<aaZK(8SUYT][S[ZF8K6,.
XZ=YVO><a78F\+T7c,VURQd^CYS_LUKHR[W?V2B[-80YKX(WAR-#>/B=JUNeV&,\
MFbLK#A]>A^R8:\S:R/E6gWb[0(W0Z2=;3B@f]L5[:cIJ13^((dY9?&Dcbc9,8;E
D2K<g6D0e2E/Q&g>eNf981Y;JM&RM->,[Z[217UL/WH#eZ-3G[C2)?)<dS,(;WYQ
:\H>[IfCe4OP6fMGe>U2OK=H)fL2[#0G2M)\X3a/F35ZbNZ;P64/WdP]8V4SFf.=
5DPfQ=dG=[@PW^G]<a(&D7XM@)4:#>g.;(P<JUEad)?K917NMG[#cbDE@e#+WY9U
MNT_GAb-.7S7PFf#W871J?dL7;Y_<d#<U,LTCZ&<-N.;:>C2Wa1Q)-)T88;+eIFH
<O-/F&]ad<feOPbR=A&70\WPAe8_(MeU2X)WHSJ[_.((9[ZgR9F6PPAK(=D=?C]Q
V=cTY#LJMDaJ;B7GF<M\=HGWI=E]M^6bKJWO^EAYMW&X-0)P1N=:Z.]90W,IR4Ia
,26W=HOWG).<)_(<P\\799PR[f:XU)=4DP;Y6O3^A67f9eT3^=H@&1[.1MA5a_F;
RQ1=N)7PeLF0#-Q6BM3A]gM[V_@G2JVc(9fNPb@T+DA?;1?,Za7,0TdJVc3G#eaf
8#+9].]L(I-\1?gcgd=46,-4>QO10T,]EWRMdCE-3Dc+D1;LR@6)+]S#CYT@I<68
e\3HJgbK7\-2U9[EZSH/eGF-IOPVB.L5D?F9[TbaK=/95<?+EY@[c0gN5D8(>DX\
@]LTXISW\/?_?6O0aK<abdG>C3d:,:V&)<58WEV\[Wa;/OV40@Kc;=.M^D,A+7\9
dUALHb44M9:8CdN0;^J#+N4.J4DbfNc@fW#A:5\6\<EX:@?dAK)J57SAFTKL#.;6
=dM7,>O2WW=1g+(DTA),^)88<GDe#ZF8CMW8eWcD._&b28ZA<_-9A/K)I,U&2.BS
@B4=PT]L80&0B[IKId4HeO(Ug\/#?TOe)DWOQE3Q;SeIFJ9;e99&@A(=[WNM>e+f
H(=\)S:3#1??AO0<,B_]Hg+#;EUK[5BVS9gZ^1Eb4CEP<<V>PS7_)_AeU[QOR7\f
0@4gZE<2<FTKcYH6<1d.MZPXcVH^X6/c+_[.??4^@K_ALTCMA?=+/W@J/6Df47JR
[#KXXcbGe+^VO@ZB=.97\3J.FO=1W,O8[QY;CF2:<HK9d[fA/5Z&f>K-b,,U<6\P
]NLADBST<:PA=?/\ZMQ<1Y0&\aU?-5-XH9_CG[<[K^CPSb<D.WY:?F>K0(J@&H>,
#2a6HMJ(48)(eD:<M@60/f&a_ee&&Ke>NS3;.^XIaQg][#YJ5G_14(6?>WMMCd(4
MUP_3:/5VZ6[/]3)RW6,@KK5DcB]^R.c:;\MH8ReJBI<KG,7IaTA52U;f7H7dF\O
<ZZd\F4V==,B@HT#Cbed+/)E-<ga@,W,?Da>ST;>:d15SR7bB-/bfZ5B-;C97,=a
F9?\eD\26C.KKA;MLeF3OQ5+XQ4YE@e)(^-,AaD\0,FN921d<J[9\O3)F@_cLEF+
U:0[)YeK@C6^:XMQVA1_#2:A(][bc1\C>g;VVZU5&ddb/8U6C[GYA2BHN9).HaNM
;GO5H&X1=UIe@T5G+9M.P.K[GU9ESQ3@>H,f:H&^+Q/LK#A=06=c^g:7<#/4g@Q_
)G@M,]44&==-_aJ4I7\L<cd&a+E/?ROPTb2NMa@_F6a8GV2>+@,5ZgNN<&5dgI#F
<]KX&+>G:Y(IFQ9_2ISRWHB[.Y1+gI3:2-DWL-66@=;8GMS7MS4@c2fEbZI.TfPe
MSW:,aQEV^3MXH>4JfQQ-J3?+DNN.c;6_G31UFIc)gGE^D73QA(R3.8[..1JRI,J
cH/>M&&XNT58P7HH4ZLYN&K[45Ee3)+Hg+)\#<BfUB@=UJB?4=U>CG/Z-T]ZBY_2
/90R&1+bQf?QAgbS1RZGJMQ55Eb@\H[7T<4(=fJC<^]F[VGPMPWXCCYdaF-;Je=M
(gV]MAK)GSEH/a/.d[PgV&]&77?5b7>)0IA/J&afI5b,_OT\OT@Kg,aS589.NOPb
Qd0FE-^cWEeR4IDZ1:&P+0V3&/]g0N:^(9aSgAEPDR:9-&Z/2WgCL)Z?6U>C<H]S
G].fB&DH05B=7XUGVQQ7>AX7VZf(#SNEd7aK+8J8cW?_IF;4[E]VVR5E-g9[N01S
DeG=I<HO@9.c>SS)H75>Q)VHC#HENSU;I8+g5G1_3gE8J>T&^b5@8@CdY>XW&4K2
>124L3/A^F^@Igaf+X^Vb6FG][85FQPGBM(]XNI)9bX[7ZDYAUgd>[fY+<VKHEg\
9JTHO/fSb+@.U0H]R(4(_<3JW&NXEcNI1R90WX/2aQ<_:VMI5INEbB?Le\c-gc98
XI6Z)52#P7:O^e/3\X5M[b)+TF@&+=P6f32?>3edKJ]P_T,\J9FS>L;RbQ<G+Z/U
/fTD5\MCWIR7Mc&#C,E[7a>0()aX5R(b<Y,X&2?O5Y>;SUE_PGYb#6/de4Q/JSV?
-L1A[A<H5e(H;X&BQ3,YcQS/2;Wc0C4QGf>XLA>E(Q(F2]2g.R<FL/W:VC&(@Kfg
S8&VU&4-L8?C4abWCGQ;/H,PFC@&P;e4;<<R&8g]:YC?fX:[3Va4cJFL1/R88G&c
Y2Q9bY6F[X_fHS/Uc+.QEf:T<aW?&=)\O-YTMLOdS@,UL[1@S9>fLgf>G5ZL>2/B
\5dd4R+f;-H&dfU7N1U4S7NW-YeF7W7<RLF-6)/+1?49A);5\SL8A+7_VBd#W/==
?E8\NReCQ^gB[(<@6@7]&LRWB_9;2PTAH.a@/NZO,:DQ^(:G5JbWJ\A(T=@2PO]=
Gc76.P4b]>_5>B<]6K#YHc+[Z80P+7b)3NTMK+AQ;Dc#SHgSN[998Ne\Y?4N:4AX
74.K+=d\][dZ;0ME5bO]Bd<>XfDHHA1g@:gP/.MH;Q,J6+XcILZa=QP,8GL5_LCa
2#(UA^F=d5.I+RH#O-?7V:LJ4c[<Z,CT<=e#4/<1&@R5/Kd)7#/T2QN/+VJGPeD9
dC\9ZYA@O232@_gGBe?^TQ#e#8W#HROQYLI0HY:J&.1Bb-;/5YH>:WM.5]-Y0ZYA
W/&BW@9/WcLHAVb=Jc4=_D#>\].QL25<ZUS#8QK=]3XS/]c5X,OJ>d^&@g0\2W5<
RLQ?Q.K-M_]8_6]eY3;_TZ#,:,1867K@CLRU\3,@\@J87eKLYf86NP8;?Gf&g9HM
<F8D<X;JLZXZXR6g0TXXS#[bDgEbYAMNXT=U51+FYaN3WB=))U_K]1>>(4&V?V50
<+#OZR[C=R0^UBcg.8)XTM8/Y+?.[#,ea5L)Q3&OAT?[7=K\^&;(<^?QQ?:eZ0U-
aM12P4SAT4R0?BQ+S\,Y\U-WL(L>JKJU\<MP0L+CcI3\1g/[eCJ1/?[7CI4AVF>M
HUdIGXLP-59O/gT@,9f6FdKQ3]\2#/b.&&?&&/67]e3:VI7(WL?7.M5eB6PgO?-&
(:BYJT1(A5SP;4XZJ1aT,3gOA;O?69AOKGFP1YU6GF[gRF:d-2R=eQdDQbT=##,P
G=Q_-;0)YMWH7_^TM-NSV\g.L(LR:V9]4+3KG949;)IPc<H:/==YW>8PO;ARgS&4
KH?cMF4SWd=He+J=^<_5?7ed>BY8X4AO<C>08bB)KVB])@f><QGNTFP;)dQgOEO\
=#AJR(X^1IIU;g,CFLI33b6(R1BVD:;T1L@@072HQM)NVIS)b2ES<MZ@(HS_R9-@
U^W&K6OV:JIWQF]-KLc&<1^WZ8(g---]8VU5P]>F(>\df6YNHg8)Cb-./=[Dag,2
Ya<P;C#=4fWg,3L\&^-.b.Qb//c-SUL<\(12PNQR56e<Z7ANf=)Q-bgN6Z9Dfbc;
^C]RSEKLf_/;73fZ9Q:\9)cC7cE8LRA_F6bUC=GS^HGI[GXVO:O(??O<fG,VD&]>
BPB16f;3AUeagagIKOK_P4.0<_HCB692Bd>M5S4J)W+R.=G[,@Y70Z\0Sa0HP82,
S^d=T8X,_2@_:B,).LL@X^,VDK/6g=OCRI_-UJ:c?XPd7\\_J3A7#V77f8W>&W\,
^Z+J_QB&PK^YD.IAEa?eW[))Y</f<FOOAd@IAeF>2Y4@AJ_4L3C.2Gc130g7[8T_
S&6E/THU-H&c]>>(/:)[J+f0N9@=8P]eJEe?31LBb1(a(3KV6e)1XWPJT9)\25gI
<Ide=+QQ\b1]SNcX>8NS,?UHG618Ea51LZH47]^?H[BK#^O2O>g0X#G99FV8^.dN
ISE_UJ44ML<+JI1NZ8A7^1?H[A^T_L@##?SIJdR9N.g+&\U40&&#KgHaF,N\7]0O
VgHa7_cWV:.(\O2gT[b6cITa[6L^BX90+dF#+^@Oc)_4fQS>H_9B.69Q5BS/LI1@
H@a,8.F<_(VI9#QLEa(7G(IICF8O_5=J(PP[&5\d21a6P?fN@Q]X#d3Y]TgGD3cO
QK_a[e^9)KJFK2TZ,EgPNT_UW6H]#KEd(F,?0MPba^2[cR5TFGOP4--K/f./cFBX
GUeYP;>g\.MZ2O&_@K<08R(3#Qa#VNU9L=T#/2YTgA-N7041/.&d4L[KC,bW:]W.
TfH@277X2S_0)A#SJ1=MWaP6EI+S91g9^g;]EMZS>9RA)fY]O)a9T5AN+N<[OJ]6
0972ReZb.,YC8M=C)2)K&KCWFe23SUA\_FKHK<8[^@IM.e28QL1JM>D;N:X[;>f9
C4(K:?=;]/g&[aQ>.+@UHC;VMdBc37FM8I[Ba]?bbP#8ATZKE8<4(F^-<dX9F@W&
-dd52C:O:4>[d[2O0ZXa59&Q(N/+):(@:@09LQVJ6-1DWP[+,];M6PBac@^FXA_P
H5G8T=3cVAXSaCcf;@Z#K1OJ#NA4RMgFeP#1>6WH93?cLU^E7gVfYFJC/[+2,9E[
YP,[FaT_TSYTRSBBIZBYKeC-6;5eLf;J9d6(Y.#.aR[(+@]89(A&RIZG-(aWgg+@
[=5#_V2EM:5g/3M#UUCJ7;QYcN+5OV#BF=g]0[f-dYUZ[EdU#M82HCXI.LO\N1,Q
.9@d9?ZOEe[\g:)GII(HC=U1515eOc=Q#/0A=7gQV[UYYK[\T_a)b&D^.YO0M@Fd
4Ja4;YK=SZ=/=DWQeRO(EN8c<3_/)H_G4;]\A9KO-[<^f051eYTbL4LA,/cGF:,E
ZHG,V+c)C/T=:<g.\.a?MY]=YC@eTO^\/;/Q.)#.Ug5J8;0>@KS(#5@QP[-Bc\UF
A.8RcUF4(X3)GDY&fNeO]/X[O<<P>@;/JPESPT-AA]c0E1a6@;U[UK,^GCARNROc
NS8?JS)6BHRDg0JdJA]/J/dJ4DOHM48#(7aW+S4YVET<=K,=B^2T:F4Id/F.B6H2
4&HH-C:c:=5H(O.=Zf4(+G+H59(#:AOZWR2BDA_)4C\<I7b1FLF&c82JK7^L565K
\Z1M-/<Q@#YDM1K\U@][:9,P:JGdG;@(B+4UM_G>R,C1F3Ac&-)[TFcM<]g=0<=M
U9UK^b_A(XAG3dB^QVN@7[d7F63SeXYZG[Z)XLF[FYd(;;XW]1]4P15Q[(@>Za^A
@3#+_=_a-L+#FGcU#?2cf0#@1Y9D5+Cdd&@.AL61#Z\W?aFgF(:DX0+)1,Se=A7S
:]^DHKQ)C]6UAET.f]D76/PcF4S0Ze0Q,_C^WY]6BQ&:>MP?)<7;Z+F2BH;IM)d&
P/?W/HSA>4c,^^1F0Y4EdTD(<&G7D]NHaK-HO+X1CZL@-?JO\NAaCQ1(N/]H3eUb
HL3=b-.-fE:Z&#DV4TW;a2e_YK7Oc3#_S29U<\.;NbCCBK+\+eMVPL2b/fdN2Cd:
Z9NYB_@8^BNTQW-@d3@2YB23GJN9B)WK64]F=\4-@00_bLYKe08UTTM@YCdcEfT-
7BC0d[,X#6gbZ6W?H+cI?JFdJ4gS>U0(8L-A#UbKR9^T_J[\;SWQK/]LSV#;3#2,
_DIQ4;GKTfKa&<BTL2MO<@\ObI3c9:W;<f&QJ?94\A^(,e^Db>TAFU&[(<ZZ(GCH
=<?/#1SX1Xa;-TS2Y;W]QVA^@X1F7=^_ebU)>1]W4Dg+FCRB?&GJ4M<1S#::>JV\
:FVfIT>J#AIaM)15K_^3I3He=9_gK>WYcHAffN_XZ[,\FEX:N<6(>[;7(=e)>DcM
A?^R..f&AT^ER=16gVB0QfOO2JR<Ffc=?eHBfKZ\#,HUY]e78^^Q1bZB^fKP;g]9
DgJY.8KBS<I0CQ3;S>/N,2>.I(^b7Pc^e:K\+We@P+R+=dU9C4&\-EO?@Vf5b7D^
I1A3B/:NNeHH2B9))U:NK&LFIYM]^V)<;.=aK.SZXV<UHX+BeJYNc_4=g3Qd&)#P
6@D6]N<2b\7Kf_?B##5HX(KcfMR?ZCSCdc5VZZ1@UDME4+=Z/fEX/>>OFg\23D?1
+GM5(I=EED&b>6K@BJU14A+/CB\fW;5G1N6RT&N3>aG0B?c^1(9E4F]5XM2T?<+R
-?[VCMa[AgaXUBHC<L59SX7:;;96GYb(&C0=JV#dX^+c[dT3dEf008Z[W3O?P77c
VQEA=1cO<+_+U^_/a-P^R&9.?T2U2->2N81)KYS?W0c/\QZX(6YgEI\[,WK6f,g9
?>N[I&9V#N2@Qa>R9Z:5VF0FD0HKX4/OB](\5BV43.EB\-A3(+D<T&g9R0Y0b1a;
#&PZ/GQbD90Jc0#]d:Ge2f770HA#CBPZQ/Q_dZ,>F+WA4a6RO/.<>C1DX4VT67@F
\:.d]@6;&@[1MX?+VL-EWdC].AJE;Uc.CJ8FQdE5]5E4DZB8B,)-HS<#X;TZ6H_9
Q;Q,==WN)QaM9d-HZU2OdE5>RIKZA91TW/LNP?0BeGX[W0NR)6J2bBDE7LNX[?FP
.4CXOSDGL)-4RVbfVZ5UER52HX5^EaAA@\9TDX1^c;;BO;OSK]FVN7K=QN/)dKI;
QVPG996HARK(W.e(3e662;P6cV7VZ5)RWHBV&0deR_1GB@gRG@KJ9>YRWT#1-Z91
_HLa6[G.=EWIVANe?ccR/:-WVC6;eP0>@QAe2+WG]CM6=PEM6GR/_-OIF8>B91B=
a0AH&H@MaU\e2[SY?0-THP;799,1#0<72MSIDFa4CBWd9&14TI:b)?Z>QeB)gD;^
6L)4)MfX#9)L]9N]fOE@e]5P07Y&-7aD3b6ZUVcf:]1Z6eYKGXdVT)YM-^90U@Se
fM;3R5.TZ9b470e<?Q<\K=+J7IfDP1203H@-:N)>&U)I<Y#c+UfD;gA877LP)4g#
KUD]7(b6_\FdQV^=?0+/bLf/e@NeE0#\APBN_V5X:U8e&;741+/6<gYcQf[YL+?R
X[Vf+M8O#N\)GRVNVZM(,/bUbW;EF^#34edE1acHCOU(8>RLaWFQ@ZbYQ=(BMaF1
-LUXV^X7YCM09+^KDJ54S03GGI8Ka70BRINK5gUPI--#ZHMC<0[\#H@@Q/\SMG_A
Zd3KR099e=M:6X@+:9bcf=d&I::H41BJD[6/a=Wb2JbSI/@-3?G-W452a>:9]RV&
7[9Jd7B8+_e3&ZVZ:#3eJ.O(bL#X1:;[T,25TMA:+1NQ,,)>f9gCH=EG8+H4/JK2
K?[L>K&eZ#CK]LQG\M+32AW[M[b3MHa9F0+QBc>BG&d>9JF(GMfTT7CJ17XJeMCV
fG4E233(a<JdP9B#+Te1MefGKQKdX>@d))#ZTGa<RXVAW5U6bNF0F,LC?W2JNId&
QAAHN13S).c_JY0[:#:e]Y+U[B2aLb)H<5KcNAV.]WT@D/ZF2VTT(G9LRUQW;Tee
)]C@1;(-S[]=&;dJMPTGg<10T96BG9QWc^6c(6UZaVA/Z_\(M^f3+VQNL,O<5XKS
gA?&E[]:0D5W22+:3@Q8-[[bYfg4A>dRLf(-]Sf&Eb5VgX/159XR@W=9EGdG&R6-
U??Be4ER/8eFU<#bCfQ&L9C-HT\NFF/:#9C:G-RBJfRE[RcVO-A^_gE0<)T@H.#;
[=bX0VDd,f[cJ=\+HD]+P8gKRHBGD0Bf:HgECKOecJ(58CU8U#80KQT4+OLH.[79
O(LU:[T\TC<MH4@=B5([V)&D^>:LbULNA>b=gZ;LOK[/B\0f4:8Ifa+eGdg\/88>
8/&3>g)d^K>>]4_\a-L],cPU(P&.8\#@d(K&==&X)IeYO85bMZ[[fD/N>aIZV2X0
-MP,D>=KT1]Dbb0Z;G_T&7-=<eP1c+Q/A\gY@:)>b8_)Ha55BIK6ICD@98LYR)Z=
^&RdW=N\/.):CY;2Xg[Dc+Z@Y:Hb+7ON4M?W0<4AcbA+X4D4SO81H66b27Qg8>;1
a6Ge<S419[H\<-\W^K:B[O0fT^b_dYN.+N?2>6S4Nc4/8O&UX:48;:YP0Q2NQ]H[
O1IVd3647H>g^&+E]GIU1_6:=UCB&-E6T.B4TdPDcE9aWB<>D1^,[]R6R5ZC/)@6
D0:OgTgYY],>K_dH]ee2K8P(dAS#A8,X2Nf&;.9F9eH]O=><F7YVC@5S=?J/bQ1f
8SZWTJOTEf\Oc3g.UF\]FDDS#^Ke-6g\cL2;54+1_2T?=\/H)KKDHV3?9-a&F>D4
&<#?O4HMIEO(9U12]&)^VSSX+.cC38#gZZUO&3+R]4>A4f8]ed1/AAF@L9XP-+CB
83_9ACFW3&@X/NZ)(OKJAY>X_e6.0NUAK]:Z/bT[V.0-+Zb]LH9>Xf\URP(,Pb3a
;3?6S:ec?(gR=7aYDb@f/-MZKZ3Uda#/R@:[X+\NQ/+Jg=I4\XV_6,5#OCU\&()6
5^_^Of0>agRG2F1b2-BHZ^U(\(^-D6LA_2TQ48cfXI9@+c6be3RP+0GHC7Dg5A96
)gd\7AL)&BD4ZGF7fQB#[SAQ8?8<U(G>P,\,5ERV:6bNL7L@YR:b3;1<dM#YXH-&
/,WYUcY19B<VT2JQUGL3babN7DdAQ\AMIU955ScBB8]<4GIAeP,gN=>FR\bU3@E;
T,HO#6<JK\)G#ee2aYT[(N9<.>6TDVHe>@>+8[ZVcGRFF7^.>C&8>8IQGN3C<>,a
^Z4.0eH;IBU8HQ;T;RS19d^Y6\cBU/VWa?8ZAI;C>E1(@H&WVLHDXTf44-@Cd?T3
SQaF)-CCK?/.7)A.U:(]U7Ua\R9W.)=4S.^<PCQSMYRSQYD0@5R&-O<MGIK>-@aC
g@@VP\5E-eN:K1D^>7QALfZgN@_U^1=]U\UV)[GJ52W9;=5ROE08@9/DZ0,TaZJJ
W--F>Q=&=.4<L@E9QdLQU;[daa:G0/HT,,#eR3X3L-3GJ#O<#J+NXFa14Za)_.X0
Yc>GB[@dYFWO9M+)H>VT^V-6MNK)=DfPMGI0^JM\M(J/=?g+]0RISHebZ76YNN88
G>;(&V6c<1I&2,UOTU+KOWgNMG,MH<O/@U;3R<V-b>(5d?#)fCOSP=VXg,W0FC.7
A.4[;NQKSN)>g5bEH4[Xf=@V6CgD8T_eKH9ZFc^)Q_=WgKPVTG4)3XQWd8Tg+cP2
@cF7V=/]=)O+V^2C9SKdT]e>2>Cd;f&+UQeGJPZ:YA1bDLMGMD7FD,8WNB/Bf:(4
b-EI2G]>b-<=C];ZN0YM[W0ZL[&73)EfFfX>D^9g?Z(E6K?G)KGU&VLQ<;I0P(H9
KgYY7J<W2W.R4aD>ZJYC2d_,;=?#8YS60HJH1<V/\Y9MNE1\L=>]LXBN^@E4P>#)
,_S^TBI2[KaABPF+^6[;_PNQ&2#9IOLc(-OJ[6U9be\PVHRC1c-Ub1:V66:b+:QP
_[?K.<1E:IeYI5>-X<<LT[::-5O44)63QFgIL0AA_&,GFBNaWN7##U6[I>M6&Ab,
77M8X.J?5_OZe7V4fX>&b_Xe8+YEc.YL[C0;V:(6DWVB&GSDE[O?c.c9<[NW].,D
Y=D[381Q]=?)DZ;aD>]gPXV#UR-=DY<GND>KFK20UIY)4FP0GC3./b@S</Y_d/M,
2+/f<T&2RH5b80MPb<698CP7+bSP12BPV)3@E@Y+\RfP1967-;3d&J_cT1MeU?&F
PJT,?@FGRY\Y=[:ZX.G3F3N38/2IfIM.5^ScIc#0\AMGMG5eK>fOJ^aPYND;M=b>
e/4NfU)ef,E+@6N4S9.dH+L:25=X4e#CO]_4\(V3L0=bI<8RD[fM+A=-M^YJPZ+\
<_gb_1,5]0&EB:fgcPW[WJCMf>NfC]0Ocb6I+VM#]3K.&,b.dJZIZ^:(32:B,)b\
_aU,(:7;(KV<gcW.Jf_Z9bGKJM=4E(T]dXAKRd/CR^?\C(ceU+^RD(:)4TJR8,UC
=M<7D;f9TN+(@9@B?VcgZOH;P2@cdfVKRg0?C^F=I#+;Q[R&3QFWM;4KMgE1C?2(
,c_M1+8;:R(S;(X.^ZQ;Q/a8N;@)U^FRd;JBbSILW#cVH3?FAVa=Oc+aA]3ggOdd
WVL5R42SI)d;5QWc:Cf@&;_CQeI82BCY7/5c\6CdNPAcd>43;=HBd(M=>,[^&7Zc
/1[X:DN0e[=E^<-RZ;a[Ng37#Z;A2:S3<VSC(UV2M?FcTHH-]0Y1cWCIP-6X6#4P
_8#33.1@X^E_8J]JT=?R+:+EI3M,LGAYI+eTO+N9N\-83^+(N30eN6Qg^[bN]W(D
\:BV/-e23=HH(6.:C7+gE1YWQ3Y8M0N#]URbD@]dNK9b&4PI/13):CL@JIDAbXfL
R^51?f?E\I]O&23^;DeM;9BB.ABMI3C:E1QCIZYY@MX_96_3g(Z&[70\9RN9GQ6L
2>[J3,==D[IM]+eeB:[bXcA96H8-V2Z#<E+^9H,(=LI8e0XYTTFVfA7^KGF0\U&J
-H32SIE(X>c/O29F1;8Y0Z,4=Z]#U@JD0bQ>I8A?Y7f0/PZ8O5+/&g7<Q>dRE^Da
GX96R_/IHK5ScK@XQPU(aY4@EN5CF8[JV1Q3G@[G50+1^#&KF/5YDU);OLZa,d,L
GbGLA+K7/7FGCE(5-C5=4cO98JKfZ7HRe:^1WeO=Y_I).C15.E#K4c@W;[<e]Q:N
+LJ/0#gOUf@5H]J7aUE#<?)aaII5CF.,-MR.=>D\bBd]&;WEM48;X&RCQd.SICG[
d3Mc:Z)<-,+IT@/X;R7-V[D_P>U@Q,Aa:[c\@U?CUSK-^;K9MR#G4=/O,<=>T[_[
]K2]7E)d=5W&^.\G,[a[J&:>-B;MdRK:c.MFM,Tf48S(8[,HH:0Ra=I+QJI9@TZW
&)420+_P,_HXO6;.Yg<]^6?D^b>Cb(;[>B\L<DP3(3CDdMg_^#6d@G\&eL66IXa/
^1V<Ig(ZY(,YO?X7-0;V2TJF@.L:.J)L,P^K2>8_NY@E67^XIF#,25^V,)VKE^KO
J3/]<]K=XaNK/>Q0_^U1AIGRPdAYV^@RPTW1K(1\[AW3O.A7BHda])1,G[DDBX^;
I,Z^4@6P)(8<5[WQFgb>55C?KBNM<9E7(.CL:U<W+&M4bdcD+67+(@eX.#=UWX:]
D5>/9H8WYJLF=,2>ML0[GIe7d+c?Dga7&3-\a)KI@=_gKGaG6B;G@3UZY&R2E8?4
WbM<D:@T0OLe74e^Z+N,QQ>?OOcMS3A\:?^fg-XOJQD-SIc+c,[)8CL13#^L=M/^
LaO0JU<Yg5fP]cY@&MSFHT&M<8P(,+T(Ob.EGWQbYKCIM<VI/VQXS/WYUFBD+e7T
H6=._^UE4/J<MR]#_3Z><E]7/(d\cR>0ZV1<XOUFd:-N3TTBM:N4(0W[b^GX^7A.
Q&YVN09=E/F.6D4-IJ0<e<[OT93P+>Z0-0O3aGg(fMJbWQ)(_CZ?O.D;11cQ>?@8
/1-YUf==&J4B8Q8P.>G2:>-JWFDg[YN6S)>;W_Ya_VAcNGbaC]>e,FFEA-RUaN7W
KeARTFR8cB#QE0>Pc/(3UHPH=&/35Ug<A6P(#K\]^f>.TMTM^3INF6gY<2KX/>/.
bA4H,EJb_;I64WJ2?fW:@agYJT9d;=W[_D4FA5bX2CCX^[@G/:KQdSaJ4@a6e5Y,
d(g<_O^I?HeFBcP@EgHXOQG1-XRKY,1NH\RX3a+AVZ-N]ULXU6ZM7YUbg>A?6eM,
Pe\WF+YdYKWMdH[aXM7S55eL3WJ/[/9>M0A-A[HZK&)ZMLB5=74-9,f=UJ.cT(3<
H:)<)bdO2>DV+,J_6=H\)BJ\89NSQ;4XeW<c[+EU,GJ]12#fLGA)ccV@@6FLIO</
)2J6+FZ:,L]E3bfF>#UIS]JD<H&#W07R1J&^1WCK?IH>F0PO50_5&ZXf4Xc/^L0-
fB#F[^a]AXNb]b,XX;5dHL=+TZd#,.\U>+([/O;QLYe5@K?YF0F52KeaM(\098[4
OCMWG+DEH5fC:d6RY,CI5OT6,;aYMLD^Jc^V:H<HgPQM,#[:U]H:O6HT]0FcV#C/
&caR+TI^I)2R^<#/0U_;/Y?S9Y.g;1Id=FARI3-3&NY/QfZ>cPX3>+4ZS&O=55e^
GdX=eZ5)?K&I[9f[D()E1RPS9CfBQT00F=_.^IF6M>DV5F=HJfFVB4GG>L\7+6XB
]ZN()H5[ASG\[>NEQ-T@4gM;Qa(BFdZ_[J9G7#QA1R39a[YFXO?UKK6L1&.;585H
Z6Z+4.G3-PCXAMVFXSb[bZdbM+0>L\c1,-LeD_F:>BM,@-E=>B\DMCPDVK5GWHLY
-O#5UA\daJ0f6O<,R(4AB:NYef]];WX_/]+=03aO]bKR/H_X7FJ9M[BQOMKC4?8S
H-D;SS^>]LR?\gXY^6TUIFRfN?I_Z>)=_^6OJg+eaSA:WXg_TP&)WD.U)=8d[Q=Q
]A)4cNKIbP11_^O6[(]JAb,;g<;7^9K5:?9Y@48MaD37B-K57^bPB91:G-E7VDb<
?V\^)X8=1eM,Ica]>cf9XH=a6IX.<L9SdfJ]N3Q7gT&D9#&S7(4P\B6=??&#+c[Y
GdG-.^5^]JGH#]<=>/JAGQ@Z#?XF<f09XF<bSL)#GF8Ha#PWF+.XN6/8=Fde6c=E
2]]7&Z:5NHO6be<XI>Wf,J];]F&#X0\_JJ\E6\f7M2/[7(PEY)CB:?<D?/,CR2=a
B5FZ+L0R^2B+]81]CZ\AT>#6T@Y9NMTDS_gW\WXN=.>?UXCPL=K7Ucg:EIZJ:EL(
9TC;<]:RWU[d2A:#6g_IGT@U]aWAJDc8^,NT]H6XQ1?_R1e/ff^;GD-&(<WK1ME)
>O1FWg_.F?3(=[>c5GM9K#eSDIX5,=I<H-(a,?=4D@TI+gCTJ2g02/fW9MGQQIa&
5CE?2.X1BOD^X/:A.)<?6ff.O]Mfe_YbWfB.V#1SR5?H@WV62<P;+&\TQ\5B4[g@
KUCb1DR,_>Y_#d;XQ(.51aP,<JD.#VNR]9C-U-AUPN[-L]0-DF2FeU&OV?S(G<:R
:@]3.:UOQTO;)ddVWcBa8B3c/WMJR?Vc(<\@(?CA?5Wg/=N>8U8XP<GZ<^[4G2#g
N\.R[H)?LP7.84cbO-TCE2;:>PX#fJ@X^@77B(;d&GSYBUTO&f92@.61UfJ]^gI#
fJVQYSeSfL0Fd3c9UW2H7ca_c-fd(&cF8fTRLJ/NI=?^76^:f>;3gECa/.8LNR?Z
BI?XOO9YHGPAc03_[-a]PX;?1=PXLaBQ-G6)0OF63-^RX21fTVXZO[bN9=eKY39J
/2V4L,#5EOUQD+[d/YTfg,(3,V8-89JPCV5Pba:KbH6EQga#YBXW23V]9@V^;]8&
_+;FWO99\PV[&(#H@,G7MRT\=fU;bK_B31dFSR2YIA3YWX#J3RPeUF5+N2B_@Ub3
,JZf]c_9O<cfTW;7BX2HS<PH9BZ\N,Q,\;c]5RVULHN,SI_W]2KI\E:.7[\)L83c
I?12Zd[0:Z=#T<K0GL1()NWJRKP,a)K]#X(>U\4G[;Z^@1].P\36176;D<]gcbI8
Y#:9MW=YJ@d.-T8@EENNKcag,9#(39f+TPPd@&Cec?F-CRR???&9)d[;O,BZ;(VI
BLe>9/P2)aKZB=9RfX.:DC\P1.&I<2EC+4RI8\M^]cf;X-cO.f<3Q9b(3B64;aee
VR;/D6W#3QN>QL)+aZY[:a/f<_.?O3fDYDE+Wc:1ZTR_g&\cddW>B8=+aYC8W<8g
0gbHGg#c?M6ZAN:@T]<YWGMPJIHIYgcK:(UDg=Z_2L_aN2&LZ14(@S785A/F/f_g
(,]TF3U=b#Qb2CPUS9dP6aIf9UU@7GYY3/Wg6d922+=YAJT./A\I=[Ta#HCaWM=G
2^(2Nb[L1c-M\/G4+3cB\.3-2S>)+6IE1A-WGAgR@4:-H3RG2YW4g(?;._SJQ[T+
9<_^\-bV[;,R3XKXgaBJM2++/g\,F\a(G?P&;@W/RX?5;-R-a3CG;)3T(=4RBC4\
7S0FB]H\9Z07@KX@)ce#GNZ1/4(DHAKO1U3eNO7\&/Sf:d3GDW/\N(c6/WM3QgeP
L)BA4d(\.7d_eYc2TCK\_ANZL_5PPc_H\:8eGOOVI[]W3J^LST8YX.Z@)(K,a1Z@
J/acCN1gSU3KXT8_Y4.8FC3B6W5fXXb8DHMa&4bc?69[@X9=ASd::\B105WL9C57
Y2(B[)QSB4):gBCX8RS1-dZ0C9_PYKM]-g;JeEB91U,30U:f9OIX1+POIHU\G8dS
_>VeXZ5JDK(#_e_/N)aX^8:8UHLW.8-5[POK,ba)]U&]gf@AZ1USedaPe#F8WFR/
1a.WS,RW>U@e1UGd-6OGAf&8D5\V;bGd,BFeG\>=fM4CX,XUV3:><]8EAFa?AVH#
VUa:FDJCee,T1RFc-]d-U_11bEaD7CK#6IHR?cFUHLJ4E[_&4V>VDR\[EL@^VT?&
eOQXW>Z.S-D;W,a?>^_+^HFbgY\..T40Q=M4P?I(L:RbG]e7ONH1#Vf)ff)Q;VXB
a=,Md:?KXHHQUaB<\bPfZ+DT]V/L^(eA?/>4H@,MHf=8_9^@+E^2,\>F5E@IJX=@
@:JY5)R85[X+9DIXMM6JF@8(<NJTKGF=A(#7/F>86E2cF>W]76R?V^WBE31&a&a4
5&a@XU;FAK+2-dRLO:H0&g@N^#c@eI>B((Kf4[N0]&5+5+ead>FFb5BW;(Y\3.,1
P+c-M7HWR7VG^B>gJX7OAV_(I6<?YU;;]+4.c1+FKQB66SA\0C,?PfBC+H1)QJfU
^_g)WQE^CP^C3CfZDJDbPb>CSXLe;X=&]7e8[QGZK/TB86ZYGGF3g/#D<N,(9:\]
Ye?ZW864\]?E)#b/e8IB9d&/&YE46g=:1NZbB7.8,W5<ZO--&C>3R@JUA=RJbZ9M
Wg,PCX,.E#H#@?g1[&+^=X^)Raf1=:@AOWIgS.d,:1B4MDfKA6?5]PBc-;97^bEC
;6S:EG\35)aG>_UC@IP/>W&.SM(VYB(>?4^HS[Pg+@O8E8.[&b#[\&eL>II&OGg2
cRKGXP+)[#.M3C,K@8ZNLQV>J3-3TW)0bDZV2<a:?HS.NM&:6_;B/:&eY-_.)-cN
KYAG\;=?K<)<bTfHN3N\HC(^E,gdJb#=(A8DL3QEK(/HT&ad<\77LJ^f7MATSLM#
_(NK<ZA0c2MAN.B86e/4RS>BJ@T_,a7J-;[16Ue2D#KcRSVdRO?R?I5+KZM]9/O+
M0Y1dAPPT72;.1ZZd_CD(gY^=6_NO[Sga.2,JTK\0IH-I15&,6_-_V;Re[d/:&R=
H9BRJ-g\d?@fDXGHb:9^,@/Xc+YWC_;_f-c:()>8Y/_+0Q;Y#FN7DH/,N3]2bNYD
f_B:dZ3FP?=<;ZQd,UWcQSJDEWbaG0MCZL<\13:Ib4^g39?Ra+S5UFeL+4:8DM=J
JY6FUYOD2E#f8_Q;C[7&^Y>H=)a]X[?9_TB3eHD;N]&7RIZdNfge0SDG/-(58[Oc
=AVDcf2HgOUeU&N8e.#/NU(VNHJf4e<ST8a^7#^[N)O+I40VFHL_N-9bAT>((=8<
HN7g>;cL8I2#bgP^G0#PW?S@I(5b0<S;^M1>Z99fYP[WFW5VS^Tb;VC-]1L>T(0?
(P7?#_Q2U):\;WEF7JO+.JPbe/YYf4E<8Ze9BA>Z3b()G=\c<X^US]&aP)4US4bE
RT5\1F]K132AZ^cJZ,#Z(0[IO]/)BUa&Y^H?<b_\TgM_Sa(AgO=^:U_==&A<>(c^
2.WBUCeLQKN:2LS;.W[bD/L;N:EANZ;11WdJ7(U8K\.;FO=]Qg-UPdKZIA_I?Q=)
AdX\SMAS(_)YU(0..)W>M_EaF((T]dD+_BTD.9ZgD(TE:K?AF-CB-L48IIa9OE4H
NOeQFQN)0UM/DN#a7g>;+&]M54ebb9SbBafD2d&#LM=-<YL6@22@g9VGgL3eF)>0
U0D:K507;0aFYD6L8b#=2N(+e:7)1WS25BKgI>>7A,9#W(LeS#X<AQdNG/]:19EO
X[cVRT(;SS(UA;MGYV\O2/F@;f9QJefeX94OgS34_IYLG;->7_6I,a;/NNWHXe=c
FSZVZCRLeO_EHN^O4BYS@Q(QX1W#C]+QJgH@(7<F3D\&:IdMUP1e>Sda<cQM2\0?
,#<O8H-Q>?dXKM;_,/YaN/#H.TFD,A>2?;R+E<5.a@Sa8RY3,OTTSIF_[V_O7Of.
CPN1IFUEE:T:9_3Vf,D:Sb\<Of4<::J.22M3_ZaPFcMO=L9Ue7-/V<bd+VdR:=.U
]=MN.R&1_Tg]H/L62-@gg#_,P5C-^#b)QUES-BY0cEf]^;)fS(,9OUX&><Na<\GU
d=@^4,eP4_=;]/KKb=0GKX;G)12#6V,C-4eEf1Q:#U=]ZeTPG:-YJW(ZUCOMV6/W
K40/O:)eR&Y844TO?dDb#/cKbe?6WX^(1[M8Zg+e6S,.G?99].U,IJKegI1_Ve)Q
\-M,P5a_C^g/d&0]0V#OEA5D&/:E.0[BE.;3VC+XJ]/bQ/NFN5+@#D.-A^ZDO]E_
K0C_=aeN89T8K1TeMS\50S#[S6BRQTZ6X=@64__4d,?.P4D(-73MNVObZN0O.M:T
&B:Y4/76Y(2W(U>^WZEBLS^8C>-/5W^-N(+59;^/V/7^1fLC]VZO:C4T0P#:O\1[
X(aLZ;,BGZ/b/+XQDS(2JJUEF]C2IZ5bV6?T1/:fO,@)>I5B\cH3?</9VVNd;aKL
eP@>,4URH[Q1DA(WcPK>MIG=#869UR0:8;^<XO=\0W>8_2VXSQ<K>H_T#&B7][ZR
<,PX8;DbBfKQWX7D6C+aBHQ28XTEK:;3\XG@AG06@1,FZGGN2_8R=-<Be.QTQ[=J
.P2,b&0RD5X@M#e[LZ9HF:597:=:,94]3IJJ)f2N.82GF[]=ZSBT9(^;.VDF,L#&
f2CE#gJ-S5+V@,0L@Q]UJ6-K3WH^MV?V]P21L#[:Q(Q:3d14AcMGI8D22D:\XaPa
B?[B]H(ONB,(9gU1->XOCFZ4]@9L-fDDfM4[1eOY6LZ);N:XWf#?gEHNV29&:FP9
#^&N17ag6T[#S+^R<b8IDaKCEZ>3D6cS,X_^YS55Y_W/7^@9_A6U<BZ4X?3-5O0H
]&GgM?d2c35-&Q3SHVWC_)8NB4,U9HgVNd3(0:X\E7?@&C7ZWg?VS=1H[b5b38\G
88>5_XSYJXLPXef&0[7C5QcBIS>Y^7M:\FaJPHd#)];;/XKS_aI\_R7fDREB4aXf
1NM;GYHAg9aM1CQHe7<^1RT.O\TK30_&&L[BN>AIg)[X@feY04g?C8@(3?IXa@1J
;+M6]BC_(_>C@MF652BP:P1fcB\)2/C>QXTT@Y:bOXQ4=VOaC,H+>I.>02@d?:Z=
W[H)?YPKI-gb4@I.N=E29IBT54</WP>;FX<TI(W]@JFU/,&e\L7GRJO]B0dEL-Zd
KcZY-a6CSUg1R8dBI6-6Ibc2JBM1/Q@)=acOYG-=2)@-KFgEYa3DWJ8&U1&L-=NV
,[=^KfSc[U02XK5^R_:Xe0Y<M:RWdPZf5\6:XeaU)N<+D1G,2-V:O#1GJ3LJ?^(9
V[EEfI>c?f\G4aK;4;#KFGZP9I-\#8CgEMMYIC,U/:)6E@<b/JE4VS6H]/X)>B+#
N]?Vf]_f<bF3YUPE8:U-Z8c[GfE8Q/IYBN_f5Mg@:T+>X/a)5_9J?(RRT:<ULY@7
)PWRfd+6(ZC4R4dHDYN+0/-?YbEdf<dSE1(:_c^B<Pg=W7X-?N[94/_CN,_K_.>c
c6ePg?gUU7].(XVK2>MWOYe.TJ^F\QLDU9_b#RAQd.9Na:bf1K\<3)1^^c-e:/c.
W8&C3]_@c^-G@N)g\HFN-,YNWfPN[N8e5C;B8;:DY3Z\<eS@HIeaP9@<J.egVg8+
aDS0IK,]0cB.WKZS+#ff\>2]<AgM(.\a4ODB@7NTbP-WV-UN0.\e-O3?e[>@1WZ4
@T6bLS2D5VBPW:[D@=3.cb;:e?2d6KARa5GP<]_ES;?A,/,#A>MK#54#0JaDO2^7
1NYEPQ6V817G#KfXTQ9(fJOWdW<W5MD?2:S(A:\FV+bQIdTcZ0E6>.CWBQb7^94J
Qec^MN=PVDV&K+F?_]Z6+c@YER_Y<\gR>ZR+#M+U+gZ6GNWF\a:^^626MUL[_]08
)\)2UYe=?cWT(>JBY;9aR)H(]L9O?;g:)4GaC:gQE9RTKa.Ld3^6)4FO=TgLbUg7
:30RKZ::?#U+5Ka(75QQWK_OcY_;B_8N;1DR_O&FFbP6UV6a\EL0fS:5Y>)/&SU(
U^]G<:WadECEZ)9GJ4W;C(Z0L6MeC/2CW4+1>AXN9&>#ZCVQ<18:_4IMMQ8-+(=0
Z,RG>RY04F>JJ,6H9[<Q(7B8-J:I4(OU,IQd[,PF<3GeWYTcdSg3<O,4d8=4=Xc9
=Z;&+,4?VQMZJ_[X5FMVeAU/U,U[[Ba2G.S;g/L@BM/SFYZ>4[fZKC_6;23O1F(L
E6<IY0cARU3]NQFXRVg=3_0LE[\>&L,3Hfc)Z&4U3;0d(CJ[W1](E+Db#=SI(NV4
;7[59_B5<7QSF]1aO9NM6[W4Heg02,f?E3#C7WHYdUWaK49Ja-#K+Ja@(0d^43W1
Mb(FSC2K1[E3.(V#7<1(=/:Ja8eE=da39?@1OF1D>LD-6P,UZGff.]WHU0#be4S-
9VT4K[5GM5dRMLbeF?f;06&SORH8Rb:9\8b=f<DcXM4d[[VJ6/9[4]T2eYd1W4ZF
EY263e[8(?6F.]4_50B,R3d..IgbC5BY3Af&)?O?=gS[PC0I#c(Gc-P<I7VQb@ee
Zf4EWbX00fT9&II&b?EGaM?Oa[Df8cEg,C-6G93RJfKI,Q0YOY8KQAbfRG&4b<^Z
>MRNBB=^RJg9_)Hb/H\_,UB#<D=/UY\7\YMGP8(4,I0Y]H]Yf-T2,9Kc_,6EM)43
P^TYR#_10;89VM-LHZ1dK[P-Fa+.Ga+4_Ec)8[K-3JXT@0)cXPaEH3DX-LN(b08N
2+b<e3[aX[9S<@7-GQ+WF)+:6D..I?M):3DE-29Y_a:V[;]G84ag6SY_8-5LEX:H
6ZdGTK:&0)HY<[M[X;]YV&PbJ;0_I+H21BA#^L_0YT14B:+CPRUABd^UV_6C,#<A
d_&>YLE=E)S=YFX;8D1[QN+5MbLLEAGHB7A.(FfE&17e=:N<KY\7U?bc(9f#F?E5
,@Y8#X,5=f02:2B09ID:f26_QJ.3XbJ-g.-FAX]A3Ae<91fW.CL@<#fbZHJ[L9BR
:T8CXSQ:fa1Ug[EXURP:\\@:C9A.:F>C_Fd^eN8F_/c2]F+f0ZOH&]<K@O8T_KID
;+-=)6K3Y0XgC<E_8MVMOUA&HLOI2:9Ie)30&dIA[Qb[Q+,T<>Pge(WS>I32fPM0
aI;cA>Ye\(e^Vf6K9_BR54.E#GJF,29(K)QM[:S]:X0gGGZ&:ZIC^TZ-+2@L<BC]
eBETdS<8ZH,8UC<Tf]BWO1=1Hg=:UTL4_[M>d17:]Z;9McC+2Fd2-3I_)#@VN\RG
ECCf_DY1Ic.U05G;e[e_\.^1CH7_01Y#]Z+O1:8C0YA2.QXB;+YI4-C<PJHO\K88
0?:DAD)4Q[LFE<<S^b<+.;)G]&[\8PC<93WHKA)>^YEM5;4aZ+V2[>8\Fbe><X;6
c=-,^9\;M)MeA#D<EWRH]N##3BW.S)BcIE#1<.W?GNfHUEQc025/WN^#6U&H]E1C
Qg/?U>>MLE&<F-;M0SWS&KE6XaQ4g+KJa=_;--,<J5HWg_3Z@D\2JRd5EH2MFS=G
:-7fM1Z[Ofc.-FL1,E5KGFH#B)/VJYf_[6QV)OJZ4S71-2XT]C&)=1<UH&8U/)GS
@_E08LS&(\&;:BS;A136.2^#OVQ>e(UUY9T52d6e(X[ceJ;1Oc(S#5_I\(G_<#L3
QA?=W3M\U#@#ZKG2:2B#H#=P2>+#E2[Ae(Y2fFY,)<AOC]YaR4I[1eQ/M_FBV?DO
FF>=>TH3ET0Ad<\6KL4=d\LABB?Va<#P:7CJ16L),:QOfda^D&g;DJL:V+;]E+b@
;-B5a[,X@8AG)VP#XV#eS:I40R5U[1R3YTb\0,&V:M]Q^C7T5@Vg5Re40OUe9J8<
@D?+gKVQ5d><>A?95M((]bdPFgABdWA<N0CJaS?;(D.f7Wb5:]RI<Q+K<-]5M&/P
W5fLES&Q-^X:^AHC()2WXAX3(@1;99MMC:Q#M#+f8_P-gHS4eb^_HgTREedT3[Gb
QCa6FDA2VVaB=X=gW9VcN=B5C-I4Vge5[b2FEZ]Q[;81OOT8X174?]JJ<D::7eL1
^G(U.Ee=/3>4N1\g9H3/S3gK=2PXJ\NVS?XPWH_TVZ#_N<Z+E\.KW;81/-K3]XfC
UTcIO_E?&&Wf]d&BLN5^)GfY3I<A5Q-HS+&>7)SB1O03DcV9&E)96V,:/0QPEZSR
(WGO,c05N=A=\WQeP=XN\@.D;bQ8Y5.QBU?01@,1Fa\\KAB3(@4cH9AV4J@#a^7G
.75J0H2OAT[DVdL.9OR6--1#ZQ_OM>GT&>W[(KRO=<O/@+PT6HG0U;3Na^RF^+-@
OM=e9WB/_M[:N/O(9-P<g6S:0cd9RfR))@0Q<b^O=Wf2\C#J^?;P7ZAB9&^Vc@1\
NW;O0GS[T+@UV8@]DZ=S/(TL6b\0H@>R,]:P3/C]I=c_O&>\JRO540Y)9UBDO;g2
CO&#\HZ6NZ&8+3bfA0@<\\W;-G&UX)3-I<Z-O1c]QW9[O+L&)6MF4]:9?DWC=.J^
f[d7P6<O\3\#XO:OEM)ZC37a(?J0a=IRRcLd6c6ZRH(B9]1?/4SYJ264NRKOYL[\
@N\&ZcaGL0KR;.0gac=2P_UKfDe3^V<-8K](_@6A+eS.CgAX48<4&;6c332UP0Q4
.bMW>[/S<X[48+\?eZHA7RGcWa?,;N(4eR&6:BLO13,=OMbWNRa7[N=IJUa0H<Qg
>]>f;#^&TW:8EG+XM#aRe1-R#10F9SK3eTUf/V]<,.GE1Pd^R6Nb7g)&CV3fY)^O
]126BfO([DDG3,7//N;VdgGK:R)G[H/ME+ZI5UC7E9d:Ta?LJ-<D1UAFf(G(gPYg
0/.+&18F=K\O_2B_FGYJOg[B\\(X3C8WJV?+5IZ<0].#5A.[+LbE0Y]I@0.M0>BH
1dEbf-ER3^L:DS0U.6+CH_PWF;gAF>=\=[#&J/_H9X+3g4=3FZ3d:8Ea?\gHRgd:
L9Q2S.ATS#571=B[#X.2)[5.c[^f</NWI1b>EDTZ)ON07B_Cb\Q;=7W,Vdc/1]U<
d>7IRSXZNW:XV[b^A1JBUV#J+_:P1>[Y(<9#N4FMGZWG[Z1>M?N6aP/Be3B2dP3M
/>)+<F,O.9cJ5[UccO/#P:+L(M_dC&g86]bS:P>U+-a1U,&R#=JH#9g4KHF])5^X
Kb@eOLHP:O-e^,4F14bF::C.8^5-5#I@a0-;,;MVCYegY/#G-NIGB43.M,12UL&g
cfZ_OE,K#ef[73IPXc<#)fK-\)OV#^a/P=5;+#:HZ&:VR__CG<9&1[a+^B@=8e<C
H;=L/DT3:0X)S3bUXb[2cLA&aCa@11OHCXR7FSYb9BFP<2AH0G;YRW?41W/32Df6
U4E;.=];I]68UP-WR\H#=HQQ0X8-0CfIW&(>I/fCR>UaTE-RW^CZ9-[Y>S(P((AP
HD.ILAW?N_+-K<?_);X?3[?,<e3+1PZZ4\ZPFGM?ME[d+ZU:Y:H5E(\fJ]gIfIeH
V3&&;6-<IX(BT6HVf4=/RP(L<CQ8/=9&GE_I67e>0BV><Z40IG_)\DBNAN6O;D+?
[;0YX]&XG.=[DY]\Zad-]fgW@f/VQ+NeCfKSR=3ME.cSH_)SI\<;()J,e@-]=+0(
-@eb?e6c3bT0/NMHHIMM3aI6#Hd7U]3,JKYP>g9K,OWV&XB7O\AM&_D&FR7,U>._
D;F,>8.T<.bd_P,_&>=GF_K.NX_?KSabfKY=WT&]\@0O+AF21e5:gI_<30Eg\QY-
5dNC:V&6R[bCQ5c0_f\V0;a-^1+f;+E\Hg2DQ:&TXLPEB)?3E&:+;<b?)CF,0/]+
.5B.F88=3c#)SNHc3-8_Sc:Ee:N>L,.&9QPb8C8LSK9dId;DVda2G-#Cc#,=W+IN
<f>[[7-LWC:SaQXJ.G;3S^D(V7GVEKLF?)e@8I#3[<0<MG_,eS6GEfcc=T5Me9eK
BgUNWS-;W#&Z+ZQK7X>c3>;/L1R5W48#Ze0K7]WXgJa4T?0fS2P+NV)J)80D7f^_
_\,@5:9/2I&CG:JMA8@:KVCKBE58fG)^J<\Q/CB-)X\>QW7I[^BDDfg^=1EO\)4(
??X1#N,X[+D8@Md14->ZJ,#bb(D/M5cEJ7N=,.GHV5?d1fI(ES=0OY<+VGN?V=_P
@8,:HcK?2I]-G\JV@(7?;\[(]C4XM6BT>W>gJX<JgcB9Zg)gBeH5ebSXfHecCGZf
c>./OK6U_d@F\<>f/(=_Z,WObQ-#Q0Z8<=O;^N56#_Pb7UN-P369QS25=3FXY5^S
C9TY]XfU&5.g)M2aI70+S);MaO,gW&c.^[KRUO:@fZeEUSdbc_Y#Z:K>B#BL3g(c
9/0A)MUD#2VW+/:=OfRLY^R5RW_#DW;Z\@/6FbQUa<^&V&[/G@B?La#BD@&=Ee3M
fG@[O2c[5VgQ9,;A2c7I/BO&7UC-WVEa)BX1a5I>_=#ED)1I.:(+LA?4/YbO,2,6
X9)dAK:.7D8U&D4._Fa>T8-@QTd?,>HYJNR9K:6P6QLeU6,Q9Z-PMXLSd,4+:PR(
O&OcTZXReK:.T8@:a4@Xb7.d]FY36=O/TK.7Y=61ZPZI+W=HA8T(g#<40JL18<?W
C_-HJ2:c8ZZIbJLdP;.Bb1fcK_^:Nc&ZIV:RQHX?cFV>dR9OFRO0^cZbbA90YObd
^#c5GFR53bU7I1:>/ZVRda#VW<KQ.4##7)Fb?O-.S^+6\1F+WE@G;>;G?VN-JX:>
YE7&+O5Gf.2NKZ8BY:^6\HFU+eA_6?a):(K+]:EaC[^=<B[\8dR5O4,8AG]e:#ec
;@Y[A17cFaC)=&g725,[TZA(.Mdf&MZ2MU&g6a>0IWLNWXP=9MRWIS-9d-;_5?<c
PVHCN.a;ZbO7BR#g5=,V4e2(U94P]1S241Y7C;7I\#NU6VgE#L@2>g_C=6/79B&d
67Be\B;VX^A&4NRWI]aAffLNU@aU[/SXgQ705MH1?GM^VFYLAcf+,aZA1=@/gTL^
dH<>=SD)@]0[@(S&4+18PI-06B6N.]5>87Ma74?(OT+db@bgZ);>K:]]I=NE49>.
^YH6S8+d)<Q<.bKO3IO+QRd])W(dL9N.0?WYbB/]<CR,V3#06H,fR(/E&0@C5McQ
beK42e+-Z<_eB;6KGYP\+;XUWT;Y-+D]]X2Wgc=?ZU_8L6e+NXd6d@<&;4cb==-g
cR5&+g\\N+]g#R\eG1d8HZ57HZ=3aQAXafUa4YL-QE67R(YRTNC1TP^ZP,39G?B<
IBFPE6KJEO(^ZIB<I_X+L&g>VP#V1[E57MOE6OO@]@?IONaOSc95:+-D.JIV<;?D
F=LE07+DbO@bR1:X_:6/FHf0(PF8#BUF95_C_bG5B;X6@TfH?B(49CZ:@\\<;AXB
(M6BeWe3Rb/32?NQ@2bQ=B&+K<@OF7]Ga8S8BdPS/]/Z>Xa8U=a[PL.14O>#13=L
=TWSUSWEU(:KRB?cLNBZJe+LMgb\72/_F>\=b-XbD85S(-=,_6AKbb/MdW<PXd&6
W(SVKBd;;;N=80@_<TUS;W6>0/Na6>_EC/RB\Bf2^Q9Q_@d3_OA=?U5#e@a<TgD)
A9\6#_fa2W4E;E9F5:D[?dR57?Z];YB]OUJ-,S4XUf#:fI6Zg6:ab9YN8LKZU)WP
(&cgP+)d^T46Z\Kdf(-:gJ<F-T<P(^X\abI2BO#=2-1B]2gQ@@6TSW5#-;/g9C,f
OC::F#I^1#1c_RMY)HP4.Y(6:)Kcb-N_&5.afFZ4WN]0151dT-JRa:;WPH2^/EP8
fccFII,(XQ&QJG32S5,QU#G).+>_Z19f)(\\QQOHI&Lg+NDWOBD<IWEV^.]@36b8
V5I;ScQU:NI5b9[313#M2L&&)#=U/YC)F-9I_3H1Wb=^5,806Z.?>/LOSV[#:&K_
H(\D>e01#FSc>;9,\]Jg#N/Hg.]d:S<>ZX(aUAI.S-9Z7JT:[K3-PUOeZJ9Y\4ND
G=S-Ub]a\N@dS6D&Mb?02ZQ^:@Q0\M/+_89gdS:0E>VR+QIb?Be2&Zg;^UeH/IEE
f,V9,&>8Q=\5X:eeK0\ad\;bRAc,VT4>/]GdbGgX&BD&EWB0HNP;E&GP&=_AC25V
AK:[<GS:?2)I9.BgVPW06#T?\^1Ob@>U:X#XC&BI&:OZB-/M<Sb@2LbQgHRf3dT,
/fM]e\.92M0HM(_S,_&+d3)7S9)@AI#8fA<K[a9A8GZ=@-2X9:Z]L]AP77.0A])9
M_1+6UL72/FNf<gV#UcR6;&?9ME@Q[Q/+Vf5E.aUNb[B,-BbcJY0PQ0V#.A=,a_D
b0K)I6BS4NUJRXfGC?cWfP>L3MHCM+,;UbMYY-L=]84O4=/(@-Z&THZI&^+]R=)_
ZA]H8GSbcIZ;Y6e,dc5I,I(2M91-).=b/a)K&(1UE2>_9IDIUbfLX7F8Z6U2ZaXC
]8ITC7d:T;)a>^IJKL.JaG5B<<AGHQ]5&X-ac3]GULa_RH;FSb=AWWK#9\<,2,FT
/c<2H<DC6T^WS-=HZ^H3FW=UeZ/#B?HKMX_8NRAKQ.74abS9eg><Y^2/(=P]0_#_
6c^#/BYPH9?7AeV-IP#O[03ZcTSRLG6HgG6X4?V:-Z:aPc^V-d8.9?AUd9LD;.7E
G#>QP4:M.c33R9g70-1U&>aM1@]eQ-B(d4)ECg?dV/cZ5:))>FM&W.KYeT00)8P4
I,Q@O3/2HKdGY>V1#JGGM-2gGH,LEM&&,PP(=]^Sd_;,VT8dC+47ZQFVC8QC1<f5
#-:E;KCSU<>>b=Df2,MRIP4OS672_dVGW=E5T:(ETUA\[J9C6#gEGS(4=WI;V_\7
.Mc6K=8.=9LHWeAE<OdB@Z#(D+]7QQfJ79?Z&VCZ_MCX]E]C?OF9c@QPT_B<(9MN
8EQGdVGK@C6/N4e]O)-DWF_JQ@FMCO+G>V?^PK^Y#\(.g?EJ[1++;>[Qf?W:AI4^
4e60d?4QDHBXb50<fLYC]E0[c5RGc/.+d6,Zc<3CG2:W0I1_CLQ21OaV-)7cG5))
0Ffc#e3OW[NNgBSfWa]L6#T,O[S^>[@74EJMWFL2M.XbXeBd)ZD4.FbaWP_(W6ZT
L==;IaS/g1)Q>]RIS.RNJdQ7Z/(&B?DBAc5G_-\W:=&7V#.T]HW>U;U->@Zg<fU.
2KG>-/fCI#_F?e/G4=DA>b5:]RMZ>+c^+9SV5dZ6(6\g1DGNGL34K.&;)?6SG+:=
A[-TU]4+559LXb<e]BD-QK)#(Z=gP4?W#=#1Bc3VdF<;<\cEN9S<H0)VV<48gQFe
C]9[<=6g_4VF_&FR/-PY@@.8DAUBXE5R9Z3^O(^M+;6PR,GY:O(-b?:@/aZG(VZ0
CH4W(@-d#96+?,+f.I&@20@^=\gR6#5CMHS_MgPHSXMU0;+S5bX&DJHF33.-2Y2E
e52TK?0\BF#A21K36&#.\T9=O2DWUVcM06Ne(BX11fL\Z;:3D,9\BBYcWMW<9\2&
Pe6^DXO6(84#V6FC^]LV2HSGLV/1_bWY=0DP+e7TbGY)>M[(1CX\F25V&0_V-57Y
YXC)C[68(<N6A9-<aOT1fA,E&5_:a4#5P0;#\aIK3MSY2>03#)Sb&0[V=N0T7eZ9
1IQ4d9#Y)fOA-[FaYPY^UMG&<JU?\G0C;)]?0P&F23cMQf2@eHW?WKS2bT,UV>AV
@^&3g&>JaVIVV4WeSAeF.):BKIJC)S,S1IKUcf2R\K).^]LC8HBG>,M?ZPUCY3=W
+TKG68&6P\C=S977OgKO7W5;QX)0+I\K+P]5Yf4Zc4[]VO&HR@9dRKR:/&=(6g<f
^R@b<]a]N4Nb#>0\6G-)(NX?c/]Z<V7:3)G.:<>d#Qe5=.YfG&->DO6e)\,_cd=a
X]D2_/]#B/;g_2HC=@_N1=725[#e,@:fY3gO_5dcc:ZI04a.gY#@5R1Y0@cMI0\Q
TU>44QW/#<;</&aM=4AHXZa3Kd/<Y4Q(Q4BK1B+LF-03;6WPMC&G7:VWF,=dbP:M
g+R+b&g?8F?@[P><53eY/05J0-<#O21N-H2\EE>+TM#e)/HfBL0R[Ge\F@FIgM:g
-ebXBCGg8cW\],?<eAYRV@=?[[-<JZX?^??:F@HSR2U9d+4E&A(<^RIAf-[gD=1]
H=ge5c)MWRZ8Ua46.IH<SO<V^AeM-M1\65<<J7=B.6(8Y)6LK>OA(NR1FYZ+_VFZ
[DIE/G6@^_f_.V1M82=0eZN[W(RWgd:aC/e1]@c/d_8cWY0Mf/cZO&&a^H>JTE&=
SDQMDHY?):_E&=T>HX;=WW)HE8MJGC_HIMg0]#\28IZ#SGZ[Z:;UH^N5-BW>QIGY
@egbE^QQGEAbP9S+0VPWH#V?)BV0E1a@QXM/HR8bL65c[J5L;1,C(7F;I&aOBAB(
K/[))B@J[1(+L1/8?RC(Ne_@IeG4Ab?TVCfLMO,]8CR<^I<H1_7Z&+[WN0HZV+IK
c-49JY]A_5(RTX(,=;X9CX5T39^PBd^T@;8Y/O/>D\+O6>Y]HKMNP?&F(//33]-<
e6-[g>B5/fY17;b?66][#/(@>cJ8&CebRaaPbT^B5Fb-.@PNbfgLI&UgY<@9)I<M
K>UF=OLd>:aA&?69_,?;QCAe\4c\&9IXTf8f6-(Z_CZ8K^a>&_V:Ye/<5>WKC20K
(TfCT;HeeeH8?0cfWfA,IcIT)XR)<aF/dUS6?@M6;]/UHC@ODgPBL31a35U7M9NE
\(a]^N\;<YNS2P5Y/;684T&L8e&P7LBBT&FG.SK[6a#44@R<X2g:AR=EfZEC#g.A
(EGXUB]#1W7eI6L6abZ\]75R)FXcBZbNA+a24/\T2a-=eL8,KO9GIRMB([eHRdNF
0+==GVdLYEP32BcE^G0K;5BVR9PW5?Q;P:fGSGF4MT;VV\F9F3_T?Y5GFQ0CB_E^
[O.^NEXP1UA@AX0;//KX.NT,?7PSI2V@WK^3GQ-TOE>\;&<0#495KQE&>J^<_L\)
@ZLSF47QR>^Ga-a?)\bRO0Y63,CL=X@\0J+&5a]\Be3NRUETaS=#<W)gSI60-?Be
[)/4aX+<?(a[RBWUVIFZFb:-)aHZcB@geb\H5CSI)EA=f8g).8Q._/O3G_4B\X1A
VFZ8()8-4K8O=6:Qd(W@1=7A2cZ4BW?,(cR+(59=Q/C5aZ^^7?UgW=)Q.5^0Z&ZB
UP#X@6^6++RQT/IeF)QBD:\;KJb-+VF/U?F-)-#7L6K7Z.CC=.f+f^J6N&28PFI6
TO.>#3](+<BU>7HM-9Y>)e0f[b=HZR_.e>T2:CTJRJFP70O2P99HI19J[T(+5,eK
:1TPgP[YK3T5WOG7].3&e4eDV=&XL/=d-B5aVB[FKA12J/Igb[J^ID7\VFeE4-1<
I8X32Vg0TX1WZ/W]^#ZI+KNb=[JSC&X+gPLSLMN/,;=A4^?=C]6.-eYEQBDCda@]
bg63ZKOQ;(^B;<^AUIbVO;LeU+D<1/4B27,9Jed.]M3&98C.4-dD=S;(2MJQCT30
0<cF&==H+[R,&#HI_\Le[;7Z<-KUU1]9JbfM-\/e3ed,2X]>e2Z)VJOE;J6&eP4_
g7DH?egHKO0D;Eg.&W+gP=DU[<d4PQ]24fY4Z6VG#8ED[L0@SE[E_YFGR>W0(dW(
[c:e#MQ7ee^Ig:TH;HdNVN.Y,4OaH,5<:>/G]_3;@A.)@(/0e=I;63b5WP\9_@[N
HME,::^?&#<FW=]+9=?>dRDgU&=7\EM5^^IN[TJIDHQF_S5J/J9=F^0ZLbNaGfc@
O>^)3&GG0OHRdfW_5[RK3+09LOM0IT:]_-]E7NOf(M#\2DT=A,5P_Y>T(Uf.QTd>
]==5U&X#I0]NR8>5<(?(,,92)<#dZ=4+Ke1Z5/6I>1_VWPLS;DD:?S]NECHO?5??
-T2_f?N^fCAa0cJ_I@/,044;2=_IX2c+),H)N37E@O_66L[WQ;-:7a24U5[cdW8Z
STW^6@&S4f?/g_4J=bZc6-UZJ:H48B^P0=gaQ?\?JOON>f/D.2DM)^)Y>D.TK9f-
)\R7:SP80@]Pde2+Pb7@,T@f(IL0c(58^\@b;UbaaeU67eS5^cZT),_YE+_#gM61
5?N&15]]X<EAN#DE^#Td6_+;?F\,@1F:\Mg3@1f<gY>Z6/JR-+^VOX60Z?-<-D/g
9[A2L.,PGE3LBTDUVIZ5QJ>73Pc/P=eK+f#IHS3(71ZPIU_NMgX=bD[Q>-=5YQ&L
OM1.;YUJ8HE<N&,C\;9UTY7W2:[+MaC>#>+&@X/03NHLNH,edX^X[8_)XK)B?O6O
>4I,)@?PBWLI]ULJ[^KMSO&gbU#7OJ5.H:3\#SI+cfW[Y_E)?DEP<S:^Yc\QC^?.
K#041VEA<#_\^@Hb^]63YB:Jd5S:IcQYA[M>/b?)E)[F(B^:@H?RSb=B60-TY:;=
873JO)HY+CCNBf/@Ag51@C9C-9U,HC:R-J-4VRcf-^VC(;A?OLYMgf.ZV?Ab?NVW
?fH7T?9_9)[T158M@TOE<&X)?.:b6-cYVJA<7Hc1(T8<R1Y1)J66)_JS_-IXX02d
(22VPYM7X?b.<]<dR.+Of)P@)T7S<0eTJa=_ALKL532]7FJWV=+;XJ16B._73/+K
E.84-d0-H51EE9\7IKCZ,.>T_>5^MNXfX-/dd@+^Q4@=;WCRU@aY[f)=SX#O0#ZF
3@8eQR=?=]HG)>1+[(H=XY:;8MQ?^50]7PEEc8T&?M<fTG2@4-f8:[N+@VbUgGcP
ZOCQ/I+4I718?AQ=^5,=?;+f]Iae]KWd]Y3CCNFSSgYOO\WTG#<a_VBZZ8ESf/?N
ZfJ&2)Ga]HIC9JAdC^<N_S?HDLEN2X)a5@I+8-D[8A];ZaNDdcT3>MF1)dIYaT.M
CC:<aG&UD?7&VW03O5e,#.K/Ea]]-^a;?c8dS4dZ.(d9>6Wcg)19VW]Q^5S:W=DL
?6/PIBAe_Q.(^5<^Vg>HRF)4@-d2C=Z8d7.15=I97aa&f3@HUZPE21E6VJZ?cd^-
A4K[aRE9b/(@U]\_\-CZ8a\WZ<FZa-T&,J#?Q>2K^//I1=-d&/JMc[7cI,\UG>&W
Z]>#+5+f,58<SX-VbWR3f8W7VBce.DR#d_PO/CeNa&@aQ<[SFIV:SH_#+a9ZP]-F
Y//9RcJIg3cN1(+90^STW2:,1gWK2FA&fU5_OD5Y\Z[AO)NA]\#1W&5S]PFQ@)<7
+_S]&BFefUU4V36VVR31Y_dTTa[T_7\]JWJW08<P8^I<#0Y15,aDKI&T>eAF/CPK
\R<,3D2(81,KBfTR_>)TO2:3C\c>N;b[O;UG,(YV0.ZJ8KQf]V&eCJ52]N:PB2a<
6VF4^<3gf1#K2RCC:U8AUC5a+.Z[M0Q\f7\L<Af:)3@<MCdVJG^?D/7PbX0[,OfR
,B^P_DN4#S_VbB=I0)Og)#VQZW6@OaCdFA.Y4Sa+)?MHH9]@((8^JW?4Z2R98@V&
/)IVV[-A]fRdDGPH3D7)+H@Zd.JPK:dOI@5\LU]\5=+g9cRMg9+6GU-#&X-.L/;B
Z@7Og8fDR5TZDA.B.7W=CKbK@2Zb]-gRbQe7X&Q7YZJK)5d7@fCMH_f+&=:SMNB(
I\5_<1WVG6MF4/H68REdC](Z@KEaa()(RS7SB8/N>QO=?,RZKMHcaHQNeNH,bNC]
R0_?eNNP_,6[]#;+]_a^3F\1=K?3U4Id=7Z:#UMT;NZA))c38W^J6f@L;SPgM]<4
9&ZYf_e7H4PI1NICR).QKS6dG[Q>3Q<BHfR[U1=QTCfOBc[f1)YSfGS:/^PccN;f
TM<_&-gCP:1F>ID_,_9d-\9>S4<0e5]Y5b(0cg]2#AGD<25R[-1<3=N.]B?,9:Zf
4:WVXDg[cBE]5\F0BF3_HE)>A1EaCOX[gGa3=4=4^bO(4L]CZ/UI\+@55.TOIO1J
+99=a/X9M?4F/?U5,&[<&NURPb=\[WDEDXAgA8bP]?)N9UK.9d+4C?J/CP^29\^a
IH7b=6)I:C.KFLaZQ<42]?(C/G>g(EV(Y1.PLNQZGOMC;ISBRN3#MK4;8RcZPATQ
.f3[VYZ7G@N4c5.3e>YG>F]-=@(+=1f+)ZH5EIMZ2#_^\<]U&0J[,7_Yg1]?W&QY
66A:@@=KRDVULXH\VeRaU@bfS>LJ?B?<H4PU5-0]IL:Sc)@1]<-@]0]67I:XMD\(
4Z;(;cNT0?R<eSE(e9FEJPa(M-B\8g&;L;++L+1:]f75IRLKU8A-_cF8;#6T?HfK
UFa,\a_S-dG,fQ@]=_MU>[FfNK>^^ONSA@.+]<F8[#.c-0OI,c8;HL1Z.)#<9C_Q
L-4A5.,+EP.P7a26c+>B>M#6MdeAOBg8dL9d7#7XS?c.=dN2BRF]XH/Ce=F&NWQ+
f-5G2ZP87BM\0<b)g6[4bb5;VW;?[<=LQ3NM9R:VfR-XGO8S(_>fa@EfDeWD)&/#
^:FB5,)(:U==bULf0WM\)5G?Pe_S&3N01OOY=YKX&NKfGeNadR\L?Af&65>H3.XT
F.1#5g4=F8^b]C8G#2A?^,F&8X&O[UIGM:[=5GT:25)^/M4=5)Q4YW9FYVQO)751
A73V37NeO^#)=b)1>0VEX+.B\CGa1MX1<WGb7526dWZ&_Q,Y0X?;HOJ?(=R/,-Cf
CC;/2^geL(B:W)TVXR[PRcdDE\1D(T?NFI7a3IMIH[XI@X&AW:?bFM4f2R,)?Ng;
@#T\0\F;8Y\DN._8^b)NJZ/;-B5\6fH[(6LdI5N:faDfa:X9NW3TLdg,-;\#09R;
9fc6_XIIW,eTN7)TZ9L/QXJJG=4K:J^[PE17Tg8^D9MY,-I]<#aaGC^,=e-^Z.]L
bHKH>A@4^4+PK)KQgIWD=YL2CSD0D3H;AN]DH,b6)E4BHR34)Q-F+gTg1J5aB&M2
L6<_ZTfA4S#\NM^HLZ#VbX7Y)R2.206f@6.I^+5J8?>GT5Eg0dHGTU2:BBP3JB?J
@:SKOS,J)@2ULSDQ;@W-F:_2LL>(0WT/\R,5WSV-O/.?GWZABI05aTL-U0We8=e;
.?I>f(BKdHJU-d<_+=PfI&0?2dA&Pd>67O5,G6J+bFRYc(b>[F\=K-VFEA5^T4_W
-B;,K(VKeS:Tg1-^]ZL0K)FE4dg<.KPIVY-BF#@852XOG]?bg8QeDJ-KIU[KU+LB
Cf,H:]1E-4c,UD3FX?9a[NZ]\0).NC.K#XQ]74D=S50-66(fQNZ06Z;a#=GLV<[e
UYIg5bV,MD><I;48,+,d>,(cC_\]2[^CRPZ:&@V==TB6_(X#4Q5[ANNI.QAP+?Re
8L5K>VSd8T=4)Z#9YMB6faR^Pa-N.deA9W7g6_,O/322DAE8X>aRT2+bBS#UaaLT
4=)D9UK#G>4Qd2[0SV0L/a(4UUX:-3K]43T]TM=J;SEEO]XZg#gPH.c8T.fFV@D7
UA.=:5</+^G//G[d]Ucb>dF6f/+Y@Q<.[H,b2:8V0P_FPS@DdQ-6W[1\GDMC^_U&
]<DcLH,2T#PC?ZUR;?.6;FK;a6?GgN>_^gX56V[HOe#Y2K4UF59:=FH7\E1S3_NE
;<T6A)27;U]L[Ya;aAQQSY-C48>GCZggST&EISFFB9,f<[1)d8a15E9Wc>fK/6D4
7P]7,\[.?)\d&.2eWOM/#>,/(ZNA+J7eGT0U.:B#<eVd9:4^Z7ggO5F.7&<FCc?K
OB3?(ed+D7\S0L/^X@:_V\HTVb&H(_gNE]Re/U4AR35c\A_BT3H/3G]gDfLQd7[7
2>LE;5\7,PJ-(A0e_@0bQ#eKX_b\aX^M0HCf3H@:QUHX-X<NK[9T+eX\Ed\#NTBM
4C0\==EgOJLO[:RZ?XCU7#/U/[T;SBCQ;DFKUddDSRfFHT@(bD)>I4HOA6@0IggX
&:V^L.H2N9MTD;6MVM^e/c#3C5[-?8CZfK-K[?I&&@2YT]XAO8@O4dLSJDM<IE/8
93d6AOK2,79ZDN3LJ);gOT+USCFc(+M80Rb/OXB6>0[dfPP,-KIS3LXI:PQC,P&[
e9WTWC^OOF4#@dVce\c^W=f-/#5V6_19RA^.J=fPM8dEWD&YT/U1DGH^A@c&<+S)
0^BfXd\AAQ,J[Nc:P8LgIP+Y,5#eI2\6897=YP3a6PQAJX@L(#c:<<G?HT^T4&4d
Ycd]NWIC:PLN3J\@V(#:(ER(;W?T/ZY7Y^ZF+,#a?2QJ<cI-BUE+8&_/(9UI2-N0
\)WN6[H/OQRBDX0(b-E?2-4A/2CS4KIML/CWLM^>VCDY)#dYb.fA:?M?&&F(HFf_
P.0;fScaNaFAUL,G(f&H6V4^.[8e+&NY>b6I\84V7[F@BTI#G1d@f4cUeZ:P4TJ&
?Z80b+-&DB#cS.]/^V[8JF\.O)LUO=cN=I>?M<0Z^TJB&2?d1DLPO17RJO\c[]EQ
2G@<>&]:,V=5V>G7,@L7e>WB_OXUfF5LO2_6PKbNDYX4+A,g)##e6S-[KQ@9cb&O
-O8QWQ?OT<;2/^;R#7.1TUQ;+B0L8:&>HZ;0_eS-#(0bU4Yd#)\4J=O9=gd\gC&a
2[E^?]QOLJK=GP6)aVe0.48U,@S#HKWNOX[^_I4Ke)32Ha]]eRK+35<(AgXCP-[J
BDKDd@0FF]8+NPUX(+\Q+0M5RIe14c@Z4J?OVBNMLN7KMR@P6Q0BdG]88N95.=T^
?3UZ3M\&B2_OD0<eUF#RW73.KRf3/=S\^53,Pc9YAA[#bSg;^2d7Y,PMRR2U-8).
8^d+V)P[YG^/3U2XYO.=-+R?6e71#_LNFN.P]RNE;(cX)6(.+HPMf7e-RM<(M)f8
H6;]HbG-\6CO+J\-FJ5Mc8C]-;/AROK(4PC0[IRU)[X:8JIgSU[K4;J+\(Nae)CO
<HI6\_&3_SAL=J)1VDH@GTD]#L20E@(U]GFJE^b,.0L>e;5<:IG:#OTb^NZHFdR>
T5OPF7&JJB?E_.6NS&X@g.4dZ;CK1H,I75Jg\U10e)[,+DHM7A\d/XIWSDPOF=(<
YLT5E:R6+FMfL=ZQbX6f0+B:[IDG@W(PCNNDa;;7^16UKGK9dcC8PN97JQaR51<H
L?5GgP4+?WF@NWbeb/T66.,)bUM?&.5_F@cUdRZ@bUcMLCb96+O[;2L/J?=JORb9
@NF64NK@&,4&##cQ0.5WJdTUc0ecKg(Vf(PaeE,<-?W^BQ32[ZA]#d@_)/eXAN_g
L7I=E1[O2FHaI-Z3ARFY^[L-RAQLTDO+S]1\FbdH4b&]1[;.&X1bZE=B,@<;L8\6
->g]9d/?J_OS8;8ZML8K&N<1S4JW8]d9Q0M[0E-#6Qb,&SRI]N:BT.AH7[U(3^RA
G:Q<7/g)P0WJ:H3:-@&,e=71&P]gW;236T@T;/[6)8,1Y[[[DcS5c/JIc=/e2S.5
_U/Aa0R]A:,^&WPfQY[KPXKN/N\S<eb>:;K/:CA)?J#:#\^1R76,,]=c@M;f9Q6c
BRI@US=a\fFZbR:3Jg:K7ff_I7?FG1_NbL:WffY]=DIMe93G,-J-aHY>Cgc;VAc(
TEPWQ:D/DgL&E<DO)2-aEK@Z7@DbZ?Xb3gc^I1CH#Gf2b95V^LMSgNKV73J2G2_V
c023#W?AU58.:T73^feJDE46(GFLDd[d#/@DF6^;B,[)70\T>K.,ER.S?ZcP3^-@
]gG=He23Q<_UfQb)4GaIAeWcIF&(U+6T@9N5M+I;-SNS,:>GER8B:\CL+TFMX3(Q
g>T;@[62W4G+2H?.<3;e&:3aF<#[b0e#?e(F=2E,P?;ZI_:-Pe)&=1X9=LOI[EG^
P>](#WG(WLI:&>G-J5P&_F.YQHbP]eTd_,.L:[2f?2CGDT2B?ZWP,U^&f+eO[+[,
L-+=)>X=UHAN&2=c5=J0ZNXKQC+->QDQPQD[a&5M&O9DE]a5@(-c,L[cPYD=&EO,
+Xa958bQW/OZMdYg<4]bKQaR#]eOB3_LPbI-.]PbJ_7@c<2FE@2A>DTb\[<?fIDV
5,OVVa^PMJV.9J1:BFZ-eaA0\c7NcT\9.fV+[^LZ3A4.QQ\D3B8S[+6Aa]US&EE7
&AcINT&-fD0>#aRW#J-T=)(\6C^NLX04YU\EcF7WE<G5LL:9)D5S4X+a]fGe&Z=G
([]]6MGU?Bf,DdD>X^/G7_+#F<T6a@5+^4I&K<L3^KgNH;ZQ+E?LN\1X-b63RS14
cKOHJ\Q7#8)R^4OSYb>4TcJOZ^ZJTEMe]>?-,;Cf=/E71g7+YJfCG?>N>7K\TB3a
HUF5HM[I1e&f9dD[?V+;9;bfg],\IQ97JR18KA5\,<OT.D0][cce-TDe:aE<>0.S
f924\&UG<eT8e-=IH(dFb>cbeF3c?-&.L\#@&@T\;F-(^L.GX\dD8Bd776&483<9
6AVY_:T(b+[,+GBQJ-c/0WTDb@f@Zg1DceE<9HET#X4f2E;UaR9Q@9Re?ZB..8)S
M<\:L=,Ec59#(O3GYb0=&ZTVI(S>J?@ffWJSDQ)P]/=@7We7#MS8\B<=P-_IeIZ;
TDXA4Yg\KXgT/+f8I9gW0b[5;NI104A7-@>C_.B7F5Nd:@Z-TU,\CI5\Ga#1DAD0
X([I1_:2.H3>g)-3J99N&X?N@]eAR#aR-Y0:N13[#ABK6BO@;\W^g9C[];MU0+Sc
T3E1,[,T@?e_Xb(,WL4_gff1/GCE\ES9&]bN7VS=6@H4Z#6HA[&=;gA&)3;/=H5W
f8.+I+NI:WVDDZRXG9G-+<+C>B63A=Q?E;/^1H,5V3VCDZ)f2UCJL#?a3Z;9M8UN
9OIb)R8)&(,@67Z2+:f@f:R0A&1Y@)^GT\K^5SbW:eF#3Aa+H3g,>):>cE7=-bE-
RFXE:\GN/g7O(L+7[B8X3#C+I\(U2S7R)/DR;XKfGL4cNO237FHPe^Mfdb@eA27X
K-_Q)=(J#/DdV^N<L-3QN7U&E[-F;0B2R0/EX6DIc(/]:e>/S3JQ]7(E+2<Ha?[a
2a=+-Kg#U0MI8UgG83OPT=FDA_K#Q(W110dTb;/^aQ<464(M-N?;@-D?gaGf\9ZT
T(#I[R;,A\b:=7JQPFATgN5&Q03M7Fdc/L3B72gUBBD^F@]^U>7SS;X/UB#Y].EB
;aN(FJYS^B^/[X@AB8(6a56[T##WcT.Jca(S)X>):]QfI0@D,N@<P5Y^J5ANO-d-
4Y5FZQcf(Mg5X.T6L0ZEI]C4EcO7Y18>I7OcYBE>0Y,+H]35H)GCSJ>Zc9\+-T=[
>VcD@@bTAfY/[,3O=95ZL;EW_/ZF?:4X1.=9V=,@(ZP#H_04FO15NF:Q#,AS:A:[
F._35IMgNG&H#eP4?[IQ7NOT?2UGUc2^DJgaHCF9(dQ1GA\YbT.2@U],-L_UbK#0
^:)+agdT6d?-<0U^SU5[]#a34:8<2C8<?aB7fHK+VI)dCM?-)b/]=S-7b=B@b3Ca
OZ_M9>VVfK,Y:MXI69\V;&DO,G<0Rf&I-RO01H;CZ(;WB@1S.ZUW7gg9b;Ga7])d
YIEePe8Q0N@0QJ4JZVffZXX0R9LQJ4_RW2O01P37FfP<W241#B#_3BU6/02.;eZM
X3Q_I).&RYaZe[aPJNCPIMOV+Q,T<3A;HH&&]=A;/09J0=KGRSYGLTEN0MTN.Y08
d4c/#)bNJ5-HE[adI2Z7TbbA29YX7;<.+>AI84LTVg<1?;K>DVf2^IL0//8YJ]aT
63QEeHWX-4OL(SX\FUQ:ESf=DDAC=Egb8<+MBG:YW@7;K_b.Wb7YD8-Z]^)_aFg#
1MU?&M?IBUH>+)GD@X&g)JdL8N9]?<a3L0Q=//&#BOS@G52cS,S<OK^WT<1:WWQ#
&M@BKX&6,6)-OXYW+FJ_]4/6+3+\W1dVH2W(=2WGAH\)_-_CHca@ES:VQGgfbOV<
C;X[gQJF4DMaag[T9.5L@gR-1MA29#60L&g>DbaP7TX(T)OOdJcQc@;Ad]#AFd+d
V[5D@g]-5MWcGKePHcPgV0OLF64VS^6]Y]P7#d(;5YQ@-80^M+;3=LI=,)b9SJ+B
UX>VG3ZNWK<+J]&MFPCOJSH:/BP\U4DaA7?(H50:KTH\JQJ]K&OC,I#6BRR7^BZE
Q69)>eXbD#&Nf==S+Q_HNA]Z<7CJDR2[U0&0GT.(U[NJM8SW(C-O5<TJ#8S\U1CZ
Ec&,LEY=FRAIHVcKd(NS9X@_X-8F8JJYD&g[K:JA2E9Hf?#dEQ0D=+^P[((D.E=(
[K0<UK6HW4[-U:/<eaH;cKf(^)?Oa/W\a_Ed0/9&0dF.Yc3;dg=&0<_aVCV5d?Z.
O:B1c9.5(4+aBC#W<O[C;11/)VC93c?6fTUINA5@fg5E>R2J9978:J=V@VB04E<,
1UY&E0QMM;H=]8XX=]^X9OWH2YCf@?#K&A;W^-^c69T43..^@:(H<?)\aX&6P3)_
;/.)ba.P9]6ML1=?d195cCce=UE7aJI7fG;@L+QGNBMBY=)I]0b/H/+(G1#[#8fT
gN,2RKQ<Z<1L4YW0BT1OIJ&Ab\7.,P)7^T]O7+UGSQ[ZV[X\LT,X&,134^UTYdZR
Y1J3LXgLJ\GBTC.7W6@gNFb1\Ac_846cO)8)GIVFX4)=6NC4MVL18f0-CMECF>CV
1S6^(S)TVM1&F#6)U<83?&,MS;^//gb:^ZB5B>\T+\I;RUMZC==d@I@40/Cg[EKe
03R(^O1R71aV1W[^.Y=S3_P_O-3^AcH6+\IQT2>7f2A@9Y&</Z=FHRS<[\GT[>_:
J2aXK&Jg/UKCVdKa>,>\dLY6GK[NPgeYXO/4VW,[1?#I_^Xf.6EPdJ7A&K0LC#a\
Se@Q.X[U;HWT5W-++bZ9PO:c5YU4,.188X2Q,UOOD?49@K,SXNXD+_I[S1c?-8Z4
F:4,-8cgVBWbK@&)JJa\;3]aK4d_-2JDIBfIDA7G_1O^7,&\E1&<TbB612DccT)1
(Y1bPXHVd?TD-38;DSe^&P8d^1-/VB(W-Wd5fb6I1=.1a&I6WR@:UPb=ST(\_cHF
;E8-?&VA#F.T+L4Q@G[7S_2]B4\X:O=fc3HIKH(-Fd^-;e&AI4KbccO_CW^]0#-2
+\ebL8N-geUc^BA9RV(TK5.d&34g@b[@B#=P9B,Rc\OBQKf7]gOWEb7.P>#AXG0g
;8JKF1Z6:KVDL6B<Q_?DNCMZPS[_#MfQgZJI:+E^FUfNM.@Oe,\>KO)8/,T@cRVN
^4cIR1<S1#M#,IH-e]#NVb9\ZgZK(/-9RPKeO<&:HLc7L&G-QY8P#NTV<5SZK:,;
0KHRB-G\Z9\egcOb,3OAU[=1ZAL>8RKTOI^1_8I?VT^63_BAHAC2-T894PGKI@N,
?0\Wf1PB_1(OIc8SLMZ+O]W?b8Y@.23<Y4BgPP?YcT-@VYY@OG5APNGY+:2AISLO
>M8]6_L@#4-H18TPB/=\X;R^+dAGHf9V+63\d94/ZSO?c+C:Q/e-I(VV-#b;-UMB
BbPHD.^+S,aR&,L)D6E-_6fC-3GVYYP(8G/4Y#)d<f0:L8(4L_;GG_<#-07TE,,=
8gG(:GaY2<]S]>-d@(HU#KUZgE\eRLNdV]HH?NXW,\VC\1RO.\/Xfa\1@?-+gEQ2
]Z4aH=3P(gD4IeB\06Ga#[NVD43_U9BJ5/<=d_CD(.3;5bY_4V9\R\eZ>edEXWcd
4J:0QX)=N0UIMD0L86.U#-1\F4MWXa<#&-7N<ZQT4:BO:P5IB/&7QTV[@ZIIENBS
@\abVIAD^+@g;AFbRd^?N?A03(e@8VR,.H\,@SL?K@g]X78^GL5FE+]W70J&SD&d
6->JA&HGP=^P=DBUUM&d:f7H]2^7DK70#BIIU>b35>cS:S0-BMX1A>FUJfRRN^3S
1Z>,6d7T0N380-?adE.##Y37PW#V;=cd<[ZP,4LBAP^U&F9025b1ZFB[\CM&I^/>
#J2-g:0Fd)N?@I7X4-[[>^E5-;RVW32<bOA7V)B@E:TdOKZ+Jd1_G,_WVU\F1P3F
I[9O=\\@TaR2#&WO8JD@/^GDS.+f-+)N3#F?d&cAe[ZBU;F>OR37.T8FeU(C+2SE
L8MFR.)0X6#Rf]8dcJbfR=6?U?Wa:b2Cf+.QR,K#g.8Wg<N^\^MSF?D4+EKG\5Da
=KB&>K5H6A@4cZUc?3=3ga0e1]b#ARAb?FFWU&I,aQ+EdBC2-gMP[9T>6aXda44&
U3P.dYIM_fTJ;AD;,J9#O,1KUSKP>e5H1XT;Q>a8[N19;36@7W?I<Q>[N,HcgHa&
^JaC5aJ)YHAFYS+Mc_d(Z-R5)?.OV63ZGD>d-O/TQ_1MC>OaVEbfC@Z+7ce>I9Aa
^+Y[>ZMGPZ1MB&@c(;=EZM7<99O[[48N[&ZDH9+(K+<WZ@eC?0X=]G]TTY^c?3a]
+E.<g;fAUN<P_V=&d^K9C@c;PU3Kce[XLSDa[>dRH(fLL^)(ZN,E,)\\DEe:A;M&
S?FR7DH>Y;G@35XBPQ\RS4>:NT6Q)70PSW=WM4XI[bA.[gS7e:A/;@R/DU[U)Y1X
f3A:T0d=TYWBS@^ZFDb.Z:H=<7V7V]D<:WLW382\>NMU4K55\&&Y9>8,4A0d(MF@
#BUVfY#H,/]6KKEF2ZS++FJ5f;e(0E-L-FG\GS&TgfD(IJ2-@OV_,@@OdT4e]SQ6
67K.4Sg9<+cAGN.>fJST9C^bdKI)=XJ,18QGR,BOH-6Ka8]U\<:/)+AOPH59P&ZD
(+(5:XWc;dI0/OBGBd/#B94g2XNeZ#gL-d+;4]cd2+KMg5a(g^f#d0@2NJ08@6A7
gJRE_W5;[2Q/4IW<)GX[AQ>?PQP^\Q&e7/Gg,M2ANP7:^RP&]4PKJ5O_f<EV?[Tc
393dD)c6UbP#@>W_Y/&<dQ,Ne<[Q#LHSY4:\dV)KL/(AHL+IDMGRbOZ=gXF&SAN<
a[eZ#)bJ2GYPBW8;Yf+X8;K?3,IG.cQBS)BL7.:\gW=O#DPF5X_TAYKYM#DEWS;.
dbBF0/FeBdBFW..R38eC<faL&E4Y\Y1(=6Z^4B[23=Tf72^B4L;5XRaa/.SSL3a#
gGO&TR)X]J3;+0&Y.=@@QI7+HSTgIbKdaQD/YFX+R+<4/NS8]?4#_DNg0::;QI)S
G?J4R=P8CeAO03T5WPER6ESV=^BG#K9DL6VJ4eG[V&;0F0-7L(&E]FZ./WRg^EX+
C>@;.-&gA#LCG-<YI29(9=Wf.EA@OM87)+4Z4^DE/)TZ-YT/Y24cZQb6X;0^_eL+
AJF\A]YZAfS\83VB))XYB/6G.S..83a).Fa6#6g&&^]VG;@J[fO;eXZ63E9ddC_L
Q#NO3,+(#IPO2#Hg;.?e:BPEfQf?@FZBNg_CLfK@B0dFd7F?]<EWaDe,3Q;b&--Z
-G98QU4,Sa:e59<\c>7_;AU3X[;I8)J#FJCJcMFVM)FMee@>KZ>ZAQIKf,Y#]?ZA
\C\+V._b9MOeW1^V]LY)^3--:IOIA2@C3L+_V<X8)Z5NUZZVBZgP8I],9P])S)-N
]HB#e7,dO@dD9.[e_:]HbSc(=]O3;X3gb#KS4MeVeI)<a3cO=aK<gc5RC26Q>U<]
[4adRdEYf(U=2cR#.FLL8?f5ZBW:W.GYS[\d9,WUf7B-[]?=>)4U0[gNG&MN(M\R
XFLRN.=MG2]e[d-RA:#\[>6^QM&;T@R45ZC-AdTK3R<WVBO]&[[;7>0H7:aYT^6<
JRUM^BO^U]d;>1?ALW/VE)SNWc5R,bCLR-6SDLMd@2\:7@^)&S7C865eJ,\RW/F9
[?>g.0[df+5]6dc=&5FOf#B8MX\@;W=3P#2D,Zf::@Y>N32J(IECd>X9GVGN3(Q=
5=6;ETMGBe+X<>#db]56L<R-&2>=D#GFW[ILEM.KRH^cN+[M?/1ad7AVU]DC5[S<
/1LR-KU04:,R8J0-.TAVN<>JK:F?T;?cA3a^77@UY2I?7ACcR8HL__L=N8c_W3d@
gf4]I,1R@4]L5Z]S.Y>C9^&&\95+SHDeJJ/;^Y0eM\#Q+HFPd4D3##^)XY0f&?->
3/1)N9dYR&S]&5)\95#,?f)9(R3[ZbTU&]NG17RdAbA)T#U]&Af\XAJ@TP^6VC\=
0?0SA:?B=1#;_LV_2NY(+40PPZIP=aK]d[CP9QbV&)D.8VV-[g1><0/bDI.bO@FU
8)0F#>b,8(TLD<GQNDY@+9.J,BN?TQ_T6@D53.<UZ4^W+4>L_<0^249Cc004W[0:
//7^E8XYZ09^Y2cMMS^01[9dK2\#+@>^LZ+88)-O6D7TYQBLO3PSfLX&X&cKEKA-
VaRSR90f\Pc5.?3_dc4Se^gYS=::A=@++6a;1^\0_4S@:HS?TK70,&ZY\fE_+#8/
[A?KX4.VbL0I(9g=YZOKB-7HKQP2G/YL3;OaU[=BULKWBTJUNKDB+gFIF8&:Y8/Z
@P<0.#BN_>F4=6Y4d2P4_fJ4d>:J\SY0\:\RSYg<V,RQd4;#01QFS53<I[RI[XS(
+GQ60dW[eNXJ44(:89G[R;+1_HCG=?#4(/GA=X647gGQY[G]A#PI-GAX@.@./1ge
Eg[LZd8GPN<9ZUL7cRC>HbNN?Q(I@d]KB_1+NS0,MLCU:/9eaX]W8Q0&ON6ASCJ&
7DS.:8)VKJEgG&/J_f_FSMN=_C9eA_.6IQCffS=gC75.J:OX,)c(RF--FcP_F2>)
@,O)b_-(N<7@;K)GZIabH5IBVd)L_/7718O^a?&Ed0+IG>&1)+gRc@V-A]3(gLTW
(8(#K8<RfO.Y:,[0\VESO49dUbE.:Y]-7LD0N&K:N)W^Se/L1X\2Wb\L/?DYQ1:@
RQV3^^-HIIXXX+>4<S,_OEE]ef)85=Y.e@RcX\-,/D+dXC_1[K]P1&=UIK7Z&/S-
7=958\g?d:65:J^NQH_LeWA8#gTb]2JFe^Q-_WFgL6M.=9S.95R79dFd(+AZGV3V
3G5gbCL#2bQMea#(HU4W)HCg<7.=Z)GBVZK3^S3WN96Za>=M0LfcEHdQ1E>bZ;=Q
d-Me]>EFDI7FD^FbDbDR/e[^2&M3#+(\@L6B(/V\FP:4<QD]W^Z,c9-2&)S(E,DO
OL#GEL^33GcC^<<8Q#.[K;3PC,a8?XdPf9>Of5=8=M@JTV1X^aQ_-W\=I89IW1Y/
@gIZP09)f:C&=2ASdCEZ?VFS5C,C4WSD2d=3H5;#UXAaW#M:@Xfe375DE<[EIN^/
48ATa-5D,\PA-7,dNQUe9f@GMfNcF#YJSAY1=MPW37W#(#8RQ5df77@1Y[\(Kb_V
J#2BIJKRS(,eTdFRcS702ZCD4=9<cW>7bSZW]5fV86;3(M+G[?0?HCPP(1)WJN=(
)9J/6+8Zc^.JRM(3;=Q3dEW2,/9&0QIVW_dSSWE:5K99KGeED7).:Ia6e1fPG)M/
\U;9>@b_YDcZ6-X^RUW/R7LOgSU\W6fgFUeOC1NVH2J43cT#QdF/[D7G,9TR7WXH
FXN5?1LV2C#38QVO)a)X;53M,/RGQWLS+,4+ZFXM1dA4e=B:IXG23LE(eeG6eaMH
]#NM]-VW0b5F=@<aKISY>F][FBcI(WC0=fNR09H6.76?,.A91,V4]WTXc2&G31(c
5QSA-4/))fQX]eK[+7Q47gd07Y<1IGEag&PJ4\68b<f1:4g;HHfRN\=RE=8?bRTM
;f.fJ3RU^gR49KN]@JW&f=#\d#GF;,^#XZ;AXVVOEA=7f:]/P\31[7KKagTV7eBK
E1aSC3(a?93Z7]=<dU7f;W/Z:V1\B,N)d.&NSA_;SD\a<FZ6I<84UB+H)A9FQ0;,
FP-&Q)^?\,Q^.fO]WQN8[O]f.]@>^W0fH?g)(8;AQbAgKO)KF,HIYVPH9UN6I2MN
19XHSg,XefZW\YTWFQKNW0N/bD^\V@H)UZS?])^bVAeKRLNFgdT:>F@=dP3;?[;<
^[C3aLW.L/?L>]79)C6[D@AN7HT#VQD-7BNWUJQWRRSd)@;EW#G9N;E<=7P_N8-1
?WWHZT^@F#9_fUN,5.+_Y=JUbQ:(X^;)d>9W,J4-f&DKK039ETa&EW[)Q@Ub+B.]
6#I3+[H,NS\WFX:98Cf0aD60X#[/AFD\+_9];O\<-A1ZNgSU-^Ug@fP-3&eC,QXT
(P+;ZG07Z>Ib=Y3;=BX:dBRDbCUfL<CIQ1;L,&#8//KgFQMTIcNPeZ>1[1;HUU>)
,:[0CDR?+D2<4UXQ\HSQbSBAK2S&fZD;T?8)?].-E2Y,/c@,bUa?X48:([9HaX[M
0)W,GZ,-Dg0^JI8fc55JE,d,MR@FB&KYJ^V)OV.5[4=\Q0_&TLWN?,?2568?(Q9(
B:A?/7b,:45S9eKDYYB@4-1K1;HQ>WJgWXKD#aI1>W[WaF7HaE95\Ab#KMW32g5<
+YRD2E6F83C-ZgVIfc6<9D98@9LcO890G6/b+9aZ6W994Z-LdAb20BJF/Q-KI0J.
FL9;cQ:<BK-+ae93][#PW;HWXOXG^)HX0;FPWOR3f&-B]-4:O4K)CKKD.5b-dEAS
DbdVe];)CEXFH=Tf..30IEDbU.GD:\Eg[3NXCXXF.?&TBE_QL/[J@^O</VY]LY=K
d7E=;HYS5eL7W;R8-7+L7a22ZD#Id@RFL>)0DG)M_TEOM&2fQ+/EV4_e<CXZG,MX
H&IVWK6(b(,2AZ^3Lc-,U(&QW(adEX.MdccePJSbCb+#K7==1&2#GDFIZ&<PG6W/
BMaX0K-A;-1d&MP>3?cgafS3_\efUBWI;7__-/@.gPJX11YTb8:J3CCa^XKgZHN?
<aV95RTK_0(#^NK:3=CgMd;HMg2Q]3FMVDW?\0@.YdV>-\/8ZO>6;7?R53<-7:WT
<PeO.W=deP,SL5:Ca9#=F,,)[V<WCE)f\LA(,IM9Hf#dJN#^<SW+/H(8^8Bc//7&
U(^S4\D^BQc@)D575NGRG3J,N2_3L6e2;^/)(b,TP;8,g8/)@2f.e7U1[W4d\#e[
GQULfU<&20R7d>&G4EVDR;JZIEaYG3L.9GZagLf-HH#D?P9c;^^d]fJQJ4ZK:I.9
H_MDT8A+Rd(W734B8QU8HUYE8VX5^+>5?Mc<=bM7B[24F.3FP&fHZV1RbKfb(NNO
PL>L1F0AD-ZIL+LP.3FC=4&4d8,VQR;bI,1(B66N1#-FBEFM]_=EK#7)K,=,[MKX
:(d+]0,2\K49T&.R33YO]01AV0d,6.-NE_R47:+B86OXX9F@(6M?&G59?[&(KNZ&
SIL]I1;1eVad0-?VQIHR-1S5NH2RE<?a);)bbC&XE<XTgK3)e-XR.CBO)c9=:EVS
/0O&SPG,A9P\Ffb9T4a&P5M).80:ABOTL32Se0_E(6<YKNRAZ5UZD94H):afU9cH
OQ\>R:CF<Q-]GI,4&F3^E341QTX]5>-DXV4/L74d.E)ZH]RZELKC<F._aO,W4E#I
MQ@2GA:5OKQNQ[YI\-<aW<_g1-O7:F39974-Eb02d=_fXY5,EECU[X^f]<3.F;a#
)OO<9E[?JU;9]J&Y>DaLAI1dH&XVQ\b7=dLaC4aI0(^(Z[e(gQL?KVB#4G+1:SE5
[CX[gF?bFeHC-Tc4YF=b&&6/HTZ:4KFcaUa<#P.<J,2gf.)^_B?I\VA9&+Y._U.A
cFRR^&Ue^fOGHZbaZ&Fc7<-82ONM4QW+f6W-&UODIRfXCCLaefV=LC<N1+(T]^e)
3VI+JU/8TTIP:31@fZG[bS>3^2_CS\T:J8OB(OPYG[TZfb=H?2-RVMGD.YP?X=+]
0R4ZSJT26,JU.-JFCE2:UGcWKd)<R/3D@SYX\^GSRH=gT0Hf#=[XHV<UJ&Z:NW1&
PLU8P:DCaR,CPgIS4CURPKR-RgR0RG[:HNYDe-M]d/9H@c<Ra_:XSCTBLCH3SOFE
Nd8P^AY+>:SI(81ODXJLEbTJQ1]);4MR.G?+-0^/YVbV=LG0CL2Q2,F>7ggBI7I#
C[<Bf<W+??I7K;^0\X3DE#@(B2U#6;8AH^N,d5A=BB=Q<99A6SKLF7dQcS3<XXE#
Y,9fD?aT9.?_AObH0AC5B.L0(eWRO+YbQf2RQf,1T\H0[0e?5YFf15]T@?&C=FKZ
#<C&f:e&/W^&_8+7b53M6D#d]IY)P+G@1Q0aJ?;:1;L_?0VYM2]?5;JQF<\,-WLP
P_?U:F_SR#8J?1@D13Qd>0@#P\9PE(P5>^7/_a,.-;C^TA?NPHRN1BG1D=/GMZF[
6/QM-D)QV8IcX,Y<[B9-#5eWCM06.,]2/c>-R<7+T.S(f:N)gFPe6K3cL\Y40C?J
T(-\U<K(KHO+-cQ>&(:R2&3Y,=S6d<T6b]^,7,ef[RM-63RP@VCVfJa)0HKIMTS_
[T[L&]?3NPbJ)PZdFVMWcB.Lg>3W>G7FL_O\ZDdE,a#TIa#8(/[>aU[XDdPFfA(-
LX;4;2?TaG_gA.dOS.^&J1MG(P[.cOBV^]V2Y6VWI=>DSH47[9QNO-[,c[>N?=[;
b[F(Y=D5JY=Hd2)1O=9,bcPATU1C34c2.R_C04Y4c0KbgW_].HU@#G]Y:U(g)K6N
4UW#=B>>:]#M-YXa?D7JB9Z7A_=I>M0N[=BT:F^=I6#fG&>7QVD1U3-.OUR/4:..
eR^3aXE:OA#OZ==[b9KdQ@fD-d(^ZZR?ARB0P@d)VW5,Q>b=&LdBUUgBY)Ofc:&J
6S;R-+:+VBaadIJC0:A-JbE9g,)9/V>gZA@CHBSM<?B3]\-<KQ&/ZLUd:F>,R5J>
4=S&W+g_XG8NG(Z9a9G:F)>@77FMT<A?Vee.fQa8F@cG\_Z8&VfdF3[7T/#G6,DL
PRWfJR?U77ZEOTBP?Zb:g)JPG-20Fe\=dBB5>I9VIeS4ZC7YcVOKd,6-b-KB=654
_98eT?7.W).HE(-C\/DG\WR-Z1PeS+g-.IQC,WU)L[=BL^LdgL]])YbU2&S3A;82
B)c?AbaUO&3BIZR/?RFV:3KcP&WEZ;gccQ4XVVbS1M-O6U;D5RR/B_Q;<00)Fa_c
#5<17L\:^g5gTT<OQ]FaU@_R@_N>]5/?A);M4gC.Mg#f+cJ@Zc=B85-GG]6FUKb/
P68VTPEJeC#K_bN3<_bQ0a/c\OEQf&OQP3MVIP\F@19A.eNdZ;4H.D#B<X)/?L)S
&CDUeL3@9S3gDL,gB.Da6B:KfEa;PX67OJ=34-:[GI3/V;/-_CV]DOSQ@.J]T)W>
Oc56DKIQ2][?XY>e7E]XV;N@XJJ)V7(cE+UM69K.NPP&,[b((:-Q36d/e+MQT3MS
dIc:@7S-5Sb@R2]],N9E&cPf.(/@?9;2:GK(;W7AXA;F).VcZJBC7F_eIMUE?9Q_
HgLadBTQT<K,a/O@+SM&<K88_]5#Q&W7Ga7g4PQT\C>Mc911)X?9IXWS:dXQEV/#
C(MS0NNAae@,X?^CRVA,fd6\e79K(^,L7_2-1+^&-G:=#PD0I=gf7XT:S><A25T6
ITB0VF_Ub;CDLT#[^\_F/,\cGaH+7e[OLL+0&?eaE#.5OKG3N\Z(#e.&A>Z5e,b,
4ANPg.\6K8-;ZTDJF6@V&OX+^MW5Q87((KD^3J1MS]TT@TRD_<=6A@g9YFTAQGK)
R+dKg:XKTQ]]3ba];Ba2X,:XA#)GT?\];<d3P[4,1XYf>.W@&>e^a0A&eM(BA0,)
2B.R5<IG42(@B^HfOH-90W^\OYQ=SH<[-T/#?#90[;FV<bQbU)[NLGcZd@<5b,Z@
4W-N-gE^W=V6KLX>&DNH,\<5GcaVNRB+F/&H_VP9O.>B(Z037MaH(1_S4]M(>CS\
_TD6>IWg-&TFM<R),DJ/YC86K?DY[RX6,g81QB:-=QZc>09#;_R8Y1-/#g#L7EU[
P/7dM-R419RD3DKVDE/5aGX_D_).2NM_-L;(O&?:Fe?]F]+ccFT?KE71Q?9=f(@3
JJ&CPWZ3E^O8[2T\;(Z&=(9W^BJNPY36:W#I4IB8/+V/D?\Y-@dG4JDKO1K@7:VU
7^5KGb<R/BDQ9O,(_7G-Wc0]I=#+W_QgO2Z,SAG9)fS3N#Hg4@d1fT-NL+QV@?>Z
S/M<T2UGVP=bL@9U2Fc:g6:@077fUX@7(S0]<KcaDZ.OaNCV]HIO[4\>D5?g47#N
gX2P32TP0QD4<7+g/=YAUbG78R6ORQa\-cS,=JcIH)9,2AA^8(/H-0/@c053f:<O
H0QQ]aR6G6WL>(J[^>+6RDHFV0MV:+4X]FLgXFBX@f0G.DMBI0P>,J;?@NH[SN1#
6)II/6/5X9[IS4+fQY<X@V6=1=C@H?HM6[H[6)b+7d7(MWE.FaC\AP6(_fN4d7DB
VQV(]OVH2)P)<f@@LFNU62-HMS8@0BVX0bM:S:^7AYU_-R4XL;2-MW>)W)BfWKOg
0K.]DH\M^N1]UYf9dgX>ENZ)]&<d\O5LLO:8HQQ39?.DQ^13>0)O;:Z8c_?+BX_-
O+#;McgbISQS]>bJ2SLbRQC2,08XLLfQ(Pg43PT[9K6/Z/SSf@XXLADJPL8]cge:
FG21G]_J@JO4B?bOSL69GH2Y#PA^=L0),+?H\LdH+R=Y#\VCF9K0#TIbK,.E]]L9
gYe<:;1),=cPf5VUNeI,e&2X#)(5.0L,Bdcd39O4_U8f)a,#TRX\Ua=/TKEU++Hc
V4dR_HF9[7b=9^@X&;.<X@HcR37Y8\#X0)P9G=UOfX98[AX?[>,NVXY7fNaP]e_V
I4:5DC9S@/@8<D)^8_dXM;g#2N:+;,daDDB\9?Tc>?)-I-1d9E[FcfVcQ4.[BI)-
NR+(6Y7&#85R-Dfe7ZAG^NMeL?>Z4?L-Y13]>5P^LYF^aO5KRCFX2^7IOTM)KPPN
3CU+_PaK-=b.-,Lc\_Qe6\SY7QZNN>RS@OJPFB7HAZ+N>\YINF^7=@+KU64,7MXG
:VM<]8eVUe6\Y5YSEM:UF]MbEJOJP(KK_)(ea<5Xb?8Rf874_/_BK7UCeP/&<H+g
.FSSDfEP0A:KbAC)^[VAQ1g4>g\1H^.<S01;V8a+^?383U-L2Z;aegZNH=)?H1>X
;>@=-b,SUW3PX3N0(@6XF0fKUO0M-PBH&TN@\Y92)ZX)3aVcFH#[-EI,cK/:N(24
N.@-f[WFRMS.4__^U3+G?L9]<E7CCe87BJO&&#faDVQ2]KQJ;8O:<87-X^Sa84ZS
CaY:684AWcTE(A[KBCOW9Ve-Jd4<B4W5S:KPa99WV8=Q97@0C+)cVUP\+F8B@bDX
27>56@aH;e^eU]0G0?)>N2L712\3LXP^6dAfV0HM.X&U6D(,c.VC^]cGf_JS/Z/+
:;9JNgL/Y?,<gALCXFU=:FP+gb;/G5.USAT/dVFc]R[Ua-0AFQP-;_DMD;34gPJP
URINYS6S23eP),/4GJ?)AEZOUb)YdRAB;:DP;7;4\PP[Q2Mc7gPA#\Lc&bR]+K/N
?J-/.]_PEb5\d0IcNPX9c--+FK2I6SS=eU7IV)M.1XgA1+UBQUL]F=fO3720eRTe
F-&J#I#W&+.A[1)HFZ7QI,Y4cK^e@(ID&Le@MGPS3)XEPZ,cOUD)A&HAQL.\D_0b
6#[@>DQg[We8T7EB-/4K52E7P=WS@4Q9LKE2PI)CTT8a(DGCUb,dAab@>GdJQW=D
=^MgaP&5:d&>WG7JAP[L(EZQ:e3YXb7#a&AMJcEMV^ZUQcc^<;05(TA[;.18,3cL
9OS.9X88bIDc2IKRDV:a#C]g;LC778BT>J_c.X[B:(QUfV<-9)-eZ\A.)7=P?3<R
IeBg=C[JGF1f7be^M4L-QO+TSG;(42T/6cVTe#PKK0<D,;:L8ZHQ/fTA\Z^GQgK.
a69&@VO+Q83fgV86g+@Z+91+NXT<VY,WfSM693;1@48fKDf_E&YW&A8)PI_KXd)f
?,[PR7CQZ(;<@XMM5A_KYD4BA:(5f_GgTe46+KdMSMf>8W,N4SSVT-9Q)8Ubgf#D
DMZdUFOOd74=:Y)+:DN?KdMX@@X)_5-^=(_FZA5,Y?+.Y<FX-]6SJP7INJUEb\c<
W?6^0UY::<P\A;&V6TIaMR:Y@9Jd7^/W</4VTT-L4Zd+H>/[Gf0DM#Fe/YZ>EgIJ
JNK:[4c2P\FP(SH@N-=V8deR?_5ZUTVJE/b=a/:gM4gUOfFD,I]K<)((2XbVE73]
-1LE=.,8@SbT(N<0FCLVPS9X=?cQMUTQ&C))H4Mc@4@S&e(_E^,.HEFVZ4-?<8?b
^7RQFF,[P1M58[FMRR[FY7C/9A^W_C6\>Y,L,B>b]eI7;&(H_BCU)\HdTJ7WbQ\_
A;NL3CP[7C7(_dD+X:-#QT8[6FBSb_P@RQXg63#P;g6QF3P1G42-bH),e++dJ#^C
N.6L>O<N:6>T4W8Q<Z0CFSfA+,V/LS2E.;B(HQY[F17OK3>U-7GMJYL-@f5TS,90
92f6Jg@f9/DLI/d9C97>fPNE8SIL))ABW@DAKBU(#DK2E.:AHKNB(=GMGMNRIGFH
UN[#79_]]B>S+UJR+L-12VB)=_3],d(CKUd=J0dBf-3]#42R(FO2E6G8cAB]L[gI
d7FOV@a0/H_MV.#0]XG&eBWDO<>34=\_AP6,L1OY:0=64d]H?cW\):.aH0/1BaO_
>FUQP#M,7,OVWGE&J4cV\(c[A^4VNO3M\)5[0T^YF6:_0\J[PAV74)/L@DGCP37/
fYU+8NVaDQBd?WLQ2NJKMMWA1)d6E@9[V93^8W+gO@=Ded9]?9@=KEIagHFXT>]#
GPKQA8B44;0f?7+V-_Sb<fTAZdY8DbBe+PYag?&Ya[41Y4G>+&:/4EXB=gLcGgCI
[L7c[AK-@R8I;WTL3eI^R5T6Ub[T#&-gN4;-C+C:MTR]H-HaO([-2L;WN[)f\?:4
=-2M?TaXNT#7EG80c;d22/Dab@WZ>6IVEC2K17FEOaOY?3^-54D4Ye7/5>,)<Wd6
<YaA^2==SRD[c1MdI4bY71^(KZZf1W]\,PWD(/5XG3&(4dD:=aO4N0dQ2N]QOSZB
?MF=<+#T?\33<[7,W\cQ+Y7/:X>_XGZ\ff,JTVX+JXV@R7A]Xe6Q(fZ=M+WHL(dB
\;F47_7C9;@M0]YE(TS]@Y:&,N@U(Y/aaH=QA7cP;THcd2/Z8O<Q:O5\T8/@YVd0
Bgad7][aeHKLQ?YKcXbdU\_OC2+T?2_a2C07JO]_^dBB[T)M21OWR^B0ea6Y_IP@
?YS?+J(&F5J&7E?OJP:N.-B#a4UJN)0@fafZN2&OIOBZe5H#b3RK2)L)PBW=K,5J
TQ2^H6,;e4B)AGX6bS8F#<7&LSa7H2c7ERab#]9cVW[e^-)ME[VB)O7/;=4WM+]E
LF:3gbX@3D+FaO9KC:ZTL6A[gEV,.UBWC,TWf<0a4ScBPJZW?OZNbNDH6[&0Nb9Y
E\G-A27Le5D0.gW;2H)Ce/&L&aLbH/\R_B,_)9+TdV6-/JaEN@a=2Q<]cP98>K6&
/9gBA@Xb?&I#>4A]\BY,8<#CLE1:6KUe)+g-?,359C@bI7&Pe8BagMbW6ODe9=Q(
/C90@NfM88]T1:11UN1&=KO?QSD@(3@/9:KdSCIM>)T:bGBT?2a?N;<ae\TdY+30
[0FAWYXOHdGALeQC2d[afB5G)==>-\,TD858/==78??+L4I2Pf[E4MF>-<PIL/C>
_@9b3XQ-@S9\XPE6A#?Q#]Y2+B8G2=>7)ZL(FKZJN&Ug9D5e/9,^WVS;fAJ2F[bL
BAF.X]?4F8LU[XS^)a1+6D3/XQI/03/<O8\SJ9\.g]&>Q4e8[Ke(D.YLJ.5gJ09@
SWYJ)=e4L+d4GVZ9EPUV:If;AD2@>C->@QT?E8ZHaI(dB;HA4fQ]b[I<Sf_F)O-2
,/9=Id0MacTK)7KW>>Q&Q^,)(/T#9M/.a0[d4WA5.GV52-_US4We9T&8363[SMfE
7N4KQ5E,^:FU?6ZEY]fc7Kcg3^3HPK[YBa0^1U-[_YQY,+#@R?26=-)8b[8\4e1U
OR-HR5(1-KS\cL0@bZ&<W=-eD/WJS,0Qe:b9#]JV-1&\d10&d0ga_9+_BR(Z5<D]
@g=ed4A+EMT]S3deWH3?QAKG_DP40#UC>I[B-R9K#+3HQVE@QcZP]9]1FWdHfAc]
(da54DHg>8TR/7I\SeXag\,;QW_d)Y@<&SL@gXS/XP@;@3A:?V4,1)Ob-BQQD<;G
W=C1+2D<c1Y77e.#SIN42+LR,b]GDX;IMT[bIUH9DP]^^Za(U3[+3[6D?48,N&,\
>HSKWN_-OX+P;6SCI>925CAE:cObg1CAf0YRZ-K#2ee1U;D6^e(>Icae;K?;0P7>
]@6MC?\VZ1cX==TV4<8:?f(+La]cS?D]L9B9/A-T16GCCN=36Ke]c?QOg9_>;T-@
/:6#?,)(34CCVX,fDJ6<c)X7-dM>7ZK[a/,TWMQd4IZ#)Ib0aL:?cWWR0:(#QXS>
4H(X3^e34GUCW&7=4I#IcOC^&P9g=+;_g_,512KH)B<,L_f0=B\T(d11LF34eVU;
Z8eGNWI5^;#D[35d,S#IQ<\]C(),dfZ,Z#b<G]]);d?[<FNREdA6#OOeZ;3+(AGC
;WHaANSVXe2Y5&)M_-7+FB^?2a=UHKJf8IJb51e=39=&]>3C9IV&cQ=P0P<C?U_b
RdXKgY/1\LZ?(5ZGT6__83G=DV9ePAaF.(:D:3:W-e>P>XaSP6>VXOLbCB@EH@?@
FKFC-U5cZ2BTXA(f-cP286VHPZ]K/<#:W#aEE,519MD(bNVe?[6f);^<HTT\_S>F
_?V6cC:1Ca?>=X)^A]-D\.N<gI?W9]94J(3\QA&D4gW-J8^)\)bPEWJV@XI3^ZD?
A8NV6X14U-W=TW17fYE-e.-MGRHITW_9P/Y?,e^3N<83QI.K_UHd(BKGDdbI>Mgf
<B\#-U;-KHcN_[4b5KNK>FQ1\I1Xd/R#SJJHf3/1;;U9UT7P67MC9(W?=O::GJ#a
5,4[+1L2,&e15:6OJ8\1[PaH[]5Pac?Z.dZ,E)I0UL#8I7F#<7AX7:.2c6I:R]/<
A&?&Rb]<<HR0ISPBLVO=(V0+acQfLFV^^W2QNW(\M&NR0LT+-_>YYMN3A[cDcP5d
MdB[AXJ7#=>Q7.b\20U]C6@HMEYcYN]\eGJC6E;L_c3/-FII::=Nb4H#>=N;-8#?
#Od<D(M(T3LT.G>>2E,DSHS0<+93\>5<.[;HVW1DK8eN9OH:;]65O^?gc2@3aXY?
QVANTK_OeB:TKE9IEcT?1:S<E.fJg>g6@\LM>Q9W\T,M\>QM[Z9:]<C8W(E/E+SZ
KT6FX<e5\YZMD:VaT7(O9MQDBeb.D?MJ[-.AL2T9C&I?96,T>P^#_0MR(Pc3O5I<
D)T-C^>P.d=,FOS3E?La>dR3RCCO93V)/?=4/=NC)<YPJ=cP_2g@)A75<1-/Q>>M
R^WGS.^Ud,BNKM#,J5S_09db@P+WN]3gXGb&\f+c=9<)(MJ[6T.3E0?<&2/0d@/a
/@<2ga8U.baSdIX_^d1X5d,?:588LW^57GaaM&8fY-4YTc-4e)3D:/7fM:1LLERP
JQO-FgK73+g=N.6I^:g-\@O3-+,C)^PC[[^;^^D0IH7(#UK9OM>Y.fTU7-4S0WU(
EJKXecI/(Rg:R>ee0A#IKNP35>+,>TJ;YN,eT1.bT>QSg2KOPN?EYX3T:dGC<b<?
YXDV7VJWc-(Hf_^\aRM3Ib,N4XAeZD5WVRb<<B;GffD79Lc27-(1d8UcN1N_fc=2
+^J8;)fK26@N6]8#[[#6ND))E6>9S;bAR__f2ND&X+Yc<X_8&7ZV+#I^)6#84&YS
TJ#Z(SXeCbLfJ?_dPG^4LaKV8U+8efL6GV[-;I-(..N#LI.K\RV]]^2W=00\W5=b
Ae;a<d.g9A8a\VdNZ>5R;,cagY_4bDN,6b,CeDN0M6]3EE2EY^0NZJB::E@@.FF5
C6A&3@JW#ZBeF<TB#4FK5_,-\GUJ#/f?#V4A9J+UGHXCG\;DFU\3GZcX+g/FGM07
Z;/:344_O0KNV#F3)fE:;SE13/f:Q[AD0f4WNFBN_N5:V>_,WE4KWNJMTFLX[ZRe
<cW<BZK?(KfE5A]Od59UBTT@LVU\U^M7GOJg&;D&-LC,Dc8,IcO7\SU@Yb\.SJfH
A&.V3e;T>e,\LX3V,)ZD6KL4(3,[/YC,RJJ6VE>UW(Q#<D@D-+_7HaV8-DB=b&P5
W92A@fbYA5Fb-<7Q->6?(g.F<3;=Pe7U<XVdd\Y2[eYT1BS3S<O4fRQ??#QPc&?D
@UcVN2)J(7\XH/CR^:;BO:9#6=b<cZP^;9-/bZc;CJeEWK3eg8\U5V:QYG2WP3P7
<SXgZ6\XV:ISM^_eT[5>b56VQY)@+B79UA<](6cCa5B4FO-6(Y9WSV[(^:92JfEG
&3<Z=A3R#dSN749]O>,\JE(@BHACdQ=BPU=,K[<>fE62.X)OWG3+a8;S>2(A&&N]
dA,;,7Q9F;5SaMd5(<g:B;4(00bJH)GMf52.SVMVb\RP\Q@b(1YR29IHDG>FRCa(
S=UX4c_3>P)_de&G_.AK&-K-aHZ_?BfWXbTU85dD4Z+4J<MU?T+][+d[9VN@A1DH
#Z1K^L,W3:d^XTS4C,\R)1OB<YfW[2?TaP6eNKZQ,e>ZSL@X^f7aP35R5+=Y1.V9
ZVeLOT+@3_DGb]\0c::B=a<N@ZS_UV#AZY#&S3Q&(Wa2BLM>c+#^5#6TTBC+c@3B
N-bS>@CC(Gf/fE696N\8@:1cfDK4#f4R\8/]BR/\RL=eHCZ_R.H.MEY_V-;9Z=7P
]?O4>-?^Nf2US=70=U)/2#B&?ND<N&)F^Q.Z(6PL&>)I@1KBFN-)GYOgb^A5YC+2
BH:[ZBN-7>,aQ\M^G;X2?648KFe.(\f5(3,GZ2I]e5g>K^EI+]R^A-FI&?A\JfYB
Q:IAW;;MR8K7&e7@>K>]O050Na<QEB2:YL5L:<ZCIT,6<M),G:OQP\;WM/QCL)0Q
\IgQ85SZXe]/:1J05O:_-ggL@YSN38C#1BG?053GC>S=)C:[YVMOD>[L8G+ebgMT
=U02eTJ,fU\(A9Uf[=.8HK/73P>WBQBY#WM8^)S6B_()].4b],Rb#OC^55YQg)6J
OTJe8,.8:X3L[SJAZOTb+<dL=L:H41E-g/cM.>9^Kdf^P(c<5_bPg^WS8)#UBYN,
O.Q8-K=P9KA1T.(00\I4IK4?[N]cc8fC[eCF^7M3<9NUJ+b,7P(+:^()?<M\e4PR
5J(2/M[MQ0ZIfU[BIZe@aW8]<agWH/cE^YXAM:6IWMI^f>2FH@ZU^#V5K\O9-/ED
+@=aIe:_CI42.GGO;:<MgU/d&Q1;J;\,5:JO57,+FSMXFTg9Q;_/2DJgLSZ_d4(?
;&_G(\@H>C.,V&Ef@B7Hc.04OcDQ9VPS)DcBIa?Kb[@56>0IFT)/AbUd.Ha8gOK9
0(ddFF6A=]KEe;;?&g2\a3]Q_U&OI>PVI]I;\1/XB7IF^a4[UD7]f=SN7HE6eR@\
>K8OM926WIgFcG3X=3cQ&eB5RX4?0@a[>J27([C,Md^Wg9Wb<?DAQe:V[1]IUYK-
NN/gg[:dTV^P]B23]J(L:2VIVI;V+596G\1bL8+H\J,@^D2J&a96aZ,OL(\>KAK;
,(\55B=#>T>g1g2HY0:H2N.1)3O:?CTTW=Ye(3@2N7G6GP^MO\PHeBXY5PMAWJ8c
ceVDT>PJ5DU/QB-XNDDI&95V?\?Z8;e#IC\a;39G=20TK?5VT<<@9JPSfecOf)Q(
JXWG5bcgR42bc@.cU@S/\Y>f3ITG6RVT/N,N=e5D[QD7=14OKH2^aE(?+OC[@>[^
#L/8:ZO,.9b7I-J=QKY][c<:7V6]I&+L0=S/(b8_QfTKT\^84[P#aV17:E6+b6KP
7T:]0;YI7C-dQ>?ITg+&Mc<W;R47;QE/.PaI)NWF]7cOUe+=E=\cZ.e?QX[KZBQD
]<[fBN)]6e3^N=DTB-[TD=@4-\B2#IASgbADR2PFP59eV(J>KT3VKNXVKW:5g#/+
>f3)U.cDY(7#1^UH5]YN+e#NN5&U88?G4Z:LBQ+9O>+\a0]1KIE#3d8UUaPDRV=#
O+1Y1,fD1;\W991/,B\<[++2X)BXL2#e91V0_NKeH9E8#RKZMJC:W+DFM:>X9B=F
^.3SH>+L-CS8;7+?V<^,5;)GZ:)#S^:6g^&c5(514(JEU0KW:c0[>;FOMR&+X-/T
&7&GY<HZR;9N4ZU7#E7<RB?a[OcX:BNMdV^gb7bG2)D0BIYD=>/:g-QKaVLS2eSa
>0D:42UdYb+\L=VcWH]\09ZdYEY.?;DL)PWP=SgVK,XgIUd<=]:cI3Q51/a<4IQG
QPa.B7>XYV9Y5=A\7-A](_,Oe2K?e?/<W2]-;7)O]O??U&1;;eZ<N/0.RRMg4aEc
(/].NVGIAJg4<MID9P79_X3I1R6QA0DdE,XSV\LNM3D+-03\J263TO:[c5.1-Q;W
_CZDcV9T>M[E>V4/dN2dUJ?))<UJG#VJgF.=fGQc2FR3+<<>Rg)3b&g5?If4P?WE
EI7K29fd:BH4@dZ-0e6NU(Q,U:E0A.2G:EKP9/3d)Gd=5)E:+,aF&(7.ga6RN=@Q
,0:2R6QTW#3D48I^5=-;WSe9D,d.&H>1;PCLZ?^IUAAY/P2((W,^F,>D]-g[g_;.
O(I0O7&G3R_Cf(LW0FUa:P,HWQ)gK\]GPGfX]-JJ1;F;dBO)S?T[b<=4g^1LU+I@
SVNS>Q6SU<0&:X#=)0g3M#&G9GP49:Ag36RCfg4aG_C--VF;^A6b1L+BUISFUA?6
S-HQVX&.GNQX1c<#=93#>U3@5[.bX8P+OTX.NI#dPK=6TY,aa[6A1K)/Mdfb=EVG
Nf6IcIGTW(C9=&M,FZOZS+ZN>Y05=70?FT7N\RO[[&d&A4e58f96H^XM1/]]0G_]
W9de[3)^/?MB4YW#A1O+GQF5cMHI>JbQ_Q87(>K8-c.=6bN)GHf^J#TG;#F[Y>I+
>V?UW\8M?bF-,L/#/8a<P.cR4S[?BAFd9GL+5XEf(01J+J<.LZ@bA30eM#f-?)<V
.QdIO//Y+fH:g/AOIV0[4)K>WBJ++/1V8X9^#V1SO94Q/:5RJ.1QUKT[Z+E5aM[c
XT.cRYOFPN(-S#?\T0]45fEJ\M]NC@7YJc=TT5:PeO+&\21M8BGc:(Sc:P9<^#UZ
9.=J[0_4TIDK^\JFE;4V\3f.N;;KbAV.3NKQJF#N(GgH-X?eSR&Q-E]/WbdOKF:\
L9//)8JP)HP][Z2:bSgHP=d.Oc]gCMMb5SEBXcdZ59-GZ:]J=+@4G)Q8eA9/=&P?
3B/34)6QTKBCHTH7Y;(XaXW\g8H4E;_#e#?\<9?f7A)fE\RfYG3:R5T:2P)fK+Xb
K?3MS#AM_Z14578X?LC)0UW>/eMU4#SKK4S[RScQe?&HD1<MLWgP50]4<_f,8L[]
J>9#1Ac.-PQ[Z-F4(T5^,1P,P9ad?@e\U(#I.e<5UbbGCfQG/[O^F&I&faHGA9LP
<7HF6>P=E1d63.VcHTX@VP]Zb@e&#<#LQVaX,U2YGO_L8C26I+H91U32Eb]P?e>P
@:B-]T.^XdAP\@S)YLK9<L^Z5?6>?faJEeA?BX+W@+F5Gg)\)8.TLc<a.+[\2,e4
Z^Lf<RdM&(MV;Q39R^Ma7@5&-c713D;Ccg(VZ,7,S_QY1-E<Z7OREJ\SY-b/bC,d
b>HPYEFdDNe)YII>.^dD?SLVXdfK8S_\ZeFIHYcd=A_b+TD=#:Ra?1T)<V=@?9fU
#?6\eZI\.EZg6+C<N>,UW\f?g5gTFIcUBFbY@&:g917L[IOJ;/]L#?6^IIAS@Mc+
R3.?AU(1N]^g_-B;0-\S\/gIT+(Q:QSAZ=c8N8;K.I#?1e0=?HT:6XOC2b>AXCJK
AMFRB)dTAGPL4Xf2DGVg<4?QVG9/\F_&E1+?K,QM&M@@7@&>[IXgMTEU?CZKE+aT
,2=,M:S8Za[ZHYHBdBZOC7-C41FbWb3;0Sg.I3FFS\JaEUYL0Z>Lg01UJ5@85<5=
T9eN:8aT7[B&EHW<Hfb8B.>[0BOV=g]DP7#2O1)CLe5@Y64TA\LS0[:5J#\BA<.[
TbC;3/L91:OTHPf<:bE^\)?>JD5fDF08KaHD-QQK,)0Y8IM])gT\0=A4J?)U;J=e
VPF8R1f(9&GgJY-(@<:QQ8U<+Xef.A)[P3[b6<9@XB\XNN(A5LTJ&dIRQ+J7]])0
X5O27?MY?TL?WQ-F+]O]c.dggg??PQ>]S\_E&Yd7UfNH9-a._fbKJ)Zf9C[eTA/E
^^?+;G&WB=_...KY,A=GBaaB[6>0M@:^EKBPQCeGPA?aJ&@BMA(D]BZ.a;HP^XAU
MX7XH=[P_K1>7Q<PMN+(5=c3]?eVDa+08AEQUDSM(&&094.KRT:ALP1Q2=c,UE)b
CAd7Z\L4#G(YQF4OVN\a47JO+a2AI47V>)RCUFRb/KYcNV^5SJPdKXJXeBeV3C#)
Ce0X[]MM_R8V^<0,H#]QSCZ6;J=;CL088GKWT;9ZO^P5eb>9_-K/^)b13XA)SK-T
B6CFB?_IV^4M+SXJ\U065f/)_F1:W-#d+<e6c9TeE[>ge=?5M0RDEKZ+Oa-/-D^<
\57#eHZc(J.3@4&1c_KE5FUZ,]06aPdY9#_6X@=(W3Ef(3#OB8<1fL),GWTK,A9H
.=Xd=R6dY2@0@bPLFK^eLYEB8#H+O#,1T9J]B6]b]]AN4I_S/&/_]Qg+V0;AH^d1
fdY/+2:OT>6>d1&:2=;=ZI<32_MVYc0a(.dANDd&K;>C^]4-QT=ENCB6I@_>WW19
=38f:fG.B3T3DdA3HX?bBLJ+b7gV[c5@a5]Bg1^<B=N5dB<a-;(#SW)#4AaS<a1=
48C;8[EYG@4LV:HFM63V>_E,=F1@Y-[a-52cFA,[5MV6N6IQPQ<G_C[],6XTA=f]
g0]I\H4a-)AG<-FRGB^@NR<8^CTSd7\GBa9(B6If-)9-cXYRc&?0TD?)TZ[M_Z?2
@S&bIfdXF:^-QU(GcW9^/,&SgDd[b],;=V#L8a?cDO6;D^C]C&_MS>?)fL>R62BW
(UMCa)+>NN+WA=_HRF99K7-QcfR7DT/5-cDTfe0B<D5]dcPZ?UZf+.)-=P:KB)C=
fLbXG6#=g]U?R;M+Kb=#fN#d\eY>e?6=X@;g+)/.dU.Nd[EBPT0ZBI_R+D^Kf(Z^
JHLJH8?aNXH]Y2JbU2N_\\QT+M9O-QZe>W214FEARO1eHELL\AP>8A_;dDOdUWNZ
Y..1MM#([CT1=?L9M8PHJRQWJ/0[?L2Ge9defdOS?Y-5DVSU,STa_P#b/:+I<2N^
gSZ6QDT&UYS0+5bQ0GcMK??7gg)#AE.+M-,2[^0:AXMT,QdNceJSI/XYYfZ_JaUa
^E4a,PC1Y;M(^f].9,D_I>#BQ.0A@EEU<YT^>OGY/\P;P_8\X9H?X>8eg,VY#FG?
@I#(C9BaBI5^c3_cg5gQ_X)c9aQ5V+T-(EI8#b\\\(>]EN[[9//>;H80ETeP;11N
.-JSLR81Q4YJ4B\S\[PCQ>,&-aX>K,9f&G#?K0&AaE-3FW_T;gT?O@0a=PP.d(dM
[e)59J[[a#J8F.+^PS4d0#HKY-=aZ_Z-[T2L]c2DYBLDIDCdAJBa_Z&^5AD-,3-0
ULJZFM\6cCc=<,?X<b->SO(,]SU#3/1FCM#K1Lg_XAc8Q3;L?dWa2ZQL,6H:8@4E
aH<DVVd=#7U]/fgTBWG&+;K(;c5/\[4814E]VHMW>]2BZCcV\>(FF6be\^e8f.8b
AS[,6f5#d0CaS)Y=ITdXCA#edBeRVHW]F/\HQ.d\G?[+QPY-6.4OP/+dX5:;]]]\
d62LKg<fG0^Z3_\)[><e@.W(JeZZSG&9WR)d&f]8#5OF++23g&cg#OT+L^9PbVV-
P8^/(dW=?B4a&CF#L)G:fF_6LOE=VA;]_aUYME11SWcTBT?7GV]TD)M[?Q(+(H24
,R<Y_O]^_(M/<K&[^3NBLCZg]AL04d4dddMY@Q4+SG31\\L+4TJ@)a>PC(I_bHL^
0/C/TP[6V#8e+.^XUe5B:^H=?-f6WI+C6U[c).[gB8Z;067:=S)CTJ-g+8K14?B@
VI/:1R)GPEWP+K2PM@Y>1HBW&QL;Nb5A:1D3SP#[Y44QXQG3GEBJUF3ZJbY+\S#\
D>H/<L(2Vc;Ue:92.ac#8\)c[1GJ:MI[JJUQQHX-O,1<&J1dIS\]0?BdSL<?RI/V
Z1>GHJGT8fQK;UM<=GQcQaeSFV3TS9ZF)_61QD&?+L_C)Q2&=LU#U6G2d#A-D3U=
gRSKBOg>TYBb1;7.V#.9MU@K;[1ad(CR<[.^-e<d#DY?D.8gV@EY(8_FLZ?-EBb,
]fdSK+8TYD1e>JX]eL8-bQ:CY8].@IF_BVe)g]f+(]QQ5eXbN,NMab5++^Y/J\@M
eGNM.aR,b@8P>2UYT2.(gd4DdQE):Z=IaaOKXK:=g(JGcLW<CZQfSV)HEd52,<7C
CPLAF,dC[_58(_VYE[65G;e4\DHD;L(\[HC9b:]/3EC_3RFTdKJE=/KJ.ReQ8:.F
:HJW7.G)JF7RMN]&AbF33[BC[@:VVJfODHBO>S/AAcBJ_c9BWK_UgT5#BHN4EF^J
-BD-G;8)#aH.Fae-e9cD7IU)IRI\X1.>DNU9bF2<gQ65.6X:PF^;<UGad=d>C^C_
;e5Mc5Xf@FGG>XIFH^+bS[=+,,RJ:E3W/TE.A2?ZL8E[+NC[\]L4I69@F5PY[Z[D
T[,I#MV:KI(4M)39Ne.4+K:<@.D(b6D,=X?SH>/YK-)S-,_]P0FHS@+N#MA+&eEg
VOK(,71LXAOF>BJB^0?#BW7Z5-\g/0T,.9ge=Y[N^2WQKPR-WCYEH@e>He[V;99?
VX88L\2IKEVM6OF#^fWSbPV.Y)^Kb2[Pe)cg(V4K6\M8J4<TM-2KgI<?[G0?QU8<
<e[\TUV:O\##-@.?).[BU(K@U1a#4e,FE_=R_,.A^F;[((D5.^gGM2b^JfGM+KLg
[I/[([+gEUMB6#6HPB.>V#<&D+DeFX0N.^8a.SX94SX\(X-T-YW+8C;QQI6&Z9La
G#MN2+V:+-SEGTI]VL4A[(EZ0CbaH[YPd[LG<Gg^?@/33Ka^]OG[8\H4RFcg]\F_
/WXS6-4ZJ=EC#UXM^,^XAg[K:[@_LMc-_.BWU_]P+T2QL1@N]E0:MR@@>4^(b2MN
^:E1B[efe<bC^7UX)F(M8009bY4^083Ve.=-H:7VN@_#9>.#0UOYI(ca:VeZ9[PE
SfRFWM[0P3);W7fee41DZ<413>D_Q,N)E0?S#I\.HZ:7+&?#_?6TUE5N63[M/,H:
^P0<7Lb?-IDK1/U#39GR5N>.VfIY+:1@=@^1I?2]Z3;?GSJ3e0-</3#64/E/f[/I
3)YJ13XXQ=[1=a(M;5\]fEY(@B2eWK-+G9eW_3Df^<U_6Nfba&(:;)9+QOU16.;;
F2ICN;R5A[G.C#.I<CF1J5YQ7-a\3/<,8]UKXXMMS4F>M?#=GL.B=BgZb[(,g#HD
FR,E2PS2gTb&DQ5N.Y-1ad5OZL+GA+=HXe96T5>&F5M0/c<Bd1.>gSE+7#OcL^Yb
5Eb+Uf)-=M5>dJM3E4NN:g8Ee<TIL7b?aXCL],TZ^>M<.1PXNbec?8fLZ=bT:M7J
KCbY_U[GY=5<4c(SWKGZ\f=Q50UJ]2fS#@LO@JND]=U]A#c2R=Xd08+U_?c3C^R;
;E0^V10Y/O:_:e\23#V[\,BKA^=_73af[>67=#0K4@b^@gCY406IF:N?:1Z+#c/C
3UGa6(,aVMa@^K[WgJD:STFT>CBcE;25]&7NIN:&e[Ta1Pe3^6_V:W11(L88e6-6
Z?;AUU#=+b7HA<;QXGZ)g)JFUW?<d3K_CT=DSNW4@L355B/#<C?:87e#-SBOCTcG
WK#_S)DQR^_YFVJ^1<L>&C[T?]CGS03YJ:g8B,8M@e+=\L^4\\\)O:]BZF)8VNQB
aK@4]:QM@_?6g#WHccSL3E00Ka?dREA]FdT+,NR)Ta=;Y5,YD[_<F)5>-f/\T8)f
8:V:b4O\.8E&3_4^aNCJN/0>1)+4aeEL)2PSf+8E]KQ=b33,0cVZePYXNQ/<<K&5
&O;T@3aWX1\PUTL)QT:58dTX[P&.YC.)25B:a@P,^3,gPeCLd>cD/U2(QP@#1BOc
9_=:6.6c:MB1N+UPX[Uc<&(IL\deQV@S:-dKbY9+4dX=G9fA9U+(MaaHD8K,&L1K
bFG]gXEV;I6N-+BQZ3G&XA)@<R?9EUZSg85KWdEXI)QE@:9UDBV=M@Q>EP_/<(RT
E^PI[MUHgA1@.5)X1(/YO]^0F?V)]8F783K>N?OdQedA]6:c.D0+&\Q]<+M-;&^(
^=W+]49bN7Y0B\<QcdedXfSM.W9aMYd(+2Xf<>,C5]-:=X]4=Q^L@INfU+C].9SP
A1BJSO2B#:1&I]FL^;HILQ.e]R7fN8\;LAeeI].4eI&F^[0W1P7(/g923g:f\KVZ
L>V[464CEN[CODTRBZV>23BaXR(g<BT^8-1D_/_C>N8C(CKcgUcd\QF=#T<:>FAZ
:X>QP.RCNZT)0b/^PEP82+)-bdXE48eZU1DTM]E;P9.e06WAKf^A+TZ0MG7V?SPS
GEEK:Fd3&5E)___(.,aE69aK-(K)L\Wf3<<(QBF:e)aNc)dH[)@GC;=1T^#I5GYG
FND@HSB02EL/4E3V98J8\G\3O)L/W^b2K(C:B<A+Q\B9L,+(2W;#,Le14U;D]P:4
84/3(P6(XVNIPG8@26JDM+PBC-c5NQB,RUa5N?(H701/Xa/Q]0?&Y-A^)+8]JH1@
F[/LQ)MSAF<ZD-9b5GITN,MWISA9VYZ(<]O]&YQP:W.(3I+OE4?abQFF7>_9fR0[
E&N:bI0B:G\/BDfeFG9B>G8Z\@U^L#:N92]Ng8B6]A^0OX5?_U^9I\[\7A<-d8TL
=VB5GU_;HP,g8T8/T=bHGR/\RI#&Z,+ELY@>Oab0WD=#R:\Q58LBdB&#ed>&??5O
5.M6.HOZH[N3^(+3,M9;:M?G7@)81Ag?^bJD_I_3&Y7RWfNe91-Y,3dT17b4?M)+
S&@X=B?OLfY2AP2EFTQUQZP+255]AJ+:g41aF&ER-)T#7Lg>[URS[TPbL=7dS+49
V>g1CfbYR0E[;\XE,MV(^WPB,:A\-g/-TTb+(HL&EU42ANf7T0FJIWgHEO#bU1QS
YZZ1Y#6;L@N/U:g<)XdM;E9/D8eM&O+V[beH3Pf[3K4+O_-PD1?X\,Z(eA@P:68/
7+#UH[<^Nf=9N=DGNF:^T5#26RX8L(-O3RIGCQD.22NZJ<f^T?93KN@c(.F_.Ae]
Q&U:#c/fL2BMB9;A)&&e3[@N.CDT?3WN7QZ^3R\cJCgZJ,D(UM:9_NJ>>_W#K1/9
?;OR<98([+;G7P];Q2D;\@9QC9JAbD<C(b[B[O&N\a^J(HM8G>P,aVO2cO4S^2P&
=(5L#4&&)UH.WX,)#T#Id-96H<b:a&===DaW-SHM#Pg@^B+ZRU]U:S0P4.SO:9BQ
X]b51)=U@)UW?\_O3WJg6A\8Q=IN)_#5^g24+cB[CRAS#\B//D;T]Y=PK)<Af,>;
G.VaZGcOZXLgC1>+J/SZ>Da:BOS4cGIA>=(S_Y+XgS5SaPS#B6<9LGg4;902NZga
_[=P@F3.GgOY?3A#G1L0CJVEP.^5/><)MC\DIF5Ia[;;.,UZ@4LDSf_6=Q2OABI-
^Bc?g[G48dS?(0ALYX,4Oe8VVe)V[XQJG=JE5JWH@6?TM-L/7d^)QLCUFNR6WeHU
ZbT:]@F&)gJLJXBV/V6cfX?O\RJe:PDH&g&68IYUCB62..3)gEGPAB<4N.4g;RG(
X=@.QaW9.SRCHC#^=]XAfI7/YUD=.3Q;8H>ZX)KXPWZT3X/UbaGc:BY<IWS-]E)9
T:,d^+=LSL&O_AIC]d.V.g>\5>5O<b?\?6B@U,.\,8>cJCK+]/b0/bP6&(ZXf)8\
IX1FSf^<.SI)P,gMQ#LFbf1a\^XE(+HWf,D>W?3BO?]NO7a.S[/632W:XYY]a:K<
bR4ZF.:X-W02\b=0IO9g9?4H+Q)^DMe\EK0^6_:_3N#,KH>+F:GM?@MSa_I(=fKU
4O;/BE[6T(V^0/W@\W;bYH+.Pb35QUTB:0H9^CX4[7&Q?T:XeNLHT0:&aA9HE1+;
<-dJ+6577L2,=eJF;Z#(>Rb5[W,)I@F=N0WdF(TEGI]N]&0bDg5(2aMP>.6#JO-B
PVOW5YKOVZ8e7]<<1c06G(7LAV.@HFNcN^.7-NVOFDF]Td5J5gSf>Q>J]LB=Zd\e
MN=A4T.U?=3Z+C^CZec.0BLV[L1C][FN-2GaY_<L4S2^W>A_22K6E-6&P/cD1fe:
PBLBb5R7/H3L,BU[b9UU[A(\21ESVF1.gIP,.6\T<c_5=KL<(I8-JYA><0e)EP8O
2JXBMS5ZU-JLXM:.=&K[Od0e]CV:,VY849.^N=#:P\5M0W_C+,UOT_QK821E3KQW
^P?YcIgUE/87IUJf/YNIO8U@.7LP.<-P,5?.?gZ,f3JRUd6NYG80+#XRWUKP4SJR
3]=024]Y0(Q(RAdAY39Pb>06I1^A3<M+3>R=M\F0IfC2<=YgcW_d#S\@0_)&QaRS
CKdM]Be8D?Z)KgGI9966eTb/)05FD=EUX:DYSgIdSNX]?\ZfJ25e\^dU7SV#1bT?
0UL?0#2OZ6aV-CC@<gZI8b;><E_J_O#C+DNOd=CFT9;BEK]Z.ZSH=#?YCIXVNQ<)
FJ=<a(XHQ0I,]c2V8F1ZKKE&S.+3bRM^.H&&Ye,(X^70cFQMYS_/]1R3BDZ-5+=.
]T.>D_GRe8OB1&^NW]S2S,Hd<HT@b)?3-Sd4HMGeNd[f^6S<YFKbU;9K>N)fZ^]#
9X47?AYRX&?3&?Q,Lf,a?c+RDW0P0-I2EP^[+caI)D-J5LK:TNWGF63IM?Z29L,S
]LX1FWed?a?e,=-6ePb\J6;e16_d0UObS44,V)8d-/S6N?9.4Q)3H:TbBB^X6Mf:
3ZAa)^@N2Vc&AA@K9?e5.OSAJ]c/.3RRA._a@+U[^85BQ0(c0VQ7.@R/:+RG&PE^
\e1W;P8Hg3=e7IA6(TfgD-+3-^3S-^&E\XR63I#S[^YT57<d+7S,_eOcI;]MKdVG
U)[QIe=5R>^?d?O4F98-MM\?)(J^>UO27FP8?e0VPLeBU:A-2N+cf5YKG>G49-Qc
/b9SVM3@N4N,(5B0477B^?Id+F)^/aP)Bb^,E14,N?L&U?/1:-P&,C<01N+VU1)I
IZ>CUM2B[;I1G,,8eU17Z]_Y3IJ8_:=[,4)JZ-J6C6+0agBa.17_a(30S<0RP/OI
YcEDY\2VFgL>#Y_=#774=Zf62M88#YgCg&0^3\PVJ)0eOC[bE2A=cg3ZZBVZX\N+
KDLGfPX=3AM?T3Q9L&;[2C+40T;dW3OL;eG@04.?UCR<GSPDMQHE&Y-QLO\V1<W7
f=VeE[c34QY:(dW0ec\BC.5XbO>HZSKOHO4)NU,KTTAFD]E^MbCgAX7\\[]LaX[)
&C[7&7M^&T-31LYaHZE^5_VYKZXaT+bUZHLT195M4_HTSTPCMD(dC2MF-e<DFPT6
D5/2d\PcXW+FFf6D8A&dN[=H^+_@DcQUg;JRTO#1&S7DRD9.L>Uc01^a,O@3IRf_
\0_4_X[bBWL0e]eGK98H-)O,UA)>5>XFO7Nc,//1U1&aL80dId.U9Q<f<I6>cTD5
U:EJ7T/&4S1#JFO&fWGC.fYKEVHZG]FSZ+#ZUQMc#,IS1F?M6(E8.@aF,X8/XJ;;
9eVVA4f2D1-5<+-#;/G^.VO:])Ub+,EgOOZ^K):5KQ=D]Q,4IC]HRU\O\a2<?e0]
,T_T\8ZFEL\b-Y_B30SQ-ZAU)db.-XTY7KbCR2XG1IcOYg1a,W(gEO;8c8?O1GX&
c[RV0,V:T:VScU5RL@a7gDK]PZ_M63fX><OD#1[04Kd-V)A=BU(@72H+g)6a2Z,4
X57O^/\5ERCaJb/A2bcKbaNNc^#KfY4(Ng=G5K)[1)D:E/@;d,a=gGF&79E1U_bE
Y:#,2PVYYWX^fR.]/Nb:MUdf2)BeZ,?.QB0:_<Y&7X.1RgYW1d)<FPX^bUf/YTW^
NKIK<(=>)S^RU0FC;J40:KSfI/_]Z6H((P7R-8JZ_KPE8E:g@R(N/F)KF=.&6(>#
Kd/#)c^J9<=\\]OR\d],f6U.8@dgSCBd&L<N?-fMN0./P1dT)^(<eD+=7(A7D\eH
_OX#7[T>Mg?E^2=dPVNg5(J<YCZ7B9APV4(:bK>T<OH0L>F5eVUZF4SZ9A<K2S)g
)fWS=5WD+TYL9B8ENDZ)W#>1KJ;6\79@3a\g++?G1T463?ZWQ&fL:D9geJ/ROF-K
(_[YQUaf>,U/>-Y=#S\BMJc^49,UXLCE-,SZDNIU@Q;E(DOEBC5L,aFHIA8EU;HZ
PD-W:fPK:>3R3LQE#8Jc3(H#9F-2LY/g80b.LQ9f>?+8eD105g]M@GAV-D@GPG_D
]Z?(Y4)c10.bE4<GA1Bee\^2^JaPOBc+6EYZ;>VY4J0#9[)ILKWD]#cUA+Z73)ca
Xa)Zg&R.U@8#QA0#\0.7g+\R>B7RFE<O^fKdeYB#94?N98I>6BM\3)]YGKfKdFg)
[1IMc^)S@aeK#PdS1B/9BMCFBK48:UCfWJHU9(H.#FR39\fHgVWXNPba&B<:>7If
;Yd7S36bc,6ALd54^7EgPW<M?/3fFUBZP&<1VR_c9I@f;-(DeSeGF[#FYMJ#_\#[
1LJc+Z[;)HgVQ@fA?JO#/ccWWFg@:UDJ,I):4BZZKU@^6P3(?]@_CFJIY-D[A,IE
FbURH_7a)S;LR__Y3\gKW>ZHB0)fD4G^=DA:)2:]D8N6VNBR4d:#+ERb3_A-+fX(
6=#\;HaO3cGTAQS6dN@B(QT5eXCUcVR-M71b\81[8?ee>)^M>S5D4bW_)M^EE3\I
[64BVYC):>UITI.dXKB0\?]24CT?aPOc\..B1WTX7N/+PU5/,PdcN-7eJT#(eL8K
\@Y+Bc79Y<YE-70CN#WG[TTeGZ7A?4V46fXTQ^-HgdP3b34]cgFWHII\D5_d@J=P
6)WAOac1P6]-WD#?-PV4@J@c<&2RdFKZc-L:A(O,LM:GTJaN:8[gB=&9&Y.,I<Na
3cP8\MLQC)^U2I)<D3&=^T:eC]:^9eC)WLJ>,X;-d4D.P<_Q]2c0g0P:g:2K7GNJ
_#H+-(LGFJ<<?1_:/?8?AAK,+99MF,7DFWKOSEP3_:DYd?2ZPcaK>R;FJP@0g8de
0Y+VB1RN3F^:gV-)^0]&A-[1LfHY=8&2?57@J<AYA3.U2BSZWNXQPRPJ(,LZ7]-V
7_d(V&M7(S&G^dfB)TPMJaI04M5H&E._+&+U8&7)J0bIY95L#b45]6CKTW;6_4aN
TV@OCZIgdNWV8[C:>A:A[d#aWdB9BeC0:P1)6e5CD0aTd/CNX_a;a\]\ME#HCF(\
8+6HfM1e2IfY;+_cZ>A6FaB:VU)D32T/g&G>D1KF]46PfcBU#E/Ad,)ER-WeO)RY
UMX15P9M-ZA&H>I>d79H8+:&L1D[g.FOUI+DfbdB:e>Ife&E)Cf,MF(&3a0BB#(U
EE80]5R[XN]7/Xb2R)=#C;cOd?KCVLEG4R^C+6F;>(>3CSF6WAENJZbZHXJ-:9Gb
c[+/;(RaE@&J)GcP(EF>,&?NJcM2P:96eI.OMNN1a[ZH8V@8I?562a[:Oga@[Z3^
b.Z8/NVBP8Y/0(2FBRF7YK+N#da>DQa,SN49HE\c0dBZ:/gVJgf3Eb\QPZZ-YLID
Q4eJ^b:03>JF<MHS0OM@9E7F]_5PSc7@Yf;ILTS(:CJ3N#&a?dUEC-&C42bf.ZYe
]T]#C0)Q3GBJ?3BM[<Cf?HX>]aVW7:R8ZJU<B/1A-2]1cESH@O]@P3O<9J^SPcaf
0<?-^\0U-;/SSSQT0]T)U+c)(CcW/0?Q@Bf8IIJN3[-;#9LO<940c<;-9fK?.HFQ
GGDJF_QaO\dT1F.V(VDA/Lf-LJF;e2T/DCTC2FF1AQf-]R&@g3<KK<EFFH9?gS2-
G):f]6/fT^b#U(W01N2gW,O&.Y[HUg2&@,JHd5N8a=-Y)YMX8,+[)-gJ(_b4ZJC<
+@L3TSHZGZ6LEKMPaK&3Ee)42T?e#@5)?-L(.3fZ@&Sf_N?P6BN]2-)R@UYK?>(0
(V2@X?S)WZafY\eOYQ?MB^PFCT]]DY+CJOgO#>>N4?@KCETWNRB2056U\_ZCJ[FY
+E.CCg@5bg748XQ[4CI4LU9OL16&4MINJ./H;&-:GBQGX\[GZ\]E&OP\9c[GgNOc
BFB/J#Z8;13@UAK>1eC5HR5]D)F,91+7M\YQ_AGd[@#ND^F2_R2IM3A9.2O01#&f
>2^R0N=PW#R^DSE(Mb5<07JWEDA?Kb?&)#+/,D2>Z,?,+]++_TD\g.MK3H(cbC]&
1SPfT)U,,#M5&Jf>6bG(-=L+)#;a(dg#LHP(A,c\PU^:E7GRHP@Mf1-C4-MTccf)
aOA-GC><J(>b\(DO4D7)aX<eRb+C7]QS<\IQTWW^S.?TX[^),ZQ0X\=gC>;4Df7D
g[L<0>P5P?&)ReFXZ+Yfg:9QdRAg1L,Tg74<]_<Zd,6PKT7:0EGe8JGSfIDb(X=Y
96KfHJ7E4?G\TgM/^K><,C:@d&70(Y-FEKSEKgK[K>RLW-D1Z&H&Kc8\4WPAELRL
@f_^&:[Y48gOc,Y@7OJ^Y@5PLdRg\^KB0-(@D2.\b\D/UdQ(@-7d.I>XCE7^JHE>
669PK^U\V:7-e\\#C7\bC=B+-ZAL\9^4#)a?W4(1Te3_90FQW63)3,SO1R\TJb)<
@X?.2W:51;0/<RJ[[Y_C8WEI-5Y1,LPMXXa278TK8#6,AZI[fOU/f@&>YRf171KR
R:J&.M(A[?P3L\CB&A&V+#dbCKeC)XfE2JOH:<CYI96W+(WA7A\TUU893f_>>P_:
;KB/=9#-U_:1)7d74W]5_/CYaSBK.=TQ6,bFfAC^+9;aba,:.VY0S/6[8,LcC0NP
(KE15GY1STbQO7E^MK;MF;g_gC&O-9AVL1[)^c<&3bfCJ>I[3SEH(27ddQW<O@N@
)7LP(IAK+#4OCHXV:(AJZ&&ON<g:?9&;T5Da]WVgGXG\W_GO3cUBdMa[S58g:Rcg
HOPV2VfZVP5NKTeCMI/TfR\\^ON\]YY(FL[NNQ],_d54/-EJG)<I#CPdSK.^H-C+
AT3c@[LE.PDPbFPH;S+C=](_X2ZPLb<WW/\/VL-b-O@P;cCLQU,UM^TEO9,Z;(#3
(YTd@S]=2YA3Q\JD;\L]>A3V;-\V-#,=;WSY;7.4C0><<G_66Y3?EP5A3)7)5gdS
e?&JbDFNX^6G=^\TM]E+H4BfJH(U?SfRJ+B2_NYKCK2ZVERa[OG:\d+2U45/(G#D
.TM4O2a)S\SYX=J[:&)X]K/B#=H+5(O_b.,MbXU_UXTf0L5VL_@.3KX?ME\+J/e+
F^WVQK7L(JCIEK>d8A&3^c8;D26@T/2B]LJP^TEWgOZMMCNe8Q+<@MSE@(AQQ.f>
#0HR5A_H_9e^KYX8XPHSA[K21VRg,/\]HGSA\5L-MbL-g<^0;VUGXAgccg)/2fAO
/(MCT>(>Cg&YZ_Z,g6B#VP-Mc_\I.b11U_<3.O9B;_eU=Rbc0-cg0G8-N4/0YFbH
0#[1B1E-B/MQWXO1JUYM+#HHKM.].bH(CN93(YB\Z9I(7K5VN@LJ&Ub5UM1@_]Ha
Vg2#D6G?BS^0@aHTeJ+0(ZP^,4C^N?)W?>UX8E(]/@D#TY.WG2Rda](acOaG=<UX
BR_[&@8#:1f@0XSQO+2XSc8AJ@7&3>^RA:;&;I-NO@5JW6:-NW#G3^f>.UOHOQ<_
<NIY5L@M1^L)#M;7HIfR_=R.bP@D3TRf7OQZE1S^DOVAd#[Lb2^SXU=e2]K5WH0;
c8Y>P><f4O\3O\e:/0eHL>P@IZgVH[PETXeM8\?=WA,\9Fg=dF.48ZcQ_K10I?a7
Q@Me2+H@]\P]4a;#W(X->^Xg/7MX9=S6-D@Ne1&G?BNS27DT_ANX<HN>97V@Z7M6
D@9:;8QdNYWCTBVIOHN@R[,V,,46OA>=c(+6L,BEg[=LQ#[2D_EZJN1fe<N^d?+/
/QDZV7->H?2YaXC:O=UZ?-DCN]MKF37LfdGe?K39<4QL;VW.^:1@W@2SF.[eeF:9
/DA;RO\=.-+L[(DS<_WE(09:I[;/<-N;4Y#>(+&a>NFEbZR3<TAggRC?)+FIO>1C
;BA9+.CG[D,?HK_^)PIJ23N-\..1+f<[<5eU.<K2,_BVS@S+P+ZN)&/0>2ZLXENP
d#Q0IS(L<3/T,_fX@==Z5cO:Z4f]0YZ#gae_:]+0[MSLf^0\M[ZeO5#L>=V+aC8X
1B2MG(BT</HbL_R,>S3b,]f8Z^19999c[QCX&OHG,MO-<PT<e7OFg8RAD5bL+:FC
aG&C5;)3R-@DeWW00b:a&.2D6A<>-YA4L;63=N/-bJUM(F;>^[X+a)&76\1C^RRf
Z@:(A&f+QPKc;;)O5E<0,F,-W[RT:CKSD#=:EG/g9=#V5O(03[R2DdI,I;P&G,XA
.I5-_PXDWP8X=>;7W?)@&>,[58NVPG.)-=,Hg+]S(MV-2<?G>f4g#.8d#O<RcF</
?P-6&c7DWWLgG\eX/BAX2Ug;ZAH)EEHG6@aAVAK81d5=gVLW#KYSKXZYSb@ZgZ+8
XN2GX8_+JO+Pea_&YdCXQdPWWF2^7[c@XXIOD:RZNM1^+LW0=6-K8XTZ<5SR8^WR
D+MNU.20b7UEG/Ed#4KQ30P#Q0K.Gg(Q6f9&IfL)ACA+UK^6[ga>A4a3aH9^2B1F
(UHI0/)UB\[d;^7[\.50N6[Y12#HN:C&&ZM9f8]VV]eA1N=:2_8<T):AXI]@ca,+
^KSX#c+?[P=.LX2f#e_ILc_I-4@dd#L.9[Y_-CN=XMJ>cOH]&b7ECI6(MIFYd8^9
=aI;,<N,TQ.B>:3H?cdQ_[K@f1P5AYL^^eaBPUB)M0/eXYFSgVa9N@Ub#<@\gQ)Y
G?FBga6F=XbO4.ZX-I)UL>[#?aHd;?<J#aZ21B493_7+2a2O3fbU91cd1eOS3dCZ
O3XRJO<S-G>J8#X):O=T@g^MG&f7-[Y\<#\GI/W<&Re.eYf?(GU:8ZaN>WX#9d+A
BGWF:73N/:9MP&4bK?d_?Ha#Ug>2ZA@J[;5Wg,Q,b?2-0MM4]Wb:S=ZP5Q>PX=<8
#.0K1JD)\MBIY;,3@[gC4>(OZ;7Je[OSJ3gLT,<3);)O\;^(dgZVK1,W#SIVf+c9
QRQGG@1N5(;4YXY951<Gd46W<+#9_HC6@+SSPWEP0W93^^f/9BSaJ5_^UJ=3]W?C
3Rbc&89QND58B=;,AO.aO[G+_)/-.LCH,@-2Bb>?dFdeD/S\@BP)#J4P,VQL>C;Q
(;7X(>;\4&]D9?cG&f]b_8D7WDL4d>\N2/EP(H\:[JbFMVb;LI-/()g@^R\_)7/S
DVc+C62^GcZPR;K?>]B)598SKe]LcO6+4bH\E3OAeEfE0-,\9&N>+1;7V_+QSC0_
MVd3ed0)bT1HQ4e0YJ,H:#JWX5857RPad))04FRE9c+75\[BL<fJ6HcJMf^YNM.;
HM,B2cN55H22(HT^Ff[8/;QddXD11UdDB/1H=Of:+DX+2X5+S#^O8fd_4g,JGaA>
&c6>cV7GgV>M)XcKUN75LTPa4b&KZIL9^6HN9D0=^&NC:\PJB?68,EZYYX7c?3O(
JUO5_.R:WW==OfHVc(6NT@Hg>QHWF1_@NP4NPAJ6E6O/OW7:D9=_]&NPXgIIG7a@
&RfJc5\D#[#<U2P;F,GDCM_.ACKMg]:ZMWKI>9&28PIUY3EaYDZ2XMaZ@\b]/@P7
U_>?]?&K+5Y=BbC@>gP4P<5QTV_O8YKDDM8]8Tg70O?#I+>g#Q]MX,)?>#6XDZ2^
_gXHZ?SG2VWYda_Df^_aaM&O<2<a96>-eOgR&5TBg,N&MYT;68,RBSdKe-@0/-\T
AKEPXg_\TAT4@#:,GFaRV2/d6843Q@c_e?=9/F2JC2cFcGgG:H@5Fb3TPYJ&@e&X
V>^#C>1+V0@7W7+=S4ZYfFK5A26Fc:HW:.XfUQD@d&MS6<[N?RL\6N?FMN]:?FWE
F]X7d&_XDB[fT9Y2MGEW[Vd\&.Ef]2\<)=+::d)XX#.N.,gbM;d[eDD]G;Y&9BCD
=X](AAW-@1#W@@>DVY(,\<4+M6>NV<?TX1,I)eNa_f7+]R_<g8,-56_;I/gHX)Z^
,Vb9<Zce=BcD7c-Jd&.a(OT1^]DDF[S)ES:#dbJ,&(RL[/d>Y?WG?2_4AKK))gcF
1PPYYfa<+\).FcXE38<2>a(9:WIF;@g//Pf&Xe(CYERCZCe64+K\9URSc([8XO1-
^\V-(XNS)ec5Ib:4WZG&PDI8<D^U&1^Kbf709ZWf#9QFNU<-Q)@fI13GA<WeHN:g
[MO,7M.,)O4?P255ITc7R\JXCeX7OK_3L>^ZM3AFR>GKb7O^gRI^[(,;R:M8O@/K
3<NA(;L1#@cg7<d<=M+Yda31+bUYGH-g0^ZGc>7GQFGUfbQ&VTeC8Q,=YVb;1a-M
b&QF92#Vg2>MLH&2\cgPX]S2;DO.La,G2S[?Td[g6BF9JOLT?8M-Da.fdEX&,1OW
XML#WA7R<\-_[8-+W>&@90dT01@+6Y,Z+gPAeJe/QA:+GBI6;NHb3JFD@-gMR;L<
7.)fGNe@^B4V?PXL#e53\?R71/LYBe[+?+6J2QaO]6]LED0a)HS)TDQ>9NZ3D[3\
gB]VW21BIGb1=<W#Na_<-e_LO4^Eb@QZ=HRX:]?0/>47(Ye8SDQ2NYB_e-gdRUY5
XC@2f(N.J\:QE\RW=1;LgLQ;#S2aKH;_VOg=0bQ-\a1&>[SS+Q0B1gB:eL9D_PG+
eHLUg2YaD/g65Gg-O848CdLfUPOZDIKJ^;R/>1bHN-=[5B/2,,Z@6ad77Z6&OJM(
NHf,]7+&MfI:FI:N9R8/6I2@55=f0UL3G^:=@g=IK[&W#X1Z-7T?V@LS>0#<&LT4
c;R_@8E#IbF&?-24bL1GD?./U\P=O>8,>QH^[6M:010)L54S9#S+D/>>dOSAP[J;
XfYfS(M.FTQcW0@PCS6fZCU/X+c>;ZN3,b0c]T-S?a[<[38]Za>OA14H#DV=G&>e
=FT&eD,Z37Y(L\AA_T]XYaD_e_[e)e?(4cX1ZH^.^_,#__9MAeGZ2E893]Y:_]U,
X.D_Z0;8E<3DfCJ#SUI7BE&./H==Q#9?=).P:/=/.\NS;^L\;32.HCKOX@dPR5T2
d@Ia.3-IZBHX4Wa3Ja4Z^Eb^^(VG#GI@QDI:L.\>-L/8LXbf19C:=>,N&>RQ1Ed,
9J:1Y2B1N\XH7e.-G2X.FfGXOH+OLCd4J[G#VT\=LNQ-=;H6OWaVT#UBfccGOa02
:GH2?(116IUD[^]O)Z0)M<fJa:/D4HW_BOVEfa@\b2?MIZM,DF]:#8:,TN>&3U/C
#+27H27+A]U&#TSBT9]<5Xg.-M131.FPa\7M4,2cM?gVfbMUc-@dB3I374]ZfAa,
3dEZBM(b]^0^A1NQBP.HK-U?d)gR0MZK4;J[./R4;G4KaI6[ZFb;]T1<SHBXSB?(
:?;b<f]fRXfZ?@e[eWdF3:6J+30d\,;TaDZCVF:<ZL\e[4>8B.7W>QPT3+615aT/
;aKD/Yb;8ZgfQ[d8/,)+I67+PYE8ENJ>&MT;d?ZR+U7eIP>^SG2NQ^ea8C@^N+4N
OLA0^U4I^gG[GeIPa\5B/c<8fG^7_eA#JL?@cF8,35K8.,I>=ePBb#\B#8?^SIOf
WA>0^JC)^/#Q;=g^/OW02T1>K+a7=N+7.b-#_>XCg9eI20M)861DA:FAP?V6)fP_
8Q37&]L56eV78TAKS?eKY=&1FDS])18a]92::ReJf86\S@,5,2P#J#+g15VLW0gG
gS[YdT?/CUOCDe7?\:>UO=C5;NCEd3d@48.VQ/QSVgac.SYMYO>&Y/^\BO,73X@)
66BX=2F8#=>3C@;2+TVI(]_I8]5B=@TeFD)OFJCAU2V((QO-<0Z;AWGS6^H27C6-
bC/=Y]:EW<EXGeOFUa3D8W3aZ8KSW[,@;eFC\DP76IG8cQa<)QZK7^6I5d?gLIEU
P7;gM?Lc7:T0LE?g;R/A_+]1;Z8U#gPN#QA>0Z:H?[a^++7E;]1/U6HaY?f+-)>L
WaU.=P]--FECYW#cX)NF=X=(ZXHdbMB8fZ?J#&^(H)(,a6f]]2(E0E;d55_FB4WU
U5F=e(X0O:0#Wc7KQADdFXFM;Yd@@#\^/+.FDaPB2Wb6&e?VS[_&.gM:;,C7<1O6
MVSAL1YA>E[[??K8aGR3-@\ZS];dROI/f,C,I[AAbR^.O1C/[A-PM&&cbfbe\aF0
0RVI9X.EFVfTD[+QZ),H>JF<1,Qg[R8=.O@/2^WfD#/2\aO^]:be]1#[5_(+a;(M
8:e_GSD63=0.F)BfBZ3#=Y,VYY1fJFG>\8LI\\7(284V4X/g(YOLa[eADf\8)SfA
;\<MDMK_DT9-D]UMA9gK&.bPe282]6MM?OR+4>?:[cB1;]R,4HX#X9A5S7eI>,H8
6+-A.Uc00RYLPAcgL&]M>YV._3S:7CATWLP=><CBF3N(A+@Q]81+(MBMUWCCBI7+
)8/T64;HXFH8F&HGCba,]C7f2]S>#TL=,/aN.+0abY.SVIG,7VYAKX+V9<BP55#.
ISLMc=2P-;V:C:ACC&E@XedG>C7(T,d.CW36F=X?BFT+>c),T&77H^IZ@\[Z?]4?
.)D^TRL^]49>g.GH>#SD]H7.LO\-+1LN,WD9H[]S<I6,/1EL>f#7(SD>/eG5E+(/
Dg)c(T/^QL<^DEJR/3-TXL\G26^WIP_F-^#3S?]5eOKR?:]Q=_PW:R5-d+QL)^:&
<-5F<,.=1Jc)d;60dXA^E40S5)7HK@+bUdf&a3MBN>(ca@]B^WOZ\4.4X&YI:J]&
51I>)KdUYf+-^,EbLTN[SIX]6#T298<-1JE]&MK[M=G8IDYgLN4]0N3?SN)>KR>P
T+T]^]6K+N@LW+\9:1+M7&TKT;CE9@cNC#V7T(,8):V,S(F:g4&dQ.P39OH8?#QJ
^18:f(6_M=(:CLcEB-X]R#9H[X\T@CS8gH;K23e?aF8HbSK<Y2;1:-2D]8dF(/;X
@8CGXbMY0;ZR#D+LU1Td[Se@S&B\4VG_=VW\M@_gM.P5G&)\5Z4H&QR<WcO<)I6P
5^<,fQFa:B4A_5NQ&WI=QNM;J.SZZZ)f);>82b8U998MP#8F7AV05K3:VIX=(?>O
SOeJ/18IJH^7Ld#2::QE])-e]bO:=ZR\E-2AX>N\.Be+NVNg[39HND:.07Fg^D?A
[bJ&Y<OP1,K(I=DK3c;g@cN[+.WUH5@1fZ08=C/T^/^0Z,:Q.eMe/eK;1dK)A5dg
#gHYPW.MP8#Z&TDNP#@7+:eb\VE567Ab1@B6G/1Wfc(L2VY)gA3f39\HEe@F#c9[
_)gRZ)SUf\Mf(@^9]b3V8Yc^Md)C&+Y&DJAE&0;9_#FJYV5@+g>(QHO\I,;Xfd,R
D0X_fJPES>,K3?4SEXU^-e)9F_@F=1Q,S2Bbf9EX<YXC9ZXM9ZY4f?COC9<UP\N#
Ab-YUF20Ee^;)A^@e((C3OQ=QSEKTWTe44;f+d&QAWXJW8;\E+@cI5S&I.WM9+Q8
FG07?3_A6G&P(^a4WeATa0WP_?V<U1Tb;C#KBbX>#L,S)+_e)H:9+T6N0LV/:W\a
TXE[I.FJOL5g:,0POJ55[4<#8X>0L/9R^_RW]aXR&ZS9=Kf<DIebbF=WV38bOMX^
EQJYB14ZG8W3YIRe2:]eL0GZd9+NQCW[B;=)]e>(2;YIJVH4Wb1CJA##C(C0V?H5
8QSfHL=I7ZUH9R4=_a@EVW1IgK#,a7HCVJc-_PW]Q:]B1R<QZ9?c.;QD:Y::CQ&3
99.^5.L?[5H8UYAIVe\+D2J[aS&>bG2gM#.cW_^NT\[YId=?6E<-D?Z[X[<^XeZV
-Y_1@9WegB(,B,8?;B)GEeJH?gDZb?)FGUOa,V9(TMHb]0_[]PIC/):eO.+I-;98
(a\5LZAK<Mg&-MUgaL=5c/OAU,^Q37+@\X)>MeY&LP.AcTa[F=>VP,8H1>(\RO,G
-[_]H2Y?0e4QG??S<fK@Be1:96;4#<Obc^BSG(Y9ZDBPW=,A=OY:JGH>a,b[:)L_
6(WT=c)3-8,c9&F-Yf>YbMWZg@=Nf69dfg_ZA3<3)#+dV(6]7#>?EeFLZfVX^aFP
/^Y<=gBfO0=L2V.FG4(gfPJPVffYJAVC.^9W4(/beVI9bQ=;OT,;fOXF&W=6EfR^
Z,a+U>9[?N<?M]J;K.d\2cJW+\[DBe/6B/;/OX[LAS=QJ8WBAe&d;TTJE4N6B,28
LO6CENUX5-XPH_9]c3^Y5Fg_T<DUD3^F>e?V)W6<:16673aGRVP^,JRL0MD;8UUQ
UAgR.M1a.G6dFfa(bWQW(E^RC_e+:W61dVKLQ]/YE(3WC:D9=W7(f4O_DWH5VCT1
04]LUgSK@VbG8ZYg9<82^>7P?F6>D&2UJgWAF(4f_K0a8=,-=L.1H-(cDU]JDAX^
,WFLK:=8FP+MBd8-4]?H>Ic[BaDc,#)B^_L4(IMc8=KW^2..N9#cMM&.;UF<_E7U
@:=TTeK+EggdTEXU5KC5)Z>/0Ef9\8XAW.PW&O6+5X[/WRFAM[a(G^+PBWF>bCUD
_Mb1_,QQ\<9BHVR(L6aF=?-(I\J7QDL&)Vd=P<O_fHXVY::+5M7QaGK10G=:X<PB
,2D_&7K(0>cQ;Xae=X=SKGE8O<X4e&KEWGJDC&;aP.=d,7<+f6b=3O.>/1G_&=be
J/S)0^D;dHggOWZ2EQXOCP>T_]]W_cBLNFO]\[4F.@A)FQJ59C&\g.&WS=^BIMg9
B;[_40HGG[?K0(P\[Na()V^7T3MA@X]Y^LIg[>KG(29/fMLRC&ZL4EOT[gC4e(OJ
A@MHQ\58>)JR?U2Na5#+J<(H4e]668@S91?_e^fd[]UC(\;4bPY8#U_Y=a/[9;a_
WGEIB])K2;:0Lf_UfURIYf/VK\H8I6LBf^EBfX+.RZg)a\d413a?8FRCDNdT<V33
P7aW9:>X)d2Hd:7N;+@7=Y\2KP+G/PIP>&E-eGSLGK>V=Q+-J/.(D.X@2\63?)^b
L>8Q(OC1VIdXd3\MNY7X[L)W0-gWY2Z4Q0#.f8Z\U;)\=DGcCbOdJ>(\N/6;U)EK
&@WA-AM^U28gO(]DTcJ/1L;+2@@K+^cBPB64L17?35(7]1_ZC)1W4+)?]>ZMY,N&
<RTTa#06[]_80RZR2C]K2dG)H^EMCLE&]aUg2BLbEH=Ia+7AEXN/-O(VdgOTaMCc
V8X@J;R.BWTgMI_F3<[MIA1#448)^3[YA^aWdMR8-#]Oea@4E0.CNTDQ?4P^]E>O
5W)3I1X1A5W?We\NG0UTWVERKPCW;_R-@&.,:.9WPF@ag4(K=EAAc\W@Ag?9HPW@
_89gMW[bN#PH1f-e#:f/UM_&W:093[@<3==I-:WcSUO4&eJIQ)O;#8FHGZ[1<(^d
AJF@+1@+g&aTgWC:SRB++8K+2eHD3P2&E&O(+C;:<?\cQfNG0EUD#R^5KTI?I1(8
=53V/,VM+.<0.>J\YIUTTB./#VGa&dfWI-JfI=(2fU@/M4,HW[b8bX?3.:CRXXKa
U&Q&J_?:cg=3YZ;XHcF=g-BTY]8,E5a:d_KFN^=APCU8/cEf;?SQ[YEGZ-6R1+b;
LM#VXJ+.PY[cHIN;/P^bIKO>:KWcH?e&LZ8INK2b?&[F;\gg>HXX5H.9H.g6_55Y
RSd.U]dFDg1Z>/ZZ/\,_(6a_5RLbDf:F,&LXSFEKRXWOGNbWJ:XgOSMV(+-FO?a1
:Ed.?);>OU)O,fD@:\KS0fa0fP#+gWZMZH9IV[@DgW94R6]3CU?(V-BE[H_-ATAE
UN]53f40I&1/_YHQ25;:Nc1VO/K:O@0I/XTMAd2g3]/<bECQ]e4YS9N#?Vf5_KdS
-,IcC;)dQ1M(XBEdbdZd3;CfY+d-3fZNEJg2[XYD0UaB1f)SA7CgA>V>7U,UAT&T
X=[O&\HUf2&4CeCaJFWfAMX>5#ZO<@O(A3eYOCR\KANG;NSGR:4b7g4J=WZQ.ML)
KUKWV5NcZ)1+2YNa_XQ/0()9dBTNK/D,2bF0..bPd0&_H;]&,P]S]T(,NYG1RD9f
5+U-?B\YZ=DF7K8N]Igg6Z>Bd-OE9OeK#NHD(bPDT]B<Qc/2_bS-B2f/b_+\P:45
>bUS#7KF8f7J3N0C\W-TJ:5IFV-/8NbP^B0Z_&XBFY@<3AT9,Y;2LXW@&&(4g1R]
N@d@-&]8KdJQ>=PJ):8Mb9[;C@9[)(ULd1;b5R[3@=Lc,VFK>2:7,(1=292&-.@E
^VG3_e]<;/cP^4>IH^E>#?AAHO[:2ObL_3PI?>^\L@bG>-MKTPabKEJ>^EDa/d(O
)/cBf,C0N47b2:(<e:TY1JDAVF^/46>;YK26b^5\<X;<W@2P+VN:(2:f,.SGfDBC
L0QJ.f_-C&LRUGd)cPOC:U)>QP6ULKB&0\#.T>>g[,]5^YD#J,Y>_W&5(PA.(\K-
3dDLeLIT5[dNZ)cM^E_^O1fAQC(2Q\c,b31(CEUR,d,@6NMQJ?B<UdB/&<9Z:G.J
PSEKHg6X5??-ZK\/QQU70+O,TN=d5Wc568,Z6_WKPQVAGe0]GVY<BL-?C]_g4G.(
&Y;1Z9L61&Q-QSa\)e(7L>-A4\D/RKN.<(#70[#+eIS7ODF0K=CIYOd.QF7LdFDd
FDQEU=X8O<WA:_U[13XF_G@:XI8R_-#YdWPAG3Tf:]PHRI[^_g5_K(-)4+/VBbVJ
_0^&1+9CJL;HFG1I63^VQF[UCB;=E5LAaG>b)KIS-7,U+Yg5Q.F7>aKXdX_b3Z.@
NUWA^a;Q=P-YPO_@>8RMLDJX5M8,7Q+IffC[[WT.#1fM0d.bL(.2J?QRE<7(&1^5
@PYc8M1/c]TcMP7<UJ5(<A1HS(WYFY0f+19;^^QK]9U-(4TT5O08>C#]-f]C]HU8
.fLFZ8@U2ZMF+f?C^Q0TJX&G7@Ye@e+)JgB;ET.VWS;cXH_Pg/5]WO6PM9,<6NTJ
O+0D\US.^JEA/IX^,Db[K;Ve5Rd4R(8V<JBO-DO,ZJ3#?,-Q.AW7Ib&>?Se,9Z+@
PLRdT@g@?QD3F#S[VDB4FB(1]0?MU4W8>>27=,>Z25bdS4ZVVP-.-&^A6YPT(K,7
PbD<54+UF<H6(8W^)Nb5WVL]Fg.(#^M3F8a19LZO@NCO&=Z9Rf#M0OU;E3+K@W;2
.8Bg-UHU#06NYNMT8(_1=f+0T\A3^ONVXcHYaP7#I9^<_(->Y1c-DXLZM<I\58df
I(=266KDOd7N5L\FbD=^=_SeD[;g_e2T?5P^FdddO5D&;@C1)IN0CYTNA3;&(gcJ
]BePE+I@4;3F_I4&JY9].?.#Z9/AX=PQ)aRER/fJB?=3>gQe232R5O0ED785QXVF
07FC9M5AV=cf54#GXY06?03]##Z6#<d1LK^SAI9bD)RV4015L_fe9V+-SQZ9+#:D
X7#\(>:ODgQJQE^C;]+c8d88O:M[#CVaBBGOM<@GbeZ1a7Y7JK^c(04=UB24X&d_
Kcf(Y,+ONK^FC1Bfd3C78<Xa;2+f-:Q0_\EaQIbBIXb9YcA@[bC[<5MLYS/[f9/=
?-S9?JgVGXF#-CH=CT?#cHf<7H2L_1dT^gf(---&NX)fd@WVTM=B2]R,fZ;c=AYH
QHAX.bCH]6>3=2\A-C\B84?FPeb5<\-g9d1W)GN)K1&Vc6Z,(TDV]--GQ5bT_@0<
e3AK;1B]WW+G@[/NZ5?[_2@@c0g,K1<C9g(EYN@8?:Z&&54>V8S-[ULX;DC[_/c;
\e\_UUTU:fLX[U]L7D91]6D6aMgO8JH0aE@:PDK->H=Y^XCCY:fILf--8PaHK1Rg
2A5A66B:UV<GL#gABgF(TNa3RICbLc<Sg2)ga9,Na[#W:K&,SeWP;0fN4N>=J@UX
1#X;)]#B/RO,:2FRYV7-bZG[,dYF4[05X1f)]W7XN6Y2[.:bB/b2H2A;H_I\I=TH
0S3@c\###<RMD,g@U:-DZBP^K/;XRZ18(<&\c7L^81W3^TZGEc;K#+/cebf4?-dI
OF\_8Qb-I>9?49g)M;89.+H</G>>@1TV4^F_b@Y+=LYTOO^g&+?;fV2FRc?4]O=/
RaM8/:SI)Hf\TKYUS<1D_=;VBM2AH4X3/R;Y<KV,MJN]J0:L[:=_\O4FJ=#>@O<Y
I4_PM6-ZHNO20G#^df31<B@/08&4c#;G[K9(a;)44,9N&DNBb(a/JVGdFK7M2Q[V
ZCGMXT16T(3)eeA[WXW^3T[:#G41LZTYTL9bL([9&)<b[1#\R/G).#bU7d^.MH;\
3UgH-c@GPI3C8C.WM(THI/9X>HRSR8+:=e-^>+4a3gL\b:c\F=CND?<8P@+S\38+
a)VZQW;2_7E4&>;O:@8GgHU^]29W1J1+d+#,ee[_VOO(0eV.>B]F0/<<Vf:A;:-Y
KU<,7>>\YB0O&3I>Vba7TUT<A+9@M\d+UZId\E(]>E:(1G;6+NY]/W3\5T-##H9F
FebF<cF^#LBA0>gLB?dDcA1D>TMeaC8:0dMD,F]#d0BeME\\>X:22E<^8Y)4:#L+
c\<AgY2>cIHRJ;AX[:@[FNY@8889BF]]LeTc48=KHac4M;_ZR)@CKGC3R275D;@;
)H9UNe6WT]PXagPc@O82PN^FbJg]8Mb8R3c9]W?;/J:LSbX0DF47/.(AI^W[X5^b
37F)8ebV3P,W0?5@1aUe@Ggg=E=9Lg+PQCe?MUggNPYY?F\Ob0/+I26KdbSN[:aG
KNV\-B0,UVaU[E3L8(<FC(g&/B&NKLR,O5cU/7b5]KR:JQB&G3Af0bO@gJ3+&c5Q
\Yc4W7Ug4,MZU([SDB2@+=:D6_5>ed-->J+4)X#^&F^^A76/N/=(3>?W.?Q<)T_0
D?Y\E-HX[aNMGXX:eB197_6_(T@8I3P4He^EY1].0M6A6PPDD@:^ebEU<E9#[Y3H
0Vab]7,5XG>>AW)6W/YBQ=JYKN]B0SX/F/+P+/KL#FRFM.N5.Q&SYL#V/F\H]MXZ
Ib7\YR2>a#-XPABdD[N:ef.[-cHO\CCD_?ZL>gFNbJE\GOa5PUe?R(BAN&3OF=,8
JB7-#\a@_b2C52dc4dP?8H6]ON9X,@\#cV3;?46R9d(:CX7aTIZ2)&U-;.YQH\<(
;=NbBG-V)YP9Q(D]^3M+1RD+>L?7gXD&+PZB]D2P_:PRWg0bGPMb@Z@5;E+(I5;P
Ef7B9Y0KTJ/>:+]Ng5A(279_fdE9:)&[VQ>CYDAV-TX@,d\KTULJb>87DfJMZV,=
D;&DVNS/F1Ld+I-beYVZK8\FfQ-\@Z/E=^#,a@Q@]_S[M_JW9ae=\0YFQRKBMIGT
a]S@/MT\?BD\:R[C4B5/@M^K,?AV+FMI4d.;I\Zg@+9ec(.8I([-8^<MM^?M&&_d
(3)XS?N,33/83EW:/R>\VG)(a<>#U,-N:EJ2UbGg+)^OKRgAC_/Ob:PFA[4N,5(/
1DX63PLg@:C.cL3Wb;gD^DF<A&>T4@-ce;#QI-J.=G^Y#>:/:._I(aDLQZQe1C/a
a-#O<5g1A+A(K<bL8[:#<ZK&RANVXGDJU)WC/L-=S@5P_#P_NXRN-:fE=L88^D7/
.9BMCVF)B+H/8gc\FHfKQ\ZW2Q\@(6QKS-JE.7#LW-\UC;IIR]\Zf?gNba2,.&/C
L,^eUDX8L5D?8b0fWH=J?OfH0E;YMfF;IUX(W0.LYd:2C/VH)Rd@PXgbF:6gSWbM
>Y68W#d;58T88NDa0F_Y)d^=IPTg8&46D\bSJ6a?XPIB,7e>b[2Zd<ga)WLLWTXf
HDR_.3CE@+4YM@QL,D?JaZ5Q&EIAHL+TY64,DKgX1E6g@V96d5X-ge(4V_)<RX@R
-f2?3b@36JH1fX;)d1e=U+X1g(>T@-D=J/XC[P,Vg4X)ecP[e3\dHWED>a<T]bUQ
BYX2fbfSg?(_MYKI8-BcfSgA[]KeG>&f].X2.,SZZEENKZV2UUAfG>8?(KLKPFV2
U?T<1.G04B&-H)X)5N9g.69b.])9DE>?KCgb&(T_.__M2RNE^/Z:cff2gYDVLeDd
B:(PE9W,_[BX4>gD;>-\[:=(>DUgAD]dPV4a-c/QD^(O0]DY3dE+]0A,dbVK)cT;
(I/CH?K6U]NfQK44=LRf>61XRWUB/FZ:Q>d:Dc4dG2.MO@b^S39a@FVMG1BEA^EC
,NWg:W=06S^Q:EUD#+aJ.XPSE\W[)F4Za8NG8e,81J\AX2ff4M#e0HY6DV-KY:#-
174(_+S=[@QNHa:b7>F(FfU]S?XQT(8M8-]f+PNWe\LT3_Ca&e8K^/GPfBFEQ?V5
?,A[b1aN&7Bd>9UR>g5(@bPV5,88F41)DeCZ(_E(K2bSPgZ]&O8?Y_+9.1eQ+S4I
cRJ;AP+]\,.<#=IC1U],)>0078gOV)MP4ANI7OQ^BC9@6LT;9d0HgMUB,?67IcS=
QS#=G\\FRe_UEW&DgD>WF?DG>dUdHQ#O(PU;.O^VD&LOf&PHTWHBAF;WYfN<Qa)\
g+F-23B#O/31(a>W88(Q<ESOKX7#MM(b)1Eb@\Ze2g_aV1#,-:>+^<7X&6X)]bM)
5f[Xg?:2:>Y)ea&W::HMBNZe=[PSNLfDYI[/Pb-LX[9c>E#4T.ReJR##3M]/BR2K
bXCL#e;=YfQVJ<QRdV<CZX/73Tc.A4YgF1[E06/C^.MGYdC#Hfe\M=bT\5GT@]I#
b\Ve6K2&QDJ5N#bU.[1MAS7M(QDI-BLM@5:TR45E6<F)f_Y^1@#+cN/&Xg@Ca3].
:[WV7\3IRCNOH]-^/a@V:Y.5\,B^>X@#L6]1R5JB=6QIg(@WNFd+J.DJT&bLeUMe
CPNAXBG:ATZCO11O2)aCM8gE71@RfGfA^S27;[4TU^O2N(J65+dXJG16=,3]?LWg
P\+X^c/2VEQ+Cd3A&YU-BCDP&&FRg..L>RL+2[W>a;W6+^f;:;1-YW&_70^[NY@K
_48SNWARK+-cE^E[-UdA-YF-9)Tc?5U&8K+K)W4B.0>:ZE^,@/gMM>M\>RdSZ:2\
)<V3[WB#X^dY:>_?05,0IX13H#^=)_g/3>D^[9-C;=9</aW;#C^.708<_@3VXEE1
W\N,f;ed/WDfbRZG,6cae[a5<e9=1D>TOU0Me+6.VCF0]SXH^(29g=fUNgGP)Z5]
7dGKZ4/cC>OPV9RJ<Y^[)?,KL-(R;8E@6?](J=Q;O;OTP:KP0Z=_BK#(@]HBPC81
.6K5Z63>DXFZN+C5)c@7N2_fNQFfdA5KRdegCYE9TJ.7)5&<CW_T02-,(Z2V2cWa
ITfadNAd8Y-S70&GbKeOQ#1K6dZE33e,MJQ^M65J5U221KRg#N?.)K#1Uc2&_84c
<Q_?X.M36_[V^>TE=2A^<(,L7@g#;bIXY@,@;H<daFZNdBMRd.S,BCB<7AM^NV0O
KA/dM[@We(1:&Vc_AaF\36\Kd7\#>Da&c\(P]e\2))Gf5D&Ad;)_&aF6+W(LZ.;=
gd2P1a?B>5JP>Y:1eZ:])VgPO#)?-^)XIJN,;I\AR7S8[Z.#F]]<&/H#[3D-+)^\
f,R(-T]\Q[^^LdYf1^/>?.4TNQ6)W#A0PA#]#NNK0,3?S1RD__L>ZQ<9Bb(IJIAd
J)Y>V11+Ce(^HI(DD#g33fbD:G^=@>I7Le>)=3=Q3&?4J)A9:W=Oc9J8UJcF6N<L
(:O3cG_#e?+=?;6I7I;AWYX;c)J753(FD_J#KQb[S3L==gX/Rfd&?WP.dX_/BdbU
gH3Q(Y\c<=>4T;YfLC#P9feXg2#PI1TOd6K2?6RLOC+W3NPD-8<H#S[eeabe6HYZ
BXKb==5&BK=)>JEI1E0[BWM3(&KG,LYC/0-E53XE@GX_?=>a.X#&3R,W1)J5[_gK
VQ\_ER-A>^[U^YBED=B;RISBH+TCI<Mb2Sd6ULQEe2gM1\]7a3eDU,FJ1QVVK<\?
1VdLT@MdFgR#4J<BdNP>Z]Y+[LC4V1,D\QP_]6[,D<;5?gE@R?Z:@5/a,T.Q[+b_
L6=dRI00..AKD9D^B)8#KI2Q(\C)^J9+NUKG&/3(gfBAD2Zf+3<0ZW]K.;@KBBW.
IV=M[=I;H8>YO4Ed[aRM[]B;/db4dM4>GHLNf=N_BaM^H>PVCOB#EF[d4Jc]8AUZ
F#XPQ@:f#T2SHL5-H[K;L9bbQAQ1(9Sd5UZ#R4,EAN^,TL=,aA=TOTH@RfKV6.@.
,J)@-/1>==M18Se-7JJJ,^6^aD,^.&BO^POI6A&aV4cX;g]ASdRIf8)N.4/PLZ@T
a(Pc3(B8UA3<=\@g6>bC:A:N:c]JQafU\<4<b156D?6>AN\C3RZJF=<Pb1O&egHX
SVFNOGGE[COX&W\Kd@Ub4YK1fC:^Z6C\-EJDI1ZQ\@[#Q6HG[EDg=TS+R^Z<A11@
f]N9<<\U\fEEH>O4c-8b@V3B;<?3A.D=&,#Wg0cC(bZRMMP]<P.8Z8.0:/QEdMcM
R45(L4KAYBYbK[EA#[Y@/CPIB>3EV8)Z5C3;&&@N,:64g<\X=@aO7QgT1X+AIXRI
L]9AJ^YLBdg#&6N)715aJH@;98.Bg91+F_,?-.\V)#Q#a[-@4./N@P61\2TWDB<G
87<S0[gIG:gNd8P=R/cdHSHNPAg0>_FC/(5UN)g-5L@ZTWB[bBLWQ]9M[PV]?IK]
\GK6;D\Q5&@L@7ITf2a]Tcf;C<L10]dN6=>X9]X@H&bTd&76BXMf_a5>_c0OINM]
[U,_aR&F45b=A\W(F2XB+:?=&^DH+M.5.^KfUPgGO/R1@P&9ZT)4[CV;>KKT]Mc#
;)/C7fQ39906@VA,QOWA9,dHS8/AB31Y;4EdU[=_M>QCWe,1bZPMZ&M[\MORLZVf
4G6E\F>\ZN@1[<N5g&YW5<J&07g,_1=bCC=Za_:_YZ)\d3<\gJQ<SV,7,QCH>__9
P:3gUO=F^L=85PW[AB<N7+dD:Q6-03-\IZWQV2V+=L#T7AgYRC^bfSW]]JK01\@e
bRVf_IZV_:B;IRfSP&)CPa1d5R]>R?JCB?J,A^JG^Sb1WF/PHa_aOF40,FDA:OHd
?(D(INAGLG-d\;75RI6OJJb]a@+8E@T:feeD#)^@T=_R(T:L2LHeMC#1TK\,6Da1
=\.+:;1KJ6>&>ES/<B@-P[Sg/d6A-cbW2#R3R67&^cYNNPGQX66,\,,19=>+IWFE
JE^H84^--5Y[:#,Y:.)e3fS-Y\?VgY__XB\#Uc_NbEXNF-_-&)F9NOS1fH@ZIEU6
b:WLdF)P7L<SL7b=dGM(7&RDQ]BCS=#\41OZfg4J?b^e)S&&BXQa^]0#PK1dKC>;
+Z6GS]eAYM>P&E/X9]OCaf+Q>gg>N(^NNU^QQVVHSb0.<c9MT/bKa/IY-=NH3Z4-
4@U^P[IH1O2YUG>WbRLH(YYL?U4U)M/-E<aQ3R_CX\_;K@L\AHAJJTN)>.[958a(
MeF<4X)@dAAI)Xg4J:HeNH862V5U6&.=Y]54?e8JdJbS-:#,VX95UASIQ7O,gI7a
>H^Hf&D5>ARSC7ZQ6C=GT0=,PF0D6:/Q]U;W&C)^OXOM9<8/^ORK:-Y=JI0UdND[
,f5IVKb(]3EWKJ-=a36M>#;8c)0;2UAa\,KX2^e[][.<]6bZJ_fP1+5caNY4NfXO
LUK]:CW0-gc-OD::;[2:VLS8>/8W?\QW6HOD[:PMQ+ZD^LOcZI9KFFVU+G@3Y]HP
R&OeK=.K5LF)]fcM[&]J3+?g\^:f(HQ+:01<eZS5Zc):8ag28CA,&SHA<N0&,IdB
ffdU<HXH^MgO#1dJCAGH>F[TJPYSD8g[W09Q1D\f=:;QfF:3<-GJ(N.f9ZH+ZWd_
/#.372U8IV5e9)S<KHV,.fg?a31MZ6/gR6g_\=Cc@,,A9@4^<ZM]_F:9&Wg\:#<2
_;A&YE0KUggEM+cZ7B.@BY7-Y0M7AJS@O1H=1)G#]XVJW):c61=>714+[g.6<>J6
RM2,13C&@G;A@/2_59RB9=>/MV<_cGHPFA5_W(/+0FZ?(bHPNGF/6NW?/8#EVF&.
MER?c\Y+FO3PA/]+[+0DUR+Og^]85,/gM5Vb1ZTN?Q-0P,)e=:\<#c?O=Tcdcfc]
=N?9G\KKd[PQ@V8Z]AKH9Q_,_;LIZPZ91]B8G^^1+Hee]SbKE0#b^P_e?DR#?^_1
ZQ(Q@6Q-@N:^RJ;?Q_R),VSd>I@LMEWJIZ(L;SUA__BY]J3N,28MM1g;OcB5U<R1
Z<4eV^HYC92?ZYc_^R2DcK9D?A[9G].gdLg>G/#):B;I7(;=IE=?JJVP6d7_DQdZ
R<8-:<4?CY;[L3&P&-@aa^BaD;d\P=@1+NX=EY2J\0Za-e4=&,gBfg(C#_Ca5LDd
L82;9-2d6:(7,ET(WM?bE5GU;bZ:<68cLeV:=Z2WeXNS_89c67;Q?\c(d3:.C1\E
&_&a,6D^<;Y]fFG,]_HfF#5[--c=C<&:6aEa81Q_<0;6]B>J?/:cI[^4;Q1,IW+2
d0[^T#bgdcD,R4F>XfHKOJ3LJ.eW=7UcQXMNR@6O1#e4Ka,5(bDKQKVYXM[F<8+]
HOQdA1AX+cbI(X>NEXXMW@+(4:K-@J01/CWbIB>gY\2I@[>g,12#)CRICG#QFY;\
@^PI2)5(8a&>=fg)PK9RbD)+;J>#8]V=ZeQL_8/>PR0,-6U?L_AC85KWI,O1U[3E
eSJ^WQd@Y/TGVFK(@NQTDdNW:g1JP>#FKDI,YV+\P:Y5M4BcXL;Cc_;c]eIQCKXH
G#V@7fcLB[J(?DKIIP\NCS9.S/f/6^7JK.V[RWZ:;c7G<35:cbICd8NHO5&+UM1X
5\W;@I[T+?6:VVfUJJSV/DR#61I1:[[,)@bCc86BCPOW5A9&A^P?0FZJbVI7AXNM
ZNgVH:UU<UEV[_(RV&./M2TX:c4JL6ELS-SLKcU]+74]:+=GQO<(Odf(;PbK6<C)
RM:SAM,dJ[[()R13aD)^@&9X?QC<d^/\+,LJA@.XU6_RW].EV8.dLKe))T2b64UX
ZIJ_X@3RS\=:N.O#=PN_#&LL3fbWJH0LbEaO\\^N+c@dcbX8ZPd/<69bC4DAZI+I
JARYKHcgLQ[R;K,T.8<e@&:/bMY=e2[099[L;<?LQHBXRAZC\g6L45>_>dT9Z2/Z
@:aO7NCH@#@<SD#g1)]S>2K&d,VU1DY&16R(D41ASA:3W&,/Y[&/B?AUXeX>K^YG
J6&5fL5,(=g3@bfMF+\V[M@>HXFHM[I:ML,0H,TD;IK12B>J33AY3c6:,0\(2?@b
=\Z<]\9&S>\Ue9b-][/H:/&KadJ[UfNEE#/Z2:9SB,(K4Ma,4:;.U7L)Q)C\^W68
03=W#?H=.e\G2&5?;UUT<QG\]#Af-,GH<?R>INY3=5.\LRN\\^6,dD<XA?2\((_B
K/=9P<K32cDdgXaFSab3)/PZ[b,;TU9Gc6d0_#O)ZcGI@cIf@SA^[f#U-M/]OO1b
.WF<PNR>8Eg9]bbNF@H/9,SZQAEX]45^T^Nc&ScGCH;HUO+1ZV3#]6L(_ETbU:O&
+F/dWX)0Fe8HT^0LBL@+;\B0GXFJ0f0]Y,E4aYC^-Ea8]:bM9>6#Lb0@SK9W\/]R
^(RaEgO/J[IDH\IDBS\A2HMLADeVWY<eb6I_BdZf2[RL5C\=/aYE_B&_#42B1F+Y
N.9FH4-/KNU43Me):;KDE.TgEL4E\QI2V;([QJR-QC:BSgXE:9RcfO5YbF<3K=bA
:KV87:XIf,.?EY[4^XI.+3@;FXQB9V=g,0O32#+RTL&H+a2M,1J(Xb9/7cIfbEd,
;M5_[e32;VWFDAVF4>-K+EgY,@[JWec8Q?;bS^U.U7.c4VfbdX55HdX&)a&gX(&3
@Q;8?[ZF8M_E#gA^NMUe(=WL.B]PDXbeDXZQY,9D[3P,=;CS&b)\&E5OcCa=)/E#
L(SY?VAc?B[VSTR8Z)W\21)>H\G;_.\RDcdNY_,>2gQ<\3YJY=3?LL4EbY?DF5U?
aPdDWA+)Zed,EHKXMc_@(61AXGHWN)1D7>_\Rb,TC3.=fB?d2g/)XZcNK9-6Bb61
Z\9-9V#TIYI+-9ZDCaX>,&WV<[(T25L<0,\X>[>aR^O3/ZIB^Vd:#M#.Eb\=[E2J
.V9&>cYC<LOQgL,ZdX6EL.7K&dOMNEQQ:OW<6S<Qb2MAL+T##T(cB<G2KTg9;A@&
=U?-<MOHUQ?I/9J&+#<W:G6e&??b](&:UGg//)LSYc2a:J>=B=:6[L08(2PD_E1X
YgaZ--=Q?W/d7AC,_2R^]1=/A68,2:\XJ\\=d/WU5;T2;DcfTFGbaeAE>dc#HE7I
I2W8>P<V8XLI,/;P\<.2:LTJ(gW=VKNMR1RD0IWb2Vg<aTFXgY72UC6W>gO_e\5U
LgZ<f_K:?MB82<4gB>PZ,[PNQ?]XEUO+P&W\\,+9YV8Qe-3YIee2&V+9:@VYd#RQ
&^T0+dW@)c=eKYga/Ef7#7IT+A36@)&^\C^.FgB7_G2-:71/T;=?CKIIMUAYVBMA
bT@GR;G^ZRC.=_TE5LYG#=NDJK38C_D]-,\8/,ASfWJU#f\RF32IMgQ=-&SLgg/.
6QGR>RVaGOQFV>7Tc8X7T2N<KH:P5C(S(P(1X<]=7O+KGG(M>ME=]S)P9-?FR4ED
Q:9,#05N99#N+=&)6^AeW3Q:B&S[IFcPCT+(=YRMTZ2:Gc3A^6H7H<GO)a6B?:Dd
:XOANA,YLa8@ccBYMXRS>2I<++>D/_+)L@6#G=K.a=C2,?N#3?d5MHROKQ.D69M4
:[9SX0R+AKaP-R=#9[QA>I:I_7+&KME(0P=CCFg/;2,9R3fDVQW#U=_d&OD0&U&F
X4(+D,9,Bf.@+JD<//J0c8H/_b,.\D=&PUca8g1dBV0C-.UH5d_;9YaD7Nd8f63L
)UE2479E.FH6gE](/f4@SL,I#SSST5L7e,_YRJ2+Q>7E(@\5(N>>XOGf2-.MHNNf
/:=2XHBd]3NU+D=B+SER@X.EBC?Jd;P9@&8cM@Z#0]UXeDI;Yc>6)@U+-;,aeb?#
D+,I.8[;1+][L3#ADJ6SL.X1/^WV(E=JQ2Wa+<Y;<KA;@9c.C+?J[cMHF)5-D(=M
C9_Ca:Y]E)Q,C@9#6X=+\//LQL1gDOROP.Qc\b0UGAV7U\3]Z5TN-=bM@KHYC7:C
33#?GAL\,GC2H\cUH]MGW,U@=/:2f.&gB0H:CZbVd@L5=]:=cg&c>:_>J#0UgW\E
-NRN22;3);aX=2&V5])gL11C?C:FQf:c6N&K07\WgFEb_:PR<3?e.5H-&99?(^a5
bRB=g@URfML6]<LgOTF<E@BM)8-1PJd?-Z)d#aJdG08UQ=@U-0(>5c#:LR;/BDc=
EI_SPDKfg.V1NZEX2C0IX[&0a&<48]>FR(J\gB7Xg/+;C?SPJ#OcGHO2WJE[X^6K
+[D6XETC=E,7QEJKAZL5:G786MPG(3M&c\YE.bb\GPUSbW+aa.:]a)V_M]Bc:e>8
MfXD)L:OLIUCc=g0N9F]EQ,2C@T,.d;[:V(Ua2L8HG8F^L?TYAZ?0S6J>G/Q?LeC
45XH2W7[MK;?R/65]_WM<\4X:RRN(7U.H4Rg)=H(K^R6e+G,(1EP(@Jf;9NB6QGf
gQC()1GMJ-5,E48HaQ+VV/@cLQ)&1A(<3?-G:8BADT=[e/EZLR0)4(f60aA2MD0+
)V3PUBW>f0YgaC,K2cYR&.0Z=4]/+dT]AUEfa@/PJb9HS(_.ZN7:aQcKY]b^c&9A
bL=Ne;WZN>bH@Faced0H^9+2Eg9ASbNA-B[ZRdc?GNY&G#H+(5-BC>#G^aa2bLF8
2\?9_X0B&a4RY(6GHg/0?/PKHB-\X8GUN_HJ)E;Z\B)CGPGK-fU9ABQ?-#/Z)]cV
G^<XVGL/ag8D9L71/SLaI/&#9[@P]C3+[E@K?548]&1HaCL)1:c(8>HNgD_N#@_<
)C3).dI^Y<]PV:,B>JMcU^5]>]f^@T[gFD3WS(F8]3>e720;[U/RU]#G9T75_7[;
X9eP0TgRW<]R;ag2\30K[8b1Q8V,f)A0E3/0?fg+2OD::d]CP3-4/ZXcXLNJ>]Gd
,f7FSg&_-+Kb_2@4Fa+77e2DFaf^d>+;W6FA&+?Ce]TIU5@V,^+W=)f9HE@;DB@N
-MY)]1WUQ\O(_b-A-1L9R&f:c)5I@A7@4M7W;[J7_VV,RTMN:[(Y^OD1WA].FFEM
QQA8<6&a_6SdWLV?+7T63=/EPJgbXU>#c_Q(5D<6WeR(9bf+V/SW,91?#<)\W7F]
+6PNB7?HB<NLC#B>cC+(^,;Q)_0NZ7WTX45f@2Y#\ZB;384Q@5/E[5LW5ZRGX1]e
ENZ08]JD2+eP)V/MH++d:A2UCZ_5HcJ-XB08C7JVS[XA08RUd(aRW5@_WE7&g?A>
=1d_?>2\dA_e<d;HaR[1&SgQc0>>gX[Q,NNbf[N^)<RFQ6KQ0M^D/F]9gd5Y4c-3
P;.B.51GB[A.@&caL_N:RHNbcA=YaCcSAfBW;&aA^&W;28bG?YS06adXYd+QONH-
G)bYZ)YG7XNAR[&4J^YWW1==f9Qd_d9U3H]O5a@J[H^^^FAM,dR0S2IEPQU.RI:R
V^a@,fVf8LdZ3[RUORWU9OSW^,](B/cEWaX3?D1eP\CfNf=^=N6?aCJ@HaA8]+JK
X8,X2&IeC/3EYAP66[E^Y1ObM\gYWgScXUK6(Ed-JD^O:IYJO2Z1I7\+HUC]<[bK
4S1F3MQ.H0E+Lb32@6c>(N+VdeETLC0_L-R48D+\:_7YYbYM2RbHd1NY4?(_G:E=
\<9@a6@XdQ9-:+3)cceYBR3652@_;LIfWJ#Of;SL1MAVdb6eQB9QZNdZ+,F=LUD<
M#+NY\5&LWV?(+>b-3&F9_RE^C.7bd=a4OKaN[BB=.0(9A>O]C@C,fPZ4@TdE?+X
&>^O/O7g4:525RcC9\07/GIF4gQ;JO@;^cP6:N6+@fC0b:g3-=[,I&()[g&[DSVM
0=-4^GYU@4=f&VU^-f=@P6/5H)9L\S^WP>,E3/HPcM6D3#7-+>BS?-]P,\N?GRf1
-2b-e#><1c0:^VRgRK+RP5E&PE^X).G/b/#c2O&[_6]eU_cAY5P:6DUbbM?G6\J(
&AJ?.I\cSDGN0QTQX;3#0A#<W8L_U80=Ng>b4U2=/_SMN,NB<5Na4.W3eg0TeT:+
<YC2E&Vef4OL+04aDFb\Bg<X_-J]LZILL&Xa?FCKGZ=/).?(M<d_#\@;Ie(8HWGf
cUSgWOL_VD3T85ZW,8K)JKeYA:a8YE4>_(O5>PD_?:C(,Q595,C2[?:,EK<<LfO4
+-Eb2F<c^LYaJ.LD[ZLT:KK0M0.Se&?ZXdV\7[ea-)U0J]@-C<6])3<D.E:\IOJ4
\ASO3+&@8?_9=J_GEKcC=&Ef5,CP(186Z:8M-G&69&\2ISL4K>J0eVe@N8bQ?I\,
U<(A1JZ:a7H-\/>7^@@K^X.c-2?1Gd5C_+fgaDZ55TSefbfF;+cAZ:L2U?c5[=L1
:.O]-_.(ECJ6.8CUg175VY+D0a0J;)GD_.WKBE3[]D9VWA_MQL-HN&G(EAC+&+e.
+23^5^dL+CA:]^V+?0@7OJfV\a;73-Pc/4@1G#G>7H<b0O+603>+O))D\QV]Q@:Z
VW&IA@Y1-5abQR4)#Y#TTdU47J:609@^dP<@.TFAbD/8eUGa[@@I>P=5;>09@Z<C
_G>I1SLg0]3[aN1_[GC=-=aX55PG29<AVFR#Z8O;,>=aK#FWCIba(\<^Y3a5&gcW
=-5V#GU(#6L]9b#A@;?CeU9YN&dLFV4)c:/O#e4c&a]^#TF>EfU_<GVT6[T^B@[F
U\IZ?1)f1W<bJf5;3ASU+ZZT&VVU;MEX8AYFM<&D/6b<B-_5U=(=IQ;[@BFSC\41
#[cKUL&Z9HU?P/P22bBZP:#S,T^8@ZI\CO\cKU7R+ZBFZGU01.EM,3S35^DBV#:6
#G\g6?):03Kf9(8GRH+49),-VA;OM1EU+FMf&0dP=I9G]5_=G9d;.1/+T8:JA+_-
-L(-4+,#T8^C++TNU,F(#eBC/@FEH#JO,<H&F\EbdO4B<a\XJJ,J\<\\<J^\Z-S\
@WG1HcW@CK&B/]e/>4+;7cPPIA?Ib/A_dDG9_dV/BZQ>;==4]5W]aa8eZ:+1D_Re
<XJ5?7_9(d(R22[I,^f0K1a<8W#87(Q/0V(F#Gc?JF:a\.]aJ^954S&/^/O?;NaN
@03H6N3-2Q#V[1d_eL+f@-PN2NMS#Zf/+XM>UC-dS0W+CK8V.Va.4e]b0Jd[IK&N
CYRUP&aV9C]#?A>9W65MeH^6aUfG69YZ<\H\OLQ6KBg#D<FW\gCAQ5(=KeUZ:9V7
2\Y=c53;@ad+>Q=F,8IYf3IQ&9-CPeO768X8G_,BKWHf5&+M[f,.B#.QFbd@Q:0(
\J/JM^+7/&]OJFag#D^[;=F<DH<d3IUM&G=MH9AT-bba1[gI;B=59G.2XDRNQJ.&
6Wg[-V?74906#dcggD:W^-_2eTN9e\C<].HTQB,@.@#_X>2?60&VRLS[3PV]YX+]
fc1W?FD+MS=RJ?f8V36K;M(O.2^O:EOP2O4X_-:eXLN>\<1GBg9SDH25e9/5BZ0&
PM.cO^JN=0?.6.(S94,H0e2RDL/4fI@gNG.>Fbc)NB;,++?_\TeX7[)eNE(??a]-
OFg->1#0b.45.1dV>a0:D>-a[]a,=g_3f^X,D^<eS:PC4JP4JK.)X;[-TP>X^?[@
,K=_WbWNW)ceM^+Z[6TWe.&\RF2<M^_N44Z?0ZMB_+O#5U^_WO6+b@^_\L(<8Kc7
NgHQN.-<fJ<RDHJE/#YWY=fET#<MA=3GG:S98@b>/+)<)&>/ZB,1ZB3L,-K<@:@#
U6^<QN69[7W62]A4DPN=EYV9De/4D;d-K,-9]/_XXb3R5I]68^MQN5J/aYSI[P^d
geO5,U?2FM@+1?Y9N@LVHfR2A;S:3[@CTB?WA3=R9N5@.M#78:W5W?)#T@SA;5I<
@a6IPT/.HQNfeg#B+FXNZB;16Yc;Bf<2)6K=#UU\71MaF&Eb=BHa[P?df^:G6S#Y
IG(&^SebO^KI(OXIS2)5/RVF62&b9,a,YJBeX,RO[,Z@922_[^Q:N\e=])Z6Hgdd
2]W:/bM8JU>KcEE9Q\04VI&),@<3dgMGVY]0@@S=/@@MS9GgJ(LW==3,-7Y\1U\1
+9YVVU>XAccIS.H\H7X#T30gT1^D^91&G2M2f2TZC6;P&Jb)50^)Z:7cfL<TFf(G
/#67)83]1,5(e@WQZ7_XJT\e.R?AZ8ZGZ7F1;^<#)@;T#Q#>If;8,V4)eEBX_/+Q
UgWM)ZPH#Ce9bfWA8GCFb:)W#3WCG@bXC;39A7HP6M[?TRQ9EW[0>@+83Q(ffCV,
8JK4&#.8:(]DK#Id8,>-/D@O;2JAeP;O(VVAM2VaKVcQ7#R8W\/WPe=3)H/J;QLX
F4^LT4Y06>T:g@:HMK<6J5J<1P1>f-;?V_,&d5g#C4)S-c8Pd9AL,G;>V>a2J4LG
((1AU0&^XbeZDV(P,&&PYBH7J1[41UJS^?,<IX8ZCOP7V(T4c-aHJQ#+:R:Z\_\b
S;-2)M:1^GM)QKZ_<MQd^DGcYeQ7c^bWK)cH62.CNZV]5g8,1;78>UF(PR=e6(G5
5#e,X7L(X+XR]_ed0]]7Va/)7g?G+JVIa^V_8e6M/H&[H7;<D+@^D\GAHM@I-UEI
IE:fIbG<)ggbEa]M;6bF5&HcdZ]XV6ccdTF6:/7Od)-c]?1384edFI0CN056]80<
fM-ZQ+C[GUF^b:UY^<_4\]WYR;eF5(-a3b6)76OKW:#CM\(CENZRJYP+VdIH,EJe
6/=QG2I8#e.JO?D+UGSJI>H+CC48<&L&=Q4dF&Q4(>WM59#US+16bIR9,UKW#fO3
22CPg;:H5H93]9<-GM2b:M2NA>g+a:;9<T&gFdN_,\,72XM>gTB/T)6:(XX#7=Ld
>N,Sg+5M24P2K+MScY<[33QPTd^9)\X&Qef#85&(GZ).(C#:4^MR?@DP9,1Z_O,X
,-OYQ+-D9Nd(Q;Y)AH^.>gJ.9RPK32eUQTfOA-6GVU#=NW(:>[WE&f=dH6/_W<S>
97C7-W/6L);]X;Y3#M,C)C8,.;:Sc+C/;AYU1.O2c/OG-4^((/@@2Yg;KT0A/[RT
7>gJeA>O1Q)?Cc/cgf3ZWYC<X0P47KW5<T?\CKT^a/g?QP8dSQ05?e4],aOQZeA)
D=H4P9L5fcEc4b5VdK?3.Z?0e036ODN<YV9</A\].eR4OY4.0e6BbZ7W87[B02[2
@=e\Xd?1-PW+A](CM7He]B,&@<&Oe[=FUKHDb8RXN)F31HAb(:8gLAX.8;eM4?G0
B-Xf=I+0T)d&\)J5#1PL1a4M01:3DS9bOBH]dK#?_DUW1.=L0[YZ;1.f+/4^8GD2
4/4N;WB2S>BAg,TE&T#H?dRY6M@;CC5X5KH/2O9XQ=)HGCNSfCS\EPdQX6MKM<@G
bX)N+SLS3J(RBN3DefE+7_NI8/GO7IcX8EG9ggG-.ZVUCFG09(^ZJM>d3&c@+^c/
FJU,A1,B+gQ=CBCEM)SAV&C;2F]171=Q9CM.Bc<6#L4Oe-/6VBFOR&^gM50KN.dB
4K7TUM=;-d1E6EWU?;ed1U2DQY4;(Va6Z3EW?VH:.1T2B1543?_C#6UU>D<SL.NA
Z4\D3bL&ccE560FaRaLM45Fe>=[Y1bOD[=MF3KM2\C:M,<(QXbJaQVfK)529>L7>
(U7:,ZISS@=HgNW#MW2CBAWg^GCM]=Dag?,,>&?AK9eOYO)X[PPH&0I^:)^62JLA
>9876:1/S[g#g4=]<?S,.>\D179&&Ee:V8&UL-#6Re3[J_1>]XVS&[&:C/??Z:dA
f[LF_+eTFDX5FF]6Z2X,C\94^>TM6,]N4Bdc3Pcad:C-3Q\;.a@\#:cIe]_V(FRd
>@8IgMCZB7ID@26gBPMSe69b=+S[:YYQSbD3W:OKb3+J/();9\U+N6[SMPGWBeTZ
-^+ASR;)AWK:eJOfe-S/Wb<C,VSK<#@cG,/cQ@D6W8[(]CH5a_R.S@5+E]E;77J6
HaZZPL;;3K:2].<a]ZYeYO<WPVY3Dc(44+M<Q7]0TY<CH(HT53<SYT;U+I:]BTIM
2+L\R,&7KQSDS[/1fa)^>Yfe[49YOKKL0AHE1DT,+8SSOFCSNefAeM1XF,8JGe\C
F07.=YL<Z=?Hg>dPNaN7E9,1X)(e)>XAF(3/Qc>HeX:>f^&:N3C]@S&-Z?(eMKO9
f](eJ:\;&EAC<\:\YJ=aV.YY^_LZ_@Y9/EH\c?C5K9dPL:B547<K5LYE.U8+B?:N
U9KeWRN]RdYBa(@9)R=LE<gd4M&:SRYeD.2\12ecd_M-IXR@XK4EJK8O]21:)<O2
K?Md,OSQ5=+&<;C,,-30/5=N:Pf[2Ra[b?K-5W?Q2ATYUVF#bd-=F\[HLDG;COMb
.2GQ3D?/F+a8fJ:8AW=5BB)HW-)@N=[;^M]TV.e,+L3;cLDQK;/O#-6XUT=5)N7:
UTK.E3PY6&EB-/ZFKgC<DX-]&]eUJ^X&A+Rdb[I;2>TNc2=R^H<U)9#ZaBB/1L=;
5W4a48c+MU+aA9=1I4K_A#Ce\:.1LJUJI#SJc[Kd_C(GRK8ZFD5>-P=S/VQ=M55E
_,5N]DF-TKX?Ia(eVJc>.Z[-Gea0H5b2Rd-=5&La5+^bPC5[0dgCc#Z5A@6N#TdT
.8(]g/7?FGg,47\g_QTBZY^UGg&gC4fMW;dc]XU2D>O?,ARL73NN;PF&40;E7A3H
@G@=M=+2ZLD<K\bQSKOX41FZY0EJR<C3K(]b_@E3#b5?3Lc+OIC=eEEW^K1.,&0R
VWEJd[VA]Z+0d(=E)8e<,Zg=;36SeM27PG.E4#WNBRF-S:AWLEUP[FgDL^UO[PI8
Kd/17^9_0MZ,;G+d)KTTIHJ&#aYN17C>.M\Q:PIJH?K1fdL98c[NR]-W_Ja>R#1,
?-UL(S)9X?P^J\34Fg0A;^VFQ3HNWOVJ817(e,K63Bf7BL)VU=SJM1Mf\,REaG&D
__@KD__M#28efL>C8F.Z,2JOaWJSGe(5-+1\afOcBP6_bcN7]bE#PB7J\afQ=]EY
>&4@OUEO@9]WO(_>e2JP///^0AC^L(L@3WJ&eVUEW^O0RY4X??dQ)8/^T7X]VTO?
[[G#8\G+(HGc\fK/LA<2b;J+#TC1#a>TAMKR#_fJLFDEW7N,TTB^Jc;+5&f/be2:
IN6X_A?dL9eMK1X>URJ:G@g?[_AR=T[5HP.=WMUe#5FVgO/Q#;EHeN[I-Q3gBW@K
TZO#bceVQ6UX+WWc5BGM#22^L88SZQD&UAO19AY60&f<WTPA\D_YI[<aO3:>e=U3
2/c.J]Y.G=f-[MEGe0X0\A)-(X3Z#5(;UD:]#R-gd^KCCGK6R)LB.??@FFd?6.bJ
NSafJD#ANPF30ZOb_Be[J]_+SR\)?C#7S:;3A<ZEdT/gF-Z\+0)\3IMB\1+W5#NC
CZce9V8\XMBE52]\;GKb4_L/(-3.JE:dFFA>,2V.QZ]AB&6?<DU]+V82V3ISO7RE
U8Y\O_),FM^VR1QQNEOTQ[/ESXL2.0I>CNPH@II7L:E2Y63HAU\MKM^ADV,F4c,&
IMHgS>4XKJVDIWJ?AM=cH(1NBK&c)af67.9QdA9b5-]9aG:d.\QU?-d6L4V[KOY&
e?&-RSIf3AG<ML1B>f?=fHK\?E<N0344S>^_S>I(2B&.V2VIHC7g40bRV/XC(H9e
Z#55d)-2RO,<ZAbe,;/A7N=c_8VXZfJ[Nd9NK-69?f.X7\4\WB3[\S]0ReXa07Ob
X<YDHcZ8OS/MFgD#+31;H@YWM.VU>TL\1CH(HIV;1L)+NN-RNe/L+\f1+6/d7K@>
;?1V?eQ,f4GA1[^W7c^9.0^7(=Y1#^Z>]-2ZLU8\71)XKFK#UOBJ)Z#c[e-MKb(@
S&M97?=.Dd-NAB1@)P==G9(cdCV5(?F._eMUgH?#:[c&4A]a)I\#,IF9S1.U00>B
QJKdU]FJNgKc/c[X]K(FRWREPGLc;,c)4;fg14BS[]7^<gQ8/JI:Fc_T&f,g#4:]
L-P8+R_);K]):g:5)?]^#bRe;0#[J4/EeYU5V/BW\#ca8#=?A)WCIC11ZO?1c@ZX
>IOVHW?;NG[;-MMUK.W_#(QUT+J7D@&0)^OA7gP-a)WcT+.LE<AF3ZgZ2#,?9ZGS
+H(7P=/3A4SY#ALX\\9XHf;f6[+TN332DU#?4g3AN3-N][]BK=,MM9;\TSe-].Ud
[:2V18?cO]:IY4M9-8R>][U8.b4U+ZO;D2&M:?<d=1JT<K^G=H&X(QJ,H>(&^KS3
6:;WSe>W_=F#<B=[Q,3P&2W9DZULa?9Fd12U]44eD@_E]SeQNF?6)9e5cO1SaCg+
eNV?,Z2?2AG43]@Q&H.U=3f.a/\bU,c/J]3bfJ.:_a6/616BGNd7BVO(3M5a]H84
>QXP2HL>\=YaeMFf+CMB6DJ=V5#7WMPS#?Sf8[4b^:.b>6gS6c0OW>@d(GM/@P)R
,N=@A8JABBLQAcEc3CE<;BNC]EU1)G2&GUQ(MZ/CL_8:>0)gRB9>?;3=T:dP.6bE
Y<#^Ta8HBD2dKOP@9:c\dJ=Odg_>_KH(aKc@#NbLNag;&JX5>&ZcbBZ(W#cd^Y?#
b4)R)M+\T=QG]YSFANAfKg(]7H,6:O6SdMKSLQ\6OKY\0R-WR@@LJ1,F43/=D3_C
c74^Xg1X6L,#S(B:fXY#>3_^Y5@GSEG2BPJ>H\.L1)US&E1f-IB99:8X.7^aK+9c
VEGCgb@cYYcV)YXDVQI4I9I#Ke^(AH52eJa?)P)21?0&,(6X[@YfJUbXA?J9ZC7-
4<1(7FdbdE),]Q4(=Q(Y#:\gBf;D^PfgfB5UYOKC^<Q+K#CNEOLU4b@U+FMF,8HD
TRfYd/\fE/T6F7=3[8O/@JVBJJ:,\QVF(:2/?UPS<)BR?SHJ+BIA20:DK&:K^8-1
8eb-a][Ga+?MJGN#AR&+fLfWQ?PV@dg\P00c#0Q)=Fb/SBI8/2;d><@GG/^VF-E9
M#@+MD.T&&O(Q7g7@;^d=dJI.OE1E3/@<b/<_A15N4K:]7VAL.W,A9ZQUCLY)(V(
9^B[WMW^f5=D(2bWAJ>+MN./V?,-/(ZC(7]XYg[U#Y3]g<B)0:[F#eA2S&X,Y+aE
;\X6,3FFIXO=Gb+fUH4-bRQ.2KC7GJSF9/[S/B<.c<cXVbM1[)[O54?[D,9(Z[4b
ZYeH.fCKbYaWdL+eDSgGIV6FKE2\Kcb0&^CN2+7.G=].O=YV-/S4E(J=K1PQ&5@[
))c(O7Q^JH,-),POQ<ZJOOeC+NCPJ+C6ID>9FF/1A]4^85YQL-=,XP<D1&NGQ[f;
K^TA#FU+SQ@JPN);>PKQVL:,d>R?3I54S7<Jf+2QOAL6\5+ZcD/^4d6Y_#[Q0///
&g=bN=@V?VfZCaS2\>D,>K:O[8.Mbg_fKO,DCM8A>5Ld\Y8:V1b=eVEfeDbN42\L
N@=b:.6Q6BX,LDRYA(]2bXb7Ub/2.&^2a8R2>bd3?c(^NaH=7E2eF/3SCQM1DS-;
S8G0gLdSL014#CHPA4-N>FF2U;)PX])STdX(a-PYV2IP,DbXLT[]7V=#b7Ie>?FG
)BJ<;VQcY@JL<e-R6<D8U(D3KZb_>R[W:7\8VB)?a?f@bSSWRAKN7VMcODBc#^IH
#IXJJ;dY[VNJ8ET+K)_^</=MY)5U0b5<DgR]A\;;C_VRe)3K@_R\XAPFT69]cX_E
d_?=.f(W#.IAS551&=T1P&HSfFZ7GA1&-ceO_=QMIafLT/fRH4bO2M.&8RM/D<Vd
+4]A_>40-X_C6.46+.^-@IZO.Q2-)3FO[;<Q-)d_PHW^7eW;d_;b,XHM)2;5()gd
]F&0<D(d6IbUcHQ,I9YP:dd9f/J_O#B.WD&[&8;L4O2-RgB05e7X-ad0I85ad^C.
U=W/WH5MM>EWOO<_ZcF0\E3OM,5Q17R]VBB&\E56F/fO6-2=4fF2DTB4J?E/9MW]
VO9cIGOVS.H;CVULI\Q=+Y9UXJCK4WX\#E+cB?b00W+OY<T.JYGXXMFe=D-5L>+J
@0,/7<V[/V?TK7;H&/(O(24a[:\ARd52ZU11)7#F834I6.XW62]N^0XABW<M:B[B
(\<A\1&Qf6W43T3_<RbY.W3@UPOafYFd1Z/WJ3=VgTBe6O=e7@4M-8\G>EE6)X/]
=bNCO#LH\eUXVOVg<YN]+W/HAC[S]_dO,8?C--/H7?^E[T#<AGZ3-d4O-L:S@SdC
U4IaUd+(5Of1V/QRR3;.E\;-<E60g,:_;X8eQ->K42#-WY[f-bRUX\T#<ad;T+=?
3SR^6M7gRKLeK2G#^g&V<-,&6H+088c<KBZI<C:LA7IWY[7>,F1_&Q_N6?3DS2^;
G^/FYB(<[SLNK5-696e^;2<5K:=>/2,PBPP)@D+^D6&@D5IHE97LZM>K+C85\XV3
f[]]XJaVE=_.GT1a=1fU(GMXI8M)F+,#)(64I74R8\:BPf/Lg?d;F&f)S&\-\=c.
701G)0^4\6:-VIDX>aMeZYcANDc[4B,dFK[&8JI_(SJ^O3QWbCLJ0WE1gEX[@OdC
Gfg[52fSV;afDbL8)GOg/GeY\M;JZ/+H+CZg0>5?HbKfW=8Y?MGI)GBe]WO^O>W)
ABM;MUKVQcV/^7>2L:e069J/?-Q1Z5T?<0^3B:ad3JK?8I=c?3M7bf,L^8[9/P9O
EF_LJ^?&>NWb.f9Xc4Y544ZMRA&P)K]bIIQCLK7]FcQaf=gGJW92)L&IBRM,QC7B
YT5867#&FKcC;M6_5PY\(8]BXEW@XaC;ZZJUVH&T>@J03,2X>U#^6LFC(JX3Mg=g
-L:DJ+#f(J)NQ27b>T6[9XbBKTEcPF&=E6_,g9_,I\FU1d^CdXgXML-I-4I&6:J&
@V?,I/f\cEVC;;([GfD90TGUggBV80UI,d,Q_.M4e&61SK8YFRWODC2_U?3@/TVK
gbZ9@a9T0)30O<,gX7NgL[H@-8N0NON?UORcODGc\&ML)K>#S_[cBB2@^#Ab@>^F
MUG]JIIaX+N\NPN);(bcUGPdDWLg0\gH#EUH#QK&[IG&<^eeO4>G/V##+C_Ba]O2
X4QW;#\8V1[FGX5gAZf^d00/Xb)U@=]AA6eg>:(,OT.IW37<+g]Y>@e/?cN&D80I
_(C8:SYe#N3ZASI2Bf&Nd7&K?_]X@4S3QTaZL-00&GeI(=,?-42CJWdI(75YHJA0
?:_&^CJT-4BMN@44a.PI)c;1TcA6gQC>g-]b7eIYA_QQ?F:7-HeQM3V<_(=S]H&U
\#?@,+;\[Ta?Kd8NR+W#cA<6eSV>Q6fQ/W/NGTMY\e[/42g>Gc(F@AYEI-J=e@7(
/db;GOO&RS^:W&:^EcF_F/X5a,aCRbBc&dSR[4Y&#BM?=-J[>GW4A(Qc_1AF1^0(
+^YS?^&Z_GXLT)cZ75\8\-55d[31U:\HL&a^-HXXNgD[CJO]L\[cV[@A-,c(4F\2
gaOC2.9K73]<UO59-H-d8Q)S&QDeBVcT<O=?6:\AR_^ZGMDAP(P^;@^+)L.WH:fD
>J1]+UE,J^>G(3-GVR_CLd7Gdc:fK,DTN;XfY^4B/MfR8d9^-+J&2Gg59S(,-NR.
]c>3;@1X/):XAZDY)4AETJ/5[9OFU-0[E8WMdce^+>P<@f7;P]YMOIa;N)JQ2Q7]
\L62P?=N1EZ>[cW<ge+MCfb_\#\R/<aBXASPMWV4D9]&WE9LD_.\DOaH]OQ:WCb=
+]/3F]UYR:6X:g-5c;U[JG+K:Ca80fH7-A=@N[B@3E4A?-LGB,&@-<A@<QQF@406
:IUA&ZdHEgMUSV]HY4S8a2FY<fPf5a(aREFU1AS&gLUM6/:2XA++aQ2@J89KOX_3
c&?ga0S)>ET,;.gVfRZf3&LPDCMMEY:4<.?6D9(;F)Ybc@gJ#M)5UfCeJX>7+C(Z
8(^PV[R(/_eY+1VJYLQ\HMZ[;A[H(&?J8#2PN/F?ML[L^H;dMLEe<.WV7H.20;a6
K<7d,<@R1OD9).K9G[,Q@18:\BaX;VDQHZD1(F8GFB]HWDHWU/504&Z?:7S&)B-g
N\G3]1:G5I^<AWX<D/CU8G&S\-c5)_OG7HR/H+F+2cPUC<<_K)GQS4)].;3f-f\,
AN:O>:.baT]a)IL0S223G@Ne3?\HNC=8bE4NIZIF+99\#d=_3H,VDQUU>W#CbMH<
6)c]=]b?&b8D9X9;.9D@Ra.HLS0)F3I-C@\H^B=ScVWcP0@35#KPcW98(7FaO@W@
Q3e9Y8?-1.9>@0Jc.I2ZD(MCg11](\?V[)H#<8e7eU>OfcfHTWIO-RR25@Kd9,d1
L(06VE=d15NW+X,V72H1EC\VQbD#R\(-4PBM:[TGGGdS[7]a5K2RfUMa0&d?[YUP
9^5P5W9eA(GU]VCYgg+3,0ONg-T@^ID2^&1G&:OU\[<OU@d4C-aTI>:#\&P/(X7F
S+BgYZ^b[0=510@4gC\a/[H:1HdQgTQWK[-R;/Uc2UO\+R5c<>?^[:W_K((1WdVg
&E7?_J=@I:&6H6X]O7e:-aL@@MAf,XSO@4E@_)=aTdZXOa?+/T.&49U_-5^4ZVDB
d6\[2b&Sf:B]-R]>IfX?U6&TF8JM+W^[?G37GbGf\4\^+XTBG;7=F4.[<R=_6B)B
eU9HFMF(..E#?:6Bd;:c;5>JdZO(W.)67Sg5HcTK,]UP4NS(652XG]J&?NNY32Aa
YZ\0D&14TRE#&PC5);9fcMHY8W6YfO.Lbg6KecC:eVCf:..S1]b-?2/2OCE=GJb2
F,,+A7?-YW;9WR;DNDJE<.+RPQ@R@ZK+_-6D/)cQQ=+6^Q#-9II-DFC?FQ\9?A,_
S[^?PcQX#\cH[R>^<BTS[/\_2A<ge0=eTb9)D2e,Y>@NE>-g8fffP3<^NgNPYSf(
3U6AN9[3:bLfU+B+?.AOA611IA[YV0Y9IILI[AgP=H,:-GV/L]^g#b(X0.O&JQeg
5]CV8.0J.@)YgWF3J<WF5H&c#Pf5A.BRQc#He2c/2,6&91,d_.eS141FRe+]=@#@
/RVJC]aMEeB&&MXc,fMQ/=G4G8ObTJT85gPGeTV?Z04cRS\&,O?:)HS\62OETE1a
XOcfE6CK8Q1>AH9>DN.&75a.475f.E):9J36;=LG07)N,IaTDQ_J\RK2bSI]@-&b
E^BJXJ4D#>/Qd+&geCc8-dN#T/#2ER@_bcSGP5&eA.McV,b8RVHVZ0DG;efdXX@^
(LRVIQ.:_FJ\XfMcG0IJB,O(OHY:I&J9T>L26.KCXe>?dQ]\1Sd5g26YCIgJLQBG
<?+)ZBW?.-e-;PGCb-.CVg3VW2:T[L+>5_D/I0VYZOCFP\9JDE&TX:f4HC28EKF7
^JSN=U@_Q@7S;?E0Zd&ac\QPS(F-<AU1Ef2K/OUR1O0>f4Pb,GRCfA@36MT(d=OB
ZUM)UWZM<Y#4e^U)2Ze,Wd@ZbR1J2[gZV<FO8>C4.Kbb30E2ef(6@;agY,(Y:@HE
7HB-^H<e\4C[_)CAMU:c8,bXBVXM0PNUCL?0O[XR-\#M>GgB_G>KAXLFKOb:M1\=
^a2NfL5YTOPBD;A==886(M,bL78MMEKJ,UZN4:2bJS:^G/eOJ)>EXOUWH.W_/IPB
JUEZ?(7FI;7?OgYUM[8H^M;_ddUSFAL5_I0?_FTBH3B0/8e</-Z842<S6[XYJ6:V
<PJ:bUW7IE^:-Z>@;>ea\aO0&(@KE4MP0_de?021&O7SbcYfV-c&T0df/XBfRI_S
g,P#5O]CVTH<[F01WfW\\afWe\#TeZY&g1-\T([@YS(;SCJH<dOU4GE+&M\QXFM0
46&PD>W,1e:Z5CN8Sf6&RD8,#Ng&e]Q;WfcQXCWg.TO;4F#1N>U]J\PPU9]GJV[:
Ge/e3fL(H0:5f604O^29c>R39\5X7V)N6cUH.@TU=\8.68[0^4,_a9P<(((;a+/]
c58-5BI3X<9L@0T#ORT3))>c/ePfKP=:d,]GUPPSCI;?(RN9)8BMU2C#9NZAQ)5Y
G4/C.RcJ:9=cVAQT_\;7;2Z-=:25PR)[g&?ILPP=<PHY>ge.X#VdV7RHHS=G=b4e
cRD)2EHIJ_Kb5#a>GFB7HG2\deU;4e.=2+7<KF:(#-_C,LZA<AYRT((5N0TY5g][
G^Uc1L3,Ld^)RFfO)(J<,P]PU^X=89=N3)Se_V5T@00^--bDTXM2<J;a2?)3QQ:>
U67a\)eI@\<:#?8QaJ\e+4PQ(Hd@LaFL2^UWX]ba(,#.J/I&-6V94XP\X54/U6]=
YFZfQ03:Q@e[6@E4:b:P4(X185\EMaM_1PR8Ce0@<(O,5)],DLOB;Pg=8eY#TN>L
7BFZ?J7FGaJIS>P@HMRE.TW]e39H,Z54,NNDUTL5GQT^\P]f(&4/T>9<]3aHG(Y#
<(>W<ZBb);V4M<0N,S],,269QM1JKc43&VPK9bW)6]XX9GC=6^XA._)GMEa966)B
^.6>U&7V,X+_+cc0E^>3=25A:#RQPI[gH:,J?fV>5WAAbY]Fd@M)PGIA\R^)HeL]
NK+N798Q+3ESE^2ReFG;B0;+.1B]6/9:9^-P6Q&UgRH@Ma)NL6;X7Fd.gO/?)J97
M8-G:KcS?d67ENXMW(3FQ0&IRG#_cL]G5VL,5&a<14\C[?;)A_^B0NO2&OZD?PO9
MT(I=bgG4L[7PZBd?:aHT4D9c7C#:Y,+2^WgJ&C,(][<#;&MAOB>HI#eOH_S3P(^
,TK)Y:L6=dD<)#dcc)_B9FSeLHU><bJYg>;A3DGI:a0T10\7Ga7G;,4a\0Y5XS?2
HHgPZIM3WLQT005MR@gS5>NET__gE+83-B.6;#T8aTM[>5)62O<QP&d@OI?=4YC>
a=Z-0g0XV+Vf?K0>4HN7FZHL+/43FeU;YPC],R7=S.H&ELb)BSCB+[]>DGbdI7<N
3ge(DB[1QFWYgRgKKSU]B/J3C&9/P<A=eH.)0==Lf:(,L4GWLdZ04@Z^2T?O)Edg
J>+@-)dIU2Wa421?E&Yc(:4Ka,\=LS;\.UG=HZ_dXEIYGMD&DgIPf=#]Z&]LQ7fQ
1CXSF7TP.Y/5\6>K2-E9>ATIO6K:C0gMXWIDQSbC>Y0b/PM;&9>JZ/D^,;QQF)?J
L7fVRY,E=60@B3[+OA^46e_?D=&S8S5_M=bef+,3:E)PNF/]O#@e3PQ?4<f9g^&8
(=XW+.fD;aOI>^RWH^Z)\5L<\O6U+Z3ebc\KbIS,B<A\^(WWIGg=O,[9M:T,AN[<
\,M-PFNJ2e[V8C7;gMZFU2X3KM0M)I,3RYf&aQ,a40)eL-#J.--R8N&?Q[<?RPL/
/ER=2Xa37@_[U,4(a6Tab0-[/[c)be-1\2]>AV,V38.EO:4_MeO@bP:-.fBKVUa4
?Y(:]@O9QTC1,@6_U4SLH6ONSad7FP2B-_<:_K:bd+F=J4LBLH>U+U+aDUK@-O;d
fdNW1,/3HL&c2QQX_T6F[U3V(48LF(G#,PB:CR6F;@AV0Q.0-[2JY#K=K(LdIS:S
b0f&FbELB](G0AXf:f8J-6PXHH<274:_VQ6(XN5R^XBC4/GM8GQ&]C/PZAYD+4(&
)4=<g6-FN#A@0bN96N?Oe)IM1FDd2^0LG=.<:XBD3TP>6=FX;(-:X]=IfE+18XPg
5I<,>G(4b-N]\6KfQ6D_6;HV5H^:f+U?IM)]RO0]g3AY?@ZX:62^#b853.?gL/gA
OGE@2548OL8c-R23dHYf.QCA+L1QG1g[-9JL_9F/e\>f2c,UD4[6GF&a#64O=XaC
[BD)g,8fG1=2779F?V=3V=O9Z3[5eX-+YOeP?Ue8XFfZ?4>[LKSOH^c3gS57IL>K
U&<VB@\G(AX;6a,McP<(UXJ^f;Y+=VXb>?+A/09eJP:_C\^#KOU,A7;(@=(Y8G\_
<PDMdfGKV^.-BWS)a)S&>(=g^aWW\R?OXBP>J-3\K&Q]@H_=KC,^N0<805[HLR5c
M99(:L28NYYO^K[2EJ1/D<^TC1\RT#AN&&:6N#O1GbCaC+V1+;=AH[EY9VJI7S<Y
W5cT?^@Y9U4\^1f0#MRF\S].S,C.Y(E?b;cXPY=4G5E0.SZ4bC&XH[8B-#PW\bWQ
JB(Ka1NXRZHYMM/4e7beP<^89AAMcO@4<0f5Ta-\,HE&L@G:0cCL5TcZ59g,FKWR
d=a+1e,G/+Lg>;4S]<SfNGc5eK>56L.I)]=<:]K44TF/]MTWVJ]M>d_aW880_0Eb
DKU+Ae-EL4HNR(B#0B0[.+7T+[A:]Dd4]a@@22V?gZ9VJ+^dbEe9DO_C1MC#SCXH
dXV:Q?1XDIE;L=^QR:;\R8SWIVQOO3:@XQE?>CS4_U._:>0)=9]D]:fN9NY?7Y>A
SFM).U29d\(H&/M-Ogd@YLXbM[bS#8_FHa^FZ[]=5NWQHPZB@HVAPc@T2ZM+ASWR
7UIP#c[V</1\&1E;PKV;.4be\CcQa=#3+YNJaNW\1C>N<;XN=,eNZW)9&DT5Z-fZ
<>8A>0Nb4MDO4UYd68Q_M(QGZDUM(=JOPdA,/83]^T/1YX8RF(EWeLQZGY<+XIO6
^Df3H]8VP#]2SIX6@B63f8QZ7]bG43B&<=1M.FR8^8=Y79I4T:^=Q@#W#ePTTN5^
aM1XLT(@^@>;Z34J_30&+g=\S4HOXNJ8TQ8cS9OQ-(TCZQ/_HFA[^9a1TDC#DI(D
A=A:VcS:f0P<7BdSJT&ZBH^7\b0_JF3NIVULgY[HG#MD1]-G?_Qab#bQIMXWT?DV
^<QH3fIMXbU&RQ5YEED1L&Q_N,/&3,LED>:-;#I>C3]^V]H(J;:.BbH8<M[U\Xdg
;6/^TR50;+cVJe)/L7)UM&DRVc\;7>:.HZZ-JdTZ9G]V6#C]A:HCV[<>?5V7Vd52
4])?UbTGb]VS18XAc,UPAEVd\]<AK/8/agQPD:JT:^R(BGQBX4cK/B#B;AHH_&VK
C9cMLP#cJIFSNW>c_SD&PJ\?OYaS)QQR:_3XcI3HJMANRLb<ZGOe[[/E9A;CEK(f
_B)WO\A+7YC>2(b]JM61FNPZ13&](<(g.]:66dHH4A[G2NDJEAGaMGL9CBb#F9e[
EG6B9RMa9VfOd=Q_;WJKg9]56(f?V9,KH-A;OX.#d>,H1VMaRMGEDFgfGA2VfBcH
-/&7gF9ZL^&<C]\EaED2H:NgZcMgYM_?\_?2Ngd-U^VdLD+090B=eNID0RV\(9:a
3-9XZ.<BGEM=a.VM7J4W1&_T-YYfP^HF1,O58#@-c2WTK:=?RRPD4cfF]dYCga<,
aF,Jd5AP]8R+;RWO6GgMVK#eK1RS)Y&ELP\)P6Z>XV.847SGJ<W=[bE&@B2):U2Y
E8^Ff5GY]?MC:MA.;5>e4NC^#^(Wg#PQP3WScgSG_+ZS(>#f&eD_LY9b8W\MXP(8
Y#;Xe.K[+S.4X,+b572SZ\F-G9#AP,<(ANc^)T,cf&SVQ+ECV3HLd#MX56R1,=<A
c_EFP+0YS(,KPN@5a?(585\[=5):HIQV9Q@ggdY[9;3fcK>f]Z[^5-48-BW=WOB\
fXU.VB(_+eF:1=QZ>=afb&GS;B&F3LB(A9_M2FM]ZX(fK,R_CIe&]YHc8Q?Z:):@
\H^b\R4E:U@b::[gNL:,3(T]MTNO]NL77[(\XLAJ@:b7:S+4:[&ER0#bbOQPaH9.
;4NcL#Q91Z&bAg/E\;^R&;fSf,::ITa<)e[U5&A@28\[5eY\b18gEZfFD^NFe#gM
^6ZTbS,^+bD@Yb@EKP3Nc3aIX/)\,_a#0eg/Q\08[((abYK];9Z,g3Y5T4B)3aM-
,[R.0^0H5FQDJ6RQ.X=d0@R=4f.UZ6bg.8M9eFc[Ldf)]5AWZ?9dOX^:-E3b56e=
]TdA&\X]C<J7K,&DGVF>]gL.WL<X;R23?\<9<;<O4>.Ea;Rb@2/UIfA.--(P_&78
aMSPL_H?a.H(ROW]29DH-AC,,^CXSfR7H2K.Bg<JU;>/@5A3FJ_S@NL=M54d,@W1
aQF\I30d/fVe_;?@beQDe([93>(+J\gILLEOa(dACM/5S>#AGMHSMLc+_:YfL,]>
Z;cH>a^0S]KTHYBCIA(B0cW0#@LW.)HX3ZB\RRJS8AA-Pc<1QU5NI^=/[>ZYcg6b
1@?.MB9PC6Z;a0FTBOO&DG^J1,MJdJY<_/[0Z_^(L@XU_]Q,a1N9I@#^YLUX\S8Y
-+\J8U-Lc<OYde5>eH/N+CP5^5-]fRHO5egK+59432F5\<CBfHVV\c1YSg5\,K\I
4_F<T]eb3P4))WFNea.;9/9ca[X?DMB5N([O-U6AfYg#^\Z,MSQ?0UM2>(S([0]K
4Y.A,,HM911Z.:K#ca12N<SQN:I^/&4/:2=V@NE:I2MF-GaX#b#fF(gWdgVRNYCJ
S/1gdE\^VVa&BF^554,2[V(+_RE,3PDf.\>Je\8/@Af)=866S/(D83_cI\2HD)2+
5.L@;)N-Tb2=#\Y_1Y=/J/)E/E@RceTXZG=_?9+H\_X/6e)VZS65e8&?2@Od2]N7
04I)<e^^@6EL(LKDgQ-a1TI_RJIZPM&5<[[YcI,Q&ZS[H2fB)RR#^D7CGJES?ga)
W:Gc+N?Y;aRTW=c70=\2dQC)GK]\9[gBC_MN1V#]0_2T:(ScPb17@;F)&)@+@D4O
<4@DW9=I@S(0Q,cV/YDQ>IfN#)1(bE?I<428:-5I<O=#UKQ?-].dX^_I7.1ea>Z1
]-eQ-ADK/0=VCCR<H&Xa5aJ4FZ^D)6&).D.SE.c+ZYWAGTd(XX&LF?=_H&,]]/=^
CH>G0Ce=/EFPE8aW:F+R[g(9O91c[dB/D;cU0Ne#CS;Y\#_1E:7:16_/g@:+@cBX
-7H<2D_B^I9YY(:NGOfcN5=,W=[D(\]ce?3RMBHN?MX:G/A3GQ]0@A4Z7=dJ&@MC
C50=>aD7HI[9,+N.?=Z/A=.8L8X)Z:3[Gg=bdV<XWSR3B9YHZcMT)?#1GfUTY)+B
eddC/22_D@\YTcM,R3b8E#@]aCJCA7/:/)=20+X<cP@7ZRDK2:Z7+VdS-P30)26e
EZ,R)?F1(&=1<A?2SB?SYfU06)+>B@(Sc3IAQ[1=TA?C;gS:<g9,65UQ/0T(R@AO
#B4@NZDd4_2;PNgdX9?SFXQ&HF^<TN02_c<_c&O9<b.I@@C)_\N]<8/Z,Z;)e?f4
^N588XaJ?F_(JFD3b(?BNc7TMX5F@g428_AdOM9D@O&?U-FL@,.Q?&gKJGYGbd?F
Db:^@(>8Sf&+b_>CFQN):\3_U0[Me6IIZ+C2CZ8f[KO+3[37)P:M<eZ8UW=9bNG^
P(,6cR>;&b\QP1cV01OJ1KVWI1M8^KQK,P8U>WX)?;_b\@UQJc@)+M.Z2LPcc[E.
F3Pg#:_#06cRa2<MX>b&=@77SDXS?U7M\TD(TAB4[9E:)K=U4+dX3f9H\80>fWFY
<KP7HbEAVdC^[.K_Z.^EYH7@R_gW[(=+;M:(SaK,Z][dM9JS4a>fBaYO2S\(XUXS
\1\P6a4LKLC53T)+Ja8BL.cc-1^fHbFDJMYR@Q=TOPGT(3X@9-<5[DYEf?5^+,6c
I(H-;X=?)YCO4\S6#FB4f7Z<VP(gIda4G61>ST;+]LP[T@ED=BA5;2Ye^b=#M,Id
&d//GBS(=WICD/N--M:fGB(E+<]HYMfD0bS1XJ_fP\a=V.F&f;2b#0G)IN2(+g8P
W&24VVDD9VCb-5F8F1TTcRYV4^[gY0EPKb11+N9LU=R+;8DJB61W6Ca,bARA#Xb3
]N;0dPdd;RHHAY@6f5V[LU-6:65Bd(7=feE1&[0a_U;JDA]V_^--0aIK8B#UTDX[
B1H8C5XD,73N4#O5a7RF3#;E8MYO&9\9cKBOE#HE)+K:ePJ-#Ag5RFYX^<)e+2d9
8>,X.UfSTPMbW,6M5A+&?>B5PKSR:GY&(H5H;(@E\/OVeQZB1Q,X>YC-=e[7Y7d<
6]bHT0A4F4EJ+:c<#7)FcM&7[S,e>9UPWW\X&@-+@L1E\AP^3CZ[JQb2L:P_NEN&
&KA)<,Ig&c,f^e&L9a0[g[4FIHL0N)SEd\Ica\BI_LL)(Ob^;@<-g8(@&10&JJ[e
-SB#Y#<^>(+YKd@2-/LO=\f6e9[@:+_EAQb-gcAFERV@-FZ<[GF8MBS+G-8bWI2]
\G317d;fBBP=1PTY<5e.7XTJgMJ?VGSe^eK=2\S]@Z-))2\eD7D,/\LGX=LHaV8S
U7]-X_+38Q;LK55\2F?CRMF=AZ&O_WKY/-3d\.#R;[;ec^c0^42Z2]^IZUc+VZa(
&H=N@VIXgKg=MU;cYRa@Z[UK^Z:b\NE[?NAd;OSYL\cY.-BSCDT;Vd\#;@LH9Y\S
<(9bZ1R;G0)UVHKC+PNaf]a#SA]5[b9dZfB^S&E8,L]9&V-29XRDZFR-L>-:?>R0
S>\5#.D8:LSTLH8R[.?EaVc7a_X#_88.@RMZ6.+B]F42.@YDc\I,8_EOVB7b2fC8
eMU?@>TQ0e7Ka+5K3)\VD&+1U,b5ISCBHG]+H(BN-N=[[c4[(Fg;OE_d18S]RC,]
K.e17aVKN8YOKD[Y7J^OMZO\G:HegRfEVRf>A=4PABdIdg.N68XXQG/6V?5gaaM_
F_GGO=L2gIGX#4e/bH)1Q3a#ZMBOE/8Za0I:>0);;VOS_O>_SY@S[\EebCJ>g=KB
>R<P?F,A/=G6fX]_A7IP_JNC<gC<UdY[(5[Y_LYK1W3A>XY<>_cU:?\-6I\P5GCG
Obf?K?]2=d=[9FH1(N)UP:>P>fHA^1aX0NT<D:<d6D@Tc)9/CP+V^6PWML@L]31W
^138F?\0]:Kd>]e1:Uc^S=3R(S[Wd4c;8-OVELeNHQ,9bY?dP;O4F99;4^S5G:;;
A:HHB-\@+]^JbS/cOg#NUc_>\:+:cga_M#L9bZZG,D^.g\Ba9,Y^O=Z,6BH,2CDA
a3bZM@CF]0dC+IS2YI5bS/(_::<KJ;g_11U#KLcAUATDLbb;HX:[GNRHVdA9ADIR
4_#]4bB2N])9-/13d0+S(BDZ#R9.3\D.AQ^ND_2D8VHQFKGeWRG_)7eO_:N,<.F>
F>79BQ<_eVHaM.5@d[#8<Z[eOgIdOfF^dTS=&MRDP#12\eV.9B(O01S0@2@I9Z_+
YPb<1LMCJ9^Z6fb[\G\LT=BFVRQ<X8g9H?)V7_XeHbc.Y6<gJ^F)TQ8HP8Y-)FfZ
bXZM>D\5D:8V,dKFM80gV4[9<DXH,58#2=PbE:aa23O;^a7)\RMY8/V3-W3IA:&?
[]Qe^6H3aBaS/aC+[>4T9C1g]S#WHY<=^KT>?F#Y?)^f\#4EFdfG\1#cfWMZCV&R
)\X8(8E)MODf#?H40\[=fAMeH1WL#c214-@]?9-=YVZ:RJ4;JZ9ecYAZ5BMOQD3/
SW[fGbNJ15^Y.<RJ#QY/>47Z[5\N)N&fJ?/Z4eg7M6\@6cN&.WO^^Wd72G-&+>2C
ANF_?8N=Z7)0<O>3SA#3.IYDdPeD/EYde]aIYTA^LWRD;H3QV3I:0.9Q8f@,Ue2A
X=RUL#O(FBAQ<WfJ[E+8[XcP(&+cS;Dc3IFT71Q;\Y=C=\=MO7T[-3P057&^=MQQ
OUgQ@&6W&JEg10PT+DP7)18JY]DI90f8-UVc6aRTSe3c-9,M;I+JN]L54W8YKN3E
.0X<HSR,H+3HZ]#d]c]]?JFgU5ONZ)BC@96IGd5F7gc^9WN#2Y62aWD]2Q#S2:5T
E@0AT&Ice.e9_C,:WMXa&5dFH;97O)MFY=+AcW6&572UgH6&6()3-7J09\LYJX:N
=:[:7aPYU.GPUIC^7,U;,+PK#_/@MV<_P^?^/XR/:KK#Q;\M2X;],\D&UdPa9NN1
S\3QF4SFLXQdg:SOTZ0/#1\ZBNXJ7UX\c7#54G6S\0+ANLe0U4a>Of)bGGf[-M,B
AHfEae2K]?U]:Gg9GJ01+B1K,@Rc(-gDN9BS3+9B^I3<GAP(Y8+AJ\MASMDK74@\
R6B_cMN6&<Q55>09,g1F:C0J9X?92A^QFXT[d+:bK+CY9.>\B\Yd(^.eE8+-M\F7
Q,T3PF[adM:SX:<4BDL^=2^c?-\03B7-:gX>R#K9Yd@e)YL@<Dg:PFV7#\6aO@8]
PBE-,E;ML>J;bW1=L:+-M+[#7,\M0gc2[4eL?/0F=ddVTC[MWLR+1X._Cf2QfL/-
7TKM<f9dYZD8DJC1W#\/]e>;LNU\+I@RQeK1#af;)P\&I=E;\+8#N__LH#MZ;R6.
WKH?e8T8DM,M@@9(@Tg>5Z?^&=bAK+D\Z4&T<.aC;HLCMNXBKTK1VAAU_D_E<9ZM
I>&I6Id@GDNL?(6(@LcTZOY9bU<S_JDYJBF2eF1ELRXFP,4A?O\d]/X7ACW#?@O/
ZU44?8F;#12+ZA^JSBA8538UI[;((ZM^)ZYJI9OLER\a4(>fH0+P<f<VV5M;:/76
C5W&cJYLA=OL7^=DH=]EA_[d#Pg[DR(52eAY&BB(O5cg>Cg\TKO1Z_C=PK^#O;9+
X&T7P/SY;=.2,=G-R_QA_#\)2LUQa?X]Wg);VcE(OSMg7EE=9(W4^<<FMU6?+[6M
[M=-QU?<Sg,CQIA(5@49\H&>SXS8D7V6)Y7]RI+.aJ-#_4[YU4K;_aaK@5FE3E=-
][T)4/5,dKaPY7,WU/Q(GE)DF(WbI^6;_(F8D:=(4LHVV^X-aG</b0Hd-M=EJ&HM
cdV-[J&>cEM)Y>RaSGe<3\A,V8.JHBQ7a>,Y8.Y8(\S=,#?&<&>0/dY:_We2?Y\a
dWFXN@g3CdOU4+RZ@-G00\E9_[g0-aYXb+:23ZZTS>PH[f69K\U?VZ7_XeTS^AF;
e-Nbd7:WcE7KMc,8XN3Md8ZA9e1?F&g^>FV\1A9H:@5N6?]NK)#gBRNC.ERP0YT:
+Y3>2cfCH1g(bb:G.F92Ib3G/;G0;3#ggAa:&?6PHg7WYJ3d,BOZJA><KS#3=/Jd
LgY.(NgB_XVR(YDeK2^7>)2cE\f])KN#>VgOR3RKW<TWR.(9L^<8@UQgOCQOKHTK
7MS6L0J;Y9(\>dg\QdfN-#SD+_H@?:W^/9&.B_T/0O^7M?>A1;^[V8APT6[&;(eS
I>L?@B57X7_I)FJ;SaQYI^,CNH0c<6fcF9A1^&C_35M2SL:0IP9LC6C1eFc>BJJ\
)]9Sg&3UVE&OC?X(F;,OWfI,<D)]S&Z/XW/D2C4b4/6A3A1I3CAVc4U=aLZgB#N:
CXG#)E=Z/NV0MX^_eDK[6Fc6UZF6\1N2(dH:/FVPFBGM9)NC,_]e7gN:E#<;eO^c
f8R9NGD0[(C&9AYTba_[ZD&M)@^H)F</_QbM-(7FAS+GJ<J\RR@K?OG<5XV1cL1;
,><fC5.HVg:\V4A>S]&GNUE0KSQUQU=WWI]HSJea>UK:OS#=V^a12SV;X0B@CgYY
F53XBH/V.>W>LQ^?3^;[=,-0R@7<]6,bRLf+28&PAe#NSD58Y3TH)^A;XGMXD3bK
4:7XVc;&HA2WK(LZD4@MNegSGU.\JH@[Y>#LbV[UDG&TWC&2f\DagN80g2?6^(2c
g]+KF7].f>#Z(bCG9J[b__HT:>g1=AB?UAFU/Ze&HT/f,Bb7[)7b0XM4R;DX-T#[
C644Zc/ZZMa@GY?dBd.8U4RR+-IRgG]+<:5GXUH]XV_.HNR;IR-Dc6\@L80HZFQH
JM^Xf^U:f[^A[IQgf3R3FPc7T]e/:P+JI9a5W],0?84.-)&IBX_KV5./=MBHFJ;U
L)VQgc@LZc>/XOI;O.3fO+I5d.U1\>7C>E9:K056]R.-V/AT)@1K_I6I[+6IBEG^
4FfMaPVIJ4WdV\/:70FV1\2+[ZeG61(Q_A3gTBY([S?3E7=SQbJJ__GSd\Ibb12I
QP)=.E9M4d&[H7eS7JcP>/Dd-KUGC<f^d@L,B?[eV).0RFCgE[.>IWEB/1W:LC7D
a,SEM7,e),^42QVa\bP.:CR[>G10S>#P>>W;5B&)3d1OU9BK(PeZL@[0TN0f9A@b
GbZZZ9#Y4Pa;AEeSeYG@JFVEaL7I,b>6bd::;T75+NS_&6\bgD16deR(VTXg\W?O
]c[#H8(4dCEAHTA?\X,5a2LT#Kcd]M_9fQ7&7&_/+67811WRUb8cFdd^(D1c6IHf
-3PXD<I4GP?TG2#feOGE033DTN?;:_Y4)Jeg=gD6+cQM#U])G]^7C9.fH8L\(680
cd)59a#IILE/^ZF6MXRCSb[R135]9c=WR=8DA@b_<ZC3[@[-S;9d27+/7b\gK>2S
^,EAUO>^?JF@\LCf9f.C,.O7(L@L8H\d2X43XCe[UD\MC@(g<DZR&IW+/R,b8IS)
QCE\Pf)FD/5MY91MP;cA;CD+PP<RZUI&0a9N-[<a/IKZ2CDdI.Gb,TfG+^b_0)<W
aTd0fN8=Eg^9#BIf,IH?L5+O->5E-ZcD:LWb5[/A<[Ve+9:3L121&ZZ]2YaA@LKL
^H^XWJEH@VQcN;ALA<FaJc02dc7c48Q48S+UCK>D<AQ<dW^B(:Y^.3>)W3a>,+A3
3@Z50;8,.@NS)Oe3Ma;OgBXAcT^-aMZ&QU2T,P_+8CQ.5C5I+T5/d9QZ4ZQ1a8aD
JOedbIC;CZUb9bI-H?/3JXNg]MW92&dCY],2U@6Z-;7_O-@5P6Z4V:NHC8/)F86+
&KQO2VF@/\,,f]3U4dX_2c.Pa#A)<\&TW^):>Q868C,T@(50Z9TY25SRH5TW+1/f
5GQc?eK6&Vb#Z@W(&S;P-^Wf_afFI=7I]5bRf34N=Mg8?aBEIAIWKa8/8T>d(P9g
JECN+0B8LdP?FWb;DVM:c5(7/L]L7Y_>..,P:YX3N-T152f1dH[;8T(P0B]SRGON
?\O^@2<fW-4T#[L_G#ZBF_:#gTM+D9W\7]J1T.Q>9F7?LFQMF@a:f//=0B>Sb3C=
;Z]88?SI?3(:80OaFbA/?bCb,d#2.EBA(?3g\0:(B<A0D(7&:Ddfg7f#4UC1E=.@
D/G^8@)CRM7-@37S>U8+&P4BIEIa,W)FdJ:eRTJNc2;ICMV\\WB(Z;?H[0>\C9EW
V&QBP.]Y1D<5_.0)-W4=7-)W=30b7^I,fHIL4_BC47dT1)fSF7):712]V4_MA>&c
3HFQ]Q?9I7):FV#KD0fNDLe+=aO^gSY)U^[_KIR#KSCREHL7DJ6_J3d1BYH<EAaG
6UE>C2SR,XJF-T(/g0H#+5bZ,<KYX>9R,_Z-N&T\,0T8T6LC2)9#;R-/#QZ0KDNP
:8\I4D0LLT?8/fgK<WDBO3K+4@W>Y]<3=[1&[?:)dWZN&6O=4T_5XK\@2GU<6aQL
DRXJ(>V1);)779TS>4Pd6Z9a^g+?_T<Ja1)9bJg11/T9V/?OVLDXb\7(#g/IPM/0
f/UMc&]^2-ZU-IfQ6QbER.N0LZKUP-I+>Q>C8X2ZcF=LeN/CFT)I(LORTR7<+A_7
),_c<OKd(5Yf=bW7S_SV4bK[)Kc6d>^+AU<-dV3V:,KceGL]g5NA--=JO_K><B?3
3CK)-J1+@V>(bLJ8@&74V8++Q;dS9<3C2R=Ae(+A>\:#18J[4f_7YGMTH?6YM5c9
C,[2-SffO3DMKB:c8XEMSEK+11YL&)E1TM2c=C)^,G7.;fAc?W>J8E\eL#d^Tb.D
>[LLfIc8RT?(^(B9G)eZcP1NYUFH#XEf9#8f?Q[K,5_<.MJ^V:7\F#=.EXOScEX+
MD>7WeIZG]PXQ6(Y.gQW6Q&Z]PO28V.ZS@5DSHJ33JATBI0(H\XR+9U3/g--S_MG
@ReK#:I=d6#,^D3(e0YgRW-6N3EFTV;K2^e7_(VI_5G5f[V;F^KK_)ZL3&#Q4B5?
aAMd1O=b@-SJ?WT+7H>_T#g2W^-gQb#8R=H.c9UK\(^OdHYg7A<6c<X=_;[R&.U[
&8C:(/<TB:]Bc04aR#2OF)aP4BA&G^+e&bRL(&^dQ,-FW/D;CQ3<]ae[#aETHG[.
dH4\6aV&/ZSdceSeBVY16/0#;2XN+GKMS+FK8_0#=a.=be?8>FWE0;SV(&P59-JU
6=fAHZX@gMgJ6JU>_Ze1I5+?XB<RCGW/F.1U;-&8OT-C+HOBAVK]/gO(31_1[#bd
Qg1,G2IPP-6LIeDOYPeH3&0a(W6&H@\R>2UKdDdeOJ&fRLPZ&DPc9I<RQ1&.TT9#
JB309O^I]FMb&C,Q.T[XU^15B^Y6U9.W?4XWAUaGN^/P&MD>&GU3cC=I&c(0(MC8
N,H(S(H3\\+7Y.ZXdbMDg3]Y9^RebG5RZQ60T/]4\B3SMNSd>YWODX_,Zd7BTO&^
7SL\^H6\#P>&+KU18^?6;g;AbI]C&^PWZ5#AHP.Kb\J.RFCMY>8ULaQT]:^/cC(T
\VbebKS6T5;\TPb):7AHPYGcDOb+/-1E+NX(O?BWYJeB^DFBd5O3#G/H0:^OQIDL
5GQN;^-V7VbQ4NGP5G1KN5X;[/;6X4,A0IQ;0R^SJ3fQ&PV7FL0N]e7RgS-O]D6;
7R[a[aH,Y/QMPc#]3VX1\FJ)[e<G=d?+)^e2BMaPJ@_K;]R<gHd6MZ.&,/I7L6<7
U8gD79Q=>FEe7>f2G@PLCW.B?g?>^_OfC62P@GFAKGKPd6K]XU6G&D9K5/dUFL4^
M1[cW?F1@116^U-7Jde^89FfYAbHEA@10MBL]@\IbU.AI&PP)RK@SK\GNWTA_^cM
MG7fgQgO82<D=2G592^X7Z>8gCH#Q>fRM\V+PW.+<T/DJK:.@MGa2ANHFU1-3CE_
WUS/L77\H/aYIG6e^TY7RJcH&<NIBI/b:^=cc^V(e.;&BKG=C4,\,34JZC55I,3O
EXJ:Y:UX(RW#J],A8R)Da2ACQNS=YS/>eQ>B<0&Sf.6)5@X[,;5\b:XU_H+:5M+O
C_LBFSW;Y&a-/5U/G)8H7M8:6gZG\\0OJ<RQ4Ga133822K5aeKa13_P+7RU&5YYg
_AgZN961H>;A)Dg_b0P.,9EV1NTFLW8^X4g/2A.eK[Vf@?8B+SFd.[KbAW5NGW^M
(PD<:337L)=dOFUWKDTAGLgge/NFM?U.DZ0cQBFM<F#YLNR@9e9&eb,W#7CO4:7?
E5]BF.<cC[AP-;RD9WB8P..OHV_b7M4=TI,L2<:HJEP]@\Mc2\F++>74H5_=4I)M
DJd2WRW-3-IELI5N<&TVWRP2&B/B]e3+,f8N>1UM#_Gb]a^NOL:N[/74M$
`endprotected


`endif
