

`ifndef GUARD_SVT_AXI_TRANSACTION_SV
`define GUARD_SVT_AXI_TRANSACTION_SV

`include "svt_axi_defines.svi"

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
`define SVT_AXI_INTERFACE_TYPE axi_interface_type
`else
`define SVT_AXI_INTERFACE_TYPE port_cfg.axi_interface_type
`endif

`ifndef __SVDOC__
typedef class svt_axi_transaction_exception_list;
typedef class svt_axi_transaction_exception;
`endif
typedef class svt_axi_barrier_pair_transaction;

/*
`define SVT_AXI_COHERENT_READ \
(xact_type == COHERENT) && \
( \
  (coherent_xact_type == READNOSNOOP) || \
  (coherent_xact_type == READONCE) || \
  (coherent_xact_type == READSHARED) || \
  (coherent_xact_type == READCLEAN) || \
  (coherent_xact_type == READNOTSHAREDDIRTY) || \
  (coherent_xact_type == READUNIQUE) || \
  (coherent_xact_type == CLEANUNIQUE) || 
  (coherent_xact_type == MAKEUNIQUE) || \
  (coherent_xact_type == CLEANSHARED) || \
  (coherent_xact_type == CLEANINVALID) || \
  (coherent_xact_type == MAKEINVALID) || \
  (coherent_xact_type == DVMCOMPLETE) || \
  (coherent_xact_type == DVMMESSAGE) || \
  (coherent_xact_type == READBARRIER) \
)

`define SVT_AXI_COHERENT_WRITE \
(xact_type == COHERENT) && \
( \
  (coherent_xact_type == WRITENOSNOOP) || \
  (coherent_xact_type == WRITEUNIQUE) || \
  (coherent_xact_type == WRITELINEUNIQUE) || \
  (coherent_xact_type == WRITEBACK) || \
  (coherent_xact_type == WRITECLEAN) || \
  (coherent_xact_type == WRITEBARRIER) || \
  (coherent_xact_type == EVICT) || \
  (coherent_xact_type == WRITEEVICT) \
)
*/

// Transactions which always have 1 beat even if
// burst_length indicates cache line size.
`define SVT_AXI_COHERENT_READ_1_BEAT \
(xact_type == COHERENT) && \
( \
  (coherent_xact_type == CLEANUNIQUE) || \
  (coherent_xact_type == MAKEUNIQUE) || \
  (coherent_xact_type == CLEANSHARED) || \
  (coherent_xact_type == CLEANINVALID) || \
  (coherent_xact_type == CLEANSHAREDPERSIST) || \
  (coherent_xact_type == MAKEINVALID) \
)

`ifdef SVT_UVM_ENABLE_FGP
class svt_axi_thread_specific_svt_pattern_data;
    svt_pattern_data pttrn_contents[$];
    svt_pattern_data port_cfg_exists_pd;
endclass
`endif

/**
    This is the base transaction type which contains all the physical
    attributes of the transaction like address, data, burst type, burst length,
    etc. It also provides the timing information of the transaction to the
    master & slave transactors, that is, delays for valid and ready signals
    with respect to some reference events. 
    
    The svt_axi_transaction also contains a handle to configuration object of
    type #svt_axi_port_configuration, which provides the configuration of the
    port on which this transaction would be applied. The port configuration is
    used during randomizing the transaction.
 */
class svt_axi_transaction extends `SVT_TRANSACTION_TYPE;

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_axi_transaction)
`endif

  /**
    @grouphdr axi3_protocol AXI3 protocol attributes
    This group contains attributes which are relevant to AXI3 protocol.
    */

  /**
    @grouphdr axi4_protocol AXI4 protocol attributes
    This group contains attributes specific to AXI4 protocol. Please also refer to group @groupref axi3_protocol for AXI3 protocol attributes.
    */

  /**
    @grouphdr axi3_4_delays AXI3 and AXI4 delay attributes
    This group contains attributes which can be used to control delays in AXI3 and AXI4 signals.
    */

  /**
    @grouphdr axi3_4_status AXI3 and AXI4 transaction status attributes
    This group contains attributes which report the status of AXI3 and AXI4 transaction.
    */

  /**
    @grouphdr axi3_4_ace_timing Timing and cycle information
    This group contains attributes which report the Timing and
    cycle information for Valid and Ready signals. These attributes are
    relevant to AXI3, AXI4 and ACE protocols.
    */

  /**
   * @groupname axi5_protocol protocol attributes
    This group contains attributes which are relevant to AXI5 protocol.
    As of now read data chunking and unique id identifier is added.
   */

  /**
    @grouphdr out_of_order Out Of Order transaction attributes
    This group contains attributes used to generate out of order transactions. These attributes are
    relevant to AXI3, AXI4 and ACE protocols.
    */

  /**
    @grouphdr interleaving Interleaved transaction attributes
    This group contains attributes used to generate interleaved transactions. These attributes are
    relevant to AXI3, AXI4 and ACE protocols.
    */

  /**
    @grouphdr ace_protocol ACE protocol attributes
    This group contains attributes which are relevant to ACE protocol. Please also refer to group @groupref axi3_protocol for AXI3 protocol attributes.
    */

  /**
    @grouphdr ace_delays ACE delay attributes
    This group contains members which can be used to control delays in ACE signals. Please also refer to group @groupref axi3_4_delays for AXI3 and AXI4 delay attributes.
    */

  /**
    @grouphdr ace_status ACE transaction status attributes
    This group contains attributes which report the status of ACE transaction. Please also refer to group @groupref axi3_4_status for AXI3 and AXI4 transaction status attributes.
    */

  /**
    @grouphdr ace_l3_cache ACE L3 Cache related attributes
    This group contains attributes which are relevant to L3 Cache usage under ACE protocol. This is applicable only when l3_cache_enable is set to '1' in system_configuration.
    */

  /**
    @grouphdr ace5_protocol ACE protocol attributes
    This group contains attributes which are relevant to ACE5 protocol.
    */

  /**
    @grouphdr axi4_stream_protocol AXI4 Stream protocol attributes
    This group contains attributes which represent AXI4 Stream protocol transaction fields.
    */

  /**
    @grouphdr axi4_stream_delays AXI4 Stream delay attributes
    This group contains attributes which can be used to control delays in AXI4 Stream signals.
    */

  /**
    @grouphdr axi_misc Miscellaneous attributes
    This group contains miscellaneous attributes which do not fall under any of the categories above.
    */
  // ****************************************************************************
  // Enumerated Types
  // ****************************************************************************

  /**
   * Enum to represent transfer sizes
   */
  typedef enum bit [3:0] {
    BURST_SIZE_8BIT    = `SVT_AXI_TRANSACTION_BURST_SIZE_8,
    BURST_SIZE_16BIT   = `SVT_AXI_TRANSACTION_BURST_SIZE_16,
    BURST_SIZE_32BIT   = `SVT_AXI_TRANSACTION_BURST_SIZE_32,
    BURST_SIZE_64BIT   = `SVT_AXI_TRANSACTION_BURST_SIZE_64,
    BURST_SIZE_128BIT  = `SVT_AXI_TRANSACTION_BURST_SIZE_128,
    BURST_SIZE_256BIT  = `SVT_AXI_TRANSACTION_BURST_SIZE_256,
    BURST_SIZE_512BIT  = `SVT_AXI_TRANSACTION_BURST_SIZE_512,
    BURST_SIZE_1024BIT = `SVT_AXI_TRANSACTION_BURST_SIZE_1024,
    BURST_SIZE_2048BIT = `SVT_AXI_TRANSACTION_BURST_SIZE_2048
  } burst_size_enum;

  /**
   * Enum to represent burst type in a transaction
   */
  typedef enum bit[1:0]{
    FIXED = `SVT_AXI_TRANSACTION_BURST_FIXED,
    INCR =  `SVT_AXI_TRANSACTION_BURST_INCR,
    WRAP =  `SVT_AXI_TRANSACTION_BURST_WRAP
  } burst_type_enum;

  /**
   *  Enum to represent transaction type
   *  NOTE: IDLE value is currently reserved. Currently not used.
   *  Note: ATOMIC value is used for atomic transactions.
   *  Note: READ_WRITE value is used to represent transmitted_channel for ATOMICLOAD, ATOMICSWAP and ATOMICCOMPARE transactions.
   */
  typedef enum bit [2:0]{
    READ      = `SVT_AXI_TRANSACTION_TYPE_READ,
    WRITE     = `SVT_AXI_TRANSACTION_TYPE_WRITE,
    IDLE      = `SVT_AXI_TRANSACTION_TYPE_IDLE,
    COHERENT  = `SVT_AXI_TRANSACTION_TYPE_COHERENT,
    DATA_STREAM  = `SVT_AXI_TRANSACTION_DATA_STREAM
`ifdef SVT_ACE5_ENABLE
    ,ATOMIC   = `SVT_AXI_TRANSACTION_TYPE_ATOMIC,  /**<: ATOMICSTORE, ATOMICLOAD, ATOMICSWAP, ATOMICCOMPARE */
    READ_WRITE = `SVT_AXI_TRANSACTION_TYPE_READ_WRITE  
`endif
  } xact_type_enum;

  /**
   * Enum to represent phase type in a transaction
   */
  typedef enum bit [2:0]{
    WR_ADDR  = `SVT_AXI_PHASE_TYPE_WR_ADDR,
    WR_DATA  = `SVT_AXI_PHASE_TYPE_WR_DATA,
    WR_RESP  = `SVT_AXI_PHASE_TYPE_WR_RESP,
    RD_ADDR  = `SVT_AXI_PHASE_TYPE_RD_ADDR,
    RD_DATA  = `SVT_AXI_PHASE_TYPE_RD_DATA
  } phase_type_enum;

  /**
   * Enum to represent the coherent transaction type. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  typedef enum {
    READNOSNOOP          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READNOSNOOP,
    READONCE             = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READONCE,
    READSHARED           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READSHARED,
    READCLEAN            = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READCLEAN,
    READNOTSHAREDDIRTY   = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READNOTSHAREDDIRTY,
    READUNIQUE           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READUNIQUE,
    CLEANUNIQUE          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CLEANUNIQUE,
    MAKEUNIQUE           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_MAKEUNIQUE,
    CLEANSHARED          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CLEANSHARED,
    CLEANINVALID         = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CLEANINVALID,
    MAKEINVALID          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_MAKEINVALID,
    DVMCOMPLETE          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_DVMCOMPLETE,
    DVMMESSAGE           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_DVMMESSAGE,
    READBARRIER          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READBARRIER,
    WRITENOSNOOP         = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITENOSNOOP,
    WRITEUNIQUE          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEUNIQUE,
    WRITELINEUNIQUE      = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITELINEUNIQUE,
    WRITECLEAN           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITECLEAN,
    WRITEBACK            = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEBACK,
    EVICT                = `SVT_AXI_COHERENT_TRANSACTION_TYPE_EVICT,
    WRITEBARRIER         = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEBARRIER,
    WRITEEVICT           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEEVICT,
    CLEANSHAREDPERSIST   = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CLEANSHAREDPERSIST,
    READONCECLEANINVALID = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READONCECLEANINVALID,
    READONCEMAKEINVALID = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READONCEMAKEINVALID
    `ifdef SVT_AXI_CUSTNV_ENV
    , CUSTNV_L3PREFETCH   = `SVT_AXI_CUSTNV_L3PREFETCH
    `endif
`ifdef SVT_ACE5_ENABLE   
    ,WRITEUNIQUEPTLSTASH    = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEUNIQUEPTLSTASH, 
    WRITEUNIQUEFULLSTASH   = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEUNIQUEFULLSTASH,
    STASHONCESHARED        = `SVT_AXI_COHERENT_TRANSACTION_TYPE_STASHONCESHARED,
    STASHONCEUNIQUE        = `SVT_AXI_COHERENT_TRANSACTION_TYPE_STASHONCEUNIQUE,
    STASHTRANSLATION       = `SVT_AXI_COHERENT_TRANSACTION_TYPE_STASHTRANSLATION,
    CMO                    = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CMO,
    WRITEPTLCMO            = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEPTL_CMO,
    WRITEFULLCMO           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEFULL_CMO
`endif
  } coherent_xact_type_enum;

`ifdef SVT_ACE5_ENABLE
  typedef enum {
   CLEANINVALID_ON_WRITE = `SVT_AXI_CMO_CLEANINVALID_ON_WRITE,
   CLEANSHARED_ON_WRITE = `SVT_AXI_CMO_CLEANSHARED_ON_WRITE,
   CLEANSHAREDPERSIST_ON_WRITE = `SVT_AXI_CMO_CLEANSHAREDPERSIST_ON_WRITE,
   CLEANSHAREDDEEPPERSIST_ON_WRITE = `SVT_AXI_CMO_CLEANSHAREDDEEPPERSIST_ON_WRITE
  } cmo_on_write_xact_type_enum;

typedef enum {
  WRITENOSNPFULL_CLEANSHARED = `SVT_AXI_WRITENOSNPFULL_CLEANSHARED_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPFULL_CLEANINVALID = `SVT_AXI_WRITENOSNPFULL_CLEANINVALID_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPFULL_CLEANSHAREDPERSIST= `SVT_AXI_WRITENOSNPFULL_CLEANSHAREDPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPFULL_CLEANSHAREDDEEPPERSIST= `SVT_AXI_WRITENOSNPFULL_CLEANSHAREDDEEPPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPPTL_CLEANSHARED= `SVT_AXI_WRITENOSNPPTL_CLEANSHARED_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPPTL_CLEANINVALID= `SVT_AXI_WRITENOSNPPTL_CLEANINVALID_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPPTL_CLEANSHAREDPERSIST= `SVT_AXI_WRITENOSNPPTL_CLEANSHAREDPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPPTL_CLEANSHAREDDEEPPERSIST= `SVT_AXI_WRITENOSNPPTL_CLEANSHAREDDEEPPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEFULL_CLEANSHARED= `SVT_AXI_WRITEUNIQUEULL_CLEANSHARED_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEFULL_CLEANINVALID= `SVT_AXI_WRITEUNIQUEFULL_CLEANINVALID_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEFULL_CLEANSHAREDPERSIST= `SVT_AXI_WRITEUNIQUEFULL_CLEANSHAREDPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEFULL_CLEANSHAREDDEEPPERSIST= `SVT_AXI_WRITEUNIQUEFULL_CLEANSHAREDDEEPPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEPTL_CLEANSHARED= `SVT_AXI_WRITEUNIQUEPTL_CLEANSHARED_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEPTL_CLEANINVALID= `SVT_AXI_WRITEUNIQUEPTL_CLEANINVALID_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEPTL_CLEANSHAREDPERSIST= `SVT_AXI_WRITEUNIQUEPTL_CLEANSHAREDPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEPTL_CLEANSHAREDDEEPPERSIST= `SVT_AXI_WRITEUNIQUEPTL_CLEANSHAREDDEEPPERSIST_WRITE_WITH_CMO_XACT_TYPE
  } write_with_cmo_xact_type_enum;
`endif

  typedef enum bit[2:0] {
    BYTE_STREAM = `SVT_AXI_STREAM_TYPE_BYTE_STREAM,
    CONTINUOUS_ALIGNED_STREAM = `SVT_AXI_STREAM_TYPE_CONTINUOUS_ALIGNED_STREAM,
    CONTINUOUS_UNALIGNED_STREAM = `SVT_AXI_STREAM_TYPE_CONTINUOUS_UNALIGNED_STREAM,
    SPARSE_STREAM = `SVT_AXI_STREAM_TYPE_SPARSE_STREAM,
    USER_STREAM = `SVT_AXI_STREAM_TYPE_USER_STREAM
  } stream_xact_type_enum;

`ifdef SVT_ACE5_ENABLE
  /** Defines the atomic transaction type */
  typedef enum bit[2:0]
    {
     NON_ATOMIC = `SVT_AXI_ATOMIC_TYPE_NON_ATOMIC,   /**<: Value that corresponds to non-atomic transaction type */
     STORE      = `SVT_AXI_ATOMIC_TYPE_STORE,     /**<: xact_type corresponds to one of the Atomic load operations */
     LOAD       = `SVT_AXI_ATOMIC_TYPE_LOAD,    /**<: xact_type corresponds to one of the Atomic store operations */
     SWAP       = `SVT_AXI_ATOMIC_TYPE_SWAP,     /**<: xact_type corresponds to Atomic swap operation */
     COMPARE    = `SVT_AXI_ATOMIC_TYPE_COMPARE   /**<: xact_type corresponds to the Atomic compare operation */
  } atomic_transaction_type_enum;

 typedef enum bit[4:0]
  {
   ATOMICSTORE_ADD        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_ADD,     /**<Atomic transactions AtomicStore Add */
   ATOMICSTORE_CLR        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_CLR,     /**<Atomic transactions AtomicStore Clr */
   ATOMICSTORE_EOR        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_EOR,     /**<Atomic transactions AtomicStore Eor */
   ATOMICSTORE_SET        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_SET,     /**<Atomic transactions AtomicStore Set */
   ATOMICSTORE_SMAX       = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_SMAX,    /**<Atomic transactions AtomicStore Smax */
   ATOMICSTORE_SMIN       = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_SMIN,    /**<Atomic transactions AtomicStore Smin */
   ATOMICSTORE_UMAX       = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_UMAX,    /**<Atomic transactions AtomicStore Umax */
   ATOMICSTORE_UMIN       = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_UMIN,    /**<Atomic transactions AtomicStore Umin */
   ATOMICLOAD_ADD         = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_ADD,      /**<Atomic transactions AtomicLoad Add */
   ATOMICLOAD_CLR         = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_CLR,      /**<Atomic transactions AtomicLoad Clr */
   ATOMICLOAD_EOR         = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_EOR,      /**<Atomic transactions AtomicLoad Eor */
   ATOMICLOAD_SET         = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_SET,      /**<Atomic transactions AtomicLoad Set */
   ATOMICLOAD_SMAX        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_SMAX,     /**<Atomic transactions AtomicLoad Smax */
   ATOMICLOAD_SMIN        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_SMIN,     /**<Atomic transactions AtomicLoad Smin */
   ATOMICLOAD_UMAX        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_UMAX,     /**<Atomic transactions AtomicLoad Umax */
   ATOMICLOAD_UMIN        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_UMIN,     /**<Atomic transactions AtomicLoad Umin */
   ATOMICSWAP             = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSWAP,          /**<Atomic transactions AtomicSwap */
   ATOMICCOMPARE          = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICCOMPARE        /**<Atomic transactions AtomicCompare */ 

  } atomic_xact_op_type_enum;

  /** 
   * Enum to represent the Endianness of the outbound write data sent in Atomic transactions.
   * Following are the possible values:
   * - LITTLE_ENDIAN : Indicates that the outbound Atomic Write data is in the Little Endian format
   * - BIG_ENDIAN    : Indicates that the outbound Atomic Write data is in the Big Endian format
   * .
   */
  typedef enum {
    LITTLE_ENDIAN       =  0,
    BIG_ENDIAN          =  1
  } endian_enum;  

  /** 
   * Enum to represent the operation to be performed on the tags present in the corresponding DAT channel.
   * Following are the possible values:
   * - TAG_INVALID  : The tags are not valid.
   * - TAG_TRANSFER : The tags are clean. Tag Match does not need to be performed.
   * - TAG_UPDATE   : The Allocation Tag values have been updated and are dirty. The tags in memory should be updated.
   * - TAG_FETCH_MATCH    : The Physical Tags in the write must be checked against the Allocation Tag values obtained from memory, in 
   * -                      reads the allocation tags will be fetched from memory for read transactions.
   * .
   */
  typedef enum bit[(`SVT_AXI_TAGOP_WIDTH-1):0]{
    TAG_INVALID  = 0,
    TAG_TRANSFER = 1,
    TAG_UPDATE   = 2,
    TAG_FETCH_MATCH = 3
  } tag_op_enum;


 
/** 
   * Enum to represent the ‘Resp’ field in the TagMatch response.
   *  This field is only applicable for Write and Atomic transactions with TagOp in the request set to Match (TAG_FETCH_MATCH).
   *  This field will be populated by the VIP and must not be set by the users.
   * Following are the possible values:
   * - MATCH_NOT_PERFORMED  : The tag MATCH operation is not performed by the completer.
   * - NO_MATCH_RESULT  : The tag MATCH operation doesn't have a result.
   * - FAIL  : The tag MATCH operation is failed.
   * - PASS  : The tag MATCH operation is passed.
   * .
   */
 
  typedef enum bit[(`SVT_AXI_TAGOP_WIDTH-1):0] {
     MATCH_NOT_PERFORMED = 0,
     NO_MATCH_RESULT  = 1,
     FAIL = 2,
     PASS = 3
  } tag_match_resp_enum;  

`endif
 /**
   * Enum to represent four levels of shareability domain for snoop
   * transactions. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE. 
   */
  typedef enum bit [1:0] {
    NONSHAREABLE      = `SVT_AXI_DOMAIN_TYPE_NONSHAREABLE,
    INNERSHAREABLE    = `SVT_AXI_DOMAIN_TYPE_INNERSHAREABLE,
    OUTERSHAREABLE    = `SVT_AXI_DOMAIN_TYPE_OUTERSHAREABLE,
    SYSTEMSHAREABLE   = `SVT_AXI_DOMAIN_TYPE_SYSTEMSHAREABLE
  } xact_shareability_domain_enum;

  /**
   * Enum to represent barrier transaction type. Enum to represent four levels
   * of shareability domain for snoop transactions. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  typedef enum bit [1:0] {
    NORMAL_ACCESS_RESPECT_BARRIER = `SVT_AXI_NORMAL_ACCESS_RESPECT_BARRIER,
    MEMORY_BARRIER                = `SVT_AXI_MEMORY_BARRIER,
    NORMAL_ACCESS_IGNORE_BARRIER  = `SVT_AXI_NORMAL_ACCESS_IGNORE_BARRIER,
    SYNC_BARRIER                  = `SVT_AXI_SYNC_BARRIER
  } barrier_type_enum;

  /**
   * Enum to represent responses for a coherent transaction Additional read
   * response bits that provide information on the completion of a shareable
   * read transaction.  Enum to represent barrier transaction type. Enum to
   * represent four levels of shareability domain for snoop transactions.
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to
   * AXI_ACE.
   */
  typedef enum  bit [1:0] {
    UNIQUE_CLEAN   = `SVT_AXI_COHERENT_RESP_TYPE_UNIQUE_CLEAN, 
    UNIQUE_DIRTY   = `SVT_AXI_COHERENT_RESP_TYPE_UNIQUE_DIRTY,
    SHARED_CLEAN   = `SVT_AXI_COHERENT_RESP_TYPE_SHARED_CLEAN,
    SHARED_DIRTY   = `SVT_AXI_COHERENT_RESP_TYPE_SHARED_DIRTY
  } coherent_resp_type_enum;

  /**
   * Enum to represent locked type in a transaction
   */

  typedef enum bit [1:0] {
    NORMAL     = `SVT_AXI_TRANSACTION_NORMAL,
    EXCLUSIVE  = `SVT_AXI_TRANSACTION_EXCLUSIVE,
    LOCKED     = `SVT_AXI_TRANSACTION_LOCKED
  } atomic_type_enum;

  /**
   * Enum to represent the status of coherent exclusive access
   */
  typedef enum {
    EXCL_ACCESS_INITIAL  = `SVT_AXI_COHERENT_EXCL_ACCESS_INITIAL,
    EXCL_ACCESS_PASS     = `SVT_AXI_COHERENT_EXCL_ACCESS_PASS,
    EXCL_ACCESS_FAIL     = `SVT_AXI_COHERENT_EXCL_ACCESS_FAIL 
  } excl_access_status_enum;

  /** 
   * Enum to represent the status of master exclusive monitor, which indicates the cause of failure for a coherent exclusive store
   */ 
  typedef enum {
    EXCL_MON_INVALID  = `SVT_AXI_EXCL_MON_INVALID,
    EXCL_MON_SET      = `SVT_AXI_EXCL_MON_SET,
    EXCL_MON_RESET    = `SVT_AXI_EXCL_MON_RESET
  } excl_mon_status_enum;  

  /**
   * Enum to represent locked type in a transaction
   */

  typedef enum bit [2:0] {
    DATA_SECURE_NORMAL                = `SVT_AXI_DATA_SECURE_NORMAL,               
    DATA_SECURE_PRIVILEGED            = `SVT_AXI_DATA_SECURE_PRIVILEGED,               
    DATA_NON_SECURE_NORMAL            = `SVT_AXI_DATA_NON_SECURE_NORMAL,               
    DATA_NON_SECURE_PRIVILEGED        = `SVT_AXI_DATA_NON_SECURE_PRIVILEGED,           
    INSTRUCTION_SECURE_NORMAL         = `SVT_AXI_INSTRUCTION_SECURE_NORMAL,            
    INSTRUCTION_SECURE_PRIVILEGED     = `SVT_AXI_INSTRUCTION_SECURE_PRIVILEGED,         
    INSTRUCTION_NON_SECURE_NORMAL     = `SVT_AXI_INSTRUCTION_NON_SECURE_NORMAL,        
    INSTRUCTION_NON_SECURE_PRIVILEGED = `SVT_AXI_INSTRUCTION_NON_SECURE_PRIVILEGED    
  } prot_type_enum;

  /**
   * Enum to represent responses in a transaction
   */
  typedef enum bit [1:0] {
    OKAY    = `SVT_AXI_OKAY_RESPONSE,
    EXOKAY  = `SVT_AXI_EXOKAY_RESPONSE,
    SLVERR = `SVT_AXI_SLVERR_RESPONSE,
    DECERR  = `SVT_AXI_DECERR_RESPONSE
  } resp_type_enum;

  typedef enum bit [2:0] {
    INVALID = `SVT_AXI_CACHE_LINE_STATE_INVALID,
    UNIQUECLEAN = `SVT_AXI_CACHE_LINE_STATE_UNIQUECLEAN,
    SHAREDCLEAN = `SVT_AXI_CACHE_LINE_STATE_SHAREDCLEAN,
    UNIQUEDIRTY = `SVT_AXI_CACHE_LINE_STATE_UNIQUEDIRTY,
    SHAREDDIRTY = `SVT_AXI_CACHE_LINE_STATE_SHAREDDIRTY
  } cache_line_state_enum;
 
  /**
   * Enum to represent DVM Message type.
   *
   * The bit representation of this type matches the encoding of the DVM message type field
   * in the AxADDR AMBA4 signal.
   * 
   * Used in the svt_amba_pv_extension class.
   */
  typedef enum bit [2:0] {
    TLB_INVALIDATE                        = 'h0, /**< TLB invalidate */
    BRANCH_PREDICTOR_INVALIDATE           = 'h1, /**< Branch predictor invalidate */
    PHYSICAL_INSTRUCTION_CACHE_INVALIDATE = 'h2, /**< Physical instruction cache invalidate */
    VIRTUAL_INSTRUCTION_CACHE_INVALIDATE  = 'h3, /**< Virtual instruction cache invalidate */
    SYNC                                  = 'h4, /**< Synchronisation message */
    HINT                                  = 'h6  /**< Reserved message type for future Hint messages */
  } dvm_message_enum;

  /**
   * Enum to represent DVM message Guest OS or hypervisor type.
   *
   * The bit representation of this type matches the encoding of the DVM guest OS or 
   * hypervisor field in the AxADDR AMBA4 signal.
   */
  typedef enum bit [1:0] {
    HYPERVISOR_OR_GUEST = 'h0, /**< Transaction applies to hypervisor and all Guest OS*/
    GUEST               = 'h2, /**< Transaction applies to Guest OS */
    HYPERVISOR          = 'h3  /**< Transaction applies to hypervisor */
  } dvm_os_enum;

  /**
   * Enum to represent DVM message security type.
   *
   * The bit representation of this type matches the encoding of the DVM security field
   * in the AxADDR AMBA4 signal.
   */
  typedef enum bit [1:0] {
    AMBA_PV_SECURE_AND_NON_SECURE = 'h0, /**< Transaction applies to Secure and Non-secure */
    AMBA_PV_SECURE_ONLY           = 'h2, /**< Transaction applies to Secure only */
    AMBA_PV_NON_SECURE_ONLY       = 'h3  /**< Transaction applies to Non-secure only */
  } dvm_security_enum;


  /**
   *  Enum for interleave block pattern
   */

  typedef enum {
    EQUAL_BLOCK   = `SVT_AXI_TRANSACTION_INTERLEAVE_EQUAL_BLOCK,
    RANDOM_BLOCK  = `SVT_AXI_TRANASCTION_INTERLEAVE_RANDOM_BLOCK
  } interleave_pattern_enum;

  /** 
   *  Enum to represent address delay reference event
   */
  typedef enum {
    PREV_ADDR_VALID      =  `SVT_AXI_MASTER_TRANSACTION_PREV_ADDR_VALID_REF,
    PREV_ADDR_HANDSHAKE  =  `SVT_AXI_MASTER_TRANSACTION_PREV_ADDR_HANDSHAKE_REF,
    FIRST_WVALID_DATA_BEFORE_ADDR = `SVT_AXI_MASTER_TRANSACTION_FIRST_WVALID_DATA_BEFORE_ADDR,
    FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR = `SVT_AXI_MASTER_TRANSACTION_FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR,
    PREV_LAST_DATA_HANDSHAKE = `SVT_AXI_MASTER_TRANSACTION_PREV_LAST_DATA_HANDSHAKE
  } reference_event_for_addr_valid_delay_enum;

  /** 
   *  Enum to represent data delay reference event
   */
  typedef enum {
    WRITE_ADDR_VALID                           = `SVT_AXI_MASTER_TRANSACTION_WRITE_ADDR_VALID_REF,    
    //removed address handshake refrence because  of potential deadlock due to following reason::
    //the slave can wait for AWVALID or WVALID, or both before asserting AWREADY
    WRITE_ADDR_HANDSHAKE                       = `SVT_AXI_MASTER_TRANSACTION_WRITE_ADDR_HANDSHAKE_REF,
    PREV_WRITE_DATA_HANDSHAKE                  = `SVT_AXI_MASTER_TRANSACTION_PREV_WRITE_DATA_HANDSHAKE_REF
  }  reference_event_for_first_wvalid_delay_enum;

  typedef enum {
    PREV_WVALID            = `SVT_AXI_MASTER_TRANSACTION_PREV_WVALID_REF,
    PREV_WRITE_HANDSHAKE   = `SVT_AXI_MASTER_TRANSACTION_PREV_WRITE_HANDSHAKE_REF
  } reference_event_for_next_wvalid_delay_enum;
  
  /** 
   *  Enum to represent tvalid delay reference event
   */
  typedef enum {
    PREV_TVALID_TREADY_HANDSHAKE          = `SVT_AXI_MASTER_TRANSACTION_PREV_TVALID_TREADY_HANDSHAKE_REF,
    PREV_TVALID                           = `SVT_AXI_MASTER_TRANSACTION_PREV_TVALID_REF
  }  reference_event_for_tvalid_delay_enum;

  typedef enum {
    RVALID               = `SVT_AXI_MASTER_TRANSACTION_RVALID_REF,                                 
    MANUAL_RREADY        = `SVT_AXI_MASTER_TRANSACTION_MANUAL_RREADY_REF       
  } reference_event_for_rready_delay_enum;

  /** 
   *  Enum to represent response delay reference event
   */
  typedef enum {
    BVALID               =   `SVT_AXI_MASTER_TRANSACTION_BVALID_REF
  } reference_event_for_bready_delay_enum;
 
  /** 
   * Enum to represent read acknowledgment delay reference event. Applicable
   * when svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  typedef enum {
    LAST_READ_DATA_HANDSHAKE    = `SVT_AXI_MASTER_TRANSACTION_LAST_READ_DATA_HANDSHAKE_REF
  } reference_event_for_rack_delay_enum;
  
  /** 
   * Enum to represent write acknowledgment delay reference event. Applicable
   * when svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  typedef enum {
    WRITE_RESP_HANDSHAKE    = `SVT_AXI_MASTER_TRANSACTION_WRITE_RESP_HANDSHAKE_REF
  } reference_event_for_wack_delay_enum;

  /** 
   *  Enum to represent address delay reference event
   */
  typedef enum {
    ADDR_VALID               = `SVT_AXI_SLAVE_TRANSACTION_ADDR_VALID_REF,
    FIRST_WVALID            = `SVT_AXI_SLAVE_TRANSACTION_FIRST_WVALID_REF
  } reference_event_for_addr_ready_delay_enum;

  /** 
   *  Enum to represent reference event for delay for first rvalid
   */
  typedef enum {
    READ_ADDR_VALID               = `SVT_AXI_SLAVE_TRANSACTION_READ_ADDR_VALID_REF,    
    READ_ADDR_HANDSHAKE           = `SVT_AXI_SLAVE_TRANSACTION_READ_ADDR_HANDSHAKE_REF
  }  reference_event_for_first_rvalid_delay_enum;

  /** 
   *  Enum to represent reference event for delay for second rvalid onwards
   */
  typedef enum {
    PREV_RVALID          = `SVT_AXI_SLAVE_TRANSACTION_PREV_RVALID_REF,
    PREV_READ_HANDSHAKE  = `SVT_AXI_SLAVE_TRANSACTION_PREV_READ_HANDSHAKE_REF
  } reference_event_for_next_rvalid_delay_enum;

  /** 
   *  Enum to represent reference event for delay for wready signal
   */
  typedef enum {
    WVALID               = `SVT_AXI_SLAVE_TRANSACTION_WVALID_REF,                                 
    MANUAL_WREADY        = `SVT_AXI_SLAVE_TRANSACTION_MANUAL_WREADY_REF       
  } reference_event_for_wready_delay_enum;

  /** 
   *  Enum to represent write response delay reference event
   */
  typedef enum {
    LAST_DATA_HANDSHAKE = `SVT_AXI_SLAVE_TRANSACTION_LAST_DATA_HANDSHAKE_REF,
    ADDR_HANDSHAKE = `SVT_AXI_SLAVE_TRANSACTION_ADDR_HANDSHAKE_REF
  } reference_event_for_bvalid_delay_enum;

 
    
   // ****************************************************************************
   // Public Data
   // ****************************************************************************
   /** @groupname axi_misc
     * Variable that holds the object_id of this transaction
     */
   int object_id = -1;
   /** @groupname axi_misc
    * Variables used in generating XML/FSDB for pa writer 
    */
   
   string pa_object_type = "";
   string pa_channel_name ="" ;
   string bus_parent_uid = "";
   string bus_activity_type_name;

   /** @groupname axi_misc
     * The port configuration corresponding to this transaction
     */
   svt_axi_port_configuration port_cfg;
   
   /** 
    * @groupname ace_protocol
    * This member points to a barrier pair transaction
    * associated to this current transaction.  When associated_barrier_xact is
    * null, it indicates that this current transaction is not a post-barrier
    * transaction.  When associated_barrier_xact is non-null, this current
    * transaction will wait for responses from the barrier transactions in
    * associated_barrier_xact, before it can be transmitted.
    *
    * associated_barrier_xact can be set in the callback
    * svt_axi_master_callback::associate_xact_to_barrier_pair. In this
    * callback, user can associate this transaction with a barrier transaction
    * pair.
    *
    * Please refer to User Guide for more details on usage of this member.
    */
   svt_axi_barrier_pair_transaction  associated_barrier_xact;

`ifdef SVT_UVM_TECHNOLOGY
   /**
     * @groupname axi_misc 
     * Applicable only for master in ACTIVE mode.
     * If this transaction was generated from a UVM TLM Generic Payload, this
     * member indicates the GP from which this AXI transaction was generated
     */
   uvm_tlm_generic_payload causal_gp_xact;
`endif

  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------
  /** @cond PRIVATE */
  /** 
    * Object used to hold exceptions for a packet. 
    */
  `ifndef __SVDOC__
  svt_axi_transaction_exception_list exception_list = null; 
  `endif
 /** W riter used in callbacks to generate output for pa or verdi */ 
  protected svt_xml_writer xml_writer = null ;

  protected rand bit [`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0]  addr_mask ;

  protected rand bit [`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0]  addr_range;

  protected rand bit [`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0]  burst_addr_mask ;

  /** The maximum possible address based on addr_width. Calculated in pre_randomize */
  protected bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] max_possible_addr;

  /** The maximum possible address based on addr_width. Calculated in pre_randomize */

  //protected bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] max_possible_addr;

  /** The maximum possible address based on addr_user_width. Calculated in pre_randomize */
  protected bit [`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] max_possible_user_addr;

  /**
    * Used in system monitor to indicate if all bytes of a slave transaction
    * has been correlated to a corresponding master transaction
    */
  bit  is_slave_xact_correlated = 0;
  
  /**
    * Used in port monitor to indicate resize and aligned data status
    * in data_before_addr transaction.
    */
  bit  is_resize_and_align_data = 0;


  /** 
    * Indicates if data read from memory for a given beat contains X
    * The slave driver uses this information to decide whether to 
    * drive X on data.
    */
  bit read_data_contains_x[];

  /** The maximum possible address based on addr_user_width. Calculated in pre_randomize */
  // protected bit [`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] max_possible_user_addr;

  /** @endcond */

  /**
   * @groupname axi3_protocol
   * The variable holds the value of  AWID/WID/BID/ARID/RID signals.<br>
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_ID_WIDTH. Default value of this macro is 8. To change the
   * maximum width of this variable, user can change the value of this macro.
   * Define the new value for the macro in file svt_axi_user_defines.svi, and
   * then specify this file to be compiled by the simulator. Also, specify
   * +define+SVT_AXI_INCLUDE_USER_DEFINES on the simulator compilation command
   * line. Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_AXI_MAX_ID_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::id_width.
   */
  rand bit [`SVT_AXI_MAX_ID_WIDTH - 1:0] id = 0;

  /**
   * @groupname axi3_protocol
   * The variable represents AWADDR when xact_type is WRITE and  ARADDR when
   * xact_type is READ.<br>
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_ADDR_WIDTH. Default value of this macro is 64. To change the
   * maximum width of this variable, user can change the value of this macro.
   * Define the new value for the macro in file svt_axi_user_defines.svi, and
   * then specify this file to be compiled by the simulator. Also, specify
   * +define+SVT_AXI_INCLUDE_USER_DEFINES on the simulator compilation command
   * line. Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_AXI_MAX_ADDR_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::addr_width.
   */
  rand bit [`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0] addr = 0;
  
  /**
   * @groupname axi3_protocol
   * Represents the minimum byte address of this transaction. 
   * If tagging is enabled, this will be the minimum tagged address 
   *  .
   */
  rand bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] min_byte_addr =0;
  
  /**
   * @groupname axi3_protocol
   * Represents the maximum byte address of this transaction. 
   * If tagging is enabled, this will be the maximum tagged address 
   *  .
   */
  rand bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] max_byte_addr =0;
  
  /**
   * @groupname axi3_protocol
   * Represents the total byte count of this transaction. 
   *  .
   */
  rand int total_byte_count = 0;
  
  /**
   *  @groupname axi3_protocol
   *  The variable represents the actual length of the burst. For eg.
   *  burst_length = 1 means a burst of length 1.
   *
   *  If #svt_axi_port_configuration::axi_interface_type is AXI3, burst length
   *  of 1 to 16 is supported.
   *
   *  If #svt_axi_port_configuration::axi_interface_type is AXI4, burst length
   *  of 1 to 256 is supported.
   */ 
  rand bit [`SVT_AXI_MAX_BURST_LENGTH_WIDTH: 0] burst_length = 1;

  /**
   *  @groupname axi3_protocol
   *  Represents the burst size of a transaction . The variable holds the value
   *  for AWSIZE/ARSIZE. 
   */
  rand burst_size_enum burst_size = BURST_SIZE_8BIT;

  /**
   *  @groupname axi3_protocol
   *  Represents the burst type of a transaction. The burst type holds the value
   *  for AWBURST/ARBURST. Following are the possible burst types: 
   *  - FIXED
   *  - INCR
   *  - WRAP
   *  .
   */
  rand burst_type_enum burst_type = INCR;

  /**
   * @groupname axi3_protocol
   * Represents the transaction type.
   * Following are the possible transaction types:
   * - WRITE    : Represent a WRITE transaction. 
   * - READ     : Represents a READ transaction.
   * - COHERENT : Represents a COHERENT transaction.
   * .
   *
   * Please note that WRITE and READ transaction type is valid for
   * #svt_axi_port_configuration::axi_interface_type is AXI3/AXI4/AXI4_LITE and
   * COHERENT transaction type is valid for
   * #svt_axi_port_configuration::axi_interface_type is AXI_ACE.
   */
  rand xact_type_enum xact_type = WRITE;
  
  /**
   * @groupname axi3_protocol
   * Represents the phase type.
   * Following are the possible transaction types:
   * - WRITE    : Represent a WRITE transaction. 
   * - READ     : Represents a READ transaction.
   * .
   *
   * Please note that WRITE and READ transaction type is valid for
   * #svt_axi_port_configuration::axi_interface_type is AXI3/AXI4/AXI4_LITE 
   */
  phase_type_enum phase_type = WR_ADDR;

  /**
   * @groupname axi3_protocol
   * Represents the atomic access of a transaction.  The variable holds the
   * value for AWLOCK/ARLOCK. Following are the possible atomic types:
   * - NORMAL     
   * - EXCLUSIVE  
   * - LOCKED
   * .
   * Please note that atomic type LOCKED is not yet supported.
   */
  rand atomic_type_enum atomic_type = NORMAL;

`ifdef SVT_ACE5_ENABLE
  /**
   * Indicates the endianness of the Outbound Write Data in an Atomic transaction.
   */
  rand endian_enum endian = LITTLE_ENDIAN;
`endif

`ifdef SVT_ACE5_ENABLE
  /**
   * @groupname axi5_protocol
   * Represents the Unique ID indicator Feature.
   * The variable holds the value of AWIDUNQ/BIDUNQ/ARIDUNQ/RIDUNQ signals.<br>
   * The Variable is used to indicate that there are
   * no outstanding transactions going on with the same AWID/BID/ARID/RID respectively
   * and it will remain unique till the transaction is completed.
   * In order to use this feature, user need to pass the user defined macro
   * at compile time +define+SVT_ACE5_ENABLE.
   * Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_ACE5_ENABLE macro is only used to enable this feature and signals.
   * The Signals can be configured and enabled by VIP configuration using
   * parameter svt_axi_port_configuration::unique_id_enable.
   *
   * This functionality is not supported yet.
   */
  rand bit unique_id = 0;
`endif

  /**
   *  @groupname axi3_protocol
   *  Represents the cache support of a transaction. The variable holds the
   *  value for AWCACHE/ARCACHE.
   *
   *  Following values are supported in AXI3 mode:
   *
   *  - SVT_AXI_3_NON_CACHEABLE_NON_BUFFERABLE            
   *  - SVT_AXI_3_BUFFERABLE_OR_MODIFIABLE_ONLY           
   *  - SVT_AXI_3_CACHEABLE_BUT_NO_ALLOC                  
   *  - SVT_AXI_3_CACHEABLE_BUFFERABLE_BUT_NO_ALLOC       
   *  - SVT_AXI_3_CACHEABLE_WR_THRU_ALLOC_ON_RD_ONLY      
   *  - SVT_AXI_3_CACHEABLE_WR_BACK_ALLOC_ON_RD_ONLY      
   *  - SVT_AXI_3_CACHEABLE_WR_THRU_ALLOC_ON_WR_ONLY       
   *  - SVT_AXI_3_CACHEABLE_WR_BACK_ALLOC_ON_WR_ONLY       
   *  - SVT_AXI_3_CACHEABLE_WR_THRU_ALLOC_ON_BOTH_RD_WR    
   *  - SVT_AXI_3_CACHEABLE_WR_BACK_ALLOC_ON_BOTH_RD_WR    
   *  .
   *  
   *  Following values for ARCACHE are supported in AXI4 mode:
   *  - SVT_AXI_4_ARCACHE_DEVICE_NON_BUFFERABLE                  
   *  - SVT_AXI_4_ARCACHE_DEVICE_BUFFERABLE                     
   *  - SVT_AXI_4_ARCACHE_NORMAL_NON_CACHABLE_NON_BUFFERABLE    
   *  - SVT_AXI_4_ARCACHE_NORMAL_NON_CACHABLE_BUFFERABLE         
   *  - SVT_AXI_4_ARCACHE_WRITE_THROUGH_NO_ALLOCATE                
   *  - SVT_AXI_4_ARCACHE_WRITE_THROUGH_READ_ALLOCATE           
   *  - SVT_AXI_4_ARCACHE_WRITE_THROUGH_WRITE_ALLOCATE          
   *  - SVT_AXI_4_ARCACHE_WRITE_THROUGH_READ_AND_WRITE_ALLOCATE 
   *  - SVT_AXI_4_ARCACHE_WRITE_BACK_NO_ALLOCATE                
   *  - SVT_AXI_4_ARCACHE_WRITE_BACK_READ_ALLOCATE                
   *  - SVT_AXI_4_ARCACHE_WRITE_BACK_WRITE_ALLOCATE             
   *  - SVT_AXI_4_ARCACHE_WRITE_BACK_READ_AND_WRITE_ALLOCATE      
   *  .
   *
   *  Following values for AWCACHE are supported in AXI4 mode:
   *  - SVT_AXI_4_AWCACHE_DEVICE_NON_BUFFERABLE                  
   *  - SVT_AXI_4_AWCACHE_DEVICE_BUFFERABLE                     
   *  - SVT_AXI_4_AWCACHE_NORMAL_NON_CACHABLE_NON_BUFFERABLE    
   *  - SVT_AXI_4_AWCACHE_NORMAL_NON_CACHABLE_BUFFERABLE         
   *  - SVT_AXI_4_AWCACHE_WRITE_THROUGH_NO_ALLOCATE                
   *  - SVT_AXI_4_AWCACHE_WRITE_THROUGH_READ_ALLOCATE           
   *  - SVT_AXI_4_AWCACHE_WRITE_THROUGH_WRITE_ALLOCATE          
   *  - SVT_AXI_4_AWCACHE_WRITE_THROUGH_READ_AND_WRITE_ALLOCATE 
   *  - SVT_AXI_4_AWCACHE_WRITE_BACK_NO_ALLOCATE                
   *  - SVT_AXI_4_AWCACHE_WRITE_BACK_READ_ALLOCATE                
   *  - SVT_AXI_4_AWCACHE_WRITE_BACK_WRITE_ALLOCATE             
   *  - SVT_AXI_4_AWCACHE_WRITE_BACK_READ_AND_WRITE_ALLOCATE    
   *  .
   */

  rand bit [`SVT_AXI_CACHE_WIDTH - 1:0] cache_type = 0;

  /**
   *  @groupname axi3_protocol
   *  Represents the protection support of a transaction. The variable holds the
   *  value for AWPROT/ARPROT. The conventions of the enumeration are:
   *
   *  - NORMAL/PRIVILEGED   : Normal/Priveleged access represented by AWPROT[0]/ARPROT[0]
   *  - SECURE / NON_SECURE : Secure/Non-Secure access represented by AWPROT[1]/ARPROT[1]
   *  - DATA / INSTRUCTION  : Data/Instruction access represented by AWPROT[2]/ARPROT[2]
   *  .
   *
   *  For the above conventions, following are the possible protection types:
   *  - DATA_SECURE_NORMAL                    
   *  - DATA_SECURE_PRIVILEGED                    
   *  - DATA_NON_SECURE_NORMAL                    
   *  - DATA_NON_SECURE_PRIVILEGED                
   *  - INSTRUCTION_SECURE_NORMAL                 
   *  - INSTRUCTION_SECURE_PRIVILEGED              
   *  - INSTRUCTION_NON_SECURE_NORMAL
   *  - INSTRUCTION_NON_SECURE_PRIVILEGED
   *  .
   */

  rand  prot_type_enum prot_type = DATA_SECURE_NORMAL;

  /**
   *  @groupname ace_protocol
   *  Applicable when
   *  svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.  
   *  Users  who need to bypass lookup of cache to determine valid 
   *  initial cache line states can set this property to 1.
   *  In order to randomize this property to 1, the user must switch off 
   *  svt_axi_master_transaction::reasonable_bypass_cache_lookup constraint.
   *  Setting this property will enable transactions to be sent out even
   *  if the initial cache state does not meet requirements set by ACE 
   *  protocol. Please note that coherency is not guaranteed when this 
   *  property is set
   *
   * Applicable for ACTIVE MASTER only.
   */

  rand  bit bypass_cache_lookup = 1'b0;  


  /**
   * @groupname axi3_protocol
   * MASTER in active mode:
   *
   * For write transactions this variable specifies write data to be driven on the
   * WDATA bus. 
   * 
   * SLAVE in active mode:
   *
   * For read transactions this variable specifies read data to be driven on the
   * RDATA bus.
   *
   * PASSIVE MODE:
   * This variable stores the write or read data as seen on WDATA or RDATA bus.
   *
   * APPLICABLE IN ALL MODES:
   * If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   * data must be stored right-justified by the user. The model will drive the
   * data on the correct lanes.  If svt_axi_port_configuration::wysiwyg_enable
   * is set to 1, the data is  transmitted as programmed by user and is
   * reported as seen on bus. No right-justification is used in this case.<br>
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_DATA_WIDTH. Default value of this macro is 1024. To change the
   * maximum width of this variable, user can change the value of this macro.
   * Define the new value for the macro in file svt_axi_user_defines.svi, and
   * then specify this file to be compiled by the simulator. Also, specify
   * +define+SVT_AXI_INCLUDE_USER_DEFINES on the simulator compilation command
   * line. Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_AXI_MAX_DATA_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::data_width.
   */

`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] data[];
`else
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] data[];
`endif

`ifdef SVT_ACE5_ENABLE

 /**
   * @groupname ace5_protocol
   * This variable represents the read data for the atomic load,swap and compare transactions.
   * This data will be driven by the slave on the read data channel.
   * APPLICABLE IN ALL MODES:
   * If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   * data must be stored right-justified by the user. The model will drive the
   * data on the correct lanes.  If svt_axi_port_configuration::wysiwyg_enable
   * is set to 1, the data is  transmitted as programmed by user and is
   * reported as seen on bus. No right-justification is used in this case.<br>
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_DATA_WIDTH. Default value of this macro is 1024. To change the
   * maximum width of this variable, user can change the value of this macro.
   * Define the new value for the macro in file svt_axi_user_defines.svi, and
   * then specify this file to be compiled by the simulator. Also, specify
   * +define+SVT_AXI_INCLUDE_USER_DEFINES on the simulator compilation command
   * line. Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_AXI_MAX_DATA_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::data_width.
   */
`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_read_data[];
`else
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_read_data[];
`endif

//---------------------------------------------------------------------------------------------

/**
  * @groupname ace5_protocol
  * This field defines the Memory Tag value in the transaction driven on the data channel for transactions.
  * Every 4 bits of Tag correspond to one 16 byte chunk of data.
  * MASTER in active mode:
  *
  * For write transactions this variable specifies tags to be driven on the
  * WTAG bus. 
  * 
  * SLAVE in active mode:
  *
  * For read transactions this variable specifies tags to be driven on the
  * RTAG bus.
  *
  * PASSIVE MODE:
  * This variable stores the tags as seen on WTAG or RTAG bus.
  *
  *
  */
`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_TAG_WIDTH - 1:0] tag[];
`else
  rand bit [`SVT_AXI_MAX_TAG_WIDTH - 1:0] tag[];
`endif

//---------------------------------------------------------------------------------------------

/**
  * @groupname ace5_protocol
  * This field defines the WTAGUPDATE value in the transaction.
  * Only applicable when the Tag value is passed in the transaction and the tagop field in 
  * the transaction is set to Update.
  * Each WTAGUPDATE bit corresponds to 4 bits of WTAG
  */

`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_TAGUPDATE_WIDTH - 1:0] tag_update[];
`else
  rand bit [`SVT_AXI_MAX_TAGUPDATE_WIDTH - 1:0] tag_update[];
`endif

/**
  * @groupname ace5_protocol
  * This field defines the BCOMP value in the transaction.
  * Indicates whether write transaction is observable at the completer endused for persistent CMOs on Write channel.
  * This is used to send the response to a tag Match operation.
  * This is also used for persistent CMOs on Write channel.
  */
 
 rand bit is_write_transaction_observable = 0;
//---------------------------------------------------------------------------------------------
 
 /** 
   * Enum to represent the operation to be performed on the tags present in the corresponding DATA channel.
   * Following are the possible values:
   * - INVALID  : The tags are not valid.
   * - TRANSFER : The tags are clean. Tag Match does not need to be performed.
   * - UPDATE   : The Allocation Tag values have been updated and are dirty. The tags in memory should be updated.
   * - MATCH    : The Physical Tags in the write must be checked against the Allocation Tag values obtained from memory.
   * .
   */
  rand tag_op_enum tag_op = TAG_INVALID ;

  /** 
   * Enum to represent the response sent by the completer on the corresponding Response channel.
   * Following are the possible values:
   * - INVALID  : The tags are not valid.
   * - TRANSFER : The tags are clean. Tag Match does not need to be performed.
   * - UPDATE   : The Allocation Tag values have been updated and are dirty. The tags in memory should be updated.
   * - MATCH    : The Physical Tags in the write must be checked against the Allocation Tag values obtained from memory.
   * .
   */
 rand tag_op_enum response_tag_op = TAG_INVALID;
 
//---------------------------------------------------------------------------------------------

/** 
   * Enum to represent the ‘Resp’ field in the TagMatch response.
   *  This field is only applicable for Write and Atomic transactions with TagOp in the request set to Match (TAG_FETCH_MATCH).
   * Following are the possible values:
   * - MATCH_NOT_PERFORMED  : The tag MATCH operation is not performed by the completer.
   * - NO_MATCH_RESULT  : The tag MATCH operation doesn't have a result.
   * - FAIL  : The tag MATCH operation is failed.
   * - PASS  : The tag MATCH operation is passed.
   * .
   */
   rand tag_match_resp_enum tag_match_resp = MATCH_NOT_PERFORMED ;

//---------------------------------------------------------------------------------------------
 /**
   * @groupname ace5_protocol
   * This field defines the partition ID value in MPAM. This corresponds to AxMPAM[9:1] attribute.
   */
  rand bit [`SVT_AXI_MAX_MPAM_PARTID_WIDTH - 1:0] mpam_partid;

 /**
   * @groupname ace5_protocol
   * This field defines the Perfromance Monitor Group (PMG) value in MPAM. This corresponds to AxMPAM[10] attribute.
   */
  rand bit [`SVT_AXI_MAX_MPAM_PERFMONGROUP_WIDTH - 1:0] mpam_perfmongroup;

 /**
   * @groupname ace5_protocol
   * This field defines the MPAM_NS value in MPAM. This corresponds to AxMPAM[0] attribute.
   */
  rand bit [`SVT_AXI_MPAM_NS_WIDTH - 1:0] mpam_ns;
//---------------------------------------------------------------------------------------------

 /**
   * @groupname ace5_protocol
   * This variable represents the data that will be stored in the memory for atomic transactions 
   * after the atomic operation is performed.
   * APPLICABLE IN ALL MODES:
   * The SVT_AXI_MAX_DATA_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::data_width.
   */
`ifdef SVT_MEM_LOGIC_DATA
  logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_resultant_data[];
`else
  bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_resultant_data[];
`endif


//---------------------------------------------------------------------------------------------

 /**
   * @groupname ace5_protocol
   * This variable represents the swap data value for the atomic compare transactions.
   * This will not be programmed by the user.This is an internal variable and is populated by the AXI SLAVE.
   * 
   */

`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_swap_data[];
`else
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_swap_data[];
`endif

//---------------------------------------------------------------------------------------------
 /**
   * @groupname ace5_protocol
   * This variable represents the compare data value for the atomic compare transactions.
   * This will not be programmed by the user.This is an internal variable and is populated by the AXI SLAVE.
   */

`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_compare_data[];
`else
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_compare_data[];
`endif

`endif

  /**
   * @groupname axi3_protocol
   * MASTER in active mode:
   *
   * For write transactions this variable specifies write data to be driven on the
   * WDATA bus. 
   * 
   * SLAVE in active mode:
   *
   * For read transactions this variable specifies read data to be driven on the
   * RDATA bus.
   *
   * PASSIVE MODE:
   * This variable stores the write or read data as seen on WDATA or RDATA bus.
   *
   *
   */

`ifdef SVT_MEM_LOGIC_DATA
   logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] physical_data[];
`else
   bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] physical_data[];
`endif

`ifdef SVT_ACE5_ENABLE
 /**
   * @groupname ace5_protocol
   * This variable is only applicable for atomic transactions.
   * MASTER in active mode:
   * For Atomic LOAD , SWAP and COMPARE transactions specifies read data as seen on the RDATA bus. 
   * 
   * SLAVE in active mode:
   * This variable represents the read data for the atomic load,swap and compare transactions to be driven on the RDATA bus.
   *
   * PASSIVE MODE:
   * This variable stores the read data as seen on RDATA bus.
   *
   */

`ifdef SVT_MEM_LOGIC_DATA
   logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_read_physical_data[];
`else
   bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_read_physical_data[];
`endif

`endif

  /** @cond PRIVATE */
  /**
    * The data array in string format. Used by psdisplay_short
    */
  local string data_str = "";

`ifdef SVT_ACE5_ENABLE
  /**
    * The data array in string format. Used by psdisplay_short
    */
  local string atomic_read_data_str = "";
`endif

  /**
    * The wstrb array in string format. Used by psdisplay_short
    */
  local string wstrb_str = "";

  /**
    * The read response array in string format. Used by psdisplay_short
    */
  local string rresp_str = "";

  /**
    * The write response in string format. Used by psdisplay_short
    */
  local string bresp_str = "";

  /**
    * The valid_assertion_time in string format. Used by psdisplay_short
    */
  local string valid_assertion_time = "";
  
  /**
    * The ready_assertion_time in string format. Used by psdisplay_short
    */
  local string ready_assertion_time = "";
  
 /* holds transactions that attempt to access same cacheline at the same time current transaction

   * does and started before current transaction started */
  bit overlapped_xact_started_before[svt_axi_transaction];

  /* holds transactions that attempt to access same cacheline at the same time current transaction
   * does and started after current transaction started */
  bit overlapped_xact_started_after[svt_axi_transaction];
  
  /* Indicates xact complets with out_of_order*/
  bit is_xact_completed_out_of_order = 0;

  /* indicates how many transactions blocked progress of current transaction */
  int num_xacts_blocked_progress_of_curr_xact = 0;

  /* semaphore to access num_xacts_blocked_progress_of_curr_xact */
  semaphore sema_num_xacts_blocked_progress_of_curr_xact = new(1);
  /** @endcond */

  
  /**
   *  @groupname axi3_protocol
   *  Array of Write strobes.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   *  wstrb must be stored right-justified by the user. The model will drive
   *  these strobes on the correct lanes.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 1, the wstrb is  
   *  transmitted as programmed by user and is reported as seen on bus. 
   *  No right-justification is used in this case.
   */
  rand bit [`SVT_AXI_WSTRB_WIDTH - 1:0] wstrb[];

`ifdef SVT_ACE5_ENABLE
 
//---------------------------------------------------------------------------------------------
 /**
   * @groupname ace5_protocol
   * This variable represents the swap write strobes  value for the atomic compare transactions.
   * This must not be programmed by the user.This is an internal variable populated by the AXI SLAVE.
   * 
   */
  rand bit [`SVT_AXI_WSTRB_WIDTH - 1:0] atomic_swap_wstrb[];

//---------------------------------------------------------------------------------------------
 /**
   * @groupname ace5_protocol
   * This variable represents the compare write strobes value for the atomic compare transactions.
   * This must not be programmed by the user.This is an internal variable populated by the AXI SLAVE.
   */
   rand bit [`SVT_AXI_WSTRB_WIDTH - 1:0] atomic_compare_wstrb[];

`endif

  /**
   *  @groupname ace5_protocol
   *  Array of poison.It indicates the 
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   *  poison must be stored right-justified by the user. The model will drive
   *  these strobes on the correct lanes.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 1, the poison is  
   *  transmitted as programmed by user and is reported as seen on bus. 
   *  No right-justification is used in this case.
   */
  rand bit [`SVT_AXI_MAX_DATA_WIDTH/64- 1:0] poison[];

`ifdef SVT_ACE5_ENABLE
   /**
   *  @groupname ace5_protocol
   *  Array of poisonal value driven by the active slave on the read data channel.
   *  This is onlyapplicable for Atomic LOad , Swap and compare transactions.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   *  poison must be stored right-justified by the user. The model will drive
   *  these strobes on the correct lanes.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 1, the poison is  
   *  transmitted as programmed by user and is reported as seen on bus. 
   *  No right-justification is used in this case.
   */
  rand bit [`SVT_AXI_MAX_DATA_WIDTH/64- 1:0] atomic_read_poison[];

`endif


  /**
   *  @groupname axi3_protocol
   *  This variable specifies the response for write transaction. The variable holds the
   *  value for BRESP. Following are the possible response types:
   *  - OKAY    
   *  - EXOKAY  
   *  - SLVERR 
   *  - DECERR  
   *  .
   *          
   *  MASTER ACTIVE MODE:
   *
   *  Will Store the write response received from the slave.
   *
   *  SLAVE ACTIVE MODE:
   *
   *  The write response programmed by the user.
   *
   *  PASSIVE MODE - MASTER/SLAVE:
   *
   *  Stores the write response seen on the bus.
   */

  rand resp_type_enum bresp = OKAY;

  /**
   *  @groupname axi3_protocol
   *  This array variable specifies the response for read transaction. The array holds the
   *  value for RRESP. Following are the possible response types:
   *  - OKAY    
   *  - EXOKAY  
   *  - SLVERR 
   *  - DECERR  
   *  .
   *          
   *  MASTER ACTIVE MODE:
   *
   *  Will Store the read responses received from the slave.
   *
   *  SLAVE ACTIVE MODE:
   *
   *  The read responses programmed by the user.
   *
   *  PASSIVE MODE - MASTER/SLAVE:
   *
   *  Stores the read responses seen on the bus.
   */

  rand resp_type_enum rresp[];

`ifndef SVT_AXI_MULTI_SIM_OVERLAP_ADDR_ISSUE 
  /** 
    * @groupname axi3_protocol
    * If set, the driver checks if this transaction accesses a location
    * addressed by a previous transaction from this port or from some other
    * master. If there are any such previous transactions, this transaction is
    * blocked until all those transactions complete.  Also, the driver does not
    * pull any more transactions until this transaction is unblocked.  If not set,
    * this transaction is not checked for access to a location which was
    * previously accessed by another transaction.  Applicable only when
    * svt_axi_system_configuration::overlap_addr_access_control_enable is set 
    *
    * Applicable for ACTIVE MASTER only
    */ 
  rand bit check_addr_overlap = 1'b0;

  /** @cond PRIVATE */
  /**
    * @groupname axi3_protocol
    * Suspends a master transaction until this bit is reset. This is checked
    * immediately after a transaction is pulled by the driver from the sequencer
    * after the post_input_port_get callback is issued by the driver. When set,
    * the driver does not pull any more transactions from the
    * sequencer/generator until the bit is reset
    *
    * Applicable for ACTIVE MASTER only
    */
  bit suspend_master_xact = 1'b0;
  /** @endcond */
   
`endif

  /** @cond PRIVATE */
  /**
    * @groupname ace_protocol
    * This bit is set by master if a cache line is reserved for the transaction. 
    * Thie field is used by task which unreserves the cache line at the end of 
    * transaction to filtering. This is to ensure only command that reserved 
    * cache line should unreserve cache line.  
    *  
    * Applicable for ACTIVE MASTER only
    */
  bit is_cacheline_reserved = 1'b0;
  /** @endcond */

  /**
    * @groupname axi3_protocol
    * A bit that indicates that the testbench would like to suspend response/data
    * for a READ/WRITE/COHERENT transaction until this bit is reset. 
    * This bit is usually set by the testbench when it needs to provide
    * response information to the driver (the slave driver expects the response
    * information in 0 time), but the data to respond with is
    * not yet known.  The testbench can set this bit and put this transaction 
    * back into the input channel of the slave. 
    * The transaction's response/data will not be sent until this bit is reset. 
    * Once the data is available, the testbench can populate response fields 
    * and reset this bit, upon which the slave driver will send the 
    * response/data of this transaction.
    *
    * Applicable for ACTIVE SLAVE only.
    */
  bit suspend_response = 0;

 /**
    * @groupname axi3_protocol
    * A bit that indicates that the testbench would like to suspend awready signal 
    * for a WRITE transaction until this bit is reset. 
    * This is applicable only when svt_axi_port_configuration::default_awready is set to 0
    * svt_axi_transaction::addr_ready_delay won't be applicable when this bit is set to 1
    *
    * Applicable for ACTIVE SLAVE only.
    */
  bit suspend_awready = 0;

 /**
    * @groupname axi3_protocol
    * A bit that indicates that the testbench would like to suspend arready signal 
    * for a READ transaction until this bit is reset. 
    * This is applicable only when svt_axi_port_configuration::default_arready is set to 0
    * svt_axi_transaction::addr_ready_delay won't be applicable when this bit is set to 1
    *
    * Applicable for ACTIVE SLAVE only.
    */
  bit suspend_arready = 0;

 /**
    * @groupname axi3_protocol
    * A bit that indicates that the testbench would like to suspend wready signal 
    * for a WRITE transaction until this bit is reset. 
    * This is applicable only when svt_axi_port_configuration::default_wready is set to 0
    * svt_axi_transaction::wready_delay won't be applicable when this bit is set to 1
    *
    * Applicable for ACTIVE SLAVE only.
    */
  bit suspend_wready = 0;

  /**
    * @groupname ace_protocol
    * Represents the value of AWUNIQUE signal driven/sampled on the interface.
    * Applicable when svt_axi_port_configuration::awunique_enable is set.
    * AWUNIQUE is asserted as per table C3-9 of section C3.1.4 on AWUNIQUE
    * signal. The value in the randomized transaction may be overridden by the
    * driver as per protocol requirements. For transactions where AWUNIQUE may
    * be asserted or deasserted, the randomized value is driven.  
    */
  rand bit is_unique = 0;

  /**
   *  @groupname axi3_4_status
   *  Represents the current status of the read or write address.  Following are the
   *  possible status types.

   * - INITIAL               : Address phase has not yet started on the channel
   * - ACTIVE                : Address valid is asserted but ready is not 
   * - ACCEPT                : Address phase is complete 
   * - ABORTED               : Current transaction is aborted
   * .
   */

  status_enum addr_status = INITIAL;

  /**
   *  @groupname axi3_4_status
   *  Represents the status of the read or write data transfer.  Following are
   *  the possible status types.

   *  - INITIAL               : Data has not yet started on the channel
   *  - ACTIVE                : Data valid is asserted but ready is not asserted for the
   *                            current data beat. The current beat is indicated
   *                            by #current_data_beat_num variable
   *  - PARTIAL_ACCEPT        : The current data beat is completed but the next
   *                            data-beat is not started. The next data beat is
   *                            indicated by #current_data_beat_num
   *  - ACCEPT                : Data phase is complete 
   *  - ABORTED               : Current transaction is aborted 
   *  .
   */

  status_enum data_status = INITIAL;

`ifdef SVT_ACE5_ENABLE
/**
   *  @groupname axi3_4_status
   *  Represents the status of the read or write data transfer.  Following are
   *  the possible status types.

   *  - INITIAL               : Data has not yet started on the channel
   *  - ACTIVE                : Data valid is asserted but ready is not asserted for the
   *                            current data beat. The current beat is indicated
   *                            by #current_data_beat_num variable
   *  - PARTIAL_ACCEPT        : The current data beat is completed but the next
   *                            data-beat is not started. The next data beat is
   *                            indicated by #current_data_beat_num
   *  - ACCEPT                : Data phase is complete 
   *  - ABORTED               : Current transaction is aborted 
   *  .
   */

  status_enum atomic_read_data_status = INITIAL;
`endif

  /**
   *  @groupname axi3_4_status
   *  Represents the status of the write response transfer.  Following are
   *  the possible status types.
   *  - INITIAL               : Response has not yet started on the channel
   *  - ACTIVE                : BVALID is asserted, but not BREADY
   *  - ACCEPT                : Write response is complete
   *  - ABORTED               : Current transaction is aborted 
   *  .
   */


  status_enum write_resp_status = INITIAL;

  /**
   * @groupname ace_status
   * Represents the status of the read/write acknowledge sent via RACK/WACK for
   * ACE interface. RACK/WACK is asserted for a single cycle.
   * Following are  the possible status types:
   * - INITIAL               : RACK/WACK has not be asserted
   * - ACTIVE                : RACK/WACK is asserted
   * - ACCEPT                : RACK/WACK assertion is completed
   * - ABORTED               : Current transaction is aborted
   * .
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to
   * AXI_ACE.
   */

  status_enum ack_status = INITIAL;

  /**
   * @groupname ace_status
   * Represents the status of coherent exclusive access.
   * Following are  the possible status types: 
   * - EXCL_ACCESS_INITIAL   : Initial state of the transaction before it is processed by master 
   * - EXCL_ACCESS_PASS      : ACE exclusive access is successful
   * - EXCL_ACCESS_FAIL      : ACE exclusive access is failed
   * .
   *
   * A combination of #excl_access_status and #excl_mon_status can be used to
   * determine the reason for failure of exclusive store. Please refer to the
   * User Guide for more description. 
   */
  excl_access_status_enum  excl_access_status = EXCL_ACCESS_INITIAL;
  

  /**
   * @groupname ace_status
   * Represents the status of master exclusive monitor, which indicates the
   * cause of failure for a coherent exclusive store.  It is valid only for
   * exclusive store transaction, that is, CleanUnique. For all other
   * transactions it is set to EXCL_MON_INVALID by default.
   * Following are  the possible status types:
   * - EXCL_MON_INVALID      : Master exclusive monitor does not monitor the exclusive access on the cache line associated with the transaction
   * - EXCL_MON_SET          : Master exclusive monitor is set for exclusive access on the cache line associated with the transaction
   * - EXCL_MON_RESET        : Master exclusive monitor is reset for exclusive access on the cache line associated with the transaction
   * .
   *
   * A combination of #excl_access_status and #excl_mon_status can be used to
   * determine the reason for failure of exclusive store. Please refer to the
   * User Guide for more description.
   */ 
  excl_mon_status_enum   excl_mon_status = EXCL_MON_INVALID;


  /**
   *  @groupname axi3_4_status
   *    This is a counter which is incremented for every beat. Useful when user
   *    would try to access the transaction class to know its current state.
   *    This represents the beat number for which the status is reflected in
   *    member data_status.
   */
  int  current_data_beat_num = 0;
`ifdef SVT_ACE5_ENABLE
 /**
   *  @groupname axi3_4_status
   *    This is a counter which is incremented for every beat. Useful when user
   *    would try to access the transaction class to know its current state.
   *    This represents the beat number for which the status is reflected in
   *    member data_status.
   */
  int  atomic_read_current_data_beat_num = 0;
`endif
  /**
   *  @groupname interleaving
   *  Represents the various interleave pattern for a read and write transaction.
   *  The interleave_pattern gives flexibility to program interleave blocks with
   *  different patterns as mentioned below.
   *
   *  A Block is group of beats within a transaction.
   *
   *  EQUAL_BLOCK         : Drives equal distribution of blocks provided by
   *                        #equal_block_length variable. 
   *
   *  RANDOM_BLOCK        : Drives the blocks programmed in random_interleave_array
   *
   * Please note that currently interleaving based on EQUAL_BLOCK is not
   * supported.
   */
  rand interleave_pattern_enum interleave_pattern = RANDOM_BLOCK;

  /** @cond PRIVATE */
  /**
   *  @groupname interleaving
   *  If the interleave_pattern is set to EQUAL_BLOCK then this variable 
   *  is used to define the block length.
   *  Please note that currently interleaving based on EQUAL_BLOCK is not
   *  supported.
   */

  rand int equal_block_length = 0;

  /** @endcond */

  /**
   *  @groupname interleaving
   *  When the interleave_pattern is set to RANDOM_BLOCK, the user would
   *  program this array with blocks. There are default constraints, which the
   *  user can override and set their own block patterns.
   */
  rand int random_interleave_array[];


  /** @cond PRIVATE */
  /**
   *  @groupname interleaving
   *  This variable will start a new interleave from the current transaction and
   *  informs the model to complete all the transactions prior to this
   *  transaction.
   *
   *  Example 1:
   *  Interleave depth = 2
   * 
   *  Requirement : 
   *  1) Interleave transaction 1- 10 with each other
   *  2) Interleave transactions 11 - 20 with each other
   *
   *  Solution :
   *  1) Program start_new_interleave=0 for transactions 1 - 10 
   *  2) Program start_new_interleave=1 for transaction 11
   *
   *  Example 2:
   *  Interleave depth = 2
   *
   *  Requirement :
   *  1) Do not Interleave transactions 1 - 10
   *  2) Start Interleaving from transactions 11 - 20
   *
   *  Solution :
   *  1) Program start_new_interleave=1 for transactions 1-10
   *  2) Program start_new_interleave=1 for transaction 11
   *
   *  Please note that this parameter is not currently supported.
   */
  rand bit start_new_interleave = 0;
  /** @endcond */

  /**
   * @groupname interleaving , out_of_order
   * This variable controls enabling of interleaving for the current transaction.
   * 
   * Example:
   * svt_axi_port_configuration::read_data_reordering_depth = 2
   * 
   * Requirement:
   * Unless all beats of transaction 1 are sent out, the beats of 
   * 2nd transactions should not be sent.
   * 
   * Solution:
   * Program the enable_interleave = 0 for both the transaction 1.
   
   */
  rand bit enable_interleave = 0;
  
  /**
    * @groupname axi_protocol
    * When this bit is set , it indicates that this transaction has updated 
    * the AXI Slave memory with write data and other properties.
    */ 
  bit memory_update_complete_for_write =0;

`ifdef SVT_ACE5_ENABLE
 /**
   * @groupname ace5_protocol
   * when this bit is set, it indicates that this transaction 
   * performed atomic operation and the result is stored in atomic_resultant_data.
   */
  bit is_atomic_resultant_data_calculated =0;
`endif 

  /**
   * @groupname ace_protocol
   * When this bit is set by user, it indicates that this transaction is
   * a post-barrier transaction and that it needs to wait for responses
   * from the barrier transaction pair indicated in #associated_barrier_xact.
   * #associated_barrier_xact can be set in the callback
   * svt_axi_master_callback::associate_xact_to_barrier_pair. In this callback,
   * user can associate this transaction with a barrier transaction pair.
   *
   * Please refer to User Guide for more description.
   */
  rand bit associate_barrier = 0;

  /**
   *  @groupname axi3_protocol
   *  Indicates that data will start before address for write transactions.
   *  In data_before_addr scenario (i.e., when data_before_addr = '1'), addr and data channel related delay considerations are: 
   *  1) For programming address_channel related delay: awvalid_delay and reference_event_for_addr_valid_delay are used.
   *   (for more information, look for the description of these variables).
   *    reference_event_for_addr_valid_delay should be set FIRST_WVALID_DATA_BEFORE_ADDR. 
   *    In data_before_addr scenarios reference_event_for_addr_delay should be set very carefully to
   *    FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR as this may cause 
   *    potential deadlock scenarios in SLAVE DUT where slave DUT waits for awvalid signal
   *    before driving wready signal.
   *  2) For programming data_channel related delay: wvalid_delay[] and reference_event_for_first_wvalid_delay & reference_event_for_next_wvalid_delay are used.
   *    (for more information, look for the description of these variables).
   *      For wvalid_delay[0]        -  #reference_event_for_first_wvalid_delay
   *      For remaining indices of wvalid_delay -  #reference_event_for_next_wvalid_delay
   *    In data_before_addr scenario, reference_event_for_first_wvalid_delay must be PREV_WRITE_DATA_HANDSHAKE, otherwise it will cause failure.
   *  .
   *    
   */
  rand bit data_before_addr = 0;
  
  /**
   *  @groupname axi3_protocol
   *  Indicates that data will start before address for write transactions,
   *  even though data_before_addr is set to 0. This is useful when
   *  awvalid is suspended for write transaction and respective transaction
   *  data is driven before resuming the suspended awvalid signal.
   */
  bit suspend_awvalid_to_data_before_addr = 0;

  /**
    * Indicates if the current data beat of a write transaction has wlast
    * asserted. This is useful when data is received before addr and it is
    * required to determine the last beat. This is a sticky bit  in that
    * it remains set to 1 after the last data beat.
    */ 
  bit is_last_write_data_beat = 0;

   // AXI 4 Variables

  /**
   *  @groupname axi4_protocol
   *  The variable holds the value for AWQOS/ARQOS 
   */
  rand bit[`SVT_AXI_QOS_WIDTH - 1:0] qos = 0;  
  

  /**
   *  @groupname axi4_protocol
   *  The variable holds the value for AWREGION/ARREGION
   */
  rand bit[`SVT_AXI_REGION_WIDTH - 1:0] region = 0;


  /**
   *  @groupname axi3_protocol
   *  The variable holds the value for signals AWUSER/ARUSER.
   *  Applicable for all interface types. Enabled through port configuration
   *  parameters svt_axi_port_configuration::aruser_enable and
   *  svt_axi_port_configuration::awuser_enable.
   */
  rand bit[`SVT_AXI_MAX_ADDR_USER_WIDTH - 1:0] addr_user = 0;

  /**
   *  @groupname axi3_protocol
   *  The variable holds the value for signals WUSER/RUSER. Applicable for all
   *  interface types. Enabled through port configuration parameters
   *  svt_axi_port_configuration::wuser_enable and
   *  svt_axi_port_configuration::ruser_enable.
   */
  rand bit[`SVT_AXI_MAX_DATA_USER_WIDTH - 1:0] data_user[];

`ifdef SVT_ACE5_ENABLE
  /**
   *  @groupname ace5_protocol
   *  The variable holds the value for signals RUSER.
   *  Applicable only if svt_axi_port_configuration::atomic_transactions_enable is set to1.
   *  Enabled through port configuration parameters
   *  svt_axi_port_configuration::ruser_enable.
   */
  rand bit[`SVT_AXI_MAX_DATA_USER_WIDTH - 1:0] atomic_read_data_user[];
`endif

   /**
   *  @groupname axi3_protocol
   *  The variable holds the value for signals WUSER/RUSER as they are driven on the bus
   *  Applicable for all interface types. Enabled through port configuration parameters
   *  svt_axi_port_configuration::wuser_enable and
   *  svt_axi_port_configuration::ruser_enable.
   */
   bit[`SVT_AXI_MAX_DATA_USER_WIDTH - 1:0] physical_data_user[];
 /**
   *  @groupname axi3_protocol
   *  The variable holds the value for signal BUSER. Applicable for all
   *  interface types. Enabled through port configuration parameter
   *  svt_axi_port_configuration::buser_enable.
   */
  rand bit[`SVT_AXI_MAX_BRESP_USER_WIDTH - 1:0] resp_user = 0;
  
  /** 
   * @groupname ace_protocol
   * This variable represents the shareability domain of coherent transactions.
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to
   * AXI_ACE or ACE_LITE.
   */
  rand xact_shareability_domain_enum domain_type = NONSHAREABLE;

  /**
   * @groupname ace_protocol
   * This variable represents barrier transaction type. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
   */
  rand barrier_type_enum barrier_type = NORMAL_ACCESS_RESPECT_BARRIER;

  /** 
   * @groupname ace_protocol
   * This variable represents the shareable coherent transaction types. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
   */
  rand coherent_xact_type_enum coherent_xact_type = READNOSNOOP;

`ifdef SVT_ACE5_ENABLE
 /**
  * @groupname ace5_protocol 
  * This variable represents the cmo on the write channel.
  * Applicable when svt_axi_port_configuration::axi_interface_type is set to ACE_LITE.
  */
  rand cmo_on_write_xact_type_enum cmo_on_write_xact_type = CLEANSHARED_ON_WRITE;
`endif

  /** 
   * @groupname ace_protocol
   * Array for the coherent read responses. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  rand coherent_resp_type_enum coh_rresp[];

  /**
    * @groupname ace_status
    * This variable represents the initial cache line state. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or
    * ACE_LITE.  The initial cache line state of a transaction that is driven on
    * the READ channel is populated just after the reception of the first beat
    * of the response of a transaction.  The initial cache line state of a
    * transaction that is driven on the WRITE channel is populated just before
    * the transaction is started. This variable is updated by the VIP, and is a
    * read-only variable. User is not expected or supposed to modify this variable.
    *
    * Applicable for ACTIVE MASTER only.
    */
   cache_line_state_enum initial_cache_line_state = INVALID;

  /**
    * @groupname ace_status
    * This variable represents the prefinal cache line state. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or
    * ACE_LITE.  The prefinal cache line state of a transaction is the state of the 
    * cache  just before cache is updated . This variable is updated by the VIP, and is a
    * read-only variable. User is not expected or supposed to modify this variable.
    *
    * Applicable for ACTIVE MASTER only.
    */
   cache_line_state_enum  prefinal_cache_line_state = INVALID;

   /*
    * @groupname ace_status
    * This variable represents the initial data in the cache. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or
    * ACE_LITE. For transactions driven on the READ channel, this field is 
    * populated just after the reception of the the first beat of the response
    * of the transaction.
    * For transactions driven on the WRITE channel, this is populated just
    * before the transaction is started.
    *
    * Applicable for ACTIVE MASTER only.
    */
   bit[7:0] initial_cache_line_data[];

  /**
    * @groupname ace_status
    * This variable represents the final cache line state. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or
    * ACE_LITE.  The final cache line state of a transaction is the state of the
    * the line just before the transaction ended. This variable is updated by
    * the VIP, and is a read-only variable. User is not expected or supposed to
    * modify this variable.
    *
    * Applicable for ACTIVE MASTER only.
    */
   cache_line_state_enum final_cache_line_state = INVALID;

  /**
    * @groupname ace_status
    * This variable represents the final cache line data. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    * The final cache line data of a transaction is the data of the
    * the line just before the transaction ended. 
    *
    * Applicable for ACTIVE MASTER only.
    */
   bit[7:0] final_cache_line_data[];

  /**
   * @groupname ace_protocol
   * Indicates that the data as given in #cache_write_data in this transaction 
   * needs to be allocated in the cache. Applicable only when transaction type
   * is READUNIQUE or CLEANUNIQUE.
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   *
   * Applicable for ACTIVE MASTER only.
   */
  rand bit allocate_in_cache;

  /**
   * @groupname ace_protocol
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   *
   * Represents data that needs to be stored to the cache if the 
   * #allocate_in_cache bit is set for a READUNIQUE/CLEANUNIQUE transaction 
   * or if the transaction is MAKEUNIQUE.
   * Applicable to masters in active mode.
   * Refer section 3.6 of ACE specification.
   * Writes in ACE are performed by removing all other copies
   * of the cache line so that the master that is performing the write has
   * a unique copy at the time of writing. Depending on whether a paritial
   * or full update of a cache line is required a transaction such as
   * READUNIQUE,MAKEUNIQUE or CLEANUNIQUE is sent. Some of these transactions
   * such as READUNIQUE will return data (either from memory or the cache of
   * some other master) and this will be available in the data[] field of this
   * class. Other transactions such as MAKEUNIQUE and CLEANUNIQUE will not
   * return any data. 
   * For a READUNIQUE transaction, if the #allocate_in_cache bit is not set, the
   * data available in data[] is written in cache. If the #allocate_in_cache bit
   * is set the data available in this variable is written to cache. Note however,
   * that this variable is overwritten by the data that is received in data[] prior
   * to writing in the cache. This is done because READUNIQUE is used for partial update 
   * of a cacheline when a master does not have a copy of the cacheline. So a user 
   * can actually populate this variable after a copy of this cacheline is received and 
   * not at the time of randomization.
   * For a CLEANUNIQUE transaction, if the #allocate_in_cache bit is set,
   * the data in this variable is written to cache. 
   * For a MAKEUNIQUE transaction, the data in this variable is always written into
   * the cache.
   * Updating this variable is normally done in the pre_cache_update callback issued 
   * by the master driver after all the responses are received but prior to the 
   * RACK signal being driven.
   * An important aspect of this variable is that this data is not driven
   * on the physical bus.
   * 
   * Applicable for ACTIVE MASTER only.
   */
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] cache_write_data[];

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
    *
    * Indicates if update of cache must be bypassed for this transaction. A
    * typical use model is to set this bit in pre_cache_update callback of the
    * driver based on response received in the transaction. For example, if the
    * response received is SLVERR, user may not want the driver to update the
    * cache.  When using this property, it is the user's responsibility that
    * system coherency is not lost, since cache will not be updated.
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit bypass_cache_update = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates if the transaction ended because the requested data was already
    * available in the cache. This bit is set by the master, no action is taken
    * if the user sets this bit. A transaction with this bit set was not sent out
    * on the bus and therefore other components in the testbench will not detect
    * this transaction. 
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit is_cached_data = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
    *
    * Indicates if a coherent transaction was dropped because the start state
    * of the corresponding cache line is not as expected before transmitting the
    * transaction. The expected start states for each of the transaction types
    * are given in section 5 of the ACE specification.
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit is_coherent_xact_dropped = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates if the transaction is a result of a speculative read operation.
    * A speculative read is defined as a read of a cache line that a master already
    * holds in its cache.
    *
    * This is a read-only member, which VIP uses to indicate whether the
    * transaction is a speculative read. Modifying the value of this member will
    * not have any effect.
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit is_speculative_read = 0;

  /** @cond PRIVATE */
  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates whether the memory update at slave end for overlapped write
    * transactions should happen in request order.
    *
    * This is a read-only member, which VIP uses to update slave memory for 
    * overlapped write transactions. It should not be modified by the user.
    * 
    * Applicable for ACTIVE SLAVE only.
    */
  bit update_mem_in_req_order = 0;  

  /**
    * @groupname ace_protocol
    * Indicates whether the required checks for WriteUnique and WriteLineUnique
    * not being in progress while a WRITEBACK/WRITECLEAN is in progress is done
    * Applicable when port_interleaving_enable is set in the configuration.
    */
  bit is_wu_wlu_restriction_check_done = 0;

  /**
    * @groupname ace_protocol
    * Indicates whether the required checks for memory update transaction 
    * relative to the cache states are performed just prior to start
    * of this transaction
    */
  bit is_mem_update_pre_xact_xmit_check_done = 0;
  /** @endcond */

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates if the transaction is auto generated by the VIP. Transactions
    * are auto-generated when:
    * 1. The cache is full and an entry needs to be evicted from the cache. 
    * 2. User supplies a cache maintenance transaction and the protocol requires
    * that the cache line is first written into memory before sending the cache
    * maintenance transaction. 
    *
    * This is a read-only member, which VIP uses to indicate whether the
    * transaction is auto generated. It should not be modified by the user. 
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit is_auto_generated = 0;

  /**
    * @groupname ace_protocol
    * Applicable when svt_axi_port_configuration::axi_interface_type is set
    * to AXI_ACE and svt_axi_port_configuration::snoop_response_data_transfer_mode 
    * is set to SNOOP_RESP_DATA_TRANSFER_USING_WB_WC.
    *
    * Indicates if this transaction is a WRITEBACK/WRITECLEAN auto-generated transaction
    * which was generated to transfer snoop data. When 
    * svt_axi_port_configuration::snoop_response_data_transfer_mode is set to 
    * SNOOP_RESP_DATA_TRANSFER_USING_WB_WC, snoop data from a dirty line is transferred
    * using a WRITEBACK/WRITECLEAN transaction instead of the snoop data channel. All
    * transactions which have this variable set will also have  is_auto_generated set.
    */
  bit is_xact_for_snoop_data_transfer = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    * Indicates if the cache line state needs to be forced to a shared state even
    * if the actual state of the line is unique, since it is permissible for
    * a cache line which is in the unique state to be held in the shared state. 
    * Valid only when:
    * svt_axi_port_configuration::cache_line_state_change_type is set to
    * LEGAL_WITH_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE or
    * LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE.
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand bit force_to_shared_state = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    * Indicates if the cache line state needs to be forced to an invalid state even
    * if that is not the recommended state, since it is permissible for
    * a cache line which is in a clean state to be held in the invalid state. 
    * Valid only when:
    * svt_axi_port_configuration::cache_line_state_change_type is set to
    * LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE.
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand bit force_to_invalid_state = 0;

  /**
    * @groupname ace_protocol
    * Applicable when svt_axi_port_configuration::axi_interface_type is set to
    * AXI_ACE or ACE_LITE.  Forces transactions which are not constrained to be
    * of cacheline size by protocol to be of cacheline size. Currently
    * applicable only to READONCE, WRITEUNIQUE, WRITENOSNOOP and READNOSNOOP
    * transactions. Applicable to WRITENOSNOOP and READNOSNOOP only when
    * svt_axi_port_configuration::update_cache_for_non_coherent_xacts is set and
    * svt_axi_port_configuration::axi_interface_type is AXI_ACE.
    * If this bit is set, READONCE and WRITEUNIQUE transactions will be forced
    * to cache line size transactions.
    * This has a dependency on svt_axi_port_configuration::force_xact_to_cache_line_size_interface_type. 
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand bit force_xact_to_cache_line_size = 0;
  
  /**
   * @groupname ace_protocol
   * The variable represents ARVMIDEXT when svt_axi_port_configuration::axi_interface_type 
   * is set to AXI_ACE or ACE_LITE with svt_axi_system_configuration::DVMV8_1 or above.
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_VMIDEXT_WIDTH. Default value of this macro is 4 based on DVMv8.1 architecture recomendation.
   * 
   */

  rand bit [`SVT_AXI_MAX_VMIDEXT_WIDTH - 1:0] arvmid = 0;

  /**
   * @groupname ace5_protocol
   * This variable stores the data check parity bit's with respect to valid data,
   * Each bit of parity check data is calculated from every 8bit of data.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] datachk_parity_value[] ;

  /**
   * @groupname ace5_protocol
   * This variable stores the data check parity error bit's with respect to valid data,
   * Each bit of parity check data is calculated from every 8bit of data with 1bit if datachk.
   * By default all bits are set to 'b1, if any parity error is detected the that particular bit is set to 0.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] is_datachk_passed[] ;

  /**
   * @groupname ace5_protocol
   * This variable represents the data check parity error is deducted in a
   * transaction.
   * In a transaction if parity error is deducted, the this bit is set to 1.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit is_datachk_parity_error = 0;
`ifdef SVT_ACE5_ENABLE
 /**
   * @groupname ace5_protocol
   * This variable stores the data check parity bit's with respect to valid data,
   * Each bit of parity check data is calculated from every 8bit of data.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] atomic_read_datachk_parity_value[] ;

  /**
   * @groupname ace5_protocol
   * This variable stores the data check parity error bit's with respect to valid data,
   * Each bit of parity check data is calculated from every 8bit of data with 1bit if datachk.
   * By default all bits are set to 'b1, if any parity error is detected the that particular bit is set to 0.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] atomic_read_is_datachk_passed[] ;

  /**
   * @groupname ace5_protocol
   * This variable represents the data check parity error is deducted in a
   * transaction.
   * In a transaction if parity error is deducted, the this bit is set to 1.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit atomic_read_is_datachk_parity_error = 0;

  /**
   * - @groupname ace5_protocol 
   * - Field that indicates type of Atomic transaction.
   * - This is a read-only field for the testbench, and is set by the VIP components
   * .
   */
  rand atomic_transaction_type_enum atomic_transaction_type = NON_ATOMIC;

 /**
  * - @groupname ace5_protocol
  * - Field that indicates type of write_with_cmo_xact_type.
  * .
  */

  rand write_with_cmo_xact_type_enum write_with_cmo_xact_type = WRITENOSNPFULL_CLEANSHARED; 

 /**
   * - @groupname ace5_protocol 
   * - Field that indicates type of Atomic transaction.
   * - This is a read-only field for the testbench, and is set by the VIP components
   * .
   */
  rand atomic_xact_op_type_enum atomic_xact_op_type = ATOMICSTORE_ADD;

`endif
 /**
   * @groupname ace5_protocol 
   *This field indicates the value of trace_tag
   */
  rand bit trace_tag =0;

  /**
   * @groupname ace5_protocol
   * This field indicates the value of data trace_tag on write data channel and read data channel
   */
  rand bit data_trace_tag =0;

  /**
   * @groupname ace5_protocol
   * This field indicates the value of btrace on write response channel
   */
  rand bit resp_trace_tag =0;

`ifdef SVT_ACE5_ENABLE 
  /** Internal field to store the atomic data trace_tag for inbound data */
  rand bit atomic_read_data_trace_tag;

 /** 
   * @groupname ace5_protocol
   * This field indicates the node ID of the stash target. 
   * Applicable only in stash type transactions.
   */
  rand bit[(`SVT_AXI_STASH_NID_WIDTH-1):0] stash_nid = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field indicates the stash_nid field has a valid Stash target value.
   * Applicable only in stash type transactions.
   */
  rand bit stash_nid_valid = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field  indicates the ID of the logical processor at the Stash target.
   * Applicable only in stash type transactions.
   */
  rand bit [(`SVT_AXI_STASH_LPID_WIDTH-1):0] stash_lpid = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field indicates that the Stash_lpid field value must be 
   * considered as the Stash target.
   * Applicable only in stash type transactions.
   */
  rand bit stash_lpid_valid = 0;

 /** 
   * @groupname ace5_protocol
   * This field indicates the ID of the stream.This si used to identify the stream.
   * Applicable only when untranslated transaction feature is supported.
   */
  rand bit [(`SVT_AXI_MAX_MMUSID_WIDTH-1):0] stream_id = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field indicates wether the stream is secure or non-secure.
   * When set to 1, indicates a secure stream.
   * Applicable only when untranslated transaction feature is supported.
   */
  rand bit secure_or_non_secure_stream = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field  is only vaid if sub_stream_id_valid is set to 1.
   * This indicates the ID of the sub stream.
   * Applicable only when untranslated transaction feature is supported.
   */
  rand bit[(`SVT_AXI_MAX_MMUSSID_WIDTH-1):0] sub_stream_id = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field indicates that the transaction has an optional substream identifier.
   * When set to 1 , it means that transaction has a substream identifier.
   * This is used in untranslated transaction feature is enabled.
   */
  rand bit sub_stream_id_valid = 0;

 /** 
   * @groupname ace5_protocol
   * This field indicates that the transaction has already undergone PCIE ATS 
   * translation.
   */
  rand bit addr_translated_from_pcie = 0;

`endif

  /**
   *  Represents port ID. Not currently supported.
   */
  int port_id;

  /**
   *  @groupname axi3_4_ace_timing
   *   This variable stores the cycle information for address valid on read and
   *   write transactions. The simulation clock cycle number when the address
   *   valid is asserted, is captured in this member. This information can be
   *   used for doing performance analysis. VIP updates the value of this member
   *   variable, user does not need to program this variable.
   */
  int addr_valid_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for data valid on read and
   *  write transactions. The simulation clock cycle number when the data
   *  valid is asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int data_valid_assertion_cycle[];
`ifdef SVT_ACE5_ENABLE
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for data valid on read and
   *  write transactions. The simulation clock cycle number when the data
   *  valid is asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int atomic_read_data_valid_assertion_cycle[];
`endif
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for response valid on a write
   *  transaction. The simulation clock cycle number when the write response
   *  valid is asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */
  int write_resp_valid_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for address ready on read and
   *  write transactions. The simulation clock cycle number when the address valid
   *  and ready both are asserted i.e. handshake happens, is captured in this member.
   *  This information can be used for doing performance analysis. VIP updates the
   *  value of this member variable, user does not need to program this variable.
   */
  int addr_ready_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data ready on read and
   *  write transactions. The simulation clock cycle number when the data valid and
   *  ready both are asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int data_ready_assertion_cycle[];
`ifdef SVT_ACE5_ENABLE
 /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data ready on read and
   *  write transactions. The simulation clock cycle number when the data valid and
   *  ready both are asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int atomic_read_data_ready_assertion_cycle[];
`endif
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for response ready on a write
   *  transaction. The simulation clock cycle number when the write response valid and
   *  ready both are asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int write_resp_ready_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *   The simulation time when the master or slave driver receives
   *   the transaction from the sequencer, is captured in this member.
   *   This information can be used for doing performance analysis.
   *   VIP updates the value of this member
   *   variable, user does not need to program this variable.
   */

  realtime xact_consumed_by_driver_time;
 /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for address wakeup of read or write 
   *  transaction. The simulation clock cycle number when the address wakeup is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member variable,
   *  user does not need to program this variable.
   */
  int addr_wakeup_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for address wakeup of read or write
   *  transaction. The simulation time when the address wakeup is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member variable,
   *  user does not need to program this variable.
   */
  real addr_wakeup_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for wakeup of idle read or write
   *  channel. The simulation time when the wakeup is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member variable,
   *  user does not need to program this variable.
   */
  real idle_chan_wakeup_toggle_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for wakeup of idle read or write
   *  channel. The simulation time when the wakeup is
   *  deasserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member variable,
   *  user does not need to program this variable.
   */
   real idle_chan_wakeup_toggle_deassertion_time;

 /**
   *   @groupname axi3_4_ace_timing
   *   This variable stores the transaction consumed at driver timing
   *   information. The transaction consumed at driver time to begin time
   *   delay is calculated as the difference between begin_time and
   *   xact_consumed_by_driver_time.
   *   This information can be used for doing performance analysis.
   *   VIP updates the value of this member variable,
   *   user does not need to program this variable.
   */

  real xact_consumed_time_to_begin_time_delay;
  
  /**
   *  @groupname axi3_4_ace_timing
   *   This variable stores the timing information for address valid on read and
   *   write transactions. The simulation time when the address valid is
   *   asserted, is captured in this member. This information can be used for
   *   doing performance analysis. VIP updates the value of this member
   *   variable, user does not need to program this variable.
   */

  real addr_valid_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data valid on read and
   *  write transactions. The simulation time when the data valid is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real data_valid_assertion_time[];
`ifdef SVT_ACE5_ENABLE
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data valid on read and
   *  write transactions. The simulation time when the data valid is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real atomic_read_data_valid_assertion_time[];
`endif
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for response valid on  write
   *  transactions. The simulation time when the response valid is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real write_resp_valid_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for address ready on read and
   *  write transactions. The simulation time number when the address valid and
   *  ready both are asserted i.e. handshake happens, is captured in this member.
   *  This information can be used for doing performance analysis. VIP updates the
   *  value of this member variable, user does not need to program this variable.
   */

  realtime addr_ready_assertion_time;


  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data ready on read and
   *  write transactions. The simulation time when the data valid and ready both are
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real data_ready_assertion_time[];
`ifdef SVT_ACE5_ENABLE
   /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data ready on read and
   *  write transactions. The simulation time when the data valid and ready both are
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real atomic_read_data_ready_assertion_time[];
`endif
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for response ready on  write
   *  transactions. The simulation time when the response valid and ready both are
   *  asserted, is captured in this member. This information can be used for doing
   *  performance analysis. VIP updates the value of this member variable, user
   *  does not need to program this variable.
   */

  real write_resp_ready_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for the data channnel blocking ratio.
   *  The blocking cycle for a beat is defined as the number of cycles that
   *  valid was asserted, but corresponding ready was not asserted.
   *  This ratio is derived from data_valid_assertion_cycle and
   *  data_ready_assertion_cycle, calculated as sum of data ready
   *  blocking cycles divided by sum of data valid assertion cycles.
   *  This information can be used for doing performance analysis.
   *  VIP updates the value of this member variable, user
   *  does not need to program this variable.
   */
  real data_chan_blocking_ratio;

  // ****************************************************************************
  // Members relevant to Master Driver and Monitor  
  // ****************************************************************************

  /**
    * @groupname axi3_4_delays
    * This variable defines the number of cycles the AWVALID or ARVALID  signal is
    * delayed. The reference event for this delay is #reference_event_for_addr_valid_delay.
    * Applicable for ACTIVE MASTER only.
    */
  rand int addr_valid_delay = 0;
   
  /**
    * @groupname axi3_4_delays
    * Defines a reference event from which the AWVALID or ARVALID delay
    * should start.  Following are the different reference events:
    *
    * PREV_ADDR_VALID:  
    * Reference event is the previous AWVALID or ARVALID signal 
    *
    * PREV_ADDR_HANDSHAKE:  
    * Reference event is previous read or write Address handshake
    *
    * FIRST_WVALID_DATA_BEFORE_ADDR:
    * This is used when #data_before_addr bit is set. The reference event for
    * address valid to occur is the first wvalid of the current transaction.
    *
    * FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR:
    * This is used when #data_before_addr bit is set. The reference event for
    * address valid to occur is the first data handshake of the current transaction.
    *
    * PREV_LAST_DATA_HANDSHAKE:
    * Reference event is previous read or write last data handshake
    * to Address valid assertion.
    *
    * Reasonable constraint on reference_event_for_addr_delay in data_before_addr scenarios is added in svt_axi_transaction class 
    * to constraint the value of reference_event_for_addr_delay not to take FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR.
    * User may swicth off the constraint reasonable_reference_event_for_addr_delay by setting rand_mode to 0 
    * incase they want reasonable_reference_event_for_addr_delay to take FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR.
    * In data_before_addr scenarios reference_event_for_addr_delay should be set very carefully to
    * FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR as this may cause 
    * potential deadlock scenarios in ACE SLAVE DUT where slave DUT waits for awvalid signal
    * before driving wready signal.
    *
    */
  rand reference_event_for_addr_valid_delay_enum  reference_event_for_addr_valid_delay = PREV_ADDR_HANDSHAKE;


  /**
    * @groupname axi3_4_delays
    * Defines the delay in number of cycles for AWAKEUP signal assertion
    * before or after ARVALID or AWVALID signal.
    */
  rand int awakeup_assert_delay = 0;
  
  /**
    * @groupname axi3_4_delays
    * Defines the delay in number of cycles for AWAKEUP signal deassertion
    * after ARVALID-ARREADY or AWVALID-AWREADY signal handshake.
    */
  rand int awakeup_deassert_delay = 0;

  /** if this bit is set to '0' then AWAKEUP signal will be asserted 
    * before ARVALID with respect to awakeup_assert_delay.
    * if this bit is set to '1' then AWAKEUP signal will be asserted
    * after ARVALID or AWVALID with respect to awakeup_assert_delay.
    */ 
  rand bit assert_awakeup_after_valid = 0;

  /** 
    * @groupname axi3_4_delays
    * Defines the delay in number of cycles for WVALID signal.
    * The reference event for this delay is:
    * - For wvalid_delay[0]        -  #reference_event_for_first_wvalid_delay
    * - For remaining indices of wvalid_delay -  #reference_event_for_next_wvalid_delay
    * .
    * Applicable for ACTIVE MASTER only.
    */
  rand int wvalid_delay[];
   
  /**
    * @groupname axi3_4_delays
    * If configuration parameter #svt_axi_port_configuration::default_rready is
    * FALSE, this member defines the RREADY signal delay in number of clock
    * cycles.  The reference event for this delay is
    * #reference_event_for_rready_delay
    *
    * If configuration parameter #svt_axi_port_configuration::default_rready is
    * TRUE, this member defines the number of clock cycles for which RREADY
    * signal should be deasserted after each handshake, before pulling it up
    * again to its default value.
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand int rready_delay[];

  /**
    * @groupname axi3_4_delays
    * Applicable when svt_axi_port_configuration::toggle_ready_signals_during_idle_period
    * is set. Applicable for master VIP.
    *
    * Indicates the number of cycles for which RREADY should be high and low
    * when the read data channel is idle, that is, when RVALID is low. This
    * property helps to toggle the RREADY signal during the idle period between
    * the assertion of RVALID signal.  Values provided in even numbered indices
    * indicate the number of clocks for which the ready signal must be driven
    * low and the values in odd numbered indices indicate the number of clocks
    * for which it must driven high. Note that the values provided in this
    * variable are applied for all read data beats. If the user requires a
    * different set of delays during the idle period for each beat, the user
    * must use the read_data_phase_started callback to change the values of
    * this property for the corresponding beat. Once changed, the values will
    * be applicable for all subsequent beats of the transaction unless it is
    * is changed for a subsequent beat. Values in this variable are applicable
    * only until RVALID is asserted. When RVALID is observed on the interface,
    * this delay is no longer applicable. The delay specified in
    * #rready_delay is applied before this property is used.  Note that toggling
    * RREADY during the idle period may lead to situations where the RREADY
    * signal is already asserted when the RVALID is sampled, even though the
    * value of #svt_axi_port_configuration::default_rready is low. Similarly,
    * RREADY may be low when the corresponding valid is sampled, even though
    * the value of #svt_axi_port_configuration::default_rready is high. In both
    * these cases, #rready_delay is not applicable. The size of this array can be
    * set to any value greater than 0, based on the number of times the user
    * would like the signal to toggle during idle period.
    */
  rand int idle_rready_delay[];

  /**
   * @groupname axi4_stream_delays
   * Defines the delay in number of clock cycles for TVALID signal.
   * The reference event for this delay is:  #reference_event_for_tvalid_delay
   * - PREV_TVALID_TREADY_HANDSHAKE : Previous tvalid-tready handshake as the reference event
   * - PREV_TVALID                  : Previous tvalid assertion as the reference event
   * .
   * Applicable for ACTIVE MASTER only.
   */
  rand int tvalid_delay[];

  /**
   * @groupname axi4_stream_delays
   * If configuration parameter #svt_axi_port_configuration::default_tready is
   * FALSE, this member defines the TREADY signal delay in number of clock
   * cycles.  The reference event for this delay is
   * #reference_event_for_tready_delay.
   *
   * Please note that #reference_event_for_tready_delay is not supported
   * currently. Absolute value of tready_delay is considered for delay
   * calculation with respect to tvalid signal.
   *
   * If configuration parameter #svt_axi_port_configuration::default_tready is
   * TRUE, this member defines the number of clock cycles for which TREADY
   * signal should be deasserted after each handshake, before pulling it up
   * again to its default value.
   *
   * Applicable for ACTIVE SLAVE only.
   */
  rand int tready_delay[];

  /**
    * @groupname axi3_4_delays
    * Defines the reference events to delay the first wvalid signal. The delay
    * must be programmed in wvalid_delay[0]. Following are the different
    * events under this category:
    *
    * WRITE_ADDR_VALID:
    * Reference event for first WVALID is assertion of AWVALID signal
    * 
    * WRITE_ADDR_HANDSHAKE:
    * This event is applicable when write data is transmitted after write
    * address, that is, when #data_before_addr is set to 0. This reference event
    * specifies the write address handshake.
    * 
    * PREV_WRITE_DATA_HANDSHAKE:
    * This event is applicable when write data is transmitted before write
    * address, that is, when #data_before_addr is set to 1. This reference event
    * specifies the previous write data handshake.
    */
    // removed address handshake refrence because  of potential deadlock due to following reason::
    // the slave can wait for AWVALID or WVALID, or both before asserting AWREADY
    //
  rand reference_event_for_first_wvalid_delay_enum reference_event_for_first_wvalid_delay =  WRITE_ADDR_VALID;

  /**
    * @groupname axi3_4_delays
    * Defines the reference events for WVALID delay from second beat
    * onwards. Following are the different events under this category:
    *  
    * PREV_WVALID:
    * Reference event for WVALID delay is assertion of previous wvalid.  The
    * delay timer starts as soon as previous valid signal is asserted. If
    * previous data handshake does not complete before timer expires, the
    * current transfer waits for the previous handshake to complete, and then
    * immediately asserts wvalid.
    * 
    * PREV_WRITE_HANDSHAKE:
    * Reference event for WVALID delay is completion of previous data handshake.
    */
  rand reference_event_for_next_wvalid_delay_enum reference_event_for_next_wvalid_delay = PREV_WRITE_HANDSHAKE;

  /**
    *    
    * @groupname axi3_4_delays
    * Defines the reference event for RREADY delay.
    *   
    * RVALID:
    * Reference event for RREADY is assertion of RVALID signal
    * 
    * MANUAL_RREADY: (Not supported currently)
    *
    * This event  allows the user to generate  RREADY patterns, in cycles, as
    * follows:
    * 1. The reference event for this delay is the beginning of the Address
    *    handshake.
    * 2. The rready_delay[0]  represents the following
    *    a. A value > 0 is the no. of cycles default rready signal is
    *       driven
    *    b. A value < 0 is the no. of cycles default rready signal is
    *       driven after toggling
    * 3. The remaining rready_delay element represents no. of cycles to drive
    *    rready
    * 
    * Example 1:
    * For eg.   RREADY  pattern (cycles) =  1110011 and default_rready = 1 
    * data_delay[0] = 3  Three cycles high (driving default_rready value) 
    * data_delay[1] = 2  Two cycles low    (toggled previous RREADY value) 
    * data_delay[2] = 2  Two cycles high   (toggled previous RREADY value)

    * For eg. cycle pattern  RREADY =  0001100 and default_rready = 1 
    * data_delay[0] = -3 Three cycles low (toggled default_rready value) 
    * data_delay[1] = 2  Two cycles high  (toggled previous RREADY value) 
    * data_delay[2] = 2  Two cycles low   (toggled previous RREADY value)
    */
  rand reference_event_for_rready_delay_enum reference_event_for_rready_delay = RVALID;

  /**
    * @groupname axi3_4_delays
    * If configuration parameter #svt_axi_port_configuration::default_bready is
    * FALSE, this member defines the BREADY signal delay in number of clock
    * cycles.  The reference event for this delay is
    * #reference_event_for_bready_delay.
    * 
    * If configuration parameter #svt_axi_port_configuration::default_bready is
    * TRUE, this member defines the number of clock cycles for which BREADY
    * signal should be deasserted after each handshake, before pulling it up
    * again to its default value.
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand int bready_delay = 0;

  /**
    * @groupname axi3_4_delays
    * Applicable when svt_axi_port_configuration::toggle_ready_signals_during_idle_period
    * is set. Applicable for master VIP.
    *
    * Indicates the number of cycles for which BREADY should be high and low
    * when the write response channel is idle, that is, when BVALID is low.
    * This property helps to toggle the BREADY signal during the idle period
    * between the assertion of BVALID signal.  The value for this property may
    * be set when the transaction is randomized at the master or in a callback
    * such as svt_axi_port_monitor_callback::write_resp_phase_started. Values
    * provided in even numbered indices indicate the number of clocks for which
    * the ready signal must be driven low and the values in odd numbered
    * indices indicate the number of clocks for which it must driven high.
    * Values in this variable are applicable only until BVALID is asserted.
    * When BVALID is observed on the interface, this delay is no longer
    * applicable. The delay specified in #bready_delay is applied before this
    * attribute is applied.  Note that toggling BREADY during the idle period
    * may lead to situations where the BREADY signal is already asserted when
    * BVALID is sampled, even though the value of
    * #svt_axi_port_configuration::default_bready is low. Similarly, BREADY may
    * be low when the corresponding valid is sampled, even though the value of
    * #svt_axi_port_configuration::default_bready is high. In both these cases,
    * #bready_delay is not applicable. The size of this array can be set to any
    * value greater than 0, based on the number of times the user would like
    * the signal to toggle during idle period.
    */
  rand int idle_bready_delay[];


  /**
    * @groupname axi3_4_delays
    * Defines a reference event for BREADY delay.
    *
    * BVALID:
    * Reference event is assertion of BVALID signal
    */
  rand reference_event_for_bready_delay_enum reference_event_for_bready_delay = BVALID;

  /**
    * @groupname axi3_4_delays
    * This members applies to AWREADY signal delay for write transactions, and
    * ARREADY signal delay for read transactions.
    *
    * If configuration parameter #svt_axi_port_configuration::default_awready
    * or #svt_axi_port_configuration::default_arready is FALSE, this member
    * defines the AWREADY or ARREADY signal delay in number of clock cycles.
    * The reference event used for this delay is
    * #reference_event_for_addr_ready_delay. 
    *
    * If configuration parameter #svt_axi_port_configuration::default_awready
    * or #svt_axi_port_configuration::default_arready is TRUE, this member
    * defines the number of clock cycles for which AWREADY or ARREADY signal
    * should be deasserted after each handshake, before pulling it up again to
    * its default value.
    *
    * Applicable for ACTIVE SLAVE only.
    */
  rand int addr_ready_delay = 0;

  /**
    * @groupname axi3_4_delays
    * Applicable when svt_axi_port_configuration::toggle_ready_signals_during_idle_period
    * is set. Applicable for slave VIP.
    *
    * Indicates the number of cycles for which awready and arready should be
    * high and low when the corresponding address channel is idle, that is,
    * when AWVALID/ARVALID is low. This property helps to toggle the
    * AWREADY/ARREADY signal during the idle period between the assertion of
    * AWVALID/ARVALID signal of this transaction and the next transaction.
    * This value may be assigned during randomization of the transaction object
    * in the slave sequence. Values provided in even numbered indices indicate
    * the number of clocks for which the ready signal must be driven low and
    * the values in odd numbered indices indicate the number of clocks for
    * which it must driven high. Values in this variable are applicable only
    * until the corresponding valid is asserted. When AWVALID/ARVALID is
    * observed on the interface, this delay is no longer applicable and the
    * delay specified in #addr_ready_delay is applied before asserting
    * AWREADY/ARREADY.  Note that toggling AWREADY/ARREADY during the idle
    * period may lead to situations where the AWREADY/ARREADY signal is already
    * asserted when the corresponding valid is sampled, even though the value
    * of #svt_axi_port_configuration::default_awready or
    * #svt_axi_port_configuration::default_arready is low. Similarly,
    * AWREADY/ARREADY may be low when the corresponding valid is sampled, even
    * though the value of #svt_axi_port_configuration::default_awready or
    * #svt_axi_port_configuration::default_arready is high. In both these
    * cases, #addr_ready_delay is not applicable. The size of this array can be
    * set to any value greater than 0, based on the number of times the user
    * would like the signal to toggle during idle period.
    */
  rand int idle_addr_ready_delay[];


  /** 
    * @groupname axi3_4_delays
    * Defines reference event for AWREADY or ARREADY delay.
    *
    * ADDR_VALID:
    * Reference event is  assertion of AWVALID or ARVALID signal. This event is
    * not applicable when default value of AWREADY = 1 or default value of
    * ARREADY = 1.
    * FIRST_WVALID:
    * Reference event is  assertion of WVALID signal. This event is
    * not applicable when default value of AWREADY = 1.
    * This event is only applicable for write address channel.
    */
  rand reference_event_for_addr_ready_delay_enum  reference_event_for_addr_ready_delay = ADDR_VALID;

  /** 
    * @groupname axi3_4_delays
    * Defines RVALID delay, in terms of number of clock cycles.
    * The reference event for this delay is:
    * - For rvalid_delay[0]        -  #reference_event_for_first_rvalid_delay
    * - For remaining indices of rvalid_delay -  #reference_event_for_next_rvalid_delay
    * .
    *
    * Applicable for ACTIVE SLAVE only.
    */

  rand int rvalid_delay[];

  /**
    * @groupname axi3_4_delays
    * If configuration parameter #svt_axi_port_configuration::default_wready is
    * FALSE, this member defines the WREADY signal delay in number of clock
    * cycles.  The reference event for this delay is
    * #reference_event_for_wready_delay.
    *
    * If configuration parameter #svt_axi_port_configuration::default_wready is
    * TRUE, this member defines the number of clock cycles for which WREADY
    * signal should be deasserted after each handshake, before pulling it up
    * again to its default value. 
    *
    * Applicable for ACTIVE SLAVE only.
    */

  rand int wready_delay[];

  /**
    * @groupname axi3_4_delays
    * Applicable when svt_axi_port_configuration::toggle_ready_signals_during_idle_period
    * is set. Applicable for slave VIP.
    *
    * Indicates the number of cycles for which wready should be high and low
    * when the write data channel is idle, that is, when WVALID is low. This
    * property helps to toggle the WREADY signal during the idle period between
    * the assertion of WVALID signal.  Values provided in even numbered indices
    * indicate the number of clocks for which the ready signal must be driven
    * low and the values in odd numbered indices indicate the number of clocks
    * for which it must driven high. Note that the values provided in this
    * variable are applied for all write data beats. If the user requires a
    * different set of delays during the idle period for each beat, the user
    * must use the write_data_phase_started callback to change the values of
    * this property for the corresponding beat. Once changed, the values will
    * be applicable for all subsequent beats of the transactions unless it is
    * is changed for a subsequent beat. Values in this variable are applicable
    * only until WVALID is asserted. When WVALID is observed on the interface,
    * this delay is no longer applicable and the delay specified in
    * #wready_delay is applied before asserting WREADY.  Note that toggling
    * WREADY during the idle period may lead to situations where the WREADY
    * signal is already asserted when the WVALID is sampled, even though the
    * value of #svt_axi_port_configuration::default_wready is low. Similarly,
    * WREADY may be low when the corresponding valid is sampled, even though
    * the value of #svt_axi_port_configuration::default_wready is high. In both
    * these cases, #wready_delay is not applicable. The size of this array can be
    * set to any value greater than 0, based on the number of times the user
    * would like the signal to toggle during idle period.
    */
  rand int idle_wready_delay[];

  /**
    * @groupname axi3_4_delays
    * Defines the reference events to delay the first rvalid signal. The delay
    * must be programmed in rvalid_delay[0]. Following are the different
    * events under this category:
    *
    * READ_ADDR_VALID:
    * Reference event for first RVALID is assertion of ARVALID signal
    *
    * READ_ADDR_HANDSHAKE:
    * Reference event for first RVALID is completion of read address handshake
    */
  rand reference_event_for_first_rvalid_delay_enum reference_event_for_first_rvalid_delay = READ_ADDR_HANDSHAKE;


  /**
    * @groupname axi3_4_delays
    * Defines the reference events to delay the RVALID signals from second beat
    * onwards. Following are the different events under this category:
    *  
    * PREV_RVALID :
    * Reference event to delay RVALID is assertion of previous rvalid.  The
    * delay timer starts as soon as previous valid signal is asserted. If
    * previous data handshake does not complete before timer expires, the
    * current transfer waits for the previous handshake to complete, and then
    * immediately asserts rvalid.
    * 
    * PREV_READ_HANDSHAKE :
    * Reference event to delay RVALID is completion of previous read data
    * handshake.
    */

  rand reference_event_for_next_rvalid_delay_enum reference_event_for_next_rvalid_delay = PREV_READ_HANDSHAKE;

  /**
    * @groupname axi3_4_delays
    * Defines the reference events for WREADY delay.
    *   
    * WVALID:
    * Reference event for WREADY is assertion of WVALID signal.
    * 
    * MANUAL_WREADY: (Not supported currently)
    * This event  allows the user to generate  WREADY patterns, in cycles, as
    * follows :
    * 1. The reference event for this delay is the beginning of the Address
    *    handshake.
    * 2. The wready_delay[0]  represents the following
    *    a. A value > 0 is the no. of cycles default wready signal is
    *       driven
    *    b. A value < 0 is the no. of cycles default wready signal is
    *       driven after toggling
    * 3. The remaining wready_delay element represents no. of cycles to drive
    *    wready
    * 
    * Example 1:
    * For eg.   WREADY  pattern (cycles) =  1110011 and default_wready = 1 
    * data_delay[0] = 3  Three cycles high (driving default_wready value) 
    * data_delay[1] = 2  Two cycles low    (toggled previous WREADY value) 
    * data_delay[2] = 2  Two cycles high   (toggled previous WREADY value)

    * For eg. cycle pattern  WREADY =  0001100 and default_wready = 1 
    * data_delay[0] = -3 Three cycles low (toggled default_wready value) 
    * data_delay[1] = 2  Two cycles high  (toggled previous WREADY value) 
    * data_delay[2] = 2  Two cycles low   (toggled previous WREADY value)
    */

  rand reference_event_for_wready_delay_enum  reference_event_for_wready_delay =  WVALID;

  /**
    * @groupname axi3_4_delays
    * Defines the BVALID delay in terms of number of clock cycles. The reference
    * event for this delay is #reference_event_for_bvalid_delay.
    *
    * Applicable for ACTIVE SLAVE only.
    */

  rand int bvalid_delay = 0;

  /**
    * @groupname axi3_4_delays
    * Defines a reference event for BVALID delay.
    *
    * LAST_DATA_HANDSHAKE:
    * Reference event for BVALID delay is completion of handshake for last write
    * data.
    * 
    * ADDR_HANDSHAKE:
    * Reference event for BVALID delay is completion of handshake for address phase.
    */  

  rand reference_event_for_bvalid_delay_enum reference_event_for_bvalid_delay = LAST_DATA_HANDSHAKE;

  /**
    * @groupname axi4_stream_delays
    * Defines the reference events for TVALID delay from second beat
    * onwards. Following are the different events under this category:
    *  
    * PREV_TVALID:
    * In this case, assertion of previous tvalid signal is considered  
    * as the reference event for TVALID delay. The delay timer
    * starts as soon as previous tvalid signal is asserted. If previous
    * tvalid-tready handshake does not complete before timer expires, the
    * current transfer waits for the previous handshake to complete, and then
    * immediately asserts tvalid.
    * 
    * PREV_TVALID_TREADY_HANDSHAKE:
    * Reference event for TVALID delay is completion of previous tvalid-tready handshake.
    */
  rand reference_event_for_tvalid_delay_enum reference_event_for_tvalid_delay = PREV_TVALID_TREADY_HANDSHAKE;

  /** 
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   *
   * Defines the reference event from which the RACK delay should start.
   * - LAST_READ_DATA_HANDSHAKE: Reference event is last data handshake
   * .
   */
  rand reference_event_for_rack_delay_enum reference_event_for_rack_delay = LAST_READ_DATA_HANDSHAKE;

  /**
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   * Defines the RACK delay in terms of number of clock cycles. The reference
   * event for this delay is #reference_event_for_rack_delay.
   *
   * Applicable for ACTIVE MASTER only.
   */

  rand int rack_delay = 0;
  
  /** 
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   *
   * Defines the reference event from which the WACK delay should start.
   * - WRITE_RESP_HANDSHAKE: Reference event is last data handshake
   * .
   */
  rand reference_event_for_wack_delay_enum reference_event_for_wack_delay = WRITE_RESP_HANDSHAKE;

  /**
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   * Defines the WACK delay in terms of number of clock cycles. The reference
   * event for this delay is #reference_event_for_wack_delay.
   *
   * Applicable for ACTIVE MASTER only.
   */

  rand int wack_delay = 0;

  /**
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   * Defines the delay between reception of DVM Sync and transmission of DVM Complete.
   * Delay for master component in terms of number of clock cycles for generating
   * DVM Complete transaction after receiving a DVM Sync transaction. 
   *
   * Applicable for ACTIVE MASTER only.
   */

  rand int dvm_complete_delay = 0;

  /**
   *  @groupname out_of_order
   *  Sets the reordering priority of the current transaction within the set
   *  of transactions that are allowed access to read data channel based on 
   *  svt_axi_port_configuration::read_data_reordering_depth.
   * 
   *  This member is applicable only when svt_axi_port_configuration::reordering_algorithm
   *  is svt_axi_port_configuration::PRIORITIZED.
   * 
   *  This value indicates the priority of sending the response to current 
   *  transaction compared to remaining transactions within the depth indicated
   *  by svt_axi_port_configuration::read_data_reordering_depth for read transactions or
   *  by svt_axi_port_configuration::write_resp_reordering_depth for write transactions.
   *
   *  Note that the value of this attribute should be within the following range:
   *  [1:svt_axi_port_configuration::read_data_reordering_depth] for read transactions and
   *  [1:svt_axi_port_configuration::write_resp_reordering_depth] for write transactions.
   * 
   *  If svt_axi_port_configuration::reordering_priority_high_value is set to ‘1’ then, the
   *  transactions with highest value for this attribute will get higher priority.
   *
   *  If svt_axi_port_configuration::reordering_priority_high_value is set to ‘0’ then, the
   *  transactions with least value for this attribute will get higher priority.
   *
   *  If there are more than one transactions with same priority, those transaction
   *  will be processed in the same order as they are received.
   * 
   * Applicable for ACTIVE SLAVE only.
   */

  rand int reordering_priority = 1;

   /**
     * @groupname axi3_4_delays
     * Weight used to control distribution of zero delay within transaction generation.
     *
     * This controls the distribution of delays for the 'delay' fields 
     * (e.g., delays for asserting the ready signals).
     */
  int ZERO_DELAY_wt = 100;

   /**
     * @groupname axi3_4_delays
     * Weight used to control distribution of short delays within transaction generation.
     *
     * This controls the distribution of delays for the 'delay' fields 
     * (e.g., delays for asserting the ready signals).
     */
  int SHORT_DELAY_wt = 500;

  /**
    * @groupname axi3_4_delays
    * Weight used to control distribution of long delays within transaction generation.
    *
    * This controls the distribution of delays for the 'delay' fields 
    * (e.g., delays for asserting the ready signals).
    */
  int LONG_DELAY_wt = 1;


   /**
     * @groupname axi3_protocol
     * Weight used to control distribution of burst length to 1 within transaction
     * generation.
     *
     * This controls the distribution of the length of the bursts using
     * burst_length field 
     */
  int ZERO_BURST_wt = 100;

   /**
     * @groupname axi3_protocol
     * Weight used to control distribution of short bursts within transaction
     * generation.
     *
     * This controls the distribution of  the length of the bursts using
     * burst_length field 
     */
  int SHORT_BURST_wt = 500;


   /**
     * @groupname axi3_protocol
     * Weight used to control distribution of longer bursts within transaction
     * generation.
     *
     * This controls the distribution of  the length of the bursts using
     * burst_length field 
     */
  int LONG_BURST_wt = 400;


  // ****************************************************************************
  // STREAM SIGNALS
  // ****************************************************************************

   /**
    * @groupname axi4_stream_protocol
    * Used to drive TDATA signals. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */
   rand bit [`SVT_AXI_MAX_TDATA_WIDTH - 1:0] tdata[];

  
  /**
   * @groupname axi4_stream_protocol
   * Used to drive TSTRB signal. The strobes are right aligned and the model
   * will drive strobes on appropriate lanes. The model also takes care of the
   * endianness while driving tstrb. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
   */
  rand bit [`SVT_AXI_TSTRB_WIDTH - 1:0] tstrb[];

 
  /**
   * @groupname axi4_stream_protocol
   * TKEEP is the byte qualifier that indicates whether the content of the
   * associated byte of TDATA is processed as part of the data stream.
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to
   * AXI4_STREAM.
   */
  rand bit [`SVT_AXI_TKEEP_WIDTH - 1:0] tkeep[];


  /**
    * @groupname axi4_stream_protocol
    * The variable holds the value of  TID signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */
  rand bit [`SVT_AXI_MAX_TID_WIDTH - 1:0] tid = 0;
  
  /**
    * @groupname axi4_stream_protocol
    * TDEST provides routing information for the data stream. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */

  rand bit [`SVT_AXI_MAX_TDEST_WIDTH - 1:0] tdest;
  
  /**
    * @groupname axi4_stream_protocol
    * TUSER is user defined sideband information that can be transmitted
    * alongside the data stream. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */

  rand bit [`SVT_AXI_MAX_TUSER_WIDTH - 1:0] tuser[];

  /**
    * @groupname axi4_stream_protocol
    * Defines the burst length of a AXI4 Stream Packet. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */
  rand int stream_burst_length = 1;

  // ****************************************************************************
  // End of STREAM SIGNALS
  // ****************************************************************************
  /**
    * @groupname axi3_protocol
    * A bit that must be set by the user to indicate that this transaction will
    * be sent to the slave driver from the slave sequencer through the
    * delayed_response_request_port of the slave driver. If the transaction is
    * randomized before putting it into the delayed_response_request_port of the
    * slave driver, then this bit must be set by the user. This bit must not be
    * set for a transaction that is sent on the seq_item_port.
    */
  bit is_delayed_response_xact = 0;

  /**
   * @groupname axi_misc
   * Indicates the value of the source master which will be propogated in the ID field
   * of the master and the corresponding slave transaction.
   * Applicable for users who want to correlate master transactions to slave
   * transactions in the system monitor. This parameter is applicable when
   * svt_axi_port_configuration::source_master_id_xmit_to_slaves_type is set to
   * DYNAMIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES. This property must be set by the
   * user in a system monitor callback issued at the start of a transaction
   */
  bit[`SVT_AXI_DYNAMIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES_WIDTH-1:0] dynamic_source_master_id_xmit_to_slaves = 0;

  /**
   * @groupname axi_misc
   * Indicates that this master transaction is a partial write transaction and this
   * transaction will be split by the interconnect into a full Read transaction
   * followed by partial Write transaction to the corresponding slave.
   * Applicable for users who want to correlate master transactions to slave
   * transactions in the system monitor. This parameter is applicable when
   * svt_axi_port_configuration::partial_write_to_slave_read_and_write_association_enable is set to
   * This property must be set by the user in a system monitor callback issued at the start of a transaction
   */
  bit partial_master_write_split_into_read_modified_write_slave_xact = 0;

  /**
   * @groupname axi_misc
   * Multibit array for different usages.
   * 
	 * If cust_xact_flow[0] is set to '1', indicate that transaction should be drived immediately on the interface.
	 * This is aplicable only for AXI4 STREAM transactions.
	 *
	 * cust_xact_flow[31:1] bits are for future use.
   */
  rand bit[31:0] cust_xact_flow = 0;  

  /** @cond PRIVATE */
  /**
    * @groupname axi3_protocol
    * A bit that is set by the slave driver to indicate that the write response
    * of a transaction has been provided by the user through the
    * delayed_response_request_port of the slave driver.  
    * Applicable only when
    * svt_axi_port_configuration::enable_delayed_response_port is set.
    */
  bit is_delayed_write_response_set = 0;

  /** 
    * @groupname ace_l3_cache
    * Inidcates that current transaction will cause memory update transaction for the associated
    * cacheline if it is  hit in L3 and found to be in dirty state.
    */
  bit clean_l3_data = 0;

  /** 
    * @groupname ace_l3_cache
    * This attribute is supposed to be updated by VIP indicating to the user that memory has been
    * updated for the current transaction with associated cacheline data in L3 cache. This is primarily
    * used along with clean_l3_data i.e. if current transaction is expected to update memory then user
    * can wait for this attribute to be set by VIP if user needs to perform any tasks based on that condition.
    */
  bit mem_updated_with_l3_data = 0;
  /** @endcond */

  `ifdef SVT_ACE5_ENABLE  
  /**
    * @groupname axi5_protocol
    * Defines the chunk enable of a AXI5 to enable read_data_chunking. When enable, slave will send read data
    * in 128bits of chunk in random order. If disabled, slave will send read data without chunking as per AXI5 protocol. Applicable 
    * when svt_axi_port_configuration::rdata_chunking_enable is set to 1.
    * Not yet implemented. 
    */
  rand bit archunken = 0;

  /**
    * @groupname axi5_protocol
    * Array of read chunk strobe
    * Each bit of rchunkstrb represents 128bits of read data. Width of the rchunkstrb by default is 
    * `SVT_AXI_MAX_CHUNK_STROBE_WIDTH user can change width using svt_axi_port_configuration::rchunkstrb_width 
    * signal. Applicable when archunken and svt_axi_port_configuration::rdata_chunking_enable is set to 1.
    * Not yet implemented. 
    */
  rand bit [`SVT_AXI_MAX_CHUNK_STROBE_WIDTH -1 : 0] rchunkstrb[];

  /**
    * @groupname axi5_protocol
    * Array of read chunk number
    * Indicates that the data chunk number is being transferred. Width of the rchunknum by default is 
    * `SVT_AXI_MAX_CHUNK_NUM_WIDTH user can change width using svt_axi_port_configuration::rchunknum_width 
    * signal. Applicable when archunken and svt_axi_port_configuration::rdata_chunking_enable is set to 1.
    * Not yet implemented. 
    */
  rand bit [`SVT_AXI_MAX_CHUNK_NUM_WIDTH -1 : 0] rchunknum[];

  /**
    * @groupname axi5_protocol
    * Indicates that the data chunk length is being transferred. This signal is for interal use to calculate number  
    * of transafer for chunkinig Applicable when archunken and svt_axi_port_configuration::rdata_chunking_enable 
    * is set to 1.
    * Not yet implemented. 
    */
  rand int chunk_length;

  /**
   * @groupname axi5_protocol
   *    This is a counter which is incremented for every chunk of databeat. Useful when user
   *    would try to access the transaction class to know its current state during chunking.
   *    This represents the chunk databeat transfer number.
   */
  int  current_data_chunk_trf_num = 0;
  `endif  

  // ****************************************************************************
  // STREAM SIGNALS
  // ****************************************************************************

  `ifdef SVT_AXI_QVN_ENABLE
  /**
   * @groupname qvn_parameters
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to AXI3/AXI4/ACE/ACE_LITE
   * Specifies the Virtual Network ID to which token for this transaction will be requested.
   * Same Virtual Network will be used to send current transaction as well. 
   *
   * Active Master will use qvn_vnet_id to determine which VN*VALID* signal needs to be asserted
   * to request for token and all ARVNET_ID or AWVNET_ID and WVNET_ID value will be driven
   * same as qvn_vnet_id
   *
   * Port Monitor will use qvn_vnet_id to indicate from which Virtual Network this particular 
   * transaction has been received.
   *
   */
  rand int qvn_vnet_id = 0;
  `endif

  `ifdef SVT_AXI_CUSTNV_ENV
  /** 
    * configuration register used to provide custom L3 or interconncet based behaviour
    * [0] = '1' indicates writeEvict can start from shared state.
    * [1] = '1' indicates no data has been provided as part of the read response.
    * [2] = '1' indicates current transaction is a block linear request.
    * [3] = '1' indicates current transaction is auto-generated by VIP for an origninal block linear request.
    *           this bit is supposed to get set by VIP. User doesn't need to set this bit.
    *
    * default value of all fields are 0 and it is set by user except bit[3].
    */
  bit[31:0] custnv_reg = 0;
  `endif
  
  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  local static vmm_log shared_log = new("svt_axi_transaction", "class" );
`endif

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
  local svt_axi_port_configuration::axi_port_kind_enum axi_port_kind = svt_axi_port_configuration::AXI_MASTER;

  local svt_axi_port_configuration::axi_interface_type_enum axi_interface_type = svt_axi_port_configuration::AXI3; 
`endif

  /** @cond PRIVATE */
  /** Helper attribute for randomization calculated during pre_randomize */
  protected int log_base_2_data_width_in_bytes = 0;
  
  /** Helper attribute for randomization calculated during pre_randomize */
  protected int data_width_in_bytes = 0;
 
  /** Helper attribute for randomization calculated during pre_randomize */
  protected bit[`SVT_AXI_MAX_DATA_WIDTH -1 :0] atomic_read_data_mask =0;

  /** Helper attribute for randomization calculated during pre_randomize */
  protected bit[`SVT_AXI_MAX_DATA_WIDTH/8 -1 :0] atomic_read_poison_mask =0;

  /** Helper attribute for randomization calculated during pre_randomize */
  protected bit[`SVT_AXI_MAX_DATA_WIDTH -1 :0] atomic_comp_read_data_mask =0;

  /** Helper attribute for randomization calculated during pre_randomize */
  protected int log_base_2_cache_line_size = 0;

  /** internal flag to track if transaction is part of a multi-part dvm sequence */

  bit is_part_of_multipart_dvm_sequence = 0;

  /** The channel (READ/WRITE) on which this transaction will be transmitted */
  xact_type_enum transmitted_channel = WRITE;

  /** The xact_type when port_cfg is_downstream_coherent = 1 */
  xact_type_enum converted_xact_type = WRITE; 
  /** @endcond */
 
  // ****************************************************************************
  // Local variables only for internal VIP usages
  // ****************************************************************************
  bit [(`CEIL(`SVT_AXI_MAX_ID_WIDTH,8))-1:0] axidchk_parity_value = 0;
  bit [(`CEIL(`SVT_AXI_MAX_ADDR_WIDTH,8))-1:0] axaddrchk_parity_value = 0;
  bit axlenchk_parity_value  = 0;
  bit axctlchk0_parity_value = 0;
  bit axctlchk1_parity_value = 0;
  bit axctlchk2_parity_value = 0;
  bit arctlchk3_parity_value = 0;
  bit [(`CEIL((`SVT_AXI_MAX_DATA_WIDTH/8),8))-1:0]       wstrbchk_parity_value;

  // ****************************************************************************
  // Constraints
  // ****************************************************************************

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
neqHt4zg1Wx6PK8KmGjA/kFn51Hh6+a5O05MVdt6uDvk7xWqAo180WH49J3NwfZ9
P6F/koNwgQBm3AO7fAjuKjOzZs5By2tpaphaJ4r1R3ij9betfT/yL/vV9SV9KUkN
Z7ZkIRyvUcSbYqHDjs0DjSsP+eL0SPgmxmU6l/bpvN8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 329       )
TXbUNHeTWIIir6HxugIp661DPVkX3lzaderDgbhQhlmjqQU+klMAW5FCy7X++qPV
yXZIyVcALwrb07FZ+3EoXVWFYxrg3S4PSLsL954dQeiy77h97fbDfeXBVf8fbzdR
P4rJT/oZIfg+trvp812SSTTtM8Sy6YxojBJ6P9JU+u9B5thgWuognhdVqBbXeL4o
DMPGFwWuTJIiEdNfIAb1AcHNH4VtmS7ddAeL+VbvqtICCNf8P+fBew0WxD5d9tDT
DEOhpo1WC1Re3Rjzig0vFOxff3I3Hy1Rj293jygMh54bDaq5891KyGpYi90eLC0H
lQVeC9v4919r/bMi7nQQ6AiREIJS0BftlELKv4WG6t8Qp5lzAc4bkPtGEHnod9co
kvdv3u2SiActj9JooL9Mw59yqASDCSbzva57WSTgVtFtKDJiDrJj7qCZyNP5pMTn
`pragma protect end_protected
  
  /** Re-organised constraint blocks based on interface type. This will make
   * it easy to turn-off the constraints based on interface type. It can
   * result in significant run-time improvement. */

  // QVN Constraints Block. These constraints are valid when QVN mode is
  // enabled. 
  constraint qvn_valid_ranges {
`ifdef SVT_AXI_QVN_ENABLE
    solve xact_type before qvn_vnet_id;
    solve coherent_xact_type before qvn_vnet_id;

`ifndef SVT_AXI_SVC_NO_CFG_IN_XACT
    if(port_cfg.qvn_enable) {
        // -------------------------------------------------------------------------------
        // Each Transaction should pick Virtual Network only from the list of supported VN
        // -------------------------------------------------------------------------------
        qvn_vnet_id inside {[0:`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1]};

        if (xact_type == WRITE || (`SVT_AXI_COHERENT_WRITE) ) {
          foreach(port_cfg.qvn_supported_virtual_network_queue_aw_chnl[ix]) {
            (!port_cfg.qvn_supported_virtual_network_queue_aw_chnl[ix]) -> qvn_vnet_id != ix;
          }
        } else {
          foreach(port_cfg.qvn_supported_virtual_network_queue_ar_chnl[ix]) {
            (!port_cfg.qvn_supported_virtual_network_queue_ar_chnl[ix]) -> qvn_vnet_id != ix;
          }
        }
        // -------------------------------------------------------------------------------
    }
    else {
       qvn_vnet_id == 0;
    }
`endif // SVT_AXI_SVC_NO_CFG_IN_XACT
`endif // SVT_AXI_QVN_ENABLE
  } // qvn_valid_ranges

// These constraints are applicable for Memory tagging feature
 constraint memory_tagging_valid_ranges {
`ifdef SVT_ACE5_ENABLE
 if(port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER){
 if(port_cfg.mte_support_type != svt_axi_port_configuration::NOT_SUPPORTED && port_cfg.use_external_port_monitor ==1){
   if(transmitted_channel == WRITE || transmitted_channel == READ_WRITE) {
     if(port_cfg.mte_support_type == svt_axi_port_configuration::BASIC){
       !tag_op inside {TAG_TRANSFER,TAG_FETCH_MATCH};
       if(xact_type == ATOMIC){
         tag_op == TAG_INVALID;}
    if(xact_type == COHERENT)  {
      if(coherent_xact_type inside {WRITENOSNOOP,WRITEUNIQUE,WRITELINEUNIQUE}){
       tag_op  inside {TAG_INVALID,TAG_UPDATE}; }
      else if (coherent_xact_type inside {CMO,WRITEPTLCMO,WRITEFULLCMO,WRITEUNIQUEPTLSTASH,WRITEUNIQUEFULLSTASH,STASHONCESHARED,STASHONCEUNIQUE,STASHTRANSLATION}){
      tag_op ==TAG_INVALID;}
     }
   if(xact_type == WRITE){
     tag_op  inside {TAG_INVALID,TAG_UPDATE};}
   }
   if(port_cfg.mte_support_type == svt_axi_port_configuration::STANDARD){
     tag_op inside {TAG_INVALID,TAG_UPDATE,TAG_TRANSFER,TAG_FETCH_MATCH};
      if(xact_type == ATOMIC){
         tag_op inside {TAG_INVALID,TAG_FETCH_MATCH};}
      if(xact_type == COHERENT)  {
        if(coherent_xact_type == WRITENOSNOOP){
          tag_op  inside {TAG_INVALID,TAG_UPDATE,TAG_TRANSFER,TAG_FETCH_MATCH};}
        else if(coherent_xact_type inside {WRITEUNIQUE,WRITELINEUNIQUE}) {
          tag_op  inside {TAG_INVALID,TAG_UPDATE};}
        else if (coherent_xact_type inside {WRITEPTLCMO,WRITEFULLCMO}){
          tag_op inside {TAG_INVALID,TAG_TRANSFER,TAG_UPDATE};}
        else if (coherent_xact_type inside{CMO,WRITEUNIQUEPTLSTASH,WRITEUNIQUEFULLSTASH,STASHONCESHARED,STASHONCEUNIQUE,STASHTRANSLATION}){
          tag_op == TAG_INVALID;}
         }
       if(xact_type == WRITE){
         tag_op inside {TAG_INVALID,TAG_UPDATE,TAG_TRANSFER,TAG_FETCH_MATCH};
        }
       }
     }
  if(transmitted_channel == READ) {
    tag_op  inside {TAG_INVALID,TAG_TRANSFER,TAG_FETCH_MATCH};
    if(xact_type == COHERENT)  {
      if(coherent_xact_type == READNOSNOOP){
       tag_op  inside {TAG_INVALID,TAG_TRANSFER,TAG_FETCH_MATCH}; }
      else if (coherent_xact_type == READONCE){
       tag_op  inside {TAG_INVALID,TAG_TRANSFER};}
      else if (coherent_xact_type inside {READONCEMAKEINVALID,READONCECLEANINVALID,CLEANINVALID,MAKEINVALID,CLEANSHARED,CLEANSHAREDPERSIST,DVMMESSAGE,DVMCOMPLETE}){
      tag_op ==TAG_INVALID;}
    }
   if(xact_type == READ){
      tag_op  inside {TAG_INVALID,TAG_TRANSFER,TAG_FETCH_MATCH}; }
  }
  if (tag_op != TAG_INVALID){
  // Transactions must be cacheline sized or smaller
  //For an INCR burst, the last byte in the burst, as determined from the burst length in bytes,
  //(AWSIZE x AWLEN), added to the AWSIZE aligned start address, must be within the same
  //cache line as the first byte in the burst
  //i.e addr_aligned_to_burst_size + bytes_in_transfer < addr_aligned_to_cache_line_size + cache_line_size
      (burst_type == INCR) -> (((addr >> burst_size) << burst_size) + (burst_length << burst_size) <= 
      ((addr >> log_base_2_cache_line_size) << log_base_2_cache_line_size) + port_cfg.cache_line_size);
   // For a WRAP burst, AWSIZE x AWLEN must not exceed the cache line size.
      (burst_type == WRAP) -> ((burst_length << burst_size) <= port_cfg.cache_line_size);

 // For INCR transactions address must be aligned to container size
    if(burst_type == INCR){
     addr == addr >> (burst_length << burst_size) << (burst_length << burst_size);
    }

  // For WRAP transactions address must be aligned to burst_size
    if(burst_type == WRAP){
      addr == addr >> burst_size << burst_size; }

    cache_type[3:2] != 2'b00;
    cache_type[1:0] == 2'b11; 
   }
  if(tag_op == TAG_INVALID){
    foreach(tag[i])
      tag[i] == 0;}

  // Transaction type inside READ,WRITE,COHERENT and ATOMIC  
  xact_type inside {READ,WRITE,COHERENT,ATOMIC};
  if(xact_type == COHERENT){
    coherent_xact_type inside {WRITENOSNOOP,WRITEUNIQUE,WRITELINEUNIQUE,CMO,WRITEUNIQUEPTLSTASH,WRITEUNIQUEFULLSTASH,STASHONCESHARED,STASHONCEUNIQUE,STASHTRANSLATION,WRITEPTLCMO,WRITEFULLCMO,
                                READNOSNOOP,READONCE,READONCEMAKEINVALID,READONCECLEANINVALID,CLEANINVALID,MAKEINVALID,CLEANSHARED,CLEANSHAREDPERSIST,DVMMESSAGE,DVMCOMPLETE};
  }
  }
}
// constraints on response_tag_op only applicable in external port monitor mode
 if(port_cfg.mte_support_type != svt_axi_port_configuration::NOT_SUPPORTED && port_cfg.use_external_port_monitor ==1){
   if(port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE){
     if(port_cfg.use_external_port_monitor == 1){
       if(transmitted_channel == READ){
         if(tag_op == TAG_INVALID){
          response_tag_op inside {TAG_INVALID,TAG_TRANSFER};}
         else if(tag_op == TAG_TRANSFER){
         response_tag_op == TAG_TRANSFER};
        }
       else if(transmitted_channel == READ_WRITE || transmitted_channel == WRITE){
         response_tag_op == TAG_INVALID;
       }
     }
     else {
       response_tag_op == TAG_INVALID;
     }
     if(transmitted_channel == READ_WRITE || transmitted_channel == WRITE){
      tag_match_resp inside{ MATCH_NOT_PERFORMED,NO_MATCH_RESULT,FAIL, PASS};
     }
     else if(transmitted_channel == READ){
      tag_match_resp == MATCH_NOT_PERFORMED;
     }
   }
 }
`endif
 }

// These constraints are applicable for MPAM feature
constraint mpam_valid_ranges {
`ifdef SVT_ACE5_ENABLE
  if (port_cfg.enable_mpam == svt_axi_port_configuration::MPAM_FALSE && port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER && port_cfg.is_active) {
    mpam_partid == 0;
    mpam_perfmongroup == 0;
    mpam_ns == prot_type[1];
  } 
`endif
}

// These constraints are applicable for Write with CMO transactions 
 constraint write_with_cmo_xacts_valid_ranges {
`ifdef SVT_ACE5_ENABLE
  if(xact_type == COHERENT && (coherent_xact_type == WRITEPTLCMO || coherent_xact_type == WRITEFULLCMO)){
    domain_type inside {INNERSHAREABLE,OUTERSHAREABLE,NONSHAREABLE};
    atomic_type == NORMAL;
    cache_type[1] == 1;
  }
 if(port_cfg.axi_interface_type != svt_axi_port_configuration::ACE_LITE){
   !(coherent_xact_type inside {CMO,WRITEPTLCMO,WRITEFULLCMO});
  } 
 if(port_cfg.write_plus_cmo_enable != 1){
    !(coherent_xact_type inside {WRITEPTLCMO,WRITEFULLCMO});
  }
 if(port_cfg.cmo_on_write_enable != 1){
   coherent_xact_type != CMO;
 }
`endif
 }
 //These constraints are valid for atomic transactions .
constraint atomic_xacts_valid_ranges {
`ifdef SVT_ACE5_ENABLE 
   if(!port_cfg.axi_interface_type inside{svt_axi_port_configuration::AXI4,svt_axi_port_configuration::ACE_LITE})  {
      xact_type != ATOMIC;}
//   if(port_cfg.check_type != svt_axi_port_configuration::ODD_PARITY_BYTE_DATA){
//      atomic_read_is_datachk_parity_error == 0;}
   if(xact_type ==ATOMIC){
  //  data size should be equal to burst length
     if(port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
      
      if((barrier_type == NORMAL_ACCESS_RESPECT_BARRIER) || (barrier_type == NORMAL_ACCESS_IGNORE_BARRIER)){ 
          if ((domain_type == NONSHAREABLE) || (domain_type == SYSTEMSHAREABLE)){
             coherent_xact_type  == WRITENOSNOOP;}
          else{
             coherent_xact_type  == WRITEUNIQUE;}
        }
        else{
           coherent_xact_type == WRITEBARRIER;}
       if(burst_length > 1 && ! port_cfg.allow_multibeat_atomic_transactions_to_be_less_than_data_width){
         (1 << burst_size) == port_cfg.data_width/8;
       }
       data.size() == burst_length;
       wstrb.size() == burst_length;
       if (!port_cfg.wysiwyg_enable) {
        foreach (wstrb[index]) {
          wstrb[index] == ((1 << (1 << burst_size)) - 1);
        }
      }
      awakeup_assert_delay ==0;
       if( atomic_xact_op_type inside{ATOMICLOAD_ADD,ATOMICLOAD_CLR,ATOMICLOAD_EOR,ATOMICLOAD_SET,ATOMICLOAD_SMAX,ATOMICLOAD_SMIN,ATOMICLOAD_UMAX,ATOMICLOAD_UMIN}){
          atomic_transaction_type == LOAD;
         }
       if(atomic_xact_op_type inside{ATOMICSTORE_ADD,ATOMICSTORE_CLR,ATOMICSTORE_EOR,ATOMICSTORE_SET,ATOMICSTORE_SMAX,ATOMICSTORE_SMIN,ATOMICSTORE_UMAX,ATOMICSTORE_UMIN}) {
          atomic_transaction_type == STORE;
        }
       if(atomic_xact_op_type == ATOMICSWAP){
          atomic_transaction_type == SWAP;
        }
       if(atomic_xact_op_type == ATOMICCOMPARE){
         atomic_transaction_type == COMPARE;
         burst_size inside{0,1,2,3,4,5};
         {((1 << burst_size)) * burst_length} inside {2,4,8,16,32};
         if(burst_length << burst_size == 2 && addr[0]==1'b0){ 
           burst_type == INCR;}
         else if(burst_length << burst_size == 4 && addr[1:0]==2'b0) {
            burst_type == INCR;}
         else if(burst_length << burst_size == 8 && addr[2:0]==3'b0) {
           burst_type == INCR;}
         else if(burst_length << burst_size == 16 && addr[3:0]==4'b0) {
           burst_type == INCR;}
         else if(burst_length << burst_size == 32 && addr[4:0]==5'b0) {
           burst_type == INCR;}
         else if(burst_length << burst_size == 2 && addr[0] !=1'b0){
           burst_type == WRAP;}
         else if(burst_length << burst_size == 4 && addr[1:0] !=2'b0) {
           burst_type == WRAP;}
         else if(burst_length << burst_size == 8 && addr[2:0] !=3'b0) {
           burst_type == WRAP;}
         else if(burst_length << burst_size == 16 && addr[3:0] !=4'b0) {
           burst_type == WRAP;}
         else if(burst_length << burst_size == 32 && addr[4:0] !=5'b0) {
           burst_type == WRAP;}
          } 
        atomic_transaction_type != NON_ATOMIC;
        if(atomic_transaction_type == COMPARE ){
           atomic_swap_data.size() == burst_length;
           atomic_compare_data.size() == burst_length;
           atomic_compare_wstrb.size() == burst_length;
           atomic_swap_wstrb.size() == burst_length;
           foreach(atomic_swap_data[index]) {
             if(port_cfg.wysiwyg_enable ==1'b1){
                atomic_swap_data[index] == atomic_swap_data[index] & ((1<<(port_cfg.data_width))-1);}
            }
           foreach(atomic_compare_data[index]) {
             if(port_cfg.wysiwyg_enable ==1'b1){
                atomic_compare_data[index] == atomic_compare_data[index] & ((1<<(port_cfg.data_width))-1);}
            }
           if (!port_cfg.wysiwyg_enable) {
             foreach (atomic_swap_data[index]) {
               atomic_swap_data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
             } 
           }
           if (!port_cfg.wysiwyg_enable) {
             foreach (atomic_compare_data[index]) {
               atomic_compare_data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
             } 
           }
        }
        else {
           atomic_swap_data.size() == 0;
           atomic_compare_data.size() == 0;
           atomic_compare_wstrb.size() ==0;
           atomic_swap_wstrb.size() ==0;
         }
         if(atomic_transaction_type ==LOAD){
           atomic_xact_op_type inside{ATOMICLOAD_ADD,ATOMICLOAD_CLR,ATOMICLOAD_EOR,ATOMICLOAD_SET,ATOMICLOAD_SMAX,ATOMICLOAD_SMIN,ATOMICLOAD_UMAX,ATOMICLOAD_UMIN};}
         else if(atomic_transaction_type ==STORE){
           atomic_xact_op_type inside{ATOMICSTORE_ADD,ATOMICSTORE_CLR,ATOMICSTORE_EOR,ATOMICSTORE_SET,ATOMICSTORE_SMAX,ATOMICSTORE_SMIN,ATOMICSTORE_UMAX,ATOMICSTORE_UMIN};}
         else if(atomic_transaction_type ==SWAP){
           atomic_xact_op_type inside{ATOMICSWAP};}
         else if(atomic_transaction_type ==COMPARE){
           atomic_xact_op_type inside{ATOMICCOMPARE};}

//     Address for atomic transactions must be aligned to the data size
         if(atomic_transaction_type !=COMPARE){
           burst_size inside {0,1,2,3};
           {((1 << burst_size)) * burst_length} inside {1,2,4,8};
           burst_type==INCR;
           if (burst_length << burst_size == 2) {
              addr[0] == 1'b0;
            } 
            else if (burst_length << burst_size == 4) {
              addr[1:0] == 2'b0;
            } 
            else if (burst_length << burst_size == 8) {
              addr[2:0] == 3'b0;
            } 
          }
//   For an Atomic compare transactions address must be aligned to half of the burst_size
         else if(atomic_transaction_type == COMPARE){
           burst_size inside {0,1,2,3,4,5};
            if(burst_length << burst_size == 4){
              addr[0] == 1'b0;}
            else if (burst_length << burst_size == 8) {
              addr[1:0] == 2'b0;
            } 
            else if (burst_length << burst_size == 16) {
              addr[2:0] == 3'b0;
            } 
           else if(burst_length << burst_size == 32){
              addr[3:0] == 4'b0;
           }
         }

       if(atomic_transaction_type == COMPARE) {
         atomic_swap_wstrb.size() == burst_length;
         atomic_compare_wstrb.size() == burst_length;
         }
       else {
         atomic_swap_wstrb.size() == 0;
         atomic_compare_wstrb.size() == 0;
       }
     if(atomic_transaction_type != COMPARE){
         burst_type == INCR;
         burst_size inside {0,1,2,3};
        }
       else if(atomic_transaction_type == COMPARE){
         burst_type inside{INCR,WRAP};
         burst_size inside{0,1,2,3,4,5};
        }
         if(xact_type ==ATOMIC){
        wvalid_delay.size() == burst_length;
        rready_delay.size() == burst_length;
         }
    }

  /* 
   * 1) Constraint the atomic_read_data_trace_tag to 1 based on trace_tag value
   */
    if(port_cfg.axi_port_kind == svt_axi_port_configuration:: AXI_SLAVE){
      if(!(atomic_transaction_type inside{LOAD,SWAP,COMPARE})){
         atomic_read_data.size() ==0;
         atomic_read_poison.size() ==0;
         atomic_read_data_user.size() ==0;
        }
       if(atomic_transaction_type inside{LOAD,SWAP} && xact_type == ATOMIC) {
        atomic_read_data.size() == burst_length;
        atomic_read_data_user.size() == burst_length;
        atomic_read_poison.size() == burst_length;

        foreach(atomic_read_data[index]) {
           if(port_cfg.wysiwyg_enable ==1'b1){
              atomic_read_data[index] == atomic_read_data[index] & atomic_read_data_mask;}
          }

        foreach(atomic_read_data_user[index]) {
           if(port_cfg.wysiwyg_enable ==1'b1){
              atomic_read_data_user[index] == atomic_read_data_user[index] & atomic_read_data_mask;}
          }
 
         if(port_cfg.poison_enable ==1){
           if(port_cfg.data_width>64){
             foreach(atomic_read_poison[index]) {
               if(port_cfg.wysiwyg_enable ==1'b1){
                 atomic_read_poison[index] == atomic_read_poison[index] & atomic_read_poison_mask;}
         }}}

         if (!port_cfg.wysiwyg_enable) {
           foreach (atomic_read_data[index]) {
             atomic_read_data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
           } 
         }
         if (!port_cfg.wysiwyg_enable) {
           foreach (atomic_read_data_user[index]) {
             atomic_read_data_user[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
           } 
         }
         if(port_cfg.poison_enable ==1){
           if (!port_cfg.wysiwyg_enable) {
             if(burst_size>3){
               foreach (atomic_read_poison[index]) {
                 atomic_read_poison[index] <= ((1 << ((1 << burst_size) >> 3)) - 1);
               } 
         }}}

      }
      if(atomic_transaction_type == COMPARE && xact_type ==ATOMIC){
        if(burst_length > 1){
          atomic_read_data.size() == burst_length/2;
          atomic_read_data_user.size() == burst_length/2;
          atomic_read_poison.size() == burst_length/2;
        }
        else {
          atomic_read_data.size() == 1;
          atomic_read_data_user.size() == 1;
          atomic_read_poison.size() == 1;
        }

        foreach(atomic_read_data[index]) {
           if(port_cfg.wysiwyg_enable ==1'b1){
              atomic_read_data[index] == atomic_read_data[index] & atomic_comp_read_data_mask;}
          }

        foreach(atomic_read_data_user[index]) {
           if(port_cfg.wysiwyg_enable ==1'b1){
              atomic_read_data_user[index] == atomic_read_data_user[index] & atomic_comp_read_data_mask;}
          }
 
         if(port_cfg.poison_enable ==1){
           if(port_cfg.data_width>64){
             foreach(atomic_read_poison[index]) {
               if(port_cfg.wysiwyg_enable ==1'b1){
                 atomic_read_poison[index] == atomic_read_poison[index] & atomic_read_poison_mask;}
         }}}

         if (!port_cfg.wysiwyg_enable) {
           foreach (atomic_read_data[index]) {
             atomic_read_data[index] <= ((1 << (((1 << burst_size)>>1) << 3)) - 1);
           } 
         }
         if (!port_cfg.wysiwyg_enable) {
           foreach (atomic_read_data_user[index]) {
             atomic_read_data_user[index] <= ((1 << (((1 << burst_size)>>1) << 3)) - 1);
           } 
         }
         if(port_cfg.poison_enable ==1){
           if (!port_cfg.wysiwyg_enable) {
             if(burst_size>3){
               foreach (atomic_read_poison[index]) {
                 atomic_read_poison[index] <= ((1 << ((1 << burst_size) >> 3)) - 1);
               } 
         }}}
        }

      if(trace_tag ==1 && atomic_transaction_type inside{LOAD,SWAP,COMPARE} && xact_type == ATOMIC){
        atomic_read_data_trace_tag == 1;
       }
      if(atomic_transaction_type inside{LOAD,SWAP,COMPARE} && xact_type == ATOMIC){
        rvalid_delay.size() == burst_length;
        foreach (rvalid_delay[idx])
          rvalid_delay[idx] inside {[0:`SVT_AXI_MAX_RVALID_DELAY]};
            }
       wready_delay.size()==burst_length;
    }

  }
    if(xact_type == ATOMIC && atomic_transaction_type inside{LOAD,SWAP} ){
       rresp.size()== burst_length ;
     }
     if(xact_type == ATOMIC && atomic_transaction_type inside{COMPARE} ){
       if(burst_length > 1){
         rresp.size()== burst_length/2 ;}
       else {
         rresp.size() ==1;}
     }
    
/*     if(xact_type == ATOMIC) {
       if(burst_length > 1){
          1 << burst_size == data_width_in_bytes;}
      }*/
  if(xact_type != ATOMIC)
    {
       atomic_read_data.size() ==0;
       atomic_read_poison.size() ==0;
       atomic_read_data_user.size() ==0;
       atomic_swap_data.size() ==0;
       atomic_compare_data.size() ==0;
       atomic_swap_wstrb.size()==0;
       atomic_compare_wstrb.size()==0;
       atomic_transaction_type == NON_ATOMIC;
    }
   if(xact_type ==ATOMIC){
     atomic_type == NORMAL;
     random_interleave_array.size() == burst_length;
     random_interleave_array[0] == 1;
    }
     xact_type != READ_WRITE;
     converted_xact_type != READ_WRITE;
     transmitted_channel != ATOMIC;
`endif
}

  // ACE/ACE-Lite Constraints Block. These constraints are valid if the
  // interface type is set to ACE or ACE-Lite.

  constraint ace_valid_ranges {

    foreach(data[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        data[index] == data[index] & ((1<<(port_cfg.data_width))-1);}
    }

`ifdef SVT_ACE5_ENABLE
   if(port_cfg.atomic_transactions_enable ==1'b1 && atomic_transaction_type inside{LOAD,SWAP,COMPARE} && xact_type == ATOMIC) {
      foreach(atomic_read_data[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        atomic_read_data[index] == atomic_read_data[index] & ((1<<(port_cfg.data_width))-1);}
    }

      foreach(atomic_read_data_user[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        atomic_read_data_user[index] == atomic_read_data_user[index] & ((1<<(port_cfg.data_width))-1);}
    }

     foreach(atomic_swap_data[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        atomic_swap_data[index] == atomic_swap_data[index] & ((1<<((port_cfg.data_width)))-1);}
    }
      foreach(atomic_compare_data[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        atomic_compare_data[index] == atomic_compare_data[index] & ((1<<(port_cfg.data_width))-1);}
    }

   if(port_cfg.poison_enable ==1 && port_cfg.wysiwyg_enable ==1){
       foreach(atomic_read_poison[index]) {
         if(port_cfg.data_width%64 == 0) {
           atomic_read_poison[index] == atomic_read_poison[index] & ((1<<(port_cfg.data_width/64))-1);}
         else {
           atomic_read_poison[index] == atomic_read_poison[index] & (((1<<(port_cfg.data_width/64)+1))-1);}
   }}
  }
`endif

 if(port_cfg.poison_enable ==1){
      foreach(poison[index]) {
        if(port_cfg.wysiwyg_enable ==1'b1){
         if(port_cfg.data_width%64 == 0) {
            poison[index] == poison[index] & ((1<<(port_cfg.data_width/64))-1);}
         else {
            poison[index] == poison[index] & (((1<<(port_cfg.data_width/64)+1))-1);}
    }}
   }
   
`ifdef SVT_ACE5_ENABLE
// This transaction types are not yet supported  
   !(coherent_xact_type inside {STASHTRANSLATION});
`endif 

`ifdef SVT_AXI_SVC_USE_MODEL
      if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration :: AXI_ACE || `SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  ACE_LITE) {

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
`endif
     if (`SVT_AXI_COHERENT_READ_1_BEAT) { 
       random_interleave_array.size() == 1;
       random_interleave_array[0] == 1;
     }
   }
      if(port_cfg.ace_version == svt_axi_port_configuration::ACE_VERSION_1_0 && xact_type == COHERENT) {
        !(coherent_xact_type inside{CLEANSHAREDPERSIST,READONCECLEANINVALID,READONCEMAKEINVALID});}

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`endif
     if (`SVT_AXI_COHERENT_READ_1_BEAT) { 
       random_interleave_array.size() == 1;
       random_interleave_array[0] == 1;
     }
`ifdef INCA
     if ((slave_xact_type == COHERENT) && (slave_xact_type != DATA_STREAM )) {
        if( 
            (slave_coherent_xact_type == CLEANUNIQUE) || 
            (slave_coherent_xact_type == MAKEUNIQUE) || 
            (slave_coherent_xact_type == CLEANSHARED) ||
            (slave_coherent_xact_type == CLEANSHAREDPERSIST) ||
            (slave_coherent_xact_type == CLEANINVALID) || 
            (slave_coherent_xact_type == MAKEINVALID) 
          ) {
          wready_delay.size() == 1;
          rvalid_delay.size() == 1;
        }
        else {
          wready_delay.size() == burst_length;
          rvalid_delay.size() == burst_length;
        }
     }
`else  
     if ((xact_type == COHERENT) && 
         (xact_type != DATA_STREAM)) {
       if( 
           (coherent_xact_type == CLEANUNIQUE) || 
           (coherent_xact_type == MAKEUNIQUE) || 
           (coherent_xact_type == CLEANSHARED) || 
           (coherent_xact_type == CLEANSHAREDPERSIST) ||
           (coherent_xact_type == CLEANINVALID) || 
           (coherent_xact_type == MAKEINVALID) 
         ) {
         wready_delay.size() == 1;
         rvalid_delay.size() == 1;
       } else {
         wready_delay.size() == burst_length;
         rvalid_delay.size() == burst_length;
       }
     }  
`endif // `ifdef INCA 
   } // if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE)
   } //       if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  ACE || `SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  ACE_LITE)
`endif //SVT_AXI_SVC_USE_MODEL
 } // ace_valid_ranges

  // AXI4 STREAM Constraints Block. These constraints are valid if the
  // interface type is set to AXI4_STREAM.
  constraint axi4_stream_valid_ranges {
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`endif   
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
`else
      if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
`endif
        random_interleave_array.size() == stream_burst_length;
        foreach (random_interleave_array[index]) {
          random_interleave_array[index] inside {[1 : stream_burst_length]};
        }   
      } // if (port_cfg.axi_interface_type != svt_axi_port_configuration::AXI4_STREAM)
   } // if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE)
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
     if (axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
     if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
`endif
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tid_enable) {
`else
       if (!port_cfg.tid_enable) {
`endif
         tid == 0;
       }
       else {
         tid inside {[0 : ((1 << port_cfg.tid_width) -1)]};
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tdest_enable) {
`else
       if (!port_cfg.tdest_enable) {
`endif
         tdest == 0;
       }
       else {
         tdest inside {[0 : ((1 << port_cfg.tdest_width) -1)]};
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tdata_enable) {
`else
       if (!port_cfg.tdata_enable) {
`endif
         foreach (tdata[index])
           tdata[index] == 0;
       }
       else {
         foreach (tdata[index]) {
             tdata[index] inside {[0 : ((1 << port_cfg.tdata_width) -1)]};
          }
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tstrb_enable) {
`else
       if (!port_cfg.tstrb_enable) {
`endif
         foreach(tstrb[index])
           tstrb[index] == 0;
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tuser_enable) {
`else
       if (!port_cfg.tuser_enable) {
`endif
         foreach(tuser[index])
           tuser[index] == 0;
       }
       else {
         foreach (tuser[index]) {
            tuser[index] inside {[0 : ((1 << port_cfg.tuser_width) -1)]};
          }
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tkeep_enable) {
`else
       if (!port_cfg.tkeep_enable) {
`endif
         foreach(tkeep[index])
           tkeep[index] == 0;
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tlast_enable) {
`else
       if (!port_cfg.tlast_enable) {
`endif
         stream_burst_length == 1;
       }
     } //AXI4_STREAM
   } //AXI_MASTER    
  } // axi4_stream_valid_ranges  


  // AXI3/AXI4/AXI4 Lite Constraints Block. These constraints are valid if the
  // interface type is set to either AXI3/AXI4/AXI4_Lite. Since these are
  // basic AXI constraints they even hold true in case the interface_type is
  // set to ACE/ACE_Lite.

  constraint axi3_4_valid_ranges {
    /*solve burst_length before random_interleave_array;
    solve stream_burst_length before random_interleave_array;
    solve burst_length before addr;
    solve burst_length before wstrb;

    solve burst_size before wstrb;
    solve burst_length before rresp;
    solve burst_length before coh_rresp;
    solve burst_length before rvalid_delay;
    solve burst_length before wready_delay;
    solve xact_type before rvalid_delay;
    solve xact_type before wready_delay;
    solve coherent_xact_type before rvalid_delay;
    solve coherent_xact_type before wready_delay;
    solve xact_type before rresp;
    solve coherent_xact_type before rresp;
    solve xact_type before coh_rresp;
    solve coherent_xact_type before coh_rresp;
    */

  foreach(data[index]) {
     if(port_cfg.wysiwyg_enable ==1'b1){
       data[index] == data[index] & ((1<<(port_cfg.data_width))-1);}
   }

   if(port_cfg.poison_enable ==1){
      foreach(poison[index]) {
        if(port_cfg.wysiwyg_enable ==1'b1){
           if(port_cfg.data_width%64 == 0) {
              poison[index] == poison[index] & ((1<<(port_cfg.data_width/64))-1);}
           else {
              poison[index] == poison[index] & (((1<<(port_cfg.data_width/64)+1))-1);}
        }
      }
    }

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
    burst_length <= `SVT_AXI3_MAX_BURST_LENGTH;
`else
    if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI3)
      burst_length <= `SVT_AXI3_MAX_BURST_LENGTH;
    else
      burst_length <= `SVT_AXI4_MAX_BURST_LENGTH;
`endif //SVT_AXI_SVC_NO_CFG_IN_XACT
      if(port_cfg.ace_version == svt_axi_port_configuration::ACE_VERSION_1_0 && xact_type == COHERENT) {
        !(coherent_xact_type inside{CLEANSHAREDPERSIST,READONCECLEANINVALID,READONCEMAKEINVALID});}

`ifdef SVT_AXI_SVC_USE_MODEL

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
`endif
      // Constraining the Delay sizes
      if (`SVT_AXI_COHERENT_READ_1_BEAT) {
        wvalid_delay.size() == 1;
        rready_delay.size() == 1;
        data.size() == 1;
        if(port_cfg.poison_enable ==1){
        poison.size() == 1;}
      } else if (xact_type != DATA_STREAM) {
        wvalid_delay.size() == burst_length;
        rready_delay.size() == burst_length;
        data.size() == burst_length;
       if(port_cfg.poison_enable ==1){
       poison.size() == burst_length;
      }}

`ifndef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (port_cfg.toggle_ready_signals_during_idle_period) {
        if ((xact_type == READ) || `SVT_AXI_COHERENT_READ) {
          idle_rready_delay.size() inside {[0:`SVT_AXI_MAX_IDLE_RREADY_DELAY_ARR_SIZE]};
          idle_bready_delay.size() == 0;
        } else {
          idle_bready_delay.size() inside {[0:`SVT_AXI_MAX_IDLE_BREADY_DELAY_ARR_SIZE]};
          idle_rready_delay.size() == 0; 
        }
      } else {
        idle_rready_delay.size() == 0;
        idle_bready_delay.size() == 0;
      }

     if (!port_cfg.wysiwyg_enable) {
        foreach (data[index]) {
          data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
        } 
      }
     foreach(data[index]) {
       if(port_cfg.wysiwyg_enable ==1'b1){
         data[index] == data[index] & ((1<<(port_cfg.data_width))-1);}
      }

    if(port_cfg.poison_enable ==1 && !port_cfg.wysiwyg_enable){
        foreach (poison[index]) {
          if((1 << burst_size)%8 !=0){
            poison[index] <= ((1 << (((1 << burst_size) >> 3)+1)) - 1);}
          else {
             poison[index] <= ((1 << ((1 << burst_size) >> 3)) - 1);}
        } 
      }

   if(port_cfg.poison_enable ==1  && port_cfg.wysiwyg_enable ==1){
      foreach(poison[index]) {
           if(port_cfg.data_width%64 == 0) {
              poison[index] == poison[index] & ((1<<(port_cfg.data_width/64))-1);}
           else {
              poison[index] == poison[index] & (((1<<(port_cfg.data_width/64)+1))-1);}
        }
    }
`endif

      /*
       * 1) Constrain the array size to 0 if xact_type is not READ
       * 2) Constrain the array size to burst length if xact_type is READ
       */    
      if ((xact_type == READ) || `SVT_AXI_COHERENT_READ) {
        if (`SVT_AXI_COHERENT_READ_1_BEAT) 
          rresp.size() == 1;
        else
          rresp.size() == burst_length; 
      }
`ifdef SVT_ACE5_ENABLE
     else if(xact_type == ATOMIC && atomic_transaction_type inside{LOAD,SWAP} ){
       rresp.size()== burst_length ;
      }
     if(xact_type == ATOMIC && atomic_transaction_type inside{COMPARE}){
       if(burst_length > 1){
         rresp.size()== burst_length/2 ;}
       else {
         rresp.size() ==1;}
     }
`endif      
      else {
        rresp.size() == 0;
      }

      /* 
       *  Constraints for wstrb 
       *  1) Constraint the length of the wstrb from 1 to burst_length for write
         transactions
       *  2) Constraining wstrb to enable all the valid bytelanes depending on transfer
      */
      if (xact_type == WRITE || (`SVT_AXI_COHERENT_WRITE) 
`ifdef SVT_ACE5_ENABLE
|| xact_type ==ATOMIC
`endif    
       ) {
        wstrb.size() == burst_length;
      }
      else
        wstrb.size() == 0;
      /*if (!port_cfg.wysiwyg_enable) {
        foreach (wstrb[index]) {
          wstrb[index] inside {[0: ((1 << (1 << burst_size)) - 1)]};
        }
      }
      */
`ifdef SVT_ACE5_ENABLE
       if(xact_type == ATOMIC){
          data.size() == burst_length;
       }
`endif

      if (`SVT_AXI_COHERENT_READ_1_BEAT) {
        data_user.size() == 1;
      } else if (xact_type == DATA_STREAM) {
        data_user.size() == 0;
      } else {
        data_user.size() == burst_length;
      }
`ifdef SVT_MULTI_SIM_ENUM_RANDOMIZES_TO_INVALID_VALUE
`ifdef SVT_ACE5_ENABLE 
    xact_type inside {READ,WRITE,IDLE,COHERENT,ATOMIC};
`else
    xact_type inside {READ,WRITE,IDLE,COHERENT,DATA_STREAM};
`endif
`endif

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) {
`else
      if (port_cfg.axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) {
`endif
        xact_type != DATA_STREAM;

`ifdef SVT_MULTI_SIM_ENUM_RANDOMIZES_TO_INVALID_VALUE
        atomic_type inside {NORMAL,EXCLUSIVE,LOCKED};
        burst_type inside {FIXED,INCR,WRAP};
`endif

`ifndef SVT_AXI_SVC_NO_CFG_IN_XACT
        /* 
         * The atomic type is not exclusive when exclusive_access_enable is
         * disabled
         */  
        if (port_cfg.exclusive_access_enable == 0) {
          atomic_type != EXCLUSIVE;    
        }
        if (port_cfg.locked_access_enable == 0) {
          atomic_type != LOCKED;    
        }
`endif
        
        
        /** Address is within limits specified by addr_width. */
        addr <= max_possible_addr;
        addr_user <= max_possible_user_addr;

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
        id <= ((1 << `SVT_AXI_MAX_ID_WIDTH) - 1);
`else
        if (port_cfg.use_separate_rd_wr_chan_id_width == 0 
`ifdef SVT_ACE5_ENABLE
          || xact_type == ATOMIC
`endif
         ) 
          id <= ((1 << port_cfg.id_width) - 1);
        else if ((xact_type == WRITE) || `SVT_AXI_COHERENT_WRITE)
          id <= ((1 << port_cfg.write_chan_id_width) - 1);
        else 
          id <= ((1 << port_cfg.read_chan_id_width) - 1);
`endif

        /*
         *  When the burst type is not Fixed, it must be ensured that burst does not
         *  exceed 4k range
         */
   
        if(burst_type != FIXED) {
          addr_range == (burst_length * (1 << burst_size));
          `ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
          addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << burst_size);
          `else
          addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << burst_size);
          `endif  
          if (burst_type == WRAP) {
            // Make sure that the max address does not cross addr_width.
            // Need to calculate this from wrap boundary (lowest address)
            // Note that the max byte address is:
            // (burst_length-1)*bytes_in_each_transfer + (bytes_in_each_transfer-1)
            if (burst_length == 2)
`ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
              burst_addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << (burst_size+1));
`else
              burst_addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << (burst_size+1));
`endif
            else if (burst_length == 4)
`ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
              burst_addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << (burst_size+2));
`else
              burst_addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << (burst_size+2));
`endif
            else if (burst_length == 8)
`ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
              burst_addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << (burst_size+3));
`else
              burst_addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << (burst_size+3));
`endif
            else if (burst_length == 16)
`ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
              burst_addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << (burst_size+4));
`else
              burst_addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << (burst_size+4));
`endif

            addr == (addr & addr_mask);
            (addr & burst_addr_mask) + addr_range - 1 <= max_possible_addr; 
            (addr[11:0] & burst_addr_mask) <= (`SVT_AXI_TRANSACTION_4K_ADDR_RANGE - addr_range);
          } else {
            // INCR
            (addr[11:0] & addr_mask) <= (`SVT_AXI_TRANSACTION_4K_ADDR_RANGE - addr_range);
            // Make sure that the max address does not cross addr_width.
            // Use aligned address
            ((addr >> burst_size) << burst_size) + addr_range - 1 <= max_possible_addr;
          }
        } 


        
        // Resetting all the bits greater than data width to 0

        /*foreach (wstrb[index]) {
          if (index < burst_length) {
            wstrb[index] == wstrb[index] & ((1 << port_cfg.data_width/8)-1);
          } 
        }
        */


        addr_valid_delay inside {[0:`SVT_AXI_MAX_ADDR_VALID_DELAY]};
        

        foreach (wvalid_delay[index]) {
          wvalid_delay[index] inside {[0:`SVT_AXI_MAX_WVALID_DELAY]};
        }
        foreach (rready_delay[index]) {
          rready_delay[index] inside {[0:`SVT_AXI_MAX_RREADY_DELAY]};
        }
        foreach (idle_rready_delay[index]) {
          idle_rready_delay[index] inside {[0:`SVT_AXI_MAX_IDLE_RREADY_DELAY]};
        }

        /*if (reference_event_for_rready_delay == MANUAL_RREADY) {
          foreach (rready_delay[index]) {
            (index == 0) -> rready_delay[index] inside {[-`SVT_AXI_MAX_RREADY_DELAY : `SVT_AXI_MAX_RREADY_DELAY]};
            (index > 0)  -> rready_delay[index] inside {[0:`SVT_AXI_MAX_RREADY_DELAY]};
          }
        } else {
          foreach (rready_delay[index]) {
            rready_delay[index] inside {[0:`SVT_AXI_MAX_RREADY_DELAY]};
          }
        }
        */

        bready_delay inside {[`SVT_AXI_MIN_WRITE_RESP_DELAY:`SVT_AXI_MAX_WRITE_RESP_DELAY]};
        foreach (idle_bready_delay[index]) {
          idle_bready_delay[index] inside {[0:`SVT_AXI_MAX_IDLE_BREADY_DELAY]};
        }


        // Data Before Addr Constraints
        if(data_before_addr) {
          reference_event_for_first_wvalid_delay == PREV_WRITE_DATA_HANDSHAKE;
          reference_event_for_addr_valid_delay inside {FIRST_WVALID_DATA_BEFORE_ADDR,FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR};
        }

        if (!(`SVT_AXI_COHERENT_READ_1_BEAT)) {

          random_interleave_array.size() == burst_length;
          foreach (random_interleave_array[index]) {
            random_interleave_array[index] inside {[1 : burst_length]};
          }
        }
      } // if (port_cfg.axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) 

      // For EXCLUSIVE access, the address must be aligned to 
      // the total number of bytes transferred
      if (atomic_type == EXCLUSIVE) {
        (burst_length << burst_size) inside {1,2,4,8,16,32,64,128};

        if (burst_length << burst_size == 2) {
          addr[0] == 1'b0;
        } 
        else if (burst_length << burst_size == 4) {
          addr[1:0] == 2'b0;
        } 
        else if (burst_length << burst_size == 8) {
          addr[2:0] == 3'b0;
        } 
        else if (burst_length << burst_size == 16) {
          addr[3:0] == 4'b0;
        } 
        else if (burst_length << burst_size == 32) {
          addr[4:0] == 5'b0;
        } 
        else if (burst_length << burst_size == 64) {
          addr[5:0] == 6'b0;
        } 
        else if (burst_length << burst_size == 128) {
          addr[6:0] == 7'b0;
        } 
      }

      /* 
       * AXI3 :
       * 1) Burst Size must not exceed the data width
       * 2) Burst Length for WRAP is inside 2,4,8,16
       * 3) Total No. of bytes to be transferred in an exclusive access burst must be a
       *   power of 2.  Max is 128  - Section 6.2.4
       * 4) Burst Length For Idle transactions must be from 1 to Max Idles
       * 5)
      */   

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (axi_interface_type == svt_axi_port_configuration :: AXI3) {
`else
      if (port_cfg.axi_interface_type == svt_axi_port_configuration :: AXI3) {
`endif
 
        xact_type != COHERENT;
        burst_size <= log_base_2_data_width_in_bytes;

        if (xact_type == IDLE) {
          burst_length inside {[1:`SVT_AXI_MAX_TRANSACTION_IDLE_CYCLES]}; 
        } else {
          if (burst_type == WRAP) {
`ifdef SVT_ACE5_ENABLE
           if(xact_type == ATOMIC && atomic_transaction_type == COMPARE){
              burst_length inside {1,2,4,8,16,32};}
           else {
              burst_length inside {2,4,8,16};}
`else
             burst_length inside {2,4,8,16};
`endif
          } else {
            burst_length inside {[1:`SVT_AXI3_MAX_BURST_LENGTH]};
          }
        }

        // WA(bit 3) bit must not be high if C bit(bit 1) is low
        (cache_type[1] == 0) -> (cache_type[3] == 0);
        // Reserved values:
        cache_type != 4'b0100;
        cache_type != 4'b0101;
        cache_type != 4'b1000;
        cache_type != 4'b1001;
        cache_type != 4'b1100;
        cache_type != 4'b1101;
      }

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      foreach(data_user[i])
       data_user[i] <= ((1 << `SVT_AXI_MAX_DATA_USER_WIDTH) - 1);
`else
      foreach(data_user[i])
       data_user[i] <= ((1 << port_cfg.data_user_width) - 1);
`endif
   }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`endif
`ifndef SVT_AXI_SVC_NO_CFG_IN_XACT

`ifdef SVT_ACE5_ENABLE    
   if(port_cfg.atomic_transactions_enable ==1){
      if(!(atomic_transaction_type inside{LOAD,SWAP,COMPARE})){
         atomic_read_data.size() ==0;
         atomic_read_poison.size() ==0;
         atomic_read_data_user.size() ==0;
        }
      if(atomic_transaction_type inside{LOAD,SWAP} && xact_type == ATOMIC) {
         atomic_read_data.size() <= burst_length;
         atomic_read_poison.size() <= burst_length;
         atomic_read_data_user.size() <= burst_length;
       }
       if(atomic_transaction_type inside{COMPARE} && xact_type == ATOMIC) {
         if(burst_length > 1){
           atomic_read_data.size() == burst_length/2;
           atomic_read_poison.size() == burst_length/2;
           atomic_read_data_user.size() == burst_length/2;
         }
         else {
           atomic_read_data.size() == 1;
           atomic_read_poison.size() == 1;
           atomic_read_data_user.size() == 1;
         }
        }
      }
   else {
     atomic_read_data.size() ==0;
     atomic_read_data_user.size() ==0;
     atomic_read_poison.size() ==0;
//     atomic_resultant_data.size() ==0;
//     atomic_swap_data.size() ==0;
//     atomic_compare_data.size() ==0;
    }
`endif
      if (port_cfg.enable_delayed_response_port) {
        // Transaction supplied through delayed response port.
        // data.size() can be <= burst_length since data is provided
        // through multiple transactions.
        if (is_delayed_response_xact) {
          if (`SVT_AXI_COHERENT_READ_1_BEAT) {
           if(port_cfg.poison_enable ==1){
            poison.size() == 1;}
            data.size() == 1;
            rresp.size() == 1;
          } else if ((xact_type == READ) || (`SVT_AXI_COHERENT_READ)) {
          if(port_cfg.poison_enable ==1){
            poison.size() <= burst_length;}
            data.size() <= burst_length;
            rresp.size() <= burst_length;
            data.size() == rresp.size();
          if(port_cfg.poison_enable ==1){
           poison.size() == rresp.size();}
          }
`ifdef SVT_ACE5_ENABLE
      else if(atomic_transaction_type inside{LOAD,SWAP} && xact_type == ATOMIC ) {
        rresp.size() == burst_length;
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() <= burst_length;
          poison.size() <= burst_length;}
        atomic_read_data.size() <= burst_length;
        atomic_read_data.size() == rresp.size();
        atomic_read_data_user.size() <= burst_length;
        atomic_read_data_user.size() == rresp.size();
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() == rresp.size();}        
        data.size() <= burst_length;
        rresp.size() <= burst_length;  }
      else if(atomic_transaction_type inside{COMPARE} && xact_type == ATOMIC ) {
        if(burst_length > 1){
        rresp.size() == burst_length/2;
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() <= burst_length/2;
          poison.size() <= burst_length;}
        atomic_read_data.size() <= burst_length/2;
        atomic_read_data_user.size() <= burst_length/2;
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() == rresp.size();}        
        data.size() <= burst_length;
        }
        else {
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() <= burst_length;
          poison.size() <= burst_length;}
        atomic_read_data.size() <= burst_length;
        atomic_read_data.size() == rresp.size();
        atomic_read_data_user.size() <= burst_length;
        atomic_read_data_user.size() == rresp.size();
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() == rresp.size();}        
        data.size() <= burst_length;
        rresp.size() <= burst_length;}
       }
`endif  
       else {
            rresp.size() == 0;
          }  
        // Transaction supplied through seq_item_port but when
        // configured with enable_delayed_response_port. This corresponds
        // to the transaction handle that is returned in 0-time to the driver.
        } else {
          if ((xact_type == READ) || (`SVT_AXI_COHERENT_READ)) {
             data.size() == 0;
           if(port_cfg.poison_enable ==1){
             poison.size() == 0;}
             rresp.size() == 0;
          // WRITES
          }
       else {
            rresp.size() == 0;
          }
        }
      } else 
`endif
      {
        if (xact_type == DATA_STREAM) {
          data.size() == 0;
           if(port_cfg.poison_enable ==1){
             poison.size() == 0;}
        } else if (`SVT_AXI_COHERENT_READ_1_BEAT) {
          data.size() == 1;
         if(port_cfg.poison_enable ==1){
           poison.size() == 1;}
          rresp.size() == 1;
          data_user.size() == 1;
        } else if ((xact_type == READ) || `SVT_AXI_COHERENT_READ) {
          data.size() == burst_length;
          if(port_cfg.poison_enable ==1){
            poison.size() == burst_length;}
          rresp.size() == burst_length;
          data_user.size() == burst_length;
        // WRITES. rresp_size should be 0.
        }
`ifdef SVT_ACE5_ENABLE
      else if(atomic_transaction_type inside{LOAD,SWAP} && xact_type == ATOMIC) {
        rresp.size() == burst_length;
        atomic_read_data.size() == burst_length;
        atomic_read_poison.size() == burst_length;
        atomic_read_data_user.size() == burst_length;
       }
       else if(atomic_transaction_type inside{COMPARE} && xact_type == ATOMIC) {
        if(burst_length >1){
        rresp.size() == burst_length/2;
        atomic_read_data.size() == burst_length/2;
        atomic_read_poison.size() == burst_length/2;
        atomic_read_data_user.size() == burst_length/2;
        }
       else {
        rresp.size() == burst_length;
        atomic_read_data.size() == burst_length;
        atomic_read_poison.size() == burst_length;
        atomic_read_data_user.size() == burst_length;
       }
       }
       else if(xact_type == ATOMIC && !(atomic_transaction_type inside{LOAD,SWAP,COMPARE})){
         rresp.size() ==0;
         atomic_read_data.size()==0;
         atomic_read_data_user.size()==0;
         atomic_read_poison.size()==0;
      }
`endif  
        else {
          data_user.size() == burst_length;
          data.size() == burst_length;
          rresp.size() == 0;
        }
      }

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) {
`else
      if (port_cfg.axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) {
`endif
        if (!(`SVT_AXI_COHERENT_READ_1_BEAT)) { 
          random_interleave_array.size() == burst_length;
          foreach (random_interleave_array[index]) {
            random_interleave_array[index] inside {[1 : burst_length]};
          }
        }
      } 

      addr_ready_delay inside {[0:`SVT_AXI_MAX_ADDR_DELAY]};

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      resp_user <= ((1 << `SVT_AXI_MAX_BRESP_USER_WIDTH) - 1);
`else
      resp_user <= ((1 << port_cfg.resp_user_width) - 1);
`endif


    // wready_delay[0] can take positive and negative values.
`ifdef INCA
      if ((slave_xact_type != COHERENT) && (slave_xact_type != DATA_STREAM )) {
        wready_delay.size() == burst_length;
        rvalid_delay.size() == burst_length;
      }
`else
      if ((xact_type != COHERENT) && (xact_type != DATA_STREAM )) {
        wready_delay.size() == burst_length;
        rvalid_delay.size() == burst_length;
      }
`endif
      if (port_cfg.toggle_ready_signals_during_idle_period)
        idle_addr_ready_delay.size() inside {[0:`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY_ARR_SIZE]}; 
      else
        idle_addr_ready_delay.size() == 0;
      if (xact_type == WRITE 
`ifdef SVT_ACE5_ENABLE
         || xact_type == ATOMIC
`endif           
         || xact_type == COHERENT && 
          (coherent_xact_type == WRITENOSNOOP ||
           coherent_xact_type == WRITELINEUNIQUE ||
           coherent_xact_type == WRITEUNIQUE ||
`ifdef SVT_ACE5_ENABLE
             coherent_xact_type == WRITEUNIQUEPTLSTASH ||
             coherent_xact_type == WRITEUNIQUEFULLSTASH ||
`endif
           coherent_xact_type == WRITEBACK   ||
           coherent_xact_type == WRITECLEAN  ||
           coherent_xact_type == WRITEEVICT
          )
         ) {
        if (port_cfg.toggle_ready_signals_during_idle_period)
          idle_wready_delay.size() inside {[0:`SVT_AXI_MAX_IDLE_WREADY_DELAY_ARR_SIZE]}; 
        else
          idle_wready_delay.size() == 0;
      } else {
        idle_wready_delay.size() == 0;
      }
      if (xact_type != DATA_STREAM) {
       if(!port_cfg.axi_slv_channel_buffers_enable)
        foreach (rvalid_delay[idx])
          rvalid_delay[idx] inside {[0:`SVT_AXI_MAX_RVALID_DELAY]};

        if (reference_event_for_wready_delay == MANUAL_WREADY) {
          foreach (wready_delay[idx]) {
            (idx == 0) -> wready_delay[idx] inside {[-`SVT_AXI_MAX_WREADY_DELAY:`SVT_AXI_MAX_WREADY_DELAY]};
            (idx > 0) -> wready_delay[idx] inside {[0:`SVT_AXI_MAX_WREADY_DELAY]};
          }
        } else {
          foreach (wready_delay[idx])
            wready_delay[idx] inside {[0:`SVT_AXI_MAX_WREADY_DELAY]};
          foreach (idle_wready_delay[idx])
            idle_wready_delay[idx] inside {[0:`SVT_AXI_MAX_IDLE_WREADY_DELAY]};
          foreach (idle_addr_ready_delay[idx])
            idle_addr_ready_delay[idx] inside {[0:`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY]};
        }
       if(!port_cfg.axi_slv_channel_buffers_enable)
        bvalid_delay inside {[`SVT_AXI_MIN_WRITE_RESP_DELAY:`SVT_AXI_MAX_WRITE_RESP_DELAY]};
        if (xact_type == WRITE  
`ifdef SVT_ACE5_ENABLE
         || xact_type == ATOMIC
`endif      
         ||   xact_type == COHERENT && 
             (coherent_xact_type == WRITENOSNOOP ||
             coherent_xact_type == WRITELINEUNIQUE ||
             coherent_xact_type == WRITEUNIQUE ||
`ifdef SVT_ACE5_ENABLE
             coherent_xact_type == WRITEUNIQUEPTLSTASH ||
             coherent_xact_type == WRITEUNIQUEFULLSTASH ||
`endif
             coherent_xact_type == WRITEBACK   ||
             coherent_xact_type == WRITECLEAN  ||
             coherent_xact_type == WRITEEVICT  ||
             coherent_xact_type == EVICT
            )
           ) {
        // The reordering priority of write responses be within
        // 1 to port_cfg.write_resp_reordering_depth.
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
        reordering_priority inside {[1:`SVT_AXI_MAX_WRITE_RESP_REORDERING_DEPTH]};
`else
        reordering_priority inside {[1:port_cfg.write_resp_reordering_depth]};
`endif
        }
        else { //if (xact_type == READ) 
        // The reordering priority of read transactions should be within
        // 1 to port_cfg.read_data_reordering_depth.
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
        reordering_priority inside {[1:`SVT_AXI_MAX_READ_DATA_REORDERING_DEPTH]};
`else
        reordering_priority inside {[1:port_cfg.read_data_reordering_depth]};
`endif
        }

        // An EXOKAY response makes sense only for an EXLUSIVE type
        // atomic access.
        if (atomic_type != EXCLUSIVE) { 
          foreach (rresp[idx])
            (rresp[idx] != EXOKAY); 
          bresp != EXOKAY; 
        }

        if (
            (xact_type == COHERENT) && 
            ( 
              (coherent_xact_type == CLEANUNIQUE) || 
              (coherent_xact_type == MAKEUNIQUE) || 
              (coherent_xact_type == CLEANSHARED) || 
              (coherent_xact_type == CLEANSHAREDPERSIST) || 
              (coherent_xact_type == CLEANINVALID) || 
              (coherent_xact_type == MAKEINVALID) 
            ) 
           ) {
          foreach (random_interleave_array[index]) {
            random_interleave_array[index] inside {[0 : 1]};
          }
        } else {
          foreach (random_interleave_array[index]) {
            random_interleave_array[index] inside {[0 : burst_length]};
          }
        }
      }
    } // if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) 
`endif //SVT_AXI_SVC_USE_MODEL
  } // axi3_4_valid_ranges 

 
  constraint disable_constraint_first_wvalid_reference_event {
    reference_event_for_first_wvalid_delay dist { WRITE_ADDR_VALID:=50000, WRITE_ADDR_HANDSHAKE:=1, PREV_WRITE_DATA_HANDSHAKE:=50000 };
  }

 constraint valid_poison {
    if(port_cfg.poison_enable == 0){
       poison.size()==0;
    }
   }


`ifdef INCA 
   constraint validpoison {
     if(port_cfg.poison_enable==1 && port_cfg.ace_version==svt_axi_port_configuration::ACE_VERSION_2_0){
        poison.size()==1;
     }
     else {
       poison.size()==0;
     }
    }
`endif

`ifdef SVT_ACE5_ENABLE
    constraint valid_archunken{
	        if(port_cfg.rdata_chunking_enable == 1 && xact_type == READ){
		        if(burst_size >= BURST_SIZE_128BIT){
			        archunken inside {0,1};
                  }
		        else {
			        archunken == 0;
                }
            }
	        else {	
		        archunken == 0;
            }
        }

    constraint reasonable_ranges_while_chunking {
      solve chunk_length before rchunkstrb;
      solve chunk_length before rchunknum;
        if(archunken){
            rchunkstrb.size() == chunk_length;
            rchunknum.size() == chunk_length;
        }
        else {
            rchunkstrb.size() == 0;
            rchunknum.size() == 0;
        }
    }

    constraint reasonable_chunk_len{
      solve burst_length before chunk_length;
      solve burst_size before chunk_length;
      if(archunken){
        if(burst_size < BURST_SIZE_128BIT){
          chunk_length == 0;
        }
        else {
          chunk_length inside {[burst_length:(burst_length<<(burst_size - 4))]};
        }
      }
      else {
        chunk_length == 0;
      }
    }
`endif
 /*Reasonable constraint on reference_event_for_addr_delay in data_before_addr scenarios
 reference_event_for_addr_delay must not be set to FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR as this may cause 
 potential deadlock scenarios in ACE SLAVE DUT where slave DUT waits for awvalid signal
 before driving wready signal.
 */
 constraint reasonable_reference_event_for_addr_delay {
   if(data_before_addr){
   reference_event_for_addr_valid_delay inside {FIRST_WVALID_DATA_BEFORE_ADDR};}
 }
    
`ifdef SVT_AXI_SVC_USE_MODEL
  // **************************************************************************
  //       Reasonable  Constraints
  // **************************************************************************

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
EWTJGaG/60wA1yGypQs5YBNDlO5p/I/wcRzBmF8k8ImZX2x/ity/Rq73XMoUbEPE
TKgn/foj0gl/k6e0zWYi4THVibwwyO6KNWTNvpeFURr/pVhdCFgam0Q86PwbT6Yk
iE9gF2+0X00QS8xs6hIqg7fOGUctodMRPG1NhOSrfpQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 602       )
Mas5LorPfMNRzoKsnqX/Pt/9FHlqgrdXfmpb80E5hRywV9M2YicsYueaMYyfXr7e
+36RpFStnwzh2+7R9grlg470jeOXTQmwhf601FIqQywQodqAqiuDhcL0MVza0xmj
dkNo2IaCHrOZUGp6JmW0lzhikfulNlGpIwYG1eurKLlI8qX5c9b2zgvp7ofUZlML
m0Cc3dOl3pENRfBeq26rLt+4wl7lN5VVpp/5sVq6cleOt18o5fXAZcBE91hyOXQz
ORyjYj10PNZe/PCXZ5nL9i0c7TJJdce70zrQdi9f9b1kBW0URNaG+eodDsT7PoLB
15955qQ7AZQK1IJR3F1H0/e9W4omcpRCcr7z9Yl8ofekopEyzukuYcwpt408j4Oz
`pragma protect end_protected
  constraint reasonable_burst_length {
    if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI3) {  
      burst_length dist {
        1 := ZERO_BURST_wt,
        [2: (`SVT_AXI3_MAX_BURST_LENGTH >> 2)] :/ SHORT_BURST_wt,
        [(`SVT_AXI3_MAX_BURST_LENGTH >> 2)+1:`SVT_AXI3_MAX_BURST_LENGTH] :/ LONG_BURST_wt
      };
    }
    if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI4 ||
        `SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  ACE_LITE) {  
      burst_length dist {
        1 := ZERO_BURST_wt,
        [2: (`SVT_AXI4_MAX_BURST_LENGTH >> 2)] :/ SHORT_BURST_wt,
        [(`SVT_AXI4_MAX_BURST_LENGTH >> 2)+1:`SVT_AXI4_MAX_BURST_LENGTH] :/ LONG_BURST_wt
      };
    }
    if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI_ACE) {
      burst_length dist {
        1 := ZERO_BURST_wt,
        [2:4] :/ SHORT_BURST_wt,
        [5:16] :/ LONG_BURST_wt
      };
    }
  }

  /*
    Reasonable constraint for cache type.
    For exclusive accesses transactions , transactions must not be cached
  */
  constraint reasonable_cache_type
  {
    solve atomic_type before cache_type;
      if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI3) {   
        if (atomic_type == EXCLUSIVE) {
          cache_type inside {`SVT_AXI_3_NON_CACHEABLE_NON_BUFFERABLE,
                             `SVT_AXI_3_BUFFERABLE_OR_MODIFIABLE_ONLY,
                             `SVT_AXI_3_CACHEABLE_BUT_NO_ALLOC,
                             `SVT_AXI_3_CACHEABLE_BUFFERABLE_BUT_NO_ALLOC};
        }
      } 
      if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI4) {
        if (atomic_type == EXCLUSIVE) {
          cache_type inside {`SVT_AXI_4_ARCACHE_DEVICE_NON_BUFFERABLE,
                             `SVT_AXI_4_ARCACHE_DEVICE_BUFFERABLE,
                             `SVT_AXI_4_ARCACHE_NORMAL_NON_CACHABLE_NON_BUFFERABLE,
                             `SVT_AXI_4_ARCACHE_NORMAL_NON_CACHABLE_BUFFERABLE};
        }
      } 
  }

  /* 
    Reasonable constraint for interleave_pattern
    1) Set the interleave pattern to RANDOM BLOCK for the user to set interleave
    patterns
  */  

  constraint reasonable_interleave_pattern {
    interleave_pattern == RANDOM_BLOCK;
  }

  /* 
    Reasonable constraint for equal block length
    1) Constrain the equal block length to range of 1 to burst_length/2
  */
  
  constraint reasonable_equal_block_length {
    solve interleave_pattern before equal_block_length;
    solve burst_length before equal_block_length;
    if (interleave_pattern ==  EQUAL_BLOCK) {
      if (burst_length > 1) {
        equal_block_length  inside {[1 : (burst_length >> 1)]};
      }
      else {
        equal_block_length == 1;
      }
    }
  }

  constraint reasonable_addr_valid_delay {
   addr_valid_delay dist {
     0 := ZERO_DELAY_wt, 
     [1:(`SVT_AXI_MAX_ADDR_VALID_DELAY >> 2)] :/ SHORT_DELAY_wt,
     [((`SVT_AXI_MAX_ADDR_VALID_DELAY >> 2)+1):`SVT_AXI_MAX_ADDR_VALID_DELAY] :/ LONG_DELAY_wt
   };
  }


  constraint reasonable_wakeup_assert_deassert_delay {
    awakeup_assert_delay >= `SVT_AXI_MIN_AWAKEUP_ASSERT_DELAY;
    awakeup_assert_delay <  `SVT_AXI_MAX_AWAKEUP_ASSERT_DELAY;
    awakeup_deassert_delay >= `SVT_AXI_MIN_AWAKEUP_DEASSERT_DELAY;
    awakeup_deassert_delay <  `SVT_AXI_MAX_AWAKEUP_DEASSERT_DELAY;
  }

  constraint reasonable_rready_delay {
    /*foreach (rready_delay[idx]) {
      if (reference_event_for_rready_delay == MANUAL_RREADY && idx == 0) {
        rready_delay[idx] dist {
         0 := ZERO_DELAY_wt,
         [-(`SVT_AXI_MAX_RREADY_DELAY >> 2):-1] :/ SHORT_DELAY_wt >> 1,
         [1:(`SVT_AXI_MAX_RREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
         [-`SVT_AXI_MAX_RREADY_DELAY: -((`SVT_AXI_MAX_RREADY_DELAY >> 2)+1)] :/ LONG_DELAY_wt >> 1,
         [((`SVT_AXI_MAX_RREADY_DELAY >> 2)+1):`SVT_AXI_MAX_RREADY_DELAY] :/ LONG_DELAY_wt >> 1
        };
      } else {
          rready_delay[idx] dist {
          0 := ZERO_DELAY_wt,
          [1:(`SVT_AXI_MAX_RREADY_DELAY >> 2)] := SHORT_DELAY_wt >> 1,
          [((`SVT_AXI_MAX_RREADY_DELAY >> 2)+1):`SVT_AXI_MAX_RREADY_DELAY] := LONG_DELAY_wt >> 1
          };
      }
    }
    */
    foreach (rready_delay[idx]) {
      rready_delay[idx] dist {
            0 := ZERO_DELAY_wt,
            [1:(`SVT_AXI_MAX_RREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
            [((`SVT_AXI_MAX_RREADY_DELAY >> 2)+1):`SVT_AXI_MAX_RREADY_DELAY] :/ LONG_DELAY_wt
      };
    }
  }

  constraint reasonable_idle_rready_delay {
    foreach (idle_rready_delay[idx]) {
      idle_rready_delay[idx] dist {
            0 := ZERO_DELAY_wt,
            [1:(`SVT_AXI_MAX_IDLE_RREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
            [((`SVT_AXI_MAX_IDLE_RREADY_DELAY >> 2)+1):`SVT_AXI_MAX_IDLE_RREADY_DELAY] :/ LONG_DELAY_wt
      };
    }
  }

  
  // Enforces a distribution based on the weights.
  constraint reasonable_wvalid_delay {
    foreach (wvalid_delay[idx]) {
      wvalid_delay[idx] dist {
       0 := ZERO_DELAY_wt, 
       [1:(`SVT_AXI_MAX_WVALID_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_WVALID_DELAY >> 2)+1):`SVT_AXI_MAX_WVALID_DELAY] :/ LONG_DELAY_wt
      };
    }
  }


  // Enforces a distribution based on the weights.
  constraint reasonable_bready_delay {
    bready_delay dist {
       `SVT_AXI_MIN_WRITE_RESP_DELAY := ZERO_DELAY_wt, 
       [(`SVT_AXI_MIN_WRITE_RESP_DELAY + 1):(`SVT_AXI_MAX_WRITE_RESP_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_WRITE_RESP_DELAY >> 2)+1):`SVT_AXI_MAX_WRITE_RESP_DELAY] :/ LONG_DELAY_wt
    };
  }

  constraint reasonable_idle_bready_delay {
    foreach (idle_bready_delay[i]) 
      idle_bready_delay[i] dist {
       0 := ZERO_DELAY_wt, 
       [1:(`SVT_AXI_MAX_IDLE_BREADY_DELAY>> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_IDLE_BREADY_DELAY>> 2)+1):`SVT_AXI_MAX_IDLE_BREADY_DELAY] :/ LONG_DELAY_wt
    };
  }


  constraint reasonable_tready_delay {
    if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
      tready_delay.size() == `SVT_AXI_MAX_STREAM_BURST_LENGTH;
      foreach (tready_delay[idx]) {
        tready_delay[idx] dist {
         0 := ZERO_DELAY_wt, 
         [1:(`SVT_AXI_MAX_TREADY_DELAY >> 2)] :/ SHORT_DELAY_wt,
         [((`SVT_AXI_MAX_TREADY_DELAY >> 2)+1):`SVT_AXI_MAX_TREADY_DELAY] :/ LONG_DELAY_wt
       };
      }
    } else {
      tready_delay.size() == 0;
    }
  }

  /** 
   * This constraint insures that unimplemented features are avoided during randomization.
   */
  constraint exclude_master_unimplemented_features
  {
    xact_type != IDLE;
    interleave_pattern != EQUAL_BLOCK;
    start_new_interleave == 0;
    reference_event_for_rready_delay != MANUAL_RREADY;
  }

  //--------------------------------------------------------------------------------------
  /**************************** SLAVE CONSTRAINTS ******************************** */
  constraint reasonable_data {
    if (`SVT_AXI_INTERFACE_TYPE != svt_axi_port_configuration::AXI4_STREAM) {
      if (
           (xact_type == READ) || 
           (
             (xact_type == COHERENT) &&
             (
               coherent_xact_type == READNOSNOOP                     ||
               coherent_xact_type == READONCE                        ||
               coherent_xact_type == READONCECLEANINVALID                        ||
               coherent_xact_type == READONCEMAKEINVALID                        ||
               coherent_xact_type == READSHARED                      ||
               coherent_xact_type == READCLEAN                       ||
               coherent_xact_type == READNOTSHAREDDIRTY              ||
               coherent_xact_type == READUNIQUE          
             )
           )
         ) {
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
         data.size() == burst_length;
         if(port_cfg.poison_enable ==1){
            poison.size() == burst_length;}
`else
       if (!port_cfg.enable_delayed_response_port) {
           if(port_cfg.poison_enable ==1){
             poison.size() == burst_length;}
           data.size() == burst_length;
       }
`endif
       data_user.size() == burst_length;
        foreach (data[index]) {
             data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
        }
      }
      // No data associated with these transactions 
      if(`SVT_AXI_COHERENT_READ_1_BEAT) {
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
        if(port_cfg.poison_enable ==1){
           poison.size() == 1;}
        data.size() == 1;
`else
       if (!port_cfg.enable_delayed_response_port) {
          if(port_cfg.poison_enable ==1){
             poison.size() == 1;}
          data.size() == 1;
       }
`endif
       data_user.size() == 1;
        foreach (data[index]) {
             data[index] <= 0;
        }
      if(port_cfg.poison_enable ==1){
            foreach (poison[index]) {
             poison[index] <= 0;}
          }
      }
    }
  }

  // Enforces a distribution based on the weights.
  constraint reasonable_wready_delay {
    foreach (wready_delay[idx]) {
      // MANUAL_READY not supported.
      /*if (reference_event_for_wready_delay == MANUAL_WREADY && idx == 0) {
        wready_delay[idx] dist {
         0 := ZERO_DELAY_wt,
         [-(`SVT_AXI_MAX_WREADY_DELAY >> 2):-1] :/ SHORT_DELAY_wt >> 1,
         [1:(`SVT_AXI_MAX_WREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
         [-`SVT_AXI_MAX_WREADY_DELAY: -((`SVT_AXI_MAX_WREADY_DELAY >> 2)+1)] :/ LONG_DELAY_wt >> 1,
         [((`SVT_AXI_MAX_WREADY_DELAY >> 2)+1):`SVT_AXI_MAX_WREADY_DELAY] :/ LONG_DELAY_wt >> 1
        };
      } else {*/ 
        wready_delay[idx] dist {
          0 := ZERO_DELAY_wt,
          [1:(`SVT_AXI_MAX_WREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
          [((`SVT_AXI_MAX_WREADY_DELAY >> 2)+1):`SVT_AXI_MAX_WREADY_DELAY] :/ LONG_DELAY_wt
          };
        //}
      }
    }

  // Enforces a distribution based on the weights.
  constraint reasonable_idle_wready_delay {
    foreach (idle_wready_delay[idx]) {
        idle_wready_delay[idx] dist {
          0 := ZERO_DELAY_wt,
          [1:(`SVT_AXI_MAX_IDLE_WREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
          [((`SVT_AXI_MAX_IDLE_WREADY_DELAY >> 2)+1):`SVT_AXI_MAX_IDLE_WREADY_DELAY] :/ LONG_DELAY_wt
          };
    }
  }
 

  // Enforces a distribution based on the weights.
  constraint reasonable_rvalid_delay {
    foreach (rvalid_delay[idx]) {
      rvalid_delay[idx] dist {
       0 := ZERO_DELAY_wt, 
       [1:(`SVT_AXI_MAX_RVALID_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_RVALID_DELAY >> 2)+1):`SVT_AXI_MAX_RVALID_DELAY] :/ LONG_DELAY_wt
      };
    }
  }

  // Enforces a distribution based on the weights.
  constraint reasonable_addr_ready_delay {
    addr_ready_delay dist {
       0 := ZERO_DELAY_wt, 
       [1:(`SVT_AXI_MAX_ADDR_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_ADDR_DELAY >> 2)+1):`SVT_AXI_MAX_ADDR_DELAY] :/ LONG_DELAY_wt
    };
  }

  // Enforces a distribution based on the weights.
  constraint reasonable_idle_addr_ready_delay {
    foreach (idle_addr_ready_delay[idx]) {
      idle_addr_ready_delay[idx] dist {
         0 := ZERO_DELAY_wt, 
         [1:(`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY >> 2)] :/ SHORT_DELAY_wt,
         [((`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY >> 2)+1):`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY] :/ LONG_DELAY_wt
      };
    }
  }

  // Enforces a distribution based on the weights.
  constraint reasonable_bvalid_delay {
    bvalid_delay dist {
       `SVT_AXI_MIN_WRITE_RESP_DELAY := ZERO_DELAY_wt, 
       [(`SVT_AXI_MIN_WRITE_RESP_DELAY + 1):(`SVT_AXI_MAX_WRITE_RESP_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_WRITE_RESP_DELAY >> 2)+1):`SVT_AXI_MAX_WRITE_RESP_DELAY] :/ LONG_DELAY_wt
    };
  }

  /**
   * Reasonable constraint for random_interleave_array
   * Constraint the random interleave array from 1 to burstlength
   * If the  array values exceed the burst length, those values will be ignored
   */

   constraint reasonable_random_interleave_array {
     if (`SVT_AXI_INTERFACE_TYPE != svt_axi_port_configuration::AXI4_STREAM) {
       if(`SVT_AXI_COHERENT_READ_1_BEAT) 
         random_interleave_array.size() == 1;
       else
         random_interleave_array.size() == burst_length;

       foreach (random_interleave_array[index]) {
         random_interleave_array[index] inside {[1 : burst_length]};
       }
     } else {
       random_interleave_array.size() == stream_burst_length;
     }
   }

    constraint exclude_slave_unimplemented_features
    {
      interleave_pattern != EQUAL_BLOCK;
      start_new_interleave == 0;
      reference_event_for_wready_delay != MANUAL_WREADY;
    }

`endif

`ifdef SVT_AXI_TRANSACTION_ENABLE_TEST_CONSTRAINTS
  /**
   * External constraint definitions which can be used for test level constraint addition.
   * By default, "test_constraintsX" constraints are not enabled in svt_axi_transaction. A
   * test can enable them by defining the following macro during the compile:
   *   SVT_AXI_TRANSACTION_ENABLE_TEST_CONSTRAINTS
   */
  constraint test_constraints1;
  constraint test_constraints2;
  constraint test_constraints3;
`endif

//reasonable  soft constraint for cust_xact_flow == 0. To support default behavior of cust_xact_flow disabled and overridden by user to enable it automatically whenever inline randomization constraint is added
constraint reasonable_cust_xact_flow {
  soft cust_xact_flow == 0;
} 

`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_transaction",svt_axi_port_configuration port_cfg_handle = null);
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_transaction",svt_axi_port_configuration port_cfg_handle = null);
`else
`svt_vmm_data_new(`SVT_TRANSACTION_TYPE)
  extern function new (vmm_log log = null, svt_axi_port_configuration port_cfg_handle = null);
`endif

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following
   * 1) Tests the validity of the configuration
   * 2) calculate the log_2 of master configs data_width   
   */
  extern function void pre_randomize ();

  //----------------------------------------------------------------------------
  /**
   *   post_randomize does the following
   *   1) Aligns the address to no of Bytes for Exclusive Accesses
   */
  extern function void post_randomize ();

  /** returns 1 if status of all relevant phases of current transaction are assigned as ABORTED */
  extern virtual function bit is_aborted(int mode = 0);

  /** returns 1 if current transaction is configured as secure access */
  extern virtual function bit is_secure(bit allow_secure = 1);

  /** Returns 1 if current transaction is of device_type */
  extern virtual function bit is_device_type();

  /** Returns 1 if current transaction is DVM transaction */
  extern virtual function bit is_dvm_xact();

  /** Returns 1 if current transaction is cacheable transaction */
  extern virtual function bit is_cacheable_xact();

  /** Returns 1 if current transaction is allocate transaction */
  extern virtual function bit is_allocate_xact();

  /** Determines if this transaction is a CMO transaction */
  extern function bit is_cmo_xact();


//  /** Returns 1 if current transaction is of device_type or DVM transaction 
//   * Additinally this function will fire an error if device type or DVM transactions 
//   * are issued from not allowed ports 
//   */
//  extern virtual function bit skip_port_interleaving();

  /** waits for transaction to end */
  extern virtual task wait_for_transaction_end();


 /** waits for slave transaction to update the memory*/
  extern virtual task wait_for_write_transaction_to_update_memory();

  /** returns 1 if transaction status shows ended otherwise 0 */
  extern virtual function bit is_transaction_ended();

  /** waits for addr phase to end */
  extern virtual task wait_for_addr_phase_ended ();
  
  /** waits for data phase to end */
  extern virtual task wait_for_data_phase_ended();
  
  /** waits for write resp phase to end */
  extern virtual task wait_for_write_resp_phase_ended();

  /** mark end of transaction */
  extern virtual function void set_end_of_transaction(bit aborted=0);
  

   /**
  * Returns 1 if the specified error_kind is there in transaction, else returns 0 
  */
  extern virtual function bit has_axi_exception(int error_kind); 
  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************

  `svt_data_member_begin(svt_axi_transaction)
    `svt_field_object(port_cfg,`SVT_ALL_ON|`SVT_NOCOMPARE|`SVT_NOPACK| `SVT_REFERENCE, `SVT_HOW_REF)
    `ifndef INCA
    `svt_field_object      (exception_list,                             `SVT_ALL_ON|`SVT_DEEP|`SVT_NOCOMPARE|`SVT_UVM_NOPACK,  `SVT_HOW_DEEP)
    `endif
    `svt_field_object(associated_barrier_xact,`SVT_ALL_ON|`SVT_NOCOMPARE|`SVT_NOPACK|`SVT_REFERENCE, `SVT_HOW_REF)
`ifdef SVT_UVM_TECHNOLOGY
    `svt_field_object(causal_gp_xact,`SVT_ALL_ON|`SVT_NOCOMPARE|`SVT_NOPACK|`SVT_REFERENCE, `SVT_HOW_REF)
`endif

  // ****************************************************************************

  `svt_data_member_end(svt_axi_transaction)


  // ****************************************************************************
  // Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * Method to turn reasonable constraints on/off as a block.
   */
  extern virtual function int reasonable_constraint_mode (bit on_off);

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object used for logging.
   */
  extern function string get_mcd_class_name ();

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Extend the copy method to copy the transaction class fields.
   * 
   * @param to Destination class for the copy operation
   */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);

 `else
  //---------------------------------------------------------------------------
  /**
   * Extend the copy method to take care of the transaction fields and cleanup the exception xact pointers.
   *
   * @param rhs Source object to be copied.
   */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);
`endif
 //----------------------------------------------------------------------------
  /**
   * Extend the svt_post_do_all_do_copy method to cleanup the exception xact pointers.
   * 
   * @param to Destination class for the copy operation
   */
  extern virtual function void svt_post_do_all_do_copy(`SVT_DATA_BASE_TYPE to);
 //----------------------------------------------------------------------------
  /**
   * Calculates whether the transaction is partial or full cacheline access.
   * returns 1, if transaction is full cacheline access. returns 0, if it is a 
   * partial cacheline access.
   * 
   * @param cacheline_size indicates the value of the master cache line size
   */
  extern virtual function bit is_full_cacheline(int cacheline_size);

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   * @param comparer TBD
   */
  extern virtual function bit do_compare(uvm_object rhs, uvm_comparer comparer);
`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   * @param comparer TBD
   */
  extern virtual function bit do_compare(ovm_object rhs, ovm_comparer comparer);
`else
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare (vmm_data to, output string diff, input int kind = -1);

  //----------------------------------------------------------------------------
  /**                         
   * Returns the size (in bytes) required by the byte_pack operation.
   *
   * @param kind This int indicates the type of byte_size being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in a size calculation based on the
   * non-static fields. All other kind values result in a return value of 0.
   */
  extern virtual function int unsigned byte_size (int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Packs the object into the bytes buffer, beginning at offset, based on the
   * requested byte_pack kind.
   *
   * @param bytes Buffer that will contain the packed bytes at the end of the operation.
   * @param offset Offset into bytes where the packing is to begin.
   * @param kind This int indicates the type of byte_pack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being packed and the return of an integer indicating the number of
   * packed bytes. All other kind values result in no change to the buffer contents, and a
   * return value of 0.
   */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Unpacks the object from the bytes buffer, beginning at offset, based on
   * the requested byte_unpack kind.
   *
   * @param bytes Buffer containing the bytes to be unpacked.
   * @param offset Offset into bytes where the unpacking is to begin.
   * @param len Number of bytes to be unpacked.
   * @param kind This int indicates the type of byte_unpack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being unpacked and the return of an integer indicating the number of
   * unpacked bytes. All other kind values result in no change to the exception contents,
   * and a return value of 0.
   */
  extern virtual function int unsigned do_byte_unpack (const ref logic [7:0]
  bytes[], input int unsigned offset = 0, input int len = -1, input int kind = -1);

`endif

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>read</i> access to public data members of this class.
   */
  extern virtual function bit get_prop_val (string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>write</i> access to public data members of this class.
   */
  extern virtual function bit set_prop_val (string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
   * This method allocates a pattern containing svt_pattern_data instances for
   * all of the primitive data fields in the object. The svt_pattern_data::name
   * is set to the corresponding field name, the svt_pattern_data::value is set
   * to 0.
   *
   * @return An svt_pattern instance containing entries for all of the data fields.
   */
  extern virtual function svt_pattern do_allocate_pattern ();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB.  The pattern is customized to contain only the fields necessary for
   * the application and tranaction type.
   * 
   * Note:
   * As a performance enhancement, property values in the pattern are pre-populated when
   * the pattern is created.  This allows the FSDB writer infrastructure to skip the
   * get_prop_val_via_pattern step.
   *
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern allocate_xml_pattern();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB when a full tranaction is to be recorded.  Note that not all
   * properties are written.  Instead, only properties needed for debug are added.
   * 
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern populate_full_xml_pattern();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB when the PA channel is RADDR, RDATA, WADDR, WDATA, or WRESP.
   * 
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern populate_filtered_xml_pattern();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB when the PA channel is "STREAM DATA".
   * 
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern populate_stream_xml_pattern();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB when the pa_format_type is set to FSDB_PERF_ANALYSIS.
   * 
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern populate_perf_analysis_xml_pattern();

  // ----------------------------------------------------------------------------
  /**
   * This method returns PA object which contains the PA header information for XML or FSDB.
   *
   * @param uid Optional string indicating the unique identification value for object. If not 
   * provided uses the 'get_uid()' method  to retrieve the value. 
   * @param typ Optional string indicating the 'type' of the object. If not provided
   * uses the type name for the class.
   * @param parent_uid Optional string indicating the UID of the object's parent. If not provided
   * the method assumes there is no parent.
   * @param channel Optional string indicating an object channel. If not provided
   * the method assumes there is no channel.
   *
   * @return The requested object block description.
   */
   extern virtual function svt_pa_object_data get_pa_obj_data(string uid = "", string typ = "", string parent_uid = "", string channel = "" );

//-----------------------------------------------------------------------------------
/**
  * This method is used to set object_type for bus_activity when
  * bus_activity is getting started on the bus .
  * This method is used by pa writer class in generating XML/FSDB 
  */
  extern function void  set_pa_data(string typ = "" ,string channel  ="");
 
//-----------------------------------------------------------------------------------
  /**
  * This method is used to  delate  object_type for bus_activity when bus _activity 
  * ends on the bus .
  * This methid is used by pa writer class  in generating XML/FSDB 
  */
  extern function void clear_pa_data();
  
//------------------------------------------------------------------------------------
  /** This method is used in setting the unique identification id for the
  * objects of bus activity
  * This method returns  a  string which holds uid of bus activity object
  * This is used by pa writer class in generating XML/FSDB
  */
  extern virtual function string get_uid();

//------------------------------------------------------------------------------------
  /** Sets the configuration property */ 
  extern function void set_cfg(svt_axi_port_configuration cfg);

  /** Gets the current byte lane based on the current data beat, address
    * and burst size
    */ 
  extern function int get_curr_byte_lane(int log_base_2_data_width_in_bytes = -1, int beat_num = -1);

`ifdef SVT_ACE5_ENABLE  
  /** Gets the current byte lane based on the current data beat, address
    * and burst size
    */ 
  extern function int get_curr_byte_lane_atomic_write_data(int log_base_2_data_width_in_bytes = -1, int beat_num = -1);

  /** Gets the current byte lane based on the current data beat, address
    * and burst size
    */ 
  extern function int get_curr_byte_lane_atomic_read_data(int log_base_2_data_width_in_bytes = -1, int beat_num = -1);
`endif
  /** 
    * Populates the partial data and byteen provided into data and byteen
    * that is used to write into a full cacheline
    */
  extern function void populate_partial_data_and_byteen (
                                                         input bit[7:0] data[],
                                                         input bit byteen[],
                                                         output bit[7:0] cache_data[],
                                                         output bit cache_byteen[]
      );

  /** Returns the address and lanes corresponding to the beat number */
  extern function void get_beat_addr_and_lane_for_data_user(input int beat_num, 
                                              output [`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                                              output int lower_byte_lane,
                                              output int upper_byte_lane,
                                              input  bit use_tagged_addr=0);
 /** Returns the address and lanes corresponding to the beat number */
  extern function void get_beat_addr_and_lane(input int beat_num, 
                                              output [`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                                              output int lower_byte_lane,
                                              output int upper_byte_lane,
                                              input  bit use_tagged_addr=0);
`ifdef SVT_ACE5_ENABLE
 /** Returns the address and lanes corresponding to the beat number for atomic compare read data*/
  extern function void get_beat_addr_and_lane_atomic_read_data(input int beat_num, 
                                              output [`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                                              output int lower_byte_lane,
                                              output int upper_byte_lane,
                                              input  bit use_tagged_addr=0);
 /** Returns the address and lanes corresponding to the beat number for atomic compare write data*/
  extern function void get_beat_addr_and_lane_atomic_write_data(input int beat_num, 
                                              output [`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                                              output int lower_byte_lane,
                                              output int upper_byte_lane,
                                              input  bit use_tagged_addr=0);
`endif

  /** Gets the beat number corresponding to an address */
  extern function int get_beat_num_of_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr, 
                                                          bit use_tagged_addr = 0
                                          );

  /**
   * Returns a string (with no line feeds) that reports the essential contents
   * of the packet generally necessary to uniquely identify that packet.
   *
   * @param prefix (Optional: default = "") The string given in this argument
   * becomes the first item listed in the value returned. It is intended to be
   * used to identify the transactor (or other source) that requested this string.
   * This argument should be limited to 8 characters or less (to accommodate the
   * fixed column widths in the returned string). If more than 8 characters are
   * supplied, only the first 8 characters are used.
   * @param hdr_only (Optional: default = 0) If this argument is supplied, and
   * is '1', the function returns a 3-line table header string, which indicates
   * which packet data appears in the subsequent columns. If this argument is
   * '1', the <b>prefix</b> argument becomes the column label for the first header
   * column (still subject to the 8 character limit).
   */
`ifdef SVT_UVM_ENABLE_FGP
  (* uvm_fgp_lock = "psdisplay_short" *)
`endif
  extern virtual function string psdisplay_short( string prefix = "", bit hdr_only = 0);

  /** 
    * Limits the data to what can be transmitted if the address is
    * unaligned. If the address is unaligned, we need to take care 
    * that data[0] and wstrb[0] are consistent with what can actually 
    * be driven on the bus. 
    * For example, for a 64 bit bus, if the address is 0x7,
    * data can be sent only on 1 byte for the first beat.
    * For a FIXED burst the address is same for all beats, so this
    * operation needs to be done for all beats. For other bursts, only
    * the first address can be unaligned, other beats are aligned
    * addresses
    * @param data_only(Optional: default = 0) If this bit is set the 
    * operation is done only for data. 
    * @param beat_num(Optional: default = -1) Applicable for a FIXED burst.
    * When set to -1, masking is done for all beats, otherwise it is 
    * done only for the selected beat. 
    */
  extern function void mask_data_for_unaligned_addr(bit data_only = 0,int beat_num = -1);
  
  /**
    * Ensures that valid x,z,0,1 all four state datas are calculated with
    * respect to data_mask values. 
    * This function is called under SVT_MEM_LOGIC_DATA macro define only,
    * to make sure while masking valid x and z state data also considered
    * towards masked data.
    */ 
  extern function logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] mask_data_for_x_z_values (logic [`SVT_AXI_MAX_DATA_WIDTH -1:0] data, bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] data_mask);
  
  /**
    * Ensures that only valid lanes have wstrb asserted. In wysisyg format
    * the constraints leave data[] and wstrb[] open. This function is called in
    * post_randomize to make sure that wstrb is asserted only for valid lanes
    */ 
  extern function void get_wstrb_for_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] wstrb[]);

`ifdef SVT_ACE5_ENABLE
    /**
    * Ensures that only valid lanes have tag_update asserted. In wysisyg format
    * the constraints leave tag[] and tag_update[] open. This function is called in
    * post_randomize to make sure that tag_update is asserted only for valid lanes
    */ 
  extern function void get_tag_update_for_wysiwyg_format(ref bit[`SVT_AXI_MAX_TAGUPDATE_WIDTH-1:0] tag_update[]);

  /**
    * Returns the tag_update in the tag_update_to_pack[] field as a byte stream based on
    * the burst_type. 
    * In the case of WRAP bursts the tag_update is returned such that packed_tag_update[0] 
    * corresponds to the tag_update for the wrap boundary. 
    * In the case of INCR bursts, the wstrb as passed in tag_update_to_pack[] is directly
    * packed to packed_tag_update[]. 
    * @param tag_update_to_pack tag_update to be packed
    * @param packed_tag_update[] Output byte stream with packed tag_update
    */
  extern function void pack_tag_update_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_TAGUPDATE_WIDTH-1:0] tag_update_to_pack[],
                                          output bit packed_tag_update[]
                                        ); 

  /**
    * Returns the tag in the tag_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that either tag[] or cache_write_tag[]
    * fields of this class have been passed as arguments to tag_to_pack[] field.
    * In the case of WRAP bursts the tag is returned such that packed_tag[0] 
    * corresponds to the tag for the wrap boundary. 
    * In the case of INCR bursts, the tag as passed in tag_to_pack[] is directly
    * packed to packed_tag[]. 
    * @param tag_to_pack tag to be packed
    * @param packed_tag[] Output byte stream with packed tag
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void pack_tag_to_byte_stream(
                                          input logic[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag_to_pack[],
                                          output logic[3:0] packed_tag[]
                                        ); 
`else
  extern function void pack_tag_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag_to_pack[],
                                          output bit[3:0] packed_tag[]
                                        );
`endif 
 
 
  /** Converts tag from wysiwyg format to right justified format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_tag_to_right_justified_format(ref logic[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag[]);
`else
  extern function void convert_tag_to_right_justified_format(ref bit[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag[]);
`endif


  /** Converts tag_update from wysiwyg format to right justified format */
  extern function void convert_tag_update_to_right_justified_format(ref bit[`SVT_AXI_MAX_TAGUPDATE_WIDTH-1:0] tag_update[]);


  /** Converts tag from right justified format to wysiwyg format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_tag_to_wysiwyg_format(ref logic[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag[]);
`else
  extern function void convert_tag_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag[]);
`endif


  /** Converts tag_update from right justified format to wysiwyg format */
  extern function void convert_tag_update_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_TAGUPDATE_WIDTH-1:0] tag_update[]);

  /**
    * Ensures that only valid lanes have chunkstrb asserted. In wysisyg format
    * the constraints leave data[] and rchunkstrb[] open. This function is called in
    * post_randomize to make sure that chunkstrb is asserted only for valid lanes
    */ 
  extern function void get_chunkstrb_for_wysiwyg_format(ref bit[`SVT_AXI_MAX_CHUNK_STROBE_WIDTH -1:0] rchunkstrb[]);

`endif

 /**
    * Ensures that only valid lanes have poison asserted. In wysisyg format
    * the constraints leave data[] and poison[] open. This function is called in
    * post_randomize to make sure that poison[] is asserted only for valid lanes
    */ 
  extern function void get_poison_for_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] poison[]);

 /**
   * Simple utility used to convert string property value representation into its
   * equivalent 'bit [1023:0]' property value representation. Extended to support
   * encoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit encode_prop_val(string prop_name, string prop_val_string, ref bit [1023:0] prop_val,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);

  /**
   * Simple utility used to convert 'bit [1023:0]' property value representation
   * into its equivalent string property value representation. Extended to support
   * decoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit decode_prop_val(string prop_name, bit [1023:0] prop_val, ref string prop_val_string,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);


  /**
    * Returns the encoding for AWSNOOP/ARSNOOP/ACSNOOP based on the 
    * transaction type
    * @return The encoded value of AWSNOOP/ARSNOOP/ACSNOOP
    */
  extern function bit[`SVT_AXI_ACE_SNOOP_TYPE_WIDTH-1:0] get_encoded_snoop_val();

`ifdef SVT_ACE5_ENABLE
 
  /**
    * Returns the encoding for AWCMO based on the 
    * cmo_on_write_xact_type type
    * @return The encoded value of AWCMO
    */
  extern function bit[`SVT_AXI_ACE_WCMO_WIDTH-1:0] get_encoded_awcmo_val();

   /**
    * Decodes the given AWCMO value and returns the transaction type.
    * @param awcmo_val The value on AWCMO
    */
  extern function cmo_on_write_xact_type_enum get_decoded_awcmo_val(bit[`SVT_AXI_ACE_WCMO_WIDTH-1:0] awcmo_val);

  /**
   * Sets Combined Write and CMO type
   */
  extern function void set_combined_writecmo_transaction_type();
  
  /**
   * Indicates whether the current transaction is write cmo or not
   */
  extern function bit is_combined_writecmo_xact();

  /**
   * Indicates whether the current transaction is write pcmo or not
   */
  extern function bit is_combined_write_pcmo_xact();

  /**
   * Indicates whether the current transaction is write pcmo or not
   */
  extern function bit is_combined_write_non_pcmo_xact();  

  /**
   * Indicates whether the current transaction is writeuniqueptl or writeuniquefull cmo or not
   */
  extern function bit is_combined_writeunique_cmo_xact();  

  /**
   * Indicates whether the current transaction is writenosnp* cmo or not
   */
  extern function bit is_combined_writenosnp_cmo_xact();  

  /**
   * Indicates whether the current transaction is writeuniquefull cmo or not
   */
  extern function bit is_combined_writeuniquefull_cmo_xact();  

  /**
   * Indicates whether the current transaction is writenosnpfull cmo or not
   */
  extern function bit is_combined_writenosnpfull_cmo_xact();  

  /**
   * Indicates whether the current transaction is writeuniqueptl cmo or not
   */
  extern function bit is_combined_writeuniqueptl_cmo_xact();  

  /**
   * Indicates whether the current transaction is writenosnpptl cmo or not
   */
  extern function bit is_combined_writenosnpptl_cmo_xact();  

`endif

  /**
    * Decodes the given snoop value(ARSNOOP/ACSNOOP) and returns the transaction type.
    * This function can be used for the read address channel and the
    * snoop address channel. 
    * @param snoop_val The value on ARSNOOP/ACSNOOP
    */
  extern function coherent_xact_type_enum get_decoded_read_snoop_val(bit[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] snoop_val);

  /**
    * Decodes the given snoop value(AWSNOOP) and returns the transaction type.
    * This function can be used for the write address channel. 
    * @param snoop_val The value on AWSNOOP
    */
  extern function coherent_xact_type_enum get_decoded_write_snoop_val(bit[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] snoop_val);

  /**
    * Returns the channel on which a transaction will be transmitted
    * @return The channel (READ/WRITE) on which this transaction will
    * be transmitted.
    */
  extern function xact_type_enum get_transmitted_channel();
  /**
    * Indicates if this transaction is applicable for updates in
    * the FIFO rate control model 
    * @return Returns 1 if applicable, else returns 0 
    */
  extern function bit is_appplicable_for_fifo_rate_control();

  /**
    * Checks if the coherent transaction is DVM Sync 
    */
  extern function bit is_coherent_dvm_sync();
 
  /**
    * Returns the index (of data or wstrb fields) corresponding 
    * to the wrap boundary
    */ 
  extern function int get_wrap_boundary_idx();

`ifdef SVT_ACE5_ENABLE
  /**
    * Returns the index (of atomic_read_data) corresponding 
    * to the wrap boundary for Atomic compare transaction
    */ 
  extern function int get_wrap_boundary_idx_for_atomic_compare_read_data();

`endif

  /** returns lowest address of the transaction. For WRAP type of transaction
    * it indicates starting address after transaction statisfies WRAP condition
    * and wraps over to include lower addresses
    */
  extern function bit [`SVT_AXI_MAX_ADDR_WIDTH - 1:0] get_wrap_boundary();

  /** returns burst size aligned address */
  extern function bit [`SVT_AXI_MAX_ADDR_WIDTH - 1:0] get_burst_boundary();

  /**
    * Returns the byte lanes on which data is driven for a given data width
    */
  extern function void get_byte_lanes_for_data_width(
                bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                int beat_num,
                int data_width_in_bytes,
                output int lower_byte_lane,
                output int upper_byte_lane
          );
  
  /**
    * Checks if the transaction crosses the 4kb boundary
    */
  extern function bit is_addr_4kb_boundary_cross();

  /**
    * Returns the data in the data_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that either data[] or cache_write_data[]
    * fields of this class have been passed as arguments to data_to_pack[] field.
    * In the case of WRAP bursts the data is returned such that packed_data[0] 
    * corresponds to the data for the wrap boundary. 
    * In the case of INCR bursts, the data as passed in data_to_pack[] is directly
    * packed to packed_data[]. 
    * @param data_to_pack Data to be packed
    * @param packed_data[] Output byte stream with packed data
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void pack_data_to_byte_stream(
                                          input logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] data_to_pack[],
                                          output logic[7:0] packed_data[]
                                        ); 
`else
  extern function void pack_data_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] data_to_pack[],
                                          output bit[7:0] packed_data[]
                                        );
`endif  

`ifdef SVT_ACE5_ENABLE
  /**
    * Returns the data in the atomic_compare_read_data_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that atomic_read_data[]
    * field of this class have been passed as arguments to atomic_compare_read_data_to_pack[] field.
    * In the case of WRAP bursts the data is returned such that packed_atomic_compare_read_data[0] 
    * corresponds to the data for the wrap boundary. 
    * In the case of INCR bursts, the data as passed in atomic_compare_read_data_to_pack[] is directly
    * packed to packed_data[]. 
    * @param atomic_compare_read_data_to_pack Data to be packed
    * @param packed_atomic_compare_read_data[] Output byte stream with packed data
    */

`ifdef SVT_MEM_LOGIC_DATA
 extern function void pack_atomic_compare_read_data_to_byte_stream( 
                                                               input logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] atomic_compare_read_data_to_pack[],
                                                               output logic[7:0] packed_atomic_compare_read_data_data[]
                                                             ); 
`else  
 extern function void pack_atomic_compare_read_data_to_byte_stream( 
                                                               input bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] atomic_compare_read_data_to_pack[],
                                                               output bit[7:0] packed_atomic_compare_read_data[]
                                                             ); 
`endif 

`endif 
  /**
    * Returns the data_user in the data_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that data_user[] 
    * has been passed as arguments to data_to_pack[] field.
    * In the case of WRAP bursts the data_user is returned such that packed_data[0] 
    * corresponds to the data for the wrap boundary. 
    * In the case of INCR bursts, the data_user as passed in data_to_pack[] is directly
    * packed to packed_data[]. 
    * @param data_to_pack Data to be packed
    * @param packed_data[] Output byte stream with packed data
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void pack_data_user_to_byte_stream(
                                          input logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data_to_pack[],
                                          output logic[7:0] packed_data[]
                                        ); 
`else
  extern function void pack_data_user_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data_to_pack[],
                                          output bit[7:0] packed_data[]
                                        );
`endif  

  /**
    * Returns the wstrb in the wstrb_to_pack[] field as a byte stream based on
    * the burst_type. 
    * In the case of WRAP bursts the wstrb is returned such that packed_wstrb[0] 
    * corresponds to the wstrb for the wrap boundary. 
    * In the case of INCR bursts, the wstrb as passed in wstrb_to_pack[] is directly
    * packed to packed_wstrb[]. 
    * @param wstrb_to_pack wstrb to be packed
    * @param packed_wstrb[] Output byte stream with packed wstrb
    */
  extern function void pack_wstrb_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] wstrb_to_pack[],
                                          output bit packed_wstrb[]
                                        ); 
   /**
    * Returns the poison in the poison_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that either poison[] or cache_write_poison[]
    * fields of this class have been passed as arguments to data_to_pack5[] field.
    * In the case of WRAP bursts the data is returned such that packed_poison[0] 
    * corresponds to the poison for the wrap boundary. 
    * In the case of INCR bursts, the poison as passed in poison_to_pack[] is directly
    * packed to packed_poison[]. 
    * @param poison_to_pack poison to be packed
    * @param packed_poison[] Output byte stream with packed poison
    */
  extern function void pack_poison_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] poison_to_pack[],
                                          output bit packed_poison[]
                                        ); 

  /**
    * Unpacks the data in data_to_unpack[] into utemp_datanpacked_data.
    * For an INCR burst, the data is directly unpacked into unpacked_data
    * For a WRAP burst, the data is unpacked such that unpacked_data[0] corresponds
    * to the starting address. The assumption here is that data_to_unpack[] has
    * a byte stream whose data starts from the address corresponding to the wrap
    * boundary
    * @param data_to_unpack The data to unpack.
    * @param unpacked_data The unpacked data.
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void unpack_byte_stream_to_data( 
                                            input logic[7:0] data_to_unpack[],
                                            output logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] unpacked_data[]
                                          ); 
`else
  extern function void unpack_byte_stream_to_data( 
                                            input bit[7:0] data_to_unpack[],
                                            output bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] unpacked_data[]
                                          ); 
`endif
  
  /**
    * Unpacks the data_user in data_to_unpack[] into utemp_datanpacked_data.
    * For an INCR burst, the data_user is directly unpacked into unpacked_data
    * For a WRAP burst, the data_user is unpacked such that unpacked_data[0] corresponds
    * to the starting address. The assumption here is that data_to_unpack[] has
    * a byte stream whose data_user starts from the address corresponding to the wrap
    * boundary
    * @param data_to_unpack The data to unpack.
    * @param unpacked_data The unpacked data.
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void unpack_byte_stream_to_data_user( 
                                            input logic[7:0] data_to_unpack[],
                                            output logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] unpacked_data[]
                                          ); 
`else
  extern function void unpack_byte_stream_to_data_user( 
                                            input bit[7:0] data_to_unpack[],
                                            output bit[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] unpacked_data[]
                                          ); 
`endif

  /**
    * Unpacks the wstrb in wstrb_to_unpack[] into unpacked_wstrb.
    * For an INCR burst, the wstrb is directly unpacked into unpacked_wstrb
    * For a WRAP burst, the wstrb is unpacked such that unpacked_wstrb[0] corresponds
    * to the starting address. The assumption here is that wstrb_to_unpack[] has
    * a byte stream whose wstrb starts from the address corresponding to the wrap
    * boundary
    * @param wstrb_to_unpack The wstrb to unpack.
    * @param unpacked_wstrb The unpacked wstrb.
    */
  extern function void unpack_byte_stream_to_wstrb( 
                                            input bit wstrb_to_unpack[],
                                            output bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] unpacked_wstrb[]
                                          ); 
   /**
    * Unpacks the poison in poison_to_unpack[] into unpacked_poison.
    * For an INCR burst, the poison is directly unpacked into unpacked_poison
    * For a WRAP burst, the poison is unpacked such that unpacked_poison[0] corresponds
    * to the starting address. The assumption here is that poison_to_unpack[] has
    * a byte stream whose poison starts from the address corresponding to the wrap
    * boundary
    * @param poison_to_unpack The poison to unpack.
    * @param unpacked_poison The unpacked poison.
    */
  extern function void unpack_byte_stream_to_poison( 
                                            input bit poison_to_unpack[],
                                            output bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] unpacked_poison[]
                                          ); 
                     
  /**
   * Does a basic validation of this transaction object
   */
  extern virtual function bit do_is_valid (bit silent = 1, int kind = RELEVANT);

  /**
    * Sets the suspend_master_xact property
    */
  extern virtual function void suspend_xact();

  /**
    * Unsets the suspend_master_xact property
    */
  extern virtual function void resume_xact();

  /**
    * Gets the number of beats of data/resp to be sent.
    */
  extern function int get_burst_length(int ignore_exceptions = 0);

`ifdef SVT_ACE5_ENABLE
  /**
    * Gets the number of beats for atomic_read_data in Atomic compare transactions 
    */
   extern function int get_burst_length_for_atomic_compare_read_data(int ignore_exceptions =0);
`endif

  /**
    * Gets the burst_type of a transaction.
    */
  extern function burst_type_enum get_burst_type(int ignore_exceptions = 0);

  /**
    * Gets the burst_size of a transaction.
    */
  extern function burst_size_enum get_burst_size(int ignore_exceptions = 0); 

  /**
   * Gets the minimum byte address which is addressed by this transaction
   * 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Minimum byte address addressed by this transaction
   */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_min_byte_address(bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");

  /**
   * Gets the maximum byte address which is addressed by this transaction
   * 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Maximum byte address addressed by this transaction
   */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_max_byte_address(bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");

  /** 
   * Checks if the given address range overlaps with the address range of this transaction
   * 
   * @param min_addr The minimum address of the address range be checked 
   * @param max_addr The maximum address of the address range be checked 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Returns 1 if there is an address overlap, else returns 0.
   */
  extern function bit is_address_overlap(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] min_addr, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] max_addr, bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");

  /**
    * Returns the total number of bytes transferred in this transaction or beat number
    * svt_axi_port_configuration::get_byte_count_from_wstrb_enable set to 0,
    * the byte count is calculated using burst_length and burst_size based on
    * @param beat_num Indicates the beat number for which the byte count is
    * to be calculated. If set to -1, the total number of bytes for the entire
    * transaction is calculated. 
    * If svt_axi_port_configuration::get_byte_count_from_wstrb_enable
    * is set to 1, the byte count is calculated using wstrb based on 
    * @param beat_num Indicates the beat number for which the byte count is
    * to be calculated. If set to -1, the total number of bytes for the entire
    * transaction is calculated. 
    * @return The total number of bytes transferred in this transaction or beat number
    */
  extern virtual function int get_byte_count(int beat_num = -1);

  /** @cond PRIVATE */
  /** Converts data from wysiwyg format to right justified format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_data_to_right_justified_format(ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] data[]);
`else
  extern function void convert_data_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] data[]);
`endif
`ifdef SVT_ACE5_ENABLE
  /** Converts atomic_read_data from wysiwyg format to right justified format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_atomic_compare_read_data_to_right_justified_format(ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] atomic_read_data[]);
`else
  extern function void convert_atomic_compare_read_data_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] atomic_read_data[]);
`endif
`endif
  /** Converts data_user from wysiwyg format to right justified format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_data_user_to_right_justified_format(ref logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data[]);
`else
  extern function void convert_data_user_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data[]);
`endif

  /** Converts wstb from wysiwyg format to right justified format */
  extern function void convert_wstrb_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] wstrb[]);

  /** Converts poison from wysiwyg format to right justified format */
  extern function void convert_poison_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] poison[]);

  /** Converts data from right justified format to wysiwyg format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_data_to_wysiwyg_format(ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] data[]);
`else
  extern function void convert_data_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] data[]);
`endif

  /** Converts data from right justified format to wysiwyg format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_data_user_to_wysiwyg_format(ref logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data[]);
`else
  extern function void convert_data_user_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data[]);
`endif

  /** Converts wstrb from right justified format to wysiwyg format */
  extern function void convert_wstrb_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] wstrb[]);

  /** Converts poison from right justified format to wysiwyg format */
  extern function void convert_poison_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] poison[]);

  /** Turns-off randomization for all AXI3/AXI4 parameters */
  extern virtual function void set_axi3_4_randmode(bit on_off=0);

  /**
    * Returns the contents of data as a string. 
    * @param  xact_data A byte stream array of the data which can be obtained through
    *              the pack_data_to_byte_stream function
    * @param  xact_wstrb A bit stream array of the wstrb which can be obtained through
    *              the pack_wstrb_to_byte_stream function
    * @param disable_msg_info Disables information regarding message format
    * @return The data as a string. If corresponding wstrb is 0, data is marked as 'xx'
    */
  extern virtual function string get_write_data_string(bit[7:0] xact_data[],bit xact_wstrb[],bit disable_msg_info = 0);

  /**
    * Returns the contents of data as a string. 
    * @param  xact_data A byte stream array of the data which can be obtained through
    *              the pack_data_to_byte_stream function
    */
  extern virtual function string get_read_data_string(bit[7:0] xact_data[]);

  /**
    * Returns the contents of wstrb as a string. 
    * @param  xact_wstrb A bit stream array of the data which can be obtained through
    *              the pack_wstrb_to_byte_stream function
    */
  extern virtual function string get_wstrb_string(bit xact_wstrb[]);

  /**
    * Compares the contents of two byte streams. 
    * @param  xact_data A byte stream array of the data which can be obtained through
    *              the pack_data_to_byte_stream function
    * @param  xact_wstrb A bit stream array of the wstrb which can be obtained through
    *              the pack_wstrb_to_byte_stream function. If xact_wstrb is 0,
                   corresponding xact_data is not compared 
    * @param  ref_data A byte stream array of the reference data to which xact_data must
                   be compared. 
    * @return Returns 1 if the comparison passed, else returns 0.
    */
  extern function bit compare_write_data(bit[7:0] xact_data[],bit xact_wstrb[], bit[7:0] ref_data[]);

  /**
    * Compares the contents of two byte streams. 
    * @param  xact_data A byte stream array of the data which can be obtained through
    *              the pack_data_to_byte_stream function
    * @param  ref_data A byte stream array of the reference data to which xact_data must
                   be compared. 
    * @return Returns 1 if the comparison passed, else returns 0.
    */
  extern function bit compare_read_data(bit[7:0] xact_data[],bit[7:0] ref_data[]);

  /**
    * Gets a single response status based on rresp of each beat or bresp.
    * If it is an exclusive access, then this function returns an OKAY response
    * if all beats have a response of EXOKAY, otherwise it returns a SLVERR response
    * For normal transactions, this function returns OKAY only if all beats have
    * a response of OKAY
    * @return Returns the combined response status of all beats 
    */
  extern function resp_type_enum get_response_status();

  /** Returns first data_valid_assertion_time for read channel transaction or write
    * response assertion time for write channel transaction
    */
  extern function real get_response_assertion_time(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] cacheline, bit tagged_addr = 0, int mode=0);

  /** Returns data_valid_assertion_time for the beat number of given address read channel transaction or write
    * response assertion time for write channel transaction.
    */
  extern function real get_response_assertion_time_of_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] cacheline, bit tagged_addr = 0, int mode=0);

  /** returns id considering only the bits which are used by exclusive monitor */
  extern function bit[`SVT_AXI_MAX_ID_WIDTH-1:0] excl_id(bit use_partial_id=1);

  /** returns address considering only the bits which are used by exclusive monitor.
    * However, if num_addr_bits_used_in_exclusive_monitor is set to -1 this indicates that, user wants
    * use specified start and end address ranges for each exclusive monitor. In this case,
    * this method will return exclusive monitor index with tagged address attribute i.e. secured/nonsecure
    * bit, as exclusive monitored address. This models the interconnect's behaviour of monitoring
    * different address chunks.
    */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] excl_addr(bit use_partial_addr=1, bit use_arg_addr=0, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr=0);

  /** returns address aligned to cacheline size */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] cacheline_addr(bit use_tagged_addr=0);

  /** returns address aligned to snoop data width size */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] snoop_aligned_addr();

  /** returns the status corresponding to the status mode value passed */
  extern function status_enum get_status(int status_mode);

  /** Outputs the expected snoop addresses. 
    * If the transaction does not generate a snoop, the function returns 0, else it returns 1.
    * However, if include_non_snooped_xacts is set, the function includes WRITEBACK, WRITECLEAN,
    * EVICT, WRITEEVICT and cache maintenance transactions sent to NON-SHAREABLE region as well.
    */
  extern function bit get_expected_snoop_addr(output bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] expected_snoop_addr[$], input bit use_tagged_addr=0, input bit include_non_snooped_xacts = 0, input int cache_line_size = -1);

  /** Returns 1 if this transaction type generates a snoop, else returns 0 */
  extern function bit has_snoop();

  /** Returns 1 if this transaction is a full cacheline access, else returns 0 */
  extern function bit is_cache_line_access();

  /** Sets the port kind to master or slave */
  extern function void set_port_kind(svt_axi_port_configuration::axi_port_kind_enum axi_port_kind);

  /** Returns address concatenated with tagged attributes which require indipendent address space.
    * for example, if secure access attribute is enabled bye setting num_enabled_tagged_addr_attributes[0] = 1
    * then this bit will be used to provide unique address spaces for secure and non-secure transactions.
    *
    * @param  use_arg_addr Indicates that address passed through argument "arg_addr" will be used instead of 
    *                      transaction address "addr", when set to '1'. If set to '0' then transaction address
    *                      "this.addr" will be used for tagging.
    * @param      arg_addr Address that needs to be tagged when use_arg_addr is set to '1'
    * @param      use_cacheline_addr Indicates if returned address should be aligned to cache line size
    * @return              Returns address tagged with address attribute of corresponding port
    */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_tagged_addr(bit use_arg_addr=0, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr = 0, bit use_cacheline_addr=0);

  /** @param  arg_addr Holds Address for which untagged part needs to be obtained
    * @return          Untagged part of Address "arg_addr" will be returned
    */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_untagged_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr);

  /** Sets transaction attributes from tagged address.
    * for example, if secure access attribute is enabled then security attribute of current transation can be set from the tagged address
    * passed through argument or current transaction address.
    *
    * @param  use_arg_addr Indicates that address passed through argument "arg_addr" will be used instead of 
    *                      transaction address "addr", when set to '1'. If set to '0' then transaction address
    *                      "this.addr" will be used for tagging.
    * @param      arg_addr Tagged Address from which current transacion attributes need to be set.
    */
 extern task set_tag_from_addr(bit use_arg_addr=0, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr);

  /** Function that sets xact_type as COHERENT if svt_axi_port_configuration::is_downstream_coherent is set */
  extern function void set_xact_type();

  /** Function returns xact_type as COHERENT if svt_axi_port_configuration::is_downstream_coherent is set 
    * If not set xact_type will not be changed for the particular transaction.
    */
  extern function xact_type_enum get_xact_type();

`ifdef SVT_ACE5_ENABLE
  /** Sets the atomic transaction type */
  extern function void set_atomic_transaction_type();

 /**
    * Returns the encoding for AWATOP based on the 
    * transaction type
    * @return The encoded value of AWATOP
    */
  extern function bit[`SVT_ACE5_ATOMIC_TYPE_WIDTH-1:0] get_encoded_atomicop_val();

 /**
    * Returns the decoding  for AWATOP based on the 
    * transaction type
    * @return The decoded value of AWATOP
    */
  extern function atomic_xact_op_type_enum get_decoded_atomicop_val(bit[`SVT_ACE5_ATOMIC_TYPE_WIDTH-1:0] awatop_val);

 /**
    * Returns the decoding  for Endianness based on the 
    * transaction type
    * @return The decoded value of AWATOP
    */
  extern function endian_enum get_decoded_endianness_val(bit endian_val);

  /** Returns the inbound data size for atomic transaction */
  extern function int get_atomic_transaction_inbound_data_size_in_bytes();
  
  extern function bit is_addr_aligned_to_total_outbound_data();

 /** Returns the masked atomicop data based on current atomic xact data_size, input args data and byte_enable */
  extern function bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] get_masked_data(bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] data[], bit [(`SVT_AXI_WSTRB_WIDTH-1):0] wstrb[]);
  
/** Returns the masked atomicop data based on current atomic xact data_size, input args data and byte_enable */
  extern function void get_masked_atomic_read_data(bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] atomic_read_data[],output bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] masked_atomic_read_data);

  /** Returns the masked atomicop wstrb and  data based on current atomic xact data_size */
  extern function bit [(`SVT_AXI_WSTRB_WIDTH-1):0] get_masked_wstrb(bit [(`SVT_AXI_WSTRB_WIDTH-1):0] wstrb_);

  /** Performs atomic operation at beat level */
  extern function bit perform_atomic_operation(input bit[(`SVT_AXI_MAX_DATA_WIDTH-1):0] masked_atomic_read_data, 
                                                input bit[(`SVT_AXI_MAX_DATA_WIDTH-1):0] data[],
                                                input bit [`SVT_AXI_WSTRB_WIDTH-1:0] wstrb[],
                                                output bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] atomic_resultant_data_
                                                );

 
/** Unpacks data into atomic_swap_data and atomic_compare_data field. This is applicable for ATOMIC_COMPARE transactions only */
   extern function void unpack_data_into_atomic_swap_and_atomic_compare_data(input bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] data[],int beat_num);


 /** Unpacks atomic_resultant_data into beat_format to do the beat formation */
  extern function void unpack_atomic_resultant_data_into_beat_format (input bit[(`SVT_AXI_MAX_DATA_WIDTH -1):0] atomic_resultant_data_);


/** Performs Atomic xact operation such as ADD etc. */
  extern function void perform_atomic_xact_operation(svt_axi_transaction xact);


 /** unpacks wstrb into atomic_swap_wstrb and atomic_compare_wstrb into field. This is applicable for ATOMIC_COMPARE transactions only */
  extern function void unpack_wstrb_into_atomic_swap_and_atomic_compare_wstrb(input bit [(`SVT_AXI_MAX_DATA_WIDTH/8-1):0] wstrb[],int beat_num);

`endif
  /**
    * Indicates if this transaction has poison for any 64-bit chunk 
    * @return Returns 1 if poison is present, else returns 0
    */
  extern function bit has_poison();

  /** Marks current transaction as part of multipart dvm sequence to avoid irrelevant
    * check being performed on this transaction.
    * Since only first transaction of multipart dvm transaction sequence has control information on LSB[15:0] bits,
    * it is important to set this bit to '1', before randomizing the second or later transaction object so that, 
    * second or later part of multipart dvm sequence can ignore dvm address constraints for control fields.
    */
  extern virtual task set_multipart_dvm_flag (string kind = "");

  /** returns first beat of coherent response of current transacton */
  extern virtual function coherent_resp_type_enum get_coh_resp();

  /** returns '1' if current transaction matches expected transaction type i.e. for coherent transaction
    * if it has matched coherent_xact_type and for non_coherent transaction if it matched xact_type, otherwise it returns '0'
    */
  extern virtual function bit is_type_matched(int rw_type = -1, string typ = "non_dvm_non_barrier");

  /** returns '1' if current transaction will allocate a cacheline but, there are at least one transaction currently active
    *             which will attempt to de-allocate the same cacheline.
    * returns '0' otherwise.
    */
  extern virtual function bit has_overlapped_dealloc_xact(int mode=0, svt_axi_transaction ext_xact=null);

  /** returns '1' if overlapped transaction between read and write channel found else '0' */
  extern virtual function bit has_overlapped_rd_wr_xact(int mode=0, svt_axi_transaction ext_xact=null);

  /** returns calculated parity value for 8bit of data */
  extern virtual function bit parity_bit_from_8bit_data(bit [7:0] data, bit even_odd_parity = 1);
  extern virtual function bit parity_bit_from_16bit_data(bit [15:0] data, bit even_odd_parity = 1);
  extern virtual function bit parity_bit_from_1bit_data(bit data, bit even_odd_parity = 1);
  extern virtual function void parity_for_xact_field(input string xact_signal_name = "", input bit even_odd_parity = 1);

  /** returns calculated data check parity value to data */
  extern virtual function bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] calculate_parity(bit [`SVT_AXI_MAX_DATA_WIDTH-1:0] data);

 /** returns converted  data check to pison value */
  extern virtual function bit [(`SVT_AXI_MAX_DATA_WIDTH/64)-1:0]convert_datacheck_to_poison(bit [`SVT_AXI_MAX_DATA_WIDTH/8-1:0] is_datachk_passed,bit [`SVT_AXI_MAX_DATA_WIDTH/64-1:0]data_chk_to_poison);

  /** returns '1' if transaction passed through argument i.e. overlapped_xact is found active while
    * current transaction is found active or in other words both are found active at the same time */
  extern virtual function bit is_overlapped_in_time(svt_axi_transaction overlapped_xact);

  /** returns '1' if current transaction will allocate a cacheline else returns '0' */
  extern virtual function bit is_alloc_xact();

  /** returns '1' if current transaction will de-allocate a cacheline else returns '0' */
  extern virtual function bit is_dealloc_xact();

  /** updates num_xacts_blocked_progress_of_curr_xact with number of xacts that blocked progress of current xact */
  extern virtual task update_num_xacts_blocked_progress_of_curr_xact(int num_blocked_xacts=1, int mode=0);

  /** returns '1' if current transaction is not supposed to return data as part of coherent read response */
  extern virtual function bit is_read_response_without_data(int mode=0);

  /** returns '1' if current transaction will allocate a cacheline in L3 else returns '0' */
  extern virtual function bit is_l3_allocate(bit is_exclusive=0, bit is_partial_data=1);

  /** returns '1' if current transaction will de-allocate a cacheline from L3 else returns '0' */
  extern virtual function bit is_l3_deallocate(bit is_partial_data=1);

  /** returns '1' if current transaction is supposed to update memory with L3 data */
  extern virtual function bit is_l3_update_to_mem(bit is_partial_data=1);

  /** returns '1' if current transaction doesn't cover full cacheline */
  extern virtual function bit is_partial_cacheline_data();

  /** Returns number of byte whose wstrb is '1' */
  extern virtual function int get_valid_byte_count();

  /** returns '1' if current transaction is determined to be valid exclusive type */
  extern virtual function bit is_exclusive_access(string mode="", bit shared=1);

  /** Sets the channel on which a transaction will be transmitted */
  extern function void set_transmitted_channel();

  /** Returns '1' if write strobes are driven correctly otherwise, returns '0' */
  extern virtual function bit check_wstrb(bit silent=0);
  /** @endcond */

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_class_factory(svt_axi_transaction)
`endif
endclass
/**
Transaction Class Macros definition  and utility methods definition
*/

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
JCYU4R/6ZnFfuq2QSUc/ieJLarREoDeboPvGKMHTHGyuuwQm8Vb7g16D8ncVhwEo
erxpQeLy73ENSZsq++jO+aGmgicTf1+neTMIQPcxLAhjXY9cVgOgsVnF/1jZnQ32
BCE4ArPOjIb2zJWXuMkGy2kDf0l1/Sy6MIXfckcgy2k=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 4321      )
4IcIUoRu4tVw+TPlDFJeEqfLtWz5I+sUQXE3TpEknNYlsDKldX3WY/CTkD8cMjYT
kOm8baD74illRfIvX/wii/MF0sdiI08JiT/yugrqoe/JssZcjD1bVUSTDbaBaBM5
x1cCzZ3Gvg9dLdGH2uXqa6oh7ixaZMvHhYmZqDbWsNrzFZpBPQTRpP82yiFy+qlK
XltbYTu92DWrTtB5vOzR5tVFvA8VR66kn3bL/N648VuatPv9h2Mzxhgbr/FI6MBW
Fqd1N/wkqHzA11OiQl2cR76IucBc/4LZojLoXOic8mhlGso7VfJL45+A3xq9R2Ni
KqdBc6G2Yfrb6K+u6i8+PRlD2zk/rrzu5oNCTLC6HdlLSny2mpfs+a0NXzhwWopV
kb5Pnm11vS2tK0MImB102vBQlkd1VN9c6CpToJOwnwlpKeA/DC14CMe4ig6AYk9N
1FA7NzJ2yP6ofo1XZElBdveVFNZpKJEP0fLVUpcEBriT2SpwY9PvfV2J/bpJcLVm
KqibchFUY69G5UwbvtLpOQAxI94HWAdVPb8w3cD3pTO25SwgmJ9YVYnvp2pHUq8G
ZTOWXl/pXi43OXOPxvqE8Dn6X/9v1n9FVZgCsG6p1TzHJUn0sOngadCYPfpbGnPW
HxB+7TubgkFu8pBRTRrBB1en8WdLVvFODd0j2YeHsYVN/AasCVsfJRzAZGZKIRxU
F20WQ7IuxTRfCtnUSwobfIK6nhAvL64f6g/73mPz9X/dyxxcrduAfMhmf3edOItz
53OiD1FGkQgYpUk4HCJWefGTkTHga9Yg3VCgp5ugxPQ1gB7nmrovg32szKFopysn
vQZfgU45Ikzx9uXjiBnGcixya6Cxv6U+BOC3th3JmaqTpfYX9w4X3xtAExfZ3CtL
AsAvjf4GrRlGc+JAkBbouWtcr+8EJJRFtCPsds8JGW6D/5csDuae9QTCtK6kyZuA
ONE4Emt34GcSvZhoB9CnVFfucVPyrplO3emE8sILBRT128ktDS5y5akiEkLd0FCT
Q2SKXVZcCSDOqFgttJPoW+hCn3HXFu4wUZPwjAEi7vaORtvO+f+Q/f10FAJBwJsJ
EJHDZogyltgw8dXm8VnvjYYIi8uasQQIaNrPJgVzEktpd1VauMp4H9aneX6ipxkC
Y+dtsuqSwxGgRF3eq5mxZn5/jqjBPJsXFGIdOGFG9FvHzS6Jm0BL/Y8xbP6nzpX6
3z5BCsIXj9TWaiEWasS1q/cKpM9mP9DdHUH4Rt86Aa2N1DELPrLjWW02Pp9omN/o
Rrjn8ShcWmO+VRUHsrhVxZY1pJaAm17BJkbd6DXyFutM2CtEPxvr4qnwln7Cl3ic
IWaDrlxSXSVTgXju8J1cpA4ZSWZ4rruYDfQ16AZ+tSVQT48B0qYyhN0gZ1jRg+Il
Se5B8GaN3WheLaRq4qnaZ3dQu4jipvcfAyJ+F93NqZZ5OvlpnkeEQwtnm6wt3f4N
eraQiEXbRfFzedDBU6t4lTn5abxgkLI35CGucZgaZtFQNff1MiKTQjjJ9C9hJe+A
ylH/OGlz7CjvlPKMxHeQ0aTUBjNeAr/R0Kw4urkQIM5XRlGe3oIFvEXaJf3QNlFU
0FH8hETqdVt+MH03LX7cj1PHEh5sy2yeWBTE0UEZLqschOl1Ts6hnaAE4GNnnt9j
FQERdDswBWkIEJGK4jiG4DO0sHXq3TSENanCT8iZVLsaPXxr4w+goLfLEvOrUTqE
6bx5fp94k14ZQL/lmEl3FzZoPFxXsm7U3OYdooYvm9pPCccoiX/TO6L8AZkvzP3A
Xb8PV0MtGPenIzcSa70bOGGIk0YGhBAVeem48YMroZFyIclu151Edv9c8yRC0yzu
T8JXpgWxol2QovpJpa97QrJPULdMcQc0+4eUyOIbr8OIxS701TysI26Y3OpmnoAr
mz1axvCAe5snpvFtQXSmWbQOnOhiscIgXI4jO6m0I01sd+od8nNHYzaM4Wd4j+V6
rXhNrGQw9+bP8zNQgTXXnzxbMfxpFnuk+vRDagYmFCmpJxwBkUx/hmUaEC+sanc/
Yy/PZ+QGYNUXKzk9SFXHzTy3jSqfvIrMmJuVibB9xLEx6Rp65GZEX0HBCuVy+ORs
GBp8L+mao0B3L9MSW4fHWo6cX0ambU9RR6K63RDeL+DyZwk7eIDNJYbhHz0wJlMy
jBRvEb+HuXtbv1pPLFZEOaSy8+W9dqJ59sdSR1CE3bi0pxKg4jae80Q4foPmMTwm
lAHJo4UA0/wfIPOxksAaboceqUEUOZhUZRXdWOVpGeangbln62YRgbNVG7m3KO98
YUQ80vUgHtNiG2XdxjBYqRgM6eZh9Zmlu3tIfZ3d8gFePjTE9zVL078amdhxIfOD
PKM88lKUpzCpEmtyfy+Rw1yvgkUOAQhS+zv4W/4YUNka8eig9Vq55/2GLu+3CWb6
PBf2LlPXkngv7XORwhEbbkaLCXYvAqumVYqREaFHdAs+2BYyWVWLgoPb/4Z3U13A
Hhhd7kEYHqWajac9UT9zFVZjv2RWXDV0AFUcRIZDD6CXvIVgt0mbcXDxEOTjm0nG
lNt9s9xzF8OPVZCJlSClyD8Nsw1AEYs8D4/nRyViWIABDLd7Vf+azsbFemqOBaEa
9ei3Ra763O9wZb9+/8m0+VGnu1pLo5ZVbDEBOD/lSZWEQV9/o74Rfjtc8w/9EfY6
xM339ORt5sHH6hmEMcVrCxSMuFNjiF1D6QlrK0fuHLMK9bcBML1S7JD0L/pILR1/
9PV4K7J5omf1EDb+jxfGcKNj6hGfHW0+lOI0kFJ01UBNeomUWdhodQQgJubZiuz0
LX1BBugD+iRRI1Tg5U0EP9d1cr9Ogc2ZkJI1OZZ3uqf9RKhQeczCNAGwFE3JULdo
+0w0TDWAZZDJTmnYl/eWI3zcQwxSfkyc+EHRCYzAmz3HoRRtfp/6oWXea2YZs55t
sSSL867+F3O7J5Nm/DbxANhC8+dosAquT4tLnwt4K68vxpVQmDO27hu4cmZRKsBk
EyuxFkcb/w8xmf6HAi2Q58Bs1wgAp3qBRY1ZLi6nGdNLGRl7Koy8vkHNPRoEeBFk
eNCHZT2RDL0H+Knk7TcVnkkfic9L0QfPcFHKTnP2NL3juUmW31gEf/yb88UDBvkH
Bhixo5NR1vQxkgTxorOMUHg62O1rqRmxLYiE0EidJLTyHu4zLpZktNw9D6tV9+M0
VfdfqaRb1+N+LuSY4fMtbjF8dIIhn/3H5F/RGkLYnUFko3EgbNHOeM5AuBeS1vEx
VC8BIDsFLsHpj9jhzpbRHSm341fjkxB6B5AMQETUAY5GpO/HqPz9JNVs4prVZRAU
X5wvWgySTFT6pYih+DhGfk8hJ1I+KcC0lYxCJG2cmPktfmM0SDwwFidtnSklENE8
RvVD97Pkdzw2IbuPD3EXr4s8OaIfp5xtZQHn+SZW7pCKSP38bxVeflWqqhbuzM1e
RImhG138fu3yFCOE3V+vJDYaqeJmaqujd6C97piaIxp98R0VgjJv10OkBUFEFets
nLgig7pdoybYalHT6CcSNBi+Z1FA4gZSLKdXi8cH0uIaCnc/WbU5rBQUE3e/qFTn
emRqdroVRiOyTrc04LuQQJvi6RCkCkXJikDLnYCeEeo4mcFbEH6gemVFvReup4yT
Pr+ID4Bk0/89vUSfdSQh6+5pvufzH8jHozhCJ/imL6x3ZsHw/rXgB571qCKJNNae
puqjmGQo+uzDvzEUpOu2S3J89agrwkije72ZeCf2J0Ay+MKZKPbNXCihUz9Sz0AS
nKznLON8kmUTPQuz2c6B1Y8x+xa37ePRXFCt/Ef826THhNfyYuu+V62q6PTjul+H
swsZ4XxbZx9/YbgBZRZ/VzG6ds+K+ZL+Yciq/u/E9jYU5SUAcZdc7ycUmCev07+j
/QMdB62TjfEs80sGyOEB0FGqtIaAC2NcX4cPv7du306Vbt03/DudvhKwJfUJ6DW9
7Qic6RfEfQf+tWAN0RWcFmgdJNUgaq4FPpk4gS5Agrs0yeNlY3BQO4/K5Yp1Zi54
68O7c2uwBgNbgXs+myGJAZkhZ3r+A7giIiLPPhrcd9+gm8GOkW+Md7beyFrK5+/X
eIxULtNiOpXSSSI6mElD2Vi8JTQrUQyKYyLUPztYC025GAfYPXcp40icXau/fLPc
aMfXtZxgf6dj6iFyHrGdOWSsr5noYZHZAIN966Op3J1OadQsMG69+W371VzNvun4
+qHjTjg3A5+nhQfPMYgmWuqiAElnZc/96iy+R73+scyg5B2/YrR3StFuqmgVP/C4
fwvriK2aLIygGF/lA5T7aSTs18GMQZnFAZ0sD+VAKE5GrPXC00B+PELk3wbAjqSD
2pj5h65e1m0tkoYB/hGlEMKyZuQb/K/gJc3+tdF91PgAXBah5726mCJV1jKuhz0l
gDg+JxFVGbDoGCtjtWVJ5NuusMKLpWRXBEnz5uCCwfSJQpWXqBVXByNX1yvrfSFy
vZt4LnncPBD3cDTzVHPbCshzwfmKy/uP0YDs5lPu6EaYTXNxnpXUHgCbpOqSf4gl
LKg9QGnmrBLQwMLXN9AS28MYW9+BA+TmyIyHK54GweeXfRF9UwFnod7VSbNv0n9G
jdPqi8BzNypTFSzCtFfsQL4Yuqg5rlFiLyEl8XJgnrrTNKQe/uTFcbVqZWeRdWM9
GOPd/Z7+9LKec3pz54SwByCJOIC/5LpC2693Jlp6BJ14zHtVTLU2IXu+8kle3YrA
B9IjtK8HEpJWEv6EhTx6aE1GQrtbSvhiNPuxKQKwtYyAcaTDfCu+vLuRyB8nqijE
LZVWCJEqD5opdVJU49L6ExXwODB2aNR7TM6e2GWtjmz7JYuG2cDmBQIoYxzw90MA
3mvQ6QjJvsFCYxaDHuZlTXaMK7z1hogK/SAGbjViXiVX8uQKUeNq+FkN3zQuBrde
41yyNMZ17n1ENwJJ2Gjliqkg74Ue7nGc9P1N3cNKaX0=
`pragma protect end_protected

function void svt_axi_transaction::pre_randomize ();
`pragma protect begin_protected    
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
pQBWoxsMLH9175Xn5MZWpKvvihAePQHhutX98rT6Yd0UJ2uMs+cNzslmGgM/RjBI
6ns/HBoCwdOq2mVg5yFnnBSzd3/p/lenqHpjbykOJi/FvR+W/IrhqFK4GvWrgNgy
VeP7idnK9BAjSZB2MoYgKHCCZG6XEBz34BpvzWWeh9o=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 17471     )
HZwNuzESZUu7Jj578iXvcphbrDlhy6Pi5YCN9TwOyhUe/aDDGig6SGsCP8wX2ZNE
6bmILimz/cOPiRm9858jv7JGssty1RR/n2FNUp5kmaOWh5RLUjp5tz2n7b0eoEmP
mElOx0vYZ8pTs0oA9a3Ur58sfs84Mnr66NCfHglBspVy+cYwOYcxbzCE0irIJiiy
+R09q5z5vtfxL5Iw1AQoi4inh+XxjaGxrTn4/dHS67W7OsxchP1nagAvBY+UsSnW
EorKEmLUS/CzlUKtZGx1jZTO2hBJs/VMe7+rhsr+GlqYKG97XChgLuOqDs0chufy
/V/VE3ICfjuct1S7vcgB237lHRWOCr/1HZULryyvVztLkCWEyRCKTaKo1xA0S+Wc
9qX7SksrQaOAcQZdZtZ0MJ/1H4s5LzLovrt3RfwCE5xCJw/p04AvsDypuW/YtLrX
LSY34u0DbaOspXlgVpTdwTXB+WtBavFoRXhBdiUIgyXorcESIQ5VNLlLEOIDV+kC
YsUJiSoHQxBV3HNZZMY9UF8FhPx3D7sIqw84If+ml/Ds2ewYpm2hI/ZhRJ12YeDB
vFAzy7gj4NBfalmAmSMIfdQCghczNxUChmCr02rOeeEjyy4O9jQFelklXRFtRc19
Scv2GYmwdgzRpQId0EExWsxFtfAwgPISAFKPx+G0iVJm9L6zZrRX5GkugNfKkxZF
rNBlaihZEc6yh3Hg5h39wdqeNcIybZJe6KJiEWh4KF4zLakMuE/g9f2xrPO84Ncg
XVJ/EHRIVpINbcz05Db7aWBVwn39AQNes3saWfVG9HZmDv5aIre/s8J2SGqaxgb0
O7kaLaERm8Vzm24H+K7dmQxSu8vwCXJFmrINky0NjUCD/vusjU32Kuk6lYEQnQSO
xtPwe5UclRBs88c7d3E+pTMkHhW6YrLjEW3ks+OyE4bbWrDVary2/TU2T0HWrX6j
lH24Wy/v7ER6l1RWDWYiLFWkSSoQd04s/ccAoUpRFVTk+hbz+R47obqK2aBndiov
mkBwN+oFSicQj8AfomBILi+eN+2y1a7/4pY4+ei1nTe+VglGyvFF0VrHFK9SQFDi
NEaN4sIo8G0gxMxwcXEDo7Uw/fvaGozOVaccmTTx4ZfIaKMulqd2KT7W0eW6ng2F
8ZpaATgJ0UM9O6LtB5Jt+gAHAwanIUkABCUOWi0EXkRVhqbzf9XA94uc7FxodhEl
yVGRdfttTPVaz+PXQ/ZenJMJtQPjaldyMOOPPgklFOt6Kvwz+tekTSclzy5eY4cq
1f1eL1NuiGoYO/jARGkQIN8axybg0NMAisj5wW7UAXXDJL3zNDp9TktxV6fCMQkD
RQA2o+ncPx2/TOzzrKYTpRUtt+D00gYvXkLUa+7N7kOjACN+7sMoWlK92qXkcgdu
RAUAqINRONTQC/Cwju7jLxLfq8GdLphAjRZqKo/gLqv221I3EVUdEfETYLJQMkFI
CvdFFUoWBTYhoCGrKOnd1+2r3dty3RpxYdDdwA0W/XTyhKQH5MCEuqp8rgQ/BEfw
UCHCzgV1Y5ICJmSfucLIbMjeYw0ef9w2YzOyAguO/r1lDX7I/3CFWLP2PA/Zb9iK
fzmQhBDKBWUhRNo/UmIR6XIUGMOM9cfwFuE0k31dK+TySDdxSDJlksiknY/TTt3Q
Xcj4HLtgGVCWE9o23ehhHrikZRZ7hzI3DfKKpIlwfZt3XQzHs6mvbmtJUGakbZfS
TURWwjCONuDKZ19LiwjqpRhaCJ2N24Q2KaGRv74sRbG0/yaT2dMpkzgLrd/UQjwW
ZNiQw70l+EnJVfpEP+ZnlZnvh5UEYMLfVD6Uej7EELjtnsjbp5NT4l4oRS/ZF356
lRc4d0TK442fnAEODzqOwaJEaj8on/sh/Scdb7OImQkaIkrzj5K+9hSqBlgAGHyl
pUka0PM6glh6ioMazMUtOxyYHwdLS4nJaMiuZxpkJETb8y+UrbtWvYdsrsnsmE19
kqkVG646xAHGOb6wArAzDrxWd1II3hhT0GAA9fTwS9yGkbUS2xV9eqey0a5Z8fJS
y+iwl07QqWJ+kyNni+JSx2cthgRnY9p2F1vxgvTBwmWZTPTtKoilGwR4C0t5mYUE
ZS1a21GqjdfBJF1/rLsSsJIJqeAuGtw3zr56/HpezQC1WnEJ4w7e84cY0oqfigZM
ZclwnAm+K9FG2F/F5yExE2TORmOxqlDV/tfIMF7DzjYmIDrfsD9/afUIYCqJll5O
5/o9fMXFBsrChEfiMa2RzCSI8277A78sDQPWfpDFd428aAW0HUUSGg1D4kTTbEPz
kUR1BWPk3Ex3YeAfov79gUBKxXTHd9tWgtuBijqbAfNsGti7Y6Jc3HgA7xB+856Z
stHES8CBUZ95Ql6wSoI7L17/hcHFz3ZKQu1AUl6xoDGOvv1vZmvAsiZMVvFSSqci
psoeYiJVQ3sv61b+5iZfLjx3834SkthZJlbSAcmLoshrL5TFp7q2sUJ6hfIaOBIQ
kkVqkwY+RA2GMObhRofnguH45TwWTavos1JJFFClsnF6rGSfudNH/MFUe9HdqQ5T
El4CLlA/1iPBx2tyhNwZhYdhtkz0xZnlI5iJ6Ttpw6oF7lxn6mmuUGHPv925DUJD
1L7cOHn2olcOTwOKU22S+RuJVZb76wrU0r9FzQlwJZekBI4jAlOizb118ycNFcKY
3gE47RCHNhiRdWE7nat4KFUQS5E7WOG9cAyhdhP3C4J0ZocMAsB4weaRLTZI5qtR
ovFTzeT7sNdIWHfWUBhkdFjyiZ5plAI2ENFe0lxAsyajOLXPpyFWCRhclqGt04MP
7iocdGZhItLAGs9zCy5kdps26Pk56BApQMEXLkxr/m3DZTP4F6RXbU6mJPX4VzJt
XNIN1gg7bJ61/NmbSYW4G4wVUU4fKoEb7t6dmIIraxCpnUi2n5rdT6yRqAB6kB9I
L8K50pmtUBvgPR8FiHzeV4bTiRuxWYCvpFup92D73qc2vPn4LFBv4P9ASkTxiaik
BAHtc60NbNXEbERpBsjIcE/CaT2BUFHY2wEKCxtjnTVv/0VjLEIqhbs69Dwdq4GC
RIaTVb020aY0G75LRveGeEfe9AgGJsGk8iP4W9fKEJuUKQ1u8B8MsXOUVsu7o/Pr
s3eDQK5vbfD1yUa5piCut5rNdmfGUvQLHBQ7i/wtlLo3pJ9i0ptuff4kBgeOaGR+
N3BgdWK8sXOU2qPcdDdHLlpyIevLCdaob1qoaQnqdCgPTC1LrMiziGgwMNfuRte3
MCGVQvkIFzrgESYqv3jQUmaGwCc8IcoyAOt9/N5yrVpH3YGjx7BsbubBABifNk50
j5a+z3hI/VDzUeV5dSqz/dbdPun+DljDR5bYFdiXy+JgDgyW7KYN1LxE9jq+ZAye
Xd3O3oryLdbF6DyekzpsuiGKAPMM94ExwGWWEUVq/xiRF5J+GI8nr5dIo+sjaSAY
YctliAtRBfkBR6AuOTvFOcmGaPJKBO+d78MYK505UuLFK5ALU6dOxdqh0yd2932T
xgNop9eXbagsDBvk4mvalbXVPyCtVwF5+iipn6DmUi/oYjYOir/UB5P4deOcrZt1
okqeAT+QuBBmZj7sM0+IR060g2p5D83wbZhWGqwL9FPh2+DkBKCGozwa0SJFL7mx
3f1BidYNZJ78dmUG9TbjqdE4LZrn2fDo0lpu5vQftswPXAvkb7g5FiuMsTZ7sRis
YEuOQfYqSx7+srALvRfjWsQbQX0+f5sua2paT3/AGG79S/C+qJ1IhguJuBalHrTQ
qvf294TGWNYfSS9jiUZf64J1/1WHBZ3Qq0o5sfYdJgHjBRngel6Q1iRMf6yujwn0
0FqxZ2IsDZ/sOb6wLoyQ0WSwiJ6ZEcs61z60h+YbeU6QilqWweNyphFjFr1w06zV
rZdyK+eaQLE8dQdZoyZwxsmIZDjuHuC7EaV21/4oG4aPn2ImrIQOYU0fF7EwYmXF
9YvkSlD6vSSHrC8zlmOFC9DNBg52oX0wv6QGZ63Nkwwzkq81lEY9Wx4hLk3MNucS
psEyjZBxs6ufWva3j44gS6pkBSHnITajls9ObbxKUCRy/2x+d+dBiKbEGyvy+qbo
o2DxnNnsYrxq2ZpuK2YGHIaRmfECazuThPzSdFvq9p5d8V/osuhZ7oKUkk0t49Qo
elhRliYR0e3zAMh8Cz4S2v2hMu3bp/6qiIjBJVq09Mz56AGjPv7ARE7ss+pHFD/w
VFEBAlWkCau9vJJR6n/X74SkGoQVgmIMLlQAySchaQ4nXg5zqO3m3IWiHrMbsFdS
sKI8mKAbtUcpEisN1W9F7ILowx0oFLCAMRb+qxgKPpZ2FEZpPUA/PW417dUbXl55
trlgbBpP0baKGEzg0Hh6CsPG/5fO2w/AkrTuT0IMogl1ohHHLYY77eJBNjeJ6dH+
ufELZsoYvpBzwUj7RU9aR0ryG71fWFeBXMFWC61MzEXE3JutBeYhpuqsWRhWi3bh
9j7ioW70YA6SygyZwVfy2HCsYs5qvYEhPoer5Mny/e9Sf8iYdmzYDMYSNyQQaYBe
WCodCOL9xmwfJ4rxhjR52dM+KeTLKGW5YBFjuv+FV/mr7VHcv5ivtsvIrCjb4N26
go5WH4l5nJ17kfcWZPHoGXpQ3OD/KIo8hlJSz7DJDkGGmFCSQL8VGPE2NRG+lSRd
zBm18XKiNOiM5OyJ941wuZnPuIlhzJU9nwUz9rIMeQkpNs2+HNUZ8ZJGsM4cLHyg
0YDuYLENOY4YwLn/Cj9j+QEgXA6jfMQOYgSjG0Flrj6FNxJjavXouxc4ID7i1f8o
Kgr8vpuMHmmCo8QFLlzd+2AbLbR7yJTnpD2lC7EOkrWm51+u17qNOjSnnArq4Th5
krV/7eP1mYWryEq9Lh6VE+tyk45XfHqGPUbZX8HawYMJS9FaPoEGkxKTMdoWDLm4
gPw3S5a0GQsoEtiulrRk6YjKVpIUvXJi3NCxfLvz6zSlGo5Ew92w7Ol1Daub9HmE
UA0BLuqHXkSFgHTKlykRcXsBvSbWG1N41jnodWbntCTor/L+rOuudtI/pEf+YU3F
Z9LmeGP9WRu8Yy+fHF/RVnzHkSp7lpQxal8JYjpeHvQzlQv2Z8c7z2KAUNwcmteM
4kovES0JFGpuIwmqfqMOsQtce03lCQq5LkFoOOXocu3BGIMOgpwAx5gJu3+8rOLp
/bVV+ESb/Jx+2uMLifNiUeAMFilk02kvC6tlN6DpXM+sFMl0sKPdkIxFnu8UgDq5
a23iTewgg6Z5L/0/CSC/PHcz3VeKAmYY1qy4kNl3yvAZ26pRVVTBIX7YU2KPmXkk
kEue3EUHBkIsF1jih5YGOQwVP2Q3trHJz24yrN9nl247CaJgq5QUq6/451Pbkneb
xYqI06FHNxMtSFwjUprzHY6+nAmtJBdC8bn1UWzE1xxY/Z1H/cW7mZteulO+hgbx
B9WSttMqYzAww/Jafpmz0Kko1b1v1/VrsZ7BTInVMSDZOV50Wy5ryPZhYRfZQYwM
dZ+gh7voMxLxp3qSBotALuWEbrqF1z462uwnYOTGyEFPr/pxwrR9DvX2K3Td1WDS
5gC38oLqnY94hEc6Ua9inWjjULSgsaFtGBm3P7wq0z2DGcy3qbOwKafPVUyuar8O
XsR7efnw9eUNVfXkwlNU5441v/NVS/wS146sn1BuH7AECpQr/h/uSMxaL4SLdfTm
h+1QejC9dcKqM5xmxvN6NezOdQMsF3AJ75pj+nyIhJzqh97NbU2RmEuS5ESnO44k
bnF8tzQx3gMdm93y/oKtMyVzy45WGmrbuguvodZDpxjeGYk3tIwxDIwd1XF18Rtr
pu+fBXnn4jYuXg2CLvYAViOKdItFiXG5rIxEZoW8PEnKDEDyrSJSczFI4BPz2U06
XlWPlSzQYYZklR8pdTe+mCExnVoun9j7MAOHGJGLCt9Yx1wIfRG1A0V18RHlLVTZ
6W153BlbbjmhzVlGqbScsD2SsIhEoIn2egNvTEZX8XLsLzTzDxQsYgrRjhz0PKIM
WogN+wClNVqj9xgcyaRDkUNvfzl8Lut/3KMcJgfrCUq7BoBw1y80Re8NQHXuh++y
I72fxM+gEk4zJNztKBd/Kr0Nj60lmCpNO7MFRCwyKY31oaVujeEY+nBNYdFqpPO/
DHYXTWSy+O8STL8evlK28jI2aghqXj50D8sxrOcsJt3BxKFqi8iPmSMEEY4Jn8+j
cPk8+B0C9azYt3jVp9KjSKBNRniZSO/Tm9omTqHTmdrxLrZLaGFwya37AeAHoyGq
yhSJB0KEOesJ/FTNY3FSlbDRyGQvweFApsjMDlYRybGraoZSfXREAevtC69Kg7wR
FaChWkqMGX9U6i9ggO1JXmzNAoZsYBu/gVv3FjJBznpFxPNIe2v+njnYn6ysCN/B
O3SijaKTJMlF2BwETYKa/4sb1k2BYV4HlTreXBfEl32fkiEvOvkcG3tWjkq+68aq
Ycue8URRwnDliTD07PWKHB7Vg+Opl+xFZ6V5+Brytn3UUy3TvfgwpvfWYkYitAXa
t54BR/FPsW8QtL524NrAvBs7AFd4fkyZ2pYrNSkJ9LRhSHigAnDx5i0G6jGUzcnx
756lHKlHs3cNcnc3GF+aBfNNTEUlonAPcbZQP1ZM/Z8NFmOC3XXLhh3kpim8sbGO
/NImCDy3XQZG6hL8+3XSygjBG3f7ftwb8JCWOG24e4gKJOvMjPecynagwg15Cyxt
DaDEvONqUmX+VUsHiYgWzJWPYZ9/nzusn6n62clTokibUOIMQTmX05P7tUsFghCL
ySsuaL/iZ73vm/PrAHJZP2H5FAj1F85AmVgaQpWsUkM0E+tlN2fLyg4atT9iKbv0
OUgOGluCW+oElUKcIw4J9tGeNxtYOG8MDIftNOGQkw2ujBr5LWnbX6tP2ZCRLXMc
BR85rru9oud/jj3Ak0jMyPIHKp/tMX3NlOackqvjHEyroOhF15BbXeR+nrggwcRH
bpv3F2kAlNFGuf+1bhWKE53W0WCSWmowvKfPm5xrWy9SSeOEuqW04mAbypGyekkv
NaDBdgCq8I/pdMVFf46/vkErqkmJrUn8p+xvZrlEuGGbXOSFAz8ODE4nuShmBnsn
YjeygK8dJ8piV/1kb2DbPA3xjOJQiLGfYJkO1YzMHHMPMjcylrPxn6rV139fbzd9
phPanpIFHZBGNms5Pm/Xjl3XQMCdsPpVyYNYlQNWGUYmaKqmzNvVqRqTvxxUY3H3
7jszZAHh5sBW91Tl3ROAOlOwVdlkSk7iOHR/zSCYnwQ8Pr13j1NuOZPHwmagtah+
cBwGo48LxHheZhhKhDy4ByZF1TV7r1+FSDF3Y44F8xgAG8zpt5bznGQLYEkmH3y6
Nf3wQgJrKVdkipgxbsoNw4osGeiGSAzpYHIV1vga8prt388Lc4+ayWN7/3HMvEdn
OyWPYj33aC1n20X9aI2Y7/as4xCaotb6xAB/EY4i2BLL+QUjCaFCd5JAHZYA1MK2
x9nYEEY6tP+uLKChjf3Xg0meC/vsuacUJfWxmJrbezABCIkjSwh6AGplN3UU6uKP
dXBasuTfK6UZSTVWYInYRdLMP3DdaaewFGVm0ZyT+2tSdDcFhq8KydfvNqeE2Cb4
UF1bOEzDy4oc6wdPYVbXtwNEoHHmjPDZcavGIyYMexVeB2Bk36gqLjUbk/pMz1yg
Vs9Hau0xtBeZ0lSGQ39l/z8vHmMaSOnjBiIcfYmLqglYg2M52fp/mZdq46zodM4D
rot7pM6Sa6i9AZ+G3GMRcIoma+0ZOIXrbw2BpYcWnqElxCIwnc9Cf+ewzPp55Ds4
BQUXpiA6QN67CsqlU6fVe+1DYGi4gxPJoWRaYm+2QXJBYWyQes73qAs+lt+katEg
KMKd2OJjXTIiPBIUGcoV5sPnPxcXvJFjSBXucROIamqgRseOIUckyuJsikHjlTgX
donIN37+wZaejYZGt/zIING1N+8XlS1P0BnV8GtwW/tZ+B6IR5IqtpF7e89V2yud
VpJYUVu/nm/s07sVIpZbOZk4utl8rsx9V/iDvXcHtbPttkWfWkc7pFTehZIo6MbW
YtDIZ19ReN7QWWmACTwfgwAGeXIde4Mvehsa9WYCSt5T16cKrmf345TkkfQiTsrZ
W14kUTSw9Kx0uwHRY5bh6VIoNaK9ver6Yt4wCglACNxSK16iI101tNEnL3foKM5B
lmQQw3UnGjlsUPmWOmdcgXCuGmU8ICwxfkyXeSptHnpEsNYe7fs8svsj6lwbnsG7
4JAbGcMgNfHkEw2G4L/4eoHQQmGtfxyaMMNirHfowfAWyOO609DrX2dmYaug0lad
0s0RKR0FeYoxASiIjTdz2n/KfX+eoUHKMDmhGcdarO+YjgB0Kh4KhsVBYkIbPMYA
8d1dCN2fAvtwm0RlU57mL6BeWXGS8OF813LSPh121gVxVDPKOWHcB61ZM5BkdDda
C6/hAQMUO1D6Q90iNfCQ4FnlZK5+4lRIWszbZKTe3z1YYb6QLrYFKjeBPjR7E7aQ
A1rnWpKvJXsLJx5HWzqcjRT2RuySBH6Rmv3HiX93/Kr77vfbR3iRsdwDKi/ef7RE
hcTQTmq9fWzND+/R6twpOq2Cft+DoZx11cLLoCDz+uWr/UiYW80/Hj9LgCPTT+YU
RPSyfmcOfPrb572Fcyvd7eHCAA2b+98ub35UI5VTKmGdp9bFY7yND3ouwq/JDaJ7
vQvP5Sgx61kBhMPQ8FBG9rMkFhE3ngdzZkqc74aiIRgj4h6Q2CT0El8DXFHfPu6d
uKuMEjssGyP7xG2ZPShZRFROn0Tq5cgvVcgbbK9AkQTW7SxDkc9St9gSpYhEayIc
TvDF8H0OZRudc3o5WVePKhKV33MVjhPmL7Km44m1rT5zrzwJqxiA5uHcdxqI7O3z
l1efPStnopYQLgwJYZZUuD+G1AzQESxnw3kPZ5HrQ3PzJscn0BMGA6hldrJbzwq5
r3s5+NqwK7Gs3v88A0w0y+r1x6nm34R0TkLrGEKcrc03XiPoQSk3XbvMMuD4j0zd
Y04Otyc849h8lGR5ruif0rQg+Uz/1zvUI8fEstvZw7lXat6aKt+RY5TniM2vrrs4
KAgornRTpbFfwULVFfK8wTW9OJ8daoPJCsoOtbSBkY8P0I2sDHBGs73v5BCpi0qW
JgsJ10KD2v5Z16W9/B55JcuQu1WfJM9ATUTxDNQ8+sPlERVeBqE1Ke76IzYOymFw
QCx64kAamV9jf8XstBY4hu8mmJn9nEcozJtNFsRqlZ/2UkflpnRLIGropYwNJvax
lVnvpKE93tJvq8LE0nlXJV0L0GrJLVSjDCgv/hSdO/eUoeO6b5funHA9kjsDthg9
fvU1a6REHlyzVHr2GXQDKrhLJDuh04mzTgZrVZ9ZnGW8TahkBVENN5NIY8OajoZG
I1eRBEy08LnXid0ugpmglcgnuUaMVjGPUaEtHlXX8OabNv5z0MM3QY+ECznrZu3d
7OYxsavaWXMDlfBAJwltmQEc8sYty/UzE9zZQmlG5mE5ClwZCM61VEbtt8N/jPQA
rBnW6IhxDd1EMRyMMIxxNQDC2YyeklWQTkCv0tp6o0i632Ho6m1QKLyPThBsvk+A
FqA1JHunYNFmcKDaR9XNxhefwYovbqOHRP6S8yaXmWXgkOR9FEI/xngEc3zv4F4z
hAlcEeCDUegwZ0MlOr539WQIkaLiHFhTu0oHm6/F2YlKRz2hPpLA/6fG4nDDxAQ4
kyyTdcB4bWNxDN/r0xnwP83DneEh5JT35fMcKgjl8AF0ABf3zPST8hAsQyDP0/oZ
28+XOLIAmsbvxvp+lBxOu8Ye+j82Ubw94uQjW4NVmgiTGsyGVvjLXG01SY1UDSTE
Z+t8rwE38Vs5xe/c2KPBLmeFQwEFkAuQuC4MkHXylVaMuIf3P65sOU8CuFY2Bkox
mFm5JzYmuDQC/pwkxpNM+kJuQxJ9hUXx4yJ0+UIcG3l2PJQ64eInBm8N8bZzuGRq
qunBQjx6WezijSLKzreaL3XtsTwqUZw5IDt8EYld9xyZywOaspRjpQw/xPBetML4
QN/hqbSSTG8HOZylkPOBMggu16E/tHCaGOJGtJ4weZSJZxaGLhpi849GSz7+fszc
9RqyMYoc8PfFXNayBun0TGx8JpoG3Eth0FTRri+SbdS62/cPM/x5Fm7Lp6PAn3E8
DbGQ1ecFOrFf8OiMoGC7JrKcG3L8TT64z6t2sg8hPL9WmipNdhGW7vayTIlU1vWo
0Mt+a3UPzSDhsDIaqAuDiIeuv3lMKiJrYjiPavGsVPwsu2Jj7FW8P66lzL0hwGvt
yRSqbW8mSP85YEb9cSJXG9MKVl6tOzg6sPWJep9hrb7XbM017bOKc2YRZES45lWp
aZQOsjzaJA0At4NmZCRbb23lcHJs8EExvGtgBwYizo1S/2u8MOnKIKc5TsZ9Syhg
wHZV6la0sHX6fxxAhAxdj0FjNq+jeAWSPvWnD7e3ObYdbkZhzEAo4vStwXpDGTD1
STDi0FJBkCl8u6jtnmJJ9lIaAfjdmmcA1XU+3HmUDQRcpdXnmqV+fj2v++joERHv
2PkZAkVn+GG1ox4YKQMrl4WbAfnC7e8edZ3kGU4KZ8RvBOhr2VYsWOrzpsc+rfPj
dpVD46GCixvv0VNhtH+4E8XH4HAwwLm8t4j2UfMatYjQHK8uOsLiaMCdD0CRF7rA
SCOsjQbDMGSukOpYEMeKfKp3SRc1TWa4j27YkAmadiqYi09/zyqCn/+SkRsx1JbY
Tnb25NNVhn7lBDhIZrXJYwYI1EPhb52gOQdkPR0MjrjQG2BNRwfm8Wyj44REldXj
Kei3iE2s9gjGgA5qyL9pAIeZhzBEdjencJ7tFlrVkQx4hKWKNXvPLFeveRKfJ6us
i1XScAJ2qb0RXUczzmGc64KFWm34n5tpjuPaDtsJY00Ionzj7ZmVxqvA808wVP8g
W4O1GnM9vVgp57tdTJwF08TOx/IgCjQyhWu6CQRjBG5zdvxajUFpCwwYHAAqtGGQ
FQkGSnpouSPQFfLqZsSJ2CiwcikEYMExqJN7tG5rZ+q0ioB5OEmqJGZRuVTZu/li
/UR4Ja+64OiiSuzNc8I1r6/v9zsNPXgrZ32czBRaAYH2Wg0+x5bPE+tmxmbYQpgw
vSEN8qHbM37837WF8t1IIlBexN9kxbq3qgckJZSUMNega0p+HLQgUyVafVSGjeNB
ZQp/USvlEj3BrgGbYkMieCdGLzC+PdRPNuLMC/Ipgl1uiRDKWntrVCDW9fGdpSai
Z/rkrhMAUhxg/PBNjdQcW47JoTLlnsEDwy+q/sohvq2rJvQQsdYtZ6LtuD41Zb31
q49vmPH56BWUU/h3h4Z+ldnjiWFIj4jTVMaCLt/WVZfZRTWdhvw6j8zFDGEu77RD
oRWqtfYNF/8czjRy1iLIQjM/3zKoruxGXDuZHCXP+h8FatjH1W0JpsQOcMXGrKF3
FJdxKW9UoOOvEMAyJ5QAE47QzC0DvZKtWw0+v6FVoaIUxyv9F5MuWDCLst0732lm
WavyoSwaOdGS9R5A2Rnisy8jhNad4e228qFhUX77aAiO4anuTreHOtksEobvOTqT
SZtwIR69mMLJRnELa3QGFPEZhbYhvJD8AqKAnJ3xA0GOaRVooMH/auyPBaCQpy+f
w+vVaQaWILI3nHURXxQOgxcXpI5h/omLwBHwmGitWG4VhsdOzydqkRTdlNODWeJe
OSgM4HtfU8+R2WcxpYhfIQ8q2+/dSh1WJoGMIOJl3gEMLVGtQ3SyXIZj4ELxHbzx
AgX6EPojq0xuTTnzpSq3/ogCc25ZJsUQX4RXtTjwXZwWok40DJB3Jgu8S2V6/KJl
rK+r1IG1E5SvEoy0AtEI/XfBCgpXHiQKhcYf1G5pVojCKb0XNB5ZmCNTtWO0Cp3v
F7T5FtaoUq61AErh48TxgF/OvlwRH1R1G62QKdaVuhjhcd2oJZWHM2cHoSUdMLZR
gtQOUPRnAAjSdAF4d4AQrwdus9S2WZ4nUEB8R2WaViKDDLtAPK04vkH/UKbWzR8u
KlizMrtpknhYOBXeb//VTQIVNysyqCTFS3vWNEQMfMamqX0ph608fv4ShicgLwJ9
60wveEnYDvtWQeVHM1MncGS/ZLBloc0Xs7X57vZSxKjgVhW3dR6EQPpYvbBV0z4k
orvBJIB3J9e3SJywqUBK1RyMZ8d9CAzRAm4D57qSwwVacQWIHw1gu2CKD1asSIAQ
Ee2kw55UdUbcRhHi9vRkiaqHbO7jHgJNiijz+tFQBuGFIMr3o9mc8hSp5anGGBUO
tcaRW6/wbxFfUw3TF/ovr21979CfEn6xS6X/wcIDp/V5AJL+CIjO/skzhlNCJtcj
FlcIOy2Rz8yxfQU+DXqmHOb0leZdjjILBOQo3tzhdzNM4utNeS56ahxvPNrt/lBB
nzaMApcjXSf6KcF8x7MoBzzhwaCpydoktTy67dvSZ+7yXY7p5m8e3e4+7sarLp7O
dmkcr4DRu5DqzqY/DT/ORqtHgmKJU7vOjaea298NP22Eh2ZMbphuTBXdLwXqwvKi
8mbF/CuF6ViWj1XZKUTShrIc9GfNW2TBiESS34oSp50mYdgY+yMftps2ydpXYo4C
5CUCllZJ/rrnUUf7NhtpUhz9s8FxmiEa7myIVggiBmA2ZaN0FmUSLVF/6v7t1JDd
BTi7xWUlvFYU7/KQvzWfhsG3gFFGTKlQ7cnzCc9WNIlXBTakZlNDoMN3AF3/thmC
u07036YAi8Os7UuZGvvxgymWlhdY1yLABmIqGYC19JB7aJEMby6T0ocIbJUgiBAC
uPabcWag/UmMwJ3l0/yKSF5KUdTqXiNRPqieK8Ev1A2qqI3OUqAPw26NNuil9MRx
ukXwr6vmYyde6Y90OKAtOvkxVFk3Z7fPOX1oiKyiilYkU4eJx0FHzP3fYJdbu2kY
/2LRPKJ+INT6a/oR3+QC2pXTNuC7T2RaCtO/0yzS3HKmLBcno8ID8/vlCISos4Vp
a+suQ9qXCYeRhXqXt5llhBFTxA8Io8eBTCyivCLq/uV4DDDy4tOLgtq5+QDWoxQ7
s8bExfR4d4sPz9uuAYe6shhwpmctG+Gtu0IIwZWlMN419nLfEwavTzRNeHYXYeTI
X/oTQEHHCrpPfzTHTtcK4Q+BrhTa8UGbzpn6Fd2uyM7Vdk/2sJuxFuDGkRBEj36A
2YKSxgzV44canYB7hLdEiG/XsqrTr0EPLpkOuRqbHfmXl+C85oIY5wOVgSc6Vxww
PxN+UGKu7Ehzl37Q3tY6QH5uI+CXUm/Yf/mp7UuSq+Ndn/pLSkk70/6AGseCmWTV
Miwru7uRAR0xFicmw6AqANr47t9j78Qtrq8iopMigKlztSIUKJfrOK4DJHel6Mhq
iGjznThqiuV76sdQ7zuKREj48D8gaHqeHT4Q3a4/p65j2eU+uVaHq0FX5vU5nrcF
o4EKSbHcqgWIn/oPv+tlQlQ0tkP7ecf4vDl9c3Y/LhhuL8Yyz+6HbYHBZ1JHLqDc
Soi41TsQdV4dU73+r7ebBqXNQ85VnXeNZfUlm1R8pVqNTFoerorhK3eTDKJAte6u
3MrT5A7qHe2DlYucFWN0Hj9vOHRzRip5JoZBhqCA1AnovTCtUIdpUXmSJ7Gp70uF
oeMr87pPiUsB68k6C86QZsXQ4/BDWrDL7gO8lmBXp8hB3293w91ssCW0x1qjuhhy
ZNuLpFYiYp5AieQagZibPLdWf6nTKjn1xLYy2/0NvVVsCJBetTrA2hSaQl5MCi31
zw/yyLDblkqegS2E47d5wW50mJrxx0D2lAW1FIx1C5dn52Pz84Ka0I/xfNyu508y
SjFq58+c9TVNvo8syMiz7JzkKlU6MfwhG2q3ZxGU9L2iFG3n0DeK/biMclwuqiJG
DnsygtSxEuZIS6oxkJoIsjguvaSwRjTx13mlxB+2zDxq7NpoFmhIYQprf7DfVIgl
o/AbTmjcNe4S9bTCJfvMDH1HYvYuFQufJlEakMjmmc8ceqluQ3BjLROmJSa9HRiM
rtLAZZyZ6IO++A7eI1hct/HWA+S9mgXgDbzmxIgKF7DFYcBhvwq5uPeoNbVD4ek3
8OSWPdWr38c2bTJjrlXfROzDQqS2buF5WXJzlyFuHu+KgUGvfMH3YTJJ3l+Y00CD
4xS6OzegVcaqtrPXFkhpQU0obe5AeQi/vD/y3eZAybb59kUBxCbC3Ox6VVl2lU88
2oxpPyRXaJzD4ck8/FZUYi8iF9zxhtnkRPbn4SMSGqME6YI3PhBSkaT1ImVGrxJz
nzqp1W9TeA0zPbwH95akES3q0DuXaBzH4TvugeMPZkKGjpThHfbSAOnQMgXXb0jR
p3ZRBfz672WMy+9zGJSxH0aJ/J7eEZnGp/0WS2rUayM0PEBjY2gCp+1HOe+WHAW1
sH5z1i2wDiLvJKt7YM9Z221codanbaup6aH2wRmkKxCzGWAg3L6f+kIt5+GTYU8E
p7GWLC4oR1QR8vY3kPjCLq6/YOC7rU7hGONRTKDWRtEtITMaldgE5pX5H/yl0WNG
uWcwj5mD81/hAWAt/soCOhWVMUwMChT0iW2SQ/24BUlul3PJCqe0i1sUqZXp5By2
ZsnMH3YLVS3g6+hfskdy4oOud7VoZNheJz5fNMaDtN3HF/CgTW8s1y7CKYJIn3yc
F5kB6+BRchloxdL7YJjrH1Tn2H1Yo73IgRpt8JuHHkAoElRJTEdF193Qfq535B0r
bPPthgePK3J6pjDZ2g7lzs5yFPyLQ5uQmY/WHiiJ+qDrZdQsZ2W1FTHjKkg2dNZr
KFZilM4WXUKRSuiUAtuviB4PiwvnqXGB3BUMc0E398tmdYS9q5Y7Ee1rysyKGVFW
gHpuVj/4yOUFZwhT7VtXbTGLF7D/v4gDoN0kKTm5DVU7/gJqssM7jSUhatDxga0O
Dky+xdtSsbqwljRAStgeUxrO+qzUFFN0QMhk92tHoQRZoJmruofv1ioEpBdPSfSt
yITLDMmD4pgX0LQ/6TXvZzlrLLLdPw7l5scUl5PI1RovntOmJUzpe3EDpOh6i7T+
MEKLDMtkW1Y/7M9gmhT1QUd/knJEU53+K6SGPTqFLVCozeLGIiOvEkTWmdw3Vw5v
yBVJ7pHjYA6E6wSNYzwUXoy4FSaO5FRcdm0mssSprlYN/O5XBZu95+qxgXCtmb76
VtePf8MORO43/r6ZwUBTQGDVl7oUoRXW8M+vxjdcveNyBwD5N2KfWSR1x1BkNHmA
Jnm9e4zUburg26B/IS6+wmLdd6gtwprck4sIyj1tVPCtuzQcE1PeHbEED6psXEd6
E3Dji1a+xOEWEdlcAcij6Dc6cW/PEPBWHDISeXzLmIDBK8FbkgiG6+Mg36he3SyG
S5wc+B9bfIQaA1md9nyOZ+uAmI8+ra0Avhiwjzsog3cyxN/9LN7+sHY/y2tpxKTn
IsS8Ce+hCuRJuJJUjMtQfht89K7lZMF6Rk5+HYFyANBPAsMGKe20qZDmsCTmB0G4
5FhBqIc6sD4kZ9MZWvi2XxJz0CZ5yACH8l/f9Eno07gY3tosrlqm86OSFg0xldre
VUPxjM175MrrTYs6Y1bDzP7jl7VNwfIbDeUhSnPqrHivQMpIAErjaXsWlYLGYQPy
c8OaabnyIjUt7sHBAHXTI2rV8ymj/JrMHPiIr11Si5qtFH6ZvvlCqLaFkq/nKM0z
O90vuuea4S7IbKtLR+j6KXVmRHTWeICWu7a9+OXjcX2vO1DyH3/80fsYYqtnTQL9
0eTwYD8xzIiX+wgUHvrgiAURCNVxQ599n5liCzLVU9G5+XCmYlTX3DtoBYnicXr/
2JXIujDWMZXheU1keVkRmW9x+zJObp57jpIP7bshoHGMNQvpewtoamSZSRIj9mkq
Zyikm9pQIt1+d3/ZkWp6IO7cWHQiuwo9WVHlVkU+/ZEzD39hiYK9+TUxZSfBdZ9r
2+0cSbNDnc6cvwgP3aMjA/D0KiREemueiAbVRTC2HAE88lg67vNTsmxk1yLbnSfY
pcFfqT7ttKxfo7cgqVi7AgwOdRiT/e4Qu++BfKFyS7ArvaOIz/rTdqGDyb8r190D
pix2rakMF9DQpRwfPSJOgY7P/fXCKY0tKAx1VBMWTqkv8HvIphZrCrsiDS4mL7dV
V2q65qwfBGCSiDrZFOFElOJ+349atxwCj/Fqy5u6u6ViijgLdDh/Jf8GJ+Uibi9u
fLDuHYPgz7Oj9nS6jS2RzOHFpU5rrVsaAIiLYCEyoDMY67RGiiWnqhAWKXcIP7yu
FVcRHfGd7EuF9HpBIsN+2TZl3bk2zCn6MEQiE6oZHx7lNA1MaP3NIxZnSsTZtzIk
V+FD/X2Vb2jMj6ek9735K+lluvxo7t1hwQYDLFjeuqqIXwtXwSrkcVLSrBuMcdG9
OmdulOvxZI4covzn9fWNfSLH6CH5GP07X17lRAHh+5s3p2wPhxfMgkvBVOfJ5mKp
eaF1dlZ62muQjxUA++6+BDAcz5ycNyQP98PdGP32dXRmDozgbI+KWP9A7XoRwLXd
hnJhQYl3zm9DqKDxWzfMJpmXA/bpvtDnc7xRfEEyLwcubqAtx3CXVM4SzJco2pbk
Q01dwAGcRKz5P4ta9XjCPC4wY8vSG3ZXm2ADYr/K71jM5JMxnbxqCPquSkmcdhjj
G+bcCdDyXVeFZt3UmvOqPHGF9I55I/dNAl03IfotjxVTyefkVoxXjwmKuYlPor1W
mM+np88S4vXW/HFOsfPuEvm45EdvM1ogtVmT1EAJZx7iX3escyexY1kY3OUG1XzK
7xLbPXlFrQcxUDP4DQgKPO3kM+7TN3xhTquREX91A5TWekYmqAwN3FGHnhUDboNv
7Ge8871kjh2xItNXzLGlkvvIMX8UnFTjr/WJI3NK2aW+BhF+FLEFifdOhrOEaQFD
HRDNcb3WLRFCqEQsvzcowL3SKHz6mRHsJ1Iq7smpYeTkYhhGybyVzrX8xPq4omZ4
+W8C6rNsGE0QYhhFj2nct0hhoYVa3vpIOHXN27aqiW24wlqdzzVJxkZmjkGHT0qd
tyZy3+ES4qveREz1lkMHBczpimnKnqE25mo19lecjmHd4lbsnn5n9gDZlp2ZrfRL
aPOMxHKigB5iae+attQ3O6V8Y/yN49cpFtuaSuCFBkl+1ZeqE3XIfPHdhrbUmzdk
k+RXupaY6ey6IAcX/qGhGRisCZVRD/lKunQCEZ2WdnkBXFW5jxijPUJ+sFuw1YFL
8W+C1J4GoUMtdKvWCzFL9WL6lBUMzbSZ6Te+HpGl/0ePTkExEmgRr0dwHYbnSknr
WfqdQbx1fOFCp9k6c1RJ8Uh1lnFHOIIzkbbjPJ38ajFc+WYsAPG6g3EPPlFe4I1c
Z06hQB9/g7ZTJhoalffP3Kn12QlMhmENY95g5c18FE2cSGAPE8Fs6qtC8E4nJGrm
/aCVWG6nzXKCqdMDOGbfl6HEV/xZ5dx4nN9Jcs52jI/7r86T//jbDiFKEPlUIy/C
i3XnwuXJTu+O0SItH88sKbEBlRT8Xx6+8vaOE+SduEbf85e010Uyl5S1/19n2/7E
`pragma protect end_protected
endfunction: pre_randomize
// -----------------------------------------------------------------------------
function void svt_axi_transaction::post_randomize ();
  int log_base_2_total_bytes;
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
aqU/cwvPFd8Hfp5tpd+dpwnkAVbqVB7vA1tF24Jak5ap6P+GGul1wSFW6w7orDCb
rKv3/KPRrjtepN2u75rUD3oLWzv+B0zXQKTGENk6PPbJVCVmLccUhtr5zc/6eR3/
PilfZQAx4j2X3uBEIFIazq+k16fZeduc1OGEtT5aQgw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 25838     )
7Yg72BF1FbMtqnAwoNIoFAHVMYM9GugRMcJWCU/lMEVQUjeQhNcklehNlC8LBBA6
fVEGPMt4x12KbUJC8ondUCJdXKFdmQxOJRxqrEUcD2nvn6+IwJIZ/t0Isc4jemG9
afST8Lp/L4UN5e0GLim5oHmdEgft4HZmuK7AQfUeeJnzP3+0GNFJGbimLrMk3ZzD
qqJWpFzqAK3M/pAYNjEBTrlfzc+4XrrLeWYk1LsuDHeXSjecyV2hjgdQW92xxp+A
v1KdNz9z4uFmBs/7i5qKmwVqsJmbfIePVqRnb5fQeQFoYIyRnlANoFY34D5We2Qf
QQ2P6Di8mLaG9fUvorRWas8ui9GOIpEAE6b1PwjVHKo8A2GqTUsuH2l2X7Falrp2
eXZKrqZVS5HYRnDkIBvqZg1JykNVLJRR8qb3ESoyb54ab+7PnAAXrhu+Sz1y757D
f7PaP+D4Zc5/p/6ojTTX0EkTdjrgEmN7TVjREB4H7E5bWUci0WKak3x+eK+gHAnU
8g92JMwQ9WJUwjDof7MpA8XjNmZZ88DL+1EFcGO04ktNCi4sx5cqBwHZfEGLOgRT
906kCiG19Y/lnQ0TXRYTwCw25ukA5sjVD0fdvDRTvBIVK7p2pXb/uegVuOUDSPbK
KazJmT83PmNpG644MBwTcRG/+Ie7my9IQXXycI6p3Gd+VQod9MOwjOf2wkodoz+K
R34l/oOb+iC30Ht9RMZA94sgj+U2vT9ODi0FbGsQxU1RX2n+KwOIgj52L2jaJ5M2
j48LKVpfNNkjl9vYstXr0beroBdDuw4XWa20ro4fqFCNU5QVCjVjF0EQFC7NeZ9Q
+Sm6Zrwu5KKMHL0nBstICeuDmvWVKIWilUjfgqrKOGqD3BsmIn/muDYXsz1XJBKa
5RAznA81ZdUmxHRjqIpFvAFMBzGJuh3qFgevuESpa6J/zSmudbsK/AQPACVMNYHp
hP1t8Mo08Yh+BfzDsk+HEHG+4xVUxaKHNxfS4Jg87Wr+XFrn35Y7jPTfaaLXWmxd
8oFaV1L4LEk+bt9TxOKnpOsC5Uj/1we95y6X5JJ6rc5POaoz79tuo0VKGuAJ8zvK
7PzFgKGaL+p4vjvZ5zcpLAt2mwaebthgXOjZVB1xai3nCz7itBeUB43S3PNLaoLT
5rgwhkDlLjNHZLvD7LsdaCDce0uJDTVGQTWD3WUhBeAPUu1UUFw9bu7aXZlNFDnN
MjBRV7jNj0LSgMv1PtgpfobiaWcqOeDKQlt8zy16gXcQ+4Z5Rakq0VYMbvYUYtZq
8UKYI1tRPOWAu7fGVH+EXXP+clDvk+BEGWMKLPAtyT88/sIseUoQyOciwozjzuED
ii4yShBDkgwEAw5tMWOnxhowcU2a3XUY3ipL86cZM80YTm7Mf7HcrCQtPea6TS9e
PmHYw6JnaRci4evDSIec2KqEAYjTx3Ydz/LLf+ta/am8Uj1I3KW3WClgFSnFUrYn
vRy1/trUbUy66EgVHcNn52rfutyrQBHn+PZ8gKYFZVdCXegTdK+S+qBBo+oz1ZGr
5ZgypvuU4w0oc6gsxSlLCgfLjfo31MXZHIt28KoC19WHxxQ5TDisdAvkbXI9yX0T
JJRqVz5XQRs7ZH8ez/f6wexAoBBNaxTXnKnPKa+CLMsntlDkCMVg44couBX8C0Ch
Vnhd9lDCDGXCc3K0bEwX8mfc+jLCwz1EJDQepSjmyXnXck/Io1aQf9XiAe7SorV5
j4kDvetWQEj/QpmRufIA2Uw02zI4WwcpG5XdOBbdEMehpN3F27WlihGQ3M3YBVNk
Kvv6XOdpaXddciGfLkrhRDoqPfpXTlsn8MRT79c0wLNxHRq8NR2CLF1FRN+F1VWY
fErpfSRM7C+7bd417t9vUIfObQvJnZE7PVY1k87oVYh1ZfhCtEM3BlBRp1hwzOKK
y8jFhxY5yb2UpyWdMvPPL7JAs4Rw6r+0qw2kXll8tHFJ3J6H6CsQCyGytK9JLJGw
/+X0YiGmiGwJTwDT1dKfUZz8ihrcS1hUNhRxILvQmch0iMZyIoXLFvN6rAk9r3Xv
0qlRbdm9btOqQpebIv3SrXnqmY4TssstfaM8N8/QOP+5+zadYWN6kGQnVMK09k7F
7y3RccIVDsDOQb4Oko2/Wwfw6GHQHg6ITc4pi52p4o+cFBniRLAElCJ6oYOaY7id
598YDcthne3u+paJkDZgJwcpz1ZaLbmskRyRR4E2pj1n/Il/sVyYYn4zssevPXXB
SGftzRrU8B6zFzSVtGP4W478eaB7Z83nySdw1MK4eXdcpwtROQqlrJPPNV/F40NV
84xifjtvUWCekjkO6Meg9Ps7mOSqAkAKw+aY8y2id0cgNrIQCYCSZVUg2fUIV6Y6
wRVwkeClNpeICwhDAcd5zpRH+OhMRD/i5zD7S9V9ak1dZRM6dy1K9lSMGOOJbXMd
sdLwf/lXeWMzCsoZLY2Pzc8gDS7i2hXGmZC9Ei8QEqenl6JRAXkMHygmRVU9LDPR
ZQpDkPowsQ91dK2QGHmCbRqE4ToqAiY73k46IQwEebOF/nww8X4DrRuOLdW69OWZ
0N0w/9FlBDjujrRNo2ueePmxv209Z855M8Ou3vVTLhh5zmxTKLfDTX/SGY+OuSSS
tJ36jJ3nE7P/DDNM4LVZ54CAKy1sypWHl4GJzSNwqewpc4vSBf8XOz85XnY1egfv
5uTOjy5u6tGjLJDaNMiWlB1jt2Ep29EEmh/1egT9Z6dTPDn9hc/evIpuut5NgYxr
M5YhsAT+o/Hwrw9ueIbdJYk4umYMwotd3fsgGUQi8yLv2pzwSCZkNcpWixOt0rM4
Cm60RbAdXMxll2M5Pm+ug4Td57XW4hT/nUSuKm7CNQNE4nkJH0mgquk+I+BnaNN5
nCsworLQrzEOX1cDltLMjB7isWSQJQrHQqD4COip4mv8n1PGAgLK6sUyi6ARGxzg
rl+243J02XEHXkES459+/FEr6DtfbRwDRa6nLPUd3T6xTI12qr+93gU4sW7E9v//
jMM4nyL1uIy4DJUUo4b7cDTPPTxPEEr1SHim6oEe8fuCYEB4VZVwcIHQq5pKoqtf
vu+QESdxCwNs7eoAAP0VDKSMzmljmJLhFSksyGHtDT2HOZ46TPonD+o2A+PF9KPX
MbEeHUPcVx9skeSHVOntQo0/O9nZ3PaewSdEiEVryvTMiqHAl4eEHSNj/vIjc7Bp
ey3/6kb+dzuoFcr89hx6OmpFwe+aM5s+gYydQ4Sb0KW+JGryMwwtnyySy42qVDQ/
xvK042D4ptPokGmsRj9/chKHltB6s0veHDgmXKC5kRrVILEyVQvHcn2ikoAZM6Lt
xnxZa1vD31cbcRStUgiiw9/gSS/HF53Z0BMYUd0+GULZFI4J8J8njRajZYeFQMuh
1WbxITXI1ve40suBiA6G0Pz6d3TP2ZJKjuU+6h+A6etluou+5SDpNTn3gZ+oht/e
4MIfUy7oYVEW3cKKTna03ZI42alhVcVR8GNBFe3uSby9JJP3Zv7xFByfc2QuvtqY
YSvF49+Aq0/oOmR+5JNtEyibBC6lqdmvSFTRoY5xSvqql4HYIET8td3NWr/Jfp59
29BUUs9/uhJqlaOLvv78mkar53U/NLGV5iS13N/W88qx5NR29QCAgi6V5N4KXgR5
NWpI3JsfxdqC3R9phhzOEAjdhi69hJpRJWLzA2b/fdoQeGlJ7UrZ5yqNReXSf5UR
o/SDNt6/Np/CZi8p2tpCjdGJgN5zJA4i08TGiomrEnEckqOi1ATkBKZQ1RoZDgjh
z4llj0o4dM0zmLr0ADT8QwfR/d1xz/kQrLsHM7xr4peNNrcVMDKkNF8WN4npXlME
KLDPuvUjUVWcQ/I+6yRL+/VONFVXQ73fHCX4vkuySVz/wZSjwO0+F6IwQCdA9/2S
FCsJ7U8O4DNhj/7CbLPaTLPpIAPO2nUtrN5RWrUipSMUE5pc0Ja3umBwdixNdZpT
X05CZQiq1zKzbiHOl9jMRZ+bgf8jK4+eDlQ+UTsEufhfB30mRzgOlPFLTVpKmk9f
XOi1ocXVs6y5/fDokiqFe8ivEsxYSZ3v1vys6z5AR/uKw2mTJFobCafllOLz4FCG
894N0/sCa+JAK15cNMSEEleJHIJ19IIboMpGthrYHvRrbdMk3mH561FviesU3LEQ
o27dK5SO40KoBv1kBiF62vB/HooLIVP5mrQiED4mqdjYqbKoy+MvhhxsR9+9zUdv
CPxi+cN+oZPWUV8/CVxPm7Fdpz9PK/gVU7MQ//M++bpYCnz+37hHUwRSyy8apREG
4WzDlUiWR1LCD4SL/rxh/ru7h0X/kmEw8pVz+DrgSlus+CNnMfI8cJGXrVcagOnC
cVfxYeSQZD+m+5GyZJZuo2bFOEBr49q1OyhKN0dTZlstY5uccia3HKXmVq44Y6Bk
P1nyHNoLneHlmG5lShCBVgEdV7L2z0Sd9JdT0UOlRwy/OyjF4+YePXtK4dP/ywe0
sj3eZvSdxPYzYTYWTYKc4+6rH/KyjO902KCDTRn21lh+uZqUWU1h3L5Zm4ghUv/S
XAlxyJJkI1Pmb9eLoivL1BCV1sRfh9nisUjc50RgYb1/SJaj7agIDDZdwlWzJ811
fmuItnBoafFxieB4e39uU9GkhKkt7xnnZfPs99KY9GyFO4xK9iSt35N7q6AmDgHu
iymHB1DWRo3Hl8+vDYVyd+z68motDY1uyHuSoRkryA5B2XgYXloRQfJn7t1PM1BS
LfOQDzD1vJp4JuADBh8QxewFkzl2tXtu2jQMbu7s91Yjew5VkFWEifdVFJtVo5Ta
N0RJsvod0O4iKjJ7UYugZOsomADCPAkGUOFnf2nctseBZ8ScMz7d41JLE0Ssg9q/
MWrWf6qmfrBavEzIgbttjQCwv2uVjIAIITbWjrhru9KWbvsNyWz3EdxEcE1Dbab5
izpitvAehmsglpUXoKIF7TsoVzQKtE6q9DXIuxelryL4s9Sk4x8vsLHljohf8OWv
j99MwlsqZp8j8ANg87GqvjfPuT44Zr1kkyLt5Ys4HJFffIOn8+lTN8aVTFYbhrEg
QU1cGsAfs2pxn0WMnGRTOjuEaTiBoLPrYLZndyKDNEKGzvWaiNErOTTuw/xfeS3b
NB1jeMKhoZEuQNwCvqy59Aw7DTAyOnkk7w/An6/J0/FqAbDPWicgrcsPdymmAcpU
+w208SnfTa7qIaYDfvpuYSM4IK5xq4oAVoaM3L7LOzBv72uudMGkwqy/KuFXOSZ4
dIIofAxqyFlZraSlorWq+ftNvo11mnGbqrrRmDBkmlXpH6gL3OtrhIszOFXdBhZf
Vi+/213bDPDHZW5HNcDj2HL95JmXy7K5oHIBIE5zvGDjXP3jsZSJi7vUOwRRFl3K
uRq6Av/ulpQicLPB3ESiZF94C4BpHTPhxl1iOkivauB0ppRnxmdncRsZIDjgidWC
P33HmBxIhqWLrIRLxx4ROOhqG3D7v4HUCcNlZvyTic33YDzj4+Pz4RwUpKYP45hZ
dSVwR3uTSianG3LA48is+cqppJuyggEj49tfCsC7nzKM7KkP/RfjKqzSbFBMqbuR
W2eSSMPwDHz/cg9+EhCFoJsx2Z9l6Y2uAeIScfnrO4xa2mUtXY+jWfUNmfLOGe1t
uhKKjP/ZW1CdSzJdnrGZTTJsIAPShETDCVAGR6bzw28j8Y0mPVnq7DBIls+mAV/f
8GR7mX8YuWrQuH8Vj2HOg0DVWRRiqOKOL3yA+IoA7yrPs73eI+cdgOfZMn80lJe8
g5pyyLbPld6i/Dq66z9b2/L5nX59xl+5uzdeqbPMr28u0I+YQKuAOl8Kg7NC5Dlh
GZtTD3j5xsy4pVkbTqiJkkjZsWkOp3X/8IONZI9VHDgFNEAbFXPdSnHgSU0QUiyq
am85j/YUQBoJRQIcf4R/llaKr04f+aAtJW08TnLbyaZPP6OnnbZjyaSUo4q43nFv
OAIp2t9RSW7tXM5ps9WXs3O8DJgPZNXeMzKkqEh2qtYgjsMIv+KtVUYMMFodJH8B
iXVgQ48VCxiY40I8E+gJ/SGudVNXXDn4tl1AfQ5XTS8PeXZINm1yetpD3BSYhAKN
Trm/Q1kmVjvEReEbYiR22Dm95wBBgMiNhWSZengLSmhuXroVMDlgoXtV215xnl5b
Zq0GaU1A7QQTkFVgoYbYgMb4JbmTZxfNlB0aJRVX1ev8Srb2zTkOU/+Md/gmo2/z
xcV/LrxLzrv5jBOTA9XRhH61ByLQeo0yRTQYfP1jNI3y65FbhXTjr5wd3TmaCP1C
jL4Fof+unLYSyyFcyFwNd87XAM4mabZpAjZ3FqHvmLgS+bYRZ0++HQtsBkCiRoI1
hoRGBkb/WJkGj2TkkeZY9dJ5JVi/Ub83xShYpE6c2iHtPBTypLDK3qWfU5O1E1At
Nv/H/XK4tiMLK43Lj8o6TxgR7lHhceTQtmXmqBDKLe5MtZpJsnxRDrjW6VwSPuun
J9xnw6Kg7QAyNmWCH1E0L3O++UPaA7jaqiWVzjchLp+8pX5Tpni08UidkqdHIzqC
xJ9yoDEfK8RnNa5qteTAHgetBL496BVDoofpOPqLsfD/t3sabK904SNKf7q3peLK
u66AVzXFXJvWLytKNNhYIG1sZcylPpFOEwuKvcTX0I6nIyj8S46t3jO+SFQbGNNJ
8x+z85lru27JyqNJ28LU+Tr7U6XmPDWACeRNTKK9cpIntE+lF5d7O2jjESJjSoua
+HLDknFluHNq0H14q9ZqTDiyNhujbbBRqGdYpldUqRdHyTdUHC/pcu8GFENvqBTD
0LiG2fmxEtbjarfCteljPq3UZw4NWllLfJlD4HvLWbNnZciJw89/W+BWxn2VXJFp
setsSgcOEcYcb12laGqT2yTqYdrcBWdkzAPqgCFwwwemXdduDRA40k6t9/EQvNF5
nP4/YfdtnhtyIg12uZ7PVElDF2gu1trA2USzLr+wSEwUOqquJCN3BBms+bZP/tFX
0iPEzudfD1l3UY2RQkb4lDm/olxOVtjrPg7TnT3T6yyuslZuK1dVR23be1PGxXv1
p6nsKYsJp+x9k4NZ7dkUWKOLLOyjy0D6DO9wyJ/5Zhv4ZjV3HqrmfkeIe24iAp/q
g6WTJmUadUkgea1HfN0fqch1n4iY97RlhRNsekgZp4BQKV7IcHyYzAX6Z822aUco
OU8rhBvoFukqLqwK55RKKLxBJIhnJsIgTnkXV36/xPNQrMl1q6dd6Th0Ln3LfxFz
Brg1AzvKoJ76SpbuHhOgaZD59DwCUcD0f7CrxRtTPFAGA4Utio4j7HXI7FxyGakD
hBF2Qf9H4ETZuxSLB0h1+Aphu2laZeCOMRmfJe3VOSxW6S3DcATtkYZ4fAMJ477c
vmkpYHeClIep8h8kPoePUH7Tf76KR3xhvz/0MpH3eahrLUHx2/vXoIs3EKg9xkgw
IsafIm05rxV4uOm3wIVU5QKoOeTkZCnahq/r7M1IfRDkGNLyr3CMnKZBYdflAxeS
HmPOgAB0kec0citKPNn+J/y3ZGM8MvQKu0SB+3goIhpAGQnKSsNRjo6Ec6UBerUm
kk6ni9YJEv/JDH8NTGxqPmgJvnGv59i1NykLvyJJgwrn+TttS1FbvO5c9SxY+3fJ
4i+AIMRkiHR1QDuq7pqi4qpUfqIAHk5p+a8UtW20dJ4MZ+mNno78Nq+2A1dSro0x
eAA8Mt07Y2dCgcUDBLlnNmkP43D9aimc3dNwe75SOi7QTwTr2X9feetltxJT+47U
Nz/rjLZTXX7jSX06k4DX050AXeY+x+j8esGzUVU1WOZA8Ax34wfoITZW2ZyXeKZR
JeW4GKHfYFJHwTMb4GckLIJeENqhzLIxHKIeXSkxq7YqU8cVDnZtaGBIX3B9aQNu
SrMQ8cR/MO+97eZpm7RlAtw/YWP55/dDxZd0PQJihReg1mFZGUCIFStX7jAudATX
3cOQeNNOTjUjtO2pZHdEIlbcbSrHDJ7RvwMCajdhdh1UmY91q0HXndjsj7VENYHf
zXI5YvQrUF7CWEzGi8YwiuV2FxrblaJtSCQTwuIWG41mfhVXErnfB9ewfNMgWHHJ
LBdT7AVyp2VoF5Y+saI3dl/U6v1qHw/tM/s7UbIVdvOHd+/c7wCWdQJYWFlvGUEa
n+DFnBbLNbeZMRs14+AJiyTJeepPcoD/Y/ef1g6UDmR9Dzvd2lhDh2InPi0lp/T9
HPGqmOV4C27zDnD4/Z75k/+kEbUM8E8lMTmQ9XLrOJA+LvYHOLRET4/VuI2+hl1A
RiLn4GHs06InCQo5gtxhPVWNbpTGLXXgQRYdn4UqDmhoeyFuWfG9BWGRyljNE2XM
oQROQgWcCDoz+N0eqG8aa7zhr7XkoYt413hOpr6zLvYjbNzZcqd2SwcwShyVAknF
VaDlr1lmpf+5uzKnaXpeOOB0t/8ZWaR2NyxAG4au+2sZAzpUWm7FOFYJPU24WrJx
tgTAOgICqAhDu6c/6C9dNCq5o2m5yDr6CobI7PHKVQjAU795cfwo4Ig93FkKMATl
NeBBXHICplBDmOiOmKUugExsGreYfIX1lM6set21lx1vbLIxJuyd4kzj20+vWFaH
m3N3Xtyr53MlNbrhz4Ro1a33nzZ2tY1KgZosNqirss8xeXeJ2a74hrQT0AJmu7Dc
/+y37T/qK/hPSZItlbLjo73wpHkqacSvVwA+lcPW8jBIr3CsnzHsFr9sq6c0vuSx
b0BZ3jxmnxJXWt8+STDhe6OLJyfrRJ1t8tgiMOTWW/kAVoFLaddVGIsnXIArdoXt
mNNaqh+80FRez/EGpNZBZpf5e2ii6AYjyev0FiDxDI6PbNROutCdYHMiYMd0XFP3
WrheMUPnGFfezGAF87FJO6ZZbLYY8rhMDVslucaGNEKBbLIf1NGw24r9hCa/q1rs
QR32kPc5R/NP/gZ3uFFrheOGndPdBcsLsefhhdVerLexOb1JptcUj4SwfTAPGO/X
nL5fhGJdsXKzlBa2sgCZNVA1/03tW3QxAnOZOd+yDZz4kqrqQaZBGiwVbVZxnPA4
pZ5Y7i7oxL5ZEG/x0Ibv7VTzup3CGePdN2N9Z5Dm4+EKNyZ5vlkaUt0h+svAg1Qo
f5QsXq7v0DOUO8JyY7Ku8Nin8NED47RGDNprNYiJG8G4NpiAKG1XHLGx1uPBrwtn
Cy+G023ykmKzer7C6Y/MMghlen3Y7eRBEhMbDWsf/+UO5LLL3PZ3tizeoKmjb9rP
6VcIbsipO87sAhgYXhXi6KPKRd4Oo5/xtqinEM5GEl0m8kE4iWA+AjutUXHga3mf
7CjKHNNPAIJzj/CTVINCeEbHL51K/xvY3EVY+I5useu+/tknFWb08d14bIe1OsWw
SUhp4zUHB5IA/q5BVbLt9chE9ipozqDkWulovor9B1MtXhVsmruZo+3ZeoAqgFyh
E45UZVf3HVIkTtscD6SIPLvQy2mwsFgqmJ/ugMKJX89OKQXxD8bPs93GFxyoGuEb
ebJxrEypKh2SQyDIWTw8M6JPfJic4I4jH1MfBXf6lBG/SxbHuQOHEzloAp3dT0PV
W+MsrA3ap8oDOC+/IyuCQmeZSXvuIWiLk13Jfq2sODSyJu01b+V8md0c3AHBNiD+
oCG/dO9a4WAnmwJKb4ClScZOYoadcJO6k4KGt7X36qzcZI+Kst7XSBetpsS848Cm
maKX/lR73LVoInJWlmbNr0pn35ZmOR4ExGGUH/D4Q6w4MWSuO1PlJ5aDXUv9as3f
WLwsRwmRkk7e0wmublqCPK9XPgHwuZzDdfsLFuLuT7kGg73r7o94U7TUJ4FBxrZv
uBA0fcccfEmlv2lVsQldfrRbopvlYTgyY4RH0n4rZ3rLcnsTDJPrEakqXe6t09VL
NVb/IShxAOSa81w0DQcy+zcwMCzO3qtEe1qxPAS/EKB9LsY6fGXYkrol6juWkuIX
3nzUVfja1Ss+fp2uBNf4/5tB3MoWCt2cNtdAl/0i75Wlfyuu1fFvGj1S3U8NYV72
zwAe7PSiSOl+bPEbbzC2RomrkKXejek1aXPwHhEDD4M7M8aiI0AbQ8AAbYCxUtgW
VH4gyMweonPt396nUzS9A4Zxp0JZlgiEVGJbRD+/SL8wn6tld0vRqhyJK/+g/tjn
QpVwwlqhPnbEsKCk56VIbDlVDGvY2j/SrVeoNvnXAHPgYDlKJx8FXP/SWv3qkNps
hGMcR6dy58pKu7d1C88gmxre6HUvN2eT8v796aH4YoBZm3pigo9wk7FQ7njTE8pZ
BLZigFdS2sJmFRfbJqVPT25yZOqTZUAa55Sl9mg6LMA2A0wkc36GNboFNb9LkJ9q
JI9OQRBjWR5NTq9etr+DyeABpWns1fPjWSKouLSk91rBJy7GXSrJzfYDEaxBOWb3
PpQUmAcJHUOj53xVAdYd3BGO7ofNNnt+6VBANjjT13dt5cNsoQa1huLfUVKQI6Jf
nLFbR1N50TUCUMaJpEMu6cYEjgU5KVYASBSJLWczSKxa5DY3G9LevfKIJB9yPo4s
3icUc334Ows/p0k5npWy/EKLliqne0UbqlzztHQHZP8jDTnsXuZ7a1SAtD9/HLp6
TViHXlmk3SqsGLFm06bPYqqbiOGJY48mx/ckPfBJWu1sNQ5XN6MRlW16/nUKrqea
TrxRX1k/tvFAQ/k4jRwNT/RwAxTbLtvpRxiEvYHh50MxASEv8uBJXUTkdj3eoiLD
ZEEo6kK9llowIy/11CiRJ8r5i/wh4GYSfBbDCtHz2Ly4vsdq+/ci9+HSKeJCVXco
RLKwk/Mz5SQSV3smIE6ng1wfSGZ7SY63yn27TCMQRff1oQnFomb3DlETTS9fY22D
0cBcgz3A+40yiESE1pkQx9kDEcJSG5LupZvt0wCLrES/BVfkKWE7c3chvG9+9KF+
mqdQdrUZTftGqVZxjcCODHA55LiqL7TNZKhEAxaUGX5HQUriUtgrbrhBnmuEl8gR
91G6ZlBAaKxxAlaFj/DoAtwv2RWL+d7CBhBg18ay1fLJ4twdVxNXE/Dn/pWhbqrD
3w21mdCB0a7LzegW8FFZflbVv+xbhGnteuQkMj+xx067UVAWtnb2DdfGAAef50Yt
SHogrKACzonvdCzr0U0shYeFO9m9AcQEfR+AxoUAv4bEweoPBnTZob1l6y3uHcNx
AQpCuoqPWi5LJv9fnelhfw==
`pragma protect end_protected
endfunction: post_randomize
  
  //vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ZudMxFE0NhDSGuMu4B7dKUeSAZg3jwHXiaPpDe2aN7A5A/7hrwdYW9jd+kUjYco/
iFQ/xzYYDevxliceONYhggpRLgWqIL6fJvDAdmrNPDPtL+AVG5JbAm687bdj384F
PPCNBHCXRAVUB2R8w3mPmJuAEIFXmuSiipCVH5whnZs=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 26427     )
+q0c0qYqu8Qm2VrGOHgSIdwOTcUDhWWXtw+K0EGTse6hJQQpI3wBBtmFn5xR6Lvx
YDzDtpD0d/eDmCTypAVB/DYY2G0gg9dC0j3Rv+OXIYiY4R6y0myOCjp1b7c5aCsQ
fp+oa79t6Kd/f3bq6z2VA2VPfL9kKmruD6Pij3KPPM2x2QBACJM21ACqUnYpMUl1
lVxRBloRzPvQwHpNVVkOrF5dHw0B92MgpZ6Lr5Xu3zr1U8+E0U06q5xjfi9bniY6
EGIFh6FDd+SHzJdFDLU/1c1X5wnht0kV33EDz9rm751FZ6uY8/ucgqdP9hBXHEvV
HnYQO1wXW/40ZXXdM43IWciu9pNLk4EW66fe8LyYstO5WyFJ0LwFPyZcS44LPf5n
0wm0frLYLDCu7SJ4rFDGNe74NMvUgv56llUojklhpqybJzXAODPYvjRTIgsb+Bob
xK506bYaEkZN2uOlVGR2jmB1uqqaHmBkyGEJ88q3ysv1SD7a50YZIeoqSWuxJXzx
Ob2CqKaEjFVvehvpR4n1DEYIAkYT57FxaP4c5HJKyr1pS2jEwc4nsSmasAcZApGa
dXb/6EtYljolHdBkftvDnP5YRDHJsh8swLj1budEaHoM/5AIdnPjYsq8nsEEWsUp
MNouBQ/CbtkdCfLisWOCtdiWqebSo9Tz3ORNjAyDyFzgMIgBdq5vfQqnH3zzdJfk
BotyOCT8zuujSEtzd0KM5Wdry5ulRXxBea7gBmH7AT2KrdMCBAVTR13ui7GpMEFp
3RRR+ii49KACW9aR54Pkcw==
`pragma protect end_protected
  // -----------------------------------------------------------------------------
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
X2LxV9z5FbRh+z6JbigD5u1ATVXOh1D+RxKTri3riwqea57Yt7VCxQl0jklbHbik
q/oKsCT8bQ9UyXTLQsxaNiV8Tpf2nlYxweBQCUW96EpeRFncDHxd3/BEFZpbjMtL
GFJOwzaVciZS6Gt+xj2TF/whLIDCxBoB98d/v6L4KOA=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 26620     )
7ywR1UHLHO4o0Fet+HneAYK2VTZyRqYWqudmFY0YIfPdL5KDM3El+ol3oRqlj6P2
gCfVG5Qa9W2Azdd+iPkPpdSrAH+1nZMTClwBAgvwdcWLZ1Zr+3m5/cKHOMoHWQG3
mkADdAHMqCDOtZTKCkx4PjBkIIm8v+LRmgXaTx8NRBe7LTkGqDi0GvqzXeEh5KQn
szhXTzQd/kii9mBbaHgGRRPC/2JDTe491DiXBNkfEGNXx48CfHhaqe8EjhRl6zsz
S45XH/MxwcTQz5z8QGbowQ==
`pragma protect end_protected
  //vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Ww13Nl0w3MpW7oRDboSnMPHVBKS2+AoEp3pcxM8l68FqCIaPN+/mxZ6W6piP2xAo
iMO38NT+DPhqgrVwDPDhyF6YNstuuVrApVlfSdit5++CqZ7hHVgWF8EKCMxcpJC9
ItLJbqLhzBef3ie+fQkgf7j23GrT2Qc7nBVxrPjb/DE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 67448     )
Gw1mJKFdwGoaTU9D1Mjf1Ung9VrZMDYu9NPapO88iOEIggwAJdd9Qku2DFKyi7c/
bXFr+jBJ8P/+Xh/py0Yv5F5uwD06MxdV6BWAbiXhYpXDGdWsQgXOgOxx9Z0nbUyp
buCJAuUJWigsoWs3li8KEYGVkuKZPSezzwlsFKFnY4YSQHHT1YEwAYuxL76GMEn6
VBLXHuZ720FC5nzz/hpO5GEQCZIRj8sUGupw4K78OcvIwRUITrsSm9dJIF8BAIF5
fpjXg9s4GCeIhYSvtIZMuuzF82nj5Tzo42JVk14P73wB5JfGGFbvtviAo2hpiZwW
qPlNh808IIOFwjg0fQ7HRDwYVkWojskJqybHcMXWXKXJFxdPmg5959bUWdiQy8lQ
oG9sWTEGBH4KRWIMY1QdIDZZo6g3OFzJu4/iAfdSnf1qocf4QK4hDrRZixjC/m7Y
+OdG1GN9hAhhgz/IvMJaBx4F/rFzpWGAa2pxWMTpm4YI55XH6It/oZq3qBLYiThe
powTNuymk5vMdUFhwT28nlRaXLbDxsjwdhECj2qCECMvFVFgbCeT7F3gUpbVWBp0
mDhrR3AqNEd1dqOvVGgbTOs3FTLyKv1ufpiFgqYTJcrHp9JVZrBMDmhVmt1h1NcR
dBrZqmsYaghgHbPU2hof1wWUq3GoxZHqKGiHxvkUZuJ+EIKTY941SH3DRo1yN2Md
Ox1ihceVpWfxQ36tG2D+UJEFNJZNCG/gximJETOSSWsRlKdtCd1Ko6E5P/Fxuo6g
m33lWOlu4YH6lE/vFGBiXJv9sWZE969DpkEM10JTMb3E9B5CyXgieMOhSjkf3hoH
6Qe/V51m2XNYuYWzHYW741178VEKNVsqRxReC044NrWshpGl0luoG/cg+rLqvGub
XkyYjQ5yl5qDD6h699xKtbMmWIjn6q2Q/SD8IWgZin9w4bdmH905dZ78b7/Qsu8j
vp2KmJcD99pTSDlUUwPGny9CwwEwgcenwC8LlppNpueE+l5OXFJ6d0Hs8Vxy6F/I
3BfK0PbtGQCblGtu3flSedWyvZAWjkWGteuv5IZUWkJJD/bXHUhaxpUhhJCCa69g
UCbBG5cR04kEzZRIoJ/fbHZhiyL8PgqkLcLcWAi1NhksF0my+H3+oplkxUrHmd0x
FLj1cy0EeykL7F1+b+/g/HhDJYgJZOOSH9XdyZJWzuM2qzS4t0y5Ijn9sBSmJF3V
42XpkUGNRF8A4Frx/wPAVQVhxZ5QcGoQgHenM1t7se9aSrtaJGAsBsBHGQkdYWiT
OMP2v3bL0P/a2LUyZxUFXs2P5slAozvJ9mar9onaVouo8hBOxOh2/O2njcrdDBR+
+6zDz/vQKLP88sUKrluVWqW4x5DFQzYwYc8dAjhZ1MFsYpUBffLBBKxhlcRffsaZ
Bx/E/tnTZGUwV08VPAsI+T2C7mO0E6xRp0mzcjuQtRAYheOZnadEhJ7pL1pkVkso
XZdQS8221Ahsjw+n0zf5Yz7vfJ1mGy0wnqOcbq2RjmlL9yzWC+GvVRydWBrsMaAj
jmW3PmYgo0eG0ONA5mQd8HG2UDSmB1dBJVwGhZl6sYM/KBg4muOrmWs2bXkLl5WX
TJGwA5xCz69HLgaKu/a4II5ldVf1/G/SyGrk1eNbMPBXYovfT8fVc5yDRWtisTP3
RTng/G6g3ZRr6A11BZfxclLyY3PnaQknB+9e2JO0yUiDHISnOLtYHaQ8kjSs8cR4
uabL5t33TQI03++GhrjWYTwnk/wxRSQZf3HY33BHw50V/GfPZzAMaIf0x/HYSpWd
aDg7swOLt0M84OkVePJ5deRtnFzUq4eyEOP70A2RF0qnvFWdtSAXCg4lE3IRtXWa
18+FKb1y47O+V0pD5qUxfHISjJsbkI7t+Ug6CZjirR79wk9IPIVi4RK6xUs4g5Tk
iUzPZyHCUelk8p3N4GNDb9X86/l5pplsGXQ3xKSbkgvhcDTAkOfVoypl2He/I78p
q+aIiGcvI7yBMK6h9sSHrn2nyTwfpF/cRtkisMJo3GxfvAPV4sKv/QgZtkypV3QX
+cwc862cGr5ckukNdmvwoAYTU+cfzk6nINELYcQ6m6XEt0P2HR8g1nVhzQvDPvi9
HPHPohxOK0V1iubWd2tW17ywyLQhHuIdym91qC6F/dPm3U/eYtSfD0rnJz+3hJTA
ujWAmOjK4qv/W68ic5xrPqCQtvcrz5bg9GU5NTRaiSc56f8WjPZllQPMCqnyJUHC
JeBvip4vO7gfjpJKtjivW+JqkozLrgRElZ+jrf+m44DxI1q3Wky2AUBOZOtHQ1rA
+ee+6kxf4+ApYuj2zjqwMHJgc1lcssTO+aFPR83l8IZE4IuHG0ixalp6FGCIoiCF
PDslUu9G7MB0Z03DgMJ6WQlwJNm4NMHHdhjnuhX59oUyCvsmCMbNLotm0EhSkOJX
wTgyJEmHNMD7coLoYrU1w9Zcnmi9KKN9AZVMGLGf43cHuoexk1xm82DnH4CDeIxx
aNRED20UtwuGvBaY8ahXruFp3dLJGZq8FGugbbUSOvjOu1KbgIstOeu/paOMIWI3
O57oqTCyzsySDdcFzB3WJjBgc+u4EYjO4t/Afdg1Ybz5Q80ktLKkWDW6kJCZC+tU
1bnvFsdiZUgl2yqqQfqUqIvYHvNpBsVMkcTiTEABDcM9nijG/OW8rJJYAqy0BQ+P
Uqf5eiMBXrpBVcfukFy6lCWy+MzzI4lrff7kFDk6DP/heENFTbw3mIiNByKeexD7
hj9YMxgpMSIXoOBh+ZKNe1B38IBWoO92mUOjJ2n+/wEjF1S+zGWuSyV4eqG0YvRM
nwGA/uGSc+MpWQ9EqUY9pbd3pYUuD8jwsAht9ecgF9LQhBcsB6hJmqN5xd150RlD
RdL1Vbpo8PLIG5EtfguOXLrxF1F3S2Mw5m/O3Wip1PVs9oLT/A0VjwgUA4WFiAih
HNmMjaQ/lccs7jHCLpGrZJT52aEixFy0SY5QMzw0w5mBF4IFBzTrvUQQOmaAt6VI
ZIQ4quwVNuL8lQ9v88gwe2Wdp93BNTBqevDcY2B6Zo+8kjaEF4f20k0y54nHfoa8
ELDpBDOjbWUmHSj9z5heYQUd3HkgyqkCPJBAQ7BMsESVSA31zY/VVGTbdZtn2PQZ
aOR38jmWvx5beeH9OLVK31r3pkmTFTdRf5c41cYKBxxRIbJML3t4dZ3Kk1b10i9+
YPPKWZTu40XIPp34lL348F7f3LVkLUWc4hO9mAdRMOVEW9LQ9aB93DQwIauNKT+F
w2nGpBCW/uk5KwYrSKiP+Bx+NiqCR02MrB3pAX4W8kgnUKqLoongBH8r6u4+rgRn
NZjtrIb4lzrOAxflrRtL6YAXD4XCJ6ZK115KBF+HnIAc7yEZgRGzacDq818qP/6w
jKKcyxUD0lCB8wYoR00l/ctUE50KQaViuRMFYEI9UDyMhMa0bODTMNdTD27vSorS
Y8XFgIgCwrnMYI8bPk74VdZT0nw3R/5QIAMFr1O5t7siWarHa+sa50QJnn1QvULC
oQX1QswpVWfzIBIyqShnqkxam/XPUe+wIaxIDi8vOq3HnfYwiC6RCvQEoS/3anDf
YRkKgL1VaNkLgYuyxIi97V0I4bcEZ/NjRUf8TyFHFb6TE5QAz+ettZKRAanddbIA
g7+P7kAbVLUhMhW9U9pUZAkwPy0o4M5A2G7f/fqKRNRu9XzgRlg4RYYO+4771ZPr
hdK8WuW0yyZM3x4w+nbhy+u9c3A4ujCPjGmb64KJZaTnOhtNfDihF/wPGx5jRsuV
zc9NObUmvYG/R3SodOsLfq7/eMX+UsqiahuB+Z2VwHnQaasU17Gpq3/t/T0kRJ1o
nh4vKnFITZrQc/t2ILtYgKJqZnUgs0eAmcmFXSBu3HSuFWuyxrr53CM3pV18oslg
3YhtTDQzzL8S2sGEScTi9pRzHAXjtPHYm+0FZHKAr14qHNSZ/UcCcukZxE69pLXx
nLvqKXFf2ih+ZX6J9IKLAE/6JDtl/wRo19SP/qBh0ki94BDFcAFpHcLiWNmt8w3T
6Ke9JXoFVGUf0UVcspHvSQhOf9EISbQNmWAKdhAj+Bha0y44lwa1OxNohqBXtNBe
O5Q8nbg5o0v5Xn6vntKGYTn4Xf5Ou8/8EkHy4osXgXUgtAVMFF5rLVK91XNR09ds
CgtFoB+fywGZPKBgulR5JbUAAom5s6bxXfLs//HI4oVm3h+/5wBLRaDsdc+0RBu0
xsqEOOs5urfvsXXk+uwURdB5Fzne3ZVmXXLkvesgLhYVaeIaVOlWh/4GrYSnudsq
78B1GwTsQCiAhU/NgNnilqw4jfXcFNLReOyfV19JRBhFdClrPxfKdr/bx9YC6o7T
tgivS+luyqBbEdXJk+k86pOInIftYJ+ELOtIOlgM5NlWTSW01kV7XX2sZCBCToaV
p/4U5myORgBQZID2DiIqyyVMF4EaI7xQYOAmqFohrFSjNHhd7QhJxXq/FrxKXGsW
EuSSjLseGdJ/p9V2NX0D2/V55Vr4LRleHWDkxsIzaDSgfLQ7YAjLMoY7GUoGVaQB
4EzvzWRW6JbECkk0RWruxGp9+eRcJnFer+cXS0wEizFoGf/wLBWttXB5Fv7juKtA
LO9S56lx6l3lS20flihM6Ae4HrwagpmJ7c86M9PWzJUTcGj+yhDXIdxQgEBdhh3w
VySUGHm98m6IMFG2B1iKiL77dxjK8ULNvQroDLPKEyruqkQl4bMfayHBoqiTUWRC
RtSsOgJn533cUCoejWJc1z3+yVD0c5xce5nHAF8wm6OjD8PMUuWHG29MsUlhUtTj
WwIkafXasZMcEme4FssuCP7B1M903CoIr4b2sgxqOAsge6Cr2AzbRgZ4GrZ4AEcq
MLiExT/DzU0vy/T9Sh99Zja0iWp0nju4EtEcpXhzAfJzc/JZ0JE22kwYJ/vPfdjv
9TKBC2ANpS/T2lNWoaMVApaKWssW+JR51cHpuOD9t3MHN4D0fEMLcke8FIj9Mpj9
hFL/Z+tDX03WChbJnPoUQQDfRT24gK0toWfaQybqZ7fKPEXSujmCKU9okY8eA08E
ZusT2bUKBFdn06QkMc88GIbuwwHM1vDU7sgz0xh7LSFvJ2F5vIPbyBofZvWHFaRc
IwlmZYKWj8uJAfDaqLlD+LZJw14/pRjjgoDM7yb81an0oDBf/jjvM6br/WzEyXec
qMdwKg4VUWV/PDnHogoulhcH4cpqc5zIEdvEjpEIR2pz6X9FTBmHsnOsjXTgFHAL
DJbItz/fs/saLV6Nn1a0P9LZ9RWICMWhaZZ4QJQ4nwTIPYZGjtxgNSt+b0+tbVLA
J0zNCACTNqNq9ZY+gthjB+XNDZoU6dee9BsAgAi9HPekst/FWrtQY3o4q/dcymoS
Ijs9j64BDG2B4g26Bwt+dgMbu5OvXZZuCUW7t3Q0kUXb3eCH0rCqHWwWiMToXBNR
M5z3qLIkAKJgJBVWLVxazwJjKo5BEiYNnrLN9m2tNGebSrnyJteh54pJiCjfIDbE
sgSqDKkUIC4yoNDGcEUBuscdSkTO0KjLkDNcJGpFGS9HlOCuSM2OV0rD/Tjtc3s1
Tal5l9Ke2YmP/19Pu3zbR+Z1LO9UAEOeenfRZ5y8zYYlQnATbFleD+1ymF+Mqxu8
3JX71v5FS3vk/DvyBZ5h+T128L/tYHhYEOyFibixoWvObXwrgLQR0jbE0HHx4oGF
fNNFWF+OGoG8bATfCQy6tgJYA0VMZ7/UpXk6+yazVhSr9DpdCD2vWTXCUbmNaDzH
X9ovywQ5a3TyCapqUGdJoNV86r8MrWLGBJfJazQKqok1UmOCfXJyYXbJrlchJVCD
XbR4AIVe+gjoeOnSRNjQNj1Uxofcjg2RThjEjJKSLwgCEo3o2u29S9GZXssAVdX8
NDCDbFoTO1LiAkAHEIW1k0yJCL59Dcsz0Qa4h+9MzvQQi9jln8N0qXyeeWFKHW1d
TCFIo5vU7MeeW14sb26Anu/9UgJ7sXasYpKHSPJtC3LoDUXvykx0aBo30xAabDuV
LPL19r5TscBDU72QhqIimaB5dYlMf+5rgmUp5MYqsWVtd9odq71ev/wECh+Yyn10
xNetjsy5SajXUlxpiDi3NLRooRZcZTPJgYdNtKRG2MHcBxpuYivwMGmRMjt1TWuV
Gg9khCZQourDYUIc61Qk5CccE4EIjtoyNjS8Yk+4Lx4LtWHczv/TiTx12iuIRjhJ
IiPrCKC8JmU9K2gS7ihFYZAAepM4r7afl4u0byMelelgZNR1UcER8a+f0Hdjr0Kj
EBShCjYWJKiOat1dfgtjCZuW3Y6qxakcwyYpVfSx7xvZ6LwCeXGf+dgVyJ8/ndkU
ypR6SwTwAWIUYkI6YvjefIKqL/n/1GWKUOsPA6nd81sEj3WMfa2bgS+zlemi12tJ
hWhCSNmJP/zeDFnfzYk5aSm3N/8apUyNaRb6CIQrdipPdtojvEqX1PJYXxuoqFlu
gOkhdEBFX0g9C3PwPrB+5kTPoO9tcK2ovgq9o6r5oiqQgZlfLBaAbl3DNeYK1wM1
iEUD1+fvPsZP78FjLkfqr4GVtVEK82yFlk59Gnp0CSy5h5vI0Tc4YEiK2QDnUC55
GbnkPh4bmk4S6IK6qEp3l9510CmrjXq9GcmRu4SNFXI8KGr/gK+GSV9TZ/tbjkdE
VgSHNRvu3DkGcZMUdaMtumzfi5PzRWVuPYBQSglNveLAp9eOfCOuYXqqWZMh/wnW
/oVelQXogo4JCu/BJrFSD1eR2eNoDwYmKqB63I5SYfmZ2FLKC2Xj+j0AmVbA6HF8
MuvuhOVRqEjdGpxw00pSOtREHSAgaBJNm7xg3N+lwSEB8dHJj25/g//JksWXrRxy
XOSDXNVGGbaShT97qro5o+czPps3P3U5QlrS99NLajhhABy5bavAEMkXpKiX6Jjr
4qXUaOdvIkWRiBzidsVG/Un3yyjsoLr2ClF+hpof7tESoX6u3T7ZUeIpKrO+cbyz
EcYlHBiWtYMTe11e2moTsq0UASziJkwxHyxKU5mrPDzVXpEwlodBJ/9MA/arC5Gu
nkUDTkWHQq1gFXZC+EfOxq+PbOnS9m5aOxtxM123ufQM2taKc9QvSATw6dfJR2O4
UbYHJQg29eWU7I2ooI9y1nVm/EGRMrNt9luA2EcN7+mB+iAzvrNhXiI+6XCsqDgj
1Ppa4euSrdAxgnLZc8foBLU7NKARIcoK/6avLM2OoW6MTPhCaHdI02pfuYtzBA+d
U14cyS4JvyYoDFMytxBHM8Xk8UdMKW04ceoMEWrOCgTUDU1Rkta4/iUPftVDv0x6
vGrmTwk0oJ/4bEf7snGCZliS6YDmmfTpABjVDag8hFCKF78amXv0k/6J7CX4eoKw
S7WutJmQ8siwa0qcFfHJCiNeY2rFIylpNY9q2JkT0D/3P/y21KDF4pqJiF6dI/++
Etzj6Umf2lL8o0AFH4SIPSK3CLPOMuWA0Hk90PyGGBVE5ajoAh51aCZcNfQr0Z9g
+5BnHrAjULacrxeEkH2Em5yvgIUgvzuS/xXDuCqg0l5Og9yOv48SccgxxLo8Gqws
7pDfa7kxXxTECC/ax9PeYgXlyzpyfDjUik2jjACqKirkBFmRkS9u1DV/OOI+eOS4
48iGKEltYs4b55K7DmM70+3cPJrymfWw9s0C3FWbjqRROF6Nkl1J6NvovRVhZOxX
0Goxvt8exuPS1UcfmQmNyI6LlshD6p207IVOOh6OJewdvM/xtIIlXMJeQ/HWMsHQ
thN0LwK5439ZYliCxGXhanK6gMZ1I3uRJlss14jpmnyrs2m1o2ofG8QFErYijaTR
tYMdI3IQC80b2RaHTtPvZvQZHQJ6UZuuW10H0LBHrifV5Cilmt9y8QIfMA4+Ebij
NPfK2ZtaOZEM5eVtvrWGrEgbEWCkA9aAl8mYolPYxQsXekUWGwdajdF10oKeFkX/
4xc5QCRMmQI+HgGFFcdNEGhWUSbNtOOLS9CUPB9idan6O4GJBneansU/SkDE7Rrn
QmLiuiFMKd3Aftx8rC7KMQQxXOjSSUEHlgZ7EO8qiKsR4TSA9U7XfKLEu/UHIe3/
UeFajsOm6YhJw5jS5AO9l2gr+djm1mf6CsB7EL9J7JNPfTNCXn9XVZnCdAT24GHN
hdXnu00vPfW5v9ciA4XPTjc0ioorURvQvud1Q/gUU1J61qefYb1wpSxnBCZ4Ku9Q
p0n4u4npWVKnVlU+lN0strcX9AAzrGcK+ZgxMcKeQzaDHJsFbMh0QP9Ic6eLBp6h
35EkB7VUduzxYnU1SAUT/f3SEYbvQlBhoxx80loUpBJlYixG4LcSH2F7VyOkmbrB
jELmtG09yqxB0UjKolglP/jSYLceKh+TLio27X9hIIIhSqgp6XxuFcpUtS5zCgIT
haNDXMgSoPOyAhRZTpVxO6KRLmJxdzh78YgqA+ku5rkBCZ6QJvbTP6e8bWx59AdN
XX+r+VCCN6kNRIFZuR40DA74/bPS9CmbEaqW5Tl05BDO68f+VcsocrtFvikzzrMV
CpFJWNYmR/+AKtkj3gKxo4wKOyLj8F46MbOjupdjRpeyZNdaouPYXII4jBDtDG37
xQsbQV9Zf+3k0+vPkY6z0kfa8oInMDkKn7xe1/QXtqaeaVRvrtkTc9tgo0eSmjpz
RkjJafprsANgBGiRzQeSJlxy/xU+hbh/N7ykTPqrVMqfKXI8rGpqM47gxMp34ukc
Q0NL5oD5h11r0dYsszlImxycR7gxNLnKqhADUFRHTcuXbdEZlZP73bWuXO3MXNas
pw8BRqQgeGnApz4h+IXS41vvpqHBVA1e3nXERXpQdciTRtRjR6Qpp3SjSD+SPUX0
6aVyZHO8OUC5Ar0z3WtfeVGIDki0EAHS284uVsJbOCL1Hr8KaK3ZMqR4+w6JmCs5
viLejzdV+XXLZknkuSX6+2MQX7aUV3eS/wwsObZVVZ3X29zAkv9f+gAj22uwUyFz
g6BSYdKw+5rO0BMtliZHrPRaKEsS6FIUF5B7ylkoHmk1vSowBnUIfoVlJ/JnH2n8
3+3OsbWpDTjAZmO+NjwIKaJwmiJlwNu6260YsQJvDFLxk+Jbvcs3ToYNwjiye9D5
KG8S1zNMxRb57jiOjnt3SOLYOF2xQtoE1wMcSIOfRW2SpQklVhO2lB8xHe4tIIRn
w75K6uBFZvXT2WE0WrLHkPK+Pb4/PeBx/85CwuMklNil4JcOTO68oEEWj0w2w8eB
/U2jPCOEqWK8f2XDOzdhKT98vrTbK6q17OITAwCWw5UCqEWDcXqP3upl6UIBKhSR
EcHLDpLvcKMBOEupQ6erfj5sar7dnKjUI7/6MoZY+liXJb8V7NrT4hs2pfQBuIys
yGoN+Z4XbmCZLxK6TKmek9DtW9PMu2Nc8REn3dpEliA0/AfeLXDgM9m0del1f3YD
9q7cTxm1aLavm0Lro1IEPjsLWWI60TAceEnSaa2/jQ6D8x1JLZRGx1meGzMjl8VQ
TWODWHnN84YC4en0G8W0mLR2UJ16/VEfVPjhjeOaJVBQn5eg7bersc87oBTXbPwE
qaVB4VQ2N4qMehfAal9ZhFTEND43JcfWBBmkSmeU9W07v/Z3p+supOurO1nJ2on2
6SaPZoGzqA/Dy6k2tFBgYOglGIGb6eqDoPlDuSk7m06PRfi+WoeOOLWvO5LF3ajC
AiTMowHPsLc1Rq4hJVUgo0+I0/rv+Ouzj/xD7BcVcTIEDhJLJgfVq98h0u922vLz
6kma+CVn/Qg9SGyEqTQpOR7b3EdPVneIqKSuYEt+TknByi/kYiBancjakhtAcma9
f6bVNbLgF2aqmbHMC/qRzsoBSKi0mNsS5kX6kPBsC+rbr+FAvEFI8w3L2MyiXWwS
LYgkwf9GW0EojjiLTCIi8IDmFpAbMmji4r2fKM4XPnQ9ZJqbrbDey1SMNuwdnWiV
vx93vXF8EZGiOYqtLlRO3Dj3FAqDF+3q5wIskflUN3KEuSBVI9zMp3lSK0M9lVS3
iIOOwj0oSBLZ0Zb7o1dRZPu0Dc7H/dto78Q40doQGJRzIfsLERz3pt5j3mqmiUHn
vJrVyzKhdQNJtY6QakvpS/vmCjQYuevaDXi4UBQf+pRrJixdM12VDfiqs7mJR43p
soI348T18LYZ2Bn37KOXJZA5LUUmZsk1WHC36QXnW6a1ggKgEtouxaatXFwpGlyf
zLlqqCU/O6Mydq81UD/isqMQ8T3Qw1KMApFr89fgRBh0Mnik7Ze+/qIfmeWK8/sA
IpmyBlbFgnS4uBUweAlXp39Z6cdmURPig1PGiQ9R/u+UGZMDv5eScmvaVApNEEGI
iC0xDS35SaZKK+wmVVTHEaWUpB/gDh0MFhqczCVH0h7Sdx9g1YKuTKCNuHw3sFOy
dEs+nyn4vVhJdUKZJOB986F3MzT3DmUPiSSlSCHuJMSb+aRpn3sKWULxHvuRqoN0
QX6xjvbT9ka+d3pVQnxwO/xrEMMTF+93PrYun5pgngcEAdv/bX+ZryQqjAq8mHl1
D7VphFa3XJhgksCR0S+9qi0rmkI3YNVL+pz+k/Po2FQQF63YDqxesn5HLQ+Mm98r
hTqln/Mjnxv/GkxZbq/Q+5MgBvv4R+P5NAvkkVVgOQ1rNso0u4PGfsZWbv9NEe1k
3l0qJ7gIUfKkPzzohLdtnx61Kw01om7KRXuZ1mQEtCD9zSK22iymT7sIPj3hqn2A
3MDH71rlPdflnPdv91hGh0vXnzx8QeLB+eRvCDddbE+B4OFicRlWXAthB5cNGaCb
ofVk3Cb7dUyOAsAxx6A2qpFkQn6ITD+LJFvgNkJFfcE45efXEJWt7to3Ir2DC/Dq
u18cnx5b0uoa9/z7KUBGA0y1ZYxunpuUqc4/rVy7CEyMBpSLH11079rRiHLSZOqh
lLu96atgki+hSEbr2wXtfom/z+v7Zs7x7o4c1HAUT0Otm48vJzsR51lH1mkVJst8
zh5lSLfp0iH/pYJERTaRlG2kLB+GngTK0tUnUaiylcwVCyqKGg76XsT6zUjc6SMn
V4OVfC5SJyfy5pw2zxKb1aVxQJQd5rUOzxC7sRMER9XUFzXzThRR3G2W85vkfLtB
RXZ79k60+MhElf7Wfx2wYfwszSdoNqdqbUGbN4VV8OVzLi1AmrPU76tIuOdZu1m5
JkxDnwJn7IZqZTcIjdNGTmHu9fCiKYJ5sTJAozmaWkX2UOe8KTFEPciYku054tYH
VBv5YsWaa7/+J9BWMp8OD5NlleHQfQ7KmYmIpCVrwydOQ/Xeuc6CjEda6gKPAtC2
5q7aZfO2hPl1PEZgbEaCgyKrWEvOoeIWtmxzolyEPj+vxXylwvaoDul5vZ5UCH/m
0361AfFedscDxin3psd7CcifsUnHBTGERkJaONoeqvOaFO0jEZLQMcf6WC44v4St
nFusBJwdmcX9h4ECHLOyPZ60QkX4LfnRlHeJxAs8Xp2EFQ3lySGkwhw5B5BIW/6M
0QdwesWjCK1sz/Rwi21l+fOOQFiVOkMl48SidrHPe/q2cNiC4BneE6rRfDD7/L5B
eWkfDHmNLu9ODt2i57jyDTkL98c8AMTHCD2FsGrLXLTYvSmHhBdZU76dIWwYLrZ0
WMDtSg2g22EN718RTIwy/8OWtgiLw1c4TYhxb692ZXQUX4JaMsEEwyigXqlHJGY5
HID65AuvqGzT84ZTKfvynTMbndl88aKga/vHsZDvfrdgxE9DAKEZ35bWUw2TZltf
g5iQ7GrLViJ7InOtCFFQr/AaNUxWs9tXvbD1flfMyht9gnJUuu2ztaNOmyLXaMbB
roZjU5u/JTyC1+kEF8dZyNqY7HnFGuhCC+PXUUEVeZy7YOT6Qj7cpeadvH2HW2kE
3iO8aOLxHzmZq7otYCwsu8jdhjLFV4TSzOGd9cuTahJ7dKtgxVGDmm/SEZS9Hg5Z
z9w0rSB0p86n35cTF3DStSw1mhDHGSEQ45YBXelUVPi0mRDM08Lf6qnaq9M3Eqrm
BMmGSv8hTsGEMwafsZP/PSZ3KWPlzVKO7G7wFs0Jc4LkqnaEPBbJ+sFLr/eBj2jQ
rhdBTzXIt7sj0qZey0ruCnq06PfDCgZtCVUq/+6AyvbVGmhHq0nDngrv+gxDGt6m
oO2aBb9z8ODlKPD2DUdXQ8IZTMXfII//NhjDUMfW1Vs40RCWKhStX8d82lK7oCag
d0P+K2gBFLCCFj+BizheIYJuTHx/0JMiAeqQzgceOv3dot4d0UuhBeumEd5wfOVt
8Zi8kj9alawIKk3nPk5w+XntFmw/jWvYUpuiyD41CFCxoTt6f2xoHLoeHX516+N5
C2nTB9iItcCOwFhr1Tt4CVDSkqNSR6cvi3jCyWcsYgqxCwOO2de3LZztwZ2KHzzs
H6IvB/qGBEIfrEQmQ+MdVJLN8JdQ5rBwTGBQ5kXgqWJf96IjhRG0Z7ITP+dgAoeU
rZvBBjXtc/bEdYfgIrK7wYj9Z4NdMYwa800+n5x9QW77kN7zWquIzxzZOUmX0Nfg
XKiZNQ9tIw1UVG4v3E5RPJewfrxYSBEawuYwVHYWDkD4wqyYY2jeY+cWNSFCQb09
Z0ZX4pFtsZ6/20sULZKcw4XfIFkTWweWdgUYYnMCFH9u7Fa4kz4w17pduZnvdUTd
A/xKGMHgDXcqnQRAYMnA4//zx8DOrYChd7JyoVnT65KvLnUvH409Y0kAcHc3fTQ4
dFdJB7ZYE0N1XVNt1af4IoSBcbeBCWHCkN4fLI/APwPow5/Y1/ohJZRdJsiKXE8U
uZtpO7C2kMoX0qfuyQykveY1eEJCYVzkoM7Q43MpwCcF6TxyHGmfIoa5fD9phalW
GLZ4DwXGaY141q4ueomXXIUe0ghYNQh15vne1DGNnq/gBXFywTR7bqbqclrlHEN9
xGJbzd5LYxvPxF1hsmfmKXzt5ziBJnoTOTtVgX+qnBdxBidN58MqzflSmfTM7h5G
EjDMv07WqOhsnjciOL2DVYjwup1XzS8Hpji4nPTjXrTGuo0+8voqKn18bGfdTIGT
1r6+xCasGykdqCrtaOhpjdpXwwr0rzA9AD5PmP1xm302ILgfvrx+RO6Uc7RI4eIx
yB/a8Nb9rzOmgrqSQljocFOYYyvioE609v8MKTGIBANi5ACacD6JNz8SbJn3inBT
zpUbGhUOVnOYNXyelYV6sAZsSizyW5hHokw3ZYX42/aU3usf+w6Q5ffbwlB7XlHJ
u1tNmkKwfa3FfrSPHu9xlEh2R9/bh/zjBburnY1Jd8jDyk0jU3rvEtsc+Tdmd99Y
obnEa/XJSIZIBLsPBEs0vxhHLDHUuzn1avTOQyCOItbkAvI836sGnunXmneMVoqe
Mgshn4p1GmapB6yIgYTru9gqF3L9GQ7PLzdVmLL4J5Bl+bU3YCZlGKYC0VUVj+ia
Lm2aR04Wb8awDj9u0iyaPO1HmpCGzwOiW3BDeXnmrS0xPoVY1B9IK2p9IJg27Zfa
uTGOPjwmsKkzenUiKwhgj31EJ5zOt469JpYbbS9o5SecnadpZUZxMgmr7rIZEbdq
DWFZ3YNnZMJQtYsZa/gzU9N0Nv/6jmEhjsh5SoKFy+YdpWCd4yqmvp0j66oe0ZIR
saA0GroViYdZ2MFpZFD4865s7tg5XEkyX3l7CsPlG043Y9P1jZdmJEi9+d5v9mID
hLAhXqcI4oQKaryixHwiZX8p9p/+Vsm9TwK0Kbx8MWLMxAE31K2GUfdtOwjQorkH
UAawBBg8QMUJv5XdKvSU78ru+SnN3CFDAMShXDSjaJMAVle2hsItWgdYJ/yQpi9l
iVVaJ1QZfTOa2BgDeEY4Y8XJaGaER0z4OZcGNSgjePXztuGujjYsVOzFkegHmFeg
NY/yCohB3ZbQzflIx91uGamYYXLfz3dlxSRdoR3LgrmvPLhVQvTg+OyZlKdFV4IU
FRIOrDZibr3Ez/D4s3KO5b2+StAqHMnWeaKz4fQKjD05Ajd3TSzI1t8wu9KthE29
t097MsRE1CpfX/323a6X1LrYEWHat8xfYzYXlaA6na4Ef6VlUxj8c8UDuzfHNUcd
evqSIbK2AE9nrojcDkcDWe/2Nq7SeMnynVBb9UR4otfzCUmcfETMOyUCvLZQdP+0
wlX1eOPYAcFx1+wZ1tJnZXzTts/oNIXeLwYzBQs16pSQ4hbc3+VIK4Wvbf9tMfqW
S1Tt8iJtN3i8xWXron9VPJbx1A3Iz0JeSAnsv4Ov2SmNlDEMkbbvRqD0e+33S50t
KCPcB6rBTBT0DEmsHz2LXJj/MRLVogok5C44AdTABguBrjwG/WDecycekOC8S9uu
XkujaTPuSecS7DF0KW57i9Fjng8YS9zy3H3velZ+OGaTD7S1G0Ac/pEo4pAZksqv
eU6oRETgp4fSaJziozcimAzt09GLIIxIhKzpuBXDnAuR3jKzv2oawse4wrYklpLU
UStk9t2Zc+yuK/9q5L32Rv53RJATPBooqI21fawsMONcP3AE3dQZI+PfxEtnGgp2
b3cJT60aDiwpgX/abdmlEruZwYI71YvqJ1RRp9lWrLdMj3nVBN0tDji+ONyzgkIB
ep3EsIKSs9TaP3vka6mvYYSFlK6T16ACWrB6bji8twHYnBLc9Xf/SE8nVDhLn5cc
FlD/5Xy6y3HsJLFq6lxBherOd/jTG2YAhnvcGiGbEgm4OUTzzuNDS1Cfdf1lBiGO
qgbAEhRc+fo6ZPLS/RmZ0TyKipFOTUuHD3K3f+1w5pVFVywFOlQZZCSl9AJxORAE
OKCDSag+lrgouK4TMn8Ymwk6EI3zeQfNBoK2ZyOj0PDqLKtbKZ0j9bVy0LIkJUxO
UnkmXvfBFaQUteSbHt/vUi6Cr+8v5Njp+MrJdZKERZwGtcAsyW2ErKXx1kW+jApb
xKNQaZGkiBHG91kdNEIxLuEYr2zQ3Dq8o0azViwV5SdLa9usrlB2U3cXPIabcazF
yGWBvfizBsNgQ7KUA/fqFIxSnVloBmunfLj8QvO1EdRjZIjL8uOxsorNCncwHEOu
AQx+4qxeOOAy2+c/sA1SNKRqMDtJRuTGzPCy9+EMKI0+2KCyccL0g7jkC5QeNFXL
gsp370is3WlAjahDhWkdjkyDr/Bz9AsellKiNVwWLjaJjNm7zIoO0F1regGymZoK
Szt1pXPejIzPiuXIcvtzFPyjay8Npw2hN5eApbqS0p57SrEk4cx0lo8wfYD/RO2l
729BpNP6MtGNxf6L0/Nk4RVx4ddtHueXveiH7EAqAe4+1tlCYCzF/gZtKtohwhwr
MS1tdoYdJtR5cNge30r06QagHyU82/1Z/u1cUY41lSQyqD/Vt0vDyPULw1HzqR9T
P/KVa1KySwYEzN4NvBy0McM6fKIL3U+Dt27GrsYNXu49KEoz/fq+YMQ1HzawR/5u
R2DPnCcqEBPm835OtxvRn5LFw3p2RyUyrh0611SHefdi8Enx8VKUDvQksgnKsYZ+
1HKTCo+CN19SyeRRqcnyrN/xQ94g6oHk8h/9Kaylt58WIM7uTOnsRPbeNFIhDLlh
iDQZtSKx8OeKhYzS1lgvo+xbSM657r1zDjSRY1iXOW865RanIMptcBlKiiNbYiqF
HZa3aZDZLrNz0vH8Ju07UshshVcAKatGyXIEgJAWbZMgOell0EUwT5htXB7Ksxad
2ScMGa6e7bCQFvAvrWAG+8M0o/vffsF4ATcyYx96ht5Af0dSsW9MmG6O/oGpjZWj
7TCoDRGd/2z7ZLjF9dfUAXdYt9GM2ZXkF5KS/DwCyTeSyjgCbNgBtuUby1xYXxqs
PzaQAb07k1m4qeqx5XHgR8gjLcWwvtOz6sTFg1hKlh4bSbEdm+PNrAA2dJSYIh4O
YUYZtuf3UJjxXdBgG00bZuvM1iDIio74SqmFyn6iAf6+DFxXvZ05q9P8rOoQdc6p
DapKKvUBkzkgIcZCKE0gZ0VFHh7wZd3jT2ZMeCimRDywg221CgHvE5Kat30biV7I
mDocDpWNvdgmotbOtMHoOtD7h1vxQ1wZ9jfyGKY+lKux6MRFdXiyDvwS/E1A4c43
kKUkH/Z2Py9gwaYAeThZyreky6uvofedlXSEWEZHMP1OumpTx/ZK2fSXDx2zoWAK
YkMOCq9rb3IUy3WdE51bLB9NRnZ944iIj6TSSEoKT11ZOxaR+aQIuy/bWpfzalMG
MeKdLD0c+88DiSC4YapSs7NZ/ZoyfD+S+9SExVOT6F4agtDNsDPTcINk6UnCra4z
sljM5H36XI4hGK5tDXnshPXm2DECEMERjEEo9COM0ELSK+P8tVmDCBcshA3j3YwE
lZudrt7oyS3A6fA2ETO1SXgklQWOzoPoVmcZDpjhrB0yz5lw0dyn7wc7zGinkzaD
T02FzCZx2TtnlahPuStwNN659Vl8kBFhX/YIRMUBrP3VGbCo1TGpwdvSiWKBPaVu
iQoXYYXLzF4g/xP+c/EZ6OfV4c7HX2czL+KPQhX20gciJ5NViLujrbAu9/ysVBQI
+DILL8i70rANtoq20zmjp4/ueKPuAVkxh+XQtc7Ft7kCzspbKtRRjp6zelFEaDl1
7pzfWQUePKUdTow3LgXrTc95nbshWzlvPvplZL7XbNUQV2NZKFVQ2/6bkYkHaswD
krJiB3ApEA5Cj2snjhpdCQ1ITra/h16NVgCgjFN8Oh64vjHVk0kyJs9BTdvzrUAz
1DrZSHESBeSGDG9+7BCm3L1Nocj+GnTx6Nc1iac5O+mPK045FFin24YHr84Vtprg
71VfwNS55XLQMMN0LoXd2kEq3ahnrL/wcs0Exd999pYJFm8mUfz+aPXaFuB4NS0M
QvrUu0N1zjMrdi7hg273/OsbvGJ/fkM5FRBjZYJtN0lBYFMCn7eixbcPTb4SHPYx
CM5NP4XkQiFMy2AHt4hsrhMx1oFhOqh0Ln7GE1sUUMkdNKHEoavXohk2ZRRHv7CP
qpSQubiryrIRcWqQk8xCazsA55FZWk2gDF57ReSdxyBMB948U2xASIFGxKqTo77c
2elsBBUg5pYeq87T86wrHqman63RiQuWK+I3j2v2Dr/44AfTBqYV+XE6MaggL4fA
9EWF2VGrnkIdMyYraxK4uUF5nB+Ws6E6Q9+y6NLpJ+VfUp9HUct4ERBum2OPrtZt
2QAXgPSn5zQu4PiZaYU2NVbnJ7BPqcXGXjlFuiMuGhd+2p5kXz7xwHj9nzFLQp78
kqv7XGIcenOE/wbsREehOFIm7NKIy6mmhK8JH66kyf/xlCi8cnJ8zBxPrmb2dxQB
uMEpVTtCdpH0DpqzsHXW3pQvyVVSynD+uUlJpBJnE7G0WwocWK0t0OxVkuUHAFm4
6PyHE1q8pZEvahjNbz9oZcyTyN7eVebukq0s1wT1Ms5J1+IefwhYUhz4D915YLvT
F4onZ/uImhIP90qRgAw7uW/4H0im9VyA+GeM6GKKvyGB7jEeW0lZcVbXK9aOcf3b
CTfmZYtdTYENPrkZXeipusyG/sH1dfofhO/Ns6/vwIv4poWIslrdmFe0cQcfQ9q3
uIp+PdXXB7q+eP3hSuo+d5VYRm6rqfhfDbHAuYzISaG8z8cq9vc6u1/zxtaT2lgB
t+IKf57SVKEgMSkTwsjtTMa1WQ/GGVVHr2imuqr59j9Wgv5MizxHLh8t7ZYvuDgX
j1UsL5L3g5jX1huc6TAeVdPl4brbY+0Anv7FnP6rwOx8Zo8DBanY1rJaMdXrKJGO
hA1Pmmqj/B72CsVvJLTPynUDsV8LaRk1M5NegiolGJMxXr0Izd5grtu4HILfoaQV
orr2fPo/K9b+UQ977WCT+VfQmVzgMevFfBKmFPOcllMESpiQaZAjoUeUPEm7YD9k
uYY5c0GsYj6LAnorZZkq8AF+HVZ2i0Y6nSFcQo0QwCHtdkA841bfbwQDeq9dfFBg
M+g1+Y/PDWvFPhb1F+HJEz6mtHI5tOPbOCgw7CdMsZJtCIY7B78bRrpdt84uMBKp
oLE/jZE+gNU0yIweLEF0ba0R/Pyjc9nssSCDoW/lfEtIW/xbg9caepvwAqkUnFmg
bbTTAvdvVTptnm0N4v+kOjSvCvW7zqFYsDTJgK6V2orqukycUgDtVPkm4ge4aLTH
KiqEcPh2+sgdWxLU+KQUAYQYekShtw8s/YKBoJK2UnEG0gtL5SxolgMsq3RC5hjs
k11wawrzjGXlZyLIdvf2Yv4/kTgSQwqHaru4MJJDPot13r80JL58+FH1qtHRIArM
rA1/WA8mG9CsurK1VI5VSz+8kSNcVSh6MhORMxejqz3zugRReUvIpIHt/P1oJruD
/MiOxcDZ4mBWA6OlqgkdE70S9/F7P87q/SIXF1dJdTbTqirfQz/AdA70ugXW66sB
hOGzulzhS6lY9brVDvZucphOgy/TJuOdTX1PiBVEGIxPaicMr5Ak9YTb5sLx0bP5
ExbWcCrtEN2gBXVZroJSyEcnowcDXRJvABJd5eGxYr0pB800p0P18t7psMS4xVU3
pjhK/dP2iTZYdlEiyXyOASDpciNogIgqSYzbrPga8t0VKE+GRoL8qPP+OpP1iJQI
unFc5s2mrQS5b3+AoaLuHJ0ZRnuze+Qrw7xZ0ekRkdNZka52R+uFxDb4Iaeym21q
tdcE710W818o1lxwdOnijOQWTa8NnDH83UsvCyGpD+bvdhasV5FbjrbVsqqW6DhT
KVPKEFpGcRPI/Y04rCQP1GnDb3I2eRP4LjVAspW6nU8EkcDoCWkF3cBIIaFVJfNZ
Jx/enVV8nVa3jBhVDEDawJk2ekubmcRlhscEZyyZgbPxfouvU2NYKZ/SfOSu7sh8
yNtZj0wSKk86aw18kBkW64QTgCKJw0oXS2C7DYIE3p7lmG7PbH7Zh2XJB6ChtAbI
x+aqAseA35U/r7LEzNvArnQgh30answjV6TEz45o4k9GaXxt/Wwfx9+xp/kc5Gwm
ITEHjeP0cUeQqVnDXx7sqV0SvpNTe4wCfVxEhIfG5ayfigIR8Xw35RBhQEpaz8+m
M9dBSM8jAZE2oPLO4xofL4WPSUHDw7M6Q5IItgKJj+PQvzBBeapSK2Ay0fNLtx/S
FjYHSELTIPN6e+KzZDP7zkm1+qweUUUj5SH8zG7+v2DcOI6zvL2qXABA1MfLvEYb
Fx3kaFuneyU8l8RNaDTmq6J5ifq1eXlFoHqdKsZRqzCNgscQi3TtUlNFgZIasbSZ
sRUosuAeyWnRgglZUW79tPbjOfpq1Lyuzq10E00e6Pm0qbdQ9ZLG6tiSmvqQcMp5
WxIZuVsumqdJ4wGTthGJcUNf9AkvV569z9IA0rIhBNHshtexNwzqUKuqLG6EXVPX
IV9Ka4zG4lYAlNURHxQuqLPz1FhAI3urz9QC2RCIS3NKd16pUlcJMFePs3aV5nca
jReEdf8+Zk+csC/TKLxBJFnOz8xeveJrJzKkj6RTUql5Zhwo4x+icuoONJlJtDVJ
uRAS+8UqbR5Mokbpx4VZ+25z8JWN02NcbHDgrAF2ZuTLvB1RNqit0M9zwgvQSoYM
azeCGvXNgRKACPY0ABeDXweaTz2jvm1hZih9Ofrs/xKnK98HFn6CvRY/G2fNZoTz
IitSEYzOq12EDpenKjQ9UbJLvssNkrd1653PYam1mE+5C+pRIvRJWPa+4JglcRQR
Kuxp7b0YO7e8z1MtN8LZ0njWrzEWVFIh4+wftPLNJlojhv5Iv6iOnVawpvf5asUg
65mZzOSJzxMU7/KST4GXcUenGPSMuzbl1YAo88FiLocjMFMiOx24YIg3pyvDbLHo
sL8rToJ1U2ib4HHi2t67ICHuIVnEmfBaJI/XPXra/z9tm7PZaZXw4RtDPawduvJR
AqSYG67CtV8ZY7OlZaJ828zxj5kDcPM/FfC0VMys8H8h33dVNKxV7zCkaE+UyQdP
Olie5gEP10brSkjOXNPBB8gCGZTHie1HquiGJXL6Zk7VDboVBY1586rCJuI6Z1LE
HAmlrb3VOANhJ/1ZnWGRSv5FFrpYaJ8fl7MxuQzrqMfVjBSZxObFnJqs/SdoLsne
mApp9x7u37MveOpJc2V/pMN/h6aOVKPdmHVwJcxmvBpQypt6Zvy/lvEB+JiHeb27
b9x0LeA6qkdp94TMkHbu7TwHEzUddtjTsyJP6/37GbR2MbE2IjZFx497dWjMxhYs
In6T/fEGP+6akcFgbRqMR2Ia10WzGZiyr/BFaeIf6bFYKTEnkEP5i8s2BWSZEGM0
4zjQWJdvioNVB65kC1Q5dxS1nMoj7tX7FysWZs0Y2onU4CMv/Lv2iTAp1gXdqKOE
zz5qk5p7m5BPgn018BYMhywd/DfKkMdgCPINQZ7vgwiRXD84cUvC5oIgj4YTlD1M
7e/6Tej3xk+7wxWH0vFhPkpstJLeYLEjhD354f4o+GUjkb1SLrJ1nJqKeEkPrlYh
uBoaTnlKv4D8ovTB5htBJoPxz0LLOY8OOs4VFZw0iZt5ReCx/zOBjMLX6me+bigI
SE4HiE3QY8gmw+G+QmmM63KSIZBDkR6tPlul/eH1RPg2Kyfm2unueMPgIXT31fj+
2YfOr8GGWBH4iy6heM2iHYD46MMPulHbRIik3XIr2Vd12JWxjubKOavC2ie18hm4
rMUr4TfwoT2vCD35vjVjApMmn92wLFTs45OLHQ8nA0rG3/iBZSXxH4aQRhTq50RK
Ua/0f5og5OjJzRx4Ba+QfEl9r3ML3VxCAgZVToKMMsGbEnGRVMVitcuaAn5Sg/Xq
aoW9xUX37nCATnC1kRpm1rSvYn2adEAEA0mfsMaNhTZ4jWhnxchtkxvMPbOQxsbo
hJ9mlRDOslYMAVqngcl/7jbzOAqSuvWizIbB3Kq9QpHMqGpU0lx4F8XhieRbZfBx
rDOC8tf5NsrtfkCsw+P95khyEy54qR5owHjHiEXXMFDx458FsjqvoCR1PEQFqE36
1n23MKz46FbzFIHw0nFCTRI48C7H+GnaA7Z6hcT7Ry+6k4d+4cy/kLhjxKZRAbMi
Lf0HWrFHNSb+yqvslsqpegB+73beLU7LHEGvhdzSnQ8XWcdGVQ0Mx6eM+bThHWAi
7Cv+/5WShSMYy+U9dn68vlHtm/SHnWPms67Rb7ZnmFFU2++V+hsM7dElbGL/2KYI
6evf0Iwf/FwBikI1ASDvHEQYobT7yEAJYVn0B/E1FyMeNZyvikd417xD9YEyzM39
StRJgxfJvCVmJHOBGJmAk4xcMwCjhE2hd3m+x1Br+rYqWSzWAKz04iu7XOPWieAq
q1NhSVPLMyWwbVNYfuM06sWiCeKW6u3UzZzmVb8rOfZYOE03V2D8NvjRtN8RLwuv
c4hM6qVCRUA/HGFPB3G8MUF3kxi9ucG6MZGvmu3tJsrrTqu4Q5AM54NUMfbw7Bw7
8OEg7dJMj5JkBysaDpKWtS5psszg4EYvAlLJAsuYv3+BFMSPwVM5OAv9/Nsw15iJ
BXmOqfgAt9+K5ywXNX66d5jjMe8oeie8y5djsZrM2yW11ZIk6Ph0Tkxuqolxh1+H
EyPG6vpvVLWuCcKT6nDqMXxHLD049lNPrgn2vi5Zg6qfDRyI+qhUlWU6VrL34+Eb
nO2sCmHM3j/rL1lIq6sNgCIf7ngi3Uv8zPOg1NqKc4JKPUPz5u7UFwCed/iJOFfP
C+4NkRcMHUrBfF2UOVJWOrzmPEZkRTEbBwfuZWa1FCyYfgsFzzaeudRZlRdpP+op
sMYkmn+rynhNWwafYlw5n9nvbWNxM1nKV6mjtf1bH7yC6MArNlQkZfJRecqVR/ZN
SIiHQj2tM1x3ZgpoTBi8lHU+hvrvY5zNdr4UiekYT4Dx7tKIUHejIKf/eIcYMhg4
xCPhM1ay7Cyjq8/85InXUjPA6vz23cvdhcCQTFEfk6LVqvXD9jjLinWmGD4ffqhl
GD5lCEB07/WmPpbfc3F36STKf1gt3xQvyuVqZ4BZ5uoR0pP35yXQdB0yUzG7P4tU
dJrade5cW3n0WkMq8haTT5lngWL8ryNNVLzlyLNSsZ+L2W0L32YFTSVTZ0rYlNdt
D5nGMoHJ5grU9H9jFJGrBzPrCJKfwbHXdzz699xc+Jv/GgeN7UekAOCFRLAvrbVf
qUzS27a+o+sG3Q7HfkND/959DRHXRMKTCq5WBfJdXrq8xgIAI2xK9EXbeFvWIgbi
gHGbj7BPCczK8DfPCyWHNDNscfV7VevuUDruihK1sENIIEewbZYyV2UxiWx08Mv3
aw+zy1Za1bUM7HPUe61KlHeHtdJZkf0nv2+dH+5qknaBtihsghmmCPTyCLn1V33W
8HLX4Gw8Ljp5ajaZMJBDXMh/3vgE6DB5093HnwRylT2mwifzyW6Ym6o2MgfoT1B/
txLhHa67akxRTjiLyXC/lO6/+yC0AnTkvOR/KK3ntbZB1K15X0GcX29paoyD0SC0
cr4Up9X9M96Jn2G1l0zibzi4yZNpJQVUdn/V6gYIoUsXPquE4HQFBBtbgaY2wt3p
duJdmX5+tCzNLOXtaWZ3icMCyfotUta4JYpDKGgdTlt4ZOpuSjW0pW5rRYN30/Lj
nWzIm9M3j+x8VIKUGxal0dj2+CVgP+lowLgle6DgdSEZdLBL9oHwsUD8ICoahdjS
TIvFcEFrk2PCVvGzGRcxbXQnld+NalefYi2yZNQAiPza1pWbolAUUV2EUGAMG5oq
79UisTx9LPfpDsaaFa5ZEaZZz+quXAYmkGXvC53Dnd9Go6R6OMejGb1aW1lU59w/
++DlVqHdyk1sZoIr/PB6gqpxxhZMGLppGk/cK1vidBtySlSN5FqXPpILHDyL0hB4
/l9NC5rrW4PlD/mNY5UVRhGgcMJKk962nNdiZpuOISZbeauU+IbFDvOZqns33HnX
/pK1DweaSft4y9voY7AfhmE72j24ta71YflZBBY5gwRIarsY3gjqUjpS6fvpm8er
j3hXflUEWJ+98xEJfrMXqcCcHxro33Okix/07Pzx4Zt6BKUoWTPhCMJldyA+lJ93
8/xqnHZxBmhE3hBFKGuPNuIq77FHrIHvZ3b/G/R24mvhpYFoyDJwjttrGXNngxrD
gEezp5j4xUtLVS5Zzbfji8uE12LVm/b00GpyHTJLJq+m3tIfWqR5ZEmKBRAGfS16
QkM9etidguPdQayu2L4xLOIiw8yopSB/3JwcZWf711bRd6tGVaT84/aiYGWHYdXM
IFZmTRpQWXW1WGf64WBMj8tIRLnjK6Agfj2WcwHjxqXstQY4YTH2S+y+LNZmL17d
n416f7TApzhu30ZZA9E90ba0AMIGXRjnK7H2akLZiu8nP0g/FOQSDQ2jioN1L6b+
vBNX6UB8KDGLalf/ke1jDleghkhqbcm3a6ts7m2tn4OU3Vz3Op9znUbrbJB17+1I
CQqwJSptAwIxkKhe3Jwgfx+2ZiXpk8piJ5Z2F/lWf3v861WdOAb3u2hFsBtFffq9
P12RKnvDLvP9N2OSwSZwZjvfkmQvJz6Ymup4jxC1Xs9ssjpVbVr66lQ15oUQxiRd
bltE9XYbgHWhalXXwNv6Opj7DEHGlDHz8wA5nIa7CkPdc2dKIGbW7JyF61ZNM5CZ
ndQDbc5d/qk3aOr7B8pekNCqXW9eqs75h8euns7VNpCzjZzK4RUuv1UssJRIcEGz
eW7Af0otcddoxoJGp6fpOy0j22YBQiMjmVBMEmQpg/baAqx0UTcyRDohECBBgaOX
8y/qe2vp7Rk1Edx/USW7Hh9i4dBoHU5D6jL7/IvnW4xmgWx50KkMK3f9+N4k0ObH
f5YhZbVTLKxzyeoM1qiqXjxl3pqIeIKETG5qECCCxo2YG4Jei7hkQTfWGMVVGpTA
smCZlPoMzTuYA2uaHbyTKy26v6CcY+BkHN1ot2DLqCBwBd53xXWDKmeNGv0Jg4zJ
1SYKf+3e7tgJCkd57zpXZzq8PGVc1jaSvmZrbXDjZcwt6XTBo4tfizuHpPO2MY1Q
tJF9gnTCB2oFWDfd4tzx4Bwq0+AUOf2ZkiS50IokFrYJ4Ja2KHvvHL1WpOw5NrCy
KdMnGQBYIXVbGrAa4gwdN1s7ewpCD45s/Qu1k1H/Auiwz8a14e9ABUCv2gW6OJLd
ThDtIy5VAVWxPJvE9j07JgA6myFpMvPqkrt9gt8UFcIjA3BE+vYfXfBhMBOvNFd2
6BUJGxVni41948UgVe5bGkJKPkMudFCoZwwxMgN7FoDe699f36y/0yevHsTLKhAg
ZZwR/wxLgJ4PdkKI4OjqAGjR5dfr5MXRya+GUWcl2R0e/68wSy68O1SYOV0vAsMG
SDGQf1BplKRj7t0vxBZgfvfoH1C3m/wQ1NxrUbdXUWvbx8kTzPNYki0RH2z3nLp8
J47lgHRWBdeQuypdC+DA1bP6DPE9JVMeA8ejG2Q9u9QPll8nXBEzRCkubcVIK14R
DpEbozmwmLNijFPnR6ppA3tULWzuLuGhrdnXp+c5WRllXxUOgdu++SoRCINKdukr
8dFYLUzsS/KK1eVP2Lb/Vt7zVShmgkpGp+fw5WMBrEP5M/91c5BHYwo8pocDQyk4
6rAQ37vyxZNkhUeuxmqTUcsgfuJGm98eYn8hYLj306LOH7n0kyoyb20+AHYqE3n+
5I2wwHWKFQuzxJUI7CitMIDAmXih+aJtZ7/3ZeqDuWEZOUnd0DheDr3Lcqp7+DaT
E75IHENyVqhtKF0PZDg608SBlX3MJ5PmNHs6zDM71UjU2Y/nf9N1Tya8OudE7f+q
SaKGnesRZbgXLjExeVLVK1VUQcnc3EcT7ZJFqQp/8OYFwyFnUnPDSD+bC+pBmKOG
2UELQvW5h2l7/nxi+3QbV6U3I2dYWGSx/8KT2ccGg46e6N4ZFXdWg3UUV/GgYFYf
jeUQGaTPkmgUhOIzCdZpNOPhDSw5fUB1Pb5LvPVxfhINqxQhtnEfHoEFZvahj841
KAV6VLC+XM3n8iE3g9xijp8clkna8JkbVohp2WmIX/HlcQcFFFAcgOJrmz5J5AHf
wJ6VxAK+8ApMj2RcPdGlAbN3HE8jAiQJC0MFpbdZvxErko+9wrG94rrpx9SGU5MB
2PJsb4XxbM+eXG2ILEjWUexIldG+DqWDuhNRcnQZDf/ovhbaW2RvStB2pb2GZk/+
0VVm0e5K7JcqCAQEhfSHLphV5otPsSYFt+F6zTKttNauip0iRAmUecT5xfk+aIy8
4deUdqFRFdtWoNHqa9NNZAAvhcYhXKHNV9ZMN37ci+XXhMRFUWG09UR6sIjgVQys
Iu0O5Sm0lhwGNuismXNzecWZnNz9lGKs2A75fqJYDhfH7QK0dj4fc8gee0toin/u
AeK74ToG4FlgZp4hPXjfidcIoO/3QJLfx+kYOBK5b6E34IkR/I+Z5wKvIk3Y0LA6
pshWoMDlZ7xujceYg/gXoNnU9zZ4nyc6P4imUeXgBr6qjA7xGKsZEjCRDVtn/Lpf
OiuCzTyG5w3ogQFNWi8WqkKOS5J2aCKYPln/ygPfOIWzyq6J9XjAB+5//Rz1OINt
QvEHLsUwfSGn83ErOuB0Edq7xcJ5hcEnzmDWuQaLbImD8zjQBkBvUttUiTAzVm/l
rvLgck/QjDqV0ow8q7/sC2eQtI9rK2Ef+58qp7GFTIpwNzZ18YC/kHHJnS8769HJ
MGlKvoQLFnXnnOcWE/l77ZcG7RXusFeIJOO9+70i91KFso2Wbl9x/vhvQYhhnAE2
qvcWzPnS1qPeOU63tfwfWmd2rTCotv7eOOjE58OO6JW6DCegruyP5C9zVnmd1Y7u
dH8nfw4LNTccDHtCpI+GzuNQ+cvbF5qFlc5JlQi3a4mOzwcLSVC6I68dv21Ugm1J
LKQYlaGJkprr9NUep5na4a54QJ+KUFpDhHAqxqOcfHxz06JU3YXmdU6fg8OliGhx
hqFvuengDsju9/A8v2pANga+ZNzYJXGfaw7cgqOAgNLDykppu9JpWG9THdI7teYl
kZx4/ya92KvYoCavb9ddYUA47O6QYY0dwUp83qd92GxEwO97m4Q5QxeoxqLsQgLG
jRd6Okm0RbSHGOScnZAGDAUBy9FYVO9GfnoeuQzM/i1RHqxyp540WCEuSRI4i20/
woj3if5JgIy+5i8eLu8q6SGz+bhy3TjbGRTxMJmOrq5H1eaP1zo42NpO/vPyMIME
IO1FEg6mqph9Qxtaz6oJecvqc2wElxsg3q6uN72K/VmicrxVaEdlWnlueQcA4hyP
9YG37dbOuc49fh4ioIVkHuXxnjMmXoMZgjXHpgMVpNIkUzcpY6hdp/lOjilTzYN5
ELE3aW+a8WcNnv+3nBYhjzmz5nx8oqS7ufAPmwLLOI8mRTFXlctJ/wteVLg7V0Sy
2Yi7wiB9nbY0c1+YlM1BZeNTltw55y7TUqy9ThE0mMt5rnNM+7XX57rFdxiTYOHF
c/Q76J84nSCrrcn1ReA5LYB4jiVry8nxAZgNLcuJzkmJwWH06O94ayigA9qPfM3d
RDFSa6o1tP5icVxEYit1pyGIx4PNa5VP0tE7fDK+XuT9QTguGMBN8e3AfqJVic1N
Wn6w4dVMksezK3oCjwRoE6BYYTm1gmh/qwa6xihhi1A442qfj/SGlyzYyVDI+7pn
Fy/DQr+EPkBcMZyO2c6ClDwdSlJ8C2fV6be/6W6svjRqhrIv8akiTjSSX99l97z6
syHfxkc4UKYX9gF5Xs39lJcv0zm/ZPujH9wEON5Py+vN6sQfATgMQaLHRvQBYECk
R4jdpPvmZbeSYNEe4oAKuc6BP1k90lf2Y7tzRm791w9A3o7Or06cJJAxuNWZhYYd
2M46OOvlM/uJ1qDXVro2OuLeW3k2Bf9g6Q1wfmLHbqeoGd1PHcXM8KSuN1rsGBdo
ayHHeNP8PnL+DRODF8V34xH56FriNDnSVaWbwqCPOPP6S2tH9pQezk2ZPQ76W34O
z0YEMkkH/NurlFalOhffsec/frg2+UgD9VNRYH/UXnVXchzpGmqgGOAf+ZCM0CgT
if/fS/KtOXS8eR56Hkavq64DB0pEIFwsQLyUWJ+2su0oSrjOQ7ui22ZPdpW7x+mI
RIB7bKTKv9yYMNXbGFvN54LJnKxFTvha071E4VtxnL5hvgv+RT2iuhN3dsg85UfN
K5PsIt9VLaAAilB1UoE2eWJUyNebHF5mL7qn3tJ6+5Ra8RM09VR2PpeT6hFaL/uJ
fazwTcxNfVVgOz3XoIQseMjEYikKAK9vdR8HO6QqSJk2Wu5VgJUzYieGQTKh08fr
7AtqFauCX3oix67KZ2ba6R5bV6Jqfrud0sYIvA99gkUXVXA5qpQPn+j8y1hRAWDz
hEaRiIV5hJOe7SN62yf0D00GV5b/XtgEIo3iipWNCvCeE3iXxTGu1DYsut10TtJI
SyCKNY4JheT5CZmoyD5O7svrbnXFEsgO+sZRCACetes1yzUmBNOJo9YMn3IKgX3d
Q/iBOuTpBLi6EzRjyTfg8y6nj5elFB0FnpoZbsGQ1jUpGDaASGczVGl+6rflAIm3
EVUD5aIGHM34HFTTGJ/oCCeI9LHVZxYn0dJ7/mIfMgU2VkVnQAFyHySxdjjgoo6n
samkaUxvH+SNSN10Sf21G2yjGrB26Y/ShW9WksjZyjF3lqvvHhjbhiekfGGCQbzu
NK5KEEyN5hg/wICT1aePhX6AXwADBLq+RdR2ijFTItB16E8pGpv0k+K1zc2yk8rV
4AHcNpTdAXRzZckECSmCD+uUn7Yuk9vx7K7LjIjhfVXQuRx9aqPhW4BOZWxgIX/v
S1+DB8hNuTImCWZ3Y9UAMqaOtwe91VU6kTVlTfBMsHl7oJIrwRK+umeyJiEQyzcx
6HpRExFMDNwiBq+Z4/kDP6nWY3alrlfBCiqG6Mdc6akF99w4ejZC40dGe9wkubtP
Td9es+lpMLC3dFDouq518mgtbpACgPqChX6LuXSPDLzvXOVfv0xpKikNhtHHFpz8
JAo0tW2Q8rymml1gH0V62lQx6gf0awvm1gihFwZIgNudEQKdH2EXbw5syNVwWWRj
nbZwFrzbLLKalOJOVlzCSoOiCvlmVMgDevXfxCInh8Ia15foCsJ5YKuIRR7GD311
oz0+5Wp4cocjFiagGm48+aZi1S9dXqyOtR60cPqwOo5kIQHHFND0prSKA4zoUt2x
ak9lgOdC3aMfcwq6lKEMnRqVogl7D1Fp+eDfeUyPvdIO3IuTArY1+5JEg7QeGC6M
Qrh+qF4ktJh7OUvK48zFHMxHyBiLNEF+PqMx9I+qGMc3p0kq7yR69km1U/jQUDgv
siQdPjHV0yHwa3qjPzgcdLgAmOz7fkkcTgjQr9QOB3pNCVdUFVvhi55nbAau5bKb
aaX0bbkxQyZ4mKPRdH5mJVmjXdEdhge4eIFhffMHGEeoYs3RNMSnOJORagV+0pXu
0QItbUxK7GfKmxsQ7ukmwNczCoYK43zlgle0TW4HB1sletd6x/SKuJd7GYryxZBl
cZesPolKkbGQdshWYsK9vr8MtlVl4qXWY0jp6zEJj5DeP/Jt5FgMyBC+zKTSxjBj
hXBfpa8mLNi+fOb4P/q5ceKIaTVofyUNm9uVb61Xn3I5JcHPS9HmdlpfAzq+IEok
mNTIM3hq+IxI2OhLM1puTn/GGQzJTpHfmCLAah8RAixg7m1nsslkgSKzXgmGRAh0
d2lqeRcOifWxBFNHQdea6f5q+OppVUu2I2etxlnNFqHK5FCAgzwEKHpYrFoun/Qr
RH0e0xqzSP491k6LgZBGiQh6vck3jIpbmGt23ZP7gmxBophi93YjiNcgRt01N/nf
+UUPvwiccLDNqS7iQXmmTl1VLMh1kcihEfgklObawCVvdtRheuD/6Hg7qiOqOb8v
qTubOWWwvyvPb1CjniBP/xpBY+7p1/wTE1KEMnIs+WcLeGQBaEuN9mfaXVXMpfiD
7ZcH1blHw01loGm9hF8+BK6lkEHdfgOS6pCAiVKpcQG8M3vWxethwJ+FBHbCVxnz
mqdRSTfE+ithalXJpLwJJuJewEXAIyNafG/G+UXDOeU7ti5KUyTIYGtwZKtgyVp9
XP3QJD+CXOv4W1u0wAtwWpJcK6tTesGsnKB9m2+PzWm/oeExHEXCTzaQQRaV4Hd8
LxEZyhIhjqpuA8YBchRAMrJPaHl/rQkZjTII9lot3dzsOA0YGVur0Rpmp4uArKCi
yxdAmG9kcTrQlGG//souFTsPs3q+M0L+gG1Uu8xRM1q6H1JvRv6ixur7x2YCPZZQ
917nCZHZBiXZhJ39mD5dyoUXWMdUoT9626aW6fgylAAs1PQnzMsf2L+MrUTvgtYd
uJhXnhTkY9zD0GL/l1U2DrYtildohEwNVliDJ/lkm9YxuWOfUc2VBJ3BTmY8+qop
32VYUvpo4IViw10VvXgOYTJc+/gGxRYbOCGKdppOQzdw3roLTmFQPe/XsYSyW89T
45P9Llb7rrTXC9RmncunKDrgAiQcLxtYQ4HjyFcFPnQKsxtqJhB4MC93h2DKRzar
n1qbQ1JgY7Qvjk0IHy1wVEB9CN+XiW6ya3liM2EGE+OOOl0DbS2bAvBIQXzovkDp
MD9bER+mKayUdvzVIkbJFkMr5F/rcu3vZe090E7VY9BMfHWtViG/lPlwSJGgwjPA
bR8JD8P2azUzQdKSAAoVAKZHm4lM2TcKX9YMAhKf9VfSRR8z44vUEFPuryJ1C2pC
mcCmKyqggPXxofitgw7bsVqS2Ex7H1g9cWU7c5PgvkxxbyyHKfSxS38p8znWUgLJ
xqqpB7gHMVODjWVnJU7gkHp2IO4+egV5x1C75E2NeEf3MP8pcLk3qLQGDyPLBpb2
ETbHdCReHrK3GTTng7Alhs6yccA1XF3RMmmyS9WV67LISDZ9C5rRs+BlR1hNBCPA
HcZgm50Wck0lwAdZFK9QxumnZJ9Oj7phRWOJJPLuE5zQW8GLVBWxgcFbWmKx/nKy
EDxEpDIOLbJTcV8BLMFCqb2T/BuyriYLWU1MElmo1WDhrz40nXqsK9qkW8jNyOBd
iUXpi8E9Kvs1agnR/PGArP6XApcMPeCVEtj2khpkd8bdeq1YoeHcJpLWhr6C3yO4
MMA/j5gHM2Ygnlu8xuk9LNfXUUPo9j0qtTUZAhqcLqsCvBBj/a1DXzjuKkXCTcuW
/Wcm98UAz8pkoEAQfBbp4FFWKB6JSUxHcrMTz1NJSUnb/TDx1Tyy62a2BM3qCged
dzDQXXjY8lSOZTzXC5r8BNFaY3f2EZeKIKwWmFkkghTkct6845vdiv8Vl8LBJiWP
k3Sp7lfm4S6bvGrPCvh+1tGPaBsQjEoz18ytMOAd1kNJ1dsDT+8XGxCReGQVFwNL
7DLsb0ZlgTom4Ho2x+nN+I5TMdKMTHtH1+lXMoHuDbkZf6o/hTu8LZckzXLWLTFg
MvkB7NJv+GMjSnbXxKmxlxlkEMMydq6XR7lL7lMZ3uZ4EbbMZjfebv4GdJvnyRqV
mqhW325ID6enSSm610opU5w3Kn/xwTHgLtFxCo7PzicazDrY9/DXRBKATtbnxdv7
vCDDadtL7ZWOJeBGcsWUr9coUfM+dafxjtAxVWFfXuT8vMG4xqk5x4ChVlLjrmuM
b4gA2aZnX/yXveMZnKYGrpc3CH+IUkMl27xF3eTA/FV7ycPOSMXDL+O48isUSRyC
rOGlK7hVWSvPUW9Fcoi2nAEK38qPY7+Sr+t/sZ1NdV0W8yfHd7Ow2qGGFzE0FDLl
9WxQTbe5VdQJjBYb7LYO/KuyQgCAYT2CZ2S5bKgqZUzjxrS0dysbkyRB0ObfBQi7
47o/ly4zVssVnOAkUlyj/52QbJwA0FrrjvXMMFrrKyQ6BniXriaDFRsSfMBszOKp
bokLzvFUwfLHrg7RBCJueejEVrSYhUS/N4Zdb9GgVeSABPl1dxTJZ+5vDvvwepcX
tO4DPf8CnCRzwHbGUanpf+2GJxVyIE3dEiDBUDa54y50cptchhK6zUfIWDL8IJOh
Hk6mMm2Izo/1L3k4LpzrRaI5g9DCI72H5+9suMEPZvv5Y9flWbc43OnlbGdC+j8G
tlxuPspGbbzoXBPYm5LbNZ32uow7bPuxJpUS6IWNJjhbFv2nhzMqW1KTO7cZWXnY
WpB609nxVTBbpIRrFMkf8VYo+eNQRJxBXOlE8UOYEemXAmpAG6m7rjyleuO29jtt
5r6HZVX+7XMRT1ztWxbyIFJoXpmmfA82wiFohAT/9FyMLzayxQddRNLx37hl62ho
7fdLRuCYf1X42t/BxQHStGPDjrUzmV+ou7OGrqD5x9B1nRd5EpwoCNk1F6IauLva
6dxO6DFw8eDoHF1S3vI6gWHRi0fsd1gQlUdsX5yJ442ec97Op36YH2MNJo+Ik2lf
jqq4DVYVMHwkq7LslP7LEGAq0IWvcNLv/+pcXMigVR9hk6kHXbuwlUNPgNJH9YZ4
FYOtDOoFOyuiEOUNzgaFazr5Bpxj9sZ7n+9out2a3Ppx8WN0iHGgZ7m93QyPAc8I
pMUzTu3ZA1U+w+p0AgdLUNcQL1P+JH6baWHiFTjaLDWWyetiW/40rArox7TGyGQ2
u3ic5GQmgTyb+jkBsXaiubZgdoMB2RfLRlCrMAzYPlXYK6RZhw78BuDwMrDSIMBS
F8PW6dYcOMo3LBWfQOIcfJ5e5omgIbRGI6RL+BC1Bx4z8kAJVCzgCoGSqNX5XPgP
NFB219FHvjI8PC+YIZvxzulfvOZsv78yk9HAVaHCBmw+O1lHCSLCM69RLcoHsgFi
qCaDku4VFKIQ7h0yCUqew36Pam9Xtw4eudwpmpmI2O8X5X0fumjh9MwujcyY2eMn
Z6itHk7a3w7zhkpUJe5oR2uzrTtT0PBS9xPnLZlTpmsliyHBz6wu/qoTjfREP+5v
wRuNgUXUhJpcrzI7kySRReyEWsubHqm/y95t5Sc27dYy4j6olZfslusAA2K/IsQg
KIWZiCXJbbRRhDtwAlNSCEMpO9j7fb0TWzs+f8zQ4i+uv4Uh6sG6+N1cPNif5uyY
r+eF2OCzpJI2zW9BT6vMB+nceb399kK982kdusTLMwYFt6NThnzqqSSPbPzjR8zL
w+3Duqs66C8s2hjGbwf/6E92fJx5Q57NZHaZXiFiCLNTq8WiNp2pnnU9YCkCHGaY
czQtPnHkJ0ydFkYSMR4FVsXUKonDm6dX/nJOd641NyEQc0NzRQD3jo0QPxXRWiGy
oGLv5E56n0DRqgF7qyBloW8N45dmdGfCVMNPx+7uZ/MsY7caBma48rGJOGovZ8EP
YiQQXvgmYvccyLCLX2LtH1CwVdbaa/lrFj+6oWGwC32KdJ95Z5HQkmBSuPrM5+6h
HdmHrsBMPcVcqM0sOOYngiUHciaUc8IlUl49wEVlW/TSCB4VhPwq0YJH5b9il2fr
4ZeIIcu2sKmd/YBlaAvZV7hvR8g38jmpACKdCwCRMSJI1+mk8sE9t7+VEagcMP80
7mbbjCZkQ9lwjikgpGxAamfP3Qa1Gcu9dHb8UbTxnbh87sWSk3LE/M56hlF1rA+s
mz6lcTGN+7pDDYkXC0gz93lp2jWlR6h84FI6YxVJFqKBjBh29NLLqHT4h3QM22Y4
tF6+nAqNsubMDBfcJvBq40iPxbAbPWaKH61qj9cFSaiYjhWZKrzG+rzey8+OYQyR
Sj0zEtulIG6wcYZY8IMhE9iLqR79dV38eyD0YSY01kB9T0mUYNriPv/L0lcVmQCH
DdRIPKgJtzmUkDjsSNh0L7MqIDEz1VOB+06A1whKbd1bBKHwk3VpqrC7eKkdCAlS
6uuDYdLJDGO5pcZkz12MGyL8FfBJRCiFku5iT6ZCw2GhtC8pEEM3pf07N77Z+B7f
VGeFflsTkKUHTnJlkWaVODk0yl4w0owIEezpx5IkpTHJPqyWa2PPiyUAmmPtKhCO
7tfFXkv6ykADMXeR7ROPy0sGOURaTCV55cNSlxyr4uLIgT1l7HYmjRyYud4cfPxQ
kg+hgrlvi7qc96k5SCSanMDu50mOk0V7SSvUeN1AYIkutlUvWLo9xx1IVgUREPGl
Q8uNu3h2UoUHFwT6CvEfCqAmk5w7uOxoWFpwMkdYKYw6epUL/VfrwDkplJKkXI77
VPI21g0V4S5fSPqn59t20O5NIMxpNtbWWkr6rfGd1edN1+ZUUvAr7YaDHrxoeCUD
yl8Q+O7QckTt0mejqP3AlUquf1mAGAQ0n+1vyC5EylUT0CxkCBiOW/bjAzYZE8jX
e3SS/P9PXsnFvp9FM/0fFMcm7A5GdBDwn6Q4sZyl4RTSw9Gxs+1EKnOamx7hoKTA
dvPt3mEyqDaE3uBKPJwgo7gjkqvGwEKx7ak8kA4pz33B74Kz/K61VcOb5NUwEtSV
aSzk7B2w/2VVwXp26oQa5F8Kq4z9EHkXYGLNeukzMMANFSO/VqhyIbqbBYJnkYPl
lUZApKppJJe0Ahlw/qfb6ZE/7/tUYNWFdYiQyx+36comUNMlKv//g9LQvBkgbzVe
avAHSBispMfL2wfJVRISUudm3XaTEN2gibQZLheOTxVPLFAtVlfx+03HjwB7yFY8
7UoJh2G7qZmL02jWbfZyfQHImHrZdhNzTATeeKsCbY31SJPq+XEAqBaNN+HOBfEs
h+9lUXnW/9z9gn6unkzCl8oKH2I6jI3CJ3lFQrFusCMQFCv2GWTZ/MYDAbrDoprQ
2j80YE0WPTLCSkzaoGov1Ls1CsdPvq0Fxj5EeiDuRHODpB14mmdZOLrpGKGCJher
/vzw65GkpykdiGDzP3EllyW1JfhIj5CqCO6+ZkDPG5xH5qvZ/ghbdYgB3z00BY/Y
/2JszUph+lCJLI76ZLXtKFcJY4SP0vgu4bqChRf+e9ZafnFH7rUl03i/cRQyaYCN
fgqYN85gEZutm669tY12F25/fBLu+aLW9zBPwNFtpza7fHoM9j2d5SCXabzGbTbG
l99+RrKSRRPJ0HWMpRAWHI3Y6kyg2/07ZnAS16A4fG8QKYVZOnAu2BFIaXbR1VpN
q/YKB59arD5KSb7G5dahrXe6eHVBH+k6nfIX3ZMi7IQ8AiHxuAaLg2rk5lBcPY5M
XJ5ETDLnAhGA+TfZcrYCUwtU73mUAiXsSBfIhKlTO30VQjVaPinDvLBly8AojQK1
9A/6QxwPfoCinrhPiTJjQRvjF8ngMstX3JjNg7vi950YlvIOQhIxEdzrxN0O4IQN
ri9l4gdbVaBnVAZHnfsPZ4z63M9NTjhLOrw599r+NanaQ7h40tVoQqnfzQvZ9s92
rVIOGyI2OrhGaGxlOVBot3j5aSCWLBHOefWbnWW2C8GxlJpSAuhr7qKSp2e4Jm1z
skciEaNqOV/vgftJ19rW2eBVBuV5vv8wHSowt2TCdtDzOjQ5AqfVCNUrDP4t62IQ
LYD1anZqdrc+WWiBg1kAFbme863ToYFEmVOjsF8n2C/i9G0aNbwOkJzPoi9xunP5
SVje0vAQUHA0tvYIAUDtkMOzm9V/y3eVNyDcn0C3qM7SNNRyr3PXzqV0FL1KL2kd
SgibajsmV+Rq8tPvRajENQXfQsw+XOttpIfr/nr4fDyCzXGiC0AxVjVw0dCi+fXj
xUeeW5VpDaFr3EWnlnvH/X1HVVj5X/c1JxqEZePhVa9QUBlIeIxldN3bX1+A7a5Z
oA9dljPjvwd+z2rXamUO6lrOhqR/yTG3qdDnmd+aGfnnaMhPTzsfNw/LABq0BTIa
Iin8igRY8lMXDAmOWoqHWhIyn4HtUK/4gZJFz9YemRKlV7hBGh6ljxQ73adjsb8H
X11o+JKSv2z4VJupyyWEkh6fwbTXal2b2O2pKgBx5ens4vG+KvJB7ldGcbHguF6+
awwj+xFqrPxnqr5rxc1foXWBCBVJhSz5dJV8ES61iNijwSaqaFsrz2ioLcstUBs9
rpVtTUT4odsKdteZXXNiXcIS2ktq895aok7j0i2necwmVQTuBbZy+Ouh042AEIs6
cmV74gJ7mCAJKzcLWu3LcvNZGkIpzsqa+6GJrVqR8fysrtRhCmndil8r30yTkbPI
HPpFnlAkW7gjK3AX1fcuFc8VV1+xRuF84bYK6vAHJAhKxVl8K2+qDr8zwY7Wh7aZ
YWIZeo/09Vc/i1K3VBqKBwhmx+Rs6f0c9HqfbG3SakXkmnEfOYR1fRq6XycPVt7V
5M3BNknHw2u+kp4KzcBJRSZF3FbmDQTA3K99lMtMpN3puCZo7WrcScbt9nUCRbfS
XqdkQ+v5ikZy9QaVciq5XM1WuGO0Z309r3RKkigak5Qu/LjIrwgCRckJwoIP9KfG
cbjYUqcQtVZ9OHkXvM16kneIUCcee3N15s1PfzfgzC6ZBRUgvf3WHjRfL8ibZPvz
IIDEGrymeZr11MdzoG8YRZl+NTaIQENJCcLCS6kMr6bjaMNmbSl2/2m4rzCKCuQJ
PpryeiU2CoUyVJt+E+dXT0Qf9hUd8McVv0LgRcLWQ2NHezvknpdLm6bAuOhiQAfq
Q3vDDGm8dwVqbJI404L5b59Yn6ZoZGnH2kzOrmmJCC3FowDpdrjvYJnTR85IbPM7
IWEcXtfifmTu0A7bFIYvNYCU0uYtFaP4FCrLXWBjKAQhMkcZuM2I1rCgyYTQzdTZ
AVaE57XiNZlxNmxKPM13NHa53ApteRGfwZVH0qC6+i64zlwd1N3FXDQj6zkJEYDI
mOjO/Al+VmZWMPXdSeAwR+31uRxOIzWDZFGj/F1Nut7pcwDHniBcITwMKjH+8DqF
euuyEtBaLrEbJNO7K7SmqxFrNMsWY2W2fXnF2IFcu97eZM8GD7V/7uQOAuuJFz5C
t/Wlvxy/7F9KR1JSpZjnEFh2XI70ybPJpRoqpGC6xwwS9uhALSIn23k0uyQwyf86
Qju9TWJuUCaLv0Anit4Xm7jUY/fRN0WA587Fz6PMDnsYXuKiLiLyjOTxr4rNEvI1
WhRIFbd5iDQvDClrQCfzdnn8enT3gnDyL6Uhir1dMRZDFTwX9Srdnh0GfAtfm7/F
JauJs80xzfVQkmU+u5K4RkKV08RFsaJf4M66ZoHaSiycmVvSjng7e1X5FZ0flp7h
DCpOxePVWYfnnjVObLSwS5FnJ3nvuf5JsXVh2LRv245NDQvwfY7BHw4V+1bd+lHy
a2GA1iC/fe3UwJg7MjlTkyNQ//G9g931HlHG54Ha4739R6g6mHVhlX0cJwVIfW20
VRSFzlemUhThl9FpDY+q+GtcFS3wwq9K5QfjslqkgpjM6o0Zohf+ZRlgQrUS+O5H
AFztPlTomQ1XcbD51bZqdvpLRj95KpjbYianZrWdrMdO2jWjbOQZ1AGMDI8GQpP2
j4FDpihPIEKtHJ3SHxH1hvG1ufVosUREFmshqL0nlM75xMBM2pYktVvMz5zbWwbx
f1f9dmfTdzE+ePFfuuSz8NoGgk7K5bNb/cDJW9xXhoSE4gDhVh31YW2bRGqOMA9q
+ZEwnecGAzZ3cZd91rZwxJ9S28lN8jd1vixZlvE5Jk5tAy6iam4nPQCjIyMHCxvo
0nuXjYmgQ1bbjXVnmdNlr5qFqHRUaLi+myuZLXFfvoQlkEcCpJ24/6lOzoEXooA2
eRmz3Ps9bpkv19uOPkMkBXwYyCKuscUooE8mf4UT7gmh4XM7IRWWydcjveJEEIMF
tnxQqzpZpjxNf8eR4waZERdGGZdcOl8jl+LQxgP1GMK2kY7OcDUI7huetdZrEkc8
4MGe/+GwUkXxoZ2xxwoNrWa98mpSrAjfDgT2OmXUD4us2zUW06a3AgqcIBCCWTU2
gspfBEMHXjUQH9g3N+SwOd4bueC9l8MzI5SeCwR9HGl6KQPx2zFzmWxI0ogKJapT
V08PM1iG4WWGnmSink96DFx90WDe623EKun9s7qAdGnijDtxHKm0HZzD4I2spULG
PQlm4QuuskRynbl9y4Pd0+ucJU4Kv4vC2xyFoccfFLgkV8xKB5g6zDs/8Jxrd/tE
dEmWU39pAMi4gZKbISrWUO5/G9kjLusZ3+NGb++q/pma1TWWEM7G74/AMUx3tWi7
cOLVseE7ZpeenptIaZiQFyRJihD04UsDE51BVp8pablLlq6UE2uc7OztUsME5q/p
E+y95hOASGe+5dOlD4Qgm4S5oms5rMfkeLp+5r0AxFpzumqSo179FrR853bkSYs3
YzS36oHpJaZVq1/sjd43b3cDnsub9CyBuzZV/A7lFCWOMSHjmK3Jd9cQ5NWXUKk/
9JDHQrG/JMcEDh/39dNIuc0E0OBE+8gwWuj7sEauzyQYslg9JTf3nt5foPYd5+dK
8Alvvp/RWQm+xQGQpXhSsJTvJM+zHXviUAZRDZboHRULbp3hlQLFTd6Q4COUyQYI
1Ocg4PQz2oB4YQ2AY0CAOyrkPZu74GuVWbmzytcdvTkrgpPCs+cKwwf4q8VZPTqN
COM0UKqjEVXkhNwsTFecObA5ZM4u0L3Of2bsQNyG0DN+lOKgV85ZNQVWbt4nwGa5
ae393m0/7C8tP5ONByMPvr+AYwA6GsgwtLeDEE945szYFF311wYn0ZCSyyqPm/GI
fnKj1XQT1bHl5R0h6aveAYG1/od4tT+e8Tn5Q3uHvS+pj+N+3q8UYit07yOZCfug
1Ye8+mz3go0CbVrS0BwGcoxW584bZpmiUPUTpW9dNY2IF89Qj0YRcIy1Rr2/hHJL
Sua9woX0uujONXng+nag/nLm/XtngKXn+mPVHWJ4MlO3whZPQjjVvf8ghPlKB5H6
/Rzt7S155+iF4TODKMTr/VBsQYgzVkuChSodEOKZIxmCLK6d+9Lt7fBOEBfn0BVS
7yKXnqEwG/RDi4KgACkglg9anic+4rt4QKsn9yN6dhXYQta5BTpkUWKQzNAAEpi7
Dm15F3yWxz56UIetCm7opn7LscoEZ2xSYQJT2jSRXAP1M6eiuDvMnTuB64hmDIbI
5GS9VycuRLIZOBhdry/DM4A8TbDLGsGCA3F4TB7hoqKkQiW76TBAssi7P/9er/j3
EwY7B8DkRZL16oZozdZENQBN/KSo7Y9eT6hizGkroJseraRRYSJ8hPgoz43uYoXj
8964LxCR4HgeTLMBQ6qFKQeTj4G5yQGAJDAz9Ymu6aD7lhFzpfrdgKcdZYLSVw3y
h2SicrswF/fYn+ZOPJfOEjyMLk0UMb1C2VPAia59GL8eTojdoXv1ysfe8Koc/Dkc
DNWhv4Z2NoivdGczYBv8Ve0FyqXNiCQU+UHOauJEyEgHmX1j8dKngYhB8UCh6t70
bDTRvuUHE+auj2fX3J2VGyghKiaNI+Y+pk9cBngRb2x5gOx1FEnq99XzwsgWkDE0
e86HM7NYuofOtGeWGEotwbOWuM1AtNn3pG8Ql+Pe9z97BddmDNn4kPeGOGLkFYeY
WqfkNictSclzgItmrCvB6dM1USNIaQthW/VeYC7oe7BkSRICrmILORWmAJj8QDzy
KN1U+uozwKrCPtcqvipsByXXxbhT36/9ugdbTUXExzn6QnJ9x7IrQ9io17xDZOuP
gAsqJCA1e9MiPFJEJKrM0PGqWCQM55u/+qLfdm357xILBog6e0th+8F6iHX+VPqK
MzNfyDVZIlruDqarIdt/cimNIFbC3CwHRx1ColDGv9CywzN4FF1dcwiCdoxjiYf9
A15tDxbWQ+od7kAIFiLcJpTDGVVtS94rYeVWTORx5MgqZVoVonve/yXh/3fAnyQ1
PcPNINkV7KbicJutdCDjmRtsoh64gv5jhXaqPScysIpKZFzRCVHZ3f/u/3EpdQY5
JTM4ysluNVAAfPaUWHqpf/gmxvUz+3ledlfJWM9KJ5LzNiPwy8NMAjEF0fXvUuvZ
GatkBddT5hZWN/xnFTabxQL9y3Gsk/HB9+bi0WNL9eYgk5R3CX4bWZR5Ir2l2Aj3
u+hd8CFzFZSExxKQwwGuWkizXIh5bj22Nmr9pBNHWeR+n8t+5n2HYZx6tSDIHtg6
j4WyW0XPv+FLKG1rkCL7xL7Farq+hzf88yieTMgJTyY0WFPVOWj30TuVq5awIlWr
KoQry33cviBU9StWq2N42kBEprFLcQ3nBxK05yQyIXwOfOvVpCsKTegZZ+T3N5LB
jlKaErxbHn84DXvkGU1kFnU1Lano/uIlhkB5FKKjwXIEfR3Go2au/5LNX9Y277Vh
bu/fbVOYBKjRM+1HeILdZWo+7nTlitRLQrvoIiiQZA+CC2dwYszGASBpIPsn/nRm
ZJeGBdLvoCKdZaPNJIACQaEuFrPNZC492lIuEWJfLWjR/PgPSrwSTt89E33hE6Ev
bFnv95FITxMHPr+oj21hA0dLiMkbnrGVAFqpiLaknN7xiZva+f87i0x1R0m7ElkE
/bhnYQdQZEJtDNJ7BjX6zq7EE6QtugRt6rP+zagU4k4ErU9f8T3saYPnsnkYR3MY
eYiGTHn6BZOQcNHZQXqPT/GhfMZDUH84+p1tUIRvKt8yBIBAwFqom2IcRaREEx4B
FOyaDId/cnvVBln9r67D3S+e9eEtFdRYKmYmkwzpY5hkK7D8S7+SYxIeuKPUBVKy
9dtt9zkEw3PNqcU7kqrx4i8kFyFrYgO3az5iycKhXqUwIML3icwcOp775R9NdIaL
Orz8lzVKPlN6L4kQ3xobncmudOajHcLAC9fSQTN0nqKMBUR6A4PsRp4Ez9RdPab7
eA4V4Vh7yxHODxqVZTxiB44fKpQHr3eXJbWtWMa+mDZ1jZla9LohIXjEjfdydUGL
rXq5NW6npw/QOUGXINg1xoDIPNah904HMLJbpltJWP9/uPfwDWB/uFdIH3yDhPCZ
BIqj2ASaQa6TebH94KDYJ3AUnGWm4ctesJUE8LEwJMgSXM39mWwqq8MBj8+tfWwj
Di3Q1oaxNVd1gkIXuxKx4YNGd0jIqLRIEMTSNQpC9ZtP1XJylmN8TgE1lKG7q7Vn
hMqteMZUJe+W6SWiGURs/BzRFrQM4kAv0BzSkDste7FDB00cyWZfM+lqmvNOSb2L
6Ax+cBB7ezmm6o1MD/RJTdJd5IEfD/93U+j9OdPOXYDkhMIGzCgqP08tEOpOMXD9
kjG+bwK2qE4acldD99jnlMQC5wQ5wtHkXxwCNL0Et0F6wFhpm3inG6wvGMSzXroR
J9K5DRQy8K47uss3jfVxl7hoxOlZskimVb98PN5UQZXM2gipsh5UO0p58fgU4Dtz
t1I5uFEoEjnizTPjE48/b2Dshy58z68ABvUVmOKhzXdktL07DDdNIx8HbSy9UxTK
KktFpP3R0bLvDAAjbFbNF94hs+OzaiQ+HLO5F8e8a+JCCG3t1B4FuuNhWVsXPF/9
seLDy2vfj1SnMFdRMjFT/DAjSvithQde08nOh+schXyiOg/Lgts5qsEgJ+PQ4oYq
V1iLPOMJbev6Ibr/pwwZ/TiOk9z2UeiL1Z/SyE875n1wS+oy8CW4mWX9gAjKCAU3
SQrTHlMTk7CJiMfgtkqtumlHBJl7mLnoBK2XhhLTFrVA+ptR0myhsDPv68A18SeF
MgtWlYXnVvFENYNGgC4AxZz9LdzFND9a/z1iloEKAH/3nS78BVDkJChneJVTSgHr
Q4oOk5Hzkt+946PVJOkSUkZjt0Az/Uo+Pw3QbDA9oSSPZhc42vyMgYAbcXGg0bwr
XkJS49xeZa7yzpeBWmoCTP13KmFXKJrtFFxuSVIkbszk+3eyjCo6gq0CoHfDDBJL
MtT1O/I+pDwWrZcnhrbhvgviaIGNMWlPsEXqwvSvxwn+eRyaQhPBev3zLXBkT5RG
JQCV5oDDMGQ+Zdp5P8mv8T8ZuGn12tg8lfhu3tX1P8Rqy/IPzImvuHqZNgrWYics
VA8hLJHqKpU6VxwRacSW2/XBzFK8oU3lf0+23Sm9QiTH+YQz+uK28KG2A5jVzCyu
K4R8Oo5QUfNHeLB1bj0yHuyYVTW67Hpv/ahfGSsvG2JzNO4i3ZQdXnBUYrwpbJ5u
ejvkgaGIhxFN1jIIk+fSI/fRGLcq11DvT5qwRtATqbHXMYrOFwolOG1zZFMfdS+/
Muw6ZZVKriQqfWuKJMcYXAbJanufg6moyYpoKED+hLBY4VN2s8wW5L94ITA5CAox
RqRF6gOGQ6lAK1iJbO4mhU7BhUhi6ENY6TfwtxroRbHeVRDiUN+R98ReKibojMoc
pE1a3CUCv8Hzm1XY2rn9WIpH5U3+kUN0depxYLoGEJy7e7N3YNWZ6d+HihT1Wugu
xUShtQUhF8DYGgItDhC1n3UkSOUnv9EFbdi+JaYzvRiziaLpoU1OaByxGK4sPnA6
LkJlXXCLq2HiOcaWB/PVmIhgH4g7kpJJk33FXUznl+cE5YY60OwrOpBv1+C/nJ5G
KWUUvbOKzxZxXAtzBdWufCdK51PpxidIBrjn3+RfBesj5f0TDfjKJ72f4VvxITAg
ihQPkFOcJSw/981mr9JIkni8os9YMfpCYb5AnCzIRiy0IwSCHljZr3ny9BEb9I5Y
DUk8HAZn1HVsuq4hYZ0LHsgoEqjKZX/5ezCa1quI+ta4Vi9TY8x3eyOZXCCsIOtN
OfmJFLJV8D+iyD6eTNHRpmHwyjVXJB55bWWF+f1nM5lWAQj1yjg9GRZyFTWHKOyH
PIDyyMcoRC/oPV8K8Laj7RO0u/oCILmjO26cpHCEv74I/SeCGe5WmacNxm8FXyy2
zHAfVc2bsJg1P8GINNWTDAcEygxTPfmu0oJpGBWmmcSEGEROMb5THvb4AKSNogrQ
m3NHr7jaDerwBIyr3XkRWUSP4ToLi2fN+XAO/j0KkwmtWEvkGR7T/7mPzH3CCLTl
D9eEYZoVJDGWuaZTKqlXIGscIwcYpppTULGZPkfEAItKCPXkAnrWqVIdim13aVu/
O5RTfDMjjQXE4BTIyfVYYNE4kRYpjyNWLeu6Fj7u/LhqEC3CG43zHhwDucVPW69j
fPobxD8U2AHzgIzG8I8XS4Tmtdo2AlRFBCsb7LTMBNg/fAzOsFy8aZeaIKuKoTNx
o0T8STVgZ6QaOWmsEqk934m5Rz7WdrWxFfInL0ilrVCM9aJz9BymHBOibyNvHJzH
OKOOJ+/6BRD+HogAS4i3t9CluChGzRfW8KVx3tN3DSLRQt6QBM68HQ+zn1UfiSnh
FUR5lnYgr+mhafISm658Ri/GF6mm1w+ePn8chNdv8JJlujQWZqLWvqxl5dlsz1eY
+TzndD1haYPNQ4KROwVFYekou9VVIOTzdPtXKCj7PBUO/X3HwaR2pnLlmzFExMLS
vzZ8JKCXZgIrY1jdtLjdnN8zFWGzC21Vs4a8UEu9T9VaJnRcyFrX0G1/owD6Ta+3
N1EVVugdq9XfAduniej5cx6tdyOAaOu/tVRYMWXKWREPWhEY5T73OdBS7CwVp5qh
UXIojbDmOXlTY4jawToLh7gar7KeGRqSX5MCQZpDvf+GG4/ZpFmbUVdGrVKxvu6H
psSfpobFEUByEAEQ6S0fCdfXi2+0T/ejyVwtFFUiJmReu/xvTYGv7DNZnRj9RcYd
iumhYFg8Huj6PnPaX5SYL+/dqi/eeExbgNg1ffKXewlbSs4Udj+/FHAc+KfgPr7q
dz7+4kzLtJSdjaaSBhz52U22wD2HNyel8VdcHg3dVrTS/0KK83zaBiDHqLV4TSv0
lbBYQuC9SCrd8e2n+fMfvSzMeISo/uW3Ixaw2GFEmBbqW+mXI/tE9Yvc8t3TKWZn
7puU5ryA6ebHazrUSiOQCHf8cDCi/f7DZLx7fZgFmGYBt/5NxwDA00kI4XvbKhr3
NZ8iLkk9KVSV28/zgjT/4Dv+vmWjUtLVyHEvgWh7o/Cc3+/ZFaOmmyUwnagDCCba
HsXTLLb2dBYg+PjKW80aoS+F4xbqx58RBT429jlBeejFU8e8j00/uQnFo+kV2Y8T
Gt0f2Zt49LAFH3iT+ZShxSzk3mfkMOYA+/WffcKu6uIQRASNYAly9yGs4/ka/nWn
chOkiW/18VaojN6LzqgP0AdsRp2w3AC/gTJWatdKWvSncbfK7eVJixmldsyI+/+f
BSJxH21QknkFuGMX5tKStZWh1EugwZ5X0nZGBb2gP4c9fz+beamYtLZCF1J1YVyp
HbPyaXQ0p7Medre1acqirhNqK5SDKwmz1RZ++BhP1/vyekPDMhGUBi3GLc4FSh3J
wGk2dwtwBdxb+7e5kCt5cTbVeTHy4JtbJtFeFjMt9VQtnfNVVZwP2z8XIeRT0DDJ
2OAGc9em3reLgutfetaFqTJx8rLfE/A8iw2PzDpUrp/l/EmOqD/O+bQFyr2vzcHg
KiNALtWk7ALP0NLioeVGjdrjijoiqFWPcHIsJg74nLB5RINUWu8ojqiV7TOjAl4q
7gDJDCEQEVZOnQO1BFrTp7HtGWcZWt6BhwPMNkKDcfnu7RSq5dN1c6x0KwDaRkHP
709CNSav1/rjkTS0ng4ZXBurMx6p0rMsAmJUo75LqOJAHIAw7iBngim3q5i+lCY9
aORogvYfTtRbsVJIalgWv6dvDR3gBmD3jLwiG6MSCpgvKabsuFJN1XL0paSOeB/L
z2LZ9mc7TKBUBkWLueP4rpzk+zMdvuCt9kvqFOVOO5NITlI5d9mJEZwzzQYAEjwZ
M6N7L18N2inxije86BQIMYpg5as+/Av/62icZob7CP5Qjmi5C/10ZWevGH1PZ1k8
5T5PyHlu9pj+UBwwC2jRDCzKLsDefbnpoqubCmGR/hjC4NQa1UwaQt2mPuTVPA8c
shaxF1gyjsSQWfmAwOlcDv+QdoBRU6vkvXdJZeCgJN/ug5Ak81CvkcvGb0RzM4jc
eYaG+cZudsT8Ieca2xV7cyFuyNynR9/NZ612E6sIBxE2gZ3HgIWFilKLzlTnCkI/
TK2N7EfruycxtI1cXiJvQR/TiyuPA5PHOjRlii/WzgmYTHs4mmd3xv2Wpf2O+6YZ
/lKCVIJbBKPGE1GbhIdKson+sKUEFF8iaVlRHICxp88Y9eSiMVv0UtvgcpSCT/mZ
lvGxUi91CkA/9KS1OcDQWK9AUvWVUEQ2AgBkBHYeT3oTA20OH9wKYqCL7aOf4QwJ
48ABoqIDnhI0r8eemA3jmyxahCkDDn13ziyy0a64hggTSXN0DO9QfkjxAyrWTJ6I
li37OvvC5RGgEZUcr6z03/R63ET0VGeMf1Q/LA6vlplhcv05ZjaMIWHCfFWU8tEP
ojhRX4ZIIz6UF+Nbyo5F3F7Fw65lzbrUAbmqKYR2Wd4VMJLVKqS6OIGEHPO6J8oX
SRxr7Kdq0TVNpA20YTvE5X9q/nbfKmEsi2tzvCmdgmKvKp8dCLi96S3TPIYygBav
rkKt90phiAH5zvexNXbaCYT07uQem69xi7hG1WfV94DoReDu11WoG9XM9FapV/NE
6BwsYkrzHt/lOF8yMa2uCYfX3v8U5azUa/tJIdaDItStKBe9k4KQVsKJf+9G2FkW
zE7movqyHHaNgI6RAX1u4bVO4PrkHSJB/Av5XUL2JGvPoDUO86rtWN8SKkjzGsyz
aEGfbBhmHs0Y4O2oDhOkBsImglfYmdtYp4PJYbI0Q0Wr53uwo538v67sirZZFYtI
nrrTZn3sJJpgp1zt5FOJnWG81AyOJJkJZJSu4DdriBdyQjC02bsqWFdDEd7xpxdz
As90WwuTU2Z8dhCZRMK+DsSNYhiqKi43y+Be/NyRlItx6uTYhjFZ9Ik/Ykxv1mJl
Hda2fc/43/rYOGUXOzZmId/pZ0o3u/xDweDPMNZvt7WMDcLcSgkO5lQ++wNjkkeP
Gb8xH0vPu/W93BpFjgB9+HomLzG91cfM7kexmLsPULBZyi1ee6T0+RWFod2SWcyN
bvFIUMUqNkgr09x/qTTdKPS3eM7C9FnsUKwAqL8FyzSm2ap+YVGhhCk7pU3CmblP
y5/bsW+Bbg3XQ59m/nvkmISXWoK1N2Lis8zTyVkKaZabRepdEvVxF4NPj3cbAk85
xzqStEF8n8ZOt6WNVix+vu2imjmOkVI9Zv95Vek2mra1w3m/yh1HFsjthqq7RyGr
09MV3G7U1vc90lT4jz0dV4eu7MKQRBFDMaRqmJnJbjhxyNeRnZ5IrAK8xbFeaOZ4
x/qnh6oIDtZslXeFTZJ6FjzKS7X6PQEIfijkGcmCyWIVmNvUTx5xCYU8D45nSgqu
h8acHkunSgCjlMu/sqPftyjpLRVaB0JX3eRceWwLTmePZAcS+UdqBFYqvF6xJ87L
BxNgKNREiCHWr9lETQJWpe2iU0U9JQYDzUF6yRaapdTdFBwAZoJuZTPAJCKcchsi
moymWez4WzCsA4XQOFMqzXM8W8rZYzfrNEEA+2x/jCM8iWlcYrgt8POyDhbl1q5k
cTLtAEuqftHB21CuZgxWPLQCWB2AMTXIRo84QdzaF/MJcgDsD91YnV34zMSh2Deh
uVKoplt3DhyOrzS5qqifEYsR53kcQOS/1iNVRW+/7cRjW0wCM3b9b5Mky/ZyZyLU
gtv7zoYZWSe+cgJTzJ/3kJlfVFRiCUSib1IhyOGo++VoXCH/tKxCOxZzSUvZkOHI
gNEg/Nypx6HsmyHlpy3XHHsDkLALNTZ2lMabwsHGOrdFfDez09e11x6GQQjnMXdi
nV/9E/zTJDvbETIzmrdxQoePla0nFkLj5KbtsAy7ADu1yjbsvrkG4ZIQ3AgBAQCB
u4dRI5iGrv1El8z86gf0582EnHSCuWZ/Ih1y2CU2GWqkJV6iY0FOc2543Q5LeKBE
SPRxMh6hIzDC3GUFBdtCBXBxmQUImvfvhqabn5nhIk1UyHK/y5UwyX+6Fd6q6mqJ
8f8aZ7ZGsQONvjXFTMzHgygvi0WmXxsX6Ta7q9/RnFNgNbEnVPpjJBjHMgSOhyis
vhHtswjRCWBmCkNhKX8HVSJjMwAXRcs4lLm53fZIeNfX+sNFA65gADj0LdWMU4TR
Ea6nD1Zn3HBC2brfdggFT6V8XJiXZDRklhiAZVfw6TwfTzy/fL0zdz8lSKjb5uCk
DVOzyautQ/UnYq/XeySwAAA8hSiD0ey0D3/nY4f1q0lPUQduQva3K54pGW4A3XEr
rZli1neV81DTZF16aCodKl6z9BQt0tLIcE795RmBZAY2oLwv5Jaq8cTvQJaTvdmj
COfFZfh1FIO+QHF7eHTkHfj2HsCcZmERRUvyzsSHu76uI/K6mV1nStT69HZ55XO2
mmGb9BHnb6W/ERD83KGWHLBHKKDOhE7QO7yiIWZANxuCv1g9ksn4EEquS7Dzn/zy
f9+kr/OTDBtJXlGUK3ae8eRfKQF2hi2ZUZD3rzDTHBiPrJWmXU5Orwp41cTr7p7x
+tN/pxJyQuBrI3HoRE98Y5A6IpgH71v40F15UuXBzOceMBnURy1nVUEKqOuMQBDQ
WnnPmMbGVozeDbbBETM5QNPugLugETVyOmmmQqMa669lr5eq5ec51fvFY9oMso5C
N3PtYJgtyVRzfI/txkGDxuypYhYzpkSeK8N3M+9pOcvQMjxJp3S+FZrKT7pegRKE
vHLs4tVID312I6rdu2pDv13cJJw6npfPsatrqRwY+HlK6FPEJTwDbxTKTn3GhmPL
6qptSWvR/7XL15be5LIbpjli/Sbf4V88BNdgf8OstirsJgwVDelhQPHrURdV1sY1
KXOUrLQHrukidOmA6t0rksMFpoEku50Uom628mc0waHT5+hCOk6DisDr2QofEjOE
hevP2C+iNCDA6sCLCKH53UIocf4VBO9Dq1/cx6paPhYldl5/gXFcae1HLi9hTq02
5WzsWBQh5Y5NoDlLTJbM19HpBxKFs6fkcEi6P+0vqQ/8YtPQEIRfb11I0Ojmt9t4
bmrZ5nLnW1qLANLbQf18xYA5IHT+bnJvSsAIzmty19yf51cYtNJkmRgH3nRZF+kz
gRLqI1uvo0l2Z+kIKgf0d+MUgAwqX1Kkmi0yZCxaLiU9ofK2viyOF4pTUaMl3l2b
IjFxAfL8DlnzOLLoDVKRGFfYEdussPmEa6/3COb3fpjN6AgDIQUWbjiESJkg39XJ
gjp7cIt0trPvKkn4UFmoW5s95vX2JrdgHCL7/psSBO0e9AfMOieyMjH3q/RrSVvQ
RtdM972NykitvTby4SMJQwC4iHkTeMLNV+QMtQkNfi8Akd1L0MP1+rWFvmkdm2AI
Sj2L1yD7+KpXW/wsAxHcYR5bGGHOpQv4mDFpWKtViSir2tJlDah94qK71tmZNIny
/ZMhSTYYoasUO4RtimBU+w7vrQtCJxeUZtwCu4CxHkHZRSS9xZoTXcxz4Qk8RmN3
saEBLa1iwJDArAoMVyItS32ywpKi4ZuYQWyf0w+k7sn/HJeefKip5BEyZ0fP0I4q
cB29FtsRGb6EBzsRSJnIR0m38xPjy34h8foWTT4dTUiAZ23r2/QbEIbs2nmO8A+i
2JhBjFyIgPYoax8S/M8XSexDUTTrBb61tscvD13MvLNfQ2gYUkz36olFZS3lmO39
zJa46Qpcyy0N5Fi+hACxsB2G3oy3Z5ZtewhT/tRXyLLPGrqY9u1VE6Gj+ZppUL1N
Ahq5tx3ird65BlT4rYp8Xnulu33GGXqKwUgTiCRlbeXhu9Jq6orR63xCHO11eUpX
BAry0lS8PJh+PIpXJw+Jkmm75gFBC/rePsr+ZHwkI9qUSjgsLkIXTo2IK5ZowiBW
lOzL56ie+wpuq8IAX7b/gFHM6i+5RtTwkwSQtfSch2hebANaRVQ7ksVl8zGXv7yd
4MnzclrM30ZVngGQAgESYYhBOPXiX9qoDp9kBVG5FXt3LKgQM5FanAWdbKI5URhw
YO4D8h4IV78ecflDBNX9iZYds0oLvPCcP2OXaSbAcNCTU0iEgK9pJBT0+s4q/Okv
70IJlqSgsJLbOqiE+F7mR2ct0WEy6+qxZx/zOOMhLVYyLwoDiM9PV0ofxsSeRIN8
DYT/4ROwPNkFv0RvHfjZw/ZVF59//ghdFBFTrGyq/Dy0X+RUlOyes+ZFDRRbOKLC
BvCaOmHgvJ2jylZJmJV2mJaAeaFGTTYRNlHpVraNmLSLOEN/NiHjN/2KSqIU1iJV
4SJTYwqqE2rOjRX/7QCsdZCYEDP1CJMt69cLGLfT4SXk3S1StGQmjB0lJcjkfZC7
7aicMSmZW5Vh7Pa+9Z/HER1nMbIoYcnGVhXQYtFLm23I/CdIrxktGNO9DdB8CGmW
FeXr6RFVYA83hlUbCHzyrNwZroSKKwIbNt/WVyHXzGzplmD2Lh64Cy5zTbz3M5ed
fYTMkUPBafKZD/NdcMRyI62IMyJjSuhPfg9HWT/58TGo2SsxBAGWINbhPYYELnPr
pOxj8gvl4KROoObDiDKza8xhrN7upveekPM5chw1q/8rbG1r8Ctzjj8HMFqDRv/F
VjcsNUNBXpj/G3udrqheaduHNi3dW/n8qICDtJWtBTyiX+0sVwS73ZDiqaqskNnk
N7i3SfCxpOZ12f0x8kYnXqnJeLdIiRjuZPFqWswAWHrSGD6Lh8NvhwU+zjWrlcBX
DK7OBCEalf2EAvD0uhnIZdeTLOKtMq+Ii38HzGRE5oRJcWxz76Hjvdtc5x/RnMkU
viaDznQ9aURvevZhdBpql9bZ82sNOyyMnl2Q0czc77GQ2qm4h5jHIl3attmFg2a3
i/deiEeBe3pre9eYR2Ci93IjMYMPdGonuR5NWuwYWO7CPpEKNnIopEKyZYx1eE7H
6uhoy2ZHnqYmM/IsGNsDHc4001nRMXfHaMg43WBFkfld76ElyR1SHVshS1ThRwY5
Sf+P8gV6R5uQY4t2p6G0qVxQGWXEowNPasxV7payG8gXsGj8h33CFo2Qy4q2D2wu
fgmo40ko0EaPJmvL3gnh+jReh9tyQgktXu/trfb1fBmthGwToZxZJejNm+h0TlQs
ibcsIDB6QrmR+qUogsK35mVMd6Vxwj11QTCazHnKyqmpQ4lAxL1pK6wyNN9rsrgO
jhKI8yMyyfNnCsXP41tuvji8k+hL7NWQIHheDdTQYZOhY/eHMzEBTQ5oZe4FXOM2
ttUleOrRuBhrWeYLfneYzyApwkcOwGE/D0TggoVOiJOrxmizee4CrLD5nw+yTqdB
vWfkakGlBs/wOuhpsFGe6EwUzizgEUiW2Ph5kg1ZPstROPppNzJEF3OLeNVqecrn
uLIm7aAy4Z3sK4idMicoORffawfis6wJoAlf35Aw+v16pieNW8NaVChsDWDMPJ2Z
DAoI2ALRWt1uHLPPE/cmY7RXLQHCT+0ilsyPB6gJ84aM/ETVZefmBmB2g8kc2jlN
ar7FNDrVTXucSbjar5itTW10cBjIH+t2CxMLbdS+e4NfJ+anyTmOt2dGEEjXjGSt
zRrO5thbcdIgjg6aruH68BDJUmrj9/a3kgUXmFcQ9n+5/b/t/0SGT4u5C9r5l6Sc
5IxrrJBYtxj6zrQFAwPywWqivSDrIdqgPvd2UaBG6mHk+G1afXtHMf8Z6zMEZMIM
aoMmzkgpQVVZyXUb9gpnCEHticYoXQvYLnPvjsmeSD/y4OriUJIEK5kh48CFFqQE
17irRhjPQj/HMxagER7vynAJdjCWuwJ/bWSDdvSPq8RuYI89MQI4VRAxfYGNVssD
e++lfPmIK9enlmjwBm1dwniBe6gJK5ur1fV4+FK08wLKqe5vH2G7nnrXLhTFnd21
iaJzLKgOYvkSZXPIKh6dXn6rwoIHfjETk2rZFs3ar3pCEMMQw0gPBPXnEvUzzbJS
JBi1txI18QHlRWn9xbY7K4sA8n8cBxk5R8pyYcJv170ruEr7yyKgBOmtF2f1IIEn
ta7yRPy/89h6P6SO0sXCukTXIqgq9sntO626M9fzaftUVidjfu7VnpzYsGUKNkFL
TFsNf4X1VGaFmhNvX2CStVyjDyc9AFEK8tlkiyqOrofmjTlJ3lfKFzhopq4OA0m0
ie+xZHx1CLT4+QUZBwIiQLRC7aomgiQ1i3tFWKxfOLDUnPL0J1axvTJ4mxZcIIwX
LykV7sqkbfpDfKYzSiYpHugRm7f+4Xok2h6M37pc7Hd7L4KmneUqQDJKGNEJSSuD
K9T66o0eNkASrpECARmbajvy1KUSXeoK5ZpIRfDavQWX0GIOb5oZ25KbWq+77RG+
LgAvandOWcGl/ZIso0e/fv1LK0Va6lihetOPZzRhB5NcuyPeOsdT/MIGrzVYjquR
UyqTbK0pYwcIrsD50H85NNqgcvDrrim80AHUrmML99nLZutRcPWYiRNt7tYKzOE7
r7ptxjXy30o9FLCSnGhE0h7pv1AATDaIKCBGwqg5lI6cLC+VlAdSwEhbVrGdl56J
3xJWGIiINWvKsKB1HynBEEpTwqQgSBePcCg3scEOzvBU8XALJe9nishueEb3JvCw
cBDcl3Q7zDFhGtT4aviKYBCFSyfArxs+mGQw5S/FgByQFKPMf7eSuSdl+S7noHgs
SYsbO37Mse/lXadGJkWhfL9ZhUZH+fA/dSDbA8K2zlrXRzLJ5XCeK+HcfBm39Fms
HZk7E9sT3uw3MxMals5rQtWkxEvqokJGXzm2rK+QZo9XX+KiddAQYiNX/IH/bOWj
2YUIadXEfJrxJGDbMW4b6SWUzISbxhv33k1CC8cU3Gbhh71PBw2hH56Y4sh0+GOM
4XH0T0VfRgmScywjiUgTygDjLlSVWTjniThQ0yAeMo0YZ4+hmEF1YN5J+QJkoGdI
1qGTRtf2cIXEVjyG30oYLMm6/T03RSC8fVD3WmgjviakDjaD6rkYsKalOdqCZuj4
vRtJalNHeIAVb7DwdUUS59WQSmj9WGD5uH8c1yizZcOfvWnWmZW6btksq2X2u/xM
0Evqw0zxeojkR1hwFvKzbMBgM88Hx1SRyiMjxuGCV1hG/I9L0BoXj780Bx15vZ01
3mnw1LPoHLc4tuneJ8f9qbToeGIZFdmhPBgoLz/PTf6h47IhhMBiN9wgayCLrOJS
iZzVdhqeCkTkkjm9qB6VdEeJV4vzNqMTnMBHSheB1daJCssQdqL/n0pMncN0XnMV
2/SCLDKP00jwnP8s4+kJKeennsjdPksKqllBRId32fYoAaZXY45EjfwlfxrJvgpH
6LQqlhulY57c+oMkkbTvyaTVISGUA+7MifY4lsc6YrWKtHdKPsUR72vAe6mz/Tcv
pDk9Xoh+CqpCmYOVGrV1KEJvakYU/0jqp3Oovziiyv6U4IVWo4lqDN6nFI2n/zV/
1eSiLrx2ilg87qYzMZ/RMebxhpGvMUhgBGvMBKV1sja5K0OKI89QEfLcaUJaWYsv
INTZxzNAteU4hbLT7/yam47JV0JrZdqcW75CFQAE3PuT5wcTMZTZj4kmEKoT6MCb
wdxe5w+fbcDtbYMPQUNSfSsbdfCQFoEaikEOOrsdrWdx8xszbWDpDgHDdAW2N/LD
3R1OFL5/7arPjcGbasnFtVyTcvhbgNS2Y1velNtzhuCp/JXhRFMjCMtpNgKl/QMl
a1Sm2hpR4xsCb0ePQv1xpv8AnE6DG2KFwLgpag/1zdjMl1PyjOKeVSVOXMujv6sR
HPMoYJn48eTZcI51fOK0QMdGcsPdqQjMK9t8lVi/PJSzjEX8d/XvmpTPs8eoa8lY
4ORRob59ixItfv3a8QqQ0iS6Ny/lj/1T32S6UUwNM4C4TRU/DHmuya+ikPjNzHcQ
Au5J3F6d7mzCofbAGUKLjXKSlf8LhY0KG8LBruIx3IjspYFS+NfFeuc6JvJvhzrf
PZcFYa+rBIxd3ugcW90Tk8nvAeJSdezfgmsdAvtBTiqW6eR0N4z8HCLZ61IYxYwv
6Rccskdi26sH6KSEUx3TOOZlqZ5/hyfa6Xzi/DFIrCWjAoEg3pgJERNyHdOML85n
uZj1h0fr0rj82EDDUSerKyx+Uy+jtqAA6/Yh79A5koUNbbDFfDgeyrcLEpY+Edm4
VXGxLuBHtQINXlIhkxByKyQoGeVudrdrABkc121+wNFePdjhvy43YOjVLUH1i8t4
aT2bA1cBdwHpKEmcgqRxIgyZoFa5Lxsu0mYGd2QHT/a+MWl82tIE1dBN2q84NMiu
4wx5JTXyYWKJ9g2gtgXZebPJNcZ/dtcQjlprd0BWvwFJMYB+NAoMuuPrr733BJG/
43TDXfea4Vf4IDXNsvB9l6WVjS8NGj+/uqZVik7rvOuMmQWpAf6Tmp9/1+zw8JdK
h6OzCl+VAIx9353+6GlghWwVR/Qn4O8zwD9qzzsZ86OxMR3uEAMmipxFlizYKqy1
wUe/hRjLBf0FlS7GOiZV3kI4XtWDoIJ/DtqAyt1TdWt9eM9aVHFq2LCgNLbOey2E
QBHpchjsNjT4pxnUXrb4GTUFjzZl5Azi4jMEFNcfOcfRLPJs4jPlzJVlKzOCVBU9
qhrNOPqAQF42aPt2I21tPojpU8BzSDIxnL5wXZqO2Io4dnOA0tSohCTUq+67JBqI
1NWSekMipl4hLnIzlzVr3ZyqmgwUtOc88y7m5mADjDxxU9D/4DI0JzI6V8+Bz/1c
m6lbPlMI2OPB8SgK4bncCmm11iZY69y8WhuJCo9fYe1Ny7JKwTtcZiL2EGw6Wf1F
2Rngkds9YHvJQa/TvhFWIZK5Rald+UB+BjGTMrnReoCZH6+k7jNNnQt3IlWHmxYh
fWE+kTECoLSfQKI1ReyX2/e9+A0+GPcgPGZozzy6iRKPm/5c+SwyXtjwUhh0IChC
PGAWaRoXizRfAQtbtOaujYTYKLl0EPVhC2kWAVGyddXCMvGq/7T07pKf0+SFeMOm
DdBW8J1xmO97aTeAnXfCEUm0qzGgEHo/DY1mUoAqrM4XMMdHKH4EXa0qj4uIJE0+
+mgdNHXIlgIrYAu4HFpxNvd/MCSms+oFOQbsZPXPg1efIr07WDflxrt52kJLx9e6
qSQQdqF2kOr9zh3FBi/TE9DS7XPRDqcQ8Pj/8ZQheuKUrNUDx51wTp179+EOOEra
j3T3f2PCIj6sTw8+RYfsODoiiqfOKzHMRRQhRUk55EYXliKjBMW8rkxJEDzgftA+
dV50ugLSVCB6c045GvP/WYhZdS5zXDLDJWzi6CBM4GG1zQvxTTlI9CZ5RQyUMro/
OluOWFPDnB0UYs+hfbdbmeQuSnDl0Ts/ISzdpUxIE596ImwuH9SncskFxS9VI/3o
TJDP8OeS8j2gVcVv7QpbudVyeEN8g0dG3o0kZb9HvZ582xWeLB+XI0z+lnr9SRgn
SnseKw6vQ2GtuGbeqGCgqh8pG4MyTY6wyuOyhLBFDpqKjmSdLX2DsvOWpf9T/dIe
H2mct0t0pongww7dgewP2Cgm8HkXIezIx8sctj+w6SZujztOL6Gr2/JK/sfYF7QY
Ct/4KYjhjjuHrLElbFIljcvihfYgu1aLZWf+hTfkD14wVLrF+wO0QH/ND3HZFgnz
havgyt1SVqOuMOSBYjLPvY4BwC9uQcU7g/RT+dlKN74NkAUsk9EQr6apSZpSReeg
umkrs/SLdPORKRZDHFvLlEuKgBao8W0+oU0XsfSHNEcfCGv2FOCTVRHt3elcRcSw
Xt6QfVmC8H9Ywr9uTikWf7Wlb8O6N+0jcBCn4wVATHAaVWHvxbKQ363WHYfyaYDl
wHPy9aO/C1bbVjjuHppkzdZ2MX/EKeaJ+R4bAqJLwNW2qgjAty98cAQ9yHUvmVMP
YuhCDwxxMgwNJkO14l8gMAIqcwrWa1AShet8gYMcIn1T1A2hV4jBFYSv6ZPd8M5o
WlRCBX0lKfnSzg0TMBR8JIY2D5my4BhbMyalHIsOpWAP1uAwVTulW50KLjYmIcs8
SdBVTjxAXsmvTmZ+SZPkSICI/lqvY+2vup0j0lP7J4jvFTJCy3leJJG4FhBvGXpV
djOiTV0FszfhmWcjsQQGZNS6kzC6ooRhFTKGgCu2+PxDJr4GppBlXj1TgZ/v4EIN
DNZHemXshEjEjD+JmNZfAsv66uiQZaq7qhsF4oStgn3szMupYCXmu8mZ8EeqpiWp
G4fNbMuc3suYbrAn3jtsnsvAhWpcgxOsKaJJCkHk9cmfD7wvS1u0FhcF/351BKHY
TqD3/VZ5ML4GmitxS0CRKLXNuVZUTrpDkgCXtGuH67fSsfdfUf+S1SLdkPSMpEuf
wC9qNL12nakiyjsmi2aBx3CoFKoVQ/Kluu60EixVXmEP2/faLPQIj/6Gvjb+H0vS
VIh+5Sw6xF9Tpl0ccA+QyTR/jObthL8BmTAs2CTNLnqFUIpkuDShyZqoL0ioVG2E
pKJGREQnHJFV7gytEZliswdOAIyCz8XhrfIksEa7lAaiQeh4qOdxEiHXRcmOyuNs
3Zvxi6xjlMnAM+AR99Uk41apQLrCgK+MefXFY7WBFpGmkl9Ud+RyaW2cn84JpbJu
ZjilcI5gFbNi2/Ios3nWtryh/udXiNgpkDOSLJy2a4eU/soJ0D6HEGMCrbla2btU
drq1Bil308z+NbPpcI/oS8HCaAlJb10XvNeWkg9YittXArpQeJbELPSEmvGS0WJ1
bZTl+L7nfKK9fjZOXoDEQL55A1B2BG0LRytVU29hl1divKIBeqe6fQOz+g5Bmy8D
WORvMcA+AZsc7z9f0Sw+qyJuHrKsLzmxHgmTlfKuAtajUtbPyYsm1n0v1XPebUpr
xXxI5IbhAy/50XLQ+Mqgb83dtq+0/wM33cix7NTmnbvlJQ52vAETjB0UXytuP41u
0YeK0ngzqdQUP/mo6GBkHMZ3vZDuRzAvXt+1qOZn6iI=
`pragma protect end_protected
`pragma protect begin_protected        
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Y+nQuPqgYNbXeAO4RO+6gcAnovDyRBdwL/eb080jdHN0bbisiBxZO6XLy/5zO7pD
yVZnb2rAjuBPtvLmfIBODnL/ilbnTq4Xxub5OEXQZyS4QlHBt0V0PWy4nBZ5Elyq
57Ao3WE3uq6gEBlpBLe6N/se8pBX4UCB5C7pvJo4xVg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 67633     )
ngBqSO3shTED5ng6DX1Aeri8HpAsUJArX7oHAjWPp+U4Fra6V3GXa1cViq5wBqDF
XqldQrU6GwwTCGddo5yS0EKUl693kvI31ZV7Lf8S3haOwB+v48/4AEANuBLkyu0F
0ZYVJwqw7uGShXqi7GVkcRxMgwQx8bpaDEsYmyHTNL/uJHrzBfECnzwyUL3UfJQ/
B1XXbXjxFMEDJnTmfUUJSDq6MQNek4zDGgwPa4THy0EfBBLu+UKIAL/2S21aHnUB
`pragma protect end_protected        
             //vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
PNWQhM4YNtgqYDpqQ2QoJAKQL0vzo7XOgNM8Y2jNKungBx0W4dW2my4MxOt53IyI
RDozGfDSteH1R/rT/XwK5uJBOTIWQPQzTs/7rO8LioeHB+TKlzLP3u5+ZtpZoPzi
njKaU7VjbWD7La+8OdVkhQv3gPThYgzNwIWuZjP7j34=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 380103    )
nDRK7DqUbiovnWtnwidmL0BXisJA/bHafnGnUqazCsLxTHyfDEAZtNRJGk64ZbMV
6cI90qZaHd24P1c+1Jz+GPmLeta5wtcLT62QVNDiSvvUOOLc1bExVO26s73Rtxbd
WJXodsrrmDaf5fmGy6bn+80lmi/IW4U1Pc9P4lFqeCbWIEkbEUnC9ThDgVKhvmX0
1Wpe2wqmLiBakxGwqMejyTxePpsfIT0S5FnVa878J2NETySCTTR+VaWu7Aa3Ebxz
W14wga1dpl9i/usMMYCwDB8e68A32A23ikvKNkQK8USDqTe8KVpBEis4t4LcxysO
2h61RrNFe9krBsLmMK1innCqZQ9hRCfUGG7JwS2iujBpoIf/YlwnHpe5XW3W+0BU
NsDBPW743j8jMJtpuf7RBySViPq0svM6IqyaV6RgOaaxDwal6zT0rpSa6o4RJkXm
9iLRPxBQ7ds3XKIwb3kUHzqQjG98f2uu55swkc+rGs+Hak9eBEYRdRvkkuttIHKG
LVpfXfbwbrY3cx7siRymjGnc1rL6vsxF7uMl/ahZC/F1XDsMGpowaK9gMrlNxj3l
FdJUpuG/0vu/wp3zvmOrD7twftpE+3uibac9DMgplHDhJroIfv5N4SyCAQSmrgJA
6ckJNgd6ca/ZjjTSKcnBv0eiLS5bE7scr8LA9jvN+qDfRncIM4oLgJMtx3UJc8cd
D+e4tRIn6HjNs0fAq/yY3iK3tXg99MQjjON9a8yRTMlwYqDV3V04qXPLJ2rzf6m1
IOJSkua1O26MA2G3Lce15pgzMZ9WnnVb3A0KbqDTNEwDVjvQJoJF0YIssEeXlK28
+E1D8v90E2udnUvmrx9t5bMuPCcuDlZx0o6Blg1TZN9B7KGKnNLanunTmU9rxZSU
UGscaHJLS7pa3HSWESRzxBgiDGwDcR8WEP4ObJ9f9PBe264oohTrosKsMnPwK8++
ZV9q87sjQWu+FB91OHMDE5lvFZ0wIHRQ2s91IRiIBjW5apola5OV8w7dj8yN0rRR
LLnc67hXh9qEzZb2Cy3bYhaxWhdTJl9QSPCvQx1Gjk20ZBK6OSpNvf1Q4ibw5X/p
DPs7UY7EL6flWelFBjUs2dWjvmkRCaZn9PV1RfBBqrXRdIgjM03Vucl1RAAeXHGP
mQmu4vqw30Mciz6PFRfYI++Hxa5z5fQFi0AGr2tb2v/fRDxeMebLeFbOUAuL2+pD
uloCbg1CveLzMqEPSaJO95JP2tt1UHCABQIHov7F7Wuamtj0XPpakcjhZWyExV7K
FdiHZqU7fy+F3Cphiv8k4krCRq0SzJGJ49wgcDVZRIIMaOdbjjbyrwcGmxZ/HSuY
VOnsiUUZN/Y8KeMy1zRT9ITJFj7aS+UhEIe7/z9lMvx0SIgohlWEySml8hk2gY1a
3R0t6SdtxKFPsvuuOs9E9utHad4mYYXa8iDmzXyzkSMeTCALohEwPoYg/SdjiaDv
Adx6OUmhOxHqwH2/JCtIoFvUK3k44coUzm8xtjh4UNJ7oW3BrfxNeenV3kK9nkHm
57Ld8erQGc5vDM52a2cZyptgaosXXv+iLedsgZhgxSPoAT43FZmb6+yP/DNg1z6+
+CYM+9ndIhhHyILjFO6JLWZ9RjVDOMgNG/RxaZ4CSRohjdcur43pAaYD53q8k6Ff
hJLp/IWqIs5Tvh9EntT6uoVk6VoCklQsOMfR1B2wLbS4gvHc3h54UY2jS+Y18TIL
75yIDOOXiMXfAEJ5vCqZMd9niCIoEAwqvLATJXfTUlCy/PmCMNNz4sdOKSZKg2zj
E+b/xPEZkhUE8hwRoCcHbC8qTefQdu2S/bqHZQWP7eHjsUpNFVQU44eaDfUpj6OS
bjLC0GQpXXroSQape9PVigfQIFONLuh65o4Q0Ah1a8WYNOBMiHZ6L2zQMfBNu3KA
dqTIpXRSfwBLatBygW7Klvz5f5fapbCkSISswKN4MyQJ83EHRiU6ejAP4hKl2wVF
uz6bLs9Ai3X91z/6tF9jrCPZFoRAJtz02XD+V4AVKxpy3xDSWBiDeOzWnt2Mm8qX
NUKUCZRnzSggMtjR0VeEd2agjOjiPCcmB6My9qE6bq5on0rpCRHBTfT3JUnhNpYQ
s8VMpChYaABMBgMIYBn+Ci4yVVUVRBpPOVrd5D79kQ8s63w+kcK1m4vR1gAD6Xol
kWItMbSIAE28vJX8Zd7TYTyFebHKYbt20vQk8gMyrG/zyp7hB51N+ZP2sfW/D08i
0O4uqiG6iSlaiD4drX8m2UmNYlUfQWr0vlKmTrVlvG7eB5kcUb/tXYRWTaSbvUu9
7qav2D8wao8FmxDcbgCbcnfZFeUHXcdHtEJ19kcCzjF5IdbaB11z0AxPzEvif8YZ
aPIKtDzeHQ/mU4S9wHvATdf2rx+3fxcxbK2iEY4pE3Uya5Nl+ICXgZAGJo7MMlaI
8hfgeKonKlWhlyBCdKtY7c9tVyqhu6K01oGz1fEm29sZeDyjYS+p/mBoNu1Qq4hM
3CBUZ369b4tN9oKOikI2XaQZ521IeDMJ1xfKiO6PJzwcLxm7PqtTDAfwU2K+ER5f
HZLYGSnAQ6/XldqgUkB6mxcx7TeRxcZjqhitKi2H0jAxhRvaStptYn6nSq303oP2
m8iqNqbZiOkPEHVgpqHeo7YnJEWvldNH/4C1OUiAirMhsuLAXZAvi8kXfhjc4bGz
HZzXf8+qh1udIJyuy5V7h4OHegKrk8lZTZNtBYoKMHJOZCre+hcJNktAPLH9nErg
ACoWq2bpaoaCyl7Grb5RAK1FKUk5FJTin5buXbvabRDcG5XwWWB8JgRhCK1SNrGV
TP+Wcnf8djYMz3hfq/ZtRDSY6MrhBEKQ5pST7QJpydECGfnmjRox5LsoLs2JgfTM
wpEKy+avI39nslS33mpKG9ra46YQiNn9142nQaTTk5nvlxISFlC/bzbXfq8uzUxc
mJjF3hlL7t1RJOSK5fdFNiGZ7C5AQ2lRyeanH4phWexftSjqQ46V5NSZiX2zWOn0
7DOKaaFj1szsGXcYjKUQUmo3R3K7wAtiV3Rzrr4cO4t6LaQNlbFMu4ovc2rBcj8O
Wgfq1unJvwIStuXDQIBo6cVd4cS8/+rq24xzbz8lOvnvJ6BfcIOwoZxJcWM5UTuv
MJ/yyTecoF0kzSG36US8TuWmzWBQvU1dspkDBvyMy/b7oBYsdmk9ROnp972TYx/O
KUGKYvzV866pIqwqXymWihQftvuh9Aslvx+7IttGOv4RIyzjrgVOepWSH7CjGpvu
DYkrotazrZQ9rQsJcU+XsiyoevWbxSPQ8DihYeALfGh/3C3mbBVNNTrva0Dew5Wz
Zlk04E4K6KT86Bisxm49hVOEnDgLg0NjSryYOOl+8nHt1g14N/exe3xdFHXBt8rt
TypmKRWS6KRIOvL0mMwILKGUuXE4TqdIWiLmY5kNS+JPPwIVHzaUgrzGzxcESkHg
WNzpxgCC0RN6XphRzR0qZrA1Raepca7m9Z8lU2DbzHKRtXzZEiRIvxfcY7ZomxHn
2+npBiG8r5FjThv3O6sBdHTgK7RHuP9bZBgU19MCFBDHx8E9Hpw4TozZrAAReVZ1
nKHQbbonl0aUH+U98e4gg1ll56vPJQEI9q59l+XkBgHGiXteSQL6J9J15yGF2OQU
CRn1uAad9PWJet5sD/TGzCKn6cMHxOAnKOrkbodNHnaZfaa92BJrkHJr2e85yyG6
t0RzJjw4NMOQtkmtYTpgTIIE59cw3e6mjEwQMHuah0OO0c34Y4gB6Itqujo+gtAf
YFtpCBxIgqxVKoSbKxmDp+9KDjmmtcvsBHRbmfzhlkHrxwW9fnAV+2Yr3FbEVfMg
aPTdTjWeZ/GXLDYLNl/vm+5od5gVNVSLhKuXy5ge38tQSf7PYDrROwYAyo5pfgjm
ZY5pgm3L95NtKmJg2PzgsghV8c9KmiCGP8lM4uXh+VdsukoKXKVWN6wCRtuP9hte
lE9J9RIZ6H8kGq5bULHgBtRLJZnY5P2FAXgnPk2LEYSBI7hpUtETkqnmKwc1f420
O5opOpKuA46CMasfoXuoHOU0IpkPNYHPVPavFlvVs3sKyJm/Qmx+jg5f5gJa8TMk
zxrauLmkxryYk62peAlhBZFOD1lF4cCTaZ0ks3v+CvzpNGRvpr61ndFzgwsSf7e/
ODiyzv9x5bXhlgZ4sgQKl9Xk4jhFL1soW84FD3kvixt+jZLKDmPLnK1bHxxIUtzS
nULjR3qAROvyw+i4JM8wDeLFvaZZZ5br4fG8kuTwiIwtpLiqOeT1Fv2zJ89q3p8v
2bZWsAPG4G/8FpbyRWkz1Q+fQjm2zE1fFPSFkSDfEfaR4NuyjXViHPaXnhDj82uN
gpagt50rxI/NYhffdhA7WKpf0M+KMZpG7W4r3ynDvCGEi9N9ZLcggBysjhrFCIuW
Crhtl28LDQfTkSeGzGN17zXKa5bLRZoUb2ts+91gAwumqmTycxtfpBIbyAOe3xVE
blWZtWvYExjWXfp//uRiOrC8uzRXnH+lBX3cfojr2KamhIjDwDYMwW8c0Pd3AFX6
BQERVZOJV1gt+N8Yv1Hgh6KKOTfqI51qWEy6UAdH8hl2i/L/I7GZSTf/ynQ3JCZb
XTIfUrGtlFa4CS0qjqNrkb0rtwA2X6sDPcn5BwGyKLNziljDChyeCNNW4UNTq/W6
tkZJsgiMN3xCBfqkPMJ2hgdbTmq+tvTfvr+Ah3f0/m6CIsnvQn9wB0/AyDTyqbNQ
ZaAeWBXalMszPUYST3jC5aTlKOd5mgorouCP8B3sCnyYxM2ac1EmcOJ+qf/pyY5A
6LejKATscjr+K3+pj7gHw5H1cNLYoS6G7YKqu54oR3hdt/RLiavVhbxu9R9YK7JP
sIycDOtjCm4oG3VlO0r8Z92UvdLYEavI3vp6s+JHSbfAqP2BhW6e4A5nBDu2CrpL
Cwoy3B85wISxlo0vP6SUdXb5zUMcrQTH8357tfZ9njzA5gpuUguC4D57+qu+3U5l
39e4bGFVN5D1RcVbodxlwnLlTDED8U+kIiULcWPtDP0av828AwSPZjm1h8AHPym4
qTn8JLvI1SOINIPE/k+svQ9F4s67fpB1VE1i/nvJzcpomnaIYLCIb3djthp4WtiJ
AmSO6x9MsnwtcYC3Ojab56wJ8awfC41WFOPvqqOX2LZ/voi2HaanXMS48uGRHKxy
/qFF6jmz5DlhL/8rNfUePKTySWzofknq5hb5eWJvKkVlS1EpY3ECAaUPpy5fzvh3
wdkol3V17VtT3TOt0QNF7U4J2OtXjqsnDnIV41lx4v8gvJwrUUEXDMUGcT7WbHIB
Z5pjpTtWqx7xJ6mgwQpLiTqIA42BygyI9BMFW13yslc9vYT3Gm5R9Js9uEHyQtWw
dJjGMYm69KdyilIHADMPXCFnOyXJrI9jNln6pDezmSGVQr0wYKjnR2sYSV9go6vq
snUqLnC3xumd1dCLbf0tX+SOv0H2RednDgpwi/Inl4NRgSQsi2ppvweb11s9YtKl
PaLpwS05Wbgymsi1tmM4sz6SMxn5lRSB2zW6vlivcCUP5Yg+fW0O716Kj/1TPPFK
K5mt+HtXIVDNc19BlJ0ZZnN7Q4OrXj5V1jvTUBXwzwTpBK0QslSyYUhqUy+b0TZ2
lBVWbykI1+v7L6t/MXsq2fmeBuiEQVq1cczKUP/Eqk2z29cAoPZ5A+I+m7XA+GuE
PtyYg0BUKT4LUwcMWC1D82cstXvkWShxzNF/ZaAhdrdjjxKD+Jkm+in4UtPvwu2i
YrmSX7fA+SNdjiGJKVGWISMNXBcualKzQDoY1A9dqbfFL1KyKE+2LbHZRp0qiSbn
zXTRXI1GjGZZtvjPrRQg5QFjFa1bzf1Zjaw9vRKnRxBRLimvM4jz2TwBbKAaQdOc
gHBu6v07tAaT169l92T/TFOn6l8+aYgzOdNOkCW3nFHMBaZAbBG+6DGEgUUyGzl9
ytJJd0pM+YCPCakOh4JcUZq6437mIni7K4Z5+4k2OB+R7SiEs+tEzUIdhjPY9vC2
jqrlUYp4qOHMQd/a2PTPZB+tsA8jGXooWFMMdUvcY3g9k1mz2bZfvW0xtep6eaTB
29hC2lDY+T9p3sC0gucvtijRKzv3ZsIz9LowncRxK9zxchKXVregrw9kW5YbxTgE
WCYuizYMf42OrGX+mw2PkE0/getPF3IJ20EKZH9Hmjf8PvH2l4hGGsC2Ym7PV9vc
zc42zdMEbhYh/Rp54lmia3ZRCdN4HBCeABzKPLsfyVf3lVfkJ3IGRXQcbC38EH/F
Egikzt0Z3Ch15FCJDY8uXSTpKAzInnJYP9WxCxdypi9Q6Eiq+rnHbJ97ev+lSwnA
YgU7l4PbUzSMlNfJNGKLSwnIZyVoZkwqAt0ThzikG1fw8+CowuuEiM4ED6upS1Wz
6LVCsa/23Ojlxanu1UTaQap8NgKspmlbDweXLbkzzKVeN0tayfh4sqxCbUZHBPk+
nYzNPazV6BQnb8ApKRX9WcTURzqdfzcOdlz7LDbkONzxy/U2Nvkn90tfu4BneA0o
z1xHFcWDpGGU3nBTz9jGf5dwCpl8otMeYKEknfcWA227OYsu4fV8eHSYo2SZc5fW
i38PpzYbJ3WmfExZhWPhMZGO6OthwFCxoNvX+Px9Zc+StPmT3SmN0maBDE8OZqhF
mVwrUMAfzK2q6MNjxuTaHYMLZMOTKIVCpaBcCaEzdJ7cB90QBHfYSsFHJ3NT4fUP
En9FwRidY3BeCZcpfSG7CV6kWnsF3NcxZukMK1aPSYvMXkaTvL9QhgZIrGy6jd8A
pvmn+I8+iCjuci9BnMitDuqhtewL7qaW2x4j5XxwiCuwZMypL/vJkgBbSwuXxpkn
DLLJUfIGLb5sFV4TumEgtkFapkCJfvYHVRnrG7QHqNQBj71E1/qysmE2nr30vxUN
JQNIh0cavRl5PT5SbRPFtUXvG85BNHrPdvoQIMWHCWq3e9nhsPaXF/DVJn6/sRTE
kRRILjBNuRCg7BkICDYqv/Q2CDkPDnSyqSGuYToSAy8hENzwY8rHp7vqQTRj9E0k
e5c3xySsJstnmPIHW1uTHQCYLR6PXsvRgNHuCGh5nF9dSbzaWEN8iTCYsVKGKwCN
c5HJ0ZEd29h2K4ZAP5xatTYzwp2Jl6qyc09qR2QBeCnyLZoHDwPWrl1sBPX1tQSA
vRIOccaPMUJ7Ns7czftcEsK3yEFve21ymLzZCwL3nAJafBUPxI5pTY59ZazpGdNq
ldVtv89Et9d6w05/J5JJAFiqR39nk2gvaQKzQHQDZSSlmTLLFRItwmlBp+2U8zlb
m1DsjLTZSCTgXIZMPZYQuGnrBrAQtpL4YFNKEQVunYD/QND1hIQvlGcSjFKS1kG1
YLNbq8OzgllGcAtF6e7eZKEN3YSWxi3WoS37t0WSl+1V0cQOmJdwPcM8KmfAuGFI
e9z6EuiYN09ap/MP2UduKx2AVMDE/wfQfA+R3Yd6smJm3jjZciF6NXorYOHTTda+
DhKLJXZZd2nFfXaosvG3OpHxOfu0yXgXkHo6FfYT34W87ZnajzBpbbguxw4hoT6M
OTVMhjDShNqLB6L+UAfMKCO2G+57yQdcOY0zGlj9USRlglzz4RqSEkzVP5EX4OVw
RkgYp9WuY4sYvaJLczjweIR8UzWWJSM4XzzZ6uCjyXU6TlLrAFpSskfj8SW6s8d6
pVjfRPmJeiIFPHPJbXGyHES1zubUXSBP6a7QegAjFxikEC8PGRp7uny/GPlVubPP
xOicFqO/k3LEU/mF0SBmnW3Z3EAq5UoeAo15VZ09JCZ45qeO0qZE89ykDy1WTlFY
+aAYDmkZH96/hKdiqlEOPZ8+bt+RtUyh8s/xspLDA7TeUYc2unQw7m9z0+XmWM+V
++MpiJxU5BsAQifuiwGaM+zn+wH9krfmwkCGkY5q/H/fFSfNaWe/oRPatwIfEXYy
habYIhG6y0YTlBvhInLe1zxWQ8qajmWJW1OYzNGCp9kWSDrh45ibkgJULCDdesbp
hry7Ca7F9Z/p7YlVep9ILTr0et+OGCrF18p+Y8OZciKe+DwF9aqdjmPqIjIkhjSG
S8X5l/iU41oLkKRGwMkngxZaULpPbsCRmyvLoRp09zCSJiUaPAxkSLv8pFGXWDrZ
1tpq8wXxM5I9sHaFJYkZ/p5TXeCTxYx/7ECo0gVTYngxe5AHpAoKabKol40pB8Jy
2LrCnrV65nh65FkjXrGaOOqj0cuZlKOr+2D01FgqZf+3oiAuhq/a0rTqqfFvAybW
1h+tudQ7ZndKclhAmXey5nyatXav62ZgT4K4SgoB7Gg2NfW77H3FK5m211LSkbzK
GpaDlIL+LhNih/kWj3kg1U0ItfDpU+aRBmakp2edzxb70SF2bl8Q8orH7bAK2CGi
l9XtrhjIZ0LSW7+G1+NHcxtdSCAXl3YAfjdoSDBRhi4uXGQOPzZYi259vWZmxQP1
uE2J1WLuTFrEYLjz1MSmVk+tB5/IPz2wV+zIN0ZMOWF/ONlVKMZWAA3vgw9zKTBs
sGc1dyn3KW0cnfK037RAGvve1nFAcYkQ2Y/N9AQJQC2WSNBKCAsmf6nbOO8er1l1
iNnk2a9dj/GGxAViOu56XZzP9pDKxyiQxPxBEsJbYhT5AfdU5zYe0EKb0aAQA89o
A7H5TdNqWuH/wJAXynCsClqZ/B3W0+h5qQDS5OHQzYmTu9VGnv4fVDTjWlCUc5oy
aj3VvBvRM+38+uBaqbb6ubjamFhv2O/0NYUqFYDg0wTd8gvnK00IZS0a48GYgcwX
tMlb1bu/oDsguEDqAuSfMKGlWETUCblgmkW2bAasJqcsmzRICKhWD//BDA54MNi0
xA2TfXR+ovJvn37IbiybBZOnpZ6S7Lecbz+asdX65pUhkkX56SPDyWe2vBJMNURE
USW57VNoAXCamyhKgdUd2nhJh0WrJVBrPj/SMy+0IPkC5gUs0qc6kZtdjD/xxBgD
1t9ZRIkJCAJRpgSQX9qy9B44cuXaMdp+LlBsREZ4DGjyV2COpsPtGdYHN9LhPUqc
uJM8QKecV+tGpjiYUNlQ4fq5vCxTY6Ij/nKCcf+T/j7WP72+Y5sEUQfhbExFBSY7
gn2ECvuqhmUun/vGwmTZiOCTrjRP9+ifs9mYvAgmRuVz4zUObcFuRniHFYPxiwa7
RnFt9clp9nkOfL/RRKME7j0UKtICDeDYfiG6qjMjgHbi4Q88eC41ftSHEBvXvwYF
p6xVrMjcRJeW6q0inJ2P/sbfA8FRf4YNKMMu+XYpvA81sO38truEAtJ5H0Je4emK
QSFHXd/iAk2Cu5BITZJIPNMbNKJ97QAsJY5COgo+NZ652TaxsVfZ90u3ZD8gfV4h
B7rUtiPKw3B8TfZW6L03ssGBxricerAr3QeNs8xyIthUsDKu8xdsXOBiVUSRDPtt
rMeDWlLZPuqg+pZ5+63H1LaVP9D2e6kK3MTE/TwYAk7seRe3MP05i7peAyOG0IT2
dj6+EqV4TXDJx6MBuGbeq7VQgS1iYHu9jSyR4/Ue8qmNkowI6Y9UMbklXalR7qo9
seG7L176fMQVRiwtCHT/YQMtg1h0BzS/ywbMHt+FZP7d+Z0YMEOjv37NNDa9EAj6
A5fZR7TcpqjtyCzLjMp/LCqUA6WpP7pA1xTW0S+rauHLQvMsMWwXOs+LBX68hgMD
XXto9Gz1YjHZT2tCQ9DKcVkGkPQJT/41W1j8wHTVdQ+BI0HF+34gfKRWVSv+eH59
0ZbNM8OWNs2BBtudqLCrwu0uBk5CvDRYwJtRKt1X5a1a7DJJ9E+sbV0CKto1XH8S
0rtFa68upabTt42X3iQf+8c3tCNCeiBFc2UkCoS4Xdo2bzbF+Tq8tZ23pjCfUidf
sebgLwGLJRlU/tIGoqWGx3eEKFsT9EIkKUGB/tbep0x7JkhxnrFiVos6DdvwTKKU
2vJekjWLv3bf+9aOU3a7VEnEtBPLzlAPnhftk7/CyTkSl9PT7FO8SeuIdj7wLEjC
ZbeqhEcYGwh69JVQHLakJ0kSRIILAhbxL41u9PN26P/PWR7J5muninSGjFIlSV/r
OrbtDs9GSjpIPDenoLjvhOt3MayomKdk2d8cYPfUoyVq8ySQ3xHuSQzopSAmV45V
1KXp6AS/1eXB9i4TqksckUnZR6vdHXhgdIKDqypr10poCKUzgbt61mgHCnF2f5l/
CHHD9FedWhlA9V7eg3UEfrwwVS6ojeNV2LSMCb1GQsrxpZ+nBUvrPKMhr2MN3129
J4lZpMRrI2htTBPoKl6f2L2WkLO8XLwplx9XqFmw5mMmP3lJTPj3g0RZx5XWROVA
aR2cMJW0OJR+ymplmKjxLsmbkPN0Zh/iDbgxrObpBdkB8vwxhyztSfBHnG473Yy8
qjpEBQArNeeIHllMl5g9Kcipg1UyD8T/eJSrRJV4uSMbgscMqwxZ49ZPJqmkIctJ
akCgdPFjNYN1uLIKq3K0QfopWIg+TvHHidc5ELPBh8//MBbe9WcbypEAbpXjd3a3
xfI8gsUy6xYTBFZk4Mqcdd8BhF3Rn8m1ucj862mZ26UHlBkB7udpkw49FoaasZ3Y
KHnRcyWZbNHS+2vfmG6YJQ0M8kDEHQGL82lexg2QcOlj2VuwuCrqX9wCG3qivrki
dZD4HvFN17xzG+eU64dTos6tzfolFhOOVI130gWNqnvXCJpn/tP2gnv3y0r+B8Zh
8r0lrpVrp7ZTQliSqIGtHrnn/rU7nlq+gXZwB5ac/mIl6FbP2bUXpTNewpDzodoW
T4eqIYzM4G0gizrAH0y9kKn3n5HGVMtRVlLcNYb4hMIjxId/9MxaMb3BpQMINBkP
xqC0+4aPTQOwwOHwnoF2ejJB/B0mLLWTNnu5Qo+/aQltErGUmuoJlCPXbRVYcY2H
eOTUmAoj1e0pFkuGJzRMUhlPquBhlrusAL3Y23e6kOXflHut8SSqtPqp5b5UKgk3
Rxge0hd800n3hmifzV0KDJ6MKF98XUKqMf0RI4C4QlHJ44+1o8PntI4nRNhGzoJH
L+UwEXbGTIDIxrYmwanScVVI+H4REk4mxlnl8nPKOAH9y9SV4+WX/XFzyT+VakyK
WsauqRr1SdB4OUXJtdGSeU9s/lsgZwa2Q+S7lhYflbZ6hGapZNiXpeMv9eYKEAzt
on1VCKre0JogsSP0O4FsjpvUrE3Tv1Bm5L8gWuf/TztOMFcXRM+SApeFSg1EOSoU
QWttF1taNac3jG3NVbX404DYEyDiZEBrDt2FRhyaG5tZTijORyPmEzQ0Kv1OuBeZ
IOpF+h9C5MWh47XTm5N1AVaFNr+Ubp9kSXdeq96UdigoUePTSgPLDxA0JQiVFWP3
0lvflncCuGHIKfD8kA2r2rFm2LI+2aDp+U1kYSYPbwV6EMXuo9jWeYf59FhXusDh
UWF3bzzKTRN/uOUJuld+9wLay7GnYnwRbhjoi/y+queLULhA193Oscdh/ve/gvjN
AWaV3x3SrQDyN7yiXmDTKWyRfTvuNtMrT1Mm5xowdvml5lbzUjxoDExZo8cDcEbX
cPPnxLw9GqFBBNFj/s1HzYKQUi+u3JnAESrMs1Jqb+hH/iD8ffCZQjS4M29e07OR
oCc5rJ/woVXYTgD6Wv31oOkEr1CcqmOeNpUvgiN9MbPnJUuX44KM7Wc22zyFbFje
H8/tUswpRsyAVx+K7lOx9vRkavcvaLuoNE3tMOEdnkXwYmH6uHlfHKzJCAJTcImo
j+zFuSQQ5T5v8wNfvMiZtsXxuBOuuLq/RlJMnh3/1U83gDWVCa+iH48PFYBq/NcH
kZyGfq9H0hzbbtxjEgudJcnbiEl9udEyyxPQt+7GWNM+uWsloAsYkS5uctyW+nPI
o1IdONCZShfx3QsF1rfcJtY7U+9zaUNQomYnBcFDnqBaJW+B190Cj74IycTz18SF
Qu3a+48p2ah/tX+BW7Srz6H888OHtJmgLZIf0aiXAPxXrBYKayxpDGLut1hgpFpd
27Pkb5g3XxpK+XpOmGmSubwOSpTdmkSuR+9vReGUT7Y35e88ECchFAd9+M9yUNQV
xNDy/C6WA1y3hSysj1b3LpvUQIg61O2sgxyXzj22/Q26ey2wceU83ew9jEglSNwL
RLGHgx/OpOZZxLwlrkRneSPLov8aY8thIytDaz9GnBS0Oi8Ca3y2PMRmEU4UCeWE
wJj/IOde5G56E8ABfzjPdUUCYd3GmKH3J+T1bDBNYhIu7yqBRda1JwpL1ZU9nCTF
y272a7hLi3eJN5+cY7/hh97P0BX9trtqMUeJooFf2gNMupGHV1kaGgPV5VkndReA
EeSd6cShPiV6PUPurKZkInppcrow/dX+DeEHDTNmKWYD1c1o2vEiEAwjMCKig9wV
quvZwUuIv2vThzU/gmHIm1CSX951rfZbb91hfZoYJ6Qm/iupzFpgyt5NUwP+focH
BL/sep4Jf1Vy19BngRwj4WV/WwxynxuAeFymsTog9lz1SyAwrPTpEzpq3B7NGq+6
MvuBRVG6fxbstU09/oB8lq6BiBFyOorChthc+ShUSI0K9WFfOoyLklU3WJHooGv2
//sNyIEDLDRTLTZfgM3gFYN5JUaM+t0U4dtJRfzaYDefQsb5erwh41M8pXWO3C+8
0DmoqgdzXLlI+0NT0rpNJRCj8fOGt+h/cZvSpcPZ2FnnS97wtPyqADi1UG1j8eNL
im6rULUJRWVI5fJldgF+6cE21b3xYVnMAytoiLmI3gLABrS8y88hPhSlMiCHkqlP
yZtARfeDVvJaq/wJuAx1HwCMjLfqQ/rE0omzsU6T70bde1BzSqypYXFOF3j2nmKe
iCoGDXn/tdJh9vnwSJGObdC6rRjbA9Jt7eEWpaHnx0lP8d1nE7OueHDx+ZNmHueH
K+WwALue3XF+/uwogXUbqR1PIhtTHQ67V7GMMRgwQMAgmFeaKIookuNTth34I5yS
PHSc5OXfF4NH6FRr+0DHVJz1HOkqUfdGG0g/Yl/U3tEAKAM4HaXjuEJIxXY6zTAx
SC30nu81eM2kAMRIHW9FG7lCRBZM1Wcws7OCbtwT1hIbroB3et6U1GMTeiRzIc72
qhLEWcm5OA+OX1Gwj9/RmM8TGaoc/L0Po6AflC4NYmuEpGSxonmNyJ/1uR+p9C7v
KvU7gWIYLvca8Yy5bGRKXKn08xnOANynPTp8c0qHI4VIJUqx3ZYkMRpTef6beFIf
LVC9pcjO4PzP6VD4rZ08zugV4x4Q9qB+Wctf4UsMW/E1wkZEmpnsistAZs6/bI+Y
ozGZY+7gV9s7w7b0mLfuxAGVldlss75j364rcnWNfvN2oWurYN66nB6h1WbBDm6D
0XkgbJEV7MH8wsBbhGbeXNaA/UBnOX35FvzbCKpU3DAVIW7BVYAS4FnKcPkPD66N
VyCFZgPx9mCwJY2uCnI6o0j3uyKbuhwpHwRdz2hTnmJVDGX84kBUSUyG0oVpnZ5B
cw8ONn3dSZg8nLBHudnnZZbDoXAJEE5XQK/pIspFY07PunVBTaFVCKlMqTAOSQoZ
CvzR7Zc6BbjDSWZcfi0fc1rBc/eUoDmUvqE4LXmjRigT3fYwRLKpuNePvtbMRCTk
RcJPPHaZ9I/YEebdWBNkVNWfUfbsRChugyhbgtxqHxjFvy5X2GRHu0WrkmyJvfHL
SzBlKwUH5QaFouHQhKnPE6jE2tN6RikuqbRzvWZI2SU/EbYqzSFcgvTB+toBS0eS
xZUdsdjRLd2tsLz+13tWMMGowZoCBvzeweUDQ3CtFFDzrsFpNwhm35R4Oq4GWs0z
O9bLVKmUeYfHK4aFZ1Xtd3p2MdX1G2EKTAzoBmCG9JGA9P4Gx7RmrduYGlxOTwE2
m1O1hcm3s7B2XQgiiKWl5Gs6U99KzkA6DXiiwhvWKBV3+ffxyW6xosbGhzjgU39U
fcLkLpYNQXqz0lia5KcGh7f+E6RNnJyFK9rf6lztNiguoQi5NK0bezqP+A09iEYG
M5etiOKe7LA2Xh73MBCZXsRsQ/GgWT0Irrt4z8YRfYQOTQGbf4532yLlTqWEeEtH
zNS0QjfiLIUwoEBqAKTyMbbQrkHxLlej6yKYEqK6PDHuosqpT6B7E039TBOHO++1
X9gcKySSblK6sR4R0khrHrbs0fuefn/IlyJrMK1YK73gsIbVxaAl8zojIC/52Wp5
mfJ+BozwEK+qil5KOO21YcknenLewNLpZyaK2+4C3Ta0UhmpOBtmAGUKQm4iphg6
qqt4Gwe45IkMeuJw+fpDkY/vK9dC0eZxEfzz5lgUL1eZrnFYjvglGOu/7U3shnJ4
vjlFPr6KlZ2dh+yKMzqggoVOCc9ZE3yZFMqte7SySSf7AEYW9G0n03KHmK6oUxkV
Cnixjpx2mKmXgcFkjn8roz9b6Oek8DMgqi/ts/iAV3k4JH8pE4iPrXhzeXTKEGlJ
Al/vj3Mbmk/24esVRi49nw1GuBaSleuN7q4ih/53Ko2rdeMUFS/NgkjE1LLjpLP8
k176x4kZHXmsBDBTL6JZ0Hv+CZZMPer2enhpJIB7w3ex50oSc+cR9/6e7XYqZ/eA
nt0fzXaH1hf8XxtII1IR+6rxu9ivhHoj0jHlJrLyCXS8khgXzX1gzC6YEtU0StfH
sfE8tHLwQq6XiEWAeFr3aTZ9hG7t+7fwR2VMV7ninv8HsIIloMUmntFMMlgYLNJ+
24l/SY1mwtdD7Wkrkp6UEuny+D0BAP8s+KcqIZtChhu8ewE7mzAgZrSWi58+xgtO
LLG9EUvXGeXYwx1+vyhSl7I06i3XAskuBISJxYlKQzOqRm+vi8rB6QtTcJ09qu/r
lFXCgFxevGKSpTfNGyRc7PwnzCZqofDqX4sPzFPBGkQ3zVgih0ybYTxGTAyynDev
jn4+wMl9FLH5XZEuH+CetuhmwUivw1yiWGeSWRzzp4vqCZ4UiEZxn5nESyYKzYaH
+sYNpcAA6c63cc3AYwwisCZ4fR8otDLMyyzIP5AsXMNwPJRkrvYsEP7bZgBICdjO
iSLJWAbmN24qFYqVCyQyX1VWnu3JZ1kNgztapet1bZv985Ak6a0HYUHnBoX99v9e
y94plERqo2PnqQLDCMdl8pk2w8Q0Y1ODCJ5M0oOWpQYdbdLMK7k72AU4ExLvBmsY
MAnVz/ozozW5WIgueLNtlJUoaYMAfNpdH38qVlQoM0zUbtlvNK8iOZL8f/8c43/q
g87/hhZThHa1VX0eWXDKAJuHNHMjdM1+D76fwg/gbAnSo8aw73TxMUv0mZT0MSOJ
fmEYLM71Z+hHIQpgknSqLxbmGrmOo3sokX8Yz/iLL8esF1HqChnGvEfrQpcSAvqU
pJ6sswbmADdAqKcYxMFsOp+r31SLNYW5sQp0OaJR7cnZpBVd3AfFyvh8JJOlxk7W
XimKUrM0YSgt0QXCQwhw25aq6t/Re/TvX42HafmG1aqY4t/oMMezTUmWqGE1DU+t
iu5vP4ZsmI28O1kcmgbDpU7PU/0VUS2ch5w3wVJwjx1QrR+IgKB52AZmYhgL8SqV
gJt330XX0IgpzXPmwZ5NCmJENSPB1UthMVAnD1oxLfJQWL3o5DndU736hPsrfn6F
QAJR7sBLwOd9zMw8gzKArc449/23kGEK3J6xJ5AV0dyjK7BABolAp9eJhehF6S4Q
aRNwNQDr8vhIkL4eJ5NrYPxRaSCU6Dg0qDt3bDU9RYphKtwxuAVJXCn8sU4p1WP8
nUmq7tOCAEEQtTRM05pcL5DTJd3pSpP/qiVOnYvPVU/dRioP84y3IpqMTA+SUV8M
sf/txM7etZwa3jqK2mbF1s8cAAdaye5oBxXG5i1gEpzJHWG9XXoG4/xLF6NM45dJ
idK7M8ecbKgDVFdSURyN66XOpVOmoZU7S4FBD95NyW4cgahpNaLkbFR5BKo0yy1/
LnGenT40LNEo0AhV9r3fu8ahxXUJSMq+XHrH7kOms70XNRTNAa/KhnGl2F13GutH
Y49SdwZjWsA9T73SultqqxVcSIkje1VgqKpjQCLc6z0t1qj1SaW90BxJmQvQhekK
t9vtv/XraE+4rbt8YRZeL7cOKntWca3jmgSYbifkcl5wNudrkKQWoMWXN+T4+4nY
aXnplUlGi35Faa77vW0ruHh17y23Le1nzrwM/uFuqu0XIa+0WZ14hJb/e8SKfYhw
XgL3rtBqc6JVB4R5qfACNxWUueqvQSob0FKc4Ylnf024ACGdX02wJTHUserQ2NG0
DgVtSmyMWCVuZ4lr6Qu6okJzNxXLUjpjv8yuMZtsetnJU/seMlmR3W1Lrdfk/XKw
fwCMpRafQeekG4+4BvlmoANdyKVyOMWep2nkH3APGHSWn+fcIivQAavIPVKBfYQA
D6hYdlsVPYJz0SSjWRbcbUtsnVNNWaHsUoBONvKLVthuzmrqbO46k4/eOIFWpgx4
xAJiiOG7Fz1NtBW81X2+/o4x8EkN3/65w7MCtgqOe8ZjUEBksqRF4Ep6LaIcxPsC
2tfs3sOe05DiC4f2/A1RbgDOv/y332BTvJORGqL4hCfjtpF3dCnurRgkKdMxJ9Gr
ln9QDZndPGu1JTfigjgijU8QPZMcw3A/zg9G4uDoyjPIhg5Q9u4BZIJ/fG5K43tv
y1AWSDp0o5vi0eYdjTv8xpczyaZrzqJXOLY+7FVjIjEka/NMrXnXfbFDs1+MGQxX
fbcDlim/ZeDzg1ipYx89E8YUd6689e909BYqBbKGFhZ3FtWijOeStKG5xMKnSKe8
U0bSJ/i81X4V643ovqOHBTIUECCTDFzbiDQfKwuOnv8NPy9tE4lW/LQZeJvd6xIL
LIgBeXOn3oqafL7h7ffrJ2S2T/3d0BBaJQBJ6g6MP3xXbG7j2NA1c4fLSFxBOvuP
Mdn7miMNa9iHnZX6I+jjHsq4+E/8s6tmXWbquj5uhaG2/JHMn6GlZhFtf0ZIWpRn
pWIu2Pr6xk0DXFRyJ8YxP3Pt8kJCcR+30KqtMocerFwxR9jLkU3RCLBc0YC6ddUq
LX1K0qsQktOH5vE+EHupdrZd+F14P34rZtOKP4Nf9YmhycyCwGB6aUosTqiDVj9s
WszthTW38g09+wTEBgg/gg1KZEZ9qyYybcgTvhikjZEJuGHiP1s2aTCdwYGf/4rU
wfrO1H7Rfa74+/TVkhRK8sKKx44RASi4BG6jMjFCYxI/ClypAkI19eyOvCoJ367y
HO+G0YsxYrTyw9b7caPdRT2JrFB2gsmQMgqf0Wbgu+Asp7h1X7B/5+prRwg1WZ6c
xWZ7Z9GCEeqaHbAarFLtnvn+Y3zEHAVcttckd87PaVsLLixpWXrylFD4ClqoSh9Z
XCSltNErzj9k4n0GgiO/rJqoiEQ2D/qWi78N9TCXGOY2BvQ1cvrR8R6BkvD2W1kX
Q2ukoadBxiAZQcATPqnwD7JQR0bKpusbDRJADbHfdsRknxmMlTRo4rQuDCxqU0aM
QQ+VdC0sPLQqmHO++7OYZh1W1hgUxnzTNnWfj7N2asGa8XQrM7MI32VJ9AWUi2DK
o8vsk6xAhpAQCDfg3xyGcaWat1xdLjpK5E+cCtnK0F/gLlGApDxf+VN60AdeSlbq
Twz1FoFfrLQRAO1IbZfpElDwVMm91Y9X+9JEYJtrqW1BfNHxARYLeDn5f1DZsIFD
MojGj8CGFKf5TEj0ivBPfpoMfQjPqa5Rnd83NtOTsmFdXZvDmG01TGtSxh3f5p4h
yv9xzvsqLsMvW5SSbOHoDa8bv8tNuLUMQ1U64rktpoEfamgMOKy66iO/x9RhLNk8
hvPnT+YrZj/DtRgQNPT1W0oEmq2L5A3tSxBNuO3xbg1zZNlTDujTUctgiiHfGwVz
zAQNjb9YTHdCPWGnxZVWssU2jRj5xgGInmhFcQuMJCkv7PK2fy7NOmD+08aJXBJa
mh0JqdVRwm1LRThebsW9nAiIzxhz+YTtCAmajbWzpQJFax8SLg+dyDQ3T2rI5GAU
iOUbrS12X81NJ2IsEEU0rj0CqkXzxBTe/Cigv3uiuMAyXYbT0WKrOxSAAFpOFRVh
VraFtRCqdq9aCKGqbAi6jyzT5uw/QA1foGdljxa+qgp5rys0s7C7KlxeK9va6doa
ox5DwxGt9n7x+/wfFWwBJ5lkzMthB7LDrZGlphbhvtP1AbFILDD8lKJtMO0/cXmL
NCdrNqQGVBQy12r3o4NFi5d9Y21tVpqk2P52WzLJoNYmAo2HL3hJxxR4SjAQSyqF
u+A3xft+hJ9sGxs+KTSrONbQsq57K7dq8ZjJ8FfyoXUkJCBuCimWa/rEWFM8P+yq
AABUIgRtz9xlTMOT9FFhZX+p87fMRYDDJIDZeXjKEJbcl1B8vAT5xzWhSJ3+/qpI
Se6tZf4ng4aGuZYaHtWUCdIZf6uwiOOe4N1ULnTaSEF+HUJnE2m4Y5yvFNONIcig
PvSNwn/OPQQJKE9p2lUAHZJ2bTpO8lqpa8kSBNmR7aigFVK+PMAWp3JSBrORqskq
CferK4BVuc9DboZHjta4u9gz0rZmQbSDsB8sBmPmxz01oWDiPT8QtGSyM+wLKa1w
fPEmsjR8Lryd/iaXeJ5bgnYAG9invUNBWMintv07QtzowyVpJDimKUiTENwpNxec
dmRa2nkBcBMls1FK6bZLp8fE1N8/Nr/Ek29alcEf3LR1MUbI9m0QzwEm+5Dbba2m
0R8L6zNfA9z86Ueo10VdnFa5lVSfwW6/IYMsYNva90F9z+7kgkP/6qD1vye3ftML
BHnLQyp3RPy0helrtc4an6ar5HbRb4V6xl460nInfGTFz4NToeGMzdNtDJhPur3O
Se+UboYIylbSUKcuYeRFBwpmgbAMqraX6+bT/tqi12hLByDyV8vYcBbwjSU7K/n8
nMxXUjfluDQ/vaLWYwqdnSBzdhhk15g7J5CPVrgfyIrduB5I1bKOgGbxEucVSvJO
Vr1ZWlc2CCdllUVIoo+9x0W72BnoLuX63q7SlvnJPahjjSUTiadiziOwaZGRQOl8
VkeJFxOwfmYt+h+2sHmlw1bjwTurQ3FqkbX7q4zLCK/CHi2yhBY23RZbnQfVjDdS
usByQNTzAdjB2kvngFcYlSdHS7apGs+cSDqJvw1vxjnM8doCS0vkifKJdPgj8e4A
o1uLqiLSZUuov3kcpyZc1TA68wQRyV9+anTr+P/aWcHr4u4okJzYvQc9+oWg/eeh
ey/urqEtQaLScJ4pWSwGuS7ZiRou6CQkJMnal6CZcaoSoEUAzHBamuq2JgISBWGL
fzsyhIGVv9RI4kp1oR/c3zXClHX3N3P8c/W7nLXFJxJsYnP3mmCmyv2aTc6P5DF1
VOAA7t7cg2i2JR0vecrjCptGfAVVTBWxPD5CivDbQqkDEAuQrgGB9/aCs4u8EA1V
qVVrYymglkZ/YcQs2eoJAp+fD8uarUlFwLZKSryueeDLEhy8DoTPJfBnlNlEYm3O
blW1Ck/RaiX2yYmXHfHMLxrRXsdaw3pmJTtCPupKOeIILywJ9gtZh8hFb0HvyBze
twBF9luLFLVw8veDkYddtGVh9PubjpmLZm+gVjrldw2h8LcfXNsDMTcXWMggd4nB
nEkhEg3KGUYdzF9iHSQKqheLAUrUU6U3W6niAG3+PSYOjhl/EbgHVMcbr+MJsJFc
67VHe7yvfQ1xGMzWD20iHIYjoDXqXLrAEE32l3nidLnCfXkpvLMVyKUbjE2MGrDw
mUDfF90lIltt1BYJFtok+Lgs5z9hpZm+IdBh4OAwXahIxFkw5260oD2psL9Dih76
DE2QNz0I1VKrEqceN15q50kWv6e1xKviowEdXqUX7VIvTyCJpw8o+QkO0OfVsrBg
OCSv/YE1yc8wTn41hQOGQvI2a50FL5tGwvTv/yNOTGFcYviIF+4psBA/hokC5etO
eMNPSse1K3d5RRu+wF6vt2MFnZ5PXednhgOTkvFoUXcpgqoHArBGIChEWzG3pSYY
0zG3R3PmdIi93kT7IIM2FKWl+yxk0XsMW8Yhe8DJPVDxhLzI1PMnQOj+vv9bYpYA
1DgCJjC34Vn8WujKo6vSY44bYFWuC5GEXPLJcX3gUGa3jeE+IIHXhYnQMaKhP25w
6dCETrtjka8NoV67CHMlaVLPduKumD71Keym+EtHwQ66yfnJcVdeFF7w6Tdzg2FO
nShMcRUb0zyGBzLD65YQs3ukyYvSnBehtALVhf0w6FYXn8yc29Sm4bw+V5E2VU5s
m+m0lN9ApbfORmq/XH+z1jEnY5c9lNcNTGayoV5XUdKDriOEbsAuiocURqa1RcHB
pJVTJQ7jeoTvzrGW5Y5xGwErWd+eQgQQep+xy/22E2mBq028hmOyrjYLsNg7tDSb
oS/ud/P6mBCPhd8lgL0Qa6IPja5pHBFHE0NAbk1DFYW1mGeGztudTFhrZfT8vfYv
hAgjIi8jtuHhF5G4sdMQaEqMCm/kN/CNeGGbcN1sfRHtV7vwUFeuS6EXJRAXB2/8
yAZKYyiGqHBnVBOxj9vExMXeW+uJ9E4NNEcD59PiEMyzNFHLiRlLn6uQ9I7Jw7lD
z7KmHGPnM/bZ/LWkKv9dHiIf+W8YAocRAvzGTZC2JitA9DrqUroWSikloD13GIN9
+EqnnbSe0aROZWYOIdu+fxdrv6rXHtEndAbMDWjWXm0budyGp8eCEbVlzgkt/4eL
+H2O+jSqHE6mgqYshIiZ7Zk9P1LrUzhi0YV6L/mNSfJPkub/c3IcynQKHfqSIVY5
6AC+gTxJQLFMdrhWVn2iQS1X+2qIAxiT8c6NBdUgiAHvyw9JN44XkND2BtjfgtQg
wZWxiOilsgv3PFM3tvKDF2GpyF5cSzOqaCMdnQyROHZVdpxBOzf6qRfmj/cpXc1+
0tAMFcyxJEvLfCD9HXF1kQDQ5OorDtUwqgcu4MFFRLcetsTWYtq+QGIaDX3syOZM
GTuXa2dXtCGm+M2C+qx6fX29x6VL31VSpfTlq1x/nO/qWPmru3H5VJf7MSV/IK6m
UV48xb2dZ7uY7cBKmXEdhm7pQF1CUNLJLeVGxE7T1x0z38CXi2Txl7KGlsSNi9Mk
++9fy5mgo7gfN3ZjJZ8nLDlI+veR6WsMEeabnhGPjn2QsJtZ+WuSn+tPu5t+8k0y
ofsFE1qdDFcyKZsQ30XCt0IpfsRU2HB0A19UpjKNN2i2AGWfTNljB0d78LCEV48L
EmUmJprWkiHNm0FZ+/kw2NvMn1M6UURjbalTUUUgOegxZMhZ7VUVuxMX3dUun5vT
8tVDjQ0wdwxnaj65duFkZlbeR0P9Xpg+xmdGsnjLv0qTv9B0uSfsd7RJbUnBHBmg
eKSaXEHyH40vQTfmg2W2yOcxNvQw5P+RKhqBq86sMhuyKGQ4KapNr522tiE99AAG
OUrX7K+3pTcxhL/uE1pQPysBEh+FKfqcmKoy2n/CzDBYUgeZ0zuvCjm0k7G+xYWq
cSmT3Tt7bKDcyxFn2GoSIX/NwqHmZQKjOURkGR5hQMRkr5C4t/L0e5fdJWn//vrE
TLE5dvrowZAuQMS5Td19UAmxyznAidPPMDWxQ0Rz7bwZmJa/jitBHdvQLQfcPkAB
reJbAAE4HdYFvYVf6y2DJDRLd1eEuVKkMxEWVRKcUSkzKRl1z++H/4jJvEi8ebvR
0/NxJBfP/kqdUJQc2hl6dTUfHhWwckDjVXRAskjR0yV1t3ki4u9jM9qNGhDImFpB
wXR9SiBAOs+8jWIF+t8k7ZlpJwYkTlSSYnS/wFSgydL72ksrwQYgOn2ZV7xGDf20
5zH93mhXnMti+p1kfbakmAdBOQZ5hXFJFg7gIr9GJ3JPHMmiywzyeg3DrV0wJxvw
Q3sMUbci+eCSjiZGBv+zV+M3UFAhe58clhyV/49LqTzyOd6wMy+PjE5XsC/9+CUI
6AAglliuHT4fV3LQQ1XwmqnTxKOpeZfIR2gIAiyFfyLTtGSQR4yUMo++nYk8ZrlJ
h77dUt8WkOD3+1BvtdC10sQSRnYHjEywrv2hzs1GyoxgUf/n0B13x5MVLlQBMebd
jr66gYFimUNLa4G7vIuUoc/lIOfbbxX4GzzGkcaIFN+r5i9Zbr0KG2VMzoGNLU1l
A+bnFPUOUetN5J34O5U+X+jXZfO/UVaTZx9z1HTHX1YaNEDJzWHzhqbEJA+ujkdI
Hue2wyVFbbok+94+r+1TbGwNhXaTMFfLp4xSZxJv8kFkrMdDZe4tfyivbkV3zeAO
bOcIFI8RUxcpsJkvcBxNVl+WtR3fA5VlZCfzKZ6APX8GBFyN1Aa9h4jc9Wltigbo
7N6cZ+ej4INuBc619yBpGf3b8bayURJsQHXEqAJx6Ts+n2L3g8pFbBbaZvipF4RH
vWQr6eFQbo2gugRKEHEDZl+1rUrfiG3SLKMBw/bSx3OhxQrelX25c0QIV93FdTqM
R3mmwnXgudg6YNj5v10jOa9oZJrHjb8kRyk+hO6jPAjUKMiuEUM2s/Zd8v4qeQa2
LW1JjSWBTCfelw5JhFd1uMy0fLnrpAsZuMBe08gckXrF5vIelQnuplkElYAPHR9m
hlcO0A+sG/hh9IP8tOlayrsBPOc/5go3CB2Rznikc+4ObE41SYiJi8ukPuu7+8w3
KqRlpSbd91m8ZmTTQAoO+IsX8jr+R9pYUFlgGoo1+8JzpMCsh41WW4XW5NGty9N+
RpBcfpW7EUUhsu/F5tvIpAgmTiJpVh9W/nUWoBCagJ6bSg5ke3sN89DneTC+tIGe
z7fFFk1uzVRMB2XxerioJ9BnxPuOX1n3t9HqKCHATAh5qAk/6/oN5gXXXCO4hGja
VLMGy1ma3R8t8AvhqwWHOwxbHiO1lfrQKes65BfgmwNHpP+6n8LpBa0i6m/lGAeA
PGOe8iJkyxZudR7o7lz1GPEpBimFq2iKo011T8IeIqfEzxSoi1HLw8vE5vq+rlt6
+PgpS5kWfu86sK/ozE4ZsUKmcgqLKNLTH9/0nTkd/hFFUvOqrc1Zj/fiS9yYKaWQ
cYIzAvzhv/88Jw/+LneqQjmkUk5DvGJtK2w4IFJ4ZjLstyakPScojVFaEDyxzC55
p3aE0QBW6RAZejiDDvzy8WhOkBW9Szdg3vIOWEDdudYcs/QOJiKYS5OFA98V3tlF
TuaheskjtgkhcUws55mqXUdBkiVKN3dWZJQ2A+e+Wh06bhU9Ml90MrUA2Djzz/LE
PvbcqjTtslG8tw6r7dRgdoestIbQt+B5c8sMVbqNBSaTNk22cnZIBR2PIpgv4QKE
Vq0iX8Jxc0lSYcJ/6z9kFyvvSN8nxnp9bfPWxo4peidZx2vaPPaN5WXEvJkf+V31
pnnYZcYLCqGBeaxIig1bxyd0qo/tqmU/bCNE1M8r5jjUJNWXDt5Uz4cJMMiCc6d4
1v4KWpRKBbo2489BJRxKGxF/E8BDf91VNpZUO+Oa/4Xuqtok9zNxn5YlttZ4uQV6
VfNIc9b1PVNfl0GtFWOdsf1kVkI7OGHxsb/Sz/vcWzGg1THeDoRI43nOUX5AhDMc
uUtCLbjjdpvseDJZWr7bXc2s1LhUnFHIwIOCyp4NodCUsuIYHJgZMHFpVzLeiw2k
G8IFtDLIg+jGhcbMndviZVx4P/MIvxcrF7up9+ASgvvKYH23VTzE48mzrQiRdtph
Dhgy/weWHrAkFSRukHuq8WAEUbFZNYYVkHjlgtXw0c+1TonSFodFTRPy12cPKq6A
F8jTu0SU1Mo+GzBmHXw6p360Mm/EFrT9Ckd+YuzOJu0NR7mMHs1NNmqJ3SzDN9Iz
36IgEq0OS5yFDTF9FX8GlMGcuY26WJJ5gxF/Hk+nPo0D+DrDJloxEWGcTfDIe6cQ
j/zqip6L/ZL5rPotKZfCc7SR+Vuyo+73Uw8XxZ3qiWFGOLQZoyXwcK3K4M8M9ttg
DdVRypDhKHmWPuLxDbsVPDtxNqMHGGWcjzFFpB6JIzCZf6QU7T0cpJP6PqG5enu8
Ej0PrijQuqCf/VOUFJ441iUQ0XSeaWOhYFvx37/UiSKwaA4D8x5NOm1DAKrVbwLm
0VxnVvBIkCy0jmjS6rrDD5vbyoSaZ+HHud/MInDK3I4dl3QDjYfipmiTACzOi1H8
pkkx1HaE2v6Fkxc2Z1ef7kdqE81GERKwCrS+Tl0nPqSvLknv8wjWc/fLIL4oV397
W6MqWAzKcnOmOvJcN+9yv8A04cSt/sIX76740KqfGDAc17dckWVQPgHpoq7cHOfr
eQtSBtW41grq8OwL1W4lf/gzhZspzsu8tIGc93WHaScDUDaiuiHzzC+mIT0ukvTO
96j8tKV1h5ye6kA/5wfM6drAS65L8Fx12AG1o6zseofGZ5+AHKA47XMnCcrUvU6i
MzlOjkP8St1L3KUmYsfPGCKIi502EihIdxQqloIhEmQne/Qq3tLKoGKZReosyUUc
owp4Ac/Qg5JDuUn5oKH+ajPNyj8KQqRjROi/xgUQzkIKcSAjOjsAV9Jz+BNqx1s1
B3uusEctPgHHR3RvSTuKfCQak62WWCpRl+1H9SaJ0MuYKL146cnLpCADI2oXrVxr
C5q+3nas3NkHcKuKzWlUEZT2qIcf5M1afy2QglEMLOT7xYxVf2PqqgxwjAL/SWuE
Ufwl7/Rh1vvAakQuORsfTfnco02JSYFKuLjmO49z/Uj89Z4C0veegY7K715Bmw6v
G/PQKA+leVqataEafLA2M+/jcpi/jJ5CJHP/HIHrl0SZeskbO13G5gMNlXezLowK
gyea3D0O2FVjwR/kqOz1ukmSDwImvoKR4XZ2XNWXXB6awvktxOrs+aSNK5wvWcxb
nGZHzXvPuJ65h9CuG3hcsHc4AOsMjp0w7ZIBSLd50kPg0IASNaFWvOSgGFPX4756
xkWnHeoVRO46tngNVQIphiEDQ6rEkGv+f/dqtH3JdOlAGO/QMFaVI/s//TJ+VDR0
mYEZ34nKOaTB1iHeVL4k74RtvBD1PXx3hXgia9vHKbUCsyhFVymXnq0O5xhlgnn8
NneJc+DA4NpHfXbPPgIAxurwpYjlRXh85DQyxyuiKtgujHCX1zE77M0hkRWrUjfj
D6wFxr9S0m1a60VbfqvLzhIT15j4X6pM+acKQkxxEd2nc2jVhda4qdlzN/zrrBxm
zc92+ZKgwpGxDgz8EybvUM6TwTqodwhnyDKaSY03Fcnw2wpF4vSumSkYTuLJnvaS
uDB9SAvq20jXd2+soYYVwLggn9Z7PMpk9ahwniRcoBcIaDPzSD85WnOe+8ZpNr3S
cu/8svqzDpsIQfayWb+1f4IuzwZeo370kCT4PIx3GPZpJhH4kr0o/12ZbxGMFanB
n0zIdFcL3u43bCKLEuifDLGIhsV510PxNs8qxR5GvjVwiMJRT0K39gzyk9G3qizb
RbPaD4ZlzeJwzHfXEcs/Z8wsOYs6GAZLLxrWvpbyrTV4eGPtsisSYuGqYuZkJo4T
RwVkaIuU3BvXKc0/6G4QC0VxDP2w8IEXCLuta/hAqmViBXdqZMXBV480zLjTKLU8
o2rUfXpnMyjcvBUB9Lnh1m8abBxiD/dMWFEhsm10JWaNNCVeJjatmrZpieAFdLSc
2s0nueFWFJzpzwdlSeSXM2nuzrIJr45Wy23hmFEC96fUPzUsx7xtzboTqRA7vCEp
IPz8v1UOUQI4W7CYKrK1dpyDWwt0fM0BCD7uu/8zFK3n447kN4HVGxXJDl5FfWCR
pu/hYiqWqLsI4H6S0Gwy93bOCyFmHg6+0xOLmpG4uM3qFgdxzt3Ktes/cL1Y6OU6
dqAc0v1wou8b5wPoK/bFdXtp3gPxmb1ykb1PNHUuseB2HqSzYQ6ouoUIwOtU1oI7
UyCSMkT9cNZVHXLuSZJf3WlLDas01NGzenNdcZbnu0R6JSu1OCWFBcxHU/d4IXoL
iRzWQh+MzDZAjZMZxlTLEmffWbmOzfOasUzO6rTp6WVnIAjtrgCkNpGc+bOG9K0p
vYmPpVXWdG8NT8A0lrZ2uL/4hZw0fsHjeWDnSgRtO76kxto759HrKG0ULjSLvDoK
x7nFlOnqyotUoZ8wzQbWv/GPyHhKC1Dq3G4HR1TE7fsp0MUCnyqcC/z53Fc4tMQ8
unYBMprNjOxfRqzz7/83Py96BemEQJwFNSOANYsgMDyTcwPoLWJzTY+GBXv/3LY9
0V+sPks9zcCezSqjjjr3Gpxt63ga9fl1UiOwrDNhPljg3cpDfHQGvDf5ski1eK0y
aYtDa9x2RQJBSaas6sYnf4rZ9ARa7MK7p8NPZodl4NnWsOu5CSpaf2akvxur/17M
gWYBUx2DDXOyo5e2aSEArTUwbWkSKVymOP8TQ+pFChw761Esawr06kmch4hB0Mdv
fIC+AVhJMebvlruondZSpsoXDFB+OjavZgjBNvKQdj7IsfMnXu0cmr3tXTqqYZt1
1XPVWVxTC/WKcCeFbgs63toxQ3YSIBImGKbsVaVRkjrGVBMhGq0yUtlRusbVYoYC
YsiFFYaulRmKwnavaE9CqNjy24UADx4FU9CQjv0VxQVB0Oh38ck7TcSFUDEVoEoP
clchFT6IVvJBNKlFIGrferPRBTXhb0phlZXqxF5DHhityyVlJmYwLjYtpR/BTNJz
AJtugc4ir0T8oTMQ/0FmSn05VNB9CeVGaIcpkmfyid6Zunvrterq3jOCngJ027al
gLpHMEzNbkXmEVwpurwXwv8qh6qBbwYbhWmk/TkK8J3dtrGdZx4G/Oun9xUBpaM1
a4Sg9+1QdTVZkOFw5jLUkdZnm6lp9TbOC1B/5nZqDaQfy5zfau0eWTRMT3OwgdwR
/Y8UgijiZKW3pDoB0/FMzLcDbjmy9SWcnktbtaoiYf8d7jsOSqnZE57Mzj0QLkZc
7GZN/fDIDq2TcLObiD4eoIhSnN2awgpN0xmpXZx8lZP1u5X6shXgPf/dUi0Y/uw0
3jKvbV683tBc5PRPGdp1DvBWJUnxY/hpwej7nC/DmSgYaSQsaehcz3EoPOSVQmL/
mQbSEs4ofqEOwQX8mhOtVWPi21jmYOj9+rVT5e6xyFtjicTqfaSp9aZpyB6pvTJX
qx1avjyjGN5lNKi4Hv2PeYZOIb2M81ETxwc8w/nIBTbuSo2sjtWW/XJUN7CqYGMf
cjh64UDiKMCFD3yZxjnQZmLYlLk7cT0f7Cghj7T7loVzs5s1iq53K/uFCXcUhq7E
bgFyXQsW4hRw5wYziSCuGLigpzJvhtSI+26cR+ynH4J8JGmfqeM+bvmCtDPsK8sa
6ytiSS3UzL39/VdwvZCTwMpTzKHfOiWCgP5o/jdn1dT1z6aXZw4eJgpVa1yor3gV
RR6Dow5xDtEv1MBPt9xX1vqH6F4iz+jXk9j/7lGVk9VK77bLfihdeaMSc4ylSNol
nNCalbEvwcVv1lGTnPUZ9u6N4HBIg1SP3xCCmLAHgAyn4FywdvtcdLUR6YidSogf
l9w124UtT8vCc1Wh5AzusleHh+05kJBz/yayYYrA6aUHPLMFGpi7awdw+WNieaJC
4hXcYZpPGJuvOHTAsoU0vTzJbNXNU0iP2yqrUx48GNWsVnEyHX3sRjv10zxfFth2
7+th2W+xPZDNOo0hjZYrKFzOGZdTL3PS7J71QbHwHubXdu1KjmRrsnjRJsrCFxcw
SU8n9rjdzky4PaGnwEmcMqScS7pP8gOPgp+kMLmtBAg4+UBS4bXORByq17GxF2/V
WWaqTYSRcFL0Pik0rgUz52K78UGJZed0gXNm1BSzqrs6zGUURhL9pRgUMoNoXAhR
ZL8AvW5UjyVYypWt+Gc3Z0UwSo7D6WySdvKszEtxRdppjtqNPbXhzjotY75Go1Ib
ATFlu89dF0ewKGjtWt+cKJfv9rNKxRNuw57PJxSZ7l9vSxVueVbxk068mo3GtqqX
/hE6WX3/Rn09bdPokqCjtjo+Q+GupTPclU+FOT3yBzR4C0O2GLmz8DuehL3IJ5IZ
e8RnDvGM4eo5vNjyG9D6PnPUxkDvkfDkQPOsjoNPcn/IXdqAwAPNfFvbwY3gFIBA
+He1m3NpOJepy1g8xisk51QzejwS9he8SdVFddCDYVDLm7wDth0V+nUpGw27j+wv
MvwbZ+kow1dGvxlI1DOium5FyJ8k8pF4xBJNO8jREXkx/WQFh9aNzGGBQAeF1cjW
GI5ga8StvArV6XJ5ktUGSGm3wm3keLTNbPq8grVZttgFbRV4qiLtm8qNVLfdbvVx
jUzEE3uJDJrH0aqfJ2rMA5Y1lxALmFRBlXRKGA6R+jm0EvQOSucI4WB8iooDoLZU
iVYWtOOS/WCLpZ/lL69ueoHCsLTALpl3JMmOQrZp+rTXPpJDbE9mSKXp7gdorMxM
8ZQTrdkfghkpWfD2/rb9YdlET7EviRDWaIeS3OJVlrwmYNzOvQ5cGp2WAc7ug5HP
Sa7ijzsXu01a9hxgt6p6dDTXsz4rxjC4bXOsqbNZetPG+vAVFj7tzomjoOiyx0G7
lAd4Hco5+Vl7Ueyv61FvveWrU36DxpDZMBz0WAO2xPpbSQ9DivbMG13gLO1UFmL8
l30dEkEKXdZdTivpjZJBn1Ya4Hu4c16K/EnB3Ph5kHYC6LJvt7m/w3DyJ2nAI/jL
wQpbzFXB1oko9NkLQ3zWM+iigRxvDuiPn8i0UuzMhLgm+YW/kV7BfpWcqFeDnMYc
OZEfowyaG+VGq8yhrxjVMvJyzZuFM6+F/PsQYDY9BdLq7k0kih5sojW8I5+wrDdR
t3wjBaLscu0ZjvaKYL7Bm2P48jfKOvUoC/b7KZgQrCIDhAsm/GhAFho6iKupjgVz
brqWU94tXgCyvTLT60v6EonES+sGMrJUJLhE4vMec/IKKOkGazoXR8tdI2jUxdbe
qPsw4fpAwYI8WUVMtfGe7gQ5YDby/HSLqqJzf1XPzyrkl7ndE3HKKBaDnqJO3ygk
fG+otvTlMuHjX7D2uzybloZqGmHnseMJU8m0/77Y87xTeNrqla/EfevfF+cJuRtC
Z4IYxqEVi4pI0UHdPNXIPRQZ7oh1MRVhqnODWfT2ZlEoH/PkRxlINFf31FDXCj7r
hrQCF+UGFcjJE+jdsUNRx0AcWQ3z3Sn/K2QPqLkDyDcW5A/7Hppqu5nRZpQDlQod
k4vyNoi2f4YViMja7VgC9EGCIj90BW7ze4pX2UY9LKN5EGeP4IXPsfQwygNm6EnX
sWZ3t92GgZaTdPWFWRnFmeqiSFFwoILJYGC5KcfeP+bTNXhMOzC7xkUoBBGGvGbl
1whpgqH/LMbyAncIwpxWym9gRxOVFYXGTVb53VhP1NqFoapzJ75T/7WXuvYpJbgI
Xr+EBOwFXZRGElv8oeooImBOYgaC1p1Z+SL5L9y928/pfpidakE0RMQk7h28kvDr
9SeDjFd16odcdEdMmdMaIbANeebwo8FkrCMEjUwPh0gU+6HRdry7+e4K3/o/tMh9
rApzZlPXI9UAfxw9RYnMLwUlFBB41ZRR6/bZJsbOe34mU5nKQ+GrysPdc9vvrxuS
jScqD/jiSd3qFLbny+0ZeRzesRIfnR8rQC5MndLG23PiZJxxia3YnKRGclwK0NVg
Km4dcHBV48/JLJm9LYVQvYToRlROdJ4K/QzKPEMopM0XeXbGw2zV9gEF+IHPQM+9
0dzBd6DJ5PHAt9av3c5bpK6GY8MqIGcL9z4vtYhR8+/C6pe2r3zaJXzAeq8LmAeO
PxmneWhUucf4Nnrz/wIckPoOmaS/Bj5MomvkA31b3eaAVlYoD4f2EUstkl1g6rZg
K6TakLtGoGpV93tc1rv35STBWZdFH6oaw/9mRrqWb/cx/FHi0TOzeeF/LLERsr2R
iwa9c47qZnwjYbU/8R2XhStriEKT+NBSdFBGFzCw40EPuAHsZr0HqUQxqe5k5VXQ
Tj9KPSwZzCr97A4PYe0c7FEoBt80EiJPIbGxlp9yGC61XDecFoUXiQy9mr0RBUOx
vVCsal9clHbQIQlVePzIvcALThbrE32+WsmfZXNYQ2YB6p0yJBzxilcoesISfxGK
aVvvNwI9IS9dvHaZCtGlLDhopQKnFJ0YQpgHq71q3bEg7J5wQ4xUtOD+MCJCnoth
rdikc3ymc8y6f8gAaXdD8Rf30WNIFqHi0ROe+R9Nwczlta52FPxaT5su1BQ+8T0b
cZCEmkAer6ySx0wTbSmfviF6I9eVAFwk7Jf177HPpwnTjEaNKhZ7zhl8Lh+QWjWV
BGNCEFanwNsXdHX80p0lfNbYDR7f1em934uyYowZjZ/RneYzml8vmmDPvmI5WtYj
50cJpjbxYzQrHUuDnBFZT1O8GJAOJYawb2tLMDMD/jJj1z6SD2AjvyJFGK7qa+cB
RoKEhY/qqvkgeiWE3reZEUX8FqfAHJP7rx+nNvrcgkZeIMxB38k5ea2l+yN9AbOV
xIOa3WA8sr2mwRsEl2ZCuYF3ROjRKU5Pe5MvY8N4vWlVgtvXtYfPBJhEhXa5gvc7
neDyxHqnccGiec2P3XS7jlRkPBdVbYo4g1K2dGSRp92MeH2Qf8DTY8azOqYD6z2k
/MK7Esgq5bgmUpyn95y3TuMAKWYwtaqTAmOL3z/o4gBCa9RlOMsXkv7Hbxzpjm/p
loWA3gu35u4dHNjYiMmgky/Na26hlPElY0x4aHRTKaS9l9Iv8vt4nJLCLhrEVQbz
KwG+ZQwRyeMNOQndlD3EnxFTHvtALlkVRb+dMZ/NtdZtB3uzH4L1YblCs9xB69Rd
1zU0mox9GMw99hshR3VRAI3hkqPVve3s3bwp6bAANIPOWfGRBN1xsoL3dQLBT6sp
B3QtB3VmsduTrg+mLnQSWNU4UMqmOzqO7zJlxKwjzDTAy/FqPIsXZfSh+Tx0wcB6
oHRnh9KTy1UU7jchW0eNqQ3R3tBuMOYqIdO08I6vCNMp5q0KkER61MhA6igqUfUK
FPc95TCuThDUb8kUvK3a3k3g/qOHChJ/gOQVgc+YEm8TPrxAPwwR7o9JGMWdMIrp
xbj2oi/VJK6ArtzhRH+aJuCdtlmLmrW+dS/MvldWG1p7fh6KEz0fIaqF1+tHAhRv
nrVI8v4TEJwz3acUE0R1WIHIOa7u9QeGPWLneMo1cqqngapuSAPkjk2mjInzGB12
JDR1D3Ykc/xeIS5QSoLoOnUC0xHu/BGZfR2M7RL8Nytt5d32vTPpy9czBwBTGC7h
/n3Ui9mPQRxper+D3Pyt95JKbERYWYSaJBAbr3n1hRuC5hHrwpIfSVLgQxI7ftmi
C/wlztsKpxGtJaj5soQenv2rst64a/Pe5BTKpBPsvmY5BuMaVieg1JUP8hO46hzD
M/FZoAJ0BigFGheqf8V/rWs4TaEsaDDUjIhzeyT8sZTUcZrYHKLWiiUuIQ6mm6Iu
SazR2VWg8J6j7GraCFwPrbhxfMwmMXuZcMCsap2IP+K9rebdhPMchwvxwlncOIfs
XJbLWhgiOJ7QxoVGUipwv9BYch5eJHHkwpq84piQP2OlljsOlxphLidJFqcLPhyU
MrXwZHMlfz2P3WIKwCDAZYlm4GxYbXrf8NzDnSlCtnH7fJ2c8lxEFZcO9WkCgwKn
GX4odTobAm1ps+fIIdBmPIOiWBE0TXaRcR7eq1W20/9oDqQu9XwmfyAdmeetTR2z
tRxF9/gPSgKtcJ/90YfYYp65Ny+ySdC9CXTrp93PobPwHTPKHZSnSEkAnzGElrse
TRPevNBIe195gW8i7XzVQ0WPt96N0tTbRdYZt4lW8jCseZ2Abzp+OOrbtAaYAmKE
DAzW/nKkxixPi41VLJaQVeN+bN9L6t96LTP/8W0G2PVdaC/hp59JijddUWFtFJZv
DtA297dGxsZK+ehtgjMvSa/Myn3ZWl9HCo8moBXt77PSpzQfci7yQq9jDoN0EIGW
K31SrMxooRnEvFdpenrTqOEiJ07BVUQQo/0cES8o4h+8JxCN2HqJhjbvPg0Kmxns
AORcmyuVpzsxtRl/n+tWPNLv1w04NGWdhY3as371+58I7f2m184jb9BYfYe6ox2Y
lacKhHCSMv3OgXhBrLYH8eg+8uI//oqVGVYwsR42GqJHLKUQCm5y2tpJsxFiP2f1
JdindmnHDIRdu5/G3CwsmWN8vIfktQBkljiQUwwRmAhnb/q2hgrlsl9kHX65mNLk
8AXya14laNKd7o92SaR/XsDHqjoTD5WXKn/2CfCHyNJj6vJbJhIWu1BYEp+zcBXE
LDRIHhgXZnIBbwTIM66xx6HASg4zNZNwEQ+btuH/zlPOIKIzNuEQ8ffiu2Tyi/Ef
lvlfo3YMgngEPSHY5sdqwtvgejrMRYjehcDwreuWpMnHu6wlP5evT9qsGYpHxJEV
4cgySGfPzg9vTaRvlv0/rLPXrSNfJFXWBNS1dhM4aNJyjKih4yTjnLGl3O18Npgw
Xd8Cw0monjE5mYh4huBQKoiU+6yRkiir5DBYAbGa3iruLagQN98mswc5UzxCRZhk
//ZiJwQp/k2xiN8IsxK/YwbL/jy99pnrGkwOgrLF+3tDvU6gaviKJXTHO/QK86yh
PoasOsvURfSboCl2rCsYdyzMOEu6z7Xk7IjrtXRwA5fOYk/8cJkOPlDCy2VdR+3B
Ub/3jvMmqbYvKjCLVEaW19BKIoPR35cuMMU9EdKnhTWd+R/6PKKNaO0MZ+XpeHN4
vhGIDfGVNowExtfpzL8GJneWR5u8NTgN++Bams5sw+qbmXKXdbOJhK5oGN9TTVU7
8iQ3FweKgm0C9Y1vH1xIq3UKoQaN405sp5GGIJlfwuctUGflIxusbWLgnU30ccJP
cwyXb6wQcUPhTHJZlXe4JLyXJ32Ac0aKbF1d9Je6Dw33ZqJfavHgpOAQ9DnWiqef
4INtokjOtCHW3qzPXXnCiX4RZ0OfK3t54b21tf5sdWViSEFCjHpMfTXLSgBCIxBe
Mp1ONs/U69ZwjQ/MCOV+QCqr0x0qaW2PVYclGhWSRN6z/CEVei8xrsSk2F7LuSzi
d577iyQMfbkHbieldH+5etdf77hDKSrEcuZqGSDRqZBKKj1u6IfURz33PR/gCNt0
TshMWBYY9CZFbCsKhc+h1tnkjv/dJj5j/iQsvD0MFgisHZGTKM/zBIBUu1k7H5cK
NglkD++Ex+2vRYtWzJTmkCOGfzWOEcTHcd2tHz8iKRj+usleLucirCBSowZT4RK9
qzOceKsrSqpkKT/vRVZb/3WRyBMnRaSTs0t89Z2K6XVaRGAYrW1BHtANrZKgXjiX
rOrUzJ0wrtnUwdOQ9rZh72U7WnvvAu5K4uKOIL2uI7uDIUrWj9oRBUQgyv22B7Mh
3QJVI7a6qdd+SIUEwQA2l7QlbVVaZInFHdldCt2Ykqp910RwyWSoA0cYL1lbT40O
Iwoy44mrW2MDjoaAjZeK13L0ZqNathNmYabnxn5qhz3YfuTrNOTKu6SnOs91oVHE
Ya4ESgHvsFN5+sqcqwSqmg63Aus3Bi7esIhkQA4sj10EMdZaTmQaddIawYGI3skV
gLmB+sTv9igikPJ8oBfWKz3rfef6wZ4GNUtLCcisVFy3lEa8MM6JEm9gW2InHRCc
VufoE/JzIZbLt5vGBxthAUghDXe2C7PP84DUxTqyhyno2pdsEjze0+c4kTzeAGEP
vfzNi3UJsRkDOCQW0ktuk46REYevdBteDJjvZaSklmHbrCmuGcEy8r3wP8TC2u+X
WhlPuRi9zZzAcmH80OwWooP+O4SSzh+fI1H7SazyRqVR7TlW0bbk66fBLPNI9j0y
TCP2R0HgkpKg4+wTcNt2PNJ+lFJG36DRTyZroZ43o8y+oi9gYZ/Z3VpDEGqzv7hm
vF6lxMRPLybZUBdeY48mHN9H2DPamgHvQScPhLNRmqtEZIwjWLKZbpONwYwevdiK
R8DYuQH/XLritI0yw/UqtptcVciN5KcpSeePktEZ5QnClCA6hmwfSkPTEja2aUcV
Y4wvJyKDc9aWjhcH8ycG7p6EyBnDdYIep06S4o4G47i+oNOzg7O2N3dlEG3+H10L
e6rnn4yADJON0YxhJW+1HQUH9MrIoPab3fwIDX+uE6+1/dAwbT08E1EpFc+XH11Y
byQPijb4a3kZ60lXon0ScStAHh+59RwoEJBqXGGnXDQVfZNs4Bw8Tfmtz66lj1eL
Wd1txX7wedZcE6y7zVFzPJV0lbycbPcgCSgdLsXt8n9zFpjfsCWl3Xvh/OTbChZt
UfVsUohLwKb/jPy/o3UswNpiCVUiVOheXy4SshC3dIitGhHKytYvpHGTPCgarVuV
625IyqBrNj3Cb2DKxVqWpj2K/Ak158nNhaUh7JykQpp2l1XZfoMClVNuCfpLhM6K
SN8MKdC/OFmq3eBNbZT2aJTMKt2aDZZ9382In/UvzoZ3/pw1AUM6cI/GmG1Na+7U
jMJefKa1Kcb1olCzCsg+hoW9uiv/dDptHA8hhpgDBrK4KvOBgnKXcl6H92zIVNfC
9NzQVp5h09UCthn2giM79Vktcqwc7CYpjMsdm+X81lrhtaJcAwRSCQJp5SNvOszq
QeY0J4WRI3RVZMJzSy/OFnmBP4UAuiOQA4fYhvPB5418VJDfT/72DAuWBHmqEgkv
8LIhoeIDaPSN0LTZuqfYidRYWOjoiska3EU5i+i6Xe5ME8vnjqkzLnoFf9PyGLkN
C0z5XNnshU+nFSZIS83x2ZpZcl5q5o5YokTJJVqa2HSlBsR/WNtd5Ym8xEdF46Fa
BEWmQvp2YmwLRF7uxbeb/H2eMy+W6U2PzEZCpFnoiNCgQTpHFPtemfXJxg9jF2kr
rvxYdknyJ5hKV+gpUDBRalo2hAxTErN9kdVbAbUCdVKHlOKrolwxKzFi3ExZLGfY
YT4XpiL3SMP78VfpU9aHZks+Cg+AdalcrCT3Jpk/dyahM8j9r9x7e889cqb73sNw
60Urwnp1ZulzkQA4JwdeExHZcO9GlnDkvvX6ADl30KM8Oea5jbYpndkextQtG62y
r/bGMX/Q8zTzxwuF81JGkB94wMdFyE0xyV0KVG+vGF/qNmn7TIxLhu64MjOIaz5d
+e3DX+6mCBQern89Mw1FzT2wboLVDDgBgMhKcFxERahnHInaz/EONs4APUATSjzZ
YeX5vVeIV4/mzHtb47W02D+lEmRjuOpSdHh4cq7rYaG6icvGAnW7P+F+6HE0nif1
4UrtOlP9yxejoN0BbPJcyMaAt76BzH2zAFfvQS8LIBOda76/aztPsz4QpLqJKx10
1SiMFLc0da4+fgGBYUAJUF+zr9zZvnJzn+5PaMj0W32F9LYB50pa36rOcK/sc0Tw
NW0HKKMPKEQGjmQlwgNT9U/it2+HZ0AruYydQw4nmknvk1MuxH6gjGf4G/40BFvs
xyiN9cxhBhqzFhUbWdl983BVl87DxVbqWVo6fxKt9mzhlamOc82keLJKtfKw5Fhz
lElrg2Qn17afVTz9vJEU1G1DaxEDqM1Rxr660+lYwGdKNVSutUpWL3BY0YpSrWVz
RIaVCL0pg0IX4z9tN5oyUGFLYGFTY69rGru9HDlvskp4eAixR/G7RvEGokJ4qBWK
DQFBPwkZ1S4VDY46wLlzx91qjufBSMrE0YJSUNs+k6Cq72xE3Z909IabNL0KsEgB
xnkqzKaRNTvjMTQLXiLBfl34Rw8hFuQQIoV1PRnmH5ydB6TfvsumYpl6m7gCG/DI
NhShVU3AezSX9r4/Ui2/zKOPkKqTErs+2pBNzv9nwVJsyEmnatrfUn0h2tO8QDYW
cf2qANzuIz11q8APS3xaCL0w1GQLi23uucgMuE+KV8RBpmnGR9NOYFQGwOdpJVzN
EgA1LFDWM2Q+CdxF9j1/u6+OeH/uPrfdUw7b0eJHOZcIZNdbd7yC2RxfBW/itBCW
3zRD6KVQB5JnqdEaMe1NVIpQmaZOz4G89Zk1MDS95jscLG86Scp6sk6+Ik4Q+WpJ
t2gYmiyaTcYuprtau2aTGRzPaoUiJhDafn7xiqGzicOuGqDXSnZLo1ncQ5yo/qzB
GqzXD6IhlYxraquE4Hsxj4LGYIFti+SB1WhlQcp1nzJVNXRU7elihmusb/Uut1Tf
VeFMuTvJqf7abmUyFBjAZNZGm989FEzyS3wqmxcTCiZEpMZL/ccjLcfkOP5+l1Ko
aPsz3J3D06K509IY6hM5Yx1ym8F2VTpgLpJQqB+9/q8Z+wWOYQDG+AcNUbnB5XKd
b64vdq+4+cVBV/bWONdka8Cvx/kIV3Q5p43jhfN1Kw+HvTgS6pjAll+TRRgCmhFw
9JkqynyiP1Sucd0e1FB+i0RS9HiJApgr/v8XXZ79iiG/pt0L+qSAenEFp9AE0p9A
OqYzmDyLbjAckaNqzSTJ3st8EydFSeeEsQTHvnJkz7CcHXbS2DCtn6hH+AZBqToj
Cw9LOAaBuk8nlll9p/Hy4IlYpXo84MBbMkduaIPC0EA5z3MatC+Wg7vfgs0KNzsP
xmhISCbrmS4yrofeGFGm7eGW7RdksGOziP3Cx2Lkvlmp+MUsJrOtvjiNY6WY0wC7
PofYFpAfF7ttLZccyZWhTGYJGIMpQo56yFEVg6iTV1A/iRUjV4VXlrPMYMLnmE77
pUbpcP38uPICTaYAb17MbKO11ouNLXiHKWCmlxL5SrNHsmiD9hSDvBXjGG0CYW/9
/V+FTQaAvs7j1kgUzvTOIU2UnNoSi8C7Sx6TOfCXVRCgXcdpy+89FQwSYE77KI/N
JotoGnI69mir4OX1hLJ4XeXIy88Kuivj5BFe9O+ai1mVOCzUMuOruM8+TpSjDjKB
rKetU7vlEjQmaenLq7RpWenS8fBjoxKW28iuX/g7SEC5MXh56zDpDVB1uybC3tKZ
y/VL9XQCCbzjwnXjkDIVhva3qSkEejlkzE7FYkuwbeDW/6KSjWxMnyJiht+edCBL
rHzICGgIOd6fu2hPvWITGHOIePKw6AWBt564dUJxXVXbeRTRXgrVWfDVhiNne/hW
JJCPgWmdVksjWK2VmNQhciMstNTJ6FCfM/dUF6wPseuAhHuIs8xLEFiv4UHcmsPb
tRSx2zYlsjn419lbgtMaOzR+IyXHLWG9XWVytX2Ih4NY/hywuDHOUaUp+KtpfDEC
LWHjPyasxR1n+lR2yKIZ8OKTFqofW6Tt4008qia1aOCtndNZtycwADM2ivE3IHbC
HvJFccRWFk0FvFt+VPRHLXWNaup/bksdQJzte7s4/1vloKVKGulYh2xj3plpNAL8
McRqQYR+zLXJd8cV09grq9Oz81ngVDO6qOhTAQxHTIcX3vnnf/9TlflDL1QA0/we
GtYe7P/TolH8gktGXPstXOBhmkpZpQdoxaDPJSxqupwcBMkFsmXMlHmzIesMRTQG
h3XvvIS0NpcqBpm9fU0nHbwwDqXErzxYORCEH6xkbUVJmpTZJRO7EOO5CJEOf1Ry
iC7f0HjAea9PODADs62C8cgs0obcGm5CuwypQ0295vt6YRdyPcufxWPlmZy6BVOW
hNeKmpVK1W8jiIALiEKTE1FbHpiWH8Vu4XdnNfNSaO8hiyaxmoxY+5HlrbhiL6W+
1kEfCwBTjO82OZ4fWKEd2NrC5I6KA4CgaKlffqbfti2Ju+vNa5WbaGz5VP2BH9Ev
rVT0xFP/umzXJ4Z8IbNcypnIxfNYj6zDoYRzk7+8nCnKhImRXLf0AetaP/Ee92ey
BH4SJTOM0nm80Lplf9Cd/XLbGIV5/LYqkjJ+uk4zMQzI+MJbnEz/hzxtopng9yXh
9z1kw5UTz8ik350a8kgTxAZZ210eBHC9ttc8Xgu47zoZivCmTfwoWi7lYjax8KCF
bJvlAGZVylFnt4H8Okpmj4cpkaNtFKeaFy8jiou5Yu1MEmsue1+JmrP0KJAUI94G
1tvMl1iOv6akruM4Btx34ga5V0UoQZQDxpzHhGhlUnZQY2n9/m9LHA8QHYMYaLkF
fyUWnlP+zpr6eaNYFGZMy/SvNRJ5BjImyiKxZrnFS9xBUgk3h6JrVsrI6187i3SZ
6ypBNEbU98CF+m0bPofgR/t8rdnnvqGIDYFZhq9QzS3EnvtRlho5E08EmDhGCdmO
ZQe8moWiimuw/pd3r+zTzwxq0V13V387lsRbxjDxj562DKwfLJFJ5uQRQyl1wKFs
LGG+gk4pXrJpQIdQJPg1Jf0MegnKXYzHyaSJkr9NKjKlxjhTfQxLACXulxy50fSt
THib53NtVs/F4hvPwBhf1K8afTSbdXLdlun/B683eWXEqqU4QgHivOAreQaYkMeo
KeZjzUPwBreprCV8bPCYMQzbyiUnlP2lFdLtiE7x556+N0uoULfP5PhCDpYNAaua
cBtk3sCMXDgaFK7z4lzdMe3G8Ev2+w6C6p93RgkiKWswbt/m2nItrYPkviOKO+n0
IUsNQ4Zq/lK/oRNS6A6i6a6qXLu1x1MhlOTjeQyby9fNHPs5Y9VwaQChw5ulHEv/
7Jcz7GdVRVZf862vdy5pAr7uo1IiGkcZpFSjxSqUFz6ZgHerFUowHA3jmhWHBTAF
AvfZ/PKoah9AAKbb4ENLdddPF8hQUndj/yJg2mwJcqSZzjH5KW24ZJBh+2JVbz1P
ds3cBOu3B3lNbhIyAav1Q863GRVoWr8uJJ8p7BLOUE7maLM9Eir/hXk6fEK/XbcE
8RwxQdndfV+SafxzxNyiPK1XbXf9l/Ba6aD11+3lyvsbAliAbY0gLaq84ZCTtElZ
KvbQ5xv4j28GZWRZqBSoHzsW6qYIeennHRHouEn2xUpotucWrHVQUEIDt+ZzQwUw
/Mg6BqIjLpGTA2DBaDQi/SQQ6NjGy9oDopdmi60kkZB7P9m6vW7tPiRhxA+OXvy2
xO6POpXZ9HjeIvRLtuYirRXyumQZ6PSDIAmRzbQizGV+tRmFG7VS2sWAu68hUOq0
BDEEg0Hoj7smmjF90WeW5qO4fOksoBV38U3cVIzHXhx2Ibvmt5YCoFhF3LJa9ind
LmZiDiyp72OFK4Qc2BE8g4GZqi185NZDJM7JQ46DCB0q/+mnVB3EyYTK8TyrV+tI
jnC/rSphdDtDB6RUpsK0Q+2jbJ38CwzSDbmRYZO44CRrRDsKZBGO9xRIWpI+QR4j
a5Ql1RP4g5mx2InWmPdOXho6DE7mv3XAkL189aPzJfV6/TDLc5wHTi9EQKyVgwYU
XluVOFnMLik+myqioIVqavj11tZy5+TphjDYMn58Gob09tpeYwxk7aj1M5EPkF89
AkaB49dmH0xj08fTM5st6p+2nawr27AdSMtwsznA4CYuYlu62+i/pWmFw+Iypm1J
483MnEno+EaJgpUGOF+Bi7gDrXMOBxaZWjhQtvqoz6Sev32O0m4snhCkJ6lt/SSw
kW/lhU8UpXVwwltAQ3lloTkk7N/IOY6iRUARho2iZji+irmhaCrRSZkv+zR3i2UX
om3XF4tVtKJXHakvamvrBm9/w2/NLadJTorq5h0rvJD9YBUKpNuCMHq/A+tM3On3
lqTWXNYfkaUMWCz7RHDCoQ10Q61aQKX0XgjHFyQ/czmmDxNeIAvbN6IV93JrYD9m
zVmoAsaStN5wjeIyNDrXYqh4ObNW0EZGWadMSDqE49pS0wuVFe6VSD6Iawz+4eMw
3FwMbNZBUEMg8LbEsdnoVViFHvoNivi5FMugSrqhElfqrPKH8mpMrMsJdFHC33IG
MeKgo3CUqaBP3nrq4zecZ+QI1HMjGUq+ZMv8ec51YoMRXoGrPesZ8HHsYI2y/3C6
2Gaq1Juw4la2g1lp42Q7U48YPGU6t5gacue3B0FpFvj82u15jUEce4iAAlKEtzEy
e+TGrRfQ9SiHgpxh+0zjYzg6qykqt8UTAPn1dFK7EozkTlCzQzLs/lpVIhw3ZrWu
Ov1IOMGRcI9K2viW0n7gd+5tlhN8br3jam97L22JMovg9m+5N3mt490R995Id8Y+
sRuyG+TV7TsRn37OlSjC7UH6c10FjFZ3p2j+6Cs83899b3s6CQjUV7Hv46A/SWsF
WI57xVYXdH4KT1LqAk5bZKuY+zx4X7mtS2eMK7p6Wi5UnaJbbNezQjc4rQbJdHl4
+CoVMKbeY+hs/mVkKLKR9Tk0huNN8jC2+ThvSXBo2j1JgMugvfasDsi3DIEKkR9A
+95k55W+kcLjQg9+tzY1w2e3cXUci8AtQIh/B00gedXIqBDlcoE4QSTW7GFmHALh
OhMZayAhZL2aV/T+SfprB1RbuR9ABrHBBTbnW4Mv0IFbCbLoi0bxZpcivMB9CSnd
13smzp2keF5IDR1io1E7ONrkqbRphttTLpZghby8nGSDLopqWGvXyA4arKQINn4U
bdvkoKkqeosuaSOLQlN5/lNPs2M974MuYFwWI4rjg3WbIOTtP1zFnWpyF1Z8P/Ap
hlj+h2BSSzDnEmPp9iaqahOCs15jmiDPkVvy6yYKENZL9TOfjbhFw7jrivuhsXd/
I3C6GA2Qh2FC+WKMItXrSb/MAMy1UjF2UMWbpFO/9m1zurnW0gqFCYJjQ5HR0XUE
h3ZKdGbCDAV0sXyXfIGYSb6+OlHlrDoIv+o4XGqQEmmSVlq/Xw0kwPhdsU4eTGo/
QilEVj0uDjRzOCjoZdylzF3cvGI33gJ2a4Ks/apjTUVF2XQyGay+Mde02Lh3sHH6
1ZC9iTeYSz2l0xmcWyPmNFribY6zcIJexML65i9OSkZMQEX2Rfc2t0Bb0rLBFDwS
BLMslo7C+fjY7ALcRnrXEeb11oG3PMqtlM9FeNx01wOTS1l6/MN/gR+zC6Tpzrr3
yu724Q/sTdy99pjkCGN19CZjnTXsSTOhJx4oOfD36EydiX+s7AIuoVjTk+cC4FbX
UjMlbOLZ1FSLyxvin38jqd18J0LaKDwygfFXrsX+1AOk3SOPBZue4Fsa24HzutSH
8GVZ3ij17Zpzws+BZrqXZ7yjF+1ntKMfVNXAHKgxvU1HdS2dTrZzL3yMh6S1vslk
XKcZnhersHO6gpRKzeT2c9JG/nWubp1nJPn/0Rd/hHM41lEQwUWOLbBj/eJjOifx
sLy24JeD6+m6eZNpvA8fVAGkD8gL7aEr4XKuUk9+r0lt/klvP0V3Khz4RNi1+fF1
2wOI1UPDxoKn3++Y71eVrbC7STyKXjRmkhjzNWUYCmz8i27TJ0XDKeg+7uf4eYlq
zTFBJOk/DRYy5+qgmFv+QWyCFGLlA1/5the7BW5wDQncBMg5qrowPSbZUViZSPtv
BXH1fEHiMLW22hHW3UBlJs6Z9oOu5vdcxRWmyEus8wq+v7ASs4v3jvfbcOHkBmpZ
CV0va8faLEmyjCMq/GP2gwLXCUHV7U0MplnsAUEHePPC/lNsUzDpsk+oAOzy9moz
4otMGqObrZMvhL2PosYfiM4/nmig7tMTl6kXSMN4FvK5f80/ORhN8TpKHaQXdPJg
KZPNCwVh2vhnJrmcPEb1ZyBr4gECrGYH0QBxbKbjs16GbF9a2PTRQDircuzWQu86
j+NKWwNqjIsKBHw+0D5Dz3iAiOZ077BFrXxgNx0xJSc/yi1qqoQerYQ8eceaBZur
DUrgqcVERTXx2s1DEkxw7dAWM63hOijV3+Q+7JgDzH0Cv7Nl7pRvUjtSDAIcrVF4
gi4o5Q76TGqeZIBjBzrX8EvRKaxYy1WVT4h+KubytIHzEFudXORKAkEtobHKw0ei
EQ6kAuDIcOjeJl3BuqhCEvTJ/40+i+yBy2bL2QdHP4VgvBl5gSY/rCwTKyMJvwuv
iFneAgsag7mD0KWQ7IptMKyG9q9OIegGkpYaVWIJ7zHgKYQkgPqMGCXrpu7mPSQt
2A4/kaBqP/QwKTEJCacxfj6u3/DBYQQDU4jtLBUj5ktO7s2n3DpDOkHN27hU4f1F
iVEAxnBF0eK7BA6KUg6P/V18pZi/HlwN4qOgJnabg7MoYnzxRrdjBgaQydIeW2o4
x6H87B1g9ekzz22lW/pqsAy0K0CWUZzNahaVgH6Sku5R+IFrlUjGZwHIUMm04/fE
QfCCTNZ6GbwiIH3m+yBHAn8NUNQW41DvVfPWWVmaEA1jGTfCeK7/Oi5EeQ9v5C31
xH3k79e5Yr9JtpQ4TvewcCo1kejdHxnJSvAt3brR/I0eqDPq6pG5eWuUjTv5YwQI
hLHqE6N+smhbWxbCx2txYRxN3jo72f3wpezvZob6VUtMnXxQcpkCUS505nCLZKAK
RFJCZDbW4es93aZQslrXR9n8ykh01X56oSkbQbaKcDt9ZVVnYbiKHnfa8C6O0XKe
xm83I9T4rFYlfibMhSnzjhTka5xM9uoChQQkEVtfKvHQeU1lfS6+bfW8mMPq++8J
7eVSLmFyYUWDGaUAoP3NHbs+7DLugbvxUpM7KHuwaeVEOCESeaZqf0ruFtTofAio
OkWBskWRIFD2Npj3qwFAUdF/fEGi9ecXAlz5GcvsLZWTTVbmtPm03kAunspYBNFP
/MxeAWkRffN/bywgqpimOOSaN70t4QC3nSKurkiUgMrw1XYrSBtn/7RNKazkqxQq
kGMMUHNYTbcSDqsI2E/L+xuQUN/2fn+LfxMv9R5qqvBmI2JXxMOe2SU69qLVpTW8
jZOSIizGWsopu+AQsvwKWXzLclLOuw4ZbXVIlJ8gzuSQu9NwQnx36QpFlj22CfAh
21tU0XjATF4INTgKAySenkxAujAKd8om9kldkSFJxwQx6XfYbZJdBUGzAx+lP1jW
+whNxV4Rb6aKBSlhHUi199RHkd/S33gSTkFHwQcS3ZWql4N94peHpi4tqhzNoZom
zBJ+NJnsa0Qt6QiqXYiHjBKtC87LLDJ5gQWxALKrQUM1cbGagLvvliJhbPF0pSUU
QJGeLO2lKByS4sdYbMQgs8kD+F3qySl8QrgaqT26EJ3R7QgRSvYFxN+f68O80KVk
2jURDv0kVhnydfWMuRNQQ0N5EL2wFYXfSfwO9UG96U7J35Fd1L8oKa2KoGD8loF6
8gZd/rVDvwzjE7FvOGlY0GJ7TBkjKO2CLBoVDcH1oqI+uwwVXGxlmwGmNiGjcfJG
YOxzE8TcnXFD3T6FQsFTkyOmAkLGuDgCpTEEC9xsOkqocTOlrnUiE3I9aZ/4KkNC
y23FhATf98x7bNcYFx9nlScjQQamrfKDa6J10h4PeNUKF7KosFsRIhQZZXREi8Kw
KlodklGZDIZdkA2MXnKY5n8onBVOH2dcE8gaoQvBrqDO10CfMbrVLfulPcTP1BA1
ry9uPugQwbDvTBIiqeGSynGB9XTCHO/8qliVTP8gk7/J7WTZLWCO6cwHNsoVtI+t
2U/B4KhE6QdKxNHzDloA7OaFJXGdgaL3Tom7v7WVxtMacNWTakabkn353LErjC0n
xBhA0Kk2NqATx0j/bvMoWFk2WcqI8ow0jFEUmKySabzCotoDNCfNUKVD2n2Dpd+c
x5bBGeyvPhZKJj9WYKXuC51Iv9P1PRcJMF6wp+UHWxTpM3wXOt4HxiOPfSTq9BT1
cjFvZyTtlppGyjrL1NxGuauYPOW1BqQ/Sp/CioCDBbYFxomsXOtWgXnJcETyeS/W
6drhHfIbsatM0uBZ2lhjjl/rF/SmU9nImDlTepiRkNw53ZqC8MNtZnERbIV/KVAd
kiM1QLYZfY/ubRN5VnJa2y79tS3D+1q3mcFskY1oH3fllfKd1tNxFSsxkm6hysWp
7U4SRn9MOm05jvQuWPasGke3L+//IFiKVYWYYYcZIE5kAVOKYUpgZm0jnjlsdHks
20A9TXerOq7CL3QkOWkr/M32mf/2QAN5E47ixpr2O08PN68JvGA6l0Q0xONwCIWr
M4mMNBP4AwixB7H3Obj3xhGzrv8GcW8a+M2P9lyASHCCwXEl/jAFFXVnw9S1lnZu
ZV7sel98fqrxz7v0fiTg14Ld3XH0JWUmklgTlPq+4iZk5W5yzr0PXkISCD0xWXNI
lMHsR68n+inVvjjyvvEAiaefZQ0Nlxj69WLfGFMboCliYr7AYyGobu6EhaxhU6N0
+LIB6tQR6Z00i3cRp4LO75SBi6ChqKRQPMa/xguxnCkHwmz0Q6kijLXN/9Tj6Hd+
PglAdOqTUYf6T6/xpyugql2M6umtJoRiGnIaniRvau+MrzUVOZqiYcNSPcp2KgKi
6AG17RAjXE5gKdorsYSydAn9vPIZdxshpU3eYhPd/fGZ1ZBiapm7iu2UCv1ELE3T
LrbkLTozOLQpd/TLaR0Ku4tw/wvwB1PBDyspwZhLNc3Q4ltvrcsz3OoCP1huNt94
wWEEMKvv88Zdno+uSQ/d8TRpdWnBcV3rl5MCy8Tdrm++0eScPhPuVGYjN6qZbaac
oS24Up7unD3/1a0Wt4Xb3/i9ZEqHpGNxFOmtQvqEoQBTY8XXseu/eoYTxxBpuIvg
6mCMyUdYat8/aN3XxKx0tZlR0xYOS4AoRYiaaN07FjoAIkI5W31OhwMAoPS969bu
qY4jBriaSMOUZC55/DkvH1fJG0HsCI1Xo4Ys3EW7SwuwWvDgp0Q02iKWaXgWUpbo
HvjXT4z0gUznz1zPaoMP1Z7UFfpvxTJYRFdDVMzSRzP7JbYQ9x7cKk6f71k9Oo2b
cKr3mn0iy0XmjXqQcP6bln7DRR6LcAgruaMM+TN5RNy8almFZ9iS5qPERPlzMTwW
ACwnIk+wn+jh8lJ/6YBnBBG29e+e2lLPYk5B0U4vuupAoQYrMvI0HkLGZUmVBFvP
+D5Arj1h1nCw75E9lqv1l9eFQ/ArzuywXEtUxBRikroPNS79td1CJjjwBdFIXbAQ
RAjzdIQwVRqKnZfNDfGcYNRHXTTZ5Xp5TEh+Sg0ei5QLa1ZnlQRuLzMIGS3B2ZPe
7l7k7g5gJ53Hix7/FI4K54zVN4vHA1ntFZdqtIKLNiX6eKB8UbjE1vN0zTQiau5+
TOBM/FXq54VwH4bYhbPf19Ts0VKzu7TqL3hq314y3bK3wtzXWVMw63UNkNM9kDin
xokxck/ulBRQ4BICXNVgnO/5hhIDs87Q0GaiRHF7tT8xCNVjywyGZWuXeKSl+KV0
J7pZJ13Uiwf84MNTGLi31tDObDyN21wC1Dy+JrCMpTX9jCXAfLzGL0g1JsUc/rfp
0Z94KAsTFdUZyKY3vZzuLcySuJ1wffCqZ600GJifsYyqob8DUrvsrrNAF0rXiRF5
owywk8ZaZxNR9UqEKq55UAXbu+qKiwn2g0a/wyIDWBD9pxctwdc5kXWKCWtrsUXp
B0vt5KrRlsS4250lB5zRKTkPe9Ql954HOpFL52fYzlQWdpE2y3Bx8h4DB/mG8Phc
rsKJJdqJpr8OIm/53EpHbPD0c2VV3ttBxfYLBGZ98TodFgP5F6bGckzmOIktEWPO
YUpcsSGCOLx5Hy1XQmHq9pa3glBmJL78d6R5msfmBGjGc5fmetNVyN9O8FZzmH1k
1J8MPyiwofCk43dLmDKYNcTCG23xXnebVEcObm/4LVUnKOIS89uZIKmbVVG5Z3zR
o55O1aG+ajtRkMaYE1lOH/ZONuXmI44bPbWXRbYYghDbqSOCO7v9WEDKJKLcaVwb
3UICO0WqRPMex7E+45Yvjs9bww4PrhizunbisaG3HQvLsVgw5kuq+Eqov/zwTOyy
H7yXDRbUxZTOcYqvwZ+nDT1AlqpsLfUtiZZuQm9UnmmYDWlCg+mYJHdncHIYFpyr
4pa97OJHzw/QiOliONSoLCfwcESbsx45XPWgvLiqSZJlOIwWuQojhRiM79XAiyak
KXodwjrmVDtFcfa6fGu1U0Oz9QXoLLFCAVcQVrj8WVkaitiMI7ki2NlSOTdLaUh2
PVmY/hAz5ovuSbgaOVJ+NhstdIYOfohno3rFKtLws+xRb/eNrTscoDpiRk7YuuhU
jYU2ogymr3QDgBemMM2hrSVuoOPg3eonRAH55pWKSEz1zTykdwVvU/KGP7XuAiH8
cP+Pa6rp+vTWw/NY4YP9V5JatFWCWBr95gwq7u5xhFZV+TDWO6N+DwwlEa+hnFc2
2G9LRnyRrZW5PA/zwMcqrv6pn2P3JIu7MquJqVjSmxzG548DRLd468TmS4CJqbQb
jG6Uv7+6+rFnGbaa+SslchHzqklDMyGueCUzEiC0LKL7v1Rq/XRO3Xj4NyGgh+TH
nCH7kL40N9QJvNWrUnLdWHlTfVwT9BMK9dIHyEKMB84ubiIJKz/ftQ/zHf+t8iUO
a7sWQtKEaEheiL1IMlTKm1XcplALWO/UR/uuM9XenNEvE+LkGhm2DTOXEQfRx/Lu
gEnznDfd/9JeP0BTmQridFS1JrIEigHi205go9m8+Nx9t7yb1QBT/I1Is9ECAYz4
WQR3K4PY958FEhFr1TQIl+mUTrY7Xuteng/ojS5B+pFyq0Si8pkN/iJgJId6jQAe
BKlRMNWGh+EyMgaRLZMAH/9tKDY5SW93vUnuZR2+KfLqGIgp5HCxPZ8TxoMSdp+V
6wr8bpD9ThqQPDV3HxMBbMJ3yaKaiDA8WE1eHbUCLTa+bKdmjA7biSPHweMkFZTG
GfoH47r9xhfU5lMXl9FfKHLQLvSCpYwPOw1fvdXO6UqvCsHwOJPoIj4XrZoR8a1+
bJsLVsmAWVvyffYZBQNAushIUz01FRBcTbB6f8BtwaLfR4niH70Kmk9hmdfREXY7
moEcJRMbhxo4d3NnnEAhsnfhQIiFnj5gPZettUIpG4DGg7T4L2EfNMNzgddISRtB
J/U+M5gVmp9fv2KnGX6diQ4rXEp7Hy8+C0qQzviHlq3zr17iDcWAdjvZXYJInc5m
K6Bj53fLuwT49z11OzSDEsHApEO5titG79ucAZJsoqasgQhJcyZmR70Ss5nyO1yh
nut/ehrh34UclsPTU6yKUByEDKb9EDB8AJu/+HqN432JUA2HBcw+s9rOzygi0iHY
cEmX8fmghxpA/v3vM8tWO5kilFabbjtLY8IPsw+RoYUHYQJD3ChxkJaoqpUs3Bl7
AawHRG4bO8vi51kbs5qqvBjoyRCSrzCpWu7Fru3bD557kR1W7d/4QeAyjacRrg7Z
wBgZ+nNb5+CK4nFouQ6tOey+XnQagSe4qH7L1NNDPd4nyjyDku+ufV2LlHXdrfW7
tBdZ8fUzB1vK/upQdxuWG4A1pg9/HKQppPKYvCAHbEztauK9OQZNrJJQNjF8uE7i
Tpvws1JSV7kNRBVsvXixE6bMNezNU4KIqjrODltVTBnMuXHgsXNkXg1QLNQ8wXUo
7TmG734xTHFl27lFyQHLcE6/iVvJQHSia+kwuG7jNIXKYq3ltXcg40OyzGa5ehou
kIkywQrta6gZ4DytzXYrbrZyeZHakpuioBrvvusLQt2k+LzD1PcR8Xj6UDeL5cdf
4ztpa1j+kL6TtRPfiTapt87F1prtscJshIOqNW4LNvp8g9ssQb+Cw/5WpVgWj+Uv
EhpcHJwi5BPt1iO2AzCpAvqzeQiXbvFJUjRYjnTv2KXvs2td1YnQRNLkUlPjCGhf
faJ21I2AdiC9qjdqSBlJhEXD70q6/urr8NgPjr+WtRt9/V3OUWHCXCOCihPa343A
Oan3aLIGKxGa+5i1wcFkttbKbytGcClG/r+5ICVanDQEi8FniO54D4gZ9eie7Vg1
P5H0y9hrrQjsPm4w3wuTDJHybtpSFYaiVJ5WX5padAO63SFTTMROYGfQzOohRcxi
tqjgBF1AaFEWS19jaDfkxb4D1qqdvuknXquva9v/nEDdZ7TMwabV7jH0ZbrpqIX8
1HbeRyHHhbDeZMdLsFOPFaDumQ2NajKPA0wcnndIlWEmxFhN/9/0q6h7INOKvBtW
4DTSnjd2ergNy+r5RKtSbeotmudLlGma2Q85T7GUCW0rvjwSE6H++ObP2enwNrqe
ocNgjr6MfXms+40adkNeN8eUdmCfInQ3McdKsKQlfKMwJMnrhk0phhuyIbmPTl1M
OubPqlTcT77azAGA+mVFjlVfwX68Oz1cD5eOeW3qn1Lb6dV/Zv+wWWCJQkAiJ3j8
av7ujLQSln/4IieN8bYJjX+3NQBALmM85z2qGk5KBhAkrKvenxF8QuvYR8rbqrps
uFwJiFQ7K2Zgf4nqz4EevmQbshThiNuY1VEDLTX0q0BJLDrrl4etdQZXEyASG+tp
qGCzQro1EC7bzkkONOPbE3DuRnSDd7mHuPk+T4+ePWXlqgCBWxCpZ8o5Ep1fNY7x
ixrWY2CF/lj7po/AtM7ZkIhtbaUCZ5OPzqVop6B4oDqYhgbasgicjcTkhjA1TXc3
hsnJUptFK8V5y4V4QmWxcuQ5yEX2HEMq6QklpZ8O9p7qduFUGLhIGjsH5hVi0QMq
5+IAgK1rLTW7r/wWG8OAT8gIUo1r31lC9XZq7vo9GL1qYvqnUM4srMTVdTPusNo1
+4Piyue24Q8fd0BQRTk1sfNZLFBjGzi7ib9gc07/rve75X7jS1FICY9yn3INrbk8
hggW+8e30KV66NfxUVF8yayPGCHAfrweIBPPzm/8rW4EZUcKKKSElAD2UP0ov5YV
mNgOtDvDNOAcQRJmK/fAgKhzEsL1V24DOcjvRteq/EAiIc4Vn7uywjeSPIKiUnua
J1FIASlj3qqtjmvT4PY84W6jBhA134V3COJV0ZG0GcxiQaMdebhmBqEUDhnXN9BI
LF0gMrLQlOsrLHVADsIQPyKmd0pqSmhEnhDK1vgKnjwq194/y0fF/XMn2YW3psoh
GGFNnMILi8e79nIpwyxCQHIkHkIGw9wf67NtqsPTUePrnzEpXvf5b+hhnMcPXQCh
Ld1lYFpjH/JWLgtKc7PvoVdnvbtSz7TR9jyj0WdeL8W+/6Fa0cnShjH56oupneYP
N8LcpkCkNDIEecT25geS80urFQtKm3JhwsaNqWTJh/VZridSINHVjEM/BtHP/pIn
L1VvRexREhhKjjp9OtJ+2CfRAaQ7OwQQwDkcPdj6hfqPCc5FjDNU52VCfiqBq+xc
H9kHWqKmhJIuJ0PQP6827QGoWQwu7u4MCZO6QBWCR8Ay0c/ehv9m05vxxhe23y1Q
e/r672vC+k4zQT9keeUASXkWkwS7w/AbRf9cuO/PedlEDHs/Od4PGHQJxSp11Cmn
L3UlzXfJpr/jgS+spCzQ0E36Zl5GiGdaCrIxkJleHpRgNjPooBo2HrZN9mga1E2m
LsYmW2DHB3mGEds+GZMwTUS1TmaYYVEiwo8cymZua42iFkhpFbgrtEnwihPMd06d
D6TygrB27xHFOTsvC5jjs4A5pOJNAb8PLBMPijOqM6slCatE7406TwLSCuOjWgp1
zh3zgvkZdxpgOcODcj4aduCKj+bR6buwpQRf7uzxirSodj6rd/qiFLs2uiQoGlSo
3paRCq7iooyVmtaP8odyz8SsXGbkcdUj2IVkMGhKqUEVUnZ6d/IBzIJs/hlW/VPg
0DfmgeKn1Y/KoC2y5m4LSBqeqxFryzTWKpqsUctdN6A6E662zfLuDCU5K5DDJHGx
dhbz53bix73badMfAkus9eZNrqW/l8djqILgE6v5D57sqfXdyzfs8hDRPjQhL2Md
CvuZAHmrOUgaDboMHaklZdzEvQUkO4ZTtojB/GZGTx9X/g+OvaHHIGfWl063GvPS
GT2SzIrSE2WoccwbMzxKewRSnAPclSj9e1Ux6Rv8pch4mbjpb/HC44yoqsHt7RO3
rUy40ydnWBPspO8GsOWbiH7Ici2whikeRpkYf10hW3aX+03saRb1WtSJfWlNMkhR
VN8Kn+1M1cwJPBK+jFClhE9DSzlAFEji/xLGGPB91uCyfiVPfi9enKdUy9Bs7p4E
n6J6pN5StoM/TyOgZkonSoKvPvH35Rzos5hQSyB3ovrapo00pAWhf0FCHF55vd0B
6O1wYkSjzIQCdOYCKp/Y/aqg0V49rD6OAjvuu+rOfY6JU2rFHNIw1PO+fbUsP9h2
rGteDBJbVn3V+D1gQUhFaPqlCw55LbMSlauy2KHZkWRNerbkhtt2dtgwwg10gqzI
11fw0rXshJANFlHU5UgIJxVzSLjRzeYMlCCVpF7W5jAn2F2sgnFoFYdGWt28akve
G2Pj4ZVMdyZrH6UvJI6Qf5Cnb1YxkxQfoiw/x4J+f8SHv8M8qZIwbNuS2tzuaPZF
slm3pv7zEak4OzvQslUJDKrtTPvdraSmawNarJOEo8Ws+X1xNy1xcYLqWH/+iAWs
8iW8qL0s34KAzF/H99n+BLzgdbnuWp9yEkjjBeqBthcuGOoWb3B4VeJixh6KQHZP
jpQ7Ix+TI0i5kwj91lyZnQxyh/BRLvYSJ+db3Z1lQ3I/hKUhbov4w7DUSTNLb9SP
yB5tlfgMhtjx1w7NXSGjdQ4vVXGsmXs5u4X90BAzW6zegFVpFD7uQ4Ge09YvBMVV
Xvub1VsOUrFaztsnZtjKS+IAObi6oIZ/4cmVSMZ78ymlR/6HrFXgSlJvBGcMDJOT
lE1jD8daglku5DJ6nx8PYprFfaXivK9xwENx1VOCgfrlenFaUL5ZVJlyB9HiSSVd
s376SROxAaWcUpFIqi65zNixPOPqIlVLSBSo9ij0C+DIWzMLWYAVJbmOrPr7cymA
ULiZldoXwX948TSkaR8iOQUUy5//eE2vvmpygkgt0J2sOI3UJCYVRO3RNFKnWnaK
2Q4j3ngcKi/EzWosRPQSwMqDlfaRCVry5FVaiXesV6c7oQ4Lb7rRBANkDX2ZYWbF
s0sEtn4y0vx/h4NOumx6mxijfXW5DyHX6jR+t/jogvjwdfph3E1hcNgvgf5IZOLA
RgMO+IT3pBLhxBVNVMh+tn+hiREDWIIN674LdYmvH1L1VtclNle5e6cgVHnlwf7M
FKEc76Z85Y0PN5hh66fj36FM/NSrNgo8JsC1TRI9jtNNRLOTUifwowEoAkaQGZSI
UOT4xe3Hr9A0yFwTjvz9WQrtJbOHKr3R6xXHssFwFYF2GEo1HsxhTV8F3zaGSF4X
eyuxqkIm49epPoRixXTQTtgWUYlv9ja3uHkHu4u5YEflewsv/uGYvgUfPau5QVyG
+G3eQyS/vqhYiwdSx9QhdDpknm0CJNNom++9beitZRwyU/zgeE1ymHLimiyIWnMs
UdJGQwX1uV2UC68VlEJs4ZEOTGq+r9pRjX9ylPd/C8jM2oHLEpQ/mKNMUUxld69q
cRx8/91Z2Qu6DeChXtlPoxSA3+4RL850U1wX34h8P68jjHeM3c6fvOHtqB3PzNSz
5ODeCKO5AL/ufdB0j2XGPmNIcEqNf8qulyLirthGovCcHk0lXXivvmrKCCTeTXl1
GEdIa5cPNn5WMtZZ22P89gfsFMk/WpAd+iBEscnCO5iv3gcna2i6lsqJQXG+h0rl
2mTBRWFfnOZsLI3BFIpbpHewAAchdqLBz24qjxdrifSEHYu8HOhzuCHvrgnkRZpq
KftXN/Ydc6kGhpe0Xbr6PWZBHRkhq6TQuSSXIKQSu0feoqqPSjCR52WfAOkyoaPm
f/UswP1dwa/8UOCWq+cbVcyfzZefH9PaeH5XqgRiGvnlKK4qTlgg0Zb4WynF7S6P
Zx/xSwFU3C0PnP2P/rDDouiQDJG7Fy4JQL2mUG4/2wdBl7RbFdL9JdfsDBV9tdx3
VDFTWyzoaAAJnGan7OuMn1jV/lghSrKHQhZi5OIn6jZaFRjMxrpeQCmd+aA3mWu2
lfssQo+yWTTXXEztpj7T+fStVmwyUIVL5ymOQt7y0TT+qnC0j6FjD6PHpIsv5YgI
wJGpBJQINY0yt9KNhCymwijXIu24mUYw+tCOca3p1rp9irB3xk8d5LV5MW+m6Xu5
90UM5Bf9pekST4YAMRqK87OEc8TiFDRdDGz1LnXyWPZgSBgw1UBM1WI/c9IkeJMo
PN/xfNz9dl6n8dwe1+UvItsKBKgXBj+e+1D3A72BkqRpbK2epbZ0motPaGZyo3+j
EOQ/L7yTLtbFsxs5vBwOsmuWZ2l+Efg/SycWwFZULV5ycl4Bt+xP+E5qBKpvNUAP
z76D/fgUS2otBj3u/e+WH9RPXtZOOmYunJA7a5REcgrPONLQ+XNvaj7YC46/xKei
nJbecy3tP+y4cPIDVNtO5T9Uzf9cFYQH8prmgY2QT/PYDkFT6XTc1H4RxulPYmX5
exFv0tkBq1TYP98bz7zYr7+7rALOd62vVdg5x09OpU3QavAxhtIJBxB5xc9niWh8
mNqV+JIhKx4i1MJQFfzgpt+/G8dRuFMRXd7USjj+I+3TE5N+08GaiKcVSAR7XDkN
qOXK1bJ0ydlqFM2JlXguAQKHSNsPS50xIbBmMe/cIEy4BYxABGSuBmS0+MDjEJGF
ualNJgu3/7J60tgdBbqGy0Fm8OLTg5sFyVcJtwaRh7zaax8DFeppvRB0tEkwjBE6
ivpg/t0Rvp2eAzyBQED50XM+QFkejlq2xuPpIWR6hJFYvlesYWGCkeE0j/g7m/fq
fpmhwTINNgB/Wag5s6GpjDF8k3a9uEeA6H7clQ88X4M6gzTQURmTAQp8AMC8upMo
kVTnC1TJniWILo/QlqWUw6XLUTcOlf5xPh2oGBNepF4Xb24Ongvqu1FcDMgdrcEX
36v+4s1z83Rgs0lwBbAB1tyqjdzeMRTyYw37ew9K0oYTAcFNdKNq9tN4wYt6Tie+
I9M3TkCeinWK+p2VvISkeV3NsAhef9Lkd2/bISysbkwcqOsOwrrCPDy4fTgoq+lr
gVNlC+/IHPpYKhf4qa7LxmimY1WdUWNphczWDnNfPlgLoBVoGMmvnS+XHVkMpqD6
gtQn0VM64wh3x8SqnFuJDxyn2GXXjkcPL2L0EQ4DXSuFWyfwor7pWEOKNYO2pRcl
/Sy3Hqx/uWoWQPN/A9+HsJJoifxx+/IH9JxD0HEw4z5eAnIPm4AsWrFyZQRESDaf
aS77Eb0eqActafAOqiPchsnGBqeIU4wSOZVWDQDb3Hubxf6rbDDJsggaJIWxdTF/
3HRabVc71+0cgTB2f0DG1eds7H5gR3srScpvEBBLmu+CLWRkByg3HGDbtvMHeuP+
ZbbJOjzOL8QDVt3GxGmOyPkZzwefgqzwp3ygB9X8OpC6icPyKV/GVbj+cr/pkbAt
xgdqhjt8bYDpwIoFw3EvL1I1RE6AwdT0g9tXt2R6t+10VW6+W43tTnaWHe9K6YC+
Ybi6Y2iQWt7/XCcfTp2WOJmRZ5bkiGNsTjpHV1p0CWk6c50P4VUxOffIod+Roqpw
3vf53d3+spd2V6eSBzsVWJwNnqQOBDMOUNoIMAp2MG+UYXnHZb+rrcrwBDhNfa6f
sqkZ9udiQwRMl0ah4Glgf4TVxvNnbNBwVRP/8gkDZUskZMx7hkv5XVMHbXUefcEZ
SYSpzBH57dFfOLA7zOrWULftMndOYOjcNWoELw9fxmcJ1HCbcZMODdPX3RXYp5BI
nu0huu9K4EV90sNfMOKTx0aOBvznBzts1rQ+XW/0JZOd7iKr8mvtfp1OXbvxgIBA
Py746Pb++mSSyRBwN2wWRalmoy32fi9pOTdE04iwONuTQsDjkEuNcrm3KEtLQFkp
g4XujlFtzr2wuTMwEF0N5HaHsgnfNiajpDVeB5OU32arqNfn30BDLiiTAeGZDwfu
JblqRRIC8RRkHaZJlhEJLuiKl6m4Acj51R6XSfhD1RvOstaFTG+mUstKZUx1SCLd
ruqJHcCvWcfIC10Ri+RaHt3Zu9/J0uE0CY6hpYo/jxrXBNB7gOKowhmo/eJjwf5p
FIrDpkgSnukqy1Hj8iVYGek/+Ps4CUvEJ2JQwt2t57dWWaGyAlfTotRLZHkEIM2Z
bD+ttvBmLzzPB3PoJOBatwtIUisZwyDnblqkEOBFVkYI8mmkFzRRZzx2eudmRSUs
TEOiCixcdJxzYH+DxtGbDxxj+q9CWfIK+D9/1J6AR54HdgtLki5JA8nqmUTLNs/X
dYnDmldeXA1iKE2XkdVHQf5GXE+esTgQvF9f/3L2vrXof3k26prvk17SscPwDt/O
TPJhsPVCS2Ce4KIlLCPGFxBog89Skq/qzl3ZXy3zUFAikQYrnhpKhSq1AQGvl19p
F6R69MbfCIGUND3K5HFVLblKPESWvSbmf29/Vwc5OWIsfvrG4RL+WyG0RDpFQSG1
VpiZ6tJWt4/Op6Vf2l3G1WfxDODJS3ZdojiNhOf6VXMVqCqniZ2r20FaBmi2CtBt
1/NoMj+4OJquoRiwCAgWsALUFL16KDTweXAJdtCrE2Ms1r5fPmmQrPDTlDkYigFG
q3RijNWBKTLanKf5Khx/SX2ztPE8iyloVhKY5YzhDrQWbsqUon0L/avVvh1xPt2K
K6FFHTYruWaQiDyl82sYA+4rhG7hzWtvnJPaeSrLHzJdFodqAPnL/soAqDmepjLs
GTbW6KVrubO/x7so2yZ2WzFoj4HYs7co3HPE4Vhiihe5XCTzbasvH+OqzlpgYX4d
mrf/VMcofVrgmqE508Q6KISkLSOoJPicv9GxGTOv4kAzDPXyNAh0NdTkFphS3SMn
4M/v2GDCvI8B9dBzIF0DsSGsBonApO7ugbDhVISED9LOSV++17lkrs7FwCxFDzPn
/m8FuI3lmU/5UP043S0kcFsbEAjXdTtifO34hZ5gJliegkq8bLwbqRmQoKSK3hDh
IZKkzQ3Qz34F9bW3XG9jN7NUPiM5xXnUSjJEGx5ZV20BUg+rqyxksoRr1Oy3Vr5/
DuFhM8vFtFwSPHSjScrtTtWIv3rsZ77AKIRNaEPIAj6w02VgfRNBw81Q2tUTW670
O9rHbI5g6VRxnIfRwKUPUFWgbBE3xNX9zPIXByu2sBTNgI6yc5fO8+Lw2FsA0X5U
ZFoNJ9xhANGGMeD1lM3NqMLanHajkZxAXIQaW8Ys7JL5Z3A5JuBc+MwAnP0vQiSG
biVmwpnM8kquavHEIvu1MToTL+Pt4XTOtQGZHyY619DgpOsRFWZqMbbfQJWEaNaB
tnWt3PikZ+WAZnsvB7Q4KqLhkveqNhJ2dH/PZJ3/HQP6Twh4K2lOOVuyXAvqdEBs
mONVQwDHThyNWo/DCrziji/W7WoitwF9WimNM5hIYT6NEM9j+Eg5w5HYseS/Ty27
yydenhDD2vj1GdZKOdlAuYjAqBh+iwaJAuqxaKKoHEVsOdrTy6W3zqCFBPRZAHo0
gTxbvHkNsw/CVSloJPaB418xBP7QTtBOGT9ih+je6F6to3dNWH+zVLWjj5NgDA/H
e6/2ObPl7DcGcal0RkRekJnQwMogSHyDr8kUWLhnNRlRc2IlJ7fJ7lkgvq4th9wJ
6eOKuFLobiN/q7Tvxo4U3FDJgNOKmvRdtsRpk18xFOrxQBr7f81+BIW34qrDgtL8
iZnn/0Wt0j7NYXlYCRSEhqwYvl99wlqdP21mRMQooOTl6URoWsUO+eGKQ+s+5ulK
81MewHurnUloYZ6LD4GZf/q4litrAMi/Ckd219lTS09KPH9g/ig+2XR1OXrG46oS
eywDyY4miIxzxs1V0wHCKa22LAUPtNj0+A5VtuiOHtq2/do05gpTgDyk/6O6FEjo
JFq5Ujy7VbXy5IDSU6jTIk1QJbOyXGofADhWn5Cs7Ct/KHYiJdHaAXWl7rgZYGAi
dR90kPAT+VfMDtA7sAZPyy3e7/cKNYAezHWQS1NWclJ7toGfNV83pfUwuxmzjCHa
TJdm9O7YEl19omAgYL+xetgo03k9PuXc7JjizjfgX0BpfvsE6ZA+yreD8kZ08PUk
6BUiii+sgbaI3gbf3GvbL7oVkRMHR+AsUHK7cNO5cIVMjVpLEtnh1JL1mu5D2Q46
O6Ie+ocsnoE38GNG2EEN0BOxVK5eyg33K2sPbATZKzYf1jJG9iQQepiemWIFerwu
ce+46+J7RcmakGmhRuC5ijOfR5mqfQe+IHMN7QpAaVQZCfKrtE1HKhya3/Yeyxfy
sO/hKwRmAIIFQaIeiLomsuSj2ELWBurBbgzeUvmg/CNrFADs2UoUKY+hdMxKaXWg
mh64wBKpkYPTuxxbYnazQ1UA5Wo9dH+bH+ul01f9iEQQMNQioTp79JoN6XKYOZ1l
lDkrwQB70X3g6iO2Tb6oVrX02Z1ofxbP2Y0oBD0flzL+zTVDI2M0ZZC2pqr/Blyt
zgpQw3NryXdx0Iri0DcxVwIE0U/WW0gnwM6odnxYRkrpew42Ld0MijtZNvNoeThv
Go6HIZ10wsCXtPHSiFf32YoUqgYfnqGR/mT/bcdGYJcefZqI8X/5BZe39kwsxwPV
XpTIH+udGgMA/xQGZpNVN5AMCVoKILRX9y5WZtvMA5UG8vM+tkFF2kaluGxck09M
GRiYrRIHx33wVh/azT2Wxixo1nxrmI4qEnmnryzVY0xzirKeimhE4JGDPVsZC8gw
S2nMdwRWvXJSatXYmiuQ5LEX92pQWLJ8KP/3ZsE3jGI0EfWXxFjH5dJ96sQswFQR
teVXzSy/DrSadHP2aegoSGVkXeLlo6MRyEZ+qP0VxAO4VZ8wTruZToDWkYtjDJzQ
8yxFBJ60Kdc2J23HspUqxoQQY9txrXaCLskecX7Qzf+WqoJT4qN+kVKkruUgCHmv
kGrjuAlh2st8rbp/D2F+xyY0DcSRXK4ywmagsSpV0P7FPt8Vh3J5QRUahGP5ETQF
dhISusOcGeYvXH3CwiqHHDrgbTi8PwQC8CV82qHOG+086dinO9nZSbqbs9UOshbq
mA+1KeVagDkfEV6Z9tMI8e0f4KEa8jh9JlkvMF+6+Kzg1Fo1FjwB60QmoQPzONAR
BRyxJMLovPoj77crrKniYDWQ2EEBYpWBAI4KAY8OOSoXN/UeScOg3eZtKk+5uGY4
6QSjWQowRu98d/t29grYrauBShaO9oaCNTI9xRwLFuPOTjq3HNTEAnc/vBBFwAWt
bWJFcXMdL8DoAKaCqrGHzPJ9J1FVeRerxCg1qZi3EZ4mz7Q/5X+VXuOc4QsX7b5r
bWliGm/TYFrRuwImy3J0TjR2gNpngBvJsCbX4/KsPxMoZs8niTIKEGubBLAAXtT2
S4Qvi1dcW+3XOFCSf60TlMqtzt0rc7OZhg1iDTbrk8QAOZ5euwdzYerqI0AlXuf+
lPh1odO3Od9zkxiEUF8KpVKGNuUciLh6yqE+LuzyiD0kPkNDrDQ/QoTJ7rq9CBOx
BwcVncT677c87kkAamqhDciszXztiIPf/12d1Vqrqt6/Aj71tHuvQElDuWipyreQ
lptqVd3IdZ+bUlXi/AULabUqxtMT33RaMvMfJELMoPPSIKfKPoScpIrnJ4ULqlCu
Fw73RqU4DsQO+zBiGJZwj5QWyPqPXWz0YKjUd9AGhUqQ3tXiDYGRAw+YDwj6ZK/Z
rmiR+5AKu31U3fvw8A/riOh+GwIETUWMkSuHIVNa4jnZQlftX4w3NLgTA06HbpQk
N/bM0do0bkWV/JtSwOuOkUqZZVlk2M/KsU6NO4VT6V9c8FEZcI3khtubeSnGoyHM
tKj/+KlXMM9Hg5u9OEFr3EYTSylUmg4LhpOVr1ERrnSHoia7LifjIIzOXnLcwtwk
lsimVy6j5hdHQhP5U5J8UHlFYTHoMvQ7rVUhwLzMPFdSeeuTOh4MqXtq9hR2ihcT
cZqw7klppL7W+8Kn0JUdc03qDYdfutUZQSEQaMHSXdCKWtxHdlOd53ck86VX20Dd
dNIHbbL67KdSa0c88uMLRoR8NCtDyeJ3b75VcaXDTweN9H9n/zxBRhSGQKDg5UgB
Tde4WOlyRqoG76MYoDXmTOruSK3bmTJ7nEIVMjqqwlXmJj1syGRdB22Un/yGGxNv
i/LLzYaivqRv3BVY6AkQ8V2VXQA0v1qZTcXM0XY7NkjpaYBzA0NzlbB3EB7d9y5S
cIByf9n8oH4/HR1brmd6VLsXiKJei5OAMEVBp5bwFiu9H3o5xnGUViV2ROuMo4aC
Yazpphp59vu9RNPgjFckFyrQMD7fIPQ1JqRg2HmkXGqdbyOLZ2ziQ/07iDfWZNuf
16uEKtVdPfqxafXMgbqxwUDZCdEW5pqCICzcNbjrLZMORE5A/CsHr2vJvrY1fUUy
T5OkkRoyDuqICEi+mkUibbPCZWJnsn6IlZPMgrW+YxZYBxjngdO/EY1WfIeKza4i
4mUnWiBowGKvPLdfrgEwP+fRX6rwYlwWb2xguvjL+ztt4U9CPZUchMKCsT9epQMK
tVbIVsR36qbis8OqsTkaCc9tNdibBasTE1280MWoKQH8Fc3AA04/n8K3mIdiuwrT
OjvXbWNdtnjhR7/nN7v6xcK7d3kMZZrTVdaKlFFAloNtJNIkR0J3p0E97wXIkbOY
4V6SWGqCHk6Y56YevjdI1K60f1j43E6NQTBg5YPzNb2JZtJhDQFCLJPpZZYMY8yx
UscfVpER5NJVEHHNeq7QFAv3uPb+WO4CVYOuofiimceXwdnXce3/OqdY1hnD0qv5
YYfeWn7fv5m8BSn2A3P594+PrNXBcKRdJT4KMsVzG1gsQbqrmWox4VqGkuJJeHaz
a7RqwdptHFw32994V8rNR7rfvhKymmt7N+01EuU4BHCLwEQvIxxc5eSJLX+ZC0HB
fkOKh6coTYgjh5rm8YNvUfSvUx3+zrB+JvximJRZdHqOk0m4h23AeAIFdll3ztmO
gZ6XjpSTAZ/vVF79+3+ifmv1OZbv/aa7Ti37s1SY/EDONX6LUsd14ESVIGo/jMU1
/5lCkSi2csQ3kdoF5Z+6yjv6d0eaXbhzl4BC6/A+Vmh3KKDIQ5FdLhGev7GjGVvn
CixhYYadY6g2S/e+FEaWGA9XS67yQY0kTCsbVjXXDt1Pm+wfdKsmT7nrOiu9CSNM
tpfjzQBflcG3zRd2CVv9wAMv0lyP5pKVsf6am78L/qjQy0lEnWiFSllKyQuyEwYw
VLMEXEzg8MbL1BCW4sWJltRDnrQmg3j6Vm/VfcUeDmHxbqN83yGRl1twEBzVjjIr
78DzjX/glkcQB2+f+RTRLEIcVxGZmOQ1f1dCmcYNM4zy/Rhg2/AWB00D+OlfZi2N
suZ4A4YYkraiTK/GX+iHDaH4+jpbc7dpeJQ9AefO+embmmOglo5/KmL1oC1dl5Xt
ooJnCBmgt+TiGqLTRTXYmYMbmVlzV/Zhlzx1d95PRKT22uZU997Z1uhfJRDL61/a
79oqDbkQgMxLRyQlqPU86dj02x50hmiaulVTV5k/m+mHYdGNF6OJsKR+4s6PNCiA
v1H9w632zFNzHSebTwQqeYe53u72cfZPrnqaFmgIZEieK2krtAcfacYI39vNAte2
SXpdUD8pZGuIrRy/4Zz/iL647PQq1Ws9jvE5XeP38+//wTImKMd14ZttVF+3RNHW
tXj8VqWg4lknAn0RQudLHNqCpymg6v7lV8CiL3xWfH9MarcR/C69U4bJUkURN63K
nNR0TjKDg92wt/SwW1+wUJ3D5OGFrdaDeTWq/STbPoWLXF3cjF0HvqhzyFxdtR3n
PcFYiCM4T5GSlL7wh78vUKp0299gNSBhjYZbP/OR6QNmfkdtqGYrnPrZEyDTLBaQ
nR6w9iF2Ll25CvIC8w5cyfJNjf1BVrd606Lzi+hhESiEVTUevVh7NPGQa/Etq1U8
CYtYsxm3blRKBCBAL1EyZ5AweZp9a/ajcdyjzTNYcVFeVarP5XPkEljIlGyOvcwZ
GgYqb0H/DeAsrcjqHyvTY3pXAm0lVVUz+FJ6ntXRx/+yjHE41TT+i6hhFbPDeOGE
kUAU+UQFqthTLtIIKrX0x7IWZ4aI2na0U5zvGuzZjFqi7kXViowmhlsB0gKBhnSv
3TeEXd1NRK4n9y+xQ2rFMdf2VK9DwwbS/t2gmHd7vlui1xPBHXXfGGDUZ8+QgZLx
POVUs+tk0fEt727XLyCbUXkTHvk8jFldoNX4+Wzxvs6Uk38g/z/3NnYiz68y9/e/
rvYHAhohKYfId0xoGQmMH5raDBmHA2qtmM7SpZ1GSU54ukW6ma8PscDXcCy5WUIC
anNKhBepOwy5VT1Hq3c2DyOwXVFZphclZ24HtAHglgkyBrGUmQwzi0O8s0hXTHJt
8nCQTE6+ISfwRM1iUHUaGwxAmEW9mSzGL53CCE0nJ8ULsT2Bs4TWrX0IBkkEam0j
9pIXYBDtGrv2t+1YPC+v5f1vz1gi8EX6AmtEblobUksf+wujQ11Ps9Hn9xcdRDHv
jYKwzs4eHkaY/umIYfyGKbpCQB8vrNSe9hz91fhheCeezojeIUsJWamH2nU4DrUD
j9sjcv1zoRelCYnD+ZP9MRLddoODERJ9yfms7nV6z7hof5Fuzwf/Y6jmim3WLPzw
Q9WSxQ+b/7x27TvN90uzhbQ3BVY1j/793O6n62ZjyRqd5dOGYj46a2mjuDvaH3yC
I4sxfMds2yC+1s2kamvIAI/EiXwnEzulETLbHv9ECYYzLUoDZYAhxcQDnTx6cYZC
Ev20LOEInutSHrWF5BuqH54AcXbZuxvxlLihVzeIOQwztGrb6EgMIgNVBO8J+S+d
R9rUYmjd+vAEP/1wd8QQdMaRqxilUfGXDbiOh9dCqbxLwjkddFuBBlzlQyiOGbaK
ajCYm1DJ5haoTb/aj0axleF1RZ6xQjkS5Lx1IBUXvGU5u5EQrLdbFaqP4cVpFagU
dvKXUY725nQuyM37Xabm9mGeTUU1wUejCqjcgBw1Ne+Szhj/6XFN6Tsdbj7JkNvf
ekEfeRXUY7TAml9RdxEmW90ZPry6E7OEH5ocW6THqplgP8tbPmMj3EgaS52vlEv8
/JJOKJC0eqOjaBVoz9vEQkrDAahogVtialjC0GLRLBpUNT3/M7YPVZ11DuKxdWkH
Q9CiqBZDGfYNhHH2Qoue7aqwxbydSaEd8+6irqdvMshW1T1ybtt17IpJYo6mnIyO
ZCZ3S0jfynm71sJKpf4+aHnAl4ejNN25B7yCVsVYYRdO9Ir4C90anEoz2cf6G2Pw
FZ8Zwt0YCK0LU9X2jPLMxiR7BlWGI/1SKvfUGbhMpw9rsP1+Ba2V6qdSog3RByOR
WdSZwwfMeTry30MARb7QpK8QRgdQZVsjPnNJH7Hmn9a5hSMm2GJnQ0dWUHMpkS+N
lJvNbyvSkvgBRLHSn13YFaWyiwjU5GgKd0osp1S9wFMjH3pWINzkt21pgC+qv2TN
8KUaCkT4fTB3cWLaUhN7NFhSZbq7hdpTK4lQBZMCXucBkVKuprQg3GVtydjMxjrJ
r5TJJKbSxVDci8H+nkJ9IkZjNPX+MfmWur+rTOtNnpRPof1hnuxgk6HyaP0r/BiW
Wd/hih+g9uS0gm7IKnASbw13WWo+fAWOKfnZDM8zMXao46O4BnB42hZRg/WJor/O
fHE/tSIBguzczw906uuZQeppXEB/fnSABc9xVZGAg4RLJbxYeksOEGJz0hfZwk8z
xb+FI37G9jAtTQAA4M7cGSXPY0mjFwnfbCl2yx17voxweao0A7mNj+Fbvws9lCgF
LTFg6DB1m09/VEi3Z61VBQcEcE1RDgTM0494IaOF4Jn+sUZ0USYP/3LY0jRv+zWV
qZYZUn7QOgl88nInNiiTwPOW0LcpXOj/5jjrziS4uzs+ZdIqL22pEdWcnnPaYyQX
PzKbWkIthrYDzKvey8XrAV5PXGjzFzPaRb896/cYuqhqhqpjsM0CqiY18QjrRE/3
Rfd7pFHn9H4Kj7+Mk84vSaOxYNtTBbK0T5MeV3JYZNgsbQ/Y4Dogv0URSMJVqtM0
ZmXEwdkkM/1dk1wupgXvsR4aNS7j8gzogyg9Gt2YbPEgOJCJihjU7B+SP0lC8UbU
kkiH5SR1OhlWt4up5+ZJymaPnVP+zTolmLa6V+f4M3KORVLAjTmmk4JlHQ4LuZlw
pMeswYOtFpaGURJL0FSNt4sqLQ+S3gWuFmz5yPnwy128P8hcNj8DJ1fGfxPQCZ2e
Vdh6HFHqgr4jCsEl6vfSwlkQf3jPyHUEloB8ToixN63AH50ZcOiZhsc19k2q8xZX
ILruS0TJhw1ql+i212oCgmFiWhoMWkENu6HyP5UcZLSX3KTuWpzMTKR53e7LCY0W
YxnD1Fu57ARgrVRSeip3hqSfINGvg83k1rAkqL7IheP4ncpDAcv9EPDN7/fzUDAm
qmDGwnxT6PpuYxAfB2kelZihoXMgTfqrloT19E4vfy4VNmJrZfC/AnO3MRB2l1PR
pGzItARydE7pnu1hmZJxLgu3eyb30VmJzJwS7jd7QEnG3iwqSCGu9MU3MMU6KMIj
JXaxub/aLDtDaO/9nAEY7Onja9Lyl3Gi+Zqd08bFcQeLp1CfG26Hv/Xu7J7ECxz1
uQM50UaKxbMvk7Xc9/iOxqrI7nxpqdckUJp3Bz5i9ak2zBONKv5HfZz7H3tfzrRv
dOplsEQBV4QsZL+QgAxqP9IjcaIuv0/wGcTojAzR0olGrcScYRLHJapVN8rV8A1j
aiKA3aWMCtQTYCX2h1oAzLlONTmj3b0IZ0mv8KBk23tM5JGVcKO9z1uHyPVRi/nQ
HtdwW779Dn5BqIaFmH1QG90gSl1RyeN976VN8sirTXaulcUUkKSZOxc22tQKFfsf
CM+RoVmOToVw/WuOmXmRO6QnHlUoTNtt45uwTH7f/dJuBwL39pMTL3j75nDK1u8K
tYlX7xL3RC6HyrHKbT4eTutZLCYKq4Eg+UsmTo5IIzsB3m2U2SN6q6RZdhIMrifh
HT40sjQM1HerRJIbujhKIXYReTseDJ9VXo1RH2RQtnprU2GN6e6TZPRotz5rU/Wp
et5Kv1qFop292NOLXYASbFdqZHDksCTSMWGSb9A09Kn2vgD4n20NioTxN4PXK/aP
ZcWcE25DRL7jd+DFPmbg52nE7sdFSFsB9luxQgKsC2fDqTS1NVCwRUz3olFYSHqX
R0W0TYz0gEpxXAXLssdGzW+qjHBBB/aeAh07KbPZzCjkkal2EpOqcg0XjgiTm6Sm
E6Zvp6jF24sCCvocPErmaG5p8d+BHt2q+WpuRCnQqPPzNM97nmpvWVqvVWNkBRLo
uStq/fEfOEwEAoued+HHmAyEPdf9JEcDr/eH3Jcq7qq/nhG2VgTlZYS9ehzyKiEP
SnpO4KhWZ+2HyWc+/I3ud43ymilgpFUToXUyw4oXv4WBfhLhXUC7Ei8dLpxGXEpG
4NjBV01t7mwqiPU1bAbHkbrZKum6g5V2UNwxHGhbe2DPI0L+to4RK+HLb2jMofks
VHDj5ojt1G2ergWWfPHzHUSN1fHPW4ZJUnAqUbjg0eLlnt+7Mkh+wHV/6yKUiFMq
UhTy1NsrhJZAdEzA6WMuvZUP2U53QjWXlKSQjuU3cDl72kyTFvncjJkf3XfefwMf
1BtYlILZJvtSuRLidDml51UjEnGbiwjN309wDWN4ysdsahTHnfnd6MQ03gELjD/V
kUfsxcVThEnF6ze8IDtb+Dn5hvjVGg3yy0mGIqmG8efzIX73IEQ4p83AsT7EaFCc
ILCpFfuQlSD8Nvfx8YGqveRVtjGfA5dP/uD0tP20FiFLQYaRQKTQ1t0VJrR0bJMD
sJXW++YP8AtkSTwD/4PlcJD+4BLiG3Gr13gOhx45Ca30sxzGOIQlSxJ5/WZwIkeF
Jnxrn4RCoBkYOxvj2DJftVTHb6hmwix8IxcY9qETp7QaLu/DYA5uoZHdFiLCenKZ
FIi3Id/oQkabw3cPU3Ssr0O23MuXHBi/H8EqW7onyp/fcEjjEkH/3v2XYUFV2e+S
w8Vwj656ti5cg0bVw4CQq6uRLUlAJ6xfMaAr1Ot+qeyRdwAn3ZTz2OktAKP7VMQ4
bPFWeZLjjHoAnzGSboorLo/jXPr6Bsy2IEpXFe70P4roh74wQOcyLurf5ZzNGzFW
EGUoqWmwgsAFgNGJO3B35Qmj9iv8Hrq6O48QrXrwlSZ7/CeBi1UlSQQXEZ1UD3v9
JYmef5bLQqG/ExQa5CPzZ0vD+iNKwl5coRu4uC2R9Dv234lFUkYhaiu3E7+oY2W2
TVrOVxtiVDdxko3gjJsW/LqvtSRAA+45HPkUWK9evAoVihzBhVsGSY+nS1HsNOpn
tGcCnoQTbf2c87j2CmLg1tek/XDUm+NDLx+nLDGQtj8KKEWoumgqdUXhS+v7rieh
VNA88HB2WVpxzHeT4K2/X4BT0515qaqT5VAZ+BclI9+IWzE4vzhLgVcnlhcRnQFO
piaDckZw/gkWGVrwqDi0/7majLG3tTu/STse3XozQs6A+UbmoQnn3d2Ko326t+jr
g6doUjCaabWwzhd9JFtVK+neJHWVZzGES12Ftg0tvDFBYEflh6/49eYLiM7gjpVV
JUHFuh8BwWRW4eesMk3HkkNtt7VbZK/cn1BVSXIm5t4aAbY7jQ4iH/KT6bq9iMc1
Ma1LV4Yx+4247vc2PwXsICZwxiUJR8vbASYUxP/RR4ZwpmIkSLX5t5+4fB0eLg6p
AsEdMM/i9vlLpKH+qH7acgfWs221nsYoSATCVYJOtTRw4GsEdZlyuGMLJSGx6tHH
I6j6GLWBOaczaZCBNvQ1UgqnZmmkLc4DuDQsdmtnfRDGQaTdvZwS5luYmxEhanlT
saXBlLswmOjYu4f7c5qUxtcl6727r1CXVNc7r8Xne9T8fLvCdpbJMfUnHtm5hT4w
O5CseCJhcPQJleoMPIV8D+d5FPCZK7OMoIyBd6Dqaq7CNChFH9855jFVPLOJnuWG
un2xKaPYFtYEjaBk6zpoxfGFUvdeSoz6gF/bEDWFfbl9EADKZwhwsQ1EKPsSD4ns
lUTz23jswIDKPuTwwVacwj2XXCe7nBdBIMFO29qBTijni2xCxqRpsSAzpHoikXg2
Af6nmbW3bEedhIxG06oOf8cG2EZvAoXysirnH3z5r5pL7bFPf2cjvrsEMkCt95rY
O3rSasK7uXL1K7H3D7v2kjgt1F0peV8KefIkX6WdIlg8Lm69UmDUXcJeJJDPnBy5
JFrtnvjCxGYh2w5PhUqMo4e9DvvUTqwJls8qhAF7kFKO87ObM7zojCaVejylyp4Q
VRLn4g0VeWgowFS2mCJFed5IdaJkGxuIN4xOtiGBosXvf+wz8VtDk6cxuAbhPmgm
la70E0iUbtH8qIrZqvz/GCxx7gEjIKtY57UNr0Ne/R2peaOdNpPYjjqDTM4W1EV1
GjchZOaC3SaHDoy7eced13sjUWUz4fzCl1EpHMudYTadh8Dbwg5hVGSuBAe8aStO
CKc42tF0V7mN0dHw+ijbPCigf/okISiTjqpkL2HdytIpRfqb0uK4eoQjqpeDJLue
4vVCkMOwp6O7c2LM3MvxD1Urv0XiASEO45OvY01inFctdUHEBmEi7OnzjjhFKKGe
5R4zGSvTbb9f7oywaIlSddZwbxwVlnfud214Gq47EcqqGDwbMCaZPm6VPqem4qh4
ecUN9dBkpXuHzOi820xp9bSwSuF+WRxvlyIGYFvgdxyY1bf5WJKql4GnSYpYUNcd
ty8722zqXpyd+i2a4l9HPE7y4W7nuDwVo+PMJ+F+sG2S/S2xfze6aTvjZOUBDHkA
DeO7FKTit0Yvx9pGCQ1SKj5jICPtg4UIHVmbMBi/wg9xw4xBCN9LvTE6dl0ZqarB
UeUaBoa8hUE2ZiU1fLbakboE/mz0mr9+zJihEui0I1Ou8vniH3qmHqSKkDUhW6xM
K+9O2Jf5twnC75lXm7Llw0YlfC803WrubYuM4H5eQMfrnntR/mwX2Gc7FPAHAt7a
djkHh4lICVp+lYD6oe6Mcc5d5aBC1CBNAx8PQNCI8vglCfdrqWc6sL1xqONYqwt0
o3amXC2LiUABCAZ/fPgjbrLvwX/RisXd+CFCdfg3c2CiIL84wEt2lGn79celGMw3
k4ukhcxiX+nWQhzw1jafgp+tzKqrGtE4/dS1R9/uksF8dVIqDwX2Bt9yzD/cRj5b
BAUjmJx/nOztUWcsIasAeOIBpL9Di1MVmVX1WVlY/wXMCFZ9ka43GzBMLZDKGLqf
XYVNtE+iS0oJQDNqvz3gq7FJMqY3l0eNJ9hlu96PD32PqObeN+06bDHVqzeNfC02
+UjnDhs7o83nGg99hG7CuI0oUqHH2wW+I3/vCRuR3zCCTBaGIW41KojfyHPuPPAV
Z5KKCpgoE09zd+/M6Ti0kPu3SfQQI2YuuGVvReBaiqowFhaMnYSG/uXXFGJYlS9r
Af+F4/yJ6XHqndVrGcm8/wIpIV8VSGsX1oL59kqjUa6jsaHqOZsMmih1bs4ITU9S
lduwekFtrQ/kipIrbnVCXXPZLMbJYrJ27jVSqQ032+KDnOAJLFYzLs+urXIPsbr+
olGhIev9abNf5qhEiyIJpxAGojadOdaARJELAAl4IzuT9R3tDAe8P8X+6XkuQ4tk
jAcCVLYkYqqdq2bJNyne77qzZ7II8o/4cEDrUB+tUm/QPN3aOuARfZLsVni6YDnM
nvHWoPvj/FgTaCTHq59EiqFuOr6SxlMgNx8mnnaG4K48ftdUZ2W5l66sA9N1NF9F
FGMVsb7OFgi+NWJFSQ0Ss5l1+sHMPQNI99Mu3SvpT3ixILYT0kKNp9OpNhRrSgLB
MD5dB4Qs6TNKB6MUIg+FLiCNe2Adaw0ugJMZpghYd9g2NrOGeMYYLXsTdVFyFSmE
tUBSJZylX0hX3yg9cnEj2gbLb3lk4CGbO6aOjqVDzbbx6SBRaEpOFGsuoXmwjUe2
2CzXK/rTn6iSjQK+a4l0jmqVjSL88PX28g1hiYNf3zXFaCOcQAmpB8RY2caGtVLz
eO1DvDIA/NV1GRA6vFLkPU2QgiaRCDHLtQXqQy5Mwa1GIIkoqf2FRRIRbbZLjAST
Cy/FxESDsQ4KtYS2ZB9Cwk5RGw3Z+OuCHdl8asWG+KN78OrsiO+9iTFQ0sObhCzm
EGsdRPi70I48L3NOEAxNrXFV9keSMOj3YCEGCbR0WlL2oy4OmKu6HtXd5MKUXVBZ
lWmpUj+YOOyLqr6FRZdlFazehvz1IJq+VWh0ULZDC+6pkS+/91sZlJLKua9RYXB8
9fWD39Dre//dD7PQrHvgdvWBZaaHKj/iyjyPOG3H9uHdwURrHx1uO1CIoiQR3eYI
mnSeZGyaf8gJ+lOhyooyBvCV+kzl5+ksxGi6AVeE7f+oNiu1OwZaB3VqBKQA05Bv
HN7GZ6qJba6VrJLng9P3oGTSHpe+fQY89Q1ktkOcO5AebE4GN/MwwfgJpkEr0tG5
WQXqNteyEz/DZLklv+3yw+wCT4t4EKxZYdSsEaoi0C4DhEqZS6l3rVNLRLPiVI4y
FtAruoMvYWuA5ZMXyXFCczqWG28NJA/4aZNAgxzWT88Fcdals2092xTtthcnAB/F
dDd5zGbHG1PjWdaT9LYrbMQ2nZTjBrnqcd5ReoPM1j9RDKaqHVXFhhMeY8RYacgj
m/9ulfx2lwQrfBkkKdem3uUh+KXNatxXLxzx4Nxcdq3j1B+/JQThAgPpg7rlOJI2
qaP7g5q8bWluy/MirPw1G02mBwipC/fs9S/6teD9yP/hnuM6GVQWQY0F+GaiX9QL
4iEXFcSZqR4d/A3cVZam9/YPzFP7Vxw5g0nNOUYecGaQ7rYBZDAlsxZ7OoBsQL/I
7iRgBAxwAPuW2jpX8Sk43rTYdGM6ZpDAxx0p0Vj0jjzxvyZQhQ7MByykvOj0eMJk
QGTOQB4VUM5x++Jnp385nBwAzpvUvZT5we68K9J02KqwlowLsRJ1NrMoBoSAdwLc
UTxO8IO0u47e4Q9eJFGnMzVHv7DVeOxIvt0I1b7xXdEHQk44lhp8ojTEvdxD9vKc
985Y/mLYEJLiuB7l8RaEWnsI0qtdN/3VQE6vcBxiT7OltqMtZ+0KZu6SNV87zHs5
BrO6rhngQJ5cfIaoLebvvwqfGyD7JDgY5aAel88vdg6IvPrlVW+SdrrxRy7ol9T/
zluGMVuTaooASivQlj9tqt4g+4W1zbLedOufDxhTrd9LdRKJMnyNGmQxqo5SFpM/
TbFkpKvGIgLeslIbnEzplknSJBosH1JzdBjEDnYsNQVr6WXAuO7OyWsrSNzmCoGB
LQhqYMPhmMUpqH5Zgypu5IVqIT4kc8fQ9PaQalTPSeH3agfgGl3NTRtfJeuvgJ6Q
B+vEgD7x/j5TcBHddbmymTP7Fa9B/zjCzr2o2Iaow+GS1M4vGQpOOlZ6dk7gOfgm
DUu2xZwN3vtK5TInRE9BvMx05jv8/AkLAUk9l0E9iainK11w/1E1viQc6JXw3fo8
pGLXRUAfkppy2Wxbfees1WBQ5kuTBpIb10gbX3MXXTotvEdP2wgKc03weutChPI/
umeo58HSRzCMV1leDhjI9FXH54c3SdXDyy6GKlFvFB2YGoE9KjrVsEl5+N9NdKUc
J9wxdGlMvdUaUH35oSc4WIv30QCXMijW3GNFmP3tv8UGY1k/0erLE0+cDeHaZ/VG
oG6RCm2RwiBB9UVPlPmcS0Q56D2flhFsrl3OHSv7Jfs4PyFglCFHm8PnJ/Qhq77I
6QcbnmEsoc23otC7y8zrQwGb6sjdm+4EY8QSLljA39ijJ/AjZJlxEetsUauncFzm
uKNHzvQd2N6vwq0XdFCAKwxqnP2C0qxadBlr2Xn8uS0N3frB9DcwJkgWtAoxfL2Q
JjZamYOd5SIixPscf0gi8tyCytW3eIbDK9trQMKbDTHPfXanfsHnyUn0cwlXAk4y
iklznrvObaAQ1GVIbvEQk4ACQbqfZVY6gX3Mu7jNRxKx59OxulWFRT82OIsonDmy
EvdemIL5BaXRJDw0eXMFzOFz8r07IRuxQtQva1VZLp8pqC4xOp6yCb8j9pS9fasA
0uY4gaZxjfjf4DBSKUIw+4eohOanEyzpZGUlmpB6/Kd7JCc9kVHYK5AmuLhceuDf
Ogvmuo1/dYaiGKvtVwECGZ7M3xASyMEMwxs9/746LCWqFA2huKj4C/f0pup9e6vM
BBPzen1T2q2BQj1Jf9gRb8Bkdem0IRrRzhRR3l7jPweUgYuvJTag0YZHO1xvnL+u
AFfzDdkC0BqX2YV561+DmigRT3vBD5iHWYj2tyNfIOFQttTUK0mflB1C5IuHcmF3
E4lNe+bv74jOLEAqTe9HgaAPCq2XzhypypPQOQEIYMuAGWeFbboaNBwnNxA4Ye5j
+WDX1zau43yXQK6bJbSnIix/pNw5WfqwxDMS2ccvrFFpuKrKZmjZsEjwt9s+FlDt
ODeRpfZo/OSqMhPiT0jXwoeKeLKldmOLEtIh4zddyIbuavcDLkywu0N9XynFmpKY
hgi3OlQQKnO3f9KmjoXO26rBzb9FoPPN63d93HRatD77R+8o7kjIBnj2w0hiVFqG
vcDHtkdz3E3guww+Rv/zuv9ygF0ZXY/tofRyYNj0VpLOOX8AXhaB1/JKKpPzWU9q
PwhnTLlfxt35IFt17NHCRYo9ujzHR4sSQDNAeDm/Z1lIuv6HrlKRPATljcpBD6Vr
kj+iQA0hoa7GUeBjtQb5buRSSXsbQ9tyoyDX5LpzArMJwk+oZOVjhtEPHEtSxG/F
kNE580BlXyKhVybwlTV13723bdmbfNgKO7EaJ8gjxyq6RDY08QongbIxdsMOkf0/
DqG7+y8/Tswm/95ZYn/9f6ijWR32UqBuHD9pVA1avFp12z6Mj5W1J+w+Ttjdyv0s
7GqhM0+QIcQGKieG+SjxTQv0ADKp5VhPp5CEwM/SAJ8KXmG2KYdkjQxzmxYNCV6X
zJ9xQTxH6rarZFR5mRJarZCKZpklk3TyvQ3HUErIbgCldxFuGkAqYnwvx0Ii0tj4
55oxXEIhGe6W9GfbWXkyqzvefCOv96kLB0zpL9r8nftWhSApgLDm/ZsBap/LaPAW
+6Z8ugq1mKW+lFNWa3aJ4il1gJrS1KenWnO68/VbbrLwfT2QLiWAhy0zNEk3M2zl
7ZAPyDaKKdpDJIMs6wnSon+nooL/DHO207f7RlJxsTEB6ELjwqPK/DMJJZHsoTJl
wDkfBCbbhwcxVsKPKZjwYig2tvLcNN4uYB1Ks17apJNg2Vs280lAMpCF4J83QDCO
uBVyop+bBQVLu2qz1i1h2IoOpjXMAqDM4tWpBwAnkqmDwx59PeQwq2cZvyLa25nd
hZANAngEQW9Aq+jVZXuHaWJxh23sT9e8r2myelfMMPmPSBTC6c8wswSfD2d8b1vV
QxHwL9WErNVy4lQL8fVafBPrVJ45fP8SWNfa6hgk32gVk3JLFX7S0FkT34B1MMdk
NEOONn23z6rKSu3QfJDc9RWlQZniPztCCLSGYgF+ziiMboeb2z/X7kWHBraIW4VX
ismu0ye68z6eboP+/MfWCrYVkPbknWgJE9mG3gyFCLSmJgyOrB1vllG/c0773zKt
cxO6RKcH3VAWn8aZ4Vu5izqAlIKgM4ZJ8TwQrMi0qC/uM3+ioKNG6O4mXfDXTKqo
gq6N/X0NKCDG6fWUSAmxHNcs8/oGyDMdo1rteWWHkK3gnygsDbbZ7GQ5F3mjincx
85vv1K8ib/PDXGAW7288KHQkXVsTIOd3DvzaEFaLzIM/T2Sn8wlBHCkAQbfN2l5F
OpBy3fr6l+gGKfv/3l0mLDN3O0bsY3mJw73GVcncs6vuTfKXzvHhf9fsapQtqgEL
5d6IHPFf7oDyhlO6iHvlMarPtIpLwqTmWxQ/spnebgNGLnqN0RMaqQkAPle+r/ic
Q/v+r3Amp4g85lRZWHSVodrgk9gRwgT9xaa4tOmafs2M3eR1PvXvknMWn1qG2ihe
Fg93PQpdpatiD69Skrn/ekj0xfh8S0DNnjFqs0PhdDiKq4QVXEoUNo3HFRnhRY6l
y08sMKeIXStu5hSiYFp6EtsGw9le91IueFMVythpXgpO4RnvD87XbsgVmISRZOpf
QEM+pXjYhmvbwXNwZ9+jiYKhFFI2xD3P6Z2boGv8/v5UJ5avCUsrWTeBdwU7CVOK
SWwrBnfvUHcsGANpzgHydtG19TypdiPCNyuptOY3qDDxpgF3d48Wa8WyqTFKzFBK
nWMj8PDuior2Eg+FCkrGqDSmebs34CjwaHce75UA4O1MSrG4lXQAmC8sAT5jTzxk
djBfZZvpPPYsTTGfZVyHXDVtNYEOLc74lblWQ5tbEZpNceA3qdqyixsu8fFJdLxI
UdgDR/yyyHfWfpS1Lu6END02Aj/2I3QNm3IwCBL/2+R2H06j6bcNiysWcIYhJVN1
v+nHX49VnlIWRnRzynEKoh+crwhnI2G2WgOfUQi4M0L+js3EYZJYPx2gz5an3jt3
UB7ZI/cHfV5PLagDAY9oLRh7YfpBwsns/MRHEq4DVJz5A3LD7AJ5zKlbQNkujkKJ
bx2QL1xyq4/Pxj6oVzBn3XMcdMhhqJc/53/x9ST3H/34VCxej2xcR4aWdmVgStM+
3xr9DUux5/lHriWKoQ2gbkjJSnqGR6oJJ1f2addM6/CfURv+Qt0MVzkDFw7jt8aP
zoxEMBZBdC2UI/X8tyw/ZwOTeg19GY6MzHEydlKIPxyE7q6PgYdkAJ+MKA1NIUZG
R+w+zXmEF4/PUfITRG7pL8Cf0Xa4NJygVh4PTodM3mAXZ6RHlfYpoOUSDXoWmYIT
3iK1v4vA4SvC7wTG7XFnz0+Nve7VnxCNTU74f32xS7hsXDqienUM6L8J6yQW6PTo
0n3O/hwmMAsCUuhAhRfgqEYUv6ijkoclM2sMXPSLaRH1VogTaeH1fhGY0mVsQ/O9
wUeBAuGYlyfCGB458w8bYc/RTXI8b5cmNjK1BafJycSyNar/Uv0fAN/dmZw9XhvA
4jgk+ucGN6UgR0O9Z/+6PGbsn2U8DIjv755PmjAN7UrrCNVh+xzF8Djc91wpS2IP
hMvMQ0nefK/1I97rbhx4Lx8tKSFcI/NUO+1OopUCZjv/SW9Qvcx84uBmy7y8WXiP
8Way/IEYGGcGQ3/5GulVxnkuZFQRsogrOdo4TENzlXaVH+AxURnaW+STzJAxFMhN
Rm5UzcNZnmwabXbDsW0HKX5R5bPiNOW0jdU+M220/PduGGFUaRDh+Raib2fcmCxo
kuOta1GbTeJ/HnM2hIiBeY4gJWttngWJDyjl3dY3ams8PstwdYzwyyXAnsrp3nlF
3gCyh0bDQEwb3Xlu+977PVB0jD06PuXToLgti5axeIlbcYyKxTYMmzBknPF9fHGZ
gpkNiFzY02XaRM0nIBX4iEcIRRghXWEGgzROOxrOyhnonnVLwMxuL8+4T/J8u/v0
faMFDU0PYj33hJBX6NRVT9/X097TJaETZgtImcad9Gn4Qwb+h5/UMDLdo0fDT/aw
KIVKksXyINo9Tuv1+U+OZQRYeSyHVu3oKVLGcnDf2u8u2QQXcPzBW2AeoE49LHag
bk30oHDVHWOWyUF2Dp3T57jQW0S4fV3XTP7uVNzxQQGfjd1DbwmQI93lRCXLHoDl
qlcMSPXoOpLcTNO2aUJcudCkshF/HPBBRsVPDLiLNIGILcboyonrd07Si3udqrS2
Kohrh/So4oyM0uVXWgQTW9WGlN6TG/LcFNn/xhRurIkAm+1fz5bSIKXPVzpeZRXP
UwKdgdzN1sZSrbrC8sL15Gy1TIqRiXLrP+e8Ipb1Ag34mtEGgkLZLmTnzWTlX4wz
ymy4421164fnHBK5Nca9c5RLm+mRUmFru7GEmMrb9snt8JlgXOQevdODNnTqt482
RIZkU0wT3TFjOw+OYCbOEkeNGogQMknrcroAoJAJZ77pzEC0OW3M8Bkpi02oaYlH
eJAN8YfyfGLkJEf7FLgMu0uqh6HV8PVoMrIEvFhQvNLBVcHId1x1e1vRcUsHfstR
0xyZ43nK3+NthpKkHWMRBWPhEh6MKSWrzEmzCDTrNKD/4861oH6C9HI5hxBd5V6+
UxD5IdNG9+YuU6Zb+jQfbZ4f/OJJqty6z5RfAleAtSEQ3d4Yx5REOFVCzStsGxeY
94g7hPq7Ve1rpIGWv+44aJ9YZK96CDHvr8c6yJui6zN+/wzHQvKxYVI4hMhB5OF4
uxs7PoXGbUVFuidHw3eTm0M1XLW/1ikKLqvGlWloP3ZSY2Xh5n+Lhexzm6gq3VJj
8W8W8/TorW1yPsnRhEDa7HeCMp1qM7hXa3A4njFBM665hKuJicx6wO855HhAZCTA
3WgqP5bve8l5Tix2cskb25cOIhDpNTqx0Q8vyWyGAdHbyMweav20MSnySgvokhm7
Af6l4/FajfVUnifgGt9bvpDy68mp7b2mWku1WCv/mEDJ0pxrUWtKNWoBw8xDk5la
ZRmMPVbt5rWrvxBcmXqXoWvqLrsV9tqN1ocjKdGuRepX0BfE93lHc7Ucrr9kDXf8
Da5VhxINugqk7iXHNu4Mwo4yeiDRzCyaU8ml9+LtrZlEogONbK5dNTkAMHk/x8l7
79vglsSmA9DLb0S/5ix0Hn1gNvDoB7wQgG71uvTyApuv5gJHTCC9uxkTB5Fu/uB/
IC63+uyakcGVq615QHlhP+iZOGVq5TFRdIt6AEgSA2cjq8GUmAwwLOJSoriwIAEX
XXY5URg87H4eEVMLdxuyoCfiCQrgU98Lv+v25I0i9H6E8xAYVBtCKnTinUlRUxz0
VgC89ur2ygYJUEMY+QtLxdvCBU8x/cbXogwzShNi9CU5echiLtg3YkCnvmbW9g/f
6zDiSQgvg+JsOh04jAVAqe1UQQNS4j5Xxkpe6mFWYGSGiFofAZ6jSjSLDWWEbFhA
gPw5ZpbDPrCf4pQh3OoQ21Jrq7fYI4uo5gebXohpbzuwV6fwEO0Cp9Tcit85RiLx
z6PDjd+h3PRgRePTGa/CkLlk3Mi67/mNS4PUYo3TNYeUJZQQ19FRbo0Pm3tBa5x4
AR++/1sWOeIUcTdnxLyV8k6eWA7BWGzlw86ahnro2qOOlY7OE0Ya1p2dO0s23C0o
8qNdkQGKFfBQzLLGP+iefKzGv4eQLmY2a53n5CQsmhKkrseRrzyNYZpNb3RTQKNo
kDxaXiqyZbcQnqlA1/jLcGGpVt5+AMi6+IdRMHGainkUdBnTMuSCVtQwDh9NGnT+
m+uO25qNgIrTchIJIpSnNsF4qpVlCCLTUiuRCN6TNFzmPphRcAIpmqO/qx+Mzq2K
kaA9o40EEiVsFCYMSBGCVnVocUJgByijdfShZ3YcHvs9F6Ybba2vMN10pGxyearE
15gBCNxkr3gffIc0nVz89xku3LNSXJoEpMlMG4KmE560LJjk2E/M524mZgUoYRYp
7lvsSc3eDz5GTJQSX50Gyd/HDvU4PfgNnXBnbtT8TvGYOEWAUFgGDBnUaWIreryI
lLiUbWCi+QnaCbWTiDipZ9oScapmr8iIpZBtH1SMzbA5zsjy+RVlTd5UyNhVr7t0
igGT7zLoVnQ69XX+LeXVyZrBb8NRjjoqPMDz6Jb9lyQkZFFbXRB5iOak3QNhwIob
q67+T3F7DzfwD0dYAPsQzKOE3CPC50vcIvWz47yhEFmnJ798jHNavYZZnjL/qz0g
Uy1JhW0B3pdXz2fTusFBs4H2rtLsrC2svRxqXnFFVX7BJ7M03TwTQny93gl6zKlF
splkPv9Ott3/BeDk5/8lmsPM9Zw7GUmslsKvahtj0bRNorHY7hYflZ3PtLPk66M/
NBRtIEIvzItZpfCAiGbRfWtO9+Z6MvgC1nr+Q+QeSAD/4lZG4fgKMCQKLrjdj1Ka
L4bbToe/fueCEGaqbI3kREy0/06F61VlM6kXxc442HqYMDjNrt/M1pzFztWsoQ9d
U05oo290YPa31b7XOHV508eFFgbJ+qDpGpC9iwxf5nhqBvx9pblFBVClcKoi5Zrc
qW6cP/VNVIS6ZPIi2xOJTwkP0HWQ7EiQiJspaHn6EbH990fViOCkV4Adse7Ge4dN
pO27Itp+scP8JD2/tBdldx2dDy9gqV3Ux+BtsyziiRBr4X1XBlFFK6Tt7MnEgxjs
FWH0AZDZaTKn2fnSjbQ7XQohcwEN40Ut6tWp0ga6vReHkZl5j1VU6P9Dzfj+ovSt
uvVd2yK6PpDtkwypxg7KkoIdNGf7t4Yv05tvTll0uOI2ba7TG7RVyAXpS86fg5RJ
1yN4mXo/OIUBGvAXWJhrwsCFdBidXGKQhzBFqH3f7RAng968pKvribP2t5w2SRsq
I3xjzmEdYlg/5VUb/5CzC/ncrAXK0ASeO9jtE/LE3mHbcV42L1GGij796MQi8cLZ
veTaKR1cUUSEL38nSr+8GBDDa9pmGe++lINSWFtqaxqcqik+G+2dFTEEw0vFLCk5
4E6EUvavA5WBODLFX8wfjMCY0lmq0XYGLvVH5EMA+kmh0UaGIX88mDhIglJwYAtL
naVG2lbZb0BF+xHqqwupyDVqJJOZoVhw05wAOASRI2pL38eVKBP4g7ig0BqQApdg
HtHGm3YNJTMPEkc5mdIVEa2kvb2XnUI8l/+GxfrZgewpAg2PVqg+mRpchsQzy9cL
9fVdGYYk6fh5rv4q2velPQfbOISkPP9Hz/iTawb2rip9HL7S4Z+FGUDGV84hP0PS
ueQSE0ELqrXd9cD7FAXbdU/hi/aQyeZnPl9rbId/QZ2539SutIIBxX8mpJa0IDHh
MwsOo8PFN4OXZ29GEHL8mtvtWq7GceS3EdTQAq0ApKk8AMUiCctGSV7z+eKu2160
16UBxLFcCSNqCqx+I2aLdltHUgI6zMMGiup8LYvNoiMzwt5dc9dwlZFzoSpJOs7C
BP9lIh81NP/8UzpQsxoqrCqSyvtf6N9jwQazdi3blGMhk5gMvgzCICdM9o3HEyjr
NIXdWeg11C7e64+lL/mFSjaU6buX4Y/hATLhAP94t+qR1Z65oHerlPWP8qZ0k3/o
Sx2+uhm5bRFfzrNXnR7/BUA/2YtsDUL1dFoPjOHBl7M/OjagPaKHA2DM8qILgr53
IqDoWJ/weVG2faXNytyK4QR2P/wNz08uMFx+AEmkmdln1dMhJ6rgxEZ3rmY1x4oB
fnz3xYZN1+hQQ9TDGsbXI/SZavcKHGvnKUcdfrjGltAffDI/pTb/+lFhYk2WDWKd
R764QGf5XE3zTJJuX9xeiyJd6FrQwJknNJ6z+JABTq2r0XA3TQGW1CWeqlyJx5wV
JPI1XoeuCW4SXd4TvAwJnuUNKWyh3ywXEtlRw11cAsgYrP/ksbf+TxHTvDd2hHF6
PJ/syWyCwq8Na0q87V7x/9oG2MO7uqq1h3qYEKqVCpDS7gpFY+zzbWLQJOvZVaN0
wMAraFyp2fI179jzOnsASN5+xlYmwxXsZ04OA2Q7v+qQX10T7pj3EWc6WVguXkPf
QV0wF2biBTEVYm47lVuGQl3kB+n2JeHOo53mlSu32mMWzj0+iwVm/EJSaU6TNBeH
rGQDymRzpreotrTfLXB+i9VolU8Gkv5f/jLkQ9WNfb7z3nTqdVuJ4yQLQdVHu76l
TMx0wwHgl6k6wdfdc4/CvNedGu/I9GJlCif4SNR3/Q6QStG6vuK+YLXZOweZp9mH
Qf3LZSfZk+zJCkr1bViCDLxqXaYR/3VGhjc7FPIxN7FToQX5W1vq3S5J3b2Jlv6L
AV8vhJ/3J+NmUirPtN8E9X8km7F0M9v9/t8C5q0nwI9al7zEKGIGIj5wU+1JkOaq
ipzUtwbfaHoiqZXdQhvDKtaE80ZQl5hQ9+GnAWsof4+i5xjzzTrrs1pmdhDrNrzq
RlYijQrY5Ud5fQlUKUdTyfbvTExZE1AKylCBOfeWz/9IV4bTuA+UhuurNy+A7W2i
z5UUT2HGQ3adTe+WZs9+SHJCmckNLg4ROL1Jwtdvie5nidQxnWMkNEieD+FTeYR2
9uQrH0NNY0eG3doF8TGzUYGs33XikM+pNB/Ca6T/k393vLXMCqEwVk+k9bVRwwXf
dDc1Wmcvws0HXrr0CWtpjDr7FtH/r//uivOp5FqmUwMx27rN1rCLcqOtEr9msXqx
ivUnSAk9bc8AGazSolLSu49cR639Zg8G0SdeD6dP0X4sXcGZLYPYVhQrclXYcvaI
Qahq1Sk9PWczextEYkcq/JZ4dY1JqvcTZcxHAbbFfOlFYxoSHgncMtD425Nh227U
S1ePKkpjkIpKpBqnVB15quuLvtXJca5fWfWA2lieTCF1VZ/SL03oDr2pmexuDQip
Rmt94PoTDNZKIml3UmJJEPRrPVp99TJ9zUSuUxTW+u94jBuVAEXWdjgsYs/DbIr3
tEky4x3oiZnbSffG1w0YvtDUw0KBAUqrGQOQ+L14i9GLPyyuAM1iSrMajINxXBq1
L6uHrY2cbw1eOoChs87rQR/3ubesR47kKLJfvfmDe02E5sQwxgkHF8PtX1WzJMJg
riOHagpEst3ADYgqAqhfKpCy6w+yWvG669hkz81F/kdqTd8yqe0YEdIyw8OLEIHZ
u7sZaMy88B2b0LZJ+XM6At4kgQhhZaHkAVDPshFOPbAccZjzpD6+KCVqr2Zu89nr
kiOAbY1Hd0Wb7NP+OBFeJrtkkRrd3xAm3HFyY2g4Fcsi6dbM+n4XMPBbjGOJoHuo
Bi4IpUKuqKxD4mysUJlqe8JYjWKA44rggGEVYiAo8hOnBMIfi6fYh4mP92nUXBGw
dtxnjcmKhUi6tbVi5Pu8TcNS2XCRmGU0Blwcuik72kHhu+6rqktyQj/80kdP2brL
wq190oGlZhrvklJvEwjth4i5asB0zUxm0rwenYVK/rEdJvG/lv8F8zJ7Zq3XCzAY
BtkqAL0lXfzbiWR0TcYxmww+1DHvP30U/iYG+aP7fX02mwzk41kggLDfI5joYl66
mKyUgfe5bI5BJVv50duHr3Rle3hbWjQqVY/UfC1rNaGPVy7QhEUpvQROqKRT1881
BXQAliKFgggX13HqtUYw+hrQ5B5zSyP7+5mEuZU0psTS5JL/27Q0NnWeJCOOJsPI
NXdHhnCtfPQ+hKEh4cJM8Zk1qcffVjF9ytPNBU+8CfSyKf0qSr5AQE4R+Nu/nKb8
MzhhTtgBce3k20xFEoODAQeGj/+D/piay9Y6b8qAkkgHjdDg8iE4h1LZvEo9AUUQ
M6xHXeZyfri4CHDNXZTU7pBddeauofx+5kxZZc1kVWmnIkI4/rUIw6Ivfbj9wb22
1j9iQybKj0SZbg/AlIQUqLaDJLTgzSmhKywa3CJiHAATZnqFYIYRcfZQCcmz83jO
r3tEz/ZvVL2sWkqBS3FV0bXZqNisIXi10Ndi3XKwmus782cBjZqbbVgrYqg0f9+P
/+brsatQirNFvY22G+mA0aw2yThXSEIZraW3wHKd4gjcDLPSPCUiT7jhFErh6IYq
56x+P/m7mYlDcqpLUPdBIjmV33cOc0bEkkccile7Bn8ZhjMZtNNm3/DQGpNsfVTX
f4cNffQStNF8H5J62bqWMF6+PujhcHs1oWX5HzNXflK1ntAzv1bVg9AchQSAvH3/
hUfzscjpkwRQnIEPN7o3Lj2VavRc5kZFK9yP77gT0L8dqSwLpinRNR9Qsjeh0jqC
jhaBONHesdLHBN3HINTzmTtHdn7je/7V61in24mzqUN5LRxGEKXZjAcamVPbYnCS
Amv8X2lW5JqNTyuUtDScYpTCgXw5dUE7iVzCHNhwMUyXrYXBtwqJsW52d3AZlbNf
1aGwKoC6e184mNB8YmKJOpzI+kaLQx4MN+JLbsosd+1/yA55X+4uIrzO/obPCICX
B9ZcMLGeOyzPIfd6UEJ7rL8C5vxsRGUnq0G9XcqvQIIZFo2TaL9YF9Agq0uBhPOc
ZnLFosUV0TSIjQZR1ycp8GEyxdUBj7xuYjRPV6b79msTk44M5thwI4YBA+jUjNNo
DfmsSj2TL+29BKQtOiybEpnypeH+HZjIVq2Te/3q6jPUwhYP3qVRroopvYdV/TGl
kQWV9AcGM6L/nsvcQegJXy/UyB0AgZZIl73uScoT/AdfEyaaVREwhzDjtFRoMhra
TQFdeWykCUQu1vqgIVZllpKtkW0cpHvJRTqdI+/JkyQlQ2+KzHfSkYrzi/Ls6BXH
5toPpPX9pDMjrMkBvmx2OHyunaO/TogaOUsQBpqQHGn+lKu1QYq95aFMWA0H5oqa
jxS1oMuXMi0VBoYtAXvlBBDWYLtN5rOc+1vG8jWgA9ttndPX0XCPNcH095O2aFFG
0LbXutOrfDTAiPPlFCtgBEw/ynkYE9ljxR54/SXij0axxT6W13J0wVwq0tgd+raF
i5Gb+2vL1p4F/YGd2nLNXd9Epzy9wsdSXL76oGh1Ih/63Ju9h9GBryqmg5sYEmn+
ak1yV62FWOY4kJrK19+UeVuvJa6wFHKffbWQyxkDOylFiYs5SJ9eVigX8C1/a03F
2Wd7R6zZrY4RDBjYWw/gVUMSb2bbkjzboSYkglCAwg3mQXbi9fG6QhOsM6TzbLTR
FMNGFjtTpRyBDt8Ewg6gGxb+HHBBwYjU8CnVvuUgL30RlWvQd1x3cr2SU0yTI2zH
pSDzdBptiwGxpAPtHXYNYGydVA2cdpxsuQ9paO/40+tmtCpPpEOQbCAgNXGEgNMU
bpdiybkCpCPzfiqTys1pJ2cxuBkPGcPS+7aL99A0Sxv7tnORUE1HDICVIzm6bFQX
YapplRMoO0jiYBs6DnoLmqzk2yloIcoKBQa16AQGDT7YkfWi5Cpc8ThKmbCfnPc5
pPI1UIFTRsE1Ge2iIR+nOtQA445dlOg8wISftwvtdnTrOb2EweM+SfbnO1Er4lEx
BPVwiZo182gVwcBOVj14MvCuw8e0AVjrNGRFvtk/cvTDbRkN3gXdBKaZAXi1HaRD
4uvbYqwABqkSBRwxxQaX6MtbDO4/saiArK/NHwzCWhXX0XxgimG51qdBbreZ79Ls
88AFpFHjjJKZrSO9BxTqWuRkykxTtyXiua4cIJDAkxszeK2tYKGj3xLnc9o0lS2Y
/l8N8McqEQEol1GsnwY74G3hjMqoFfSPURPYglDDKUN/0hXjbOL9Y+lEaHbTGkMh
T3Lx6cSBM8eo88pp79ZGHU4TNaxwCyCthX/5VkvXnnnOsKpe/FiIS43YAu4g6Rzx
Xqgy2NJ445AIihcYgiTiQaPasbFCinqMymdYZ453EtaVH3DSUTHE2FMwfYe0hkaE
d4ZjGWVrTgFyn2UBPDeHae3/yvSnBYlgM/AOVVrODZmlrz8QVQVQM/H581t5qbTL
1YwC/MEupqW2RYe6S44sg9K0vqu6mC/vQWHBKDYCpXB+vLCvdi6Avr5Q4YDkmxtt
YBqjUTGj191XDx69HvCnuHTDtWwrNeUB5tE5yKZj93gPhFE5GLjKSg5/bUhFdsd6
BWkFd8CezctxrtB4w758y7WJWVmX7D/Eo52Ngufr6mWHEjBsl+s/fDD8sIZ4f3Lw
FET/6sKoMRP5ptrGkftn2fpQuvG9fmqO8lE27a82X+BZ2yKSN4pDyfstSz7MQEL1
be6Zl0mk7H9t0pTp7sGfB32XyByRKSOowzflIt4dsfLGft4nelFodmYHPkIm4ZmS
WcJAudlVhc2Zjj/ujSOeNZ/09b/Qa9sEQtQ9tMz5LsX08eGxV8XP2mXYvFhQ4Nfz
evGexyzWNRXT9EL6KxYGpfdxncLmZD4omfnb1+TCENqT6TzZNAT+PjJWgOWDFQsY
BgtKqwO4lUYiHIMKbgAgNEkRIhagaRmRl9Jorz+FsEZzWnOm7yEPBVMt8yE40s3X
Qu+p4owMEKneiZuqla17wnI302QUQcacMIlAFFl6i/5dyZt7l5qG0P7lI+wy3TCN
ZDBnu6leITMgjvJ7jQhby07pcc/555TyL2zRNFnHpUyqdat1WWPTFhrL7xlIS7C7
Tl1q5Yvg6PV8KFignomYr27oJNjeEQm5GaXmO24xGZuyveUDa7k8tflTbwHPVrio
NE99p3smB29SZH5LSXfqXvAZ1V8a5k7dVQJpN59XZfOQVyhx6Km02XNjLzWlaFIj
QCGrVpSvfH84sKukojr7dUrtz6gSPnPfcfbTx7joV1PNMjJBdeX/4SruxD+Tx0+7
R+2oEpWn8rDt2Q23SEJbOVjtiEUw0GIiVD3VyenPYyJssDgYyYHexb2/aHgb9y/F
Hd61NUfZ0oIbkRoMqzb5XrFQ0k4xFKmpt6qqvzq3dwupENe4aP9Ee0iBvLfT6yIM
liiS249JpJ6G1U3R8lAOpBcPyhACAmRGbLbHLe25BjtCvHei2sD+bDo21ubN6f/9
zPCTUmo+atJn7XLfnPla+RZ/r/ztSRfJZlfjXqs9vCKaGYFx2RkDvuzt5mtiYIQ3
v5tUqPdu/uU+Z79jCqzRY/h0qFbrvkn56y1NGfABwe4XkELy7oS0CD+4Gs4yk2Ru
pdjRGKVxQFFUjCkVkatkxnxjjKr/ohLVKTA1BmoxKO9NQx1TbC3admW+9Rr9kQEj
d4BZwl2c/CgcFplUEiXOkrwolCqooxjVa0JH1bDd3oSy8PAAMs4XXxeMMHF/TZnM
ATXX+UK1b+NU/WS5T70XMovKt7Iurw1z3dkkVebmv0pDtpGxTpwBTiC5IoVvl4OV
gvIhj9ln8W3QG/Nnq0QLKZPXGT4uW7um9ghLcPMJnU9m3mblU7LHex238cIdFGy7
hdbI7touLXTrSa+tvWPnJ65LM03XYUfxTFZ2x8pY+tmrl1gy+bRCmh8/alH+AyeB
2HcryFaL9OKjuw5Mh4YIddKoHEeLBLh7dJ8Z5oBEdcp6JMC/ksA6gsSu2RZYv5IJ
AJKQMr+cYVIqiyiIFRNMs6QrvwjrYh8y6K4pGLCMSWMY/puw9qNHwox3Y15Aomqq
4JOW8/7BmTB5VdJPWMM6dJVbisMogi8yASHrc9X2AuC06nA7tgtaWeJysHmgPnyE
qByIkqaLogd9GRzAhIG0vrotGQBnF6Ts0DGMXXzPNCn0z9YEOYj+G0bmzjWbsgqi
FFJu9nHkZokMIjiaUbpgrL+8eHjaDmrIJLe4ENsxamRokXZHY6VL7jryGZgYRMHU
5hiPeaDc9SpO2rVxKvW+A1g1ykPmF99I/1pzRYFBp7D3sFtarth+1UwDjD2EKhNt
6Xng57412in2I29D/dOlj9mVPXhy68lchcFWHmGZWpXnlrZkGbkaPIhs34WErnBl
prDN1cmXqt88b43lah1H35JFxFzO2rIHdY2DPUmpfoQwOfs06nIOFK6gpTS9Gorq
11MnhZUiRbnvjpZPcbuCAtZU3GccpzE+3KXqZOIskU2BiA2n6WdL9zg0M4/QDS+l
Yei784IOg9rPctrFhr34DdACtBO6jTtuQydVGe1bPXaGZaE2PQxpJ8THBGuMDgGg
HhZkCVhIasUoETJbKnfhgIahxQ9skhjX1Snsa+7GF1gSaz521H3tNq5lefQrOXuh
JVXyuXHrax0N1v7AR6ue/O0KPw9JhCN3DOQkijTRp7NGtkd/PJxfkTGehdHWAKw1
k4UlSz2BZsPFBcbpAcdUuALCOsSHt8ftlYfkzWG9/pXbzD1DgNN2nI0JeFKkMWs5
BTqIQXYWoYSSGUfatV9ZoOhazucKkX4tBZYD3fgayBY22H+NCQ5DnF2V/cyilpEH
LkFOwaxT3SXvN9Uwsqbm/3anYTRUYFK+Rb7i8js5V8PZ3wpEmI/pL9Zm6xuTq5SY
SMqKdumz0kWTc1N5bIzSxn//CyNYXAZEHAdzlXey7m/0SmrFIzlK6JS9Kc0L1Upf
F4NluvgsxXCxCaNwmLIFKMHJPB24zEUaoIQmM7/wYnv6R8BcJ4/urrmxSLsEAEKT
s2eTcXTrQO2XPlC5k7L0LkjrLC/aYmhhNfcEB6wLJObU8LInyVplUtaaRpy+mJEl
/vMFPB6Ln9KsMquXGhUbsjvpnYfpH0dAkUAr4Aoyk1QAo+ZZsKKORb6DlzNtdEWk
Q9ZyPop3yaFoSVz0Rh/ZZNt1ePS+wCxVN3OFBf1km6KnsEV35EwgiAk2GBGXJV0H
K3ZHeoh4N2FMpdmcaM6AvLKxN9/fkWxYJ/AwZ2aVa0HBuNsWqrjV9S/uR1wPT7l7
5n6ghvafTIJGR+KpEg/D6lV923G89PKxTSH5YH1+Ye8yhmuzf7j4nyHi0CYbHpxh
DQZ5vJ803/BQi4CL6leejVkSPrTzEEEh4FdnWBr7DyX180Ao9kCYRjFZ9U0xXmYQ
F9gopjgwqKCbErgbZNYSDqs3uIpT/8Ch1hETFN8FJXeKw5EylpbG43h372wfDiyy
casGCy3YRLOFbq2npmxRxWchgRcOGoRoG+4gEq5B2aK3YFJ8OYFmdn9jLB2pPXvR
4yXj94o4ZUbkcKeW9/uOVy98okgfTsICDp0nQIbIesqrFUytLJK7j9p5yJhsZeOz
8nob6nRd6pZGwVtk84I7Rl3N6eS8HvNKkoendRKJYSZ66r7QNn7lVmI5yvrsWdIW
lRl0ewaJB1c2chYEpO1PnsiQ7//CYqX9jBYjMTMmFNBg3TlCwkL3HC76L+ptnB3W
sfV4Nt3sdeQPEI+tgsdsxTz2li+NknvYnN/GDU4wHOtk5g6IpXum5zNSMJwKcJXY
WHXaeW+/xhfBIFsCq/n8MTAO6imOiW5lgBZlhPauQcQ4fkbbHPBohlut7dF2Y6gZ
Ci7xsbjiA5ILR9JbEPmocu8JCzUROvjfc9+Zyzgl18z6byBkOEfLzCg8qUcZWkVj
pN3ZLylCBw3I04uwt3NBfn+7/eNPodY+URE4OSShjXtWsD2Oqa2Pf0P87hA/4Csc
8koZAptCbzvV1C2eADJCC0HrzFseFPY2BG/S6tUVc+cCOsNwX9fLanEuj2iz7HEp
UZf5IodHN8V97W+7/fDxyQWIwsJe1+JqJWPY2eq+bzK4pYo00wrcGzhDmExo3wNi
JK5/jKUJSWx+VeRo61PtBVI5WQkg+cx8mIWyZUCrPeWX98RqFrTzLCtEf/k6BTIE
g2HqreLPTyfP8gbty6r5A5GfuUD2j4NudiVaQ/9YZGevWMLSOOY95tpI/QAs1wG6
6BnFeWLqNCAY8KVmQmMzGekPNyi7tLALM8XJQguel76tBEvEz0NR7uu2LtMm4whT
ydB62EK2iPD2D0T+2V4DOe5tqvqE6zp3vSVb1J/LTXtDCFvgo6fbRMqBnkpUE3Bi
ARtzgU7qSb3bv/LPQ5R/DIios//IenqgS/5wNf5xRq3D07Ax+C47uhVBwxbugDbm
C+OtaC35qmeBPIthD2EoYEacNbfuVI2YG0UxntPg6zF7D+3dBU2ZB2AqYhdrnkiF
LUGVTUTKQQP8TpJqswl2iL4U4qhdfa1Ma0LLN7d4SDWtCicGXK51WS9H/IO1g5lP
0mQwgi6NlrPx/yuWjk6XW6syiBjEDgzoZvxp4gT/0QqQDrxvi6y27bKbW4Ot7Vqs
DmTEPOgbq/p57i90IZFspaNJ1EMlDwiHLXvTUrojliyUiyjUPT6Is8rM4tU0sQ1A
N38mATA/DaKntlJ7sVL2nK7MvKqILQlMIsDm5Jg9gxxtrqR23afRzE6mU5Lf5gN3
iEdScPFYxiOQNl+YfsELOjTOwcQR4b/Y/dgw/MMuFrhzfjvb7WXZ9FPFJibiUJz/
uGQq/hllrXbm7Ndr+TaKBSXMt3Evg4yAjLnJA+gPdmV02VnWULXIaq1ziW+TneeH
yFKI3EfukxHo6rCBfVAD4HwrJREJ87jrWOUu8p+6lrc/V70L/OUN2kuxhV4hVEAZ
oL9pobwzOu8SaPdbLQDLxFxb9TbVrgcOBC5quJiWKs8rwDIAFJjDzqNh6b+Y+q4r
xRHRNwiPYg1HhjbW16sfohvFZIgwdlniDz3RH3dkNKSArlqpQudEPoqppe4e31Rw
w5pzgPzvx6iZo+z1TtfHJdeTr9Mis3UTNkx/r53hB2iOmbhleucMHqb3DG7MdE1O
+AoDQkFs+8uwKtmiSE0P15GVD3GinjQqLyWxPjo1DMycxXNtmnMKGuacEyWTiOfF
xMKC9sxVSp3RoqTNB8bOLrUmx7XZFTJgN5vi7sQxtLT1ZKQFYTWoQIbeJ2hXlU2W
Vlvpm9Y6gwJeq5T/rMsmYg0FlQJ1S/IFzV5rOWSEusJ4iUK3Rv5PyyFlCnlyFP4q
SAXB/a/6icvM1oelMSUqznrXAtaggat325StAAX4QkTk/t1ZDsxw+5IhIHMxbXOl
N2O3rnBIx2ynxB0zYFjvarC8C41ZLcz8f63uLd5J+evdSNE7yf/hYVp4sAUtaaxN
rXwRQETLDiolwaFibTyYdS7NNYtTwzEd6aJq2eCVCzze0QVoiMWTn3WQ4miygvKe
YfgM1USp4+zCY2ACk4fAGrp5texhFDpz7OTMM6gSCJM3CJGHj+0J3QPShBge02Pq
PlHHi0ftMAWStIu2hv8BZE71A72AV+H/5x3gIV76zEHRE5XX6KHgWE9GjGwgbyal
dIkRntyFKPR25IolrrehxAQ+k7R5LVI69HmWrzqL0F0Sz4XcyDEd738HuFqv2ELU
r8b8KYvYv2GanmP8SdIm0laxgbi+iCfkyMujcy14CII0ZqpWwGoPafCh7gewQFdT
6joSzjM35ypjzafBNAapvTccP7UZMMKM1AFubHWs7J/e7avJqBG5AZBmyVQt/+6y
u2s/qprNKpx23riVtVirZg6xyUP6Gq1l+ZiRQidQ8RYRhDYdzrRrDvadmFiNMPkE
0G1qLBmp2xPn0Qjw7Cxgh4o7fMalmVZV4Vrf64NT0EA3A0hn50TW5z7e0es1P/Bu
4qvKYptswMQ3W2HKvRJ/7YDPoOa2PJT8ZJRqoheONc2B63eGGvKpq7v/MeiKUrAV
n97SbT1JohMClYLFjAApRKluFdvlDZsFZpCGPvb2QABmezEYXlBXEAJfOMU6Rd9Q
SJXqvUmm4fm0fI9EWt+DyKttNnN2R7zbbAKVXMgTpgViC+W+8X3C20d3hKr3KPoy
9I36IqRkDTExYLBsmzykps4tjAR7KicJyHHQjXwSjNps+h6lMBt5PXixGrZqWdS4
arqKMjld/mrZmTzQZO/k/9z08IuNGa3vVCSah3X4wm3+X7SjjyBCK2nkAPNstYml
enrzs6xVq2X+D4G5khEzZ4TDzdcJ9z9gmKSXoE6HN3yf7iVc1pPlgSrQZ2OK+sW6
LKJdfL0rPeNa69r4ezesBCQmYEClAop2pugo5PyXl2DN+OXTXzlBE741b8cISdJ/
JYhYyUnjtpPjMN/486mi3gmhPuWDS/DtfjH5GoOo3eG6oa4N0EoaNl+zuMwbFzR+
LqizfiWZFcL+A0Jijs3j9KoFOGj6RNfXw3fgOMyCUH+Wh+g7QEHg72gv0fYZqb1V
P3WqulxndQ8aKRLM0OLYlzvX2hUTcl/0yHrW1MGFU6zA+2q+5u8uGjEzt61ppFou
Yd/55qn4schKlK+bRNZrUaFVdMlUTpklGcTKCnAqiQAp/U3XMQzbDQ8O0nPQ3sGh
YHHNAcLcMYcMmjZs8HP7oMlCs4jeFQxHnwxl4ioTGOD8nWazuh5Je1zhCnYnJfbM
T3DsoyZFw8M2UZeB/l/x9V4C4Ev4qWARkw7H1VleCEkEgq/VqDABpJxWR/SVWhoD
MaVfQ+2DNuCBVUQ637aI06lsgcx4vQf42QhU1xmLsyTmMFxHXiO3M3d8RWATQgKZ
sk59YQf1UTFEfVAJOJhMaA11+itqW0ObImL0lkbx2JlQGPqYoARnDniszm/jlPhO
OhfMqmzdWNh8sfYqRO9HKUNYNP532OASWAY8Vtgc/Y8/INRKhpUCcT/lekNbNXg+
S8oVkc1QFtQ0AhcoZ49epBCB6N1PtEzuxV1Lz7eyYHicNfzKs9tc/ZiXCC7Bh6h6
u3H3MmXm3CbERHbgvVCQhTFQoO8lGlR21FwVegUOQ7Gcd1pBiQ1BEAvLtYd0J/kv
HlV1W5FGh+s/m0ofuC7BBaN298jLI2LRvQ6PYP5HQQS/wdcK8YzCcGAa+0mVg9Fa
oLJaQ1cwhPJGEA8jOAGObWN/Icge2TRXYMTdJdb5Tmj0C0ZZmcFSjJS7rE1h3BDm
m6JpuXWuhBG0W+lPZCr2Bad7iPq+OxfS+6S0/7It68w2w5d7+4qyjAYblEZfahkL
X7q3CVuu5hOEfT0pP6lFRdAoR/QTnTAE6Y0KGJ659Hs+kUgnQbfi1mMdFGcTwk0o
G0jZ2nKWQvLzwOLoPCRbETc3l6SFxevD/qaMYK7Yj+F6xQYVlY3VbeyojNl10DHA
8X8EAWzKVMnVpVIlM7dzSDIamS48emTmjxkWRYXW6pORUSOeH2/YXAF3ZgmXXWKm
jZRUxryN7M7mQYru1xPpsdQpCEZ6BSZ33wcDV0DrXPn+lp+NuZv2Hf74w3JY8UL0
RDEAYpsZ8dwLObE1nVQbnUyoGVYOIr2JsjxPMqmqFg+aiSpIWYop5dd5m05ciEjR
gSNYXDFwrX7ODOjsIJWy0GqWiThHYM7iJFM1b8+tXCOuXcqvhiJNnaGssgB4sX9a
LjGS+CYYwXNV8jXhwrm7UhR6vEON42crO+UkakMj+Y4q5auEU+El3Nj67eDfpAxL
q2HlHf4fZpL2lSeCY9CK3I1qiFVFRaoJ+iUkHrG9tqPb/wtu30GB7Bv+2px0OhdU
3Lylul5wkBU/VHCgvYcjp2LsfngWSRSK8hcYtnP9fYY3FZTt5RfSKQ1eWCaO+pkf
pCoAe3IVJe7L0xrnCywa2pStzwZa39RbOYlSVeAHU4ktibKy1V+NVEntPE4dHGGm
YEQ21atwJd8VYwaxWz1gNp7CNKDO+1iJo/aIsUILnlFUXbaZSa4NbJl8spOp8Ho9
oUtSNArtqRv8eHtjwqoZ3xK7Thz52Zr4iSIH2wPNa0PWFEwQgnf1UwbasW1jCySl
k0/NzFvvTksVSTHC91gRj78QUQFtHoeyV8WVpB7Uirz9CbfuMABZt156HH02bldc
ZuKPbRYzc77tPbUGLjk8otZOyNDKM1ezAW0QOGqccmxQIDI3KudRTceALT7RGu0J
bAwdAuTg2yV+mPyfERKGvyG+vf1lSk+E/O2rPCWWRubpxcq9huuAn39RgchII9gT
1gr9iWj2FqqYv7Ic23Ec8lSxClOnycimSNrNQUxknOvGObV3TR1Ou6l++BDeC5XZ
neaMXs5O4T6FCM0o051qLwUjq7t6aY6y50ljJBv1T56VclVH7k3aasaXNqQOBPLH
5sUpJd3laSnzs0AOFiWgUZP2rVQHG+8KITbtSN/ey0IOMaraQOu+BBDBFZ3btDCt
ChUNMJy5Obt5wN/acGg+C/CTM8mazKUSMCmuXciYiiCDVqcVOj9o8PqeWCwk4TUw
PKlOVHjhte/qcZ38TTpGGpg7yYkcE1DFk7EMl3eNM8TEOukWIpXj+dJMwPVtoHHX
5nwwVhUCFZyfNginWS6QtaR+qjjaVJuGpYxb9TkhQPyRhRUiWx5ZWxdLp0eIdqdj
i0Ly0TkkVM2UkLqTwwH9XiNBgwJ2zIwO+XbnAVLdQDmEzTLSmZYkVzYgeqzzONl8
hnFdTuXCo7BK3TFEcygx3PWwMdKAbqwLf3gHFTaFtYBE81i0pNyqieS1j/1EpXuG
HW7V7GxvpgdIjJv5TyiAiyfjXfIXGIbGNGHSQSDJ5ZsQWlAANFvYa1Bsi4aGvVfJ
xcEBwHDIUXzzmT0oTpgwFVDJ0v8Z5sXx8PNaK11bgWDTCuO/PIUmbkdCKBl0oQTM
9AJnf1pU6WRtaK0SCjRQkbIo2X7GkFHwOlXgEZGtxg1j85yr5qQfioZj/6lb4Av1
AomQn78a9lzJ0XozQcGjWTsrnmLE+VyKHnT6JG6AWhnqOpsv90xH7qSRUYWICvUO
3itbZRQAXOmmBgyfHdon+90yYk7tepzrQ2Nj3IY8n1awBWe4aKlR6C0MswfeIZjr
xDrYBxOEqesKMNlDKHtBJ3MlHAmiiO2h8XJt0Q0ICYkTEPWeb9mI/MJAJ1AEjDVc
YKz+gc0dy1+hfd2GKOBCS3j9aKAVj4pWNYaaBzPmIqx1GhXyRFe+Mgtdk5WeiHVx
7Wh134qA/ruEWS/ky8rlpisqTn8+LBguVp20c85AuRca4QghHH3q2RXJUtBjElee
JNYVb8w1AOJLjVNQmUE7Vd/gdd1sFwbbiq6T0/4MRYi6bdpPaZMmztygUc7LK2Qy
piT2buuzBA8PNnZFyS0akdMCD+h78QDrK7lf3OLWxytAntfe+u5Aa++2QU3FULdk
i7XlzZchaoXk6Xsa5+2S3F0b/XCpK6k8dz9S1Ipm0I3A9HDO+dKBgzzOsgR0MkSm
d//jH+z2J31iW6xbanlZkWEJ3LpBwl1cl6Udv0aGvoVgUnFmdMXpm8VP0c6moVuy
3MQbvZlWBr3Gx0+5xalMo8n/ejDpmPMCIUJtD6sl/hnxHAew/rdhYByJXO+SvDBN
QTd+ENIIWd5Qq/5c9Jqx1fvZIR5tqyb83/Pj8RBL8aPdZ7dcVZNaXHvKRLu4UT+C
nkZYGfzq//zzS/pJwc0SKvpx5AA29w+Bdnl11CVqBtHYk6DXAeuVhQthKvDn8Zgk
WBUu7wwESzfXx33EtZqzmz4GFlRvQ3Ooqbuh2VgIAi0ZUx4t7BH6xiNcdEV4dNA4
DCN4qtoNMr6XUs7setIblGZM692i1d47u9KnKjspSLlNfhb/ejgR9G85KwAVP8BO
rrXu81FY0+Qz7ekPlgmqF7LvvQ2OXOTfjkM9bFHNWHi6E5MV621GkjareEseXBJk
xST0eSUAR+PS51USJIDKWs+IqbEmpFFzMewOLBtYBnPXYoftfB+KJ1Q7x2p7bSVu
oIMMRiOnZSE8F27UfIWhxMKHqliLei82oTFCc8C1frprG42JnxBMcaB2UQSEj4Ne
RwpInR2HJdGB+os+Udccvdt1/gLCQSMu9Mg6DOp7WfpxEA1KNbf11KOK1jtaOwGG
z4TBYA60FqfA8iTvidh9ueBKusS2dgdxivanZpJOBw2z5Z1cdJHAK1Xl1okSDOMf
E4LqRCfg1HEKqaY9DTo/W3FJJfEczpGWVsTEZeyNzCAC3CBd7MfdGziCtGrkpODA
7BRhjDkWOQNjoMcZM3THIJ9uOw4VJ+E4IfG+0SX0KZ4sFz1ixL7kh/hR9kxTvcD+
Duj3P+csG7l3n1P+xfPDd5blO3reumUSocAdAWmlkV24oJwZ8ktvA9AnWz37mWJf
ilIW/tZrVQm6xEVfhC2RD76UzXA0uQXbOic2eGpZVUGKiFkyGy8GmMzII0G9o0vI
dTOJX24dVxxF3MVoJfWug72WdA/cAnDO6jEbH+uCu60MED2z+kxHJy4wxjtuapkd
1u0QMEVr82/IOVZTZCVbx3u7yU49y1roIr2oIPgUoHno7AEvZHoYUsfXxHRnwmqu
Uw9dcszgYPx+R12818KgNMy32JQ1a/Cg2/ZMGLVuHv6FZCpZqNnQQb+nA9RopdUF
sf6p0o6xdfv8VM9NLz3XrBSrWetfmB8apejLZaZpQ1L9yxnwoKjUWB0keN58DlSG
esLTHRnZSsYjz3xn97Q7syol0K8FVc5LwB4Hxaq9rziOIUmwcbX60GCeKHoPxe8t
0TEfwJflk1dVebi5Loac42XzGJZVQdX8KETuUNTkaSvH06KVFjkzl8oqQxd2Ok5v
PorQN0EuH9a7a3sRUiJJPkkRcWBsIjdeoaqxElREbUhJ5HbYd7CkFZj21zZcbDKs
INAEiefLJinCRdkOJEY79Nbrzhp3rJodlRbpF1uWGwdWfmX/rdQ7zcTUGCryO8YP
RYYZiUDorw4Ac4EZlwIjZDGNFEjqxMSkAetlDIpuTEwcKxLCPR3xYwU6oGi/+VeE
EuMHsxkHeZnjGnvAiX0slDpqWoK+apWsPjAfaOsL4+H1/sEUQnLRrhUBKUDmHL2I
ciS7TqqhiyC3ax/Dr5Qq7gDllhZMpmeVlyGbZUK+GS5RVbJJhIYjp/zwEdV5zz8l
Ou6T01qNgrqULpKXpd2xfQtHfCN4v/yl5YdIhc1wIZJXsA0zdBgi3uZKtrRp1R/f
sp55izlv0jlz6GJAm0rNHVd8yyg3XOdYkaPHc35NjTJLk7ZuVtmQSDWSLvcSkeLY
DEwlFKXMmTptuBchYBDR7CZ7vCAFpPu81nmKHrBTCr/fdAI4SHIEqEC71mhebs+4
MrXfp8DZOok8IQjoi/6I7upFYgZzCcJnuOglPALlmOqER97xKzpXjwMPqVAz2U8j
nVaA+8x4roOoDXPazBaF+KDArjHwbONlsqauiqQKymx1MG/3uv1hlQM1w6CJ1qC3
R80MK6a3TFhUK56KK6AspIoW1Wk4ahKCljlS0LdYYiUSAtmclOWTN3VYbFuVuVcT
zeuK0KCVvVFOZrnU7IfNBJn6EaD4hcq0NtCEznWQmAgFvZOYuZeONyDk6ffUGpzu
jrj/RYLdzwLW4IrU/5jWbcXGg6quJjqntwBz/Oqdp2Xa6tBVS81o8a3twl/2ExBc
h/XP71qORdm630QMBMKsCHoqmurjGAplxGpLKzKpfw5zJ0bCH9/BEEmDQEnjbwBa
ciJpUdgF8O9z6bl3DckPOgOrWxUN3WgHFGM0EiUO7hEVFOG8E+CVk/oshXVF6tCy
ExeSzqxchYnIFWa+vNO32yRSz8Y4wRD1nKkwYZOCb68tFdyrvZjVTvFoyUfqWppz
J96ZttEH3FeI49upGfHZAF0QqzvvEycweBWwYBeHb7rKo4B09fQ4ebFrzgLHxSx5
2BUkkEK1DqwkHmKZlO/743sp+cXm53BxAFC8KgruMmy9Zga3yG4dl7IYufZUhouD
f/sBOP1q8eFqYkOQ82TQd0/bjd8nD0VS5xv6feinDI+ndpmGFhHyC9VwB3G5vPcL
W7RNt/9PDxxlt6SR+BaQ/sXvgzX5atvjdXg+j4ttceXgtACAYeOj53DWs3ecWSLQ
3FmsB+29hUEx0ynh2vslxUZIEA9VDYBxAccO7qo9rUEYJVYK/JwJpDLSFYRnr3hb
kEm2udk1LcHEqFOKsZfYNR+HAz0+UmTuKCRbFTaAtI2TFjbQ/nqirXa8Pa14GzSD
xc86wVDbV8CG3YJJYBHwPCsJzt3fPHoZJxk2pZMOFmR3zjPqkZoAJqwUBTBM9tAb
lY2/72iMvp7BlKkgaNs5xxPeMnKRT/CEIcGf8RMvjPnxPWld43AfICGxHBl8Y38y
vW3TamDSc26cjAq/7s1wjNQ/kwvxEer+39ZUgChFIgZk1Jay/22qepa6LGW77uPa
NvCqnADjKAqez5A9blOv+m7ICIO2u39ShoNkFTbi3RYZvmwTun24MghfQ+tkJgQi
t8w6Q6VJTw4U0lo8kPTq0b3dAjCheiCkbai6LgonpttE7Um1HpKZRWj/V7gXdPz3
7UQ/6e0CgTMgJprvxjtDIOfzEGmGRlQ2t30ZMUEyPVc286KsXvR2KNb/cLr2CT2l
eKO51K4kDSxNalPiLsgSMvbQPfu2RgdG5yagWH2JMxkF5Asoky4hXJRPJiGb/rsK
3vdroxhQKaqehgGfpfJLsY9YiEwe+mvK7YkVPS3JQT6Udl+hA0t5z9ReKvEDQRYZ
TBLePuLPm11V3b0wvJyfRm/3qVL2D2YKV1O46c6x10ZWPQebSSCK5pdOoKOEJw8V
j89eWEY02b+LeWyQWZcr+OtxJ4M89yTErpKZ4uXN1YhgVXy7cTzo/twCzEXVJTW3
MO/SZAt4zu8XQ+nyW8J0FjdTuoTHDMNgJq+E/nysjfwwHbbRUq+fg54FBXL3/Umw
KVs9MX7f6WAsyrjU0ARPcNOLHLOAmcVLmRQCMiLzkD/VBppMlazfE20Tgj1+rRTX
RgEp2FToqzPc9O7HWgsgJptEUn3a2VSOR4ewHMv34wYpJyze4Bc6tlsHZ573AAZh
B4k4+yONhZ9bFoMu6DfgScPGPr5qMJQe2eObtGlfyrJV65MCod2063A7LodlpFNR
V+IgN6QylJMOXJ7xkrhi1WfqxXO+COXwW1JGUVTSQW9nFLqdIg432B7kV4tiv7JV
0wPocBMKTAi5GGlQU72LhVQJug/M+D4pYXkGZbdcVQMxRfbuGSdPRy/T9mWI0Drq
FffB3kP6y3+QXwT/ACdQUMnBbnKn4W/IFbKkTIjWob96tVor5+6W1kta2HZx6vTm
BPwEJ8cRnmvEeq7HCvrfZOdQZ1SsDWUoudNgHzj2zuLLBY/cjEuSr1SbIE8U3mbH
HFIzC/4MrPaf3CSFcIKWWlgmcnn7DbO+KA43uEVDB39suj/g7sSWM4Qa4hpg8NCI
p2YELWn7xmnp+HMwR7weZcSla8W4YpEEOOMMBoPo63vj5fbe2BxVAsRO5fPz0q8I
TDQdgTIVlgVatr4eu2VspPwyCy078N3u88+qYB3wi/NCX7ySB7ECjUmLBDb0jh4o
ak8FAJ6Rr2fI65faVSfrogLKcVl+feNWdZXSS9FIR5Xbjm6grVNtAtIvpwJiHkLd
ntn9JDavXjRMjI+jmIhs+HtVvmL0y8Gk8myuPhW4craUlI5UT5sC5s4Bys6RRoml
zmMd0QjntPUIDZvErlDIOH7vV2AR7cNxFuxYXg9CC/la+N5yn0YEu316XHmormz8
mCWtSP/D2mPJqIIGF0FFA+OUEN0KiPtOof/sLnnRVtFNQwHsRlLy6jHOyl9bh13e
VUDnro1HNA9PELFtX0XMY3ORVb5AU4vb9mLz3kaI00rBy2S++OIiTMF5PwvOdn1t
iMQGPj9jD84sEvk5/lhZ8p/S3yDZkLhmrqJFvJ2VpN9qXzKQ6gBrSCQV1iKEI3Ap
UO3U4T73zjRM1MIiEz6HOmAwVCZO88G0lF1ir1SsehK2qxWvceu7ePqE6VjksN8t
W7MLjOls2gdnNhSv7OoU7QGKzU2vsJBsjdFXIAE2JJ4+OOB6/EdFAJluy9amGIhI
oRYotJZgkHaFNq14IEl7nD3MLe++c8KZu5DFfD0MRl0ypzZazuwxDiyHXLUjvKx8
9UHHSdnmrnc6t4cUzddFCMr7SzhmYIyyHXv2kDion5Ev2Yrn1tpjoYsqv77WzIqY
6ghlH0S3cT5FpTtP03sOWpMLdC9McYvaOe0XmQcgSsXJA5J5mEjTEpQQPWyQQF29
iO1ZdxJF9BYU7CwBd6tIBpJWVOXrHheVb8xo0/ENEP/syp4Ds1fKOqC+gbB19SrM
KCx5keWsRBoY0NaDY74zChI+YQ1QR72bp0G2m7LKYwXBC3hhG372Q0gPwVhXEvrM
x+Wwxj4fOHbm8CDVzysFDvVfg5WOBOj7hes5o+o9/rKPykta6h7mAl5LtdlbfzrQ
4358dq95Udcc+WWxM7c07WUwXarW5ZfKqT//z8uGD5bkAAd5F8vj6lwt6YHTOY5N
I5VIgieqWDHJSX586sirRs65a8gsS6AI6wbugHbZmNB29tWsrp4D84WFxxmFTdu5
Dz5zONG9Hhy8PX1rSirJH3yqfZ1Z8+ZgwRwOcgu41D8nvULQnH9c9XOKmE74mWDB
smAHmZlstsCF75Vfto3CGANxd2cId5YH31jk1ta3mN8cwrAAQ7Vcpw4MXPzmKXiA
w/4A8+XCJxcSnquHo6GtrNyxyvaI10K5/dSEeiokuTG/XO43+rb4nzawg8wGFXGy
Ph8ZDI5VF5w6GsaszGOWMSfg4mRwnPNdfejqWgOsytdMr/UnbZaOn3xKBR6G/z9b
Y+G4CZhCdrIaNmH6n+O96RTnxq4THQ0Jato8+u0ZhZRGf05JxWAyewbzBW7pG4cq
y0vRzi9rSQR9KVxqIdLr0+OqGzTeRWOLbdkqgAFSHVzwARhTO4NwScidzJY0HLXS
8qJCJGd6vaetHaSVMuaScWyqwo/tXXASsZMthLjXtWp0AsDRu1CwmoL+zdx1D1+C
+igvZv/AODspF4vKI/sOPqmtGAp8yHPDps4kghYl5CP/abRTthzLKio76pCHm/QF
j5VRIUdC9EoaGEm1+nT4OQ3N1NFzptrikuGKixpe4QT2wkS8XIjoPrxdUswYh7EA
sbvJsY7W4C/jKQYTRrpVkRYrDofJbZAZ9gNQgCd5EICZPQpSHOdzQh0XwdSmFhyg
t9l2OnFYp78XfaPRcN4v6T/smBvWnx5gByIPz6G+CR52KXy3l8GfFjjMFbT79MoD
JIVi+AXBGoZZb9dzwEXI5IRnyIg8u6menyJ7+bBTPopRC8sBLtd0zlNHLtA0wY52
hwwO0deccKdHyLUuSeoWcJLXi8jAySo20XTN1ZJqtxBcMQDcRuTkCmSibsqRqpGY
QAWiy3rutTbIX/Qb11IcNB8cq+TvTsOM+LKkH1dp90HZlkNvf4HzfYE+HlMj3H9E
kT2Ujg5SIRu3T90pUDkzRk8pXDDy9ELR24ABXmAwT/CFukX1l6J0cuF4DdBcykM3
VI9lTBOl4vrVgPQVt1aaAdpuWXuQYegJKXwcFdJ7EMlh2p/RItvWIyGG8SziVAgE
rG7zq/cxKa+9Nl45jNmMcH5wl2rb2m4YZo8oYZlQOhyDqpdjVQ3NkQ23Z0WC4KkZ
q/hxVb4vp3DfeGZ25IrrnKMaED4Hm83eNaP6gcDflyjziqT1ejmcPf1TV+a88FxZ
indxRSUlDGOZTi5PGfcxBGxEJy2VIpKl5JrDeZR0vgySlmI+mUroybHnposjDHGY
CLApIIlMUbLLCtFL51jCzRG+djEfnGhj5KiuZfmjWE0WR394yTXn9yuU/TPK0BpW
pqAmLnus64xMCmbbnQj5cUmBIvP/zjg2ydvhI6t+oF5TRRbnIbXMztv9ncXDL0Qg
PQdwr5mRqNR4dXTbAE3MHgTEWBBLh5h3kapDCr23N2MqG2CXP2jN1Zr/BHv0WPX2
zp2FJTuV/EcADRAihD/DNZQff18tCDNCfiETlTGNSq/KZ+Ew5KX4ke1pPD4rqRwB
y762Q70jntapqxaEOHPIo+wmZz6qsg44HlYHncbj/MxCuU8nRU5+oy4dEg8LdfWi
h8I7P/hgy+DPuCKGKMdrRiYuSNuH+kNslkacikrKwTl/r4cIWqyM0Xgwieukq59u
9wZdmID0Xm2Y7K0y54bkYzzKtgP77GIwLRIXemszKm3EQh3DRTu2rqYmZZKe5VPe
Uf1GsSCFa94GRNk0mBpKcztHlQBhQs7y4SwRPFa5R1dqQ/O+mCRZ3cHKsP1WN2ng
v41Axzfmy7d9eE5AN9oEmj2p+Xg+Y3KWoqAtBLEudZ+j2xC4grbDI6jHBArFzUP4
IvbjLGJRQDy4zVL1Dui87Xabw/6z8zHm3W42Bj5PW7yIqmmJvE454rw6vJUblA00
htzWm+sEvQ2P7ZNC0kCJzFVdVuq4tLKaQLigSGeqhxZtQ+83jLqIEJayVIpMhAGI
bm5fz3YDJa/c1sqVxZdJXekegbEDSYwveVelqAmsVx5rkVGPqgyLPO6jGfpiM3Gx
ULvxEBhOnYnB/3m4pDK3aGdyz8KlMdMEIcXIJiY4X5dm/Kwtth+8H5HQKIkELLUu
SJXfB6poiFe1XTrCvSt7qjganLcUWFx6uVuhZ30plybim/XJcpRVUqlz93HA1b4w
L4NQEohs90SBSNWio3mtStmsMrhhhXeXmpvkeJgmpg5UYZ06ZC/RxWT7j2zacDs8
4uZv2pMWZpG2+F8ycnTvM8fjENgpheRQVAN0awHo7BlSzGer3lBTTfdseF6iqkRV
wMU8yDXqe/ihLagugT4rIYK09n0Iq0HEqxld1lslvXiy0jkvGtBsKrkPwEOsAxu1
cJyWEWnoqZWAlc9gWMRy6EHfmUOiPRAYcSeUgCeF0j/1XYru8WuO+zjeK4qRP+ow
2s+Mxp0+Weruj0EmFm8rfl01smPwuyjC8HSfekS3mNursx0fRA1RkAMWB4yQuml7
FTkDJf04Hk3TrY7wCcZDvZkN1XySszttA9kEGfKJIItDzzbka4HMaS0c53mClwwh
8n/FT2odvAuV9gf14Scotakvs9uRhMqQo8K8yFCp+59Qc2gVR5B2T+kT9fNtzT4I
s8uJsNKZTgcCxW47i3LCvVV9BhhdF7NyR6Yvfnq0JaBpBrejKuHrM1HVVVoYpFYc
JLGcFXGa6/JS4tmyJo6xvl5XVg68+K/z0908mdwBoVCXk193VjidBW//egKVCX0F
EkxVxP9q8FfmYrSI/h1dENUYYIAmQqnO4FEzi1U+IHh74vg6ag9CqMuMPzCA5DLm
Ijfepy92creRBkmzRCUGwZnRkFcYfDT/AToEjjy65JX9PTgy2KXnaaM3VZxMjB+/
ZuEs+rG53vwe8A6LcvI+uwE3hSxqVeXztZTKNCYH+67GGn8wOjIar2aXMppUUakC
iNo40j7XTGZV68hOMSsfwCXU8ogYIPKJITEFqk0iy/yEqoOA7RkWjbpOXD2Otvtr
F0iMWwV9tpKsuB5gEUpXDyQK8CmbuovF7Bh8hbxdUo4uoyP2BrfH7cU9wjDm+eqX
w+T7aP7U+/f9hnLT+cPFDzB7v/feaBFa85P9/hh0QTmtaoX2CMzJiOJfDI8b72S0
mdMJeQ/QYSX0LcgcnlzhldjEPCjE/439lzUe7s5GrImFAwKjhvVU1dh5VbCLHJnm
2sS3kYumMfF0xB1rWkSza+ju1g2+UlUlQaJ4Elvo/ovTAxzznUkxAeQD2dM65KZH
JMlwH4T/CRBOdiCfVwLCdudkxssitTZGkE4K+bBfJsOtGM4DOMdRUgOO/SNwdzoI
d3E8XeoKCNW88AVlBYEeymVbfWRqR6gujrzhwnIio+CBkuEfi3zSWJCTH+ZZmxHx
a8feJb84rk/Cs5Al2wjpdzAjeuwB0zqOD9tByiTzjJwI3KdlUKfzd9lyRPenNpbO
GAPTdqysK/IPhEFlVAtZlGDqbgVObyk6m4+YQJC0Ag3WgOpyYj8LLfNYuWatBPpF
uSaL1hFk/rTWS+14hdDMcppguJhY2y/RaO0bgh0RrUgmDknQe6ZX1JpZyYQQpOEm
ncHAylpotUTbE0jtL6at5jbFgp6qIAim29NB7bFmk6ni2sR53ZAHkjTvnbDqYBDU
RVBU1wmJS4vxiPjedyYw5CkH6StpftlCxGCiYz2avlhs9Y6Evzkmhm9kondzQdo3
eH+h7cEsSDf9hVnykrJbyFPpZl0hnGeBQMyw/vlGoKdXLh98GB4t7Fjs2PtWcYfs
r/XJ4KrnWxhx4UVMCbCwvtfVM1hjNDtuipoMkwAyevI1Zojs9iXVHYJYqzGQ7BbC
XMvXwzsTYow94RWCjO2dvozh2YBW0FioPfRPo0pV5mL8gd3ThyU5uzpbJ1bDrbAO
ZQVY5tGdJYHkxHusjGyc2SixF17yukMbajCJFF3vdRLJUJ1tw/Nb4IDI7WRt4KZM
ihuqwOqN82A+UOuy/KyF+HMpZ8jUSFdUZwdAjvKyM7H2ZzgPWop6ILaesBbETYPu
hH6TG/xXr5uOD+Aix9VvBPV2B0R2oeZr7Bbws8Lh+K34db5o15ypJ7wRaB840juW
9fMeGfpgHKKsR8OF2DLN040BITVUlfsGHt49ZqrwDXlqbwoEFuBjjYstZ3xIPMPX
ZXa2yMQ+tX2gPRwdg+nCGXxlH+cjHfUXxA/3eBZzT9m0Nh6sskwlNh7LDBdetE+v
6wNTcuw9GbWCTTUSk/eKajCcf85j8cz8otkZj51OENw37deuyQfWTYxfLM+vYQ49
uLXyKlcKcdrZR7Xkd7mq8IVciwVNAxZqMEIE6s1W2q2DHaWFBdlRtj0exKvmaX3G
q3v/nvN7aAgAlTUFl/7pRZcAvZnom00MZ+i6RO5RAOcZ66HONKLndjyRv4KNZPue
SUYttBRDWI6BjNS3Ks+/cBQXJLMdU9JkqFsaa9o6DC9CxDOFg2++v/Hs9/UxNQsb
VOQVD1/XgdU7hX/k3PYejdP4KdlRI379mA9uqE0Dg6u+8Rk8RZwJuzJMO/6etzhf
/N7Rs0+m2h3O9tfk9dr+ctEh872WvKUgClFPUQtYkHNrPjk3B8yTKe3RGzzofsvK
J51hy4n9VTr8/RXoESyjFoh3L4h2bOk8f56kZhEu/NlN429n1Q2Q0y1Np2OjHM/J
Mr9pJSoUGHYN3YGYllaX3SpH5urxNcZ7Y20BfSDmcasX8IVP9VZOyYj/UVOOJW25
IpGiD6ZVLtI4PNdxrZnzfKnxk/nEeu3PnBoGKimrAhTDRzlqOGtgqhZIEXzXI9Ap
Y/7OQcM4NnEzDY79+z34+lQBIAda4Flmol80SOVW0SJLYySOHfEpcGF8zMAPBBo5
4nQWmKZyCvQj7juJ4NQCxUW2Nlbj66s1dzZ5PlN6w8grs7ZmLZrkj+FTtwXgA58U
Pi4tjh/FIj1IhUn7PJtXx7Ucl/FF59kPeP2CsZs174TJguiq7pIOvVvZijEWBJVk
NJ1+3ze7jFSy2FeQ4NcMfHd94kn8i391wp6AirrAHdbZIbqUIgwUITWydRwhsXVr
32MrOKXRyOKUG3n3QXtD4kPLkVlaBNLCu3VNMFJNHEZ98IwR6elyG1rBC26K52BT
1M/D1fox8A7opWf4XiP1ipma3+I4a1olk7S29fXknAOYJJ7kytpqQeeecrLGzC1X
o/S+eVYhNPY+oC3Y5KOE6WBkSjx776sjjZ96LJ7RqPibxBUh6GND1ikBwUGvHWUt
g2BySqQu2EApzjJhAaoHlRmYpdY42Ql6HoztArNde0p9vrAPX2/Zc7xCKSUNQ/3f
z5LXKftGBJnDZ9BOc1qMdnD3PvoB+A1vcgDZAOPULFH4KwqSWMA8RYQBPV40PvUQ
DkmVp0KNW07hAgR2NR7UlpirhweJOdUUlNAoAj3AYB8lwOeOxPv+CBcn9ef7taim
VzFoUoA6pZQgF4xyBj7ijuiMRimOLuh6SQFLnptq1SYSEQrOnzzE82TTAnghxIrb
21HKg756ZNh4wKNly5iVPShrUlecwQKPguQCKo2oaqBF6VXf5Gd3YEAXX4o/nHbN
BQaSGWFZ86kngIB58n4QGPM5bqOFnIiO9hdUm0Wg7UnfiwcHlbytPylT3KX/0H7c
jjIVU0e5PKDYd8Ot28tRscI3LCxI4J9z9aRcjHndtmTpfn0x9Jq4mJSTzWUYyYpR
cviLxjH/FicDlJH/syp7kl1+qIPWglt/mWHZKfepGanDX8VTG3qrOORnC8lWxwHw
vxT9CUsBO8Qhj6AROfDvThzQom23ysFPB1XtP1NXmCBJYqkGkOxuDLm+cAz5kiGb
jwTzszGTEmOPtinSkTrTeKZl+5Jyv4a8P7UuXIIux8U5oY2XNVul/2fvueDRYDVB
hf5oCvyEJfOCJ8sKXBh902cKC7cDU9vztzxjV4wLEoPDFgCfoTaz3YSqTwK1EUcc
ZJ0x/cXxj9GuBWNCOK1M24suORm9YtEDQrq2HLHVGh5viJBCEY6qzXz1R/BK960U
lHbzcI+Bu/iEQnHzftf42hPLBwRCsM0/y5/Sov3Q06XUAWa9XRoyA+pWxurfMZnh
1eAcmtoxxdvrswHdFzRUe0lmnpcK/cY1s9fnVftDLRYDdtyZnw/s+FvzLA48eoNd
EleSCLwhdi03caruCuYLFg6gpofyWwM13XobzJ7DiIKHDAGrFbTSk8THKm9IPh1V
4LnCK21mbfmYQfAh9kJasUr0nTi2IsajgSxKLODebFlWWY3SG8GlFt2EK+gUKnKr
HjNZTriSftSkPw5j8og2PKt/EY/yh2zfErVWTw7PRAByWth0tpJuvZ4TBSSpWcU1
rFzSyuPYokPCCPuJce3VU9Q/hViUDOnM1AIKoXaYQxEoGSOTG2V7joQThaljIAky
h+q5SqgRNPV7EjMD85YDbZCZ20O48UrltfsO0FUv8M9H7BLIl6UwDmW3gVdBcANB
ItBENf7IWwGdvJQdzsMcL2xW3C/2oPeT6pi95OmV+W0ELAfMXdJMio7OLsyZKLLQ
CN5D0PRD3if/K1aFvwvk61t/p90oe9xto5MfMJ1WE6qoX1Vg/S+hvjtWhVHp+8Se
IcapeMNzWORVm+9SEpqTe9zzBUB2QHg5vCB0om//IMDNRIArbJzo3c/RAlSAfmN1
ofQs4VNqq8QnfgNriH8bcKUu0DqVq8WJ2+9CVCRG3YofV2pwMHoDDRQD/gGp32wD
1ASg+7w5hHrUJgPsUBj2BSqCt+kG0yV3OuyqiIzsSVa/wLoLfXDESqlnviejS1I0
+dfoX9eShUQ/sNhCBtSZpmQsSfgS3EpKDfgQg/vNGPlqn2GqLhuMJZbCJyG8SJeu
xtLKc0AwnYZs7XaDYM7CaLdBHErzCTLIyPFmWCSbAmaq2iMW7PpbVbRAkRRl6Bbo
9OTXjG1uzUS2pS6NeKVOyXdsstlJ8KmKF8RLl2++l4pP9AdNrGTUKaoqfkTGQBXd
p/qrgH3BLmiZ3FgmqAKtrWeD2CwY5fzQ3JhAWY6IoSr+CYfbPNRyU4LckcqPBv8l
4IePzVrkyKP7k7iwydr5Fplmxki2nJuFJKQPrRQSpPOVynztKYsc8OVzda/n0XnD
w5yXUyVglPCRWmJY7S/u+ZmkLyKznrxLXxa+wL55KNzOxgdS51dH3pZzhY0ta81n
jW8iZ5sQu76nz/NFiHMktgC0fBoG/6GluoVzPrVaRgpu+ss/T5svVmXdZTRlBfci
VTz+i8TLsDBKcjH3ZC6r6uVj0UAbNpUhuZvz+etvW8BhL385q/zdPymobSxyvWhI
nJAI13fzu1cQWrnidI56Y5TJ1TM74znQmaRMAmgnJdTjCNEYCXydCUYnJM7Oey6p
s0MvsDSu3a5p4jnopwH8zbkGQ2NJbYnEtfOjnWjsv8KfyJsr2TmUS5R0W8ml+7Bn
gj7QMhEYtMlvLuF6z+ikbT9zS77szWNyDhN7KacMd4JOgNWZlcXiTHOUSvwhiqY8
e+UPjVa4RJI+xzoXeZLkNJsJGrB0GfD3l8KNc5i/kcW5gyf7hI3UFCq7K26aUao6
0598IjYp3f5nseAgzkvOcpn49KKm3F0cOisWBJup4UZjmxVuNrzkN0BwA8AMZQZG
8MjzVDnUXX+uFx6JX9K7jboi8ZxDTopFFhHHICDfpZ714nMwUFMRJ93EqtZJff/O
taDph8zP3Fj2x/9al9odStOoksl8CGZ5xZRSXQMOtPpDi5ejGud+3k5c+VHci02j
JlclevpY0F1pVtLrUAbG0Ml8pDrVlS/VWPyWtpJ8cNf1r/0GWvtEdRgDseEW/FMV
Yf/4WL6j2b06Ksso1ZKF/47D7m4yljQ8Mkog/pdeRUVRjg4ZhZv5Rx4hcUOcoxA2
eneLSATUFReZTTKhdnu6YEXL3DwmyP3ejIAZ481reWp1kTlEjvIv1hJMm7O+25QL
t6G2kBwb3eO/fD1Ud6rHi0o/xKCiupnJQjlPLcryGkweBYPhxt/9lZyA0fqWVv+9
Ul/nVLmvaGk/YGNaA9esMjVPzaAkLqKF+T8yL2i+Qeqag5xO/o/Mr09PqqN/JmEN
cqlYraZ8EbhNf+QoaaQaKWmnjRpdeseFipeLyKaSyJeHRcVJ7nMlPksrBtzx5BRl
WE4FizCj9Qmgm299rwIQVFsIzzUC6XRiCnI4JDRZHhtaGM7gavcqzJm+TQ7lN3fp
Zvedi2tsuVzd2bGNShLkruxAN+g+tc/MsP+Y66PFT8PiTCSVqQHohr77Wi+8OePg
UyM0L405d3xJ2Yi2GESoBs2eZSsIcVDoLcIWigtE/KOYQxM3tr+jTL8ZmHFpI6jV
nOp+J02LKRopYmW9IYaUb3Ltlxk/LNIVW23bZZoNFPy3a1CjvaMV5X1pde2QswRB
CmjlO/5AIs5zUuAtuouc0ESv1szt1UtJ/4+OCrpnLhyCcIVfCb1a8k/Y7c2pDuwv
iDKhsJG1h1nvr6qohdTwfj3yu6IDD5eLkCnNc8wOSPMD6ju9oUQCiuSHUGEYB7oB
XEuP459dmBcShUlBBBIgZRwCTQ9Dl4YidGFBcgwWSZWjc9agt7kHPnemTJOxX/zM
PbLOtZtMIcKHe+Lsm11p7tb2aPz+5Vg08rjrTGT9oJKeZ1djpDaKGfMPqpMnmUlR
lnjJ5dkMh5HkX+fOY+tacFrSr3zNKQNmhkHMDvpBbGxFWMpPdeNZ34+dYuiDjMCm
JkPjONluFYTqRLJcgxIfMg+8si8NClnn7qyQA72cxYNAXO4IhC5kRqumjcFw9CjD
txE4qZuXFrtSPWck4DJJGt3XegZOnIybHX050esMWoC5mfk5Nd/cRGgJTxAZygfA
LPHfWQSrAkE4YQld8Lo3xrPaSq5yqFAaIGKuRyEeLq6mjC+NU1ArlHGnYQyKKJkX
Tpqf9kgFumqwsFND4EpcliHkLIRSmSHibwacBLSQIHOpat0g2ViV7yb9/+qgf6W1
/YbH7bpPiMXdLYDICp4tn/piu3aSPwHJtyzppf+CCKD0/PllkUHN3Rwd/flNtD15
bQoax45JEwAvmJBBnOPo7wPfbT3BJMkpHm/+WbOf5dMD0Ft/9yP9ukjVdMtScVcR
dn/kkL2nw/Tj6ZaNYTq4jkMCZLP9VI70nQPYtMk1EDEc0Gt211hFsUS7NQVbxoOz
Hqq1X5ymFT72XDBvtZYwFRW/wbk4xyp29utAdTVX7bRvWw/3z9jhScSavZx6X7Gb
3kSNFYrBDXqn7ZvD+U1c/hBQakELZ/HD+HMUnU+/ZrhaCtG3uOTTanz8R3aNJgw5
s3uKj9TV0DriL4b0Bkc523JJkp/dgz4Lr4gBi5d+cnaQHqbjqX97Ey1Iwgrgif8x
NEk26vkT+MoRZnS6xUMJL+e9JeV3Fh2wcjACHQpNGls3YkrsOrN8YPIbZ2Hgy+I9
FbkxJ/wx16O4TaDdWJfm9wdYZnDounzHfwa+dErmOaOy6V6CBLwxf8mZ0z5DzMgu
ED19YNb2Reg6QbNZX+RsiqhdLk407koa900oUxeFBftYr/DUDyZegSm8g8LmHw7J
yaLX2cjyX1E+XaAtzL1xJfyCOTP/nmOBfJsbK+FzI12YXhQEm2VFtMwbbo2o5irF
Qn47NATlJWQOXYlpWsSywtMTGMbpZp1B9DTksCAXuDSFxUsJEb3+VKd9m/nkU6bZ
iY9jsKD/tMCgGLex1rX3BvsOJbZMkOJfxJyiNSykl8ng8pYcxnet3h7dSYVmIN/z
KBxW+RoKLvc8m2Pm7jJXDuApEmP155bs8SeuQBv12DjQTP5+N4C5s5cRyIkl9pdN
aPoKTbwjX5c4QYmFBbuNIHzJzq6IuAjMEoq9PCh/UcYgHcLzuaMV5QFMnpvJueWf
Ar8mqSitVR1m6OtJk/H2LgP7ZoodlBtzlU+FaAocFaoSpjsOOMqI7HJdOSUJgsqR
8xqBAEA+57pIYSvyBpqij5JeFL6RN/AGxBkRQcP7Zhg/FwTs+Bqz9CUug3DNIMcG
Rnmv/XX4jLxc2KRg7fny4Qkpxrsh2YA75TnVmU4e6tQUDkmNnIPAVOIHr7bSZSrq
XWSrRcWdnB8P4HeBczk5U2cxON33IoNGGCO3cqr3Vl+xqwavIXnn4tPOrWWpPnV5
4w/6ROzb6pQDiy8ZtfEX7KZoa2Wpoahy11BtnHv4WUsaNawey8oVj6oyqDRnmLux
mpMD5Rv57stP1a9iMXTgbgA5byYurXd2fsqb5qg7DucEqoVlkjj8B9DE9qCzEgoN
RTYdy1IwjAEyD4zvzpHd1gv+BeEjpyozA3KPHfzfxHZhgMWODLCD8gEcPseTKbTF
ZgpExN9F3U6hy3X4Sn6UvN9EANDe9vXMgsvmcWidaA6vSBJEgd5R1L7vlgTnuEov
KVtGctBaWR4KIkDd7IXEUO0eo2a83i0Aa8tgGmvMcAZnqRzv/1NRluf9z0VPT/Tl
m6xMbt+nPZBt75m5mI+c5jKc1P8BPe2aGPufgi1OM4FykCrltPFRTsT4JIWGYzyj
uk23qNBrNg+SOg97vu/bbBOUTs5bJqIP7Lzo4Wn82o9IdbbQxAATa0aYA5C4NfKP
xi78uL6m2ZsN0gFrvKVKvfIscnIyHKAfl19eG9Dcrgq2eLgrm/tn7IzDVCQA4M4e
W0ia1PGHMVKD8PbgkmrEqTNQyeT/Fo8pWcJA3CiQhUbD7rt+152Dt8l/BCdcDodO
3lFwvL913GLa2K5UXvxWuW4/1cVy1obXqpSwATQheduUthXMWHFiG3wR6g9yHPEo
76ePxEsnaI4FxkKZ2WcsNqAiFlqqPSool9jl1SLQKMpxvHhn3gqpY5oZlXuQv1SF
GbZLmsYmm1ykt4KYDTI6Ss4CbhBJqtqWjQdMrwp3o1kvjkVZ7TLFtZsPwwAKrOZR
ujj//bWRs9mWAWdm7qR8veHgh879VqKFPY3NpFIv59W+mef7pyT/kcglAOWPcrl5
1hMnd6t9pG0lGf7TRliyG+a2VzMHXxwseAWvqGHvPDqYbXJbVtFYfNtp7ZGVIsWT
s5wBdfABZm4fDT4RDN6IidmslHXZgFDizfZ8NkM6L4dqJU3973l0a+NcQ/fn2lKG
2W0mWwiFhK9f235gmVpTQebdom0rEwg1nf6yx+9RJ3D/lsVuzm/QNNvlzylSumCD
GpudZEpocmDn/K6WVt6ZbQrK71KIN529VexRFDjnqSaafF1p+Wsflq0HTPmy0Zu8
/9DMgrf8BqYIwONW3GLGP7rhsBJYcE6aGFAP0BfFD+QQqbCXUlxhAyx9ILAO6b2e
fEtNmnRWglnXvbrA65xQ3M78GfuDImOE2bweYBE/MiYGhEDxpVFCJLy/KWlBbKXO
zw+9PGO+STqgzMAScSY4ZmWZdLCgdqVfA/K+aXl3/tbcRHSv1KuytwY4fvSPMeB8
TbkN4ZUxFmqTtDZAnWfnJHKiy5vd5XofL1Aa3IYHovPDWZhsx0rEmPjs+jnq4mYK
qTR2f1jiBiXMH3Pn/qcZzxFt9Zow3CanR0IX+u5aMJpJmIhzBNlU3EbHmZpcjAv9
Drxw1tI/LCaGsIqkT+F5XG3ZzRKjre6NeQKj3e4boUcdku9Jz8owa5OmJ5cl3elr
hJ4RYJHFFTEbpVcJuEcZQYd9Odibcv7Y10fszYHLvIA0goSuLCUP/VL3KD17CZoT
2KgTh0zoxdDj+zaMYgzP9wQ4Z2Nu6LApgv1rvy9s3KIiF1T1CWILGhUnY1DSBKV3
lkKyRDGb+iLxfLx9HKtPPILG3L6Ib1XVSm0E8+TLXI4yRFc7Sa2uhK8ntJqVPAeU
qOT+KNQ50CrCvJMA+G1FXv+KZhZ1Rl25WSTqre2/XSiaokcgoZgiMKGUMPVdQ6n3
7lLNjayJlBUfStdKQW8zOxwKSZHcJEJNyb243eNX7GqUzO7FZFdy9gEpNqI4wIaq
102m3hBDJbBn5Kd2WY6GMkIyN0bTSKR5uZ4liUllWCTRUMlfaGFYMZfrMiRsBlbB
7JMUlLE4+scsvKg+LSaaYIIPmtjuiQg+S60ga9zHu+FRk/odtHVh8dLmWexzpou8
Do4mF6wir8rlb4vwjL/5/FPMF9dkQBep0GkXlMOKP/I+hiM/DCVhPV7pJuFtXjST
/JrMZWGhopbMmkbnX9SiBiqn7LofvxXEIF1CwSBQIVA01Sm3l0AWNKpQoZ+Zahyd
0ucDGmD3csM7Ud+c2GeM2UEJfeI/BvY2KVPONDTLT0z9G1HKGBGfAVYq2aClgZX2
IqvRJok9ox1m6/clquhtxcW0FOKtrdydSDLDyFbtDNwMT4R0pgnUZ/8VJDc3wFDM
ATPZRiLWiYOHxqL9zxSm2TfHfOgJQdftdeAfEUaKYnQysTLJNg6N0yrZbbFMQMQq
RVgerQgFkxh1vf01PqvS260m3WRVxDpuND1alCvlPBLxiHSXP6ElP5x8149JmxCx
zhwmQA2S/zXkTl3r+XFxo1A9gxyrjEdvHpBqW0hh8WrgFJHAv91KpjWG1gfc9e3q
vpfhl7CMhCeM3xwRGu72vD5fV0KIF1hC+jX3o44MsfbbMwexT4XNEZ6tMltEEK0t
uwlUarMgFrGlu2t1XN1VU0kwOoLWV0q/2TFVcsOSF831B3CqIoq5CjC3NZGnQiY8
4LMNMf2TzmXFqSh9KS2iXSOMRtXZEc+WXPkfvmUXDQb2RnbagH0EdOli1cnwTtwy
J+W8t5rMOwxk7/wRgKTCA5NtJ9VBLTQvzAWcxlEkwdvlyrvyjLlv+7Onxfmv4j3Y
iv6ffTh7LRpTmNxJCj6+A0REPCHR8t/92yyLZYe6sW3JuvklidNnEwI80TOcggKa
EZbbdSp4oSvBYbu5YkF7TXby6OOU/KAr3aaBJOolF+7z9S/P04aviAlGJRpoPuCF
f/8yo8HTtxQxWag330KIToToueicqJaeVHRQcaSiASCfo6+Q13JhQyeNIzHh07T+
aRytvAntXuuo7XLV89TPHnQrgOdlywdpl4REWSQH4UzTTwHIM5faipCtyvkWFdgk
x76GrsjDbDaz8AtuLDWaU2DeV3dshJ9/Mdd98Ok4xXw7IynKybnCKSrkjWq+8H8h
y834D3hBzB/IjDrUpZI664Hv2StPd8TSvtqoOfwB+CtCy5MahFwdOlkjtotDf/H4
QiuT9dBrxPUJUi+KQb6zxEsslc2GzISdLl2yw/JJ9H96vm0YWgraOLDDnScxaZl8
izuU6rkYsjvYGZfiVEQSCgWiGezKj1HjLzq4I8Fv9l0vR82LuCAcwLU0AonA0gj6
qoZ6dLL0tpDTZQwZPl8dQVkVWc2JzmmG03MpO1i6p1TUBiztB2hzK2mArC/iq5IO
Byt2LfnS6HkRukLMEQn0Kv0jmJaBDJIqTmNYaPEsDp7QcZLU+26+qsSKfmkoJQJm
v8Oxqm41KfYSOdNfLRBZU3LzZrneSWjLo7h0l4oqoQBY6Md6vjlbwI6z2g8NRLRJ
AyyCfZWkPfT8+dAEy2sMHYCxooxyCerLOg2JOTd/R42RDWWLUpRKcdesEREtVHV8
bQtfWdyc3nPL9nNcM8yW873NQTonqdEaKUZKbRWh7dOnDGjyVIPPBICvKN2Fc0v2
71zTd2xl9A0Q2IKR5nCQa+xYe+8L5dxJ/iHn8pJr6Sk7bnaBvn5+GFgPxh8GpOOx
71sPhYUFSU0+VQrInj/nG2jjiWC7FYUad8vyP3f3UTGA3l9Tdw3PFw1uigt9FoOO
iFl28aLMucgNnQ8f5nwUzrJuNIVauGm0/BOG3zSiD4vVQXjkiaVY3QxRxB8sziyE
hLqI4PRS1LCgfngHVtZxiKk9gSslapE1+/t7aTWuCYBzu8AMBetcNQ9VmrORJK0/
9LseBRz9KFI370gbReAPhZZ1VpIsG5rxK/MiATriP2obzaF1EZcCisHl6+yFFu8V
RlkMWJapbt2UTFd9T7PTyMN0gr5hpW/ZsFpYY2wxJd/W5ewYGsKc2jpL68gm0FaM
G5cAYUwzBwp9Ns/75Kh7nxohDVphNewWWoQni5dAEEpLpF64RoKbvdPp5v4Bq080
0AE46yqyJcyJD9ha2i7Ta/YHE1yxtkAGTiXYhx88D/pN1hp1DUNdeVrgIwVcvj5a
BzT6YrboN7rPslGUaJrgnOPIamweWO2CXIDwZ5PPKKOy4WSBjiBMnYHr3R2dEeng
vH7AcY+HSdQAZBwBzn6r60mGe49NhyfcmAcXbxQ7/wjMHdGdHYdSEucJ65z5qcBJ
cBunO6J9YiKNSGHsFsVlu5lJFzxtlEhHhEghNcs89/xJnW8fog/JrDQAIB/VJstF
y5x2c7/5qRz5EHqV5Y6h8Cg1OaMQkTqIb3FmeqPo4p8+1S930wxVpKydLHGktzRJ
ttslLMVX63xvZMGNvhFPTPKNgtuNtnPmc4HE9i8lkPOhFBkdq3ElN+AFR7g2szWl
b2drF7vW7FVOibFYcgr0OH+eL+m47/JNOQd3wunqmJPBfa5q17SNni0TaBfoC3yn
CdbT2V6dLULaPnmE/ADgcZWCIZ2EbAtiEl3z8gaJy9aveydccDBNlTGSrXrH1BtF
ns0u5qlz/zftdYo+nHnOtqvaeii7FJ47DnRhWdLzvYM2FOX8X6FEpJu8znorQ9hm
1q3fbpImWRx2jnd9EIjrDqaxPAXFKgZIp0kl/zQuXdxG2qrr8IvLgGSybkHbE1w3
hZwEMWpXkvgSVTgOFU3FUxKlR5qFuolgF56L6aKGUCv2xt4UmXomVpLzABiqiIdU
Sg/EcrblfK7utm32VteBjl3ttJ96jtQ6a2JHLvfie2HveQirxzv7SZU/0KQJgMdD
0awOz3pST1MrgWJ66UfCNzQa4gclrK5anXFe34dpV6sVnzHsaHfNbXsLNGg7hNyf
TuybCb/DGr1azxNetNRhJG7QLB3C9AZ0DdHRGIGbUJO79vARhng81lrvMgf7RhIj
mPDMvqQjh6PjRLzItppHDB03/oN7u+O1sNzDQRshg/NwKLnVSvRVaWNxqRxVGfvH
4x78yfdpIVL7JH+qtDV5uTuyXkNngJUUWH1NRFMTC5pg0qe797FBfa0QJ+t4jX6d
BDHkksmXfP/Ut9bBMX5MHI+A6wy6YjjlZKtiCj/Qrtl4yf2LjnJcgunFHYrdYuBq
shlKWpG6XdySBbLYRgyICXYpH/HKHYga4UMEF8SFJGxMIELNHVuCEJ5pfWP9aYQy
5KbanEDOeYzxmtGeB+0aVVBiQkmnKsIRETlbspp6mYfSwtgDrHL+EWc6s04M1Ot4
7Efj8kYlQZtcpc34pApLuFY5ZOazT63G/KMR5UNSrJjpJeUNsLM3Vn+9jukAHDx9
arSJt/bLzTUsfg4Lwd9l/LEN9EwtpoyOVnAyLd7tvcZrq1iMj1vOHwi0102K6538
BKSRZS2W8Shymp8jYf+pRpIL7aQY4oUQhuipnc0EpqBO8H5eZ/UOA1bJlIh6sB+D
foKsB7IN9UyxZ2t/fEt+0hEHPxs8Cm5ogcb3es4yrGjEpqDIsYDHGwHCk5vaJPap
RV/Y7fcjw8niKk7lq6TTbOhM9flV7Ah8B0/5IA6BkFa6GhEpkRVqWIdc7bW9jB0l
JRKO0yMT7qZOyWe/k3U9G4MYoqDEsy/aOi7OaMfkpdq7WGCpBPr7SLw1T+MrLJLQ
ka/GMisLDPQWIf2lOWbJ+WQl+1vq0uhc55IFDIN2NcMwFHLAs8z+ILefWFX32ing
5O5zyGD8cRpSc27USEmxEQAkABWW3eOREO608Cwo7SaLX9pxLz6zwnLD1EdZoNDx
UzLAgW77s3YjIyJmVCej7FiXuYDFm+tAPdIKmaS9U+NptfuTeUg+mbMGuIwUa+3f
Ac0s2IAPEIVSnUADDxnle2TzYYj2AEBAPAMYb+p5cVv6AJKu2jeo5MpbGB3B27e6
anuw2pmZjuFVKwd//xrk60p3e0h+PoMNy8UjnrXgZFEgefFwj60Y42aZZIVv4L1t
6EQuGNIcqa1Xt147AtodRTYTJHm6NElKQ/84Q3tvO4z0B5/pnZz7PSYrQ84cvqoD
enPoSjnXc4FtQJ2vUY/hPsippReDTCJFe9D0B1SUJDinDEFGWJPkJO6or1BA3Yhy
ruwCmyi9xprkBs9/Siw6wyruEetrUPZSlIW0i0D1lZSxyv8U+PE31L8DKh9QNZMN
eJ5THjoPKHdNTLOo5UjHZUTYX9f3yCtl8Nb3AEKXxUkcsZ9k9CQ4z79UIPLITpL1
JRewjASeyItab2gPnme1Cz55d3MIblw3dgv6NU3HdzS4E/C4nprOsZKt+kH4hR/D
EMkvsQkE6IteVRDyX7xHD/Kg9Jp/C+aQhGNWowW+5WqmuWvjXV0m0G51dlmYwa5m
4iNallEsZqs71hIEHZMUaUAiD/CLRm4dDfbAFRDvA2tigB12zdKFEQtK+sQrnT++
MXgiFYL2zR/xea2uRyHw0DQ7/i7EmgVuDLAKrj5U6qCwd9d1/JdSkEZMKQApzdWH
z09aEJVcJ5hwd0SV4DtWAufAMuPCcXgpvQ7ILg0bdKBdVTgKzXTUrnMRwx1jhN/q
yPKp85IVwiTL/6UVpGMaE0pZebv1u/tUyuE1W5pN0q817B577nCooB0YxyLEw4bG
OD3fqvKqbRCzZtOMvJSne+f156cTLB+Hu9kIc8IBZ0QApgF9FDk9hDYm/Rl4cH+x
UbhWitGZkc1BN0CnuNkB70mF/vsOK0fxfFaK2AQRQFd8yNQavWtcMfqvD0eO/mOg
3ElCyo9tXkKUOXnJqS5ESqyZ6APDMBNJSEdWuT2Jb/1T+X8v9mj7rwT5q7raDu/b
z2EQmDX03D4CZZWN4LWgNQUEgbjmqFW0UGAI4soLkCqF5V4RaK7c0/ijcTmPK9g7
z4lRXSvgfDYbQKdDYjatJDTQCsQeD3XGA2PahcC/X/n6mNepVzPPyAefgHa461Bx
c4LaprYrRYiHFsGm/HGxNxFPY/Xw1o3hDnm3dTxuejPGdJhMkiOOYHaspBeV7gK7
DiaIFEHoAqmLZrNTYgwdppSn7EB18VOx45fzc1ENOcT2z+IZ9oOdbOnzsQrTs7W1
zQ2iWz2RyUmOZgmak/GjzkUdqQ/ZNDcchz6qvCT1q9MrOIDq0Aqe0ns+HZYZWA9A
glEDJXw4B63F+FvM6IsvLmKHCIGDQ0LtLlIW6ZQUOxtVjnPB+BD1hbgoCiHTpwUB
RUiyTrU+suu5HJ/OoFu3hA7MtczcDRpIeiL5NioYExhj1Q0dILKiun4IdpAigS+P
Xz88IBR0npkeC/6sj4YwnaucuPEH2s+lLnghxmcKQDd1YxoZKCfDVjy/LlepsPxB
w8hCwC5bsAXnyClPn+s3ea2aMsiRF575uI/Y0hqRPX9s4mISKdEKfsQTcqAfFcLW
j5oN3ItBbi+vTWBM1c0djQxsNsmOgoLbTszR5E96ObD+bPAOZxAKr5fgzWxaJejt
r87F9w7burAtqD2VlEMWixpwz4tz4LGSCUDJVPHWBwgYGo6G9XOSK7jRhHtvXP2R
RP5LWu+C2LB5rYZT8QngJcfbyMvdXWadrmBfzxptUz/B59S9f64XshHn6lozrrUN
z4dEp9V/wxhblpdQBY2pz5/rGICLQcOQSeWNiycUpn2vUHKKGykSUXnoylH3J/s7
gbXfBGy0HCOfrfamBXYzxTuo4wXh2p1r5nnpvRIzkUH4Hb2+areJt+zyQLJ2cqt6
WjR7aWC6FF1jcnSKXlVigBkC8ErvFVcf81eyCRJK5e3pkGEK0JwUjmWJuDNg0z1Y
bIwYpv4A2pIfm/R2YRgc5ZmGFlxvwibiMFRcNIhc1wKx360/zyM1z1+5Z92Rbuz3
rrH1XnASyiklTbYVLIR4daJAB1ioiX0h5sPnwgyLCPrCHAIPvy7BQlY2PJiO8XZr
HAGAtlbj1uLprQXrdhDiEbPLoRqO/ZdbP2tY6EF5m24VIZNtqJ/kiaUj5972Zm8T
A2Hzd3TCGHr8b5L3Pt5ifJfxErhqkeRuJuFU28/zGwC5DpqZ92li2dQZyGBcpwDr
uhHDhzshKIs9SXIngOI12bhUJLlTTcbN7gE2wd8jaXXymgAsEDSs4Q3bL6X9boUl
aOoe/JLUENUzXKynH5WfQuZhY+TRJ62q9CCK8W9PSF0sR0hORkhTmalhmnqvsinh
7MWZYf+SDjdNj1g1jDOCDt0Ks6xWIfbxGbtlrj01nypw23Hn/llOtTdwTvi4fAL7
VmP+Vl5nRJLwYnhecIDbKmqe0dOJkZrB3b74Kc5zL/YXA8wx7brw/iAccfEzvFBG
oO4EzeaQkJtm/iDUFqi04MDDRNGO+9VrlWwwUkrgUxubTiWcEiGjWq2oe/dog67o
tNVZpVskLb8XTYDZWkzvFyZgCdVE8FhuS9oTdnCGLUi27l3sk2+LV2eVILKEAULI
3gttnFZWqiO5GpykNdOmfC9JpvI8igTgDC4yxE+UkExus5y9j5ED7umtH6khLQqy
bt2rT+5PdsJmKWgjS2G2NWdfM7Q3mVTnQqsy1zNJ6zcpIYP+6o0aOxnt5if1Yhee
Bt+LpjiWBrZefibSc3jIZ7+eZUQUUi2P1yYm5YHUp41uPnLp/r6w1MSR3i5QEBVA
MLEoFcDvPqPRKAAowC7Rl3RUE1TDqzFyjjXWkentOwZN31NFOqB2ilOUZpF3QLZ0
M+lCJEKp24HEH65ybtXm4igvE5oAcAMMNGSGKwPwp5fayUItvWDmsMO7Nw/uVPvj
8Zpt+TaAaf9zI0KWxjx6mbI3GmJa0SySJpQT0U1mToGUqMRbMr+V0U4hCxiStEHr
byruQ1KIp8f2i/897sZCvkYAOhDN1GD7QYcTGYbhRntbrPZlko2nuV0brj4Dqxsc
YtM6wk3356DB6dpuWlIrvRJxmWfnM3VQD0ofpE3aRNDeSNmzvbLSx2sovdQHiJaU
FUQIPm4cy7jwKttLgiNEaklXQjRcYBggi4W8JXVOgIxsC97n5DJN3ZK/nrhUe4Cn
dmYIzJwsw5mNL5WSplah+ZVsUw0RaljH8UeWVJ+cQbGnwcZCHKcK8FtDIhn5Mb3G
1fYiByHTkrOR0wtAia3YoiepOZGi0WY6owbWLEpyQEX3uWbCRrBxk8syP/+nMlIV
xJtOZxTOJkVvEhJSNtcoVJRDzawWQgLxaSZhEj1axiZEQrIRdWt0LVUM5m0C57dm
rVZ1niixmlZQkqOaAdlfQrMljUmTV7ilCq/wbfsWRgpetWuX6Mi4KIDBcbWYqwdm
86TR681IqXTMy0sdp/HWnOIsvzIGqA8bH/i50i6NN1FJkDsoF5PH3mHW3O8qoATE
/gK4IeXFzrXMBrDfV0q6WQoT1gKpjfXjXq9Cq72OZ/4HMnwjqO9lCtCZwquOxo2V
UjYI2+NijX8GUA84MFebqBNOqVd2U26XyhwU+RRi+K14jipw4MHk6FzGvGOfzwAJ
LhNrZgm7OfGbYFodVvgQqd8BL6pDYeiUjvXZgmlXyYiyRafGlYOtJKBFPY82zgdC
/K7vx8XodIW+JsxHg0/Enbd1j3mJixxWa3fBx/uuyB/2nHyEkZzlFWmgFDVuuw0W
mWoFtQ14LodhZkGCQ+FwYI6eIrGzdgNSqAWb9RzVvQXzR0ekGv3Z8VeYZsxyd7I4
TM3U3OOl5mSi9eXkOPW5SxD85Og6Hehig705WBOhq5tqsDpzxHaxj8qcXtXwWH69
tPRX7tR9hI+w8YtXahJhTUFwrILpJm4QOWCh9SIPr672IGmF1mKpH2pt5VAB+h+h
6edIgXN5vUmVvvw47MmrcSulRDZnrtzmyJ36RYYdnzuu9FNnPiC5vWvu/rfTHaNq
k6rqC7yGxrwegS2uvGZmzHE3jYxcOefPY5lex+NbWY8ZZ0mhiVpBuPzRR58w0O96
FMRhRj+on1gMvvtvAoA9HyX0wIK9Lt3szj/V2EAdJmT4pBy61KBVhJe7aoSVTahT
HyfXY7dR2clU0zIgBfdtUROSUJRAWDPs0nYcjycX2dHQodNp55ZMLhdspBl5u9KR
mq8NI0kjFLb4AzLHmV9AIqHYuluA/ZNe7IODWGWlwx7n9vvBOKUh9YdSfNbJtktS
c+xLheC9SyYNgX3Q6wXRTmsJVHabcPD3AVeGK6sInIVtZ5RfIRmm0PCJ9z2VHIsp
xX2aK45fK0mmA60/dOdTk2tfLnBQGKaucA3sNlJPRX0wN1P/JDNDqWSBzJ6BEaeL
gL+6vEZuKYYZB4jtal3AyjQfQacvKaU/E4UxyIhqm1B938TDtOhdE2w6zFUiSxLY
7kv8J9JwikOExDRYS0A8i9J69LwTMwbZWC3TQeaPQVHZOG00Ys5tCMTJdP7mDVCJ
i96UtYqoB9bsLu4RVk/SdH+J51IGQehepPW6YT8MkiD5rfwe0Dp3s9wx9r5qH3O3
MzQcFR1QO/vFubeBM72G7K/zaiQq74eQgX7nky52zLBQO1Np3g79PHvmV2xQ2NDB
6txOCAUFntgSUghsxILgYKduea9q6GvZvqk/tY2prtseYuSAmT/g70J2qiU82HCA
aznauMBtF6H8HPRGGH8/eKNKgaBNEazy5s3KGhne0h2igxqyk3uiwofsluoQl8np
71pIO+ixzSu2sKRlL3WdR7udZonyX+fVXIhj6NnUcno2/IPl9+L2/ixLF3epH2Nt
/7pilUhhraVoYBNlAli8r6VJoC5+zTOl4ZV7Sk1Q/LVhMgWQ1cNQkHUYdi9Xf74w
upY1jNYw2JdD3FR+rK+e4/g2Bc/CvEZignBNFDd0eDxStSVFV6NWICvJSyQDLLxI
dY8idjd8/HDO9ndPUNYd5Jq2gWp6Xv6PPwxuFFiNSYXUPlo1QXtofuUOmf5vQAKZ
D30n4ylmakKcUI1FX3XIk0ylfhjIQFmnLE1svt7yzEc+vrLQPV35gaV08LQ1ORoR
76SSNusJsv1bq1Wi+5RhvRKT4GdnLypkRQr0EtMQeKz4Cs6Zau4I7S9i2x2X8Dn3
FAQ2IsW5FLvxYFassCMAjqsATTP9tZh3g/wigDKZmR2TX1RMI65eB4YnW+PbPab4
Rq/zVQ8VNrEwvZtwIGJkLaVktTJslZXhsg1jZu7l4lzESLFA+l3HZItBJJuLVgJp
ImAvqfk15pZs4Kfwk4yIPv/w0cBKQ4SPWvvD+vKMaxiat5VyeAVqY0VxWM6KP4Gi
KkCs77Cw/EJu7EmI7+cPyixsBVUotMbJBnOJZAkbhFO6csV6OyY/kAjHK0UDWdrL
KrvKMdJkzOmsbxr1XGaFD9mwNlpCQgl3GTNArTi5dyzoeIdPApxhpHf7HTPaSMyl
Fw31Et2g7MZ8lu6uR6AnbYLjxIvjOkUEUyPkGj6l+mclbbQY8WlJuBKY8m1zjhp/
AG3XtAWYL3t4SNuFqRiToPoOZ8z34HMn0nfpINZYn+P3lBdz9dxEon881gzhTFHj
2sLqLjqg15AD4joxzX2Qjopc+Yw9/Z1Uj9mxy8EnfxCzH11LKA1f21qcOU7FF7sM
yJr9IvfiWSYIbMgWwf0AFXNYNpHnApLBDvSmM5r+GFU+tNYVXT6udcHCrpRZ7EBj
y2GtGT0QovsT64p82pYGB5HO8OIf1w5tn3xaWe9Z4MUJI6kksgunzu57wopKvn9e
WybzEZkSj+1dwTJNBnCPMY14gMcoHmToc9MDB3XM/jopcggUA1TSSUKusi0tdzUq
U9P6AHFDqii1n0oQCaLAA6Se9mt0th1ax3F9uLMKyLjefSKi4HdFQdxKy78jWw7v
K+EI6JW0EtvitxGYHLubb7v19ZEn/iXjMP9wUOBTeqbMQAyiYlLgC0S9s7I05l40
qzkTCz00O/v6FimeBYmI0RFTVf5hOBrq3CaIOSuWKT/E0N4DyN1ZBzP3tfge8pdm
EzTBpi4w6dylZYN1zkOoJGRPWJDM9vy4hvKtd8xfjqreLj3EkeLUnVRdS14wFaMd
GHqIBnzXRiSEQ54aCt6L5LLJKZK8kVZRvi82HD3onvVtVNzNn03O4HGioZLmGNqA
MT28/dCaD+FKESlpMOkjPCzaJLg4/nqXK+mDFl/WLkYoR72gLGFIypuZAnkXBChA
tLv1ArbYlWYKGVrHxjSeyF50LIISNMNHMO7dW6iES7tWK5HOPZkDwiGPxJ+xVNis
3EypjdVlrnKwhWvPJqBcz1uokHmCavsaf58C8Y4V//x1iisPFl4Gzer9Dwq6vWLl
nFx5dF9gDFvTnJI9s7ahvKr8hXg/39lCnhfNq36p3pbkGI3ChIpdTGhQTp41Zm2z
TRjU8poWW45kLi8I9yyeWw2mm7IL25ZVptXzYCbpwXqjr5DRJGXJVeGYWoWjaXP3
HGRWB/UV2uy4oOFdXPI+34Wuld/1FNlkztBHc8IHcDk29wkLgYLisu3P0l4EzQUk
/eqYe8mTqsCNAgT+hpLittTu7OvWwy9f8t+dyxfMUzq9O0NEqiKTohqtusAzlsWv
fem8JxMiDa/K2FniS/lHMwBqjt5t3D6d8hBV6NdSdgxuTAMx2EsYPTjJakXoGQa6
P8c5ZfTJSk+YX1CpU8M+uEYanUrklIsBaq8T/K5SxdkKZSjx5WfPVu1MCRvUqT/k
b9fN+7I4MVyla8gEW++LklYiTt3elF+Rt+vmu8Cqy+Q1IGgAC8mSSpCEMw8NjMAl
aAaOJegQPJH1bA5CXdUwoES6hzi2MFiEMlBb3wwicKu7AfWfBW2qxZxLXWjx4Nkp
WA8Kxo+5KH1UKJ5UeatnSxVcj+x5h4DXIAFbKYgYBijWaYq1aKFEU8U1R0qpJIC0
EW1x6SeFgvCmcG8pL+Q06nQm7BdZfJOUMJwKnZZRWsanofjxxiOGYGB/2uEvkIcU
GMoeUXBqY3WVD/t/Zx9s9eGUHtuR1KOK5lukaqaBt9gpPpQWEoucIWqzYJ1IXY2N
I6CTwq7RynrHwPJnsVgXmBRGQlURvvfK5S56lmUdwuwKGUSVzfSk8aasckyH6egB
AZ7IvpEde7NGnGZMrmHBV3KcEKi8Epwyn4IHoXohrLyZe5tfexyk62S+IsBOawz1
ksAnQ7VH5sT1XyOrMWJRON83f+lZNwyTq8abakoR8xn+1lctSlEhrPZD4HW6EuVh
WWU7mTKodICq66Lv6jXWOJvDEh13dAcBCqBXfOwjmyfDPiNUa1OBFY3mIkRJEMHq
XmGgjg3gy/5cvoNsU3ZSOtiWzNSuK6HGuMZree+nzxMabJ33vxEQLzVVhaXUsve2
YnzRNhs5DWg2klfWIoL0DlAuZWkRIhCi1wPIgUMvcg+g/klKucvcF7Ouv2+wfdmc
lnOJl2zu4p0V19V/r4+KNG0MRCpJQfLdzqJNmaO8acq8nSpv4z0DlkSP+0f+88lZ
24/PlbN3zGljfB+gD6yQx6YgpiFqSbnHmrVYClRnkAaD2b1Ky3cFyLgT0WJ52fgz
o39/secLya7SfAJdiLqnDMVqfUGeXP0YZfzPJjydcGlgnnpu+56wVyGmWH10fIZF
Eq6b2BSl5qsNyQw81bD2zkQPVDRoG6+yynsIr6QpiLqnwNB2hKpBKt27+X2Znf6R
OB3J4bHDFpiBq3c0xFngPc7RfeSzHpz0cfddxqD3pIad378wlzD6RRbIPC+ah2xU
0P9dMTzJpemx0dkdagOPF6vtLE1kNxbZfzT2cU4nqfEW8RiG0PtzRIMZ+aeYG2fO
gxW/6OJZYd0izyWCye81BI9n/grutgWKWAxLmSEi95ai2R+vmAcvJDblguzBy0nS
8+ASEVztAZjZytb/Vub1EpEG/rhl2/N1GaYqucocMRG5LMW7BFIidwr8xPGXec2P
NxbGKeZDv88l9RLktpZYlIDk31KGr5m7u9z8SQ6cZwnmrlPnZk4VZRbhLFzNhXvB
15bt3zPJSh2eO/C/mmxgFzIWAGxOn1RBpaTNArUIt+5hd7nh6sE3niKa8rNXgk1X
Tsj20KyZR4CH/DSXUBxl2qif9HYsS+N3DHNf1H5koyN7mbbScn9vL6QcpsHgkSiC
LLUSe2yV3X75AgE7CFm1yIFIHcBnPRsTvthdRx603hQGI+leKGkSZsoc8RelXypB
5f27cM0P5b46mSMAnvRlcPaHRzqqYcuDkiCgFeQN8b4qYIrl0d1F7HUmbikHLHlD
Cm2V+B63O3PjFP58yW8FqGGw8tKo77P5gHM3FVhWKvWQQKy6va87A4rCI6nFPdjk
lHor+HaNbiCBBlYW40qfTlsLntjdzJsTFjfBWcUhKsylJG6sQ6AVQbec7Qvz0USd
Nv2aaphEOBMm6LQHhd+acWH49jcwEhqX2pTQD895VN1KYLCw2vErFDO7w9X4azRR
qkWoV8ErqGJe4eyCvfZ3ZUhlBbgMWf3tTO8Q+diAZQpKUqaLMeIymciYDey/2tAy
1EN9tZyXn9mOSV2PiY9KKX1lxXpRtqbjRLTdQUWoD6rmv3Ij5bOqlcLCkKRA5LXB
p6V7JiIvj9Of8fDH5nZnXJXIBd+mtYLVYqLCtk71XLeWlJACGJqXHawho7H+AwVS
na/rrDNE+yYFd8HZg/M2JNYceTYgLv5wTOvfp87XELYFujcPfrD1yn0jjA9RAYgv
XZi+DZax//4LIxGYynm7iBR2MSHVdlU2wzsi0tJnYFgGHb5ltl1M7P0EKJ5okKjx
pdXf7PWYbOw25gv4YPfKHMxfzpIUpOhG7ReOQwRZOQz+XJl0jKv3A1XxD6qxoMy4
tqP06ipKaUGi1W5xBB+VypJgS3qOXhXFvTGYVouEulzwtp/CXZ/I1ZjjHroBbXS7
0bBqDgeCzUXkZrqn8EuoITG7cmHA9pRgVFvFU2NC4qPKXjkcDy+qq7jGR/oQ1rul
f/dYn2aoKrz0VKj5UNPAqchvm3No7DrLmqAS3wCRjkoAqJCXlEUjBOS68R2aI7Eo
Rhpv55X0kR1a8F6sUTT/Oioz6/v6bF8KR3wN/+flFqh9+cENLcFWmFnUSQ2VeL0k
ZUz+r3qz5s3XKfnFAeBLfZJVl6wO/baam9j0obGnXR6M0wWchSPM+ufkFdITTa7z
X9Zu/zB9VlgsVEZMfNqr0CuAOHew+WLusb+cgi4+ViwVv6AXwNwX0m8pvTWMD2Vj
l5ws+dYKXouIPBUp1wDViOcyiSPqK/LUtOjRwsBcRxLomIpjw3cq69Ec/L44RaaC
bCiGt5a25TOu/nTc86amEHIsgnA+qgMNS8ceDXE6/qA356l1Sh2MVSC+1xBjT1j3
TyYu62GEh+KZj2Lzu/V/IJweCSU21YD588B/gq+/MNCoSBYOhHbZfzb8LVTClZ04
wKH34Nb1665doeHOBNMjL0aKWZdhP0rPBWHJfVZ7z/uVK0+eEtNTZso/Xhnw7knq
70Vlvt2gs2/ksso2sdEQBmEtFpKljAXMTiV0TheRahb5V9pZLM6c9P0R6Vzh11Wa
DWUCplHNGs0rbn6BSSu8ipP0KlKd4+8AxVKuCRoFkUr5uDwPqSiJG8ilZ323AUNE
6/3VmlmZO0YzJ2BuptCIiAQ0gxcO3tFdqlCK8UzfMg62zJ8QEx7JbdaibjFOCc6B
FtqNhQ4IOY1BTnSw1NPYprRlsa3A0zHBctRtblMyi/HTyJASLmZp8UFUbDVKE7Ug
VJ8JNNb6EUt4VmUKXr3f49zm2s3/SEJGuzP1qK50LcLYN2QJcKfkkJdRkGEK1NiY
Efz4Snu+84MRDdM6Be+LvAwKpCi6OXc0NF5Abfl8WSqKNuPqszAPZjlfK9A7aKjo
t2MVNkYGiQ6O04GsRUF2Q3x+QLazjWJePQbfJ+5IoLM4Cj1+ZH5L9QDm0McASkk0
MiBAxxDGP/ZJMOrl/lZiGok2gNL081DqNQNjtM4VPknxD0wOVYIVNj+lJXvjyUDh
OdmoTWHgeCh3iPFwObectO4CIRoOhvJxsJhCNw+5Ep9EXThuKD5U1XuRfzkcoI29
sLRAMmRhFltQSstqEVU9OPjx1KUEi+AzBOg4F6lryz573KZgxooFGpJi+LfFGYPs
dwu9vbpkZTPZ6TaTX+Xguwx3dzx+2U2HJoeVY9iLePXMnsQWuqE2ECjhYygxEBNg
9O9+P0pDBG2+c3bc3JswTwcjrWdvGwzq/eiSbssxXncpgsle45wcf4RURs+Zw0Lq
sKwbzn3pcVQ3dS5AFq4LY0Wct5eZcZgOlvdoONdppDr0dzFUknCQ/g6MlnP6Uxwg
AAjG5YhzEsCeWUk6fkyytJJv3dxnDJpXYNcbQJb0Ldjp3fPsBSHGsVjGeVjMDEjq
W+3HT79e42mg6K0NKmVfqx1O7soUx4Lz+3lWZE2Ad7Bn+Cis76+IEJcgM5VHEHHd
QIoHQ7hmgI7LToIC56jRuI37ZnWC9z7aCwX3ph3zgQtV34QEmdG5W+LqB4CNRpEK
p1iCmxg8WFmazZyS9uGdLEqhzu60vypFbWiEavR9bdmhVb8mJgwox9KwjHmg/lj5
+DHXxWJfVKZEY0igHH0Rtjf9E6yMYru7ebze5Bu2N5zKjlBjh1/TXxTKFmj7VZow
EEgJqULub88jW27CPs1q/9RdPanWGiIHPneSpID+9MF/rUUT9pj6kBD7Uz58LSnu
madW5Rof7IzIpwupaEzzVN+jSMIiMBUHH3IQwh6DV/K+qRmDvQoj5XFBLg13Yk6B
qeGeQU0hzJRRwIkLz+EsQ3Ul+Bko8poJ6D+Xhw9+6fdhpkWj8+JlVyYNLmuzaqpq
0Ik5uNdUBxqHlU0hZTVGeypsIsDBqlysW1xHv+fIzQ7JgwMny02UsX/0N9uFzCGL
/5IOMuOvQGxr//K/puQOAKdHCIEPn2fNbg44ITbP83sEreRXV+UozPy0ZUS5a0fG
hvUC7S6cT/xB9l0VvfMCrAmt1rkoHlhizBMdCN48WSak77/oHDnPULnKcw7Sf1Zc
OCQw3EpeKrBTTxzNOEhDNdTGV54NZg+EbvkwIyYCaTfxBtRr/pKEMRu/GFSz9AkH
N5qB8ey0crwweL/b2yMJlXScuplNz8K1AM7K8GSQ0uAYbRkLTYsyupqY06nz7/zp
YOQRRUNoAE1FD++7nm2KC8RbbwZiWhmCxG7ltkjlqi7Z0+v3jE8s2TBf+u9PphL4
Om5F+phG1c+hfGGDIBlKcQ6ikkpXeguxxaQBre9x4PEANCMgkY7fYyCzm1/zLXZK
izwwYTJeCMUZNqHJe7C7JyP6vUEB12UY/kjKYhQl+xMrvNVclN97YesUQEOXNGdk
MZEdkJ+/28UQXTQgyA5Qu81c8LkQY+p2BGUt/yuMGjq1jHS03QjENjvj3+2gcfyR
92byIGWAhcb0beCDuDgj5s9XFnTVkzytRmsF4hpmrZgw8Ca8L7P9Y8tfvcjJ0ufL
eFriRgap3Ysk0Qp6fxAaXr9uEQHTMKY5EDCUy7d8wWyIqJBS3gd3a1OJtQg5jEOr
LNyLkvQRhhEkIFDekPfFAtwT6FRgxzFHJrT6i7N0lbwGOcGi0Qo2L3/Wg+IicdJz
SCGLeHBZJbkClUnb9MfELVeh3bmkaEhbh6+dfekQUsVuapxB0bdULBk9tJF+E5wm
Xw0LI33Bz3DdU9LaVCNxVEpVHW/FXEm9gRVxbNWRXBSADQZ2HgcUQdN5dae8zNIc
i/n7l5LsJhiHYBMbaJEGzZKfeZ8ioQnb0KXJCiMoWLYJap+nShVDCj2SbriKVKnk
wzLjqJhzs2e+ihjIa8HX2ZTLVDqK1rnpd8VHRBssnHjk0OaLvm4EoggILvyZ0Kbg
6HT/GkJKSzWkXXQ1clUvDwGv4UZR4cmb9U5CdQcyzaxOeiCg0zbBJYux94lnO2kg
8r0qg0tGY4VkqCPgoEN4rf1T8pHSs77rZDgVjVn195zNj3Z7cHWYIVtsvEScpErt
fkukyT0pVxl5XFZWndwolWLHrDBrX6Xm8GPbPlTVAPDoQdz9GvZ826hmZn8c/cA6
pogDf7k+6cFyR9UnDy1fIOephSMTU6Bj7GsNRshN4mQJTIEct36DtcmIMbjpdB+e
oWU09LB+rKRPnqYoPPXmrjVUXsr3D1g/Hq1pQ9pBHkpkyV5Qh1V/tZp5TUY0ufQw
Fzix9e69rwUynjVCLB9j1yL0vCrNnFeD+KR+XHCWq3aYPPlY9xQjA0odOyTy/11Y
j1lEDNAHrHet1lWoZy4WLAYyVd52glBz8gzYPIvWrcKIqd1+IPr+9qOEqaRYoUZx
8FAqr3gdEimhiRJztYVZMr0Ujo3YaLV7jxJJu/vlm0chYNBObx1lHyquOpNGTJwL
+WLCrLb2p+C16OgM8RSeNZCwRJSFv/WsAu4UwPeDIYKOsPUVmhPDPOolBWvIs05Z
b8gL2OOPTsryQd81WFA/GfgL9bFXqD48ARPhJXDZLwGq3BUS5yBBFFkQXV8R2WDF
6oQJUyZ6t7/1KIyvZuGFVshsA3+NZKX+l8iPi2TtSesZedjKnTpsL1lAlfd7fEec
GkWmZzLC/c4lWCSyzHqP2Qkw7N+9GVicsGnzg411jCuqSqmDImtJFdzY3NPk1Amj
SkggWfNqCdkGktzbErMA/PmzC6cLTKiN68FHnXL7ZCgX5Q9ZQgP6EG7P/fd5fbAw
fLbeOG3vJFlKF5DFDQMnmuv4x5btZ6NkWyq3FAJvpSrH54r+/N577LzuFLpmiMay
tJO+1lISCy4ViovFL8N9UlEZ1dtKoHFu7xsZ6I52xjRbEaMtwH0Xua1avM3wWeCq
6/B3jq0DZDkRYl8P+8B0irWEh9L5l6BG1X8Kgot6+grV8oq64qGeZhKSjsyUSKeS
FK3/CakBBQEFaPq+0vi7f22Fd6XqsmsPDGFdzl76704fhkhYgpgQv59KDaqdSntb
FML5ewRpErURK+JfhQyCheXvwYVoJ9zYkzLicKSlH9nzo8YpJUaq76rdOnN4BFu2
mzxcUXlhKK6LGmmxX++4VbPef7HRuDbIDOmPwi7u9AquYQcQgNfZm4eKLjmnJFvb
qCLM6pIMbSGa0XEU17SqtvE3Bxs5xWL3GQ0a4dKnJ49K/NCD4jfcXH2+sPCSNRxk
eN8wXEf5EVDdJaW88a/otp/tN/O8uw6eBIBFQUKfXAF1Hw/BHT2CpwRkZXZnnmJB
6/nOPaQI+PRiKYDbs2qFqRIGg6KlDrNgxKwu9etW1nDLRQgG9HyRMstnlVInNQts
baV3Ce1jC3Gdbx/h/0pV3JjeSeGB4DDrg8YBFDkZfxb3nVbesPSQ5uphaBN8ex3h
U6CgiwWwGHsB8dIeIL0PbzUrU1auQ3Kz+AFx1iO95Uy06X6VHI36no4f61IQANSF
ocPVY6NAQuEKnYCwVxgYC2i/AQIZfhxCDYhzquxmOSKefPh/zmLf3YohnCpFess+
P+FFb6poWdgEzOV6e9aruZKU89VJBUr03REVMbICKeS/eUfojLGE9LFu8CMzR6uu
rJjUDCv5kN+cKfIQFrcZufV4J+tX9+qNSuk7LDYzSJeSCwYIlbX9XlhMwS7Z/6lV
kFWARh+6tMRyGbqTA9zNa++FwtYLRDBJWmSXDDkKov1pHN6Q2CQPfo7+RTGknQE1
d/12GnYkwS1s2J/40rf8laqRyEEaCfH99bqpwpS1khvTtVM12iSvS3s9wSeR1PpP
e9hBZ/YCqmk+u2x3TqXtYoz3HX+ptAwG7MIKjgSAldISFhivaJOHVF4BGbaQsXL1
PLT5e2zq7jHiiU/twIYWoPe2TCf2rcWva6jFPdOM0nIWs/3LGdfW2x/T/edTeFSX
VTkqC+te9ALa8bZ+Syms9/t3HBdAsVHkLPHgcWvLyNSNn5okJPba0EU+IxCH5bUH
git8bxaV5CAKikeOEZJVztIdrUroR6/ovYyC8zf090tF30NGHCW1Smt2TTeGqQAM
W6eXiJiENorDy/s71g3n42RGK1wuzy3XvsKLrmgrQudom+0ukw561vhlJTVD5AJB
2cxGZiwrdJxx2X/xLO/L3Bm9v+HOnxyxmtXwJGNaK0DHUy0N8BO82ZbHW7z4XpCV
Sp2qZPUUFjwkjLNPjDmvqD207R/2Vbm1gMeZ4gBXQpbWRQvWABR3FyQF50l5BqAT
nWv46G4CTMWo8d4FJN5PFJDYeK5/I3G/oVmWyFeRfdF2shWHTkBx30fVcENtFSbM
PTxyJwUrg7V6fFUFZIn3z/eymVLbf13tDsnWt8nupUFEjqHrewWl6//GRekDrjth
3LOf0tf5W7SiIJ1UwD2lxt4KTCz2HHDPsYD03HmCdlex04xT0Nx8ypSqPURGnxpo
0V7I9IBc1suvyejPq04j9L6NNBltmWPzCah4QHarGZWB5+SnwgcSTv6AQ/XmWaLw
rZQkL51ZqA8hx4+9SMeYKCZIN7L5Yopz/4pcJbixTMflrjkIzSn9AWH0urC4eHZO
aUZDwVPCRrebTxpHm/9Iu72jJNAb6w/VesMohxEfxM0BwvbwP59xXMiokIvUX342
9xKPkngcx8Lz2+fGtlfqrCWX1Hj5qrtgmZXFblQVNmKwd73AoWVKlmhGD58uc8iO
RCPWI+elqQq59KO3nF7VkuQ2xMoEZJEvqFlVXf5QRP0s1+xuZ0AxeOcp//bTaJiQ
ji9TmX0+Xge5zwzZ/IXD0+N5VIMS1PTXSjbq9757D/WK4U06u/tWaQHYI9fCEn2E
mgRivfdDgWYkogHZBpEwYkGKFIpJge1Ey3sOE+pR/EM31usDb9zvZEEMBhEPYGtq
Bmumx/m9N6H2GDgTJLotUbPJBjbNHafcsi94OY1vBYJXLZpwArgef5ZfOZkLLdL6
YvtZR0v+b2OZM5tygD6a4c47BdTDi9l152AYeH/A1WNpAE0+y+9NZFRxn4wP1F7l
ZpgMtkqT7Gww5/4ngMIbGZPlruYPfv0iKYSfsHRweExf99o7BbunjcHji66PTQpq
k7XH5CiHnHyFdgAi18YRmBLqEHDMgvH9ysV7TmDOESrfuZeBerV8d8KvQ6Tm2wmg
xyxRyHW6CeXlToIEl1redGFyxcYpF+hD8rjOf49kP7FMlUqOD/SSKhWNFCTKc3OX
+4rrKhNarYrLskGhHV7VJSzDWqmlmUrmX1S8LfyfaKB30RuVy3e4RJrFBfBdGnLU
45bpbTFbz5YEz0PsewsSV3DPnHrNagKhX8pFK5um1MYsQU3PXjwmLNdc5bKRpOaK
C8MhPxnnRSSm/VEqq+pQrFihUrIyYBn0YK8fQEXexG/HQtCGho9AvBYBpDMGmIi7
u4kl6IkwzHWVjeFobKRyNZvRTGV46PwVq1AeTSOYhcZogl+YwkuVhgGi1J1GIV3f
z7Dn98VXBswd9KiCwqxYsrpVTsFdPRDLykAIqDoiPRb/FtVM0erwNdPzgTR1jBtY
hYGrZ++GDPWPMP7PhunY06Xkf4WuEcmS7+5gHcGJOuN6eTSzAZFI+1iPbM9aWNyO
pFKRZ+0m6U7Sj5MoTyEImiieI8x0gKPGh8wbwX0MA4DYn5yQlw6e8HHVr2OgCnM7
y3D15O6HHW1hFgbWe1yFj5j8AgBrWeEkq5PpVkUsRXZTnom6y64w8RnoBG7HFU+j
C89K7HPDnNkSdZpMl2CU8byj4SiHLjZRQHl8MgcZ9l6zUTFRx2xRRs8fQ0aVnfUm
lULiv4KC2kCWI2C9+Pb4wD8Kq1CG8hdyCLuzhrN7bh05vOkbdDJoEBV2/CI+7v4K
e2B8+OeX5U+P1/dwewX7rZ+81KOjKCbevE1DFXMGbB/xI3AKL9TIrMgi+qrvVPHT
TmF45K1TlSJtBdbzfmSzhqgEsiLgRxCLQCV5ArWyQDch1tt3xUo0JY2ZoQVrgnrs
ZyfsbSBapYNmwUUSw5jgRZoNek2Z6mzYLtBf5ZNDR3hXbHeLUOIrj//WaO8JnQd/
jfd8SqrbpK94MUFTiy15TmFVi0mR3+A1RwXzs0EswW+To3zHV9uMOBEso+egBhpm
nn7F7aMGaiEnKs8bEgrGy9ayl4uJv+vImCA+A5nOofgAdqVWDU7LSN5iH8m5ITwF
uLMcHs7lDGQDkLbtT4JVp5pGVRKjoTN2z70UE1yHher2tRUgRTxQGBNyOjSiu4Td
cWx61leWXeKCgoLiDDCX9yAyAGMqi/Tm6lGn7G/rN8EsOnB/8CxaQCn4eUvE3EUK
lIX0CN9YW/75Z+wYQ3A+/OWxoSzP7WZcPS/cPojn5NJe952C5WxRdYulXbgwnu0P
u52XnVjWmmuHy7Z42GsRC3TAdF4eNyiK1Jdzmju7zjEEDJAvFruNKUcvXWrhkhLa
huXU27e2EMTDNuXCwi6T9i+3M5l7BaaG/TtjVd82PIl6skDa+kKAxdxxdSuAip/J
R2IZGfZ03Te0bHQUnRXz9zYOHSMbHooaG9NdY24EGby5IEqExK8xJDeGeskJj6xD
gsQl7aEca1b7DkiM7yzkiL9Vb79hve1j8EZtDsV6n2+WidiG4MwDNKOuVy5ZUJaq
wOrSK47n0xbINhcU/7i4KGDbFZfoHVq1YSia/50Ola0H1nh/kc6R5uVL7NPIN3PP
vfOA0a1J8Xc+C8zzw456bFbxAMWVDc9z7HWC/C8IfH90owlEfI+h65kZ1uYAQhtm
RI+AEJQZs+QE+Bo/qqpYMBlqNflT4w+cneZG2wwRTeje/FJezQ85gKsv4dK0pDi1
QSL53C1/zcETmtsBZ9VL8YXn/yCILjlLYDpw31boakJTlFfNcl7CrHlaImKJg74t
rkldMNehi98nV0nl9yODkPJxvMKmuxgM5nT7uHK9bCXZi1P7+qL+zUBfEKfLHBUV
bXA+h5/Sd1QD5RizYiRaKyMOFPHhh+h/Cw+FI6F1JyDuL3lgtplEpYdBXP8cmtVp
2lwUHhQ7KrjU3G0orm2Edrvqu56G3qQio+CaKbzUwQGqNgQboI2ktpsVh5N3IXvD
xfEkWh5LWTf4UPyeXB5bYO2APoGE0+CDJR1H4RZV1Fb/ZdI0JGS1gNog7xg1lT6I
eO1q32KGy+LSUojSlc01S+X2Zb1GawdMECmADyNT9FqMEk5Mh+bwB0LKE+TaHSrO
q5uWcyMIP/wT0AjUz2XfJf6U3LFvSe4FaaSTb0eCbbo/l8xhvqvKyLq5429FRMlR
yb6OJGPqTjtgtgetAA6kX4vwgNuLENeGrrOtxnFE+CzxGI5NFGzlTgcrFQHlg5js
XL80TBBUDA24wqXmXAYrO8WrBHLfm6J30yoWB6WpDYyhVu91N48L1QIKIN6OU0Nx
9O68Y6JmFJDA0KtZOXzAEcmdIlNjfoWc10hrhQv9AQ1wkrdtlA1p5qolimlIGWDn
EaV4QijxV6tfiF+roYLtcE1gndSIdaS93jnXV2YKU+bNPuL6SDezboCF1nSvrG8u
d+htAx3zRIO6VKlOqROqmYjZFJLCUNEO5KHLOWXFEicUPrIcXg1sBTMfugQUovTQ
Lh3B27P0m3yuaK9D1eJFbHkrXkRZKV5bTsuSI9hjSBMDDWePNQLD/UEY+hFM4d7a
gMJPW0cFTBB1gkN1wz/ROoeWgFb1Ns/BJtsSXInAhVdlcckI63tFDwbobni7aYpC
VRXyiuvItCdxBlQJMVoBBIH0baCtPmgWcAwu9Ccm90n+TwOIZH/TuSfsfN0Sl2SK
Lh2LtTzBYSJFUIyvjHjAM9s9Sw4o5Z3U4HgThmKvAjXusB/0tQ7QzLVSkZmKejCN
XLDiVX3Hmu+ub7nEPu5V35wkLGOIfeiayFXQKVH3Sa3uVk2BohCI3pJAzCJ4PTbt
tbz7yNWBTDInU03KNsfkE9WDDv9FzyZQ0SJ5rBD1gA7eDvSweVT5F+wsbVIvflY/
0XaSovpuCxSHlMJoPqzBpXkIgyBqmydxL+epcVV1vV30yt1+05T5rCm2JFIYmhTU
MXi8Yubovoo3Kwenp5b4AAoVkkuuAmnlsyvXuh/H4spCxWECXOdxGxSPhfE93Lai
xbYIq/ffZ2xzpz6Zfq80VywpWDUSbyFxhsYUlxMucJuQWI3Bv1telGFB3jFZ+k7O
LFTOH2mcTeKloEk7KyGBXqHv6ouItQKLmnYRoFmOOnZsxsfxb3HpL0YsuxWQ65YO
kZiFNin5fJPjlYmxaOIX8Tofrtrb0sOA+Np0OdWnAUF3pqT1+GanlmahhBiaseTs
TK+tc2HX3u36RwmhoXw9PKwz/F0mZ1pFGcneaw7YPI3zxZqm+YAFqmm2zquqV81q
tF0D82ktdH8bwQhzstuARxYcCrouGJt5RF/RWKJblMTDAAMMsuNEInIsO4PWRCiB
VqzYXQira5mSA6TncHS6NFp0Nm+vpzi5SNrB1tI4jBl33lJWH1JRy2gSY48ni5UW
/jNL7EigXHQBaBLEsTl7hpjZEhrOnXRYJv9Ycsqz/SAz5/otWgsvy2+uoNmdHT8y
N36D9IWEnaSKCSnoiqVKneocGYi7LydriKOPBS4udD08DErdisKI8fF3cMJQppAu
9VCKtUxLsyEeG9ewoNep2Tktd2fYRFxO+P9RdTRo+K1Zx+DNxva9KcUycnlyHE2a
s/an51sAqgRtAVan2nL0oqiQ4AceSuaANKW0nwZw2ImhFc535BTSM77+sw2Ck8PY
M5SUs+TFZo8hp1dFUcPOAtIL75O/9XQYZsc57sZThulvQ9dn5mwxqysh5yYpV7dt
ZCHsHS81SroltIQSs48UvHIr8jQiQDSF/RN8yCYKEXr9DkYPr1zlELzzjYGuddIl
PcQYpoukkCrER8QpPOD0cIe1qACzA1xtA4L18+m+hjVEfEVaUoWl/aHnKzCLankM
WO2CEP2ZTpbHxFsa3LQjMUIqm7IFkXTomqydpsIyR6qdhm2Scbgehhh9xYaUDsTJ
x4LRql2fOqos9wTNx8EW+4kOoaUB6cftvEcXJHv3pqyJ+ThDOhG7J0yITNPna3du
GdiLzkjQ0bq4/c3OQPcg7UPfScQOEtBtuAX/6O9Dzlvw1/9sxjtBvyW+HtqkTXYz
bPQpi4dwoDYnOBVtLGlWc1bLe7nN4dvpihaAeUEY0iuzJh+ZK/gcz6hYz0PXYCgP
1Ddl7VzEamXUmUKzbCvUhDwxb0wkS5ltEj4G2pUwM1K+3KOvt525ItU3fZUb+g64
ScXd55+s7ZBr68YG2q65en80mGJwwSKbHyyquIK/91DUhoAxhrcSft52UeOXbYuP
V9FvU+Un3epOGKtQTu1ZVCSyvdrHaSojAL/ta2kofFv3ZnqYa16Hk5shbRmm7GF5
eV78pMCEQA+Ru7SucyXX4eUCGdF6N0AP6ReZbQvkKfoFU13JmYOruScHnZ0A4wF3
G3NlHNYF8yk61N58sDV29eHJVlseIMl0dD3CJRevwkGqlIqitP1dfieOSgmsGBjc
hwiaI2q5n7d5qg4mex3jfmHLBqDs16b9eOl329Svg2+BLi8VUlLZUac1UJrC8D1/
zSLRkfDW5RytIwmsP8zQ2Vfdf4xLR40I0pxyE7vEgjdgofmYfI+mPpQKjuVTeoZ9
htz+CovjO+vi5NdCYpwrkJEuYT98HzZuckGhTN0nk1FkDESJMzLWlRp2Z2bgOSWa
dGsOWLNnqVyKs7lrb7QYIPvhbhxaVsreDPp2hBbxTT2Gp01A+3biBvNBy8gF1Gc/
mY4/o+SXPQPYi4HmC6tjvda7d0k7wIH0XN1Ne7pcrmy2P0518qFJgvgY68wDfOVQ
msLhPYY2TMqPbPkqSpNTeCfQlgTdd1jfJZ9kmL623iCLk4yYpL9Ux70vugQzCsV1
aMa9mtbMhrlyzojSvjR2+7FAlBNhurlj5sNwZIK1+Mnk92u3KwPFBhTskGBCMl1D
Qn+nW1lMhhHY9X7a6xsZIekhCQk1tKS29aVC/6Xgec/3OOolUS9GQB7rSGV2s2Cu
uphilyaE1qn7Z1Mrv9951aTDAHrtdblu6jMgT0dQ90fwKzohYbtdoPOFM0v5YAWM
KPVKh3SMU8fO2X5A2poNvf6pm/oaxvbCb8IDcjKuG/4BksBzsLv+YyYwRVC4YHlY
0qLCZTHgpeT50lxJznRDjTPvksSpC/OggGkM0S7e0CRHBdRzSNq1lzVjmDgHnteH
xsiqYfB6s4lxCBsJ5Nj09Fn1AWPE6BiCh08ylYY8hve6tr8CUFWiQAjvK486F8hJ
jopiAYw5h2b/45w5jRFX4MKWzsqdpXBhjN/yA+BPk63x/quGrfcPSHWvdIyWppag
kj0019KZBSQXK9vR433Ntq4oAMxS8htu1zWQGUAVCpr0QeBtARWS71z7EqsXMhxN
7C8djcXNUQPgLd87GyM7bxoJo8gbCkNtNcKvWoEp7P9yBwrgbRuHe0f4dEBoET/D
nTOx0sjJ/PwtLG4q3u5Xahxq5Jelc73ELHmU4tsJ1QCtKOVXg+AAvbdVqbZD8dmN
xG3sZllQE0c7Wxr3lX/D/642h93/IhnxR6oRU9qg8qIh7O290i7pHTL4qHZEdPEI
Q7ywHT626GVBgvov1iPoPn0tzgnCzev4FlYus8aGmTbRxUC3T+d4CG4uZ9ter2Be
3QVj3BuciBV2SteSJewQBRR+/b3awQSrXlJFttXtpPGaaWtn9I8lcac+cyLDCbfd
gEPlxtZtdaawbN8UA+HiKx8LGjpHS7LRyhL08lGI4lsRH5YFq8tRcqtqaxQl9ED4
zusplhrbhtElFpsnK7q2t5nVvezMr5rMH+OvP8MDf6t4Q31x1lDnGN9XrJiFLObD
3aQXhnkum3ioqSGNaukgh1KK5xHllzv8+0fE4pOqI1nHd5h30OkF1VU+oiu0EX6u
BU8X5qBUalhWSf8Q2mA2prGrzK0+O4liPurt/WpnLvYiVIXiT6/A7Z+ESVPjUP50
mBFWjPvFGM8L5hG16Gv7mu1IVv/4I7ZMd3Q3jyvGvs+8QVCDQckx9wgWzT4B/tAN
pesnBadsVolN3lgOT/hFnNmh6NovOkQQu3NvYk70q0KJkNltCcyotknOpDyEeSAd
lOeMmMOd0ggNwwX1afikfsS6eoBOxfwmtjyRlpXjiq+jJNjN7a41yDZgjCvHN89C
9BP6hMhuooav/ckMP3jbQoRDwEpsBzsJjQS5JOZ4mIWj2FaczNJEkBPUGCnF9ZrU
uC/9w96oE5vtl/i3JDzLq1s+Gm0BQBI+R5ZjZVywHI5nQqqGa0ppZGpjf54JEgf8
mnymidL9MRDfNh5yPOjI3Stk07dwpKkvzMeiTf/GYuXXUihkJ0/KvUkkVvR0TULw
Y8k/TBi/RKogtOwRDQQhFyGic7XetQibffHmx4YwzZTeIs7+FFWN0S7I0jqCH7V5
92D3F0q7VorJ9pleIBv6yl4SjhhmGSYHo0mE2oL8FM9k+QfNRNoRDdT3jdQoUoj8
MbNAJE+cfpPgpxeIc0UWSBeNZRCCgIo3sX49l4OFdDq/J0Jgyuod5CJBNkmebY6E
6dsv8Rmh/srPgeRclrdI2uk7Y5GsgY0+H7xXkzVpGNpqhibgezc/lWY6UlyCXD6Z
MSaEuDp3Q0+6T3U1GXg7M1OglKAWeVpiPSmRpzBcK5WdhymrafqruPhN5h/T/su0
h017o3TnZMMYsxCy598aSjv+dT4KwkZZ4Ud3fj5ayMixFtpNxaE8E4HEIe0T6R3p
D/pF0jmuR1W3GRwyfH6cwO3YTVWjmF2ymwcBzapwdoSfhcjmmMBX9TIPoisQzaTH
mdY2XWnvu4pYDLH0AmDm5oglLAmxxFK6c9Ml/TTXAR8fRwif0DXxTRetCxAPjmV7
b+LEZoWXT+hGRH3fhqN3WlsZGvgf8F9h7mtjT0dXNhMAlQ4/QCkBi+uxdhuS0lCD
2cU16/vmZvD1YqcuNZt/YlDRyczgh8VDI3ntFni3OSbC6RkEf8VtAb6GXK4w6iCY
Yafn6seJ0alnkySL3u0KKE8jrEyMwEtRnMOPbtMg9HMt5ag1stp0yDacPw4dmywu
uJu2c+YRuoR04pcZs5UoA3ZoCD2gC3djri+q+cyZC/LhytVpW5Ifxb2ATLE4OotW
gp5DxQ2sHO/GiGfBNy+dV3vfmBQ5h0Nm6ryNtUJhOkb95Qs3qJJwGLGVdq3Yl/Xv
x8lfPkNyzuamqJ3MoxW9RdpgFdINq6SJcLtAHNtqrAl4iSneoKzUhx43wbXxOc0v
xbXyNRTvYBE5uW+qwXSU3J78NaZz45/ozFUz874VVvChm/YcTNmJRv/OtdOxK64L
LOnHeFAVc2Git/uxIyNzogVbw6L1+Kl5d4LX3Sj00wW/IQ87edTTh0g2l2BhfJwE
IhGbmG+P3puXhD/WHMcb7H87FmrAgObNMVh9nBJjAsOkrwL4Ieo9uTnbwFOv0OfD
tBkk0uT5H4WELihICVRyk68kHuFVXDBuMSiQBoLBVZAOYKgPA+7mlLGKtRZadwQg
WbNtN3N61W/WxunoCXzc/s2X60toG9kHUsOZJ+142+r6GrSkWhwptafN7kFYhQQj
LbQvxpr7w8FlOdu0OJXr9iVVbWazsD8c5dG6dW0EX7UjahgG+Om9kg3DAjOf5hWX
hDJJ8fgqyQ5GEx+AMK5HUJPKMYkmvjBUKQwgwb7rFeNU/snGaD7gf1H+PVuRTksf
xrTR+dZw3TxAOEHlAK0HRCmwhbA0wh73fxCcihZKQiQAd/kEOPhQpTPOoqHWhofh
KxxPX1qoSjB+XajEAJzzT8I6EnJYGc8VOepnTBzVFYDYjVHp91n+m0pJyFr72Mk2
kVtoVNkSpHYQPUgLxK53VOH1lnI5bFrpHwsQb4hs57EnT1F7zvqfF9JXMOSs3DTt
aDBs9UX1wcQGoO4PTpa2zawgl7RRqNfz8zds6fBPaSxfais+vszT7VYu/7pjqFms
92L5bBPE1MgTcrQDogD6kdm0BJ9C9agyJAuwYyiOr0hZT1FaCAxnmdlTtVecK8eJ
muDy+KmNrwLC6SpIhLCf/o+adIu3P9ixDQaZbaEyo2h6pauGeYCZfMxun8UriMmw
jcKyQomr5ZVNA8SYqTGNrbYjKyDgaosH0PqkO+o+z1u2ArdgNW30BeOjFZsJc524
NeCn9yxfb4tWgzjw4g8eGF9c+Iw498HkjZnxg5g7YLELKxsNGGdj+e+Qf2e4+y1B
HhbXfCCY+ocZt1FejGD9rjzQtxrZEm4k5Bhga72pOcKqEQxSFehhaoKg/m3Nneq5
SdVF7X8ezdHUzBOSqunX+LpVxqyZlwDmUowoFWVFhal+iZ8BWHvy7MXk3PHRw8g1
UDx02EqQ/6Nhqr6qkTfZJ1wxu50dBf0ZjD8DEydJJaI1iR5zxJBPfnbV175FlKBk
TJWUlk6rvGnVt2JKyJ8RfkhXHBHfgMEW9c9wcX2K+Qgow+meJFZWJmHkqiohy+RU
Ud9C/HGW/VlFBe6H7aY5Zan2TqHOvuM8gE3WRPlukD88Auu/oqjq4Ojsjr9TtpMg
TKaomwp48dQh/RuaA125ud5GHAYOhedwCQ+HaVPaaPyLLDadLMF638kqBKmkIEuU
5Uu2pi1yTMgMQGgeiE2xkoyhoeiLbAj4Ov1tTtkbV55D5FmJS1aWQxCmuDcqZh3T
vtywuXZ/f1S4gwtfjSSx4HoGgwurW8u7hU0yvj2S/sBgSb5jCfmfgJaVwAf4Xq5t
UCEW4se2eeMHmKim4wiHqy+f7Y66xasrhfhJha7nivMbeIkdlJGSB/jTn7Skky+e
7BRMjugxBTGMilqIh+hKniIpuL27kRUPEMKS+rQQ+ZksUCEwQh36C7ZRYp/T+hBS
vth3zlJaseVhMx6fmVfXJFYdt+opli4Zi4LBPhjuMTB4/V6t0+WcJ/E7ljtXNUVG
RDHOg2f1WxiItLriDoRLDaBaXUEJ3eLsmgUFF1ABLNeb74SgUROF18p9TtOKwK+t
ShtvTbbIXjzEdYX/UzTUsqHmwIE1yZ7BWhteBtfmqNCR1LwxNIVcMcLLJuDEzUi2
CQmF5w2iJfVCtBek5GgFEB73lFawR479ow6RxSxStbXWTDEnPzNBekdPKh+7UTUC
0jFTwDUqCJnYvoym+uN3W2bOUC03O5k97xB6xj4H7bLAxVxYBf+l+gbNBVjbJ+5z
1YM41VADcLowAxx10cHAVIuXBpKDcffLMTTH/CxLnZs4oTIC06r4NNHKzzuAaGiA
xzKyM6bkD+hzQHTT+dHOmTmOPPOx1UinJ6tOoYy2CI3ihg+MTJBnEXs2vp6Zm85o
7rcsxZLT3Mue2gXU0nTL+6sQJ3d4/5ZPQYbeiM9zarrEE/GXxKZLCKkKzyo0y1Zw
lYtmwUfIChoQLphcNMrwi4zcl87hXsKTIukcFsfuPgQ92YczyLSXmNg+qyOOERQM
SswEkcRHP2iDmrBdrFiaPkyoJSveIk6FGOSiwqhluKbs3agw5LTyR6T8DYO9GynB
SWIJaDTN0nQOut50vtNSmfxPI7+pjpL5VF8WSiUA337M2+1/IYpyLS/pkKzZUP3p
SOF8PYhSDy9pGHbFSfjsHHTVT6yQJTadhbhMqvFsixBp391z1oW7sQuoJum4P1Om
Vx2j3noW5f8eObZ1iIMrvQQsDb//r000XwfFTvCl86K2gX8X0Hxn3e2AAMXYDMjO
pdiiaRlfy00CcO5QS3DEZybLeYsy4N7g3WGhDP0mpyn8azQeQ6MCXUSxOOkl762j
t6Alvf+DK3oHlvu8TcG7imRhTl7SZXJiJqqVeBtq9jO9nfCvKa7hl9kJEYKI2Ipo
s5sJrgOM+q94eb8D5RuDn/rHQGs/Y5thC74vNs1nVZcr6o/G176/f1Tx8yEktpxF
mtGdu6zAQqX29rNdJny87j1uqBDbQ+PGEQ0czQpXhFrCq1ylQ2FAIswKe6CBi+ZO
4vz9324st06SYspzy6ICna7EUX+SjMhABbI6G+tQvc68PUr33fuocBOhb08gRzh0
yVzKE3iUGVY6aD7xKEXokSOauYb6X7GvSnc10q6qEaJy8ZLduftP4m+y+euazP0w
/7fHv2L0toO22OYGoGLh+QZ8gk9G7nqGs6aPbUiVv8NGXEAux42vtW3JqLQS9p3o
Nkn7O63RgUZFlPndo1ds+DQMnPYRh9UnSd9ZJqUU8o6kFmXTa89oAH4IWrHyVulC
MGGht0y4pH8Hd2l1qIbhmRXBTppbnShx80i3c6NibMaph0McIFkbuznZTz35v26t
5P0mpBsbpVSrlBS4NqcvlVHTpXepUWUSJgC42jFb8Tl1GEqD2RtTOASUO9bh5Z1W
ZurDsuZjUv4y9bfHyDhvIiIHzaN6rN1DImnX9NgOcMy/mjSUx/ZesSJZ7Rqhd3bo
H5PWytjK0nW2b92zcEdYncStN4yXiI9C2BAZbmMb0tzkH46q0VcnPgDihpZu8OdD
T/PBVDIJIRt115XaxpbFXmQ7jSWddghgIP6LvaKaoe0ZodzF3NGa4R9bY+lR2e4u
pXwjLzgBXzDM8arnvh9CKAhBuR9QRsRYFTGEw64iqaQAW5VeFcRUOfGAskwY9JRd
rzIwwsZBKndiMl2V8VosnXU/ot6/JOuuKTArJqa6UxfnH3vkBOPlDfqG8+xm/u+F
kzera/uMrl3i/cHqn2Qm6Qus/YoJDnCU8eugroROTaARYe08aMTF5PulUtqZWSda
TAHV6i9jSLVNLSO4619GtE+e5vYALM+RPCme8uLLuNwZQiXTtHerGmbPuiZ0sxOG
HORMIJDAGDI6+Fjl3W/z/N7DmrKnKYB15KSIq2wgC2qqGUSbCJsvATjT0iK8nKW4
oEdM2sXBHboR3N+PBzJyGOa3khg5XcH9dp9MJ3PxKY6hUtEbpz3onaLUye7d34N6
Dy3AdyiD0QXsiXaZIEeGwoBWyNQkIwVrj3m6ZtegnQA3DJDQhJBL9bupswsk9y5q
BsO8qyEckKxP7yj2uQslcWaXj5Z/by7BeOsVLza6F9LekDwbCoRKy3wC7Jp2TMh3
3dz3918a09NeRje2ncYvzx9Q1YTXP2d5UR396pxED8nOZqm+iepAGFZhlh8kEx5f
4pDf1YUzSxMi+wuxlpsD5FW/Wmy4jOam49GUb43kia3xVrw37oEbz8kspMUEctw7
5MNgq55B8YR82lkfOgetvV4BiIR5WMiG27KCQvouuHkP9g3tA2+BIGY7TBW/fM+f
e98krR5od+XgOQ1Dg08Ey0KkD6J7y812KUXftOZjtpZPU+nvsP/ZBQd3k0E/BN1r
dqsqP/qXHgQWa8ihHt7r6/GQxMU4ppzSoa32XIpRK2IDnXz0coFor6YYA5QkJmIO
WZ/7i1WmrT3isN45LSDwwPtgBDEZYOWNKQnLIDtj0XCjgCEyxAbzEZhKH1D/9r49
NSGRGl5JavFOchRayxvApTJqUiwCMwCLB0akEGZodUf6IC4Uml+BVj9lehDXgAnQ
5RWse872fdbxBksqCwF3lbbjVOcUZdw8Z2DH/t/iMVg7Nr6uHec4C/XurNwKXmJ2
2S5TlWASJivX8yw47TeYVHPj4yjTWie/0HjF1RVFOJFUXnABJcnrd6Bm8k8jEWxL
YvgJZ0HZdX4w/gkLNvVdJGf3k47g/qofy7uCaxqBB+HFr6+V9lrJUy3U7vk0iD52
Gp4UnQNP6cFRlqSX+N6kTwu7RyCt/lQOd4lKU1idwNk2XoVLCn/AjfqdVrXn5MX+
V05rP52C7d1Z9L3kkrd5xbKYvzHVWCG2LUjG1L5fX+6J41MI5GDIH7whePdKSjfS
3tFsY8Sbz0ARqDvI6+cdJ5r+8rdkEB+pkGzjvDb1KKhHW8cxvVoZTWM5rMhausnk
QMuVG611wj5HwrblVU8ts3HTUNWuH8nMdPHDC3K3fvWtFrq7tM6KUrjQ7/yMNVhf
803pZ4owARGvL/QMvEPue9t2kNbztt5TT8PVRw6zMsNzdgdlo3BmOdrRO/J2S7BR
xlaqXXGcfvO2pkk4Se6lkFIG2n3Nbuqa+AUsS2EwC+5/ZlRLcHWGv6M48oBxQNeJ
oPoFSpuL2B9x8H5nM0fs8DYropsPwEsFVB7rGI6m5uMryGwwbNYaHwanNdBi1bqp
4KAxs/3gPIJgjWKxKMbT87wjLaKVCkJoHQQKKRuqBj0+L8DugHhZffV6fBbr54/A
3n6zjVdepM0mA/7CUvVx/9XGBKr2p/OWqeNlfxo1jjT3xjZmr472EYEwJBRyFCdq
F4yDoggcZN0MoCWvtoQltHgTe0rEVY/PAfIq/Dwngk3jutoao6IwfKlCQa2SnIV8
f//4Glhy9W3QHCSakm5hz9bAfyuzrST/h7ea9McDMLkqkYm0kSqtzo0KyLldz5qJ
DiFLo/kJtBo8nUI3F+uwqAkY4iax7XoNRfkLR1IiBXqfib4VlWU3uCVW8kwW+7X+
oPiVwuGXOGse4bIiZKJDo1FrnIEgSy+mvfqFSHji36dgXA5LB7qA7Ee/5KgMJtNk
Kxa7cloYCiRDslJJKOekSyH+whkfQmZzoV51f9pp67nwCjC/e9nD3YQgHFwMflBa
Z8IZBmlkc7tnnua+RxLInMbAzuNgv3CXEOAXI3mybycpEDkZB1BivsX4VhmB19Vt
hRimLK8nvOe+SZA93E7draa8fNMFnO0Cmbht+w0lVPU7UDGXQrp48U44i3oKpATY
3ouiElHQrDxUCIuakbyqhfdwrX9Gjo78ZCnxaMsA4/Whdn8Ge6dMFprIaFjUdZpf
kUoe1Uvod48qxMFAsI+wFV/zz7SPA/yBJ87Jmfzplr+VJGxWSSLU+43pLwJokwBF
oNYMI1CQsyOodfRjAS4yICuMgBdSnDtkQRMqqgYjzuT0rX2jS5H3a8Guk3eB4v1Q
eGrkPcrPZlB74TZDCd6bo5iRPixyvQ3+lxjLMMV84Eqql/GlPWyfoRYDVcGwUa6Y
tX5oDQhs6ePT3JkPLRzCo5tfKUwYsye3FermwaZw/F08hgj9OFwzGbQ9BVNzFetD
D8IMkuIIeidu2Ci9iK6rbFDF0S9LZHrMbOuxmf4B5zQhcSpcvZm0iFiRm07ylMgj
SurDothm05X/pnU+lxRQ2H7yxZMY9AA9R1+LkcNNPZML9UbfCfaM776AGtu2j5Mf
EQSIM7QHrODfcwjv6T16Sl/ZuOXn4p7/MUJ6ZQnV7SELZHb9s/Ks6PGZVXmqUKTU
lYKIsqHURDjWM/DBeDB3k7hBPNBtNu2kyiCSV4d2z86l3RPenD1QlrzFKLqnZuUD
JW3WxY3jTt64Vvt/mHwx7ay5kIY0YR2o+7SGXoNNBA0WSXkdolFU80WZgwnQgAP+
KzgaHePTre/gc7etzq+jQXBslltKCeg9b7CLbudQ1+MCPY3AIh/nvelYpY5kwp6N
iJQuko9RgrFaMRLLI8QjtLtzxx053m90X25TG2AwhsbR9ehyUW2oZrJSB99iTpka
WnRg/wWSBOmt92geHJI8uzzkY23TScNmNsRsqgIOBv8K2dnP9j5HTlR93TQ6xS+C
E0R/ClEXBINoIos/8HFGuSC3cbCwqt98jw4qZ8M6s8gxajTXE6gWe/l9r8u5lpRK
MwSO0vji2MkwD7aQUibwUT02f0KD0vKWzgQVGgV7Ns4bjmqg1XeovnWpoa1aiqVE
HS6D20kiBVw9AzSyjXmGvAu241Ltg05I7fsVK+u2cAEatAeXYvEoFYdYKlu546Pp
Ol9+E/cB4WizyGUwJgDIEJc6XeRTdxIZ5KCEd6gEQRTOqdbPKvzgH/WJlYgswuYV
V/HqhWfO43kPMs8fd6jnLQc33JX/Rkmv3OJL88+88x7ngzLiPcbWpXP1aNzohy1s
gf0Yo7rk6aX2i49WQ2NGUQ/jFd+UaHNvi3E6uGM8chzxfXboA7Vho7aW+20PTVKs
xLxpzJZRr7Z/H4za8hWv/AQHWfDh2c8Io5xHlEyY3FgMfi/MYJMEgasSErMLM12g
4vJY4oetF0BBZZXDS7WoUr8WUZYvXkCYTn8aFI/cOCpXbOCIMukFAJCASv/gqKPs
uv9HrKZH9wJo5b5NSOhzFB4uAIixS6EkKQc7hDiZsdLZglNkypd9OB1fPududQfU
u5EVyc8JrmL07RTG5JOSJZ+v+aU9sKHpVA49CvPz8ZncCvqs88F+A12j/6dUOhdU
wqh5OkPdLsAXqCXCrw/r8w5vN1AqXb5hZAiapVHJ32wmPpMtMVq78sIaBiZHQW2s
dmiYF4Fg1SslYQwrrxz3PlViB4T5SWSYXOomYfcMZ8sJ5lGBROfwJgvMxhgxWLrU
gTyio06yIgqmPh58D16vInwj4tRD2Jvv7THe7Ppq17DEcVDJQPvMSa2169b7Rka4
YPaHOI2w5KhK+5sFSu/7jnkqOC9lIYmHRtrZQ3BV2qgohZdRBWNy/xtSxgAJeH6k
wlpy5/z/FfprbAlPB1m9Fx38DFMkS2+fts/0dZV4nOUdyfoW6tEHHdckO7Mr1qbh
JfpeCBxaMH83wKfe+sp4rQ+HDnDag4qkDSzZm+5hsfCLYGZ3ogRByZt6ffWJrbu9
W9Qwv87IyQ5eqCfI9yXdFVumlDPzk0PFwalkStgJIei9UhwHaBBNFILBWTBgJba7
3MUHqfzHCew4sCFqMz+3EPbgsnKpdlsxT7Nm0bFBNtEL1bPwemqkvwdqq/QdzAvI
Pj6tPGMa4vB4seUnCLRdip9VuhBx2WwwB9HVu4ytl/8HqUTnRaHzQx4NvK+yrjsh
5UeXPeFFs2PbgNgQnGqULAzIg4hgVzyxpuKAV2yoz34MnVJvp7Y46unt/D1Afmwh
dev7sdKkEG5V9QztFNAzxuUj5FF3+exP7u+TfV/D/FHXoYNcxy2XHNhu+o4Ez7WK
oPty4o7Re4L0M1idyIAEKscQ6BIweSjCdRhyBM7jfRCsZbB2XHM20FuElsUu6huc
vweogoPb82N9GaLmeYa89RimngXDg8NzpAyIeQ2YWzgjdm10w8hJzEshVwGxY7Vl
HgC32MPk8nkzd9PoiAFoEC6oNMFwukJR7n7xHQimbiFSAKXDgdrsHsjx0mSD7eyq
eptYIqKSH/ZKJ/8G7pCx27AdibyfTnHHbeIdr9SMI3n0aroe9IsU50n/TTLDHLIY
yj0XwC+Mdq+zflGvvfsnDRphLQ9tnbu8J6W25zMl3L9MNMfzmeGwhGW4fphePdKA
XXU8tdxkw7KjkFvihEYoYdZP5HaPLR+iMdfOenRfVE2NgR8k0Dnhh5p7M63KKpEe
EKN63qOlyNOgn3BFIcY9xmuyzcEPWuRotS7+PCb4DJVy2JitD2bbzQLZzEuc9BL4
Z9xColnU6Ft8KKHfCBjK+0xREJz262LeZZPtgCRi1/x77bKRSU3lCP6QVmDgvRQQ
tCts6y8Ka2zEjkwj/6LyUpQdTudXd3NZZpInBtEbC8QG0Uae9m7mSlYUfu/yXNd1
6x6sppgy7JOkAnHCHCs2QDKTCazHFM20N+8lApVejEalvfkmkgoIM57sKnpnBu2Y
3MuUsN9P8qK29JkEx3rswaSGX3qUyw7LN1NFZHYz28X2Z6hROcUM96Sk7hTrBe1h
bVX/w2fwxr9axq8jHt8vEr59Ez3Sw3RvUowowAJVmYuZSVmzhOQANwisaXISMlwK
p1bbojxmCCBlHohOrVnPYktA0Ava6h6TxjEgEpGJRz14McBrfltBZf0fy29An1+m
BlE1HzJCNlle/NmrwRnwMWwnsgaAtsO1G8ayiBU5tHgcFqhlYyiLIEKLydcY0L8U
qbPxIbLdpjc+U2ndWasqc3IHhmQfRHdh2Pd/JdDCxnEFYHybP4gZ3mduetsNyfvK
So5CYkOyBTyT1fgEqsWKgnZeng/IbFUySYMpcbsKT3Grr0pwOX+Xc6xXHgvF0T7y
IiCKMNU1wxQbP6dyOOnViwb43k48He1jZLWqKGdPOQGMLNt3aBiZJirRnYh/Htb9
lqqEFK/EphD444kIChEipx6J1jbIH44jYpeU7ONeULZv/EGXQq/CG5t8jAwMSjw/
921gKvpLH6QCkP9wjCgJJ8A37ASUPczkzZ6IVFE54viFxYSXJgXkm/G07fQATDDp
YiktHgPFINMB45M/ptMjnK21HPE8j4h/syLZ6ly2D/1SMUd2hLmTChpo5rn8eyzf
qZea6326omT9rdZq7f2xmInx8BazNhP0JjmUOi90qTOPXIIJsqfu/3nnNIlN4kUS
bRiW5zwbCpxB9Ir9FrKTgAPRZV5qDyJWnRZxUckdTvvJRbs/2y25RHpwrJmcA6Rf
Rtb9KfZB6OwvHJa6kas6Jp0+9AGoHrWq/6X/R5sXxTn28MBj4F+6LyxwOuStnSw9
rdrpyRc1dMVuMM+DDSa+j4Y/PjhztYsxrDvcbJ1IaiDp+yQeEe0spm+RFTg3U1nH
ixSeIXOm4j2o92ofv8ZmX8E8gqvt8Ss08z9B7S5uqB7k4qqpSGfq2y609xz5L1vy
FcJOKJxdgzoOJ0unvHF7xtJB4k5FO/IMkBECajbiltLrPN+Oez1HVc+sioDRGdzL
XHrxVKIaNb8MQVVSnM0Kh5RbnhUbf5AyWxxaPZlm6i3gfNdijsxPo6xZ2f5ZDdRr
HcejSPyCi5O/qIbocQ8NDi/3CbkM3UTn1oyl3DbRX58BeY7Hoe3rThhqZVQeCOAS
lbiB+O1clElR1hMddEo95IqUndjgz1h4muycLAh06NjCDMldG6CufNzhEBZnt5KS
0PqsK7AzaUTga2S9v4yl0tWfsM0X/x8BjOHKryGEYhrTRekhA926jIgbtciAG6He
wkyIWc7f2hQKlno3D11BPfqcTrwVjw1Xl22dPYYLeWx2+WWUy8YP/rCoIhiX7zDi
mx8CSA44lguokcgD8/pC+i7DwtDp+0U6MbyWOPIJD5943whSsZJ4G/eBD43KITWe
ZeC8JS4qJtdAnzyazttBCW2s8ExUIpDiheD/LGO3tP2KQN+sryUQGwPiWrnIZyXv
i0zOqe2CNigw5DqWeqwWTvv+5kPpiEIO83lMCcmRYIp5YH8QMdhOb+z77X7rhGDj
COsztl1lK+9v7DZGbIMvwh+403vLQ3A/3OeJBCd0ASVPU4Th4wn+GlJ07gF55wv/
danC51Y+DUnrftiHiuRCf8mSLc89p7K4Dr1mfb2tMUYrPbniXpAoN1Ich2y0O0Ag
o9c7IP79CZNiLGdOoAGdyetfs8+VIsDJSeWqq+tOpZrKnV7q/vYlkucXyq0f7+Vx
pWvIi1AZfiLpiF5lBPvw1RfiarhX58O0pdgf38Idgf7aGhsCHMaYxpHkld8sPFtB
b6Eaz4A/vCC8yjDJ24MKp09FeozSCRN9pfp4aepW6O8CfrQQFd4iaj2Q5PUdeJdc
js82ncbNIMdGfXVwQ1Wnq7QXD4nK2zxrM5w4mJmEZf7TJu1PtAWVrFQa1mKc0qJ5
+GXksJfZ6LMv96oWHj179EaHBhunqlzQ3GPnlMAQ6PhUtGSzcdos/eP37wEra2bj
S461pfyWtyMVJgV2U69rD6xIFfFBf4+bRtzEgvDk6jIh++P1+rpcS5mdETRHHZI1
JaB6ky24r7PsLK/CzaxnQMq43uqZ55zj1Nw3dQbymGmeUeuNUX5NaD6Sk2EwP521
0TTjvEwWp3NXNBqCrNMM4VptUkyO33IwYY7EXaAW5vgPkeU+n7LZ6gzRBooTTxp5
HU4hp/e4VVi6f8xV+aluP5UrKbAZwo4AcijJTYjb61aUh8vojCx7CLsdIumbdNcf
WEE8T0WaquqOggmklQxhCc/zjoUXpa8w6lieRrxG12pzmONThJm/76CA8oTOv3H1
mwog1Mcuxc/PzMaVGUJIta2XWTBVyLE1wVN5sOT8LnQWxQuwnHMiwLfj0rEL9Dw5
ykic68bLxF71HCLElYZ8FHrJafvsvH1cSBrXb0bt1CE5Y+tFMT1UR3Rsweu2A8dQ
ZpK7JsQkpWJN2hAhXBSeYogQxB6ft114m3r9Ob+hj4g0nHzAB5D3VfCka8ZMie2D
HOZMjqtkNTbYlWQh7btH86t9qFXJPUWaiboCJyI7qF+j7igthE75/vn7niSmB5E1
nZgiBcmAwaf8QN33xu/puM7w4kyNn+LQVkpnz2fL+RGNamiN56grz4eCjYYRDO8U
fGYK5fhoO5g7XzYRaq4QxCRgTkzPyXbiaagekUzFwqpKL1CUCn0v7MpDEM9pL1UL
mxoJO7RPH2ReiDJ+XDwJFjJugvM096u4ez+4QZ7zhGp6gsArAjaFtpXRALzO0C/J
QLdf6LL8zcIBXGR8/XpUcQ4UzdE2Tu1IQH+5idZWz/+0eufyJ9kJ8vnUtdTRO2nG
lPNah6NitsECVJYNHJVdeqsbTOJK9Deu7l1joiHPNFd0USR1hRFt20s4koEmfdLf
4NUpS1Nd10rA+ijcBVY2KsOaq+9MwXsRXD43DzAwgmSbFnnaTs7EbDi0acoeo7oP
kd4Z9qcLDyXrvhSx0YG2jklekSW4J5l67BKcv6gjeafyMph3mfLXmyielM6HpXva
1dT9Q9w30Z/ZhAD9GiCLXw/zffLJBmQhzPEHf00JVWz70bl8/Dwjt8fhRZxFISVV
vhp8ueMcdArhUOOp7/pwFmGCrlPp2ZkrwkzXBKu/jJup+8/FKLVNSkF6Et0k6jyg
hmn9AlwUutTO1BJYJCtjHGlnRbdSUN+1hHgo5B0nv83qsVUvVpgnf+bTJWdNynva
BDY9AFiM2sSYs3G/6TB4qh+bCF1SDStS+KcVDHn9K4EnxhRhywFeqOxqrIi6bU2d
Tcwn3baMtgWMvXAdUVmAAVfKdlj8HzTWYlyiw1giqzWU4yO65WHlt3ZLULCrqXQS
14C9zQxpmlcrf3MO2qVc76NC5j/ITCMynv1JKU7jNygVDT3GlEf/JAkKvQz9UFSm
tqsAlLgBEhXMWKoed0OejepcPCh7Kx18mZQky3aShN++W1ksb7h6Ts7Mys2UL16E
wlUWmr9NXCoIl0N/zWHrA1z/T9180LFb32WXQiwze9YQJdJE4891RedxLbtA6ZMA
g0ffa+CuTwYTHZ2H/p6Cq/K/nsW9DbTFpWqZT0MqvbRpoLjYVbsmQq4HFAzHOYnW
ZTuMODkTFGQDuEvs2TFyLCEVDZmosQKfdwh9PG2Jum+fwqld9SahVuoL5JDXm5co
T2mYJ6N+zciFN50lJsdI5mj+9qzAe/8C514xAoyVdUpYcXEHs+gnSKIQA1wEVfma
drCTMnoQQTPLLMR8luHQmCKAJ6XFDXlKlVgAd7k1+OoYQ3GLjFCeq+Mpk/rbfAlJ
S93HFe9OlZdb2Pc4X22l9EO0LlX2uPH4fP64HqDlPU/r6DPjvMOs03mMThOxmFos
WIBlFSxMFHQa7iGWOJhR7tqDQ/O3pbxZcjittCt+XXItZB7kIzyicJKZVL83vtqQ
SAj82BZta8mxNNfshCv+1WZSQe1PxLDZgzMSYp1uHATdpj/LGwsesQYh6FXlnBof
1+3etf6yuXZC4rmZ35c26CxL0Ek9eNxVXOKjHCqp2dEHYMWQmOrF0SDsCMpiGKiy
ciecaGCax6/Gvuq7LJ6g2C0ZBTPSuoXCrAbENrVrR2buWyRWD5JTIsFNtl7YWBTH
V7pLdoO8MIhnLMTdkmH9EZu8BdPym+0hqfrbeUTiTjd0Pj58JVNtxAPkX6H5IxkL
SxpwjHKhFOuLHwGUi4eqi5J2lNNC65E0jMhWimJHEqjIKd/t0RBh+jCFQ5k7kr/8
jgFxzX46Db+R49qJvEZAfFd8HAKSwnok+EF8hqKEq6yZ6OZbIhUDvyRHRY4KUo0u
JaRRo4J7aPKct7tYBH91P35KjO0NdsSR5TdoTbO8/4alKdYd3o+6u+UDae1u9ulI
6R9Hdeho7ZeZDbXcBKg00Ol6e2MKflPMbRf6OkHrSRFU0zKuJ7WCnML0L6nw2PVN
2K+g+d2juVv5nxdNm/tnmo2EdMsqWXGgF5mxq1EURXn/F25+ugCwSYrK3g5LwU4F
2uY7mUwpCc4LhpkbASWLKY6xECgJ2vaI8jzZLjgOuMSa8C8Kd//0H3ZiBnxKaFbI
v/p6Xlx43W6M1XwSJVoFh4gCCtI/QnKe4ZlQ6PFu0OehaMeVP9dC23GjCsYbyd0S
THWXyiedJFkYlyYUjsdstVRH2fW+BgJqzpzgGslcbYG83SlxkmXZobo2hhHfGHzi
D7MqvbqljCIfKidfbC+NEN+49d9kupwWFbS9PdYN+srEW/JzrWR8eYjXepsyyvDc
duLcCbULXJdxgbLA1p+VZ8Sb98iRTcThCfBegCs0KHPfIQzQgQv0tLgua7d8riOd
VJZel6VIO+4novSnh5+kBMJJfvxJAEUT4wuJcxj3CnySFz5Z4DSXRxZMlKI9Axh9
M11EbyI2bF2mjyF8CZAJx5DR38ii7QR500D58Lxw217cXpEQj4bW9wyUgcRZiqCE
VddrG794UYVdSX+HkrWUnKVoNkntqgbpJZ8Lhtejv3oyzYYQTsVNJUhvLmdTf+cu
xKIHKGEN91PEa3UmHjnBu3718mSVdca8PaF50rJ01qBr9K1qMGNzPeDzavIPmUgK
KgBXs72dWvMvVVauUKhrtegrdwcyJFKTb1rFTfSoRa577KmYn+W5pbyvwY+ntyCd
bMpOH0vEZSc08TBwNBqWj+G+I6bufxYeVFPigJ1a0Dr2atpVLxoJ+E/wpMJc1EEJ
W7TuQpMG8s/jhRfjBLQ8x5NKFPIuxcyp0ZSIijhiQz3N4g13pm2PU+0fDFSd9aME
LEreoAQR/plSjT0wnMfO3wPu80He0eEG1MHkyKaToIhiC28V+Jh2uAEN2aKqPZCj
QIKtbuS5LZ8u9n+AUiupyjiSNV3W+XEjxUO1rIwDWVu2rMXKVBjZcgagqgOARmi1
KMz9493GrDmPwzn+LZjxsXfibVtygpceUzp2t2UTNwSho71GGxcTlISb6CJKfhRh
g3N31Xhfbo6PqqKrgCGTXjHCz+kT2AUdfHitURTjcj4o0OVzIBj0dJLOavouEIiU
XjWFAmSsNl19Sm47FzhDx5UxlFq2CUjhdhMd8V7DlpfCJWAqnN3SQ2OhvsVMufI1
P48U1aJN6LPdonNrBs2/LLchFbgbgueU+D/NZh8mzJDD2Bev3hwhC2fqYCcXmdfY
QMYD6PhRiaXxyssyPkSC3Mkogl20zu8SKrPC3t23FYy9XQmEdLz26kIvi9a1muo6
OeVlc2Px5u1QfRde3oKirBb0q0WislRw0r1Qdn/lTUQKvk7Qh380fRLevRYqB3+A
f/AahqCchkipXx3NM6Ls2hb5hzWrAM9MiAvAMyEjRJ+BEalkKMu1x6qWHZQu7TCr
1v5ATEZlBASS0cc94vYW9T1xAwpvwEy/hqALib5NfM785QXgbc27gYqm+b3KeKl+
lKyaW/gRZwy8aGv9XK120I4zLM/6iAlDegVdXTaovDQ2gAzKyjn+X7g/0a3ir+cI
s/R4G9tNqfqVVcCGLzKTSKRQFPqzbabzAUxJ2o6lZnz4y9amojXptCIiXht1B+02
XssLVJnoiMqBAzK7gJeaZVhs0CjzbRJ6g0Qal2VWrIJQPI3feYFRRSaFqFF1xtBv
5ieG1Pcc1FKnJ9nSzs/I3Ev0oQKCn4KpnD57If0o8H/7y40GKQAtLqbEWpq3fy6X
uuRZ5JtkaheXpEz17RKkjK15JSlD/gOtSF4+p3QRLYVYhBW9sQ8VHkpIjLwLrEQr
aJq9VXfUgSejK4EH1HhEWsXYEQTjNvSHqmZIf2FyRA/rdM2KK547/5RCPjwTfU4Z
yvrixaNzp0t2kQbePS9tirumnmitLZ9IG6RZSNriuMGhgUEP0U8tdOTWN5obYKCX
k426G8+uz+XzogKzhBpdKXpwLkNKavks+mmZP7k3eo8PdPW8yrtJ5PJN7DM9IXJ3
Nz7ih9lvMUFSsHgcqGs5sAWcKZ7+/iiGa7s46gonorcL4Uo2rucY+0Jqi55AI2my
8lNl2SSzLQ8j4cMLfTctP5NeNAD+hTTwcWb43r0b1dO11f7epFfjjyK32rvufpq7
zR3dHjuPRWUvK7Hqxhzp2ohPYYzBgHeFoFkBrJPZyUj54KI4pgwjy/x3LpUtHBoz
ILxYW6gqtphO/PPm6xMTEH+Wk6z6usrAvVY3IJijoCXP/dCgF4ipT6WbkH+GGm9E
yp9eITosV7kyK40Ffb6mNMft9l0Qc0E/FVj5JUxk+ybNFx8NN9DrhYkHNCsJwMrB
5CBTbVCunbobwvlOEV+5wHmf56e3b4XQLAfZhGKGRekRHGZJY9kNphjpzoGvCx4v
VoBkjlKa/vxCarfQ+0cOF/ApjgbOYU+MHxU85loGyJrIx8DPTiO5Y/SLluM0KXKz
MI34BJxdgN/deVq0ONbQ44vlrQean4XnZ3pnG2GjCAOX4edl7r45tJ1pslbzN9oJ
xL/FfqMHlfnohJSSy3EfJ5UPLZDbGemQ5oYBVieGGmh8a5v75kwFZZY9wtjP+W4s
iXKNKpKtWPiY977A6MecfbTMeYonHHKXwLY51uas2P0iVZarV1hGjdNM9NE3uuRp
aWOQkfHMG4/9ryFptYPX83zo8qCTnLEbGDzTtAcCalt+/JbGvI39IrXAIEHmClKH
dTk9QrUcTGK4dsZ86EaPb96v8c9uyqj9IBpI/d+FBcXqRPUiPRXlwiYuV4MTMsPl
DgjVyuvTNU9O93Cz6HW27aTYI92DiKCyQpvWQ0br5mkeJbTcorTppdOy0VNLU7eA
6yopuziRz4MkpkNRM6vJPVP9XEMsTkjDwpPHGScJZO4LJDuTgnS5cEzGbA6oW21g
FEqLo+WqYrPY2PHL6CjYAGq1JlEp/s7UDSLZQfhW4jjEnS6Un5OgSZkE39Qi6cTn
3S6STA/aannuP58y6Om/fsv6t4UEEJlwew1tuzW8m+lq+qNfsti4JT1UQXiKYrLU
v2fkicbhSxQjsK9jz6YdjX8r08ft46cqdISqo0xHnk6ckc32zXB2x74wCoNbnYoA
/wZ6OGfWZDjQQwgIFrKhFf7qXEtFw8BfU5SGzikTuCcosOmyDwofKuQCH6ZpL7ug
UzfFsT9HEIGMsG6RWDVqj+Z/HjDlAHz+90bFARD6+VhN6TOD2M7oJXDpHUb0oO1U
bhsCw7CBQsnZzINoeWwNi5OeoZQOTIeF1SZl8GN1OQ8OmzwMVTFqINJR0TDYFaYq
QFOop4wcpN0wV2JFevTjOmCIMwlvyQhmlqTYtG/WD0ZgvVc0FHmEYvrnCMroy7Im
xRKVj1fIVpX2Go47JaAr6vuxf1r4dLkiSLCEwW22OaXfAdyYnoeSIjhfrpND7KGU
9n5ii/HO6CpjQVVvRSoy/ahYszYoS30U4o/sJaLJ0E16Wk5yd/q5pSX4M0QrkTuB
WzacvDN2fussnza2mbj3bKlhpbBZ4SPRClwx5VIw+Y+10Dmu71ktm4VYbFfBQqwo
Poe+DxuecslXuxD0dj5ZpRoNTUePyY5liQFwnwF8atgdsjsa0gIJEG9hdjAJr7Kn
ZQDdx4pNwY3c5sWrE80FJHD45K13qf5SnbHTOz9r1266WCe75tFnSdAf6DrOMxYv
eyXnxw8mmxcem8AI41vXxDT+ZIq3Aie68Vahz2fijq4boWzPU0J4RfwepvUgJe03
rJ61LLZkOOlwFRDjwmtbQPMSCScf5deZOFAIxzfx7ErSe5zdJ10zYi828zQpwkB6
xhhBtlQft15JMWJJd7X8F5sLAPsm1NXF8ujSCahGUyjctmjOkOSrPuEZP+WkGXxM
hI42i2XTwytCHB4C4YGbDIV63rYRlvEqCxAAvmTKUBcUUtWiHxd/TA87UDvOCqRQ
Hdsr0YQI5iOOvwWAtkV2gI1CK91h04PB+wA4IU8ix3bfi0O9NnekxEoZflr9fOHM
T7CEiYi8eU5/OYkmNC/V47bmZ+RCAtknYw5u1wZ6q59yrUn5HBCcTYjIUVYO8wSd
/uwInnuXAI+Y+L/HZxtPwkuL/3lXkoB8BBn3pBgpl/waCsvjb3oTSCiGkvkbgKu/
xbZG2Kk8yeyH5PuPFfuCI+IbuwFDlorE5fh8vTyZIQvVjt+Y9DXuwZkEBz1J+cQ2
3iMmIkm83OSkc1Xqw91PEyjRoGSE039Tzrbi2upvneZgjkVivY3HRJAe5mbcuZ5S
RMJ42UmWfqI9nNa7iweD9mdjr5DoPky1meFkDZlThFMdgUhVr+SXRdIihVxZNefl
NwCGe77epMxvcKYtzc0mKTnHZj2C2m66+LEZTw5tYnnJKCeu2CUTGs8FzwqyzVua
aan2CWxSNdwlJDAGDa9dSIUlItHEEaVOxlRpftwK567B3ye/fKBuDHjjk/aiJVi9
2xt+GKWH0LoCW1Pt6I7Mp3hG/C3EuTovmH00BuQ3jyzVXiQmXlH4GbCRft3NOjRV
bRJ8GlQyyhFkfPrctyIUc6aEInkKJc1MfB6+NJAnZ36r3MLpTj8XaLde4U+Oz91i
Vwo4lx4b3xKrm1holj9vfpEdV2NBRFC0D3+VDWpEOH6Wp4Hpvbv8FVdKNwd4L2iA
nfbp8cgnGPwvapFvqi631eXwL8uE2mU6nR8sKFQqD3jx52Kmm0k9sQf4sSs+cqcF
ezrFDJLWJlxVNz6c/cOvlg15JCP5kpIA22fTk3HcaB9KyBITNZt4YdZCPjU9aBJL
swf6vDh6hw3CWA+kMNy2VDa8DYsENbLhBy+RBX6aOl1qJ9Un0FGCYVDOYzkyray5
g/NVrutxqoSDMYowa81qfU5SflPpwOLJwwwx3MnNLZrb6TIFmYfybb2HbG1eJ3Yp
yX5ywPnyNlz/JF/YgDA6k5pnfboVKkeDDUKJUOuHgmx7Flfk3iVQS9o9NYPkShIf
vxMCxBl8RQU7+Ljxk/kqHfwafN9WArGR9UUr/pCPdRZWXfd4pHgAwLURbIlkZoPt
2qlQZGYn54vH5OYvZcNjCa3RowA3/0+UTapRHzUJm6oDdRCEet4EOie4/U62Woin
sQnsYAcTkWeMYNwScWKTdhsAFQlN83smy/rozWCAf4SLkoVsec2hZ3oBP7sxu5BY
7Xn3BCxAvtFNTToXLohrDELWuvMa6Y2eMvY1Z51paDq+oMy2z2dlSdB4UAPPQdY6
0gMbvkFFwCdKBXFe9AjVjjmc67pF262owBDeU3F1uF2rn/SG9/FzRQCrpf/KeZKl
jGjWwl+htfRHPuP50efQUf6Ex+Zs9/6s+v/h381lO08mPta++toesRoiQFQQypvx
ZaYw5i9NEQVZHxkkpC0/fmGuk6kdHE64bQ0kgA3v0/mq3Vv+VX1puc2V39C+uhGb
PQxj6MBEHC63d/px1Sd7mKcSlr2zrC3RTQl+VHGaQobn5tnafG0Kqbo2Ax1q/bR2
kZ0r7Cd9RgyI9911nLrQtoJdp4unnCLDW27R3XhItnsCprP8a16Ao+2rvY0m6kLe
XQi/q+o9GLbOWsz7E+LFv0W3mDepZNMgz3fbWVkP+rIHVAiDyHIeSXf5We4pqpp0
Gl3Z14ZTxOU42Jc33Nr8/sw9D/NWv1ITbIlviSSjbxT3gdhPEBnM7LeW/Cveb286
Af9TxvnAuNw3FTBO86biTxOaFzTm2nwACTUEKPzPNJNG6BhZA0/wK6ax9RrsNJJd
58fmBicZhhAOUXCrtwccPGaLd5J0eXjtK7uXphJNCqFGFUxFrgyoZp4tf8HTzBdB
hmMU7gwkOJ4Ur+jfGps0JuxiY7TtHqDlx+8njwa6Fj8wUeoVWpH30UN4e5ni3XBv
4PwfPKPmwo3ign4iO3uuBzhGaRFBv73cMlYSCv5CJy2dn7mbM3CPi6kBjCLQ78vf
/gX371IJ+cdUCNJBNtW/NhQoiRkdih+6sapiPmfXx+lqkLbyq6lejmw3oXZAJYcS
lf3gPhSrYGUUcX9P9pjo6IqX0PB1E/f+woqFzyBxSUR71KbHMAvc6WSjdHl4YNDn
9sWeKBf19fy3B/7l7b8Gr23E7MtKymnUKpV87o/2RzPWLpsftyXqDG+jQVtWt+EC
TyJ9/OzwKgP/IbiEyWEVaan6Z1ANJdNkMSuPzqVW2btnk3Db1BmzbVVGgzWCIoOV
3dEKIo3WmtyMqwhQAdlAZr/F9Wp5Lgc0/p6ZGFRQHNzelgxBpElSQmw6NYAKntLl
bmjuYnbnP2yFV7jSWkEA+/cG3xw+B+Py7LufPaCjsG03ucni7/k+EFcWjVPLrzWU
EhzuJcS445zLQjNf2Hw6hfOeVwD9s4U5QdA+EZxsS9Svnbe+QW0fCEW2wN2J/YbP
azZ9+8hwc+mJzETl1jCaHkwG0WcmqBuKKajROK1lr48QvA7rp40/dUdIRFrqWazn
cOklzORxUoSPbhkAX1DmFn/6x8eF6rHcxphSS2dNu1819OCNQOBlFqt7HMohuL8c
8i8x/oWYJW1SZ8+PEnB6geDH7IvDIaXwAgOmOR0IfSHvH9BVBtW2JW6wo2Ag/VMN
tB0e7xfItm81hjnrlLMIzG5eQ3Wg88AK26dEwO9/OSJMLwKu0aC5wTjjItucBuLR
HPnq2v/eF3615qAnrQFBihI1W1O631OauxIx3M3u9NjOYKuTIQCAHoz6IoXADdGu
CJ7iD5AiHVwh6wyENsL4mod2QZUUhXpuzfCWD2cCeubY5UMQA0kogfNBL4i8OHRm
TTokztCJ8jtot8Wqde5CaLodyZN2oeqoQvLE3CW8iXVE3aLssoU2ZEZDA+1KjV5t
4G38/gc/0mUR7RVopxSyqPxIdCQ/DwCL0L9mVyN/s3aQXTWS9P2oj5gChVmwthue
lSHLI1R9JmY3GLg0LJ27KOE2w6ChG0H2fcPgz1TNTm09sdWDvuSV1PowLanj+0AZ
dvjW5eUW8DKQuT8fPMkaTxEsZ99bx85v1tAyzkMxnOjijv2TTUP4aDjpDEHLfZKo
Ca/ObWD3uwFnk8aJqkWRhlsyRcozfJIb4pBnOA4ksM5nf/e2EFX7C+8c04wWsOcp
vqoJc4rSQzA5xBA0UW0bDjhZqjnWthICSDck5J9ydGvSUy5ZbZ4UDXDf7lwTVuBa
KTaJ3/+37rTOrcawTCh9yTiqLGHSUtxRvtpGCA+t0chG30m3sZlHhB/AVQC8NMNR
woC+wVE2tEJL4duYTM+2FqkkTdd5YbX+S/I4Syl6d4DeIWE/mUoYfyN9qLhhvpms
Ubk/blYUnU++pNHbN/GRfiQcNTlF0eijiCbk+AbSpr1s2VHye1WT1TLY6yvYXH5N
QDZtoCo7cmhlty+eRbOZi9A+rKnBsRfRgdJ7q1smFreJhpLnOcGW8aFDzq8cYFtP
RDQjzlN6YgiVH9LX6fyd0Co3frHpDBc65G6wr5VIFfp++Vk69zwmxvzd015ic5SY
ppzJcGHnzsjqMCHKXlSDc03ngQY/dU4Rle8Op2161UvENmKBR12ewXDC0gTlaogd
EnfYruOBB8nPiCHFso6NAtcXjJWX1aJ3S8YCFvRlgU3Cb/+CuW52571Pr0LIczQo
HZHyhnWmG9TPgTiEcmbZi40E2+Bc9G0Tb39ePhJfBkoErVERAuzT16k7lox/hoUl
IygspxBSj7L5+bZZiAX0vjLG/Q9OfrThQ3p1IXdmwuvbgOF4hoAU+hgzSO3uKaBV
qycgAllq1cs5NU05aNIRTYiHoFGCV5cocZlnO1YJFE5QZVJFb262ebQpaRJ08q0d
7GH+OXYWzhEgLu7ceNFwWf8FbBCeIdlcwBXCBXdo4E5LJTh2QDnr5aY7y47NKIn/
BMLQ/XffVSvB+ERIQQB2nJVJAjUjMLlf0+l7lrd5l/dHM2c+9hGUmfLAv/PVvfBQ
frxoyIMNk3cmFtFyoYUicpi1/RDS2spfdi51KQCRyyjrPqu3KlXGk4GFGhdiBhWy
XGWd9WeiuW9ZURfLppL1rMBdB7rWqdbd/eIYzVkwXUFx+gr4ZU8651mDfFSbgEwQ
U8qQoJZSMU5eXDKT6tGf5gMcZSVvlC5l18C0jrRndDUMgivwTdfD/qpAf+hcVb7v
YHVwmh4ULdJk8+QKifIFGlfADxQykrDCCk+iu+ZM+5CpaTy9SDxlwhx3nSOcAKUP
vJsnQzDPD4m72+HhvCeAY9qyrKweZrCQNogV2gcCsGuc2ILqXgVuTdTROQbqvwDJ
p/naS8crqjdjssCcJEkRerzAfzza0i6Etg5AJnL6hzKNHX3U4CXXuY00dYnUnCKx
mXcVbZ1p2UR7CHPo+cXgo2x9GHjlNfCk06kH7HPnuyEUg6W5Y1TfGF6ztV2ZQKOd
ivccn/IwDO5+lNIVQigKbgB3gCbsOqk92BVbUyzCwafkqW7kXgLfyuk3d5Kyzs0A
6haEiRAu9nx8Wes42NG0+udkskCqFjsiNuO+fNP77Yn9bpVp0lqLexVqlgHhXmYL
QZ6eQ/Cz8z8OSasoO0WUy63UyndnjJrrzDBNURUFQryo58qaRG7L3kGU/teAj5RZ
5T0jZ0JYzkwCIvCMW3niFbQQVhK/CiNzK4BUj6eiBGYXf54kQVxkcRtb0/Y75LmE
KEW1DJWVOc77rLYimgaR1eURCM9E4dLrON3ExEFBze5WyINP3pOo5jS45qvdyLT0
K7JIaXIl84hSqmIwDRHxumSu1LuHZkzlNpt7Kv0RSVOzPj9mxzPsbQBt5t2lqDFt
OtquZOpbuPNKZlENw3w+dO25jxLMGoKmUbmkFqtIYBEbFXerbkfoWLOcPbFgSZsK
eJDFLlCS1XvIPnauDzAvSPdMzB7PsOABQ0o/0jaYlAoouLFvXMh8nKPEmRpFLQP4
OwXmSY4KSjNSWCO4qMQK3P0M6jZvz8h7g+4UYag6+wtmROlWBaWh0ml/zGCI8RDL
4tP+DQT/940sK/CPsz4csHzY95NpW/BhT5LRkia7zyYcToSfRCqpj1qKqMzk/aTu
OUio2+ngWD1Ii/WdpVM4rth/5aXoU8wX1yRpE9gdtrC5+kp15JMlQt/Vz4DlegZA
5znnB0atjqbvzF9266+yCB00RdofjfU+NK7FP2os7OhHihfdKwxU1Y5JhGmlo10+
jKFJMb44FRj7mryPu3arr30OydWT2R5JOAKHMse2LAHBGuU7yyZhi0ArCNulNGri
i4AH90EnoBMmYUDoydaHru4Ebs+lO5G29DagdHBAUZbeOLQEAfiCpRh61AxlFzT7
o2jHlBNSU+wANFUzts3PmkuKBGyE2R9bKQjRCF+awoS9diUB/TgyDpnuDV5FjJP3
d9SRx+M+sG79L/WSCe4+DcdnexYy3BhV/iriAEHVCEdwCRyQG3Ucq5YtGOKCmd/8
hOPVsBkUAxCDK8NthINmJXiyDBrKNjEbGN3Y/FLcOEYZvcsECFDMoXZ/zRyIZwMG
SwO/w9yN0DcVcrUjpwC5KNwJX67t6S/KPt5zeCi96Gs32f1jTAFX4Lfzn8+t6KWP
DV8Jz8BKkX3SZG7hG5CmDRIGvdgip5nEvSw2IYdOqA+nJzbJjUBJGYqE4BcfwwDJ
sSt7+VH4T+6ntvqNOUm1bZ+IcDAmMnR1/fb5ExpJ1VWuXaR6jpkq7PZJ3ojLZqJ7
aRQ5aAZUPWd7js/kie+rQEELQG9JQOwTrkr13JOMkd1drPWi6BgvTMsXnyjds32/
kuQXzoq2CibBmf4HL+USfl407x/KYfZO1FtxFotUED/YBIUfPlzV726/R1Uby/p+
GNJGCwG1MVUChQXhdOFIEyvMlte9328h8a75ytQK6GvRJK17y9M6ElcZWT17nxYZ
pEMiOJnz8mjEu13cy4aScTNI3Smzy2YeBKjNralHH2NBLJclRp4oaqdRMfkrqvFq
tGkNsERmT3W38rTAfSc8MxYIrBJGZfr29Xt6I1yXcKv0sEARjJNTrJDp1uv+HLOT
8uy2TfcwRzPR9gckth/k47K8FYkejnsWL0pQa4qsUQrKdx+gKjExPJ8xIk9ubVD+
BtEvHmTORccQJYjitZuFu3NHDQOi5Bs2wBBbFwrvyO2iOASsKnOuLFKofe2Pq6/b
bn5zfIOMd/ZTw2BbboTMsQvTe65/rIUxrCXv6zNsCiCd+mRWDp+XYp1NHF2egyVP
P4hpGmp/RNOAunEStR5ugcz/rlztcojzHAKp5OMCJFpvEt2q5KX/bLxc69fZyyk4
q0BVt8RHexE95oNG5/qWUHHNW8V9V6DDPyIRzD9CMeUGSW8zvTPr3e1cfio2VVII
3LqNJdWP0BWRlBWc0afDsNtV6hC4J01QlUoNZby3LpSY5XxscDk8kqii2AQpqnqn
Q8G7V93QAoUyiT5g3s288kPoA1cjAH++hq6qV5UTEz1VvZOL77ZFiE912AaqHXmG
zR7wPPEQC2Rq/pO+ti9ER43F8IeoC2elGGRnzzOI5+TWQbKlkqmJKQPcWCmYuvT8
/RJKhP4bxQVrK4fqjVuTBJUayPIj7Hcvp28vbSxelJZoIGyE6eZXp/9HnjwbcBtO
xygvIeuF/OrmD2sbE7AO5mYbjU/zisyr/X+X03see5CjD6zwr97S7sVNMKUT2cKh
tQOCio5Z/hRbTLUOlUg5Q8d9/YvQGrTR9jYYunXawieDc5ir3Bc6siqV99aeba/l
OjeIxJt1FFduI9YtCgMjDj7H2mLwFxNtjS7CeVdKVnLed7DFLYB1m6kYdR0tFR5n
67EsEkk0KAGs1ylYIXUp6Ru99Rsrka7UxfRjHfiBtTE8zGmOVNm8dP1QfKXogmoE
zkK8Hmcv9CyAvI2THnPcdpjIoUCDO0P3LAKJITvjlFD9SCqelzmnyIsPt0BJ7llf
tRCtRJ3trzNoZT+fjkVkWnShD/9b5Cf4ovucXIJoBIuoeRR7lrskblWb2GV/EGSy
vQTwmlbrPECQkqnJp5GoWeHU2DOy6DFahGOuAo/Mk0DX8V5QrPeUT9vvyYt0VUab
CF0yidM3iFPWExxHYMMJkX/LOIZXJQqlI7womq0htESQE7Ri1dAPVkfPezRlK6Jn
sw4/Zu9GK6SjQF+I1cTz6aTPY8DyeKkQ5tvFaMxxmiMbPRyKn/A+HoTyo6BKDz1r
zUoL/LOfsqHlVLejreZ1AcvFwfZOZD6lISOl8/sdyxiDsoGlaqm/XEtcC2xHmd0l
v5U0CzIcMRTzQhQejQxRKydNBm9TmUTlqdGI2XlCH1929qJSnd3r0WWhSGsKXLzt
uZzPRGZXTg9Qf88ySRGzvXLVl8APtRW/n4yt7hLw8WtJuws9iwSz5Gq3v7buM5bA
ilZh9LO0ggGlvR9vWS3svMO9jXJWEir0tY15YTd3VcUad0RoWZBImsfloYU5icKy
7j7eZc3rbGtwgMaa0PHeRS2wx2qdjTL+jBCBece/Szp8qMpkWVNXvRrMa4SeWEJT
LdFgdC17AZLfEr0uZoNsFWYgxyLF2tmCU2fmwwAj9J61CQHSog51pnjT7RSrSWvD
h37O8Yh2/NRwWxXgJ5ngf/RkZ+r0ZWQsz8PKoq1mvblzaI9i2+Rit9jY1OcCzx21
FM72gmnEUICTOPdAxhjD5JdnIHXGAJyl0LOOmiLcfS/pHZGhwco5U5j5FQUIzpw0
C/Ql2PRZD9ku1CovJ+tufcK9P4P4OIsXaoEhAQVWzkHzdDgmKmFkMFknlWPV9rI+
5r9ChOLZmdaggMvjIAOzwlmZJV17qUtA/BOsDmpChxQQuwaI38a94jQXTfSNeUQA
kLzIoFkzUJ/epJ18WHkjpKeek0ZnpN7pfU+Rqjm6JvZvnBa4pXUQrN8a/2XvLyh6
kuNyGmv8nqjzTKEGdF/wa6zP9rhP0e0j/aSAU2VMcmIW+S0M6Zt8r0zrdXTsFhpc
0909cyp4zcLMuBZl4SFQlm2ETGInGOzhmYXTg6pUCcTJfLhlOIQLJkOHy92GRjTG
VFx/XeFXJuuz3ovGD1gIkA/b71EuWhAGaOa/JCbeLPT+FFsIvDpAKJdIe70UCkK1
KlhtWcH96A/yeF2mX6LJ9M+iImCLZwIcy71q8Lw5fF6VFmHpwJW1dzGEBr7J3XE0
7FLD7nJtQwHwJxjOuJJFCz2fpZgtxI8DsSwHChy5M0i8dUd37rMQVSMubLFLweSn
N9mZsuDoBW5YD9YWJfyRm2/LLadnNCBPcNpiPXOjn66BYHC3jX1+ZjE6R0ZR8Lss
M9TOZaf902fGm8zqW9CB+b60kD1pnDWgMuEvbgcq+3dmx+T19lM+8iYR5yBZMplR
tV4V9IHnoXlk1W2ckHg1baHSARST/dsiBUNCZ8oHn8Xc5+74dDhiUsONc+abhmZN
LToTGG3YrIS38y/0XZCtRaYqL5T89yb28O2Ee3JRy4JT9227C7YUCn8ct8O6qdGS
gi68eclh78b8iwATkHhzdAxYq6RRSQGK/ZXqo45c8ucO/HQ6meVVpzDc0Tr92JEE
ItV0CxMGyEew4IFGU+/v1u2iPRXKRO6/O/2yF0L1DoFbIY6Q8ONxtJourFQHD8O+
0RBpw9WauBkdpkRs+cFU9peotOeTF/WNYSNvdXp73bbZ18ajOfuc+y9dso6Ric5L
sacpiPsz4ceJf+0UZouvWH9l+mJUcZAafv1oK1TiuYb3eEvfT6zHhztdHcm2VALE
Eh6v30N8WPtJbBky4VDZTQKw01MN4c/vd8XmDtl8Qg0G8VUfDebcaoOcst0oqUSS
CNurk+imUPslxSpkFXETNuXQGo8Sb7mypmW+OaHLIugyd4bTwxee+LCDUYfWyEgY
wvJ64pV4uLcqeXiF74/aM7hUI5p9B0V9ZkYNVZQzhMaKUeVVJkrCxBj98TbZgvE3
mW+bdTPBXYw4k8XzunXp2URHsIBv/2MeIJc5msTUCvx9mGaqY0np7FEA13rfSm39
LxDlK+joYdkftzXpckn8hJWpEzsfPeLV6lg0IL6Gn6cx/+mAqbS+Hno5LhDTcJqZ
W+ri2F2n1OgCu8LPK3zwr6Oh8+HXfTXu174lKoXzDnlGqOTI44+e+1RS6PWpTkDo
841e56sVCVxfNO3cpWbrBgGLZEWm3P4u5v6L1/m7rvQzpdBjIaSQZ0uzKGCVUqP/
zw60TA4CD4nsbCR+RDgGZejOk1YZ5gsEuPTXBI/1Smkg+x/OdD60IbYJD6UZZLk2
YRp1W4j0fQYGYRQyrGnN/5bVZ0u7uLWAjuXZWJev6cAl/HQsMmTGDvrnmRuGouXE
IDzMGATeJt5zgkr9tHeKMNeN4NkLVY33s9Gj8hQZZvqeDH2qsMeqtUFzvFkPtTlj
clgkSdxuQ1yCtg81G2d7L6UIJZSffPascEt3Se7wzXnq2Vx717PzgrgE9jD1Lc8C
vjy7ByLjQzg3RpzQ7Muji1KcvBekiHXQGyvOx1EPwK5CuxdXa+XL7vKtA00If7jY
R8E/6rFCXhYOjEZ82rb8OVr3rh5/YzQEWPlc3jICuXaxy2C9vR98x2Ar/DrHjfwS
v0+XfK2PISFK+WPCp9otmlq1z8dyCootQaJWMnCnvSiiPhIdupTulhQlWIL5MKRg
nhTbBiS8Da0q9yGgn63mG33RZ4uTBKeIfJE0t4oV7dDMJ8ERRhy7o0odpUhdUjWf
EBWC3nj8QlbpYEzX6zpHt2+LB5hTG6tiDkxzFW8gBNLMjxXmEGjYosjN2BuyDFCR
1/gPBNfbKPj0WUqO9RwdAheyIxquFnNOg+L7Wy68JjfHZaJdi5GBUeooRW/sDm26
n2+/rPDkuP+pmebLC1Uf+LmQcR+NFqk7TgxSWdEybMs4hDXcCWFk2ZXmixW/+har
BnQvlJrUN4MXzLUmhyd7ppN7KVUvYUQSiheDPp1gPX6sCTbwLvfJwfaGDshbuxPf
WsCWa/L9TfcuIbXqLnvacqRGkkh52jCCN7sbc59vd29loBX4yodNbFO9Xdb/VL/z
gUGkQH3QuoGCBaqO8upU/uytvtqY7M0RtVpqlxID5dwrRnXD7cmbV8L/JqxIrxpE
kYSm/DWSer8LJJLMnGsz+GBJBd6bngBjf/TmpBTLoBNKEClNLXw+eU1CqbVjNnn5
Gg8k7HP/5CQcnFXOhIcHmYis2uXTett/zxpPRTYMtZVnE21mXE+bmjv+855YQFTC
HiCPnJA9XdySAfskxpzr7yimLqVEFVteuQMM9EMejmTDRdPt/h4HdKsF7SSCAssJ
i8ndwBhlumVWIn5368na1JUaCbNv8SXxdFZToNQjLbNoH6AuO/eLVug6G6hCFnKL
/c17O4/gp/Z6CCtviCcWC1OmRVTENSrPL9V7j+3oak46ktaMM48lFcnsMkNAySjt
GIVR5SowWQqLUV9O+DVatLeWkV6HYatmzxxsDAZiboz7iZUmbo3EPIPj01a72WHJ
+K7U4t4DjofBFshhR4pvJh52GsrFypoO7RJO/JttjJs2AZf6518gyCS2J3JjtPqf
3ajph3x95hDxZ1aHNCe9882RyY0QXWruwWx3Xx9Ulb3I7GQIgZUL0/DXDpzy7cIM
HiDRlQ1gHUArRQRUIlo1jWM6N6X+5YRYrUqdUdxf4CaDnx+Z86mVxmpCREZEp2vz
Kh8tmqR+dk8F0hkYOTxcDO8PVoz3m4bOqekfsKW48kB+H7EFYwNSOHxYnmQe5Q8B
xI4zR72fwh4oQpqKJtThDfEJeLqLHNUj6VhIXNyAiYkGmZo+HIXnLFMztlig3pdt
hLmbXKTbbadKRXjXo0P+K9IB7veC5FYlgZxJ6e95MTaW0/QUpU34hWtREvNgERJA
9ndSSSlrZxx9Cxrk3UY6npVvlJwU1QfB2JKEcjki1ita3q+49kVDL+C2SWwvL1hH
2d96gmBUsruONRg2VfrPIADuz35saK3/TI9QOKRkFVRYuntYAkdrKFatyswHdQ5n
YHbshxDjvCCkptK3+Rk+Troz5uYAb9kYoLC1DuYkUFMJhl1NaAt6EGv3ZVyr0eDl
CHr4ueyMy5qghIBNg9UYBoU7FX/Q0sDOMaHub140q7yHNzvjSnOPKRa2Cx5Q9yuB
pOYoYofdsnt6HdBEVnwWMA39AF6O3XB7ZmHbO0/6veN0AfcfktH8CxZ1MtaYGWzi
0crnLNLB71QJ5KNH0/UKIxqAx2AYpAGUxjSTV3auaqWHUhb/qFy7Rb1BKl/XzKpH
6szq6DbPzM672ZFKgBjOrmzULf0Ekoc4c0zo2ucWfVn2XgS2Z1Brx1IEmhlH6Y97
yl+8GBIcQx65DH65ujhF1g9cqTo33GIp0t5XUeIWZ0euBHvOJsBuAAmxDBoZO4bj
JOTDWWzVW5Ghg7GgEPDMRnpzS5iXE08ogbFgYf8kVP2bEGMuZcKnUDsQMZQAER+3
Yt1538wQdPnB6xwK03Ocj/NTWEon5zE2/0iZq+9h5G5WVefQQwYLNVhzEuvCVjw2
P9dZ8iesv6vw7HLtRlhf14lM8W/i4RVt0pCCF3YJrM9tWky0mM0xVNIMeEGv5dVn
Z7E4xhVGBjN1Ders3vDQbGbk705lbBuf4PFDnW4xj0hsovG1fGBJIQxQYi927T63
TCvviIP0BJBB/ezAjwcIOFlWlLNIf3f1rCptDHQXD/NvuTB0MKdvynOfOMDxRRMu
C0BgxOurnVQAl5Mt+qRCHvV97lYQ22y5j/H6dBwpgjKKOi4XJFkmlIzeFUKGQIQg
iK5/5HLlBxuVMpd0ZaGZXMAgRnsV57ZqBNmXaG5iWN/7yTxk/kMt+dl4VfbM7pMa
ohziGJbNS+e6Y2K+NY97P5kvUT/inBHQPT42RBhl9MZIcANsO74BIPTVDVfniHDd
jfC5xfVsudnVG/UytphXzmp8d4tTCN+dJTkG3/sMjD4j77ZWVIueR/munkRiEV2Z
4wsf55weMqh0LEwiEwztGevCdHtRLZ1z/v8tkxgsPA+2ZVRFRvQ7rZLOE5e1+pcK
MOO8gtAGrXUCXIQNLzSp+w9UD4LvnpAkv7Bx3HXmeeFFaeAxkD//9prGadgGKsxv
5zE4pa1FKM5D+XbWNg7JtRiMNSEVA1oddf2F8Tn2T117a8ThcOxVMDITXP0Sdkeb
wFdyMmhYXcdi1OFm6nk5XiZBEYTSrIvJl5QorTOV/egX4TPzxWKi4XREgM2Y29if
IUqXnB2j6Hi+NAUqndXW0sM44Dh83bx28foQi+n/ggJXfoiObk3B8va24LxwClM+
LlOef9BpDnHpDXhpiyZajldsyWcgchA2RmBwjGDcYGeRfseUzYhvCMdoSZnGRXy6
FdmyeJkMSzRWGIy6VHgHkq/pmWPKnQ3U4mKo9/0vHvpF8dSui+BYAydAaC+LMgSE
xGqkgB022gt0X/Zr1yaZOKfeq7z/jKgzjrDR276Op/JlHPW25ytksNkNDr7Au+LI
mgnrtoEa6s2xJr2Jpq4QSbeuMNpjiY+ODW1rzXnuSXjsLRg48f6BGbyA6WbGrEzm
rxPysInKN2UT9MeE/X+FXw0+Lvh5SjqRF+8FC59aZoVblGC2O9nF6ExfEDkFeBhZ
6hzYa3faOJf9BwjRBZDrnqmvrlB3wwU9Gk6CvyYypiE1uhPL7adsLRgR5I096EPL
aZGgfMVC4Ii6VO+kBMta0XXJ4bX0xm/zADwOuccUa2z6JMlb52brnB/q7ErjEbxS
Ju/lCxHL4L6mPy4kwZNeH7RYdpGf3VXPGvpx8VR4GtRESLDkdkMdVkk8C1GoTGow
1CB9qKaBknwACwozKZ6foff4m49fnkVm1IpcXS+UburUsmHB2tYK8hc4nEj1HrN3
ygqTKnL9Hayd5NZbmruPXpFbUj1PA0fAQ5ivWNI5y3upCTTJljZM/bAt3zGq+nMV
SZ5aIvDSIQ3vhh0nstGkH6tLmdoR6klDaU+8u8FNkLOsn24WIRqOZ0y2I0ZkvSM7
SCnfECQMuu+aLrm3Qb+UWolfItkDLN0r7OQZx9CrSWF3MWHtMeasRq8bc760hXOT
wTqYeBGpxSdL6NFUAlhwsNXB18ogYoMcw6eujchlsOZmHyiMHjwuSGOmZHjbGbGR
uE+WQRO6Se1+wpcotGuXM2KwTz8yeH7xm9CtUDyYGESCfGX+pFWwm9SYgZ5CS2Wa
Eove/3JcQ+lSqlgH9uK9HlfRrexEsbE3dBRO58iBvTM/dr30qZrBuSpQ9Gv0ZaYA
gmZ8I6YZcDiTqV5fzBJrFBXU8a7/Ac/c4eywHxT/m/FNWuZi1HMpwXUrhxAWY5zl
FwY9CeNPAKR+Oexa8RKI4/vZPOaR8AuxM5nu0dk4rv/E6N2fXK90CXdR5d8sp85v
bNC2F41Zblj4XvvBEYFhAHiuSddUPEu4PATV93LIfycVAo8RIgm24BVFGguZB6AB
q2G5FpPsjqtHnoundgA+JAg0RrbwKZ/9jqAmZWubaGjYWU6njs+thPxXap6jy7+D
E5si/gQRprEYdMCDmyGO5JXkP8pai6zQdm9dbyrcXb8Vj1h0wZm3b1Qrr7LDq5LB
c9cDLAG0feqmb6Vwk7RfT9kDtAxcRij3/vepTNnh9b84q+dS48snESVD8AZIGWk0
i3kUODMA3A4Q4sISchZ6NEckaKWNbnIbu3zgzLBHCMvydOwWloZkn85TFHRgT5Zr
rmp4zLwdIjVl2Cxl7M2jPr1qGHP3r5/vD+0mfHGu5DdDR4MewVgzlx3NjdstgvJ6
zw5q85owKnpD/NaeD3mjznYSqfDvSNqs7QRZbvlH2+xmXJDm7pE4CFTyh4RSUcgr
6z1Nwaj7P9BxGHrd1VtDBwVuAwcu0i7FNDgYTOMYAG3cZ2CZdU1HEfrDc7Z0cULJ
DVUgE4OKPDQcJi7JQE9bJKsLOeJAwuP2pU5E81sA1VaMOr9u53V7ZUxVLd9ENJvQ
LWOXmWJDH3sukjM+3K1+4lLtYZXLGn2iNrYtN+LfUCn7GGZ7D/kkouOnXsewrsr3
MJYithj+WwT1wdV6P5Kqr5PalinGCN+6f/a6WM4K2sWFaoiG7G92NEeyX1bVUOxq
C2lCH3jz5s8SglZ9NCY4siuY8uWFpCz7J+u17FpXE2m78ddPrwajBHQW3xw7H7jn
bSHsNIDEccddKLQMZDii/D8upO9iCy8bTfdHAJbHSaU7jce+zCE4UUsLc+q2vfjR
3j+xloUubSM8f45oQUTOE8qivziXG8wgGIdVC8KGh7mhVu3WCyTZw1zYxiTB8yV5
7gDvc0xhG24BIVLhY2xa7t1j14HZuB69RU0B2Es7uvlY+R07r0q3YCuJyw3awNQ+
CZc36XgENJqUI8sMnnNG5lnmzvfX5X4FrY+p3gCAT6vODIXL1ONIKmm2DNuTMqhU
UZ2GYjH7Z5fklkPKJbzBRqRyGpXQ5auqwvxoD+U2R2mWD1hfQt28woCB4XdEI0UI
tilhkCuUCYwLr06xLdPfykwg8OaHzUHCjUiRHyxuuq5VsrRTkv7mbICYI6wqMZkf
UZxNKGjsiDeZ8jZqoHPszsgS058SbIVFJRLdswqivz5iTadquwBGl4Wr45fA2CcS
awQL0+QlTPbIyU6HMtoxkKTJVYg9Pfx0TDYWsoIsQmV8k91+MIodPaoQO8izQw5N
5HX6NTn/OHBLBA4I2ov2Pk9M9wSLrMaDzIyQBaUEuY7lnKeKciaGBXwE/aKmgBVP
s5j7TPg+XKKwu5zTcvyw4IleNSImxzt396Zflp+xPZWaEY4+dBmq/12RgTc9ev8E
ZbROtgW1WndLv3iPbNRQau0eS/QG8ofCfjS6dZ6MJlqlTY1ppH2Lzpe32hTnP7VG
LDF0FPnJ2EQqRLaUIVeTjcIUK9zTucHxVzsaj94JxyAl82p2b6ukJF+/lfbaB2rc
SuTy5RGnH0jgkhrohVyRauVHd9K9u96TEAALeVewgwP1nDCMs9lsgjCYlj42tqm6
EGbjIILgZl1CdYkgkGnxksCNGT4C3f4E9InIdqFvOKrn9VnoBxgnWQ18q7Y+TWAI
WfzZwcuS5sFFZzp2F9uLeHdnEWW5ca06A89vmrG5o/oQmsFFiHIDaiHvnFz3FUg5
38NQxJtnUDHbyD6ARIVd8zuokY6IQEFRLt+F7CjF9ZtkA1145EIEC3MSx3pA7Sdt
uvmrfdTYFhAlKyps29yEzb4I9WYHcCpHEuEyTgxADmSaTcRxymoQ7J0a4InGDVzM
p9znJieaHS/cT9w+SWrVSsg/nvpO8pKkU8N8Ur8qGOI7ajidseSqrg7fx8S5XNGm
XeiAC0N4oYVptiU8/+Tx7LL71bz5K1RheUgWjCeNb7JKYGCE/vb5kNyJD1LPvJHO
LNsaTqGKgxX43F3L2HAX3JfeNBnx5It64gxmmvlIJtE5FcCgsCNNkIoHdKA1Kj41
emNgj+b8mYbtSe3FMFtZH0+1iy5xrpuh3TR9g7QnwrmOQTGcOG3mXvt0vLnOPdjK
hBHfrTVNh4YzlCowaMh4fiR5oOMHx1nXUSkUnNTV1rIhZlwPEFDFjNR7wLSP+P+7
tcA+M/oMxsiRLbedgq6F+Ji01RFvARJnoJDhhlrldYK3N2IaDg3eZuA4iZz1nYSn
4WR6+DuqQnx3rXcDuEWxNO2RLu8G//fBSyjDuS5bdxhMR1OlOpChQZ35Eo2psVrz
/Zf5f53fSkLSah09euOgoyWaDT0b7YhQec2dZtxy5HiM8QPjCFHma1nVIlOihfrV
qnnICkIAwSW/mRUj3OaOYEdDzE08m9zKQPgnl7zfhm9eIJktN7n5WSioe4mns1ap
GVd1P09DKaHUB44Mpd35bE+kEDAm8GId2IE35nr1ED/h1FuAzst3vh+iR8wmmzSK
WOAWzX7eFARH8Z9LPG++ShJWltGZmyvoW8V8Knf4Glf9sKkU/WOADHpLPm8ZZ8rg
NFbAYXsL7UYIk0pJa7/f04lT2cxkXAtnzdKdJYPMXPrHJZ2hmuVnWcLmTUzBqDeZ
jVuvd/5aJsD5hCiejwRE4q1p31+Anqdsi3LZ0eKKAMQK1UvHlVCMf6w7ENzh876j
jtfsyQJRSMWTuCVNzwI34C+feC2H2IawYXsdw0LIppmPz9ONuwgDX1RrqjyyQ9q5
CR8Rr3BU0N1ufD7riMT/ysVPez4cjs0P55wEqHhtFejTmSujht3GtEK3OQ9IvOMW
tZVJhcyUTf5/V+bZ0Dr4DjiIqW1pTEXK3ynsDpdEikNsKZ7Ny7MWpCxy4A5ZDwlx
BKe1iz5hgerDylkQYztEhMOMGOLarwEaW6GvU9p3nT/8QnkPh5we2IgFtSGRyHYz
ly1gvdGXE5jXrfzPxvvn3fTAnI42pKSisnwR4hOQ1vvWgy7PgWQmePYRyTo/CRVE
FscuUFk+5UHtmAj7jxhpAuXKmckgIDxru0/HY2oe8bOeIJ+uZ2JKOufKl4LGJHgb
DG2N+O1t+BUPjaEnkIUKF6szAhz2bowjcAmWFiFgHSsdYpjWFfyhHRyty7yaJoDh
bCMNR9dxEc+igqBIL9//QtP3pbK6fkQymi1K8ySE9qyNd8zVS1lHFfCY7d+mBuoF
m0q2M+FzqwXGGh9NHUQS3jOizLIpZtoLEOuz2JzIlzmP3GEnzAqnrWYaoC2MdgQX
NEsKZ95wHV3tg7ErctWHaz2bVHcCuAKVs5ZC7F4NEO6E5Nas3Hni7rf5wCJr3sNk
lbhtCFa+4xovQ1L5jJFFeQ/r9ieSiot2Ytrql2QJIPZ20lpna4tdl4h3B1251RZK
uKp7PX86XFct9akWVhaVYjzI+xzzR41JzW2WGNlG5RUzEG68Wmbd0nm9nqZULvz/
U8l9fL4bzUQ3sOf1TZBgj9xnCYaYCfLaJ7/Om8t2Q0tU4NY+BWJtjwMTrQ/I0Wvh
MQtMpA/elmWwurEHpCQ4DX7Ovwb33uSY5J88+fdoN20xPrsCldZ95qUO3hfAMpXS
J/jvgIv3wuMObFN87iz0qQU4aNm7HmkkccYSAO4OlgZXQcmE27c4vaE/d+nWGY5p
x56DYpovHwXQ2eFwlIUZCsT3HrRLNkKqG/kIUcL+pRnDAXTeJF0/CVGlSVnpKdSY
0BjUn1lEXKDp9DCnJEtYi0U/cIrBxtF91B5gIZcelLAtspyTxU1NGbI5i0HswNEM
dy9/effllo6EaOyL6sTwJqaQqCFlpAg0HXnFdiX6gq65yOyZEmKHsEAeUY6w7q0Y
1WeUf6wyoP9iRUuoWsMPOzCAXU0AlSeKDrwpVtQ2LYQvegUCJiV4AkItRa6EvlRR
FMMJUOMGuRv01yssCxHLO+07CujdHz1AtEUf+gxl3wjpU5MHnoIz4+sCELzcCtNE
KScbtMAzm/tYkpphyYZBbZs8GxOWVb/bPUmDWFsHOaIzJkK96HRw96ZWaTimglb4
gMMWq8H03FDJ6zWHcmiXpgVC9lrj+ASac8BURBmRE2f8+ytzukrtEZwixi27Ewv3
eEjTmTKz9EqwZvKIauE1mvCN6/hRILxBBtArG3RoPTzWHnUus+dercUP2jicrwQZ
MhtLTHk3Ce5qaZyKjWvHQ5PDM52DV3lz7H2Jd9Bch0OOyL9rGEWuU2nVIDOL7HFI
mbAKv1rrDiRS6ro6jFnKSPes6QrDrjF5NoIjv91QoIKVow2TH4VGr+fqthbQTxnJ
6lO9dBjbFpU9BA0p+4owRAnjJZaXg9DekJkLQKnhl/mc+71n1xQ/wypSPKLi4FRG
UHNhykky1SMImzZXdk0G5H54Ga5lirlsbyqxgLPOES1m71OapvUbnDxzIaI/Ubhf
COtcx5SYr7uI9JiTS8izvMQ0e8UaWFqzvdrzn7t+d38HVJU3gpNEvG8yDVEzRIOw
WT2WxT8pMhuItnhlSIQOe8VN4NLQyKGndpNNcGuChK/SikUMm3ZbdmYSJYeVlin4
lAwoF8aFePKCm7Bbr4rKN48fYgYWg5TEEOeWjMdyJo4up4cjoF8vQXwOIt6FPSfs
mJVQCqNBZ1/Wh27ChDssgc+myteKxbNpSmsJe/kE4N7jZ1F0bizD44R5NNy2pl/H
eUvfrdwbOQ0GSllG81UQh69C0+X7JPwDifUhfHrpPERLRM/XrMoI6o0dJx9aarqp
CLjK0BduH66VQ5AXphWkyay5wJx19phDMEJme/LVwFdfEK3vl3ghM52tAlZVgXN2
DQ5w542ohBQDwTcJanvDF3MvZHn+4L5UFafxxarFkRG0zeCA16H2qowpp83PNd/P
vxpbJIdSjBUGmThRVho/qiGtyfGZd6xedvce66E+nnX2VhbOs7gOghO3p0ngE5MH
9JaV/xRqCJqxqbP2WehcvGUN5WiCeej4yuZM0ksKYJ92Umc4KmxqPTS+wTlMsxpy
bMT70oY/Ku6jlSYSEl+OziGRelRfuOwKtEMW0BYEr+IfvbHClqlwOC4GlGb3AkG3
k4RmclZbcB3VfRpAQCdLMgltxJsPNspoppB5C/KpAWW3g0Q5/sL1v59lNEing1I+
E3qOt7jj5S0mdJ5mBro6kxvc0Pz7O2DMzwTRAurCMb5a+m2dXt+TzK/4yIIxuLPP
AR7SOdcwj9p22N4GNQoZz/aigs4dNloobVoTIOWcm04NYpbMHuwIGjq+Ai921INj
cXu/6fTnGpCaExFa1E4AkqA7IYX3xkj11FV4ADvthuDmNQ0wpMM9ICoDT7O5cXBV
o/uU0cMwQXHpln4cCcT5r4Hr1afeqhm+PGzFZrl+De1bpW+La5D0wnTGsmhjDinD
LkLGZ3bKm1rnB3Ihdhf0xELE8eHglASN18QFjeuVAAV/Cx2DzoeE0e5PTVTfpGdy
NCHytJ4msG3VK/PX9D50lKQ4pbdl5wWEexdWTXJzL4332+b9mIv0XR1Y9iPNaHxk
qt5Z3ww9HkQk1Wh3Kmu9sNYJC3dZ+TWDDC3ZWUiktHXREKbhnVRiHsJXspFqkONR
cmgMkFRRNdOmZZU4mcIGwIe8BepWSxzs0E744SYQ6CXCxcL05wWTSsnpY9sVHDJC
vklkdDzyk+meNIHaU8zhVRld1WrJJ/Pj2rE4uUaglsDZB10Wqfsl5XxqqIei4QBc
uD5SSdWkgB9hA1rufwgAmr5BTRPR2NBFgEhc3R/DKIU8D/Gt2meENKwsSq8uCjpa
ETPNZvQlk7Qk3buJu8r0UK18PMcd1l/+fcigHlH2dZNNNaJZbsoWAD9i/Yt3Qzd1
UGuFrCsVaY66N0Y/6opE9OIoszZ75MqVdHz6Kou+qlQcswlwdRSzviItnk+MhRUs
2dJEbOGiYuKn7KaoBgzmK3nXQr9zM2dfeSpHpqjzkcak4RfJJpucD90CLzkUbFJT
1Ccvm3hDsyOjGmTDfUf/le8fhDecSykQ2t8vPIKs87XiqKOZr8c2DjyDwnN6a4Y3
zggUxYDUT0UjUTz1R6W1JAYvWrvwXYuJvp1NGybt/yAUO9ZKbuEGFup7U39foFKX
3wlK+neZuDBWXUm4i04UbpRdoMjN3/++zs4FEEoDyq0tarz6+OVJ6HReLqjViIFK
KD1BMPaI6If6A3mAaAftgcPwWpMBDH2w94MvbgNWyu9m+7XzsG32gR1VrpT1Y5Nx
V4UtVpn3h+YL/Iu5AP86riZefGVy4dMGqHaqlde78+CUyxugy7M5dEBhvxukb+pc
F2hg3hlSRSet9pmDIYPYHmuXrQ+tV1OKf30v5r86722e1ZLSck24LJ6xZb+wpdD/
/oGC4os3ZhJ5ZSbpOSNcthwEBaGqq+S3dSDqBnBIhIjuGGK0rsSDwHw9/21stWMG
FOqu7qILwuX+CSJL/JjX+YFfJpO4L2H1pDcWBJ1K5BXvVSsfUMqXgSNSBan78aCD
k6E6K5z+KA3HI91qGztbjDaSt7azqorewkolkW7shs9RiSkNMjb9nppstbgzibb8
DymINWc0pKYFz0eJEjynhNKqXPunFd8OrbRsTMRxslKJ8CzR/OUYiTeRLn5W9K7o
GoC2AlotKU14TAG6FO5gjqSAmiO+UOGysb3j6ljpGd74uuQolG07ATX5tPHPfZRj
c10YFleTut86R9h5ACiGXBAO3mHbrYqsSbq+sUNlKfH2PsQD2/oo+SFHb/XVwB0K
CTKaa0g5rgUEvNK0yf7TTL4hB9rUKNoDdXIBBo6j6j5hlE07rcWjsqPe73lhXSDV
44Sy0tU4PwN3mh1bKOOEZ0SF+eqzMTjJ6w16yCOJv7/MDsBPtZ9GXD6iziyYcxUn
rz53McIRMeNsUZlJx0yar7he8iYSn9nL9955kkZ7SVQUbRC7WxSu0P23d4wqGDiS
9H1ZmL9spEiWl0Gd8GNIiON69tIoMYVQlJa1H/LNd1G2QDPx7DEmfaa6/An8oPB3
jOK6l2LU04G8JeRAVKaGEm1WNSf0vjgka8vrH8JYHyg6J3rTCLZof6a1xv+5uHN/
V+VbfPMkgvNaBjLVoXxbxBDwpeNDs8OPywcufTWuRFRfSFaK+UMjh5stYYCiiItR
SifJj+N8siWfLeSbug+pQZFv9GdtoCrylTiMTgxOHTurh4oYhfGKDFZ/f4JltFuG
iKZzwdTO6zaMn/xtVDAKLqFpA6pmRAwIzsGZOZSjjALvQGSZlALsJ0uGBV7c64EJ
eOjU+9EmI9Xbh33X9yTw0NM9FArnM5yWm7g6h6RoBbVrWSOmbgRKh0K9RqtrmZ8m
l4kfuZTQezniiQG3BrtdO4Q2tz1OpL4R82RXZjoX5yU9XtBlrTOw6BZdMB7Y57nD
UnZ43Xj5BET/FC7El9A999jKasVgvq3ZRftrZEm8es1eZVym4LGa11+W/Jsl5gDk
xJuopF7H/CPlYpJseUj8YMxU9vO3YCt//3OTLQxdzY663scUP+PQgPP0fd81Rv6n
TzhW+VwxKxlMiNbcdNj9q8oK2RfCnb1SMhlk90yPjJpLE7cA+OSTCsPJmhd8cJ8v
FnYSW1SOmSVmlsFiBsDvkfquOmwWEqQwZ7Sv9/oknlo9GyzZwuBohiEdR76+3WGN
Ve6ZM+xcJT/l7LwMHr0hA/aQjalcwV7peFuqtddgSX7HZKtSQl2YDZeNOXxZFQ/D
PCguVYhe4LozQFFKfqvFis8a++KXWRotDhRIEgnr1hH0Q/w5Al8vqxgqQqRaPHbQ
+JiW+CuxfLu8b1MU4sH5EPCRV7EHOXAmZgMUTGGu+K9Fx4+yhn0I75gq1W4KgnZa
wkHuth9l1yicAAZcOY9DJJ9KT3OvuoWRppyd5qIEHnsaPVjpHP1dxslNqaXd0ooV
nA2Zm/1QEEfxO4vlc+QBmWssPDs7O1JPEiR638bP1Ue/SpOwazRZvvMT4Vz6V4Px
wdFIz6/LdOkzLRo+3y59eOXaFIHxBneMjwubHxcD/55JEOzWHD6RMoa2JDVrugXj
OnXTBFGvr8pS7QzdP98PnWCECJNqrYbf9vbl/yFkBnIgif815ap5Za1U63BkMbHa
jCPs803COaU3qPQLpHNR6v7xjRvBLmWiHxan1I/sAPyfNRqP0xyiRA3jRQqFhyq0
8lNVCY00G79Jw2DTCUcCtzJr5EJJ7QYs3dkujJM46We2+CLeV2tZni4g6BmqO473
YVAY4/lvPorrJLdHpYukcYXodQD7awllkcQE1mUioa5T+pnTkaMLuhFo5JHT76WZ
ArTrCUl9cHl7Ba6rVOUqc4qrUZ15T62XW8HW/QnN4t+r1mpELs6vh2zNvH0YOeFQ
nJbCldkcJS1KFCjX2CuxOpJPAiKbB2lTrRzdRbWoNUCCJdCpC8Khp+qSv1VwoiCd
eWvp4Ci8+c/lqXM6kWzG46wK/flcZvza7vbgqA2A4f1XdG69K0AI4QIhIC7Q37cv
2VaDmqrYBVuecqSrdvGv9L/2vRX8HUJtVU7df2h5MNGF551GFr1JR/kEO+V0F2En
yZNDTj4jw/KDHa6h7ZdnXL6du44E/c2T8lwFlTqQW52NAcE5RAtdLwUS96bHUh4H
iu5xzxpKk6037wmCLhTlxjXVed4vEE/ij582GbyiUdI28BMN2KOe7eYtnvhAuypK
D5+CZD5OwCId5a4QJPxng/vbCrRJRQtcnsYd5YrI0CubQKOQungdQJOKann5Lx30
zUJ4ciHEkKPZFu+NTxTtYgVULdwNloA7GPTpyJUUAGXvUIeFzqbps2/bCyr8MUBZ
DrT3TRKq48rlPFWuPf1v1FqoYv3E/H2+pE7g/6+VlbA/lLbbP/SS3XUdDxK5bTlB
vB2jW4tyvXbpXUm9wl1zb8ZLZcEvjVSI966oafmMbYrwZnra4dIfUBSDT9d0UTvq
bmh13DYFPeu9UkrbGNi2cg5IN6bg0aoYkr3rDOmSQKze3q8ShNYT7DnO6FVcqN5j
ntu75HYRhYDJbmrleyyi+6jd2xP4/hictlkyJRAnEqF8FUgBpBXMZZeNJSsXy7P4
InprQBGGB1ReiRpEyymUQVFuWZNLlpLfz1nyrFAUlhCKq1noMx8zA4Rq3YFscqZH
Bv/BdUfCEHQ8cY/4r24SYhKjxSs4tjl9nwKej3h2GC+ITZXx2lME11lqJ/Os5yoH
np6s5WWYpQnodELsE2wUh7QQ5Sw/V4FI/RlWL4WRcGmFdOQ8yFChgKTJ02BPqZQa
pWmq2W7n6VlnQpaAT3zwMt+U9U6Y0q8ncZtDmS5KVmy/LRdBL2XXjjTruNOmoyJR
mz/3w8tDI2CB+xv9carZwd5rqEwRx9QXkm5EnWu4Zly2sfqMzJrCwtXHbfeEFH+l
X7GiGKGB34zra1wfCBlu67A/CNCRrLra24fXrnSDkJfXcNofHw4UQcMJiPbcDcVs
rQecEn7xoH2zCklJ0DHEbrWnFtK40T/saTGvg3EeOgdcjJlLpsPBdyQ4dla6/UUa
10kv3jlHq54pSdHpg3Mb3UX3spUz1+ravXqTxIjnE/Lp9r3dUGy+tqg3pcZJfguK
onHxkHvQhkHV6J4ItAyrZ+qPzW10YJP/B7vQApk5l6+1geQwabg8FlEDFC0sPBuO
LDr0woJWjEArDM1MDnlVnqrv8TllNiy8vzlEmpZb5mU39Tq8ruAk8f7/+HXldYdY
1LrDnyzORlVkV3S6/QXOgwW/O6z1vlLk3qazbWbdx3dtEPPf/pKm6/HufxLo4+d1
P2H8TThvEUxgjkItu5bOPQRlhfX4CrdDm+L+MFXPjbBNBnbEMbp/uFjR91EEjE31
4ClAJaFputNqDCm4Dh+NhRKOshq2KZUoqhpq5a0BoNnWCY6gVunxnOURThCeQQIL
Lmqqo74kmiHQWxwVAaJwBht3SsfoLMFASNPX7R2KUZCxKP9+gR2hs58JOox/JANe
SCDnv1gEtI+MTbv9uaZVhULHIRG2my3LSYYwoHV3163m9iCc3tmDkQIbAYU+EY9P
/ziV5E8Pu+IFzIGVw2iYXhNOf2Sj/tQIpnNN4YkQH6KfmTSEUSGhU42yAKhEs61T
kTztdPaa0IaTam3pkhf3pItXlcGDEDd2ol3E7AOKz4SRgL0+v2X2rSkTcXS1xurO
5PlQjEA8Vy0B7fnc8xvLa8v6hFt1Qbad0k0wi+Tq0QYMMBXqnNqgEbQphbZBPhkO
wbqKDunw0FmXpTQ4qAq4D6RLOO7zoDGz4G1hgQV4+FMZbb+3Zy5ZtmDaSY82kiub
UD+59oCNLQbI/pG70U97546bygJh6/by4FhhUsbBkZAJ7NIVvDU09sA9g5mdUvFj
rYdls0wfp40FcdOcJ+ljXam+m8S40ScnFVuPryXvT5rbN0JUGq960SlzSswtAlQh
b0QXJUJIOtGbJi+JK2UJI5EFaBPFSQ0PTOG9r7bEorz9KKFOyPTZGjO7wWHHBaM2
g6kMRYjINslJw89HSTcl0ZLuiyox7OJPhDvbRUoB6evyQ9tfwr76A/Z4q+/mS4nO
DsPmoGqZ1XmL6kw4t6bD+insg+yq6EoCefZ7VhHuHsn1NXNpWLYrqrhQy14sRplu
BNnpnDoiVCFym9gudir1LV3tgjtUMoeLrFVpnImf41JAynCsNEzF+M6Impk16TJT
0KO+M9QXfYgW+YHvLvYuE102LL6u+T2x5BUTNHcKaHMb3WYzpaXN3IzVTiCGPoGj
K/xu9tIiJyiY/iu6UdCLJwek3I9B+lk52Gb1pJRW96Ul0gqoCotny5ofmyMTW4v/
/U76+F53KuijDZbe5h+ycvhtwrUuXg3g9w86Qb2lDUQ0ILtpT2y/dEpJACJDRMDb
94cNvZo32pZ9SPLodC5Vrr8LrFHPrgdS15+YJr6GYVC4EjIoPMVAaODmJ9Cqaq0j
amvO4tYK0sa3p1UrdZGQinL95TPlKeL+oeumKDfLN7U0CaVFkOCANugAd2SSQiIo
iV4FEhSiK7pw0mrs83/iK9zcBHgR3GPRlZagMoqqXfeBLfJloUMT8t1snD7f/NSH
GkaEmh4JpVU85LMoR/l9I59edAML46pooOeHCiLIxvH5djmD8tcIfyEtgFAAekv0
g+czDQui61/2++OC9imzlAShs3psnJ44l8/G1CIRz0VAanSfU1OXFu0xCH9bL2dU
kUVdLJVl0hj8pipJiXL6L3JR8Y14ChuUaOQJMVbUHmVay+epiHRi5IKisZwSJy57
vMGiQ4o07NpmV0G+ZWCmu6XXyPE4TP87eBTtLJOqGZyEmGdRsEPPs+GhVKtrsvnv
PgGrDbo8XRyY1jVzPZ+7+WgpQYfA8TrEotQctqD/h9UpgRoo5OyolgDEsTg5TXaO
Z6uP6fzDoQEw2Zu/bkkx2yucr7EwU6S6Y33XX8hDpqVTzYGmuzNot3pBEfKV7Vuz
CFVA12+69BaDp0ESF82Qv1huMnbNOJEUSGqjTZU/c07wPqX7fafv4tPVRZmOavoe
1ZuPubW2dD1Dm5xJ8GR6SPYn889leoUgZTbsriJHArtdn9sDYagn5BTaBTvZx56j
c9ER2yVNCDXwDLKcwm/Y1YAkr5lx1uJwQBIrMamhOAWRZhEap1qY3nSCDdhJODwn
MsYA6CiCDOlIsNVtZa/H+/NKbBtjjpVyTd297jNLMwasDjpurIvH0NvMFyY2Y3np
o0GtP4SBZQiLhxaSUpOoojlMcmoT6Ue1UD8qpsBVj/uG0jamsb1W23e0+NGbhGej
eqO3dsOX2xmDWLQz+5SJPxLIIH/RZo+Gx5pnILttUiCZ8lHRr6rxFhCYVnXrqzjT
PCske7Xg+boTC5RnfBHoWl42HYeRW2HOcGWEKrca945SxpuP62llZOAvo3F0m+Ub
9nTsUn/2obLUU9JK6phqF+VEoj99oNkn5xIQbsis2lBLFAuu3LmbfJTZchLPob8l
cKiHoLcTfmzLoC34FfKajya61hMYROjcsSWom+jvgFO697zKBBk1n0GnpYiY46w6
EJgaGfAm4F2B20FS2O5tU0KLZ/p6DgjwMden45Tj/roKbQZ/6ybWo97cSA+ByQ9Z
y+J75orcAFw2TLmghIh+ivJ+HsS31YzcfUlIHbIxjYZyg7/pWYU1aTxJ/iyU83Bq
YY0tVkEP8VxVEvxvzntzeosavG9WqhFyD1/nikAXQJKnAerfPmyjkjoc42l7t33I
j4I1CvHnUUbnkhBDXfiydmkByMjGisKekP8JMu+vqZX/mU+liOh/FzixKWTM37qz
CavBX2tvRCHnPuaXEijkc5ubGCb7+hRWcue5+fmBarHK1vsHlDPksEM+ZZzJDFK8
MTRbUq7LyPlj+j9BcUkGw/R3MLZ5GywOWcSr33xgQ1Pv9BsRD3JRvD7tHeqckdLl
5I9oBHTpRWvQRUUdnOenLGxwllAO6rlstcabvjUIKqbyfacxe7/0KnlSt04CrvEJ
guEVk+wMkT7BZHseLTyC9+OyTse9id9vUnC6UeezcKrIkU5XnJDIPITKuIDNxb2v
pi9Yd3II8UB/ttcnHkIGFFccUbX1U1UH5Jl7BSkOl3H5rCgqle4QpfawOy8HRfVY
5ZiQtXyyvErjcNZxomYvMBrrOx0YANnGMPOoauuQjBVpygOTuBCwE/UawhRFaH5F
stWCWLlfGT+N9ZxHFc2KN1545bvrgIBNnsIuZA3o6Q4O4KDfo1rg3wiyb3WmFQSx
ccT4Zx6GwN0YmD0Pa66NW6ndUOa7qBpE9ufuL9kYuM9/SMBDwDC5if4iWwgM0s+E
4cTPD45t3QZ3GQw9l9w7Jd56pIYgaZKP27BZKxcJBiiejnivI/z+sx5joNDuuqsk
CQIlP8gFVFaJqtAymoL1FiAaA4i3eeXe7bU7fPzhvcaxrczeEwe4uLvVyApf9UXv
muGe7SYKMv1J1c8+sdR8qB5903Z9eoTBIJXQktjCLtKT5jQYzq830cB7lBsswljY
VYr8IU+2aFOsmtztLxe4+ceWa1qxBTL3a2Xs2Vo29JGYp9Qpenxa5ROpH3k3pEM4
MAiip8tnAKkkSBJGsHFMpy9KuBvCYzD9Hpn/3wgXCY1PTamU8+j1dA1vn0YcNLpo
uwt2ZNwmT7hWd5MyVWPIS7n7RnqETsrCXaLA7mFK8FyYPMA7WWF9U3qd+ECsTOcZ
aSkOGbGSn4RaKqX7ckyi0BTDxB4KmqmyvKsJwgCDubN4ulz1J3eXJEtw9Vx2Oz15
Au1x32ae2bBdNcFtbH7wQOXd6AUAeMMRxKmYmXVg+LXGLMw0lioQpgGXQvL0lUZ1
wafTuNBDh9vqtczm9004TmRKhZoVgRa0DqJbG94xV3e+b9vLeWUV8h0i7vd7RK58
J18gxruBcAV7pmk3XtUy5aGy6yv7OnCdXmG9cVhLSzABAreebFkIkW/ujgNlK67O
LKehZ21Nywc9VAyE/FvaZdkwJicNH9decV0wmiJ+yEusAV6OlNoUoHyigLhd+H9J
Sdyhks5bqdyiKpYugaxezcqV0JsdfYlWs/3xQDx7afj1bsGIKDRT/+5Cnf2N7x7U
4UvjYhKzcw38PzxnG1fxvKopi2nrWMVYHaDUbhaOKxV8TFSnSGTHyQIVsIjzbi0C
w8T4x7SdOLC15SiFTOcgF4bLRonGqtKaZOOW4Zqzr2g6iXFC90Q4F7wdxVsCndez
CNmQ8oq1kyxHA9xoqbDSsPvUn1cebFHhb9w8HrKID7N30hbt1agOIrwW5k3A352g
bLmgihSotaqZ3rAV2bfFiQteDdchCSzpPgk+wZim1wzuVFpwTlLYsTC+V1ApHXIP
OCE12sIReKALSExF+VBCZX6mwvgS1T/CgjET4nbQogHPWyYxVQDkWHOkE3btRGYu
Xf05BNOypK9x4CxPV3Qen+l1ZfocoUMDjZxpgMrNoBbGlfYMmSknwdIqzrjXpYPW
8zAlpKYrfoDWVHkisYTJOsF5lQBT2GOHiJMrvtEKcten1j6A064fSyLghcgW7f4V
9px9j7qLAnB/Q/75GV02BeGTdfcHzs7zYLjSBlhWp7Y29HgnAmNst3RvNDERIsk1
9S3nWAOStq7o0bwRdbbp8qP2SobdA+F2hcsgOJ8mXv3BiAlZ4YaODQhwUzwyX0KG
7rD67Yn00lKP4eUhBX44INx1TN7sF0OYkpnnNXsPSp+i+xGIgKvTGQD1+dZLW6Kw
veTQoZ778ETEIzzMpGMNN6u1OuNY8OxMsD+j+0d9Do6q0u9PIB3iRN4qrKqwSi70
q9q3KXld95tg2lUrV2xG1srnoDxw8zkjoUwzWhkpVdlcXQc6n8U30fWBh/lI4SWa
cfe5Ws2eFS4DzSjcdSfxXwnwqGFDiqxOL3dtfXmSaV0d6u5vG8KJHN8tAcIqm7F+
oOj2zxSdcl2Ub79lAbKWvbCHCcP5cwM0DYycf2WYLQ0lruwy+TqYcLHUHl18Jytx
9YLUsyTfGHTtJckovhNlz7Kaki7QqMwJ5CH4/4wpX63qUG/5r0IFvgFnaw7kpqcK
HAL0q85lvMC9RhaxlAvfu233y2Asg6Yg19n4Qysg2EE0c2IwOdPiaJaMXrTE+LVk
HxPNBeoE42J8Cm7IN1z1JELTjTEje5HNlxn3HBhOVVBC5RcL8768BuQA24GOXnSF
6qD/g1ByByXZv6oSwgR+rolWfwx6GD4poiB7myuIr49CFaaPg0RzIVPep3W9DUwf
j/r9L1SUdJoeYLWp4+z/vgFzV4z2OSXHQfxx2UmYMtYxmyQeKdxP295cUlXt8fn7
Ft6BgAZ7F3FGHIsZcBKHfMWm3BRoCGZlKfa5SM2pGF5nASYT4yAkRLzx0qBZ5U7+
HpGXR8HTLa2dHY1B7A2pzYX4LKix/jMSVqDlmqjWrllEnxAI0+oagCDantfCKIyu
giIFRe2jHMFoRErQXNa0JVR6TR1f5zRy0Bf/4mBqiIKZUHfyz2f4IvAf0GMtsdPH
O5tdC4bDWG8w4U/OVR1eo1QPLjnaAfaYFslVg6awo3X/F30MlzUkiXhTCtBseg5a
rPvxq4hmLAgCdL1n2WjhEa+zcB0hIHQCQLyQ4PDKIhYZpnEAc+99RGup8USQ4SfS
yYGej+ZyA9qmpUlHxeY73lU0eOgtZrrfoSVA0qXYBXS+ml/NvmGMyvM4i1aMEaAX
3nwVEiEtrq/g2nHLsL6eneu5XlVqwpjoZfR5qiTqIWWMx45LXdmHO6kNWC86K7oh
fdAOGGSYdh0Tb0IrCXZxV67KMIDOd7/YCvEZu0RnZZ+EEnYI4APp5UD/DOBO6BRc
qMF6irJGv2UPc55ecCk25ZoD12iho+GKJB71RVDPwU9Oq0lBqApa1EGVEeL7Papo
pMJ9wwPNikDDrUlKE0q6gA0DEOZKRdXf9vYazoqXbOYgYjdn1V0ZKhi3qlSs4ve9
jQMSQYdKfsZx+rWEdSH896q7Pa5fFPdlSAnsQOyUN4nYCcOv7CUIBP8RYuk+WzrC
kd9c9ZSLKlqBiSBlflm4C+g9iDh7lQTaDDpUjGGQGZk7OA4k6HBgjfvn0dOQVXIM
wdGmu08N3f+Na/FMr94Rjw6qScVvF55nhLZsbruyuWJvDZ+CUxTpgITzsVESDm+6
lwLN/krWL8ePU6Z3j/fxQy/n4c7t7gINZYAy1+SglWsAq2+UM1OIuFqIBj9CH87v
uekw0EUYK5HgxBaZitFsP0H+gp0ELlUFvXK3yoqdSq5abBZzIWMnOJkDMBsvjoUt
SKJcTe4HIF84UuzpyL9f2ToYFUh+F9nIPRu0sIe0PYoyustuSx1BMg2ruo5RqBkj
1Kd3hBgFzQeIqjLIQoMLirl4FeTarC23k/1/hGRYS1YdwC+LgXwhYsVoNXmgqJDH
RJNfOiXrGRJCT4OoiyiJ0Jw0qFTBC50JRRvWVQ5mAGrOYugj4W0MMO/7/wAvlXMc
eUENyHzdQqkxEARJVDMa6Ir4Ac2vjvVuxj6T7mAyMCahkrjiWT76IFWpW3A+Htsr
zzEyozVuPRu08ebPU/itoepn/XvjyANcGRIaD97GJ32HQv9LqzznocTeqZdXUUn9
sWzDUeJG5IBIXSddxDgzabbD3u884djTJj2tm7qbND4c9KpZCpDdvD0h4I+VI0Ob
2GKA4qkNZnLW09TcFuLDsTZ/Du6v56iXTD0Z7MOaWTCgMUG2RAtZZmNHP/Gh3LtN
3ky3lzxBDK77Iz9o+OWhzKaOgT3V7xz9ikVi4fRp6GfQ6u7Ws6XxFoppMDOKjlaU
GFpWJ0TbRZwR5ziimT+N+KRmDACovBMcqGzOF5uL23GIHrCKAXDi6+Dh3pIjQnYd
0KyV5uxYnVmqL2SrcKUY89QqGhVF2r2TQ6y3Iinmu9lMcpdnUfQUoHBaZEw4xX6Z
dGhR+Km1zBiiHFqlcp9fs+LJvgR1Wdwzc2hsdmlxvG/ciVIC6Wfkuw3QcoPIidtP
vZmEWDAXE+oxHjw5IhsXfuYKVz/A0v7UKQhm+re7cNmEMwSWKAFgzV56nSCOPGiE
cdaqmO93U9I+nMg4LjL7IdaZ0J+T6r+Wy0+PFu0KNY8evzMhcS5q8U08Fkxo8XkW
G4oe+mTEdrzmccFvzwHddYDNoSK9aDNomszVCh4+Be3kxwwVVtdr7HjkrSeKKL1D
28bFdS3746xWpidRhIh67mWBaAR6vGblm6SlR3GhKX7eP+pyPVQHu+MIwgfrbz1z
D/Ng4ZTa39le5sJWs+wUqmr8jFYY+1MX9WTXtVKoI138yaA1K3krHtfJt5sywsAp
WKWV6fT/6HTE45tnSnaSz6RGZ+ECu+nN375KW7oVe0x9/X9NcGSg2nk93HZmaGh7
DbOWqDNkSB/t22pIe9fZgoa8bCzowOd4dH7DCm7fy9mdv9UWcEWG3AW/HL2IXLdI
qQI/MDadL2ggxQu/1nLx7I2W5XrGoOsBp2mp/7glxlIInT2lhwNH1P5ZNDgpojaD
UvO3IsJgAuqCNf5D7f1W4heShLqyOnGES4pFcv77iB+hpGWQPhWI3U1sHqFK7m4J
48PcoxbTeBoFl88Y/fSALxCarIt69j30BdqwhNeC3rElUGbt/e7pKv08PnJKCSGu
fOOTJyYZi+6hbIm3SxxvkulW+AFvAerjfltJUiFxIiLnUixa4ZORtLZbpHs091r4
TyulFRU6dyTUinv7Sa9w0OvcXI1U6AsUj9jC/OaT7mX0qyhDiJJYACFQDp8pxmRJ
IBRYtscc5RBZqFx6dzKf0kJNXH//Iy62ZWwwbpWNwvjgsEDPcWWc26oi9S9qnWxE
BJztV3/wofYhmuOgI8PlGnlUzVyn0xCJP8H1g5N5xjt89zL8D7meuVOH2pntzOHC
Fgt+szYGxu6QN8iUH59ucewfpa0i9e8RL+zefY7TNogxxgLSWo3kWjDfMRQyr4Qu
+lbc+Sm9Y1Q/dTAfVAH/ds0eQSjIkJf+13OKlHlG2xuapKzi6gQwmpCBWSc24xlX
B8uKFeyi/cqm7SifHrNfgkDrmJ96/0cYA8M+ha4AlHDk8Q+EYDdldbKKb4yV65Rg
tzIPSVzoBHplucpESfNQdnEcbBlShHUW4SBJ5P7eCLDrZiRvRWy9w3Fkn3IAV89G
wPCsguHMpmyL5fzDvMvL0ciqMglcM4Dbam4vpIT1KI6H6Uw4t2q2e7xY8CwV6z9r
LxuVGCd5y6FZCPYCtCj/pzhSlYGvrVgUDAJLKpmSMfNL5Q/CLJw5o/9x0fdSoqOK
6tokggd9Lvc/QioFw2M9TU1npbKExlGJJMRMBDMJECDnsj82pJPs02+wDfnXwIgI
o0/S5SXaNNV99xANTScJO/bHZiwZ0+M1hgsVWM0IO6+YdCoCylLi2ol3odL4RtXE
sFb0MCH5S2YhlI40ls/DtZfVLAc1NbOWtsCzXxrgXItuuovPrT6FFPEIkIkiULre
o/9wzMpeKk8MRDW1am6XvRmlTPCYJyfBxylGqXeByNnt0gaivx05krpnwXApLtBH
4EW6NqvZCt5rI56SrrTJfQkWNubhKl2wZzuTR35TL4m7IzznVnNy0aZYoVmOGXbD
9tFT6YX1f7INVFK0abzGwPIBFsF2FfwTDr+8D0opQEEgjn3bQZuVsfLOuc6Br5YH
/CWV7O9C8fkaknSv7DMaKO4jdGoPAXX/wzDLTqm/3tNyusl48OVBOhKmzKGbBKSP
adT3mbLCLpbQpw+kFKKaxmEm6pOcipq3JJHOIMBMPEfvmYelmqHcOQ0z8ni1OhdU
Ixu6Yy151Y7/Hj5R1DdrDQoHwjYwJW/JD1EUdotm9drZeKGwDUVhvYeJ5r3CZos6
Pld/6TB7L6Ajl63gr8ELcFs8B82RGv7bj4r4GL65vz6PhHFhCtRH3QTr95StB/MG
ZF0OwM/W0QFhR3F6MaaBulUGKn0gPCvJvaHqR320LOcWfHex+tc0Xic0h26nuZFO
DVXF1M76JEEsa0ssNbghOLpbO8XWo57QeMxHzWI0KG8AWclzcSFTSlg6W89A652z
y0YwaaJealztg9MNxFNrpYbRVdLDo11UduCHcdV+FbC2Z6CTz8+j++zxy2+E3n1+
TzaH7K7paEdJ65oROF+np8ZOvTyEnZSgP9Quo2ey6qaJTnZevsSFdnERRFoRygkq
OPdnhdrZiWCqzBTcT5lWPAcA7sLUcasumKT2Uw03SfW8z9T9BR7X1i5Uooe0AOj/
nh8phnO+FZHsJrr2fdDAY95I+TwXC5ira5hz3iKhEAvIw1bi843mt//FE0+4OIrz
8yves5s7WZNNN1VWALNardQix/iNbpi3L8X7ibOBHadjWwhFwyA9De512pRuCDMM
m8rEp8aCRlmVes3CuVwcrJ+596t09vd3TCSfe6N/tXM3NnFWyMXMgD/qfKs6H9RN
vSWykF+1hdE/UxdkCi6czytMYCx35jwfiExTUTSJzZ38Qr9Qg108mw4lyO0RDyfq
OpPwaXIfrzOjRIvpPqGXPa3C0+zFvztbDnVRi6fcEMj4TEoxF6LwV95Md2JJs+js
/UD93IjkSqUKCAl0VomRAMcCxg6u9g8GYuJAZUgnlKnbS2p6rf2A9NGa7rJzuFLF
HmH7eBvNRZNzoR3cATvv+Uu3ekgmKhga87WP/KHwUXAfgS9MZyM68GqSFebuDEpI
/61Ro20Z5ZlvuW8RftDMhfsArzVs7ULfAd/aTzJ6pGYe8u8nF2vcjKUFghzE56IW
K9cVL01v7WOeOmAKuo/FZTawYwmEQltKgn37e6iG42MFhf2qZ8O0nJujRUOLT/LD
tn4EsfTMr1009D7WWTQ2wzLkupVDNAjVrclxrzO/KVW/yXsmvYJMWNzDeoxQpeSI
vxbXlW2GGUPKC/Imp9kgBN11MGQNQDFbCwu6Km5qknGeWcjm0ckP6w2PvPpWmkqi
DzEV5zQykNwzq1Dkyx6SkAbTh+FtmHjTaVDffVin+tzAUy/8iUsw38CImGaGahc4
uZAGIIRII9NFG8fkafEhwuayoXsxuhg1hkCchwY3Z01nZjaC1WK/foyLM85eM9lP
yNwi0CHjM98QtlOOyf12EsKt3xlwM/KML41GSmQ3gVv5F3oUOnl30d59QJ8rLjS5
o6Om1EFCWHyXnWCNr1YoasNNsgJrnfZamyIVr6H8bzsvIClTdk1Gr66aWh5EDpEq
vIHxk7iizOmTbbOhzWXwUkO8oln8Xi6AkS8oI5HCNhsOQjGyt9ek3tavtyGxSs9M
g1VZdycbu5DawkN/FacBmBebmxGEnSlISCKrwjawkaVBuSqpq2B98KpEOYyEGt7r
9ZgU4DueQFpV75QhGSHCp1lcZKHRh6ktUpuAHuV1487qQ5+D+e5eykfq0swaJlM8
1XXWk3ozhdJhmJDgVk/Lbrm8w0DJrKG7qdquXQCEfqS1PWILnvyFsiN4ew0uyFaa
xCSNVSj5Q7vT40h550IxcR83V1/p7Hn9ZkZLemrldlTRexrZ9Z/JtshbUUA518/S
ROZqL7sco8rmBFJwZECUfjkXDhuCw3/rENKE+S2iHzNcLqeWnUiJNeVVhxOEEd5c
d5A1/NFAqu74kh9eVejZtPEqFnOPLbxDC84AmAx5gHOiPnm+2Vx8Tu7VBkUvYuBY
3BcqdKCy6/4Q5ISsAzxRsJZxfaehvbuoy39HRqMdh3qMbgTZzimi+ddoZeds7KcY
FScLSghTuxnjznBm8oGDPaPHiVYgK1GK9nUqPcAb9ZOTx9MGSC8CoKMxOnL1ly6k
QtxHHYU2OSBjqkdGVdYDG4g65fPDz61nabDiQRsA19D0E6sWU57Pg+HR5PUQ1Efb
U4YRFQPGZqmM6ndFyG+ubOzetGTwM/sKi/1p213FmDHDOCvk0ukqZ6wkCQr6VOso
OfLyOseRksElJsgjmvgY79Z/bXIZEdog2+3X/oihrktTjNA0oGayKPyY0GTwgyu7
XosrxRCii7I7DicsQNmicgmcLnkE4IR1ZXxHTq8Ay3Yp24jl/yR9viahcnIJfNtQ
shViI9eSYrzdVtKhvRbVfb/XmxxRIBjciumIzSf7zyAMWA2yg4C4lUeH3t532ekn
Tv4bOfNUj7WeSeyoIEufxMjbpMlHEetWJ8YQSfFM5Mbsxi2q+mNNzBOhtaayIuUW
CyJ3tjCTukeLJ4MRi5IQO16S9sSlAW1uazlnr949xQ3HYwWwQ0aCuRJxwLBhMl05
DuXWe7x/7RtFeuQzRQZwnmZiFcaFPcLkgeCs/eG8qSbbbrkSL/2k4G1A/oTBah+t
QEsjFbp69XT+y1zrwgh2YD6NSEEf5kxuiWbpoRX55Mq6QcM5xG2FHzF2ofX3rd7C
L3bqECaTp7H6Rz2v1TwmaYYxfd6S9DW/xhySJFMvHjwDT5yx7dJ+1pt6okeJvAdt
w7htITdV9jK7u4PAfET9Ztb+sJt+ykZ/ECShX6Ru6gFnPqHvf1NrU2Ddh7zsk1Yy
C4Z3SLQrgxGEr/4jOAPtMKBjpUAFtNIOr2PlT6mlPbDdjKMvwBwu5KnPcS0Q7Dg8
PTH7Yrb95hYO5RUDUDQeGwslv5OUOoE5OGcafrPCfU0VN8mosPkAcLtWGbgH5Ndo
tlbKShaZ2CPKYSZX3UtvIfwKESHlxFwu77n9bKOPSLqDeAL50gxIHaaaqw6kcGEb
qrafW1kEjeut20x8gv0NDGRYxbuAFatHP2LIaR8BeNlVUrROkql93s/nFrjlvBwG
pLQP7JY3Oht/Mtc8RI7OlmBLktp29DWKl4YLmcyPvVsmBXpSmJVRpxyhiFO1Bl+S
bWRopKcMDE60Bcc83VaQgbvNdJCvtOE6GnXFdSIN9SINPk8kYaNoX9VNdCF56PjW
3yQTadmDtVfNlPC5iSI8LDGpUf80m9YwvlHKGjFdtPiTwDgPTxhG3CQ2fgjNtHYQ
c4SMHgMCZp11yY9XkEHlOuo3FQXnswivOUPO9f5OWpmHqTkHcJqKwVv3S3oT5Kiz
WMlkJwNcCkR5j4rqgkWMvAd88zfR4ggP0vsWV+SRzLV4tCRj4BAFzaiFMPfpfSnj
03cBMgJwk7u+DAKUVzotGHD/0twRJDrHUf78wTRKCD7/dC1uswnprs8h3wYIzRZn
oHRqWUWmSu/rKAhiS+2ZLF5QlCfsuhxJptAV1Y+GtTpf20+KOOG+o1H4DDWskNcP
h4BA0j4dkBzfKrC+LLp9Ct8G98rKS7XCAoA8VU0PHCjSs0h+xHBthnNfjo4L/tSt
5RQSVTi5ZRfMdFMnBuJmZQu9qBR8x8cUnyGNTW5BIk6eAMztApgiWQsPLoLUO8Qh
CWWuGcsYwwSDJNmphfyifpNkTPXRo8+VbS+mJEGrrmYCbhAjhATSuHSJGcEzPyoy
2eWoB9kNb1X/veD8gsAyafljAsPD3g9uYpTEQrtj0unFDJILUthNjNYGNxFczCSJ
kaIiTprgcIpOXRD5ll25iceEO6NpNFJlkAphwsVFMDnC2CumsuNEPe/uZn/hZbUd
ibLpjhSuDicdt1fKJiGx4W5VVl/yh4ePjr3N0eA7Eet1STKK9aw4tY3MmIFuuOwH
Xz7JftwbysiyZrBGDl9S+8ojBRfFAdQedOnpdM2Bo8waB807Sjb5PALWhTSrqvPj
yRNDW3ASPL4bl0bhSFx/2kQndKAPpD8VGG0eEwKtuMeiia+t+OE7CJXGYkpmSN7y
ARnhSyl/3Bl4tf4jp32Qy7d2g4IY/ZrZJvB7HpphX66hYab4eZnXsJzI4/3w92Tc
CHhCOiqABycf0Otifss8LI9sgMzbbzEzYKViLIGrDxASfXbg4/TenfRmUe38rsOh
n/kigGHgKAQ7/XfdUwtU2V207MVHPvVSBKB6N0s9FltfNajKeWF6KL29uK7tsBEN
y+AYSXyuyqtrkjso2H9u8KOK4m+F9rWHHuA2ApwOhluTmYruTdVMCRfGJNjHam3H
btYFE/f0GgRXfXJzXn0p6JzkkrhpYIokJW0YUYPo6oz4NbGUCE1sM0CSoEaKqehv
mQ9xFyx6Pijlvmx93EJQt6Y6UnBGdohE7rCVJDBLMNd6VznWdNuq6XgZ9lwQrZN9
9WGfDIjd6FUWDTA/wnU7r4EThZ29OzwElzQ/2qVHuvkdW9/u926Nmm11ezaZI2+J
kvTx8dMO5HK7tAWYWNqOGJS2zQeUmLkjViBrZdeHBIDHUP95UITt/UVQoqW0TDnH
4mTe8H3oHK7Qi9snlxM2bmCoZnaaVWNEDjineJAH2r/XkaPL39ez9ySixJuQD+W+
36VT/fEn/uH3Y6j/7ukp/6Yo6VA1bqv085Xo5jmz8mXRGYv+JJJoSJY/xvcnd8UR
6/z8p1lguAVB+uAaY345YGFun6k7sLsgjaDpbrdCZwoBkGur8VWMDJ/vEKFSgqRD
26Jypc/o6O8IX94ZAddAK8oUVvoVucXNLFvT93+VAWknhxoHmB6Zf5qNOrlXmhXi
T/v9EEXPAI6Gt8Wd6rhzHci1EWs7m0XPKOUPRr6hQ3Iy0lingSzpnOlK+aacbQ2b
wwv0Np+wBJ8JWe+bfS+dHteGeWwwg2ThVBns/nAiP46QCPezGdeeDk+kHQHdJQVi
Yev4SyoZuF5IOKkvKX2WbYqqPK57djXVVTCDjHPhiW08V+elDlHNGshSRXw2nTnA
BQqPLGu8cJWqa47kKv3581xlMWsXzOYp6EOAwrIA2+0kjBzjm5EouErLAosd3liN
iZlNzQOSmngtLRj74TBNAEbjnpCd2S/k01b1Qc/QlFgcTSbvU9nU7COrxUr8Ko/4
SMYJMSXMmq0boUW2TqX/zapgIlgbPhckOVfK6A4YiJuaJX5nUtA6aGYC2MLShvXP
eTaRqksLuWJXbka0siNuqucr3neb1mCSVcyUdBqtQ9g0H1fM8HvGnYZK/9HYlvYb
vPPuSzSt2r/ygO3XLjxhgXqeAp9GwChYwanejvR4WTQjnnUZitmY1CYVm9AijcPR
xMsjPRyQ/ema7CScbkHq5w3+atOgCOHlPy1DYJckpMZddzQSIX+SUMLX8eajA0bJ
LPjZxPzqqvYSBv7xG4Knc9G3W+K/NN95Kt6Z0W2NpA264bMqGCJnbBG/4TBpkFnc
vq/wE0KxEvnAZdG2quKXngTV4a5FS/jF5+iFDCu/s3BvXUz7SuIw2ZgZb0wwT38Q
4J1QBTHMYJVcjELny02pVF5BKb58y7qVw5Huz4COMlUpOcFFQbLL6gWeAgwlZOAC
Vnut84f9EIu3d2h51nYWIHKqC/I9JiTcq4e+x1kxmNAk74SgPfwYMLxKpRnMV7ZZ
XXjJSbtn/SPoSXTjJNafyrXYuo86PMtj0uTs800+Vm+NewYa8tjbhB+iezaomsy/
6TW3nQK/YoAHo2qkUmwg5H2uUvG2LNGshk64gSSLuEnM5WzjM4VflAtTPWkNWeJ4
GPD/a/mrUpTM0HOhQ7BsSWe8o8339qd23Vx2tHSjno69fqszuULW8BOOpgJ7yLdS
7BYvf/QvzkJyZ6aY1bdZiaI4JMAv1GlWSkFbyBQrh3h0Kq/mAdOUysGpj09yvwGe
f2PvXzJ+l5qCI+hJ3wlarxEUI/d2qltmgHqHedAqAMs6Gp1LbVSjcUukRARRhrik
HoczRPXQXSNJAhpP/ExEkv3OT86XnvwDX13+yuPCp2UUoPtkWn3ySygl/XWd2oxr
82mGLOqqy2SGl8rnoFFoAJ3LkRfDnuWtSFCKkRcTEA86DI3oRYK/aOdi3aPed1Um
3OGcVBskWGxeaMD9TXR6TfSI8mnmLdh3MCCxzbuGIjmJti767PnHVjKlEj82/exT
MJ62Rmyadkf2c1c+2+oYQi/zU+fyp/7AT4TWOGhrXtHPuIBzwPwyxJdwkSsq2yxx
azwrjuGw5LTn8dG6WBCqQ8+fvCeJhcDxBy7J1hB60H7lyDhDBolgw2ckMQh+sGvr
z0h0jNookgj7pvn9hvOfFOKKeQZRu9ojbzGjkqV0ahQXK5GRcTvntBznhibbElxj
+GYkQEpd0KDr07knnugveBZOK0oSr+bKg7ac0L7a1BoZlqFS5MjDfEGhYunNQ5rO
Q/sVbQZMW0eXVyRULvmnoK1NhMiuu6Eo9yktm9N9PDQV1cWHFw0HvH4wlDoY6qsp
u75fUHlxPzyI/6tJoxwPATxkLd4MWFCosW3O9OiKBRqfWTl8dKsYxQci2nB5Nbk0
XXH7eE9L+TtOSRI0C4qSJdYaRloBripBGrKE99zPp7wCOcQAFeXQcMlMVUjCg3mK
4QYZcqLxnF5paY4Pu3SacckTnHOfuJpgwanMShMNHSX4kIC7mO12md25WY/T85Iy
Z0vOC8HX37397SdmqwqZ8w3UvhU5S3dspvPMyAEcUk8Jqc7KKDXdmwsrRtCBYBq7
VtGGNkgFSXCSJ9a7LG+rHVS3xlObfAVuNPc22eaQFzGKlnwQ75IK/HOaqLZ00rTW
xN9FqI2OgdSGjcTstVoUn+zTadzgIfwIdAeCQNFXm1uD+N0MqH2EVUpZlYOyqGe2
5oZrq/wPKSeyATwILukr1PNh0n3TOTDBCQTlYIV/bzaFGzv3TQuFLUhlIYt1ImAf
ige9Ia3hoTKUf62MZrda+ERH6F5N5J9tl26izDBN5BprRf7dzEFfMzWaKZtEYJ/r
s0vBlZe2sRlg/Kho7dm3cBRHohViizT7j+RTT9HTJWAnH1MsJEgSIa5UojxFn6PQ
Pd7U5EJD6skjXI4Ir1PVs08+bO81W1nRe58PoLJTAwNbd8yM/gbIDQT2ke0EcFso
USxMciHD8/A/yc7Y/AS3+5KlnwYXTfevyoUqgNjLOtvHyHeuzebx8clJXY7cECZ3
t77JBBO/oRDZLNqiX0/24Ba6Aj/UXJMTips7uV6EdduXBc+RnHzQBRZvrnZDCLnI
mPZOGo0uRNWpysOzWYGwcy6ZMDVuVJqhcB0O34SN7c/XbBe2ZDJZUFAc653W0zla
nShUQM2hX18XRJfR/T56nOPqGdK87BB6T0e9BrlULQACE49m46F1VcUi2vTSR8b+
vR34OiI04/lLj8UTjbKgZ5yVdK6oSGrCwAztSiS3aAGSy4aKKBBcJpfzIZKSXQik
DW7DyzX++3gqVj+aKkfR9O5dm8SKYqShjvdyDQw/rlgT5RgiD1bh53/FuThKr+df
CveNvRds8de5mT7bXdSS7vLk8ol+HwhoKMQt4AdImqvhPX4l6bL8GVGaPNSJs742
WLeLvpx6rl3jm27j09/+zC3QJnghSEzYovSN3y6BmCk9HM7clYmqjZdzEe+H8cA9
h35QXKxUH2VfX99byuzbGBH5GIjq31cAV3GmcFYyAzJl16UJlVaCgrf/doISCTdE
W6m07RWH9xfAGGA8ObZwdaZ7PkY8u67na+DMMgQEcEaSAOUabckgvjgwp8+2BBM+
mdXWsMXoAuTVdps1/eZYkPoFPda/Gl/v+Km5C0c1N5hMNUhbQhQOoj6YKDBrJi+a
UqMFJ5nqTxtLFCDgHFsM7NUFGkEUg9i0NPAZOWRCscrGb6CbV0LCvaXkecOUwEkw
QwWYbfLX8mPcwo4DYw/VIeXKHX4NHb++E6JvAJLv61XSIBUULi6oFDhFfDA+KZ3P
8Fb66uJD06Vby1MGVeDHD0SsucSh20RIv4QkKG9DWOyj/8RwWdshBSQEapGG38rD
B1QQ3xRBRsnRFHPzB9FQh8JTg7IhAEuMrFKhGyFPagLYdC5zW05M3jYvtboV3vmk
6091aXuPK7UH0KNE/lUHzb5Ez4+iLf5nO8Thvfj/IJRRr0z7GS0p1jY15kNfrlk2
wpVbUjWqXdklUOgugUnZG90vdYd9uXLvp/NCdxEkD+uEH/dl2EzItJaiWUc34VBh
z/lsHbyBZCcDqwhI3BzvOVotydpBYGK/lCNCdMKsEMp1TVsORWIBgFbgQ/Lv6AHs
51M4OE/u0PvZQWhdFShXugqfWfscS6tptrZgPr48paEX6tCJt3BsMMJLf3CpJQ6f
zyzrSa/AWn7gHNtS2evd7LHdjjkEfmBJpNLdKGhBBT2hUw3aDWvg1J7I1B4DjdRM
uy2frxVsytN0Xq6HzxucbqF9dpWYUXzPeGM4CxEqszEH2GwYiCvBfHjiDifdqBuX
8fgLlKqzw94Z0VBni+Zjr1ihDKKKmKk6bGaae6WGho5rwkxdzRiOg5vdhD6YVqWG
wqrMNZka/38jOLEm65YFtvSBJvXb55NHR/9Xz0uX3gfIpL867kZq8a3D2nv9Khk/
WidwqSAxtlFOdO3o+DiERb3hTYsMcIE+GB+mxRYy7nlczAhCeXqfFT8wEBciVSk+
wXsyM28kZsT/piJXPJGJIvb8d7p+VIxTs2exBwrqIFIYSjs4Mo+g8WXWJUaX6UNt
3UFq9qGL+ULilFXhi/unpketN4Hx14+DKt96YaBei8w5Eezm4eAifkHG81EOzDeK
ySZIbIvGqK5WlKAqeDSPVHb885EFJgxoDQJvvwKcjztw927NuGkdGDtbAPu5wDG1
sD0LOOKm3+YE6soio2dUBafmggNH048IG6A7rosN2x1uKqmb6rBX52iaRPcD+K4f
bq5CZDIteGWKN4t9CsMV/c6GBDYT2YIFYgVk99Tr9TKNTo/Dh7R+Q3NrEk/rsF6M
BeXea5IDqRzsyzDhS/+yHL3tf36cqmDO4bvqM/S3SqdEroe+mJtKSB6NrS+6/7Aj
VouvMWB7/x3dcdPtmDGUYAuFXegHcYZOmhYLjG5mAYIFu1jieolbdj3qo7bNYk6R
5HRBfQd/cHtg5Nn0muHvkDGEmYCN2oOzK3Gz1eGazD4A3UkOhYyGZAF7Hk5jE4UC
S4GTYgUzpfh3eMR4KJEsvIzsi0Yhr1XT1upmydUxnZkSL9Yns++72CHFLxxKp3/g
ODYE4E7Bbnpg2nGum9QIeCkys56I2myUxbq66o9BSj07jqSh18cDSWId8r5ELEed
vDZXECC7u9ylyIwJ5CEKBcj9yezPtvQ9umta5fzDd8yESo0QYjtfzDLserj7CGRI
RkpFmNHBaZwUKL3Dn/ySb1/EFAL4um/1IiVayAsP1iYIkjTAslgxk1Eyin9o/vCM
ud3TT7tBGSCilEBbIfG9PLHdKKWNwXKtsOZzvsu6go/QW+zdN2wC63c3Nw3bwo8V
gnDCEG0jTenxi6jQimGH2VujWggGYw5Gko/NdG4wPqa9Gd4HewbHDK0ZPDnfYec8
GWNwc+QEicH4l1l2EdG++vADa1hzq1TPGZro76ssAwatNj/jk0UjiwSpGgQDrKsG
adUSL7VbxchXwsCfcNdjxiTcUzGe6n6/lZMpj+nGikPN96dhp5Z9G8uYgG/9mBF3
WyANwfUFgOJsc4EufrRuFHjgZwFPmLac8bEFPEWv30I9vJB1uqD3CFoiC3MO3DZ5
VUPPvNovZv3iVFU5tBK1SsWo6m5qbvXvK+dm1iu93FvC9nbhbTS0ZcETpRKFTFJ2
lyeOynRdB5q+mQ0xQqEClW9x9UDsN1H69NgWQOJqfYDNXVbxrRYXPRVkewnAYGVD
rV8w2xEP8UQfUyNv4ZYeJzGd74bWrs9l7EvUmo0sStmfgyuh7nma9WzBe8G0Ap6j
DTB+LhY30PoUFg+GNG/wUYezBQDrKpvCcYK6OWkW+XRxWEX+MFU/Wk8TYTtwFa+F
7FFmejyWTV5J8v77vt7peld81PLonNGCetZWPAsuo1JrA0dVdq0U7i6hfKaH08dU
1TWR6TnZKx6r/EX7QqbBZPJyqD/yNI0knkuLJKNKgOuY+dGHqitT6VddtzXxTXNn
E+mqNoNheeYR5lgN4i/+xJo2vvdoUomYGDBpez1lq9iBPZdhg+cEPy109oKtgJb2
Q+03zdIZYqjpZ3D8RZh7X9HuO6mIqKoS/bpz9G0fmj5VOyg0F1NrPeCGJwN2GaNW
BzbSIepmdYwbPA8r9ooT6XsSSzBJq8KGKuPVUoOg4y0VJ25HxOyAKIyZQn2Jc1j3
BmIHeNgnNWEP/zsgIqqpudjleFm8ek+OUaFjKMqG28662qm2Qpak/wjkxt9vpjzY
yJkoHx/JNYvV2maEG1kJfom4Gn6b6qcB52PcbQ8Zi9svKkazrCv2lqlnmRQUoDwj
96l+K+68/BNdJ+wbEyqzWgcBjtiyTr/BdIcEGONE7AjXxaGdT2IIGefpXRJtzWaE
mw+6lsAdRjk709BLNnrprfObrtgggiNic/f3p4mZ/v8teaeTDX2wKLN8HrY0KKIz
11SYxIhHm/qWD3x7w5/L2nNpL+EHG7ix+9EFeC89WVWUFpnahVayrt1qZ6UCWgJJ
Xd6080UW6U+Hrtyw03ijKOEasv5v6zTtg6zrDDuuG0YD6it+pG6UT9u3TBqvSfMd
spcsD+x0F+GI3/78OdnjChqEvPHqAyZE72vSVvsqCaFmoavL/JBcTkIUN+F4NK1S
GBnsAgI9w0r1ckg8jNo+RMGekd7BkYd+/DlZlXHrgXS1gVNuZqCptQBug2amRXIK
td8uA72cfeAlx5sWBEjwMrrVWGEnOpbEfYZ9l8LqnAzQ8VA1HqPPkZj38ocfec5v
V6+rU4ij9JJIGVD5kl2UpEZOLjSvAVDhZMoXP160JRsfLNb1WmwLLFE/IMOto8d0
UPUh9aJKfYQRBgquFJwreGknc3wZyI3qilumRcBHu0Y1tfBPbtqjQz1FBF3dnQ/s
VNJnaiA/3cLmml6f7MzfbVdzhZMnPbOe317I+p8Zeuy1bAC7fRqzAciosuEe8pI+
oc4KaUkQ5nJ2dfXVAauLDVYcw48WIT6bNI9dUF62ztFUDSfGYWAFKI9oYL8/o5tF
jHvwAMZtRltTiJ3FL/V8C4sHrsYKor9dOneBJz0iwZijpHQeI9gAFitdEVMchNUT
FAYFYJt9TxsyV7K0QtVX4FfFjmRHdQacbjw3JABez/sNGNZYhHczWUJw4ilnSypH
S7JOYCQaTFReeefnSRnNSb6IQVD8zJfjZuJXSJosgYQTFWQCUUCcRhwanXSqnU/6
TS9iXDJCfMCiLMCXWEJSTuRAPGUUDZ8+KLfP6+XxUoJfzwDaahCCTlz9hGp04P4y
U388SMbT9SxiGJau8AuQdHG4XlKXjYw3UGbYGTpdN+7KV8iC9D4GRQJV7VVv3Oq/
ibF2gxNE3Ss2+RkRC+bVSi95bL8GuufxZFYZkWREUgwmHfJTzAGPmAXwTHIL70Pd
ogBvqMmHqOxz2tr2KzQwgLN5I9wWZpfEu+LFBq4YtikWwebXWVrPTPbCFt8X8pR1
m+hYdv5mIxy4IKyT4utsiOpfKpXX9UqR4pF5LgeoKHkNGY1ND2lKjIkjkhx79I0K
f01FvkSgPJYmyVjcQBiBrvciiektQVPSfeMtYOVM+yuquKprHTylRUbl4x0fkDOH
pr/2/aycvKdhacAi97ASgpW7jG+gaormr1rTT3V6/TIHIQpyr4Ev4JCFosIrfe1N
cN8J7zjaS50eGgBjqaZO6iz7xE+8Lemacqye1wVmSVAkrKbBjjsqJysrA/1e7BgB
mkdgGZQj8qxp0x00NOaimo5bip3zbGKf9Y5NC3xJ6vCMrrDDWi3EcigcNDdNZg67
xzvTagcCN9eDx3Cu+ulLjXbhPwgSE/h3HioueylRW97ukFgfWxCnUjy6GEOP5grd
GesBnogiZcTtTgoQ9tvqgwa3W2hVk7YG1ElW6P7HAXK9i54MYDeMgE0a8byCU0Ot
Tssn86l8Tw6HzGzsD1JuS2mvJyF8Y+ZpK0VAsqFKLOGjxJx151IutYXrB1Vx740X
Dlb4U6eKTdo4745XjrQIc9A3jJZH+h2nnenFQYclppfCMRkJlEh2F8czsog4b5RZ
5K0et5VhV2FYJZloM69xizWsx11Zn9R3SxI+TA/k59QpYuWGIB/ws2JtXYQWNqxT
hLU3sON1JfhusUgeye0fx4mjeJia9i8k0F4Nh+WEYMrbc9fX63VJ/+NXxqu24jmB
+k6R5NG5acxEWAx+P70/J1dhXMuouh9VNu6xYuTdep3Fk+Z5/UTr9cXy5u9T6kJi
sYeVJqz50+XgbOuVMdLW+wbTRNvuN7OpH+fPaSf+jmD1SFBmjA3TlSqDCE2rg3p2
1O43uBFDYDFZNjhRPj6KPy2db9S/3/nQjI2W19atQe7iRBCaIhEnGMprw5mWrXse
grDfSWwz+BOsxhoCxBSSD5XBa7wTOWfESqrKI0dnR2cEXGQ6mu71tNdKsFrgQEBq
j34ghyZwCEFEFVgY03a2AB/R4o4Pfb2uFI6JKyoI9eklVqz4ri1/TRS5LDp+1u3w
ByBm6iNHAWgdpudMwZPfKENYDMOfcIuUJ2ZIZvB80FUpYHEo2JPid+vdl0L6XKAQ
a7UC+JeSZRPpjUyo5gkZI6EUA2t65mGafDKfclSHc2oL2kHnbaKrFcxndilOygwo
cspUbqKjK9Tx3phHKa7r9b77T0NQsZddTDzKwdWJaPqED5MKkVJ14cvmSZ5X5mg1
fUEAr9CFJ15+Is8s8VVUN5tldHcrubpr1hCV0PI4jP8Po5UJpfISNCEnFU54zr4M
ABI0rDmCqZV4n8nahYosc2AzRMGDLHsGHq3XvaRFGy6h+LJrUoVVgR9x5ngpSwyh
GRttFqpnvZ9hJADZjW9liHUQEOxlzG5deL7LTP4vYUYTxjYbGmNirDW9TZSkSmEG
8DZSlXHD1bw9IV+YN2ZDXt5Gf5cVag+qkzpWqHxgB2aWO8yx6D8uh1Sj85P6Co9o
S/L31LZ7+Mue/HeyJVC3WvrTDcHNYd/6AnWGgl0FG3pef2+zuRVPBLjEwxGIAs7m
j++f/kNW9Q7CFmdW55Yls7pMndxi/5yq/SJfSLdUj1mcF2WF09+CICzkhnCpQbIn
nAUiT/8zSvMzxvqoV4sB+bmeFrkdfyQ0v6FWN1B/PLTYB6dMW/dmlZCkqaLpWcaq
IZ2aO4WzS98qBUFiIr8sqrZVyqH/RGAjZP0eB2HTA0nTIoXcikASuYTz18W4y66F
8UFzO8W8j4Qty6dFXDp74gkZUDZh3XGHI4KZ7GKVP8ivq0cTjUoKQJEbPYCeAqkX
EiJ3HQwgvTie0GX4prKQygiHgrfy21TUyxQrziDudcd1QxXATqlUjJFv6qctjGaf
94O82xl1JVuoWbVLQXLmKYSjpOqNImu0/ZeB5WRpBBEogFD3r15DscEI1z69EjDU
NUsF9YZElsWI0PvoHrNJBlxrApAGOMrXJopiaP63VFV0n/IdxW2E0NanhaShA6KW
Yh5+pIeMy7B6TjBDZDlKO2PXKrb9w/ptNltxECW69bfQ3wvQL5O05XEv8XJAWWhC
Q10HDzyQxvgyizkZfC8SH3uZ7i6jrXboPyw+jjUnthzKEafGLLyIAOVOsg3+BQUJ
FfaaM8D98N5sK0Mdsq1EsNA7J7DFwbK03Orfu/cOQiGUuSuYmiV+TYa5WEXNlguS
KssN7J6AOcbYjL0RT2D8JygCbpYmWcjtjjriSGj0QvR7OX+iZl3aP/+oNl/YRab0
XNsOBEmDOK3ucJUsU8k502nXeFdxkSQbRQsdEIsVIgZckUl9B6YONBqAs1u5GUoe
lBK4YpfczbzPs6pjofhSSpp0LnKySn3pw/JFWHkE4SvZavyizvU4SXtdX2EmSDYY
PVvVPMDefduQXYyAyR2mdPttQD31CG4uEvbHrcehCKXdFnsXsaXDwltThEtQNjFV
zvLcBv6CcQYFNmHTEACH9I8MfQwxEv4ptCVWD+OdeR3TzGHx8USCRmYYKpZgSHuh
1DwEmK+J11x7g7dUJbE+axwVV94BJYz7gjomAcARLM4ql9SkUvldUNxsYuOZmul5
fAHuT1bMd7aFuqNBUdcADHd4ZVpOqJUVKLm6ay8K+IppF9rPpXy4xTYSJyHB96lA
y8vu4F6KO8k/Lyt678jTuO4DlAWMBvlLWUm+eP2mS/tfRgHoxLHLO85vbPHvCKeq
DmScYTKoWAZ9oK7hNQEXKFpP6xare87YXpfvTWkVjsP4sQutcSkSzkKHtqjL1vgw
lzBDxkNeJCA1LSZT9cdt6CGtIFuHgortaIxKqaMSLXVZ03zUNfKwW7a/HB15u+xq
g6IB3BrB19x0b26Gs7CWEHq+O87WCVsZLqa4+/8JCjxFrjZcHqo83HrszKHic9k7
YIUtrmrNR3EIJWti7uvVOAjEVfF6+SCGEAgXvEEdjdavYBMYjZLObnUdmoZJMiJ5
Ql73I23Lr3+EPTielmjI3RSVfwWUWG3nccbZZp49aQ5SlFJU1pp7+RaZqsqDL/3V
GXTludDY8zNXdmjgZdcaUSl6IM4a2nV4aYQ17PrXUPFyz5xPF3VQMX0WiuIKMEyR
cRXyAH0Ovk2fIWbiaBDQz9OZQrIXs+3AywptXKW2dsY+KQehE1PB3UBGm37b4ZzT
LKEpYMP1jdK9gFcLpbr2bXw8PUpvFy744SpZzd72PZ+LDKgtq9DzhkVOLCZjcoVv
d60D7hEBOpGIayeriJC3HWXwOuFJVSU5eF8Tf9U6th1S8KDk19b8l/qHyaCU2E5p
cc49AhG5S6l4DT1YuSO/j6N1hbqJmdVTil45OdGDh4wQf1gUTuY2rtHJzROHRxcA
5GsvTeTaNzCb5bqAfa5JjUnVTsM3ySzEkAtsK+m3PLEpZJgtO5QxRmgLeIlfDggG
3YmZ9xaoGR3lSyJUprz4YfYAuQXlHDKy+eDZ/n4KB6t9+4vGIuRjDy++iIeUo+z6
6i7vhPas3MFeMBHn2vlm239ob5e9fVACbzP2aS0O9VVJ1IKTUHKI/7pdltONdwQL
m1XVExsUvVnidLMMktXiK6EeRJhBhrIEIzVXRziZpQjam+e84bfYCLL67WEM2SXC
fNLXSCwnG1RUJzFFLp0NcCGVpAhMZe3efMIDrleWRIUXVRsBTs8JUCHLCPWi6VlV
R9iC+IiL48BzPif6B77Da860vBXjTZ+rI4lhZm9Rn8tOgBLS3foGHYuURSnu8rWX
3FxGKmPuC40NB+/rBf6gXPno6LJa+zgK78ZPjReOzoiG79MF1cQIyAeoSqkgbwi+
6O+y0M61PuerrlABZ6WP5Ebj92pPjq/+mgd2lp6eYWPd/QVceCnv2M9+mPDxLa4I
IykhIhwi0cNvKfesAoKqP9MpOKZ3q7nn01I36UMbMga2EDuUT1z0SPXoHavFL7zD
GIPFCzYD88VEhpNLjgcBEWgsSExZAvbistT2jWQKTZIkZwOG+coPHGPTO+y86O7W
I73bLjkh8ow18lk1+JDd+HBSvvXGr41IKCaAMz5t+4ChPbpvtuviJLKLrGepIxmG
GTOZxlS8uuLO5jJUtDIes2L5tRwDlqD7S0Inl5L3rk3jQXYmBbIQPQS0jWgM8URa
4QX/kJ0ORDb4YspGbmsUdfqbKn3oRERUhHqOc4mn3gqVfmuc6HGWbmNW+NTzb7Nx
z2jMrwEycjiZosNSbp96zUqZJn40DT1ZFxROoJjuKZUeFnTVk5OZbYQI2hUiYtPI
5p61shartyV+5iDYbc/4wawTdRSFJfBrF+bQJf0XSF4msrUG81pCt3UvGPV8PbKY
4/prA2ioxN7+79F/oqJIuToPbuEV5RqGxDZaqE5oyiIu5jL09CH/FURJR0CUHSLt
GnHD7jvt3VpNDb7zSq4UXFm/FdzjSM+mReCyZu0GPcEJvwab2SFysqYDh44j2a7F
RwnNLXkRwV9zjcDl7i2Ky+QBYGwP9X2QvijHAIRgqSH1e4jPvVIp3rqBi6GlBi+m
H/Z0j4ZV+HzPGIkswnwMOxCsC44tONlMB1a6g5EW54ZqRVwrA0c3OG9wHNW9ZEQh
h0HZCxAVMCVzUcSvm7KCBMsYCtEaeNpfANnfru+2hvyFrjYSQfs2xn57mFZJ5+ic
Zzpp0J1N813QS3nws0ZaAVcA3wjLppzTmzesW/ZoNKZQaMigZTmrin0fDlolol19
FBk5XaV5TpSkDdvGILfqxaFaC/wshrfe1UkCAAm2r9+6ybgUC26exxD+z2r3AnU7
c5bKEY+ebyO3VG88tUAleF7BWy8AyRqlKKmtjhjnvc0RQRk+Vt1jvH1D9wPJ/Gt0
cO+o35EAB2B3cCPZp14zcFEKmOinDLPixJiQ7ZalkmPhQTerInl1z56uVbgAlu7h
irzK5gsK7s+TILwDRKDLQBnJNhq/0xplj1wd4gcghB6d5sBz5E+pM59esTv/Oo8r
U33MYeIxNcaolWueaVRLEh1vJwVlM1y6p2xPG7Ik4fcugtTXE20AIeX9qRKydc+z
4NTcU6nH6lUQ1JD7azUDJkn3BeMppJxHtz55xo+2suz1ggNWC0NGYt1fTk7NgP+c
vbHVgSOLXaVSOuyN2gaX+hzQUdqBHKHp/aj8ckoSap365kLWGzW5f/bamzoENdWS
9zBJGCwP6IofVq48JeEuFkoQaKTqQSw/Mk+i1FkCxM+tnt+jNgEh0zAK+mdWm1UW
afAIkP4FXxwPclUGQMu8kwysMciC9JM7azKVNlxdwwfvzPqF0sYzqG1lRBRRQoWv
AogKeQBix26dkMz3whWoy/Wy6lgJfJ04+qZluP28KqmlwukyrLMmuu3AK0Atbtbl
4UpVOgaT/0iC9zaJlEkSjFW5AAG/BLg6d4jBgqoGLxl1VO0/dpo+fmf4L7ql6tHq
cUlEpcWWeZNZud3B2hiaWMmMHUSJFYclicxNN+KgVzjZCYu8QXJyfkIZ/1wRdfTz
CaxVqE9kWqT+naoFAKVgrgsQlF7oapOB9YnkPvaF/E98pLuU1X9Cx4HTYGtPnMI3
nlg0y0+7DFFARqL2TQ61P90vs44cgZAh5hWLosihEt3BOZUYr6xQw/HcKrbNEY4m
SKBWF9umbolmw76XhemCo4BvCoMqKJyVwhIGK/xc+NrXtEXOLCZntFPctmeX/tD2
0Fp3Tqre/NqdVSqSC7wW7eQMwqBq7OLW6eh0xqq/d9mxL2jtYAFbhACZV0a8LpOr
MmpfQsn8j+QxQ22N/nHVQ7QaO/e/QFRlUFtMZwstEJlEDXaQL0lQ3lXeuwgawXRc
i7yY2bqs0rvkrv8VZqg/QQ6c4DEMixnLgMQgS//05ApycX+iIT9wJf0HZ2oyhSGU
jFwD9j0PoO1GsvdkWYxDCXLcmCOF6YZY6eoR6vyAAJW73G2PxkvJts2Pox/tyaxw
+f/ReAdaL7rU2hBxkm3/7xbApdCdUby0aLEU5J0gju8oFiqJGHkqsv7b4pLu/1L1
OsB/iMJ8uXRl4em9mn1/Wr8ibgi5BtXgzthrQ8I6B8UcD4HwFPuW7VNQq/6Fo/Al
KFEj7Z14O1Ws8rRu+fBo7kaacyCMGuowUiULp5n7aYv5QCcbed8kIEWWJod2RPYa
IYGzQMr+5vngCYANz5kTerZtd3Fat67z6n9zbtgTXk6n6NvZeETXb+MJtCRKK0M0
jrxbCQ94rjbpCR00f7EQx9TQ7+wu3i+KCWbEkLNLVLRxPM4MIzd2yxZBR5rlXd76
R+G75tqp5RWa6vy2R1QkjiNRA5fq7+eAEPznG5Aeja4T/6EgHDp2Ds+jv0Y+pDJ5
Sxb80ZWi+8CzJorwpyqTUQJurR8N4Xij5E3KammYxl78uXVvnRziX4ryKB+2Xgy2
zHZJp6QDkK+6+coYk/mbjL4hRNLDu/OqouaBsErfNM7LtToJHTbhPOwSD2FLUCGm
vVEcvNHq4dMkgAmJmwFA5aQYsMInq4arVskW1dFEQ5bg5azAGpb06NgAG9P+6g6j
y5cl3Flsdm/EtQtN/kEBA5CxDyz9LUOvFfW/6qPi2Cwesx4oaC2OEyYSb6k2dfJF
4F9GxPs7m4nefBbFexqPVaied9Y+cyaoxmbPqDWeeuGCDhuUo27M+nJmJ5X5+qjq
MtS/TbD84yt9ytJ/7qe5rOEjZL9eh7ZQtmNApa8uccIrvIdb9zdGZ1PG+ugW04MM
wBd9oPzSXIr/TBYrKPhT6E4Szzni8p3mqRHPveWWdago89ss69CsgZvFiQ10q+s4
ee7C5XdnK/dCnyDgXFoChVNKZrj+QVS0CLMf09fmjpCHi4zIexDXg1lsTmQY4u8S
8WCWIHRaiQp6d+dtSPzBZp474qViqDS1yORUN6nanRQPCvIgbUXYhobSRc4qxw6E
BO/9KN0mBpfi2FMatOn4jsvJAlWTDrH2DG8Guzg30c+UzhSmDREfVx9yuiezLYmo
PPd1LPzG8TgrWKsjSe3IL+NTwy0yY+lpFHjewmN98vtTk6WW2vs629YOvPTxcuaO
JE+LaF7YWGKkRlZ4npca0b/tgndKFkNIUEcK1RajiaV1WQ0iRGBTBXjaeA4PCnCJ
5PTKHB65EagH90QCCaBnkDedNendU4nEC+to0Q2kRcvVS2IdZ3rXiPNH0Hd3Vgjz
/mcl7274qrtnbPmaUsHl5meFlOG6YGARxz1xD+I4EXiOwkrPN6QSIrmsQsnzLMUp
R52ATkO889xpa6TONlizLK92BZWhQeXu/Y9Ko7hMPUMafw3zZaDa7p7SLwFsDB+c
/ssKTLtxoDnJxmTddx5zbhClsP++Y+frvpBDYdxJRbOxuwK0aKzn6HBBTKX2jBm1
vfAz3tsj+No/qn8Iu4R8ped0liTdvJRZT2eW/AnwpifmC4Bc4UJw7FYknnZ1sepv
i8QEDfdCmqyG8/ocUwNF0+C3GfYtRWtUFVAEDaiu3F0vIn4Vpb42xMalzfrLppop
mLDNafiq6/Gjt28LLdjc+trLlaw5KFv0o94mfAd05i78w3ly4PCFMZw5wboEXmjX
kXIQ9PLPzAc5HfpPN0zsyNPfllhGQzTaoGkuM6GduhoNJpN2gQT8ZdunYvahmXsT
zE1a5eiKLTemLPLbe8y51w3qL0AdzAKY9wXli9gHjEuhxBfGTBwMu3NC05l8shta
3+CcEN8voNGSIRZXmmqUpF5lLPxuXMMEdOsJi0prCEfn/10jkrIJfB6tW/WwCO7E
xsWkHFN1O7O3aFFaz6gDNGkM27xjlCXHq3ZV0Ghvax3tOaAIxj1rmLyrdYZBXNzm
acVHlAt2oI7LVJlzDWy17jAW6dlx8ZukruScHDa0w+LaOQbfh+nlBbDi/LUtlWc7
abY+9xgtk0OnEe/loQemT/7ITYku+JlEPE1j9Jokb0d75iXNopU0g6/QUCzBqqdD
aCD1GhduVQHMtfDf4CN+7OHjBcPnrzSYvj6melUrmVYLFRD+zFUySVnwcugz+ZsO
ErCmNcowKvzL3/txZLcvmrHhBcPkKip/VV/2phXcs1ZoH3NdXNzHa9lRPT+WwFtX
IVCuUbYOkq7fY469ZlCvb+xKCeg+hpgqegxHFy4c6WHZqpsOZR/E1xDUJzPUrjjT
+xuaXWLHfFTRR68YxrDPkFpKSrQF4vQiJoYK9rMgg4nwfpWwWWafw2F6Jn9kxLu9
G/+Cc/jA1ve6e9/Tp+V0nEw8ZvDUAAlRUIlW8Gbmscb2FfOKSdHT1EW/tVb8uLqI
Ra7QJU/bldYVqi3aqOvtL5fkbIbDwWl3mmm+EHjzK3u4/HVaevrEeV3hrX8RUC87
N8V3P7L8Ql8gmy+MBUxUkchGgAdg4nEq1vjS/YFAD3v8u+xb3W0R7M5palxqDSKG
tR3oj/WkMOoZwVg4ZOUCM37S+OqJ0oIqjhiXk4kuF7XrFlvy6UBJZnHJHNSdAkV3
vkG1t8OMv9ni+fBoHvV4P2Zc9NG+RfwS1SQkx7ruiF6SflDw3iyTEVqYGoqgi2v0
+ZAVr4231cX1gLhE/ObuR81GWG2TmvtvF2oTF36RAGm8/XlGYzZi44QJAooh80DR
DN0Rq/dfMU2z6/CVXh9KSHHFhBWWk63kjquBmJH2pXiZEwKvSLNWjb5vZYv/LkNV
nFS1SuK6rPtfSnX2cPzaoD+Qz1aGXP4CDHFgeOGz7x4tjsyLSyCME57bzOV1emT3
J5uIaYr/jdnYgUdQTLSp6rX6tfaQECkrPD2XB1l6NQg8p2liSAEJePpnfiu0+MPB
KLqa8sCQE5SU6Yqjrp8Eerys1MPiqARq2a/OX5uzPcWJ6Mw+nRfi6z+XXCRuIrPV
bz1eEy6g+Ks0mxLUxmxkqj9oGk+YWjtSoxVmNZt54v9FsV5xD5cevSQTpEv28PWh
duErx+TlWHuXZlAa7Ms/yfpXfJ8ntow0HbjzF1EA38JpAD9DTf87XeVcy29uRSKi
WWwJczPcVQ4PBrbJWgVS2ChoMB/ufIEyHZVH6mHrEidwsjcpGHfBrfaXQO/WFQZt
IVcNJxmcrNp7Neuw734nX8XQooZMVfvc9w9Qs6XEuFQkf7UGZ9AC7wb9JkXMoLoa
tl7eUs83S6i2bvxsFpIIu9xFR5/Biro6yw2hdMLFvsgoy9jqFseBD272hAO/T7Vz
8Th7G2EK7W8z1b+cQXVoOFa8TVDQzPSUYIOpmeiK/dGtMmUBCQ5te1LfM+GGUUIb
vbdbDx0Xqk+7AusX8K9MLDZSyZ7bKG8J3ZF/xCOxu+Atak+pgEhvkbwNHBpekOir
OossBmdaSkQ7ZPnct2uz0HN1KOdnGdPwMkJrH4REXpAPR88+BqXuS/bR+RJ2wERG
eGaLABUuULS7Fpo/hIYuYcXyrNztjXexy+Ct7WYken96TsVKSFz6qh1e6cy839B0
l6fTczsfo+VH+J1EYbPsRdX3ymQLK9Jq6cS8JmdPTvKmHeymiNf8dUbKbDT+rIUn
6kKJengCHntGGh5yyB9astbjAKd9fsWoFmz7clqMm3VEUVvCtqu96gBA66Bys4SZ
BKraYpUHB1JwDp41gHi9JrrTl9BJUZ0pWB8D2NeEy8K7pecdGAsj2Vj8I9/cdxH8
OYGDLn5lUqrV79GcTnRegpuueb1Kn/QpHaxmMdacNUllaQDYd807vsiZ5lZ+3SzM
bWPzDCslK9shWdE1OWUed3EMVfzEMGBz05TnEpoITvxHSJcnUzCPVd8HRco1O22d
iJ7uYwcO8MTqoLrBNjj3E3FP6K+muyKxLHyXHyIKX6OUh7k57tLwTKWvI3ZfOMQC
xjmkqxzMUmksreA0QvFAb5i94zOtFlU6nyYkjVAI7cPOuyFI5NWwIFc0z3vQhRm2
E79a6W8JTalNNaGIKvtvwbPPW3IVOat0RRoTDEb/jqvEBZh3SeJWBnqiNY+STsAV
5IaNadR1Z4ktZ2oluSd1h88Sc9+obA9Yh2IVxFGEqwGI37cD63oggyiFQLqPemoP
GYkHKVJmKmjF3W1+8g9Y+BjybGxPaPQE1HJttwE392qUOchmSS7hKBcbzXoVD8e0
WBSsfyZnBETTxXBs0ZYgATqCwB8vk7OHr/OrhhaLClFpgGoFYKbH35syIBMfft3x
EqIdwTL2WDX+l2twDkhTZO9THOfV8FJlbCRe5icUbtoAOFWouQHSNFfWis3H/7Fl
EwV8C2pCWttDScUMpIQo+rfNFzvU/qMHdsmVQguypfPWpD78Qe3DC9dxoxlFu3ws
x6Dg2z9uzD6dJFGBrYdQlpxyFSc4W6ubqCZEgydGqMne1prULl9buvB1vVKEFjdF
veArsRx5hZ6m1j9sN1FYnTR/uFX4mP7k3UA8hoGibSZjx5hxlSrhIIi5KY38HHLL
vaJpuIIDKQ4ZrCZ3GKtI10y9wy0TIfj0hGCpOCefJ5TQYqZ4VeHcYeMz4Cl75dhC
3zKc1vN1hbV/Q8zGRxLzYGHC2iySHE42WcNqfU343OUNDlmzEhYfskG8F71vcYZu
gScwGwJxzgPC0bRCL+1Ws7nnZjm2CJ14VsAZJ/F/So5jVEB/gfKb5lYA1KZ4EksD
EycyiCdL5SXfllR5p7cbeoWRFXIAthIZk8WsNNCZUNPX8WBD++LAWMNx4VpPPSeg
7OujwkVug4uVyB64p8rQ7AIBiLpCJnAKJL1vljNXymJNoDkJBRu9OWH0rbT2wCdt
IkcmVUp9ZsUh9E5P9BJ7XkKskv3yNn3LSoZO+jj3Xr7D0L51bIozJbthLbQTs+tZ
/xPuYsX9E+dJxE7rE9KyTLST6mKQlClSJt0Lqy0X8XUY/mZMgh2UG6JYwfzCJwUy
jIhxI+2WycVpI6r+CUiDnhgq8xGPYZAq1z9XHLwoRl1vbx3Ya1iotzkfwDGpvDlG
ewzLs6Q7LwmtWkRStr8d2J8Kp6nh8bVDfJJFCxrmW1kUPHaKdo13rDKK9FuvQA/j
I2XFKvuKEexKKH+NB9ebalXPxNpY+YNQtD/W/vIwwwusUxPF+d80p+DURoMleoq7
q0nsTFVHiN43kzET4I+8Xw+qMP00X+aHr4nHL17FrvGwQEADhQuQT8lwbxk32X5L
Ya6pe+MzKoxwbQtP+en8CuXQdutfnP/IxRfNYJmjAZqjjwrVeb4ZiKvSQL9vly7F
AHIoMQrVUFyCfO+GZlXbYlYM60cCfAxj6WC8aInw2Z0eCWg5rRtKtL9neSpAbc0n
gkbV/gYwmLTHGDmalTdNs5kIwvzOIe6wv7aunVlP5E24XOtSk0oxKlBSMHytaKeH
LIqRxz1ESekvLRbtZ/RL8wvmDAPLKCOvqpF5znA1tqCNbSKgb9gJ7gfqS7705yA4
xTQK6hsfqldOVEEJf2eIZ7g9gv3ZQ05ONSNWHqYAOe260c/TCH+AZp8PodGrT/49
lhG5gtkv14ih7iTPySgQP3ahFtjQEpIZMRfvMvR9DoZ+NHKegJMqcVzldDGfY6v6
MAmeucfz/5ectGxqn0jbUHBjKZldlDJ7pwybqJo6GCiURuxXIMH1h7w3KLftI48q
tgxi1enHotYT4LFWys3cozx4lQsUP6ECEoanDxgc/CVOCz3xm2i869SjhERAz7o1
cMIxHbbsJU3jMhl8gMwnbAPrArqXj8pFQIIxTaEbWerQjQ31eJ1QF8ok17xecvwl
ObuS3euYmtB7a4Eqij4UMzFFrCa6fgSPLXP9mSl29zu51SKxpHiy/dgYADVFIOVe
amc57EYgQQz/ALTaBTkhokJfsUtOMO6gJ2BHS8P+TsVHMQnrfe1zZDbqKhzExSMS
XBDifl/D7G9e0UVVXKZKLd3xjoPTI8Cp0kkhE7yA6J0NeVEjKzZfNXM81bdaZb3j
RA9HjZW40DyrIRwAfKDZcVBWUmU4vNVjH8ZySvj+YiLzBTkDq/S1ep6DkTfNJx6Q
mjJgnqW7MmW5CfKt2Yy6MXk2zlPFhG/2zCxEloM/dg766Lmo/JvjTkJr1ACEh1R9
zPC8F3WKOZu14hDOGRRwT9/Bglb+2eZ3S2MWKa8SZuIiMjTEK8XLOjWE2liX2X74
/3F0nP83up6UvI19QASNcLB4PT6TZtAX85w5LmQc3gzH3p2vnD2JH6EoK6nRfnp8
WG7KtBQv0qLjXOjO23jR35ooTcU9LfbjA1upf2Ii99sEQhhiHIsd2wVJMDPMH3vz
RYBOEYtQcB4PpPABHnpGB1d+iG7CyPpLhC640Csrfyd9iA3Lrq4jhsRgxMkfMw5r
ousJzuQj3A232TvVi3VlGNB/6lK/iETnOZcJn8MGc1tnpWIQmmDnXgRrqIyagMfg
Q6cqd4Uk3wT+uYSdyhYhft47L7+RumZK47UDshSDpsYkzsJPFtHxH3Eb6bpl+hCv
+UER7gOmv0N7iOzJ1WRTuqm0AYMqBcP2JWAzlbmUiX/x37clEtg7hok8p2yPfiEO
Ft3Yqoiz58BgVzUPpYMyIF8y/gLFHvO4rF8CTAua9iogF1Vqbqe8GsaBZuE4ZcA2
5IALKlkOOaqUpqom2tiPMZjQW5t8LLiX1SmUwMKS/d6JVAqhPDtLvFHDWu8x9Egn
b7zB7vWtUdM0knsgXFe2b+Pp7n0UmF1GINHyioh9Aa/HsikA9kTGmrJkiZA6rNk4
KC2puaEy95o8C+visrXQHxd1b+OGGgAOiy3wMyKHB/2WeNOdLDtb14WVZ1LHAK8k
1nMbQy/CeWcuMdHliufy2oCoI+2nhibjaedTdLzDyQhbDoruRx1DWE4H6cmd8YGb
krD8/pWRP1LjUcUNGph0N/Ild3/bg6O1468z5zx+PbCCMHLgcqHBEwvWN0s9Rk1a
iy2z5GXz0eQma+GxhPsNC6ktwxjDF08NA44yy/0RcSztgb82vwRLQo/bc0LcjaQ+
IcFUjfj+U82fFTdGa1Lqfh7z8XTQ7uukt5kDEhoirqgI5tQVbtCtdp9Q6BNNgRa1
ClHbpTbrW6YkoGocK2eK18ATp5FKNVdWWVmTAodlAbk/bg4ZZBXv4lLI1MOHQ9ge
iNlKW6mifCtwfNAFQ3/pSw4FbJaBiFmapqim4+3vZSFJgGve0nh6ZyPnhNKGtmgE
j0j4wOfVfV3ttWGCzCgATZqvCrQwONYAgz3lKhh8ARXWrC3psXrs4zjEmr2xiWpJ
p72e1tD/z/jXACjH6qoCjrbaLuCquMsXpGVXlCc+LUXM70AqPi8mFPt8k8nPoYx1
XSFqmXtdWeXfhgNT9iz4hbidrHW4jUJ6F+OTlix7LLk44x/A7yj8uBNv3QjaRDGr
rnwjmKNwdGtVRxS0UlhLAjOhYGCwii+Gdy8v00ykjgZxoaE+B+ILE0lmR9aJvKVB
M6MWCmX1yNJrom++5sDPzej6I7DEztASTSpmFafwkOKF5AbpF+FFdj3JEj3BibIv
TVcmqYKoUo71A+F644DcItBnsIq8a9nmK/p0ZyugYAEGykDPZPVtU0vublDvD+RW
juwq79u+aDDiCMfcy13PkHGbsKrAykvhLBS9jgkZAPLOmtavdUOaZZoh2LQi2Ri8
l7aHV0lbaJWTixIBkDd1HMKd4/vMJw/lsnJJVjt8vFGLfsHzaGO88W+3rmo2crRH
XMucSCy9f1IGSOP9ax2Eu8ftTnhkkE6NCWlhA8tJGdo9RD7qI/f5KFxSXcPxHn5F
vIvQAiiYGnqaR2sDvyNlzd4qHluNTXnmqFleTtd611FKzGhWB83R36r8gLWFwmqc
YqtIA2jMMkRqprfzST073WA38LiyQBHlnQfs1Vl9HLYTzNTZ2ePx83ywt/p6jqEv
2ZRPtvwE0CW+1fid8dOZ9hwpacAMDJYGNVuaWZrECbz9vHjxW4R6Tv14cvQ3sRZI
1AwWO0CIEK2ia7Kycp++SYOi7epmxa115f+YKNRUyWK+YGRjM5SbNOykEav3kf0w
6a+RmytIWQkR4+5hI0D+LdP0oJjauDQoult4JUgDcrTiD1nmobjjXMg42eUV09WS
3ZS4gjaDowHYUS2dkmMKhMQzqL+BSHs/NX3/BXDQbkxq5GfVY1pZXNHkhrKoD2RV
f3RNBZSQYIpJH26nM87n+PGbbvwF5z84lwj+NVSlsxdON8ZTisIOOm3h1Tb8a5Yo
hsSgnDptErubY67+QfLIW/9O8CO95qqyOd02VRHerGi5a6VuIpanh+fw1yd7Lcsc
WdQfFEO40RAUJUb0yI7n6Fi+ehXAHgxgVGhLjVJJlQ15YJaCEGMkzbtLxgp5e6Ts
nI+RvUPKE30wezWf5uAufez0OXdpfbwxQj/B8ryZ6eo23hVhY0jlIKl7734+G8PN
FYcg2dTdkDjAWKmFLkxc55zld+6hbEuOMmVmJb4AT9QKPrnEEOXeVd7JzKlJGl6u
2nP70b3tds3ZZM19PalHTwJFHtJEkiKf99JNPxRizS45SWcrx74UXOmLtSMM05IX
N9gkQz3aGbYsdU6X32hBLCkCqvOricsErOld3NHVkVmbeciq6lqbFhDKMtUht54X
MVggoHfj/rjtkdqgnNlsASf+HM9jJeZrkrlWXgeeFtwIvGfrvmmJStG9T9Jq/8XJ
N32FyKE4KsjhNstnBYdgFm8PbW3k/QPkvFGs7jRxK45E7UHcxaw9ov512dgMHACo
sjSDJvtzRS4rRQzmxRKm9OGCK3vp38+zlhr8JxA3Bcx1nYeNVfg/1ELYwbMKqGq/
kM5538/W/cClr5+yfJTxDMrD5cxKrtlsJfwouLUCEwCS3I8/QqstNQghXOwPhfNv
jZ489uX/UUn3aEgQZ2FXH+ttiFVp3syrxHtGGK+9NtbPe0eNZ/rxBV7hZ01d0CKJ
nDSs+ey56eQmt8E3iHO6+8emoqZPebWpr6ZL42dRLkOk/vrchkLx9QSzrnwhaI1n
9z7wE5TFgmuEh2lCywxKp2cXCDVYKvdexs7m9/IFWMLftiHq/cw0oGuKIBuEDdDk
gnJuRiyQJKKznVb1Lv3QKDIDyHelJsgJPig/BmmhN/eApXaLKg1AY/uw5dgYfe8J
pgOYLiB+zLyv3OYN4VoTuLz6crYzqY1J+YQEiw7KdIgvdQOZJoCD/UK3pSNMR4N7
Z3g2atwtnPsmvkfyYXGrNVTDxhlXIyK8iqJDHXyE7N8rkof7z6HXzP3EnENHSQsS
O0IkkZgdYAhBgC+iyxv86ygLHhN4VUC9+AB6KNvOLSsE/jlaDAAbadjqiLQJ46o5
c/7YUSP/FN2FyB9xAtCC/psiUpyVkKbZYtDAJwL9hXiYFMS4p6/pR4Qo8231xGot
cFfm6z7gfAwcEv72ecZBhmpJcFfJIPWixnRMUSnlzAV+YL+gkEog12f2H9fGfuXY
+xWR0KePyTRWILHA/mZtt1E40eNw6pAGZs4g+0Wz0knViBkqTgLMlIU2EoeSqIL+
P058NZzKzMshpaqE5P0ArK4fv8bpzOIpV7OlmUjZZMU0+XaCzi03ejjowno3qFon
jqBEj0jo5rg5qdEzODHM5iO/1EjPsDOHeyTkb5xzUEAILknJeSMN0Kvm9WNq+jM8
MonOy8KO3AdGFL5maqSTUCYXTrBrEwzpvJ/+T/2IeQY9qpC4RId+EAeOOhg+MaUA
+++N7wThy7FOjdQUWTgVazZGGoEMFxQQ2digpzxEaz8cmdxTARSi1cTT6kz1Rmeo
rpZ5UeapJjyd4Di7vJgnfPRAfX7IKTiF5LVYGoc/6sFt1/MB/Ms7pB1nPFlBnLiB
NUCMC79JsDtCe1Mymy6KgArME1J5tnKNK4f3ppbERsOt4qhEqr0vca8tA/URBGDm
SmSB+VsZw+l0AC4SexE4bfAKPPwZSzXYNHslDd9wEXJBfbdh66r9u7rP/uboUehp
0MQRS4dayObfScFOsGwQWnaW9kxxCkN4fBeGreR2e0k2lqFdXyA7uR24Zd0qLfRu
q+VLrLmXz7UZbro1vlo2p+B6ibHOH/pJCAqaSOX+azC6uGmuI2+nAt3y+tA6QqYG
MCAWoPczvKUMC2vBqQxJSSm4OW1ZqPjkNt/3qvbGX5Rjyq7rPQPDyJpiWp2FsnU0
JJobXvcnYGYV78GfM9B8QY/h40sQGBy0ts22OrMgI3EtiV5nBTyEm60xeVzGsga1
Q789Ufb95yVdpy0FlvJcnrJb8VJyvS/3AfRo2dMIjtOq2u219UujrOBZkSP08cEN
flqsL2PWl4PUkwf+xYL4QldoiF6+pqZMRjR94wJ7PGKfpomFdVrEXaPQPpy5tqme
Uzl02jLU7nhbkeLq+Bhnva8zNcbIVn39Bcvuc8eWvXVrWtKUGCGG5vYeGOSa6iPJ
jXLAx5YUZi/XtiNjnpBEQIe6dXJ9egoHozTU9A6JJyf6/o2iJDQ4kilenR2kuSXu
v+oILY2YObnDypGw7H3+1RdNg8febjZX9EQ9cPDwnPWs5MTfsgtHIAXRDDva3d6E
EmLv3bgUyRlG8th9EwaPkrBJdawMknDQWjwAlCf6LTE/IPHUbqtvwAsouhA5D1+T
d+vs/rIwSbBQWPTXxFxJ/KDBrhteYU0fauz85zgGvXf6QGi0Ry/4EtBr96fmb5oU
kgDzoPyKnnE4NZctnTjwFQShfnfRssWGseTiQBkfDp7QqxJFJ47WUKnbWcXzM5qc
wzsIpQgcm6kjVKmMnUpFIA05xvM+ln7qPKM+IvtxbMTIe1F1A6MEumwIAPXt3c9H
CbvtgDKK7XVA9NFSAL11eEnkuP9fqQtmQi/FxjFUORh2h4Le464u/mTEqr06oiox
7vN5Zo9SCEBqfRR46820Blqrzr4Ea5PwAcLYys+mA1v9Mvg3x2W3PeOJgRTSZk0+
O/r128BybVUvUCwxxCm2pFpQOTXW8aQGdtuUie3egF/7nv3Q7DLjXzAd4UgEo0A3
H+bwVIHAjpOrMjhgwZ3kGwjHr9l4H98Bo+MmFTV3Mk5T8eosOqAGl/g4HwhgFwZr
F29XRseodGCYFkULcrt+WGv2FjqoOyFry4ybHEu8zWlSRkbepC47JaPspD3SflS/
ZQi4Uhk085dND9vb3TIBuh6UrdY7haynLVgVnxKC7j1eht5EEooTbKY6++AwiYLx
NpZKETqBytXx85qsZk8CeihhIBSwIagzbIPxQITu8/vMAW/n6ztk+sBuc1ycsK2m
/wEvpWzBu2uOiyB9pykkJ4P+cj6JOvnUv/wRIYoZzr1pgEd71RlTC+w9heh/1R34
4CiGTfoeirADw9q5wKXng2arS0djnWp78E9O5Tlk4ESxluBl4Ww7AJo6wqVT+/KH
TnWsazKSNqgwcSxbf3ZRXif/ARRiEXdyuooorKpKDVLhCHjyeg+oJAWyoBdngepP
CRPP69YFRgmhnL2fz7Yx/WszTIj6KLYfM02blvxs6+0xvdvlRVAo5Gz91Quq2e6k
hPQ1W0nrl9zoCumvaEJs292V6fUyye0RdaII9vGZzVUO4ZgRKaGtp5G0h9p+Jr6s
I7yczLF/ZwMV8kjTripXlsQ0LX4hA8USb/qxtq3QXG8w0YD/Nrdhgg8QZJebHNj5
9njrqYB6kPxZS/4CfW9FGKkrGCSLKDGxNLksgFmljISX3fnSmpenk9K00AcUjeuk
xnZjf2RapxtsjUlpv/sKnBetq4YWVS5hZ1yzTBLEfD2H6GlhRs9fwBrVW3jl5yk7
mbwP1nsO1b0iL6ahpPjsxuue7K/kNVe/XCvdOcCmjYUAdjdmamYM1b2WoBbuozLG
UJslHpV9EsPWvoGZ8r59ElVkoq+MPVutPp8t+j1TWzQszsJmJuKWXPGQhER56m0E
55ERDuFAJ8mheah8j8enXpDtdi/RbXPImWnGuzWUBJhAx8FgRRsHaIZKbYmtxJZI
RSO30JPM5REe1vuRDDxAhTRAXBy06ll+gMLozNpovD9/am5nlPvANXiJKeV/7D3s
mY7jYUbVXzKUlq+wFZvBaefVxHz06duPpV/FhDZPyrTHo9eAnZ1OPab++3r0eUff
w5LQ+G/s+ks0mD19b9zXf/iW1RisVouPn0UFpasbnWRWnHTg06l3kOzJsmW7ONAH
MtEuR7VgNO+/yuC8UF8Hbn1a5vxM0K9FXcoooq6kHwSJMGc5rHGsaw80qOUFvlHn
0Q/mH7amT0XDExuXiuT6wEqZA026f43AAgnEE3So7KQ/98LZ8hYQJ18yZykYv4HG
K2xWspym8m7A45wyTiuwEqWH383ByRNOjYWOaZWH64ZoYBvGhmc9wjypI7hR4FnM
lQCxGt4X2hVT8XfDWarI7/b85w80cWAZbPd2Fw7tGvdxbR0jsNCSP2H3Nl9PqL+7
yqLFDoZbrlWapycoSFZcG7MjoK6+fq4UiZEs9lc+eVJ7SUI1lTIQ4nQwM9yNvDEb
MDB/5aUNuUIWzNOnmDcagf4M2kOfbt7KYaqjcNdna9Zu4YjaYb5BkkOahvnvs2LV
/1sfLdVM8vbCwtq1owKxxTOQiHJU1EhA8IJ51MV3/rYvgL1Rv5Dt+ooPQyOCIZuY
IomhdiwIg45L8pTNBZZvzcuL2ZlAWUZaR3TA+9WXlvw/awlXq2PWqnmW4SZtLUtD
yixRX2noW7zHLCq+2mVIZ9urOLTfs5w8ZF291ne9N/ZNTXPHz/bljWhyc9nU5yzL
eCQ1bvQGI4+M3iewR65+K44xcZ5MZx6y78NYIA6JGqDYN3FWYFjmr3nQg8xH9C5/
rOZgg/vjPrGJsPPnIHvs/JQroNjgawCKSjzrkYEom/NaGolLahnnWFQs+t+LaGGt
hHKV6cpJldYl9anfiMs7BsdUJ6xgNGwqFywc2sHJ9W1EAVU/CJ1UG3XVAhkglLdU
4WKFN4uzg+TF+923OUoEjmZQqe/+TLIzQ0z+JO3/it080ia9y8Dr4y/XjwE3HzMH
3UqZuAKvcu6x69BylVFyNsmuWlPDaB5BWgOZ5TF/aiOvB9+r2JNv7rTY5Gc5JCSu
0B2t7y7qPZWhW/71BABCPicVf4xLBV+3jXt1lpL90ai/D6Bs1WSkf3JTN3Ys4pgG
+q5Dml8OXU6XsjmwdXJwWi2rtvuXTTrYvC2gWO5uwrT/uSkWfGUSICiONuF7X6iu
PfNdifdywTwqnUnXtFNXwOY9oB4Uc9IMzOTfYj5woJSJO10Py7b5IOkTjC3rPrQH
iygf34j94vJ+iLyoRsHzf8DhZO2689/FczVkcef0G3dAVChRTpvByhwqINg5hpOh
yVIYVga5/nuxEVmT0owqX9VGhNGh3LrBSuyn/Hu/7IzQJGpLRTPdHf3dAfClemID
xkNwwtScBIyF6IDZrU/S+VUaYxLCZu50EP2yo2o9w0ixsErCoX0PSyXU3ZXcS54S
eFSa5jfup90FuX/j5K7vN3ZW7eiT1HTMtfeUZ7wHXHdigVOvk53kwywyzQLvkw7J
m6itJMVOLrOSQ5Xkcs/Vl8w4J96pfrUe0k+eYM/ERPnO7OfAeP80ANNxQPUADBQv
K0DQbF0WZiM0F5AeGIR7n8IoIasYj8Bq+RdNxGp/svu4jufWjTunVAcBXvlj8lnn
kxvpl24nh0SUpuBH4qOm07UKWnwlPdeFl7kFUFIBj7AfFXUPlnGRVWZGR6rk+yMV
FTjITMf7D3Dw9Gflh6QI2oUTqNpr4/PBFr7yoL06zLIJoayo5EthFL/SV+7iXwTQ
EpaNOMJXV9E7cicr9SukKf7N8oCU5LO/8+YZwU1yrqw63LhWpwRBdZvPTgb1p6Ok
pYoT7fbb3tscm0fI40dt/Ypr2A2NlCfHDQkmzA6KJyc0FWO4X62720UdmztdeCtz
S7+fAxSHmoP81QyMtnU868hbEk/IvhbENx6J1MhplOzrJgpyd8srTw187J5V4MVg
u5l85gsYf2O2w7qgw8/6pZHnVS6HDGW8lzRQRuFfPt3mjE6tbvAOsBDMIdqFiepW
4bVO2bJnndm3Qzw7I4z4qef9XS9I/fXJR5HYAkBcI6u5Qw/nCJQOYbcekzEVFkqn
6hRI4z4728KbWIxYv0hskvbbz+3LpQoPGObeuc+gzXfc/72MFBcu/6OImEST+/nP
S+XgQ5LWEU9E7GWlo7HCwxdsPzKbhz/GKkGmyPsfBBhnVTZrO42xCsqPVojlKwq9
KjHaW8DyTDEQyYvLD87FtrsSWbJtk0An5ByREOM6rXYbqXpm/LRgg8JGTSVL7Dk8
4avoNs7YRyd6ZiSv3gVSDBs6YTVjSV11ZrB7eyBvSrNlhT9sufgRNfMryoQAjE2P
oNNmubxZeueemtFtQuc9u3ce3E5TByMFSjMXNeSbQuQwKq4ZEQ4Aon1Wk3Qoirjf
NFeqt0JQ9Zd78AZtQTBnGhqY84njDXvHS3cC7L6MjEqHHj3DjvD3t+McTknPeUuu
+ZnvfjoNeJo4LiDxxirDlUFMJTzKGBYOO7zhiwOw2SS7LgeTg1uqa14gpwlJDGh7
bQOsvGjyPCq59Chs4AchLSZe8GAuJuRBBpJPZnuAXIwWRndIQ6nL3+7Y/xqX/0kv
2R40FR10LWXL9XZABr2DQF+fatusZI2EePkAJPfN/fSrrilxtT4/M2A7tI4HBZm8
pr7SHYYYWFTl++zs/tYWE1l1DOonNY9J1pS6+ehliIMiBJQJaoL5mwlPC6C6Wj2n
UxWJNOSmSlbFIJMU44nfCgjvflfIaNgfPt9Y5uAP5xrltSCDgkrYfYIMhNduVjMo
bcOyPalv4keMl30RNEQYp3V6i9WJO/BYRtpY9dxUFljdWoRIezq2WyRvRX7eTa9w
uL6lcH3XtH1PijRVMxI9+zhGXgnIGG8/cb94bWzGascKwOTtDSU7fFXb+Hfxa/Qz
n1k7YloS1wi2ktb76YzU2jhWIgK7fGMSKuW8o5VMDvUoeOzLm+2H1ZcmP/9EiIWi
SRnE4DpJdI6Pvxagn/7NwkJrpk1RFxEy3ZW/sOdr6pkec/o/onckwot79+BGKZ99
mRnQGEP/RjJnJ6nfqikhDrP4h8YpeeD1Do8ixCyCDjHKYwofDE54AXIsxPmJQbhU
zEPDHL8020yyCf9v5JiVsoDcDZAjhjKGOgFp698nKfgXAikEvaVg3k+7sMtmiiMY
/FXT4vFzohluoqm/tj4aEwBuai8ZxKasmdTyHuPhWTdqIwjqM6M40W+Bxgt7LLif
5ybRp3J/GqQXO+ha/xA+DZtQLaKjTpD4rfPWvYqMaCwTJ5evAYVVEwgCjUhjp3MU
pk/daUp1UF+Gb6VJktRWohV5IaeoIRZSrLvAEUkZUcfP7Ik6g3VzjW4I2VUnxj8K
19pphPDLmxAuxTODnZytj5PCAAkGpfiQjG00aHGvh1ADkInPaRaMxPXO4tmEHQB9
yvlr6XlPF4f4SgVKNhwumOJOCTYhAalQiNz+i9/7//7SpIVMV6wyWgjkQeVHlrn6
R97MkJxHVLXgxCkwfMl0PiWu2HuE7IIA/1qb8B6AKWZoDx1Fqc/syAdTGOC0M1E2
xoWbfn6zAgkBU7hd5fZyAmmwn52unWw1xyDzuSm8Z7IYq0MsN5xTLGmCBijJ+D+u
8Z+96yG81fzs+vb/JLbrDR9di/+or5nxQqjFcQdybAQMUYyD7m+zSOqlHOiWR0YL
tgkYX3LxOIYHVDdwGzg3f1Ezhh7GDv3lXLxbTaUJRTLCrxudb0K+IXpI12CTr5CW
PUNOMDoy9lQLWXsZxfRVmIbK/C9gxdSVnpAfxwx6GN1hTdGsqHuWRDiJWPS72pFe
PDMTpoTYtp26vAwyr2Rws2UY1ZTenEC3rwp0hvKyY+8owaY9kXUwJK5cWGoagb5q
Mcfq3Q/TTz9gIIgXY/GOWlWlaHJI2ARCHmzG9xNCT/+JiNuyRFMoPYcKQSQhvcoa
O8l33aAqzuRzJ0blhuKCeNio8wAgLz8nwQiK7riNWFmcrD0WqaylT+e042HDFhv1
jzwBcoA8y6ZXLr0WZIGFtqTGLP3nRv5Hx9LemBMQsU857vsmZDHq7gR3Ox2M96JT
NYw+7BlGHIW6TEHBwjPOhJZDSUmhJXQxA9/E+8Tau/htUVxGI8DrgT+H4+RLhjPG
c0hVOAvUCRS1/GW27g2CIFvKu1EEGnxiGyhVYC/2kv6XtdQT1989GmMHYhqvoL+M
tLRJDd8NtOEEyfP+ZzDwQ4zGrf40xxCoikTtny/nWV477HLO5TZzBoceZyEtPqd7
aBVbw97fGJrZk/LI6bAioItQI6pWyHaaiA50c3hKocJdRm/w+thmOBn044AO5MRJ
+ShGCxsB7ToiiB3L7yitl00mjZHnalAZ3R48hgTBEcXLH2uRfbY9QmPjX70FgGPm
7NCaApDuRA5YwsjLKbFHzvj19+ZvRpvolmfIeqTP0B2tedADcHEt2D/JzemCeo60
IVHpChudeHF/IlnUHjGD8Znq30s/+UI8NhGVo0kM0pN+Lrr/Hh8oN5E0diJdRJcD
6/eDYvuTGKmKU+DmTiWCjZXIqsiM3VW9E/OYhwPkiHAnjyNmWr4tBGlTfVPAqIGX
xrS7SVT7CWpsCKGlot/t38NtEfp8LV/6HwYt7PgWh4N014sRT8PjOaSVuyIWCx1G
Xgu16g60RxBKNkHqiuRtlszB/yHH4czSD/vnN6EeBZeRsldZdhS+wSDn3JRvHnvN
tFdTLagXdS11/MbqUhCRzckurqbO0SQrwhSGAr/zMAtq+PSvjGD3Qkr+X7v1OaC6
MiqekHxOgq1UQ8LCYTMMhg1vRbpCjixw+Favj78OnUVrYYFNQjCv8E5bNoLSme7a
LVqNJg2+glRr5hI81ZPOYzyN0+XcK9Gq5Kt5nr+SNQoo6Di50D5STvBiPOVUlicn
TDM4GMvF/k+eOWzwsCdSi33lDng9lC6tmPBKHVSRMMWVB2DGIp+ReO9u2cX6Exhp
jxPTPpXcie+j1HJDbMDJwmv4dptOH/alpbCq0MkvernxJMuaY6622nh6gbx43pl4
c31r8KLTnJyWJ3Ep0Pe2k59YqJszuWe782T2/0HvzuJj/diA2imZeZQHQVqicxMi
Isupf7DyJRSMX9Tb2gS09qttvTAXPjZCPeGuv7xJEcw6nVePUFKVQQ8Fj4Uz54Wk
i0n0xbLXLUH1QDd3M+uLpfcgQ/MfN4lorj0g4kq0ReZcM78kwwOdQLd/qN9hVR/S
M4M4FkavTXCIDDrn/aH5m/O59KjPzV5OIs3CqeX/C+oLIM/TNWRjTaYLhZ9KNXo/
NN5O/LpIFyOCCIDJFH6RTMg+hi2N7cuctFFXQtslt9rMYwMRM1Hxsjr4r+8uKxS0
+/pBh4fciGgFceISWQxuBSI3OPJ0Ks+u7Gly4M/0KtI28sTQ7cZiB20GWYDUKvqE
ghAKWKcGHkF/yXa+oEVTgdUR7nyvSBWrdStG+45xLp0nAf4gPf/qPg79y/8ArGS7
Y+NppmDW6Rn+M6cUqQrdzYo7eNctQssn/8XoBBBYCF3K2jDNv5SZm3pMak9tooQk
dGmfK/TlLZ+6/0bdZrzfb3Vr7NimUeHtZuO0FPpSS3++y2mTY/92eE5yroWvDyHt
sNre9Dve5NgSnGJ2e/Jz/+bKwX6qFyFoXLRdXSOCQnGHWNHZaO74z5bPdbglpVYM
MpEiBPMfE7GitS1Xka19OfV+56MnYtrvhXPmbGz8pKwcb+pau4CPrYv6lIZyfcXu
z++OOWhi6WFMd/f9jc3Hap8GtYM8a4d9EwlRxMPE80FompByqLX2xC7EVYfJN4SB
kNav3Prpyiww2p8cdSaJYdbMg5wSQy8+SSyHpP0NZggpT8B6muIuMH7Wh9gKpj4f
YhNkqaSEN73E7dgIdKXwUIuckTZ/iwqhHZyXH7oo5nyI0aV/sEtlER5t8FM2/6f3
LcpRhIbHjAVDWQlWkx3jVsKuhwLfvyzdhQuxbHcxNOYHoPeBhdWSBXil6z3kjd2b
Y7aE/xXu3eNe2gXn+maYNvWR6V2wleUDv6zm5mSXV3POV9uhB3NQMlaOy5Z9iUYK
tqR14B0jW84+WzKUDhtjvDmjXhRbPWyRf5IfsTAGwTGF3i7xUfKue9RIRbx6fHNE
PWdMpQm3NUX820H8jhVxCQd+hKxpSgsAXfhxAUGPeDi+nqDbm+zF25yYykkLoTPl
KfVFoyhMhJAVkjK02FH7M+d/zH6wu2vyRHdjnz9PqsLxS1YYmifyyr8gkLv/H/40
mt1UCMesFOvEkaCNANVQ8xY9DFq59Q1pfOaIyyql9dI2FgSURc9/+4VWoIqypLGQ
ET9kZW6K9cn3Wfjnf+kTDSCMhTAS6ri30OBQwoBvDWOpMbKdDMsBK6vXzDlINhlX
WE2KdQ78scMHArtk6yDSFeswITx7T4ZY6EfHGkW/sfJUrjBRpi125P0PijJNC6KR
DQi3KTJ/fdbjprTjZkLZHvWqidnzS82H7fFNLABxeX3YqKgXnydyarnC3O7ckgOd
9Uh+sZEQZk0Ry48l6ssYA0xg38US6uZcbyuYIWN8f0LFL6V3V5hA3iAaU1gg6RsO
cYAYJ1O1KZ0+uwooQi91r4ROjYW5ObKT4TqaYFsCarRAtTdQ/4dQoIjYuYpfeE9z
cK/pwadKm1ZYK2F8a3kpRxBDLGQ0EXSnBW/R8YR0+PSQ0nMNtMOD9x9WLD07R1e3
lDjQ1oLfmvb1j7JxdsNa+Qa4Kr2cdhmddVQTk7otUT9r15T+vyotymNOeKsUSnQj
xs6MV4EhArtS0r+50iVwZ2sYmKfD1jLHUxdEeKvFI0AA5bxOkBVimGdixAWtIgo9
KSkfhQhe5xcGULV4Z7fS9cMr633dVyqNgSlYdUVfpSOQzlfvluRUzk1Pf3A00KCi
pWBK/cwqtB2f4tgQNtP5tJ5QEQc9W8g2j1BdNK67VVmI6JDNphA0kUoQJPwZG+X2
BkZOM72/RJ0lSfebu15H+PZOuUSg3D4LC+TaZKDGiNB+Pw+EA8k+aBbrTZgHODsD
cNY+pyNkV+NgG7d/o/Tpk55OconmDKyGZt3bIxMJEn9RkfWKvbDGjFmK1Rnc955l
uzcC0eEdYNHT2r2odpotmrJxxQ/QXKBqJne7MFrK2Gx7ZrLcx0cw0LCL5bbtl85r
Jy92wz8mU9iR2QnEXhfctY8ibi/g0EmkH3+BCBh7d29lIoqia86gG7C75XlOOWyz
O1xXKmzvSQXvg0JG9plgLfyjdMnjkKkOuQWYM6e+hfCjAir48EK51+KTb8dq3hjy
ZTRn8SWtPNKmIO2q7AhNzOxr850u7fsyKwi8t9GtdQrXB16E2PoQ6KKzgbR1lnd6
sBHhVxs2vdqMzrA2m0MyTwUykZoVHlVhiOJvJ8zSJuMp7aoZY1m98QaZwZAgqm7t
3enoVzA5T71MQEcKag2I8cdjOOfGSsTYfV0oH99KMVM5msEzf4HCOurEhV6NP79Y
LkI499fX2ZFoX87XuEf6XWHAunPPH0mD5Drl9n66r7VFn2FFM0ilnUfz5n7ouxzJ
P1LGEbvsQA5JDr/qB2CtIbi7Ubgdglvqd9heoNgGVdWEA6rdBaKKEDA8b8Annwuv
JaQobMY9/u4aVNCj5k5xZyA/TtzteyC3U2z6VL434mRpYxOdUj45JiTDzwG5Pe0E
vy1K9IGwrCpEGqovr5PYNJv2ynEIkXKSYc7vALxX0Fp7FzbU2FAwGJVt+6KzL4/v
kOfacZYG4v4YYnp8sR+z0aPWKYafim5FVwKXsgAzvjQ8PUVM9l2he3ur4AxL4YtD
qsfHbk8H76y28Ck3k37QMAqyuLZL+FIHu3WMGb9H26MczK/6/Kc+omRGCTSbAcQ5
dblZUS1x0/6AA//jM847gI4yVLCPdMInnsFhXjD2BmLawkOkusYy4GvS00x9dzZt
epaBPHpGEw2u3MYEpLsXZTI1hEHX3J9C9fuIbjZgNTp3nFErue+kfSICDWg09c1l
Q58NDRaYNwY6SmeGnRFbNM8rutnuNACBNFNQKIg2iuW263V0f5h7h+aExYRW3zwi
YmJqW/qmQIuoTkR66DpkUZpIZ5KKFfjH70ac7CiCvxnBLCw1oWwfelshPEYlY1b1
BNfBkAJsbi59m+DWDRpgivIj1OLuSi8enKfjS6dtCOkmtGalPxnVPU9JbzifhG/K
WkbTPl6eg0H+pCatb4l5orWOAGxBfdxwAj3qCDVjff5UQzqkCS4rFwgi2o3JMw0b
/cNQSFwv3UdVVzEGsYbRY9NO86SH0GGfuyuhhBZ/HCyxlQW7CVBja68xTiFiLqVU
nSfYWN3rndG+3fNKVzHCTquNhNK1z95eGmgdd3uZMNC/AN9mfMksvV88Jwe/IZc+
mHWdbrqLjy1oijMeKngC5iaP3gmCCSqwHq37HLv8jcjhcf0ZwKNUgchJ4HzXl6TH
LPrpFyP1U4vT3NJSi080yQ2rCS+N/uVN5JpEaVau/D0K4BLWLISA5bkRcGhFjDZ/
IGiReQVEW3mKdLeGxzysW7ypPQH7j9T7e+MmWMF8wI3Q064brd6M/tX5SIt+LF2o
imqYW+4gOiA1I1MTRcBjW9i/lE5fGTpA00yh/a6lt2pN6P7jVEybMuZxezC+5Jrk
PxK3tMTrCZQLQaYEEySjPYUUhASWOsMtH+DTovCngA57cEVh0e6KVPaSv0K9gJ6+
t6IikwXlNo2vy/3gj+GHJL0deyeklayXABIy4SJww5hLbLcQuq78P7TZCKjN6Reu
kp+ZvK5CYn9dpYysSk0r7t8UuEtvjC45Cy/pxpPXjRe/JMnXuXDj/bxUitu+chim
ZGUJGaCpeb0inNrMsiNzShZZDRl+o7vIdvCbDdK4V2j4LQ4Y5z7c016Lxg1kNvhS
JpVWNysivBlbYM4YpA0K0rT+9cVltCOQl2NqCwaa/OOsm/7atjHzDSngaDGrDgfO
Cz+9QbcGpJbi13yek2w2MNxsDBvMGzvhcLWo8GCTbYYl/5x26FHRXwfMwHHHsolR
ylzUdkV5PK7jqm6CyEBphD+jng1woSYXDInHiR4/auTBmpFTUTMyK0A0QyT+RX3j
iiPbYRfC/j1gjjnDJucsb0KHxZ3AfhVz1o02OHPUU1QxA4Sl9H90OWsVKkilpmv0
4ihxO+OgEGP8zVEem7M1EpH+Ka9i0SK5bL/RWAGzrTBJBjyv3KHFik2y3gIdjie9
W4mPw6Wb8MeEhhVuHMzsKbcLD23SlDhDgvf0jd/efJUvM97TyaN6GHn2cIhZXgB/
qFUUCNGqjB2FKXL65rCxILCIBbASNOLu1hEXyw+tctxcCO0ySmD2pl6Jq9bM3yTu
PKcsnxj7OsYKVnRu4f4g3z8U10/X382sqjrowg8QuIcpE0HQ18gioVOyT/QaEyXI
CMBx4Rlz+9tkqCJX9FpILHxFz7grReA484CsqGONqGkG/94UczOcw0V1xih3LWKR
uwNzi7GKYIPhsqISYO3fYGozZStSumuqT/5lrpmWaeP94wxUxZeC8ESp7XHGST5i
6d4Yg0YN1y+OZkhvtbw9SB7qj60SvbDycdPd2vLb+7XAjtDVrIUnCdZ79DPWs37y
WKqbAFuR40yn3jVuLSW2yXNjpGJhrLW0GSjRssGSe5f2LDHVoipulj//O6VUjiUY
nDo6/jpjbqgSwYvll2bkl9fPYv2jZBsF70ukVGXDsK39eQ1LBRBiJ1JPVS23rya5
xypAhAZkY6MA0M/IcPpHazOEaYfcZE4J9SbdLUyjU8dz+IidosD+XaeyOm3TfzqW
q3V+xXjPE3zQCqYmx5earp/hgnLQ8Zd1skbo3Fyl+fIQAa6LWVlVHS2Rgoy0gmE/
Br/UGvXQU1WIR8Tisx2HpVVRmimNIQHDrF4+R0RXYgxEoTxM5v8KuEtTQfu/ThVL
0fL8FAe6GR6Cn8xfhP1UHgHvG++VatUMVYLQxwMcNsVPSl6c+J6UkJj8IGsIW+P9
XMuq5f7o0EWLyeLq/no9Qfa/sh4kzNn+Qw5UaiepgKjofOkkoDKNgoAan02IPXlh
kiJ4P2JCg7dHgBluEpseYnYlDcV6WFpMrCDSGKicPJXORCKJ6um/1Y/aKInIqGnB
Pzd3ZFEQ6zmb5s0dV3M77gC9fI6hIGIsum44Fty5L0wS8vmYWBJWe35Sje0bZAjs
Jqv7oLTB/UJGUrFOY8N0aa/GdC8dapwDsCJLli4Fz9fS6SgLWp3oAciv3cigthWx
zMavK2KQsDfS3Pr4alv93i0huB1C+t/1fJlOMCkIvfvOEfrY0OvhvyS+gui80Ydd
Vp0j7bbBx/FK8gdYmvnbj2wyOUdDY4Wty4ebDMJJH79NfoHT2sSTdnaIzSL3l/8t
qZOGgGGMbddnaE2obGWX1x6Uzf2M8sOaSrMIS5N4/n2rTIsmU8xFJ1+q0o0DfBR8
/+zOOSsRdaS24YVVIEY2zetWqdhH+vxLzOd1aU+gEcnnoNv1dvAzLsH+XJp6z6a2
OQvtNWtBSy9dB30hL6pk449539bYlFwPKsmervCVbr1XHq5Nleh66uFUlD3unF+u
8i0wcSCcDcOpGNlhLreGHZ0GzOLRKuVKjKHLyE11S/o9OrM3YlTTusZcZJqkHsW9
jzsbrxTlqCl/Fgfw2VshoSzP2GSZrea48Taek6RQ3GbiyNq3VpKpkJLASqUXK7K2
3maqonf8WDvKLBRtaKglfZEmdF+22UmgHLEEHXl3TkGu0dzH1ld2wBKy7/O4mu8B
UvxoKJ6IzaXS2IddsacYC0XmilPGSg39S5HynnmdZR07RTL/zeo2TcZ1rx8RLD4E
qHI0hnpBoN+xFG+yJQJjZaYOkYPjS01P15gvZtEkGS9uTHKO6/doNYZ/GCIV2sM1
27OyqEvhn/govPk11N77WgMYdmxOTnax7xRbVh7LfUXd5lCaSzx+/tDSKiNXvorl
L5EGHu2Hfh/YxBXJMTJpkOV6t5DmBDqfwjfYruurIXgq1FTypJuWKnViOrbXWm9g
eglE147dnAetjapmlddNag2ETATyw6ZBVzQVHE322DuJwoQwc2kJTYSBJH463Epc
47X1wJUyP19gW+xi20wgWx+bFBerPaElxsk3ENLCB7t0Dwfq5zhU2P7yed2v0VQN
ollY/vZdoLULku77qG4MHWQ2NhMypVgw44tEKwjPm27a2HDm48kEKq/hrNA7QQZf
JKsO22/yj/5+X1zC0cmlJPmH+bU+3uRO6kirTzYdWUOh8j+oggIbUrc/2kJVmpvf
iy0xlBRdbH27KSf0Xix6FmzHZRvhW89I9KfZXIDq+uo7iWfJH4eoi5VkoQjmlE8V
+u2JEeN9edpJu+GRrlKoh0c79h833V1+AgsiXAx2pcM9lNNgvtPcFV8uSDc0/9fi
7VEybZdiGtm00wYwW2mCDsWOKa+iPANoR69rR2rzDYV+2CNFbM/dCi94/5fCjwBQ
K8fAjLA3W1qxbLaa895mJprifca3hvQuDytV6D4qrL4Dmv1FCTFWQDbTQy41kXsp
l41qj1gLhbcvP00d9UdGM+zaZrTEI4fx0Xcr9o9j6Cyc9OCNtesGRDsQgrvhp0Pq
vyPO0LZtVRQ2d6OgLfl9RQVuULZMJ0HNzF1jEjDPVdbH3uJNmgRJJCGesiYK5154
So3sOnyqEtvG5YENmLc5mdUr830Z041ZSltZhRmVLse7HQTnCzMC79TOLgaJ8HhW
eTdu13AQGizUrLXF8P7KY2Av+6xgPCwDdZU7IZ0CpMEGPjJ6qkEpRI6iQDuEXSVl
Z9yV5wqSwqPJsxcJ9pP/3PGbf2D9Leb+ygSRktYfuoTpdW9yKNJFwdGAPPKN4s4C
5Wk1R/w+0GfoU+uW8YCyHbZlaKYc/ghjlhMJQittYBB/MyyWFglzTZaAEoepSDm4
/XgEKyjr/rVx7yK7xoN96LlNRhdbcgBwP+i2xMpYck8O56HbpnymN6bHW+YRulJh
QYV0leSgOL4gF743CI++/MT+ZubkffwjqpDgoHmqDRYc+xsZoBYPGQKmtGLKZtV8
SoOhFeJuBXgdffR0D/G00BHsN3pzvJLYF0HykczxPUsEWPlkJzGhPRxXA6yWlmOC
WeayfLh2Niu2JhFPm9mX2L5AjEDpbtGwcCEaLTj3EWwbY8hl8hE0KOioLz2zMltV
mJGTTKpWRLws2ClaWJfX18pLYHq5z1ZGd1hUVCJLLS/p+hRsFLzodZw8AC2dXfny
R26iQooVupizrmHH2CATpwbA0CKT04quvjLM+l436ekHHaRbuoQAQNT32Vr36Kjh
RyfzT5iUP0uN3eFQTRj+oDIEn+sXtVg4cxVKHwX22Bzm42vIEVpVahuyodIke3RH
v3fwerzezM29kqLf4pBK/ZLhigv7f3nF9kBhPQG6oAEy8LdG1bxQuzJ99keTKLpN
EDSuoRD8FtzrMhikVUW3Hzki0OA6aKbhbKfTydm+Fe5QkvxtCqEevz+nM68IzFs+
ONNQvOewPwwxO6nEEQ0xZLG186cTexCm7y8fhTFEND1H7xMgRAA2fwTsUK0fqCTi
p/t9k8giUjZLe1kPPtvgGse2fP4eyK8UGvqwCVgWE0NI2H/pIT3dpa4QMSYgXENb
qEplXnLm5u2keQD1bQWwAxD1qRn78yVqT5pIlWhEnSd6c9MA5INcV8mDxk9ppI0F
IsJoJny1rtzzRm+9AAaPRVBDE/IPx+V4cnPsxRmaz3ROavzN3hmQVlzUnpFDSRRa
QgeETPTHdZQvgZwMv/HnHQLnVCo1SLZS7/utC9pNFCInqKrdYJSfoPrIPTl62PDz
awXPwsX5ln0SL661YJXziuL1dzUnpbRgguzdrgDNp/JKZCF3ptN7U+NvGdaHE04n
l14s99VSYKx0HtlYnTbRy1p9ZHEYiCSvjDqYCEGB1n5S2ADniIu+krfkHDGD4A2W
EdkB80cv30nfLog5U/XuzBJNivB+8wzuramLH1yfo35xWHTJFsT3P/25jseTEU3u
1WqeDnfzSW3t1oycrShJQbxgVeFwfHcaWWUGtb+d8ZIC8yr5zcFErorU4svri2T5
v+xPEZ/0rRQ0dfLCwREqULWzjOJy0WaLMfyI2U8oJdGD2PBTi6LUSmKqgBZAnWXS
DgEXdNZY1THkCeHHw7Gg4fAge4Lf7ExTjeq6tjSTLYJeCWdRht2/zfCfKhKw3Liu
LqZ0ONNHfNvTTn2vi/EykhlXcA4VrHP/Jl+hduiZS7G4M0Z5/CdbmIAR/cMAdZy5
nPat25+uLCPc3HvwjHFn0p0movF0P64o+jcT95589aUsaa8S7MFQy/0TMkmBFFnL
o0aD7XvOct9vyf1RvGZxZ1uR2qN0sKUfATAy5D1IuC/QBGDGxCsag7U/AFnmwTlc
uFvw7XrJZl3Cp9UpDtChJwB115Sc31jkSUXQS8WeKH82h1JP58i7LIaduN4PKprR
qG5RntFZBeSjaYA9wmt+URDTQiMxdPRA7+mRef9ncjim/nWCC+sdozlgspRK48YX
JRm8ZawwraeAFxEyB5tyO73Zp80+XGUl4lQZKqhPqS9Ch/HHi0W/5XIi6lJBypLs
xFz8IzcMF5AjHC3TNo2BBD7MqyJ+y3UOM0NUV5yXZ5ldAtPSLgtdZee/s63zwC9n
s1B2a9Fp2tiJfX/grZAcvUTRf1YmJ6wdq2AxtJQARsSiqAQqS4O19+SziRSq2D1T
foskrFq/KeyBOGG2TwoDJJ3yTV18AKohSmWhlhTRMR9EwocC/v2xSOcOJTBMKsVT
+k+GrPl4+t8dbeCCc9Pz0ivUSBxP+ZkeMnrND7XqCnBZumxSduFHTsLdpJmZ8A2b
bMOjQ79IIUHhHQ1ZzUP/K0KWqv+3dCVTB3Aw8kDCGfJihbwstzE3Shnf0HeYSiDD
fA9ukUYnNTmG50UXYKQPJCB3VYHAJ6ZZC2QruqRmnpLM+WrES3wP77YxWYH/BaEd
c3dNOHqZ3AuwOo95bGkeFAuYmx63rOrELLSPS3+PnzXKasyK0uYp93NaIJ2JCoJI
y2LUyhnVnclolpgOpaBqxFjgCInQ4gPQl1mNaTYJ8VV+GCHznDrutKOgxK80ac+t
oRV8WrfXQMZV2tO0PI2UvrAs9NtZmNOKP2bGFySuDtAvmBGVKKEsUqI+t7x5hyqB
urbHAGMGZFAI9eH1+8znlGRqg7kvr2reI1P6c1PO3tsBK2ggFP4KlGd+ihF46BwJ
bGxwdUAEitoZXPPaob5wjKGlvfz/x+M0MhNWLOJasVGsAkL1FmXF0jl1MYZwNGl0
U/ESkMRgyd04PD25+ig40US9HGvNYJHfAHXUiVBqTnXIGdPmX75B5+S7i5VPlyHL
G5HDfLyQr2NvFyFo4FsQhwSMUEtCE9yw1C1PULAaEIBOF00BO4AQu+Xi0KNyzxDy
nGXcNE66vMJJwp7w0Hvc3I6RpvCCmvnuXCx6Yqa1eVaErMBKFgAgQ33aVmv2BLnQ
8CkfDMDxSWXYNl2cK2kUNnJ1yk5vynXXFzHDerrbaecoe2JRLtktpljoTwveHBik
nAOhavPEk2Orz/4nsZ4/hwWtdwp4jOUUKFxIFJ0WvSEEenRfCZ+CG5O5AcFUzBoa
jN4lpURDr150U66LBdWY+fJKJZneKAPgSUB8GVVxIpuSwvbVYMsq9YUDgDtTnuVn
GnM5/z9BYeg3rrC058IF3YrHVAnlDPlZfGe6XU0u79fWjbz5e1HV53z/NIxgz0D4
s5qx06noZe+z+hlEFOP+HdH7fIOf53JF5qHUupGesLImS6OjiZu7QKhrzee47pUx
PosBu9V2emcAnmu7NjnL91SyEARirFhs8YnPrBdc80qN7u9kpmH87r2n+3csSWlr
JbFpfcyl8WTDGRrg5K4lhk8Y3cO5nKhBhbkpBX6SDS+NSPjJpYiveDbtCIdAO4vy
FvXuxBWR7a+mELdPkEoKfzZDEpMGArsuCefrhSKiGHbu1qYqUbHey5YnBRHNVNf/
6SuTuYP+M0Du5SyhkiR0Cy0IXPuQqbw9Zmg5DKFEE4QrZnHLlsfTuPcWQJ+mhNiL
bIRRL4nZf2buPHpYI92+EWuopPtyqM75TfNzF1i1X004KtimDy9JVrq+SXTMU9mz
0Vz+WonhOBzYg5kRV66SkOgEZ2HymBWsa+mJZ2T+CPGzEmeWzJqSMUP0PycKvA9D
dfuEJnzF/hjwojVYPQ8a9hbeyNltA6jz6uD4k0CSFuvQOQhY+LdKBXsda9E6eON9
xEwpdlKeNNZkTVE4YGSNhtiiYaMHfWY2IVJxsIP8OmHy966yT5j1nMvxzVhUcVtH
W2Bs2mdRah1HXdlBOYdOei/AO5nLLhFn4ESdq6AYCToz0sndCBUMKQDy2zH/M2bp
G5WGuqeM7CC0XRyFpsn7ZUbWC/x3J4q45Hb/Opsg5mhJtVkfHzpIRj/YL+sXQnRb
4hRAh4kwrdwuLp9/EmJWCyMGremJ/UDN7ZZPvUf/Sz706tNSfjso0OLvkCXdaVcF
LdFpb07Tkm8Ig7JQ1LtpodkPkooEqx+HEBrlf0ZovqblNcssWNJOWymeABToz0mr
iUB30IwaIjAtRLZsS4XqD96B7Ti9IQA4Q0F0vZhbYHMXxdjvK2s+xN4ntRQPeS6C
/sB5EKdWQl9sbnj+eEyASVYM2pPsF16pRmXQZ6glxz8NlqjfAbKIMw3E/24utv1U
p/Kw+ImHM1nl7nHA/f1f7Qwe9gQRyFNlJktdINo2vaM0G6uVPGcWiKlq08Emv1IN
kqne/LOqq1o7nmd2c/T+ESbDh+nw9qjafVHfQ/VBa9C4L8nxD4WAB1tDf3VX85Y5
SrSc2a+DY0otCjNd5aFsLN5SuQnbxZe3Teb/m0g3/77qlwxjWLjJ5GB5uaE90rEC
OITpEmLRjaqPVuK64g+ssIrVDUE+IMqodPqllVHyyS8VygRc3t5fwGwyDh2HpSEt
cesRnXw2IMt0QxuYAP2uTy0TwmNcUL/dCs0TB0qum7tAzZjIlLLmohovkSF0x7r5
xkDMKe58QzciSRRQ+eFwxRbB+L9kBHe0zAQXl9yN9jj0BSw0q4fgzPyjnA6FtAcj
PjIRF3eQ/cZ2jd4/6Hx6gBsrVY/y6etDOoVryFS2TGa+M/QtwR8XM/muC9hd0mL2
8ILLF8k9SAKpmwbiSSpFFIMiHrZPoV+0nsjJVKokdy1iqCnoJOiiDVXRrJ5C9y89
TSjE0ox5pSGLPWrCNrD/bbAPxXY0kUVmK/TH6sy8qVHuN5qOgYEuB1WnrvYtAKcL
YpZLJTtPUxEeiGE+KZ4oRQbJFd/8ciaEW5sHTkRLEPmnfp7a1M96A9zYTsMdSJKQ
0WpZMEwvd8W14RiAiCJTXBcx6Bc7CuSLLcqDGh+VDTdRe8AABkbQ7Afs22j5HT12
i71SodhByj1PGVMGaGEqo8bwDfjexS2xSA4kxbSfA5hbdEx4CnNbLmzFXT8hfdix
R8yQVQ9WcPjhyVrk/ink1Kq9NKiNOj/T1TuAnsbmvL4Y6YtjXRo5dXfisXLXOxO6
nMKM8rYGzIDXr8/p3beeSMPdblqkpihs1dke09b5Ha8F6OHGo2HO8DunMgLyy+jE
B1QINJ+p4FS70uTC7fhifG/c7nepnEeubIlfXsaEAbdQq6zVedLlahXM0UVifbEe
stgR5qfsEx6MYRgv2XXpbqHQof/jtYsxDYoufDa3+AN++ixrmYM4uqAc2ojIpXCz
k1wNYN5IwImI8UdYKO69f6pDk9sYeK7QsGl8rWuqbc3kVsCCpIIVpnDr23Fq2/OG
4H3KQWNdS8YK8WBrcCx5EouU4SfeyXaLrEF6vZGVzql7bTNybNOtv1b/ZASbJxRC
I3YYNnz/e9y9CSnQ/7vaP+pHtmonvgXyJQ79rGlKsxJFxaZGvww/4X7pTbZ8//in
TWgTH1ZWDy9zeKfH/ZG0s5beq0zF83t897d9b3lgWrUT+xrJVDtxHKrFqH/noqpa
m6DX6DpU3L5fyxL/37zTelXwEd20EAjMZhpqY/pBw7T4wH5bsyq4+VORH8CNTMcF
hKq0rUONxxDrLdzQwq/RVWffX2ZZ8/sfwBVkB412fQLs9vrIRISOhbrbUDx5PNFt
An1dX3Jj8n0uEG3KtcvM/Vvhc+lmgQfnlcYdRls2oLCEgowJTfgdYKYIpzKP6WPM
C8QgzpRRKAHfFgPf9r61Bdgjx13Z71ElLT8R8ikN59AFGSsWTQQvW5Zg27RBnXFB
BGMNvFiSd/fEUmK7ZjTHg/NVACdIszB1ffCwxr841TOJHBqSM24UIiX4z2jPTFYK
u3WQb1+DeosjXsdt3xg2PDxjUvXvUu8DIo5MTDeLwE3wqiBImjxvPvo/kDphbdFg
1oGgPSnMWTST4FhcIIF7SRPlPfKZvfrnFaWOWzEx+H2RYw3PYgQq4fHBF721mi/1
Ze/vF1Rhy/74QnsVBB+NgKu06IB8iFvepdrHaB4jvo0GMuwAJi+DNQnyydrTE7vd
844ybxdDvMOCYsxjJv6yO4CDwzT1LH68eNc1WFJmCdBhsVBu9bQza8hQ1+9RQ4Ot
q2rLFC0KdIBetkR0bjzS5w/iYaCKVo4STGvBjJqtlCK1GLJBh5KUCcx3dHxyrNy0
SVRSizNIWOeXyYCev9zFt+q/h3wL9pcrKgkjYZzXlTXu1mBCIviOzO3x3GLjw0ok
KKcPxVRAXCGwYLPTTHIytX2Hy3kzY2lSom+dHe13t5KlRUDcEwCeVJkaIATLgRC2
CgJgJvU9Z3WTfJ5QC6oCu3viAI4+W9uAVYYgEbQ/NMSVEjVS5eJI71l6ndW5Mshk
x/YG56rVpBT3H5FjpXizK8m9fhcVqafP+nzNCB6VaxV+WbMY5+luW6qjKRTvC4vb
RfsKd1qgnfgbIplUFzxoRfq2KvD+MtY2hae4ePifhRAKfqpw811U8nHl/36QD6RS
90oQoZ+totce0UpJ5z0N9yN5/UlC1M3JFxo5+JYcmCzbs6xFXS5O1IfQhjU+kyoI
RQTQ3nm56XC8lxUmv5pc+oHlfyffs9nAxBjzuXpf56IFcdSXTR6GnA5O8yuGYtJr
cpX8H62ZXnQR/Q7VFbUwVsze1xOPujDazpsvS3a1IM8vpiK98A2ezEZcCOVuQn9e
bUfZN+HOu6A3g0MV2Z5wsZiY31Rq3unzVSNEhxxg81FhmWEiOB0eJ1wfQoDcpZcx
KGB36va6SX+KFa9/57rQrSYpEZrWU4aT4mwAy3wP3JK+h+zcAZjGb0WOEUOdKEKs
UXF7YsB2Iwr1R7UgtDoEg00E10pVq81d6DK6YDi2A+0EWNrPnDVs7vhgb6jRWkPb
mL3kp6aF4Z8s++ViyHyhbKqSZZPHjEWaALUMYm8aoUdDKKlgQeS499Fvau2JGI3F
DHOYlzIJcMou0QwEdRfRovwcWN/X94QxpWkq7gtAJMf5+gyk83/uj8g5i3D4grHZ
+dJWfl2ZRYRtWjLwBKaL4PleW0hO3jxdyUkq7qyK0Q0CSRftpg4XoqBo/IK2h52y
k5EqaAsrzSNQdeDJ575tr+XYvyqF36y9tR29eNn+FsheX/NCTj7fWiODvlHjl47i
l7RzV6tYCFEJ3+8E8tfVfANZME7pi8NSnZhHdlzmE5y5mXQmRClpheJn9Ut26iDO
tLOOcLUObKSyZI4DZBqYdoAJ8JT6hFEn+0HuVqWTCm4jbaXnY1PGReEBxAKwZ8oX
qccPHepnggrG0+z9BZ4wvX+Rte+TXrYemNuN8l0e8euzADG1UZjemvzvDXCW4gou
q9c/Ckjgvl4Sg+V/m+DM810Q8kazkduVbac/u8+RZ1N01jadD+yOqwF6dV9I1H/w
+XSmmhnkU+yFzUa0j5dK042sC2LSZ/hLDGoQyQraEFl2b345hJTcvn9FBfnWYdMF
pRYBNyXQHvnmsxk0NOeFJ3ul0ZQNSicg5Di9sSu5lDugHmGTvpOFuDlGCI/JNRpv
xEWX6EyffIOIZLNLsiwjdmDc1FOGtRHm+cQFQQiiHxHt3QvhGtc+7nIQr0zmMXyh
XDwqKrxrxkGxObDyeK7uVNzNpu/xYu4eZhao9MP4Jjdr6efPOpQcv9z+ZjwSHmth
h/iC8V2bpQVuU3Tq83EMDfhBmGt+utGjZebBhFxRm3PJR13/9QIgK+vyviogeX+/
mHsW/l4TVxUH3rWUvp+tVBvkoz63+aKibXI64DkZjRCuZSl86UlDUgr+vVOrcTmk
UVG+whDZ8Gn7WToYv2h2EAksVtmDgo/VRM9WINuITvLrmwqRzPOhKj6oUFdGhl/I
055z/ncDeNrt1HiA3Dk2ud0XYedjfkwakxCU7gwVRl5S5BSXFfyCKQ9Xi2yW8pMo
N0YGLlwmEU5QOMlS8zSaPUpqaP/OsoO3K7Jrv88rqyCR81KKwrgdnc35/1P7XdvO
3PhPFfTGWKT6E8KbuW1meqYVviH480iEkaSqGTmb8Jt8qs05VaoSC7lUA1+Xp5bL
IRONE3rjoc7aBk27njVy+NWczNPUvTs7te0eQjqMNWOZOWrZOkonxwZF82PnbHBs
EnPVm4ho4nUL6Ju+WZ18oRdsriDPtN2SNw2AUnrJaMwghUEULoCE9oFytMcJ0lQ9
b92uwuYv6CK+J/K7uVLoucntFNEtkfc4q2TmyiLlmq1kZPLqQmOEv6ldfiyMm4ds
YZHXwWIYhQtWhNtpxfSlk+yCGtJqmbOOpzr99sqoQhTRy1gwNX4CXxuxn+ngE8Lr
ta2/JFyrGK0bB1rzls9ihDRclGNUp/XWTCGutFFkUo7W+j0t1iLr5S12MDoGBgpS
58maq42meE1OWbTxFm033Y4/KU513nViJaB81aW5Z7MorS9yNR+sMt0QLc8JIQhr
kkxtDvaRrO3ywKjwmA/r/kHr7tZgstV8DaTZuG7fnG6igI7WknfvYuJBz4pUhv8C
n2+bDcowWTOCwtUnZmGdqTpYxdAljTMZJc3+pQBy+xGtMI40gDllbWOPot3W+amO
rxr89qGrpyDuwkUIVfZ0Qp2eY2DKl2934+bfHZ5KNO5DUsJZTsBuoIYCOsERVHFR
I7aAP7orBR5LvYblOEM9e1r4wH4IRLyZiYPwuDJC628O+BWREOKRxZ/vJd2FUdCc
QCwwOj0juwXA9n1Ivx+IaWVfOPuWK5C5vZBQQZidXyN3bSVgJmEG3pBHgWn8kymv
K/rejGqnDP9w2pq/K1giAR4zbQihHkEBOR6qs//YhQYDs2rMhjsod8AsjQ1RpDEg
SzKBMENP7bfz18QQPeb4hQDxtibJq3Vb9qOgSjlBOsAw33iEjdxbRpgNKkdZIRUs
ygV3AuB8erXFcz2QsZwo8xmtp0zhcXGKdaYtVsMQi3X0kox4fQNgIpvYC45OAXdR
zd2t9Qs+BzbWwkKYWD7pQWzHqfq0rf4n5m59btn6NS6fNk+7s/hXu56s+kMDeeY/
vNB+POlBm6JcZYArJYuLjpPTw3jA/A+v3elWQWMF6Lsf3SWWLxT2jz4pRm7+o1CJ
/oUAXkQygHdZ6kOcM2/7xJOSwNJGoCWu0RD2ssc+/OS0VHS3FBITxYvvLDjeZcEm
CJLyDLSYVCgZYdXSybPjRJTQi0VIZ3vbg0s/Ev4m1QYYnwUG39LyZRleQd7kNWvC
Ml6Fn+YFJ+pmo6KMYfkINzeQ0Ni7GjmgtsFsLTXXfrzqX7DJJECNewTDJci04wCQ
Dpw0oPOTm9ZX9JEaE+e9wxxV+C+4oivbthhp7LJuMgyulwSJF3MpLfcSU8fhSdC/
F54V6KD89/iuri92QS+OlIqKwJUqUP7c87MXmYmdf6/K4MqFNF6aPxInrftBSlfT
mTJI2ttbZQ3eHZ0W+TNOtXcF4mlEzNaioVdbASFYqHnInzWNyEnTCN5tiwrZOkay
24SczLZglgXC43IEwHLoYvT3E9Ea943P3sJ5d+e06TyNc135xLXMaEk4DT72Y9WJ
OIXWwwso5rKfV1DRV8fjAZX9eS6KqQyoVBgUkovjZ45dqX2N3Stsmjy+zqwLP0uD
a+j/kYx9RSkIPUYlOaQoQjh21hqFGB2gzUflKTQzM1nNzQrq17GyxLdNLg+y6D0w
coH7GjO2jI2rjZvc6T07CZmUmCzObmv7wNj/W6LuVlnVIO0UWtOphK1U7qenu9Zu
VcSU8EovoFSn+omXQMPhTLlhX4Zk2yw4wym6bZ+HUns4P4oNDB5ZlD9EpTuy1gu8
VJUGKU4TAUz7a8E7o9rNQEeEmUMmxowzNwQhqt6NPxbNHu2k1MFASaW4jOtqq9qy
TOPsCYKRddFBZLnFd+02BRaKlZnz9YhAJHNo8vGASBNmgahDOkg7Z+1cyxPX250T
PPrDa6EpaDUeWJXuaHVHFlsmZtV75nyDu+rPD2/kHWM9/sFoHzadDVOpVlx1yEHM
vLAaCrK+B/AtyS2yXYFwKe0Ao3FlNWyMQcUgqRWWdwMnOfnVwD1c4jwuk0R8JexD
j/e+MqlqcAHJuVNvF7OyWPWlsJb0wfTDxnNGr9qa0g1MZn7jTeMqUTsneVCUyIAc
XIz4GDHbnh5LByHWKDEnwgN/Q/Ly/bdGFHH05MZJmKHZ5hJbFLN6FWm0jy1dfzwW
Lq1j6Xc0aA1U6v+qQ6/mA1XGAoqhHWxBG2TogzYC5zttgu9+6Q6pFLPSNpSO8ddq
03xmsIrLaqbSgibPBB0CiQQHBy+mLK9VdWcsIp0eZysDh6sSUEbIIpReoiGLNqrR
9hAv/yXCHwZZOk7KIjr/FV9dSw2Z+cHY0Lgo9fvqVq0NHHkrm/DYm3bSCRD2uWza
Z+zr6CcCBYoogNGOT0BLmay1305Fmo3FFn8AzKL2ndDnhq4oQZxihrZ05TeTdOlk
fB+VviryBpFSjz61Rt9cxGZ3wHJ43731nn8Xh4OPzn/2JGPML5FSP419Q5Ysg+w0
EZKHtcjWwlSjQ1GsD8o0d9o+63VBAH4erH3aefvWT6ZwVHjC4DzHfaulHHCYv+Ib
x/M9OQgiVE056zGMlmJguxj3TQLOKdCNR5VyXpQOe2RXmID3WWdpITVPVHvxiHas
H+lNyx6nzF/hf/k0ltO4y3KX8cqI8A3/B+eoiqEWCYn/g2XQ4butQFi/wmPwanjk
TjwX7MJl+V9hTy6smR3rZknoWWeVdZJf0xWeAu35vi5Wqahahk4Zb4TbVZvQ/7h1
MajF4ETRn4y9tCVxRTwfP5/q9yXWazYLPDZ/Z99yTJ0v/rkuZc+Fv3vFl2OwXpMc
NaE4UEKHvFke13Tx/PN46bcEkCLGCoRozH39bWWgYmNxbOsod42OPGxSFJH+I0eY
+WLLBFuJbxlhjG9G29t8HhBGqKH51XnpM1Kn4w3tKnbNyK/GensDhL+BsJ8UWZWZ
4Y9BieBHQMk99gMKUI0EHBrU8i/ZahYhUJ+7PU19MQxXzrFJLPEWDPKRl8dTEvzs
CM+XUNDKZb5I3Aio2KXh7BI8ZkIcJzOUw3s/yoEvXrrb6Bk7BUlN2uTLYQa3dhqb
as4OpUDXXZaSpT/GTMwEmZD3D5hZ0lJ82dz7wk76maPDCja1+FFxpVWKYxNF/H45
YF6ubRkxXEaiXpILQZEkvWUZ3BgbkVQeE/gfd2Jc0nUOwc5M+M/MYQp6o9H7BjBP
LaaKdXFUx7VRYYrOlHqp+lDB+c33k7D6tCC6l+6ehjoNv35iQnkLZ663YC7xxi64
VpJUR1e35WQd1fBW8FXyiCXT/IsDl4NtWWMxpUNI+mZOwnbE7bymqsn3kfTjqxuI
qbWDHC1oE11pTmQjr0EMFBlVvF/BArt3nfVCSNC7IUgSjJmdVGsmAM2uh84bBqs/
UIok2/3PrpoXZEg10spvto/PXRMwr6ea6V1JtwPxASOGLUn41CUNrAWtLWlv88Lo
MnW2ykFhVbE3qy8V6cn09yWei3XBhzOaUuNFA8EW7xIM4RJo6Y+cHZOHdW7OXtN1
MNnJBihN0TfoAKuyDvQBoYED/MUgv28S3iK2YtsGtwUEOR0JBFJb406Oo5TSuxwq
9RJukUfwNj674Da4khAbMxeAt7DsyyS7MKch1asKgd1ALw4MY+Puwc5Soz6xSViL
+qdR4eIdWWPyegAMA9QWN2kWC0Uqr1OUr8SPO5FhAnOH6gyJVCInC7SqCDC2Ugjv
FN35y3KF8xVBn20XidtUJ8Y7BfzpAVDTmYHzOAW1uiXTS34TvFTjiEe0ClKPDP64
ByQCnSCV5VqSCv51PpJGGbnaw2IVXlzYtXslwgNPfIpRAx6z9dPEImEwOPa9tMDK
ld/2atRb4bdfDit5k1w8kW23B6Wl5eRsPaYCxk63ceyHQ1PU8s4p7QAv+07pij2S
7sGDkEuKuugfug7HHddUi6IHFQI6E5moXPK1tTq9KeaekIn7D1ooBln4HopmAnHR
1zQQpTIu/zUB5cKZiRm9oONBZNnTtObHlW9qA9FQVvNIcC6srfiHcQ2BECieZE1z
tgaLfRaZFRSh3TwKEUWTWxy4M6WnQJint4epWtKa2Ryf2OpeF4NYua9sJA4ZJWrC
ZnhRH+S+Uz+lIlwKGL+wvdPdR4mbGQW4uC/qgYWCCvt9z1Dz52fxEHOzSigNhARD
nI8GIP123iWSw/K0y9Aad1AaYgyAVH/UX8+s7LLKgGyeHPSCZSb0+rF2r88dh4bc
Dn8uUWMQO6W/wFmvjJutm8RvOZ+i5WnSpJyIRyDCen4eUxmp8ru/gjvoWJLJCLsl
+gxejhQJkjJwmHTCZw1QZreS+vCc22gn/Nw5c4Mfnhj8jJl06kY49O9UguGvAMwn
Muof1uftHVNbkn1HSP8u58f+WaJ+daQPWTAeQJ5vBR3zVOC30mSu+u4yASCsDWtg
7JMORo3kosVg6u4iPBFp70hROHfMOLgKe92JPZNez6uSqedQIiHNwYLCcDfmlmds
cTvdKg1DLrFSftThwyXG/P6NfzsKAClCeow6tQh3BbZiefRd/qvtZsHBJXda4nJv
D9zAugTh/sWfRQbV8ZaKgZM8QcEKl4xcxroAoec+9X/PrYhtM1UWLQfE1b9OvqrX
UVBLvKDAb5OGUVXN3KhnTBl/lLSn7ppKliu/OTwaXPj3L8+8y5flf5i8V/Xsvg2n
RBCPBUumtGw7HHv2C1o40M/tKqTuU6m9RJ2IvoYLD/CLbDVVKUUEufk55tpPjLHn
YsYf/r75Y0ITPxZLztsGM6XRgghqp3GBbN3WEq0+9i2KOCXtqgC8MS9ZaCUsSUh1
JCyj5mM8zNWssnx4TlP/IFYLZ6EUeYla3BsPA/TfxhXA7jRQv5iz8lky7E7p/qzq
QF6oNZO62UEiEgMyfxNkU+o2aBrD2MLbwdwgmrgVqtPyAnbGvnjP9gCYT4DPS15S
FPQlZDJ1ORlmvfsD71KvS6yrlLpVmUl1Agv2swr7gs9v4YcccGtn3DoEYwNTjr3/
em6tIYql/8nOY438o+2ZR2PlbJ8O7ty8eYXU270Ui+LHM0u+7AvmiZ8xLM37V/TL
PN3Jsw9R8LWgUlzISKKAPxHBPWb9VRTHvY1NVtxPQEl9z8JSi/ich4U4SnaDXtej
B+uUk+ZowQwvjRdrU9HP/qJcML2feUWxJmHWeOETaNd+uDByebn1LLEhFsCeOR9h
exaNfJ5i8TmdYw45sWsj6OnqhChoLnf20VNJslCq1GbL4h2zAUh1CaHKTXlTdrXd
UBOV0ntS8uKHYGAHK4RcHgIQsldrqiWwLZ9RMtpDxoatUDhImwXN8kHUus85FI5J
fcXO/VQzALSID4ZFoDAJ5ufmpn3nsiK9XsqzC0OZxjiW04YrXsGy8w3OoWukMobC
lZ6OOGJDSkBFFXhDAjcLRgGLjawXwERLDhn4dbcpHoObj/BgNLoLBO9dsLhfqv49
0urmyzA8c/PUzzgJU/SBHV/xMW8HOEMTMzzpuBDK2pgyt9Gbd8o/QOUD7dt9YppD
uFGk2JF5vckRRVJFfv3FSyGTsAosxe32Q0L/uS3NlFCAFCLvq0qUeGTliTKE2pXy
HBpcx8RpEFhAf9CBGLyHL8LT1fkW4MlJnlhNl0CJd9c4Jnzg9xdg/ZcUNpfrh7q0
95EYYH+c4AJgO01FTzCYPOpUzwAbAhekt4dzjzxuzeI5hGJG6INvWhIjlK0E00L5
6ItGsnSUr8pGj5g3HWjI9U6rrEm/nbtixjitISX15bJAZsJVT/AnDkdbI/UWxYsQ
svOW+yzUaYAgVrNWvhPqJXePMwy3bdlGEh6amTLQX36JUTOSuYVteP2fn3HlezFa
PaNXF+EGAE54HWsMWd+qCkCp2yJwdy9J7OjRNBc5CuBqUWagHElqZbTGz2JUcCKr
G7gA5r8B4Y68UWESevNghagqMRjlbiPbNe2E+51gJEoHfm0WG9KMCeyQcsG6TwE+
glyyBeQ8vfj5IfANCMMf6MHnmkOsZkgYjtofV5QnHM2+ozj9c+9WF7JDpu7ZiQnV
4TiEXmIDqEqkcU4wGKYYlu6+HbPnBFAX3AdONMv7yW1Ke4mX2FmarW4G37LuMAIS
6b60LjKA2fB+PQzZT7oVDZB/nZaeYeSiSimw3JChK8LQZT+X8747TyydrdarQZFx
tvERb7SyXUXk0BLyBnhsY3hGlecK+VED/FalabuBmrcY7rAL0wW68hsicRv9Dztt
PWFYy8/dnoqzzyiwB4WRMhBBcGTa1brAydrnqNebOB7cSLKdH9LEwc6qEFEbcgtx
5gdVY0nfJFXQhDt9IsFtCM0tNoypaiVVMk2HSvJZPawumYo66kzD620n2p5Xqbev
VOhXEkUl3+VNixqv3nFFRfZVAvl/TSncuQcFRYezyfuUWy2f6qTLJjfxKFXb1Bn7
nGbkuANKK73lZEYY5yHD8DQn5MawN4Y696yjupg9/dv1m7GiNVRS0pj7kigqoAi7
C1acT1jHz1ZFqWjl99hl0LD2/O5lEERBxngcpHIkcIR9f8+Q4c2gBwS5VoGovxoc
Ilnl/jXkCMZqpgtcbj3EEHYVN/OVwZgFqfo4KrFM3s0atgitqAa39gG7xHKbgCof
GU1u8m275O6w9erwzrpHU8w4N2ENNoLSafLE/fWNnoa1THVmd6H4pyagDrsMG/3i
yFDqXxAI/bmRU7LPaW5zO+Yv5e5krRlWfbK/hqbNQaqXKEQr6iL8GGtyK7ur4hg4
WshrMbS3j+ULiBkyanfUEKcbDjNG1UQXxyNreJzEn0KVzjybpblF7uvornq7i5HR
hORtQX18zKHJms5kIqKaAb1Salr8BOXtVbDNnjyMdRO94V9PjTxwknF3C8HuG/Ou
lmn88bKkWnNLPqCTV9fdRl0k7MV9Hg1yLJvKNouwhB7uZwvLchBibqHeXuqiEYwN
1s+AwuIYkRDxc1fFXUw5u54je6wAiVYO5vEqjKbeJWbqfUULiNe/qsS9ym0PYm8x
kvM1jIoMc6gFC0UYX7fwAAYHa0/4MD0hnOcyjiVax1fveE7Q16k8tKNGBwydtcnN
Giiy7Ty5SRw2jJoI0H8SFecRdPuuK8JSKJhWscjRB3cVT1CK+kKyldQfMTy0AiDX
ZsyMH9UERkPjs0fNk+Ws057XJPisRMxCFDKpOYyG/bOhuea6y9x7gfgd8WVY9p9H
fwN9Xth0vSyNukrPtPHUtAA/YwWwowmvugIbABSetQiHjKAL+cfa6bgZCOxF/o7e
Y8FJh1taAZeYt7fdqRvxOh0Yvqd4KzoQOt19EHrk8Hzi2qypDtJCfvyczTqUKpGJ
Zik9Zv7Ehzdx8CFdDnCWTenY3GfTh3tJasciqUzJAFF7/8rhmxo+cTnnkH6RsP2h
R8z8WQqaWRzKXYWcLEKq7yKjEkm235KfCvuJ7tRIvzQ4Be+xpBC0EBXdHYlw9fSN
64067yI5wlfLRGRdEwM8P/ItAWG4ZcakofTe64kejIjiQeG4stqMD1jrZ5BzbI8P
yUTqqaw7hUelbOkBGbdMYAV6BrZsSUFXJZ9FipxDxIacs+JJ2C+47MUYznaGn7JY
WBiKvwyRSduqaKbTONhZbeWgNsUi2kHW+JwW/SvOyN+Y7JONZNsrJ1Ani+fQEB1C
z7k33+8nKV4/xVMCF+NgmuHpzWSFCX/I/MsSEQHLKkHMUQ8hdbf8FiulKl9QBvai
Wo8xJOSNm+ELQ17AtM7V9y7I1STRqD0e38LJU2FXjsNaZbT24Fg7Y/2jfMPNPDNJ
NvoDv5eCD6l0SX1+Fo/eT403WNKDRutWOa9L93AMHaxlPxjlfThy0Y3K0FjZkA6B
QteihJ1Dua79PZIDDuwe/191GWwCi6oTo1OIBOcaqyiK1j4js/R71O1Di2smK4+o
Gh5MDa9dy4lQIc3tpft8UQ81SnMtA1mAhZC54pwaSP/7TPKx522eHhY689Pgxt+D
dESj/Dr+MhmL2oYLxo1kDDWDv4FnbPOSSp6MvABDodoSm50oBEsB/5ZvEwIv6S14
8s7YzGYSlMhR8p9fD07VzGXgVXjok45IuIBDGhZW1gAKCeNriAxD0+o61Ycz86YV
UOeGfeVgdixkGECh9TIki9/eIp9hQ2gEQ3XLM1YBo+D4smGLKLItDVvgBqLSH0Aa
RyEnpmRy88UH2yL8EsKyufadW5OSymfqXKKPwixuF7R7XJflnigJ1SOnHzfUJYjD
xBbSUKby9M8Lpyf5sUf2VGZGi+m8H929xcsc1hQCUYL2MECbwKvrJyDQgvWBYEaG
EQ15Odmx7GTtM+B/b2/+pMYgMd+seoeB04pfRE2dAa5A/kemIvSqhdV773RomhEp
NDDZDpPEb64rI3Io/FAAke+14kVFFrVazp/emMbGbKZ4RO2UTWWfDHMqBz5C+56Q
MtiYIcze5O/hDB1iA80UgLEDTdJPJES4mZFJvjN18GhCh3kuWt2SCKT87Kg7gCWv
T3Gi+phV3XR1uSebIFTmhzztgq4Tai8grid2P5Jr3QzytKVrLUgypsXWT8QDw+6L
oKfhuiVF2dhKGEq+7K42xkwNlfMXtZax/xDOADDXuQS0EPfHZ+C0NcIQMQn+PHgg
LTo1qnW6UfM7+VhhFXJuTYlDytZjdCKzDJepeH2qE4BHUv4yES0QmHAecXWCYFHm
vdqzbISvPaC/4sZIadcRbNB3D8njfntvhkVJHf7kvggql0UhV+J1z3Sye5dogcNO
UlnGQzmE5YvaRODU2bwkopZj49iDEyFJ93XRgGZcJIJ6fJWMFxYz1iHSxc1LPaWg
StTEESL6LlkCgbi9yde3EkpH+NdDKx74FdU1n3LpY4sMhrjxiV+cp4SLFTGJiBv2
ezD6POfHkDzg9JsKq/UU1ZwNn+SwZrrk63LZs791N9wojM56PA6d7QFdguuVcMDc
CjP1sR3J94SJN72tfFhbHm/eDi9pkbsbhryYyil1qwdXfFNOPEeKoZ2dPFgpFREA
WLAq81ER/zG0UIqgH8bkXX7+fnh8DpWCuYWKRHEdJiCIpAy9QsBo4G2lV9UvDlb5
dZU033EfgPgpbyDLCImWzwwHDFU4Mm3pH3bzV6qV4vvyJtPA5clpbfr5oaK+IRUm
coDTsXqpS8/odXLoaapEvaB5JAs/O2ybLZecz7ybVZknwKW9ZxNhHgkZPBHwOzEI
Gt3N8IuCrMUH1HPrsdLoWx2xGAb51POnMomNRkno0uAe8p40/ppIMiD/SOXSc52N
xhfnkr1mztF6CpoW4oI3JFejONx528cI7SqTN3MRKAWURaBqXq9vsTHkcE3CnwNx
i7ZsOIsXhfAN/efyWE3Nlegf5KugU5WNq5cgbqNctMwsZ3I88NSTG410aYYbaPgz
GJ3674nbiNB8D4Qx0rI4NJFDayUbX+gXQ395G4vnqgS0VrFVNR6sm1+8Cegljh6q
79jOA3XTE/DjdZ4NxqR75Xu3xjDXZtN++oMU/WExLh4UZZbvjA63OofkdcOrTnv6
RKnllnDWgNXu4iHoh20amrwGOdzxWYKmMXQaNOEI6cVB6GMGtfVx+LnxsgUM8oN4
Ak4ZKPDTlIghjaTgCxT2ClNa2FcInjF/jR/KK1csM9npwtyTUqABmfvwj0z9g727
75dFHHfMf1o5epzzjaXj8+71VOubuAxdYzwgRbEy3C4xMJCvwc5XdtX1/pSXMYC6
5HtuhQbN9sjXvj6s2EmdKtrHZM7PGq602+muLy40Z7bB7TLey/KjtcTo/2eeTSyt
l4nezPUdBzibUrj+H9flroBvqsFEicUvY4PxLF3THlx9o/LvvmZTAySX4OEJ6GuE
a9FLoYiHKcROB7HugbDaFK1O+OxUR41DNOPyaASeITZ+wZ+JrbjPHhr8B8OlNhEC
PjYt2+j6acBwD5VQOtsnxv3J4sosxxIwflHn6AkQxd4Ux/B6Vi8Z07DyCmkffjWj
wX5tX23IUiTcT3Vxv01ZUDdwx0h2RWMfWBUoOedccT9HNl5DeOLI50tRP3lmu0zu
WWTCFI2t+9b9kkBlMVzy4IbM10LIX5P5EA5La/cuOw4I91S3nGC12Y3AkIHZMlGq
TuCjWLx3TOU9K66dXOgpCAmndqw01mECG3Qiq77gz2YKwpQyUh7qFCkg7hLDDfx3
R3uxIE8+V+lx1dBgULriZWUj6v0hNuipl9AOZ/qmZyySFycjuBRPkxrQDKXM/iI6
blF+GtNHBx1WERXwyh3qiyAELyoeYGuDCqSzno6E9zhIFyumGmLEggf/ve2aEje/
w5ObioGsoVttKSho7Ihd5ZWzhGnJnYxqOe9M/74KNeWitV5KU0KiXYHOEUsp2QJ5
nuNzqFiPlB3TIPHo+K/dY30Pp4J2pUtntOC7Dm9ZLCwTvRXfNmQe90J7z9rP1/Lp
qgHyJpct815E5/3gWpxqQBBovHRaXhJVJ0QGwFV0Q0NpeT0brseqZE7wvXw2lvvc
yxaAAA16317Ym5kjMQDg04VHHbEqE/yPzjWpoWsYyQTrU+IaWWpLOhHq/yhgRrP8
kWiZynr8DvggvDFoOfFE/FrLSft1jwLcYtHONHnmLcyjZgruYY8U7Aj2hutn1MYb
+PSaH255zk1PfimfGlBxOVxt8gr39Y4gfHe2B3uxeScuqSLHMswl4CEFPdQ/93C9
6FVJVBuTJ+aYU7mYpL+Ygwkc2urCCetW1GEjCmznQTiHeN4bdCOrBEv/OK7gFT6I
X/zxFIXpBZNu1SdPi3CeE/C/fwPpWST0qZnqAJF9+u4Cf6cuHo9L/XhmOMIkpK99
+g8e9u5Xtw5ZbIq5krLjnzfjp80snQRnGGTP5zR8UwMRZA78f8KxtUSlKs6X1Mzx
A+3ZX5iZWoocKnNwz8qzWS8AOqXoUxXIsWW1+eFtnhOvp4NTk1YdkEykAlVj+N2M
LvazBV7nVMrX+mydOf77dS2CoFgVBazGXxz6W7fd5X14PgukicKJkMZFOaOaIrvM
0m5AYNBjaU/hhEPJxnMMc+U2fU2mAstimr/qHH5Esh7oI0u+8shawBJRZDiy8D2R
XnWEBdbKhyLh4LiWpaJkUkpvpldtvqBNqziPr3xK0cVg6ta2+KC/JWNB5TNEv0s2
bnf/CYISLmmNXc4o7iytaE2VmXnXxQgzFRBF8VVtfJxK2FV6je7PLZDv5HjYpzOT
XKimQ49mvN0YPcz0MlBE68GhJlvjiC4FA4EiCIQ15o5XsLVYo8VyLh2e91af+WGD
00rSTuwwsEFe7thjJwAtMeSrqYQVRczHYfa/qAU86RfsFxChAqUHV3nBpfLZWM29
OsNlGCX78XgNWMabLGWnJng3FhA+p0IvDlQRRfDbRh/dCUDOuh7fYuAcA/kIiCWN
YuactIAypLq2NbsSBmj38nEGiVkXfML71MiwEEkgJ6VIOe1cLS8ov64cAV3LP5if
/1EROjbPLXZVKTX34BE3Bo2i8/SCkm+rPCWfsGCNaEIDEmf7HljdZEgobnfx4JX7
sncYu+zz5a1VOBkmpULqR0UCP7nSY3cM/9hkCeOjbuly6ClVOc+tnCgpN/QPr5g9
8QbygDmrY5SpIM5BrotEkyfy7svIEaUKXsefmKDronFaaiCYLql6Oe9XJw4YuqBV
hxDjgUUeJiQjvJI7pU5OcAqyrEDpWBPKajwAm2tOxlNaxVZaIj6tgap2/RGPv2Gg
OVoQCW0PTdwvKNLHxajrNpqaGVHvXQOhCRX1u3Ns0HocM4fK2x+S6GFQsdjmVBkW
w1ysYQIotKkp8gTn856sZRCLzHML8VV0BNTFH9BgPTtbJur+XHcw3l49UMEuQroA
x0MnHCFJQ50TCZWhL21y7xYySqgEaiKiOKxMO9s1Jrdy38fCFSvjmQO2lgqf7pBe
7JcDWWNV7yY7v9n0yq4ERNh5oikOb53z8nPSpN8Cz9SktpmQQ8xyMTVN4rQgRX7k
0I7ye0fJT/MyvHzp5MmfFbH6ivflV+rNWEMu9U7fX34pLiOr0ou0IVjdRfGZ55p5
bp+XRaPIm03/+zjXVEQOOCZ7ezem2laAp+g+j8zl0ytCD8nQ9caieupqtouGwRee
NRhcNgJAPBG856x17GoiT7MiVMMnLAArGi6UcMhc8Cr8WmTCE3vltIzSlopKarVB
nnuIl3A4bb7JT1PSa0hgX1qr2PnNfrKPbcou5itfo7/BXclVPMbKA+gJRmaQ3b3q
4vlrTj4f76gw2NOrOemdYbJD8A9FryGnQ7MYdHnkmqlpec1GccXtI/FjSrhhcPiY
lcsFDYAu3NemjWNwVwTH8lxtQdgFRDii1Fu42nMAR8j394JHVoLixnqQ0mLcYjOK
+/fwMQxVGAGLJfMaGVWtKy9lH350lqAOjoVcaxGfWoyRx/5xjxQIwRIwaAESFN4l
QegnUqoifhSJrq+gPvOdmz/sEkULxN/s/I0/qFuy+dFM4ujA7oNnKZUwHmGGxns6
h7Yq5B1bJXaME+rUJW7CDNjqK43h/b1eQox7ZqvRX+br+C5lUaBPMQ2GWVEYV4pW
YJJDFikGdfLYK1AfNGytPx8KFAp2LZ1oK2nCf0vbSYlct7vZgNa5fmfNJEEq/iM2
fj3ypOYUPO7UeHsNcWM8ossInodJto2Qt80c9JL1BfDlPUXZ5ojgat4XDTtsstP+
ib0YuATDT4rUgXe4XVdrHhPLcRwDHtGnZemx0dDcLAPAS34aMiLGLU8JwMj7JK6Q
7G9X43bQksTyvfcVTEgGIfZg72bzCV5sDa9m3+Qe2R7Ofi6UeMRMNraA+eXa5jB4
QC9t4M/ETNdIs2rzFmWXKpL7vzBoR44R1hbtu+d55iAzpF+ErFkMjPOTeIFAWZOe
Bgmgte6yIW25Tt/Eps6xRWmQcr6FjzLL36cIIglBS+bf4ave06K70chHFGWWFmG4
g3wobAnzsxlGFt8Cj7W4+Ygka8NdBoNu+67MhP1N7dnAw8Rc7uffxJtNHQMOQuPW
Gd4WjnZWw4jIUGEYAWtFSBAl0KGuB7ERqUNPb30/k+PXKl1U19fvAXZx/kT8jrZy
OS+dM+AMLmcwaQr5l7CF6D/rQShotkkdyEYcR4TQ3iw2dCy5uB3S3MJRf59KD5a+
U57TGltsFukwBGfQGFlxyXYrHg4tDaqer+Via/0RaHJ5JbfBuvGUhkLTqf+iyCLn
YzPwLKWVXq5gNaIfPgzD4V35dzyeHjvjlA7UdHKt8p0sCp63r4ylTtMGkCSBt+vy
spr7ORSMu9nIe4sJb/3Z2VeSglDszDseq86I6Aqtc/T64SRMMymOYfWkmwElZgT+
N1dLeznX5ShWON3pdEabXX0K3FFuN123JL71Fi5ozBIu2WnPWPTRKx3JaYV6kKtr
lxMicEmu5KRJ6B3izISHu/tJhVGWcf0y4xCdUbXs6X1D1y4ZENzbl8nYNXxX8rDx
/wUEhdAm5u6uTm4zss9ZbYdwlFFOXjTptLJLs7wqkAOj8tLNBtzA6xhe1iX0ufv3
nx6iD1d2uo4XvUV/9csvff/QSfwbGKX/kYZQZ7cTtY9Gw2xl0w9lfbJDpVHKN40g
ZvIflAA/MDA3vLZgHalu1RESLUddrctqfeAsadym4gHI4QP6gAvCXcG/Sqbp1B0d
LyWTWG+nusDhRJXfQI2p9mjicGr6lFi63d0tMEwjxUizbRIdhlFz5WKTmjZwOw3X
9qTzgTRSC/4HaBZyKWSn4UnVwxx6i4seCHpwD16bJRNIFoQmUlcCdgie6lygMrNX
RUDlqcNGGsXPxNmjDIWGF60vIiA5KqAYWyw66ueFW2hoo7jEjzjKyDar6nnxZUcM
+X2cxeT3Vrg8Iooop180+31W+WoVVRM39usPm2wBnvrHvN+JhMaa/pY3cVDRv5H0
NAakiHiyZPencDxvyn5DFKp1cLLB79CyX81M+9DK1ISvbNeMMtaI8ByOVRlK1DVl
bcz9qd+n+Bu5/6ea+LElAhALkpuGE9KqbdJ96HKRzRQF1lTg+WSHGTCD9YArpO1y
A54KWz96xzVDUQw7maietMgORYvEFPTVkgukW/5TDWZb+B08fozhpdjo0h1Mkc8I
pKrN1mwoDr7XMCMQR+Cp2y+mkqNhO37EMc5R8CjFLxYP5J11Wz+6p5rT7+X1q1hh
v/DNcqDDY2JlV5XaHNQO7ZwNt473U0JoG9BxcdPSezkqxMprYP4MLh9f+uk25+rc
yCxsc2jWrdYcEQmNCN7XiaAO4WfYn9lc5aVPF1W4qxDl3P6uLq9q22G5qXxjjNPu
+QuF2D7vgGQH+RoxZ3eB08xI7JSn5VSyDbRv6JVELUkHot1Bxqj696Qk/GxUQqYF
dW7Cb/sQeX2P/RerS2VPbWOnQ5ujeGVoOTPWG8I136i0rfRSAcqIeqEcrommoUtx
J5ZjDVtBQdNwz0sXTV1VXGRJxOM0dS77602X8AbE2F4gwm616e0niz4p7fh1lmqT
wyFPVvkhlEojfI7MKci5tQsV3/mh6ezlUScFOyL59spfNXMQdXZYuDW83PWniPj1
w+SW37v0gJKZ+5yQsNx763LqckXiLFnUjPNv2VbzkyigQbbvbEDbsZG89DGyCGTl
59hf/fTXVQLMW80c12wdnIOBRDIqch4T61ibnl+UIxDMrtY/0GFkQyKAG7Gr3NR7
oVWABbP8CJHwoo+DgexdG2FuaOQsSX6T7+j2SOcwFU7GwJrNNQOtW9y1dtxCw8Rr
gQJGIX8jwb8Occ4eQMVSHcMB7QNO8IH1zem4VzGIyOzz2Q7aLnrUt+sZ3lqAHiUj
X6TaHncKvvfHTXIVG/ZUlErSKutBPMIobCXkZJtDPcehAf0ItgzEl3gDULqX5WRo
Ez2IfLGbO1MUXzI7kfl205thWQ3iU4XrbsX1xGEgeDWSnbBBm31QMDDq7LtaPs0B
RunnUFk4nphSWN0h/6w1hRmqldusgfcp/3ZsWicV40xGIBvxgBKj4DPlcbelOUWd
ONne2okZMT2DydU0OpZigAVNKkE3xElW4PFFbTDYE9CfeU1QHb7I67/AdcpJ6U/w
5eVEeMMTFM2c7KT868bE4owQgBU0xM2uEN7zCtHo+jhG/dQoy0qgAqL1ITr/ogBP
6oN5OfE7/nvlpcYb4kLrgydrI/wWqgM6zErPg2LQmEQgLlZrrp5jAtREtxTnuYAz
FAXSF1YA1qYh/qxJtyyijOsUJ2pZjlF/9KMNT87PDV+vnaQZd0aweAtEQr2n7+Lm
12aZRI6FGdT030WRnb4DJL1nnt/cHiq/SWCDspN2LRYjSk3JtP/4b1SUgnPno734
fop8bIPkoQzKBNuYyDJXRxsfqqtxdgFmHK1FZnL0TXSPl5vFKuN4PUhcpaE8PqC6
VW8YQyAP5tOZFa6BSDk7H03ViYm+fg/8z1/X6AOSG8W60aoioHX53+Y/uKxr8jzh
wJWvj5zjX0AYyMW+GirJJ8Dvnn4NjRcnqTFHKBjPMZHwkAAEFsayDd6Gc9VEIfF3
yGd+mzJRay1kYUHUKt51wPKirCUT8r40CwhTT5YFc74Sp3VRGpCoDVqnZJtOC2yX
TdgcxRHcMHDCVV7OtWmV8fvfIINsJgbFegDwgAT5OEL0RKzq+KN0T0jfcPA7yte6
L9akChLB7RVP/D2az+DeMHFr2McOrQUc8sJZMt+3o6sBNaO6+e1aS6K6l6W4c5Ke
ZfuLG2N1eCrORLApbhSHN0+mksuZqiAJ1g04MbLn/xEFNFq072IUukgAvmQGw1dq
R5vwkQ+vKnxj0kfG8s9YfNDTkiL0ZiVYZbSxQey7OjW+pSY935UxI2nv7bPwWVmF
9iWq6ViYlvwWJ/9AFDnMrUAhrprhvXFvpQZ+iv7lH0nMRrgq6D+L7OMLW+Ff2m76
M3Blq2YA75dhds+hL3HZpuvZakK6DNWqxtVTNq7EGd0ZH7PMk815Vb+zxwfyY7qe
ySgGQeUq2YkO0iCQL13jwKFMwhqb83XTAeE54kbXUtQrrstBD+06QeMZSgEIchZN
LZ5EfyMw1IeRv+6ViB8IU3ro1ggfPvHXiJ4/2mbLauyQPn26Lsc8iLUpFzJo6Iga
xlZTie5c7taWGLyAePro0Wpko0aSco3ZPOmFxsiqdq0XTphwcAosA10wXKgz2C+y
ks3uSo5OdTviaPLseg7Zpj+SJxhjGsRwyGEzRMraacAu/uePqqb/JeImYemzDVSz
QkAVg4j1NDZzTvDWiO0nAjB8OVtfduK8prlQZusNOBVoSU7AMFsrrQghW3Fkwdzz
/AcGwKSLBdJTJnOjzfeqOP5WTfY2rnlYRWiiD5JEeYZts0w3Nou5W7SOVFe+juMa
bA1UBwSkOYduOlcF06cmS/6FlsM6KV/1DEqpBH6/RjtM/Gqm7IedQRWNJWXHVyxw
zCPAjRLzXLzhYjtO4dEw7ziTZLQGFp3aPyXOuFIL/VVBxE4YsbzUVVYjRFjtW6UU
IJuobRETQ+Nk0J3gN5gWAWxqP7hj8d/Lmca68xzzx2zPUa1CNQjN8GJjXUa0Tyhw
us8q3uSlDC9csqIOlTBmfEpPs899uvcHQ4kt/ZuqkIFgaFXhDA67R3EneJiHg+3j
Ji1fgEyUt2bLmdMXoPFErxjXKWP61FWXCSY1kQCHyScZ6kYkK7q4deZEiTnfoqso
xaTYAQ6Jup70JtuTiKpNdYPkwKTNvDp0aJRdvXNNzX/0i70WCSRaFBefSZtfwrW7
RKZaLXA82Ibg7E/21REPNcFWXUzvZ8KP3095rXeDpP6dCGpqgBqfVjt0sUIONtlZ
uVT7CDUY5qJS8oJivPCNBVIpOekA7EOS2qKzlKkIy1h26hv2/ieg4mbn8iPuhI9j
EOGPpiRan/TRmNi2tMW0NoRBHOOgEVBq7GbfpoRng5Pqj30cXjZvWv+o+JXIJTCg
FUjR3rzt6x/Th3d8fpPjd6bfaeGihvb2A8i5kl/ZVBrMluS0Iljqx6VEgtQ4O8YV
xM153ku7EiqA9BwDsjbXAkPu13H4hl6csu7/j5yfajw18gFQXfMN8AUNbVcd7V7b
BXjNX467pr3Ul2Hf6bzDJnfSGjwH5TPW1YrCRzEY6HeFsLZwvPoGAhONRD78Fune
vlzCHgXJ9O1YLFTxeOCtD5S50agFArlFdwiBxiFoLsvVMWaf/5a2hrq9MRI0tGfv
B6pHdWQslwyK2OvJfWaYbzmr39PVKPXrSHM8sgyXvs485IrP1mosepED1fm4BQ8B
kRQoUa+V0+M69jOile0GDINu4fthzXqFVlV15CXSKZ9X2mGb1MJxOnurTrgOE37t
70rE241m8ILxq1epY+pdl1VFc2t61yBt+ktpfB6li/BpH6YdnjGxNcaW5U5CISir
qQ0kczt7BjRF7TwKrTJbOvv+VgZH74DgLbUAFVkBie5A50tP8M60THTFNbtj+nAK
3FdrFGR/bB0Rv6SfyBeMkIePJa9yzT/z/Itjqgv0xHnQYPNW+KaYVVyZyWLxnQEU
xIyjO6s3d4u3giraaiXHpFaLKNZumoVjSqR+kXgn5FQweyycMjEvF8LGwlVTHmfd
8oFZBgSqm0WZGUY+Uk+5RJXBEGCsZlSurUZgo09PpO9Asic9u4y0vgb06aYxCNNV
10whHc7srxYtCThpY6ulP0ANqmFfG92Glpz7R1Ktin/h3/sUzlX5IPIrkIIaEtnL
d2z7rvMYu0+Cm8Fjfao7+6ijlWJwrdIUzO0zC9PUiqeWwKXQEaFdK2cstJjO/8Qz
UJlYwNDhazIJpnu+Kyn13Swhk6+fNwBc/NkUDaoeAj6ryEaiRIK4A746ShLLLv8+
BRGvHi81zsF4T+lK7d/Rqj7vXHfWjywRoguaY47kpOkIESpM7umyQA3bRXp8boIH
GFX6cRC1SfbpPTXIOgoTkW3HbvdpbdtFsQ8gecHegLnZ4QwBiCje3GA0K+5zmf2Z
Z6pumRo2ffytT15sphcKRtQcRWwtOCa2M9VUWkQWF7SkT6v8uThkGNKX7gUDb35U
DvmvL3K8GHkP8Z2a4TNAPi2Ka+7WNJIQRoyVNnbcLvR1ktX6Nw3d7s/+6lQohK4f
TqHgcBPmAls1oBEi1yTCeW8ZMYxTXnBkYN85BXKuft1q7J4AwfKHj3DTQihRnk2k
3Fe1cERfCM2/ThokkYTfqjAb3vjTr3vBNTP2Sg2o+p56xM6HagHShLA5VcmozrS/
SemKycTkRDPk5kQvDupyjZVgUoh8kxh5zfTp5o2/iDewHXHRKv+3abwFFUh7taoY
YqGq0SfTv5wvYxaPC/HVGBX3va19vqeK25pmwie4JsL4FYWY946ux0gqerytrKhO
FL13F9H2Oxqqog9VflUQg6QddgLvdTzF6PqFHgvtijiFf7kR6rd37jVDnuwsWtiW
1ZikGH2HuISmIpxBd1cSWodvircpMI8rQETTMKJu4AWRL2eUfb4gBH1RXzMC/jwe
nWFyh0e4sr2BzvKnAA17gcxG7cTdbwKFhr1zEk46MsP5yKVwD1N4EtyFyZmS3tyg
sj6aH3rXGdAvqy2eKYMcwGuj0E2QhMWpnskowUryYVT67GadRjC0aBU9AgpFJACy
QfHPaZRBVJxZAKwpL8ErHZ3IpTm15cgJAbgQUc4jynaUfAZSxlmi9Cvfs2QiyRAB
G3te6yDwGDw4cBo3e2BeVLkeamnzi/YGBjaUkqNdM5bSNIs/pQ/JfPvU4SCMm9ef
Z2m4MePdNTJPQA60DZQPBjh1YUUxNU3UIJYAaAu5Yl6488bSZFCIaLuEX9TPvBap
LI9MM5jlrsFPgEE01WxMLTjnT2fLH5GskWjGq3AyHaLagtEBTlQC+szIGWKmkcyr
HAEeQNNSJxvGgRFbS6qJS7CnK0ITRYRyXDDok4P5lJ1eYBZRVWuuJXYd+N0whPe0
2hKy9qtJHPY0w0h5gYtW+EXbLugkPyk7eFAnfdwzrH13XC3RJQ7s2NujHA8PeNG2
dx0EAfTG3bYyXnE1SWKnn5cEc8AmRlZ11rIiK+EB7fuktaBcXtS+3tk8/C62ltSN
11HeOOVR33+AwXn29d09DP1jEyNRGTGQVMtoO500HgfEdnWeC4ZwiNsI2CWGHTyt
58/obnOPi4crJdi7Cry8Nui3pJcgFogl+PWuWZgRoSPRdvBydZbU0x/EDIVktHGq
qj/pU7NyPni3CHQMh5SA+bfgNGk64pxqnNxfFc4wJ3zXpltBrIPLybzuDx2ACsfF
LuFfazd1HzJlBFi0exPEdHxYCwOslLOx9a6+Dmzabq9S8ja8srKzpMa4VIB2zq6T
Ojv3hOFx+/atUooNrmIL0rwkIG8/dUfi5rcJVMewKP1oIXIEAJL9ZjoToSxt2q0b
cEyxRIWNp/Qn5nlTu6JmbHosGUW+kmSFpDbmUud/1jLvtuvY7UeqqjvDt68YCsSc
6TqR3GeOjGRiVzyiNw5HrI6fijJgKBznAQqzVT9Va8fqZCp9IxUrMjlvPeWcyOfC
7cEp18QbVNYACMHQvZudBAzTzVNy/zINy36mNPZlEWAyo/ZEhPPdTRDWWxCVc7a9
oONwgP6fuLmAs+dXhsPOaGGyfWjc1OI402M49PsSxbWrGVjLLrRYl4tY/Rr2QS8j
Ziewg7mLfkogKQ/yzGm1UTRTS6vVJ4p0TwMOU/QILs1hgTlWpeZ9BMlsnymagNxP
m9oWOpwlj2z2YE3kcCiCNwYaBhPRguZVE/StTJhKajNhIyQo/6zamkiRbLcD1EW3
3FSW/p2gk+MD2iJl+U4YF5tm3wuuflRA3ZjpN+8z6ErsUvPY6G/BivA589JhdR+7
cWvyRZ7T720sZCN/NqXSKPdSJ/kh9GirakqKqgozMYsB+L7qCzYvl8zlLXsS/GRq
6wlQNlVRbFJz9xbEY6nIYBwuFSEezT0uRWr8Un5ZcTMLhMcwSaPRyS4TXrz2MVK/
OvcMDGcHhdOqN1iFX5uGm3yz0+yoHC8PWMEhlZtFdvNdV0rMlz8gGruu+fn8zG6S
2ZsOK2ep+sI1C3BbEUim/rVRuxIEZOgsOPw8I5qYIQabM2kn3NNU93v7U4M5S7gF
yH7g/+FaLHtsB7HIB9y7sck76cZyz/vayLrTYpXdmrlFALuUzm2dry8FzrChaopd
KOz1oBudY94bHijZMVzQ/ObU70WZPIhzJReqU67O32N60luzW5810lzGbSF5YlQU
1WGBmBoNfdqMNDYGyoF1sfo8O0WJYKgM6wqqNuzi7rTUPHR6ojyf65nyz4LSFQbc
Xzin44HZeHE43ekKlFyCw0VZLQZrazavMAoTz5+HJrgLqGbq6oRnM2namx8PCWdR
yOe0x9ztJlPwFyZTAu7gpuyOXYWO3/tRVkP8DuWXH0yL9+atArPeBX2KQA4SrjjF
utPQ1NZ2G8I7IvRR3wY4C5GSsQuc3fjEHueyRq/ci95fZU+FkJUO2VpBpOPp9NXz
P+qZa3doGUGmEmaHd8JLbPQ2C0EzoKYKl9SOcpuFNH7sr98ImOnbkpxMaujYaKoG
Q1uNrFFdRpNGhtLqem3WwITAVfHHIinmvuqMczi+UJvHK+AIYvS9ja/g8tD81gaR
bJn/ibSHdUkDs6FQBt/JscOIc/LREHBvMCXAM0O6YyzWkBIasgUYuPlM5+xz041C
7LT3ABxl08Pe09TknkB6EnDrfmyvKsfbvg/q3+ttIa3fGmx1iXbxKAK1f0xzUCye
2QpfoAtkhvaZv2nDSG8W5KmhTOnb8EJoH68Wbu0zSy5exGtIImFjk1SpZWZLJshH
Y/G8SujNz+ICkMMBH0l5gSeAn4VfCm27QFopMlBLgEHZQyiK3OOAVYyyri8Vogaa
mq/x6XDBgnas+sQHMqio1kP8D420/YJc1UnLdxg3mExwm9rdLUO76wW3LBzuhSN4
HcxCs06Kfo1NvfANjPOxCtOhI56ig4s9d+T+ncHDPK4Qvgq3SyD3JDfYxOPVJ5GJ
NQdtUTm1D007YSkOf05Peg//uClA5vfgrxD5J0ukl9wivhdWgvDkEgXN7bMoC072
IobG1cFi4PadTEAtsdy47Fa2/Gec/VYH1OZbMzbEXVOoNg0EKpcEyALl2C19okSK
F4zYUSaZre4f2xzYdHCntF1TyjnBeJmWbMpCw9tl78S964ApL+u5l+JoMyaQi1BW
FfmlkFM67DQX43unQR7rFJGpGMwZ7MO5PGobZpHEDSqHceBkV90oZYBn6K13mrs1
EKLxgxjR4g2IHZVPadkHgX5f+HR/PA3mYu5l7Ge22td7eDlIMULB6HIH1hLxji/i
pMix6s6eouJQIi5Oe2U+7DrgyJYiVBkTxQPH8ppvxAKLCAG6AsdbnLPcV3Y//wFN
MfJrHc4lZRKWhcQAjMxjgukyiwUY+w8ATEAt+piuGXY64h7ukqELkakyi/1WoowE
sTO/nu1nz9mYrsDj1ZEanTQVYYfDcugAkyWjdvWt6PScSP8c91MrC9DysiPxgpY7
61V8BKLeJYLYQlWIaBmDTQLmyJsI/SO2WFcphcnszTPH1+gf7JWkqkUNNdpm+VLG
BS1f75VlcWYQlfrY1CC1LY0hkc6ir6ah9PgkBqvoypms8TLGWlygNmJz/btoqV2z
H2liTcCoqaKhQAKjw8LAFqGcTWxvWOKLRnXrR4RpGVt2IF6I/u5/sWFOxyKOz0Gc
R+Oxh7ZYBDq4k7o77/ZOv0CmRwJDisZnXZ6XEtIl0STIWWdgsfrSbxuHIw6WVgJI
F26kLe/Pm/tO3bpN2/GbOhJqX8LqUdTocSjY1z4PItuvhcAMrCAT+phi1FY8ez61
syMv6/2+BJ6SLOaC38sjRIcl+4+9fvgrgEn3ds4I5u5rpCz7O98RIk+IsmqJ+WWu
dAdZh/4Tf8EDzHZt6sGa383EERi65SswOQ6KPx2AhuGUDrGdHQwrvyX473arfwZ9
RN0g/wSBnate7FHCpx8rh3B10eY4alnLsEJDFz4KEhEgpbGbhwPieRhKPFJnZBfF
cLq+/WefjS0p2uO+pdJQpuU9dVybVrYrvAPmAKVnWPOTcHc0QyXrI40EiNIqbMkv
t9ebboMxFQYSsKOTfa385e/ThUTkxDrOoLW23i19EuMqeFu0CiiRSEc+WTeXLU8/
qFr4supd0D8OcM7+w27m9CH+U4AQ3K3ptxqUX9BjQ+a7lcC04qBGXfrp3UisQtUb
jWLVjgIlrwSlXMQSqhZHVHCGbX7zxz+j7NfkxcAZqts3mSya84pjgpvOjBb169Sa
scG50Kh4EUMAVfA+X18yIb2GiBqs5E6V7HVh6GaKKSV3Q4msnZzH51MeV4ptv3TY
YnpVnIt4uWfcNgVepEPgoHuT4xVBiKof/4JMhkL88lRNf/ucOHDe4tcZ2NDyxTer
rZW405Yqz2jSL9Bf9QHtFk8IQo7oTn5M8VEKIh8m9uXDY6NCVv4T5wcVLdohcW2U
N9XCdPb1Df39y9+w9cdHnVyFcBLLLc9nwHo5biyYuihT4fuzHK06JARPmmtvnCuG
AqyaJoj6aaC0CtHeWO83lzYcbpt5hTc2g1Hxian0R8IXFQKBeEYew7xvCpE1AqEG
k8bhpqK8uChfSa+57C4AG9XeUGpzDFm+DGASpLQqKj9sYvmnR/V0+Mvhb0fnDlhx
8l5oFzhbNpy11jNrhJHUM1q7pd45nePXI/Yht2hmNNzGXxGHV8XIwyYebNSnuBnA
4wcDEMrmbcE/UtL8bbdN1M9xE7m/JuDicbDW8s+q77/bzgIybbh/d+ayvRe4w6S6
CkfTb20/dV9vT7gjNN1JD6NXVormqGboWS4bq4UjAfYnqVkJxStlaUE9U3K4AbDd
K3sxt1nC8lOiRNbF+y/NYyEKUluQAKYOcRu4GJDgh9ES7RHqOPQVktdAd8yiPbx8
rgN1H45bd2czTMnlkhpZ/2KclntB79zhmFjCn8dd1ZTY94dEcP8kJLHMdefyoodn
EV89Lr8zQPnh4lDMZgpXvIbWJl12Xgp9hVi5LP+jDdpMNVzySDc1mJ46qeU3tUJ5
L7E0ZjRA1RdnzLqfNiyTzAFvnHAu/S+AP2ODJflIFV282RFU+m3kt6ZoPfPaOLE5
LBkY4Nd4nE5IIxAPR3JjQD63HKGzIyKxBELgnsrz6QyTwhyGZkGq8zqGvRz8EuCD
0d4bJyyO48VmmBWDhZ7d57coWe/wc16ObI8gdqvZGqogQqFIK0bDRirQqA/7YhZA
0ZVBQCM7N3aLfhYyi9tFK7J/ma6Znd7KANRRVEZhBajQDSejxQ8wNA1E8nLQ5ul3
gDt8tR2Rsj2C6QhjfdKJS6+JHqzVxTQ5Gd/JTlwiGHVEKQqcbrhGZEf9tA+9FI/8
zdRCWLvtiq9oWJweVjC+q1cXd+DRzFPRDzUlcegKN6E3es/YSvaBjK1gVovmkVuG
YvTUiQ8vUqyWt+LAJzmacr125p3TjWeHZi1yg7OUgupNUxasR2il2duI/QpU34ti
Estvz1lQGi4uvt4dfuBwb7zlOfMJpsQy7jnHXhpx16dxHuOg5/BqA+eqW41pzSgw
JQdVLX3HBe20HwdWlSZWXha+mtt0g7Dn/ysxrxQx1w6PYup/b/kYySRXWo2odqqW
u0Wqg77mvTNCT6/fo2wsCWtxUASeeqw6Tpr/6DI83+YhHk+nP3Pe3lvczi7Yocs+
PKaLzghTweuLiU+V+ZU3rJQ8D3HvU0UgVPsioCYVLzgItByzkl7bl+bUrG4sIQBi
1t3y885NXlHBvAIkPEJXQJ2fSHF1awrHlGNHlBYaaIB03x5sXe2Sb85XEaxHAhoe
6MH+kbDUaeM5RywvdVUfLQ8A9qSIH6FdXKK4pDGYtyLQJSJqa3OAnxPqYQ+qPWNa
15DLUcYyg58hfmKH1nlgTBu1QMuuiU7UmPPWjpC36sqeyzqUzjXu3juqcCR+Ggr2
A5u9qO7jJ+zuwbi9Vud6YSFTq2qlgxIk8NPr8Ti49wwtJyM2pJqCb1QXiS34coom
pwxhUO+c43W420EkZhIEPjQdTSIq2EfrnBH6PtiNrIO/hGRpHmYwnx+jhlxM0qyY
uPEJ9nTpHenhn1M0LJlzSa7yO/7ZCTnq6YyQvmwgC3wxn6CJiX8NHM8FT/vDU/dw
0Eif4j/WEsOCzpaknxHgJlL4rLC+/ZiLY1X4ubldf9TR7epWc3zZP/BxNvfilF5q
85wtJg8E5XdvnxuaDA6yboFMh+M4ChlG5vzr41A7tGrJ0nuE9PvFCayN0AIHd5gO
jYAg5okuENb3G2yTPn66l1XyU5/CXHclgzlRlalBisHKB7IrvNfs3dZeg5PVGEWT
SU+e+QRfjJAXSXlHYJBzty561tgPQEgZAPCgJ5BrhOnvNk7mGJRLFnTFyjbalSy1
swY6MCiEnyWowULpwiAAUia+/z0HbkhJxJGC780BGiLGLiTF1/Vf6aKbwDCD+ibK
krA26qf7Z6uz7CXwibiF/IE2XmAKvKwFcNMRwGeCyKMMdhcNq0Xy+T4i0EiOOcD9
xRnJNIkcXunWatHhwUZhlN9FatOFJeqtCQ+3253Qo7apuHFv/HXFoCXZ3l7Ahj4m
bWCIaQs5JWPwTHrPJvoIUom4/aqVzMj2nms+fa49F77FiO/uAmq2gLg3ZJkDcx+V
ZjgB5n+4A7p4Pbh5zdliGqXxuAxFSxkFrLToSf51Exn6jYFI7gXaRfeyfEfTBP/c
NOKUzI0Df95PSdIyqz7g8Wwo4pfhe5lsL2Z6Ep6wOqBtG65OpMVFdQUDN4sQUsLO
ygEmpxjRvIFOJhdS90jxs6+Z0uIK3ElnIAmtX2b07x2Vz9Rg1Wi7eqr5mcEb57su
llBfeq/TdY7KdIH5P784QjxSLAn2qAxxg+JpQFJhtijqhprVc2HRNCxUYloLIHll
B3p1CZQHZa7MVZQZg1f1mPK+8Nv/sF6pJtdeskv9iXK3VBK6xiS63KyBLytTEy+Y
GVk0j6QZCWNwNhVJ1BXuAeOXY8vfhKk8cbm4A4ESv4YA/Woe88XwSV41vb+PwFCC
+7c8Y1nKAltmQqheTHL4eIOGhA9akVzVHXYD1QOZKCFYuwJYXWgJsC6FKsYIbLaE
1D1DHRsHOOJq0LLycdaaSZBYYx7N4ktkR0otmoa2WAx6AKf72gg5UsKCrgTgxdX3
JxzkuI2YStKgxrfD/dgWYH7WP8JdU4quUw3xIbWKJlYoYS3/l/h1siTIINtimK23
0LW2rE56YhrKgBhLyD9r1tUBVJO5xqAf6qE0DtH1jbnyBLAhY4FKDJwWnRRdcxsg
ywiq/eszkwZXkScMY9ShFwOcQkTitl8VjTVjMj0gjzLNS40Svb82YKwYZHFvJDpi
ZpoYzQaNwyKowZ9wu4r0kJXQHCDXTYpoo6TmjEvEnviYwkdPUSACroSgAzgV5A47
YJp+vLadCRaafS5CRh3howSqB7DbB7wlnIl2bsbQdd/agrHXyEndhH4A2bORx0Ng
28RGzoJACxpc7RXxrAsaPXMlBeb6MIm4LUp6KGt89J1VMFGV95Rl89oQGYxBrcnT
JqD8QP/SHVbKcsAjSO27nl9lKHnjwJczRxXTqPz2NbV7ZJz69ZsuHru5ItyigFYA
t4hNUSrPRw+wT17SCNH2QLIbysv0lZ6D68ogDmGuB+UsoYtZMNl0Db0JMA+Axc6H
7CGSkWBkgRUx8boF+Oy12w0tJhN1mtOm7wXnjFcaeQVIRfQzH2PZn5uRbylAOt5K
cVwC51C7sCiuN1WUAzkZEzjqr69uz6vsh/GI0OYtxevFz/C8iaPu8o12Uny7Ob2J
0vgi4+v6QRsY77RI287Jw6LsdB6BlJTpLdee9bXqrG7VIyIZa+ogAloem0NW7jgC
ZAXjp54+F4VFYVhnqgu/kOL9S2mn1g2/cWUPQcX9pqeClYK/KTCMfy1eBNQXi0qA
M7qO8vRhr5r7sJLsHCYvn8Xc120zoX3B7HSX2rFFESvamDh0W5mbiBcOYvP3mMo9
/4u6ef4Uy2HydztEoIyflpMMZ+e8pXY/vTGY7tlldqBomVc5gPqRYMUTGyep5mCG
T7NLAo1/Nr+97BWek5RNRJoq5ppshWoQTW7S4rp8dYa+Br1wBLZoucPceyvF05Ro
iueRneX51VNgw0CBlDsyU42f1+a2Kn5hah0fILQgwFRziAcfecT0S1L+znLwo0Q9
4lVgt1oX/iM1E1Lhq/dkfNRj8txxj1UDhX0S6yPFnvmtd3h6FJEMK2t4cwlb3Uzr
sn+CrMW3V1FZ6LRIhj6EjcaSQWNtInRlaitt7dSyqvwq+RdFb4VYmh49s9/yLe/2
3BKhqtz2L+f67H69BpAsAFVL2WQeHh8dN3Rgh76wAG3nDDXOWpgnjpnxz1YX6ed1
9LjP0YoFsPHYLVUEv3D9BN+B4uAGwt1VRriUVbqt/XB4wKKJ+mFwfidn28yEgspd
te5iI322aZI9Xtu7Qzm5Ly2KXjS7rngSyj9U+CSX6bSF5YJapRY6xB7Vo3/LE2ZB
bEfHm6m80vcTRz/8Xyl2X0IshsZAoeEWFQoAX0PTrtps+pYyxQZ7PIJW7PFHeFRl
cSgHEI0F8hu7i8LzIpMOs/R8hCf/CVRRvsGu8ZkR87PGjFdQ77bg8r0Re+T8J1Ae
Y1QQRr38kPiymnRUCs4ym8Xgc7mh+N0UAol8zA2l0hpzwfzUURZJjEpuSaqxQCuN
kXtjekdvYXD64W09oDlY7qKT0Eam763ENyrxDhjTQ7sgmKkFnATW+nckvWoZzr9r
qx7SpaF+Dxgv2bWf+Wv+jyD1f7JZxsdisw8u1F5Xi3BIfgAyUMGnf7Z6IMp+LtP9
ndFLprXu4ZwZMahxperGeSG+XvHcFLq0hyshnSuGChXux/rzx6Pj3gfpaGiNRtcR
nv6fRzP4tGtR56hs+kR9hR/hfMQtU7Z/dwObI1vpjo2xN6REwvWzWLJSPAxifmrK
KRrqqLDaN7v0REUdN77T6KyxTuDaf4utNdoVZkTLgOjXjX0hjQ70eADWGT1pYW1u
Ikv1sQAFElgC5Rcs5JPh2i/EqjnRktStcxW2A3ComkHDOiamvQwefyuzyDBeOOqI
CIA2Gc/+HS3Lbb539c3Uyy/ukyXfeqo9AeXM8G8Y45XBeuxbHVastA4P+T2DerFF
Hjubu6u3vdKFkmLcyMySC9JiDA+VGX9aRNsxtewa37vrx/lhlwncAqleJKlCMzMF
YVz7Y4rnk0BQx8ZXwQpnH90xHvD8h8NSMfO2EVDwO7FgAnEh1GexIS1qYRw+zFo8
2TcAGo6H/ROl11nYHxeQiWldl3WwI11qmJY1hCElBcLtTkfRx7I7eLo9Hj5WL4By
WNi3oct/aQtuM0mVau3tP03wJqN/57xX5cGtq6pdbSd5HNJQtEtUBzwX14TgijNJ
VwmE7xWZBu5BD4UoPFrAB5ho5PsGDYodzmGSDWhfF0gMajxEf4sW/5QzvvM3rmkP
i3vIE/mtEDP4wmxf+SDlsvoXbDBNJx5ehAglCQv0tAQEtDp4e4QRQIl0625I4qdP
wIV/FE5yB2LDuqpS/t1dmfadgmkqtDY1smyIjqxt3nJ2KTTx1FWVpXHgyF9UrWVC
ViaCgV02ncwTwQpgP2oCR1jddrr07kFIzTzEIk2/16m+vswQ+CmU9eDD9NGc9VWT
rCB2W5C4TysUVntYQ/zmPXBmd0ysPhaimRnYlMXZty8ilauOm2XfSPLa/GosHw5P
DseRUVhe7Mm+aoeVvUr+ffi0BwMl/55UQiQcBBbKPaDAEFooccL32Oc/Em5Xiy0C
/liwVsjE98An+YdEQm/eBK6Hc1JEkPjyF5RQJna1BwLi1vOZji/lqKjUKWUHC/k+
zB969nGqO1Jd6BzDdMpDrwlsI2/GQ8zT3XUTO9xeG/aINsYPKraaf+3PO8nVcF/M
GJoLFfOEGMdj7Ahc1CiKMJrxeAlcnFx/cABh9/3aemEquIzQSE2WZ9260vSQwzlO
vODPTqGNwI8Y1SxTeRBWQeLfbyuA5pS1aNFBB7jlTPHLeFnCIXGltWqMilqWvwwX
iBbRBnodHDz/+JMpzAq73c9eZG9xkV73WZr38lDbJP1p3VhO0HKILe1H68qKnLGD
mUU5ye5htR7h1XwEwPa0JFk4LxRR3BYBbBgnP4TEu2mgDMehgjE5nIony2nMprlq
WMvnWaMN6cuPqUhC9dHIsLaDmyNUS+P/EcvNOsrU4A4h6iTmiStJksrbRSBUyDok
wCFxQiLJfv9cFKfxNKTdbdmaFbqz/fiNsyrnE85u9nW7o8eX55ZdeVKrMLuzfEw1
mA5qDHb++BdGT3YGRilxC5jMEKL1jhtBIrcCa4ZwMhxcTVi9mzg/9YI6dWR3jkMB
8ZR0g6Q5GpWMRAJBsQUaETr2izELnr2J9zHqRj32CQ6HHmP4C7YX7km7iGi4E6WA
+jJprxX0a6jcchmgX/yvDSzubBa4SSs0GT+RGB4YQQk6Jcq5mAt4P0lMxFiAGrXB
tEHvJGI9Tl8nTPh0cFPNxWNo6ZDTnh+Hju3zYAJoaaBvAIpyc1RsF5uetQp93EAV
RCSRh/17QmScoguvtKVNmBObZjJ+ngS/rif19yrhNVFB99oOiHpSdKciLKDYRSZJ
Z4fXHT1feiJ8G+LXQBLRkJ1vTRtxw7xbLU+kkNxR1WtoHUWNZCC+0hqrwvCTHetD
2jA4e1+encgfzj8VYAN9AVDrCVNJ88lbiDAMtDzYhb1+ji3nUIuEAxibicfs6lvn
ZKKYhhLpiPGFn97lcBT6YOOtXhD1NV6/YNf6+BkwEMYXJJ8e48KmrtwRlGzGF2Gv
5WcJOXhmbbdNd5TTcRL33UUBYnetZzXr4V2evt1WMBFighJvDTYXU7Tun6KvPjo2
tj3k23lRESNG96g4iBsvDa30ISCtaXzc2dP2wzlQwArqvlBzOtYcEtXWhk5BrwRX
2dUHLFJQHWrckzKDU2Ymy0/0eDO/phAu2T0rMHGVUfxYxO0ax/fQaabgNGn9vRAx
KF50VLyo1kBQ+X0PAl5U31+KuFksif73mhoAnayHEl6FnRXctjugCr8tLZwslMlk
C/QUVwi73EijpAdqsL51kmms3YurIusT5DVMJrFGeKRjKyeHga6s1e+BOXnADsW/
b/iGn3zDpxomnLZxfGJaRSuaarAk5wsTusTOUvur0Yz7OP0P5WLVMVu8AZljD2tw
8eum7iX5WGBJzZ080Vo9Bws3GLRfV3saKhoigb3O2mYir6D781iukrjeaYopiqid
59oEy9/yvfzO0YvF1yoeCSbMvGsX8LoNhlK8IOy2Ye3vHCD9l7/AfbVshRyha6ow
eiRHoseYfceKiK6ZCCpWkztA5+69pUBWCwZdL05ieV+mLY5qM4zhcGlz5+Jg8sWE
6IG++JwDmzEHpYWOpDbSw1Nkfr+m1bdVH+j59mx2jZEy0vCSq3C36KdyVGcNJNis
9UMhyFfVsEL1ovj3Y8wSVKvtFMRzdldVs2NqFn6aoESw8eNDY1NIHxPYuTPvPkjn
+zo1/GNG4yAkgnyGNiyNhX0wZKcc+8K/z2C6Xh1oFRLe/E8cl2Lw0DH9GwjE44IH
f7dWC0fcapGdvkK4KsvqjXqlYeb9KeBFUqG+HPvWkq1J00mKljvR6DOU4znqdYCg
VwCVWiJTo+/Eo3US03KUW85B8xAy0fR0S3pdTX1uiuv+jKgK9+mIGoLO2o3vi4xd
k/WQ3daj6HHJGVFMyF5Xns+in9HZJadKxqhmUd5rIQGar85JU8TlOxOCexX0VZY8
agZZfhNifPxMT5BXWG9OnxVPa5AiEv5YouBqbYkbfXaMb4jONugq3MHT+IS0QDVT
q4UGHfZQrpAXnXJ6X7WdGTJ7KJeDXk1AI3r9R241PivnILZFoxknHaO77/6KYuA3
kPHgdolqC3XnwsVVC9hA5yb/2/9D04roqDeWGuB3IZ/wzOblSrXg6kfh0ljBA2Sr
cyDq9T4XP/PlU6bV1uaH8LzMOaWfe3Y8wOpYXmYxTYUnTmBUgGhjd33AJi1vzHE5
x46Jo/+TInrTJWbK+Qf9tHcz/3vMVxBSK4AItXbDnxnlO4pFTmXtl29D4pMYMqR4
NxEEe93PUx289nkA3mhWkXDzl4WsXVLHUlgODvEGv3rh/v4eq5TW/OJdeskZ3f8/
6wnjSUzbBrOHSSpJReqZPPlh6rXcXf+avU8YhlduT7xUbSDtZzVIZDBgXiPKVIRN
uZKbWUWMH8ZmNbkYqYnNmgSZRPAIrTJEjatuh1ZpxKffPapcsJ7dy7RnJ0YC9TJs
381Mycm+sbOY/Sv35nr8XexCyAbDsgRf1cAuIlaakuwVq/Lobe5znkyRNoIawFMG
QNjwSh3yQRWGPLsC8UwvNKHY718p/4+Yrf2Bbhfncw8SifBGYGsYAB4XhAF6UnTS
kw7hJoKHo6cUxJ+pOJ90R5ZbW5R3pvsWs5gDpCW7b8tka2FJH5zBtatSdUxb/66c
KhsvWZNkHKTm3cLIql0qBXhG5E6kYTk+tXw8a1HzIEVq/BjXcsBHVHpcck0Z1IOa
mwPVoMpHu5jxtEZhq6jHExMwZMDdG7pSnlUaTlyUZu1lzsdOvOBzuRkmJxaL1K62
bCPxHpuh2aQ1eLhNMzzaJaKtrE9sn61Y9TZK244CwH2zlEYeQQ7HUfqwIftAIZec
CuUSYhzhkTxvTmLDpx3JE9va4G4HWJ5gLmWS4EQ3qgzzQzLhoLcEQupn9qd8QIzF
W9/CsECSvSTqIq1Ik0QnqMbUbveNAlyyJ7TAznwAJqMSDY/KCgLf+ZYa5BlHIceR
UEkQDHR5zfpsVG3FrI/FjI9gqD9jlZeSNTMoaysh4rEkrt7I4BcxhFNYPu/a+K0J
5fYxlPIAGLeMd5NXrqX31aNJkgq0juH4h7wCvzoDoN5XwnYMqul/FmTzpHFsq+3j
4tJ6CeYoqt7ogBsD3s/fRBWDpSQrjuGw8pxmzbr1smSzBhHGW6jfJ1ufseVBCnF5
Bf5cPZoLWiloeIPpGem9YdI3YQoHlrNK+jznOuw+msZTCRg/0twcNtOJqk/VYD0j
b5SWILhH/Jm/UxqfD+ti7hxH0z/6ZjIRN6/fWLZP7gHGUEm4CLJL/brnihG1qbfo
45B+FRFxm5knmzRzANgHu076MPAqd6iD9GXwlS5oWflpwqg8vr0JSXauWS6O3U5d
wiStP9bE2amyJXSXvY6airTgOBZGbBVVSruLbmzXrHKb9darrZJtkQmia50JnuIi
ztQq2dG0XJCChu/SFSFEnGgysslb2gv5vhTq70732HqZVaM63Qc2v8e+D2LypZLt
7kywXh2A8H1Rmsu6ms7RL89ZjlYMXfEEXxaG1kfdjfE7xMVNqVE9xNuGBLDLZg6O
8QXvEg6vCdxlIvw4Azi6kQlph8y9iW4ILvv95iblnEHwgOSQ5bUKWKfDWlMKU7RP
1gIL6AHDizklEnAV+hgYVF3OyJGrYhB83kGQPbP59ms5WTVU/twaWFjawxDVWx3K
7zRRYw3+z28Y8AW8Di1UAtD2VOfLyyDzvwyBR1+YdnJ8bO54cGazhkPqa7e/3Sdm
4868DBlmzBCvzwa4dCYJLx1Eff3YZ6eS7m+dmXrlOt++RzdkB9SM/yiTNfU53PmI
v6BkzddYhrqOp+8BRELJRVx1nQYcYPit6tpkVQFDfPouSTqnhu7udWRizNgI3eKx
Htz0DtPn9yZ32gOluvGfO5xK7xmeh9+pyLZ0DMi47u34VlYgxoAeiLApExighrPs
HpNCBRtvu+c9bCC9yg1fEhURJAVUZTObv6Q9GzCM3vQfLrrXoBRi1oTn4joVtzol
SfhTKDR/HoEoJtSAaIRec/+blCleixgNFdDAQ6jP/QsEU+FnMdAxABtB6CgC5ZHD
mKPiA0hPgQqOTU2slbmuDmAzfVwSXPZxsGQQRN7eRsFBFtPL6tUukg3KLzomAg4G
XV+O5M4X0hv0quDSO9oqFk1pAZp72Me2YpxNA0+XO0IaEer2UvXwJ/O3t4GVT6V+
TbMVHcwloOzefN871Me8zASuT9xCQ1hSSIeLaeHpudPGj6mbo3ANX97/ITwFU6FK
bfbUOXa9lsuL9UtOxiKJqPb1wMNJBbv1EIMYjqq8bH6w5r3gRF5HUaL8LwftHRe4
mWQVKehQxRL5NOYNTu35Rg4hotj629Kim1dw8RnVJPx4mGfMgX6jzw2DVLXzLutU
/tJ9a3aXzjJlXWxv7ZOpzAFb+97LNo9r5ln4D2hToreEMv2XLD9k7X2fM3zsqqkt
F3m6/jRyjvpCUR0kFCuOBy6tUUP/+mP4uHT0KykSLkl4+9rT40PjGS5O88mEBnMo
uORRIjMKe/MrrdefX+LlrQsiE7D569Mp2PyjhLiFoa0h8M5+2vpK1Nk+S6AfIj4F
ZLLPyAO8Xltobzoh1ByEjbV3jSZzVZocARwNNDx21Ep+BK0XXcMjHKfb5swQJeOB
RQ8xovf020N2KVYzy42BM9w8OKOlGUCPKvhYOhpWCZt76/XBU2d3D9rPvX+pWHr+
7F5tgEBh17+FT2SEnjNmdde+3ErpbqesSfxkutfyPT7bPKvVYIwCd6DLptUEZ1on
9gGERlVDlcVF0YmpTAIO0X5W+adV/QYPMSf9mj2S2gNFUrAhh/fdcIEqZPRCRm+f
2zCWJ9Im/tVk7eccnR5Ni1OIz+NY/fDP+rXPFcfcj2SpbmXWNC5AC9pgwfbs8U8E
BQqxwSwE0uT4EAWv794mm/IkI8zAO9bAPZITb0vnhbhHtBhKB6ujzywvrGIHDkIj
q7OqVDRrST6eII6AWzLKkOOL+VkZjrt8OwVREio4mSdWdRlM8zz3OVEW2u28mORs
rAIzqikOQDhHGVvOuo448cmLGb5Y02c0NgKhi47l1qkXYe0v1AMz1prPnsFlZrtN
dYFPt0kpdkDXq/p7K3oFa7SwwWLdcKzv2cyFw6GKE4St82NOO36uVQeaflsJKLT2
9i42LPEFGzMahMuT+BSlxWkxB3GMLTp5XW0CdsNVx2s4f9LWKV+BX/K/Bp6d/qDr
0QAcYNntKeOj9Fxq99LqKs+TIQd9lymUHe/uD24MrCVt3a1kGSzlyPCCoF8EOtGw
/1WXkNi0CUoK/uGoU83+nmZnPOT/CcLlcGhcDOpm2lHOx8HfLh0wjjVU8UF+gk/q
/HytwuHxSPxYSAX/ZapkFU5l45X2OdETtrsoU6C/QSjjeQ5oNvLFenlR1aNO1Hz3
elMk2ICD+jSLwo9snezXDvgpHPAKMh3VTBHv1N+HCM5H+uL1CSF5VlrQ7BIHnrWT
27nMCURzgcY6VhVWdfPRSyMCQI//HBkUK3g/tkFlx+OojwXPH9XsE8BIo3vKCG5q
cGWAbPiYGZxrOLkPqZMTmNUwDhwQ9U07ui0QQvwrgTqVoAF/ynsFI95VWC7owFOn
uyXoiZ4x/6BO6eOeO0YEsb9s7B3LxcfmPLXPFh5Xtq2iuX7WFojHVipPsLRDI4i/
uQZIcT6Qkr55LvstdgEAIKVuKzxOPW3NQ8oK0fvmqy811zHqpRdfjU/rF8b+Rlbo
Q74cozidQDn3OWHs0VL0l46D8hJVTB+33lnMwrToEWqdVBX+ktA/vQpFpcu104Tr
44asGNJ68ZKyKBdeuhRyNnz6IITC8Pw2hripoqJr59wAKQ/hRMRdRUxZ6H/8MNXr
Y8nhYCQlbhWfIvPdVDthxQRkKqNBT2GeGdu0vO7ThzD/D1XQPgpH5z5xq/OjEDgw
sYm8IaC8X8poGmMkxW23WyOBkkp2f8glsguVdyHEY59R8wPHzF8k3PmTPYW7m5lg
Aua3EjXUjv3+Ni0riEjhUXBJa0eAeph9USe6NO9Vj4Nsd8tIut1vF5fV6ClnrJHq
+a0s4AJgYTJzsFfTn0gw75KwdsfcGpKSpi2a+DnpmXsgplbDYOy1uZGzDVLPKsJG
rME10n9Uwo9mgiP5YRQT8LEvj2WGvZZTejAT396x0ZjroA6gIxoDnzFc2LpLCDPp
yoeXv9IHwunTnmInNIzWDVNPwgY1Rozgvua0y0zrSLj75gA3cpfwWHRLEI+6uyEh
4dMf6/vKRvYm+JYQAjJeePF2x4fJgQJtD1jZfCS0dLG6DyJvirnnXuhVu940NdO0
l12JyVT8zjzAI8kq+JMtqLIOZTvixU0KQ7Lrra6SRGcrCiHroTgTElrrS1a+5PFc
dF6eOoGfkytLDr3TtpRuGeJcECIwptJLR/lnvWdps6JuZ4rqWTJPaRtlIRlp/mZl
M7Z0cs3h3P4pZ7hNAmb6dI0AczCVrW4cZ3xZvAFE2m0PwRm3gGvYRg0kvz0AGvDX
Outnf/6taUbHLUh7a4+WPCGC4ZIyIPVki0jnJ/VQE2zchAoCDulk9PHbFDuf4/8g
B/Qr8pKGqSF8tDTUFcRwuVi1BLgDDT1pQKW6bp0nUKQeiFgPrHKbGBg78pH1JWbu
gRMFQSTLZtUj7JcdnPl8XZjXLj5rDU0VMzJb6WLPs/M30wTjHNwWT0reAeBoS+74
8x+MrhTia8fp0YyTakTxLh3S1pZSfniN3uQ9XOoVp0du3HONzUpoprcYL5f9PvJY
BfN7it+A/uEzB8h5dwb1dCkadyn8k28s7xHYFq0tmxh2EQQn8ZPWAliZwAk6nXM8
sjpRV+Yogq1ynH+/2jH+t/C6MlDLoHA9kWjrVVteRVB5FJ5dNE9sSPEYyzqbwj/6
rpLHFF84q6f/wvVbWLekzpSB7tqr5YltH/ZlMmVqqZnfcGSm9TkvV6PfJe7aw2eJ
nUBi4aP4eBMjKzTTYsCuhIOpAgvAzzd/whxb/epAsmo3POJPVPEAHvqvSqpVyWqf
bDXa3ByKaujH82IWRrPU3ZHdreReQdxF9stXoWsxKwSaRKrXBz6K1neP0YiwkQl2
RC/7ru2+ZkCQIiPxUbBhOT9NRstvJEBodtgWxgbF4fpgDdrombkUk1JlUkVQyQDV
1Ub5Cr6myEF+Bj66ebf42yry7PwBuGDykqS+Mo+Rj7+2E5s0C8x05V2rV08nR5/r
tvWAaeRKirNUrIyh2Wh6vOsocsVhOqZ59y/uYBIYgMhdm0uI4g3YRWI7ltGRa9ZN
1B60YOLFYCCPTFnFJw9yAklfuCnMipoJnJU4nTEHFV8yFso9MGJDTEhH1EVDpWES
eSHll6+9U9pL89lhURGS4NZsFxPXhZ5ZEXs6u53EVaQCX1+wouSQ55tqYXTiXL5v
0dUhIIXvgEH+9j2e3X8ZvazqTQ8hPmyQ+z3JqGM0fQSb+5gyjL4vNlOTX3wpKluJ
prRVysSWIAhGgXbeoYY+9My7HEOH5sd6qYcyTRg8T533P/+1hAyWM3+QptltFEX8
WQzstTjtHQFtHxC7rN8NXis2H2fTrtqxFyIf4WdF1zxBwTokYlPeqZbjf8bo7j7b
p1ubhMQV2eIWIiAlikpB6SJxsjgB3uI52MT5rl2tIHya2q4oJY7VwECMnDssqaIb
rZY2m1y9bmrWGhIpszBpua0gr/PRT+XJJSQkuBsRigZbwaxt8rj7zIq/1K7Wm55o
q1Xyz0KbBU0ihwME0lamrE6l7V1LmD0djn7q1jbtAqh7ELMbbJJfq78jzMKTP7gE
V6Fa6KrMDC5S9szcEhWW+lqqlogBY1pIk7Gh4+eoA1nLb2ksmvnDAv4zRDvvx3Vs
V9C+NZ0ZyxuiTLnpQru0zNbx+h3tqtE+UGF7+f46Hxt9dw3u3GjGyB90m0Ka6Vtq
dmTa5TRAoZhidpViSkfyu30sH+gjM4V7S9KEYe9mFiC1ooj5ipyuxlPo5gZArWx+
Q1VbhlvW9dUkoMbiUvzKyLYxG/RwZNTvdQmTGeQsujWLDHSecynonVeUZ8rV4vHl
uXeU2sL2upzsj+MrtZHlBNK901wRtTEaJyl/PNjgrEwAmM47WbInc8AA86ltwH+V
DuYWyD5iRT6wrxlHOrkOSqOgUhdRL/iLEYFVwfd7S9w/DxQfLtVH9XU5o9UB1fO3
7YzjG8gcRsl6Kz5wQe7wJAv1qVKE/zDfXLe18oORy5NuojNJJfl4keDd45M++OJM
k6ZA8PRO19/M2p1TUMaJlG0CoezPq3wejPW5fvk4nuiRPPikmrsX+TDDEugOHFlr
RJJwtjSOJMxYiyNGdg34WbzB96tHKoTu4IEZKKJ7rzODrsSpcQ9sroESYdJBb0Jk
gXSPusFcmmssxDH38xHI1kqIisdyqBCrKMUGz8Xl9EcLmKGBlmrzUCu/KOsm97Hw
rJqMc0VOcuafWgWanibdHCoDnpD/ifsmmqUdSticZVgcqYilfSiVR0MmHUeUMssf
YlRcmN4pqdD4hvsjhd19FwszZAdeB5lsBVm9GYTVvoHv3GYBMtF+mRPRiNQduzzf
YPlZNeuw8OoRrSen/PUZfIDWLhP4pJmAXstCT+iVZXaXecqcJ4lPNoLt0HQ4OMgQ
wU2QYCOddXBK7p09083Y2P8zvT57Zm+rEnVcBPw9ESSX1K5cBfKdMfo3SRTtax6L
zeCDlPN3POFZmtmmTdsJnJ2zLBkRF+r6n87mdQPvMyRggoThGSsdcnKDliCT87P1
vYNSe8yDhJTKLyILuSTa65EXwtDEbI7GkUZL111T4zKAzGaMjM8gFbn9u3LzgNtr
t81kb+AvguZ97dCXTlgOhDIrszk9JDTHGbQzDJoiUPg2l0sp2D1fYIX6rRlDb2ts
tVy7mkIdMlgCesctF5IWKG4ziBBzcMrRY/azIG8JqOytYqRdLXCLc+5SkSnjDtaF
1hRcINTBF7FukfUj2BpcdWKKj3SoEhHNyMgq5KBxrZ+JJWOoMxGUuQ8ksvMbgKof
jptsIklFEqFpw4OFvd0qaejWkNt8QWXDD+CgZbZexcAiOhQIzEz0iBr0K6LJhdEd
tbvMRuKCihK4rRMOKERcb0fpn7Aiv2L0UJvJmmD5pLzAv2EaDCVi00OrJKaJA1OC
YGZRAPKM9jtH83P/GiXjmbuTGxTrNdFmVIe1ybDi/WHq9FB+hmO6a/NAlGv7U2M5
hEW8RhVD/1vaWYKYwE/7snJQ5HiA+ibRYi8AL3hK9xehn4gIT7g+99bnT8C5bpjj
zPJtV1exUaTx7s8XGhfZdpUM9SJx0Nby4HKAG5zzRaMELeNAs0uZ+EHPaCpgwcD0
oXBqcGcRJV2igluyjGyHRxn9nJJBKlgYTQ1sb28Ax3RCLQQ+f3UsE8YbcalPCXcz
P4YXn5SBSEFlefYPW7HjoTKbMsclUyoVBgEJSi/GH99ZpXB9cvWMmgDDmkVzncgL
fGYWkTFRnuIeS8hX7S7LzvpoE14u8PUwN+el5padGGOsA04kDPxn9HJJeanBcb9L
sin2UYTaHufeQPCgFtcimdemQyKsQ+YPijCMyEXX+dSI12nssdfGVCccdk1pVSyy
gFHChZpql0kbkv2ScSVEssRkK93N2cSdpNMbrD7Xve9n/CHJf+SyjXlRXTwwDcKk
JaHVN4u4//24oYPrj0zIS/21nFplS3wuvakFY5kgpPkA/zjfuWPSK1dJoOE1qL+6
8CkOTeWSjqmqQwLTmkNfsfTiBvpHf7VAxxx4tDt3HsE15Hr7RurFnT6F4Djh7SWq
kRXJlKwtsE6Rxq09mEV/KM16NkGX/0N2IotvWP2HdE6K+YUvfcTcbWHi68yAvDEv
ugfr2ethQPveM2qqBDzafGfgNsGYE/Q6muHOEIh4CGVB6yptz8iT8u0Us/MKfYN4
ThI+di0J9ev5ir9DD2+dhiUBsBiKev0YLaQw4FOA9ry+WeGLPX8aj1fzvMhP222/
W3gDlE81cX3Lbf4FJOW6h21E6wALZJfgP9JM/t57LCZTjgVtVecaw51aJn4vP66h
znrSX7f7v+AeHWeJsPbzMRECflMbPe6CKeLPDZiXsbAfufMGukXGrDOBYY6HRhaY
rC+H2w4TQDnHFtZw9HpUYUr1CS5vsfVvVgKrjJ3296chSbAizAd68/UPMc9A/Pcv
4ntiDiT/7DPsFjPPaRrmXahYskVt08h3MlH7DVuEmVPoEOujR5KG9q70Wz78Qame
H6ZJkzPhzVWIp/5Vfqg4cPLktEzWuw0jZ9hqyC6Az6a7gGiuqDvrXYKoXHDTQX4Z
C6eIxNBryLBUAjzXdWW7E30LANhVQlRquDWqCTArg68EOMcI13dX9BTst0zVap5X
rQ+gTCPrnPdYRpA4n/qt6M/CMHY6d4DZNII7iUGwKv+dGa6oC1MhYIHzYejyz6Al
CywITucXUVwUargzNQBI/DL5FMnQ5D5V173UAXTQW9gnWF0VzBGXGbuUL5uk2ytQ
i5bfHx7uMrsei1k2dLGcFJQu6buoSngJ3QmysLHqoQ9plZf2y/hR51s0T882iKlA
IkV9LI1MAbzzcYuSgHFaLJzkPBr5Mtzlns6jhsJm+jV+4Tf1zAQODahbLljtwuvC
rYRbDVzAV4qr7v4XEj5LsSgcq8fVpva+bXe2VS8M4rnzKj6O6PatyePEvWkb8yAD
kdq10y8s8UQbl6Ni6hBj9baPy71JYMF6z51oJzgC3L6s4n9J361Gj0JM10FokkaQ
9UmSJgneAFZ60CcLno6tcBW1Gctbh1s+ugF2PrvP91VMAJ5fuYSYTopJA2Ho6enn
zI5oCcLxEqTxj06QUAM4uXhhbPAFZBcPc01uXdVUGENZ2VOcHtQU8f4kZU9Bt+0a
YxNIwWpBRiOGKA9r2iqQyev6qgf0fXvrkJiwg4Com+E8xAj/2qQ24U5xpbC8+Q7n
okks7HxhJgHz3ZX8Fwh9wEEf3rncrDjpsti+VBiN7nAkEcHXDvQZXPWpWbtFE53r
rINDdFR1Mr3k9dasvF8Tti0geHCIOLrt/qLDFJQ9Ynle2LCGf7GzgFrMhpvI0I3j
VXJ35DGHxkulNU33crRoVM98XY9Yl9edCceie9zhvOxI7UGHAXIs0nFCdgWxUWDy
JD3qa6MWqTommeYBCoyMyBfTc/mBEUai533+itPLmZ/JEpdt6eOb9OQM+JTixoyh
PdMhHZXEoc8VxUrbOLfFSlKya4YVQoab+5068A9Ri1zWuZ8mXqCrrndSE1OTFTwo
sgDqpU5h7hvB5jRPXao+HIOlvpVoO59lhqla+3xxQS34O34I/Qpfvwl/bdXgt7/M
1M7TTRNDyrVmBgmuigM4wT7+QOFyHIXJ/NxFqVJVDi1g4oraQnSBNL7aLPXuJGaX
hkQmQQisQ9bPCblBzLf05MZxCuATtnSNIb2O+Eg41zFRMjD+AQ1OHCb5cIb20s2r
TEk6oPlqUw4534ZpLjQFq7cyh9byH+K9ftMDcLmisDGe75eMyzglAc3SIHaFD1Vy
Mi2+jVMI3PlvGC4iPlUbri3r8r2yTWZj35lQsYCh6+tAFzfOan2493eNvTT52Xtj
G+SuaWAWf4NPdprTOZDBlkI8s0L9cqxR4mOfbUqjTGjaj6N5BJ1MxFJZXmGpx9PI
Qd9OxfN4ZSVQ398IiweyVYfEP3FurHjuYq5JGF/FubXl++u5Ry5Di2bkHs85nXWg
fGZH5hF4DP4P8pkciAtuQ5m1yiSOrAUPJRcMo1NVvMp17iTBIPe4PyvTd266P+6U
+i5dppnBEay50sqMaJjPn4PZmgoH1EaWpuYHpawWSRBRzSYzNdyzFHMYHk8r/aqS
cYbh8SzYg9LLZ0bDEK4VaF+mGPoo2sW60gZ6ynoUN0bYoUZLI9XKvpX7J9T21cAJ
PmwcHhPyPfpBQHCvvQkkqaFn1UMHquZiImMLk6NfeqtHMkigt7wDfbQNh3jBZqKf
H04PqUiWpRS3nO+g83SCg9gSEYP4FIf/bzvlr+hj6Sv4yT3Y9FNunLyZLcXZJQPR
nlofRqpr01lqBKpQnabxMPnDO/rODpFt3/Cf9VrENYXdv9tTVjeGuelLhCbMJqlY
fw7eBhXCa9sGjbORCY9rgpSpvCuj63u8e2wG7iXsrIY8+OGAMUaVgcYkSD4xh5Tt
+gcHkiU+/wwGFAaOkQLoKGowtK/3wV85uyul6LRYAoD19755AC69AY/eAP5aKDbX
hfiLrBnPj/bupaYVmyPg01hKXcJYfzef+pwyn52qjrEHsT2B1LmJOUaD85R4m+oE
NsukFInmE5h0cZgrsNtL5q/aXoSWjBtpJ3HHaHZikSBCTBykBynbmNBXvPwk2U+9
62UTXQQFLiaOUj+zqJmxNHFu+P6HQ9JANalOSafbuh9wv2MrDbIQ/nFPtS9jnWtc
JAwmj/BBsXLPKUPAo/XeqDWhp8EyadQNXK0FfZINxY5pj7XbmJTxh41DvTjnzu8T
sh6vtTjh+LrtuWUv13uhPju1fg+43E2iGNJS8ksk17vEEVOqUKpDw+71cxeD7CTQ
L93uzVlWF2eAYgJRZbLGG9o2+fbmjYhxTF6zk3/+1HrGiqMMOvJq/YqEPp1SPW4/
KCVqHvVtAG1ToJWWA5IAdggufpyCPdaJ4oTG9ZdZj5uSmG4vfowwSRqEngGBRPR7
zTRVNasWs3Wf17a8Y9FgjbFCSBFXE2CKimhDlsRoJ6pb54bhmGO1nZjmi/jhOp5Z
DnxcKtRuaoQnv5TsbqJj0OSecrSyKVTxd7O+tX9BAoiHvPJ0CODZNpGYVh/BWfFe
7KOExThrrIqbd2JEXe+FCjwkzOJa1yMKURmbHfCO3Wbv7owrUbjBzHM/IlOPSuja
2DCAYM6hk7/BGtuR7cEkLO6JeL/cw7ePH7S0Dg+Fd+YKhdZnj3lLjLdDakwBYqK4
19bffpl+mp74WwjHVxyKsvWu8YzRs+WAHIpTEiE/EbvWJIXSDiCqDi3wUhBOjQyV
ocMVgRl1JVH4KoVd2/VlUuDMe5TN+dic5/3l6JPlGvyAXhKi11R0m7bQDDzh0k5m
NH66fyFeXGR69GnXimasCHeFh3T3fUPtPAccJ86/MBDJ+z5KJXdNc1yNQIJ7q5DT
Nl9eMifZQ0lzNcfWI9knN8sf8j/uEV0Tg1zPWWvqyiT5AZR9ATd/YBDglYd7yFYX
9Fc3nBkYp/D69ftFui8OBvMvwfOKZATXpsOaneQfeXgtmzmHyPluG61DwG9FtHD+
TrCLJuoiOMvDNV6h+7uKZJAIG8tvfRVZO9M4Q6WA0k0ZGiscAs3DwZ5O6FulZMOF
omGRtbaqSYGFGXw7rUObYxC8iYW9936PaIlTvTjd8QTm+gc+lCO1AtFXbWCp4Kae
fAB8SCoH8WplYLnxzQKYqt56/7QXgwKaHItLJAEDW30t455+t1GxSnw7492kRfFz
6W+wCmwEJHwHM780vItcPvKtoMo/l3eO9FIW7RWWKcASvT2vjwYMvnSxBbNs4QhK
YZBgvhAGGsT1jpuTuo7KE6JUxZRPIZNfWxXiy3c9gsgjme6SDYECldkSg3t7xE6f
XKdBIP0x6AuhRmYzOIpGbnr2DYmtZYWiEPTtOTsNw2/7u3a+iO2RWdKOUY+DtCIN
xGMKLsqs6Ln8NU/dgAQXlyAHnpr3i7iwP2ZUr6X+45VUzyZtZKeBtRVRre8wg8SG
QuVjoB8MRuTXI3BqBcG12PMs+3ggLBfVjQ9tXbgUbf844iWTQs1G8OJNfRqfPszf
2ppSM6EEUQJj6jrcikVrTgM6XETh0UsedNYXqMbmeyF/7I0G76p330TbTVepOs8a
icMdTSXde/qlf4UqK/RvzKQ/H8HV3lY5guJHr9uC2+s1z0jnmUoozcJkYdCnyban
jzYrSP4G8jQ+TJl2uOexYTksAopwh1/nSxwyGGegpRWtlMwVLwplho8DxWyd8XLP
9BaAQR2CrqPTbwV+5wgAVey8fg2B6e3Wr9H/Ko8JaAmeFIffzRIkc+TbCH/q0FQa
y9EEh/uF9afBcurwIx93rr/cwrHn/aSsZ2q/hY0ZO9t6FpILPp/wUTX/wiqkW419
oYWB69ZuXEAjh1LucF8NzyHy9KoV/UrU2UW4S11H0j1R0X0s/Flj05WHpI3wPeuk
LcRTafkIDaKb4/MNqPVXyodHpURi+x/WsJ2i1Ska2rEvZj4Du39fzJKbrNwbXqbV
gy29ZolswHv2+QXVobB/M4UtwyopqejhG11twPHnhmK9WfTBlRzFCClvkGZY1utG
W377ZgO7rJJ2Os+sAHgAKnDSeZq6SWkSEEcyRCuS2kyOXpMHPNHa78/OMrBViKGy
/M0EtOKkhw7ISkV3icXvMMN7ONqst2ThzcCEUPZ1XDexG+HiXB1bQfyRpDN/aUXk
MzqR4x4RXxY3ducUtsj4vIJtzejoAh/Pl+WAIF9wZQUoqJgKZV0GusmPcd9a4xyp
6cY6s9T4Mq3kOnhhmf/0EK45WyfO74eyiQq/I5yxRHoZBw3xRsiQXLo7+hB/JnxR
oEc3PmLJZaEuzWfw9B5uD2U1NavAE6cdL+JwEOa+O2QTzPgF/dhnZxEyOP1R0LWI
00vUIfEn7E/WoCV902XIqNxSWpsL0Vh0EQ6DaV0+iSlI6Jg2Re3G4OLG5r3yRMMx
Ff1ggMj1pw7G3W+U7kfYls++DEbuEl+v+cWw31iYQrPAprdvIzOk1DUsAz4W9E6I
xwlkhrsO3f2vQIkgLhHt0WGdMowGMixcTi/ywfVL7sL9YRpFZeeiyA5kO2K/RFxj
lymroCOqiI145czlpfNx0fpL3+lDUuDZFmRY453YsY9xdwQtNEkABvOAqGPo9IBR
Q49Tv7llAiEzK2JV/vZAdLnALT0+RXvFY7LqHJzawVELFGJy34kccFRRI1i93G5Y
vDRN86VfCFowf/iNdHt8i/zCQREC3gdtSQW7I4/JnH5J5nOBOsaa68lmFXMSP6I6
sSQQoLB6DfwIqx/3sOJaAAC4N9As/auaEZ0p/mn53CzOquji5jPAaH3Jxgkoy4RF
9vgC+UlJ0ODGji+duvAYt/6knApgu2vvXKaOpJxka5z9wBOA4TEeeojFr4baAPys
5VpJIhCjEQbR8rB04IdojgCtd4UPOl4WpY2U5zX4pe+7Jn62Aq8FGNTkjKcu1lMN
5/bxSio00w3FVvDS2HheAw79WMJl2lRtcqtK0uC0xO9zdj3VMmAL6mzkRJscgqAy
Xrselbdouh8ZOiZqs8BYzWVcs2WTuUMffxGM4IzKIgXVZfz+29Cr3+fiU09l/3/Q
XMbxLRsUVYUkztZJxLQMZr6XOX9eAY/6VMa6x5ro43kUhWWAk6oVV1d97lFTGlH4
2xnU/Qebsa330h2rh0nzMEQMylxkHqTK3mBVg3ujVRP2nm/nsxheOwRPHVJmlrPY
k1+X5mULPLEsbf1f2Pl0SQpRbIRlEekCVSM8UlKNvk+T64r+ragCUirwuwP1GNuQ
dlJYi+mrGoGqhwUROtW7s0RNNqs+ADErb2YX5JskIl9WjpKTE8BS5PHnGfOfZ4WC
OktIhkeBLlxTEYcDoh9OpiA7aS19AohLS+pfWj5IXMRbVxbJg+7PvjN9/A8XE74f
9bwRnHbtYHo0UyYCcpmMGsSastuvUleFNAFjlwKsiSWX1xe2qphcuFNO+fEswMWo
bdViCFOM4N+kK/uyrrJffhk9mBE7jjvgYMT1+/QYcofv+Nb44/BExw3NslBpiNT5
WvobDVG2t3DWL17MNmtnOjMUpslUfnCF3B0sftVUfbPRu4jGC0QdqmJG/CloCtz9
Rc4dE2Ztaw7TVcwMCpzqdt7eMwCjTOT19125AMSXDOqqd+bnJUsHNHIQmYsKEVul
WVtUB+GLLboFQsOXQ2nHvJFUPH/0EtoSW4Zc+aBQnnyIs7ZdSpwTuRY9accYRqJm
xwM1hTcC8lPXwGtBfGXlpYoVnc/VgjqJuSDoq5qKK0PK+oHZ0g6ZlRlJS2jdDTPz
nF2YFatEC+iVTFbk14SmkREdy3qJRbkxywXYv1Geh77SygwCgFL1g3hGkjAtm6/3
apPc7Cd0A24r3Fhjz7I6fu6mmcYHn2/6QSwdFgIV75BPIipaoE811/QYNWp6vpUt
/3XEIM0Im/sPynd4ZW4+caYJEC/CtQHfg45XMI+xs8HxKGU2PiJ7s1DYes690FvR
5h0byy17ETc4oGILG81jNd5JRjlH00gcn7gt44/WDPgqDl3tQdp0QxfZ5vDYe5Lz
KJ7/NvjunYQ2AeJT2a8OMclCQxtHP+uTilCusGeQEhq3PFQv8Q0LCu4ITU+xbmkN
IMZA364bL4VRQMIoI/nUJejtL/8KSJ1tQ8YoZZJlan2aD2+GkntvvFdBY47ZUc/Q
Tfuc6ndWuc7cbNiKFTyMNPFQf1qQBvpvASch18zjuMxx7H01MdO7KclcoD/RvaPf
5poJ1XXCjgoUwLO9vNrG6dhGJAJVJjbSSMAo6ZNco/kBuw7S2wZU7GSnE7Qbcam1
9pWvXoolE2ZxeIy2ReGYYQ5Dy8QDAoyz3koUXtCbYvubTFm0+GzcpbM6V2G8Qrf4
snYX10V/9iBWKJiBZZFW6C6m+QqcHmXyCUUUYBimyZ478wuVkOV3Fh96nYKvIuoT
k5+mHcLzA/HobjgB/p/kHgbL1tT96HcU/hydBpdBfTSZ9KysDDM1d+vSXwHWO+mm
F9AsMqgrPJ/oon2mNLOH2vqOU06uP39SkuKpMBDVzPf+L5QhwC3bhgPUKrvTBgjq
rgr5XMi8sNCBC9kdzGiAt9Cscm9d14gXE3p4iaQSq+ok6CbqkB8VprMcPU4P1GX2
xeftH68YaOF+EAQrXglyS8kwT4kzFLUqOWHuK27D1BjKs01GYkp5HlqIsZUeHx1q
HbaTd7N7fRXMat8x3hKHXQLS60nwJBtmF3xjVpZ9lkcauichTI2LUc2txCoJl8D3
wJSb5vSG9stjulJEF+GWqqFBzVomEplUTZGpBTEVJuKEOZC1sZPC7CQ0xbkWwHVn
gP8Ewm6uRtyoJ5w2FlZe6LNfzKWFf3QpPXASWZ/y2BofLC+XyyFLHB6PDq2ZPtjd
q7QOxbU1DRHn/EpMKiPfMiVQK0npH6iKCmSfg+9+m00/xu0MXl1txTcC44DQUM90
WIHHdsamRpdaas384SMeDxPXjGg8uC/F/oJZc7SMBQj++sLlSRlTBKh0SF1t9V/i
LbDPrX/+bHGoJCybaIR7we0+P1qHodPY0ZL1JH4rSBp3F1kEYlhxuDnAQBfo6Z7f
zT7FrGJoZ7cbaA/lwvpicWMJHL+0ryLq3TGUfmcqCB0/Y4K0BVFvkhMIVvbPPUvP
kTHnqK6HOv65vKqOHtWjoF/xuMr6OQozuw0/167HgEWYy2gyzknGPuQ4TAXIZ1Kd
HiPRIG5RTeH19JZbOFkRW3X6lVnEREI0ekcdTSogWpTPMMLTr33PL4whWQhxSF3N
gE+lk74a1hyY6auUok05p1TNywZDog5EK2pWm0I3OIWf8JAaee8d26P/SaHnRTIZ
AIA5oooMt9+EzDUAhn6KWjhnpIfRjFjN6dNb3cram22jmgoNdg5z7Gsa1hrx5AzU
9KweE3sIdboF3difGKvRFxa98Ffd3tez4IRfbz8loPGp0QbIQRgqChF00DqU4poM
89DbmW+o2xCYzJuyeaTBTUB1vJsCXA+GPBjT9h03Nq96v0JeygD6na8h7rK746EP
QuQfoqyzv+k+9daGYQavqZBes37l5BOPKQIi4WQMXivWk2DN/zOexXzattJ4n45/
qzSTcsrq4AYx02OIQPXlmbyWECxYFjvXrLfY5ew4424Zi1gy+biONkwkNcoPB++p
Qe1dIIJxqm480MGTjSNAtnxCoqUyiorfNtvl5g8JMiHIgn5ZY8y0M89Gzk1y4Pqw
6S5WOBNC6z/iwtcfawqQfZK6X1OULlSw4rz5BSt6ezYMCKaPV8q/62MY1c7NtVEW
fO08g6XL2t7s2uS1W2dE4vTTDpjUFxXfYbMCpR003lQYZHR1fng6cxPbIB6vNRTU
xzUXV4xkggjjepVXRxS2S/ZGo4o8TNbd7WXXUhtTT/geL22yLpIf7dx4Rpr2K0sN
C3HV0ZnLKVAqahiUSEhhvsVy6/AUhAJPUPW7e++Mb4+WDmlbLhWctXPOdA/+we77
WGgKm7jMHLsxtvU7pq0ddZ7iDBJffrV9FeLhEMVAIthb9ivZE2jGQXGXp9Jkit2i
PDiWVlCsFF3klgmpdNPt8sH8Btd3FbExYO0/aQU62kiIwk2hCFjMzwLv7fh6r2oy
EmYyqYF9eVWEROrDVrOzlI94CA8zgoOXE2SGiiAqWyGLqG6od+VVFP6R4JrQGx2U
oh+7mhvOJKuC3glYmDudkOrWQbQzxDsRCXCxpRMa23Pe5paoM1NBPqiCSVB9f3ZL
a5+VgzcgYqfHRQpy2MgDWoWSJRoFSF+30A0hRm5TGKKrc1uNjuxULcNWx+OolDlN
MAuLwk0MI4shn/+lmU9aDoJ28jjK1fAerav6X/eEuQKa7wYWq1S3ttJcN8htlhCT
R2gXT4g7XeSqgkdCwvt7u5UUxEcbXRvFtfhLdtchiIWKPU4QkQ3i167XYFpr8TEd
ReW+9sIiwXJ7dMm0bwD8JYKGE3oZSvbVkHLmpuD05baQpc2kB1qVN/3BIINhOqyO
DdpiQvSgPIWc9R1z5xlXpEYXO7bdHlyia9qU6MBgRqzNbaHlq7zWOcvu2PaxWFpD
H1WGv9wveRxV+/Wx9bAFok70WxD+iUgdxTj+IMa+VeNjrTqVGVqeLvMw5kLTFzRE
uADAerizBsiYseKHOprm7MxfNM+xngnIJ0KQLkoKk27zpEiH4GrakVjESDECvrsu
NFpCrRQpr1Qj/4gLO/Qf9xxdmzOzNk96NY1HfZy6ZoHjaW3P4SAIiKHD47vfiDOC
unGgX+He9k9iCzQ+vEn6GMQFg9I8dvMmZpZfOfjMa6ZBal4BQq5mE3oiaEe1DpIF
ivc3Szk6E8uYZuVYSdlrL1DLQn1t4jtJInZQf1sanKKuZlFlTdpms0y2R0jKSpUj
Nr06M82Go0kq5/cus9jSLzFNV2Nl9QDmDJqrNXoVWAGyYwpvMIEMVTukA3Mxfy9x
AbXWueplBaXVARIuyOeS2G97jrBa4YpzwdgHsRHqDpoZejFGiWARFLRhsHj/7Yhy
bje+Y/oy7iWs5v9n2PW/Z7euFsdUrN81sMDiCsehiUpRKupbFkiG2JpiacKy59Np
EIrWrjSMGCyMN9EQqEh4OonH95wXNSU3xS7vMX/EWZTWM0wD4hBVzMfSq7PVMmt5
pXuvAnNgP4NejlhtmembNGu8xOAOFbelhd5D3BE0+K9WvRBs9QzHUtPBXpZr1WBu
cgshDngnGffpY2Sx7RGkIXI+flLUu4XAu8yKaBh8svwTTu0iiti2XKJw9UEFXVTQ
s30lV8XMSNtC2a8Y71+8otJH6BrGEJ8AAo6CAJLsGZywXdpawv1sDYvAmXI6Gi1c
VyjyndHj4X1yGt2t9wqGdDVSjuvei5sKFZDSGDcem1/qDvCSFa9WEtK9bXHhqKcb
Vh47Dvemi3h8+WAw//ReRW0nx/gVr2ikHHENpRjY/IF3cvdYVaRQQpuPfYrD2u/N
mIG9D2DreQLlkkeaHHw1g+tnm1Peyo6ekzxUjOdFMCQr2Q77AtlLEmU91KEHl0rb
QzvJFJvYd7DsShCqaSHW6AsCD3LE/hpX1gLTLqvlJ2keLsvjagAoM2AmGlG2G4/E
5kFU/bF29APkICwME4AdZsWeUPsuqiJjqJ2f910poNulYpG1l1dspJVviM0S1X9n
JJ+ZL0EHCkJ+S9G+bfwxCaOjjvRgXwwRdWi60CIYx7s12ZVT8yQdi5c2u6gU9Wz3
/+rOcIG2ocSNEEIgDbbCHcjl4+hJ2aB1eE0gGV4XWG5S82lpEMeq30Bf1F19VzbV
CdYRs5wYmgSNH9/fubgj4IXOS6iWXOJbEA9gVDWfYru+aVzUsVyZDVmLdb4A6w7C
6NCA5B1jsYT9h/xElJONPVQuc1XvBElfwUHuzBmeosZz8YwdYm03VnKQdufNqwb8
5Z1e5oSTq+/txnYdI6xLJ6yPadeK396tG3f6LUD0GDD9gWySbd9ZKZ1fnTFysaTs
zmKP8MXjRSkT038MkvlP3yztopooNMLlrXYlI9G/B6cK6OEvbsAWQH5nczAmDRK2
rMQa1zMTNqcwKrmX+NMDf628TG6kceAXfu+AtmrHH4CgsH/D5jZGWVsJhLkXspIt
dcJ8A3hrlR7EcxpyIXkRUHOOBnqHniSIHnjn2oTomhC9frhUWj4mDexIUVE3mPRa
0AoqCL2hHd5+xpPqa1pBWNCx8kBi9RPtZBVuZlgo+5NVSVX6Y6k7ymxMMV/nyFLy
Cy7TuL4e/JrEPj3HwlHZVuVvA+BPyvJHeE6AhMyQsDCSedNyB7yl/Ml/Qf/2n7VG
cBcRbFpYatxSIy/wZ+DXfh5VqS9g+ZeFrYrLmHxuWlKqCwMDiShZ8guhgucy+SA/
Pab4H9im1Ap6x/kHEbOUKxgwE//t47alKCuoljMl6h3hikSXshjg0VZ648r+JUcb
j4bTRaLiYXlhB5gADM89W37sPrksArsxmqi8wiIc+wL4g56pJ5AgxHu3x1rxe15G
tNTzkthepXPm6OTKk5zy878S/xolU2uaZ1WT8xu17EAyBps8LHplrYWXyZT8TBDG
e0GVsjDsdczXvLzm0l3TvYaDNQ54mEkpMaP7lRssgpn77jnsvsKR28i8aRtTh2Fy
F4aunIAymQPnhRVzOymDFEDm0jBBwUbtG8IgD0sSNESyst73KC27XJw8+0+QPE1+
ew3SNbW6pSNrJUi27XpRAlhzVuclaolhEcbTWvoCOQb7HaaAr4xwZNqqcciaE84E
DPJyQA/ggP1G+D8iwWl06m5Re4XgqNUsAQK6XyR5ik+TkbFv+B5EmHIomTnvKBNt
oCFRdhkIifHFCVb7nP3h/dmpBs1HaOQUbgApxlAzMouA3vddF/u/ijxZ4BQIAOH0
AXfetIGaTCzBWsWZGGH0N6pbFjOd8B2czWngB/Jq15lXoJaluwX0TJIEu6E4v28a
H226PP3UvWIYAyRhf6fQne5fX72bpOqTanzOUlD57d2yMK/AkJ8h8UwQf3dCuLdr
ZUfH5u9iHiAjg92uyiGkjnoQREfbWKtIiYufEB4ET9rg8Sv6RBICrDIeXhQD6SMu
CSiptfKBOn360xKd+CjzuCaI2xjp0ldQKFiKgi3yeVfAe7Lx9zrP62b07Mwl+sa6
5c/EKumP3RVimcjnI/wrYf9G1fUAoMPV8DWZSqG9ThjnWZJ5BAgLqpUCnY+Ps5dj
R4CxEKGaFJlu9JH0QnW0srgct92GL7W9dXDBVtppNZ6moMi6ncP9aWobPj+PwTxM
mpgz+p94CwqPW4x/gdDetflH7gIMnQTf28GPkhvz26yc218aFpdfn/zHXUOVLT11
WeBSRNOF+rKHtJq2OawCeF1kX0+T78PyeZm11FGvJ8vpnLi7nB8rzOlt/TvhA0i3
shwiHeBO+hXifO+14CQCytRA2sBZECuAysbB5fzeqY6C1skC3c62We1GD81dE/IX
qzVHQsAu8BqQzOCsrS8A8zBeCZgqxCHm6+JyliRMbVDI6YGZrzoNzYmNxMn9SvqH
qh3afZAVArZTUW3gEjHnCNS2s1d57Va+AhWYt7Yurn6f3JxgYwEf2PlzFcXJ7gKi
YdO5dOKyKetVFya/AavGVoL1UdF2eaOJIIgoLus0YNMXJNRCQlEJ6kxl6ENl8kSn
4xexoxrYovmctP7xtcJsn+V8KACkl9JTF2IGoEfhFoKCuY3EU10QpbWUa6rn5Cfl
NVsxXR0f7Q5s+49RpxH170HLeq31i0SY5JVsaEV/jCzVoxXy+ETxr+2uzOowcKWC
+B7VFb/ZQ1J2C+fAdVMiOq6zT8c3SfUHQSw5sqbHfE4A9a8yobDJ8vmciLbbXi11
PBbX94E4JvgDQa5wgCohkG39c2IMHpqGsmLYMvNMS5XRmlZ49h7TXdl0rozAPuxg
5+EKsNMRpFi0CnCjo8JnvAnHismtKNIfPMnL2JzEI4Eu/3S9R6Eta3593SUt7A22
HYiS3I7FlQFsa79iHIuDMY95z6Pe0kHdw2zpEh5xOlHqG8EfPyBpiLU6rdym85UZ
2MXgZ9MXKkAxoQc7gVXHwu1I33s+wdNPqgUSASRKfzUGbTomwwqymiQUq/OwYQXt
vodomiGkT+DGvzTjoPFh8l8kEF1aEMDjbDcFEyQ+Pbis5p0POVRWIkVZxnE96BkG
WbNROh8IkyU81lsFWsaVZumehTHNg6FvVhfyF5vDrrds5HnfQft4l3wCKiEm2WJy
CYWsPPSXylOFzzSzM2YJvuXMHFsgDoRSNfTCqy8GB7QhdspexJMxxyMBYHTVc8wr
CLRCWqC+tHcO1nXnRSzetkogUGb6ECzXRSxVqoTqBGJFRFJVBUuJiW4MeqvsTL1r
awxyJaGshq2MW7XNFZPE1rnUOv5rGU45kE1crVyLgxFwHQOMf7vOfEdKRv/S7Ss6
whKsRH33HhPJ2wQ1BlmpIOOr8nuJNFM5gBN/l+fTYGI2ai3kOos5yME261EjLSOm
bDp4cZCZnH/ZruGUKa7d/DVlw9EqMcV1ovYkXbn2Y1roeYrVKB+VYNbdBg0XrKvG
t3Ubhh2R+WkovliQ01R30G+HqEwVczqkYxFBlAZEplAuIct8RFiIzKItOwEG4nLM
Wn0BTk29QsKfu+XqWGGRD0lKhcOpLO5qj+BsJu+4hDuxCxdrhwD0znBmALtc1en3
wG2llYuJdR3NCIAD6zWoDbn60L/oZ15olDrpnehqAWGJyomeoKkRdGUNqEqJ0v+T
q8pPyOAc1zJwEk5PDzjWMxt9t/ZOEMvZ3vtbNw4TL2xlrACxVJk09Jur5t4OtcNv
ss2kn0lHuhbLBD4+9dcsDsYhlLwfrz1LsUzShQrFL5ULdSdwb4suI/H0E/ph1LZ7
EgZruvVb+Fs+PKI34lZk8PMSyvPLFIjawPddiEGBPfOtTMY5nDEUMoRvynQ/87rE
geFQC37gUJP4yXXidkgXjsZKhRhIP8J+rHXu4PCqeisMk/k5qBSGBgZN17kUU940
A4SzlTkpY/0N4VQugR3leWBeng1B6D+htPFsCWZ39Bo2PzyD57mpTbDCYTghMuSo
IpZcRqvYA4/GlVm3RaOkqtNIqZcc+J1ndT5JvrZIuV6UK2lfO4fPnxvJbhGibh1s
qkOhgEClZVPtqGH+QXyEIZmpPciPc5BVMumkCnMYJoOkJgbIvENZgRNFKSMLs8ue
SvH7ZKYdzA3IBmtOyfgPyVgpPg2pF3eHvjS05G5FBfRjEJ5nl3X4QseNQ1BASu1o
6IpQSBuZ5IIUgcIuwGjiouuZKM3WifNzAeyVyGWCmDcwfiZwqB8ue3n+I/5Owrg1
qBycq+uys9UZJJ4whDVlhgQB3AniVzKnjrTXf2zbOEi6OUyScQuVdhM3/xQ+OxX5
00cksR2xFhJ4e2vlylbGjeZgKOUzBpGQsesOBQdt33QoCVHicWN4aakXbgeL3X3E
UvGayhEqDZV2WZehOfhuIDa9E4sVmyHD0KBnbiFAZ7zRcgAXMclo3yPibvoOmIOg
6QtUudclsGXFOf4H6orEzAtEbniWa5hjjbCnZai3mU48DLAGWfgWyV9S/Rpj7ZAR
JIfTx4uXyRh/1hNAyeR4Q51Lt2TCfXbr1Vmc+VUDVMMthBlt+X/nW4sS4Cm7NrtL
caKIytFgnSDe7FN+91qqrN0xUFOqB2Gxdb8qzKzsaIhy8WH5yOC7jIYBvQk7kIqZ
Z+Re+xjWf/4ocLYwDyXzXzHBgEtqTft7cpgtCC8J7XNdQSvhug3QL0hQuEugHmZW
oKC6QBSd0NFPpn7sj1XYzB4AFsEY+SHSV7r/ApwDPtO2RCx8rWQZAhF9bBz14RHi
LPjLjuFgg3/2fJVlxn2WRC6BaSsyq7HFXzw2SCzySmA2vHBkmbQ4kreJqilStSen
krv+cZ0sdNNg3jXIWUfhIBXgPs0zqLQ5sRxOzS/6/VdaRO8kv0lYIuQqIfcHoZ33
diQWoNd0ZXU+W6G4cb3uqU3RNtqBFp7Us++ntVfCuYsvXRczaVWQwwrcKi+bWpQd
hzDBMFl5XFlYFsJwyqIHuQ7Qj7kkvtb+Z9KJ5tWxvaiE32IX6yeQpKxkSrpOLqFF
PsuTdlPSeppN4Aphmd0wFok4i5R15PEQYVyzXGOKK730iU5uUKS5dUZqKyBZ3mge
C+KC4I5NImzgCjPUqML2S+nnKXgMdG/0jqv/6jW5Fyjee0yrSUwp3EQ5WvzA0rRi
90H4ssGuW5TLZuTkNYSVCUvyJVwjtU+0fjBDiHRLnTp/zznP9s1yqqtsoYU+DAvv
fGfveuH1X8LHk1uD0sNR0hfGsWpI/1TPQ2/7z/xAIGeqcigNXRZXI3QY4tZ3+CQ/
i3As52tNtA36wAUxQ2emQs2L8n/oPHvE7pJBizkW8Ef5cpxv1JuajaTWIKg08K7p
boyELcY0PGGVTQK+l+jlIEh/cMnXIlOWHG037Id/mW+ErbmkhqCEjrDFygT4ueZi
H8pU63ySKGpsMFu/wGQ8tjPbVwB0rGneoL7bWlknfx5EO6J0u8z2XFa1MkBplwll
m4XmRoRCkDvyLZ/ob2hZqnXiUu5Kc4lBYNQYX6My2gKhcHyN/sAHtjHDejVcBXhs
UtisTMVAw4uZCHKA6kK1sSwqIxVzZzeXeuPVL22NVVDYioTa9XKkusfo4wiDY8tx
0rmKQivffkNQ6IS+K30Evk3ohde3s5eRVIrOtJt1FJCKgDx0WTARGyszYy24hk3X
4EqQ63M+iCN6FQClTj2uKMtKP06fJk5PmIj35S6jjZbREvL6W8YwmE2ZQQahxXTA
mQYkXCd8azoZYwgj822+wA837Syi/BENHiQS/Q/32LZwosKwEiBif/kCWGMKmM7w
pkcXcrxpx5KqMTWVe+WogrtUcNDJizwKJOkzfV4zUf4yzij0fjDglQZSQn/Dc87I
yD9YXOhk6P8n8qlSsnZS0DK9SpnI8Fm/GRXRX6xXDEdl9xk4DvHVKfUsItWpMyjY
hC+fYSepJB1peDXID+CymHeETbkBXVoZ+KR64G37TJaS2zEPTSEuk/dsI2pm7/b6
34PBTd1pkNH97cw1u5RFNPkAnb3kf7xCiIP5HMODRrRTYsMOAdBEYLCnpd0BOUbv
jJEjOX7wwayOG3O2roLCtgVDbUlJ8VqZa80lBooos6vSr0Mi+WenmbOxJThxDnF9
MA5jkFesOA1cYFfVBXjNGHtbyy/kuhtQ73YTn7TIG8FooVl4Eqw2gi3dCnhhMMfQ
AcPdSPHOsrb6LRnrbm1i2KCdlUHK5MSO/orUKGASTMbI+1YdqlbALssvuFqgrvLD
dmjxRPmnXwEVtZ3VVGUB8GH1f2dGt4JCMDNVUZjjjZthZCix3Td5JlROroe3tj0G
lVzwMAkY3szn7z2VH74OzDpEH1nl8HxQjc0t3XIbFK0WGATy7cT7tUiXulmYqtal
A2k/hXHesFGAuoKC9Ohr3jJ6bc4KV9GacKPBGhy8gEiCmVhnwfhgHdqNMrNGMMRi
wO+hJsSxyiu3Ob+PBgGQvAypG2h9uoIyHxChplyOrN97dYGMp/JG3Rt+vPc6rMs/
AhgneHjFQ6L46VY6GMoEfMjkKwCfJ30O7ZRj1qXtrgFW9xAMUZ35+r5Qv5VlhXFk
miDEoR3dV+yyMexDgA3bRjDfCvvh6E5Mk9dmvmZuwTlKj//RZGfVQZdT+h8s+XLJ
vKi1FzNLKsRTvkYKuVvBjiwZl1YT//vA4RwIrLI6oeWC60xAgyl8H6uZ9nfga09O
V0xMuX4X380t/s/LjuEk6GJYn0GH7sLOhHxrlmHIPt4ro5YxAPyr/JmqFzfxb9aO
KIeS17uRiyA6OPBOeoL25ewqcdxdPDX/qpo1fWvmn0kO8c6/aU6QyFAq/50h8q9C
gP/T2OX7eA433eRdwkr46GYtw5PBH6K59eVJStjG3bT9zMnDFs3mxCBhFUpMca5w
XwZwEJWOoHO9K1HxN9OBD/y3GlsdEP8h9EORuEczeyPDa4uvhty2or02On9nruc0
wf+N/ZLB5ij6exfQIno4Rm25fpH9q/jyGgIX8CjJJNjus4PxcLhx+LEfa5bEkHAw
Nh60Qq9PXu62AzPuvmFyam2M07C5EfjPX3bHkKwydHVY4p6H570ID9+EjhmVp93F
BdAQ5HvcfFTilH7oIZuhN/0rwfSx+gWoMu3rfT+i+A/JLtQUGLEdtZON6IO0yeQx
0vun8Eno8Bow7ES+d3BMAIbhKKNpGGgQQt57L88PdDpBZ39cITxn1bb+Dgd6lSts
c7KdxFAYd3zehAxKWmHlV/cXN4oaxhU+UrLVl5fCUEDk8uZSF+g0SueZenNOA2XZ
9AGzWDvhkfosHwcYTZs0oDaNVOy+cVzO2JjXKWnJIHxaji71IWaKhS8iSmH7Hv+u
p0e6az2pa+73NjFBZ7XmTRS/0trAKKq9LC8q6gLv6yibilVHkgsk1F72H7VsR5J1
QhsVCRNZOpn1uGJihC+AavxskVD49WJXrfIqpLZBlpcChWQhoPtn5m0W+6vUSt/N
UuOmZxbgXIcpQA9hlCS2nVhFf8C2osSXIVPo/Meo6xcGbtrv7+WP8XSeGDo2k8eW
F6eqisdnbpDuHxRzbz7nuRRC4W7iFYPwOY9of3s7GhRqjDlC0rUdY+kc/GSH/7ua
HT7bzpl0BJlVAIe7+/b8njKtFfbG2v2h22KsqM3mwxIfGquK/oq3sbxgB73FnifI
VXQgaMI0MsCIa+o+nXWZk8NYrrrdIgYu7k/bgZwE8cVZPfQrbuNwU4Krn7Wx11WX
CIy4y0cp+ycj1npi9nP8cTqrPVygJBo/TqFSL3KjafMY+7nH/6DehnVURILJrecs
YGqTJ+/EeHA8QUwMGTWg8H3s+4kO3gVMlloNa/IX7JDb0vC9ShcgHcpbbBWupC8q
M0wUYbmwxigVeR2/H3r8oTmNYHdJl+eXDOm5NG7dla1iEoWGP23B4rbjpZ1fAWoo
KVzwo+gF9h7ufmJbXDQD1gkqySR4wbTpFXpvk2XgXF51F751swIH+uym6ydVBRY8
IZHFDaLyTgZe+OzVNiabC5IW89EMzHmkfrrQhroZS9pZ0IS77NqKWZg0Pnediu9y
G3OsX9HPMD+hOw/Dm+XCjYY/HRJoTVeN9jKcW2+OE8/Tfc6Yd7SpFi90efNFHNX9
1RdfIHJ5648NIl5p2S+qnhP9BhA+l4e94tknkxX61f+qALvZZa8yJskrD6qBJUpr
gRCfWZsnuu8mNOlEhyxiOHlRBlzCZ0SFU0txTrx+qkawgrPxmuGz5xtdmFQhEfYo
seGHBDYLkdi1fe6WZj1bjW9B5YxwRv1O2UIDORxI561cHP9BfEE8Fla3BiK8IFd0
Rx7Nu+yUr+f6eZWlIN+VJ4qOCbj5TYW01EpToLuEPiwMpvjZNb1fS+BEhYi4Lhts
PEDbtEhSdGDnGqTPij+KerwyIyD9YZsauqaJM2UGmr6dGHddcbEQ+s/ivp8yDD1U
tYhxGn41vusqMqK8tnbp54f3ZiokkPYtEKYUvX0FdpliZApNzCXq++Tt9W0WgmgM
shBkEMj7U4UOuZxFyGn0ubqkC6z5gki1Kp+/NlrBMaMYvrhXik5zPyr9yfocwDee
v8HeU3mnHWhi6FWZsiaj6YBKuqPYuIZXdPyxiu/C62MiIFkpacEvDdIE73u4SFcC
VhKgIDl7O6/l+DSW/8X38LdmUIr67FY17LVo/bMZ7tfucHyd0464A1tR6RrqqMC+
8tCQxmB/nrzvTaBUCTM6mddFBDP3F8ih5s49/jiir/18R9rEPCcFLsM56KPjNhPq
SMQ5lBSdhngZZHj2prpr40AbfclVK0LN4BlpwLfsHeRztZm6dbyW8fdTYs0iFtIy
cV3OhtWjU1AM+lZ8kizxgPkjFSkeC2FYR3oOB2qfO+BaOi5uCRWs9ZgHMibrESYE
wJLXntGdgrHVLV0HHx4jAGaP7hAXC8igFVuRoAx2tcI5VJm+y/89kz7tQotLtfOW
JTAVVZqn2T4UXR0VFpSWV+6l6Vv3sfZXKvfxOFiQ+YCfPpQG9cy0xB6ef2TGrHJY
CX7KJFAVnfns+uATVJhv2Yao3BK7VEpPrgByWVW9j/eYZingsjIIXWjTipt+Ruv2
k0vysPyNlSBpUgKmM2MPNR9czVKigZ9Dk+P5saUn+wwarsDr6C836+zyd7qjlCxj
TCQ4WrLiRXsvjguYioLOly5f1JRibqcp97Fo+IJvSBpNfoGCoQkVm+5ipa2pmtnu
G5FaB6wTyqLuC9h+xaN7Cg+gtE9UtsXWZC7lN9ZcGWlJoGJ2gzj/v3GGae4p6Q/1
np9HcETG5ZuT70c9ynHklSX6RCunH3lZZ0DQ5auuIf4EZNft5Pk/Vmd1PFoMiN/Y
+G6xXnBVUAnqaAhNUMz7etXb2cN45imxC1FTGtOHCLszNfbnsVSa+05JexPqDz74
ZIB0VtGUwYT87S2JV5lmmw1/eKHTF41XdPfgYLOSkWP55Aj9Wat6j5yKuls/SZyC
rWh36jYftvCCnkf3ROmZ7F3/a0OezwihccY4xaGhUlI8Ub8wBynxeg0CMuYBUk7v
8jc5mR6G757N87AT07QsET1E8+WibEfk99BE2LwwQIeN5k+pKmmi7kFOhdVFemjA
4M2Gnj2/IDaa1bCAStp99wfLVL/HdOc1fv9akdmDEN6jbj7q52Brqg/hpPF0BLA5
yCjc/0pISSwe1XuOJOfqI8azx2u84dDFJUyGc26zKSPEYHKoUHjOOVAHO/eYD3WA
WNWU5t10Shict/RsnzXixxgkm7jnw7FkuKYFZqe3OZqWaWilyfRKobH4hG05O4MG
nTnUZnefXpkMl63DYs7F1+vRAPus8EhpmQ4LggJsBUtVzc4ZnYR84vpYjD0WWTrL
VSOOWT7SSaFsCxpaa9nhxU0L79+VWyI/N5DHDbOIm139y9thWKQdIQimqzhcs2Nm
s8ys1O+DXHxTG7J3V0erjhUFCciteqM7lp0O0ScSspH0xInr0CDQWnEHGvhpdvej
g0bMsBrc0MAoB2NDqfAWzscdbkmKvqFjbdrIVC0DtAjM30+F/6l7pbaqkWU0/huc
1bE7Y/kFgiqaQ8WqYxgTiB7PlzoADjqE65w/5MlgjKXxoM+5vDGQKF/6eO5WGABd
/CfLQWHjfCGrpcugl9enu2of8SYxY9GTkOm70rmMWhwzm08ua6AmcQz5kLsVYVdZ
WvikpwIRECHDZT1MiobC2DWcSalJuIGshmw46Q9RoF77e/ttpWh4DxXOlMZgOhWG
eqczmjl5CDbUKLLCptD2ESnPSBQmrH/xJ3JQ5NRxBeOh2iqcPIJNpTCHXRdfxTHd
QsAOmvKewfZ77M/SsmGkTHhiZGaCLVB52SPbz14p/whfv2VHVJtEjGyZhOOMF4LF
cYELK7MpFUkr2Kf3ucYY/FuJKmcUDrrGJOh1styZUzc76bQpr61y06KaM+9NCz6I
a8zwW+E4ipAT9RKW4Yxb6mIWQRq5JpjaikkhnGHrWcSvARAA0YZ+ZDhDqiv6Ee5e
tnNWrCga72k2fFhWMMjBgruHIdBJoEeDnClzfWO4Rv93xe3aCZ1DXUeO33F0j86X
9sonQNYszKpAFj6xGULdT+WG1ArIh0/5F7gdVd8qMD7kJez1aB35QAq9bXGs3ETa
ld2qwfV3fjFn4Hr8+smjFBXHKSLH701pQA0lYZ2XsWiQTjNCpAmpkGRstuyVxn8J
wsjflYPwBoDQ9qVlDfwU7qPj1OufwX6BQSlA3gfDd2kZb2UCfX18U4EJrIAsnrkZ
qOI6xlcJAH9j9cfNUSveuCvRqtLWrEI0sV1bxr3tcTr3kRmpuHU2LyIxqI363put
dcWTDgLxViz6i3KSFgBGV/g9TCsjAUsF7KgdwUgxz54j/8d+5bIvhZihZXk6IyxX
+0HZW7a4Z3wiKCCfJpLdWCVklapQZ+JWaL19HVDGZeTTe6S0CNFoICwld5r9xggS
bT6HhoxoXDkJyS89thTBL2XKpXZVzCF1G8VoW99V8dRC1aHlQLo5EYLhxP8l4DKx
lvzMWmkU6ix2+JHTAAaswT0HZlSyARTHwPJMdKQpyf56rdzM+2R0p0aCkyKqeUdL
r/E5mKcEWD7ac9p1ouCK5uTO65tvSX7nl9CD9Qgc2mqD4YHrwAFAhdEX/y0reGsj
PKj5iHcIWmhVH1ynEVEpvRVFhjVHqHvQgowf4jOyyXv4Z9JaYPzpnaGZ/ErGaK6p
H8IU1CZDpOy4RB4wEFcjhZQFvLUA11+ZKfDOVPBP3xEB8B9oteBog0CRU6QrcsFP
Nix+WZbIY43rM15X4lkJ7ErxMp+MQpz2IbV9S94zK+KzeiblY6vJIfKNWiBSxFp5
lpUk9sCVUsxgqq4ngc88DwK1wc2wAc+kJLiTpzqQQU+l+2YuOH4mc++dkWzHxiYX
lqNA5IUVRJmnHdTsgHeLPMMoztpgalyL185dS6Qa4fsR9/TuI0eARcgQHMRTw88O
b/+RJWU8Ehh4+4nWoh7/YFfGiGrw9ZrRYlgUygpZ/8lweiyVJWjOsNzftuzBCG56
c8heqMKUwFgrzvD3pi1efr0DhEfo7cItQhNQ0Sy849xd8jWRQkMYZptiXmguOqdK
6MJVYYufR2EUa2AlpFae0DmaA4CXnvN1okoMrACjjTDvh8fAVDL7DprS105RQ1DY
Rhww4JRGWIPvNtVZTX5a4+phaqEkCCylddypf2HkrSFlsesIJio+dmvR9ci6+B97
+npEzH6U+iQ0AcaungIMUS0SDJ61aK6W8p7AqJbg62p8MzkdMd4X1ZBwif3xYE26
eDJtQbdCiQI7LmdTVQRvEzaFnNo/guMLxB07NxdvwQG9vspD/tAgYls69IYtywB7
LwNhDN5qXBI44gdtGdAheZX7JgfFoEryc2kQXIFI6vN3xct/K/pJRYirvHAPI+CI
f4X2kxvhUnCuIB9+FtKj2W2HcGkdDmREYCLtO2WTdk8hyIpqrzd2RJfQmDrQhmy6
QXG3B+4NIjiUlHtNDYnE2AcUXp4wLheydo/xamRixvcvpaJ9XJpzXCznYeIBaUns
dXVqUg1kSn+p/BNVXBsUD1TTLXSmgNxUVYRZnKQbLcOpoHJlK7h276jxT0xfwWbi
J+lhP7Gtpj5vjomevmcivF8DodVHiGf0JWWppOfmwvwEhYHPRAS86nz8k/TVezCb
NO6WWuT+hqRpfscQXfiGU8HyvLcLOYfF2vEdExOGJyDG1PVFlqyV3iAzp3SRIBPW
vM9ROPYyO2av3htBFoxY/oSV42UkRyNRLUR/iRtbRk7Wk3PWN353Z2eF4fOjv8bk
BmhIfxgNyCFL4/keG5zd+yjU08wPTjh+6+AyacvWEVWXXchCuukahraW1B4jtzOg
iyjFDVew8fQzs+vx1dD9uQ8ENSxmmAUSwIFolXeHIg3w6tACFBG1DnQ8lXPPdYos
T2be8r+kCN4zqEhaoAeOOs5imwEZ02rPJZkE5/E7PsPAgJ3GRCliFlRk9UArrQ/R
PhcVeBFE7AU7mT+cDVY+oVpgowkhmBhnnq0yoAvoFaQTJnmQz3se6Y7cL8Y7mA9E
a9YQUmSLUJKpcSkhZRJK9r0ldRNdKT2Ea91Qk892QuOHf59NzUlmhHqYLzuxbupk
OKzVqhDMpWW+yfXIs/XXJbpkyhCED7LTmx2ydqvXiJX97ehJ9MKe7eNp/WiY4cv8
PjjRTMGxjzwmTbU0qeetljKxfq2RAVVa664aAH/NOMtDKQF6PH3mXW7HjgN1y8Xv
q7Ahprt73MjCQUhlrRl9ZdvEjNhZWyj9z5ZMA93i/ct8KdgYPZJZNIoRqyhCUHu2
HiCLHz4qfioSFEnTDJTwP+ONjNAGgwtiPbd700TWa1Ah9yWKmUpVKP3FyGbxHBlD
Nfv5wxeYJlAh15DJ+YFLc9SyMafVoVpSgIkxBNBhG+7eLfEjV7W23JK1ZcnEQn2u
fac5Zv/BB6/gQt+mmA2gAcrSZwHeZayprTRQaPuhlF2Y2pRLb70OGuNKoILYU5fG
c7M1UfHzuHSjBO5qM61WlqXVbTJDBfNmE4U1WO7KElQRRFmkB5j1tERd0vcVQKvh
3irVBUAo4fd5FzcGAh1cJCJ7tXbUo5ovJWGbw7DclPUaw+TJDt1V+P+1LwX089Wd
rV/Xc6EYTibtHvUv3rXr32LstXPGdmtbe/loLaTurFyy5n7Coz9aw7oCuBKeNZK0
/vCxlySfsT4cHR1Tr5kKjZmJ335LTsnw45+V65H9Wm30BbGN+d7bc582JS3BGgmG
tNtyxS4cERC2M5b+xf76go+egu++XhakZqau81iigG+6wBses8YcavNZu5lkrAxM
o4VYc0uCd6qWh3G+rNuJdoHEEL9H5j0nfgWewZxqNJsRkeXfhgikqyGGoutTHoWW
hH4RblEMPj3VOOhxNllERGInj5AdrMOzwNhUiOEVjLa0cH6bSExJJOe93gu+Fdlz
QLtMjeM95LIiCIb6uusI3ch5vuLkMPhPS9seXuPJDHxXlL9eSMoirgtJxYmUwH74
INRut+BIl0C70vkn3VnujY7NuurQ5hbTONEKIZwgQhVmCjgAzibGb/QBAnISx/hS
Cy47lB7LlbzZYGWN1Dr6tKdpeRvwiaXTBcAs2nfnr11NmtGupS7k+qEhc1w27nlf
tyi6NlxHCeX7fLOUUGN+zYJ9tqWHGLABgFPw3gwr6Ad/HYt+6mINbXXKShWO8QIQ
N+h9sNYp/7+MJ6g274CGkEo9CHwVwCLdRTqI9L+ZW/LgmmI/fOJz8krW5qhG5LAh
32On5bQ/EKDdK/fITE075PgxaTGitoRt/TTHiavPmlZH+FvJgdgh3XOKyhUXNtDb
uDr462b6uoG0n+wtWL+B3RaJpTLuLwM9frwa408zMFeHtJjFMO14JjT8HPIRuwW9
vZqX7W11zjwcgoojf3fvCFeT6ZE2OXEzkST20Fl/eTtxkm6WVEK9+20FYkHrvuxX
UVJBRGN1tFauuxcpvFd4tzHC+IjY/J1Gw+bfNeJHgJP83IYaOtHy9E/jpmcCknz4
oudI76hjdPOvpwWqiFg5W1Yv51rg0koXQU1jQDgVYqlxjBx8wqQXxA6xKACtBUmc
eaUzI6X4tbxnGfTB6UrQfGLnaJnfxGBM0ABpEEHNB0+kC6fzdV6t1D6z5asRnyCL
MGMJi584vXZ2LXl9Qv53Qz8OKAUrvkxbnA/hTR4mfeGgi/35mNZcmLkChW2Upmbz
MngF752EOsm3X0Zd8iN3itGiW8RBAHfCVzZV+E7UQVv8jBXa7OcqTSNcUQ/lg7iO
dmHqGDwEdY6Efw1J/R34jD3mIbZz0VVp4qQHE8sUPG4LLo+2/VGOQ0UMYNTeEOCl
Ue/p1WwdAKdg1Ejus6mG4ac03XywYtlmhsgdCamuzQVxv3Zxsulryo/rVya1dg2J
+4oAlWzx3q5ylVh8HvBn+FlzwUfOe6Vv6NDLxeqlPuJpGTm+z8+ZuWDOVnb9dZIc
/2M6g4niqdEZ4f2ig/pusMwGLh2ktotbyyGZ6VaMCcqO85Qnmw9k0wATOeR6T0lF
lzFZoPltZ1qfQBs4GpiVtl7tjR3/i1AUsQbC2mf94Iz7eet6xJsc97i/7F4GB3DG
cTNyo2CdXZvX+eTqO3Q6YNlYKQ6yKwpZJ6onXJORZzfxyNYnHEFUgSz+/lZDsHKy
Bz+ZDuD3GX88NmjVECwFdoQI3RZTizJ/qNStdZvUVchg0bAUNIStUxFR8ace1GL1
C64ORcGK3ElDo8Z+tzREkfQddp1AmuvZn84mwTv21n0X81HffuIMMoo6dtJU5zxE
CqXsm+Y0HkpC73oaGK18xB+GDj1UCD2K8sOb0Au/ryefcXlz522lGxLXg5QAjKtE
PkfdN3fKByx0XL5wTD0gYIUqz8OeL2GWCXJxbe2CgIW/0Jh3BlmMVEIExdTkqYxt
K3rqFhTbJoXjl2p5Ia+rJBfMdk/12J5cyfgGWzdSGEVdMo29C6ScFAlQYUyfETso
gBi3OtYHOnyg4bbg2ewlklRKiTzzyUYVXkJgxn6U++9x/k1cJxjrePmmSw8t10tX
A39mo5FY27d+ZagId41JXCfyV9LDzSueEF7M+euAQOrpV+UU3ghxfmA+30+VzsVp
cbvgPM/aoAjVHsQAqAreEn0hSsvGRjJ0Hr2bZw3rtaSQCtB+3/Stmpg1ijeJEr6v
H5YlWrSoUqbABBxfEQeVncasOIBd9u2SNH0hQ93Ot/lH1N2uKgkTK88ePZJFS1X0
0u7Xv7Q8BWp5+L3dseDIf2W89RjnO/KuVemDy8e9+iChx43LlVD8Dn/ywDu8iGEt
mzmdF/ToCEdF1tnpALopKv9IF2wkDbEuEiDumWPdtK2TxOcmkBSQU6QSud9Os5MX
0dMu6bL8neeSVWpSshvflqwlleWj6Sol3mioYXoqUWByxV7HEq1XfuRdKSizC72a
Kt5UBQoMfSMHTgkL21UMPLmwBVxE0tbLt9N8Mi4w+uj/hvdJFBRqHLhehmL32WTP
rNcC9uqkn7+HBDmnGGY+eBdTuEnMtmcAAUR43XnyYsQf8n3gUyy8lIhrq3keO/S8
gFKARM62/PRxf4eAEYtmtsI01Qn0TMxPaEQ+AF0wI7Z7poqTOMFykU7oxFV428nD
mQly1NlX89r1ErrCV97z8kGGdxscQere0jRXF89BxkJde60z2XF7UE29WrxGHFmT
mTG76Bb1Gs+oPLgTLO9leBjsftzR7GEabGZzUM2QVVOOntwrtOmR7cvjlZwq653J
xllJLW5ZsSVg4R2gW4rOw+HPTnsztMgriXCQmgyu6ffpKf1+ZgiivvyimHbUy1xv
Z206g6hl0UHpH7/qcIfn6+K0JdDVzk7e8YIlek7fook3VZtOuPml3UVVGEfHclXW
S31wSgaZa8jmoyNuKJcWQULNrDJv6E1Ptk+uUy84e8eBfZ459mmLJ2Z7kooGY1os
aO1QyXZoaULedXzDwR72+5TyWywcLE0TViZLSv4uFySAhy4bE0l55afJ9VgZjKDR
+8KA6KC7FMHxV82el3BPM8heGT3ZlBTSBBaDv440meeE7nBQaZZsMqbsVF4Uaa3L
w3p49jUN/+oWroR7MxXEuwe/Vs2Q6QSsp9gu7qvY55TCmkiqtbmAYYM1CH3k6u8u
e9WvNvFQRZ8gfJ7AJPtaH8yDV+O439DN4WzEBJOciLDEbgFA9PHgde7W0qLx9ASz
POJddsadUYXBn/JGmy4YF/yr4Mw5jhmLA9UB4tEZWs6at1Sx0s5sO456/e/mG2zz
uIw7rOTs8mj6JfXscMZ0UuHVH6LRQbGKpNgfxIjO+rPhVDAkOkZq07kou4L/7p3m
qtDhD3p6ZGcn1na4Hmjs3BCwX/CJw1Gz7UYPg3KhCcw4LHJrC1eC0UkwJYCS3MpJ
0yfftNqtQlUND571iF8DPGEMxkBZWlNG3B9daPpCApW+EjbUj5/YqOLagitsdn90
/KOj7MyK/3kfrrjwZJC5zGN9M2FlDRRoYm8WyE4803Z8nu+0XUafy/Z3H4VUHZX7
JSoE1bmIBIdsxXHBumiszhYOD0oRzO2FCacPP4PXTll3PjEowFEvMIC2lmGKlQNY
86Mh4MWqFkAbwbuDhCcygpTED2zKjstt6bKofwDN4Canv/AwoD8WJvajAvWaRrMj
844/47JMhWxdnT4vzlG9ekfLebXDpnhqczaWAku5q/xvYEOL7S3TfGqTvBHkJtx4
pFDfJolKvirlq0vGNQBRnb5mXRWQ5vZHmOl5HQaVVRwJClJlge/ONMcZO9Lbk1vJ
SZgLzxIV0hRkniaSvfx5OiGZUsX3IpMF4J8Tu/1eREbL4aZuAyCMgDf1KttvqYVN
O6J5u1oo/T/FVZ0Yo0nw4rYC52HV3p09zHkqxxPzvx7NjXDYWeJ1r6JE+KA/fFxE
ta8KJ0aXpTvNBAuTEw9BiEV0N7eVSlb86ut8aK9YJ75XrqVn8hxLzvlK7+WwBNQ/
RHRgxYSaIdYhf4BF0njygLA6NeSXaQ3OBj/Hmx7UjUy7pHFRQj/roev6PzwDzeoF
qL/b7D914XMmgDNMR1JMFis7qN3OG/B6VLgTnYTWWSDcWULw9x2tA/ZQmV5PeBOT
MS/ZfBgovTtosNZlIiPI2O6n0QCHIJDJrlYBzZ/4wQf9ITXVItr3Vo1zKibMj/Qq
LtdUEzrHPP0iCXt9HSncI2AcAjLYmqX85o02U6s121sm0eEdh0xuQUznUglIW4wC
ud0mgRIIPAEAvQNQ3CABxoP3Y+djBj+rv/9Hoc/uXxHwXFcGlYMcSfvHWtFF4qd1
r1nJDcDhtD+FXv5POkba9nMHYcrKd3FrQnL1KFlrNMUDhbUCJgf/LcVEH2TwiCdk
tcSnpWn4Ilhhf/jT7U9Xs/e5zujdMgmkrk4Z7f4pwnlstwyBTAXunMnXQbanEhrK
2A9c8g+89drQ6aCESxEVKIryfV2gmF7sb+byXF+DBTjz1L+jj16y5Z561BymdlX6
NdZgmH0osFJ9RIKQCoXz2//iVknLRB2qsKo7BXl9phSyC9ce40JwbfFqE0Fs3dw4
5DwmIgSq79vfHbGrvLw7ykDECYzMWPTahItxPo6hd8hVdb8LG3t6uqSBFHr0Li8M
qM6VJ8Pmd+3PSWeeML1w3ifk5CBr+VEYGAbR2R9n24M1JqWFppViu6aO2oNRQETO
H52XllOQDaYfJOzDszoj5cIFXEUEFMOCmON8T5VveChEWRC8hLC1QOoc4tQHjYLh
0yyXMtIMa3uN7s3X+3oIAzPNkADx2Yn6P6t7cg+kamUhPMKEySWG7LXKbPouO7Dw
fHnURy35deNLVFkHfrjx+vuEVTVBKQOU2LVKDLtO/7ln5Z0wbxtv/Torm47MgkQc
HYNjRWbByLqutkpp958KRIFNkTfUOrXYmIjcNsGnpbeqOY62s3n1hBvFeuBr+UZp
oso9wkAUQ51OfIgWuZHI8kNYVDVEDVgLWW8voMrePnmfG1l1LyE/Q2JmJykl9UlV
hPgIgFboSwJtMH6uQ1HFPRWBuSpJ3pggyBCWt33E+n9QRpGa9VmK7LeMTKMdC8MJ
ySedfAxd3TD2b8FVhzl2em1VhK4oeQ8iQyQZeIEtUOnPqFOHmhP1cDx+SyKQzdpF
Ivufso/LfJ1f/TtIYL8G8ZztMIgiiYvucBD6DUFCc1rbqcu4j1D7DM0qm1puN2E7
BRvb0hgtWWc6/LaeGPEtzfKfCh2cX0pLi6JZ4HSSeCsOelyxPlgT7GYVVBH2tZXl
CdAvMf57Q2gnS1qGaX3nyiM5AETdhfKIcP/SKv4TCj9/su8nNdT41n/N8ayndOj0
lHJ4aaC7rb7E17uVrQSAOfv+65P21+R5MkYnPICG5zR2Xz7/JRNiitUq/DxRuhrF
ZEW0Ht5LsiaIjvCIm5fdItpGceZADsYFunnBONHPw88NOjPeQbYN+ZtoH1UoBrSI
UNeuEE7fI2q8amlECDoe6oq5p36eRcP9P0KkOLSAKMY4L44NA8C+aXFSroJ6B5za
8TqaFH/lK0vMRrfJX9lcGI5v9nT+lhfpdnLc8qbBJPrgO0qV6tscsDteV2vO8Fwt
z7tm4rrUggfQQggskg3yZT6OofCbTRacH4fPd6+fQrMvhcLmRh1jR2foY+IQpcIM
xzKSc4Ig+Qkflw2SaCx8Sg0P/5MCQyZ6tsO46dl/ScbnifjGJd1KhZ3at1OFhzSa
PTt00J8fJyxq+oORremx5JCxrZpLburCx3bYX154SmXLjo2mCV+dd+m9gJTUjRtc
LhP3pffERbeXCHXnP1n9j6DHytPnzS0pdKu+a4K50xokpu5sFtPIBbRaMFsZq4/q
eKXatbCN6YUhIjioIzEPY2AUxC7LpXtdrsGyCCi3VyoaC03M9gZuAVpZWGCqlGII
iZ9+/yvIJ7t1tUeb07YX5aG9Di0/K5LhN0NDVbZ/ph8xSFeTrR36ZjdUXXTwI3j+
fO4Kxk0294b4BjB0/x6LOBJhLMKpaXeVBhP7N2YT4/eRWUaAk76pradnYOwFjGTC
by/3FctiEmpRZmGtlkpd0voKsyN8bM01U19Ot3i9gWbp8H9O7PEu1ozGzs+s3ESC
wuu1JlAxjx/Rz3FSIH9q03pfgm3QXtkYhFcv15mJU7Hl1cxAZCvN8ctDifHzUwtt
DQInMCM+7iXIVfXwLLfhpdFF695PeCONhbcI+JSm1+pkLRk12ws3V9pnNvKi7Rk3
Cq2K0JFqKsmwlTVgbgA9JfL1cMa/DX+roieXVcz9hOHkYgP1WJoEINGZ8Gbg7zrb
AFYKV1LColcV8L5cd8lSqRHBfZNkbuoHX2BzbPjmHO4EXMJyeq3bmC16TwJD8s55
A7BvzSU/DgJ7dRkon5/BFLxLu25N6iQktGAt6P855dwMsGG6a3EFQQ7eEIHcgBWs
n0PpMzpBica5U4IN1r4Bd2e/3dqRR6Xs32zEved71vBN3bB3dm1OFnq9g3ilrJyk
hejIfNsJbjibIf6zrABz6BTcXGLPKB/i70zzJemgw0mrClG4kVTtOCwJnj4RsiTj
VPJnG1Vhu+QoxI9j/hH7JdORQoRNvX9v37WZT2p+puZKGgaJxBkao9In2JRQBHaU
sbZlaNaOhI+MMHK4E/v+OOXkDtRHSJRz8jnegF8V72LKqflWDRLFfUz9ocirDY4F
WX66wCZbFtn3M8+kM+65Pah1agxp2WCLHqK40ZNiGxcESEklAINOstt3zhK51Ncz
qXdKtcqWoqsjhXULM4SDYJSte4AuEkFymXZLRcfeQHvRcY8FMbW7ShCdk4zTHm0B
TEV5d5KJHpdyiA8p4c78t3B/x0fG6zSL27465dGBYJ2abl5Z4aNt6sBpUJs5OJAv
PN0OZDLXr6p3cX5JmD931BoYce0ycCgGWcU+bTDvdDDYv8q0DA4ziiV2lOrAUyNm
alJJz62uxT8UZNIaYPTvcBVl4m3q/gYkdv8Kjkz6pFywlLlrshebUR0nMU5NdchU
Lk39N9qxoJEeQS+mmNqcjFo8SqTjaJ1K6DvBRrOPEUKNJept2Q2Zf4nxMMrBumxw
/2dupG4ggv6XDCASUT+Z48tUyH6Z1Wa14X5f4IviWXpQGnfbECInnPI2tCg35JVA
427hyJ9rzXsBcxcrFE6rJe2c9moOIlpA2kw0fCjNHrwtKLnTUiWTu8L6hOdjhUnM
PP30cwmCNFjrNc9dRSmwnpu5Gl+Gd9ThIcWMZjZ1VsYdzJB9l68SaZs6+YLlAmoj
bTARi3fUHmqkFZy96+TyXGZ7P49ps8WVDcoj5NgOca/yaJiG4oVRZdBwT2Is1/tn
k9rG1M9FAX/eojhCQ2QI0gwSLZi6xk80mf5Uggs98M+fiaEPhYOrsG0gulJxa5SN
0IIHAf+KhVGkJlefUvflDSmnUaBg8v8T7qtJek8Ap+Hz7gwMuxI7z9lJtK6qQ44M
sHHLzZP4TNbVLmKdheABQyFcCwAuY4L1SI2FZDogvmOgGex1bk2evmsiksOlt4zn
4cSryuLubizMV+zoseit/P3X8BZtlspYwtq0ksx+6pmFl5fVzAOvb+zq+Pa5wsNh
JcKyK/ysshHkpTOq8KW2xOaH0vxaDKFYqlGJEjPm+uZiyLX8HNmED3TbjqbYUB4g
4ixvKtokqJgMQLlWJ/GOo+y2/2llRrN2+NTTpgcPPGjTGVAxBd2tZqVrHGi7d+Xl
paeg52BEbXT/SaZSuOR/gEjfiTeB/xtDgQdTqtWZ8YaCHv9t++KF5K6ojMsikLnl
SijhaD5lO59Zf6EKrfhoWTuJ9trpfIyDP6gf7PCd+2yfoz4nDpsN9yffMxl7ju2J
XnbpYyrbCycfehuz83Fkzf/2qJsZJnCYNhRvqP1ExEV/VPoIeHG0lnAb86jRNis2
Ym8NKUp1PNeIggWGQz2DzgcMIT/QExFw+CYPtorwj9KLgNUHc93KPspbVdWLqfcN
xfMmax9USFW5Ifk9j6hzQUf08UWs3QYqTTyk6BLmpg0O/rDXUcijhvpbd+DMQRX1
d3FZX2UeFarlmzzdXfUDPYdEkft+W/fVmSEENWDpXcqDHzRMLKpcTJ6L+EYE/gxN
X3A/9E62Q3wMXk50eQUHvpbKHJUUY7xVEVn+agayS6YcRebtLFxNjoOYljP92G2A
4NDmNfrkqSv05KVgot3VjZz7APrCl8dTJ+rhtcchcycRxt/tRPi4KqAShL6B0dXu
oDCAEMpqXTWxXStDd7EVSOVX9ECzJQXRwOS5r/+hvzKioCZcwxTWIcw0qLJKgmpK
/6pgiVOUXW3q8DgGUKF4/3ZpIvDM8QofGhKopxf+VXGAfP3vtpVPWWH9OCf4Mw52
URRHkj3MdPEgMxDBKwPrzTKVK5oR3ipSvB4PZUPww0LM4Ek1TwjlR3XgdlPyQ/oQ
vHJO6ywaHAJEXBpNiYkrwzuoTdn6oQ3cFY6AmUzwzKGZfNUmk2zMKhop9cRHtOD9
tRKq8T6/J0zSXK5Q57K3XCD0zPzEviKE6D+ZsSut3WPNRQyIaSW1c9KSbDIduNbj
AMvKRYXutsfM0yXIJCN+zJLGLlpgNmT28u+Qm0N5AvGHgPOQlh4c/IdhJPJ43xDF
jUJ/Rry6qu6dDv3a2iKcmqSRzxyGk5ghvGdPZI4HAoh+2K88A17JcVnF7tNSBNR0
9Pp0KNsnVvpClHiebklYJTi98mD/eOsFUou5T4m0ItjdZjZK0gmzNE+4n+A0CPBm
CnHQZ/UcJ6BXqsRS9KM2Kv/UW+egYRl1d7PK1Ovnc8z4CfJMo6sFb2eVZkMtuXTf
vTt02UXZVvHric4oF0PcFqmvAUn9TIn1VDB30/jwNnhbAnB7HosWbYma4/Fb18Kv
VnrqOGy5kWXBfMdmA4wbjeJXBjjUTZyRqvhN2X9D8jFurxOMv6X5+4CkPtkqBBYS
9PLh4QFLkFtgOEgbHxe7OlWYbHQ8WbiYChclSXiugbpm+ciTAsruLPUKExpQ3uYY
y8vyC9lVqSVccPppNN4dFWTTYLVdrYjIAve7LgyHiCUitLkQu/73Nmrs++hpNBgj
A+jLe8q1LH6YGFc1tLxfZxYAQYmT8Wo7f3sBbcMoy/qZM60rxhtE3n88sicjePYJ
l5bL2FdwlRNs54wvWj0hOOJC+GnRiYbphJs5BNiZjTLO7T/jVHPZARsDY3XGdk0r
iUZR9EtkfQRjKFNgg61pM7lQXx3QHT6raPBVJgE6H+KE26Pi2Z7R5dMvMDE9W6WS
AejXNk48hfs7uQDI9EC6x6OtOGENOoMUSkIFVtvghGUJlDdqxFHbwPN8Gca4YjNp
W/m3KWUmqUZUir+4INtkRjVcaR2HY7+j1EoE/VnMAV2Yt2sNn8DAEFMW2uzY4WOi
uKlp8db+yxsj6M34lx5iCSFW55NU6VbUIif6fte6p3Wy8zi5Zs7zROerwpBmFwQO
XnlOm4Q3buVeFLvnlvflCdc8aNs6fxD5sY1Nz7jHF+UXlguMpK4sKlmJFxTSPG4/
v7hvVpSHxrwGArS0hAIXq9O138h5EEOLMv6nT2bOLSG2eV7Fbji/luE87r3oj0p1
n3AIMy7zYsR9oU7sDD9FUxOl0wk/7jRHPGtZE73nyojJmFVT1x6e6dtvz/Y3GNpQ
94krs+6Q1Ah4OrDhpu+GlXicuPFMPd55UeM2oRs+7h1Lqz/x3M4ZWues+w4RlJRW
EW+z/8yPphMtYVQQmvvUVmTW9+4QK7Xy2yGV9bAxqJ8xd9d9CG26OYxnaCZV6fuZ
2NPRl66721U1hIZ5BDGvqCiYYtRWxUObRRKGJvmQfWaIYU3ZSru+rzjkqGXRUPpr
xPQw8hwPoUjzD1ebtFYUchYgzK/kmlJMJofjq6ann+lEix3hD4hi8u6duSk/xDWz
bbyI7nu6HavewE31NRRigqggXNXMmFGCih4w8Irk0+9gqcb/4ZZiAhQeW5GGoPEm
cuxUgtWSjYUnfBll6Vz+Jfx4QyaKukwl+ERF3zHZSVzympd8oz5lHyjrJteLFRss
d/BR3LbDaFkrNwoJX5L0SWfjV1I3xbjKE/zashmxtdbLRrr6ph4zBXi/OMk3JQmL
Qm28i8f/h4RWD+9RmlJa4HpjBamMt3SstO4hzBQPFv5RfBpc8kUR9MErN9mmvBBR
okuEs3wH+byHwhgyae0y1Y9VCSS0PknXYICBMu+WhvKSjX+0y/tXW1b5cV0P8LVH
NInzqz/qfA61KeEVuD2zTA1/MMIyHJjKj/0w7Ke9RrshHBw22jGzX038ia46fryc
CHQcJXi+kfdiMbazg7ux/6vu4vnqOFsZXay2an7joZEEa5zxIZgOdqDonLBsQkyP
Ui0BCNgCT16NuTbXDqGl1BKkqx70/FHTo8gxRCVcSBqgXb0Ih2/ihrSfRtJlZxWX
AnxED9emsvRSkrD2yiBd/GCL4xfHY+13/fFTCDBP5h1i8uESF3E1ZNNivXHScvRy
uoPSdBjxLxQrkbgm3hpB+Y0MzPzJo5RjZN59gZ48pP1RstVLcXsqJddE9pmXVrns
kVxihLc0aIpeZ8hqeEMaaaJlYCfiNpc5yTZclUUclF45dPSZZzWPRKilgbZ0whvb
hCdjjUvy36Mc3WYzCqCf17JIIU4wmDriMtbZUca6o37z47qfF3MjshD11VZd/KJn
Kzow+3muUk2ZHdjk3HUM8WCrDUpgmpTyItvpaLeVxrpggIK+lqL/CofiwEo5370V
2udrSPlvxkXdYbSlClt+CHGuRjM3Kb7BKdlc21hRvXvx4uNfcboSw+v0DDCCkhWg
9uzs0Vhs2b1Umd1YQdM+jdvWNL80T/eR0CiaN7DXqeWDphAb7CRkCCFxFrPRqbES
a/tUtcLqC0Bm8JAlQrTTCxco2E00brtqGfZyUhlIWdoL9RenKVvYBWmebymyGch5
+GKqmP5aDeRNvZ6mcYT2AngJFCE2t9COjJfgP2nJ5UJAlJF7sqLZg+a33jaH1JP2
d4rr4JYWSnnK4Z6mdDIHUoUqjYFD5NMH5YLHmy25aTbrI1y4K1k8/p1Y8NGI91zW
zNuNLJSykIwUo/6+OI5ozWUki+wf7yiX+RWI9P/xtvFmwUno9WcW0Zzn5wG/ezj7
ClBJoR7+eQLvJ3TSu6+b53Qy868XYwzB461JLwQpcDtECX3pHFQlJZSOtqc7P11E
mYKx2UOaonJo+/EkIXg0HhWtIqxq2HgU4kNqGLWq3UB8zWRV8K3z88pYlZmF2UC/
ls/3rmMNE5y9aaxvVGRcdaRYCPOAbm13ZWcUIog9wTqVYQrKCJdIdUyH4P4rZtd3
jddmYRn3WwBFK8aPlbe6t3i9pCpRhOWNgjRuU+fNxXlEy1kI+ekaxOoBtpnIstsm
J92MBaiJ/yzPhaM/QPpu4bTweK2JRMQI+7RtDi+0yjedLmbqp1NqfhaZ52H2/qO0
EEN66oXpM1YQw6Y+ZU8cRu9OR9hXNKXyzu19RbktVFWnFUDsV0zpqDy+0ghx0Nzs
J7m2EDtA3PK/XPbRr3xFMt4uGZQtDdGVMM9AAfWauGYyZ3FOvEpNeoeVG9ERy/k1
HXJCntFU1DUlroS7iY7MoWQnhPl0B8gTozeGvJ4eBNJWuvI0xnpuzPtvu8VPznH7
ykxNVjUY0dUChK71r0zbWy4a56P0KgF74NdHn559ub1hQymbqEodDIyddHggTZSE
6jICd1LLdlGEMIuBPsMWGZnFB3Q6iOOjdo9K7R4dlvKVaHAYKh5sDMEeaE9spgjl
02UP0s0jP/UusgbZtuh4u/1uQkM6QH7KFO5lj0SnUJEqLSq4ziEtSPzluirylKL8
SmziHGAq6LNYwBmsATHyoWy1beuaW8M4ci+V0/kBVJoFwAFH3eAJLMaB66G+VyIL
AdhJ+KCWnP4qh+I4SH30VOOkzj/fIRHeJySk3aYeRl8KpqtHWirQ2Z/1kE4SU4H9
LJcWbUcHKqJobeOJzJePj324sCv/9c24xJv8LMe6BD2fJcjMthscJxD0u/itLFgD
Tr18xfwbJUkvqv4yExSOOsDYDGPg203rDRt2Dns0tqJijQccQC6aejII0ynMUUa1
dhH6FWimmf9Dbyp7JIzoCNmtSqcnhSSO7xfED5Zdw1DFQpDoMfhM/5+fqGxHQewb
p12omSXgCf4iO4iK9nAXdHydvP+sm93XN8+yrNqzjatIatMftGxk+biNcpwd+ret
AjsSNKeceUYy/rQLWDJYA8FDGe3Wt2MKEDx8Exa/imLY7tNNKGJQq18c3ccslsZx
8Sg4gzrtMTQvjV7SIJJmmHSZzWyYM+cZZkxLX8TQJG30i3PZfVjFeTZrxbeaaxsr
7TGJIpGf/aLZfmyKQ+EHTpsrLmVsWAgl2F2RmHLgaM4iazQjPvQL3jQZ+65KO/hR
gUx1lFqtO+qrEUpoo2WUxkb8FBjZlBSkHsq9NJwK1k8M8dpXiyoppuGcajZqOef7
MGbcPrzlOanZoHrawuGEkvQtw/Fctu7UNZcWf2sAFCaPvY4joiB8PZsYj13/X2if
8/THRpmoldXULTI2Ebn9GjiqEOY0rwrofpqKgKe9ZH9dUZ9Lf7mZ8LTA0rqXSJDR
6mOMNoQ5Jx7WoTsaYNgLuOGPTYMuDRbEv2Fc+aifPsvuYIJpmoCiQ/U4meoWA2UT
WuP1qz/OmtoSfd64EqY15sIwekFxjcLxTOieK9BwQNTYKb+sOVJiB9uR0YBTuEhX
4bquEDo+M2v0i0Gvg3SKEWNSbTF77Qk15HwXGTFzNsZFtUDNbLkHztFqPvKrGtoI
UhAIT5Pjfh0TPvz88PFBbxzXm0NSsPwYd8VUeCpBVtIKbNZ0CxhUVNK9kIYDbMbA
jWTC+oaTMA9M9G+c3f5GwKBN6nOHbuvYi67vhYOsZnD7rJeCyUmavRjIVBWQ6gGN
RWzQsgifGW5FP6EorDSY4a6BOU/2sBvA2EipG9UoYeM/UPpOtf4ARzNqj9KuG7El
2pCGXRrbKwI66WfLwBI67GXMoarVHC2C9Uoa25f1SLvS0sInYgv9aaY4Yis5EumU
iH2kAkp570CeLgeaQ31eu+RCz/IOoeRAOnZNkzmeIKsxV1xv181dj37MtE1Vq9lL
bVnM1z61coydpGKFdbwH9dHhb/5qKdHN8vb2YLULAowS4OxvvN+yE/jZlqFOeP3o
48RvkZpd/4irhmsvaH4yZ5hscyoazzCdmA0fTGf8TYnU8oZ359h+z2oGjbmKU6nc
nURpls1EhTRX2YyKEuQpVwA2bUjYz1rfUF/I2vOqoJM/DEsKCxz6Lcq0jt1ZiXTG
f60WJ6vOar7ThcRGDvjRsRucl3BQfybRV929pFdv9wn1VrR396tlJRhRTZPido7Q
2099rnvU+w+RXoIxwJ2sJ2slaYrnmqnhDPXkjI3elgVvTxlK2aqow/s6cQy31Bzm
tLMUu5RvmA1St/QogrZslYo7rhBCt5zzG+105+C76GMjECyEEOySqQ//LhfPw2J9
1yA5kjl/cJ5TvRMmTcKg62l160FzIOoOhWbmpVE5xDqynGx7LCyfOawWNyX6Wpjo
RJSsqkCMJAYzP3UbL6kUklpbUc6YWEspGVpLZxhqiLnCA9PbP7qfOzm7KdWMyBmL
GsiTVwiHIc2sS9xylLCnI9mO5HpGlnDgTiAn0pZhjkerFiDZVOxQHRja2bsO6Nom
ltgCIAlilRV9aw4okaUvWpiZU6Lgn0P8a0t+sQU+JlO5okNGU8CfmnqRD1BfwmHR
LkmlkfVPIpGB1AEDL2F8mgDojtr0TqK3g6o+pbGWfg8ZRX8X2sRxLjHl40zgbsYb
naMX13OBqcE6rD567PYZYgVBOeQdSjpa0uMBkJzEpTCw0x7Sm5xVRfoflEiKOTk7
el6xmot9i0dN+ejkgv+nbmUPcsrABbDn/ek2Tsbdc5pWhLj0aHAw8s4EWmz3tcXC
lNQ86tuXIzGlpx8XN6uZzL53sYXTK7TQsbiHnDc3df7noA40+75lHxocoKNF6p+P
Xdj6rIybCXwBQB9/SbAjxJlBe4XlnYY5YFGyoIm4yTMuvKZ9jx+1JD+pv3CmNUIQ
vvug2yQYz59m8KbB0S4Nzf0m+iSPmZei/VncC52Sd3RyaxqxN33LiHEQrboAW1Jg
piWe2YhCQ/Cm14C4kR+/RLxjNwNewZwKdxayFj3PqkZuOoxgLqKEzv5B2D7IppWh
nrBJ4PSor1Mi0XoU45n6T3TUn2aSt3F8bPSiNtcMU+Gk94/GptrP+RrGfYppCEir
VtfxXZkYq72sygBImmSpyezQfGja2txwXAYz4AtmicTTcD7coL8VFIpe8mX9aA8H
QLWj3vIjr96e3uB/Xg84CkGiINt+PINnHXRGqgbGuOWtHX0vbzSEVaz3qkgGZiRW
cVOrHpbyuyz1mjk64uMY8coHRMlucZ3HjHP2PbC2AGmr0NNktVscPG9HkyLJZInk
Nx2cz4MJqx1j/898jjrlb0vx3SKTM1+UlEH8rfsqTDJ/nTrisavgjDoile0l+jE3
JS0b5F2xSBzbOE08T27tX8pMbe9X2E3NzPWeeFjVa4dL6jtd8/JkAhXzDoLoM378
RHdRsE4ekIJSBo2D0CBtZaBtmoKzWkYvia8JTQZhkAiLLE60M/d65goP9j+BcniX
GZMaIQkwl1LCtFv2W3ORb4adb0CO21w2BjYnaZu95VDVQr8gJMJYiz4OM+8d9028
nlwF6N1cylV90pkZrdPt4QCRmRcanUjzxjdvmAeDrCD1ZIOJm72FkNfbGfQbfT3F
/gcW05O+Ww8tP1Z3BWPYF/ps5QA35moMsS9Vl2Ayn3Wtui1J1dsP0ol0Wr0411ru
WlLa9g1A/fN5d5KRoj2nHTEpo4Ueh4Rb1W3iOnMneqcrJvROJ2bm5lYAaMFMedRI
9qrhmYwY6l7T7zZCLvlC25WgIq626Vhn68y01gYnVz5FwBm5Y1lqWI+ynPClUT3o
subRf2g2duqgZa+Uzcnx4xrOyLr+j0zMcumgJHmyBvEtanmYu/FlY/8AepX8KjPa
8pIlGYyTCbjWSOzk7S0VAyEhWlYECItcZQutDnq9T+JWvh6ZXCaYhJhYWhFCqubu
tUnkN7tzld4qbYV503bRs0AM8mVsM3Nu7Y99Z6f72m99grPNrM4WMVc6D9Ity5tW
me5CXI86Aet8FFVZJIxVJsmtptJA2H+SaQWz7BX1h8eB8f6AiCcEhqovJjolnvFt
ZZnziURB3P7F/AtbFEqEPrivrrkRIUzebHEEsOdVtfJaPIjVFlq5pef3r60RRcP9
Urln9JNjxebHlDe4fhkApD4lidvciTav41qMGAmps1xsuRjr7UtxlJjGIVyvDzSG
yHj+DIhM5q5yCIAXOGHeAMa2DKTEnuXgS0h9Q6bl9jFZcdTfTrc2dYjFkn7DGd9o
NO2OQmDYwvQXYgiyl7hIZ4NE59SURNHeYyhzXwkwHbhiLw5H/6hzNK7WGBzGDkAS
nf9GyMuelM8iu0kFw4h4ZyK6Q4/v3hlFQZlTsEHyf3Pg3SMUkPWQMXrLcEmCKOt8
n2Tj3SJ09bk/pLWDB+y3aBAaYf9fFZfqd887yFLx64rPgASphOHl83VbM3VAxODc
jhHyZrCpNWX9gvPctyQ9yASCUJ65Dedxlv4kBNtJa0OAZ6S8RC9axrnqjopgU4UC
sWUA7umD2QHGZN/bQEuHd3nCfqJ58P4ZDIybehJiIP8LYFTJQoy9NqrxdputLNPu
wuxH8DGaVgvErntn67VAZUcT5R5Gohvct4cPHATxgwCbauZ0HTcIvVyn2Jt1uc+j
nLJmjr38zvZ0kNLhY2mCd6kY8LmR6x808rcCM/8254nvWBmVOtlr6bUDSilncwX3
93p6Gw+pOKAMcjaEy3FuH50DwTvant/sNNTmHVqMJ7VBlWJjrPPbSwvRb/NL4c4Q
UTzw5O3ChgPHJ8eu5BBItnkOKhyVUFGtOZhOwnsW5hVkLr3GS3vdcMFLtHlsWdce
5tMXvtN0wHD+ilwi12n6l27/+F/pU0p5yM0IjaUuPS0AaVAIDYyvTwStSZ+93nIU
4oG8IuMxxsHVARU9rnqk4zgR7SlGdDDFFA8P+Tpka6nzlti6YP5WuxY6QFxgTcZ1
iEtoq3bv/oHX2HGCHRYR0csvT0JVMovvjkH7ZwjjiS2F50+Jj3y6HZXRpUEsUVFf
bR1qYf20yI6UUsFdwXYTMojwzBa3MZzqXKz7Oh37EUDHd+nZTsZCkL6I5BjBy4RJ
bixEiKb8kzOVQjY3xzoWvg0hy5QVyXPXRKx9sbhWMRf7S+Rb3Kml9oZwhY0M/yfH
XAV46+o8tPKJhLoRMPkJp7ehULBRtMMzsVVymVmqZ1mZLHTop4ZpT1SQ6KfIa3SS
uy2v9lgE3d+lu6YlJcQPCGlFVcDpip7cieby50gjcwT5p0dPom3Y4BBmyMWmQwiF
hipinjRojAZ684PQiktnYxiDbhhE+EiCVPvgbN6QmsVLObS4Q5eFuwptXUGEEPNY
Df90FGzHq0xd2gLW7vybow/fgyrmsGzrhCkRD5PYS1/XJDvkNrzQLQBrTB9V32X2
XnUT7UvmOeWaYRhpobxCMGPPyc9hFKN7KUcD+pFut7DfEUsamBwdCHu8g7TkUrx9
sK5DRi6VGj/aeDjdrKU/VqGjCNiUOCtbs52pYAT+O9wrHFfcEEkQs9HDD7V/KN4C
mKnuFobPEaSHy83UQ92YWONwgB7H/MOVPJg+DW+gAcVaLUTg4vN43YTX4Ux/wOZE
+aHFiKoJ/6PDoESddpKy8vfyvMrkcn8aAOp1rCcjS1nGzmoMQjGKVuDSXDzA9JeQ
B8pynLYoJz3R1Ps/y4vD9JX1L6cPn3DwP6amhwLte5ceuhuIy6tTfhhl9tfjgENe
iACjjFT/h+oERpE5uACa3iTS8sKIYkjvNjhC2IXCl+uL0Bub+HyYBwZZyTT2HHJG
RdoNypZUXs2QoIoli1QLGBAl0MtgmwxfDxVEs5NNzjWD5eLOIHxQAQ4wlcP81qdr
nbKik4hlKqpxkPlaaQbLa+lnXp5j2LHcEBKXXgaRxIXQ6ulG/wXY0nxlhQeRlzhC
oFAKgszx9rNANjttdtQuz00vaTzHh9FxcaDeZksfNRDd4kN2M08oAubROKhNO/rc
FrRn+Vd5VSrXWPFxzaJqO1sOPIJxisOqFlZRs2Jq2oAjG7vPhTA9FivrRt3pd5H5
bCZOhrXB7zGIemf9ILFIeuAM6XxVDKDQ2uWNCZV9rO9uoQQDfo6/LECF7Xy5W4/S
DladABiMMBTjZopkXAFBOpIfzuwC5R92LM9X03zFHNiJINtGwP/+RFx8OYfzakmF
LOtN7Bt77q0Si5VleoYy2Cnitg2Yim9YKGCDmd8stsRcdnDVb7X01MwfpLi+RFjp
WpYow/JhpXzFioFHg7crsacYVxzABFHU42t8OXbV2zNwhdBexjz/DFO1pjjOxmbQ
K/bXWguzJCMtu7CRFX7NcZDOV1iUMZWC1+KUQ00e3Mon0XqZ74aDnuZS6RcDHvhY
SSSW1bVt2L2XC+smELNCUqnH90sphJ7EC/Yi6XZ0tJBVo3s4DC5sCfmg0M/qBIlR
6kRhO2GjDNzi2vksQ3RpcPc8+TA0gNJQ5i2eB0CJnR3dyKOytA+dZqwstV+hojrE
7CI2vPf6ShwVkF1ajvLVM3q9nK0wmlRo3Yvp5Oud3t6RufH5Nadc19Nge32u//nT
v8e4+maRUJP049pI3k42bm4+19a7vzaUaJa7xgAqDN563grqxJbKyY/mAr1xnKDo
2mplteRO8u2iyaJVY1AsJXopM8J3HwHCkxPr2+DpZjC9AR5IXbeGvAxDBZ8ftn9a
VcRnQCA9h5H2HYvFSKYJyfkozbb0z3T/vgFl7fL2v298t6JUjKlnwoUuqOmX+4ZQ
w887BaPrNRfdfw0ZL9pl5kY3Rw5uBdC4r+fgArwxnRDT+hgHeET81ybd43C9Tadk
/i2G6aCSURwF1nI9px5N8gm/f3pU3Kx73QtdZSHanbrfD+vSL9A1bbk+tKzHpmUT
8Elf+HVvVxe1hnUDtvwTmsHGlt3Uxhx8Bva/Xm7ou5mH052ljT8CninH6VgMDQJw
rxqlmA0W5dd+B5ZtRfSIWVnBLsNByOQKPxLUSMCohDy895/+dCg4Rlvh/rzzRDp0
lGDkr3vUXR6tuvRXRKuvPW8NikWtNmfjjRHkeucmOfpP3IU9rwEf5Kon8ShgQ+2v
fvyslZhv+4lKHeITTXLoHHDcY6uPfAdrL4i9/q5jXa63p84v4ntZ8TPoTBML9zym
U2HRbibVKmdyKv/Bj5/2RswsUa4ccZn+tsDFxkF4LyWvF+9oSFvcvhMc7HlK3Rln
xXICtG0V3pRy/eyMeyXIlIZKi5Kut6BTtFLLrb2ePN126Z84sZppwO0zG4HWjR83
f+IYtY2FxEV6TipAdVDho1866LKMc/FEzbrEMyBtDRyw+P3i6T2FzC8H4AAaBwGK
hnEL5xscdoYqFbQUROi1VUn6PBQwx0HGeTEM6n5DhJy+Gy23vrvLv7/G4Ogi0fLT
2dvKl9YdggX9SXRN/vOhv/+yjQ2QTGvuTKfoRZR8xLX/7CxQAELH4P/v8bfz0QiF
wpiz2zaHS+wWKjIM0WI9TrUsbbTIDdk8IapXiibrDSaXSiw1ZZX+un8A4Ih5FuqH
LCP55LHKUe6mnVOuUzkMBfe1ZBoZW2BZrQ/PCA2/PNakofUoLppkvd4zMeXMqsbf
pemaAe3iXzoCsxxY7BxMionXxmEEG/BWRKsSuWS5lJ8xxZRSl22sXmHmIgZUcumo
HuqqBi0puNdqX9KSbFHt8XW6hr1KS4VBbLprGAqejRPuxdKuz2RtVomlp/PHJr/e
3FNzKC4nT6snyJG6LHAa6HOIKN0JzOopfbl9zVprJnkEDEyjLVf04wItjSTW72pQ
nWCE499gxk1c4pXxr0qNOmppks6Cnx8DrVcKSIizEPWRU3rdUv0ZPkhe5oKfF1xE
wBiQkclAT+G7gkHnDL0tSBStIKFT54ot66dO1jkh1xxMGTi0BmKWPaTjRTwDPW0j
yJS7ae1DkpfO5H95WTrvofWVAeHdanSvTcEwm+E7E1AkubSq4Pn6/xG4DUPyGjgJ
xzd05O/J0CaUFHUDYN7cZt7Fz7tSNu/6NVUXLZ9XQPj0+YxAl4KQYOcOGpRfPrAt
2cD959SD0EuPWMf7g0RT2bkW/uYKAuMTEI58ycj8/bwL8oltuDN7q7WTTipGF6C4
Ivvry6/s4W7V+GG+Nx40Mb3DD0C6z6Ch0HI/IczCDq78/qBqi0njUmnM0btw4lU4
TzXf885HhY1QT0R76LravFLQFmkjdfHNHO2o3mntVumldcimsKnx9ijxTZFmPPEK
hKQtMBhRFHejfOLqdXpYldI4hRsClbOdI2iRO9f1y5dD/g6nOZgMV/3iiNowMMZZ
wELDkYHv/0wrCwKcS3zM7rim9N90aFVD+pxyoGGPVh6Y+kX1eo5oU8V2HPBnoWA3
Va6BLeQRYJs808GPLgHg5L5/aujkgbdiWMjNhyFXKXZ/tDt7Sh3AZEqvgF/Qtf/u
78kXjgWpANIc9MCqZqGyzPBoz8TBrsWP7pfXReaxIYn7rNw1u5La2IxjWmG2l6s6
LWJr5/hhvJRx8KOQ2q87VGRhkAVXxsVm3yL9OHltbLD/w70GrBXfqtXXf5gHiXJ+
mHOQusn3xIilIxfBn+83XpM9KwW/izNR2EERjF3N0SQZ+sGPkdUlU+eW/oVPmHVN
u98i9WUZfidwkoMSnD/JPGHNkhTTNhHmlHHcY8WVpA//Vij1Il6d61z1CJ3anJP3
Kswy+VJEB4EmTawic05Dl5t//hkoVmAU0Mol3OtDPhfstIi2UztAjUfkcepDOeTk
AhnKslHdm3DNwpD9mO8yo7bw++RUc9DkXDpw0XrVMnWSCS+k4CyNqCTbIOCrrTCE
3fG+k5mU4PRu/JJwTtyYhfye3HhpHgypLMebh593ojP9eVONDfhXWJNpWHx88ofy
k/V+0sM/f+QEw64F3Irg3o6AXOH7LvxMA5vCNwC5aMLDHtaEcXgzDKSAn7DiK6V5
hWnA4BC31CoImxfQY1OQIqzsjTr7a9Fy15aTX1VXhJLLb4pjYkvhWpEjHCcqMaoI
vbuboT3qCvfo5nT7tu/N2gQKHHkV9wTtjR8ZLhmgDKgvS/NGj9ioviRx96cK2Nhn
wk6XUS5wpQJulnDYLWK0P6q3t/QglI95fgT2rpoaahgIuZdCuU4rpqCyvR//G8er
XnrlZk+NKHsm2qhZuBKc5Cqw5c5rQEpWELlyHQbgDFKcpzGbMpWZx+Gy0pcgmSue
7CRnuqVKscXxI2ZwrtLGN1zYrYlL5Oxe1T5C4qJtFUVRDmk4sdG7IAptBOeN3pUf
Ln+tW3wVttzsEsrgcEX+G9rXHURJTJI9hKQ8FBSynAswh/0lUpM5XgDJN+xxC1BX
HMEAluoihZGWpaGIep4v4DiGDVqz6Iiq5nmva7fRT4irkpA2yTXHW+ddHHMv0CSg
A/KKo8wUhR49IB4lZLzBEHL9YT/ylBk2CaSR09WBmsWsO5OWlb1O/P0pqOKmNJLL
cAJ3Lb+17K5YxJkpfek7QuPhx08TCsgYA4qCQS8F8GNCnuonFOQg1OaEeCXnK5nO
gDzJj/njBW32gWKYKJfYGTJyKeIIC5m+6Jmbh/387ZLNS2+5kcT7O2IM//3yZg4T
sq85ZJlTLkvd4/VFp/zMKfTw9ZeEckv8Rp8ftsIyKTzH3LUxHkTeM9CvpqRp3h4O
8SALbYM65F+GpgQOSbKbZVNSFJcwFhoE6w+41SwB8oqxFBFk20Jacenj7ApLqTjT
S92NhhNm1aFXetUthnQU2JU6FEf7K4ZXQYL5wEFrF/Cd0BqlfutOS2OwgvvMjyI0
1rxdyj5XYgH3Ur3o6gNIJwHYRdMLIgLw3frankrU/fHxV6HqHuzDVOYguSpJd/hs
EMRTERnuY2zWLpWCNBDRF4wI4pGKeb4ndZiQQNT25GxYcK5zlwcJ4fh4yVPbAuU0
MCGvxoLclW6AFrZXIG4Lk8FbeIgBWvsY3EGOWMetTyvPZqPT+Yf2hZmdyP0N9ZHP
s/6+bRRyXrFr0QF+6c12Iqc3z+eGs7ZxQA9yQh/nkL/1AgaU9Thq6WApqWRy64Wa
rALd/CH09h0FdiSJb8eQfueQxdP86Rsr8k3qGHQWzva8aBsHE9C2qGwgIW1G3WFJ
TkZAsweNJ0usCjtVygqjvEi7Nw4MMqMrhQbkf7+ITTcGW6KmnqJJAfxU7B7PKmgu
YZuBOp/D8lFp0xsB+UYkkmBUdpxSdnhh3V+cGgjodtuac+qF/VK9Edd1RgeMicUR
OVfJucvJj3gvgQkZt23cWvvo0uvyo0vnsiqMNBUjG6taxh7Uw+7+oSX81H7rqrKV
vznMsGqe0+Mdng9k8ItZMjql+0J3GA4LhLjFAzhBkbRAD85h46AxhNcBghVlZVJi
0a4WEFhDq8UkYK2EzVwWNlsYpmzvXEB77iW46x4L+r/eIXpYxa1dyZEjx+n0Sl5e
10ipxI/eOmL04Gf0PFQerVuj6f7qsBEYnqW+X1O3GWlVFVEiGDl/y0CecRbNvWfx
/fcEppH71LA0vjKSFFnDItMwCDmgIDd2ZgMHYL+zdR9DFyD6nSCaMsEc7lhLQJWH
T0/AzmsJKnfrieoZqdCivgyvBAtz72dLA2SqsJSGKqG/tVa+u/hmxr7oKcAozuJj
pxwCkSo8vJhap4qHrtoemuWbnfO/jcF50pSk1APwVrLb++4g3e0J7dFBoZOvwcNo
Lu0VpoCm70UgGgsVlM5chwzZrX4rzy8NKd+3QRx9cjvXKYE48/+9apRka1LPrgD7
mbobEf/hRlKgO0HvAvvyiQS2TOAaxM5i+B0R8qrgb5QyZVbufTNG4XeqinGN1+B6
H7aRevBDKAgyW4fuEiYF/u3S+L8HuL8NIqXNmYvaSlcrPl3Gp2rbeB2xUUgAkEn3
uE5yrULSYOnTsv/2wDU91XcNijnl9dLmb6nnrgX08mN++UtoMYT6a7w+F5m3xYD7
9jzTShx6FRFOzSNT5I4Q0TypvNl/mdi4ioMBhCQ5AF9pyk5cLU/ZV1bH48SxDY3d
DaEV3tvo4bulduUiUQ2JhPVC2jmm537D/aVFfxFxItfJQhYJUGZ+Sm9kvBjRKg45
l6BUjXgRVdmYFcplEPWuYAdbUMjfmfn6U/cenh45yMG3Uq0HY6iNJ1+LI6pQ4KzB
RUJpln57wb2Q4ORHhmw2nXKzbW62FioicadOFvOQap8j3oKsD4kH5Ak8s3/23Tw1
7NLCC0QXrzPeTLJrawZU1YK4+xpL9qWAgmCR66+G5wCdrKLe5GAx4/9KoczqOpqH
6H90SK26AojDttiF5attz/Vi7RLGBcp7zwFLt82Q8LNwTsM0aIr/IZT2zXAacSDx
xYR6mFEnty/HAnpCPecNrl5ooCYU/Z1x2g6DrKgp0rFS8ND5ZsArZSxibxfD2uxE
toDTepg5lcLzaVOH62V2onaCv+fw/f+kWaaOjCQnjT9n16oZOWrJxF/+LrYo7qTI
NkBuga2GY3zszSrE0aBYjiyQ+6QwzV3tsIvgrW0V92ysXqXkwdqI1EnnNiCvSCd7
9tMM4op/QWQLCvLNth3JJcramA4eXINeJNKcCkdViLxbEyx4UZSwMwLMGrlqgIYt
HBLYYhUbE4suaJBa0K/wi6SNcSFXtjrgTUn5u1ki2Q6cnSgbDnFXCRES7nTPC7Yc
VAMQfiq4g8YdjTE9ZgA68dJfItFSmBvfCkf7LtNTfl1SbfFwrtNxL2QRumHGjCgX
MPVSIealuBT/8TUqYBvvjTHT7jKRhCO21kBZLaw1GeMImePxJCKAqWVNmRsNWL79
9u+KsSh+qiapKRUk1S6A27XwzYEwuKByM5nwFdoYJryrYg3C5onhUA2HFdFy0C26
oYfL/QQfvbMsH7eTvxvXz3zE4Nll/DIozWCJ5gmNvIpTPA86249+5XBYzfQdoPlI
iDuTLfdtp2egpkClHmYqn25seg6QU+Do0VUz8F6IbF0O132wrB/4P5QNFPjHgBRG
HCfkmPboQ5KRzwrpr0nNsqtyA9TnsxRK7sWJ0IXveedbTX0IbzKD81OgE7YZRe1N
i6tbKZncW3pOphaRRyEdoaix7+flXJW1pREbOfTokQ4MTQi5Yk1QE6dYvwIbKNm8
BDd1Ed6I+GvWlaksfBPzOndHarJgI8m5y+NHVF2tMOVLd9bnknne0eie2+iGB5RX
jQn5sdlugOLO1mLeZAhgp/ypfzbIUxPliPvdDt6aSKnmBXg/q+4Uxc4oLeej2IQ3
b5SxJ3Ul3Ndja0yER7cmzaJv/cHldu0ePeXGq0NH7FYJWBILlSFaBc7iSBLWJClh
pKnsbMmQAz6secYZ0Q7UEZmwBYJ++Q7OjjV/lAG3YQ+D6XEh+VjDguy469owIGVS
ZOW1k0zK8M3coMFFLrE1ijQkOx3180M+oL5Rpjjj5gRW+JHZ7HmBY88c3VsP9bhT
9xQshnQTGLXhgV+4KUVb+KTjkFVp+QmCJ/8SNIQmwZJlEXT/esxe4LsCW0RNd+V6
L6uWpqhDETAIyxtDhycSbZSn9SIMFegudKuWmw5ODQRTKfRZleR4wZVts6Dk3Hri
nBH2LHNj345AdYhHBQ7rM2ruhVBuwi7H9VcBBEWzWJYiyGEg2O+1LT6vTd7uhi/P
klIkDhtyigSSrBqwlLADPAGKsIP/qr8hT/3d2PE8V44tY9jvDFLW2VDJdloa7/oF
oynVYclKmH/poetN+Vad6fU9ZO3TCHdjrGvi8MsFUuqdNXvIJZ+rXk4JEr1jieSY
Ui8z0EL4tK8zNa4sOtbMjLA8FBJZ4zwabUO5CVuiKs0W/nmKzIEIkke2YpyceR2M
p2sAzrvvV5FTHFdcxywnOckPfesmavIgJFz1v6Qsg8HSlrTCW1DRH6WfQ15ye4w6
r5pr2vdbWUDWvvJWskTBBgCKmOtoaD2rcZuqHUKjapo9s9Oe4p8m54pIN632nXQP
VQkQ2nJ0QwSfB1BIiOlwAkALv7bqgUIfZ0CqP4EYxA05Ll4PYjOBO+8/jW6hMYZ7
LP2eJPpTzvq/9xTIZapIMbwZWzgm9b111D4eQ7ob98FuoXTvT4BD9E/E5PAwwtMa
j+dSo4j43JyGDqq3prZ2VH9BtmXB6aPcC3DD7wAYT0aY+SzegAltv4aLDcmgv2j1
VmFjFl47XtTBOlnyeo7CAH8W8UYrNoer1svYhzTy6mHTJN3eWTtU4mVey3DcMmtH
1TzG26WPBob1L6JFBCiTvgWleQ8/KQk17vFP7xHewXy2N3pkKlgaPtY3iS8nt+G/
vSsjS/ZACcd/top0NY/PQecX0PG1ANmrTQYiQXNMurI/jGPTEiTDMbKmQZSW2M7c
6O/WQq+frvEK4Ku9ELT3KIAnXEQ10UcEgI6boKPv3873PyzEC8tDdJNAkEVLMPb/
PTeMQYGFk1IULKKL8YOcCGpLvVilJWuxKt7rmpZ6t7pOuETHOf750irP4pdi4afB
vRpHXTYVQK33QXY8aSAQhZwipTHDrQYZSEv7OyNNzqg2i6iszPsMyh5WnbpX7JYm
fiIohdxESVkKZXzL1be+UxwrZQhFOj4HQ2HyGOGBucVjGsBonJYttGEkXgLgjY+q
yAar8JgHNHA4bi8dfDjWPrz/Hfrah5n+Gvjlvny2G1q1SJ4ujYYvbqZiJiPKPeT4
qHWWtuOcrYKiTktb3rV/idy+hN4Y58OmlKVAO4TjK3nFPz404lOhMGHM4MKMC2i4
qvEb66ouBDGa402hCZP7bQt5UK+o/Fj4JpRcCOOf6HEwSPv0/kR3MigN/YFs6OE9
FzMaYtopLkmw+bdiZwM8iGEAmbmRtNhjjlwoZ17TTQNkfKG4UM/Z8myk6bP9JmZA
wLjOrT7EL0MkKT6xPSep2uPKge4zWgcwN+TIQ7N/wLymNyOX8WZtb2czMMmJnUgK
hrQfQB/qCpx+QuNM+9upj/Mpv4d4S8PknXzZph9umJ7YPCT+uS/JSRFoucPnk0Sm
6uLfh2godcNslrgfFmF0bW8bLg0L2DhcfiSUBFfWHcV109My5FhPNP60Qjqg5UC/
+mPY/gQQ/mnPyXAVZ7YvnknZ+cQWXzpqxORX2En8+734FWo8HtL2vTHyb1Vccdra
8wk55RMrUqDfsoqhMP7J9d98PGwb+odEBxuDoG8E3KHvDxwpw8m60LJiA0Aumu7e
oc4HBsYjyFQVH77ROrI7HIc7pIPRp/Vl4Gp/O8JvJbOkUyF9ntXkeBIrIPIOdWPs
XJFk/Ib15Wl/XYQ0cHEabLxCKNiFAFlSj+6mwf4s37+gF7zihdc9h1Ld2GOMr2QK
9Wt3UvbaLzbRqfXQJww35BtXNvvLWKd4CryRUVAcrb4e4kzumsw/tKLIPsMR0w8N
9gMr13L0pHIpfviUw41T+ZAxSyLTDwiw7QJCi5wFhjiBu/Alf0hEC4I59XDOmrNi
J9F6l5H1IiQy9/NA/SV6qzTAJDG3c4qGF68xcKUj4Io85Q1imp8xSG1LRCcnSfTT
7sF9fkP0+S1/kVxKlCRuCd5xhO7FKM3Vy07xxwtlSZNKaJ8GuZIdk43p0S5jCJ1x
C7Qbxb+FCltRO1PFotizoun0SM29QZJLy7+ISqp82c7Ot/y0n+vsV504sBjbCGc+
nhsjm+njpwcLUvJqJtRsUwTwHp+Hx7CjLknyyUhUOqGdR5IoJJIhxODCKflTZ6wJ
3dr9RDUJfKQ0NMgaisLQLsLUGHBaYgsl26XcIKg8qx9HV/gLUB/UQBKIpOixDqHo
Y3BGi+HnEYTiXT7a0a3WnJAO+oXBiM5eEaxFMyh6OVVIiJxEq/VJEuVW7jN/F++L
9I4Zpmbdt1sKflUCoBiIWrlBUCt4P4c1itNdL7lH1B+S1QBjfgUL7N6IFV5JNYuo
UJAYBoQxNeEHhne2EeqTLwgy+pLz2Uq/AFoMsp9bV87JXEIEn8yPL9k1Y37IslBy
RzeS4XLICIIFYzrCQiL00EusADD6jTetKiHm9baMkA9Gd0b2pq+b+Jr06ocvn9ud
wLroRkDaWFhk2fW+iJYDuX//yB1ibMCAVhlGXkuvOpfnZzbaZ/MsvfD6a9C2ZKBD
eHPoDDesydJUJ1jNj/ma9uXOG3i6PH6/M9c3p8cWbEncRb8BVaBoAgOUDiVpdCR1
CLKtTgh+luiDVQcS9zhrPg66jman++KRLgDFFc9KOKcnSo0I0n43S7pTxRwx6FPM
iJU9yvITeT6fo5NOKlPLDAjNJACW1p+GWLYypbjRmlZ4/bBgHDN/8kwT5G/vg5LF
awlE+gAu3pIxbEBf0QgAaw7aB+X9pkhXQUx9Ylft7oTVKOFfuJ5GWQodLdfA9I/w
D0JB9OT/k21zvBXpnBs+oLsv/BvWniAmyhUXy0Jc66VcfEmBVfNpzMeHe3tXx4l7
mfBzb1cT4b1tZprrwPeQoPkyfFPixjeT0zuHxrp+S/ZSzmw8z2R8RnN4cRWiQjRB
jR7UzNwJt0qiiTse1QcZV/Du5Wg6nr+B8CAttgXX3wDdgsPJ/X2JBu4a2uV+tVBt
X0QDqad2Tu7Dpcg2HmDmmOxK5AbZr4VRXgzYOxLR1Y0QoQczOzP2nZkjEa+3Q5fa
vyfQv51BWZ2LrVaN9kXEzHhVpPQ5Z5Bh5mJ11C3D0Mf/r+qItleNi24X6hJtwfUS
B1cupxZSFjFHv6H8DpTU3jaR+aPA/wDjxDF/TSVLiuqUDzPDmZ8xioNgm4AKnawF
nB+iBCAdWpbCXf/2dYCA0st5uJnMkRWEgwIDBbpg5jbycH430pMUKuMYJLctgcZS
VgFC/UJ0rYUnUAHlyao5RC7kGGTdBntFkxcMtY3CC1LcGG/SrrQEH7BJuZf6oVNt
0y/SnCrZuItQcgSX5J+6HS2cou6X/vJlr9Jixl542/orKP1PT4SsV/+68Zm3rLwE
okmNddDgp0g61m2a+FIbM5msd1HI5peWo97UxC9UgIaeCx0ysnzVEvTxEW4j+KJv
0cdBYTBPIglCDzJ2oT5pzG87DV0ykFu4vxTK8lFK7ubH9Hu5TkjZQkx2cdNDJOQL
CABY8XUhyjsIl5cwVQG1QY5ON7/ASH7wneqlE1all/ut3q5o2W2ADNqGceP6WOoC
CGfTs2eKCqnIj1wyE9jdglht2JkcwkNYpP5VbkPtO3Y0jzwYZY4gUdsEx1XtyPKt
jcDEviWrFWtfl9X3o1teV6FaVY3TLH2obZrQyi/MaZKyRiai+Qnup3ojZG8tpM5C
/ThGLIJdCR/Jdm6OESXnQxPDzhL3tO3/qk8hxbOtayOGG17OX4VBnNqdyaoKlf/O
kKMA0fcs4Qsn7j49bkWaYGb8isdpeuovAxDG2TVpR0K5IOndPb4jp6X2Ded/FAZD
lwilnBRuVYHqgKRJWcIAbTDc+eJQo08Rsp7BsNOoWZ+JHc4CduDsQHthTe4MTBDO
ql7JfCg+IyUSK9dX+tMHQ2lY3lr5bfTVV9lh2fjmcfnpPmWK08s8t0rcrDO+DaUz
vLiEh8JQFCdKYsMagHnYVzUC639eCwoFfeEp8izMRP1l8pHk4Ab1eh+wJuncqvLa
TXn1w0x24N3RCN4TbRzjbBLoPjier8QD/KKwh3RVYpAtwv1Q8FWsMyLXUozF2YDO
cNZOoUhLiRvg/SCbOgRKvyRHA81BL2seRT3aB6Dcb3VANkpIS+iaqCEva7wwxaXE
Lfc5V5ChoqxIzsM0uBn4HeTcv478OwHDbqtU9cSzlWelRsUTFfm+wZmtgQAmomMs
mHX8CJVbyBCIPEJySwwmwXR21PYp2xfKm3oU4B/VhQW6GUwC+ruhePzunRPF+PLN
FFjrD2NrGMCOnHkEgaa4e3q/emyglQEh+TbKJDNMFIvqxtWQVmeo0tsP625arRkt
Rw3GucuGaxvh/mtQg7/9GvzTOOK/BiQSQpvYVRf3LCOeecAPgBT3ZixK9oQlhyB7
Cip64aDpGxXdQHqyb7YvY9FOsPxcNJG/6e0zmszCNWdnZOQ8XfhdurrM+FdlmjGX
7vH6W271lnmw+8VIhyLyaimu5wCH7Oo/RAFg9fDx468EKBHIa1mC+1tjywi8df/m
SBzoVZsd2jhbzCB9qcmNiGVP/taxUHYm7V7368Ve/jEd7Rkcc8qkD2r5GkkjNv/D
81XPeBY3dcJSRJbsizcm4pwi/FLw4JxYkJL0ATcgJuMRhp6K4pmJPrjEL41Ei27J
FnYmKgvyTc6hjDJMztgdTWZOIhzyE158ilJtR3Vq2ImckRWUIRVi6rsoAByTxaBc
wEIjvXFmiFc2O++EAZ5BJleRbSo83v7oMGIfKIYCHAzbXBDqPtqcUhPSumwdhlOI
xkaZXlXyZzDeh2AHH6gQtxa2aLtJ6sCu2kPb6y/XCSJUV5s4ON8uLOBT0SQXVYmo
gvadnIteN7uOD79TAMm0sZOlSifKmJI3AC4+a9tGrJg8HlEoK1Ge3Eb3AgSifVjn
dg1hfTB4avjXtFyW+3+ofV9LbTx79oj2yu/59jSLs96ZFdYZEdJdd6CXgoUECMjM
xXH0AOFyqLnaGLAV44V4ZOf/F1WYGKe8iYkI9ycthoRx5oDZfFj5IiqOtlSclL5u
gtHE0nEkN3Czo38kmbexwEQYAuJmW39xsTSE44kA1B/aCQh9wa0pGQ6AFrJ3xhId
+shNcwi3GHFF5N4apUaGcPIWgfpcadmvKUwHunEWOQlfqszMtNcP1f+giPC4bx1J
oQ2KHI/g1olOrj3WL+FsUUgTbXXiDVAWWoE1qI8/vVpitCCkjtsnO0SA+CbpJ4RL
WWJ/FHkzkM3OAvaozZRyMiK7pddgpiOQBsg1iKvScbDdQW5OGtwE1YXJGAy5BcQD
UajaCeYXMxM47G5fLrbd2JaBvzmhw+EfhTFzjyN5S/SrVTEWgOtnO955Jko7EdQm
Hlff/t+OrAcz+dEQ3FhNszLy8uwGKfshnedFRv9uuRHQNIYf/vnRDoBFdMZWfHwM
pPf6DOV7Wa5lyyML0APhiFrIhHQLdEMtsb0by36Gk/EIUxKD0C7bdodcTw9dKfO1
SO55qBB4id0lvvpilej8Nd+N8qxZw98FIcmjeWprJizaJQa0AtBYuT/dvlUeGT6E
f3tlddCffK58vpFvL3ywqF1ImKsmEwrq1OdFpzfsX7SGQ2HoSQ6FHk0VidBms35E
foBaxBbgZpyZinM46wiwMsoe8RFTrDbVToncKlX7lIiqHmvCWaZnMVQgOgdTacsq
DfqVzxk2EZnpTpg3uy/nndF/kF0rbaHaMmjzMwtmYuSuZpFeh0/0kpexAqpHne86
YUzM0GpmdvtFpYyumQjE5odF/Nr1XuAW+3Nw5PQmF59LdI+/XKcG/Tvkn/jejyUZ
jOEFFrFUI81CI8Ff1voTwCWhppa7BrfGXDGHu0lehGRtafaUJwJOHbZkOulO74On
Y93lcv4PF5VipUWuywnIst7Be/stPY3zu/JVWLCBmVItosg2fbLyuSid2Jpv1onh
HOjaHXx5nEXYjAA48buS/nPnuGVF7KYErfBz1ggE5UOeUs2FxUBo52XCb7f3JqzO
oaXhDWP1l9wndwdjhwZmatBfJtmITc/V9Fv+eDFGE5Ge6L2HUVJ925OA1IVOa0yC
2eBYpFfiSQoZWo0GdiG1gCQmxf8sGkzOMv24Nk7C734EPBLcH8+qAv3L9LKiuRBg
5mgRH0sv1a6qt4QlXt9BBxH42IfD9kiX7Ay8wrAksvARkW7BDd2sy7pRM6J3x2Ek
BqHZmG6A50HJRXLJ8ISI808qhY5635FCjfnh55gTRbeFQE3h3Q1rx7yf+vvcaRZR
8zDVgoQJP8jOBYM1zFEeVYmA9yb7lvZsOTUNnm2yqGpfUOvkAY+KcHTsp1xoFDDb
xgDGOPgzBIC0jQ0if9JbA9Zl9K0hCB4kynWVeBELDI/xzxdUJIqC0hcpoZKHb0OD
VrA8SmUlU3ep5ti2W+J3CqbVT2N1H9P6mCacztrvD/9P6IoM0qYf0CslkgxF4AD7
o6gH035DotySLXQqR/z1GM2Y7N+c/ycNxeM4uTAQm9VXwtOCD9NY/HAAhYZ1nwn1
qVRV3ngF8BvMgK7sXR9WhHH9/q+9QyM13S+VIwTLcEufiD0/LHwHhnv+KH2cheN3
W58siJO6RQg8gpJSxtzB406lSLO46PM8IOR90w4EwPtmCstgz4TwrqipFQIvPx7y
Y7BCFuCmspNC+F4S54nrO9h6VG1BVlpbfFJPN2rkRMwAySPT9TrBJiBrXC0NDySD
Rf5xTPcP2iRif+F3alQEIlz2hBpxSQSQLiYDDkRO1lTkuxiEeLhAh4TrL0S3w4ae
6131nvOnm2t/L2Hikds2ks3pqIq3F3X2viBiDG65z9TvLIQVxNbi7jeCtdn1wxIp
804DXM2vjj2NPejdHaHfMDmWwaPntjuAVAZugMOLVV8T3QuciwymLgtiLaua5fMj
RhHmghANCx8DYY8a/zoeDnCet1dSdBJET2NWPYe9l3yrKG2Cbm9vwFdiXk6iJPJ9
r198jKppKQDqxjocDfes78dHUGGXR4mnxsKwc8cl4TrwXXsRNZlAqklQi1KLrycO
YDEc1RmSL6hx9A/ry6GTvWnRC7QmCfdYunh+WUgqzBgflby8ZtGiRMYc55CjSPWi
YLCZEJZLSg18DIAPyY9vsS9/E+KQmIxTtlpNRaOLl7/qF7RiZLoF8eIHGMVP0esJ
/XcFKK79Mz5wYNt3QRNeLkJJc5ql7p59NTwHLOTtb+kUkdMdvjYia7kXhYptJIy9
yH/UIt0r3DpMM6CQnXfcRz2pS6BPeKaNLfoB4M82uqlzpwMAT/zsByB7XsDmJpiO
KcAkJXb7ilA3rMEjx+Lub2tl1GPYJ74M0SQdVJpmwZyL00gipx70Lwrwn7HEsuic
DddDbNa2CLdTWyG808x9QADL3v43yGvzXMIQox6njClFt9qA5wRw/dLMyZanWFmb
liHMvX4i0DVyCoWP+e4TASJPSMxi8bU3qJgQgRJ1I2M/+OsLp8MOrFYnFIxdX6HW
oMP9y0O6t/EvTM945YR8QkMzPBd6kp8uz4MqQynI67yOMPZbORRgwo2IRMy0kvu4
mWQViE+HJnFjxMFEbU4VEnvEQQNqVPQ6d0F62a+n+EXOcNB9kfF/uLJVBRcPwDeq
3YTOLSDgnDgO6Pb+cmWuJMRkpf3GpFR6mSMJcA9i7llzuVTPyoNIzMhnTk6I6pSE
C9YAaJj+apOOe3llwnuBuiaSRl4WaDpi98PDHWjQfhUaIKZ3J/Jiv0oj9mfZwNQc
SWhJtVsjBelFng9aKlqlR94i+n+Olw2JVGsiZdoYRTbyvo4X2mAdHCkOHjV3uSIx
ywuHmH9LptO1NWl8IYY2oL4iAjscaNu7smQPBulANRiVFY3Q8MQmMkHwgGu8dgk0
eLgmAC2n6zZSb4zB0EjCiJhbd0IEC1KUdsVWhz53M/uvQSfpex3uGs1Tik4y9eI+
Fs/Uh8BxHy2dPJMGeJN9Hme3W4chsra7uoD1mhWM93zUGmvmTQGycefo1qhEKs1t
RiLU8AJHTJ0m/ZFd8EAy1YJm8mPjljIiHiGLQFxYEd1UTKFU5Xs0ShcQxZD5S6JQ
008o2GM63pXmBjTdxPc9k6elbFwqI0euLs3StwwyrU/OfGVlR87TyU5sQr5QSMYs
5JLkjDLOsr1GRNLnvVhnwFlIdRzCsgWxmJokn48xdIWvd11LRBlapr3Y5zrP2SIk
3QSdkhyQs1iyte3VQ/gwkoT9tEENyJjsc2snch//3/tFTL4++LUGcEqVzRx7+AzP
QPtSvh9ZRf2rHuMaIzf5DBqZ3LOScFykocoxV7uFdy0hs1ijis92f2fei1L/0Im5
Qtb4lzXX4Ex/GOTlri+683bJo+nZHn0uUBwuKMaC0MzujkDxwWVd1O7qJXIuevh6
DPrLVWqQTUBhEcIbCacMzH0ECnBe0SKwRh1FZwndL2EKAfyCQQA19aoJnWPJ7uOr
jBQpICHanukMWwIny0eUOIEo62i99gCX1aBfatPlw5xkz2MY6pYroObN7JNUhjLE
Zjnjg0NmnkWNmcvoVvoTOMN729O10TuEXDMOF/zqEK6vCHSOB/VYGS/xWuZDUlHw
WpUUFABzajCcxnTkQ5EYyE4yrOU29rqC9vbjJ68pAFb45J94nR29VBt4xlYc2LAk
dNr9AZrf81m2Ou44DJos14tqWqk+uf2bkQ1f0JLxFMPO+YkmqtAcXcYC3QFDrbQC
VkQ+cOf4f0jxLeXWxgRcE7sMdxZbnlH21HqqpmE61mPMbRTUC61IRRa34e72r3sK
o8lHYQdlBvGe1HekCIJ0Lr+bAVyMfKeThPW0eUmYp7N9chLSlAZM1SZJodlEpcbI
Yl/EIdshBBDpUIPCoYNLVErMKEpdl19OI20d8JjgSt30oDb2xROV9hknzARH34So
PBd1En14zDrLPSqddu5CdYvitdzs0/CG5F4zBRDsmW64kwJpi6NTqhS1PtVBuHBt
U9w+htfmGasYDrcaBwgCEPks7iG1QRy6pVk45Nzhr2Ig708pVeBee5aFCrq6dB0w
KEhObFjTeRdgpnKB48+xIeSwP2tShcCPF8S+KCswFCQ738TlMkJ1W7yuBq6i/aTW
znGxzr1Qz79SbqIvtGbgT/Kl9fuJrGR2mZOwpgecva+T9FO0NFKMXCfcDvU9Bdiv
FMjDt3i0+h/ZfJisZpLxY/o9bv3TH4tutgJbZ0kl4qIEN16/mtGOfhxThfNdhrO5
VLnNntqDud8X1c2S5QtjLsDjg8Z2G2IpHRsncM3yXhez2SEA5U2b30uSwR085keH
zZoF3/HukLoDDTzPaUUlY4268lvIHrz+lzIFg/+jwBpuemZOzS0/OOrxUovtMWyz
XoEVwOXbf+CTBuxvxunFHaRWxq7Cbh2QvGPxeQVNKYhgdS1V+BB8Dv56cZJH8Rd0
ynYKwDnCtEeGsi5Ia7/8Th5Pg6I1vlPyg6v9O9l9RqFh+4OIPofUKcoQMsXvdPeB
GldbSclyVfgWCnKmLtwL0UZ4TtNs1vth/nseRMdhKQWLbm3eCxi3sZLyqSrhLuXF
ZiQgTgyZ7j1G2TjXY2//j/pugUQxdSApkjiXITfHUycSTL+oDxWCLLxoa9vQ0Y00
LsJd7CoJ4Gw5FEHM1ybmhqd6YnxhDzYPvZwnSNsImGhs+j3UoEqBdsyuU08t9fvE
Fr5TnohHrdIn+aL0FGqSDrf+v/8v3YCxxg1IAKvaCdYRqkqMD1PWbBLT4y/hqFu6
oqLYB+00nQdpULgdtjs5KLeSNUNKfm9E63SsYhxdDTWxAyhj19VlfTzQruQJMAUL
mlDfrbhyKp5M6Z8TbvDeKa9N9wIxABpQkCWY5o8CA+jAhaCBmhuJaCVpr4dO9ndB
6v97thfwCWDBbNeGso/7nPipfxhoPYQGXRHY/7+hIL4sVz4D4qAhAGdr0N1RhVgu
lMjBQJH7t+oTuBzNGlmsj9kN81kU8UDaDMWwKRRxe6vJza5Txo/LMMYop2RQ7RgL
yl028SF/yvl0pBYx25anEGUV+GmdQJ/9n9DVZ2VFlE9PDVljgxFR4oiYjh2qCFwk
UpxDhKXsZj8t4FRRe6n0KA2UEP0IgwTzk96ZPeNePeAdwlos/okI6iNR08P96n5u
Ua4s5EvrExYpxz2WQKuZ4F+vuyN9A8mZXMtBICcIZPsbzAjGcnw5qZBs2YH7k5SQ
zXk16jTVYfSzBdemBjIm9sqgAryzrZNdL/qN4X5O9Br9ThO8rAM2HRUXCdcqQEP6
eEVpar+l4tY5Tto1zw0IRojl8lBy4Ks20edrcVqfEqwSfHo157tZM5ku4LsrYGCJ
xBOsjocIj8XjwdPIs5tmnL2Dl5sdqaL8R7da/IoIseFEZqoOnjHKjJf2VG1eH7W7
M0XvB18a1BW67ccNIxOs7SQVJBcZHWcAZk9Q/gCRWiqDD11HeXEqt3R/EsZCSvFR
kJp/AoB9pDUdnVxEzg7r6ZEU4dk8U5l0UtUadc9+ca2eNakrapPSmlPpF03z8NtS
/aNBeZQ0r1VrXpPaFBE+eAmCMhOZElLYQthmu5qtbEUPmYxrDF/aC64X8ttycoa0
k/dLWmhkQqYN4EBtUVQfpX9tgZlH50mGhskupEtf1Zcerd9lt775Jx5+7Cm922B1
g/ijW4+ehLcnSxfnUrB+TreXzAM7c9Q1fP0i6PL0AX6bUQ+2Ygxl1NNqMf+AvORu
HX4Rd1y8OrXAIBzfs/3mnz//8wmLqmQUfM1jVAPjrjwQdRTy1bZrHjGdOnO4VrS0
t2um10Kh7NyoG4PO5BeI4kVifMqx5X5e9y0vtacgBt9PSPkXATuyeARdtLLrfd22
6/LlD9u/LyeJtkTEgosK4G9qgJuUnsa6wZZK4cd0qM524jG8HZ+gQHQ+fP4lajws
UXWOTld0Z3BRvxlqVNCprGo55/sr8DpG+NDIx/mTg+zpMlNuT7y63vcRAzwhyI/B
2V9iGbOfJuC64UMBd3JEi53r+NNJ1r+6eHKPQ/H0ANeitETTYJR/hgIpeSN3f7/k
y3GvEW/2pu5vmACJFCPjSs+Rv3qTSVagakkvtufgyY2PwZe/czhm1MDdMuKBLT7M
jDDYV333X3AgheEkzsACuQqUQ7soIKFo2SenNumijSu8UzdWkaNWtpTAK9KOUBVR
S9LO5MmqW1kKjTPOm3gtwmUZP41fsEDNjsRUi7fJvi0k16VDf9+ekV3Em4BPkw+t
P5PrOW3B4d0wCcO/ReBQ6Cls8LNL+SP//CJk5pKeyY0g8UkY+4aCBviCQ4C1Yzfl
2+w3x5c9dYP+8b+imwWEN/YxdokQdymou8FeYWP1Fug2ZeWWlObWiJXDH2SRR+uZ
wArc5jZC2dK5Mz2xtoyx2fzHQVcxLl7qbEhNIVafGPpJItNBd/Gi8m2rvDPkSzGH
K6hdz37tLk2/abKD3nhVwWfoIf7ou0+dZmIRx42I0LHIl0bLOlqicAQh4j7mpaiv
YmQd2OFU1EAmK2THLWgTDhc4m4AYOSWChAZCsIazC8F7Cn8l4pC/wlCXFZ5N10bI
osXVCJVZAm1bi4a8QVrTTMnP8I51bYzc76QUxjjT7GiYWJrhVNdw+kW5JDDZsu7X
6LH/rHuYzMeUWNR+/31uT+mJlUU3DEe+IlVD6/3M/R/3Yo7MkVS0Lk2Qp+GZpXQ5
RwoMVjMwgup4U89BISARIcmZDlZVURlnHJhYiGF67wGhz2b4rXH47vXzRkhaT4j6
V6bUT4h0Ooc/UA0T5NGJeusfVRqC8Rhlj1BZen+XEC/7Mq/jvNRrvCZMfPtSWliU
1rvvOawVgcM51UStkFsEPio0KTvU8coyzpfiL/anjeWXcEUY7H73p7KH1Y7zT5jP
7Z8Jdujr/gwgO7zaByJfWD92KP3xCTwnS5lrIxyywkJxCWbuUwjBl1ZHkUNdBD71
20FfcEW+G5+1aWrJb+ThDzyfZ7+8BKFTtLtDguVseo98llmsFiGr3QcXKl0Cipox
g7uYRjAZyBYEwfpdUcLlxpp1dl9HPXGDmrP3C1QKl9ZRNzHUKziWTN5bvN7bk7zF
2qSCfORBjTlmo6nNVHaQfTTjbm6XsePveOGxGMfnc0LKuyO1+woYZgpAhFhIm3DL
5yu+U5Aq1EvuQWX7q9pZ/0QRU1C1OBxVVDeR4o1KMjiVPh5FHJlaRDlW3ppUjcOP
oOjP/Y7tFwLCcMm3JnxOtMDJk/uJWPGRTV914Vn0iwJ6S52zUkFtpe1h9SfkPBDi
lJjWpFfAKaohzduP4l+64qG8yMz9jNtWDgWJHgBJd6S5/S3/jFmuniPgjpjZbrq5
BH95mevj85yQgYKvkrfFkGFjoZesE8tC+W63JMwT/UgvpPTG5cpK+ZQAFmTAzmlI
0+D2cWO51LY82Ra8XA4qboQPq94aJIZ7pM6dEJnC5flNbA/38ud6RMaOJMvBfD8z
sY72IJvAeBXj5N3XMS9z00eVm25b4wJO6/56WpFDuDw4F9IAWYLlWNQqpTk58s3I
ZlKvdqPqMppcLg+NdajDwV7bvJDXIbuQini6VnAWw8E4Dfp4S0iYtPwXvCOYzkMJ
74CxR/v9qCx13msfkowCvzEEsMKJujQs2ymEA/e+dXn54h+Hy/t0/ISun3IJpF6j
NA3IkCcknD7FOf9mRQhzQ9sKAz19Hdo8UGvd6HekQUYgV3oCRShpgAnB9dbOjxqK
tG7Yk/argDZ1I9/dWz9+W3Kc0rA7tzRd2nnwFk+9u49hvbyB5qo4HIJXIZpB5wEM
BcUWtc6xOz8pv09U/5pN7EYP5NEvzMTl++u/q+W0RT35cpeKvyzK19iw5R5Zz+eJ
HbgwvXIvnSaaqxeQtNRQ1dMMDT2rlOMy0tz7KXV7uXTBUYfsz8Y289ua10Hfe97k
dEuaRyeVFKUPXdXUS3/S9V2WiIey4XwwtkYkKYvko2XfZCAbplFF0JY2kkWHrfTk
5+6rTqoi41Qtj7nPK8UDW7cAOSPx9krGz34K1zPvJIuJL0/hLrcQXUF0MqdxM1lj
e5vTnEJ+xbXqcwf/daXgKaE4rNVAfdngaWQn35iThdmlheTvQgKPnetTAXTMKNO8
HjmNgBKcO/D90oerN9FLThXlRxpYKwKcyBr7V/pcJU0aAdlVPJjpAlSDnBoKOh0f
D3FXdP/p9yG4XgKVHfRP3bnjEIyUf8GywMCOkr6JCPdhDjVCXmlmxC06IasFdf8T
5xtPtTTQ3TRnKWGxNB08ZI+s41JgxwrOKSGTXnA+bQ481FhzpV8CaIoSTN1yy1oT
d3956ZFnKDLJO/lQiS+ExMzImZX5eovckgBxRtidDlUXJHgVIVk8tOBB0/FeG3oK
2SyvH3MWCVeOFyDTJXain0LWhyJyIJViXYSy2FBYSD6zt11+kj1dkYXSfd1CCzF7
Z8is8esYTbVN+YPl27owDVMWEzFZZEucCq4eFdpKac7WsLoytmMOVItC13Ju3LSS
dOv86FwM/IXFFJKeB1/GB1w1dN9WEhcke3879Rys3up6ahmpLsMzysC6xmR1yzih
FVusRq0VgiDiJL/tZsO2+pchLcYMtDKiLYR2qIncVJwGo0ox7egBwbDYhyqZw7+8
w8LN2jK6BXanSo8O5cDfGWT4a91Rcd+ercKuay7KbabStwML267/W+zX7fAANWtu
hj3++IdqIN+fN6maxDS0yVrUIslPNu5mBoIxupNVNa5JKV2IaA/ZLwEzla7CRKEI
mL4pBxNGZJcAmgcQHyVnHjPB9cUT7qOV5oXi3g1XAiz+8g9CV9js7RpnSIzXsLu3
wuE6ibanD+wwvARdO2Ed7X6uOt3T8iWky3GIyMnw3T0h91oaLFToynV729DAftjc
5SIFNBXtXLAZUYLGWPtUECsIVk/JUZRGuZuCr9fTX7l8bOb4NTa0oUYIqYFg7ClA
Bz3KjCrcojsaGoXgb7CkR5lSiKdh66umpoBhhZwHZJFav2PODIltidgruf9o5fgD
AdTbZg1PaiJNfPZusjM2E7+KI5ZpRtUGsM4u0PvThV1r/zLQp/83wGFKsIn27IW6
vUAqYi4PpNRvndj/2GYZzTCRS21UROzUMirTPzifiRbgfICkZYYgmjlOrDLdHkWx
efX8jGj3YNgl4HDdkrY9Msk/y2yFRNR7mSwfCE0nqSK8Nd2rvqLAGp9Ga3n7A+Id
N26w5gqWoGC09auN26KWC5yStGZsNsi/VE4xdqyyErKX7tBibRAjs6QjZGIr3e4z
TP23PTNoaW7Dh+UqbklSTcwqT1q1qkFclENfJ/zgw+eZBVwG7+xltkV9H27cArFd
nmw2E3yi5RcbRucvjoBrS3awq+20banEdglBJHzMoeMeca/om6FUCqAAP8cwQNAX
K/xiojK5BsbmaTlqH8WEAoRInDddysQmpefF1R+T0bGGRBt6aphxyCk9DNZarfvv
+1XPaJeb/FmtVK9Yzhv8fKV1SzfaC+dmY2kFCaL/TWPyVhY3NQYi4VWPzI2hU7OA
efjIKVzOIDc/GnuJIGd1IGA0d4OgdSnNAd+Tm4sVabBqVK30u2dDCelvUJrlTcJd
u9tmkobsU5rArzWHLoNZ0bDxj12DagT/iC6fGjx9pl6X25jSxwBTsRcsVJsfPdfN
tDvHA4seD06wLBi3Ihzk1rW4sGSLHAxymCfnwnIquKe0avGo0J6eQI4ZrDUh4f+S
o1F/CibmrbRfTVwdQRkIyQfSGGCvAddKQ5/ePxulShE8PbUMK0XnRkiibAFveI+n
ZwT+vK0x4B/caLN5KXV2lKNN1/B5vkrbHCvzbnxt8CQagqoahNNRZZo9a83sNxa1
R+sLHiK1ewwdpkEjfDZg8T5zPj/Q9ZVr7q+c+lOz8TbUlubQbSP066AvKfnJYjQe
sMPkcc5iG1/dE3ZpoHQRDbuY9Za6F2P2uGOOBnCfOgfN/W6p8b9SRDa/j5gacIn4
r7ktp7BIzzjOkFax2m5kZj416RwBEV7zKvgBXyJlelZKJUUUA9IBprYo4QbR/aeQ
TYR/i5Ngd8Gmnm00dVUhyPmTr5U11wozwMxU8hZPMwzGPqgubd/RvkcbvDBNtzWf
SGILxAz4BYqlYlkmBcC5/hH8Vo3kSL5mZlAJfA0RhICJdyWpsHOSCXhXDEBl5EGS
XBx06SPzFr8NdXwsNKbBv1WoGInpiKoY7VZTfuyA7Ek7M/BiRUTeesWKcB7wAXNO
cSbm/O13goMY9vOTMpvxeCKOvvxjLBS3N8rJEowhHk4bI1SQR2xk6hZIQKXpMCAr
6wlRBLzGNz84nl/M2r0CANeCbqMPLZQIYe4nqAuMloEZa/4wiW9rXaExDJwxjz9Q
ckKp1Fimyq+vXtnbz8iRYt3r/9n1VhwLNyTA83gd1+Ed9pizhfDqLC+4Znd9Kk7K
KLjOtZ8Y0ydiK9pP9PXQjK1ojy/jwgZAVd5op2+8dOJTChfYllrEw94DGKTtUL0l
cnYF+N3D6FZJ276GYTr5U/ccn5Q6hF1IgPOLmkXfBPcfyIH5/MveHlKJRNep7fym
Mzj/waNZ36dY2xS5YmHYKscOttYJE7lcN27XVbZKVManJ8nG+1yRZ1xd2MrWZrKn
LSv1VY7wQwOrSxt3I7QpXzZ5Ga9RTWHB1iVuZ15UgPYbRZNm8kMf+ObwiTc3uH/L
0cuCyYxPqgw53eLdH2L9cI5ePQcD0ID3IbEmQaisIU0vBCQPU9r5HyyU9vS1mCXH
ULU42ZFfe3QsTsxUg8y6ohM+KIQKh7brS6hK1U2DxO9SNHO+H8brVjWvSlmLDwf4
HJtUhGz+GImk1VxjegGrBff3a/jwfcs5cv4FeoNAK+vZanZP0xKFAB8fu6AzMjvn
ezUlzSb4nmCS2wgaeCsM0z1c8LxMEv9Tx2b7Tub1dseFvIoYSEqNXbNECczypLtr
Q2/rNT+TFwnZFB+FupLOsfzZP3dfLbrHVSq7aBkklwQ9WBBP5EzXqo1Bm7JBQpF2
YmMOmoNtwhmyodMI909D4xV86j2KKHVaovpBse83s0fPYriSk6P3H3paMvjMnRAq
4qAbM14IZeTc5SJF9p6AKb7rQQ7/qsq3SBfWrCkX0qQtdUealDqXdWRjB2qKh7FX
OEieE5L/bcZueBSi+bTZO9xaOxb9HVVIpVK34uWxgJ17CnUo0HymuEzs8a+uixa0
2sglmCLP6Dt8EsbFFRVy/ZZKnA3/YAYxEOzHoC5sWZHaFvTZ39i+9JXVEzvzBlsg
/fftyKvIrGzjCoOCmvFDv1ZYwJHrdlerCkNV4xihskNo7s7fu6WbIrA/G8B29M/O
ICD7nuGMxoHa9mfGdQrOVydeevEykls/rJW5EQU1A72h/zWI8PWpg0NSlWhF+iDn
wjsjXnVKi8QbHOTFJtr50zzk/GDfi9zhVbPpQ/Qd4yC5AGKQduxGrY4Y0AurtE4q
cmOPAgsIKXgkpaVx3M11rIjNH+iAXq+lRut0nt9RNpUnVrA6Y0xtQnYLXt8qfK+a
4ZZITqcYS5fFdgOgqQFxy+FX9beUmBtULSk1A+dPlYLb+FxvfHfkPH/Zs2VNJTb6
EZDCdU6NCznIND382Vn218N0OXtHBUKMaHxTEcILHlpwHnYpp91JtUsPZI9IVpLf
hvHm8rJDg0aYfqAYUKJgR0qR/q7Q5BQYn3mNpX+s5b1aFw8ykBQHAO9jZgvaqh4R
Y9BPy5It97uzFZDyperwRU9dWnLdoZPWQDL3DOCI62I574kCTw5gdpBDhPfWpfwg
oCPwepzSG0SQMTTEOIWK9kv35qd7SkaMwdTcz69Z50hDUS1jVUTnPqC/VeZUeah6
Q5zVmCH1prdDrYQS5zGiNaxD3cthnffbki/orKs2k/S+0y2CikZEMiPugizbkMvr
v0f8WTY/0VITvqCg1JNb9CmU/VZsyEVpMJSl6PxQGpXQX8AQasZi3WC14Rar2UJ0
nTL+rbKNb8a2sleWahex1ByETBHUEflDdWsi/iAzy5hVJeOxCxd8NjB5w35Y4hm8
ViYtKfp2S6I36k/KUdLLECAmfj+OiT8R0wgVbfLbb57xwh+EVsQ5XK5n/0eq1M27
QG6EdWhHdu/FhjZGHcEgAmaQW+qk6P2woIBNK6OKzMkkxAmDPVm2mmmci4OJ8Cyr
tKakBzTRBIvS8t/yAkMcZcpZt4Kp7YQ8JftBOzN/1sijgcdmFdK6f9H12qI5p67y
hwl5bAtWJmHEdpCwU2qc2thcDUvfPYWMC39mz/S1QiO9BwXPVEQADALW5nDnFfA7
aiddI95GyvwLl8ZlUFdjd6Jx2sLSzCQwP3SybUu52EWkpsSXwmeodCyYCkK9Jc4m
iXEa8ohNDM5FaWAkwHnd/Yf2niFTiZC1alhm3CjXnYwXCN30WhzfKf1GXG6B1H9m
MNUbpAXaLKA/EGUNEdaeKCCd9b6nQVkrjCx514zkvMrFlB89CQ1vcrfB6J+cr0Bz
vm2djv+bxTxGVkF8oUbGyOslsEKVncga7XUut3G0LADSXndLCmwMttiYkzyzBoc9
aDmE5MNwpEqX5tl1tLO1Pg89+ctzE+QnZ1LZMrPrtz7ezL59dVS8bauLcyptmrP4
NnUVyIra0BHB3IVcey21I+JEg2vgLb1wu2s7118VeJV3PPNhH2p5KWbaCvE/Xufk
jB3gd2tccEWg1iIKztaE2BVMNpcg6tusrCl3wQ1fWxv8aLll4ELhu9M5nTlJsId7
P0KX25EgmAD8mWx+WM1tPaymS4lBi/hILVmhWNT7kQcju4NxNh4auVEIxEYi20F2
NCIYVxHqJQ0AuMmVCniBDo9Q9gPDq6d2MuGrC/6cbzBQlVEh0QLDT14E5qybAU1q
dRmwyg1FXL2xE7ElFSZPHGM14jVoRHRY0qFSROv5ti631yY0TfTwuwB+tsmQ53m2
PW8s1yyphR2XISCm72cFCTr/Ob08xr+ys+pd+Q+I8Pfdv/RODm8ciRfP4hfLGxTk
C0xa2n0VJaeElP10zOm0bSriadrUe6T1JAt+3gkAjPm4vCLyNIQcm9L81cT4GJRs
j+EimUxbqVnFjjPnQOVeUZ8S1Lh5kL7a4hOof6Ka2BJuIRrFx9tshEWya2mwBozV
2OQEOdzJH/scxKS4610hMifWTDsVe3sQsHQ8X9GESMpnd1ZMx0StYq8rqR44Mw1S
JZssTH01WtXkL3oQDUPoa+OVfLYBMwRTITe1tiyHERzsIXkLJtoXjGOCX4PjA1Dd
Vb+72yZYzhIYUYZRL/4BqapAvNC8TBi81eU5eogKE/SVwmyG8zoVZpmK5RgSxnUk
QImDBPV+xt/C22hDnAlErWpTe7gLFx/hxLqIpSMpmHV6KQFi4qnaNlqmOs6ksS3A
jCmwZwo1LL8Hj8HlyNTQJE45CSS/ai7ILEFA+j+on9yW5WwjGf7fiiLL90W6t99Q
pn+rJQ4YVW/wR+BnXyC0Y7NbkxKMigsOBUNjPwUVnND41q8OqcT1cjDIBxaTnL7A
D9S/HjjLk9aXNnHIr6JYDYWly3z7aGHhkToBKG4kdKwDw6erSM55Xu5P28xD+UTa
OOgnn0zV/+9e6GA6MdnT8tC6cCC7md3OuOGHtnrlg3oUU8tTvO9Ip5xWY+z844IH
HBfcVaZZgNVzhbwjgTxCDf8Pq0LUWmwlGQMjLCl/M6Vg0UjeHrFqHjoX0jdl8+1y
FzCaeMREISxNLNGgqjgRVAVu7mczeBdaGmsafXXqofDO78FFkMJzyyG05jS/yldB
fV/scJ9LZ29AmBUz8CIaPJcOaK3Ac7ZyyRwWq2xSyvVE2+e90d96dTomMDwx2pe9
dSrxY6FxmC9QzmbPTdJm6GvVP/9WJDss24zEhQkHI1PHvo1JYo8u7PpMFpiNndKQ
MWWqinm+oIkrQADSvDGBfWkg/hfzgX7bMtyBUAgYXeali70Ewf7x98YgKWi2sfNf
uZboHbE3d+kIzL+2c+5tSAGkPBUfLVHE9Be+NDb00lO3jygWRcY9Psj1OKC5Z7xY
eoXEsiIRKREq1R/19+obSXHko5YeNft6PIKJz/eczI5Y5emmH8S41jUOkqioAYgy
mmnnmBBA22MumM03T1Y2c5mQXRXoNeujPOXhl697iiHD21j2vrINS0IrOvSKukTh
M3NZN1zv4iKlo0arO4UqZS3xnPV7ktNagdOHg1DkWSWL9pSzKwJXer1r6vc+Uahs
ZASSfGwRjxbLjt169E0XWbP9S9pob9z8Nb/koVby/9n59BQMpefXyy6mRSKcPdus
mz/hW0fIByzl8A5Kv5nG5AXPp9HYY8cnbqKHSKWWvp4qlhkpDrXXJvjegQUMX7RI
G1XKjGKFkgbpKw+rTlWdNlTL4PzJke7HbxQei39D+fhAL5vVGp4alc78gPRxKE55
Rw1Itb0cPqf3Tt2HZNl7JTHN2YL59gE169Vj+C6w6Rb3rfUPPDkA/22pUE46LTrb
Cg5sLPNfew1m3QUIxrqtqXV3aCqvEJP8G+V9e5VdZQRSJEegKwlbopQ0DyG98X0B
4EfOSdoceJUh9s8i7p9ovtXfdrT/Nt6sMy2rbNE5d0JONHvmIVyUZYl751kUlhpE
KUdrEMqZm4X7YqPkuJ0QaAoV8bPXoqReSuDJjGiWdFL9ZsMRaqwRIFT0b/u/ivIt
2Yp2i87idN3mk7NnZfUcJE+cobXf3iOaQYfrgPQ4DQtPWQKzqKrBgVqt/5wq5ZGa
aRHTtw0k8izfwX5+Dv5MoLI9EXn6dekLHLx7XYaKeVaaNsXJtcqCfWwdLMLbTxi2
ROOvXhuNm4I6ShqMM+I/6aeQotC7aF9zWBm48m/UfhIOaBlvzyDI4YSgV0WLNzqP
BrXeKTXjPAWKd8Il3iH/ULs2D1KLf6Q4wML/DinkJ2sDr9Dn7svpt16Xxh6schEX
faU/wgWSVrehDlevjpXRg2Fvb4Buy63v7xhm0fCSdu6NP+/i9IwDVCA6oHpE7i+X
tMUDUOuwR138YfW2F5LBMuDdt5HxIY28F2w1+XLT7ycsUhSfzRHUD9ek2zfyV+t8
498Y1/YPs8tyMGdbk/utEpweKm7SjDClB07lnFf6IywPRzWmQdwXpxLcjrbuJcz5
9qQ6jW1+SuTlpnX/b4ymDpPHMNaxr/qnRZk9Cu/kIV8qaVmSTVX97mAhkdVfD9NR
zUnV5Ub1CTKQqfGlf34EM9ZVG2zKOSySNI3OktjO9VgdjQ79neYbXm0MmWIjrTDC
nqHo7iQCYx6pOd6zmpg25O2oT4DFhfhVi2bP6p9rJRvDawVd7SubxeBJ6FQ+U1Gh
1JtEEjEs8USrzYxgdd3BAu+jI9ZpuiZWIwTp8V65o6JD6vqyFX59AjYakEVCWVfz
cgAKAClUZRadA4ouD0M+nfb2iskbtLux3QwsjEv+SGCvCa12Gmu9s3yJDiYEn4Xe
RicQei4Otmhfv8p6LmksuicQeNiKb3eF21weHo5RCok3TrvnOw1tCKC19Bd4uXC/
6bYnh3el2jBcgVD9WD0MVx6aAP+8Mze12B1W2b576wHA5zTvenMqkpDgIqWvMpMB
BiELlONfvOxwcv/9glE2yzqEpZuDoCgIq06I2tduWlpKsNY7vkmLKEVydozMUzBW
Bf5jTTQDGLOvJfHVrLm61Td0RwEqn/2wJQfyAlU6ytG6mbkrvWYKzsUVk8Sb8VLe
c1Q/u/8O19f6Mth/b2/XM+qLFQ7m3IudLOLaHPEokmd3pLBqwwf9/4wFsQU1ma+a
ySLO8efwBfJxJMuJt8IoAe2XDJBsDetKzxkZHDqyPW3nqVIEh5vkK0ouE0ueeckE
3ZPBF17d5RwrJJ+uO1aSSrlALliPm72JTAEwRQge1ULmnvdGNb/bJwSpem7kzZ+O
Y7mt2IYs3bIM67faiIghZKgbQKRXlgG4oHiKXB3XGYMGhfxhE4KrmgJl4BlqOllW
KkaLIlz2TXkO4GhJ5WAaz3wgkXoQXr1oGBseYBcys0BFPRIozLuDXNf+LJjiqiCn
n1YTX6zXFwLnFmOBh9+vb7o52HC1Dn2YrnMeH5W9AoJK5KdpR8K6knTZpAjHsZzu
M1uSsI18hUpyqJrflkOCjNL1l5kxJpZ4oXAFbK2G7TgRWL4yqvQctb880PGXNl9G
fiCgdmtDj+0H6CNzBggMsHrsz9M+B/K0MlEU7A/oY8fKdQ6A0a6kWlEa3mNc+WY4
PCmpWEJbAhUQRugidLpdQk8qs5XHPD+FlmhbGOtuqB5chc6V8+sf+Ojtq9Jx8Mt5
WoOT9G1cHBsG30KtviwYeRiQRfMxRAwyLrRxJ0Z5kFcjkaRJ5ZQK/vRSuGMD9dZe
vSd3Jo19ihHSjG87aNSpal2tzI/WTAfvSXoJJg1cuHK4DoGQiotVkd1qqvaMDK8X
Un23u3lrdWgyM8x3u1JbUIK60qMlG1uwTOjcvbDwnn3RAqZ6g4vQO2j15sglpk69
XCkyGm2hCmgwDwJ/T/ybT51WsiCMgbxj6JHqveipMYMUyLcFh/2CYSxYbIOQCqPQ
Nu62wrLFycIsSq5UkUXbsVOenCjxA6rNLo2gPiHQs5zDOjkN6AGUbAZuYtXtGKKQ
uvYyyoNzzls7YUro/JWg6jpRriavg9jHfzxdRnFXNqD7ucQeZf+GmDTeXRMaVMQQ
J8MmlT0KPrk3CKAWqAbiFbeNb6L0SDV3Jwl1Wtp84qSMYHqDMsrUdmHAnK5IjSLD
Su9uT7egW4TTy2eOnHOHjZNPP1UbAuCB4dRP1iT92nwQvqi9x8xrUU2uxywuV0J2
InL82LNKmej48d98P+atPoYQ/gGz2Hc/GqL1hAlnwlDkNDz18N1WUo6PjQdaKPnb
88Dy9vs+pZpHI6/jpn4p6TnvDJ4J479/0/7++g2Wt6RatdKlKlEb74xew/Bjz9ev
Xcfxjv9HHwCM+SEOVD/6uH/FUVGnjuWmJudQ9T2vjpTGxUBufqibGgOfLMzCVeR9
zZ5ODGJgzuCiUHVYaM1P4f24OVO3A1o8r7vjBS2TZ/NBPqLLF5wug8sC8dz0HgBj
N7bZNa28uUfPVxmP3CT7Icv0WhlldHTUs/VqkfXVPS3Q7OYr0wW55IQz6CbPyC6q
Fz+XThcd7lyFT7DIAVL0ve9I5G7GrZyhqocRy3c6dL4CIugcq6Tkw/zDKIgsxApC
vA5ga9B0yzxstsRpwE28T9e7gee+cbB2842QJDxvWvwNSFm5afPicOUcOrCXI/TG
p3KRpMR3BRXTwJJK+a4L1r4Sp1KtcOWkyr8u1bOoYnzbzCXDawVV2U+T5YMbJXWO
Fvcp1ktOjwyusgqWkVGIBWVZvFQJWcUARpX1caI6Q7GD556eunN3jK53tjhfzpda
sHJHybWI9RFQ9hmL/aAnvKN8qPasjeV+1ZU0HRFOF+ZGEURaT9TgP4rqGl0TVE9H
QOXJGkXpE78vRKozXvqelnHGFU5KHtwzrpJuM6UMftrzrghz7pk4KP0Y/BFol1CN
/nrK1+P9MFZWWS2JaEnJwqzvml3A3dW2ZViad/Frep7H57ped+d0BncTr8D9Q4nu
J0/FXWwhL28ah36lMOz8t3N6XHvOpqE+wXsXbYHYImGlsJYCjr+Xj9rNoyeaHFrw
C1nmCktYPPz6Oa+mNBLDRcx1AMfFEBzQ1/Q0ZtoyHlmlp/efbUh0nbjKEzeAzSW/
vT/ALcBibN1uTE1Uhm2CNK/CRhcO9Lr9SrLS1zvpmK/6BGaGN+WRWklyEBwii5Yr
KlvgzgAMsE8JeO1bECFtsvujMzgiyvMxjaSe/LYF7FBVBa913iHZXC3ZBU6WIVHb
ZXrMF1kVplJ/NHsst5msP5HXExQapqBmytA3sQj57Pow4TOrt9GlHMDik6is1uFJ
ijibxAB7qjk7ygydxFiI1HQhUzWXwnxQ0fy13PEFmv0Dnru2wX+7qPnOIP8caD9Z
yBbLJPs3MKjWZcR6U6AE8zr85T3kkaM9xWhrqZJIoGXIf4V3VfV0sGpZbdHc65X9
AH5+cBAlhwBv2E00fWhDbq8/0vlevpP4WQT9qSAt4CWjSFXL0CXtZNpPjh11Jc0y
qGRhd/u6DsJsk6BOXGb+PzAD56g6m57CJbKfWGCF6Hta9R2rSbC1SMjsb+3zWlum
t8gCph/5wHcffJXrtFn4QQO2RoYp5b23/+mbJcG7mooU+smUTj/Seho2IzDHMQsY
JtNX7/yPedIPBKBuMuOnFwv8nn53QMynwC+A98vGlEqIDXD4uFrCdyX8KqqYDbP5
EFyJS9NJtGUz/kOw118Dz5pYGeJEHv3/mW4P5uv2MJhrM9ZK9JAA9s/pC/dFR4dN
mZkNFlamZtgWs7FcwBCo1Xxco/RhcLVP7LwvlnJVeE1lY2PifkNQy6fvxuCTRUx6
NZpph6Hf4vCWNfVT0kdBFyz0CaC5rba0FRB7+25xJsk4ksZ0nGMCmWLqqIM89qyI
LI5+JEQiiEw4sU7xomJFmAObGKaGliK8Z0DMmBtDGNIW5cRagvvbDLi77fCbU6Le
rfL53w4cDxnVbs79yvIgIkUyVQMlWkxg1pN+b1s/XZWKgc+ZS1SLez9sqyZE4WRu
EMd1F3ZjLWQ3z1DNVqwtzh0lEPt7TgV8C4R1fVm6s/ejVRE9NchC99RRLz4vcgun
ptNOJxS9x350DAnGeL1xxAtwJqdOUrWU4Pg4G/f5xUmLci72aM2CzWLSeLjzjiJi
05SAmlT5r18me3+/MpKB5gf19tZfPX/3rxjGsRNK9TZMwJNaEhny4xxjN58ajpC2
YMB9r/4/TmLz9TMtNQIQZkZvR3LfRZI6euWKjhNM0SnwG/C4crpT5tnaHAP6dXvb
kFZfy1f4lfnlTxBmQspii3gMFyvt7Y4tH1wKN4xKFviLUFc5kCjHXuGHKXx1MxZD
1oixvmcfxLDgZ87ivEiK7ikTZu0ICsUgM3Cc8O+dWQF+2r6kNn1E/xlApDbd/80b
u1ca6ijNPa1YKfjJy/VL3TiX1A1/jJxICLWo9z5K43fS/O+5j0MKs3syFO1tIRSR
1tjMJEisXFZKIx58/CNY+ye+Qasa4SrJrf9Vl2JrugET8JZAkD+Tnna0lU6aXOlW
VrYaRQuwfqa6W6YWZCjK/310meMe1+JRBIZVOL0zdxKkYiPcgG34wwUcHIVNV+uI
C7NAfds1EMoLSGayb/XPjPjc6Qhnr5mGBoQpOVPDw2yZ0ryBP4wCLcQNeKZ9xbiU
srkIqfD0b4i8A9/0N8RJtgfOTuxHGfaHhnMhZY1ju7DVT2fFADHKrDsfC0Y+W9bD
p0E00knNfxcWy45Y7+2SIHGNLBJkL9k5McyMt8oR0XNDPFojfspj0PooyLHMoIjh
bQLHB0eth8n9e79EOtJHezFAvTUurPiap+zl8uTn3nlGW25do66AixakccVvjiA1
aG++4uGFzZoNUF76oC+XrZOCVj4TRssaizrKfWVJohlOdNI81rSNUEBXz0l+OxN8
t+hc1zpfoDHX3Sv5c1zZiIOpeUyvhg+sISNbFPaOdH1GDzg/daw2LKzOJITmKXtM
qsvUFE/90Gf4BrmxIQJO6FSRn0ow6SQ9T6fwlJu1qBibYR4yeV3CfeSpjSroFPzL
GG8pngugRQIjs5LBtrYkAkP0iP1R1NN5yfmn2pWTMlrNEyF9bLZr2I7C7k830N4h
f46SnoRFsXaKZ3vgoXeBG6hSFBvT4oJdW4AwNxWXIIGqKAoloZLmblSXi+Ji8uHU
roXl1WRUdaE2jDm/FsqYURBN13pYLGW4v6Nx0hZ3m4MYB0hRaQ50HXaYliyOOux9
F5Z5sIi/jTG5kj2rMCp+1xuPM4KJQ5A1piL0THE96efDB46gGkmwsBzH7/4SWUPh
FD0eOXAwx06QSkIi43Zx3Zjaf/jI5dUuVpq6WqH6uQdB2jviD6McwX+w140WQMau
7FRrdOJpagDq01ORpgAjA1uwlIruUsPfOhpDDawHOPpUQcboQ8EvB3Avoh9qzsDl
OSShz1y3Qj0qMcTybZ3eSAAe8HaO2R+gCf7fLQ3DBbBo5rwaf06ceXqAaL8YzRhI
3NE0q6sxk6D9aYwbrBATNlz6YkhoEZbCeA4FEs8RvIh9gP5g2RvDtRkEh3p954BN
z2kwm71HqPjjc8bSLYEAaLDmI6zhjXcGV/oKuShPdazyKCN2s2PGh3cvIEEdoTbW
wXIbIHgxJhTR6QE6BNNpE5tyTPAdTprzFD6WPRMqTId4XYQgyHy9/AyIuD1KNil3
nrVitrmHkJFWtee13UdXSECPU8vXfotZ8r7c6Q8r7PF6WbiwehXsYPkbB7d8hjRm
Sod4TaWERgGm19dAk1Hzsxx/cmNdtRAd/YePVPU4NDwvfRMkwsAe9dLoW7jiy1rf
Iu8KIrO6DySz9g6anl4WjJC660I5CdGnrlqaFypelC7vYPEbyUrHgKhynwoHCI5+
rK12foL7ZnMf8ka5zMmK+1N8qcUet25kuEI+A/8TLyd/IOKILdg4tmm1yrhYVvrR
dfdX/gRxwNmVWN0e9qYQ2MsHXdt3G+fUVvQn5sCilHneFakPsZLrq3JfuKA+5Tc7
j8iIOOKjKRru2cFLnJitqjp97dkDBltqIM0QzQ1Ba6OrPyeLKjbdlZ92P0cBvelr
tUS7Xm4g2FesMUsNHQ9Lios1q6iN1ombHcuihTvTeeyQjVqT4fpsFDEG4Bwixb7i
eE7IWWQahnGeMuo6ljmOU3nN2io7VW2sMAC3SklVT5ZgevZNesEfnHHmEAeYmveo
gEuYgKv4fSUcHDuaNGvrurP78tCdZTR04M043zCqKWkdmEW5ojyo3Kmkz8QqCfuL
PTHIDCelwrxqylKCYErj71MjfLm1ye0LETsfZkKTDTeWJ3DQz0JOjIuP23twZ6OQ
aKXb7RKCwAjKxPHs/+SUhfjhtG6TZDSz4cPQzS6pgUhgGtFtp6fS/crKB7F4oGsS
81qEy6Yb4YhxOWr0PgQvkt05oqJzbrQg116v3H4DXpZjA/g1u+sjESPmrhUuLhlr
XNmoPyxfmOv4XhgrKV5Lc/ZzTdSlVyAhjCfXNIYEv//CPfDuQshYNgoofx3C/TQR
5gYizv0qFG8XTNM//rmfxnuec1qud5tlFCGQobc4mWH7Qe2eMUze+Q0e/I+ocMJE
8AdcdMwac77mIMqRZBh2xfBNqvNlcErMP17YOC72lG0jOqLexfwI4ifwOlO6xpTV
eGaXyFsQnNRq4WQkfk35t4OOL+Q8zLsfUUPxgShe8mKC9nAmwrRHus2en/HgLCVB
VTPjwkp/18+8O3N6PdgB/zBciqVIAR+eus22uz8q0eTZqSdZfOLUJeG7y/BLOsDn
VHwFamTF5hfX2uP1Z28/CyXzCCoEl+wWJg113USt1yx+PRbR8Z+UPWdQq51uQusC
+k0/beWVwkFnMsPsERPOlYE5NEGzYk+0rFB1FxiYghgoSulmNYGrcW0KaLZ1rmfn
jzIq9uqrs9jSwRUNPU9tgSQh5F3aufx8PwfoEY/5Cun1twSlIcVxFaWyTCO5KhSA
OUohLef4XEPxNI/VVbDiLpXXBl0GiK9K4DYrCXQLtvkpP2sflqvDr5g06Cdkavm9
ZmOoYJq5+wR5ApINh8cWSGrt7qNPMPTG1ZES3x9r/PSZuwxL21Mxj6wsHXNYDbO/
8BjbcJFZ2ebzEP06K+vlmlRPqbuOj/Wm1xKX72QryFRWJX3bsKFbJLZJZftlVE5y
VyfY0Xdi453sBATKhJQT/xUNBZxPvcKrMOyi+1LIHyjT7vF4nIzNaqi6IWVOK2ho
PKCDSgm8smEuJHYJwC+AhDC1jXV06jpRevOpM1MkZc0doDHXakxeqy6TgAZH7Oa0
08nGpAd82wio0rE9D3/QU5HqFFCbu10QQ7V7FPx3Z1IOJ9ebkXE5W7COJY7T+WLs
X4mu204fEArv8Un4QdqSR5iHY5o9MGpAlXxlL8nPUBEBmoRtKLwN7hv5LUbTrX6o
hKeIc4JUREf3u2LZx77DwwcGSY1+ToPYluhdRfCrWkhcmXTndaaVjXMM0CIT+5zL
87Hk39NqeacX7KsDdJDaAaW2BAwLxFNBI79y2+JsipVFQjXAnWW5xF7J8PvoBxU6
ZsQwgCaNsEPQUnJcZMoIQM4/ujp6gPD4+IzC15T3bX+AhoR0FpXUIE/9yOkSDoaf
KoSNfAe1RBo9wB1g0/c/Jeam0jKk/grL6OZf9wXU02E7CE33CXMv+XoOoAwlWfGW
0rANPfQpHQaaMiCY4pxpuuG0pCa3M4k5cCH6swOL95ZJrkM+vJR6643H0wBLoYoA
VAr7Wnnqmqv87pFjkMhkU2YhvLtyh8W7WUvuLje5tYodE5dN03arULbU4dlpvmdT
tJJpvnMXUy7U64tlKIPj3xD6bSw5AlsPfDAhoKO2ZPJoUhEopOIEjoh647Np4/yQ
h6d7DcCR6CRtDeyprDE7auN2O5Bw1rYXhPMAaJIY837Mx3i4KJQ77I2xEt2fBG++
swmZmXYfDAnjojTUwtDjVnvbS+HMm0+driDSbecB8CJW7724aLVwGrCa5M2IYl8V
ONGPf29dBelFzNTXPrugNBlo//GV0ImAJ3BCuDB7LTFZanmgY/nOotTjKox2Grpg
6FCRCcEXSFQj8Z3wvxGi5CD/i8BL3XeZzt0+4GHOhFQ1DXjawom8RZlNgmbx/fuB
+vvETqBXi8tYb6+oNEoSlw58amVzyU+62zdoM1nXZQT8d/SLZ9+24WRbQ/6ojXlH
B74pQ/89Rg5LPHRh+wmiRNd/bXNGJiqZWSxxLxr1yGkE6W+Jo95S6bGpsD/wryTy
/XVuWLjGz5DDBDzvgHcHTgsWH+IAw0bQJOcbb/2umN3uOC/RKrTr9nFCkcn0MigF
wLz8msXXNbglNwm/uc0UYFSuMhtBmV1kaB1v+ALP55kX07HEiNY92TBO9Zbrk5NT
DGMjs++8mLW51S1ZCNHIzu11n0yTT/HKTMjGAJfzRPmy/pMLfIDTF9XECQpSPVGB
4vhe6FT/P8QPqkBAxOPcfb+SjbykZt4NDnzmmyQUfLAWBGrw59Rq4P0pEHU1Pg3i
Oatuo+3f/oEV9RFJUjKjJylkxzvLfssQ1MG1ltnys1rgOcjVRu5ls3O53eUhkSiV
QXf1kTBMq/Frf34a+O6rejY0TWdfH/oHw0RnyPMye/9rpzFT1ownHL9LgYoQDu6i
JVTc79mjict0HQJEYnCf/0wA6HKbktji5Lea4xlC0pFPDSrwfJSQWIrY/3VGr3u8
RYjczl3Ox2KdNvVF49g43x1NWevs5jk3GY8Lafa00tj8Htop4j70uVjjoKJtTzor
ls/2ba1JxG09Syui12wbqZV8cM3HSXYzEKWvJplHeZalgEm3pSSFdSmMl6tNSX+9
K17UmK7ZTGIe0+okK+h7Z7MXoTcByeDSQt2IzLQSMd6khD0i/irUF91XtFFM4SfL
0dhfrmTqIj6cBqtcxqzi5kPs4WAUXzv4+LLtf2PNqgHAauhmTPxxms2yliXMdqUp
I2eB9AA6tm9JmILhKezH7eU21q2JVATUHcAScrGxLY48qGUO9OfojQhDlGLdZCyM
RP25rSQNjQfhpNHiYKZQjoWgCAIiEh/5UP0B1xFMArBZRCbJfB+TSM9NIgHGo0F7
uHwZ49CCiG+0H9qvSB8MJXTZ24tdppKt0/tR4iPHCdDmr64G+K4hav4GWmTnfkIU
goNDHpGgwJDnzAMbsebJEquy3wNRTWQJW/dzFsU7GgrwpjHVfKX4bR2FcAsGSHrC
+tTXMHPVNpBT9OENAYNDr7gd/q63OzNrFoDYy0kQJBYdWB9rs3poUXTJkFwlK1+M
fu8xEZx7WvkgVXUDaU4Y0eoUIX6vwFYyq1EBkJiEzzotkW1Vj1vpuhCTQibL6g6a
wQv6oRFq2LhPgItYSdHFqazmdIaZkqhuV9gusR/BGzxE+ByTSO8sdro/8ncxdJHG
a2g/ENnFDc6vZqk/VAYFGoCc8x0oHgMKH30TuXA8KurjE6+ygIJvpS4aEJKZdgTV
CheMqBA/6X+KPcDqsPvv+j26t295J/DO4Qwac2GMXU6Wem6z2nP78DTMlkqeEcJw
9sfveygTIUFpPZxcev8fA9WY6QL5wprdi+rPeza8b5HOct1TdLrrwtmKpPxdZtR8
AN9wrhSsWm2ZcYWYMHX7dh8k3v4J9PZaXlmKeIOGe2i8H/tWdcLczkMlyH1vRm88
sy7yZbPBNRmzWg1TdCSCRQkGo2zijkuFbLPd28YFfIyUK1Um81Ei1crAbM5MNwQR
MTEqbX2VdtKNFtbApKlE33NX2G8XDsx5BkZ5PRIAZngYrN3E/4DGqG0KIrbsjhfN
3CYgS524OkBJ58paaA2HbuqKtZ2B/s8aNSFB034l8qLzrU6d0eSTgOkCjmw9NFPR
mx+wcBsk3jNzpcKvT4F+5YYqMiEABOYWPlBb0WrOk7WkkWlIuD6WMZTnPYmCY4FI
KEhVV5xg1o2Jv/zuVwb5COBQFrRLshFFiu6LMnOKI3xgNoooLmuLnCdl8UzQVGtS
XA5yTOFZGV/CqvuLfucdpfFIcWCIVI3Vdz7MdTsc1ZlPLDsnga1V+NHvQZN2XkAE
W/7xGen8GjdL2Dy2UkmP9HW3POY9PQ/hAYEjtjNpKP1rs+Evj3Je0LuePAXUOdFQ
lx17DIat+NXRRRS5L6fKA4kwmFZTd6p7xXhjhgs+MEA+d1YCV3D91+z8/UZPCpHK
5WSkvgZaC/bg9X3ezOMb6Iv0oN8m0PMZJjwnaWqKDwPNtDGRFOGhUOn7gx4xFd6j
H+CCobdhE3BPqMEN2mZMP5ySOaXR7GBjRtoM8Kyy3lEx365DLFwAJQPtEPxDu7zk
8ujZ1lHOfrAGhiRJ+ZPu615t6NVygh8adm7StYV7hgr2SBpGFQBqo0juITzFJ6k3
jHED9L/eX3PIXmzfxD9qnPJFemCHuwjA55W8KWUhBqkUDUqpZpROdIVyniF2TX4V
Ln4QzdY1PCaE+TXQtKysHXmTurGpmImajRk3uzWDBpv/hHH94YL3PO1eKSFvjzsC
LTH0KLjSJW1VGf9PRaUtFbHVqHOHzKWewerw55D4ZhvzmeTshFlkB9Mjd1mJh/Nk
MZJ3YZqpFHUUSuUsFyqleyr9GZNe0wgkG6bXlUK2MKaQ9dCiwre0ExJqRA4TwzBu
JNl+X1h/rqiUYLWd/pmA2ndfwM+PcMJc8cYYk54M7xmD8VvO6bMr3HdIzVACK9yp
fXoBn+e3pxP1qaQD+MXFVBZuNANrTbUif156jwBr1fT2HuDzqEUy8c21GL7tYjns
juSOlXbwlQ2tzMEhS7m5fpZ/Bd4VSsKThoYUWNK22j8AvnOT+lBk3xMiabpPmlGW
+OS5oEw+bCzzOuhzGhtjz8kuxTUl2Io9R5mAV0tN/CQprYKAd8pWLre4Shw/kDru
CtWXbNqOBcKjDV6gHx830aKFpB0eMeWwihFetPCxdvpLNRlh4jcBSAeKBTOGOv3c
V6qUIJ4SkKOchQpR0naxZjMyGvyi8ZChceQ0SLbOLPNJhlBQWYqyFyTD2PbBdxL3
JLd/eqF1Zz2Xj+7NWQKV8upd77GJBjQDdFb3VrH159qfhby9jD19s4u/Mj2a4HGW
zclcPyl/MGGiItPbhU5DRJA3BiDvFyIQS9A/AqRf+6sV8ijBeSiBPpO/oO1/lAJB
rlQPmeyU6CiAgjDjmh2hwxo9yJ4HOylw2i6FnDunU0kuwf6/G5QpVS9G6YgaNnvN
FvNfEUHL3rkqYqPBrYMKWZY3VJd5+yXiQGYf3wtmPtMxNA40pQElv7DKLMY8pFIX
tUkq08PDbwGm2CR0y0n5KT7ZO6Rpt9cbX6v8Tg+pJYogmnAkaC4tSv/HG0wFs+ce
4qvLzAkNtyk5xBhjjOxte0I3TQm2uwLlYqS9GBj+XXESFcOgcJuIw2f1THPxH1XX
RkMzWknDFOLtidP8uX0hyIgGrpCVfWg+bNbmD16pOMmsf1wEt2Off2QlUzIkbBEK
mKIg2rWYbpheBJwqeVemrqs9Wrf6Xffhxrx5X9vNFJljIUwzdbE7X/k/ezJL3jyb
0s/J2agOUNGkDF2mBbG0JrRq7p7D91U4uDCA4HSMSmQFivMhJQEfwuXtdgGiQa96
VQ/2C576SVXBW1LWQDwnwxpFUDMwYpM9oURz+xLWOHuW9T4QbJLPrnxR6Yq39SUM
DvRLsBVud2N+q08l4rkhLlKX3puCnYXfGtxqCE+dY1r185y7E9h4i2xePvLHb4Nz
6PwEg7qSYe7Cdvi7Toze8P+azUG5EBkEQHQDy9F2hb0jmi8Nn9iqNGeAP7O0EwXm
qDjKw3QTCppr4L5TADnVTxBrVEVSNUEwNShloOqlCK9Fe6uOjZ9uDCWO3iGSX3qg
EUPMPB5rVSQ62ibtmFKjmfU8RfVKRCXkYDF+jhhBxUdliP//RFKFGrrg5EVn34h4
eJhnHQLBIy3qIUSqhYSFaQuJ4/qKDoYaj/ncIRucujwFEaNXWdWeVLySbArjJV0w
icQzgAn9PYPeOLToWAjX344h3ljtcOkdTcqMeTCPskmIGQ8epKrCjHCSR441cQ84
1zkznIts1LEDdZSZphgKmPfzvkdpIHXTcwsoppaMsRelP9/i59zfbOnO+5FfC7/J
Cb7X7Ct4P2Jk91/cecCqZhaLjSug/bvXcrMheuH3k41r0Xe3p6I0ZkPe+DNrobuN
LSqrpZHznEVc7mCBUHZXiz8TDvjQyV4h9rwYPr35YXkNa29T5jf0Y1R74OnPlSzS
VDvty12gl3mQGteCqddQ32Bled4krZVMCCWsEWJf3TkdcCUxB22+mUwAGcqE7kvw
7exT8UUJ52OsHLQ6xYXWq9cx1PwJgNc5dbzhl8QtLvDGvsOf8GV5AQy2pfkyHKW7
Vb3QlN2+6F8lh1mixjRcprpSRBm4mcxUGgiz9RMFlAwNIdjYzB4zE/pJ8NZhmkfg
7fsZr0nVgTm0FiUfmoRmGwH+9/Hn8VSULeKPKXBZFoztZ9rAeHAq/8INGJu/WEHs
tdWZc46RDvyksvYdxzCFg152WoyZhYfVf2dRVBS9C7dHy3uMawuO9U2aydjDLInJ
U4ATWuCm22d489y1vUS8YuCrbF43OhRsfzYBvnTzzhlePn3IGKI4gVTn61GgS4nK
mTwgZ7/PeToXq+FpfTcjkCvm8YQLHGNSUu46hEGE4GiIqq25snNMXqU+opkqnBSl
jg24E2RWwI2nwRPyJmRlYf99WDlA7EzH9gELt8SyFosD4qg971P5Sli/V7NEY7z+
wXWLz06443ulBwCkUaE8H8hccZ2brJW8CMspSx3ix2CJtSvPUSz/3IB+esj9ooMF
M82OIHokX1/eRb2TBim+T0VqZHLQgd+0YxLmhXftrJ3kMMpLTFLfC3faDV+djr6Y
XY/tMwRG1e1HpDCZWkPo4umlXafJMT+id9cK9QoMsBsYZYA3K/LJ3jmpV0OHUXUU
3DnrqzBZGYy7+fZlhW5o1yQjFaS9VtUixbvhKK44FjRsZKPQ9ks8l1sPujsM8l6B
LcMyTqvIOXdAr3DQxOHapN2bY9NzAAPgQYbS8jXaUdgwBEtE9PBkxOILOzDPpJS6
78mcZfa/tA9LUrvgQQiNqG5QetCAHM8D0DYiuwyJZqeagKbQrjgHoZTzgVo2KMg+
c6ZkNn0FdZdem4pApg9iVpwfjdHUIO20FdFTArSLgTeSPwZWZq6u2awculx4n7Gw
kq8TSL/+c+sDVPnGtBATv4pLK/dcbeDsjt8YhoRIo+Pwh33hNLmWk/edZLdeST97
wjnTjzZwv1gBKkMlbman8yPP6CeE3bUycBVBTEj7s/zyD74WkVBGScCuUycdvrN9
PvjNWFNwefQLM8/SJnOoup1mpFS3Lcx/BaoiQydoOL4Os1y3zrBxsK3/6cq5FHH1
3EmT+S2xi1gs7YQdaTMlslYeoT4T3TNpbaxgTYPzGkuii/ETUXxpl4MLWzjLx7pU
HfObTAIckv78xB3h7zZuPBWYBBKeZ5fMGWfY01nrLhOc76rdF4jCmU4OURxLm2b2
6Y6wpv2OyLLDwGI7wjHED8OEaOxq2b5TTyj5LJ4a71iarqNwc2wFVrlgfyMtLNxl
Aw7Ohp2gapE17fjIBaPO84Ka6s5BjenDdDRh0FH4QkUvEwE+qC7hARGRAZeHDdt0
zPkZcFYw8GotrPRFY5b1p8jFF5u//+F/kfRFCMvVLnwPeL0MMbRXwXlHhsYqWI5q
4JVQeyqIv3BFVmsuj7WQTsiC+zna3FbTGmc7b6bGH4WZ8liQeC+LjTzwTy5MTRBS
HvbQDCloO10oXs1EBtHZqgqyIpJpQK++c2HbYdY9IevoI3fmAzf7fosE8/Alo2dh
aEegDwrLXg7OYM35ICGOmT7WfTn9rxosJNUyVCVJeV/O0jY5OqHRR6lyuS/RwaP/
AAwPyZW3CtC4UhgRvMFXdMIWc87HoGewwQ/4hzMHVl5hR5swNfIRrpAr4qAQEswS
XJHeCnetmfxI8KmE27yIIMVDP9yrBBv6L8biw9nESg9QFDhX1BmblKvrY36LHQ3c
b/itxUevPdSHw9OvodqS1I7Ecnjq9Mx4Z6JOZ/ECXsXuGw46hYf5wAm2xAGpemq3
wFJ4wMUTXRvu77qBeKqcELmWKxh90y78wjt8REw8SR0RVLX6O+KxLRunV7ldgFzh
V8r1bf2bi/HcL3H0SNkKiccQ6giJOAQtAxf/VtVCyjUryUSwmq8fx+lyl6xaGJZP
F5w/Caep1SNyqRE1Ou37kATZetnFuDXP1oHBcxKOA7I0Q4dxTJvoeDOqDjmz3u11
g8FJ5EOXXwoZS46rYeVhmDv597zctOr0xVVQ5+qG5KoK/xg0QXzt6Qb63yx645bd
7GIZG58bK8FkrXFzPdPjsQKLeJ8ZF1lWrZrYhT08Hl00hS/oA5JPTSWiAAAf1IP0
MDZ7ZnMG4QNN7XpcxsTTzqvDJr/0PgXyby7R1Zh1He5Dj1Kt3nVkdpsi8+PHvOXH
ayPqA0Tk3OBgsh3p3Jqk1LoE2FBssdeN4XOyO9Z/RmJsEQzvmxLP71ocdiWMoQQ2
Ds07e7Lunva2ymXkkAn2Wz6LTS8DiByQr51jv8E7+M7MzqIi2+0gsViUO9QdLyDJ
Xp0WQ80aTB8KBrVtW5dActBLrM2cLoUqF+3rXNE/LGlRHQgl43uzvgAx77QWyIKn
mE3+xFwgbzDB7LUT8WO2TZcLaJqU0VphyEUiTSvm0hn5GgLG7/XFNyBHstpwsKnr
LVrIPW1y1ChIB5jZk4soNJKhJ92bRZDgGmle/asxAtRz6fjeLpoo5sk5/8Mv61sr
Wszmzq9YidOV2tHwdYsZcs2TdZLHcTSQKGvljCK6nnuoOh363aWRoLMk5tU9OHei
TC7WIOffU/wGsiggLBi6dnhhup8w+mZjBno84DPJPj+QqfmvRgL/k1yjFXvV2jdw
tuE8xwbV64fUNoCwFIyTai35U7ZPig4T3sPa7hnK7WySI0uUByOs0QcV/WfOpyfv
tOxOsTUjaA+FBXTWRm7QrEn0ow6XCBbb0+L8gVKkAOzc3jyG7AnfRQt9ptQNGSl9
tClukxCH4wi84p0OnnE8rMIkQxRJOXmjsYmlCVf2G9iN5zwOLTE20yFqm09wBqa2
tQFUMb09IsWXofMyxITXlGqxz8pHJlYXDvc5rnInIlJ8Se1XXxaiEZOvt2txcLFc
IP3WWrnRS97rWT0MaxcBTmB7tq6q+/3520ejCujCZnpKYEsT6zMQdJlAw1zK8erg
or+8gLLUQ/i6ti4Ij+/JZDjAz1N64y2YAnLi/qA1hLKr6EVQPDI6F90sJcUa8uqC
KGeMnPoiYK7VnBz6inU3Gs7VBEOVI8/gESahfBlAL35mXPv0+CUEGQlVrn469xhP
qaNMxk6hlsntpPgX4a5+2bzUqibHcYNzngsGWAVskGxtRNkqONFxQkn0ZwppzX5d
OzE/YiFfTj7sThZ77vUkcqgic0ymnkO14GEycXmsZSPdCxPsWhrtt9a3zgCmWJHl
rBj4FTDnHib1xBnRJdE73xQlwi5m43agYsQ4XnRMAStWWYxZrQRHRuHQAjsBLCYX
Hikyo4hG3xsKw66CdebxbqNPaPTYRVJwccWDuJqxTzZbSwPGszvrf5TtF50RexqL
WXbSnNK/sbgCNTNQHn3DYEbetI+rLPJBtA4C9W3JR9ldp4baeWUOmSn34oGxv47A
eJmJg6RpqPwZOaRrbNaaTsKHIqdEB2Bxj6fmNY6lwP3eOOqOJIyQcxnw9LfMc28d
S3RNkFgViBJOIiRGX4n+1fSp6SZsyGoGrl3B7ECNrmV9wVPJCFlKdHqaD6inb/U+
SZz56nG+U92ONDPmv46m3Bk+6XASVJJc48FXqxr8qvxdjZ93poCPBy2WHBCGq6m9
a1pmbODJ3EuV6gLJ10jvixlvaAlNsz0W0/+NDyQYMB29u93+2hNREez5oHJano5I
UoEoHD7GDY3r75guyBaQtI4FhQxaRmG3VzKeA3653nvrzHzcG3Ze3H++x3VWnD2w
MzJcqrBnklDBxc0+s0p1nlUGu1ep54htXmw8MW6MGOs+fIkz4KyebAkR0HfQbl+L
06VwpQvrvQCKDqQc4b7eOMA8hVMS4z4q5xb7EJcy7K1ts1/lMab4D2nQZegWN7vW
O1j1hr36BLPT4TFOCUiazxgGb3aJcw7aAgcO0mqUBQzMbSwakiQnQpo0nUiG8qrZ
Qq/cAl6kL+N0awdBfKx3ySVRgJUjgEgyMiSCV9BlUj7o32Iw0bOeynl2JWyQwFNf
oIcHL+kNndyAIJvZBnNk1QpFwb4pE1NfmjKuKN6l5UpTynPVNsKvYofD+Nw9Dcoz
XrwhBv9zPdWHLUf3OW9wFqgFbe/zc4KMxHQZzgrFwqI/YyL6CNDXoVwzA3KpzEXi
zUP5wAHjWApwidsc7j53Dz0VMBQmWePsA+XsOPdOa4HUEPvr3YB9gE7x2kjXXYAn
QMCHJOTO52B41NvwiVNF9hHmxBFpT32Lt5yGC1hLz35ZaU3leQ08rGf2TGMTjVVj
WuR1pkdByKNtJUCtEaqshhboA3z/RAtWcJnvSRlSDW5Q+50FDSZW9jaFBPkzCDO0
eradWqS8UsPljbWNrSSf6uglVt8V6ldQii/Ze2lRhvNTlsLTBQugknISaQW1XGd7
/e4hvUTkFVz8MT8C7c8pFKDKHSYlHC8XvzEUHOpei2Qg0/hdZKbZg0ZM446lDg4f
AaDC/aquWDFEt3zs43beSBvAHnRzm2R2IhBK3ANKcZa1R15rvTN2Hq5f2znwPi2d
v7v6gBtM+ZQtzsazcXXZuA3/hH3+TMLNw/+AJ3gOiG+ZDDmldwobxSszGf6PnM6W
vUoRRVo2YqH81kBy/Ms9F+YbiAv+qkZYV8Bxj1zgmpknvSo5Klr50o0uIDQLRH6o
xp98SgKeZR1VZp/pTfinfe+YpfA4ucExdTsSyyOBsLbD4IOKCovyVbBDJ6XtWdTz
14dyat8U3GPMhZRWgMh2ycpQRApGqwi4CmHZ+TevhfHAf7AfA/jWd3CCaJs7yPW1
41ICrgqyy3psWHX4KF8oE7PVkVpd0BSPM709Tswi3PyuknAnoB6QIJHozJXDOzVR
QiHSBpiQGvAr5XfcnfD6LObT1MryOEZgEiN6e6+DbHNbYjSDv/rFDLTZp+E4OnK8
gzwQDeL8roydOHC84LHYu02mYrRQcH671VpDauMDZIEg+PZvd9K5c8xGP38O5k7Z
P9HBBslDmYEjkNaALpAp/XOJ5mCemZyDTvUwmqGyKwfHgywSKHh4TIin5As2M7Yf
ZTf1ksMsgJIKXMJ6yCgH+s/GUsWvD7v5OSB0Y7zAGQoPANwYCzZ4sXZtssg68niH
2NZw3gAVz3nDTrIxy+LwcR+gsbCiCmbQ4v/xdQPS6eqXa+7XknYl5WpVFOqUx9VJ
B4wTGWrXrNPZC8Ml2pUyyXt5zJbyIg2KgYcxNJj90it2pmJ5b3KB6tnKqxuFUF+f
skoC3JCkguG1ApVRvhaPXzZcN6dxeeP8qLd8+N0n1aW94O3VMaBFS3/hn83Asg8E
A4f0Cs7irhqiE3u7mUwzysF7qsKLY4lZT9gSRGqwCcMJLbk5cH8/WX9ybnnQBsEA
ow7lUu+9yyuaHhsQvE2stt2UQ15jT2Jz/CLmqqwsthGvGa1dI1ctUhV8G1oF1nCm
BQN7qgFdRC4DG+prNEpguyYsiQNAxGG4W1cTwC+A5fPM1q891s9Am9u8hKRuMGcv
nlHn5dPbH4VtTHB8GNW9hOq5Vg+NZMZklcYuKflz8qP7sZMmUVAO6PugZOguFxcP
4M/PTFhGLeQG8LfJfhIO1yukXaI9IdzGn/h03ZhYwRoHdPk6evXE3I2ZHA84TmYP
muztnsDrXHZ05kRA0rmrF7xy+otqRuseBS5BqsH88FY/m9NPtDTcVXDyGSsefPSe
Z2Z8BYpv3s/igNN/nRJ4Jx++m9KdtqMU2JCHKXEjreCisDKPI/SUoyoOm1D01/ON
mX9O2FGKB/lmXNuxrCx9h/qcdnjxyMBnROzwrN+KT+t3a+cYs9jaYm5UR35ovqHP
b4odLszI4Yhz8GwPNG+ZCxKF/eFeNzzndIiA8OLRc6mD4P/3ScSZC6eiWP+M3y2z
yF5YT1T0JuC+x5/3sLRaXzTEEPxDyadj7FfndXgVxRFf+NEIBJEd4024cENjlp5g
Xrbdlbk2AsXehZR9uaWxMCBpznXjAQdzInjhQrFo6DIxW6jsSltqWYxIIQSFTcfE
SKFvPOGsRfXBfdL9loThOFbBeCLG2pgtDI7KwCkJci+PX4N4Gjh/K7+7IVeIILYB
yVb58t9l5AJENeBpdO9yhsZUwEBNBoD7VpvQfXC87vVVuiJXQY76v3MetF3poy+/
6o2DDGRZYXwNhazA2II4NyzMgIIjQP257kew0dGX79YbKWs19DB2tP8cplOOVje1
EFSEY6VfIlypGcxHIrKISk+N9HDVfwBvzYrgXEaqBlKaGW9GwIocPgfExljnbBih
dAQ58IuYutGjaC9Se7iwvoemVB60DmLWPrGukToyCEWRvZsna7nUYEHFFnEOCMZa
vg4dV4aBXzaLBgjv7/ZnwuYuuxCnDjm2H42IjkIKgEtcFZ/7EGwG+bs0xXN7qhV7
uDd8Gt7kwfDigdgiHPU0jqLcSNol5ElUUTJxjG0Eb/hemEaOKWqLuLKPHBk8vS32
UIiMT1A5n09YdP3xiNicxZCxlRf/Sm5G2Lia4oGO0TvJUlb7Zo/LttMDLuDWcsS/
++WpCjVjzCdg++NW9LrthiEPfgay1A/W0xcwDRSo8X6ba9VJEGSgcaT5HfMWfZib
csy/sP8oBHV0F4f3/0RvlSbKneTYCXQcXSnPguO9cDahzTXj/YQSrThwXCxNKegK
zIlw+mH11z2sDg9IwxkQASz2wQjiDxTkUY6NXUYYeqzsnyTL5DyszkZBbrQNh28o
7NSHckrntp4l5//5fPHY/t4X0q2kQklUTfzHtLItdKvTRG5fA0+kzAJqjh89DKoi
izGFb5mWqeFj5jY7suHMEVSI+fGzDRGseWnRwX5IK3T3HWebNTm20zU1HANvubSy
0VjbIWN4Tno0YEZBeoVHnwMOiQ5XTMl/oMbuCIOAcEdufkM10BsWbK31Sx2XfJ4P
LzEFjyTcbUslTugtec7L2AYCCQif58dwvPWHk3/cZ9wTg/VCANIkUJA4SUzymxFs
1DBHYRH0aBoFzTbM21voJ+lE9TZXkDkvg/sY4rrPmIQ8l0SegK9JyGvsieR3rl8A
5ALFzwbUqdvo2YOct4xl+Q8L/6Tjb6z3kpPBxVZ4F200jQaC34wku2b4tynGkkbm
DcHIk43bu8aI6WiUkS2NYECCYIwbTl8GCbTL5v3ZjgnXH1TO4jGF+bF2Rh8onwhr
Lk9NieCVI+xDjvODMbxw5Ys0CBFLYTbxE3iHZaqHub+yzW9jshVDybqw+zHU6FoW
QFTuhFUFUpaYIrf9Obvg+U9HI0+HJkJxz5dgQDtY//m2NwpjbRNkxQQSSLspehbn
/cuc6hHKuMGOHfWqVHJBLhNW5EPD+hxb3F09eeNqmBqMd1B0Rdlrs4p3HmX7FuU7
cxYMi2Mz273HcHSgaZN9QToJM1nJAYz0p0wU9ObWaglGLK3Fa3MaB5GYBj2LojtO
aZRRvhXOREvbKI3lVnOrycaePg0Zb3BbFr7aPt/TVUaLzw7aUnhfo98r4koC0a0o
UNsqIGfx7qUXhpQSG8DjFVCTUPd4Rnkxameyici8icJ/7FAy9Og198VeVgT6XFd5
KEpmaVHJlfz80dcDSoICBswIlbc3KsRsbC3hW7O/yal3RDm44/KEr5QqGmW59/i4
z2J+qClUgpNZvjvNoK/CXHOpxtL/a+uZ44rSC6JiALVtzK5iNOKvYrJkqTS0zsJ5
bk/HIwYxkd7s/GGl8vIFFjVXWAcROggO7DBLMNBT/RJpvWZrbc7Aii8f8eQcdHwm
azJqnBlni4uNgzgDC1HmbxeUAasU1kKPzA1glBfjs/SpWu1v33Dh2CyfuVlpv7RT
j9RGHZrVFKXtbZKtI4R9PCdC1Ub/nok32MdQyqV3cYYde4TDT4HzKmDhkFkc1zVB
w9EPMhKkXCM3QQcwrtGaJBU646ZGaWiZL96qfXhRO32XMTBC4aJRpXUX8nwNqQ1D
7fLzyEkSAqwGbfWLAn7krvREQdc4k423L1J2K1OX9vlq7+PbC7yYG8cR/CzKzAlw
MhotjTOLcRCVGBfJ7jIRkdUnryzQABUdYncuuFQlsHIkRJaDCGKfGfWJ/nntrReb
ZQjA3XWIuwLQDUfPYiT5pYpYLqgFo9c7NXhhwMfbuMDPlVG/5GRzTtrO/oXDwuAp
IRl0AG1pQdbtfjoZyr0BsVMSk45PMajwZMqdBzdTmmpbCAPHCpOR9kYzUXAsfwCc
IjbkiOm2wEwSJkrd3VAIkPdhQWJwKpiGmyEGEMc+VLSr4cuK+X46PUErmoC3TD3h
SX+ThSOVRbd4Kz3j9d5duIOivtzp5BhlPRdOzu8/Q5aVeqjJj82q7hXKdIwk3mcl
tY9nfCvobKE7xpqrEUYbMEqNVESY0MCf1qDvt0QEZR+il3SpEtTvmMOlaLPOnISo
IjuDtWE4eCfMXRBFxRnPP71ia1k0CsXd7X1f9scLa8T9wN8OrJTn4MhumITrySAM
xAMl8eP09BdDNH4H+2v6hBZ9KbS8TNuMSuo9xOfIFRLU1cajY4joBdk2qX1lq525
ZccJIw8tNQhbnyVCtcT7FPp/KCRdsS8HtY71zQMXKMaRTx971U0tdTPlekwfwq+4
V8OKyw3Hnls9NADIuVmg3OwQ1DTrjqbveUMjuIpLkYFhziYGs8qgiVoWWknjUCQ9
ltk3THO4vj2Qjgb9jdXAixjw5Uip3+rg0aneh9UqU7L7xzv/5G8MS8dHBCqiCZ7U
1+gJATSPFANqm3rhgF8aV3j4qDBiIjQcJJgdLlCoIT5FFn1f78AvCOLjFH8h6CBo
WNdwPWwlcZeYPZpycANS95fblk8a98d+6q9T8UYp0RgMbbKErLTqCKbYRhsRLgqa
v8jRVPA/CGOnM7u0QNLL0iuuBvewVCip3H8gjJ0kqzEw+Xb2V2R5Ky95ZaP8wUfb
7/HagNnGHz6R2Jannxm84WrfEPWmqP6Oqu19LA8Bcur5bPczkQw/DVsALx7lAQIm
BbpOJgV8AD/wthD7A1Q4OMVTe7Zk8dXlMpyhaUfckAKGyAIksrSvr0A43TtvBeHM
JDwP3ATF3RsO+7TTfTCqWm/g/k+hWEjCuJMWrYQn8LGemxwZl/UC5iTtaDVHOZgO
54bFv4jFnjrOzSx1XCp2qSP8AgUwjoM1pEqOJpPSD/ev64gDelAln0w6nWzwpOD3
YJEb8Mqkx+c9YSkz81Mb+L995ovcs1gZbljDmTpJKM/kWV4c3NOL/Yi72kxgRdne
r5U+Ov4G1OhgsDFu+0S+8D3cpd11XWsa7pKA0274udEjc3IAtI7z8ZYDASdPa2Bt
GCvlHZxzHGTwtnXG+m4lScjPIey0vXaGrCFCgJ+29dKm5qqMp5SU2bMd/7M84pdm
f8elfewHDfJSrmX/OGr73wW9kvRbc7xPat83rAtPvsC9LA5FCDV2yq1qot/XvfkT
wpZONGbUfRTtu2sYET0Qx6zTmltvOQ8n/Q546SrstXXmOQZro2ZJ8VbjzRPsxGRC
gLdxxi7tM3+FWbIpBB/tSOIHn54aWjMXdb7lJPzkh0dA39LrgycbmpYW9hPnWBlr
d+ejF593lNWhAZ8CpFtQ//6rZvnKY6C8ds91tpsuO08C1SFcmxUfuWYw8+HM90xE
3/jLG/KNW+owin4Dpw9xYoLkSj5p10unfUmu/I12/DoP5NcNdYLXVqhcmzj/ZCtR
PQOuhyoTiSGPCEdkmXxNmq11WW5PpZ3pooztU9WoWi1I/yeIQ8GSTwtWsmAJY+ZS
H6QATGtePz1jyA+KF1vIkYcbfK8ePQL6oKn1VtBY2um5+B+SSnGfLNKWFZqNwbIp
SGmnHNrjjI+gf1jfwkAR8rKblgBQ0q84zTkgG2GszT04A1JXlKs82NrmKY8netsY
5Ms32DaDS1VJm4OGYulu7zSfpMcF2VTWQIPRUTr18eHGBE+OiASLLwpA/pYkR9XV
19743dVflnAa7PkSshmCXbGHGTIqbBySisoFpeb1YVFY0LZ2boYTX44zvirURBls
EIlIHtmnCX+A092+9I5FW2YM4TuRnsK03HdREXyAnG8NvitrcfIomq7Du5TMeCYF
k45qBKBgp1/gW3m2RQkJhpSGNM0vGwvY1UBea7GGGm2io0YopHQXBb8JJj1KMKLs
3pM7cwhWwnEZIxt74HR9mbKTn62gZJ1pzJl7KeIOS2lLV196Uqv5iQO1Z8x6ItxO
oagQPBJnVF0tIEhy2uMX7EfqzAvqhLMbi+ib6sblMkndwsKOCWEvQNBwcMWL3Wac
S7lLlqTvQ++rnLezGx+x2+K7iqP+1O3qvW8+Tqm7OWTCc8GeO/gVpJpTGc3DxIoZ
Oq5q0NSu4XEEJPhYYAkIjYb5nfIjDGR3iFm7681PRYwK1vZGDEgSqY7RV2q+GXVY
kA3H7phyStf093G/k5P2fRty6o4gCAqRvh3MCdHAhSqW+rSir2NaCn5grJQwk+t+
iWKNnRZ7c0yVpAmCDlDbpDN4gsSPFIDwgwrolmTANZVvn+uBhJJ6Lq1RXjXu/6CP
P4V3um1MNcMIbrm6Du7f5OgzswpctTpqmCMAa5kaIlF4j5RyRX6sAiVgj6nhnyBz
V+QNa6auFEXg7aBvrMhepwKSpjoPhVP1IVtmniySMg+GYHyWP3eJBY9ivtjw3n9G
9dZPr64emiTOGrMxmnlIjELvnal9dxoRF9h1f79hAYis2DOnGTPipuqM0p2V6GYI
NKLQ3tUtK5mtRfadRHf0dCG+He3djCZ5iXS1jIQJc/OFL+U7iOUGIm3cNTGvBd/S
CY4zoZeXqvkIPdtMTIbYHlAX/00BZ10CRnO0GfRwWYHIyWCd1Gc9NZ31xzGI9yLJ
4FR9UCWnGt1M+Mn+iBPWceNojcq5d8Mr+Gbk9yTUm8xwlkhDBdDx/n6unx8aMEDo
IKjMIKmmBqXkXEnMpGqL0IiiFZEQkXexgt1QiiHv2RBJDWzB+FO7KQlIUVZJ5U/w
VmM+u0dLwHeujOBr+o5LTYgxim8QUvT2d6kq2HHlyq1RFeqeKgDyY2ixVBl1ExkZ
buDvDYmxQCBWnIAxcLPFBFHPfxsCllfW/W8VZgkfQxAQb0NL0tUK0Vczi0nZOYhK
0IfLAJpH01YMbI4eVOOzpzLIvf7cXLFMamfEFiXhEcvApSmiIw0yuvK+Rtsp+JR9
FrRQsSHm8Y4YfIXzUfPYnHERnA997hAQz7tCZJOqdJTkxCv5na2hWIu2wP/3imft
RQQeauUzkyFThOfyL1ivH45wAtjE6MGV8IWPYEJkSxX482XcyPDihi6pZjivJCnI
ro5JKGOddj9x+X9UOV+QstwcRhKjU7EIzH39egUTMv8f+StYc7FGZ6JJ0hGihhIV
+uW7X3F03dKnzFyL9FrBFQe9snRjuKuf+1AchCtTrcdnDjVNeVy34BtQLlDi1uec
O6CX/IjK0wxracjnGQsAX5eCg1PqunUi1KqC4ZdCV3LYQQInRyIuDoCqV6sYQiQh
CulTZBdOCYYEkYWOgdAfc8ecQAwxagEcwwA8SNTzVkzJhSFmXys9hoR3xbofu9d/
LANXk4egNPhaXqjg+X/zN5EKeGb1DyVciCNhF8U1ePIPkKvwpIeqV4S65U4JXi4f
gNDtOBkZEToX2wTK5tRh0zRFDu1UsNI7yrMYuBM9e3gsVLNumFT2PIewXwbsd862
ABCh9tNjPRQzBjkARuhjuYO5mBA755atOdZ5u/BZTNo2lJzucDfUVzPLcjg1FV+b
szo5spL55KyZmWcrKmgtTPENk6Vz678IdSuymtbeGM8cRYIdZ8Ogt9zcPyKswvPF
cUCo9SjNpy7keQSlkMtLMTe57e9jwu8ZgihQk/dvWJVzQVDodUIZx3L0gz96vI9u
hPm603P67OXU6NP4I7M1PQ1HaOT4fq1qx9C+KWvHlRvpOsmlqSs5JFndkTW0XCHd
EetoGzuPpxCvxEpaPAOGb/URhV1VJ9sRWS1SQhrDPpxu79xwkJQ1eIi6ZtsCsq+r
A9rUiwyVE+2LeTQ7HxQaIOMBF2eo4PnQy2ikufZ+SdQUVonzD2yM3jZvbe8XCX72
+e7GDQcuRNAVNZZiWuuGeW7FXoZe6bqbIPMshtixoaraRbiIpL3u5RatxxyHSkFF
EiH8nZ8NDf4hb3McYa4S7M72rGWcaPCUYfsRkaBQnICpZ2fLVAurVEPGepmNE9y6
0u6BJ/lSXiPKZK4m87OKZ+VuC4sWpxHbljewDs6IfzV03voTQTAq+Aw/e5GDrvMp
qBATUdgIzNhqWPLt6jECsu/D2lL+yzcws0Sqk1aoJ/nblThTvfoud6xXWJGY0pdW
bVqX5A41VUs18Fv3rJ0QSOF5hB4EPOVKqZ+KtKC0QZdIwS9Ud1N4E+iBpByayMuL
bR7gJVobRMwnXw8Lzu36byG+JW4BdKfAw5bHrdC01StM6GjvJmdODnD+QRxMZWd6
p54FVpXq43ARnd+eTiS2iNf9SpVcmyodiKfQhlj/v8WbnjRUs4Fi3taUfSTWRmyz
mmXIZg45fbnnJPtLfAv0RBNLRKtkiwVqWNNDnL/VUfx9baVGXPg9Asq+JCvsOj3T
XUpCDTbPUkL6vV8Pp4ZUUOWqBqGzf09JocXI88RpFnjB4ow8RCSHU9epyb/Y+el0
pFcxjF0ZHQ4C5FAgG5VV+gqMoU+hALfK4iZ8wjjieXd3aPHch/4X2Y0nVxRXAJDs
sikmmcyfAX2JEZmrX8K7K1bCQbHmBPxwW7PX0DJMhQoOomGlt8CTKdpwau0A83SE
XiyAWRXkecX+daBPRLq2qcXUv5owBXXPyCUokPR76RB0+pg836E+Xd/9Tc30ajsj
P2zra+oONaWnKGIkxUa19MKnMR2BvFz+EnHYRMtcIJgVuSVRhlJz2f3T/5qEPCf2
RaDf/AHW/KlfHUV5DavPxRlK06/DM4Xu/UoKMuGtOvicHEsEk4BJhTIpsbjvExdu
k0Vkyu+hJ5iYOgWi4/BX7p4yNFf1QsFqj5kkW6pUw9Bk+3L0Kj8tITLkIarKtIhw
v35ZqImavW7NGH6A0prPUzNul33homFTvWZNO3ZolPVz6BYds/e5QhIOiwYkLWEi
hnRoc05scpHFPC1jCwANmLQScP4vn3nWd6tQhYjPSs/JCY8GG2ZOW58im0A/LGm5
pUGUbyfXEN9vSz4jVbvo5rSBHPErqwj1FYk9z/cZtQfF1SyC/A+XQZ/y8HuOuy0U
+AYPMwEl7tDWkB6CRy+Ix8DAmWX0McRXKyPHhNpE2w25Bcwck28UHm9qDYzuYlGx
2ZAQMD/GZRKIheS9vpj7UtKvgXZTFn6ObJ1lySaQlby9WKgoOge8VXu/YG5qYFxY
xj3U/zSRiHSvSlcZW9x5P5t17Hd1fOsWHA+tIo4vXwgcTCeFb1Lf1jbgn3jiz7Wb
+xYNwZIM1Cec+fFq55oySWFUFchqr5tdYjSWnJ4Qpb+dDpDoxZQTFVwcFifCBcc+
SB1EP786dmKA6HxYmLqrl9JAHCRwprOD339WGvXOJi1LZ2U6ZQI/ZS2pL4tWaqB/
GsWDRQyGhK9JhNnFfAwxGNCjXS30Ez10bAayUu0WTwZ272/l1EiSf6rMutrijIIa
A9OYoceAo/uQDyRYxJWqIhmFEUNfHppmvVLnogFdlHs+4rvZzCXmaD3PgmPKFTeU
3T1nko9+O2xwzU1j+zqWRZe5FW2zC2GX4whXjkhGDayTa7AjwoHv591FyYBjJN/u
OEFmQPbsky0jkVVZUE3n4JwRcdXeSQEpU0bJCPTK3k+f+em/gTOqh0/haYt1FJRO
D8m6xiUvk3ruUnFIAV8Hpqmr8NyGgo6bOMO1/ifHulFhdz6tIxbSKhpqUiGnLZ24
iriWGoCr6vQU0YUIAOJCfuUVIps1mUXrbAiuMhVTAOgtdmQpVQN4UYWGMD08wvsW
O6CBMjH8X9UIm1EoHi1oX2mhQGb0jYydnIG8qT+NZwP4YAJvJnbgSfs3bIEYOhBT
G0s4kpPhQZKZ/zaLNaZq2FkjA15E02MTz7xJbLONE6Fe70H7FE4nFGX7msOq8jXT
UGnnfiM4XxsjgavkpfYcIFW7hB/SFH32HxtfYbcp7RyatdWBf8/Jv2tCLHq2rvAT
QiEO6zsx+CWpHUf3Rwz3HeX0L8SLumaCvDoZH2X/tomrdM0sCzn1m0LZuWUzh+XK
tAT1VtxYE6KW91ptJT8hcT1kzma0RmzCRwnpVVB7ldDVHrGLsLefs6CKZlFybXoq
9ct0VTrWuL3uq4A727YXOMPh8eIoCzx22iLfadKsrm6iPP5f/K+MgyXIRLx0pO4Z
icRpo0rDFRJqx0Rf4+ugQLiD87JLDqWqCJurYcdah5WRgoh9A+1dso7Kp0E7rmHv
LvGo96CJCqn3imElG4lql29+6so2Uaxb6oJSbIBU3M9HWoMqI4MWi3RlaaPdAT22
RKu6zCHQC/Bh4f/yif+P9kCuo+1jofx4AydWtM2gU5ezTIDe8bDFWs/KuLO4pqRz
KHyeRss68yhH23ffnUGZw87IZWXceoN3eSssg7CnsfM/4enUKp1KDgvYA9M/npYf
b4AsBUQW4Hr1r7k8F4EbcDC49cQU6uCAsl5pdSyq0iwe2fkSK9+deEjL0ckeTYEw
fY9hqr2ClRVPbRgTNGPnfL7c2n1omlZHmcDVq1b0hs3rlKwgNI981Bq9uKEHLJ1y
FVsu9IZROKxLJE9WOGyOWsOfpVcltEUm7Zov08eDDhqnBPG2YbxI2M4GnyUwpLUX
uA64iJIzf4WF2PwMNr5S9lo9hoRbzihctJDjLWi8uLI9IC3dlMPV9nhQVnkMxGs9
AjyC4EHwff92jAIx1StomMJcUUrlZc5dnAh2ZKYmP/D+jN1EefULIhoXmT67UWlo
eFGlDtFb0D6HfGsrVCtv/X5OBc5NV122FR3a7uqDd+goJMcz92HWZ4A6OwBwFb1I
+eFmwg0nMoXf9Ju00dHfQiacA54X4jQgNpHchZ/73m2dYcUZ1fqdGA9xGjWm0ksO
QO6SUTgCfgeVlpRNniBki6ImfCfGvAXxPwcTOg0I/4Az5cbX9hxJ+oLvhADVGfT1
3umtWQCRBFNjQPXSTlYAk69u34YcyYBDa5HC/pgvlpDjayvOI06d1dTOYaPS6Tse
RopJh3JXV7eA9mpUr9QzXPNmOQ4xC69QvZ7bQlGLdSsNcw39Jpg4ju5/LWyOaod7
J8uozVtO4qnbIxVdANpTKbGiOkMgja/MaNN0Go4s+HAvE1XM8Q6TOeEBkY7SAso9
/u07REMaoufnUM7Ae4LheOCVs0WCJySa3LthsskWw7dCiYFtFPtdOaMHZA0Z49cM
dDiK6uToKfo1ZZ9pMd8sNDzCCM0fOLN+auG7Dxv+OkHU6uAKYFitaj658u2s7P2/
prgaheE56XJ7icHh9BaxxdftXo8Xc3MZsMeb0hDqDdFBWaf4DnYr086bOn915Keu
Ox79i59Dqldt+iyUmIA7EYplFOYOWXJlppcVm1E4NqKCbuhXUsWB5sZ43KRpBkQN
FdbqgQOiYXqpIXS2QmPfdu1iykUBcbDMSq7EcQHDeUKQ70g4sR8YbYCQZJaZze4C
uQk+0WOFW0j8FcVHZmVaWcs2VRvZd1tFzqsGWMXITxGSameF6FIbIgQv6e41FWko
5tI1PSCLujvjJQfyUoQhUYOgflt7LcPFNuQF91x2no297M9a4aphhGRvx81IUuZ8
bAepMmUQqL63c++renfPcMUzHg2xCJWjb94ZqjX8+jEM3zDB6S4vbyiWf1166moP
kSYqqXmLmZlD5kH69Ic84vK7TdXHCuSoIvlMN4JFoGKyXZXbO5LqZ2FgRJRTPZL2
07WmsMc9PMHmb8TL1i2mTxUbW1Asz5NyR6wd6jr1r+kAjFB8ftqunkTq2rxdoLFW
LrxDr2IrVLhY04Bq7tPJOCEsWGVgG6Yva3lS5H7s2s36d8Qds90pwdWLf0Oqfd7L
PSXNKgT8bWJ7P1fJeVtnse/iCICzLBz1oAutWvfMZ1W1uZ1MkV7eoW6D4g5aUdFc
gB3C9xyNMqwdDnxAchIHkPs/jik7nM06AMMF7PXG1hRoZZuz1wAhY7d/OuPvdKX5
Tmk3yTq2D8Htm8BdG9HN3AjJnFTkUwwitbPHUxQXGsm9IeeEL1J5LffEwSSfqTi0
6Ax8FhMQg6wLYYhVKRwvUL0QM8UIDwIno4PTalW4MtZqTABFcvjt65ucWzWd7DQQ
Is5a1h+unnLFs8+UDKp1/5LmRsm4hn94O4FRiLvAA7Fbr7vY8EGM6qtZTv6o8Pa2
8HdWTFhgCEY/mWg3UBqBfIs4d+maq33W/Fgo37L9RK+oF3hJ7X42ua8NpaOgRPFj
GuBfSsldfQuekR8I/+mW8LCAjZLDNhmvCT5RRH41L3iRmawPeslazAJ4mKvxtDpS
CxT+qX/lG+/qhTHy2hKHbzVbDYjyzGvvBv1UP0IGtzXJNqLlgbcIVBcFv0KJGOb5
4Fjqsn5b3C2t6Q+K/QZ+v4qm4h9SghcnoPGeqIEqMM6tg64bzdrlDkbEwIEUxWiI
FoNMdY+xExRwBeAE4Fpqt2YQ7yPx/MfErFBIkjCCUmWGnfgqeyRvPhG7Q8hdr3Az
zR6cnaI1YKIYoUNnQgIJZPBGWz32SSuZC8EbdDkpID8BzuBpFXZmfv9O4zeSKK4i
fqvvVxetb6yQJFRV4LskLrZ0M6uotOPFXRSP3axs/OQcyN/f6f/n/HUA7RaoL21y
OBqAxaULvVI8JslpmxqED7ABC3Oje7ZqbUyflPUBIewd/4cfnPSx2suUF/+8tnyU
7kDc0yWj0rhCSYxqpZAdEfiWM/O5hd/IhFcefDTRhAHPawwWCFFKigyzMbgQJ5bQ
i3725xKmYfwmg851F9xWTuVo/FdTXFXfZHs7ddm1JXkV+I9xm4v8gFwAWs8AGCsI
L/IyldujINwUQjv/fYYT+Oi5yIhWfGmwHRQ9JHhPoXU+ywz2CjV252bJWKlgagop
Lkr0knCRLqJ2CVaikRGzQs5gt8cDNWppl0UjBMFzB1tnAUdedXfyZEdW4Ls2oO+v
Pi8nWoGweve5oEThY3Sn14JEfeMKx8kihdxgdZduVdH3JroCn2DtvULODw26PyQF
aQyOogE+3ArBmk5fZJMt0bskRt2PE/N7fvOr+RzWuUDGiy1KQa/AIGkEXJCcoEcb
mKckHcKJTA27WLxUMK8/BjcuO9mBoQnBMGTjlacet8LqlEfswxFIsJ60/djlHkNZ
TytYvKJ7OYen778n7Xol7aFTIQlqRRy7K+Q+8+lGahMPf31ObRdx6V83GmxEom9p
Bx+eyVTfkj3Ri20RzHvwQgHRthaO7n0DFhlaazLXaHZIGjsojPk1d4PFtuTPwMv1
roU6wVFT0WZtoEoAPKtu3UGIE8oHvQDc8ntNpxsGa+oQPJdkdbC7e6pK5WVWOyqa
g7U9xesRgluarrSU1MR3ZCR0uBpg413YCefErxOMwFvlmlWHHMHCnWvVlkwwzW2V
AdT0np2Ak35uC+NbnovllRa2MZ3vYTXknb+P2ho70/J6T9XdJuJg/U+nYc9+k7aR
CKrA1bmC7Zr6zCqhrBYtPDibuHA1sO3mmIcUnE7B2OyUwq1EFvD1Dm9GXXSc43jU
QWGztC3bt3538G9Hc9760ZAjqLToZ9VLB59PgLd7VT/my0v8FIdvCQvl3vixu61i
zP4lR57utlS9gYXXGV88V4g+67HF+rC/rfK1qyrpOJ1qVfabv8Mlntr4b+X2R5d9
y6MHUv/rGOBCN2D4NxDAfxJREjQoCDBB/wcbcsaC5Z+pRIsVCI5c0tNhd3QNMpwS
vQXEpLIEv4DBf04t/UJpfyAVcKBxosZ11KEmJtoUvkMJ9qWV7mARIf6Gx6OugXo2
t2sP9stsAHu3PbJjXGVCZp/v4RRmN51lUnlDF8pfGgmmddlqR0OItaplvk6EV8+l
ACIcBN4HUjuJ9Z6rUJ782J/RJFRR5yxAWdQjONOrXvmDb8RZFcIuJkRMPHxe1Q+m
t2IHlblb+pkNrKy+NQAcv14qa57JwmefGPg88/cFUwW4mSJT/0KSd8LYqqGx8XRA
dE7w5oVd5kdU6xbyKGVn4RzqsmgFjrn/oE8dLU4DK9sZx8+4UYlRZt77HeYg2FgW
OZPiOw/8FwWDknf2QRQNhCg/A1b2itZ+9mmYJjL3Vx222K06orpVsBUxXPfVtwAz
lnURLlPXkiD5tPpy1DJsyPyuvGQkGA+O0zLWOsIKh0HS1HVkmrDiSudW9JOgzd3G
iWE1ac5yP2nbkxrwjGf02FaYLLJnC/WYhGoV/mQGUMV3W7WOUIf8HrDhgvqHICcD
FZkqqEtZn3J0JGW5vwt75XYZigsZCXQkxazLcdbcyPsNofxBLVoaU7Fi+2Z/IZj3
OOm58DwBrfGJh/0bJE3uN2ITf+UGag60nFIVREMgYwPnKaz30ACc9uu9fagMRpOS
WFhmr5Fs08Iy22iE3Q5G+eAxn2fhbAnuek1+2J5X9JYBl6yl9Mi/quvwFhPUoMqS
0Opcu3gNFh4PRxlxz7vnhc5FA7/++eoz8QWV/IpfV9RBPxVZgWVCsaCT2MNpwf7z
W27vsO7FVkILCZIbV2C3J14q0/7eOuBAgsUdgIy9B8XJpapECvu6VOqJJzJAcuKO
FuXLt0RQxKjxcphTL/9zhuaMcjH4uJ26KKEUPKHHL9USDygw1BUf5wZzgVl3sw4j
YU0nPDEiPPeyXqNRKxJUGPSbji9Elnk2mFyp7Ggv3xwU6pndp1BhGV/MEVn1cv7E
ClCQkKKd8abVc1fDpSu9E2ozSZTbg3mVa1I61Yam0snYqEnIW7MrfMbDPacuXG5q
0G/BG4xomtxWRsndKp0pgIuL4qGPdQ1w8Hdvst6UHygEDdCjbG03wjRaEHiDXf9w
4bJ+xjMcXVUMpHzSmLGM7KSS/IDOHVIWYhaaJE4jDSTNjSq6HHexKuLiebM01MNs
cddYakqmEmT8TShbdc0EhQpMj4LFMKS0BS1mTUV65qNRDdIH/TplcsjzHI9LCOtI
78mtx3nbobrhl7S4ienmhfyWiPRy+4R8rldNuYrRoAc7pbzFKoKyj1PfCDV7Mfmz
EuNcLiJDd6IGvhyRnp1Ctxt/2rgRmwCfVvuYz6BAUayKPTBhyN2K2PlYO/dnInuw
tWjPjS2olx2JBFbdZkWI69sIQT/oS7sVO2q8PxYvactsEffpnaiQaPBokpkSkg2w
QGcruVmSqMjXXmjzkK7o85wH5PRh3AQ+zpJJbZ6aZj8qfz+QDdBn1hfRXB3wVE4p
IxDwtcXUU15w8zjMqrHmn+Iom0X5H2OEjUSD8KNAFLjEFSQtyT7yxlq2V+DTNfsd
oyMClcUhUr1Dnq0z/Q4u9cuT9HsphtHH4OPxzHQEjwDA6kZUQbOazFBnm5HTU3RA
CfIoGZyExDh5u+uVgDCnkQzFyCpoLZUyeIQVfE1VQ+GjXRtOXuKwGcliTyCSDNgq
rQmorhTQ1ETN0AU1+JzXiHCAMfFV5SfQCLuCp24jTCj3A3kaahM70pl37/ObD9+M
jy6EX+UCDHH41tOmJsi6tzCNW1CFNWmHSkj/WyH2yOFlDWVoBLzAlvsHGAfKoTrR
v0m2H0tH1cIj2i4VFpr3tlAS4J2VIwl+MH/We3FhuOPLFny+bT4UnhOLZrULc6c1
1R/dpXE9x6LjpZkHeRtxYIgKHhnf6yQFCjqh/Tp8xjRzxHE3mfyjbH//jmsqlslU
Ff2BpjYQ+JffT0acib1EwLJ4tlpI/PO1385rQnoSP33KMdOlzS6dWUoSfbOTypLw
/mSQyxb8zPBTTSFGgSdW5XBep8RnAnXGt5mqpswVixL7kEdwhZRi9a+LRezth8gt
R0BtKWIzeMzC6lkqOjGtXgIJjdzccEaZJkmfZGwRuwjXdWqx5HOVETUg4tCZPj/8
8XZxxzMh8AGxzesaGZ+M01aQSJSbM5PGMD7+muzqlCGzmabJF8jc1KaBsGphxtKq
kaLRTLnaD+rLJk9e9OAxuT2bSrjBfcIlIltnyHlWi88Q8zaCWBxeOvtZI/HRtou6
enXnDwUawxMciEx3aC+ZgEPSbuwJL3RbQWXDQNMcQyuoaEncouZVOKLlw+8YsaaM
9oBvNRODq6E4DocmtewiVRsdWDnpDS6U9/bNIwkOZGQ47nQJ0H8zufkLRuZLuBuj
vpL3ycYgv4Gtnwgw+rxDkMeaRE9HXHQmEmvfdBvuTk5wdIEbqaGzRfV/qxeQewEh
fU8CMsgY+GrQcdJUa50KVIeGTQQ5QW2VaAXQGqGidzbxJosz55m7a2ThpZmlv0/b
4h307n/xnnoIqGERbEpVr7aqtn7mgZhKrBJ+t3w8nhPU68fjo/GtOI6ILDvGiUHH
F94wgLEC+78c3VKB821usbJPFKcqTVeAH6LYQWICXouy+9qWK1+lO2OPkgs9MeIk
fUTHRlluKG9qEAsxlSlKNDZJ2Jp09HEpxsqRE8smC0eI8765S9y72q7i5acC/Yes
uYKReOiXS9vVNGeHAzbHV4E0FFUOM2ONPpt3WWFx2THriUN5uKNdBDZl+IO+FwpG
HCyFurn7FcFNOYk/qdVpSNcu4qxicJJFrzjVtfw1k3XtazIYSYFyxZBECfL6BW0d
mf2/mcC+9zt8m5+quGk3KgVlgabKaju5UwIX5uHQa4oXoMtJwbiA20dH2ozQq9Pf
OYouBkWlttJ8bvAumNKHlR9hmULLRa6zyvJ+p0pEfJwSHX+NPeAPc6qTaXGsfV9f
n4rCTK3lS6yuSjd2Pqkrs5kw5F3JBWYs6uo1sL0MhWetuNsancLOUg08VE67Mekv
8RfoLjCxQCj/Smdwl8oIvSQnXHDfcHDX4UwWhtzGPmkh8dqEVliXN3RM/GHSwAQW
8k+uh3G0GOtThQsO3gfGf2A6bDlW2FRMxSa5o047nnd2ATsp60vF/DNMmXMVOGVG
PRaHuW7+u46HVKuXXxuKWhTvpJ9ECqFpuOnjfLuzJbGc9rw7tMRmU2qeUWsiOIB5
jGyPJyhfOvLA5/RlFk3Os2sTucZogS1x/ixwq8OI97oXRuMHzbmNYQupcXbPqvYV
mIvYfcmhs51Kjz40YvXzD6ZpZ5y34CgQPEE+wfyBP734JOcIZrItq+imkV2MOLBq
0z9n29Cl6bN2A+GbkAzn+sO3C6NGYv9/YVa+71eJ4MTeF3LJTyEqnCNV/UyEdoTK
laFeTULLx7IZMDSQFlWZZzIvEgbgPRVrGDM5iPtUpSH1eq1easw5cgyyfPjgQQYR
w+H/cvbhAq9+KzkXVWp8uinkQDCPL0mebYWrqJDzZGXEGzs/vqHWvBu6p0DNpe0Q
WrDRr3gXj+iKB/kN4K7KfbLv8rahwpJQwKIU8Et20M20qCw92/Rx/CYPua6pCGC3
Te4LtQ7H5OBjQzEcGfgeQ4Qm6Atjf6/4pbXAWEFbGSDtcxxMWxKusXKbMUf/tU+h
THExT+LJpia95rvQB5ROT0ENWs6/JmWQc1RU6wJ26jWPkL2fzaOMt4K9uUFAgZNW
002r7q7+R3+/1LzuGHqivUa7CnIQKPZQjtBsWhBd0zyuHSmTFII5obwATey4Vrp5
T509JYmZpUPU23qCLpUa3rF3/9mKlS2TnelxkGu/u4Zbwo8gBOpAYYcIqhXI0Gg7
xpQ5ENMv5NihkUvObjMHnuEuVAk/bzHObI0h0nCKDXDNirKmyj8v3SSvoPk1334b
dSTHHKuxFMae/cnoqr9IYiNCbnWxvp0hWfkRZMNji2+jVLRAff8g0gHIBxel5mfP
6oiSFTJuiqglkr9kiW8JICj3qU9UCWYTUpAqgwtHGvweRsdz6k3dkERo+9JBdhvz
rDrbfmwf9dNQeqFUHtQecl2BM58JkxQHfvpTxGxXM2lZkJDwOO49ln7sqxNgx9NA
u/TVwi+ntm3TxVXSQbR49IU5308w0prI0U6jSXz9reW0YtK5uFv5w2VemRhP5k04
OBp8SYj0wwEOsl5R1ZYEUjYmBiZFmINE9vI+s6PZFXUgVDm7tqQY8tx7tXN3UHq/
s6/JDJdIoPfwne2wv0Qvb2slp1xPgrzMuwky7EW8Fmp2XKDiFxgy9upjQQyUBCrT
jdXbF8kyUBorIUEz1o4XUwz4I3nsAS9ncQJXkJlqb0vV0AphE+wd83FYjws5Thdz
/8v8uiQ56BjCJqjZqdxI2pcEwJwSsFubIsD1rLqAxqr+lxSdvZrNIlyyBa+GmVXS
mQ9+TJItkp47gkBQd9fFe9C2pT886q301cn8AxcL7cOpYPqEfYX1JjAYeIU62JYM
8icT8m94gl6KWqHCCmpVwbSY+A/ducMrrlCZ8KvhVkgGawT0sp3fIhxaZ+YyHKX8
MoR2IhV6ZeeW1EuLTHq+5WrOQb373INRylguYtFSYJA09qAiqDyiKcTjNFKaVTXd
RR4E4fhyWkWmGeh6LocVFlznLsovcPwOW+yhJqXlbStimBeeSDTQM4e7NYBhr3ws
t7QGE4mITXer9NlOmDHKlHBfI3e3eAU+uf3okXN3Hg0F8AIq6feQD/ImvGYD0kUP
Av8gi9C2hrEtOmDQf6cL0oqGz0rsne45K0tRFW3biszC8aJorNschm40TsoeyO0P
baHpNDgLKR0GATz/c7Xot94kWdxFq7+H5Xjroe3VwwEXb024rBovUal4x9IhON/n
kvVBbae/iWSZ59on25QGNUgtUjHe1l3+A1/rJ7JLlJs0XhnbQ5sn80/SRLDadrqx
DGl+L88wxrtlR3WY6i/p5Gvrw/DmjibCTD3k/IjKsVY2HgnQRqE/LnvP59YpyfZW
80uo1yDXkISeQaO763SfLlAsutHwEgKt2C2xombvESWuEHp2ySmPc8IJ5DcNZikG
UXXIjEIv1Wze7nMeBbZ8+yYxsw/47v8DoSXA2hXKDxPnVogpH8KeIgAUyOO0buLs
BosWo30XALI/UkFDfCNdEVekMC4b/CIAb7l6kmcgEPfpe1YulmSgw1HdQnvcZfj5
n9j86OV92abgIqfl+a1sM/xrNlYV9qVu7cluvGi7lp36RsOKpZKdS3PCPvsizpmQ
NR6Vp2F4E/fxkpLpx58DSjpCaXDJCUCyTouJlVpRiCMU47zhHO3zd9cRmFx2gaYe
wUFDWjWboS8a7ku9DbFn2GdC9zW78jFn0dgIAuQ+/GwPraGPqLLqUPpzIaLtWwir
k9g7UIU0xhLXNOfUBTwSgg4ktQEOrVSpZ2VVpDUtxXFCS37zmJFuIb8fnhBr1WUW
+a3YjCXj7W0nYWVPOi3U5OYHl6uIp8NaJdlURGsOfjRqhcDyb0ozw3l4i/iHbuu8
ZA4e/HIWh5+K01pCoo8Qeaaz7heHdxjQkiWBRYRyQImYR4PdDN8yHrrdRhCuZFsC
V+7zq2z4rD6BJvjmNHP1GQVhShwceoUuNdv9zBAw9UupiC9oTTR3S2OkQB8Enlob
yQt6P0OnAd5cWPw0jc4UKccJiH0DbfzbyFE/oj0OK4rFTBIvjvfexJ7FjySt7obH
ljD4vD3ppow6eFc7fibwsAgo4zv2pYioBwYT7bJ03VhE9r2xC7tHM/EYLAGlKgOL
W8Cfr5uC168W9fUFra93iWAnmN5Ay6HSyXlLVoAyUojAobOPYnT2psQgdO3rmtna
uNR/jvDe+jPENTUwRT54bme73zbr34kf4jVqsJa2tudUdZ7NJNvWrRP5jO29DecN
6OY79qgRK8sU+cdW9T3McCtRGHgEqxaI1rYWkcedsxJ3r9vqDE0Ii7WW6KcbKw+N
1KyhSKzH63YorX3qPgLiiRU0mci2lSHKdjWvrugWkSkMjXH8L5X/E5QXgIOHc4lF
FDWDmPPoNt23tyuEpCRsMWaROfVRv5dIgjC3waUNaipGpAaWKr6L8EgUjJqye2Wo
gg+X+I1onqEPC5WFC/Kw+Cgws5p7SORqANjBuAEb6a1rFRpQMz9ugGO7y2VfEdPW
5XxNh40NjSEDLsRA9kUC0vjRXMFzp1aatwd6tyZfyL3D+YB0yhqgTbc/zoG3dK91
1FaCK/dcoly6pezpVjAfPWhOAh/j7fXWm6fUaO8axnGNL08MAQrNWL7FgHgbFbps
L7FUBj0ZP/oSwh02B55WhYQbu4JibcwUR+byxidRXx65cOiruQO36oGTBTb3kHsz
niNYKFvovBQqpNiPBXFVYZzIQJ2NQhqyBf1A71dRTGkGvSBihVyoxLwrYrLG24Kx
p/G/0sPt3J0Zlt2autkAh+1Y+UmTCebpiirFDXBD9f/qBV5Oh+0CNnt4zxng/5yJ
0RwvbojezhXelTBMRANHcpPqVNnoTfRPJBQg3qHwldtM3WOXgm0i8bOKSVxH2jpW
QEVa3ME6L1WZCCDpBR/RHOvpV2RyEUveYwB9CR+E5vn6PUiQluUdNHrKAKfNxLdc
hOKxxVvh/C88sFX88cSbDQPrOhGsb4pMIk0F3IrEvwBmMhfHrAm62fzwgsIgmwqy
wyOgLukzjzp75Pci/7OpGPyrFG/ANtAKHICVl7IQSDndrDzhbQS1daux55J6iIpx
OXpwLdGDkOZ0cgLMcFVBllOumIKtWqZ/bRmqsvB67zZaRppo92I0ztROU3c1UgK6
+h/aUV/2UuZnFhDnwkYk5Ho/9WNbNkvIZsZFdQYRjpBA2k0Gqa2ecOAc7Zg4x2KN
LUDC9IEi8pZj6tNFoKb0sOnk/tHNpQAkr0NEugQFCe3FziZ2QDwOVu3VhrKVDm6J
GHRpELUpkmpZEGLgOW7TesfeRT23ViEJpb4Mw99Sh1LAM89E3oQRthC+vq2phfdj
1UHuFsVAyKTThNYPJZgU+THvwf3HlG9DM3SITRpYuwqspDadY5SrPfHMMXkgD3mJ
fylu6AzNLqVylSg5Dpi/kG4JXeRASekeftRJeuvKVujK66l+zprKAXV3B7Ap/vDh
lGa6CWKcFrqVRrV2CluicjRI7YHRXKMr//heQSg0w+1bG1sgtNlowsIytqL7D4G7
mj84V5L3skaiiQXNy9pQcbhqe8zULoYY+RvzevY129izttzv7xY+jHAkYsv+w6je
Rum7E6SuWd6BVawLgVxbuuqaOqkrtf41QXs2HUzf1bkyshf5FLlCYzud1hRKmETb
plxkBfO6qoVMFLtf7KPQfd5fp4pZJtpECH5DzDsCUJD5kcKFD0+a/FJGdvz1Gowr
nPrZs/50xWEgCiEuldgDuSwqmcbesxRfgUm9PFN4Q7UDZhxYgbcaKclHthGgRBsf
vQgZpoTiHl+Uugir5VxV6wFhpZdUvdpAmbRtLxPiH2TlhndozyvgZeNSgtjDwN8Y
iDfXAPXvtmJzGErlzNB2yDl8XAAKX/sKcw3OW6GnpJ1GDoIFD5C+clS6nNFHOBqL
GNqh1PxbDFit2oCIRwfNgJcs2JAi0/za6L5gfBYH5ne5xKTR4fc0JP4DKHBDBjbX
AtdNwXYHJ6i/6EvdGo0Lye1N3vP9Jvfs0gywHhHyunR0qvM6ckiCB2GovYLKNXEi
AKdEJX/mMLElIEGMw8zm6jtU1b0tEexEVAiUlWa3OQpzNBCuyh91XkKDNSKHJE5D
xPyrxLZN2lEH17cqkPLKcplc317N4GC9h3h/rqSajKEh/b/hE33ri85nPDYsseSU
zPbR1Zjkd1muPv3n4pGEkEh64CYlGZIXyDG/VPSc6sAPxgsicJPbrq5ZXhILNcn+
PNDG4Ixj/PuIzVikiMuRGwcmqiviElmivEud9ZLWJZRcDKkPqjlyuZzrl+PX9/K0
eNvZ7/3EjY5jFSeUzcGLXbAYNR7OsVFZUXQIKs4AmOwy7/qMA0jQ5sMSxcUQVXq/
7Cjam45Z+PBNseSxXMtpr76mzEpwf6qH4uVC5CNkCQj09utqQirOvUoC/FDLWm+x
v7hJV7K2AUPfNGDCSMZIptwv38JbosJOIlQ5ji6pW+3rNhUvSWNNxn6wHTVJbtoP
g+2LdR6iHpdUsKCQd3v8jdRJZA+jG5BRZAkeO4bGNOqe/G0M824uto2F4NfUvtmX
ZI1bT508cSvs7ExNDzuIAPdfO7jZJv5ElO2tBcAOhN3qP4BZyXsYgXBuHz1ri0Fb
974kKEvCQkumHtBdfyGXZRllIAd4nFH6P80IHmIcypGPt9iKkosXO7Df8XLFQwNA
GI0qc/v1hoBDFIVZvc4mXQEBW8szJejYoVhIiOhY1k814ule0KC5k33dMSIpDMSe
lUoyy7oOGLIlQ9XY4SWHL5Dkt3gIs2Jh3tDck9rqlAolLz0ByxHxk7YSGgCEW/3N
9g8YVLx+Or+fWFrfKINhbm6mOyHsBaAiI/AGkJe/IcFLcFlfuWhvZmWqgJLjsZ05
9XnXKLLYxqlF6Oow8IABLDpDO2pA5hxiE6pMAec14KrQEK2PP18sTi8OvJHcRz2z
nDTnFAPBRJ7mgcVhjkfUEoKAOI82a3lCeMvx6Su9/4aSIKlIgjzAP66QSpbkG4I7
P14/2xkPliJEKSKKGkRlhOhDZ+y+b7YaADZ30vSgyzrgLoIpCs79pEm8kqSHsIn9
KUp4aYXNFMitD8WhZZpmeKdIq0V8ioWKBhOAJ6CMH/p5dB8sayBu3lZkwkBRKsZH
lr+p1d0Zb1EtVzt5QtmAi46whMDhnZiPxSO3BEcP7tYprIEVFbmqjLHysiMhNFLN
7i3wDT1qYR55AgibEjZG4UG5ndSihhdw0PSGXsoNZFMfk/2GUYK4EUzwcuhYSqmi
dmhB6Vhx0qeiuMiIObxKs5sblexf9oEzMC7jpHj0xass/jdfluwqNCJVO/kiusiD
u/3G9wl3d9LM47yDYZkgXcsgEZ7pYNVFZ7bB5nk1NddhTPQESkMwQ0C1/tYhRth5
WH0xQI2nzpk4Da24WA5M8PNw6BYB4MPUih6t/XM4pxkkEbHYQ2+NhCOK6cdAJ6Tu
+PefR5f4F4mOkfMra5Otyr+R99uGktfb0PU+GcmUhH9n9uyUX5uY4h9U4q6EdIOz
M0xjBaURVBrP7hpsPWKHsfhtBJzdcxmp4Dwq91R5J7HzzmW0cX0WcMTlZJs7Fzya
X8lBfsW2i2kpssWteAcSoRlFcSNTpjjNUzl2LR2sL2t72Q6k1HNpfbRF14l3h1Q6
DxNkqHVb4dpHmtm8B5ZRGWvqHh+a8Pzu71HV/N+ceCgMhea5Tb0fgkOYddcvIO89
xX5eLkkKXCK95krhzDVbK4k/yOCrqutfci45P7lS+Q89Sv9ioi8TOPrZg1qrDc8q
IcQDv2HnUVfxgzj2iKgQHRzbKS8ObpOY++aHCuZx6sQoOw9VoaTs3RbJCou78V8g
T1gxKnvaP9XUOhRLUAEhyacu/3Q/0JgJXXGvXvSlD7f/MYmPYQC0nTv6vMQdNEvL
a/YczNaOXOJOr8miMCKH96FE0pi3DC6/VQ6j6r7/H01tlDmGGTdE6agEtvK1HALo
dR8OhC1g7RHOM64v1FkbH87ZnTpZsrfieWYVq6Vsmn9vzNggKpn5YaHgGG5yZ43m
GjczOWRLLLd0cpa7/UpCcvpb39xXA0CJWyehg/YkjbXqsvPiAcNciJivFqGlyJQj
soF5kzrJ1PYWKQ5fjmTODEtqZa5CU3LxTLOcC/jgfJ550ZOnljum8ItUjumqWQNY
X8RdwnubcN+XBbtA8fTFhea30TaVWwoswCPn5EbrUZQY1SKttiYsNBjyGGvL9Ztg
98ihJ1OH5+vovcVRNL3xGKVpuXscJSzuA3sd3KX2zVvNCeg3YqquL/9VowTuGlMC
hHf6C+fmrmwMXu0bEkhgqfSP+2ihxLOW5T6pQB6hVW/wVhOFmCgplWatRodCAX6D
tZ5MJ5Q9OiwkyRuundHmnCIPRdm29IbIvpwtSE+0kzq77JknbJlBIvJ2Y+9DTG8I
xJg7/w6W9TIe5tUByCkvsP3fpkjfBALQG24Kujdi5NbyipoiMOMaEh1WlwHXLCus
seiWTtTKrGMt2O6wAC6CajMCQDEtCcWpHL5vAIxKgGaZriKBoUagGVAVSK/hgeOg
oWT2PwP99bJaPz+iavDiUNzEebq/R7XyzuV62mzSRmJoGxTS7aUmB8jpza9GV9Q4
1RPgDlvRQfmBSvUAil9bkhMFo4yIs6wcShbIX8UEqCIRicclJJ24tN+liknUmoGY
fRcqkBDzndVwAzfBDqo+JYB8pwyKJ4cz/fhy78ecUyuF8hofU/UE3go2z5/i5/iy
IYGoma6JZ3zas+2UdIonfwB+ElcqjgITTo/qcfMSJXyCewE/JDBwJQnsGX07bmjY
dh/NBAMYYjw5cHRNzGC3VngDGdwYv6Nc68LuyNZ6v7ZWTawL1K7bxLNjPUoEChY7
HHPXNGmF0dKgDiWWDWGOeAlR+geBqJ3YpIDnC4BuugGeItXHpneBko344ECin+KX
XoANa9L5r2ww+3cLR/T4sQYmxMf1OG3V0ZzYEGV8I/Zt36OcwEaFTQX+gekvtR5P
jtMlXXRQNhv1ZDuCqcyfJyPFVEwQLqEH76ieHbwk7u0jOmbVc8XooIEY9GnhXpoH
s4vt5JmpmIcbtuDxqwI7zLqYyoSprn6b/VdNg2GKrMi3CVpxpOQ1MeXSoAo55M7z
RQeo0A//rAiArArf6FzIa2rgmMO2Xd6kU8q9iKRUNgC+AhZBAV6/O2ZrrgQ6DQp3
8mI0PCUsBk8ILtD6XFMWRK25aKKJfsUY8uFImRCvzmNpY5nca3F4oYlHSLI4A4+j
FSZ4GwUt6uMgOMFarT0nPCse++tBTgSMRxVzgadlEk2oPFoIbvEjz/GFAqT0LGTK
7Z5shUWdNfPpnTvft62u6/Ny1wtwtCeNQUa3foyzwCNiCvlI4ZLKwi9+Dd8ZkAzA
w0i7uavV0JY5uS4C7QJ/DMKjIXlTQL+DXSiwZd5BANc/4+RzI2NTyy2rNeyrbgrf
Cg/2nyPdL4+nylAjyx/wLbby4ITEobuhMgzr3fEET5URf+geWSUdkSXnMm30dHZX
aJqY64kkpnzXAelnHIYUksrof48d5CBVqOue0M7j7mxKytOaWT5R78g9Fc+xs+fb
nTzvu5oaVtWT7QCMev8ePwbyYAy4mHdQUZGSK09zQGCXoNLs2MGIA91UTPmgtEKq
U5hcX9EnFHjB3/Q9m2vduL+7T6IVtUucXF+vDEiqrFiFgjBqkLRcsJjeLRlleUxO
LoZtM5aDTuSSCsb9ZEOqP5/mMRMwV09B4MKRyJeVYw1w6/33IKTVLcsd+CpLiskv
NlW+ffZjm35wQ/3QzcWrsbj+4jBLECLOvaj/z3KZ2sz3B13FPrY8LogIK8qY0lDr
2bULQQpJNqxqxd+KyLySUYKHLXoAd7udTwhFtqMzgi5EEdbGhWxWcOkkYaw0Nh0i
C9nQ9Dz4cFXkdA56pLlerX4kHAASZilEiiFkE6I6F1WH9xkvmY6L2nJmG3wmVcuH
0FkvXZz9ilEZLtXyfr3jXauCRGzJN+HSSVq6Wz9+jReWArJnLAaSiwhR+lW3d/gD
5Cr7LgaE7XRhJCNEzxaqTM/rxqKwyvk8j187hyFArdT9lQskh+U1C9yNmGHi8vAg
4za9UUmE1MHbOemLCBRVoMYz5oXV5OjcJwmOYBfMTLKfz9S74tb1129oI3T35hSh
tSvZ0k4ZsbxPFfU8yrVhXc3DKn8483XGq0tDdK1tWQmu6+fj8fnueyC8gPpZG/Fq
jkA2eiGDtMpSFrwPerdPuzvj9ASj1zZvVus2AxQl/wSXF7Gc7DEWRTGcItx2LolE
Khnrnee2t4wifinsaG+D7nzFv0XClmPqJ2KEQu9VD8grarnAXat+LKymja1gQWfI
sjeyMkj3OtHaXf06PZI3Nr9y61ccUvMqp1vlg/b4gpSEoravzM2ZcukUL0e3xT0A
eqDsi5qcrBg8BEqUEkud74EzbVypVHs4ODTS5ilb7Hxrqrw4CVq3NftegEIOFtjv
JXuuKG+3V3NkdXnZqkl9uO/q/FERWyoVGlyjO0ylkFhEHzMkhuthsaRsoAAW4xqv
l0SYb/pGtHKSgcFYqcosbov2cwbkyTNICfQ0AAZiLKOeDua6IQRGdI6YSHghbbMF
/o3hm4WfXjorZEqvBGPNNzQRUgB4w7lGn4W2jgwfBqzyedAOz02tJY9qQKJvaE9N
zPmlJlajrdf/3mFK48fXbMG++qg/59lMnhiFtZo20dx9sbp864icGPR1heYkQUxM
92YdZAuPQDRKE6NzEBxf97cuIrEU1o3vuEqAvcX0siW7nkFpXyvIVFo6hY7LmOx4
FBfCT3gBgYm4T2IEf07z7J7S5/RyuN1KnEUzcIGEmDCemPsKAOxP9S4M2/0eLYuj
9ld0W80wLG3gh5r+qBFQWEHbMNngMy+wAoOB8VXOHgT+Nb796OORWoaw54OnqB3s
T50UndBMRa8E2zv4HF29EW6fmZgdzY9iVVI38Nhjous2ugiBqwp4hWBd5Y20NgG6
d5e1LBpyxMylVIJWEWOq76cH0PjlbBHRQ12BzeNQaeJ8CkReQ3SdimMUBbLqIpbK
N6MpaBHiIN4NxF81nTQbAmDGg3QOAPgs1s4wu4zXTZo42P9SaF9NSheIH3Nfdn7x
zuEWTVsEp3IHWbgf1DwG+n65N3E3kDoT159Qsco2WAwEBWIFQOvrsp7AVyhja2V+
rx+KeLY0BaYCeDVjqOKO3ZWJw8uEYJQ1HipvrBxjBIa/67iIgUeaSl0rXJfCKGKX
3PDS7EJwFU09w0UD1X5yLLv1Pv5u51UAYgVcburC/5TAM2oWV9Ox5GVEm0JGP8Cu
M2IqsUqKHbFQrve7YHNtOt8EQAeCWAZebqNy+IqbmKbC/b1ro+oBJuKD29XVMDQw
lXF5gM9BZcRdd/g5KTIdLWxMM3+8GGEQdRHYovdanMxjFba1wOC2uFrfhcB4CdYU
cGZM+HmzoFHYRB+auXUG7uDLu4I945/2Ye4Y7B7aQ4KXnYcGtlI6x1wgxDnjenLL
Xt8qyAk/v+eakAd6qCYTfnWimXIgk9KoQAyzWWxsC9Ye9pgHb3ITfdFilBHDO/Q8
4z8j7qtTUECpHVTqjLZvvFwL6AmSg9xnUvcDE2V8+Ju+IzhsKSFioQXM06JL3oEb
o0VaAg7lnl8P4QRyaGus+Nn1fQPTkqBFCGnFm8FXbM0oc5bTmddre2I/J0twbQX1
izzeA8BjgmBTQc8FEQu5D0lMQgW1WKgUMNl14XbbuO524+DXEZ9pqdFSAEmoX9Hh
ipfGTJSu6OwCfmzd+L3/hM9qcQktBfnFXEkEOINFba7EGnuMcVR0rkq7Z1g96KD3
0dQDUbgVy/AY7JVT8H+WYA5lGcHX9zZGjp0ubU1jwOG6QOgf3LM7wIJxn6bF/mRj
dR+5km2N03jJvL+gEevPTCx9t2SUmzHK0zWH9XZUXI75wGo2RZDNpdh3Gel4FbFP
84ROgfvDSY1IhfY5XSba1HNNzy1l73dSnJoAXErComFZB0eZyHyCa10aV3/9do4S
ZHf1nGUM9Dz4GRms4/f1kFyPxMld2+wCwO/c75ZWXEAto3zzI0UAAUZqgAoRfx2Z
qBPETpa7/sK1s4il5v6Cy283oDGgFiTTPwQmb8ABR5vcuLCe2CDn06CWwAqkrerq
82J1GL3jJ+vi6i8Wy9eZ8y9qrqz1dBMHTUjETnjQFuEUZHu/NO0EW7kXnaxKY3cP
wK94xAAYRTOuAbx0HGTZoAb3evIEy4Zhlk91adkzvIvhuPPeE4nOhrFMNtrc+sd9
PtyfhP3EONMLY+6WVIEOLGpxsTsYeu456ULiRO3ajGsHV41ddU/iXRG1mMCie1gV
LHsoTyn7laX2BqgQB7EgEkxN7auKw1DGbq5/EndckkBfzQfcszxQsoic+lpkCsyG
BFIAGmox+xuDmVjyCOSoNg/hcFO9RwWfAwu0/cmBhuD9Z+tjYtcdVbX93TafxIaK
PhXguNKgzh4hahgsArycYJOHLTcwY4SNL9XnYnqmBJf2P9ZkFEoPrCzcboSJGxV9
Si3A6wct5m4PziFCKIlI0YUN+Jv+LacIVlB6BatJ9NvZyY9hAroMuTsXzKmsR97P
FCoJl+dIC0QgCNm6x4Ri8iPtwjRk1eD7SyZEQgqPcR8PLZlSEGGcUsEY4kaNJksy
PyszWc3jvsLx3RMFwX7oTJZwyRr8BnoGcEW6DavfTQLxU3GqapggpZ8UxVJBgCvP
4CLa126p7e9ZKDrqjKKI7CYyiUuzjNaNUB08kBHHyL/aUtOeI3LlnCvNH02ZpNlJ
SaydHMEbgKx5tlnvD3sW1bNus2KinnKyO0cDKhAaMgt8eSgJpNPG0308wesA4TIq
n8BZJoTsIP0pk8uiC31V5I1L3KeR0FxgxX6yEbQfhBgDP7dEe0+FsAJwBXomWt2H
Gbz/1nwXN43vOOa7yCb/meQYTBd32O/4olHCiLSggd27ixRgN1TaEHlx6qY0Phxf
z5AVK7R/34I1AImtqeBU8z+YRQLXVielM1RWV2sV9uB+CB02v9jCLZnXyOEA6mWQ
xk0disWLoro7V1hdA7nmFfaZOu8mwv8a9xngrPRTueoobGdtIAbLrR1LBi77gguu
wUYm3Me5kHPkFooQ7Z4Ww1mYBCp32ipkB1/gecntrhfEZ792T4Kcgwr+g767QXcC
7YfS4WqSLoQEpx+vMKXM9AaQNhmyiSi54nRvYOvGqyWWTqUsh/bjzCGLAfJGWTe8
/X0PU77+PSjyOKdySkmoLs/qDJSr3ANiDcGrUI42qg0ZoczkHX3Pa/1Vdfb/WO6v
qF07Z+e3YjKJGBKtQrjCvn4lJxQMn4tCX9XueN+Nk8ELgya0oe13QTfsd58wETyL
8wFv3m4Pra+uDhCKeNft+Yiljv6FKtLKmV4C1wTufB11VNhTg+VBWC2O6c9v2jmS
CX/3mU4CcXRbVS35o9GRGC0yH4lJbZ5XEoqHoSpTvrREDhIHsm51ZPVIi20yFAK8
YSwTqWICCEbP5Q8z+1NQUl4vJlsej7TyjQgEadMdcLjxYXE3s5LGCq5f66kp/AuX
UtkvREsaHCuBd+xJFLhccuGaKwbQ3guWiAD3edb0FmQPeGHMD2gOTCjBI6vYYYzU
NCi9oba573jLb3u33BDrqooidpwFLDqXI6jtgwIrVj1N0LDLgpq4l2aHwNbcUI0p
UDhNwA+PiuKPtXMd7QbzhmN2FUvi+cwtxodoexehfkI6STtdOBh8owkSLD3I/oke
03MDY+uUxvWTwH3TOtnmRG7bm4SPzct6LUd+qf28Tv08VZwzRI+tAmos4cj4UKto
f6v/QrVYxzZEGu6njO6hjiFsKtAnfh/LrhsajLsV0dimvvmM8LVMxZgeRV28Zif1
JrGvJRDM25rUNt7JBqvRDJhVuI/S0oVjSXjFbqwSzzjMenajdQMVahgJ7EGXWBUP
uFH15ZhDndf/YNTMi5fzwMrnpJMzBLDoIlU4R7YNxtAYxJ4qPLUkNbZ9TWfwQwSe
Xns5EvZV8bcpVrvbNopISVxQz/fvZ9cjhVJqlmxOoDcyd0eAlRShDix/uPMMIlIQ
I0J/VRUKTero/TDeWfMiDV/RbkwG4F/sz5t67mRJhcpCgVKnwxrTbjKOvOfeAa1V
G3AoKcmgE7HfHwSnSDVVaEP90//A/tW6rz7PS9FYqOvc4kGniYNOqnKHE9N6llZJ
/AVmSJ7RqzNxxkzC+SpLE8MrJTSJvNGatBmqECznaGr38cdoyRa6IhX6wa5DxxJL
xv6ZiQ9HO6zcli002n8LpGJyt83yYz4CLK2GPeOydXKyzBl9xa1SQSMs8FFxeHQ3
fB+AZytAfmqBMauEmYW+Kz8TUqls0y1GYMU5mmaRQYPZ0eOR+vbPz+Pia6OT+W/E
PXnvWUt1AeIe7tdIzf2We80GIE1oyxoteOkMl+c8sBqFHB+Xt41CARqtYkP/Y/cu
KyQVaVFDGRXB7dXO9nAdpK0PjqYWdnBiLYS1zDuWaOId1BEU8Piq1PZ7Toe2sWjA
pWtGnPYEptXlZCAHIzCLzrRATDBvWRmRJd+umCdH056iiXh3FjEQoOFxWAwZIIMa
PPpwqIZdiGrCGDH+ZPRXPgohgnEUd6tWgZzPN87YcsaBoGEhkaQcjet/Z8/TyMXe
MCZKrs8b5ndhry921c2sS7l4dJzAC7qYPEHC9SZhqpAwHPXY/5AFVgUB3ADYvOqD
06w2SXf2xy2swobPz/Pbor7hz+LH/tQgqE42MLtuz8hH+niJIPkQ5TrKon9MMld0
55Q9Ftx+OYZw1+gu77WhosEOYK8doxA5yaDN/ZdZLd3/D64W5/rjZ7COmiYBBr1Q
FdWfY0kHUIED9Sf91PB4vdzEqIqwYyrIQyS6sK18W+NJoZNBX2FbPgGGZ25in9nj
FMCS4WtCwvop7fUHKwJd2QbNFegkFOq5FxqZUPnt/KTe4Li3hiHZZ7/MGjyxdx1C
DCyxIQ/3Pc7dJRoLgCmm6dKQUZBLReLn8YGTpStsVy7hAX5FBkyZkFXQPHC2GTvL
uj05P2Xmlp/Z5iXjoSbSYB4YwJI9+/CRgMFEz9TxN2I6advdzZccwn0WM2qFeyq4
/56o6ApYrH+NBZgYrMShFbiHRGWxZXuiWWXUKdw1RjIGkh8+jOq6DIalruTRTceT
rVpWd38DfCq1iS3YckS88WioOahykmMd/TWzysQdE2pGx7P4tGRQ6FOZ4uE8RUg3
bFWRHiAKcLoYfIbLWPqIFZIQ0HwKx0SNgrK41SBsuwz2OfGHFhqAdslzeNwVu2Cz
Nw1DYdMfbLi7tYNq9OKhVCOZs793Olh9n6lsRWPwLTJqnp7hB2eKYLr3xxGE8sgJ
LnYbL53rxO9RhvIL1mcLWb4GsbEP92Y0UBXOr6uOc0DkyBkBHdbwq7Swy1h6LMed
WPy++Rr4FMxxvZPTCpwZfAZQCaxDapqBjj8qh/MQRlVN5Q3+VIuxqXbxkInqnj5o
RNVs4O/BbPuqbmb/MKH6LBhU5WHBf60ER1wPIBepPNLo4PxpY43DL6qq5a1bJTk9
4cGRq5IAza77XmzUTRFP1mhSv0OITsBu7c76jdavONZWKkIPV3WtUI7OsPc5tOkm
KmIf/bIacrw3EEh+ai7txsEYbCmYWDhU+au45KyV5Y9JCnagDM33GTzGmffWdjwo
3r/BO4DuGZyz+C82vS0T7dPmNX9q5v5N33SHiiexTPOMVLii0SlI5rfiKZLGEb9Q
ZRQM1UlTF9yjbSsGlwaFkRE13oXJ150viu/K0KXwjWLUMfbjHN0ghG7i8kzAXNPX
UoeH3fPjPyuk+MyqE8lsZUyem+/8chOF1StmMRucSKjAgz0Ndma/y7ks12Lv8pAS
f2RGPoNLWkOvxN0uC10wAzYImogOfhGoTRyQKjYY0TCZTnVCq0Y2Rx9AbqbF5NFC
VWGUcYilpI2igBrezDMs5iD7qbkUBYr1w/jyUmb/Mc+JxFNYD9Au3fsUH61vNzNO
L8lWSRmJkD0j9k9/Af8SQ/pdVTLnSICoAlIuf1oDUIije9eky4R1LR3Pab2OJO/P
joFOoB7TOWvk2LT7TGXiXVOZhMCW5o6xTPzw2YsqDPLWib9asIdqgy9Tj+H4Qmj6
DCA4l0f4HcxWS7fdVWe14VWD1RIPeBX8mf8ujK7+JCIu84lGe2InLl148rMH37GD
BHJ+P9akSsrtsO45Rdp5khUuMuJIGLy6pYVSNvCdFFhF+TgzI6TbBcg5WFR0Zhjx
COquBEedM1F1VXNqcShk8xfdWZ6+xVEx3hAP1igbRz0BrYvQendduXV4GACSt4Hi
7WyU0fmcTcpLR+vB3+jUGXY1269z/bvsNAq90zH417XC6J0MfpAc2wOzyc1hE+iv
gh6ATAXONFy9v9oy6Lzi/8B2SRs4d6XjSD6jfRVqlJGpdEBvKt79ChAJAqt0ytv4
I+tBPC7ts2RskJ/C6+bt+N96eF7WRGoqD9duWCYtdeOF853GFZcWpQTTYpowWhhD
jY1JkECiHOnyHGUxMlVFgZewIZui3mG9IQeMt4dHlVSHcc9c8f6cOGOtZ2BaqhLF
ezc7GCSxrR3uivn4ILeyZhbrp6Gy/MVPgmzNccNJFeJLWJJfiWyZJs2eXGjT6tLt
qXeFNX72DyNQS9obVBWg77vPCEYIss6mMP6vtqbiZyQQw9Xk8Z01rgpku6qDEgxe
vZN9EDlDvV3EZxCnl1xN4PbFlEeA0DxykMIJ76+av8b3MlqoPTSNhIJwigKJFEl4
0TFiOBn7xUMv9TLUYXA8rAd2AETi4Tj5HYF5JEIyfVeKY1OdXIol8KZoBxCmju2j
7uL/Z37QkbWxqdqCkGflSM0yGdB72IcAXb0djMTnzjuh1UZVdJiTZaQpTovKoKtd
KZSFbBwZDRGyX2+tcwp9lUmBEiXckJEKaRjvMzYmgu02UJF1NLcwYsRUI9S4cwKa
WG+HfYKSqa9g+QzW/GSLiNH//xJJsmgIqYbLfV7Xs4ljUug0hswumJ7yExgLk82P
zHAHY4Tjoi8dmAQwYonufCos7EGn0811oEHdd042bvvGfGmZuHHYouIFesUeX/Gl
scoMIyhlbXve3nxBG/8pcKVKTt8INnu9bCy1e76cyNKcxz6yTl9iV/t4BobXWSom
f3iRNSVn/6KGIJlQzPYyIHvO0/8YLGE6stilLl7zbLVOIWx0TMm8KtcwXigh7nqh
f9WbCE+urVtySw7g7GUDOtg94+ZVYemaFBkds6xp+3VDhF4gyQu2OdMqbMutDXoF
ijYJ9W0W23wi/ehESHYjHSNWZ34Tygdk3V4DZZHmzd2FTVXh0MOLfFhQykKkYGW+
JaWbEYdDa8ezPWMeib44W0yCXoWlr+2YlgFQ+NaIsuJofzndPwyP/q1HxrP620v6
QkoAgJvAlu5HvZhkP143OgH4Ua2WTWCWJLTXxV+EWYQAtbq91b/py9In84UCP7Yj
J/xgnMXuZPTyMb0WxgIun/5xN493PhbheaYGzDTZuZ4wPd24GiynrtaVBlhm47oh
WFoFycoSwRe0ED7JPJGgOKcUCZaiu1f0WByGUVxaN5h5fQSCvrI1HdC+/QveBYQp
FUxRnxqYL1TIvXEs1S6zo+36GXUH96c36IBdCC6iYQ5cfca62wWL8ElhAwP1JlTi
ygIbMvk8Hz3z5RIbO7D3M093GAkRPi9nmNiwQFOqmOcW38wiHtOHBu7LYkDn19Ta
Gg4CZisOOudX/L4ruthiEdpVgEt5M85SeoXKwwLdzT+/ns5vQGRbVm2Aw4g3ezIc
FNx7JQ7WafJaxYLtR/DpqmoZYH0RwyfBZsMupkvI4bqSUsD4biov+3cU/d/VFUyQ
7frQR0WprudMgSLlg45fqFgxWBQMII4+ML26VTGjKXQr3fbv3/jAvOjTiiC7ZWCK
OjigfvNFugni9VZkUSyaONCSBuVJqvP0fR9RQQmqRiRm0jOjEQ7oRw3XLUbPJKZp
zZ074p6SppgCt8q3WMOEX6WcOQFjUrPVy5Z0Sjq3ZdZvHiU6H4Zl1RR3J4/OLY/H
QxXyhEKU0VSDVP/99Jg0nsT++5hMTbmbzG4zFW8nNv6TApavs9Qhb7fF/Z9bJusf
Mjgoej71MslZqAVRU1I4pz1dBLF9xf0vJBg7FbPih0Kuvw4RfiqJgjL22blEObZB
dVxnZ2VtJhS1FD7SLvyYgekUj3hUTJL/6YFxBxwMs9fwBM8fnjcPzF/iOcw9Omt7
5PiU/xtZYPO0kGxHttWJGMYPWgj8Izpv8+i+SHWt5YDzA6pGoXQdKQXkEGnOV89e
JgiMxi0yZtkm+Z7jpieE+nhG/wyxTT6T7Kh64Q+KsjHWytCMk40JjDiVUkabmXRD
zV8/ZVdAHzcEPRtzSveQ9u1ubjx5C+bFJg5aLmOTBjSdMZoaV0aJZMLAdd5W9VeA
qaXwcmFk61E46VwgYWKTyFpIuAl7D1l3ZFtYvQinTpoYyIx2SbQN/HQClXAE5nQI
+n8h+BGb9xfOXi1q4eJj3APUUQM8jdbIl5XHlWoJzyG7JN2CDkHZUtuc2PKlEkVp
qC7Qlhb+ZsOKp53tREAJSzjzzjb9aFJJanO7MwIAOhB39MoiEVcaej/QqOfKhbXu
7naxauZJbW6z5Hn2ntDh1VqhGNNU599WD3t31bejkNUU+cmKezrYATck3iqBSZqy
sIQBW94BnWxyqJo+DtUPCGob+RC9PDeLHvmyVAqN+YEgbbL+QzGiH4Q7bZLyCUhf
YOqnCiopECACGodUUgAyk4QG7xRIbhwnnc+tcsbupAMTmJ/7m6l6hWDGITEGnmwN
pkLQieIUUlbkdt6BdX0uAsKtKa/slPHtRwqEBgJF+atNWd0pnhgCgw8AS9Dsp0uN
62XUOgAQAWhE49ylvj3gYbYuXK5lQIQEMv6XefYcWpAGBxfntmuVfzQ5OTL+HWBs
rDvYX31Y8DzdTW4PbJjSspWtxxpoyjUoMf42sXwuYG/nbQoAi62GJa9YvORyFVV+
Vkj36GMjcY7RJ6B4R0cQUwnlR4lVr0MUpftB+5tw2rCEa6q7cy1ywbf24BVLnUB3
mBZ5+AnvdtOU9SPwDBl27vvGZV4hp6Nzu8fONAywikOO30EI75+Qig/OHup/oV9d
UPtuY7hRDsArkzYyKH9ERw47EtpWUqlrz+qV0QthU2tYzf5vPY92lkALvG07TOYH
Lav88rgqwdLs+5iJ5uhFhbU5eg2i4vZd6OdFUbKX87zYpFSH+qcBBfzsZbU1E2tr
HAoLd0/9hx8asvEYc0l7oed1z6P6oUSnHcPwdui42SdhEvNm1zRi/357bfHrXTm9
wvDYbyI+9/Uo2nhkp7DmzIIy9v1KXQiON+j/VG4Rug8gyvvs20Ial2PIYngqDqft
KwyLXddsbLxh1wzo37Fd1XOUgwJDa1QMncNGY4Rsi0OeqjB4CZxsO8LgLv055kSV
/Wg2nq1+cYoXgT+gzGW06NT7Erkya0/5Ap3XkRnuaWHM5neTvYEd8DJVFawsPzBh
onGyR5Ngsb6oNqTkJTAEc9MCc66I6b5PfNlDeMj+NZyIl0EmvCAvTDWn3K3pjo6V
awSoIE25TrwoGJ3oNOEKyOJSVp7y+eWP+DHfvandlbs1TFx6XCmEf0cKRNxuRFvS
XiT0g7gbvG61f8aBuKaAZPmGrrjIKL0PFDIvTXOIMhRZCz5himxTjbGvG0yZNbm+
YAO3z3zpmSpwVrBvaR+Fxd5CqImAn7ezS8p6Z4VCIhIA2zAWmU9sdLtR96Gsk24z
0oDZ6qQ3ugdkxPmIEdawzK5zCFcPJCKugXcTr9Cs4o+NyZHSOQg6FNEeUl311niY
IBVbDEBoJ5Eg0bfeRyF2YiyGUQWJUCRCEsrrKKUMX+ueshNnQ3wTgc9leeoTTcWD
MfVKlx4E6U0i7r0kBFdD8rrPFu37o9x9HDrLjN5WYXw4biBtzPm6pxIWutaq4hPk
iIis83/hN3ntAo6VSBn3lHcPhcF0Ly9kgMzgMRlxKTMof+cvtTgjNJlH0cVTQScE
Om1zbTNSIVr2SziIUf6V6pGBgJfdD50rH92DraUMk99cS7J/E+IEplko+8MJ13Pc
WU2D0fgnsqq3m9OpxUgw8NKjc7ZEWnYEt7KZGK9FRbOBjRrFV2dOzcxgDDdnyLi2
9NvuzMGEMJYhMwjmq0HWmjIVtIifOfLpJWbTApdeVHKHN/0N1x4OeA1RFwoRcnAS
jW6VgDJZ6FRsuEyMFRBFxLpDsvFMQlShMQ5oPInlSXKwgJJycLDR+qE/mTnnIjnW
6QZzTiP22jKiGmR4q2NuuC7gkGFvlD0GoyAx1Lqy/VwjjOuFmhf6gNbDjuI+Mxeq
0WdM6d47qQcMAQmEeWMzYCQNLLcPtbY/XExn0ot8+jEscVTcN9YTa5tOAZHBZ00L
W53XS5SxPu8SyDO+IAwUHn/H6RmCXP8W328bskPRbj3nRMmBHskYMpV+XlCvA9Od
x1SjpVMdMIjNf1ziaubldAWo6HWjxlVvvCnyjbUKmeSXlAujqsv2se5ZJL+c7TRI
86enTUMb+WGojYVgv9XjktnvyeZhbIWXPx7VGporiZGgDhHyRAERrS84cXpFbyip
EOV9l6o/JuPgva9brYvWznz5eqPyWbk9+XM81CA+Itmz9sJW0zKYBic0ueF85qgX
21QJfxoVV6Nfm8EvDg/1TmU6S5+N9XRqf/nnsvMRrl7F3jqPaDZrYYelehg9/tyO
GzrR49Wsz+2lFebrEUmLhsog6czPd5dgFMkjCVV2AWdlj+QiLVPlbaH1QTvcofrU
XlBqqrVTx3mxBPmrQ23oeFJYDIArNdnPNndzekeyItiAWxCSyoNFqw5/vLcwNT6T
tfR6t94C5GHhE0bWJ1IeyPKZBIuCTm2Rlsnd8ZMbbJfjW7vIvHOkT5hc8iDgtaGU
qkgGehsyKpMFeyKrUVTgDrU3eWajg7QNDCIGkNceXqYYDWzMQ0uCKyk/m/oGR3Xy
Lgw7t2ZYSyoJFfccGRr6eyB6GBIBbDteYfk3uJxw8MbGkbt2OfsDicGV9/GRt1Wo
78WxrwHH7DZiv2bqerkQUxfPZUnNYnvzqTdfxOhc1Q5OR7Err3EJ4ddfFZ1HGmbY
YMkmMTlBtcyFQobvWoWCPpZ3V9AcZNy0QBBp9DvB1nQygM4WWC4028WV/cLz7C2J
tDHsaEP5WVLNWRzJ6u6hFhQroW6C29FNo6IDuQ37wDBIvGaa4VX3e0WC64QF+35C
PX3dmoXpx+B/4CspEro/0P4B0nWaz6n7WUGhryF9Le+NQSnZvIWdFJF/q4GlPvMi
bWY9myNkhqfS9wpKkLBXRfRDYBPsskld7MFVC7XyYpU6/Cn5Os+y9Y7mXZSu4/aK
G9mH8saHk/iiA7dZZap74CgL9Y2KHvWvRV4pXhA1B6aamvtJt8vOySaNPhde06tA
mbEabdop6Jah0yDNk0vx7OSj5T/WrM+Zj5Ft2Ds0BS1M8hveY1EctfYzxy8xL6Op
2rVOAryxVvU4TSRlSKAwedSRypLDURWs87iuy2bQZXsCTUZ8iqrHUs3SLUawdc1f
8utUHdpzF0KR1AdEA/jllDafWn0pNlDCJoTrU1YZbKtDAPJm2fsy7/gZJ3Z2OahS
32q4g9Efnp5o9mHzjiZfbbujWtMdxVlKt9JgP9G8fVXzxTNS+cIIzA5hHtfg8Qyw
J+Sni5pbc/ecdnPw0z0x7JgNshenz0zLfFCIQ2ELF7PGnU/3Gk80iRgKjB/xkiux
35pwNjUoboEw0FW8PyRjTSFd8VHmfPkm7nhPRaW/LvyKFCWvkObX6LvjrkkBFgRj
OeIob4umn5COCtpeikoJeBD+kvaoStfZqa0rMiNSk5eAHsRGijZz46H6QqHCyPuA
MM3SMoQawVaee0IsDhztS7EXM33tQh1YEx2fAlan1M2OU1Ax5JbSF8bc68HqSzwE
+wOitqHY5WppIzVubxHipw804ziwJacJnGAGoovdezsu1KKaZONCShK2rRnhjRBg
9CZewlF2czZkazInJaH6PFFB97sfuvdR4woZYotgZdzRvUEQw+oSWlR5nZVtL+gM
KongSa4g/OrqgUQuAdnU/zTlEmR2m119/69DJ2L+1eCF0jv9WQY0/e4r31hlfbFj
qMojQ2+r7PGhap68x/mYQV0o5KvzFSxtuJg8QnOT954ycmDV1e8RjOliPuhgZucY
0nkHoL103u++yHOnpV4NISjO82JAOuJ3KJydOWTkoSwz52lcg7OIRHApFrQtF3rV
OuV+7NRrbpXUGdlwyCL7rMmB1w7hOg7wkOe5Qr1YMc205sofKTQYfpVheXTFYPUy
RbmOpvix/nrR7jytYtzqDSD2QI/acCHOAfuF/7+VBhcKoKVEGpmw7wijyKWz7jGg
HHpcDFnoUuTi/Epb1+xaIhyIwKqqqppNbjoHGTEDUeWVapaQsr4vtnBGXOdpDE6W
XRFFrT+Nldw1nGE1Q2ESca94JqrKCOW3W+OAc5Md/g6oxNS6pRFAs3oXo2POhMrF
jnwFvoe2SPLAk7CHsI5OqK9d63ES8lRZY1wDa8YcJ5UHhBZU4fgw1mjoQm00jj7u
1T35BPeWpOQlIhIwKk9ke6t/13baqHzHKnJ0QXqH7L8rfSYR+CYQFRTDUJpWldYy
WCz6o1u7HiV8F34JfZAuaQCskluehAOGX0sWjR+GqFwakD61gFn5UTO9xmCyD7Rc
klZ54LVZmBGn3aFU20lc51eRcIKaeXwZjZpYkqp9MjUZ4BG+FMJm403lz8BZ/ejv
nO13Izct/kFXTYesvrMklWVavP/np8pO2iHH1RYNAEjwxZl315HBZsT0KhF+YYj6
bx/JdyasG5uGTTABSHFJEj4SnDH3K0Dqo1mtuGQj5JwQOYjFZyRq8KBokmSy6kmU
/Zqx8BnNEwPa3gJmz1jxs6RrXlGJsrNs7PEF4E3juMEa3sc9YEhY+CxERNrzRxYV
v6uQ5S5yhBEMBRqcXeR/DETsfqN7WM7/8fOUhGEXgjfFDDI227WXHJMBi3AH+cnD
ZExMEO0G7HsM05Q66FshZdJQ4N1qRG2tXEcQAe5fmHKKEKEPYgaDLztmzU5FzfOE
cZXLD6TJaiunYRk5R/ZWzYKUf9ulQMK+6P+5eMYaMLt00vKEshzkp0O7U/Mv8Ygz
QpLArUf4RKtdp9ObwK4KfVISlUbipexT8NS2hTEF/N4TYm+nSCst8DX4Ysda0EcA
4AlFb4sIsEH5ET0G/URBnoboUvlO08+XbOWGlkmPJZCn491Yiw7YrBA1/iOcpbC5
VKw3I8pIQCVTiijEFJ9WiiMc8XleyH1FR8J/+9St2MhwH2KagqRzykBStYdayTJ6
QCXcU8BpEbXrBdhSeTTeeUyZGt5LGGtrCQ8J7E8vVZkoWfsWLqOQYx1bmj0ZMolR
+MzYegFb2FmAvblUuLp10kJAfEAXmsVJmB9YBxdeskU6qN2W6ufr2dovJaRXwka9
R108PsiPebNEaG37sAZKdpOLRhjb1HtLbnAorlRCwRv9F9sxFvuH/9vPtyz/H/4c
jUYVbC6rpVwtOQinvck8TPRy/He1S7RnUTdANB9stLnizzsqVCbDi5AYlGKbdzqE
N3enVK6IKN5TJSaDc2dlG+EG4VI7H9Zlsw2RBXVDiF99uQBypRx2ryWXPZX8buFW
/yxEyYaAgcJ9Ma1mypdRzQKiUbLnTgegmCJV+nvYCOTrZP9oBvVgJY3FuaegZPY+
85cuKO8iAVlYaK1xrj1732hZ/UEEd1Cx9zKywvmCn064ejiA9QIuA20v4ZjfKHeg
Mcp70LQpq4HkO+4H69xY4UH310nmEc6Gkta1t0dqAaiRTEiWzkc2Kr+rzmvgjFDM
kAnfwEBQ9hXrvBH/4cuCEtwejhR/qXyEdZM/vWyhbe8f8R+fb6tL0kQCJGqkQEZ/
jce4wTytUMpvXc0ItzbyIswlxrPPH4Rk5d5l1wc8f2f6Hz4S2LtspZIFa+eJV2Wv
dDmbS5cdmUMb3XydAg+/y6G/OXgUKs5+b54XzslgpU0treBLhs1muqDTmOV8XjQ9
UvEKLFGYy8C01r9+gOJgMN6Y4bXN20fXACbdUaCMVH4mXneICMBhe6gU71ja5thn
A3CGDxDcoLdcfNVEVKbI1ecSdC7j+tdnill7DO6uAT3oLCUGqulk33tIDtP5cCS7
jMy+bsA/owgcc0/igdE9m192pT1e2p098U9v67KLzc0SkS65C246FBk0VALqtxY4
wpeGwABkSIg6fieCZ8MmbGw0pziyQ9waIz9P3lSYz0ofo1r+dORhDx0yyarfjDhr
5OU/KsReyFiQ2uooTnjjrY6BfcILnqAk4JkE6Nkj3ksmkh3qSbEa5JKAtsMdP/3z
YNN6GqPfM//FDEcs255WwUDYWdrfjUSglycDdV6WoZK9Wv1c89EnRkfdjM9jlP6d
kzOXDnVr2W7v8kiQB0AFY73NxXChu7RAiETH2uMBhj8kVEreabCtv7gBS5kVXywh
s0oMU62rk9VZI8/uVSylz+Nkh04OksPM/W1pK7X7CzTaqE6N5k8X3p1N96f/muN9
ZL1f64ZOpy3J9tadHDzLDcr2KLJkyNChlHAcSPVCp+u0nA67mpZGeq2K8NQUmaRL
gd1bznCWzWV26btaqnI1ssE+KER3xoSKoikPfJrz1qUnMsPvqvkF56dKevll8zFQ
G1NGE7moYb5bvh1/FFkyZo/oPVU8T0Ks6iSyUkD2g947R/AevpxZk2u+9tk11Y1G
Qxu0lEzxKFobmfhWv4qpomd+fdzl5cPwpWqgkX0TEp3t4xcAIU5FJ6eM3ulTqOYf
nFqDc+5Vt4gzfFy2HtSnVc9kYpG9MBNlCWqY/MFnU1G8Dg1Rbm0u0xQ/BzquD8rc
mueWn+Ka4OiKFPr5yajBg5yUZoIbwvkZkXoADfpafBuO/lsPMe1Fi3aXg8iN6iUD
FY//VrbWGN2zSkM00u5oB6vMMb0WX766eR3WI4bA/NizJJKT4Dv7ZZjV80U+JG3V
qknsErd2myZ2pBl8RariFzO76q6d8CUd5WYgr6rl8utts7QMARNGazXpLDSXmpgU
UbcEiaApTXB/ykerW4DhbSgyoKVUoGFeua8NM4clZKSWe9aFMEoj2uhQnwCcOQaC
lmjIybxZHhfu4IMdkyllq08UQqYVtdJDdCiDp5woVZhsuOnxrR/bQXyUZfxpGTvU
tI6voMg9QlNonJJW6ux2ObmOTwFZJYENPxABm+5ncBzPDyLMvzWZyu//pUl5QA6r
9vYfO94V2qXRkRMvdX0qrbS//hB5gdO0NTjV64tYY6CnIguz9CSYlGyyCHaXcNZz
pRij5sJZ8OabNoqED2e8XNbRGb6tSyW3azFCK0aXg5koXvW7tinDRipP3nBrIfcL
Ex6FeWgxfGD+ANQaM7UV33QcTivltVMoBlcC3g3EmSTaHYsU/OPIR0gOlr5r1ueF
nrfF2pjtTlpoGbT7zC9CO3ACsPgDvNO+Hnysl9mP60xozQPc3EU4T7REvFl7WqrT
KrDeaboo47hmSrrBohgloTKn60n52lOVpZQOtTjE8mIiCvcICeFzTZDN8TEF6DPT
DNZ+AYanH7vHcYTIJHRRugLkt/2JNbig49lOkxiVvzVSA2oLPe1eLIWXLAA1ZXbV
S0/Z8sGSCy7Qr0v+oAPZ4S6ygMY5nfSdEGamsfLRpOKP03H1c/VbeSpPlztz9C1W
rocFI+wML1Iw6sQasg9eMliJE4R+RO4/1UegoLjv6hBqds0V3QGEMLFgGj2bamxj
bas6FaDXm6pysCKGiQb+qeF8BWSKIwg7RG40YOJ98SCqNnv8USFFdnCqeFL2Qd+6
a6bv9FusdX5XodSeTvrVpwekAAGb+1UjxMDTSgHehNFwCkSWGFQytrdBV8sDCJ5l
bc8zopkvHJU6C7TQ/s+T9r+YIRw8YZafNAcOCxA4+8PZ3sWqBYXx2wKx5jBmKlVK
/bCa8bNGNZ5CvZ9DnOj4kufXS+IotfuZA0jv5yUbZYqLP5Y2/3jKRcLgV43mu4x1
xhXhylA/KJcGuHrmBsuqHGXYkn8pT/7PlC6QXmZZXaDSAyGHjCZe7YvV4UAZdX0U
NlGSj5uLuR+v0C8j7DPccQPA3x+B1GsBsh2ZGBOIfOUg0xTR3dPt7WRCbGqfY9y2
3W92lZs6Cc0Kf1aVpF07xYzvmnO3TqIrxVi3sh9qkMu4MxU34eZEfKwzsSd9ndm6
rD/mx+aZSytf1S68I1UU6/e6mYGt1mzjmTag4Ht6yqRw1uVXHucfOe+myp5kTNtz
oykPngLYh4Jl+hmxtF9YpT5Q27obEWp5dmaZceT7ZH3IWhh0h5hKo6PGOeUnh+gH
LvQmT0LvwZHAyCEvgGAMxNUwCzWjdqFslc5YvOXJC8efjpfDWkVHdKDmNC8qg8he
wM0mJ/Q+tHg9jh3y+rlw9lh+deqCbgec3+LCdpAbSS4u8aIWjtS7VwUjIB8EMObf
a6cKFpI/TLekBhkrmPZYAqB1ZM6p12XUL/XsuSEEUXPCyrWf/hnqfneq5R4OyIyu
cDnP95/DGi3ZPz/TtQPQV844dA63f0vE78YbBxg4hEm7AtqxOHO0FsdZIABJ9nFP
woto3edMZmQUse4LW80Rf1lBxmEA3kfvbqA3t+zqczERUjkoq5orSdGW2V4z4vb2
w0zCmyGL93Dji9zItZbrSvwiqDJl0kkgXDPF+WHkNjOkHPUTpamSibBidWtZDXM1
di/dqkljYgxTnp3tjrUM5zZPkSkhNtFesg8ltwKWcRFIv3iv0onFdSEtPdjJc21u
Rl2N4XbTqkLMD5XjLn4OBmozo6hdpnCxzeuRfp1GsiEQLftri03dMmaCXqMDjyYL
hp0M26DeruyQRHN6xNtu0pZy3Z/kYxerxm0llEsXxB1Saay+zJ2w1y20MgCm6TWO
StHDE2IlnqkKC4TRrU1tfNd1ghTyMdrzZXGWO99zfnl4XFFArTexR8bwcMDfr8d2
nqKnu3SzUFduCFtfGUPyD3K0uTpdi5nlWwgXVvZi2X8dalt6crPiouT4CAGdOtWB
4qrXnT9xKvqMLuJ4R3d7+dIIepF0hdjDzubeOPU5sL5C6nrOKD+5VqDvbcBTNajB
FpjevjXlOLD+1W14pGKUJFYNyHc3ooqd1ef7bitNOUT3QYpUGX76Xw+jr59apgfj
YaA2oW5RjKPl9gq1wwpezBg7CIfmOjhggs2jGnNOD3pr+/sGjddJdo6RSysfxCu0
wAtLbix5bmdJ7Ve26bl6k1oLlb2zErIVTPBuEmSzoxdozY49r+wygDENMp5ycgAe
gAI+fmooXGU72J8YO3KkRZiBHOmjRp0luDdzLlxbvOYrCbjF1in0EyxE1+L2DU17
BUhqKwIp6YpFzVYEMVeLIGhe8r6td6jQVufX9CPI0enemJs0OED2Nu0zStP3O57f
VYxuJVkEmoUQ7CxTrj8dHATuzD4DemVkndzlf409bACPaym7GBLAbK4TYDDSgDvT
YQ7YjehMPzc8wbI968pMha16Jk75SN02ICjn4bwYQiMrryopJRsqtXU/p7Ck7w55
WPWpetKIBev7gH+FQDAyKVyhx5MF842oylemfTZu2Q4LN0P9PZP0w43ZG16sYd8d
3ROTYyFwTrjxFV7OiyGScmI4m+KXUhZPtap1Ky2z7GWXDuCdYy9Gtse7t/eUKW1u
5tvMjCaXiK390rGjjd+orcV6ZvclGaoPBc9S/9o/5ypfq5HFCQxBM54uUxnvLUHW
WFJ4Ah9PwVVi7fZ3Lhgi75Z8VvvpSNtkWRL0hJ/WOsGXLCYQu4dqpDxsmSKdO118
e079jq1fbVKiHvUu9exppmHK1Lwme7MZbeStumOhJ/azQW9GZPVXHE7D0RnjLXfa
mL5KC4j7t7cKg9lJq2YQC5FxfHZ+lxSI6VEwfJexVBeaIHVEZb3B2uH3S8ErBx+F
wIyd5ukET6czSJIjHPnuWNcMPtWrUqtLcVkW5MqcnmEjbctPQS0HKsJ88wA+nFaY
2NZTE1ruE09PGBF+eSG0rHszfMllyoFm8+kN4rQMG86daFddO66nRDX7rSnU05LL
tsJpFAtAecw+YP9x2U2AlOZ2wj7MjDOf3rar71z7l7rwPNR/TS+BCKhZes0YjXMB
PnjW8obvBY2OMWgRAm8tzHms4x6ORMfoFSGMAQaRqMUjCj1WQmWDR8yf6ToeBlWl
dGfl42p2bJsdvsOSEqujMt2TY8m560KgPDijyBumUxUTOATv/+rb4hYuuG1lXHBY
UpZrGhP+2Oi2DASggbNclpY4yTtlwi8du36okCCgEkopgjTKHfFCos0P6t08OMrK
qpLSda0Psa87r4GK1vzvL7Zmh8tNhBiYVSGFn0Y24qXsMD7qzEe0xfd7xrTjOvpS
6uDl3S3uCFVJFsKAL5XMLeXPBRh896NSf57yyHrYqwNraqtpy1+IXPhnuqALia0h
VKy8xeSwX2juk1UCKCdaWWsKHaCJ9wSFs/YbJD//yYyr41uUSIO3t/UogA4y2uW2
KDbQAnWkHBiRvO9anHa9SzeciuGw5aTbY4wpXT2+DdWqw5ZcXV3V8ooZELtIIz0r
ixqaRfs6xaORVCnF+HgBXQZ2kiK3nEYFcNv3s0K1zc9bw/n6dtP0KkeZRtw3ign6
liGP9SLopE3WYTAIo7P3Slm5a+VXPKtwSpUrjPG6wh1KsiPbIZYVxYCJ432Gxmxt
oqmQoFWX4EtguxjSbHyI+pd0KiWYwa665KkBWRh0JavG1OH02zMV26sbAszkQghx
odeAIZ0kEOZxD34K2538/USY/VUvR+FVcfO1of7ImeOvRZpqwQJRb6wN8w7q7+g9
hg3srERL+0DXLhyMPO3AZnVHjPUYF398i5bIVjtyvqgDHfb4bBFEnIvI2cYPVk15
hYTesxcjEC/Xb6tl8Z/y64hyhnmVkToDldVoD2SRNlQKsaRF/Vzq9muFw1E+meXa
ttvXoLZq02Hf9FRaivy3ile1dSo2BNUKGkLeoICSHDuTaLmLFxC+PEtN350p9wYh
pRqNNVSkm4+vTpFQw+TFt57oF3V5h8s78MzT0fT/p+RT5pn7XNM2V9mmCsySp+UE
Exg+q9Xqga3jznzplHTBRCRHjPxY0osvbYXW+htBxOQwZuK+KAEe/FetcHwpiUda
guWhrihLTywh9yKDv+poVux5on7Vd3NcA5Svq4LLrGC42mmdxlwbPbcAe1SA1jzZ
qbG2addibd8vJrwiXID1uOO0pO0FQ9128UmyZnuDFnL+6KQHG1urngtk5XfA76yD
XLqklOXj0x6IcqJKMDYTvThOBUUVL4I6Vq2+//zh/fP7rDxqQoRRpvPcsS9vwsfh
m6wbhhXja6xClfP/JlsQxqYa6JsEGLiBevuS7Jms2T8mQpRbbXvpojFAV+juvauW
bjYFlZJVm6n5zO8ZZJYEUQlMBADne/SRlUT4OgeD1n4NdqByydFsMWEkwZ9g5ipl
/1Z/uT3klgOWuWgdnjzPXYiliOAytxeQQiwSXe+R24JbeJM1s5Ym3HYp+UTy/8w1
tgFcx24UbSBWd0kOzGOI4R3R+fVpmoamxFYPi/ra6ZEdwB47T/uwOC6fwWCFDIj1
rp12FDexqp3xVRovVdQP4v0r+Vph7EgGaR57BlYBjcxWVDLiCOFPUHPHk00tw6g5
j2Bbu8lyMkgMy1m+8FGMP23N5sXCv08yBoU1yBXZGw1uFxqWDtjB/a0HiUU2qoru
GfKRX8pdq19dMDX9//nYMDYJ54pRbjajncMqFlgZPp/ngFj0qb9Xfl6hfbVlZasa
r1ZheLgp367JKoLqlkxkfyrwS3Co3hm8RoUiIfAtj+nl0LPGOLPVs+OntaXK1Ryu
4hrBjJmpIo0T/nUyzhR3IEic7yUc7BdAn4qCt81Ag8CQbZF2vPGKXrLhZKFRaCLy
Tqi8fe0Y0t18Guxt1SxA5LxtiR5sbmuaJ++zxX9o4eBeDLnLJkWsL8u8O7Cf5D7o
4g52cHjjgVM73aS0PjxIz3RJ4CSoebztI8Br5jc8QGxxK1yZlQMauEdUEHg2Rxe3
bYIzof4mNjGBN6ZrqBjSJpeEtYR+gwLCoVxsImSAILBE1fIArERIt/OVqes0LX0d
Si8BjVUDk7K1TfuB0/ebC+sc3u1b39BZDMlkkh/L59VxR60GM9KW46Jc8TjDqyWf
k3N73t6c8dt0thEMNyeAs+6O27kH8LPlPitlvEw9gf0tKKGIFnUgsagz8rU0RYW6
4DscTMb+Ers9fD9rAS8KV6ed7WCpkWKyzcFCNPmGwaqLAheh/Exf8nu/5kVlYMpC
2tm1gai9Qfuvtf6LDMLenRWDubjG6OAKNhUaD+bzKC7SQx+JBu3JfWFgrqACNjX6
jB0bJ4vlkMIBTom90pszac5uUp5f1MaUqNXSto7hkJib7y2gcDSRvLcgbjq5MtJ0
v/m8WZgTsuK3yvKHUM/Y1vTtOSjSgvlPUydzbE4LfPlDQg7aNaUmZgDc0j567nDo
+mGSnEM9zENGiza6Qr9U4o/L92oXLJ/qy7yc+Q5uhxOpEK6o0JtW+fbQXNhy/b9n
LFxHSGgkwNeS1BiSrT4oNmWtkWhNrQJwlMLIygREi7HsaLbCbHA+KSr2wjUgtQHT
r0D9b//18mmlJ5/K3/ri/dN4Zq4bd7ruFc8wzORPRsSzzeufhpTPndnUhzht/bzq
Q3NE8+PSQpkxbqgpam3SnrGrsLX2qzpp7Wt67w+wJZ/32aAreO2GjxsgsSL9dkeu
LtiXbdQqyF5xtMKgIEmv/k/vXmxKMBZ2AGFwEdA6j81x4/BnM5/rf5SnHYTT1AwI
OPaKL0mxTlfB+HMJykLfXV8DI9F3Ow/vmnJsnX2J8DrPG4vTlwyb8aW0vmj9+SaL
vhSaLLJr6dnBj8JPKzXN4kL4VUKqbs0qfALD7heESmoW+KJwYMCYh9/UYf18pstR
Josp9CanGkrhB+P2ghxSeoR9nw4LY9BFEvlDMesqrcgfCHQoV0TAf+pYWA1n2Xif
NsiZk9CiwSRRqt9fBKM1LBtwjtzrNaV61QpSaFfBs1wBmHgB2KgUMx3WCwrh9pHi
lA7jnwCLlv5l1KU65XLOTCEi5lHL3WbXf2zfa36gUPEjPELeDD7ixki6APClIkJd
rRiQWlp3NxxcNuBhyr2cz69yFym8xyfnUtsXxVeDmIyAh66zRccf73RxmFwMx5Ki
+c0wVkNgKU9rRVOvBR5NWSZfr7eed620i19JcluVtT7XhxKPFX1u+zOsC3mzaRuP
dIq9/i84X1DDHqskDabY4gwCX1djpJFYo9uWbzkOqXymQRDkxI2zSk6GV9BGTkCj
vwuCpA+nSzD8n1if8ax5ibMmCcW1Ki8tcAC8K1oGA4zXvv0P6vAYIkqfLbL5Aodq
6/w7BDBlmM7lC6RrAfiuwJQK+JbnhFGoCUiSZo2jAw7D8FOQLuSHlkNf/voUSNO8
QTbSRq0Hi0P6mYHuMyIiwjsdpQ+Xdq8w5V0M3uZisqWUpI3gcBCFrvx/i+X3m62K
5GN0UomhM05O3anIl2YPI6B9JvFr1+L73IxFNyrMUzrHKuzxVvd9IwgiEHYiImSA
3a7eHAD5rOwjOwOyb1XXzq+8DY+gj6J0vVJ1TtqC9ABJPbUitsxyJLTOh9hxDkOI
kAn8RaqLZGsZCwVTJWKHRb2U8NHS02UKkqW+kTHvaKwmTRAihNt34p8YKjVQM64j
Y1CWXzoceIYJODIZG/lXHiJYOGQ1mEdhvYbg1mLoOC9WI8ayOHYogEdiNKdNXbfd
yYIKExfW94/7Yfmuo1WVVZoCFdPa0deYqfKtw0oFQXmSZSVXsE+2j8gxUWySB2EI
u9sBCgkvyco2E8kJ8a1T2Wrv1ruMUTa5N2OggScsKM42+V2AnoyQ+swvfgj+xFOr
erOEGPAPfM41zykhyVSOdRueV7u3C8swFNPNMJrVDd//YloQM2F5VEZJGj1QcfOX
ipKD28bbR4gfGqrmPsb4f5d+I40POrNVIaIz+edbKYlzZqYlmOgB22iB94X9lREh
KI9nwOh86icbqy1BM/hfQhL1zDuriOT/a/AoikNqwtaeyxTz9lfEkctGgq/0bHnv
wdAY1XEpgUFNkAFI72B7yOeDOqVfGxUaC8KDVCh2uPJmbhyAUhyMNPQXEgWTj0gQ
eO2kPQ14flNhs0F6/1IwI0wHzlzIxPD1SbvmPBN1KnhXOPHBfEBNMoXP2wj6BHsp
kwz+b6kmvhE4X8cHi7h8QRsB3Secvbu57Lpku7bZztjFsMVs/ug3UL0y4BP0ZgIk
XmwK/CWZBp3j87K9+5w/wCMo4S7dVeeh/zaOMqCrEW/8n9Fp1YaU674ZzJ5NCJ9c
pr41ak02IEyv4xE3NZzyBvvlKWQKHl4JuQr4sJEUXM6qKokHbHxnDpGGZjWOeY6u
ivWi0QHwLsPqKIlVwo8zE2gSA8S31J4SefoUHH0sOHYxLJfEUb8uATgub8kGapHB
wUgNdlLdsyQiSEM2/cU4R6Kx78PWlPvwZi3Z9xGd1g3J+1AVlW7zir8jrV0kFdPI
ppsNdpwCdI4N7WWUyBw7V5B//yw/kYXFOVq3p8BV9JaYtOMiIR7+fpqehljiPAn4
sEQPeMfspNn03HJ0R3uN8eRnNkh5cjdtq85E8d5QtlYtlnsU+/FL52/DISsf7cpk
a8jR7GM/4EeEhnOHejzCgYcPIjiHcT4d9ghqBPR6nD8AMmn6xd/11v1dh0rEnfr/
MkK1q6c1geYbd8x2zCXvMy3kUbOQejMtbscJmxzIDKQIDu2TGVRi3kGVNw8RT6+r
vs6kq9CxEj3mfSZz0anQRalm0171GMKWjuoEhox1p+lVkZEYbaiYxJZg2Jh8rFqY
tPl6J8nSq/t7hWG9Tnl9ZbZMreazaO3OftjVxL43WRrT1YTQStwgwwAMHGrnz1bz
QMwXSoGHgJIwAbOde9VlXWxuHH4WC4r9BtiMB6TmWftpoLCtofAb45LqBaQgNrCu
GLP3fceCugXwRNmAt3hrp5430WZIpeLfbJ1JW3b+8IR6Bvu8tmT8oYJuHc9e+Gl8
RS6zVwK61s2y/Vp2+hTWIJ2eCmCdqDtnjs7MV2vV1W+tebj87OduqrGjEYrh50bc
xiA8+yET96sC4NTivkejaVvmsvKEFN7Kf3yG5VXMyPOePF66rD6RAuFWPhanmdhD
rYoG7KesJN5etCvjg4PRTpD9clDbc8c7AZk1iGxUiHrxEr6Fsp7Y/Ubr83I+jdfG
rMECNrB/mdpW/3gldeWa3c5/brc/IjPWOQxNalbiZ1wThdeme1sCaRykfTqEP64U
v/NMWgV0s06+D9lcxQbYvAyfcvGIyhUees23QaNF+hSKy8gHox05H6c3/16hfDgl
msXtjkeDj51vtgTzOKx9MCQsAyj4Fhm50ggt0E4uHrD0u8Eha3eYf2LIk+EmR5m4
g/DeudDVawbC7CwID62W5EMogWuMq+hgbHAa488fifQo5E4gnLxzSurDl8ANCk2v
F7VE5SVdpIQY5F2Tubzpc9hIW1PehleiU7an4qKpR2TpNldBsJrstcXUtUsETeTZ
D4kjhj/DHzTowujzEDftuXTO5w6fB2inqLGft9yt3fCkLEkdbGJYo4UWbw0aUJUc
lex8OcW0V7bSLr7Kz4oh4cTxkivc9wvDTp02OpN97a52mJt+H9wKTdHrnVwC+zZ1
ivXXsfZgK+jlb/8JzMWNkUansMaWExnaI931PdNAs8DJK/ZRIBO9Blwa82TSrIjH
FM2cjWYnriVhsG3CXDIUqwnrlzFNMQry8nrjZmmEMo0+lJigg4Hi6+ScR26olNfq
9+PpTyvqNNCHgx21xWRWqYISFJQsBAMb9Ovs9Bdbc6Xh0BxEOjvLvHdiQZEE3mIN
hTnstabpeShNAVHFfC7UMbhPzLHd1LDGBldQuR82fa3/trlLzJHGIl39j+wR8HeW
LFJzmEyiMD3QRwS5OfdlpaLmosHtpBBcQ4XDcLoaHb1CanzlZMJW9m/Db2n4ZZZE
sHirNrGEFoLMjG9HQejaxMyrqoReM1YtHy7glSfDdF6bjzhtXIpoTNioirwO9qxi
V99pbxP0e4sZ4LXYJfl9lSCkGRsA/nYcVxLV2CDmNsa1Wxwvq4urYwQg3OasoQtb
0k6zErLy5bNx/duFJoPevi4acRJ/Z/FKJlYO2gFZXvYFnuhEIHXjnoE4/PoPEqdI
T2aXDzw1J4RiwIiQWmiOaGLH6F/HASf306s0o8VdCtW24NyiAPvfAbkWDrwYszHg
hCubcKBXKJ2fa7Ump+2p+dwEEwTwkmsXTUazB2P5QN2yNHWkHwlsAtONvlIlHPpQ
XOUZc/xzWkEFktGqWm/oi2Cf3SslBkSxOtsfB+kxo9D6ygaNXFG1RMVkaH24wCnG
hU2xdFoG9/v4sAB7RcLcbqv9dORA61wcGYODCIJDo/yCoAdG/a4xC9QyhoC40tkg
JI9av8bWSRi7tu5L7/Qde4YAC4sXBMIt5opR3/RdiN8lKxI9y98MnQcwz/eMH3N0
2na/ZlExp34kGjUzP/GttN+VjduFJ60yy40ohgudW5/m19z65neQpF7AIm2MUaEd
ciRUvSJartGb2KXLkrcjRAiehzt/nal++hx6vAgzDUwfrx4VEPWgwyj9jNyH3nCx
RzhqDHB9QSiV5NlL6kVWe27IZdUjaUzG09XcsWWAA73uSTqR+VwtJQWL//kZA2f9
YKVbGjSLcOOtx22UnDGNDvt7Hrm4crd8jhDzHk0DIJjaUe8ezLTqrzERALmlUXPD
diy2bZ9e5zaTVAL4uGbwtV5RY3qWISRO2+wMZOWSpTPNJFzCYASm2U2n7VgdPb1h
cqKUMjjIMz1vH7/ihuI40Bw9YiVIt5Ft1wsOWEg/kIMF5eMeBFLvaXjJ275/umwG
OtGLRvl87o1dH4zFIxDsMH+m3mS0aBpeR9NbkILksb1SmNkeWOn8mLUGQblCZEQN
7tSQn91/RFL7LpT4IOfmbASql3miv30wAmuHLmjjzfgS1+XX9AWF+PhmhPfXhGWI
FWB03P2TADEumXazWcqDJXoXjDpiwj2HiudtcFoNw3vDMOIrF+8ehLZNw+36BCqu
mr9qOBHgrExpc5fX9VHYF17O2mRD0qlS3S2WCiqEdk/hINdcwrE03D8J55LBt2+c
doBpRbJAqY8NLeCu41wKyOdLbxsl3yOEPtOHioqJLjskTsVN+ra8jdapfrvafqkg
QXxOz98gHRxNkIdHtTpi1GK9Uyczw2F1x8wns/dan8k2L5Qq5yz4Y4Rx1JuSdGeO
v881u8YeQI21GaUuRwnoxuXhTQmm9iSS5BTbUB5/xDbPUzvP7SdneBiPyofPUWVd
oUEqQzqEWhWRDJbj1FiU4286iU3pKEGQw43P4t4jjM3pHrTYsFv9DYcN16/z8hd3
GeEDbU0BsxYuZpu0QBXCoSQ8EPtlEPTpItZAUkYGnU184GlbhuSmuN0DAyVvGGxo
DYRcevRpSmLup3jjZCrfgq6dh5r3TffhVMpY0hHKFstZ74sF8xsF0wWHX5f2acgm
LaZ2cHQaw2Ra4aJbqfEWPMto3dBVhqgI3fgqG9eswOsAFKUnKWiUdNVdmW7uWYZi
JNEE2jnMf76vB4+6XVMR3Dfj1dJLteXn9rjBuB+hlds/WmPl1h19k9w9T4hHmwU1
t4oKkzSJZzdHzH1SSVp5YmoZhV/X3QZt2Q1MRSvcEPoK1BvTz4nNfl0hM3PpenKL
qHQSkz5kRvdTm1MhKS3XJTxZXs+1GEghYy9Ilf7dgobTjl/gAm6YieiLExnQc46k
P2FZiEClcQn7NLXrw/l5kg1Hxs0378X8qSR1eCBh/bRLLKXTkqpC0hf02w2SdtXB
8O3+4THDi2tvvCTeqBba3oKjw71phtJgbWXGIhDM83wWgbTEzihUNhkMQf7AEApB
hrGEjgzb7+7Q097Dpj5awgzUJ4d/0Ed0OPP9lz5zV5NOmoFxiElqNjdLNF2bFtwG
wvdU9uKKGoybMNkRbbezTOyHbexrJ9uClMgtYRsedOskd5+Vib+qBf5Ojxy2NDhn
GpICJIxlSDgSaYnNKAnV92YEgLTK+gw85Qi5hvCy9eI+3WW6/jWr8pufxBb7tlzY
spMEs8YTcnNfJkmUAOW/Rg7HdKdCmO2E8q+IftBnmDjgvOt9T0mVwJ3pW5fOGVv8
b91p2NNcVqUGQ0McTa6p1W66/o9A1ATGSsHqAipsluDJTItFhinAKLd6taCt26Mn
A2ha5idZgyooxrRVkLpv2NYpddho3nDdlYQOsPqfH7Nw9ONjBC39CxxDf27hSecO
fL7s7DwGD4a8bHh/2LIQGJeyp9LH2iEc36eN4oBGSfiBnGSzTnPo09Vn98s0Oidv
vF6OEE1KmNnHzQOh+/nB6RaohcLFXhFfHxK6D4lLgbXNPAQfelJ2tYNIbfrNz3bc
Ql8kwlSjqTiMF65e4CCDyobfqd8j2dg+3KN/k0zB1UbLIcPItxoI2TIMEKgaBTUq
EVegBlz7SWqukJhFH85GYwVl2pq4vXBEJpE8of0vp/1W8Cz01hlvwKbaa/w8liuY
Lnt0RhV7BCkS6eY34eI6btFRMojoJ4gxS2tdjJzeBy0ps9zCcMeICs+wiup1kfks
NEwqhNyVFHCYpJ3o+yXDLLOdCFxBsAvu5ckmPJiHnh4rrbuzaM7AMZZue3T78ZuW
I1o/gzQq4fp11HfbXrbjKGjQxkxknzWfpA+GWfGRC+E472uukIwRfbzv+mEl/4Uq
VRZdlH9zcSGuCQxG2Me/O73EjcQRegayHjIYVX6tSt2tf5uoVl3+bJp8WLtrilkh
xfCdTTLo2jvZo1W9fausjbf2sFJWo4hYtJG1JUyQLhMkoyK+RjdZvm/Mf8tLZznG
xWQeysXOSft42Qp/La+ktXDRv7xocc8TFXJhfy/ukl1Bc7oEmKY/pGQK4577ocjL
KTU5qjU0aKHre1KFH+PfKe2+rJSI3T/Cy8e8htXn9NSpMsMuAyQziUM0oOMOqspy
E4mzr7xslzy7wO8WEO41v/QWZ1asgrHZE39A1MSG9Y7UX6hPjtx1K4FLeWPziUfk
61ZsleFeWG4ogBVGZrw9vJtETaTN4sLv4MdH72+pHsXR2iDijNYjEXvHpMaS9vwC
rgv9TNv+nBNJ1LoizkccHnI6tdnCx/qqsUepAma+8bCmFFj8D/D7cxe6NTAeWN2S
jqbzN6KGONmPyYDor5MrpcHNzP95L/fPoFEbxuVToZp8rzz7RLlkeodagdedOGLG
m+HgsydOFTEClUalzV9JpokuYqm9BuqtDEEPiwwrGFaviPbeX2d1rhMJa0m5MAEg
tbhqhbYhgNr7Wk5iG8kZWIoSBsqD/Gk/hi9TVB+VN9nv8FHi9W3OkOQ5YNcTqdbw
211JWO7Yj13Rs+4UrnrSzph/i4iRiaiPJ76oKwFQBcWk46I+lSUIZUF37k06Y7l6
zxiEpw6hQIDUQXEONB/xo7fli6nbn2Hnis1leDdYLljz0wB08vNHxva/XC6zvRq/
sFtDDUFhg5yKnFRd5GeIBwMBEZcvevfMMxRiQAil0ryD4sR+oNQTyeSRNTRzR19o
qg5oDS2vH3Yx1nDQhC0uSM5qKGgGT0R3X2jae+OWZQAWt7eZ1AoTlMPW1xO9nYtx
i7cCW7OEs97tsbDNFn420z65C0a1rbiB+8f2+7bBeWAtiJKLIZGANs+a0bVzMTfh
UVLDUUzElm8f6rvjKW3eNdFsh/bILw/BeAeDcE9ndpDfh9wRnwPk7eo0/YPxH7XB
nl2FVd27AZXa+y8eNYCmlSyzyMZqxrReFMSB3seU7jByyyJlCGrGeObGJD04jJIE
dKpyienxTszlkjkyOCvHCV8mWoYghY16O24Jk2iP/KrkD9bH+UI6vwzCr7G9kirC
H/Ma9e3rR40NT7yixHnMtavXAKDirr5wBd0KnKawNpS/jom0c4cjc33Xg/UBJepx
s/ac7qU9ZkYoMKqLP4RXovKhtrPYdnqsk+Y3lbJQ1iy5bXLwEv90o0n78UCLGp2n
qwmlnNdCNWG4GfkZ7yRjDOOp8ahUsKYCRAUzqO2jHjzQEniCidt2t0zxcKE11l2e
2RDsYClsD7Bzktlj58fUTqLE/V4pq/KOdvIpRbw0hxPn8Cp8pMIBnso5kmR6Xpnp
Qu1Bv+LAerlz4fm8MAZNOdPVoQMkU6XYd5bQnj349pfEc6q958B47eA6sFCV8tYa
oo6dX5By64zXZ9Gt22dGNkvXXBEdLTXYZV2c6fAuWWZl5IOF1HLKhIgpyrZ/u/s+
MWt+QxIXd6/XTvWH9jiGTEO/be/zM1vfahrQ3DxdKq4XScX7+ANLQDjJzhcIkKk4
BxnsivPPt3gNNVJxa1yd27YLNlous0mG4+ygpUu69wvpOkFONdVVSrrHCgahfRUC
evuUDhXFGHss7sCyTSI06s6ocQHNCIODXk54EQmA8DXnHCoFwXXp/c0RdEjHzhCG
OxdEEuAJLWdaFElJg74Zu0gF1siwnM+vBpCxmFPUpBdrpbOTJIqH2io9Fx9CBk4v
XveS0IkBkyz0DrWe6+QncJWfaZNcr31/vYULSVym1glRpReP4No0IuOJzwpOI2Ja
b25y/9wcFFgVS5WP1f03n9wD8KK7+UOSg/NqdpNpjtrCpqavMBdn8CannEQLpQKa
GPDP6+r8zHM40TgpL3mAmA1QUZcPRGER2IwApqtyoSvi7evgQO/BZgoDokrNT/g8
nNux1wuK0aOSMuGP3ZIBQJH4RoYVSZSawiangMDju2Ahffmqq/R1FBheRCKI5hk0
OHwtzsMaE1l7VvU8s6XLilrTJF2LTklodo2VIuRyLF5k/r4NL9uEqn64ASKIUGJ9
UfyVOivG71cWj74/Pj+93WbDPIQJA0q9dVuzVcqs7p4qlPmxbiN30XbSFEbGGQ/T
+R97bbeSd/rEkAL65qOCyyb0Px3+wEQmUZfDu3zQp3HRMBopulglW6eI31rpchdh
qv2PZzPm9hXU88QF/A2l9datZQKRm2f8nc4qviCuTczx+5YAyyUoSNNJAyLxcsrQ
NWkUv0/2GRk57UQMScR+U2eI8mbPFElEUR66950NcUd2qNMGdKurp3DYsll83vLl
E2YMeaCWzXAEj9PL9L9mHdoEyIMPUjnI9QnG0PkVRtUPgUMCNe/LHpoXplPYpc4Y
DvN/5TSVMvD0lvzo4Aoh8eKFV8JR2JvPZOaMtQZDcMl/sFugmByzuVfESdplZgTh
7AGuonrEokudh9pTsh9j34jhv9QSVZwmlG+zLOJVZD92DHcECCMjoBUaaSTeivju
QXr22mlFI37wpKlw8Qxub33A6Lk1AVPeUqeLKEAQxjMZ7VvegsNR6u/zHhAADJiv
Os1fbCPPB+OzPvuw5tiYD0AuGl7CWJxAqtcgrW2wqphAxpv7lm06nheWLPHFBGwv
aYKBkWqGCwhFuUxToNmXmO+tPtHiENDUvdQ3IHq9urR81K7G5wdMittiBNZH0LQd
M8pNRd2UVOgHvg0K4oNjZebA2/qVPbcyIh+Ll0k/DYW1CVaR1As2W6MfEXR3fEfi
+kyaYhVo5GuEDiMpY2zt/3odLdFWqEP46sEx1CecSsTni8d39YkorWg+DhoFGPdz
MrQOjK5ST7+VmfisKQEEYP/y6LyLADmEnV7lJC3AVmhVF4egnoWpzzuM35DYokx6
ImrysNMKp5PZGbJd8yZumxkz0JHk7IxVVlLOM13yHcNWzPgQ0v4F+S34joMc8/3D
uVbrt3zcn68eFxa+/V5RYp3qPKaDip+QBSIXzOrPDEerp+lqTdyUbgRT3vwF9zSv
Gge42dWdd+os0cAcZKeZFuVZ8FgWs9OMCXl5gp/jghF4OYQDVg8AUiik+IK5m3QH
SISmAx1sKgGkzIhSQbFoe21j1fBy9R91rfS3gZCD7EvBs63pOgfxPAr8wV5B+n0g
B53kf79vR1bjR9FnL3chhiLU7mEsUVAufoMdZ06R/WjiXZPBwXcCKRIVONSZuPC1
x8vprD3MnlwW+Crg6ifU6/xcVl45bB3Sj24YwhWtiob8qn5vntWCLY4XVGfx4SJS
Zvf04V2pWpn3mdBpVdJiZTsIbZlNhRFwWtMLXhDG1P80Z3zPIr4fNJCZsJRwSILR
cEgUTBo5cSfrN4oBZpPUstTCP71eOTMVbm/rwncNmZlscpCDBdzW+NCWk9nBqj21
dE+HgcrTkdg/VcWtguS5kDnvoEfXdcmqVp08pvimYdryUnsBOiSR7oRjoU2VDYds
QnqbJEUnU5njqQY9MRwm1xbk1Qi3RFzaU4xTohFOGUy5uSofz3+wvSTSZFwYDrbj
TwnstkJsmSK0MGp+BrIh6o0uKAeaWQYB+sgHwzfMaifq1D1O4oxgkeodmr6HlknX
77l4M7gvDw6aJE6k3Y/EeLhssgIRUwSJSie0Jg2hBfmaqvhzRlCr/oXGbvdjGLyr
ZAvp6Rp3ioYl/Z+hWd5iD4s1bcwD+4XyGI8yA2AQuJiIu+Zdpw77LxyaqX7P7S2E
UBPR5ae8QY5pLLdVD5ELVXSf0nqZOkNhWBSBW4K+qKXTETtUvvNCcCDMQG+Un04q
b8lB8tl3oxiS/e4QnFHa+mhCf3JPh52HNrPgQ3JJBeIScR5plfl1GUMcIjlunQsg
Jmac8KQR6BEQWQgRdpYa/zYWslYeFm6P7WIsmGwJyGABZsi+i6xPqcR+/I0PXHbo
i6pMuRIos+DiOoMeTaIdGnh6T//STd2K63IsSdWsqD5undHpeX0CvjxpYuZ2tjbv
q2ObS0FZ5W8KaEP6h8sIDNnYajX9a0+tNCY21Mwso9x9g9vqCm6oTMgkyb2qv/x9
ls7naKy6L6WxzH9cXa+gl3D7TGJGpWJYbKW8Jpx5N1GrfE4idgMkHy3cKlbEkX1J
iDAv4kt0r0C7dQMpDdFD01aOauyLZvJ2gAOaI3pM3rxI6EWtVP+W3gQEy/8pTdnD
8fhUvJEPcWZdlbtLwPQZdmVdt9iPb9Pnk7QQdrEw2o2itPRHLJkzEypBqNn4F35j
L13I8KGk0aPjTYB4MWoT8JWk4an/5VtxSMo7oSfVndV+oYvyShRWaIesTrDD8ayu
sw7Bs9GutDLpGrox6g4MGKk6uELctOTKeRFcY8qh+AFb9Wmf1uiGqdANcyL93jEN
GZm15Hnf6m+PAL42W0A3lswjQLDPA/y0h5/eWvJjB/xTCAalgwLn4rUXOC2le2cG
a1TNpQOgGpY9mn5OvndSU74aOdeTXDDMNg323WqzNGECIyVnBcLO2SYMdC0egj1f
Z2c3EoefGUeuIqbhtL511KIzY3F3dRgOxpxjLLAoInPZTSE87Y9Ccd8OQH3QTBWr
I+eoZ8QimuhZasR/tSJKfXwoMV8yi92VTtV+swjeSTecyMB1ViXeKLjhpyTtlIaV
Idc7wYc8aaFpLo1Bb3gIAT1CHGdp8zni3GTqfamGy3BMLZ8pWFI3UrFRsVuiB+m0
/oITBtNavYL2grkI9fAylFgNYGO+2KatUICyFTDZBB9RUuabi4W0g48zCKxh5vX/
3PvkqWgELVb35BAdgJLcBwsdkySydXDyQ/7TCrxnqDHY/mfHHqpsrFatMGhJxiXj
DSgFJSf83MsSdVky1G5yQNI5Q/D/e4gLpnT6juR5pjKRBCpt02hRTHI8CSqV1OJi
k1iWMBLWIrSbbTqznOLdQeEnixYlgeekOXftVyNQcW0hsJBJgKjKoRNDFwYX8TjJ
XgutjJTSOKN6MZiSyw2DfgDJlRJC4e8fO4R15Q8CxBJCOjJE/iijj9uMhdTICd7M
vVSSJ0test1kScCcJvbEO6XbnTo3uoAUTqFDiOP4Kl/pzmggEamfI3ub9LKmjv1Z
E80g5MuHFU3FpraYpm4bA9VnKjMOFA6FPIzYBte2nc8cJq+fsuuzVdV9/gNmuX2p
euVq+D5h6o9An7t6FZW29IdhWQ1aAnyhf/KFnHb+gYdKKv3OhrbIGaJuayrDESV4
tob2FIRDhjwgFAn76F67mEqtyQ2pHGyb6Hf31N+0vkTvFN+NRIXcsuP32f1cvz/P
jWi7sWAGJV1w+chlR3/35OAmwENGmMwz7xQNZ7VTs2N55JXe8btoVwGUu8qrPduH
7oChEKQx7EUrzM2JBXRYEud3z3Z7V/bOGNSrjfFbFrj4YhjbLMgT8PrxRmwHmBQq
dql1NBQAtX/9R3jAjV8+adNd5qCUMOHpoF+duE1zNLaSaeNCpd7pcp2xIz+HS2kW
/E1niC+fmq5KqQKXZltLP/3EzjjkZ+F5TjNpysDNnchOr6N7o/N0krrn881SGBD6
2xOnWKzVWsiPcCrqkmpy86mmL6ZTJdGC+nMFhUmyJlVEmhSP9SbOrUYyYxJAVzou
313mJlOtPmplC+03YJIsK640Q46XuQmY7c5lXcoLAvlOyrAj+Xc9S+iIBbUoBMFU
kWlVVXfJ6jvoTyMs2QbboLCnvKM0uCsUDuI1581l5UBvGa7bLHz5QVeNmCqd5I5a
GgZPnDIbSuP+4xmuSnDHXfkjLdrrdDlIPG1jtpMiCLsgsn6bBeoWq2NTHuyM82la
W8uH7uNwb+WvaJSIFCb7qIuMPb82z4a5b5kzVVADLt1cxEFCuhBEJCbHWoxKvAGU
Z+IUVbOxQJvUT8aeu8cFGbWg7D+c4/lhrsq+6h2u9Q5MiieMuumxmeAe/uxpSRPn
CJxF8US9zxpN6EcNNO3KffXu8MthqVm3pImg5eX2bQ9J+4kkgTcOUbERpwRmlLFL
BXtRyYwegNMAJaqk9VT7rUfEuD/mzvqMnuUiA9MeU0mvY/7vkEUyr1GYJAT0Audh
ciBYQXwa9lKa9vZ0oNgMO6clUtWhfD9SKo9GCGvv2vwiEq9DdKmRYDRtLjpg4KVV
kLaz+SB7aoo4CJJgiPgeaG52PqmZLVrkWJb/DXZiBRM/E3KpJ3bBfH4no63NHR6G
NKdfbHwck+O/RjZrKH2VmnsqJD6GG0trzTs85IqPWYo3rcgsXVPRbqFUedZpShT2
mqr7KQt8cHR5/U8gKs/pZdOGYfp/u3wERmCbDDX00R5EivA1Ay9ERcd7KAWGE0L7
JkceMUI8Ic22JOg6Ljvs7TbpnnaXa5We1awirgOsKADhNIguhfLMRhvIlvGDN4sI
58lR50fr9BQFnP0QpPhqpseuKAWswhzyPxog4QXgVATNRQgRCwS+kFLy0v7Iz09M
0eW7cDBGYlkZbPzg0MzVXCNV7t+NlQZXpSw5weia1/kWQ+5w3uUB9iXmkqG5OhH2
Orn/rVZGVZDaa93pG3Ekc9MElxPS4R9mzPNU2fKnZYEjf9zz3f4VnQ5YAYLnflqZ
tmNQyT8fXErtzZrElvUcDxHeqLXpfJK6KB2lgEXvOJwvmQD0c8VOA8irepaeO3Vv
oZx93n1oSOhLqMKr1a7VxLDgIFSnC/9q4f7QhqgA0FfsVCaOQ0ZbqELDNFpZsav+
0Tf+Tk64IrGw3CFpJ/lxGguUI799Q0oAEl0O8kYsI544rEOKJLfu5R1LPdVMsFnA
2wQX820MNY/iQ1Vynv8XQc5iSVpBKTACvQ/9vEf3g2gNhR52qD8V+0LM9/3T5+Qo
AX16qQZNvBwUs9hGcYYVSrn8hAs0qm7J+ZrwVRKdkRujnimL9MPV8oLUl/yffbp9
Os9V4PK0VVowuQ9RsW6wkfZOcoMZeNILAHKOJK+Je1hRNWVe/fiuYASC5tVPmBXt
FvtMR6kHCHRs+aNyWGvc9PstrnqPqx5MCBxy4r66SIMe6TB3EdmI6E+jiP3xvucS
9FpbCs+VjSwlBmtHCdmkuX2K4rOw5e/y31bA37+3LxpBXg0Av2cgpiKLr0bFp5ic
rHu38MUUHBEW+/PUWY9+57LS/1gh9FafOYjChkwgX1Ny0WYeGtVg9rv1YifXfdw1
Jp9ELhk54velRDhZP1bFyWZbkc6cFCcYXp+mMrYNGh+1UI8NPJ7dlA4I6NYNUaib
ihSzJ72YkE1GIj4h1nwJbpzKAxeQU1G7xfTsVpKDLZN+8c/MfMT+zr6ODUEjH+s6
fb10uJEdAoVd1dSyBPLVmfajJteMNReCqjmFGhwPP0F2aRJho/nAZYf0jh3YY13i
4AxDVu8hkralajVXZAQnE5mk1bBA/unGaviZbcO4iqlSF0FFFpWFeBItyRwB2tQF
Q4Gxpjkxrs1kwa+XykPOG6hHbFqEFnHOi7wXf4RyI5MO06oUZ9I/pgcN9C3I9idn
qnBvvGF0WOxBTnZmORg8IvHWI79pTdxsarHIE3gixwtm3lpm8nCAjG0mcq0w48ie
kcEVcfpMmygWKVYQeULv4SQgwwttSbpoT7q5FrOw4/OUw9xxU7kcewB+fcIWqfuT
OooO08+op7TWWHcgD0wMbBm824CnvAgXOtPJF5iTF1mtPAWQVGwt9SU6oWpBv9U/
azetQH1yz5J+iGPUKN8mxehNCN+f/3HpXMKGoD3/i1eVrUoCzF6dh+tZha0ofU39
IqNDXyFdZehY+q98eZUKkbuxHlvKpz97vvGRfyCrGENR6OUBFR9u6wkPRPmPgLmy
vXnPo5xsFSWm/GzCBIyUQ0skIa/X0NNH0rJz6iMpDeoO2VcyxQpCHnDNgpmSU1nF
4kd0PMLUZx11rL8cy5z5l3t9cxjt7pDkVAS7E0sfOy7v2hZwytPCM+CubHZhN/Ox
zs6BObulYhcbKRl/qNv1DhileeUKqtZDOP7oH9zxumvnyznEg5zZV1OpuaiAn54R
n9H5zcJAODv+FUNfU4ksMojuxF3q2bDNbrJUFgTvTU8W3Fqcb07v3Z2l7CqO8zB9
rpIwe9GzAxqHRP/hc7oh0QoUb2eyukBzsfeY1KdsJDCccV/1cRUIBfpDl0Kvb4W6
JkXMaeQyjackBVtWi5G6e+uzaFiraQUlAEx1jREeyf+4Lj0/7SWsNafQBbrR4x2/
7Xda3DwHDexD/JtgBvu8zsrbGdgWDoNjncBwWiWEegtzR11QhJ439GidRYjHb4pU
BPtn+8TJjxkdnPZXvZavPZVpg6PJZFo4ZFyRPv5BfVmtLGUxsVm7SvP4a0kOWAta
8jzisrcWxgNI1GT18NgFtImKqGgNNepcCXKQnptOr1ziiqizKtwV0i7ijQmmlaBs
jT2nM4l//nZelzBWGuhPi0mNrow6dW8qyPULihxN4KwdlgayXSLswdaTLt1g0Aex
Mt96kINvfL3cN8Qd6IEwYBYx0WOiaYCdzpxV4BCxspnFxI1lMTHbjNs+QDbrL7fq
h5OGtV6T/D9sxT8XETMzyUp5sCkgwme6AbDwiVE6WzEkCbdWMgt8yEYe1TzjMadA
tVS+e/tk4fuVehd4+BfQCeHkjfpCQcqSutR1JnS8YWmJjXu6pE70L7Gpd9+aaXx6
PaLC/M69bEKvw/vJc1qZVQ5l1mEDIupvjVEdNgF6vRSfKWsqbbTXbW0qK2ITJ4ib
v4H4xteulI3UHpF4A/kd4gI4XYatNMSh0UfIHOSIf0XFXkXdkPBr/9Q6D36iKK5y
j3eJvJ9tKmSfHS+sdF4rFExZmN5N4IFVaSeb+YCwPSOrQsaJ+IdH24XQm/Z2hOHj
nI+5nMQfmq0qx2s1W/ivReHP1UsX1AXbbXX9eQf1rINxolFfDzDHDNAkOZMNMX5+
7aIzlx87BOVAtkZXu22z/MqeJMoGoL1Ux5hZmuj9elm1WMrrSq/3xjec1qED3MjG
EGszr11q/jTQtC0AUi3XWfFB7QhfmC1PdJUPPiPxTTSCXSl9vKGqycSS0A1WR6WL
N8FTUvRxoRhQFLWTMlZVKjohke9FZhSEDdZUthrXr/bH9Qw1Xi5gvLE0jiWdgU1R
D2RRIwTDYbvLHP29Nu8jWA99hZ3sWoaC06YejINq25UQFx9lo8mMKEv+QGzoOJJK
EF3HuXLb9fvQpiqXk0ui4piqXI9vs3GxAXBJ0HBxCO80zHqWtVtZY5YdiwCrfc5V
IPmW56Xyg1I88xSVM56mr3z56rq51OzIQcrfovf3vgwBgMqRF1Xf73kDOLtZnIEA
JsXBHHTbh9g9moOvigIl7FdpAFFNdVPtW55Y0uFbza8y9nGwi1OmjpfH+2voINy4
ZKP0ORhh4qQWb0X+nwBnB9kGQZAM3pzV7XIAm1P2EuIx/1KKO8dMz87UVLX7ULwY
YV15eVy6zyuBo0zay13Dop1AEJynIEr5FWOt9Wugd7JgR4BFjuvuhyqMi6M6/JXF
LvKFuzwjbYGvUmwU9S1HoxtOYHqAjKaGxRE1kWIthwpY6letyex7aqKjP2CbTr/a
r5p5HZaH3cieWFyTTdzMirZeWzBnr+Va48LOYF9zBnvdtKspmv5yk7en/mBt3qDc
Qn06YzGtBUpoY6o3bDqoV/29hLcT3e2glVINJApHwy0DykcZpiBaAYJr8ofjmHvu
QCRbzJQRmYG5IEnHCrRhv7p+jFd4kI5SAb96l66tnPQLLhTQKNFirHW0qRYxmrpe
N4MdgJlcR1SKdVOBRW2LxxUw1d5rDDEUdjoLsRRAw66IhBzMymy7hF85msNs7Lzv
Rxkeg0g3OnUB0HbAlwU1nrxLHVpYOu8+2Favee3+JDHbfUa6otCh0o7ZzGr+kZHv
RP8IN5p2itzC4xp1eSdaWL/m4fYv8KV+5tykKxcJRLfY3g666abopIM0xk27Tkew
AlrxWGPgwrVodcuJoYFkxygOSL4ksGjgO+gXzszLwrQeaXXABzTRjioEUWCiMdwE
CPJF+oF3B6KEbRajMXUyFxjMhcPWhrdJ82B1qemsNpBLsb2mvuNDkjuP2NJZWO/u
huUo8o9aYvRLhRllP0ahRCVUWwrtIHDOeAGALfDf8Kh9sDCTfWzAPuPK59pGFxZ3
f0mS5NeKU/RHoIfNlhhppUeFlGCJ3XzIPsQfdrY+H5fJSjnBxWxDS5gwurswjukS
wBA8EtkGy69hQeOTDENHQJVTtN258et203lgxU7WUjVVHIw8m34p0i3zaGLiDsLU
CUihmDWLoh4nscd411jrDgKQHTtk4DIYL4XhIyRZlbiKVKSRINpp524XFwLNEb7V
eTT4ucsDY7jcYmUu4QOjrcIDDZM8q8jpEGC0muALvl1mCyGWuYXfW2zXh2/QjENz
yYI9uqpqKgNZ3pV9nNu2zCHtWCaDJYxdFzffNWU1Gbci8lUchPrX2NtudsWvkJc9
QZBJdJ38X1BOqmK3aMYmpsqajUQ8nBNmezrM+HLG8FqITgMxmihfY+UOPFNXG3rc
0nA+ntz9yS5w3BJyFkPss0jAqzandTHQtlKJWnkJr8Op1dN+nbcv9pzrgi0hytt6
xG0E9+XvAzWzL+jX0UgUQzjS6yLOserQBfmdSP3646BxkF6c9DfCfWB2CBcpPWme
/J0S9tIFrw2vg7EH1v+vjlSKmNS5TBFPwqRFlFOxFadl6IFJAIDZc0kc79mb6Wuz
ZMUJSRQnj4Bv8MlWnR8K8WSsAurq5CDvG0Ieo+HhvRGY85Bblpf/EaoPdG7cUk+X
+QdRHJLiCrXkzaHXYEevtPWQAyiUlpjS6buDGB8m+2XEBXt7DnCkWN738vMTyEIb
npOTK2KGhJlNGBIfEM51UKCdk4DobqrZXj27Do8cmDAbEBNbvaxwzfIHTOUYINqT
3qrivsuXnBM3Zm60JqkBnCrD5RlmNh4/p9YoF+sp/TUBNLHtbpGHxCrTsXylRhpd
NTWMOW9jJ9RvYU0lGoisKuOa+CrdReFQ+xMa+gpKC+C0FTFxyfpfvQb4CYfOrEl7
0Z/AvitpHTkODianbHzr0HuKF1tzxYCD9HVrhvmR2i9iRPR8OMrcB3R8iUr5Ef2A
eHatxuEayCE6UVVj3fSuvcDPvFBIdyciF2EMVTGsF5lGu2CMMrCrCJ8DncMk3n3V
ruswChtE3tRCr5b8Ke3RdAqTQ7d9bRDCKFyN/IDXS4lTOH0NYrOPY0w4x6hkxSal
fPeoVUw9D4dwRVu2UiOA/mT+cYjBYypdPXnJGm+f2ZcyocHXUAdLgebBAD0OqYtS
xz8n0ovqT/ukqQKzD2bEbjBTUygtnK0feDrboD6DeVs1IEdyrcu8vUEp1RysMjMH
mBFPOznu4Znvpo01hz+mgNT4PRG0Np008YBvx8GVnGVf2/ueNjyDjSro4mjpX0h8
tzz2Y8rZfp7qeXCz7+v/eYKCT/gmkWQ9/eAhAZPgxi2hkVpEFGOctSeCGAePEsKG
/o4DLCenwqcYSC8M9L+TkY8NufrQ6Bq1pZmRhYPwgY4xgmhYaObQmI0DbI/kNqXS
p9vJmCLrlSC6+1fY6qJUlzeRh2sgFpvDXA6lAbocuU6ndcD6yLIW0nfOq4kgcjI7
N/Vd0IIkIWp3PZJThLLIlY76VNXvdzD7hoKV6vpiVi50BQkO8U/CM90x3IVZEPAL
Lx7jGk+I4ULCSukgIwm0IpsIVDLvof+zzhYjlpqig6IG92rnFC4P7BUIpE+HXQsG
wYehYrxvDZBMzyhiIpj3J5obSZ4UE8EYl4nr9cy7W7bgrfd9b5cgE6+MM3VX88Ju
0EgVw5X0QlDZbtdB4/Pp7gHphbbJHWHzYx/OoLwBJpu0NwhjUOcw/XPtLMKtmd8g
OtAwCoY9YI81+pxHGleuHlcqdNtTkYtNpAFJcqGAEuA2UOsZ1IJWVWUZUyfvMjki
uDwUXU2hMsyqg3buNvdFi9pbqc82TU2rj1MIN8hUGSoSWdxbtbekpJ6K+usQsXWI
eksjRAuuAaK8zGKl90n7sS4D+nIu1vGRJNL4I+sXIfIJuvGktvzTkAKG0KG5zxGg
gQjALHZAPL229cZOk8GXnWtuD6EF3IPCEFRaSLnodC4OMIK34A6D3zbySpf4lzei
Ln8IRQn24bdrd5tIHZW+grsi2fdMjLVO+oHxcjUd3czFh0do6UBS3bSE+IVfsYX+
AoMfR2u4fzTq0oR7a8QPsCF6WI/4ADW7w6NJHIEMvYrAyvLwQcEbMuZS7pt1Bl4b
3HyKoHafRfqOsgztfLyEhotUD//MQ2BnVFZ1PvnB6Ql1PNe2kn9Bf2KPBJqz30la
V3kGcdYJZ29iGL4MwERAarTIl+t3hvCCh2L7sDPqBD2YwtS3NCbGprB5FPmw1YJX
DTbjShcLabvPyAUmTVCOUJFhQvZ9CDx+wpAqRMYxHsE3xwGefTicX5z3hqtLE8GA
D4i5vS4VaH7aPIz779AbXmZwfcLihAIuULsdxZF+kuatB3oAHsbka4nev6dxjT71
y7miOo9voyiN2PuSD4Z/9Mnqy1W2P6vg15oO9n58H+KIvFau1UvIyG+fpH+cVdWj
5hIgn6gFYXZdFvzV28pUCKnlhy2ge6sBr5xZ4J9SFRQAF+TQq8mBWMny4rxvdwyl
vn0vhrmuu/n6sMgCdw6Jw7to/ZxRQwHWTBjsZy2eQRLC3NK2Jlw2WTsUsEyZF1il
IzdZz3ySm09hEiJ5mGeI3kYOG1wdj4TcZAoPvbg/h8/1GWk2/qSjI9DlxhbJdlEJ
rAvhEv2si8HiNys63iODtlXDfdZLDSKODtv/x3BH0yRsac9v74p9Pb71+bPfrFbV
CixS2vyb7Ud0OMzVUW/W7oWFGpyuqsx3s7SMAJSKq1tp5a2qx5v6s969IXQHJH+M
UIA5bpWD5HmyfRRGEaatBj0b7IRooAss+tPfjeOIgprshl7JvhRudWhSaEmSuqaP
WUqw7EKn6/svIfNhNnnf7Gz9wPpDcXUSVDs+0dsCfC8FCORop9LLkS8uGR2eQe0g
qUQPkThdbSr12ngTLMv1MNbKU1S9jrulI0HstBAttR3SmGH/1k/2kUpT1/bdY7XP
zUzNFERZtZQPZnoMs3+na3X4bRU7HyiRapXieLvM75ahGCyRDJuft6rmYXnm622Q
7URaAn+p1SEkCztHGMQyKZtXtugkiExJOvDtXnjR286nMS/+NVCgBRPhEluiYgvr
c+6DKjEDGpxaSQa6K61iBl+AtUveboIbQ1DImC4gDa84cbxx3gsM5rEax7o8wSkl
5ZYNV1IsgR/r9mabtgaMwu1vPbKM9A6KvqixBcxVyDqSbp8VSBYS1XTj24O/Rkz/
ThoPDalZJUHHGe4VnylHsyXD1+V/4YtOa1s7ABLOJFjMmE8441PSbj5PltxtLaZH
kzfZCmV+vPx05aYirnC0GNdGebqyc+GHc6snQRMQjOFhCljivCv+lDssGDHhgsrk
oPMPuuOb/yVCfBVQ1ui1FAwfnBp6SEcM2qMULNNvDfCzyys2FuTd1i9EMkT0PTKD
Fv0rprmaOaDrvhhCUm2jT3GxCtabpFCJicmjTzsTFSoGeVi6DdQ+WH3lVZD60R/H
2jQ4pUd3s7ZS3ntuzhEkaFe1zDhcWjU76yovOzA30bFXWNIfioeXIz7XQqBMZmu2
c4A0FdmyKK3YwaDHIVFAU0eyiwo4lDERaLBZqF94uCg3voY55rYB9aaQ+4OrKlB2
3mytijSTH7cxA3maPX5NUHKfTAdNCMlJhGEBG+VjwT/HeV0L/GpyPsPOwNoSgWlo
RQJKumJ9KjBcH4c/XD+m3qKpwy53Zjej6yipg6U9/SOio7WokM8TOw2i1UrpHXpM
N7PMpC7QNofgjjy9ZlsBlG+RCGHfR+/xh/worPRXbBMl+8bAnfyTRMR66PseAvr3
TBjpgCDChbd+YIHjMQQca7I4Rt6+bkJRfDCVy2AyI5zhksRAQxAbgUN/RxhNoiOH
WVKQxCBNtJo9jCgSwBBszlGAyI+ScQUX5i10+tl/j1hChlN+P9Ygn59DI3dBb3/A
kFafv8yIZ0BbZNq6MEmAR470SR/nT7Ulfh6irPCVe+r0nPI9aYReHNDY4uwjL0lZ
NlStZxn6sVoZbQUZXlEcegCgUnHHzLLk3XWiC86N6vNHQhIN29c/JifS6yjgruhg
Go1tEa/iI5j7AOdcOM7jDOc+YBojNFfBBSxpuNlWc7NKE6jHn3hXLZ5kvS0l0Hf+
aB4VCJgAVDWOxvlsKT4MCH+8qBAnhdvxgFVaPkfpDzhefH7GVyqzy+uKqC18xZmK
zFnIwO93G+gbQrlVYbQwe15xvGMyC4bbYVeoOHMSb+0vawL5DxbZczNAT6lVHYDL
PdW9G9qIVpXVuN2vA2RzdJrGzuZmAaV/7UC+Tl8unijjlWHPblO9650dhgqlyORt
8aaQi3cpc2p6RJKK2cQNvjjTVg8OuOXkye5RUY0v12oM8OV47Rn7Roetua8kplrh
pOaqbjZcKPB12eSV66nkVWzF4LAZiGFrAfxi2etwWqUUFvKrL4z4Xl1x9eVXpfOo
z1GP7xjp2huLtdbVSVS4dlLCHJO1i7qxNcmuJ8DJJmYB7++fVMNOyGp8DLLNE4F5
198GKjR+rbT5MHiPrJHudFdOazCFoPaR74CGm1WOxxLsCRG0KWYEQJDP1xssHLF9
hqOhk4AU+I2X+XdfRoyKVK9ra39mcMtkbqe3y04ziOFxw+w643iVlhcqwW1LBnQs
W6vd1fVx+gn13hr0iC4tZPVCsAufkkBFXtrCjCDBS5PKc6G8tvvCx+K7nanwxS/D
ZIaK1q82eiEZjbkKOKNxwb4hUsgaB0uX+SNlTYMfEYhzNROFPioPGR5IhVZhOnPg
dP2NZIcTeZ93MLxdJLwoLcT3croWhZmkdJplhumL1T2x+jMH9ZoNzFRGYPx9k+vJ
QbWqDDKvb5QYaR5WkCmktRkheil+snxnaecg/MNoc++hDiPBCyfSmw5bVCFTZdvU
tqNANBi9CNcbzirXGzAroQ3EMynVi75vLyGW6rjHJd40i/O2OS+cZp8Ef7h9yR18
7v/mpqbT1Kb80wmPMT4yvPOy8p7EoXNDGYyh34rLG4LrLQ9l5Cywf4AcBI47Aa17
h5gjrVhnt0wKy8pm/zBNOx/Vor1kgHkqjsS49KPAo707AH6qUDzqn57k4ZeHxBXz
FusRrWm4PIjqplfqG6ZIl1sq99cFH06rJt5/j+2jowhcu/4u9nnJhE6oih6zT86o
SnAKII2wMPJ4dR+mqFquv+l9RTTIFFIVPzhNPDqw5RxDCxi9jneqglMjOXnQgQMS
O8C4A3TRe7uSSM2dKI+tpa9erxNLsc9L0rbvj0FUsGEgK1NCQixyPmXAtjAoeIyE
WonG1m5gjwT0oEaw4cIJ9X8iRqzH8zcxbE5jv80B7rRlu2uoHXNtxVfU9thUg0OM
SLH/v3xyviBmMMOAY8gkqEdWf67Nx6E3ZISkbNC4MF2XRsshNd5W+/riJ5gAqKaq
Bjd2l2zufn+EfzquO+MnzDKEhBlQtHKo+Ktqbn12geo4+o1ApY72qbq7ABxiPoLF
n2lzVFcBkBsPymYwABSNEhBP1e3BUU7sUNfoxVJrZrhruYRqlKbElOtCmRSuXfDO
cDoYIGq1C4pR+tamhBMJURfW6vAMbQUbt8Wv6hkazM5cuo8PXLADiyeu+NWg/uHs
1CGgzZfez0fRIAFL6UJlONtZtqoeZaZLpM1BPbZh37o3iGiYYYjaacJA3twg7+AV
WidJrfiBxp57m5JvX58b18ES+kiYtqU3JsEEyrlXry19sToaHMZ3KTLsxYyjj87k
Rg7fX1zXe053+D3wGRF+yD4s/d0avwckmmWeC48eyyMhTHneCvfYp5cwUneXmKkP
gy1KDSQjta1/VuTccoKNpdaLCNeGO6kFO2D5ZN3V2YXVXhGevlrSsTw9JDCEVU2r
Kusvi/R0uyFnhpf59AxJOF9/A8/bwhEMGObO0sEzPezxD9xGfKWMTkFBNxLrtSsp
SaKLIgSf82JmhRsZ/pO8QAPtkWWDp3p0DDpSikqgX4ue/0WqB3ttAefdpjOOV3oC
pCxoTHHTF3WTYYKQ4mI6o1NaW3LVJEWS4Q0knrWI0s5WdtkP7ROT2JW/Kcn87Ftx
CWl9fLuLpko8Lw8LJOiloA2uK/2yRBvggtiuoZdzbLApabLIFnD6LuvztYQA7g7B
C8PaKgcVznmF7z8kfKmkklMG3kFf7viYcjVc4lzFw9sY+eSpZd5u/WzZK0dTB8P7
YlWJLqD4n+r3bqt39NolljibVIMoyHvjYUFGhPmuOP+CvP4HgJTEaAAuH7aP/j5y
0hMs3YLDuoBOz2f7dy9kdvvw5U6oN0+pREOBer6CkFR2b9Oi/WL6kJjkO/H9mVTk
c2WC6MM7BewqKoCbdDkorirdK9CDWDOR2KgafuIm31FkuY69Dd+LQb7PJrF0PvYq
S61LI9VaaooriZ6AXMOuqYxoeIBzvVivrq2X7aLSxmbYoUYHrZ6r5MYq7m3TJq/h
n6GKa+Dm1xGkkLyKKsKLPJ6De2OEFDSKDCapEWhQIoeWsL/M0qh7zbsemY3JtqR6
N9oMdgOBnSUnV7rJgGQqv25UvUpDDumqSs6Cm6ObFwqOeu6xDP0TG0YBLKJhmH5V
LsrScwbOdyun8PVotaCgOkQhijut9Y8td8u9vnDsFqv3p6ZvfoVkNmJrg9diqNfV
lh3qc8Bv+qy8ftfcB0wCeZt1PvukdBpqqksZQIAoXiJNU25OAEKrAhOuQXbCRF+F
7lMiC22jiQDQQ2mOPqxcNbEH2n0s/KFZaEMoI2J/sigF6pZBV/zEvLK4N2aLbu59
SFr+bQJSLioQJ9CJzycxc3jikElN3WP0tFtvOwqQc/iY0HDNv8gF19rpcubVRuOT
YKbsR/DW1EI8+bidBkGEiM63Rt7f0BCgi3Xm9mELAPVDD2Lj1yNLrSun3muZX7dl
cdf0VOWaM+KvvJWQ54Vce0otlwJLLH7nS3bk6OfmpeBtzdCmVvs5IXuBmVkfrFSn
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
JUVfuYJJTRI5lraCf7ePo9t5voPhMWCzCYZAlKqwb6XVEsmjW8SjSZuBx1uXotMJ
fn8r9IxZYV5bqqo6yr2mC6Sl30EznTv/zdQXRG5NnVb+XSKPeGIuuSYKcYzXfCRD
DBWkjekY9jiFdKjDqxAxCp/XYGvYiAb2dSQo5WTVsTU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 380257    )
Lyx7nSyFnSCZqe5vxLC9nYYzBLnhKGGiaov5OrUY10M2NgY0YvNsjV2qfQw7euTh
GDjM119EjA/mJ1XBCIXJh3W5qESib4yamW6BDCizy/1CycjirMopFYFHStTJHFMS
1HAZ3DlcZ6KxkF1HpMufKnYRO1MNl7wNpgjxEa3BQ6ZwIBhfoddeYEMjNkyKdjm0
RgcG06UYb6iFrY3komAPCw==
`pragma protect end_protected
      //vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Egd7PhydEt42glR9TPRnSkYpncAH55mwTWe/qVMpmPSk1AlxM0LchSzADVtjYFiJ
F/fgJi1+597h4SocVn1PP7bUI5UTSUwdzw/NDkSF4JEspWmWa15mti/G6EuxZyn5
eFhcrlhey5tLzkqoIo1AzJ9dBLXpcH8Id7pG8bwXrrQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 454128    )
GyjtMW+E6ZY2zVXeByz/b88p2lEg9Vj7683zoNWX9Ezvt3OCiIzAfj6UvX5VWNdc
bikVt6K4rwOz3YAUgA4bVCC1dAEMkPKVW4NrEVTU5Ey4lBkYMVjPc54FD2BAGGWu
d/LSx1bwSZrSQTvHj+SC647Hw/CvCZYtGHI3iQLtbgrFemzCiZf7nC3rR8/X22zx
gTtW8XbLS243oZUzAjbYT90MEL+AnU0SzXuuFDrocr+dqfgGPGPvrv/nBvit5KlX
eMfJf55ODHqMDf1w5yRvw9i11/VU+d0gKppe63PIXR/f73dVqhewJeRAutFigJIA
A++8/foTqxVX6Nt8Ghq/k39v4Nt9MyFlTEUBXKVquz0JGvXgxtlsqd1F4zRG0+k3
caB54Hws1WXEn+3J+pglx1GTSxiXUFwQNchUjYGyxfntYAqPKFSn8UmMvy1jXPsr
PiHfalkOUb50LqfZDz/G8A7Op7XD/Zq9+HI/cfyRHHfixZrc+Mj8V1HUSwCpuqsQ
N5UIUBzeuVC4VUybWQv2ZnAXhvFYwCVUpJGGke7fUsCdXh0o55T55+uhBYQMK+OC
AA5xpihHGnoT8tqLPfmfVEn4j9gHbSbyHBXgQy1p6oVxqgMh/BktMCMrddMKDKIr
22eabHpA4hwnEQLll4brR/oCBiE3drpj4cr6Gj9GACFhtar+ZdbFYNl5znwIagVx
KwHN/LCxcebHKVkriZhS7pEz/71otIy1ncai1KZrGQjqO4azr+4ZZ4wjWAodIzxq
nH9O++OkkoWUubwC6LSrnEkIERthtErisYLNbngpKkqPlC9Zi6HgyIdM9Ctu7rtI
MSRHZpsZDsWIL1zZVuFIXy+3w3G7ilBbLDtYkcHqfE6I2pXdfrwrObbiEn8KJCzq
1xNQio/7/d8P7hKYTn9gqeLX0v48L5OHXXCbYzOxR+RrGGgJpONLfoaNnpkT4QWC
fVltZyxtfTMlXkzb9xV2ABNw7UeuxHx0qJSRPTkPLkOQQdQiIn0n2f28xnVei/l0
QFC2yMC6Duo9kwWYDyVC7dhmqPnmP00/zAopJnymOlGoOGBZAr0BVM1v2BI1cWds
3CWEfY90m4qRgzM9itG+pZSsQyV4XIx5Pj4vgQ7fGd+e1MNi3xTPyTScIG4BYdeG
oGti1hT1nFInKt4AC+ebdKY82EKDq2daH6+N4fMbDHC50b0PIhs3cTQWNk8EnybA
KUeBstc1gBudkNsDW9qu4nxLywKdSgyI+CXRYg1vzG0pxdyNqCH5ZgF0jmrEVQYD
uvxvivHRf8xtXmeuFr/GgAcVCqT+VrqWHcEp29VUZ10TCQLrAc4Mx3SPSquCChvq
oC9uBBB4v5NZNpO3YBCSnZcODA80AATm1xuT1aNkyk7MRJuNAmt32RtT0d+0r1uK
8Mxiv/ZFX7qPziRrjYXA52Bo62cB+Rit5ZzMelKzJANv8SyAow4JrIenG1kWZlDd
ZKtt0AkwQVO08uAh2t42QPmhbAd9BQpsEb3Z/tgxGIlZeauTyzkN8Ujka+yX8eqw
Hhh+hAY+htJGh+ibgv7tBpKzGj9L4SIfkoGiuTo2fwaVI4geZiUVT2JJGBeHK/Fi
T/ZMtUAQIVoMMU0z+9gBFkhzQLUnegayMkaqIHLV0EoSjuKchFWD3q3KjDsfp4+L
35ohpV/HGUZ6Q3PKuBrk5SmG7SKZPaVxwgMBJPY2g8edNfyBU73WFy4gEN4lQi3y
DQEb7moysql/cZykCTRqWwfWszo7nPk8XbHq6xgSrGFPenuNjc0tCuskEz4tftVS
PzL2otqjX0puvcCTj0ZHOmRW+FpTxv5/QClUP+luxHw6jFs3qKrk0Zt+51/1QTeV
3MMtg03OAVIvNNMhMP2IPHEJhB/H94L/FcmgVWrVxrv+jIph8OhNlCSCpbNLBJmk
InX5xits38tUU6cWFW6/OyqP8ywHFlzI2Dq9+/Z/ZLlagX87PNAkWutVpejWPMDd
pdnA+k877LfaEfdTlW784qtYNlr6P9o5hvwhrxC0IxtYY7SUL9zsnptzrFkWRxG7
DSmj3QbqyQTqS/OdhSWzz8cQyipq+QbOKPvJmhRRnpylx/VFHRTg5hrGzFCzVDlY
3qZ4XL8KjS7HyPQ6VMTXeSqTEC8ph7ki5EncEk7UULBP4UC1RXNUn4+9P2GDHMBz
lyrxRWzLun6hXsEBDo7RnUM4Rfq/4y0KHJvxOZgUPYx6x3VzvH3jvLhe7/BzMOVf
y0UOku7xtuCIb3lrYH47H8FFj6vJsmmoo6r26PLbl/Q3in8iJLfmysLXVtEckV5J
xTaSRxDXD8ZfrV1MHxL1S2z3yRbW7HycDL44AQIIYnhSnJGPaPV5ErgV3J1D7ECa
ayVNKYjHysW6UxQiobncg8/1w5ZLtgwbTk+mRu7c8Wixxwvsher0MjxIk/hoJFL4
tZrzt9j913ECVpUHZ98GR6ZYnf6+bJDN4xyPCbkyswqVZY1OaaDBLWwpKtBrCwfb
SSDPAMee4sY1jTjaJ0LInvFz2LaBDj9xODHLmIehnnZxIcn0LpTl9BuLhqoAjcYS
YGlErJyOYMfKKaCO2w+Jf4lZ2x3pfzmkNbwegG09kt07LGWfJtaI1yRD1AREaYFH
WHp/aiGMjg1gwVZTmuOMx8yLhdr6YrxdNZMUTZTqtgJIQnnnVT5UBAz0F7uXc0df
5h5CcIiJEDO5QcPDcwGV6+zkhnNXVu4+DfD8/CwkV32QmqYb+IZsqByTB1SzLQ4F
dywOZN6dTrcTHvJFCW6/zyynarlU6PqQF2pjZDCxv0mygR4bpNToZ43yUIfilCEV
4FW38LHTbBQbSBkfZPMf4igZoKrRLgbHm8f1+xtWAD6sZ/CZs9WlqDJ19ijpV+ln
KZcCbfTIK63BrN5KJ6oF3aMo1S40cRfkIz+KqVv+2+CjPmxzNwBC0n9kn7IpH5sY
jugD/MjTFk98ze99++CVDNT45HqiiD1VASwnF7grVSEbajynE18XlV7nfRjTX5hH
OoZpvQNaSP6lfZ6J2gZHfCINy4IIEIIv3EFuHHyztoo1d6NbHNl4WcCzCX4Pc/bZ
SCmtIvBnkfRAQxw7+MoqxOaaVZ2UWqsUcsOKevtF2eEQ09UH/fWSbXwhBo1651WL
rnJhZMDf/8AZKiNtHuYrUqSXs+14FEDcOu7GiQ+DKx8W5u/3OgHku8J+AzxXcY6U
jalfSsZSD3wJxH2oOucwv2gR/THBfs4BEK/2W8u3r9OVQZ8GdTGh5goew23Y+5h0
PkYzOJpYIEq1Q7Wkhsa8qfjF4zLjG6/4rieKoj61Q1cLgQDSR+DCMo/zr1D+5VNJ
zsL286C+KbRNTvWI3NpwBHM2znLuEwInAkFGe9mxPbSb3CvLv4pVybyKm7eYFqiz
watHhgQhsSm/3P4fLZHkoS0qstje+tpvtupoSXpe9+//4P3PbwnePOtCgf+09uzJ
AE/xq5P/Fu7ozBknN4zQZMgZgUb4EFWTltmChQ3uLiHv6xWD7nSN1Y3w0DsgsHAn
0QIk46yMIynRrATgwnTMYTvFmiNNXjKEwHFCthD6AIHzbIEC9QguwnIL0tPO2rEa
kRUXNpjFNN12UXdMCo73URPhRlVOc8PsDfYA5eMMhbEhw+rcm8oNPR0tQBTAsB/T
Ov4G54SjzjN7RVsMoGj8/qp2ETtTyjaWCWQ0qHZR749jRTGz0rJD/ZEXW9JB2a9x
HJBgIb+nEO+ev+gFJNf39HXieWzg1iL4HSC1OWVsDRiOo+T1jGKirkWocARnDbZj
0o+NHjL1DnuRKJssT95jDOxHqFSVGACdMAcgcqDeeR1Cna2cv/zZxDeUWorAdkPB
fU5IKTZJfReN6OOJGz89sOiy6RiI7LSKzEEWKkB989+0goh6IEtQ64zWoG/W4iiA
VIr/SrmZyLMjow2T7ElRI0KWFtSpmEb/MdQcJO0FkOKpbiz+aGxoHY2iKXp1od0I
VGqe3TP6TMCuZzpdsHfmJTkX4JoFxqqtg34yVEwrd2qIzbdxO9uWfAXXhapxRyoC
thXUIatiquoYLtw26CVrS4A39zejC9/B5iF0MI8noMLqnJlzesIqskclB7RlDcLe
+8uE925isKmiykxgiKFw51744FcmXYmwJ673ibcBpAJjvF2ivGsrZmhF49WFRXcq
SiTTXD+d2AwwoPcOvFPVYKgNsYwXEmSc5hwDKfHMol8ddOE3uDASkZUPZTBI/JIw
TYqJBJPKXGsQRsa39co3NxsXD7irGvfAAGK2o5lpOSiLsGOKHLsm/MjLosNLFkvg
7fUFAalWZOpKBLlh6h7Po2kALnA8sofy9VAehvsSOwRiJvFKaikPIKJXzufX2rS1
SPyEXObjb0HgDL01MEqgTtZQeZHDYjiWw5Si+tUDEGnKSeh73JqtuOluaGxYNlJ8
SYu6MQ2525Atsg/25pY9gpIptPeQLThksjE/fVKAD3lUgSwaQQ6HIAd+vpCKgtxn
2WFDMYnvnVXKcoNkNox1Xorp/d/59fGq4nuqv801CAEnf2qk9OALQVr8/4iRc5kq
Iu3mXaFsMuO7Q9ZhfBenFeOaVBtruXlgeEs31XkJ1zK5IjtLAU747aif9o6Biant
VaA/bYwTtIkeh70dXZqJWX8QnQTB7QMufhPmarXM3XDd5oJXjEF25gtuLS7YrClU
6j/tUddyvgghIZSpk/5OmIOLS10zVj7Exi/aSkQIHPtmYk17xhyhyM6KqivV9UF1
af6a/34sadbxNNhRT2Vo4zHFgxNj6ZlR14XDtbAiwQnk/9c+34l0lKuAws2ovDBu
J5Fzt6q/Q4WSx+t3ene3ucx0Ag/olzZA5ESNSOSgBffmJWXfM6eAD76Ka4Wr+DR/
HJJr9K4/M3jOaAQLlU9mc5FJ7RLvdHXhBGeQ7towLBDj9FnA6KvZOihW7RDvSzOK
lSy60zw9BLqbX9xqJqFdXvTQcpaIs5u/hl+qR5w9hwrWgkxPmZmb9AF6YqBJFYvh
zco05kMw8eWD9P2DbBHQJWtG6ZoGpkZWLPZx7l/nEIwipJik6K/c0AERZGPHzbTT
n8NO0KeDu33M9tOjB8IfuZDDQKZD3fqFbwmWKNpm+R1m/B/5NOlJ6VcHaLdJDsKP
k47riMjoWh3ZclOmcOJzUCJESGgXsWEmKtXPuGkGtgbOYDKqCXKXtQTlPnbN+/lC
mW4UzeYgUZrkJQSRb7FL1XZJSvNxs8dGAYJgnVH8X9jy4VV7yngjqNs2VdfHkDEb
c9lpIEMcOADjuYg5L1fAyfQ3zlc1hTsz/kGrC9imSrqGcoJyendDwRnBGBXVmoSZ
a1/IoSA3PL/nXoGPEDbAbGGt19CHuj1hY2j57eY5YBh1Q4nSH6lvvuMfXfjQypjw
c8mXOUU0jBkxrgAlkFecHJ+Mezv4O8F3FCPTOwYOS5Nw/aMj/Te7qJVqkoWglNdR
WXKcNhq1mX1GHsOg81DWXZyoykD97t23J3AIeXp5YG6pvMpDaOwn0YrNkqKsrauU
zQ2CRCnIrzA9EtlxZZr1DTLU3L6P9LngI/fBqhF7zx0OBs9B1PM6sjssP6+vV/F3
ioyuqqOXJm7W7VeJE47OP3k41N2O22v1bTEApt8sHGOclk2rqYMXnydlFEbqqkBF
aHuak/kz+L90BbGpMXF+e5KmU+DgXttRsaumjMprvpJf2xsoyTeetiL/Iv/zuL6k
aAqmHmRJTvRDDrP3RNEMORqUEQvdfYOjWzyw289QeUAZduWVtgMsE6fl02bCYELh
pshM2ooGdP/pA+m01lwy3T1/sWFJobbLCzkgmfWmtIYxjBTa5yhnwpEy3Gt5nIbb
u9P+Jl2/gnaA0EuZdsRApNnpn1/S98zKmr0f8vMJiumaCc5ZPnCnTqC9EDIk5coZ
vyDVqcF9SPUJXYiz+75ym7UHQOH+1XfDFl1DEUq0kLBrzj0qh2VtmCC9mO3yuFfh
xv8qqRnNFUYn9uyAf2ftjR8MMPQvJ7OZd9+x59H/tx0w6x8OIVxOX/GLBuG86fqw
XRLjHswpmUqYe0MzKeXesWKkQkqvhgO2oBTFb5ytAH9avMXAXRneAoF5sJzpHAaa
Fk1G+WcT4Kb2UtFqsn6NzeaDKAWcdbITIinwlcI5xUEFYB1kxbEtxzc19ZHr2loa
+NkSNciunT36459wXv4xL7C07XeMV1JaCM1KDAd5doSull67HjI//zPGUj1H7awl
J6myiFbyh/DsBk2cEBOgg8xrPUSEtNxdUaalvsf0PFLtFzpu+FWYp8C21ehmGVr8
cF02GzIQrmCj/52dpHI4Igp7UmYmcy6hPn/k2hS+f5AYIJkRDnOUKdtODIZOT7AH
aUCXIc5xxXovh+6Yaq/KQ1YeL1YqexWYWYXkBrmYa6qkwwdHIfyp1XVYSTwryt1k
KHwuixlK6CHRJnp5k7yZXZFBSmxgMu5cvtIWisljn3AMeAkPKgy16W05lWOwqtg9
28EOnEHo6hUiRDEx2cCRba8VSiU5Su5YddYDQHwMWqCNdW/dlMfYp6wYKZ2m2Mde
WA+6v8T0A2JK6mTn1Y7PmTC+EMgvWCE76ldJOYh/icgEFtk4uQGKGnCAaXBwCeiY
ntiSFHEzo+mSZWtyeLSVTyzJaa263/coKyM8lR0w+FwEfo6jUiZwRhQjB3Uz1vKk
8ucJ31wgPxf8/4jBjk10x/v6TY5H99k9q3SFx3/ZVVuvPbC3meRgXf+RRUU36SLj
+kCyRh8x+TCeBhysmDBp5PNYyJlkslj3WDjDVd47WLfp7qVMK4MdMOlC9fhzZnkm
XRtlMyWWUxLProdlLD7DZ3Y2X9An8BFpSJwbqZec2QFzSGhP9zjEzDxh/qnOGQjZ
78T6fxc7FJ5cxc7WItvHNyTlAhCGOpz2zj7RIVowEoZPRRXMNUreqCNaetBBcai1
3MDXMQ3pADvjO2F9OHG08CVPsHpnWx/USIflHDJIivwV7ajEZKBUo2KvFNh/UbiX
6fzDDYMB6rdfCzjJmzNDIS6pBgN1VRaXTWl4XippRv852fUZxYiUpOcWMFx59av6
9ixQh+x42cTeolzGmIRvvh5G5AyjIdvQhUvSVejvVl0zhKUhqBBPHKR4Xkm4ZH/w
SQPydbgoxFmNoEUB1aNc/AxIaH+GF3bkJSfv3xTLE+wJjIyUJT9V9lFi0w6VPEF6
wBv1+DtKoX+zpnHAp3Jq7FqjQmZqa2JR6jlGtzsDArYKEcHQuzGeDSEgm7lnFgeW
q+uLVQEdYRYXPR3z4rO/KbLho5+X+1p8jetSRmIvfw7PLvPLyWePYxXeWuwb26ct
pFy2yJtdrXskcE23biO4ULoO93i/nHBy1RAhUsEnlqpYL+zYozhc3Jik+rFaucDP
8mrXj1zZaTNIKTt1W/4KXsGMGR5t4/i4oon7VmvAoBPegmeodINJ1xBEs9rmIfHg
MEjTb8/4DkbPHzZZ3xJ8NwdOyBoAhdOqcCYF+wzhRG3ZgKn78u7sTVtmYH5wUsXS
QD85uOramVXzmk5jl068bR6lDK0zN3ekzzcb5Hwu2mAIyufDDQO0yDexrBTxz86v
kIs4aGvQhpWgrJqbBCjeynBM3KdCVAFS+Bbr+gukDeCjd9qkhCTDI+h8BNuhCxtt
UqAYIEiQgC9jYrPMp2aI21deZK86zd6VfwIwLvAwFD0ROpVrAOwA525f0BPIngy1
n+ASqUrePytkVc6T/3cn9QDAOec5Wp5K3jSG02GxdhbBi1xQR2R3irhB2UKIl0h8
WgyD7vJC4FdcYhIBu+YJ5gUqI/IquXWHyFEBJe1SsY0YTM0VrPED+1++ZLXO8Rag
yC8hQHlF6t8yCFSNp31Fios+UtS33d7Clmfj4bGTCXAfLLlxHuoQBF0FkKCTpM8K
Hf7BEwBSpgmuCM6NZDt2DYE1I5e4Ec+ctokJiIhWvahcywV1zVwsZz0Bau8/Olc+
ZGMTMMp2eKSr3FXzQeij6VCktl9tx5lZV3WOKa/UzBiDioVLRQ+gtx4H4B7F59dp
oAs1/vLS4rCXYnon+4WeVl4h3zblqM9InZyAaabB+pVA3z/oPPamoCKljl1egj/l
fIO5iJvpAiEYQm9Glrdt4Lm3ITng1Ro24gsSKgg3lA+Xev4hfzEol7FCc7sHYzrA
9+yzb8eRIszsi0gjKIRSfvub95Xj9eSoeVb/zs+Vmk0D2LaUJTxkf7kJWwNWamf4
YKK2c1crulyHk+H1AFwOk36cN/+uvdb18NGw8xtywwx4zkR9ap3pWTAvTWC8rJZx
7zihilSW9ANotAXnGUvXFZDYxUJGVXprq4ZUk4SmelEcNkEJ39A9EU/0Q/GkXtyN
k9wh0jn8qFUJwF0Ux2GdviB4iAo62gyUW3ngWczZJ/3PvcUrpFoA7O8eMsBoJuVl
k+/AIcjRfKGGbK0go2lvpIzC7pRk+LjaaBAj5MKkX9tfXsNHAAXSHhH7MiCvT1pv
tz/W6zDqCzYa8JuG0IV1adXnv3FrEUfDV2bTI9haiq6p/YT26khIrMbAZEjDmKwK
4CZWOr05drDktf6GHqdxP6XOoVaeDXZkvvBrM1zsGf2UpFPajY2e1p7cfF3YaXwG
W5kMJwr1/9yzgkfmj83BkxQ4XmF3Ma1IQR06BQPfWZvei6VeALyq3BanttWHetzB
9hd7jCcOiqRc90lmyR4U0u5iaoxwbYEvtfG6QjB+LHCJPNLo4aCeUhH5c5Jxo8e9
qCk/02a2viv6rQa+b8dwHV7BLIyhOAmW8ThTSxogsgW2b69nKsijjRDLVFIw88Iq
PE2po2yVsyAwLAauyozbBwNAZqULkUXqHeENuSL3/Z+OSc/NRBsoAxA07QEza30X
l165jtKiU0NiUNfKXR8c/zmIHw4PDTJ6hKm/D2Po/GUREAuiXAXWmFxMl5U0qG0J
C1rdZ4p8nnnzlQ3tgGH7insLAs/pCo4D0+mWbZSaRt5nohpImlu77cMLyyES4UQv
5H/FPZUePHIvEkH+G6pfBjRbNyUxFMzvxKF2tnL6o7fIZZixkJ+MIjAsJNM/Gims
J6dW+diqZW0rycgaWWRXiMUfZpdNrGtMo1EYnkEnYKuOqviKbyPp4e0OJYx/8Xqd
yuZ4/lCq6l8FZZ3hWp57EHYkCJwMdCVskHSGnw9NduOQMSYU2iJW58B8t6Rusvq6
YCWqMizcrlkY1r5oSD2cA6K6pk2XjzrNgkLp7t2uBsZsHZUofvNcVCkpzwMbOWHx
SkamqEqARM25QKMnUixNwlDPda6w9V9wtDjUiJSUw3vWtonPtXBgKETxrEaeds0Y
Fr1Drs6AxUMpN4IE0BpzdQobHhFTwFuCHd4j2/87w49FRRcTfqh6ko+Xs8pi/Ppu
/wiHEvDf4ZYG9vwdmIv4xyMUsEKzh4jpmsPGb9rEVb/NE5ToutUcrOpf1zrMMbMo
UI0x+7t11Zg0+6y1AgEiBbNklUEwy0urMeEmQ7a1sr47jKIWLkB7TfwY84dcIdo9
9KqPnMrN53uXrSdr1xrCv7hYMwBog7QqHxIQW2jMD/ZyaSlbQDux0cNjoEWqNZ3J
lbcCJe+lTeEGghDEuLBEgo4+F9ZT4hQPDDpUXLv44+p29F854BNXuY466NNXDH99
j5/vreeu3EJCvIQH/buVSUAasCv7ZmN7TN5SbNzXSKWgC+XJ5sCymYg2CLe+tX9v
oCtD6tDYHRpIB2VDmjB1u+ejb+rlZ2UvcT3Z2DzsBAdEMFAhhQfxny4++JwzkDuj
isBf1MVgV/Ik5BtLBuD1X8FiYtPVkVTD1vUazUk1ssiDgz77nc+HzI7xKhoGx4Sq
9HdM2eXryU4rzcTJL0DJG33cntVALa9f2fJqs3XMRv5Pe4p1sG0b3qptblZLPWEd
8JKJ4YNTL5PVwVXKIeDIbIO0Ki0gp03h/PcDuAERqHOLbO7Yzdcc4bRlKUlaQHzD
yHR47bjydyEdPQQF3cqWq9/1m68sUXjFKSKp14VPB1oIlLivFyXKbBAPsjBO2Ugd
lUJBhPXGYc8dEC61M4jjGUciY4ednb0fL/L5Tu0pqwF7Y2CXcmEV4OwUoZybQaGO
Dlk8XBktmuC4HBAZRXe6uTOzph2HCV1pnnvAPUtIpgOIp2hvwsqi5ZAqxGLeswUC
1OriA4HO1EOei4VEsic11RYtJc8vxD6HX98e4j9LrAOud3y1oZQLVSlzZ3arkV6z
ubqaclVcSjEScVwtDJcKdl4hcbzHBVoZrYcgoJzBkuJkcNRc8gfOCr3TfF6X7C/H
c9PvAmGMQZL1Cd8kcSGI2FR51betKhCjX1MwjFgfUixv6QMW0wPQllH7k8B7mmEF
gFulUgHoORm7rxCGKdP2Q1L5cTTS0/xjzo9vf7BIGTxrT2thWUC976+nPf1hzMJw
El5G1ZVDDGg8h4WRz2t7kVipvfzImLaUaLwBNlfNH1wFZ7miRxa9UHoSVwsWN6F5
EVjlXpOxKXT2W//ww1zJ1l5+qIhZ/pw7EA4HjYLBg1nIJs3kmG9i4KC5TEMh1VMe
t5rxN1MNZgUbsyFod6mb94WVG9buUEc4nW257y2S8OGPok0MeDmDMRjYPPrH8YHu
2vdMvU3aptWZaBjkWNIljrEsbPrCzcDXlqZFk6+PAPIZu0JxqfJnyyoO/JD/cu54
cFlbGD2B/hx7eyeB0SchgqcrC0JueD1uSdfK2szC/8uUccGXknE+vzDRiLTPz3li
UycYSIhkesk1NUVGubSa/Fpzf8+wqkNLPfdx9IfKlMhl8nlCCUOxmgrSrWeQa6ya
YSbVO3dHt5jF5AlAXwIy1JL7ouEF3sS8ildsfkMBzBt/+LEScJ0T6rXg0i7S1NiM
JEP3nArsqwQos8pgAWVZ/D8VPaw1bDAmg1QrOK6KCNDAJW43rP5tXkACINhj181E
Djc2As8h/3r989nisNwSg3hH+7Nv9MSlUjiwcLOMNkpZWVYtD0NygtvNnzqP0itL
xLAIuUpSXrOXCR2+XJSlefNMTKP/PbRoPRVZ9DE4CcdPBXbiycx6LJz4duYf4BjH
wK8ptZHLJ0COz9mvJJxuTrLX0u/Iwq2Lzu0mjQ8G2mh5/phityXqbs2EC1JMJ17P
DuVeE2RKV0rvog/QEKZ/7FC6G8ralnGYerB7dZLamcHq9Vh8DWevJZd3nkwm63YJ
sP/VE9JPaT7nHGFYrRKi8wytKHGv8JUjECmDtvx4kwm7Qf/GWhS8AkPKL4WVCFr4
A2Ttl06Ok7Ltiu2iCnqjF3MLc8JxGuHY6PA2trKY3DWFjrl4kSNARgVlWlSOe4BD
geMnn1ViyIzjybwuSwolX28p2IF6JDF11wN/kTzbMCU+U47/yrJS1KzdrzTCvyTl
WKPZqA78exwEF1oyjMmmqj631rG4/QK1s/pS1eWiXzIjuujWH3vjiJxZi7G/pN9u
HSpw8XjQtnX8DtPyuSvLw+3kWhluI7u3SL160PQEcrbKiEc/bl9YrFr+LTh8Qdjl
k1DHAcjFLwT8RiEScbs8h0AqzGTtIZzWi94qxcTTtv173lPhzHfr+jittL9laPou
ja9O2HZYCVnU7+IogyNbfN9Jvs5GXsZ6Tfly44cqwxNnnhVvdz6X3rt7tR3Jnzj1
D8zLsh5W1+wjfoFkywRuHDAaVlAFjQF+PN3D5inps2BDBT0JmdkYMH7vRBp0F6ga
ahto/PEdLzFISqabw1kGQsXH46OWJDTWi5JAugxAvRyImfisdbu1OlcvJvQ5uJ0A
u1ZZTseMkATXX1c9c5Xqu72PQKQGDFHkqPn1dpR4RpVlg26xN0Jnbukcf3UqT1MV
lxi2YklATClY+vxjlcWomxGVEzjyw7o8NFO4BjKjep+h6+pA3KNQu09gDiRRbP3+
+U5MUrZIqxIsHEb29wbm8fejMHQ7UAV+zpmwZ6HqLxGtJzGEP9WNsEQK9f3pMjdM
B0lvyhOK1XvPMKXGpJzeORXHm5rOIlr6yyzuCDmKBP2+R7W8hNe/cXrOT3fCl3N2
adCdEd3TcrFE1esvWIwgnvo8ZFb4Uj5YtjbnUrc9w45pTgo5h3hUzufC5J+hKHSw
sm07Mhx8NNIMXP9rYsvL0u19yCFnSTJIiecuIRO8l0ccSrjmA7bm40UoDjoqubnT
NcZWuO39dSGirybYvsmSlsR6ppNU2xZVxqR86tPxJaG9W73y3TqAxRv5geRy7mut
EEGzg13zqu9vCePlqvoX7I46elPsSPsSXutDp6UGqXkaC5mcavjKmOEeyx8aV2WY
r3H5ds6XrQK1jWjmby+T+TvRUBenhVnVssarzVJQ+R8a07HKw12jGDstaTyrgUSy
XmwQjTO/ZANVAsNxsBfXPmJG2+MgNc1Qu9OSi3d7zS9JlSPYUYlUXRugNkdIxpQE
0AIEZDFV8BoeLi6kNUSQk+D9F6suQfNijYuVDsG4FmNiBRV1yb2S36/S2NO1q24r
ac8Wvdq/3YUHb8ORAkO+skPclmVe3SUriKh+tyLcYa+vbVAnYLlcPO0ypcHg0v+B
7D/QavNX/nxNfSestvPLnAgFwILMYODj4h+xRfOAvQAHyiX/aZ7v1tQEwe1485Wu
LpkJfQ5GQXbb1VPYsu8XNnMm0kzK0LdxByo469tb5P3IqGJnoOe7fylmPBAnRi06
ADJNajFlHVhCqU7xVJ7cSkUe5ho3olVHhGUs5BRqtVXOr24I204tNgwlo+tRwXlt
dem0r7rWbOJs6c+FXuWlbFxeO/YNtL4gwcioVecivEErzy0iK1lo//TVOcVsm369
A3QAroOL1czjejuFPAPQUCMHShKTKaBCDewaD5hCkTwukbBWKYf3y9GLACc3n1JN
NkQ4D0sQM1RtloX/aVofF7SQDePbVLJuLaxqtGH9DnL4q6imDuQJ2iaHz8m2PaPZ
Z2NmFESCZFER2M3+PXUPZ5Poj8LuYZ4qYH0woHZ/rJ2BSncxZLzo7rm4O4PDXts4
Eyy5Wx+p1vBimNvTqMXuJAGtUTrRwhXrMJOg66TwQMwm/MkTIWUEPGzJc+utlAu3
6QkAA6ksPisADt5RWMDNY2a5ooRKO1imidJAl7IEW23guLt5iKC4SdhNSSHYMc6W
iB2GMS7t887F9wfur2vgqdTNYUFtyeqAGdTYsPjorbQKYHLfVqA2qFHyMt9eYQIt
NQvElM/x/bzVdY/EYcTac9kdDFxYXZr54aTZ2hldF9BtCYINTIY8YigN+m9fgj2o
JA5FkUEtTgU/fZ34EVSdMTu1wEPvdF5tm2ojNhuL0W6wWcrfRVDwKpWF9fuVcxuq
i/d8hM0qOKkih1ZbUwL9eRf8lO5qF1sDxwuoJHj0pYATioRlpcFVML4fEgOjSysM
tWYutjKmqt1Jhxvy5aMyBlDYvC4bi4iM7CtoB/FJXxfiDwdav4ozvWdndCKfdWDy
ZZKJdt1AKPuqksYqcT7aPHpngcDjrBxZspYK851HOscspZXFPycW/nHi0OubfPrO
9V+WGQECXWM5hDmm4QpNP8fMXdyosvYFAxv95wCmYPNp/mYoXkVLP5bw3u8FePhZ
24R2+xqAV/sKF3++Rnt5348epkU4eRyTiOMEMkSOI2KKEcEw0BBI4daEZzlrNS4P
yb0qmbTUGdfMDe+brP8C+FIPqV4jmP+mbE/kczyxqe0B8i3FjbSa3JfzJHqaJFXh
sgaV8N5Q16GkenFYpCxWhVLi9GlLqxOZ4FlsSLoZWBgUtWWnqnv22vjpQ2EotFkU
8DqSwPYceW26mnKr9R8zGHrFcVAFp70+M/qTBoiJI6S3VKLwKIURKKeVCNSHhHTh
7L0vWfN2j58oPWr3fcqSpYrl3wdWeUQ0ylbhiDmfy8I9IIJ0p9XTXkJkYcD7t98E
+ngT8UA06yen50ZdQq6+dmd2pkXeSIr2SG84z5+scjnsxAYgtIOiYq0r6RZP093E
BN74k1+HFcXykjXUcGeAhUkokZ6u3nVRHMi4gRKXWmbeflC+HM8jKc8ji/aGSEHn
22X6iOLH6yFLpYV71k53X3PzQdMRFqna9x3CC+iLU8xxw86vl65h7O21Eh8EY6RB
B5EStXUGr4HYAhTHLjqbdy8KiNPMZDiVrLNRAS7N8S24EvaTKcjPsICOcOHCmR/1
rBdhQjbd7k+WTGmg1ueY0wmaYzizDr8R0JVFOycvnErmfYwiMWf/C86TyqWV3f0g
OGbog4mEBxDpYNopaGMbkzEWI3Q2pgTBJ8Jc/anz/U0fuZV0Icdf3/slMzl6/Izn
kHa7YgxN36F6nRtpzDoC0pDBzLcklwW4SpliC89nQW0QrvqokO/ClKRb3y/ObKj0
MGaFko/DmkXh3LZV1E1rvlbuhS13SlNaKCEG1Vmys38dDeGDHvEa3F1t0uvUQF3y
mLiLic3VnAmw1SvnuE9YERYhtcIrLZfopCkpeSy4VAtwfhb5IzVHz87ykAINB4Qe
GL5CRhXJ7gCzgQzG5WNfouyhZYXOyng/JQ1ScqE0OpWUOSwfxkmtFIxzNaJTxYf1
ZGD8ZmyKi3jCfo42bYDyd9vW+J46+gu4+7qxmV0L/4GBmAKZuO6Qhm/rAsP5IDEV
pDfiFMPdgT8NKUZTqO5F6lsFTdZwXOtXUWIjLkQuYZsu6EkLJVaer8RucpjE3pbZ
M5rzHkRYdnE9icd/rOgMx1cTIihJri8H2n3pmd/jDvWouzW0b7o2EyOX/rA7690C
3xm4nXFMHxF+m7gWa/7rPVAT4fQKX5dB9bHCLu3n20CaoEaXH8FA/I5ov05qim6c
b2J6vOFf8tL+k6CD5m7PssHySQwbtfl1ng1e9IXFFQR+JaMvq3P0BBmds6jds/+u
XbLwBnOsYppCV5Iyv5GyMmx2l/Q+psu4EFZ/RoZUhMLVsVFrWwx7SbYoaQ1ov7ri
GdHgO5XDfO69xIHh6Rqitou7/yIVsiLC4iEa0eqMKPJe6OouPbVtaRhLdoMKz8tp
bgbLoQJOg0aAPpYC3NhnO4UyoYSzWGGxJhf8El5Jr6TTw9wgqMnpCS7gEiAlQypx
GsWwZA7PF0E0YMKApWO/4T/oeFH+xEjKZjxUoqa7VSrJgBVqn8AmFlpEwr6kaiwh
P+K5Vn8m5aQbbFUvi/0FFh8CHh+ufje3KtfwDzBKa85vAw20OQiPhZBoS7M3geH7
n8l6gLXJJbU668HEugjj7MWhu5jR2BFeMa9PJOA0BU+i1ArafC1aVgubwgVlFlBO
E9cAKgZbH5txApLCx4S66PxPEPo5Ocjk9W1Y8qZfrFCb1sxCscOlC+TqrVFBSaJM
yrLVQAIYxkSCt/vyvJznPvGX1oT9W+LL16iu1UuF2ejw3bfJLZqUg7xO7T3hhI9Z
lSR+0rzIG4iiZSydz3iq6qJeD7aI31NVPrnGXld9sgxiwzPXWg2R9MzQyqqXjmIQ
hPEPxMtZgl5lOU7ZDSakhWClYbW2yoZKKncU5BLEEOOabhmdUwPzKR4fpFImicBa
6UQpXoKwCq6Mhix59bn9OP5pnKoyuPBG4F0e+5ORAgCsAXFuAAXSaeCoyJ3K6+VS
T3Z+j+K5CnfU8vLfsYhvgMQIj78r3ZuBKp9F2c+y0x6B+gohDNgp/ZpHB9qffP3v
1o4sw/kdGU8xADDmtnfo+vXkoD3mLgXzTFFxox9je99oJMmHj4RWSDV/Kv4vDrot
bcqajDeilnWgrVq1X6Wa8ZWKMgf+2mgnTcYvn4i+t0t+UijvsLclxlj/OcB6QYML
1Bnt1Gq7POsRa1ViWREzyOWwlDQhAEFMSz/NDUAWEyEk9eIc362lNU4ABK72KW54
Wck+GJDvBnXgfwJH8Pbo4lNLwnYCiOWxZJx64d4F3mpEmjo9Zg6xZRhx7K2dD62d
CTAkmHrEOay74j37Iijn38dmd5BqVFO79t33KJav74udvRcx832CF9IfVBrA/S5j
RNCIIdc/tjQl62loavV2eHUBHE/sSrrnMVRIBPwDsTYANktXvC7Zt8qarpcKfQ1r
plN5gbHZQq+AHDiEYlutA4r5Jd86BNS8kEbCkYdgRmqeRpbLMdtnJ/Bs9nH9S1Ti
39St09UxXGoj+YmoNPbnee8LhAhI87HHd+/jbOJ2O4brKJ6Cbh4Gj/gtekbPcMSr
W0Atnla9NC06cEBtVOal2/INn4plp7e/f3vHbPQVyq8ZMikdjZRsteHoCHHklZqv
XE/uFdJq12hFsvuB+f5vBiFlM5dwdTghHOQSfSZTBi110h9KUFT2EE5jeGgJBf9j
YasvFjm654DJn7hYQi16Ky1QmG689v/poj5U1AiXCiJ1Pc9xjymd5e89tZ6H7C7Y
2+tL6Wd9OKo6qaTxuLycyBxgg7yGhJIAwpxsvOvVHpiNCweeX6fS9jWaQdwHZKcL
il6kY2rEf4zVbNTWGqu14xSc4IlHIqezijstqmIBdBm3EPlAvFY2yxqvGlKYftjJ
0gzIDSdRQ+OHERBJjYGG4jiZyOlvi1GETrwUt1gUQNWCZQaH/Y6UTPVEOhqmH6Y2
6wn4Km6XSkmiM9N6z+Df3JSvGK+NAiM09tgQbr7oNAszNy3XPbUnaKflxblN4hha
cuOv55QpRxCIo7qAZSUseSJuf75zHE8cmpQs15JWT4jn8j6+sSNsq2ZX7aScAlhe
fEeyO7jq3IDdplDu420r2AyvrRfmq3ggf4HQHydNw6rdibC4qcGD71NYh8Slfe15
PhdEUpenOgwSwmJgSdCtrbF3PmPLFGIzGCb+XkMxPtFd4ve9VYef0cADrQo8RAr+
afPogQ0C+8fbPeYxfyMNZDCpWg4ONo8Od8ea3Is4KEjK65z1rpwAKlJ79a0OXeTG
r6KeQqW4zRTzKP7p3k4cHxE2fHYKMKZiWR3gjpfAQSFA7F5yzPw+n9DbRdRp+WTw
wmYNfQYpcCq6pR3USRVW3m2nPkpzQeS/Z+58y8No412H8QQCVX8cKNv8Gosuox2h
sC1eM1pFNV111+nybEYVEeNTyZrBZfFdTax6zszR7UjMyXYXjq6EOPjGiHn91Cb6
uEZRnpPyh8AykMXgd1ipzhZ7aVKlaT/rrMo1Whjejn56jTIHypALcyTYc+pVvQPV
xKEc8KhtGwBxDQqGPyoHQWB2C646EiKeXMUpH7yOvXKe5K0tW18y+hdDdfE31sG7
0Uc0yUNl3eBSQnAU5vHHyTFHoYm1zRxMUrf2jXuywbEDLdzRaSBKEoeIgMvl1m2C
+ZajbHPzJFApRhz9bQr3VsNcJx3njhEFVI7x4fJ87f8YQeBo8ghGnmBxqyesQYG7
NqjlICGt2LdGXqAFM651/YfCZtsGWuDENjyFBTlKnOKg8U3de4ldF8JhQpZJhLBT
M8l8iWWg652SHEgD6wUpI59rk+gEYXAl8pHORLDETXgtaNHc3+UUXg5XasQzmmbM
vr6JBH3qv8y0UgDwkpxQ552KsgwhSeDW2/sCq6O05wBttlVWLVXYq7fUjaKoLY2q
fSQvxDNnm63UHN3N9qQpo6jZ11I1VxHUcVjc5LyNbkBypExr9cDRi7oTPhDmo3ry
uiQHgrinwmcr2Tm9ClxY7qZw4Zpy7bUS/7h42A0ac87jIZmALjmQFpYXCDEj5kcH
sd1wqhebRZLCShqvj5dx4nQUsHmeStPT80YPhcEwTz7mvBo5WpU7xrtPYJbGFQxf
XQ6XJsl+Kr4ffO8w+pRHxENLRAb/0dUMQC0ibl7WWk4sjdgTSqdkfkSKJkX+1Qf/
uQt/1KdW6q/PVSHQFf/0xUyiS9Mtr5P6r++GM3XcQ0yCxknhOD0PqA9PhCBwQKiO
ZpCXolMgpoAQZ9AQORCLLu9ahG3YhRmlEqPb9V3eptfBi3FFJbwsC2KFvDXfnXz5
Q/UkQ9WoXOwqQ6BLULC/oltGIouGG0lnSrXtG9PpIF0KDZfcDniO81pa9D4NV5XB
nL1+chZNXU8xW/zUGvdSU1qZ48wAeYJkf+VV6rzc1zKKmEZ5PONltWLPXZxMy/w1
Ui+lSIdsZlNhdQdYqZFEMSUQZ4/1vLlPgZnvEnosXIlP6Rvp20do7dl127PJ3GQa
hSWeM4rV/S86nTjaAr8lqUaI+aw+c0qaFAULrEyHghwPL021AOCqvcDcg27LE9Uq
o9mleuNuZzCAzZr2s2kijddXP3C9a//U4fQslxTmvQVrlTMYLjX6mMC2nBDiSIvY
nhBK7uwJj4AAwGtdib9QnaNFkpgswIEnz+zgkgleTb94sB3zK7vh7U3tM/Q1Xy2r
2K6fFTlYk5KtMD0NOvTcu/E/8UbGarD2lrSbHI9Se8JVHUvlpkjtz/NYdjkoZ5mr
mYngpAXBsYzSxbREZiRMstRi3yuMX+QjR/ffrBc6oOuAduhJlBw43vu619QeF70T
1q3sCrnR1kA7ctagXh9xzQXT9iq+xP2nu40ofc/QK5fh7iT/21xijG2RW2GWkHev
s0sHd9qmzZXVhsUMIB4EsPfm8VmhU268epQqv/CjVwo0p1CTmcUYWbAaPNvCZ7HZ
Z+saJ7B7dlthVsaaDJ+x+6H+0b0/kopajJhiHRtdTvUM6eL5qXUlHfcfroYq7Dcq
e+kS8RK3qbGzO1IxdFwfCA2WQujetOnVDFK1b312GMkJjZccSggd+oBiMXZEJw5J
pZJSYDOM/BYkbC4K9VYX17qeO6PQWspnsu34ROxYXnx/FHAnJFtB2O/Pjz5DaMZH
xQuFg4jEJfNix6vFYtX/wueOC2a+vtkewt5mpV1xepmXjz14OPgYklkOtlHTeeOK
byTEhX92PHUMmaLHJL+PG4sh0dRGDW7ro1AuTXu5901VvN2TaHmJ5q7wn00tMB4S
CuZXrgr4IaZvyQoABrNV0q1AumWGc3AVAmEVsQvKiMdmjnHgFXSaSBtCkjK2UAQQ
Y37mQgrrdsv7e8hXfz+UloqVqXnW1zK/Zm4ZnjPKoAEY0GbPoZgQuzBgTLXzdTKV
x4W4bxvQsC1tGOErlZup/IsETxst4BPzvhDiIasOfH7YEMyHTNI1YwwqU2Eqh8w4
BXKcIrH5EdwSIchx/RZx+1QbpV4mYv6hh/bIZqTjDBA3Kz+4P/urkZ9O0yJ1iczG
l0QIdnlLJu5RIkbrxZkhUfZKws8LHLvTz73DpHZ5UgT7/rA8TYUPdbdJBKy216CV
uwp6vMeVe0OJZ2UJtVfssFk+2nCmi5GZwy86unFiJCLUGU5SyYlwC2dLssTxf9gE
gqacbEhY2X/hEuhbo/Gs0wnY4kd0Wdg8u3psxoUs0LSqNipd4IyqMQwey+jZ9WEW
u36c80mwb203Dv9LsoF4SLbVHGGZFTY0Pq93kNMNI9VMJLG4HrWNXMUyhcEgIVdL
kX/HMMoi0oFWqmVFzw9aiatB63dQyvOg1D7vM+mqaN9FurB9HtheFzmAfrsGMjjN
cpou/Yah1VbF7xDQuwP99GuzDbRjU55J6WjA/rIf0dX2RuBN5nMmEOPDGV9jRiVW
UAOtkIfmjlkTgxeJVVhWeFi8RkmNAPGC9KfXvG7+kSbzsM6kfkv7hfKqWmh/0AJ1
Ahy1JMNQKp5/ZCTaDKTx8NZ/4ZqIjGi6+yGr+wfz/RXEkTXa1NcRA/Yz5J9jhGSO
vcgq4Ct8dNVj3Nldq48D0W50UQQxGi7vN+W/4cTLbMezkr6y1zCf82xxVKTUASu5
k7VvrePzyEkaCbGK7h5neMUbOonpE3Fz0pY4nrOP7e5hoJ6xwLQCGFktpGcjzLZx
9Q75km3PoPWGDHSbHZs3eE2YdHI/NA3vvb2nVykVgk9iAqiMzlpTEJndMzfZpBIW
F/puqWD/IOsYhtLUb3BKoj2pvov7/Kxfz+/9xkFDKAoi2acgv+LdkSk35notn89L
RDTwQ9sqWR0cd12tTFjiUr39aP3bRyUSeaP8Ql7AoKTpEa/ADuo4LqU8kZ/XqikP
8+nqaC1lCFq9shhqs4yJxi74qa+CeJ1wrsPrrls7YxIA9khOL1qrMJfqf7Fzpenx
59p7ITKDKq0CC0L/o4ZuHcduRAjU8rv0UUp+w7snwxZXKQsqgpX+He6vQFmXIF+i
uAfjdVLMpSC+GH8K5U0bsmIm9qfJMtfiOnQiaJeEKANcAjcfNeliEuGK+l8fgGkM
KloPGCQOQrCIvbCSknqQdSU/rt2rwFKRqChMZAzaY8Uo1s2AwQpmsSgnaDRGctXX
8k7It2gk43iL8bcteRxTd+k7/wyDjFyl6sfgFGeRlK9Qbx+CLgrSp/3V2AQibniH
Db6XAwbscN6HY50TTPMr46athtH7+Qi+6qrI9CdpJTRg3jJ98m+KMTSFo0MuLeyP
QXPJF6N9g/5n6ke+opQvFduubwP+ha3OHACqEoC1OX6fYrbsYXEnT3xnMUtFGdaB
Vy1QM6+rKjCIICJzmCYf8ahoGkLo2shIp7qnE1Lx+z5TuRYr8mWEGKJTQ8vp+rDp
03ZbTSiJ006qz4+a+ADDGlXbfIu0hBXmo1NhfuhWaljkQpOFZHUSWAWVte9jdbuk
ug+SBwpSzOhM6DLhlEsS3tyHXc8Md+z3AZLwrrWfUlj1kyFIVGjkZMUrYzGKxMku
hAu6MW6V2g7xxDjtNnNCR/S9lKlDxf9yV67DLbzdRErNTee0svcbO8oav3MSyyVb
wgWGPNlutdzvHRebAHNxCkf18kCr55OVDThRI6sho0AuADvn38jRTP2+dFwuNRub
L+xzeph5cp5fKGQA9/I6tVL02KJ00cp8UsbjvyUtrARh9P9fmsfgmAFLPQmphwuS
PbC54SEt2clhELaFRQ/7dfLMYrjF3BzUXkgLiNdGBKQDQcVBCS6NixXGT45WWE6C
tiOHUWHC+NWM5BY+kg4T90zenqdmFsIj4b2n9QDRcVJkMNX127Xq999W6sEH16+8
++pjXqj7YaDZW1BCWQ5+CfPpTiRl5fnTvXAN4rceSocmjAx8rBkQhmQcah1E2MXa
Q/6zi1p2qXP0PV2k10gYVAUrod3o/mmYV8e0AmBqm3jAH2TEp5V1buOrhkxKfIJS
4yxbuQJiGxEg+nYwdPbrRlL3BvfcgZre2ZLvwlzA7s7o0Woc4+ZINkmQOXZU4q22
X+6IRSAV2Bsd7m+ZCK1laYve/kpqKF+bKV/DY2VWCoVYm/5JT2ipLhb2pBOREqAb
+GD8CXNu+SKHb3BkrOVl5qA3GdvQGKvKQeklkjfszVlqqr4B0H2TFKNWJs4ooqw/
lOf9c/wI9Z3BAg6PSxjSg6COeoEGPe5DEEbsAEjLfXqi1f33WQHpXPN8qwMklOFU
/23v+JwHGtoCUa2w0nCXGPQBLanFjRL/WAOkrB+gxi+2c4XWyojO0p8w6Gyybpwe
raOpMvNzkXVnuRlUVtxtDzlpzx7ds5QDlV5E2tyNylMs6o/+5xaXhN3DLmECOHJy
Ws5A/BA0HZPC7YPthBUbgp1QNccqQaEqzeDH+l8fmFimQdPO0Qc4wKRr7trPHfLR
TAutvzEx00xp8YmrcSlFQTPsCYgoJsm3bY11pD1CSpBTHYUEyokKwsvdejOwJPkt
mwDoh0J01iHc+bDIw3uC51cP8kfxmulCwHQTErNkvtMbvnEQbh6zbFJrKz9YFpkD
/KmF/ut0p9K7LfY/x/mJa58urnyVbdrEqPk2FAvWZRKyG0YbIVIj8jJ+oUyCC7pa
KeA61bob+6WJMfAGm+twXBX6eJ2MnTnrlUtSopMwzGZPoRPHRgEPjM+DJh43pFAj
a944YPC1XI+l3LD0rwvI3YhyYbSJbmY5iPS6dEIo2WS4Vu/XxUJ5c/O0C6raefYy
GDhKPDYPCVREH9aVEgofd9wU4tY7vma50VTJnU73gl0ZW9LJgxu1Aj01IecsfYbF
80qZMMSnZvQHTLzQKAO6FtZfLB8GjAaBUIhfgOTQHrixbrS+l50h3tLesdSXi13z
/+J4HXrbDSrG5Hpq6bWbG4j2hnZbShixAjZ5oomlvioiBvWxn34AxnmqPFwCx8KB
C/XBR4Lo+aNxDmMwXjLH7DgDsFez47Yb0C1w0VfuV6ZCffZD0oh3++/ue9aY3DwU
RwfF1gqV/ZJPn4qO8rhp5F7cI1cofXN3fVV12APaoUnGWS6mN4ABlPpTVrXlOAn3
0RSbQyQsl1yn0Yg10PjZYRs9PVs7WiKhcY/kCTBMVo326q84dXjN3e2L8QllTaHc
b1epJw+YrS8KC0QRaMTbPrSqR3XkI0d52rPu3vBS5bIHGt9kfJ+ZEEPPPs+rIwnG
XgPMh4ColjZV18/VW6Y5VYAd5iM7sQbMtvoPrh5+1F/y+khJlz9ddHAeJ8XuePqr
fMu8KGmzzbl8bvCVHeLxOzXFUVgra0xcOLBHKETbH7MtuR00fCznpScATTQz8yia
rtOzQq0n+jrHU2mv4AYfU6tmQcGc/0xPbIzBDKc7NvP27IDO/lUvN88FbCHiN0y2
6V9vjq7AZ3wjrbBEtfYpREvFG3tt0A/YhRnvi8nsNIg9LE98B3cePvjVNfZgWsg2
9iFvQ0u7wBPJDvYszj9T0GNk83ab+V0jYqISD51s8460ob9a3Rhs7rvKmjbRn0i1
6l7GuQCViAg5/LQv9isTe2K9iyHFG+2rGvQIXmS2162u/U/OoxKfPpZ1ggT1bi93
SvmBELdnTREwWAACihHyI0YO1DqiI4hkYsm6MNwA6Rm7vrcm1z9DveL7D3fGQIvl
a4zVekjY9q/Cos4MpeADozo53SZO/70Fjpp+xYabvTa83OsGv0/VQzO4IVY4b6Uf
8o/ciBdgSsvclCjNRlLZVRwF02xEieDDi9HDwowyyNYq9J2/ie8K7diopPqB8jyS
nCeiCiZ6D74Q9wxlEwtq6Due5vG/cLq5zGFzLU4XAXaxjgXgUHfV77Y8RafttH0o
sDTKT/5B6i4D+XgXNiHbvg8tLp1LqVHKrkNMxqL2C0muOK6zhvdjAwpxDIuLtbgO
hgEtorQD8pgGMVGX3ohrgorLvQj6jkkq4Esg2XcPHJ4ZsYXVgfjDxfk9FUZCjNM6
e0RdqIhASrxlROcV/ugCjNyHCAp43u0RkmS9ivtc0wlA9VO9Lq6UBCOsDe7hoMLL
+e4ocY66x7GRlL9S2wZysIko9Is0tp7UmE4Yb14drPaJMHYxH7dA6ScCRZwj6b00
x9n+OZEjHhvgyA4l8t9aBwbPm6YxBHMpAUxfV5Ph9f4h5j8J5rzfFQ2FJ8J7Lpfp
zucQrWjYrdem/A3oPhaRh8Wr11b4OywdlNbSVAv33SFHEj5x+N7c3pcuwvDLa2Eu
oRWUjeqRggIrjWWKr54miXy1sKyhALxzPFd6aJS64IoTFGmFO6nm/ZjCxY6VAkR0
V4pZHleXnVdUEJtKb3gRPww9zj+P3VxqN7s5eY4VYsOWNANAQ5aLbUSllAFwuqAt
8TlGXDqwjnFvV2Hc+k6VtF+gHgmis+sXpDsluc2P9BMtmSgAVRZeN0F+TfiinMe5
1n58YeX/6M22Kz8jJi94xnVt0CR58VnxVcDlRX1cye7Aw+IWlb0/QwgNRLS/V/dv
8yrmQKDwJVvpsxmnzJ8atHwXolEgrT8oRodwQ+F7bQhQEr6LkzLCv0C1+Mtel0kx
hoqNM+xDkHkImFk0K/7S1i5/BIRCV7DwfYcL0qzx44FCbh1QWwCBu6mEQc0c2n23
y1N4PFkKOUZRg1uAXAWus/Trv8foX/Az3QgDwg0wkeulAfEeOJicXR+ONz76WfpK
yLgR/WBNNFdjprhpQYJZxjm+aP7U9KhvEJXbOlT0JCIQimXIu1I7Ql1hT26Ajnyv
9vFNQSUeA7BgMMwQbXNYn9LEslt+o1doR6uLZbXRJo6OVfbjpcoc/NVRjJn8aBPZ
Lri2TcGU8fr4u3su/wWgFZ1CH/HI8WavTF+KtMwUR4gKxB/YbVwYYZtB6/3Dp40X
e7XWXyS/ngu4XDB2y4kGr5eahPEySSLLA53bxVJMCJ1YZB864wJBMV5jJFxSWjy4
AdiFrWAzto5l17n/dBg82n8ZfqEJJF01aOs0G7CiAog2obGITdxuSioCtTDkq7fs
l5HNxkkDeDQ+7tLqC9EPxeNVLx2UdtpwAKFo1MhPvZ7nZOnu/FTEzqWtYnmLA7Ri
sV9uWMfdssWU90b99G/OO1LVvWaH3CdJ0twwWPNMq1jezyCVX5EDK4Ejp8Ztzo85
9XrqJitn9nDmB1lRhJktfZhi7wKyGLpk9Kn9R4bAPeOL4I7+oq724wtwbimZ4NSj
NoqzLkTybl1rHLOx7qOrX/sxPID+hrm6bsdEUOdMieZQkz1Ab/mgrzkaWptlP4/Y
tqXHONfKtp/r9b8aDrEf8SsklEeNw+rqJCYeJBe4xEdNFk9rdOEksPQzTTZggEtu
9JjUWLHHFgcQsS5FD7/3ns5uVzN0dPIF1v+qOVaVPVvcbXUXn4eK6O401XFqkqp6
RzD3k0Wg28CHSLUocwARKaM3JRgijIxZkTsyY8OBQf4v+O772h5VZMcjrL8cvck4
UKb93G4+Pqr4J7ITE3DBNDYV1/scoXmHht+lWH9GxCz3p2lBBksacQk3zf5/1Ar9
zvo7pv7ONAjSvGLJZgl7pBgKECYFabBrhQlBr+1CibSFpxZHg0kUPz39B+GfezyR
3/0rtWfO5Dp8WmHMbWa5OuKhifBhT3IXXTNLd4JIQHs5Qpj+MpEvQxjOwDjb/zT3
YgaBaK29zhAuAOzBeVJrPh9asNwUUWvR9zKVjrurD4If0xH7j0S8vHObqYnnsvDN
w9qfbZCZFW6JjToAZpfv3f/a5P8rwJGGZn0n2I5LE167QLe8j8LZf+NF/RGlsSUe
UhOxs29NhZp4Fl5fok21jdBNiBy7DypP6/t0kFvEaG5xTLf55QBzq94tbjF0PzqE
XAzPBoou7TDjZ+W6upTVWJVuBCs0rV1G+HV5mNeKIJmwKP9rql9PR11RBkkzZMXX
sNkr6AWu2aJKCycQroz4CShZfFbMOErVheKyGxOxqAEzZZEVpH2Qasq8Ii5Gcuu+
uZhSV10NkMPYVpY9XO0Bu9HxHn/GeaN+XIu00H346TbBI+NMiVvqdAu8FFXFXLMH
pL19Fl3gny7w6nhPRIPQP/+i3SgZDj4GJEoc0uVUAMnMByN3r1HNKMb8hHHZV/3s
eAHKusXtTdZKUMj4kj3y/zl+TmV1wbZZ/5G2OYKBz9tHmC2eAhavQMLkKVtTbg1c
xMxcI+zHvgLrg0S7CleWJSn/Lo1p+pg2lt47BxjJ0HbXsawBA4rAV1h6Pk4qBw53
Qtqczd5s/Oek7T3oGS4lG+ogUrChieaXpc0DESwIIvULv078zz8nfheKNOW4S0X+
UhMu0LwCibRbEJyZX5GZkkY2QxZ9PTLGQTnrRDcq1nBIQyjtbRW0cBNAAxXZdHxl
XBzaKU7aRgkaQ3Qqp4uG7XoGtIYdd09Wd7VdzONrBecoxRGvzkMsThUh2CG2RQF9
iFX0uUUJSbeoZmzJ3PrEuZT0FCdaDsJIWzmcLZut3wt9ETZ/MUsd+RbsjQq8MK2r
eyKN1bZt5rZvoRkVySuOG6RlcOsWEuNH0RGjs7bNwpwt85ESpMjBTpqn0sHyWDZG
MNOogeDRvtvSXQgGrl/g2DkMgBo+Oi7SGl5f/PUGAyWYaT0GL8278sFkWWoo7H9T
BLGy9jh20uhWv6B4UO4GlIPU4zrDqqWMRK7Af4YiHHTjrCUrqBZvgRptc7wmgzjB
+5VaSIWGCsdOkvCbwIfUaaIdCrs86J6+ukO3X6xjKBTY6IAc7BZ+A8ZhsCpZhwn6
11VBsdiu7pJkHRVaa2ew9cyM5NAwe28fMiUngHOgieMJXvUt+8ruvrwt159BY/sv
Mvppw5vO1ZAs9s6pdVZ9JAM5AmFobUj/rDAY1brJKD6VKnZWSIjwaRTF7I/SlDrU
J2gDSIID3Yzqj739SRiDpqSLPlq8Le9U77NJXHf2Dbjg1F+CrAhEGIUZGk337MXH
anCT2CBwxUX7IKiXl0ucvMvbYqZNy49x85rkbXb5q4u1jic0HA9NQArvSkqlTDPX
mCZfoCopbHIYUd3bXWGJzrupqpktJnboCL7Ly51iwQVeh4UMICArwnWqNQ60vj8o
qyVViGxUJT6wBQpt6OJQC9G1hOttTC495BgbxzugW8W6bXeZPCpQiDayhcvOhy8F
oiGOq86ivCj+H8/n3MQq7I8bbO0ZucJVZmA+e3Q/xlrQd8uHfb4W5YipyYjDrH6H
+EM0H90Yk5s6LZ3QvHobwF6Xt0Z8rQ7bRoqyk63HR7uJ5ohjLFVOPFQcK+9CIdy0
xngtEZLDUUmQkm7tFQIitXwLuT7L1vmdKaR0dYjSuhUsw0cIghpT188cWPTP2Lt1
f5QksKiZJX7FDgRk884BZPmLhjiyeLg0zwhLJAVlQhsE1EApoPBs9kmrcdUPxLWF
/ZCh/IAewSYMRdGklRHiQBwDA7Sj9/P9BjslAGaKAoMVdTXUtwImuUOMYamw9Bqj
3hAY+9NwXPJtvp66RLdqURgkl52EQ6pwi/UwED4zvHdFYqK8OkgLBcVyXTETgwpp
dMb11ZCUrkoyjKsYw9OOaLVWZ5a1XTA665Cga3pr2shm8i9yMjwlwHjm4dHf8+OF
+d2RXWyCU0i6IP9l0QhT0Uu2OlljwvoTdnFtnMamV2hbVi57vVD5HFRwCVwC4VDA
0ao5c78vausj+yKvp/BTpxIAFR8gdCznHOkdxeoZ+tUNHNDh6bUNHrMV41ps6NRt
81R3Zb7HObME8aF5FDkf0U4/jGi6TjWJmM4P7BoSJ3rFZQSGLD0zKBdCWfcAVatq
2NTKq3FyyEVt4O1ECn39z6oIuq2t2SuuivnsF/NhB6jHInUpR+lV24w2ElX34EKK
8IQifo1FGfSqjSBPXacnietpu4Sbxc6ApK8vtcEJZ0WV6hYGnwLsAxNAKmjnsQJV
OLmGh+zp7+iPaFubuWedih1Jk5pNwDwqI1SoZS7EvY9u841A6ghyBATbVB9Rx4yO
2lFZpxz8OEthWBUlUIZLGviVtR1nbh3vOf6ZUl9zWxMzGZuHjSHHcX92qdhMoNuH
Z5a8egXlMQ9UDs8R//PC6Uv2Pyij2DfIrtlHFT6nFgmN3f8EPah6znFn5g2rGnmM
vDcuI5rgVDkX/Wo/jG6WAmZNWh+uWTX66efH3kR3cpMqLQ5Vw16ZPxZrP1GByVvg
VkulZV0NxNoukbR4tQj2rJVXqAoX8MZC8+gcJd2qMlBof5uWus3B9GExpMQPjA2e
DpKukXzVT1HzPS6kPHdcqFw43iFtuSZO1LFbzvLRC/l+fn42UHNpAsEAI8A+iEy8
DIQYLS69RrTEp+W5k6CaSc+KJITuJcRQi7XKXHdpGmevdr7LYnam4/62FPudob0Q
LvzM8Xn57GOrGA6Zp/tXV1cdliFSFMH+4cry+4artBhAZnfd7GdDwaelcwn+OT+/
rXscQLZG8XcSlajaocb8gi4p+ZNIoR0p6pKn3pVQ7PGYi0/jtAEtA1FnQTgBu4xz
U/7DWY1GWptS0cRfRZOsvr6wIOdLyvAc2GkzcRN76gqm43Dm//mCW+iyOGCsVsTD
/D+JqD3bWX6Y1Y0y8skjEw3zSTS8CwWszIDRZQT4omse4xvmJf3HtNyhjzPgIXiV
sAniBw3Ti4kWljvtd3cF6ii+ljdQEH9QWMMxz8cRq1gf/vQ4XAEkZkWvQYN57d4A
yE9aK6WulKDCvfx9Y/VjuUANdyuhkWr0Lav07zycpsGd61d6AmYO9OH+FOB7mtu7
cUABBJhEaZTi39pLdnNYCz9Op5pqIEWQ46SOwJk0NJdHBsHu5acx2dS4A0CiqlJd
uJxKJM011WefHMdAGMg57MGsCByjbRcrrb/qDELwRCODX3rDvhWXqOh1Q7iuxjqO
mZkm/3vnqVz4u9YMG1XdIoCUIIEYqYN0S+KSIAr5aGQKAJpF8t2lEu70J2gp9Odz
PpqK91jDonmJywRhYgG3ndq1Oo5zOP291ldOA+nmd3XM2+3RgojnTSsRzlbNhCok
VFykxFubXdYvSbVY7aMJt0lVY8j11TT0JYlBaF4lwcBu0gjZXcLN/lMj60kgOONm
phWTcUfU+ptjBgZ8qhvlvZeqjg/Mrza9mLrfVOGORZI5foYvl4UEuBFbj4lGwrhw
EWzYX1WLlp1V44iZEZ41KxyDsPV9SAdTbv610BIw2ve/9wfzAHTdrAmiviV2rIDr
Bbrgl8JCtz03Dt8zUF7EfhJAEXMmLS+paZsezDu7ugDidHUH3Q5vhPXFq7lTOKqP
sNT4dwJTbM8iVsuUuuGhKnG/KBIZMQ2GouV3ynGH1XrmeRjQQCt5/b+OkrCUT+FS
2w2QsrqQlrW17zkRlrQNaorSrNx45cBPa+UD59g1T6lGBZXyiQhggPBu30lajG9X
kSo945FQYXmGmOGJrpu8k+AxwdLkExkbE3shfe578WmOPYUhvXobkFL5tNuaokid
qTPu1K17nDGGNXirW1W1gYLkCIh4v9L3gUewicuL82gvfup87Cv3ux6z6/RTnwV0
a4jD551TqFI5w4SosnmRxgdmbA0otBAskoWoS1vDkz9LTnyZDjZGzdlj6hi70WzF
UDz9Wa1FXTonNlncuVvbNnv9JbMMs+NDGFoviNV1Y+mNCqAApQb2aAky+oHOwkWi
shYAcF099qTn3QVvtispMLwG1NFoGDoQwXTusXji/3elzS/g4zkcSUjjyB4jI+nF
Qxccr6tBtLS/zK816xBty7E6RjWdMKdyGw0ii/rIdLhMjq9pUfSzkQAX4/yr5CNp
Zk/WhonrAQiQ5QY51q1pte39Ip4xuf5kgoLMEbl7VvhkuZ5ar5T8cIQPeDIb/wnG
8751K2zj58p1DOesPcxc7JTbgi64A5Hi36ywMH9B7b11Kwcfbh5YoHEwAMLC7nSi
iIZDbWW+QuEK/221i6sBLHZSi0l9QD63APagnt2TTuMD/+CoT149C1CBb3y8TyFO
vNZKDt6s3hSUdau7Y/zl8u6aSMAOcMg/EAFlwmIu/PLAAvBohl7Ph79K9PYxJFE1
FuhID/n0YF0wUVnQududQ241SoMtYz2mMuVnD5J+FRhG+q0zpKj7E/5uHj6xCpmC
arup+ppitT6J/IBpXFPmnw4bGK8CrbKpTglCpQE80LMUTn38xbP/Moj3CqcNzXae
1/CV1F2NbqM1mNVihk9Rj6oN8Iw+n/hBZh+gq1Yknce4JpRmjgx8btHQNIgx8i6V
cex7FlekHfIeUjLML4xKvcpgEOhqgQQ6cxsrHiCKv+kKcCmJBoBCQHj1og8g98zq
S2tZFB3wkVsuuTX2hSVUvTWw++iRUYxxMp341C8bYymBbBPvT34mqbtNHSgjWGVa
Wp0LPFU0N8mPCMERWzd3ChHeFRTVCLGZx+tTWHJhCA9+H4FsHUdEkJKYresCpwP7
VFBBPEuMFut8XzJNs6JvHWwgkYvmyfSNtjCUhhdK5uHJVqwB1nlUFUTiFaPzpqgc
AE/SqrSNteGnA6WidpXGYTXdWXKA/+u7mJasCkYadQHQjbhcFTzHr84yxPpWEaGZ
FrQ3JN/HD4ibVPtth7mLgPpIsT3ONJNK+qGtNFvVc+16YfpmQSZslJ+PWSIp/+nU
UjuzJJdS0BHjLS6eNRD6kjxK2C94cuIMLkeI6TVh349zsxsBLgXQ9Pm18LrN4Yxv
IF+Xo0KqL/EkG6/IlsIaCyKmsU2q867i+BsJJcPKsnvJMszl7428qHd5rihoyy73
9YRX/w+yB4KIRjywP+scxrBTZ/0N2IQTa1bCTKHlvENo7UesfIEUnwx3fCB6TLxD
rKWStG0A36KuarMnjJe+dnIdqhkH3QD/gRk5TReszAKObm8py8GvJP0Ar+fqvqIC
wla4USoesayUCtxN3G09OD0yUc2d3EIdWGRsFhg0wDG5FU+tn13y7YaeD3Mm8N4i
9yyQXctJwQi1xAsuBaJHFzKNGt/utjZTpm3c5pLcBXfFuMt1qq0+jgrnytHYHtoP
ZKpopA090KNo1yXw1UBa1cjlcv4FBMJhclLeTR9YP9PCJ0G32BWnIY7GguJcPR5T
YpL9YqoKGArq++D5VoLf4MJth+usKB8cORk2pDR+u4R0WTLKYr2rkUfcn+k/WNnu
mZYZBb0vzfPL6TYhTWdSNSnbFbg0yGbI53SUG3czXUlGnpC+TTvTXDL6F1c5VyFa
1OdZmhJtKlt8J7DOiyP21tizhOI49drvfGMx/Ioy43vv1rfBPY+cyjDJMEv4xyYQ
8Ou8e2vmJSTOEPlWNmIk/XLwjyBU7BgKeVxPPD4+la7GsFXW9DN2j7bV1wSMzcGV
zBULeXrvug8o77dMy5EiaXXQeATRxB/mxwL0RUIYtmcR2gsRV7Z0TsXQcUYfyU1l
lUCgVkHXmsa9Tp3WcobpRZmJJkhFNtM3DGF6e7sTybbli6bZIM2/J8tK3ElgQjUQ
m1WIHqKYVtuoF7IRCgZp2uWag1Xu+9juSPBre2H/KL5J5GenpJFxJV3wMzcy6Hx0
KVp8inTIr+iZoymx9rAJgVMY1RQyW9Mi0L4OI0Bg3vluTXGgW7gbbQXu6w82L/QU
a90numg7eZlnvwFp/L3q2/oKKf7PLWKWMrJKOrp6N1Xyl25W3CTBD2VqlW7vyAPu
zDsmvvBH1NTYcMKG7selx+ADQX/oHq3Zu7pnu5tzumIYEkkM8kI0BFSLfDtM63q6
vsVcQKa2HCh4uAKwvJc6X0DbJ+evEg2dGNgo/segMCtO0dd65NjXqkRl1crOAgw/
uRzyIG7bo3GhdOuhgK/qivjd1HmZ3qExn+ISZDdSq/eLQbaU7kLeY+x4wmTnJrlV
pLC/or6M4eEmHpIZsgegn/iHWIqoSQ34Ojl4pUKvayZvMVFc3R22NZbrS/HolSOR
cFnTbFrCY0Q2/Wa7InPUy4ykZ6jnXAGlhlPYiOR/NYGXXhX6LgKhFuxC3AHrBhW+
RqE//78kl0QRYI62p0dT/Fcj7+W00P+K0YHJektUIQlaY0KTw7qZawkdKgiATqXy
qVd/FlWCNUmGoH5u1aqX3B4RqTo2t4Y0fqnIildyiG7YMiaxybT0v6DQitpsZgAX
D9UbUH/7DRSF/GVR7u0lqjoJHIo+Rx23mQg486GV4Ry90myAegwmJtmCfO+gmc8P
KuFfNtrrEBF6gJ8zNoJlDO/4hhP7oJLdMnyEUqeKmMyqMtiY/8USS3AfCmPJC7IP
wtvtXIkXP76rtgN03FS5RpbBwFI3FixWg3pRL85eVmDnrhNN8xQxGTi70tfrH4d1
24mNECTYHpdt8CzlM9Bftgxnfb/SrKHw2NIDBXrH2ytvPBKpSgVvxY151UMOdjp5
TetNO1HJOqGX+BbPJfkQMFOUau8cZWAyQoNsCGQ+nsYz1ybnUqPOMJKTRy/kkg0y
RXAUPHEGmPUCGPIQu2oz2E7YKfF/oIGQtgOMo3O/XGswJar0bUqcJs3BDRo/PFEi
qygxzZNC80SfB/f9MRgUBi26oZ7pLLdJNILPRvkkUd9FjWPqqBGVns6HCeMNodAQ
SaLz1jXjp+0KiT+nALYRRaZiTdcTVOyHmRSmQMbTlruMFKZCMB/vSYamfE9gcynA
4njhqsaWu7SD1hEpXouFf9fV62wcJMmoKWgJF7DQNumfMxN0RL3QPk0Krn2f6Nan
TQQKdoYhTrDZ0SpH5qgPOqCIiCPFpNiwSu7BkBqtsqlAX0/C3fVZ3DYj/YWaYZTV
wMnqwjoJT+djkyeYzAKd83Mz37gLBq4TgWWN7h5R4h0KsCccCRLFWyLDbWWZWPvc
pfuUPVcdEHkxo64VnLOVwalP1W2xxXBSC3SodYAY7RPL3fYbbNb6j0Pky7O53pTh
buLvMefg0+oDOiUBlewjtN2OE71rQu7wLIcbUujlEhrHr8EZBHjR+/s/g/r9E++O
av0Y7x9qY3YrgyBqsONBqbWL/s88ZvNnSEhjfwIrQjCJdMaU67CXL3xEP8m7znzZ
NAPGBNMJ5QXMhDh4uJ5jd/XIgyTf4epErq+gGiU7sN3HR5kCSFUw1vYL1pQxp4+E
k0eBsCjy/y04I9dYg1q8GYW6rLrVZ2vYRZFEYz4yDxEK5uczMqzR7RiC8m62HH5L
o9vLv6STed6kY24/cUeKvYU+XNetMZyR4cvrSqxD+2obAVuAlnmspq4X8Bw0jIQV
bUV8bblQ8cjthYTHxxAe5wucEMl62hyzGWb++aIC0nQ6SotCaezOi7sEzPLz23D8
2wteKywEMozMD0rwDhmU5rMg2vuvOZtWb9eC2s3hO++FW9TWisr7rAvFT2ycURET
6PJB7iPG0x3HCnBE3zbQI/+9G3oNAk3aL2dBD1q99LByx3VxYJUD+P3hRFIGmVFb
tbxwg4QT/YMozylU8g4hB0aStUvc70odKJ60jfTai8YB4nbtACDtjDZDhdaNHOgn
Iq3P0O8QMEcFVcQLdb3QAKk/r3EaVEgRscEbJIr97mpJsLTtpxwbS+gWbPAkQ5SD
GMGfNX1cyYJsb13RDjwxqi60eqBbtcBk4d87vAd4Xid9+58tmYCXgTrAOH0nnVXr
UdlUieyJgvofHj9MYx8HKpYt4FWjJ7qn7NGHYRPsCnp+671r78yYcH2JREC4mOtn
AWs6DPCXsHMoAcGgVtJNZDMcs3/w5mp9siqeE1qx4cJCz/CqiRPOz0/61jCo3I/P
vVJITxOFffnkRSM4l6T3/6mDvt72cRjvG1qxFuscl8XreY3YSIYcuaBneMhimgOV
+cY9A0f//XdjUZh8uKdzEP6gLV2OjeQcYuOReh3EBcQK8gd5nqWgqjIukP8brJBl
EwXzeLjDdv6WAWdpSJbBZ4RuKzsN/cpZ0CIqyrbcO7QOjs0iVSgLjSB5mIc8t4dg
mWRbPucOVVSouybgIZI4tMgJzys7Ua/xlIAv85jYBO/QnVX8nfeT/58JbNqPRA8Q
BA9bNCse0Ydt2mrLprpmjKAOyGzvgW9/aNI5ieiAZsJyfzZZgMAUIgvnECFQk4Pc
OACOYui94bqQwFYeToDHo4L3+lrXsy//N5lFyfLzeYRxBnZQua8TOU2fWV+dyZcs
VY8DKlFJR/62u0grEIngHkA8X27NQUnrNsOdsvlaqYPSlePqHZCbPVIwYkcFT/4T
viDKst3u++wY14MfZsHczJXoFCNzAlcmZSEjpbyVufczJiZmVvcGrtkg4XQIxLOm
Ha18+IhtwSEi8KagN4fZX1D8vVPQdh00UHSpKwZXW9Ka9rWkLmyjM2RgHq+f0jd5
jtrRhQu30iJjpGVQHjlMWm9ucS12/aYXz9ay0lcbhG1Tbo83bmXUFhFeRrBOdJPa
TMMNKKtkGCuEs5UtESxBA5PERfbOlgfKozpbteX0oGiFydKInr9Le5eZKj0qb2eJ
l8EfDqZSNu/rEHy4OljKFhGk7KDJYfVI673C5t9wA+u1l2f+hVweeWwlY0BENKZ/
q1eLfEf+zL6pdoSkwxC/JxOBGOGwe2mKZ41QD/beMQu/ArG31Nwi5oCtdbgQe2dv
pHaJAY7aiq5xM/q02KStY9EILFWdC9sduufIWTJl2FAVMQENEeaPmzJqmSN0xHOQ
01U4FpSwY2ZSjA3GAMVThZvUjLE2obti+uCkzsISaRILHZY2KKdEIM7BIOmBnEXy
BjkH4tc7CIxz+iJY8zurY42dMs88Iel0ZX/iNtxZlA/63Gd6jXgdNKmp+7L074Yp
MhC+UTP3jDNAHi2srv/3A/swNB/SlfgZu4jJIJCSj3rnZQaO5EY/IHlTc3iL57BO
dWzQj+BcPLqEhI1RpS/hwmBZO+a3KtFyTjLEU6KbHD2/7v3ydvnSHVuR6Q/qw2dy
ngFrZ/G18eHYGn2+zHNWbmzAR8s1MLJJAhXyazhdcJmEMv6S4V1BAPjR46lo6kp4
zRqPlFHcQ4WDpZXEDxYrizecQAxWuIjTYM6EyWA0XOFsXs0I0K4yYMshCz44lrFR
v6MW5JTzfXJ58FIY6pAvK3ClpnrX7jMMrii4QLyByyhRlUMm2O0Zkj3U6eIR+rEI
Puh2vNmSlg6biDNM48PX78wzxaWq9630u1m3/Uryai/ViHRp8RNlewraNzjP6Vn8
aDtbQ4/a2YU3lYBFunkMoVoDItMGqb0q9ocEFWCMLT1Zdlu7uMfISWLFQUhN7QuH
ywR9NNH2GR/91qG2K6xL0vXLKv7ap23D+uDz3kW5LHkPdgExLmBUpzDqnRSTyzGN
Lyk0KYJluVd4Dg/ml++C5Qe/JdlfhY/2rOuckVZctbdREOgOD2VLGtYCD1726jaW
OstOd743xLnxXtuB6gqG+cQpSZjzMI579iXBzdOPWpbXmWCKmFVakmpEov7tZsfD
BMDl/Pd0GBYKsOSjdOWH6JRjeTlNO92oWPMGBWUr9HSVamtJlpsQctmiA9dsl66g
X4pJSMpYMfGgc6Uyz5GZydGBsYOBlEg3tlo7tyDiBdb80CJMCTU7/bBo7GmEWT/H
GFLxlMD1W0nao3FN3WSy1ToyLD+Co/pLZHzJFWFX/NNwg0iUxLsJXLZogEQLt+RT
3VXbtaOGgw1+dtrOr0X20JU26upbo6scOrj7Hnw7ufCKb2Ro3/UzOHb6IY/n+tsP
N53jzsVfaIjukFJZ5ZsU/tKduNftfW8ui8/4WwxloVLm1tXmKFSpGkPnJRL1m6UX
KQ103pm4/WfguKIHTpvsk6Xt6BAFOLY3MQ9evwTUHqSHWr4VNRMicRItzbxdXJK2
kJkTWTx4riFnXP4BvSW7cnq9/hchJ0c+fuOX7t5AqbA4B4ERV3Jv+55SPhhFZkhk
rPEYJlA6+OYbH+Xwfdpf4i0N7w29bkHMBfef1mu4ltyHdh76Vp5nGOG03xGfFK22
Mr/8FULe8k55+rrT+d0+vaB4XVM6OKM4COMKf0B1g793sxFSixpNjvBwGH42WICn
Fd27UyU371BWdSnKPd1tQbvixltCMuxqCga0uYoQ9LFfMvPTep682D7N/LslFzfn
SHqLdnBoFyUXHPvMWhOrt/8jdWDCbh/uT+oumBJMUKeI0xDi5RUsxshgeFbU55QB
hKBdQfblqHjAxk7idhoKFT8RvUkmi6acN0sUowFzbnIwl2Di7koCM6lDACHT1gOS
qgRcxPtKQbqUPtTlNz0momCLZ4IScLfDbEQskMCLr5gkIn6Ijjj6vdtPGXYFilkA
765fJCbyeBdO909MLlVyKkK+7ClXQ5yVDsZPwiySsPorlStPzSts/bqiT8r/FEjO
47gSAc5tLmOWe15QZ+Jh8VgFe8dyVYOcNiUs7ZH9+cRbvRb57Lij8rRL6eCSRxT2
288O8ax5jh3TN/JjCByCpqW20giY4LZ55M74fGlDKZ81tKM6F/AYJCfolXu2hcHa
0ZM0xTgdc/vCefG2CJfeIIwEUXs2E1YPSiM0zOF+AM8Bv+WsvEArRCmEeA3o1Y9b
VMzgp9q5nhiwgLZXak1y5Nva0Ix/Z58GtlsY0upgZXUvHQc8Ihotw385vxG9Irdo
xVqTDElzzW5kM1PL2rp5GNGdbY5UDg46z6xagiUYwo9zzi0J4tzdnSYeXHRU+xVY
n1hM3S9OEbCmBhNIScDZJKFI9tMkOgyiPUzhhOV30UgYxz5Ga3j4SaQseKf99iKg
LtT7bT+pZId5Klm8h5DQrjVCEhNzmxgedZGegaXg8YHkZpmYlbSfJXpFXLC60Wz3
PvKTqO5vFsnuiJJpikBHebOx9e9CSCg8ju8HZuei5VmMvneeAEKx5sp80w5KsohX
LO8K9XMiQKLSfcpM3z3yTxo/SnVpSaAb/9xTt1hnMnbyNEuIfFki1ePwM489/pm5
uRhvQRW6Ip1axoAuot2FEMZTRZI4cEqdN1gPHH2YCMqDkeo2FnkCann7Ee7bSOX5
BFxWxcQhnoN6MvfVBTXuofoMR7dtf1Spr2JEFhV1H7ZJ9xTzJmVhEp1+9XXZxJN/
GqnGifwdmFGC+KPLdjNJu7mpwx8L0iKXqEBbgsqq2/zZNKW6fkRreB+xXbg2lmzb
uy84RgVtQpK2n1xJ34Y00koUMrYvUCXKdCL9paAG+ghfkii/aaUyhBgLf/paAvHs
MBwNo172hbxwx6bMmQMPDj4Hc8wAx/OA0WZOy5LnmXdiKeutbWY/wNaLG2fkxBbF
1Q2fo8S3DAlpPWRqjYTyHLxHVM+32o1sI+Xo4OSqxqeBQOqbupDR8lg1yOgK5Mzf
D81C0j8rRR5QMb+Q5oya8QLRdsKzxeqIb1d3NPRWDLrmQAbE0OKAYaY7Uez0ospS
5wkQWvEz3m69TwMV7bHUPk7xb+5tQMVZMzGAVQJhsXtyxru/BhuiF7Y25hVHVUV8
5UiU0H3R6Tia6p5yyv9hvskCpJAz8aEO1Hac02SjsggpsSZjQBQXoJ69EmPRvPQB
0df4hMMrp+tSLbMZCSGFJ2sQieiBCVL9f2SoFbMzCcY/byZhBkcPzMZy9r8BE4oB
T1iCHatLF58LFiEyaJwU/q+oR+32o+n0NRbaHiP2qY4t1HYYgl0W/ceHq75ou02C
Sp7NPeupA5OVUjqWe0WgICYRFGWfZc8l9f41ogHL2gHNAISGZ1fwcffJost+tCj+
KytgwuUyWBEd2GBg1i/0LtL4E/o+N/1IDj4oX6iV8do+8gF9cZKqvvwiCmc4esm4
lfAcPLitz8IqHX57y3uvdQF3Dh/Yx+6VRsI3T6w/gsnLe+JERCG9TumWzPHbHIu8
6eSFF/LeQANxmXqfWzZ236v6YvUiIlXArUQzDPxBeDEb3/onkYzijXhHgyTW3GNL
xla5NGob0EB71NP97YCcgdOg9VEseAPBdx8WLzD6kBMvIlNKqJ8mZ25kyjGfAKNn
tvA437w8e7Xysa3AgNSYJIA3P3a4mR7CxsvANs4Ikrc3ht6XgOHfOMevVTB5SdpO
Xw5O1TszH9dQy1jDM/CTIY7Qu1ob/2gZeGaQq6WeFXj+y5e0ExoYAsllxb8hcHHg
SbJ2xI0LL0G6c1Jo67XRKNX6TW+h6+/szxTdSwjsMB1Cj+3b/BNMJoeogBVhoPrY
INSHaqHLVDofb2VD1l1eXBD4Wrd7WHF4qsj0b0IyLpjdQ9AjHMiWHcVc397dVwW1
saBQ0hDNim6ZE15WYhOZQ5LYn5UqoBQQ0X5m/mJP35FK+xxmYx9L/9jDy/QpMycH
gMUg8hMeKKAOi8SOgA+wjuYDyhj5pJACyeBxni/CYlRjWgeSm/wggkxNYLVpPswu
WGoYzkwStJlVlXGmexUIJBvwE1O5DahSj5B6B5ibk3k5/TVDfjCmUQ5Il6E9Heo7
rqD/87GT0KyOtkYpcx1wFRXnkdHQ1yEFe564BApPQI090/Jbb+iYQ37BCVV9GBPF
wToiWX43GzscI07RdD03rccdjYF+BxowOhZTmIccEatJSoq1bt1B9W1LAsSC9Zwx
fmq3AJusM3VoXSbI+5bfNNk0QJxkujYAao7mcJPm/837uLfMbH+n56EHy7JqzPZr
lVb+jugJw2/aJt+YBsyS8VqUHjOehP9Texn37pDWGySIYd3S4cnceaPQk5qTRHSd
SrQ9Wu4YopsBSATho4oulFSsgng+67viuB4d/XMePYcwfiN19/x4zYHYUuEJDW/v
QkrYbCAWKzF4eYzItikGHIpKu8YOPj7n1/gLdWDyFZBdWpGuyNXe+V63U5ea+OPe
YmPL7XLVHfYC8LU/V6Rp2qQzhcFxg3brRVTWSSzs0O0neM7SOwIcb7ctJezJd3bR
8XdjVena3EdmurtQP7MZbmv2GVj9pdX59mG7M5XCXJpf8Lg4jGzHN0BIqi0XKBeF
o3r2OjnHfcTl3quZ2pRSYOTrd4WiX97B/9M7tqk83t3uCUGId4FnE0ovoevqqH/a
rk2O3K1wpb2KKdY3ls7JMMue8laFq+tXOaoa5LgGiIRwwzK4HIOU8NG3si9y5wcQ
/UIoXFvpHOfDNB0Cv6badFR2uf/IJFlztSZvLcHbMv662B+fTC796UDZZCKGf7sw
7ua2dLJ08RK04XLnp8UbDSehyZu9i6PAF09O3+3mOsAQ6YM8AhhPSu8rCTBG+Ne5
oZYe1GXcKto6Ca79pv+59N/qNgv4lnExQbJtrruyjEtKqe5MHeCMIdFzUbZmatTD
MeODZnVD6cRf3TnCcRlwDL5QJCQ0tp7GNQSAvECfqe1VALS3YMvVdpR5DjunrqW4
jjH2VMXh8igy5niWPFYMk7nYMdedokA+Z4BlT0MlrPxijpGX8iMFeGWU1ySL56gY
uVaQDW+328qGNxhL49mb5hXv3xwrCPRut61gi5HpXCTOZIdTILAtCBdggGkJooYz
8FfkuUsaXQMxSSkJOtdbARj5W/WNa7YXs1jRQW3imOEoLNvpBQBzfQ5ubmVSsY8h
fbZQNYELOwpnYJAbE0/Z6cbqiNOxJ96ruu80EeaEaojxQWn1/jHOwzDAvOonDbPs
wn2+bibNf7OrQDjJV7OTHx6QZTCxLBevjbqmpILw/AFGtq88DUa+fMC4A8xe4nGb
lOgVx5Qa2neaB203KOKrRwCC2hI9sRpeZ4oHMJ4sK1PmO/yuPyJ35ruQD5Oy9QTt
RRrNyaRlAG5G882i4OXaBLJbzpS93k44pTdsdP8K2bql3vjz3N9J3JyAHTU3KN0V
FMVU8itYOPCH/Ec+FuPT/xejJ8wqSIpyjj7nN9YnGswIIxK6v3UBnBpl6ik1yxmQ
kZj7RI81wW/2ryk3+tdOr9U9KxTlBS8qSvl5Ld5XEVB+mZ4y3koZJVsAxSgOgqYo
02uYRebLRNblUwMhxlpRN7gS7SudMrgbFID33MgcOaYW75yWIAYaY/xFNin/QrpB
/NzPyMN6t3px0Mv1nRPodUW0bQ01SfUGyfTzmHAigweeBv483oSKwHr0gm4VffNN
OvbC9qBVUz1ieZtxsDtq00KxoHdttGCNr/r+g/gg63daQd02cmdx3vLqsO5rBvBv
iJKqOnusrBaqcIsqmFmBTmpxi6ox2PhUS6BMu7RSYBgoUcLfZnloR6CYS74TE7GO
CP3zk4QMPc0gKrFCrvKSu+7U5+4uUEQ9zIKnGJV1TM9CMKl2e2lUXy3uRVQ5+itu
AeOItUlydQo79McQJs2ASL/XY0UrZ6wBnJT0LvGV0VcCpdlia7dzzNq1qAcazeIg
lU9D3LeVWdCslZet5kGOCkaCPZd2wcIw+BQVBhfyUNfBXjZE2kmJRMfmv+If5+cl
XeFWxO3tdrzLJBSBnxc6KnUWqtoKf3hOFv+emQ/9oxqthqTZUO+azcEHLDUiWOzm
trnjO7sk0cpJUDug0KFTa0uGHMFA0a/oGmbCh3jqiOUrzMD/UphA12ukuyMEzJsZ
E6TdymrnoL9i8FNmq45oWITCjNz2uz4paL2k65OjlIXpnSkP39mZO2zoneucAAtC
nwfhFjmSVMes6oXCxPLJBkx2L6TyGau6quNVXZL3sHiJMAGH9giT5gT17xf9jyTg
d7IadcTKLGIYsK4KeSu5TG1qNwNxr5SpTvkxonw5QFX7vaSkHDbLETBMiBqetnSO
4bCku0RrdJEp9iGZp5d5scgmfUsEsFLSnrI+HpxYmc5i2kmXOXMtFyyWyV5CavQM
ExvVjyOtBJkz/VZp+Px0pUd/xrNwAZ1J+sEXfsHVrhYqrdyWzstWFvoP5BRHSKVk
IToEOeMXRmdakMHLXu3URvlQVX3pvaSIPrcdMhSfI3AJl53KTUL4ozPi7ruhsBvh
vSwFjqu7MQBPNKpiUZpVzyxxQLcq5qXi8a951gVmLJd/O0LIFip2imGgGyP/2a7B
WeWgj1/hAH65TzKsOwztpbXIguZ+kX3+7FNSyqd4EPx1rW1sleNKg2EjslJZ/+Lv
oRc78G6ioa22/SPSNgKcOMoAp0igK3XGx3TsO5FwpqpCTVemJblw3mHyf8+v6O2H
URSjGAdPMA3ylNlvxDTa2LydQ5ulh8WLJE3P+inn1TJl9FCCzm84eM758h12KKg+
d2hYutprRVBHy4qe8+VyVu6qk1bSqqf5wq0cOFwxlwsR2YHpq8BxPRA5e0aFv1ge
ccOD9Ll+H+ZN6lmetCh9GoznTb8zpkllOQPDujSFBkpR74eXFmIGYHDe5ZHrSY7z
zco5e1szy0ApErBc0G5Z2zbG6Osln6MVIbGPp0/tlcmtxgrpfe9L6ss/ZsWSTbaC
lIoTocuPqYEBwMAUQPGDobFd5iB2v2xoIiXD1x2kEndIbyERzAV5mx1qxn2Km75D
Qtg0ZOsy+Ikw1OkwHG/M0TH+wfd7pfORR4pJVek0E6QCuI2/xFe173lnCjxqPKIS
lAeooB4Rh6W7u232oKnM6Yo20k1zcZz6Uuj3KnlbPMdzDHnBAmo1gu3EXNVB5qNd
U3PiOvL2R4HFKqSX4XWE6FldSzsaHRg72R7tpqhLip3VkLGGGj/974/58uObi5UH
rZYtWl/P4v2prx7BK2M2rb79BRRmJ8fdHC1dQ/5yJhU1dhq/eEfpgk0LHsQVIPWI
MozJOLTH1uoZv5NVfEJ87TNjc21KJ1esSutdJUeN6btzxkH83kBYw2ata9nBnCsC
LIPLrBobDJ4sbWGogvMwcFRD3SBe6GMJ44iAtpdzqiE8gJwVTSNPYpf1M2A6P3wR
HeeY4MWvpTChNXFj3W0MYM6crb13UscxUysbCJF1zoFUpeVzxzvRiKr/ay+mmd38
sfrUMR23j6tV+hGnpTJ4D1Xxb8ArE83xDKLKsZqPkc15bU3vt3c8XhGlsjmtUOVG
A07ldorSNK5U3YloTfw3quLRPoFeWX6gKUmy7Y7cOwVRMhPjY3IyCkMkYhDRjq70
FOKrct55WqCJXRGyxK1sLvwkr4zCegi0XiirdqHqKegiTEu7XBxa1Z1TFmmMdYY/
M9VcJa8y6rZ8g3NgGKzUxD6Hs6GKTT4aigBHCXAYgxBnvtXM/Vqv+geIzTZ9WqZZ
RahYtzHzddTIouI81cMd+tDL1Y3nHe+FBGFAb9cdGueb7MYWfTpcjxOrYHYBQsy7
1PMPzULkkl0gmf7v7fEhRuTKUnDAkFzBKcWrwtEIquHkYcokEEZe/IBA5jqhhyCt
xlVGpsv1maiyCK6sIsLBUl7WSYYlE9ks7bYTPCeGFd8P5HF6+DMP8nJJhE7eesqc
puR4tzkh4aCGVh/csl1379AeDIYe5TA7uROc2QyuRdzHKq9yfmNKH7SlsgXdL9/t
7ocZDj+yXgdHv45l9g6esBG9DVB6FAFRvXEtmpE0ZuFGfJ0P2v5Ilr/JrOdD/c+s
z035gmNlFkSRYmFU7FV9icyRMXNafDcPcJTj0fgzghUCxzTXi/z3hvPqiOZT8lR9
VCyBYLk5aKEg4uXwEgbhpSeNX02MX3V0V8Mmst2IB024v43/aquVR+9eGrhrt0fU
9EuIY/VWpMiFWc5J47Q6Bpjqmkw3HfPN/TA0oxejI1ra3GB96qKV18lwsQPfvC38
zD3PZ2scH3wbdRbeY8nvW8Cg30hjf7/cC7scb2vaUadEgDLMKpeedQ0KSu3g7HUk
PknLyVMoSlELViwa9BDq6KsHF4SGmzCzlJt8jdhABEBgK8/ukGIi7oGloU8Bmlks
D3Vl7cOaVsmefABttvmOFP/eIR1cuYhrR5wUXATJazf2jMqqN1/ym+uhX3C6Pm6t
lxfo0aAV9xq/tJR4GsK6OxsOSd10mdaAhdeolAnUvLz0BbmWrDYWDrmVsGghaI1d
TOiHzRQ9gzaPmgJ61b1j27zZfMSdM3NIWZTkf/yIYjodMe7RzVx9HE+uusfi1yiT
PaKwqLg359iUHxf+ZZmp3fW5rT9eoFjPdMu5G4SuA6e5D4c5iX5hM3fNLKJBpkUS
QsTn1yaXoOYxrqmrDE1MukdTIvn7ZNwBS96LEccJu9RFH9Ck5RFQMrSbUnDNpuC6
O5O4Tqmpz0dn48kaXcgh7uAvFtY7biWJwc/N5fii8EWka7Pl9wLKA7oXKVS2pmS4
jaM/W+9pz4kd1UekBOkwRAlopECgQA5kuaDUFt4Z2RXObP3Fx9ANfmLkgH/Hgna1
uEXECFAoyKrsNJjI0wYeAZgI1lcDymCYXr+pblfp7b9xj4noN/du+iFSQ+BQ8B57
hOZMjQ5ye8h/nJJX/ipfydL7YjafMY2qxP1pc4mT6Lfa9jl7Se55B3qRWvgx/8kJ
wcGoMZyiNlNYM70M4FEismPU1hhM+kVMRcAtecvjCzS+w+9p6FCEF3GpGiojug3P
Ic6dd3IDPQXo4Akrd0HIU0IhqMDUUYtMYoUgPfGMtD8+IuFUsk6TtHDvW9fofRLx
FakoXYW8thY6+Kzct4DMNsUPpYqB7VQ575YfT8XrX9RY+sTRR26YkygFtyDwaQPr
YylcN78Az/Rp6boKcld4SeHCQp6N+PyO6Ir01IVCIBKA5bFgfLYh4iAM14VKEJGu
3yaRCt3kbGNYNk9cjxOuJbAaxiT//EMC7/oHIxIgVf0HlFMTvLoJFrqcYS8m7LJe
00aijDDDYwqpFn3aK1yErNEyOuj5kzoTAtp5XBnkY5aXhhEybVrSiC6vG9DGpQjz
uW3wNSUCF6OTP6xqI7xTPcjR5T5pcqxHZgIYWPIe/Li/H4mgeMWiwKEeLm99X2am
jSaz9AZtSyaQPa0qrLkm5H4NbVjjATgoXg1XtZCNYbo8psy7/0utXSOFi0lQyjnp
Heu7UXPdDk1rmej/ezZ0YhBayd97+xo/jPON2DXLY7pVZh5BK+Qt3TBWfkpz7Shq
wBJaY+pztju6yhWSz2/xI8AKLbzTRDLM2CkxwKNkNFns6ZlOLrKA9gTL3jOvSJsr
H0/n/8CJowGOeNOb2H352YRk4cMaMtjob7xEdAKNuIfo03+JKDdBRF2ebevwLr2a
gEiyDEgcODF9dQ8pSJXSMZfezqPufZqr2XUR2XW//G7ON1AoAP70I4BJFK4yTC5G
mVDqR9EF3aIwi66bI+wbye+bPOptRwMlzDaNpSD3i52Z7eujp+45q87UlSn5XSdm
vPS87cHgTUENSK6xNBX4+TKlQCDmzMWlwNCVvPsBY75/QnySD8xdFZHRKyWplysA
mVITc9KsQooW7NcVOwloTQ5mpIGjspU5ZQbnuR/SA8+lDn4Yb+cdzGaV/LgpGQ/L
7iKB33WI8q5v4a1Vz1J5QpHBweQ6noV4TIIxwMkbDqEOraKp9jN0myV2Nson/Dlb
WZzlivM7Op4RjMSwE190nmTPWhesTr1Q32K6mO/TgR5EJYp/HUw99ur9S8fJh+VA
ZnYdgzTTWwsSf9eeForJTbJV59Vqu5g/sR8cknG+4zO+1AlBtWVWAxup0WZTqepl
nnCFJ2oWXyRHioN+e8nsNtsj73kxo5/sbzEDsi6DG7e/MNZ6HPm1+hLYM8HPSBXN
KVN7nZwmnFsLlf4S21ZtA5DLQT+hSqSToViDrHwYvMVL6kGE6H3E1iPSR4hb9vEn
+T/jQmXXR3dIKv+JHKnnqeuJTXfl3/mleBAZ+DIcU3HV+Q7mbgh+REhylv0xDKHR
wBP4UCT34viArmGvFrUMYhjAnOK9NBhuXBQXCAt3MOEpebHDvVecpc2fT0J/bTye
rBmxCK526fFbod41LC/syv4p/Krr/Pv3BV3hL6uIMooZuxmWdTNVo+s1pHt2iboI
UbyGIxq5a5gJkUjvbC5VWJ94fbAE6kZHRVz5zBbAKY3v45MIJ4GRE8/YxhDWp926
Tdfy+E8/cY6iurZTiW779NoOoZku5d/vVExEr3FnavmxAbbV88KM9OFwM49h98yP
kNiQd5e7ZkjENqYP3cUogjT3dyPwX0OdKHqpQG9EjdQkfYj10MXt/nQULqN62I04
rU1Rn7qZj8YWOmfBxv36dfmgrm0Tgs0/3A6fAK4H7SRUclbmmpq6/OY87RCHh0Cz
22UJChrjXVDaSrEyM3cqbFcwn142MmwLei8f20NIDIxeO0eFMwqhtglrFUQHXVJk
1GE8XK+RWxCrurAb335FgObntqIBXqUrngdMSd8q2S/dKhgJOk+9pT3Ipc1xee/1
IBrhwOoCTYRke2845hHMKz3qQIdMIvovyHMRbKzsu3ouzMjyopZ+Sq6IHao9t4X4
KBtGJ1FEk8ftY4CKqmwziVbxHZX5cJEyuPJo7V4Wxw66HbTTWoq3rzQTKqBgc7Dm
/ieWNKiVR+l3Gny4arXlzVqDTl5nxp2Z6x91KGBr5E3bDCZyRYbBVhunzkS0eshC
xNeMU6H03La6DLJiF5dXBg7rbXa0JBP/SWvPYorv/3WbWUqgFIJS3oUE7maaHhi9
5DwV4pnuA4pq5l778BwbeX+fMDs6iESHOwpzu8VqK0279k6NTn7ArzcdPnLl1Z0T
bQpiLMFwmRD3xaBvE4RS6I6zqu0kMC7bv6H4vJrbNvgwdWxsFbKs4HhifLBOtUt5
94A9Sb9IOe1G2xEpmKMQXbecds2PK6J8Ybaz8LCPBACo6ToFk248jvhlvRw9f/YF
FT4uKXK9QK4pIMPJxJ5ifv+xWiSsQYVutMn5gPhiTU/3As8mJT879XdRuYKZbAWb
w65KNa5Psn+E+g3sPq0B62DEXnQv10QhzshVITl3uvGrLgZHJ/kBy56keru0U8pU
qlgARZqUEmRao0p3qsQcgBMHG1796ha8H0c8hSkQaSOEOZwUxHSgHWStCSDRhe05
CgSEDGvJm4fhiLzLUOg13emDqslwT1LwuU11fNeBJLeJjpUgoKBdHU0OkhKvJKPf
I9Mq3+ATPg3CIFnIIMgx4R91Kw8QuPoldai/cZs1udSJEEC5mqVUQtSsYOKc8J81
CqkM1+DkN9NhVmPfUKXB9ow7VzFeCsbxmAW/INVroucVD1Yw44Uc24CEWvQrWawh
tgmwc+RwsuY8MkaH6s3bkSUB59c2CLGqwUezhSAPjQlGHsgEDaxQ/bdC0TePr2Bn
S4DYZoaK2EqOJvdp2FF/3QmYPRw2+SNfwmGGNE2gV9z3tCoNvA/FiQjiOmG63JRL
YzeYPNJ+1Uyb1aFXkDfLOwfEjV8v18wiAKdXTHXTh8SLxEZDKGtSEpnNxDWX0U9h
wfcHuLLcfaC47F8c76YpIcljb0LtyXHxUhx9Ciu7cRp8HheSPwAZGauDdEfvBjf7
BZRPDceeu+xgRKtw+Io8MLAqYeuE5oejaMDda/XL6gmwTh8J1yW2SUtSmFBbbaLl
KzjSI9tJazWxeEnBixWA0j0GSWJM2tK+l3Ns5nNLPd3a8XcwwENmp1y0YY+j8+HC
SszPRhLltzFtCY8ipK4u0tvSV4VU2VO8zJi3I1SNiE91W2AQKQA3tnB3Smr2rK0L
goLKNagAHQJMBIfJcFgl8fNZObl38JJR093zNTfGb/Jghc/sqGJfffNqqZuQzAa6
pjOtV6z4xTQ2CM0CfgeStAS1cwF3Qq8EY0+WbsaWjD5+nKTckeD/GcoMJ7z80iXc
lKLAM/P8KLn2y5g+6ERhLV866uZoqksfOXzgUrl92CTfLLb/ufvD5zgOf+dppQi3
aZ5DD0muxO5S/pYGwb888GCjm2UHXDKCupSAQFmb2xtY1OQl8xpJRlPlppZL2Y+C
vi3Gzna3Z4PstCVP7dFxG+G4VwYXFQ5iDCxfkjlhSdrr46HyaSHs7FihIC16d7i8
tDRSpk53ID8vpWkGUsQe5cLr+45gakHh+j8+9zK7PGU3OlYx2L3TqaJuwnGuBNxG
JeSPcn6ma88odilRBOO4cp0jPoU+9IfEkTfr4AL8lFHYs5hSbTfj4CLPaLGY+qiB
a/MZUHxaP/Tk37nr51AWm3bA0wAaJKiPHMWB/4vLia/Ixq5d9f5U6zqFi7VAJAMR
VbS+KiJZPmC6dUtjWnRls+wqecE6Mv3Vet97tptepsueWKs1CaV6dwIr85mNpmtQ
+SUu3mcA9TPvW8AV4GLljTX+XtHjI7qR3UDG7jpVtKrdNcnXMkhPxo68Is6Vz9go
7bng5n96mlx2E2UMUWfik+AOiCDf04cBjIdaLOHz74YR/Di++2fEKP0rADMojhWt
aC6XQuzBpsrHuPN5SymRtwDiR2ThQwvgneVKiuoGXja/qyEKxy8bU73LYxvvz3dy
wboxOGVi/4MzjBOMnV07gZCPJ7YUJTyeEQjXMElk569lUaGjLlFyb/eGXIkuntod
dLsowQKZV+fZ5Hk6jqNsdQgW4Fwuqb/v1sx1dLsN0L8Q/j/KcK2KiEBtx7Md8rp4
wRWilziNo/KX+xHoqaEf1EhK5t4M02PAP2B+2LZ8Ciw7YNQbZDqrxMZA/bO9xGWJ
fKLVvZNTysHJWA8f4KLNzJTRJlhU4ZFoKOdPCCcNjHzP/MFDr9yFnTWnaPMhdCvr
HKEgfYTp0htpB/8zdo85G1ARmsLkrKTAcAqWWL1hNb8skKyz/GJQY8uOB4yzRCdl
4LXb9hZvlR4KPqGwk53ySjbXwBoSWLJ8nIqHtcveqUyfII+gKAof9eC1V68KM7ul
ilFh77sCnpUbIQoO3SGB/qD91t0uPuCbwpq3KX8yCE587rchq15d0iSLwHQOPXoy
8RveAhrs6UEp4u1ANtfdpo3T1HIe038KjnQCu/mmPWr+K5pJI7zkhl32IwvFvNri
J+aJUAPy621SzpQTkmiK0Ze/uby/781TC9Ti11KFtk+uCIdjsiu3YAplmbS0J51c
FMf6U4kJayDEYbPpA8gRofhpI1UOoPNXQ3t8mFDCdBFnkfNLgjJOsWgb6rrST1y/
SpIJ93HpWjh1wQDE6Y8150L5rOSzGaqwSiC0XtqG+MHNiabadQK3eXKYbLN1CDD/
NJpimk19sxiCH/Y4l9Gfmpyntqs0yCpZ6xrFY3kUbKy7nybxj4SLTXY32LAeJ3rV
0WHRaBUQj5BVhYiHyuq8BtPdDNfER8rPku3uhnrnYZasGEOibEEvNNuhbhLjTQG1
0wj10BXFTcCg/oTg/QCAAAMukVIoDjlaS8vqnoJQdrmIVGHYfpxTtVAfXy++Bynq
lU1/LB8xsnuHwQ393T2IJEs5UpLjtG4EFcaAsNSQ3wSfKT+R+e7u/p03PW1R1z0b
WDV0HKYc5NenIYFVZZMMeJGvudVl4fmq2BNhYDndrCZQt2ehtkj5fVkP7QL/ogeg
60g150vKuGuO7v1hqT5vHTaxDe1oi3KzgaaY9TivMSONG/jSoi/Eb6fnyrLPYJrA
nTe/ipEPRLxfRRnx5JA8CnlXEQQgVhoFE2HHA6dGgojTUsmJGurRrvU3AgC8srv3
/uMPrkKdh6RICymmV2s4/QbTx8mR8XbQ2ZSzM/5BjmuMQ6HXSmxjKMoEi6dFXhA2
L9OvrgbF58yVF4lwvZcgw2/tjQElks8m9mbaP1hVnRxRDhXdfYv2V08k2kmXiGa8
4dZ4xkZUqlq2Wj34nosBxZsrvIsLo4IYcTWZ2TvadMHx8l6fXSD97cKZC2bXMr03
oIB4J/+qEdLALVn7lHhmJpAu9Rfrag+vjB74HoQZE3rAhXCgmJ/aQzfQkEy8fIdL
N5io3wYiH0UKBMpP+cuudj1ePKd8tkkl0lFCTV5a8x82Te9+YdWP8ZpbFt7flV3N
X7JbfbZ49AW7AnsnlSNKPcxKgGP0QelJXSQhzwZkvLFY8QpvEIqvR1WjILN7zMYn
Vkyv/JWN2Nzdftp8Wp2K842n8Qwj8eRig8XFnAtWGdafw2ZURictAi8ZgA3+fRYu
xMZxO0KK0e63CVzf7kZ0cI341+afLxbFTKBcMIKw4K4utDpVmrr7m5g9qkfrPWxc
driJgle70c5Sy92iqDxvjvAKZpNM1SGe0heQTNEjj3WQGWRtWxyg0tppWRF+0Lqr
cG+jZ67EvViS3xvHVi0n7c4BVbTdPLWeBt/wNJL8QH7aVdK344gMtjZYpzVkJrIo
nENR9O/Na1NM3uw1LN6EnjOQHktPpuArDZu1tsFKb/3ImE8lBUZ0c4B523q4gsoM
qyA3d6OKjwba3Uch+Ug0i6zLMClYJVlhp30VJVPk63Qvt+qt+16bFizI9jcAA4H8
5ezdb2leD609YV3VNHzr0HeBHUYWXokyt2vSfHmZ98ywBdV4/vpiqBOjfdXODvGL
+Xt7Q7GkW8Dqd0WBXO/PbzVQa7bQKFntC6uvcAOjLBMrZxptUoFvWzNLoz7Mb0lv
yf1qTaFdrvOFpYhDAFRsHcltRuKr+KnumivkzQb9P1K0je2uqZ1nFf/Qk41F/dKI
mZBKs4H08zVw/TcLUFFmwC+9w7Le3rLMmAdDgKtsWZxm3OiUTq/k/MrEqjFzy6QZ
AIPXN6Lrm0X2yfxebkZr+y8ery02rNYli7MtkHCHi+XkvZ7s04PPyEGgaUIfEUYg
7eixG2UDENpn6AikZXe+V46V5rgQJnym+fvaYHD/R2eUIkXly3I9Jcu/Ktc1YY5S
H/+XR5YsxOyEnrBgt1axKztj+PVlATPp7S9g1LFhngjizlpGrVxNwYSprX/E0EY4
6aFBHfCXXw47BnhJ7Hmdt0Oqp2P+Keaa2FYMv+wF66JZCV/cP1mDqNDgPIw/lwrV
Z2B74mp46EuDTcuXzH78GJgex94/4Y0+inQdxwvqXy8nT2ZTrOOHhLwIVMWYea7L
ywanazwLR1WGWrC/r2UmiM49U4/JE7mQaSiM1GR1RHo3FB6GkzjKW9WoWX0OGZrv
+2E1ZqmpnhidiWlPHVUngkYHs/TaS1GX0O4HLN4H5NOpDKRrlkqGaQZmqF/gADwO
80gy3LYBBqKL2Y/aCGpm29pI46SLsFgqbqfTRBykZNtxfNgqWmLmktGHsSjaf0L0
AWUTWgMdOp5CTK8r5slsfv6lCl5fOe+2Fqz8jC3lmNQ5ta0YRvtBHrqRAUsD4Fhj
TvkBzMdEKnVK0l7/VWv5iKbqSS7dpwE2GEqu7a4ogLlkwcFf6D+ddt28uHQRV7KQ
BNSbgZgpKOdRdaeent88ga6jdpS1shaSZSN5tItSU5AGaVW2pLQNGAR9ee8FXk+3
SMBXpvTjuxuBhvjHj/onP5nE3IdtqvCiq6jtUpbJcbFMdsB4jKApHQoY8xvBwk8L
yNZJtmTh/LGdWfowRJEWWi/c2hRUxxm/OGRFuv04LtFKrJFm8DNexL+R/IxawtOR
SZofuh5k7Vyh6796D+T0vFY7VP+ovJBnu6peaz76k9hruHpPGoKtuWGRJOfLaPUo
7kPqzJrhhjUlCGPuIMasltnztawIWZB3C0fpLKVF9Ewe1kin2T/nTy3ilayk5Zq8
ATZWsToRS8lcosTlervUdOLron5K+P5pYW5Mqpj3CuAPzV7WQPImdIhbQmpep1ny
vkm5lgqHdKyENv7rD/ungKxqOFW5QJvqg+hBBbovPbFEvlLFU5HqV4BW3E7V1onY
DuVRP6c9i2yPkiY0+uI48FpGw4kSpuk+GkzM8iZvS2//LpryzTtiHvSX9N8l5dlh
nMnApILe3sTH0E02bizLP0ohZdwzc2oZE+9pAB64/Lb5LlnRso+AebZev+v05ELw
697N6KO4r5NJlae8Fv6kg4UF8YpH+TJYMZKVcKz6Ee/S0jDXEP2LdMlhmO5jQCt0
XS87ZGoYGruxKfFj2F1x4Vyq0wtz7MKB2ujyVF/uMSwbVGWYeoSmXxvlYEcznDM/
6alPslH1wn/KYKf/OTX2Vf5uFzQZgu+gH4J5OKKJ/9psuaXRy0jGm6gGbfJu5QPH
9kgFOMIJ1PKksVEWZnrcb1ZWsumsuukrdeiAZ7eP7CGVLy24lKWq4602CUMkM7lM
mWUssZlwWY25R+pPVrsOWDz9ucP6CnyR0iPsMWrPFdoWxx8vKs/gvt+qPaYExgMn
tDvjpn3CyPJw2L6SW0zrlJEdyE9U22pqeuTp9hP8Hs3LyyT4IW1d9xeq2mgJiy8w
huTxSz6NZVzigPHI3TVnoi6bSKM/AJbOpt3st6ig5ix1ZW/lrwMtiLJVVkysYhAX
YCeSthQXc+jzaDTeKhAfMf0dWgHUM3bGKfxYkPKYU2ieX3SvmcX4ntoOGzyz9tsa
1Kv8iISrOOqEGCzMinQnuUzvb360ukgRYjjhP2hbVKNGt88yGbACaLmrCG7uUXp2
je/en95D7UdMgpy6REnFlTeg5CY3+yYl3DR3wgjrzMoF58y4t0m/QuWqJ3EiU/1G
qxY5e+UBbS+ztLNkXwMRWAfhMiA1HGNdwZyqjHcFaXxXtQ/Kjrv4ShWqX0pWAkUC
MgDSsDvNLX8FcADcx4adb9RyyS4vslumTUSySycaqzBZhwy8bI7c3dNjvByhShUa
Bl/8tAOSdZ4+KIE/lgjiYLijc2h1XI2eLZXsXVyqn1FtzeNsLNKLLEt0fgnX/uZm
xSRQNdXPPL8a3vzwqMrBeKlxz4mthPhCTv4pksErb9clnKh6xi9Gg9NngrwQ8eSN
B3tYYPZfPaq1nHJTyjjOelxJO2fccXgjSpbE5p5xTBn80B23pY30Trt+8obeDbPX
p9rAqzouBIGSmw0dGn9KFEsenXiQscK9sN/Gi+1z4V/KDRLjVaTIZ0s/zLsiGhFc
isQUEmEDx1W4z8uxHMBuYEG6jOqxs4Mu0lupcAg5sKhd7hVNYgiEAIc3p8v11t9b
nYOzLabZ7nLyMtc+W8URm9xwUfq3GA4qc0tJfKXMiJFoVK/RosVHlJvMCAsIRLj2
JP69/7018dMr2Cb7/N5Xpae/sul3FVWlMEg1OKbcJjAr3CGnTF4kCM+Bl3cxTqfZ
2vTBrl49NEZorHKk1hToN7LwlbCjBeaDSRS5p4UnscQs+AKBaW5RuEWxlNGRoVgL
0fyKXxKnrCz3RKf6AddlJdKDSbVh2HwbyLLo/z7gaIwbUlqK/4LYyDJ+Hjv3+Z70
sRKtBs0lhEasBfsjfOTp6e+qkLanczGXkFQqmDrlFQ/j09MEgJV13ubKBUp6BRCr
urz6OQaNmH3TJI3EXK6zOeDPqZ5YpqN6r5+xF5jJIFW13siZGmHkmDTejVTaSQS2
XGTeX6QurtIcdmVQSaz2akTictLNUx0Z3oCtIa/vWdImoBG6Yh1aE+oTFILoDbHd
LICV6fFNydi0krKcZp5eTFCoc1TuMyafUEZvEztwE3DLn9Qi+eCMaldulEI7QDDx
NXVn5SxR9GNASFOqn740nWvTKR3ZRSSBDyB0N69gMuEWvH0PNN5F5WO8zk9pG279
eD75ihwQsIFZrVT2Gpyiaqx35XDFEEVC4Wo8PeO2LIbS0m/Wepmv83/jBkgRMm3u
GManvE0mfehn7kik/tCfa/ukTgRaBnKzz5+8FJUh88WHKH/L0jYhPhNxOOtj7vee
fvZ54EWFWaeYTcPYRl9ApR3QJ6KP93ESuhT2h23ORH8Lhznf5MGAvPBLeer0fs2h
vMmsukPZYc+Ja/tIujaDtLPFhzkQKgJv4TTXxA/LiPhPyTmFE5Q5E3dLvCBzbzbL
nJdI2b0kqBlnHjOIaGwV5YXolqiZHsq/F1vT6FrErNOBT1t0VBO4NXDgmcLkXA8m
fpj4wOelcUBky3YJe5QlEkLaZCS9AUPEgqvvHaEHnRmOXC63DEFmftMJ0aJBbGwP
/hJVyTqD+ukmKVakIrCyPNjhrTIvbQREoIu1cdWYVTi4sPa/Oq8m7mIweEdhmn3B
3JsiqPdXfFmrH/bFlcKDtVWtxHRocMnEpyQPPjNcNoFYF8sbtxMiK3l43mSsII6C
jddIEduaDyfZNEPP2l1EPHqSkA3vYw3FN+RgMmM1NPz0oDrTeDByM3jIS9hqfV6j
VcW+wQNffYs6C/PPQoQfdOkFRmqJaSI2jezhHH9jGQrNUTmMjY6C964ndMVbnta4
uzk12Ef4IHUFfEOZ4f1WrWb1KpDigPxXVOYrKvUrFuajt26WuovjHpijFR3Hnh9G
ZJr2/FY9kAwkxKEnNaDuNJm1q6u3g9I/9/HH1qfzxe1wJbldp/WKLv+dyGDS0UvN
Sx0DuRG809YJbJLNVPclDI7lKV8TQLHqr3lq2L4rwZg7+yTsbcWmj4zxji4fdU1+
dmWQGQw7uk+qfB3KnowRZQx3WKdljTCs7oMT55cof8oQI0cYCnihB2As1G+6PIP6
D0my1jqAt1t3POdMaYE+W9Ne5gFPDirsAW2Nng+qv2UGehjjE/YbdNgkl/dUhjqD
KFPfnotnQeqGyRX4SlpcZMOli4cpZmzfhw3S4oircc30251UFuPuD6oRDT2atbTf
OCD+JxE9u72ZoxT2w4/63Gfe/sc5QmjeMZRnxIoF8U8x8KhmrfGlBFOt9V7x3TwP
LklWKPaWX9RO+nN3l4vj9XPFLtLhshzwrpRhTmqjccXiWJYplkfKjUhHcLexFH4j
U5mRqNsc/CHTIaw3D6vxqiSZLygUywTT0UV+u69HMAGCa9eEvprsNeN0sOUm20Ng
OyaIUe3CtOTaq6nDlzG15QwWX3oT7HPI6umSfV6tkuF3xRslmKxFd0XbCUyTNeAO
1KMPRm1uJb80EajteutVuwAFNhJAn1M+Gpb91x61SFB4z9x/5KU5nb1TCO6Qzvkd
OfYAE+rPyQxX7WCIcjgVO8kzwiQbUm+/I9l7EnZhLPXb1ak8fQ1cBCbPEg2Ilqal
BXWRcer7L/2YwEY1npO/rt+CwuZGU4881AL7gjpZvAve49eobDVa9nmmurtBvsl+
1tXpjjXKCb57x0ApuU3Q4WO/T7r644kaLHQzUNzJNpajwaGTRot7KpSYbXtpOHj/
sSC6yhPC3EharLks81Yxa9i0UjLy1tUUmcyEQ8VIa4YJvBClf41Vog4Mkk1Sp6aU
iscF3j6V5Sg9lmpE/0VGV+opuRA0PfXkrNVLJxCiW1lkAvRPn57jabtq+I432pBo
vE1s3aZ60XUQoHuqGR5FfpUMi5tkjCJU/GK7X10iEAdbT6nRWitRnqTLYjMZcjd9
ExcqqiZqcygN45rghavcUV4R/GrDQu7k7FkDZi/1FdnDxGwVvb9ZeN218l084av2
tXMJOcVvIHBNfMPSKg8mY90lKxWHAv25mICOIQ9BsFulh+fUz0cuhPMFYbagW1K/
vfKa8wo1tY/VHVxr51BLDtuUn8VyIA0AupRmXXFWJlDJzw9ZGHM0H4UQI4DzH2av
jFXk57LtcYVuxAFqB7wpcYvtrjTmv6E/1YLt5sM19XR0YurW4CxXVXvrOnfpUsh3
DV/X0Whvi6EfsAS0JBHFGMoL7SyEcq924hJJ4VEIgzBlACc+orNzjiM9BSHmTHZn
8PHcMLz6QEXRx4Y/P8Kyg3svkOw48/btuOl3nh/Ly7fT9ilabyxubAnb/XcHpzxw
hbux5gbEDfF6qUz5kHk4ccOga7anCm/BGTfEReSlhJA1Z4NQz5wV6oWvpi0S+Boq
jrb3Z2fiCJd4eih8IBcpGOGEqH5mR4O6w0gnQPFQXTU2QJjE9HqvDdgVKrSjYc7c
qoSbTSBnV2zCAgeQGkyr8EiMgUC2i/MKZZmCgePyJWGwKZVaa/I2lAauENSHjmyM
lh7afHWWD+WT0M4PLnQDhEX7IVjVvPPrCXy7mw/IfQa4hRtlexpY9txeOKohRs0k
9NVk5+XS5WGxrFfzlJ2GNNWgVqVZH/Q1Hq2UuyxVN189LURpF1pKQmD8W24T17Ww
z3rMvCdhPXZie8dFfz8XflBFr6kdm9yTZcOz1vyLKKQdUijqQMzLip7QtHWZTECt
D8C5b7xMtfXpGczXuFccduSqSknFqsJSWjEp+WANdOorsee8T1/LvUr56TZp8vLA
vMao0rTfPPteHqWDNq1xouMLDwJRkJja6H27v81huE874rXRpwUnlEcLu1v+9sbK
q2vOKPuxBe84xnzNzSmx6CABY47mqRGK4p8SLpbL1Za32wpWtILSfo88s2PmTlPm
0P0L8m3y631oFSyLEqpLWt/Gywgx7OW2LGKQ5uTHUtbUhIy+MLSjKtKdaXXgW5YA
bc+XqEb6ivlBFbP9idni3ykbg9TUmNOEtrsuu4qjo8u5NUR08VOp5FckA+7cBQ1t
mz/WCcJz8vYLEkgFBq12GCtanmVqXd/yxj1Qm05t1swjVDXQxgnQMdrew+GLg5xp
vGN0f/sq/pUDz09kHmhwC2ymzV8whIGCTtrNs+Pja+jJMzWjZHlMR0hAZEHkWtzk
681FV3gIrlNwCiIzNi761T2V+Lj0h91JXfq2NwXtqf9Srg5VXbrz/aw7qDP9rwnv
F5Kr0UHZlM4cdZBDcMpLQqA/z1NuBjVYM3mcdnBaGHHi0V7nmHhsN+gppVy8LxJY
3HtYQ8WA8jPSKAKa/ORRLJqxIV0Cao5xm1yZyWvzZtPurlfUUk/RCkEO3E036ZSa
ayHFx5CrBz9JlFyikV/OHiwzhTEv4R2d81Sr3W3Hfuy3HBi3evJ6xg2umFd6R9hp
/7gkDWusiSJAJn06YlvBcfCNZQ8oQO2SP+nx5yxPkZg8XsAfEEkHZkO15omXfn6g
vK3+ICI4iRZ0Uk9C9t8SopqbL8TvQJY1cI7sYLrSix/lwrfcKyqr5rFQJDIs5PO2
XIaTE0++OdzVKRUJUXWpkuLQ2BY0FkqDHhCo6FX7SdcstnCkZvmzVWu37uudPcxY
xuPmU9VTXZG/AWY+tmo+V5hKUMXANc1Pl0LllT/LJunvA8UgrqCQOE+P2VuoQ+wg
2/g5rIIDjnnpeCzWVkU3ENTN/oU6COwU7x+wRHKwsb221AOxAjdM2Z91lUyI/teO
ihkaggv5ssE8KREhvE0iLExU+0M7UqzpDqXe4bUsO5Eko1H7v72/CUWmKzatntbb
rJBBKocI/YrFEVpbnGnL1W+WK35lBZtXPKYFmt4gD5AXKgVF27fGeBrUmWt9LbhE
34qyGIcFxCmcPIJETMZe1JIGF4Jv0QUtNLC08XabFtfW06NjBGrje5seKzmCj56L
g4I3LNGyCPnzikeOms3eVSbM/iCdxa9QwIsmqQbiMEXTNB3DEWhASGQvmeNzhzBZ
jMFdfrLuPL8F7pRJ5Kzf9SZmGJoDBeJXQuVzsugqB4gTyLDk9qKnIZ4QeHhoBK5D
x+RA50AtD9llPWHUoUE0t3TbGuLV8xUiUHHP0XDjX7H5Jk99WllXgFe+jx/b5wQ9
hd+jbONihfT/aQpu811hbdFed3Erm3n0CUk1Zxh/Ja+UWoI4se5vq8zIK4NXCrh+
wy2vleexotyj8ijjN14zk3xqL/l2KbTAxeEJ6MNkk8xFY4jhZKdRCA90nQSsixsq
8r67xfJdddZVBl3pDUzYlD8UfeNFZRCexPLFDxb3zVTPuR3Hjm5T9FquFIzCu16G
J8SUTgDddLOm/4hQ9Vd6kq8FkqTPCxvRk1JDdjqdILcGUQqdI2IujJrDhlV4/62b
qYyRMWZenqwy7uWouq4Grwk1Ey/3l5xuIO8VSK22vZmoHXeeIES9ei0zzkrTZo4J
bYV9+IsxYjBn912TsrAM38a9RpUSHvPrTAgyj1WXLBUdKYEz4q1IhfL0Il4ZHpjo
Naj5TA9bcTCKuLRod+XNY46+ap/aJr/RbXc28UrYEzEecaZePO4+MeRIQ1M+AagR
dd0dpo2gHgrlxIFT0ncEfknY1PanM0A8hEF5XT7FevV9gsLo3+mY55/KiF7B+mj2
w+3vvGaUOiDA9XJQmuL+hMJ6XLNOumzJ3tKu+buXJCIoPfsQaDvwl/yDg2ou6V2I
+uAhZe04zSlRIf/2A2ke7CSYwFDTP11KYvHm+D1tlnGLbd8OyDngM+7ulu1xpMEW
bHzaD7POvSvbuxYzCyY2HE7u/KM0gpQGgucxjiUoqlTl5LlssVqoL8LzzvvgsVP9
NGJ8hexz6Pd9j/zX1Iv6zlQTbvayVp/2GWLXCpCSwSMouXfNkde2Nr80pHChf6KC
JBDETvG+0qGlDjwP+4k2JPf1BESka5ysloDkvJm38Ocjrd6z/whSe5HSlUKDebdD
3FrdoRa7ek+KDnSIsSmC9YLQJ6g3qkr6vEVb2bU5Vo/xLHMmv78L+GyH8nhpKuHp
zWbpW7lQx7VWBhge9UXBXkLGfDx9SE/E8H+lxi4QJfWDrQfwkRMpR1RFR3se0JBP
6XHAZGwf3xLJRGWwH7SxrhdrQlZ54fUqALj/8JDrc3arqt4iw7z3WWp1KlU1L97n
16PuT4f8qH3qIxg15AJzk2yFkop4O59SriKGa0bharetwBPRCPT6mDXkHHpp145z
BmP3u5UQ4EhYUOA0zsOzN2eIhKZz4htXW7R0V3jvHXg/qXtJ0dJG50V13+GSB68k
f6cXCI2/kf4DnKgMsuuXHD/5mNDeW4TJm1YhRlnkE3xiJiT6HjarpfjluZhHcInL
xPtJ6hko32KZocmPhlv5cN+OQXL6YQF3MGEGJT2QLmYRvPPv5WA+SYm0NSfxMLSy
M8uaOD3MI2MIFntCA20ik6omPtiUaNM3t5GcuI6O3KDFGPZgtcMXL0USJJWOLJtU
ZP0pFhmX9+T/M0JdEMF97+/pxnJ7eb3iqBks0tfwJWIyqGE3KbH4XmNdG4WYRjWP
hFFUqQAMp/+u0773kBGheApdHPQX494xqz+KRZS0qz+K4aLK2sT8ZgW3vdf2Q3+o
8sz8c773XUTJc06rmK+VR9Sv/zy95+IfDXVNS1sBs/OIUgA7kJfc4nuicB8i6lnK
cE6CPOiBjO9SD6CXhjZkMWMF9sIm/GRNGKv+yim5IJL+K3LtrSsx6UO+TfMZoC8O
LgQjbkqRuoohiWG0/AD4OghebtVYa/XySc4nDWZMldh7ng7PcOVRVIlGEslghQDn
KdKBPU6HDP1qCfzYTAgS0XemAkMuvkOwt31fd0kfA+Y0AMx4q4DAnd6zBHEcKdDk
9F9ZUEDwSaqPJk5uroA9eQalB5uWkSTNWrb35wrAuyaJjdVhChtjtZiWFbDTCX+q
m4DK+33tL9msSCG9aHrLM60+ECeMzZp9YyDE/uwTQE5h3mMHhHGWSyKsh+Dui3qu
GmzNnb/F9K+XcVC6LdmInlTHunpSAXfDw2BX6hg03qM7hFWCPsmxbQhsEnjkdnbz
nsOlZ4/Iz1nfZu82Z5NVsWG3/ZckySRwIR0CIzpfAwIZtZ9Lkbjk5LjFXlzYkU7z
A58XEXp1BZEgFsZmAyguBmmhSYRIlLzqAgDt9CzqcgVMn36qbrYDxlgfFP0qWX3f
5ob0Av1mwYJ8MErFoJjcECY97weygTjWdTTFbBFVIugb/VQYXlaFngfYJ1IG3G1z
KWzUtWj+vwGqg2KxNfwUJ/Edau7RHWRoV0g3VCuWgE3zYu2Nkn46XVJtTnbB+tjp
RBaye9hWe9BmrY0izg+XumVsmBqHmTjxCqgW8mAPnD5vCMS4ehnyE/EzRCeFrh1M
Y2npR+aXNuxF/d3Xhz2BmbB8dSim9pYPpjqDwgxuxwut+ButrsZNvN6NvrqIYhKa
cKk0RHjsrUxtO4AvXvv5qs/u1tX8ISlqCCcTquI44ksEtJ8/gH8skzWfL66iepIU
7NhI0ZRBw0o7JSRZ6HX63NjXKVXb2jr6NpPAfNGeAakc4nOebEyUxixvW3gh1/6q
68XrwXP+DgI+OfkC9PGslQo/3+W3tUDQ6DBzAXPsXW2iBb8a1Z6QzlaBqylrdbHU
6k8AsT0+N4vlah0H7ZJp2gV+SqsZKg7Q6UTrTSJnW/admETqdy6T7GkRLOaV/VZZ
nMBg+PLB61b/iT8TE6ikaJXwbSlulXK/OqBtSPa3gCEED46hJRzuZGSl5CfCZOKU
4ZEozu6rk0ats490pqka8te1LPHlVMZ+5daSZg5fEMblX8D+LS2VNOTp6DH2pcdG
dUxbvS4K7+Ibmkl77sESFM+6dOIQRfK+m4CM1jFkf4a5ZcyFpzktl0i4SAL876MD
iZBWSG+IsClJUGGdY590N5JPOo4N7Q+Y4cB3GyEDuSJUMGOys0TcS2aBgBt9FvRM
dzGRkk9L966261WYtzik6C20gM2nf/oUNFGGU/Ize1AmQcYxcN2jCcr+4rv8Trl8
iPVi2Z3XytoPMaAPglkiDQ4+N2/eg377lukWtRQ0GXSpqVXF9/f29p/D3OxqskXd
DZqm2c/TTLArfzrwceG6L/cfRmasJwVu5Ih+z6bwKkTiAEFdAQwdFpOHo/Lff0nm
gJsKFixra8aSqnDpD0LYOpQreQ9bvyAV1PzJfqLcFCs0avRwfELNpqB1xVL+hRFD
w/tZDiBtByGhEyVEqUbQC7xX5SaHEfdaRGdw8gFyW0hyGJ5Ny7U6kCmDjglpYMnX
SERtd5kzgcBg8rfXD9I53P7as221J3+8SC9k+nLu+uW85ezZ6qjLoM4lX1gSTfCH
VgtP0Q+g2iLxm6h595f9+PwkoPsYdhr/f44ypNduW67hsi4QQFCv7t4PumN+w+kx
TCwrhNnoXQw7o5jEMGwEeOb8oUwv265ZZcN9AEeBTrqsFgRfuRbSluxfSEoMS7tt
Bigv9NNMCtmCqYeogopflbr/6GaUZD898G0LVmO++CEK7ttLWwmJMzealvYG3gnr
GdgY8T1V5WPsJqz60hV67ktaBNxX0111UhWGQBC4QxGwmc7m/Fcg0SERmE9bsyA9
AqrOL9vjY4UbBBGQ7vBAnJVjf1det/ePU9T4PUbEniTRjaxfwjHdqFeKlhj3BCkS
ihGz73wYB7S6kQ5ycPKTrjDCi4nLB9I+yvCQnNT+OX5dwyfa6f5ldx8lmozqnY2T
XbjzWfVTsgKOwdNxIrKyCNnLhElCb9ZRR319ekA29DQNpjUyg6iopzVEJacLSyKy
fGUZUXMok6ZY7j13kmhQXIa1Onw8ZDlKGplZpVDXRO+JUky9WskIQNyJAyncWsTA
wurbvXBb+OKJoVmh/w/R6ptYTT7kaFDcl78Q/wKerGK8XzK25T5AF96n1UwNP4Hj
r1qplMOawOO2lj8zN1EIagvekyFujo5TrqavE6MNrbh/noL8+2DLiNCrUZcQbSnl
hNpHUL+rUf2Q0650QqOXKTUDSLbP/dthN1GA5m/oxmHAWngLbXNNutNE1P/Ci2zf
E5cbUEnZR8WUeWT/pE2fX7pLkrQ5fAmhQEnP74Y8oSmC13Fbnx/jUKB8Lwf9ToxW
b8McFJG+JmxQ/CdktDu/llYvmJzfy2sj2HDvBr11G87j4Ul84SD7o6vqBIHBLiCB
GVhGLLu78/0U1hl2gHEh6dZWS2knFV8QL3tmqR2nFmRXoMWrLS0k0MDdKKuDcOcD
+pkxMCdlvZDYOc5nTeiWldtgA4pGWVju80p0CTs7sNp3NnRHySPtJRdEXXrai8pZ
R5lbUo9oRMXFXENyNZ86fWsrCEyqBbO5bcYiy1CPOoZ5NFsdCJx7dOC2cuYP+m6A
b9dztr+Ed3/lPRnnUUbG7FWQ0D7+sahjsRhDEQMsCz4hywLBerfj/swM+vBReWfC
UFQlRZ4GUq/JU7bgjCfnARIxC4xaYHLL64M1tkY61dUVuF10kL1xmbMXddMnIVmC
FHirm466caI3DY7dLwY5QohEi6U/+p/dHarnvPluU1Adzf1SILrB9XsAqKoYN1bq
Dag7IOAn71u/4T6MmqG5I2ItKOCfHOZ3TZWVEgRRg2WxLnAqdh6dinPMHMqFaC5Y
zXNCfrpomW0Pfx4wQHxiVPDuKsylMjGK41dR9XbYApmLXkZ9vE5Z/g504cAx+UOJ
IPhazKZNIIRjT4nl7JeIFphOmyNeTjvopAm4QJAHkx6wxreVbJrxcZMgWZ9Sjczq
DzzX8g0y9abvbQh1Q+VM76cKKJUX931Qu5YSTBLQaNmjcmEDI0pUNqPV9QGLsbrT
vB4sTYnmNiSoh3U5z/h6IZqLaAQAw18qkdpiq2UlPUMlXprEYm7OA7kg78pC+CzI
AvUjqU/lqIxde3ERYxyFkOKT61GxRGehNbblPuqJ9KwhcteHyKtDec6fPEzIAQdp
vl3LWU24JTnAZmQUgyOPANesbX7MnNISQg4fdkzB4dl/QlkygJmVeodiNVRkucr2
sucCAu7KATnCrK84umGTpnfZ/cc+uNdiRTZPS1Lm35GdrjGDR8LQOjL4Tm5fXK7E
+kviXuiY+NJmD6zsdl1ecCrdI4KYrWsAFuBssuO94yolJZXemUmgvaM4bqfSw3AE
tbe12W1SezDL7j2bOnpjKqa9RLHf/7WLXi2eb9P6SoBcq0Rz9diNoJH7W50/8phH
E5uVnhYxYjAFlw9PA6PebKfD7KoNhVX0WKDbzdH8ff16wWRpzbtYeiX1wHkLfgxz
VssOZE0plLPM/It3GuCBvDGVlHrlva432uurOcAbJZVVvewvECoAseEULNpZf4bg
0klny8gvYGj/GM18py2rM1cUqRdOZCHZGbWsAQeELCnsQqz1xmGk7hT1bC1zM0QQ
Ows2vtoeb7C22l+6wo4dFoZ0W+RN9LdzEfMtQb/teQnDMKt/c+sGpvCdVgJshCQc
MiHLBvyLJL8jExljWw28NeVvpmSHZLEN9SinrCZF4+ISZqvX82niFLdwcp+0TQzD
y5UVAbgZJvMhAripkbzDP6sug3Pz5Chs/OJFQO5nCNOhTb1bgWS/MoYmOn/FPaP1
vflHaktzx6jSqGplXDCJDXSFtt3PSIhEu3ypgVjbyHAfL5oSgE1mEa06NCgzwYe8
eRlGIA5d2vfwzccU0ZWtwZ7/7yT7juLtInmCt7MySM9bRKfEyG0DHyHz3GCnho93
GJWgU3Uk95eH8pHriX0D8uRl5dN31+OPiANlfgRFRIoTw+j1Ms6T0LGx6RRDIMaB
CThzSk21DGJPlifcUzs/uxY4KIqHjxGVaAZmdH7rwMgjmkY1i1vUNwhLvg8vdki8
/WPfqSD2oildEEASQA0+WZevO/Jo0r/BtGaRlrAPNJ+26CWjZ/c9mw6m4Xy+rvnX
B/bAYQydBJtMqm3eZGkUQZWQgMsIHAIE9Xk0vJw3dp/CFuIlKnzc5OvBedVjv6mP
pMh4LmBfxbRimIHjUXMu7ElMln8vZ26vy+2LrWRnKia8/NI0s67iYlCkOkHFJjlo
WGQF81P5fi10v5eEGMEG0+jWsWqHv39LOwzIHS/8m0v7Catit0VGi+/zUMAvEE/i
3xoPJxEFeKc8uNdA6AZlRnz9kRmw8g42sfR4gWAjKeY+zi2oIs80q+lq51IJuYkC
U/u93Vzty6cJAPFbQLl2HgSNfm16HmwQNgqoH8FWne11IpLE6tqxS80dSHV9/9oK
FvsVjT4tJMQwCzpI0zTG4DZPaVOFVF49XitDVyrEB4Ti49JNW0Q8yqaByZYDh4bu
TDgT4BMCcbEItSudobYrP8DTs/LC7iYc6+Yyv7zxgR0oZrF4jDW1e0opQ5au7YpZ
ikZOuYkAZ8qTqe2SA9fx00M90r0X0EOPg/lHrN+Xqe4VO1E9aT3uFDznASoFX4Fi
yaKgUfsQqBolTvpJFq/htcci5ow7mPpdoz/hJPjsc7mM+FNveWZ9Uz28JwuxQGIo
Dhcg+t4EQy3yNLygB/BVnUqXsvavnrYk7gxRhDFmO29Ch0X8D0Yq6y3pVE2IriMi
7BTASmV812v+9ZmiNhYeYgYvx2zcHtKdwhWXkxohrbnFkkJamUBtnVq9xcVmL/bj
uHnqUOrW9f4W/jzkC1Kg1aJJzWjd+Fsz494u+a+C/tk7FlcuPwZnOoQmKkjCEUN7
HaCj+YYdLfRUo4wuQ7TNPkb0b77RX5JhBaoX9gj1hLGrakoanYYuqILlRmKmemBc
5ECwZjfYf7MKOiG469CQ74SzkHdUqy58HF80GUbGjBMdvDrysOOg4MxDM6pJsZPz
Egm3YZ9jL6raF0mazxNLX9VCwaCC7LCV2Fj+mgkICDaV2Z629Orr/ioQO4NYAWem
fmsZLkJpLiiA3RaM8KejsbEXWwClrbnsW0/BmqgvqHDOCws1cABu83b1gcSMYL+E
fD0YGjynhbFV+8rj8N6l0big4mi6W9YRsMyJO742E2Ym/5GmzVZeRnPAqoaeG/hx
bFx+kJJOE4ua0MwWbJVWlnfnXibiKUU2T1EX70M+TSiu9blzg6xEkBrQ5XAqtcrR
YuIIJhnxdqICy6uju4a11hZFG61SJPH/Oe/po/Go7ZrrK5jprfej6o3+38jTbEJO
W+Jlmgv+oOizTvZPaGUs13/yHkIRgO540eoHU+h+qChdvk+7O8YzhTXMkxvhIfrW
uD6UTYSbI0sx5R8GrlPv2YKMSizBSEdGPetX/gAwpjd7c8qzeykrV0gu/mjDAj/I
TVvutOlEZrrO0V54kk00Yv4lDcbflPCBjOoBXSn4pWkPcbF54uzrvdmDCXr/J1VN
5s39lWULBUlpO2FYI9Ci9sNDbpuh5dBRAWmNyobjlQsW8kKQAogvJGxNc8m0Rb6c
FGyYXnXk87X53deR75e1jlRQXaOc5jurtnpDiTeM1PgzlH++MEC3y9ExSldtluvU
MZY0eYH4MBs7mdEYXlec7VzOO6SoagvcdmBcvxwHZI/n4EElxDgZ3IuU87s+Wa5C
Ztaom5PeLAlJob0Su3WNEdNyzzKJ/BgjxZAMbKHWUxWulXqgxgSpoMh89RbgHsW6
FNS8w23dDO/gqHnfwF2dKC6ERRKmQh+ynqp6yuOT7sAIPbmSbvE0TSUI69a6Z396
Yk2YKgqDaCndj0g8iY+f0SRz7jBngeE4XqT4KLXCdI3AHBKAKIYQKVxFnyD34wDu
JrmpvMOI1kq0g+V6QP2129ufNe6w/ieXliG07HyI6nYUH6T0vBgqUgAckc7A+BKO
caqUY7pEIBufq6FmzegEejD+KnU4b09HiGDOVNrl5uWbdoG0pbW9h6rQiV5YVThW
Js+k+EInyVTioanhvAV9CpzhyJ+0yVaHLXGE7siHXzNzyizeVyPwx/dBtI9pp16u
53L7Ad5SuKWlOGwOSbVqE2w0INrcWLXJPaYMlQE4Sg/bTYk2etW/smkar/yN1n/L
MjywbQyffO85pUFtDloMl839K322StlnuR1qS1EMcZT1+ljorNShm4kF0VT14Mvr
LqJMj+XFnH2wUdAyZx3LOnpR+g88bxuftRyOk44/ckcSgxjV95/NS6wZirbGdMnw
io2ULDA1VE9bBIaS90UPnmVcchYs0Ufd96COzDfOgF61Jte2z7nHJPAmLG92n/Ib
y/M6GjCEq/ObKBmUlkb+NYAe4GWQaE7QS1jkYt2BxrTuYosfp4rQbHk8U4n1QdnD
gaBYitylLaWywiwa1q/T9BX9OaBgxJJFkcnioJ+qQIwNdwlfZmtwM1zGkv56QKPh
vJHXyOg8XcevCLxxOBMpF6HSXk6hh1QsF05AxUfaONkx/lQzaS95qGdq1s3PX7ic
DK5UwntQnWe1QL9WWY1UHt1MfHChlO9ytzxSBXuXJY8DometTmam8gug0eVWXlnQ
T3abv8ts4Gp5Ikwtc4wk4dR5CCI0IAQqmxXmtv2HyAqZrTQcAkBJ0O6UHEdkegGU
km4UmEGHWoZVvYDFk23M9UTnbfHTHRsIWEmbmwaxf3PFrjcuXgSwwLtCK3NX+bm9
k3dbRHNVelCsFcgzogO8USdbNVjyQDGXaCKwauZwFSulSXEolYCrIytoF3E7cEsl
2Ic+uF4awCj+vTF410VGznq3jPCB1u6mJgcbu+c7zR4WkOcDRLsIXfQszl4v31lG
TyZop5chxHPKsz12GT1LRYKQ3H9gc5AXw4PHrb5gT0GwGskQY6hgACgaz7WOFugM
jsz+0WkXnpgXBUV1lzkwS+kirPcMHZiRRC3o1Z8RkEAtIru1b4BRQLNdGaS3zzwp
ED6WFt1G7LfQKtqtKH5HA13xSNZFlE6qDpwqLLJBK+Lln4KEzlDlHt1opjzEKbve
gWohlwHbEwRxB0pzgRQNGQnomaelnHY3ZMnZ+DsUnW3nmblE82O0uS6hOKjvJQju
Q/TkuIfDWXJNKsYNKyAhaP/uN9hdcMgEC7dftoCQX8quuKmx28TENJOMuf1AM71P
Mr8oa5GJ27Kg3ncNkUxd2LlJjGaXX/iIu5AOumbXQDGylq1McYB8RVfdnenDSIs8
z1rNYYN3ikTnfYS/Y8F1KJQ/3uqaWZOfNevLMFF6X1VQPj6WVyjm5bRfobWlgmCb
QmujOD1HeSQhGVh3FoE+1fHLB0JVOSTt8pChjWCibd6qRpqmqPPtsNdsO5UNKWPN
VC2aOOzZ8+n5hbNLKVHFCbP10nDC1EpFsYGZOVlVGXDhEKRCRcQYbNQOeg5ZzQ/n
BRTZmTh68rfPh1zJ9YQuQ5+wwPOvJE5gMxjz8GY5DeSSAoAb959FjzBqM8CYuJ5E
pVwEV8lSN7hBW19Krj9oj733GlaeiiCDYd82nBKvTXG8kS+2rukh/tkTalHdBnl3
5ZYKf3d0Y7iH27zw2ugNh4fWa3Kp+VyKD0R6liKJz+GiOeeSOxauh8+zKSPAiVYu
8dnxRH8tQ1flckMpuvaNK4RJDwR6ILIpjq1IaUK04SvRE0cz9Lg3K+jWr6rmz+iq
qk1eIDKXKg8udFgtv3PDTLnjtdfw51Rm8K42c3BT5IUM0fCHsXsSvq3j1QlKybL/
QuKyT1OjWOBzRlG85B0V/pmAM14fOjlq3oZ9ovstDNN2ug9j/NswMnUvuMI7zhnV
PebNLJ+Bnv7XI//CnzdHM5tVeMQUcXWcwUfZkpXpRse7hHV1avpmpJKox3ljZ3O9
/QibNAkd15h949pi0jKMhnzX2+PDVBkyi3sQzmRHZkZN98kS60ECwv/mQ+aKAZCj
z2rZMZVcUiu+tQDGHh195z3CC2QzxwqEORLZftb6i71VnqqcroswUTQGPCGZqlOO
VFVJ5y5aqzXmSBasn7in/1pappSf4AP8TAZh0s2+ZPhP5gRnWGN90T+wrzlhS5hZ
oU6xwRI2iYGEHlliEUnzhwcH1kMSG3IOfszJRzdya8uGC2UKzEJeEE7CnI6mqyxf
pfN0r09PbFxaY41frtIBG2O9gVBkqFTNaWvQ+HaO5gwWTfhbHSquz/Og198UwScB
POnF04Hu+G4ZptyGQXtgDe+r+YFOWmBEtQzqxP474ZCOmQ2Kmpo+FUOYu53+oSwq
zy/rlAzkxq5V7FEsbDQ2r8ZDg63U397rZsyJeX7c7wIaSTXjuBoByh3i51mFTjlC
OxRxYrh+KLm3L26sHAQW6wmQZ0OFjMjsrVtT2lUBMleCbpexeMh4u7DWKviMVEgQ
F+CR0lerrMzFDruQbnPuFTPaIruNvPfNxOlL5HWdofMdYCGS0KLi/8V68eMmFKf0
r4IMQlysH/x8Gd0I8gQj476yYz5o89deJjzAzwTFJOnpU2weMeVJlmPSAJEJg0N4
sZb70lvhk0HnP6wcMyYlRzSITLWzzEhuocphITaOa5TabeCYb4fEwIWORen1PGkL
qciJ/g2TpY4KqpXikXOvUotB1V3ZJ4vjr4+YF2h0aSs+HZu0Ja6UJDkVcpOBQ0wX
gvempU/Iz+aZt9qrNO7WbdLUfKij/wl2TArckGSGbaO0eUuNmXlMuqHRBZMVBhWk
v7z5zWZs7Z+TaToIn4i7478ZVE3W4C/iSuDGFWURIJcoUNLtRFM96QHyfOcyr0H9
TUPvHNkgyGFbWvirzQgDB1OLqwYKxtFdtDutXP7eD7XcrQo4rugk42PFMZVD0LAu
CyVuwQbtwZcqcDIcXeyH7i1t4pgD8DDPklX+L27i6PFP401kAQnYrvcT4tXzN1+1
bN4Q9izVmv8yzoQN0kaThbbSjgoYpo9ZIPJi3pclrfaAFdZVQ2CxrK3FO44ZDHGe
yA5fSWmDHOLHHcJ0GDh613BQ6Ef0ReOCkDVuR1SXYImIRtGYN6B0bLVn/9EJuj9W
qUJAa//CA1B38XASJtt+GoL3GwuAzSbZGfMWjzsw6YNUXnMZIok+3Gwkh9QNsmcW
bSarXeT9lrLpG6r8kunfHPm9g3Ohlux8GvRHVFcCu6oVh/vVd9KXJlg6ftm0D37c
9Jzi0StXGAzOyqLX2tG1lMXWhYCXd1dm5THO/xNNsdRw9nOGsMKFmAm3Y3wQSLtU
b5KXkO+E8EMc5L0wVyH4YIVQFkGdEU+mZVbt0RWVsI7SVX6cM0h2GwN4XvA3f/Dj
+e/6gWtaxX4FXyWBWL4KVMbmBYxbx8cDedXn/UAO7LrENNudBgkdHMmLa5AWGP+e
9zuE3DZpVp5LCuxk/S23ZmdCU52BaQDD4C/XDlYlT8tIxsUsayN62I/cnZ+zZNrB
1sAaWOedZjelRoVMzeY0Y1vaMxLm948jTIsxQxxbVL75/6nT8PRQizdlfqpTUTuv
xqwh3hbOxIlvtlZWfQfVxq35BSlVzGxu4taOzkBOuHb14QVZdc16sjXI80Nq5vRN
wWuAG2dK+6S9agVF4Z8QQAeNwY8wMoKJTQWBCgqv+bOT2K+aV2P4PpQlybgPIgK9
AcA1lN9Y3PQujaBBu7kt/ocIfzilKHItmbgKyCaObBAr3OHIXtKB96+y0VuxAbxt
QgQH/NZO7t2ecqRuVMuw5gdPU2YicpXKo8P55WHghK+XEAE+Wqj40gYVRrHqjI3k
LJgLaFrlPCabQjeBYM0HXKpM03LNJqhwKrrkGVxvicOCu2e9YbC/4XLj2ioDlVuD
F4/9tAVp5NiJ6vJUTl33LmKJIlLn+E2+BVmk6zCsS7OFEUe9uyvmFp/3/byCrDTY
oM78fqig7UWnmRiRQ7YWvW9Q9cmBJ1G95WMgUTt2kkr9SxHeYH6F/3Vi8DKGwlvx
07qLdgrfd7rQNNmFxQhDggByJu1iYj6588j06P/PAJ011mFdl0tLydhwDxWaRbBW
RCaMHLMNkXMnS9NFBGm4EMaeaLwkfkuqz52zmLivCB0jdHIlcTm/LgNs+9MSMmOn
TRFDiHut0ZavNzZlytODlaXQBdoCgS2HTulh7ejeK4a7OjoY1zGSTXl4BGfI7rBv
v3ainBzwVJhj67o7btNbZ2r58d5gqHItPU/zlioXQmiYF8wLdSDdpUpGtT2cjWIy
H9Ma6K0j4SRQPk8Zm3V5gRI4IGMlQwSmNi2gwrECUEpIYrqH6wP9AqGhY/D1coN8
15U5NK4Ts8mkrAv3V1tNWBEBruT9QmbtmN02jJU3pIBSGn1qvfc3fWOGJrPjgtYX
OfXHLgOlR/5JIRmDo7sfqy+vZXpKHQquSzLHVHAZqpvCLOnqK3TR6QnnzZ+CPSiO
MUkQH1/5qqxAbVFe61ALLn7Qvyf/ElIEeOa3slen3tYMcnF8sOqir8CKJb0SmyDj
4H1U9pzTEssIAtf2lZ7su3xAPhU6acZIuTSnAUT+FPirp+WuDKL2URYfnK0QHBU7
CbjTweXwdiPlbOrBXbUKJ1ukhBWck8zJ6YN7Oa5G7tVgqRLiMZNP5w+Kycj9lCfx
2cwtrCGjxjXrDXLxX8X0qhw247N2mIAE/7bHwn+01MypwQ0j0UfrBxbmrqJJQxSn
hkXdWkblVvxj5ljtLpDYXTIwJhX1/WQcJwSRg9zYNQZCcHIkwsyE8+apkb88OBRH
CFn1Oq2Iv6putQ/xCnrGITZs6AXIcKH8CEhHTlgE4MAFxESAFhYWQgpmt3yQ1ga9
1mJHKG5qQXuf7hWLny6zAlU0eEprLFERB+dkadzp5ifop6RTuSO633RhD5O4fd6W
82yjqHUzhyz6/lAoH7bIvEee30MvQLv0kZfdbWf9RUTi55oMIQG9JvvFYRdgwrWn
H1KV07zTmGLY3ah6l2VIUbaQmPIPnM0RHq17HGWgpd4bF7cH/aEx9/i3SQ3PuNxB
DFIwEreDfULmwReSmnb9WDaG/k/51IZoKZ/OPywCRzNtCZfwp046gPzAAN7tQE1+
FS4oUZR/I9F0vqgdybW/7/XzFUubFyJmPNw/oas3N4T9NC91UfuR1ZBuQTJYW0jh
H7AlpmMvH7HYIOXim2yTrnLgARRZ8eius2gjGIURwSliB9yDPMN+fAO4zoC8PPhk
yhdkivOhmi/RamtEWwuIZsUfT2DuQCL+4wG/E519CqzveYnhcAL3Mo4ho+AzTpWz
l3hRSPpwjcijqBUxAYEjuDA1Q2K2KQXz1AtmI9OfX6ZhRX8j8rs7tgceImAnsb1R
mIyaFQBEqcMmoKxcx2ZZt1AMHWlB9r8CyUXOjvlo1/kJt+j1wJoTTT0gi+v7+z4p
i1OpFmwrtiDqfpArJnTzxjqp/zl++TA7Zrl57IXOWowrWtC/nuSFA6gX7D4vpQlQ
9aN8zDMrwwE4gDZAh/w8IeT6PlIV86tl8eCY0tDjtvmXB3Cr75vog27hIjPwi8aG
QNYnjBwR+cG/drH+GqNQBtwle/MFcZRGewUbrkqE5JE1WTY1PCAlx9Q4R8wZJo8i
r4d9k93HLcSpVda5Ej/wd8yWll/qCBfjG9YTso8BugVyrwx61ph6EZoOo6wVOlRO
KwZEPbDtprpUme36yjqK/+b7BUYatRDIaxSuRAGKktoyElm9GWJoOccra2xyZvVQ
8YqMmrvF5kW3O63XQpGiqqakwW1qwYZvHGZ0ZCQPFOEpqv41QpW/3+R7XgG+2H8z
ke4XMKUlGTe7Is51RpITXGgd0N6hAKG4+3VqD0RTQt8Bfz3CFpNKNCPWjKScB7Qb
hy+TbqhNmDT/lI7dKb0tu22zLeN6T2BzF9IB73HyMXFBfxhl9MPQoWiTRuo05vau
4JAKsj3A/UngHq/5GVxnhawgUy1dI9Cv1/L9Qdcl9XVE30WmeCswAqzlXsQ2Mrjw
Ti8eWCRokUUqNRKM19jYp9O/0v54/opgSBtWYNgEwvb9LTpuVmXN5JkuDHX2Zk3M
2XzrsEe2IM2uXlVAxsfGm/DDZH6DBE40ebjo6YjMAgGz05RJa9DLOnqW+r16GedX
ScWz7l1nDcDMLiLjSRoufZOnO/HFWnZ5LpE0f6zbVGwTZ1X8Z728WFJT0ySBlkMj
mJ3/lOipHkUFBNNYpejCK6AUfuE4D4atGGakvAXc+WL81C2P5c+uYu/WekOq5QC7
BTraOzs2hczh4rX8g3dkvaILFU/+ymTt0uMaRozcZhW0uoI/dBjwC78zRXV9XbQZ
jIRE3p4rwhKefQNmDG7PsGInBLPEotN3QLCRNHZrW8osTvoUS/he4+GkOg9yDxnN
xDKdj98UlUm1vcJqK96TKE3jj15U0bxcGrzI6ggbsb1hqjOzZs1zhPox1c9SzWZy
nxn332fksKgYUr/phfp6sB/POhUkDfK2Ildd2BGXBci4uYRs+f0AasSpdlR7uv6v
KwNmibAaUuvxkso5OroNexAG2vUHOCOe25Lv5Uupa4Lka6JJoxBHRrXTO+3eKx1/
/WZTLTWmqLbzZtKI/j1qPR8tz1HglrOmU3KbguHY7ZpBXPNhq0dHrev1qtx89ail
HlFicTboe8VDiujVyYon0Z1hVV3LpCz+XrjdnXwXGZ/SQNUuAeYZ1FTto4eakfrW
8MRk929CQ6joQdD+dUeIbCKoc4YnpYUfRfCyUelrN8T0wUDbYCXogxdPjK5h/f6q
VT66Xppz6SsNOCXEWQQZs9QOaxPVXr6F5NDq8Sgma2pOFTKvJ84THagjsouiaMpu
eu/MQqKYP/HylVeexeRsfD6k4HbtuyyT5HE8qnpr1KqF5L0LgGCizrnF1zG3B2AZ
xakm8KHUk2FpZpY0ZhvZUnhkxTFrfvI9QIoKAvZIw2Iuz/KZ20Vw3HGxO+oWBzf7
UTj132axUm+E1RfyZN7215hyI+bo9z7SnQ3yacccIdcJ6T5xGa6arKkvJDnhNjWg
taeWrJlRbU1SGQdd+1TNDENuXvz0mqhL3Yio4UDFm0uyNQM/x0/1hSc3fG+wiBdK
NUhlQljhp8DL41pINes5c+99KWc2ErhH4wGMaqgPsQq0W/gGi8sgK/cgLAbJWcjk
H8Ld5esW76yuekiR9RENMj13gwhIPvXyLTmMBeK6fsQAYH69gBuQVHD8lJsUFTIG
X3egSspbkq9K5axUoDNDpNAGYM+KMYX2eZaDatwns1/s41SEyJ4oKkOj8nWEA50k
QZOrOZgszIgcE67wgedqSoaYNv1l8tG8myybM9zKFGagBCaYTgUCGEElK/fgYAkB
KW1ppOP2ivZkSqDb1qkVJE+XEmnwd//2UbNNnDMP3hWCyhld0+IbRwdON+1IPUf7
nhcvS1VPc/BD8YeAgviMbz2V5LBS9vpLxF3WuV12rC9KITAiBk4Vy7Ot0ONY0pxe
q0FJF/FQE68ai6S3vhlJSFhT8hyVTZqt+Vwlj6vokTyIDMPGKId/OooSUBNq3PCE
TcUm7FmQwXopcPXICWC354jaPDuu+TOttG5TNr2A2Dk+Ge6t2TRGamryP+0d5C0p
9nyMhlvRFTs0e+BwKZyry5/Tjj1yfov/bdDbU/fs8tIRGjH8O0sBKzsrXcpV2qS1
JJU2+i40IYQmrQ71e6MrNtWX4vA8MiYzcbZqxR3CY5OlX0pm51tiXw2x/xyQyPtk
sJQ4JWpnvA1qg59O8JCG+ehV3VFqSknyHNCpuXXS4Z6aKfAZt3RL7FEZrl1dFZwH
fWqWVreVQVQBaqvXvwyMZkCxROFxnUj1hYErbUMq6cYb4J+ciebLJmVI6WJV4Ah1
x4LEwDa+K13ND59JdHpkZzju9IznR+1FEBPu252dv/NdQSjAAV5uodySu46OQBR4
SXhocmBMOkK7HWQ7+oyrvOi90M5NUes6so1LsmTU0Mbw1de9hnqJmochyfOlmvyd
3r+dCqbP/mn797XrojfSUtfWlWuK5vl7aquz3c5uhZK0cE4BEzgFzk5cmFR9iSCq
7O7kFzW5peuoE22/PVGpq7y3ZQQr+A1nWcQvmgec9ykiJemubytFOEZpoDvLvddG
ngk4h8drSrDIzBdilzzrPtci39TrG/QkHT1NqxY5XCvdkh+r1i4jAu59G0CMv6bT
dWUS/orXcDIaL7P3xRWz+PyodDNR5MzLsngDhflOx453VGF48UCQDvLKmGGexn5l
6o7E5MjnenmKD9GhfO2F/dUYUf/dLesyh1CraDM2q3YndikQG9ESVwyURmRbJM2L
riFMu/rOmJm6B02oawTnMneDlsimaPpUiGtLaE5DcfLDp90lnc9zyHgOzHKRdogC
9ELNt1vRI6u7G62IDVd5BjAseHii1TdV+FgpdG4E3HiaLHEiMqyn5YbbPep2oA8z
JuJ0/s1/SlJz+X3hLzZe6F8IlTIwC9WbzKNlpH6+hOQWItkZgUDw11T9HJ1aE5Cv
Rii0seMeregdBfrFAqGXGkdLUhwC04MAoJ/q7gtV5/ch4qYlGeCijB260pLT8XEr
9oCzozQg7VygaZnvSbMn2OnUYHjPdkKu9rNhYiKdoHUTSZX+EW4XGO8DX0cZRNmW
zR/tR5gmaZpY5ICSH/WWAe+l3jsokqeynQ0uA0pzcn3iAUh6XHbGpTFAsQL7qKM3
8awdYDFOrgQdyAXdflbGFqIG6nnIx8KCXufzFbw0G43HqOKPN3i+SztDgK9qL/OC
fJ3wvmaGD5JxQA3XGKo6Lk3zi8hOqEggGrc/v4+rZcU4uDU4hgcTQdPHIj9NOjSD
xIqYqZ/Mn0qJ684o/DV3S/ebzSv7hl6qg0jPqo99CIQ6rjmCFzEcHKujFLbr/B5e
PQWC/pV2o0K3998tatOXiy7lUC8o6Eit34jNU04aZocskLQmhl3YgbIrtVaPt0sw
TeZZ8v8ouA+tHkYyPoCvPyuPamjoFERfYWbeXayhtcOQYafdDzB+2x7eIwyC09ud
7Pee55x2yh9KW9q1LA1YKlT/gm/b5ir6D6/d50Lev0ynNywhb0xLihzT92x9IViQ
m3XnFiOvI1w6CanKq9crkPeEAAixbKQy2/gPyqC70O3LZbt/XCJ55aPPPGghjVtD
pctLbeyVEbQ/iNJaUYKwJgEMsU1b4R3FeK9sq2j9ju9pRPRB1MfdTd1uJ7qSBdsQ
zuh92q71Pv08YCKeP7crn9puavNwpU5i0FzbatObAytllYOO5s+e9akHVez3qKNG
UeyyuPBY/K1s1GXnj7n7ANNflyuBTtQQMCcTLJCzK45K3BglLsvM/O8OPaD/Y7yE
utRtGxNc1ZzpN8/SgrxTjN+/rFw1JJ8Txps4g9IqpzjyHmel7wvoQeif+tTljvBv
l89+mD13Y+LSoj1B2haZ4heT+94RqgPh61OUj/m7TDJuZskST7+sLJTmzYNEwVR0
HN+HJR8XJZ661Myp/1wx6kwFEFp+0IQpIPQnQUaCwxUIB8y/XMwQ2hNmS9WvMhJQ
7m2tDiTwYJOTsyAndbU9u1NhUvJpu7nw5Fa6DUm1HQ+Ao1FICXNVyVJOuVycoF+P
aIOA9sMqDJVNBBrzIoKndPU/0X8hz4gwRSpQDx0nJFiQ4riLTd6B2vWk8MkP2ZEi
xaHtlRteXzzm0UhknQT1MeRCKv6bFRvr0k3QY3eFgT5fVKrxKjXze8aP4iD+CxlY
6mN++BYB5XbW6GvA3HWlKjJZ5+11r+kM9DXKKj7gazPWulfs760EQMaDm5onBlBF
Dd1B2LWcyezuz/aSZx6EhYf4DUjePJ8wEHrQ1SuGNhv+WwtNpfnVTbxi/2eSBnkO
rCbjef0oB8FdcWzO3JPe2GfZi2OGBFSazpPvkpbezTCCA02clbZgWPsdnf06WLAZ
bqmrVwXfYVvO3MUPOQg9bL7Tv1csVx0HWBY821tPfRtCUZTreWjTcVPuvi7cepiM
MfLDOe731taGDFEtjq2v9raww16rSywb+woO60zH2NkY8C6gbYR/cnpiMVCiLllg
x8h4jAbo6kRm+5Wl2kXM6a8pPerFjYaUTmNom7SGXSCkcVJVZbVFHIyRq3CAUN27
lEXNPs1OlHYsbvSSSliK5eO/7jXHN5lCSap9gHKkGfQ/V+mRkfeBC5ravFnve8Xb
/V5s6whDd1/xzGY9JT5jzmVKBKRWjMVgKulr2ekG+NPS4GbJoaA2p03tPr9LjeBw
e4AeZ80/cWcybd37e0w3nxGbEe/CPzCtHD7SoTBC6eAlh4FYRmuVioXVUGCJ32Ui
ETOdB7r5kw6zEllWFnqj1EuL7gBvSuGCtI6jzuWjqEu9eJI2M+D+rnK30FoWmiYv
6EpxVtbWPkHBBjYVAG4cpg9wAXT7S3FpbZL+bmg0bvNg/6HL1E+LYU/THpIvTr9+
BhFJmfFH33kPmLHh9e9Vd/rQLupRvHNr20KYXxa+omw6SozI2MkqyeDO53WkOIck
pxS9PPw+dybOQjMBw4CRJDE2Rs68CBY6+HihVEcM7j4Hzg26cBivvRFWQBaEEGCn
pAdW9dZO4dKST5Iu17oOlBAFVUHmKguiFWP7n7F0RRGnINI0Yl8/7C33dI3gg0lb
TD/GZuLMUZIrgyo4Hk7wFzPF7jE9eLYSToxAiGD3B8GErbUr/FCzWZau2IggZ5Yw
rF+r5PJ+wJHeuQRmSeBP2+qnaKNeAjXikCHlc16/RUBE9PutQiEQv1l5gUEDCEza
p6TuBIS3JUlazpH/h1T9WiNdCobc18si7D+pvID+sz4KfDcgRPx6aXPG+NwXruid
QyAJlvExhduE43m8D0Aux+AZj3klxXuzkKW5KVjKIy/4Kc/8ELJM76iUqzPddi7n
VJrqyQ7sfblaVk0nG/cBWwq/IWpPkvoYNBnGEkYKxcXMVjES+b6nE5RYAnWYqBBm
AtRfSh95vhYSyMYgGyHebu4Wj+TiDnVYH3sNzbtFT98khmrJVJNAd5l0Ii+NoHFs
U3fximNZdbTlvg2T1+6pYWu1b3S2h2TnjSxIpVZh3nHlpEjmw95aCnCEgUCvk0v7
cFTkcz5U6jHNWcmI1CXLVjB+7QPdzSo9mDIww6i9VJKcTuBUDKTPSqjXGk+1ir/i
B6cqEqgkaGXyI2d5SgICIEGX3Gki9snPj5BFN0dNhbS079eNjPWh4Fgpo0TOHYkW
m1Q1XU77MMA1yFS6J6zrtlb1j6ey5Gqpx/+4vlDuVkLYHl2SHty7RdZY+Aiztwkw
TwITC9lofclf33EbsJJuCK8VoBoQB2uFKWe+pWlQQ0HfS//MaBkhJUvf8924PPB4
QOBlmrnnU5HMg3wS1cKMxp9d2zmIw6/R8udtJlEBVZ7IJ82SkEkleSLAWhNc3BXd
5xV/34WW+9h58rZ42wrRSaX0MZ571SK8nkZDHnn3DQnR9dazWXC05HqGGq2H1v8e
M3ilHuBSIJkI6+sCCN4cYgHtPiL3+d1IWEzikb5ubEQCCmgZKqztNCU6n1JwR2FW
+yQ38hXHMkJpeUnxBYcki1kDxeOmHLC6FCPmKVWzo8oOOGB31ZwZu5fHwntz7uzc
dYfMAPzDewkWUimQCvwLXXmnVxxkZXfuJGWEjymRnPqjSxNcmtVkVJqyRMsBJTw4
FmPxikzPnVhcANmyCMN0HXXq1TEPwjwrC0kIWUFkrXFoLefntpyquL0rMWZqUx0+
egEWE2H4G5hDkl2uqxqeVUMFWVvM8Cqdgm3PHpBZSOOnEhsTcj7gzPESdaa8/WQc
5B3okzhDCEHKL9zDAlsKqDMB9LJZofNjNvt43jeANHbdNG5qyy/VjiP461hmIcw8
q9LZvOoERZ7kMFyXSsiArDWSflgoZgNBYmPpUM/LT9cnTtEWcEaQ3z/jk9/xBkHJ
16vf8b0x2vBwpTJ1iCaaTcR2fknaPywYCOm/u7ixbk88lYtNvdBX5x/sy1neK5d7
02Q/XpfgoeU/IMhAggiC83CeuzO8ck8Gx6/Yak+gGqMPV8eJDiB7r4x8D76nZdgG
VMaREfrQEOTy15udou0C42qsaS9Ykq+cc2qxX2BSV7euG6O95XLnMSazScotNKPP
bkLU3swhM5ozHNkS5fd2hPQpPa1NKzu5ob/xOetu8xW4d/zkldFt9jqw1zulZfay
CxJU6VeJPqyGw8QS20cvdlbNyz8kLqpyHH1J1CuLXKdm58LMcq1DA6p3G4tdYn7D
ayt2YmnS8+FNLJOmKz9t9g2MfCcOlcIPVUYFW06ZgaOjyx/piJ989UL5GzEBry+T
wZt7RcrLXOIGMOjmM05qOYfFlK9S1ikadIXsLE5K7m+umQh0raV3f+te6iI4WtHr
MOgQQD4gA/uGpIKAVcT/Do0QRBpYz/ZdDPaAst9eoJCZZNvFbrd4wQd5IR69PJJp
kk45nEUzA1M++3+QF2A8AjxRgYIDM5lbg+lWwPLPGPVatO5gNLOgMyeam9f0S17N
vjAKzb+ckjCI+lpgeXJRIdm4HchydKyOMKPMMwZ1EaCwnNW6gsPFhY87gCR+qbmx
nC0k0kndRKNjSQED1Zc92ArvksPGuan9upPgEJagF8Ks+iyw5GecrxDtcTVnCHKs
VaSC7THRuwQO0QAp08svqXsmbPJ/dSnipJ/B+3e33O98Cg3C9hqFjE/YfV/AaTeI
AO+whS/C6JWA69qKNckRoZPrFbe1Ezdk3qIkPPCAp+dXWKAqQa2Wk/yZ01z5AZf0
DgNP+AS2QpyyE8j0jbFa9uMyh1Lhv8t1m+JjIltbunhPNCRrClpFUvSRnVwu5nqX
ch1Z7+qHkW4FaarH9ly+wHzIRLzD0BbwAQZZf2NxMut6VloXk3anNwqSoTBtd8kT
lz0dGWxr5DRc7kOIwxAiMsE28xrzPBqTfuOjgzPHe7HhNsLbOPReukgl/0Vj69Hu
o6b+z/28khRoWn67cNXre2KYHu9R24B6n/2eGU0gjT4kyfJdchSj66gsEDiPtpP6
y1VRjqcsc/rLvXuEB5WHJ5SKYWX0ti9/lhL9M2flaUVRVn2nq35/Hrx6Hb1rGDyN
eGIo+nFSVFZy0eospBBOhGaavNBfd97PSCuSobZrKlzeoCR6Q+sevcARKzq1yBqO
vgC75zbATnA1OxMBiYuKVz/Nuy2I8/44DGQFOI6z4eWMkCXsS92F0oXKkZokloeE
FUB891WKZKFlVgOco5Jno2gpsFqSGnuE8rHK862YqoMX1cYt5bPFJfxdyz5haUdd
eZLIXnshSk1TCYGkQPq4FxkzMRQeYQXV/IzyGc2MprDWCEWRlkcoPL/949Tya+yA
9kh1i+Wogar8B8XgAH4bZoToVMzQLYj3kN9F9OS8Dt+mO7I5bpf4ZqKt8VjWljge
EmEWmfgY6NETxqz6+2oxthkapv7AjUPwhP61Iy0tUkQmWytxfD8SyNizTjMRMZFC
iDEb5tqNjXwdvwoP8WbFNQqN8ItC+18fYmA6XZU5i7s6eX9gumaMxdmrrJpiObyl
vK18PDe0seXLIr/uhXB0q5CUWCEq7Ira+2OGyKQTMPQQjEsm57khixCtsEBMzrtI
sEuWRS71/xBGIVJ4wlXxXHXDPHw33ORghxKl3GaYSOhHLe1m3rrPABx7mHC22eh+
0TDhH1I+NP05BYDQi1DEVKHP8/cRI67r0u1RTHi0zToQ5c24iiWH7Em0RrYNfZu6
vFC63rw3I/D/E8cvi7N+KGrO5u5oQXfMXCUu6k581ovglARlR+wdGmvbxvxOQXS3
2OI0cDUOLtIt/BVM92xzxxgbtkFM3lESE7b7/6MPhh9Z5hoIsRSIf285sxuGuDyw
UMzeGHY2jISnG9lO36X+mbNVxthZNBsGif8Ksun0RzgGOEmM/hZZKrehntoYbG9t
YA4Ve6aRSKYfIttbMwHp0dfIWItD9StsDl7jwIFlYe+Uv8bv9vAWIRDZzT0GX0s3
QPn7d33I+TZuGCK/5UBanZk+u3HSy7RkOMeVqkkzn63K8JYh+WEx/BfaN1YwtBwF
iluWjJTCnPwS8crvNsml46djl7ipM0YoE1LFcOkn5wCoslv2r2XmJr+2GXb9fo8K
/veKFqAuBwsUv5SnppYx/VRz/lZt0frSpk0n4rGw6JdLr0FlveCmXiFiaWwOuGJm
GB2JZDxg/Bn/dEKm6WZF564HO21y70tbaAAdsZv8cqdzO7PTxoOKNjb+hNb3V3+e
WyS79UBHGX649gUVqJrgIvbLRu4xghp/rFM1xSWfV2UFX8i2t5OTBRBbwUyBEzI6
ThkNFLJQmjt88Dp84eu7dFWeE+KEL1X4t5YXUmK72vw7v/iTe6M0a3VY3Mcr5wvu
KdhvXpZVPCAP1NIgflMWUBqF34jN3LUbn30IaEERcWcG2EJYbe2wpAFhhMY8I034
0v6ULagw520uwgaOQmIOKI5orRz4UD2D7qKLPx/DE9/HHJn0ntDANpy6NkON0O+H
PRtaXCUrCFh455g4HE98rJg5/d5EDGddZKClv2/xlZq9WEyknc/Bgxo/baZl+BTx
xQEffKIG00hFdA0YnqytVt6j5gCX/TIdq4jSr9cAi/Ic0diYfcaXMhmVtDO6n7es
6njmS9As94FB92gLRe3ZeMZ2rOwTxS18ap45PIz5haMpKgxI9KG5fuiZMR53yFoG
RgcAQCov1ThJ1xSIwAWjXYiRe066bQgi8h1Er5gR6RqpkDzOiDyz+NJtOLw6jVzd
SkHa+hnIILSXtBcCvO5/IoE7JCKHwkhf/BHLtibqkILGgpOsCrpX+aarDVRtFdfv
qUp4mfTWy1DKpdtg8giQmkMiAY7LATLv+kkZEzyUF1bzCyNxKvQlteoinz4fuVBE
DeKLJbbQt01yeenrkOOxLBFKAUYTi26NFmgRdL9egy3h0k8PwwHlMTfKxezL+j4F
jM26GEeNvgfUI6oXIQnAYVYcLzVR2JM3ecytwkksRB8he33ZVfwIVSiibBie6KzW
6a6SfY5ihGQiWQpwjvrUcuC0Pdlo8ARU2XWjQDOuoiWk5deft9cPCFHzf2yvk8Zy
cOT2Zy8ewAxPLYd9YBRPtBDMckgYft0u5AXCHgGRXbhRdmMt3t4uEo3NbtL+SpqV
W3GxrSP5qmedvRV9X0UscXCdkSNdUov2coxqGleNzu60MnwOMm79Jjje3s/hwRua
qMHOTg09WGdgIPgrc65AojdB0dkMeGrJoVtLC1dV5qEPXf5U2qX/czhe3WrcjuhY
Nzbg9DASBVfuNcHXJlGhn2FqC4oA0N/sZ1Jg5vqzXKbKK6iPerNdyDC3c3zz4sj1
pdTbtXZTMOX38KyhWDrjc8vURV+04cLr1bvIaSEVV7fW0DqtIpMGEnz3WJPWBGAw
SYaj3RMYwjgSXGjyjp930+cMnFcPfECHx/6iMYHX16H6FYbMUyT/V7+Y+GCVCUWa
9iApDsLzrjb7Bf4EdUTnBvp1X0sagIreY1chMYsYLa2wwistBzMJhDLJuLzxZeoj
sYJvrpm+vosMZ7qDKneoqzamu/XC228NZ/jIlN6rvl/mavLhuhG5/RuKFiMv6bJZ
3c5fWzpR3+VerGqY9Xr1zr53c6sDQiYrD5BTWwc4DsEEVS6xey9JsGjhgG0drvp4
gLewRlSGtOtluUhlMylZFfG+aYMR0yDXDwft55CbVQ4VqMmDKOy9S04rJRk/VHwf
yquSH5eMkQ7/sLKDhvzLVIdbijU6WMyzNU+DW+g9KkNW3B/nwrAxzYDHDY7qOYlm
YcanVRhys6LyJp8GNZ96h/0n446VQr6pflpyaMzWXrTjGsMtrEtXcVJfE3NXuZ6G
wieSbCLhfJ2gcurauBVmkS/vf3PXD3G18SQMkNTVrMPoS75b5uLO2Xnavd/vcRyf
jIB6FPA/hT6BRlXGfHwpkdANNKAgsDyN0oEO/WSJg3nZZei9AdoxWtoEL194r0ul
Tddz4gW6XPgf9mmrtxvUmVxyYfqxZkhsYEsbCTOBNpkzd2lzVa1zLKme2UKziTDe
5f1hgF2T6CCdXQcI1ZNEyvOvM9SLzp+VqZTivoyI0KTNXRh+iRwHmq19t/aTa4zK
ERZ1jA/V6t8l0rsncvcanRtOyMYMhG7l+8BQ7lWgEHDTMoaNtYoyjNeAf4UjdSTn
FSjD8mWhtbI6X/U1PV9KITWObK1E82qcqdkEcZx3UxIURqYAs17392JmKAHpUIbo
0llMhDrI3WXWfCNHCe1mhP4wQEJnHGDEknYVbHMqBhcRccGftirzGOaaJ5OiIVt4
/Pbw+95gDKJv6789Y0KIv/bG+gpa1jlzCRHnrXY0H2UTcMu/aPykdYpWyxOknFxX
09MsLED++16XupNoPZVufcWnO1O1j6O8VCznoVNlolYxw4dNViFyGVxL3ODFk4+N
hpPz6dhcq3UjdO0sEsmW4KLVZWl+0OMuaGxSIGlqGfTtX0U5Fa44jt1tSk9OKxPu
fXjkS1eJXYtZHBsgDYS1FmR60OABVr/iLk26qg60BTHhAK1y3PgqF736t45GfYSv
RI/lGtLRSEbiJ9QT6tiz5nG5qiUhGpyPtef+8/5DMV2CKkZ9qCJ100FII46k8kWx
T5SDcDLYuYhg0j/mhVjpeGPoWbXS0sYPgs2WPSmuZ+4xkyP3nzz5M/99F01YdkZF
dnWXzCM3WGDPoIx/yCMMrEwjyl5Mu5gnqsS06GdMbg7dwoXYUOF0TAzW+O366GTA
hvcCT7x5nAhB+E0PiHh2KLQp7OluHcoPHnbrTuN3/JqYosj+wNX5fqogPsJ3jpuT
5jDjEnjnaHqLkm6+nCoKPnB/DmbgX7szpXF4p9ZV+3IVlzKQS2TeJBxgBezNE8cI
MBav41J/fB1o3BsiOT229VakYAvG4aZ3SlsJ5rIVNAMx69jcQFSNFwT7KrojP62T
bm9asZ/QJ0WRClPPYlLrU8L81fP7lge+h1q8M+b6qmt6aTsg7GZT3NL7WRPuPCky
b94C9+oyvbyGH8K3HhIHxy8dPqeDnq2IpiuAIwhYb0GRNVQia8XDMym+xsi+cUP/
Hxv8d2gwW0Ef9egyQSjVAq9qVqAdw6VweK6euTp9GZxyDE+fBrX45ZIdr2m2nOS7
kCYy+yvvSfNOxnBSGK4W2UjLG+VClMSuvU2TKDtp0cINK8xdl1GU+NUGviB1n3Mz
shdCLvv0o9jV66uszddS5j3iajjECxRORTHI7AfIxKTx/eL6EptmqmJe/HpcilPj
JXibC5KpmufcYHwKdRv5fn0H/Q22qoM9eQKrp+u3HDTzbGS+qgjs9vFWSL206w19
4+WIiIzDvRzckkZu6xdKTsbTq7HJMNCSqp/oIQfMxIiSxo2AN64gjCgh8qSWaojj
KZ8PZzRTiMmjTJcKQ6k5YF4vgfDjILAb7VDhdoX9AsqRFGZy5s3pPKuOLpGJFLm7
ooqX9CRIhBdAS2PAtVme4Q/aPD93x2tXfjVkbFyEOnlJpTxidLHzY/7eFUdQaBLu
pdiMoeBpD63ZMlbgY/f2JrP4kclK02W6DQzya1GeSMC5QBof/1WFQsihGssmgI+4
IJ9UL64lesQf6MuREomFTTMmJinWdLLwg7e7xXkspE9vV+ZBu76c9PKJb0Pho2Fn
jgKR2jxiFCu6t6jN8e5kfpVzblTZ5LDyj9rvnQSlwX41O2D9q91mDWwIi8e4gSKk
0054+8tB0YOIVUhCdhQvF0U/1/owgm2paPqubC0RzSi4k3Vg5awAvEJAQsYVj6kI
5MEhUsnahEb8GABg78CArD1NGayi23v/1160zvLlJWBlxbllGLfCWtSrwWY1OyUY
D4hK8LgcifeCiWxyG/1IRaKp+O6Gi0QHZ7scatnDc4kHPUVIzrI4yLlyhzpNlTbr
rj2JW+wOavU274z5CoYmmrQJy7PbcE6iHqPgJhlQTBDtk/jv0jErueH72zRqnncH
VvsMCTlGoddzFA9aoyDm7eat7ziwmHD7oyi+5A569p0PQBIWpo99N7iWhZdlDdae
oi1yfKyP9fsGncP9rSsQK9NhYvlIGPFBdyangbKWVUMxFdVC5lwDFeU98TbuXSko
UAErtvoZFhEE20eQEPpzFIoHncj1a5JbMIfW5MmKujuJhA8IfLRjpMvvA7SXGloI
xnGkg5YJlivLGvBLmrmPBWn7hz3moCfsinT/cTXKR7sXIrwwyTCPMMhn6Aksp2ZT
iOc/atjCxmj6a4wdQm5q8ROh+cyP3U59Inb+oQHB/h5LOt8N/atozOwNfLUFE0Q0
Get5zJzp/PhBkMajdJkESOtlo8PTW02aWJFI1jyAuFzKEB7YNHxXKe+V3FLUtu+d
/WH4uk9gKIJvTId9AbVg8mh1z0tJf2rL0AI1aeZBnpcc1VKDseYZOw17Oqha2Tvg
99GlGfOSsN7YzhLPncHLmfwA5NiR43IWedk7weDnDldwv8o7wqL8Hxchul0F90tY
ngRGa7m2Mgd+An/A0KGYxv+0fxyByBHsVYLNw1NnSmq9176E/wfViGiygtD5yH/P
ehUAA57ciWleeaYcwxo2Qk5mT9gSlKv+zgh088wvvyA/AuoNfPQd3vKFEqflMP5c
rEWP37embEhQN44zkZvK8a2p5H8Uxe05s5CwCWfSlI50i3bSXheXHjZCPldAu62l
k+CeDkWQmnXGfxJ+C3YwUTGj/a08LCaQQTTj2Z4lBS83cJLUdVNvrF3K+dLfVQcw
SUUVlwdoQ/hc/L5wbiR8Bs4L0IEqP89JHkvzya02qf818zPBNjHyuREDashXhspp
cENb/NP7tU9k26xP9AOpwj+pVaa+VvvEMgP2HQ9pTTZzGPDCu3i8ftA5ZnrAFSR5
Y78xE29o8/uWs14Dwh2Rs2lX2FRRflZEYesCRQ0Wtoji+B1KriKcvD3p+X5kfzIz
gWl++hyf6DLbmJnyINmTTgx2f7uZuhhBrW0456XhepJ/IpdxOTzzfKX8/aQfmEZb
Q99leo4uxy7gF8F4aYDvcy22PIDhMpy64NY/tFquMsjc/RGqaNHCtng5F0nNR/8D
LVL/KgZUatVfkxqifYS8gcQWi4gQNrZC1+ZekZTGnQ4yWCitZVxbjxDHOe8K+M7R
zne1ExSgQbqneLK0AHIC/8583XWh//QdFf9SFs25eD6oGco3CipimegM4I7RKe58
O1Y6bYUri/7nX0/DIf+Rhrdg+pPNKICKH+T+x8XMWMLh7FK17XkqZiNNDySy4kAg
6sMmY/T0wzw6P3FBPn14FoiBHmliibXnVsteSt68gAYK0bUwEIZti8bwlSsU47e1
GAydlh2UPa13L4DcaM/7Y8ocfPu+2aMVhx/1FHxce8Kaew0vQ9AxaKZBna/6lzDu
T25ombxyuQAcY9co+mS71FlSEDaeh+VvMFJyTsrAeKor5mz52gV+Tf4h74zRNhXg
ZPOEDMUj/+xYmvMwxcXv9vCFzzjM9s+V9HfzgZNSCcYv+C2Q04aEIDjp/RNPKgen
EtsfbeQZ1qt55rzreUfdQbux2f/B2FVMHUrjAlzii3x3doFtFwdLSz8NcJhje36A
FIPQW50313M3fTbfDLuupJ/7m8/84g+7ouH6a1sO8CFErBvUDHQZFNFJVoPaFYWk
+ApvsOyHrlIw+EmB4R75pdDS1nQjZ5BpItRjUZOrFnTie2/Pu+XIq6J+hQU2x26d
PRPp9MqSd88adbEWMbzOFEeQGhGgFaUGBPyJbcDWHnRB7Dk4xkhb4DG52N9PKEQr
RqdnqgImauPvoWmk0CxD/hADfzchDpX6ogq5ykVEndKec4Q9pU+ARfUEBXZMlFmZ
SZesRJfFo6b4pWc5jh4faYG+U26v27fbmJMvPf6AGl+bSUNZu2ajkUqEhdMRok56
KoEF/zdPUM7h5fjHzsG6gE7+vPabJ5gemN+A0tKyVJbtn50BJ2C57Xlp/eY4i35n
GDlVXkKdcZ1TCLbadBhYVmhzkQLZHU/gsz2bPc/YZcnUtFKqsVnNS4r8OR6ZI2JZ
4IhFaKiJZAk7/IgEu01udiUKx79kUXKecjbySTzHsbybrB9mENlZb+wk5OmW7H/g
ZRpy4hAHgL4h5p2d9dlQjHSAeYGTbczcx3i3S/KrGVdQ/NrIqTzKPrn7Q/SrY2Dp
xfRck4CvJyQfAVXPO91sIkaB7ZYv6Z6+qVqa1hXk4Q5nvYbHGdgHiAoYvTgdlKjW
H0/OXYuQONNEDXDFYXH1HWhBuSpnXkqcLLne4DIneCtaUlS6zYEjc0gc1CePT677
hIkHowlU8E5HDwz+8dV40fpM7bcWFkGiKL+cP/u+MbKY+en5g3ZYRX/CrH5A7gyt
oJRGVnyjv/ksDtC/y+Y6jXHbs8FINlT6I5YmMGTEv380Pg6MSx7ZQZ5L9mDgGzlJ
2rZs9BYVLkkpyU6ma3KbgDaa9mGy6AUCLZCxqpGFQZZxPI8evE/JFIFEAdofHhbu
L0S1rAjMgUeVQVegmUCX8mik/uLhhAjlh21HPw37SyDJRlciS5n6EmoS3upxOvvs
J1TjzTReQqwH5y6U/diE/F7AZO0quV/8RWFHjKp7rLJ4K2n8aL9rkw/5cGrLPxr7
4JrshQ8ZSxF0mkoxUjk4yBXXJt42l1/fXJtvztyJNDfkQ0Rqr2cGmIQmLmdIX5z4
36rPXRi70+sBpc6Qk3FsNg2DajJfBpLj5zUoNuk7rHc0Tja+ZLEXM0vQfFw+PAla
cPxi/sc7qEs6AAbR6+fj+xdg96k+7qMpQPOTte3M75IZBZ19LgejWGk90ADyQIZf
x398+GhZ2lL+41DemqFpD4Q7rGaBOoHoUHHJsCMQnXFfxRfId4l5JCcD2sx6+xwM
gHZ8cxm4uiGfJBeJcKpPMf37RC2GHxzSK14dEDsekFYOHgmWGZv0uXBIwobuTSmg
PcMypaGnSYY1jIXbXkFsHNKX/GgXC9OLQxHZdoHU2Ii7Gk+cu/wtZ2R0JSelb0q8
XXA/HlOJFY1fJJwhaMXpmWXhdZaYHbbRPANbBzjyzEWoXruD4chjD28jQzcRtpGF
Mk4ZKKhWOUhBIfHqLq9q70BYRlZu3cA0Gw3ZKOuZjOA/Ew4MZmWMZ6GspJ+njIEY
oLnVbOCxTPSFn4wjxgIUijKzJamzgfJ+HqDgiobU9nR7hF0W1HE3WZkQ+vgAEA4U
PU9fmAuHu8TRg/2FqsL4tkxS7jOslcA5b3BGRHjDu+V/TEbjtP0ayOhQDMIGBjCT
BvMCb2eQ0Fuuep+khoZgFhgz/DNwmh3Nu7j4eNrsd1+yuIjzARyYw5hST9nPAD2/
ZjDghhP+9J5svV1A+Jsuu3W0/u1XBnyULgWJO/x79bgDPxjweTZl5IUjyOAm7iAd
uus61ZooG9Fd84VDPzdnlPAZEi0uUBBPRCawLSHKpraVOJk2aLMD4iNbcnceEY4h
b+ndzBse3nDJDCV8qdkMHZTPbJkv9l19mu5vtRYF8WsM46e1FhYuf12OOk5WsoIZ
vPy23W5bWMBrffKsuW5j1q3QLaihgjF2xET7wHG9Utm7i9ufaOwjgB9ETrtEs8g/
RN2xUdF+5VvMPOgbR9aM+uTeWg58hmB4t6pWl7Qo5yhOKHhlA7S8Ktep8rw5FqAG
YQYe1bXgpVHPCyqagp0rePVnPRnOuoJ2jJKT308do3JVQ14Yt2cU1USHPKBjDfVI
rU3kqAslpN+yO2dd3M4DyIZJv4XOrIZuZq/dtDiHmP+tI5bi6yAR2rIZUoLv68ug
Fg75kHuxFn+wnOITz9vq92tLRVu7Slm5NroYaE0NJ48OTeb/zHW8QULyyUMi+B+b
dJAXRchrn/lLMOjG8Ir65AoAEazYLjWFexqtRfEgpyTIRjDDX+SJ4bu9aqhwJtkA
6EozdYj+I6bVRSIu4/n1F8p4lA7nHbXTK15ZQxG7NrDrBaxVEIl9eOxjMXRV+lF3
ve6d7exKbvJH5z7/6ta+pRsmjlLtfg4KLVQHJlv0kqM2+nQ9MBQ+A6LQZxf+p06a
Z5Sp0BmQ/k8hUYVeqdmPpPje0SDMM+P4gJmfmGisQNPCVj1AMmZGRrKBuZulSNPH
BBjEWRr29rXL1YWcMh69vFyLTEVMdImS4pmc/DHZMXmZGBzZ0mXXrR1p/zEr0UW9
LeLi/19/vqvXGHdMY9kfvDZbDdNM5KhCuQlbFQC0a0mzxOvwwd0wLYh06HXCpUN8
xHM2OC9GEqB268oMUqzp0/Qe3qFek7qLemDuUL5qysSCUwd4ydL8T9LrKU7CNDxN
1HmPJBj5vHLqp9UK/LFSrpIQKccV17FPDWJLBmeyQD3+k3NPrbhCqzkCROXUHJLq
cB0vol86eS90AICqEGP99gXUAlemgYC9bDLRQOj4vCco//goLHPLuP7LdEJuUTmd
T8Wq7H7OgN1lUtlXkxt7PsZ9nsObIfRcs5uQRsoRCYuio80KhVzUWfQgf7FRdrlD
2fUNOV2m+heQ32JE9oIiM8S1xrSvZuIG3jYsz9oKFXalJBjonLOEQG1BPnruu2Wq
BCnxhWGpUPNlLlUupizv0sIbz7BtpVlcRDB+8O1YXUshkINrsEU9vL7e5krpy5p0
zXAqHqRCQInNkwe/I2arLfv3+pBUPL9n2qqGgi9RAG97lzEgdE9LU/jhLBl9CReR
CxCegVmfl+6WUNVYBnIIA5F5tQu1HIZ0puewJ7NkxHZ8KB5e5YiFHGlMwirwoLu/
EFwtXJVVH1j+G6E5NrMdEjGO8+9zoQGJSI2YJ3DNq1IPbtnl0FLbVBO414/sEo9A
vin4mevJcIP9eqtQlG89eEw0qv0vPFoUHjb3OAlzQav1C7wN8pqO502rBMsnggUp
S1Z86hugvDQQj4wKEAme41Ls8SYQxtSfr1VMi4HYlf33fbeVgzFXCkfhRyOiObpW
NRrwvk7e7V1UHF/shzaOjfBpdlWbESuyY+fZMGH/y1Ws7DwJnPKELC749tSxuWfS
qMe9L/n4SHGyUxTUe/f6p9oIw1gdmVEfn0nDhGSDBabqBFrxQTeD2Kc/SpTTPLKS
b0tbGbRVZFcCpb3BSJ/q+KC1F8R/er5b5QUd1CnN2pDEKROAwrVm6uwOPuFrdaCE
WTxKyw+SkC9lbFjWFIJ9lZ02wt9yr9DRcWC33vnX0ejvjXArSmBon4dU+tC2tLX5
QKdwuhkcruz4HLDOynPpv19iFerYTAqUW0N+Stu5FWXwCbwwRixlXsKfxyKvQlrq
mwvF6WB/L2lQ3Qj9T2Dnln2+bsUYudUl2Mx89kpBsulXVQ9rApKs+WqlELXW6pdY
1oDL/yvz6AQ5ww4Bs4i5kfBIO0uWtTcX/xZuTs1eYtTvFJGp0DHg+JDO6P7Jv6b7
2CRsSh5Rrt1LBri6LCSVP9nl/qYL3eJtK5GZc7x0pA67HJx35auVkgi+tQswW6Df
Jx4mWvqkw37/YCJLCZOGjMxHg5snLiQVRgOQ9PUX6BQeMHkaaLsylvWybqTiD14d
guL3NXVVcNpxzR0qZBEMtehISOs02Eh1PDMN5nq9JyBHRS6o1NEJAOP4PhidIW2o
42Tl+QNtHbRojw7nisDprpgnRbtP7+y2QGSOk7Gdt7oxLZJXc6h5obCF7PTUqzFW
6Zc1SVMO6RpoURWbSIHTivHhIhu6/52K00y5m6q6IlK+yM1w5kFaiW3i8k7FFRh8
Ueqa4hbUkKctfcEN1fhKDzLq5uYdd2oHOm0Fevw+9UIzUwsKhZvBH0GNBYFHaYGW
GbkUD6pkWlmCKtOyO8R/RUCXRXwwY33ciO8l0Mf5DoL5SRBhAH2NKC7zZJ9p3ovZ
iIW3qveg6hE7KWINHPBL4/NdAcr0yAeWMXBIu50dqJLbS4niaRio9+/cshwF+7Ej
b5700A3eufBnL8CeJbumpjZdd0JnzoDhlfqPy16rL6tsx0ZeDp6hDwwxMGnYQ79b
Yr/r7crO8zF5EnJgM0CrzieAAK0or1vfoOEhBdIUZrmYoOZA0CEGsSYt6y2PnQwx
wCIViKcN3c+yfGhAP1+uqBQzTzVrGJtIIMGMsMs6plXrYFB2s9Doycfzd19iyf7J
PJPkYJ+rmdd2fOFFlsYttF/d9h0IbdzAcBfOErJHaHvTo7jXHKc5I2D+SgjvWOj3
iVkWWVRmpiPs7gR384qH9LpbCy+BO9vY2g9N+rrtAYgY4C1zfKrROVTSrI3azkAi
kwS9nelLjw1DFrXoTDv5XUO6/4Q7z17hBqjvpnYx/9DERqOOFwjW+hEHpjnnEu2q
Bjq0q/P0yR9KMJGdeAhzSr7+GSUJ51b4WCItciwgkWGJGjXfhTpKdEk/pGvOQI7Q
Nn0bK5UrKYsH8SBQQfUcZrEGJTjsxYSq55Z44kZeppU4huwo/F1tUrwLfBa1LD3i
LWVvFw1RrXuUaqlRGzGL6rVL9nbJiWCln+I0XKdGmWLEH7v5eYACmVmG+4SfUfKL
bK6Tviny+ZVcHvK5/ttV3OV0vBhyxNglwnlg0DWtYjpinn1EGmgOm92jUDQfdkyl
aWMv+mdC8LAiDPBisbzBqf8UoY2yLCvYd3Ba3HXBFC1jC09NS8/DlloO610J9Cej
b5hv0lQ8HYh+SQ1W4z5aVS234gkzf59BAz77XxGUXRhAmHl3URF32aawHvrGlRx5
J9kl/aKiWULStenLgR1k+sLQw2FgWAEIY/afaYnnZ0HY2W6Yk9eY+NSQRLIrCpw1
h1JZGeYvX2HQ1V4TvhwxlEEYgHbZS9lI7/PADvyteQfHJJ1rT300E5OLv+elaWXQ
5fdvUMaqGu4tMcc4WEUH2la5k13kgN9W+2XZRbADZoSxy4a5JjBpNQCoDpN9Jjvq
IDPt7XxgR7JNFsKnUsJPHeTgsyLvLeGi9MuBY+l3P/NgCjEiwqDqAHhYbuLEWCMS
w00cFlcgsJcrA63uEwYRhb9ccEhYnyy8H8464pE2EX0GG+8NZt+ScE5IZE4qOEuM
kdzqdPi1b45iX/h10ELlfW0270NUqIxk6BLNNNB3m9cAhSHx75qQ8ewTNwrrSnyE
g1G3dZTnuz6fi0i3n/u7t8aUO7fJ40yZ883eikrhb9WqdsDVCkhkksaDFxBftAUq
phPvlct6h/4p4DqKzTvjE0Wznua8qXKGfnOhZNWf29h8373BDygIlmBpRhbH9IQR
yIcUOrktBxQGxN6KtO5nSGjW/Cl9BpPySknkDqZEAKGe9LvHqnoMrPyKUk+tdHJK
Qq7q/u1j8OgHDxbRPYGklh9ZZkKLIyE4RlTp64EF7+yUzImNs6lunwoUS0P5TgGN
sAaouzNsmXG/M97UjlFiPaJzsmzUoPOVDLdNM6I7mimjwlmoBtvgdx8lAFG4iH2c
AHRPxzaMFVYjpcJOCl47zbWLuGbfI1TPFegtDVyIV3gSStX796xthpdtD0rn64HC
pACAS85G4IrtlaXOl3AlkCMVp31l5zFKJ4Xv2suddrHDU33A+WkGSnW4NL88dI4t
GM2tek/kYrMyKC08YBIgHqF/RDAyQfpCZGNv6eVlrfGrWjt/ZsmTbt5x8ttHmtSy
/FHYLRE4zBNgyAOhBEwq49aj+D9kXCg/TjTMIwakioYjUHHCwn3SOc209818LUj1
OQ8Xdb2jkbH6qAtgrR3F7UQYgJYFS5SRUc9DYjOGZb3rR26dkA1YnbOXvBmvNzDb
ZOX+jG5dVsxIO4xpgMYjitENveBaNY/ZyOcXrmrFG6g67n2LZxnbHNHMhHxQupKX
+toFbnVwp6g/LfSfttET9mDjcddkrlwlw8FTyQwsxgar6Qg1NvBpdJWgdrfspA9l
V729qGXcuOnyG0wTm4hVNMqHTfdQWyqWGgZgEKbV73NfseGEiG171ZRNK9dEpuix
qjdvkWWQAzOLhxDdW6rkmluTsvraI1Bc+HxflBqWqWi4ywxEgM9XXMYKuCfBV4tg
p/tklA3oi7WrU9XCGp7lDTkdYK+mULfMQs/BWEqB0gEUMImjayruG1Erj8HrqPFw
hWEm4kg53bii04PYyP9pifU4nQf3LU4nOrmhfJ4kgMDtyxO/2UOzHPqG3ApLKE5g
OGMaPE0TpI8woHrWgxsjPFN8DkWY6vL4gXnTp7dr1XLyP+uhskKDAhYI3YD/ogfj
PnzO2Pk+uEpCJhBpApkH7RJPalpgQO/iRCNZXUdmcQ7pgPX3WI5J7955/WZl1S0M
r3ONyz9teSUIK6x1bOKnYshrJUi+d0fXKXJnj1VhuyGukKTrkHNLujpgJkkaS13G
Xtw5EPKjaMDJoQ+WHDs/z0y2g4ITEoCSN01KcjILEvo5VzYnjQVHBME6TKjzGY47
aRnh5Ti75AT462dV+nYGasH/p9PXtL/K3zUMYrFmPu9xdwPRmG7IfBYvk+J7ZiPx
z7vVAGuCJlurrCDdzCZaTLJ6aI9wXZKkcTYRJiMm9X+BH4JEdwhXxTN7zHD9fA2P
OdSuZH6+26hdxIlct2yFOoy9j6htlFZK2c35DHrDGoKK8iOzNoAbMjHVypLSAFn8
PBpsoZrpJlUWVG8F8DFTcbOtXUdq0Q5qX4SzTAijebd80ZPFiYnHIy9k1B0MuXh4
jhqBWFs/8CxWgLEBxOIKjue2Ovk1D4Wze8j8cLtt48nzLv5DBQRP55E7IMr/rV5v
cIS7KmV1bJw8hU4jNqcMScUaPLrVRi5ENQn9U6UdwR7nfa9sDRFr/sHIyO8rwhSZ
/fBriNw8QaLCYptj4uVvvOrW1vW4BKeMSfNtMO10ON42ke6WRWkQeEx6XDQ87Td8
nyaq2pdAl0hvltcbptKvmdj7D9d1UjU1R9SSZGPSqaFqoNrVRQBcWUTaF6w2F2Hv
d5Va2AohkrdpOgGRKAvfLBvRVj5MmLASuvt9mL/KxlBiS1/RtIKgdMfXrDfF+38e
H1rqGBlfHIGJLv3pEy97Hkhz1b4qBjayKwARNn5bg0rqf2DxBmRF5Yau4SCrmbOt
KIEtlmgyHyJEPV07+w7k11LqEKWz+1Aw5x5xXNRLtNPLxaTk21K3BgH6Sd2yt+dJ
VGb1nQkiESD6n533JLMxi+uFZzLdwZ7gszIg6HftuA+kepR3fZi+tPqyIOnRHBfX
b5dxGg2tmM3PUMM+5EjQJ0ZugEoJ9l4n6l5RpcQwr4aSaVsxjMKm0eLnRKhXU6GC
bmKodrVH34FpktRmJXKma9G2wvYXCpRA3RkJTMn7OAOn+Ft2YPX9l973J9DjQJ83
kw/NfVpm5blot1MePmW/8OflMmf3n+qPLpogDA957vKQp8V0S225eodVRZDjLKxg
1iozsNFuuoxoi66xtKuQQlYOLyujRAzznbtBliNenKOnnQg4+h1tkn5qhjFID90D
DE8yeO0PofFVioWwglua8OqkfC5OyJg8DStyOG/cDeVMD/nXWsZj0uCESXgbCDqQ
i/TheXaQsP4Hr+PEF7JqNCZYqGcElu4bgx6wnhOD5TLMcjNEPIoGnWRQXYColjP6
rS8DASsqcG0Gl3khx5xgzac/uM/V23bWh7mGbhEIXTsHr+RkfI7llTZQ0w2utJwp
by3z3xLTmy9Rb2b6DuIAnO/MJwLnuNYTSbX3meNReu5IjfmuyeAYqKIX94gLCXnP
LHH5ek49jDg/5EoAWqz9Is7lxz880y7ZBRdga98w87goiqrGUpmG1WY3eRM8viGn
lpIPMr+tKGpz2JfkrwbVYhD/ywBwbTRKF53HNmgCBMtJuOgY7AmB2FDWLIr0jpnK
0xso/hNgciQhCzpHsVTAbu6k8GZ+DsbfVJSAa1fS+EzbAugWWsBhWVttQQuHY3mL
4428OKZffbXIAjrcItG5/0zPmkFRB+pLj7ZTI2KKNULQRAGsKSMFsCZqmqLpjfR7
wm7t0LZrrABMeEP44SEKLoqPH442J2GIhLq0YnQgmHfAUcQ1L2FfE65tu8yyVhrm
HrjL2CfAlX27kwKCQFkcC4Lh31nAFL5E10bX2LmOQ95iwimeue1XjmbDNNgRub9y
+6cTYeRjpkTxOJNzTzCtjVqLw1qJCFee9UnAg+Cb+sbPSnnLhv4svpvcryhTBz7S
vIW9qxfCEdb35YnP+CMCiDVZXh/+1oeXCVbnnV94hyEljGdcdRJ3GT+Gty23EzbH
G9PqwsSbjg65JxPnFuLNzjBzavV7dKSnTpKPf/lj9FZBiUN20VgXHYY2RnxU7ePk
13GbXK/Vh7phOl/B7GuPBw5OirJP9HExxQRte0A4ToXnZc1sNlyxLR7qrKo3SKe6
XL7J9ul5gMNkn5Hoz9PHCvqYGllir3cuWlCj9AQGtogV5/Ht1uCe9uQrV0ZbNED3
QWFaHx+M0VbOITecYykSJSrBNRNvrL0Mbx66x7z/TKlVpc4V60XXcXBKtI9P3H7c
mR9ahxg1Zo+nm02yVY1cEw4/HAd1AULs/5mtAU/Yk5VshaxsT644Q3yWxkyLk+sU
M8paPeN330GOJwUUcmHJw1KBsu73cPfEBOM79MflHxYv34C6phv2IjOENNfnYR+f
2TOiDuHT5FHkMKWeLTlffwAQjg3mCsd02aJCMuJ7ocv0Lc0mckJhnMXzDVAzsbUo
sawoSNzYa1D2hTPScYG3K5yrHDO1Wvgqn2blEEaqBGYhhGXp+ICIpKu1L+ad4dJU
zurlGL9kbnf3SYgJINBWXlM+vyPnPS9Z+78eq6lVuDF3TsNas21fcKaSQ5/zPQje
vg03kMtAXgKhvCTW3yJ0eRzWAW0vDWtV/x4+GG4lR4BpOS0pyLY39OZz+QgtvvlL
Xg5zq7U8hJoK/z0BW76smsRqYWs3xVWw9t6QHVIDJ9gO7kFBAyRhh8/PAX4Tccfz
UC0FUV1YcjTIAp0fxHqsqVzTmgToVX21EyB0ls3+0n+jDsKD9t+cFJzGOaZuFKSq
ZVOf1R7qooct8TeC7jhnX2PPwgT9f8dAwBa3gh6CjMIWehhv4tocWBDBxWy1nVZ3
i2GkvfHfUYc0HCpOQtR7u6fFHoeZsQEBJxRg3D/ghZXvf0t087vvcvWMDonzvTCe
/O2Fy/4VvaaCI81k1W5xAVzFqHqpNT7u1sPNFrszgNLKAzKjiAKOQ4AKb0gy175i
EMlqH210nyQkazXnT/g+9qZdQXyulvUOO1me0/MjhUB9v5SfgPi41ugVFUquT3oT
z1DTN2zbFSWOXjsDLo/Iv8aWgrXlF/4bfeOuaRhIY/xs6OubLRyoFEiIAlwUwFkZ
YkMvwdpZH9ULBnQ5xIooB+BNgv77x4rg0rIgsMjUaiGbTmmAC2KKi6aq12XkBKUB
wsY9HWPmboqfCeyIGZJUjS3fITN8YmWDsDTj5T3IcZgQje1BNH5GlreAfKcsROxI
kfJ89FATV84aOiP1cDeVim9WwpXyYks312pHyYvvxaLOjdOHXYPq0/whCobNxOvF
HOaz3Q/Smac5kgWSOtWyhGCKmsMMwjMTg65RTQUtvrpCfveb/lgbhAWW8HLn/FTc
tdd0ppSy4YT5sBmxjOC0Vv8BjRiSb8LpMBFwnGtsgMDFLybl/hJAKbswa/ZOCxKe
MKDDOwUUs8fcJk5EwB0NPnOv9G+MkOGRYUofEJwzne7uMV6rEdLow98or1SoJbM1
XSZxBSl4BpLoLLxJpeCzVnEmuI7iyyWXFy9kvm4n/YuXzKek6yn5NDy3Fcwa9fby
2aWjGHOG+PXUbjh06GWoaax7Nq/ahNQjKVutJmcbxULScPbFtOBFefyVK/4JWpVg
ywZ/doCsqE2oqbWY06R8LMLyV4TEBADWVF1ROu8ajGpbhNScfDGYLHvpq2z8wER6
i7lBaAhCEzaZtPA89bUhPdQccT/EKUHANdGn0uhPtLEm1NQzznjv2uyQYHH/Avri
0HbJRmCylkAm5ARa/QOnEAWfgRupQwY2e8LED26xVNs31C/ZHSdDMu0faUmchD1f
aZ4q7V6FqOt/oT8LRZSmBaJdPj3RtQID7xnyJXP4dZmIuUdwTQd9DVCiNPZyfx4g
/TJC2vwWHl7cZbq347IjPniwQcAfvWswJt+EGcGIpZNOkoolWfts0Wvylob7xyJo
H6wo8WOCCU3v5od7dwhDEfZttqbOwjCUmCCFQd6YixVyR9r1A/YqmIumTblsCg+c
b8FqHrN7XsbKGqx83nDkiQ5nQQg1NNLjMdAUPnbefTb9Z1wc3Zfa6VoXwkoxUAOS
r6ZmdBzBiUoklfD+hALu5c3a8YufWVE8dmzkTrOV9fdUfAihikze7hS56JAZHu0q
AdaFISi5qMSvTMWQtHM5maJrRMAePc+VFxBINeveZfqZte8hrjrwTSPQDrJO1Ypg
SwOkDpLH36cNc7yh1a+8izlYuudTb8QGjcEqEh9zzvsqQuFAWYPSg3VDPwCde17k
EVUWv5abIcWTlE+hoC/tRsdNGRIWjjvr+3FgyyKUA0XbzaFQcJfss16vVX2BfsmL
IYtCrknGiNfB1JwUp0a1XcFg9TqxlbawISZkMbcBBwMPtfkdhaz/08pfoRwCYKIc
GivMqCbYSmQEs3yrm2VLPPe7vseCrm03n/G9ym68ah0XYhkd+fs6fsS9daDWoQCK
Ale82oR+rJ7xnlbJPYanYd7TQQQbgAspCHNJDo2iIoBqUz4mZuPDW5qWgow+ZJd4
SIMwsPJBqtiMa5zM9R6Zfmj/wdraGszgMpEd3e7afq1NZ9DcwkhORcKdmvxu9ZJy
gu8vdRNWuDDEgc+rICmhPesZD9Keyxuq57YMgHiYHxfJFYPEOcPXmB3BT8wc1M53
pTF4T3+MxN6HKxaT9qMrVSPI8QnTAaIcH/dn62JqxxqYsYtTI5MZgUjbgllZv9DA
2WfXmIKmIAynHJkI6JS6PWXc4bOcB0jL7ZeNWOHV+XqKy6FDNrL1ez6Jn3u2iQST
o7+rO3s7kCKgbLkjZ9vNPyzfug+gTfQv950NfFSLq0vzq2B933bxkRJpIMSvQ/V0
ouyNim26jHtc71ZQjJvEccbKeULjAIe8Dx+bQS0hImocYL0VBEccGo1X+57o5YyF
cmQcZHPRebAiD+6jlZLJzCdRIYZKQnJYjpTlqXGGjv3xh/qa1EbV1fIkHvcUQi7F
o4CRYj9j1hycofVvKS1WjRXHLPU9wuN9X0QrnQfsGggvD2/nuv/X6fFG4XLxptR6
mzu2mIMkuT1D/a3Higi6AvVVuZY7dr42XTswwKV90g8Ae9EC5bH2xpTYqKp0xM8X
OgoHtASiM2WUUiuph4LvZvCETuaCyNDO0GLM2DIXad61YnzYBayRWeq5fR6645ut
BP8zq6DIDpONqqQkSXuKYfaNzLl2ttTm7tS9yfYa7T4nCkxVRCe+3J33RY+xXxzz
ZXHqcVaXGTB2NEDtcsyXDEicpi0mtIg0DCSVTEcQIX5bGx+mZz77et81Y/c2Hkz6
pDYNjgsqHboACNo8ucJgllif5vjqma0QFGwA9SXBR+EdS3BdmUvvGvVjvDmul+Kr
zf52Hs143mWcwkKQmwpH/PHRwDtxfgZv4qAb1vlimmyNMqYZjPyr73T0gUffS8j7
aGK07xMqKed43N+7UTil5egFyABOdWG2Qwm0HGfbZh0WzFobDblBdFgCPMLV+Oip
po6yVaTguNUHL3zFMdmDllsKJKsu/rw2Ae2zGtZk+CQgzuECUYMgotWoNbOwHb3f
qUkmb+m8eVesv7Ch2JbuvdfELKCvxhCJL6izrWKoN3eisD6eUzbvSLTSzHgVNFOK
5T8fKZhUg/NsIxXpZIl64ogEf1SRxfuyH1uj2SAyuN6VJ1znT9X58PAuxjFFuqKc
qawpyZ8qO3Me5grR3V2/W6c38l+1/7MVBsDKMHP4cECLWt8bZrJDCnNv/yvmrT/Z
JXU0B1iM6Kf9SkuCG+7hniupENsHLg0j52aHA/TZy4DlHPDKkW1jGGsgmhvozZFm
9p+RkxwpoWlBaXhEzBrPuXX7vQ8AhFw3h/DGaiT2lJa6P3zWqrN79fTtWAmIymWS
CBextmb9Yah1TfyglaHdBS8tNxiciQDxusViRE/Nu1PNLhhZFZsG30/giE08FYPw
+HvfYWpb0FFPyWvI1jTO45ISkOMQnmAJYeVZ9Sc8KO0AEhaTVI2Y55xz7Il791v0
NO3AdQzY2+BH4V+JuUNBql+S7QgEDGIP/zcYa/FkhY8TzIKL84ofSV5C7HdQhIiT
US9+N1KcM3eHIXQznJQkIKxiJedxvw06EhBvMasUmPCOSmEm/F35TxAQ0X/PNqKv
QQ0MCUQMK5cm1rv1U0UrK4PnvpTDm6zOheBGKkJ7UrocsYiO2uCOtawPYC77rBhl
xSCPmH2csHzallCF8bcTZY0YPC1XqYuHVEU4sG7bbtgiJVhJn7U0TckVXKOA85eb
G5TWLAh4TZtbCf8ZTTpzycy8mwL08zfnE+ovxLFqjbYDKsX0ARSExE2hfSsagxU0
Euyftuoz1aHJIWLc+UM3exA1VyE89JOFUAc6W9giAc1Q9oKcJtZ3rZPqBm0Hvt5z
mdIXTkQwDbWZ/Wew5WdKhX4xKDGKhJGbZA/ev6LgAZDLQgZt0JDM8OoYqP+54h0n
663LP/F7D6jNTlqA5x24qxnwMutdkToqcoYcvxY1w2YzOJ5yUqT5fZyG4I/4qcTN
1nVuszecQXAtgBraPCJSWd7AigxS4wgbyxh1kUmjY1xJ4XmG8qWMDpuIXvMgI16L
nOGKPRHT0fNJhUBzHNl22kftvD97STSAraqzzkfkcNzZwWttR5i6lWmCKrQOE1M0
sr+xZq0ncHkeNaGTGS03OncXN98REwJXtbhyiUsgvBAwC9+MsL6yrDdPvR8Forrh
U99HaOn/5/5BIMdo4rTWjemfB7PEbsbuBokOYNpa1HaZCNDg26nfw5DOfGs5LsBl
/lmzqexjgJFjvV2S6/ApIvBHjMXwyFKoqMoo9FgZ4IgJGfsvPcddkAKHcW8lHFu5
+6mAz6i1Qscw3OTXDMLvVGGWBfXQY1899vvnzoRvPiVuVdTKVH4XBvD3yDcwzY5p
nge+R9U8fUvqtCqPj0hd4/dq9TdDzz18IZOZbdWtCNWn5bkpdLKNoDEw18HzLI+i
akbhG8h7y8kBuCFr189K6AP6e8XWv1QVbpzHm33wX4o8PXTtirhQzrIFTC16LTGR
CbD0lws6nVsSdogLxjXHKVwNIIXsatYYvPVEXl47TBHSKAfTdYB6B2/JxlACQEYu
mZYEyjwCP4TISBqPljKPI1qGQSf3ugD+3qzzWO6v8p0YtSWnNJP2km7rmMjTukJi
+6nJvqLEd6Q0sigRtPS0eZUmKBA9SVOPzhy/XOr92Tq7YFTE6qlND12uHUrlCBHZ
ZpxjJLkdqEiRkwIb0J/xycqg4r/ChU3Ajm/DbTICZWR0Sn0F0hGGYBGx4SbKDXHr
tjMv1WpCmv7qKt3cXD9XoCr+vmZw4pxYMAop7f5TS/IIF8A+SrXvlp3mQLO5zUAd
SK3+VQBQ1CXK13wlPuwRA1g2le2VoV2hWcrCIWd7ij8tvIccaGDdVDSl4iOhnWOn
X1ezSWqXlJKXQa2tSITx3oY36wwyeF70AlinfT0PEvoyV7NT2OqkpI/BVYQqBv6g
eojuFc8hh1x6l9jSGt2fwEZahuUcZhDtjOzwbPi2LLV03nb+9hipw4lepFzu8nSi
DS1YA6mS5MD+HCA9rbVeIIBJ8wZylLSkfljJxecLp/bUopwHdLeGRJ3o2fLIDlbW
kWZmx+69BQTXOL7aO0YTwtyq9a+wn4bU5GGf5rjeC0MFvUL2BLDJHA664lWaQYLJ
+302NL0H9Og9m+F0HeyEZOpWGGZpZubTClgyJgGrHNxYs0GAf5KG6zVGM61Fbb+j
+UD/agq7dUs7SG6y+AL96IHdfSJ+BbemTItUcCnLSl75ts0MuOYUyFnwpLWQgtzx
81TcC3Lpedv2HFeM4joLl9aeUK+j7uicbKcwVNmZpghURFR0Bbf1nRa/HiYt8tpG
Q7SdiUuJC/AGi9i9LY4KTx2YMtX/PVltsxjDb1RM4lYyd7ciM2y5xvnHIzacJvPq
cx/ehGVl6YwMVsq66N7fPd4rpwcdVYygOVWtV7ohx9N/TLNWaV1/k/lq4f2/6H+A
59i55XO9Sr5Mb4n3/cH6gvwiImvVAfFKDaNtbVVRArtY4gUah+55t2hrf/8/9YGd
Je4LZ0Qe4Tw5o0cuM+3nw+1AaBrY/eXe0W8s8HmnCV+WTOqEGoOqBQLoJXA3nNqP
En/I9eqEa4ZumUF7jI8eDQ+Ur28VdBmnsvyiuG179UVpjSz5USWHBIejRiHBzAc0
htx9i1KO2N5hq5CRW78H7tkpYp+OGT0YkTcGZ0/n0ldtSFMJgE1/VQsPHqG3JMe6
7DY+FuWW4gVINfS0t+GaZtin2iWU87mMyWxv5H0MJUGUZa/joC0aG9cTQK9x6P1U
7/+NCXES6+Gy+ajc1AexAcMMSX4Yjg3W0z75eoWRKXpiyFcK8K+SCNvvC2HsXiMF
f7D+cBBKOpuy4IruZkdnRiF/BkhS+lfiV9E4xbx6StQfTKFPeF9LT8Qr3qn3n/sj
LlSSyGiAWNUxEo/WqFcTPVuAJVzFOUEvEfuJR4LFKpMG59tJKMBKeFpKQhq/M809
oHo59uZFmbF1H03BhB0NeJVqMe9tYaPl+fZ6q+SBg8on4S1VIhRqX80VXua+PJsh
xpionCr8fRIvMCogrcq6OqDnAAhbunc4S5c4prZfktFEgGACjJ5DQYi6s6r2JYxs
wosSfo7C8xBJzZwvgJAkNcPDAJP6kmki3sW++GD1HfxpEEy4PjDuk1rVLcknco2c
8633zJ5aCrTHSt9AbXRel0NiB7RE6RP5SftZj7fkS0qblZEKpILWEABVihNlC7oN
x2dl/1+N9swDlN2Ml8HnI8GCS0OQWWg0tkXbYhNNR5VK04g4Y2aZNa0dty0Oia6t
frggmq+9jgT3oPKGUBDXQznYFNNoRxq2MG6nAMaDl0hzYH6pwn9yu67260AkSVvl
7aSlpFEr24H0w+VnHpU+hYo0diY3CZrYT7u0NffiFgHtwJHITSvdKOSb/aoAj3fa
4k6iumNQ94PdtQvLfWJOjg3s28wn2dQaq7HlDimaybxIF2aIeBfvAz7PkTDOaKD3
4K8z4wCwy7Cbfnikkms0c03mlzEvPISMesFcFYKUGLpDFGxrIwqfqdRSByjhGcAy
ZpFws8pmIZGm6J0l59RbMflTQE9vDpSsKO6b1j51mQChPP6/BpRl1Up1D8SvjFNF
k9AGn2yDM1L7yNH5YIJbKqMH+cs22lTiBzNbo2G7vpdEabN89QQXXGhg+NoMQBRx
eJt6Fo1PUMG+uWMlJgbyM4eBHmm5KAm6ksqZ/t4zMxa5+WlhPrW2Ub7oW+D/Icum
yAOK5y8dWqTv3eVLn5/8zRto5NfCLlyvtXyaTQvos30m9YqgqwBhEXi06N5m9SOD
qStvNTehxm0s6DqDsbKXIp69ZfuDTD7aP67MhZCkJvbqErzZnbefi7Mxozi3uRCv
TdBLaMUIZGfsYAzaSibISpkH/9SQe1/0BT6/jkbFPcOPs8TudVBbFBBYpg+dvuVr
iaUWQhV9gWph9pUhcueeymOPkGLy114NZVlUYKZApxoGaUNq1nMx5VO9Ms6/S4PH
hC9Sveyd+3nV/OwR3dzu9xXq78R8YEpftXkCRSJisHfIJKaxSckThPZABJUkUcmC
kuXanak4Qg30aKTMq3BORWWzKU8xGvGRXoiVbsqW0SP2sHjJwYhQCznXLJt5qQtB
aNsecq9uGYP5+mKZ2RX4K2vWL9IWJ+AxcvlJq2+4QGCa04bNc32x/Zvx8sJ1htfY
xZ+7tzd7w3PrMzFrc+W8545/Sv3XesoyEsjdtTf8l+SdYG0drEBJMLgtQaXmV42v
fCLbpZyxr3FAKutMGV6wsUmfo3Gq1SoT2V4+I9rr/2xTieMHrSgXj9X3HIn6Fkp/
vJnLq0rFKsOgmEXBamXkAQwL5gZrrOxv9rxtnhZqDmUkmJ6J1e/4nfjFxtV6UOfZ
JPoZdMQyYCaKbgzHxAJ67mQRUVaNaqadY5Ek4DOBOKhYXEF8nWfhqqP/eJkkKjyz
Sm2KKqrJ+9YkfnVVSEd6taOdVmDh/Z3HJ2301VOYp4xcl2cSTukEqoA9njGUxGql
`pragma protect end_protected   
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
mTJwxRJXoBOi+AnaklJ3Hawh1859D3VcpTzSQGsNqVQGp/Ny+x769srPx6XkVajx
rrl9WrBZseQPeS01viCWd8TVv5edFmufdztXz4xJPPoNUMEjtYxnHJZwZC5Qkt2a
cNCgDYbbnxF4jatfFbN0jMkhEJmg2oSy+CEsxUla5q0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 454313    )
uMzReaArNMrPuGbXdy+K9vx5GDXPoB7Ppot568NWcgSHq7LU8iqIZm5f72H0s4Pp
D1B+ksm700YgVvvJ1bmdCFbhA+nSsn3pqJdoDtcFS0vf2TgrL28qRt+BKaw9D3lj
UFR9YU/yvVwdddoGAL4FLvHIjhtsV+yIaXJ/T6MLzxQcsVctQrLpTDp8QSh/DXoH
A/00fgYLkLRcCkIz+CwxZCOp0L4QZqozklqM326EdEn69fLmlee2caGH1n7JaoxI
`pragma protect end_protected
//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
pdPygj8Nh63Kno12e+WJdaae8S02E454v5wnhtVC4EyrgpHZytx7nbWFwV9Zlw8j
cp8kjnB1Ac0uIoUP606Kj2++uVmBDG6iZq664RvoLNbYlWn1XSETwOV/R4iCtvul
zmivtunOBxpWH+qkqkdj1F0fpKrANah8/uSMnz+YL2Q=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 520833    )
MHYveC5NUg0QCB+ZwaoqAr0Fo0DrLdvusADDbDTaorasSX2J5Bixn9v4owYO1exD
xill31VK6vXjIMs63ohxion8Bgvy72X/2WoIUIcSGjHYd4gCPEoa3QQyh2gaDW9n
G0DYnsovU9eoua8kf1CbQLwMyYn1wgPRVm/NvVIKXzRh7eiTkEZMJOeZs8q7SLLx
7DH6hTd9TR28Qzf+Ur3pAN1bhQ1MuWwmYPFPbNG9i/qdcAuytPa731p4/wzrt63B
7tpEqnoH1CDG4NF/zO+kbRrC+GSLhELNzFqITrjW5+0FppMXy4ncMpkb1rp/z+7b
tUp1heUTUCqeYpbhumpmtquGPDb6idYiUKoMwECFWf/NkF6BorYY0Tn3C11BdO+N
qckueMQnaFBgsjuBc7vgoP5vSj7mXyO3nszcI8nFA5gSJb7WTGDYOi93496pupBe
l3+/d7pCtpOUwdJXBet1AZSF5ldXRJNUxumOVG4UIw6ZDs57Yo/Z456xQ7qxgsJN
dKfF47Ls6mOR1dOpIOqgamNAuGTFHzxTs3VVryRo5wYlTZ+V2JaNktz+KG6Kgn+j
ApZ1oLZyzg7yDD30G5FbsPhvwgFXyLAoFX3v6FjL59qamnzV3rzxBRvXXdXnsOEQ
Ra/0KfBTJihfBHv5usY4d0WfbDJlOiBbl/kgz7/POrC7DqachH2RXrubvHE9imPi
HP80MmReAQIeL1nv9aT1+l34C2BkSyj53Zk3f/Ziq2MMzPoZfJXcIID0xnow56Cn
lUtN0w8RUAkNLl873oO0J2gztZw1Y6RP0Q3UaHliyzjLOkWwoFstHFPJgl8syMmA
Bs+51EYZlRbAgI8LqhV44iittCzpXB4idSRAqx6DlOPYsfgSJ9L7cfa56Hsa56qQ
4EEBmrJRkzgRuCBuUZsPppYGo+LQlUV/J/Nj4wNxG7WAbuYAVNXIBBwLl4tIHGhM
E1m93Cz2CPcL4S+r1II9gDpGqh8/89yq0JiltDmeE984MYyjjfrNgnDBkkmYjC/3
/5XMGvk+bcog0ErEPeBnogQou4H4nMvqy0zk91q6na9caPQ5h0Nf0UvR8h1NisLm
RiLHGfGPDoUgr/WtjT8uHtEsM5ceQdBEOHV3wABu3Ygy1qbkGKQCzOXuHDLjn9O2
oq3k6gFisUNP5FZBsTkLDKMScjj1RnZnYNjVsDcYUj/T+H6NvmhBdCFW4EKOpy7w
2hhZ7hUixxSKyG0EledWRM0wiujHq3VLTScXlYZcxBA3Liz+Ge5vIm9QACVBAc8j
lO/YNDci9jqkJBF/Ri7/NknKKx2tkENcye2JZpIscMkhDxXJF/k68iNM9a7Wf10d
+RLeN5GkU4Hj/l2b3O7VcVsGxTeCW4wZZXikMx2SY1zd6xpnUFxzAlchSh66RxLN
PHZXGEolIAape0SsDXjDr3KrTnnaQ9uVGx0xiB3qOpuzh0xF3A8svZXzZH2QD+/J
FQaaYbjuJ08KfVl0betOMC0t7SNlXEaN5W7OncpYszxuVb/0yDxRHcy5i/7s9gbq
jFI0Ia2BB+th7JuLzxeSuqL/XfO8HQeobvM7hm93+Gk1dmLq1zrMcAevk9/tYgDM
VRrDw6MWjUiYZZiLjvuNgR9Q6SKJZ8fDh9JTThCHf5Rgfu+T2DEJu0vxipNjAH/l
rFtdR+6VjhR2PSKWzCoA5Zwbm12hWgMHXXuBsnODRNsQeShhKqiEWdw0w2BbWL2G
PCsA4fnVDtEn2SiFyMa3gcIzX7vvbnoTxVnMm7x/XG6NZTWjO/80A2qYMRjmVknr
gocWJ9fmP9De5EBbPf8GEMJ+f3k7qn7DBlQUuEk1Yb0F5I0g9rSgUEnb/EuUN/ti
aq4wZ0Ta3G6l1OCKyGHt0vuKx8K3icRcpfG+Kqra4PiuQe14Tqg+nwEfyGYZalKQ
s9YZvfs4/4CT4ziXecTCbKhorHwFYTQNly3rKcxC/eLzY2AggMkFC8dupOFUr28u
B8+Vn99N4//K3gRfG8mC5QlnKnrKjbNX1q/zLDqfh/enMnsh0zTm8ixQUvy6t4qs
e3isjsOXZgDY+FwC8FFprgG05EqmcBTwa27DVCpK6DiS5MK4JrWrBYIuLukUQTYT
kikWx2uHDwbPA9n2nAV9yoOEPzltCEbIHMRfZQn7FbI9Ma3C6fpH1u1ul4zLg/4t
1RdWVXWTDCoHUjpM0hv/oQiUrsN2jIHDeSqvi/QeiRDTfDXKl8iSQo4O3NyflGqs
5q1LRpSIQqO1fSiJhF98TufbiZlngPVWk7ACNtJtm+Dq2+ZMiJKiyHahHN+tzs16
kiMmXmleCob9FRir2ex9SbXa7Ge/BiQItlfDsFUuhXk3snCSkuPRJZgGXx3xNH7Q
CHWTNqfdFMl11zXo3xjDGFcyG9mE3nmzwHuZagmGcoSOBi/Um8Vn+qmo+Z4ZkjKk
DL1oGUK+n3ZMWl2KUnXQL3nVuNkOKUw0HL4oIP4NSRnma2bPMadKbpyTiSzuw8Rc
QC1x2Yl2vd72ovXSguzhSLELr9MLdQaUm3tJLbBEGAYlht6Y1AdDKvkjX0H+zXae
xehIciAjBG9SOBJoWsKhxu09+XrPsXeZVfwBUsH44spUiw0+DMeDogDlFfP9UNr/
DYtBoHzhPH8J0WCHZs4JKORPlj0/gefQM/pJHiP3Vd6/SjLRBbkB08EI6irBDUNt
BzM4r6i0i34h3WK/gjfEJKN/BJd71yc9b+gzKQ3P6AyIgN54aGle6sXi7oce45yW
Nl+Md8KG3t5oeS20U2fHvZugWM/wTlyLQnPcQ3xtpFnXQ4Yz7U/2mU2kQQKTrJ4O
dGqecysOEMp5R/+goljVinfI+47ZptQ0BUaZkz2H7lHNrzYHJBImTNP//5uVh3kK
LnGFxG7gjJFVWOnnSm4AD1lXXHjw+L6jvkZEiwtUNbowYDnuq131Upa5wD+0qhm9
166yuoiaqXvnrlz2Nq9G++1xWTYRZ5/CLBNlGF7YZakqA46SNd1GE5sQEuXwD0ao
ASZmHk+tr+0h15V4mzCHS3wgYOX+b4sWriAUv+V+io9UhGPx6GKRuUS1tM8Q5rEo
Orkajpwt+Tmzfg0bfJ5JJY4BKacKk9DxzH142jT9cZYYb/jPiFwMosNhVj2F1G67
Ax0ppPI/9noWLJzdRal9k5uUNOB8ECy7RyWJckFaBN3SXbFeBPaOu4u4FUVc4OBN
kdl7q3MYxVMP5+uCAGo7A1UePIRL2j1C68NIVxOEZsFKbEn1W6J5Nm5xfr4Bafes
tJ++7PoyHqC34qCNisQHr/54rVbASNLKKPdf4LjCPu93aPp75EaKK+Dsb3zbPIOO
uEjBW6HKDhQcmmV3JjQufN5xj0sS3fdS4tIeSmP1VYUYBH26bQguArCbxk8jIWgb
X0SNmsbcGNeM41XguerIZIJ9Sau1fA8+cdSNOiR+H0oxZ0vrSEczxfH5PFs7F1G1
/ypPcrIE6v9XV2L02X8Ct4E0fjd8GiGwK7SFjI89vC6C+l7Fr+1iK7dcE0Yu84Ng
F4xszWmwYUxlG3N3IHLNssJ6QjJe3Dxj+WjmgA7rxaHNFf9ey7uWaNKBsVRLSIgT
z3EQ7eo3quuphyvcLcTQ6dC0R8aV5LXwBMd1mPJWW5UGInvl1qhap7wh0G/NnaPv
rmOocx/KHSwF3qGFa1atWElpskuv6BsRkt0yOCitodLwpdEUVubTvcD3Ji7I+qtg
/qYjMwfXNAMQQJvCGIql8e128LHSaORgI+qXdFoUy1YgAGIXrYXOlBtoUJ66c73c
xw4sf00yfLv81Y+8CZRRIL/6V2tOaluBlKSfVdRBHlLWWy6IYDRo080Ue4CZ7iGE
uDObW8DIaqW85/Jh0A7erDJ7dJt9Q1+Y40OAesEWHOInk6CLBMFfqz4qjBXt/HhT
DNkJgWrJBLfk/m00CAinAv1HZcZubWWlsSat9JEypHDPHSW5SIpPqzdi8OeJNh0B
wHk6So1H9OLTn34ysMEeTSa+riNVMqpDx8Y7fnpnQ3+4BN8SOQXEIrGUymaBtRK1
YKx0kR3bbnq0xw5ObvHIAn1W8aaAyl4S3Tb/jcLASCrIcuCA7JvZIAKuMKObZAhv
5rZFElmmnPuz3Huc6o0B/TInGx23P56HTkXY41iD69io5XB3/aidGlLugDqy/irK
u2mio0Vi4dPIlbjxlasFRZ5OSYj5A1nA/D+aJRD+wRBUUMgTTYwt2WylU9dpee1A
JgNJmr3weSDiphmAm/jjnj+AhJtGVVWXESm43a8gp06kLzQmUhltHRftwJQ9sp4e
lUMu8YNBmLCv6iBn+D3hweOA7iIPP+4VEOD339r09mHhsOpy5FJjZYEcQLheGozQ
wfJbRnBD6Lxk1kz/8EozaQ8H3HGrpJCZZ6+9TyQtDlH9VneOeLcvQ7tdJ3RWde4b
6WR+1lkg1D0sqNPI5GDiJk6BulYV7Xp2JAjMyQG0ilC6KNoZcqGd1dPrN8tqRLfQ
SIUomBdGh+2bWobNjrerBLAwtmPpCWvo6qXhumO664bpZ8DuWgPCph9zG+3/6fRJ
g4Jx2VkYJ9XNf+JtGSHtfZ6AulmcUvY9EDvU+dw46+liLKcHdTddSrFCohQaf1xl
NYB5B7C+2/YjLuRuUXFrpBwEdR9KMvHzcPAP9QE4NRilf7aFGF0Z5K1lNp2nweDp
vXJWgy8YXV8UeR4nh2RCC0EtNg6eL0ssIuwKySxw6dTmCdvhLO1cS1SxD5jMgknn
Z7uPIuWCdCvlfNTZJGT4adrW+kLJyCvP8YPyEXOtk2/D6uHy8mNHs+ozDNIRuNvD
Weu8vWKxLLJUhiHmX/NvjW3C8Ry4yCmj7Nqy6u5BR19BNY6uXxz4f8v2T7wZSNjC
DNAyC8Oe57eP/nqV6nRvbPbC0y2K6V2eGwfpmCB2dE2JV76DMWnWyCi8BdoQ/Ll5
Tw7Oa+LaMfpLj1M3wjnC+L9njypsxebXJ7b8Qs3n/EQBag/sj+zgTOoLL+mCI6U9
JEk7e4IJmd3V31HFTk3+fuHHgpG7XfSzIaIuMdIs/pnvv56IcldPQ5hi1TPUBlha
xHnj7Ck+V04L8f/zkZ08gr8DJDVLOw8PZr356k11oT27NSgXwy+jPiVDyllpmLIZ
4golbLuI0wOvZbUk21BDH14GTOPBbfEtf/pYfs0EVSqlK6BHzHOqXiM95bktiAuy
0SgzujliGyybX/Jg2c1jczgFAMxhRCYscqbf+cyKVK9ufaD3Bg4vttsYvkPdBDCf
4IexF/lUwagK5aZcFVkVnbZaMYW7HWNvagVq9sFlJJH7ZpBS389QwJu7G7ioWzGa
DMSHs4Pnfi0/hNhlyDIVB/c98pfRJJot5qPQP3EvoCatVbo592gnwNy3ZumcP4S3
nq6+x7nd7DMB6g0foYIXxMmNmaOxVE6opCMYnHKcvSRZfe6LQgMHZ0LczIPzMOO/
3+pUbXFy0xLP4g0ZrxOAheRI0CcIJ0w6YRghDadoMpwOeCr/7t2cPbZTxR+6Cvbm
O08ajZ8fqkSoAEari7K//BnbsEpzf3paYHz2G9qg/jei/+FjFBkkLrM/r6Wb9QF0
fWFg+r5MbGqhnTssvDuDsuoM0jkvhwGDGuOYGlWSP9303b/AR8pfzCybnS2N1/sJ
RJ885LYOs6Ff+PlDb/ZhP1i1VFisBsE4GUO8MVlG9vgqZk64EM6+LGgdEAEiZRJv
3yZ66XX4n5sZbpUB7MjHMQUfyv52PYH922/pJe7zyr99KsHCYWea77qSOVwO9XdF
Gsuk2Y8zwRjIfAW3ezMwL/FjXbpwoz5HrBdRwZPRPNnidVouS4JJXZewIZ+QnBy9
UVC+gb0czk+N2BK3Vau9QrL+EBxLBZrnSXtP6XsE+SmYmMzL0+Injp15HxdOBlWS
/CF2EXnLbfflereg+dhoZHe0XWLqZMbFmq12s14X4JhEC5Sa3KsmtKPd/3pc0ZIn
IEK+Lum8RA+igaMH7PerBlgEozLBqNXdpWQmFEwNSYZ2Ov3IsjqJ1ApcTgU+Z+fE
vNKk1a7XvoQQhOpEZ6HBj3Ob6hrPfNG4A5Tj4Li82KDxPBey0bWEWxTzy3HOKkoA
woWkfLlKPvEd4hco406bMZaUif38eD1eMfl6nKAUpw8mdLpekpY9C/TSO0yhWUIj
Kqqc43NymgkiOvOWXS85Z38EzlzoFK/QesyprAWGM1b3Guv8boLxMsncZ4vHxZYI
bPXZl8Wi+MzOS4tvf0l35EKAm/3il01KZRj5mTuOEn5qOk2kKsG5ltoYFYaCkplI
dfYUC9olG7WKmoBL70f9E3A28SoNdknqp0Z5ijEX53zj+TSXl+GYLXFmO6PHP8Wz
jkmJ6UVnhpu0Mrv+KMbLRKgOsSbnjkbP8zNQHXhgIkFl3Y6PFPldXibsf43dGo7X
Wqitaw1nvBD4Y2Zb9g0rNpKT+sR7GIfQZoxFjRF8SCCaeD/QvEcTAPE/C2adH+zp
qXd2xRxc2dNC5FYQUOvmnkDsh5vDcNTo7tLRMQF4DSNFN/txp3Cyvjwsbgeiq/oT
Snlik8PQH3xb3xT8UFBmj4pBR1CjbQnk+eY5Lwvbw3hUxpHpkY8FFmoEBdZM+sbg
oKVfr2tzn4WYAf9DqJc7TIlQG1R6o9DNJ3/irOUObdzxjbbWdQ4mIIueLk80Qotp
5bVKFemCQOmTR9LdI/avlnnbEJyrQ4iSCeLNS4vvR8SaZVl76xjGEXOiuuH03+b5
hmy0rMwKqs9b4x4M/B6nhfyl3D/DfbS48FmzqboiTgJexgc9qO6u+7/U4dMYmeON
dfaez0BEe/RrPdHvL06vUYZWH25syLZrMqXCZayJiwK81VExphGRY7fLeaK0NEBq
/yjgnHWwIrm/dkM7Atc3fuRxYerhgEDWfpHgKq2A1LWRUyOAGOghB0ZXcOPYNJc0
FAkSfSG2bD4vIxwIK7T7BXmoe2pqGU2cRiQGKvQlnukmJXFrVB47XQzawFNlH6y3
e8PCzTL7+Osohfw+Omktj5yG62y29YUWMwAGtQ6Q6Fq2eiDN+4G/+rpCHnVgcY9z
BtaQ8quv+WdKpTkn4JhOeoZ70xC2JYh5kYCQ5ySxKS4dCmtMmfbMMrc/+LxzMEcV
G/cQHF4SFqdsLK1V4+r7IRVnHaBg4iABnwbsiONxFkS9DEGUNAz7DMVGQu8EnUTk
Zlgx208P+olh8YuZ2V88K0MO7tcyrrJGEdXl6+XU5xssG8Q4IEwswny1zWcMMjcO
Df2iW9tiDvb9vH51dI7NhzDCMTsLJ0eemyhPTureZzflJlHPGbp0F71bvzz5iW2r
P25K35GDn+5W7PjCwAmtTQ5sDYqmzi/itPUpxcxOxBshD+luT0g8ehos/98QjQwD
vqmvv+Jjeuobtz+KV9BGBC1jRBV8WHsXQS3h10clQMbAGE1kF+NXSs0ZsN7QIZJG
DrFxiVI4cQHIJ2Kz2mNAkoXGJmJVX6cUVMER0aTVP12g8cWxPdzq2Ha5S0mOLarl
t+0nvWylKtL3+pJcHKBNxoHvC3aTcTaGwYtFTyXT9YnSgiO7wLWWACmkyAKhcWcX
bKaPrOQZhlBpHKp4jbSCQpvzBASljG9hSdAAAx7XTpdWWOJWqJdqjFkTqFZJ7nkZ
L/cpmB5T2GADf+/vkRRoVwldgX+tJw1igWRd4DLeczKjo6BGaxUwEEXAsITQYxZK
YDZOMuVx+0bsqcl/6mfkiA8RandOL4U8wOsIabYCa9pqjPU5rPBEg6Mjk9SCqBwb
Bm4JVGsR+rYJRKJh7uBMSFCU5A4XVBmej79rra8Q3aYy3N/7Qfv3gcRvX7i42hq6
2RV3I5RHGIGGOsHerrepVyY8K6q6zyw10lzjrYapbaAzv5L3qQPbNwuVVe2rPWzk
p+MqfUFAcGjdBDgpZNXgtsE5lxDqqp09e6Mxcsw1CsA/tsTjHspTW8QQqgfWihvT
Z92MSuocbxlcYWfgvw8VjAdzDnSshvSFTMQ9HSKcwZ6M2REGhtGW3wirH8gpbUT6
/ZJ7ZiqnRhNT/efAHc6/Yr7xLFUHaQKl3+RX9JRRH+JCiZ+I/EG5VTG6gLSN6VI5
XHuMzWpNZAsjRaajaJVdvP6RrYZAI6Dg5SbKSgrwA4Oj+EiFUofuXIiXWPGSVBrX
qDyYgTj+OchYkpyPJ+yrS18S3VukyqT4mCzQU/sQqocmmCzP72flg4wdtav7MCvu
zl3Fgzo69lmeXvHm8nbXDR3r9eK1DO0ngbaM8Ax0v3SKb/QKUIU+1jfRuAPkkgeN
/XJ00Sg8RzPW04UA1xTehND+iGNo17m6FhCunSomevj5FZDrdvP76fFT8MlsLM23
BYFPYRZeeB1KCLOfOicmhFSEzG4HYvRifCLoz2gwTnCywXnvhX8Ze5JUH3cTL9vR
YNJbb01qsA2EPEpG0G06wXEfGVkmOxcFjmIg2LAEluVX7lNqdb59t8rOYO8plMx/
erhyN5wFy9tGYl+nrIKDMUGKaMI88Twq4Nk+fbFnOaO24AXXFM9fNZoAtrfWcysp
vw9HS6Nip+ytUS1xEDOMo1Fbf2s09ne7eejvVQpvi6mpeX7ebpilEls3tHXMInBq
idettaJAaaw0bIAYzZee+whC8hV39QWTjlNzuR9U05V/ol+LsmyMoCGX+ZZu+3xK
vw0UbtGZ0EuEkqrQ3opQuqaRAd/F+K7+98+r4dLtWaGLYnmdgY/Q+C6INxmbyWDz
2BqMyMPBBleDbeTfOOb8WfMzR4Wb+lxUMqnijTa6ClngLP/T03TdctTF8MCWCcOg
vUFQQEyU9MCZ3zeyFIvWYHHnmXq5eyzF6R8wxihy/+2YZObX6J0R/XeYjONFlYV0
XXpQ+GA8vwkRuQd4wQoTA0+Ge5uxVWeB5XzRXnV2jKGSUDXWAUn8VKkwdjIABLb9
Ulz8wlkZ/+QyqHYLVYUDMrDYZzg0xDpoyLDVYkDgy0ScIWMR1w91bXJPcY4e0Fve
p1Weys99nv6ZYl91b1L6LnvmtOvErhaAwPy/R3196ixai3Z7WTXBJia0Ixkly+Mb
z81Yj1ZJGAfThfADk0F9XL4brpFXdQhDeT+31me9GOVe+fDSjGHGQScjmu2jadw9
hHe+YtEOAldeRpbidqA7nAi6t6GBImRa73bPtYvfa2KAqyWuISfO/5YQCwq/1oGI
OOAFEBZm+gGqF/0g6W8HqglvpKIS0/TPPCW1DZnPzZ41IvDpLBqnzJZlW7tzm9sL
ydYGvIGCjN1d4l8MEV3Z7jUpwMfAWJzOZSPx2OnB6gVYQxu5/+q+QovHfVbv55ud
yjHxHiDXbE6ENlhxZNODuMDBk2vP7f/d2sq6diI+XMvWKL0kk2pO629DS7avBjR4
+dTNq7ef5qODz6N9eGT76Lpfl5dmuO/bd6bdr+8r/ncnI4UtnKf2ONyVLVRSXI9w
9BTPkkTMHjcwO4LBbljCXQDbkADnS3aP3AcNDASY2BcX+pRmBEnjDso3euIgJLVX
dkj6gsvYj6taq6PY7665r2dqBKXSth9KgjxH8HnXxUcR6pagfDPyMiTJPysrSk1e
MYweECi2vh8fKRQNreGM2l97lKqYpjsviydFB6ftgGbMQORIzr/i2Gs2wfR+n409
QFhIShrF6ldwzqCHoQID2edA+WUp2Akri6BJ70JYwq8k7TImpRrL5WHROaRch6zs
ggjiUXl8RPP4GxnBGcsdNEiOtSLCkiVkHbIcUZ2cTdXIljlPIBTvK2LFs8vtABUz
d12GNWEk+G0zOGJRPUMR8uVUHqE6ppqHPDgRr9RWZyhCbeH4DVSs8MvBJV9L+WJp
BCV2jkOSRQxOZP9qCDgQaUwPDnrR2I0l9F94lTgd8UBIb48mn5pSEn8bRR2RulA7
NKHcwKVZSOSRsYAejHAlrsb7nh7ijBxLXoDSuNTECFpSPywOt+MYbdcTwQr4jFkU
3soKLtZO7ivZQz7YPlaTA79k2USQ5K2A0FSxFpnG9k6UPMiyDTePtgVcSWi6r6Zg
ym5F/T6C09f+qKHXJyRH0NHuIM6aYarirmEwZ5/yz5RWIphlhj02tAmJsnflXc4m
/D9SMBjMvs6l9iP+JtgXSVH9EL31zhalzlJkeQk7QjWG3KfX0TQAaGdZsqZmCu36
5BOlAytzZexSUIRl+VGJR6HZvDPINPvtvDiZKZ4XfLAepngxz1GKk4Dy2P4y8MZL
1PmoONVi6QnDlQbx/fH+6SZcEpJj16pAX5T3NsJwGEW6a+pcXMiXpMhoVJnLve32
fVRfgvp8wxUp0rEzoOGQtJznKRYSrn+ixhksWJ9VSy6o6imT/UtdyvBK3anzI2CK
8UZ0TdjCrOtEKWET1Keu6lOWpZDzmD0e/rYxLmMQSv+j92UERZIhyBTiGRXeFnKj
QDhpJ7AbaNwbWYdNdFJP+DCP7D1JGJRybr/3OSaIvsrlndOz+lD67eCHOFwnG3Yf
9InFFUk/AfmL68drN8NYoKa3DtJIPm894Knyqeuk+PI5W9ekdhNjObuz88hvR8Hv
kgFhzCnuS8sm0MfMUTu0biYu9rBRXNLvYlKTO6nBZ873wtHnrdFD4WkzJZ4FLtD5
vvNJf5Sbp6muLJq1/XczXH+lfKHPkVznr+/fDBAJu9dpMHjlYwBtEGxf2rVvlyhi
jFB3bkjr3aRDpdtYHkVv1cBH8FwEDevZI7Xh6FGAvMu4x+qIamCsWJLzGzRLjqn1
j/h5UqKyLmeyX8QCdHNhyv26nNCKjqz3arIUuCMbu6TJqEFVQTjvsaTjQj++T3u/
aaHrkcJFtirYc6ie7HAYSTfTVUOGV8XFAjFhhrlmgrVDa8GcmMgs16lQrOs/oF2K
wpSuTAf17cK+bwtS2bMP20/JefrnjBkvmFfAddosHLHkDtUPVdRCMX0B+WKB8Vmg
4fEDetboa4XGzBDoMnZJ5Lu6Q5gu/PaaSYwMAogzsZjVufRN/U9sZvYToLPjSRX3
td1kUVVnKZ9j/n7dvMvpsTFNI9k2DpubTfOCMnRGpIfBO2YLLHMIn9k3G7yZ83lm
31/yZICQoJmMqbEtYOkGdEDiubx8nmjo9yKIx7AbzMe1mQZ4/XKjZT79MN7tdWTm
KF9BE+T96+3AVDVk5qdO06ui8sRdvhZ7qaDJ0kgNre8plhU/eacydrEvRdUi604m
kFYJU3Tuv/Ij3jwHfVBzsMghGq8hCjHqHwlsiCotxOO/RIBSdZpJSy3bNHgJBXOe
erJ0DoG7NzZAs4bHwCuo0deRVuW4gMHt1iBuN05XU58/OHoSlqCnXJU4KxTKdLSW
KAiIA4LAlc7UM/VcVGEKsGj2d6EsniasfucrujNHwKK84prFVLaYq5dDmdAJlu8W
1Hi9FGPFAOL9yvAjvxO4feFjNGVaUiIIjm0KvEWECJ9imm3OoVnNbzP7r9VEoUeE
I39wob9dzGJ26uJNVIFsuLb8L6AmCnBSKf5XmIWhmwS6CR7WFR8uR6F3HwFS3sZ9
gPkCbQ3sXX+ry7S8+AePmvG03TihMIHJ3dnqHtAW8Zw4NwRYWPar7/nbBk8bTsZ8
ocEzPkvBdR5PUvBjU4KM54vYC0GiQ+RQouykoQ/PwALVzlyyX+Cld2uDZvrYgUS8
97tiAlrhIxcfxYHCD/+IgI61yDm5F9XWUdPG819Bd3sNDv/dACO3pvG8kiVVa7rP
8Uxz9uUYqx3X3CL/qGvvUXufIqPKgSpV3swLWq3zKul4qMnvyL41LRAHsresCIqC
J9zES04XzIXi802mm3qMXmbyKrDrIc7xxkcgh7JOUY9Qh3Gp2ygvYQ6wJ1zOx3AT
OJwcBFgKToG1eVvTdVxy0VIlFyGCbzLp5OJa2CrmaibnVE5mLMaNbx5Eu0PevpM3
NhxjqGxb0/5gS4c43UkmN7wVMHTF1U+NLKBUKLEqg6E8VFBNO+gHp4CRCxH4LeHu
Cx2DujhKliynNqjLrip/4PHjArLQPVPYSKlZWeEaqYZtoGNwA7TBccgh5pOxcxlA
jmLvamM8yQlmS+KD/gO85y58tSedz8fJaVyLBjOO5ivjvcFJa7d2xiP64x/3tJLL
rM18oA5XDIFlFyLlDrZ2L2kK4Viq6wzs6EQUO7ePgADba0i+kgIlf0WhV0JWQoTa
bXoCUV5MGa6il6BqYLs1fpySeNgWqaNf4lACDdo5JrkqQNFlUgJEzev96QbwQQdm
dDl9UCfmZ/GQrKnIub5CeEDp/CWOM4ysm5sQQiah3YGY6hOBQCCZYzScCiROiw5U
+4w2ctSfO2bx2LmK0oeJno4Ck4Tk8/rvQSP5MKEtNQZ08XvyO/IpOI3JQZipztOS
ZhYe4ZTndjWGLoLbGHwcaIX/SZDggsv/cEWnzGXBllF0yVDbX6oMjPiivh5OSDra
JKJH5LV6g/tryZJbuyNw86PmJfmKHkrRWdykRRRrammH8cqj6Ml4YjGjUJhBJVO4
ltYsqj9BdKay0Fep9oKp4MCegsjO82N8F26kn4+FLwXFtRGwmbu0SGP7X8PeovT1
fb956LZlZrqHMSYYU7wWGCjl5KPGqVmIcoUjiZB/u2jB4aNMVZl+pVxNeGjEtFve
bw9NfuT3wXbb2fd6wXdQ5OrQ/RKo4/AT/VSOvX+TElHdLY83muLRKzD3msewEnHC
SdyOWU4yaV5OLZrTjrxLd1M2Lf+6yEXEKfax7tve9DwY4XewWHM1rSo0PyGzl/TL
GkN8EI7/cfnrBWIvEz8OsonRSrdsgfnihz+AF1lPTZirK6zRZ0zOxdHdz9f4xTPB
8sIVH/FGif0NnudnqbW1ZGxQGMjU/3eeOVS0xvpesv3JbP9cTQK7QTaplChJyreK
uD90UKvKEDSrEdRoe2IGUZynLhQDnkE9Bzy7C3oWjo4U2KtS86Ghi3wJfxGNZGwh
8tsjbLTSAwB8SrLaLQR1LotDpiGWBkqCISigZ0CF5fI7RdWGGiQKzEQcg35ehrhz
SFF+uLCIKnlBMk2VtW3wJMkN7CC7HyHROqmKVQvHqNrq8c5Sz6hzQeE8KhB7xW9o
cIJl1i5IVokzkRl3nUjO+Fa5OcL95iGXvL5QZ8hHNjM34JhSeP4BR4RsxwbaW4IK
qiP/3C1CbQMtEesaeJrLBpWJ9QoD1CnqyU6pXlxGRkFnwJ4PtUFWyOnKWlH483Ee
h9bKw3NLQTDO9jXzuMraOsegVa9+6NlEPNiAuy45w4iyqxbEeVZfuqOxrcIHgNvA
f8o/OysPJZ0lta3bdNo0ZXRrkLJdRnyxGE6AoktPSiRTSWVboKHwSNXBmwpCY2jY
zrBL3j3JyUaPfKpMgTfNBIaGZI1pJGVSgQCA6g/NbNMv9iurxGdu1w3Oh+KuQWOg
srdnYG755wAR8mDjzdUce2Uo8go2mvGCzX/RyROygoGe9sOlCZ5VVZDnBWuTYf+X
9DnDtgwrtFfnCbNpRohWEe5QvUGP3d9LL5KTg6/6oHlFQQ/QaNe9RPeUF108/2ns
uoCrgLEwZN+NBbr8ZF6pRxvdqSGRjp2w0sJsOGy/k8MXHPPS0R0rs1FXGzTmv5d4
JFDDdUpDqY4Fn4P0+yfDys9YxdppCefkhMDdlnPofBVl5uPOHQn92/t90uqk08tf
xdlW2zI/RJ2tuT1bWB8MrMlFkx9O60boM4A//kuPxTEXBCAzsIh1pTRR15I5kmzV
C9q2aLDMLMpv/QPTCTeOqWjjjLO0XTCs6GLukwB2F3L+cTst1sA6fZYX+13Zb+Is
KgEcraWG4WTpHZq3SlM8VtSEuEUGvbpSvBE94llJhXCKrZSZn2DMbYj7/CVZIT0i
A8MoAt9Ei9SEKWWd37W3FudmTyPm6TdqaU+2caLtm4ejNsJEurJ4LoLs4q6GfjcM
qH6SgThI1+shMzrbXf20OuFs6lVk48o6FHgoaU3daGfL9pAvXDsSFCfYRg4fU5/M
sMfHWZkKAdyXrx0doGc85pUGpSMI1TMm8m2y1eY8IYwHOPV2dARrWw33qwHVAoRU
Wtkq5mqwxa63i2bELjnZMrplhWBhtuRq+TpJzAvXpQmDmBASyKFvnfj+l3WKTv3U
fAjoFx8PEVFvmjTnSYySzyTWF7eV9hzWfqeZ1IjoFoe45TXYdXKQelYAfuMb4JQE
WxAUQwoiXPln78/gr0VhuQ3bUdOH/7Ghd8hNVUk+wvliBsydfYwaEaDANZE+nIjs
V0rwK8MjnOMi3ll5GrJ6b3UYk+4jmnnn9Nno/D2Msz+YW4gYppOUlsAdyfmRRY+U
/qa4hLs8xmhEk2XtwncYOQV1PNu5LjwNaZkNIhthy/6j/BL5voiRSgF+fqfz12vI
lLUmXvFeiEuk5UDu6UpWWPjU5XRY2KUDmsHlMjLAzSOL9aQletaWi/fC/Lip/Dr+
uRnX+ksoZXMcUBkfBW085epSUXa/CF5asC98JEOSvuo3VPRM7zzo4weLXWOEVTnb
bEe0C7zygz7+m8pPEF9ghnCg8DvtQH4lAPIGHDDPMyfYuHqZJ7dePs2JGbwtY4R1
LpqVQ6yYaVButlw4mana8Oke4eEElz8F12TA88kYWgIGIjAdg9uGMHoUaMACYzIf
Cwl54rpoOS0H5qucpzkzRPx34m5m2q6atDsfGt44SpxhEclHonY6Sjw7SB3emQcD
TQBrrHx2XAFrIfyhmM1zkBIyasliypR4rZ+yfqbXt1RH06v0F/+LbkD6wgjH4eS1
URN4pMCDaT+3PD05bDE9chC9OPjtuBIZXfZZSt0jYX0zprkplkiY5+w7fI39BZgg
mTpTgvriH9lwikm/g2xFX5nGlctcc3OYfFM5jbr7aVuP9N+10IM/pM9UW2QJ2/kz
neQoCiRykR9Ajl6R2rzPYf9JbZmTlILkQOzbwyMR7gs/Sm69xaIgHnEj8U3N7nDp
2H35tjJHFiRFxhNyXILFr3WaG1vrFOhO3kZ7l4i6HyNHopfS7daPTyFRPBYxg+BY
1PIX7fDU+kpLWjRfsfJ4ru8bgf328xBUYpcGE3+qO+w82x0kfPadXHKftLlJ1bqg
4Dm6SqNtQSRjUbqPlu2U7sM5glNTboQi6ZFfQii1wQcAF+xaXL41K+C2JvcRA6ge
t+MBk8RybtxxH51o4dm0CJGKfaGOMq1eobli995Aa6UAnnR0v4EJAwtL1AQiuHNi
LRIhWmKlbpcPlaFVkShmeGbzi/tjngd++FWqZw8z4ByKGDK1XmVQSwQuy9jmnexG
LXNuDeHKzQAYJS1S983poPiGHDt50Z36A15xJF5CTKNf7dPOS1YpMebBxL2syWxT
8ZwqaYs8FpDvjVv4ThQzKXwFCIo73N99n8CNdAbgN2oSDVLP7tu09zEeNx4sJEfk
2IexKWkaNiM/8/j6RzSjbQBiVYIxlqYXE7v3xAfN+OUqKlj0E5mv7UPWt0EeosmY
0AGZEf9fUBlxz8dTJwGDPraC593FbrcOuwoTHIaHKtgI6cRx1WwyCdxxlcVOjDoI
w1zuVj7DFwXuw7k/MyIOqmEANQqZU2RZZ0Ore0vDff0fitzu/V8kqsjKtbjksIJt
80rNvcbCUiE1rt4SGaBJb3TDTnpXjizyLD5F86iYQT/2LoHSPYgSREmZrC4LqQGf
UUaKqzB27JIEY+7xy28veLwGq0/hk40IaTSvZ56wEwPIShNQLPc67h227VSISJVW
Y18C7b+XvIsUjnSMKJCMSxH5MY0+NdBzcTscBzu04ZDxADvN2DwfPR9Rh1ml08kz
xhFk2IFX2NHIamCCj6D1qn0njVpOFEF6OB/7dG9jQIkU4uRBUiKNsg99I+1vp0G0
Q3Eta2LQcG7QDJCJccqIcxwax589mlb/v0eFlvFXDZHLvOBaJlRZVsphD/ZmZ7iI
i58N5orHGVLWyMgN7HpIocKu8+YNfaDKUWSWI5kvkHH9nBv6izfB7kesIjUlAgGk
Z9AK6diQNcjEJfDBz9p7oQbQSiSI0/+kSGhnJXh/HbFzy+OjvV9Gmvi+56ueSdwm
wIGgtxnHBe1KG9F3dpSuoNzxSlcnb+pasvON7BNdvxTSUGbuTRUUw62cnW2CQDxY
LKU3lB0eyEUCQLIUfo7aU6WEnIfjoI0icPAf7RCDzlgS7Tux9tK1td8+kchutQSX
uWGp/4gWbhxi++w7nOF1gDtJW3gR0ohslbjj3/9QV3EXTDr7axAc0naXTqQke+SI
pKUcwxFqLGZxWrIuO5QZt6Mn9zxZLOrJeWbtYflrnynljpZiBqUVD5i3PVux4E0d
HdFCdxN8ovNubesYOGdRiS0Mt91dLVgoWHg5kchxeeR10slOPqG0ejUPWmYgptnd
3BqJm1SbH+JmGZlJ8kc46Ds+IWA4a9A6Jpg9iROuMDw7bYQFsH3c4+DL6D/0oJ0k
Pnjq0mY0Tt+pWt8ikYk/TbF35SHQUwQzS1gEnREwuZcJbArgXtqR+ZmnY2cTIbt6
nBQyR+B/ciIIyAInovUbV8nKPX3nXe2hl5+J0A4Hyxlf5dwyZiOmP39ZgPT7D1v2
7yQKWcyRl0KmOBjfHn1MH9sfVsIq7dZgo+4pSjNZPd6vf+owCzq8vv+a83hEnV9s
8y7Bik5Eo0DdS2ru7zssh3WQ7uW7i6fVKrH8KeAXGFKuTzvepI2zDNrgEftWTeci
yWJV3O4u1l6gdxabVTjUAdI+Qvsscq/6pq85OFCkj3JpQeNEJlxUzQrrKtgnvh+w
S0egxOYxq0UqrNeprP2uf1JRDa6WJ92myDnlKNQanmlqbQ5/2pyZjO79tH63/bdP
dgkXze7W4+pHD4xos6SPRPsH3PInHbOCP8TMSQZCfg6mvDZ/Xf8dsS5kiECFaN/8
iSAUE9EbXbeeYaXy5bwzYwmdSjbCnKilsjWScjQLOWcKWLDxMEM3DQBeRH1mxpcB
OuEB8BckkpLzvyqpAOVLCFbKqQsZUZDZlVEXp/n5m21T1Sec+5n1HJJOdSy4sTDl
AapliKnBzevQ94K1uszF/VQ/oiLr3f98zEdP7sx8HrfkvzQiHJEG2gbKqs0UUG5x
9Gwy5x2O7nue8lpLEqqnyJfzv042HhC8Rn2+W/wHGmigfVpaBuwi6BNWSk5oYs8u
8DhfBcYR+3Rg+OQl8JoIGbcNRCTcpfVpGZtVHv33JZtPTKatvmfZCArh0ihywMi3
2UWZQ2yRNveUDGpz7TUaJzRPREQ6HdwUYBy8954XRlTzxq2e5ZjebcCakQu4afPx
hhwqX5Ov4DUUk/C2bM+rM98Y0/N59O1Rdwfvn+r6XglFnSyiqWhw8o4WcqvsdIzt
j9TWL/FcyrzuFp2m9jT91j+oia8d7a/jSLWIo8hu0LErfzDmoZUMBb1a4JzwXJjM
vtpBIt4giAwujkdptrGUbUhLwEHSOiDKpcOpMa1V2IC/RsosjR7czoWKF9ci+uQO
uiCS23MED7mjYBEYCA93XRpqiWemqtLhtBUKtDn5RVYa+xM7SY5krwhdgIqQcIGx
PIiOrKUZF3geCzdS8hJIXj6MCSUOQTZU8e4o3bcB+52D7SYLfnNDfCK4/7AhIe8m
YeF/+s0JZHXcZX87wwafjVXIcrYZ9CsLckgCkd2TaVWlirt7zC989vPKGC6ZdqUt
lf4pxqCwEUckuK5EeBC7n3pbw/U7ZRpZxgKZtYJuklm/pIuM3897iPsdBK1bMjvB
t1nTisfxUY/7JeZjDDAB+0dHODgX1W//xZK8vU5PinuOSz7XB/L8KMRvrGAP9VCw
7gXR2TGYGvdZesNDgkQHGBtHpXq3dUL8P6tMdmU0kboAJuG47FEU0kf4YayW5L5a
U3j1n1/BMxLs63tw5Q83QA9JJKfz4MuitCZKwelgqEiqf06Vxi3iP+JeLoBescGZ
tSNwhgziUHXr2UEsV00Qhj/2x4aNRN0xM4lATRAykY3z7JkRL5LBpNtyvjQeWYVM
eqFvC30jSzY7hvPsiCBs7qpXe5o+I1t0F2kcbTpdd47Cdj9VpD5hOrKo2iNf+yIY
TXcCaNhGmRSm1aIYsrzriuMT5ZP97GbzIQtZbMZcaHM37eeuE+W+UD7tE/BE9gMU
II3pMJJfw+NZbcf2I6t5dLDvPaIUzXmeVyO9r5rrPlBUcrKYOdLsAZnQe4QkUkwa
09YlMAusLRHEvbbN+nVzEEvblQQ2jceXlcHl79mcUFq0yD60rNhuWRbzlVHYPR6x
g4IBAx4Brhh/ZEEy35u9hLDs/DkJSamLtUKArN620Bbmbw4tzTJniEEi25C0U7Gv
yPmK4ebgzIUieUodszTS2T/D1Dl1eI8D2KUnZwfRRH0dxRindaHPHs0BT885DAxC
SsZTk5t8Ym214eAgUWEynZfOcy91HfR2+XNHRpNW2lo48eHZNKt3p+yeYGkFij2A
XCSF3d/M6Wfsd9bb59IO3P5HBj3gYXtho52z+xRtw2J7b/7yiel3RjcTiiFtPHp+
kVvskA3OP/VYAqrCjrq1OrTnuqTvuttGPJgrONpnZ1/fyvRlWL9Vwz0Ix8T7YOCC
oMcAsFr8tOQN41TJldv/bATTIxxGLpmOXa4W6asYrwTxGB+jMtON0jzzMfOdAJq8
TiCJv+QgkxulfzJ/EFyIdH4oLbxKnINixEjxZKaPI8UN85GaP8tEpH1FlN7GBVCG
LNXTkfT+SAycErI/SRRULXBbYltxIuRyKTgrtaSm318RtcvEIT2lAlU8GPK7IQox
QQ21B5ikSNG6aN535oidmkz8BZFlCPazBAXRplMl/7Lg7aitM4OB4wmoBH8xMpSL
lHPpeQALF1wUIpM9bGL7hCgJv8jb+TNv5vvwI0lI0nIOpri3J5rezqdjYUsYeTfb
mcou1M7Vs/rTJN3Oj8ncyb1JTyRRc3LSLX5Z+oRKicaU99kJrm0xQd7+7z0vCnhZ
NjT0IHeDiQMKbjX2wqfaM6ypnn0gfTpBfW0nBhGEDO2gbZOAYaQwo7lg3iigCS25
Mmm7QsucntEJ+y3e+DaFfACAXwLkn5fEHR0ffeuZoy/TEvXH3PIVoNCN0EJkYM0t
utcAkhCM13WKwZi7sU1IzzXYqi2Y5M8nhXX8UXRato5O/b3aJ9fBxWEidKlH1O3f
5A1Bb3InymmYj5am+waSpGpS4iERwVk/XsUUB4VaVLg6i9B05kEvdmYZJE7l/i1G
ALNS/9dqSOUUzXzXIGRYvjSSdg9iuoIeqYHrvu4BrfkKiMhf05OpiAvqZ5YJPD3i
5HutDUtcz+GmRPC5i2g2Qjepei9NBXCo4UgKM96CCeqGB/t5urS7GO1+pR+zwPRj
j3jRMQ1/XNNzwg8oij6LFVkfwb4JAS8TpN5xsKrtXjtESNt7YzhKwiJJXjQMjWbM
9l9ALYSTXLWqZoT5ZrtRc+0uTus3wa0WJUhqL8Oeyl8SijcQw690kCGWzzn1QfHK
bV1q0tNDO5BackqDssuZfxGXrNk+0+sJ4E9DyaeZqdSxI+PFuN/LBVEZyjokbwnL
HXC0FJ1RTlA3BmsiS+3RArI8BJhS52BWtY9kdPoXXVscBilbKqkdXTr0f2AN1RFs
/xYZPiiGDPJsKPsStDgP2dMIY4iuZ0PI9RaLJunqYH6BiKmv2xvL1pPMjtEXcXiH
09RizOERAMLmIUrX8uOXCNQ/vXU2qWEdtGgdKNv87jYkvZr1fLxVM6VofyrV5bHJ
7gePKz2Q+jx6T8hOT+UZnX93lnbQr/Y0xKRMszK1Ho8Gd/r25HWFDKkbrnCLOx2C
E6sz/+vHfvJLqqJxBynDn+ZHapUcRCg6bzhfxuhfWe9c+xf4FIfbMznRPZrpFITq
7I4IVYDeZw+0T6huuY5rDiZjjRDZp7Sp5g3HcG3r5ffsPpTrNiig4hZpvrkc0gOA
DeaCIsPbBgY0lmP2PKMfV0HApu9tydCQT3qonHHz3EIPDIpj2fSRp6TOY3eXTHEv
6q1sTbZ1n9xWbjg27PhR5v8wlbEZRn2Sy7N5uPGs553gzr1rb3xdiLRZOEir+Ypi
Zlfh6EmeIKjHHWeo+MMHVesC0ysaOikJkwj0XIRfE4nTYKm04q4wekZeMbmu0JrY
TJA7AllJffOcqhYC5UjBnmwS9r2HFQMF89stsje1zYRymbrcbdYp/Q7cT2Vb20co
Z+vdrgVSyw8Kh7p5BUvyZLgGArE7fizXd28LUKbUuThTjG69rlVOwdx5F3v+872m
DfVkKcfITebB54ofzCa0mXXir+SR/VTrqLH9y9/lqx1TnP7ccqmThg9MtwqAGJM7
hZiwxHb6rYOLSL4agt48Bx9UkdA9cVcEaidkUhwocBicY2Z9w4n7gZSSH1aE4uSp
wE2qKNNuOQcUoa41OCqG6qwixDxDJ3epmu8W691A1dKti0s8QNumkQja45H5tyAd
4YXOiMQ56nOuKom6LGnjjzzlOziZa6nP01P5Ln7S6SIJHiijuaQ7WAMaQ+/bWzDb
mfYRfogRognA9ROoolM7SDx2gsuHxLOsGeIdDZuHw1plRGqodjiV2Sv2/DCuY3bH
7quli67V8QCOkmq5kgO2mgO568yqzYaoX2covFb9FV5/Am52rFJZ14yWOAd4Eeus
zijkRV9yeBUBHva0AIR/4XtLRM8eCvG3P5+hesNKb6cKflwxjTnxMADQ5uO/wlP/
o3R8kuzxg50BsFMAKH2d0vrLkR2jnbJA0XWMoOfycgQnoQlZj9JhCF+4eOIpRWn7
54LIV4hl1oNnuJtDkVFfkMPjC/FbbpHZU8evw3EacxHroviX45KkKqcndfWpMrP5
vq56KPJxnNcpYLwMcETbuu5oeilNakTMqodmJHHPPOcrf9Zi8vzOjBWrRWJGfMJ0
0XXvBdhY2lCPlGVuaLygV14k4tarh8CIj++YV+ebdlV3PqoVEGIkaGqjjIOk1YHK
RLvvZzDm2F8YBNpfz0LVglDTehc+Jjv00oxNTe2tFUn55JRKQmCkbXzbPHtzs6IT
r1P9TWKmGcXiY49okGu0qR1wL35pPpPesE+kn2tLqodPVWKURUzj+vfI1ckNgfJV
xQFWkvcYMepP8ENHtvKIJST8OVG/ZAXn5E6kNOp2XFDhi4AiiIOylS9pmTMaKl/V
A+6EfyRYYrV8Lxz92s6DCbkb3BPLfUSTZnjVp6k2wbyNTA3Qw9a5vURmbAKFG+HS
8Ke55QMaEINyuYt3TJ5m77lgDPsEW7tps4eOD6HSXQu7sHsC2FfiG3+9cFv6yYxe
x3E+Vcg/nQSbsVr9mww4V6pjqo8mr1c6DHvJHImvNOM28K8Qo3BVDSQzzT57gb4y
NNepdz3SO4308SrTAloGHAlySut7kdO7AnuzbhxipGATcFhUA+Lv3kRp3CXCYnLQ
WXeEaJr05tqX87fAjvZiRla3q/ubOI5RFSteWfeS+Clz8T3yu46ZbWLzqsX9y6kX
pjkzbCkrD07qmR2tVGu3XC2k8cUIEOHY97tkdiAmdq4w1cfALpvtzlFfDni/+YA5
/w5iGD1S038o1F1uWvDbq7DKMSoBy78sIxL79+OOT61zqojn9hjp178s/mRY453c
gz52GVWqPvdr6endEgIQ+7iNpMtmgCkhLKrCI8ZWJZWHM6CGLs7fNkBrgDsYXrhs
ogOsu4BhiEGAaHw0yUR3QYbAOP72mQMtvBZ2ghAe6lYzoMEG/vPJa/1MwFn+5uIe
dXw/aTd3tmg2nb+ITEoHS9aFq2SaqqfP03Bhr23RP+KLE0ufK35GPb7a97y63WjP
kgTbFvSyJ6cdTXVAnxf6zgJfr/VqmFyhBKr48XhMoybzuwrrisqB8QIyaWH7mlDb
Jg3osfECXUMJJQmh5BsOJBbsOOePP0TNccohVl0lTx1mPM4pknAZ6qpI9UtlaS9w
uv3sLWZrDcwmn8XAFhM7xylJtGBK+k1pRkr9wwhJ0+uPzLr3YnH3Id3g6/2dQ2xu
Tknwm6nZ2kSAm1uC+1jod/FucZTrOnv0iTuKniEOxNYh93+X1Q16UTXrUXLDvm9R
F4qIbi1gOAMMTyWAck71TqJkZoXibIUiO6BoY7r1PlxSYWBFvoo5L/mYnnUDptqm
w3CvSkxL2UxDarzyZtFE4odg3aNQMO6mcH8Jneu3Pprj308z+fMPHF9zAlbl+ORf
yWJ2P5OrNGzqUhtcpZVvFxB8FR5kZ555p4xWQMw6nKte9teblxAv4OG7T46eCNZa
x4CqpGeGTE1moMSeSweRjVXdg+q6R4l5qd6pJ1WIPMUQ3NgmukQdQ0AUJHzAOVw3
VH3ki48r9OyJ/V2sN2ZTnpcx0RYKHKgkpU9KrtE0v+JTb1WivF+DKiLCY3MNbLH8
jD/SzolDu9uIUaUzVNLF9Sf+UDlsEH6MFc6lUbgRUT7OAncM8NbY0cEP6T7ukpEY
NHLaomJQON5CDQd3QlYGc8ED28k/CGtINrDwlT0tMF1DJx4+LeMAojwegiwtgEIN
SPgaTsMtCrsIkAAuZU4QDezNlkwqvPmO1U56hV6dXCDPiglnyqmZT9yI8SPCrf7i
DP4RpouEEfWhQTZ/jHxFLgWnxXCsZMp3VPgzuBzn8NNFW6jXThzIhsFRzUFjSpxc
n7o+/w4OSPK4yCyQHtF6wqYFE6KsGu33lWe2cC48p/+fzwwDZkMJo7GKE6Ihfazu
VW53/VE6IuPJFormeFrq8tvDL2EyMywP7trjD9GnkuCWfB6LOtw4g6NMrm4JVgR3
nIYiT6Szp/aAAJdbpXKheh0diG9G0S8qMcZmaMZuwgHosvjCA0sS65EcCxp+s8vq
ly3/OwlI/REz0/YHy+lL8wCMG88KkJzccKmcSdjIom4UT+QdA1ugkFKn8gUWVPR1
6TqAnGfdJfW4RZFLx5pJ1I1Jl3rDHCkdzNZzU3cy0oJx9A0DZr9pNodtb05fWxpQ
G5EhFQhCqi7oYhTLngC1aOrI0KNzlyiIt36OR57CSlajqZlchMauk92Pex3LOsxL
Ln5iNYMW+mIRZNkBLrYtsWbIa8EDMBj4aNT3l+7tb4vAHTRCW8uE7XlNan0DdmJS
ZCuSRZYIsWAF9+82+v/N+G5JSZ+fH/1KB748vDw8bpZnSJrtoMr/URXx28dCgN2D
D4+GeCFoTGDbPDIVb8C3S45e8+1CfLxZe/FQY//ofFe20LEBOpalzaVw2u51AIEQ
ixO/mfOrABGFZhL3LQKyLx71vIsolgyX81L2as6lsTZJRhJcFMp/dgKC0D/vD1Yt
LK3CdsowgB24/7ctY4AloCqGpvs/tGlq5Dow/IrOqFBMw3IqKqUO/G7oizKS9FqO
akOYPf2a/UuwKmGKxLd5Y9hU+X2M2F5+k7WLgh6il1UDxrDbwnHq1OFx4nqMjQu9
Ot/IgdR3n0b9fEWKuA6JB5kfIu23mSoXTfrP9vAL8RJEiDI0D+pFw97ToJLxDuK8
C21nJ2qqI5GAHM9bv7KHv0IoJuINY+gcGvNH8WyrSxZYDfSC5ZID9mWCplmwRbBI
1TYzW+soFn1jZxzhOt71JTjZiMYStLPxZ9GuYeg8Yy4ct+iYUGo5YNgGSZrawwCE
L2BaktaFSiwt8lpI42Vq0paVXKKCSCkw+wKw0FjmhLGnchoXzGvO7p/crvZ51ZcK
eYl7gWlxSHHTX9ucOBMeHsCtX+ihlDvNpETBUhrd2G8GemD7x/nOmrc1ucHwf/Tu
eetyhh4gVVIa4M7GVjoIKV7RhEhV7HnVem0gEHwKjlgI4c+D/M6uFzaT/1kQ1CcJ
Zl3TbznjPxF0STeg8YssvcuvM3z8GCv6+CoNqk2Z0O282ngtR2Yt6nSnHb/5B8Vc
UN0THf6X4rsiGvhJT1tvqIf4kSLkfMgMPUIFR3zg71sot1zqf7S4Mz35bxlx8sf/
SJxQ9o1GFMzwMelbrG+MgLfK44tsPdIeVBuYjvArLhAlaKEH6cDKmllhlG1cpD31
+8M4c2YU0ZhwOVSPfiRpV/dB7nUvKLv7xongSQy6YL/+WEZD29t67m2EKdxgBVpA
264FCfUICb5eqN51uuweNrO13WyCrEWJbf6wEm6pZABXsi/9NLzSVjnuQLgPCU4g
wyMSp/ZshhqSwSRKIZrdYzdkEs81WMFn3fWj3Yg7sD0wpy/79sjDx5R7Mf/javyQ
E8KLcT0dhG4BEKmM7WXpGHzb/HSxVX7Qgxt/JAWIAmlmtgryt6pchfaQerCdEDwL
gldyCubHn2zt7xAo1qwyzp/ZkOmVeIGRpzkjDaY5PXQvWVn/o8SwGmxEGAV6bYmC
VALyV26IjIuixDVHMVN/GIN6qT6AJ+x89SJMei2A+v6Jlez5o8DcEjxrAw//iMeM
NmnYNIKaXclr9qFDfVr30nuxjrmLyUxaPfDIh8IP2dbzUpKeYHhzmcccpQq1u0V/
aG41rPJ+F5/FQEXP5RsUQc3ybYwntW+bYF2XjNC6XnIFpqreH5zusa5u3ValYx4J
8gsB+xST5cijNn1YseFM9OozyVGF4WFUe0kG/0gb4U7e6WYqeczeY3MxG3dlfvV/
NPq0gyHw2UF9OVDAbaOtk57I9uhluYBc9PnwVRcFr1rajQjuDn8jr9N0BWfEuWbE
OEWKE2EfsWA9kRrxbFvDEGD21zexyCFhmZ7eWBO1qapVBENXkSSnZA3DxrwYfJUb
uFn2yN+G1GaM6fIMIJrlZn8ffR+Y+ImpDtMLe2Uhm2XUcb+EH31lUGiEFFfEdYFr
dJ2POZN2MbHlaiqT7uDClXUejIchiCuAguH4jw6tcqcmTwenJoLMWxgl2kEm9Mnk
HwJk7j0hakVCmSn2oxSIblBVZoOD4s/R3ibsVDflla/oLn3tKF1r+/x1vdRTCrTC
KsSw9zj3T7zw4p8wV7FxYz8LSpf6/vXPUkH3OMsUu1UfEEs2Qs/FoWOQTlBIlnDJ
FF/S0g0ojqhNBy3BRt3BbfqmtCp4a1b4CXk8Ak62BT8IUyH98ebBt4uJDdp4u9aw
Rb9gfcW2B70MimdPSRGG6DQv12ekLFWLPyIICEPveld8C1kVMwf2nSfFHwMfu9eJ
xuZoKwKzs4J3tggrorGVg9IS8/pcuYvoGb4+gh/fCVaLlwZDSQNvVTE2WkoOvdaq
XjwYkhtPKu97e92OU27ZV7Ju92HS7y8niLrNogTc8osyjWyC+B4dD/Cmp41KJgmm
ga5+nfPVmVskEWEjmgpH0ujgoCka8quZfAgJhneBWHJsWFSWeBUoJoiVmzBPHjv3
YNsn6tmT2wQd1uz2v6KWj7Pp+Bck9R0JMGJCd9M8T1r1Qv/G4pQsRjboTIGxpVSZ
C19Yo3OTzMrxuyfIrahPOq7etR7OpuJLn1FmqX70RQW1innXgpyRFLzKCoXSihti
Cw8UUzpnK3XXuriYZmdpvSSfS78Hmg3QRxJcl9bEMs1JPnvJFlnHrJLYzH/M+0Na
fAI3kM8m2Xz5ZvlDYimrwwHQ6t9O2xgxqFsAKLezENMjtvs3HL1/n27ZKwoHPTkc
Vlz3ZrolwpByL/USggSWmHJPgCxs+wGjXDWLasYLUhtSF5hVTK3qxteEKnMpiWlD
BNF9DTO1oLG0L8LcWZXO7FzBjnwqFsfFrAG0cgZff7NhW1OGq4WSkoFjTQmpab/6
HO75BI0V3Qfm4ts4UTAo1BbjxyU8975wnyLyA34NjjCXD6G81bESPteR/tHFqTmK
bfLXratefSpuAPJ0jCZfnDw0qdpiLE7L8lBzLchUMhModEdAtStlwgQbwLXO1uWm
/hI+UPobbXU7hKJtrg0J1xnA28+wem7C1gswcU51F3kKue4kh4e1jrpMiFQU0N/O
ZxfRsWLPgRLnienoCB8BmhmuGT7oZdyLWZFBzXv/AMfmvDj5/WOslVO/GN1VqUd5
H0EmP1N3cpomByx51JssiTrAzBGAEDVI3currXXft5Hxak9g6JSVGCRDumaeR+BZ
vnYhZzZIMj516pZ6gDIwGHtLp96lEFzPiPdOU6mxPCZfPwrVQQ6fqwkIThzyryfL
LwdyU5+MhK+X7oXQove6PkAV/1NFXxFf3c7+ZxMsayMp2SKY27aYcUSoemvD2arm
o2CBt2xSaXbhBN2qvBirVAQ5iiTrwlCcoZLJ0rg3wLSGghO7ppIBl3Dad5cZmutW
GEK9r39p7Gn8aNAylS/D7ySMG4BbUv7uZZsH0QLf98HXsm5YGXO2HnIOdJ6XltaZ
ajzaKQVBSll6VbfALQ+Ovw4ErWtn3CuRNEFcOmGiLFI3w+gMq7eRUf1eiVCPSzpR
vOIa6UddP9/93iNP70eJoUC0bN7Xu8mX96IwFQuOLWPllaW3J0gCZC4p2Tt+yZt/
cVgoqmXJXwzMxdF411cEqWXaYeA2qM5g5ZViiJC+j1o9muAOpD7EneeIMqbX0KA0
p8PqJeTerm6mRom/gVao8b/7xieivBhJ+gIuh+rirlKDn7gNaIf5qybzo2r2r66p
eu5UN/3zmsuaY69aL2mREafR0iLpaNGXPl1qJHuTbx2rDYH3xk5aWDGz0QB9toBk
f8zsYp95LBVzdr6svwEiJCIYrA00PkkXwRtkhMrgeTLkFVzwOc93+TICjaobSb41
Q/AU4X4DeEYeVU3mYmwfhUgVyHC95iypt6Y3QlzQJ1BLxBfQz1P2rTFfAUkS2Y4v
kOdxj/7BQVV95rOOLeRXdT2VhIaba3uFh+iNV2hv0p/G1mat+4kY/Uhxc006amX/
Hjne+HGVRn+HdruBzr10QHzE3BYwuGyl4cs38kqfhSoSgq9JcBq3H+6KR1mF4qDr
OzwzLHkZQhQWY4Lq0yfEk5OHKTK9xgW8Q89K1H/R15UlDv/k1k23Q5zF6kDzLCfN
yzMPzUfcSTWycMwj0XD57fiUeRx4ko/7wZtMPE5tw21sadAryZh/tWUrQad9dhD8
6orZE3MnDP+Ca+SLZEi2Ls0FHRbajrokfQqF2lBqmLC2ho0rjbnMcxcvzZA6Gp5G
z06ZnznLUADCFiANTcB672ZsSGCWPGgMt8RI9irx4flFIGDoV1OccRI5JI5riMbK
8zryz/yIpgqXjlQcpYdKq2tv9mieDOdCtsgGueAjqdkHOwJOh2BC5tTPBX3WjYsO
znB/E0dU2g0NaGzUCEertQ049vZsQ8UQ1MsXC3HQtQK/Km/RKiXsxFwoCNZeG6h/
HFD9bPWW0oiruDOvhKv0rY3r8ENKqCV9OVYJ0t+nwQYlTmaNSYlre0ZTtrBIsTZM
MPgQvmtGaJc96sepSYaSqEXtrL3IzwIlX+k6XXq88aejXmQm7HZAg0btYAerQ472
FrvbmS5bM2+I+/iWNnwWyX0xHKJ117g4UO2PJxaVljoKIFVNrAjGP191evq3EXXL
ESxMIxGAQ9azTV2sAwt1fgbd543hIGLfsLyoL8GsW072sEVuQAnpu6r2Eze2DYS/
ohm4CxCpCag8FKUeyyd0OOvWX3ma8ZzkP6qLZZOsO286tN0bkvyvkG3Sx3cqeBW8
PK7jkaer6DU6r7ovDXR5jFV5pr4g7wm0ra8CqXlohQN4amrCGiNQVxk0ZFD2NgOR
/fKFooKgB77CQyMC4Uo3tHXWg+PTvyQ8tUwLEtXJAeL6d8WTT/RYy0gm3L7zVMd3
ogmG9lQWcyZEpDjDgk+ozUH9yfU7QTQqyZPMMv3HBeIxvzkUMLCm7/UluTILDOoa
N5h6W4PsDXj3VqIUEKBgLe8VfS4ShR6+IEWqWotmIfzvcYyxmwLtBsKX/sIf4KNf
TTfvPY26Nzh4j/WVc6RY86UGJuewBW/vqslj3OIX0EVSgqxvVxJsiENDS7fiOvqv
bX3+9Iy9L8jxuECsTdzN+8KdAOXTJM/qKTQp/4Oeys3bnQJ+2HkQxAar24sZFeOE
wYrqa1uBaW1ltBxFOyRTrQXqTN6J433hBC3kqn1KtPBfH9dGHB44XeBkiRAQwW2p
uCfufkrst1RuU3a55BS5VzdMu57AXpW2BYlqnaclxXnnRkP21DozFV06QTLPiirq
x9E7cBX7Ror2bNJF4UXYrH0SNSlaTAOLvLyzYwbniyvwj3c47KimmG4uLFioXuoS
KngWX4ZTowH/RpJgOJ7ei+rKTcIoIAw6yetsMPamAj6a6BDN40XTagtHmjS3mC3u
MccjN82BX/wEHOucbiMz7iAt3/Pgdg9cg6ZlS2gmGso/PY7W7NAsp5qB+PAiKyxT
6shoJ30EIGu08ikeZIp8RYESU6ikz3+Y7py6jrz2y0AWIP1XbNF0ON0Mx6N0f/LZ
s10tit/i0rOMW89X2UK3Qok1kwrZDrQzJJlnu2to+XFj3hGHyKNR5+xRgQq9fydB
ggTy+HXbirzhcyIg32ES/2/LySZ/AAAMHfY+QThUJ6101MHjBXEfR+tmpjXtgoDh
8l3JH/V46bRsNiJbTcbtL4XQnKFSfyTndniYPcPqDhp9gqUfS4ZkiE2S7KdZctI2
IZjqLbo7TpKx3OFbCl8r/sqNfvzwACzO+FEJ3Spir1IKyQCRzJqn/iYkChr9Wojc
77UzE0lFvVDMfgaZJqcsbUZJhiKMJ0woNZzQ2xwGGhWEyZzoM9kh/Ch8kBD8KcOt
3wFCgpfSv91WKzXD9qqhf0zJ4Bmb3noWVpM0uF6k37POq5gMmZ6UzsiX8+BkAiuW
4gZgGECOPXEj/XwpIGxZVSnmICVJrj0KvHQslQPOJ24tYfwum5nQBISrMRhO+haK
ji1B4rCNk0KaeqHALKxjb2rjjWQk22yyUvW6sbe7xLuUn2Pa0Kx9WFOh9GedUiie
iaR5TvHZe5PiG7YrumYPXP3pEUe22uosydG+DY02v/91AeYaV4p7oeuB+Ac3NAYv
cB6W69DKLOOn1uwrcrVygvixvZ3MsMHcQkRsd0NA8h/LX8MnQsMWEwd5cQvGv0F1
XQaoebtKa2F5eSXB37o6QDgmU9CpMpBuHx3OjgLsge3hL0zjk6I44m3I2JjvHzka
xjAT0ZF6rh++fFYcmzzO/TMI//oR30LZ8O7BNw19EGR139HamH5jfuGkwwZeq6oE
oAXkd1z/8j4pIDAwY+gLRf5vKRNcPU+/UZrh3ajA9bD3MrA96qswTjzgcbs/F2X+
e3dp0ZxcHx8+DPPWxpufyJd5O47kro/z6jMdakb/e1OOozxFt7KkdHHUAC9sO2in
Ojpfchw1jFhKdq0QV9jyHhwDX81tFo7cnWsxKial6eyhuJ0pDxiGpTSBOdzORSth
YlNFvzHlfauq9Y6gdgsSoV6xarKkO3lTXHtufCU7oRvvY+GO7KaLhoJngawX8C5k
Mp1wIQVw/Z1fQmCEnEy6st4deri3cduo6lqNoYgNKeB1jXrlLTDnqRx+uP1bVEBd
fYQjsKCH/wXTPrcavPoangDq98T5xRj/Or0Z7b+qsQ6Y9W3fMfItKoxa1OhZLvaJ
Ntkg08bGHzKC3fyKmCEDlTGmGBNNqSmuAk08mYh+XJJljLLZhKlhT5D9v3A1l+0l
afnFTivAb3Dm0T1MGjoQtWlbqID1NJBpAn9vxApRl0bbSQgC54G7KF3lnmsBGF8h
3RFfCTi/u7UJQOkDqt4SUeA3ijSHRJ5oZ9Y64SF4DTkpRu7IvWMjfyf3n6iGUW4u
1Q6gdwHlfcp1FLzPdUXF8y1c0QqyD2CgI7JjdKMiBnwcgWnT0nLBG/hQmifcNzix
prjfsiWpxzWFvWGUf3f4s1VXDWQazIWYwPbQOygWFwk0HOPo47Llk9haLyrGXnFE
Jxi9JaPuDqsMuo03gxkGNk6OATMlzxt24giTAcyC6rr+Lze5lTVndPXm02sxjRDm
IyGDdXXiUdIVuz4hahVxOIvmBIehSjaUX7zOhHYv6nMsHKlzodSNtMvhu8XYaW5U
Wk6p5kjlu2v1hsu7Y9EegM1Tc8u57jgn6hiPsJezigReX2rEhtsDMCURuIk+b9xY
nFk4ExOvwEvQ1LFMbBYClDGxMOVUZTjLVgs17mOg+wYFBw5XH8sphXAEJ8RxfGDs
SMAOiQ+JlKTp9XKyZh5qpIuztlBDYz0tIYnBvEOBjYT68KkdJQu3rTOF6tKln3e8
7PJ91QaTs+EzjN7e3RqnSL7FPkL3qtOzJOrLP0nHLEcuTc56mf2bMF0zp4dcGX8y
9p5ci9WW0cdD0unST56Or5cuD3o0PvbIK6pHc1C7YzoIHw8HHmWAui9yMvOvKdJE
yHWRqJFrzKs+5w7RsS8RVh9Lk3iqhr3fwFpPswlFINdoylKaBtKG0mBfoSdGlofk
Ws526FZSPL8ff1sQBU8kyk4AsHnv+vc5dcVzxceUJ1u9RMGCQI0eDwaqOInx+7KQ
FQ01t7VlBPri6ALCpSDtaY5gGWBu+Qqh8YpUSJSlA9ImqAlgAVyIIMwNSAeGDRKc
0U/SQRpX3D8l6hLHjLN6C14mfkfzX5u+4wWunYcV1oi5v0Bluwz9OC9XtrZUvBIg
WhaBv+hfD9rdT0HkWBWWf9dLkBf4RZD8InK8CHEQOZ7qmfN+Q///kj578xc18vj5
zhuTuxiuPFizabFu6gQX9nuIrYkBPpvwZlkesTt8eZxNpDhceufE0nwRTfq3bFUA
J21aedU/scR8M0y8Ugms6bbwv7a+8/T/czLBgq2o3iKh3SBwgoMMpqtgEKtY7yvV
8dVJZOp2ecKoZqztGKz8EIwAWKZI5K8INF/aXylFaaJoreDCu6dZM3n1Z5/9ZyQK
6aR6CpKRpgt62epK69nu6FNB1yuXj3okDatArZXbXzr3ICvA6wBPdV7AcODRxI4x
xgpKvge3Z68pKYspggy913wK/ghF8JLwNJlePOCE0I9HfJuIuJsgTi5JEc+Xz+zF
1MiJBJJ6N36LePaDBz6zCd40jfGthuBanJL7LcKNwsXCImkC0rHsHpaDUTzABg/d
TPqo3gAnlf1d3RfLs8BbgXxOnEHHPsVMaxZJl+ZKtMsE5JqhJ4Cj2VstczuJyKC0
Y3L4ONHV1uHivcmyHxZJrp5ftWqg83XchKeEAjcn7oFJ04kXZTJvwCQFAb+UMfas
PgQ5F5iPTGduHQDo6spFCh60LBJsMQbTgZYf31hXZsZQHTI+upoxmbgySpOJ/9l2
LKPYbqVKiia4uoT9Bpgngd3yCgJE+id14VtfKrPOpxDefUSwPzk7G6ZgW0qDpLug
QMBq4mN5i3pK+QOxd0kSVkbMff+hGJukq4aP0mly3KgtiX/0VP6drPSI3vfcx2pJ
5EBLXHlUoYFh9mnJW8xZVfZFfK2mvHGroQGFONmMk7mAiwJAdl/o3X5urf1Am7jn
vGC8DI2BQqedLSV6/r9BI4ija+6sR13Jr4Du/3/ReaPf3xCoi9txm5x0cKy0Y0AE
fYirKwYaoCk+UChXRRKQcmhqg8fu+X2wS118XEZyqz7P9pyNZQ8PjquEjf5kYVQm
a1FYadzIYEgjDE3SW+AdGjn0HyyPCjfpSMFwdaaC0U0SUrPqFkry5fD0t2yfseRw
Rb0mc7xcuUqvLPHnQHnLDYwbBNS/ZLFniqluUPRav9y8t3X4k479tgXfJvyYEMD+
fo/g/ivbiJnd+bGcCqXDmK8KZJfyFPsyLigQGTp/3nBS/zUUfHgUNFWzpIAQHh/Z
SLFj91q0LbU9RyKMkRd/V88fp2Mw/rD7Wjk8Yna3iDzkXYcf1NXKT/EW/fYEr+f8
r2kyoh6KSDGWRY4Pd5yplBtQj5lKx8mc3ckI/daBDKNxiaf3e8vZC4+cXWYvczGg
KXFGncStxMBt4jQeQpt8O+5sM6lFPR7I3ufM4jP5vWrcz7wd8+7K4CqULOVrk/bL
uExt85AnOXjh4j+aktKXCOH0wCfcc13zhm7Ry5WJE/zlxeSmLiofMspe9QzUbiSk
PHUwLVB4VgLtF1BMLuzxyDr7WHv3yz323YKTO39qjqkULMpUT2gx+QMPKCVu/4N+
eM/4adMxWPcQL0x9z9eogiRP46EdcGJXdJGdl4s7O/ojnBeHX/SVyacNs5rW+uXN
EgUcj2dV+Z8vrRH12hRjOX2n7HT88luKAm1QscOZvk6k+e2S+RmxEuXVzP+hn/i7
GuhOm+xGWfJp+lGSDjMIv6TAjcIpXVNdu/Ivby1wc66cAEA7K144l2HUA15LZTTP
D6Mrd+nW4b0XCJA+vpYXhIhA68Pw35K5WbvTl1j+ybjepYSPMyiB5RS0kdIvumjB
EtbUCU0Fs7RhxTSFGY5TloTME6jdSp2dpEw2cGYGq2HFeKU9lakLfXlLtgg3DG0H
8wqbQIGU18LDT0HT0i3BVNIb2ZyA7Nhx9Ou2ntCeGFuIgppoPUCyQw/YZ17DgCRy
RQVl52hzaQWg1PKu4JsUOhpJxnjmaSplteiA+GAjAKiX8hY0u76S6sks6ty+s3wp
Ve5ZIUh+NlKJLa2HCnIrbKW6phFYoO8dnx7wAde+xOzkkME1237oLK/1nZAgrtfL
rgnGkbVhfyffu0B+/3hkljoayIJwsTvyxk7w66YPBDIBe1hlJ3AQfsiZVu0jhlYF
qMeI5j+DmLnvcH2Eww9OKUVzkQ72+wFUSA2Yei35Ud6TAS7DL5iGtu8fn7a7n+YH
m33km+OO+u6968LWKfNOyTpJnbJ8iI1BFvV8YANwulzNIzMiV5A5/jePBOpdR+6a
AeVB0GzeNgwcXvDm1nO9q2B8jiBHGQlqur2ERZb27bUut2/QqwRhjc4wanxAYf7o
YFWCJ/pRzNRKGaHXApC+l43jy3Q3+wZcsKL1o7abpBTN3I3rjCQJL1d6ciMUibBg
dN4DRqlQ5S1AZk3TGa6xrXuEJ2PpAlaJ2x+4Cb6skMFBuavc9TdEctrJcmRp6X22
53z+QdyOkG011sQJgsuUneHsX+KAUzllhcUkYCYR+hVGhBHLgci+56E9mmiLzW0l
KrFUjbANeHyFOP3J8ZC6Z+gBq0FQ26FET7RiiAG4Qpk/LphIBl3VT909CthBaNiV
apAwDsrWahZpOiFdNIssN9Odwzn14WAUfJdgKmKXGl1vHkU9fXF1jokfJ5dHqgZ3
KZiB01K67txiV61PBt2ScQQ877p1hZIf2CdXVd38VhEBfn2Ce5pJAloaY4xjTAf+
6ZlGWc3GT33OrOO8fkEIW+5tZ1j+Xk9BAL3pmVaCjIztJ+ywvlyjthYaCYficYeV
iDAD0QawRnm+ienOgVRRUUj8sJvaKJNDdZOatqUeFJF8VfPLsUtj6rmAlVWQdaBk
dqty1ctQBqjjDnsYp7Dy/5utbKJRdS2a3VobyiLNQb6D2Q6ulqqhEplDf/uVAqxj
/3N+hSCb3PdCNBe6NfOcRrBOtvzOcGM/B20eCxly5GRy0P10LxOwXAptHCkcMfZZ
8LeD8tm/WAATbm6iBaurzD/IvqUpzYh7O3WthhUKMNMq8xJDPgyDu52x/hbFGAN/
vPfvPS70jTgOdyeJ+vbXn45A+yEBS5Jk1DAuggIhGtvDF+BSoNWvxVbqgPjVW1zM
qHAfvc7sPSvWAvudIOb90BY4StJqJfBn818pxFvw9cWpXjZAz9ocQhzwo5Xv9Xh4
yKeg9vrVBal3XlcJ2OTMIlgWhCB2IQhFv2EwE0FpeFoArX47dIJyPWDSLpy6MLQl
EoDQ4A9PTSIecrz7Gi83doF7m7HSuuUaiO5mCdZSypVc+uICIP8yNb6qFl9z/jsR
0oMqXr84FKthntylKAfVvi+o6OepKUDPnlvpta22IvBMQDQMvlPyLpNrrMDPLL5N
31gH8gkhYMIZg+cfEZ4dA6wKHX0kQlWS8H1aZcQcFwVena8NrBTxudJQfDxbhLON
OnXlOHHs/fJnRBLr2Pv6i8LrlWRu36m2paPmwi72BuHcjKiOUO83jSk/QWcMANdv
9thSYXVvOqvEts6MHQaV8r5ZkJIsTTpHQDKULqJq08P/zU6t3RYcwyHA3jO2t7sF
4fkiVKLM3I61sDr7v589d0O1y0HyEvnDjTuqSlly7124guw72+W64P7Du+Dz+p11
+yim0CEQkAb0QaQGbFG3Kji9hDIx9rsB6aOG6eH829pszfNUI3xCDHkiQqOsnP7/
xZOqP0Y6HwE1Q2sCQvhuAeW4VhHsWKn9pppjGJD96WJx0U3uetCO1HKs8PXphvbQ
pmoIOHOe0yAlth1MqB0ou9tfgs9JcKUAP5D53xvic09KTQ0CGYNZ++hMekKk3f8Y
DEY/otpkN53GFy9t2xUwsauVd7kZy7aruf+qIHU+CFuyspD2eJhstjzHYuBdaqWZ
Nwk92q6k6ovCsH8WUojaem+MPvI6Smz/k/GZ6etVggaZi8nZ5IQnhmAWIzj5gshK
AxVyt4+pUjp+r0xF922xuGKeEDGPLVZmHdQ3R8qCA7+ileW9pxnaNZpM9lbU0Qm3
/u1V2R1Zz1N4OHGHevNLIk9cIEd0o+vFDK1GilPAhU4M1FDDXZob8wz9i6lqOSfK
MJdP4wEMMuiBXVpJCmGTV7cHd9sckGKOPFsn/icP6DjlWEEy0ybTd9MT2AHK/4H9
XyCvNnhkgXJJl73/UUwBrtVWz1qjdQk0YppA5iFt7A31Wj/SAYLNL+FzpVz0fX1e
ko+F9HaJ6+wnWqX9hWvzMGR9cJuNOzQ+FuHbzrLntlsfvR77lUGYYVIDJrvTL+Vo
7TdBT+5zOx1JH0v3oRhQ//9zwJc4BtHdPIRsLXLN2dQuu8fB64BqQ6SC8XOpMYpx
pOqkP3ks0125ZV9Tus+L0aMtHR5xBUWJmkQ6/lZz+hi2nUcyqnybtyzks9BZIAOe
tWuTryhsI1hW/5y+/BtgkCcb2LwRSB7X9u9cBYTUM94bKXGqGg92D4UvKaDDTMQe
0x165g9xjx5R6rmQH4qcoy2MtV/VRyJ5EAyv0S/dg1pE8I4m8HSv3ZnZFbeMPxfO
tHMFEiB9pM/koVEmetk1eR2w8uHnOur6afJxgZB4bxndEAsxilK0UqjvdMCTcKib
GbEB1Gr7GjNSrlWOalBj3jG2IKPnuwLchPoaawLZPeN2H3/O1le+EdYHE8vPBdtx
iwSK+YkshOdZAGSnbhF0HooH1pyfbOKVvopr6xDfvjkQksdvpcr/euy5zO0KmGuc
kASBLdvOLoRJ5q/lXP1J6enuTZqj9MOpBWiF84xzKVZmie063xJDv3Hrw3BgjOw3
GlYP6N+iCwkQyvfw+NpQM4HyUP3/hyA+b3f3/75w3JvZsOnfomQX53q4sGogvl3s
GN/vDfI3a9HzBCBr96Z7I6Iy0CcDyg1rWwH1cjCFpe5bp223JwB856x7LqeXMLpN
p0/n4XEnpB/qN1z4mvFYhDOSvEWaMRghMXo+d4malVkGiWd3JkZOkKQyX3+HBFwF
Gbc0sv2C/XKcHS1xFXX44jMno1y2o0paRbBjH+vW2tnCwbZ6r1OWCuW9YXe3klAd
0B0ECsCuaIxNoEM3cw4FPvUNNvai4xRTjF3ifjvghPM6QP/zfqF19aRH+WY4lDn1
nybbfdNON2b9BW2izZGEWSERpeoEv9ozU19QUPLqlnCQO7sznhuHH3itedi6sRTn
zEVXenXC3FqqpMjAyCMcLWx3yY6Ycx7/h3eQjUq4jcM9rIhRHGTNXfWrnP/eT9Og
lnWAcUhxutFCt4LRW2v6VwtMeAlYYgeRmVMFZLaN/SsyUn/7xakV8Q5K7zUbMpA/
ETI3ckkFLfEMGuYig7o+7atDbo5PrhR1qKNDvxHzlsh1YhFNBWRZjga/QHlEoYEf
uNls23QFlst0+MZhfstpEGbgzM2OwccZuON3/cPJ2McaEs4NqZCXoQIc1z++QoiY
868j/0NIzDHTDyaV1DjO7mDK7Hmz5k3rJsnGJxp4A13eaRoX+iG+CaTAra+GzK4F
eZxmb8BiVEOOubWMAs7Hdam19xYNwJRbu0tza4n5B/maaSGLNVqtPIxqiLcoOFQ5
YFyJFhyAfvd4Xu/GCEoDu76H5zEOLYxiOliSlkU32XHw3ehIkB7nTOgdiBQ2doQT
v7thPdBdPDNN6zGSHVGYdaFfVrWXscoe2ptbWnhRKJ5v4AiQd7zqzm72Mo+FUwZb
/0bBObQsRy+Cqg+aLRAecyiZBZToMDU72qbtt1WC+Y0dqdM6axy63iRpeEsL2o5c
L1N9uiy3lcl61h9/0T4Mn+2cKbyKduj46g3V3m6OVg70t6ygQoa9/tR0Vs4dsO9u
EmkotAGa7clBuBJXASewuWWTgYP7pE33s9yNxnALwaepEwMwLz1XE4ceBRu9wtJH
OoabFIgPU/RrwdjO1gRp4Ivf9/o9TxDGGuGiWRbjjnoixHyMlTbhQ7mH2R6namhp
XyP7CMrMaBJLcl/5GpRZ4MMJ+raMeZi1mOP8YE7EVvU04GJAKVXtm4j6Ws+PZs7l
CokJYB9i9wuS50Ht9u6fnsDudaD/nhwBL/PIp+Rjxy78Eci88Vd6kdnDvpjf0AlI
WipUWS5Jo+s8yUj1WsAatwmCTH0OqNxJfFvyoX/Y678XVQk/VSz3RpbNfYrbMB8K
FR4ivgEWWSUCcIFfJ354ISHJtPL3LLo7opbkgFVAr+klzYtxkYZO2BGtSV9Ae/6c
y7WcbQeehMXgsfSiBCm9DHqSjfxM/FGvpAHlGU4IbbluXYF9Px929ty+4JaqTc9y
4B2UnjmVBhIcV4sufKskpI4ctyUliKJJKPS/9H90XGapIp7Qi7zBCi79Gwf96D+h
Fnj2yIp9GRcbHFcf6tN8el1g7NWwdXffl9JUicPwycoczbBRYa0I6uUJqh2voA72
Ev/WbQcmuyKXK/ZCTx787MfQanZpv2i4KYYM8wqWXmDrgpuaChlHyMXv4jOxsRuI
Mww9yYMePEYJ40Pdh97A5T09UqF5MscEdcgYPAblDbNJ8ldHgzZXan0TTZ5vSM9a
1Tnddij+8Q0YBQmUuUXNxFDk3yT7uThTkh++10HyxEqpySFt/cHnx6ZE2YQ7GrYU
CirNtDdRH3qlTGjDIoRBSC+PIG41QHDyXW+DXZ3U85oDd1u7jSoVW6J+sLiCgMbD
0BrrgJqhVZn6qpAMx6wbPTQPXeJQX0onG51vjQJNWXWnun2N2h+UAUsCgKMRgiuY
bVs7dN9wpFnJooPbMozuyFCYGOQ43uWb7ViT0brptzxWAONXFJVtAPYEiNcDe61R
GQsSpubGK/RBH6c+65ZGkWYV20P1yDBLwtEETffN7xO06Jhjcem/57Ys4ew6FmKk
x5vapRHrU6HBHKL8hRoQ82waZbijg+UmXGAtonuhv6DbNo7BPKDrajmmwefD9JOS
Cf1gVqLGcih15JMxRttHA2bIEMwr89+kp9DOXvrxHWs8ico35vajK5s2fzXaqNPs
TP/1Umxjrrl4c5buNSOvUWVK/4bfDp5kr0GUGODFG0QdTY7TVQg9HVnY9Hf1MxJb
Ba6i1BMmpjeItG0HO8Uc50aUdHvhaxwBRd+x4T8prkjT6kJaGnZwf9+6bSOlSF//
+WoojDs9OgHjpAvtJwuyxbkIeoa7178Gn0NozbiTFOSW0nVBcuJY5VAfsD+IqPgU
y2koyftj0kZxdeaLke2IpiCvYORHYnel/0B20yby85y1Mm51Z+I5UTOO4BMsn5UB
S9b6QsWMEJ43nCi/JFOttsIuXf92IFxw0QWByTha+H8NTolN6MWgJLB0NTTKTyh7
fY5E9Vr/s9+pSggWwWztnVrSD6IZM54I6RK/j76xeIHsgD2xSTPx8EuYg5vqUyzj
5K5/YQSVWzWdlgQ/chW/zVYCt+IhTabmRnJwU9bEelifbi7hnkQucngudfEXa8Oz
lAO13BO4Tj25j1uIAcG9gDV4MyHLNIzZb8IAZfDz33Jpig1FVL/k70NJEvJk+Fbl
Aotw7GOs0OL34+jHtK8NbJmtOo0FCzkfx2qnJhk914oC27fX6G5FRIOHLnYNbO57
BH0WQcFlYCv0jmkHQFrTimka/dRIndsMLWCw/wypbduhFzDWwIPEwYyPLtKXl9aM
A2s73BX9eg4KlHlcXK3CgOdUBgvKTRYxogruYNdJjaeHawBXFlwSLvUGhG7KsmcL
0AID7XzD3nEEWoXGhpGGkT8traQhf4HHBIVfKcEuxfdttV5rQ2NKay5lDl/ZfBhz
AqKcLxGS/G0+Vur5oL7WcuuPjw9/+EqZIDEd+gr0r3TjZzs/cud2bavnii47f8pd
iHSiVpiY7qGuwIEgNsCQp4+TBKXfG5TvO0NItDYvM3n3UjarKK6t3ew1mqQSdiT9
ECvr/YV1WQ1uGi/S+Ns3yxUwyem4yKTRFFw5yivlPJ6JKf9eS+4b6ZBjWUiuWskq
vqyeiatCXg1NKNTK840AXF4xsFygUuU0ayjUXRRb0gqwjHeXou7YZlqqxT0HsH8Q
ED2II3m688pJrC2lI5hAZBOmsNhJ5OCpNpY1d1q29qKFskwkzKEYQR/+mB1n5snl
g7l4jqcVHakCtNoSi2Uq+H9NZiW/SkqlMf3H0zm/gC7oDuBlkcDx7RJJz6RJQAAE
v7psv495+ESnY5z74oVgTHELAlrRZqRgZwJKklmbUkYsVq7GqPm1WF1Us5Z/5bv4
6a9tuOC6+aAItiUPne9AphCZ5YDLBlmfd01p4qv5M695fums0zqrJ5FzT+e2x6V8
FKBOTsZEQBTGucasr9D7hw0+DUx9oYnRjkkMVta1mm9OEqj9MHb1ASBrTS2hAUV8
y8NhsA7npAoaDPvtKlE6EtUZPaIGcpfyNTJwskI+lhswDHB31Hd3yVT5pAbDtn4/
MQPrIgY2vS6BvnobqP07CAhAwG4upWHwX8DmXtKOC6TNHOupfirT45+pdWkt+F+U
3OneUmWG4d0iQeS8d8Ol/SgLBAFB3A/edhHk6Uas1nsCifSo2Dv9O4CxbfLhEnwj
AeyPwh7lNImKaU8cW96DzqX7J76fdxiQ+5x6rGGf+UH4X9zayH5yfPEYc4v7y+9M
FGwajIF103L3UBWowNAwkaqsYoJBIsH08BGFXP3XU6GmTOgUWPAOU/ndvZLyY4z9
dZpmITqxb9i/+I4Bj/6xUAJMTqBS4cfbbxBiuEI4pXNy8UWGU8FO1T8VGY584dsT
5gB5lFcueH7JCS4GCbcZKT3R2AHHdSNKYGb5fQ8gmjlI36YtBJa/ZvZLzZc4hM05
c2dn+5TJORb5GUNSroOfyZ4XzMEvwLQU2bBRynx3Kn9j4lWsOKafi3PU8CL7HJwc
ngN8cq8/CTvIYh/czvjE9/WIHIpJLSeqWdfuyHKDA+joyOTIv7mR/gx2my5a81oO
E+on5ynttnpS8kGCN1KdaiOvpPGLIqL27i8T0WoJN0coluzGq53uilTuNZHSz/Gq
5KNXDlOm2bnt3PmVTOqVD8UYrMuuWM7Xm14pM1R0JNj37vTSAzYzEmEtVNjaKg39
j+mXhFHobH68OgkbPgQ8xNuAlvPYg6LIRW48CRmPAcKV2xYWJ8ixJIpfRuHrUsVN
nn30NOOW6OQjmjJfxVcybW6jGUvjbx/5Tbmd2nkK/slJV1WASB0NfTI8BbTArA+K
ppu02a3ty5TKRGMEM3c7ycsYP1IZNC/RiV1abNI+LpPRe74rJ+oeX4F9H/Mjg4E2
8nw/t/LMwSJCE2SkA2L0FUmbmp4efQHzY09t9Vx2ph+FlaBolgmZrgH0G0YOGyWh
XhIFT3m1tQPfLF9lZmPWbyO16zlFx/bPoIIiZi6O+dJRdmxb1UlAHzHfqudnqk8o
dggD/0kZcAnIlQb66OOecJ+zsA6UaTzFwm8gdMlJ1TflJEYOResSwRvWbttYJZ0k
BCLKeAraIuImZ07LxbWaya+oMvxSnIDI20HPDbk2zouj8PPFyJxLs+u67a6Zejy4
fjiLZlQXwvgVL4SfvhOlIw4pdaF4Q4w9+ft36Ib0eBoIJdL+pD/bfq6+5N8nRKmg
ZfvZWcGLSpNj0d3mhQS8hAM2h0H3qtK/yQbbtm7wjjNq/NblpP9aReO5lrbCKMuF
MMP3NdXK48Yar0e33NjY8dMTWcH6/JxLVgITN/Dg19LzeQpSni3cqwmX879JFMqD
jl9w5G9fDrKoF6OJA+9vCYDgnkNaRKvzYKgV+zajNoS2YDGjE+nQ8JqwXZVTPNRb
1SFKQiCQNMsZHmXbB7gPItNQnl4BzGYW+8JA/X//Xh3TqgKhL3orz0fhdc25Nyyh
ix5DgPtzmEmSXKuZZGPOcrNJmpI6jokmzxrIVquxAa0tvgLZxGXPFvCuT180TCey
Dq3SpxT+Y2HSid6Ne5DvNsP0MBkrCMd+TCiToz0u2iVIYkCyfP9nh92iWUJG/2kn
tUJTaqo7HqSGmFHes7Ool/xPgLrn9OP2+YOU1wsx9jTupiS7txCcZYw7OGtECYNo
QWadjKD7GS4pVV6AUu9GluSSNl3xF+hVVsRUPrW+Ohv/FNAgS9dypzIElXJnX9vJ
+SdmATgsXeo719WNkmp0ayp7drWOgcJMVbJVi+4bz2sPkf4GiVruxiD7kijrAC/2
U1YoDEgjkyuCjyjTynwhWCYM3x5hM6Fv0QZTrzkubFDYcB5brGhSizWcVLEVmdvz
RbUZpqB58INpTKGIxadEPatxUOu23h0PeqI4L09Jm8CcIpWUgCwRA1dkX7skUvIE
AFDYJt9yzXXCQ79ahd7JPC/3cLu73osnkt033oLy9dP7zqbOrGlhrXQdL4/DTDO6
zYchiVLc5jdhTkZdU7TdPSI82o4AuB2k389T6eBNTUXFzpaEfOYwZSqMOll6wgVY
1qBGffHw3OipGMEPc5PM8EjC2BmI2AY7OjMdw+FD4Iwzxyx6SYb8PzvApnvke0gS
udv7vh6ft3g9YOLW/xaRlfyiICESrjhdsyAINopUXMsvfqcJYwc0l9oBdvv7DK4Q
jIWQSm9xr7fCVWdoxdG1+pRm6vNZwglpQmSS+J0vBL1VlgO5P2oX93nUhDq2JppW
obwjN2I6tdd8WB3ixba9v0dinHq44kOUaJUpJSmaUqhiIPCupgE2bMuxec8Bz1bN
fAAC2jyloGb0HpmrVcwJncG6Fx0xtThTPP1GxHJYOQ6KFPBtCIeZTiMBFv6UhwRY
6FZuZow0mNpl3uSAvAag7eHZS1n0+xaZm/iELv01xRGZCk/s3RDDAgwPZRJTX5xL
trtY4SdhouS58t6nFyalb4ilq0rlFyGHZJJDttbbhamh/s1VSHjITpzvWY5KuHWo
vCeJTBLHlTqPDcBI9icNk+bd7zDscOt7dmp+DVdFtYMAaUrFSXjQrObOQEHo9d/7
528/zvCW+/dZzBoVl2UEWlHG7Gz+iN/Nk0xR6CfG3mIJ2zhtUjAE9V0ZpW0AqxFD
6z+xcO6mNiBG8iLmeVeJMDKlwgtMKhFqwnCwx+mBF5c9KoJ/Z4L4PT7NUiiuqRil
KSXdbFB06JHYDGKWgxBQbsGYzN4ikEANDCd0SrEI7tg7n0OM32lPnLUJZZ627esN
BEDiPBRUGuz+esX4l+2p1Zonc3EEaqI4bcTgbYzt7TfNvRuiqGXqEe5v9mI+KOtv
6jQL9Acx8EQZpse1f+tvKyTXT1fshSghLc8ZmLaHDE68Tzwydo5CN2QPJ+RPso8n
UHpi1XM0NCiWojruW95BliCoZO9qsqcN/gj8lhaWZgFXvhp/fcmjxnZkPevg3CJ/
gSrIPECpD1M9cmC/1hviG+X1BCIW45G/jdSeLSQqvE2UK+2TEayEra+JHlOFkTTL
MWZxBZ+fnYps8bwUroxStxPHUl/bzs2kbcHuyMiCMDY1JlCPWWUtvcfAP2URDaNU
n4AjiReT7aEJyyo8mLvD4oKw8ltY8y6DNWOSjG8+b/lBfkjxbo+betakgN/AttmK
iEEFTMLbSZnOeadhz+6592q4lIoXMobIiQ6kb4dhHfKZ92ncLUscWI+l4EZI75t9
fMaD8dEioNVbw9wAln/3NBosERspmcOTKejiK9iD/tVFDDdDNKAFRROtx6h/ziZW
FWZS+dLuj8l531dC2FwU8cfNRV57f2rvV/SW46NqrKYRFo8j5tpro8K/vz49iOYq
Bj45d0WiwPVySQ1HMW2PibpNh5PSCn6ADiBpEj90buJx0Z6SWcxhRoGxFA4RkKwf
u43ASpWa1MsjzxLeysgiOpQvAQ1+SggmJ3OhZgCL7hsdYohIbXRQR5R+e4Lzs/80
1a9hvNXggg+APsYcq0rPdwMd/wxYpggxDNCoLHgiMKPzrfgkLONdqrzCu0T3GY9u
R13usPBnhDGxLsazVfuRkgGA72E3Ar8ijk6aLOXd8/+YS9Cj3nZIoui+bx9GhziZ
6p0arS8zGAKSapcGNhokX3xYnQyzM+OKs0bglQF7J+JDnv1RToU1BnzEcDidSQ8s
i5MoXCVEyvG5CBy+vcHchC6ge36qHQpCXLE7h96Oe5fMbPdfF+ZifGuhmOymKtYt
yRDaI9D/TkUn/YIQk8lDksLRNssxxvjWQANaZf7gV4zPPTgPw3lVqpxXB8GMHGyb
qWHVNPYVFjhvtt8VaOGLbCvbpz6kt/jadtg08I0EaWV+PHoPViW62Kbdrr4aUdz3
fiVHVHRuy4F8CwvDahiTFwrlDteXHW7xG/NzsTXDOnu5UI2Ul4W1vwv8ccOorebQ
X5Yd+ncuBG7SdBUVPL1xg/3BVf6FN56+KBsT8KZQLKseBGqE5cd60mu6YXSCr84G
6ShuMob0VRsDv3oM9Q4MhAkHtIRMGDbpmQQEpbjzjgSVGbOIA6Vnjie8LdI7DN3f
X7utsbWr55mGdxXb/tiiGbOM6RYCLwDK4krdNUZyKvDBMu7PjUpy6LFI8v0t/3Es
aQL0KHn8hYGecKledk6FWCXAw3JW0hSKvAfkp+kvWLxTSH3WPWOyhVqztaJMyAAW
J7HskrFZf7Vj4lalWQe/lQxyyJYhsY0PilYr5HOt6N67fd5gbuuVYbS+httFtOYN
YhuPvYkp0cPYQ53newwOUfbCo72pyS/p0mT8jJ5C1/i/KL6WqvFAqnhO4T+iAyxA
5PwNAgnETteDekVxdbOz7Y3GzE+GCR9QkU8TcEZNOSEKw7ZbnWG+dKM8iqsyC9Tc
5YQFZ7xvuMLeTThhGkbYbEnC+X5sXDm84LoyMpv2EGr8yBvS9gBxp2Ca3dI87QUZ
6EL8cjzXBEKz79pQmdCrQ6mxSd/N+gNRisR7hf3PSCjt4cK5oitaRAuw//BlVkh6
WCTMynfE8B+dgMvJbDtWIL79eDEjQGaWcaQzPRmK4bhPZBxLPiLcKRoqbOHTG1G0
5Tj8cgSmrpnbkp7/x68HeJzM77XRIXic4ytM6p5CskP+t/XfqnWueBKEbxy39WEh
f31q1m9ZAWs3LtDUVj6+aoVN5V6UgJkF9jwzCeHZ83nDrfmDC5xdBVlYO+FbN0uV
kJNb+BU6PxTgX6j/effwqpPypmVsWAGwIodPqQ6bnxPj/iPnXteWZvEtDDKG5Bcy
LS3/rZIJtdQ/g+d3dMmDxEWg+ngpQYIKpGDXFuj2Udpeokl0ca2b8fwFVOAuW342
lpuAZchyDXU/iBIgyGQ1sp98ADX+Qh+Dqm4Mam8TOZe8UtBe5LVQzXWYfftsLnYc
21pu+giLGy6oPIIIBkyZ9Ag21rKODRrMA83LMpUzr5BMipZbnLhlFdoU7xhN7Fm+
gOg6dSm/JpUU3yqsLh1XNq2Vst7GpuNkikyAthVDR6A2lMgbHySATdQLnwG092iD
HR9nOhWN4+Yp4JybHIY66PnPv5F32naYCWcut/jtMyyt0WgNp8Np3TNsypdVevv9
v1g6MyAEjUvwnAc5QrbfNaiXgESprBxV6SRG6KLt0+MkcAwuZ+41oBeT/FAuZhAi
YmvsOtcZgql2MY+6lX9Zczxo7Rm7dqIo6whxeA1Yx7kDE0brxjGvsu9lZGZ+mUx+
G3Q1MbI0yhliabn0klPCpfkfbhuVFTio1ongh9zPrt1O36j+QneXgudJ3syph4kV
CqzpJuToQWB4JJ4uY1sgt4d9n7HjL0drrPYCHmhqhXXbvPU6tb+/4DJvLX2a9DVl
zXp9jFcxIO4eyrgh+tW/xjY+1BX3McBFXE3A/Ema0stvYNPW26AaR2ITasApQ0L8
862kLpDZVwd5YYuQcx+KBd99KLOcqV2W5rdcNZ2fHO7P2Xfdm45huEGZbpB2YARb
8evRsAkKoTVvB4JWNxXGAI+pKSmhroMY/7cFReJ/xIK/4y3tZbm7JJ4UtKY3wZvj
ceZD3TK9++SgO8+I0+o5QGPosbu4IaC89o97KZz23ppX5rphmgPGtqR3wyN1OBhK
vQGOijZbOcNsX7qKo8Csg23dahFDhYEYvD21BiSQZqjfpaxSPfFmeICFMn/Ynfjh
HsVmIM8SB9MZUTbsaThDh748d1nJy3R5dhSnaoqSpJcbRzj7rB7cS5VsfwAtumib
1a9eBOmjMrlMNlFGtgoL+Qb5SdrlX8ygguWOZvsezq577xo+2uQEjHDTxmmToR/5
RDwlXmCqAsYWSHnbq3IUHx1tEcf/LrlB3I0Gmjq0crfViz83Ldp8OGhnQSnuorfG
7Ao0rpCEJEn60xnT0mZesQ665T7sboMQkjdM2GlI6mwkn7MX0ez41a1DntZSjBHM
rVaNXqtnsZvBfXqy9BVnXCI488tDlhZqgJ5d6L4+0VxIk1m0sTMDHg3++Yi/A5W0
hZd3mtIfdMHISCPUzUtE9ydM16y6EyIVUtcntwxjN5yHWsBpr1IeTEi0NtDmRQ58
E03uFuEiY4/lsjwprbAfG5wHE7+OdyK6xqQalInxJy3n2ueOy/mHfPR4EEEZhNz3
XSxLygay0j9ji4/eRrBgyKjEUIg8MSsFBGvQnzQjiiLLIy2M7+//fajj6qUQDipF
0qO0vDvfkTRENVhRv6NYeW6w2u7CJBCDvdznUMAFwWTuTKtLpe/zilQ3VHVNeEV/
8jC2u84PqUipxdcyo4Yw8fcFVAHtkEb8AHvP0fgdndZ+mBVXDIjtZw/utg1ly+/5
ky3UO269xNpP3EUxKqAvsroir+pt2FHEWGk1414z2PikJDcJauDtkBVF3eEnAfgb
rVBwSaGOw4E5IVIQbBadBDSu4frNDAOme2NzakZyWZPbJagRnggJ7PSSjTTNkypB
FS1jW2kRPL7RXQY73tiolHrr3q53114ld3e2aa1U/rGGVVs8wiAViQ/AI97g2uMG
VQDX0YrOsA0bNw1bQzyTB3rOIU7OvYj3N16HGFtdTcOq9WnQJV7jANPbFWNTivfU
zJgbG5SICt6I0s42hOSxFNfNX7mO4zY/vip7vfGMVv4eVYpxbZGoWxB4BbEDnAe0
0X4x1OPmTDKQ/DOuv/3Ki8aT/ebJlMV43HjXKujuvlmSNWSc+LsSynSV9u5uA00k
D0anjPvuUaHAg6B6+jHM3Z7Xiu3Ww/Vm5jQ/c3Oty8l1w+NqJY1t99j88WmMszD9
Ial18eIryHcl8HCfZ9muQDkVWSzxvzAEGfTXJouTGebJLR8NVXxGR9h7pTspKRfz
iPfiTY9OQMaGM3gl/duAzhb0rJNp6+eSUTnXxd791qCs+fOHM6bc+y505ZEYH/uA
B+C+rB82GPCbLPOHvlflIJZT6zD9BgCUTWRSjG0+9gsV0FX3v8mYhTfVtCGEGBZ4
bAtlFr875lzovRE0Tckt+DHj6hTU7rCRC4to0IwDGzpqCXffpvE50tpsTOHC3qv6
aXX75N66+wLIyjSFu+N+VOqb61ZhA/fvRp6716GcUucaWkPpW1S0PLrhaRBqz5vn
AlpZliu2jd7+gBd6S+AI7ioHMGJ71l5l+VaB2/sG54a3elcgxWz7nNBwTceTJaF/
nMw5qCo5apH6mEMxjlritt71YI6htQQLcjgOJk7MZx92BGABUFQFdkqbYLB+j/Q8
H83fOhRHPEo5hvC+HNYNUb89HlRBjNpGCdxLGH8Ib7Wvyu+Uz40rCpPTIew54ITG
JljQsyR+lqeHBYQc5j5wrhdiukg1Hw5Ux6vGEtOoJfbcqWYFFf3Nxp5TpWO4+sQp
bQZ76pjzRt/+Jyee6oLT1t16UW0tWi7JznpEVWrlHf4hZfTprvfOsBA5WQEbPFOF
HMdIBcVvm+46oTJ2igrc15VzjHuCS17p4EMDc6HLju8VSQXIRhubQWp+ZlGaGEGB
SNM5saA+IGwv5sJi+wvZDfmmNEa/8HxALeo3zr4AvQLDZ9OZfwGTxb2SPrVSmeMy
mOivpCLFCyQU0YLvxo7CFsoYIIteE5VXAGRc7E00KuzkSaeQEwCbnCFv8w83EWbV
vfE1aWhRwL4rGT55Yc4rD6ZffaDTeXBa5Ggw5FWAGVMBoBHu5YXYOxC+2n2QtU2E
IAoJEi8mNrtiivDnSet6Eh+6ozqB4jcn8Mj0prwNFp1RpoJ0PdtkD0NQg0DMYN/e
foTm507rP6xpv5PbiW9OYbJRsdQSYqDyNfZvzSFnDWM16K21CdKAiALH9TFuLomj
YJZeV2WQvJXnd7GSJYHLBRVFBjD1s1CcooTVzJFmrXwp60xz1gNishiNDDLkgqn6
i6PGUbA7zVgfEmzBq8grR6hP4V+02Qd6JB5AYCFqBdI/5fxt/RpNVhWsPST/Thhd
KCO8zQNnpxapg3VOx+N+dEn64IFz1bymxc5b2z6sOEb3P/cHYlNQ1+pBvN/HgaPN
JxtYA2oKLHAUDksFWoDm5KO3oZzyXBkr59sOU30IVAy46ah0Fq0liGuDsIPwd8qM
8mPOnO72C/qWRvxuXH9G0l80NQABKFnCL87GdLRZFlFJxxxnBG+tBGPTxwqomEKj
dUHXB9OJmZDPXg8IlYc+JdHCDE+w+Z+PsZue7jZhClfdhCa6TlWZm4Av9utMfHIj
XhnIUh6vPQ9YiEAxKgEFWG5o0RaCkzk/rlo+MNru1qRCTMS87MzLJ4ZRvq9VABTV
gItH0uus3lHM/l/KgPKvKib4IuZtC1+J34iaCaIDjHEIkUNZEH1DfSSnQxx7TYiG
35ZlmwbzXZGO59qaGAIfCV40t1pBqwMjzjVp02oWIsqQRyWHbHO94S1+F8IMOBHk
Ox1PG/m+5QtMobxQ2vP5m62tLT9oI9QIQ6CNVhvHMFT9SC5KheLymC4WJOfxP7c8
lxdYfY9xGZUaVF57Pa3yGfiQGem1sVql2N+pF01m5LrltWp0XRUmzDEunxazjZdc
jk2gKAJ6LzJtTgsICYwBlWIGCCiRQRHPUJgB6pmRRe4S8Qd7m5zln1iigjwLo92p
CtPWXRqXpWfzihvtNqP/wM5A1GeyF2O/FGJq4LChfz/zfuOxKPkgU53hAmnet2dn
FMdaxj0bzlaHbQOFqdO6Cn5YIx4utjm01wZJO0VcBD5mX438hX2zPBwwmM/fNwLW
cvgfK0aaUdwrXXWcnY+79xBixSi72v/oPs7JvRLF35NWr6UpXDLdivO8uRBuu53I
c3L3QJfWiCCvMKm30mDyiep+IA7t0G7+CSFVRGacCDDM5R1/QRuMpp6kq88OoAXw
Exk/JbHkZC7zzu/SQCwUqkcIQNkKZBophQvaKoO8eOPIRn6FMuqG/pseRuzFe1AL
IqsbOTI+c2HDpuuJyjC6ZZoT1OWFCrwxwf/X5wDndrdYi22c291xia9byD5sxR2r
SbyFtKmVhz70yu1ENDxfcK4BCNbvGA+jTaEhVcJBBGzqk3VTPPJdpBq7pegNBKNl
2uQK4WHlv1gOI+eQmr9YiVbxkSlcXVGEHNcl2RIw1FnCHX0v5nmr0UmRWg9VhYIp
1lyV2LbUKTeJJA/kAwA/mdI43/dnvjjzYA8hMycOoLqwmlFf3pMdJdqj77NAN8MZ
T2yOAvvm9eASfltAonxVBg2rcPu1+Oz5Bc6dzafyNZPlLL1PSqM+ytQQyWm+Qaf5
3QdDr8122ukNABYCfgQvgXPjBxyXApzq6ohuNZEnaO7hlceydoBoqDr8D4GEytYI
xJhh1+74+6Auj+cI+luA/lTZcBfPc8gE/rdkvQduSd1nirWDVerlY0eMZ0021Qir
pTvpXespNsLkFxMtTYz40XeaS+Uv9zzNLLxZl9o8eDRAx4yqmVmMvOxxzTmqoBAj
dc7YJ6FmRMbh/NMhcfwk4AHYUcmZHpFDg48ZZBVt9oseLypnzv+JP5D16K8ORrFM
QeR5EBN+k4JkkJPuApYbHYMy2O+p+gcpJnsd4dAWgz+CZ7ETXOWRPo7ru8YAVhHS
fSmYIWFMB9syT1ohHDA1Kk7blU5s7q5zhjl4ngShF15dARHDEWI8ykrTyxX0hLL+
GEP7FM6/TDkkXL/3ClNmjWpNumTG8ZO0W++NeMutx5+HovOzO8KtemTL4/u1dq4T
lxX2xBBzkpgVE4/F6Y0nd/yuRIjI/mgJXYhITaTy8S9fKaVwpbU5G3k+KJDiarFz
R093RRHLufYoxfiMvlUNQpFYzSGDUWY9JH9pcdOmSH+wBOkFhoYmO2SUCVBL8Izs
B0rglQv4pRIcT/0SLT8avIv9FpMv/r9JxDOD2lWTW6QoNwVftnTrpieHeOEVgo/p
hNIpj94T+xloyBHlS1GOGp562rQnI7dcIDLJK3gz4p/jizrAuD2+HA3GbPzTEaCU
897Hd83FCnXp9Z8othQebjKHBO9O7G0BkYarIOYcwlbxTVYiOAlAAVIeff0fGi2v
ZDGE37MOHdfLRTDMFJL4FG+kHgEbNQc1mhBL+rZiEBcbbTAa1SAUAytP7FyRKeEH
jH6VtiJKEDdsQ/wjGW6f21c8YS0C+j2ueXfJ/9TTLEg/2IbXWh8nxvWGwyqCQApc
pCsehsEKnWeeVOLCk2RhcD2MIEnOu32PVexlxL1NDYTbH5Z5FLQOPwAXE781rbI+
p/JaYwgw3he9p25VzfRWdYjtkaEdb5RQZzyiqBfL0tvCDpYlwF/yO7W5PhlVCRx9
kTa/+pA6MzGu4h0utDUQnfgsIhHT+4+hdOmdkmImjFYJ6qt5i2ESRcUADysYieGk
yzFLT/33ZC1cNI/oGg9N3/2Hysuzy26uU17zRhuHvkPomwv0SF2iVjVQ99Eb9pFy
ubefOOGNvMuxc01zziLg++Ml1HqH+XwW5RH/At461bqMIz61WATL7EyRSrxQzSKg
ZfXjaRMKekoPsIdQcDt6wGeTYy67OTMxDFCAF3CfKz2/4BXTGxYwAlvQQJRpreHz
nOhcdF+FGKtMLYzwXxQZlRAA/yjdkf34WXAgbdghhUvf7yt6s/AAN3izO/+p9WOA
+KDGTTTqV8yeQZv0LRuPeR6EzMIiNqgE8OtIbkwPms54qVQ+Z5uE/VY2FZb9DjWH
ptl0bz8W5GfXBEEjtofaOuG0H2Gj4FiFeUEHd+mTg+6N+WvMaEvXMWxEbE05yK/q
SQUqm+nJMGvQAmGXJAGoo4aa8hqxO1sAAALRvP1WAaoytwZgCpv/ut/B5YaHYRHL
6be3PS+Y5FmYKfNsDwWEEVTGoDOp+Bnm5RGkeJkCXHUTKc0r3ZXMFel56EAfAebd
OlqeNb+fFJ26wS+kwHWtlE3iWrFL8z4dUGfGEPgdRJSeDVu+K6DkSmWB9ZnbXR6u
uR6YyFxN9SL4OsVuScw5dkxlvIksLS57xN+8/xDWvdrpjgu7cboVUbEbXRE3G4a0
Z6TJaDFdHPa6zw0BT68fVPgG2glUBY4YSFzX+KI3aTl1d9BsbX5YpdUwSfIX6phJ
vu0hZYyY9niKtO11YW9lNj0zqU+YWvIZ1lvO9JUJCaQgLcBBl2lM1IAhU2Z8b+Mi
pNP3UcthXugQFmARXz81aeZrXyUTbVbhr/Lcw3mBxWsBmtKn9apEoJ95MeZVo91X
XOmIcyHNVCgtvX6qsNt/hsHvFwA5ZNhRf2opIyeM4l5bk4c8i3S4nTz2H1EhclRY
rHFZZ3E5VpAg4ERnJcP3B9ukhSJJCz3W12XsLfK54Djaerz6PKoe0FyAH+jEvleo
Vpn7kKKuGjsjqNFilwANV79YouLr+X3WYs9eCJ5P9kcZAul8ThkTPNue+MQ9iKHR
zp6XP6oDaaTFNH4pJWlQRy8pukcZWeLPUyFBJmo3XXyt9/+hUVlcxQEBag5ZKSuk
15bfT8UAdCNe72gxHSJVQQOq3fEpGln01Tw/p1dmYp2rO/GBwWuB92t5vn5Amfk8
cfXQQ+jHB9NmVSsqdBFYOihvBkZI1haXgNrNHn6vWBe6mtqUjYs5aSd4uqSFYVnb
OBdm4mG82sO9LmqzosPU9wocR+oVzs0kIfVlOT7aFK3mLmcsrZcftoU3BIN3C4Ia
Sb8rbXnJGIfNHSz3vK6oKZpASoBLjX9K7wgBpQeU+3SEwus013JDeMRbJulRGyFC
uBf/lhRJlv9HMh2Xk79wiEcPwa6T9HAOfXrrJrbfV/deoIoTJYSgJJ17TvSVgEBY
P41vgHPv8pFdCj91ojgxo0mr1fDZRV1O5tcpu6ueLEzYQwj7hcqppt+m9myECo0s
M0RpV5IJQIfPl5hrrituC6nno1n2J2kzjv1t6DGPMI2pm2ZNBhRklAP9JC41tIdj
pXulkKS9q2hP+Isn3zyEalKPXygNT7H3wZTXFmAkEmg4dAP7LmeTAnONGN0gJdKn
qEd87Zx7okUq7aZmUOu+U+LXn8ifRUIOeI2xTDSu6YEur+AnC/vC8qIXJqAmuI4j
gmh6EsYY2l6A4XJo4FK7FeaM84JZqtDhcpgvGfjKZfYKx2Tz0C0Fuc438bqXfVr4
fPht9gL6cABX+NgDAd9n+V13N0vW9hwjRdl3rBlBccj1Ekr+BQvWl+UTrhNFMPQO
QSu7tJ/3ivrwcrk/jbB8ntFZb8Ub36iOa/ZaWnUgRjiqdVo/NcuLiyCi56vztjbK
mGkbmk4nqto5v6r95GqgPuIUMwHbbfDmGNHaQDpsqgQAI08zqzrPJsNLik5+O9vy
tI7ZjeEZiXiMKxiHUoA18AeufZyaW+5jC/0T5BG6QDcDjNl6IS3XYAXtMOX+gI9z
pA/Nn3h3G9ebz1+UtZr3jLjwG6I7jledaQBzgQd0RwiZi5foWhZmgsYARsYoHmE1
6xurv0QiBHm9fydoXFVyt3qFKWjblWYnXlAuOufd3oFPQUGx29qmtGA559yRw+WG
rb8C33PZKdKp5TyuzJpsbeeqvpedIO5AdxjBSDeLEo8vBIv1Q7L2EZPHk2MwcRwE
5Hn3sTke82t8I/YSdh6bt/L7mJ1uy3y2nj/l/Om4Nb16wLNmVdquAw2/3K9deqk/
zbxYcVuqO7FjoEWfTtkzZ73s2qPddfN47uYy6ARDVMrEhCmkrXmNIwv7w97lkF7x
0i+t2KaFI2LnKM0JiEex6p/tEFUkOAsLs/n4PYmri1LAZ6HwBPyiB5fcVHhf3H/L
z0tpcDf74TYYjItywgtOpqsEekpSMan6nElGZVpDTlkg9AkDSkBzacNzC2oqoARG
tiVEFuFYlVNIbyRNCOtDBf7y8R6al0AF1ALcx+RSuimX7GJ8P+heTYmNUJ6ot3l+
nNBdaOeTV7+9hHhSK8yM6HnIih8cV+PtpWCJcIFJo8qTVVlQQZQjUTL5estLdqun
bMiyu0EZywZNPiEHJSLf679YrKiMJluUuM18Jrjo+WQwY6iPptnNQtaT9C61FGog
jCOx0yzo5Mfhp4T6yquCJzhJW/zIbwcYEfFpGZr0bcMC+FBMcvObTKcw6ekD/8L8
+Uch+QfSOD4BovxFsvY0R88EIPS9eEKJGbJ0Icii0a93IoK9Svp/Q7cNlmkkhJOH
bHh027BTXYZMPCknYokAEB6X0FfMqe8R7AL6hRxC1/OBntZVGKgZt08ypKay6gYL
IwuciqyWrhPZ/opDrZ0EzXqTfYz/z9y6SGqO4czsUaojF6AUssv+k3rM3acGogsv
5g5ylKE0s5Hk7Rp+DSMq3bXsjjeoXzBuC9+10IAaDLFTfRqyNUOEv585uRDjRjP1
JaSMTzHsLxIbwJUp4USSIm//NM3gf/W3Ka2t4/lz6ZcduPCWUWm6jIQKZd8RsA9i
+UfjDJkqfUSQOshSn2n0cZCQF3fk2nOVAZDSgirPiYaNcaPcl8wK477XxmSD6Wsk
O9DpjgiQWV3gD1ltytGfvvnck+yFfsuEGLiym3CeWMJMZMhyZIeB7eZRT56hFMni
TCXq6vVXFErHQoBWzGUfVue2j/utuW4VzqcJIvd8TXLh1gQ+CMsq+ChX5N5XukPc
+qWgaW0DuLTDQbGwMFm/Ha1ZqyN2JNqAsqv4cbhl4oWaEv6vY2Ma7Sw3tlM891ub
7n7LRi7KtqPHTpA6kfPRZJWx4oexjJOJ+uWgrmHlUz5x13fkMzQr7zRiff0PNYrh
GKwqPlA689LuNTZUGJcUUAg2GpykGucacCJ3NAEnUJYc0E4ZqYNDPB3xpNlt98NZ
5QP5X3+F4MqgfPqouJ0IUXv7ZrGT2yVZWQ5Nv/SM3w1pieLu4C4yI/qU+0uSQWHW
WqV5pDz/nMGys5AYb13RE3Ue3YWFpWlIAYvjUinI83UAZDYtbl5AiapbKKy6uYZ8
UtEdvEBBbiR11UoLYBOz9+CUTwc2UWvPqCvjygm8AQgVVIKRi1Dux2i1n21cPnI+
UHQX2K8u7HFbd7zS5tdmg2R7M38OeB61ieKsrOUOC/t295ceDSW9dJdjUUNWogbX
QbQGVDARbFAp4N0PBuj7NwovlYJmZJd2OcYOnv1zA7ixR39t7OtH2Z2D7JDHHQi0
6cY7hiA3w9EglhfDjZgAS5+TkS4sJ9Rd4EtABBQdonW4Fa09b52Vh6+aeOgFLvjU
FyN/ZBexo3jGFKh2CeurrmkvnEMpYEkSiYA8okfoLepGJ/GdtUC4dBQaNvWawtTf
62P+YH6I8ea3tMS6ATMHs0GV7YCgtqgoIeJljsbW6lZRIUuAcQXpDjPRXAh16uvb
xlqCm9oHTMaxE3P7A+NCIHbstAKLxZdwt9B4i1vIxDcuhTcH7WMBxUTGIOgHHMq3
KCipQLY74A2wye4oFim0jE5GKQB6wa09eAtJwJuVj4w2ki1KhE9j60GJZ/O7RRrN
vb/VDa3SQwkG21neITliCnamnTgZakGtiISpIyTaPRRhjXNqcSpzF2d/53sKdJzX
1bQlzKlj/73QBu+RHDdLttILJPrXFLDMmAJlH9M4acqnuM9huaK4ssD4dw9qUKIB
6C6boxNFcn8DW15eddzbJyF9TAIOzzrPAeitdF3ZgTiwXJ3uVKOliFltHb1hU81h
JDM+WBGF2QW+S28XbGcDCht+kMkaaBBn7oi1UL6uPMOrjLVqa7QQtL4pb+3yySzt
YjD+14RhKNGN/ZIIQFZY+eFcd57lIm8wyz58DtPWDkMwo4ErL11I3L/dtSA/hmEr
pcAAt7U87CoRdLAMW5tM5bcEToaVdWbxQhkKm94T1Rrany/s7dI+uAVTGmRp3so8
uDC5MJ9SqV5m3EB8S6r2eEQng7Vc3ep4wUfMCmEsacZfmb+w22NsjHe6RVw/aaia
8PhBPHSCGB9peCvL5BIpj6Mz9oGQ+rb3ofPcn6Sgb9RV7wPwbkzRhh64SQxFCOx8
8VqLjD0gzg3jsAMeH3+6QI+JKawO5kyXpMh5Z6iWd8Vhpd5+eN0234QrdPWWdAHx
zexc+xgXN0kkK9Ks2vnYtFoJO4tySAw896n2iDkCl5kLV+GGEv0+pqBSOesrQP3c
Hg6hAfop3DUb9pechk8siQCb7cuhZKIMFSeM5a4//ES4vnpo9edFVMiTj9lzdoao
KHqf3V2aBbW60raPjM0HRqPN8kvzgj7+TmmvWS1Y/6z2oadez9MeWNuEFiGZCTIF
c7XvLRQV9PQJwCCU1SpVSOlXab4JC8WxHrQ1dZk04VBC7udstNbBTY2B2/M9J49A
ywRL3sdFkuVDU2bujp8mPzP526dKVPIFbQI4+6xs/Kae1quwWrOMGd9kbXkXkxkP
d4jjvqPzg1OYmTitny+Hb/2PJSKAabYaeLI3uCR9FP3Iuwv2TcVY76wpvbZNgwkg
fYJPlUy550WXvXgVWdNLzNXsJngdEm0NYxTwWOnvMJIudGG5cHybkDzoEtu8pmhW
mVQSap52eTXfNd2LRVOPMtnLrZ3Fs3UxAAU9QR6WitXQOQt5ZT3df+1tTSI+sYro
EwsS6D3XRloJhgi8Lz/ooRvjjFcOQySH0XdvE4elEmMsB4RQyg/xh+EZCm/RMo1A
70CcjKlpo7/mVMHQNnlYxhyF/P3+0NiKUXgv1aQwD8dUo7JBX+YTsZDVpkE2X5sk
1aAhsigqFwW8BgQ8AT1rowTV9O0iVAcxyfwVAZo/85Ci/AX/4tsfLDlUYSQ9L2i6
yniGsE2lbRv1J/vJ+MTHVCWJDM3THiOQlGKSsUwddYhWX0JpbKBYSMYt02ic9z+w
qhl0r5ragkpxn6RRVRTpEHXBL+z0chsvDkK4DhpXt0Dhhp3+5B/hfoHnrwRxvM76
oHXGdDdbhPxWT5pQyIgLedOn/ZCbTFBm1ockk7sHMPjZesI8WvfPdmmUPSM/Ku1a
nvnXofkxuK7ednBkDMsBrMtdNnJOAe3H8ZLTHtNoWxmzhsbZJU1YcsiChSjixUlz
78s3uKEd+yyceN4gwdajt0OLp10CwMEeMO87j3OjurQcpNKbtiLa1fxMiIDCIBOC
zUQpU1YFPtEx+6UUZMUg0FpdpVhTNb7wXZmQc04VLEfr0C5NIAPRXRvi6QtnEj1h
IdIKfOhwzVltdxWjx0w+3Be36uwHUA4KlPN/zxvmWa5c7/8o+/vrouqIFGqODBQY
HJNOJa8R7wQt96dwAi5Eep5FbduRw+ecM6/oA61gjiKJDxY7w6DlCRtEexVI3Qen
UJP0SAGNbylOjp07Mejk5mnZ8sUB/NeeP1rZCNVH+KwmW8BG0jsGiBkJR/IFD+SC
Kp/eADZkmqae0W21Dntn0+hgVIVGDI44rfi3MIrFZZgs+IWc/kV4koEyrp7ckJJL
kclyEGRyC5DvKt0ifQr4KtZhbjafcSIm3brpSox9/kLTq4M6HM/CvTEKMUq54y/W
vMcG2bwaEcRF46nG3LDuPDJMy7Dm9XUQCtHfH8c0BfiFAp+mlGYKBe/VJ3ptE0u1
or7y5uHn/KiyhxmwuQBFZkAL4k7P5WgYmmTN5PZeedhv1WFX2gwdyPLh+tLLK/fM
EZyvAiJl9NZK+lSQxs11SxKG2UYLL2o7p6R0Hf1ksUbgPFJpp9rCiuyC5nH6+eiv
Q8HXjAHlOVbN61Um9LtbhTD0AE9LNi7XKIrct2VHJelYKFOF39CvYe6Apgttw+fK
nAnXhF0+c3VIvgkgt8EIS1aLeO0UQsIcTZ1K4lg3P/osJRNMEYfsBDHTF1RY+fi3
GwTa+QlN5Bejk5aHdmnM1ZhYpq6GlbE5F53/R1H9evZgqnJhW8C1+e1vsclyxza9
csEgTar/rHcS1DiDQhDdGLIrLKgv7Pe1K/sYpg7tgiqOq0y5unNje9VSjviZhLC5
838XGnEqd3G1tEyds/Y8+I86ELAgAK3YgijckjbcGeeNWWjyUKE7dedMjCw9KM+k
ryp1EDuA7hkTfdbkffnUDg6STzhQZRFhLAhNJW4BMrekXOssdavwhYryG7xN8d30
I3bRWK+McRAVwDs4xf31G27I/Jj27rBRF7OHSyhQ9OPSBhlD+wMV9BfyG96ibnag
nmaT19Klh/n+EPD/40t/6kuYApNZgGqlfaBSFJxOLgtlCHgNro6COyGNXQhASFh6
hxSbMqeVduy1twYcioaWq9lLn7cnQm2hQ32kaClR0ZV/2ulp/RmH3W7AvnR+pvlf
wmggdKJFHk+qTwbANdKznxjba4TWZAETECm7Z319DSfncgIVvBBv61wEQ/CLSVmD
SuTFU7macpzvpZstUPTqqayuUHSq2s3ln1l0aycA8+LcCtsMn2xmh6M0NySVh+2f
4nQgIhOobfwGKdlPgKxpR05HHsayhJ9h83j3Rh8cioekGFyBsEcMyk3OnPBac5FN
fO2D3Wbbm826dInjSZP7YWW4OaJg+z7ftO4/vGHzeYfLk2qXh28SfWTG1hou4IMo
L2LUhOcGxnpYKZhG88FEBsyRufEYRQSaFvUO6Z0QqgvkSFYpAiehbJc23jvCJe45
YK7c4+qvhwn/bGwTXdg8EOsAa4kXoGICCAoUKPT41+sEnfD94k37CX5bzKu/Bo0o
V+SB4Hm6Tsj+9IZnkgKWw5P8Rzog6M/qP+TXXyb5VaV4kMKxiev13vo1spYdv5GH
xALDIGIqaphVBIksapqJEB5XAqYUN8nvjxT/rV4Uolk2qMuw0Hyy1//tZx7mLU/r
/8q4DV+d+zp2tXUzroVu8tOSiQWLz26rpn+PzRfZRKFfegyfAlfkP5s0aOS5m+el
faBDwqGOc7lduvNhggHQIvS5KsyGHNxxSTtVYMVPrvphO5XGQ5tJyHKzMp/xxrFA
LJpjJOXnj1KcsoeM5bKcbukIO3DJcHmsUi9pvr2eL4o7GTX+AkIR8vFZmjrXTrUH
dvSvox2PbThyWt6HobZRcm9/qQNg54AX+bGC9aUlkF+HjL09MgFhS3/PIFd5AGKT
fUcPiKG/+5UFYxe/Mc3naz8Q3Ci0kmuBju/M2m83Dx/CRvQcAgrmjJvSt5giASD5
9MUqU6V3a1TRVqnkVhrmd30MyuNGRaEqgD36Ywlsp3b8sc960+Tw3vxCmo9GovgT
CXz/x9EuZfQ8oukr4K6mTUpDKaRU37FejUI3YO3wdJsR2x5ExLdTQw03WnpT/y8m
K7qZiyfSf/teLwahO9hbcdqUYSGR258MhIJgR1anKZxa5aNIaZkq0QRkf15RGBS+
43sOEtsPp+Q0i2OXqv2iIB/J46f8SX+uWB2vpGotdupDQz3PHy4BkiVKuVc+UGWY
9Bp+LmltxRdaoxTZCAe4Yc8+xN5gYOuKFGHMV654eTulpFQLpqUtoS7uAecYKR2+
RCEq3SPUtC2HzgBwZOkOsyNQUgY8NXxFmZ8RVi2CC+z40WBa8UuXn2mdcEXCCPjc
XCXUidj7QeNjaPufPgpj35KRVGnwcfaUvsZfLPwcCl9Y5Yft8qtxaOyJ81mPIOdL
gKTetRAUi1RbDx9zR20Fd0fkpOiPdnnJXjOutT14WdnhVHNOhemjoY1DLDCQSeJ7
8ifrzjOXyjUtuJzheXJnFaVHySsrCmlEuBNg7bRCKAcYh5Xf6y5K1YOtvEYInezy
iPCWusMykTh7hdCJO0UB/H3gInSwvL/lOUPmMImTi9BPLdbGRyGDYwukyRT530tp
4lH08aikyirLFEFUCg6Q2w6J4xzxMqFEwEonk9jHqgECnie2iRlEvfy9yL/RzFI0
yH/RgdEDFxPiMjxI71UCg6ajY0kjX7y9aJ3Qy/uE5tIfs7qc+aVo5vcuIkw0+5yT
IcLIysWUI5g7Xux0zsdZOvhL5jGAAoGUSB+rGcxtQcFLaopr+3F/xxCjKEGE0bj0
kyOpv/N18j2ZAu9/atAOmnWMfoiJ2zT1J46X9+M7+QAuDceu1Cq/0LxEIHlN98J9
pfQincdXpbWZjFFuYeKUbAdt5xsdLx3lsN1EJXZPFOlhDHOrJSlLmuDRVMl/m/fB
M3WKZHFHeaFLASY3Z5dMAflA/xwYikSEJF3FD5QwavxhKIjzAVp6rhe77lQTAZ7e
4LS/mUHG4XHYMwe04yOboMBARkvOk5uu2F10fpiwJz7M8siBec0JzQNDkSrGF01T
fBcvl2XJD8lDhhzSEoUKUgExXzLOlFdBKb0cIYG6pbehN7OyaiemAlkB98R3pqdy
DB2rZ9UgskorFy2U1K+HBZdoYvZnBYY0raXcxc1QP6qTn4wemYH5PDJCyiJV35EB
d7qGuufYcbdpUA9ffJSgb5kyQ4MMUJgTwLMWCoUpo6ed4yVT6IH5MmQrAcfq5bSJ
x71vcVY6f8MFc54Xz1SMpS3AslIORXG6yl/stMt8e2ioCC8VXxNFOn7LhOlDWTox
LI6pyYG83xN0cmo2NKj+v1jxmNVenBSBiLhUdqixPR3QKf4fjKWV4L7VtRk3Wl2x
iJcx7ZY+o+qX0/yVtuqzugpp1H162wUgkAvebEX0yW1AOoy03UAe+fkQ8SE3YUEv
NsI/oMr9JI/x9sMx/tYBnCCHCz7b7XotJ5vIJgnHY4CXxsJ715T61TX5zuIyhI1z
KdfTI7/WSwK5PiwkLwlKwOUMCqxjzi+rquh1tWC/ZZtNJikSMII4bD6wd/25Z9r7
Zfsl1tCM5+d/XqAT9x2jew2A6JiYimVYd1J2ZwFqwn3/cRB9TpBvdrF3cTxeFXZU
Z4uVRcGonPavcqu4Box5az2+4FELu/NE9e6NS6aKLpZOlOuCZaPXmbt+bKjKgOvK
5oQ4j9rFsV2fVlFP63UjzUb/la8nVEMvilmtyeoJHXnRb5z6inCkNWjFpI1QBLuW
uv1/dzo0kjMfjWwE0TvUJyaPhBhcDHMmqiOy0WEbBK2s3vno3162kcVcs54vzJyB
EtpqYj/a1GGLdmWt4GqJN8Vq8vhS0Y4sJIfkXBppbFerOsTkuqqyoN+dEymBz+Vx
cIM7I+Z89STYfBEub/nXV2eDKDqvT7rt359tB2F8H0CowJY6Wky6IMcumEIXyKGA
qYnCx9Dolqmpkpplkgyz4IvUTgyA8nYSVmnqA9deU67GZdsbLdU5O/8NyMCpOKsw
YE3QdnO2zX4Yx9LjwtbKwTIDEvgg5mOl8ak5iFwrEiaKjpsJ2J1qdD775Xz3mYJp
h+QylDhIoBtst2hOc6n1MbAvL0AhYxLlGFLzKz8V+s0VtYQ3C7ILTSO8F3PahGZ9
LSBEnALAFq+yBnMi0//1ZPS/kNG4SD/iyVs1WYXcK68tsoccftTVNqUsHfBCKvx6
oUOnUaQi1dC/AU/awfbCuy7lTimqA+hg3TAc+23i7qCfMhPNoopyg6J0bKVEhIHx
Lcc3uttqHkyFT81dZO4U0lt4hhFF5YksQs/NWUmZGmZ//TyM7EzJ3KUXp0j/zPtg
dVDQELjp4dCf1+b3Jp1ZGiXLAP9rQkZrffrOFHR99VqKcfkjPnT75LwAOECTEpNV
FHy7f8i0fCBAX9IUWFV3WJS+WzCcYspwP+rmcsdTfUw4Dkq+5f47/bCERwv9lGoH
olfjp0EBWOrqkHs2lr8cnOwt2SWMEoEeGv3PMxOrwLSrH8405pB8xHh2W8jj+6ca
e/XacBH2O+yMoMPSnYLi32zT/hjxwi72kKvIRCzppaMmmhWNjaEQOP5nouzHal2v
I65WCL35jgIp5Z75+rtJFEFdvfT0iSx3KBwV600dMPIIELR/Qbblx2YlqnBjwuX6
nrq6KFUdsmb3VGievKEFPQ9wgzG06HSVqqECmvxCbOaJXSv/y8HDGJB+Dh7tG7XA
XxE+GHFrhV53O8g7XCDxUpbfjpUBEeIKugIqD5ml4hcAKx0h0B2nka7nitTS+AG/
WtiIUn2lPl4suXN9bC2qfqHLJWkbWPKeuIZSwVf+gxkehYW2XIf605z4G4ULHoTL
45RApvyQonz6eUsBsFLvlZkvh1rGQaZgigHS63RdPnzZ54GIpFVn8y1o9H/wBOIO
m8PLnoxR1il4ILG/JmBzW1e3HWA3Zupts0AJvG0yJcLXQkgoYKJVAp/64EWGClTE
SxFfZyMv8YRFHrhoPdWJX5sW/qhEgN3uHFsMhXlwUmVyUcZNWPO/8uZV47ALsnCD
+s1aKEwuala681Rf9WUQN3RTComy/eMmeeHT3kyZik1a897m7999bVx9Uzzp799T
xqzjPKPcjeoof2Om1ttOKUrGDssj0GV1FUiC4yb5gOl6BeUQWXI6818w3VSA85rn
/uRLjchRBCm1cRiE3z4El+ai+DB37NPL7VrLsHwJDqaVQnQPceq9HBke9WGgnXNM
UmQfQArjnlngDJic+I4FN4cFyYu3NwkWq104/uT7dznESzMoMviH0caFO7iHOQEj
t0PJkO6fUDD/qerRP/01Q7xFzvgQP5YJjh1tvYByjoKe9xbchK5p+9C8p/Yvnu6K
X9QRYTylv3WvxpCIe1BV5X8D6dz7b3rc7ecVDDvMtStXWhULL8m2bQMgFbBXzpIF
33uqKj569zAhmqVWZhtmeijMZLcb+CgTy9xnd6wYMdeSLAcZCx80hgVUUHZiLZk1
tqUL2b9nlxaEknX/U1CivGtjz00m8IW34hvZCvCppx9eiWPzg8zF4iYaeSjJ8kvB
08pAruA0CpgurngMNnDqS5/N/Db6fx+dXB1nMkQiI4kZRww35toq59Fn5FyCzbFV
6AcThfKEW5IiZeD5zNTrcEn2L7yoDG2d/cEsMhDAVjAwRnHqCwgzPsWr7x+iTBIj
K588Q35Ruceiz4+X3y+r0tmseTkF2GiNNwD4e7D2rAoXFEV4+uqA26jrPVpUtSkZ
NR3n0/Y4rRz/7aHTUSX3dBNtA+RKuOvDdwStXUPBQL+1hZGeD+QeZfGUkUodWBhF
eEB4mnbziIhBmCusvbQN9pwbQBnZlhIrfVhhk3j21KUieqvi58hlcMvMYhMcND8u
exk8T28uU9gE1Qi8vEGSwkjVxAY8hoKtvrs5bWaBASGE/3vYLJpCXdLdGyfLA4A2
Zy6UgmpIYvUzNVdPPyKjHSmBWbyupEnKkeOy/6tfEFiMT07EysaVR/Zx8cH/J99+
oa/UgrMija2c/soT/9Q4nrTfeyq7YjdgHZl3mZ6Lpg5fujktyrKt2/ziTrscZvqs
g6U68CUck8r6FwpNzzfP3raELZDcoLzWf3PzcdmvcVU/mLvwtPYbLnp6i93kmNha
UzCb81wyW3mfnT2v+PPrwDu+MoDH2hWq3oTooQijbvz+zm+0Eln02/tHkrnvy8Me
y5K2ttdg9QkpA0ffav1OCQgFUPgeAFbW7M98PE36ONZ8WfROffKiu5xH+ELYZZK9
mXtJKGoy4fenslglBFB/ooq4dHikalYOY02TncosUDsrexTEb2/f+qm3MNZNU6fP
NZVj5A/MsFdbxmAe0CZUZIZZmPUvpg6BPcvibHHeyQPkCOCigLtjgfhXR2pz6YWv
L7JIvt9UELcblB3BmxvUo2tKP5mxJXrvrijCWpqCFQRSGHFhxuoWgvpAJb/9hLO8
QoRndZ+DUlUFQ8cSBgSug9PcHLkrIFQ9yt7dJi8ZkXCRBCLXm7YiAGj2mAdjF0SH
o2wYJRqi3WqEpDiggmZjWKdkbeosSchG8AV+eOyWjwADZ4LX/KkVyTJWV8pU76gE
fAz+sAGRndU+5dDNGzixjUEXhGEQiEmD51n9PxT+EbRiyE+OeWMQjONJiBpY6a/O
5T/exDEetchz6tACVm8uVV/eFjoyoijO3+ff5VNtz56PnS3W28flyoYQ9LZsK+fE
QE04eJoIzLMtqOjScmFVtDu865JBFAIYDW/121sZYg7E++HBn/ohmLF1n9JQyB3q
FPJVVam0ABCVgTJVKQPsv+Ti+NkuA//oEOl4Ch8Ijo8K8/XCV78Emej1uy9egled
HuKuZYB+X+3RtuJAe23dEuwd/41wkvwmEacgJps6sAdqutyWCaNz74AwzJ7Gqd6D
FtMxargkBoNymsNLR5IonTXLlFrao8J3ejMHRRTb2M7IfLKeu/iNvd9UY1EamBE5
DiHh8o/hQ++qP7vMSprb8W2MOTjxc8Yx08eXUMMQiCB2vpq3sms0HUkbTKcrf8Zq
TYKb2nrJjkU/eg4vr5ycqPIMbbV2jvMPpzFrj8w+bu7jDidzBARXQ2lVcpGnJTTX
HtJs9ozrkMOrhOFN6IvBTBtDOJconYPVR+4Ie/n0s8kSdkB9ttnAfSNFKBLKeKny
Jz/zVUpiqVnz/uJgPMkHIFecZfZgwOQmEzcNQp/Kp29onGglO0emBi78Bp4xQDzR
EI4jZpCZm2ni4qyTTJ86CHLsfkappMemfHDepwJr7Zf+ZYkup2V7c7kQNPkdmEiS
49F4iJhA4HLnB+pUM6jObbZhtjDqlXbrTO1Zb1TbZLYrUc63GRPENnONx+P8QAn6
X080nidFoHVXP812ZahATlHzM0lERzDvTqgaL7rRsVm547IcsBjSZoHYGwfM32+7
vGaBMJ/kZr/dzyYk9W3guRL3GKVc932fl+as/xOs4PmkQ5+zb8TUVayoWVdHBC5h
4/pD8pOueypUldJvPYVM4czfe8Y0xN8pm4XS/Tp1BvUgJsLLMBy2nEYaUb2FEFVq
7Yy6vcgBlD1CM3A+kDuxr75cexVsPBr9tAUjBfqW8Giv75p/aHKbpTNj4Rmc3ZLn
rsTcX9h8mA1+qwjifv15h893tNcvx+6ampNYd/dPdUybUnUUfn77V+CcN4zUapxl
c4hVou00l7vLj5gvyYjI91qtLQfSKkAd17Jq8hyrFFDAc98qU+GB3JyJ+ZILZZ7I
oG5GesH9LhTyTVjf550Jk8Zw+dQzboUIGtFUDMvvhWDF3MZSoH0xlpHDoyePejLh
gXPE2dUeGKhmE7UtuIFlVQRlfo1GV8pMumRkZA39Lqy5cv3IKqOUApy66v6NH0Yj
RsfyCJg8J0bpJT/1PLJUlJyLJa1kb3cB4IfZ8qYr0mJVXZ9ghBNJ2Y1i5p+ttJ/8
C2lwzorDY2lrcRPqrUE91zczMOqMa/Rjm7mSDJcIRRXW99BP1u6GsSDfZJDSkYbJ
oBEx79pVwW5/irZBsoXHX6xHjoFO/asHAfTxlb/NbimQn1qZJ9mXMHPdiXxD25y2
f4eHrzqwFgCp4zffhIiNqQ8FIlHPaQKfcsPcCHfjVN4L3Zes3ub7qAd1Lo/9nt+B
wxozveyZoF/tO2oXBSWcny42gmlrnWIBKfRg1nXw7idhoyezM71VO4BKoZ603s+S
GRPefsJE8ANO+yi2UZJ9DOo3FniIhDjUETegr46eWAeRayRwPxcWySb9GrNzQu+C
uoeiHa64gYv20J+uKPJA3CUX5hIM19t/2dvnCJqAz6Pi1RpZIg6poKIlsfrl1v14
MJWm+jjEj9VMuGuKNFThvQpoamTDq/IXkur3xNWHrIGlvx8xj/ZYsljBuIL0jtzW
rYPmLWhD6cwSN0qePr8wk4FCuCTcoIqe1X2wWo7MQt66lkXVcwcpGj+Bw2eJ+gEL
ebIyJr32V6Mv8KY+mcNQ7Mq1detFSe1bUsizF8fD/ejlbBOB0LTl2UcbO0qa9qIv
sQCRJihQq0+GcrF2RZGrK5I2qMRUzSuwpe32X3H4YvxkKbMwbgpmOCxIq+obRXM4
GvPWhHnU1htvBFEz34egWrZL82MN+c4tkyup3ctlJcxQdBkFYDmxfCSP2/GAHM0h
TOxULpkfzlyzCa9vIqo0DGsMRnhGaZjsO5Jcv1UIL3q2o80WHKw0x2oq8dmZu/Fp
yGEIJvUmHDGZ1VpQPc7EsM2JIxB95YUQsTxCsrOojt6JpSN9vECjYS+ggbsXsyT0
Kj72iN/rSduGylh/ApV/9/U3Z1UokeHr7h5gxXHYhr9H4sQ09XKwe49WP7nwuB13
9xfF4pFx7TcEr51i7T4I8DKyQuCFAdkiHX6EPCkBWQHFZMqR4f7M3qF74smktEOY
pTgMWeZ+YD3QqkYkbIDCUvtxxGocymFrvJEBQZ11COKZQpVwLD07AbDQ8H6L2fK4
T+24q4Swo9X8s8tXejNdS1ulU60TKsKmdmAnA1GAMQ0I0EOtfHNpnN2nytGAVcq8
3t8wfoq+kKbZYC3cRowuXQ+15+taRt19uBKAzv9rDhkAeIaqK3sE6l4T1fLHp2gE
uhueMwxzqE1tup9PKHWbrRV87PHf03GmYjDSfpZcWH4ZtXyFi5Po9M6iwPS6KhNG
30nXBT0pTo/rgIfvjZ9kDDprv4hyvWKK8l6/2jdYbFmsWkl4OSv5biqvqvyJugxw
jcod/Z/i5tnCa/n+fNMiULncG9LWdbfP3s9AwXSbJPrXl4bqNcEsPKgFFn2s/bHs
0lhmG12VYDxqCqDDZvzjhXVkxdPrpp9laeJ1lKYSwZzKoDnLlVg7BFJGE2a5bYGa
7xGxTwu9ZPIMGvMaXYX43H5FKVzuI88zWHZRUqtt3YH1312zGZQFL5yDPrjSy3Mu
/w66R3nO4EfjvG/4wVwc6dgesLHlA58j3jtwo6CCPmu/PbTGbioRQiODDqh+RJ8q
AHSN2EsAYRrsy+B3NVPhzy1Fql4+ZFtdNIOIOBeWF1BDM8AFr6yaLutDO04ZFR1a
4WjOuBshkF6nN7s38yjDA7ZizA3CWZn7aHnGbKsm4DyNa3ddy94NBFUOjKhJ/7ti
WRrJRbJhWnKKl2iLZQ7UE97HQq4nxi7wTo8cpbpeBx/10Gzr1xwrWtOUD47gBSOp
tmYFzttmDYaAxUkgZsg+xUkcCKEIqfOPoQALfEf5qlRuHKsteNYxbDXblQVPwXMi
Us4QNyomiJ+69FZ496gc3u9mjz/Rt20qpeCdLKNMWtzfFtz/W1SKKHRgeaLV6Cw1
rvJkx4AywD458YHHotbl9mhtUV+X9nF8a8gfel1CEJKw0WKEEKnyxztOessG4Vak
X1ZEDh1ahXKeEOU1RTN2jzTs5KSeRtqeFychr/yr5F7JKMrBJpRrEjdK/Ubqb1vD
Wy9jAy4KQDgapIm+0LF18EDs34p6YlYYUcej16A+lDr6j7hPe74Sk7wbV7I7212X
QZyUDgkW+HJmmGk+pIJNsuXmag6cxDG0dSeCtktL7TkQvRkbjdVesAVc0/rlWMpe
i6X8YpuHtdyJd0KuzlXtrKC+a9GUmFcMri4g3rBLeveDlfs856B+PLFKcl25WcVG
KcjLUFCU2PkpunuisuTgklmqx2RGHhQpS8HOHw/AZ6b1oYAW3PPDdHndTymPnhfY
bCD8R7aDZavnr4kitNuZANWS5TK/k28Tgu5lraPogA30KqBZ+g0D+nVt3yWJP3Ph
JEYbFr2OudGXbWaXpojw5oHxHqidJBq0xH7OGm2UuJuI0oeu8gJ/7MRxokZxMlMT
fFItGICVxF9cE996cJZCpGBycb6gcZpfEfrcGUJQ+F1xCRNUUlMVpW6T1hfFr1hB
Z6POw92EE2D0a5Kl1AZ7RVMpopfrEyurHR9BapTW2rkk/yGP8g1Ri2guibCX84HY
36NktyBvzKJ5Hg4zm2sKyxMjQNf0mlIEvl4AyM8FEpjU3t/iIhsrDmjQ/S0gybvK
sZ+WbVA0VxSk3Xc4O/zcU2Tw9IsYf4Cl4OtS/stuQZgQHkEphD8WriJDOOAw6kw7
NQDMgD7M/iUnTD4c37W7GGVekmkW/06JbGoIub2J8iYM4IdTyPS7HTlVULzra6VY
0+LjE/T1cFTr81VQiDPNOdMhM53Q/mQKSaj2N9YZ+2dNeA60u73PYlCPPFr8LCly
ONnbzD0MPDL/y7qbZTFhN52p8kQ6Ivd3F8f1n2HL/VbSuDx/x/Mqsz05OhZnH+/i
/be+FrQTwwKN7qMgOXa2iajDJQr264Wwx+NamihIpXJwpZIEqIMo0Tx1CCEfmcfx
tarzZJRmxkHYbOJQWGPg8KMW6lfoMR9e8vzHfJLqLNx6lzAsq66lhYYusm9WRPyM
q/k6CpXpovoTSMpH7s3xzP+xQK4x/yKdqnRzL7iPnP/TmnBnQTzqOoLMa8RYr+q2
01es25cKgIXw7lWPxEYYJ9uItpgST3MJW3oHNX0eEczVgZNN6rYtZkKADhxHkfYF
HWCpcmy6krBdJ9KvwM90XHx9A0BkZibf7bnGRU9ZfmmhEodef31cGtpBxQH27cHW
RwaqTmI/xUzoA1WwggxvpTvAcZMjA/OKsxIqD2/zQUoYgKclB4P9aJjhzgPtWIwx
fxfcDfbvSj7cdQBP/mMpH3MljPxPITKX0oi0/Ou0niSohMSylErvmNcqcbWJ9RDM
maq2BC19E0ycJlG4dit54YPeOjlvhEXlC1XjQediFCPVRKxSzXJqgC7dWmMwgpX7
ADhktRu7dN1n1hGKIT/E/Kzjx7at72IakKgf+G57e5WALaV76wxjdUnRLSqfm4OQ
zDRGvP8hh4BibJaNOmefX+TosKRcEmrKVXfNlbZM078MobsrlLReN/7JnoTjbu9M
VUN4g8RjhATmKq84IfQXMm+fWGs8H9sg2xGrsVKglggXeGBN6AyWsOEdb5t4gzZp
1BR/Q68uOk8SDMu/ksLJHQiw9kPCuDPtDOObpmTjq8sPKWeqt5vyXLpRKtmKKn3s
2fVltIYlvHL+8yzrouHaUn1NomLzEjUeYyuiStmE1GdnpyntOUXrG3I6iX+Bg04a
wnbJpToBIz3FgysvjZC8tJvLSDe2aFE0KyHFJsDTH6RdoqVx8UD4ooxUT6+5aD0g
7K9wSuB8dJD9YJtjT8BEcD6rmKAnwnGOCORRzSGF0ke717EgrbkD1pwjO61ZIrl6
XWXw3X3lY1O13y+EgguGqPItL2sVNTm/rSkeSCPO/waXnFUUVjz4Iv62S4CLmAzT
VPKKIU6U2A7iTAGgS6AounK3vPGZ99QKhR1pPfI91LoWTqZogRBBlY5+92KZGGAc
ziRGzD9WSNGZOsBGLN/lv9pCE//9usuyh4TN5Tf8f9Tn9YCsOS3JHB/o9uNLszFu
/dv/LAraBMu7/qS4B44oRpm+Rzy6iSZAEdB2tHqqG4xXfjLSXxVsLRGixZm6otzK
0EI48Y+IcUW4S/0zb50BoqCMQpbl4Gz8UyE3blLWIbjp5ECPs8kjRnHUAoSD67TI
17LvbaLxRpg2aM5ocr4agfea/wd9690SvCNqVJd3ndeiLrZojtyMVEgeBcis24yJ
gE8HNX7XXIBMpeafo1/ZcrnwZFMc0q4dgWXCx2DR0KDskrZqmABOxGALBHowRXJz
KZ/UujQKgnQjKiHZVtx/LsS4xIIENE3AsFTefOXff8yOEE1LiS5Rlb4K3FzBjdzx
YePG9WQAwQS2Cb38mT5BdaZj1Hcwoh/Gz5JFWgRHdS9wa0DhvELP+eN0Yxb9nECm
hr0UhHOrvzqa+ySBWGg6ohtWZQxZEevcRpr4PAVFLeR8jCQEEzf9fXatWGNKVUPs
szUPCEfevgeZ6/gX16mTWv8JkAP0lJm6Uu0VNgpo2CtNARoYIXS2Vv+Wlds8Yz9A
NotUXz8cYWOPiM383YOBbt3OT8OJ6Mfmb5sTcD6sEn40CyagdST5ALnbdyb508MY
lM1S/FTDcbpa3/vnXYkywJn8YTc4fiqQo01boI976pPxrFvK8T1n6cpHnAaUPxKL
uwMtur8O19bJepUSSW1m8oR3u2F7ga0kmXnfOjHU+GlxAzGdjmllOQw2yIYXlm5y
AUjJsYNHOjsbq/bJ30HvL5zovzVkap8GDHcNajM3pfBkY4gwxk0plQWwfm8jupTL
/kd5phCpdeetlR+vwSiDQ9HHN7cFCaNFPBYzs40zSm29kE2K4L+H73UcS9K2//K1
0oWvNhz1IBuNY/0Mm2mzs+VSTH22bS0D5XQ/HUQSqvode2Uj7YO9X3060u4pQcUF
fs3+7xKjVvdyWAbHqWg3VmnYAWmqsKdYoxcEOKXaDxKMldGAbpAMPOFkcdAbJc0B
GcaC4QM0y7Z1LPzhSpl8bD4EH+nW6D/cJbXl+adCAjirAXrmxrfyx9/HOaK4D5kK
FCstNSHJSuTWsAB5EgVNgHHL3sYujim54r5FAGsXafwhwtrXEPhCxMUVoCm8cJw9
KIV8To5NctfNyMkhXYs4W9E5XvJUG4137PbinB3pg1vWPwd1m7cr7WJVaUjh3Hwj
GxRMM+SqLTPNz8veSrtLmu3xj73qc3Yn8ThcPR3XCm+t66T3hzH2poXjEjwJxQSz
uO5dMANu2i5BIsH0fsseatHbcOn4XvacOpx8kX6I7Z28zRQ6aEvAG6QG3srqJzQp
dlZc0ACRXmxiUgkOVZm0dmyuIDATT5qowHh81mdlO2/Kmtqf1/FsVI3ZyRM/l/S2
wEaNOPl/ji7/iJ7skmP64jm6tktZv4EBF0Zo1LGcUDNU/vZhGwvZXi3W0WzhXanb
Ng0aofIIVhx4sU+dmOyvur0JaP75QaU1d5whTi1zmpPnnDz6hGSD5/8y05DW4HYh
4/917tdPUOoXpezLvfnuwRSH0YJtxCccB/3AfcHLfr9tNXSAn+LGKCJp8a4HaaYb
KkXSHS1CSBYla0NI/CJ1IFRtjxz8V89N0SWCPnJbaBLRt88DHoImttyaNWjEf2Kj
IColTpPu76Fo9nguw6X9yeagYdfFOkt3jPQS33OI0EPPamKZK1ahLgDbdVXTpQiL
kuqYUwuT9QTTDJ63PFU6sk9jA5Q42uLqd7k2IDCqy4Hwz4amxIl3GfU4WArn6uYe
S3wl3a2Eg2t0nJlWmfwcKnmgA0Y/rHaA4sNW+Fa6bLy/dkmXGBmspVohKub9jMZ3
ekFpnI1UtVUGQT0xRQBu1nsHJvdDpZy1rzkzj3x0TfW4zjNAeH5DAcfgze2+GkAa
YbKrlb4AYOuDg7WNfVsIJ0Q4lgabA0D7vp8nw7Lzs4QNg/61Bcpi2Gs3XUEMqbW8
xKFnWs9bNvbp0vG21ODLWmURJ5Adtu0kNwKcmx5xXoUcdvHcPgyDRhNrzWDgWlmE
K+6XqMKhOYNIPtI3/VSQMb/U3Aip650JvBf55HiFkZDRjB17tGZLd5pvowlgdF/G
ufnH+pW5cNKDcCyOtvBtrcX2EuazXZ+SpJD2/bw1fRmBZiAHKDlPLj2ydSKFwDeT
wfYqIJV6sTQSCkNueFZeD9dJId+qMzETePw0p4FOSdGpC8yeXIAESmGelE2+q8Bq
89WyBqZtHTZJZdCJpYUHFReUbVrMAhDsdhmYA6S64KPu01TX2Y6rA5Ki9g1BjviO
yf3oSkLdaDmaTbgARu+f2seuK1TuY9CXqzmFopRO1XJRGlg6Ma/j3jOMPoR1xKox
ilJKdQDdf0oskmwCLtSkGmjXa3n7qYPQlU+X/k6Pz+yVssqfyvUc5StST6VUL8Ui
XJMtu1TsDg1/l0KEd4TUiM4k9ZxUnrJBdaDxakU8sl/8V4bokkyoP14ItghqU2ul
61XOKK+t4v5P+JRdTRWL7MazS4+g6tkT6JcqjvYwAlfpfiR3bOnBKEZZu6QkNCfA
o8+rNEqGt5wOMVNVIBMAqhq53aaUMF5p2zT4ajAxRu937rlMoLskMyXWUAZMKyyJ
vBRo4X1TUV8hJQB+ZuX1QsZDwlEmJ1nw2OBX48z8l01IR2byLepSHE01llStr1mn
NATCRp2bPqAbUGZ/bBXw6WUHnbPGR30yMYvl0nroXr3oW569NX9n4C8yFzRRu8aS
qFq5X4YRbt1KWqK2D81WjJDwP+Z0PgQwoIdzi/VIlDOt3PTtBcl0n5FHky0xYJ6X
Dr2U/wPjeigrpBRa+8ZLl0brhmtU/0yCTJa4nDlTgJEFe/QxN4SxXFcY2hLZ9qd7
FifTY/gJV8ZEd5WUVxfLy+S7gnfAbYzh29W4zu1QAHyF6Jvo/KbrVByFVl36xfzJ
GFYYqxX7mn/jWx3i6LDySzvAPk2d0nEoL6ILHce29pOS+XU/dzeYmDNAgWKvrrU+
i5T5Qkg61XluprG9GwbhvukCdg0juzTWxWTV3lC9qXH4Ezwt6HXspXngQLC0QD9t
K7eSY+w1X9JF4sPPmzOVpq8OzZj77Ahik5EllhzharYrjF2sYBJ+46fqATzZDIov
mb64kaXKyNPsazG7RrOdbkOIl3qNWU8Mpejda8NIyYGOCEujX9v8U/TyUsKdbKyA
OebADcjdyifOEUrZGFXiixnQ7t+0XpTzIg0ZM3NfZ0734I0HX6qLar2vawDmUenZ
syBipaK6Gupxv+IwA8qx7ywzrKRbbxlATUvwfQxxo5xx7xdW2F+Yaqrvmfycv/pG
/4QpiGnUlvdbrFOP08wXRyVEk9EcJBFKRqq0nLvFtkR36uNvm93yh/RASCRxZLxW
5gXFjIz+MxMhAtphXcoH0oDGjfqTfXF6Lcb61LpMKa/PusmJqBL7uQTWKQn3pYEx
Rsx8kGtWJ7k9zvs5CNkZopIqN386uY+xfNZUtr5Hc9HZWDraGweDqo1Lc+uPaV4A
x0zaTNrscnbiAMWbZsTD6oV0HzY8Sw3dFxFzikzHxt+8PaibRYVLx+iG/u6yIGAn
N38W/ZscZDsojM5wkeg0W+vrBtPAgyNAGT5uOREzaHWS2nAe0r7QDlNK3LOiIz3l
PkudhJ+E2z8qhXz9scDgvehKC0BM5t8fxJaANmS5FBw7EKk83FjZUhP/ba7HnhDv
9qxzXm1jg21jQA5BhUQr8wc9HCFb2lnMnH2uhK86UMO4u6ng48K1StFM+qfe2G6t
teOgSCiOaVVYLwx8ZkWPYSGS+htYJmTrGK8I2LXWpDiPxqf+rL2nxW2CRwrKuO8g
LjJeOPYoyJ+luuzVVmidQC2HwDzOumJTwfdUiNzg19QORJSYf96yB9y1iGxfcSTF
87y95pDAop03DmSCgbg7oe2W/YmRHUe0+2kaveAXWdjL87OljCPBqkxLIA5REyAx
cqs3ewAy++yjuNgDabbGm65os567CDjLa4gKni4HbbuFx67JbRvM/rYttsMuoRM1
RMms3MxKqVMTSJfydnWTsMI/ha13WVpZqAIxdO1Siy1SZ/v+c2xncn+JdxZa4Hyl
aExghH04bflKfGqe5AVqZD9ysftIRjBDRm8dwrW0Hv27LwMnwO5F4NUYOmX2nMVI
7S99lYnXcVuhkwbP4y0h12dwVkAuvTZjOoIXr0pI+gZ7UMPBP4ivtISzIZ5Pnipi
mRk0B6+dNQ6VnIOzUsYwzKm59/+v7ggGijbONWpgJct2vivIJnnbdWNHeaVd7R7F
58elIDIrklzJ97HtBY/rhhw4/06yi5iI+zsda4fZo7GnNUqTA7ElWi3RH6/KcuFh
QjyuWK5SLvvtZUktcMEOc2LYKGSjEO/SvvNB4cNxgJ63IRp+jGxXk49fwV78FDoi
maIa6sICrZfNfOkWgrFSrEaFCfG1lpQHQshxbg2MklHP90Dy/ORLJKu2vTEOoGow
PY1u4qk5t7u38bo776DGoNzaIeFEjxM107lfvEqKY94ADcYaa0KylTVPh1+h2QE1
kRcKKggpzfi6kuotcNUp74Y8LUcojTVHPUQ6pWXaIbNUMpuVpli/O8yS03j8Z3NW
NpIFomPtRhlJ7sSDM0cuRDMH3ePY+vhRDAlz8TcqegJdHEgR4TiCPBWXntQkCDqB
3awbLPDENNvBHodIiaO7kg1bh3AAD47jksdcYa+YhPjFqWgQGs5+wYNkI34URZFO
IEKKORVNttNE21bo+Tf2D5bl4G5haUDIlcFtDg2ImdxbohUmG35Kj5TQFRxAaklA
oKBwKaTQG4MUMmod7MkBIgPiV7SpKsOkS1sNWhjFGrfJZk/7je+f/UPH2SU2WvRh
5bv+/2Kc/sdBt/3zSpKu8O6jgJlaDeyC6/KtDPB5DXEzIpaTCPZiI5L6XvnAO4hH
aJcm+d8dsbxckTN+su0H6SUrw8nT57eAYMS6gQdHnM1KCUoSFo6n4j53aun+Q4Q8
eI3Kanjt6N1Dg+IVrdG/RGOYbHj3qy3Vfc3HUhzuEUqx9cbrzR2XW5PJyaJtBuyF
Y6lOeRvvlIMaR7fbDObHFgGIZLkkrKl/xOEacFrSCLS4uF31Vmg0yYh/YXKNcOiV
/6x9OnreCxRe/W4E0ddPMECqsYnrDGDPwipgoy2cYH6f3EuHz5AFkqI3hqiqfipC
GjDhhqoFpFwtOT4izAhnURshKhikc6BpeQbZl/i8i0A2ApQp29WxvEvuuMBLJO8r
/3MJoU0JPUmvHAnExW/Ks7ywXfq9FkiN9F7TwUFEewhwNpXyDpyEm3n6CnskjSag
VuqrKmcrOkOsMPTeCCpw2jMRwvLrNdOGMCOhs4164lImfhS6NUXoJnxy9g29C+ND
GzOxJiwZICO0BBnOy0QtIs8KPhlbOejmvrNdD5TGbs8ndmTEc4dZ89FBFEEtHdYH
ElOnPPVapOb61qbulbShd/by1a0dZ84HlQn5BK4KWWCPNlArss22xD/bzOr9Bel4
HXL2hrzNrATypGh4yEpoGLLDRhT5A9EMAnZvlvqx0T8Kx5b51sY9yvVV7qO16Bus
lOOgTvHnJJuC8lTrkJetUe122HV6ZIxZdfMExAromzv9F6wfdPjo6P11TNJ9y78H
AVrermc3L6aUZvEYLTutzzT1Nj8E2V6KVLlbbHI7e3aAnsCbps3lAilX5jTVgvoo
uqd/QeVx1fts1YuO4QXayikO6jqnh6LWRSaijIpbhnzBy8SCkYM6svCZ0RoJ55vJ
L5JjbsF6bEgWfema0Ky1o6P2OjiKWIiuAM7Q92LJ7VTcHVeCFiYaRtt3/ZaJCgxW
Vm7zPs+5zLxBV+JFtIzMYmFb83Lu3ERcPRKk1t2gmui7MDBJDbKzb80zL4YBglSs
pXS52G8tUkXVbNJjEn3ctsOGrRNQEwrOGfwXk5uCFXuzz2LPZdosdMKhKeV8Do9R
9p4meOIDxQftyLBganA3v06L/s0BjdtGSDpG1/Cp7Q4KXA1v+dtzT+W6QwInXa48
uzT7fYJoTBAamWc/JhiTcXIQUes2V45Hk8JWGywAKnCJxcKGBx+WrZB33L+zi7Lr
qB4R/8FrcsHIxZiJCpkSfpThZb1epJPaKW5mDWzrWSmMfpP3oMrU3jXSjENb77/Y
yNU2CEYXgMKrZexdk8Doqyup/NuvlQMXfigHb2cGDzf3+ECqszEcY/M9/bHLvuZg
rQgwlN7eymVeiy7goiRd1hS4OKuA95lisudAudcBzH935cpBdQAquSY/sY6JQv4Q
7vJXV9aqXv9CZiaVkKOO7fICwr6NaBtLV2paB7dmnvpSM+cUZoAOUrEnNutUZjqk
8pC0DXMlAD4ktajTcWexBXQt9HSmZjXo9XKCZki/Td8VePcDTUqtVFiiNlKVexeB
Cj3vl1/t/LtagjNvNCfjWRFY6GP8j/wBVDSPcdknBefUfHoCKagt0XLCFm9KkW08
P5mXk/dsuEXyHWgfkl8VafzH44f1N+Z+QrPnP2W5A4mCmUmnDhraRPEODI0DEVvw
lZig7jLt0zPqPUAQCxJQGygmTQ5Ii/MaxHLzAmbLIN05CuNQbhfbxVdWcw1cjzOn
K5qefeMrk5m+idr01nyKZrhjSE4yFk+4yjPBXkOYP8C+i9oLl0kG0P9Fw+eb3C67
HtxxrtGwj8JiUwuRfXV5n3lC3m890gmGNJLe8m8l1dATxDTucfXjtFqnLz+sdH5c
vEgJQ0HKxTh47wYD5NSYpanu7UCCQaKYZFj++bH7DI7wWHFKd5lLhMNEHhebS5A4
X7T+a+znI8SRxE8qHUZ2Lnl0wAzl1+6DBxQ/gyn+1Xd1xNLt0yXIbp/VRCHvxBdf
KzW+Qw0Km6ied0rxxSrsWx+fCbtjwTUtiMexhwKiraLh0LDm57FgTetg9noRttjg
JAT0npgMmGQlJfkhAUN2RX5a/CiJXlkvAqj9uAxNn7tHci4jRfVvSbFhxrsMyTb3
JXpcKx/4KUENjmHpMqjRsqbusqbjehsTmjpQXMbsK9rYzJp7i1STomAVH+U5rtww
v2rRwyd58ObKUqe4gzNsZMl3NX2dMjcxdE2BsS+2dbMCNUeZXijYNDpnOVpibdTN
Ocm2iFjB4546LtRrf52xnldoCVFEAitglqN5OG9EIJL8EBwcCly/o7N2Gnp0Q4FK
eCCfnDkTu6SjTUQNdHuOtwCUt+Z9ZRDmK98itPd4g86+DWxGwnbdDtlO80JObDzI
gPLol4R4YY1kd6jSaAvqAW+XR20x4Dhurxf0MRWJljlb8kUQW3mfzhZHNxJfFbiu
Xl45Fa9euA2EZJ275MluiAkJNN8A6MAO9S5+BXMmU7eDxRgcANW/VKkfzzQsKWVH
x4/USR3bJi1ZxUkCM7Uii5YxshuhhkXYUoXMDcn3SytdIW7zPBQUnacgX66WLV22
8xnhEQw1rzSzSYPlpRxwkJXSpay8oeEquO5fcdOWVs59KQjvsBMSGekigEChxfT5
fIm5xtcNJKDnT26Yj/FzFM0aU2A+DLs87zhZ8NAHZ5ZMl6YxR3Ki6NNUVESY8Ap7
Kvvfyv2CF2EWNRyFFEfEK0aqovZxoOstAAgt+ey4cBaKknB3fYVkwvp/f9irIWOm
ZUQ2ZHfHX3tedGulNSDqFEHFS7z67CBU53tSlGu+7BXKTN0pFRl2H71rD7aOH0Cd
Zao/9K93rSJMlPMyixrqUc7W6oDoQa87UGvrAuhKRL664AGZKY65mfZb1lmCni4L
mZx6T8swOUQZFvj+WBKX9KSa3nLtFmxjJiWaUFdGyoCxJTiCXsiz9bAKCcvgns1E
8kIZzPZqTn/OzCOQccsZQn4w/VaYC/FPnAW+OZeeB9EB25D+HlZOHj3p1gKll1Gg
bYv4V+tvqSmTY0FR+L3ZRG4Sv4WNfU0InCai0XlaczPHaPTIB3uCDDLJlJd2FKIB
+YmbLfjwZsWsQn1KPPGY9Izndsb2jGk05VZ8GvrHt5zRaNxdv4bC64rajDA8xYeV
zBsgdra5Y6U8jDhdy/yrndNug3ho4NffJurX4iVVCG5L2wqgeo5wAHW3X7Y+GoAj
oBqD58oRyONWujiQ42OYEwE01ZEnNsw4XM0O70tEeWKdoJHEp0JBemH7/K0b1AD5
wg3OIHZgrh7v2RO7uIYNtkiPb5hcaAgzcj5vQ9cW6NF75IGapSkH3tvyIeabdgiN
pciKdPhchOPrxKlKkPKjjiZwV/wQY2TqxiyrHViV4z+ngLOXQ0ergZIihOGt44km
7gZzHrcJM5vcocKaoCVyu4+g8vFdHgHENNliEvLfYkhhSK4yg9agjpPuIBAGXlFl
WSDz/1F30sUuWc8oaFU6jsNMgDhcBQVXopXroiM9JygdA8J4VcQ1MGMuTi35OAZo
pS2UiKgWUFWtepRX2gSZ7xCug8JJSNdxFrJ0cVwVAldBr1YCc7A5YiSuvSLQBoI0
C5emm8mlSxvk8OopF0BOoz4gl/AVbaROGQhT3Dvy5s0Xf4z82KZ2abNy4Z9ccaGn
S20FdgHbKTCi/gS0jCRFw7tMenUCFG1qyul1EcS1INuUFfoUJvjkZl32KdO7rpD7
rsgjt+jflrTPg1JhX3VwevxgtSuqOsUbi9mBjYHC+0sk0LzdjqRkJ5FSSuNMBTlP
kyQyYvRy8SbYgC7jEVqJ0Ab8rVev9fnvbJ5nzLF+7ygaYshPdvz9quOsNfc4WeQ/
A3j7z8rN0GyZNwP9MbVDZwftGlturDUiaf900CiSew/dKKWJZgeLy4tAsjfTJnu7
mnoBuK03/GRvmwR0U/QIEUoShOA4tR2c186MHbi9RoMgXb0llIlQzi/KzgDrqnk4
vdxf0Y1kH7d+BKtLUxfNwSGq4kjbZd5Ll21zBJm3BWJuNUBy/Vo6PGD0e9gdFYNU
5oI2KxS2MIvcgwuMWwZooQ91NdfOhYBuiLvj9RO/t4EtlM7B11deZJ14JVpeKYRA
H8F5xURAXN6WsWxMiqpV4VHRPwpYJ6vI7SKE5GGNo6wvSJd/4VSCNDZWxLQu3Fj0
Q6s/lxpj/36fH5VTTKsg9PqpcyMFoXvuyMViQatJ027c9sLjQSRlDkCeXOCWjbzM
KudeB9qGEvuH7iY02OiimB33+5Ts2oRbezBQh8Qw3U8sd9cqu3TmAFJwiw5Ye191
nMP+0AAosHGoAs+oHp+E7mTnWZHexMVT3sWWCr1zZC0M9MtNww2upQ8WaalAWv0u
A0VPVFHqYdggdBf3irbx35HrDkrxVU+bdb1jAp0h91BAI/+3EU1aXUT5GB7pJeBl
CR6/ealFEvbSPYyBga4RdsvHn9IMgU9s1u8Z98vsftFxi2d97JqY1eHmgcERL/7v
E91+nhSFWQ3qvI0VHRbfUSVKm/SvCOq9hfXnholKWcv9YY1u8FOXtyZKtgHfIQ8y
XpjJolYcIe1U4rwTDyQD9NrMuhtmfB4jM8fv/7PoiKrnZlOkr7IKkx3YBntVhhbR
t/LWk5aajpioEOtq4R4Cghcu0vYFEDXWAEU4zxuHYD0EEKjWQ45uBTTmLFG4Og0V
w7c9D+RA2E/UtZ8ziKTlH7hkLinASPNHU4UqulyUCTGc22EkRN8qODyu1svEoaGg
eUVPMWkTEfGELnaiZNkN8qfq8Z+zpXWSOdjZoqV7HFUZYSxPuh0y5yCztlPrFbFY
vMEaTawSEEGqkafgMgEfzfjiU+jTyGkrJs2p1r5RDoW0UzsX/hvjTQYNaBIeiM01
kr0OWocN02EOBbUgmURgKEAGHoHEfEWh3v9+0z1jLgll2dut/GfoT0cWEHf4+DK9
jAgfj+mOjtfecDlCGCZsEeb5r+aiqI8cd9+ieMAOL4HZYGiU0oDeadW2yjPyGcNr
YvHdC+treJ1NkVDzCxN3WkdMYLDH/MhOTiBb33mBZ3rQ4KCMILCzlzaWe5n7+p6w
EDb0fF0RxWFY86g2axhhE7gdHAZ7FO489CIHKm+19cXYNggL0mKZ+ooK2ZJWfj1P
3/eFhrzDEJ6jQBETz5gm6jXTsawFTwwyoOmSKjtxSAV/Uyv3yLtllGFV/BGnRTqn
jjKfU8p8Y8ZQv0bIOkgdWRvvDb7rRL3SYpPP8wNzx7D8JFqaDGqznmqy2tE5t42r
WY3TBX0tnvKQdUZ9R/DUO0+J8xAF1SaxDBj5qssmFli2f8Q9yl8fGqjbarhO4xCR
txIFa0c9IhgPYktM0QyeckFqTnGKkmpRSP8HE3ironrGl+gun2xd8LUnu5Xf4L0t
ee3dWICF3VeVYnxg1qShjMiJAPrueyZ0tC9EShyX5lZetb9g6gvULG4Nq18x+GwU
0/+yi1TCxiMq4NWH/Ljt06acTjZug2e0i9zhFM4glVYc1vZuS/IEBjwZv5I/0wYV
0Cf20ag7vqx/USBzSW62Zbx/ZCHZwFHwn/vOI620DEvURsRgqpllqOJtiXzqKf8C
AtZeLwPhby+ZUT/zxwfs/g4CrcLvmrgHrl/bNBpvLPHCKw+oIsE1geESj1PuDy7B
XbrIOTAE5qoGHQgbv2aSGfPicKLZ5a798j/NIDrRfqvmYXwCgmdEWD8hdNhEko1/
nvA5qj0dHHrsGFFVGqkJp4J2XmdlfygR8PywIJos0rrTfZRtbFrKMmsP3twkSMui
daEQIpTl1xyrcQJshdT8rLuAKsgF2UqL7D+qyB10z/DKo8euMUUk23TpPATjLei5
GQMR66HZewdi/DlfnVVlX41fE4LZQt0zIWsOJkNCIpCqsVgnsSaqJklj1HChdwmO
zUYPvMdHHcklqrbMeCjz9FZi/Cos7pW0ntES3EBc/dSw11cFieohKSZhcGrt67a9
0Vmf/d7eNqRjNb4vJEZjAyd/85b2Vvfwuos9EBERtbdlO3p+0n6zgKc7TewrXDNU
j/fgg5vI6uAHspBj6gXuYDVfrgCu9Ri1t9YqzLe2tNprTaMY4xyAk7SP/4jloOlk
hB4uRjqX3wXGXT2GwjCeiajSy2wkbmhRZ5ZGLGxz1JnKy6Pxu40pG5j5CzSjI+CQ
NBnX7AZF3PVabDC/AOhsQ3vh+Tkx2QcikP0ybza9AkohkmrBczBsoox6wUldXiQ9
MwwSyDNKgBtPOEO95HzGMKkC27sLhn+zdksfPNPVSXlfRDGLWkHoZsLE8aBDcC7e
Fahohs0dqAieCCGM75p3V+W1cKRbGvxvpCApWoJp11O96DaHhkVeCwhDdq/lGY/m
BvT4q4UimTvUfLFKDnWDjPm4KkYPRsPwXE0FN/siFthJXxny1ReqGPRUjCOadC4F
H8mZilnHcjTutF2tHG7yhQfCM5ThJ0/QjOK4436SsjjkMwmYhIU/Y67wmDieLo0T
nmDGVTxRIcinddlOVLGHSKnj5qAlQuCclqRI/NE8Q37ixKBk6Lbi5QOGrE1p1G3E
mCziiFvv9+GooZDEaKyvi7vEtqhabSCUG1JRspxCROMZni5PVC/Xi3UBCwAdhr7I
v+uavNxdf3UutW4rTuLAz6MDUP/RmmPGYG4eEaPm/O0zgnBDJfQFgIYaWlMH+5Sy
1ce2PNs3TDt22MO7WwllmK9FBOfXdIX6BsnbX/XXVWmg5BZk3VcS1B9NfbdPwJAq
sJRyUvAGKp4x+VbNkDZOyZzny6GwCLzd7rFTiYsFORKnuDgbwYqtf9U6G68olj0s
Pvd4QLYd5E2HIwgDh1zXN8cJ5mImtIgaIWOdtH7LnSgC+NOIxEJdU9sxJ9XCJpPx
cX8ZWwcypRV9ich2RKiqXDXOKAB6exPMdq6z9WJS/ZhWxkBSQiLumR1IJ95YqpFa
HdqKRcbJ+SZFB6RwbyyMTI/Yoyp21EsiHdsxHY4RqV3QSJHiBXM+YpkkSjmxYhBb
2xU4zPUy6WbMx/i0knz4K6lLwk+3234oIAWH/ETiGNT0KEqA/tWRT+qx7IWnif28
/7YpwZIPWpNEAWVvcriYDjxLpEmMBiLdchqVG0v29z9ctQUyXiGr9RbALeAb354t
tTXP8iXwD9K0OqoBOrJhNBbnK2tdNPZjdzshxXKNBvED2cpSTm8q5VA4ObMlWszv
lYyjoyl+oNcEvnupszPQ5G8J0N2T0jGm8sH3bGlwjXKNcn1fMguXsAm2ZUo03N7p
JrRQqmijcP57uHlg/Mr3E+bfizQTDNNRdyeuBEYB+f1xfMfJ01sNwFX5Q+2q4GHf
388on1rUJBecyB5Yvfxw8/uKfOz1cLcICQUfMSKYf6xvyEfBx0gHPDjW2AnWcfXD
QlvjvBVG0o6PMI3SCicB28Hfbs9aTxBkjo7lO0vMZmzNLVukZh3RY49mVgt3CFZY
RuhvQrALbayZCJ/mzOyJD9mWTZPytqdOvu08fbNw6Q+h8UqXRDEj93fnesk3fO+1
jnUoZGTlnYTT/TD286TzrynhZsbxMGgsvsRAqmq8YWzPa68ux6wxKUoc217VrZtz
rsPr/1D7PWrCkHQafQIRSBjWFMCGuWlqr23FjoI9TOv8MCX/G/Ek+mcb6lXKcQpu
k6geGhdnoj5gccggfKxb3PzSisO+m6D5SfQ7AkTbV9H2iLwPJLEepj7ct1HBAu2a
xoyNbcI9hgQw6zWOmwfDKvppk0qMSU45MUbmePKq8UloWMYy+O5DydiQhIsfW8T3
YYqCJrKNyVXXt5+zCg+qt6/6WIAjmedcuRxLQwvy1B8z1FDVY4PKk1NFsadiaSY1
o0eFcQna/S0lOQILvSPWrw2I+m5efYCDX5GLgBv3cqWSkug4SvLLpc59mHHDFk+C
GlILyeYc5/QeaEXCLYQED69I0eokRtFP/iFHk5cuHDLA1UUxd5cskLjKfzUAJaAW
449BJUzB+WnVBB0TmnpW6YyiwTxZmZVvB9krMBXp4n0IxnmcGPBWjQiAtl3pJKnE
bdlKtX238Aw3NCl1TbNh7dCPJCree9loLA5x5YPG0GDBV8yJTM0vpQ+YNxLJfT+p
XgDK+kIGEj9YYQP3EatTWr1x43OMiZMXRanWFpQZ54hs/nizzsKaH7SF/w7Jdc4F
Eh+3U9hRMyPzqBVGnuul1vqrFthvAcPr+FsOFG+P+jFI5szpLrUUkNntTF6EnOVN
wW8gvY8z/u293iys1AuplVnl24KSbd3EkzHSCkEvjWKoWPozzM06o2D/+1u5MIeW
mq2+om4o5/tBruPCUeRGn/EpJ5VgVJlmjWv7NILKiuIfx3yLgzyipvFgV6l+ftMh
w+2Jj22a2PFiIR659EzGV3dv1uj02AKhRPdHzECb7brtxN0ev1kyWMiKRM7FrBuu
iori/oyCKyN/bZ5f7WDF/3j89GG7rDZqYAqnsMJP2faxnvcENkW/tlsquMkhDIc8
0yNC+B7ouidg2kVulgb5mpMi7/RRuGoPwHEericuprqe9/tkGHHXE7XqcLVG9YTb
723Ne8GgwKolfrld0Oe657y53AfCFopztGr87ATbzCwucc9qudZH+2SwMucCUaS9
roNCIy8uZTjvJ1SXwGkfnEdRVWOqyQ2yUNI6Q/rktzMVJmKDAqEbra9KPv6Sg+by
YVcM+JOqIaAC9aFJvn9sqf6CgQnoVZ00csX84v8dkF91oumeTUMaLLPzvxH2IKAR
e3U5PvTWSEiRIkgsKRUxIBaQs44JDhMMnvQ5BxoZG+HneKZeen7ZTAIi7ejCuU9a
WqNPPWcfbYgmo4Tc6P/Mw8iJXIP+9O6cmmmiUR7pS6CX8rtct2u4jasMoA1qJbJP
7l3A7MswNA94Iue2GX2JKZtTXa9aHyUWGF2IOIUfNTbTPZ0GvPDuXcggI1i2cUk0
9GAVwxXYYcCFsV1RztUrRxP7vAI9nLTUgciZmfraLLgdmJ/iu506tifjFx8gtpXh
s9LmyswL0kAhWPL6zoDVJGvt7WWMEGSUpdSyxSQJyfuBH5m97/PILrirOX6E4hcR
1boAxuDP2msHiGKjjUyCRLsrMmtdKYyF9l16+3aPXN8VSqqwQzae2YRwOlx0z4qx
ao+c7AxTxJNxSs+76go6jBZwPbJiCPgWeLJGCl4mm0Lu9anFwYI/Baogc3F04t7I
h/qvI/qDi9UHmVhS0J26MqAQZzc97ZaeffJfboo0WiYNe/s4PXMNlAT9Dn7mzU9x
+WkJq4Wny/DnkSEGRnZtSl6xYoVURVsaC0ROmPmFh5rIN9q/hzFdt6OUYH8PLMTJ
SZQ1qS1NpYTjz1OTwmtYxBDyi5O1+f+icGBsVAyaIvCctA5HjCoU4fu5xNtGDvXO
I9pJ2eNwrB2HOx6UbbWe6qLjAY4UxmgvWoFGNhV0D6a8xntkAPd+ExW2xcfznjHo
nXA23Gt4Of4mRQCYDhcHgb2YHm0Y8+f2W8qumnyoUL+V87mGJ2ueZEaREyb4puby
9AjZHHeYp2bElIKV3KsKYHBjYSZqTpxtYe59yUMPXmGR+sg98wpQ9jgFmK6t84q/
2hphc68D9k9csMoquO1hCCZqcpO55vF5HRpm5/wRK+qVT0TwIadtWsO3gkjeSaGW
BxbDJmLOQ3X4GKbiPihMyiubVEwmFL+2Mu7HmWBlAEtsUbwUu9pOXT6svGACcxEG
DfBs/QVPij9NiwhAASX+1ZOnKtH8DaZVyatcNBdhLI3J+xi0j8IRoJNCdJUYdpKh
HEAd5hDoCiNAmJNoCCsmRtdoC8CXL8Kxhm3K1p2Rt4AK2SIWoaq066R3kW5Y2OWz
kMw5bMl+ss0IYgQptwsEk9nK4c/mnXuVQG7Tc3l7x1Op2kCIAFQgYU+cA0MbuwJd
F32p/0hwQXnsi9XfSQU8Mmkrq3D6svWMc51mz3n2USiOj6KaOpyhCQaodsSSAq95
8IxPjBFC1d9nGiBYT5117LahDFtEZhC2NnsFbq45Zmqyc4Qv8nWnjy2F0pmpw2RI
7Q4mxurFRME0O5doCXEGs3YTdP1eBN2InTrEkUmwTdQ6LEQUOHmkTYrOI6z3nR/F
mBTRWHG7LmA90IckK/ah6ivnHbT7r1AnhzX2RqBrXLmHsELkz9vVgk3UeexrbZMu
rP3erZHB9gxc3qwaENIVIQEdnd7z8+zfoCkZh2o/D9Thv+rgVa0C12vZiSrPgKVS
33Tdr0TLp1S5AHVZR1xiidCq/CYYj/ApDbNbcot0drdQdA4BTQq5ZFBAV+lPDnhI
PyVef6PhKNAkgsh6y9IfcrnFB9K3HuiraT+/YeqplA+/2dhJqj6BzQ6ioj+SWiXk
EFvIMO/aRgsSja1NACr9BPhGA4enlWAcAOQ+KidS/50cDJyr+Ohjx+mIjoGK89dX
2sBNZ6TjB7Pvzq1f0n7wHcwQwcxHRxUo/RtZqf9dfGEw2KAF0E4Vc7h2a8J7O33v
3cpSkTvFQyNCLWvGqwsRDoTISII0XyNb8FYiUpp17AHF377QG+2j+YifWXpnFi4L
NuYmouTRb2Ledc6VYwHZzNR5vG4UCSTfSvL+dGaO2SxsM52KSGpb5UeO+kAROTG7
7OZdJHrqV5tHZW1V9NNyMlOamcwPezq+zavjPk0vBXpS/yXm0MZR70cQRAuTPCEU
kL5CAXNFD/plG8B/4ioG8wM+km8nXl7HphCppyVOZGnkfVmoJvBf9RGuf4P6Kgdi
PTcJ/EA4L8iRH2GRuuLfImwnBzPcHV/RVBaSkWaE8lIj7+13D0X7oWMBFyZxbmti
u9Bo/5HlyoasJiK/L6Kjoa66+pq4xwh3Xc0q27Cxb8b3OkmIK/OXJOsPe9tEDwhs
ODMFqo6EEtB0TMT097ipM+8KFe7iqxT0qtpFAaZ0EPJyPwYqAeFE1hZvqlpyoyEU
cUvYnVIb3KKEe8W9famnCTblt6HNF0UoRhN/lIdqYwGejPMsZvmATEGsqRTMDaN0
aj7jg4scDQqfV6W9o6D7uNfv8W5viZurNuK/noIgvewEyt9we4LFYkkdcDFS/F2R
BKEce6BzLeQSBpZBsN4R17M+dKpnxGkdnR3sil+ZpBfrJTPyelTsEJOFvYyIg/ly
eIamOvDuaR75+7Fo4RbwybXaUycqLkyvoz3rJNpIinaVoHZcGTxLTuG79eZlqCjA
HcChuWmLMBaPjh9whV4dLHfciEQuKPPWrl5wVuoiC7kSqR3ugM62q288lAvPWJBu
pYhO1GfNZuaxSL1lfsAkWme6SJFLazspbtkPOneCdqDvNaZHiPxc9lNlrpZPXvyE
O9IEzV216GaqLoAa9RywdX90fb95T7Eg0vdai4UuhTHPcFdhuraRUR2L2WGMSHbC
vMLVWCaGXZ8XPDZXcF6Dyk2giCa6gpQhqNMU5Bb9TIfOpyPl0MbV++g5D9j8nFGq
RG2dYpAr5Z/7O1mYeC6vTHBLiQKom/ao5x1sNnPEscHsyioC+CCjLz0RHeNW4/Jn
qETU43ps0S3JOQN5gJeFHSuy0a0Ts4XJok/SpNz4F2Ngj2D1nhHbBJjP7wr1NU96
P7UcL7Gbn1ktsRGsTaxsNzoIBYlhiYm+Oa7yPzyrkvlNrhOK8gMh9bPDLKj63I1m
J9SorhuyQQJOsEbMhB2f20sZWhE4x6iNuWNsOtCv5wcv+GvGl+9aQKVJldzAs+Yj
rMb2qKGt5sDPzZIQAW74m0IsR/pdRPposbzD7RrBV31xXHIWfEFgu1oeQwUXBeec
kZNESBi41thz0KQwC6H+0DUO35pYHB6AS7XHNiUKZErft82fe9gfI5MIupnfFol2
wq9cL9yyvKSZc9zv+lA7AvjeEu7JW3jm8vgjNyQvy+vvt4QW3f/AYYZ41xdqReRx
BBsic0/0eeICl1dBeC1tpzoXSCQvsIdo83ITTT+iqoIBgoK77gqtgqy5Sn4qNXP1
NWMkWavXhlIGcleSdDBVCk/M44Q2rMws3T7MB4Lu65Z7U+CM0DTz4280RkMkCj9K
NsMKoQQ4rqCW9RY9JhpwpADBixUvsyDkvMajpwYqf9TNvucqFK5Kztlaw8zv3uaZ
fGki/NB0l2rB6ffPGjxD946s9qkWZ2FTihQMRclDDvu/SUD2+xDh7WHz/wpjjcNe
vUGGdIpvfvQlMcJ8bHvPyITjAdAFo9V5VeVqPr7etfT1frwXBhIM/+fAEpOPkgNP
8JPUsUAtxEr5ouHq0P2lZ9K869zUemHl7x/qHySoxndtYEutrEoHeO5TNdPpqL2H
E79WeIeDPqIVWpVAuRYO0yjSJKCVjOFljzis96/Sdx6wVUFnGpDZ2gCyi2+zxbnF
JW0ZQ174e/3J4WTF+Ipgt4EZHR6KGDpkBKUDl6B6jM64jhu417/3Q7TUAklAg6qy
4AmsbyK0MAgFo17+sU14yHHZMRGPbBprm8llsdhtFR305nJXHxqBqQlK5b9IR1wo
lVMsN7PyAR5ZhidcuU6JWm+pNpq9+PMovanVAPiyd40ibwuBswKYtix67hiSTwjr
kjPwfy+V6kosHCZfHLL/uH0tTkiNObqNvhTqi0DEO2JEibHGaj9brh/cZ/wWx6yW
ifMVdsY3dnQYN5C5YFmPih2LSnXAIHpdQLrgAUX8uwFj7e2Pc/AETgN5xC1hSqh2
ry7PQaUV2DqAGkNWWsw7Sz0S3+TH6FVf1lGkFv6pOxxNy2FVXneGyLEmghdHvvvu
cc/aEFzZPshPkP3UwknlXoiDBgde6TGPlMiYtR/ctj1Kh9dmGxmaBqUe290sOV59
VSchny0I7qKag8a+dHhAB6c+SA+yELjUAujAnbA7KMqw0FZeDBOqgcj+6ybwaLom
uWRHbogf+CQVMB8ZxOwTBvGA3UgqLLo+0IEwNsVjF98jVVMrB0o1siUVZvj2uh1F
+a9JtXEhXpI8SKBIV9w9zXSWK893WUZhIPQjRFXWgFg5LnzQjOaVxKRX18UgMHUl
STSskQ6RnY2CpR22/UJowssQrF3k1Dv29U0cHJ0BiDKvp9a0BYa4LDTAwcVoMhJO
jUnX3gkuQ7IDEWZ0Bc4MP897tkzpcFzfz6GZMc25xT0x77QNviJTzFcGAt/RpO0l
tRPpYtPXM32OIZl+Dwq9wjhl0JpY10+zdVCBtt0pJ9HfxMepcTsjLZICDbzuoA9r
20k5ac1HoXai36+EJf22nQsp+7BeEArC6T0T6G8axKJ6qaP8z3Alacrcx8gwpVP7
QVub8TRy94UXdescoroMHyRUEFzKG3njd2bsHBoLWyu2iWptk4MthMLmw3y4zd15
JG2428CB0/O/pxf1YSUm+QJSgF19PxbaOxTjkB4eS81LD7j+1VJcG4Hk36gVL8gJ
wYwHC6EjV8ajApxqwb0V4YTsNEq/eKTSXoVp1YACQoXQGdx6Bq2MlKsKFiIKaovK
OyvjWRrACIE6CSUbeE7uL1szeJRRGLc/9SGvUdhNf0TrQGzwezgWL1x3MgWEUwsy
rFqMhKovH9n/AQ8UxpaXFpKPIDaEA+6mnCoKfqnvgcJVihOYV76ZdeRpbKJsRYyU
hmfcGGc9bqOp8mYiaQv+QW2Bww6y+/0qFMPezO6J5X+7CcodJ0I3fYt6gJ8afxxJ
69BL0UZSM+V6QqVEz8JQEDHeKOOVJOnQJuXRrRDmGSb9Z03nrJmumrjyvrs4tUQy
0Wf7OGu/LbrsLBzolGMRpFGa1I1lhlybQKAOeo2Pk+KQm7OQRdQijZ9xOol6NkKK
R6kBc/RJrGE6XpfJ8qh+COmJRhwOtza5uDgZE0PtHtodWlDhgWp9WyfzWGb1zqiM
/VN6teaBTjYTVK/VItUKfyQIlayeOAa23oFk1rBm54au1IEwSHA+uViDbqQhGyGA
yCBhAaoJRmWQTONqjXoUsUCN0pxk9kLimVC6suVL9s320O18Et249vvdLgQc1Om5
JTXM3VK5P8tG41gn6hGQQNXyL93gIKjYHxruVj1gyrsV09jqIoea43WA+VJAlUX2
sc1u/YBEbpSbomMsz5WwjL/pTci0gHUuFr/UfEOGezO8ZhLQyJ+FiWPex8N2yTSx
ZqpCI9xZcesesAfCef3eKEHUJSuX/4Rtz9xd4kso3Ac6Acn36sfhG51oeoZQHrgO
cJilswP8vdh0Gp13WgGmb0JYi0gw1A7yGSKBxxKVOTcQ2t3SryrsBCLhx1sMwK3I
yfwTdlqwAF5ZiEOb38xLib3hTqbAnVewdF3gV1UkxONC801LaWm9QNoXD4Kt8N4D
gK1h3hFjQOj+Hkr+C+wpH7Q1roylG7aR+jRdct7lFDLE2bvBh1Da0hkQmt6gKcVk
UekTdjczlFLQ/LrB/GCVCvmfX38358lJfTEUa+71pj9AQ9/z8Oaj5qZMHr9tnAO7
vefu2YAz6kssiOaMfhHctATNJFmmp8uka5AvCdpE9Be3eHYTAm3GM0Ez080y386r
sN0SHG1TcfAlxsSbq/ez2AlqpMdmM5flMvj4YEx7TxqFX5Vln+27osDfNjnQv1hu
HhTdtruUHMNStWobFwuexW+GYzP3lKi9VC4gusf2P9RZExJRNpTQN6QBAqEugm82
gqibkQ39wd4QgLZo5FatVcHAPn45OHM2h7zfzRzFrPZiFgaJnFNgJQOKLhdu00qW
0K5FbpJihMSU/YBTCkqZ/gJY/zPJ3eo6KClqmTuIVI8QWBZOO9gCTlvdb2eHbpHa
skpWhEFjRdNoh4t6J2iLoH1fEH6dziXpFE8g1LTnTDUtCHks3N+3Gy2MZfKLi96i
tCVtIxMBRPezyvHs0haZPzBO+UiJZmRZRLzcP6ygbDKzfVnnaDSCiWaTR3jFhXJY
27jubbbrE04lDklefdx2M3Uy8hC22VLpIVcmBiYlh80XHaoJnbe2TjjqvrWyTbb3
wM1FZkoM5YZtPzJmvmUA38pG6n6lxl062mPKrkiiXuTxicuhPG/DA/jlUnrc86US
tycdgijIzgwf2TeMYCtcTMiHHjJTJ8pkr+fCJiQCTbR/O36IOzCHLN1t2ugRyHxx
XA6Oq1PEoJuojisUEceHGKk3K4Bxi8WHjesOPjsf6WWJUwhwDO9bOcoMvnNcywnB
rvT6w/loXLzwgXFmaBVnkFSvXK5SgF8u64Y25iGz4KgfNOjSpSUbg9rVxFlq4Fh9
LOhutrFBfbXnlKRSWTeB9PIInSGTb2WE37I/nJIdPAof+bb6F8lO5/n16WWJdfsY
OrgexTNIUksN1yLtubpAuHiFl9Mg0awifT8W125me/qNkX7oE9k013T4n9WaBsBx
nVt3xGAOxELuVS2damGz9had+MlKyxRHuB+259eq9gJaoDR5MCvU0yD84tADgW5+
iYiIwttbWlEusOrp2ARRuPgUasjdcDIf2r3lz04bW81pQL0yneTGM0FgB4hpOf59
4hGLSS4fOblvddWj93d4afugMzcL4vwBNe0ttGIASKM/B9JhpBROYWQcwSzWFXsB
sWES0U14zIm+VaGTHXz/AxsvSaFoSjfS1ztUnpelc2ZSw7A3VZOKiI18F2gxPbwB
Wj6E4Bc8ro9umkRTCBJEZaU4gx8QKkIpEPmwyDvABHfcgqMZPgX4y5+qfUk9MKhe
KOo9sjmwq8hs8eerr4FABPdHQw6j9rE90jH3tgY9yUsYXtF1YKjdchDzbBO+F77i
ad9K7oNLh6LR+aLRsbEbo5vOxQk4bmSAaluIl3qTNhgGelB1GruN1R38xDJPVmDF
UvJOH1wyjGow9UvvXphNQf/lOeUiX8PquO+FIs9X81cPS7U6JAeyVSuFkarsd8aN
44bQEEhZL7GqfldFUs6vgiz7UC2mapIC3jYh9fxlWHiRMUxbsS9Ou7afPfFTC+xE
/AGAfyHm7WdmCSqpAAmbOyZJlQMZ+WM25/gK43s0q/RnPc6FTHwYxc2EaA4BEW/Q
nlhH4lnDhSEVg1ltX4ac8N11dgZDQQgqLR+7XpoWhmh3e+EQx5FRXO2GpkjwjIRt
JdI+z8R6oR43tURsgAlkfosGgPP7NHg4kapoq8u+LE/pOOiM0zu/Znaa6s8xkhXi
SJAR1XPdmvTqEamwP7at00hSQLnPbvJe7agMK2n6Ub7UskpkamEBhxVEiFCp8My+
oTiY8MJMSBPG8/w3v/ldf/1/y5vwKdcFJliddUueZ3XWt7Gyv5ZKutH3Zx61ox1a
tuVvFqyIXYcYxNzqYzrHv+FKbTIPgjzSCtkLFhGdOQ/jLa3iKuSEB5PMPitD0SKE
XBHmCa2DWEn1rxXfDFtHkRTDXdI2nOS2vCrj3azxe4WQ3aVR3i74QTBG54NJVfx0
usyIK7oLvAmAnj8n7Rsmd6MpYn1KbhEFiEF90FKLiD4/IhUPbZIiZsO8oN17aZi+
5rfZa+Nm7OVID9j2vrCBytDiUxTSK0cNABHa6yrMaZk7DyLygpZW8qbGKVH4Hps3
F4uiaS5O2rhicPPlv5FDvkuFa3bY3MW8jts0EdNS940+krsiFjNSbJm9WtQJCIhD
KN0xPAXmjcTOGVbS3lE8jGusz9P9HciM5tcOxZikzIVtCAF845vcE443qv51aQAh
Mg9UGDbmdmPNroSkbYJkdnPEBPWRaJ9fucBxdLFknLCVOn8oJas5MEmwIeJs2ykl
bF70alZmgB19Ju1ePBXj0tcJSMAQc5jASbXP17lXoivUXT9uKkF0qPq9buROo+5u
yGxxU5OBJEsLYdFc3q3jRuR2RL39JjIZLPMXYPjYClry9Y9L4A495CqCMaBQZnIE
EdMhADsCsKL+R18bB9QB8t3rPvwPL+0sQk+uqi8yF6UvU4gC0sH5udQsXNAl6uCx
+4psU0HKUGpmOrUnawLftYrQWVhDhsymHYaQX7KK7xSQnfhk0jnzt9oZQvtSOyLo
P2QIvDVTf2kTGw6hCdTyqUINVik/pj48du146mYi6IF8CA79ZMFXv5rrMEYVar8o
hr9VhYb0YyKgYOoh6XinuY6lKLIOtO3V9A04WdKg2hYpLbKO6ryAbD5Eu+dE2c9U
Ea5d7KjoWmPfpnoTO1H3jCaQ3kgmxiJ8cf765mKRWzyMDzmbAzph6PWe9fquIMKT
lVrsG5/C6nQbZPWJqyBNNqyeOYt95DsI5WxdrlxXKQVh97x18rWAZOQRNlezyNa3
iItpaTyryyLwrU9o0Pg1xW+JequdjTykyW3EEYU4lG/IKm5DgqKwh2+rlwNNCgWx
X8uB/9/EQ0wn+AFUQOyuhAf5eE0niFu/Kgr6soMaCmbUdzteJ6Q73F2Kpnp6DE4m
uRwdE1uDndpV594XtXPl6Wuw+OyUniBQcp0Fl3+eN5qCCMQE1apzGT95Vz8rZ4Qy
cE8zqyHQ78EljrOOrWX89Pv1JMcwfCNcmn2jqZtkoWBE3FRCvS+sIDteldnfJ7nl
mDghEYnl9MgkY6747WwC0NQjgNFBE2OjsrJtiAo5TIvO2V6IMtoiBi/7n6jtBsvj
STJhYTcAhI1l0BLjdTrev+7VV5isbjL4dUv+N77TbdGUwuogiHn1Vpez/Nd7rN8P
sBopW+43eG+z7HfSbtnbK2+nlxdisS9lKJMRVohceqWALp9HypcnktiRD7TdPaCr
KZtElb088BhH6UILT76XPnX0YLJztJUBjzrf80/B/xcxXwWlIoW5Hzhyd2KjWppW
evuylctv24OA4RyID3RJkees6N4N+lrSLR0iB70lW47ryf1FAvBssdQ4JKvO8WlN
`pragma protect end_protected
  `endif // GUARD_SVT_AXI_TRANSACTION_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ZJdSTFSpbvkvguBRGw979N2U4ejyxyMTv6KO3V36UdHGRk5quoygF8DX8OS4AWf9
CQh4HZm8lvAlIuiCXvF633fqtqlA0cN/v+1Aa8n5ybPUoUfgdUBnI+yA7ATqSaTS
54G5ZbLuqq5vaQcJ/MSEBTt6+xoOuLL3PIZMS6fOD+U=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 520916    )
SxpO+eEjCdF4A+4PujAUFpaK3BwtDj8C0IjZUpqDy3gt7WzMFcXrvfQOmuIr5dlk
WylcoDPjv58TWWPVM3+omZOyZkG4eElpwy2joMIqlR9R3CAxujiOHWiJP5egmrNZ
`pragma protect end_protected
