
`ifndef GUARD_SVT_APB_CHECKER_SV
`define GUARD_SVT_APB_CHECKER_SV

/**
 * Class declaration of each of the error check stats instances using the
 * `SVT_ERR_CHECK_STATS_COV_EXTENDED_CLASS_DECL(stats_name) MACRO.
 *
 * Each call of the MACRO would declare an extended "svt_err_check_stats_cov.sv" class
 * named as "svt_err_check_stats_cov_<stats_name>".
 */
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
u6EFGTO5nwdNnOqlbj2y/NIPZkj4ORe7PjNGWNsLqTovVTjnNS1DAo6aecYCic+v
6vdyCnbUJEZNWYRGiyuHeq1l0F1mB+XxWVNELZ8R+usrm2nJy0LSibyGCbP+8SJv
w9y9gtUpP+8tZiSBARH+VewPeFQ3X4V8s0I9NPXg+eu+cAZbv/JFkg==
//pragma protect end_key_block
//pragma protect digest_block
XEQUmGKQaIQflWUQGlgP9Qvz3AA=
//pragma protect end_digest_block
//pragma protect data_block
JD8rg/qvyasqDkzYcVzRuyo2wt78JXhfbIIrYdam0z0ZFMTyo5CB+kbsJpkDz58c
hT+wHU0ZqKOfNXI8lgDYocd9ySDpvAGlixYPIxlM6ftzz6OgkB7aCMgEEneRSzhf
Tz8E7U3cYX8Zfg0cdfFguU8TLwq72rpq+KyyT6z3JXWD4cIGy+Z0wMCCGAfspdVF
ktBw+nU27v9wDlKt+3SITNkB5SehGlfAdFq4DNOoO5aJ9S0wX+tZR2HEFKZy1UUr
6OBWRiSOAI+VGk+XpbZQE8B2bSbygPyv8bWGQc17h2H0UUdTDf5zBq+ICZykS9ur
KtNDc9X6+DSWvpDOWCx7o5KyRgBy2NsTLTp/vWaI4WU+11odVHgtRL1zUfn5sJCK
M8I85kBi+EOkhFD6exo8iaA6WzoDE0gHASAO0w/S8n3d8cAubPL+RyMZw5rrO2km
oqdN7PKaNWHVTcrLsM5uyaDC8x2GOzXzz1Zclv+uk9842EDVg6wli22Qz6q6ng+Z
LUVixqmoutwAZqZ0Ft/zt6bufhubhnOL4cr0eIeeaCQL/HRST4ZFG2zkzktWvRRo
rnyxV/IBOqBaxfR3r7X+84tllx96f3DyVAsblnC/BRhZXbAJkn75IfVKNpoOdn2o
/W1DukQPW0EV/PklWZ00P8n6NRQ/Jo0eLqg7IU5W7oUAO29zJ8gMEy8owUXjfZ2l
yOwSzC7JK8Teu++G7V2whZq+SaP04EWKCn/yqKhEF5syfrMjbZiXxRbJ2lil0pRW
HURhFmIOU6GRr6+z/CfbkKR1Rd+6cXn2vzn3XLQUuAj7HOupqoA+0e7+y+/rc+cU
imq30I2vlTp1CBihOIPBOOc4amFKLZ1B7tCfRPtC5zmxann2hT8WLsGef7tQHu/O
sIklH8thSn8vBXzkz2oAujUcWW4CwYsBv2hXtoPwC95Ueu+7XAO8YLsG/DBCDPO6
/evaYN8szSq5+GOpKz98EivI4zQUGarDUXyQf0WPrybEjnth2zfeJg142xCmkhLA
xKeub7Ln0yXzTtHCuyxqM+2uCyAn6xjBlxUUWUGH4WaSqFHUpTik4v6Othjx3XhZ
cgFdfSCQRb/7r0qlq6ZQDxHJ/5JgwvXjQfMS84p2zjtKbvEcTVf0xefDWrRgUXeA
bxah7TW/TPRo1XxGKQd8mD2b6f1FxUYdsrf7HzsJzlfhqiMkCN4dCqEE2+FUNxL9
SkvNoBvx7YoiGNjggXy4WuiSYIXwLCAmoEAx+nGVYNEvzDrWRcDntEDWvR0Czpye
oQGDdeEmCnU/OAPMyiyHev2xj4RQmfBcSUFdWln0yH/tCiLEN2MHQTz/m8ZKDuPJ
RLfBH8yuhscwSA21gP/bYqABLq12kGYkeqQ0kT8461YKK3CNPHJiNRXC9VkSDO/J
wi0AydbnZgnpwCF3R3txdHUyPTf5bMF/xj2rkzDyHVB4vC8bwYuy+yGjpBChtfbs
rillSKo3lXGp+5QDToPSU8YpkAKyp8pfqnVjqaIgy3ttHtY6yRW3ntazrGGAWw2a
Wyhe+elJVJa5sXKGB/LtYxfd/PInLZW+0hS9HCa7JDUQ17Y5hFurKzuESnxt033z
J3UP9qrvVIOD+hHN4xVwVfVO6XRMdvjjebuiczZO8fEqmGAxBGB44R3j+h1h1UXY
ZguJFlIaINPoKyUhqKADhRQ2xr+OvH4EqY3t4dg79Py4Yk3IqJdmU4jtaXIt2HMr
pyh2Va3/TzdSDKT12Xi6SFtq9TeQueuj1xColLkJ6wlWU8y7lO3o1BwaRBYqus7p
ye42LtnmJ8jn8RgC799XU5Z9J/50B9xZ6kc4PECsMVh6JA2DFcIIMuSVASakiIGv
UbHYoGj7Fh2jA1VLJN5TuXLNnHi246iXSaUlVc0VKKJRFDDkv6XlvrBTyk72LFXK
8XOV8vgOT6TWkUQUIckjzGfZ+vrxQZ1kiXSGD7Ld4RCtAkiCQem+R1M0mxmM5jLK
TG8CvHMwfSL7j4ygRQbm6C6IfSfrgBssvtygdXGH2YnlN3yW97F5SCPPaS9pnXh2
ZQscAuL/qO4Op3yqLqnN6rtCsA1wq6wR71jIG5t1lBqsgKAzXSHSrOpu2PfIxWqb
ej/zXIUmqmkot2QtWKQjE8xddnGOTr0m+EFND4HtZhRQ2ZOr9VKsFRoaHKyHMFaE
s1RnhE4qLhmJQaB2WRieP2gfQ/FYjTcfX493jDhkM+yVZ6kt3DzEfVV+ra4ummNK
lQecqNX/sosSNH2p9x3YaDH3AkDlrsZ+hieD01Edq2ClG/I5J2vAhYjL1Dy8LLGR
ZTJpJ5Q8lVwEvHh+0MX6GpkbSdvJUEVIvof8VXbFyxB+uV6OJjwpRoAAv/caWJ/H
uVSbXCoEviTWuTtacX9PtCRSupy10SDCg6RiPmvEvU6cN1kdzQ22WqqR4uvaalEq
Rfu030LWrjBxU0IYysjRu0uxXaReLO2iL7GqoI82p5vtMdXx8TwfM7AQKQlhJ0jV
UV4/LyXZMnKaSjhXHowKgjlY0nsn9W1ykthPySYXQksU059ZIFPvBFyUPUDdRkpZ
RRALa4t6L1GlaaahON+RVLAvDgWZtkH0bedv+cN8Vjxi5yec1l2qsNyGgaJVjQkg
M6KAZufpOWvI671rx7W898CUT3GvcFi7NQYDI1mKfutiHzOx6OQKkQgEQWp8HECL
1oH35OFWp1lchUDmLXkgQ7bS3OkqRDTbU4KGTIYshLmJd4X0xwEsegw77b5JzSpW
rT0yStmP59AkyagiJO76uLgpW+H4gXEsleWAtGnGFvdggAg5RyGrjpjNycFtakAA
/+XAZlXuc6jRsnMRD5LAG82w7l/o07N9gidjKJVEhjU1HWpliNqij9EfvjI/tzxb
2sjyS96Njzi1cLFjHDnCwKNAKpVukyPLmMsljXult7AXz3gM85qpSbc5Rt2IbcjO
oCGoiJwZsZsap6SYgqK3GWXE51QQAfKGUS4AY9HW/E7mClrBoDvYmMRQ8e6JcCOC
EstzrM0h9ENNJUyUZNq1JO/S4YmpNF9KMlcEdPAmEHpQ7PN3E5TdrJCP45YQXxWW
05jLoJVlMm6e7tP2TbVL7A==
//pragma protect end_data_block
//pragma protect digest_block
zhJDszRIAiW6q52kwuRHF85SNLI=
//pragma protect end_digest_block
//pragma protect end_protected

class svt_apb_checker extends svt_err_check;

  // ****************************************************************************
  // Public Data
  // ****************************************************************************
 
   
  /** Checks that PREADY signal is asserted by slave within timeout period
   * slave_pready_timeout 
   * Group: APB3
   * Default severity: ERROR
   */
  svt_err_check_stats pready_timeout_check;
 
  /** Checks that penable is asserted one cycle after psel
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats penable_after_psel;

//--------------------------------------------------------------
 /** Checks that pstrb is low for READ transfer
   *
   * Group: APB4
   * Default severity: ERROR
   */ 
  svt_err_check_stats pstrb_low_for_read;
  
//--------------------------------------------------------------
 /** Checks that after reset deaasertion, APB Bus is in either IDLE or SETUP State.
   * This check will fire if APB BUS is in ACCESS State after reset deassertion
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats initial_bus_state_after_reset;

//--------------------------------------------------------------
  /** Checks that following APB control signals do not change during IDLE state:
    * - PADDR
    * - PWRITE
    * - PSTRB (when svt_apb_system_configuration::apb4_enable is set to 1)
    * - PPROT (when svt_apb_system_configuration::apb4_enable is set to 1)
    * - PWDATA
    * .
    * Group: APB3
    * Default severity: WARNING
    * Note that this check is performed by passive Master when 
    * PSEL[svt_apb_system_configuration::num_slaves-1:0] is 0.
   */
  svt_err_check_stats control_signals_changed_during_idle_check;

 //--------------------------------------------------------------
 /** Checks if psel changed value during transfer
   * 
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats psel_changed_during_transfer;

  /** Checks if paddr changed value during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats paddr_changed_during_transfer;

  /** Checks if pwrite changed value during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats pwrite_changed_during_transfer;

  /** Checks if pwdata changed value during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats pwdata_changed_during_transfer;

  /** Checks if pstrb changed value during transfer
   *
   * Group: APB4
   * Default severity: ERROR
   */
  svt_err_check_stats pstrb_changed_during_transfer;

  /** Checks if pprot changed value during transfer
   *
   * Group: APB4
   * Default severity: ERROR
   */
  svt_err_check_stats pprot_changed_during_transfer;

  /** Checks if multiple select signals asserted during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats multiple_select_signals_active_during_transfer;

  /** Checks that bus remains in ENABLE state for one clock cycle in APB2
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats bus_in_enable_state_for_one_clock;
//--------------------------------------------------------------
  /** Checks that if illegal state transition occured from idle to access
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats idle_to_access;

  /** Checks that if illegal state transition occured from setup to idle
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats setup_to_idle;

  /** Checks that if illegal state transition occured from access to access in APB2. In APB3 state
   * transition from access to access is valid transition.
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats access_to_access;

  /** Checks that if illegal state transition occured from setup to setup
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats setup_to_setup;

  /** Checks that PSEL is not X or Z   */
  svt_err_check_stats signal_valid_psel_check;

  /** Checks that PADDR is not X or Z   */
  svt_err_check_stats signal_valid_paddr_check;

  /** Checks that PWRITE is not X or Z   */
  svt_err_check_stats signal_valid_pwrite_check;

  /** Checks that PENABLE is not X or Z   */
  svt_err_check_stats signal_valid_penable_check;

 /** Checks that PWDATA is not X or Z   */
  svt_err_check_stats signal_valid_pwdata_check;

  /** Checks that PRDATA is not X or Z   */
  svt_err_check_stats signal_valid_prdata_check;

  /** Checks that PREADY is not X or Z   */
  svt_err_check_stats signal_valid_pready_check;

  /** Checks that PSLVERR is not X or Z   */
  svt_err_check_stats signal_valid_pslverr_check;

  /** Checks that PSTRB is not X or Z   */
  svt_err_check_stats signal_valid_pstrb_check;

  /** Checks that PPROT is not X or Z   */
  svt_err_check_stats signal_valid_pprot_check;

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
/** @cond PRIVATE */
  local svt_apb_system_configuration cfg;

  /** Instance name */
  local string inst_name;

  /** String used in macros */
  local string macro_str = "";
/** @endcond */

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   *
   * @param name Checker name
   *
   * @param cfg Required argument used to set (copy data into) cfg.
   */
    extern function new (string name, svt_apb_system_configuration cfg);
`else
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   *
   * @param name Checker name
   *
   * @param cfg Required argument used to set (copy data into) cfg.
   */
  extern function new (string name, svt_apb_system_configuration cfg);
 `endif

  extern function void perform_read_signal_level_checks(
                                                         ref logic[`SVT_APB_MAX_DATA_WIDTH-1:0]  observed_prdata,
                                                         ref logic                             observed_pready,
                                                         ref logic                             observed_pslverr,
                                                         ref logic[`SVT_APB_MAX_NUM_SLAVES-1:0]       observed_psel,
                                                         ref logic[`SVT_APB_MAX_ADDR_WIDTH-1:0]          observed_paddr,
                                                         ref logic                                    observed_pwrite,
                                                         ref logic                                    observed_penable,
                                                         ref logic [((`SVT_APB_MAX_DATA_WIDTH/8)-1):0]  observed_pstrb,
                                                         ref logic [2:0]                              observed_pprot,
                                                         output bit is_prdata_valid,
                                                         output bit is_pready_valid,
                                                         output bit is_pslverr_valid,
                                                         output bit is_psel_valid,
                                                         output bit is_paddr_valid,
                                                         output bit is_pwrite_valid,
                                                         output bit is_penable_valid,
                                                         output bit is_pstrb_valid,
                                                         output bit is_pprot_valid
                                                       );

  extern function void perform_write_signal_level_checks(
                                                          ref logic[`SVT_APB_MAX_NUM_SLAVES-1:0]       observed_psel,
                                                          ref logic[`SVT_APB_MAX_ADDR_WIDTH-1:0]          observed_paddr,
                                                          ref logic                                    observed_pwrite,
                                                          ref logic                                    observed_penable,
                                                          ref logic                                    observed_pready,
                                                          ref logic                                    observed_pslverr,
                                                          ref logic[`SVT_APB_MAX_DATA_WIDTH-1:0]         observed_pwdata,
                                                          ref logic [((`SVT_APB_MAX_DATA_WIDTH/8)-1):0]  observed_pstrb,
                                                          ref logic [2:0]                              observed_pprot,
                                                          output bit is_psel_valid,
                                                          output bit is_paddr_valid,
                                                          output bit is_pwrite_valid,
                                                          output bit is_penable_valid,
                                                          output bit is_pready_valid,
                                                          output bit is_pslverr_valid,
                                                          output bit is_pwdata_valid,
                                                          output bit is_pstrb_valid,
                                                          output bit is_pprot_valid
                                                        );
endclass

//----------------------------------------------------------------

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
nSoWml+41xmmKoC1eDlgAuHc/l/214+TfboTo0mfluWKYmVMQ+t+rbf0w/E1i5ck
qjMUOD9RotodD22UCpGKW1ltY4RUH8BmkOcRWk3kJsfYxSaOYtLQuKCsuz7gJ4qv
KH6GPD1PUxyv5Bzq12G08YZ1Yn+lD86bPafXv7TRAtsU7XpNBzeymw==
//pragma protect end_key_block
//pragma protect digest_block
Frf8EWBK+itDZ8kZhGh7t7NbFXs=
//pragma protect end_digest_block
//pragma protect data_block
lBhjnxrd62aCEmSnDX0gji9pxSkvyZBEHvN2KKg/0FAcHnlNbBqb4aiS7k109l6P
/Z0KtP1MoyYZAnwveggla8YF7HglTTh10CiPwouc+JNBqzjoX9xL1YEHjn50wIjM
hIL7rQfgWV3PLUUVipf6qSY1NrfoW6kt8JYboo9c/5S3BXg7zLDpzr5xjOmWXsJT
gFZZX6pWGTVgMw1/mUFqdpE/TM8MVbfJJWjbzvO3XdT5Jy13Y+wxGRojlHI5fcEn
8Gv+NlMqwVbpYgAVDfgCXUEVCanN7tLvl7GDPplcjLjqi74yzDhrgBd3Ek2r9yqR
fJ6Qb1A1mecoFUDsx/Zd7XHxzRr6oMYnTXuOee86fyTo/DlhIv9pVjFcM8ZX7tp1
Y6VwNiNRXOCuxltbJu0jzvZuUqyLozD+PaxTAqIjl8omHQP4WkMKKqZyrK0VeN11
0rPyj6fJ+q1eLq4pGPy8Yus6Su7n97sZxvYUYvT58Jee82JnJirZNlCK1qoUKV7N
nVcNauEqOc9yIaf+YFjff+/J43bjpf98SnDeDZzXqlzpwpnVVZNTMtxFQ/FVeVYh
KP8FBA8NYy5qQdT87YBhkjHp6MxXuaadINOhgwwTH3fLYyVzF7Fuhq0YzbfNPPp9
9uv+Qgs+kjxNpoDPRZrI7MbhqRGRlJFWpbO9jpJyJcySy8cwO5R2hDT+OWQ+74Ul
8W1CWqsV1SRn7zZwWT9aw7CabLLDVL3fX1r4gXMRyaTXlQ9N45w/jF8819iwljRp
35IhzF4h1hSUJSA97+hlVgbb3XBiZ4YWNhFFgbPHtC2hD4TChwhFEimlNrcFDJ82
nQY6c4xQKXBuu6L5hHQI9cptd9d/weftOotzYq9X4CkpAGaERKVEkN8bLX+7eL1D
FIdGlJU/tHpFs4Sd1RtBbIySl2sD4XMiUcOZKVt6UBvi0q0M2LxmSwCRaSYg3M3C
G96O9Qq5HOaxYz7iAd1nMVn0L2l9wuESI/fOMecqaFIDVLwB4YcBJbg+gpd1dSVE
Im9LQw0mxopTZD9B/FM4NnogMXmMDNPyafqggX/RKSpvnBGnpAhSFcGws9DsBcQA
W4a5C0UNsX1RwQtrpa+ddQKDQVvH5Jeeu5gULL1EERzBgKKY349L0L3OkIm+m+NP
JuJm9gkBRZET5Uk8mR+VlvqIIxYEo27y4NsKfTNnYCCpg/HLHzK12Kpdq4kSZxGG
3KyV6g7v0yIp5RnbkzpDBFXinfXsuBBASLDrS02aWW0Fttccpnf4kMJLVt7Xskjn
CuA+RuoMa+nw95MIfRCbDCY+P2SPmHG/5UUyc4fUIwSX7rm0anUJcvUFDrzfpwtr
EnXuO/uVPLYjD+bWlPbMtxd6b6M/BPzd6PCBwzFTW9PdZ0L7/8jRNqENhn5VwF5X
PkQACGSous42zdF+oblnJv+eH5SvYAmr9ddgCQm6KowfnOu8B3AgpyIECdtdkLKs
W1OPJs7CB+AMNOYklAQR3YIb/m7iwo4gLU/3mVQrMiGdeoK6JU4sc1Ts8N/MJXU/
zsmij2cKywEAExK19hG0v0f2QwaiaJ4cebREIcMFuv2K7+EHU0TPmv0MSLY4RrAm
NOBNM+sBNOw/WKo69kXHvD26MqBpOakoAsL90io6lRGLXNAliAGG08A0JjuQk8Lb
sKfJ0tOm8Jhxz/DSCnEVAic4yUTP17AbWx2NPUOo0gCdl6n8bhMdqIaU7NZaLBkB
am+EuFgXD4Qlkoekn6+KjI4ypZS2YPQ+dR423W7KMfshDPV9U8VnOFHgQenZYSQ9
ZSd6XvRE7Or/pzffnhiFuH7LgtEFV+Iib3CsRKOoT6BoXnsXyHRVLsFFW6L8bGhR
rHBYnioK6w+hU4jySsYfaD6wEgHiW9JE2LLr5NroiWO/DxyXdf/5faGXEVOaRkMT
0cAu2bhjJLYen/FJGWogK9JTbOeSrnu1W5TBcprKkuIUAS39QtE94ofJpLwhheNc
A39/R9nrDHTCn0hGG4xPDwOWN63pezOVZ0ddPbrolRSOJK9NhuBztpYaLk+W778R
69qCzKNXk2/ZuYfDkIa1KP/khnA6TRzzXfXgGpSCtN4w8Hi1zKilYUY40nYz70aC
Fup28YGaUU44Q4Ns9nNVRhJqpHYuonIwjlhzBulitkiEE12R6PSGpqq1yFzO11e7
O6xeIomEpQQu4rv2eSD9flZND6QfJqs8In7JJOUTYavCmNSc99XbRN3JUAiVZ5op
Ilsb+T47V/Irz4rs6i30ouiYsucGxYDKgttJvk4h6rKZnYMD2+5Iolnsm+O3++yx
GBp6Ku1r/8EUxpTHjXV4uDJ2hvqIPaIMM9ASCajT+zKySVmJfAR6Skn7kdc9R9hT
02/GTLZ1RSOBiPSq9AwwwBF1wdrefbQm6UZHaZys/2RUSI3jucUAwBGf7lPTdtLI
nLcjmT6P5C6fr0ickNdtBjCEhjQNzfKjoLhePEEH4AkB+uonol5sZsqZQXml8o8O
otcyC1tUZ0RykbrykkwyRcvjqATT/I5T3tb6O61PEniWJaAHmv3TzEFYkceo0UfD
qqFVljpWWE5y3K3yFtlPTZlaziCWR92xb10gdr6RLR/in/hlnPy0m/wNf2VB1kbS
+XiDa0XBAjLs0I+uK6/QKCH3yD68WqthePXNgAojypyowVBgV2b0GNSb424ZPwVo
t9CwRjeTYbYjiwSRxNnEJdIMv6cypcRXmcFTs5s/7fsGk7EDiGD4iY+ADByAFb/o
nDLa5Octc5JjnXdiE00YUs3q4MrbVasn8wrdvEaZgY0biJCBR9aqxEZz0BSGfK0o
3cL8tzNFaTkNoKEJeeL7e661TcFhqj6hSo3RhMzGCfSVEYleRcMmUxvpXQTzcnsx
1nAl0w5UoxmK5sCp5dq6/vefbC7IK7nHoKAd24yj6mhaQCmKb2bf6vxf0rEAmUD+
hyihUj8n+/zA0nVTYkDgB/yyD3xrEvZOONBMSaSc8q46gLxLXyN98KMZDJeOl09H
M6r2zzQCJfUqU1XqsSQHAKttU2REOfnGuIkml300Op5sbpv6NgqOqmQ/LaC63gj/
S+62cRBEbTspjcVyQinWM67CrVyvQqlKU2G+O2GIzh+zBRfYO/f2kCdveoLuzt2z
2xAQXXmS09aMT4ltz1x9IqVzvoVSKnmAaoAnW/Evm77YSQ9zUeAOHKAbZeIef7ic
q+k6RDK/q+RzzKTPIWghkmaPi+N8dHloGqwfvCA+l8SXBaAPXflXDfW7CFmwjGuG
wKpW9qFs8a/SoWQRvKFukM1nor/jr4rlCh8+1ag5P4qa0bSbKoaVlQNhtFahRofJ
Y0ezaDsFA8ktJiV8w0HvFombvU7ttv+iwpJqC8/3v8UYTxIQZYiwa44g50mLhPxJ
4BbZOAuWe0A1rmrbvOc+NYXv1ywNyi2ji7W5owfgtQuP+zOHCrd6zwXJGifloRrm
Thg5w7S/QkESgJb27SWI4lDWyQZH74eldquVjbw9y/AxK4P/eGT1dq1xNQz1C/GX
S+Gz8wQoUbmT82eQg5R3k/gu+WUxcweEx4naKw2lhgvH2W9OFB0Fl8opFET+Okrp
spSFRdJZO76ZBH90urlEOYCPm+31vD//tjoOl98vb5u2TCD1AHYblvaUR99OV57z
xR5Dkha4wwzXSOMiVV20NA5k43uDO57huP1cNb+8vsNpWQ5vOHnE6aJJ9bjIXF9Y
dv8ptwY0R3PS3dG3feaa1L9J2sFd5Qo5Aj+sxf6TmAF2Y6cmnLG6nkdxTZld+YAz
xb33pD5GKukWcNg/pfPmAmGVAFjhxxarWkVg74dX/NTIMUirTZ5CKSgKgkn6xpUJ
K4pcNPPWGpfADWiJz3nyIo9HnTQVplIxtETrob5gLfiLSXt8ZXmNIWGFlbb6zrLw
njhk4EweUV51ktAhCuq90PM2voAkq7TgQhX1Z1B0AOcnHtW77mDuHCk0eFtLC3V5
OKYx8jQeTiCdLDqnM9Kq8XWr1KRjzEwlK1/XHbtQQDXpmED8K00Z+BD8HG+iZrk+
ubFO5tWPZyC/URrXKaWa/kMI6JwLHaZ2SaWNhYGmUpmGQHgndlVhE2UJp8m1GjO3
RkRi82AzwciZgw6czU3O4Gv2Q7iv81YppSqgp5d7zaIIOKx+fWtLWKxOg/d+6rvl
x58Dst1U2k5Yr+iVv8ymy5Pmwz1gMXvnveaUP61h84wyVro+LTrvjXDaSI3G5Hec
fO4p8uz08KY2F6loocEoG1xKvbUNk2JaPy3KSy+NZRDARC/0FJB3zFxeRMHtIMdt
svjzOsPbaoaEhansPkp0T0mj3LkSH86NKdBRF0ZXhfQm6xIcRBoFATYPjqbHJiyY
LijGP3JiXkkLzi13m2KoWgPhjzb27+lHnpu3L6gjXNuXp4duQQcP17wojain77XS
rRjH27EVmmOJFbE0xnl2zCDKMWofdbPSu5/9r3kyweOu/xiRe5Ic7xnf87nMGjeB
oU/wecrWDiMNL9qRpO4F5XMsnUdosRKsgqkDmxl7p8VRAY0ZmuippJHacYa32gDv
W5+sv/ZIeSjOKMTs1T4I/a9LKqauIflQVtsBF7gceQm7r47nx1kaMs8BAXcRSH4y
cJFRKRjN+1SlVIGGLX68m5YJyS7LHwPXx6volCtt1y0XWbK8mQNVXlaH2i6PI4Rv
KPEjCo1gS1XGfS0RE/xh+ezI4iQ0CDlAubRA46Ad/e5plFQd2EWf+ayKuhmqBnrH
XzixaMX5129j+EPw97V0MRMEVyaADpZ2+IrhkAgHr3ecVvxx9/u3nYGCk1bup1KR
BvdsnYOQ+wXJ+/JrUZb8x/GBkgFNqS/66NNbKXKILhrG5oaKao+OwDaGCWgLTzMr
YVz949AoIdGM6YKsFZdN+bsNt6YdG2erIPE37EaxJU2KWq43mfv9UepgtY1ljdqt
0jfNRNsL1m+DpdlhrhLUrY3bLV9xsT9dLTgQVtaQxc7Xz20WIsYpG9Fxs9AlhZcy
fOoEijjNxzQdn2PokXOkZYgd2Y7ycTNTFghjenyUVkZnfUIiqPr28JeJ8qjxY+C+
ZgRAuXro9L7G+4Cw/bRcMfms1z1KHE3MMHxyd1E/7gMnkvMpIUS2fVQ6hHyz5kxB
fa62BG/IZttANrJqjFUJ6Eq4fZ2ss+/y2UwdwdWCJGp8Gb+lZXFAImmJvLP7JIq2
y9QTehZBCcejyz2e13B2DrqAzvn2iDbkebhp4K2AsZylIxmLc0xOmHCFq4NCfw+Z
CJjHUni064dUQ3/IWaBTOjZswTEwZ0w4JWXlbZUWE3q4wFpd5U435T9jOgme9Myw
6ijW0PkaxHLB9DoOl7b9eUjGaHDPrpRI94Sa69BiAJ2kmDDdBjYTpUPG5aVIUH8N
FAVafAVr3Jdp6Guhb9ZoA/gDf6tEDHxvj/Xnf5SI9q9dzn/OO2fYVkJtJc0JXsaE
zW4xuM8O/8Oq8A0hXocEZX8OeUoKqBuK2veFAQLKRcdStAAVjbi9UD0P0JOuszIf
qEs6RLzDTA2iEhMUMqWMXiIjipVdSPE/faXSlkCKvDNuQIqPuCarc4T62tZ+q09t
V4CtsqEyaHD8eYujb/5Hy2ORuzgnzuGssWuCM9eP9U2IM8qDR2Bq1rCDmjZjM5lT
Hc/tK+3eolLqSb7P5zjhuelwk+McLCPQbNlUkp6NwJsU2ree3l47DIQWfKgVd8RG
RAv9RAXutBmzX/dAy8rGuBGxxQCtOWNCC/i0EAEdblEAH4V0zwpbklHBqvJRUYGe
bTGfeYmQkixoqTHehdIKE4PCpxUYiZfa45KtBC365Rb6wAOOfnAM82cXtRpU3upP
U6l4s/HfB2QvBDQN6uSg1/9JPl3Fjvv/jzmLDO5Y+OeyBUQcomi4wdbFoe5oHlQp
fmFagR2z0r2kGrDDsVOI8DRvAsxafrajGONwqDPy8sSW1va66G7AjGdY41rDc7jl
lXHjvP6p9utWpQp+IS8nIz6VbUCwVo7hTQnkwS4fNsxcK2CHGfsWOP92gyhHNxEI
y4uoi/BkHF+2UrW3G2h0h+2mfvPFOa2A3IvPz/KWcvMVL0GJh/oOi0/+pAMbYBT2
GsYbLhTgFYR02eDD6r3NiwnaQ0D1Xffa6cAYu/Wr1mRzP5F0aIqazdqBh0OHls6+
ploFgPqistmVfHPp0z2sKoled6PGfoOfDtoLmGKpiiQp27mWZ5P/2Is+4jBmasgK
hRqFEgV+jIQ+s/Mit0zp25/mJazhjmRUzSBMqXh2m48MZsUBXwSSYNxhyHGlVPSE
n7WdT/RUa1eStb4OsXLfwuwbFJJ7FCje7N037KpevjcHYqIe7cz9r6dLfpKds5Ub
iYLzgC3kbSTHJxigIIYeQF5iuhYMyVILLqKPoyo9Xsu+aQbfcOuJSj+H0RTvjOyl
OVuAQ++G3VoZYytnGvt7G8ppswAJgRnSnUbo39BlNLlZLSobOIXd0iP/AZZnK28Q
I3UZkdbe2WniQbL1+wmH8ZVAQuktiuiEn9gx9Q54nInPWiSnqyOsQwdpw6vCmPdM
NqyW44DQUjoH4VNDfXvtBSRQRYObjMNDW/YAKzADxvsQ4m6mTpKVVPrAfZlwwoDM
Gkm4vaZSrxAhIvMIQs5pgaKB2FYvnkT+5ckwz0R7+ZGOOlxg89XO+hM995YUXiAc
t5z3eke2jbMoZaDQUpEPdtB09NRWgQsuYQBoYkXVVphTTlSaFViSvMp/wmLmoX9m
YDdilV5rZ/+mZ1V5Oozf5bKmnQ1gMRqFpE9Tb9RFmnWtnPm4uXb0incAZ92WA9yO
uQgM2S5q8rd783shLN2eBQ9A8AVpQ7B2DIxlwKE/5IChrjd8nCAW4SuVfhsP02rD
WdllcdPks9KNdZRH/0VdGkLffv9bBTt1izPwrkSGh3FEd7paczWod6bNzOM24h40
OxCXlk+qq2S/YFSe3XdUxwwIRa0Bxv83mUYq0Yy/qBUZykkKgj66b0n1NhjyzN3B
J/R6/DRebx3IAYNr8r99u5XSpMP8I3Ow33M5Oqtk+EZ55T5CQDwcKAUv4uRydcs3
cNtUqAVZlhSmcrIviEr8oxLZIIFgu/Q2wuvRqKK/CCXpg3ytmWdHulxzOIXVvzao
wIQrWaWgNEcx7BPwXpC7REYF3o0t9dCLErx5siE93VrXg4g3wLq+AohAKtm5oal0
FZwssr9xKkwX0jZiVCodbi5FeiOTrx3OHn9ftsJCp7vGcFmjpau/704XqbXYYjh3
lOjBp4dyYD106PIdz0vH+IfQRA68bgwwMm0v37vc04Pi7VZsKNY4topIebpJIOzp
bxzBAv9PUI3pZJ0yo3ozkGXYiQZH4soY9sAsdR5vxE30b2RfRB+vJ2q4C0LgKXYm
PZfhHUqTTNNfaIDauG15HLiGtznsldVI0M9+FwT9qwBW3V6PlrjsKiHt0X8GBwrV
RscNDoHQp+SCrnSRrQSV2ybHC+W7qHIoApjNyyeJJtJl4td6Afb8MlGYj33UkX5t
zfhp63zP/Mck82mxjapXSPANUTRYu9NGgGTK3tRd7S3D/LY9pmW6DJ9dFrP4M/gQ
hsPvrc23kEbgxhaavCygaZ087TjuZTlHKXwUE9ttzTJ24Ols60r+ABAWA4wIYB/a
cVvPuPwgfpuSSR3gctjbPM9MYE4nL3WSl6OrCO4gZrJsgL51pQwhdWCTXOrJnTs8
ck61opkYBvPXVqTFWHza2sSxmJrTBVHR1sTEq1lDdRSQig/4aeirWepo9EmNUjG8
4qvoN1R8VM4ge8Z4CYEf+vc5QEbwnrxYieBrgIO/3yy6PE64YLWAe8S4ONs/cfyk
1/PGU3DmwAiS/aMKWtvMRqlToUDcREN45TSW+r4eUJQaQiWwPR2MKYSscySiTpQF
TzmLGBpIbwDQpiIYDbFskXRQ0CuSIcxiEaKeoChpTfxxOxBL5b+Sq3GuTPNqn2WS
tW7ZBZ+AznaYlJCZvGN4Byakuz/1hLbGeualpTNkv4GO4mTi1bX7c6v1S/4Hfcp0
iIX5S9/aZevQ0IMOVF1ujbA+XebWEQQiltkzkEVhDgpd/YSrD/5Ox0TZY6wZfkUX
COXcxqUf7BZPzU67nPc9J+FGshFEvXWzSRSMgjv7FSoe2KCGygYm3l5VsM2Ym5Pv
RcmzXQLTLgJs23/kVZhuxSy1A8Vr2n6PCrB0wokfvenKcPlSlcXBgq29GBvipcw5
Rxe+Mxf51xRaNqxsbuxpZZgsOC+o6J3WZRxZ6+u5waQsbaHSqo3+5Nu44PiksZfp
krUzHGiRz8moCs8xnwrmoCOqS29BPoqPQvRZnWR67jCWfim2YvJLfs2WjSy0nYT3
EesSXmONoTUWj7z8rBNr0nMYXyFMTixdyD7SRP90P5HnnxHHnNCSmvhbREhELEMK
67O3x0dFtniUccQBmJ4hd8GvAodNaAMgK9bep5Fkwft7fkHF0hl4g0dEfiR24pSL
Vk4cCMMfmr/WA5a98AAK+TnB/LCedawk+DlIRlbaQuqq3+brpXYo5h6LlVyEkGJN
w5j/E5k6fdLXzylKuZlTA8Y/mpVMt90W0aB/fa4Mi/q7RaI918SNDiGeI8S8xEAJ
/eUInYr9NpQHdRNX2gsgZKdC76tqH0Dxj/M1+dhXJHdSpSe5AxFtQCFaZtGzKc62
GySCm2QSWyWJ6/2JfMtiXUJgkEJK/urQUZaVl0LI4kf0Bv27zm93FU90L5Nt62gL
mer1gL9xa35i233jJj8mAubi3Qiit2jfW70G7tGjq4AfSbrJxFQR0xnG7PMxFFCz
l5Ai0Zyh1IROXgMYBCTttK819NhNp/O+eGoeLE5qkixZTfDaDiwEY1ArIA4sNi4n
2Jr/DCdCEKZVFtJCDE+Wp6sIjLxR7p3KoIsGef4dComVuuNzP04+GY5hKK49Zqg3
gmuKygqZaQPDtc/uBu50F3VShme6N0kruJTD2D/URPIVZAOwckViWJ3derUfxySN
NOcSaS/+crhWx6AmeP5ScRSo6kT7LCF1a/A1ssgb/q9icQUk0Dz+q8VkvuG11GFj
EXsyaJp35Ag874URltuPzrB5Y+GXgWJLUFG2g3MCWSDtrlVmidKNO4pvgJIFOJof
g4AE1C4ythMiAp2sK21lPzdBT1vPCOZeiU1KnxcGJrUkoZXVd4a4z2ganx6+/Q3O
51O1KMjFF0ahjmEI1Jv6coPbHbI1JWlet0p6HXfIDdT/t+6y4Ul2hvFVhVvZVUyb
bCQiIUBeRaF3Ikp0nCLiftftQDZjYa5F7obxExDll3c=
//pragma protect end_data_block
//pragma protect digest_block
A4w+74asvuhLefUgedcV4XpxXIs=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+02GHHap94QCkycQhbMvvhgQXIwYPUGBV64fj5kOKlK/LwqKr3y2c2RUIup4U//w
pkdOR44vpKRuQud1+NYCvRyUzfXLKoxBQFW7rVci+5mYzyQrU/kBC6NI/ranjfam
910jxtHdEIxxm/67NWcIhPUKTADcx4sQeLGbg7bQXEKLu5vwMHNYbw==
//pragma protect end_key_block
//pragma protect digest_block
KDydz84N2fCPx//azNYwsY2IIMs=
//pragma protect end_digest_block
//pragma protect data_block
e6MwY8KxPNXtV4ND6qjRx5dT+CX4gbrIMAFO4RIhNg/IidhocHvWycAQTPPTcP/Q
HnG8NVWfGJs2RCR9qcFtZEZkLsb7jevAYKXWreUwa9i1Qx4OLgP97J0NStfrtawy
MMIpV60du1LQp2gGV6kPqXkaYucZ1HpeB30mvXRsOLH5O/Pheo4BKfqaRDVDOblY
XHozGhHmftQX6oZqtm7XcEH688Hzb/4VP6Xd1bcfCukXPlA0zRi7Z/gObbOrTAsG
zsc2KQc5ATOOOa7EuOw2GECqeFm5NuLx6vKG1/b01knSZekOzSwLLqXwpTjM1hY5
Ahde0DhXgu94pOpK6l+DFciCOgtDnTiNioV+5GLFnfyS5g+smKTNJd8eDCKoJFpW
DH8S8jMuk0oI3+xzvayXQG8IgiK2+vH1PPbGnyiA6g8S3gQU2Ewck8HxFc6JwF72
j1ck/BGEhK9Xol2YkPcq4O9aqQINzWT9mGEbJtLUtCAGPrIyKYZOgwMTX5PU0gTj
yL4ljxY7pfhHJ6nO8PUQWOXitOhCUJVj6pnJtPn7wMOutDXuqWp2Mdotokh5K8QM
XEFI0Qsf+YvsE0miSocV0kxAUDXafnXo5680oQQpxEoFOsiNZrlbW2CevH65zJB1
f/YPNiVWTW9uw0p0HhQhPngxmFtel9Yh1Z03yehdTleFSTMFUgFLljMfcTxWM+xN
f0Lv5bfS04o9HGN2Sk1mf0JFS9crVStnlEo7ufSIrPmozwuwM5dI8ju1efR8bR5O
pcukFh4DuM/JnSYxEl29hBm86QqsZnS8NUVnt4QPXyvIIPbRMufRcn4WlYEPhoxk
A48laLeRxWKIos0wj/TNe5S2fqIn5dwhP2zh1H6jlig1HxOKJqBT1N1aHdH/xQ/5
3A5nXr8p1XpqHz9x2nK4PJqbyMBF2/afnBDjvL8EdWNuEJobtUgxKPmfq8GwyGQ4
7l+0+Yk6c/NxFc2GjizlwfPYfEA+xVSa8HZGaLDnLnliGgkAg0xDkcBhMhPiZg4F
lr9IFRugQY8SpLPc63nE6I12J1AkfgVXhgpqWEhHO1gSkR9tv1H5JgWs5AmIvdFV
S6knaubq8zqVDaiT4zwBUzIl8w8uW4OVnoJH7YwG3i1kEPHWuwJbhL266VJWeZLJ
hptjhJ85dBXJnxF1JiZgbD7yKxe01xd1QqoSeS0DI8qEqb2RXPazmfJkgMBg/ELn
qjo9kmXNgtiR7gv928h/Lvv63bgkrsoL0pokYYh6v7TWqPOkVG0azcP3dXsasBd5
DnJcgXizov4PN8O5Zvixlr3wITS/CG2pzpHeWet61hcMhQvgiKs5xM2vO87mMevQ
sPUxcsDjIUm8STfYGLSxHerKGAzUMLbEh5JJZ1hfUrY5LorJagqVrfk22A54PYY/
E5UX9FhyZbkbUhYxcn7MQIG64KFkXwVdetMNGbXxZAxEeQvyvxMP1DLejdoilhwP
WIzWPhZQJr6Q0rXWug/vPsbPRi6qcgpzoNun1x/U1xI/rD4U2oWASYtvMmFAW2aE
HVXX4rtUdhiwAVHUn5hT+3hRJPeZF71vdoBUgmKTz8mKohWGtFMzazZ8c3Z0VzSX
lQd0WWlLWj8Ebg6nJcjLLTgCabU93dxr0VmAaW9tu2ldi5dCTZxzGxKRyeTgcq41
mavkEx7miw103f5E+3KBGKpSS1QJao31MqU3nOUZsREpzmlK0L6zjvw2BAzi6Xji
mSaqRNvdKMzXmlMznvyvEuJF49HMQlskblC8ef/JyfB6katS38UQM9eH8NaKFFha
2g+4shOBgETjW6SKQNhNyrJUfeX0znwr6DGQWetYhZjmrvnmrFYURLgvd3K0ZFh6
yHl+N7iaNekp8v2Tkjzii8h8eyhRVoWtJX58ihS813b3/WaXaZXein6faTAX2hGr
q+ovDkH8edkl/aaly54mWzgQThO0Bn+JzTaJPyXi0/ORs7k6ST3i9e5gGfaG02EY
+VI7morFdd4A9EwCiG+O31t2Qet66eY59mU32IHvxvw0eQzWKzAtaVgs1QLpiNQU
im/kK9U+ePnwo3TDzmhFj8Bwiy5rJi9RSZAW0DAcFMEkagFHF06xnseNI7PhSa7r
jPVb0UZhU2Bv1hMl2ZdcHAerzPYR8gdC5DrDRXrAeT1Ng15F9cKijgUtWloZcnLK
Q22bJUqL/u7h0SctoGUIwnfyFdAUY0X3ek6Qeck3PBh5W/tb0Ir5BS/snmRhavj3
22y9OnzwhC4iSjZTpSr9EEph8Hs6NKdziXAXCce0Jxva15cgZeKfL0cRHX9WxbHN
5/ykoMUoFZbGiK9hfoI+iyq+lDMHrD/S7+B01aOk6/KYeMPtf+VUUE9BuKB/GsSJ
IhL77jwuSg5lBRo/EQlKtt+hwgkaI6lXUw+/50Cq8qAwonXDRipGtZI4CC/Q7hXo
idoOeSt9ifkYPkISp8Ohxohw3TWePTUcE0EZEbtpmxvt2AYIfi2T1XoAKM89RSKq
d3YsOPmDzUFPfRmK306nUBRw+PZ1rDycvqdWWEYZHk4p5WE29tblvoJyz6vlE/F7
7XdQwwKAAA55eeTT5pZX16kP/z1M+KD3TL0uekaQovlUivLgspYG63Bf8rWfB6fs
szzGRf8iaAJfTM8cKet4xou4XaEIPg8Fsf13paRGpR2y6TqvFUo0Ym7HczEGLkWU
a11Ig9ZECB9HVsPOJTK8UPCNW4HUOcMi0cCSwGCNplb3uRy5r1U/DrClouBKtXUS
UX2MoPnoABnuWparCiM9YHQHYWBMPMoXbwfoOCJxt66mSH7sWxF+WCRK6uIioTWE
NldUXndG9K1YCzXn74JHwcciupLjqGGoivxa43NGv394zMap7fnwVeT8wSVEG8Br
RJYE0mmu2wgEsQo60xSrzt/bewkNqCfaosSL0Q0fCLVFvxU43C6E/XM/B7mNDjFo
IwSFJ9lV4w5Bcrd2xMLxw+BFrnAQOX7EOedZedd1FVsj5Xw5mMlEqsXOBYH/SksO
iQd5cOMiNC2mU7mc+5FBJw5cEJAlEtAde6QaQt2tq2BBcvmqx+Yag5eT2jkEWJO3
0pAHk33mdHdwMgCul2ixHn+V+21r0pRiJ9K7wRxZXP+4/Bo7kmeAYyPGYKxiosac
loVxWbPfFv4VvdEylg9pEW7kZmka1dtFuNPfyEXhJBPVerjF1lwCFI49mSPDlt+X
aNG5C3kEplaC1QkQVArzL9KB1F/6+i9iIB12mCyTl2M+NVUTj4wcFlfuUhCefZVA
Lj9nvl35S2E7cR0RCwqGlAyZiFl2Q4UjAoKMren9R+V6VBce2G1XmcEUJLXdNO4T
+r610/Az8U928OrZi5Dm3Te6oZ0wvq5XzW747OuNgzBTFlI8+vqaHiXCHZHTLjbw
il4ttxOon2NhoACNBlc1X6BVTjyLIucQyWjMYkYIF0iUXMQ1LS6AlCmxQW3hPQtq
yp6ljyWEouiKeQNziFNQ5FfAh84DCd72PFloll1FUQiwEOaW8R41+EDUMb4iiwJp
udSXRjoqIVozK305qg6kmbj1qF1+yb8CLHklm6n0ej/ukuNH9ZynJxlXwo8/jHx9
Ymrln2z26OxMwysd28hbPnye7lDgY5XosUCUaP58ywnQoJ9e7eURBJANQct738VV
0ux+iPff0uvkLZdA47LHg3zxfEEBt/7ZE5U2ZgPd8IWXa72JrkdBd9sSjLYKMuN8
b+wct2ds3srJ4DumCvFAWI6kyWl07Z36+KfAzcSpjzo8lAaKIu9opUJqleDBUsVs
g6wTEFzpuYYHjwai/V9yB8q3DZ0boc97XD4ix71oCNrOXdFUc66hG5LxOTOMje7d
RjqnMzxb08IE6cWLGNvjwYmU1kwyGC1/5L81rYHeiB77bOuBhhMOUHZ9kb5LEPPP
y53cTC9Cqw0A+p6sGYh59/jn2Lrk1lWOaZoF3qp7odQWGqChokTEQKJHBmCo7YfC
2Os7rKuaXKQSx5TW/Bj9OIBZPe9pqrZLHyn99vdcsyH5Im8pzUWRri/psn6R/RIv
ZtSTUF36fcWbM1J6fsax4jLM4TwILB+tqb3LLIRP3tRqlN/xUuTs9yBgbFLuu1By
BWknxV07YGzIGd0ik+cHO/xUnbr2Dl7Ko8SS6swqWn7xdjQqY1xUrbIVaPDooq2B
CCuIUHzA/NkFXxvafnvxAUSGsqnYJ1mOWV6tN5QRWS33cNcrhgZUGAI4ub2LixSs
Tunf676mMKlsXaOU/l9Yo9gu1HVdj6RNZ6p3cfmVL3+mTu9D/wevxNrkQo4SFi6g
4YAbH5aqlmv/nAmufLAbHj5MvjuvNMHfAvYy55QPFe+v3ffDABNhQ5gxmodkotiD
RC63mh4JF1IJiR/ufIFhPenzdVxwskjt4L0U+TMG5BBUQrQuIG6NYrCwKbe6shxi
0M11kvDI2v0X/bTpCD/mvMUMaBSnwxgewR3VyI3NisHKxKQGXRrrvgH6TOzssb3K
OZl5e/WjC67ypKowKcq9B19exelQXV1vxnLyqDH7zBilLbup/k7+XaMlN5aDOfkK
yIEK8u7jrGo+ZQcDp4A9gTGifRCqGxTf8Q0uL4eCCyMu5/bX2myTPtTl3Q3cD8+A
jtRBjn5PkSZMI/NNaA56MX3l+k3VQs1vAQgE4xUPn/s7Yv8Jc2+vzVZNPmOagLHy
lUk7f+3737WcyvoHfREqjTkXYs3g9Pdx3WDCos7IzVspX/MUPXQbRvcgxvWi9n5n
dakcztwOEBVp2/u/NOnCQTBSIervNE2L9M8ICup24QtYPF47omnrAkQN910jJNbC
1ibIian/NrGP6sLuFL9oIz3PGuUxn1XJKeuWx3jA1xUbPqKNbsSEfKvRYg8lzDKG
UlcTCD2po1KE1LNGcttLrIOZ2ShtAEZPlfkc5vbaVfL/yX93pHYGALGh5SJoQohS
T/P7on3ZPVLUPvLfG/5hwmb+d9yrD7hGlbD/HIOx2M0K8/h3LOBa6CT2Rg57ndvT
uEJFxdMXjf4dZQOR/l81Qlt+6rKkqN+/1R4QUL6zJr+QeEJYdPQfkH+Lpj0JkRbv
TT8umHefJEUpv9dWmBN+vBAe5/zggqzcD4L6WhrxUo3gmTu1jQw4E+LbUc3EY5QZ
9gG/HejDmBvBruFuymiLsFYwYdWYnJYnqb7Y9YsBWRommmjfjL7mQH21T29PB43A
TBXA1zZu5tGaaWzSxFe11Ic1emx/dY7o1dTshmR/iaQ2UWH7/RuORivCOywqx19y
qlI7wApC7yf6gJl+bueCrko3DhXnP0aoxUzvGknbHiKqeG9r5B7UQNJLU45DPmhE
hoVsYKtcoU0GF/PSkgMvPy+lSuG6ST30laVfqYP2u1kn/D0gEweuUJf11rbYpFS/
Eaia7MkKWgRHdndK2OU6WyiwmINOvYTAxrNbggPgCHglwEtkiG9Wc1xcSJ1K6djp
bqd7mODlkJGyjPm6oOjNabC+iRJRPxgXjTaDNMCRvn2AjZVWZvyboJSYgLIB0PqM
QmgHksLQ+hawEcy0bBznTWnZiBKxmr1nuQgbUwuXAKfRcb1dX9+O3hB0v4xx9wcF
2pQpzq6a7DyXnQPlj7n4fLMCnm4LCAYWUuYYvZ9xNp9poxMwlpr3xwbpHoBRERb2
+LNq3P+Gtk5nZxQBK/qonm6evtqwY5UrOS8kAiENeQNYnJyc956U7GOyK/uUx7nc
b1NCxommlgxioydy/1IFNE8jes6JYUaVDRBXVu/JxqJ1g47iMu7wkHmt3tCZ9zin
9o+lQqTe2tTCroX1yDb8MLg9be3aghIhKPqr3MZ/6UnaLp8ArIkW2Z3fvnAX0EXt
SBwZXm92RXJK9Vo20Y4f9kna6e+9sW/XmhmS9bePl+khmDTeRrdn3LWqDGM/dbgQ
D53eMqVIvpfNyDnBwGdONrNTosaW9Y7DQvCvVWzIwqWbaWgj5MYeQdCHBXhHfr31
fgd7lzWquuTZy/Qi/tgivVmgYnbplA1TgX8FAHzuhj5Yxs4cRSzdTjIKnrqL7DTg
Sgg6pHcVM8JkyhQU1Qk2UQ78Yd9zmUt4Hs2UZAEBio1Fu6OH1mfMXiBSLO9oDP63
ObcHT0/iajBBqfr06DsJ/SuRsWN26znQIr6A12fAU5SFzku4yXh2v6hRNUFyzcLO
7PkUqbF8fuectnKY6jx7OQ9uSZIfEFMjMvr8EXlBkoJE93g28+7TlwEkjsRRcw5g
RUOVVLmbPEwWTK6FMXdXjRN2BUcKiN9jWC3Onj7UJq1EHmN8RXSXbhmVv+Cv/F3J
dhs6T8R31qIhV1cuRMvmYTifCV2uum0EFZWLS+P5kmyi3eQuglzx2hnkL+kFyZBM
/o+1ImHY/QPwgNHlGf7NvYF1zjwCGxX6lajPYmTpCwwPIX5N269jCqjYW/hM615q
NfC0VmqYM7IJjJVoEr7+EQlfzr9ZBuFUCeSOxVrTJwu+t9ifpK+PFD3OneVOKPBL
THGmI9QR9capXlEboTP3bS3oefB6OAex96gHXJF9lZljCNZXz19LlYRMtr79EXON
9ONKz6dA/YckEdJ7a6j2RtS24FfPka7s4Ssoi867j6dIPCWrfhjOQBDIGw4uGvnI
9ETyGhRn5+CY1HQFUs6ywnU98yWFjOTOKbOt5kE64ihJzEbJmtrjChe7I7KvPkd9
Dqu6gsRtZP/5E+6KxRwghvzFNxfW4h0bBoPi7Gl2svDEvu6aEhBh0aqUH/iUjO1G
U53qOR76qdSZMpWz9z59CR9ZEuHDpW4yMIu9E7lOtM+gJew0rqaTuRhK+j8i8yim
eLftGXYUD+kbaZiOUyDztPIbAFMTLCW2dQi5T/lR1DeneV/fk6wRLT2hQY3rGoAi
PRlvP9V6WyHzQqK1PZJZ+LNXl73eUsfsrLw3HDnzjhD5CR2h/XnZnsoyblI+Qls6
WN/tF7apwH4x10sy/nXKr0FOJEg1jsDmGwNO1LAcMFzklmO5u7mvOfCIWrdNNlxU
KODG21ZUyz34GGwxxhdSK4kCd49TGlwdvQ8mUTY7tVOxJrWC0fcFR1JtLtHT/P6j
H/sCKfAOe7wTfMPyr3FTx1WmMeNG910IEjSJimp9lZVbwWBPLSpzA0xOzEWDPyve
eNmbDlmPvh0f+FfSyaHuH5vaWEUkkUvwT/z02dymqZnkeJO3EacQNx7szQ7h7daQ
K658K1VT4O9urcfbRHeWZBJhUTIv2oxIQubn3ape8isSAtHZywQs91kpjhazn4pD
Wo8vGfh6xt4VDne6le5uxfFnAiTZEBbKQFn7VwDF3ugX5vC7s1JTlE2dsdUP+dpJ
e9MZH5gDTlidWOFRSjxclpKqH7y1RmQmh2op/OVhLpgOvsyOm7r+RBI08UAZR2d5
uwKrAnYAemMH2TXBpVgSIk1PCd5nnx0XVC1M5l4Rgb53dChs7TAclQePA4eaxW55
iwYDXe78Ab0t/OE1L3QEPxGNkOEaQOF38k7f5JmDGba/kjfO5Eb4hVtcsyct1YUC
S0nLn0pTNEZkAs+7KRXfkEfVl4hZyoyP4xCdvCa6igvTItoDrHddazyD2+DsdI1a
f9cHcNBc3ho5SvsihgQa7eXNxShIQnfyodOTu8gpE5e08m3ASzGimHRtF8OG0InY
Vw4tc6fsaROiquUqyXVaKCYHXJMxf+lLF05unBkQZH2yhkqi0xVmpH93dFvfiNlZ
RC4xSmjx2DBEBAlOHHjLK0SS838jILWVSCSEoT8CryNApgVYDJzxgk+rBaq35Ev+
lw6kSY7qaUQHtLjc36XsiBY/wSesb2/rEk0Jv++edcNdttle4x12oz7LrTvSFtpE
fvdzMv/gTL2sNXpT7Y6pMtCq5Vb1Oscbr2DU/7TDHVS7P7QVEUiOdVTNxFmV+wVX
gOTI9ofIe1uth7oubVGMCmRjcNJY2uAmc+qfiXK7Mn1mUbnJSzhFZDAamRG7kv4a
aq9Kc77JwlfGqso8nMIF4CjZ0ms6O3i7nlcPKXTOYYaJn7sac6tcqzENhi/GbHjp
eLe46P+/BMvFiA3rZybw5xBIq9rQdnaGzosqxzHA+edZc3RP8OVMuvWswr9mRIaF
KPXRDRZ98nx4kvP0uDjP8lvyutC5wtVvPjfBgPlgv33fX9PbiBvb3VcuYvHabUFg
fM5HJigaDiUelnXsSTJT23kWCQR0e83doMI0AvsrTKcxOl3pt4lRsBbLxWzM30D8
CVEoVa5aqa6klLctP+8w56fhrszUpqXRf7b8ARPeNUtAUBu5sfk7hstcJNH4c5m6
OdCCM3U4X708bldDcSl8C/UyvUot1rT36fkRsWPxOF93SVYpTZkhHfWbECLr5LmS
PhJ3ATZbR3VXgCtdOqbyarDPxa552B4tbS5Y0YSOEsnBC+B0iQs2fhxPUUojEZl1
Pa/sswCEW63PpAoheb7gLIwz0s2B09NY38T2v5EUMgze5vdRZx/Sws9lQexoKzAj
bbuhkV50V90hDxorxALuzzyNZu0XasSDgUtywWaMA4y92mSO6Kd7T97gbOwL4YcU
6QH8OkoVqKcqZohy+27gvjPxN+suUa+Xase028yCKfvImhjj+zh2J8kY1Nv+LbX5
U6jSqmoGqjnwDMsg07MPt7GwABXtE/QB7IbBJzuDgdpVpuzCms8t6lDIVveh1/i3
1X6NjUKs+nbk34hshtnVPy7F0qOxn9zNZ84bxpTgjf6MCMxdFphf8A9KN6P6yHa6
rTwAk+Eftw75Ats4Ww9+Wa8mH/fArMMFx9cM+eVwPqvQrV01eELuFHkUjQeenK8A
sTrJvQOnUBB/HyLMweqayPglUIksjPc46KPa5wOkdqx2X1DjqsZi4eFFCNJW4Btx
LYX9zrrAqgexlCkT3aBht2Ws2pklWr8tooh8pDwQ1xKiimimNHhYER7+TQaIBcIC
/2zEhAoe5Bd3yWG0ZKitXUhJToRwPzE0BmThVZcyU5YK7msfeZ2GJWfW/QWRIUK5
RDAPDfgKYBJBY4z5mF0bRKtcezZYb5kLRjsedz4FMBcE16eyTXZiXk7xbTXHecck
T4j7gUDTjsQ04Qhf1VZUcAfXG2EENUSYBFMamFV6tBIaJzH7q9EEXF+PxNEoi4yk
5EfgxppVnByupeBeSLTpKGQEf1IebJ65Sq/lSRXURH+JhX6CIdy9Kqs97xgPQy94
xgf0jDIxGQPGU+qYJ5tF5V8Jvb0miBYaZX0rjsRH7VdpBvrERbP3gWlsGFJGyXJB
S2yap7mY9xYCMmRwiUKO3hxuayhr4oZtNVc0Qnr382FIxgxtxLkWU64VyPorC4YR
dmGkg+3t7rMKyb5IA22wQvSvvlWNUuNF9x06KfmUHFhl+8cXFVSjLTXGbgSfm0Q5
thduz6cSs/hIQSfwSgXK7bWD0DjYRRgrm783aTuc/yA+Rtx8uW1l5VEb6XalM/F6
GJAcPEaQAAZ8AJPyKXKl2pZWZ6KDBRpYju6H6RA0UNG2NqMuQIASG4af0I0fTCmv
iaXu2jqLh7k7wPQ3oNVrGDmhuLDBYK5Fxtme1ry01i2FjCcVuh2bY1FDl+PoPhu9
zMwNWyPgGotcZGdzSVBHvv9kahfnXxHKeg/TtFhdjJr6KnRty3b37gUDs9kasD9/
loXx3gYMkVWwlGZOf9AZSCPG/PjWtXcbE+OydDAzuKKttilWf/hAX7KzWbJY2hJI
rI+hKsJDkLiFVC6LOaqAS3fgtIZN87F0fCqd2vDjbLxRSXCUzrTqm/5Fw4MoNZZA
yD5H9AmovimSxhVKGLujIFiy0EwfN20jRwSHD6PzhjNXukkpKP47Yp7G7lqa3yif
V2HUKAfSqjTH5NceFk6jIKaWtu0h1feX7ztCSaQPoMxZRzQRcb3d2u98VLwWbWow
hMcaf8lPfX2DDeyI1wE4BvhpeBc/2d1KT0cRPL2dZ8YdPFEF1SszkvZWHw8xK47q
8QhOz6mdwaURvvXokhGupT9YsP0C9MFufBz6CV1B4oztqhNyI/bzEob/mEix2Dzr
Rsma0sh9cW0kyDuidM+HPwFbLmy+VW9MGAqkVx9R0z0FEfNqMkTJJINkTqhOdpZ8
lpJq6oJt+1AGZ5P3mlkJAA10g7KT/GxvWKX1OMC0jnxNZpz//4EAtOdfOgI8fY7S
38nKCYu19OUYpkgy67lUhL4Pm2+0w24TjsORWcKvNGTXJx+F3MTtKBdN0syatL8K
VBxBtkoYLy6/PrAXvIWx6y4rslH22hnpxw2WVeG/9mvB3GdqiHN3ROCM/trb2eF9
muC4g7DNKIPWP2Q6gkFfbjJY5tWfLmeD5xNVTRrldOXpxYTHtJoWIcs8pEi0vQny
xT5UXOt8HoMtU1fCQLe0ZALX2wx9I+1ffz4HC5/EGSSUhLl+e3ONYlJ6ARscipes
juSFktM61qgUlDVzxvbzY9K9ywi8X28riLWYGpZzMAUCaCISxQ/MFRP4Q0ft8LMo
QkD5lnUPvVsRZbF0Y+3I8MTS34qnrHs8de/FNzb3qi+vhrJC8tBp0CEsaoOXeh04
eslLBuh201ytam7RTEWoCNHt9ebq2CK0x9GCpGAQRzMtk6/CLCYXW3LY7ub2a4hk
yzLvzxPh3fd4YZTUZk84qNPcFkKCMqt7bC82lnXU/FTm26spibgyjZZByXrQ2LMK
HYStbAgZiUSZv1Q1cFUPaQ==
//pragma protect end_data_block
//pragma protect digest_block
4/1Kw/eDP15t8otTAFRf3ZSdTGA=
//pragma protect end_digest_block
//pragma protect end_protected

`endif // GUARD_SVT_APB_CHECKER_SV
