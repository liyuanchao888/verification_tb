
`ifndef GUARD_SVT_AHB_MASTER_MONITOR_DEF_COV_DATA_CALLBACK_SV
`define GUARD_SVT_AHB_MASTER_MONITOR_DEF_COV_DATA_CALLBACK_SV

`include "svt_ahb_defines.svi"

// =============================================================================
/**
 * The coverage data callback class defines default data and event information
 * that are used to implement the coverage groups. The coverage data callback
 * class is extended from callback class #svt_ahb_master_monitor_callback. This
 * class itself does not contain any cover groups.  The constructor of this
 * class gets #svt_ahb_master_configuration handle as an argument, which is used
 * for shaping the coverage.
 */
class svt_ahb_master_monitor_def_cov_data_callback extends svt_ahb_master_monitor_callback;

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** Configuration object for shaping the coverage. */
  svt_ahb_master_configuration cfg;

  /** Virtual interface to use */
  typedef virtual svt_ahb_master_if.svt_ahb_monitor_modport AHB_MASTER_IF_MP;
  protected AHB_MASTER_IF_MP ahb_monitor_mp;

  /** Event used to trigger the covergroups for sampling. */
  event cov_sample_event;

  /** Event used to trigger trans_cross_ahb_hburst_hresp covergroup. */
  event cov_sample_response_event;

  /** Event used to trigger trans_ahb_idle_to_nseq_hready_low covergroup. */
  event cov_htrans_idle_to_nseq_hready_low;
  
  /** Event used to trigger trans_cross_ahb_num_busy_cycles covergroup. */
  event cov_num_busy_cycles_sample_event;
  
  /** Event used to trigger trans_cross_ahb_num_wait_cycles covergroup. */
  event cov_num_wait_cycles_sample_event;

  /** Event used to trigger trans_ahb_htrans_transition_write_xact covergroup. */
  event cov_htrans_transition_write_xact_sample_event;

  /** Event used to trigger trans_ahb_htrans_transition_write_xact_hready covergroup. */
  event cov_htrans_transition_write_xact_hready_sample_event;

  /** Event used to trigger trans_ahb_htrans_transition_read_xact covergroup. */
  event cov_htrans_transition_read_xact_sample_event;

  /** Event used to trigger trans_ahb_htrans_transition_read_xact_hready covergroup. */
  event cov_htrans_transition_read_xact_hready_sample_event;

  /** Event used to trigger trans_ahb_hburst_transition covergroup. */
  event cov_hburst_transition_sample_event;

  /** Event used to trigger trans_cross_ahb_htrans_xact covergroup. */
  event cov_cross_htrans_xact_sample_event;
  
  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Coverpoint variable used to hold the received transaction through observed_port_cov callback method. */
  protected svt_ahb_master_transaction cov_xact;

  /** Coverpoint variable used to hold response per beat of a transaction. */
  protected svt_ahb_transaction::response_type_enum cov_response_type;

  /** Coverpoint variable used to hold number of busy cycles per beat of
   * a transaction. */
  protected int cov_num_busy_cycles_per_beat;
  
  /** Coverpoint variable used to hold number of wait cycles per beat of
   * a transaction. */
  protected int cov_num_wait_cycles_per_beat;

  /** Temporary variable used to hold address pertaining to last beat of a transaction */
  protected bit[1023:0]  addr_last;

  /** Coverpoint variable used to hold htrans type of a write transaction.  */
  protected logic [2:0] cov_htrans_transition_write_xact = 3'bxxx;

  /** Coverpoint variable used to hold htrans type of a write transaction when hready is high.  */
  protected logic [2:0] cov_htrans_transition_write_xact_hready = 3'bxxx;

  /** Coverpoint variable used to hold htrans type of a read transaction.  */
  protected logic [2:0] cov_htrans_transition_read_xact = 3'bxxx;
  
  /** Coverpoint variable used to hold htrans type of a read transaction when hready is high.  */
  protected logic [2:0] cov_htrans_transition_read_xact_hready = 3'bxxx;

  /** Coverpoint variable used to hold burst type of a transaction.  */
  protected logic [3:0] cov_hburst_transition_type = 4'bxxxx;

  /** Coverpoint variable used to hold trans_type per beat of a transaction. */
  protected svt_ahb_transaction::trans_type_enum cov_htrans_type;
  
  /** Coverpoint variable used to hold trans_type. */ 
  protected svt_ahb_transaction::trans_type_enum cov_htrans_transistion;

`ifdef SVT_VMM_TECHNOLOGY
  /** vmm_log instance */
  vmm_log log;
`endif
  
  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  //----------------------------------------------------------------------------
`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTUCTOR: Create a new svt_ahb_master_monitor_def_cov_data_callback instance.
   *
   * @param cfg A refernce to the AHB Master Configuration instance.
   * @param log A referece to vmm_log.
   */
  extern function new(svt_ahb_master_configuration cfg, vmm_log log = null);
`else
  /**
   * CONSTUCTOR: Create a new svt_ahb_master_monitor_def_cov_data_callback instance.
   *
   * @param cfg A refernce to the AHB Master Configuration instance.
   */
  extern function new(svt_ahb_master_configuration cfg = null, string name = "svt_ahb_master_monitor_def_cov_data_callback");
`endif

  //----------------------------------------------------------------------------
  /**
   * Callback issued when a Port Activity Transaction is ready at the monitor.
   * The coverage needs to extend this method as we want to get the details of
   * the transaction, at the end of the transaction.
   *
   * @param monitor A reference to the AHB Monitor instance that
   * issued this callback.
   *
   * @param xact A reference to the svt_ahb_master_transaction.
   */
  //----------------------------------------------------------------------------  
  extern virtual function void observed_port_cov(svt_ahb_master_monitor monitor, svt_ahb_master_transaction xact);

  //----------------------------------------------------------------------------
  /**
   * Called when each beat data is accepted by the slave.  
   * 
   * @param monitor A reference to the svt_ahb_master_monitor component that is 
   * issuing this callback.  The user's callback implementation can use this to
   * access the public data and/or methods of the component.
   *
   * @param xact A reference to the transaction descriptor object of interest.
   */
  //----------------------------------------------------------------------------  
  extern virtual function void beat_ended(svt_ahb_master_monitor monitor, svt_ahb_master_transaction xact);

  //----------------------------------------------------------------------------
  /**
   * Called when htrans changes during hready being low.
   *
   * @param monitor A reference to the svt_ahb_master_monitor component that is 
   * issuing this callback.  The user's callback implementation can use this to
   * access the public data and/or methods of the component.
   *
   * @param xact A reference to the transaction descriptor object of interest.
   */
  extern virtual function void htrans_changed_with_hready_low(svt_ahb_master_monitor monitor, svt_ahb_master_transaction xact);


  //----------------------------------------------------------------------------
  /**
   * Called when each beat data is sent by the master.  
   * 
   * @param monitor A reference to the svt_ahb_master_monitor component that is 
   * issuing this callback.  The user's callback implementation can use this to
   * access the public data and/or methods of the component.
   *
   * @param xact A reference to the transaction descriptor object of interest.
   */
  //----------------------------------------------------------------------------  
  extern virtual function void beat_started(svt_ahb_master_monitor monitor, svt_ahb_master_transaction xact);

  
  //----------------------------------------------------------------------------
  /**
   * Called when a transaction is ended.  
   * 
   * @param monitor A reference to the svt_ahb_master_monitor component that is 
   * issuing this callback.  The user's callback implementation can use this to
   * access the public data and/or methods of the component.
   *
   * @param xact A reference to the transaction descriptor object of interest.
   */
  //----------------------------------------------------------------------------  
  extern virtual function void transaction_ended(svt_ahb_master_monitor monitor, svt_ahb_master_transaction xact);

endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
wGWpvu+30me1hXbX2DpbIGsiAVB/DN2HH9bqWfWRCljVzhyaKxB3G07y9dtqKV94
HgvE4NuKMXbw7rZTZEbeOr8YNhGmj4CZQT4wXGLv5uqOak6MLQHDI2S9wgUiNxlg
Q17Gc8MCNwUlD9XYXkwqzxxw07zVTvPj2n9sJsmjvve44Azf4jKjVg==
//pragma protect end_key_block
//pragma protect digest_block
FrXOwvFrWpk+X1JAzpmqq+4/4w8=
//pragma protect end_digest_block
//pragma protect data_block
q5DsinwGngGFNtrPPAbqlPgndFUagMh35+qBbn26C+H9+stDabu2HUefyf0Yria7
CCjM2GnYWoQhiNCYOG9cbOa5Jaq18QQCM0ldRCNBcgTz+mGYpHZRzToYgDvLi78n
Ty35H1iaZpP7bDkntqzVGvGzYW6+ZH50/KWUPbB3TvRuDBnl0wIHByjQHhSTXxZj
//FlNLVE7o2zQcLJqj9057aeJnNfw+8UcLYnyJxAzlIskhidMI6/Yaxw2VZSAhKE
HmApa8HZ96ouW1S+HXVOADCNvcXb4NYCYBg+CVm9Rigoi9LrGoRqNC26hvlDB/XO
D5jf0l92WANkUxNo6CqAAG+2uhswrCsXdhP4ATA9PTPq72kFAGQ/WFQMnCvGRgun
mtPOGvoATHuVP5QXa22B40qX5QKFEMWtLmPjpnYUooWium4qbfD41DUpKz6Kzldg
NWTFOcTmjx+ya7uZXjRduM7H/pbnsfWBtKhYUvInvkH46lMVTKM9A4Y3Wugfi4Z9
d4BcyqgMEK7kLxoMVTUVi0mivRD5TrFYEKgyBKK3IC6i46ydHgWfNTUw9oTeIMpV
Lk0Dpt7vY3VGh8PmESBhRkmHDMromh56Utmtylje6eIJWdDvazTG3uw6j3i4FAKg
MhXyGU4YZxTXbyEVQhGqShw2RZM4IHx0oexgtCx8SnVGCKA6CpmqksKhRP2ptwuV
pHm+LyrQJqjU7dADaIxZrBWMEGXIrn+ZEXfH4jcwold6zEHfgGBP4ao+q3C4dhGm
TT34heyt9KsGxuO7y0tO1AS8GDhvKDBOtLtG4B57AapYDgfEetHk5GObTSBPWA8k
QBkr8T9CwRkllnik+cg41p4ptGqXboj6GVpnnUVCPiLs3Gwil5T2z7rC2dcTNgPU
ZwWoU2IshBeup6PfUYnCL+GRY7rhGhKIbinTpUtMI0NICURxq8Ib9+J9lgcDUxCv
5y6cvtRApuRcJxzbz/sqiuENiSy5dzx721Z9iqekVt9dE8pwDSAwBG9W27LWxDuX
yer7Jl0TfemI2jMZENadWNrT6X/Mgn0ym70MBrfynwQR7FF95qZ7COa6q00ll8mW
5aqjDhCGzPEB8rHUNVbODhMb9ZbpbydD1pSQEymGR+H7hhS2plrvbgIoj0imX2Lu
gg3Vy7nOGoz3uCzMN+oAZ3YqyaisOSDO7sxv+HewemVOZQdo50W0v9X1X7Hg4xhf
ANixpt3HdGsRUNbkh1Qwozta/QWV5FO5s+5Dc65mQy2z4njfDmTUvQ8BA1Z53X1V
V4HgPDgKWQWdhd7sOHijxAJeMsXflnjt3mtJt5NZ+ZS/aabXfCAM37vOIwotZpfp
hICNVCdBqRpKh81nFIsRzkKacDbMc5jFNfoB+vYbDsHmya2s2KW2GqZNmxsc8/4d
wzYpfFAgv7HDGwz6Cu24vHTgS+S/2rUjuBQjWBhb9n7VeGoAmJCs0I8y8+QyHSpd
XnEjji2qs9ejDvjLm9KSTSBwAmS3VP9pab2uo0U4jT3wKpA89GfisoLfAiPrmBtW
sdwQ6f2LkQskmu/Dl9rkCZdY4Z4acpWMBfNigDuwRuumXrXk3gv5v/dpLeAY0Zrg
5NtnEQTsxTC0LbrY/iLA6ZHurjVPbga6yYUnJ6PGfbiv6Ns9JsW1qFzB1ABGhKOV
nJviA8o9yxoRmCsrxQAKTN76l91LwHGChjOXhN8EF8i+XTDl2xhpS+74wpjQUrER
fI9KeXf0dpSwPHnnP6b+tUpgvhouaC2v+23JzRfpRNo/Z4kAcmPGN3NVuL9innY0
+Ol1yh+u/c6Fvpm+LHJwegysio22dB01UDe2S12mHAAcYEV4E1ozrTD8sNbXGuD8
hQRUGyHWL5JA2EWQ4hP0pVyE05jVNAwpQC63ZMcRM9nM2BUOrkibPea36Swr0cGv
Hqo24Ljv+KJw2wmXYJvUdF0OsCKczFeKF6AEAlW+vsNmccbu86MRpzB9qC+tD5vb
Ol7YjZoLukEHqGBmRUMFU69510CwviqdZUgWxVXepdzqABCTfnOSbRSI2S16hgC3
T365Ctyp+oUzKQBMKM9C+6ns+YY32fXlb1AVFBrfEM1t2rIC+mi8EeGnVVkQw/iv
4f1SjwwBm0CZi6zFD/mCLVuh1ZqrXVLswmBO50jcquO2vQxcikPEDgtnUli1tvAR
T+BFlyyVirylHiCjuFBMjlSqNpo6gOWtbki7M5JZN8RBe1NxVaniqINuXUB7Z/jD
54alhJu8HfbQuq3iDPDp78FUM0Tw5LR5ka7obqjuvrrQBl+YDbVt2YYYrYioXHpz
XsFjX5cpWJc/cuaovg3QsKnKd/xXCPIUepEOMElygy05gqKE85lDEiI6PZo1aJn3
JXnJvbvGaYxjnfZMjyzPyJ/B8RTjeYr/i1c3s0mvNDL+Ldf16XwYHkhabBzQQnPV
ZGjTuQ8KMB1DGQP8GQ9DT7qACC1ot6h8N1IqxHcfvzVPcTRZQ7JR6bC6mZSq74j+
bHceM2Kl3BnSGJe5RFem9jV2HEXeai0Gbz+fa4ZLEmXHF2H3EUU5c4oEgxVmX9iZ
SHJ5TJMpEtV6ae+7yEOkOqdJfqLibHvqljNzK6sluvH1H9bPiJe6thN8AP+Z5Jcw
B3Npox0kthPatBMUPxX6pDDjYb+AWPh8gc3dakca5FOZj3I70BMHzR5FQ1f8/7f1
OkhX56LQcBmBXZHKAWRnOXDBv+GW8Qq8XLf/EOICqUn1LXDLoVLjGjaBhv/KRYsG
JATJtcRb+0n12j2lMvH0VsToshOjSk2nIi0RALnwHAQbRfLvi/KOG2Lr9bt8wmz0
j8uk58K7W958stO4xGgNb3ND/jjVFyhKxa0caM710XDI33jrdXctnLwmHAYb/80w
hETYZuabIDD3z43QBz9Ylp+uJXYKcaZ2aKoyj55FhxE3WPkfyZEA0vYOxqG9OqSb
Yd2YuIH01twV2jgNzXf6t88Sx+j0e8A40aK6/idSVAX2vEvG2kE2fK+JvpuaTKA6
Zv4q2x/A1QMNrY6DM52jYTjbJIzg3g7uhX0kuMuSVq/9O0TdZ/+hMj4xYU9AIsmD
n7F94EzTBa3gjsnDCMEXRl2fAZMDZhezTYVkGZX6Ly+sSaywC2INoZqHvaKI26Tr
Na5qlmVZq2u9CWF5iyLwLlycxPWXNnKIdgFeGbFXZMVC6eDJHjc/+lwSAEasiZVc
dvKqoqswkl61n58cLQORVDedAYwiC4oR1vRluIWWyIFLNA658IgyVXXEiw0fIDAv
bEmnpWqKqA4nxj1Lhl67n/NMw5dUwP/dR2B5P6l45rhM+pv70k0d5dOCpOAyVuAV
c+0c4kTCOPrTPRpUKNhhwVOHyxWyDTHJ/oDVGV99fp1AvOLp30FujBpZoS0BogQU
w8JCjR8x4945vafgTEFUmfQzuVSUW/BZKl6cPr+Aj7ptin32V8lUY1R6OR3OEfl4
lqwPCVf0MQsNw7pW/BBJZKdzjIbOMrhcLSPIAVEJmJpQewJNt6hvlCOw+fDIW8ev
jEp+f0CWRNBq2c7KdCdbB5UIMO1QSjL7HKn18TmFZXguiqL1n7ea5ZLNyNBO1eE8
i2bw39rQpU8b9xI+rwPRlQGljx8Mx//iVotpeFH+2L+dg0KY7ZM/sj+RTJi7Rgyt
Wxvp7L0X1gaV2s3WLOF2QUMaFPegPI8Q/qRWhwMnXPdvfMAoTjc40tLZElyIN6Og
tQ2iAMMm5xt+zVCrBpnRidB3BKprQ8I8plTJ0FRSBsrwtTKBO1YKrTwYtwAD50OJ
Jq5fZ+zow3lVGDudf0JfIZoJ09dISX9LkUu0EcqYVjwIlhvAICFXoapNi2WeR8KI
DhWPuJ+DmKI/N7jswY4vmL9bKQX+a57anuxqjh00xz+eSPSnhIgv8FBdXxc8y8lD
j5r5YXhzdDuxJJlnL56gcLdLrx6c6qWxZlUr73ljTPR/DZqn06ULBCLYA1RxA84Q
As+9HyLpjLtz2PKnOZSA9m3ax3qJM5XH5ZIfFsoJ2WvlkCd/76Z9GXt9xcHl8sOT
+BJnxqs5l4xh6WEevIK8UAuncyWcE7q2p8DU1fwyyvz1htBm23CBo30ZN5GFBuwM
LL8QtVaK9MDRhUcGRlgpzJMRgdnXU1+z7CAwqTHDzOpSHJHmJReeNypBMmWnhWUI
WGMsKFLlAmwtfT3xW7shexbjewgxF0uCqdHMS/TKgD5kOqJBEf0yc43uywgCg1yq
ExcHkHI1Zy7u1uPDVX7enoP3F0OMcp9JrH/seDNRq6WV/HdQduzD1qj8FDllPVW4
CUW6klEa7H6jpZJXwYbwpMUm0PqFNlAzHt8pHF7O3xg55D2oa3PZGFuEpgd0aX1d
+V36GJA/Z1zAhvngvaJyhc8+5vYXgq1Lh8WID1S5NdTMIwWs36Nq+uKhPK3sLjHJ
ZHbGa/rgO5dZFZO8hqqqqaeYwBIifTdDkbGuTZnq3bVtF0J/Bwp8sV1oZQTO6nL9
/VNgswV1tA63UPOjk2bNq8aOoYBzkTMLVFg9cItkDHk88usJ/5ZpkQZy/VbQ57kw
YND5e+QhI5dIKb6YKadWV1BFrEN3mk2H7f2zRDYyIihrkDmtpiWnrIR1Qgyp5XsW
mSukjMs3WaawIsw2icC+kblga5RElGbw6GUjOy+u5NZnnsIMXAhraguK4DPVSp57
VyxX7p+Nno9FM2ktZSboWzANwdcFFy9RZRKKxlRcYlpX8h6+BTtYG9d8q0gSKJtu
ql31LFfynx4cnsmo4dyLjh8qm0JZXeU7sKzUCLL2LRQL1dQx/m4ap50AChDOMpTJ
+27ppFdu0YWXQVRJ3kit8obZfGBap9G+BWHWbxmy2Ii/SdjGdjEkZS/kN1jzSFgO
oYGowYaDXYe4EXgWIZF+dGOxVLX7hEn87M9r3YXJ1fe/yJttIeMDEnbZSKeB5EDA
hxnFrht3azOQibkIzv+hLz4UoOwuBj0wi2qCtGsNgQGCVn54DoO7zSbiaP2hXXS3
qUrPuYUytMequV9SXaFz9QjEEmtyvrrX+Sxa8NxycMYgU3chKZhmD+LWGcpN0yHi
bkAPq2hPXg6TpzC0NsU21e+VkAyqU2xFaWOXF334HhU93INq/aZ4RpHG0fVTCUYh
CdW7Uc8P+838eie3VpNzAn9PItkL9gzA471oPZXpAZAYcssTf0P52ZKGBHQEAGmn
4by1iYMv4DRP+hSBlr+K4uQbwmlGMYGyRdauINe8J7YQEIQHQM8av2fLUqOepWd2
JXY0DajqZlNXLmS3r4BtxzTWF5TgtAYgqgxg5PZcq7aOcRhDKalikaRltZX39W/4
VxlLaGue3bsy+TLNRZiGeI4Ezw7D0jtYGWh9ZEULxUPcN4n8BzE7bQAK7dgrIFyN
LDtG+ft6cmp+CRvrgqEapSWIvIyNKb0jCRt6tVmDw6fgL1fwyyRtjx8LNB81F02p
fFHgYjoXRwfBlFP4fVAtCjh+YS3GGeM4InbU/fu88BE4EE5IGI7MuCldgxjEfcvq
Vtlf/p2JERnAayUYS3wyBKmZwBIIjGf8hJ+m3TwZQ2dj4pwTw7l5FBThMDDZuWtk
4BHa+6OFfVixHSnXRW7lckMxRvj91Qdx8uSnEYbFN4hNCq9MvO2EL8WFJaB/l2lh
Sqeu9tStvl8j8cII9QbSNYiPGeqWJ/6Gf/tpijbLD/8i+HkGpFi0JjxpurZ/Z2QI
b76xw1pa3n/ZQ5mmHqxZgupPGqxHP/zpIroOAnHDxI7JzplPqxkUAIFH3RPvxn3N
mKq8H1hJopgctroD5XWXUl8yBfmKbt77WFpu6ghqD0SOtRBmIh1Zdz1EraVDfcTB
JJ3BAeK29laiq4wcm48A7rLoYGZ+hTHMWWZ/MJUk+cVP0k07aXRpYxHCjE62PfRX
FbgNW0yRTJsHtwwbN67tL6nY30VA3VmFqnKKf7DwlJ8tilXA24g4nH/DOK78pWJo
U19xtT+w9emFJn5skkiazZ4p68Nze8E9p0Wva50Q8cEaKgNu9IAlFyFs+kV4T+Xw
x4aU5QlAGOCxf+YX3OW6wcUdVsbF9XLGWpo+shRe+KqiLMmeDuav0dKVx0NIT+Pz
uSX6mRA5kz55bf9BATQnsfDSy6TAAKeDoumBOu9v6uoVjCHmuxEPziMFZNrD1QMy
iEyaewzTz3SPlru+8SpiIuKVFWPjkrUIzeE/OSvpBd/LL454G5L/SBSt65QUJomt
z7PJsmPCzSZouACMLKdIEJ4jICYOQxFdBVpVowF5TDyLvOcxICMDHxFdRG2cUiVO
iTO3XofU+gA+LRVEEBQenwvUGcfPJcVJCTMiNlQt4WulZLjkaa4JrCCfumUYjQd+
t4iwpNUUbHwony+YjlyNOpzb06VjMJpeYGik/J5VTKeptqGbaYjtB2SUVr+v8L2E
IVQ/DyoMMUEIZ81ORyofyf176w/vAg+VLAhV84NxTeLwgtx65Mra4SmIDZ8IcYIY
4rxqqela5zAY25OpPpueQFwPRsNwpBB1vx5ecryNY8YBiLV3hLB2IUoT38lzJYLw
u5G9L0QvVvHTntUVUErTlNqYg75dJQuT+L3Y5rBq9G8fCae864b7emCGWcPXSipo
QmM8FrlHAuzwHs9EfxL1sBJokQ8IwKVsKr9fzHYLYFVpPJ+aV6oPXj9D26lYSMUT
n4rDyoPkFeIgNrDEfQSHQmVZNBer7oq6F0qqZSmzs6n2Z183MPLiD1hOmPSrsYIQ
pU+2rXa6HyevBCgCwoHDhopJWLVh/yHhyDhPoUlbDJ/ILfsIvhpdZB4yD4rG4tEh
tUqkLQAaDAq0eh2Zd7egrISne7vNx6mXXaW9tkBtrTZAkX5JDpZx5wl1SGgxVl4b
qANxRDCkD6acbDKZBdXNd3UaTOnqbDEpDUQRZMwtdvEnUK/dTJmDrGCpuvKrIQ+K
HYa3Ix06XiJeLoewBLjNGeXtMsAP8km1mHljJGYm0PcD3RB48+qasGsugWcsdn5n
vd+DV8FuV42zHz/QNXdfQ/sJK0i/pRgnnR2qvSMHXQccwxEVmCsm/2ZX9zIvefVh
/bICVEM+bstDJUWeKzPmtJu16gQPCJZ6WGjsTJ2lwAIxvRod/m4sMS6jhgkLMzeN
9OCMHdwHlGt0tUHTumxVV7oaTsIr8Vfv2QEc15FktUHEn4Gia2fvTo0Usq40oFMB
FawFeCSqESd4CWNdDHyignvLoxA3n4lEVQ/APO/edeaA2QhRVhk4YFDEijVp2xd8
Y7aMsBQL60K4kDdyAvjewJY+kShLzhhwlkYONbCS2zfIs68WDZoT80H5klGxDJY4
YRKTmwzEN5LrhJcb5thl4y0vpN+JIYyrQOPiN31QORU/+haBzF8eq60eNCtc/8Wg
x2ssYaOvykD7Z2agiFSBTwu3A0bDPoM2AOlMoTcyLtYg0qx4bL9/kfCFIe8QPE80
+FEYUKwoY05/vqWYgAL76FNJoQyGF3PMWRUqsGeyMCzSyvPJKZzDJNTJfioiLJ8T
L8Wxfrpm4vjZw6g6++sr3+rJA9AeuyHyuSn+82S7nmyYAgLQnZJDc550f8c3Xwee
C4dDl1+AtwWSVxPC2TiDOaagUnZ8gCqIgtI0J2BozW28u0S7YQXMLMas8Ei2Fkp2
VWLq+S0PJmHrpSThr8TfugWeM0oTJJuV8KtO+ibVhmGMvLsP3qJXvcIwNOuokai8
WRxsmmIf2JTf4wKs+DvheVYksw7N2akW2YYiwBhxcQQV3L2L8UCl+WwhzsC25Jvq
+YxYfijt0Vm1VrsCEOjGmexKUy/jKxNi1v+dPU5iRQFCPKMWtc3S3E9NZf/FMZVx
ZRNNhxlEEjwLNiMisvE1UXhjcE5O+xtsI4RB5eQqws8XrrHa/qroqwjkIE3jK1mC
aHt7RxFGBzfk1up80jNaZB2ii1pAf8PB0c/GNqAp2o7LD9vLJ/82S9C2jHEgYQXl
hBiQNuZc2Bkd/DLQT0WMRbeNqsAd2m4SeJTJHxcH93jjYdiQvchI1jrvasRac33L
Na/zYoSV+Wh3tCO8qTbhOOvREOBfTde/9QtD/spr9PEormSUG8Kywr8pnzKkP4gD
IN/d86QFCmZoxFAZklGurCea6+knV/968VwvcKBTQ1c7aJWxaWB3l/9XIn44xNJ+
hnQU5hxhCb7AsPFZLu8epPUVhoR3XcQlGhF/eAw8hiOOoSXikEqdrsp4sRUacylF
iYbmlrxffThr5zMowAiidgViDFx69FdELuToiEmGnVN8GNytDOqU/r1od/tEipDp
B/+vv3viBqLIpOy4KjQz1utLZheTQmPNd1k6KIc+AqY6eCqTeAuu5hEBoRwSCkzb
LGuBhUECMcuMzxWQat94d0M3eE3ps/VT/P+sGHJ4frZ/jMD6w4d5O67q4izZMvdH
MQJTH/xcJTdvgk0OA4Juv+VE5hffuQZZbjFridG7VDc1d9zQ89uNVk8bcgGarg86
4HvoD0zbnZLJDqMfcodLRTA38Hz8wfn4QEtPIUgdc4lkGB5Il+ej0vjwjQ+3bTEh
GpiS6fXCaz6tLlZ82kNYuCwhJ9Fxya4JHVC5sG4DAs//+5fMmfu3ybIqe/+u+PHd
zBvKgu/u8gLmRR00DtenZjiWqH6zcLpyZ752Hl6CnpEFE7erOFjBwPEmOXsCmM/c
SnNQZqVRrrx7glHBFxjVTNNY536z/A3WH2H0yDfZ7LZBBQEV5jPNPrR5CE0xkSSL
quv1MsLqmYvKydKUrNDenc9E0CJuBgrIeQaFiV/5+g70CNk9lj3lCsRw+jAGOTIt
0hBifR5/Xv3qt53VwVXALHoLMyUJrt20zarni1V1ot7wqoaAc1HWjcEa8AM80Bvb
lRveiKYZXg1snQNrY4LrwKI2aGFsECzNP6+WeEdhIaOg/8csezxfbedgOBhHBCzG
YrE4vCnkbMMKQNjDaGNr2nnj7M7f+aEjC/CzIyVR3FnuKust6zcQn4p3Ii/zroDY
RvGBNbz1ndl2et+MOykpuMF6JZ6TsS1UbFVOrDIKOiXDsuOkXMWWy8XIaeuwNLuo
W50M9j3QUkv/y4pN4jB7FtH+Qv+lC8wy5Kmm0A0/qsVeBRCDbFoJE96wwV5PCr69
PXtc1YP/mJWXOS+g/9EFW/6oyibO8bco19Qd/+1cNHPrWeK4qIodpo9z+6u08bnn
WSHAq7RQ3kMtlcRQwKpga1t9u5QCyrXq5Myym2LbsC0g9vs+HsyCqav6PSHhYO6n
2jJXN2EIC86vDBIMAheKH0vQ7XD76RR7u8b6yce8OfElUsOsQOND+T9yIV+gqvp0
7ByG+2HY15BZyy/spyTMBSc84R+ixMkIvhkH//GdJytFCzhaV2dy1I7M4/scWRqw
2TOWpLwdZXUvdjrvKiduoQ08oTiaStUWGgjX0s1IbKD3tr/tNSnXSYN5d2+82Qxl
h6n9n/YNypskvWoDWz56c+9wYcGNpyYbMyCUQO/DePtsX5JyZ+5v4ZDyQzul4N/r
NAGa4HSlerNZZUDyDv4YFXvScZBxHQS+KSwOMR8QxSHwF1iGCN74LM5aNVJM7yfz
5+TB37p9FD3ykb4DZOkM+m2aepCRsCYJ5s2jISGFBbkAole5+medXt5McP3UMPVB
DBiX5+CzAPoJ0gbQYDWUVuiqkbB6fF12wv60BHU6XrVHay6oRDzHZfdUhEHUHiKE
bED6qtPsPSCEVfZHE7aSMQteRvfGJldqPX9nrbW8ZfWb572EhKg1yNV7fFF9be6P
byKaNxwdfOxSuS6KIJGOxKSFUHp9iDfBwsstNAm+vw152ldIPokXHoOK0Nfz9Nb5
7Ik0c0p/rXlSE/JJdBRkOMD5h/ffrvB/tc9gqjOsQOQj9VM+1uQmfXTjnjQhseQQ
1suDL2Q7oufWCdusvtGNCGEzmTWoUR0ctMxcOyHehzsl0SWoC5JLRa8y0JNm81yJ
2zmXZJeyTUtNroKNee3E/kVI/oVjUoHJps0lzmsNcQH4Oic45+gxgw8k9OPsV6nl
70NRyhMckFyg+Dq34VFYtUBd14ns8zsF7k1A/NOba2CYIfFV4CWEInUKmHyDdefH
8rMUT4dqrYtRXO8VLHyyQc3PUU2gWm6uJTzAmrrZDKH6RnIz5qzhMFeqsMFlkbfN
TaHmSt189sun3bxu4ls5qhT0YffGS+pcFbXvTm26AcjJCEota06BXWpESvJootjl
cGPEkVhmAeIi6w8drNetXmQaJyDkX+f2W2egYzhehjWyPF2VIwfFDa9UkkESkkPz
o377GCTbWMyztqF4rW9+KQ1WW3KFMybVKp2ElHDXhBEq4obY2j9Jhnfrr1bNBNGi
h8dpoBRpCvbfxUjjitRhoi6iNPyr3QCPudqX91K5syfwCRPWBsR58NjxklZd7SjZ
4CTwfC8F7evzqKtjr7RRdq/hNJvzxtPylJqwh5uyjcYCn5FqGBPYRLiAzJjCdmEi
PrLZi1w10ZBn8XlH988TyMMgazEjGZTZoROD62Oxk8nwUSKjdz1bKgxODssdr5G/
qLC0rFaJZHGl/W4TbBl/+7qY05lBSKls0Bp57jIEDX1BBIqrYxqd1xiAkluAWh4S
ZAbRbBturkt2NjBPYSMEXkqHA/6OWrCjOlrF+HE4Gvk4JQFXeIDfNAl9+Z05DKlL
JqHn6K52eUWeuH4Lj1FJrtgeAs5VqGo+CNETXa1ActbMkkpequvvaPX4ZTD/nT0/
5su+nI4MFasi92zTrA40g2prxaWlwjWAnNwjmj/eoFUtw50r9rgoZGnHIHapY9SD
9wXtRlQLLDcuIdiLZTyyTMbW+xwLl2s5q8VzsjK+cUd2EITnjPiNJ7qU+kKfZ4ki
CjecJVi46oVqaOztib95Umee+fZVM22umCc2l4vVlBC22ksZwu4XwL6U3hVIPlzC
S23zG7Zy0fvNYVVzBvRFnpJEvb9184EXcPis81yskIuMeAq96xLSgmd4gBtMQ5RZ
Y9wI38WwB93IpT0pXSFuZfjd/6PsQ772pIhxzXSinmF2MegH/Dp7i4XpJhbfDKMW
3UKdWykV7+4avwW8aRuZCHVWwuc8lJ7P9pm/9v/YHf6Oytocfzr0hLeYImBD6COo
+L59UlrFvvnxExUEQ/NuRt9bn9kT86MCzfYKXFb5xo7EN4SxRvEYdov4FyhgCzYC
D6az0kJLrX2riRr30qMeYb/O3Q0cprimmZ5/QNYPMcNqVAssLv4iNbMTsfhdFO8r
jQ/mCC/uYjtG954IGtjp0pneWNLTrUsSYLPRezZbW6RUuFsqDEuYrAPvBoUTLDe+
5EC+aU2tLXd7pRwQrCayba7avmS/pzaac4fUr/yFs6NfRcUNPzFW4A+CBIU8FYSh
PX5EPInyuOup2vh7H0ca4GlSNPthXFsuvIaCZNGRImxZwim8g0z/rl3ph+D5Ze1s
tKt8Vb7SI0IiYfIq7oFkbxs68ZSgir+KFWVclRk+Co9NMorMOZFBMZyGITQ5PQV4
sWbwCE8MDO1wwUukJsruVskyAqv3C2GxcaZh9IjZgTSbSyDg2bExtpDTak74afxG
+7usFF85JZTR+dYqXIfW2b+2fMz3GbyTHH0ur6QdKGYKlReHn08q83TH6d6vlgqv
sfVXg4Xsj9ABMdWWI6u7ZwKviuIFgQqFAk1k6WsiIwLTl/f7aZ6qupUKpWmoAIRy
9PnBGtsuXb5icQC7M6ssNa4vZSkWdeNqcwpl2i1H4jt8V0M6EaRlCcU0hjVRRq97
ZNC8T7DcWBFkPGGpJgZMIOZxlA2Jhn3/1iL9O9Fc+YhRRRIpZT3V/qIQjFg3stbn
+7YtSjaDBdMhEtJoq+6WZbYIHv9bt/mHJ56nO/gfB66kqhf4dGWvYtt2ZKr4CZ/b
dJl45V00fEjiO+vjQAPaZ4Unf9vF0v69ppriZugmQtc9DOJsMnff13RTWKSHFA1u
kMGbI2aYaXTaZ5kZ04mXbRctUFbgVnb/03pd0lCckZXq//VswQMR6nnULPTrXM2p
OXxIBe/BXdbT5c69ntQVenULhPGV8U9mEe9tiHyeIjLEwZNBikViu3reZh9Z5FUN
Pk5irMQRM/dmXqh2EtKhi9Y98q92cG94dqtpLdVujAYh7Yf1zu6qIKKbrvc7ZVVa
0QuJuM91gE/40VkoNNdJuPQ665sphiukI7yFYCft4AZjddvmC847wFkuvFXzOSjK
JsmY6dVm9wqRK5O+WnY+QedUIEr91t6PTBiPKH4+E4t5vqmT+wYxr+rrms7I/+M2
q1jHXNFaKWEW1Vms1Mcc30z8mG4Ij1yHTEbo4sw0XZcNpZHuMCgHZmfeytWj8N4/
WJsQEvysvTxM7k7kzQA08At7FrhtqoKB6vMA8QGgpbLUTwHX2D7ZDiq94UoPcSG1
73i25rXWDHdQL1weSYwY4nLZHX/w/9N4+FuelE3Vh8ohN5TRRwQaEv5kZ4lffGRF
8Fq1mHUl8O+y5nP2Yb2MaoY7bqdZVF+sGrB2Rwm9gfDI/Sz2opkWw5LqKKtLqau2
TWdnz3oP718lE747Ap/zUD9TLhjkJNraKNgpUMLKf8Df6QxzlqVrevmp32GXgKSZ
lbQlxFxS3iFJq0snw8SSnX9I6CH5tAQpoRMLwyAvWoIE9I/g8A9WLjCU91wW5yll
IOirc0re6z6J3CJr5lcsU7udcGvI8nz/KS+Y4XrwJgphygurwC5cQbh4s6+sr1W+
PWlxGDbcsDgcdU7NrAlIp0oKwSTEqLHJ7E7Q35N5tg57eS65qUCSKbkW9S2zpvPp
QQme67raMRBIHzacUCjpYAGFUTf3y5nIjFKA+A7DtH31SPJCRP/17cQj2owreTV1
1fmY0yx6WAK/kOMCevSuh/AeCrOXui2pvRgD6PxVn5PkM+foUfXTePr9JcrmVz1R
DgTW8PxCvy+oZIRYEc0NpqNyXLVPggzVZXGbuB0wE+BUsqZ/RN6rkqvtqcUyA79F
mYBIeO03FkjqsRE7/pe2yGhAFHeKWL+wvdGnkdLM0PA28+w2b5nOLLXpwiv+FE5a
vTScFjbpbDeBlATRi036DGFT2CIPwr64cCkaptFoU524LPh1lC8dFf1SiUbuj09T
J9cIpQQ8ROdpwwDgdcF2UysUGEhS4Wvahy6Io+iYWedEzXGZd9qWwRvg5HnQv+BF
Me2gaQYTiYDTFcBN/mp+p12r6RlDV3UUnYvp5fWJ2niqfkBF6DJc2htEJHKEGvMb
2ipTEcYM/6o4pxUF8VSWAVcj7q8bcRBwObFZd7JNMiEkXv2OLcIvqLK6HKRQPTM2
1QvbCES4wMzU+VWB9ii3Uc8kRhLbkRJx9G1SQFcEFWeoS4UbVcSih8S+BsTuk9Em
ES9Vp7EHDMKRoKsfEmBTVYvw5mmY8CgnNg5/Q7lTJOOzU1PuAD9cK+aUToYATRYb
iyIZRVdJfvIjQ0VlEbddxf3OCcr8LBUgyMRWxJfi2waQDuKFjIkd2GCb2CIi/RtS
1AMiBLpnvrBaeAP5wkW4QXtAij3DP/8LamA4LAPIaKaBSlJQP8LyDzYgHvQndBVb
c06RCN2U+oeyHbooEucYLlTR+ixZaZ2zaZhlfufohexWb5vRkGvgasuBj6RFNbGG
QgBm5LoqZMH/7aLaX0njQMPzfp362wiarLCM3M4PT+ZKEng5gTVq/Jggu1RbZ/CU
emXsuyNniib2O9awQyL2s9ee0Z4otNZaj5uop/ZyaCSPhL8wKWfX0OScpmaaCR0q
s+jN/IpmWRWjN1vo7lKpMh3H6oA5+MmNUsS1wi66/2u6Sm/KuawgAjqRcBofv8Tt
2g5aXlv3UdWw6B3dYRfAQgXi1cbaV0XrSCkZ1BNp9DKtOmUJElASolR6zPeQ1MEE
Y/WSIuU+OxwdzEveQJtvIK7ylUSWiUmCIZwizXjjXQnUESey9jVrPFv4QuWYavfi
STqcdNnVC/f0u2NcrN0kS0aMir/ZMYUItNn4lD05hYK3w7sLIZeyMVBAhEWnPMDt
rUhoc0zZqC/pPn2mldiUHYM5m2UNa2oBkE4v4vN3EgGbknPZVmR51GiljfCZOmZJ
nXA8f9D9aCD7JilrkiTCbF/49f7zADru4BqZPOhtsgoZrof8xOEm15x0RW8ICnXT
OnowUrJ86NO1Dkbw5ZgxB7A1SZoC+/DEzP1O9u5kImEqE35BPQN7ZH15ykNef5D8
8ttTLnZsdHWr/u708Xc9OlUPIFlMaP3sm7D5ep9iXZI6or7p/fxaiIcat/Pi9K/8
6LW/3mCL0I/J1AjjYdKFPi1sGe/Abn+5edVUMVlcEEBAk/xw0YdndrW6uB4cwsu7
wle7qkIbJo/kyQHnGQp/4L9Ozd/TCuZqSyYP8ugD3mbw7AWJRcIeLPAJ1fiJ41DF
KuuzIYZhwKij0F7N8vSx6x2uC6jNp42w53bByAJYCoPKvj86E7JF64Wg4QuMQkg5
eWTo5iHDNlqtL4NX9nsf3yVzE/U0SWCNU2BqOouAb5hECOi347K5otDY9LnpKjj5
cD0IgHpSWYfewHDL67+CL7DBU0K73ei8HWxHpFzNZUN3+0SdW1WHQeroaBnEGExZ
fI0eAryjsb8Txoe2BfskO4q2SGpNyin2kjNFY9eBdAG3SV37IgjAV5RxJv+Y91CD
/rQphIl4gd+cQbB0GbbArfBLLykcRfnjClmE4c/4EBe2Y98SKsgI6YfPhs7xP4UG
z5Ebc/xpcQm2RVCX8RfSf+hXeIoEb+VzEkSjqJaAaFGZ0sf9lyyl02xFiMCKeo4P
IX2z/Qi17YgCWx2N+hUzc+8XETtPZFZu1W3fjEQtFl9l1ZOVfADN6Gp4nXkNQE+d
L3W833Rn+pOJUGJLtCfIqClRH/0RaTFDm1NwNXvCFM/JqiS1fI12e7rSf2ndQt5B
QEEhmT8HisEvIubZj4FwayZwhgo/R4ir5pchzixTyK6tUJ8tvh2+DxY0lLtxv2N9
IyOEBoDjzBHCx5y9I+JEXlTxCyeqMROVfcfPEXc9QcXs1r6GLK/OSqYcYe9ijcsL
b7mqaIISixB3hKeh2b1qzMPqhKfAAwdPbTKN+CxpVEhm0SX+RgPulWgVGsObBzcA
AZutcBBKAPc2lZsR8YEmLM8wpmAp0yS9RX8TYDusuiCi11QEdbKIyJz5vC2aoXjU
xUSpFM2qxv2c6wD+F71TXbo6/MwSMCxfTaQpXBYQDguFId5fQu+7RN6XXT2htkd4
0t/BXeB5S7B7ScarErNv7hLa0TEk3OFtRfn3HVzabS++jtUIquwwlrz/cX0Y8q/R
0nn0+LHPxJIJLS33+YI5Y8RDkyJBRqGLkEwVKDT7fnQHNJyzjdDza1Tgbo2Dkji+
b2vpdzCLOjSNLZDDtxQfUCNMUZZgr1ylfCobAIZY+RrSzCOnjakPJ1iQC79f/+O2
96sxG5wK1Rc0CUW4kFRHMtBuNpMDO/UZ5U3LjX50Eh5lD6rhCFM7Ciuwto6l6eOc
jVnsbM5PEwyY8Z5E3zpNXPp28ukH/G8cyhtMBfUBRmxdVoVVcip9OY4BHw22/eCP
qbO6DmPcg11k75OFHni3IfVN+3/6z04+QhqACLKQrdfoWmvHs+wgn5/KCRDv5nZo
fUkl0busO7zejk6JDj8y9BqHO9UyZr2G8lfKj7iMwOglmxwqfNMcXoCuthMQBuf9
DvtlXWXoIWaiFl7X34qL+yeBhiO7dOVLCZAL74CDvxZziGvnKztAsQDBL3OS8b3y
NyMnmVJL9RViD4uo45mmah+UDSxI+TJFXSKBfsDNN4bDzbZ37UkaBjrTkBCiGiA5
H8J2BhvnwZ4eZwZ4kQAkPhFNL/wqm/4hKf9G9uKSKEZhU5sB/ojJHo/S1ddxW2aq
nzv/YRHNA/HsK1YBho+lwMkbaRf23CCslD89kipU36CXYBPj6SaPf9eYAltPJguM
7RCrJgaie/Q0Q17SpwCKuoIAxcTgev7qmOOQUf/ooGWFMy7HDT8W4GkzgtL5c8wJ
R+MDr/19lnVGDl1IF7QBtF4n4Cdr1YSUEIVaJfmvL9l94xh97iARF8ouyUuUirl1
St5Te9/PvsQt/lnqlehYmsaw45zEzWWolkD3EoBkOBBRkPtFsD5j/HV0kWfI2oU8
vijccGGZ5R+S0W0YifhW3//UgkMMvDq8ea1eRHOdiuYoLh4zav/kBgS127mA6L2p
UxdUVmoPu723D6rDRNR+D41e45VbshKsLclymHJe/o9xjJXvSQ3E6FD/78npH6g9
1BwF2ibfocI0nF/dsm12FORvd61mN/q2g7TSrKM1R/I00zQ4wV11c9q1nCPXjypJ
K+4oBBNIipnDbvI0iSCx1wXKXYPK1S/THBrdh0vRwRH+pVoilVD4aT3PuEidlTAV
66XEN6QSocUdgj3nGDz16wML1bDraqZTc7j7F5cTrhxmGrOMPsixp+xoGZJG30IK
29RbM3640Wil/ANF6rhssbznFVXXGQHlrL1rG20LyIrba7m7Zbd8X480UJJcxHxq
CZZbcRoBidyiSR5NZy0BfSe+v31Qc+7fNjuUZI+UwZTL0APjtny4m0oluB/e5kjA
IaHqj1rR/L7GRuU2yeOVUyjK3C39FnFsliCqh9g816txyh1r2XRQQ33XtR0DynD4
NftGNnn/Z41TPfGE8Nc6a+Tx89dfRgh39Afr9R4PR5yBnqHdv0UpsUKWFIeKTJ3S
oE7G2jFsEiLb3nLBnbMYYdgfSX1JZ4PlJHH4T/i0L+vagFOGFr8grQcHvyEB8fM4
Qk76A6SZmQLZhsMp5H6+OlMk+JhY9GMM0RmjXwbFu7ANMydx/1c3QvlujioCewQZ
+ziJBEMDgMvQfHNDqO4Jkz5vJa3MiBr6oM4ju9RXrt1d+adaTgITdDkpM/A9q8M/
t0a99J7EPL2lB1Q9/+3mUbn/d6z3PeEkGOvxe/vLOzjYToDUoelYGCxn5bR9rBhA
gTHlShCBWVu+XS6qPQ6Kz3yz3oTOHPb4/K0V/4QJgb/rZIuamVlxiz4bKq1Nv1wV
VO7/W+K2vzGhN8phjtm+ntVkKtqHtNSSNwQ0r/HbYV60VppkboAdTQHCLjlhTVFu
vTmGMyjJ8g9HC3n8/HhvZXvQUzkVPrmebbllhgOe/sIKHd19ptqdjwTXZJ6265at
4w7Cl+YVjUsgBOT/pLWiIxZAfBRTxTHN2YiCQdMYohmHapNcbbfDmuZ4FXkjbQ2+
lI1Y5kFn35vO/AugQDzaPJTJf+UEObft/cZcBLAHpORBWKukF0h+F7ORjmGneUpH
utwTHYsg8JSFAvCrD7gqJYv3KF9zpDLfwkOKv5Tkf8EQfeb1/rPaGZyvYUvbdVPc
nJA01cWAqOuiRl5Ep3HEZtQw8UH5vkYnfNNTlNnd+/vybA1IqhI2VHYZsLNjBQrO
qQDHTdllXzkV0pzgBQ86FE81VLplJENKnuiq2gz8rFmWnbZuzi3zkDJuvANfa2HY
jeiz+N4h1o69x03MejeglKCXJOHhaC6gLbFjFblIc//rpF58BJC15L84gltNfNnm
foAuKsbim4fyo2GLOZPCRKfk7IffZWg5a+Ok2JYqRd0w3Wj5iMo5Wu/kRtFeVP0c
yGejPJPvNF739TZzgwerSxVrlYFNU22sekxIUtqbL0NLf5a7xJbiji5d519NTRf4
KO6gccka7AEo+twbLU2nYck57Fvjj15A9TQL5CHQbiA1n9s6Q0ZEEq3j4eomFHM5
H+bjpfN/VnmUQQ92gKbFC0TChvoYRC+ufTTycl5OmoWDLPuRXgQYwOjrJM/Oi5E6
WEpQ4MzVmMpue+VhzslSYa6jsHfNSOHv+Y/9Lu091r4L8WWAl5Pb/CyNzJCvaVO7
UU0iCMt5iCBLpgzOgKrpi4mt+79H6XDLzmXfqSnbewZjjLIL37tpNcz4JgTQp673
e6DH9xtsA8rG9MQXtTer4izfKtcmqACJLdWimfOHPPGOyqY2KWSBak78J5P5f5ku
v4ZZNQlRgg+jNUT/Ys2yaIArR2zl6hjzWMIE9SZsSF2wNlFS25KDRj81JFWLUz14
ewFFaFZVJwuZ6hTO0mr+TYBv2kuYx5uNe8MkJgfr4PMyOWz7VFu+LIsO3zLD4/9+
29jguIC2MkGQDDqfXmyWLn+aHHkY1bzyh7jeqsbwwmDXR0HVBjBq3Ps7yCHtt/DV
k4ae/BsCXXLBuMly5F4WlfjJ2y+GvR53MytQHn4A73AqxIWOZg6ZeubmdvHme7gx
CZkv6zCwZRTIZLzkty3a3rZKf+kh2LXWEqBUXwM2b9FSvPa6AARms0WO5OqrnRYg
RKqclxbCYdjKDsCbAFUEHTB0WYikibvQc3frKb/in2NdFlMYuIJUymO1BJZdTFQs
etB69tFw41HT2isdFMGUuwaZbXsl2C0HK2bq2HtMZ4IdkCvpHPxnf5nQRejbpjKN
B+Gcnrx3Soi8cuPuG8oZ0zJXlmi0f6YNzJv5rF5xOSP0kC4mHgFkolVwC1T0GC0I
Dn6EkwxWOEUJHvH3KODZfJx52lCc0PlwrYYrr/UWOivV8T5nI8yGb4D1ynnQwOrF
g020bYcWmDNPj6XNhAsKKYRZRDllpIUBIHtN6ArbfaNLI4HE0D89R3kwk2qG7bBX
YixbLggmoC5ZQHD5JgUsX7hVE8LU6HdmADtZ+k8ZF146Y54MpkJejrENPsNBTPFi
JuCnHenECYD+7H6AJNo9BkGjZW6XGbTNlu0vwgA7vnxDEgnpUE2p8QedIju4YxrY
XGcoL6g6BxYrzQLb2Oo1VSep8rshzpQbHT8G+9rsMwyz7OTyntfc3FqXARjM3gY6
a4vVh3adwidchlwdX8KEX5lX7eQJEvUaF11g1tD5jh06gKI8kcbahQNv21K6QZ+F
O+Wn5JtpWx1J1SUrk668D943obIa5dTgqiLWEQkBRngww2wqCzDOQv/OFZf+tQxE
qVb6RVP78Cr2jQI2V5icmhIIQqFiAJNTSh+1KPIzMSCFpJ3lGBMzSAFlsiQRAdXC
blCg6JjiU+x3MMqMhQ8FB4F1oeL6jdLy5WUFtcjgv5SGuGBuCy4LIreE9UN0YMR0
gR2U0uCsVXLJ3grxNr+/PiSVxSZ5XmL42PCEnsNXCVGhYIDr1tF4b2F5uEOA3KDL
trEThv9wsILaihrSWpnjRZIq8TcEe/JsD3/WkUzpRHRSpdFlsaX2qMX2QnIdbvgT
e41/IgGOZH1g7qf5BNGfQbX+7X4NO9spbV8JtHE23UMtroP1SHk8kcp1rS6hjjVi
7fptxdJkiRlhIXGHtCeA2SpvF825WZHU4THoRXCkDkQjEkqVuxvJkK3tjLukyTq8
m3hlAsR9B8E5C3PcejILq7ztqMVrg46ecwyDtx1LZCKvvDCyIqh0GRp0wKFHT5R2
ZXS6ZKOGM6LT9Pm4ix61CBLYT7Y8gcwKDoJXfvqkWKqxi+OomcfH9CY/nP9V2X7G
H4G5l8aM/3H6LpyNwL+A6s88a3BbEiHQbkQ6y0v+bDWv5jU0Y8oW2tQPe9kD+7XA
r5jdd66GyN4RBEKuUXuQfX8oLpAo+cH9J/Hd3p3t3V32xgpwbaQYjloAK+5svmoe
JRxaTJVjvjwiTzFtMnhNK0OxG1TLccO6RHTzyAqCodK5XTP11KTCMpMYcT3UMmdA
8eQBMukMk+G5GWxI1ejKReGGR7XjCWxDv0Yu94AE3szDC+Ev32mljoWLL13fa2Px
4JZRhA2ZGySPPiAAWGret1ZxPdJtj2ZD9UG6iEqT87CEiM59VglWM9RaSlBLH+az
AargHII4NmxGV2WcJ5wA8Ube83ai8QxAkGOeyX/3JLlm4ihy8uxzqun8qyxCvguB
VuNSOh7vSMNL7IjcTZ3Jcqd31HG4o4yylOsfO4XviRJ9LtcF2eHyetufSQsvhgD7
pXhO5QSSw0/o83RG35UcUc4PcaCPsy2amASyvgDgMnaBIOlVsGEnmckFtCbul2hW
BbSiwuEt5mBxGbeHroWInlMV6I7yjpmiz3ipgXx/E4JBJAhf9CPYsKVZTef7LUuI
6Czj9XEyyjgg+tX/nF/Ic2/71wiQ13S/ZSsJDxLUcD5XFo56/x+JMP2dAMyxLxKv
+k6j6rD8NgKDbzxBCQdcOwHE3SSBhuYxV5BguB2SLVqGFMlz9PjopVm5TQX0fdeE
/0CsmHswH6e++ItWllBSq7Em/rWx2eIM60qzj1+ccYYUN9tftAfNFivD/ao0pVqJ
BCgmtZnFnI5ocUBDJ2cVyqJgmy+sX1xAGMBxqNUjvua31CMm3cfmuDtBsgP1YB2U
wkS88dWcHfKJXYC08pI+jubOTMp8V7dVWYBwlSj6VFHEd1czGinZdAdUJE8opmcO
xeH9OvEY+lplD3hwKkSHr3XhxRbazeqhuoDwYIQCW8uWQm0yUPDYdE4Z2vyVC8r3
GLoQvxq6EfDauVIR6AMG9S+HoiS0q/J+Eodb5n4a/ylZ5Zq1Yw/qJnmM/gHZjTAS
YcdPSpr83x+jVimqqMmcZMzKv13GiyvlWvvYiN/Uk30euL+6xJE41BkYDK7SjMBF
iE0V3Yx0VtYkFVfgwLcIrMVM97pwcV5RaOwbLgQtt7ulwxuCsScHQ9zK3TJ9c3Xd
ZZg3vA4h3nIF/xCbfopnKO/i0XzfdNRHimlMQPZ5Io3d6wGhumiVXlvMKbZqyprV
+j0olFhkvV4TyaGWNlgjJeyZMpRk8p66ZEabYBecTn9ghFCadWEpyge1PXGTEym9
D7eQ7pSX0RsWBBisyW7hAB1wVJ8anbyVpKl7X+C7MfuUyG1Q7OKY4jU2AEfObDwr
FG6xQIWKDqMsGCbEZMMqtBI6aNiPoThxKhcS1EsuGB2I+QozqD7zKAkea1bGinjK
+o4jVpQvrpUkwsm1qDRwOQ==
//pragma protect end_data_block
//pragma protect digest_block
3ce5ns7vmCSJ5R4XQlfu0nw6+SA=
//pragma protect end_digest_block
//pragma protect end_protected

`endif // GUARD_SVT_AHB_MASTER_MONITOR_DEF_COV_DATA_CALLBACK_SV
