
`ifndef GUARD_SVT_AHB_CHECKER_SV
`define GUARD_SVT_AHB_CHECKER_SV

/**
 * Class declaration of each of the error check stats instances using the 
 * `SVT_ERR_CHECK_STATS_COV_EXTENDED_CLASS_DECL(stats_name) MACRO.
 * 
 * Each call of the MACRO would declare an extended "svt_err_check_stats_cov.sv" class
 * named as "svt_err_check_stats_cov_<stats_name>".
 */
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
mqOyJWnBYY4LgnNgSbQATS/eTzzEVUY6AntbXVOJ9rCozr/obacd4Hn+zr9LsrMw
xE7rcCv5gj0b6jOUPPyxUMRRjTMouKK46b47VJ8XbEKqT0EuZ+WkFtKXNUlMvqE6
oLwuwEyA3Od+nP32OJs+HITA1ikl14LmVaYSE00PahBh721yLN3smQ==
//pragma protect end_key_block
//pragma protect digest_block
NeHH5HxtDwZpgdalwzqyPtf/hQw=
//pragma protect end_digest_block
//pragma protect data_block
ic/dHMhIG8ZxgbL7aQIPunOtXJx4OiNmjaFfekN6U19eGAoUSR9mY9O7ngkYUwGu
PKHApw4udFKpHvbOXW7ifONi1Ck/dHCh1qELaYtYpOJOz2e027jVcPu79soyQfxB
vwGL/cmtSHigOoxQMKoFP2MnzbL68KSvAq45XO19Hhu8jFRFKPlNyjm5mGeWsSax
phe6th4VNY4YNJ6qs0QOTLnUQleAR535rt2K0XVgy3E8qaqTCarCdBEqsqFjwsXV
nIc6XQ24d1iygNkuoVXRpkwzdkYy7V8wZ8+1D/qbTSb0qZxT0MgVDCjL9AUS6HhM
8Un94XX1nb9xB5BKBxP+qvhFoBRaBRWw295rXdFJcCFmG/YgT0l5LXJeyNCWojNT
C1k05PfcVv8dRY+mtoYoX0hCl1oo3vwhb9DNF/FJiaWsTrqC5LZYRkJ61VN9pXnS
Wz1S+NCMLcHzBEZvrOJtLKzZ+u4oo4FqjXyxXtjhLAlJiT/YniLsus1QopU0WUnK
avuXmcIzVaJIL1mLry1ISBKT+bcfD9Vij9YKUc8QJLp6Dh4ni9aMLpDNXglBnv/n
LoMRazwxDWZ0YjN4CSKFRshz4MPCvQp6weBXFBN9Vr6ejnX9wFxvtHkgtphL4K2v
10m7ZwnEYFCk7TQqnowT6l3LxnCpLJRoIn4c6JSB+qhnraXZx07E/N6QJMG60+jX
v7wIy5iQmi4X5kC0D5NVfhsY52DqIRaA1vhvAKNfD12XPPxZenCJkOgcc7VVOQV2
RB8PpuHvfEQjSHRsp6FMLSwOElJ7DNPOqZSy2nJkNJxDyF4XuU55acSVyVpIJ+29
hX25VJNawX+rr158FG2TBvYXbZS+corarWkaOWFq8H/FKdglHyPnDJjbjzc5P3Ns
R7l0WXYguETWRdmb24QFleq0rX9owPoRhcQU+TLvzBvT77HEXrlPLodHJZWyFdvo
HTJRXbb8G1x6CbPR69vSi7c0bqMXuzHZy7DNGCle3MauEQqWO8Z34UGFosrVGjHn
/DB+cNoPnXxCobugLfcP8vyfr+9VT6p8CrK1fe0ozBXmNPBPF/+GCR33yyDrMGJd
MyRUrAIxfX7CQZxsRzoUaXTUrbVT6m1YNx/Ya3QGkQ0T6/tT6pKpVJKtQ17u5Y5r
A7aFAfqNUxa9B1EKpmi5Ou6AyFvcYcFqVMbyyk7aPfDOsrM0mx2Mx0esVCsCLQYP
a/TcqGrmX5npZCxapjig80XZH6YfcJ8TFN8j/cnOXFfKMs/kGgZ043Tvl4PEarWE
CUqS9mbREOjL3QiVpD8tsj+U4y1Qs5c/nRTqH0xbwJtPaVfixd8XovedX2h9tN2L
8m7WiJu66pN6TebNqAA48IZtYAlGGYuAqQdY3fw66HS2vYyXebbcTKsQhws+i3z8
CmCMT8mzDYL75k+nQ6d14OQKbZ4b+4FU0PWKFq7m/pWU7d8pMSattfgzUcuQdbNH
oj91KyLx/8AydllR5dDnjDRL9VSkG9tmOrUld0Op8Q9Sop6jJbvjsrHg0Cc5ESBf
ApG0MB8w4NZ9AKaN9cpN/XZ0XVWwsi35CemoYgZcZ3Dqfoc74MiXI0msh39frXKn
SEkyVdZGlT7iPNk1AmTr8pGpYhiyTkRO+MExzo6ggNWZkhyvFEok3AiKWNChHTA8
0VxBAoU1SgZYyxCtqwIj0h/hQjY3Ha8r1YWKDpFwPx93ZDT30Tv41F0R5bbigY/A
1Staood7AVDZ5rHwuMUHfztL8hMRHSPbK3pzN8ZSTpb1Rct6lRFNKNahQ0IzMzOj
ehtfx+4bKdoF5PgQtRtyIHmC6TKRbwFt2ERiDLB3ZO/eUrANe3oYZFVfialyLSxZ
yivfWWawyIID0YaBrbIe6Wb/eB4CKPazFYLBloOR8s6BRUc5eN7UR3/wcCkcSecS
9MTEHKK7E5GeVZGK/GCrR1LAJywooPutFN2uI34ArtOFQMVVDFAPDMnh1mms2BO6
HwWA3xJToAFl0BszfEMlUc1MlHP/D/EbCWtwfhKpAuj1EgQqlkmyI/H+/lA8V71i
x1dV5sbL//RxEpCtVlmdfVk+9gmW4kkVx893JAlFOvo+7HIYH5SQW/7lZOsCmWif
2gDpRL3lBcWAtwS8PrZD893m/8CAQjwwNIc8COBnVu9p6OhpbjGTGsZrjB5bLx76
nh9h1PdsJitYnTcl5s+IncV1yAvaAQ8MHElC7v0LP5G5BGR1XZOulPdLPEwWoK7e
pFudGF4odu4uHX/U/r8h9QktI6I+efxQGOFCr7W9AHrnCBnXbsD1wAcXRQOEIyxP
XgpCsKLy57eBKHXK7ev4L9F35pqoGsRv/g5S8s5AYVKOnXiRoj2dnzjAK1CDE5RW
QxkKFVIYMF9SAS0VNEAQv7WiYVKPBTc0w11VCcVH2zxAR81MJoymMz4ph0GW+G9F
vRhGJu21Ra0Me9Ee1gxZBOV3ZF3AdieMm72KBaYwgw+DFH0p4CAEc+JssBxJT8dz
uR+xemV3YoFSkSQ6okPOtx/mpbCaS+GQ+U32GJxBYhm25ivNhzAq20879eKVmEd3
Yrr/oFAAe5g17ndUx0aaeoWuG185KwgxFJzjBwO6VKhAXsCGxXnQPihphifsEsLV
XDODSF5k1rDClTQRu1fWKasdpGProVjP88cAgMnFp8Swedz0a/WojKL23r6tDm/J
Bm9s5p9y6yP7ZnFCcOYuSZNBh2grxN+CxWGt+UULqmLq460AIvMHCA1cd0HpEA8m
KksS3En+gbWzJkf2Xq1F8HJTk4LDd71SU33niGd+SG0ApY3QS27fF8DynbgNgnoT
u6SM/5z/+No2ys1OASbWpSVdnTN8YhknEnuQSQaPdJk39lT+/FWuTLSNvNctkcbX
YTH96cIPwllyMFfHC2gs7oXq2m10e9L33FFeGmmWgElNkVPrgjXX+12YlBBALG31
yHkczu0FX2ipRpuokJ5ZlI5JNQZnWZrGqvJrvTBbQmRU4RYAOC/DGJPujwbFeE/c
+NXaYWDbp1vbMT49SsxQoBHjx8S/yclAt2Lhhp17XC+CHCVtNMJXXtvIYF8C8MGJ
L/iCp+IJjCCAGANvM2mKPvU74X+1eSIxKKDwxoKJdbowWOsxwmzxp3FwTb/d9YDd
lrPPa8GtC9AAJufHBwWwQc6deir/IVs/8pbdtIaej05tLFwvbZaTe/FK/ZI0bXSb
CaPP4hm0ex2g6mU/u5hziQgkYi3+vQPsc+pPFsMiUU2so9iche9mfGlXw0FZOdSW
uOm5Gz07SldjyJkimRO2y8sGhUNguvAsMon2SgGyZhDvzpQQvVMvicsbaS4IRpsr
YJtYK91UvHd1H5YP3gBkg8FH+reOff+40DVNgYB2H+vDRuyieWRslwLDMtWrFoK/
ebNtELEOP9f+FtHOREwzSAfdHyqusdEjxRPW16vueBpZql/IdgOXbv4wiAXhqhKK
uRL1TSn1R0BRHjiVzMT2fiIG/4w327g5TOxpkwGsQxmhhTD5n3+VhqMpvefBb4X7
CD9ZmGcgLuxhTJRN5mXPWjz2tNGJ7IEnh69qIZzqPecOAMoNb29YtVU3f9zMhw7m
Am0Qz4HDZrFF1Nr4tgiHIYMkEHSlLDJZS9ihuvAv/UPvA2Skdhmj21wUeZifJBDB
sSQsbxX7kNk2A2bB3A9SMxdzYiFIW3gGAUyBx9n/Biug/cKbTJ+HMD4d2ckPcgcD
CqRA8CuFL/fACF0qn/HTc0sKGeUu51QKrC+1Cj/4i+6y8vmi9nsPlUuIyvi5U6qK
sjYVEcOnE7omfjaqksdJpAaHg/2gZvnawtFWStrSdBEkarwYQY2jQh1+prKGNk6z
cRYdYrhYHLs+Wgm3IdMFjJW0rA2czjDPCsjOAIMsU3tbzzcIP3b4OmYFf+lkAoGG
JFbg/zHt1U22eZ0fS0YWqdiEWQFR+H1hdcuR7Uw+jmgkT2bNbjLBz662E3eqAkf7
W/NumF5+8E1G1BpF8hLrOCTCfmwTT2RKqYoEyDegaDeyz3/iCgqcke66suJSj2pR
/aSxtuC+cwgvT1SB6N8rjKL2eKJJpSd+LZLyJMhwN7ME+R0QzIwcDRXobV5oq+j6
3/s6HgwzVGB6jC+gQ/KoJhM6QDfQ8sdpdRDTsVtzYskpvAYkiZSZFihh/IE0xdWX
xCk+jr7HoQpJwLzjAFjOo/lVJOnBOExZBBUD3JYC0gEPvr9UhhVnJIhVUJ/oyscV
CpOvaTWwTXynaqCwff2Xd+dcaLxd5nF+FDUkb5LdWMZMVWznbWAEnTSWS7A0WqPw
EIA6HGTiTsnO9bQld2OJ7oEGoqUqLmLc8U+EZWAHKcMhe63XsIHt5tUR6NkOjB9c
p7nK35ChA/BeGlKcnvQavoke8SwteXP+FJcAIgvdxsN7yyOqyY4UkxOH5uaKaHy8
MnkQ5DNQ9cFJ2iWxFCPXQarCQ4tetja+WSmOHb+lMmgnUyxfhTV5OBELjVhhPYyN
K0JjqSBK0zKwIQbktQqN0ZS+d+sNQZuUf1G2Y8scPhl4aug5oB36estIux0YeKfn
56/Hepg26ZemnDmm9AF6jeqnKr+/9h9MuiDa5iji6FYZY1Zor4WXcUdYtlcqBXnU
9v2gwoGVWrtKooeww8ncac+D1u/Mic4Q8CoXOyRMyrJqYa34oR5BQ2nFk17v73rB
47RMQLkg7F4jTqcTu674x1AMEa2eD7JP+xKBuzwmyWMFrFi9U408mMZPQAaaIlEa
j+0XyLjMRMA6jiYqKmtQcquB714vMFisTFmBQ3p9fIpU5jnzvcyHVDJuCcycHVwC
0okr0EOsggPhXY9zsdKoVB7656i9UuxZsmdvH5Oi4ma5Mps5c9p8iUvmzTq9xfEs
+Rl7AVZkZJ9S3YSgdLDNhc+ElXk0Z43uNA/HOBG1HEE/9Tb2VUF885w3PWMjrJi3
OBbAFgz1S0UOKeieKIxI4negzraBCfM5pxrBARo5yymbDFZFcSWFRMlQk0wCatDg
OcUDO0fat49W/hXVEx877RO+0qHeF+V4ejRSivHAZq1K5rOl8PiW9Pw5GBAn+cTQ
ZTslFcxzRrcr0rqR2S+o+Be1Z0o5a0viGbbi6RgL9eF+U7NNMbQzc4JPP9Xvh5Qs
ronvCpY1pJV2qWAEmsjbGdoGvn4B+4kj1vct2IVSaRiouuFrXb/jpft5FKfom643
0Zj7CQaXKfhdhyZVxu8tOJZd/Rfpm+xFuWrkMcz5MmsWAXzKEk4HfJha+4CM7LN0
YS5SeEsYI80eRLOTGmjr8L27eKJ8uL/CRlLFcGW2/Jp64z/MYy32s9OvQfTa35V3
W7jQORdz9eVCmLWpXhmaKhVN3tguWLfl6y1ESz5bGhGsxDnqHcG0ad87+G2taEn9
R7z0QueC4FITvxPgfUwEXV96g3awbbuqxD7W9ZAxNfNStg5DhjUCO4IJrUPSELsC
ALrHNworsn5Y5XtkBPhm2ZBX+aKFGjsASAZjFTkL/xY9Cq2Tp1GrM+V0owwOgEK2
rSGii1RqnsirW2Z3Qzq9sefPj24qzrIwZCWsD/YNNllazTy/rulGbgzbLQcatoI2
qVUMTeK8OYQw2j14VrhUWHj+llzS9xY49k2r6XLoKoh2ToC8TPLNh7IAtAbLKfDq
ceViuFHx3ujUj8hXLx8YP/dOirE2o41zq3+H3wQTL0F00j33GpdxDUDnhM2g2uqZ
R2TTBSnXIWrAZL1dSXhA/PlujKd8wx1gFt/BTSbSKZNTjhERJ3MLpUuKqzdkcjCQ
qfOJPzSOYKn5wajQ73ALTKtwd8uwp6zRdlmkp1syafQZay5FA26VsRgfiW8R3Ktk
Hcx540snZCNBkuu3fSpftBoYIewU8mOmrKKn/Y/hofIQWFJhIC+kMJsnl2tEtGbD
sSYp2wrpCOXcP/qlUc70Obk9fM+okI9fT4nfzJbvZApqBXdzD3cjlWD2F4U9Vs9R
B+mhErCPj656234yDwbPeSV1izqQlOdGUWbgeVqzAKNWjxrA7OozwW0h0tGolfDI
5byXUtkgj6vaArh7JuGMK7HAVfgpU1ZjCkHMU/z1xT0yAtzobcht2nnkOtj5BjOc
b2FXwKthgw/BbHgAnUk2viQLh7xNs0fny6pH93VJdr/ayNv1fVZemR9BekiUSMmE
txReO5U9jGJjkwuSqO0YM9KHWxDi9Ngz17nMMhRWrcz6GptPfMcA4yV1lmrj29aN
Pp5qDq14mQ/Cu1xZ9cIxbfy8JCk+wItKB+sD5bzDhtmb7SrK6nc6xZgHw3MU0MLm
7amieI5ak1gXx0lXtXt8Xe/bpJgvS2LZXFkpu5uXPnLSmTXylNcUVUd7gixbq8Ln
9JDn++nvwAeIi+jD2Y3os9oaAY/Gt+7LMQLowVib69LQO3JDL5pMBMeVyqKsulyJ
dVzLbiLDtFKsLhLwyS7LxfxWIRF8Pw4zCoKrkLikvsdMfv/JEMxOYpo1VaRHctSC
OW74L5gTKRWELSgWV18gSfkyhKKicBlz6lAI/4XIfKl4Yphrw95ftfl+q4uZMH5F
4Rttv3oEeOKsdUh4ZdZ2ErnQ2ssYyyt6dXY/SXhl2mglG769bpjw3dt/I9t/0aoF
dn3wpSbuqB1mtfyk4N2wY0EbAQZ07Q0n51twQ7p68lsfqsfMVCjRpHZJr/VC/4ss
ChuEFWWbhlAijmlgEgLH53m3k+SmX0Ie2sPfNyiZHvIcHc/vPQWeWJJiEqMpeUkU
gSLZq1KPeiL5uHXBHXOVsCisY1TnMP08bUqpECshlECqVhW/8hnbSDpmEQb/+Z5/
Ff3S4IJwYr8DQKWNOAV3aqjtUMEqfvUIiPbOVEAz1q4X5JzHX5fvbR6XqrUaMr3N
o5mQ1APXcVgv9CjUs85addX7qsyGRVftsy23N2Jp6YGi7LAwhQ0LyTaO8vDpmgzz
7VngbRDOpkp1tf2fp/SU6PCO7GYL4pm0WztHgle9zU4XkZ6lylWR+lKrppfvFRsG
aszr5zSaM+WxqplIbf2mXo9Wo9PRTbXX5q4S79OGgapsVTpjHQPwQYfV02bRBDTu
bnatyfk3O+pNZlDjzWCE0js2zJUB8hNpTPxSMi5mEMXWbDaRVaAq8WKXc/XnH13D
h2zDrlDl+5eCnaw+J3XiK0WP1B4Cr5skdaVzaO3+oT6spggkbJ1r5e0MCYMu0Qw6
u29WNm6Izci9jDJwwVoDfx1GwvDuFvm6K56YxvvcHvd6Lpijgs0hXh0DWfNqmUE4
WaXhzJXSOBzKkm4M4KMH8fPLYRbxzEPT69b4AECbCLMJstldCqY9zM5kFSmq1ysL
dJBQ9MZdrUPfdVMJR/QhHMtAAwaEvjLMQM3KgvZr3Egk0sNzEH/JejboTARN+YNg
3vE5qI6Y6cJ7y0IVk5Mm9EHut1EmbPxNer5l+rg52X37DDkn1H/wZ5KjVUKrNGU/
hn18GRFCVZ2uijdnDyFbBHxEuG7GOqOmuM96EO6TE4jVX1WC0FijcQe9HITjs4qb
4OHc7Vah8idMxXfHKa0+MiB7N2+ja8cm0lWGBnCDnDK2rpa4Vo3En74rvGpi6+0X
NS/j6nFCJv9xUUMGKNwwqN4RXGXkH32czRrowSW48WhiwMYWbfVo1UG5FqkI9OKy
vON/Xt7+R0NcyMQcPMdC2uEng3a+1mobkYeFiAjlLjNnUW09p9RTefXzanj53iTG
I1fPv+NVn13/X5tExF/A8l0UxGCGVb67G/dTkhKDEZUmlgGl/DyIwYf+kHusRvbe
k9jbFTz47fdu0Dn1o/ChioNlguY+sSBGJqYHt8fm1tdHQHBIiALkKehETj2mvzDS
9J8ENjoXz4/M9T9rHPq2ZDXsw3GUfaIYrMAEZMolfuP+gdVzN71b058w3TBfe9Js
kgsNRpVZTG+YEXd0IhQ+IUsL4bWspMwIFTjdKnjVEK1s7a4YeMl+RgjijmShoo4H
GSbAlw1usk8eEBI3vyX/QRxPyIeOWUacHDhDv7y3oqs+O/Uaakc4NdapfxpFWLgj
SV/j66UsflgBgNF2Cc1k5Q==
//pragma protect end_data_block
//pragma protect digest_block
Q4cVYM0GjsJN0E+xnXLbxT21x5U=
//pragma protect end_digest_block
//pragma protect end_protected

  class svt_ahb_checker extends svt_err_check;

  // ****************************************************************************
  // Public Data
  // ****************************************************************************

  // Signal level Checks
  //--------------------------------------------------------------
  /** 
   * Checks that HSEL is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   */
  svt_err_check_stats signal_valid_hsel_check;

  /**  
   * Checks that HADDR is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.  
   */
  svt_err_check_stats signal_valid_haddr_check;

  /**  
   * Checks that HWRITE is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   */
  svt_err_check_stats signal_valid_hwrite_check;

  /**  
   * Checks that HBSTRB is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   * Applicable for AHB_V6 extention AHB_LITE
   */
  svt_err_check_stats signal_valid_hbstrb_check;

  /**  
   * Checks that HUNALIGN is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   * Applicable for AHB_V6 extention AHB_LITE
   */
  svt_err_check_stats signal_valid_hunalign_check;
  /**  
   * Checks that HTRANS is not X or Z  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   */
  svt_err_check_stats signal_valid_htrans_check;
 
  /**  
   * Checks that HSIZE is not X or Z  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.  
   */
  svt_err_check_stats signal_valid_hsize_check;
 
  /**  
   * Checks that HBURST is not X or Z   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   */
  svt_err_check_stats signal_valid_hburst_check;
 
  /**  
   * Checks that HBUSREQ is not X or Z  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hbusreq_check;
 
 /** Checks that HWDATA is not X or Z   */
  svt_err_check_stats signal_valid_hwdata_check;

  /** Checks that HRDATA is not X or Z   */
  svt_err_check_stats signal_valid_hrdata_check;

  /**  
   * Checks that HREADY is not X or Z   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hready_check;
  
  /**  
   * Checks that HREADY_IN is not X or Z  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hready_in_check;
  
  /** Checks that HRESP is not X or Z   */
  svt_err_check_stats signal_valid_hresp_check;
 
  /**  
   * Checks that HMASTER is not X or Z. This is performed in full-AHB mode.  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hmaster_check;
 
  /**  
   * Checks that HMASTLOCK is not X or Z on slave interface. <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hmastlock_check;
 
  /**  
   * Checks that HPROT is not X or Z   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hprot_check;

  /**  
   * Checks that Extended_Memory_Type supporting HPROT[6:2] is having valid
   * values   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hprot_ex_range_check;

  /**  
   * Checks that HNONSEC is not X or Z   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hnonsec_check;

  /**  
   * Checks that HLOCK is not X or Z on master interface.  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hlock_check;
  
  /**  
   * Checks that HGRANT is not X or Z    <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hgrant_check;

  /**  
   * Checks that HREADY output signal from bus is HIGH when reset is active. <br>
   *  This is applicable for:
   *  - Master in Active and Passive modes
   *  - Slave in active and Passive modes
   *  .
   *  This check is performed when svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1.
   */
  svt_err_check_stats hready_out_from_bus_high_during_reset;
    
  /**  
   * Checks that HREADY output signal from slave is either HIGH or LOW when reset is active. <br>
   *  This is applicable for:
   *  - Slave in Passive mode
   *  .
   *  This check is performed when svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1.
   */
  svt_err_check_stats hready_out_from_slave_not_X_or_Z_during_reset;

  /**  
   * Checks that HTRANS output signal from master/bus is IDLE when reset is active. <br>
   *  This is applicable for:
   *  - Master in Passive mode
   *  - Slave in Active and Passive modes
   *  .
   *  This check is performed when svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1.
   */
  svt_err_check_stats htrans_idle_during_reset;   

  /**  
   * Checks that HRDATA/HWDATA byte lanes are selected corresponding to
   * bits HBSTRB signal which have value 1 . <br>
   *  This is applicable for:
   *  - Master in Passive mode
   *  - Slave in Active and Passive modes
   *  .
   */
  svt_err_check_stats valid_byte_lane_for_hbstrb;

  /**  
   * Checks that HUNALIGN output signal from master dosenot changes its value
   * in middle of a transfer. <br>
   *  This is applicable for:
   *  - Master in Passive mode
   *  - Slave in Active and Passive modes
   *  .
   */
  svt_err_check_stats hunalign_changed_during_transfer; 

  // Slave Checks
  //--------------------------------------------------------------
  /** Checks that RETRY responses are not received when configured for AHB Lite */
  svt_err_check_stats ahb_lite_retry_response;

  /** Checks that SPLIT responses are not received when configured for AHB Lite */
  svt_err_check_stats ahb_lite_split_response;

  /** Checks that only OKAY responses are received during wait state */
  svt_err_check_stats non_okay_response_in_wait_state;

  /** Checks that ERROR response completes in two cycles */
  svt_err_check_stats two_cycle_error_resp;

  /** Checks that XFAIL response completes in two cycles */
  svt_err_check_stats two_cycle_xfail_resp;
  
  /**  
   * Checks that HTRANS changes to IDLE during second cycle of ERROR response. <br>
   *  This is applicable for:
   *  - Master in Passive mode
   *  - Slave in Active and Passive modes
   *  . 
   */
  svt_err_check_stats htrans_not_changed_to_idle_during_error;
  
  /** Checks that SPLIT response completes in two cycles */
  svt_err_check_stats two_cycle_split_resp;
  
  /** Checks that HTRANS changes to IDLE during second cycle of SPLIT 
   * response */
  svt_err_check_stats htrans_not_changed_to_idle_during_split;
  
  /** Checks that RETRY response completes in two cycles */
  svt_err_check_stats two_cycle_retry_resp;
  
  /** Checks that HTRANS changes to IDLE during second cycle of RETRY 
   * response */
  svt_err_check_stats htrans_not_changed_to_idle_during_retry;

  /** Checks that IDLE and BUSY transfers receive zero wait cycle OKAY response */
  svt_err_check_stats zero_wait_cycle_okay;
  
  /** Checks that if invalid HSEL is asserted for selected slave. This is applicable only in mutli_hsel_enable mode */
  svt_err_check_stats invalid_hsel_assert_check;

  /** 
   * Checks that HREADY output from slave must be either HIGH or LOW when there is no data phase
   * pending. That is, checks that the slave cannot request that the address phase
   * is extended.
   * This is applicable for:
   * - Slave in Passive mode
   * .
   * 
   */
  svt_err_check_stats hready_out_from_slave_not_X_or_Z_when_data_phase_not_pending;

  /**  
   * Checks that HSPLIT is asserted for only one clock cycle. <br>
   *  This is applicable for:
   *  - Slave in Passive mode
   *  . 
   */
  svt_err_check_stats hsplit_asserted_for_one_cycle;

  /**  
   * Checks that HSPLIT is asserted for a master that has not SPLIT earlier. <br>
   *  This is applicable for:
   *  - Slave in Passive mode
   *  . 
   */
  svt_err_check_stats hsplit_asserted_for_non_split_master;

  // Master checks
  //--------------------------------------------------------------
  /** Checks that transfer type of a SINGLE burst is NSEQ */
  svt_err_check_stats trans_during_single_is_nseq;

  /** Checks that a SEQ or BUSY trans only occur during active transaction */
  svt_err_check_stats seq_or_busy_during_active_xact;

  /** Checks that htrans does not change during wait state except when
   * htrans changes from 
   * - IDLE to NSEQ during wait state for all burst types
   * - BUSY to SEQ during wait state for all burst types
   * - BUSY to NSEQ during wait state for unspecified length burst
   * - BUSY to IDLE during wait state for unspecified length burst 
   * .
   */
  svt_err_check_stats htrans_changed_during_wait_state;

  /** Checks that contol and address does not change during wait state
   * except when htrans changes from IDLE to NSEQ */
  svt_err_check_stats ctrl_or_addr_changed_during_wait_state;

  /** Checks that write data does not change during waited writes */
  svt_err_check_stats hwdata_changed_during_wait_state;

  /** Checks that burst transaction was not terminated early: 
   *  - AHB master should never terminate a burst transfer when OKAY
   *    response is received.
   *  - In case of Full-AHB mode, the master should rebuild the burst
   *    transfer in case of EBT/SPLIT/RETRY before initiating new burst.
   *  .
   */
  svt_err_check_stats burst_terminated_early_after_okay;

  /** Checks that master attempted transfer size greater than data bus width. */
  svt_err_check_stats hsize_too_big_for_data_width;

  /** Checks that burst transfer does not cross 1 KB boundary */
  svt_err_check_stats one_k_boundry_check;

  /** Checks that burst transfer does not cross configured boundary limit */
  svt_err_check_stats boundry_crossing_check;

  /** Checks for illegal address transition during burst */
  svt_err_check_stats illegal_address_transition;

  /** Checks whether control signals (other than HTRANS) changed during burst */
  svt_err_check_stats illegal_control_transition;
  
  /** Checks whether control signals(other than HTRANS) or address changed during BUSY */
  svt_err_check_stats ctrl_or_addr_changed_during_busy;

  /** Checks for IDLE changed to SEQ during wait state */
  svt_err_check_stats idle_changed_to_seq_during_wait_state;
  
  /** Checks for IDLE changed to BUSY during wait state */
  svt_err_check_stats idle_changed_to_busy_during_wait_state;
  
  /** Checks for IDLE changed to BUSY */
  svt_err_check_stats illegal_idle2busy;
  
  /** Checks for IDLE changed to SEQ */
  svt_err_check_stats illegal_idle2seq;
  
  /** Checks number of beats in a fixed length burst */
  svt_err_check_stats burst_length_exceeded;
  
  /** Checks that a master started burst with SEQ or BUSY instead of NSEQ. */
  svt_err_check_stats seq_or_busy_before_nseq_during_xfer;

  /** 
   * Checks that for non existent memory location default slave should provide
   * ERROR response for NSEQ/SEQ transfers. 
   * This is applicable for:
   * - Master in Active and Passive mode
   * .
   */
  svt_err_check_stats illegal_default_slave_resp_to_nseq_seq;  

  /** 
   * Checks that master loses the bus once it gets the split response
   * from the slave. 
   * This is applicable for:
   * - Master in Active and Passive mode
   * .
   */  
  svt_err_check_stats illegal_hgrant_on_split_resp;  

  /** 
   * Checks that master asserted hlock in the middle of a
   * non-locked transaction. 
   * This is applicable for:
   * - Master in Passive mode
   * .
   */  
  svt_err_check_stats hlock_asserted_during_non_locked_xact;

  /** 
   * Checks that master drives HTRANS to IDLE or NSEQ when it
   * does not have access to the bus. 
   * This is applicable for:
   * - Master in Passive mode
   * .
   */  
  svt_err_check_stats htrans_not_idle_or_nseq_during_no_grant;

  //-------------------------------------------------------------
  // START OF PERFORMANCE CHECKS
  /**
    * Checks that the latency of a write transaction is not greater than the
    * configured max value
    */
  svt_err_check_stats perf_max_write_xact_latency;
  
  /**
    * Checks that the latency of a write transaction is not lesser than the
    * configured min value
    */
  svt_err_check_stats perf_min_write_xact_latency;
  
  /**
    * Checks that the average latency of write transactions in a given interval
    * is not more than the configured max value
    */
  svt_err_check_stats perf_avg_max_write_xact_latency;
  
  /**
    * Checks that the average latency of write transactions in a given interval
    * is not less than the configured min value
    */
  svt_err_check_stats perf_avg_min_write_xact_latency;
  
  /**
    * Checks that the latency of a read transaction is not greater than the
    * configured max value
    */
  svt_err_check_stats perf_max_read_xact_latency;
  
  /**
    * Checks that the latency of a read transaction is not lesser than the
    * configured min value
    */
  svt_err_check_stats perf_min_read_xact_latency;
  
  /**
    * Checks that the average latency of read transactions in a given interval
    * is not more than the configured max value
    */
  svt_err_check_stats perf_avg_max_read_xact_latency;
  
  /**
    * Checks that the average latency of read transactions in a given interval
    * is not less than the configured min value
    */
  svt_err_check_stats perf_avg_min_read_xact_latency;
  
  /**
    * Checks that the throughput of read transactions in a given interval is
    * not more that the configured max value
    */
  svt_err_check_stats perf_max_read_throughput;
  
  /**
    * Checks that the throughput of read transactions in a given interval is
    * not less that the configured min value
    */
  svt_err_check_stats perf_min_read_throughput;

  /**
  * Checks that the throughput of write transactions in a given interval is
  * not more that the configured max value
  */
  svt_err_check_stats perf_max_write_throughput;


  
  /**
    * Checks that the throughput of write transactions in a given interval is
    * not less that the configured min value
    */
  svt_err_check_stats perf_min_write_throughput;
  
  // END OF PERFORMANCE CHECKS
  //-------------------------------------------------------------

  
  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

/** @cond PRIVATE */
  /** Reference to the system configuration */
  local svt_ahb_system_configuration sys_cfg;
  
  /** Reference to the master configuration */
  local svt_ahb_master_configuration master_cfg;
  
  /** Reference to the slave configuration */
  local svt_ahb_slave_configuration slave_cfg;

  /** Identifies from agent cfg whether a master agent */
  local bit is_master = 0;
  
  /** Identifies from agent cfg whether a slave agent */
  local bit is_slave = 0;
  
  /** Instance name */
  local string inst_name;

  /** String used in macros */
  local string macro_str = "";
/** @endcond */

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param name Checker name
   * 
   * @param cfg Required argument used to set (copy data into) cfg
   * 
   * @param log VMM log instance used for messaging
   */
  extern function new (string name, svt_ahb_configuration cfg, vmm_log log = null);
`else
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param name Checker name
   * 
   * @param cfg Required argument used to set (copy data into) cfg
   * 
   * @param reporter Report object used for messaging
   */
  extern function new (string name, svt_ahb_configuration cfg, `SVT_XVM(report_object) reporter = null);
`endif

  /**
   * Execute signal level checks on the read path signals (driven by the slave)
   */
  extern function void perform_read_signal_level_checks(
    bit                                    checks_enabled,
    ref logic[`SVT_AHB_MAX_DATA_WIDTH-1:0] observed_hrdata,
    ref logic                              observed_hready,
    ref logic[(`SVT_AHB_HRESP_PORT_WIDTH-1):0]                         observed_hresp, 
    output bit is_hrdata_valid,
    output bit is_hready_valid,
    output bit is_hresp_valid
  );
     
  /**
   * Execute signal level checks on the write path signals (driven by the master)
   */
  extern function void perform_write_signal_level_checks(
    bit                                      checks_enabled,
    ref logic[`SVT_AHB_MAX_ADDR_WIDTH-1:0]   observed_haddr,
    `ifdef SVT_AHB_V6_ENABLE
    ref logic[`SVT_AHB_HBSTRB_PORT_WIDTH-1 :0] observed_hbstrb,
    ref logic                                observed_hunalign,
    `endif
    ref logic                                observed_hwrite,
    ref logic[1:0]                           observed_htrans,
    ref logic[2:0]                           observed_hsize,
    ref logic[2:0]                           observed_hburst,
    ref logic[`SVT_AHB_MAX_DATA_WIDTH-1:0]   observed_hwdata,
    ref logic[`SVT_AHB_HPROT_PORT_WIDTH-1:0] observed_hprot,
    ref logic                                observed_hnonsec,
    output bit is_haddr_valid,
    `ifdef SVT_AHB_V6_ENABLE
    output bit is_hbstrb_valid,
    output bit is_hunalign_valid,
    `endif
    output bit is_hwrite_valid,
    output bit is_htrans_valid,
    output bit is_hsize_valid,
    output bit is_hburst_valid,
    output bit is_hwdata_valid,
    output bit is_hprot_valid,
    output bit is_hprot_ex_range_valid,
    output bit is_hnonsec_valid
  );

  /**
   * Execute signal level checks on the write path signals (driven by the arbiter)
   */
  extern function void perform_slave_write_signal_level_checks(
    bit            checks_enabled,
    ref logic[(`SVT_AHB_MAX_HSEL_WIDTH-1):0]     observed_hsel,
    ref logic[(`SVT_AHB_HMASTER_PORT_WIDTH-1):0] observed_hmaster,
    ref logic[1:0]                           observed_htrans,
    ref logic      observed_hmastlock,
    ref logic      observed_hready_in,
    output bit     is_hsel_valid,
    output bit     is_hmaster_valid,
    output bit     is_hmastlock_valid,
    output bit     is_hready_in_valid 
  );

  /**
   * Execute signal level checks on the write path signals (driven by the master)
   */
  extern function void perform_master_write_signal_level_checks(
    bit        checks_enabled,
    ref logic  observed_hlock,
    ref logic  observed_hbusreq,
    output bit is_hlock_valid,
    output bit is_hbusreq_valid
  );

endclass

//----------------------------------------------------------------

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
mv3EjS9Gl7pglQXmn0v/3h0yKqISNYC/oR5lL3I2IL03PpqIApltMELhkyKips5W
Kld9X+zRjedjcA8MPFcliRpzHaYcPag3Lob0YfWLv1zer5QTQlWJoHVvmHxAyvZ7
zHGKSrpII5ogQVKjQ4nUa+ktu68awaEUuOu2Ttghh78cUb15laqXrw==
//pragma protect end_key_block
//pragma protect digest_block
HBKEXYSlBJzk+eJq2fjTGPoAHFQ=
//pragma protect end_digest_block
//pragma protect data_block
HReVXAe9O5BIH7YoEAOZEacD5hcTuQrBkWAdVC11+QYNIpl+Oany1KyoARUhNVhi
UUJzNsVo29xBkebHA+kLaZyk26HtN1P8WrDGxfH4J6VI/M3xUKaxen/9nXUR0PlU
c7BEtGkoag96kBKhGG9mDBpRODX21gINN7eZEctCRoqP22v0V+Eg6TQHSXxFCGXj
8hV/BqbpIjWZseF4RvDpPSUxQwgA6W7kB0KopyVnd9F32/ZpPo28DHrSwiNxzeV1
hXvTQQJZKcqdNQNUjXV0g77+pGUDc0fJNe/QzbElmdGKEbYqJbufr3yvcPjp5lsN
wU81tF1gbE+qYyexbPwo83Pq43uOX0wZCl0MX4VizbJaS5YVcFyU/6AISoy0PfdQ
ZdjjUN9djcmc3xiZd8jZ0eJu8oFjpcVTtE+JhjrEXGsTY/ASVQaRby9VldegLQwN
31nbxGR5Dxbmb0xYASULh5KJoKFp/DUkV7S0FEFjI+Rw5cSDK3ysoLSCYtVz1Fky
oSEV/D82hFs38PQjd2scfNxxPUvF/XGqNWV77ZwbVEp/RYRZ8UACNu8Swv1/yvbB
VjnDShbt9HVAoPLUNiLmnZ7MbrYUbpzJhvt0GOuerxBNGfFKj7mHfPF2kZEA9CDQ
VRsCsyaJQmX5MHHcAe9Jvx3l3kKhoMwoVPfEuM9PyRNk+6E6jkzSUca6lvwq82Gi
726nUZO/POo0GS1GNbg+abLpH0bEu/v7Y2XR9rwh7u/opWi4VUZ9uDYagQu4xTF6
93fYuz49iogPgBYsH2ixBpxH+mb/eqU/rc64denN4EMQIV551AIL5dKqsYFdgLpw
gWdkC3C7sENGJOwvUbtVMluggIU24qHf2n3iV50oCKZ9xRUL5RS4HRrXZvLy+oPu
xV7U8w5+1EdxbONy8gb77P9JEDX4UFxTDCSjDbpZnS3/dkER4kJ9JeoBgrnpG/pP
sVdf1HcwutWuSeFpN4PhkZw9P5tT+joaJe91N07ZTmqjM6EXR/2tyd5c3Rf834Me
ha7fApDYUt2f2ragokwW+Gwo5nBDzF4qVebuJI/n/2ekwRt21clZl45gbNd2WOFP
btJSrTKe6LCx3R+8XmCqHSSqzeoDPz9kCMwoSXWZRtNl3/ExUgA80qMQjbusubZ1
d3LnA7r4NsopH85vLecvzMPqNYnOGnLMKid7aFEQ+M6PMpdURWxsqIwnRQDKX4g2
VT1kt1VsJhf1w4TAMk8ATnErfcIk8ghWdOGCOcN6+Y63oJwUYLxkAdpW+KTD9laZ
hvd+ZczsJNAM6VYglYsdtFnMKlXhA/ysCdYIU3H48LvDupbByuG7c3ubDcTFM3Mu
0LSvC3r9xAYiaJZs7fJaO/H2UqJ5sHmSdpKycZ+pXC8DWnBE1h1o9SkNOec38DCP
cpfl9JfBn7CEWAoE/6lg6uihMkKktfrMMEKXPKV4bRPS6Sk6evrQijIMDztTXzYE
peyJiihy9p7jdWm6KrCwV8HIexQDlpv/mYOeG8LJVItEXi+Jk7clnw+RFdMZCFOF
JB2z053KzjM+uZnGr9f/k48BcZyFLi8XvsG0UUtrO8xWXVk7JPh4PkyIP9zTegsx
3zY/I6P9huUB0MhOJGWynEdljyLT7BJfVjN0bMzFalqJXVBnrVGiq2nuOZNB0ZYc
2KeERPt3n8GBeUz6nTnEacJZyMX+K0MMknmR4DkTZ6XnLRYZTGc+ay2Kv7gVPQOZ
pQ2eZMlpFmyBWbnbBjDZTDi0T2HOvlIFP/eLXUNtGNdlMY8BC13lRdFLy2o0pqIf
mHQ8g9Q2thEjBRrnB/4B2Txluiew2L1Yes3WJTkr2p1Tn+cPW77oMpSJip6XoeGQ
ZWbikD8YuslP/LDMnDJ3n4RF4oGfDFeGG+ve2A3NqVXmKwJv2f0a9KlVH6q4Ycn/
T1INLiZ6NOx9b9D0+08L/Ni0Gdef7tG2n3FMbAhmCsGsnsIrHvbYL0cmiRBRgMj8
Gw2Ilh4KYecHLlmh5ZUcAb6OtK7EjEnvE53L/9xEDE9tH9WUOe8mysT5Ez445cbd
h1EoZwNTowBaTBrxio4Eqawr8VFyRCe4w7hQUQGEvPR0TdV/0OnyZWutJVKEtuBu
+pary3tqYTp9qNC+JP65Dgk3fr/SCD3SjugIq0ChKpKC7BhkE+VJSk7JDMHlTfMi
lFd3i488xxoCo2O2xeeoIEyKEGlq2XiOpG17YyS1Ilt9TR6sdFVZsLsiL2cFbPDi
X5NymnjNPPnk7hsqRPhPH2hRdPXooGx19b53DDs05MJeEboAVfIDuHRRBLWD1JRV
3mb37byNcwxf7mJe6Q9OVmC1S2qAzIKHcc7Dka5MjJ1uRMhI5T6nEgW1QCjwKOHR
rzVQEJdPoEEfuVTfDK9lVNysJyi68lglWu0eQ2k1H81AwTyIEpF32XoztvLt+7wW
5VaQxYRDiFPbHxiMqU3XqjG1yfOcp6o2ChN/QnYtBfjiZUrcqkmJ93Xvm3BlR64d
ljY7CuyU0UASWq4AFPcjnIuYoxuYwsx8dWSSq50nFeUsyAZbs9qpzMXzxiDzG4yv
AWonQFVU9a2i28cem7WbzflImI9I9gLP/p155rqFJRUvKUzeo0xjr0oMdE+vywDl
Go/vYPXvx+uymbDcNgh4h/f4L6BCL6PeqQy9TyvAFesvQI2TzoWgDO9mlKCE329n
pPaRliGRhzqdO0ND5/ubY4lWGcP0Bt9y+3hjyEJDzfOhEl1osTNHd0JTGer7nY2z
jmUJh0OekU+XjxZsgm96h2d9EoMAsdLls+UuY30OLeTa9LtLdmAGBK1GNAqt0v7X
+q/TTHGqn/Kte1uPbJ4d+7CQwn99Z69y5cjcc1LOxLwko8+jFUxrRk2h98Mu+CjO
0Up5VXUgk2mgySnU+E5ABV21fqKqrRIYpcmbsWaF1WEfm2i4XIhO/IqnynA3OB50
YZM7KNzSX8OOe/0/P8r2SSsGv6sIDZd8drvG2PwOSHpF8uVwqIhiT0vz6F4xDu6J
lvkFujS15/gOn3lQgcFesMksb34KTffO2LJe/OwHv2vP0lE4E2I2mhUzYpoU3k9q
mUfJm6MMvfbQ5txLFZ+Qo/sBcqg5u9w3xCte8765MwWItN1CHsfQvZ9R46VtkDrR
Du1w69mS++lg2lgKOW6JcQ3CC/pQqEbX7o9MCZJK1vqxUq6EyPeIugCqYiadtVvl
QgMSQJFVrKfLP5IRQCY9/sT9rOsCFwgbgvdVNXoRO9+ju6/cduoR2T4V5QBhcqFf
hlFC+mA2hPxYO1o+8qC55ATCs5NyHo5ZGGtcnbRY8LKrHHy0wVRleRYyPUkdHAuV
71t2CCaS8tLewv0xLmEwFVvr4pAGAoTPTVlrVF5qAAFLwn1dnUNh9bCl4IP6/xpL
7+7asZELquycT6ujuH6R3rNZSjaLTPJYBzylWRea8v9MemW+6E0+kLvjzd7YIj9c
WPNASlJltmwNCEcNlSvUWXiiNisHXXxBSs3QIp4seb/B0gJLA9SciD8Q9pPUMcBL
IVKA4VBgA93g5uQCE5c7cNDjQaPoUC64VyC5kckOASkHwIsK/rEnUMJSyoq+ZPli
hKbnRKBfFs4FEhU7I/r0JfaMOocG4SrjvpEpwhSEAxDVbkhHBU08WYoywEibkgAC
sdxY+Q4aK3hmcBo/MOODCjX0p3sQAAYWOR8boBfTSTXGjXG5dmwPy/8UIPSisftw
6Dl8PH2m6Izjw8l4QZeowqmJ8nfIrW+P6mpIDuo67GqahpSFse8z9HgUTaDywWrs
QnlpUkW7N8i6mXCeg3knr04AZiY24K0TLg9voIbd+fNjIJI+ZoedzHT/lXOiaOMo
Sh6JAGPV5pwCWDbMDKAVGB3XjQ/6E08Y4Qfvyl+WbXqsa7JhAnebWdiVqq/T/m0c
XJdAW1ZcDDZhkfngWl95L7b+WWzyk1gD+X9XpUYEJUvdgdyZRAR/5ZiqKOWf3vz9
T6w12mWwj3YMNDhFrXD5Gm102gsUc/fRkROA/9WZfKmy6NhdGUkW1veGHoCKqCrT
rtQ5bQfphXhOgXhuwyvwHNQapgbVdcZ0Mb1YhSUUpJu3MbUAFPNP5YmEoFdA2FKG
wW4RKH1Gqd6fPdt12kBQHep+vtme7U5krX5ZwCDzoo58qTxPQZf8C7/q8xST0zfB
gaDfbb+iYK6rUCVFBAzI6QKTHFrW7cr8VMTiuGq380hqRbICGYuzPMYTh/zsJtsZ
qJx1BquxiaOh3TMcpAx5D4VuQaYyzqV8V9umBn33pMjVuivPIGAr2p+ORfoSXjGE
tDKKdBaEf07ZGwIc65e0B/xZJOD9ZUJ05KMvadjD5DKnFRgAZXEBQC8BGERctzAo
nfsSORLZvQUkTbmA+Uf7pngX5LbgmVHt/JrkYRadCwyFMEFc8suE1VbqYfdGTedJ
mqSdldxyiZHCxGn48onFhnGjDn41WP6PlDTZeAuOoc8W8DFfnhOwcqoLi4ZXVSmq
+wGkFmvDfB/kyDWqHXGjv19KvjH75EINUaHbMwvRr8D1NVqRcIAS7fQT+rm/M1wj
WOvhqOnqx740iX7CwGu64i08oPR7H3uGFoS297bfkDlYeF1Ax4Y+ghR9B9Go/2aW
znvZWIVMbZ1Rb/Yy+iT0MrZMzhWnEqEg8ZYkat2rG+i0BOxmpEmsmNPitDsjpgQV
vDpe9afwhxgqqyJu8Bw/bIMK1boz0PgLWJTsvlKPpCw/jVSSM13IASxxY/nahzns
IsDeDT9rAg89YNlNu4ajkZeOZfbe2yO65pV+EuWvF5OoMPKGd3X4uKwIgsKgjvgc
222MjR/ZT2/BQBNeHtayxMM3aBonDOpEXwqpnfnIXrt4a1AzDihUV/qIVf9jXT+Q
sk9oR/bRFKGKzu8lbc7bGFYNPummVN2GRldxh8XZVkRzgiedRQZOStgKt/ZZT0aN
jh6qifBmhDFkJYgRzNYX9BYlE9Qd9S0lqQIQzQ+4yfvxF96WM3smwiGDN9jeYqUK
k2M6uymzH6BWoyabeZaGoAzT0w06ZXgSn3m9vOp2YVLsaQb3/AJRO6xFqzhtcY9q
2kLWuPw+rmUxu98W/6RMvnrmLq6vYr3KF2CZ5Ma3CKdgg6wATE8zRIecdtR64802
ahaBHmSPCI5ZKqO95YhK/P8tN5FX9IMDBQlkMnj5z85JatedIYcMY/dGgbglBgAv
tfp7nIadMzRLzkDL8YWbPYBVu7CPQBolyLWhFmXnoyEU4SrS7ohYR4eZqno354fl
UZqksF9VrWIcWocGcO61oZv0qT0D1gsNXQb5EMGNC33II+8Smp32c2uEZsFU7M9b
zT4CGaAm1aQ4WLuf5J4D04jxoBJZc9Xiy/QLPRD00wYFW5ilAKmmVl7iD1qwDDR4
XPEaIgfFYadp6/jljXRRpAdcjdzuPMmSKd7MmZWQxUOQW0yP44qwUXjNfUGLCVDR
T87WFNz3DV7JFTXg63NP3G4/cqnRyJTaK65hfnY0lblLRkmM+PsvzLaw7WOx4SyS
++pMdyFwBPEQJREKOoq8pI/usb/3dTiukCbp2gSXUPYVQ3GD5Hi2IGpp8xRwQU/E
TibjcEU/XD2J4y5JRikqYir1SSO/FB69DYNrcF0YpUUcJfTR7rsqKd2if09rcS5D
x0ZJvyPrp4LUc/639bSd/MUIq2H/Re+NuOpDP+p81BDpAoIL1npvJxiSFXJj8O/N
7YL5SQQtyJheHHwKCzi2mVzaHktb0tZqLCZioqgyHQKncjniDHpc9ijJIJW9S0aU
f19C00/3d5GVG9Pat2EVgxk1HmJGjOoh2LqsYqxzZ/6JPsh0P2Oxgb22Qesw6zvI
Y5RUUUC8p3tzETs+GPCsRF6yht9UVrefbrBZ2ayLogIMNWwtYJMP/trVGtdpqhed
SOLuaZ9E8mJUGbjLP0AX9pXYYLDOdJ6havuotUIl7QDi2A5T36sSfVK7Pm2FgXce
MMaX3pxF8VaqwyVYpeaVPCNFrh8DOZw1KYvWIa0T2BTPw5EnsZBE43gC3e1/3FWF
zvNkVh8yPpFNm1VLCrv5SCrfXSrnStuOIS8c1LFeJLXrApL/8w4cFt3gXxsNp3K2
NZSW54lmg2v9SAJS+Pn4XPLkSwjrk++IOfkzLt6RWS0y9CrW0F0j4PMNqV97Qj3K
dQxU4wj7nCfwnd8nh/7KORtwL03IxfPb/A/H7Ja4zF7Lh31KO/ON5x7bMPcuZnDg
UaY8fUziz9Yyu6pddeBR6Miywby9kNxWLAWGp2m4D4w2yU31rvSfqBogXdzfMumu
QsSHHclzkt8EXhJ9h1OrLAds+y4oiX3n0QhG1Ivef6yj76SkU3ITBRIl9HbVFP/J
d+32l1fDcQl+MNmdy3A48Csm8kDseYTmxFKzIGQ6U6Opq1moZ9m099SQ4a5lWqfG
KN6dcK/mgFwZapPpLVSmE733EmEewrz8WWn8bp3VWlSPpm/0LeGXXPLAL16GtX66
7qDfo5Ac3Y4bNxp77KcFv95B1qxBCDtNNiD8mubiqZGo8XcELRsIQmOlsc3uTXfI
PkmlWdCkzyRj5j6e7YUfyxNjZXTInE9xUrweEJmg/47aqBFUXzsvE2lFFnJ72EcT
sMtBXSJa0L7en7l/KlH7ZkHSFaLLg0F+i4xjzXFO4OxY9B/9y3f9aC9Hbd+Nl6mt
HOrk8U5/r3N+9au7WUOfoScPqOOy5oIjd6SXq0Xo4s+eoAY39W9+lfbA54PsQaD9
gPSuWa93kljyo82aQRUc5dZy2dgm0mFewIe8RIqf5G/lyeh0d8uRl5eTCQwz+rMP
CgsQoBNrz/ix1Rcst3LZhk6OFhWjKMUGmk3ixc7u1sKs72w5RoUeGdfzlFP4Yu7X
kJVgt9QpWsTdwemgGCoEGRv7cTkjY8rldZERbPvBABTnlwSwrbEBG1QzzUHUKXzP
J46DQoDI/jJNFih7NM4FA4M/5YfjqC5l8cvkWBUICBKHbCF4kcwH8EV6OWmEuj95
docb3DLsZ0vsmDpph/jlXc05SM96MJy7oKB6/M9r0mdjxE3hMO1JxNs2wFwBWKme
QEL78uBi2i2tytwTKXtzQz4OShHWnrb1c2YfpB5B9jPdLSg35aOXkkj6yeIpdfb6
AX3RJG8LIRXYpVLBzSsb1QJv0/O47ymGUotTbAU6CQwSaNf1g16jS6LqDC1VGIUV
oFxZsqCpgfRwzdSRbq4pJ1Uy5kb5oNMX/iD8pvH+wVGb+pV19a7370DonW9r4RXa
I7mNfPAuFmncmx6/ahlfJYsMA67pPRFrcdAtRhsGxOkzPKj7tiwfiyfT0OyfN3k6
wO0/X7aU/eYyYixBY5psnAnYw2XPLXh128nfyFVOsG/D9Ry/UoqKvFBdNAyeHBjf
83/cxmZ2/LnyZj8F9GfQIvGCYXvCntIWmlHzLsiz6+U16U3pa8zaqB+WhQ3j6PrJ
jpJFO/U+q44FUs0iTtrL3vnHlT/kBt7eQYu4uAxh8Sfz0PSlbdhIOhmdC0kvphJf
uaLvjLJ5W2mjKReB3kIXT6hH1zHaLxrq8TPn04MhSU4dFIf6lDuKzNPxQwKj6PNJ
sZjO9L73RnM3iv4apiiRcZH5mWykYCWo5QJHvNNfHJnefrZKz9N3nJC5OD306evZ
y7IWNEA8tCEUg/nl9XbJSCQY6EWKEP6C4cHgYWxXIp3qMyo/dUopm9bv7YZfV9ND
l/yhz4qpnw6r9BiLHK36tikILCtUiTgAt3RZBLCfTzdAoEDr40wYbgOfo6ffmm2K
X2GbdMa0ZLjdsqyvuUsYXMoYV8ifL9WfXIJF4M5ww966F2LT4kUcSnk3vBVcPCQP
eyI2aY1j0MsF7w7Mv0X4qe+G/xcULmSEddYKxItLrB60j+hU2OdVs8DgcslLsIaf
Tdv80nrFZ2BcA40KQ5lc+GHg8dAGnFhH8Sc5Ira+GH4gCqFhTc2YSmUpYoCVdSIC
DaGMlyDfQwoyjHPMhzGfQ0CR5hOOZtPdjcYno0eGxcasV47wqHYXx7jJkqOI3Vz5
vx12vc+nXbuesrvyHoa/e75lQ+2gd59yegqqKt3wwD3d//M7ZrALrZy8/HlrSndZ
JBvp5Wm2I6vWHjYhzNZ04uDKlvW9ptIC3wKHgDPXMVY/TRFCpRE4PxmkULi2Hf/9
JZ2THBm39e0lKnLRUpLDgwpmbeRoxkte36dfl5/YgbPgn/dx/Vz2dc23rRYyd8r/
WJMQ7qoV0UQ5id3lnqom11gKN0BpOqvVmG0u1qyxM1ctpjrr/walrEP/t/WyqvRp
kXgm8g4NoW84YF04+z3+YutqnZBily6jPFH0lMFks30yKekucBuAs2znDloGlpck
jvT2CMSjPiz3s751qtF2qW1d/JBPEQJVSXjPE6jTJ4KIaLo+Z2P2Tu36RYZfWYzz
7jPfKgp8eeW1B8E7PWPpK6sce8eRKktbHuMstnZtA1eZxufIjZiLZu3MCDKH7vT0
4gbU72FTvXtM+6AQQbHUM9VBfscOy0vHwQ4xasiRtpejwT3H1LzrLAv0ptawZdLq
XNdoZUgSWKzhDlHEBfsst5xIDXuhSr3o3zCjDKYMC9nxoyviZx5iIA1yCnFXnpMw
Rm3TbzYgLWqR9m+XeMd5faGKULDruQdrfFQ+NLGhMr+mzopGPU2srqAwJVhZqUTh
epfQKXIBkeWWNpkhNKu9HO5WPBPo2LdVFlAQHJpjX1m5VsRjoDqzc6LRrzIeN6oI
X6VgLHBEEzcmELIslt13pa2dHHjy8RolkRz1zp5+91Uje9MFQDqDgl/5xqqn+00m
LQ2/d3fgOdLRxCQyvcm72Zcw5un1QPvGsufUoKjWH2HzVYK+1mhZQX9WsDmACi/i
DlcN5eu7eE6pLZwKBLw1EGtEv0P8q7YupLREN3Tg9UzELmEIpJGrSmcSLm9v428Z
NNZwlMd8UG7QBXbPe6lMUlp49T0JRF3i8hQUctfJcTpqitHVQeY4xD/sgrAFVdS3
GNmbKTwTZUXyx9qK/goEoRVYa54o2uJ4WnLF+eM0PeWURxOycPHG8gWqd1D9/h2t
DZG5MlkKCVCFAdm1Lg5zCpc5+idyfVnXQEmImUcz3LYvAiD6QcAlKzDibyDR1FnI
OBtXDkxtdLo6IXh+beXaEKJhpOtBKJCnDOB+4nVyqfoCL809wB/pocsXa5Hj/osb
GSK6NQFzCMA+tFQ8jHDhTTKJMvUc3KUfC/2f5EUXnie8tBXEr0am2TXSIk+5sYxh
MjAlPBWrdiddtg1jvCEAyXHiLLLV6gAVyvSjH9f+b+qVqS2aeiT0G9mvpgj0ETi4
X2L5J0YvS8sSTocWOuu3gAoQdFKi51MV5xhlG0HIHB0KcRmDWzTaRSHlAp+0h0+9
SplWxqL6MaY6MWabauGBuxkHbTYvdWZhamPiXlLGmQoV0oUMTNMXAAi7F8zjp9/G
ZlSPz7vrv/jTJhDVbEcVyo7wa8OEiXZ98aKipHgfn5/bjlSQ/xGbrfU9/Vn/iOJ2
C/U3KPOG1sKNC3rzD251TMCVGpMGK7DprYaxEZuImvGNeeGhrVxnWQ/YO90bmkjs
K56B2CuxZy9ZoioaPzMSR9elzVjXtWliV9c9V7nMADrK7ygXDTTomf+cZJ6FrtK+
GWJWWi0CYgYKNKDVnotMXRKvOz/Ty6p6c9iAQ6xZ5X5advs4/rGrvITqINp0YBmG
rtC6mSyslKIG3xMQWzbzbgJbAK8/ac9+ijHcDY4+SyqevsodXJVZ/NgvDeNYELBG
8wOzpIC65NNpWDO1x/RyBqJCQDRbaHJcwBJ3jGRQuBZKpF0px6lTyrVFGw7L6P4q
qPFXp40eKfPZ7wWT7d35U7lOU9dz3RCH0tP5aycvuvA4iT5ruTGeJqFzLl0m+OPZ
ya0NrW0biTrzsR4J3XefpOknbuzJNzp//Mnfh1ktJIycv+3Tz4HgVbuMBWZakawS
DqE5br6dEvHfJlzitXcMAuRyLuRsk4KJUaVCO3vcX8cgxtSOhhF3hzrAQ2ByuaiV
wWpuamCSrsiNjnZokGebe+9BIQPTu6ar5/rZzMBaAvkoKZoXgGHMDHiQJqpipHN/
RWQS1PKFEzekD/WUHwnZpBgBaz6RJIFWLbn8PKzrwzApsCEX0XrFeo3St1/A8BCI
aCPENjlfMiYSziKPKyjW74WFJO1oxoDKQOHst/ggnpIGRM4vsQGZ/qKdmNdArwxy
ejfFaj3T84M3kxHJUGuCxSwO9URYr4tU6fAlD+3ckBnG48FXxpJGKGiCp+5yfkjx
m1kbD1HxGol/E1WRCrGrB7VWcruOlfaos8iTb8ROnPhbQzSGSzZf7pHyIb8DXCoi
EygJQr51iFE/RDdFociAjKuJ3PDBSBPdYo+W7zwJJmXiPjPGxKFddHep6Sh4XePQ
35TvJ1gZXlRc7woy6jvJZ7Ox/XHddsIdvQSZRpEEVYzILPXywB25lbdnH881rHJg
QIkKHrWwEkmZzHh7yyDcQgfpovOWyFhhsRPk7SCdRK03qhoivvteWhRX6rYV/Muo
MvLgHhp1LkJ1DRHhsL9lJqxyvvT8gi1Nsq03Qb0fyqFujY0QuKIK2xlVQcIolh+P
+0XL9kYFBzfSR2E42mb/rgm2sKNuILYVe6BnIc52NYvYLcoWiSuRdNpPXw71rQUl
8PRVU5z49r5aYDp9ERII0dkcMiFdZK8MbGr5OTjYTnxeqXDwKrNtEIumDQ0+tBj/
IpMzVpjZAoabWoqBtyMCuHbOFqSH5++hx6IRJaSREdCvAobDOBfiImrfor6AfzS/
/EeCMhJ6EX6NdyYBt9ZNIbKIlwAvyTNE35DUiHbmZwA2tNdSRseHrKWe5/qTGUNW
X6azCUol0lb/2tjg56llfY5m9yoN2ZmPl3L50WKHNvdY2+SloA3TL2lB1YrHya4e
0rmTgNNLfKaCtNu+j5znlHLLv2pwhCfhZOENu7OJu14iKlPZAbBAs6fINZXC/Tez
b3MV/mrK/ZL22Dg+mtcRvrsGSWjcOGvPCYkmj6Shd7HKPHZXCXVzokhg0DZa8V3e
y7qAmywfDcTywT/pwzQ0o8j5Ld8eMWzz/gwzZlC92P8HZryCXQM/BKlVHxmzQHhu
YgbgvHpX66GiB9jioS5m5SplsRrXT0Cw5TFu8hn8KmrhLJM+Hnm5OzQnwnsFCS0o
hLxazPxX8gKvpwpfKHbE8EZNs+EgD0nu7ak8QJSbxNCY2RJzUakpXeKq68jXxfco
4mbSY32RLHLif3iqf4pAcWqmPJXlDC8W9O9AdXSE18F7hgw39bN+obLNMyi8Q43f
43cRqK3mK+4impTgoGL5+HunEt8i3EJmzzXymE8II0JBmga4uIyIrtL0xws7P8Ip
ukjoBIGlBDgaZQbPtZ1OBdShZ6yvKlly8LBBBBMT0Q+xk8cmjDbNtYe1gWiQDTXX
xEMWdDrfegZLnXfD0+90O2QQdvddgQQ+2fsfpqHYfJ/dJqyHDlPooWzVhrycbMvK
MhU9rSBxTnQQcuPt7ZOdJ5cqoQCkJ3qmUdhT+HmiCbXaPz6UdJzMIU69VhYmwawy
fihM7yFyHpiOgyAmkpWSG29aNmoVmQPis69mQ+WdReVP6U6SdDuzMaoeXQobXCkB
xpqdjOqdBKTIw2hY9Sr6HBMkMlbWVtod1x8Qbl7JBGLfjRhw2dEGMBgKaXWQvXZD
jHbWPA8Jtm36StwbXKkBzg8A6EgaTyRSydijxDQ9r+S3bS+auAbYDHymNm3ujlLM
VYhIaUoIMo7RZf5fFrcFGuvdXbRTCPCcJIJ9KMzViw0Q2PI9KR5O92F6IqWRYn1+
ykbMumlbZxGqAbnpvaao6f2iFez9S7g1ZFtLKndcLaJgeCka2l7sxh6Ch3seq2G8
jJEonEfN4IN6yvrALPthDvzgcdhiSgXEMVElEJfW6EFjVDSrHp6VNRvAYpQJuADK
53nTOOcJVXrBR5zrwgtHEOXLdsyWGuI3IExdy96+ZiZPfu8JpOC6whlKRCUZVyGY
llIGt7AeqRDjWvJwN2XbjNzsemJPakkiwAzy+BaKw0ffTJejJz/JhbQ9zSr+uMNP
HeCSYYsISn3htZMgGwHAL7NRfnAp97vDHTNhTnhI1+syJak5/UPYnirLdQ5zD4tq
3v4X0aHDkhR0aZChRIZQxos4VukSV2rZ7XiX7AbPrRr5pt5j2Ol/fqvwDnZFp+tR
3aGn31vglEk70n+MWQhKDV0g2piC4xe6avUkJAc/kh2+WZnM2I4YO4eiyv2ZS8h2
m2HEAXclTYkNGxVtSuXoSVlK2sFktyyuhswNq8/0QZTWoexo7RdewlYTB9xIeZ5O
3ZB4TsfR4EpdaTpNzPh5CgWTBv785flVQFLVIQyg9hk5tzmNg6l7ErmOMdixZO9d
otnjBBuHWn8GZZV5SQjrACTjV3YOaA8phiLKtP2cOIleIZiaQ7Qd8OXY/YGFkcRh
RPxECGY37GPjTBYEj7HmFqzu8fDlEqMWBu3hM464KWqdcmMmCZV1L8JwRQ3pILGq
mBiGkjiyKpSltYhXxD4KQb+jJuuyQvG/6HIawzewwL0yDhv3w2k9zOgJozvoYjhm
Kdvxclu7BXvmCSz/dito1Eqr6VlSu11mOv0YWWrFS+I5TTVnIFBexDFGegNUxnt8
mMRdtPQ+Bla/IEh+Y0YxTCJOW5wdq38+PQe70AAFJGHo0kAvsA9291KSfibG94gk
m0JFupdt818iqGRyr2ZzQ4kUkB0X0Q8BHyAkTYd+GOR92i0vfkaJmNRr03xXlzN1
Jo/tW1SDvLB7ToIg1BheeefSyNYlfgSjeYhO2Hd+e6JHUIhT5irF4PXLJT2ZDyLp
Emz0P+f1yV7Ji61Ohb1kXLPW7HPztyU4faSbewFoLo8q4m2UhF+fslRPMFFnRqMN
CcJhBMTgThm4K+5s4PRXebUWK37gUPvJ08Ot6VKOukxQZjPN6TEJfwU9KLvWjRzw
YSREp/yE4DOZh82onW+/nqJmW3vTZm2rGsZEIHogtaXQvPHcAgbSQY9GZKquPEJx
Dy6w8VALBnPw/HQ6c0emnw2xTlY7sBiRBmAuG0fjep07cy8Z9ZsJmxY+t6lmyLKg
pUwvYnkj4uIHEAq/o+nETf0ekmEy/CLi46LTrJ8Deg/rOX0+tSLxgcN8O4P6n5Sw
ssOqNBpRnRwwzSKMwBRZI39unlQmfNtuUn2FroRVeu2K8WQ1en8aQeSyGcA+1twA
bvbEGfLr1a3b3Utmp8V57FU4R80tbF4BGIQ2RAYo5pRb1WDtaZpGSJQGHsOOn3bh
7zKenmzBstnVDhJtx5mzQm5R/Avjv2DQELp957dPO3UXGdWWeCbIBbAmC1wsNNJt
AeQVU4+d5Tlup370QCbTb5bwjvpFuV2S9mslNhSegU2tYv4ENzrO62nDe7tnzVbu
LxOxQq0XSvJTWk9Gg3Zk2dUVvvYnjGgCOcJQr93CnVCDgB/vKysMGBqNkRlNispM
a+lzFWvFi9vGCEtOSJZCQhtj2hn4v461DRjR60UAkxWv+cMtHgLfYLnjG3Ilkw9/
TGIfAbqqBb8lGI76e67m/iSoUSWyZIA9sgOANyI2w4h4UN9Oa6uZXiLu5Erb9evO
BGlLzlfAk7kq7aLzzuF4qfNCX5f6IWParW+fwZ/PySvdwOAShxImR0QZfy/fZblq
YeZo2dO6hor4FWefqlB7Pq2wL5u0arDOz6R7dzicXvjGvMSsmkP7hBnu34iEf21V
fAPZoI5Jb1pFuOdZEYvXLWkuQqHoxRjJzh0IfBm76NHEwU57P6kZ0M3vbZyxIJhr
PEK/J0kqjSqmBddEUxOa+xZZILIg74Ks7gub6yztVfILUowyo+mmUhJvKNs7r4iH
nElrWDqRHxtmWYp8VIZ2rvyeLXoXLTgMX/H8eMfjwNK602acB8FD6LRXiFbsFFZ3
nrWTdUnIkzQoFa8VNDH+Uzyfvm++jhV8GTIxwnuq2IPtMNgfMIrkxoy2xoarZZ4Z
WhARM3iEyGoUjrH7TLDd0jcpnvpSdQ8FODGMnL/wVgIn0j4O0xHssEqEG4ACKDqp
nxGTvDfnTkpaCduZyV/qgdbu5TKFKpONgMtila4+vyhJwaWMKmIdRgxGlrIAviXt
jWyfjuYUl10sjTwDsas945Febgm4Oje9HIkbxIwbgPA80ZKaTAjkO9L40f6MQ6W6
WBRDU6UMgOM1+F9IBJNaesEgm+rd6cEbOmczp5ng8v8QoNyOOceZHaXreBp2S1kK
89B5Nt6nqyjG+1MsLgYCuiO8k9t6oyxC7LEgFs+mldei1fcoQYi24EGZJhZ/IGRb
3GtQ920wjsHXpxGDm3PJ2lxooIfkwwLfEfeAvBHIcW19PoMaHw2kHuteH4r6r677
BBMS/72ow9pZo4d+YSFT5aak9uXkOTx1uT0DdNXLwWfkE+vQhCnyqy2iJc/cyVNY
zHQQvAPCKid+/Hr11sxlMXebkEpELvfk8FKYY+eHxqS9XTvMFeIE06t1OyhzZNl+
xEKEwkziaD85LsGwMD+ZRMF58GrssdMCKGEJOW6sgLtoTl9spjMGudgqGz/XqUbB
9mox/wRZr93Ic6BqVk8tt6GqXIL43qFg1rC3N2xnWgCwcnUDdoVPGnHX8TyMuvBF
R2hsGkkQlSgBMxh3jirHign8pQhlPusa+6Tl56K5c7Ex9DhExKarEYTyp38oPkG5
dqAu+R/VRUk2pj1NLXTjf9uvd6VYZJoSqRgSHCnKSbBJfnJ3QMmXLxxCucnZ9mFa
qqPE7d+LAz/luJJ1wCPIPhqiTPCGY6kvoaZ3XNhln88mOZqbtlKWXtSf9b7RjiGK
EDOko4sS1UFG2QH1mNuyjQnH2InP1zZKVF7HdbTOnsWM5PlbFvIeIYs4cmgCKeH8
9qdhZl3btPLzl5nTx1UolQMDw/7R4telV0IxBnUsvKMfKivQ/4XcDLnMXlCTL010
1Wf25i5s7gk6YLhSnmjPaV5F1/U3Du8fDz5POilxYLtw0gelOOQNJ3n2+nW6IAiL
VrImek0Hd8tx1exoeYDe8bT82VQg9i/ERLc8xWN8PxroBwz/HdA3gWLWDUN0n1mc
hPsu14APZDQBAL8sXBpRV3SI1uCiJ4aO87VfziMXp70ds8zZo54Nkj1wsv9Drceg
+E/QKZri7OIKmLmASO5MtQ4Hc9AhEV8DS4zn6lUL9fc0n3S+h6fIVkjzIJi6kRzi
5hvpDKNa7b1Fx0/jB5UYhYAoLak5nxfY0HxAGx7piDP2+R0MzwwIPOSDPKO8/rRy
6va3LTWQMYDdZ6WMU5EdkgooAtu1ADrz+eHF5Jq7xCdmFWuzHtrUWm9j4xB9UEOs
PvVfZ+D05T6Zuc55mUN/JNvl+su/O3+CH9JCeifFrrojYmyD1Waqf9ee2P4nudOt
Ch/+8St0bmMAhLtfUwBvIe6kyHIq+bFi91ifYxuip94YcgI0uakzgfDOsp+6xA1E
RdkbycaDOfMgfnIOHMl6XxUFCfA8E6ovNn/PICXeLKw9lotQWIYKTXnQd13ydzZl
eF9d7zhuVaFR55bfjHDbWudjDt8ZRXqZsG9LP8UanuuDc6zLgZtINoBA/vEEmR8/
16Pyjt3kGGVofGAX2pK+yuAIajPcE/LFeLQsOtYJFQyCiKo+XUCFwqc3KWUrPooN
98C7Ez6BADlImIhUQnEVhhuBsqR/+XuVmTM5rkPKRcUjmyu9CrAGWpdryKP6UcYa
4ezoROH3dVZn5mgBaUDsMrFrOPKhHwN4NNTxFgQ4yXUroTbx1Aw2VwFMazuVKy5E
QjNH5m9fzEP2bWr2DorxmHD7IzuA3VPXVRkpR2MGoz2D6yzLHNUgxd7rrf7Dw+JX
ilowDxaqmMpsfZIAgjkzTf1duL4V8EvtKUwWzMDW+aX3rc7mo8oKK5nksG347UBf
QFcdhz+8Ruu+deADPdU4XGCdJqQmSMXlSwbH71ED1l8TJPAJEo8EIvBWG0TXarKn
wv8QXmlxKXfKAeuIOAZk/PtOa1be0igpBpoqDv1rTVLmSmKcZEIcPmnenbsxcs7p
ktRjtSn1BF3V+YKaw1tNGLAG1mJaqFK57SIVbHQfoPtc3oeHmhQ41WpUfz/OZqsb
7mw7YzOgNQp1WBYgU1iYK6yxvDyPvECqNDo1F9vCx20hhkfMi/9i5XCncLzUexzi
3MDSfWToWs1yG4KS0GgDeI4CUlqECOXpuWlbXdX+23hnpYcQ5+/O9r3Nf7AZG543
ZiPWy/gAvRfHG1dIF/p1hvyaid2HwsHnfVViJTLUFGmTf4Hs6m+YIxAUGND0UQxo
vlTT2dNGfmlXPtlbymF4xhTmL/6jKpFQEvcdWa4xa3zkZL5WP2nEDhQghM/bb1Wl
vWCCWTzGW41bLez/Rd9Beew8F7Z4kSnei1+cSqmo/uzs/RUJnCtYabtlPy7bl8Vr
gCy0JQk3waE1Caiq1CxFmYJI9enzboGN1A7kMhONxu485ZtANU5kPLtmdnMECVnf
K5qAHBq0RzVtdS4mP8CcEhaq3FWMjQQvWkNyW7th2gQ1+VvpDJmFvk+cPPg/v1m4
AvY9tBGN2HeXtwb1iEUNtXJSho4fuITqyzqv0vkI5/bX7qJppuiTjJsbSj+2NthB
2LiCRlUvr9xKb/QFovpoLuplMEOVImA7M9qEkLPl1Y8fWzRNhOntitfOXEDdTmFa
gfnVIZFzuvQXfxWj5mgaZEe0vbVitP/Q2QFRN8tMHxdybrffHmkx2td4/wPrPT0R
6zeTRPLo1xtoh2ARXM4XjmC91sKiYkC7LpyJy1+niFxxTIrFpAqiP3gs9xHRkPE/
awbdlcCYNsyOUo2YJPA2+oVEcZeVWYNAdnm3xu3rRC6juVXos5MmjSN0sXm6xiak
RfKEy8JM1QbfcAAXRNIVDEzXoUESGHk3b4R1gB1sg611P3mFRpliuy248lgPNAgP
2z8fLNXzHT2Si/0AlSw6jVfSxJo0jC3VaNpKyJBYdrYN+rIrctacRXlVLVDmLWto
XIx8EhmRgQX4l6VSZVrWsvpXE+AROHIa30eUktL9QPC/0WDIWsUA9xkST4llbEG9
Xp/nPPDmSxJnBOGdcS+0sUdWkTQ03eaxuQNqged2Ie0p120K8Iqlg56Qq16WSCv6
1gPlaJ4+8M3pJv9o/MmHCxHCXX71Hqve+ZpIRrhkPBwgzF7gBhrg3M1LJgjpuOu1
Nstqv8PiRwEskE5kUUoLxz9bRtjnGg2wgxUa2qGwy9tL25EVtYccEmpQRDFpbP/i
8Q/GgefEiO6B3jnSWj9rHaP8B67ldsrVskMmbIokgkiqE6I+XImG53049wmQ0Z/P
w8ZLZ5FMhCPm1FAzI9PbApC4FCnT/3I5Cc48R8WWTdUFitMYpl8IAmJTNcq7/c16
GR34pSqawG2DgtcUN8UoIlQ7uebxfuoT6z6OQjRw3K4qKwjgtYXqKi0gEQ3rUbY4
VOJch07H27GT515CnWObS5yDaTlVlxzw55FdpA7SzFsVDoy7eKvFUNC8E/fOeHM/
6+TXynfBsDtu1k/Dpg8IE4eTqMQhj/D4pZi3hDMTXDH+T/iqJWNS6oAtSZ8frVPY
97mUXST2kyVIyBVr5mfCaKm89FNrQ1xZpEyam25b9H+Mv1N+HGFUxfHH/BHc/sOy
uClK2DC0VsMmdM0K1QKWwsinPWgQ1Z3WC7ybzYH2WzydIy6gk5GagNKUO+YCWkEv
bunnZqV14s140+nYE3HDDQ14R1NrnJoXW5X0nCC0nwuPESsmnAnv9lT9F/Ai1ouJ
EPb9PQJrVcJAqWAMDT6pJ+JHYaNph8pk4azBxDCL41Pb2aDcSdV2arzb6NQWCg24
Br7PP65xhgUs7NFT+4Zps/hoh7sFV01WM7D4/LB94x2WnfFWMZ27OhveMaJGj6WR
AiPCrKVClBFksbYH4gPf9DJTLWHsFQaCdGBhyFNV1xvAaN4yYjLTiQgxNpXdjFB0
VXF10hpm+tFKTXmtKANae3oKxG6C2eAD+cU3nGlXi3A8mRZUW6G15akuuRGaAXJm
8I+EX/t9tZdmnM49KnL9fMT1+rGF+OAju3103UkBS9zCblTO0m+NMjGxrW0Nsd4N
wuDmuH3/J4/j/9gvdMfM+nwO19AEYDbwGeOIJPxulEkF8GsKGTRUb1D7a6aT8LHP
LPymDbJmuDCrbDsGIFFxNC8wkxTCfRjZenLi74Xth+1UiXetHbufxrpN5nzvRg7x
lNPXLQHRKkDhzWrF4mg/rA3w3EWP8P1hQHvzCIHbPLN0uF4x11QGq2Xj6HJQrLKj
WJPvpPiJ2RgtF016kRu17vK2SW2J5kGvidpgEWrOp1TjkgvLK1y3fnIRUA7BgLdS
eG8vLCHvFsU/QvZ5rfFCYC/7p+bXEXsNSXHj6NGqDLa1QNpMUs5eqPa8DZbf8Y8C
+LFAjc3AX91Lv3JSoLNZgSAh/J1oRDgOUkX1uEs9lUQqypt4n1FLYIfMNKyHKRKO
71MvRZl5iUjXXDGmfMrNQ/2GR2lB/4W60yvVneaQdMBypEs45zdS5T0Anr0Adzs1
38jtUk7R2vUEgqCS2M3/8GPoDiJYp2A2wL/5Zktp0j3WdS0nmpL5AVBrhIZj/Ith
D8JkD37mKaD2f5SgRHhN3kXyOfAiBNqrKRFN4/EFwYL3Z+OpZ6scbBuh3aol5FWL
Y/qn4RZWF0W1BKZFK2/MtB5pm0AoYoWcC/zt121OzXVUim122SNLJs4iVMgevvel
I4Dh8t3b+Y3wRGtXMyRekHaxTkEhm+wsBQnE47ccHP92fEVigZQByuluqrC5ZkkA
ZhNujgozMAx5mpsz/vgiBldKe7qcVg5qAclzNW4YJ5t36H+UwYmhO9oVud7N5/U0
5r0HHfSYSkhYxkF9WWPuIj/LdzwkAWM/b7LzldQL9J2Aa03axjsDcqSyw700vC//
j0s6x0at6o9uTYpYlDxMf75LiXwRVK17VJruCm+sUlSe/FEoC9z3UvmR0tUcOarX
YNfPyoA3QKu31FFC79CFbGLjCj916eCY+FPT145xdKtke22z2iAmaDwFBjbJ2WqT
CXRIIyyk7NNjBMEjIX84MIUzkSFsA6Y6JgjiQs4ZC7as4Ez5AgMN0p+H77Qm6K82
LJ6Br9LC7hiXd3Y2sEUWxtk0TlySy8MIj1uooVWOfPwRRtXEfZj6A0ehfAg8Uy+r
EVSf8nZtZs79OeAQV0QXXUMdIrxjvgX68btaQQUJLRg6KIkbOCjAMroGW7BvvDMq
znKaZl5U7/XmrbO9wqgooINDS/mO2K5x5TZBao5MHe3zZ7I47gctKot3Eil/QJYi
sQAqSjrKuLv0GU/atoWYDMzgKPs+0q2nfoawIOfEYQGQIiCyPNX0GZR0+mtLjPKo
iWoLXX/Nc3OCG3V5BhhLxsR7aoKbWTcsrnvhREUFd/HhcabhLoy4VTyhK3JcgGX5
lG1O6zc7xa3jnrBV7IECqrfC2i0CbB56kpflWgo7LtXBW69zjKv9pPZOFGs47lJ7
8hU1alT3P3PSSJCZq+fD8b30s+Jd63F4ci9O5atwC1bkU3jVVxI6Tn95wo3sjxHh
EsSEFhdcQVo8W1HNsTBwGXj8QfBY4bpJx2MdY9wwoH/MaVCXxhqisthNAJEFZhvq
uhUIomTOSwX7ECHm9OR7+IeSn4XzzZW27CyVo5/U2Cys5+e+XyyJm6l5LS7Glxiz
Hl54l2tQF9XV54i7xshMx1ddMIWJIaxb5grZTlVlKz7XRyRToh1h/i1Ah2eNu9+H
qf28PgJSnTT1wtN39OgV9rAQuKIRQahmnw2REVx88prF5kb2hlkVNEnkkonZhlBY
ITXNMVLkrJCGlj8ks5E2/RDAy1UmWWMYFGLcPNKLyJx9OZj/LMUL+zz9XUKNZNQD
43flp4Z4NvKO3VNZlfqybR59OEU0wfUKpq11GoUcSfjr7XmyQYcc20xpMBRjAIQD
cPPzU3wCEdpuM06k2cTbuUTipzc0s7uOy5xEM4If+KwoyQbh9oXPVpqWflo/SEOM
6iO/3RgSqKTzi983JID3JVJ+at/hfh2ye04BYPh4sVBzSN1BSs/IGSwzmYvakFNW
GIGm82wjXfK5FW/k/TwCVylmnOViySyaHXqOfQezNSHDOX3Gmpdgm20jZHG4cL+/
INy+t0V9gLR8B85HfhpfczocxFQEFEtGOdWYNNvggFp7H/T0qMbYY9xMk0LOZReQ
EGF5d36SFuumfYHmaa0QcTPQTmq3/7KmwUcm2HzpOlc5nagWuNt0+MECYYfqXdef
2OD24DipnhkjI/5baCb4xe3oAys8ZYqc7HSAkBXR+VagHP5yibxOeGT/Jdyv6gCk
54qdYtrt3i9w/c0NVDKgYZu+keSWWV8CoEArE1ET0rKUj01cBcpK0FL9BhKwcelu
mgj4c3usHwvsUD+HKamRHSGzpDKi6ZQcL46c+xeGQjue4UOs181SjqDiXS/eO1L1
Qzqx6xDJlPVFz9GWphZsvM+5XmRlxGJfp/LfD+90oydee3oNiabzKhHVgxe5hazd
LKARudx+FxBt64uO7aVBsQfxbodNoSx1bsiZWWgITEqVpwQo1dDgfEAAaMmI1bZQ
TZz6avAvCkHKTGyW+3GQWEFnOLdaK2hED0lLduZezkrYRrh/n9SKHVn1bc7wG79S
7SJR04zA+Fo981j0zoTqwS4qdDHVrHa2mp/DShcrlYvqMUkD6C28ou2XCC8RvC58
6y73zz7H18Vj10SCWNb6CawSqd4okogpPBGVMQwW+oetl76Idjt/OhGLaDLyH6xO
+w1/l9lAKHRmqV8YSFKUOdPCAg0OmxposNifUzzlTBGcverJzcHNVaWVfR2PuDpq
ntWBmifP4xRy0PYHIkdDx4c/HkIPtBW/s2jOUOn1GB+cluzxL0Cs52KUspH4dVOs
N8Av9QCqdT4Hn1T55Z3GW6MpH99ZSZ7alYoRbjH/RKL2iMlQG9TQ7ZMbUXbiGO3C
u/wocHsos4W5wtC4BlR3BKAu1JgdZ2omlVy0qJcoj53C8TQvSDNO7jBNMWc7CN5/
ckJspSi7FbBiYwhO8wKeqmQDCCWJ2XnvkquFOqcY0UvqYT7tPew/XOnCI2ddNuWS
w0Aotbd/haNpiCzewItFaD5Y3jQTy8ZDVXxoYXHf2r6mx9pNULrmSi2Aq3dszd2Q
E60OrU3RCIspteo26aEJK3PyaVhOVVkDu3ZXbKPieAVGOAUOsLIDItpNGOdcY14B
Zq6dTtC/EUrQxgWVOeD7zkW5SuBsnSD11eR2lToJyiN4mlzGaSD3zfxUqvXsKpG4
sbiQQmCsIWsoTmPDZQOPNyPBixUUfyA5tPQ42cVMhiJ8tt8ssZzR1JzMhpfxR5st
MnMcCU6BhWthbNL86pBb02TRFgSSL5Xv9cpzsMScsoo6bn7SMxDaWFtsoJUmF4Hj
2dCqN0LfBqVMFfi4OWpmGeDusWw3EQruRTUV0MUBu/v9r8io96DED8DUnbj0CxO0
QVQSRxwu9wZ+TCwtjef59ypLdgmNiSMDgh7y49JR+mIm1iJ2t3E/wMONZBwFXC81
iP2mY7/BvvVrmvjl5wfRJU40fsgroWRj37jNMlWYp1/53CE6fI4IdkxxQT6WF7dI
hwWA5WJI5JQxa6rmmvV9FBWV2LdX1e7cYsGNes/MUvvjg3gZ4dWM7xgHvjF56+to
F1+j0HuLVHOhPt9bKwAFNHDMJShUolbhx/F0Ta+6Y9CGxihtWm6klcSmSq4s54bs
N+DGDwSKj2vDthHYpPl0DSTrfhmVGxqCiKZUt8vpMkJ9niFubmOELVfrhhYl3SDf
LpYFYAI9AT3m9uRrDZQ54ZOz/LAMenFJxlthXnhDkYZ6j9rI/daUfqYSLHWo+lpd
nMXvZqs87CkXEAZ92GLhoOqQO4ih65rrnsXZYVNqHKbvj3moZ+P/XOknGabQRJSm
fvcggcGrTrbNNq7a2y6AVge0JvZk189GIPEpVY6m37XpEFbvNvF7jMU8ol3Vl8Gw
smyVB2+l9/hKyhMTEHrs/MVDnGaYKJYM+Obdn8WVFeNJmiAMv07wcjwnzZ0NWcAh
FR7utUkBgXpz8Ydt+i4quUgsB9CBXjHSE3+/zUOk6Zngr4ukGx6xIzFiSvj6arS7
3+W8Zk2whI686kW2nRFJx3LpnVaqwqk9puTcUFdrDIgXhtMm17X4hBIwU5F5+BQ9
GpoMrP7HhONXIzqRQUWuKVrhatGtQZe42nW3xg7Vykrd9mL7zM8GXBHYp7ANzCU8
DCnD+rcT4xG7tKIzLEHAokKmgKgNpfmCWPEK3EHgAmsKdVJw7sXclRYiCrewnGZs
LSCz5KzbGRZkAMHy/if7GXx9/W5XfACKlotwYHTeXox0YZZkYfNScDl6oIzvMhZq
073DES3919MuNfu8opyPSazulYNhFketIMzumPegF2KTtkKF8eugCj5aavbfIorc
R8qGMs7hqSa++wi8Kr4uKvyzYYMRvJwmQ0d3FByApAVjrRSlhqZqueDyAWWGD+47
7ZpG1veK3Ota69l14BCmHuuoLElGiKgi+H+KO6T94G9w2C5vFrIHN6svmDB8DwTW
MnBrAcjkpaoojVRCK1r7b0W6AJLsFpcD2NCbVxGBiOG8vqKqNLtitGSpQ6C9316m
bO2ZNrJMMs1KSUzRLgpI3yt/LZPBOECp3lhx6dpTjoHhTKKJvh8kg3rWYEm/uLVt
OzGwbCDJiCKWlg54kojQk4LTm2l5gjmpyqAeLGAJSD3Hsq8VTB7YHZ2BTXO3fV4x
ZLd/FZv8Tj4wzROCmfRl9jM6l8U79KERwzF4/p5W9zH584Ln1azyfZqG8t5nNpaR
MsTieIt0Dfmm+XKuMCYHCx0jwhOpoQ6cVbJ+4jJOHqHj+0cYfYze7Nk7xKcgt+lT
Rj3DefXu6SqGyWuxgXbCgK9QWLK2wHrHJ6zLAfoMVBCPwwR2FOkCakHP2OS5jeot
vl21EpZgT9iRpVLfrNd20xya/ZpP8zmDDgk7rwHQshQ7NVlZz9BIozZZWK9mNZql
od1IFxpakJab15nt2SY9aKrW6jhYkjnnvJUpcafkz5Ax4rcVH6XV+O04jbw8SClt
SkNOuE44y+3VTo7mwuYuKrO/n7k8i8LjDLaXukal5Kcvz5f/LnUPPO/Vfl1FVjL0
lVlRqwgg9isQBY044QzF/W5yzlvHxhnau5+HKRMh+OuFdcpuuSzUMdbhhe5GRF5r
i/VuWW661nWSzr/NFewwfsaIwVnTCuA1WNqeLOcfk8eMayjgZiaHbu8nrDDmU/n0
H93Hi22AZmtTs8nLX4Amjiqd/8n0hUj0aL+orFWsQCWPs2cO3HOsb+oeib0bvsOx
Mk7RYJ3fGkfA/ppRn5nZmjZYOnSVZQUJ7o/aMpvhX3Rq5FLvGbjixzdGwoe35Ng/
KQ2+V0BgX0mDZH9D7VqBXdLbJQxiEuyhBVoIMs02zfAfyT/YCyxNWnx+zTI7s9YF
nIDFRuOUoZSVdofvnvuEidZTDi7QCqwGuYIMBVoGy4Asg7mYUwF+bADRmkEMz5xR
8wtTF92vAzwx1izyOOx4fep1BE9ALX7tx0MH1je0NSLhzwfoPaBQgiwOwIKcwtFe
8/YydB7/ouZKtEV4ik1JzJRloL3bAlIJ5NtB7qdUs1e45gwKOJNTjAA04CqLwq3W
8vHxFR9WxPU/Zy3ddJtrY8e09UELQSB2CrlN9XuKYQqb13aa10j5TTNjKbCYGqvd
neXm/t/Syo1/e+0C/nTLT3CrHCRSr91leuj8a50ORILCji74aw/3RIJTWoOvGC1l
Tw/jwKlHjM8wqVTO0b54mGhGaPRbRhUkVRgRk1T0vD6S3G7j7mVvSSRv4FOm5Q8g
wQvaox3yU6Jqn/RMh79zIt+C0HeV4FLI626OOukEMcv6JBOsOuYA2HugCx6OPKks
LFLviqw6rujYOhWfgQnSrIGlmdajMJWuZA1043wMH+8IOJoSmF03mxusHAImzr5q
OXjm26xzEMBi3ze+ow/cY+c8BHjVi6ZZH9EOg9DC7CoIyvIHAf7njDQ5Y1N4oKku
Ss2puiA13dUJQLzytQHucD0Zw5O5LaXqOQQEjWZed6vmWpYQBGm6EE4I1mi5QLfa
dps0WqycXFlcVf6Uq9554eVE9Vghh007JJe+OYVMN/WyjLw9hzWezc3IdLHPGijv
LIwC3PS3KqqJwlDkEAhKzRnqeQ2IsZqPEN6QVpNXWILRzRpdfoQ7WSBSbgshVtjF
BgZkooM+33F2oQSl3RHTEZQKpAah+deoFq4BMRVgvD15x74c1Xn5DwnkZYU2SGQn
qNh4Fmo54faApc5wR6rPsFhVEi6Nasug41vynzaSHaSLZcIw1oLXuMoXfIVxWVFb
foI403TorgGPO1s24978bWxMPl3UNV9GgFDrdvHJsZui8csBANBLt+MDTm0zJ18L
CNcwqMionjjcqG+VB+jYY+Sm/wrNjLxAKSD1j6N2NsNDA4HENjKbYVLyZ2r+GLB1
7asKcCHNBy2iELRFXuQy/AN3FDxQqw427X3wxZKU+x+5UVa6lPfqOrjzXV4oUehr
OzYwi8lrVK23gITosAv4cTMAoGZr0UnaE0HjpQunFEWVlGKDjGA5ByG3YXkIkMEZ
AZiRqzSa5JvzYMZmLy4AzeJ/D2u1Ogj8sRRmkq+n1fSMFZcrzLnR/nBJNSIhpW6Z
hv5WrFmCrPvM8mOhU5LmxobweMErVdi+XjE6X2RLBuhLJ9P7X6edRI2SAKdmngyH
HMDOuTZklyvfAes+juxnitTXdeIzSeShS4DyM5QJSiS0WHatSk8qU3R95J0YrJ2r
vZuaLSMsauZENG4qAzELQAWDEAlFRZbeBWzXsTFxFExkxp02kbePwxcxq8JcmYNR
1SZSoth9O+Mro3vbF7mxmqVN1kSNwHXTjBpxwMx75iXBAS67Nwo2tpyu6VPyhu+A
t6MRdM/SK8TjO5YHtzPvLw+iEf07MtTbdr3jDzg/jHdDFUhQAXoa0AYxbdY9fUgC
pD/GXPBinupCxQBv5xKsZIh43kWmkBEV5HKKiZceauvMqN4Y1Bh1Z58CEWsDBkE+
y18xIzXK1WTAOpefoEP/XA==
//pragma protect end_data_block
//pragma protect digest_block
d5crUjtHUXkW64BZnPM9o9PF2A8=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
kmi5hvwtBxVGISDU/o96nQTuILQnZstIOKJ7LvOUBWHBX19EUIE3GNOKTrt4aYcd
dDfEF9DtxG/QhgZFXWQGAog/X4w5k/sC5l2sr8Y0uaUIhuYzqdwq681+s4Rlr1XC
HzZrTeUmwqgd6Cr/OH4ZNM/V8RqcCqa/djJDgak36W8FG2yaNWD8Bg==
//pragma protect end_key_block
//pragma protect digest_block
LXwYMHJVT5VHvUS7DX04MwZh0SU=
//pragma protect end_digest_block
//pragma protect data_block
EVMFGE9chOxSk2eB7mIvlgR26/evXal9P1jvNrZmoo3tV0wxk1hgCXG9uvVKGcVG
dXXimzr19wp3KDqxOXfbJIARV2GqJ6IA9IgMHr7EY8A4Oc14HqxIH5XvEGNJGPVb
mBClEQqjcEmeFig6gy4DP/HzpAU72U8k4H6QawqXey3+YDirc4ikpEZwBH0zuVC8
XzmQ+FJNe5iew8tI5KQDjMDoyqovdt5wDzmmPqqGHCd+o+r0iFpxMiDvX0Ibsgdd
fu6I4qLDnM4imvzCYngTHVtkGtHcznZJvl/aa8zy7Pv4Gl71GsZY75unK3A/WAqJ
VakELgzDAn6wxDTKN83pcfEun9NmDkAS/zB0jIadUuJCliQ8YsQm6nXQJVLogiEk
itxb+YKAidwA2F2BLzBowWY0cVXrttdo9fNI9YDI63iI9EEs85maz8mCnU2ZVOw1
iXMjqLytXpo5v4I8NJhXlvhMCrELT2AyL+mYwtckEwIxwCD734JcGInTP/1P1c3c
YWYwzH65b7jS0DXBFfyyrJU6LV+VfOj2FC2dfpcXNZnx+qS7gg8agPAFQx2vX1Ot
6A3hs+HmIcIY98Vku+FEcvCJFWZP1ucRDRoocuJvYF8HmEsG1Lbzwim71zzRnZut
XJVD2xVkxAdTDa3EEB8blyiiV8e0PIkbHbjXVSsXVvVdC/B2urNEcxfqJRe5LYri
HxirI1FDur4+VjpdzT3Xe2o3gs+k35dR+Z2F1JuWzwXeAi7p2U5KPk3qOv6iZFwV
TqCAAPJefhXapkkKnfgOIEsXCZS5BeQzcf2d85tAMbdRlrPD03N+FKwBegjIKStj
wVVoxmRCRoPKr93z6yWFufhWE3vqtmed+OmMGAzPqiVg2yScWQv0KlDJIDATkSBc
03vP1HHomRnXB5vUXzB4nNtIJV/zlV4M9tEoIVBMKpQ8SEHnUXWX6aR0+6xm8+Wu
87KqO/t7qfYL3q9LQUxialMg0D2XwSwSHek/R+ktwfX3SHRhvGEq4MkME9BtUMwm
qypgJpQ5W6RHyt1NSxXdY/XGkujOpaW89p/6mA47fcQDIhX6r77QTnWGqKzfa+tG
BWoEtg909TzN/JalDwyPV1gKQAb4hKyVQgW8k6HxIUwJmhKLR6gJMF++R6pgA4os
GxjA9kBPHcaQuuyShyv/l55HzcwehBWM5EDwdR9OTwJCEBowTJ2mdJIaIIgNxcLm
LgFhO9c+9rfXCoez4Y31Sn2sWPnxOx1MYpPhbYBr5ufg88dqdF9hCERH8HYElKwV
fBJY1fQYvfEDoZBI+svQfZSwtXc4fyjBAxPbUXPXRZlpPLuGa5UdYAB9M/YeXyeE
yDU0Gdj68E9n+Zz/JbrE+BWU0jBEYfbQG7oYMCdr/yGVYTYvgpofjmJcg51fank3
M9+k9KG8XJnxmozjAXv76cncPJMGLMefMX03jLGgaChx8fuhgfd8wIIvFAMTyzBh
/uLoDFnpyHTHzmpYfXkdPH+By1AtZ9gHi51quMgUDFuzv1tIZy0jJYJPScOOmVrH
bkulYkvEi5Wq5z3XzNY3eE6oxuwubZ9aE6723rutPwC67PMTXiRftfMDHLMOUJ8R
n5oCsz0AaTaT7LfB15DfdvNVwOu2cXaqREUNax1IXd4uBorskxtfIMEOoW9bq2YO
dVivmLuPRr+NpK7EjSYJ5300szxuh5jcHnAoZvTOTmI+NCGCU5xAFbxcIe4ISJOu
492wxcWl68Etji3LrmhNoy+XdfwY1JcMZv6IZJshA5UrvIN9GjmPlw/jX7nAxTo5
zfSMqRdhMlts7rGuSRGYhyXBfadIM0pl7S7e9z/tsREPy2OdXdkuMDIiiRC67WoM
Nyf6pqalGATu6IF0ax0P8mKL09/xY2azsyav8RPoQAO83XK2jVY+8HsoxCfAtt+0
FXYIDpbUGJQP3MftZ9HxJe1A2TI1ITOaGPlrTq4nEDPD7kKbU1T6rW6nAzxH5/xu
5I7Iz55e+zJNhUFaFrw90iOzjgpZhPBCdrd2FHCgQwozRvhB11vzuX7VpuAFKh5P
xZ/OO2uKWE2JbVuKSOPD00tpurM9mmCEFW7x55KHjkzp545jlMybxMj38Opl+veR
j5TVenchFR1dgCvrCmfQEml4x8YJjcMGF3CIUKzWl2mfzufT6tvn9shg7uVUtlcg
5RCHjK0i3PfJ3uxJFHI5+w6nKjAS4HPXCcRjxY7A5qRQ2akR27kWSP19yBDoXHZP
nUI8muS7JPhSO5ebUL2naMBmp6Zp7AQqQe5gP20G0YGw/GchkbEsc1yevrBCD9my
ibHALAXYXB/6gWEwAvTnCc90oIUulVgsVhcWVlzF8UjwhALqTLAX8jHXp1SVcO6Y
76ZakjV6yUIzsrTIRkzqErhaiezGEk8NKpZaGtLBkOItzbwJy5099jY0Tp6wnE5x
k+bpg0UKltSii9XcLp4dyUkee/Usxn/46DYIBKLisSMirNBvbO5lZW+E1oLgFcWR
cl/mIkijgferty5RiEX8S9L6s4YZrTM5OAtcD3epng3W9eor4ox6DGaWHaoxWyge
64JYHGg8g4V0/GLMvgJRpNq3oqVpwVPM7Gz0tWmzpvsI0S1UilOrUJSOv5+VJYxj
bOG5Hz2alalAYUVB9SDKZ1c3ZsCKQ+3YIYnt4YcdmzIjKqiLwq+TuduXmvQ4PzQo
ArElvOiz5vobLPVH4sNAXzcYL0CkxhEgR7FnyWELRqiKTBOvevIn6AMSZO5XC5jX
0gQaPVDc0UOywJrUqyFfyYu/qVXCkAIbtyNAkEBorLQO4U6UM5oN+daawCiop4O5
Ck8OzSn7ZPIazsfjBQcc+8eYoiBSft1O4hhnsw8T76NKgNNS3mLrl4uexHNCZAff
x4h/b8Ht2F4jEy0IVe6HgXTLDo2OoYY+tQ/e9xXc8dsij/j5+Hxc9k/WExgt5vQT
vucIzRLhjCfXKZARK9xveGsvW0a2XU2hYAmj5GoOJBpJuho1/5QGMSJVnGu80doH
TR/kPgEe4QEnLtq5c9DETlt0COgOlkz5/9SSUU11fbzX/EHnCsEnFNCn7bFoHEOZ
W03Jj+HqoEq/P+eySCRMa+J8ccPQJgdKMAAcDGaCyTMGybhHpz6an0LzZA0XT3rO
0+B7s13xqQlTEYy3Vzti6TU2fgZjXgk2fAcJIftmUh5Bq+moxcWoF2mZPOWIaTHY
u4X5anlzWuOJ16FpP2Al5jY+OYgupgOdXLzZtycYg7JK8YnqWOTmxMpJcpI4Lhwp
xN0i5QacM3gJWOUDrk4X3naTfM3YQsOLP/VEs6RS4OHOKhvL+L7zj8ZfwsR/yScF
XPZTiURu4aGD5/ajFnKcJTeo9yYToyfR35B/bmMMhIeUpmuHRdkYZRlhugxCDS+A
YYk33znvdeRltx3eIoNld24S9MFJRljtPKJhPpTiZEZQReTD9Ksyk9DYB2fuRSzW
uk5Ae9TYI3rB1r2b43BvnsFl+8dFO7l/OSqXNvXSwTIWvA/REaJvQFWlBr8t73Vx
vWT6937EzqtCqr5dVI1DPmNWXg1jxGbdZ2zn4NB1gh9R9lat+IfYA3D/mOXQF9lw
LstJTYfnJtP3CdzcVHpIT9F+HjoJTl3L/w0+bw1vpPa1rIY7H3WU4+kICXcXfz31
FL5Z3laLfAT+6GLtv8vZz7xyzEONiiFgJu6kenQHQdpQXOe56qZkiMBS9/5+vVcy
V2F3aVx4o9KlJlgpM1CZUCw3YzNcWNUFvcxXpAtBzZdXOQAibUXxUS3aNO9fJI9M
aoricyI5cx3Rbn3xcL84IjI62W8XNpIOb9EvEZsOYH0cQ/akljxGoRLlC5J9UMRR
wjGcT7LHcuwoIZRwj77uQZlzbTHdpwVlrUoHU0WqM/tTUrUGpjKGHYmvBKJmHPxj
VqJImVjd2T5WV6SEqSOdGTRamjTZrF+fJ7exYHMhkUDUhk4k/GdGj1LTrYUGFd/d
2Z5+jJtm3zScP5GKBLShyppe2/fO2t4DmwaS91T4iILxp7M3sIXfukEBKCScWOyq
2OGdkoHYef7qSoHyhb/VYbseOmYCXAvB+w/tBG9HP8tYnzXIM1ugovLmyHXchTYu
Z6kA7HBTwYwjMP0qEJ/6IFTD+ZoK/pADvlAjxVs1tLx0f11wfLSV26B95GwLqet1
TZmA1xgTDYcBCqi21D7lRosyntY7Wui9kkxEI/JAROCHy9vFb6ZaNwycT8SD5N/I
2IeGmRkLqWMsOO7XKhayh4DjpfFt4tweF5uh5L8xX7Rjz7+1cRt5VkT5lXKe2jAl
uVx1IkGib4/9E9hhS874aOZ8n2A12sN3sMWLHtmqYMB4RLaqWm5itLBNb0t8Ncgx
XgAga0/vIAm7XqDx6ZljQP9OvKsuAm5C5j1Y2KB//sf3Gqh7rg5pnEGtVHzhd9Ut
IlKRteIMxA3HW76uOjFx2bJLtfVBeGqnqsrlzOQLZVBLxEBFBwxS64teLoTv+c6b
SD9swjOQpN2TTGEAE22p79ACGOoGWFEqe2wh4b2pYGy5SHwS7p72f04FTWj1AJa4
VrZSFrUPwUnj2wAbZ5Vw00LgJ2tvOpRq+AoST9+aITsx8yNVSKcXwFCmciKnuMFN
dK7SSDkf9Qq0RuMndur8AAnIJUX381WC3OvwTI2mgHT+MTa0vMNeRmak8HhOBc95
nNJyWSjFpCqX6cfW/oXXgnVTCY8BUGPz9nDUxohVoBeO3krDKrpPzLFN2c53B7xi
MxkXOh0N6U+fpR6NiRl/nNG3aVUPXJNjSj1wSTyTnlQ4cFmfXKexet6NEUI4RMDh
GA+bozeRNzexMWqYk3LtBtW5Q/UUiiajPIM3M6arP6psPw3tLmTRq8IC1QjjDd5D
ITOtWurbe8kZEKBO7X/1rH4hO+76SF3Q9hc3Tfnlq0Oci8P00uD+Q718LUXbEGHV
5egPbXvMtT570NR0G7fne42A8t/JCZyPb+HTiYOS5OWq5qo+/9KOCS82ZGCa7mqq
dBVhJSIJvMmfnuGnPMWsVX/fQA0UonK7WS5hz6pvixqTPbgYHHxKoPxLWdEJmKks
emjtz2BGkTEPe7E2eAykX1FbjPW9pbhJR+y6fUbTU0u6b8uhfz19RAVYvLApK09Y
QCsfTSLvURoCFDGT7jx0hPP0tFDZRkxMe5z8lHW/VCDAREYM7vqczwjrHgCHqn+Y
+UH0JucFxgmQQ1OlWwlcEgbupNusdTByZnDdU6fVdwf4qlQ9uckinYGBnYfG9yA3
uXxzWjGr8k3TXcq1lAH1LmSNwyh0zbhzBd4S96VqE9RT/AVIJ0vG2QCWNZNnTZh7
YVeXDFvqor4Gk6rpe0sYNyUG3CHiNrX2XD7p82RdamVBD3+uAEkKicfGk1b9nkpC
2ZbUIeAMNqlLhV9cLzXEfoTWSTzc+mUEbF7hv7ln/5uuxWrfK63BUagGS/tDiDXA
VnFCc60KuuM5+TI2UIrChxA3Tpcd9E1YJrbkkTZnnTLXHkpEkN67qasFZr6l4gzF
hsuUJLy5wAsXQdPAvX9sZ/J7LEJdRUc1el9n3bze3h94H0RGNAcCECb3i1UENNFA
05Sg69/UzDc7wgem9yE6wbAFTV63vZfzOEXp7S61oGaSMtnnweSiT0AN8GOriXV7
uhR9F581XLUktzg752NzEuvnkHI0OHz4GQM7JaD6/AQvtKICQncZywu+191t89QU
jbc7sE2svENK3+Y1z2xiKZgHKafnXTx4pKuWyr79vGeMZf1L9n5yIaZVDe86FOXz
KgbvxTjm/xc+b5mg7kULAMSuvqo5We4OuHgn2DA1HPrGC35yEiwjmzkUPDLZji6G
nv2CqRJBN0dRMdfoN9EFVx9rXAtFxswlVlRxWG09KpjA1tytCIus2SKnWf88p1xS
pxNVv7EZByD9EYnH466GkWfX758xlvgftFaAGPD/jSQ37h6oPLeDWFKa93mU/wLv
in4TygYbkJOeAOT8jJdzLiqeP3ybUC1hPF+xUiIUr5isordAj0y4Fiv8xVAXYbKY
BYO2XWP554RlE2Zx3I/C7lhoGz8GbHy1w9RbobCmi/iqTUY5VZKf2ARhzeU6IG93
z0CyGfPnKkKCvVru5qnElGSEWWY81O5/sX/kbipxPaopqRBP7Yvqoiu0IhSpgYX3
tnLEI7dz0WoVHP6QQV+pXcoOZ2LJzKVBU87Gi4hmzHY4T9JULbgbaTlBdrgD1frA
+0XTweAuoEA+jdleAXA1q5UDjlsr4BnrdbwTtnH9MHw08s+zeWnFG5Kr428non64
3FqRaUv0jBIEfRtKNKHADesouS5M+Glg4XjOCKwknr1JIRZnPsX2x5jtisXjRR6b
Ap1FGYrfyUwtO//kbgmK6+gX5gLye8IJqy2dt3SwB0uKAulaQ6O0gqdY2buq1lrv
dcXfSTwr7yRjTuU9UIi7zjXZYo5YeRbJ+LVLd54na7FP26CUb/d61JwSjFkPIUUx
Eq3Z26x/A0tbwExMwCEIuw9jOl+S0RkcRE+LDfJzocdcI6uySfbukmsAIs4fKy0f
95YtfLJfcaITj+mEuqesWQVdZzzNotQm2y0D01cJhjFfHEq3KL8vIrN1MKWMJgA3
zYsIJv53kB5stHWLuKplqe5Mj9Gy1sBr+m8lSFgnaApoWXKEq0l5oUVQ+0+zBB2a
rhBGsFH+7gmm+pt3ac1CLMKrz4OENWe2r7rndh3uh/Io8ga4hWigKkWoLTxVUxHo
r2a21DqCvEn98XmD0hFGEBfV75hWabOisBir4t30JmPuwoxq0IR00BWH0DIZIMzT
AhH/lcAxlDrAqdYAPAb3OcTQ8TMtnDmQa/JHNqL08o7J5q9ZsWRUKFbw4HmYiiDp
jPVGUuHJl6f0TZihKo3fxk5kWtfp7pKFqzGvq2IL+1IbPMU6wV0KcC4q3vYWeaL2
d95JhqUziDXf+0EEwhs2BGJgTbpJgiNFv7cENYDkM3dCWa591z8X/3XwUs3AgulU
6/Nohjm6bjEzq1vVA7yraMFCPZ34oFxCgknKKbBwlIs6fecIa+f2vuzu/QOe/mKS
7pAHNxkfiYfWqc+8iN7nBT0hq+hEWF3m7NEP/IPOQf0a9N2jCiV8MT5KsHV4RTNs
Am3dPdD12vnUMVCnlVcwQu4iyveVwv5pZvvPnT7f1pHr7+4Osgi2oz6F+dz81uUq
miHX8tYutZgaTMumc3N+LeSm4McMx35CF+TwsjqNysRc3UWXoGcrgPE/vyklLypX
KGNnWw15LgD/Wr0egH188Casq57ENkAEAcnUUx0Gp5CoeONAPLFWNyBli/PxGftm
/g38XOVeaAE6Uu4t+p1x9vhvOas5/XiuROdZHfgH03+0w2b0H11Qi4SBeY4waeuP
lywDbvECzhxnltSqADZhBvXOeKYjfjKJUhd4V9cqlFM0BJpccQ5F4e1xU6UlC+V0
qZP+WCCQWMrNZ+45zy598EQQEFbcR/aX50KjQ4xalLOWmQrDupMhi7+ZIjnm12bV
0IHaEh47G9XOCyZfa5xlLfamL3BzLM1YOIjRZ6V7GP+BdUgdfUdm17aQTI1d5mcU
Vun7uRRwvNWAhmu/r+dYulvM/vVOX6IzHVgrYRNVm/QpUnKg8zVgU4ymzXLYxV6W
nZuqJCKeY7P27Kzcu3Knu1xShjDMz6KwDhJwcbJQSqC+qPXAGSXyv0FSj/Q9fOPL
jY0Jw2hlz89iCEpsLAHyMw+RVsiWANkAQUR9SIdiCmNy+LL3XD3+QuFqQF8v4+VN
HGd263pIBiQqdHdDFXcDohJawnEApC9htgUKAFnirfvxePJj0RYYOohk8ouIPhfQ
Erkdul09oJSjQFaVdtoDcoUdmFQ5SDvN5etVRAhsQApBEl5NjUlxlSLAKdAmW23X
19hbjYpUztKz7jbY0OZM3NY3TBODGs2Mt+2vNILfRt46S/wTo6YxzopJhrJMeEiR
Y1KQHQ5mhDu70BaAbbrsuk1xOroXcBL8RBZuBE3bOaSn9SzMH/wegqhH5C5C0DAj
ZU/VHQJbt8my3Nkki4RtSKD7gqphc9WUUAJ8qu/jXnBCtII7gXmQZWli4Dcascj4
YEyxVCqm3UPYAoVp4+9drghiiR3kJhnVHTqgYj/gmLpAcELqJ1UYSE0e4kcOruio
dxIa97c450apxfV5IawxuVj1jcCo/IBj2VkE7+KxjIuM7XssxEkF83oWt6QqHGTk
fsz/k00ipAAzbLL2rRGMCB5kivDmFjV4baKCXp9wBNZ6dTYSHB53bK+E6TYiWy8U
HnDTvmAYYYKASflKXiNKjlf3lN6lAlQVUGurduv+UEFL89RpRnjvw7pkC5ILc4c7
Mx72iI4X7TSp8IJzl5FKRlnEKmD+c4pLr/mn2BRh8axV9WVo6SeKKCyCpd0mNuuB
rreKMvE0MkMvUq7y9NIl1Rfg+iw2oZ1eiahg3mmuSwr5vUWZQQOGcYiEZU6L66Pp
ItKqjOrXRHODicvzVlECaVLFso/jCLfkpDoxQHNiY6yF3fC5sUPxErsLJU/VtKev
oxm5u9CpU7WeMzledgBH0WiYUp0dQMQYxkl5CWp5WYF5NPg5Jaqn+Ej2f7MLYMXY
Zou47bPTIZoJM86iCLlVJ+F6uVybNgpNl4zfXPT3SMc1udshHeFCNtAD22F194Jx
GWIX7wX81ltzBPqguVQCH8hAs6W4av7m03SxmANw+R741l1rhe6pzCZG1slMxbCe
+y2RrwmV67a1i19GV78eRRpx6OtfAQ0/t3PRT1y8fvT368KDvQpGHwOfXVvpjsGc
/+yqIvQ2/FOGAd0dvbc9Kc3Jz+PyTlKsQ5Pu9U6A/oQSHoZMp3YMThwpnfOLzPSj
zBrM9n5ayA3gASGU81/K8XO5U6LVcQSCVT0OAwRbx/NOr2gj94kz8zpa7Y2EMpOU
+SYaCV/dTGhqq7beJ++bdXXTHGTqTAffuCNQpe1dy9lOuvk/gFBT1tHQlOypJNKK
PjDW102qC2B9LRMt3SEkWqp5A5j7pMTjn2ZQGYoLaKnprkH4KKQIf1ZyD1PSVjC6
PQ9slwHy9OPoN606W2DuRCqhbp3pf/PtfqKCnK/FEbOl9faODDeKU9ERxItOlukK
Ewi4Q1QI30ufbzVivb9fgKMoyb2B0HcCgS4sas0Dg/g+BzJix4QvtbxyoS3gFme9
m6W22WJ0k3/9ZqnYcnqUQZFrj3l31X5rj6ajig3+WSzg5B/Lj7yI1+APkl5P8f0S
W3MLvbiQR/pqAAdoXvUNhcMN9F0SBUnrF4S8N8NZm1iG1WUIAvSFwet/MgfgR6Q8
ASwTUXNL+tBc6D5XLr3QUFX4kgfdqowwx0R5SL7G6jIoyZ3LefThTF9IQ/lLTuV+
rySDqNh1KShQf1HO06MWTqLRBtfGy0Jg8hifx2+NLDl23iKr+qfPM25TSdbMXtRO
i4ygG4u3vomdIyx5qW3OJqXGJnEPme9Tl4TlMIYRzdyxUb03Yh/I3C8uFPKjtFSp
zdGi8mP4was/xz8fi7PQwWeuJBiqfjBQYsvwqUya+ubfohCpl4v2qRnKtjAKW1QV
TCq5JArudX7s4lpMikeAGDsAK0irrldyoP/GNkTvrc4Bui8F3x/fkqer0TNpXY6x
zmVnu3jVpvJHWbCZVWi8MCEOBDtwgU76X5KsvXtrNnDtEQz160qS6gyHWUitt8BR
oAlF1jzEogySo2N+6b/XKUMdxJdIgd/6JxdxsAiydrTM3YECpQ1xIz6SpPppGCd3
LNgu+a3Z/oq/IXsgviBuwnDYV4YDhymUPakfygRuA4AbAY/PiDawNyM7x8M1n9cU
cx96XR3jVlf+ZLicWguEry64j6oUNZ4TxgPHxQ2wXU5BC/O1cIJY7mWIjTJpMWU0
8KBNItahTM1mEB25l3Ah6Md6uPkMidawYKsjzK1nnq/n3Fjoj3MHNjy66uXHPRCp
Z5imQKkLxfdXweZCgnWZ71nx3nbSRuDy2/IXyzDsDHlhr7257azYd4fiyDvzfGZ5
6vb8Qs3Zszv9VQrCAfKsNvZalDl4IjtYdStpNX0lZXNTBVh4V1hJsGP4y007kPln
YgwAnbG++iEngBldzoBMImxtPgrBScIrz4WgC6cS475YLTEAoPJgM7Jx5NiRxXqB
g9ks1laW7e8y4JrolidZQP7jjBkWWHYvuuCvP3Fy0zRMRTwh0xZGxsdsCquZ3oNq
+9P/1lbUAOKpfAAkBGNFZUB1Bu4gDS9jK8RegIrXdXDEEzH8NTeJGJxRopLuw61l
JhTVTlL9MyszgLhT5tDsijGkyLWcu7oBXV5R7mhqlxvFUiG2vXpXRBy7+hyvDXLQ
+y2Z05wSBBCisyiHaaSfIzD/qNnmm2E97Y31rnWDRkvyfdlC0Abz8DKeRfNuRBWL
cWCq59/s7mZ68uYxkKjWmHtlUNrxKgFqwkHCj0IAvCf8mgbCrnYmpnHCxCEncljG
W/tajuWCw/LXU+5eLJBuBCIVaY0dZBtZRraABMxKZUgOdtXq88S3mfeyI9+ajdl5
qDqdMXhEqOyt8BotExDpc8kpp56ZZc64xlPnfqsLuK+QXG0o+ofpMOKHJiyFjQzO
3QSN9zCZDpxM2wxHEZ5ptsHtlxj9Lxmmj/QlV2ZuwrtF32bTJ43k5OdRi/tPCqzw
HujRbrmzyZ9pqFJbvo0JJce7fPhUwqeKqCVnBtNkdEIMtSZOB5XCGG2llC8+Fq4H
/BY8iPnxlO8lgj1Rdr8pRwZFaIBP4omdKdRlqUvy3In791q1tpUoey/uDLaQ0m/U
L540Px0X6hEAh4tcWWRrVGiK4xntndqEG5GNDndj0GCRlQDjbQeCGodYCYYKy0Sk
pSroYdGBNni/NK0cCvpzqAKzy/+PCHAYfxWXDKg5a7U8XmW+7ezaQGaO/1wsLSgs
kr0SrCFvWp6s3miQfIhgEAq8VbJM1Yp9zvUnh5KwmgrYjxmMZKXpSj74MW0725xy
OWXPVmPp5EAGqHhSW+7izTwFTWNAfO/DeCr2uPjPAAzmP0byGjbkbC+T5BPINufc
Nqj8seCOPhgiWYtBNzmIvjoc0GobFkKIgaznwVuybepU4L2323B5VcUvZ8Z6igEi
fxQPywvhdjjImS0Cw+CN1AHy21MaXMzW8MrYGSX1o+OosgXHJ3qYk7hVHZWyeSVy
VDPN7A3mbJI4xzSss1UiBJ+Zv6YXdS/inKjaHEhcVEV7Ba1M9NopuvIw3nngFr6V
I/+gbkqGwILzDxThjIXiuYrsUQkrEadJcksoy1Weg8vrnP05rvtNENFuIirqPqfa
qtIjiRVhiovJtWshXQMCP5TosSwsHJXftcs3WpzHJR6oLGN7SoLF5igrDF7EatyH
BgmilCM3RKXVDVKg1nhXwZRLm89MEuhui+ehss2XqTe7394brXfZwevH55NdRi+d
GSiiP2vf+BWh1YPgnyJ+3B2ZlqUefjr3UjGwkV3y+/zKspEjDBzBwOZE+evWLKn5
vJ14d6P+tF45wIPwt3yNTx0iDll0WscXZl8wXpaGN6tmeDjT3cehqlsUngGsnyop
Hp0uF70yRWj4jfPL5FK6mjkr/h69kfkdr7NFeGwEE+UqGYlOxtKatwIr2InGnXRz
sRakoCutYb1J2uCZVtXh9/X+q+j90Nq3JYrMGPVuOVNqwqiPF/cdibur84p4N00u
hAKKZ6FwDCGBHQc/hBslDXeWgeqLTGYpVuEnCa3SOa2hQyOhSnupxV5GnM5Ko7jz
0jNTPyULrKgUiRFIPJiVuvU+QMWuxnNqfb4S5krdSaZIVKql+N1zNFe7mZ8w7Rrq
vkIWsxbazr/jhI+Qad4Aksj2xUifjn7IyH59UC3xbhZc688uN7NLxWXZfeZMgPIO
yczEsrITUHelwSWN3QhQLIMLONOaSuleQK8zTDNj++3YWdR+K707IJXcEsJSeUCf
K2w82tqEy4CvS7cTAlf0U8m9EiiS5AudBU3oAIH3dt9RXO+d+TZpwDl8OizJu72w
XcT8wo0pkz4yqkKTgIg+N93ER2mmVHp0HdHwo8DFYl32NtCTn8lO623t9XEvFKg5
tHt2IUU+QwKrAB4Jzjui7IBe573bT4khCKwKxR4GM/SqPmcVszAv+C+nZaAr6NPs
DEcxBEIQkbuDtCcOUlIexi3l2VA0Nm6uH+iGUH11JLHr/D6EYmEcgaZieQnvof0E
0A8oKPYWtJydVegJOPe2hyUQxQ1ZybxqiEpKteAfiit3HFCj8mHcr/dzWaxexRMu
1dkcYaUVOptGV6z67zntBKSbr1Bw9yriyXR4uqhXEHM0hf8mFxQ00spDACkuvXpN
h3PHAJQPFggzdJ2tlTuheNP9VCx+Ga/byhb7nhUpy8Mz2qqwPuxV4f3d7EE0WBT2
mUIpdEtTlatBGbWh1+tYSrTWAmQfdykT42jxmv342yPZaEPfaRZaYB1Yc1oC+Ds4
WQIiJRkocYScBGONxwHi0/pv6McijhE9bHI2OJZgrwsQ0D65bC0PIqCS/whs8bUp
xG+TxaUUNC9Old+8RtZGKiyDtZ+8EGVqpwgxGoKQ0ACDrOE4/5WQP/fz8pvGlTFH
1CwuNqOGYRV0e6R1x4ec6BXIuVElzcclZFdaK9Cn6rRlBFufh0kIBSNsQ+n+qsKK
wdz7BvrSWI8/1F3Tdd+s68hpOsGNK3hqacA8bLU3HF9IkI3JW7AKKdWDWYbRWXhu

//pragma protect end_data_block
//pragma protect digest_block
uLUAridlb3a/qV3tDfW5cf4KScY=
//pragma protect end_digest_block
//pragma protect end_protected

`endif // GUARD_SVT_AHB_CHECKER_SV
