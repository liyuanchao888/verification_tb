
`ifndef GUARD_SVT_AXI_SYSTEM_CONFIGURATION_SV
`define GUARD_SVT_AXI_SYSTEM_CONFIGURATION_SV

`include "svt_axi_defines.svi"
`ifdef CCI400_CHECKS_ENABLED
`include "svt_axi_cci400_vip_cfg.sv"
`endif

`define SVT_AXI_DATA_UTIL_IS_VALID_MASTER_IC_CONSISTENCY_CHECK(param) \
`SVT_DATA_UTIL_IS_VALID_SUFFIX_INT_W_CONST(master_cfg[i].``param, ic_cfg.slave_cfg[i].``param, \
$psprintf(" based on master_cfg['d%0d].``param('d%0d) and ic_cfg.slave_cfg['d%0d].``param('d%0d) which should match", \
i,master_cfg[i].``param,i,ic_cfg.slave_cfg[i].``param))

`define SVT_AXI_DATA_UTIL_IS_VALID_SLAVE_IC_CONSISTENCY_CHECK(param) \
`SVT_DATA_UTIL_IS_VALID_SUFFIX_INT_W_CONST(slave_cfg[i].``param, ic_cfg.master_cfg[i].``param, \
$psprintf(" based on slave_cfg['d%0d].``param('d%0d) and ic_cfg.master_cfg['d%0d].``param('d%0d) which should match", \
i,master_cfg[i].``param,i,ic_cfg.slave_cfg[i].``param))

typedef class svt_axi_port_configuration;
typedef class svt_axi_interconnect_configuration;
typedef class svt_axi_slave_addr_range;
typedef class svt_axi_transaction;

/**
  * Defines a range of address region identified by a starting 
  * address(start_addr) and end address(end_addr). 
  */

class svt_axi_slave_region_range extends `SVT_DATA_TYPE; 

  /** Enum for region type attribute 
    * - RW   - Read/Write
    * - RO   - Read Only
    * - WO   - Write Only
    * - RSVD - Reserved
    * .
   */
  typedef enum {RW, RO, WO, RSVD} svt_axi_region_type_enum;

  /** @cond PRIVATE */
  /** The region id for a specified address range.  */
  bit [`SVT_AXI_REGION_WIDTH-1:0]   region_id;

  /** Starting address of address range of a region.  */
  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0]   start_addr_region;

  /** Ending address of address range of a region.  */
  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0]   end_addr_region;

  /** The characteristic attribute associated with a specified region.  */ 
  svt_axi_region_type_enum rtype;
  /** @endcond */
 
  `ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
   extern function new (string name = "svt_axi_slave_region_range");
  `elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
   extern function new (string name = "svt_axi_slave_region_range");
`else
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param log Instance name of the log. 
    */
`svt_vmm_data_new(svt_axi_slave_region_range)
  extern function new (vmm_log log = null);
`endif

  /**
   * Returns the class name for the object used for logging.
   */
  extern function string get_mcd_class_name ();


`ifdef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);

  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif

  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);

  //----------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of
    * this class.
    */

  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */

// ---------------------------------------------------------------------------
  extern virtual function svt_pattern do_allocate_pattern();

  /**
   * Simple utility used to convert string property value representation into its
   * equivalent 'bit [1023:0]' property value representation. Extended to support
   * encoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit encode_prop_val(string prop_name, string prop_val_string, ref bit [1023:0] prop_val,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);

  /**
   * Simple utility used to convert 'bit [1023:0]' property value representation
   * into its equivalent string property value representation. Extended to support
   * decoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit decode_prop_val(string prop_name, bit [1023:0] prop_val, ref string prop_val_string,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);



  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************

  `svt_data_member_begin(svt_axi_slave_region_range)
      `svt_data_member_end(svt_axi_slave_region_range)

endclass
/** 
System Configuration Class Utility methods definition.
*/

`protected
1X-58JW.3P]]6K1DN0LH[;HgTDTZY=]W-.08:4=Xa@;eMNJdC+LL4)[B/Qde\07F
..]OU,@E]3B)Y3S)WA]@1)7H^-Y&d<_>TW<-+?OKUV8MXY9\-RRGf0_[>PJ-@Af2
F,KXH<>X)bN,46L+fPF^[P29U8X[fGGd0-;WX;+&NB)#GHMc.Pf^M.EJG2,=)+gM
>IXGSba.T;7AHJ7SR-+ME@ZBbc0S95N+6D#caQA6&?G)LT0<AdS/L0WANVTE8Ya?
ZWC_TZ@-?V<L(7T^.IG5QdV<:13K0)a4RZR[bO7G+X<\3QB,Ba\M]Eg=e_MY]La\
9S/cS0Q:=<IcH=EA7EHLM\a?:cbC9.aN72CKL:IFUb&GaEU9]BSdG<US&<c6&SG@
D[7;DM_LXSBNbcX)R6fa5([=;OdZCB9;4HG9RH]GWfDTN@PPg1aP<9I;VE7,(59D
B_;bAGJd1ge3=\OM&\6\L5.E]&@OL<eQU3/16QfKS,dZW:a55TaF>dSVG=CCR7A#
^O682dQe1\@:I&_:/.I1C?<G>gA_7J:MEF+[OS;ae7_g&DZ&Sd243#_IQP\X((>c
@]FG7[650,@P;(8Q],eD70cF;Y:&N3KKD<fg[D3_\0/TB(+67[LcZ,LRfa(0Y92a
1Xd_V[eS.QeD52W&UTXIF3Uce9Y#K0?-:,Vbg?,C]8gCEb[I6CY[&QLRO$
`endprotected


//vcs_vip_protect

`protected
=B>CQ<4/<YC.J_8B_NOXR7:FcOQW)#^K_9FFB7NTFT=eP(I]34Rf((-P>:R7f&aH
(eR\cXN90YS@5b<JD2eEC@7USR80\UW&(_LE;ABa5B@\[a4G1gAc?O(Te@gegLA9
f3:a@I;DUM+>(B67+7C>R0_;Q:OF^L810XL&Y[P>I_L/e].T3&G=(>6b@S;T#RDc
D74LWbH<ZN=]\9(;0JaHG[?b,1g3Fd]Gf;D,QJ/+?g9:6GYU.aX4f03S@2QAEVIU
fX2-<77KUD;\]GS?9>g5E(dV)+AFX-T35)ASLgCUC/MKXeOH\Kf6L9/\\Q99dZb.
^J_eb++26VJfWE<f[cQ5__0JJe.R/+)SO8EFG:O]1O.S-,,LN9R;<(4ZE/E,G6S0
B4V3U(MdW#S#HKJ5d:f9_D,EYMbKZedS@-/V:@cXCe@>+e7X9UZJDM+TaC_M(5C8
J,fW;6IdBC55dMM>0UF]/&_EgY.Rd_I-UFFE(&C+E\P,T@__T,0HEJ5XFaF356J>
X3\^F#AIfAaN77.TI(23-P<SbdLA<6F]4N\?UT^IM,6AV/_P7S-.P/G=3Wag@6?/
0d#YMV/eNXH7B#gOV5g>3S5?fKE&>>G]e@K)[/+@1JH.6gJfL@?L9_FTLF?C/bgO
Y_C_TD47M42233V#BX8ZKIB]+Q_KALM=\H8H?)gT@-MbD/Kg1_7Ef@KcV5EC7LE9
N_>214]2V3Df,\;V^XEU6#(S_[8<^T.DZ-Z2#F#d#5/IeR>f=^U:^.>3STJ>#=aU
,g]]]O\eACMM1G\DH)@)O6HfO31P]#-SS/Z]gUaO=S=_gd9N^8I69RXFHBIP\[V9
7D/Y3Z>R&aXUXI-9LD+&5^e7ddY0HDe(BQZa9=^44V&]M?<BG76+gME\[2S08gXK
R1,1b:a/7gN(=W/QUV,2,[2<eJ3=,)N?](g7b(bXJTbg7:W5c<THEF?VRJ+#XgMa
-\-+a5UD)+TXHI=G#aEePef4([(/NVd??&beeC>8&5DNV/gR)T2M]TGfcP?T#&YG
OY0CHGNL7J,_J=aZUEV#J3H4WK-_9&(O[^7PZ3Y2BZ8I<)&JFTLCK/H&JDLaPJ6@
E:gd^HT#VM+8.Ee4V#OWXdFb7-TK^X;K5HGM/b@;e9QV:\U2J^=H^;^RB]_d25Q#
WV@,5P@VM7#P[/9\28D:EADX1E^\1A@.I<R>\KBQ9S0NeNLaLJLC(&7X0#C5JCWX
B.E9/&FdPMY7#FFeMH5K:W1&Pf[R[\(W.P,?dg5P\)<+6C+C0=VC8P9HQ.DROTLc
XQd?SM,fJ6b+gA((fQfc[d\/(aWF)NUBgR=)T.b1_^21[F.Z&OZdI.Qa14X^WbV:
&^gT[E)/P0e3XCD8EP[@.@KWI3LY;W-P2Y09g#21E(<)TbK1W[NaB<;DaR1Z:XC^
QKIbH=)F/#L:dR/XWCD.B7\A^8IGKNH?^Z^].VL\6DEGUQa(fZ,=&&\d4;&I9D]#
9fG:AfFg.A;-b:H+cFbSLde6;F,^#a4d7RI^1:1NC:+[;f:2S\_Ff8D3\X]Q-0PN
W:QR[U(3#Qfe#1#8<cd.)aR.aaIIb3Z:VebaA8.T#<_=O0P^,DN[UVU0<C44T[+N
]&GSVAL?d8^QH3g)NRX:;B3Qd;1/?FHJcS+9++48/#2I.E>8A7BQ1NW4<cVc6I7_
g7+E<_a[P>THQFa:;0?IM\Y6E]JDJf(d>,g]]/@.<9H/DI@=5]EUPB#P>XD&N7GG
P/T(<de[gJJKXRJS8cXg_:;TSV,g<T4L35MJ9H-aEXE;d_@_K#C&P?d0RESVMP6(
FT3e\/,+Bfe0/).F#ZH6A+K_dede2QgGS]#D)bb.Z/>M)T,X/ED@EYJ>e+<5LUHe
#[A\Ia&CG)9_FbWF8(EFdRB4RS5F93GQIP=X9X=2[LGI6;M44A-LB+/T<Z-1]3DJ
dMKJUdM14SO21HD4\^Va?d<]#G#bePD=VUCefRWD+KKQNPEf0=5XCeQZURCJBaM6
B\ZYI(/TFAQ@EA76MAM1\c?BE@f.6(a])1^/3FfVJGP&5c;XE&<LV6^YX?0BT2eQ
0+KP/Q&C>I_<1B-,0eC.>57a\T)/DRBb^b9d<>C3OSOTcOH^Ta^dd+V8Da=,[<#Y
.?R&<9A@QCSe:V)B7:/OCKLW\Y8:Aed1JCM-\WaT&_/c#c()b8[RKN/+c9H8LVf>
?a^V8Xc9S2>Q+g83BObQJ+c</gG.;N^@TCD,.T1[6/dB5aDdYV4\SX3&0[N0YLV)
/MH>eFY.>d>05XT,VY=38=dQ9)J=NK+3]N;_&G]X6CI:/0:E(ddIV#WFZ)B2<H1V
[S)a<,?b[LIPdKMF(8R4F:HP>Q1FR-2fRHQNa_Na?#NMBY-f.OcQR6//5SF(D9Ef
2VAV<;c=O]N8<P<_OAXV7V<:_fV+@?#^gF^\13X#^\2WVDR)1IgHAO;OW6@P?@@X
^58B/?c&<?>_>XOSa,:?]_;(@_&1?[;VOE;44A0K7?H1G21I[\LKM2S&;L;gga[f
eN[7fHf=+)_Q6\fJ]I-BYf#+=NM+)1H]^5gIJ&b@Y5Kf3^3QRNW(OdNC^g.EN_K:
#L.9(&&Z&,9,\DC@0_,LTdTH9@<8]ZI?&&H1<7+d6V&,D9;4E->)S2b,@==;XG=6
4g:VR[E54&BGf)#,.OO(O#Ie#7\56Re5W^?IGa/B0A_^WYAAK(c#^K&IG7b58-K0
/T&=eY>3cfc[AMf96+O\f@EacR\f10<II[VCEg:7)dV2O16(K_cI<X]8K+D#0?L<
@234(bW\PUZDW=BMI)A8dFTJ0a<RN=Bd)ET33FX\H(\F.(MFRG642?E2&T<EZ[f,
A0>FN=WTbZDfK;U,.HHM9CBGJc;f2/^U?4#RA>\.UFB>)7XT?F84VAN@:B/]MOc;
Z;N4W7VO-T,0J55M.+00e___UZ)@?eS6W47VC.VMF(1J8;U_QHN3YW9@c=1LDF<F
5HA#XKYM.AFWI_,Xd;DP=FP^g\JcA.^KLRMefCc+23WL?55[F0DGHW529^=gL/LR
a@4]P:MZPMPfJZD#:MbA4H<@;/cceB\Q?VS]W5L;7Bec65P7P6+#SF2):K9O,_Cf
g13@=#BfS\HC4^P^PK=\B>FD6g>OaE?G;(2T4[+0VV/_,G9)2JAY)GI-Mge2W<C[
Td\eDLWYc;UHVWaaF/CdM)H9UQ1W:2IT6b5/[6(VY\d)+TQ5G3W(=JRVDAOK\I4+
:6>MFTUM#0<S<IVb:X/VIDaE7F+G?0]-5@<BD[5?;38P5L;A0FH1ae@)Y3#d_8aW
e2OXW7U4c7\c2]a;+X]&E6KZ(a9,)O3BFBY7IMV)90BH^EaRQ4(AgQ(X_^P3a5H.
W=[a+RaI.N1.I7MgA)Q&3acO;M+9C>24;Z6JA#\<QS?.EK9K,?-I2NJ5BE42D)MD
<.&I7J\TY+A,BY9:5P6L&RYWCK]7<M2g0HW9U=-;[KE-GIUF]e[Z3bEeIKG+VC4,
8#>2@Zd-CJaVRN&Y=OWf2bUURefDCf0>-KB7=6PQGH\=]>D=FM0g\b&cbHPdgUX=
PN[T8+<?SJc3K7Zb(:<9@b8.GEgLR+.KZI9=.:[d:f_#^d6?>W_6HAM;6706O4_=
Z[4EI,P2&TUT5TJ:-I]NcYb]:FRL]W)<?YJCN)0_L[7ZTW]/e7HZY&,+=B8[IEg]
\d/_B4LJa\D\bIS#b#gZQAP,(0XJXT<<)N.O=AC&])U^B69=T&KGGa6E^Bd6dUT#
4CgNa1?,F_+)@IF,Z\;<,)[)<Q#\1+KS>/+PcZ[Q-R8#Z#>PH<&XB<L0O?EdDL;M
)ge&&)M4fEHf_4P5LS>g_64M[g^e3@:6-ZG414&2?YYCe?S7F^FBdfZg1@(6JFg/
:>;EYO-I=I;ZP_]V-dV-WNIO4VQe,K5.-f-\QQ_YHVZbHGDHFH+\5ffJg>R<,eYO
C\L)D4TfI&McCSc,XcIJaKB#CR2TX6a)BBZ4,BH&L.KZ)c[^BV5RP5KE(V:e/gR1
M4G#&&2a[#:dH:9VCU?X6_TW0WYKX((aG;:&W]fVe?;@]RLLP4F=]QP5-=J6D>PG
>VK=e)B3>TK/B_H6+G]CT/7L\cQ7:+^@)B)9C?BF[1^>K3LHRP[Df>:aSabg(;d;
9]=TD^9^4?031Ya68;Ib=bV/b&KScC3KEeAdOL_-WKfd]9T[b_C<QNE9AS1NabM&
.RPFN/.=[Nd:KINJ&M2F6,2A-=Z#RPZP((#NV2&1=.PQ#;beOB)dH0L<U6B8Cb3^
P^]d/NA2<6aSRX>2;1UFEH6FTYFF<VA7OK83[MOe4Y37L.#0?<MFDe]fOdDF=^K\
;bSF@CWL[bcM<DQg^/OGI[O2bfA^9\<:3AA7(E9+)WC45gNR2.?0=cJXQ_Z)00<T
4,eJLc0Y4&S<Ab?=QG;eIK5B0T_-Y&P,YUQWc&HD<:K.&G(1?fC(,2IZW_H)/a>X
HWU6CQDH1NR=]=80\c?)>NAXKa#)Y7RTV@@E;f,4,6LT;9/AD,-PFMW>GR^8H(&@
)[]66+UP^S^&G0fgS7B+LUNUNdfU5_5X,,BgUd,;&)UJU3)4UGHR]_X&EAc\Q0g2
ZM]Z8&e(GHK^()6AO>(#UTaT<-aS/TO_2_fIf^4FEK_cDZ43ORINK,5+P,>WI(:<
1J?SIZSeOQ89-0M&]7?,6g+FL7E-.4EQGJ63/XIbZ-841?\Nd:#[D<cdOZ+E6N(#
+2-O4./D=M#@[S1+Bf[WW+>9d(G.aNP/=SgCf@g^I^D474gd.(P8BE9+[05?IQa_
NNd5a?W.0X/Fb8cBce3XK3LV&(a)HZaS@H4A^O5XF7<4#b/O7:5H,AYTQ0Wa1Oaa
VMLXBe[<\N-B#5<.gbOYc;HHW>T^&Td;\PRDV@cXMY(1==\OMFG&0BTfB>@Va^CI
OC\7(=^ZP4d]B.\1YY5U,@Ug:5=)2Qe#VUIR],N^36MMU&28PGI+@&G:_,N@.ec(
/:d14;YK5fWMaR3M4B3NG,7_R&7GP,eGK,OM)?#A#K2-V)^Kd-H\@A8adZMK.IQR
6aR/V@>[/D#-28=4bfG=TQL3M86(2V#Q(aLd;A4810SUCE7MGXMOOEMAKgP95,2(
HF6\YDVUA=CXc^)0,PedE_XG-QP1/5fE0HW<cgM,S:9=YIUIQMaNdJL#+.O-.=/S
JYURH552aD?1&M(J&G)P:FI7;G8VRA:^IdF<^V:P[ZKdY9dYK.L78;9I?Z4KDC)<
;7f6/J;BO?<[[6E8R?.4,0&-@MZ[Y(6F9T1./<98a&BVI?^ZEW]XR2(ISOAZ;@T0
BIV[ZKP^e\.L2X]fW@-fGB@M7L-[@1]=18A-[0NQJ;3^;4-S6X)K/;IVU.-=>5H;
EcGZ&)/1E?EUU4Vca3DPPfe0==g=?cIVT@7/e+b6I=8-Ie6K63:4Z)5I6^N>N7<f
8V]V_FG\FCA8BZF/3PLT-aFLaV3>7DRE&NNBaE](ff9EFY.#L6,R=^#C^ZYS2U[8
#V/[_0:)bED+>b89E&PL&:eID^]KcbI06T2TU)FS5-)8bb+cY)[\+Ud9/#VR_OD)
--C;8XE/&dG[H/?V7TP\BW+\;[g:EG,9S,.5TYIae^@JKP&ZP7KFKF6,g@A>A,5G
?K;DC;(L,deaT]31ZQ0SLTPgGMHE\[begA4+:e8(>KLZ3FW,0aXD;Zd;&0eT8H=H
RH&@][2V^,UOVU1N6@,XE/G6@+2EUP9J^4[aQd#KEgM.U,<UF7)Oa4f(_Z3A)B#U
-\#WSWa:?X3S8\QAHDJ^#BZ3J7.Ed7&7H+Se-POO_R^::JJCCZYQKb^N^/C+?2YM
4E^3WJNaPA6YeRGaH+LdCB9V[G8?25fNS9>b9K5MgXa43=e.\#+K=57SDa9?<3^O
>P-4LP<M]K<KO7b2:;C-80Ng)R1^U/?JQb-T4,f+[&HCB15EUdT^-JLSTN_1924D
ZYSG3ML+CR@OG_,,F5:=##:P>KV2Ld;;gD>cgEVZ(8.[^^Y;(5+.g,S.)6HG:-d)
F6;]ed:17@dg=+Q0&/([X=IVQC:B=gV6MH?a_OEK1B,:)</f4>4);O8d>J6<I+<D
?4A^N-e<?S[I<<#T[(-M&AS:LSeXe@ggJ@#/HUM96^-/N,:ebCRIE14Ab11J:gFE
4OLTE(MEK9\4aFH+a(_T&Vg(=8&Z:P8QN(?ag2[^69e1E3(44WZe)\4)AacKHR+Z
1K0->^Ebg>R7?>NJVbY3/KZ\7I1W-a9T4-J+=GQH(?,gV\cN@&)M-VFCQ7fH;TcO
L?+8/T]ZPVef;.7WU-T/Pd-b=5L-c\(OV])Z3Y=g@^L0)]Pc&9YbKI#V7ZFDL+g8
NQK+\48?3L19dD@,V>ND&+0S-+b:c/M>_If&I+8YGc_M)\W+30X(d(b2R2/VdAPV
X&QB3)1_8(7Q2O7G+KB(]&V1LB@0VQE[N0&9FL^TG#U<15]D/2<-b#53.-WEM\e2
OI@F;-AN6P?9CK^(W0bgNCO(\bNX=N^O_>@EIBT^NSJgS7<O>[GO:XM0]Cf,6AM2
dB#KETP5e&.QA73?BQ5;be^@HFQ&Z+&LK?V4.bZIK]NY8V(2,RP2b3,7I+CCdDeQ
JSJ&ZgTROFNAC^&6X:Z\,Q+?f.6JUEg/A3Q-]4+CTeQ&_6S:ZAN6RTQ:4&6UfdW@
fEN@++FYgcYAOAYS/1Q-Z&W4VQ89a@85Xa]gU4M]GFFdE[fTW#B\Z3GD=YYDI7VR
6=P&&F6Le.bFfa6;F23CUe1XdV.OZaU8bY9TA]^(aBVPC<,PA>^3Gb96<SgW7^^D
4[@>d,32@[:>60?1d/R?IZBSTO@_Q\&>J8O#a.6O1+Gd32I,fRINP)?/+;T/])#H
?.^L?.^:U8]T]U;beW9#55/68c+;@>=,&/1D.6MO=L3S@Z>-1LLeV#RB/aP<W8NG
XF,&YRg6g+EU]af==&fIfMD/-a2bcJ#QQQI;(14W^X.fV1a=^)bCbbO0ZV4g)[2:
ZA?CO5;WZGO:KECZSMM3AdG8^]78>L6+.>,N5DI.H^-\]8cL#1??gTPgAD<HXea5
.LJ\J?2T,BRQ[eb/UR)6DbCd@PgVN[<-\JRJ2W=76<BaZ[9g7/F4.b-L4F=ZHKaX
7_;cO5:X/dIaE.X:K]@0J3@;IO0#VLI-/<QSP\)]Pe/b9F:1)D))>g<IY_)U;-@K
\2DJ7>H:HNeNEcKe-_WONM)^1[PD[_e/_;b+(;S_C629JZg-cK/A?0/;QGL_M&=G
B5^8^I?7g?.D3.VB_JaI,3X\[bbc&gPP^1X_,0MG:7fN+-QULUB4BSFAcV<MB/YV
L/3;&R^;FU&PgDFTHAReUMe@:T7QdP,#SCRCeQ6>>3XL/=HK\CFE<<d,V[#0Jg>^
8c2<F-H0d]VN&E4G_3Y4Lef]BT?-81a4)DT]bCXE[>AX)2Zb\7;\d;]5BE/=fGBc
>JdbZ<J[gf/Y^2:56:0KJ\V/D\BHTX5?M0Pe<ZJ6I<_?JAIa>KI3e^M57^E;AB#J
R<5JZW=^^92^NBA8g/&Y^F5L]W<9\RWgdC&,:CTSZ1dFR4ZR?,4CCVU7,Ha0CFB/
[><,V#PWa\\^KTBL8X9L@f(7aVgeJ\\O/@,eKaN+ga0CbWFQ9(#\N::[P&GKd.fV
6YB6E@<a>Q::3=5T_Rg1afWHD,GM)<Nc\VXK_3+N#Dd/f:?6BQ+HBE+Ha^=S;cL2
833)0<IUG4J&\ae;K@b/1206L+T(I_S)Q=bedBQIeD2b\3aK&IWJ^AFYZ\(H&d8M
KggdHM2FVR5^ALW6]FK=ZL:Ze>eDAU76+=A>QbZX(I/bA1b-T?8C\]IOS,eg]Gb;
S_H9W<0-5_Q\Va5OU#=7PU^XB0S_OBKe5WfA.e058(^461^M2=>@A\.RbCKM^I78
Q;.BKN98/W5ETcM(/YT&b\DF5W1<U&2VA#F0WX<+//:/2C-JR;g9_Z8c;JeMWVdL
)ET(Z26SD#V:Z?Ya[5.&J?^8>bCR8Y4&3dCbAH-9?I[4cU_1T]FJS<V1RLJcW:dF
6Z1a<ab5<Sd2#B5+S1fdE+\CcAIEaU\]-_Z:.0b7V,[T09X(K=(H)WJfW<e6^UN@
b7+W2E>^4d=ZZPQNR682g](LEgZ-/:M;EOad/@Ma;e@@5MAXD&9/][-52^7FcK-<
-aH94_Af4+FRL+;8+G:ETLN7#b/NN90gP>YPJ[,LQB;#QK.ab8?]/]T]=,e]Pc^N
bT#=,RHCaZXNBKU#<@X2gTPAeTT]0/6GH.\8Y^CDZW@T@A>HRR1H4^SA?>AK9OVb
(+&.SbBT432?2UZGW^G4/b^>0[6C>eR(.]GE+)-\@+Y]?D^b;bLK4QdNJ7<bd.aY
,fHU?ZIKGUSD0S@DC5QK6e/]BQ8gH5-;0A&2\GF1b@gR)>Ob2Ld4M1G=4f;d+R^P
GH(<1K1M2R^75]OG2d9<c1]Z<IDc&<SE?&,/A-0LMQO]5J(^9X=BG<)eeFJQPU3L
O(bZV_L_K9MWcCPfVQ-\KACF],L&]-SJ>F7&+KZ)7cOU>g_ITb+BIF]Ia#a90\Q.
(-AFEW^)<)M1bL0S+7/ef:gg/^HMB4?e3YRg24L)TJR<gGI\Yb4?B];3YN\aa<;(
7Y7c=Vf-aJg)=\9)eHD+G_(^C58b@R2_M:C63d@_U3_X-g4L^[N0f-IRM5#aW::Y
\;R@/a?cOUS/]QN7gAf.,-64RJJOJIR_SG_RZ3[Qd\;8fbA@972D?4YN<b?]&?T2
48ATHA.I&1>^d+)EdGbTd.M]45QQN,)b.K0:;=T97E,@PgfFfK<M_(CKI4V3^_76
G:c731Za/20@7VaHV:<N9DK<MXcAHKE.-5HV\/#>-VG]]^3,YLZ[dP0YS^,VG.B[
;YC_&#/O<)-UbRY0C>##0#I5F5J65(DRI_=;8I77CV=B4-(cX9P&QAPYD6Z>d&=L
./dW#\PN\gfX8ece?b3V.3P(S+2<Y+e@2>/=P,JT8dMXRN;/L,H/>E?E/?>;B0N]
TBbN>X;AbRQF;&Zc.Sfc_BBE^I(ZA7^LE#DS.B0<+8BE:>B>MR54MV)<SLa9;,;M
;M9Td.8\>aTe_A.W^>6>+<YX:=I[@(f.0COS()U.39_faH@/FOM;/&T,dMPTL)8c
O2Q?_.TUX,+^<@9/A#I0Qa0=O(+7P>0>R+efSHI4^DT#[5_6/@V6ILZ<fZ<8/Y-V
XX/>?S[1JXcd/S2fRP=:)AeXeC9#E]=@N^[1T?VH9D.:EZ#a5SV+A]^_9X?87KU0
(C0?^;.U6<70=JXOH?5].S:]M3d>9Jbca;0/T8D;ga[_e9#:W/+CfU]?#=e<#:=T
N0<JPBc1\=Cg^((g3caLDPY@98WH]K6ec)<[0(^,[QN^T#-GX2OR<N6]UWeaDcV&
N1QZE2bc7H>8c3c&J7R>:O=P&7<1W2Ga.R79@>&+_)e@DO0JBMc/?WJ)&ZO8A260
Y240@eBJF_baUYbCMHcXAJe;.Ja)U6-XO.R>1IZ6URRgX(d+Q;-gdN&Q_BXZGMeA
@UUF0YU<U/UGf8:3-G1gcL\<bVMI79H&<dfQS7N;I)5dTaV)SgHYLd96+])VgQI^
gX4X;X57f)U0^_.U@>Pb;f(a1.;USZ=RN+P=V7S\<-]Se98;NCLF..YTD4C2MeC^
Qf?a?#C6DaH1JE\Efd)V2;C^86;)dMVQ5+1./58M^Q1cDO?=/5=d(,1715ga+Mf,
Z+P7Re,NMe6gdF)MACVJ^)?.K-:B.9)JG5D)<QQS^+3?a\fMGCCT<V-S(\:b4)9J
[5JNJ2L4E8<eW/JL5X[EV2BRQP(f__geg5DUGf4[J4B/ge+V<=Z3/+ZIJd1^\d#^
\:18#e3FLHbNI51_F1QM1&=I#I<>],01YG8F==eb(M^26E-gRN6_A@:;J+bRZPL\
9.AQ2geQBb.^J1.cc30;8PcNQ&3d^./<>)SGM(9?9)>5J&)CT<+4eAa56G<<IU4.
NUT^eIN]J.#;J^QX1<HFF0O+\1).O&8&Z6?/D#V0HE(A<(ZZ]+9\N=-gMFH<Y.<e
?He?bMMc.;eGGY[a)P6/]bXReK?-9-86-A(c(c<7RbQKGe@<g^da74-d(=,9ARAF
VV<]7AC/L\?3LUgVE7GY,YXMY0F,XH\e78Y4)P[3UC<fYQD,&_7Y2:XN<6XfOcI2
ZZ=CC)+.cV=KK-G<-Z-;L_U3/Y1TCDCRA7T=,\J2;<FGT&/VSQL^KSaXAfde3JQD
bgA_CV\]PdFD[P29BASN&\OP>1P?C:Q=aM<3=HPCXX\@LZHB&>U_;-OgDb361=J]
F>4A54;7R(AdL\;eK^T-/fd3NTI9b.<#S-GE-FG(gI=e)FA<]P@Z1\/G5KeS/#ZB
6FV/5FI/E3BeB[A-QYT2^2Z/N=+X]\;6B+e#<C@):D3O>,G1c<+8JS9V6F+JUdT]
PfY95L(BA]QT-=/_7/2EDP]6M6.DA.4E>R?caf,QDORPIS66H(Yb3SBAL(;_T[.S
/@4G;.+32KLJ&00+M4cK9RP+S3ZQ9G<HabW2Xa[dJPEf\D3=b+f-f.A>F7bX>R;2
ICdb5B#^)CdQKO/B#GOTCTXBK&bR=;+EGKG.Ggc\NWH>Y/?<;G5=QZ>aYAB_=:85
(H=G4Ud70SU#4g0d3ab+@;&I,W+TV0XAB>PK?4R6\9Z2#QR_gPGTN13&g[0>PZc8
bD1DR>UJ2&YS?&b[6]F;G.#[;YA+aVMY?]1eFHXaXfJSYU1c0b_e=cUc1B2S:PG&
W,,XP78^QLSUMd@+//;9>;QYD&EERbNRS6(I];08XU@b.M-e77SS]88,B+#:\DDT
#22F5WF-Q<)4c^N/-Q<g@3Bg4EP.Hg3\8LU86W3NT76Xd5&)HE5+\_+@IRD/VFDL
QVN-(TL.#3@Y&8&GH4-R?JObHOJg7A]]3;<Pd<K:BG[69],b),fC3e.SgO(&E0-_
98.^0gYB03_1L3ODC^=&MK&:Ifb7A)GG_LFNaVB<QNdKea[Kd.ASI_@].<c)eBV?
;QVG\;EJK@dFHW;8?B@#RbDISKHT^e:G&3d>4X6,:GX:_E3UV)PcA1N;V&1&aX6@
R9_-N:G+2Kd)CUQ[H7K&Ld\4Z@,Ha2D#=QSI[R9S[REQaW24P>aDN??@JJ;;-LJO
dEMLCBB-A)C9TYA;JL0caf5TSQX=9/PfN=SXVO+GOcI&(8ZP,&D;AW5)>0/[b<N,
UV9B?FT9AUc:a8(QG6O4A;bOIP3LNC.c2QR-NH:bQZGPUb8_C-:)gaW64Q7gW.BP
O2f_^1Ae&I9E)g1@eW_(d@a[S7gKF6[Y4B9)\/^F:ZP#[.?Sc>;Cb<Ja[)N=DPEQ
g[J)c;.PZS0fJ5SSQ(S9?Z^dLEfbZD9>RdggDX&6P=#Ac50-:W,52fW.A7E?3.03
3;S87Ag]T,g0cR452DGKdQ;G0AY>P_RVa?85JF1G7gET^K&a.YQ[T+I>C=K^NbLI
9ULB_?2XNN8A_]J0I(#R>C2=Db7V<78-aMaNM>J+=P[NK^_W:b7S/VL/.P2MXF2Z
YYH3O\0L60V0@_[Q8V,T=#<a&B;J-Z);f0MJQdZa.G1Fd11cgbHA;)-=^gfF,?:\
K\#d+)XI[EGgU&P[]D;F^J6O]B@YDDG_05;89ALK4>>2:;<AI>A5MdRX/]L=73b<
f-(NF3NQfKG\\O#/WOYZeF&b_IR^PV@9+>D0TN9I)K5(<G3S9<R,<P:#?&;[eKDC
0D968.ND7aKR3+ZcdSN\;,[S=LOERP8W39<ZaH]^:OIK4eI-I-_>KbgW<eb0X(QH
(M<g9#RK7H^R-$
`endprotected


/**
  * Defines a range of address region identified by a starting 
  * address(start_addr) and end address(end_addr). 
  */

class svt_axi_slave_addr_range extends `SVT_DATA_TYPE; 

  /** @cond PRIVATE */
  /**
    * Starting address of address range.
    *
    */
  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0]   start_addr;

  /**
    * Ending address of address range.
    */
  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0]   end_addr;

  /**
    * TDEST associated with a slave
    * Applicable for a slave that is configured as a stream
    * interface (svt_axi_port_configuration::axi_interface_type is AXI4_STREAM)
    */
  bit [`SVT_AXI_MAX_TDEST_WIDTH-1:0] tdest;

  /**
    * The slave to which this address is associated.
    * <b>min val:</b> 1
    * <b>max val:</b> \`SVT_AXI_MAX_NUM_SLAVES
    */
  int                                slv_idx;

  /**
    * Attributes associated with current address range.
    * [0] = Indicates secured address range where only secured transaction can get access, if set to '1'
    * [\`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH:0] = RESERVED, should be set to '0'
    *
    * NOTE: This attribute gets set through /#set_addr_range() task as shown below-
    *       set_addr_range(<start_addr>,<end_addr>,<addres_attribute, ex: secured>)
    */
  bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attribute = 0;

  /**
    * If this address range overlaps with another slave and if
    * allow_slaves_with_overlapping_addr is set in
    * svt_axi_system_configuration, it is specified in this array. User need
    * not specify it explicitly, this is set when the set_addr_range of the
    * svt_axi_system_configuration is called and an overlapping address is
    * detected.
    */
  int                                overlapped_addr_slave_ports[];
 
  /** Region map for the slave components */
  svt_axi_slave_region_range region_ranges[];
  /** @endcond */

  `ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
   extern function new (string name = "svt_axi_slave_addr_range");
  `elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
   extern function new (string name = "svt_axi_slave_addr_range");
`else
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param log Instance name of the log. 
    */
`svt_vmm_data_new(svt_axi_slave_addr_range)
  extern function new (vmm_log log = null);
`endif

  /** 
   * Set the region range for a specified slave within the specified address range. 
   * @param region_id           Region Id for the specified address range.
   * - Min value: 0
   * - Max value: 15
   * .
   * @param start_addr_region   Start address for the region
   * @param end_addr_region     End address for the region
   * @param rtype               Region type of the specified region. Please refer to #svt_axi_slave_region_range::svt_axi_region_type_enum for allowed values.
   */
 extern function void set_region_range(bit[`SVT_AXI_REGION_WIDTH-1:0] region_id, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr_region, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr_region, svt_axi_slave_region_range::svt_axi_region_type_enum rtype, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attribute=0);
  /*
   * Checks if the given address is within the address range
   * as defined by #start_addr and #end_addr of this class.
   * Returns 1 when chk_addr is within range, otherwise returns 0.
   * @param chk_addr Address to be checked. 
   */
  //extern function integer is_in_range(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] chk_addr);

  /*
   * Checks if the address range of this class overlaps with the 
   * address range as specified by start_addr and end_addr 
   * provided by the function.
   * The function returns 1 if the addresses overlap. 
   * Otherwise it returns 0.
   * @param start_addr Start address to be checked.
   * @param end_addr   End address to be checked
   */
  // extern function integer is_overlap(
  //  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr);
    
  /*
   * Checks if the start and end address matches the member 
   * value of start_addr and end_addr. 
   * Returns 1 for a match, zero if there is no match.
   * @param start_addr Start address to be checked.
   * @param end_addr   End address to be checked
   */
  // extern function integer is_match(
  //  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr);

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object used for logging.
   */
  extern function string get_mcd_class_name ();
  //----------------------------------------------------------------------------

  /** @cond PRIVATE */
  /**
    * Checks if the address range of this instance is specified as the address range 
    * of the given slave port. 
    * @param port_id The slave port number 
    * @return Returns 1 if the address range of this instance matches with that of port_id,
    *         else returns 0.
    */
  extern function bit is_slave_in_range(int port_id);

  /**
    * Returns a string with all the slave ports which have the address range of this 
    * instance
    */
  extern function string get_slave_ports_str();
  /** @endcond */

  //----------------------------------------------------------------------------


`ifdef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);

  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif

  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);

  //----------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of
    * this class.
    */

  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */

// ---------------------------------------------------------------------------
  extern virtual function svt_pattern do_allocate_pattern();


  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************

  `svt_data_member_begin(svt_axi_slave_addr_range)
     `svt_field_array_object(region_ranges ,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
  `svt_data_member_end(svt_axi_slave_addr_range)

endclass

// -----------------------------------------------------------------------------
/** 
System Configuration Class Utility methods definition.
*/

`protected
c4#>&>R7=1LFJ7#+IbKXA8@>4L3L2d+O\J=9ZY?2P:PfW#N?TbdJ&),I+cf,KS6C
\5S/SR4O8A+[VWW8>>52-(@^LCU(VA7@BH)RQ:#M,9Q+BF]G..42CB@NP/LDg1E?
1A.TV9P8J2fT-_P9[8^@?3cF@Cd]HY]CVW7EaU#d-QMCC>KPJ^W?)08[7XDL>IPg
<S0U4=b-8_IPX&G3?\DH#[W(#bT4TV(,bMb(N@Sb+<MQV7^^#V#B.I+05,ZO]XZc
dgCGYZY&7.cJQ7_gW).#.OX.^RS?C\55Vd,&L-H<F4#^#5.C^>_[I=Sb?RC1&YW_
UD+HDJ0Q7#^]Y=5Tcd+d1FH#4X927/#<SUe:d\cU:Y+4.gXIG1/a5(a.\B9;Y63.
dMYET\cDSZ]bcgPdG^3R-V8QD\SDPWX<NgE:bS?^g;FWXX5cJ&K?GAM^I2<J2\#V
McEH@<.GYKTacf/(#VbTKEZ>V^VNI/&DF=b@?83:<>9cBOGQcN=7/d_=)/,#)=##
&&@&9YH:GCKBB3e>5&@UOY1C89B60He&b;;/_@g8-8ffdCHR8JfEQGQ)bJCPGX_7
6Gbf-16>ZGI#,<QH:B/?ZT/\=?0&;V:E\^L\XHJ9BM(W[cT-7AA,OAWXP3?S^PaT
YMdfS3]D:e88I84:QeQcKgbX5/7UB9U?33)5fLV8b0GWA$
`endprotected


//vcs_vip_protect
`protected
S#JgHFLWc#IeFD(<<N;298V7C:/+)eg/FFa-JIM:<e7[d-]<BUTT6(Xg\D?:bNOf
Z_R3W/#+g;DK26-g>C4E)BW/6@>Q6[eA/869#=gX=g/MM8J2Wd4ea)Q1Hf>EO(+-
9cMR::[bU?-Y82dR[BGF#BNAP8.F(L5O7Be+Y#.;B6H]-3CSG0(<d_[LF[=V6.Q>
30IXa@&J+>)9b,,K7B8.K=01/KA&8aB7<CG4.6MW@+C]&^#=-^2UP_FDAZbgS@Zc
6X@9MI.AX7g6-d[@BSe5=)@5H2MPQ,&QN]dD@E&e;P.ABcO7U/Q^/TL->5-K0SW4
W;6cO,_U\:224;=F/B#f7bb@JL?K:Z</aH&&X.ABgF>GZ6)fd,+Eg@]?08bE-,90
34+=F5JH0\e<Dec16f#F^UV3NWK)CRU^DeT987F,@^PagELKXMFQ,DH9f:aN,c3W
K@)&,AL9D4?,LUf?V442EbHOZLDBB8TLXcP0=XJ.,e(X^db)E_MR92aD5PJL6B<e
V\F)PEU<.7GR2NAIJR3-I_8F,PPQT>ZAV?b^(R;2[=;eV9T[YGa(4ePMB#g7E7SZ
WUG(SbO1.429=\.=SQL1_/WBSGT01)R5ZBC@cNL.5NL_VFAV-J\DKE,K4__HLKVg
/H4)RW[(DSE44/Jg>/@JN3V03>3;:B6U1Z\BJO[Vb0X618\&5Y/a<;]<R_C0D+Ad
E[(Z)F0BN4)5MgaZY/C?3XP>acS5?;LBc8#b6BQ0O(6b>d_ZXR.(,7LZaFQ#Gb\?
3?DagI)B[):]b30fNd6e2Z02_DR[8&[EHfVLO=WbRA^>8XQX.f[1c:)d2OA+CM,U
&G1VTXTG14]UL(B.R(+J6BK==ggNEX1IgZ6N4C90IW<K,(6\T^VEMU+?5e\/Y&JD
N2+BI[^ef[aOSH@L=#Q4[3=9)#+;Q6/QUB3Ze6=^^X@L@K^]ON,1#P,77?YP+6BD
@9fO45]A,TM9XP()#)6L@<LV91MU#\\3b>^d9E=K>S@&_ea9V?Wg.^g/5QG;Y-Qg
74XY[E]F+SX4g5>[NSOFQ(fdeF?Kb@#cLLS#_JLQFB+W^2gJ\WcRMXFV&YTU>9P.
.>J].HN2H?WeG_]+0Gd/9bBT,NBZ45==K4BeCgCRS>+gLWN0-C,E?158&\UcH\R7
/]\6+VBeA)^d01G587dZfa-OM4^<);P<FbFZ8B;d:M#49]EgC2g1/2)a&,BF.aTX
#P\LZ4;\M6=c:_Y^Ab=K@WE2AZd:=]IP+=gRTbL](b\=AA-CSXWA&Te0ID_SA2?_
DH?S;2RB\8eB8Q5L#d3<U-HACMFR@O>AF;fD8D83NO1NF^2B_CfbBS@fA\^])3/0
EN&91-1(b<-I;.EW[^a>.;FQgWC6-Xc9X?<Z2A3YNcSY;B^ZS,L)A;\QWcD/UH(f
>,A6N/8D]e\8U(BL(f5I3XH/;HH1=Z+2?J.Y1bN>EAY0,=N,>SIVU\_ZGGJg;VAY
EO1)/8Z^4E)>ZQF5S<]65.9J^eO_?A2,:6.=COK_>ZM>E7V>TL40JN]1L7#B//<P
Q4GY-aGJIE2Eg3T46\RdLSJY9].?U,,?P4^@FTd,L3YS]E-)E_,GEac&A.[J0G\9
:+TBZO@VW?O_.(2?c74(IUU[BaCAD=J)F:JP;dP[dLK6\K>-^g<H^f&TY5JK7J^X
3,8)[57.-;A:G:(@c=<Q_e<Q)I\eAFg=01_d9K2NLR3adPQefDfZ72<=D_8@,56+
]X+Ra4M\gP8Q\DSXW8UR>C<5JVBf3D66HdOE2HM8-_A&6017&SY(,=bd)Z\d?[J9
DV,.YLE.<Maf41-X0N:_X[;H_C+>C[+d)8eee_G:.W^\U=FUAN^]8Fg-VQ>/9Me0
VB=(:72,He41=,/=0LG>#B.L:eVF-e5bAVJZMTWI_Y\9d#NaK4:dOTDBUc4+2A14
YQXN4_c>d^K[PfB9]>^IIc-<]e-OaED\A]gL8_>1BYcXM,-7Ac_WPEUDG&6/H^e8
b;EXV;(EdeWOY+147P3IDCc3^(JO;,2^XGZ=F/;MVSG.;e-V.C_],R50)9>FFXCP
5QL)]0_YBGTD3,2Vfe77^2L=75]RHc4@/-<S67EL],ZO;cFCH^E.,[>3d@B?d5R>
LOeQ@AA\T1GAbCD,A#9dC6T/)];gB>A1/K>_9]AHP@eSg_H7dMG]GDb.eb#D+Z?a
@=5UB?T576^6C5d)J)=Wc0LbW+)#HGI,0;MWCd,,#0:<Z&VG=c4Z7&1MTH_XA?+1
-6P2RSLGJXR:PI11I.F8CO\a/)V?/[1SV&;X(<12:Q.C=G[UFI_S0DdCG#^S_EPO
OA45Xg/>RR:E@;)]WSeYBf.2XA4Z01HUW(KTX__INCN<UVb1G^HNbQaG]V9OS:]T
3/C)dL_]A^e)OgS5I@TdO+@@,[/SH0A/R->6+Ib;I+=HBV(gA;?Y\L_C[KGE^6\E
gSI/@_[c6C@[>;]eUY-(;=Xdb_A3,1,(0X22^P#ac29gM45?&G.[5S)JD^FdN>dO
Wd-46\64f6d1^/-/>d)&9DICgF;.,@/eE+/964H>5>9@]-BY3GEMDJCR_48^8g6L
MbOZ7Q&@g=4+UI;JSCNT?HMMeQa\=:cK)K-Rf[N0^;5^aBc7/A]+_52DA#WV#\cT
[889N[La/8QK=5(;9:7b.>XbI@JP^AFYT+]c)J==OcHC96G\#+=I43Rc2H33J@g1
Q;Xa<^RC2c]MXQ_S;g32WZ6]/_7^_BS))6eX<5Z7\g_<aIQdbM+LN.(1YeGU\f)V
[5\LR-M=9B);[)Z(HdKF->@CM8LeCeOM)TE0b]6NYcR\RJ.fYXTI[dYaHb<QJKgg
4eb53TFCSCX_Tbd,UgRb2[+)JJ57QOKPX)OL[[?O8b107G.AX+B421S#G[QV7;MO
NVD)EY89W>ca,NH@7SW^H7fW+IC2V#R3(6PB+(55O4@TRS45VG;OVT?9GcE9.8/g
UC#3)WXc=dI5[UO(MU1ffcBdCA3S,=_=a+F0:,a3Jd9&[aDg8FEXKS?6\RLXUPg?
K.CD0;+-.?TP1-_SP5+VB].RQ#=RgFG>-UgPggAE7C4B1[Vb\U(\6:5-(^+eR0Va
5O=FT3XKT=A.PNfWEF+\HX@7\WNaa)5)#(Vf5^>;WBc3(8eI,6T.B\&1(X8I&4::
07F4-;NU^7G()0Z;,5778&6PZ8Y&WXK=Y]f=fQ73BNZO80<.^QQ,>MJN2\4,@7;U
cK=^b2AHS,>G_.E/0V[[KDK#_T3LgCbS(WJ,-ZT0;g02[@O;<LH9PNDA(CcMd23b
/UHT<AJKU3Ib\8BEZe,YHZ>-FZ<&2)2_\YRdMUES@,\MGfM;S(^a/)d03f^dPK/V
3^bd?P?Q4R??W3@Oda(ZU_fSa8#)Q#X>cD<L87F>PDLTTf:,g2^1[).FU5BVg,1\
NX\P),,=VMJ^N;FbS&eHeC\</BK_[SF=fbeTeP5^fc]C7WF&[T2KHM&6NH=47<d^
BZRTQ&AO&\.^NA?;LQ7X3=WTgC[c6,bKb9JN75,3&gHPVa.MX?7U+Je4dOHW9>;H
5PRHWDB=VE):=HHbPdW3R(TCIU<TB4@b<b<8=5_e+3fR^>#=/W^G-2B>Z.-N=:M3
=(]NB<E(=f^c?6P6RAD1Ma0LNFNRN&.SS?C:1_,fT:,U-G-^(>\<R#^0>1&HEHKO
MMCFKN#MZP5\QOX0F1IX<4L^0aM].SH[:.2A:H\G@Z4[4@[QW9HRED]WfacKBcPc
J[3UMRX0@c2F<>TVXBG:=0>I@JB-UNW&^F/0.LE=.EZ>KIg58ECHD1EX?5Dc)[7B
-9,=EU(:J8WC2b74>N:UJdV@d_1OdOV7D.7)>#Q6LS.e,5+DW_Sb<2GL:]/128Nf
[JcEB:cUM@;MB57#YDJLdgCNB_e,X03O@QS?bXY^6N_@WT;](C?@&e1(@8SD=+<U
7XF2BgB2&c]R3WQP6QKNJYUZJ_UE4-bdGfJTd:GH3QI39?d:R3BS6N4dYf_>A\#.
V[K\0ge?2.ed),eV),Lb+US(9Ud/3T.@&0L,JS749-M(_^[GDgRfP^?3>_]Q]SBA
#FS/P-P1H-O])e>-fBaRJC<;HfFBL4F?g.f^=\?(+c2)]EKfU9NM+1Y=SXFZ+A+b
LRFSEQgA+ZbS@9Fc[DLPcX7>III/FDcLfER]D.U?4Rb]T[@K=(XPfg.PCWY^5#I=
8V[^F]PBQ.EL_KC6.MVJT_<^O@aQX8^dO1INK[6ZT=QM^G?9eV.Bgf.U44_\8KPJ
L]>=BK)LG9PQ,NZO+YD)<EE=[RM]KaDED^MRB;1ZB1N.MMc_8/>L.B)@4D8&/6X)
+E)\)G7e6dYKD6GZ1JQ0/[Y_1/Q0H;?+2a11e.G1[>C)KQ8FDSIR<4^:.a[KaZ9Q
OKPB6BYFVD_1\]M1.&;0VUT?\SGKL,D:>7=ESJA1=-7>H14.C59AX^f9&(#:+9(1
cKc^3a9+O_J?C)(8b[RTgE0::OT?1P12G;&YD..S-]MfM&YUB[EMD_DHJ=W9Qg3D
.DMMMd:HEAAdU2:g)+ZIR\Qa9]8_7DH9;[;FHf?90cDC^(3Ud)<cMO:Hee3ggSOG
4;\5@B,_4@EbYNQ0_a[-YT^eR@X.6a:9Q#\TQY810,a0=g1.f.9=faYE/9.E8AN;
RK35OBe/?)Y:aJ)1G0K(8ETQW@+\#:EG[;\ER,;Y;R1ED63;81DZ.KH1F]YF4X&E
N=_2S#_==d5VF]M?EMYK=:gGWS(ER^Z:c6(?-HR;K\MEN,SH6:7J=H&Db4BN5\E8
4,L5<91/__gSc5[3g&FF_M&+.W\CHA>,fHFU6QMA1LCdI7NRRIW3>^JMA/OLB<c+
PFWBf.eISc9Ud_>][(>;I<)+RE3\ZW9Qbe<4_8#C2VQGQ#8K>(dU-#d=P/QOPQ#W
]H#DJ>?#=YSE1R4,c]4RL3[YX00XCV]b9<O4C=-9?7(/2/3V]+;/E)\;gaEg<_,9
J9Ff](/T9TUY;A42EQAUBVAc[Ad+aKZHJRB\DE2.MY(I1P\RO@\IN4<VF>0IKTF1
b&BOeeAG4374GH9YX?W:D/Ld)FC1&BgU1=dU5C0Aa9N=3931>RP2?^G]e9A0]IJ@
?dAI5<2^efJD:QR#)H?bP_>K?73PL/Eg^J67(dKVUeZQ81Gc.EeUY;&[8E#-;.GV
?>@E>U9<482e5/QFO-<-a=<JXARf<C+0f;(geB-V.HWP#VXK?MCF)eT?VYF#d&]6
1?O0.#dBD\(&OCbPP:1JW=eKQN;);DG^ML:^c.N(+_.1C5ZW4^KWb4&<N9J0a(RC
G\4A&F@GY7-2PfAO>;a<_dTKWS2/G&L&7G<962aF<Q9HM;8W]gT3;L<b9f^YGN;=
bdab@>4.\VD#<)5f#Y7O;GP9SRM^1<8S\TE@[;E^XJXC-^0,O9+c]9O._R3XRZL8
]&,TR(dRX)(:OMReW;bJN(^]3F8)DR80F.5D,P4PZdF@L31]6IUWN3G=N9501B&H
Ug>+4edTHg9;g(IPdL#8+8A?>L@V<,T3B[a^NN>0&4V>:O1R+cLXSHWgb#;S6-IU
@7,:cae.YeO>XWfEa)Y@b/EY8_QTEIA(c.KX[)KTZOX&W/MZ0aNHSWK_-fNGO&K^
X1BTUFUS,<a?HdPed.MM@YAS4g]#M2e-8E86(c&C?U8\DNLKg9e@V.#YCQ)7Q2],
8F?WZ=9F<\#8JdEb4d<TZUYHgBFE\E&94YPP_aE32E]IPT=U@M=L,4U.(Z6]S-9P
3]I?:^.\OOWKE0]EK1g2KXUC/Kg8T59gUE9Vg2Z50,eQ\\Z)N#\GIE3)\DSa3OQS
:2;S]H2fI#5HB1<f8a/g,O@P51V:>/_1+16J&&.73d?gA2g+UBQ&&4,A(5F#5AYV
&;>-Hc5S<JJc8<VOA6M<M4gEPeDXS-])O&=H]@abeFDF.MXD,gV:F3K(c/E;:#7M
WYW802@NEANg^1.@N?0PA\G&W;g@0&1f7?Y=A[M1AEZ,b9g=_cZ_\O/Z3#@eZ5O[
8G_Q=LD.ML1;FMY(dc[R--A0&JQD/C.D0=K;.d(b),QXc^H=e,6985gP2B6I)>?3
0Z3V@9@P^O:,?K&L^>G+2TY0+Y/7+<A_?-=?dADe^d&:4<5XQIAR2A98g5/5YOF8
&\HM4[+;\5dE]MPSbIC0,::>OWH):F>G=LPf)@f\?bJ\IK1+)5L(V#OYE0Y:)Of]
>B9:V#[>^@?:S413N12\IbQYd2aER4>EAcgWQO#KLbFK>=RS7LK)TX),HG2[]-2:
HAD.Y99N#PY/,+0L8+6\ZgXW4N?R=VM3[&d&BPT0PTgCPEV\^PTJ4R]?&,;8dJQE
3-[\T1MG2J08I@3P:UHf[HWefH3RU.;3.[/--I65/f(^P/.JU[PKO:W]Q+,G<9I:
.b?V0\;0<#7fIF@a1;+.D\XWLM(EVS6><@MBcPI<20=U_NN7NfAM5=F;F9O+S)#)
)<=BBGH?@QU;DVW35+NF6B2D7\@g6(CHB6X]5<F)c^dSI(QNI@eSICR:Z>/LAB<-
R;L4cbEY:3(LLe0I,T4;E2PXKIMM0Qd3D(D.3SFX]K_[dBHR<beN<>bH&e47H+Cd
a6FN=T>7#bg49:IM8Eeb>A?_^^&/d&,RK[?-1Yd?gb^7,VC+8T71;d\UKb5L1Q7e
2JA3;C\_=B6S]FK7>>8\L<2aNWD3Z5ePW;UH&0K)KXc>9+9&8BMPONXB4V?<@SOM
N,?L]67#_T,4+=5+X=_8Hc>d.W[+K;cL?cYVNSTV21_SHVXSO-bKf_5Q@FA8ES[5
6D]QUVeCWP5+8R5>F9R7FZ\M.0SNQ/7P:9H\[]7?IY,;]]\I<e1IaAF>ELg+BGB@
:M^-^c6IcWMH;=@bdF5AbeMRS1a\/F^?]X@e8&B_8+522<K-J2ZC.GZgbBWb-&#,
^(96bSXO94Z(Pa2K1?O&)0aI?Y#bSMfFW4H<N)<,XUF#[d\:&>8/La;#)Z3fd4(F
X>H9TJ@KG0>,(BDJBJg5_;DDRHY=H]_J.UL^Ogef@#c:_^fg&GD3QV8<[-a(aYC&
BUB&TSAC=Y]\JCbC=WU.7b:_WWNLV2ZF>-RF;e=]Q@DbPLea\T1=;bZ,:+M&b(^+
N7TUO@@31FNAdB<aZTKffMNcQF/#+<7.S\[3:F;YN<D.O6E,4_TUVEUP,&8K?d1(
M7N4P,.VUf?N44IAYP#@J?[D[Y.C([VO^.6E0F^J/IAVU.&2G>KffYPeKe:8LHgT
aF?g^[5&#KQ:BFIL5+.0VEPI_0V[H_EDHEV&M4?6dN;YIV@eQ/aE<:eRRf,2/.66
-YKc3DC8B2J<:<HSZ?.ILf2LGMDZT#9Ca36XLVU-4\@6#1KO5[>d0^=.C3996O9N
&ee]0:N07ONA1^KCfV1DBQ@O,5)-b4\(F)--:\2WX83XIEI6W863?@M(2YWe9B/I
D1@QP_OXQ>ZZ+b##6aJgS+Y(L[U3d9]Xc2B0&+I+=ff&^6XNe>cT@SDD[c/3df?M
[8)OU1,9N@,ID7\fg]R@VQ+&#5:G4P85TT8=L.L\0fbG@U?[IQa^Ae;9cU7]A\dZ
U<AA)9.JK5&+HZN3_9MH,QI+0.F25ScZ6)?I\;Y4]aH\/D#UN(^b^_/LK:#[f9PV
bB]gMfO1H8W).Z6/D[4&&\YNT&PB_&Pf[#3P\aTK)b,[(YTR-fBH;&eg6#^UQ9]6
.T)fc85Id[7gMVPLJ1@HRX(SVHL&cQ/T]A=U&<.C^E,R;>@@PJ,e>R9Z[g4:VK&D
#@Jdaffe;aT9C,VY<YO<K6-,]HEUfffP.[#=MJZ:Mc0WZM4d_^8=939AG(\&HCRB
T\YPDKBXd)S39ZAHG2^,7A)I:#U/AZQ)?>:OZO\\;AC/-Nd@AUQ64E+#MWLYaE3U
5(^S:3eQ))c+TB)cI2T-QIgN-9,Z]dFc25KR4M,-c9:9;D#QDa6c[&7IU.20@.Td
a+Ec-[.Z?\2Q31?BU=/5H/(.9<RF#Q>dGDM?28Y+;.WGFOL1+[\F3@L_fa.\9-<#
dcY:aG5b,;B84GMZ4Ef&aG0K]SMc=3\Hb_GW7/F[a+0C[bdZ4BPE#?\P8+@gVV<)
e/gFFe9,T^XJaa^:@b+B(Hg5X#PV:Z4K]_\Ec[Za)WTO&=1Z?J:6@aaC<Mf+QQNN
ZH@>ZbaE<(aQ?7I6AKDLPX5Lg5W.O4R+fG2;.7FS+_Ebe+g]Ta:_AYa^H)IT1B17
@R.7DO#BTYBRb))A1,#51[=VJWS.:\fW&SWdK#,X0#Sa9HNL?dN.UXC2E56@UKBZ
AZX8@&HXDZ3.-0MDeA]5TXVM525:YP@=8BLMd>+>(<9.E:.Qg)PJ.;5OI0V.,OY+
Z_W;1KRF6YFFDNW_gCJ(.a/LINSHaVgW^4#V@A<4)MRN8;D87aRI6JW7+1C+\DP+
a9U87-66I<P6.8<>M]CKT4C>a]O_=48aC)M[W=7F?-AB#bEHKdUDB<4fFX3a\Ic^
=\N52XAG2f.gbEa[[L2M^B::I,+HZ:(R#Ma_SCRM9AV,M@<9Bd@8)]W0KGU;KX<D
eKH[VA)FW[8b2Q.\4AeGY3>0VNH)T)CNU0_6H#WZN_<Y2S/X73#C1R/TWgX8Y4.X
bIYRRLcIe.R+<e[2)\P[/R;AK&7^?0O?d.?CL@YM_5J)IG6MJf,O1T[eJ69[#bF#
.[?]UQB_4=;C^6KOLVA_ZfH]ROIBMbS0V?DAW-PY=2^?9YbeBR=^1P+fSE#Q>1&e
c\a&_\#9cTG)YD@LA6]>ML@RVEY4=0@Y9a9(O_UE)>Yc=&?/VGW9,Ua]F<)W?33@
\Y\M8EOM5TX<)d\M&PY0JB_SM.-VE4BJ9#[1eN=4,X<5&]ID+d200Je/,/Qd68VB
a#D,IM5@\Ba[QU+:b@5W,LODIP;79=XI-?&88]+aK1\<^G?R#Z>DdW-KggF[[>)O
K&dd_b@c\[_gFP=<UQQ1IP5Q:CIQMMWWE0Ae3@dS7V&-60@fVM],XN5E&=OK(<3@
,/BC6K2@]@0VNX<0)6B.\G=F&1]<DV9AU3_^S7UX=B&_NUcP92<[7EO^BO<?ERPH
(aEc1>NZT_=W1J.NM/>A2OWP<D)GT1(daeHUg7<]4N?AG>1,;&3R+g)-/-.E=ea)
_#=e9RdS(f@_BL4NM[\J&Ia\F<O.<)/+ZGa:0T5Y8GGc0TG[M\f.H+@HA=FV@)[R
?ZLK+?KI/7_b?US.RPTQ0C0GIR5YZ&H(NKb01D)U;R=-F3JNTFVN<A0<bY5QZY@R
4gU;?QSRf/=/3R<D&HP/SVWRf^dG:eOZc\6f9JL(d7N.<6cJNW4RMN&VaOg3:H_=
G2VJe:5O0.(/#-R\8B?27:>J,LEMQ\C#+7>)2D)DKNeD(?TWFKI/F(6CIL=U&_(K
1DP-V]Q@:NeDeHCNEH5#9AXH.:](XcO8A/AUN6>YZ1A44F6(UIQZH@QI:bUFW]b,
L:,>64H7M1>U<eFW@Z)C#]U^5Od::aaE.<=TY)UTV-+X)a1/E9]6Y^KDRL-XU._N
+8.DZ.R+-&g[EO,IOZ>Z9M(G/@f9>Zg@TQRO-7gHFf.YAK#W:.ecL>L.HdZD0]8J
E74XVL]>E<):S-4?VQYEED23&P6e6+V9UYH:a8^.Z^dXL^#QA7^K047QMSG/X/UH
Jg9DR=G[X]UJ3@a(Y&O7\</AQ<3_&GYJbB3QO:IDT-b_aWgYLB4gZ:fg=a0>UVY^
J-&Y@D<VQD>?U-2N4=Q.-E-QHaQM=#M7B;fD&a61[H,FW=cGXX+240-a\,2ggJTP
JD\aLW]G7([KAc)4>_Pa-)/NI^d[UZ(?ZAPJTHN,fQ:_9<Q;cZZ;P,XC=;Q7G(7-
Hfe+=VF.(P:)CMaf-Y?(2J?P\.Wd=9L[&P<c-CJS#FLR.L2L&.MbX<UT:8&9O2)3
+/e\f_]-J-0VH7=C?fQPG/>_1U3G2O3L.T\7[-<I/Tf70^=E]R?#OS\)H]+@LC3I
:+0@KV(.&B?2JSPX\(JOW;TZ9F,,5ZPac\5HdA4YTT\^;64G8;]^^.d<4&A62c7#
eHZL.BL3H&U[]#IKX7M\J<?BXC)<^TEaZLO51efXPV.H;)7_N8b6ZJ1)U@U2+8J?
e/eI)a.5a:>.f?X@@<5GKc9YBS3YaE?gKEe8(>BHX9\6JDO@CJ2A_9?MIJ3\]:(Q
?SZA3I?DEEQN()=UUMF4L1YPW/5YB,IVZ8bS=YdcIKMc#eL.5U&ISH]R5N,]bKWg
0D5>\EN&:g@W-@3I_^&=5TEHJ1\+3fbZ)E6N]EUd6Lg85:V-8-bJ?\BO52VD^9e@
X#5]()]-3c_&5C+]aII]g56PYV_R&>AS<J>Cf4]&3,Z)0<C=[)A_9.fc3T)>3@=Q
:eH3HWF_ER]O<MOa&M3KJg+9,^A+2TFS[F?]fU52G?b,8)Q/2+B=I?-Q6-YSc#1)
O)&TWgP1RZ7+U2LVEFd2?UGMPAEY8GAU@>W9PJY2(-&e._.g@#3HX>:La;?,0=H0
>>;Tdg0c^WYgT>-:7G(dRD51f#g3X0_KRT7g1&REBabEg,FgcEaV6](@.+0bD^/S
:NS?Yd+Z6MOW9_ZZgLN12OeV(HU2I7#S7[XTDYe\XXAZM3OL1#;&Y/aD&1P>#B\K
BHPNE6F,51:VD)T&8fG^5U^<]]bHH3B+1^[?Oe0XF9bS(Z]cEKF#,]F0_E]#&2Vg
Tb;6J&RXEGfRXOZN.F\(ZB)gg7+(DB^;.VF,7d[4);.01P/=a/;B9e,],B3MGea5
VEFYE--/FX3)_CPVW,[75eV_dJ1/fcWZND+Jg>b/E,5B,OZ2?)K@+9LK:Q5D68SE
M7UR#ZTEfZb+0@=\)98I961Efa7>I-?8@O<6,<],MOZ9;SG@W7YQT182T=/B931F
5VfAd+SdA-\NPGIc68KQQ7/88ZYX[Od2f&+T)0U=c/,R06&6^8<b2N</E(8.V<YP
d6EGg38G.B<[dd#-6CJKPU<P&CeB>QGW_PSN,2ES)U]UJc&):)UZJYg>R)ef^6[N
[gU&[<D,NESZ<fcXcc=.TbW(B_W=QE8UC001HcZ,P@L7gSg5.V3S9>,H1RRX&#@5
75eR@Y-g[FQ[8gLTSEUeT8Mg:a)Z:KW9BL;)U:SG7)Z-@ZSOFOZa[a^e&>f..969
QEGKPCaNK_:?RMKSaU(?0,2>)ARV]=9SP:KW=9&:F;.(:GT7:8Cb0AR#^Mg&+c3;
6Ic]XG]&@FVI<3]RYP.5-e2@0T.2#?5-H+3Y8dZ,2_fHIZV/_-bV9B#f+0&P<+8f
<^Y_N8WC^YT3]bCM3U-H0BU/SX63+V+5AB2DZKT.f8DGOC4XP<X^e4>3f+,#G3K8
fN8TWAVBY00-/S9M4#0;JRO:0\F[SMMI0:+O]O--A,b;gd(PPLK^[9I1SFYI./dM
XTSPdf8[VP&ILX-<O2KZ-8gLJ+a@Qa97a5+ggeRN76;>J8XTK8IEH#^(^LB4@6gY
;Q:NQK/4EWPS)CCH#1-33+?a^B8[BSHcgLJC9[F)=YQ\fbJVDZN14WJT18C,-0T=
+UVH52-X)\7DgM?MH2Z^+#];a)PSN>>PDRF>/U43]Nd>M\4#II]-CMR;#-\W>R0.
Lf+^DM3A2U^A:JE?KB)P_cRVTGX-)1D:VLa)b]B6egX/VY5OIg5:W2UG)ZH;4dG-
c0cQQIK\_Jd2<AdS#T.>8gJTN4e9A#@9.CWU<#B-JR818?]N6V.FI.7@<A)Ca/2N
S9;SPPP;-d0#bIBd]G(aBf^T@ZCZEY[C<DVc;;B7UdD&V@B08W#:aP^H+^1@9)HS
XQZ(9/P\\Q\&1S3e2-R<&cOAD-Q6/HPAE0>]:&WOI9&d(b@0_ObIPXLbNYZK0I40
@X>Mb4;[0=6HaDXZ>OQO>-/IGNJFHWP[/D<E^80>;)_Gf.LC28:]/6,)V])&.)FO
,AFM(GD6-#RC/X^_MKN-+#H-U7Ia6A_#2bd:.g0ZT:IL8c-XROJR15T3A/ZCDTA(
0X9Z1;#CL<dSeMP;A;5Ze][[.@\F@D9/>OZ8_?9TO&4VR)FHI?EB(-?HdYgYW,b-
YfePQV>1S>]\M:\C,W3[08PX?L\^DZDY83?180<^6L3ed9OAc,>9_-[;aF<DA3cJ
Vc<&HG\cEZ)4Je;:_=3X/\(_53--B3R@;COQQ?#>4NGZ):&B._QLLJ&7L>(XQ-6_
O#F(/(UJ&JA5]Q^f_GFDHM_\XE=IG=;9EUb#MeVBW:0E^T-bY,7fC>]6OB?R@JGH
B234@QGIDH/D947@7gS5@f327B<AUTD6;If#,JDG&2QNFMAPH43SGYdX_OY5)-KY
d:CWIMJ/&eXU26JHS55PD#:\GJ3[S\G8Te32U-92XNHSP)WO3SYgdTgD6QMR@9NY
ZYY>3&;((g3RWHO@SH.-&SgYFL2N&=7FV5=Dd:<0\CT#J8a6\YZ:KXT#6CX=cGQV
&#,/IIE:@@eD<&>+&C/gV5,4?Z4:I&W+HL,ad,G=I&KNRV+;,:BQDW^YF0Q&U;7)
<P.^6\C4(gBA:7gC-FF\/e[7<(=XBAY)cJb1B[HF,Y<Pa>6RESM&L4Lg0e;AGXB)
&L#LTN]P6@HQW)b&G/M:=@Y2>N/L@7@O[(X;U)[aV^Z];;a>ZLb#7g;0g/TK1MKG
&05^O3N)a,D&Re?(O;XE0EgP--)JbIVfA_07AY1Rf-971_L+7RGQX8&(=UcT<Oc5
c)e2+ZB-Q<GKdQ-#[/-f5R(+JU>H56+UF;O]dQV7HgAMKT1>ZCHS2#B9@0fT8;,+
HdDcGA]M#ZFD4.0dR[K<D6aUVL<+<E^M1QcSU/@a4>4Rf#g&O[8C1IY/Ig5MIa)A
aZEVeYH0f4I9<@W0fd,N0E6?K^\g6OSE2.FDH^RB1JfCY[D5S3cRM8g?1XK#]R22
^_Q_\BF1AB=Ed,[ZBKWg^Qbc6b3+DegT3=)afL1MEN((>+7LNd5D/A6L\\.);119
>BPPPWc^9>)b&^QZcY@LJJ0+g:]99(D/P]:EgF;gA;K2I;H)>O3=S2^gV(Y63Q-d
HG/Rdb_HD?.L,L/<AeO>Q9PJ5R++aDTfXW_)Df.K,?EU:]#L;CKBV<U[3Y\ES@,\
?,bX\OYX)JC]-Hb@bgfGM(Lc,.,KT(U;Yd4.N]WLN0gX72::fD7J=c8Y;_ZFcES:
2WR\MD5R&(b:7.P,A6_ag)54^ZL3HU6IWa9&@@Sg2A99AfG76T@Q3/R=)^1=+-1R
Z^PL,3.B[+UZXEE\S8RS@ggAgfJRTc1JE0+)I?#0=4^gH\97;E9RgYN3,=66,aFb
SY)Dd3U1<(@J2J7I@TFVcN9<D5E.]:8.M28J8g<LAKcVHIae./E]9T??AK.f?]@^
K(;,c5JQCbXc@f[YeUSFGFVSf4@MdedASL?JP_++UP>-9Pf[Pd9>bA+]&AL-1FD+
:cP\X4ZGcJJM&J-Y,0VJ(KeG;7&B-428D,3C5:Yd@VTZ)A:OSTKJ1N70ZW>=&O,Q
(:NWeB+g?5W/:QKH,F@;@[UP0V<[@.ZL#W9b:=T<F73N>NH>gS<[ec/9=aKP[21=
719TD)L<Lf2.]gG]#MXTY9M8NLb+>M;]T95+gbUWK?O@B1dd;(0](::>0HN]VM8?
T?SU.8]---#Y^]c\[N4:M4&/S:8dEKJZ\]F^L/B5(J>HNT:cLL5)&ADLK[Y(-,EC
(UAPV<TO,1K0@<Y3MOUG6NORB:W/1;d;30B1AA3AEW-;7&SQ55BS0XD6UV9YH3fG
<ER.SC1)P>5f6KgeT;CA;3RL_3)T\F@MYI>03C/6WIc1gE;>IJ+U&J/TKfIB4&<[
VD5b9;VEZATX2TV?B=N/bf17cRVS^ZWYJ[Ie,b5C(7eJ1BA.9/:R\e<[:dC<LJ+H
9U5#^D+_:PP,0V5ZAL#.:W=AHHcY_-_c>)MgF;(5[O))=PQT7-XedGCJL@D4^1,A
Z8K,Z6^V8DD<:F>:g)RH;[1-Ce+W.UZ/G)Zb=LQ?M,60./N;F)L?(3(90,96Qae?
#ZRNK\Pa;PWab@bLc8Y,K2VdRfGKW6HMN;2aN-GD<bObfC@\RLIFaE<>X(B5+^]&
F4fUZ4DJ5X?DIZHJW+2EPIcY=6;,c2BeQD0+A=Ya2LP)GTMDNYS8.I/<_<?DCOO8
SMY663P2W>Zc6.R_dG[^C1=9+I0I5R1==>/=H#J\Z8B.7N,BIKBYODG2VY-D1OOd
bUPD.CV=&\33SgLDA>e<eTYEVTA[faW4E?FD=d6-0RE5U#\e2@?.7@e[)PGKUX5.
b[/J=U)F@TcaUYUJZ/PFEQ8-,VARM\dF1L[J(1N90b5R7,)M54#e]^8gP@]@2YGY
g?^^9XS3[Q0+:-C852MY1YC&[P+c#5L#CBa6C<JF#g4&JDLSL:0+IIf3,Q159Ya)
R^a_4=^dV#=@@:N\C[Z717[M2f]L[ZScIB(cEMC/YH&>T^-,R2G:JX[G105I&3XR
8EJaaC\G+He_M:\Z8G<7J]I-T=4[Z=RFOEL(bT+UH9;T4cbZ9cOC(V_S^83A5++e
O.?g#3edQ::^^JS[FV/9+MKT=(c0UY67NWda21/e3-#Q=HX]Q7F=OL1Y,>_X>[)7
R<F/YLJ.37>?[.c&gKC3@T)Y@36D(_96a,=f7bST=K-=T95.g]L^U0Y0YC3.ZVH\
cV#7=1Z@?-RHNUZ;((#T-fNI03]>fYG4@)-Y?)98>#TJK==.7I72).;<5IN&+RFM
aLW)9Z;+4HK2&GF2NUQ5OY]B6A70PW5]OVS_3YTG9Ke=:5c2J=A7L)56e+Q:3-A:
3O30L[BJ13#?Q(^/_bdA>De9<eQ(dYa]Q7/1]+cX=Uc3@?K--BW<XWJW_YM6U1EG
A:e]TALD2b23[gPIOEC37_14RRcf6;>F^F.D@@J^03I[IE3XE,1fX:J]B:d=03eL
bC+Y4Y(.e(R+AHA0+f#<JE/I(gIc-LEcK3N6OL@#+Cb5/&fGT(PaJP8?XYMUZW:B
&4RebPJ=H\[NJ4AWE\fc_@bNS[(IA_/]5D.T6.MLT8gZJ1/.OFD.397P2KKL239R
ZRIDbZc//(PDM+9)3Z?-CE?WKP-#@7KCJA_F3<6ebZ^LTXM^6OdDV9B)/^S&0AMZ
VI[45JZVY^539Y[)P(ERRCL@O^X/+AVVC8[HR74,>SC>bT5GEP^DG(7M[7A?C)4@
SU&gMQTfO#Y(cDPbLW^L>98Sd8?OZ;H7XIeL+J=@_FO;7GZ9Yef48>PWb\2;C0;V
@WO?;:J)@Q5KE4CB?]AD3Z>&WBKEDL>OEgR]?@.5L4ZYM&.<gOaSE#6Rec_.f29,
HX7XY8G3\Q50LH6IFY^ddCJ+G:4#=Y/dF):Y<8TKcc_6]#EDTXDRb<_ZO;JCOaV]
1#dfD.:F.WD)@Pb?T@>GO.(3e8cJa[7R/IMUC]8J>?e6#W;+W;<#RKL409Acb5>6
eD_1D/1(eARc&JG7f@7E,_;4L^13(N>CET>KRUbNgXRB5J>-bS^3aKF7>KHcE;DW
4X1+_K\UJ5J+c/5A)gJ>]L>)5e/70b76eWA6Z=MP8WG0aYHA0+&#J<1[gQ6]^\fF
BJ1?fSIYK\a89S7#:E+UUD<5DdGNG^f#0LbGdR0=T:aa<4:Bbae(2NN]H0g-TcB1
9?0]HXN4K6:);+6P#3X\,LQ\fJaF\G1Ha@g-dNJYG9&[G,^>Dc2ZRg9T]?g93ITB
QDE?;5\527QfE?WEDC]5RFJ1>#T?VXQ]4[C#F-#U00=9,50cV0#K1W]TVP2T92\7
b#[=?:\aV_Y7A&KPH67df6a+,YB1V8B=eB/JHgN:@U/2+/K6TgM<GK?YIKc]2W\>
;=;?\R4O@@VL3aY:TICK#>O+JW0g8ERBLRKK3_KYI-.3;fALDJJ?O[[9Z\TP5.EV
g_SH8R[)F3J]_;JV9Z_L-bCZdaJTC=:A-g,R7b?2#WFJ(OZ<-e64@NKcQ,W8G,T&
LE?5@NY]#&AVRC]:e/.?e,Y/[()Ub;HH-N1EQ3^[):A#U6C^Rg3G#c/#7+K-KQU6
NaH>SWXC6KW:g#7HZT3[U5N@)KQc^?b#>0YG_K;MRMLc7K<K#4g+XG&+Q(eQFFL?
]\Z>>4BZLPbGa\.5.Z-+Z90&bUd&.8cHW>3QKEaa,8:Yd^+?9AM&&&TSV0Y[J83;
9[.]VP)-P8.f./O_4_XD<S[WXJAGafB5G_9]b8>XSO2;)O3K>TTW+S#VQ.;[S.#5
NB)F]U]dAd#2=/aL,QW,A747bY(g.()/MP-CB(A,78R11+/cB4b;^416?#YBZe)X
XcaJ8Gce?5S,]JRb][\0?)N4Z+.?YHX3\LNHQA+)3e^3X:A6K)W/R?T77dV0]GgC
VJWRUQ#C?&[9FS1N#/NdC/gSR\X2I/R&CF?X=1(1J5S3AgMcMP\a^_;7egV8X+DF
E9\@X>SI,Q]?N5J;3f9:(B./5ggcA.JVOe=e6.f3VUMC1d4H,\Ba5HEb.cLQDUS5
=0<GdQg=M]<FJCUJKC=Q[fU5aE^<OBNCV9[&OA)R^--JVe^,5@@5UZf4]F5K5+?V
/4b\[c&/WP3T#0?UgE[cYHd^ELR-KbC#3UOWGY9#5/B4K=.,UO8\:f6/Y@JPHM&2
#(66,-:b@K&-Lg(TX<.(7)G+HOHH9()dGXS)TE9T#Z2=EDF>4(J04TCCA@Qc_M3H
3Yc5-RGH9Ja3Gd(JFEGE(KRBM@=fB3Lc[Pd=#T&;X&4Gac\/[SgaKJT.&KKQ2J5F
:ZH:a6\KYa-_H@F>/2OA<I>5SO(=@\:GcIB@7L-RY\AL>//3K\UGE=05?M9VHP3V
TM(2P)DF97IW+/29I5;Hd7/7g>I(Rbb[f#\6>8G?VV=_T@X.\F>fRL6;>#BM1=S?
KSPZ/Cd=f.(F4B6-f:?XK3bCBb(X:S]K9/Sg4=R[eQg=,a9X6#;2T^Ig]fd9C9\b
\Z]T[DD7Ad7/)B^4D]LE3M,9+0O3+:.X[)CSS^(:fT0\ZX6F3_B,MDXg6=7;ebbI
P9FAT+OV9+--09_Q^)7TN<@8UJPB+?(?;J(cDY55(G:Va(SSK_-dQ8(1^gYZ,:SZ
PAX-^/-)Ce[OME7^bEZ/MAW[-@>#81VV]H\]6-,0b&O[&MYI:M#N_<^O?(\Ja),d
#a3ZN6+-dMWCYeG<52U;CPDGQ0NF9#\E-(H(edN7B#YR77.SeSX[@8QN4>S;O@=.
QNA4Kf_QDJHbeE,Y#I,_eCY]6BZ/HcBZZLG,WLCS]7T:PZIL>+I/<33-f-AGXSK@
0H6I/^>/f6_5_Ob-\ZMa_gP#gP[/be.7YE^b3\7TI,9=R49BNW=gP\\Z_XOL6V[B
/QdT+BfK&970YQLbfJU4_C8/#/EC9D:R/I6/a1C9b5JP2Z3eR6Q^Z,H;bc,a;LN4
@5,T&&07D8)X6O]&ZNG1N,0>75/KFR]JcZ)K?P\AM&QNTYX]/N5aW_M?OfG#J2@?
(PEYGJaY9EO1#c+?^X34Mb(E&5[Yf.I7<;S,\<?&=fI(\,8,_QB.f@A5<>&ML7C/
BcP)ZePZ.dQ@Qb?b3C-N6[,CH9fd5?B2S^CCRdO1A:f^5NZMBfC.XPXNA+;V2VgW
Y9LMX;6G=O60&33Bd6-KegKb29Q)UaIDA8fK/B:7(?;fRUC+cRV/D<aRKcSfU^,+
Cad0=#ST4cC1];;Qa/f>K>/XJ1+c&0[27KTNfQ]78<g^[(I1/f@S):/FPcWUEFc[
2Ag_A4\4_P=-X6;eABfUX?)f&f+N9WW]AWCRZ+:H1H(e5AAbQTC/S7>8V0:F<Y(H
;BY-+;OZ3L(@?ZJg)JEd[16V<#b?[[f](5KDcLJ1:C<SZYZPfC[+E#LZYX3?UWT=
TbM3@PV3^^XY/RW+FW@M3NQ+#<=H^JbU&CcL1C-..QaQ)RbIAAXf7#MMKRRb+=C=
P=cPNQf]Z#eL,6)=NKB1WFC+b#1#I4<e^&cVJ_39cW7_:31L(@e/HCgEGNS(D_EH
#^(d_QVcCS+g(cA-++_a,OY)W7T5JWOaDRMMf5,7#1XQJgG.B=]G53GcO0[Pc>SC
S:ZJWHZ.K2Rg/$
`endprotected


/**
  * Defines a system domain map. Refer Section C 1.6.1 on Domains. 
  * Applicable when svt_axi_port_configuration::AXI_ACE is used in
  * any of the ports.
  * Each inner domain/outer domain/non-shareable domain/system shareable domain
  * is represented by an instance of this class. There can be multiple address
  * ranges for a single domain, but no address range should overlap. 
  * For example if M0 and M1 are in the inner domain and share the 
  * addresses (0x00-0xFF and 0x200-0x2FF), the following apply:
  * domain_type     = svt_axi_system_domain_item::INNERSHAREABLE
  * start_addr[0]   = 0x00
  * end_addr[0]     = 0xFF
  * start_addr[1]   = 0x200
  * end_addr[1]     = 0x2FF
  * domain_idx      = <user defined unique integer idx>
  * master_ports[] = {0,1};
  * The following utility methods are provided in svt_axi_system_configuration
  * to define and set the above variables
  * svt_axi_system_configuration::create_new_domain();
  * svt_axi_system_configuration::set_addr_for_domain();
  */

class svt_axi_system_domain_item extends `SVT_DATA_TYPE; 

  /**
   * Enum to represent levels of shareability domains.
   */
  typedef enum bit [1:0] {
    NONSHAREABLE      = `SVT_AXI_DOMAIN_TYPE_NONSHAREABLE,
    INNERSHAREABLE    = `SVT_AXI_DOMAIN_TYPE_INNERSHAREABLE,
    OUTERSHAREABLE    = `SVT_AXI_DOMAIN_TYPE_OUTERSHAREABLE,
    SYSTEMSHAREABLE   = `SVT_AXI_DOMAIN_TYPE_SYSTEMSHAREABLE
  } system_domain_type_enum;

  /**
    * The domain type corresponding to this instance
    */
  system_domain_type_enum            domain_type;

  /** 
    * A unique integer id for this domain. If there are multiple  entries
    * (eg: multiple start_addr, end_addr entries) for the same domain,
    * this variable identifies which domain these entries refer to.
    */
  int                                domain_idx;

  /** Starting addresses of shareability address range. */
  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0]   start_addr[];

  /** Ending addresses of shareability address range */
  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0]   end_addr[];

  /**
    * The masters belonging to this domain.
    * <b>min val:</b> 0 
    * <b>max val:</b> \`SVT_AXI_MAX_NUM_MASTERS-1
    */
  int                                master_ports[];

 
  `ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
   extern function new (string name = "svt_axi_system_domain_item");
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
  extern function new (string name = "svt_axi_system_domain_item");
`else
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param log Instance name of the log. 
    */
`svt_vmm_data_new(svt_axi_system_domain_item)
  extern function new (vmm_log log = null);
`endif

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object used for logging.
   */
  extern function string get_mcd_class_name ();


`ifdef SVT_UVM_TECHNOLOGY
`elsif SVT_OVM_TECHNOLOGY
`else
  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);

  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );

  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);

  //----------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of
    * this class.
    */

  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */

// ---------------------------------------------------------------------------
  extern virtual function svt_pattern do_allocate_pattern();
  /** @cond PRIVATE */
  extern function bit get_address_shareability(int port_id, 
                                        bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,
                                        output system_domain_type_enum addr_domain_type,
                                        output bit error
                                       );
  /** @endcond */


  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************

  `svt_data_member_begin(svt_axi_system_domain_item)
      `svt_data_member_end(svt_axi_system_domain_item)

endclass

// -----------------------------------------------------------------------------
/** 
System Configuration Class Utility methods definition.
*/

`protected
ZP/3g>O<5.ge:,\JA=X0,@;:8/FN<.N?/.+T&?Q;:=(P5P&&\KUS4)=.&eS].,+/
/XF#9LW[YF,\YDb_PaUF87Pb0[TSTPfI::?87f8FD;<H)ZHdP,(+86QAHM+8GC32
ANA[DTSB>c(G]IHD#2?C;Fg1]G=FT[_P(CBGPP-HafK<@2D&2X;WXY+^Z@^8)&P6
^@YH6&M.3+RXI.Meb7:Y,ZFaIX3^=6b.b^T^OWg&Tg-?2SNT0#+Ba:aXTD9g.E\\
:U&+7GF^5;7ER)LR=g8fTB<+P?;QJR\<f&eK++\(XeT)P5_GF8&6d.J1DfE99;Y&
HeXf8J>>-IK9)bCS[fU)Je:e2_^H+N5UE/_?2VNJOB<gCe>DA=&OX4Q^-F4K\920
Z.+132L-]U9f+GP[JNacO+UW/bW6FI)\;aTQaJEAP2LFaI8NU.SKd(a1[L4\Pce1
[Z,;S7aOM:_cPM=X6g__HI[Z2dILg^;CAHFN.^g/V:5_:>egL#EK4=/\dIb-KS(f
XD6:P+793#WE:7?_4^VLKH8;B_-g7Y.R:AZbI6.HR_]6+NQLGd3M/3^+VDWHA@5d
f#YKS/1#Y@=Mf_TaNDC6/ELD]9c65cEb9d<RCFO4]c#TfASdW)#)8/K=_+W)J45A
K-=b[L>2=<O2N(CSZR6)ee@Q1>D=XK?YXa;^Z)9cF2+GN)E07K2R8VK=N$
`endprotected


//vcs_vip_protect
`protected
V#fN5))9MNd4UeR\_8(9DDAMLD^_8V95f[4^UP8aSW>-_HC,9RD:2(T7/Ed7<U@P
cO=WPO6J_>&2LcVR:ZcU-F<Pf_X#eaUEG\a@-(=)V0KAR)SA61VT062,Pceb2B0D
?Z4IJ)>L#D&V+ReQ51FfZ]0<T]d+eVCTG=S9.cEW=_aDP\D9<Za,>]R4M@UAe&^1
HeGT(D:QG0N&3U<V+:0.><BGbc88:T<R^L,H4f;Y[?FVDVL1cOML^BOGc.Pg(0X>
^Uab=K-TS@A20Q9T&=_;R<a3VTW6#X9(EV^\_/[HIKda2?-b>V)WJL?O.MX4]OIH
9MK^2(MdP5B-QZE0]dVd0CQg>EZf:&QB4CL3.\UXcCA90aGBI>Q2E11;0AI]1_Y#
\D3g^7G8Z8Q[<_ObA<]1gC+]8gX9KN6^<X>-YWOHUJHa_,fQP.(JS>:IA=R+2>HI
-K6K^eZd5[10JeRN<ISE7_<GD_gL=3DD#gSZM@&b(MUc/7RU80(BPC)b:T,YbAeN
N=HVD2<JXWO3\RRE1^?WQ3XA>M]]?@B?OBAI_O;c;g]7=gXV-6)8QV5[L<V71DF?
/:JRS1:bd7,6c-F&Z46UTRD6K\MY.Q##J]K1WD7IV,<b+EQKN.^R&EcT,#C/+3[f
D:#7Q\dYQFd5+R.Z>JHR:(aGU&7:b^6/+6/J#1NdV5T5F+C+LHbQ4XT+T\-gI:;S
IZ/+^fCK_[c,OL[>cJC1VC041eRgUI[aDgGA3,Na_WNAZ:eZ;[&ELXMB=a7LFIRd
T@A,>M/;S:WT@I>)CNOG)L-4:GBN>b)J6+44#cFCXNO&]c?U5[G#P(#GQMS57g3R
IN<P\dAB#Y^>37d0U3<N.<D;]c]EC<LXXb:,X\[R;UcL=VD6S;@@BWOS7E?aY=1g
bREfKD[>cZKRL1fWLN^?(/_-HP3e45)<B^G8I-T78ROe[2IR&#_1/UI)A:Q7Y:&-
BP;V+QV#ac/5G;I;D3=,EMS8;GC4;cbB9NLR9_1[#Q)H-;\@_ZT&G671JGUP<BB)
76Z00D-&6>9/gO/9A^@W^WVbIc/C[(84(F9@d<a#140^-0<<UW1Q7aSNf?B,Fb1L
ccM_>Qd8FYT53C)ELg9V^3fBS\21[9ER/7Zc[.Pb1A,;W;e@D5WPYa.?.X6JHAP@
Z9<-bFHBWQ@8CJ86^>G<TUPKI19WRH\GgGOTbOg)TgCM<RRb@(:DI5[F8[O-THb3
7DR0N]Z<^_,G;AC5CgK0UHIVWfK:YQg7#2Q5?QGWT5TW\0M&EdY1N2A3\GOLEJLU
&-P1\VC&E<AT2.+fMO7a21QU0<&A;YH;XSdJHgVQgA_gRN&0TK>&0<dS8\:,GcO5
>b=4A,>X8>3a4II@6R9+P\MO(N28SfTLIdM5QZ9V[_+WC4<AD&JT+UT9VPI\8CC)
S.>::YC4JKO-@D7&I^J_4I+]++)1>#AE._Q>f4:96<P,1]CO-c.:-ZKH1\[2./FU
4U1Q1cH<8SJ<.4(@IH<2#<NAN5VGXRPLD,^VfBbgF<cD?O6QKYfUfWW((Ve<(>E-
120D<;)D8cbf]4AY<BIC\IfJ#0)K&[F:WBM_@:2dH9B_^TA6O=[9-)@/g2229+#d
1JX3>41X)QWT>JBa@X<QCU85N,/IT4-PCM;3KG@]d7137F;,OU?b;&/L+fD-YCYb
L)D(O5IJaWaK/=-0_J9+O>5]U06:=A-8O,_,9Jg8/?_Z\VDIJUFA7ZWJB^]MTX->
?)AY]gO-a=^<MROfPQf8RS0:N+:g93<BG:Bf[?b=H6PF)c\NGFcU(cR>aSQB_7#A
cM+g6V;XQNacab#5R6Y&=dB=2/3PVUK/R?B=?B<M2X5eG-.g1E5]5TCIS\O@EV09
fYg61A^@5?caOW+QD<44K)[+)60K?AX\^?X>>;X5QN^[YFID)E1J^;\T&3/>EbKQ
7R:&&e#a6\.F/:-,M@45,@Y0IO\9Y-/(HFER-NC08]Z4#/B\#[Ue&cCgF&W)QA^+
<4C\c6dQg7fT-#8.UZf:8,V.1+^P6L6&CO[[W.,aUU+J<F,IgX-b#H/[gEI_bV;]
79WINaGSP/XN89=I1)dEO]<a64&[d3b;bL.R&P(,)+4KV(@,TYQ.QU?M]Me\^(/-
F#P5<H<-GIH7):94a5bc3\AGb)E_&0D89dVWcd92R;4:5<^+a7F_-HaODY]N)WMM
+_c5(F/0IFbMENL=\FH7@+K7VLU3GFEfJ.^XKIPFQ/O20CL6VCMb;OSb.+TWZ&CC
D0;9EU,O[gfC<<=H(\2)[F@<J+K&&_#9,caCf5P9;UH5&3;&.VdgW1BJ,0gTD_Z5
F6MLg-W3?IC=W/YU><E;dLKI?L_@8Yb)fJ36ZFOA#5?)9/2K:G?,I?#0?9P)]4J,
;fPRIX5BcL^+/O>.W(DJ.EQEDHK\GEWa7e@Z4@OOc-03BO)I?dBLFV>I^RS/0M+\
YW77X;M)>BQ?]#gP3T.TTea4>@[03]KSPaGQ6KE[[0&M)bN]VZ[7=3,)\d)DaHg9
BMW+,c17NEGKb+Md8PUY5Z_SN35WSJ-L.[fZ,<^]0J[,E8&8T0.dfBb/?TJ\CFN\
.WQ8T)8_1M\/+T#4-c[]K(EH<_B_QgPe^MI6NGLSEMX-SB66<7dZGOVee/]^gT)[
64[La-efKU#>db2JM+gSMZ8HOeE#0RCV]MMV2I:X,1Q4@R.)7_)e9GLTA#&@Z?gD
/AfCCY[5Gfb>@R(4XcgSW7Y+6OaZE\C&HGA-44D:K/dRGNDUKJENca\:9GH+5L=&
?)5eG3#8Y/f)DK^P/#E5L8eVJR#c,0gYE2b<dC4\6]#&1-BV#;Y18HXGQ,T+d\XN
C8<P<cP=.OQeYd@.dG),G]fE.aYQ^9>=7d7OO+RXP5Ha)G.>87&2AZ-HJR(K;<HH
SDZ\Q?1Z5)O-_A06XHY+&RXRIXNP83Q3;g/8ONJU8Y>SLZ[,f1FJY^86UT_.Q\c/
=_bbPaf-,[/GGFAYQP>]O.RTC[Y19VfGO9BW]IbUY>_1_]#1fTS2-9G(^\>Z@[NQ
.F7\eIK>[O;,1]?=WV:eU+MNJ,e26)))bHF>3V_L426Jc/B[)GGHO2&M&Pf&c>#,
=+JHWF3^&Z.WJ(=U,,2<:@&I(4R_#H#NE[=e_N]V,N;JCEVRc/\LHT09WBOCbP6A
ZXJaN>)W2E04XB5fZE_<_=WaAY0@g[:3=bWYC+e3]e8>aM=gg:ZDK@@278.LCXPI
cX_U\HX7FX3Y,c#URU(,M&)C(\Z/R]NKV]<F_E_#b.5&#dOB>JRU-YX2a\>?/9H=
YWe>&6GCcC-]M6;CK\=aM(C6DOZVIIF/X<eY=@]cf/Q1Z.AVMZKV&@8==RP7(8\X
?b>S9DXZ,YTBa]TB0968fK4ZK7dZ.OCKA\+gTEWYM32-I=D=-0BfB2EY]Q.c=KQ#
LZbP#\Sc/V:0M+H@#&f0\D?D9Sd1C:N.Y.4FU;J1)4O020GU__G@/YFSE11]):7R
0cd6b)6;2=GY>_A]QcUC2?+P3R@=,DDB-()[gS_#2[R0b]I5X]G:1L3JJV8XD_]b
MR[TY8?F1b=HY4Xg59CV?481LC_a9Eb(_>>&MbW6(-Z?,91FZL]R9E##@^UMO258
T;E85gd>;a^MNF./OZBD];]K&5g]96_?=-/7Z,O+(+CBMe+P<2K#MIM4g8VXA(_S
P=5/E->RTbFWR?2V/_F44I23XRF0b/RfS@YJ:G/X4?c\;&S>Q]V@-B?-E1>8V[Y0
727FVd+JbV_:/5>_3J[PdS>:\b.XH,&a&_D4gcUHfeV]+cGI\466A^92eAJCH@:Y
-@EV8(4T)Qa?OA2I)0Z3V]deLEgI-PZ/92HgAXF?\0VTIL9ZQMHD00:VYC-)><3.
G9YBMaC[c\[[g<S87eS[8Ha+Hf6JCNPS1]+Bb?J8a=2T?dQBQB\?TU6&(3C0[V?O
Ga9VVYe7W^^H26&5F139g2-BXaPC]5gFbRR3?61fegLFFC[IO>JBeFCZ]X\Vf134
U=ZbO]]c<4USE]5d;.cK]Zc<WE7J2gAIe[3T7-cC4TXa@6Y6_/LK8W+V&4##U?/8
UdWd@0VF[3U)\eKeL+U,9?1FQ1NO/Q>8+e&JI\;S(5SD4HeE<?]/2L[<@K]6Z-gf
]I1d#PP0d]4CSMC2C&C=?IC:](eF?E/VC/a7^eL/_WDN.Ug0gLKf?_K7Q#TV&6W_
1_Z<-Y=^?FG_4+KC5K)DC>PO8-N,)K-+;<A-HXLLBUc8M9;DQMc;6.)ZTZ-F?)\:
(5L]G.abO4PH=dDK,b+0J;@C.M.B\8L?6;IUb_T899bQUZ[[\IJW[VLcPT:\gNQM
F8_aLIL,Z:;&\EZ3ccD?)_2ae=OG.NS<IO,AN2aAV9&7+8>C,3.O40da_4BCff&N
c-[Abf<V3PAa5;T5D[2[0E4ZfgFFUBa@;\.SJ:[CWa3bUP=]Ve-XP@be1#PeIbT+
.R&e=P^&-[D8^OMZVEE8[[dLL&TS2QSXCg\WG=6#XagHBe/8b#B(_BZ7bA;4OB+<
F+>Mf3:+gN7c+52QBWL+7?LU39M80SDE/e,#4-L]JH3bWCQRe?3H;aVdXYUQFB(1
d<XTKdQa713LbgE9b0@\+,99WQ/2/f3S25Redb6D58Z@#J+8W\5cF)T?6M^0LZ=b
Xgc^I#UO/Z/WNV)-Y&04/HJCDVU7N-3?LF+a?A6NX8>W_UV2<Qca42EN?3/3A#=2
XIeF?^-J@]RWV.I=e>B-30;\U5a5CM0=U591:J,O^/8XO@+F[caWXESe?PM+de0I
b>(e(W93EBeHR=,RO)>6c^72UVD;=T/4;5Q:9GG6M00b[I;NLU]^3aY7ZC^#<&eZ
BG5A6ae.aR)E?c,RaXU97F67^U]+J:RbU<C1TO3+K@CWFb4:F#?+SNHcKaXUP4XG
NdTB6Dd2=QAf&SgTb)R.O(feDW4VX8Y&H\fLPIBC[VJB/ZJ>e:V=38R#.[3f)VU8
PV)F8VSd;]_G&L1Fgd&O:A_e;QTf]:_TDe0<J;JQE]43/H-F=MQ(7W:HCL>UWVRP
gbPFVPX15e9a=IM+:MJR3>a[OSe>7S,WLd.g0TW?#K/&)/4ARSZC>LL;H)4DJ^ZW
)U>/b(.E<(AYa2eZ:4HcbP)DeQ\8cJE.K:3F-9FO([_+]?T7:21dUHR2,Y][=K]f
D?N3=PRV0M[>9L/QcfV8H4):&EIP\&O]T[-4Z>N[URcP.I^HV14=/Qb2F@/^FTV=
6<8Q8/d0+d&.1I:URg+J;)^P@1_Z1a-Aeff/43-._]d1O[Q)^:R]dX^4]@<H<b8)
FN?4OFM]0_5.UP;URJd.UWTM:+53BY.BLFD.46:UV2KNS9fGP-Qd@_,+2,.]bUc[
I=7UH;Z^2_KT7S+FUX.5C0&.6&g-6.b/:>]H><+?Q)g#JA2W;e_T)CQO)7ca1W&X
QNH^PRP)5C0W6g=?]9P[e8,#AK\a;\bUN0:3H1\JRT,B,<N4E8ga[;f2\/@,0=e+
df6ae-U43Z)+f:0CZ6>(_HL7]CDPDd[LKXV:.QWR\=CM&U?NVDH4TgV1KQP&a\16
[_L7H/a9U)a7<0F1=1)]#:1@]>\I\f?A\6B39DP1(YT7=f@5:T@-)@.E?,+aPV@9
##OX4-W.D-7<FIc5CAgeT05]0DWS?8VT#?G(49IBIEbZ&P81V_T\-1N[1UA51G2H
R#(/41Db]I<AY@45MX/E)V[D//8959,(0-Md0:<--0#cV8)QIc/ad>AfQfC@M.2T
b9@eO(RXZ2QT5SBHBd^RA>3L&M]E>Q#)+5Y>0ZXYDf?QJBZ&/#:H[(D?)g,UFGM+
1H)KecdDNMXLaTBeQA/eQE3VRg+2^8.:#TUcQ3QXQ]bC:^E/K<FP2;UdVM(_A9-F
,&3O:)Q4dB+(SP:S<NQ8>cU6eYM@S[NGbKKATd6H1N762:3F7f3\P3[DBODR&J.2
\K\NBF.eC\bG_2\.bNd][T5&[BHL:86@+>6fI/Z8OVbP/<25)JYFQb#0X5X-(9U\
H[:U+2HM=\F+&G>SQ+)2+^S2_)OL1V4)PSN.AJ#-dA:6c?RedQgY0=cY8fS>,V4^
]deBbB6NT]CEQ=<PXec_4>HacCWV9^BD/&VA#Lg/VcEP:0)>V99?QR^1e^]B05gN
)XKR=gK4[Zd8b._/^(E()/Y1c<#fQ#b&)d@2UYfb2,2ONfHd-0V;I_A-ZeG3+g;?
a<^2g/;>0LQ3K&C&#/]DfdZD+8&(+#4H:?R.WLa2(?GJU10U^4LW?3#9X(/3&PG:
FQaP75:Ja;d3Q/AgR\,O-(M18fW+]U^.+>(.GI+U+3_bIA7f#8P?e/<UD&c8POa2
.a:>WU4PVCM^XKc<ZPWUc[c7W_GRP:Q.)->LTY<^#B)@GD?Y12?HdOT+HSbgJDJE
>])@AO#X7:-1O7cB/UX3H]fYRefQY\K,-Y1R_0FN0&5TJ>ggQ4JCbR&-^X7&V<R]
:)c(-_1c<GT?b=3bbcC;QYdJI;?^#W:^eX072?Ig@-^NDc+FGga2I]gGE>GQL^,#
UZLNfR?/@X,DO1Fg:\cO(3LLaH]E0)f7aM,AC5J?1bJe1]DI/)@HANI/&4JJ>_D]
]W#1YaeK#)D>bQ#\,)HWa3\4Y08>6MZCQF)\d-G96g+dFea5[3)&Z1bYNM3I3?B7
H7?b05?7(^#\1SP2T<G(?Jf4JN;S)?]OQP&B#N/U9#]JK-W#3_8.JNBOIIJJ(@R^
S,=^]/_YX7[4Kb,ccM)WY7D1?H1J]a&+?MXfPF0M1c2#2Z#]UO8#:;@JBcJU8^/W
-+YQ;]8J-K9(Od0)R.eISMgK]IT>MgV8],I-/S&]^]:a)@f0_C&5#KD;[;N,VJ9I
9^YfRD6O9ZPI71I<P1^??Z6U((W?I;B[J(fG1+29KMbV]RR7R7&C1XZ=fGVg:X)#
8-^M-R/0EUD<_c8M8Y(bQ-B<84X+3^b^E7be7Z]<9HcG-W9K@d/@beV7M8())A;=
H>X?T[9JH[IgIaONgQ2]bRSC9\6f#=?G-S3Tea.fI+ZMP<OTRI.[38aIA)=gf=W^
GI]<RP</C<T5(U-\#KfLH:Z.abP1[K=Sg8Q=L+1G#[#(8\G@IDd+5AWT?D06aC.c
bN&&KOF:MgV]/ENb]?>BC2[)=?\U\QH<AT_W+\=@FUdCg(S.&^Z3P[3AW6YEP()P
eVUE@faAUXPdK?44@/Q@HCaQFT>c)L2ZGYV).7(LE-61^Xe))R/\&5/7TfY\Q<>/
e/#-,1O?1VB-GQa)U5-S:f:MK.aX#7D5PGM>0?32=98_=BdKXSD0M:P1d26.3W])
-gM1_-.)c?)gQ)2e/?2Z5:<PSJaX_9P/P8\H/-+RM5/#ZDWZ8WM&V;+Z#X_GCU6]
SK@^=:X;Y2][H(@?^.QTY8(6\LE70UY:TgDUdMeTSeDc(K)4J:+2MfE7cH\<d;Ra
58X,H61gKR-MEPMU[BI)0))2XV#1C.>b^R=ORW.b2+.f[,#S9N/BS_VW,8e7eMgZ
c1eP#([9e<3fE]O?^12g_PCO2D-3:51/RFSEC[97TN(,GcBP]1OI-f+Y93RL(]\X
J5D&4[]XK[B#9C7JT,edK)M4+#+dSJ<dCZ#Lc-7EU]Qe-<a(F/34\aW6G3A<@dcM
6Y_^4W<T<,Ka&>[X58LPF3^=,c6C:^(E&&P/PF(bEFS>f?+CYbT@E)Be7CJ6)4_f
B08]f^>C_&>-J.O8YfQ[K-BZ0HN9a8=QDP\OGY4:8\&9@\P\6#RN]fgX3VaYD#P8
cN.M_V14U9Z7R0=S/8(VLGY+NSSeSVY;+-E4Se::a2/G@ZSW(+J>><.ObUW;Fe#f
#ZW9O0<1R]K+:W@YF+eK50=@\(>-+5B3M4N)Le8/58^NfYF3WNddU50,A\=TO>cf
\:f/K)TEfM_WFc;H]R)6N#VZM+F^f+K45eAJ)0fB[W=>?a1<Qd/#f1=[_8Rc_dcZ
&K6O6\ffP3Vf]53cfFF;aAV[G:Y+?U->[[6CRgLDS2PbW3D_BE_HHBD=BE=?(:?O
S(+88W?R.?AB8PHVEGB<V@J3,O[+M3G5T@<XA7;b@KJ_94KR]Lc)O[JZD-Lb0cJg
EL3Je;(C2+HFfHAIV9fV=;AS<V1=G7c9f_5N-&,2)ZV0aH5Y8@=+]Aaa3]CE7+e8
_g3O,E(Jde977X176X_P@e.FO6E<NdJg?V5d-Z/WM,6-JS-dC)Ya4<bEM9&SC&HD
=)TFR.STQ-Q)L.)5PfCdKU>:@b/>ZSYR0IWX@F0_50FW4>f<GYI>0..5I,,V-CWV
Yd.Ua/Z((?8aaNH9FM\_A&KS_+&XIO)d)EX#g-JAN[Y(7LXgbcJ+_NWQaG1AS#;T
_QMDIRKS\9E-X7CB@VB1ROP?b-CXCdXM;NgS9XI>a8J77RgLUL@V91W5;+P@SCfC
[95AMR1Q=:M&3Z@Q>2H\_BHSI2c/Z12C5=M7M6KH?gCV)SfAf>9/7:?U9a1+SRdc
O>XG>Y2FI>KeJB[##IO1O5V;?cD7Zd5V37U#]f,C_K]2FVf(e@MP1<Of6G+g7I:3
<UZ.B[39f&KF]S0I,ZKQIR1cf;A5FYR>QHJLYeUFLQ>P\Z2X([)+=bUfUSX,YbaI
\?C9N)(71658.UZcD?DX&K_7#KGCHO(3XE82236/=X;K^=J&.f9O:0\)7PG;X(P\
V7CID:LA_#?W3OT=OgP&+HFPOBF1&1S=2[c-OUcN]TN#2gN?HE-F;D?.ZV+6\gfD
Eb@HL>A0cZ/e_9JC(4@fI?]Z[7aZ@\4CHYC1@B2KgeD2=.H29Fd<4G(L6MW^;K,6
(X@UF9P@]3,gC7^+(e3X)ZI-JOU-=5T.5f+W9@GRD;ZL:T_SI(V)[&3,b=H8PVeb
ffeF9OF,L5e3)UDG+ReZL1SX5,RW]=(@H+#d[,IXFFQ0?c\:5d@(JeV+0))@U/BQ
:O5U\1Y4R#g-KgB<Y#5P//S?U>3G6B(@SeXc@-](Vb>D1QMMe^7Y^7O9]6Fa8I1O
BI+=0cJV3(abfWdF\<@T^Wg87IWeG?T.#2GBa.FY0;2<PJW8.eR2>W[58fQbJW^^
cJ-c#E4GA(_Z<gS:+AdeSS514ffV=08(]a]A_c/CC6c@0Z/a@gFNML\V(;SNc-MQ
OMeEI5)_LK+db7b6/:E#A_3b0<C1ea,.H000c0&N&PUUe.F.a7<4.eMbAP]Pb/cV
+gPNV53Z+U4XR3C9X[03CQTfK-eSb/@4NB12<7g[Cge746B<SVF.:feg0EUgeaD0
>[R@3NcT^4dDZB:^]Uf(W-C[S^b@H#63(g=U/&[C])gX463+E0@&=.0a0AG[H=MS
VHDN,#0[_J=]+a@[49?g=O#3E+)bXZ76EKFY&Pd?^+BEQE_Q,49O^<aRF6FcX0RF
IWC+/-=P3FD,e5(MQR&?<1+)DERG/)1:I;8&(+N?EK8>N1>^ae41K34I,OUSe5[d
@WO61QS6H3Z9E\WZ^eN(V?[?)4YP<<?U]JIa^EN.,9&^,3Sc7=2[_DKQ_9<MIgTR
59JK)VK(Wb;XJ2;EIF5IX)>HeB\ZPRb<IYSH)f)BI?VZ>TaPCI\),O^UbcV426C?
dD6/HL+>,0@d4.:g+\UT+35+RJVJ(SRBKRIT<R:Vb6>,aBgJUU04Ra77MR0X\^2-
1(bESPXe=G<F#=&R1FJ@dM/&(H15gaN<?JMf=-_RVd&UCZ-\D.S6S;A/Y?8@7)7K
NUXO,I8BG?O\5,US+XYU6;a-ZCeB[<b=WNMREF@2QYPO>3SEDWB\fPU8YCB[Q/>J
#K/0+HAA&H<-Md+GDVKRLT7G>c5^KJ:-S:X]_]3#?40]=DI\#23D,9+XZ[?OUc:/
7.(/3fF669=e/R<\GA\)(F;:WBLF?G3H<S8,G.8-8@b;dFd&D_N9.7-Y5\A)SS.?
<UdbSc^C2RW)Bb:e,4c-Q;P?ZUD/25eQ<SS>Y:EV\IaP_RCRPI0+b/X_eDU:>0Mf
G[.#(22L8(ZHU2R>?2Bb@A6;2=?UPZ?.5ZO)e:(H+f+26&a(Rb_PL51B3B1a;[3Z
T[UA\T&4[@,]F1S0;<B<\11OOJRV-GR#S=G9P>N+<G\S]R)g79<SCFg2GE([gd52
GbfB5DVVIg?cH;<78T5D,XYXK;<UQ_PQ.7\2ZS[-;F)[[I/G^6c<Q4f]VATG(M,;
a2<54GH>4ZF]c,S=C_]?4=A_&K\4gfXWa[W<MaM/?\VJ&27#<=BO28gLC+R1IGcG
KJN@L_c#.7dZY55X.U,DZST1/L1..CT0e+&G?&,7<Y[HgV9#?D_T/:4-_M4/-0&U
C75L4ecXA6c3ANa;=3+XO0HT6].64LEQ=K)-(GOOR-TAdg>[@g-_W_-<@->c\?Wf
C>;O5Ce@FR,cK>GWCd5@R\XbR&.Ug1c@2_dWc9C@4RVcWF^eCcD8K3XHMK,bUf2G
<TDfS)g<VaZNXRG5;+89F7FLf<-3;(/R+O-:J>QJEVT\BNJ73Ncf],3c=H7)Z1ZM
O3T8FX=abA(?KJWU2@Sc_C=6bVg4<^C#D:Od,FZJS:[E5-(AS;UY[Md38[S#AL-@
/RgZ)Bf#_K[MI<Z1&L:Wc_fY[0#XbN=NQXJbDN]#;C&U84(e)aSd7ddW<H<ede4H
3K\b/^6PObg0gbGYGY2YS^[^YBL\+ZOOIP?G7A/fB(ed\?^dUL1J[E9AQa3Va&[.
^-E((<cG?W&PO=B_.\0N96<5RfA^6[_FTEce10XM599W7a1e44@.S&5]gT_:e);5
=SL7Y5T)UcIGS;UEcc9fR,XZ]3XTR/0d,e9Aae(Z22eUPRWS7X9V5]XJDHPA.QM,
)QX&5D+#KL2AJW7(J^7,<^K9TX#GafH(5d9[,Uc2IWb,\1Ag>S:#UPU=McNP)NEU
YYd#_7Ca-/;]_CHOF5F+OAa6)>7<SIM7L?@[,f;L<86T#[dFUJ[MJASQT)eV[W39
(1e=Y),_7.d^[++2f;1;D,?N@/]83d=POY1HRacEG.5e@OV5)fU2U4FA,[bU39a4
RGHLNXI06FgBN<-aEKI=R&E;/H\-Kg,U.YJ>28;bT(15AD&N@a=O1:7O31F+@L5S
/BJ>fF4]O&Z;E\^GOU617,Y:&X<\E/;/T-=DJB/S-D:5\CHMT0LGV?#WA;JQYLfU
XR@8H&-8GU<B#gN@S->P+OfB<74EJb)fccM&KB\,c(\aQQHIPQ?5<E6:]HDPcEPY
H_AF,KX.A33OPBPW=e+UG0X04.N(LM[fCX#I[Zg+&J9GRI6=C0g3<df<8KPB8T^(
K;D[8U_P>CF:a<<\[8#daE<W8.N3N?<</8?/YGb;YGU:71>bBETJP0&b<a\AfMK&
V/d:4^L3NO,8X.#41NEU?0R:4]L)9^;@N.-T(cZE9fZT0RV4RY3C1]&6<=BWbfP\
H(O>NY>MV\G>^2CBY=>/GJVO;]G2:YEd8NDCLKbBEPWC([5_R0J+VC_=VOH<6b&&
E=0KcL[H@+,B=V5dfDU5SPOb[O5#?c[M.#gJHX,LdCHKN>b]ZL5FSXM.2d47TR\E
<^9^COX)S\d.E8H@OTUZ=eRa?WU>KSd@WPddBG?W<-5GSdU[_JL3]8V(Y;W5S&N9
3Ag6E;S?@M=DK=Eg@VF)-If2(()H9K7N=]g]0FBHfg)(;/,7?Xg]a]b^I)UZHf=I
K2>9Q^QXVJDG#SC-8XUW\0?)ELLY98CX5_DW^fH8)4)6Lg1<G+MQ\a.c.E(?Z1:\
5C/VW]IbdH<AJH5UXaeQZ-Z\OT(ASLVZ]g<+PC9MUd&FAJ@8F4;=8\S#]LGae8,7
VdMM_C-6?cPCN_g70<F+XYQ=d5L3)TRL+AC>(JZ<E);NTXYL/L;^[f<X5b?>C&F_
?+-KK#C=R0I1]S11aXdR:[=M?[PW/M9XE06WARgg96fET)c<7/W,?(aXO^N)_I75
56I;IT3.<bO;Ib&.e:/&PFegIYU(-1AI<QUTB.QB/=UE?U2KVUe_.gP]7;IJ-7/)
</APJC<gaLYF>dDW6+/[OR&_Z94G3Yb0Y&e9eM,:)EDY52UBALG^K-N-,#Tg.<>J
525a)NG2(45LPR<T(?VM@AOK,6:(312F2dE#?1X69Xd2\1#+5AZ#0D86FW7,HFeM
bHU3gD1>OE##-C,aE_LbI[e;@1AUGGaGJSYDU8F5RI;CKScc49MHPWPWJWOd5B1@
RYDb)<RSa&9WR2V0[>W>&?NeDYd,7ef5]bDac9Dg+0[?\K/-SG,W60V/)W9?)5#&
_U-99&MG+UUJLPILA3_?/T@bXB(G98;-Oc.43:[3I_BLSgD3]=,=-IO<50NG[YYA
C?;5LVL&#-6)4Vbc,D0/C1_))SX=be^UO1VD4=[a>GQ?S7Db4?SId5PfO^&=d/>W
B;G/b8@Q-dI3&=U>=<=eddPCc]1_+^f\\MC2Xd29RW;BH(5G\VJ_,DaP3A_R2A_?
5]>2Qe10TWN,BCPBf1/:S8SW:<PJ7Kg+,;Z2ZaK4RC;DYb5A)G-;gX@c.Kec<_D.
/B;ac[:<f#[\(U)F9C1d1^^X>7#Z(B&Q?IPYd<;a_c/>U]BM3,_OOI#<_AY8,DEd
9=4ZA[DM)IM>#fMK85Q78VA85I\/][Q3&9_&UL_0eZ2gYP<6;IV\a(eA@3=45I-V
cI-0@E0_3:)93gB-7TOe8]A82$
`endprotected


/**
    System configuration class contains configuration information which is
    applicable across the entire AXI system. User can specify the system level
    configuration parameters through this class. User needs to provide the
    system configuration to the system subenv from the environment or the
    testcase. The system configuration mainly specifies: 
    - number of master & slave components in the system component
    - port configurations for master and slave components
    - virtual top level AXI interface 
    - address map 
    - timeout values
    .
 
  */
class svt_axi_system_configuration extends svt_configuration;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  /** Custom type definition for virtual AXI interface */
`ifndef __SVDOC__
  typedef virtual svt_axi_if AXI_IF;
`endif // __SVDOC__


  // ****************************************************************************
  // Public Data
  // ****************************************************************************

`ifndef __SVDOC__
  /** Modport providing the system view of the bus */
  AXI_IF axi_if;
`endif

  /**
    @grouphdr axi_generic_sys_config Generic configuration parameters
    This group contains generic attributes
    */

  /**
    @grouphdr axi_clock Clock
    This group contains attributes related to clock
    */

  /**
    @grouphdr axi_master_slave_config Master and slave port configuration
    This group contains attributes which are used to configure master and slave ports within the system
    */

  /**
    @grouphdr interconnect_config Interconnect model configuration
    This group contains attributes which are used to configure Interconnect model
    */

  /**
    @grouphdr axi_addr_map Address map
    This group contains attributes and methods which are used to configure address map
    */

  /**
    @grouphdr axi3_4_timeout Timeout values for AXI3 and AXI4
    This group contains attributes which are used to configure timeout values for AXI3 and AXI4 signals and transactions
    */

  /**
    @grouphdr ace_timeout Timeout values for ACE
    This group contains attributes which are used to configure timeout values for ACE signals. Please also refer to group @groupref axi3_4_timeout for AXI3 and AXI4 timeout attributes.
    */

  /**
    @grouphdr axi4_stream_timeout Timeout values for AXI4 Stream
    This group contains attributes which are used to configure timeout values for AXI3 and AXI4 signals and transactions
    */

  /**
    @grouphdr axi_system_coverage_protocol_checks Coverage and protocol checks related configuration parameters
    This group contains attributes which are used to enable and disable AXI system level coverage and protocol checks
    */

  /**
    @grouphdr ace_system_coverage_protocol_checks Coverage and protocol checks related configuration parameters
    This group contains attributes which are used to enable and disable ACE system level coverage and protocol checks
    */

  /**
    @grouphdr axi_master_slave_xact_correlation Configuration parameters required for correlating master and slave transactions
    This group contains attributes which are used to correlate master transactions to slave transactions based on AxID 
    */

  /**
   * Enum to represent where a chunk of data is specified in a signal.
   */
  typedef enum bit {
    AXI_LSB = `SVT_AXI_LSB,
    AXI_MSB = `SVT_AXI_MSB
  } source_master_info_position_enum;

  /**
   * Enum to represent the coverage of system_axi_master_to_slave_access.
   */
  typedef enum {
    EXHAUSTIVE = 0,
    RANGE_ACCESS = 1
  } system_axi_master_to_slave_access_enum;
  
  /** Enum to represent the L3 cache operation mode */
  typedef enum bit {
    ONLY_EXCLUSIVE_FULL_CACHELINE_IN_L3_CACHE = 0
  } l3_cache_mode_enum;

  /**
   * Enum to represent the version of DVM message.
   */
  typedef enum {
    DVMV8 = 0,
    DVMV8_1 = 1,
    DVMV8_1_ONLY = 2,
    DVMV8_4 = 3
  } dvm_version_enum;

  
  /** 
    * Enum to represent snoop transaction type corresponding to
    * ReadOnceCleanInvalid coherent transaction type
    */
  typedef enum {
    READUNIQUE_SNOOP_FOR_ROCI = 0,
    READONCE_SNOOP_FOR_ROCI = 1
  } snoop_xact_type_for_roci_enum;
  
  /** 
    * Enum to represent snoop transaction type corresponding to
    * ReadOnceMakeInvalid coherent transaction type
    */
  typedef enum {
    READUNIQUE_SNOOP_FOR_ROMI = 0,
    READONCE_SNOOP_FOR_ROMI = 1
  } snoop_xact_type_for_romi_enum;
  
  /**
    * @groupname axi_generic_sys_config
    * An id that is automatically assigned to this configuration based on the
    * instance number in the svt_axi_system_configuration array in
    * svt_amba_system_cofniguration class.  Applicable when a system is created
    * using svt_amba_system_configuration and there are multiple axi systems 
    * This property must not be assigned by the user
    */ 
  int system_id = 0;
  
  /** @cond PRIVATE */
  /** xml_writer handle of the system */
  svt_xml_writer xml_writer = null;
  /** @endcond */

  /** 
    * @groupname axi_clock
    * This parameter indicates whether a common clock should be used
    * for all the components in the system or not.
    * When set, a common clock supplied to the top level interface 
    * is used for all the masters, slaves and interconnect in 
    * the system. This mode is to be used if all components are
    * expected to run at the same frequency.
    * When not set, the user needs to supply a clock for each of the
    * port level interfaces. This mode is useful when some components
    * need to run at a different clock frequency from other
    * components in the system.
    */
  bit common_clock_mode = 1;

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * Enables the Multi-Stream Scenario Generator
   * Configuration type: Static
   */
  bit ms_scenario_gen_enable = 0;

  /** 
   * The number of scenarios that the multi-stream generator should create.
   * Configuration type: Static
   */
  int stop_after_n_scenarios = -1;

  /** 
   * The number of instances that the multi-stream generators should create
   * Configuration type: Static
   */
  int stop_after_n_insts = -1;
`endif

`ifndef SVT_VMM_TECHNOLOGY
  /** 
    * @groupname axi_generic_sys_config
    * Enables raising and dropping of objections in the driver based on the number
    * of outstanding transactions. The VIP will raise an objection when it
    * receives a transaction in the input port of the driver and will drop the
    * objection when the transaction completes. If unset, the driver will not
    * raise any objection and complete control of objections is with the user. By
    * default, the configuration member is set, which means by default, VIP will
    * raise and drop objections.
    */
  bit manage_objections_enable = 1;
`endif

  /** 
    * @groupname interconnect_config
    * Determines if a VIP interconnect should be instantiated
    */
  bit use_interconnect = 0;

  /**
    * @groupname axi_system_coverage_protocol_checks
    * Enables system monitor and system level protocol checks
    */
  bit system_monitor_enable = 0;
 
 /**
   * - Determines if XML/FSDB generation for display in PA is desired.
   *  - The format of the file generated will be based on svt_axi_system_configuration::pa_format_type
   *  .
   * - Applicable only when system monitor is enabled through svt_axi_system_configuration::system_monitor_enable = 1
   * - When set to 1 the following callback is registered:
   *  - with system monitor: svt_axi_system_monitor_transaction_xml_callback
   *  .
   * - <b>type:</b> Static
   * .
   * 
   */
  bit enable_xml_gen = 0;
  
  /**
   * Determines in which format the file should write the transaction data.
   * The enum value svt_xml_writer::XML indicates XML format, 
   * svt_xml_writer::FSDB indicates FSDB format and 
   * svt_xml_writer::BOTH indicates both XML and FSDB formats.

   */
  svt_xml_writer::format_type_enum pa_format_type;

 /**
    * @groupname ace_generic_sys_config
    * Determines whether cacheline_and_memory_coherency_check should be 
    * fired as an error or a warning.If this configuration is set System monitor 
    * will flag an error if the cacheline_and_memory_coherency_check_per_xact fails.
    */
  bit flag_cacheline_and_memory_coherency_check_per_xact_as_error = 0;

  /**
    * @groupname axi_system_coverage_protocol_checks
    * Enables system checks between master transactons and corresponding slave
    * transactions for non modifiable transactions. This involves associating
    * master transactions to slave transactions which can vary from one
    * interconnect implementation to another.  For the same reason, these
    * checks are disabled by default.
    */
  bit master_slave_non_modifiable_xact_checks_enable = 0;

  /**
    * @groupname axi_generic_sys_config
    * Applicable when #system_monitor_enable is set to 1
    * Sets the allowed set of snoop transactions for a given coherent
    * transaction.  The specification recommends a specific snoop transaction
    * type for a given coherent transaction for mapping coherency operations to
    * snoop operations.  However a list of optional snoop transactions are also
    * given which can be used for each of the coherent transaction types. This
    * parameter decides whether the system monitor will use the recommended
    * mapping or whether both recommended as well as optional transaction
    * mapping for associating snoop transactions to coherent transactions.
    * When set to 1, only recommended mapping is used to associate snoop transactions
    * to coherent transactions.
    * When set to 0, both recommended as well as optional mapping is used to associate
    * snoop transactions to coherent transactions.
    */
  bit use_recommended_coherent_to_snoop_map = 1;

  /**
    * Allows the interconnect to respond to a DVM transaction from a master
    * before collecting the responses to snoop transactions sent to masters.
    * When a DVM transaction is sent by a master, the interconnect sends snoop
    * transactions to all the other masters. The specification recommends that
    * the response to the DVM transaction is sent to the master only after
    * collecting the responses to the snoop transactions sent to the masters.
    * Many interconnects however send back response to a DVM transaction prior
    * to receiving response to all snoop transactions.<br>  
    * If set to 1, the system monitor does not report an error if a response to
    * a DVM transaction is sent before responses from corresponding snoop
    * transactions are received. <br>
    * If set to 0, the system monitor reports an error if a response to a DVM
    * transaction is sent before responses from corresponding snoop
    * transactions are received.
    */
  bit allow_early_dvm_response_to_master = 1;

  /**
    *   Indicates whether coherent interconnect should perform back invalidation by sending
    * cleaninvalid snoop transaction on its own without receiving any coherent transaction.
    * A coherent interconnect may do this in order to avoid snoop filter overflow.
    * If this bit is set to '1' then system monitor won't perform snoop_addr_matches_coherent_addr_check.
    *
    *   This is because, in case of back invalidation coherent interconnect sends invalidating
    * snoop transaction - cleaninvalid without any coherent transaction. Since, this is not
    * directly visible outside the interconnect, system monitor won't be able to find any matching
    * coherent transactions and may falsely report error that snoop transaction received without any
    * matching coherent transaction so, this disable_cleaninvalid_snoop_to_coherent_match_check_for_back_invalidation
    * should be set to '1' in order to skip this check. By default, it is set to '1'.
    *
    *   This will have no effect if snoop_filter_enable is set to '0' in port_configuration
    * 
    * NOTE: This parameter will only skip snoop_addr_matches_coherent_addr_check only when possible
    *       back invalidation is detected i.e. cleaninvalid received without any matching coherent transaction.
    */

  bit disable_cleaninvalid_snoop_to_coherent_match_check_for_back_invalidation = 1;

  /** Indicates whether coherent masters are allowed to update cacheline if attached cohrent interconnect provided
    * errorneous cohrent response. If this bit is set to '0' then master will not update cache if it receives either
    * SLVERR or DECERR as part of coherent response. In this case, it is master's responsibility that it informs
    * snoop filter that the cacheline has not been allocated in case coherent interconnect has allocated the line.
    * For that reason, master will send de-allocating transaciton CLEANINVALID at the end of current transaction that
    * is supposed to allocate the cahceline but, has received coherent error response. 
    * However, cacheline needs to be removed only when master doesn't have the cacheline but, current transaction is
    * is supposed to allocate the line i.e. current state is INVALID and final state is supposed to be either UC,UD,SC or SD.
    *
    * If this bit is set to '1' then master will go ahead and update the cacheline if required irrespective of the 
    * erroneous cohrent response and in that case, it will not send any such de-allocating transaction.
    *
    * NOTE: if this bit is set to '0' then VIP system_monitor will also not update snoop_filter during such errorneous
    *       coherent response.
    */

  bit allow_cache_update_on_coherent_error_response = 1;

  /** Indicates whether coherent masters are allowed to update its cache if attached coherent interconnect provided
    * OKAY response for a exclusive read transaction. If this bit is set to '0' then master will not update cache
    * if it receives OKAY response for exclusive read transaction. 
    * If this bit is set to '1' then master will update its cache if it receives OKAY response for exclusive read transaction. 
    *
    * NOTE: This is not going to effect on behavior of the master when it received EXOKAY response.
    */

  bit allow_cache_update_on_excl_access_with_okay_response = 0;

  /**
    * Indicates if the interconnect merges dirty data received from snoop
    * transactions with data from coherent transactions of masters before
    * sending transactions to slave.  If set to 0, dirty data is sent by the
    * interconnect as a separate transaction.  If set to 1, dirty data is
    * merged with data from coherent transactions.  This variable affects the
    * way transactions seen at the slave are correlated to transactions seen at
    * the master. This must be set correctly, based on the behaviour of the
    * interconnect for the system monitor to correlate slave transactions to
    * master transactions.
    */
  bit interconnect_merges_dirty_data = 0;

  /**
    * @groupname axi_generic_sys_config
    * Controls display of transactions debug messages by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set to 1, transactions debug messages are printed by the system monitor
    * when verbosity is set to UVM_MEDIUM, UVM_HIGH, and higher verbosities.
    *
    * When unset i.e. 0, transactions debug messages are printed by the system
    * monitor when verbosity is set to UVM_HIGH, UVM_FULL, and higher verbosities.
    *
    * NOTE: It is possible to control some aspects of the transactions debug messages, the way it will be reported.
    *  - if it is set to 2 then all transactions that has address overlap with current
    *  transaction, will be reported under heading: "OVERLAPPED TRANSACTIONS STARTED AFTER CURRENT TRANSACTION"
    *  - if it is set to 3 then all transactions regardless of address overlap with current
    *  transaction, will be reported under heading: "OVERLAPPED TRANSACTIONS STARTED AFTER CURRENT TRANSACTION"
    *  .
    */
  int debug_system_monitor = 0;

  /**
    * @groupname ace5_config
    * This attribute is applicable for ReadOnceCleanInvalid transactions.
    * This will indicate the snoop transaction type corresponding to 
    * ReadOnceCleanInvalid coherent transaction type.
    * By default its value is set to READUNIQUE_SNOOP_FOR_ROCI. This means 
    * ReadOnceCleanInvalid coherent transaction type will result into 
    * READUNIQUE snoop transaction type.
    * Permitted values: READUNIQUE_SNOOP_FOR_ROCI, READONCE_SNOOP_FOR_ROCI
    * Applicable only when svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
    */
  snoop_xact_type_for_roci_enum snoop_xact_type_for_roci = READUNIQUE_SNOOP_FOR_ROCI;

  /**
    * @groupname ace5_config
    * This attribute is applicable for ReadOnceMakeInvalid transactions.
    * This will indicate the snoop transaction type corresponding to 
    * ReadOnceMakeInvalid coherent transaction type.
    * By default its value is set to READUNIQUE_SNOOP_FOR_ROMI. This means 
    * ReadOnceMakeInvalid coherent transaction type will result into 
    * READUNIQUE snoop transaction type.
    * Permitted values: READUNIQUE_SNOOP_FOR_ROMI, READONCE_SNOOP_FOR_ROMI
    * Applicable only when svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
    */
  snoop_xact_type_for_romi_enum snoop_xact_type_for_romi = READUNIQUE_SNOOP_FOR_ROMI;

  /**
    * @groupname ace5_config
    * This attribute is applicable for ReadOnceMakeInvalid transactions. If set to 1,
    * it will allow the master component to write dirty data to main memory. 
    * By default its value is 0. This means by default it will not update the main memory
    * with the dirty data.
    * Applicable only when svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
    */
  bit wr_dirty_data_to_mem_for_romi = 0;  

`ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname axi_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set to 1, summary report of transactions are printed by the system monitor
    * when verbosity is set to UVM_MEDIUM, UVM_HIGH, and higher verbosities.
    *
    * When unset i.e. 0, summary report of transactions are printed by the system
    * monitor when verbosity is set to UVM_HIGH, UVM_FULL, and higher verbosities.
    *
    * When set to 6, summary report of transactions are printed by the system monitor are
    * loaded in to new file suffix with axi_system_transaction_summary_report
    *
    * NOTE: It is possible to control some aspects of the summary, the way it will be reported.
    *  - if it is set to 2 then all transactions that has address overlap with current
    *  transaction, will be reported under heading: "OVERLAPPED TRANSACTIONS STARTED AFTER CURRENT TRANSACTION"
    *  - if it is set to 3 then all transactions regardless of address overlap with current
    *  transaction, will be reported under heading: "OVERLAPPED TRANSACTIONS STARTED AFTER CURRENT TRANSACTION"
    *  .
    */
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname axi_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set to 1, summary report of transactions are printed by the system monitor
    * when verbosity is set to OVM_MEDIUM, OVM_HIGH, and higher verbosities.
    *
    * When unset i.e. 0, summary report of transactions are printed by the system
    * monitor when verbosity is set to OVM_HIGH, OVM_FULL, and higher verbosities.
    *
    * When set to 6, summary report of transactions are printed by the system monitor are
    * loaded in to new file suffix with axi_system_transaction_summary_report
    *
    * NOTE: It is possible to control some aspects of the summary, the way it will be reported.
    *  - if it is set to 2 then all transactions that has address overlap with current
    *  transaction, will be reported under heading: "OVERLAPPED TRANSACTIONS STARTED AFTER CURRENT TRANSACTION"
    *  - if it is set to 3 then all transactions regardless of address overlap with current
    *  transaction, will be reported under heading: "OVERLAPPED TRANSACTIONS STARTED AFTER CURRENT TRANSACTION"
    *  .
    */
`else
  /**
    * @groupname axi_generic_sys_config
    * Controls display of summary report of transactions by the system monitor.
    * Applicable when #system_monitor_enable is set.
    *
    * When set to 1, summary report of transactions are printed by the system monitor
    * when verbosity is set to NOTE and higher verbosities.
    *
    * When unset i.e. 0, summary report of transactions are printed by the system
    * monitor when verbosity is set to DEBUG and higher verbosities.
    *
    * When set to 6, summary report of transactions are printed by the system monitor are
    * loaded in to new file suffix with axi_system_transaction_summary_report
    *
    * NOTE: It is possible to control some aspects of the summary, the way it will be reported.
    *  - if it is set to 2 then all transactions that has address overlap with current
    *  transaction, will be reported under heading: "OVERLAPPED TRANSACTIONS STARTED AFTER CURRENT TRANSACTION"
    *  - if it is set to 3 then all transactions regardless of address overlap with current
    *  transaction, will be reported under heading: "OVERLAPPED TRANSACTIONS STARTED AFTER CURRENT TRANSACTION"
    *  .
    */
`endif
  int display_summary_report = 6;

`ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname axi_generic_sys_config
    * Controls display of performance summary report of transactions by the system env
    *
    * When set, performance summary report of transactions are printed by the system env
    * when verbosity is set to UVM_MEDIUM, UVM_HIGH, and higher verbosities.
    *
    * When unset, performance summary report of transactions are printed by the system
    * env when verbosity is set to UVM_HIGH, UVM_FULL, and higher verbosities.
    */
  bit display_perf_summary_report = 0;
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname axi_generic_sys_config
    * Controls display of monitorsummary report of transactions by the system env
    *
    * When set, performance summary report of transactions are printed by the system env
    * when verbosity is set to OVM_MEDIUM, OVM_HIGH, and higher verbosities.
    *
    * When unset, performance summary report of transactions are printed by the system
    * env when verbosity is set to OVM_HIGH, OVM_FULL, and higher verbosities.
    */
  bit display_perf_summary_report = 0;
`else
  /**
    * @groupname axi_generic_sys_config
    * Controls display of performance summary report of transactions by the system env
    *
    * When set, performance summary report of transactions are printed by the system env
    * when verbosity is set to NOTE and higher verbosities.
    *
    * When unset, performance summary report of transactions are printed by the system
    * env when verbosity is set to DEBUG and higher verbosities.
    */
  bit display_perf_summary_report = 0;
`endif

  /** @cond PRIVATE */
  /** Indicates L3 Cache is enabled in system monitor if set to '1'. if it is set to '0' L3 cache is disabled and not used */
  bit l3_cache_enable = 0;

  /** Indicates size of each cacheline in bytes for L3 cache */
  int l3_cacheline_size = 64;

  /** Indicates number of avavilable cacheline entries in L3 cache */
  int l3_cache_num_cacheline = 1024;

  /** 
    * Allows different L3 cache allocation / deallocation policy to be enforced. User can choose different
    * modes as per underlying interconnect's L3 Cache policy.
    * ONLY_EXCLUSIVE_FULL_CACHELINE_IN_L3_CACHE :: inidicates L3 cache will hold only exclusive cachelines
    *      i.e. the cachelines which are not allocated by any masters and only available in interconnect's 
    *      L3 cache. It also enforces that only full cacheline will be allocated to the L3 cache. Any
    *      partial cacheline transactions will not cause allocation and if there is a hit that will cause
    *      deallocation of the corresponding cacheline.
    */
  l3_cache_mode_enum l3_cache_mode = ONLY_EXCLUSIVE_FULL_CACHELINE_IN_L3_CACHE;
  /** @endcond */

  /**
    * Indicates if the interconnect DUT forwards a WRITEEVICT
    * transaction downstream. A WRITEEVICT transaction is used by a master when
    * a cacheline is evicted from its own cache, but is allocated in a lower
    * level of cache hierarchy such as a system level cache or L3 cache. This
    * cache could reside within the interconnect in which case a WRITEEVICT is
    * not forwarded downstream and this bit should not be set. If such a cache
    * resides downstream of the interconnect, this bit should be set. If this
    * bit is set, the system monitor performs data integrity checks on
    * WRITEEVICT transactions that ensure that data was correctly routed to a
    * downstream slave. Note that the interconnect VIP does not have an L3 or
    * system level cache and therefore always forwards WRITEEVICT transactions
    * downstream. Therefore, this configuration attribute is applicable only to
    * the AXI and AMBA system monitor.   */
  bit ic_forwards_writeevict_downstream = 1;

  /**
    * Enables the system monitor and VIP interconnect to handle posted write
    * transactions. A posted write transaction is one where the interconnect
    * responds to a write transaction without waiting for a response from the
    * slave to which the transaction is routed. When this parameter is enabled,
    * the system monitor disables data_integrity_check. This is required
    * because a transaction may not have reached its final destination (slave)
    * when it completes at the master that initiated it. To enable data
    * integrity checking for such transactions, the VIP correlates transactions
    * received at the slaves to transactions initiated by masters based on
    * address and data.  If the VIP is unable to correlate a received slave
    * transaction to a master transaction, VIP will fire
    * master_slave_xact_data_integrity_check. If there are orphaned master
    * transactions at the end of the simulation which could not be correlated
    * to any slave transaction, it indicates that some transactions did not
    * make it to final slave destination and VIP will fire
    * eos_unmapped_master_xact check.  It is the users' responsibility to
    * ensure that a test runs long enough for all the master transactions to
    * reach their final destination.  If this parameter is enabled and the AXI
    * Interconnect VIP model is used, it responds to write transactions before
    * routing it to the slave to which it is destined, provided the transaction
    * cache attributes permit the interconnect to give a response from an
    * intermediate point. Any READ transaction that follows a WRITE transaction
    * and has an overlapping address will wait for the WRITE transaction to
    * complete at the slave interface before routing the read transaction to
    * the slave.
    */ 
  bit posted_write_xacts_enable = 0;

  /**
    * When set to 1, the system monitor check interconnect_generated_write_xact_to_update_main_memory_check
    * is enabled. 
    *
    * When set to 0, the system monitor check interconnect_generated_write_xact_to_update_main_memory_check
    * is disabled. This is the default behavior. 
    */
  bit interconnect_generated_write_xact_to_update_main_memory_check_enable = 0; 

  /**
    * When set to 1, the check data_integrity_with_outstanding_coherent_write_check 
    * considers the READONCE transactions. 
    *
    * When set to 0, the check data_integrity_with_outstanding_coherent_write_check 
    * excludes the READONCE transactions. This is the default behavior. 
    */
  bit include_readonce_for_data_integrity_with_outstanding_coherent_write_check = 0; 

  /**
    * Enables data integrity check in the system monitor across master
    * transactions and slave transactions of an interconnect. In order to
    * perform this check, the system monitor must correlate slave transactions
    * to master transactions. This process has a lot of DUT dependency as
    * different interconnects transform transactions differently when they
    * route transcations from a master to a slave. Typically, this should be
    * enabled only if #id_based_xact_correlation_enable is set, which gives
    * additional information to the system monitor to correlate slave
    * transactions to master transactions.
    */
  bit master_slave_xact_data_integrity_check_enable = 0;

  /**
    * Enables end of simulation check in system monitor for master transactions
    * that have neither a snoop nor a slave transaction correlated with it This
    * check must be enabled only if
    * master_slave_xact_data_integrity_check_enable is set
    */
  bit eos_unmapped_xacts_have_snoop_or_slave_xact_check_enable = 0;

  /**
    * This configuration sets the behaviour of the interconnect DUT when
    * routing master transactions to slaves. This information is used by the
    * system monitor when associating slave transactions to master
    * transactions. This parameter indicates that a one-to-one mapping is
    * expected between master transactions and slave transactions when master
    * transactions get routed to slaves. Two master transactions should not be
    * merged into a single transaction when routing to slave. One master
    * transaction should not be split into multiple slave transactions. If this
    * parameter is set when the interconnect merges or splits transactions, it
    * will lead to incorrect association of slave transactions to master transactions.
    */
  bit master_slave_xact_one_to_one_mapping_enable = 0;

  /**
    * Enables passive cache monitor. This allows VIP to track states of cachelines
    * in cache of passive Masters.
    * if set to '0' passive cache monitor is disabled 
    */
  bit passive_cache_monitor_enable = 0;

  /**
    * Disables the secure bit association between coherent and associated snoop transactions.
    * This allows system monitor to bypass the check for the secure/nosecure bit between coherent and associated snoop transaction. 
    * if set to '1' secure bit is considered to be checked in system monitor. 
    * if set to '0' secure bit is not considered to be checked in system monitor.
    */
  bit coherent_to_snoop_secure_bit_association_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * When set to '1', enables coverage for system level protocol checks
    * Applicable if #system_monitor_enable=1
    * <b>type:</b> Static 
    */
  bit protocol_checks_coverage_enable = 0;

  /**
    * @groupname axi_coverage_protocol_checks
    * When set to '1', enables coverage for system level positive protocol checks
    * When set to '1', enables positive protocol checks coverage.
    * When set to '0', enables negative protocol checks coverage.
    * Applicable if #system_monitor_enable=1
    * <b>type:</b> Static 
    */
  bit pass_check_cov = 1;


  /**
    * @groupname axi_coverage_protocol_checks
    * When set to '1', enables system level coverage.All covergroups enabled
    * by system_axi_*_enable or system_ace_*_enable are created only if
    * this bit is set.
    * Applicable if #system_monitor_enable=1
    * <b>type:</b> Static 
    */
  bit system_coverage_enable = 0;  

  /**
    * @groupname axi_generic_sys_config
    * Number of clock cycles interval needed before polling any hazarded address.
    * This restriction is typically needed by interconnect which may get into
    * deadlock state because of certain implementation feature, if transactions
    * are continuously sent to the interconnect for a specific address which is
    * already hazarded by other transaction issued by other master(s).
    *   In this case, if hazarded address is polled continuously then other pending 
    * transaction issued by other master sent to the same address never gets selected
    * to proceed further and remains in hang state.
    * <b>type:</b> Static 
    */
  int unsigned ic_num_cycles_interval_for_polling_hazarded_address = 5;

  /**
    * @groupname axi_generic_sys_config
    * Indicates the total number of entries of snoop filter in system monitor.
    * In other words, it specifies number of cachelines snoop filter can accomodate along
    * with the allocated master port-id information.
    *
    * If number of allocation of unique cacheline addresses crosses this configured
    * size after considering pending allocating coherent xacts, for which allocation
    * in snoop filter needs to be made, then system monitor will expect back invalidation
    * snoop i.e. CLEANINVALID snoop transaciton from the interconnect.
    * <b>type:</b> Static 
    */
  int unsigned snoop_filter_size = 2048;

  /**
    * @groupname axi_generic_sys_config
    * Enables support for tagging of addresses at masters, while disabling
    * tagging at slave. Tagging is set through
    * svt_axi_port_configuration::tagged_address_space_attributes_enable.
    * Typically, tagging should match between masters and slaves so that
    * coherency is not impacted. However, some systems have mismatched tagging
    * capabilities between master and slave. Such a configuration means that
    * secure and non-secure accesses to the same physical address is treated as
    * two different addresses in the master, but as the same address in the
    * slave. This poses coherency problems when there are
    * secure and non-secure accesses to the same physical address. It is
    * recommended that secure and non-secure address regions are completely
    * separate for such a configuration. However, some systems may need to test
    * this configuration with overlap of secure and non-secure address spaces, in
    * which case this parameter must be set so that the checks detailed below
    * do not execute. These checks are disabled by the system monitor when there are
    * secure and non-secure accesses to the same physical address. When this parameter
    * is set, the system monitor keeps track of addresses which have accesses with 
    * both secure and non-secure access types to the same physical addresses and disables
    * data_integrity_check and snoop_data_consistency_check in the system monitor. 
    * The system monitor issues a warning when these checks are not executed.
    * cacheline_and_memory_coherency_check  will also be disabled for all addresses if
    * this parameter is set.
    */
  bit support_tagged_master_and_untagged_slave = 0;

  /**
    * Indicates the mode to be used by the system monitor to co-relate slave transactions to
    * coherent transactions. There will be variations in the manner interconnects
    * schedule transactions to transactions with overlapping concurrent addresses. 
    * This variable helps to accomodate these variations. 
    * If set to 0, the system monitor will first try to establish an exact correlation
    * in terms of minimum and maximum addressable location. This is a one-to-one correlation
    * between master and slave transactions. If no such correlation can
    * be established, it will try to establish a one-to-many relationship
    * If set to 1, the system monitor does not try to first establish a one-to-one correlation.
    * It will establish one-to-many correlations, including one-to-one correlations 
    */
  int master_to_slave_association_mode = 0;

  /** @cond PRIVATE */
  /**
    * Indicates the mode to be used by the system monitor to co-related snoops to
    * corresponding coherent. There will be variations in the manner interconnects
    * schedule transactions to transactions with overlapping concurrent addresses. 
    * This variable helps to accomodate these variations. This is not expected to
    * be changed by the user. However, it may prove helpful in certain scenarios
    * where a different co-relation mechanism helps correlation better.
    */
  int snoop_to_coherent_association_mode = 0;
  /** @endcond */
  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------

  /** 
    * @groupname axi_master_slave_config
    * Number of masters in the system 
    * - Min value: 0 
    * - Max value: \`SVT_AXI_MAX_NUM_MASTERS
    * - Configuration type: Static 
    * .
    * The Max value can be overridden by defining SVT_AXI_MAX_NUM_MASTERS_(max masters).
    * For eg: The max masters can be 450 by defining  SVT_AXI_MAX_NUM_MASTERS_450.
    */
  rand int num_masters;

  /** 
    * @groupname axi_master_slave_config
    * Number of low power monitors in the system 
    * - Min value: 1
    * - Max value: \`SVT_AXI_MAX_LP_MASTERS
    * - Configuration type: Static 
    * .
    * The Max value can be overridden by defining SVT_AXI_MAX_LP_MASTERS(max low power monitors).
    * For eg: The max masters can be 128 by defining  SVT_AXI_MAX_LP_MASTERS to 128.
    */
  rand int num_lp_masters=0;

  /** 
    * @groupname axi_master_slave_config
    * Number of slaves in the system 
    * - Min value: 0 
    * - Max value: \`SVT_AXI_MAX_NUM_SLAVES
    * - Configuration type: Static
    * .
    * The Max value can be overridden by defining SVT_AXI_MAX_NUM_SLAVES_(max slaves).
    * For eg: The max slaves can be 450 by defining  SVT_AXI_MAX_NUM_SLAVES_450.    
    */
  rand int num_slaves;

  /** 
    * @groupname axi_master_slave_config
    * Array holding the configuration of all the masters in the system.
    * Size of the array is equal to svt_axi_system_configuration::num_masters.
    * @size_control svt_axi_system_configuration::num_masters
   */
  rand svt_axi_port_configuration master_cfg[];

  /** 
    * @groupname axi_master_slave_config
    * Array holding the configuration of all the low power masters in the system.
    * Size of the array is equal to svt_axi_system_configuration::num_lp_masters.
    * @size_control svt_axi_system_configuration::num_lp_masters
   */
  rand svt_axi_lp_port_configuration lp_master_cfg[];

  /** 
    * @groupname axi_master_slave_config
    * Array holding the configuration of all the slaves in the system.
    * Size of the array is equal to svt_axi_system_configuration::num_slaves.
    * @size_control svt_axi_system_configuration::num_slaves
    */
  rand svt_axi_port_configuration slave_cfg[];

  /**
    * @groupname interconnect_config
    * Interconnect configuration
    */
  rand svt_axi_interconnect_configuration ic_cfg;

  /**
    * @groupname axi_generic_sys_config
    * Access control for transctions to overlapping address.
    * If set, a transaction that accesses a location that overlaps with the
    * address of a previous transaction sent from the same port or another port,
    * will be suspended until all previous transactions to the same or
    * overlapping address are complete. When such a transaction is suspended,
    * the driver is also blocked from getting more transactions from the
    * sequencer/generator. By default this is applicable only to all
    * transactions in AXI3, AXI4, AXI4_LITE and READNOSNOOP and WRITENOSNOOP
    * transactions in AXI_ACE and ACE_LITE interfaces. This default behaviour can
    * however be overridden by disabling the
    * reasonable_overlapping_addr_check_constraint and randomizing 
    * check_addr_overlap of svt_axi_master_transaction to the desired value.  
    * Note however that this parameter is not applicable to WRITEBARRIER,
    * READBARRIER, DVMMESSAGE and DVMCOMPLETE transactions in AXI_ACE and ACE_LITE
    * interfaces.
    *
    * Configuration type: Static 
    */ 
  rand bit overlap_addr_access_control_enable = 0;

  /**
    * @groupname axi_generic_sys_config
    * Enables mapping of two or more slaves to the same address range.  If two
    * or more slaves are mapped to the same address range through the
    * set_addr_range method and this bit is set, no warning is issued. Also,
    * routing checks in system monitor take into account the fact that a
    * transaction initiated at a master could be routed to any of these slaves.
    * If the AXI system monitor is used, slaves with overlapping address must
    * lie within the same instance of AXI System Env. A given address range can
    * be shared between multiple slaves, but the entire address range must be
    * shared.  Note that this doesn't necessarily mean that the entire address
    * map of a slave needs to be shared with another slave. It only means that
    * an address range which lies within the address map of a slave and which
    * is shared with another slave, must be shared in its entirety and not
    * partially. This is possible because the set_addr_range method allows the
    * user to set multiple address ranges for the same slave.  For example,
    * consider two slaves S0 and S1, where S0's address map is from 0-8K and
    * S1's address map is from 4K-12K. The 4K-8K address range overlaps between
    * the two slaves.  The address map can be configured as follows: <br>
    * set_addr_range(0,'h0,'h1000); //0-4K configured for slave 0 <br>
    * set_addr_range(0, 'h1001, 'h2000); //4K-8K configured for slave 0 <br>
    * set_addr_range(1, 'h1001, 'h2000); //4K-8K configured for slave 1 overlaps with slave 0 <br>
    * set_addr_range(1,'h20001, 'h3000); //8K-12K configured for slave 1. <br>
    * 
    * Note that the VIP does not manage shared memory of slaves that have
    * overlapping addresses.  This needs to be managed by the testbench to
    * ensure that data integrity checks in the system monitor work correctly.
    * This can be done by passing the same instance of svt_mem from the
    * testbench to the slave agents that share memory. Refer to
    * tb_amba_svt_uvm_basic_sys example for usage. <br>
    *
    * If the interconnect is enabled (by setting the #use_interconnect
    * property), interconnect model will send a transaction on either of the 
    * slaves with overlapping address, based on the number of outstanding
    * transactions. The port with fewer outstanding transactions will be chosen
    * to route a transaction. <br>
    *
    * If this bit is unset, a warning is issued when setting slaves with
    * overlapping addresses. In such a case, routing checks do not take into
    * account the fact that a transaction could be routed to any of these slaves
    * which may result in routing check failure. <br>
    *
    * Configuration type: Static 
    */
  rand bit allow_slaves_with_overlapping_addr = 0;

  /**
    * @groupname axi_master_slave_xact_correlation 
    * Enables ID based correlation between master transactions and slave
    * transactions. This association is used for performing data integrity
    * checks, as well as for certain functional cover groups. This
    * configuration member can be set for interconnects which transmit the
    * originating master port information on the AxID bits of the slave
    * transaction. The system monitor uses this information to associate the
    * master transactions to slave transactions. The AxID of a transaction to
    * the slave is expected be a combination of the AxID of the master
    * transaction and a specific value corresponding to the master port from
    * which the transaction originated. The information on the source master
    * can be provided in either LSB or MSB of the AxID of transaction sent to
    * slave. The position of the source master information is specified in
    * svt_axi_system_configuration::source_master_info_position. The number of
    * bits used for specifying the source master is given in
    * svt_axi_system_configuration::source_master_info_id_width. The
    * configuration should ensure that the id_width of the slaves can
    * accommodate the additional information transmitted to slaves. The
    * specific value that is appended to the AxID (either in LSB or MSB) for a
    * given master is specified in
    * svt_axi_port_configuration::source_master_id_xmit_to_slaves. In some
    * cases the value that is appended to AxID for a given master may not be
    * static. This can be controlled through
    * svt_axi_port_configuration::source_master_id_xmit_to_slaves_type.  For
    * example assume that an interconnect appends four bits in the LSB to send
    * source master information on a transaction routed to slave. Consider a
    * transaction originating from master 1 with AxID 'b0100. Let us assume
    * that the interconnect appends a four bit ID value equal to 'b0001 for all
    * transactions originating from master 1. If so, the slave transaction will
    * have an ID equal to 'b0100_0001. The corresponding configuration in the
    * VIP should be:
    * <\li>
    * <\li>id_based_xact_correlation_enable = 1;
    * <\li>source_master_info_id_width = 4;
    * <\li>master[1].source_master_id_xmit_to_slaves = 1; //Specifies that value of 1 is appended for transactions originating from master 1
    * <\li>source_master_info_position = LSB
    */ 
  bit id_based_xact_correlation_enable = 0;

  /**
    * @groupname axi_master_slave_xact_correlation 
    * Applicable if id_based_xact_correlation_enable is set.
    * The number of bits of AxID in a slave transaction that is used to
    * indicate the master from which a transaction routed to slave originates
    */
  int source_master_info_id_width = 3;
 

  /**
    * @groupname axi_master_slave_xact_correlation 
    * When this is set to '1', "check_master_slave_xact_data_consistency" check
    * is skip for bytes that are already associated with another slave trasaction.
    * Default value of this attribute is 0. 
    */
  bit skip_check_data_consistency_for_already_associated_bytes = 0;

  /**
    * @groupname axi_master_slave_xact_correlation 
    * Applicable if id_based_xact_correlation_enable is set.
    * Specifies whether the bits in AxID of a transaction routed to slave 
    * which are used to communicate the master from which a transaction originates
    * is in LSB or MSB
    */
  source_master_info_position_enum source_master_info_position = svt_axi_system_configuration::AXI_LSB;
  
  /**
    * @groupname axi_master_slave_xact_correlation 
    * If set to svt_axi_system_configuration::DVMV8,it attempts to cover the DVMv7 and DVMv8
    * architecture recomended operations.
    * If set to svt_axi_system_configuration::DVMV8_1,it attempts to cover the DVMv7, DVMv8 and DVMv8_1
    * architecture recomended operations.
    * If set to svt_axi_system_configuration::DVMV8_1_ONLY,it attempts to cover the DVMv8_1
    * architecture recomended operations only. i.e it won't support DVMv8 or lower DVM operations.
    * If set to svt_axi_system_configuration::DVMV8_4,it attempts to cover the DVMv7, DVMv8 , DVMv8_1 and DVMv8_4
    * architecture recomended operations.
    */
  dvm_version_enum dvm_version = svt_axi_system_configuration::DVMV8;

  /**
    * @groupname axi_master_slave_xact_correlation 
    * Applicable if id_based_xact_correlation_enable is set.
    * Applicable if atleast one interface is svt_axi_port_configuration::AXI_ACE.
    * The value of the relevant bits in AxID for a write transaction that
    * is generated by the interconnect because dirty data that is passed
    * by a snoop transaction couldn't be returned to a master. The relevant
    * bits in AxID are the bits used to indicate the master from which 
    * a transaction originates. This value should be less than the max value
    * possible based on #source_master_info_id_width. For example, if
    * #source_master_info_id_width is 3, this value should not exceed 7.
    */ 
  bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_interconnect_id_xmit_to_slaves = 0;

  /**
    * @groupname axi_master_slave_xact_correlation 
    * Applicable if id_based_xact_correlation_enable is set.
    * Applicable if atleast one interface is svt_axi_port_configuration::AXI_ACE or
    * svt_axi_port_configuration::ACE_LITE.
    * The value of the relevant bits in AxID for slave transaction that
    * corresponds to a WRITEUNIQUE or WRITELINEUNIQUE transaction.  The
    * relevant bits in AxID are the bits used to indicate the master from which
    * a transaction originates. If there is no specific value that is assigned
    * to WRITEUNIQUE and WRITELINEUNIQUE transactions, this should be set to
    * the max value based on SVT_AXI_MAX_ID_WIDTH (ie, max width of AxID in
    * system). If there is a specific valid value, it should be less than the
    * max value possible based on #source_master_info_id_width. For example, if
    * #source_master_info_id_width is 3, this value should not exceed 7.
    */ 
  bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_id_wu_wlu_xmit_to_slaves = 0;


`ifdef CCI400_CHECKS_ENABLED

  /**
    * @groupname axi_generic_sys_config
    * Access control for cci400 interconnect checks
    * If set, a VIP will check transaction rules defined by cci400 trm
    *
    * Configuration type: Static 
    */ 
  rand bit cci400_protocol_check_enable = 1;

  /** 
    * @groupname cci400_config
    * cci400 register configuration 
    */
  // Since CCI400 configuration may be accessed by different component for
  // register modification or status update and system_configuration can be
  // used as copied object so, it must be declared as static object so that,
  // all system_configuration handles point to single entity
  // It is also declared as "rand" since set_prop_val tries to set rand_mode()
  static rand svt_axi_cci400_vip_cfg  cci400_cfg;
`endif

  /**
   * This is related to low power monitor agent, and for entry into low power state. 
   * It specifies the minimum number of clock cycles that CACTIVE should remain
   * low, before the clock controller asserts the CSYSREQ to request an entry
   * into low power state.
   * Configuration type: Static
   */
  int lp_entry_num_clocks_cactive_low = 4;

  /**
    * @groupname axi_addr_map
    * Address map for the slave components
    */
  svt_axi_slave_addr_range slave_addr_ranges[];

  /**
   * Array of address mappers for non-AXI slaves to which AXI masters can communicate. 
   * An AXI master may communicate to slaves which are non-AXI. The corresponding address mapper
   * needs to be specified here.
   */
  svt_amba_addr_mapper ext_dest_addr_mappers[];

  /**
   * @groupname axi3_4_timeout
   * When the AWVALID signal goes high, this watchdog 
   * timer monitors the AWREADY signal for the channel. If AWREADY is low, 
   * then the timer starts. The timer is incremented by 1 every clock and
   * is reset when AWREADY is sampled high. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   * 
   * Configuration type: Dynamic 
   */
  int awready_watchdog_timeout = 256000;

  /**
   * @groupname axi3_4_timeout
   * When the WVALID signal goes high, this watchdog 
   * timer monitors the WREADY signal for the channel. If WREADY is low, 
   * then the timer starts. The timer is incremented by 1 every clock and
   * is reset when WREADY is sampled high. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int wready_watchdog_timeout = 1000;

  /**
   * @groupname axi3_4_timeout
   * When the ARVALID signal goes high, this watchdog 
   * timer monitors the ARREADY signal for the channel. If ARREADY is low, 
   * then the timer starts. The timer is incremented by 1 every clock and
   * is reset when ARREADY is sampled high. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic 
   */
  int arready_watchdog_timeout = 256000;

  /**
   * @groupname axi3_4_timeout
   * When the RVALID signal goes high, this watchdog 
   * timer monitors the RREADY signal for the channel. If RREADY is low, 
   * then the timer starts. The timer is incremented by 1 every clock and
   * is reset when RREADY is sampled high. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic 
   */
  int rready_watchdog_timeout = 1000;

  /**
   * @groupname axi3_4_timeout
   * When the read addr handshake ends this watchdog timer monitors the 
   * assertion of first RVALID signal for the channel. If RVALID is low, 
   * then the timer starts. The timer is incremented by 1 every clock and
   * is reset when RVALID is sampled high. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic 
   */
  int unsigned rdata_watchdog_timeout = 256000;

  /**
   * @groupname axi3_4_timeout
   * When the BVALID signal goes high, this watchdog 
   * timer monitors the BREADY signal for the channel. If BREADY is low, 
   * then the timer starts. The timer is incremented by 1 every clock and
   * is reset when BREADY is sampled high. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int bready_watchdog_timeout = 1000;

/**
   * @groupname axi3_4_timeout
   * After the last write data beat, this watchdog timer monitors  
   * the write response signals for the channel. If BVALID is low, 
   * then the timer starts. The timer is incremented by 1 every clock and
   * is reset when BVALID is sampled high. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int unsigned bresp_watchdog_timeout = 256*1000;

  /**
   * @groupname axi3_4_timeout
   * When exclusive read request comes, this watchdog timer monitors
   * the exclusive read transaction. If matching exclusive write
   * request doesn't come, then the timer starts.
   * The timer is incremented by 1 every clock and is reset 
   * when matching exclusive write request comes 
   * If the number of clock cycles exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic 
   */
  int excl_wr_watchdog_timeout = 0;

  /**
   * @groupname axi3_4_timeout
   * When write address handshake happens (data after address scenario), 
   * this watchdog timer monitors assertion of WVALID signal. When WVALID 
   * is low, the timer starts. The timer is incremented by 1 every clock 
   * and is reset when WVALID is asserted. If the number of clock cycles 
   * exceeds this value, an error is reported. If this value is set to 0 
   * the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int unsigned wdata_watchdog_timeout = 256000;

  /**
   * @groupname axi3_4_timeout
   * When first write data handshake happens (data before address scenario), 
   * this watchdog timer monitors assertion of AWVALID signal. When AWVALID 
   * is low, the timer starts. The timer is incremented by 1 every clock and 
   * is reset when AWVALID is asserted. If the number of clock cycles exceeds 
   * this value, an error is reported. If this value is set to 0 the timer 
   * is not started.
   *
   * Configuration type: Dynamic  
   */
  int unsigned awaddr_watchdog_timeout = 256000;

  /**
   * @groupname ace_timeout
   * When the ACVALID signal goes high, this watchdog 
   * timer monitors the ACREADY signal for the channel. If ACREADY is low, 
   * then the timer starts. The timer is incremented by 1 every clock and
   * is reset when ACREADY is sampled high. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int acready_watchdog_timeout = 1000;

  /** @cond PRIVATE */
  /**
   * @groupname ace_timeout
   * When there is a read/write coherent transaction which has snoop. This timer comes into picture.
   * After address phase handshake for a coherent transaction which is to be snooped, this watchdog 
   * timer monitors the ACVALID signal for the channel. If ACVALID is low, 
   * then the timer starts. The timer is incremented by 1 every clock and
   * is reset when ACVALID is sampled high. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int unsigned acvalid_watchdog_timeout = 0;
  /** @endcond */

  /**
   * @groupname ace_timeout
   * When there is a DVM MESSAGE type transaction which has early dvm response to master.
   * This timer comes into picture.
   * After address phase handshake for a coherent transaction which is to be snooped, 
   * the timer is incremented by 1 every clock. If the number of clock cycles 
   * exceeds this value, dvm to snoop reassociate starts. 
   *
   * Configuration type: Dynamic  
   */
  int unsigned early_resp_dvm_watchdog_timeout = 50;

  /**
   * @groupname ace_timeout
   * When the CRVALID signal goes high, this watchdog 
   * timer monitors the CRREADY signal for the channel. If CRREADY is low, 
   * then the timer starts. The timer is incremented by 1 every clock and
   * is reset when CRREADY is sampled high. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int crready_watchdog_timeout = 1000;

/**
   * @groupname ace_timeout
   * When the snoop address handshake happens,this watchdog timer monitors the  
   * CRVALID (CRRESP) signal for the channel. If CRVALID is low, then the timer  
   * starts. The timer is incremented by 1 every clock and is reset when CRVALID  
   * is sampled high. If the number of clock cycles exceeds this value, an error  
   * is reported. If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int unsigned crresp_watchdog_timeout = 1000;

  /**
   * @groupname ace_timeout
   * When the CDVALID signal goes high, this watchdog 
   * timer monitors the CDREADY signal for the channel. If CDREADY is low, 
   * then the timer starts. The timer is incremented by 1 every clock and
   * is reset when CDREADY is sampled high. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int cdready_watchdog_timeout = 1000;

  /**
   * @groupname ace_timeout
   * When the snoop address handshake happens, this watchdog timer monitors the CDVALID  
   * (CDDATA) signal for the channel signal for the channel. If CDVALID is low, then the  
   * timer starts. The timer is incremented by 1 every clock and is reset when CDVALID is    
   * sampled high. If the number of clock cycles exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int unsigned cddata_watchdog_timeout = 1000;

  /**
   * @groupname ace_timeout
   * When the last handshake phase of read transaction ends, this watchdog 
   * timer monitors the RACK signal for the channel. If RACK is low, 
   * then the timer starts. The timer is incremented by 1 every clock and
   * is reset when RACK is sampled high. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int rack_watchdog_timeout = 1000;

  /**
   * @groupname ace_timeout
   * When the last handshake phase of write transaction ends, this watchdog 
   * timer monitors the WACK signal for the channel. If WACK is low, 
   * then the timer starts. The timer is incremented by 1 every clock and
   * is reset when WACK is sampled high. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int wack_watchdog_timeout = 1000;

  /**
   * @groupname ace_timeout
   * When a barrier transaction is initiated, this watchdog 
   * timer monitors second barrier transaction of the channel. 
   * If the barrier pair doesn't appear, then the timer starts. 
   * The timer is incremented by 1 every clock and
   * is reset when barrier pair is sampled. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int barrier_watchdog_timeout = 1000;

  /**
   * @groupname ace_timeout
   * When a DVM SYNC transaction is initiated by a master on read channel,  
   * this watchdog timer monitors associated DVM COMPLETE transaction on the snoop channel. 
   * The timer starts as soon as DVM SYNC transaction is received from master on read address channel
   * The timer is incremented by 1 every clock and is reset when 
   * DVM COMPLETE is received on the snoop channel. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int unsigned coherent_dvm_sync_to_snoop_dvm_complete_watchdog_timeout = 0;

  /**
   * @groupname ace_timeout
   * When a DVM SYNC transaction is received by master on snoop channel, this watchdog 
   * timer monitors associated DVM COMPLETE transaction on the read channel.The timer 
   * starts when DVM SYNC transaction is received by master. The timer is incremented by 1 
   * every clock and is reset when DVM COMPLETE transaction is transmitted on the read channel. 
   * If the number of clock cycles exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int unsigned snoop_dvm_sync_to_coherent_dvm_complete_watchdog_timeout = 0;

  /**
   * @groupname axi4_stream_timeout
   * Applicable when svt_axi_port_configuration::axi_interface_type is AXI4_STREAM
   * When the TVALID signal goes high, this watchdog 
   * timer monitors the TREADY signal for the channel. If TREADY is low, 
   * then the timer starts. The timer is incremented by 1 every clock and
   * is reset when TREADY is sampled high. If the number of clock cycles 
   * exceeds this value, an error is reported. 
   * If this value is set to 0 the timer is not started.
   *
   * Configuration type: Dynamic  
   */
  int tready_watchdog_timeout = 1000;

  /**
   * @groupname axi3_4_timeout
   * Bus inactivity is defined as the time when all five channels
   * of the AXI interface are idle. A timer is started if such a 
   * condition occurs. The timer is incremented by 1 every clock and
   * is reset when there is activity on any of the five channels of
   * the interface. If the number of clock cycles exceeds this value,
   * an error is reported.
   * If this value is set to 0, the timer is not started.
   *
   * Configuration type: Dynamic 
   */
  int bus_inactivity_timeout = 256000;

  /** 
    * @groupname axi_generic_sys_config
    * Array of the masters that are participating in sequences to drive
    * transactions.   This property is used by virtual sequences to decide
    * which masters to drive traffic on.  An index in this array corresponds to
    * the index of the master in slave_cfg. A value of 1 indicates that the
    * master in that index is participating. A value of 0 indicates that the
    * master in that index is not participating. An empty array implies that
    * all masters are participating.
    */
   bit participating_masters[];

   /** 
    * @groupname axi_generic_sys_config
    * Array of the slaves that are participating in sequences to drive
    * transactions.   This property is used by virtual sequences to decide
    * which slaves to drive traffic on.  An index in this array corresponds to
    * the index of the slave in slave_cfg. A value of 1 indicates that the
    * slave in that index is participating. A value of 0 indicates that the
    * slave in that index is not participating. An empty array implies that
    * all slaves are participating.
    */
   bit participating_slaves[];

  /** @cond PRIVATE */
  /**
    * @groupname interconnect_config
    * Array that represents the domain configuration of the system.
    * Each item represents an innershareable/outershareable/nonshareable
    * region with the corresponding masters and addresses.
    * Use the following methods to configure this easily:
    * svt_axi_system_configuration::create_new_domain()
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when there is atleast one interface in the system
    * with svt_axi_port_configuration::axi_interface_type set to
    * svt_axi_port_configuration::AXI_ACE or
    * svt_axi_port_configuration::ACE_LITE
    */
  svt_axi_system_domain_item system_domain_items[];

  /**
    * @groupname interconnect_config
    * Note: This use model is currently being deprecated.
    * Please use system_domain_items member.
    * Array that represents in the masters in inner domain.
    * Each element in the array represents a single inner domain.
    * The a bit value of 1 indicates that a master belongs to an inner domain.
    * As an example consider 5 masters in a system. Consider that masters
    * 0 and 1 belong to one inner domain and masters 2 and 3 belong to another
    * inner domain. This will be represented in the variable as:
    * inner_domain[0] = 5'b00011;
    * inner_domain[1] = 5'b01100;
    * Applicable only when svt_axi_port_configuration::axi_interface_type is AXI_ACE.
    * 
    * This member is used by Interconnect VIP and System Monitor VIP components.
    */
  bit[`SVT_AXI_MAX_NUM_MASTERS-1:0] inner_domain[];

  /**
    * @groupname interconnect_config
    * Note: This use model is currently being deprecated.
    * Please use system_domain_items member.
    * Array that represents in the masters in inner domain.
    * Each element in the array represents a single inner domain.
    * The a bit value of 1 indicates that a master belongs to an inner domain.
    * As an example consider 5 masters in a system. Consider that masters
    * 0 and 1 belong to one inner domain and masters 2 and 3 belong to another
    * inner domain. Consider that masters 0,1,2,3 are in a single outer domain
    * and that master 5 is part of the system domain. 
    * This will be represented in the variable as:
    * inner_domain[0] = 5'b00011;
    * inner_domain[1] = 5'b01100;
    * outer_domain[0] = 5'b01111;
    * Note that the system domain includes all the masters in the system.
    * Applicable only when svt_axi_port_configuration::axi_interface_type is AXI_ACE.
    *
    * This member is used by Interconnect VIP and System Monitor VIP components.
    */
  bit[`SVT_AXI_MAX_NUM_MASTERS-1:0] outer_domain[];

  /**
    * @groupname ace_config
    * defines starting address of each exclusive monitor.
    * User can simply configure as start_address_ranges_for_exclusive_monitor[<exclusive monitor index>] = < starting address of exclusive monitor[<exclusive monitor index>] >
    * Example:: start_address_ranges_for_exclusive_monitor[2] = 32'h8800_0000; < starting address of exclusive monitor[2] >
    */
  bit [`SVT_AXI_MAX_ADDR_WIDTH-1 : 0] start_address_ranges_for_exclusive_monitor[];

  /**
    * @groupname ace_config
    * defines end address of each exclusive monitor.
    * User can simply configure as end_address_ranges_for_exclusive_monitor[<exclusive monitor index>] = < end address of exclusive monitor[<exclusive monitor index>] >
    * Example:: end_address_ranges_for_exclusive_monitor[2] = 32'hC400_0000; < end address of exclusive monitor[2] >
    */
  bit [`SVT_AXI_MAX_ADDR_WIDTH-1 : 0]   end_address_ranges_for_exclusive_monitor[];

  /** @endcond */

  /** 
    * @groupname ace_config
    * if it is set to '1', exokay_not_sent_until_successful_exclusive_store_ack_observed check 
    * is executed on per caheline basis.
    * If set to '0' then the check will consider exclusive store transaction targeted to any 
    * cacheline that is yet to receive ACK i.e. regardless of the transaction address.
    */
  bit check_exokay_not_sent_until_successful_exclusive_store_ack_observed_per_cacheline = 0;
  
  /**
    * @groupname axi_system_coverage_protocol_checks
    * Enables AXI system level coverage group for master to slave access. Note
    * that to generate AXI system level coverage, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */
  bit system_axi_master_to_slave_access_enable = 1;

  /**
    * @groupname axi_system_coverage_protocol_checks
    * Applicable if system_axi_master_to_slave_access_enable is set.
    * If set to svt_axi_system_configuration::EXHAUSTIVE,it attempts to cover all
    * possible combination of master to slave accesses and hence system_axi_master to slave access
    * covergroup is used.
    * If it is set to  svt_axi_system_configuration::RANGE_ACCESS then it equally
    * distributes all possible master to slave access values to fixed 16 different bins 
    * and uses system_axi_master to slave access range covergroup.
    * However, if total number of accesses between masters and slaves, is less than 16 then 
    * it attempts to cover all possible values and hence uses systen_axi_master to slave access 
    * covergroup.
    */
  system_axi_master_to_slave_access_enum system_axi_master_to_slave_access = svt_axi_system_configuration::EXHAUSTIVE; 

  /**
    * @groupname ace_system_coverage_protocol_checks
    * Enables ACE system level coverage group for concurrent ReadUnique and 
    * CleanUnique transactions from different ACE masters.
    * Note that to generate AXI system level coverage, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */  
  bit system_ace_concurrent_readunique_cleanunique_enable = 1;

  /**
    * @groupname ace_system_coverage_protocol_checks
    * Enables ACE system level coverage group for concurrent outstanding transactions 
    * from different ACE masters with same AxID and same interleaved group id.
    * Note that to generate AXI system level coverage, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */  
  bit system_interleaved_ace_concurrent_outstanding_same_id_enable = 0;

  /**
    * @groupname ace_system_coverage_protocol_checks
    * Enables ACE system level coverage group for concurrent overlapping 
    * coherent transactions on different ACE masters in the system.
    * Note that to generate AXI system level coverage, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */  
  bit system_ace_concurrent_overlapping_coherent_xacts_enable = 1;

   /**
    * @groupname ace_system_coverage_protocol_checks
    * Enables ACE system level coverage group for coherent to snoop transaction
    * association.
    * Note that to generate AXI system level coverage, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  bit system_ace_coherent_and_snoop_association_enable = 1;

   /**
    * @groupname ace_system_coverage_protocol_checks
    * Enables system_ace_dirty_data_write covergroup.
    * Note that to generate AXI system level coverage, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  bit system_ace_dirty_data_write_enable = 1;

   /**
    * @groupname ace_system_coverage_protocol_checks
    * Enables system_ace_cross_cache_line_dirty_data_write covergroup.
    * Note that to generate AXI system level coverage, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  bit system_ace_cross_cache_line_dirty_data_write_enable = 1;

   /**
    * @groupname ace_system_coverage_protocol_checks
    * Enables system_ace_snoop_and_memory_returns_data covergroup.
    * Note that to generate AXI system level coverage, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  bit system_ace_snoop_and_memory_returns_data_enable = 1;

   /**
    * @groupname ace_system_coverage_protocol_checks
    * Enables system_ace_write_during_speculative_fetch covergroup.
    * Note that to generate AXI system level coverage, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  bit system_ace_write_during_speculative_fetch_enable = 1;

   /**
    * @groupname ace_system_coverage_protocol_checks
    * Enables
    * system_ace_xacts_with_high_priority_from_other_master_during_barrier
    * covergroup.
    * Note that to generate AXI system level coverage, you also need to enable
    * AXI System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  bit system_ace_xacts_with_high_priority_from_other_master_during_barrier_enable = 1;

   /**
    * @groupname ace_system_coverage_protocol_checks
    * Enables system_ace_barrier_response_with_outstanding_xacts covergroup
    * Note that to generate AXI system level coverage, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  bit system_ace_barrier_response_with_outstanding_xacts_enable = 1;

  /**
    * @groupname ace_system_coverage_protocol_checks
    * Enables ACE system level system_ace_store_overlapping_coherent_xact covergroup 
    * when two master issue coherent transactions to overlapping cacheline at same time
    * Note that to generate AXI system level coverage, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  bit system_ace_store_overlapping_coherent_xact_enable = 1;
  
  /**
    * @groupname ace_system_coverage_protocol_checks
    * Enables ACE system level system_ace_no_cached_copy_overlapping_coherent covergroup
    * when two masters issue coherent transactions to overlapping cacheline at same time
    * Note that to generate AXI system level coverage, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  bit system_ace_no_cached_copy_overlapping_coherent_xact_enable = 1;

  /**
    * @groupname ace_config
    * Enables the get_dynamic_coherent_to_snoop_xact_type_match callback in the
    * system monitor that allows users to set the snoop transaction type
    * corresponding to a coherent transaction type on a per snoop transaction
    * basis. This callback is useful in situations where a multi cacheline
    * coherent transaction results in snoop transactions where all the snoop
    * transactions may not be of the same type. For example, for a WRITEUNIQUE
    * transaction, an interconnect may choose an implementation where the snoop
    * corresponding to the addresses upto the cacheline boundary have one type
    * and the subsequent snoops have a different type. 
    */
  bit dynamic_coherent_to_snoop_xact_type_cb_enable = 0;

  /** @cond PRIVATE */
  /**
    * @groupname ace_system_coverage_protocol_checks
    * Enables ACE system level
    * system_ace_downstream_xact_response_before_barrier_response covergroup
    * when a barrier response is received after WRITENOSNOOP and READNOSNOOP
    * transactions prior to the barrier from the same port have received a
    * response from the dowstream slave. This covergroup is enabled only when
    * id_based_xact_correlation_enable is enabled
    * Currently not supported
    */
  bit system_ace_downstream_xact_response_before_barrier_response_enable = 1;
  /** @endcond */

  /**
   * @groupname axi_addr_map
   * Enables complex address mapping capabilities.
   * 
   * When this feature is enabled then the get_dest_slave_addr_from_global_addr(),
   * get_dest_global_addr_from_master_addr(),get_dest_slave_addr_name_from_global_addr,
   * get_ext_dest_slave_addr_from_global_addr and get_slave_addr_range() methods
   * must be used to define the memory map for this AXI system.
   * 
   * When this feature is disabled then the set_addr_range and translate_address()
   * methods must be used to define the memory map for this AXI system.
   */
  bit enable_complex_memory_map = 0;

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
 
  /** @cond PRIVATE */
  /**
   *  Stores the Log base 2(\`SVT_AXI_MAX_NUM_MASTERS),Used in constraints
   */
  protected int log_base_2_max_num_masters = 0;
   int num_ports_per_interleaving_group[int];
   local int interleaving_groupQ[int];
   local int ports_per_interleaving_group[][$];
   int lowest_position_of_addr_bits[*];
   int number_of_addr_bits_for_port_interleaving[*];
   int lowest_port_id_per_interleaving_group[*] ;

  /** @endcond */

//vcs_vip_protect
`protected
(T81QU1Y?PdbU3d3&,SW/-f6<=Cf9b,QS1GM:A5dZg<XTF8/NQ&4/(-IT8/56g42
MdOgGT)B5L5=0_f<g-KGBW3c?ff>)AU3+B-7^&;21Q.N\f-HW);2N7a:VI6c)-&C
EeW6&W1/@F&1<cSB]bIXKa,9d#Id38D2aW3QBDJ/I,?QH4S_4<7,?]&.aQSFc<)c
@-eF&,d[JOX-B9G4_C>T1P<9P^U(cOJ/La,NM(97VZ8c&+<d6/V^+@M7CFUH.)<a
3;#DOMeH@_]ZWfP;]XX4E,g,0ZOdeHPC<Q#UC)&VQ.6#V#=BF.4;3Y\3Z@c1KAd=
T+DSc5S6N.BgA(e:]0/a@N]]aF,K0&)6aXX[b-@L0-^Y\W;Mf#YQgM(=3LK5U>,d
-;DZL([E;@1+).+g&0B&AE0GKKCTUSNeLI@73I>])A(AUON\a4ZIGeP[IXU5eTL0
aAe9_gFF\@F:/#GB_e\(d[/fSIg@>)6IgD>N[[80g54A6].f(<X[,Y0KN91>E<2+
,gKH8&FQ.IKB(^g2P3]&,W-b7>.7HbRXT,>/a>S>Qa@I\eI=ST9O0JH.P,?D<IW5
GTe^,F6>EH.@\ZY<66E-6</@--M#1\7G^J:,Ea9@U1Gb1@.8[QHNNRdEf8@2_SBT
,QS6.PDZ)DV=>VN-EKg7/b1[-^K4L.HWa9fFR#-=3F_@a1gZC-VLXO9S^KK?[#Y8
86.G&E4LI_c_XYN>K^<@O7?/7H-L3&1LD1DFU=1bOY@R?bT^=MgDf\PFQ_()V#;I
-MUCU<gLWY6HCS_:&C@>\HHITA1M-??DF5=32R8.I[UR;Y\C5U.3aL)Mf<SV+.e(
BWIG2W8D#:OX0=&UL?G,fKeJ\)&#3P&^Q[CUTZIGM.B<YZ?f9L6?c]>d]@Ka=4GZ
G/+BJ]758OfQP4N-6\+\DXA,U_1T9KN,ge6eE?#1A0<XdKTDAC\]b=\0-3Q:@BdO
PKbA5:59KZ6;AR&S3_73;RSERGU:-b>M,>\,6Q=JJ.6_@eF3846^7<\&M=R6/1NX
<,YYIP,6,B=:,@a93_)gQA;5E-@[O\:.14e.@J;_;NZGDf2@d,VIQH107,^JHY9U
572<e;6T_1gG/C<Q<RM[Q7K5KNBf5QW@IZB+Vb;973\V)?>=H+WDML/^)A->d9eV
Z#.Sg:3fEcPcH\;[FW3aHG?@DV9(b=KCEYDIHfR_-HFUQ41E;FY(RSV^cg\EcQfE
Ig8[VOC7N/O@1:Xc4-86BP]6dXS4]Wf5GW8=R^\.#NM0NTY#Z0fd9,Gb[MDSBT[3
Y^GW>E06/Oa@7>L/S(]d83Z,MO;>KMX<M1d6[0.[U<C1N>-,113Z\A1LS,0]VV>6
_/cR@=3WJMTQ.<FLF?Pf/>dfK(0cW=):59RZNRB]?@Gc5?Rf&Ea-.A&>LME-DEN1
,bNd/MIYS1T92aVTeO#C1A;SM(3Lg&Ja2NS:&Z>4ceZBaQTEL#JeM8N:GO>]/7b@
cM>C)BZ8bFDfK@P7gUIZN._2HZBE_]CeO]^=&(8H[3GW^,:MK[g]((Zg#[+EJ1FV
C-RHWCB-E@BH6.5V6N[H7f-c1X601C67-d@7UP<PL0TbBOW66N=E8<bH\2S8;,Wg
94D@FUW(KO/e>aOWME<_4&Sg9Ldc+5HOK?eUKHPeC8=X.FOCPZb4K&SA4IQ:b#bF
F+U#0L#F0(9Y=W-)=E-E1GRWa6GOI,U:6G?>gURN>A9\.7C&&gD@Y[>WN\I[XQ?U
-N)0<FB(=e8e.)O7)JYD?8Q)1>G#3eU(GLCFf,_DB3+3(<X]QFBaI1<f:D4=E64^
[PR=+RDXgQObQf_P:+FY@^e)5(_J)3CMLR]N0+cPISE=bDF#6MK>Z-HFOUV7(&#X
FWOI0C]3g+,JbDT8[c#5N22Pf+/(NNO>Ve>6e0[KI/=(gedCKU_(\DE0D.TO.9Jg
eO4b==f4MIgWcKFW[]T<SLeIMJY3)_O\2>ZfZ]4.gfXBU+>J8>OdZLBU2;HHd7HL
_F0W04DH(^^>e7/d0(E62WPF^g?KIJ)1ZTP&X#gPADLP84Cb;BYTBX0d]CI?QV(U
>,,10(=7L]NS:bG4eeXH3:/A/Z/IYaeJ^6>&0H(7:64b)>@GBASCE>gR?^#VX#]W
F?[P3EU@B?V=c&b?G&21)KLEOeQa.B=@5XFb1]<YT]EDSDI9(1D60CVN9L1[1?0>
)gZ:NgK=VH<<H+4<?W6+2WJ<WM0P[V8.@Z[U27E<F@Of/[C_UJ_Q8fOR+P>4H09,
e8?5]_\a,ZRCQYX#;I2)=+>)CX^V)D_Y@S?R7VKWdPGNg7\\W4,\6)@-Y;TQTaNb
bgS]D5eW@H_>8[PJ.#<d_;/H3Lf1RJ)>\(_CHSafe4J/GCAP5FTI6AB^H1(69Cd9
O0/R=,dG.E>_NWaMBFQM+=L(530@LBA9Y)^d&::+,F/Q&7cK]dL,3aIH>.F15O=P
RCQF1.->=BGAG8NCR^cO+R6R89JICb&-GTD&EBY-,;L:;16:R6H2N=L8GBZN\S?3
+;IST?)AK,7e.;6\X=Gdg(U.@=X5<7?g=I+:Gf>ZLgC,S/D?>H=QXS0W+MTH9W(K
/0WFT.Z]a5#NQ?VEe_E]D?[REV=37N^/;6DHF?cZN]^4#I.AcRTM1d;dYMRTOC#<
XL#6P&RF>5B0DW)+a&XF47]6F0Xc/][;3JYP--\,[c(./B8:0dba6[US=\f2(WWe
YbA_ECg@dGKA(G;=Q)dC).:0c1EYA1?>cP8XgbH@/Y_B;D=WDNe?/f?W)6TH8D24
&U;eY4;eG_)N?EF7G7O[IG\eDGLcLXeHe5HZNH(_X-7W6KM&-^>4@QAZSgS:OA_b
]=?-.Ref<W>eP+3[+//][(R]8(XeJXVW[-V/88LF#K_?4d:CZ;154+dXb93@K[c4
ICZS+X(4E(H-]Yfb(<&@b?7#-c]?H.EQ/V<e_>5BT-]X2EUfb_d,8<,EOJ:=3])N
M7T;010(=9D4RXXL1Z;5OEe:VQU_BWcf/d?+e<>.LX9GTD6\3fE7X-gPPMV-U22F
#IT<_,K9b.+b:YfVSHN=2EL=#RTJ]:8\<8[?B\2I&g6g9Ne_X5,>#00?GObI1R9.
:@9X][2IL=IEgA\:N_#?0,9b-MSG--eRX^/.O+/S[8OQ4-&7GGC#U1af>5&8QLe0
PJ^/0g5M^3;M4^Z+QJMA@=EE3KIHW^>?.=)BDaUb=QT7[KeOH5_#JL_0cX6Ff>@2
&,0];N7M7S<BG8\76AaG/Q#<)\6U\(534T3(gdada2>0(QdTa8Kbc]#>@g@->_47
)QJTXOf/cSR;CPI4Q-f^^>PY?9D>R)A;L#ZX+dUZ;T[[Nb&;22#T<5S#a]3F2U?4
B?1fHGI.#ANHEb/HOZI]cW3<821.+E<[R])KGNN>A^f&)NLb14B/VgCa75.4FXY<
JVMGe8J^E0<g?2KNRWOI(JZKB_aO-H)G<1<DH[;PTN26Z&eOf81KET>9Yc_._4Z_
LR\aL1]&aFa3S^dSR7?:TJY)SP5dYYbC\ER7>E&QU=\N67,6,;DK=,_fZQ,#@EM]
2:S47L?L2T5;9d\[_==cJ@X+SN&OCba+G>^<=Z>W>-,:/WJO9@Ac3_;dfJ.LRDN:
TYb>#6[fD71MODC?KI6Z@2e/2QQIER=JZ(G+]#P]4;ecf,/e4NT=5CX_G=7Q.@gS
U+F3[(>Y->UXJ==DC[EAX34#2Y_.DgHY8MV;2/<V.)d[9;df@;;ZCS13UIR#A,VL
:[6(:)(HYQe023\]aK@8R?>&O@gQY1J20EMTdD:3YO8=OI?5-Y=g#-&LbCZ&92M0
RbfM-fXU]FL6T>g/?f<e.X7K:F<Ia-,5eCC3JZfG,6cIZ.-91d5#2\W.f_X2&ARa
_MG@Y:](=c_E\_a&#GS9_-9_/I\)aOA0OcC,NF#c,G<GU^.;VW+[@.fCZ\JbISHf
XH48+1,bD+WK8WL45PR#P-B#gDKGYH@0@V.5fXe#Ig5C0KGXO,[BXS192/2JH>9O
T.XJ]KXF^S<0@HFZ^H]Ag5dT<_+,F1W9[B(VfA9GCfLTX+TS=S91+=)8[FT\,,+U
_gUgK0d(<bQBSLU4_acHP+35M(HVfIQQc8NB]UKN(::8gDQ;ePE&8NFMB4@<,VGc
1&#aCO1U5[IHPVG7I0E-<2H7BE\+)^5KfUcG0T08R+@[WV-_d^QJ;0-S=?.<d(GI
QQ?.1<2R-S@4I2I#FHX0G_V7I/C(GLY4ecd#K?@\;8>G&[9g9CFBU.B;(^[-7(59
@)_+-b8/<@GP83f(<fE^KYaNdYH82ND\X1\0dRaU)]DPVK[\S[L?;:W.2bGP0ePL
<Fa8fZVSKA1>^XR]D/[^f_QeA=1>HcF+gJQ20<;1U6ggGb1MZVM2)1_IFTA)&cWS
D;Y3D+GOK2BX0YN.K#eQ?BV=fG?8DT=-(>BK#eFKD0d]MA8;BD=<gJ:9V-7CPM_E
[.d_6DP61:[/Hd_664HUUc6e1,9<>Na36E3.?^8LW\V7H9dC9c27b,@Q(3Z/R:/P
4>0JOE<RC[WSXG4UMLIC_JFfNV-LfDMC)Uc+bBSG)Z0#J1TM<YF[N0ZWHET82\(P
?/[fO>8C)Ue+_<E<]Z&DF5HI=ZVI:(+6Q[-RL/U-F269G/TIb2X)SEc1?-TdOUFQ
Uda#-65>gTH&^ZKa_4ON=O45G-HMA/3TD]Nc<(_91fUS<Q-75Y]#_b:..aeLXRL&
Q#bJZ)P9/R.,9#D2EBfXE94R\_Sc+4F/4+_,a(\da@f;[Hcb5Pd+X&<e,6&Z:G_d
3=HYRb=:(D3+>=N>H=BEYS7B<Y0Q\P^+I\QKTVF^05XZ4YSfAG[SGg;4Q4P5<P9_
2,V<7#4YXT-8P^:e^\J#KSCTCD:.WM9->H6NHK#\_M<O<]GX1,0Cdc()._)d;TY#
FaKa=WCSa#-+9L@8E?dNPA[M;,#IM(gRd/\;;Tg&YPNG]L3eWW.B^G)1_[6ga=Q\
K[SH\a=P7@=2T)_Y^XI>]b1dVcJEJFZX-]YdMgLT]1:E_2/+TM?5:K2ZXR;9U6bf
I90X5.bCI65>O_;1-4<#N9dKcc9N@Q2=WH5C>:WJQ4.W4+FS^\FJ19:;.KQL(+X0
;VVe4OCIABF#GV]9/\I9aS>[,R;^\U./MU1-UdMd@GZK/:V6^g[bI6KC^#=5HcUP
5YcA9I7HPMM7dLBW4P^,NJ7;2H&;-AIEC)SY33@YHgcRdN+UcdI#-/B_Ge^:eLP9
_Ub\WCffa5-T<DaQS\A#PNV_(9<ML-.6^:HZA>c2X/Z?CDAC\:;Te;L0[K;/gX^3
8b4@)JDcJ8[[U53]N0ce>edF8&_BR&]/:A;Y>OU>0EQW4UA(878LGDI&8M>2YGZ)
Rf;6@H.8LW<6DZ.RC2>.U0-+,90X,#J[6g.b+<^f,OPMN;>2VYPS#YZ/<YKWCTN4
.QX/MCZN>5J,f9f@-Q,)=J[N+^+/=7+Q5R_c&<[>VT\]09:fR;?2L#RR-N@^c:O2
F-LNMb(F#f6Cgbd@?>eW(9?52[W&IRb.Sa3G]Zfe@g=8_9Ldb:L(?(>;L\G,\134
a3T<#9;^TI\G:T-UB-#VPOaQ[.08GV4D=Ie:_aK;5e[ZKfPd_;QE06OO7MO1)7PX
=F;9@.LQf<Y,Q-Ia3:^+6(3fRNRX7Qc(6Y+eW7;A/D-+?.>7@,;,b5WMd.8ca^@/
L__2\^(J<ME1=PI7Y#KedG:7#RW6EgK?C(:N\<-8?HT@^<#U7V:@\/0KcFZ.;L>G
=7+[4X9Ae?M5.+[H5e@>INQ<DdPeLG+POT>M?:S>U59<+GMg,BB@Pf(\;VN/@WN>
H8OfE]M2619a?Q/Q(bT@ME6eO\F^TLFYd3&T3_Y/VIYW<A9B96A,I)18@?<fJ-,D
=aI6Y]0+6ON9ga,dKgZ^S1LUc0H9)&g7dPc>8(1^UcKTA)SUJ:0+8XdbK-YMGJc=
X8DDG=CS^6B)XOc7R>fWA-2e6N4KWb-[S4Ld@=+0L006LEE)bZX0J+:GFWf^D;>;
ed8VYM/1gVFX2a6=(aQL^L3=-\A5U,EgU:/SbA93=9aSF8+M4O>gK0(I#@GDE]ZT
SDB&@K0Hc_SEHTG@#Wad55B-.Y_d,B=3aDM5)QT5)&:].QV8]MO[^J?c\,SbSRB1
\/L<4>e2]ccN+5NFD69?,eNIJXTT&]@Y+\gdDQ/.VYZABfJdW&]74dEE[-[dO94Z
cNDAAQ:T+<T4C9GZ6?@;?Ca6^C1I73FOd_Y6K[Q#08:ZFU9P5H/0F5e90TNcCMLG
cTLAQN_#2:X+(3BbQK+\g0F[]acVX@/IPV2@KI1WC,4YOKM<F_-I4=6GbA_#>TVS
(5IJJ.D55T]>.8NO)YLQNV7H:<P3,S9&S7PYQ.#<dJe^R]VVC=^7X-GF-?NUa)&=
bY+JSO.<C3YG4=T_;)L;)_Ca@HE,W,2cK7>g>gQL@AMZSI2LMb+ED1:1M8aX.@eI
2Id@2K(@+JeQQ6H<1?gEDW(R\>d(.Rb(c,4HZQI,_+D;-XfGV0[,OSf4290J_]][
dHGa)5G@&#2XUNV=QfL@aZH.R=4M=Zg0HVR3-[c?O>.A0JVR_AgRXHgTY3WW^dVM
BaO:+U.D/g[_65@9@.85FeM@c&INA[6R0/V6IM:5#gBF;a(.+MO1;2^#?\cS7+;L
0&8a=DeH13?NH@S>\aH#(D#),aKcgUg^fG;P]<YXQ32ZQ&VbS.@0W\2(E67(PS?Y
KDI<#SL3g]=PIM_ZG)2J>_J1@82WI4DC#FZ[.8e9M[-HXYa5dG#cXSLMTEMd:93>
]#8G6JfW&Q\,E79VMaR/UG&88Y9?F8&2HgGIMfZ?d4=B2RFMfO0(409bA(2VIDAc
c^2Q?LX=:1_;YG8&.),6UPeO&>16\^UB4[gg6_QS<Rf\]6R^W\MFeFXC<9MLB,L;
DJ&<\d?3H8G,9=A/E;NZFR<2cZe908CKGF-=_)(S(9)<36W@V1;=?Z(1JR;+/U?f
.__DN3B@c.^0T3O=>VP1NIY>7:2W1A^DQDcbf>[E6&&bDZ6bOW@?UGN:1IA_OB&e
a7c1F\+/3cX@40]c-1VF8-:@#Z)6[.UCR?SV3:ee,/Q^15)&AQ<:NK^Ug&VIMa]P
O(f/NKW#K^CK)3+@X.W-(QX/1/VF15TGHbID,2K3cZKKWS,>d4-S?^I7@:,A@P6I
3ZXAHZKPE4L[X8GIeeV81V=?[M28g6eCIIGQS67P?:>Ya=F?GV@PgdCKKP_#]SfH
UN&7QSO5TL<D\\N<H:Ha6B5PBK]DX,559R)+YM5O5@KW^I^QL>RScOF-@<\#XF..
S1F?AFC:2eGdgPY^C(&N=\#)A+VQU2:PC6gEYH\fSf-T+E4;6RGa;Q4-3R..C^]=
8&][<&;MZee\Q&0<ZTVTMOeaYU4T(H6dCPO?O4W^ZR@++e@e>/U:b50,AN3d)U2F
fb&.<:O))&AKB<;,9Y:^Q6b4Ue?\SIBRA(V+&]1QEF75fSQ?0/6,Z4C^9W;AC,_J
e:BQ,c4>d;J@VK9A_P]^;NBb2WA9#9A<g4G#fG3#Lg1F#J?KA02[I[U&;+2;[2-<
+90^eK.6K@USR[RZgJ(THY0(UDK0L#2>7WLVGT.e?2UDd53eO#V#AEXG1O1)?J2Y
Ac4S8Ha-@;G2eK+R^5BZ\+Yb9:GP:H@E=K&[&gE\WQb\QN2U?BXY0>)[?cZ8?5,d
T+8KGC_:3L-O^[PF&681[>_K-GY_P2ZR7_<E2@d)XX7G>ZNR:8TV^VVK7=2ZJc]X
V7>GSRF13gCU4C&>FJDFZF&DA-#3\7E#58.T?F>7?U@T3<D;[#e^=EeWO=2XO1gQ
T&QBB@,@OK?#T#[gYf,\U(F-5g(_THbW6AV>fA8IcU<GR,HPcJCJ;41X@4XP8@-?
4SWW<6Vc[RVH=.GEW4f[_D>+PCNg<9QUHB7cG)a_T#K<:PbH)5#K+(;c@]I7RH;2
+3)]IJS<K/C^C?)ee/Td-8Q5JXU6/dQ\?V+<^YUdL@5;M^Vf(8(9Db+N]V/[67U?
gcWE\+6SUWB>FE?44S7AAM\=[6KM@.M^d:30,Y/@d=dG@)C1;B4^UDgXN_9[,IYJ
gK_AF50U\N()?N,+LCZf4\UL?2+SH=S>(cVL9.>8Y+E-,LO;C;V;W3a\09-Z?f>#
+#&]0V<=.#.E)5ENUf&9UA.U.T)e(Mb;UH26@Ba_SUf5Accf+gKgY/781&-1KC7d
)LL-eRXfb<O^=6#9_\XS,DD_UE<=O4J8/EM(0D@7M\C#U)f<&KUf+O?+>;M[#BVC
KCXI1;W4Y0^cFCTR7W4DYVKMc]7](K<8Q4=&VOZUDOUd4cTAA^Z__&(;W/^:GT1S
1Z9_IVDVH:=f#K[/1?Cdg1\C=0UVf4><Ef#(V:4NS/H[<U(Q+(SSa#/R+R7O^dRe
EI4CT^+M#?O0dGC&bX?#01b^X8F/CX&[8\bHY;IU)PgG8M7^?KVCd1MPID?^F[Y4
JdSR37cYIR[g+;:-cV4;3a):)#DPcQRE\H^Gcf8K9JU6YAgC2FCfI=ZY.@ba9H)N
W@#0<OS2+TZLJNOfDS)DXO4CfS<@1>>J\cA^92XaU@KJ6[ZSC43ac^<<#-FaCHS,
Z3^55AD#V,+534c#(/B?7:+L1D1K<<\TOU<dC6/?)9bF)VC<<W5IF>[JFYa/ECTK
Y6M\b?@=[PXZV#cTBLJ=^Oe<RJTg=^e2d_HGYE[>T2Q<cH<a]?,OH=J859f&3dDA
^eH#_7+GMG49V#(78>Wd:6D9Tg5Q-GJUVK.MB7\e^K6?0.6CY;&#B)Y&c#O2Z7]A
PAC;\3#OE<G5gYZS^Q38e7TQF+D-UI7MMQ-\_<dZ[6\E#/agX6e[\cG3F6HE/F1:
L9BHKNHEJ1B\KcD60AX:f5MERZfgUJ<(78F(1W&P_KdHb5O.9>5TaG=F^<GeOgR)
dJSF>TLURd&V@8f1OPdRZCf[]=L2PV5(,9g?,&f8-O+XRIV6NZ<L.Y]7+:9bVaD+
^WD?K=FO8VaL?Rg#cbDD(S+&?OSd.g&V1A1@aaE#f<FEB&Dfd?\DJ;NNVM@9F=]<
9a([&)E/f(aP3H7_RQ\4Dd>==NP5>JXe,TXHae.&)5e.X:Y2&R=WPO?>=CFXLPJ9
JbZ@U=TF7f;F+K+WF0><IHF1J?;4_?S4AKd\/GZUcSELgYO(b>=F5[@]2#MbXgPS
:=8XTOND<6-0+8cCCQ/DHOS<_H<Q#_f)Oe1d._>[#=.O(/)F4(6>8(aRVL[CLd/8
FX#gSV#A0IU9_[5BK7RCBK+b36aVYeRO>Q[c6cTSfS3^#CC=5[5.IdZI]C5R/b].
:RAHgaN@O:YLMC\G(FWd?;\]@-0@9gDC]5B_6=;5aSMeZI9ZW<A\9bJV.EAd)TfG
+;7:A(A^C@>^NM,;A(:43(gK^@1AGSA8EAMCGO0<,BcHRdYAMJ<06SO,/d5X0\H9
AV8E7[/bE7.B)X5^?N1SUAcE8X&a7DXc]<?A8=aIfgaV_95/22P]LA0JPUYFGN:_
ab+FYI58@32AI7N:XW5eBgC01Y-C:X^AY=X.3AIa4J&cH\JUL6=&0QOOb(UZD9JC
03dT-;>WBJ.bU:8-];]aLcNYA\D1]Ye08L66#D4bAMG+V#=-\+,WI0TW:b#.ETRE
d;2JcbZ/=,dJaF#@Z[P^/+O1A8(0W[7>8?:EdKABJ(/?3^L&1b?<[P-Z^A3;BQDI
]A-/:6:F>06.>\aGP]::PDYf9.Y+Da94VU[C]a6#3#]HcR>_8[;WcM63R6;J=;9X
NI4VXD13;?AVQ9_=7](aI/XA;2/NJ^WNDL?:3S&G3OIAGSG5]@1ZH__a\UGWaWI\
QG8PL+]-1(HZ.f4:YW:J:[9\8/DG0+L^YfA<TZ9Y=J>P,0)W4=+Z-(-a(KX:_1+1
#9G8#H;-YH(6N(bWfRF2SN4J&@[a]VbA:FH:RK-B<5(]K+LO&2O#U[]?,E#a38U[
8N+C9Q+^U3JV\2ZG3\?04b?C9K13,;<IV;9O^Cb(Ba1d,&\8^?_LgLV/f.N9IGR&
J7_Q:BL;3PV7,[L?UO[>0f#W&f56I70<C1g4,L4cKF95D,(+TYfL1FD)eZ(:J=>=
UYa=L5>)Ig@b=;8gc&/>&U.[2+XR1B=3fB??Hgg<\f.S;We+K?\@EA:Hc:W/f3&B
9^\#-Pd=03N.4NM?g@WBPH9&T84d;IRH(/TB&B_8M7LD><Pc_?<(gK3Qc3(O3Z,W
[I#,W(JEO;KVaF0B(_0OK^@>KPD81eeQ)99UEHM2P\5-KREIUR=C^Q-6>POf_JRP
CAQLN_a\H#\ZW4RUKf09OIOO3V#FMMV&G<0NBRXP0-(Xg?CP;/TDC_1^SN.=.0)V
d]MJ]3>G3?6&<FCcFL./R0?+ZQ^IX&C(Z6#E+6=AKP?0.g[g==<MPg)&c.W@M27[
]VJS+S?9d4abZNJP+[J2HSA4M4KO\;;A,]fEGONQ(,]Z74MJf6S/JQ>4(TVWVNR#
0>;QJ#&8[Ke_ZRU<OcFbUT9VE72A@fXO8:Y8&(^)7/#&=GG90.NWZBcQIe(+)7L,
G_T=NX/Ia9M7-L]S;P>/c,BJRc^5Y4)D9=X7ISf,eA.74M@Z0KP-R,.O/K-?TX>F
NYPMW_1IR^(gNO7Y>5e0aP?P.g6.5S]YL7_TWLa.4YR\UI8?>[^ZH(T#\#Vc(F#&
=9Y#dQ-W3/]aU5+:=Q\945+@&M4F^(_VDde;6<#:Raed]?73:@b]@V/?OY,QUBb@
XX,+5[-Sa&/5<R_7NJ5J(IdWI[+_A5^A)4L1&.S(J\/Bab<4M[M[Id(dGe_cg/bH
7F3[E:X:;E=NRD<8#WZ?8cC]g3Q,^5Z@U9XSS__>VM/#bI#E2SbC0G7dg2I3HH<Z
LN;ABLf6/6.5&P2>3V+,ILDRU9&&K.b5>,A#4VNa/N[WA,:\Q-::A7BNZ2If,^)V
ASQ+R54&FGI=H,#?R&A+L+/ccWfBK&8WRTPWY^/f[&-NDL7a=,(3O=^&_7c,#R@_
[WOc-E>f)8d2DPHGcE^gda3;HA#?FNW[U.UQ_4R9\5Xd>)G..6L5#Ad#2TZ,)1,K
]:bM9e8R3=6/\PQ_\0@OT]&QO4/FX4bA@\13PfNL.#3D0f9GQ)T&cE<ZDT14BZZM
\\D>3A2F4U&3ZKfaFD:C<BgGD>e]\a(dG2Q+9RJW9U]aPYD_E,AW;AKJMd7V/N1K
/:PXCHLA>?274OeTPJ-9M0X-56&1Hd6.Jg@.8-bK[J>5TC]9M]&IOKW3-9O53a-+
e\/T[O5.C.H0X4:,]2D0<D03:OBY-R+\JYZ#C-6@CLQMIHCLTHYQP/I?+GW^EFDN
ReD=4@P+HYD1G,Qd/QNefHIgD6O];R],\V\8F3.X&ME)X,.0,aN+:52[.TE#cL((
?=@VXc7J5.-OdXCZA;>?^1F/dX7Da-B29PdCL&M2[Ac3ZfQ()=016YCb3W^LaM60
3<9)S)(&J?XcL?W6IR?0Y(TUQG.)-A(.N>W3]+XR/-:,FR4SeKRO5&S9;[cZbf@d
9TdDO.[-V&QY<735FfC@80YG7GUWP#H:/)OJ<ccBV@G10LAN:1\6B7>Z9BXJgVIW
.E\Yf_,&FJf>b\^2efg(OaY<J^CUU03g64=>D8.T1=Od5P6;#:bY-RBK<(fC],?1
KLG7AZ^S#+]75UH_=F.fLJ.OD&ZJ][2K(.+NZJde\95B-^((NM^6E@UC84FC7+Db
dPNTR3R7eABgKEA]X_&9SI06OAOfH0[D32c6HcZ(N4G:]9,=;ga&.6,bbdLJf63G
W/W&S1SaZ,+M>BR#e@eA]\MBS:=A(Xg.]\J[2RG0U4_+KS7GUG9^-WT_<=@5EfeX
F0U06XV<#GZLQM#-J1>/\F=b;]V+N]@[Fa.@c>A,YU[Q#_Ba]bJP,QK^&QC5+CNK
;gIM8=Yd/da6eWMG8K<<[?AO\0Xb[=>BH_N@bV8\-SdZ,3?fK)BDI?EYX64DK4I\
_^K0R#AF3T-aMM[AQXZ_S^b#88MFYdb/b#f/5>-OP4+KRSY1CW82HO;+2+<d]<E+
Ig#KLaZ)[_1XWe:H<fcM]#gTD9>L9-F3X-4>58b9B)I=NG+@_c2EBg8GE,0X3Ue5
0JY9:_^V?3<@X8XZ@(U9&/OQ9CD&NW7HSaU7JV<H@,@ebfN<F:9P;>c6QSfMRa&8
XJfQ?BgfO27ZX6<IF].gAU9eBg.U23;df;<De-11JfC@Gc?]=>JG7?N([R=7CX(e
WBWW7CBe]S#6bB-146@R#Z0b6<deb1],01S1?WF=1c],@&Q=BeVb]b>bP445N\AC
Y<85&)0LaOA]?+gB?^0,3JgGW-3.R_eL^eC@b38_SS7I-+A\PWd3=3XOAA>TS<Yc
\:OU/38_f98LD-G2.1,G8?DB.AU5J)J_G[GK8OP=B:?UR>MA-GU5dT^#MCKZ5b[\
H<R5,IAZ=a:_KPfUb5_8AdJ4([:S#NZ5b:^I\JIaP=aE)IaL_TMAM^J&FJ:E=MDH
LbUbRLWJKT@)@E5O2F6P2ZJ>[Z8Uc6OWEX@fUJ5/>UZ\?bBA\C6^0Ee87O?ENYBC
;3J,-gTD[[&<ZSdCJK+c-Q\Ve+,D&/1E@5?,4YSN(:^AICR-1D+=2SU/N&bK\([F
SSR^44&&bZ1E&CATQT6Z?Te@(TP>VEZ&S_)U2-NDcF^4W>GHA0F/>MQMffG?;J6J
?=:<PM0=)OMS7TAc&Z+(CU)V#3eHd,CGX<G6a(I\V#LR<XV5_-<2#>;,fGg-43Lf
P@FLLb_#6;8O5HVAgV_dA]R05.71R8FH\)^WQZS,@\X4(&V2[RQb29cJ4#fU2bfU
T(_BA1UO(Qg0+,F,.DJfTFZL@36CAB3O>;H_RJ5d5GL&MNV.>ET2=K7R31@d+(0c
7\V@E:]33EQR9J;D;(.XQ3[WaG,3&,43A_Wf.0DQee#9WDA(0YIS,-Z@6S@>]]K]
U\DU=F6UcI:\,):RHC2JfDBM/J3/>U@XY<V1<WV](O.>O?B8>Q(H949EF_.G:cEC
P)4UY10C78&4CLcVG8@9C].QUX]Q84,9]>gb6Q/DGF_La&=R,&C:d?8+Ke[_SPP0
.a<F1a(_I\3T[O.G+<a2(F2f.6=I#XL5J/Vf:Ig=[84c#NH]g5JQ8bKI/NgD-<0S
H#IPURJ00R&B^Jc^_)#+=4#SYF2TCf&/W&<L>2?e44JAP\.[dPJNeHE#PG\U59>:
c[><@V&PC::.@1YgB&g89f,fdT&@KMHd3RRQeRYZ&LA=d88eXL=C/Ng.&9X+d]Wc
\+S\dJT.VM5>5OXf]UH81@?OBTB:)?HPG0^D=J<6S@21H8_V#LJObcOeZU;,5(#^
[,=V<=AP]C4),DDa(ec5^RV(ZR+2C=K(gYP5\^5-9W92O2@=.@W2S(NV[;C?7fdJ
8DPP\LF;dRC9?=8L4#MNJ8]-4>+UZV_<bD+\b9[8P^U5Z+R/-gPdbC>&IQB;8:DU
6W(C<ABgTG2Z]2MJ:.5_Re#\A(84BKO+OPBZ^a.b.]M\YI7)I0:UW+R4Q@IG=.#+
_Y>SA7JLcB^aS4TZ)@1NUJNOU]#SgK38,)>\1B+AU0T?BG^##1dc3QAa::>Da-g#
BKZe2SVKCZ3Z29-eE?(?/63+)FOUCY/e;b=\RK]<TAc(=7LMdcQ@P2W.((R=ZY5;
-GNI#AfcCE4;:AYLAb2Ydc;2=Yg5<;RbT_daf0Kd3:21[O49aTRG?]=PC7QA)IKO
dX\6^^d?2d6/X9&-+ef4VEMQO@@?;EY:(^37V5.B&bQ@IPe5X#bGXFZBKe.^67[M
J0(ZZ#N6=8EE5?VWEMg5Z0DPc[ON.3?J93DR>aQ-\a.F4U^RcB:WTc:\-RGBH8.<
\_WRW\P4^,cP3\&e=.W_)C05GV1_;PFZRe;6bd)cBO:G37C[IC\?]E,8OPPYU&&H
5((2]Zd3FdRN5A3/7EB<Q+eY-Z2JE)aS_B1\?SK/S^J#5&TaLf1_S5LOf>,@W#I[
?\J^3DgCV^d08T6+MY8#-Y5gM_Je90d_@\Zf;RIL5e\^_,+\b;5J2L^8TQ1DWTfG
V.,fB^UBY4@QP+FF_MPa#R<^E9\R>UU-,,[<c\B6+NZX5dN/LcRZ0@;db?YfO;c/
?[F&/)CBJ<T_?fVXCSC]+g2/TUNUCbb9OWBc=H/Q@f18GU;cc1D:7C-eJ9eOaI=T
_)NVO@a>eW?9d^(;17.1#/=,d>#a@)H/E#<B934X5=8W@Q,)HSf97MB,^Wb7+WY8
.O1W.F>(a5;89IR719_1C]be\[()PL#QcN4GEgNY[NN=CCQ_ZR1b9VO^3U<Ya&[M
NI88[.UX,U=GD1(H9Q-:c^JceKKfBDc/IX,2Wd;WK&M?0#8SJ&#[;01M77g&/P]_
M>ILAHQAEdO]O1AY(7?cYNDBK<UOQ:KWJSVe1)ZGb@O7H>Q6;ab.7&)_K;egY6L>
G?)L:>f/1#WTaMRGGG.fU2+[Z95I,OWKdG=P;D]9Ibb8<<FYKKK])-H.Q[45U]9e
>6>JND1F&gZ/)7UKF\]1A3O0LI3CQ/afONac57+)]KBHV\9THXeW.fU7^9R0F;<Z
Y7Lc7;[P0NY_GS8agY[eYV,3b0+_]EEc/6[]^Q9Yc<UUWUcc4NZ?-gN2bZU/X6(,
GZ7\@RL4B:8gS3WDGe.\=G48CA=1d-<YK.[6b6[EbMa80I]ZF=D<J;EdCI6J3[?5
@ICESFUa]^,SUR0ZeJ#@IIMD,2-;G]PKX.NOfg6CTS_I\&<?I\8SX;>+e#-+-+(&
+f./]Q>U^;4CGSC@[&XbHg)4:[>6MZ?YgVNbWBQKcVW9eW>H@_a]A_g\fd\.(]:M
EO;;Rc#GAd?_/Wg3W#8WME\3d-(@F72#Ee3/=R><3QY+/.?I^f/DS\O7<Tg&/X_R
HbEE^VBW=b>=<(FPTMI5EN0UJFA>^<9QG]e)IT]<bKP9QM:Y0Se+b[2)8-gWJ\G=
1=-@2dfAHXJIaX9[H-80+J-dK0H<Y3^72EcJ:UKG+/E0[GK<0EYTFUV/\C=2X37[
\NgIe3W;UdC?)BWP?#1eJ\fC@?F=)Vc?6#RW847HY4CZ=e=)bb6Jf&CKO3H<6M-f
6GN_:bQf2UF:.NPX+B,C&D09X7a4_X8R(,f;F#KH>B9P2f/XD.OV4^GXBU?aCBG8
&T6U8+)3=,._4#be-_G(KCUY\JX=2;@YYNL;_O=GTaG:c>e^-&HC/A?U6><WYfFb
1\3O0<I]Y2I;a)D#WE7.[2M6Z4/ae+].aA2cZDN31AT08GS=/JWM9ScL,I@0#:ab
\RegK<fEbeQNP0e\,0f>+a7?&R/&b7>0dI90<Q]\d3Pb(<d?E09XWc1/(,I_-.^.
Q1/1Dd/O=1^[6fa&ZM)8,9JQYICKHWX)P?V1ESWJZ[KSL[adRfaNB/UURA]\K=I&
PKJBP.J-ZFH245.?RSWMX6I8_JEPbD9)>>A(6R1=J53#>HK\#4d1GQ08f3IVJaJF
g1Y19:>cE]:ad_@/IE]0Gc8G?HF5L/7G[dQ8QRY9XUDJ5Eec;KHRe5:^F^McQK]D
;bE?eBC._J0a5#>d]Vc5W^)Z-6RL1GW.PO/5b2+E+)NPF#QW;FOI6&WE<(DQ&18E
P4gDO5@E#1KQ)e-_NP_DI#7@OF#<]WeP<\-#FTL/3R_N\0TX7HP9YCK:YH9aU<d;
@+Ib+DGDTM4^)Z]fN87^8M(6<)]3XH?e#[L:BEATQ?WZG^_=gT@TDX[MW=6:YER;
FXUA=X96P;YZ^U^e;E3E>/<SM&.,Q@I[2-0[TQE<\4M,ER,J8;>DdI@B.,=:\<S/
fa44E:?OLO#]De#XRG@e+HedFU.?Bd0.gYG(_9<QV>@f?fg(K==FIC[gOPS1c1FJ
Ke0MEHeX9Z(4Z),HU_YA;fUGG.dIe3G=e?e#QA_P?3e6QVV>_G9<8_85^RD7Da7_
LMJTQM,I[Y:(FMHOGSY[(QT]B)[J#01_O>e;e[F)YO:9]2XgSP@4W3<CGPEKD;Q/
G2]#KU;37>7T&Q6E499X?M#d/g/MN[:J^76E6^&U(Q-WV;5YVTG6g,.@P@Z^Ed0+
HFQ0HT;YNMZa&O71SbW?T0QD1Y<(@Z77ADB_<UaG;&W:=TORAL2B@O5(gL?+fSC(
R@c<^,_#ECL0Xf@^T@3dNcZGB5@F87#U>eVL\dM9;bO;_H?N2&>ZD1.EWDFS(KYZ
97QNZ(WZN#Le.6d_896W4#QAZ^4OFJd#W)QE/0&fe98LZ)DPQgE;>),V?fFbK)T:
LgJ>681_^&\\[ZD-C?N61XOOU;.F]HEHKG.a2G3W8O=9[AY/>&gU>3g@ge+8.C9O
5FN#V#.U5.9e8K)-V6/IdYbA:B4fL@Jf.fXN9KAcf,5DVISW]Z@,H__5;Q-RaA(7
G3)NC@^fH\2/2P_=b,WZa50T^aFM2L@0Z]MXY[Sbd0RV_[R4_416&Y0PA54UK.R4
,-bS@88&KeWdU1[P,@GXaCHbA?#A\9-fOb53;IW3H^M^75V/O),e5D.0I<H[;A?T
LXWJE^>D<CE6;TG&^E<;)]G)E(_8ReR1Y]b<,CIPC7T45K=3K&MYEKI#0f[ZV<KN
:WITd[9fXN5.EA/+=+J,?)_Mc.fUY6=>bScCS@eE,eB30B)?dY&Z;F1+_:E@<DCf
Fg\)D<-49L.J>FJ?Z?1?/<YIHKX<5VX-K/O.GS/.)I..R^9>1eCHf0dd5OB<-Y>:
X2OJGELZb+3fWP#DHbU8(_,BbDGI9(E[S8I85TMeTGXaOUK8WCIX2PN)1.TCHOc?
^F\O(<D0eR.7\#c/)8WL:[T-Ve;_Yg1Hd9g/Q;MVXWaZEW0H@HVM^+,?bd#L@<&Z
)L]@(^Q2R\[+]F:A8XJg,^I&8+03MI8R)VND+=?[.34^9I>-=T]e\Z>_)T@VKSP2
E1AYJN2TLeDW;AWKJVZJD^EDFY#4,&DDJ8:0M?Fb\2-A:JAYA29CSFLOCYDCB_RI
O[:/))0=>9_:0GX1<a@_S>W#1J>J:+Ee&KU78RG>#,VE+acA,&3gaC9T-dPWZI.2
cC.g-EO<7?R4;L3I[LQQeE=MJg&TARXD,dQ8LKaVP5BE2[-IVQB[\Ng;\74^dB\F
a&OX2Q9G\-P)PR:=OQ6]?#D[:c:KfAR:a?#_+a:(+];Y+R.O?[P<^K2B:[8P5_L7
XFc4Og/3<:Dd8G;:9^[J;IdJHT7;A66#,ag89K-S8&7R>TK/FUXd0BR)RcO4RWb;
B+3R,R86?bXCQ05dT8C0CGZ0VUV6ELK04bS+FS6gT\cMO8Y@/:66Z4<^^FZ]@aa5
F2Z8/G[UeTN;e^F-)I5KT/5;?D[KVRR)6a6IKcCKAA^WVN+09Y#84),XJ27\U9;b
#@b&bbC?^KSPN1,M_7e7HLY.ge^5,E:<=1[dccGaK5T66eLO5Yf6Z=W.;SbU#.+9
<>O(5TL[MC8EBUfb#0-?I&@K]e:V-7T83;A@bB^DZPA)6>cJ]U3I10T^\M:@]gA-
JG\_<DXH.>ARGaa>UE#X;W15@-(f66@dMaACTX#_JTBSc6)RR+\KSf;1HPV)ePT@
)KNMV6:Q,+M+Jf6R;X1<;g155$
`endprotected


`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
  extern function new (string name = "svt_axi_system_configuration", AXI_IF axi_if=null);
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
  extern function new (string name = "svt_axi_system_configuration", AXI_IF axi_if=null);
`else
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param log Instance name of the log. 
    */
   `svt_vmm_data_new(svt_axi_system_configuration)
      extern function new (vmm_log log = null, AXI_IF axi_if =null);
`endif

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following
   * 1) calculate the log_2 of \`SVT_AXI_MAX_NUM_MASTERS
   */
  extern function void pre_randomize ();
  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************
  `svt_data_member_begin(svt_axi_system_configuration)
      `svt_field_array_object(master_cfg              ,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(lp_master_cfg              ,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(slave_cfg               ,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_object      (ic_cfg                  ,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `ifdef CCI400_CHECKS_ENABLED
    `svt_field_object      (cci400_cfg              ,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `endif
    `svt_field_array_object(slave_addr_ranges       ,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(system_domain_items     ,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(ext_dest_addr_mappers     ,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_int(enable_xml_gen, `SVT_ALL_ON|`SVT_BIN|`SVT_NOCOPY)
    `svt_field_enum(svt_xml_writer::format_type_enum, pa_format_type, `SVT_ALL_ON|`SVT_NOCOPY)
    `svt_data_member_end(svt_axi_system_configuration)

  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();

  /** Ensures that if id_width is 0, it is consistent across all ports */
  extern function void post_randomize();
  /**
   * Assigns a system interface to this configuration.
   *
   * @param axi_if Interface for the AXI system
   */
  extern function void set_if(AXI_IF axi_if);
  //----------------------------------------------------------------------------
  /**
    * Allocates the master, low power master and slave configurations before a user sets the
    * parameters.  This function is to be called if (and before) the user sets
    * the configuration parameters by setting each parameter individually and
    * not by randomizing the system configuration. 
    */
  extern function void create_sub_cfgs(int num_masters = 1, int num_slaves = 1, int num_ic_master_ports = 0, int num_ic_slave_ports = 0, int num_lp_masters=0);
  //----------------------------------------------------------------------------

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(uvm_object rhs);

`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the OVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(ovm_object rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);

  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static 
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);

  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif
  //----------------------------------------------------------------------------
  /** Used to turn static config param randomization on/off as a block. */
  extern virtual function int static_rand_mode ( bit on_off ); 
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /**
    * Method to turn reasonable constraints on/off as a block.
    */
  extern virtual function int reasonable_constraint_mode ( bit on_off );

  /** Does a basic validation of this configuration object. */
  extern virtual function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);
  // ---------------------------------------------------------------------------

  /** @cond PRIVATE */
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);

  /**
   * Simple utility used to convert string property value representation into its
   * equivalent 'bit [1023:0]' property value representation. Extended to support
   * encoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit encode_prop_val(string prop_name, string prop_val_string, ref bit [1023:0] prop_val,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);

  /**
   * Simple utility used to convert 'bit [1023:0]' property value representation
   * into its equivalent string property value representation. Extended to support
   * decoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit decode_prop_val(string prop_name, bit [1023:0] prop_val, ref string prop_val_string,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);

  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern do_allocate_pattern();

extern virtual function void calculate_port_interleaving_parameter(output int num_ports_per_interleaving_group[int],output int lowest_position_of_addr_bits[*],output int number_of_addr_bits_for_port_interleaving[*],output int lowest_port_id_per_interleaving_group[*]);

  extern virtual function bit is_address_in_range_for_port_interleaving(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,svt_axi_port_configuration port_cfg,bit is_device_type_xact,bit is_dvm_xact,bit is_snoop_xact,output bit is_device_dvm_ok_for_interleaving);

  extern function void add_to_inner_domain(int ports[$]);

  extern function void add_to_outer_domain(int ports[$]);

  extern function void get_masters_in_inner_domain(int port_id, output int inner_domain_masters[$]);

  extern function void get_masters_in_outer_domain(int port_id, output int outer_domain_masters[$]);

  extern function void get_masters_in_system_domain(int port_id, output int system_domain_masters[$], input bit used_by_interconnect=1);  

  /** Gets the slave port corresponding to the address provided 
    * Note that, "addr" provided through argument should be untagged address i.e. address which doesn't
    *      have any address tag attributes appended at MSB.
    */
  extern function void get_slave_route_port(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0]
          addr, output int slave_port_id, output int range_matched, output bit is_register_addr_space, input bit ignore_unampped_addr = 0, input int master_port_id=-1, input bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attribute=0);

  /** Allows user to redefine the master to slave routing behaviour in the interconnect VIP. Interconnect VIP will call this method and use the first slave port returned by this function to route the incoming master transaction.
      By default, this method is undefined and returns FALSE.
      User is expected to define this method with the routing behaviour of their choice and must return TRUE. Interconnect VIP will then use the first slave port returned by this function for routing master transaction. Otherwise, it will use its default mode of routing master transactions to slave ports based on the address ranges.
      Note: This method is applicable for Interconnect VIP and System Monitor component.
      */
  extern virtual function bit get_interconnect_slave_route_port(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] tagged_master_addr, bit is_register_addr_space, int master_port_id, output int slave_port_ids[$]);

  /** Gets the slave response corresponding to the address and the configured region & its attributes 
    * Note that, "addr" provided through argument should be untagged address i.e. address which doesn't
    *      have any address tag attributes appended at MSB.
    */
  extern function void get_range_region_response(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, bit is_write, bit [`SVT_AXI_REGION_WIDTH-1:0]   region_id, output bit[1:0] slave_response, input bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attribute=0); 
  
  /** 
    * If the domain_type is outershareable, checks that all masters in the inner domain of the masters
    * listed in master_ports[] are included in outershareable (ie, in master_ports[])
    * For all other domain types, no check is done.
    */
  extern function bit check_domain_inclusion(svt_axi_system_domain_item::system_domain_type_enum domain_type,int master_ports[]);
  
  /**
    * Gets the domain item corresponding to master_port and domain_type
    */
  extern function svt_axi_system_domain_item get_domain_item_for_port(svt_axi_system_domain_item::system_domain_type_enum domain_type,int master_port);
  /** @endcond */

  /**
    * @groupname interconnect_config
    * Creates a new domain consisting of the masters given in master_ports.
    * @param domain_idx A unique integer id for this domain.
    * @param domain_type Indicates whether this domain is innershareable/outershareable/nonshareable
    * @param master_ports[] An array indicating the ports that are part of this domain
    * If port interleaving feature is going to be used in testbench then this
    * API should be called after setting the port configuration "port_interleaving_enable"
    */
  extern function bit create_new_domain(int domain_idx, svt_axi_system_domain_item::system_domain_type_enum domain_type, int master_ports[]);

  /**
    * @groupname interconnect_config
    * Sets an address range for the domain with the given domain_idx.
    * The domain should already have been created for this domain_idx using create_new_domain.
    * @param domain_idx The domain_idx corresponding to which this address range needs to be set. 
    * @param start_addr The start address of the address range to be set for this domain.
    * @param end_addr The end address of the address range to be set for this domain.
    */
  extern function void set_addr_for_domain(int domain_idx, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr);

  // ---------------------------------------------------------------------------
  /**
   * @groupname axi_addr_map
   * Gets the local slave address from a provided global address
   * 
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to translate a global address into a slave
   * address.
   * 
   * If complex memory maps are not enabled, then this method utlizes the
   * get_slave_route_port() method to obtain the slave port ids associated with
   * address the supplied global address, and the supplied global address is returned
   * as the slave address.
   * 
   * @param global_addr The value of the global address
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *     mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *       indicates a non-secure access
   *     mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates
   *       a write access.
   * @param requester_name If called to determine the destination of a transaction from
   *   a master, this field indicates the name of the master component issuing the
   *   transaction. This can potentially be used if the routing has a dependency on the
   *   master that initiates a transaction.
   * @param ignore_unmapped_addr An input indicating that unmapped addresses should not
   *   be flagged as an error
   * @param is_register_addr_space If this address targets the register address space of
   *   a component, this field must be set
   * @param slave_port_ids The slave port to which the given global address is destined
   *   to. In some cases, there can be multiple such slaves. If so, all such slaves must
   *   be present in the queue.
   * @param slave_addr Output address at the slave
   * @output Returns 1 if there is a slave to which the given global address could be
   *   mapped to, else returns 0.
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual function bit get_dest_slave_addr_from_global_addr(
    input  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] global_addr, 
    input  bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input  string requester_name = "", 
    input  bit ignore_unmapped_addr = 0,
    output bit is_register_addr_space,
    output int slave_port_ids[$],
    output bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr,
    input svt_axi_transaction xact);
  // ---------------------------------------------------------------------------
  /**
   * @groupname axi_addr_map
   * Gets the local slave address from a provided global address
   * 
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to translate a global address into a slave
   * address.
   * 
   * If complex memory maps are not enabled, then this method utlizes to obtain the slave port
   * ids names associated with address the supplied global address, and the supplied global 
   * address is returned as the slave address.
   * 
   * @param global_addr The value of the global address
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *     mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *       indicates a non-secure access
   *     mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates
   *       a write access.
   * @param requester_name If called to determine the destination of a transaction from
   *   a master, this field indicates the name of the master component issuing the
   *   transaction. This can potentially be used if the routing has a dependency on the
   *   master that initiates a transaction.
   * @param ignore_unmapped_addr An input indicating that unmapped addresses should not
   *   be flagged as an error
   * @param slave_port_ids The slave port to which the given global address is destined
   *   to. In some cases, there can be multiple such slaves. If so, all such slaves must
   *   be present in the queue.
   * @output Returns 1 if there is a slave to which the given global address could be
   *   mapped to, else returns 0.
   * @output slave_names in the queues
   * @param xact A reference to the data descriptor object of interest.
   */
   extern virtual function bit get_dest_slave_addr_name_from_global_addr(
    input  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] global_addr, 
    input  bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input  string requester_name = "", 
    input  bit ignore_unmapped_addr = 0,
    output int slave_port_ids[$],
    output svt_amba_addr_mapper::path_cov_dest_names_enum slave_names[$],
    input svt_axi_transaction xact);

 // ---------------------------------------------------------------------------
  /**
   * Gets the configured slave address mapper from a provided global address
   * 
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to translate a global address into a slave
   * address.
   * 
   * If complex memory maps are not enabled, then this method utlizes to obtain the slave port
   * ids names associated with address the supplied global address, and the supplied global 
   * address is returned as the slave address.
   * 
   * @param global_addr The value of the global address
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *     mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *       indicates a non-secure access
   *     mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates
   *       a write access.
   * @param requester_name If called to determine the destination of a transaction from
   *   a master, this field indicates the name of the master component issuing the
   *   transaction. This can potentially be used if the routing has a dependency on the
   *   master that initiates a transaction.
   * @param ignore_unmapped_addr An input indicating that unmapped addresses should not
   *   be flagged as an error
   * @param slave_port_ids The slave port to which the given global address is destined
   *   to. In some cases, there can be multiple such slaves. If so, all such slaves must
   *   be present in the queue.
   * @output Returns 1 if there is a slave to which the given global address could be
   *   mapped to, else returns 0.
   * @output slave_names in the queues
   */
   extern virtual function bit get_dest_slave_addr_mapper_from_global_addr(
    input  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] global_addr, 
    input  bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input  string requester_name = "", 
    input  bit ignore_unmapped_addr = 0,
    output int slave_port_ids[$],
    output svt_amba_addr_mapper slave_mappers[$]);

  // ---------------------------------------------------------------------------
  /**
   * @groupname axi_addr_map
   * Gets the global address associated with the supplied master address
   *
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to translate a master address into a global
   * address.
   * 
   * This method is not utilized if complex memory maps are not enabled.
   *
   * @param master_idx The index of the master that is requesting this function.
   * @param master_addr The value of the local address at a master whose global address
   *   needs to be retrieved.
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *   mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *     indicates a non-secure access
   *   mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates a
   *     write access.
   * @param requester_name If called to determine the destination of a transaction from a
   *   master, this field indicates the name of the master component issuing the
   *   transaction.
   * @param ignore_unmapped_addr An input indicating that unmapped addresses should not
   *   be flagged as an error
   * @param is_register_addr_space If this address targets the register address space of
   *   a component, this field must be set
   * @param global_addr The global address corresponding to the local address at the
   *   given master
   * @output Returns 1 if there is a global address mapping for the given master's local
   *   address, else returns 0
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual function bit get_dest_global_addr_from_master_addr(
    input  int master_idx,
    input  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] master_addr,
    input  bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input  string requester_name = "", 
    input  bit ignore_unmapped_addr = 0,
    output bit is_register_addr_space,
    output bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] global_addr,
    input svt_axi_transaction xact);

  // ---------------------------------------------------------------------------
  /**
   * Gets the local external slave address from a provided global address
   * 
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to translate a global address into a slave
   * address.
   * 
   * If complex memory maps are not enabled, then this method utlizes to obtain the slave port
   * ids names associated with address the supplied global address, and the supplied global 
   * address is returned as the slave address.
   * 
   * @param global_addr The value of the global address
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *     mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *       indicates a non-secure access
   *     mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates
   *       a write access.
   * @param requester_name If called to determine the destination of a transaction from
   *   a master, this field indicates the name of the master component issuing the
   *   transaction. This can potentially be used if the routing has a dependency on the
   *   master that initiates a transaction.
   * @param ignore_unmapped_addr An input indicating that unmapped addresses should not
   *   be flagged as an error
   * @param is_register_addr_space If this address targets the register address space of
   *   a component, this field must be set
   * @param slave_port_ids The slave port to which the given global address is destined
   *   to. In some cases, there can be multiple such slaves. If so, all such slaves must
   *   be present in the queue.
   * @param slave_addr Output address at the slave
   * @output Returns 1 if there is a slave to which the given global address could be
   *   mapped to, else returns 0.
   * @param xact A reference to the data descriptor object of interest.
   */ 
    extern virtual function bit get_ext_dest_slave_addr_from_global_addr(
    input  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] global_addr, 
    input  bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input  string requester_name = "", 
    input  bit ignore_unmapped_addr = 0,
    output bit is_register_addr_space,
    output int slave_port_ids[$],
    output svt_amba_addr_mapper::path_cov_dest_names_enum slave_names[$],
    output bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr,
    input svt_axi_transaction xact);
  // ---------------------------------------------------------------------------
  /**
   * @groupname axi_addr_map
   * Returns whether the supplied slave address is legal for the slave component
   * 
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to indicate whether the address received by
   * the slave is legal.
   * 
   * The default behavior of this method is to return 1.
   * 
   * @param slave_idx The index of the slave that is requesting this function
   * @param slave_addr The value of the local address at the slave
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *   mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *     indicates a non-secure access
   *   mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates a
   *     write access.
   * @param target_name Name of the slave component that received this address
   * @output Returns 1 if the address is legal for the indicated slave, else returns 0
   */
  extern virtual function bit is_valid_addr_at_slave(
    input int slave_idx,
    input bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr,
    input bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input string target_name = "");

  // ---------------------------------------------------------------------------
  /**
   * @groupname axi_addr_map
   * Returns a valid address range for the given slave index.
   * 
   * If complex memory maps have been enabled through the use of the
   * #enable_complex_memory_map property, then this method must be overridden
   * by an extended class.
   * 
   * If complex memory maps have not been enabled, then this method randomly selects
   * an index from the #slave_addr_ranges array that is associated with the supplied
   * slave index and returns the address range associated with that element.
   * 
   * @param master_port_id The index of the master for which an address range is required
   * @param slave_port_id The index of the slave for which an address range is required
   * @param lo_addr The lower boundary of the returned address range
   * @param hi_addr The higher boundary of the returned address range
   * @output Returns 1, if a valid range could be found for the given slave index,
   *   else returns 0
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual function bit get_slave_addr_range(
    input  int master_port_id,
    input  int slave_port_id,
    output bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] lo_addr,
    output bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] hi_addr,
    input svt_axi_transaction xact);

  /** 
    * @groupname axi_addr_map
    * Virtual function that is used by the interconnect VIP and system monitor
    * to get a translated address. The default implementation of this function
    * is empty; no translation is performed unless the user implements this
    * function in a derived class. 
    *
    * Interconnect VIP: If the interconnect VIP needs to map an address received
    * from a master to a different address to the slave, the address translation
    * function should be provided by the user in this function. By default, the
    * interconnect VIP does not perform address translation.  
    *
    * System Monitor: The system monitor uses this function to get the
    * translated address while performing system level checks to a given
    * address. 
    *
    * Note that the system address map as defined in the #slave_addr_ranges is
    * based on the actual physical address, that is, the address after
    * translation, if any.  
    * 
    * If system is configured to support indipendent address spaces by tagging such
    * attributes as MSB address bits then user should consider that this task may
    * be called with tagged address and translate address accordingly. 
    * Ex: if secure and non-secure transactions are supported indipendently i.e.
    *     both can target same address without affecting another then tagged address
    * will contain <security_attributes> as MSB address bit. [0 => secure, 1 => non-secure]
    * Typically address translation can be performed only on the untagged part of
    * the address which can be obtained via master_cfg[<master_id>].get_untagged_addr(<tagged_addr>)
    * after address translation is complete, it should be tagged before returning the funciton.
    * This can be done as follows::  return( (addr-untagged_addr) + translated_addr );
    *
    * @param addr The address to be translated.  
    * @return The translated address.
    */
  extern virtual function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] translate_address(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);

  /**
    * @groupname axi_master_slave_xact_correlation 
    * Virtual function that gets the components of the ID as a transaction is
    * routed from a master to slave. The default implementation uses
    * id_based_xact_correlation_enable and associated parameters to calculate
    * the returned value.  When a master transaction is routed to a slave, the
    * ID transmitted by the master is transmitted to the slave along
    * with some additional information in the IDs. This variable indicates how
    * the master ID was transformed when the transaction got routed to the
    * slave. By default, the value of this variable is same as master_id
    * However, a user may override this function to define a custom
    * implementation
    * @param master_id The ID value as seen at the master
    * @param master_port The port index at which master_id is seen
    */
  extern virtual function bit[`SVT_AXI_MAX_ID_WIDTH-1:0] get_master_xact_id_at_slave_from_master_id(
    bit[`SVT_AXI_MAX_ID_WIDTH-1:0] master_id,
    int master_port
  );

  /**
    * @groupname axi_master_slave_xact_correlation 
    * Virtual function that gets the components of the ID as a transaction is
    * routed from a master to slave. The default implementation uses
    * id_based_xact_correlation_enable and associated parameters to calculate
    * the value of source_master_id_at_slave.  When a master transaction is
    * routed to a slave, the ID transmitted by the master is padded with some
    * information indicating the port index from which the master transaction
    * originated. This variable indicates the value of the part of the ID that
    * indicates the source master of this transaction. By default, the value of
    * this variable is equal to
    * svt_axi_port_configuration::source_master_id_xmit_to_slaves corresponding
    * to master_port. However, a user may override this function to define a
    * custom implementation
    * @param master_id The ID value as seen at the master
    * @param master_port The port index at which master_id is seen
    */
  extern virtual function bit[`SVT_AXI_MAX_ID_WIDTH-1:0] get_source_master_id_at_slave_from_master_id(
    bit[`SVT_AXI_MAX_ID_WIDTH-1:0] master_id,
    int master_port
  );

  /**
    * @groupname axi_master_slave_xact_correlation
    * Virtual function that indicates whether the ID requirements for master and
    * slave transaction meet DUT requirements. Typically, the ID of master_xact or
    * some bits of master_xact are propogated to slave_xact. Also, the source
    * master is indicated through some bits at the slave transaction. These and
    * other DUT considerations can be defined in this function to indicate whether
    * the two transactions fulfill requirements of ID transformation
    */
  extern virtual function bit is_master_id_and_slave_id_correlated(
          svt_axi_transaction master_xact,
          svt_axi_transaction slave_xact
          );

  /** 
    * @groupname axi_addr_map
    * Set the address range for a specified slave.
    * If two slaves have overlapping address ranges, the
    * #allow_slaves_with_overlapping_addr property must be set.
    *
    * @param slv_idx Slave index for which address range is to be specified.
    * Index for Nth slave is specified by (N-1), starting at 0. If a value of -1
    * is passed, it indicates that the given address range refers to the address
    * space of the registers in the interconnect. The data integrity system
    * check does not perform checks on configuration transactions which are
    * targeted to registers within the interconnect, as these transactions are
    * not targeted to external memory.
    *
    * @param start_addr Start address of the address range
    *
    * @param end_addr End address of the address range
    *
    * @param tdest Not yet supported
    */

  extern function void set_addr_range(int slv_idx, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr, bit [`SVT_AXI_MAX_TDEST_WIDTH-1:0] tdest = 0, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attribute=0);

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the AXI SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the AXI SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the AXI SVT
   * suite. This is checked against OVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the AXI SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif
 /**
   * The method indicates if a given master's index is participating
   * based on the contents of pariticipating_masters array. 
   * @param master_index Master index. Corresponds to the index in master_cfg[] array 
   * @return Indicates if given master index is participating
   */
 extern function bit is_participating(int master_index);

 /**
   * The method indicates if a given slave's index is participating
   * based on the contents of pariticipating_slaves array. 
   * @param slave_index Slave index. Corresponds to the index in slave_cfg[] array. 
   * @return Indicates if given slave index is participating
   */
 extern function bit is_participating_slave(int slave_index);
 
 /**
   * Gets a random master index with the given interface type. The master
   * should be active(based on svt_axi_port_configuration::is_active) and 
   * should be participating(based on participating_masters) as well.
   * @param axi_intf The interface type of the master that is required
   * @param system_id The system_id of this system configuration 
   * @return The index of the AXI master with the given interface type
   */ 
 extern function int get_random_axi_master_interface_port(svt_axi_port_configuration::axi_interface_type_enum axi_intf, output int system_id);

 /**
   * Gets the number of active, participating masters with the given
   * interface type
   * @param axi_intf The interface type of the master that is required
   * @return The number of active, participating masters with the given
   *         interface type
   */
 extern function int get_num_active_participating_masters(svt_axi_port_configuration::axi_interface_type_enum axi_intf);

 /**
   * Gets the number of active, participating masters with the given
   * interface type and dvm_enable set
   * @param axi_intf The interface type of the master that is required
   * @return The number of active, participating masters with the given
   *         interface type and dvm_enable set
   */
 extern function int get_num_active_participating_dvm_enabled_masters(svt_axi_port_configuration::axi_interface_type_enum axi_intf);
 
/** @cond PRIVATE */
  extern function bit get_address_shareability(int port_id, 
                                  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,
                                  output svt_axi_system_domain_item::system_domain_type_enum addr_domain_type,
                                  output bit error
                                 );

  /** returns 1 if snoop filter is enabled in any of the peer master's cache */
 extern function int is_peer_snoop_filter_enabled(svt_axi_port_configuration port_cfg);

 /** Used to set start and end address ranges for each exclusive monitor. It adds address ranges for all exclusive monitor sequentially.
   * It means that, it works like a fifo. First call updates start and end addresses of first exclusive monitor i.e. exclusive monitor[0]
   * second call updates for 2nd exclusive monitor i.e. exclusive monitor[1] and so on.
   *
   * This is just a utility function. User can also configure or modify address ranges for different exclusive montiors by directly accessing
   * start_address_ranges_for_exclusive_monitor[], end_address_ranges_for_exclusive_monitor[]
   */
 `protected
2]I6aLb1Jd2/,Ad;f=cX2-@=->K7#bP;aC_AFO^M@YUc+57+5S7.&)?)g?SdL/X<
BHJee8U5JJO/,$
`endprotected

 extern virtual function void set_exclusive_monitor_addr_range(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attribute=0);

 /** Returns index of exclusive monitor which is responsible to monitor the current address - addr */
 extern virtual function int get_exclusive_monitor_index_from_addr(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);

 /** Returns 1 if any of the masters have port interleaving enabled */
 extern virtual function bit has_port_interleaving_enabled();

`ifdef SVT_AMBA_INTERFACE_METHOD_DISABLE 
 /**
  * Function set_master_common_clock_mode allows user to specify whether a master port
  * interface should use a common clock, or a port specific clock.
  *
  * @param mode If set to 1, common clock mode is selected. In this case, the
  * common clock signal passed as argument to the interface, is used as clock.
  * This mode is useful when all AXI VIP components need to work on a single
  * clock. This is the default mode of operation. If set to 0, signal aclk is
  * used as clock. This mode is useful when individual AXI VIP components work
  * on a different clock.
  *
  * @param idx This argument specifies the master & slave port index to which
  * this mode needs to be applied. The master & slave port index starts from
  * 0.
  */
 extern function void set_master_common_clock_mode (bit mode, int idx);

 /**
   * Function set_slave_common_clock_mode allows user to specify whether a slave port
   * interface should use a common clock, or a port specific clock.
   *
   * @param mode If set to 1, common clock mode is selected. In this case, the
   * common clock signal passed as argument to the interface, is used as clock.
   * This mode is useful when all AXI VIP components need to work on a single
   * clock. This is the default mode of operation. If set to 0, signal aclk is
   * used as clock. This mode is useful when individual AXI VIP components work
   * on a different clock.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_slave_common_clock_mode (bit mode, int idx);
`endif

/** @endcond */


`ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_axi_system_configuration)
  `vmm_class_factory(svt_axi_system_configuration)
`endif   
endclass

// -----------------------------------------------------------------------------

/** 
System Configuration Class Utility methods definition.
*/

`protected
M6dFc<>417.>G=)3Ya[6(g1B.H/A&L4X,MJD.IQ3K\;BXAE0R28L()eS9P_EW]\M
;7IVJ5Y,g5PHW0U&20Y/[.OfB:C;ZEAME\S)eCYFC>c7G2S<;[?-([RNaaQc>.B4
O;RfKV(\\RDcbgM^cX-2<.LS0->.?)3BbID0XZFN(HDc1-/4U.I[N4\Q3QHIQ9ON
:EE1c,Dg?d.6(dR5Z8]XD=cDLGL++6aR[&&b2gbe]MR\.^SAJVGfS9A7d23L=E0X
(>TU8I..bScZJcC?QCMG-QD7L5W(YI4_LQLQ&IQ]38P?G79]ed>S,GXa2,K^(O.]
+8gb8ZTS)KYS43V\JEWR/W_P,CLfMJMJVA=PZaH.Z]3De=6MI0#,U7B\c(;9eCH&
7(Q6ZOXH.J598I8QZ[>+75ZbJIOXRL&C?LbHA/N<V,QeWU@EdDM[d.3+[bbS\:b7
:\-A,Q#,aV3EU@>A?L&P(XX5c3RQ.OYHV_66B<_,aOHg@5gB)VcX[7B/7gZe.J/@
QP]fIKfJeJM5>C3L#.c)8=52^\9Y1YAcJR2M1TOQb6<c;ABYD?J8.ME]LD^H3.fX
==IO-0UKJ(=BPd(L5?e&?8#gRG?FMdEO]_6DfUG9)G8[#VG81/XUO/c#O>U5Z4.+
1V7IXdFC:,#c-IPNV/,WHH9,[JGQ.&/e9gfcb>)_X\B7[4F>&2?f,DdUY8TeGKWK
)e#3>D.S1(L]T_3J[f3W&5_28M3Jg/1,P_V13NY2H:K3\LbKUFgC.=KT<9=dY.&?
WUJX?;U>DJS>VC0):9R+P4K0=5bDF0[-\AbGF:)STXWd>_QQU(-1D]BaLg<e8LB1
)Q;Y#Y>1)W,L+T4\59<9QFf&WI8[D_&^>VT9G7&1X;>/S]W;eM<aWXaHaFHd;FTM
S8C>Pf[3J90T>Q\H#7<]NBAJZ&MFE4E7B>M[e2&IBV/CJB8\N@J<G?=.CR(aSe?Y
P?Q.9Y-bZ\.@[FS9]A8CERHM7&J-Z/gY^9c44I]S\AF5X>;9=V>OTIO]Z^O+KEN-
[5RZVf[[b[<^?-eUTAT@Y:P:gW[CDY>F&H+aeC;DNONN]6E9P7C9MJ\HP46QdY6JV$
`endprotected


//vcs_vip_protect

`protected
\Z;\B0U7B]@@NZd(JeX,E6AZAEIB:.f?9XN5?5C)QY75RG6@3\)V7(BLRQ?;7VLT
I-[&aLG->4VV.@(CdG=R[UA\ANL1<#8-=OZ,YSIZ<<HYaPK6[A->\D0fG]#/?YH;
KRM1J5LH5K&1bM0O1F.bTK6DQ(=-ZH^68dQ32>MGNIDTVZ6P5e[b=GgGEX9PUaQe
LFSfUH+#\9O/9[,0+KH-:__a6>T6NYR0)ae#9;<YCD<\]#+bT/Z\PA#ZbWe[+=fZ
<VZf+4d2:[];5CD[;>>]5;;0d(Y/L\(_Ig)MNcG5U;NF8<X^<RGA-ETd,=R9c650
&#g9M#1,R0D<EL<,;?\2f>X_Qd6e/_2UEf53dJ@Ugcd>fP9#_#Pe3GJC\a;FeI#I
Q41/P..fCSE;K=I].?0X^M5VZY:S#&WRb-_5Y21c--PA&3YLY3/][,OVRXD0B+Qf
6^J,\?BV@EY=O;TV#P?faE9_Y)YcV7H>LX[;>YOPDf9R+1H;Fd0b,#/#9(JRZB&e
.;eJWQ@JQ.PLdI&ZQ,&P@J8XR(Y(OO/b>Z[cZ/XE?B/ZJ9VLMbZ,QTB4N,:1TWR.
;cD=5)=97W^(V7>)@VEQb6L5X;9Ad33<NJ_D&(&gC[=QJT4fX:?<#9YA&E_5/H,:
^XD;8:HT0eU=:7YAA>T5DE5LeKP[cO4C=,/^f=4b7FF#,&MZ@U_@^585b^aYZL]D
0(1\D8EE5H06N:?[BO3F6[ITFgP3E34=(WV@&O5b?,P6M(4VIYWS^fBKVS43DD=0
@?QA4)D^\&Za9MERHSI1RGUU_FP@3N^bWWW_8dcP)&E1:K_N2^<+]Je&7-GN4V;S
&3c=K[eWM;d(:H^R^4dBbcd-<VC[0@-RC]WO;@QeZCR<agXcO1PZ9U1c1g3\:=Xg
;FP+a3f>,c]?0g5bHG]<IH_A_#[FE9S-;4;XB,MX:_^/3bWCGD_OIdYW>J.#f=Q.
?=AGI[?H-gM.>2SF)D^<B1EFLI])(E9c)>N;8?@QWD7L/b@<>a7&K4&?JQ+UEMV5
:+VU@<:b9-cD+\)[=#21/T@;NXbHJ6UC@_,bI_e>VdD#3]7?<>TIT1+6RW([c7JA
)EOK?,RVW]Q]f]<+C6O,@C9b&V#)<;[.IH64\IK/TeVJ?KdWd\5^H6,dQfbR2EJ8
:<L:)V59[W0YIb<WgO)UHC9\1K<<^/BV\NS01.VT7)MH(NCV6UH8VK0Z^Nf_T@7Z
aB-9]b5QHFM2AQ8@W>I<3;V#c^e:Y6<=<Y63RbPCfPE1SVW>+ME4eXC^69Yg0_FI
G9RgV8F+(\YH357YX\2V8T@_)G/5UDJ)\9G8/^e82[1<M99;c(dH;#=6^4B@BV7U
a?4^Q4b3bePWWb7OBT+@WS@]EF<E(7J6X7QYCBB7GJ)IY>BOGPDa;NE88<<)3G.I
gO,L8D#OY@QI2\HWaPPg>4OL_KfLFG[[SN?)D(3FgL5&PZ]C#1TCe[OK7Z#gCWNc
X77F@Y]fNAPO+f9D7NN#4NH#,^G(,X5EfTIGA\?DGQD)Ce?_G#^BVd25V[D&3S3V
JK1U&_<(_#1dA@OPH-,?>=d=@O=@>f3I-HR-6]K,EA];8OS7W#g_QMI<4GG6J,ge
LK)[>WG)CK,3DA(LBWNE>&@bUfK#[bc=UBL\X-SWX_D]4W&f@8,&^a4a0GFWd<2M
P.Z1eI,9H9EN6^5E1K+_[]TFaJQAS>IATS[];.?^O3[:3,:CYb0ef9T8&NR@3G&e
+CdTc:Q5<fB^#QE2:cMKGH3..>4b=)9Jd+/?8P4>SeB,660Z>D@P0.X3(H6)c>7>
N^DEG1[322BBEcac;fLg&EURBWO8(=HX9L@T=8bUO1B0Y,bQT,/4^2L4;<^QfJEW
^MJ,2ggge9Y\fa7gE_6?0B)P5B1)>,M],U>.cL&LWY^Yd/[0R\#BIWPc@2&AV@<<
e/<W&^M3?X+23aY[IMcGOCZWRXaKg^]QL]c<>4a6[Q;&0EbZ:,g=Nb45;D9a2--]
Df\X<^-6R/E(\b[PQK\Bb&5a@cL[V_QILUCeUFQ=LeFNdD)gH8J>;3M&),V^K3Z.
Zc(1BGU)=:-J4<D302PQQ7+:YDb6THP]N(^DY9K:&OHS:U851e#K&UY>7BFMa77Y
+MI2X<3a?8SWE(JE]>Tca5_,UaJK632cAY0[_M@B8&&L0JPLHG/U<30KDT;d=Z5S
U#P?0,TbO=?S&#J+35,LGSJIN8?\bR8\d+/S,+OE)7?(C;S[>=Y3773&GO2HU>/1
(V))F0_O,\#;6W0eOZ?,^VScg>SJ];+&<)5BR[<7MFSW43^G[?4fa?9@+6<2_9SB
fX:,85_;/cT;I@+1@4HL7:fe2PV55U3^^E@=(8CI]PJ1_[&D5g/>:J#<HV,QAAf,
XE/@DE/_5FS5/\JX\e.U_9gRVFd/^TURWOc?2SL4]QRZQ]X2L[,E0XYYK?^L]9YS
Z0<ENQE;4?&eC]f>RJ&47ROXURUZ)^2EX<b46G,2DMb)51^:V8FB4dKeMPJTFaI(
&[,Qg<>^S+Kb=0YD7ZcDMKQH(X?YYEgQID()PI&&Wb(1aBcH_cXTb(1Kd(7KKC7A
-:7=CALIL_\0].P\)b1+gR>[=3T.^-J(43NTQDC;I&2gYLN85eS:3)7VD1dOI?#:
_M#=&V\&eUK+.YGOFVB_L/OMS84VYZR\C^d>2)7:04FX--cf+eY?]-MJ#Vd,fL[[
Q_^^R:P3aEbO0T&L(e11<KeM,Lb:aOUE,JZIFHZJ(N\G/[S-VKZ2TEHJ9RKaC52/
)>&)+G&7KZIT&&YAgVYG-5F6XL>7@Idbb79-+M89-I2>O5+6IJA_-Q+I2KR)O7?_
64LMG;:XNY)T.4EURf>_C1S5dJ#K7P=++Pb]FbCD982ONg6&K/\a_^&-+9U>dF<P
:?XE#dWJD1\+ZgJK6TAT<>g4feKX@PeA]Z)&=+54DdXZK+2D5@Z)+-RGeHaP:PE+
58B85;A;/aKC+QD2?YHdNM[B>J1KA&6d9QFHQVAYJYZR)d\cc_EUIX(>7cBaQ+Y3
-HcYJ=P\aN\gd8NY@WAe)P<-C4\,,+5-D</A?.?JGQ?>1T35/Q06\F./R:(/DG87
SUD\O7.Ca#C0PRdHS.<4^8NUU.-V5-J_QM-W\FYXHEIP7\Z;gf3K86XA>=K)XI7T
88U#[;A&YD))Z8:^B6R<LWOGQaW_@:)PaU7c,AI;.-S+801^#W5,T;D0:Hd-cZ81
A&EPXZ58[WQ8dW]6173B22+S\WZDe@?(8S@_R=[5F[EZ_01GSc<7B73O7+@;F\Ve
..e04_7\<75;3K13.8?.^G=69[aB#1MY_LI-+MFWHI\e:#^WTR2U7-D_Q];8Aa[P
1WUQcU73ZSH65J6a)\B4^MAF,;QE^a9>6d8Z1)M7WcR_C_S71C/9G6T]c2gUEGEJ
]>/S2ZQLUK8UI+bBSD?AIgD^=E#:5+S&Y\ff\-Y[;?g2e:e@XLaJ:3?CBV89G?<1
)]JW5#d12=&ZN)HWF#.K;7YOBGE:eeD1:^I<:ed9MfeR0AD987dDVM>.O?@K[:O<
L@724X;-^.4(/>QPO_[\/C1[6G/eTUBF(Z+?fNMf)/0V^<</[N/fcf\+Q&CP67E4
eTfEGSDTUR343(\5PS@X-.TB058Z:7H>b?(YaD59:.(XC)b)?IL(Bc>8EEMJ>S98
beg0)SZ]9>N6=ce:8R7?7dIa&@Q.S37TOQ:O)^eYe]13KV3I-1&e<Z7]S^\6<-<0
\OF4Q6K?ILD)7AAD6@681FffaO,A#ec<J,8_c,TB1)3B@9@F.GY8L-[DB0(>:D<?
CM(A.(O=2:V86W#\9#cceFAL+c#VUV;B=aJ)[/Q,ICM^+3NbZ++I4V)?@5/T@];c
O)]K#5<D+.9BWL@WJ)PgB\FbJ8R&&4[,d]CK/#^.6E<O3?:F5[,>QbFLEPDA:CdX
A]aN&gCUcWU0GMXQ(N&<@a+L)M2/O4/++=WG:aT+BO=XY1#Q&2gda7=YJ:L^]b]D
S:5]:35P.)<>@-M?#\da-#\b[.@=c=b_(QQ,M?d[H3>RE[BdOa19[B,]dT?WE(3=
^eGX^K8Jeg4HIS[D4NPL;K,08JM=;T/dW_JHQ/bWQU\Q(A,,?WXc?Oe(=eBHHQdW
<0VJ(##?a@Q[:@,,-(Sg0c-d)#^3c^,Lb^F,AfDK3XI/@^=#<K2b4I,EFM,M\WJ[
8fW\\Ecg\RX3)bAYV3A<KcEKdV)F+G53e8-;831EDdCg4RDAD#fZG#aEVMZ=Qc0A
H.PYL#T1O9fUWDD]8_S5>E?=?1G<Q?0;#;M<);BR11KRX#eDC-X)aU21.67[^\KO
^4<XM?6b9@WU+AOJ&[L6.Z?2ZcDaVHg/4#W1/<,7?6>:94Z@.V:DUR@GJ]7gZU[4
:YL:B6G#J@Lgf.KY<c,PD+=3D@0TfT7gH4a3-<S9=]dQ)&.]S.T:8,86gN-[)aSG
0,N3,@^:SbBUfV(:bc-b@GVUS(VVF>_bQ^U&CX5+.J0-G)4Z^gLO?+K(-5T0MD6D
2A/e_Se0H/H=c^KG3HE,N_,[@Se+P:c]Idf5(G7(CDY2XB:WKIWV4X/O8U,c8WP1
FPc-VHJSbK1\fa6?;I\(cV=+\_Mf5BCe@9dZB1E[]_SD;>YV\TO^3R9(TeM-.UVN
d6-:<d[8@C9BWCMMa\J8dDUOB8G)?B^/,IQXc7,Ae@.=[BY8+]g:?Ud/)+9_XC^H
C/]:15FN;<2>M_#..UBDfW@\=8VZ8H5=,6[G[E,-5b6B+))#bDT<f?RXQJBbS.1J
Mf(?N^]K@C]c/+YV(-K_Q3)TSgL8(ROG0)G&@M>V_T2K]3Ved^_23dZSQ:J.,(c,
3DXAA+<E(@J+I/ZU-JB5:7AX84JNgG7P)>T<4JTaX#X165,?RJL.cZBO)Va4c/]7
>#6g;,Nd?U)8FFNg]4^R]H55ZX<?A\c,L-.<^OFZOV[Xfe@[CLeA<__d9JWH[FJ2
b1,L)5DS^5V-;P2RKXIG/K&;Lf-J[b)A6?Z2QAT8R(Q5c.22FYV\(39D(O@?<EKS
5gXLP1\IbQ4cH<gIMdX10+_Ne(D.S^T^]gE,.F?eH<:RcHY;/NdHT.c]&RB(+<Q&
V4Ua/5#g(fGXca\9dTOO57G.-AURZfB9:6>)G@418Y=X,^OGNc<e8XZ1g&<Accfc
gg4RA\H^(cGJ;XC]J+R\WVM2_PCQTM6dG]TWU/N[,P<[Z/G8)dOS^\9Y<1/2W.XH
PQZdVNA5XH^bM,V>c?O89&?Yf=Z/;Q:PTI?3dI]D^b11DDCF_-9Zb.Q5BP-J,],d
\P:d7\ef^1S[QQ-D>^,N15?V=NOTD1VM6C&@UU:[YPX(1eP/YQ>,>\@f:O=)@34,
HS9O;-[MNX\^fZd.)91#Rgc[Tb<3>WFHJF@b7M\R+@b72Pa4-3/\+=ee.8>:Qd\T
>e?(=\WLN#b\Qc/&(M+D27^Df:SE@d9d^_0c07Z0?ec/\f@T1#@0f=K.MEI::O^H
#.PO.QXG7bJ:W&CKDOPdfcY8\LMbbL1>g7=cA#B[X2g>>\b,@TD,>?#Y0C_DO_cW
(d64fKU9@IA\H=;]ATT&4R.M9L/4:c7-=C2Le-H([-F_NRfZ=O:[a6IV4^HTe(C0
W3>e5V_1KAOMYO#ILa/=XIK=?.Y?WOdEXe/Jg0=dXE6?558DFLY-Hd(dM:X#&G&P
BPH+:43U4/:M,RN<NL0J58bIa<PSHE.,)d>B(BgQS&X^aA1ET70,P0E_2)Na\\\0
Q+7\A6NHU?GIK7:Z2[/J9feCRI72ZL]X-9U,(5GGS:eR,^#S]Y4]0,Y\YOUIaDc7
S_W@g8e.&H/6=2U^,NT0B:977^L2[e9dI3JP=4-]T??_S_RPR.OMTgIGA74a0H@b
0_?DNK/,)d+&X5C#>7dD@cIf9G/eUK_VGN+01^#aAS2PP\^b2g1HV;Yc+.78PJSC
6L7eW0GM1B=LaUZ)P].B0@gZ5Ed2?Y(_HJ.eNcK6KT-Ef^MF?]Y:/6#T2PS>.I_A
Gdgg4,ffDPdEUYWT#KT[e2)&VD4C[2cIKUZ&bf>\CQS:?+XgH^gVAL5^J4=bGK7-
Y\0ORG[D,>)F;ZfAYHLRIe1(?6H)J2K)BdWb46e_KNZ6R1OIdC2FG<AbJ6-^SHIL
d5QNf,(2FBbPUFNKI:.C#?_?.WB23S[U5_Mb=8/371(;6,g/7Fc)?0;LAJ-g8F__
FCA?IWLd2;=KN0PNYG3BAK+6;?>QM-MC6D8J@P2;eTDLMD@^OPa.7.XW2.96;.gf
<@:Y-/)KZa]J+QL248ZM,.9]#L-2ACTNY04D)a]L>Q#YK-VEMTC]?2#H(/^H3O=?
#@(-L-_U1/dHVZG-7eAC#T072);X-N75Wf7SZU^W<eWA<GB:8[^5:1dCUVbI3CGC
<f:AV)HPJ>[6c13c4,84c68KK^&>;aKM@.N/b35F+bN7Xad=?5_XM=/cd<D6V]ND
8L9FWGcf^fNA#cAIMW)_(]R?8<.=?bZ/AJ>PG&=3VIYB,gV&.]J6/NB.O:>L?UR_
/1:VQA@V6XFHTR51bKPN[^2[-TUJ:U&7).-Jd]b:>^)_cK\DF7<G9QZFMT3?80:S
V94EOg02ALQ=QcBU(_D?8&=Mf<)VDIG6(NSDG]X#T/A=-?-,7@.Q&=L/UM>f?AVS
cCIg1FP(A#.\MKPMANY0N9\5942cc8#AIB-/1?d^^Xd36PL_eD>W#=EU+04;/SGI
2;FXb1Ja&=]&_TC>L:b:4_E)=J280geFc/=H,e[+_8X-RRIL=UP)0:\;)Tc^=3e?
T9X,&5Bbf0g_5I]I_(I,&Y59[]2CK^fLbO8g4=eY63</N)57Q9XU;PHGXA99:=9D
](2P^<d#>7Pa/:,Cff+aNM_YegYUU3RY<8S<B\^M^2GZSZT5D;IE,.JEg/e)5Xa>
SaIEdKeB[9OARR\c5TYQBebb4=;3>L;KLPQd&\IQ]VE;5#\1;=@0#V@eP.N-VSfJ
Se=\RX[caKBa=+60.BBMeN3XU==I<E(N)QW&X]DC@<#E.eBf(#;aFT]^5?C,00WS
1I=1,=Q[GG_gG,gFeP:g[B:46DG;1)bW>eBHBI:PPS@N(1gLgW=V?b=^KT\Va#eU
T8^SX4[>W[.&5GJT^^?+P&X0QX&T,Db#<1B:^dRUL(Z)9]3TL&K-O&.4)/TOQU72
_XY-Rb^K<U^6(?ILZc]88,TE#-74?Q/VOG8[@H2fXH\L([VI+DCK5-79PNP8FWa/
8BXG+.0YP3Y3bX9-L^+C]V6O689DZBgDQgD:0@,6R)^-^/1b:/La[LJ7RJ##+)WA
;I-1I&&?QT07(W.M1A9ca799@-+R?D9ceZ4b^H>E(MNR&.Tc>/_ZTfM;9:_g4]DG
HfIECb:a27@e22X\bZ[-O-0Vc<5gMRb8(>NK[a=-#GgD3EV]BFM&HXWP_CM57:gg
.>F-J+#E8W?4UOG2e4PUU^U70?PUQ0HCI2+(5cRM.T(>29E>[+FDJ&O:6-f([_f4
/X:EALX&N.eb?/.cDdEgCW[F;PI\.O8_ACAD6<ZbN48C^LR(#b=)GX2\c6Q0W(:g
5H=@S=>e>&P9U8[R319HWW<WfI8NE[^U?(A7a=N6>#&g3V51QTD0g:J&,O9ZF&VT
?b&5:f0GbECc6/@<:4Kc&8^-E6CER&5/Ye1UT-_=>_f&F+D5)ZVG4CK00O4&5Qa/
TI36.ff1VL4;D[#C_b#Ua3bXO_\6RSHZ_CcU/1L;<#>Q9If\#7<V3JKD(#[KP=a3
:D&G.0EV.9?Lbb^HeK_/e-[-f6I=FKT830UK13,/?RPGbN5)#=SQP9A(D(-J^3OG
CHFNHR6BOF]NZX[YT)3VQ)M=+Qg8faV(\<#c\8(L:Y]>]d8AAEFJf30L5U7>#g\W
E>)=fNg_@TZ6D&:0aB5&=Dc3fF028bRTd+#[DX91M[M1/Y3OYOW4G&_4>3-M#8AU
S9+9A33U_bE;(TE#=A^\=7E;@&f\e;055;-KTb4gPLBW4Y<]R(P;^ZJ#ZP?>G29#
^36X29&?X.)_AFM=4<I5b[-EF-^UIK0&&2<I4BO7,#)g?Ha1>,..aGL&^Ta;L5V4
TgO?LU=DEeV92X=JZ)C1[I;#eIQ2M]YV\2]8fYNZ9];(::YZI0dHK^Y4SPb/:-F@
GD^b@X(JCQCG^C0a#W7W5T)Y5NABCeM^+RD7I;a:2N;Jf:67X=#6H(^T7G:eEQ2^
[B1>\YEB<.&3[LEJ?2gL&[24DfT)]N]QMFW(^=LV25+e>VCe/SA6?0e2D94ZA@>\
00/GQCKOIFF,6L4cO;TN#=8^UdCE;0?Z[+O/=]=XZQMR\1CC@A)O+1L(.-RR[;K/
<\#+f\..bC#Y=GL(gOZ/Q@NJN?/K1O<IB:R6bV?PBCO)GFH:S./\:R^,aa[#FIC4
fXK14N;f=5>RP.LQYM/HU(b&U08A7.QB]2LS[S+][)>FcCG[KUZQ=98^=VT@aLU4
(W\A#CSDJ=JOK/V3&M<,_C6&9[45Y0@E[-9W)23<LM-:f@23c),g5#C@b[;:J@9^
^bS\81J9^_TdN.>4.bYN<LAZc96SG;T??cbM0)YdNec087R&TR+.EPULWA&5;e?L
Vf25T>.I?43\c\gGQ?G-[T#H_>0#&\S-bX.]\#Y-Z-3/XLR0ST#?LRcEJCI/+d#)
;,87K&]WR_4GR^E<aeKAN#D.4DJMC>CTSdUa67&WVEYdX8.<>MA>L1=a;5Y@[^H_
2:#(K08VA1cO#fL&R>3Hf-a>A2A0MADQ[._0MOLNC;>=HRKL;fe0=O9);.]RQ@0O
L^dM(>G.78DD?(4[9S_<N^+U57E<2fc4SG0Oa/CJ36;[^IRSfFG#,Pf(G6O>cF1Z
#a5=64XeM80KNJaN_.@]MZMY+R44\;&NSZUPYT0RV_^:WD^C;6AQ:_A,&bd_<2K6
;<:UWG[PW-KNQ47W^+VU745F5D,S.8LdDK>6;M9a:]OP>:d/KCC+#\g]@ad[JBNA
HC2O>O\PEV>1Y@:(9d92P&B,Be<,:1A6.@FX:\eOR^K5GR[GF]VVGG&a[0BQa)08
)-MeEb/55a)>4&e/US>H6-RLU3<Z-9R+&UC:+(9CfCSW39TX6M5XMX;GWIIN^8+4
c4<B,><\&C#L]X3J4=:P9[YVN6+g2J^P.#8-f?J][RRV3C2FLP[UA;98F,Ug6[(^
UV/VILb90U6];^KNSd83fSa0?K4_XOICPM:=MU/_Y^ZX);4B\Xa;P8;[OFc9>PNb
T(CWLLg=L\@TDN[0UNeTE;2P:=9\gA7C.-O8e(bGd;6FV_P?37>dC;GaTZ<JN8GR
)F?=H=,_MHBg]JS3&;V7S[XGT+ROW[:f]<?N\7&YCfN?IT@a)=RTWB1cB-R<(.>/
Lc,,I/784HbF/Y8S(#F665=)^,YX_5.7LbP\eOLU[D4)g2=Q/&U9)7g(GZGVP.b2
?2G4=fDD/2]\U[/Q;)T0HE=.N^WZY7T\,7()HEJZIdC9G664OQ4f.NWaJcdY>922
\Qgd_5(F/GY<W<7Q-O31Z2[D4?E;NTP-6UWF)4:Ie#1g])bOZ8K[b0dUHU=b/O&D
9W\TS14E/Ae=H&.O:8N^H;4cFa5-RF124=c;_Ac0Z+M765a7TX#-\d.0#/(#RSIL
4C<&--Zc?=VLA6WC4JX\@2R=_?7Jg>]U&E,6ECCRYPE6-O1+#>XSBe7=>_7=Id71
<+FY8.g6Db).4GdB,[[O?8=4ME_BE-:<f[_S<:2;(AaFNG.FGKK@0>c20G2;(F;a
C1EIeK]GQ)Z:H6-[2=AZZE0R_IDgU:D8]WB[\_;QZ([>32C/XKUZ-8Meea>_GQ<@
YBMD5c1ENWU9E4dV/(7)P(I/(VcY7^2M0D2HYN5QEKWgbA]1SK(c4R?)I^1dB<?&
HR>F&TQTJ\5J=(fdX<aLS;8/91c]WGN7^(V5cO&Z_Ze.?\2AZH+-W?(J.8JaS>,E
T&-,ddFCf20AIa5;H_gDaOa469W-,[V1[OI>ZVc3@0CdW[dd7B;>B,eU))<A+VJ6
K(\gL5B=.-#WO8[^cg(5=F;1bUcBAMGG08(YEQ(H7KP7Jg[QU#^AALJTD6;3^f;/
DgQ)a52-7+>@F>:([AEQ[4WJ<37_Wd5NYG[F6a<^OgSa&1=G/1.PbW2:?U+\WWX1
<B027O>DJUL.Z+:;g<.>Q<>/?6D#fWI>_1BF6#CYE0(5P]@6AKH8;ga+&c=BGg62
Q#F;OZFI]H4S@gF\SQ(f6<cg2YX<Bg0[W6^H,?1M&-\eJ#dD.\ZE+FT(6BBWg/@8
H:BD^)d?22bRg9F-MGG?&-;C_.e6\5-[/eT0G>gA>,Y3YZOPN(^_b;g.;R@_Y+M+
^1OHFe]G?VA7M;2&gcD(+9cBJLc:eMMOVT&U8_O(I6K_1OcXb(,5]]V)[Da1(aK<
Y_(]8eVMfB#C70<=WA=gY&QP#C>7W2VJg1>?aVc\3f=d(.EGZB5MGf:].Y;5#_<L
3Rc(ZeTKHBf66NXS\PGNJ8VX(0CAf>\W4d587^1G1_5BH\F=HPW+(_82FUZ75\eV
E--0I1D;GV)3YT^&[4WRYd>]D1O&^VDHa[Kfb.WCBdFf@Z_#D(@8(^]S[T+T:-[9
cV1O1#&MK203Ted+#,W=1#Y)&#D^R9Ze+8Z,3=JfN?,4S30>8)<#fRNW;&F8JWc3
>[STSPA&AI(7GC(A=ZWJ^7bO.2a?dIa?J1TPXLQX=&UMbgb6]8[\cW?eLW[31VS5
^Y[0H\EZf7Od@^VJ9L+O0KK;eKL2>849+d>0BL@EK2A^Jd#L?Q#,8L)4/=D:):;_
C((a;R4KGF_C5QQS[4FTO#M]N[6FHR7FYU?MWRfRbOSgK1g?_,&=N0>9#4UM7Mc(
^HX#gAZAd0>-2V\6^59M.e8d:?M&Q)R7D4S[-/e7^&G:@B2Q<DSM9;&07H/b0_A7
:TbLK&.;_W0gT\@#SI)=G_b/V#A8dQA8BZ_a]F/MM31HU?:aN,8YOVM]I2RUF/dY
VQ[X5K?#;#N4(gC&L)^LdWJY@_&V:JdWd5L#@9BSW[,GY2K;[T1c(9eW:UO>QUQR
6Ac,aKQQN;?FI6#W-PS24g5[Db_VAONbO#f:&MCWf+MdKF(X;DJ_H3PFd<H&B>JD
=GdY&^[I6@aTcRL\4QP+Mf=e&Jc;VQ]?B3XX:[X-(+/39G0a-Cg.E-QBN\WeY3@O
(TONbEH3YI1I-ZDe7R=,eERa6RI,=7F<15;08U02)DD;D-Z6b(;BU8RYc,>(TgG@
:Qa;EMg7/?E]-Z>H+>3,9ZQf^f&FB=U8PYBE]NE5(P=W8-6>R?9<SG0V@T6IbA@6
:Z0<O41g^D,RS-MI?WJE[=(BQ8,gbVA0gU,:d1LJ#TZg/RYDJ._J8f3]a1>ebK6&
RNCDNG1GA6d?-B[ZUaT35<5^9Y3G^WH6M3fdIMQ2V[Z(9:3[2S03SK&-C_F7Z,:d
^.5V5[AT3dN6Yc:8BUK)[R4&8]fMMd[Q7LYHgK=T])a2Hff_bV4MDaKa>LS>#:Z1
7ZM5VX,d+)Q1P].ZgB1R1g+9FS7_)=.#d;Q#B@FOBAXAc1FWJXO[)/BQHU1I=DS5
8O6JUPFEDTW5/8@V,SRWAMKFg9,,f>dcffecSY]H,5F^R1<YPL3b0-(a;SAM3FX;
4>L[)?cY&)cIY>U-7Y]-DLB<8f5^g)PGf2_MFX[?0XYa3=3Z[AMb;+Z+e<9b:J3^
Fc@3Qa4(;SBQ+X[5AS/=80_5Td.BTD?gQ[4@_>Q]>c@&T(LNb;N3KFJYBP#+4c@J
LR/61ZHXYE0<ca)2^2:HIf^R5TT/T6P_H9<c:0I@BQ#^_<Q7PIF-N468G0.J1gFa
MC0RPRL\4Q=SXR0PI_1_,:[TcC=R[R9Y3:9F)##<P[1=]K^[QcPU<:1<f]QE1072
/a&NcOIEAS0(K;0-DOK.=27_+5HAFZMa&G?-&S<>O/.<<;[_P/fY5=eVUe6E1YPZ
VX14-W3&8,O,_)14:4R-dXbN+J6d[9S/HA130A/La5H94)F?SdOSZ9+P5XfQ4bXA
1//5S:5N1^RWZGG=O10-b\bVL],]@QVX+Af_[bAU)ZDbZ^\ZO\DR>:\IQ@Nb;,R,
BJ9HHg<G7GS@\Y\F9MM\RLJMY3-S51@\0)5V>[#;&/;4+<bYO<::R^eOXadH>Q-S
dJ6/+-V=^O)P#MPIbPg7K3JOK^2#>d7>BOCHfF2Og;MUROGYaZb<PWIJR?[/JCa_
X.OFE+0M6+Jf-_[OB@WXNb69\5.gRO[JUUUCgf8c]+4L:0&[SLNFLWgcG97^UG>[
7^W^[f0&MT]^RD.3R:6JKb?,IgQ6<dH.JgNU;W=B&(;O7,cNMC8&^/bD[_eE0U/V
1ScCN]AXdBFJdaXaf&E4bX/U/^L)8;2cFH:a=;aU[+Q7FTR\17,H>,NWC<)0?0Ye
K9G7DH03.bM@LS>&^^]YB+;c>:)JcdD]_Q4;2-OC8\/9@]&[)KcZe:I_bJa6GM&T
N:?\6467T3B.gL2\9L7@_V>3VCX1NW0eB6O,CV78P^S)RSM:N8K<NVUKdR;_.>51
;YNRDc28T+R=dO]YN#2<,AMQ_U<Y?J8V94QZ88+fbaBIbWS<S1G68dP?5><O?Y6c
9H]^N<,.S=)1O?<=b=.Q?[(,FM#^bV9;c;ZBS04ef@_BV>[d1)#J\;<)bYHL^aXf
6QBT-;JEccAWP5WQP0>EH^V/D6R]7Q6&U?S6EBRdQQ.GXgCAX:\EWX60.H[H#\#@
2#M3@O-@g7CC@KTY)D@:.:ZWLfEWfB/S(g9#R>2O.A]d7ZFU[(X\c1&&46FB.394
3S&8.MTKMIXXW^b^[QR&1[V718PHT5D_GHBeB<-O_ePLg0WdB+T[IN2,I19I79C>
)A6JYV^F6V2=WRO;GBU^J2bgA;cM;2dXc_BMY.EB,(+KA00)M5^^1.,XP_8([c5_
X&0YE<74N^RO?@PDOJaF<A9g:F=/)3ZcaLO>R_#QYO^V[e8BX3ZB(A0>1M[0-Jg[
CR(;X7eeUgg7+4\8H?G(H8=,\We#Y?4T[8e1(>=)-7I.bL,T5&BNTU2.2_,U,\3\
E4+?F/?eQ)^>bWaPc=G#89B.(G?KH[f)[:;11W==JBKGU_ATQ,0+LfL#0Eg=JKG9
-]]fIW&PP&0ICM0SQ./0T#b:<5QN,X-7Jf:X3@?fJ?N6]e,N:#<3:D95cJM9T#Tg
@B<E8F_MC;464/EF7bXQS.C^e28CVaB8c./VcF,C8NgIAZ0T<+@8^QBTRX1H)-74
?<18NUcZG@+6TKcO@C83#^68B7(JZHfSZ6<X:c>Z];37]-,5K.F]>MZHV[ZZP6M0
3U81K;dIU)JDTY(>KPA_f9NVPP55](#[B-A/g#X7^+4\E-HMN]8,L^e[JX?]BAIZ
AIVT4XQ/a@CB7;DdZaKYH,WD7c<Df<))E<6K40efHSF1AYfM9XL-\8KEJU5XJ<RI
CKBM@c>7\MR]<d.<_^Y-.3KUBa;7F3f<FIIgV+]1b-Y:6cI-:0Qf0-Y56UI_KNN/
D6_DT?7g[#AgXT:d2<5?)&M<QWL-O(T\SUeY22F,OR;C?_RYC:UcWUG&K_()Tf:\
f:T5Aa#D+M/W#]1B8bTL,PfLd7H^6\=\4J_M;0L]MfN@EJ<3+6_P;N/83K&C6R4;
XA5b)3Md<KfcQ?^9g_7eV0Z,5g9QZ#c#G/]LU28g_cDD-6dEAOb1^U(f=[G8M/-d
4#dRVefERC3ee\OGXL66a2BIJW33^YYO#/B437#J>W5d[UUDR&Z3-GbeXG6BO23S
\<.0d/^d[ORP83U7G92S=KSALO6dC>bDZB#Q&RS_[.2)H-,72\e/8.:^=>b+/P-?
1F,L)571:W5INgOYca42DS#560VVLQ[TCFNbffJA)G0OHTKAO,X49_NL#&B]&+2#
9?e^3A#)8F_)&(Gcg])J/-(M0^G6Xd#d6d)00<\[ONZP1J5,U1MR)S0g16WY,\CS
RW<I6RGRS>8/K:B6X0LN9a)UW1^eY;fK(W>FWCMKTKJC.72K575O+e#cHGG81RSY
dJgLHDXRNGJ3WI_GUBWaS5]fC#UY6?.\O)@I-G;Z_?67.aMSC<&[a(N9>O,XDS@b
1]MPECdL)O,>KbRE18,_RJP9F(a&f-SIdV7=6>d&-ZCeSd]4:V4Eb-]b@&[g^^&J
4^0P_K7E(Xd89ZH_cSGI-CQ,BXI6<N&1f2aEEM)/gONW#=a\],K_1OD?+84)W823
#)<BJVTc1QP)0&FY1&D>F?D^&/E3PfD<;[\_C@A]V4FZ2,.a1a7RDd1#bGE2M#&-
KMb,?&IX8I\SV(?gX]J4@K,/C]g,LS6OWDVLeIccgH[=,PE-9&ANE+/)62VC:5AH
IZOZ3<3/@#aBKXVH;(YZb/YB[@H3-&/\6M@^e<+dV=g6g40T]I>d/OfLS:8JRH;[
bUJ(B1;1[B/E-[;MDX#fH?,WXG9D-SbS3eg<.PY,>)K4MLB][\>A?\?<][R9);EL
Y]J4W^I2_2JJ+Kab@&6F5]W64L\L[=P42P5WH(R[+O;YcI:<0E^+AOP<S)I(#[XO
9Mf[L2BZN^,[THQI^_99J(:V(-a#?S&)+NVT0Gb[c30I:548\2_OgMKV6V1Tb5BJ
ecN]Y=O<?KIc#P8DCLWfR&<X)H\-=/U40bU4@L//6Q]F._.0:F/8:M.Z#5eSF#T-
)Kdf)0&G>E.-[)eQ+/dH9R\-X]1ER,4#PO&ce&3ABI4(Vc=/_eY\5B:aTI@S9d1G
Ga/-cIH>6T9BI(DD698DK))a=4ZNaP)SO7@=;M;;;_N;VbS@P0Y.,C&1G\?7)[PR
5D_WXN>1)KW+OW8e]XF=Z4bGfJVAa84&MTCQ[UD.&g951d^GTNB#VLQcUGWRf9Og
-4O37BP\J-(AcUDYK;BU1Z?]/:\[3<OfJ2J8d^ADeF-/O#HC9MXGQEOGd0<a7.C2
N)-fVY8UX4+f8/ATHaR:4ZDZ)a1DW7O8H))H[aJ/a6ITgd]/X[>eQ/VONP?X\JK>
ZQ,>^Y0]g09N>-(O;U/(66ERBOb/T5P&-VYODPFA9KQFQd3A#8_X+A/E9(?M2HV=
YV.V,L4g@D5TZ_CT>D.4S5.,;IgV[4&@76a_Z0V6FR7ZLZg..6T\&K3M:Md9_JI5
M.-,+6_ZeAPHY3?[d#MCL>UG-ZBD]-JZVK.P]D:Wc,gLE2B)7V&1>7=C+FK]NYM4
<H?8P2/DJ#d\>BDF8PQ[aXVW+@,JXQ,ZAWATO85+_a5+)-g]G?J],-#R..bJ9]PB
WXQ)aO6\0>\HHNJ_#XC:g/XLd)GCG;e1+RdYEP)UD7[-9aU.ffK8R+]MX3=Q:&/&
T#Y9b([+LR4[E>C>a+[Q9+,GEH\Z:]f:P&#PN4H?ZQCNKK.R#CEJZ]c5F4gO@0Q5
D=DD+P/YP&,VM.>IeY_2SX>U7Q.NUEVKW6A<T6aXNQgWbg>Na)EJY=?T^T+I+4\U
VBFX)NWe\Pd+_TX^KVA_?6dKS8>1T/eKI_Mb(&9U.@A@6RS_2P/bQdKX>Bb/^\1-
:gbTR<K(.Z(,baHb0?V:9F):)A;VcdTOX>3S]H]+0#_N>BEP_d8b<3bMVU/FfWPK
UV(eD^g6FOZSf],b9XBC94(A]2.9MDbba:1ed4G\NR<,1:8Uc/VF.C;DASP<9^GV
-+:M298O5L&3[J,J1RP)GS8QB]K)M5Eb5g-X^H=Mb;P]X0B/:gZ5]LcZGB5JaH>D
]+\K_fOKU6b^<WTL0VXDAA1Z88V^B1,8O(ULT-3b/dd=X>g]cIFB>G?K(=NW&L]I
aMPY_-<Z8Zbf#Of>ZGcK5&TO69&eT#+-1ZU?#6HB7;^Q)g5>\6V&^,[?X)Me9E,c
/eVJD<^V&)J#8LQ-\#>P:H:&I^)3@\HAZ\ad/+WaQOO^Oa5&_6gE./KUK[NfR\7H
2HNT/e?SbOHQIbb[QMJD>SK^(A(YDKEb9<g_c60IAI]5]R8]&N>691S9/\&88:=I
[-G;:<+c/WQ594+b@Q#U>6F+^K_1\d@JJWT=DG_[0?ZKN.gC]RJF9fAW1g=YVBQ;
-;)USF)EDKY8BHNZ[)K2F_&Mf,g/-QBCVV_9M-&VY0_(,Z&b)UdH>J<1TS2/+eGU
\J)>Ke6Ue@.GeH+Bg0<DW21IT\;HVgP(a&B6<P;G.\Ve,A,T&d><27RK)F+4Z2?:
aFeYAYJ[_B81;8&R44Y(4@6^7aZ#b#2FdbC7,[a,UW0e#[b(N5ET&/fgZ8D5g(D:
B1:E,W7F18g(:4>2+0ZLT3dD#L?B2:[NM6BWF;()B-R/?&5a[Z0D975WB^R50/=;
c,<DIK^>@7RH;9#.MJ(_AOZ#3_-GE,eDXg])AT=F+cGOK#G,:_2cFQ,A(R)_&BPa
3Y0L;\;JV>]aGF+M>N)^g=SW&e=d^<S<=]--<@F86@dG@31];WLG/U.G.<]H)DQM
3a-<HTYHMSc6GC72]IgQfDgC@#^S6[F?86(,a^E;T.K0@aKHW+?H?@U<0U]G=E5:
^9Y3SNgIF7CPB]NeNJ]Rb(ddCB7S5E=X@1+gSGCd60(7gIUC&^1+IJ;4D2)DfgW)
C8RE91;/IF>YTNJV+b)^^/BSGdD<O8cP-E(_(EX-cUKKc4Bd-9b6EFFIF:1FHbRD
0NC0Od1PbEgG&?c,(;\8R0\J;<GFEeIc-TdCO[3\Hd]MJ7PIYF8+_TJ]BZ=_=)\T
R<#+5dT<\cOV&bJG]JE;L<B7Y9SH:LX,LFbQ\DRPdLMfNfG.7;X8X?\:S,d:(#TM
:Sa-,_RWde^=b-RaX?dT,>+@.f0C<e6/deSOgeR<bR?D[H+TCXVXP^F;=/N71T#7
HP>cQBcXYe^NXWGf,-Dg^35(SUDH<K#8]1?K=UPU6Y?\gF2g05b3]e[fCNLEXSP0
+51APGX2=@^U)01/1P?2DdNI0@]?CA]g.Q,g);+_?+UG<gc^K;EgIZJFMZ9CJLN3
.V-DTPXfD#7[LVX5DM:aC\R=]Y/.8e#D@:75[U]0g[CBI(AI)R]Z+ePBA9,LNB1H
?FbN>M+_5)eKF[Ff^b3QZV6CdPB+QPdb_8]J=cZN;,gM/R89T\ES?(W]11[>\#Ze
VBfBG.C(N3Y11JZ-e)Z?N=3#G93^@B;Ib.TAMdI2+.c(Ka)29]Va(bdBC-IObY,7
P7_Y,7A1.>gJ[_Od-aa1[1)4Hg-MNV@=fe=VGe,;L/X8SFRX<MO6N&;5Y2:.^1[S
3W&OFKKb[)N^DH.a3IZ[O][;6/,8e>H5)9UgYO\=GNXP&-+2)bf>7ND34fH2FR+-
U;acEKIGOSWNKaKXLP(WRR@.+E>Xe)L9UOW>P;X(f:Q:Q4@<T[ARJV9GO1WP3U(F
?<E573&:5&.K&NU<\IBMKUEd\3bICH>;.^OK3FLaN7CX9>fSD6b<E2]W:a?a>(X6
/ON2_K]>4gCdQ)M^C_G^<LSEb>_F>T\1?2c(c3/_?22gMKdcT5.L.4RJW[YX5#]F
?7DUe+NE?#V(eF[^D,-6&M.V<3fRO\QJOg.JEIfT9aD)XNdQ3aRg]3+HI30CA&F]
7eK<I3QHV@/AUF6VFD-GD1&E_/DQL&+_gTDRV.,gKfJZG9Oc;:N][ESP13Og@\2I
BQR4RMF6Eb-<A>b)MW1VJVGFe^eB5R=W]D((P9(MTO,;5?<670CNI/]MDX_NT&BP
aNEeMc()^MGZ0.K7bcY;.]O)0X-Y8\\GTe4/Q@F-=44@1]1JF^(N7O2c7+38[L];
]=V@Z#MIA@agP9>QH^U@fH-,WNI)DbF)G[]2U)(3-JB@IFZ5Lg<TWM@,@aS18?7(
/.f5;&A]SS2CH65&]DQN>9<[>=<;Y44H?)^^+@gO_R[VRIb19=&O05Q)eN>@A#+C
^dJ@MD)@ba=/dPdL:KQ73Ad_,9G\<bE]7N.dGe=_Ob5?Je+e&5ZVZN6+@H=S+C(X
\bU04=KAeU9f1C_G(TB1;T?a-?4(ECXdER-FU_^0KV74HK<cU>1fYb&F+.&##bGD
82:LPQT\Gb#R))gcE.#3#@T-F_2P]a;J@:V#F)&5e)><eaaCb^556L_#BH7YRd>U
F(dK]4B2b]6O^e&dTbNC9FO.^W#MLJ7.RY\8??fLW8N-A64ZI\EZS;f4#:[CPNB:
gS2EP,66Q7IMa@MO(Ue8T[IU2(MP[fbD-/ATe&VEDJbTVX_J)4:gV.g@MD#DCc.b
\+PMP-6(#TY>E&,Ug_,CD=)E5H,Q7-B-NM4R4LKEb.P3P__<aTHL.@B?\CT]Idf_
D4<D@^\6,RBYH6T4D-X66^Xg)+bQ^JC<9[@eZ1_\RRR0GAQ:VbYTc]XNX^FCBTRK
5#+WZ]SF<YI85cZD@AKf\ge4&UH.O&2\_3J8&TNa6)7511V1dae1UEAK\CGBfeT0
QcUH&9[O3S6=WKL548NVDT>>PRJH;354.IVFQYI\IUW07#_A=A75B#YH_+<&e4Eg
BVC#N)^ABNA+]0BQ^,;.Z5+5J,R.[92F2\#cV^.70IRcM;d,H8.8;O+8U)/?_8fG
@<U7@<B<-3(?b)VYG7C#CTg<\bA=d14+S))5e0#\.27&XG>@0/MC1>_BT8Mg_8-+
ISU^XOU90a]J,39e8gc;IOG34g1.>e34EE2@@Ed;YVKHO3Pa8c/^_K<F0F\;]>NS
g.-2YcLG8K.FYV_)I)ggD#dQ^BK\#XUKGA2/OSe56[&DdFFU<IF)X3H:C>TEM/B]
MZ_d?)R5JW#?bZe5K^7/^^=X3VL+07)=8HI5Q<JGU+,,:I6LXK]a)QFD3,#bMIM[
/AHNUVO:5Cd-[>R>8XS6AMMZY20<@?NJ;OUCV0BdS&+JLUSgI5H0;MY0;?c;<0FB
e7EZ_IW@3B(I)H:\Y306F36d1G&SY@.P7JcBDZJDbYF.6WU&/X=Ia]QC&6/f2/W9
C@C00F]?:ca]\33CUW#0b+Z)Gbe2g4K<Aa4cRb6/He01H:V_NF6FgQEg+##<19I(
,CQ8^V3PN&PV(K]0JD^RU\F496GVW82G?e&M2].S(afZ4b.7-Za)JKM]S0G8+UZZ
?bPS_+dADQaFPRW26RI]GMZW1be.dIJ^g[;8Y8X?^3,S&+8KfJYVN&(X<ZEV,S/5
?J/30?X01+^H<IS;+RWI^-cNGCBCF30AK5I4S2-P>S[@d<]&OUe9cf\LOSWG[.<6
+<Q4H(CI)3>QQKIZWFG>K0RbC6gV,C\KH<>b=&_dca3/:I6/,#:eaZD=<6EHef5I
ZGd=a8d,EHab5e<BH\,P-Q,;O0]A&XPTOg7-c+KMC=W^FJTC1cBbEZW^4,YX//O5
FI;>c[T8OXO)W26eG=DaAW_3ecKT<[=0,Q<fWP.=_.F4#cUYOKd..MW5KORJB(\b
gP4;7J:CQ,17?L(YSH@K09F:UNV5D&fTf8.[,cX.\C8^9>]]K&R3aB;aT81<\6S9
_eGN+S;S6>.H))V3BNSGV4G<e6Ma0?RTYY^#TEMGJ.7UI3=SG?1Z(\_d\c<<ATQ:
CH8[-,2KTI\.dgI&da\^;]e:D4T_;^ZJAH3<<-@I_6\;9N.WKG21M(7N,,b;TW4T
&[;If.,9c5\B\<YE);DO=-bF6DJNH2)VeYZ@CPJ,D8H>]BTEGA<)cC[8J>6\X_N>
#FDL6cI;g,7FJ=;_4#^WX-7P7T@g&;JaC^KNOR=04(dAG67WW/?MVG3@&aT:+S[]
c6CB2>cJ0GDbV4;T;/c(aa;G8MgTF;c9P/4_,+8d57E6Pa<J\U[D-,V0@@HVD&gB
@L80;bM-&]QFUJIDM[N0g:HIRU9TX_CC\)J@NO>-@P_>)\9&W#[=5Cfa<XIT#8c=
aScg>V^0<2E)H_8/<X-N#@P^8b;Q.g:BE(NLE1Ld4WfM#A87d[[ZX6?.))VCgC\g
.aX+(C;#c)V_fX)X)_1R57[f41e6X05;X_0_P]WBa(H610=.Z[_X1NKeNAMFM6JN
@1D&b@F[]gXRDFG[BXGRUQf7+,?10ZX1Q^8/DUb6G75eYF3>C+])d#SA30VgYZHS
2LOZeR2YKX-V:S9bY48_L197;6EQ4?g0)b/(gSEXZ4UT&<841ET=J)DPC)<0L=0&
QOBAc9>6V4aEN7S#,AeKF4AaE&g90LCfB#cPLG<H,.KMK7_D0_O5Z_)]1B_aOW2)
]IbBf1/3bWI78O^9;G5]aFSAL2gO+W#D.0;4Le(<,4:e85AZf_1<2D8M.R@>(V1V
@&7Eef0E)C+Fbf9,8DM622IA5O[7FF[RT\[NeHBX_L2MHZ?0C?0/.B^Y<D=+U4GM
e3dF_;[a&<^Z.NJH3Ab;1CODCX>&WD8bN,VQ(gV177C/)NKW=CT2dA=e/99Tde])
0LF?.HEG.(aPceH=/WS]DP9L[\a>9./gU]M0NV+UMFP6N]\<e),6#d6Q.DO+aDg]
_?3UE;B:D^1LfGV8/9Q4RLe8Aa=UFSSV1ULAN,c7eG,A=2A]B[M[2?U<NGO_MY79
TNf^;c-^V@[M^/QM^fVRF^#>Md;V.&dJZ-1\Bd]9XGLO<+AUd5A-18c[2aZCC75e
,\&)].H8BQJ#/PJ6b9==]/5?F7L)RZ^6C@6\Jg/+ST73\-C]W\I0gSB_f.L;W\NC
Q)PX+6WI4CI#M=8bQGf64__fWa^fMU,f5<4Q)I.MGAZIP?BUgNcQ7E[J/g2?R\RI
N)EH^6dRBOIJV>-Vd&_:I8GgUg+#QF@,_2e?BU:SagbFa.@fc^KD983-/(JZ#F:3
1PJ(KUB:FP\#S,c^7b1K:1)+094=0]XA&MIS4PQd^M09;H&GS7eV()EB#C29KdgM
DHf8>cRGTUV_4a,0<ZDBLQ/L3_=\(Yd@K.ZCT8,CEXa1)Z+V#SfeO#E,M89<WW_@
6CC9H/>07B\TfE0J83\9HBc:G1AW1Q?5Q:.]Y:-A(T,+=>:NN?ZG<3Z@P@<X+FMR
SW\>8Nf/&XeH:/R:gO.Rge?<BB180&PO]CE/DKd]ZYfS,MR^/^9NTg=Og)gMQ#_(
5\d;,3cN,^T32f.(AK^@JO1_HZ#e1NT,SNL7HE8Q4J[Q;e\J@&(gW:^9GeN-c8c+
M+_AMBIL[&9Aa5N+F>;QBJYJK),J[=SURUb3H/W<9/<dWaQ-?1^CY6=>S6eT(e9a
)IIcgPW[^c(5@O=RK7E\7/.PPG[M=)]#A^K^#ZJF3^)A1>D\F2G-1YWX<b1;4)=8
c^+>G09)+1()J7X59N5+[A]JXWZHJ4D@N8E[FAgI-eHOO:dbAGIO@>ba_A2HZ+W)
bF?0Q+W;2<8CJ16[[@Y.B&>V6J\U6->:UB-9F<KZ+BY34b(gIcT3d>Ca^X9VMPJ.
GQMV6??eCYHS,H=g@Oc2c7NVZ&R/acJ>M;0^TF:3.U,O/+0HL8gWXV_+RG/:C.Bf
-+,,L^Y@15G28G3QK9J7K,dY^J;3T>EOC^PgE7(JYd4-^5)S\68+M7T\M<]P5S)W
eH]9)[Va.SB@YN-0^:/D>WX<>d)KYAZ:HL7+P[8UOef4e=cYJXKDbE2Q.\5R0S2P
g3ZJJN_>:D8/=&7=&.]IZR(_O8(O.=_H1SC\\OEXUaS#4K8FgYRb@2d&H(g@L7LG
5/;][F6CaYF5ZSOgg-X6+R3T+67_7OFZ0WM]>(BG9&R^\X0XLXU((f>34W10\#,/
b/MfZ>G^Ud/H<R9ZQYG9N_N<[((4Ge\f9bAg)eWVNf217D@:;KYS^_C17Z3\X>C7
/#?\QHON/L#W@M[dUYR34>S@#WI+LD:K+FPd,B)O&D-PZ.ceaGebf)>[L[WP,R=-
a^gU]J#]TO>;T@3NgY8(^+C?DgJ0/W,KF+f+_(:8<#A,^]FIe?FC6>d\0W-&766\
0,UAZe42)2V#@B/:HOK#L\f#V+E=>481JT(S=AI5HO[K498&&#=L5-1>dX.QN5IR
XPH]UO6.b=/4=5:MfR]U67a;RS/JXf;3]?RE)b,5gRDe]ec<2WL>3(\2/aZO]D]5
K=^BKCIY0Q=E3YCX^aA9Xg.+J=^?);D[<^2Q:R5Wd&>]g8Feg/2Ld0H\?Q8IWX-2
<=a51A1/-T3<C@AT/RS<Ag6-FLQFPP>c=bJW@U\4>aE>H&WEUEIPId]GcLY;^7YR
E;aTJC:N#V>]6<cR#NH3@F7W;+<WWCT);5V0.SYU_-#aIf_)<F&8?RS9@ZBH3cEW
=^5I3C&TgAdK8#CO,=7,C5IZb]KF#d:X..:I..\f]T27&BKgd&>7XSUS;@M.Xe(7
_&a^FZN/@X,F]/EZG\]D5F-d:VJGH.-GW806M[T_]eA>#^-ZI7OV>2_?GG)MeTbb
WN,7HNEP:FM@;T2W2O8)YK,fE<D3Je3Y8CSP_F@>&#CQgK]_3DBbOT)f;HSc<a_K
NSX<S67b_&AH&VGZI\f,8H0;Z8cE/L1@8(L@?]/U6a<\eTLNMBF;12>RQ__a3eE#
)^Ndaf(ZA[O<ODSLUD>@W&)ee7HGc,2KD?7O[UX-dETXP@S79CbV]d:/XTF<Z@I9
I[cZ:Ifb.O-=E>NC6KSK.N5Jd8U1f@@]&Y.47B<5;cELe]OaD?=bXG4=FG8#X8?A
;XAL/#8G@bEW?VFWNCG?5dHf,JGf:cRZ4cg2abHe34]NY-Z^Qa,JUJ?27S;A3@+]
Gac,HP:+aU9-@(O0PN0^81@?PN2RcRHGLJgI949[S9HbLU^)P_95]CCXQdG\U(55
39(]V,A22\IA@>f)bYB;PRKZ7<J]FHK24AN;dFTNE6)X[^FGg4(J;e,MFW?D+NWb
<ZY(Na,e:<XKFV2\_L#[dL<Q[e_G],bT<eCeI-E;^#cU3H]6QRYJQ8(Ta4<6YXgF
Y[O[ae?6_bbUXP]4^Z=P>c<=O<>ZPeT3JgV8^d2-bP&_EU##],)cEVA<5HFJ^NX(
;e@ZeS5Y9<Oe)e(\E/5dR[FTXWY0X8Q9]H,)M.5,TTJZC;9DF:de7/:[Kd_WO#3\
KEYN&dU8g.Y[EP,#;e48cJ>SCXa@-KA(cH>K[KW+TH3_R&EfB&g-:C_a)?7L0)0+
[Lb-+)LPJ7Z+2JRIM#FD@ZI_H7@X0^\-&[P.RAd<G3P7_R3</CR2eY;e.]VfIPH=
ZAE:2K@)I>&ZO>T<)d1\=1MNTg3>bD]Y<9,F9DWE]#]OfLCZ9PS01e_Bg;e>f<2+
XXK3[M.1dNDOBfTRHc-d7cO+P]5Y:g(QMA(,9,#NL;C@)1TRO];f:.8V\VLAEeYU
74Ra/JHc)8=+1,_e1H1_cM;S<8Q:d(gTb]P+XS;Yg#R_\(/K(/LC#UJ:I5;:6NTb
DB7G#&G#FN7<KD7&b,edC(&[aMGHI-<+&8[B3K3_IcEdZd14M-/@G;_?=G0JO6&e
MLSWMZ>a@bTI\[f?_OaR7958;8a(?bO)R-)LSOF4UX2Ea+7S+_#8L>M3MN:QQ_+K
0+B#=3Jg\gF(G^-M>_9((&7EDPfGY694@1HC9&e2?7I\4209R.QDV2:<4&#]W,#P
V-.<DRIUGN_0K\_5_JWL[Wde)[ePaNK-4aY;2OE80c5\P6c0(^(QHM<_9YfLZMF&
6&M[[DK#VD<FZ?3gOLQEa&IK3R3RV@:Ja.<C#1;H39[egWH9[a1)CaA\K)8Q@e&[
;BB7cE3E(>:&V@)H^N1CMZRNJV^C?ESK></9O3S7W;L_1\[((a\Q+-PGJ>/8JS@L
<2:>=/S-)POTFND>IMF2RT.>OYG(A=F\9\M-TPBN>?A-&Y7D3(Gf;W2R=-9I6R,[
>:IK_@fQAGf=IA=U8R60JY,R(&#b+6=</gE8b)=d.eScgdZaOgUc@_T2=/dI\6KI
g<\Jc,6W6UVdNX^4DKRf&5H4<,IH[LY]f?1aIVfXDB-7J.b;^Y\+<]1PMY4O[W_g
KXUcW4[gCeY_5ADaBJea@C+XE.HOBb4:Ve]gE[\K69XGXXBa5QG2:6ADZR0].(C_
Z<gP0JUgb6)E<+HHCZ@]0+=IZM(48CGcR=VZ88TLB0H)1[6R]C)XWVEWfSBNcg/b
R_H4<N>GJA9NWO]Ba<Y+c&aA\K5cR\/Q/:?[[J6LFS/e3RO&gVN#3K[R+aV/D9Td
:7WXAb&2b_,M_G<VH_A12?M>Te-H#02P6H-@3e6Fd,f[MbL9TR&#-3c)ZYgFL@N(
5)bX#LIRHECQET.eGCHbJIK0J898Q\&EFeA6D+YT[5O\[MM>gMMf<SFU=U;=E4OG
DW7G@BgTfVF+NIHBVKR\<)#db,]677\O?W7.WXE=Y#>,97.OXYKKW\f(PCTFS23V
WV+VL&[MFSaa3FE\8_-9Y:55VX4X<QLc<7)X[GaMJg-F4f?@IM(L)79bN[RXOUU2
e#ACA5V5@K=J-2>@37F[^a=US:_E[b_0UA-L?[:2=C9bc9\G[UJM(M5O5SM.>N,Y
(J2aX(X.#13AT0M5IT89RV;/=GR=X&(.J^UX,Z8\1eeBV?T.=-c@[SJG;d+b]CQS
BZd[/H+JLDcJ6/;)>3ScLD\SFQK7Kce3<9#5F]Y_V.,5[YB)@T::BfEX:TR<^Q+@
Pd0P.bM^\6\S<Sa]]O>1,2FZUBY1Z+JO_0&HFQME]5E^MO^LM:2+Z=4:?U5CD4Fe
N]aT:daO>4^Z;Z;-b-V6Q+50A<R)QL?b-FQ0.WO]^Va(_6O14Kc,CZ1AJ63KMGJO
M9ZBDLL7d3OF/M6/7GHZG3P)-bJQ+KS?Xg4;>7_N1TPb2b&g9Z(CW7JG[2KRMdU0
LV,+DX.C&]Eb=ef?ICYB=D];^L)6):fc0:Xa\_Q8dVA1EGg-e<d0>2QD@WVAT1V,
b.EDQ]3_e2DG[N/\&CS>Ug487D-DK&YfZ9X+.,,#.N;L:?/?W5aV)HJ&S;LWCJ,)
_,T,WN8DP-^HDJ33[#_BB<NTQ/4#K-M\?MLS?d8#T#QX:JCU8:3?-8YB^BWc79@;
@9?[N<)R#aDDLHc#HAg>CLK?2b:#5D/_,S^T6d\UDe)L1@R3)CR::/cc@P6-4SV-
gM7fD.9OI4KcE<E5eY9:Y0/6W)XWKe.R,f2Gae66#g?ZPD+;RRIHZSG<(^bK5:LB
(+(CH0G=1TGQA\_[BU]G.(gY_,@8(RU<ZC)4#L/P[.B>.GfX6ATHG4d>?LcYe5R^
Ze)PgNP@4NNQ+66[X8?Z1&2Pb/+O>R7F<.-?bG:8VZ=,)2eH1Hgc-2JCRJ&9U\gU
\R4[J33/N[:8/K_C4C+:UeLC_@,64CbGeKJ)g=(,PG_<:/E8fG0)U3;#f;)/I3KL
J2\]gIQ_5J+<M3MQ#-]Ub8?aS<]U^4;K\?X6KS<e&FVQg-5K#_<]M1#Q_SCVJ1f,
61UJZW,eNcTCKJ>GBD?^H9_1RK<@^TSGF^Ag&]68VS\\@fb(c;WbWd(1Q^RO?N8T
6<,]W44a/WfAOC^^KGER?RSE4fQB6V,[@F5_9ICcRYY1KX^+V7)gCP\JD71V&O17
aJ=GUO_I1>A#_@CSFUQ]9S&U6[2C>c-N4QQ.\J[OG+adZ[B(T^(g.c7-IV-BJPUV
b_d8X,d6XR/=Mf(Uc?#)H9<+_=cIH#PebI>YL2=X^YB;^C1Y[^.IJIB@O#H7DK4U
<.7c#0([4C6CI)g3Q6ga]=31[SGf&:ZT2\+(^d+(,=;5&c#e:X1g9K8&)X&.,fQ^
c(Q^JgL/<1ec]1QUO=-c-G3@KFDOE]0DaYD1H9W))d0HZQMff\Lg2-NE0-5aIIYZ
Wf:[T]IANe[B&=g4);_>/97\=-^Q@+YeQM5J>X3[/WRQ]@]Z_,VZIT7.B>U5V),=
/TDQ5AF+GZ-)bA3Z/&APbO@QX4<MWeCPcVJZ,@JD/Z>>HE)MD9-W<EB4-0ACT\Le
K_76d>2S:@CRGE5cXGQG5X#_K/@,P_-d&NK&55\;.JF6TF5/^b/<FW;.;8GI+NRH
FHa<#]d?B32ET+SSJ]D;Nad=Q9E0F<KC2fa@5YK?>X=b<S_1QYHf:ZE-)2-<dc.4
d.ege^Q/UZc\b_RNW2SQ0=2V>J;F\43T(QVc@[S.WGF[gVC\-b5([0D.1fa60J^8
F)4Z9a7LB4MR;[P^>QbO+<-.dU<78g25YCYQNG&@CNI:FHEZXL\b,PFU5D<&A@a]
JM@_B_CXQ]98:_TMHT3<N<R6OT?L<VICbcF4?DV\+F)Y;\JN\IP091,W>)I38&P>
D&^CcgHcZ\CK_-YX[[\YZ.&#7V7<##/(Ke+[Z\6Ud[>&1OA?NdA7Ae^\CCLaeOSV
0L#3eTg>=;I674N&Y[>,#?I]XU[8fVI-I#&6?ge=[@cIXNV5X3/MP^R(4A#Z\X?8
^3Ve[,&=0d)^&#KB4<H[K:5U/A&/\?a6F.8(Z&DW[gXa>U\]ZJ,Z#ge=a->4bQ,L
WA8KH5bG8,cb<\gFg=8\:O6)@eT6<)c/9/1].-Q##IBHa\TYdL:C+.IL@BCUeU6;
=S5gYS0fdXRgDdRA1V5R9X[f/dgU?F4ScZPcSZ3;#@HAM]TE@3AIC(/Q+T+Y\W81
,NbZc===(b34&99HLg-T39)L,D>X@P^TJ0bd6\H,7@OZ_5Ne&C&78^fNX&?E(HO0
#Qd(5:HK89-ECOC3BT=BfG<B\8\]QO&)(Ka9fI,dL)D=YK\ADY@8f8:1BNFCJ4N/
.;U=cM@YbD]#NRg.Eb,QU/D3G8Y/+R4a=4KH=00UBA,>1ZA6T_K3>3:CLT0#5@Ye
_5V/=C:d15E?7:Wf8H;K0N3-24SKO>aMXc<]IH4H-cWHJ&1]E^5/C;B9Y3_5ZKG8
D?<8VR#/NQ^6(SQZU-N:ee;,-OH-@OB,QP6ATK8I-SO:+Iea0#<@NF\3F(RV+BaU
+e&W;3O[6gG):^OA@.&3B9<Je-R9.?(4P>4?PJ[K_51WL:M>gSI(c7e=VIM7#(@L
J8#[TKAPQP)#CU,7.WVQ=#CI(RISGb\;FFf,)E7Wd<cNYLVHbVYU+S:Fb1O<;PMK
+7eXa,I(0^YS6;FSG(X0N0E7debea+c)C2;?=X&d_79INfI)3@BTJV]MNO?9:?2I
S0EZPEaOMQW/C+5I05UT7@;9Qd):gC-O/8Ga?#=GM\BOAGD&H#CDALVXFW(LeF5C
IP6JA3>G9E6-?Y>/YT+,/IHN3_b=N2UJ[6b?K_3/RHL^_cEQ2\UDT5,Z7KedceaS
O-K4MFF_8Y<OM)<bP3<P0TW_](G(IQRbPIJ0\\>NEf]H9L71_E18AW\69bI78:=3
BW9W,9GNE\.]FgIfO6ZIE:JU#f[B?I9#/#AD;/dFLKg^=;dFD(>g[8P.K8&b]=da
NCN5c@:NY8E=KWC;>^WEUdH6H7H/P7fPL8dBD9VCRaA/<;#,aa1K#d\=WWLKXSJe
aB6:O_)(=\(JDA)-@+MLMbA\gL>I7/c9MHG829\[KeYfaU=^FT;JR9H]?dXA=<)R
eR_)R9\9]_JdVWdX6?:R2#.7\a2#?9K#<35]TBb\Ef>31e3ABAGbR?/RXY&:B4Y0
?.&Raf(G4V&QI3bI5B.f29K_AZ+ZJ:+646U3<P&RY1M7YbF1\d>VVU.+e_e_,fX2
VN[^0^g=\UB]=O[JOZ9d@71@R:QPbFAfOF8YTL0=/I_Sf83U(ZEVN^U3@b-L@OEB
5&6^0gUe:KCAKYaNIU/a1#fAK.Bgd^d\DcCR-e/YO-^9^1NAf6(PNaDBYWJN.Hd(
_=^\UgM]7SLL10.D@<.,B\c?3N8GOJ#J]9IY:Ie^&8BK5\S;#OLY/=7P2OQ@VN8)
+\UgR0IM_T;CM7PY@ee6M#@^D:[SG]TG:QKI=XH7NIcBH8)#R:=G6Od#&<6+7<MN
^A,.GBJHA2HI0B@8S7F0<gA(fQ&cAceCQ=bQ/R1LF0<b<@69]fUODL/Z.dXPegEY
cJ2Taf_g,;AJJZ3.VN1<7d@^(Ya?^BV<4[3#2OYTFf/3Q;;QbWe/TIa)Y,89&;]d
BcEe/B>6b?3;N(K<7R=,?ZeS4Se4-+_C.R9aXc63AM2X1/(ACAUE(IV5K(WE@(7W
(N0L<C+C_F1S.,IK<N;YC;\EQO3[FL5XeR[0TXGdNPYT5@b2^4ZNEbNJ>4=d-N;:
+7P/[2(,:gK?e^cSM19XEG]8XGb(&,:MGGa>8ITK6,b^BB@aR7gZ,4fF<:c)KVIf
+<[UW&3B7\V#]9?XIIaDH3afAO#G3YS2?P#&ca(C+FI?f?PQe[EcXc7W(JR#4OME
7-S_d,5R3C&gZXfaIG?IJFcX:0@>_9G6CILUe0b726d<<a/8L@]0#e\JYdLMV>5]
BS6>E4Yd1]#AHIaBJ>X@,II>3b/&3cdB^McK=b7?;2:;0ZD>aHV[\.;AQ#JL=4:5
W=211RQ0cJ0b3c\KQY-c5+9Nb->f8\67WZGGeO@VGMZ1:]_KO_B5S8<=^ZgLB@WB
?7(FK1#3g8<85.K>.bTFL[/#88#0+e(Td=9bQ9^W[/Z1F?2>gAOKV4)GR\bG?#11
1.^?C]&A:KDNeT8YPa7BAY6DdFQReW-.gY&EG?g@L2WV.A\:7=RQ[8]8ILDMIYFC
LX8U0U(_:X6MU9[IZT8JbT=_b@A3QP5IG1-7gc?=/D)WRF4W&K):eAZd3<\g?Z1B
f?c<a^0&\NgAK:#2=<;M+16,2NXUR]g6X3II&A#4CZO1.?:11F(SgN_HMQ8McM68
VB.GTJL#MF;V(b3&,5]JDGGV&=bC(8-MMAND>I6W4b+^a]bdF3e4Q01ICJaF.OV5
I0RH3WFfHF<V^[V-)Q+cSWKIY18MTRS1J;)a.5K:RWWC[5(9I7(UZYd\)N:[bID.
\&7fNF2M=PD-GKPg66LV3YJYSFB&CXa<R;45,T=S-#bW+97[#)?B@_B&-Q^d5aY:
FMT9C?M;:bYV#65+dHLJ]F4/cOYJ&:&SV0H8dJP(;J^F8NN?)/7;dXT6]3]M9Q=W
W+-^I+2[U-cHA>42@WGgUeS4@A1H&FeKV)(dUKZ5NO6L32Kda8)D?ZO03X]4Z[f?
+F1IYFZKN/]3A\1J\=J.Hg4^Z_NK,<b9d:Cfab6Cg4_;R?F)G8E39]DNW+K61BeE
?b1\K0ZKK-\d:_Q<<I]R4OU4SN)^#Fd+51M<.[Md^=ALA[JT5\QH>4=C,^9d<8B6
gLKA(Z6AQ&\XH<I^#gGbF=]Y@.I9/[)R7W#F=X11d.9CO98Sb55=JK#HWD]GSeO+
+V?G.[fG_,6Q@AId;>X&eC<JGY(SGHRc&WNQcUe&V]]7BY4^45/X?fX_IIfKH]8_
U1KVbU(\+UY,;-;)b]=CIS]C\/],6L/DE@/WbJ,#REGf-LcC-8:,EFV5\8_bX\/O
3&bV3L5@15gRLSeA#?G\+M^<D4[GV/9Df&-(FbPQZ]RDbS1W3/?e5b+C_97_UaQW
=]S.CL3=,O5PCS[TG&VT>a_62QCQYGLVNF(H>[E+V(:E54D>SJbC@:PRHMA>16A>
DI@9^F,A]f2U[Ua/1NN2bdf(UYOag2]:&Y@QSTD7F^)?M+SMeK/ES/K>GSBJ,7A]
FU>d_LQU7\X:UQM,4D1S2AEPZSgG^7\\M,d&8L>4X/HeU?3YV;]GKa_Z\INE^Z<)
(,U^Hg;;:6)0+UQ=KV6/EaX9H6g3XTTBQ+G1+Z\K5H+85O,eWZBLP]<e<K?CXJ40
g<@HNQ&0cYH>GPA.Q/SKFLTYRU>;4[Pd)Mf<;eC+61PcY_bdNKZM\Icd?TL(UbN.
F-TO3g6>;83GG5YC#Y.Y1gJ.@?R]PD7C0=9=^F2fUBV2@#W9)N:SYV9N;4]/KNPN
FQg=A,[bcG9@dF9fXg6,JfJ1:O-)OO\^bP0<S#@fG1VH_NgW>X0[CJJXT-eRAZgT
fX)J5FMYT+LgZ-NIcOW/HN;00OO+5;eRUe<=U(5bHSYD/VaK\6Q\>V0SR5YJH)e8
V<LN]]EE44K<0<e8E&&SM557Q:(#MJ95Wf\EZM+1@3#=<c8J(RPUR;NNCU_1@Q+a
_-@AJ.PL=+]_(:e;AQ>4WZB:e_;RC?)UMU>/:7V9T?SM?CYa_9TOU<eCbEcMYf;L
_HJ-WIa;:GF_>@AO@bRYNaa2Y@/K+(,,gPf)(e]c\O?1:JYe_A@HMQ8P@=[:+&P2
e1A#221.R53eAgNO&V.-)[[&T]KT8YS==9F,]?,Y=Ua.+aPcY]K@\#HILaYa9M0D
gFNO+=OIV#2dB88><^Q_7J,A0A=\gbfM68UQ>:2N=S#47[+FK#M,Xe=O@&4^T):L
HVMfZ.U73B.[\fU177G75[PKH>?.dC0;]^7L(5gFaN<^f/gZcFE,4[^B>f>JcJ;7
B\/NN3f6g/7LS5CJGZUF=7NHO9E>WN7VgcPJ2;SV\@RT,Yd@_IK5:@VPgG^S(:JN
g(FdeFWK[H<JT9cAfFJb>SO]OeURSLFLK?WMTSR9^6)YB=>.\R7a_WAcdE<;dPcX
[)0OWX=#F@JZ(E,-I:OcbT?^K.fR?e#?Y5NK89)&[UC1fO#>XS?4NNWH9K9+4a)\
&\bAZ+1W8RL==d;J6b?.Y:M1fPFMU-Kb@E-N&.cg15_dcF+Z[OZaa^CGWc_O5UC&
U,_AQE7LY?14>86.XIBOf+O3d:,#L=Kb4fe:6AZH7&?RE7U-=27/JU_FEec)(IcA
g+T(JDf2[A2e^.J?:PY)OKJFKJ<)4]@f/KEC^V(WQI#/+Ue)+F>;S,M9,);47./f
Nb\,I/+X5AS^0gNI+G=5O-._>GCP-A6Ac3PZgN8&Tc-OROdQfB]d_AB/M1XW>M:G
XG7OYN0V)4>FX^E9M/8&ZQTNRLOF>U57f&^5WHg<@VeL)eg9.EaddC9R<>(:I7.J
?1FY1O-.F)F<b48/9U5X?&0IMUFQHR1.e+:6-S;gY6\S\[HV-YC_SRX+cbg>aQ^J
FD=X@3P@/T;WR[g\VSVa_T_FIM:B7+_dbUP&4H2e=D3ZK?D,e@9UIdDY]0UFGH<0
^bT7aL#RI:/GY2KFPb@LRFB/O^>W4P^BX\dA)UV>Za(-HO#7?9L&fcF12>Tc^,MU
[7E8^ab2a.CZ^MI2ADRG[>21a9>AH)0\NOW?GN\&[6caC;]-W_:5K\g0-8>\;W[_
X0]1c7^O;+QA&DY4PZ-d76/;+[\J80^&FPE0MNN_bCcgB.@MX=d/?B,>K/6)[GE6
Q&1.+2FERUZ?faQ<C./>Q9:0C1NU5LW_B9^:^7R<N6X]MFF[HVX7_+&(=a_75,>B
?NLLTFT.>K9MWRZKKVH,)JT0K4f1=1af.G[;::XZ,_O.O6>DgXFgK;;]+67d8?3A
X^JX((VaB&c+3T/LG7A_A+I(I\:RLM3JV\2E2@\6B>T0>.):QN^gDeBZVG)&JcD;
[+>9A^6JB3_cfd+XCV0176VE:6I?0;7=8ZPU)SZTQ449U@G_VcX)8X.ATb)K]ReQ
REIBdMFFP)+C<>C0@eB804DYF>I\/,@X@,#0=edg8cI:C9b4XG[.caZA8EE^K+[>
H-aeYZ>9MC]gJ[]T4Y6C:/b8f89P4+e^)K;@,W<gM2/L7,aB,OaXI-\^;&@2e4NC
Z<1C.0Z^5A0D2NaQY)WT72-8Q-]M28_I/0W[U<.gaB/=_g>MD3VWYLMKbCWJK\C1
4+Z>>7+ONEEYT41,R9&=.=SRN:QM;4I[BK77T@#:0^S:7(S5c85FY)[G[.:<]=-E
2#>D1cMb9@SYESH]AGPW;1Gb^3BAS=^R((X_J>MB;4Kbg7K@91J?P0IV\Ab.=PZW
9^&b+<:RFU[_LSbga>6,H]EAX89)O-J(]bY)N1<1WS)VM)7:b9263,]V,CI6C88/
8@874>:H032)c-d<Z;1,L/?1)/J\>CH+H#0TGbYTS,T^P?G-4?)__U]Hec+RP,/3
H=DWV8b03.1)?NOSBWJYV9#L/b>S<f<OM5N\G[#gU_PV\.FZYUC6\+]7?\H[QAZ=
4-G+:Q=<0+(AA#c2AU_:RD[[c-:5E0)DY91V&\S+B^W+<69HSf>UB&T9482?J.8G
O:Ec3dJS\U;NHb_e&,#H>D?1KVLEZW:7C&0Tf^EdO1e[_>dQ5e4[,64L7-gP7F/O
TBQ_X/73NV?UNe(O]6WDLM2H)F_YMB9dZ7T\=UbGN2D+a9cHEfQB6eC420^d.JO#
T;M#/R:.W-HgV0LCFZ_cJR[&&YZQ)43fU>T9eRFaFK.3I]@g?EbTIB-T55PQUOfA
(AAbT8:cI>M<g=/;2E6><2+2I54F+e,HB#;2=gYFH^@XQ8>&KaVZ908H3IC0L0ea
/QOY?ITSJ?/AZfb7.eA,bS9CZ3GS8ZZV/7),?1(=K#;.)8Y-8A/9_O>JfW3L+[WZ
UU[:W6_;]A@3XLI&d0DHR@6A0/U8Q5\f#NefDgI:WWVG.KYL^9Q=MFLA)99S:2DP
?5L79fDX88&H.Z,.V9XQb3b,^ZcNC&EN3.-PK\=E3NTY9@Sg0@5,VM[F]>(Ng.CO
S9e=R3;:.&C\=Xg5J?5-g[MK&,^,=W?2Xd4Xe@(74Y^J[+<:<VJ<DC-XgdSUR.gN
,RK4:6I9ET(_fA#?67S<_TOH+:;3=CdYFW<@PG-.S2=@HZ;QgH<7d]D7dNH/IZ[g
)D&H=@b0-N\QZSIW-P\e=7FWHeAa7b(10RSWOa5^C(,Q=;N^,\\RaM1.]<8U^F-^
4,#ECbJHG^Qb663):Y^&U>(f/:&4eWMa6S,A\f7L(0]G8JI?a5,^V.XH+6+\DTB1
(LX7O&b98Dc9#Rbe8dB?D.10Pe1)(4-gYCTBU),?K]R-@Z1aJgb]YeTXa59J4O.U
;FU)<YN&:(>W?S2,D:g:ENE_FMeWX.cfMbB+]/L15Wf@1IC1Y[D-)g5LB)Y.PE&W
M2)70)E)6U#_Z;RW0P_IO_+S&7a[()DE&1ZY>(4;IF&+>eCZ+9^\KM671OVJgU#<
5QC^XIM9Z11a@S7:4-:7[W1;_5YE_fg>WBQH7a[4D7[[0#URSYCNM?\.X[g.;)a&
86ca(2TFQ0@+IN01)SWX>f)5-5bX^\WbR^68aQ:SZeL?@\YLZK-(:;,]P)1U1aK/
LK=FWbE_PF>QAHTg3fd0#/;BH1FE3D6XL&UX>gB)IFL(QDdRA+I>#,.),U;[E4b4
aWAL,JL8#U8IT?#[Z5V&[6-<=(SN@Z]/eJUPJ.Le&A2+WW59)Gad/7<@eH9SZK5Y
.2Y,dR:G-V+bAe?2a627eJZR9KM(#1-,e@DZUPfFf:(>GER\)B+E;a:b9c63[+eV
?NL2HTU^AXXP0(1GBF5c4]OeL<(B;(85J]^>:>eX/G==M5/(3(dG84_0JYf-4:dB
c/#;OR+X4]2N@I#KZE?V]90:gZL4ZAb^+VK1A2#b1M-(g&-6;gO&(]LUbOVQc<YT
T>;,J=2CURU5,H]1+7^J&A<K;CE\9e?5H:5K^SAXX@IT3ZM^6I=9DEVbbaBC+OA@
[[X=aVB.EYNb90cHV#(EP]#?^^=3Oe(MNDfZI\C-HD>V1,C80V#HEE#3(eDg7OL+
E6#S=WP>Oa^c]PP+D^^01T383A]<R#I>?G68_:-I#Hd1](7g0#,)B>)W&.fFN5eP
+eBe\f_@59;?BLHd]G]51_3?OSJ(#O#eK@3;BK)a/LFb;M+eIg+XLLQe(?L<#-9c
,=#1.d-b@BOGN<+^0^PT405b=E7a=4(,=XYCHJbB5A[\9YU+JD?fVEP(2E13WfP^
=ab+RXL=b_bW8_C2(;EH1PKSc?@YUS/fBMc.-E;34cbTAY(C2#A,Q:16#5DROMRJ
;:d0&a@_O.@VR&MOCB[1^T3RWBMDY)>FTbG@cR^IH-/:GL0)2<02AcDF]GI[,CL\
)/0Q>\&KV?f/NUJ0Q52&^EVSO;H0S@(/7L-M01A;I6Q:PRY0RPV,cZOPd:-d9/#O
G1=Pa>3+DS-W6(9@(2U7V5)KW+b]c^L),1P?&9P9<G/5JBK<)MeO[\X\SW9/GR<6
(F9Q&:R7\L_7<6LUP=2RJZd&)J<9UHfFW&5&Y];cT0aVL3eL7b/V9>fJ:-H9&DNG
J[fJGN2R3f:HR-+K]\2&HZVHV?7@HNQ+3Y3@+2Fdd&eM,RccMWddfQ;Q18eES]1@
GeU]X[=EL=<b5B@(^\\]JLE/5V)-YV;E-2)0L69#<]-S]abcG=MCgDS-)LWfU&1:
bE4MZW)SbE@#IbF\JLX5bP6Fg_F::4B\7CC5/?,H6UQC59<C9HJ/SaO]6+C-1H(7
.OQ:+NY\I;#S_QP+Q(-7)KEEZRX\VG^GD1TV/#[?BBF.YXaX?X/5&-g#1J[\Y&]X
I-Z3<27eT:YX.^Q<41EYNW[T@f^Q/M=g]5R#2QFS#KP^ZXR\1d0Ef2aV3AGHH5,9
=HXXR<9D?@SYB7,C>6BX88Nc7[bU/._9D0#_V6FT_]V&4LJ^f_eMXf[7D9-8gg9c
7ebM5gT4<OH^c,&g<F.N;T=Gg[FG.4f-fXR_R4McdMe60I]Pe81X\^]A@RS<WJK-
O7=D+HB0dRA/6cLa7dBUa-X#2H4OMeI^\Eg2B[O,-]\N\\Oa(7fdJ5BZQ==3#f^H
V>JWBEH)\MdWK_4;[,6&M_1Qc&&a)MB]0M0<&g-A^VaW-#6-9(=<M0.D2KIb0c/&
TQ]@-LFde0NDb^VY0[L>c/J(N<K4XbOPQR7\FIcJ@?:LdL9246eFZ0VT:Z3f#C;@
2-VTU:54eV)/NV8O4WV_#FJXPQB9^C8^7fL:DVL)7[LF?D3_V2H:N/M)\I(?9f^V
IT&GPN<GIgYAWb:;^K^AK(X[.N0QO8a\C_Z[<7R(HIc^E(D8S0UL_R7eCc@3LIP[
MUPL@87DG3[2XD_2XQHPEAfbEW\TY+ZJBCf4?-dc9H@g(KYG]-;NN8K97>DS\>_f
J->/Q261eg.R_T;^f64?^c)7P./B#Ae5+_],942):9K&fOVUc>\b5@?6aTc-3FMJ
8K6(HS-g2Z&D</6-)Xc32@K)06-MI1F?0+6-B78SdEAZ;120:]TYcG1La_H],GD5
#2Y.GX?L[W;>IL+4dHHfe+ba2caCN\&:[U+DRGe7()_;RVA&ZA+E#C_CR(=]eF)F
f7FP2WFJVH;/,#)9LA_MGGF\/c3A>c8dKF)19f#e3F_.I[be#KK(b)_ZF)7a@\(A
=-]X[3.2d2[M/H/SVS&(Sd^2,)0BXK#O9.U>2798\9U_NbQ3-B;F#g0:Ac7H=2S,
3AJF7GO:?/96H+;P8]5T4A8./Sf;<?O1-;Z#>_D</_WTH<T#b4IKI<4C[Q3N,^]C
Z3^dW4Tbc1(:d<+#aXVT9])ZfNKaG?J5QMO&MT.I0YM#BDKKg.4W<?Wb=D7@SOM6
Xf8C+AB&D&6)fTCU6g@KI@0A=]a9^3d3Rg<bb_Ca]dS@]M2V8Q[aO?;2\F(><OXW
[N8)#_9C,+:ETI6PVSGM]/=^c/Q[O#[)]Ve8:54N[J?\L@]aI[)DB9QRK4KU;N\-
&I/g?-5=<29(8&_P?&U688WX<M2.7S<Q\cF#XLCeW8R2YZ+HJS73O@NQJO)W,VdD
UNc\I+BM\R]F:HIF7I7[]e\AaB+N>IdL8d9JI5.P</,;I_9-?Of\4>Z9Kc6/..EY
:=?-)IcMW0@9C2V/Y#fb.6.>+bR#8-6b7IHR+.[XGW&>_=bLac=\E^/B/I;^df=&
0@A9NRB5X/Qb)YKE+,F&d6(e[9\?AJV[BNXf.Mf[UA:TZ>_YEJg=;3KG0K;\+QBb
5PU\;:-<&CC6C)_PK8N67#6WTEdP?5[]#,ZD5Sd:WB/FU)H?#P[X>0&D(<R[4.+U
59K58g7B72<JVJD42,B;b)+^LY?9CP/d\@E867Y=A/=8a=[+WB/d,[W5Z#DL2@R6
<TNIKGM1ed]1bHD[:bgN1A(9N@^cL)aZa2F<LU0S=LF<4ad_9)b[QC#A3<fdG>Ed
_@^4J13fYQ5QY&XL9.GH[I&b)H^cDQBV&A;c.&g]PSH9YR_&=/de6<5TAUDHC<;7
D=0d&&]MH<KDX]_ZR;IgS.-ad,FgcB&IEQOVYR/RI4BB5CQX)3+eI=>OQg1QR;4H
8?]@\7F3T3O_Y]g9=YJY.M3B,g(;##,^G;<P_UdDX1^#0:8\V=)0FMEc)=?&gB[-
S4I@YVCE+AJb)&g2\FO,JJUH\IO4\XGdIJEH-6XAa]E<(=P7+EV<3A6a,HI_R:T_
A6B@SVN8GY?V40K;a3OJ]Ae=eS/JdMFZKg54V0.)6L?d[AXB02&4GQ5L:84]Z&#?
A@+T_1>e8938,A)B=7D/11NM;/)N7b4;f-L:U5@K&5?BGD2R0\^+^gOT>+S\c<-;
&1f(f(bG0LD);-7KG,?5AF7YQg=W3P0R:4K?YD\V2?IP1>;W@YR3W077e^29IZ5+
8@2CI5\4a=U?H,?10R4g6]5bQ<(?=@4&T^]<bM<V1_F8<.gUV#CV.Z7A8gTQ)HX+
S:=9:B:BM\GcHa1-&J-Ve=T/[^@D[Hb)O:G]LWX99NaYS4E@b=J#YfUKHGPR#Y4a
(QNH8T8G)U[Q0a=X2J)L;+NPBJgG@g?+1GZEVOKGIb8<(,]9[W=5R\0PJA9D>>/_
>))b&X->[N)9C\>\GLW4+04\>6M(PJEPafYdW(&Ge,dFR8SIMQ6aE6OcD:ZXZ/H#
CM.DW3bFWS^,,+;A>d(<S02,AgR/TUFXW^S9+D);5dNaVWA=eMKX.NEHL?#Z&&Od
=,,82<#0f.]\,,K>3SQ]5U()B3/HdKCX_[3cY40O,.J1L)aKX3X.M,Z8cX8NSgDW
D#Q3,R>8JAK(.UMR.8E4X:_(;1VKL_IM>6aMUS4UOOKdWW_J9CH-85ND_@_NZ^N:
TP\2_)GL]CN2P8-TCX;:GbJa55@VIOR=bUTaF1>UUESM^?DeZ:Mc#CJ9A46=)b1/
+ZKVI9J5:UHGNd_F@e8/9\>EC)J^H@TOM].&&F@FFa3?@)S/NK2+a^GPF7A[>#7K
SJ..>ag=?_>MWDG/abP]FQdRKF9I_f4T<;TFE[+Yc29E+W4:+6;]Jb^cE/?>CM-C
B5T.5cfJL0TP)EI>V;bU//[13;K_8OKHdYIMP,#A&eN(TccGUA/YSV-ET;f+\P6@
[M66\\U:C#c]^.:M=Je=KSU(([a43LJ87HQ^=]M#&c/7fRac6e0VSce;H0[-H#Ud
g8(WHC^[C2.C&5O^]HfS^5UE;GL(?+R@eYP-\JKFW@bR,G7D7G-Q?Ra2Ec_B1IZF
Ne_0-QQXZ#PF7TN_bILaIL0//f0EXe3G1fd548N/2H\M;4ZMJ[K-Kb;g#@WWG.d]
AU=fCfU5RRK\O)I^=[eNX7?c<CXWG#VB/RMZO2fZ81PT9LFeZaOR+?;Ya7<7/@I]
MKV?NOCYEO((2JMH+?QW^9X<^7(LBWKC&Y1+9?/6BJ&b)J<DR+N&dK&ZGA43aFYX
F[90_NV?N)6);N1Q:\b]a-.?MV23,UW91OCXRS9(Z]IQ<8Nc>-N-&c:BAC==ED]e
CKS]O7;)Kec0;8A-FH6b;QF+<MY:MWI3MQ&OG+F=..\#XgZ=2Z3f1?2;:=ENg,K:
N3H,72P:gYcQ9C09MH-LPIX=OJL9^;(?,Oa)Z<=&4+F?B?1IU=A[c?c8G0#@A:]6
d9INbNc8DH,\&4_-EG:d7cF+RNdW=>e>=.=,]/\QH,AQ:(-f45J+9YMULOSAX0&D
e@aT)-_=CPaDb2D6DI[P,fMI;OJS3Rf&U^-HJTC1;b2GI8\P>XL.;#8E:]JRaW([
&_@C[60N(S@HVXOeK1UMXB#c+E0cRc3#=Ge[2X?N[CSU&3R,Reeb_5;Ug3_4Y#@3
]EVY?R-+5\TVc<J/46]B:,<OQ)@67/DTO_dX9DDN(29bATH@-dVOf:TP5:J-.W\(
;JQ330GJICNZB6#M2J]T8Ve746BR#[GAe5F#WE7eR^&/_7G(W,?^W:2WJb602.+7
JfIT&U[J^c&?a#g#.L9W36SaLZF,C18a;DHT;;,4&.Af:3&T?Id0KT5(HcVI5?d:
@UeX1_e<be;aLS1JbY0N2.[S_IO7#D6>D40PXcY;DPLf]+P<BDF2@QM>a?)A8R#f
?X8ZLXB#Q>T&U7-JdR-egNT+_=\b@MEddR6aVK,b-=&Fe69WKS@3?2XIbQ;YM6-5
.X3OMPXd,D6J;]0.&<6K.1c9M2C7aS@=[<<3V+I9_IC-FZ+MPB=>TK\M@E_;@e0e
[ZK+#IGCPg/^?DJ716&QTCGAC1f.?g&(71BY?g<9/cD&I7A0B-,]I;Me.VQ3Td3@
@X/d8PdFfg<2C-MB4\Y?+O0WE+e&,&>P?H-O9S^?5J<<Z.05JL_)SJa8A>PN(>B4
7gOIOb5S9;^0e<G/M&:A7I?0)+TFQD?]CD]8R1+9AMVED\ZV](a7@\CJ(UbbWYCb
.f)O-\M\Da#PB>I)PO5e/>@U+?AUa\(+QM82JFU,a<M#^BaD]\BNaAff3SNNTGW9
6?eM72)G?M:(MW.2bgaN/MZ@U-@6^E,ADOCf5\JF;6d9<<]fST8PSH:aA:EfTGIN
]P0Wc3g)I:9dd>I9>:QP=>ZS?^AQE69GQfPQ,M<GH,_3J(]T=[TgMBL;W_1]O7WZ
-OcUEU26e4B-fbG^5^dDgaXZ;BH_IK8<L2g/0bf>^dEC@KQNSF(M_(K/FW<2O+>F
S(c[\GG6PFYF+P?gEbf,L2/UQJ=+X_=^+Ma(^B7BbSV+>GA]2fX.]UM/\GU,?X?K
K=-A:9U#D=[EIb?;),\M<cCY5XdCRUX:0\S.[&@fWDdS-cW8/<\?HWO=<]WIg5(a
R6IUSc#cDTN9(+62+)cdP=#gA</Cb(I/M]IQ9;8[SfZZ&QH53E?F>75)G>SVVgeY
):Dd,E0#dUH+G#B,Q9)N\1dC>&LYHLbRfRB&;eJTJALKdKP[IZ/+NZ)eW=X3#0Ug
_+<OR\#^g11-=gRdIR@=bO7YGP>:8)9b@@=fKe?=+FZ>+J>+7<E[;H5/U5\9>_BO
=Ld.S6X90_g8LFGb=FQHT9:_8fdK._8M6L.EgQOE2Z,2a4C/B\D?.S&ON0g^YI3J
2/K5VcIO#SXC12>Kf?DN_O6@RP&C(eF09B(Z):CfUaT88AL3F^fX0A\/]&-f@V/&
EAXgWdX.eM0=.JJ?J\<N&+NfQ\-Z.(O0-OG+>FVRH/d,8e=V@Lc3/Gg]G9VYK?\D
SDBdAUOP69CH0C5WOcUT_V(T>],\T12INH,:Ld(^@N9<:]dgU\E9UZdNafQ#^A=Y
EegOE30AA@:bJ4_4X&TAE9b&]=TE0J);-e3&=Bf(2=&VVg<:ULcH)<dEf)DR2\J5
]2<]&A-9SSV3U.HU6)+2Pc(_MQO=NI\)gYa<d2g6&6:&=ODX_(Q3^?HQa,&_#WD4
ZSg;@8_M)OWVb:cV?0gcCC/\@8D&Cc=G9S?_;9B[fIN_VT=ebROKUa8V6QE1+[R(
J.C<[IadKAd[KB-9Ig_[b2gX_@SQ<@aeWU?K]JQDg/e?b:T;UUBEHNB_;/dEY>8Q
5K3P<#BJC,2,V8,fX94)FWS04QVC=L><RQV#FH;[XH?R&aZ41.V7Kd1eJJ-+?12>
,BQ1P+CD@[6.00DG^cSXG\#.EDPL;=A;ASUb+RaYJ8?gf56;>BU&6@M5CZdT)^Q<
]T].bM/79aTI0:/9F&RJVWD,]44U2W8Q9g1=\=UP_Y=3V6+1U>G.YAOQ3?J1QK5^
4.;T__>cQ_>U=.cg-C26?Q=HGE3HHDUeO9=[,-;CGdL().Z@F.6;A+RHW3+79Lf(
Q_Egb<e)GCQ;7)FJQ()U;g?ECB5b/4(&QO=,fM.9V1?FXGGL7cXL.f#Z)&MK(;EA
9S>aaB;\,K)7gO=N#S.U7&=17b1O<bJUF4AFb^#@WL1LO@#]\VZ)/dT6BfaSVS-T
bJM,O-HJ-(6RdU/7g-bB5\>fCR&BMY;YY3\5fN##RM<W=;E4P1KVP8]G,US+7]07
a2Cf4]7BFEIQ@,49AZ9VF?<=g:+#RZdU:R0\W]TCZ6=GI9B14I6UM3KY60H.(Ee;
1a9=194dFOWJ&O?:@C3W)Ndf\ZQYL,FaZ)9FU(@N0B-@XOIVIdKUB]1&_2P7e3J5
PG=2;7F(0c67_A\CGO(>3b9+-&_B3EZ[FFDaJC3J,gZd#4fCU.a@HR2WB.6XVXEH
,V4+d23>D=F5)c[Rg^[&Z<gCVD-=]65HfNcZQE@,B-^O^1+MM8)W.TJgfgX(4B&b
U@/F>[D:EX>b2/\>eS6YX5d?@Y1TY>ffd^gESE].E3b\,[86^3ACRMTWD&bd#?bG
c6feN:c.8XeC11c@-PXK.CDC;c7X<=S80PdO[Y;7YNJVHFE1Ha>1M>(Z8DB=0M_3
?,7:TDdf6b+]D]#NB9,D?Sd8CMb-@/NUa>(;M^/e0<26/UV>C?HAeW:B\YKc&C:F
L1bB6#&VG\15+DMO31W.?U=@1d3,>6Fc32<>K\ZO;SH.)0RAY/-[9YJ2[5,8/C;L
&fVHWYY,Z3?=Ma3cEY3H1gePd<)1bH5O=GW/.2E=?B@bW@U]F;,dN=bK-FHL_E8f
A2M/c\U(eE\@T2S2E@/U7PT929^L8FE(^GB6CF\0E;.LW1LRP.C<F)fKL-42VE]5
FYdb2D(\DPU^K-7A1.BQE9/SCSfRGFb)V+9E?_W65_:,B=cN>MVN^W(FfGEA;1fE
R0O7RSbU<:IY.(JgN^3DSSa-.[\\\gS;-R;TA>K>W91DK:c:fNRcd&9&PW;.c7eR
XF<e+ADT9F@LF+X#,c7C;C;-Y\W^+a2Q:H:NReN,3+Zb1DLLa/c2CHR/+@[N#EKL
eZ\C9W81c)U8cCfBZ;G87.ZbIcI2B2c]#B6MH,\\g7B#e45@,3f4:,4[[PH)Me8H
gG[7KUI3\@92GZZG2(_geMJQGd24S,;ALLg8[B>U:b4L1+M78_JVSU5I<0F4Y73,
U57;LOK3RNYT\d<X_-YFH8;g:Jg.5@-6UL9JdN?f^U=U+3PRY;84PfY8P)7\\ca]
UHC93.:ZB336?[TZNO+CF_dXJSFMG>1J0DI7FJ3(N;f1VgXPQBWML^4,1SZCee[.
R7V(O]g,RZO9Y@5FbI@cYQ;[_B]\W5#0,T#VXgcFRF.FN2eV9B_Qg=K1>+bN\(e_
^>-Q_=KZ6NHUTT.8]-CKf?R3C=\O]NK_FD_:>J4cNSZ,4?I2;U:7ZP--AK/DBLAY
C232:e:2M>U[KU>d?1:FD\6-25M(R<NC[Z:f2>B28/De0Aa);3[DQRIZ^/]\Q<5d
.bZ>FOQR\@-b9.LE/ON:RS_/\DLEF2Fg-&D45JN+T:\&885a=HbK\Td#:/;+3;5g
8\7@^;S^DY(M6Oec_+/#-8LFA(&@Re+JS6.9]C=OYH5LM[dVM_-3@b3gf?+,O0O(
)K1VXBQSKaQDFbZM>OP9f[,I6].?AR8<K1dJ184Vf0b]LfJR-(<18[Gd9c2#5Z:Q
Ve;RgCfdCH+4fZLMXV/aT\dR<cTS?2:C&J^Ob/UZC8gXD&Y/MgCD0\EBK8),-:?b
FEI<3([\J)A-E7Y0aO,H)d?:=9+f:4-?c8(A--2SaAeN;d>WXWe<X43B9RQNd\_U
()Y5c>1B.^7=NRH36/K/Y=O\SJ=&.[bWdG<g=)XV,U:/Z:1+8^QA=OZDEK6WCafI
#<MO=c6&4(b<)7LMR(JDgbK;?5If\^7(GML_c\:RYa]7Sc,6cU&V-11+:DKXYS?>
&USZUce64F.f?)&JfdgJ:E>[1^4H1/R+<T&)VR.KED<.UX[6(@QDWcMW23/<K?1Z
UF24+_b(0)f4V]F^PG9_2f)<)QLc[4<I.6bc[c(cbBCXEJBdJ76g[:J)&.Ua@><f
5<e&_FI[7Za,5Yd6_2>C5.70D3#R4+>R#_d5(1=76B)P=Y^G+JVJgc:#<9YL[H0@
9e+fdG&]G/J-^6Y4+Y<VAb.FHJ/#f?->X@Q,S4X@b.0+2ONDcR17?AXO\_,CT-V)
K4&Za^[4D?6;EA[IY^1S-D?e-4FFZ\De)E:2M(=;;Q3M6V,6ME?UV8XBgEHXbc,B
)&^GWUK8C5LMWd]EK0-8&LT#0>+&BI#5?-E/YEc>ZG#JE[[@&3<BBbg.X7GT0:U7
9Qg?@8?=E_5_Sf(0J;]PKB\&V]ZF&3\JGFRWG=TfZRN;0?BJ,L0GLFGBS0,3<NPS
c2dZ(H_?C[ON6Z<VJ/P?D_L1DdR8HVI13Lc87E7d8[_g].WBZB_GW4bB3M@Je;P2
21G@I/fRO]g+-Q(4\4\-+KR]8RB#]UB^.^0><V-JCF0KcfIB2<_Ea=Y3fg:g1M0f
_D\Pb5?GJ4gK9,I5c?0MD]X)U^\S]Z@37d?WX,C?WF0T5U@7dUTY8U(DE.7<XP01
.EI9:#O;dX0=GZ7(87DBM6DTIHOL7K@f5f4d#0WAZ2La34&cfTdC4=Mg9[2]M+8F
LWf;3^MUG30QY)YSAD.^Z6KBfY96^&EK0J+[/SV]_/8407/YSbXY/]VfR&PaG;:#
e4T]#D@H&\bZ\-^G;B^:^]D;2VM,PG[\M7\S_g#Z.KR75:-Y,Jc/5+@2&AGLGe@K
>#H5U;J<XXR82EfFO+E##J+22=G2H>G680\gBa5e;;8<J2)C-ET@9gX+fV0YMR7I
(df;V0AE.Db@c90I5aZ0S(K37&9::&ZbU0b\VMdY438I@YKDc+fFGW8#9S_XH\?)
8FQ=KJAK(IIL5_?0-9AX,L:09-J.5JVJZN>,O(;[(7MH04bcc-YX8?M#R6WE(<OM
YWR99PX@&#II7CPbVN]VP+]]+dLKH72:-gQL\\L=U+40ad1?@_D]DU_f-Afb_HHC
c(<SX^SBSF1HeY]C/TPF:8IegYObYMU+a0+P(#,LgM7;RY/VQB;I]0,8DTKV3GE@
OaZF7ObN&c,Y0Q<;1;&>9S2G374ef(eYTOd)c#_&@?MKPWSC_f[OO7N?CF^Q_dI0
c8a30Ne1VDDY=3.1=DD)G.a3<0+Y^[0g1K]].=P,Jf_M3TWM_9;)63TQNcX\&5NR
5W[&_&WS&N>aeGH6SPSZR.1ZfAB\=EGVODL5VWd-S#MSGXfgFQA:FHb)=D,T^#g(
X7bZESBK^e393BK73\4DGAL?8Id>A[/Q+^VU+,F&fEgL5_=V+@C@\>UfPA\gY=@\
UNGS(LK\B)CBC2Z:8YV:DBSNQ/OaU<;g2c,cLaP]<\)gH)F6+e4944>.]ca=7;O6
DdcA7eD(L.C&H:1G-50S+f8D(;YQ/g/A3^_;M+V<g4EWcT\ELR<X&IB8B1]T:XG0
5ZKJR/&7;MY9L#dRSN+5].\<[g+O3Q^ZLL;&8#:?)T4/9G/:K2WK<H/<&9a?YE[(
7M_4J.UJ?W;FOBfE<<:CJ^E1:=FAMe;4aOLYX[;<CdedWYW-59eGA7H0)cOKd2a0
^ddGb<?I6e=DaTbG4Y8BU.A_Dd/_LXWRX]R,BABfDGI0,,0C2:N/8)/E1_NIT]9P
W#aI;24c)T2^B;+8CNHH+fEMFVI<NWGN963B5\L4^K6Wd7\cg>Y34<?)SPTV\K@f
XYBA;P&eMS\.X3IEd.W-JHTfPA2?b3.YP9\cC<.\Q_-53N3VW5^PH]F-g#d4M^W+
UL8<QBZ&&_\N[OR6Y/+7=RZ(Q4(:8\G3SQ+\6e<E4/T[C8SKK&KLdW.Ag0MH:?E8
+<8TQ.YT1GMB>2S59Ke(?U?K&c1\BMXHd;N\G0K67_<I;DbEgQED,.CA^<MX.4W6
E2Ja^LJ.JDLZacSI3-V3E.M]([aNZ9;L#gB6-A^F>:Xg+JM.E];S8Y/Lb[?Q7V(1
.Q@Z<+OSUC+cd4(.-<OaPgf@5[588edAA&&U@@PFD5+(C3Qd\>11+3U0Q[H5MQ=+
(HdN_Gg>:C@bb8?4WP>7+ZAb6B^9+_^ece@2?B]KAb=HUYL7H(\9@.<YLT\eEa-:
_?Gb._YFJKSQ>D]4MUEY1)WFaQ;@P-9G.V.?=/aJ/c->02AF<PJIGZ^^8:V5,Wc[
]@49U;bg.bR>/K)WNQC\MdLX,CM4+2?b<,,OcJX8+M(M+85U:\WM@F+_19Gfda,_
fN1Y8DCe]<<f>fPc9XGM1AW(H9A8]g9681YKGa_(>+R;J]N\+W]Z>G<>P_^4gc1)
JOLWD5;]?&aN?A=FM#\8>+B:1YI&G^]9\49L_9JQ&:;J-E>T+2FW9_IHF3S96P?:
:W11d5(e.=8Z9]ZXVU&e;\N;&<Eb\a^c0?-TL[.2)aW?,[(>^X&)+_]B>[0LP00,
e9?KQFLQM0</D+>04A4/JU0fBQ(2c1T-E?Ad;LP4[./2S<87aEVC)=aE>M6G?A:@
9?@A[C@d[);ga6@_a3G3DOEDLY_>48[2Uf?IO(\f,IeB?YS3)BF&<G/C0?A1.4Pb
Ee8Lbg8<e#ZefY(ERRU^cLY\0PTb.e+\8BTZV\P[dF,9AEM1]=T&&AX@TffVCb/6
2cZ+FTHYFT#F]W4?S#VDLb7CS6NZ9@_7?7#/Z4Wa)AaR#b(/D,[gJQg<5-9]4H(@
6b91c8gZ+5FVN_@6^I[9F](.E^6WJEgeN>V&X08[8X:4[d7=07_VZ+YCCWPc5eJS
WEGWd_Xe-:CLeU[MGe(@+-W\S)<?I4IY#C=X/]QKL^-JB2@+VDCN_()[DD[aV7I9
EOXDV#FfPQR:=5K=6]=L4:BC)+E=b5,ENJW4Jd]C9DG=I6cg\X/&1ABN@1(IbB&:
b0:2].H)OL4e71F46ZRG)dER^\R?)Q?KLOccf-J8MBe531.cA+UJF(W1]>?Td;6c
0A(\O7cM):1QHRQ:C6XVU=>0]454JE/PWe@H1PTWDB,Cg0f,gf@;ZIRfMCG=:a73
V6?@KJgFK04=0U>2S18S(b=H.F#7KJK^)=EE/e2b[TOG+deP&G_g@dYcdY^]QNLN
1TH>WH@]J[9/GS?HIMdea4CKNEIM@[cXaBg##8,3Yf1[9Ka@1?-1@C6?PU)H:ZSE
8bdf16V;Z1?f3<1Kg4Ab7E[5T1MJY_B)557-5AU+dK7<1\+1b\Nc<AG_YH73Yb3B
.^Z-@aEA+B=R>AA[-B=^L0;_#DMg9I[.+SP,(9S71Ee:0//&WK;NRMJb[\f858cS
<G^HKST)-)-49B+L<-?Abc2ccAZN-:5C:YLWe9JF.cWLS&G0@7TDAA1ZIR;V?54D
(N,EFU90[<,RL.0C3.&^9QRCN8)LO\XFJYJ=.0MKg\d?^#[_IOUEI0Q<0#RS+HN0
gB3#K.Z3+S&5CbO2eQLE.=/Wd5b3c7J@Kf\/YB>KCbba<7_W:d=WP]g-7;a_af]#
6=X0&2,,7bN,80>;VDd]]3^XE1cCTC6=e^T@U@W^OG>-K1JK1\bK^#cAD?YYC+=8
(d1X=cV0>7\XMSPKB9f?+\CO:_,J8/UUPDJc\QgCY,Z7)+5M?V2gNTB_V]aYB&KR
,gNKMZPOHP=CCM2a+95MA]P[cWR/E]UAC?DV#M/;P/#:a@>P,)J@H_c.2C&(+<B?
TfOaH=b[CQ+JR[IK6N\Q[T:67Z]0<]@9(06aTa^SJ3D_MO<B-Z6DC97dVRB1a\-@
M^Q6JI5F3S3QHIKBF/(I#]NDPM[Ee@TO36Y:G\HPYT8S&2#T4OI43Q2FAR^RCWEf
;UHB8T-<A>d5D2Y=(J5fVOgIYaQL,6,GM#C[8YKRg#_K(FJAd2-C-f;9f:Z0@S^0
5L8=8a^g_GLgKR8AbIg49MfNWKFCQWEYRb1?Ja+/&C?I7#NKMIU+CS+N3e(05aAC
,VGGG42O(S=E?#=#CQNX;XBUg-4H\?2Mg1P9,6>?4g:2@dGHA_X=8X.A,AZU##fe
=_SEI5:O[@D5.G=Z1ZVD0\aSTC/DD,/:F[G1gUZ(#MDR#FI>J_DEGWdOO=+(-I3e
bXSX10&PN[<BB/09=LWGP8eg6J\N-;/=D9_SW1R/[(BA_F8d6@8]^[1_BHG[1M3.
_T^@>M3>4.)L3.[:9]QR&D5gNI?VA2U6@=8>f5UPB55Jc<-1>XDKIOE5^2_GP-/\
82G6U.UYB&7Va>bD3P?<1#]#@++E/KTO@^BOVa.d6+^D^W[QG;L[+cBd9.]UY;<.
++_Q)aKQFT.YX5-Sg1M\>&-eV\@[V9TTK2.d=>(Y@3M-fZ7>S2()eZYZ+>dSJ3\>
&)^Vg#;O<4D@\_7OQ/;Ic/#d7;+;@9e:I:YcB(EL(8CEGTJ/A:C#I#cP-7+3a6fV
2?XM.,^Q:@9@c[F7#d_+7f=P_HDZ6F/-^MV=3LW>&97-6aR&Dd#0[dM3&N4OIV/3
^S+3?g5,E.HSDf/Cc/b,8QZ\8<3TQc9Z;OQ^W,O2+;6KcS;)eC44RY]0IWW@\A/C
K>bI&0^<:VZEYS^6_T@\/Z1>NFe)_)c.Z@a3A_HMS^\4bH3b_&G3).R&2:Qe#9QD
a,?3#7MGC>F8_ZR570LASC45V<58?\.de2-U:XQ-c,c0d:#XRK[_-]\G?1METe-d
\+PW1H0@e926Y/SM6^-1]BJVUPM59KEbEC,V?-.+9AMAPF^.2OK,1WD<4QDS@<LM
H[?@<745gU;&a-Y>;#Ge.a<[a1Y\DQZDP8IdMX+>H=@^Y6/+9+a,.8NJT3NW[P/f
cbEGfCe7gSHQJ+<6OM<8[g9&2,ZVGHg,W)K=1HFdBg).0>E,d(0&Q0e6e.8)P5aD
U3\&#c)U0@GBgcPPV^@?,T](9JTeA;dd4?]#3=1&GL?Og,OXQgS#0+CVP_\>T8@]
P7/R<b=/T6IL,4[((+F.XJ755QP/O+;?Y.I0^,,;M3Ld-)J\<aBHPR>?L_bO^1Te
2-Bf]1_fE/@]Jb,UbH^3O\eeWZT#UZcVO=LHG7=G\E?9a3J@/L>PZQDaST.\<I)8
M1R<Kf(#1:SZNKK@KgZ+)fG[5,&2L,f=0Uf-fT,O312]fg1^-XQ6>5U6=,BdUO+H
gRd9HEReG\5LJQJR\71GZ28^E[^WERa5)LA6a6ea;cD7P2VI7_W^X^A,<0dA(]dN
cYM,HFb^36K;FIX@YUG9Ke/3EO<8>WLb9/+8<KHa(8JUV;^1UBb4AN:ZZX=d[CCZ
OG)\#-5@28CbF@E&QHIW@2VPKM\@@EfF1G8W,f?Z&I/]9:28XgV7Sd@_XM=89Q()
8A>[)&#()ePIZ1GB=WQLdU-I^4E8CF.QT,S>+]BW8&)X-e4OK6)e_<I2e]+W6K7Z
95QO7L5?24XU7,-gU#-<O<8JY[<_OT6eeYaI=;>F.NCEJMaeWQeed=ISUUY9QO>S
PbC5L5c7]&d8b?RKOfQH\28QZ8,Z>4?87:5(VUfG4SD[f5SJ&P,I;I3VB/:6-M(1
]e.C<N96@]cQ>JP4Cd5&T;9JXO>YTBHRAd3QM&IL(0ML([,[\J7L1LG-V^02)LJ0
bZE.Q&S9LB6VG(?;,,5eT\J0M)RTKOD4;_.3?H\b)d]3OHeUf@MQ?H<_0X[/BWIT
0Q=T,3N0?VKS7;X,/Wc#R0>=)RA^X-CSXd5>ZA-MS1=B26^)\D\MX<]0=:5NK5PI
\R\1/dFAUO^()]cTDI^K(J+D,a3(E6T2C)7Z5\N0F6H.6-Q93J?KEOa2cH9Af;Fb
U&,?bGI[D2[.S>[7NI^QIMU0(>-NU.K5+;ONIB=SQ/SS]O3+.EM_TeBUaVaJJ-Dg
M<dFEeX<J#g34/WC0W#>?[_.ZC6+-^DGR&8AId)[^WgUJf^]f5^#<(X/CQE<YIVI
EC+Rcd]XVaN66Z685VI]bd5USfe<[ZG_Ye[J/SfU2e<+OC^SeD2AR>XR,Ma=YPf<
D6[#Eg<PH\VC=W6GE7ZZ_(8:ZZY:Lg3G/SCD\3^LB(H[7Y#?ge85&EO,;>2RV-S3
VaQ_PPIVV+S>:,E&Z8.O33-^2#YJ9:,LNE@e&7MF>038J9)^T02A0H#JRQ#bZ8Qg
&NZH)@3WO&aTOTG-SOA8P:WA8AI+(L9>?JQT:_((,)G5bW31Y>UcGUH;L7\\LK1N
VQ_XcLaDQIRHBW2T;@Nf/\0RF7RYEE^8=^H(g77HC,#2N8OB]-c#N8JAP>9,fJ(^
3@&c_HQ8c.9RF\/,I,EXUQ^LO.CC->b8QN;,]@Td]:SNNG+Gf++R\eW[@3Da8\.1
Y>F]W=/R:957+bKB;Hd._RLH@/3EcLX[J,4H)+Z;MI-E-BcV7bb?12,39\Q_DB<-
2AHdg;U;d2X223=_d\#Y[I3daL:8HaUYeO(R/K;B>R1.#R9O3)/LcTbV&e8JK2,]
77T92@B159C;:K/>,^RJ]2IG5W^.KO>VTLKA+4[79\30,ecY4QC9K./7@\WP)\Y0
0I>,IX3N5&7)E)&JVcJG4&7=_cIbVGIeQ,J-GEAYWAFN:/U-890K164@+I850bcS
&Q5DT-T9IF-dQL5Y7bT1YFK&2@cR&bT)2+IR=c[:-^I@P15fM]D7P^DgZeH@/D2B
21MaT#KSL4^L02e0L&P=,7?J9_I0U=#B@>Y67?fV/W2Q#g+HcD0\G0,UV-]V\Z=>
#LC^W-MLYB8HOc^d0:TXIbTVREO,T)3]2(TCZJ0Oe+AM;_9W[+=WPcK81@HX:V(E
aAa,O)<^TQ6HS18GXSR=aV@e&DJ6V#@S@(3DHRQ#UEa[.&0^DHIZ>,g-X9(339@L
+B2JBI>DLV[SD?69+A?CV3X7?/?(U]&=ZA1g/f2H^?B5H>KW[,UZ.2[f0^XHB-Wf
X5P>^[,;1AEAGb,-1<Ue=<C]6ad+_<TE41a,JIC59-S&O/]\NWQ?#ZJJ03^Q?P46
#&e;E.-0cFF8]AIE6(6+F+@.21Sed;3a_.dPP4gDT6B2NZLNW]/AAW0WeB6PO-S(
ZN[G5aVIVMS:L?D7FW<Q&CXe9=0&^a(+6L.b?2#Z?)B=^c(#?e;)8,25>OP,1?6@
IcD2>.A?eL/0<M.RNW,IBD2ZL?5@bM[;-#=3&)L,6_X(+Yb,.Ag(eB>U1I,WBQ]E
#3e,39.IX\B6VF.(2]7(JGOg^-&b^,5a2/HWH[_LQ&]+[c3PeOC&]&]8<=23HgOW
EZ],DY+0O5fS\I6,(XT90O0P9G2U3#]T-SfDL>NBO[9A4(U3,X2PG?0QNMRTTb.K
@T]fb<S?c]WCYH[//O-T.9UP^[VR/Eg;bBPRN-IQ.^-0aOAgEDW@9F#T=G8GgHW8
L&Ke@eE/I<A+_2(8Z?/V_Y;)e,O>cd<eU[-VKb_0MG2gVCY>]A_NE:\U21JU;^P]
0VcU:F.2@N2F?+Z1SbX\&L)3ZW=G[;dRMgL.ga]A\g.a_d;A(&a#<GQNO)Z6AR7W
CD1X+@(RKN.7Z&;gS[_[WO^GPCAcFM4g?M29cQQ.e.&bOM=]>/H0\)b:b8a:eXGR
7bG-7QWCXc(N6:5[GFHdO;6g_UBLX&\Y?93b#MZ[L0W(e5WV@02->].U+&+cO]&_
:C<EWF-G/Q&d7>6+M2=GPb4f[e4XaDKV/E,c\OC:QQ>:0PZ\653^geJSGD^C_7[H
1(c=d((BQBXO#PDR1]I>GV-@,OF)f8>&eHKH&AI8BfdGeb(@YEJ:+-[QB(fHTVGg
<:)WI4(K1FfD2M:.dIef480f0(bdZ\X;PbeXfL@7ST&6F_3VJ)48O=BcIgO>(L(X
6a-RF>cZ+=,<bN/71WY7JZ;Nc1f8-R8+PgLe88PA2BV-1XH,O\<#+JMC#UF>?Q>Q
U(159]HLc]K6]^>I0.]@#IR8I1)8bY^LED\b=JPaf4RN<^WYSJK8(Z.1UfMY.;AT
K?264c4A9PJ>TW9SP2=5\Zc=ZQ8#EAH[Xc4HE9@P;CDd)6G>g.B;:.+5W&SPbf#g
@Q)42K0JYb#JX0Z>O1>Gd_.51]9U=+2\GO(1NFU604bK,@:((97L?HXe82YP7+MI
)>?YX3Y--?9HfM#);3#=CLP/H#Tb./@#;S2;@J\)=^-dbaM9@Q3NC>&&WW?Ng<Sg
Nd85@M6FY\cOJ;VVVSG5FH]CS;II0K,DHPN2gY]eB>:.V;e+R0f&a&7gXFFLS644
^6X3;Sg;;5T]CWea=OM]Z.adZIJ6f7NOV@c+e7)JeC4\VNg2@;HT)>bgOXWG&695
EYbF[-@EeENJJAD<NT+K2W,J<,_,&]MLb5IKRY>77B4<KdMB.9.?T&e<?3N)7R:b
dEKQNCN>)g#V[I2O.:26NWM5C/L:R.8>888-4]/8#\G=.D(BF(XIT0eKJL(aBc-F
\d1/&6WIeIMR4>Te&/<eZGZ:Z5F-\76FeB0f6SY0CNIGCK@.W2TY;#(:]PQF8V@E
,\5FO];E:f7_+X\bNM.9]\?HdB3.8EO)YRTcT_Kg)3P&ceVeL?YPO5?CGKBA\PcW
T1(1K7\[6F][4YE\:>HLANaU>[.b8M@FHI\\X@Ha#@6R(-fW9aU4YfQKL5AB/.X@
^@(X_4IK516E&-/D])BR0TaKI:.83[W?+aGe#-Bg76Z8=?C7MDKB-Db(1?BJ0,(5
N3TN^&]-P^GP]#^K]&3B)eaT>9/e^gT>a6&AG\1A.gf)6dT_+H=+I,5USRCf68E7
dY,4FFI9)/=8BUTHEbZ#^9eA\#(gd37TBJ,>;@>daLFB9NDBCUgfd#X/5<1?CT]c
(2AM<e1ebDA#<:<_NW??H1-VR16BBZVJb4Ed#,.MYJ5;g9MdG7<AbNJ#41(^Kc#P
6WP-2fN8D)bd7^VL2CaKY-7APd^9(07&<1YN;L7HDCZ<)^9ST7Xg9FBagR[[<85[
S79FF;@3XfB/<<&):9#Pd5FH\e&?fZ;4B-5=\:COT,\-&O)55:d2-d0Bgb.JCB[,
NVW(3>1YB4Uf#Jb_54b=0^8L_fTf4/N-/51c>O::_MfD\IE\+WX&=A<WO3BXY=Q9
>P\GbOAe/5&Z0/7<Q[B=gF,>E:GaY^86b1gJ2G^BLH4=01<)=?T5N+HFEba:F-E<
Z69AIe=P8XFO0HF;,=8:0G,>(GCbVG-JgFY2G,=SU+\aHLe_F[?,)?AVM8SYQ&E,
5Oa_8L15KMB25I3R\,TY8b>U3b3?-RUY]1U[YBLC?:8[G+<;(?)c5/CZ]I2\GJeP
OReZS/gB<]f2]I<0:];gG/.PH_B<531Yg0>;RIE.GB>:4GNTASCN^NPR3e+J;5>U
&O?VPU-.9e79KD[<D]fcb.J],TC7SW:L&[e4(a<ONZ),/G2_C/]J#Qa34^1D-f-A
bX&ELQ->3cW+@YALaf/&-_?AY,7]=(G18Wd4&O,Z9;F:dS5VKU_T#[4?>>Lg5&DD
8V-e26a?MD&gNN]/Q]c27&.Q3Q-H(/=<3T?cECc<<:bJ-a?K9<.L9MFO\^@P:)\b
?/fT&O)-DH&[NEO<SB?N3^7;4g(MWg.0beEKZRQ3e0M+MGQWA>H2IKQ2.E]7)ZX]
Z&J>D=)PSF4BE6(\FdIfM_@fHe]QLK\<85@N+)^MMO47G]IZP_KX63BMP4]XH(U:
XI#=6c(fSV=e5>,Z<BfB9=ZKb@+PIKH@c7C3#Rb1.;3#\X[\?#:EG9@KJ6C#,bL>
6^YP]7O9(KK&_N\Gb?HZD6a0.82BR<8(X=(SBEg9J5RQF<.7L@Aa^59W=Nd?DB,B
0[8F8SUND?)(/)HaBE^:^IG(T9X<+<=]\+OCKV)N[>.OHNObRN<.W[8AG#TTO?&0
M2YOOa^HQB;#^E]NOU=V]PT;fMZ-gc(QH^047U\07P2UY7Z,HeP.,f#?Z@]3V(G^
ZN@bd?+]C+.H;<,9g7I;;V7I-<?-<;^1AVYdJZT5?B_-7VFR^gCFVYJ1b?WaML@3
LdH[gc1LR3+X=@dF.=Aab589_C#F34DK,6Q,PLR^E60\H,YMgeII^K+\,^&I<+(9
[F;[fWP\M5aU::QDTG9EagKa4f^#K>FCF\E(a17>OKCCNJMHfVb8aA44&TEWG#cf
\U,W8)[YG:=HC3Zd2Fa8+K5FY6L=1gE#@^^KX)bTQf8R<&a>0NB,;6Z)Y+aL?gUb
c8&^MB=(cb4.>[\I;V[US5e_BgUY+KCW\,;T6\AFHSXc2PZCbZY-6[A[[R,V<?]^
<VF\X>,TM8ZZY^,=K6;gL3;?NL(=R8];?K&,C5?3X86/e_K(;\1I0.)c@NS^[RRN
=eQ48W?bZOdVQ;&=0a)8?K#5:^_[\,+S)a-MLVZ;6ZA&aQR#\5KS\IVEf(G6?f3.
cZ0,B.ReS^VN3SVf\]_53.N4O5X5>DHRRQZ2QS,0.[fK;gbA5E83<bWg>e<>CB2I
HZI,:U?BK@T\/V;0cg-dFf9@:LKGGbdU&)18gQEGX)EgMYLeJE_P?6I\Z7<<fC_8
3_PYMc-1_9:d29b\Tc@)P[I3b@U:\^HXQ^&(Od(0C1JA+@ADOMX=Od+b-g43[^7=
abIdf8b618?.(fH)),/1f7X\bK<Z8SCcgQe@5V6JLf_=;fI>@=gX#,aB^_ba24Sb
bM6;8C227c0e)-?GeLQ_4NLI.gNX=^B7Z3cBYI[Q8(^M2,,E]TS06<2/]aM5QD9-
5a&</I+EJ@JZU19g.I)\PI<EZ)B9V>N\/Y(VAR=>6Q(9cU+F41QWgbOfa2Z7\&OE
2]63TU)9;23W_HU)IC)@=LIcd>SA,;X8aDR)J7N7B_LD]@:?7<TS1EP/4aI7d7UW
+I8DE[](QJG(V6O.d,eFc<aN1.^Ng<&dPS+C-=c3;0HTP\R1G,VV;A.9J&RbWMgS
?&PC(Y0@K1V_ZQW<]JQK4M<W6#ZJS(F0V7HI-LA@f.0gZS9e(MbAM5(W13;_LYQ)
\)GHQV56RDW0P7:LV??0H-g#;g^FPC(+^3e4<a?K:A/<a8Y=(@;JMK)VX];&#CY5
_VJSZ:_TFZ1X\AK^HMEeATARA<H87214)JX[XP7P3L-J?[CNFT8N&PXa]a90BOL]
,6f+\OaS,H2IUX)L:G2<=9^3YBC\QcW6<-9^g+Kd_eb^3T#JaRDYR&ILLd-CaPdR
Hb6a5bFT71K<[J0:AJHGGI]PJ&a,YPLXRd7D2+]#1ZNZ@cS_5[c55ROUV:+^=_SQ
<]:AE5U@3<aDAJg]8Cc[\@b;.3G\&/c8e3OSVgL4<V5)BY5&L(SQOa]84D:bII[[
^3\:N,2B56D+N\A2)9]<e/QE9&PKg\9VcOAQ3a7@b&\CUL,d]7H26deQXK5^\U^?
8V1>9,\dM,((Wd8UVVK+,Cg.#fO:,)09,2YL/BNHTfcY;SeX@:9?W@f8R@T\#E^2
2><A;VZYM<9OWUWbIYL/SGZJ)?_QQRMe/fM<PB],FfA]CDA^[ZXMHeYE3gU74O3<
+BG^&cY7)X/cQZ[Tbg/aQ8bC@cK8)D=AWAXXP_]ZO84I-&554596:7IETO#OGXF@
]H>64UJH1(MCOQP)[6,WAYJEJ;If>gdPfI73L?8J1\fB;)/gGV_Z_)=&H7aVBQG2
&4cg<QS[;6HP>XF4OXMM>#D_+9bL,+-b/3H9#1(#W9:7g9.WZ(b@U:,&>?5c>\bX
N7d1cL^(H7Z9c[cX,GDS((,bSD4@&90T9RPD=++T_.A#aeV2Jb.(-,P:#Z(.gD&B
(DO7E1b-,?=S7G[=Y(O)T]?E(7CJC,?3@R?dOa>C,Y;R)CC+])LB@eX4NB#@+)QM
MMP_dfQcF90N-S;-8G1[H:J2)WFOS23G-]=[&VZ\#Q)@S\+=?JHAe=fG9C+\Ye3;
IZ9?_CIM&2ZFYG8@,8N?@0RH#)AT-2M:2EBfJ4fC?@JGgI(00(2V>/=TM1g4)UA5
WFYIa<DM\]7Z47#X70LM)-O4?A:Ved8b=D.f=3gSIW6]8)O/,3+I#&c^g(<&0J3X
_cBS7Tcd_aee,<LB(Re>SMFU7KP?VXEQFI5fK?N0fG(J7L6,)TAXQSg(CbF(<LDd
EeE&]4\ACT^eY#eZHfFIZS&#>HC-.H=T\2R<RSdd6<_2JW?W28WZe<PJ?-bVcIP9
GJYNaLFYfa51D#0(YC3_ED+e[P?Q&g5K=_,]d_6VVM+WG2_:Uf;6gWKO0a;A]&]U
N>#,_,+UQ?R0ERG-3^&..N[;#)G-DQVbcM(WgB\4>\QQ._)\8BO?d9F[\>aG@D?&
S3753R<?JFH6MY=WI]/,4+R.TEV^O08(DI]2R+NX#WL0=?>K)D1Y4)P3PW#:@4.3
5bMXO>-TGA-S_1ZZe;g3e=06J+^\>?dS:CG&C#_B+Z>LJCZ:H_a&M^&Z>90XBKRI
./C&N2B-&B3ZDbfY^58f1c^5N]]P+)?JT=\,U^L9#Z1A0(MLTV//ZUPL45FYg]\B
H/BAWId.C>HA2/D=8?W6;R.I.T#MALO=6.f#1(d?@0@&1AC=\80ZR71FV;1&Q3:&
2[H9G&b:,aaHLJ?4bW@JI,a7D.KBGE==M)V;5&F-_S.\0@3f4(4gcY,EV:AMRWbD
OU65ATJ#2ScCI;aI+:GP,MCWg=HQHCGNBUSK60\5U>\ELG\(.(U;0_U:\6&fDX_V
Y2L^/PASQ,U5.O1eY(dH]7IY9+.Y^1aALO]Ug<U_BKY-CU-@PJdLdRe[;?8gGON,
bgG)41AWQf1_U6(//#L+JZ3CaM2),C<&BOMQUgU&P-b8+U),[T<BFSC)_+JT[R.L
0G?f6>(EPMOVK[aQPF-I#DLVO5,(JJ-C3R\1=#H<]7#)5g^:5C1[VcARWKPW[RKH
V503dg)2;:27R[2Od_UK?B&Q14),87bOgfB/?Re&@BK^CP\FNG-TCQEe3GfE;gT1
VMI8_Z1<a6/E3,P=HIDTY96cd3a??^1)B2W;PUS.bO4?RG(FR3P(bdTcBXQG=2)3
bS(?D9c]Z<Qd\9#B906RCINW^MA904JJ8\HFb@;8C@1?A.7]/:-3M/fQSc9?>K[M
&fE]=a/c8^H=.TbaE//>ZX1]:V2J.dLP>1)0EWdH.efb[LC\.0cNeH1>CI=YfR8D
Z+^aGG&.W]+2<0TW#300AZSI)R^>0I(]U353+9SEM^ME<7d:KPZX(E7QEbaF.\\<
5.[2Dg.Zc06K.S0Z\1B8GXgQ])PB8/7#PN\b7^b\ZeeB4A:WaOA-)DMWTe2OR1V9
c[V,[Q#Q1^UIgFOMdAYbP#W6#.2Ud\5\69CH;YAH460X@I3KS5EE^[?+g.,0D4fG
\CeO]&=gLR6:G0SR^P_XHA.4)efg-gCZD2HQHNd2;e6-DG;^Ta&4L?5c80Pb<I2<
2SA?Zd/g)e&LeQPRe)O0>(2]O#_-Xd.TGSA,,d6N.;N)\DUBg@J/O[a[a4P;0a+\
N)3[?OAfbVU70E(D.S2V.8Dee)V0a4GgB1_@>+:I[]C=F1EG2<9@D.Y5>Y5Vf[9V
IOD-ZCP2HJHK>ILG9^3))VRFI;1)+e[[-4FU]]A/[:??=B>NK:CL.92NFSdNEag,
H(_SG^:>SAYL]FfUC(a_,6LbP9V;53[gSeLQ3)cFgU5\MA>Q5d=9VE(+>CXX;Jf,
LN8D6KBS:=T,>^-HY+Aeg5++U(NF5S-(-afC_U,>Cb5aK,AQD_0U5_@.fT0g+eLU
&2DLV:FcgM>]BS?9(3^5M>;L4X)B-YR:+,,SKDfRJ2M;6]7#O_Z_-99[-?XN_^S=
[&[&5aL\6-P.QA-AcYb@W1?>LJfgEL2Z?=Z[6WW^>YgYBc^>TVe8g14GIMT1BF)S
(PI44)VT.(0c[dC(JeC8W^,>?/>4XPg-W23L&d^#LeC#UZ8:?Wfad_JSfYM7V</S
685<g^@Eb54c/g>W)#4ZE]C4\TPAFXT,UC0P/,R@H0Z)I4dXK^Y]YBN6YH0&(faQ
[JBbMK@J=b)Eb;T;WJWLUL3?9-.O77&B86XW/NQb<9QPbRA=7=1IUK_J9U7XZ\Ba
c0HJ.7g&#H0[[;QFQMe6NUK\^/gbE/.9Z>]aY@D)PEBbY;7YgB_8K=@SgP3AF1&-
ND]??CZ739E(QJ.DP-aXV,--<-g#9N[2;6RH[&DZ+>b?6-\#J6B+,Id\4\Qc0(#D
4:HV5d5&=VD>.DaI7a6.JK^,>^Wa9A2,X,&?Rg]1&>4Gd-R_;H3XgDB,ZQXH.Ed)
9&?[\_?bCGDW;:ONS;Y-5I>1\(?gO\=V:d][b7/cO5JYgG;1^6CA3d>SD4GX#00A
)^KcJ-FF/X&EES-5;df9-KC2E;A6HB+N=NP].3:C_dO-gS^<-,\BTecS6Y6MAXB(
G8)9cR?6B@:?3Pca1_g8GZ3UP\aS1J6SX3A(&2Ud4a\^Jc,JFee3XY&@c,4\QfS0
:4g82]Tg.C5B9cf2E.JW>,TLX7EL.2T.;^#@+#W_DF<CaH(cE<=G[[7\4^>IRZf?
;/Q@-CDfKg@CVWM9K+ALT4LNc=[F^7\KF9.5eBBMN/Tf)C.00g-LKcN07ATPb\IB
f@-8e.d-)ALZKI;_UgeOCSRZJ-YEZ9D_QS+X1:A:LV,PQ,FgZe6J^T>B0\Z>F?a:
^>FM-D<?SE)CcaS;ebGR?S2:W;A[1IUc>UZU33gCOc9-<7Q&cFRZ_>f,])3ULE@W
3b=4WI1@^4R/3]O?GdU<:0ZJ(TEC[TJNS86c1Q..7dfbK17D^K>3KQ[Z/>^gM)0J
4_Pd?>,6c?5]5Z/U=+_J;f0U,aI4IDOLTKa@<a42YPV]@K=8EJMfG4L=M=GB/\83
bUg[F[VY.GPa=d->K+I4Y0a4#eS^T;J9?@U[Lc7c0LR=C>0;PQ(2A?5<I/)G8^Yf
7KQ1fE)>Y)L.HHH#T@Y:@0[^<+8gJU1(T^Q]>]AS610_F=D?:A,Cf#e+M?G\\XQ\
@V@&KYJKe&(>,CEVXAJH[SQ)7,A?R6Y+W0&YEGXZM3AW?,CHf038afPLBdL,?5:D
8[(dIVf/&g7[&U2^2)6@-EMQB6OBXS_-;,#eN)&.Y2W):eQGe/E>0V,=7M>E[DDB
H<-@SO>/DN]ZZ=a+3]Df.,+(]&:g[L+La[gP,fd8d9dLK-=OBJ?0BTTCSQ--3G1[
1eP@^eIHZf4UVM3g7/;AaLU/S6RE4Y@(TLVBF#H.]dO:&)CI3Q1XV;U)BE(?7+1;
)UO>_=a\G6SHGJgW(eWBf\E?8^5GR&^Dc_V?)_bA-30EQ&W\O14Y5V_0<_521aR#
2NTR@NW.C+HD:?Ud?_Ec,XEY,U1[G/;e;e+VMXe(cVg2AX(QP8b.GQ\--F,U8]Yg
TKaV@74\Tgb.,7>HaLM_>F13?/N)PRF=/=H2L);&&7TPVU4TWR7?aD+0UaQ1U#Zd
gJ)O7_TEM=HUBF.BdX65TQg#]/GY6KY2OSN20MUUbF/#;><?358O(f2d:TP:;bTf
2ZACP#S;VJD+I.D<NCabY>WO9IM);>NMbB47N8Def#EACZV>B89baUJMG8+AJ5_&
b3,cJ@b#Y5gS62&G.I-6\dLgD?Wd#e:D>O]T@O8f,2HL@@;]8c=fR=fPLAe0>5(F
&P<cQ_S?H^F\AYY7V0#;:J^2YH>4XJJ7_+DG+DDRC/\=E?<RGeRg.6S]KH_-^>B[
7/@G@32(PCOG(9&2SGDA+L1b@MeVL[J_(dYeJGC>04>Y&ST?5)87,#Z6,,61+\2T
IR:c+34V]BL@94b7QXc#BHNY@#LWdDG&@@+#QP:-+3A@E?Z&CJb&E/CY&;;<IX4N
/QLb3K1LA\&&JgRQ:1JaY&6=aNdQG^Df3T(+NHRC-RS6Hda8\SU3YK+D-fN-LX\f
f3S[GGWEG,DEg_.EHPbYH.X\2CV:9)THBLcfK86M<aMTd6WTNO&P(+<f7Y(d6CM0
GXBbO>]PcR0DeI.4427^S=FR.-b#\(^Z<8eN#=KD072\IRR<0D:VZ/2UKKL]RN^@
D+ZW8XZ50C&dF=C>F3R+0^Jc_76;GDTYY,R7#S+&_)VRGILYAd[9343#/V>5UZQ)
A:R[NS3CIbb5b7:OAYS(M=&^KfE<?c>d5-]NTfV6A/DZZQI6Jcf(OB/4a8g50X(5
OV]-JE5f^&B/^CQ6A\MaO-B(b0f-Xd43).<&_0a==ggQe@)WF]\U;DV4G?)Y/UQb
D93QA^+/O&5&;J;X^3)d5\Q/YLIWSed6H]Mf-T(][7fZQ)D-a?D1D;QAD(N-1DA=
N-.3[>31<IdeK3H<eA+AV6;cQcQI0^-&99+)Z9\[2Pf,_)45-CH-146I3[G=_/US
TQK96F_)H1(2OH0+OWP(GD4R@]H?b5J9G6^,VZ,-&#O0dVLJ/e;LQbX76.Nd3@4F
<U8,NEVc#)&U/[Je02OfT8G?IV):\M>9&#YQJB]<UBV##_-f^fJ\=(:Y:^_>7+]4
MEdIU_-9U59/Pa0eU>)\#?dKSJ7)31c,-cH9N[.I>ZST-0C/AC3?[8S6F7B_aEW8
6KbE,e2D9JQ7gYeBCaW3L6[g9LHC@+fDJM?/gD7Y-KgM8L=<8(IW)e=Z7&+EV+F]
Q=W1^Hg8eY0cT3X]TOX_X7;Td><PBgg_KU_HNM9T5W3[J/7SeJXbBbWEX4G\<^>K
++Hb#_)>EB=GY(IHYg/D5<F/,dI-O@HX+;NJVMF:F]LZ\@;Na8cAC;bA;JB(TY1B
C<)F84Z9:J>KYd9?MO>@[OC@.QA7a?e=;C-\).J?9TE7M..WffO03b_/J\XA1]Z<
K8eWBe+ZFcdGe-:.Td1>K5VW08FN&AgNK=ZJJZ1B^_=7\IcTAW4,4Y[W[1:dU8Ne
]-KS[H_(#F-O.JL555WDF035,gg<(#H/f<FQQEgZ8d#)#X_MUVc[gUG_I&FR,VA@
XTAGJFENMI&NZID&5/S@]\1E[SK<65&307^?-g;4&__862@TYGKNVV[9J)^2&a^8
g/),9E3WRGW2D2WN8S9E6K)SG+-;LL/B?R;T(V1V]PXV\52QLL));16N9gW@7RPB
;>@:^f+0<OUS2TSQ=)@D/(ASaW#R6^IeaK3#RQ@5(2eY^TI]c#.Mc--C:AR.gPYT
WG1eYWY),F5e,P7UUD6<MeG@0KR[EbD^=[P/ZXT+Ag7WQd?FE78Z&]M;b1]L5WUg
R4#&N92A-<N,K65;U,MW22WfE^gP7T^T6c8]CAaW@KE_deBQPdG39OD]L#V0H[I6
gCJF7=f=c@0B8fK,DfAgJHYW5f7dU\#W&gFeC@&#K9.G+Ic/YHM9U6X7X<;^<TfM
Qd8ZI?RFb[BMD/-G>K[_9/Y(@8@aG(.;##J=<KBW8T<.Z;HDVLBDTQ[(1HS@;F+B
8)H)[8d:,QMX;W4(<g=46ST[/.0/9^K8.S<HKCf^XOO(OLZ6YILQ]V7R\P9PHUDW
4>[.V839J?F;Z#cCSAFEZRD8X_g;8K:.PB8#66g1c&;OQ8cbbdEMe8)/=H6PS&4\
7>ARb=-^FGg?CH2YQM1B:.<KMc#FQ;W6(;@J<R[+3+ZMF1HY)S.KgRBUT)Z0HQV]
_4:CJ2(TTa5d@_5XT+O&,cV4TSD@?/R<#8g=_VL^[BgGCF]0=C-^HOe+]KP(f(=;
S6M(Ed:YeA1Q11^&&3O^b+^RA>WY.>>@:#_5Y)(6:T;:0Y.bL)2<&&L/LY6-.<Le
WY&BbN@,Z=cW426c]R>M_ZH8ZN^K#7R.[(BeL(CbP3Va6#KH8NfAR#^</)Kc#QL9
Ee/[-A+C58[(4_OQ:GNDLb^E3ZR@E<C(M2S#g<#M0Z0^-FSbNPTd0cS9))[,XG,R
g038LW)]8QL\/ML7,)eMQ9<0T+(fYd&+(<J(/3=,/Y8T0+N4[a]A\_([g5Z^=WKa
AY)/;FZ(JTNc9CH+@\L\QR02gPNf#bgA_4GdRP3YgWSdLJ\,5D6^2]9\TZ6#KUaW
C7W1f0,1NJA7)Df(97U,]>=\F2+7EQQ@WSMQT2^LV>cY:dPQf;Dc#TL_e=]/93,E
\N5)AY:8RRKA79>ESXE+6VeDM\,H4A=M8Z04<)8M?b(SPK@L/@_TCTO)SLM-13#P
\U()8+^S>V-JH(d]6ES6#G2JT,b<8RbVTY]8YTQBF_b44A3-SU=?KMD]\4_B:N01
eGJ;9LEg3C)6QW)9-GH/(_e6?255TZ5YgUFb\T#KaSF7c9K^?@]IPNV_;6PMQd?B
0<Z>PK6B(2[?/(=Q]I5QB3SC2_38=1ACLCUU?8_,Y<[YN_L\@D#3^K;GUL)13.IZ
1<)D0TWR7,N\8_L#=00cA/^>-gNLegb6R7.-T4/@(+G;&H?a&M\T1bM]^PgF4BeB
1Wd5b>A6?I<&Ac&<OHf<)gf6UIEVb9V\6)/:fY59H9:b99DL67>ORK96#0V/3S,5
_^MS>D^SfQ-:V)AABU?]c<M4&1JaP@>A-2?#,JO/cIUX.H;O4FZAa[9FRdK0C2Wc
Ydgb:F::<EWF.C5#[e7EY,d+@_XNOC/f/0,I2U3P-9<US]c-+)?_U7=fM^+8@UY@
Eg5<Y=+^M^B)W(/a=W2YK>N8,aU4/D.7\^^(6A^H;:]^7<[M&?>0Ze;B6W8K:DNZ
\Y\e2^:ab4dL_79FJ=fHA+aEO&YJ>CN8JWX+A^C:B7A5QU++@XFH[V^R+0OF_<AB
[G;UcB9Pd@SC@e64Z^^eUDT4]O&f[43++S3E3_T_f8Oe\ZFKH&I+\7Cd:1(YONSU
dJ^\TJ5FdBF7^9KYEfX7gHJ^dba:OgO7UOJ)\T>77?Z;4_eNKG8@)W/&C61S9QR1
QeZHSN,Fc(d9PYET,D#23dJIdbaEW<:9)DeRZIXf;;XA[dJ^8Q=@/GZ^?C63TM[J
PV-Yf#<#GD>LVL]WCLH/QgMY5e3\ZIHTX#b-@4H.+P5J0J(RaA4U/?ac\,T)UF&_
Z[B.[J2&dBHSU0+BdLY(/.:T0W:@ETI>S^G<>7>PM&7)#=6-7B,E[>K,(,O)Ma2.
@^_YT[&Wc_f7AMF=M#4##O3H][aD:UF.+NI\J38S^5:I>CZU._HfAG+BB5JeC1cU
(>XDOCcH\G@FWI_#[YW+HS7;@-f_NIc5&<HB?K#R5_fFR69.8AP40ab8[a4E<[cJ
L<K0B4;89:>KcJJO<fJP<&J^_LISX/M1BYa1[PA#4dO-E-1J]ZF_HbR2N6CG,YSW
N,\CKJK;\=M:,C]f7[#,cXZK7EdVRVT8_2JHa6UR]2TW>=?M5U5@S5Ub.\::cH.C
6V[((?W.D6-dF.H)gK@@(QS5:c,U[Idc^>9^:fL&ZY73?(^0c([+Ue/3G/Q7T_E&
UP_I<=VK=R]FG[Y?I0f=FAWH588?[]DO-J-,=@[V16Zg/QN2gQQ[(-SWge,WU)1N
,SAXEJ/VH56X)4O8-;@D5)\38<@/\M&&SU&[^O_UE-9H?aYS.726=X.BT&.5Z98.
P6&-TdGF,VH0(A-J9K^@:B=ML-2_F;NK:2?+Af(1,WM&QaF#&67DOKS5)2MMEG#H
J;#]\fa_VU1_?K=Nb]e,CCZMcg6[IKB4R#\#Aa>Y0F1DDScKK-REc.E(G]ffVC;G
c9\/KDBc1V(&_WAKUJ:7XE#IF^X(;1AVYN6VV^/D.2VP0+LY88]0=K],(gFOBbI4
T96e2O?J]R85/b56Y-3]1[aQTP:DVX0ACNH6.1OD])TGHTF#,gAW9#V]/H0RD^L2
31c;-0G[6YG,4PDK2EE6(5RBb[\OJ?Xa\V?d8b3N?9Y.7/-BJ1:M?#Q&UL;ZZZ+,
G_6gU#HUCaJcMH(ZQf](JO)GDPU5#XP-PPH,[d>LDU<]Cg:VUBMW>?P?BH:,QP(V
S&YI#bb8R7EI>#K@NKaX:ZO+L_HPSdHf8,[Ncd#>=RJK1dZAI;-]aJa\NZ]94@)S
]>UaC:&D3)O&d2+d@Fe=H+>bb_4UdE<,Z#SbZX4gYI2?D&G4NW;M:F9\UJ^X6>e;
;JO6+ZYYI8<]FS:CYfE#cK1=[a^K)7P0:-[^d/C8b?Wf314(aRCZTd)+PX3?Vf-I
;WR608(Y=X@/d29.&7eQ_/S:MEfg]8ZNdKKcXM?Bc2eJNM^#a#b4F1CK05fW9Paa
.9g?N+CK)];LH:NH-W)TDX2d0F6;@BVH8ESA1B])&B1>H@-+]?,7L2^gUE3==^:L
8T]Rd;Pc4#QK+\7a+#UeG+/KaS\S6L8+-)a47O(VB^+281H;^]3X7KeXI>,8;=)S
FJ1e-8GPSAEHU??d33QP/A>A=17VJRPGe6FdJaZd-]#9TRVRF>X->HVL<XQ-ECPT
IRQPYc?gXcC^\6Z_6A5GM8R2fb7T\5S;=:-;^6-L^gL)_F[.J]7=.2bQPgEgR^Q.
6Pb8K;^\/?1DI#;,a:7Q-5bQD8c\@ZP+K+(CK1<=_SbWE2W;VDa25ZJOP3d9W<?D
0c/0?CGfZ4+9+I0dSLO4-TIf\RW)->C9_XXTS&J3A^E\/+-SgT:D?#PB8?&_#H77
GO[1c,bFXNCe._I@H-VdKg8+g6)1dC2K>b&_N<PeD8_,@;<8+DFf7Q:,RKRfQ^=[
,KQSUa2c&9c=b+\(HZQ^_R/&C\Mcb2OfE).cV@Ua62MHGBHI^[F:<D1]fc<8]6/b
^[RMT&KNZ1OK44dWNSc3ZDDDP/^DHKD2?]-_Nc19B<bI<fPTFSF#BCO+<XX9c92I
9ca#:>NdaV>bPHU0@L_dPgU;_-HeD0J8W962^7#_=5.)J-./[T-0=S,R[0F(.=ff
[ScAgF@/Y)=?#B]:,6Y_INgMOM4L4;YWT?RKX:aCUKI?H5;^3&3E=G(?:PE&(J7J
B9\X^1+NY?Jd]]^[6W14U)=S\-N+PF?X9[X&+AV.XaC8)H2SKR(gP0?>-X#9G;?9
+5cTYc00-BUD(a38;0RZSI<MNZ]Tg+YBC)MOO<GN7<JKIB1Gc+B(-;1Y>f5BQ0G@
e[@EfSJ(@))8?fX9-?<1I)5FOZEQ3H4BdPaV<44d@a\5;=T9SG>]@182859_<Q:]
5&f2M[E+Y/4>VVbf2LZSV-(#g+K(/W85DeW4M([,g1XJU)ZVgS9ENVGTc@(b0&Y)
5E=.RO+SQ1:CHAda&g]6aD]Z3AF_SRG^8K98E4B_006]Q44e.PDa=AJ>D91&(5;4
=ZT:<]fSdaGE/Z=(.\g08_[A_PS8L8(f]:]+U?5#@Q0V-;@f#Z\[cVNQM,0A>Y=[
Z00/(/@AQ0[VT+V5G)/J6.0C[c^K_fb^?0=3[7]H<O(AQ-:DUc9HTXAX96:L6YC^
,#cOO1Q4^aTN4ZI1eBT/@]AHe5K4]3O_E/Yd)fVZVfD]XX:::5UG1B2FW.HRO1@H
d[+7ZZ?9[?_L9^?I3C:Q=_L/-9^K70.2X,/7??SK0a)<A[J2II/-ef3#C78MLEN=
>76L\1MOC)G(2;_&Wf:5d,[P?2Q/Zd/)gE/A-M?PLP#_cLDJODSLY.d\F9G<8U@(
M<IH#;^<:+S9E@W+M,,.JMCfYRQ^[KRAXL^Z11WQbeG29KPRNSIE0@K4,O>UHeSH
/P5GT-W82^5Db0d+LGK;E=Jdd2/WE[Z)407SeH_1K)_QB3<QEM)eLL3[[_Mf#=V=
ZW-I<9a9>:2G)9@^?L-)818D:ZFRFQY85)>UO>QNEV_,:Tde12gHXaa?22(@ECC/
aZG45QPAE)aAO0>7bM,QUbW9T/Db:V<Bb]?_1d2EOY&FPX-PBX@g#NU:@AOD1B;Q
0f?DO<Q]EJ9=-:_JC(<D<>2U88eWP0U>G-,I6+GZQ#@A9[7.7,SDWfGE+,/D&+X8
+GD/\E4>^E+.CX09>Q32c].aNCLA3:JR6UXT(JCYT/I;g8F:Q;f@;UN:(ce:JW5<
&O-(.>16gVVLF5P[^0=?>MCW_)X8B+:.&HeO6CYYSaP,?V^IDaLLGbN1XIC^<BZL
N@;8UEK&aUd-Z5=T72#XFUPE6,P)a#Kfc=J2[4XW5??)>/+PR&cRcKRXJ0NgNZUW
<EG5e1g,]2H)C_[XBB2X=#^fN<^GND)V;E.6/^,(6(T)M#_RbCX&(47e8\N=MJdS
LY5RID32CG0PfY#d.d(SdG#,g3_Kg_?OT,];IgDGgMg78G3S,eL-9RDQ?H4\2;;d
+Q0_VS^CJe-M0cUbd[:8-IZ2?AKd#OU5V1-7[DMaVU[;/R:F0I]U8>D3(cCO/&I[
[S@(1ONQS=/c<(O?4JEb3c4_<bcLNSA;L5WJ3K@MXgCeNJ&#I;/C\Qd6.:7JVF,I
FQD[KYX([g;]8aQU145W\FQI7NeQb5[EI5e@M&HEU-F1Ne5CT7\PR8NT/Q)aTHU/
I5JN]V.[+=Ye)6\(J:<YD7]MP=+LP1S2BD]5A;D,0]IZ^^)+/e<9H&DQ6<=BRYKU
AJLLcaL;9OX8P^G10[Q#^,UKe/UE^LVZ-K)<(F6K#/\R9.g/3V5f.#7KBa_KWH93
f<.RXWa-+BROIP(-UaV47+:Gd:^^a7#MM>F\dZ7T6P73)PD99Y2O-3^YX+Fe]T@C
PDRNC7d4J91)S^G0Td)4)HB#&gJF3\Q&#c^=@(\X;g1LMSIN^FM<PdE>:+5gTHSD
8END2Xc/JGe0)_Ec#/7Q)\)YQ)S;aG_LSYI:C]4LL7/>PC?3]E=+RM9b1CcBFUaB
B(HL7@,L7cL@9Le(@O0X<R5eT)TRO_aJ\N^V-g:[60W_g>4@G24EX.U_?RgA];Z1
N>28gJ_f,#++\<2+:+-/AT2;&8F9)gNfYK3+[gCQS=;GaRS0+DIf2b@/844aNg.Y
:G7B#H-#:.DObEU2Wa>B7(BFDH>gfQ8NI.R@f\;NYC[B=NKKS#,\A?Y#5HI8)Y_Q
Q]>Z#+bN))SG:#=cfS8A1G;g0Eb6F9<eZ8VPI2H,[^3,d4gd9<E1A3P3()#Ia1^E
(bY95_Pd>LaDX)J\XM+((@B)UQbTGYdZVB9A-P8?g]X)1]\\PbK/.?bBHTKK#)L1
0-;L#V<2X#&W4K5[Q7<51^VQYV?7.^BM-WSP5Z5WLD)0CJf.-+D/.\12&;/H3_EW
#_]P;+96BJ89)]A>3+@ZDfPaSZ-\e6T8Z)]VfR(c7V.-DI/9@AS\SM:T@.Y\<MID
(6V0G3^7+/gZe9^Ag05+[9+E;,(UEX=aY-1F1EDW6(4Z]CgKDJ\O)9DYcR^IO:HF
a,UB7N,WSKbTJg8(]J,fY=.]MAQ[FPG7dNXP45dUb)E&]U4+6O]>^_[)U/A?gU>X
E_/^>OE&17M/W,;J&Ed:@3Ib<DOXIXHb05d<TNV>Ee,Q8/f0d#E,6#I[>MHWF<Qg
JG56?]]NP-0;f266GB/YPb@NT9>/D2]A^28K64M#7:4GK24LPD+_IHC9bcO(54QG
eYN9]5Z:aZ^?@f^8e#-[:gL>GeAW4I62/-G@]Na:34@4)[WV#GNK/]P@.G:f#<#,
S2\0M:7dcZJ9R#(=JMD^Y)b(DfK;A@0A+8a<GS\A-2ZG2YC[C1X:MD;\aEHS>4Y-
]5aaf6,S8BMaPVXZg54>S?2DF0IQFdOP]3#B&HYaD]<:g^aIMCbBO@2EQMdVRQ;b
,].U5c6V3;VBK_ROXNBBDPf+abZQ8S5#7H0b,)fZ+c^BSfO^M\gEZ3M[JJP[V3\^
^ge20>=+YT/X3XTB>O7J&VZNa;[bY1O3F[)YT],FVaS0Kd.+4VRF(O9;<WE<?,Z_
D#Y9#Wbd@SdF88TI[/G>S,Ed91+K&RaC?Q^N+5+2(3)#(9ERa_-a8C57)d9=BR5e
g\(4QaLXNVAS8FW;Y&:H\Z9I][/=2I4=7b+WC&g0T/6+4dREGIc\aW4I/T?IRFW&
2+d-AA7)SL6VY2?Q>Jf91Q]Q9L(\&\Mcg,RLBZ7&9?d<0GRe/NAK<SIV;P&UeS9N
VAP;\&0+BMX(VBbeX6\[)6+850B9-KK?=0T9ZVJ_TO4UIaIPY2\5fe[M>?<aCO\9
BF#9-f\XV&DcIUG+]^/FaT\RV^&29F&[dY:,U&.=+9b&IMF^#Recb(6JIHBUg;[#
HVO6IUJ7QXd-SN6E-Tc?FfU+/J:(I<VK4VJV1B_\Ag99\4MYZ@O?YD75?a[BO00,
.9@1YSZCc9E>\U@8X#4Tg,ISMe8>_TQO:DeRABLWX0NT/U94;BE4>c3X5)D7C(M>
]\)@+L?).J>@K#0Qa.R1[VR9U9\MU2SgcJ-K(g\Z9KbPe72PYYWdZcJIed;R;\D8
^IJBg]:Z?.aHH3G?+A8OXc_-],J8@@bP:dP=fDDS+T<b,Ae:ffgWe(IE-T7]B6[b
^O[IOd:/NKMI6bQF>OOH-cDP#5U/=5KeRKP.e(?TJ5_]&(_-b;Xg-8L3?&\U53RP
f1D?Ya0GGeVG.c0GK#[,0&+.CM)_Qd6cB,#6CHe(fL;)d_0WB;]YB(&PX;6LCAbU
CF9R0:g>J)T4BY/?>BID3Tg>0Rg_[&cfC8/(ba2/].;F(KG:Tb?148(;b\^CWZcT
g18;6DEHVU#+]:-[7@6ZaLHDS?R[FI&.11A):[6CLXRQ_W_5SYeG##^a,74?I2Z#
M\MYBW81OG.N<8.?3P-H7OLGX>QYV2G(g=N>)f)bAS0bR;+;&](O,=8Md:39;Q;,
F>dd73QWY?_aZK:0NNVF--_P5^V9>2gBb]?(a;1)(C@.K:c)_,ZR7GF<>V=RUKBW
d#e3IE5Y/[_8M&^>G5eWfX?UG:3-;P]QXC@R+NRGO:V1U+W+^(gCO2>C+/)L]D]f
Q,5I(-[<>?@?S;:/9c?JSBTBN;Ya1\;8;0Sb4EPGbS^XO.R?B4Gd)BH3@Eb9;ZEG
V@04XfRTQUNQ[1OWR3D0#@)XPI=K7>aROU[7g=P<;=P]_#>]5G&3GYceFNXQ4@YE
#b(7X5N\X&GfX=DUNP9.C=CcEX<+6=)+6]AL;1Df69[)=[+J73;PYaBf@NQ9F&J(
ZeT(]2.^@e/QcTOC@HWZ0:&KVC8ICCg8JEa#ee5N98Sgb(+YTWIA_OAC.+LRWY29
RU>.B]+4GbVI<K=de=INYC+g;_..>/9OFUU[,/,MBWICNS-:5]K)#-BB2+<Z:LPP
.(fAKaP7<4-RO##.X=A1]FEf&U8Z?CQ1/Q@(N;=T;.e)L2:RD5MfYNOa_PME5DO#
O8Eg-4[F=6XE-YQ26(FTF(2]\N#]0)0Q^cg8_c/:cbP[D;_G?6e;_+4=)Fb=YJ:&
3^QaDRB8LOWa)b(b(QXI[789#SW7Y4?/>dReA^)ZXId4F)8@GU;5_T2e=SccLO?V
+^I8C^W[Y0)^.YJ5C=K4S&ISB>A7&@Ud^1^Q0C4S@+MaJCZgS&N@?c/>:SHY>L+K
+K=c=UEIa9MbTf:LNQ(RS5#E445c::FC3=T/PQWcUK]F-V##0/dQ:O,Tbd1+&,FP
ZW5[S]@24;E+>D4BfT5O5W22>79A][H2.)c7)MKMD7eLgYC4cFECEX.,X?S-=IJ0
UX[HaNGZNAg^aX1-/:16CCRG/C1-LBW32E(HV<XD]_/NLMgZKg_8D.?\cWPCXdZO
WROI3OB@2)^1U_+/-fAQgG<CVQ&P,DXdPgg^M<?LYINMHLL]0^@<bT?SaD4O7@SX
U:B)J_3++gg-_?C]^,W>BLabGd^HJI^:[5B<_)]NI>5ggCY(0VGaN#]ZY(.\5-E]
(65(eSIZb@7247,B8\TBc<GSFaX)f5@7/O_]1dUMU9S2&#8Pc-^U=C0C;_@2PW_F
dac3K>WY00=7C4V=A>9^+2_0T2eQ<Sb3S+(g0NLOSGY>G.K0^VE#&YPJcLDd<9>/
J@FSP+6JQeVOE#UUTI0SAFX2=a,Ld3FI<7g()e;1;7Y-8C)^[YQbLUP;(&&XO3c<
DJf;OfCJ4^WK]M79LaT)<+Q?.J.#LHVMWM[;#:7MPC()_OV2LSPLA0F<[e#CPTSJ
H_4fMG8Q.P?T0.-DI.X(PU#K:dCbQDHUZEcKKKf>dDdcSBR(N^cI]#P89&OGdGd/
A<5J9H=JR,Z4/^_NQ1VHI#;LIZA0/PQXE,B,IESgFSU2IFU;WOM,AJ#-[87PXSgV
#;6A\?_/OaC2]W,[G?KTAeGbI,RcCF2>HO0/SHEBVJ=GfPEa7H98aWPbc;IWF0#F
MOSYO&SX0T8W1]bK4(3+2VH;..TG<gH-4B/-_MNO>CTY;gD#La#X7H+Jaa2+fRe[
\cPZ34Lg<3Q9^3/6f=.RO1a0[6RdXU)OJYg)<H5BEN/KTD>JQXRNU_#A;LW2+DP0
YKX?-A\UV\:2K+CaM6+9>Q+f6^;YMdGLCF9Fd79=R85EH1eAW=.,H/eR-:CL@FBJ
P4@Z5gC7?=XB;McD>5W4\<JHf;C6ceNY(/[T5Qc;/QA5AW8#@#WGPW@FNJd=,G[g
cfO@ZG;@gL1c?C3^W59##,Q1,Z0)YdX^A4?[BZUUXAaD3U/fMZb71VJ(/K7Q?S>H
&)L)M#;J[:2e2706LB=beD=_/M(cA].4[a#Y,U#D7QfKO7TM[_>HARW,.7EL\P;5
S.8S+2a9-;N+-6RH&>E(#a:UFg/==^I[J>+,^^)6T(NLeY<WV5R&_f5P,G,)4-FH
2[#(T@:6DZJS3+IIW3^:@]5=[?gZ\TNXK4S^#N15DRO,\>WX_.EgL2[&\5UZ+g;K
]-N\XUP\YQUS7@I9)(YdU;G&7bHFTEGP2>YeGRKHPFI^#1Y_TdO4+3MZ3X6g8LAd
+(T1VKPK)2(O45Y>)Y-gcQ1a\8.99LU?]XYN_OCaJ5Y@M#82;HR=6=)\)^-VI46=
bDf4FdTJ>L+Ib3>][]-0HD_Y_-5E4[MdRDe</\ND@Gf,&#IJ:<W#<0[J,T?HVS@A
Re4_@:.TIa2_P7<KN:L#EWJHd9=>2P:4^3c<KKb]4aed=:VU1dBA=#S+SV1#^^gB
Q.1?W@VdbXKXaC>&bb<bXW5(CYEXHSQ9##-+cL1[9-@N4A_B+]:<RX(NQ\ZAX9_>
D6OGe;>?(/K3BFcPCY-WA@N\b=H>DgM=U1I2U=\56<,B2](I4[>4#Z.EFZ#F<BNe
ZW.cK0G#=KNcFM4R6f=UP#b@&GQL8X^LQQPgS_)b7KDY@KXdf^[ZVAgRUMC7/(^K
e2]L9@_XTW=X-Tc/PCX?9G.#g@E[8,\HVZ=7><PRKNQ\[&J_21#O+V-VV#-A:MD0
,02>XaC.UUAW3<<-R-A/.0Pec@J/2+/OJGdS@T5GI=W^:M):e=S3ZdHVAEbeI<IS
4[W,F=(D^BNZJBe>#+E-_OE2g.Z6/)Ta1OI:9+5ZT7@U3MA6M1#9BU1;&eYCQ7B.
?>;6a+Hf._#9SCIZPC^DMK&E]NT+YB^09K\.]II=7:+H=b?F#T^VFPCaM+1FIE#@
P0KQSFD=dWGC:L/GE:Re(fO9950OM2S8]K;3WAT8)[SS7e.C7KR^^,<E1J0>E3-F
(J&eM3C1>LJd&7Ng9J\Z@3\F4eS&73f,MNBDF1V[>a&MSA65a>MYCKZ[4_1U?[4)
e/E^H@B\\V3>?Q4V:KA(E4cI4?_@=HMV1I,/e/@-\]1A]BU;R&0R:4ZNT.XC7GQ(
Q1H5-[/\&R@DA0YEJKXP@25-BHE7Y2]P/eS0J7O<,1^-^HYa&@7Z)O]35?S2:Ngb
,/<E#(JEI?7COW:NGTT+G@P-FIE@I4Ze)bHK5+6_.B\QEEJN@cRHc;Q>;,:d<bV#
0^cf&D7TKI?0/;-VB_\eT.geC17Z1CN0Z8/?YA>(Y22K9\#>H.;f@J+HdPa?MN<P
4K]GD>V;WV\;LY(U-bg_2fAY/:581S?:a5gcfB.X[I3XK&<)9UJ@0/CHN.(#\GVU
a5;MNE60S4aQQSV][b99.JRBWQI6egfI=d30&Q)4Y4B68.]^>aFd82OeCH1+U+:(
da,Hd6N<]PXZcTJ:Z,b:Z/1:+P)#VAcgG4DeB?SYPQ+SBLUEBBTY53PUUHLR2.2:
:)@He?)dHS=H?8FAN>_^JU>WOA^a+F[WF@VQ0^8=A5P13c@+OZX2WA<4K7[[c=VP
G33+3[HE2C:--bV_N(OOWXP0cA+X6D+X+e<+L?:5ePVOI+-//(Pd;TaGfOB,X\XK
e)=D.G86_2V[HDB/FT]^K&^>)3?\.bZg>0D<.>O&^3K/^S[ZJ]?K&=Pa>8<7UF]4
L2G&65Xa4Oa2=:bMAf_abU[6GgN-F(aM:TV287-,52=dK/J)#<d<O)e96DONZP7R
Y8cDAR\[dF,,/)0/@fNFBGHYc)Cgd8QL3W3&:VD+3G\5M:dMRQc,IRC@^/V/=UKC
aWaLEW&J(c+.RfD+L]G=2JgPOQKdK@c,+&_VN8V9=VXN162NFD;>H=cK:7R94[HQ
_ZR)N4<MUMgb@(WADb83^7=2(@CLBcM6EE4U3[Y=2SGc(Sa9GM^OT)Rd6Z39bY>T
69S,,[-T]EJ:NMJ,#GJe\_Y,5P8N(]7T:1/=<.,CND-&;JG?Z8JH90T3;E24.=4/
UWZ0=7BA=4CEQIXNLe2gU[H]TF7#/S5N6e)eJ<,&83]J]5PbOI&(1V_0CSW(/Z;O
@ZEUe#;&XI\_4+,VHHJ05&W-B74194?X;cH;K)HdQWg<F=(>ASE[M3++O[DDJI^T
T7Q&@C:T#5fdg]0,X?2-]/5[K<JIQJ#G>P6]<><+ON[/.f5a^VS?#)D01-aSMJ2d
8R?HX^XaM<I.fCH1,T2QaFfNI87YO6_-HDCS&]Z(e_]e.Y-XW.]R1bHCBYG6))A?
&6,^;NP?(EP:a2@=DI^FaQD^9=?I:8HQPC2aXaVWY[d/[3BU:c(<d2)5==A#<,d\
QgF-I6\GE&L09G=c_7^aSDd(^_UM(cA\)Fb[ZDB\PZ3R.<5WJ_4&&.+-2fIbW\F/
>V+>dQ8f(=XGXa=VJHaU;Y&@5a&-Va6fG,TU0RLJgGJ@c:B(SH=M<((bbbdVTD1E
dgS/aN#6)KgC:6H+ZbKNUb__eIc&X)U9,]7dN.7IT3,5@L6DZfHS,gT(5RO3_2gA
=e@U78A>N51YSK)Y/L5.(K/]MC(\(cN^gJ@.LAfG2Qc4HA>^O?+#YA6d.MgaDIV0
A)6G)W8d6&RgR:(69bD&g.cKYUA0:0+YI<@=C9CT\.#DdM0=eWR:<8a>X<[3[8:_
C&P-UNS)S5=;WP85WHEOe=Z>/f<\BZdZ+:BfZc5H6>AVJVQ9U.XRPZTd3JWS7ZWc
2b(8JDR^bbbcbD6@RIG\E]:_?L@QAef51V[.,Hf&:M(]A3Z3?>-WR^TF.Og&^b\:
ReV&L[9c(gd,8;RBYXXb1;)X5PW+4HVF];U+9F/fJB)TXV[+IMdfY_V](Q4aZMO[
^I3-DS=R^FTfB,XB75Rd[R9X[.bK/M&6WS,a);RR?Q4Fa)F<:8aFG^0#S^e>>)0T
5+9b&3009a^(@[>D_T&A@R=W]:&Og).cWBA0R9SD8QD7c;-OF=e3?MDB5<g@-f;:
f?09.6+#=[=E+\BD-3K,g>#>,&a?7Y3-JV-RJ#WN4V[X>?957=/<7RE9NGP/fUO#
FAX=\#U-\)FV#0-R?CLUM:L??a6OE_5,Z1GBEbMd\cde/8OM9-ZLPVF?;Z1WLRB(
\b)]dR3MN:+FYH(0)c@0Aa(a\_.fDRHU\+-]@3;<(a@8H=#AB/J[E<;b^\]E:;_J
;GPeEHPO:^>gOO3NH+9=..K6-VAaJNX?9[[SX.(/</__5_7GRKe;>X(U7a4fU,9.
9I1[2Hb,Q<-S/DNb9[2+Y;IEROMAZWM_JM2B(-;e#41U38eF)F\A7U95ecFEfNEK
DF1f&41,XHT9?I-OWZ5.TMVgUWV=ggWVGM1A=241VIHaW]&OfAfG-HFd2^MUV3&P
?R&#\,eI[?cTMd:^,QTT9RU7\O\(=3HcI)Y5/3M@3YF6S44?@<LN^OLW;\V2>D+0
EXUbJX9RaNOR<TIGT2c=K-21^0IPcCS33,KGP=E4K>=J]9_73RAeHF].0-QBPI&H
@fC:gW?CLUK?JeQP4N4G&7#_1aHg[ef;,LcT?\/[YZJEG)UF>Ac,?^I3+_d[E6)J
Kd4P68#SUW@+:4(.7]Q6L3.>_\8/T8a.I0Z.AA-B=2FTFXL;WQg1AT3]L)H;W>42
05]T1X1e2g747+:0_V,F8@79(9d1)77QX0=+:=S06a0Fb&A_)8V(EbG--4IG^#fM
KY3cNA2)La&]95+)M97[30F^4(TB[LYg]^:f5TZ?f#[7KLeX/J;(C/6:-Q[5A2G4
?P^?A]6J[Z4KeA@5HJ2@IC]>6K8-P(Ef;9?M:#NcB5D./_C;D<EDWd7dKQN9Q&61
.KR9If)C8X;1/5;fMQR@1g-8\L5KD9a2#6NgC(6/^<AZH-<9a&&F@g(aO-?X/eAB
OJ;3W1G;6I1=e(TJQT/VDZ>Pc3L^0:PIDR)/f8Kd1;[K&1[7G_-);5X87X6()+A]
W]V<T)6APEa#d46J#Igd?_1)11b0<g&Y>3AU5XW^NDFA6]ZCC?EbNG30\Da9b21,
Fd8T:IMF2bM9O;<&,B#G@=0I6=GN_;7:U=JA\@O5^[cA5(V+ME__)35HI<Wg==2M
T-;=Wdb]:.VaD92_f6-P^JW9f6S,.BH::gKfB&J8#SgTR1OBE9=R5.(#BIIGD2]W
eW-#G,K8&Z&DJdMF=aQV#>Af5=KJINd+>bY=U_BTNR9BAXDNG^TS/fKeDBRGZI=W
A7.Y8429_dU)7IM5R2226+Z<Y(I.BPCG;6#dL[GKFb4+FANO?DIFKfAJXWB),I#E
;]G(>_2?fVEaBADS18A2?XN=\^@HDa0BCX8^W3G_Bd_MJ/JKHa5HE-L#XZ5U=JK2
R&BQ&PL2GOI26SPJS/f:)>SKg#]=(H1J=^3OFU9GdZRDE;4+99(bJ2CUR5[L[MM5
#UT4@J\-DYX=g_@>eW+8bfQER[4UP3ea@QF]TP:(G\5/d/1,4#7H]PC;5Fb:@g2L
Sd?^H-K;Tf,M?\U>)=f79Z/Z;)HbS1)>)5^GXK]0\S_YS6[DH[Y0[=d+LO8KS>Sf
1\J;Y5.cH=XU1If9dH\eEWe+=)WRMPK@<J2:YIf905G<::3QeG/KV1_ec6FK=6d\
L?@9EEPS.B>Q,N&BgV-b6MU[f=4D6U4QT3BQI.LaGMR=^C=<Z@VNf&+RF(6TZ9;B
[We5^0XSeO7#Bc?=NN=G.RG?[g,(79LKJ(&F/K5C<+#\[V1/gYVZI3]Q12YD4PAN
J#?#3_WM#1E\(#0;LaRK:+IBRLeaH>cV)Af;a1URGeC=:g-9RCXC_,a+:6fW^71;
;2gZY;fO,I.dSKPRO_.eMIf&Z.4-@.^345==3dEf48a1QH>6TKR8_=R@,@\aB/=\
UZU#\W)9^3U8#Xd@6KeNXQP/OSQb4ZC[J?EHM^a:4UM@F-b^NA75/#L^Z9],/(83
3(J4(0FTSg4b-D5BOT5f6>X[D;.K<1JeSP;3S7Q8<7gIQU/=DPI9c_(^,N<],[S+
ES]>MV\Q(cPL9@XQ@#BedGeZ/:N93bG;E_.,+/-PgD+e.W0<R.U>M(\a<JBZNS@N
_[]a#7S\8]_Z@fH@;6)IGXJ5Cg\^SB7VZ^gARcDW8W]CgLS(b;M38:2Wc.@[SA61
_[(J#F_;d0MXb<UM>8VL@G2-adcT3E(_PC.-+dbAI^W\5Q8#AE;L?1)BXG/;[J_:
-B+G:2(Va/;8][<:CDJ,?dd\./K\E[7=R<7fTO&()-<M17VJPLXF21=0@:+DC3)8
4]AM].YY^MOWDFbUEc4LJ#7P5Rd@I-eg9_:/)>CPW,8SN0a?#X?gY3cCTNI>=5E+
W]0SN;,5b.4@PB(MBUK;N1&YEAKdQ=8W;I76P#X]3IQV]3.9:/+&a]\K8VY+d93J
K\e8K-5)C)[F:g<.b\]g=F)CQLM2A(5U7;Yd1W,g#/Q;_2F:RHcALX=dC#E91P[A
PC&XZM/\&Y6?OYd932>>:MYXLTEEHfd/C76=#gX\Z-LL80[SC8c3Z/S>9XPP9GY6
<@6^V_NAd:A]+P2?(9YQ95V+fES.@0C@^O>;E1O+_EW;=>Xg\V,A8A196W<2B\eW
@VVOHE1+,W6,_:.c:\A3E:&QZOHB.E_(TQC2Xe^N2-U#caL(I?=FMH/&:UZQRO;f
(TSf83Y[07AZ;1LQ_J[KGF3)KX(8LTQZddB88IYK0@4WN1&OHEK+_?4V<<QKJcNZ
AF=,LLNXMZD7&R#c^R;Y8b=H)aXHYRND(c]b[6N:HS?B(>\Hb?G0=g7=#]84Y_E+
M(04XKSe:aCO[<2^[V71_4bTg>#2aCJMA7PIL_ZG-dIYNQ+-fP+\9Q.@[/\9F^:@
V^e+@8bdDGN0G5EXa17CM.B<<K5IcY\e3>C7]:1FS&a[?,Q)YbE,fDM-P,JFJ(#&
<;d<fb#-.K;-(.-IE39V(IWF8]HW,8LTN#66<17LV>O1+YVP@C-C@BdR+c(L2OPZ
R95?;La5)5FRRVS#1X&W;&I>D^HUN2E>B@&Od^>&H/-#K(S=940^>P/:F,<;94S.
<d1?50;KF+XeX1>+(;,GgO?d7E)),<X.Q)NWDKL_=.>9<QP)M/7=&2TRc4PK#SXE
_bc+ec&OPPV6[TN;P7>40?FOI;M(MRT17;&Z9JH^Ue3(52N<MMFd>@<T<cI3O^FB
)ZZ_;-CgPA39U-=BA?S:MUa2/WP7J:RN1>b2@X:C,gP@]EIC=3/QYG+5\3UJ/<ZC
(58,E=]VTa),.A/G@F<G@VN5@e79O+E:2aI:H][R+g9UT1UE_G4WQ);/@98M&LcA
0J:#4Q6VGCgd/R\C,AL(HR/EdP4(T3C656U^(W3I953W6>gB2I.D2:7BeS3::M@\
6TM(g.K<d]f&8cEc9L-c=50I9T(#?XJR?-PCb70:Z:22\D=IPLG)X&D8V2E>f7B]
J9AHfN,EMI<_K#6=(X174eDY19?G\=Wg>gQLUK9RPMX3TKacadM;9;<45[H-OG0.
)]//JcOX^#3H\)6,5GCR[N;b/,d>7#M6.dfA,EBT+>TaX,HQK3ea#1F/F_FKPU32
TOIYJd#P4-),6#_;>@PO@]Sg(U=6M)&^Y/8G6.ERQG-+E6_JRX1e,;MET,C@4fIR
gX=:LZUb_^A36g]/).1-(V;C]+:TD(7gDc>+8R>BcEGg=aZaaCYZcT4CH=5A>R3Q
(:d.5a1\6]:_&V^gO^8TK^0;eV#PKF(-&Z5+)18>_=-agaTeBRgS07g(FB)+F_16
6VXHD_QE9fb>Cc8(YAbUX=d&+N_cYFbB)Y&g-]YXI=D6@,YZIR\Be@TVg+2cQL//
W=?[RAW]DD].P(M?U4VWS-;)[1cW2#UBTQPX&[Y(R33RNJB=<T&&=/L:7<60P^T_
6Ta#/a<N7M=f>33D.?F)\e)@S4(I=9T^76dS.5=Tf5Ve^<PD>fS^]J.4S<K5T2Q0
/8]<]&I18Lc2f8aOFfa>KB]6HS5/GWY:#7&[<0Q-9e&RJ&ce9YC+9(@RUQ(Z[4]\
K6c20H\E/GY,9[bTXb4e:,)1JCZ<E@518]+D.-@]369N\&Ng)8[QK(.=gSGA4V9F
C457A3X,C_K9HZ64@W9S)\Y2_&N(OH<HdF7Z06=M)V;C^O_eR^c:&/:J:-^;,[gT
_U8aZaC=TIUU-)7#XNH]&5_W=K6bB3.aB+8J?+)8@L9X-5dVUN89gKUJ?[Qbd#:J
]T3ZL:<LTI-ID:^X=g,7CRf-H7X1F10_0.c.HQK>.:1R1fCQeP?TeL\2@S[OI6-V
O\).TS[W/f6+4V01TCL(eAcgHG92Q61[;BCX:PRY8JLB8Q[.d58:W3,+fcV)UMR<
T^JPA@?QF,>,ceDAd8dNO,UHTYa</\98Jg+:#97AdfCa&_KNEHDIB-P71R3YeBM^
#g^_MI:.+:ED]=<==ZG9eVdReSL:0(@P7\JS>XPAPKf4]A?A)4?KZa&QY#4.g(M)
LE+/X6/])-#[W;6J2U-@,^1Ye>\0ZTW)aCPF5Z,R1.)7>D_g)eH2&E7URCAR/QG?
M5Cca7_@&.c40S#IQIPb\+S\MBKJ>\DdN@gbe:?cV+RfSg7I@??,;RT?F?1e\4=C
3^aIQ4ZZE2+\2)3DT(J9f5DSdV2S[b#dLDC=VDH2/>^d_b(E#4&/,a<:SUDXf9<4
2;N9a)5:Qb6UFed97=7]_b78DKG8IZW/(6=@D8QOe^W_H\fVQ.I>M&B?,+a#?^9]
O[:)OL)fae]g:WF7AAa2?9Ea/6YJ5UN<6=HGG47ebOJ0Va<B7WF8Z;NDd);Fa]5L
]&WIFb1H&g0,W&7;IXA4/egYU5/]?.-2Z:4W\,9e;<P46O(OCZCb([Y^Y3\9=8>Y
PVU-^M97MG\Wf;==<N-I3:aQB=?NBQZ0UO)K3AI8[eZ>8LY/EXU7E&54LD&23:cM
P@NV@^P553eI0J+A>LJ<a^7R:,Ua+O)-c^P-36.QfN\?Fe1-H9_[)g,L(,1QFa<5
,e>-SC3@M#61D+aVHTH,Ha;4G)gEAXAVMH_^a)=&RGWS^P7)VG[ebM9_0M)E<MR:
D?I/2VS#]UNWTYLaS=JcaHJbN,)dc,F-LTPd+OW_Bdb7,GNaIYEKWJ4Mb/:]OE(H
SUP=#?>JXWQEd7SBYeT)6KaNL4P-S.EU^V6H>.fV@Y/<CZe>.0=E_O<.G)I2ZY)_
Q8-9)6cK#cK?<LJ)KZUCPIcbKIJGV.16#dY@]/=];1L7VMG4YNa=E-92Z(bH,BI_
/W5_^6?FBG5R^G4ZX#?UgVeK<3QGF:N(?(9KCL&8W-d8,BdJC)4@MG@@S@Mg1L(f
V-:@CbQf9^5[_C^?P^N3;2X==6K3.UG@ADJ>e@Hf\c+E?5]Re7@RS315O<2.,,#W
QL\X]B[K[X>egB-\T;fM#U<3R8Ba0X.^PK5-(NE(2G.c8..[N4R;,82e^5Z6_1H4
YF2<2HCJF71)L2a/H:)&U1V64/X-1U\6aRW<@Y\S_aP,Nd^\@P0#V:fcKDBFCB\C
&gMY[IFS^AF;OaUZF1K7U<<=&L+9_)W8\(b6F@9[VZDKE10@LNS_?[>.DaS66^O[
gJ@?G3=_8]1S_PcXW]HA=SRd_cb4;FXAe^))>cQ>N\@&OKNf;3Hf<5XdEH_J/Vd5
YVR<7?,CcK-N#a\/Ke.VD0>O4Y;.X_D05D=<:48AF\O)+g7S?.fJ5W3+<ZJ/L;@@
&g8X\:+HcdDdfRSHfP89^GG]#2]A)BG[L>YZ6\_0C(JB:JUIKPB_FHH@4+7XLU)#
Q^;[J[(@gW:DEM>YQ@VETN),EHF=SGY]VMU:1P1B(JO.[BH0ZPB7;SWLDC,7@+[L
.[FS>B9F;(_aIe;c;G&/fY0EK=g3FBIKAI7/0Q9;J-+5C>11KJSAD5V]4W:]H/@f
KdG=cI#;1FX/8H3&I6bJQ-0IH>^5FP:aQ7PU5=(_d3KWWRGH[1W(G(R\/dVBL=4)
9G#2<(/1_HVaf,X0SBR?f;85NK4+J6@N4cWCTHN?g:Y&Pa6/I#];dGPG9KbB(-ZL
Y<9O@2=)O62Q[UPQRb6F(F5[G?GB=W\>C.+UJG5@-J/]Y8b=A0OEe050J+dQOG,U
G9:WOc]Of#CY:cBOIe54HHR[-0\1Z76Qf]La)HP\I_CEYTf]1d>CTDN;e]0+B8gF
3EYdBB>MYX..^&@\_<O5J5UA-R@[P>57G7H@PV4Gd_+_7)\1E[b9I:ag8.b9.2U5
fV/44ZHU7@REEKT@^d/:c6e.&QA;e<O6LN\;PK]fQ#C1WYa@_R?.N6>NIT\X1/U^
YaRW8+PbR>OU_U2[DQ<XIN2A&#+3PU&W_1(^ePY8V;S_YS-;L#EBA-&PA_9H3X4(
WBS4>P]K_2TWNRSMfb#YGKA:gbRc<2XI]Kg^(#eNI@&3@Zf+ZM[RE12^]6[ae5HZ
0<b@Y=LP2UJ)<5W3,^3f4BPB-5-05Ab>=098[YG;I#@]H,#5#(Bd/VWOZQ,XC[O9
#GZ.U4>?/UJeJUb_MeXC@O^:).2bbb.FGS(1U<>;_CGMPA\D+b\90X>gZ.La]#_a
_9GEVDW/c;9J6@0,e53E6G46f_8^8+7DS(LD1cc6YQTaU?(\?(MR[_[C/\b=7CUD
6CEOB2\[]Hcf-U(EfM6[<DD8?ZbdH_TZbb[>=2R(ca&JSeXEDZd;N01)U[Q\_f:_
\V&7K1T5gI+agaHF_;5:UDHU5E\81c96B>b+)8_TK1AGW(+<dY8&N::^L?\_PdO^
:K:#O.#4@89#=:N55^e^,bgIfNOH+;YT)=P((?Q,V+7;]32;>#8Y5g]c3LAUJ<Y;
KgI&0+@5::.c#9?M-8d.UZ<O>K?7bWCR^2CSd/D/6LPM4aHT:I(b[GREaIP\JJ/;
\dM9Oc\(6OYOa4:eUAb#8?)cBd]7R\9SJ_X@A^Z@AfV-#Z@,K]F^1+B@Wc@T6V+/
(c-]+TJ/dH)?)?ZOQL]fEIYY>e6C)#@YAC]gDT/P&E8\21S,cU@8Zb^HRM0N-CZ:
cf-XXIRF5K4WCfSS7IR5^,]VV<@Q#S<:FF3^/&bOY_1IO93U3]T^eW&L>;BU0K;D
f977I@3a7RPR&)V#]5gV4dGMVg<@#gHUR3LT^5MBP;R^[/[&-_7(f\YS#FWGe/W&
9V&1fY#8AUg]Sc-KKD&.Y?_M\#c<V<a=K3?J?<^g9:_8;&DW.X-7:3/bS)FOe=:_
J3/3aCR\b:W.R4SDZB@]T7I)4UGfP4NIS,I^A1CAR[0([CKa[9/#&g5B-?>L]b3T
5@Y9U//P,G:>7YVbG,T(V5Y3TfYG-HKU7^570.Y=J.b?@7?+X250G5,6:5T;U@XS
.U0\e.5F1S1:QHNcR2_BKW#6@[<,eEe\\T/;DK67+3RS5_TT<-c1&:GW8<FN^W1:
RAE2f7V/1[:69^C;;aLTDH[eDTP3@J@Q>;9RU[^G;B-M9D3[0]]IFNdASf@3/Fa-
H64Nab\]aU..9W9\N<R+Z0U:8+B-&d1^a:&?)-R-6gbI]ZbR&Z3Q+3Y7C#134;.c
Z0=S&6OK_E5B)GE<DJP=QB5=QAc4HK<@7a&I\.bP-W,1+]K_E\0AZ<CUSZFERDQ/
Pc8)LNb9]XRN[H-1E?,5\6K)]f/K>_CK^LMZY:2C>Cf:(/Rf7b8T3RLL.,LDN_6/
d/,/9RGP(+_Zf[[>8F)6S[XSWeIEfD&.);Q2e&P^KKQYQ@=UL?N>Jc]@2/)Eg?ag
X,WdNae6UE?^\eZ8QTFTCXVdMNOAaEJPZH93E,]&U9;JLLRaGB<3GU-3[-AF;[L\
?EHJ@CNQ0?F?,_D2+da5).;TEBe94JP)/M)K.If],JCVC9</BU5Z;aASGAU8)M8>
2>]V>J8<ff>BdZJP;L(&?Bb?beW27gL/.N51=^BN<ZB2GS_0S.[&]A>&]f3YA)/F
4M(T;A16U)T@?SBDI01RHVQbRZVK0-3>C(]PgYUUUGB.=X8J@._2K2N?OS<N=F0Q
]Dbe@^YYXDL=5bAGA_->Z(?8/&Y6[ZG3J;L.P23RI7B3dga#(b?5_?N)c#^IV;>M
Pagb#.JLHYJ2X0](A[8547@DNJAQKRFdO-/YNU,Z9Q-HXC:.\EKYgU=PUJVF=CF0
]OWMCd6[[3KB&1c\FPe[ePBK&b^[KN^T2AKfQ9Nf[ZR38;/(+L^0[afL=K\?MU9D
LgCP9?4bL[-;(gZb+,N?K(cYOZ/f^@bHdEg=0&?H)d,@L1OK.H-<PcKg.]Nbg(67
L7[-Dc(M>eH@?Q@_20>7,0DZP?-gT#>gbeZ5_TDM\[\Sg9<(+Md30#?66^\FNK74
@,;WO[a4VHS(/^6J-K]HS_)_@gA-[c+2@)-AcP]b#1f^Jd@I36)ga\P.Re13@]4^
gfRN]_F+E<]1X:H]^J1SG)T1-/519?68\5f5K)6(S8T9^T(M_4<Gd5CE5+JbORTX
[\S3WF-e#F=DTRXQ@##8:#D)U#>@@J#.6#]ZW07;JA8-CNJgS3E5:@BCGL&XW]0[
#6E;W7II^HQ.M&]P@L\NT1@6g-PG-BgW2XA=R/6+>Q^4fI8<HC\#I;H;14R;SQHF
CG[>ZX]W@T4^^HVWHJc=f2SARPQgOIe1/e:^(f&(L>,.I5bc\VB[?ee=J]?0NbS]
,Ag390](J).F#1__O9NeU@H@3aL&6[?7bVDA:.E3DJ91@_;]b_:3c/-KA<.:1&e8
W.FSMMF58gA4#@+?>L#><G1P[_WVW(aO2)>&<KJRS?+,<I=P&^,Y1?\F+#7S:+I&
NW[0U^,Mf9&5L+KC@\fHO^S;[RJP-W)R24ZM?E5W^\=41AKdGP=E489W_C&4K0Qg
gQ@Q:S,X;+L5/2YFS706JX8@gYVg1G?&G3Q0U=K;cPU?-T6[+3Q0g<(Q(TbP./4=
d5eB1Y[STHYK:\@Ve(KD[8M&/3\^S+Bg@\L8b=I()[CTS3TWV^/g+1,0:(7cI)XH
+7UUS+O2:^eR=Hd)A[dQ?FV5:.TRPT34bX-H1aVa_SI]D,H>b4,:A;@SH\<J&fUF
JXCL-G>d=O>UT[R^2f7#9LZ__/E?F@]&5DK]5&DU1eHLgN&HOEeBb0>fgSR80b\5
A[VWe)N3HC/+VJEbWV2[JOTXVKLGF(+c[6Vg.;Rb]9G.EMG;4Y@DBQg7X176Ve\,
]^71]T5+KdFA6aWWX]E##@baaBc5ED?9bG:Xf#U@1II95;FJKKfK\UG^e58a.R9<
86ZH1\S37<6:IH.YIaX=9K>BRZ4bH(8@:7B>N&dZaO+:PHL(8;P]KA85LV<;K75-
c.;J7>:KYG?5g4g_,E12?LG<0KOGA9NVQSSZ;#c>#Z?-RQ/)&9CK?Vc7EWE(7GV>
#&d\.4/R#g-\TFP<_c.Z;57fPdZV6f2b9Gb-.?;7LTL,WN44H:N=bZc6>154YB):
(5=J<7FNN,IL#>SL#e;@P6YfeYCN^L7ICMSe8SQdc>^Og4,04ZYB9HfV[-#H>6XF
(WdT4dF3/#>[-B;0X+dPb,2T:FMP2FZ<][9<.Je_RX96ad&<5\=5^)]PgJ0QE72<
),&&MaX3C01EBO^\SI?9O&O-1_<1O8L\ZBH;-V5#d9Sca<N,dJEO?:).)126ZH^7
g\<\,HX/2L8ca]#WfB5JgLbg=H2JKI2@Xeb0cg:N^37((#UA<<.;>YS-<e9_>BRE
1.P/NQ)g0]_D\)?<-=,Q1?@&X=b5@3\gbL3Y3Cf(P)?WPV3^D(fX@dPQff.MS?EF
G2cA_&0U9c:#75Y0HH19XI[Ub<b1QH4Q9Gf,BC&+:e4]@>OC?f;Ngg[Q@@)Vb?L<
>gXX6G+9&/HXU^2_9_HgeF6J3KE8ELEN&ZU]=GZ6_1Q(OEf7>JgSX>MdSa129cG:
YN.2b^gBF7SYIHbg/)M6Y.V:-f4PLbL&f;=ebA)K-d.eCD41O1O>@7\c\L-\IX.Q
@gQV^3HaKUJNY95KM_9fd\1J_;QT1.>(g;/JHK<QMCXO:Sa\fg3g\\V4R6[AcQ@<
A8E#c3\BPF#<b<U7/F[EWP,aHBYRNJJE]=NO6D1,E9D&L[DBL99(>.S.Ad2,L?K:
:cE;R@)eHD+_ZJ<Q/>gL1OPY(Ga+SWM.(;4Z?MdR6VS?2LX]ZJ(P&6YURNG=H=&>
:F63P2F3GgM45A,4FB0RXMB:&-OZ9W9J\6LKP:5+C&&eA,:4_cW7@=@T2PU:@c<d
Y79TGF=bL5K,SIV\W#V0XW@G5K@2c3)F4c?aL.\/J8e2JJE@?^Q0MUgS<ZPfTa.^
8],I\B2;(VF##^.D+ZTe+.7O-e)[/Z[#_e79eN(U:;8[^Q]-=M7c]+4AL)HdUZO[
,E]e]L85GH0K@79A]CZ1=+X/>U:L_MN15.0B=5RTW1-,R^A1cXSOK[&E3K9/G4@c
-a];5W?4D=_aWBAHH,WF799J_-b_^HF@53,TeeSHe>WEWg?9=af<?K2)TNE:#@.,
D;LF;T,E;VREI5F5-QN^E)gZVaPXJGG8[QdW\,5X-T>@V5:_GPTYRAZ.W5S11B;/
VK]6)@DXA5QNb)db2gE=;H0E:f@d=F4AGFcbQb9UOO=YOIW\=GVaRbF]0#[K^MX:
\g^61&NY2&O\FGSBc@#?BH:22BbVO5gVO,4IW9AD2T)<G]J3ES^eK=AJ,4O/+)P?
COW(X/69G5M.>cRDZ.g<;Y(^QfHe1SQE5E-MVDaS[>]&fAP6[N/5R?MZA50F.b4V
<ZVN](7F^FF.=,9C6K/_2B)WabM?)E=Q8,PKDZB2[VHA#+Xe=X^gfId3.WZ1G#5d
IZW1A0/Ic;e1X273R+[DcM#Oc::FUD#d#fCUVR0R]Bg?YNH<B^#58a?@C8QTA5VQ
NS3NO-;UY^?4g#^BTF3I8.R[LW7(>beaZV?[C14(<_a@5\d[FUQ?:&9G(&S8(3RZ
>MM_C0/e->WRP^VXCNNK_U6?;_3BNR(O5[T:OfZZ=D6J-ZK2<ecH&SH>F.2-a6Y0
CBFb(P_KH^Y#S3^>HgL[--M>?@a;V\O5V,YOX=LfRH)T,OA7<MCB23e5RH2+Ze@Y
9fR^/:f4g5EfZ5+E8BfS_Q;<LH6VWeK8R9SC65D1cVa;KXNPcH#Vb>HI:[<JOFg@
DLO[:V9=F+\N0]2\MeUW:^R@4>D0]WH]:X16JR5XSY&OOKdL:3JbY_cU(13M03Ge
fT#+S+L-R,DK8b:Z]#;/IddE:62_T+-P&G@<&>KP\NL[QQ,46FbK+Q[g)dK=b<;<
G=.U&,6YZLZVa#8F(,5YJ>7HF59<+@&=V<YRZ9aI_\C0D<()FL7:@J2[c_d9.W\F
BKW,DF4WaK_7W)(JV=QA#A4IbV;IA?SA@\&ICRCA?-4C[JSPH4)9aXf=JA]_GfdU
4_g6=P_&X4G7E]XK4K[ZK,CW)SD6<A]d):4-<AZ0UJ@;Q19OP/8cP=RC98#YM3PY
c-E2UYP6_UC4-Dbc>\/EIEQ[T_/J8g^Q7S,4IPaI9B^H0Y8^VLB=0d^B]QM+KMcA
H@V6<CV=FZ>>TB=.)CWGZ7E^3ZXZ18^Y(?4<]_=\8VR.O7GM9[SA[(1CdF&3gAc/
5c_VYIK)Ge2TSSHaRMEKLPMH&N6ZGZ(/d\b(V\H:X4b5GFS]?[eZMcaS-5_a]aRM
#Q02XZRJVS:D]R#^K>@B\.H:5f_d,UUYE>4^fd:>,Z:5;g5#MFLO[d7B2:f\;UTN
6/47G.a7&ZP<8CQMQBM2N0;&4:O\VQgJB4LC(R3]&>.Z9]1HgfLUA&IIbD[]Ef;b
eTDQNUSSV74RX4T4f&AKOe.65aCLS+Z>(58+A2G9^85F[e7TO.-@)OE,DD4).8^I
^21P=aQ.N=GZ[81ZJ9eAGC9@<[[S?RUBbg_]I3bZ:/g+J=;)68]2<<D7Q45Y33U.
0LMCV=[<a91823/M65e3_\H)cKQ,d-\S_U3Zg5fF7?CbD=1_+1]@A/LP1[E5Y5L9
1SAddJdF-./8C,>UU\#3Sf63#cZP^g?N?EHL?3Q(LU)IVcP0[:IXMXM_-^\.H\IU
I_FPJ]C6VO5QCI#O(+@)4UGOL8,VHJW#f5J/b94HB2+96#6@9g?>e5fc23;f7@5S
TC:SM@Z)JEe8+GKKB(](Eb+O:K5NA>E[cOJ:V(8->6eaQDY+;WC]Nb@D6Y=M2#b-
[:+:Ee#.+S:[8R^W0F8C?#0#d78;R<AYU_cMdb(?-g)\8,\.Y\BR@gKH1H9/Taa]
I25L_RSKcM9)[0TE>TC9D.KgTgZ,73RCS6HSE:,OTSNgWC/;UMTOT3R#U(N8IU#<
/=DD9SI2,^\)XIg6TZa[]46afLCgN)+,aM-UEFTbgC@@F]&A&R;DBCg&5,69/(TZ
RXD<f:e1KI@AgZ&_QSg@;N>V(NOe2T<.=g/(BXYEWLRUKF/]2[=PKHe:S?RX\_IG
A=C0;C@1/HM=d8@A,Cg;#SfAd\XCbC3HZ6XX-G9\ULF0(L8]XD.L;09[>RBMN?PR
>ILI,8CPde;F,#g9@LESd5S]Ec0@.T:U?L_/N^V7Ha6F;+;0/aAL+_X7^T:K?C:-
#(B?f^BF=;KB](>KP&=:D2;eI<=^f@)&U8,@f1)bFb0F6PF#TX(XSJK,aW2[L/MM
?>R7;\H3Qa^gKG5:+BE/5fZRe->&5+24T-b,6CCX/A\VY#Q.1C>_-c6T5L7SW>?0
<#()9==,6HOc&57+Q>&8aW-DE+ZQ7.ZOZ]&=@FO0ORDg\E[;@GAAUaAe3cQ1+X_[
XY#b\E\Nd#87<408F?982<B3+H<(]MO^7N([UG/1@bPCX=?3-#SbG-a=NYHN6WeM
cR<&R]dBT8Q]VLg4d-:=;T2)EVVd9/+<@aJ8[5D<+#AJ5IT;@F6aHdQ+X@DP>d(P
\40Tc_b5<f9E]??fT>H-C[WH5\H]8(U)[]]6gO@dU;9.F&HHcON3#I/?]+8Y7VIe
IgGP[F?@/EZ_ZC4]P9fPM4(>;2E0(NR&)IP@40BOC4J^bR,cKZPB3@O-E;NQJ;OA
:WIB<+=<[Ue]+\M?=]K.C;Ng#8a245.GA&RP9=.?[<+\XU:618[fFF.cCfWD-8=d
LR,<LdT,APFEad\8_.+[5=\0RZf0/0GL8.M#?9CEA(,H\FJC&,Z<^Cb9e2_G33&<
_fOF&/-9aAUWf#QMTK,Z71^EHLN@XBBKN[SDJ9]cdf?6310(X,V56.dDB9Dg8f^^
I=-/;&;H2.KcfXc8;)?/WK8O(7DYE>HFc@C+C(C,W862,NF^-EbeS&+F8GIW3^XZ
4>-dZ75-U>^=+/9bEWbPYWeG=EAD6C/+;C=35bI:V;ZJI9de0RGJP^MaKJI9E&-d
K.UGXfc)6f(<YBU.B\7ADZ.YO772EN5B_>]AES0@g]9a[a.VcP1\1XFa8@2F,,4^
BeIQ+4(WHP.aB0&#O_@3FL9W9OMa75D9NZ3CX<TSc/#7G[5cXU.W>0;bCfYUE>@T
7-_E.TG,9JYKAI6HX,D7O./8)J_G]<g=NAKQYO0cIE4&bK(>XG;\3&+]V?DL8[5#
JBD\6@gWMFe,;ZQSfC9RP?5C<V0@WC^L0-Y,U>@1G?IQ#deMdPa,40b7XG=B>Z6T
eRO25+WSF.#[:VAQJM1cR3Z<I<;9bKOYHY?E3\RX/M4W;8#+<0=#^T6LJX[AVGTD
a[Mgfg/H&7OPW>H9RO1V=b4G<1;TG,0Na(ZO2QJc,AUJX2MIg,K-4)VL:&1D3d4,
@\@6UUG8Z2RA#b.SJ[:eW[GZ>Za)+g6ASUO,g0BA84@BC<F5^W[]<MP>0PV_B0JL
<O5Tg4b_=(C=\8FfD;9\R9\H-A2SAVCUA^1\9X:Q3eJ2\(=\bZ07_#7IeY^TcBeO
D)_,V<3BP#ScC.a\7X5Q9@E0fC+^g>Z?e#F2^A<K9CEDM(cGWZIg^,,3_3da9YU:
<Q(&8Q9bfeJ2b;HC&<>;eQRVFO(cZ=6UTX4eB_\K&DXK5A=f:RC6RV?/A=((U>KS
@&A2+)M8cB)RCE4.\5UB:H0(MND9A1:@TAKBZTd0Q[42&@+(,P:0C<9UD2dS;60+
C&TL(02Afb2<E-/[C_gZJ.:#TR.^;31\cM6d\YN(e34TT7TQ9,cLfaMZ_d9aZPA(
a]:Q>+Mc0OMEZ#ENI6J/);Y4;XeQPU/(;78MCU.KbgQ+R3O)&YA_P^RX&@NZ6MN)
W2>Z\.>#U9/JbPFBYT<(S;ZMC#G7P:26d9^TB0P<-:f.gc(KecDJ?.OWI+)Tb,SS
&e4-99Z&1O8(fY9fV((DOYg>eE,8I2>/WL/POHX:K4Y]F56.ND&V)@]^de7D&>.6
BX7OTR3C#d+MPOC#Q)Q?W#=V2\WZJg2/^T2GJ&gHfa[f7Ec?UJ5g3YM;?1aW]B1]
W7d_L1a0A>O&GQ2)Q.F4B;gQ<_QK?>\_-e]OI<,,;;;+SUZ/PGLB^?F[Q>9NcRYH
67[PHMf_Y@[^+#=[T[;6[fVSL+@Y6beW2^1[1-)2&dId/\0CC\=-ZQEF,X@Y0F,7
]@<T>#B;^@-6L2H[@G]ab?0]P:VYK&)ZH.-C_UTG4H:fA1,/65c<:dbIZg]27.?Y
H&[9&?.UL(O04.TE1=FU,bPXcO_Rf8EM:96S_Q/d5af#_g&^5dM)3V_YY(,@@d76
-16+3Z5eK?-=PK6V=27SO,L9+?d=6..:b[fa&2R(7+\?HAA(M6:4Jg)5eI7D]Wfd
&0_G9?<BgGMf#[;D&ceW3OQ<A4[OYY[g[80JNe2cQ5-=S67>SDb(U7KbZ^),cYF5
L6F>fHPQb715=FWPN4.7@T]232^:[-H9ST+-aYR#)S<G>cVS.DOD#6(M8[HQ13/T
X5eVeIfQ5L52-+UcL-4ZP-Q5KT,]DS_&/8?:D=FR^_QP8BNS<9#/<4J#bK-GK^1=
@gO&EBBYV6\)A&KD0&4&]ZXS=GLURWB83R[E;#d0R[LOS3@WEV^ODU=.<P/)WZ15
>B_/>=N.c]FN]SLDO=NgQG4?VfUfQ&<W0C9+V=YYWS[S,Tf4_MCc[7P1M:2gcbAF
-]G.:XeAZF\+6:XX5^B3c]LDd3SH+a7-_<RF7SXRHWCBMB&1;/CE/@D04We08YB2
PaEC^#R4]6R#P<K3&<BYS6,A).7g^9MbafReH]F#XPad7ZS,b[3G\VR;;V8(fIQc
F;U8O2C(QGFJ8Mb1;>(aROQK.0\KKXd0^=cCV&Bg6@53?FV9#+#/;X/-18FNWJdg
D@E_;0UT8W+Y.T+QSCRJ,FSNW,9:eBS\68O9)->^OUDMg,_SS\/,,,dT#Cd@A>.A
>RI^QdMg@Dd<3ITH<^TJZNPC+QXSaX>V35f5./8M1+2fQ1K\dA?N==+9g[L=:U01
HUTH/59,[A^E8HSDd>_GUZT7@:?5XXGYCe<GC^D?H\JeX^O/88+@fQeH^>ZI]44[
>R-=@+^)@6C51F73XUK.bbCX#@U>>g(IGgS^\.?SVf7OS0]^H&,1^:1<_DVHc^#g
@QFLBZf+-@SfLUZ-Y07T-ecY&PRD+823[62S=>A29[EI@aMcAYWC-.CI?ec/f(C?
4SI#XHdd?J=K\:aP<_D([:Se,CS1NSSBN[58<TKF;<f@eJb+1>7\=+O>M_39KaI^
1<X:<Bc(S4PN2SC;1(Z1>CT>5D#\JgRXN7I>e(V9bQ.XU0]d_^4NUgf_P?QcWB_E
+Rg3^+]FPb5eeC#L\3L:MKa.FY9V?6]d>K#8&PP(a\4:[BFe+R^Kf_:2<D.&aLb-
CN,G)PK646FfU?bDa1a@SB:XD]Kdf?IAdCUUXF0[>RA\S_@)G&\G^dYI-L,@OJ,;
TU1X>A5Z(HEg7MFNfa4U2Ue9BaQQNELHM^Va81cM^TNK=?B6Y4QN[8&d^]-<G&7F
M9c8@/B)<)I]7Dg&gSbOK[(KK[cH85N;bY&YI#7ST-]d>B#=TM.L8a/EZGT4OI<6
J6X7>[)BJM:;S3DG^4_^[=d7L+<e/R@9.;7#XX8&VB6.C_:M];/#]UDg@(>#/]bX
7a8@<U68L-L8FEVL>N+O_C]cG]=d(FOR1V4.?TL^c>89U1@9AWNRUD]4[BYPaX(C
b;A^0#91YF9V6JEL8J_IeGVHPC3N&AMLT3-Q=O?Z1;CK;b0TRgWXF<:>]Aaa&J<V
-.?HW8+Z?<CUD#Fc[@O3Z&1WH2B17(]6K2+bDJF9WOLP<DTcZSUD0VPAIWbN^@5N
MUa?..,+Z8MW@41^1@6QYJb<gOE<G5YK001O;c8)0gI/DK8#=Zc#:eE(V.<-LZHG
33@P\P?NWfD.YL-HJ5+>8V5f&\:G&3:3b06Z,R;?4=Te_>c+@@a9;,@6(,=^)F7I
:.WTKMJ:cSMCdA:J]1#1H;;7XA]=@2</cR7.5Lcf(HZbg=Gf#Y=<fM@f<CEfV,W]
\.SJd,MU4[&4b>A7]>1aR.(>M2XDLbZ9N;dP;g6CZCgUC&HFTSK:(dg:g;Ha,V?8
U2>AN28H;S>A;RBNgTb9\LHb@XN0OCOeT;L[7e].RbJYb1#M7_6HFA=28OTAdW[B
CO#eN#?-]Q76A][FF_Y-L94:VSJFW0D>14VW&BUTX.D5HBfC0(D,6aDG2S,8-3f?
SZbN8^E1;WS^[dQfIG[e7fOT8g-GWI5C<gC6egG]2;\X3-TP-S\d]SgL?&(#:>4E
8OU/2gJ.M\RdebC^K(_RR82<_WF7><e#HTF.de@cFC=6c)BaD^_/B5Y>HZ#Y06F&
A(QIF;IA=Ve7?>#E2;9E3a]1bX<F^Ma5CAV_G@S^&1OED+afM7NBP\g<ZBgQ7DC+
?HC,W-^P@XLO5(bRSD-+^4]YSVJ[@3JB[P);F.g,@IEe.K(@21,?=UHS8L(;.eK&
QXD;[&VELZa-X?J;.<TDG(a/:gVIM(T<0&V]c:EOOC^c-@L<,X9ZO,-MLZ)F^YJY
?FD<KC?gOLJXe@<aTW)H3QS))LfIg@8&Sc#@W6:37_H7K,L2-\.VA>aD;M\S:[].
]\Bg,Q]5[c+0IPEWE>)PB_e>^ZU>.S:8g]5Z0B_dFA/J57:W:)AJNfF6.=2R3?Af
_QTJ-JX=7?@3U8VFZXBN(ONdb8R.RN.ST[a_CO^]GB1WIa-EC9QGKVdK7M8\J\0;
C;;aYD<d]Y,)3[WgB=dHF-6I1N\^RLUL-L(#_0R;d[N8KcL?;@J<RVb5SAKH#e?X
J=#G,cWK#Nf,QE;Q976;6aXSf)?N]NP4/A01T2_-KVG0?]JZ.;:N@K33F9GKD5-2
GB<R?[04;MUL2AQ_,5D?^K)J9):c,9APbT8TTBIP>K]A[U==;>:aCEV\HLSfG9B5
#3/.2/;&XL8+U_942D]3,]>B[12@33QL;OLcAT6+Z+\ZOT6\#7?)Re43aY\HD+S9
F)5N<<1[5ARdWdNb<R_Og4(Y.(A[GGXD1ZTZ=)M+d8]QVP;0e03([R>K.7?L92bc
Md+B[;\C=#RQK-9g13F=eb/A/3cAMD<4ZK6VPC)dTV[).1_2[1DR=Zb<MM;V89]C
0,eY-fY5&=Xdf?7PV:/AbRE^X1(;P6]+eTG)XQQ.D^/L-[^<BFHM]?CU>g>-\/Ve
?O,0Ida,QO\\-_c4GG#?>VLZXJX\#6;09-WA-PdI]BG-O_?ID@TUI55\Tdg).We;
])c8_T.dg<g/g+>f4GL3&D95AP[Hd,WG1A\C9V30GY\G>8+[@bCKJQP-]=VHI6GE
b5D#bW]-QWXHIUf#S.N[.QZ+,>PEALIa3<0QeB?LF]B2geP]eb-V0EcZV6O6Z4(7
/[EYUM,A_fHG<CEXafcV5A/=^]>E:3HB-OVbG:.G@7J)<:Y[3Ec5>B_/C4([Z;0Y
_MgV1P&bAD.<W\2Le2a&UV>\#/69&1T_eaVZOXD/P\bW777<P_S))),Y(/>BG5AI
\W_bMdcQ;_,\fT-FKF(JTW1N?fcc(CMP-=/42/:6&N.+JdVJ.41KPCG8JTPIf[0V
b[-SSf0<XC3@c:U-2=Q,(@K>D])4G1QSa@+]Z^Fg0&7L9C(2/;&I?UT;TVJb8g_[
EP4f@K8M[-VYP-#3UP4+]37/AeBe:&)4\S,MC/C2<D.HYTSJ0404Q_;7F,3;LZ1G
)VG(.#C+DEF7\XJ]-c/ZFMN_VaQc]e=NWJfKPQ?2ZN:,>WdFNKV7<VEfM&2FZ4<D
/6R=YF\GS..3WU#Q8@PX9S0]Nc/<Le.f?Z&T494Sf?&=3X>SI,TS><7c9\aIbQD=
#caY)^fcF)Y?01NU4T<W#3<Y,a5NN\X3;5;GRWf)77U4J>YI<2_F.PC95@1[e.d@
;Z>fX[9/Jg=JEPWJ85dWBU7K0QZ-ea2/)26;F4X]QLFQQ67AVb8KF)f&8P?F\@e&
fU43D+gH=US1YJ0Z9E+3@W<;T(f.-A3gRbbK:)H8AT?(R&V7(Q&I6\4OBVAHJ966
7S8J8];4eR2@&9[9J,LHAb7RY?DafG\+@;G3\1C/SZ4[N,#LLbH&4,J(10U[Ob&/
GeE:,32\UZ41F8MaFcL-gY+X7&3;9,ffa/J;EFMDMQWTX(WNZI;dg+PR=+VH.aXD
;(VFFU=./=^(UKJQ9U75ZH3AQEBBFR.H5HP.>E1ZafXET\cM1#P1^^&M<_)JBc9D
Z(Z#G\;3XM/R\H2aZ.G34W+/LZg>8_?b52K+e5.aL?3OFQIHeLE:[Y-U>BWacSA5
0Q<88+@4A2B7g@2N(SHC[ddA7MWYGZ@HTg;:ADD_#NI]47\[_-/H>[/&;5S-?F<>
@@K+#)BY^5V/XT68c0[f1ME::6(HCQH(De7a2/=G)ZU6KB&N.S4E\GC&4T4d?31N
,M7fL8HM500L+9QJO-01^M:)9/L+@58PGBgfCXeT>(WcgV2:DbEXV.Y&+SgC&>f;
=,-:Pb5G<:N[Y6C<Fc>J_YL0(3O&8H[K(EC>_<]=JKb7N,PUIJ0#HQ_-3#_1M@8B
?:PeUBD2;SfJHRY,AW#[2OH(C(eb;3XEAdV_:;(((c[NfBRaEEW<G&Da0ZGg8f[7
9^3.)7Gd&^.DLSf?V4A_PgWIJ[KQVT2QJ_WGGGBg#[T=c98OQ?[eaW-gWa>JFf.&
A&7UfN0HU.P26?VYT4:T\I@4Z@R/&-GfJUIc/+DZE;GPM^4&G73_#J;FO]AR9eIg
32L/NS+J&Kd?_Rb+IM+dL=VX]LeROVgB28F.W-d9-YT3FdX(DK[Ld9Y[e;1H@g.b
A1c5#K/#9DJW5+)ad:_CIL)c^X2MF@a,;)VdC8^@1L\3LFH,>LUH12d9OE&DWQd>
(?B@_QP8?@MPPXaXX,b?HW=;R9I6B?:f);BM7P>W7C&IF4RcHBIC./H?\]\CcKA3
AWB=_7>a4<]dJ7R7)IWG>dS6:_Q,d27,+fC]f)#/d:_9X0DTf1KZ9)#V_;<:WE6B
X]MW66PBW8+2T)gd>],D:J@>+QB^2ISX@C1[DBX\C?>LR?3^:=)7ILFD?T:2?5_>
7S_e1VcaLK>_.MfQG[B)c+WV8ON2\dI^2K.N]3:<QSB[fcfFG/Q658_^L=3@QF]g
XU>-/8@I094+G#G7]MPa6,<E)D1\DT:a\X4J2<aN+A_0gUTV@3-XCTJba8&e<W/W
f-d:K.X=)?&Ge(H@H07aQACb&7?=DU0g[eYA(^RQbDG4f;.K2N3\TL=eVW^e@CK>
LBBP[.S,,P?a29EUX;RcJLH&^bB51I\0S;e<&ZY=;>CgZ+gYSDgWb>TY=&fd<e+4
a,B#]eK_b:R#[V:d7YI):M9224<\UUX/;Kg8?KP7=6c/0GVaaJKF?;1[O]S^_?<G
CR#7E7M)I;d>2M/U>F3)@<^f60QUC6W.00J;3N3O);K&#d<\/f?E2I4&(4>#[b\[
P6c1L@B>b@(C2<X^fH0YN)b&V/@BWT5?e6f]CWXMAaQ:g5GQ#K+A,GRMSHIdM4,I
(<-\.#68N/3;L\QDC-]ZbG@(4c8X?CITF=U6PA9X6bC#-;@9fJ/F#>#V#Bd46^_T
Pf<De\]aEZZOM=;3>[BIXQ=A4.9c845fZE(?K&0.73CGg.E>E/<QG<G8]04,\ad-
)/[/^DFB_BTS)\YI,b#+/Q2&/]IL@N3OY9?^,5:&>W8MVX0XbA^MH^&75eU3U)6O
E7?0Y]eJA=JLMK&Jgg)bTU-@-A@4#PRO:1bQHMJI\CON=)g-L^^cc,B>63]<9V;/
=J?MVV[LK19)C1&HYOf71/[<&H3<FM0&b,^g3\->U@R[g.3VeC1e#K#c@_gWYO4+
&+aH0?UQQP19IbZP9M1K1f@>?3IKA#ILeB&\L=.C_5V?6DM>[dU)7Bd?GEBHE)7/
F)KeX+8HOaSHF[P:C@L/X4<<5M,8e[8\+Z+?P[^Y@UURG#=K)PbEg4^Y)G#-PTJD
W16@N<0>D[)(F-OAbP&LI2A?B=AH-AQ5PB]6+^K>.?c1ee2_S[b(N&+3Q)I.[HAN
/6]6d]85+AQ+_T/44\MMO8LH34HAZ@Pa+FC+GF0@TF=L#7<]=I^B:@EPJMA4RL(/
03b@6ADQCb25#X_F8C#8,+,+de7V)TaKaD=5Lf5\+R@U<;;<2-@[0&F+/P2-/H:7
9b<W]8+T&R,WCURb[gYJ_>BX6:0NXc:^WT0V?=:@M[MQCQ-/aVLa3.K5>NE1GG)S
8B[ZV/,K,)U2=c75?=.+a\A5MO(5ESCc18PMUO/\-Faf0DTZR>LF6;=Z[@M0?^N_
ZXT8_&_;W[3+Nc3ZKW)5+YNWLaC2;;E81fKaNI(A1@-6WUZEU6[g\6X)#KFE2M,]
EO+YfU0#.V,J2PYSaW^._XA?fQ_X29c,8e.P^;XAe;ZfQ7R43LVU;3\W6X1V1;2S
SF9Tdg.U,P#/U[,JZ>E=[LeL_Z4<dKF0(+.QaS(B1MB_+cbbS>UV3[D#^I]E^f/<
5.D170M7JRFIEd>eYa.3[#B4(^J[>?V<6LL0V06I-Z/WR4L#fC&\=T\EJXRIA>/[
WE+B^:4gO[[5WVRCJ>EB)O6=;<d^+8),d.d:/11U=c4.D(+]5Z)A?YBWb&\=Y&T;
_]3U\LC;>\LSU@UgPM.X#<?YCXa7.UBNg4_9)d=PgHNdRI#/)a;a8W305G^-:94R
\fafW(5(RaB;#98I\d1fK=Zb?,_aMZF;?:061HWW(2JV(<9N\<_<?BC>^]@dU=P#
47JBF\HcH09@[(O=H->GNGM];^^;-@eZ-S@O2\8<(H<(017/V8bJ8b<-L>D,b;]>
D+Z2WR-,IA>RFf\K2E6>;_^&Da@AA9.4d,(AgC+/J7@W/@QR2f-#eT4DWR,fcJ+W
T]:4270C<0B[P,KPaV5bFYZ4,IZW[.UL:G[KZN#121;NdU-=Gce_/f6J\/?Wg=>/
PN[Ob3OZH3V;.+]cZIFb?-(<gA5eVf-E5]X-7/3E+5>XL<=7X:K3Z+EJHW,7Ecd)
87/eX\bT5C_TI&>5E>]TUEUY[.]/;[5I]f\O#KLfRI+aN\LW;&2G=4[1Kb4G?WLN
Y_.MG:LLZ/0Yg=QCB[RPRUHGH&gScR(5/3bNEI=_Fa(=-W,c(47NDB]&1RHe+25O
\GbVVGB9V+-IAM^:I.WOcYV:5M64;LcE-+X<BDJg@&daGN_e,5<?>D261d(5g/Kf
]@)RAP/KCQZ)3#,:8ERCM84BR-RD?6S8&I=#:ORAU[^37.A#XQ;g>/1XM_aFfB23
.V=UWICJc((P1V@89WV0YK_;Pd:XDKJb@GDgHFgbED-@HKC_e+abG/bFZET:R\4H
Y=A3e-\B0/LN^LRVRV.f-B^/U05@LMH7(AUU^5JMCITa@2(RUHK.?e9NX9c5^:(+
2c]GQYg]f]3:T\-(X&8Pdd6cJ/C[_:6).bT@PCYQE+9eW)PO,-3=@e,<@S?.ZQWg
M>U1HM&Y&CF.1[c#eXGF51ITTZA#P\]G_BT1FcQb(MaLc[U6G@0WC&4+;fdXcR<6
O]BZ(LVJ(CRHVMFNNaV9/f_B^R/ZY(cfCcKZ]-;VW=G)9/P7_;f[41b?b\g;;.7c
>?=d;Y@<cRP:_3YW.dH)S@9CC\UEBc;F[E==7XWDKf,6X:@(T5f/9=e<9<#G[cR>
Y/]_AEWK;fJg:W[8[IZZGGZ)42_KQCSNS0c0H__WeN9IWeH674X:ZA/a:UAE?\)J
S2ET2HH[4-<&X;f>-d\L6L<JX6\[QcEbG2=?e?[?/cWd9b?DWR[,KIbB8a?+-/^g
QB:g8D_d-^ZTSeW4?YD62;#(Tc?0JgLf=>1L1Z[/\BbC<PZYGQI7X>-THQ)<UNJ.
&X)M;-:8NFb.Y,??#JV24PPW<C]N7AJIOb&>HIFYS]F8<B4ec;;[N-F^&)5ZaFf0
CT/72G6SY)CH3(#LGQgW,D=0IKBK2Yd/BQ;G357/5#eH7P)/#7B-1O2Xd)9,(Q1c
8+S;H&8aDaTDgXAUNHK_E_9+a6N?YF;0GJfaM#XW9P/d,F=G)aXYX=YPRBUL@Z^<
c><-74g,g?C88NR73;f5a#YD\XX[9U9]?U>dD@M3XKTPG)ZFe;;,OI:V?Je+FQb#
5^HX@_RCG_fbW_^BKZ6MF:5W/:g;WG@MA5^<]HT)821[M0QYc?8FM&S5(TPJafG[
d2PDb[f-S=KbfZCJ<KMQ?K5adT-S63248ISD&25Aac6M?b8Qd1bbX,@7&\EJ3CEP
W9&RXU&<D?gMR.\E8][\[O2LH,B?]C#RMd];W_)<6f3K,NI]Y/ZC<gT]a:[1HA;:
@[^DTUUW_[7G_I3XTJg5;W\;;7=Ua#1K38VEg(a<L_C2fT\Ia#=]X.)2[ReWfC<D
>KL-15IG+&#B]S16#>BV,3VY;QMg0V&,)HcC>.Z1g(=--WS&WIbHS25Q5d\\dV>K
gW](4c20[C?QV[JHAUQ,MJCAHO-O5cDBXfc^#\A1JXY.1+S(Q6g/^YOd4P6bYOd=
@Z^3+FBaUY#HgcT77e_55IY[>gBO>ADe>B<UbS1E24XN,]B(NC]gFHS-;e4aWG)O
=IQ\.9DGcM1(>/)H)RNJGG0\;IF=&3Va>e#XgD_;BK-/K-/@/9\aG7g=,YB1f_&7
G&g9dNMJc@LHCT&O1-Z0B@.+&<MDL1X,/LS0HbT@Gb/FQdR_#PPK\#?gX5LJfaW]
;;,/^88V3/45\[Qe\:8e:)LQ43\ZeW7NgAAQ;fQ^2fcIT<@4,B\SaX4NQ=;?[?=[
4Z^9?D/:?^,(GSVX9_QOeX0:+b5(Y2F@+OP=;cE/)9SIT9N[Qf?]FO=/=B41PVI(
[)SZQ?fP.+FDH\N#Y23IF1VKL0I&:,O2Me?X<-6Ea]KKQ.U3IfCV[0/:D70W05:@
0AIYH1)?+SZX)@8EGQRVFM5cH^F),.B0S:J>3Q\RA<K&8W>Z,E(NHI:6,e:)&\2X
1[QQdK0,>4bXOPAC)Ke6=D:6cY+HfEG)U&J76QOHSd#EG3).S4SZ#XKZNV&WCI#&
X)JdGf>d\1[YW,\2O@KbOVc9,GJ.I5-OecAU7L,^1bF-/)XcIe\.]^OVYAaW3U?@
L_1LR5(P7D58SKO+QILX^<ERde:TSP[P-ZOJL28<SQ=U;CLHDAWf9=ECc.Ndf[G-
]Gb:VB-,QD(N8<0458?ROPH7@WHPgb<BQ53.?7.[#ET3W&43B>+04/.2+STI);=F
Sb6<SbY;YQXEf&[efYY;&d-52Hd\,C,(=W:(4B[b.dPSKM8eMQ3^Z^6H^>7dO-H8
]aLYGK:7P7VaW,gDf<O<XPQBE=^f,[0>eeD.&F(-05G<+4bY)cDUZL2;7IPfeQ_N
UW=?2+U=>Q1Ac@M5E14JV@?[1LPJ;5/3WaPXVWX,N9,Z)R]&D1LF5J[P?NCK>>>@
2SY&[D[K_I,A=B8@]e2]/57C]TD5M->eI(d<H\cVeN:CI)8S-eRY;0T^NTIS9YW]
^10I_#:G7NI^Sc4_O->,7/),(@@PJO?\1&e?,-/Sg<IFf@1CHL8QNHI\b56A<K>d
2Y473S7M@5OM5-aI?fQT#:ZV(DFNM>T_3H[28dLcQ9Q@PP_9;54(eEY7.B#5>(C:
8@<gLB2f-_ZdJ5aL^\9fFM,1LWRJX@/H/97@S)?>7G=(5/^#\_0.ef5<VY501fGK
#.ISC0E+-])Z2;Ogcc43M4G+C\A\KZMNOL,B)+Sa2aY6PTDXb#bM<AN(E5:b+V[+
DR24@EE=.G:/3^@c3I9_f3U9?S-fBW@_d@6d_2dHX4:[:Z/@2ZP?L1dfI^M0ag8F
g(.2FY5SQ;RNB>AA_@C>_J:8OYXEa8.:=0#+Q\<KF/\54Zee:LO12CKC:I1BPNdG
&9P4489FZD2\4G^)=8<?O[69d4LXHUH8N:6VN9Q6g_D<a[047V3fJC,79gG91Z(b
HF,XBWJ@MYC._(?:9^/R4R?B&4?.d/3ZZ3TM4P&cf;;WYa2Lg#P?FW2L0QL454@J
ZeICIH>@eQ#EJ2#ANBc9E=T6.K:Md95[G>[?95/CBEL<U4DURc3C6aK)).=J&8=1
]cOceV14,>+\/Rc]Ed,Q0P?&.7B4,ICf0gRU;40=BAW?0:[^-[AI)41.#]&_V1>V
<:H4P)P91^dd2L;7K9FQHEF;K55L]E;=c+eA=^efE1PT-^T0]8.[K45QcUXB[IGN
_TfQ-g:MOLa0G.W[cGC8D&-Pc1Ce?\&,@?69R]dSM)#<;4T?/ZTIJPbS768NO_\P
(ObbHM4cD;\B6BV36ZGbcB,+<eO4R@)X(=6XPS,TJ;[ZF&VFXJ]24-,M3[SF3W@J
Xg6/,D?0=Wa2S9MF/Z9(UO(-CJLRN;NP8V,NE9[eE8J9:76g74P?;C0Y=F<\B(TY
&H,J\H(2cgGCcQKBAHUP3;VD9>^:VIgYQD&B?K+818MFAF\/EZW=#TZUO#/4O-I:
2?>K\??\g<#+_SZbY.M_EJCc3eG[177ZO25Z,7+g7/bVJ#KBV(e9QUV8R&MCJT/0
gR(I,U@&HYZVb.:U)_XY/JANVAN)#9B,<0&)&9F-&DGR&:QO:]@6@)).a-#f_F:g
?dER5RRKK0Qe?S:3?gG-:Ic,gQNA-]Z:/eD17cIS5/.f=9O<GR0C,0JZ1OLJ(d,>
9Fd3::eE>]54(_aOUU1MP]T7O^\TQ,J^)Hc/3.fSB,=Z:9a0G)-c(WLF)1QBQPE?
IEf#BQ6TLI::+X5_8:@V8[?\J8c/7^SI3Z.A-DLaMY46(/=^?V4SMd?[gBZD.@H]
@Zd(FWH0I:)^60CU>>M3e:B\RJ[FBCF)-K7H@F3fGR4#APO[Ogb0B#DPOTfZeWGK
^52-W<Tb3-F@G6)cA4)W&RKeb??:8BbBO?V@c[B1)DFXY:Y0<HcN.=#?g#N8X?LE
FcV3OY:XJZ2E4E:Zf__\;:_(B<<9]&T:ZfbG.G8GdE_b#a)CQGg_BH5I(gGfWd9S
Hg-aOe1XV@f@#7H>d)QQ8/809<dL@]e0LTK9e-C7PD,d6&dAJcN,<?=Q#3QWEEJ)
<KC^gO#2dD&O[IL,12@WBe&e[ECgg\=?7]OF]+c@5T8IUW=-6;+EYZ660Z-\N#QV
IS&cV5XI<\&+UbWYLgNA<D2[aG@DSaL5S&OAZ]#7fe)_7C2F6ORDF&:V-=5I50)e
cNZOWQ5PW\Da9;e[-(N:CL(.40+=MS9L:g]_A91XVD[BX3+(.F]=ZXI&#DAUH4>c
X&FKUS.bXAC]??)Z5@_:9IRS8;<QKVC&7TR6<G-1PE#J&,W5TdW,?E)@aJ\H4MQ5
:1#6B-&@KJJQTc:EIfO[Zc<8->SUbea;8b;f(gT&DW[(V+18Y807(8D\Wef3+D8[
RN?N<61<2XU_YAEAcI)M/ScBPEgY\#TJ(AEH&/OQF;RAU=G7^+39(+GB<gX(UU+f
,Z//GO@W=-STdEH9D1M-[M1T.\fD0.4#g\O7+-=13GgC,\]#+UFYT81<8C,g7VNI
Z-=2gcfE97d@g,Fc+L\-RC)2eHWb5&4#8-72JOG^T-:#fS<M[W@1&7L7I(,A1&.J
1QOZ0A.J#E&d/_-#dWCG/Zg\KNBT,b\ZH[&TXVVM?8)+X(MBH=-a0acf(GEbb]Z]
;]]W)&W)\LfH<G[)RMLa<,/648\3=2B38>^>V:SGCaIcNJQ-?2:Kbe22Z(UPD_;X
?8/DL;BHR/BbYIbg>3KNPYJaa.R?NLD+<QaE2b.0NgdaJ@IaXL>?>fd?_#Q\Q^Z5
DO#M\2>aC@Y,_bd7VV+@LEWL4VHK&?I(g\5OZNQ9LT.bedFVDABEa9[,gZfUL7.Z
>1=U7_;F&(caD&6LI54?QaH8Z<2J6#,\<44]?BX;0;7W882FIQN(d1ADTdNK2--R
7QXecVQ]X]2^C/#75]YQ(V:cEfY=bFO\S(VHFU53T@=?XBAa>YE::[W4CWd99W6M
^dA:#Oa5#)HO\f[,g_LSH-?.BE(e_86PWV?GV,[I>8)>,[gYWPd(UC2#.U2T>+4[
a3)R,-185Q_4b3Q9K#f=]5Pe[3gf/7PQ-EfR5#LG^bXXTYT]cT(eg70gS.Y:d6_I
=fIR6CYROcQ+6Efd<L/NNE\P64SKPC#RQCULFU/B\1&UGKCQB:4^ZGFd<[K:W1Gb
,PLC\Me_0+[=e5T2@fLBCd5Y+&..PPXUEV\==[+C;8Gc(LdXKe?eV_O]G=E&^&S]
9N2bA=[Y[TDb?ZU8gX6&=)VRXEUSQSV=G;C=VW&HX^gIG<4<>P-VXOHE^S^/Q^7+
7e.LBKPcN6a,;08CZcCFRe(L^MAUE0E>-SCK:ZQ2G>,Q1TX&4@9X?eT80N:A),UZ
JV:9d>&G-[,6SgObR\9S;&:Zg.Z[,/LaJW/H22N_Peb?#a5KB-CF>8^X7,F-b;5N
[)d_0-2a5IaO2(SR3-&g6fYIg-GB_a4)79c1.WE/0N=E\I)_.TC5#fOC5QH_AfP6
?)2EfR6VAdU.J(5(g=).6?5>32XdT2W[=LK^NgfefHST0D.4,[M9T-E\Q[TeWZRO
db]\M1S&-gGSa>1(94N=)JL(8.^NMURT&1H,J]1/>[D;H<H2W/7]XO2,V^^;A+;.
JCe3L>[O+(7YVa]Z=b:6T+e=JUc9,P6K75<D60BK5QZ2[U?a_]cK&&/:42=Xa6H7
Lf-HE:(SdW6K)D>=-9+e+?:0&-Q/:UJK95L1\^_QbH(HC3RSg-723e.\c3BNJS_a
V#]H7(9PVD_N&@HJbNYJ9GM/J#Q=?BH#-2RU?H=,OC400&F?UBW9#gS&3>/?@HAA
&+1W?:9)+6]aZ=)GZ>_aQ].7X-VY>72b2STeH0:CaV7@XR26\f5TJ2G5@R5X=[1b
NfO#=T>_N=/R,?X,/O0571LY)V5=)1^\bAbMbDTS;Z27Q4Q4fM[-3UP.P)IWAKBH
L:0eBdZU6-?YZ#VD@H\J_:3H5?J1K6gXKZc7Oe<1X.AVR:YY(S0;X#WId<L_32K=
bMb1Q+OfgES#TW9O,[+Y/LU8Z8E.;VWX&AF\2T7FX@ZC6DgN-J+JT,W8YAGZJ3F5
>bCV;,99U2231#,RRaM>A?[C3AK>PO>GY;S.?ADLH3[5?&HHfYHEg[[GXVZNJ[97
3(#W)X30,c(g(I#H85E1-D+/XJ.e3]b,C-J]]Qd4GM^.3.a\,0G16DUSMLXeC_X/
G@;.Xe#F[)#F2)>AWP3&H<8c3V98AX^fI9UH=WQ^.5^@]a\P]/L&9eQeb2F52L5L
WOY3\SED,6XQ[EbI0-\7Q)[25Xg\#g+e1O9R()BIBI3=F3W9B.;)36UNT/+A?[PE
Ad>A)+5b2OMd(IZ<3<5(bd;N[Qb0-F+Nb#SA)W>DIA.d4/.G+g?^&-0;MO^CGf,Y
&[[BEV66W^MUSW0.81[gQ976@;:MM,T3_,[:8_>O=)-A;_JP+:R29a\LH#AV=aZ1
b2VWEbLU9[N,1D^<,#+_D#?<M<L[I2G<UOX>f_A:[8^3RRb<@9JYGVgI^8E.^,.P
_F]<&gAW872UdR,2_<.I1K.X(R^)bT/?OQWcAKW6eNEZg6YXZF?^7LEQA\C/+f1B
MN;L6)6LEQ.<P/a(UMLe:5D/0=7ACWaL:[2>H&2>[UL,6d6ZST/1Y<<81TXB\NMc
INCg+/aK[[eJTeV+D\bBVcGV\:\Wd52X8_HeZeQ/Kg7g>J6U06b:/7-2+AVJE.(5
A,Y-ZObUDS,JZH;>[_Z/Tf@RWS5+L3db29SU&TN;H+F9VeVSLfR#3YO=FMNg(]IP
0-fDPZ-Sg^JgQEQ,aUH\fb\:)E-P)5_#=Sc=XfY][<&35Gf]9NEDSVFU:bI(_H(^
C99OO/PcHUK/]P4R.RU).=K_EH_@>0S#<[K?F2P?^=a+2KdOCP#M^KaYJ\(8SAV5
/8TD;),dH1O6-:P]]X>(,QS^c:YD<JF_GJ:.b5WLGT^F5K4_\:g0S/cCP/Z=d<.G
R5#8XIPfLLBNgZ)6Ke[E9Qe.3TP0D[U:61<P(X49Wf,C3c=?A4W:+EIUF_VKCM?+
>96(Y),/@=MbR,dW_ROL_9^Lf+8V(/[b3RD0.,0CB(VXVXDfa#2e9Gf&_(7/T9Hd
50d)KV(A+Z#AIO5NeQ,O2+R+JH)V-1YFI[aMO0R[D&//GK\N(F=RbH\WGC+P>@Mf
P8R=dWJVL>SVbV5GLF69gC^S8UfJW3,;]JPM(^FZ]I0#bbX4bRMEJ]R,ZZ:^O^A3
9_O&eaaL&<Y>UgOFUFf.TNS[ASdL\3&\84EeR1@UDGPQ09DcdO]/\fM[:Q#7+cS5
V1_=.4ROIV#K:e^\N2=\#GIOeW>cR\73GE;81N1R8G_#cRT2-=.<.cMEDbR5;9,g
]7,ZfYa<-<-\N^PcM#=J<GU\<\;C^\GbI__TQFbKNa]eSHZ<;=5.Ve-fY(+\,\N?
XGO7]Qd6JU)gg::3_I<ebCCNdBKTa9CT14PK)CLC1JY^S/R1QMaNd,gg63+_5b1g
3g-X=V)fg)=L44JCd-[(B0FS+F(Q\Pca7EI:B=5/KRN(/L;)ZG)081/<YSCX4X8B
6,4:X-gg-558=b0SXfa4I_?-g&4N+D34]8dUR,CO&G0S<UD(D@7HS:]LUfe7FPNG
gEa679V&AK[?1>7_Bbb@>UL9W1F.0;NM/7(DWUQ^]>0IX5[gCd(:S1[>d-=_U6+_
K8DCE=HUA2TeYV>bS;cO5-7N.4[#=OWQ+3Y.SAMb6(EF_S_D#9Cg29e:6f_3>gMA
HXVB)^b5C--F]A(Z.;g,40(&F_518V,W>J5M\L)1SaQ,UIWLS036EPYF+9c;GBb9
Ig]^P]\B6JD=HcO(4dR(JJ.T78CY@U&D2dCgAZE;gdNU@4:PHfbC+ZeOI#J])Ve:
]1L>Ec,5?]D#)eIULJfLGSa0LDg_ePSR5.X.=UIaH;(BfQcVN-36,dI,<6D-0S>F
.L9YcX9/J8)JOcA.8)TW]Ef+:H:L?18,G.?Y&?&:,.1UEL&X02A@&cXdBQ54D>^f
dP&B_J<;\[2H#MPOZc-P^LYg\c@E,FZ;[GP=.5D+=KWN\N3:b5T.FW#P6=#=FfJ.
de6.>X_QI]E@7W1MJ:VgGcdZdQW)5@W1N9C<aaJ.(KcWR.>KD-4D@O@4gTWe+bM@
15U5c=X[7R?#;AH3)18W)6f_OH<dNV.O\5aN5C,SaAX[WON/.Y)4b()G\fSUbXQS
C0F+gFM2K5C.YKN;c2HP[P-bHfLB(/00cd3),I,0?38LeG0QC]QAVB&JbB555\-^
eg4QSB[539P7LbWUFA:EF3R=DfM76dRD;R[cU7@_81LVJ4N/bE]&N69X@0@_X:\3
TV-\OfBV&&:3\^PW=AdfAP/E:6DC.4Sd^&64ODVIH;gg+9U>6_MV2X&bc;Q^VWa7
)BO3BQ\GL9GOO4EHF)Ld:HW21GeZ-3c65ELbBK.BD#0[+8?Aa_+gU&R)/=(J)=R]
.A^bWE22>3Z:4V)0eY]W3fM+0REF<-N-\BXP7K7R,ICWeUNPHe8CV\#?[X4fV?PZ
#H0;WPHO]DSc9+bCG2QFR\U,[U/UADgM3[GFc4=H\O2bU539,I<?K=V)D(-(0A)]
1Z[X/1)X4@P(AaXW\WBQD_Gd6E6P.83U&2W[&)M.1:VL&R8>#JDRYW_9eF0,^Y2,
<=3P32HG.WfBRIF&\)9Re)LZV,fU4A)Jc+NTO^AC;Mc0B4TcYOXM4gU<g=#?8c;D
_PHD6<[Je<]5DQ/^D]Q(I+e4YN#T2dC(RQ\Je-eAF^SJ\^_@VU+T05X_GH?PO/SU
)VUO\gKX^@JIC_gI8>.GO:WO3#C<5(M#.=1<XH]>3?UNZ>[]_SCKb=;c1^BEC4+b
A[dAc#.Q,3Q;_BN,bL_[S?3_OFOW@L)Ge(F,WNY=P@=N6OdP?^<Kc5+,?VdI7<0E
BYPJ5([^_;\bX)Q^-/f1:;GT?:X@4+GETW@dD35?]Q1BfHB9CF>;c_[J4S&X.19\
-Y52dCc,M7AX7c-eS3HZ,R?Q4Y)=NSC.f29Hf3Ud0>ZeU6fJa@IS+U5^B>\/fSaF
TWbFEMA,JgW.fB>fV(^)/8KbXfS2GM>Z&UC0:/Ud5dU9Y;4#RX@AP(JW;6)&g@KC
EVR7TaM2W:5bAF^7VbDPYQ9;_G7S+:@c&Tc)F<:f<&45I&)YLd+OY=Jc@f-/=?eL
73O5?3;BZXNTWfd=_;K8,8?YPP8E^^OIY;,dRCbO_)bePD;_;W>3LKEgOe&<S@P4
T\/c?M3a&7>+OY.Mc,Z&9V36WC_U/59N-PKTa[S\Z],TCcJ:@Ba5:d_S&3P0gZ@#
C;]IdL0)9;NZ^X>BXN0b70YH_fYd.L9Wf<AW@<\,8:[R4;+a:=cB46OgK2>d89b>
;eZb[4QX.]eeB^S[Ed9e(aQB]&5L,O<XP:]g+&M)J-;77PeJ1EO(bE<@)?/^aPQR
3C+f,5)-UPOP\b<EV:L1@S+65QZS>AfVCAG;6]ReZKeF@;RNN#0acb\b95\gLN^]
TLLZ2[UUUUMUI;9<3/a^ce3_858K(C\M,&afFUSK\P\V:S>AfK.)UF]E//1YB9-F
f\\ITNP2@17VML?T6H,_LTD(;U=geR4E?]bH63L[\1?V(,T;VIBI4Z3U<TJUc,#-
^54AC\a,.P1IJ<J,H5->Wf<I(--[NYVE8gK6:Z8X[e0.+LP(JU@RR)dGb=@>A9T0
?=R@E@3OFSMfSC4U4)[ZE?<+.SC3\8K>LGg(#.DB50S;R<T)?7_Wdf]/->XfCe-V
93QO@[4YIa&:RTU?>-F;gREdBSM-J7D45H1fOebLN(1FS80YD>:T--0B-9c=L6^A
^,/./VU_6R71BTS[:S(Pb4QaV5F^PgK71aSSP-#EVNRM66L2PMWM5_H@:5Gc2P?X
e[_)1@Z0G6M4,((2Af41eD1UIS-MfGCUUL6[=GBX3c4gMSOCdYRD757bAMfLQGaP
2+G0KNOFUT-=+:D33Z3HDc_B.M1RVR-H:M_N)<@V/M8FMAUba9XV?^aKeM&](c(7
/\Ff7DH/26?\F@X<cW32JPH.bXXVT3,#\17<^U-cA&YdQ):[HNf(IgL27<4G:Yc=
Z)SR69=Y3ERS0H;>WaTbSM413b+JgH[XbC&FR2_cE(KE+#=4DEC8T85GT3VB:W\9
ONbWCNBGaVKQ()bQR:F)H&=W,H>[O2U7B5,.A]]dZBCQ6af77;W_dF<?U3/b&:0I
c_5Zb#\9AYKOF9ERARG6FTFL,+J]c4>7BB\9R_O1QYe3;5aae4WS\L1ZaR/a0=&7
78&\g8\cVeF\:NdHV)1+Pb:P/=<AN2@,WD6<fFHKI6=ZV+/ON\]()V(F,0X5O^HR
E&9NF^^#=/fZa,RNI;#H1+YK&VV1J=@G@Y1[9aS^-5D)WQQb^b<b_g==@\EC5T(4
D@L5e>?XH)IFD0DHYE<2<]X:eE-<[C=<_KeN7I,^Y3HC2e1RO^7_\?H3VKN\?]73
R)X<]a?T:8e\;:&OG>VT-<S<D[DSV[W-9KN8,Q(\QN&J(W>/UVZc6dCKC:C=5,8Q
O._R=43N^Y54&PIR5TH2GUZT#.>7\A<b2&d)JVeRV3Zg_OLHc<+VY+Y@SbK72gA(
JXcB@U0&bV(gDWaCW\#V6:c5[#^M[4WQ^Nd)DfDR;V:V\GL#MU1FfWH1<&bAED;1
RK#_;HMMM#Jf>&[N,OW-FL0-RbG((fPgNT#;_E&#_J3Rd;YfNFH5EHHS4K3e)8U2
WUd\d3)(BSV)9JQ_RbS;RF0;P_B+Ndg>^RO537EQ@?,<6V]<Bf8,CB#[g+=PB75,
J3X7E)CJ6BU:R^+d1\H(BGGQ=8D:Y?]C56QQP<3X=1f?JN\.,(MDN#?\5-VO9@\-
Y2b=Z)N)&[gXaS;POc[eI/9K9W.QDTF7/YZ4e4aZ+bTFT2+.W@\9aU4M>CG/aV&0
bOC678-S1R6=]ObGZVWde3aP#,SgL]AVb(2gMf,K2/?>@K-=<#6?/bfg3X32VdgC
Z=9C0#E^)V47bQ+V?gB6^&-c+R5N=;ZL9XLCB00UW5PJFY-)\2,Z_059c)68_-1b
;2Jd,OY[QR?O7WSZ7BdA7G4+9X:dH#FgAPgT=1GGI.#88Vdc5J?FUKCT_I8;T5NU
;VC:[E1aSe]2dc@CAbWH)VQ=7fQ8/DN,RJ[0X.N7LA\SA^,-&-4bZJ3DXKT2LX:&
S\AX3.6.E8J.&RBCUVJbNT[BUbJLROTH4c6U0d7_f)()[0bcc<-Sg;BW,5Z5+R>#
K^G+ZJ86?1[[IHKA8]5EHOPYB#JP-ZHVfPW_^:gEF+52^/QUdCHK>RXNK/L.(RP=
U577^E0?7)\-gB(DK6.cd]K5N>b5Q4?-M?9@]<3Xa\e9R7dZRIN&YY,.FKEf;T0d
e>.IB,7W3MA7G:SK^2&Z;a(f,]cEHWL=;M/()UD<[VI3@b[A:@;E3Xe#J/C.d=J1
MU8D+@\YFGFB,]38G389E4cc^RH@,Wd^VAbd>QT7AAeJ:VfPbY:8L:(+cdZHY&4=
#\&W(4T\_,ML;>HTI9P//KNK]][JBPF9<N=>RFdP6aMND^#0A<+4-.[d>COc)b&V
eMgB^X<cFI#fcY8IeF5(H_X_#c0D(aG]02Y;)@AMd(=JQ8f8<=b<&A9c0A=06&g@
?73V(fHY<HTPLW+[17OXYQUWO=05FQN9KdcJa2MA34V2\Tc][Rab^FU2CC:>H9;S
?c+EGV/E1=dKGCgG\T]]W4H7,OOLc639EP4d^WbPg,FcV^C[V;0GDNg6O\^2g:MC
fK@T8X(a+IB+-7)BbfQ2AB742.@\^#XJa6aU[@67:ZgS#(Z)96TbdJ8)M0U9bXQ2
H/WV.?>UZYR5RbK(/04bA?][dd-91Zg]a&>P3/>57[ALK(KfP81[6MSaM[U:.b34
,6\3A7E?IcY_&;,P9NM;eUXT2Qa6bC7[[7N<BV3Q-?V?[CHg.7?[gU<MbO6+8BNG
3J6+\AbGd<X0B,eYX65#PB2X2gFec9Ca0e):MA+5ed&<X.OV:X0gGPM^3T?L>JQD
A8I[)?K(b:KC23+d^9>/<F]>9D2^IP28geb/.d_@<\[/G==F,#)K,]DFWQ=QPdZ\
V#0)/2UaZCc-2:K,QQ_ZcN6S>4+-6+1&2.S=?0U\S<C4)&CQ0S+L7N?#?(S<P_#X
S_eQ9R+0P)_>OJe/Q(-BAf2&5VFbKJW2(JgDW=O/(M,/2Ec5+@MKS9N<S0]3Id.7
C[]?L^.)=5=9>:W#.(@XZ6&CLQTV<)OS:?4:_,.W>8V^AOa0IS1<E#&7Rf?>Q;6J
G8O&ZPNHB:.C037AB[\Y3C^8X@-=Y2=Qc2PbVf7D:XE>L363?/J&2E_BN-CK]Og5
V)DOOT61-Q>8FA9YJE:K6]E??b@Ff=@ZJX>1&(X)FNAg5XD5B8;CE)_:RFfWRJZY
A<=H/4CSM561M]AfU-fIA[AAEeW>7Q?R0JA]((:=HE=aZ896f[d&@[JRgd1-Y_Y7
La\9BT.a+#E<1G5J@DRR5U/dS>&cQ.CU81<I4_.L)72UCNNdO+APS3.F_KP^eZJU
A<DK[-(I=aO^cTUa1#M8_58N/K9;8ed5>;43MfD.+Y2XLfRAC_c(K54WPCE#YT_<
?#1_3,,B[<NQb4R\bKUeN_5.BW(4_W,V8J/LI]H6G41gS4[Me2;YfdfS@53d1/^0
\gGd5D]JJ.Z6f0[5XgQCVVcOI/CVZ?>:c8(5J<S9=QOC<,?L2D)U>47O[ORE=+f1
OA<KICCOa,c1DHJWL/IegL]PPVNcH4F#Q]67SdZL_CF[Aa=C2_-63;Jf0VBO@B0c
:^/McTPWQ17W<\KE-X#ZUHV^e3,S<HU1LNE)>__&H\1:N24a-74#IZ2H4R>\-)XU
QMf5WRIKb1RLN1&GB5MTYHCTW(><JYEHO^PP<.-((&fXZVWL#+B/+a3IE6\^dGfa
8G-ERJOHG&KbR.^5:<;0N+61S9_aIP=D(-;-Tg9\Z:c[83fN6)=XRGL[OC<cTMY^
?::3(R-[O&L6TP#:b80P:=X0+22D+e8@.60bS6UDdLDRNJXV10Ob\?K^c.]d[f+,
^c_8.H;4Z6bXJVIHFCcUbXCW1T:R0>R6ZZaLPU4&X/79[(R<AVDg^W.[0.&fIN5?
2#aJ;bSB4Ng^d-D@W6#DU+[E29^A1d7S#W9aD,,N=_?1;25Ag(c#1E/57,H/5fBL
,fN;=KOQFT.X&JcS/G<O:PM+)c)..^5XBURRXJ_>1]3W/c^3f\)P0<(e(F<DcF_J
=XJfHfK:D.YS;^QU(H_0-)1E7M#4\RHA0,^gTTK-JRTaB@K-=@a5F\@].)N5=_\.
4DO>)+==RN7E<2NS;GeD?)?=N^VKMNB\MdG=a+Y#bY<JLK8(ePNf@c(8Y^)aIODa
fG&J&X;#5_/O4M<^b]fBD.J3f7CgZK+46T--+dUN.g)3..TG?WbEYNf_b;Dg?X__
KR4-UP7c>Y&X(f:6:g1+G+A2FXJd<<(#:GG2AFTN?2+3bH976S8;>9ZLVJdIFX:/
9RNa&3X3,E-daY:D3K&?]@/T49]CI/AYT/?_Vf>6/2KHY_L?F=1/([+>Mf&//]+Q
\,2-@HL?:U22e#[4R/H^Mc?D3c7YZ<?NJad5-AU.256OSH(8BW-/</?A&CbfF?,,
+?:_EWeJ0Yba(dXf##^,02VMTaQ]N/@:f>ea6YJb22DZ/-N-ef7J=;HD]MAK]f(<
)QI(+3K7G4d5]+[D,PU=<_DT9&W4[Q)2+>;5YVH\QUED5.+b?DVNE?-^VfS(+5I]
/H,>,+#.#0K+g&MM[0IAV.bI^?(V7U]a8,IU7EF#KSPBNQSBLQFOZP_4gbd5KWSB
YBNV\F>YgO6WXeKFSaSMT?K6W1Y^)(G(YTW^GHT__(b;/ZA?Y3,bMH92e/G^3ROQ
RCga_(8baBS_?-.W];U:H:=O)LFT(7ZD\8N695SE8XPeH=Y<5eC+7aRWFY,1DL+Y
.@#>M&5cY@=NLP19#Aa8FY@I^.V/Q)ObFN^E/JJ[)@_KfF@X0TAZEO#&J-U47Iea
.N@c,+3JDOeP(Qb_bX7[;f4H]fdbdJOSPG-1B<c<fKa:U]UB6Td]5K^>)^Y?V6>N
/BEM2c(XPIK-O@M_:P_g3^9^GZF5IdO07,<d;g67RF+KF0QHX,A6UDP^DJ2Y/]/4
3P@M]\N1J4=;&;Tc8#eODg-SgfD?Og(C1IDO)JF?9/@<PgfAf-H^Z43a3LE(Dg>I
_JU);4@681+Ze:ZGc;Z-D7&E;1L\QGd+Zg)+O?bAX[g(OcME5Ib&N2D;YgK,9bQ0
a6@4=O434We<5><K4EZ9LFA1\X_QVV9T(6GK1-ELDJ-\@U?;cLKA0LH]3P&[7_:/
O4:4M1g@SI9Oc;:d[eT#faBQKEDJ(]U1;<W=66g44NdH3F3;b@L(,0PNa:cO&[L1
?.C5RIC=1JJKTV9J-AfAA[?YNf+/F@:C[9MDN&HXRccc#[W)ZVd2FQfa>DENHJT?
+<QdT^N@2W\UA4W0S32FB\1S:=0T4+;J3]<dOBO+I?Ue4fAK2=.F>Q\5bOEeV<8^
XQ8I6TD3d-=G+cRRe3@g]_W;P\[>E9=-1-&DR5<O39XZ00VJ]ISP<;K28+?d;g1@
^Kg-)7-1=BZZY@393bG+G_5<&L5+90aQ(NdP9Pd@Y(NC]IKH,fVHQ(SY;M92FDcG
+,(__4A7X-9-8KU\L#KEfT38MH5g(@Y6J([J_UKE-]f/)EDRTD90d01:?CUY:#<L
FEU(QD#;684)PI5GZG_4b(f3gQD/G8)bO78D9#aH0GcaG;YZfO82e<3J+=cX^<N#
YYHH.@)D/fGc[^@WK&#.:ZC]-I_fOa(W/\aGcD8V#J]Y,Z8YGG&0f+<0c6;X;[Gf
7I)/_86a(ZXA8#M-<EA>O,<?VBa=>:cKf.&>R,6fbc?2_QO<8Z)YdP5GR+TH3,3<
\\2?AV5<^)E/Y@\0^J:^@5)Ped/f<V;,+:O98[_0VBE#FQ[TBJFCf#<e90Z^gEV&
YXS23FCJ[L>@0f\=UII7GWcJa<SHa0OAVJ/gbDY=?9_5_/#>9H=LC#>(7D5BZTVJ
fRaHM8>0(_F(CQ5UY><8gGb?2[)aVX[1X[aM&e^J./4\<a.4K1\H1R\/OKABZCW,
f/NF^>96,E@f4f4?ZA>RIX7f;R9XCBR6>(>_fFT;QV,#J(E4K2>+J=G_aQ\>)U:3
f:,7a)764E8[RC2g;.=f22_S1\89M_A6PXW9#/.5?K;K:Qd95W,dGRPEK<>8MJ&6
.=)VeVV:?+[V=N?W/<U>Ye<(.YXBHQA/I(eTJVEAE+O3_&2cg.VP7dJN<V:VPH<M
AY6Cc.68O>,T37SL5Z2\_O11WBa50(E6\#8K(E6V(LTYNUO(3UE=aDX4)gaJMXIW
Q-He,98#DV4L.]L@<UVX6&O2BWd<2NKWD.24>Lg0)C+Y?_A&8EWM@DNNWB(?,COF
@cH:OV,Q2M?5B[S4&]^b735_YNLaGEUeXa2_VM-NC3&ZW[T]=4Yc1J,dF>KJ>U]>
]dT6fPSV1AI,\2/TO+.S98)=N,[WO#G[(RKJ5JK604),G#HeMH13C@F,@+aM+-YM
EUZDS50^Ne8@-D1^K#&)AXa3N5d\<RJ[O5bgT7&.cTa3Oa&I6SXKc3b]^U1\=XM)
BZB;@Gg7eZM]4-IEOOG1c0<dZ4fBS<MPFD\9.cg>/NJ+_XK:QRNED6g8adQD2)OY
29&]#U_]6gA#WbcYUb+Ic)-SPR3;9PIO/9@ZdA^WH7Sc+_(P#1f#@bW\#0A3-.27
G\5JPO?.cMO3E&,P_US8VN-D/[10=dAb.S?8)TO_8NO\,(4f@dG-_A698?Z;G2GO
;@6\F^+^X@Cde)^8T1]2KVOScN<4F:Uc7e\Q4??3d_,GcU\3G3-Ig&Z;+D/UY[@U
&9[:J:FC2)Lc,:NW=aHAS9)+S9BbG=F+:TI,7(+1C_TSUSHf#<@c-SOT882)\FcG
1bB=PGeaDH>f;.a.Q[+])eN@.-0]LEfGQXRQ?<866SPXZcPCT?dN(/)JWE?M5S9)
APYO-4RfQT;3I?RJ;B[c=N_-.R&N_(AcAd/-291aU,C^W\L6cfI/]-5J<PL((^>1
ETdc];D:0B0,f(@HU\B6PU<A.SXAN7\#;bK:7c:g80FDV@<U]YY8H;[^C0eAHQUA
1Z^7b8]046^_KN&A(P._);\?Y@@ULgbdRd9U#5?0W=.AA=g.>NQJ<3HW\PC,42_:
?DWMS^E,=X)G+1A2?G__.=0Ea9LVF-Q1b1FP&Vg@B@AUI@I=,4/J>3:3+GA;#U07
06[e_eV3[1^d@d94#e.[#0=Ab2H>6#NZJda(ELbX1#L_Lg->dC2VFW1@+7K-WYS&
.8-,dVF)0?a_M4cG)E_d\Yb2#-ZCT/T_]8:B]HaIKg48^_f(Zb=+/A+,>P0/@K,]
fO<?X..93#3:_<+5^+dJ59-@=(7Z(H^E\bWPgNeE.4^7-<O<X;.0-5=I0LgIZUGa
^:?Vg3D\WO9f-;_L?e^#3U9Z;BS4KYOTa@<[T\:KNZ8A8HEU?IK.H-]3\2;dc5]U
29H_++OJJ)YC1+9G7]=f@PAd>@+c,28f^B=#)c/9K&-\fcCV9]#bEIN[YV5I_QA+
&JK][ac,JBY_Y:E]L3Q9c>1\Db^W]UB=JUbXN(])+HNUH9&MVe0QVbOEO^B;=;),
2aO\W&F[[#B].aNO.0Y_M0(5CgL):=b9,9CD8:IgHY9,IO<^QeV+c0UA5W:3:(HW
P_@^1VV3<BQd?4/PUUBQ=Z(:b(+Q/>\5W+X35[K.&3)\29.b=]ePYV0EJf?9Z#^d
0M&3LVI&VG,<_PG21TL\SDOWKKCD,H.d//KfeRgJ<J5_+d,NB5dID7c9^_Q@&3cZ
.C9]dWgU8\[,^abIZ,GA0bJa>\9,EFe,RA+CT(-BaK<40X8HI0b-<FcBJQNY#H2T
XOG=Ra@dFO?9)VWC]N[C]-\P5+MHe/LZB7fZ8YMc33O&GVZ\&@1#P(HaMKVQcY=]
b2NU9NLcCfb0(ReEE:1#9d+WO;889UT@HE]5-LVY6CHfPVCTd5LLT#3BRPT@K&\g
&C5d&C^UCEc)4(_=>Xd#BVeU[;X;QZNWMD^f/D14e]:+bd)?D#&7d8Kg:>Va=KH8
9RKB-/NW=^GF+=##Bb;+7Jb;TSI1f:.-K28R7_G<R8JL>G=f,b(2Z8BBVS#]aHfK
dd:1-b@UC&M;[.VA1TYHa)d@(Id0aJUXXFKL_<Z#340\M8C02bQ643C=7I:B6U6)
[P2=YL(P),bWIbN[Ob0,;&a(gIY,J@V&M@3PP)aQFfD>Ia78UQWZ/K_9KB)]d/bT
C?4D4G+1Qf@K[NAW.01d3)>UH+_TK/8fWJ_359G2R.K[3@JCe?_O7?_G,F;O:\33
_]\)8XK:.K^@G<V>::#,V,+87_-?\G1PPg2#DcJT/E5LG5APcS6[5,@IZ?@(MTK0
7O\4K=.LKXJC(3J:XgX=PBEAPPES5[6.4/+5.?406ZRWTG./^_73Za,FB-Q,CZ#Q
7W_:Z,-__f9O7K@aHK=0PX?,?4[Z0dJ/M9\4T)O7Pa71#2H9&HL>\AOG-@IS\^78
89=O5(Ja+\-M)(AA,HFFL:>a)J:CVF[:;HZ4X],)>,#Y;QV5Y[):2:d5Q@_G_/&=
gV7Vb0J=eeN\ZQ4=aE8IBNa.^ON],0@F:<LdD@9Q@>3#eU?(WAUcd[/:(-,?=X5Q
A1@K2F-9d;;>W(((4g+>#4YD_TeYYR6JIQ;N^B0K-?O_I.NFYZI2Y+.Rb)-f_1eR
RK/QJA^HE;?-N9E<@J@VM4OVTBE1WL+/::DdI-B3WKUM6-PCA_B?#K\QF0J5de-e
\ZZ&;FT\F)7M>1BWTbRNNTOQ_1Q-)+3Pa/:1A7@G[[]VZ@UPgE5/DX-Bc&HC2c9,
fJ\EbL@d83,=+V9??8XXe?&bF1KH\bPY3.LR3KW8P[Ib-<;Kg14Q=(&VBO:(^.g-
F)E?OE,>D301.7R4T::&1:5:<-OC7Q-.(Og:WXQ#)9gE)6-H<8CeM+0ELF2<0_Z(
7f;XSN@F/4Cb]D#dTb+Z_gD1]eJ=_OA@Q60+8?&?#b2F2PFbXT2U(L^^K3#U7CA6
G?J6^33g:<Da0_)CRB_&-VQ0E3XMT38cXNgcH53^T5YKBGdKC.L50-0,@45Z\0SG
7_8)X>JNQce;((MEAR9WeQYK+/cHW-/8,a>BT(9398;IV[+,MWY6W/?C/EeBL;(D
\4(U,/d1M/##eRG7S1?Z(V\;QbP5^OD;\)<eV+L8G;^?^B55Tc3P)9@F^e)LX7OG
1Q0C74;1.W#cC<F3_TP5&,G3D)\c=X:f<7[B6d3gX.>+YdUgYaRfgTB:).N)-@Sf
Wff?-PQI@7f,A[fCV_K6<3DEZ.7&M:Qc)G>#W\e^VY^VU>_M=aHg]05I<H+C)T4,
AS_#AP:d]bQ.+4(1^2S=TK+W-AA^bB;4-@Kf]#GE6R_.N-?;_cX]cA^KN&5T=U&X
CBe;/Z6\).(&B,+=GYA<Tgge_?cL&A=2SX5:D\7)MJQc0U]=T0X?.[f,6K3cdVL7
5g+&4YW_NV4=@\RMdRKA&AbRL66,55A0^fd9G\>a]L#O&19(>ZAZO29.12_C/DSa
]RZa0bQ.2WG6H7HcI5a>JbAfSeAfWN5L-(2N725OO(@26J[PHRSWR;YGA-FMgY\S
ZTX9<R<+AU2;/:]FfQTEc?<Mc=IC3L8D+\1@=0RMI+Y7Bb@]_O)R]U399?=AV&GW
B,XY6-#TDJYR.g1_9AD[TRQfFU^^9O/b\\,MUDIB4C3K0]d>N6ZV)8(\DZ+29Cc1
-KOdaA[Ha(C/1>/eCFJg]:R<BJZ-B;UeI5FL_&+Q3LU6Q3KWFa.V;BQP(XT1S)MY
@#6T6LY/LTP74BgNV/fV[2Yaf1Y<:09d,3D+cXcM0HSdB2FHEV<W^U_;ba&[.Q8N
]Q#B?.b9\6)4ZYE)J941g^B&2G\UONcDgZ84Y6g7)ZDa;EccMZe5V9aC:]<E-UYA
-@:0A+]3Y,VbF0^/gP6QWWTGBf71.@N^H.gVM;+gJc.g_/VFWa7/@=(7N]H,bTbE
=b1=O7I2bGcX-=dLHRWLMW;)/3?M@,NFAD@=,I^,GS.QYM;K40@9.<_HAe&5I^1E
,&f[EDFEb_G:T_3OId0IM#5OHEJJaDJJX2=a9U@CHQ]]+^R8#=:F4,8-/_Bd<(/X
fT>K5#DE6-_B?36(O]g?ZVCYDU9PGP40^(@M?>OPR7&#7V.7c:PA6cb6,1Y]12\)
^4HG_CLFC-]L=F,SP4+YUJ?AM0fU;2U4cg/WAaF;Ne<1a5.Y4,(S:VR_SX3J\0ZK
T[MB+<WZg.dQ>Z?>=5AcC]Z1:?bWRYfZUgE@X-c2b+S82cA>D?M@gC;-N);^[#M,
T2<Fdg&H?>6KEJg,9\8[LJK:fVAR+253RK_0W\S7+DZ3CZNC@^ffU5dO6Q(L1)&-
\E<c&/9V9bKC-;M[5=f-=1F^J.>4DDFJ4;a+LLXdK)f]^CNfg9#[K666S,GU@)?G
YA;]#5.Q0ZYbVfRJZ88^5MfH#cW^XE.D6&T72648gP1AdJ#G69e;63WaP3+8ST7.
<Ae3,\O)?_.9N65GY1YdT2;d.N,TMNa;HCO\KZJSOD#,#5NC^+TF_[0L8J\>6X5@
0;.ZU9SLcLC)O/fLQNRHf^V>=+,H4g?UfQXaA5^2(JUeebXfb<_>T2S/.RD#g4+#
>4],3cH2A9P8bHW3)V[U-0f6>NBGTg?V^=,3A@Ff)F<[;e&Ka9J4GP0BJQRTM:ER
6eS1[XW&+<_<4)<;@b)DYJa?RD3+eBBfWY2,^8FXOBCM[Tb9gT[>0#CUYPQ5&Q;4
(3:#_Z3/=#2gI@=BDT3;]GfW[e)-,KP#N00-W1UO1SL\[5RYNN+A6=_fd8^[<D0S
#A[Q_e-&H8=#(;R2]bXLWL<Y2,X8_5:d,754M[<S>]g/D1Ia5O<2Te+E]Of,P>eE
;Gb5XH4@U1P/eI+GIW\ED1>@\:@Y_)[&./Q[+;>=\EdD[\XU8b9_U6P]YMQTWJFd
CUT4YY;4U7JE<@:WDE\]86I9F0+<R#P6_IYgD3)N7^E7:^?ELEHCa?fTNc>YBTg0
gg1H-)ZQULfbKN;CV&@4QWR<0S2&_HG)#a#QZcUG__S=1RFU3N86)U>e8+cQ/#Y7
b\H5\;fC8\CIRg8_c\TK0eYf0Y9W+gDVc7>C@a>O=#X:TX1=N.+@D19MUAgK?/NG
e9XD<B7O&\P#=[0T^O4+IIK>IL+D\>M]F7c^1D:,KWCF]I;42;<21M5LF/ZMeEQ6
>4<f36W,RHYdbcBT>G^8,2-64B24>D#_F+V0dF>EMNe=<1.<MbAd/P0NF)b.Qc>L
@)?e:FX4aWVKC[H@TM-N,X04+@U5E6\L^DMB?Rf>(H39L82)LbE#FF>HHAc7QQ9V
aF48NZ7_^KV==dQ/H;fb87K\WBc\<83)M\8c(V?I[:W@GXc5<)@GORQ:RaV=Y7\6
HOYTceEO;+FDGYY)+:8?fH;LHMV9W?N[#LH2W)E1-@S.M.6070.D&M?3f<R:.eWK
GJ[_+VbOFe:R-YINOeMEQ4a[e:7[EN)+MT:UCPO2dV7(Y>X_SE:D/.e<T&L5\+>,
K#QL7(O_^@.2Q9gd6W=+\0)Zbf>H@\D_9>(#_HBMD@)BCK7/+<bUEU1G3<IaCdgG
FGEIGV<DBUNB3b)aL<J[)RcB;M)S8L,8878X#8f>6O66L83E@FbX&QfW1c;4SCE[
<6,<8Q40I<L3dV@V@DJA0++R[V.##QHLaCT^P;\<baBK<QXG<d7&fRA^0<aRU\G-
LX,\Y6;E?_a71NAd;LcS6?-]7d2P#3G15YK=,@E<GdcgD354I&-T?KNVN<B#LK5F
b+TFR1>]KPeMdH:NdM&_N]:g1<dPg18b&GXTbK].>-;Lb8P1P](&^@:.N,aHX/D;
\429R#c?9:66J/=7<.6PD[964_<F329++JKPcY24-154:=2e,dQWAVa.c7B]52cF
9S+?\+@RW<7PAH?5@[)^c7eHBT669S[/;fI3a_>YDbPfLCM#)M?)N1GdFGecTTa2
b,#]&5Z)A]U=4R0g.IW^Z:8&JS?YX9,UN_U&UD3CP10Ef8+&d5=E1-e;RYLFV>[O
AdY:[N,/.>8&53?590[Ng1/Pg(&dM6aCadcg7MBK?]=V,-W<=W0+<PK(eP^@MKK]
d<bO1</\A>PAe\@;E)bE-C8:OVI^gPM1HE7HG96Y?QS<2YPASGSS5c.YO[U+[.Q0
B(/eQ/@NV-4Hf)GRWH@XTaX0A3(,=W9g<Za0O]BLVY[>)YGLaW_Vc2:g[[d>DcfZ
#[LUTc=UEK1=,b(QGIAcLgZFY]>)=1=d#1LUH/MNO1M;-Y2:f5g&:#NB>Y:+&6M0
[G&WJ@-H26;Q9c\:1C4;VJRbaSLXWJ8&+fa#)1R5GRS+fM<JU^8AO2+)O\L1YE75
[(EENZ(.&I.Z<B.4(@:91aI^WeZOg-B+:8A;e\=2a;7cbAE#IQ(X/BG-W-,3?MC]
C)3@[SI,C)3K1H>4\;a/Z(^db67N[bE=9<2?/XA/N2JFE2<84YCH[@cZ]B2<c67\
X]&eQG@e2>)(5A-RWJ/EBHf>8KUBVZCR+/OW]?CET@/J&DF)&0=eB[H?00@eXY69
:Q=6AMK@GR1]DI,C6L6CBRTP,;EWHVWTD=DgeY;9T18g?Oc\B)&,M?4JK\3KfdY,
FND/]5X(HWF;XZ&=AT,d4dZ+?V^C82V[L>]1\L.\5f?Ee9K6S>0.E)AQP#@Cf3aC
XJ#cS[[#PJNR(29O9AbAN2cT);fVL#OQdLaA#g@fVW_OVZ<XHESR\=d&<K2<K00A
dJaf@EE9?7C]+<1?;&HC^#TbF/)2RAfS7-f19&V4E6-:[]UDbUY]ELXNX,T?HV(W
I.IKE+@-.,=XFeH#b:X=QAdU/(eaG2\A4gP<SZ/P)5ZbSJ+S>d(Zb=&g;GF^EGKB
OH081NHfQ9(_f2F;.fQ0+PJ17]U<-YG2NYJNPF9MKb+A,J6E_0U8^:=a>#b/A?PL
SKF#a/4[I8,B^F&=H&.+U2d?d<E.3;]4gf2]LQMeY>7TDd-\X@0LZR0Z2[H7SDbT
MSD0:IGZ(&;8-fWCQaO&A.?\PQ?W;GR[N6TB4V/+4Z(P1[>-YL+TB(8gDM3TNQXb
J;67AVKMg4/>g;OIW\>g+HL:9N,J\AWE(:#R58CW9:+UH7Sfb7[4P^;e;TD]EOc;
;P=gRP(=<6B303&UU60:/&<(I&LQQ>[6^Z&>P4)#-,45S@77:[C4M:J^AUODDK19
XY3WLIaDA]0HILJE#Gc^OJd6Y+A7B=+_6I\GB^VEC>]U]^;NG5PM<G5:PUI,0K\#
E?;08d_WLfB(c;41Re[(O,bKaB-@,?N?8,8\Zae<P\8^2Sd944Pc@3[_+SaI3O2>
=PTOLBNI]]e)HB0XK9.NL3+(E,3M(S>(_-_FXf2dBILF89=+#J09L;UAPJ:HT0ZJ
F?&49TI:6)6YcG#^fC/YW+SU..V_40eA#W-X].VAI&cdEL3JV@;<)CO+8YD?9g;X
X_4V#7^C]-JV\eaW1287d0IDF@.JSWF0?,-&ESZ-14#gO,7ZFW9(SXU77WEa4g?N
WLT:OXA):3UUL.f8GRbZZ?R[gH.^>N;aD>[AM.AV@7=5)2Q0cP+4=/CYW)4aK7\V
8?d4<XM[NH-\ZcY,=)d#MJ;L6Y7[,=NB73:0I>-d332KA:OYJ^0LUZW[0QffH.[S
]45OP754RC^1:+@N>V.e=SW;-[\AU#HVSW8:P0B#;>[ZUHI]CW2X@]GV)1eeE-72
e97B.P2dBdSSELHf[N)M_2SX\/df+S;I_)Hb#3J6g6JaCA87ZT,T+))Q?Tb?AGLE
^0PDS2N]:@KJ/KdIVEEg;1O0/PJ2WF1XYZf5NQ=^4NE8Kf4g[GYaab_g9AcSE:-c
9)54\JXS6MWT/C8W+\3c;I:JI3eT+&>OB/(fI69B05)S0(M/#cS>46af09\/=Vb+
7[=Q#c8;)7]9ba3d3EcSX,W\O/^QVORXI^]K^)Ae@X&aP\UaE-=d-1I<#/1T&><f
a>E;>?U7E2\D6B;&1FJR-Q?H^6=eXE#TKI+E6W<W<3P/43)Y)4Va&.-S]]aOJ.1Q
2RJX+E8D+ggH9\;^/@1Y<43[.J#2gB_AE;VE,+&8U/dfCRNG?e-De^SbP:9CKQY\
2:b-6Q/f8f29T.:2#+Z4Ua?Nf@WCfVY@?8_CMW:L532/>];cW[=VNPMLZ,KHZ97N
O(#MFM#EJPLQ?9T\^?(?g)>cae(O95@M>NXBPW#)F02W#^G8\SD4_^,+?>a<4DE&
cgZ/UH^\+986P;1[8,M7I2Of))cE+PgMB+^V8f3N1)O75ZYFU^bf4EF_W7O9a/4c
Ygf5Wb0]<9DAR_M=?FMeW\&#FcS;Id+]=(>^>A-;O:g6_A:QT6RUS?7P9+F7=U5]
)Ze=H[5&U(I@:OXW,L#?-eOP;Ea-e#4E;_31/:g7-ce(3JQ\O,YcX.6fK_&:Z-Q\
[+=A;#/4e74bBIQ#LK44d0bQ;I@EWPAILg8JT:]QK1d?\XS>bW7D<LLMH#YU04_5
2\,E)U+1>[DEQ/e<3R9R9]4=S?V)-3=#/CBZ0[1FX,1RaBBYJ)=O3YAGEJ4HOL3?
A;(0,3=fQ1U4BgI&cF0A<7U:7Ld82U?HHTa?KVX@)4Z)dRdU]bVW\U<9d2d(U[N2
\<Y9F-0;/U6GV<4PDIB?YS5+3IYcbV5b5N92-.&.(@<2Ie,R7#XAOJ/RHU_Xe[Z1
C7BL1G:N6S(O3bVFJ^?L?b1O;+^<>=CXc5;<2CW^AaM?5J^_UA679F/]\Z]@AY1b
BZG+-Q?fIgUBCWYfTDf6b)b#]9VbeOGFFJ6X^)e704CcN(H5[A-L5WV_VLa2,6Re
,#1SV#L^I-eT@e2(IY>UV,Sd>e_HEDBEK5f(eOX&fQBLCGHJ+\IGM(_-M5G>?L44
:)@ESR/9/D@<,)1#MY.e[@=a;3ZJB?R2/8\MF-TP7EU&>M89ZS4012J)PPM^DW^_
XQXY&J/:D24=3VP#<NON@THUG[@dXU[I5=g&H[:H#bf751gaNL-P=00?2O/NZKXV
-R\;XI(]1D]HPKQR<UGK-HY=5RI:TLO-K1V1fP6RB\E_X9OALGLg3]L>5>6BdA4g
S@32/^OPILf;Q5bB?MMF0>.M[PG+>FbXc9(e9-@(L)ARfWOJ1U&4Q\G+DP:HD^9e
\f&J&#Z?R&R)f(Z&1F(E:H1H,0K]E[M-7#>]+G=WfGScXa>A]MWQEE5;QAR,9_(d
\H[)B>(M.HNHFEX=]RY/91]AZJ[_>QZ0B];Od(3gM\aP#0VgNE5ZE&,J=?\+I//;
(e\d]L7[L+/A[TacN8255)edNI32A_9;\68(YM@W36K8Bbc^TcXNZ-WVU5#IO;B.
dF5,B]^OMP3EFJK?gH<3;NFHGf5YX/1>.685AYRR8WCH\5bd.5ZdfIU/==)P?;G+
Jc>,WB(&XSE=E+7?B0;O\dV&8)6dE6M;>^7aCGdM<Se.H:&S+0:ccK98T8_Q8XE1
B(P-Y13bfO6/)2bYa?Kf#1b7BXN=eXS#VEUA5]@[TBGeaT8E;DD2Nb7>:JVI&FVB
P:4\dQfIeb8)][74eV_+O@,I6#63/R[eLF2Q7LEFf2V4.)->Z8N:6_/)G&I6/]W-
4M[K?DdJX0)EcUXF5cV4HU/(QdZ>&9B<ZI&EPLC:M;cUR:UfRT29E>+Pb&a^[732
H&GcN=5Sg)R\JVJeG8Ug+a3V2(]KNCVENg=/aPZeFDMB5A[S:Y2&)P3.HOT&V>97
+(259KQ(^Q-G3S(XA[CLOI>WXHV1V[<C5L+0GP#S,/58D3)dV@K0W#@7M&Y9eFM;
3PWD.;JTDR@=ZU3>.cLB,DYb[ANBB_7=7HK.GL?5.;79(<LWBF)cY]AeC5/KZ?9.
7C_@3A]X(c=\\AQcfM;-c.H+JIM[RPd0,@);bdR]3@X<;<UA[(PXd9J[&Z/I;eHT
J0+c.d:X(<^Wf[SLHba[^P3JJZA\ff4f\V<9G(EL9V3E9cb@TX6G.;+a,abdO#NN
;QNAY0T]+(.^)>Y_dNI^Q@cOVK]=6C5[F7,(I>DJ2_>)=K:MGXQ(NSD/2TZde@8I
W+]84TdQP&@FFW.^f.;E[G?<>YSe7&L8<B7^T7bBHW-=-/[:)2^MK&)<3SNXFAa6
0>\b3<E(a/baZ^-6D9;F77f-Z5Uf_cD#FV6TM.H7fYH(dTC69.=CfXgZ&L1SOB8:
(L12)<L<)e=D[aLa1#(@R634ZYg(=g5-N8R(I5<>[6XHQ>DU<F?/OF=@O/.MMC/I
=Y9I##0C0GICECf?,<FC40_JT^9NQ;]G_B>d.dOYV[.g5\cf8-6:@,X=+G=4O<Bf
\eUcPT932\eR<Y>BQR_;cBMNU<?HCCC7<4#J4T4CX(&8c4^SD7e7S/T&+?D8KB5F
5>ZQ7PTWU:LDF/#673D54BY<\AQ8212-0/,+H5S[;@FYWN)WQLV14=.H>:5?0^MS
f)_S[eX;S.9\F<@\?D8P(@W(GPMG[Rc]EY_[&T&;Y6TPH5Tc7b\a]4BM3TD[L@FO
8f<Y2]/D(.U:1=XW/8EYd^VHVFeaZc\,g[@ed)6/=_N6Cb+4R,6]e2><?F6c[?9_
?1Ca5.+/,c94RPHb,&gCbH.+S2/P)5LTT.J-aT(ZMG4GH@QX/bVC7KIG7d1?cR0U
/@R:BZ&)CPJ2geYUT1AFA-CXYaJ]]cY5\EcK@Fg2gfg,]b<X<Xfd+T0U5KH[dN@B
DNPYH([T+\L;Y+O+D.MJ_=NA3Qb/g+:ed6TFgJQNKL:dE80NHa9cJM@^Z\NGP0SA
G&K^BH#[FeW@HDa.XKE8OMdW6>E/]^L.[FB[IH?e+\EVaRMbWfS@a4dN9gc@9BIT
CQdVF/3TRC3,5D&7O72?,4?1FP=.&6PUUf_e<2/;W).E@XV?P<9a@KAKO.)cW[a;
GS<d.bN\f4DY5@_,;/>RMSYT:b?^][Ea\O#TD>R5^M/a(,gg,QB4K6N60W\L?a2&
J\gMZJ<LU?_bM[.FAaU_LRTO:D<X=^2B^QVXY+:aO2d&&fZ<ZAD.M-=TI(U5Y3C+
88\0WY<&(#Sf+RW>aH9B/Kc#/J8L/c1O:)9U_Y;DK<QRdVP_)D/L.def.2O+2@aP
=,bdCMDH_93PJL1gB=TN:Zbb99)S-J87CNOBc938WB4YVMb9060ILD2E@aG.;OD@
I6G;C3>VVC\g>fHU?9<YA^PRDC,0T,cAYC;S8Cg;+)0=Af)]]T92.dfbWcDUI+Y\
?&3+;:6AKLN8JVRPA221??bOZ/YY<+eP?#__2;JB\fIT4f\);1>MJQ8eOWMOd]Ee
2c#5e18:?,XP1?Y/6\((E&J1EXgaTKYM#1GE_A<e61g]Y_8;abB-d0[14S/LK)X2
GEL>E^/T&PgF#&,I;?I7YDB3d4WegU&\JC)N:7D+\>P8cLA=0Y<-N;B>LOQ\][&_
]OY9,5gU=-8f/D/f)X0S^b<SF//G8e_LHI3.M+O1CJ.\63[-Y5S-Yf.\Q:0[0U?[
Zc&KeF#+?F;A=QE4>_5_ZgZ@:g_1[/BE0AH,A6P?QIHZ,]?XXcPe?ZN?[)<CJ>Cg
Q4JIQ@=5OUSTG7V6()=3f@d_E4[b1&ABV^]6)Cd]XPFX95WW7KD]dL/3FJ:b>,5,
&@Gf?YPb0Y5ee267fga>\S@@D3#__e#&EQCe@(=dBbQXKX+a/UH7C9A/J/3(4N;8
,/\UUg(a3J\+SJgc=C;),aIV[#Qd;.^?RF@FSHG:9+V9Z;a5#L7XF(P:/9eE2_8@
ObM;K0\ED/[65_68TW[__QG-DCd>,d5e4THGEgPJ[OD>493-VE)f\3<K-DU6H\(#
\,c/Fa?N4fO&^<3-\PES@EK5\+f?]H)Gb4X>8g3M:XS,7+AK.,QbEe0-9WU;eZY\
&?0GJ;J[./\4>?a&&)XaAd+&KS;Z/fd<M3S@E4;L&6E^5d_#F:,J(BVbfQ8CLEA6
7G0U]Da[@\@Oc8TN8C]7K8@GG1VI3I7b,-GOCX0@:>GKf>]f+4LK@V8P&Q)IH&^\
cVBZSCXgI3G780[\^AU1.a4_^5/<VFF1Pf.6;#eG1Ba7K26(c?+_2G11O=MG52:>
)6L<BC9G&C-:)-62Va5(S.Q,+I:C:#H56]T6@@VJ:_1;D@6d?X_GN2X9SXRV[Td(
CX+:RJ7_O.J2C^RMSc@3?/)W.16XMH,SXa#\YEY:?JRS<DAB#Be5FDW#6CK-_b(X
MW4OOF.:UG<@7K(8P+dA@fEWN6YFcA^C_5_QNMKe-+OcC,8LHe?6CRdY\S8PIV6Y
>eA=(&4^<WMF9A4f4H.#G^Wa^.dSbKGgV[1.SO3F#27-gVGIe&91cG?bXNJ2J_&U
^#1[VUMSDI(@;Ad9HfVX1QOJFHWZ#O4E)a99(ZDTQ(T6/@#IK,1T7g-I#,^/\c+T
[B=NNNVVJQ:^>+Yf3N^7Pd6X0J_fL\POAA^C=7H>,EHd_&;,NMUYFf/+00K5ZWE]
20c(Z-+0S&)/cEbeTVD2N&?8B[4eJF);[-/594cb#>Tg^X8(3RXSU>=/BePL.-&F
DcSCbZPcRJKAW4[1Ja+\Q=DF-D.a2HbdQMU)FG9VYMF[^HgF#1[gJUIC.VDR#WSV
8YCMcBgR1W5,S872O\O(H63N1EM]CCAP1@@>4#eLbSgQPc8LVE6T>J]L\.U-T1=_
._QMc.DOe?c8gTdcgQ^R12Yd/9WYA(^M73<93BcIBJ(/1_+UK)-LLQ&cZ_Gf0fJN
Y,7/4:U9NYLC,@Q1OYQ?([(gYQeW_(+]U+_6aPVe/:/.A<PP=VH>d)O=KF^]GYP(
^&FUSZPH5^Xe.WF\C9<IJ9gSFEdNR2g-SMNAF[[QWUA1S9;4JR:HM;T9E[.BOOCc
ecJ&IWI.US78F5@T^YVBMGRc@I<[?/3b(#d5ffKdNf7L>e9-/#7#;dgXf0G8bcQe
f+.#Y/J^[42PQ&UAb.B5Q\P3D[\II)^471<RD?87K6_2_R4I35AC6&@HLJB&SZ+(
UX&V(+M]M^U)5(\]FF#Nc(U06gT^&XE[CeKXdHJ82bJA:^ULQJa+4g#K1Q)):FX8
;E=PMd?^=@65O3S-IgW7fQJ.L5K20=J)T[Q4ddU5^TG^JJe[B>H<XcaLO^RZ82aO
-1^Pg^a?+\gMV[0aX>_;AeO.SXHP3J&E<_Db2GLWPbFUGPc:D=AWJL/ZWg^-0OK(
^.#__]f?J28CFKDT2N)0OHNFIg6NNeZeG5a2)HAAfKM27@f@PGB5DJebSTeYM<]]
-(\W,2@Q]>(D>3I3#G22P7E6L@[;W(FZC^7C@VfSdd>WI)GMQa.+[+N:fD/#K4#A
\-F9bF20)KB:2GfH/](4<:A3D/9?Da.K6KSE_+^O3@]WC\WVNFV>2PJ0TJ<PT^<#
;?[Z0)T1ZII\=5DR)D=]RFe5>(VY@#NaCK2g-4:/W/6Gd_>80F:XL,eYFK:4TWB?
.9QgZg,,AV78gM?+DB;+NF0-+baK9X@)&&0GUZLC9KadHLA40VDN;cb;6L:AWU,d
W<,OUCG^27-0/D@YM8;XLA7;0EP6NVUS0M):g;B2I_FB9eX3.L=P3QDb?YSN(WG@
MT[MgaR&@10=0&9,1EG6XeNN2SOA6M/=20M>ZC5b=(E&C8d6<e64_QM;O6X7D4=V
DW(A^+2]_<HeI.ZOX^:#aDNP5RZ9Ef?131T4gS.EYK<KN/B3@>aA]ITY\<=Z&R8#
_1LV9Y1f[&B9(LKQ8SSZJ0ZL.F6MJ9USQLe5W>0C0#EUg,A-9#Q3#cH:_0^_<]]-
)7cFMF&ffB_,48YUNPEd1+#de.He3Yg0Y55_-[8_#,6@.QIN)&6cTD1eEBQ6FHb-
Uc@52._K]NDV6L&M+Q(]VB+T@6/1HB\/W3;16Na4I^W]3.8Y77H.,.J\Cg#c@_2e
5TUUG:b7+WgNcbIL##L);Y?\7-YgVZZZQaX=R@Q^,X\U>c14R1,OJ@ASBEL8;,OH
8V8<PCafD[6&gA-R)L\]e&GMaL\gfJY(]N/MD:OPRZ8QATW&de25g;+YVPf/dfa_
b&T;N0Y.@<>-+?@1^=A=N^0@-KPIHNZPS\8D#@:c)#=_0+<<?T+Df=]cLRF&1@R\
AdA5FQ[\775+U;IB970F@A\fXK1aK&;,V>ceMJVJL(SeLF[V33MC-LK:?MD:@Bf5
2,WXD=@c?c#H.NN1^:76;7Y0G_1B7>^(HC6UFU]6XC5J(a+QAM]e39dJ\+=D4:(]
[B@[0LZWAN.,=)DW-b26)(<Y/2aHcF\HJ/6GRB\2=H-dCC-<C2g_.abI6L&;4?1T
\ZY\>bReU-&QLL)8D8^;3^I118=e4=^]EEQ[ZN@]ILE3H\P^c?X),:fE8;\2c=7V
<Pa^Q9JK6_Y3/)E9fdKM9>YV_37H8[gD99A;dVN;[.0Y-AH9+39/.?)Q0KT/T9U_
XdV5WZ6&/EXUA+]L>T[/C_.FFd.2QF=(g.X<2DEAZ]+a?VJdfb<AH6We5.]O]>&E
:Sb[QZFZ(PV&,,ABF3cWRB?)=d&eN#f8F=L?1Kd1?ZNXY0>T5RO0-W9<Ja8[?BfN
d;IL>QK#8#\IXAL7B(CER67]6/Z1X8#d?,EX#eS7/=NfEaSJ-T=-X,Ib-WMSRR@&
F^T;U:2W)f@-+gR@D&gd.E52/]C?510-2(-_:dG5d;(K)VEA;de1S96N0_#@+;bd
XV36S>b&[[fEXf<L2NW\14<7DgIXC]c,QNG5APH/X)7cVL,b+?H30\.KV)6>I=dV
&6G(fF[:Z/H59V<(Q,^BMHZ3fW-H=.7LaI1TE7JL&bZWPVWQ,1O01[/HLY@S.:KI
Q:>Hf@aA4?F20S_1bEO9?NgEUSK;SdVRMOWW)UWF<+4WaF?[>1]bO+07I7>T[ZUC
3&B&?J;Wg_.^[9VS&<-cJQ3e<cI8/0]U2N+6?AD:47caV0b0F?;b)PXRGBE:<TMV
f\gG@?4H]QPgNOVLDfYS\@0X-O6;]^>K>TS8aaf<&J#TW]P7[4f(KX,PM0XUH<0e
DZ7.,d]:?f:NFVg5_N<:BOB?2^TT5\:P0]5R.YN.ZSCJ-fA70cR69C&N,Q=ee9OL
KEM0VS]&8c&E?&U7O\RBbe&#]<fZ]a2V7cQSJUFO^8(3RR1[Yg&8cI8T@]GWF<UW
f1b]b52CEPX)Ve)DVUI0a9Y^a/87U:TFGG@Z)189Ea8a^>WE_3I>6KN_:2&M2/G,
7+Wcf#(HWGR4G30Mb0@^^)4&WG<b,T1&;54L?EXT&.5dP,SUDO)(1[Z>&N]0DTLD
+SbDS-ZJE]&XJX/HG)b<UU1+6RC)&?#F\S^(-dN?Z@#X?AQN>LBB)].,?3=/M6GF
f)\=<:@2JeK)fV.95MM3E3f?&.=FeXJ-I>=D7AMMN=8bK1,05:0L_HV[#,Ma?+32
b-bUHU33JK(HBS+c)NWD=5#R&B^O;<;R?A:cUD,H<C.LL56(_MGGYX]<D8<&R/P^
2GTCA(#IGY0_KBXe0H>&5B0-b/?4]9Ag5EVRAT67AT]GH.U^2fTddGDZ3RN_QC3F
fUN)b?^#^DcYHg,>H3D:XJQ\TA28(B2JVTG5Ge/5&FP<QE>GfOG1\3@4\3Od3\^Y
a[JK(D(_/?L_G\IN>C3@QG)KVOFd^aDCMPP5U+gffGN:)G@</>YWEPB/ggUM>d>)
SK]9C++d@)cdG#51B>,?@VGOF.66I#422GTeL)SQE^:gT=HeJH2&>Y3+gQ>]<;bG
][HePH9N;;(((PA=KWO4GcSTFJa:.TLFQ6eb;/YSCE<#RIH@=WWRMf,c6)T9>)WO
KUB:Tf(N3NL>#HUA+UA=W<3b?;2LBWbNeWDX3?LJ^0fSKE;E<]:IV_\ERG/[I040
Lg7bU;-eT,dZ:A_&)6/<IcVV(g-=RcM^d1eBSJ8W&g9dM4?^fg.4U#]aMc)]AcO;
+Q0PNS31/AIKB55OG<2HeUE2#eW1@PdP-MK_ZX[6eL)Z]>7H#dLIP7Q)5KZGa9=8
/aE@J/45b8&(2Kd+D38d(RY/KD<2@F.5-0?&HCJJXW05A4eRBXJ2+MT&8.(O7,Fc
/be./4/(=HN40VI^79Z1Ha_QaB?eWNAVZR2S#L4OZ@;)[]Ag7QWgFVFJFP0DU,&O
aaSXS]Y0EX5SPbC2@O_+<20A8>>V==52a^+TIB?=2Ra2daIfG9>=,bU&8ES2Y\4M
2RDZ9f7Tf@1UI-(GWH,OgBdgGM@IO:KG<#ZBSB0)N2#WKQBX&7_5R,8b<25;CEC3
0b.H;Vfa;.F\02SV,a[0WQK>T=1L/S<?QU<<O#_<E?;S5H\c@f-A_eVN+&ZO<N2G
ZTF8?3Q;5g2cF5/K(SHR)c:\:#,51HJ?^P8=b+f-HV353SIfXREMY:/01VOeVI9&
I-2VLb_\Ne+Eg@e?bN<R<[2b-ZEPH=eJ6\[RCR&-F4W-KKeAb?f]_\@IeeE1[\V0
>@:HE(F@<+71YM<_>7Jg76ReEdOdL4>(3APTAeW1g#BS:K@C+0_:,?RM618e>QJ8
B:BFC_+1@?cA5NU[+,4N\H)YD9Z<55BA]dcGU+@[SA18/Y7gS)<MDeWQRFLD93ag
A(bNH5.NJ]\H3/VWX;eU5@8DDBN6Oa=[Z3ON5bTTgZgRVHK\0G@3_H3I8aKMU/DB
da.D[P_6;\<R1H8H9M&MOe&6OcR]5Sb)?DPX6gG=aV48ATcZ6YHK&6gDLf9#fFSg
Z/JLJ_CFEK3+SBIV3@F.+O?S_[KD<JKA[[bAY25K@)-@e@T4689G6F(&d25N^BM=
U8gS6LA&BAM#TD[F&>)Lc=9]cWK?;JC]9_gc+\PGRVSE5aLfU><dB6/NXC0dPa,[
+WE[\2fCDRFW_UIC:87->bf.S@CM^P^BIdF58[B\T,#9Y\J@Pf_NTUfZ;OFd,H[(
,11S1]AaE(Z1+;5@TA@(IS8-g8I27gS8_=5,ZR;/_1bRgNYdgVO^4E\B6_-Sb-TT
d+]3SF?5H<_BL8d0TeQB(=ag,K)Uc:AG0M5AE/M#KW^,6<G+N(6#7L9NG0;@SLE@
0-H-H4KH2\&bUfeOJb=+@e<<@VAS7?>ZJR_Z/.GDIP7#DTRYMRF+a&>IAA/L(9fN
[+Tb+U]?@0N1DW;V(5Yd0g2UW5J0X:e#D#]3-DXBcfg:B[\R#XARa(cgF?DL2]OZ
<.AD>RKOXU=R^.^YQ=#HDfWT[c^6[[FX=.U_GT(E\c0b-AGNMHaZS\\dNA5V_1aT
PN#dJ\/RTPd)V8MM/W]_2RZ;.e)90d)Y()\)07K]<DQ1eFFPNFCQSFN0\f5XgR&B
FeB/1AJX/7?VHa3Qg+FZLf0QYPKG-^(W7g9f6RCI;V=M_DM9Pg0BCQI12b:020GD
GSd.U9=^Wc2G7NLCZaWB-f2P>g:H.8OTX:+<MV10E:;^KTO^S:9C9U^XF9O.,3N[
Fe?J92He4D^__7a-,.SOM@7Kgb0cU9141X0@XReeFV5FJc607S&VQ[Q>WFF@\_bD
.;JR8)aZGfI6TM4X)N/L7eGe.21=?JRQA)D^O,G7Y4IYI;cb6GFP+)EU@YL#5UXM
>99(FYQ?e0c=GeG5&\D2\[EfReI#/?)MO(gHSQg:2)O+_2=OHZFOK^&Z.2LK8>H,
M,0gBX^#+)HYOa&P6bH)d\O(SRcZOYTE4K27,T+c[b2Df?/gcOZD[23]gGPM:+MJ
[K,CBG/fP1RfS6-AVQ0QQ)URbEN511>e.[:=+8&eUQMP:2[PP]?]/<<e8DX5YgF7
Z(]-eS+RD8_08Je>^E<Z-;/WL7TN2U7;&@dH_,?]6KG05Y[:3Q1BAF#[2.8SP?BJ
7\eVfP;YS)0O1,gc@(c#=;[O3];+gL5eOIf0[BM>S5Vd(=:Wbd,N1]D_MUG1HeaR
/W7GO0>=IW:.A\IE6.V5UK>7f..fMZXdY>EU@?eO9;LU81<6HX>b=-d4_NJ(fY(D
KU;9(8H_.LcYeb934cULS/5^dC5dG;X=f>YTJXF2FPUL137<II)E,,HbY)JZ8WS?
^7/dQ^-]F7\&S,^Rc&bUGO=@ObS1DNP5HZ?7(IL)OD/dd&f3;FTOS&S\g-0;SVUU
Q>&;8SC:WOR2<g\fdf;bJcVD40?KY6V[P,)78gK_?BbEC\VH8#^08);M6YbbaPO^
e5?W=9G\8I(eFD(KQ8UYRQc8[L9f19A##8W=);d_1FPf:=#.NFI>#NMc7Y\J=3+A
QJMPf8<cdFWS^.:4MWE=&(6I1RD&g^U8eB@+fd=gI2WD-?KT>;gYNd/V0I)^?U4c
)4^IdVf8aYK+//\(TB)_,<e=W3I<UGLg1B6[4KFM;4YOOf5DSN9bb&7#dX6Z)&IW
]:)N#6]f8DO1WKOOb63)2LfbSOKceaN/LG@E_N33(4<:;@E;2>3WO-\S\65^Pa&N
[2gF5=17f4D/WOD3=8e.)DEQ.OB):NN3K[\JZ9DB\eY^9,0()W<)R+9C+)2TF&D@
K3e?L=]EV;YWIVcI6-NUV-OO6L6ecIE6^eZf;/-(URT.TPgJg7MZ]b+QZVL9abF8
f],=L&OM[=/0G]9JSV1[8Gg>P;5]ORG[FScF5JCb37O5>)7b)MX@)cY5ZAL@1?7b
H^;?_(VHJ;E4[H;dQI8X_WJaa-ET8:;TUF8G.Hd>,DG7;9:\7\M<&f-.Bb-TbDK[
L:P-=C0D.+#a>g:L&W87TRPcW0E3f@1F]]aKf^T&L(B74D\Zc>06[HI)6WUHD;W)
UL+]3d&c&BYT^K+HUf]PL1FD-)cHT)X/)H<?<,?EgR3ZK4DZZ]b/F-0WQ3PUX1EN
U25I2UNF.6(G&2W)GP.EV6879A+(2Zd:@ABREGf2PeZV)#^cM)SGXDQ]ZL/0XPN+
17I0Y+,]/(FEe4]TB&07@,>Y=c?Zc,>6_5S.:>D7S84?6I;(^/#ZLJ1ceLe>X>dX
cPK\:PXDNHG]9K&gTT6BS#5Q05e]-?75CWC+YOLH<DL&M[NaTO.R[1->-XbUD60F
F4UcMJ8&f;CKE[&I(=;/4OVP4d,Of1XP6]_DL.,V1N;+,<__Q+7Z=1c?/gBC9Z..
<(-I,H(>X;M+b?dQA=_&TH@P(db^5UD1Ac#BVdZbcB@S__I;g<E3bNO<X&gVN8P[
KN3KN9\3MQf#0AFZ;3(c:+?<RABKD;B\\F#B#\NX3bSR/G[dB]NWU><8_D(KGg_S
B_Q^Le^=EHBQ1H]N@]^Wd86(^c4:6>CcQM30+(^<23Q;3d0?<dD?/>@Z/g#=MQV=
c=]CeUeO>F4Wc94M=?2gcS9DAb9G_Wa(I;,dOS1??/N^SE0^VQ?X6dLDRSf35MIJ
UDX:&aLdA,@#N7\)HQcH-WUHTW1=>:NOD+JC=H><NC2+T)a0P4J;>5PE_X/;/0b<
R/UUb?a=.5b?>f:<Z79B+)a;)c[#PV&&TRJXMa.BXI?@FT6FC.be(N,7Og<,;E3[
WJ3@\+_0b02,.?8WB(5V+_R_>dL6G:(4e?<@VRTgEgCY<c8fP(3g.FHTY5APa=7A
IZ;MMgcLXbR4TJWB@E(9QC,-,d2#M:C>&)?4.5=08F9LJ;&4]KL33(7\GM=g>F)C
TW?_gTS_b76Z/.fX?KIAT,;<1J)]d2+3cO,KHKF7A_&B1^KMgRWeE:_JF/:#cD]_
UYP0<gP,D]aZ?O,Q[UY6\L]&?^K98X\dJ?&@0=3BLV5+XI_BE;_XJ_832/]H?d;@
WG10[Ue2J+Y^YFPcJ2Z)>RM\2</E@>b5BEcGL=W&9ceb+<)(fQ/IeGJ(E.><9e;Q
18H&<V?<=]PI4/D:\g)W_]D2Ma,KZ]WcK@.F=\>;16M8/Uc(N\>EU+&U[9.46/;c
8cFA;2aSE<=Y2<&46DX8eTR4=:HGd1Q5(K018.IX)5b=>TIF]4D:03N7[&;Gd<,C
_)8@T>2E[@B7B^9=BOG1XUSHNb_W_cc7&=V)G#NE4M+X0.\ZecFCQd#aT4]7g(GE
KYK;SA^f[5(^KKIb?aUA+Y8;bKbN:g,\3fJ,D<5JMP#K0^V\_6R0eR0D#K42&=]e
4@a6&:6U^=N\)X2[?V28B0Y1cU?0@N]8<Wc-K@\B6\</E;?2]?(F(fUaS=PaCJ&/
C=N\Z#E?A\XBP(3U=/(BdWH#gR&:[&?V4egJ@T>YE,JI#@HU9CFFXVZcIeK>d?aE
7[IF0UWV28OG##J[3+SQ2-Z4]>?-Y#.KGad,2[K>S&Ed7VFGS&<0_,:?f_J/E(5H
11J.P48C#NA.K^LQ40S>QC\FGVVb[])CM-1CKgf]Q4cD]-N_cCa4f1JaVJ9P>d&b
@RdSK5:OYW@>b<dUGdeED6I8/:FAc5[-/\GP=,:^=T>J9S\P:>cD@IO;0ea<9[46
P/[da0F(/MMB:)b?+fAB.<5Q-:PNJ4E?<(7\a6AQ79_.c\#cBR=ACa2CFD:T\1c#
(c@(3Ge6cZ:B(L#XJbC(NEVf]-8W&Sa2>d>KdD@g>-V,d;WV-:DWdVO_MXUQ=&TS
26b[P,_(7(V[:G)8>E8c;6.CT+T-Q=_N@#[/O&-AVE[:RHC(ZNFgG-UfBeJEZ>/3
U91eH-M73AR1>2c97Ef2=7WX9>,6IVZ/B/=WRRTPG>gJ];BHK#g^+>X7#_G0\;TL
\c&SE[/EX+6d:[Oe7@GTDIfM8bb/2K;U^SUCVc=>GBV;V?0,APR86[BDXU6<#LXJ
S5BJO/C,&9I:Z(8XN\DRW9JL>YD=QDc#FNPaaIS>g^F1>X]@HTKX^eZG?5/5J(Qd
OT[#/Ea5c@8U=J0)\6JP.<b]]\VcE^QGVA;[<H(O^5+dATA&J\COJ=OWfe[D0e^X
D&E1\(88]=T(a2YPcd_Wd6,X4ec_K.E0[NG8C<QEf0BIA^/Z[6=M\FH.4(b?HT&G
V/@?;KJTAQTOYf32CVWKF-SeZcM6I^EdE4dQgafA(7CA&3T?bT(<7,adN5N\a,3H
&43M<1XdN=Y+e\-NYC)]6)T7O-(G)EB.UefG)ZX82D3.eBb/K;=<3=#&\26W@6O1
U:+ZTMdOd5XXL@_KEMS;8Z[9B-7&eA7#bOP[[,NP]3__X7]+4G/WGTO4?5dAWR>D
8ZF\+LbBOIaNE.:GM.V_Q17bS.-).=5eFLF^dE_cd+;Le\7O)KU^35;Y8,9#&b00
B_9@D:?\Eb=?^?0\6N/-KK>@5Q1]e\LOfH36D#JgQ3K:J0e2HZKT=39KX@39^,g-
;>H^Z>DVBf\=.F/TUOgCB-?,=7HRCGFb6OF>IfFPU@3fT@WIMB35:N:^f7SQ)[Eg
CS/=-RL,U<P?7>:55cGA04g[C9HC,7CcUXfe8<[IaO].e?WFOK@TCd_<Lb7KdLFM
<P\AR6SM?-1MX)#:7315&.L<M9/QZPWUaB2PdUTCYS5YKMb.5;1[>,?:A3Q9X0DE
0C&g^LLJ\)TOSC[F?aY^ORcP)bI:/(3F)2Y9Bgb/M-H?[PEW=5-XK3D5eaNgN9a1
S/0\XXEfDJATF8/FL>>\>?a4,6Uf5Q3+=<OR@844Bd#)^-]+V7/>49(EKUQMRA6d
3L=EOF#G>IdU+WYC8EfKZ1:#gZD(B8-5>45VY[Z[J317R:(I?PLJKM]6KUHMZc^F
OZIT5D\dd1g?Y^1P)--<aMUQQA[WY/dcL)]f<^GR=M\@R=/L&/,Y6QC7)UTeRba6
_N:g:5IW5Eg&GJD]IJQIPb_#9T^1HZCIUN-e_ZK(2TVg(ZVGUJ5X>,:.d^WTYO8[
QZUaA?-e>Y:20H;=4P&M@c6d0AMHc.7PWb@P+^3Z1;c1&+R5IBXZ<ec1J+gOcLL(
,bW^EARG<,N:#DI]Ef^Sc-\e/-.[b-+TIbZD-\TI7TbO7\MVd)L#5G]3J#V8[b&b
#AI#ZXVRX/KNNJEFT9I\QYALR07>A#(72#aO=/c3D]&@4,f?^Ad6g2FRNYF;#?OA
c?]Oe])+A.W4?)8QHfQ<a..TIDOEc8f8Q>ZO+@>4;LRYI24B^g(XKIW.dRP?@=[[
W9[g2VGc]W;804W2d^[SDaJ^R,X3YY+JK=6bGF761cNBX)(0/S6cTDJCGJ,463L-
8<H.bF8@0N,0I@>HVEgDN+#.O?aaU4VeCTN&4\#/@Z@CU339MUVL:9)9C\2/T6;a
MUOC@5663Y0X,-e2V[N&U;e]77gWUYVaP:C1ab2eG/A^IVQMK(RQ7H4.^4CE/1)^
L7.P=L7B/aMgR,c6UT-dgaO2bfYbC6HA?dB^c=>NbM,S0]6AO1WbfDWf<ZN;8R:_
\Q?,G,afY@GGIM,&I,.e\U,D61QN()ZbE[;)Z;=9IWA/T-G/28I^EB?]2WJO>B+Z
LX+>G_.,+<GNIeg47DYdORV=Y(;JHa:=3)5JK?BCMM?Q/JP=K,51C)NXLH-a/&g-
(0^JIT[>,YK/(VQAKLZ0/Ef..IIb@#3RA<S5WI_?&);Mb))ffd:CbJ3A6D_FcY2(
dd:#056LDE0HCTQJ\BLH/&BSUOD]>9WXdK.S#4WC=N]/L/-V3IFHKdEUc@82^(]V
e/@JG5H35CY2O.@<]9L)/dAV,N:Ggf,4:KWJ8?\U+V8aVg#\N\=6FK7E8ff/YD[I
X8_a6BC(-dXeULZ-3IR;K&V@TJ?EJeM;cAIYL=-HPMGED_D/<TNB.SOZ3VLRT[Y,
IF[DG_FBDKZZ2eW;1[]bZPL[=SG<OD[LTX=&9e(aTQ=K\\GeK)58cSbgfeB?XN4J
f57a=.YI6_WbJ:bHM,LI0Y/YN<#_)0HM1&YTWJcE>-U;:QNf^5&ELDeTdc@d/GLI
P>0=0YYPJ>>g&L4R>.[OI_d0HgcOS/WMLBU]G6Z+-febc\JaN(,1cX[D5:-=,<YF
V\(cAI-[UJV<eAH,//S5(eRE>)a?.6&3NIF_bcA#2F_fdcc,)QGSY.daZ6L4a3<E
HQZL.MU?Y^Q:-Ue1V2ZT+K-@#[#B5.VH349TF&,_a>Td()XW?)WVf<]Y\QQ^-V=e
2H8;Jg4)3V=-TYfW(Y7CVdYg)X(PYNUHIW50Z&WRf1AAB<KJ,;]ceOXK:Y/0,SNN
L<cQ:>R5Hc]<-R\W2O>3?H@7]D^d+P1__(>?#9O0Y00=/Nc3]J=9KIF3NPG#C<1#
bc3=B+W,@P=)4^dSG128:^aLK;ILc;>aJ/SE]gD6,TUd1_9+:O+ERTM;])Fb#\JU
-)bI8\e2A.O/#)<ad<_FPR.8H((JJ;WP#,T?[=QB]YIBaf&\^XEGS9J;SDIT/Ug5
V[g[I6SQ5;W#f:09[+8>S?a[FU7NeB6BTIXJ4?C&1T<B.7fS:?\W:LC6NbL^JUG]
a:W5>2a0B->;U)88TbXI4:\Qc>7G.96+/D.2ba-C-CBVGYP@@a;++CGgAC8_c77B
=+UgE[C6UA5HL&,<3V?TPS;R8:Lc,\R1fSQ)V#U#<<&.bUgbC=2\^a/PK^[OX1U_
ca]#4BMB,CX4F#\3;FVCPYJW?,WP>0\46+:KG7R7MCd6_IS@A^F2U4>0?;-,N]98
@_?P-2HIQ/]F?-0G[gd01dA#BKaa6-?PP+SZ-#D2aJN&4:#;>H?0cG2:L#(M9d-c
N7(+]]X,KP=XQe8Z>aRL#aV<^?4>).YTW2,K[Bga,05]?eAW8XLBL,&-bO/\^LeR
aN>N@_)=6H>X;P/9?Y->_3K/5.BRH;<K6^[^00J[_FV\+&T<H@G,J=MI>7D-7:<Q
P1(8,g:@AV;BcbL(&7#Z.KFE,(UKf2FU:dACIQe8RX0,WY)g#BU\():,KJ,2-eaO
0<XUMQV;a)EP<eS56[Za&_PZ0-<.DBHHT=(a?AI@M^)]Y@a+W6_RgG7]O@1PI/7d
3/Bd)R2ZM;Zc[<J5<)cM@VAO;M)b71H@:K^^e5\K6?6DC].a@FV304N7(7<U1,9[
<LJ4DH.K.FT219>^A^4cO\(NMb98;<gM^?b3D3WPCaDeOb3;?NB\[>NMRZ6A.Q9c
;V_+a@3R1OJPK>eV9:W4aKIJ]g1G-H9P+DHZOEC<I\\W5#/TYEf]0HT?D@24..b#
]c,K#7<UQ5>NN/=7>XCJe?EY:c-b]&II#M]Gg:<J]?FY8AD/?+NDQ;aEYL;TY\]\
N=2W(^b38X+8>(\87#GJWYQ9=Y@geEJ4J#bXYM\<I&DcgY#/TQ8ADYO:)HS^Y\<.
F-L#9;#<22\O3AIR,/cVGUcDe7(<+U73b<XQb2gXS;E1YL1UJbLTE^7>;VMf@J:J
+UF@N;=[:?O>GV7AL9N62]f?P]Y@d,?D1GX-\N6?LK@1YE6[IIRNf?MUFc\b:JaT
0^c6TQa>eNTgQd@cI?e+[Sa-==d=L;DP]CR7J;_(=9M)2R9>/RTVeTV:dT)Z-#_4
\P:S7/JG--]@,4W^=gKZJ#?[)FVbB5EQ1L@:1,-8(5.8Lee0BI.<N1cZV;,4#\8@
?BYF/N7fY(#?95T.Jg0-IMb@5b(-E:+[bF\(.78NaT>-MINQCO-G8(f>T81acf=B
<[Y.ce/XOM9OX\KK&\<8^YF_Z3]X=P70#.BeEOQ-K58Qa2bbW^9a5M5#-bIA7PgX
=]aB^-OXRKg=[gC?J/?(GG,gfU]VX@;6FDN\.g7b+[b8,&F,:-0<G;4LT^GZI@#,
M[?\7J)b?AC_\/e,P1>dNPB(@LSRK#3QRO(d33I<#<F^GMKUGfXXL<DCYO1e,/\X
0<G<326[D-8Q,)NcOXIIFFX:b9&VKeW)61(2\+GTIZE1P24RPb\J9_FYN3C&eAJ+
;#^e=A?=0JME:CEF-&>&X_BdUN#BC1NS3P[MU/F8B-VZKQeKF<,/S>g[67NCP7?B
3E)987^Z^a9;HK,?b\ZUagGYC95=56-8IbYOFMJ-3^c)@.8\1_E.7MR2F1N>_I(J
3,6>eZdWP1.?b?AZ7#V0\)_0HD)A53K:)[&PDC,-b^H,C=]a+:_5><BK6FFOQLE#
+Ve3&@cXJ3X).geP^Ta1)@J^8MGMG0GX+S;+DZYJfSdU1eGO8:S8H>8,R:RLa&_F
a.BB-6RS3YFMLYV\(EdQ9P\PU2IC\8^H7FUY6\#HCNM7<.M+44a5_M[7MQIX@KgN
T_egDAWG_H.L+)N0><F+3S@R&#HM@O[+)EF2,WRSV[f9AQ(,Af94):O4)-SZgODC
?cK7S8Z:dDa1H@V6OT)3#^/]<g\9c_MM9>dX]QKGI/;A^4C[5Jf7(_7PPGJeS8K?
92K+bHdaTXc_)S[?+R),LH>>DP&>JPWeEB]5_9K#^ER8GVgE,>_&g:A.BFCP,^5-
8a0DM&F<eWE3Q>aZJ^cYS45T<@NYN^c[K->R2TV_cVJ[_YD]gZ-R2^0@F,=[fBG.
@S;&SNE^NZcI.3Td0NEE;fYLc)?8d:@5&3J8MTS1c2LMN_78Vf4)<e)DTQg^Z9_&
c^E=Q/1=-K>IcJ[+H.c=AFg0HRI8.RIL0@9].IQ->c/:HB9.S(HVL3d^cPISG?:a
g8+4/<?-94RD?/ISS^B:U2<]bC_V1f:3Pf5S:Dda((23]Q:5?]0XL4K7ZE[WgOUN
5T>N-]G1gB?;)CdZ)gd^B76OGe<IJg8+)8C7@0fA/W^7Z/KXQIWZ)PPaXLN>f1KY
/IVG,Y(C256H2-_1XY>=e?Sd0^,X@?XKRga(WSJBCd5=UVV;DF.S)J<A,a(gZ2YE
;6&J;?\Y:.Pd/W0OQG(M<9[U-O#a2C46cX1ZK)^f4+Y3SZgd#JG_.8Q<B^B6Q3+T
NZQ2>[4N_7=40_#\>CEcf=_gc4[eHgZ[QU4(T==OgF9LU28/3KV)MD[0EAP66]/M
TZ]XF64LE/G?a#7BVQV\_A7P64D1,BdaEQB&A]eWCW9]7/aK&I[7,O&M]1I?b<?Q
\H:_=(A(+(J2#)OLf)^R;)^6L8a1HGg@A9IFF^@g,:0fY;YdB<-&\8<<eg<g_@K<
.I[3eDe_@BLS^@5E3OLK&=_^29<LAI9\SX3ODQdb&dNU9ag.2&C6./cc,NAP+Za<
RYSNB<]D071L=(R#.<.6-0#b9)cFD^#IZ.dOY;8G(A.aB=V,/,R&=<O.3D+BH9Nf
#;?PMLVZ2NXWAPQIVbWfFAJOCCXO1c&b5.,/0a?R\A_&bRT:9\#>C+W:K1176)b<
+_;(e1VdVG<J99Fb4>K.LHUQCG[UfOHXT]@<-a;X/Mf,ZE>0/0?;Kd#7XRFP70gS
-LVO&7<I:D=4SPBKg,@0J4-8ZPQb&HR/CWI[,_^I:[KD5ea]95);/PIcbT=Ae?+=
\TbR/D^M,(T9:8:a&MC+C8,96DYZbLD??L60N7KT#=AC,4a5df)2ZgM)f6WO@J\7
NR.#L^Y0MUP/68f(^5T8QW?bC30G_N[a_A/V:]_<N8a(G9AU5#EZdRaaG0[fYaNW
f^ZeCSZWb-8?F0?A&fPS=_gPFf2,aeH5ef0&[LL08FUJNDF5^?(U#.RMa0,BOSf?
RCA_J)IKa4::KGd>c>K5??c4J&O[YTR#HPCUD1U4Y<:_VL]b;fY^OEgTU^e_OY]T
_M&T3=#K,49REY&A.He[]BHL>6c]OKZ=6TW[#SW)0MI>=#H?9f^f;eTA.07b1=][
e3\X\?459G2KYX7.cWKMZZ.ZE7Cf8?19)Je_+T/[dC#0-OC>_H<fXVX?X.=LRY,W
g,R)Mfa?4_(]?<a05ZaA;1KSJ=>FYF;Za2QA0I_Pb2b[UM2?6bYd;D_JSS>8_\1<
df_<]O?0TJQN(a<DTFDB3ULdD?BT,O\YP7Fa;Y][>O99&H_RUaBK8I#:((#1V23a
H:e>>1GY^6K^>fI)#fdFB;5VdR9[.UPP7G(T3(DIJ7>O43;XM^2]VU/S[8:,?N8c
WW)0NS:NC+FJSd/NR3.]0>:3CEW>_+M^6>ALBddJb9WYe=RLD]2HZKO9<.+._V>Y
8Z;KR3c_>@P\eM/-[PSH&S?:>QN3bB]>fT2[Ia))B-63>P1J5H=#B\5=Oc+BX=b-
L6fg@+g&A?<Q&T6GEC8c2Q/T&(Y[ga.Q3P\[](S1Q(22M_<6^,XQ,A&^/A0/9=g1
P;DD+?1_LJO[H63PY9:FcVJ(@aI^Zb8:f+eHC^RWAF,\?X,;Y&&,^S8J;[e2U1\4
2RZ.9;(>^RTZF+5W68QOPgcIBcVLM12=4\0Sf9;,H6)gUA(Z__U+X]gA-2,VHg>Y
9fSbA+2C;cdaS2^8L9&b1A^fdMeS;)-9gA=M,F/^(K?ZQPU<;MB/71SLe-g[VN4C
eIL:]=V-[cP<NG7O)W5:PQXf-?HXYRA)KK2)YZT\ZY(VK.8.-B&15^@;]2D[DA7-
<.Y84I]#&=9EJe.6C[egf364TSQ3H/9BIRB/#6#dYL_9CC40-^U:7)5B6U71-569
[c?:LI:)Cf-WQfDB-fK>;6Je6Of#FJJ(bW_:f:&KD5#Z0.3V^-2;faWX^)_d.906
([Ld#JgPOa\=a5_=S1#aMJ2U.G&WLVVg52b4OA_=:-]F\;R+,\e@U2bgZ>I(7#4>
29Mbf42=ND@bV3/]T48:@MJgb93d.7JOA3a(e/F?[.R2dL&6d);WQ[dP43T/[g.G
.[eE^CH/+-7D,C<.;HK7D45D+X\/D:DDJG&<4JLKR4(QJU+.(G:ZafL=>I>>PQR(
X2Og?[E92]Q([9g+_EBf&CHVV50cI7A.Qd)5CS,A.TKU/&SI]Z2GC0-34)?4<9JN
)P4D/Q4Mb[U^T=<beZ<\5He2#ONFMAN.6@,N5I,9O6/-8@J8NWQT04271_(Ogc;c
LES7aJQWQKFe#95>BDU8VFIS)./4QC>9>UHGILN2IZ@(N4Af@<c]1BdJ_gS7NR[2
+7ZVG05K2WH,P:I^05=T.TF(]3[W7S4A=eAOE&2[:&S:_W_GOUV:U;,).bc8#R:b
3,LLES?Q[Y6<VCY3[c&>>4E_?XL9\@K)H\Xa>;eR=f<R+_)Ig[TFAR#0H>Qe@(1_
2ETL+>QE#1IRB>(_b27GX?b^ga7<D8/aG]D#>?Va7RF9R2bDXP+-e-Ie[ZTD9[=F
C1=?YL?\M/@N(DbA(]XdaJ0EQC)6IW@T.G)(#^0Ec2_fd0Y7Hb\::,\H+Y^2LC+9
XWe@GU5^QLF&YbKY0Kg@?JF+B5O8??K+O:#]1WE]eQQ[e4R\=7=(@OfHUNeD-?JV
[=7IR7.,/g_4N2-U>bfU#-^/KD,#ACW]3;ea1?=T4aB=MI73>56bNV6/^DHb[J7B
K3I-8aB?6;.6DZ;Zc9V]-a4@=B>c@WeNYO:+Wc0G>IBc+VS095O8R@a;LbUS>EP\
U)JVD@.580:.3=[U(:>8)C@J)E&6.6B;eaK_/?TO/J0=_^/b&=FE<L-B9BC.:W:#
<,H#&+>VPY?E^H.#?cc#J3,C0U.^[f=PRfUNO1[K+R/RYU)4gc2YbGC5[+@SQ9Mb
9\(SR\gM32F-4BAC<6#-C3R7f?,W#4-c<]9BFd(bI?9F,S13Uf.#3X&EMSJ:0A@M
MIZ]LFW6RX8X1\Z5>O?DVEA0.UP5:J09[,<G00JA(579S7[.0OR687JaE^3V(FDN
=2\S/8XgY&@:OZL]]PUBZ<5/8T?66^B).[NafQP,LS&ZSW@B6=+.BB_WfC/=)3Wc
609W)[A9(>faPU@RRQ<LVWD^XNX/E<J>\UB&ED1TI94BbC>.Y\.,g@dQ=>SOEa1T
.,K4e2XA9ePJ@&Z8^[J^L9>]1@+O/VC5_084:W\:/1SGa6QMa)LPRVG9>bY3>_eU
Q6eXA9LIbC:?_85@]FWI5V2?IZ)ETP2U.90#O&TU.eJVR,@FD?Q5N-G:T[)Q6dKM
a=-,FSdVaUCeb?MV]8[OdVaed&2F082+996HZ.gH097Z\2ZH#7T4_YT-3\)U-S1Q
HFY_Q-.48>^8V[+I4FGQ+7EBS_eLcRb[VVa3AR[N7QZI.-2WJ8:\D,M05ED_Ve]O
QD08A:46)N9>CbTb83X4P:>ga/F(9MZ_g4/(=XH)/g/8-eU+--3-+eIb7T6P=>;^
PK[EHJH[PfRHE-:+W8>U:DK7<ONe9Ta93.C.9;?-<d,5#L9&eMO0&e7N)S5\gI:J
8FZS7dTdaC#V:(e_aQG6HC=([=V.Ob4L=)<)^EM<&g.WcU7B@#gLcD:9HaV^L)eg
1PV##aS89VU.XZbg5YNaS[(f9I9R8IK7a;T3_\Bb^,R-dC_W6M/\0F5H7SED(Q>8
L]7&2U9@V@dS^;]ITbM7C0Ka3SPV01)UC[K+8MSEZ>;=D6&XC#e]PA>L7Y<EFEa5
c?P[I\&/U&3I):&(92a#g==P\X/@QX827#G\c7KE,IBRD]b&;JH12bT:F4F#=+Gf
6X@<:2HDIaaZFI9<G3VGa3T>PF+0<R]YJQA;d;_97IP;]^NISRJIIWVW;Tg\>9EI
PRg:dK\b_6Y@]KdULXT?(B\Y>BEbLL1A@G7ce7B#KH.@T/MY7H8)LG@WM@3HQdHP
K.ODD/KVPWP.Y3UAWKVf3<-?@5f[&TE#HJ+7WcZ(9_]Z&OQ@8D6:.2APRSEIDZZ4
6-H-2ON-9J-^UTAQRW&#+I3.>NXHN-0f\RHGW@Fd+O#RSHV3BMa]7U55#.X-1bFJ
JGB0[TP#bT3\YfQPIE>7DbSJWS:&bMM[9Hc5H;V6DRE5e4SA<\1U6BL4Og:1aOI;
.RFc1J@PL?_#,[WD3adBgR#VN78a^,e:Q&J;LBZ]65JB>g)ODTSE(cE)cK1I\C8/
W1a2Y8_bgN4^O+7G60Q\:5ZNYB9ZJ#9JKYEO6V3a0]a1KcRF_@L/1\KN-7XZARcS
+EgI>P<#+7?WTWZ0_ZZOM(^fPbE>S4_3c@7NQ>g3YNfc_@Ga><BY@E-8VF=<X3NJ
=1J,Y-D+0S:+McF-W=IC1XBa[=X)XVHW/0(;3a[CRQ&e\ABd5DD<CdS>Y<Q>U,:A
[&-dFbOUDP5L/Y:T6:G\bDeH;V1L6c=UNbeWYB5a#+^EE+I^Z:&#HN9I3(HI\C<D
BGgf44#0_TSZN4QGg>\9N5M\EZA6_b=c+9HbYLdJ(FQ@ITMBX^EHREdU=NEL(-Wb
g2BfgJ(++ZHZE?L?dHH&X;K(A\-+7I2_fT#N137H,]OD81T.M2@-2+N@-.037\IO
6^VL\C5?&^+6QE,e.N&&)La]LHA5gIM+=RD][fdgRX@6423R4L/E<F,(=8^13Z,7
9dCCWM=U.3;]MGWf(+I58FE8[2&4VP2K6J>;Q0ZFM#T;5?GO)R<006,UIg&fDKR3
V1F+(BEN,52PYXeO\+KA&^e\0HXbbXM]0-Laa-5_ULYU]8TL.MN##eM6HS#0-1Nf
dDXbF@AKHSJCB+AH[-AFWd-^a<+TT=HQ0BQJW8N<QAW#&dW++VD4:77JWV<C):U^
2;)V.[BYPK/U:d+/O>.KH;?8DQT\^Z^V3?f>gbebcgRNGc/f0Og87#X&-YN4LD=3
?,3AI4aaSSCWcX[,eB@ZT8)E=_R@1]g<W>=fMg):ge:F7_GfQ,WW:67UZ\&;&:9(
M75&<b(=7M\99IY3]7d4JXbQCa&Ob5a-,&KgVBEX2g0Y:6BfR3Y/:0[?T&D6PI)E
)?@,WJ@\5>3dH;2T+_3<ETV(O:S?fffG;cFO-7M2;dGQ_YZe82A>#0-D;bIHf:FL
6Pee-J_4XD6gDK><bUHa+<KG8L[[?O\IQ.ZWES-cZ.-TJIC0.+N(7WIYHL[),a9d
QZ5EK(/7@g\9bJeD5ZINYg?X86/60@A)Q#66faA<fJ=\P..gZ:fbY?Q#7I[P9A8A
B2NM00beJ/-T\VUCPORaJ^dAa9[M[RI9(fa>I@Y@UUR?Z6O2TB]Z:;c_CeBQSJJX
3CR=PA)b_R44[_:_^^KYeeaVDANF09=1e_0dd&#O7R71#T)I\\,V=I#HT>>eF)H+
):]@&)@GD^8C1=K@;:61K(^I9OfL+;;ZBR3T=Q=<50Z90BX]LEa(1@[^FJJ@@^\_
E^MCJ^=:;b.HIN\QB[Bd,P67M3Ff)UQf/2d5eSU^fDT/\Le30.GAG@eJH&^>&QLQ
KGTc?d73,K3<>;/(SH&<_;0W@+/K3JM4DA[(AGVd>SU-6_T8Y@,WWWIdN/bAFFGC
,>VFB0#KGB(_0YR@HYUgI/#KSFXac>VILJ]L?(c^KIcM=daC0A;:H<L,--UF-YN=
^XLdGUEW#K7VZ4;d#^PE?G.M01TTDf,)>=@8BTfdF73>V^L:a\0RHQA7X^X\];#I
(7[c(91/=<F;SE1GH[-)U6EF>RYKPDcK&6^M<=OgeKC&B6b(dFD=:-3TbMa4;=C,
JK&c;+H,FQ3d^[_CF?.M7L0MLCe,SU<aJM#@)(I_?(fV<Z:_.8)a0#@<d<6#87>L
eONe4);(<FM2+BX;?#RfJ6BZ)U^]5_0fJ)+KeC(cEF07ZQ(HXV+PVT3CSJ+Q4&_Q
=/XZ:8-Gg<(gO8IM3?LJ)<VH1[KC&T>;00R@?I9,?/egSGWbLO\Q.)P4cdFODfd9
:WOg@]>e(=^L\)QULffB?2QZf0HC?YaN)(S[&\T)ENEF4Dc@#3.)U;Bf5C?#@NLQ
A5)^?+ZD)e@-MdIg5E=e1(^H4cHA8S_6,\8]0I?-d.L-Sg_c@MBH:N&T5<G/.N[^
Y-.7:DQ^8I_NTHdIC3OcKGT/=5K0DAXeJ;O<<7PB4d:9.R6F.OC@W)>@>8#8NA=Y
aYQ:HQ.ES)_EKH+M_R]cYCO_NO<EQ,X^(/AB0&IT:3>_<a08T[IAP?f^E^W#/QP:
YTM>W;-RLG=]W&MI#F(W,5.&6+HVJCP^a^&/MMbYGU6#QIP@7E0USFE;16-E\+/=
272YNR2<58YZ<-X=6&4S4W4ZgQHVH(:)dBT3;c9MEK\W@+UC(X_fEXfVeNAb2dR&
;N>UIO47O_UYbLe(Z^VB:\;d-@e_TT#][TO9C0PH^FaX-+H1;B5^(>QO27LTB/7>
O@RAGA#f[R#GYb2ZLDQJ/>VD^XH4<HMEF3Z(2\gN8ePa1]NeVLUY=H4QfLVM7]M7
S+GQK]eN5CO^>Sd)X6J^ORQ9bf/@>\_QLK8]EQM#fL>AbfTL,=b(/LR\/Tc(2ZCf
JfU,&Ae(#^GOOE,8@1^cW:>KeWC,YT0T-/9P[6V?N5A=[WY=2IFFA.2aP9\^^Nf:
P4V]&]<R6_]+TOa+_26U==7#0E]3AgQFE+??bXdLYBDA.I_dO??M)eJe.6TN<XXS
eW)US&3V-BM#31(41XC(WcU#P_eeT;fMN+>L48F1IDCVIG]VWaa91(SRSIQM=J7B
^XC<9RD8_TRD]3M;/+22H4GS>XWIJZK8gS;cQ89+)e=5=N1?HX4cL8a?SK@7&/OR
F7OH[R?,ZEcMY41<HLH[Bf(FTB<DRa^U@IAEVKC;BL+6^@E:2=XLS;BZV;DcWeTX
ddT\Oa59NP#1S6;e6e=E]Xac,OJBd#&0U/-/bX0N1Ba..849&#g/fZKeGV@)]g\9
F3O,T^28Vf^Ief7]?>]d+)dcSe>F:D7G3aT>/H+Od:@^)fE[8A-Ce1Z-.7L;9U(B
5g7S_HUWUGKZDB4;[GZ8ET,d@=SYX\]5-F0PbL@(ZP,A8N-gWWJ79dO8eEVbTC_g
5^R@AAH?KN(TBCIN[-N;Ab.cC9C>YcdD;\b[UG>9YZEfc()K^?U@>]2;PW@.#09[
TJGg_7-ZO@[T0fW;gNHUd9-I;<8L)2\ET4,H^2&30J-CJ72f\AYDc2S6KZ4HBRfI
)1FLU[UKY>;B&:-8H?L/Z-WMR:/B3K5^^&E.NQ+M;VS@X#EH?/dc9V1\V2)JcA0/
RU,M?8O>?:7VLP\Pa-RULW)[4SX::QY3R_bM^4K49YYPL,R-7B\R7(d9]eFIEE4(
E,8NENP,>W.JE)SVH+VU3U^dEHg<>DOH,f4W,DYg:SP(;Z39gf[:gD?@,\RFZ=L<
egSCS:M3H^0SF0S4JH2;+K@_6?)(Z#)G^T(e._4S\8,LH-a.G3^CYOV6@+,:V^Q6
G,\7RaG4@.DX6DcQ>8H/8K99U[\B8gb-<1X5L0B90AG3OF@8H<3(TFN[SGJg6WIK
=V1O)b62cCL(b,:+K.;5IIU5g=P(beSIZcE[Yf8?&9?2OA?^+N\C,PQP(XbBeYKO
CM9W=HZd7?[\DBT+O5F[B)+D#2O9E_Zd3U=7g.RKM1EgT_U+:Rf;FPT+\[H3I)1G
d[gf7+#<(CG4,<8D8Aab+MAR2QbLG^,>7D3EO8X)P:#<NHEK[J>@7K.QDUVY2f>B
G.[ED;A[Q2<GH^)UQ&)CaJ&O#O@V;gRBCRJHa&#[)RPJ/(WD7([a:&9cD2WLKgJD
)6VbA(U)_DR(>1/IIAeH4X+5Vd=4#][K+SA1RR&JN;?PPNKe58)[c+f&FM2[1;12
K+gO&H=[+6,.93b+bF#1K7QNG4g6XP<]#eKV:LX3MT.6JTYR>2,^NE0D.Q<VD15@
H^RaL(8E.#[44D3Og:Jc)<IF.ag+0-f@,:0;S2&71MCYAf#;.24XHCe?WbRT[NA^
HWd?)W;?@435=SRKPUfQ1>GK><f>B<A;1U&aP0\UEVX5_/BRRMe6B.gf3-:S-1Y0
7L5ObM2[8\?3[dY(+BXf\V-M[,,G8YAVZ9c+MQ2BC7gV4^9F86-6#13;3P0T76.]
E8\FH]7+X\0W\JX7)3&O9aJ8Z\0d9E+UP;Z9R&X\B^Sf#^7NS:..Df))9=f58V\a
+=+bHV-61WeF:eSCa?@--E:C6a2;[2X\JIBW<V=>G&A;[AP]RFSVIO^:VIVP9LIW
4fDKe;/?K;6]M-/>/a-&59YWH,DZF+>2MTV>H2eH83&6&QC6SJ.2L;)bX0V2]&R]
a..WKUP14f>a+(J]U-JFI.E^]R/#H=+aFcQN[CQ\]^V[WB=I_]MV1^VbT>JZ)Mg7
)6#C/\-a&Q&OMa=NDFZ4F1?-]@4I6R6)d)^U0/#(]QT<?@T(P02bTAZWTZg9d@E=
SMCe3bLRb<_Dc9ed6Z_fV7/F6.d?I;aaO]GC[GP)KZaC)13)4aG15,Ob(GS(Lg-=
41T]T/?1AcI-:]b:,)_:KQ?VE<HFfe2/6:[Cd.TA[g>44EQ95AfE_@d/4W1:?5&\
2VW:_/)MJY.f1&ZCD6^4)3=^EFaVSf(LGO:A=cNcOACe)E14<RC+d4ZIE)T6fI=0
CJGaH_8OV#\.Gb8A1cLLg\PQ/9PXKc/D6?Gc(f#-QB?SQ_?e-,NIXHN5U/1J7^#f
1Z\SB22N[K,Y_QJ/OGV29DfGRPB@RGELA8+^T-],gE8+/X9fK=NH>2g@9Z^.(+8Y
:.G+3)E47SBfXP?XM:c2Ngb(RfI8a.@Z+c;Q7-b[.&ELCLZ8OGJ9<7-227cbWd5=
;+>N3HgaWZcF/(Q(]R=]bQ,F0.C.TGE.K=J1O0Cea-+W1T]ZUF(SA<@Z257[2[43
((80FK2Gc=J[K2aD;PO9E&)a9^QPFY-NK6f36U+2DgBZPE=CD1W^J&DP(-+]cBFJ
+RCLc[E1dZ\Mg?\aTNDMVZDL0dfd+JNad1+;ebK&(_WH3764:2U[OTP])4\9<ZJ.
b?0+dRcO]aC8WdMWSDCJ4eS+E2bcN&.SH7QVDV_HW-C]?)P^BdcGF]2O#.9E6U00
GFXPf&#gG(9A?[S44[>Xd([gf[IZMN,HKbK]R?+PEWX,CHD@0DW78]YQH]YJ8cR2
Tb@:A>+OLIeXKcg&W.S2P6PdV+Bg_^/OET/;2SI)9GMQYb;,R>11d<]_I^d+4g:]
[ZS>V33@.+56_.6\cB=e06^cNP@LGS[(4f(&NR(N0PR@XS@.a(BeGLb8UZbG[TI]
cfA@/\Eb<=E-EMbR#L0E&<3gF.308Hd-b5(V\/4Y+5O,dZWX+S>[&)2385KHMO.=
ab.XDOf@BgX8+U&UP.62bVf]N=fXFLO8RE>;OaN7LZK>8A:6JFH)3XS:g;9P_6,,
SJL=AE+1W82[=dPZ]73FRQ.H5@##62^#K3PM(YgXbR9LU.]J7f/:^\RO_B9Q&/If
\Y5f-g0KY3Mg?W/@ET#</976+;JB\D#FbI4,,c1Y=-S)-^VF2(7J7O]d2-\#]]SJ
_?=\OKg,46+>f=DL5g>3-I_bVHT@AfG/8W<87DR,TVZJ>-bg)UW]Af8V#a6=S]bg
A>)3@I.5]VP<UD0WO+Z=\BM@8;;#>C1<=BY&6]D&4>4[H04;=2##?GK>68ECR27,
f_X(_d[Xg8-b;Eb1PXQ&R0dAL-8#M(L=QNL>E<8D+)NM1SQL_6H(U8f(4S-Y;8:Q
Ig4[[]Obg0g\f=K0>e7GC5+G-7=>ZNE8PW_KbKWV<IG.>)RF;EEN\95[W(+-B.ZE
/;V&_(]gL.C6ILX.SI;H^:SR>JQ.60#S_65;:EW:AV/_WS\.d(@Z&Uc6dT&N;J2W
gTe8b1b[(3M0)G3aeFNCE:BNSg9)d<9VR.7?@4gOE:H4I.<fSJc@9d2V_e?YWfc^
DM;\PU(3)9ObR0V@#2K_D@-B/^G\@U^39J?5d+?eRBb4X];@Pb+XXdG9DUF/5Z8-
GMAd@46Qa_P]FeW)eFP?)fLeb[2441I-&WC+EX&ER>(O0@1RL33AdYIQaMdG<7G)
+_IL2JPV+:G>9:AUWG]MM@&.)HKM:QO25DGJ\T+ET#C#6N3-\AS-?52J8215AaX&
(:T3b.](Y2//9f]S#d[.YcL7[DL;P/RaMP)eW56M3Y=.PGMVNaDF-G,UOLU9fE]/
=8@OOa32(QC\_ZI-2U^#496V48UC&\0\MPdT8N7RKA:)d(0ebcE@HZd(73<Z8TA@
T01]R_[dBHdaC=?_3OKN+752A_(dUQSAGIW(TS?K5K,FCa[gYQ5T9-b_ES4d^c[-
E0AII@2?_@9g-GO1N23X=77(+9V5DWW;6T)FSbfc?f^A>^I4?I?\#bea9eCQLL^+
36V-b8<Q@7D0Y]4=0^A(=P\?TcBH>-X,.S5cR?ROC;&VZOY+Z_dVQaAHG,Y8>UXA
ceF.bfWa)Bf>@6(^F6)[UL/G]H15bbMUZYSDA4I7/EIEg8]8:\IATMF:(5-84/S)
J8-PQMKL=W.,ec#/?[[5fZ:?SE5dTZ,/R8U>6)#[Q(N)^6=8JPC(#4=1Pe>-2IVV
R\b,.A/U2UXgPT#f-a\e3;]ZJ]XY802RW01M]WCYJCa4W63a7&(S(/7FUPA=49U=
X8^<RQ^Z9+CYAUF0X@53<-#4J66&Y,;BB.(bY8:f(I]dfX7^g1HOf+>[)G8<F(>P
DX(?3@OSS0J^.U:Y>,PN3RG+RS)>)0.5KZ&P7UQF@C+BC;H62R;9,P)&QY5V411J
L?[J-M19SRSFK2W60/.TGdL6g>=W-faV<FLM57(N/N._G8+N-OH]=?#;2_f,GaY3
+B6ER5-I3A[N8F,2ecY0)KcM^H5PKRFQ;/_<S0Xb-&->[e6.YDE;]dBBB>RW-P3(
\g(VP8L#5-GaQS;?,E3)C4.SBNN&4(8\&^FRL)7)(R\9K1BRE_#(&VgXL+fge[4U
TV8OOIL3[_[NR@K+SJG)U?^dUMf(B,RE;eaga;QZ:b@#Q>eTeZ_E4O#6A\0g]^LY
?=e&3\4-bPXET5^HB<\,[-e9K)[8_f>HT14dOAFN)OFTN);PPNL6OU?f]/Z:=^RN
K<FTeFY+V3KVgf/FSg@b-YK,E3?(D46)VceCB3N/Oc(7DTgBA78-6G.,&HUQZH+D
KGTb(<4X.RH>9.?5(0/AY5,9LY+<0X;a9?BUJXIXKf),9D+[Oc3GQYY@._\ZU,J\
I((;b6W(:@A6ZPcDUQ&eTDMA#=XV&O3e@;^EUCf5.[EU]Hd_W2=K7IY58^95FWLN
[]?[c7LZ66WeJ=#Jf0/CGVdg&7]GA^dP-M\gI)bPE>A[H4J7R@]2ZcQ,QdLUa:24
C3AR2K>[BdVS-:KObd&8I-+2KG:dQM0UVS</g18/N[E/Z7+;>TJDf)ZPHNg&ST>O
P/5U7bCXS&FM&bHCYL#c2UQ3^;E^^E05ZD^VAO^-LVC0WFGZE<X^.L/eO(+JC]GY
/JVI&&>0fCG4b05[<F:9OPJK;5YRG3MFT6&X[D)B4\9NW.DH5[\b7QQ(0c/N)&7=
=556-?_Eg\34L3?FO\#[Hf1JD+JSYX\9HV9cR9GZ]_Z(c?3L-.0-[10MEU@Md7W4
MAD\H3aVGS(SLV]SPZ7D9IWLgW#:_K(#Z\.CM7YPQ.]8Z[H+DaS#_G-:PM/a.5??
J+fCH6aQY,:Zf:ZK>TB1-#PY&CRE-(NM-KT^]+NZBW0Ne[/1W:48VZ#bE)78_>?Z
_<#6/d6RIWC^Y4[8PBY7=3CJ[K=VfQM@T.f@QRUaH\Z:WPI[fH#LS?,Ob+M,I21>
Q8Z8HYI,Lf[E3CR509bfP;W5ZgM9VAdP@)<Sa1\S0eQS41-VO9MX-FIYJ3M\+P#?
faA3JNQKde]5[7&>Xf4<N>)\JLWfU11TcG:I^I+P#6FTW@SLV[RJ@b23&fUIVYQ<
JX(fDeZ6V0>W3CXJKE_1PP2eeQUP.+I3d;-WA2La0F4F0_f=aIYI,P8)7?@W<N7J
U=bZJ6b1.PcZ0./MHJE9HT)+),gWO2:c8;)#ZB.Y#6R\;^b.G62WW&KaE/E/A999
Q8fO5[/^d.\R4K25da#IW2b=8a]cV(+D(+e<.5JXTLD\f7P(K6[D?^(DK;#+PK:E
DI5TU_;^-?MLe&?(E?AK+ZD]Z3:dLg-(W=N@F[R\.WYU55dL_7CQUSg,Rb8]0,fB
e7E7,B+(65.Te_F>f46F=Qd9(9?DME(M8dc)325J0/?V6X;#)U5HBSCQe1K)K5D&
GI3IES\0?ZbYZE2VC^Ja0)bXLM]]?BR?&I6NFAgM-b;>FS7D.<56P6<7)>?3.2[[
H&>^Y=A3LQ6M8)T]J=g/W_91-:4e=C,;Q:?@c[(L\LI&6,Ce>5AE@P^-DIQ4<(HM
,D&R^X&JH/D>c3CZ=/^C\VV3c3#A;g7<Lg84RQ;)X2fQ5]WV9eYe05e]0>1]aULR
&.1Z0>;UQ6#YAQL0GOS#?BTI)SP84DWfG.YJd-M1eN>:>?U?UCJ:KRH=YBFYA3-e
[K3C/_^8J^FY8@]?HK<=Fd;g>-1\AWWJ(N^D5;Y-[K.cAN,H=K2[BZGX(5LE-5EE
+HbD6JW0D,bONRIGLJcg((]^/fNL)eRQHS41NPM6K5Y[HUZ7RgQe.25\,]BfER4T
D#H3XS4f-a8G9SHSFbB[CFGR8d_8H^?gfA7d2B?:LMYM\UW0Z8#TO4a+QfccDeXT
fJIZH,GQgUD>d?T[P4JMQc,C2M989O^.[FWT@9T_,S]/EO+G-C2Y_NGeR68de]J7
TEZ.UQcC#2]@Z/U,\Y6eMZ\=QWXM[:95@3_R?MHA[GM544R7[0C9da^PSPfS+RdE
+,@g)J3)BMOJ4a0BXYRb-IS^._dJ<SeE^;DO^9J&?YDE^1+3_PT-UYFed[M41\A2
FbN^T,<)N6DNUNQQfY,]V?3+aa]==W1&4PA4T4ZdUfb@:/@1C60aaNIde[Ab36/:
KJE53A?CWFWIRY(U_7],>?TVd4+AY0CQVe:C7QZU7:IR\F)GX0S8=e:_A?7\;^b]
R.,EKZVV_H.DZAQM0)+c@GNVQHT<ceA)g+IAdG4M:>CO1UI\Ub1PX7e3C>dP_EUL
4UZO>/-QJ(6E9IE><JCB>I\W5-EK2TAFeNG6F^M/-7>9M-7afW6JJNZMI(BEI5cX
e(HJX8SVTKG-^N1N()I#M:T3GM/IYP+6W@YJ;#:<c?2T7B:b.84^1GQ)86NZD]/=
@#fHQS#F@g_cO&DG\Ne)>_W3)+/;XC7;[\V[S7,M]G0Y#LFIGFMg#46SO?D_\3X.
e]=c;M23E7Q#&=DY^_e;R.XNI,_g&VZ;IbLP9,0131?(G\\VNXS.^a1A25RT2:9F
92La2R;fZP:gF-ROdA-GQdQ>VB#SVNWD<fHSUVUM&0fP1R_TYNJ5F5K73g@cU(44
&Z4Va2Z:F40,eP();:,8GS5D.[B&55L3?Hf1>_NYEC^5<Z2WK+g_,RNL^0ZX-(27
-P\RV<bO6HO=GV6f@Z\g[R)8S28DHOdE3GCJFH;.@;bAGF07L#)cU^8A>PfM#HE+
>c+NRg<A2eC[YbZ;7I[AHU]U9Hg#-bIIS#;ODH3Z8,.FK?0Q4O,KW-4@dRQfP5@,
NV,H3WN:@.A3F\#a;?#I6XZ?_6PX\DF]W7N[D<VDdKY[>>Q;g9,IZX.NQCcBgBE[
AT33fA>3OHLIR/S115@DWDY2Y8&c=K;Z+<U2AS92BbA3:?.K,eIEL_@SFV7PL1\;
1I[aLa_3J<RC1/8H6B<.U;9-fCB:>\M+^GUT5@&Xf1OgQ78CY3=_c+fVA[UaWd#X
&/?@..G+RO2M#O([93@&D28FS-^N;^f;QX^Vc8be&Uc:Sc>X)X_S1KPgYMSJdJ7\
ZRT(Sd@F5S[SVOX21DQICI8aK.4SMbD>G:cJM/^)cGIJ9e\BCMD(N2&1G0//fRe,
d/^4WP?]PUF]ZTR_I7=H9[H;/B#8=?bMKRLPT,I1U^I&9P86Y>PMc&]ZI2,6^]XP
;eUc&]3:dOL@-_F5&b/51OQN>dNW-Ma:Xb)_E:I\=][BKQQ>VHJTI3@Oe&:P_(6,
0=.?5BF)a:[bX]Q;ef/-G_fR-(^eQ_ZB70SH&M:LP?64AO;G7OZ3Jg4)Xc<M30?:
cT1[Z/PO<\Se_bLHY7=fLGMENC^?QHLW/F4c);HU7KJe[CcW+?a=@C\X)Y-J&2XJ
YZ]5TE=P(BM<V7XZc^XA,7C<_F/21T7ff&&HJD#>g+gHCaLAg:\SH_@8^DdI2X_W
b\6D_26<4.BOb^b=4).#HKU/KZN)JQAAd=EaHD3T66VfW@0C4O?Jc&8Zc@af9^VP
V&Z>75EeL4<7/8LQDB(WA9Y?U\YdRWKK9B,XCZ5\C+Je&8@2T,=U[5W-^SN4.M1f
1#I.HPT-)Y^4ecXBKFBC[(VXKZLUO\,\7=d#JceF\>0b86R:;N6d322Y=_H9[CYH
\/UC:0+84,EePH&ZFf>&CBEaTc7/bc0Yd^bN,#\Cd\GL.\cUJRSS/5J#9/^-<+-+
;gJ,&L6;eMeT:e+^Ja0GDJNWdI_<&;><#^.2/SAeD#)JP1ILcfP78AG7^I91)+2R
MT:[FMX>fY3-b,GWP93IeX\NR\Z<?QfeYCV9\L1RFW;a-;D185VO_)Sf?OE#-]DA
AfKLSB3A474K,[WS<Q3_7QA1S1YO8He8adF/9T:\Qa&,a+9gIJ^f>0<T1;3:T40G
<9=(SJI]^6XFT-eWN/JTd)/E?^F\;;a>2N3UK<Q8b_^IWF.^BUfDH]+>2Ad@ad9&
\OKAd:+YU]4\-I6N:?<M)]fK:93EFHRfIY]3Ac?6cdP[?2I54OZ-[U;:#=L];1^U
WAJ)T;C6,U1;43HdPc\<),K;c(_=)KF2C:LMCFVQ>G<2E=3[-VX=/?Z:U\D<?.,3
V5\dI#DF@_Z4CJ^XX/S_#(ZQVM4^^ZAaU2QYSLWH?I8_5D5gW?+9KLM(H=AgDARg
<:d;CRaBVCeOPROT94dFPDTE@=0)6[G17,JfE74)R29/V.WR2I(D:S1,SMZdK,g1
WAOU?1&W&P1Kbaf5@Q0<9XafGT>K@(S<e=cAMG+FDCVf[Zed7&RWE.VR#A3Y,aHR
I:IQEHc2E+<#LH>gXNY#A?8BR86]@KR+9+2S^7G:MEb>SKZP4g.VRTaP5S0@<6c7
3@QV=N&e6g1a_VV6(YO/@e>+F0EM[WC_J/f-88edHA:07R<I:UB^U\^-+.4Y5O^+
VO7V31@]2R23;b?4=;&fb/QJ(a#,IbTf#QZ@VMPU(f6.7>/;PRWDUeP1K,92M7OD
@27Y82e90V6.dV0HeI;(1Y1M5;/GBZ2ZIFM+),GP=e?+dU_98(A7H\S1N(dYLXPQ
QY2:VXR+L6YV^b7R@\fM_U7C7;=UW?@b5NY4AD?U8WTE=Y<6V/G;1A>_WfY75Kb1
I4OCHcN4KR:d3QOOB2/6\Cd/=X.^]G<2V3S/0B5&-82W((#0AbAYbHN3fFCaP3R]
]DfQN+;g9&[#WTE/WZ3VNDS]d-36_<d=IGCDbC\cI)Y.7O^V3dVA05GQZgF\A;,?
)]^Wg_M##fBT_ZX910eR#B<9_b)4DIB#(L,HG?E4@A)FQH4V58T8^H2[A1e1bFcd
1;(Q)#g55WPNW<9HPFXd1GVfY_3F11[VM1&R122>D:fJEF9WSM36+K\&:P,F/9-?
\ZG)=>\@L^\S,FH@L#H+TSNEUV,0U\I]M=AUWD#8PSU\b[9MgR-eaG+V;AQ.>b[Y
ATUH):aUFM5C6_I1/=W\VdgPYcYS?#Ta7YV^V&C(AIb)Ma;#U/3^R]Q6I6UZP4gY
P7A:USHS&M^cK0,&>?3b.:WVW7Z(6a/=;HZPL^09.F@PR]K@?O)2H=LGQ+0J9e0B
WYHXM_L/1LMXcHaH^]:3U;>Md60g(+N8Q2?e7_A\FV.3&O;&FV;K:W>28_7]ffe<
g?4QCX7C:Z]-fScZ_E^JN8fM:ZVbeV_5<3g^3^FBPJ.BLOc<5Z3C?YB,I8<P..3O
PJ&AG;>WLG^Wc1^M7,&M&(.SN8g)689ca5K,3+5LJFb_0f-L1KcY4ZQ7d?TZY&6d
?&L2D\AdQR#8eOX6cYJd02:TI,f:#1X1;4b91/)Z=eG6fcIRT+-7CK=5[CQIMW3G
dXdR]D(#XNLYP#7A_,WWHXc&6,G6:CVS@J8/KbSdAVK:&@>gI^I=Y/-3^(O>;3gC
BOK.XL-I@VTD:^(5OU4N6ESUK:)\<=HSTO-S.g-Y;#?=MX2D&3LNab5)00@a=YNC
KPO7RAD-_fg\LZf32d9+X<d;MCSa26H8[GWQf&J:+_^Z7(9U:bJ0dVG7<0&H^:M/
C7-H\8H)WbA&<T,/7IH&N=XAgScd2VCBEeb(eCL&#.3F?XYg/3,FC8^PHPd.9cfJ
N,4T+GP)1RaM6R(\1H&1G#[++7>X<C@#c<Zg:><M,CGLZg>Z_^ceZ\1MIegXBVe#
S1EdD++d+2M<Y8X3N+HL9N5W>/Oea=,Tb]b6C^,bS^]J2@\-+5@]AO?Z>A\MSb(.
E+,Qb.O<2aPE\5;aC7Y\43.QZ#AEY#/c;^_GK4f3NG[,N),.7SgcGZ5&@]@,=eeD
G55ONDZ)eV?Q12)fNPTTO8a-AUHUZHHe/D=+A4#6Z-be@d.C/AT@Y=_]))ON-A8R
J7NQB/LD,4FVQNC>LB:I?YS4\QM#Rd&D=]T]]D+)S2@)LQ6B(WD88O_G0E=eH^69
TI/S+DEXR)dN7)L1L[HeZ@Y7H/U1?FX:.U:9/M_TXW1O89P+RJ&@4Q0/ZM^Z_RXM
gS4\Df[M\I5(C37P^:7>I)J=NZ=9a5Qa+&ZKDOOST;Vg;^1N3UR);W.MYBfgc_\,
OZcV2+_bb+#=eU>IC3d?F2H8KN6U@,bFa+5Y=W9-?dZVCBQd<\H3>Ya2H@A-Z\?@
3GG\cK;=YB8T@Sb-T<KVU;5S[?YSb>T:gGEWZ3a:#-+[-^P]b_SV6I(=OF(:K3F6
6gJ8H5a0?QgXQd77-\cK/-^732&VVBI?NIDZVRb2&=_U2CC)GZF1>5VHK/D;:HG\
]G#FG7=2,XFJ?M=SSdNKEV,HU3=acCS4(,#2b=29cc.(TY8&C40A#L;^aaFe.2A:
9:PH\.IY5LT/5[Dg3Nd[J8C60P2^M+U/UZIV3J=_5P7bRV+9Z>HOe@UafRMHG\f]
2De#^KSGG1dGQQN3QfJ.9<M=-Y1<;LNZ0c(K@fUEI-3;AgQ=J2aYP3_>\HE?B@_R
F#b_8M&2@BC-f0^,dTOM-GHg0=VgZcc[)T^&-,E3-S;:4.ab[\QMASDeE15M80-F
aeZGD]\B>M)INSPCNc8J1\A5-[0Ng&?Xf(LF(OQ<<LYQ0J+L5F&+5(aA:(bfA?1E
T):2?.LR2^NJaR_=^CDbfDT9DYNWd\EG)PV\8WMg;V):DdBdAA#)XEeRg&)\Jc5B
CC7F&T#WF[X48L<<JRcYL/HVPSG[]U+CUgEGZ?T1Z#9N^7ORd&/fO)We<)XK?N[W
84B_R(YPSb[+CYe\LeSQ6aF(H0?gPd&(]WT@[[&#ZLbe2)ga4Re(FIR+M\BQ=FA1
G,P24KSaJ87.1MURBNdH\_JZgDNE>NT98#DA8)M,eMcPZ3PeUfKG+UKW[N+#+N#7
(TC@HLgFQDd,T&[^bM4Q/[YKX]W;)bf+3,R<5RZcR_U^@&R&+5#0?ET;9:0b&BfJ
ZD20H1ZN.,\ABFA0\,@_DA_gV]MVM7@gf+JL_3\POM_K:;X;[aP,KeG#>\8bYaCQ
5&YF-ISc#b[AXFZ?>6#;6\c(dQE_<a.1K4.0e-aVXC0\]0:?5@.-RJW)H6=&,d#b
&LR2.GAZ;)]MOg==9[EYAdba4MQ2c8.PCF&ca./VVBeA\.a)7g4WN=]P;I?QYF.=
5LD0>,RCX^IaIF;\9J8LZHSGG>WK?.^17N,@<[Ib9&JW-cAOH-34;F(eVcX2505P
e&<,1>c9T1>_/2=V)90S[C9HY<)^_=7=MSY-E3U+M,09&gOKF8gVYIQ;7YXY[&2T
3+VFe3B2E?G1S][Ygb,Z?KW@2gJ@Q>@HM_4^V9;a>eT&2-E.?dbP^a-1B=J)J(QK
&TMY-&Z,>RA?Jec<87g@bQU9c1Bb8<.DZS8GVZ]9TO0:P^F-OU@^7Q,[JT>WCfG2
ZVVG&Z#_SLY?8A>L9695bHF?++7@A=720/>b##NJb_S90S_3?>18V@=EP=>9GF1S
L\8aF(FCceMcFPGRH36;bC3JcYSF&-.\N^O;UA7+V,D+F=R.8bYe^D,Z8A^]8GGP
GbCSU:-d:B44#XLbGBC+I;G<(N#U@1<4GCQ^<V?1>T4[4>S60<?/d8+IAV2\_Q2&
:4UP\&M\8&#f2(cY5G-dSR@A+&TQ>I^00^fVUd4cLL33bOfK[B(55RCcS(:beP1Z
g+d.3FJa((Q1N/SOdBZ9XP8P7G3CT])B\M;=gSI;fQfXNM/ggOb>>R43Veg)LAH_
EcI=S@3@g24-4^/,@<:[TR+LRg67QI<JHM_)aH^7]-=)=K)b&FZVD?J7IT?)7?NL
4EC7-1b&@bDFIANR9bUZRB^7B>&VQBM6Q&a(IM@]M1Q]G6>K9:)]W76gD,Z/7Z^4
IYJ]4;bD?HdE.V]\1XW7TFe0/>;aDZ[ME(H(BeGL^=<S/aD8?fb:FaA^3&;JYAgc
0aKO2ca;Ke)V@YVHB?O8HBPK]EEUDf@,^MEE\6X1eKc=@&MAB)?_=A[N;N\>O<WZ
+F<[b7f2cII,^)U6QAcQ+Ne_2b9bJJfR-6e1]QB^>BNf9da]TC4VG_c4WJ5E0;c3
XIRVW1F=//?3<>D+_[T&AcDQ66gVE+P>WGWX?EF3^U37?+P]2/ZbXcT^<BfY#+8@
CZC+I_7+OGQ_1=EXA01^3PZ<@[L\SCSOM366fc##&9bHX()_D?,^a.:KeBcXgGR<
N::WZ^6Za3TYY4IGCRW)5+bf:TN7D[G_9V69C,De9E(dP6fdL<&/A/^)12LXfPPX
=W,#VA\5UYfdBPM<J+J47Q-^?g)a?VN?P8KX4S(JZ?a(7U;M(8(N-63G\Y19f0#R
9GN+NHd7C;4N3_T@Y50^[]\BcQ)@8\2IXg[Q<g9AN5O)]4eb<=^[O^bCC/?0?1>D
KN#EB:AV^fM^@&[]c>KN?>c4\dH[cKfZ>)7&<.F>3gdW[Q1GE>]3Z=H<5O=D1WFd
M3YXdA_9OLgB2HGD&R8__YV(dKB/C6+&Y3F[/KXAR(7D12QYSaNGcAJ>?Y?2gF8.
=1#-R;BQF;\DN1gL&]2X^/A&2?:.I<Pa:0(C=)f/gC[+:g.82QM)HcKU-1]TVT4H
gWHAcZAL?:3_ZfX0ZS/?04gEb>WbFOA[UMC@<1fg\JO=EQT1f.897<B61PEf->_b
&cI3_)N>]DX<TODMc+8+cDWX+9NfRU\W[fO&c?<E#D7aK=PW5J2c\>LYg3\?T=JF
4bG0Y(L02fAa.K^[Yd04/I:VIF6^>^A9WYg5_Y8V+Sc5AZc45g_[.Z)7L(L96>QK
KE_ZZ_c)R549,WB6Q-_@Ra.2]8-M@M4W,QQD4R;b<fJMNWHaG<&FMTKWZV[IW)BU
LdJ(=?)>5>_(bN>W+50@-,TLS1We5./c6?g0XJgE07I#REDQ@?B#4M(]DAOJdgg^
2MD&_7GWeOdAIVKVfVM@T:V3(+<LMXOV2]=;HXN?f[GYeU/Ag[Mb0d,:PcF_LQcd
26&fe-CR;1^NCcUfLMe<+6E.=;P_aFM=SOVd0><(:_/MP;O@#7D@4?bcLY42f>E5
8HaC&YKTLDe7Fe6=:B6gC^J._LJAP>P\_]bN2/>ASVb7LH#3B@7;DGdd--+TIBfI
Ed/gMBH_2<AYf344ggL>XeE&?c:0F.&6,OfF#XUa:_g8U@P4>+NABcO7^1X2EA/W
Ta+HU=+gID3bf5<B[9.)c4H0FX6TZ[;N)],9JHZN6)Q-fV_3E/d,2CXOfe#RHAMV
KW,R3Q[DL_FBTM=)]&UW0@0Ff/C_L1GfK1,]dY_OSI^NCI/d=[g-YC=P3=0/_UO/
P,0U5>S^M8T&\07,\caN(Y7L:P<7f\/S_07E8C5Ud[[P97e/0]<(R+WQ\+G\M5+4
]5L3GPU?G][V;TcL0aL/((H#_7_O?_R:X?P&7M@cXU?#I_@<-.VJ(\e6/0TS(a4Y
#A8cRL#bL@VCSXG+ZCLC-YS@3f4:I5V^6cI6C-<SbV3:24BZ4K6Kg7MDE\83#U5W
8IAX]K&MN.^ed+d.If>AA\WIZP_YF_Z3dG@YGEIW[Y_EPE:EZA_e)K7T(85/+RSZ
QfQW:GQ>16[Bf?4fL(<92IAcX)].KLY\?XFM_A6EE./TM.<++KGCS^&KP:(#:2^M
0CRWCe[CXTJVXR)-gG8fIRLML9OVMB]&C,Pcc_7(ZARgd(e);QKOW2M9_QBN@(];
Y3A(:QEf(,V4K0S=2/:D85:&BVQ7FCR,.;1#VcVKZ;]73RO450=KW-Ub-fA+RO7B
DI&@/(0#KH;17<_U37IVUR9Ee)gSD6T^\V&+b?CO4/#faW1@F3\FSf_@JOfR#a>U
d+)gJ47aKL9@c3E&_<^c6+c(1WFS,d4X8BDJ@I9,fE0P\5#B4MgM=Ad)KB?-#Q/K
MZNZ,C#ebND]bW_W+XgXJ19[1dZHH4WK4/Eg2.Ub;MRc&@8K:dd.#=+U=Xa=K2HJ
GLKCH_OB\MFaEI9??,XQ;L26IAD56,KI>;LPZ7=DWIb1#Q4bD^&VOCMR5#F#M.Z<
2>R_c1D7._fRAG:N_dN.W2U&C+5fK]8=[Y[g)cd[e6MPa@V:]Sf5N9cg:<Ub].aG
\WP7/2X.L<I7,2]g5\[YEFDV7Of4+J&6([M2>/67(Gd\[?U&,3_MS)e_T=J)8.3;
\,U4TCSeS?MPT>c.N30D;M;\fMU8b-4:T&Z#Ec@+NLVS5J(N)@-ePS554359A66=
/E06@a]YG50H3?-Yd@BS&/&A@Af,6ZZ[@,2>LdPb,RDNFI7K)SDJNWA\.=<<]VZZ
IP1OH=Og[D560O/;/>)Q@FO^=QTE]aV0D+FZG](V#G8Ha6LFRR_B+^?I^XOI]D-F
?2Y3.I_dE+fRBY4a-DWZAJ1eF7T;58\ZGg7PIXBg\dLOCb^6I(c9G9C\f5D9H)4(
BZT]CI7GcK0.E&B8MWDTIcg(>J\L&0Z^Ze.O<#I.Ke^IYGIGU?GbDP1g+]V>V?R.
QGHOL#,GBRW.d=VJO8M7LP93.REWQf(HVTFU;0g;YP-(fKXW(Ha55[.GW2PUK>/V
M43/]TV:A@,ce@gG87MW)J(:3#FF(S8X.FR@7&R/RG.Z@\d\,+K+<-^Z1-6)03A-
N]FUQ[dYfa[>4M-cWM\TeZ#HFJ&eZ<G1B7A]L\6VK^dSXD<OgZOP+_DJCX90L77\
GH-=]gQI/SBX[9F-;[/#Sf)KAS@ILC]1,aZ)+,Bec/U)LVFT+ef)/E)0?[]>?U\)
KXX[1H/&A8D@aW.K<Y:B-T>,FEP&3?c=OJAYf0Ja;MA6#\,a\XJ++@A.cY2U-8C4
7K:OWFMgW/T_GfW0R>TH5_/g54I]2T(SgM\9N1P<LQ5226T=^I.JdEFQebg.fFRI
.R@O-SN0NJO7:^IYA,A7>JIK99^C;&He;7a3gJ/W_GHPe:-6,S\L(4Pe<@\IXK[.
g&^G3)?5R0+.V\C\-#L>YSJCaA4#-T7CZSd_I8I(3[(XD:]\J/ZB43>Q4J8>[(=8
9aC[?AD\X#?NF]bF:eLV/\0;3YK:3;cBZ;c<7]b.+8^OH.SCTG)[b@R@:#QME1NS
daBRO3^GXDa::LLUb9CDDdga;&?E/LbSQQ5\O\R#?H\I?;@YO+FI+VRZ2X<+].9\
A^AI9]82RS<^8@0CYb6@OggXXZ.@QW+7AIIe\>SdQUK17D:Q(-F6XPaDU&_HH2?W
K)JDQ#eOUX>UFGD/Jc[BML+4O?PL9#L#JY2SOGb60=6\?RR&[b.]1PcKPA3AK6P5
\R-)<Ea2G7IT/IQ@.44TF;=EI7eK0(b-IgM,0-,V9+^:W(P+_N0H_3,-4gTJg83B
\\-1YDJ0eAJ)T/YV)ed[1RLO,68VR-RZ[2U3dW>B;_C5;FYR+&1Y[5=8HGY9:\JN
</R.4C#ZO=ZW1]Id)PA<<:e?34IL2R[()C>e[?4T&,A41A..R1JV6/P2P037#K3D
:-.Z4Y4>=@=F)TN>GNaX=Qd)-I@;9?caPW4]-;_Cg#D^&A@>Og\fe>>0X[PEGZY[
=R3&KD4W=>S3U^YN7G<0Z[RN0aX2FDIAN7A))1I>M#MTPC;@Zf+9ZY,C2D/c7<N@
KF[\TGR<&c1KSGCCL0IC;N:dH8G+:KZFF]F^/,J,eI->B\4-cXK#>N4(LUG[3])3
TQdX)6@aa^CJ\AEW_V1TPC/G4cSc)4<ad9&_>B]HH3<]ZO?.ORC<_^gSOBdbFg9M
cC5=VW@R5@U\#L7FG-d2:b-D[fTT0[]<@I<HX+]]C8AdeBB/F^2HU13A^[#/C@be
(9_B?]2RCb<E5Y\QbUZ/ZE,:gDRc_]\agB#IAAXI84Yg(42&,V=ZbOOL:VSINZAa
aUIAC422\5?@62:QQS]#-cO3g,d4aZF5f#\b;Q(2BS=Y:\[)@T1fQCOLbI#gOa>O
&;PdV25U^=1_HM#N2&#:B)=f_((@(/5=d@J--R81GD+3](EVD?^3>(L@)3-U0+V:
bKHfd[^^a(NRHI3LBAUc8=QMR7M.=,#FXNeKE9I+_Q=[3:/.2@F;&6?-2,;Vg18[
-&OU=2c(B/eR\8?G2Recbae_#2Hg4_cbD3^^]RdHDH+#,.<ZQ2.cbYUIS(8ggL6[
Yb1=393)f6/&-0VdW.;GEEEBbNgbT4C[UgOCSWMa69C_=Z=P1D<MQ79?V]7KKX+C
5^GfPKJ6=92Y:4?73&DXbY8L(SCY1-0fW1/S^a.9SGT5&b+2.89S]#<,;8GU;8:_
#T&_)4ICA_(U6cRe7S48PF4c>>BaGI+L7Q7.-SC&[9M0J+J:S+],3+&TDc5PSOe;
C4.;]&)OMFQGbS^KB(^>L_KA=H)G_3_[.8UMNX8(]F7UH+)b\WTYKIfIUEZ3)NJW
94K]=R^A3KR13R3H_+7ZG87SG[cA0b((JX<#43Qf=\HK6@d5LOP=gN,KS[&Z0/A.
C8+]=)f?)WLK5R&C;^g4De52(7?7E0CO-,VO+.V.MZ/.0560b\\-ZJ^BQHZ?V0GK
B=C.B(8Ua^(#M=O7KJ])=9CIPYH8EKZWG_>Se5.@0&M&E.^@9eQ3123L-+NUCA76
2N^,?gK?[+M,ZGC3RWWS_G3IE\HY#\HSQ;,65HD[\<4D=BZ0+H.H)2U38QWOVN;[
&YR1Y#7I\M1eS[_d.57P:d1Ta[Q5=J&XRW[+?D44O>OIS;O1+E134@d&REZU^?4^
e/R<ZQJT\gZ2T+A>A@8>KU5Q5\<WC(JeU,S69T6;3[d^KRJ]6D2D;0/dSN\g1SMI
Y,KAKLSFHM0bURd8a2.d^bUf+BB;9,04;/TSMb&YJO2,Ddg4^?:a0TWJPMB]AC-E
[YR692HXWg-KW?+.Q;-,@;.5b)>C+bXg/18+4aSB2JHFY?.#,_YR[H/1.)cT;.\g
I/dRA@7=Q2@5,(#H,bBBbR1dcgJPH@SEZ;J,)8&P??7P_aQ(?CFR?K@B^/.X0H6R
b6\D8B&WZ:0/.4?_\3_4YH1;TXd_=[>;G#8T1&<T6C6EXHKH0UaaCX6>5[C#gMDD
<LW2+^>=E.=M-U7EZDT3:2LI)G/<&JLX18dHd14;:e#F-4N)/#C]a/=5-A4&f=K(
]@^O<2f0(@J&1EDDP#R4-0^:M2E/;^L06e+^Y_(TZWa8)=2+:8U[KG:O@WOaN@[D
X.Mc5SIQ^T@Kbf](G=,UF_:1_]7_-[@DK[e\XEKU>E<CTZ\gV2C6E[Z:(,#^E&^A
Q6<Q13(8/2Q)2;c_O8a]E^(V@UeIL\32_VgQPg]>XFDJg&)/04SS;_ZWaBV.)C64
E,GW[2[=S[+\ReM(:F#74Z0Y_<H;W3&a#H:9^NV/T<U^AU]+0-20?bZI8R68(+SB
)=F8E.9NQ+:IM0R\.0#VW2DA^T-0CFJN)5@52d&6VV[d^9+5^V;(Ab\X5SW>K;7Z
IXb_d+&+)Tb_f4.[FFW^#/eZ/.M=#c^.b95B[U6faMc-D-4:ZM-@E?#W^P6&?4NU
\M?ONK4D30N\?NAa(7ES)Wd\[?R7KPHIPXf[_7YE<Y\@C^W(?Y7fMASD,4e#\I#3
TQ-?>([F1-F:TB()Cf>.b8cNCR]ae<cd\BK5KbU#dd;ffBQ<8H.LaD\LOc;_CeKN
>Za\U>CSA>[4H;3cXbAO-DF&^BRf1EYC=))91GVFPD--B0_3E8EQK,c;#c\>-[JB
Jg8T1+JZ,3XT^V\/PI4P510]<LL4Bg^5gdM0?^F8J@TMG70X+=fbN<:/ba(JBD4?
Q0_Fe/UQ/>ND(45-O[7DB1;^=B6_<gL[7.KWeV&U(59cg)cO0,EZFNGDKgZ;LHJR
RfJ&ES0LULQ1EP\BS1Nb?RX7Ac])/&#HVBWCK0Z+C;5-W67<cbe>UQ#QG5YdF5_;
6O>(d?R/804[QBB#R&F29KZ<W1/[2>HCMLd=g8B7IV<5]M3RVNF2BfZVg3(54#?C
V=(+H9aeR=6;UC<7.>N^MX9)R5\e5-F#6af+H?8J+]-&6+-.DCa1BDR_05B>dDLP
DM9>;G(5(F&.KF/?O0H1?c.gE)N?cC][5+D,H1Bd3f]G#391J1][>[6,O/]3B0K=
>SJf]],VgRFR3.MF+75a+PDREN[BG)C+U^OQ6O./;0,1\T84C&XA)U7N>^BVg+?+
>/;D,Q<S]2&JV(>8H9]a;dg(LY4,LIV6@9@OHeB1eD-8QP_<5[=(@d:98-W(<2WM
O-JRYA1=S[@eV-2Df1-M0d>2IZNH,[T]N[Ld)C/9M,S-?eKP/5B5<D2@,PFaZS@A
VYP>FW-0N3CTCJ[B]cY0:,@9FT.J)BIXI@aS31dHF0b>@Y&S?0J>JMQMTGa,0TM,
e&-JeTPZM><[-2898I8)bfGU02JD->:Yg&[3Q0S]F:7V[JWU:?__Jb&dI1e;)->G
2_aW[BV[7T_DX[,f?:UAeKZd+bKcCCK,HJT0E1+3=.SHL]HOf,VgZY&0;^f8aHSU
BT,FG9)5<HD<85)7c&7:eD8>HAM)7I[W<)E-U^Rd2(T;I0\?d9-cb0EI,<aPH-N8
Q87=&LZ3/>T?Ea>K[X9@<YC5>1W_G3>,2I\TI]KPgKK>PGFZ<+Y\LS_1+GWaO5OU
3;2YKLSHO2UG_L_>^B)aP--XENfPX56D/>U9J.:=P^Bb:_QFSC71ZJTF)2[;Ya^W
>R;ZOT;G^dGAOaJ[2<@E]2=Df,Q_</+YQ\-OU^WZ>6bF[>VJ?RfcGW_VA;c[A<]7
@+cS+N>@S_6Y59#<f>ac<][5[gU3Z4@#ET>cN(?H=3@K=EHWVB]OS&0Oa=?cF[N;
<>Q:QT@cF4S5#/5)<JK2=O5F&W6<:?206RQeE?9I;)/86@\8cIFFO<e&MHK._O9>
[N.:cSZ(Wf((]V>/6C&[/8Q\JaeOZ_]Ya<(B^IQcB@40@4Cf?_6K6)#HID+-fK0a
2NXB53Be4BEfc1XQ146XC\&&fG\1B(5D(BPGE^<bcHV:H8=ZBHLZNLdT2OCS7L6]
NbP)HCR,CX(GeGIC>BOC16@R^3G1-4(@ZU;-8)-cNBG7L5TH/20&A(^E@8QDgB]F
+S6P&^PUI,JP.AN9Q#?-aeTQ;OZe0?RZNSR4B:,cYW1cD>XU?LZ:#NdTE4cIUWdb
L[6YGOWDYf,M284G2LFM<ASJJRN^71d72C[bc./=bA8A?U<KVG6Ib\@1IUd.NUKM
[HEdcab[Gff4=fS4S&DVM@T\HFS,ZdB8/B^f?I^[(VK\SAR\N)MgdEIMZWOa\-9[
WgI6@0Z9ZAM3?/;\fd24<;?bZ\&ZAG9OXOLE9XQ)2336AbYH26b[C?eXZ(S9\I0)
G,[HIZ#SU^;W#).G#aRa,=c>T_(;>;Y9g(aK;Tc5/RM4-+bb/6AKBZ+T[-MR+4R,
@444_5+4,5f]gf4&K;:Y&f(dZ\N3R57I\a^:FgV_^IfFS563[a<0]^D\K;ZZN07@
I5cMK#3=5gDYeGaJ5fL?AUC5(FZWTG@TQ8.E5PH&2&N?IbNOWXBO]2QI;W>6,(@2
TPI?95LbgX,8.#fQ_XA:\0;YCCDV1V/;Jeb8)74>,VW<GN^794(([G7+R4O<4ef5
KT+e1/N6;V7BOMMVK0V;#O0QL).^)22UHgXZVZOO30;J]gcWXfd75N-H4beM1caM
;LI9]@V^HXg72J>G&(B42RaRf>DV3+1IFR+2Z>_=#\37AC^[Qcb)cBPR_P>V;M(8
(N)1b(U&C,&]9fMNXWb]MV<JHeKF4SUX[L0M1JF;1T&2fLWfRgWQ>[^]0fMWc.^2
f2c;K;Z]8YOT2dDB++b;]?dA=TBW[JWLQJbF1U5.EM80[7E4[@bXVI9#EYF\-3?B
FB(.3IFITSXS3H>CSd5T47_[,>V#[LXW9\+/HM4.]ad8&LdB].TE1Y;<O^&RIgb6
]A]20[>&<fI>U[4UC1]53(<a1LWL@?e:-SVA&bZM(2G5#APHQROL5g8eL+_\VCX.
/EF=3d<QP=6G_FZF/C,Z3.2LKFe@HfDRe;US:(K;;6HPdMONH/(HG4<X.ANCBRIe
:3E70JJX27?433OOG+FK,LYF\@fGJ^[4a,YHdL;)cF5Y&9UP]:f&<HXA=X=-S-fc
caaf9\bQV/7ZQ24XWe\G;+TeYUB#=?7T)J;A4BSKEQL0-;/,U(_dY]bY>W;@3Hg,
08N8=EfWSH[_-O\a^#C#(;6;V82IQU8af=^+[JKNV]1;@SeQDO;D7Z,WDCS,7N-G
ONSL?\=OI:^2gfAc.4)E/,QUdV61VAJI+MF06+9Z=</D<ND9G7>f0_5-=Yf?6fAK
PgSe9N&V[MY+2<ec?e&(4C(,GQNGXX159G&>3+a)FBH.aR@(Ge/:/-H?eA^G61-S
6?/.-a=\(/V&KF=&T0Pc+J_H/e9JaN(IS<49:5L1f^P5Sg9:1>BfPNK59Y<^J;MD
/T0\+L;ZAYe4ND?NS:O>Y/eO?MQ@_0#(>JOF(HWGP#P2<Ag@.Z8AaR[aH&aDL2>X
3_L2M,bE+B>Yb\8a=;0(69^b=CI2:^O^-H;Y/RY]>3IN/e]UAL\5QV=/5>D#:O9F
:N_#f8,X@]QO.dKcM34?H@Q.?APX^gYX0QNCC-]66KN@J9J],5,b,:AJ>3V/(=[V
O#I4<bCJPea)L:(bO[^/(\6:A^2UF2Rd0fABgC^[5UPFNgSNWe4LaILC>gL6CD;,
/_437O,M40\(8:-WPe?\:a/;<U8\_FE&b9_FFZ(;TI:ZO^R_Y9GV?.2CE:1?/:M/
R-gX.+_QNKgG37+J2GTJ-@O+F9_&dNAMg&OZ(Oa]U?8K]5=PC)4[bKWZF1U(G577
-<]-G[&BY>:S8;U6#6A<a-R;@a[;Ke_Q]e<4La;?=;5P>VRPC6;P3+2.g@,I<IaH
914T^>>4]6bO&Q4_59+.M6d]IXdJJTA=VBf?EC7V8)F#O&L9aa2[Z[c[J\RAe+F+
V4_&Bg-9&aQ>OW;84BRdIYTfDFBVG)+0[Y@I7^_gb7@/.<-AeZc^=G8.Xf;HB)N2
WC.E=#:+5\WL\NW:f<-bde#@&U&D2C,@b<V8MY=55N4867_3;IOKVZSH47fEMS3:
A8X+LQN:Db>dG5Q475G,2CNYS<Y:18)Z)])eD<W#8\=Kb^6.3a7:c\GSAcNV-HW[
U6G_H.PMV2YWf6BYXQ@EF<[?U,S5)?BbVTCY=-F?OE[Dg,RR??TeY5J&d^MfVAdG
7B.E1b\B:0eVMg?Y>7^RK)\=DN:AX9:0BRIVJ==G7H4Q#MH/<.@d\=.X(,=c2K1d
,4<<DN?9NB,bTI1.[X?-(@7GWNaQaE>XSWHYdX3,OP>2.A@MRN,31\AVfPa8:1BS
5>M0JHJCe53/#^bgQM2.)UO,cG2^EK]V?CAI3^W4fQ+&5US43VHF8VQ8^>8aJ_=N
;)K=Z;=Bf,&cT#XG@bP8\e2LBMX=:5bS^_/OWFVIJF9_)M7,[8HcU+;QZ;BO5Vc@
8dBG##[Z1+8Y4_AGGK)2R[D=YK@EM3Gfa7S?Qb]9UB\R&[LYW\#JG:RX-M=?^gU1
M1+6)Pb_YNOFB3EV[ZQT,F?IXDJD>Q+#LEM8YV]2S_Yb72LO8I+/RE9DDQ@\,Z0B
SV&+)2R05BZ0@=50?K=eI1\g->)fUM8fR]a[CYe]H>g/DeXO_)0U43:KP,S[d:KC
?U.L]?C/JHTJKQWYc6_M6H5?YaU14IaaRL_CRc>O1.2c>L<?A=M;DBWKb(fDbf4N
aM:+A30Z8D_c7VXQS=M;da@C,_ga4;([<(0]P(gE0_)SS:-f63^+#]5IBfWLae5[
b\ZFYAX#V)TFE?+8#INQ=/aA@P/A]K@UZ-M3cEKR/(=84./HM0NY?/NLa&K([0UH
FUZ[(GM5=BN^Hc,SJ-fdT#JdR]Md,g4MD5<Y65WfcL[@=5#e</GOa;^c&@21A#N&
7_TNFdGX4&DQ(B[BE#U9EO0=Ne1bTZAPY..XDa)D0ET__E7Q>X7X[X)#VI#XC2\6
F#[0\(]f0.575C)ae-Q^-;c3WaC;&/9Tc,-e]@P@M\cH)=Z&&I0[.2<6<g^;5J)d
Q5DfO4Ed=PV+a><FAHGXde./P1UBDd0If6W)cA[D6Z5bRHW&R\,(;g_L28PaD<.Q
HQTMC3b@,^J,^@9[F<FeGGd7Z?1[#2H96Z2J--/Qg2&SDUb;7-J?4.3R;A>RH&0(
.ROgPL.K.F+T,gFbY,:/9g<U_KbM;fa+FF7HHfP\NB,4TV9,SOK\R+.\_&@g:_]Z
^PcG1MZf=D>aU[f1-g/d;f.X2HM0&Z9>VFY06GF]\0[J#SQ0OG2<B&3:Qe+cRLZX
U,^IMJLTS33ZI9JSbZEIS,[>gDdEE)(+Z2D]f9K^V,9]7QLT1QbX(JYP8H;\IWGd
.W:3(>LT\KB/EaY[)^f(QKX]KPL/&<:c>YbB#fA#=;d1RBQ.S]#dOD:E50,cfOb0
/VbGe/+AZA+5-<NBJS.2C4D2TRCC[9G3FMFT37<.EQSg?ZDf:[KD@ED>R1<8[K^/
&f0)UA9/a3F<e7S)a85UC3@^3+b/X-A+MUM+<-ZW6Xb><+TB8MY(+CFf:]6J?#81
F5R9>R64/#61KMT5QXgHc@g;>[-IWb,37C]<RHZ]C1@a55:UUHQ)P;C-#C.LM2fE
\Ig;Q.Cb^.G3dd5+FHWC3Z5N8cMBYZX+<4/E3.=^f@X9EY2c\&2^(V8/[7.f\YE#
&-#L:2;gfNS^MK4@0\/@U/.9_[YdQEH6QP,HT,HMNc>OT;4Y#)e?^D&2=;ZGeIN#
<c.-QOT/fCA>a>eY6J2eOB=:Ed,IWAaY,5-;_0-X<<KII/HF0\N6\/?KIf/Ue-Tb
aCWCb;#KefA+X^bd>YK&E=PXTbX\aHH.ST]PFUXPeGUYZ/[f/EZ8_W5RL;1df8G=
\M3LGU-3DdZcRXEf0(H:P[,)<_]8YLXZ2fM^E>R770UPe62cG&OU?V(_Ia(:f,VJ
[[?&fR-Y>P]FKPIA9-;^7M&X6W-6L.C(:b\RfT:>Mga=WJW8@@Ud@fH.\UI42P#G
:EAM63O(T7E]R3E<b,ZF=,O)XK3e/^S@AN=Z,OX@VRE_@(a1)g_SXACV]=<bB(ad
J2Rd])daR6R(>SM^_J<&UO#N>1g/FW)?5Z&c#8IM8VbDdK^QEB>2aQUOU2aa&.8<
?)Q<:Od3bOceXeQ?)LDSW-\/9:#c@M?OeM8(=DT0efJ:.A]@)=TLLGMdW+1GU.b2
Ce_T@bXX]P6O-2[I7O)^\VF6YEZ9=Vb2b5d(-^6V6Y=0VZ&W1AA0S,BEG,5Xe]/V
OdL(2B\]&Q:U_:5<?LFCd,eG@e_4KA#fO(c1A<0+5=a[@dU1E/C4#gU\7fHD:Y4Q
d,BJD0&2KZ6TC?O.MQDX@U:ZCDYYOJO/;H+0C.e1JW)1=V,fD\PCQc.?=V;T^B>(
Z#+QV6fgFO.M?/2gNP:AQa^Z^E4JZaSS^[98dfaM2fc=J5BNC4^2,GU>CZ/d=/_a
NTFF4328=:]A.ZH@7FZK6BH??4-Z#T:[OA\IfGdZ5U&RL5[c?IP<8CNe^5FROY0V
OU98-dG.bdfV3;B2EFg#G+6/A699D7e>cKX6L-\5RFN0]VL=_U.RMI6M\JU[RDK=
;4.H:XM_0RU5\XAf_99KdIW0g]]?Y=TB&:g7/V9]TG<.Ad@+H3^f[c[TP11b45U6
Z&[LV\G5OgE)GO:d.6UgVO(>R-9:L#C];a0)+Dc<&-6Nd9PJ#gJ?(3@b6>A:V3FU
?bHaD2#0]OG//A:Q>IMGN3_;&#YDC-35,-8W+CL)YAPdXf@HIXNcUd\GaSDWLL(/
YgY<\60(EY8O)f>P&fC=2<EFc5MT<M9<gg,.(bOXd12APNPW+bJ9D->K60]Y8UUU
53DSV2\4G1YTO?f#XHXYE0<KG&4Db7NLM]W)TWIQ2L6DR1[aRM,#>HFg-[XMgIQ&
fC21SS6cMR&]<^,KN#_KN:RP0<?=3MPZCU9c/@d#QM)STNS1O@GJc6X5C<YDD6bF
>VG6ZF1<P&PQ1=>0UdMc-Z]AU_)L)##WXbL.-;5N73][9,U<F/NP#Tc_We1UV:/]
XFAO51);[[YLRLP#XeJaIeg_4Pcc5BV77HZ-S0WACK]_dV^d.&ZD.bBH/fJb[C+7
a;46:&(HCDb5@>/N?WgZ68eGFO=]8E-I6=&,DbV--Z3:7U3&;SSGJ<#JeD@NR><]
41ZYbO5L1Ie5BL:.7RL441^_G>3T^SRA[S[OfZ8^.+?B5:bL7b-@84>?+:_<>M=P
/(+H0N:Od5fTGV\dTLQ_aFJTcMM]-WIJg>@f<:6g?56\]8<8H8A)cV6NYd^;C&SX
e[[&AIbNd::D^+a@7AcL]\dO1?VX[GV0[e_bIID;\eT/g+T^;_0e[f^\Q8L+1(-X
7\JSfS<7JNBO<C]TC&:;4V-VPgb?B]1,KB9gA85_LYM>,_d2Z?V,BL8c/U&0)&P\
Vf#Z=\OWEGYY_-ef-S;?H<KYJaW=11(PTe;T_Z/>WHSN>P>4OC5;A;BgQeE(F96+
0dU.#?O\6GgNg1>6;9_BU3bLUQQ+?/\9]F74cA.6;#.RR;eX,J6SRD)R+cRMB[U.
Ef_;8<&OIMc.WWHNF?BUUSNPC5X]<\(H,M6/2L\b>X(5KZW,T+G1R#);X>42O20O
+=E_eG1b<HA<Tbf-[?eZge;?OX,Z5=<]eMRK^e+^[/G81WDgEgP:YcVG,;--cDdK
d][:W7T,YBN@]f4ER+PU.15V^9;RWHP\F]@:#4&g9@?+fbK7R73L;GeXXI1_OG\/
I4M,\AfI<KF4&FY?F.Pe>Z;O-]0MJ2+(W]7C#[4.V)5I(D6:GY&-_4D162KP@SBK
UbE&J]3F>Z#cS4PO3FOKU@&,/]Qe3:CG/+B\7_2eeIH_)EEd.3QY.V<8,C\S/&gd
(<f\N<NB1[GU5cZ7E^c2S;Rb8W#I7=fa,GU0?:Z,ZL;3)92BA^BX>;V=fG(bPf-B
-8<ERO-].#<d\J@@<=+^\BRR9f+R=JEWS:-:5dg\T]Y:A-\-]O.&-+(<,O/:@;>S
4KO=.P2f&]Q^P5L?R6CBCE54.I]INe;4J-ALBdEf>=CVZ1NcBLJg)Z_MB/G[#<c[
2BZ@VHTJ2WE,c3-b6(f02?aNg0N@>Y4,W0FI[<ff19^=f:RNC1A/c;&YAeOP;C<I
[4>X0T,.g^7055M/.](W.ZD7^4F.J2SVM=6ZA7PCRRQ+\-e1QcMRgWLRNfXF3J].
a3H=(\MCD4[4/a[5JOZ=-^RLOA2Y=b<([,25Ug6/0:NT+#<CIB)E)2O,HK&CE[O)
C3O;RE+.[0F3fcZ=Y_b=>H;=#]MOe#(\(<CBR#)&\[:I;I9)Z5c,DCfa1(+<Yc>H
:5UbMRGJ2YB<^_JCP67CA1_KYa2P:VE@\c>#9a#[PY>b[)J+HbY]\W42EUVPA8UG
7>-F8TN.FACXESe8[KIAU2ISO.MB+Y<&EAOKFb/R2_.K[UFEW,6O/RfU-1bOUWHd
VW26Tg5Q5/+>@@J#fQP77R)40]QWVVaJX5U8L,D^88da\VfHL8VW42,NG?DL/NaJ
X[\V-R7,,U3(3K&2<^0RRVI;<0?U<(&K+5M<70bO2@LW9#JbAAFJ=M=M[D95L,+U
2NJL_]35_aE:4(WCSFYff2FG\OSARA>ULaO=ed(Y_^O8e[dOC(6_T_=@S^GJ<cQ.
Ad.,4X_6SW:Q:GM\H:DRD_<UMeO<K-g:BLa26>R\X2b=^:eb:29aSFM,33g]gU.X
XOC-]\fM=Cg)1DfLEa0&fPB@G:?bUgY_bZE\WOIF/IbfN06K7_DDU4)(IPJP(/Ia
DO7M22>R<#ATX-0D&PNV#0L[7I,N&5[0K\EVV6324,dGI,cH)@,:\0:>D,0=7>=O
6Y>R]K+GDN6d/](Y-I)HIP75(C9EN87deD:5R^BA4VLWG(G9_GMc8Z7_F??<R3B@
H#[=c42R:dA2D;U/^-e3;+5FGB0NN;?,PM2[G^KgKC8W+787X@4=6+6P(-Q<]UH+
N,HG5<6cd_S0+9E(bSG4HHAZX9Ue+9:Z,4_b/&N/\S0?VM0_(Xe2&\,+3f9(g@b#
YGN0O[.78WZKafAS87K>(I/E&@b[b^gWQ;8\:gf[BR\)[5689S]P)X1.GT@;cc0K
(.F&)Q2T=H];)7[?US:>BXb,H4VXb+XO8IH?THTd8PO3,E7EFGIJ<G1g7CXPeU3H
.K]fObGP+g8C_G\AgD;b<PVQDd74Bec55+]Y5C9T.;M=HS+NU#C+9XF\/cT+[S+a
/M_R#8=V1Jd^XU[R+)\XgB@ZH9/^e>9M.&fT1S<e8DWI@g:3)Q[<Hf5=/Y5dd3/#
#WLRIUXG9fO=M=1d;X;\RULeI,;ADfdDRd;TgCX,;UX=-Y14eW99KC-(\F0V>P-K
-ZD;LF##<#fe8?gZ.&Ve@Dab)@J93HIUbXgE.A/4?d?5<<+Z9@DPJ(ELTGf1fL7G
54Q1g\7-e1B6E&_.4a/SVV]=4b#&Kg5bAS@Vb5>G6\ZeU1gdCS&+FG7(CB<GPNG6
Y45S,FU:H=M+F9K7.7\L9.UgR+W;(>UOU;V#Ha]@62aA\dMWg->f7R,8_]<O9Q].
eGH4EV40TWW>Tc,fg7]d[2YG<aIEVN#O=QQ4Ta6eJD?d_&E>WL];QM5/9f)^#)I8
U)XZIB/9[#C//D32TBG;DL4FS;R9gXLUb:^b4W+9SUU1[QZONU\]+CE=<OJ3SS:\
OE&/IIS_RJc#ON/aFPN]&T#)Te])K[Oc\ZPRYHHM,f.J8/5O]:LA]UM\W?0H:PIg
JgHRT_G06A]IRYc1f[;Y#[OgbG,MU(LGd=d)FUYg2e2&?9#e&M8;)X6=[Cg[]_cb
4^VQLCE/FOP^GdQ9MZ5ac)\)H@2+b;\>DD:7FXP9OK4.I6YYX88N&NH=3NZ6V-[(
Y_/fIJC)2ZaA]G7J\PS0.g=L>O7]-E6ReD7MGC>P3WM6ZFGcXNT5Y?Q/4&C^?#\e
BZB)\F<@LB<=/(<NeE:M4A)26EWE-D<Q\^_5V\D#BKO^],Db[d?Y_dLR4J0/-,C/
][A_4KQ>1#;87bQ3_Q&(?+dId-W1K=TcL;+\Df4,]UG8beSHD\BJB6F,DgUH7f5+
/QHF5D1,?>F)OHV>V6BeHXdU:_Kff_3.>>4X]a4EVdCP+NQbR8PegO:07f4)HK5&
D#2b;15,X7eG):I/IbFW1dCX;^^_A?0V>(-Q(><+C/8/:eH@:_^L)1Z>E4W/LLeH
P#+4HAg_8C_@LPfXUP&@O+\a+/@Ha9Q40_&68KDcIN10Z0393[#TW0\;:9BMb,)5
2Of.8ceRY(a#<JgfVNQQ=&@.KPU=b_29-Ge7U^Y5@XRKQGW)L^7Y6AM(U#W]NFJ-
4<UAVOE=SFg#c-8_fUIKZ;Xb<J6@3K7#KBGT#S@Q9Ea\EEHTb9\XTI4c>G&A4GO0
^M=/afS598WAGCYTVLbgLfV-Y9T@/O>aH+B_I_\V\17baYBffWO5cM([/+QRS,UK
6E/Y;5^c\0?]e.ceVLVaR@HeR^EICb06:FOOM.c8;897c8.^,UJ1#6,5UUU]^^Zd
.ZY_f.HH8\VBgdQIJ<JP&U5OLW9CZA=^P29N_)=2MC>?cR@A1?d:/NDAdZIc5C;K
A.<&^fUTIY=8)(V26DDXB.)FY&H>(?)[DQd7:Pfg>\#BORX94Sa<aZNWHFL.R2&/
>K@]YfID@ST3H=RB,C@=6R<B\Q83J:(LYK7EJQ=Y#3c3[UET_dSSa@]dV2E)aF6c
?fEa69;Y#1dS-Y,)(bO#@?8KJ;F^J2T[fEeQROL07b8N,cCcdMT&X2Y9X_A22[dP
OD<BaLO1?7F;5O]GA:T>^)9#f_]>RaXG.](0,?37^Vf]B_>2QaAA[1S2+N<HV\2U
/JdV/=LXb.\9gD6;B]F]feCAe(7Z>)0X>&0Z7NBDNS[,b@M\B=6H8Kg,5GV=]@M_
?Y+5C>]KcaE.fP08]LT#G4\_52J3BO66TK87eV>]c6fBCbI^^5d?_N>2G._^TB@N
NggML#b+#HMgE6@bg1RXXZ/S9>MRdg=Ad1<H4^.d#^^\9+@#O)5L-7]_b3)T/fe-
C[/.QcX)=BSR>90HQZ760O4\IUM_N(>O6+BB4)#SV8a,ZOE/83@?MUaO\#JO1LfT
IF0-/0BYW5c=@[d3f2^(,JAN1?(1F;)I?FT^[cEDR3(KVNB6=f5TJ.18^)\K=2#]
:?I,E2,EGC32K2S2A4(E8LYUcHEYHI+5#;.J]b3,?#2Lgb6[W4NV=RT3)G3L)aWG
E3RI@9([^:WIY^BS@P5JNJQ;@M.bHS2F-96,FbC(cOY>\_dGZ-]DAC40WD71KU&+
/bQ&+FSC>K&#gJR[5,@RZZdgN6HFcc.fcCK?VLgEZL\0^3S;F/3,D8GEHRbF]-Qf
2C:XD[)@XUQ8U:Zg<E60E/)b)P:&C(DMMeOfe/;GaeYH]=@@7e_;&J82-abY-LF6
Sg,e)#IIWI(AWQa?CbM_XAD1A)&_L;aKN29GFYNHL_O);3H_)P0cLM[^Ag#:_+a-
)#a\PXFD\CJX;N__b&VAU6[VQ)JR\Yb0^+CYLef(GT[[c[#D=D>LH1Qd2.6.VF:3
SI4=D0&/>E^Z4)JP-NP<-a/V<)U[fL(b\?f08WOZ3[_a<QWAe9>.^MI5&]G&dR;;
8S-?SGHGY>BS#a]Hb-d?bW&aB:)00_3T^Xe8eaMa^G7^6B/X6E&F+/+8JIPVV+g,
&;M9NUc-CB6c)\,^S76&^D^Yc3?QFS?:fN,5ac9&BPULbGcefb-K0dfeHC/V@2bT
g3#B=U/N5FFN290WfGYU-9D0c^=0_&e9()U,1[ANHJdWM7bI@1g^FS8I[+f#4]R;
E8V7eH;b:#?e=2W:LNB&b:?J4<[@O5=Gd=.,/c0O#@5Z.YPWDfHFXS<_C;UZHY+U
VJS4aLBecR@_8:c,BVY2L8=cJGV:6U^Ob&>HR@4>ZXDA.4H2fZX5>[\(-,@\&W__
3I8_CNSPfVLaQP.80AL\G0\)S?I_KEL[#d<HYV>+a^ZAb3,SP>)J)5RRbKI[I8_&
4c6fZ6->V43EXEX=9eW>.>Y_6,<6@OYC0UT5YS9Qg,MJgW))CTLT&9UH1<cF(4:R
/cI+bVc6M5T^#AN1H>8WKM\0K._cYZ.1/WBMg8>V=:fgVQ^/E=#-GM(N_I.XEGS4
FCUb[_E=e]A(_e#X,G2HeYFbg2RD+=dMS3fLdg1+UKHaF&S4;8f[=5DWcHQJPT9M
ZFS&8I(Gd^8eN>6XCOH5+\LMRI1C;Lg\&Z42>N\J+NZ5[21P,a_/GS7I/M#KXfV:
-Q8P]2@#^]2]5SC@QWB71I9gC0B?CV:AQS5LJLG9SU#H<T]=Zf1=#EWSHgGE27Pe
1Z9LW8?]#G:PKf4X2e<G\KU2)9)NK<#aT\VXXe2:60;@R[MZ4c=PS7]=X(8L[\d.
^aE-d)/@GQW<4#a+3_I<]WLQSWTbXD\QPFCU()?(1MLWg?ONQC=(JM2,(.)L:@BD
UB2.?2)OF#gTU+9=QWXa)dRVMM@]R-9f&Y&U;T]^BfE4[IS-N0R_\\0D&223/(WC
XZ/[e8G6(d=(Q0_gDbN[DUWN.cWL\,CYD.OfFUW)DZe3b4052^64BREL/.PAN_;0
d\84<4E6.ZN-PZ;#<d4fSEKV^SQ@CcRUPM+8ELdfD<RaT4^bE#;7^@U<@ZR9XcfF
]6<@<Hf:Md/?AA#;2=,@dNG_L9_7MKb/;V?_:6c]FF5B=b;LV12/3I/HV+=\3eYd
H\dAdfN=:)S1U?KJ=KS4g4G3LM6=VL?Ta+0HaF6WUXVfM=[-dC,aJ@QHNFe<+2C-
:PBd\E(bDfLS4X<KgAdZROgddTMW697/JMC4TLDA+Ff]TZJM9Y+b=f=\;35#Q;93
<29+P[[7M_JIb8ZafJ<&V/YZ;4L^V0&U/^X.>;KG.]W(,?NE,ccV2c&.K(YQ:8UH
F?73GJ6MEQMNJ#E9I@4Re?T/,&OaXd+baQR7P6H[0F;d((Y+PfQ)G>GUP6FK5;b]
(,N7X(83DJ7)@,+geLWJ5CI]e>:RS?\/>-cU\+,8P3^&D_:cG;UJFVf0J9Bf^Q+J
gD<8C8PKDEgeOMHI)MgPgJ[DN>4.(ea>Ea,X<V0&E8\(.6N^J]M5IC=Fe6JHHG^\
W>R\2g8XTCbE0c(ZBbMAE@Y2YWLV/?C1;gFATT3(F.5H]8RQ2Y[1LO;dDWZ./\P2
4SD?Z5I877V/)e9OOQ]6+9=NBGe(_)PMD:QBXL1)(/9,8-11e6_0M;aA,XJ0WQ6_
TU;),_@UP.0bSU6)?bYCf&?Q&<;7fc[2UdIcY=g4\1V#AG#<gQB9IfR?2W52_5]M
D)]??9R5180UgX.]+T=,LR(/5K]VXF[e^L9BK/:TTM,(A#W1#25SgRUE+PD&].a5
L8-ZMXV5K:?c/<YU)G-e[eT+H@.f:Pb3/fJKM&MWX.03P&bP_:OOc@)]/>QTW](O
MO6ZO[1ZW<9&TIg:,Z0Ae#Z<bGFFTZCg0e=M.-g4J68BF]/KTX+a(f:1T_4PP4MQ
b]g)XC](g)DU3#H1aA#X(-0V:1WWI_)f;e#1-BdFGc_YF\(SV?\SWUXV:FFBW/^L
K@&PCcHO[aA[JGc6bYPH,g=-CPJ@>Hf.dM@9f\FV,Q-K7-&CD_29E)QZ087I147C
8HWA9\fPf^Q;.B,W7D\GR9LCH<.2:1:4NP5g(0^/Y9>FCcTOAFeA8#3\g>.@VI>:
5T[PE<FNDK;AX,f,)D&#L?PW0a.3?C4gAQ&OF(VK@VR;N+-4@8(5U&UHA6eY.[BV
=>dA[A;4X)9.fE.WU+:1V[;TYHU[gP9OD&&R&M&cF(?0K55<\XdY/KU5(GVXfg1L
8T2DYNH;<c1BK+G_X+2?-3VdV6N0C2\]T/[U[fa)7;[F/T.7U7[Y,T7:T,0NJNIg
fV,9M.ZEL]D#XaE;N1V,Gb;3+W9>JH#]X1S/I>ZIA[Q0IFQS8H0dZZ/9.(ZDR17>
Ng]))abSFCHC=FaD,cB:g6KDc;[3#VeZTGP:QPPQPb\[NX^Jg^7_<.2Xab<WfPB7
^+D(MZaD\@CY/<&O&?N^e0KXC27J7]+cP_^)I-A107c?>+1SE29Mc8[#[+&58OVW
>LaQXbRJIO(c=Q-Z>]HJS1-6Y_F=O?W?D9I.d5RPQ\OUaCA;T6<6(9+b9L&.QZ1-
&&GVE8)D02GH]>CFf.VO.Jd9g;-_4+--dbNTcg/]b5\LDF[>aeEJBb@d\O4;XK(M
)]a=GM:B2g=;.R\RCGKKVVWPa7QB9RP.(VS\a&dR^\T^b^]#B&SYa0P5[?gR.O8J
UT6RU2Y3&BMFTR=1_T:ILB0W(ed(2ICdA>=B8Ygb0HQ\?)(_5/HGA^#cd>C5HC]M
[&M8+9UK0XfY>PY&@YE:Gc2-DDaO8I&JD<@N9O7RCGE)J@&d=]YLQHY<8)gOIIa]
_#^.Q#?7:P>ZS#b[4M3W\ODLR=L3?C4);gT0)Ug<K98de9aJBZ:^=KRDTIAVA[)4
VCK]87&6CY@EQAYRH:2S(<NFS7=>L:M6bO/EV^V(,HWNaDK4RXaad?ENR:aX-1DO
Q5\9c]GM(,</PW=Y:<f6bB&W8-P6<UGJT]G[ZD=R1^fELOE<4JCe3[00Lf&/Mbf@
HK0b&9C3=9EBF^M8=+/Z+0I3_/Y4UTH026O^A@5;I5,(E1KJfL>Q]FM-Pd9_:b+A
NfFZMDLA^:/P=M&IR2SSM3A.&BTJUbH.0^<=,U7D_Y[T.^],XXfHa8dM>?afLM;+
fPOQaAHTd<X<7T[^G)8K)35.&-K4EPOf]aZ&RF2&UFCHOP3d)Q>=_YPUf6-eI5g/
-;30?&5A\WB:_0R[O#)=F=EU[b7/K;D_G_U8I94QLb8D>IbaUD,DVP5.Ag1g5_/)
aL.Xe03@52dX-GLeK11+@#3<)?#];JbHA@^?-1D9Q1^LcGB,8^^1ASO(cXL6dAKP
1T<YO]<Q8WTcF:_&.[BX2Fb:cYAb7)0=X42OR);I\BH,eaVUE5PZd_BO>[LL=RRZ
B1;=eTF1/_HJ:[g:MK3(_T)bg5F1@agFf9a@IWZ1OS967).EMNMUS,IIFY0d/+4)
]GSb+WJ8P(9-T3W8,f^V@<[-&@fSFYM?66^LT+.O?SKV[TaG=2.(MS@(H?VT(REY
RS;TfQ9\X-2fDHS+#cOV2FX18RB[2[P1]aV<BU.L-F)bB(E2-:JKQ]b^OTKN\J#]
BL2VR.P==_?3cWeJ-GPea:NJ/XdBS08W<]6cL^B+217\)b:b:/DL[AS5//Y+:QFB
IA/0982Wdb@da[/I<NZ(7S.D[g?-:HE<S7dO6I)CEe4AF9UYE7IAY,c9Tg#KLNM&
UAS4P6S+MVS74@^dYb5G3GBFB&O&IJ9;&1H?NRG&ZH7SR0MTM+T_0=0@7b7_<I02
@@:Ke1NF&H,[=O@/f<WP0K1(c/NCWSFf>#;e6QIGW;cJ#;5SPJI@W-<MdBFF18[G
Wd>10cDGB6>NAB<&Y=]g,_QZXOb2@.1Da^SDLb>FU_#_DYZYaJO?LOdJ)N?6LVTF
K-GV&K(FH:Q>2\+TPMCT@3&Nf27H]SZCW+OSE8_5,YL]>FDRTG1_)4S_L_+Z#<7:
Q0TXeP[Ub=SBdea9/D<LYGf7#Z7U1eG&F+.N:+F;#L;M_Y4Xb4:?FTK,3J#cIJ3L
1^Q\KJBb1DI-2.^,0.2L_E@-eKFI7E(.>,BXIFRPS9e@JET6Ce2\=[AC75M>A(\D
8^NEc-)[>[?KC1;9Y-VOK-eQA2+R3YfU.C[W[fLONMPOG-MLeH(^,&B=N,=[b#62
@MHK]QC4#<bD68P.EE+@D1+e5JUdB)R&^\T6SPVfc5^PG2LI_Ta;88=X9^Y4(>H&
:==3X5WBb6@KZW/&EL=GE91GWWCGaa+&V[/[#0NQC9\S4?A#3OK.C>f^Y+/[KbEU
JE<M/MVV]H(LTW0[X70C)@]K2dGGb\O:=20JCE35MBY#U5?-W-&>VHV02=Y1P_aL
<C5R]NZKU.D_\PD\_5R0eSGN.YMcXH2JTQA@U072&eEIO@+aSL52I1((fc:7f^6/
-1-V8e4YV/(ZW./Gf0X4RdC(4fQPCKQe+3@c7YgZB4/4V+=R@7GIIZ7^Y/R,308#
=e\T_5HGg7A)Ad:O1,9O@1b3W0e[(C(f[d2&UP>TQHB#agI8;N@4#dUQ7-^JI(IJ
5XS.abB,>IcD0&ANZc_]>[.RG_:XURA8E&b&9IdPKa)H78g;FOf-^d>=[Z1#:2ZJ
.P[VZUJP=GS#g[C^?2,R:A@WUHQ]_c/S1Ae.a;1PY_Eb_\\@BB<34d<N)KS/WTV;
N(MJ4GPE0N][6fWZKI5ZJ1VT\9Q8QTIV,:CRfKS#)0S.R4/E53NA\cHc,TFd5Q?0
MQU&1)f=MddX>d?T]4bdf<6N(a&5fBRX@G2A/dUY6:]SUd>^Z7FZ^AbU#2f+M#P8
R_g5X86J(a]R7U:A+D;3c2OB[)+IDQW)f3Q)B\7bK\-G+]a^LPRcfYTUXZcNX6E+
[L,PgFNUW.g7gN@aVf+CZ]7YbZX\^@6C2;OKAf7e5]U\R-MgY9W&M?W9.<C2UX4<
gJB/T6J,\5+2M:M:?I>MDYSdef9X-FA2Y..5M:\Yg<F1[A<&7)aM-aI<FP(G^1)U
OG0@,D2ZJBfS6>01D;)YIEO:M#^TV(H.BbG_G+M/(WH+7?>SS^-:V>^,2T(,F#;0
3^:ReY;T]SaEPRB\5@H99ef47N7W7W@e60:_5[EZ(PYD=7_QV]#,:M<c#1VR@L9c
A/S84E+5)8QUWZ6acUQ/;3HT0IE_CLMRW3M]U(P+9gZ@egE_5F/+_Q#aU(NTZd5d
=d>MZ\KXWGf@0DRObcEeW3P&S;,.2+a[.LMeU0@SCT#TLga.RB_daS2/L6Og8V=/
aR9T[QIV^JALGJEF4MEE\@@&U6?)^\Q@6L?>#6W>c6^(Q3RRAYWT9B/\/&RHC1Ab
A#e[[L;A.Y#D=A@Uf6^@B->VaCL<2K^#]6EKcIU&>:@G)E9>-8:IP@47DXF^MHfE
IM,4P(JaNL4F<8@>_:==^T9AG(3(BWQ5:U-fB#PVd<aY>V?PH6C<P?Q&K;N6U88C
=6Q3HHS(SM4=+IePH)4TSP)[0g=?HF17]9N6]Og0<,NENE0d5McOIfQF(gPE?A<)
(@bb+RcW>WP&?dTS_0[)=[5H50^6::EgK,V_/L[0AH[edcfM9XT?eQJd=&<WJ-d@
g7f?-S7M/S1G-0cQP2ZD^2#QcJTA@O;E,5GZ-XdfT7fM07Q0-fg>CT9S^VI2g:aG
Be0d:;]([=cUZ=0/f04/U,EJ?g[GH:dJ>F[[?I^>,=4be-?@3M2#&T(bb=K)[2gF
YQ\dHf68)\SA^](/>(f+43B2CQaO,/CRN\7,?]aR2LF)#E&-]^U:4T7WW9C)JJ+S
4.YT]ZbRJd=1,9VIJH<<<A03=_/L28KX=YS_>d:C<>#(;/5Xd^L?RHXRacS8V11<
>D:@&[O2G/F51N@2RG]4+;\IA@C[7R\7U2-gMNHIbefAY;(<06gDJ=JA+b9)LBQC
#INU5&09\<(KYR#.Ea&:Q5dQBM5POB\]8V@83?_-9f1(fL1@/:V=IROF/dV6)\+X
-,V8PfC[TJLP^V9361X?.#VI^_9ZES:4\fOfZ&)<SVS50EP.eLc]7HP[A9WNg;0O
-MO+,U9JG+DZUTAH5Q=<;f(U<c^TB/S;2Q4N-c]DP?1,WNF9VF:9GPD:\4M[Oc&L
21MA_d>T/Y#2V)BWd)bRCF^^88]3#E,X//:>bQR32EV6,ZDR_GX9/T2=e6Y5IJ:_
.RI(IM]Q=<(_:=4<VA4B5bKIIg&Z.P#EHO\Ff_PIb4dL>=;(YZ?_Q;6^G6:BgFe(
+dV2EX5NfcQ>TJ;\g?_M?SQIW,a[M+11bR/+I(ES?F69..NQ[?A0>]GPI=WNPR<)
H4gd]IPR+W&T<;[(3aLS-[SBJb])#MJ2C@H6E-O.I82(]aMK6eRR)+[J]^.C\(^^
8_SXRHFaB,QO,2?#L_X^>#)Sd7-A]8.CCX=G:a,ZNeM+0Q4C-IPcV]Dbf+XCOP><
^-;73VIC8U0H[GNK]5(ZID#7Og5E/I#T4O:XHPb--cY][0B)EU3Y@^O/9Ked1QLM
#1fQb>aG5c-dX0&ULR7R7&^U-1>S]@;F9V3EY(E5\8)#cFgD<2FC:EN874DR=3/B
@YaZ&3?dZ9CQ3OKK@d7H,I6N0[a;]+,DPDU\;>\55Tf2EUY-UP(4[E9V<PF;6RS1
dcG/U3-HdE_G\#A#CPD3>eGD.YVg0<;>[8?6Z234aU6b;=4Z)@/[-RRCeUfP=A82
N.P\9f0ICd:\WeV&SH9M?MO-=21WGG#WJN/C>@S=M=df@:Ic&7TDeW>#eK<7?;e\
/M(Q^eT2f/X6D&#GFKa2:>OBM>0.@S?@Kc_6EU@/:_)cTR3;;,;Z/,PZb_4W+1OY
ef[#&I89ZZBf4S@OL-6.4e]bdSG&CX0T\U6,5(/SGJS.Ycb5KOgd)ONVT=@]Pg5Y
N1F_KMF[b3OFfI8;.6^VEO;GQUEAGK=R.:ac@M,SATgaKWXZPfe)G@LPT1+&I?HV
b)\UgQK6#0O\IAG2=F#aG,.PfS:XG:NgMaQ.b<Z7C;7dCaI^+@+<Ub5GYV,L>WZ,
@-MOX;>&XgF:H;T3G-.WEZ4SQSU1MV52#C@X#g3WE\A-=?_&>Aa:P.8VH[@P6@c\
F+LW)gR8TU]M2A8<_>N#(P>f/^RAAScKB=)eB#g/4LgTG:B&:c/b<:ERI&P,D23[
Ia?]L#EF=aI;YH5eACXc#+-WCgW^Xd@I^508g_Nd>L)D<,[KW+E&:O+@I^)RBgA(
RW(d:dHABN6:V/EU6+,_NX]+Kc9G4d2XZ8fdca=,M28bX]1gX@=Mdg]&QYTT:eSG
U:/]#<O?2g_FWfBe85??&H](N-T.(AAQ<&L^D>L(f0bXHHO>E^9Ke@+ALaG/bFZM
[\L+D8A@<>I1TZ5d<=H2N#<cbW/FHN:<1.MI/G,B4A1CF+D.D&5ETZ2\#3/ZB\L?
I+;V0A[W7dHWZIFK7J>I#6IWWTSKZOWLDGf^B.2ATGf>&L-JZR0g1=G55?O9]#ge
c9LJ0\?(>+4bZ/(A]Id<+6H:a,b5ACeCMHO^N4_XgRJU-]C7?K1244VI0[?BLV]L
efY8)_);,-F_G>SC?9QT+5SQMQ4FN,AW(-d&c[RQ8Cg;&&A0?A:Z>_2\XVZF9-a_
+J/XS&8[CZD8=C?CCZ)Q<G#^Q4^RD#0&]3,L#4DHZ;K?EWBWB.X/COUL)@cb5CSW
G8M(^bcG9L-UE]#[EK/Eg=VQ\aL=++?[8=B60I,T1NWAXU=d#N[5bf0EFd4QP;)e
/4TUdGS;.UBDce.3:\ZeX.=:?;J+B,#-)H=&6W6,5;baPU-V8)WY713VUMX4?WC9
V:,S2-PYT>BZ;_\UQ)_+\eWN?,X9?,_I4^M6K/2:0E5VY(Y[UJDa=A8L0Z8-I@31
2Y.-4IC57ICgX>@cB0LdN;152JG&RNG.L88@\dg_E8QH[:2FGMB@](c&dE=Y(SbP
CgE22fIffO<ICNPX2.S\#P;BHO==GH3\=I)UZcgN4R3c75?AC?^2#(&[T+4>E?@6
BX/+L.c#NK:B;=(#Fd^LL3/8IA0,U+).<97(LH?VR4]J81)ZG.f#Aa>W#X-e-f7&
Qa;::(.CMS;E;LYdAaCAOKBS<U<D+#]W6/0D=WMXG-O_aZ@<aS:B&1Vf\&eHQLIA
gE7+75&\aa8FXVe?4=F7N46I__:E;L=,XY\,ZK5eXX[EW)[4LX]IC&c2dQ\e?=H^
ZE,gE?\ZMY8Y8cKQ/7GP6&:<J3>U8U,WLH4a;;U+0H=I2Ta7M-.DQc=cN[K-\WD<
OO7D)b5__(MI;Z+^\Jaa==[\II,bKgKe8+;)F@W/eOI15XMSREb4(._JY&WFKb9_
;Gc&)Y67#-MG6N@N)^850Q0ZdK[EM2gW.c+R#@UeP<+1aP_G(/(1P\Ya7B+MCEb1
E)Y67-;.URTBLKQdA3ZU/^bXTReb\OY33]9A7;d\TM-VZ-,15e8,:<;=9]2OQf;?
ONIEd.4=:GUJ@QU;#.(47EIQUaK.P6?g=]JVcGaf&A=&K06=2/>Qd-K>:g#U)B#>
S]U.?5_MffaEVWe9-9Y5d;Af=#a)]0FS/LaTKW2D38)S6D2F^_H&_33\OC_FZEMf
LJ3Y]cKGK41Z00=@#NH/EFKKW76&U33D#B-(T_8?(Ad.L)R\F8MU1V5AOY(T6F+c
TM]JWP8Z&J4KZaLI>#R=\,CF:/VA1<D9,G\2R3GVNd3b4-[BRO@5706cdTUN?,Bd
baZ^45VT[_?=-R+)L4XEI<MYBA1QB<)IT^AE2+]3R3@8)\LO(?)G3bN1)IX\A1=_
,4a7APUa5+?SZa(9YXd\g62+K&e1TLfI6=9>-[P<W\=G,Q>bf<JI+=P_gaWV\F?>
:?7)]\KA1@8AdTfV&GJV#AFE@H?6:b#Y/9RQOX^g3MRZb(cN.H->@EeU0SX(#^cc
5)#>0J0O9LPabQ6C]]<aV&?e+X7.RA]Lf>S8_c_4b4aT->4,.V46+XAb/^dEZ6N#
@a[K5Z2<U_1IP31Db\KC><.56;8DPfHf\,W7#K0+/6cQ^V(VF.P;4OQ#6H=,X[E-
-\9,N7e^@(QE[XZIbZB<HPP=)+/7Kc=Y2Je3H>CBSIScaUaGHC0;XB=W6H@f.<d9
8B^)M[0M7MZQ_G;(L:S+SQY2<VZL]1dN+[<VN&-I07e/)Q77V:H9A7[]4756#[U[
_=?,,KG(aYJ6/]a6(TPI4FQ(C)1cN2R:U>7DIR,6#C=A3UECETDK^7ZN2??@K;B3
dHRb,X,8QGF<.QV\6]:X3L;edc5dJ9G_Z^I0&e_Mb9gNSC>63-T]:,61THCd.<[5
51\eG;1b>8YYI-\FI#^CPe0^GBVB(Z-,0LG3QET4H^2#C8GYHf@78g##4.RK,TV1
=be7SY[;#D&\/_YPbXYM;D=TBag\B=5e9TP)X=,TC1N<7bQHMMJRFOa=NBB)f2OK
D+6-T?W[&QT[=)<KH:H7HN1^\Xa=EU7QIW:d=:?)c^GPEd[;<)-S]_3]([J0.WPI
g#<N3MMB>+.[gI8?\R-6@7HKQ0@>\2C2ZCP034=eN22XcT\CZ/eEIF89]GSUaJc0
bE@CZU1fKCHfI2VWc2.3H=JRR7GJ?AA\]\Y.>G+4UUTCPTMUSP[CL@G:(?.=F7NI
Y;53aT3aU-A04=S-]>QL5@)Y,abQ[7CT);@8Je.HAdaE+G(RQ]7Lg44BP74&cHP=
:BU#H9?)G:I<WAa2+D7XG&XD)3W./=WIQfd-7^)OP#73f=N\A.)g:d,/2]72SD@^
G4U_7AfS=Y.A7:-C5+ZW5PFS92KZCMT[;c6>TRX^gBML7?+#;\B0X@Y?+fc7_6,1
E:=0.Ja?0Z01;Z?X1c\[#3a<4YCOLEYXGRX4R>&(3C>5Xdf>MJ-[BXC&aZ&^76JH
)[A)(A]Y#_c1O:g=,W\Z?RKVG6XWW]LW.-FFJIBG5=-@,EcX0(4/7BE9?7]7b8gC
.>W8SRQR1O3gJ9,?#M^B26S#J=-VC+>@&Q;I+MF6g7SFaMd#IC:6_BGbPE,Y^HW7
eM?N.TDEE=)IafF+8>>M?;b:IFcb#Wa2Ab2)bI)2S53GQN?<?DOYdZa7IgVC@2NM
gY:7,D=#<8=4g,P<_0SMVe(^CefH_KeGfK:8YONTI@+^)?N4\G4+2(dVLC6QSYbU
496+b#AEd/^D4CQ)9,]]=A(3VCA.\X^67U:#fUa\,D9DW\R.1b(_YbN^LKMU3g86
d)C>g[?8GOdL5=V5GJe-U-1&B??2Z&EE^O:2@O7TZ]e7.AFAf2UA7bfMP0gEecg6
CN1E-W\T<[&6]GM&d+HH]]5gY[HB=a)]D+dF_gO=6]\M(,_Vb?OBN1R8,\X:e(Xg
VG_>6OZ9Xc^1f^(f1H12ff&JUSVGA=QH0,G#&@EW5+gOB\bA/C+33f((UM(4<QMQ
T3P3RZ_30L+-IG725;;^=Dc4T5D66bOY(9EN0e10&6f-1DW?0<5bMQ<5CJ=C#RI9
<X[-Og\[K,M&B@(-/P4F^=N=BG5>:BAfH.J>?gR4Q],Y@HIVbYUFVc?U9P,4A?B;
&Z>ObOd=0DXC@YT^1&T/D8&021NE3^AY@M@-XU9-:eHL,=I#\?C_U<^;/6<Lc.cF
,0_\QdeS]@.,6KCe)6\@-0MG)Y7)<.X#=2S(2#+Q[IM?cB>0QL^1>&1/G7VIO,2K
/c,M6YEIWe.LTaT@Z3X,K,4BL17/[EbGKZ[[1PZ;WF-I[5Zf^b\PeSYL+42?bL.C
&0<4]89+UIf<6#H-HP/d7d5T=J;[CU,45@Q>C3:R][.bC,6J/DA\WF1\:WHMC:e1
8Y89EZGKWM)T8(8P+YSGE@9c</d[3gP&,K:VJJ9&7AH8[S&XL,4Y^50KC,K1@+:,
+/.YX.HaK7.W6G91Z;Oe9<&aAW=<[G3Bb^LF@>(P6+=a=a(fdL)>^2.WFISYZ=4M
T46?-82bE,TeLeIA_[<Y-9WK9#1aLdb:1?;-e[LVZ6OLW3O9-8(1\PZc:D/H0[HR
_7:SA6V5DU^>K=-=IT7PN(C,)5H=73Q_LM.+^9-B[J(^f>1=9(U.+]KD<X86S>69
:4-8[1&@g:[DN#N&-gSHT+C1,-/BZ#;6YQ]9>EgB&(6L9e8SL/Z.F6DN^?cWa\U@
J/3IAaYFS4OV&_2MZR0VF<A7VOZca-THG9Y5=YL9f5W?=(O<3(3U0A)3Ag3F]b[;
MJB2.&1f[3E>WK[6K0I955I)b#JDTMPNVIXOYI)J=0C=@ZN7-L.Ga45Y_3ASX(MF
_50Y)A,HI:/<E>-W413<f\ORWF.#P7&fAb[O)?=8+Z.]OZYaA99B+O#FI.3ND.A<
<f&HbGXg2d15=&CCM.6B]^U<)Af1fSNYKIFBdQ032KdPPS,1V@/fB.C)<FIFJg?0
abDA(f9>D#OaHK9GR]3B1K->AK#<PP_2-ET>.g-<Y\H:IN?gBT:1V)UIaY2S_@@X
?#+CWd:Nc?)7LIZ@#SQ&Z.dHa[\4S7.8IB?I04+gR^De:e=[X;d0Yb0PIO7_?YK1
?G0W-A>(-\B\QZ=3-[-,].I;Ge6B:V;Q\.1<Y3f&WGURE?TW@#>QDE_F)>NXUD=H
,K::N,?=S<06e(GKL,;AC,AeA+I/?^d[&:?;L0HQ;^5aR_P=.8326OBM,e[gL;b2
+fdDCR8.a2>_)FP&X,9+ff?T>96T,?CW/-=FeM);A^e7f^NCH#@6W/L#EYX5D[Jb
T-XGbWW97DVaGae7^=2A_L2(B[YU[M?(NfPSA.(KN,#+[]Q@g2KINTM(+L,5EPHY
>1)_7LN/;^8EH741@cBgI8AaNNVQcGU9F7WP(MF_TSC0GDQ:@a3T+@O/D+SN>eXM
04M)2AgB890HYX;(e&E9Yc1Xdc3d\(6AfO?.9._@/YB<7(OJ7,,46Z0)]R8g5N]M
==:SS:M+W7PS>@=Q/.f]Pc79@;3TLG^F.]Xb,0-.4gJIfQ#bGIe39W.H^D6/,D4/
K,HBO,b>aTZ.;_S00;P>T\RIdg@7G=>FRM&dfJ=c+,63c1J[+Y]b6aYHb#LYDXc5
4fZE@9?ZN\GOC-&1I>G(93dV3JRYe6C?X<Vg#AHg1TdQOg#D>K[FeLf;V5<<.6B7
P,GH8T7[]?+LfcL\^V)Z]f0SfH1H[-?ZX;VKA\b59K1G(9L/:DH#=?FKH=2+&RF5
GBB.7VaEAFRdeH?cUNU8L\T&gB?;/^CI+fRJN/)d_\0OUVQ1<W7=2Q85B^#]1=UO
O&ce;6W9#J8V3_SHL?=O>GF9M^RAf(=G+L3Ja/7#eccWF0dK9e.QAGFJW8+;<8F&
L]0KG#Z:?A]\0[.0)>T^;<3CWfL4=5<V_e-^?9=f0_c7@>;^9SOOZJRZA;-[,@>@
d>_1?K\C?PV-,WTGb\544R/6(D79T<@bM>MRRE4f(>H[V8)b_38QKZb2]S23]P7J
,Q7\:N:-T,.XNS7LbO[;,#5S[0XGHd]FgTK/a+;g)g8I8.O>IM)-0_1Zg#0L_[SG
a+FN-HC3G,H7fJVd/RGL^8L#MPQ.bb_S_9:V_8.@e^E2V;ZC9f9/L<6E;0C>ca[:
_<=PHF;=UC?a1F+0(5D9R0M^;KdCJSZ^OH69N..M^d;9VMDQE1U54<PP[1K9;7[4
]YTPV0=>1I:GP=M\@Cf2IM.<4PTCH;XcUa-]VWY31@T_=g/\Nd/dSF5E[G->-_6b
K&[:>8:L&S&@1B#PGb#1,?VaU[ISPR@1LIF6LdAR<\Zb:7Q5H>AOe1QYQC;2A_+G
\WF7-c=_=?&-<B73P10@J?96OD\>]^S:aR(P3&TK^ZY[Y\d0CSA:R8O1Og1,5W9=
3T-NNB=_X^KFO74L.gV@MIE3fS:9/90bE[ON7[(;W?b0PbA#LMS.&KK=S;,g)4V[
>S[SS9ZUC0?T2C;^3Z(^a@SABYJUgU><B\\_VRD:B-cU<4)dJ3YBB:?6,)J^9Y_;
fL.0+UVT)^e&6C1]KJ3W<6GbK<F.2bFNZDXZ&JHF_QB&W#U;Q@R7C<8BE:5+41M9
K75YWN,L7.^;+G<6e4AVLY[cg6&fXZQZ3Ca1(PNH1XY-I/eD9gSbMWa]<+b>E:T0
O=&QeFO#Y)Y-f<=+[@MG:=,d<1dHVb:B(;-G_AVX>ZKKJ4,\UI@G,Ba1T>W063D4
76\T6,5Q4bV;;<JAE<20;fSI3;2YOYI7D4>OQ=,NT+FPZ?c3:B1=cK=GbX/gS@_B
Ge=Fb.N4K&<b:55-#O-X6OL8Q^d@S6Nfb&C0D\1A^F<\?IK45Sf5K..^]ZQ-U?cK
;3\/)#JSX^6F:RbO.efSJ^H>[2SEF9R>JU_,dP.aY^9T4YSD=O>^/Jg=^O@Y.Ng8
WbQE>\NLY;&,HVO?=ZXC<DZ0-K;VJBWV^-/@+S[baJ4fSKG548:V@7cC7LT0MIa-
_TKf0ZL9;^Y0T)ELGQ@];S/C[5c=O>(0U)XEX?87>:)a7KT8fJ:0V:B+A,_5Y:D4
c7.dLZM2Cg>-&2_VMe.V2IV05[8@aW;KT,a820PFDLN&V7GY=@N_(0,/-8QN#;2Y
6QdPCB5[#.7TCZeTV]?eJ>0aPTgJ5K+F-C/)605IW,ee[,IW\F-,J;5_/aR-B4aB
YIB.aIR<U^^f9IDCNVZBK:#.Ba.XMZYU#TD42UP8X>+I4H?JY8cJX)gN;F?0:gcC
Pe5#A;f&?NfYUH-&AEc._1D/X=97R7I)70Q2Y[EdW/N>VX[c1&\VA;VL3Z3H^e[\
VbW@[)XbD8L<\_@(7G7EObH>]ZV[3PLL.K1TM^U=HE@M=B:Y2>SBFQ:D;(VO+e50
PVGQ:V?1G+Q_DE=VbYD>gc#___g(@NMfb+b9e_/3dL.1N4AY<(HUB^BAd0aQ91E3
f,GAd(7W2M:FgWD+S5f:FbKW)J0=R675PD#=K>)PV@H2G^TT1BFBU1LZ/NJ6f:<a
:2U>,8FU>Q\EB)A)233YBN#G7d?fC@)NHOU0[&cb#8OKAK)78e??^T(Q79IF10Kg
Z5OM)TLc.4cXE2Nb2[I+1UZa91TNa3#\#QFTSJ/,R2(+WVT&0&1C&c@CbTgXc;7M
d\DN=@(Z]ALD-[FRcRf<KaY2RgQQ#[?b-Be50&6.(YaIR]@Y@GS1TT&R5,4@(g7M
B<d?/HfPg#AYBd_EZJR+aS-c)gOMLNb5_R7/KE5f)A-&A)=C8@@f>A;E-GR?33\a
3G.@^fB#[b1+K_&L5M4Re7U.Oab#(=KQUFK24_bAU[3,/<2-L[X5>UVG-ACRZ_[g
\4TXL.;4MceLW+_IIFQd2R_3)JXTI+G:03fg2Ff,SLE=f&Q)GK4eN]>W49Bgc<M[
3@Z50X(.LAQQ[:>gOVE\=b+gTK2X9&6g7M_CHD]FX4=I<CISObAO)OL=fJFXI[^+
?f?NTK<9@f5A?^9f9F1;c6<^FTXe=N#S>b.QdL[ZcSBQ1DY.OJIP^CeOH;_2(V3O
W48NB0:A1-4YE04<F;8V>Z9(&@NLfT?4701TY7Z)4-=<U:JA)&(6XZ#BS<ZH6,@(
&O/7e@d).+,Q55Z50T;CVU5L);5>6g>,aCY-&cK),AZRfgD;,@f/c[:c7F\EI/Ue
V<;F@PZ&:;6E:5S\_N]/-;,Xd_K6(BKNYUD9bNUb)d3L_P4T9@C->()@eMZB)+;=
<D1fgJ\OR5<G>3O)4<POE;2CRF\^NgT2[0I0O2\Y?Xb<2;eCbaN1d,NW9OX1?fA+
Z[]fC-abd=&/DLDM)Ma-IP(@[K5f^L2AJ^eDJ,3(3EW9NC7HA(H6:,X5XXOCOO+.
/PP0>gA(g[+RdA]eKGHfCC_+2LH+P63AQcB/H^-@V2C6a.3<CLF=C48CUcF#?/^5
9@UJV/FSPDPW@W#,-gJ(=Fa\[Icg<<(;&O-9Q^f.;K4&5FgC6F9[>+G(48#\fHN[
[@<?F2?)O953B=^;YFWP0,EW0A]AR+&?U.976feSdYM](1^PMY]2C:]G,K-93@-Z
5TK8635A\0(4Nf+XQ=7&WJK]Q-[2^2;Q[UB9X(Y^\@P;.5:.Pb<2#6/6DV<[;01A
&gJB\cIc=6GJD9U].f_VV#B,JL\AH]&ILQF3QVYT<TKNB-^3F&70#5OP6a;D,H=^
)/e)W@1N502_)=7#Hg1LTR6XSHRe.<:]7T@23J;3^51[M.(W?7YEb@\/NWASU:[C
Fa8QXDWFT>=E(?705eGUX0G2F-WO(80Vf\6:7&@G&/.eF9>>K;YV/KL29]a?&C&J
()eC9L5NF#G)ZeK4+5DP,N]TfaAK1=P^]9J./7/<e//K[R?I/VO069^cLg@,B-R0
dEXeL[\.AL_NWH9cP_/F?ZRF4>.1=F?RXW_<=BI].1?L+YKC?HE&Qe87[a,eL@+b
d]_8C[_XR>,(]>JXB\?,,UcWMX0-CI^3/BX;+/)T5)#N8beSWJ=F;YFg;>0NX0b6
aC<MIS-R;0P&/7[CF3Dfa9eNS4HOLF<Dea1LaRHcZ4T;\)CYNM?A5[R/6;e8gDaR
;f,XG;a7OBa>R79EVS\DWA:cg>?X4W(]YGad_[F\UKP/P,eN--g)(PgSf8BKGFTG
K5NK\LTE83e<Z#.=L;b/8Z6EP.-I9@K7+/@M\=U,;&LafK1c/<(a9:XF))YIaDO<
a+<FXSK(<\5&/=COUEP[NB40\50b[ab>@WZ_L,d]EL6f4M.A.P8=eLU//L=7AB25
Z;WcV[VU<FQ&9?T>b-L-V7UC)-;,(gR]f:)L\J57.+-?\ZBPLXZS-_I_/CQ^--\6
Y/K)#RfE(N_2ITDDU/MR7SM=?DW+Jf1QIG,<0;YeD&DdB8Xa:FP0<-,\-b.Vb]Za
YF&XO^VN^.Ge<.a8\fJbWO2K.MW0FN>#>4+=A>V^3Y65NV>3R#GD,T0-2&;6.Z&L
[[c;,-?4@ag26\fDHJHH##ID[3_KI1P/T8[Q/[P0<N8+E)#FDB,f=/:=PVC<Z?LZ
-@CYUZSZHBY/&-39cFY\eXUaGCHG2_Hcc,[a]5?U.c/fd3(YL-5R2GgVNb:N,QE9
2@\cRgdg[D=0GESGD]2SR>G7WGL^>=T>RSVb(egS,TO17JgC<=R;J,3\J#H0J^<+
-ZbGd??e>)EcabLLb+LWF2[:@cOZJDX/g_Z1aF/c+&PDXSN69C#G>[LXZX-W3EUe
>@5P(QZ#=7dd9#MZ+CE#HDVc+BC07L)AaP<6Z:X_;#-V,e=Mf0>I#X7aFN1G@eK/
WP400NNWTgeL1d0P&H.RS(F>Q?[2/H@7Zeg_F:_adV6<,=X[#Q;POCXVP2gEg5P9
3Ob<>;,LE7E=RaJY#ZHOKRP;Y,X>Jd2b?aAFHMTJTUf/M1:&Y2UVfN72)Ab5DW8#
J2/IB73#]d[X#>U)W.D/+@_RQe72FNURW]GcV@&P/)?+gd2YSYbe&>-W7Y6J>+>e
]S[(f)/;HfN9T:L,WHLPObWD7ZN5dD@M_GDI]=4cc.UO:C=H/B#M204Y^@=XQG^I
eE:fHSPf@_RD6a1-179/YNE0&URZUQ<^DRX(_^cMR(9)=cNg+LG[L2ALA,[\)Mb6
aWU@G7=DgPTN5Ieec(XBF8P<FO]d[[HR)QQ@c>4SIbD;,N/G^G,dd78^3c+RCDBB
-85B/]\7:L_>\GOA&QC<GV+O5RI@OfCXgb-6-E8<6dH>^V[9K1VMH18^:^Rb&6ZJ
KA0C83<ZA;fN<ec0+:CICD;faWL6C[#VV&/8:F\KKS0(>M-6D9_1C-:a.PPW>L24
&:BM]AV#Yf:7]WF)3SZ3X=E0<Ce9e4;YHJH.H,)0T2L+#H:ZB07/<&0\J3END.Q+
>5g:@8>4HHK:dcI2/Z0=.CPMB[F>EC05(W9M\DJ74BgdXPMY[gH6fU1a)&YfTVIW
KK73(N]>_YUJP(D04<Y1F:aT&&^MC;TCFT[OW^Z#?d:XS,/GAc.4J.@6@24gTAHg
+C&aN?@S5J98];e@Y0df=L;XA9[;2X:^G5O:@Rc>721b?CbL=eUTXP.4YbC]THR<
C7d6HO62:9#WL<F=R9/63WM;#U1[(_C;/6<NCP8a^3(Q7H=KB0Q1eP5c/)1@c45S
0PgPCP89J>/f_)^@@ABU(I=?gL\Y0e<fKAI.0YDAF=.=(WIB)cb<^dd&R@aB=D,H
R^?UZQZ6,=XZUdbCYG3NTVCWc[EI/fV&5Y+-GdSg&7H4T1^W[g#Y2.OGQX^Rd0K[
(dUK=fFK(8B;14ZE]^5-.bJ?RQ^fR)90VMI[^4J4M&KO^2e>[)fZ#_I)W_E^^?a4
^+F=337QC6f,-U,2&]9BD9_XU>/Z#ZN:(CX@L)1YI<K-/2(FRWYAE>aW-J[-C9ZR
//YgA6bPZbD/]bd>9b[ae)cNAXD;5b@=F[7]X7bF,UOeMZLe_7b7UgY[LM92,HPA
&F&bb.F#SU;__H\ae\;0Me,SA>\X8R2-KKEG9KN>F_f?@QLOHSAeYb_CX#ZAV>d&
UbUXb)8L?__.W018DQWZ2U3W2A+]/\IJB1V\JA3++M_aYFG90G^;OP/H<Rec@-Qc
.<)J5+5e6#;e-8AJ,\@LZPDHbABK;U-FD)]g98ZOc6R/(dD,@RP3R+@bW)bb-XL,
dbILA6R/:8-^S_-cE-.ODC]<aIUHV=1FC\Y5S<4[7bO=#TUO>.3@R5<b\LbOdU0g
Q?3f[)N&5-YS6F\<La7.VQc>5]Bf?_SXKb?TOC3Ed\L31J6b3N(5S+;>gD]+85B8
]P@7T34FPJ781,>GdFXQ@UJ[_K?C9VPfD:C0f_^W@?P<A:T?KVbSIc;b;VcVL-.g
//cN2L_cJ3<M2=8R5aC@K7Ma0@L@1D;[]P:1/\BX/-K(fG#Hd/\MGFFW2g<ZH=,;
-QC^L3JBH0(<,Oa<U)DQ4FIEQ]8_Vf465R^94<3_a:5@65(Re=5YL291J7L<KBLA
eZe9TQT=Y^O=/Hc(Z:3(RQZZg=Dg]\e<VM3Le/WZVUZK2+&6PVgfbMM4;)1:L4.M
R^]M=L,f6_cW]URJT9a3;;^=LLM;4FQ8IHK>Cd/cT)8L.>AA@768gXM4a3VH+<XV
ZdJCBLeGH[Z7eeUS-]ZBaZV2eFcPFO2H<GOCE;Z#HKc2;Oe\fY,Q-^6bSKg-F?O7
L4GA:-)\;PF=E&06]?N4F=Dg6^VUK35bLe0)b_b25<O1(HU--5\78RfU__TRe/\/
+QDSU27H?+A]I-CfBC-L6,f)9#V?SE.DDJ0f:J-d;Z,gG^=;VDA.-[])2DVC.2aI
]X8&3f-#>VFWeKE;@F3Da:48[C#LO7ccRR/GP+cV7NI8@_OURFH3Qcfa#IR30\Cg
V2UU#eA0#+L90[\Hb5]g.?=6E?8N+c@_PA:U)WI9;_;6\VPc(UQ8H[^EN11ALOgS
\AV?+--KV75(eA4NOG+R]7U7@4D]:P&E<GOV;CY?UaG&RH-e/4G0JM/Q6>X=JUg+
K_M((E6d)()bHK1DX3-XNWNb=K^PN:D^T>([^W/7c86TD5Z69OdJAXKR7a.S<bZI
dP1Z.0+H@IDX\5L(H]I#<P^5Q-E6X,NI+fS:;B09>C^E62E0LgDAX+2V&ceg71=#
K=e:#WFgD&(P0R(:)fLVCD?]&14K<M[Y40(J5)B^@;N[6Y\AS=K0PTa0UYVC\C+I
>P2C:6MaG0g2H^-E-/X_37=RI)3.W8d(,>GE#V05dU.XTE^=]TfCVVCZW._LZP_^
O&g;4Ke<8M&WHF36H]2eKXBdf7_HT9-]D:XT\F1fX;(E9d>g&f_7c,6&AG>8+_ZV
c7IC^N<Q-aKc56B/YNU94N:?MEO52<NR3L_/@BKNHD/Q1VIc9;Gf4DH6SOM^F\+;
+LHPV(C4D3T<.C[;4;,#c1<2P?,BcU^US=:BN9T)IZ6MYWf&8:/5M>Z2^]c35AD\
[,MX7>UEUbaA_E6,B26W)PHGZL^0=OYIc,35Q9a@LN2+<[Ge@_RV/53RIeGYBN](
LJXOc2E7HaELYIc\]d)<-Od@7#N0\eTEa:VU(3.K019RCEMTb2>:?7#?F]]#9QC0
B1[8E_X/&KY57K@eOXOHCTIaA8D7;&7G3]SZc19D;S;G/]?WEH/CaE28=;OW?6/)
^]8bE\[M&YE[O8]eQg]I]RD&7.IK0+KT(9/Y)b7^#8(2YgbM2=SR[S:4O((02f[e
<b9E-8LPX9aNOUP74U1c7e?(A\0_32M:M(#1L?fP/GNa7dD,C-O7WKPgbK]T6.+0
.)6?HP1[IC5fJ\]K&3W^_N_TD5EO.C>fUf<47<4^8(KF5CDb@=QC_UTVbSE?:^T3
25d7RQMA5\]C_7^UgCV2e]Kd+24AY:<FD&(,B#SN/0.OF_46)2UX=^Pe4+RgH(^^
M8Y_QZRP;gg8=\gO\Q(@Y;2)F=9LVL/eU?8?[,?eZ-I-I)>6.QIK125TVE=/A-KH
2US6-56@I8JgO[aO3V,3WOOK16F?R--Y=#6=\Q,3SFSH)Q2ZSW+]<gW^+#bgT;@8
&?[DIU)-5Q_8VR8U4EPC),(Ac7/XJJ@+8^V>>&J3eSUITe.798^,eT_8S-U52)U:
XZd9PZ\<MgP7f00H,cHcS2\3BR0<:=Hg0[]UKP/(]c\TU7eL,?BX7)PP8]PPg,JY
9_\Wg9S2QYBd)GgL3Od<Je2>>UPX\b[g5(X.Ed11J]G76TRPB?LIZ_8bC5K[K[d>
>^ES50GV<FXRE9M3e>?^dH615<[,Tb+b6a<D5G6H091[I>ZJ6Y1;cA?9X91M<c#G
N01/CGRM@K6Nf^@d_P9f:/+gb&gZ.#U:AKcWX&/H7WN(F;A/E,1APEN;=@2Dc<RQ
#Y./.7XPI.9?/E[16\-M@gX4g4UBJgbSC;;9?.1G-D&_YQe\A6[NDD:PWT)7=4F?
JdPG5+NA(W3bGF7STV7S4@AZTRNJNeXAgfIAQg(0(dD>U,Z;Y(CgFRN:EZ-2]-6I
GV)7cga@UV\@D,,7Cc0<QLQSB(]IPfGR\5:22)eCWE-A=#6NL>+8RgX_I]d8Ea&=
d)Y(Y),Y&Q]-gKUPb\cT-.b[<+(K,dgE<:)S6ETaH<>^eQ=/4<1gJT-PYb7(]cXP
5U/JUeJgAR7-MXec[3]OaQaE41X#9ZV[=,RNZ-QT)DCgb3CUXQK&F7Q67a.SRe8c
\JDN&KC(NeZ,,JMdeVU;08E84]5P2O7>BU@J56<WTLNF.-W10F+;YBB5U9b.bb+Q
=H]8Qe#7I0MJ#+_UNF[_=Ea0KE:1cbDG>12F)W7]/7>3G/^?0&Z6F?8NgS#,gE6N
J8?[/.\e0&--fD&,_5X?BJBOB]3@^[8YB+TQP]&.LW&[FFgg.CMN(df=FFUKG26L
:+dE:H8RV2,YNRW?A2b^f?NfD72S8#10WcSB5M]f>GU38B@g80A\41(2d,g/UQ9_
F<1+OgFVH5_6WZ>2#QE<EY)U_N@TUbLC(#Y#23<e8;7C-T=]aQ)4O3EHe5Z1-9dA
&B7gJA2L)BX)2P(1_A<^L+=]W,aS+8-K/OQW0fJ<&_8PZH44C(C&CXcO1)R[C&4S
IA1\O4V:?-d#B1bT5b1970,1L[CJ\<-Y;B06A(RV?Z)2+&-U8R_\CNAD;^Df6(=H
)7_S#B^_>L=6#(CC\QM5P\+JK,0AX7MU6CaX_=@;MK+L<bAFNYK#][ggdA?P:PRe
<6cbP[WU7;]W5:b&VcQ4012e;2f-H+@B\1UIQ-b4=TYSJ?5KYC+8YXZH(:7[BfOM
>[?H?6c@e,WR#>?3edQX;B6PEP2RF9RKT<)[,J9F>4Y>TL^g5_71c()B[-B\6\Z@
H700)dOP2A>6IY#H^bZQKR@2#UD?(B+g=ZPA?VXbFKW_Pb4HK]-X1Z0:=4VL=2UA
S(c^;@(PA<BOD41;Q6GENGGd59L7Z4&UR_^d0U,W?VG-2PR7;ccO(6^&56\6VWQ0
=)>]<G?+U_=RO7a;=MT^Q+U^[5>#A1:PP\^^TYWWL]V[#.W,K1Q]f&A63+7g8>aI
#<2SJD_<H^@N7Z[Q5Vd_cd.Md/f7/@C3OeD+(;O[+TBLO^cZM4W##<J;3L1(0J9;
5BBKO=?HRN9L_+/=N_6H1(1,=9U3aaSJeW(1ATVR\^E#SC[X?^,G]8DGC0_Oc(<Y
ZSWe=?a10bGFP\.+9&\5A+R6BOUNfZ)Z>V=.3Y[bTYVHbVKKUY^>9Of-(-6FSI9/
XYT_aQCI.YC22gCR/V=@I+SS-CeffD+#H-,P.EPOeW2+3OCaM=6?0/0>_]4&Z_Ge
fM#=CR]BS]][(eCBG_T)d,2cG64g.-e^V=5]d;0gb@B[O?4ZUOR>DB=XKIO?&c]F
X5Wa=dMO&A:H\]_\E9.YGQaBCF>9[fX]Z=]430_:\9,<G;,72P9:OSB#T(aaK;L6
5YJ8&?P?2+DWSH_IBF?E)<@E99c>fFRDYd.9-[dX2B2JLR3M#ALF2YQSe0Wfc8+(
2P=,KbcHUAH=bN2G]@_b:;^VEg3D9NPZM+51,55Z[:654e))#DCGFPJAO#[fB]V>
BLVF@]L4B>9J;.Ccg8IKB;7H@9bK=:JI9Hb66\PJZa[:Da)fCcF_P&]+7gg=.S_4
2+66c+/XF7R4g8[\@([22#H2EbQQ(_5>,U6aBEQdKO0bY114:D\:[^@MT<a.dB2M
)XV#Hbd-cI-c6/-\&DD2>@4^0+O&-dJSRTJP.J4BZQJ#(WT4c77/QdcAZ6#3O)H_
G=@O)L]J..7f_FCEOTde2_6GC[(eebO+BSAX_Hg6c8X+C_8fG?ESASdX(@,H=,7f
E-O.^Ec[-g?9fV@XCT1TR;QS&V59-&I]..#:3E_;J8[f(2GNcO]>U[4gQe^G)g7=
9KfL<cJ;>_8@<E1F;1a(M3W@2U>J3Ja[9X;Xd^QE<.,,54UFec@-U61V]D;,ID6+
+5=>)NfLd\::PP63Bb/=12:,/L>c89WFY<1-[5gL+N2^@^TYO\d(>B,eCFT,N/.e
R?_eaE\0Ff(c/F8RI,0XBF3SK&B,a(MT3?IZ5JB)>K(cR2TFK4ES:^aITIeHSR>4
f->,#U-KKZW2OAN<XXT\.7TgS=fdNEVTAIWIJST2&BTET,]S]59;eQ3EQA50cK&E
V;JQ?@:Mb[/7YE<WEdQ](DLe\E&MG:E^-2O-;VXaR\dZb=O=L=CAd=6]3cU5)JOI
d^1?XD_^4/I)43/R=ZBD<@_G?:)]87ZQM&BYDLb=g9-2D=7PN/,PK)QP4GQ\:AU>
-OfU5Z2E4Q1@5W-R-^+I)M?:)4JHJD&NB:cH9QBR_g#/;A-(N2a=Ncd45HZ4@<^C
TD5)0IG1=XV&Z,1:7)JKKP])5egS/Ycc^IU\A<?>ZFMUc\g7]3C1Ja<T8X4A6P[g
>)S:8ZC4QPcN=eQYX.N3O-3R36V#A:9(dWaCaD4C[LDR.cF\^;Xa<XK^E.cReA-1
R?G@LEbIWP3)gD-+;AAG38If^JVd=@<g)E8KD6_K=IBP(B_PI(aXF]S=EfS3KCPZ
.K4)EUO266VW;-8DC0;3c<5d&>edXg+b@BH<@#.F.^VC;c/=969S5E(YWdU#1[Y0
XVD/,+D7?<)eZ(BbPA?gSP#d3_D-R+-X&3_R20>f.La<(_cJ.9.RU,<WZ@Q;KT?K
N[@cP/,AYP3eJR;?(/TU=UHIcS9T0&GO9J@TU.EC;G-fRR6+a][:UZI)=B/N>OQ@
[ac>\FZF+1MG]RGNR(,&A;(UX\=(9CfaQ>4,g4H-NJf3g4SXTVU2UTH2&0L)4b;M
d_U]R&?dM3GVA7H0\+N_T-(bO,ZK^#L-L9J&XF^/81WXL[a7fGWG0JR_(M1T<HCO
e,&8T/5WAXYO4g2&WN_18:9E)55[Z1KT>X^PP#+\:Q6UCO_E2d8E8[USK21=d5Md
MILKN]@6R91[1-##.NI?=13CUYX4-;,b7TVR37.bLJPdR;RIB\3]34,[B&OR,WYN
8:[^4dXK[g32]F5R6^T>NGR[IR,;b=;W=U[TYU:NQQ2RRD\)A(HE&S-92J6.f2LW
4e=Yd73-b[G/7OJ,.+cAg\QK@ZCJA[XDR,N+./RSbFC)<g_gPe8]c-,Z20e6_65P
Gb#.6WL[\_39@QPGd,J&EQ-.(a1GBRGWA9KCO8Na?:Y0?[O?E=62I\7;V-LWHEA6
Z(,Hf[HdM5E0Q/aKR<XeU?^Q#HIe#a=Y\;dM)9;fQ,&R#4L8(bI<;D#SeIU_1(;#
24-RJA\4],b+)XP\.ESdD\B9=[7U>I8Af0IJ2;EgF)MX9YZE@bYdR1Q2T./&4<PV
5\O.GE]Ua(K]TK94I8K6&.f=__4SOb5K/NWZ?D,&d(MA]L^=gWAHQ\T@^;Y60/+Y
R5Q2f40?AKb])LZDc/&JS.-;E(6)GU,R&5RZ5L_SAX65/N1FC,MXF).H7Nd^=.eU
;U9.R&N(Z\:RgcEB3(:R4,/FDGV[ZQ5N^QMa7MQU&4YT;V1H-OZ3>9[#Af^feRI5
=f8-bCg?4=-84EO>G7#K,M>E(e^(K,0LA+\T1#C@fB2<6,J-L/aS=+fY6_W-<@ZO
?S8A@7<:CEZONSE-V_^^[+Z/SCR../?QR>I74f)GE990>IXX>TcgO0,JL?T^HDXc
5dEX^[9?F]TNYg.XTYO6eP>TZU>S2V.LcCJ?7N7=6UD>C^_6Q1[J(KA[]L\UCIF[
1>ZA;S.:2].L;?:ZQL^CK-a@/T^64d,a2/@-HFU+HVGOVgC#W5Pgg2;WRO@@7=cS
W=d0-?T]<ULWaSaY-ZMGXEbe8B_O1)(-bbGdD9-)GLPS><@\@4/fF#:]XZ6.BCY>
=aBK?_M^<YLe-<b(K#_#VYf35+D#]HQf6?eeJB::VeCDYA2RQRWbID124N?:7B)6
,:)4+5N4@J1\02.HD6VJCJgQ3(\g1F#\:K//eHTO?.g]Lf1Dg&3NNKRS,7A:@deY
9cQ<)g)3;XV_@gfGD]2[P^,.AC>HW.fa.Pf3d(I8E8IZ&c3I=Md\HYf/R@9_6-TC
W>HLIW;Fg2>/TXF1.(G0LcNLf-b,^;LceOAA@9NJI=_YB:JfSOLS]9-RJ\Y):9c3
-5g[8NGN6_GZ>;:V.)V92X794Q(9NRI_]0DC>-fDMNA,TM4A/Ua>W27&bBI6E2\A
<#C:8(gaMaMe(eef0FWgH]Iaa)^ZZ4Nb_#cF?e1O.gWVOb]&M8SZ),&LM8aRO>J>
Ca=TGV.&2-Z]&bddYTXgbX,da6K5:YK(9,1P,7LaOFg5+F6E/&MT>KLUeX>F[.8R
DcGH(bT4DX9\f&@WN58>\GZW0H\?/E[_QX8g3#_U55@d<DNUFW8J1\a^8L;4<,,\
[dbH2S@Q8DMCDB57(/c^]/I+F<R>T97/+\R/T9a31UT@70,bWCSR&I7-4C6C.)g,
LC&/^C4C(5-X48BWcY):)g>\=bC[DK?_#f2D#3_AY/=,@7S;26\#XNbZe[\ABKW@
DQXB]7c04K+)NL[?A#-Hc)JG)E0KDbA;I14U0MKP2,D>^L.T#T7B@J5E-8EbS-V;
1P<eC5d1SV:)9]bS591d\(dWb809Xdd#+YI@GVASF\MZ_;DL<(8=R;LT9[]BNZD:
a@[H(/1/;\&3NB9de_]X.f(A/P4L8=245dG#TcCWRJ<V\M_N#(EZX\OZ\O\K<W09
QI(_bRM^(W,HU?:0,8cE^14W(<\#Hf^G_3631-,<d=cE4@LV1#6FXHS3Q.++&e+O
CMa3]\&HI:#HE(Ka0)Wg-MY/RbZ.61dWT.gfE(CJ2dR/)HGESOcaLYFZ^&Q]A51W
/UP?LB<0//5<X58\]HG36DgRMG=FQTQaUMRSKOV[RcJaIW<FZDcdYB-0>HYe,IHG
2T]BQ2f0;OIT387Y^Z_IAYMAKW=AJ+MZ7H5NOMbE_^+aGaF8YX/(U7:11AC]S1L7
#6X.;D/#Q8K44E53/<@9U/^:a1B:XMLd>+,Vf+Q;Z]3Q?+;@W;eE6\,@9YNg0>W=
QVgY;JU+9P\USRE/VM8B&+0b@?#:b2J.d<BY5+3UUG1IUF1f]^9/;?]/#NL)DY<2
.J5OQ_MDd7=NPR4,gDZH^Q@[UKb^I[@=c7.A<S9eLG.9/^8?&./3gDH8@Z]Z.HfY
J[F=d0IcDJ)/4@\F=(U8Kb2Saf(5/gN5C/0c,0H5VJ](1<LAA@K,9eE4L?C<M5GF
bg:WI7g7G#g7W&2\?6+I&HQ-U.&9O\Z-.Sg[B@+D^+(V1A0M-R_\AT]KH^UH@:DA
APMIF]SOBW)&(+P/B;)LVZ4L7R)]>RX5dD+]E?)Y&a:=XIQ&ZV&Me6DRJG,.:9OH
d]LTX+V,DD@:bEIb4eGbHTbC6W81-<H;-?Re7dHa\^3RB[e6(S<b6QJ.MRA(S([_
]e.]dUQ1DRd5B+KEQCHR?;OG\[G^TLYb3LXV-aV66<<CT7N7Kf^(^5RJcGI,KK_U
G:]eKI>T12AX[B_Y.H08PL\J/ZVUaY2W8\:eB(C;><MZ.H]B#=\Edd,_2SH3R;-g
1eXfTILWO5d^:K)H9DZ<9@a/^NPQSeRM&((BI;CF#2:::]-D7\KJCf_c;;&]H8(F
8#\2X(#S:bFAa1Nd&H4E/gOJCCQWR&A<d=(-e^/J7L_2>^Q7O@C]b_b_>87bfaK]
1#>/F+gdGWab6D0#e0Q(^.U-1P5]c498VL>ZbdW43<L.S\T-0]>&<(gXKLAUXOWa
C5EL::&YO;?LMFg]<(f7c^/bN\=N9.\LbT^#[SSOg;8[F1g,1]c^.^,](SU#-M6\
E,<09WFHR[-,,7CBe)c:GO,++_A281A]@836=4.\]ge7@^4_5>5:K^3R:-H9OF:f
RD6g:Fde.a;3:XH4;F>GVBJ9\N[;W87I=ac^AX_5?-/;#@.9<]GB)G3C:/EDg]^<
.AbIHQ+b]\E?CC<8DecF87PMJ7.,[;a)Z3O_a<3=X]+1-B_b1.Ac9MQ7]4aQ3Q;^
eMR=D1SDbPA^_N_ULf:SaP6VV>aWYJ6_<>^c,R+/g.NAeA)TJ./>Sf9SCF62ZF8]
d_(,?1P0FR]\-AMXLMTA^Of,)E(E4()\68D3H6YMEC,CGH1I\VTMWWdKa8,[,+5&
1.JEQ)cLJM(&B(+RKf0cW_@^K^DG.:GY/e?QHBVP5P5ZDDU&?F.8g?D(+/FP/^21
Z[IW)_cZ<V?4DB^LZ3ObJFYXEB(XaN[aGb8e(2N_)XYT4ZOYZ=PM#?SRe,c:LIdK
:\@f>6T].5KPR,7J6cSX+eJ2b::HQZV&OL(AI(/N_WPS0FCN4+E&][a6LK5Ag,G>
<>:^^PJIMY]:^;?L1)KE^6e:?^f/>MaTH^+C5=.Q;bF9S[6Tdb-GQO-fUFI;WV1>
Pbd]171#[H(4Q6=0+Xa=cO-V=@@0cDTfA3)0V\YO_@V+@U9@\K.-?0J;>ZATV)D<
S.P@_VYcR,D)=[gdaY5&E9;SC6E;H_]gCd6BD/:P;GU&gQd\dU.J^TNETG;SPR[-
6IcJ4+e#cdA2A^@DcHZ^W(?TF#PR1)NH&(HW9)4Ff;&gCJDP_[\076IXE5c7U)e0
&5b;X_80Y2V]JCQ16CRf\#=QH;NMJD&<eDP\=?a&_e=,?2:K.6Ga6_TMTDXLaI-N
8MFAH?RJg3BLd6N>;f#YER,Z_J<5@)5#+,1SeXZa>-^T>(QSU@+V9:P]Ff<Za[2P
^Sc,,XK-L9HB@Y(X9T1=XN=#&ed)Oc#=ccRMC-G??RD&1#K&fDQK?&UC.PB28&\b
1+[UP[X&bWY]Lb-NO#FKCY^>?Z6H1AJ_OARWgTWe?E@@Kg,+)YWRW93U-\M/BL^a
]2Y3-.&BNWQ^_O3P+O5,fXR(4f&Q3KSG\VP)RbIO#bIW071;UY.UgQGQO?M1MD1,
GRbI8eO3WN>Ag-SYQWB\]e\.;#7b+e^cbe)Rd;H(Y@YZHA[b6=NQN-9#WRV8\+Q#
0:0;?#g5IcRMC7PSc5&N9YaRQ&g\(7LV34KbY<:-&ZFE604C8(E1Uc[HZ0-9&df5
;aOYE/3N3)KOBJ\e&TeU]HKE)^@FV,.SN46#>>g_+2??eVX4?7JX167.?cAQW9;(
)MeT[e96gg&f)+L7>,.+88Z&H)R]SFM[:DN]LDbM0fM:&D)48SA#?@_cICfa4Q=#
(d7:Ya-I4e7>Q?YaHC7Ue&TV[eN7V>Wb4c:SP2_Rb&f))\HRJBSX,>XH8XeZPEID
B-LF\53T/1e@<PPH[a<aRIbQA>e2,_\PV,Ld8<[77D:SG1=_.QZefc0W3S#,Q.fD
Vb[,;\gDa[-3&PT<81D5_:8YgOB\5OQf5ML8?g?KI]>,8>S4<Cf_F]V;[PX.5XT,
]aKKgVOa_,QM=C@:@0I_g][/08P3KN02[6]f?3G8X>F[fTHJ=O<9dLM<>,H=I6<K
/ZANN43.BdF^eN-J>&&^D/cQ)TQ=.])/7_@b@Y>7M+FNI>5O>@>(KIRRf\caEQCO
^PGCF(Y<:H-bF[?(<;4NP(1?f7c;d@3,aLR@)UGCW@^U\3<KUH71=YL>D@<)10&R
Q\X;CcO]=#[(Q+><BR;/7dQN.LXI=@;IA7&GMOaIFH-6B0,(c..GI^R2/J^L4P&7
Og^F?:]gH0L1)1/)ReQA3=^,ZOV#0e2QW6#b4]<H9(JOe^;@T].&a]<@a<?Ub[:H
RP62CO:ABZJdDSgY]CY.NARA;CZRTb2DZ:D_7_C5IJ]\,JDKI<>L96@P^307AaeL
8BDdC&Ef9/W-VII+^.-3>L8^@#;SHgUaS9I8IOH397E(g+5X9O(03BN&J]cA]DD0
BAC8_D#E7=MFJ[<(Y5Q_]-#;=7<;#g=+M+Q,7E3?]7QF-g.;RA[@O)[cOR.2V-+Y
Y^?.A=@XeW>_H_5C_@R8AcUS40OMf&PY[>+[ULY?4@&:;P^EYW-)6=F^2\eX\L-f
TH-J^6@^W5ES-:J/7G+,e_NF(aDX?@GK9LG6(PMWSLa3YZ9CW:AaFdF5)/S5^d-R
Z1,=TNG.LVM;G>@f=F^#,K2/,=IRZBZRC^gUS)NO9Y_\gNA#c3JLefD#<51#gQ8c
=CU;=),4&:L/#(TO08E=8<PbZf1faUPE6Dc#VRR0]Q>dLHBA,/WCg3^@;L_.8/3?
2WN9+7800@K5Le3CKS/6V:2gd57CFS2b8,S&X#ALS6VFcN<0>>?Q;0Y>P[4?)Le5
dLYM+:aXCV=BSFUY]IANS23b[)TecRX;C/DJ27gd.g26ODFdZT.?8]e=1-LU94VL
,SRNC>?E.bXQL,N8N?\aMgeR10A;_AA/#23ET^fQg40UfEdg#[O&_:HH9A_JI56M
C^MVgcWWLX14H3Q\a+?((7V4SIF<60Q<62HNGP\][?d8]L6GgJY=V:N>g;9O7e]&
cZS>@EZbHJ_e54OF^2>H.e[&2?ZHHXD5Tbd/=\dEBF;]@.4-5cYEcT;.1eCD4V5#
R@@,Y4,G8W_-FT8V)=3P&_4QB6W0]WP46g@R#==_JM\Uee&2-@[BSJ#5]b#QOV/d
8:\6)/>2d?R4@DLHNf<<5+.]I4Q9^15;=BH-\JF=B3>&3RS/NKReMIYg:.@aS<eE
=H0(4@>WUK>DCY<7P0dQF2(O5:XbP4,H[-JJ@#4?;@SNb8FCC>^9bdF0Cc8<?;E(
WQM^HV85?];,X1<(\,?da5?=R#\8b+T=.]PZP=4(24SCM+L,F0((DKbLBKSO4-_6
5Gg#A[E&S5R;Z1D:]RC(S7DaK7\NF-:OTY/fSS\&e8+M4]-.Xg[J@W>1U.WL\@+[
WW(W\f#89SKf\.ZOY[KNg0&OP/HGRK?f:B[H?]JIHIcaM\JY]PWTM?/ILIMPb;.e
:=b>(Pe/GCI?0L75NB?fWQ.0Z5)f1=HF+1R]N5)>c:_SKf@[b4bSD6eYPGG-/QD@
E@f]1#GM.AV[ef6[XLc->HI<b0/gc3e6MG14]cWTK@4\cX#:<4:+1OI.,AU-;4IH
8R69X&^QdfH^8=@/K&(_J/O_BaWITC?GXR[SVE4<O]/YePVPD.H\T(NLGJ_?^9Ld
[Icd064-?OVQfb&)?-F,+D_YES-?R@P,+9GE#C:^KfT-aN1e?_&G09B2#f.M[UI(
[Cb3^#AfLg)OTR>((@P+:[f6D\P:S2ccG7XJB@7PX;4SA/6#1]WK75<d82c9fP4[
,NP/89ZTOAX9=@(G,Zd4OUa]a]NWH5,>[Z37>J@31&)[=-ZOM]eE0(Rg05D:Ce]^
;A#X-e4_.dC?EP_9@&dO:TS.HPBFA6Y8-+WWR0e_D]B4[F.^f9bU]WfIBb56\@Pg
fN,(deQ/C2W_/6@:W^UW2?:M<39.<<cN3[f5YTJ/#]a0VU;e57X\4RRZ5Y,/+;^0
S+^3J;c,V6e&[YD9GO>FSa\4e,LZB48d?e0Q4O>Q@@YX-bYdITe,TU8d2PZ>@>9:
]a[^)S#&We8#UP^N.GKC3TEYAaE(aW5ZC:DU2a9VC\_>T3b[Y&Q1NVK,[LH,3a,+
GXe1_YM0aNS+MSD>cfY^@I;e2X\]g0F923MR1Z0FO9.XBF4a(ReJMYf_eW#.?9[Z
O#CGY)Y:>M<-8,.IJBWYG+4AfL6\eBc1M.T:edVZJg=TWUJMfNTCfSI91U;W=Rc2
LaI[16WBY_2J3(Z=9^<9b;gGg3\[EdcY1E^L5Dg)WdX#=4.F:KcYUBccFIBE2T^N
>K7WY0-Z1#8#5+IPUYCX_5+VeKb&>,^OQd]0T>F4QP_)9N0cWRSA_1ZJeV.&+^K8
3,gLG+O[&7?e3-0Og-LHTDB/Y1TYSBfa-AH<P<2:D?Q/E/K?<Cb]_->/40P6;+D_
D:O,AcQ&ZMd>TOD&ac.;J_D2HER&QJU\ePB@M<<SB.DGES@Ze1[>MV8.YU\ZDT8S
YMQ);)dU<P/C?A8STT(D-Q?&;K(R7=7@Na(@7&W6D<ad1HQI?^I13B@&1[F\L3fM
<\Z>8@f1LJA^JZKSZ/X0S8-WD3+QU^NYKA1#Vg:ffW>6\&V:Z_,V7,(M?G7e:f#_
G+Q1S)N:C-g.;?J91@-<=Z>4.3e=AJ&Ne(dcJW.@>)Q/W15:ZgfC4I\R8^dH-eDK
OU7KCWc@bA>/\B02CgQ2:^HOE(2B-#-1_G:(fKgH&NLM.4Z4EOE+K&;M?cYH<#H.
BDUcS#L44[R(,1bRE&gcb4fagDF=c7_X,\eF_J0^@-+&cRXcUW:\8Ca-:YOQbP-S
1]d=YCeIQ-]R,@S_g7R4J?..EA,+G#(YOMA7@GW<5c.RAE5(B(N?g7-VSZ=S,47N
Z7S+;Z^cS[I0_BI,-S.A,]>/#,(dfFb0XPI=gWZS:>d^GUB0_RVV9U6?F]A>TYff
g]VFRRE^:5]U)UcL;WC@;ICb9b:dG0bBcRcQKZ798UB>,0DN=;JU9P>a(fWfQ=RX
F,CD@Aa(X@+S@,^eE@4IdJ=Y@-ac/PK?GJ,DQ6]8NN=QWXN[RC#Nbd;E-JZ;Q:\\
?g(X8ZQSV++,<&B+)HK+cAQ3TC,50339;JaSO)2cL[.:PSK&VQWZ3O?Ocf32gKGb
2EF2=\#)B=U_#2X3Q&-W/XaSXBaV>QV+>DG/VE32\FH8@JDg;@3RR^HaQ;GP^Lg?
O/O<QQ?DQR=R:NDP5cDP60ED#[7e26U0H[\TVBJV94Q+\Q3=A#eYJX./fA;(2[g[
@C(W^NLef]QSOe>Ld:8Tfb)[<Gb:6?OV:DDPf^YD,;D@C_TF\QJ[)N/7-=JF_;df
EY<K08bUV1Kd.MT3P7/>c.CS)8d7[7I3H<T4&4cAWJb[Gd=-3g.VI@\d#GWe=6A[
gA\W7)4_eVAG=PL>>,[\,6V1[6YFfb@=V5K#3F2QYg<L;Y(-2[&e?39e5[/&D5[Z
f9f&3>dKgE\RG4EP_<X\;FX]5Eg4Jg;RW>5@T5[)B9P_#Z=9V\SSQRRL_>3R8\>P
T_&,8IDLA<B\1ggAY)C_?GV];:6]g[b:QI3UeLC,BX83>&@6W##XK7KLaF5PIGYe
:NW5,>4.BJc+fD^K>ZQA,a3E?Gc.DSZK\_2_=NY\9.H@Aa<,T,R.TVa_(V&;SY5&
RI<:C]8D/c0NQ6BUP;?Y#S,OQFLaXcL5KOB3MF9BBGSK:YO\=g>SXE,P0-7GT6#1
(FVG[Gg7FYagH\e_.<0+&=?#V&#(ZA>PP[AG,SA(?0HJKY)6]TY<3_f<K:;/Q5=W
AgaOUc;gR0dO>6N4MP&f-D#ZPT:>9^DG/)e7gSHL31_/60]9<:)3b+;^[1T8+O54
5OT=A,b#c7#ULS#&SF>QW+7VP#_W2O-UPcO.bNIX#7]WVG2Aa8FNJ;7AZ)fUJ4Kb
A5R3>@MTU^?A//:Z?0.,<1e^EQ8WMW[=&017;=[EBS_[cNB_7VUSOB=1Z/P_&1>#
T#BZ2YH#?VM1@[/PG;^^7#420@=/[NZ+@N9YPT_I6fFAZIcb&Y2?N;PTY1HPg0D(
HeB30S#UI9G>7F6O2IOWg+>MaQe?Z5:X]13BgYF7Z4ZH:HZ\XcW6AJNJUgV[;A+A
\4+&]<0:.</5_\ZcRR/MG10RS=NN8SJM<;C624EIS0#VbY,\(>8f-+&/O/1Ce5O:
E&;=QX7aC8b-CTB\:HG(ZQ:2,#8B>1,<BbS?1#<Ta(/(BC7&0.f-b[B\ZeFM-CI2
?,d5B<LY^6@39fBaA=,W2<IC@]50[Oc#Ed1^f85JDT+K-@a=AXVc&eP952,DSWBK
U^E]8>H6;UN6E;HH[&>-406\S\:M7OYC\#X>9:<,:NUcW_XEC-PDO#a&_2RG\U@?
dCJ2RPbMFWW7>&6V=+1-91ITFFFXa/gJ3@#,\>P&TdA\,MQ(=3R],LZN.>:G&Qa9
_+<]g)cB^FF:E_9Y(7a.(.GFWQ_;b[PXb(ZUa:R97B+dcEM(&9<9TT^,T<1-V8UU
1?cOX94=R-YDZY=12\L_gDR@H]F;IBE9.MMC]NQ@]bMS+9<,DZ?_2.4UN4G@Z,RD
:^cd,G91HedS10,P1)8_O>f39UI8dF5,.6Z[D,a0E>:0Y6G[]EY,9DJ5R+6[1KM;
#F^f>5UeN8bJ(J)0]&5QIS2\OB70H)@OPeU+:Kd=gHVTTBE7f>O:L,?9,4_)(?Q2
-:O0^a@K(CS+HUSY(]4DL-#,I8-]BeP,/#7&dSYO[]]dC06G;2?SCY0J\E)&5>F,
f6;aAc&>\OC\O_+HP\)<(1FASa&I-T:GFSc-\JDG5(WfK8SH_.D^K+JIXJ9PH,(B
cSY]<T9(X0IC]B+HXK=M04B-088/.E(/GM6F/Kd3[b(:FGO<:fUA>Yg]fI;V;8LbS$
`endprotected

    `protected
J^^6E69fcH1X?E&2-F[\D[7,\gJTBP3-Z3]DdEJ)\2[U)0K+U3H;-)NfcD,Y]8^(
&dXc,/?TAR55M(d_U[Nfdf7,2$
`endprotected

    //vcs_vip_protect
    `protected
dd(>P&XC1&;I1G-,7G6,BHMf/O0/dJAU#H^X#9.NI9?NB)WTb?V@6(aJQ+@X>/_=
0Jf@=;>eS@c>Z[T,Od]NBERX?Q8+ISg:(>a?^?:J4^COKXK6I=]d2:XSNL=AQ9Q,
MM<g.]SI9DdP:@b8Ag4GU+3dA66N85>aS1W@eV<SB(g472DH(5Q8eTe.V8@IF1-M
.bY,JZcA\-VIeQC45ag;;EGB0Z8GWc6(VRV@IFG3Hd&,@-62>4?2BQ=G=,KV+.GC
D24JR@(9V1:WC=\eLGC_5K\#Z^;W[g:D\BKOX+]fU^SPDGgDFRL68LGV2YgWePA4
b.UG6dNb@._e-YPT8Q?[,)]BS&eXdY1F)Of]PD8AdB7=\@e[D<KLP0HJV[=I_)HB
<RS7(#?M.]DA.VO^&QT94>)^&=@JHALRcL^Lc+.?98dF1+HD))TRbR5F-dQHB(V\
a=0;P5\#F>OMQT]g0d;f.50#RS.#]4G2RZgQ5=4T?(/)^G.#XN)MHVY[#1=_fH]Z
F>C1,&e@X#)\)e_e5@TSUbBGG=beHf=IQCV895^Ca5EfF@)DKPE^@N-W@AAR=.R4
01+WS:WcC:FNHPb/WN/4g]P.GU<?_BfgEV[bU23Y5,dZJ214dI5\Jg[CQM^,S0J+
?(+2V0:A/cZ?EM[-79B^af^8=ERJSHCBBfLcX\<+TDR9XEcER5a7Q8FN7APZ;J9@
Y-1FVDY-U7_N&Kc4Cc0eD8XNOFR;/@Zb(W_\eb;L-P58(cV2SZ+GS<C>,)L+2N=-
HRRJdIa0(Tb2;b\[@2;2DMRHPAUV;_,DWVQMD[2A5<bGgTNQVS0BgFfKUK#g&3FT
(7#WK&WS55Dg3,bG>YQbZb6T0LW=\5EC,-\fR/.(3V78dZ)OH3OKW-6G,d_d#<^2
O>[AK#MTX][#b5GL&&],W0eM,S0R[XYeQO8cLGVe49)JKXOY4W\-MDOO^ZB1f\]7
TP1<5fI1O-8?])PXXG?WUUCTNWI[)SOd5WIAa,&/N0\0JeP[?PI2FA[YQZg@Y8X;
OaL74:PYggb/?g.KZOACab?)1-RN9R<NH+?Y=V7KVNI64K)L3@OF/C&4:-MPRK9U
<cU2:f4;9TR3X/Vg#@-6aJK&:XJEH]M:IW;I(^(+ZEgWJ/OP,3=HP3#M&1AWL/-B
]b+3HN@C5\U3aI[:7-Dd#@Xc2A/U[Hcf_:7(=744[OVMM>;a0#?GbR#Q,VEY\8?/
YOEf+S.G0-DfGWNP7<)g8(>F_>T-DSZJ#-ab/=c^d=+T@[EH/AORMbJbFK(\&5^T
<?KZ.W=d5VeWDP9Y)4?[;^>N+AL&-P.2D6LA:40-/Xc-P=]-)2^8L)CMG9BDGO=)
b:Y,IC194XeC<YH.ZGZ/eg+SDY)/LQTJM&KDeXb<aKPX\g#gE+DOL>.-2fB)J@Lf
I[Bf&c^]Gd0-b>R8eWX55(M4^b:SBP<)>71Y,=3UGAG/PH2#/A=&]HRe65Xd9Z3(
g:2H?=b)MS._YfFg:fa7aYCHYZ/1TKVF(c\3Y]Bg59>#;)-:5P<NQ94;V7LTDXf6
.d.(MI=4Z0d(fgB[5&JO@-]81-/YKQ(_\7,V7,H2C3L-WbbA/5+POJY61BE5Z::#
FIM48@TU^D,C[3M1+DXEGR?_J4DCLC>6\<XP@S5U?eg]02IY\_9/WVH>?cI\G_8[
HE>a,dU3PXO^L3LXdgFH^L?)7Q^ff1@.U<]AVU-PCVVg,.7]_C\;>6;aUDSL#2#/
6dZR;TZ\fMA<#><LUQGd>cQ@-D5F6T(8NP,TMY+USWEV6=HgGLYG3]b,2-)_W>UV
&T0e@;9LT.e^/O2]7:_?+M7J-YGdYF+>MH2F5<T7U-(Y^cX.9Z(A1:C4/XfX=;gZ
>UNN9C&#FUe[<JJP.X8GGb.02T5C2dA8;_0<6>R9/;8>5X-f=;0A6f>PJL+(.VPD
X\Y2TCb4/H16.6bW^QPKGf;]a;#/]fI\64P/#(C<_Xc9&Y#4:^#gKS>QSCdD@PQ@
-14gFVP[WR3;YF@1;_0DF-8W/8O0F:(gSP1/SF5XO:]Z/ggKU@<<:0487N/9IG]^
(MI(=G].c67]-&F02H@<c=@ZYZ<bF#e4K/_cK^9V?-45gfU-cO-9)K0HD.:DZPO.
[W&Z]9B^2fT&cVLI7-fVWQ[3g_RI&ZT6Ac;WRgHZ4c4J@.4d9WGMH2J_RAC8>Jb\
:c7XaFXHfJIO5;)@.<YD>A,d3,:a05E==]9LX142<]^]<d40c46_b4]^MW)N1UEO
f#JR:c)=3)VSdG0L6V2284R_FIfK\D)]-L.F1_8,@D/a^^^XXL5QVdgUZ3?3a(O]
5A&W9C0Ke./cZY:XJ(BD#SZE\2g,)6U.YY5FKV5G\\&K,B2L-SRfIC>F76c->V9(
++cORTCcKCR?G>V0;ef,+-/X3@(Y3L81[BXNDB5-7JG8CcIfd:&H6<C(6#eBXQbQ
(M2faceAG8+#f0gI2-RNc31P\a8Z=:+&29YA)O,QeY5Q_(gX&M<A-:Y^Ye7&7388
4>P/Fg3;MKcUMEU[<[EX?>I<BPL,<:MH,2.=9U;7V][4Pa.8Q?6KOLOdM\ZC5_ZC
WcWbY:[_45R[[9[6d.<]];A+eNF9,+dE:?LY2/GBOJA>=MJD.<LaO_&0fT/YWGZ:
<FI_9#1ZM3?8Og[Z?9A+A6_BY8^1GAK-NW0;1+VM)T]/JB,b.,b(@;#O,+b<XH&C
Bgg>?F7T-#[=A=P)^B9^#R_cag=_QPQgP:U_Q30]8MH8=eME/&&9W\)?F.]^G]D1
IHc]\Zf]-1X/H2_.f^2,]TE[@X+FJ.:d0fIR70?[gR.MZF3#KPb7fK@4gE8(FOWW
KP-)-c+a;5OZ//4gJO__?D1)&[=@ULH)IFNP_8)fOI3IW4=3E[[gOgQ6],N?VE\8
,NE7I&6514)Xe91]+@.SK3G[J7POIZ&Y,E&9;f[_S7Z,7WZ^.YWaDfQQL\(QA[6#
RS:,PSS2ZbdKE:6#ET5PUOF0IRJ]faY>&@5@Qd[Z[;7[#aR-Ea(F8+H&gab,eC:G
?LZ<OcV.#+&7591YI]I.UR1YGfC69.7Xdb10F8<W8aU<JgBHWIZYVSB+SQC#:8&)
MgP\W<DK-&]H?L/AP_]c,)8HZ2RQ,Bg]^>9?Ag&g#)=IRdQd^HIZaPf/Y1&AK2@b
a-]G],\@4D@G[UM/860&3[-92aa7PIIT+2:X<[F5HN#IGda\C@F:Q>S0[+^JN1DM
Cc7=[@?&>2(;>I7J5S_ZfJ>[)=9S3-),1AO2JE7\7e^J:.&E>D5RT^4+],008A6(
TaOR1KcUM//W4&=I+.V,6Q8[(T_;D-=(5F@Y_H_fKUbE@7-(c___[.&2e]HM2f#b
&]&NN@ULV0+9#YdI>0&7fDeBF5]0:G]<H;])RO/bB8XJ+GKCZUbT.+=gL4AUcY+W
+TAac=]+4eUcM5^QI6]Tb#Q4Z>d#FWORRVI,20([bVKUaZHCJUID<>f0gZ&/BAA0
.9L&56W[.T1HeC5TAPL1L@A,I+6Q=H)TCTGb=H820)_#N1Q6IMUKg,eGV<cRSW>N
TP>DH7.^-)#dJOJWd:1bKK/eD\dFHZcK-@4]QAORD)55APP#2O>JDEa@+9]_SB/L
LGce3-Z=c&/dUC+&@eAY,LMD(C=aID#2DL;69[7W4NZH<2B,B6T\7YQV=?PW.HV@
#L1#9JJQ;dROVUT4QcCM65eMF:-#MD#CW5M4C,?LB0gd0->&I?O,TGeE[A1?R4+a
#11dH/?28P1-5>_Z&Wb[@_J\eW^bCNUBMR_gEK,(WVNe?)GRC?b98E#<(+G[c1AJ
[9-3;^9>NJ1fQ+PA</RN/aW:E#&a1XfE=N5,(-?4:J@,IM;fE#9d)Z5+IDYe)SK0
Wge5@WG<1^e]g[U-F,0?eV)I58#bKP_4XE,KUG\PW[L3\d?P,#NKKN5?H[_c(+[.
ReLD\]-(?;&0dSP0Y63a0>1_YNGYF08M\=-TJ>HA&=M(87\2+?37_KX,>:c7[-cK
K-ac#&<FBN/YBI#+XSW5W]?B2,7aUSPZ_&^WH:K.?T2P4DTb@Q,@>,Tc=29O^NYY
6f9?bb92C3^XT=6\J3J1fcX^=e9\=Zd\,\U)&9?(R1JgV;+Ge4:^e8DB6-\CF7Rf
WZ&:;CTXZN&F@],6X,fdR:1c6H4A1S5UHD6D&f]4bB1HH^?HH.=#<>67;/I-5^FF
PL9dHH0>UaQ>C+IM]daSEL+94YBa>NH\.1=7\;V6<F:[W;O6=NVDS_\ZG649N(1I
)DKG)cFeCVd=H_\S#b5S[aMD7c57.QNWX4KD=B.BXcYA;MD6cQZgRXa^-<gBQ.2F
(@5OW[3Z6J<I:G32C=&Eba^\?D,B7F;B<\VV&;H4RAe+OJ/6GfPG?8TD,B34;[Hd
-537\E5I)@Gd>Sa,HCJ8NK\,R&U6FS,77IASO4A?V<[V;;^3O86NVQ+FHXGVFBPb
4g_+T83b#;;WM[?4S]&=QU<^)+4a=:B=EXC1+)KH8,WGD4K.<LKM+?d_)#B&f;RW
HY+JbC#JQf5:]4FIaMX@<IT(4M8PaG9+C]M-cBL,2c<NBL@#)OWdWMHfVXd&#HJV
0\T31@MVg_JD-M4d(>5<9b]]Fc8g./[I?3V<F;XZd?>UJ2?bRJR2B];WJBYN<&):
)eEN6+ebNQTR3Y8M\\G:QD6E]d,fBG-@8CZZ:NF7L@U@?T#<)d@HDY)@_@4H+7+g
3=2gX7@F<?SAPH<5@_,DYPg5R<76YJA.=@.#8b[2K22^F2Z_\QG?NVJ?:=,3_2S?
BBdcf&a7bJ.FU4N=f+23Q=Ef+NdN9TTE?K5-9)+/Q[+._U:<J]Ya]ZY\Y\N#He(3
?N:+/<TT&.R]Z.KX]W<VJ/X.>cdVaIE4dZR\Q127XE?&K?B^8P7X&23F5LPgf7V&
5V851K8.1Fc2V-8WP=)0U6:E\U#fc@Q:(1E]HT,I-_I5-RR>8fbBI\3BQ;]X[UO?
3V(ZUOXO5GaMW,_S6?I;#[c@7?\\T)-PN<]HFV\JH#YaLZ^KJ51(=29M-N<,geTG
2L?>R:DTT]O-AGQ.]#;d8<:N.O@UP6E9K=[D@M]7PK_Q3]G#U9@90GU@3LHb1K];
5049OM\K[07N@VYI=+7=D[Vc9H:G<g]7.,M=6EKW+a69/6Z-44E(N3W80I>=_BXS
FTbS.A6#KQD#OMKU-S-ecfDD=#5-=bE?\H+GM2/-TZC394_/cJ5<+-NAW7>ZZ(TZ
\S8\LE=ETVWXVMN\L2YEN]WZQQ^bP7R<-QCBFKEN,a@ZVY^#.8TMbOG:)N#HZ6Yd
2239R>;X2];[Bg\gHW^)GV=SPb]0I7\P/+__UAEV8g7ZBU4YP=U.GLZ_.V:P)cDY
=gE6\C,[eS]Z\P^>B(M0R(C_/],_]VPN92Y]Ya76DR1WB.0.C\R_7WY^&PJ,NX>Y
5.Q,FJ1Ob3DT:WH^DW);4WAD>_?7[=8cR(SJE<SJS?Egfg2UE>>#Rb:S^,_aJ8OO
1/:-]^Y_;PG[3H6(cDW;ZMQ]>Pfc-[Te_P0[3dD?MQ@C)&8b=ed@CI@Ga:;CB[N1
HGS9L0B8-bSI[PU/OJ^A(La9[?7_e@\a3Z,[,gO#O:=D0(0dQ7.GKSOK+_g>X#@F
C\?@C)^aPD5>LTT-c+dXeQ@+E/fb?Y4/F\PC_]a9d+)RC;U]X#AH.4<;X&QPBddU
K]5//=37bN;J;@PS#J/S1GXSFaFU,P+c[VF8=cLL[[IVg//34eD@F\N:8^1#bXG[
BV\DP_O?E3HOLD/aLf4-.66X<P_+I;.S#T0BVTZ(A5CF;#CL^)d#(;EMcgQAWCS:
:R0bW@.)7a<F;JOe1=Z5d/]/2(3Y2VIQN,cO@_?WR8&,?-V\C0OSH,VB:1FWg&.1
_.d[8HOQb^4U8&&W=E1S5Ld/QST-O_LGR7>)R?C@OY9PQD(bZLd;7T<IXWfIa0>6
3.Z:@4WI]&2N(R=H@_FVQCA9G9#Z-Rd2GL&Z\70Kd?FC@^-?#6P[PLaXFfAM=-?@
12Td^1IN;AB8/PYfTA[ME3H:QDFcI29Z+_(77e4D==IY0RBIR)W<WU>M^(9J&RP&
E5TWa.W[M..K)c4VV-U7,_eAL#ffcK[FW\TNVON]:/&fJ8;+T)6^C>^g2RMTM-2B
?[cXJ2,]^6X^RCT[3Q_c];5=FDPWMP>#:+bW(eX^TCH0MLF2JBLC&)CNT?#3^.g=
Z)9Q8W#-AMJ&JMUJ8Aed#;/7J7GV9_6Nf@4N@3N5L[SJV)2\X1EH#-G+^-_;eRDB
R50]V8/[QgQ+\PK4VZY<(^^a8:85L:T@-aHPD^S/QV8E^CW0Q1_7>#W(0W(H+M9b
QCa4#GFZ9/02bAHMEYDEWX;]aa3O>FD2=UX6P7gUR);9?)V-.\>R65eH^&I;/A:b
P#]QDRVD[N=Y93/]GA#[KTJ1KQWRU]@;+?)Y,O5L^I?L2?4\M8I^=Z[23OI#2E2I
?L5C1J0E#PYN8-,aNM.B.I=6fb]217H&9d[N\dBNJa8Qc^EBNdQ/>W#GcIG<BL5\
?.XSVeb\f__4XJ;X[61g4N6KPD;]:WAJOON5;f1^Ag&Jb@aU<8>VfXSW(H[S2gLA
bXL4\adcF:1=+:@&JH_IOS,2>1[U_RBIAOdGb3?25C/M1=/L=;++;(H@P,c^B+8)
+FL#I&;@BL@L9W3b#/ZF5D)<.a.:3W,61+Zf,B/JZ(&Sf4BN7I;PB+)STGJg201(
T9(EKg4cLFA1932L7S9B6Cc;R/P3a+eJM,A:#_NSB;09^;UBBHGA53BKH]a<b>Md
NOK?f8]_U9B\aG;57BT^C16::XYR(O]H>G(N@WbAfHBNB(+^2J+eA74)N3E\aVN_
.SEb?5:4V;NXZfR>_T?OIOf&?Ud?d#bAAF6M9,8J_#-6P&G;W,#2M6?1ZM2Z_OV(
]03OQeGVJ[N;dI>bf3LGW2?>X-Z<[@aH-1YX@/02G/#,7]Ygf3C(XAQf:XBBZFda
#M0-@O_9UTEJ;K(?>fQE\?7eQ&/SRL<XE<)/@NY^.5M2<I-ge;6@_6PU,#>US@2N
a@CO]fb9E_.+28>ZVPB]AfcJ4YTGC?Y:YaGV:.c8@=f<b2]gBgBWZ/=L]dD=UD6=
2V:8LfKV+-FC5GcB_;YQE0cR:/E1f4FEB22JY3R,KJ4cPKDJRM)<TAK5_X?JJc)1
).U_84^b_MW1&7]7]Q#W=gA\O5?2>AS\-f+feXga9?4@;[e573:;);A[OKMB/HM8
QS].V/Q-F;=>EdFNOMb2,6QW4Z1gAd0&>5OMg0AOfEX4S^,[:7R]_V;0F>.fUB4X
;RG9]@GZ+M&03(,96H:YU(ECBZ@bXF+QF5(@AB(>XLa6MYaM_:dQ24U8-3PEB7)1
_0.fJD+ZX/\GaE)=30+:I[<MNJP)72g;(>MR7Me)[.U_=-9.;DV0AJXB[-5M6K\J
d9DC;6PZ,CQ<Z_bA--F6eWN,98KK>,2UN5c;GCZIDacBI=dUK8XB@S[OcBBc)F2f
A10S.8?5(9>K=5Z6gD,db8G:bQ8\cVc<d]DQD,\[]QCJFX(HJ--1W.6ecKUB6:=O
@[Z=8L)\eW^DdaM:[.)0H65U?U&UW=:Z/+0Y#(5Dge8;7CFC^L\I-]STTTM;H,EH
6&H6BG,7bfd[fb0?5VJRfI9\1FN^8]=N[;FAaRA:F6ZP].8ge99g\W)Ia>N@+:(/
_+O-2^IQg8-^,2CZVM/O1Jc86GbH2:SIR&K<#SC@&<Zd9IP-Y4EMZES,LU;1[Y6G
#SL-24?P9e]a\D\EHYHHH4g6/&T?043Sdf;>Q&HPO\C=FgRGeSU?L5HBg]3X_UT>
ZIIE[Td32[La96-(40P+65&Q(ZOAS2UUUggI@)aeGS6(X).ebPDQ6.(SBgSO5Y5=
gf.3W0CZWXM#-HZceMLf(ZGO\+aO,@b2CVH[9FYL;CBCD@c;IE1M#7H36]I@V,5B
LD1Y3&N0d2HQ\<G7.SW+YAD84[BdY)^O+C]f.#=(H_MR7O,=0UgHOd;K]QMPA@-a
@VORP:THOfRE]2KA<I0YR<2NZ:S&/a)A;>.PY8Tg(b.^(GT_Y_XDOfG;M+.CZ;2W
dcBKCYI^R[B0(9?NO7CE[_JZ3]-5>ZR(L;7]1Pd4QbObL\80=O=P6?LB7bLZFfA=
^[g]_<MPO[\C&?M0_[8HJ\&gE\:[DU^DZOK[f<IS:OWWN;.Q(<F,:R,TN]\+(6JO
fCT5aW868bK[MLDQdRTbW8/g7K(BLeLfM?HV_0A_2W;WK7YKTQ=.]MROcUf1^)?g
J>aAfA_[.5I1Pd/7#R3W_H[1CfUNHEH)Z2e^I9I?\FPDMKO)4-]_KfXW:)^W\bce
,5-H2c1aQ=V>?K4)S6T9EGI]2Ee/1)BB;O#HLJ+T7KLN9PDG//c?:1_beGG;20V:
Y5O+P6eb<CdI3RC>Be)GMAPQ8+V8:T9DEFSRBSXDR-H9WT+,6VX1,V>M5ZO]OQ#=
cO+?;Q.:C(=.baYLW+@Og)A/]D.Y2(]eFFJEF8g40f</a[YaO@1Zb,1=9^TF/3#e
Te6fQ&8W1gP,<gE\,8,Uf9^NGb,]U,bXH)(_I?,fKF[2&aUGZMSe.6>U^7Uc<]+Y
ZZQ_Qf7Y3dd[Ob1#UO1(P5.(gc;X+8@^E:L)H=a5JEdFXMYcQE=41QO_1D6_c6^e
cE]UYI5XN3[O18Zf-cdW#_T==99(#=ACg^Of\KRUR,TcU]e?gC?K=N<P/AcT;g)-
-bFCQCKf?<bGZE[&gcG+PEe.(#Q?fgQgUQ(4aN7,&Q:,=bQ>f@_2PUe#5e39PWbQ
CX_^_J\dT]1ZFH]T0<0G=EZPJ5Y_?,F^:Pa4@V,&D#cA#)(aD\+-_<6&O3W6dZM5
N2\J=O73&P[SZVZ@Z6\bQIZ4g28582-bPW-^SMdM\XTbZ,UaGc3FR9TVg>@?gXa5
E9TT1g1ET<29E,6=[cG^Jg\<QLCXC.1[X2&4N?_?7[IG;)/CT2:@42?^C?V5(eb-
fJP4Ba\<=8cRd/B5+X0?,,+L@ZDDd3UUVEQb8&BUcIZeSd1;<8OJV<ACFX@OB4a3
FU3_#;<S5G7[.7;&4RP[TdM,_N3]_b>MRZYEcE(e;N:0EZ<G=gX5?N60E>fCIB1@
K[URW]A7f/W&2RN@FA\ePW0YQ=I6cF.YVG8&.aYU3=(&LQZ8?M3Sb0<W^>eUb1cH
9P/0TQbDK4L-A0GU<[Z&7P8);<\I]KL._?T:2ZS:K_DWL[b5N2&E^/N[V/T49A2W
\P<J[ULb^5(_90H]]58-M&IfEK,.:8cO8g_UN(.CVf1:dfYN^Nb0bM;IKHE,8)OE
W>Y[Xf[03SG5LfIA1H^2_)R<;^eBX5c8;]\T+9/aX9HJ+N&,/E74GQ=&b+[(07C&
C//#6cL\JffB+:dS<?)Yb9c:R9ac)4G.0B0?EXQV&eD+-eDLE&_^<PdGXAXNf(F5
K+E[@a#MfX[eHVP=PfGAA7[@?f#[Z(=P#&W7P.WVH^-1>TZ#@XYW](//(\EA1U\2
0?^_,F/4\Y>U3M0VC1PQMVP8AS^d7P#-A1R^g52W:bO.R),ID;KZ3Pd5W4CM<gXM
d?4bXTX[V9:THAS2B+SW:99D.EF.@WQ1^YUXGPFY]Wg]?3c+_#ZYSAJZc4L<I3JZ
J7bf]5IeAS>g4(Q/@c^RG3]GU7g:D-3/]QHcP:O0W>QY#7?Mbb)&_9edeRc5UKNb
TF+3Q2AaV9B:HX>VFf8D,8[bQ95<a?NF@W6cFc2d](+]e43adaf[5gX&J#6eeRW7
TOeEM/EMN&fUOKR\UZMf;-LGUT?HU4B+2ABQf\@NQD5b-QM4\6a/2FAKA1af-9FW
R,:d0dRD6_a::;AdHYB@/_4(Z\ZB/4L3&(57/Z\cG6_EF/M.U55gMXSL1^Df1A5(
baWg3[P4A-ZX=3,=g,8-]^<TU:9R\X@D\6RAD^ZKf,#VYFGbcRfL+]Q1IQ<JZ-_K
OF@OX]>]@WB3F6_CXM&C]\W==<[J](W^,\QZg@a(V5=H<FB?B[74dU_[P[(ZOL](
[GR,WL>?+0_]=FM^(Y?AB5C-#&UdI)F&,(&Z7W.(O]LTNB^fRG4MCg2<B]G;W=5I
+[Y:[-19aa@3I^&AfPCNNgBb_[4NUT]:b9<O/5CY5g]_0SS[<3#TTCH[8?>;I/8,
N&2fC[B83X:<J])JeS5JL_]bbIS1TOeYZQ2H:V=bIGGR7I\([R<[6gf78;d4#&7U
K;/]A)7Vf@Vb_DZUPVE.]1fN^W>T(@c^?L=ACgJd.],?6a,ZY;=a5/Q>1)]F<\:Q
6<CQ2dKO=5R@?#1^&ESW9/M+R]./E[->01<P/dVLPfbaGP(2QZaO0:]Z.N;^,[G#
)1D)Oc3e9J+@_)-3872)ED,C4)?VZG_A[e=BWLM?)NXJFK+:T,T,L]-//ZN^c@@:
bQNRaA,Ub7-OGP7]fH6b9RfMb4P7Y3TIYJG9-.,HVaG<6ddQV0<eKcR<QMeAXV#_
/-=;Yd60PRg^KE&^.F=MH0(YF&>O[f7/b<Q92(a4:I8^&;9TP,FV2^(.3T-0:+)b
GbM.Z4QPS,<C<9KW_]>DUPKQ0Q=Kc:c2RD(&?;5P[GVf;M=PM(FY-FBf[ZZa\@,G
0SR&C2>H;X&eS;NIU/T-QZMS+3E+>Z-@bf>cA[L1XUe+VLf]b78>]fI=Qcb,<?BH
cA<3M:HIR<NcHXg.DF)N8,28W?cCQZZ3ZP>+GX[0GW_;CY+E\LGW&g-<A.]Jc6CS
d(WNfEf.AUaWSR;,;6OYda)R;Z7+Sd(eJf/F=/0\R1.&CAI,VL-@XSCR#<S][YFQ
B;KNd^\[_-^402GPGf4/]C;DQ]RWO,6]4I9L/agKXgM>S8QEA\\;ZZ&F3#G@La>?
KMS\b[@O&:4=,a/?4M?D?56O+]7e<T5#c3O1WVV/GU0&e,WRJ>ED1G^S20SZgYUO
2]7XL_(f/3;:@&(V9AAd,\\\NbdO1R#?PT0B6N)=c&-HD&dXg^:=d,@Zc-R5&36G
EJ6N:WGTXIZ9Ce@#c\:QL?\\3$
`endprotected



`endif
