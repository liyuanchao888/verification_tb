
`ifndef GUARD_SVT_AHB_SLAVE_PASSIVE_COMMON_SV
`define GUARD_SVT_AHB_SLAVE_PASSIVE_COMMON_SV

/** @cond PRIVATE */
/**
 * Defines the AHB slave active common code, implemented as a shell assistant
 * which basically just converts requests into VIP Model requests.
 */
class svt_ahb_slave_passive_common#(type MONITOR_MP = virtual svt_ahb_slave_if.svt_ahb_monitor_modport,
                                    type DEBUG_MP = virtual svt_ahb_slave_if.svt_ahb_debug_modport)
  extends svt_ahb_slave_common#(MONITOR_MP, DEBUG_MP);

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************
  //vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
vsjmyNGm10arJoCMXT3RNUhz6nRwLa1C4lirNSBDrvcM+rAKArcooAVX3Oc5/2dR
yn+NFuKILEaRvg2m+B5vRaNGwhWRRK1Mvnco4pBiWsAsoMPi8wut0fM9FlwPLC7h
XXbiuh/BuOe1BBQcT+5gTxcC0g5SgFhgLF/sgWT6tHeAdMKIxEVloA==
//pragma protect end_key_block
//pragma protect digest_block
a4C7NxvKm5XedFUi5p9qTOVHA7w=
//pragma protect end_digest_block
//pragma protect data_block
peyQ7Kp7iti1MnbFhJ7U41LSnhTjHJxyeYaIl1FpuMPW3CQdk5nR5T6xugJew2AV
2pJZ8ZA7uz3PBgSW+H5y826x5UnHXYHlE/YHe7ZffR18i/2nneaSPvwQCA9o/WFy
KPUDED2ePJCLXsJW4/yPs8KeSEkwuKxF6HjgbWiEuFer7IUnQvNDwyn8loUkhmyp
YWei6ygps1Si15KscE4OLXYzXv2CSKOhU9ld1UvyKJpLepZPqun8jg/PCEbdp1ro
7sGs1rS/OuissCjlpKLpKjkZHwStbfs8SM9Cp8siImqDepR49YfaqWdC7Gr2NuTn
g7yLSZpT0YD5B6jQL85Fd+SzSB/laUvk0embjr80Ds3ccR88SL+PFio85X1v+ywG
ZaRznp+bwtrf21JKdkJcnvq1lOpLeLFW3LmSMuTgmknrLsBKMqu53TWirPu08eJg
SAGFg/20WCTXeCaIkQp0fXTzL4zRzipwgyg7KvoUpYzplRqR+ywBM/OsH3qFs2Zd
c8268ukWs92SIK3I9pdMaLtEC+E7MbeUzSMLqLNL7rB4oiAdYhedjsKPuYwCv5ic

//pragma protect end_data_block
//pragma protect digest_block
K1r/+wh++MiOpthKy1Z763uIU7o=
//pragma protect end_digest_block
//pragma protect end_protected
  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // protected Data Properties
  // ****************************************************************************
  
  // ****************************************************************************
  // EVENTS 
  // ****************************************************************************

  /** Event that is triggered after every sample. Other processes synchronize with
    * this event to ensure that all signals are sampled. Note that if a reset is in
    * progress, the reset_received event is triggered prior to this event. This will
    * ensure that processes that are synchronized with this event will be terminated
    * at reset.
    */
  protected event is_sampled;

  // ****************************************************************************
  // SEMAPHORES
  // ****************************************************************************


  
  // ****************************************************************************
  // TIMERS 
  // ****************************************************************************


  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param monitor transactor instance
   */
  extern function new (svt_ahb_slave_configuration cfg, svt_ahb_slave_monitor monitor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (svt_ahb_slave_configuration cfg, `SVT_XVM(report_object) reporter);
`endif
 
  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the signals which the slave drives to complete a request */
  extern virtual task sample_passive_common_phase_signals();

  /** This method runs forever to check that an active transaction with trans_type
   *  IDLE/BUSY receives zero wait cycle okay response.
   */
  extern virtual task perform_zero_wait_cycle_okay_check();

  /** This method runs forever and performs hsplit related checks.
   */
  extern virtual task perform_hsplit_related_checks();
  
  /** Update the component when reset is applied. */
  extern virtual task update_on_reset();  
  // ****************************************************************************
  // Configuration Methods
  // ****************************************************************************
     
  //----------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);
  
endclass
/** @endcond */
//----------------------------------------------------------------------------

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
L0fWaq9YbdeabO9tGjJdVzAbNg+essjj+jaZdekTlRAP/FXvc6oUW3+3deAtaGxn
CFj0Rq091dE0G6ubM082GPNb5f7OhO7vNRSL0z1AZdkeZl/Cv87JBMFseik9Odgx
K6bYmo2Rx/rFzvH+78ZSiFQzdXttIIrVqLrenEQmHKYcuHEN0t3HhQ==
//pragma protect end_key_block
//pragma protect digest_block
jj8BVEM/g6vEQRhn3gBYHqtcWZU=
//pragma protect end_digest_block
//pragma protect data_block
PLhIZvLk6ruFaDZbzETtaI/3N/YrIA2wgL5W20JntiMflrW0eNITMBJ9Sq4+/3o5
EE4uztmxzhNvs0Si6L4+nopFiB/DOAUhOAlan82EwyijBenr/Q3Jg5w+4ENU0ysX
Wg2okxmAlAxO0hc9fG5jNOc775EwmbIes+EBGaAyEmVQs+zNnLdkIFEglfq1wJWh
WFngg/hrsmCbptJUjUEHw/vjItsu+SUcuxn/XsuyW5+aWKNlOsEWBDrlx+43vLJD
GwLvbFxWvtO0SJcJnQsFOskBg74lB0TSkqvPGQBf9FaKUbPa9GFzw9NukMq2llas
g6rpkex+oO8WT75O/AjnUsof+KsXn7nPRajqYRZ1ODuCGixazXeSlRdIeU5phFgS
8oXmpkX3G0PWvEAYGa1fm2i1gVFKYCiSE7fKGoKqwbIE71QCk0ot+OS3+NQtYq9w
xcwEax+zdVBXRVOHs3WrB1Q7outtdemFWUPdiyJ7IM8hrIUbejTWc0710KlhosmX
++04871EjN8+AQLDiDmsRaxDfx3f6h/hzMjyXJaSq8Xd3itdOZ+BuLiu2i55Tjl8
B8WoSvU5OGgM3BwhI7Afi6eUR5+N8Q+Sf4R5HH+DZJPP9ZMtWMalLbQudJNhsZ/v
p9zXNMJh3HLTbJBOsbBZshADRLqSjQIisZvgQNw+Ij620XWci/2/eYxsIG935Xcl
6aUMD2RyqUtiS39zsvX6ufqmSJXSsLFIeVRXeGgkQR4LE5A0nWeY4ebRdQVWLsBn
S1MQODpRUGDoikS6zLC+zUCRy6bs7sgZ2KsMN4K2ek78eEWHFfEbKaA/ZRn2bKD/
XbgAzTzkSq8uS7oHsE6SaqOXmg9cGvOxOfoDVkMYLHD7JAZ6jVrfRnLvEHM+vANq
KsEJgTSbZNc82cXnYhWXvNWtSvwzjUlWJNM6FQhEq/yz/ZIH5SUfgAtBdIzJTgOg
Cq3MITrKWDpCtKLweD59Ek4jlIEFZkbgCVg9c3Q1oW+ISMdt5qJ2ASaz/URIrDoj
FyeG8yzN9IcK/AYL6y4wMPkrTx9ZLaeTVkOPV81GOaQeHyntx4/B4hS9zdivHB67
7GAkQcM6vvc4VulxzaqFtxrY6hpXjVamekCslzTnUYiUPUEy8Rm7gBUVD6AI4lJu
Sop3H6eFafX37788D+4KZvTSNkiyOIqTnTzCaQK0vpruJ/Qxn+wBBoK+8H1jq8MI
+ma7PwbPjO25gC2X0hr7/E+RPw+7w3c4EpMClug6SKPSUhFyqRVQ05NT68EhFV3R
K1R6EmwP/ZQDu3iIaKq/Tg==
//pragma protect end_data_block
//pragma protect digest_block
0hXEnbAKbLVIdNE70Wws9IIPmZA=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ZjZL6oi5Iww1145HHj5qls+ktBp18qNnK9CmLP1GTPEGZZu40O3+FySgYVP9RDfH
1wmcUORP2z8+/16E4XDJ4cdd0QKPiYZonFlGXD+//bxCKnfrEg1DXuLBen5rvNr/
fpQq91ZIsUMSIFBdFqzkxnc+URofJhFFNIQ6n5QcsMWzq5MbT0bAtQ==
//pragma protect end_key_block
//pragma protect digest_block
u5PSse2HTvD0vGJGYcSrrFQz5G8=
//pragma protect end_digest_block
//pragma protect data_block
R/zMz36Z8Fcl8cwPoZuvWxlCktBFXsOb5gyPgBK50eNdDvqUu/WwQrIrYCro6ERY
taAZMb+g1BJcQuRKgqZF2buLaYK3T33l88nSUJZLYN4L3PsEBircwtztry8QFMpP
N/U6tZDPgLHs5hu40Bja3kQDSexrraa+/y22Gixwp1drjF+d8pTLVUDMnWFzb3+8
UwAaFR9GRm9GDAAVe14DNe7frT8c4lzMd7gXOrlyB0VmCZ4sOSefOurDxCbdr1u4
E7b2j8p++P4jURFJCKCI+8zTxMzlE3PC/Pc2wm0I6DW2zsTeDFlqNRmeKIDURzYl
oHfO35ZLDt7vht6JFJpc/xBdc6UyMzmhW32Y+peDF025UO/y+NSlcMr8IKQ44qVi
eTtEA4LSS5qU8fRBKqlWHQNXxVa4yOzXAxrPsrmZfvH3Rl/25FE48cbFkMo5PYe4
Ca/vrwSVHfo4J6bOXw5XenNYJtV9iNRSdHmVPiri9bN1ARr/U1qebTlY/IVKwTXD
xZHtle6p7gq06b1oR8grAGvtBTnwHRPK7EJzIZSFG53IAxrulMoZamX9eizvM+ku
viS8lAB7/LD7l/vrEew64aT1J0wIulsZvXXBsVKn9ryvqaO64Fm5UKF5W/Zk4LQD
0R9BvFSzNmu2sMhGoIam+RprMx1QiWpMHOY62xvVA2euBWIGh/DIIBRwN7u/1fG2
gjiolDG2d6jEaLi1EFqcd/Ag2hpH7dY6+L6JaWu2CBtp2pGPTrzRZwmmzmvjsTvi
8SSS/tU3kec/98H6UqeA98a3LIIkCJVaE6h9RH439iSMLASq94qHScip9xbgbJHx
dwG/eBpfZTj42LthaUm82arn7FOlNoc7Puv51wrRfwffOVPgn6vX6oTSm2yGa1Np
AneDJlV2KQcGd+IKqDtcR6iyyAW+9LHUAL6iBJI3T4MLAF0kO/7EPg8tDai6jTY0
vNPT0ZvBipZ0hez6LHKqfmy72D4124WL5CLWE+zvaJaAGu91cCpUCgra0Z3qooNp
eGt/ik6dwf6mNP1valiH4X8HFHQzjtvDBzVGITUeakAy+O8fXsdB1YZ6GzjKowMK
WHbV9y0/svaB4y2MQMUY5NHbmy4CLPVDvqAkhgBukHPoh89rSggcadtOrxruYSYa
VMm9LFBxzs3bBi3lgc6iusFR66jTp9UggaazV4oCsgoXlbZyCu+GlCDInVIhsMes
BUjcGdjdbJtWeuan7FmLMrpOYLMvHchbKyIahsCmxmiIBfqzcJIWeuEZf7qSidIz
FP3nm7e4C2PJrtC4Cg0kU1IGN76qyi6vMnEv2WHidOot74xPJsygOln1xwpNdwPa
Xpmt3gx4J9IDmK0eSzUpdEmwVzHWc5wI+y0hUtYgOyBgI47/dhczbBQ1abS+JQ6Z
uSjX6iMI+5N9xPdFDge8X2y5vuT+N2vtLsI9lzV8FJj7FzdvMDicA3n24Jc6/Cam
hVa775b4xktluIQQ/aRZ3i+MSIx1DQnZMKMyy+B4aRHkgfHsZmBR1+QRHT/xzhVl
87zC9iahDTjO3wGwdyCKhtmLv990VOxmLNEGiXpseL6hACoT7VtDSRNyxfft4aTi
4XSzw3GkunUM9go7opvMkcXZc14SoyKiIA6q/RXALCXi0N6lnFmvrlpGhL1yfDuW
xadDNDAa/g77cFp7AstTPz4Jez2exIbStjvN64cfW9KXOO6ZBCA+S7oz3nRvVdR7
NxIhALtGgwSH+GCYsOWs+twS6ZvmmGnehQgguERMTHRdOnnpmciw8O/rKjOKahd1
YUWoC54DOJVIcTxVeLfL+rGXLEzH0x9SSjEyPDgv9GiPkBn75GzTUPp8U/K4sEqp
zT7tRzeJil1gLcKOYbwKPGM2bF0E60uWZNkdR2Zy+aZM7PrXPG43JyW/Se9cAabX
QK2uRC+UeRzSm5ajZCopPlFObdO7Od32JCJTOHzqRXX7UsHPuC28Dd1UTFfAxME0
/BWK7o/UcjVMuHmSMGh5iHB/F8AL1aJHP6g4Mms4ZC1IX+AHcpVnVAl3TRx/pkxl
/sVXH6l+9HhHy168BLCYCTz4VKtWbZxwTJiXqERyT0Mhe+V4iZJtvPPHOMqhY2ex
GowzV6kESwavvk39/x04K6RNZebwrTYc0Y8Fsa1+eTKl034/nicIDlL06FO8W/0D
CDOJNNp40MaaZAE9vzAkO73KcoeHdzD1QAnX2fl2LJADuEcpSHcHWnG1SS6L8Z5D
r407Aq4fdmfP06fZ07KIfQEff7Za6+rXmFgtg9liXWddSSuEdSmT7wVnjXbjw9Pt
UeEsQRa/FjdvimrJLH1da8bXNS6s6og8HYu6/LPLQUJ+fXlFIOsQWMB0k69EWfsW
xay4e9Gq9j988ERlwdhIA5wecNFRXFrwnqzOiPY1pVQ=
//pragma protect end_data_block
//pragma protect digest_block
vJ8PUdYKQdd4hYuf48DcJaDECHg=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
adSEeNR1gNNNUxh365zcOy+V2GF3yD4Wp+rE0GanrMXqMeMWDDAquyGFVAwDfDaD
WVKdzWT6D98hnT1Z2B7TcaDQeaUUBoFSCbDr+RxQyOh3akUjon6kJ0+qnJ2FmwRb
sIhzhQ5jtEGDCspk3CYGdrp0TwKX4xU/VwYQqzGwbnwW0F10EBC10Q==
//pragma protect end_key_block
//pragma protect digest_block
vznVR9s5Fonq6rtTvmGnmAa0i1I=
//pragma protect end_digest_block
//pragma protect data_block
zEdtPqbfPVQigHXu+K4lbXoj5VpltsXXPN+XHZEg7bw9AIffK/KyEmjqN1odgQ/3
X4aiEPQkpzqFAksnN74YXfXZRe1CCpmJrGm5LcmxK5PvFoUyIBObF842+V4+1Mnu
rdHH6iwjwq/8Y1JuiPRXrOJrqOaXr9vKjmbG9DfHyf1tMtLFuGk00gM1c8/WXQgH
927G4fShK14TM3J6nx/11MTY+FcJnTckRPE7fpHyV0abSW7Rr8lAGV6dhfVFsqUL
F31Pa96x5/h/qGih8P7DGabJ7rN9G//8+CMSCV7lujkwLV5WdaZHkpR5Nk5Sbcnv
0IkxkXum4/LvRB5wNBmohymUC/DEMuQERyJg0QQmPeKAeVUAKIZ+zf8y6w/4DmE6
YbUJzwUw4r8FdrE70dAqPnIZdkz5z/jyjDkDU1U/r3MDsNo+d4+B4LobUSnGYcVk
e5yWQozDo+63bJGJN3xTiexGwbz24eZHL0prHzlNEgPSZsJTWj462UHW2nzu6FFA
5RzoolAkEkajXqbnsuAQftA5SHYKpt7q50MeLbo75KepI/90FfGP4hSsLlL01dIv
P2ETYBUnbRAF2aABwruasA==
//pragma protect end_data_block
//pragma protect digest_block
1/SP9NXg/b8SYjKfwBCMeECW3P8=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ORmaDIqABakEC1zrtKetQOvt1SqzYTCMaYgTRyhvDr/CwpuomLJd3IxivRDWUtBy
VP+pddhLAuricSKXJIeTrboh8qSGLEPfvv/vtF7uQXoWtF8oO8fJxEGwxraichc0
HbpROPdEW3O1Z0/71qGnlk6deAD4DMPjBhZ1WFGK+/+6kb2QnfMc3Q==
//pragma protect end_key_block
//pragma protect digest_block
k8nl2RbwjlOEWmIgUOe2QuSKeII=
//pragma protect end_digest_block
//pragma protect data_block
mhFXcPWTwwYGqxZ4zz/uzTx3G3PQW4Hj+PWRQpaU0NghKPb3s5qLZyaKhLotO98L
Q0liJd6eRvz5lDIcRTzkYqrFnc0MhN+YgvD78vdHBZVkdjYaQNl3p+OvhlEui79u
CyvAN10K8WgPnJINWCNtY0w4x7ijzQpjcOipe6P7tLynf28+BYpQeK6Hagq4XiPj
12t9cKw6ALrAcBaTifIjxstr/G1/MPG/iE6fK6qV+mpjE/GpF+B7ZuuYrlAFtgTr
JJ4nN2Fcm2bEQz7gpfJivHv6oOn+TslnMFDYkpTEmAwDxkdGFc0goX8fwJ8T/9E6
CaZUTxhYqxb50dswmC7EwWxZGNroU7f34fjLBlGbJ753U7FbewsvkagsNtL2fwEH
TWGP65GtGcYfepZ5KctQVAXTn65M50hA0iYXFBBQEr2PLpkjtcPUTNKsQl02Mjx6
OwmREIM/lkdoP0hpqf/SnC5D+Phbp8SqmCWHyVaYsdWVE2bbSJafRyqVPR23LFsa
qckSggmFPHuaVVuc/CuUGJCC3keCBCyWCf3qwMWYBqlCxFgmev04cMb/yIRZ+11z
AYx6PoyNaki8OGarWkT/M3V+oiAlRZLit9WdEwJrxVbaDfBt0jgNlZC5lJDQaEG2
tovSJBo/wiTBfHnjkhtgpHpfGusQv5RvV+am2+VK+Eo1pM3t9VqHdqNyvsAAVcMl
I3bAwBzGtWFh2C4uSaPuT9jNVwiG9pTu+iqaMyUaGjxMo17a2ogunKTyht4V6Xs8
sfUJiA6zMvphAJf4w7kxXQI4pGRn0wPfmKpylWKgg/os78hI1bFbAideD3J/ytMR
Tb0xfk7dMbpSLsgpOyEkU1A/PdoVgVVpdQW+1yJfI2vsVabiKWUFVV+rV6YPSa+L
8cWaFrt99CsIZJ7/WjiW0s/edVd/rd/DiHPxT1ALfLgYhBzVOkUQmE6YHKdGPP+p
L8VERRDUKaCZJ489/E6fKNupQBAsD2D3cnPQNujrXB0axf4XP13DpOVTRTSi4pzU
8evst+ikiM+KzTX14rXEDQESw28DSDzGs+apia0pwJ1s3VDuIbdaWEH+lff6OJdk
tNkpolpXeClxDHX8iUJht9TyttXkjqyzYX9x/kU0EaDglSZeJY4JG/skO3sLCsEX
9C60PoTBD88NAGkuSucMGEACJmIodVdqakH6QHDdw114yYhDuJRuNcg2n/1lcZKd
S40kxLPHnlgPyOzzewuXJZbbLEIz32tIXlbG3nU6v2QD1g/IIewJGS6AUAqIS6qs
9TmZRWtu3GgYV8KebGbZ3pIHdBuVqQN8c1wgJcWH176DFeZe84CivR0CL8YLjHi2
FSxF42d/OZqyE6HrtRrkJtKHec7qBplGRSagVz1+g/+E7r1ZYsnqYHXM2O/DS5gH
7FKiVy+IeZLcmGUNocmUt0z8tAr4KKf/mSn2U0kChrXsb75fDBZn6Ooed4o1aKWB
RzwLyRjuxHkyFih2w6blDK/7264dmEKOcaZQgdKOGH4DyYCdNvGcN9n0ZPFRNZz6
ghIIIE5clmHUSY1C1h3oEsnlNCxAVo8doZtjGuEwdyTHhXX5t/WscI86xZAUMpfg
ubyjSlrKe8EFe+QI31jM6IwCTiannPdf6tw5bSLwK41aIKh7C6v/FeErbheNkcvT
oStZItdaAl2WOIzYY9CUc9JVol2JY2bN25d0GdrUzIMI1gdpQ/T6WI1BJWur7x3+
q8q70mm+9xnI+dPwvW3IVH0OB3v/09EkkhFaIhl5qj89nwMNsAEDM525Bs4Of2+q
UMXrhm4sFDnAPp4OTztIeNHuiGNsuS9pjgA6aBYSm6JYvgM0HyJerIyIFkEK5CeO
cAI1OPLN0yS+BqQ/8a639GBNK3b+q3hDxeQ5gdHaHNbz2AYI14AwtIsUyWOHb4RA
0pSGgTzfYwtFo2E4GyQiLkr5lBs5t9PU9lK1FLJGZt0JPwJZgaETTWJfC/24X8jI
qMMWHJk00gh3zPJ+ADtJikv6RfeYh2fHgTN3OnpjU0TEBF/gv1xSzo43yqdpPZq9
h+VK1WGy0qtjprhjwP4e6p8C/+UjSzjXhd4Oo4rradrmPlIafpoekhsopsyk2qhY
L1M+tMiJzYuL2iX9huWs7xvG1znhoUE+DFxJcjNSW2OJf8eJNXxXJFj8p1OWkYCq
mcDz7hzmmf0xPjb0ndECDs9lPJHf+Ld1Lcz/J2WQ4MaxKO6kfSCfNAfiNcjJJtdh
FbDAJd7t2BQB5jBGl25ckN3koy4S6vslA5UUIS6+TAzCSFTCbuwDqFyDe2IfcWA+
loV+oxrx1uspgPihC3p1blIt6bJNf4S4PBBQKmWftt5pwrYcFpHIuGxBLKlUQcKF
15hTDMqkh0y2RNb6zPrByT51aTy4MZn6tpY/frV9sLH/FzHGzBW056vy3d+P0yag
8+/EnQzjCcJKv8H2HhRvoOjYlLsHPvzZZQFViqVtFSLKgZixr0rx6iRLG5zrLDVJ
Pkb9R1+ZZ0Do8SBDJFihVfaKfTOIeTNF1MwHoVkeuGh5D4mGdF+WTwnpfnikSDGT
TmAotMPZfToBJZHdvjNW7UXx/uwtda8cbFGHNJpoTjsSuW8GOMMvywWNOVLQimBU
TXVdPHmejKtd0sJcWzP2OImJWB4cAze/74qWMO479mSZcj5U8gwwxcYabY2J9vRG
SfZGp5EwJVmO0ywOgRB86Hy8t4tSaNQ/4qftxfJiA4X8JDj3/i5az+rhib0ARhQY
I42OXPuIVDRTuxtCkMddkRK7latJ3Q450j/GMpKHGb2bbBqjuXKL/u0/Zgg7XYdh
bTI1cnAFASGRXg7f7pA3mRgdCAh6Tyx4D+Qra8Zz3QgPRwYlPLYLKpR4ny17WrAB
W3P2x/tKk/knOR/MloWovJZ0qKDOeVspyRARYzAtfQX+uWnT+EUHjgG92ASl3lDV
G+Zs1XIfEeAJz1s5JR2hlBF/mlOR2mPJMvINZ5genXkudKdLIs49gJAvzlGorEv0
jZNYNr4/a+/m5UVPUu7QfctQ5KH7nhYGH82oAuKn677p12wr6eLw36J09jIiQs6q
UVLCeThT9mVBhtb+L22PVckMmFwDCVn5kGSbbowSi/0mLRHOSGATHiWR9sa4Rs3k
k1Avy5+0TuPyc7GZ9HdhOEyA54SPJtqJjPmekPmnIzS8i3JewkoTd0XBlM33CcZC
Oc8X8BN+cJCYTREQqguRN4fryAQbr1Bd/nlTpyL1pE91Wjaefjd105NFa+7jGfUl
jerkCaIpaJIjlmLJ2XdjhDlIq39H4D/zqcjMmUGbghPQAJQmLi7S1wT/A325GqF9
lmsupXqCPmXgcelQffZcYLIlyAGzEz/yxeFn/edVG25ABnysXys9mTAHSp8SNUvy
drN4wpG69JrVWrRg+CQAT/esYJO6qztmwYaqAd2QsiHBZHZ3hxVS+c1HZ0XSGmuA
64+SJi0GqhHF7G2Bght43S0YNhsj/9WBuL56ermWvq9+H9V6VK46MlaPlkCWSwtN
WcRmKOyHxSwpQw2bJuT3cdtokOPHthSzDCdb3WrsCFjbBfP+VR68caNZFbmem8Rj
EX8IOzBjjU5W2VG6vVNQQT4i4yFbOPRCmTNRt+bpu/UCv2Fxmup0wOKGXL15Rm+s
cKnwAOYnJQKFVIqL1lWkF7WkOe/7O+PF+sN0c8YfiwgAZ0VsuqEXgnz8N2NIBFuZ
3CTnwklCHPI5A+c4cPIhaLMuLYON5JGjob7CRSkMnE6nR4XiA+e4IXcvfU7zxLYK
m5l92w5u07jRA1qffPWo+WpEMca8jrzZjg5YMrdSFFZk463l7pO8o/9Q6cf3tySs
YTHKfhshQfHFB4Tkk54C2G+0Wdf7BRS9TRAey3Kos+In+qstBZPlNHfje4TEi97D
oRcP7nuPZi4AI0B45Q3dbNiTXcI9G4IfH+7JRcCjI46Inify48RlxUOBdSH7c0dN
x6Jpennj1SO+zDR2ldDF9vuKU8au8yrV5VBbS2y0pmpAyMySgRF7njeWbtd9kaNp
P9bofrYhsBiFrg3ALXLIh4b1SV6LHfmdb7r6YPYPcI0oU812nDxIOc7dYJ2kgib6
8pA3jTZBTHh5zmZ+BgYdMBjmWsyRqK1a2RiORdqBjqFDMIr5XWtaHBc8zcoC+zJm
KA4bT/1l96Yzd73wTUUNQKmTv8ofx/w57dK5HTMwxVEZb9tRFuX2t3FMZTIKnfcJ
TUCfX16eMzZVgFfLPpNq1ZesplJ3YVKbKgQXTeai8GrB64l47LZqwhel57EpQB8O
stO0J6HOTdeql6BmL+16jvAr5sMvXDY/eqzopDwNLR8hG/pN3T+novbLwUzGvtQu
tbR8HdCD8aGQ633dE+EWIjgBnrzpgFT82IvWHDYHrs3PmjrrVTU77fHKmhn1QNO0
m+RxlSKf7lOg/E0Oq/5ZayfdYxznemA+N29fJGv2jjSLI6CYdteJDt7gmA9jC5ja
0laxseMrCD7dhcv6NqDqOJ03xxSRfTOIHTSgw08dKyhXrC/zpo2GrTkntXDzoIIT
tuaPJw/mPg7t2F/tLWDQTaBdUVKAOSN3+9OqIYNR+20R+HNVTdOGDBZJtL8f45Rt
CFMtNFs/SFVLEw/b2gEahpY9VqakHgIAso/3/+BNBKNU4jr2/COo5w6Wtjt6I24u
etRNTzdugNCFI6Ap6DMrDRQuppE1pbfwwWwXQqdLMsbyfB0jah6bI74YAFy/uX7d
nmufzlbichuTdg6yFTetQm63EJxFWgKA3XPltHDXYFOuNRhOAq4TBSXLC6IQO/kV
ER+0DAMl8aSTMsjBLBX2Ab12jOKAorhj/0SmE2Etc6GIfCOkZT45fFZBPcTnlQMF
TPdqjdcbQjCUIFDIfUt6dIu2+LAHyezycWnYV460bDUFiXXLH4gfKfwniGzWiW1i
3k/BaorVAnQ+aIxP7ado749h58c4HpB6hCwA/1gZgeuxWjMNcG3cvFwr3cu7cX5i
fTkUx22cDpEjeFaYW+7+C6RbcW3qpeTBr2vsJiVyRbLbAFSDIsTlJVlebsmr+BIr
PjZhm0VF9rAN9zJG+BKWFrnpj3TC08pD6TMlRzHqbxYT9UrBqAjL/q1rbRyoD517
owe9nh+wtU4CG1ecFmAp8MQDZdLys2v5bDTJPdXYZzraz+T7G8WyJHFNwmikbNZR
MGh34uldPP8vhZqdzUZXoq4zOvHpSZb4rck2jcbIXNSrYRmIBPqTgXrO9TCV5FAm
PG6/z8KqP0Dq0ba8LUUgFenSx/0Q53+LhQjohQ9ZnWL8CYZGXajsI71U7LvYB0n/
pGS7Wqmse0iLx8eNcCpyV13Rfy4MIHUw/oAFsKFA2Al1HywSW/I6mfNeWLRQB/wy
1OBmxsJtLMNnKzQ0hGGmLgSkIGJ2U8HFs/ZLu1O+4S8vRfgjBo07QQ8I8egy+N2A
boy1zEJHb50n3Dwe0b+JsD3FdvbuVq37NOddmRiyda3KjYcXTfYL+V3zMvzJDqJ6
34zxWE7J5jJuSJfPATB83KQRMzQJoo8VOMHvWBYKZ2L+fjBQwevQl97mL5YnUqxH
6I+eS3N59pSLLs7oAUsUw8WkGIg/dbzn5Sa/+/TMS9pFwlnerNr1iC2xTToysUey
h9WxQfn3+7e9j5wBaoN194adiKYHpZKnr2kROSHYGxfFrg6IxyzBnJFEkOlsiSnC
P1aHaFM28XRz8Nsc9tJZmfIVjMNTmxMHthfhF0FuUIGLZGpy/6hMLqGf+L0O3oWD
9ywew1Y/fhxq3aXZ55XxVWyxFgtE7ntKzMI13g87oi7+tHnrwk3rN/SIcSXBENSS
ZQRJAXvcHUxORrc+8gPaOGXB0ydgscJG04IiBCxjLcxu2L77WPdVM0Ap3p93IACo
ERhnJKxw2mtgS6soRL2fMXqAsiu79qddssMg8Jq5QhFYh6AJ/23NJzDTL7r7A9c8
4Wdyy1/DJWQJoY06eNO9InbAPqQ/prfvtG5KuF1/EkCOTiMx0tf2i2Wq+e1Izg4S
Uadx9J1V9gkwAaMKQtM2qSE+u/Is6ySdGePLsa79M+OCeOx6yAzsGr4Raux94uch
k/bOiB7OkrkLSPX5firEgbaaBGvl7MIafxuA0PSrvNKzUcTZ4mkFtHQcVh0GtVK2
Yy5oFlb3dPvLEd+8K1eKsfmOw2GE93SI1QHNVIg/ymB5WFGEY0LyVGIG7J8nbwhs
G2uMjqEnhSGb91uvvRLb/pUTNVaon/TQrFbnp3a/WIX6JybaDdYmpS30FUqF2b6W
+sMnyGE76VIGSCp2o8UL6HNBfDDA/VAm9Ojr9troBsQl31x8hVdleFAESXiaRR/W
8th+y9M+MLUecI79QDMxDDFsgVOSYA2hmnlRNmRBZ822yOUpEHR95ZIrKcVLd/uQ
rvq73ghdp1jPZG48oV/9m/VFcRfdrV9STFOA44E+bRl8qxiYAfqcu/T98hxST2TY
XvyGVi5y/3oJF5PoB18w7aprpWjl2WvLRcpaZfS/3kmMVrj4426CRaTcz52vSoxQ
GZ/Kp0lcDvJ1S35hdS2BbwQoXhAfLLm8n3519u0wM1bbAX5FsLiG/tN7XCYMWgLz

//pragma protect end_data_block
//pragma protect digest_block
en7q3S8jTvwAIfNZtfce0q7Ew44=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
lx8GmIJUxiz9/oj8bTTJOpj1yJcgYOrmGh6XbgvEq2GWEMErCpOpf+uI4bJotHia
VesMqgutQafSAtYhD++3O6pWzgx76F8yFPv5V2jUu6HAK44THT902714VcWyBJnK
phzK3F9rmLprWzVaRr1CxyE1M58Ob3OVTXsYjhhrZqwSxv1DPzqLhw==
//pragma protect end_key_block
//pragma protect digest_block
pmnAzn+53Z8vtgLmjsMstN7PRzA=
//pragma protect end_digest_block
//pragma protect data_block
vX8UiFfUIop/Gu6ymgi4i4+KAEeP1mNkbyMXHNLaeVoet8gPfcXCCvWx6j0Qv6ky
QmF9V5JhzA2VR7Au1EMND0NnH8soXZ66I/uaQfNxPeQPplOfyISCzgkob/pY+hgo
VUgUskm2M1Ni6U9t69tjwqUBqJ6FyS8a10yyJ5McW/TDytpfg7UCFpbFYJn/x2KP
79ebxZ5LUABkeQcfsDlrU4C5fwxsOyPv+oaRE0wzekbjkTPxf0ahopuf5Ygtct6Y
awTYAy28h7h3CtKRgsC5mTv1jSeAMNmMEniWZjaIQ01YzBffTyEKudruX6JS+4pb
pjBkk0XQTKenuCqvZ7LLSQiQ/NZI/B+8+BWW1yQmTFjpo9UDTTWNsLnAkIPtZ76d

//pragma protect end_data_block
//pragma protect digest_block
Yw/BUgG83s8AFY0LrvAoX5iIx3I=
//pragma protect end_digest_block
//pragma protect end_protected
  
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
wdN1u+V0tNb/+JT0BfL05I+QoGruTiRiFHVZdzNh5dKetq7CK3T1KZAt6Y16uUpT
x66oB4/W8t7aNCZh2et/wpKBWXUrGrzgRbA358PLR0X8ArGPwReCJ2OA0aP/YEDs
UMcMoSLqFOSNvl6lHS+x73TpKqHNGKCHZ8wM7rUyHCBer5AUK4dozQ==
//pragma protect end_key_block
//pragma protect digest_block
2B97DivTNp4pUYdyGH3PmTVFrKE=
//pragma protect end_digest_block
//pragma protect data_block
4J1VL2nRTvTVJVaEow8hgtdkOBSXlpWWO6vlQ9gdomyX2byhjchXUGmp+hi16og5
A3ig5c4lUgJPB1ci2Zqizf054Fp0iriZQeD+6hh4BEuiV/Qhck/gCX5ZyDctfEY3
Ii/O1UvEtO6o4klgTSPkgxhvJ2NPlLysoPZJXEZCDihfN2GD35p73ITZZnbqHjE8
4tH55V6p8j10yKq3VIYgouZkXzr+V6ZyBiu6HX30w8wK5V34ZAW2aUjr7s7TX7qw
hPGDPBOrcIz/57eQiLwaZkvB7F3gkSHUDKsrOOt7E1il0iOdar+ckGwJMf75+1E0
M8S87LwFcTPqp3RaUtcIXR2OcYT2ZvvZ9F3WqHPkitd5zZZhLNgEzfYJnQ43YERy
5oFlzcYP28YUoxjdznBphek4Mc8h5Znvb6HeayJ6WFD23x4jeOhi9gJxoI3BEXB4
JWGWMGTT6wak0kPx8KPGkHF8QA/bzLa04IVssQSCS6RaGngHHPmMnUC/VA9nJApm
RkpW1sAGGILLNyUphSdS9Tq8jygTGIzrdh9LFl4HrGblT40qJ+KjutdqRCann5Ul
xrBWbeoct/C/8fS9SLR5s/M1ckvCIhH6UMP5ExG8kkiVY8fq0Gw/wKz30e377Qu1
7tbZapHLnDbIhGL7BzZI+z0x9Y+zPcTKI8Y431uhNvjN6CQfEif/jZ1z5ibIpVmO
j40ZSqTVmG7yQi1WshYM6B6vWZEuzMzuSqPpxbZwwvgOWL0+j91fP2VQv3a4w+pz
s45HL4pnGxpBh5ntIQwgZYw8yJzwooke/1asQyG0s8mwosEAgLsBthKiGsYr/GUO
SZ/bVnnP05pY4QZmS2HVX3yunhrs4yBOd23cHi21IxFtYl8obX2UhIIeI0gyxl63
ryWt35cQg1279/y5ibsYlYwSbC4YjwHT7oH1z1IPXfDHtu3+dbDI6n1ElDa88wTc
+NeuQRyEx3dIbsGrTA4iFq+ni0FvTp91OS5jC9iyqDnhT/EERuAy0O4uVJ3TLq4t
VT6n64HAOcxMyxBTdSz+ZZCJPbfZRjkiX3U9fvMDcBmdp0o50eKBBo3YJO+kD1dv
iT29ckyCke3dVa8//hcncGk+tqan9sqcQ1FXW/qFSKLqTC0Mdcwczcm5w7M5w8Er
757UZgjKcATzu7YcMaA+Vs4GNYM9jI0xr1PNvsjLDdteb8Q3Qid4yS/QDEjD5xVe
xpoiRcLmSl+/WAE3mJKisQJGsqazo2k+wDe6cO41Sb5XUXzyWxJd3rjdHemqbSQO
qQ4Qtfq9lvJjnypKZgFygz+6YcKAbRO2wEqIECv7ydhKOpGC5YU/5M4hDLBwgxS3
WfCAJBBGAcAfklEDJ9sdrb6JLX+9u43bPIJCxvn+O+5OjRw/FkbQSXUfip6Qu+VN
TJcSrjlZ/HLZQLEG+lU8Aqjn5Tkfcx65u4tacxljhnGVSRp+f1lMfXUW2qwn+oh/
sn5tbGqh6G+QD4IPH/TUWodbFGsBXE6AGRZQlk5sd5zMUWGQrCCjJ+Zv+tQxQI4/
2CXMHwsyfeVNeqIypdPnQrQfgfFepPuPiRzfPpRSuKQ6RoxPCAKbVU9spTrOzrkS
N1lrfKGmhKlq8j4CgbL6ux4GcO/BzBZENYkW42vmO9I0yypusFU/4lzQb7yesNVZ
kR+ewZI+Pka3FzKj65KYbNiqT3KfU9FExJlNfIj07zQt8bwESY+s1M5b5DEEZHK2
V5EUpEsflXoskLvP0gUBd930JQ1QVPFBjHTxHhipheXG8l34wI9iv/EC+3VfvHS+
/928k3g/M7A4CFwY8jmWxZGp3GtOKbVrZOpZCSrRTiNu9CwvTt2MXFd5MdOa6Sf9
iv3aputXSZUAHeDMVi2qSuE4jC16icyMVfA/cr1DpNrX5k+1Sq/FjgffUcSdKCS+
nitiiJS+/LBQmESPWGs+Z+XAxJLrJWB3mOqdRhY46ElQw9C/Gg63MP/EKFsbwH9o
iAt7898cdRNyls6JzmyOPhdpFFim+jbFJWY5CbisE9RGMDCOk4NkRph5Hhna1XwP
/R8hZ+GjhI3JyoF+s36ujKt44gfqOVlmjanAYAmXP4qjGEnKa/9yGcOyM4Ib+xTm
Am4ehtZC1ofrqTF1KFSmC9MaS6oq2g3dPfe8DDVmPHKysrzfj2wFkGtXTI3tjNYx
bteT9ZebfAylK9F7sIgtbR7n5Ee3jK5CpEifmy4MEKE53hhDxwheUsoXyhhUObsY
vNx2u4hetpR4Qti+mUMev7LIL+AjWuoCp9bOPedqM0Gs7/DIzHaHGbmXqv8jyjLu
kzEWzhkxvvLYspta4BnFgPzx5SQYgjGLcs7C9m0nI/9xebIf6DySIBCFQyvF3E1o
zUkXgavUUJcfifVy0e7LOsohdFzwu9CaHoWUArPAhTX4k3g6qYZPjBlbmS74C9/e
cUo3errewR8Ibo+daayQHjlivZuImviaqifXbqhDlnE5XC3eidiWEKLChRc4b+00
N7l/M7ycpfKULk2NC1cZPfge9qw9wpSD2lcyzpnMUpAIhtKbzNH0TL6x8JHytjAn
a95LNPSU+wM0hqBs26494R6uhGjD6kA8hrA74esH2K3BhLqYrnXd3uARmdEt6V25
MNiZ0/P1QIuUwBFH2xJWeEOnyDHLTEwb8DUiNldR+KfmjrRhX91PoCeyxyWZeok2
Vbn1pUlnfiBdLKY0EsoPpgb0L43aYMgVTMcIVksXK9VZY5Tgy9B5eTvqYjHO/rQJ
vHsjqH3b9Exqo9rzcF27c5cSrv80HUHihCd/mazpIqf9B0lX7SKkzp4mcdFZ4AQB
9VSE/3aMNzT8VYujFUrZ8zo5uOZIFIXD4PD9q8CS8Lg+oaySa1R7OocOB/1iP15x
NUOuy4sJTIndDX0xlFSBluAcZqqaX2LYrCyLBMPvyMJYqj7aT6lGNBo8difQQXEa
jZP55vJYrVjwbgpn5/qBRlTzRonClvpv5DNBqFpeJFx9BpPPHcjFngPsuRGcemWg
itcDhPPliSLdS75THAMNKFJKuyk0dR9lebtGDnlgvuoixv9JxanFrFQ/OjS57nMr
q1/vA6PsePAf5ZPuZxKSQlTz3PKGp/qjuWgd4pPe9J8Nn0At01CO60Z74yMyPdOz
x/m5L/j95xPV/RQbkpmrVKTSi4/6onqSRQowX4ehFjNBxUZ+xyUqhtxZ//RKmQtN
zj5slS94J9rWNlqDxy/VHEM9jp0m3P+267LZ7dmnS6WvTpXCEnEvpdrAX3utdrig
g+VPbkELRRl7a89r90GA4KagaPaAYxdpdKiPp8OfYn1hpSt60DtCmbjJL8t4ph08
/ksyF0kOlVz6Qp8Ue/zKUQbcf+MtUGi0f6KuuWglR7YA3ggEJRHQNwHbOdOib8fb
DMRKatGwHkQhvya95s4lqoaG6KmDDroVLvmIkqFQxpprCZIge1nXqUfyVBIA9/yC
fU1XmEPQjgdwNYiOXlbTtCJLAupTuuTDNjeOon6ABj02x5pi0WjcmJp5lzQ/Al+1
mIN8Ya5Lp+FlGCCRoc8wVZwAh+S0se6voi7O5H334OJSmzsvY5rQa5YeqVbk4mmZ
PrCSD9Jk393UfhurWRERaWX36KiAHU3NlW2eQZWnAwYyfxlSD5d3c3IdhwqBNVq3
sUDWXk6SHdBnShUPrUQA44j/hdZ2jWjAjeMYzofw/cPLyWeaJLvxpuI0SO78wuPN
E79Bk8voyLGjGEQoMHwiAwqSsAfr6epRzBnX/DhdUobuOZ1QEAp5AT0iBU59ZGfZ
PXMFka30SpyG72x7ThXHGrHpPM7VlyBrWZt+lUtXQITLvYpIz1AtpPqU1E9HaD+i
Za3UDSnfpYWCJJ/eAVoxknj8l/FKpiSXEuW0QJfC5TG4zbiPN2YP4ilmpERhWGpk
TWEDRWJBP/0xi/lj4oRaliVdmPoeD8ojyA5njej5gNyJShG7mWlzfr1tsEBViJes
FmhwdQw6nk+EzBmk+kVB4Ym6MBLYrACtlTiVb0nXxrI4fOKSUos7iAO0JDwjIxo/
6U5v1HULv0hcSTTdaHEEJiaOWe9893yYYEzKls6ZwunzJ4UmH5VClOgUh55xwsFb
qUI4UAFR86FU+wFxqPcdUWyFrTt3z158GeaKFfYqpwIQrO3dKIPGBg2IKggzcZ2t
ISC1wXIq34FbfnyE7GLFpbEs96RM8jc8P90ElNC3a0NCmgy+zClhm8bTL1oYegKi
bNZvcGS/o+K9II3FJ2ophw6yyCe84JC371ZsiP9oHlCLaT62QhHkS2gQeJIJSeJX
81MG+PXUuKcoWXSn2xUdVc4KMwMEO3NjsTtQCZM2xLk5XqRhM9aIZi7n+NYBSxML
np7/Gr52DIS6NsZgsm6saIxPpsUtSedhmRVExK/02KXmaoPStWDi2F07ZfOJN/q+
xdEf3jf+AQMaTbsJTQSCCmvPsbxJvhw5OdyXtofi88IfhQ8neOoGUzZGHsQ9xDqL
oHPl6iPMPub6QBFUyqTb/ccdDY8vhgqpAkjjiaEP2P48MS4lMt5uqh0v6b49IPv8
L5nK22w5AJQk5JCuox2MT5RaTyB7v4kDXF8ykcJnjJdBBGJNh8Qnm3yGocdzPjOM
mjhDCxqIckXHg6whhp/jKdQMpJt3jPXEInadqpI88Co0DHUg4+WiBOweMqOyQMC6
APqnoW5SIogj1MQ9Bhef/6vGGyijxF2orTGRZdLq2MoXQPhyTArDY2ozfPuWR9Cc
0NSk1IpmWjQlja/OVDw250L9wT0F+XgmzMlq+s0HQGhDsXU96KMfDHcrov/036GT
Lvc831NWcAo735NS4H+R7Ho8+zYQzioLbjCgsyf4b3wOpx3TmC6zFmHOej37uQkU
XYOtJh8GNi0iUScOcWqpYPIAdSLUz7c0G1RvdvadcAFzLsqv/QpU7QGQ/SqtO3kh
CHzPvJwbokvvVnxYF67bAidOSCDZ1ybQ/pkb6bisZABZ19NmO4IPU/9sk8aJpkyR
JrpOQtUL4e9+0o/+N6V9EJHb538H5OHY/x0cLUA99fSDXC+rGOLzNW0zvRTuh+05
3LQff5KHIdqLwpB/+0FJMQS9gwO012fgDFrwBgzL7u31JcNumzFkkhPx3VRvrZtk
W12vyy9qLmAp/NwsmLl7mQJojSX5vPFaCTH7hRGDD6xghbECsvXIkv+UMdZDP5yW
GX0ANHJft02Zg94NCXo4pakEpTln6WYSSRRWrF1s3xlvgjqJJ9RLahVja7NWVu1G
Ur9IE4Hg3SzrVAvM6fwE96HzYbuMCM0sWg4FFcUbTI3sTml4T/eKzbfym+j6b2uQ
WyixFPjHVrRb3P4vM9j2aOfsz1RV6Q02c0RetPHzexqzWmZQzH4ePr9sHRVX16Lp
CEIgsFZVvrlRtNbE2q3xhH3z4MNneu9LcVu5rF0ERrsEN1bam/3k2PJmt072ZirR
jtdRjm1wlxSpcYae/wflOHg/xZqp5qfJHeXmzfmQVgBBFRJejfFkbl66wzKs1b/w
FfkhDGLj+dbwBEJ8UT1L6fwuty4ta+YoguSiWlkDCcfTxGKr6zBcGP/YC4fxHFsQ
kqKv6q74oBqhdPHdMiJcUHHwvy6GccEQBDMd35vp8GCeKUKKCtjEerJno4+VkkDO
SJyW8RNvSooT2spmjmnmaV6P/qe1Lfg+A0UnASZNRrc3qAM7JtcI6FoWIH8XupXS
Bx3TzgaTRyVx3rKMoZzsaKse4oKNp1kXSvQqheLffy7Sj6tYpuD0jLFzzS08Ot9V
Kjk1gdODTJ+mV9hhIWFOrtC83JDcyEQtycV/s2/6MQECHkiaN8BmyvOC6WcFqPGK
oLpIh71WjTbsHPZnp9m2jCqyPZZ2M8Bg3NsRXxy9IcqcOemyKG63BA/xI9RSXeUy
eQ8vqSdUQPFDvJUasJ3+1aNHN/Df7w6fi1N0fd0QHdLtAL8ohCDJb+Y9VAwzfWv4
S/3FKF8nilQpBbSyIH54mo5leLl48fsfz4CHbno7IbNrYagQdjt8YK2JcLmc+9mx
KDZLjRBFFB2b/5a+7l4JPO81LpniJVnVeqUR1zyjltLCqwXR+3OsLjsKfKGwLSmF
YoUrUn5HzvnDcpr4dqU82sarxpMPTSexL5LT4bce5UGrYq9gFQV0pc8zggmLfOUI
nsTdBgmd/Z+y+C4x20K9E6Plym/wG4gPl3wl82zyl5FG5nshpNFeNG5IngVVjj3W
NWZH13VPGrpZ85r3Vd3dISrXrorYFqUErnKIUivKlVLDkQHbLOxUpzmJnSRWqF89
CtnjI3MwrYXhKMZq4CgR1+URsbvxDomN/B5TjP9MC1g27UwYE7jKd04DE5+DJG81
S25obR24Lwj9awN0WJ35xxPYSJ4gOUtAkmONS8LoFTmDrqitd9O6XpeoBLd4hpZ8
AY4aAAbmpz3p06g03IgnCAgVBOGOW0X9eZKjPGsOx+hLhMhBqEH8vU8lv9TDDmU3
29avGqq2hBApeWuTsTgQE1P18L1lPYENH9CEXCnewirYAhDOs7IBS/p1Wsm6Zdt0
OKiacfXn+vvd7xFgW5Xd8q17Dn5SPrIlMMb8ONAQcK6lgTpHCCUJxxS9p+Swy97y
6Swm6JAP96PbISUHo46uR5V4P8Zjud5TwskasVCw+Hdv/3RCh4P9QRkRIqpMRff7
ZSFp26+DjIZmoaFFbeEi2CMWw0Z1du73qOnDcVjxB7ry6pXInS5/2p2jKTKj2Ylf
41KRMjKzAhUh4iPfEJ5QEN8J8AiiAKiQQX6DkizjxVsVLftU5EywZ7NK9lxIjiCu
Td+Oxbf66DTiwY1NmGY7rORjG0iE3Ws0bt+ITEtyJ6w24IChEkNyvinmjHY9BXF+
4nzgplI/neBWERXAKDmzoZ0nOGvXDibmQD5wNx2F1O5vrSK/kY55jgJJZ8aO9SPi
Zv3Vh8Zski9pfipT+Wy6ui1cgSMjIGNKATm+ArGIMaZVDxtc0n6+hdffNp8yZCN2
oxX5QLbTtfjsfMkps0ihhwzR/wYmNkQ5XF3P/LwFfUdnIlB23KzKS5f2MMmKkK38
XUMMCA08qPwH2apGw6FwNhKZO/jytP1a5GZ9l5HIQhZa9KExzzQ8THnGeIjKb7T8
biTXVT0PuHHbCypYeDLPc7tF3vPMKKAfkohTayq1vRnoj/CiQFfPLGAUPwCJ68Rv
/hvva8QwqAt320q+pIi2VuUUUwIoLAVByzUjFKVPStXegVoWrN+pNqpP7a2tf2Kz
PCWV8GyxAvfnt+6oyzlg2X5bmEDp4lxiXOBYlJ12O6JhCvKcG6Ys0hL7Hodb+DVC
7v5efZvlhLDSQteFR1Swq8WgrQh28I3Hd1jI+9DjTzZ0qHRNsmNMYejufVmkv9jZ
iuouRIkkp+Nba5eQarGiLXEomnmJ5V4xqNe6JM7RfeI+RKGatmKpPZig+r0CT+Er
IHUg808sd8YaHUUd6/WGlxjsUjyiJxwZQef4TVzzT0wa9IY687DyzXz7Qhz1GDnF
Pku87+t+Pz9y1t+TVfvpQNx1iIirPvjioKfETlBJIDl4R4lzbNQggB3J0oY6Jsz8
jVDHMbPURIT2fEhAyJrJt8wlfRKILmIutfMBZMyZ5lBPlMXQPYcINKr4+J/F6qso
sP0+UGX7pwehTX5C+zbcu+Mq/49XanxOj2M7z+3Gu//CvaN/+fj45VYzATXzXW+1
ye4V/lWMuYHVVel9JdqZ1xGibiBxbyIRgn1iPRiVBVECgYO2RMCzie/paJ9kpLyF
5fHE04aV53ZhEKNhnHdA026dfl9k2D500sgMfS/qUdeZibKoVeax6bpxYE+xHZbI
1vrqeFf1XYSEl9OOfjRn4/Ng9DNyHZspu/KzeqPgaaRdRDFWnW4dwJ10GriebKfG
OjsCQbaL61cKvgS3iWAThXf2I2Lt7WSATzF8iTl6H75Gr7UW3PaEaWKZcURC6e0z
E5i+JhMAN1hv2Avv3w73k7l3fZ/8XSIlFV7Olh2GcZRN4MRpIksIZup8llwwXfzr
++bLvQ5HSKQaeDm2iG/Zibq+1Q0euVt+QMcsXbbRY7de2N6N4vHM7TCtXkd+JZcL
ZKLaF01mAsX4yTNP1G6UkqlVdhuXP/YO/+0opOoT33jhsnX3RI8Q96rQzbNvWnrK
i/TMQXSNNv9ateD0OjzScLQCbo7N0rCGMu8qgxAc2JbZ2eJKSiyf6Z18WTfUjdil
Sp66dOugo1jLqHrJcijjVb19uolwh2b8gSojNWe8dEVASmIiVckbSjS5lM4TbKgP
AxHDBxdbLgNky0UrYiyfAzpeHJQoaZsZ9yHZy6FH5axt406+k5QJs74z4TItHePx
Je+2/JLS3/+U14WHk++7y5gIqTjIup7N97TOM/powcQV8GMuRHoVST8Im6sdOhzE
j2qp50ZaGul5fs2UBDialctyJkwhzuLOvflJy/v4HzMjhkZUW/FAUArfLKaSUJW4
LCL2ssNaR6l1VWdANn/RbJuk0MFhtZDaDAuXQ0xnKL43Wk0BQO13usoGbQt9XT4y
23wnnP75FGVstpZsDXJC7eEPO3978Yo/Xrb/TPW+lrvnfSb0jWLsw+mTTbYv6X3L
4L9SSOovuzHK2d/u/tgJKpLIKS03NKWOJ9y4MOsQIXEOG3ibh5bZKqrQeqIXwzur
KDatO7V6YzFiSYB1JaAimLCr+gstEpVCuiHosKUHFH79yVrFqRlF1DCpIZhR87kE
Pf4Bhb1IXvvUo1YVQDv12gw2ydRj3V4BAzYnEQZacoPRw6qpJQhRQf1G+K0VFzoe
Qb4mcgidfmG0JdzM/sz2v0uQwRi4cYjXGU1d/fW4T5bWwOx+RVlnZOc219w/iIUF
CpPr3WoNSN2g6ufedXXbRuf327hXRqorfzSyZ0A8a3FSVWPLPpuCrjwobAComSZx
k8CrMJn1Jmn4HLqDMcLYucv7hNqiJD+Nj6Je6z7BYYl1Q803FNXdXvqZrtIc75G0
jOoGCCcIovLyAMO2FxUUvk+lPFJvI7in1De+bKKUWXiKRmH9Og0jWYtrg/AtXyL0
UDquYR+k2xUXTvyUJGJY5l42zFQunK79y/CmmvW/+hDQoMX9lLcVHyRfhXMlgP3U
uc3oXrH5/NV7xkIN2CvWOLSvoB0S6UFkoAYWADHKuyDSJViqP3A3iC2YB+iut8Ro
FSbDVh+kKRKTmW0Fv3jIGXUsUpyAQuj9x0xAo1UVBQp9hArQb4Chz2dKvIfdaiC/
8l3D63zqlclXfdvnYxd2BJ47Mckmkr/+89NfcwTfGezAHUx0j7QniH0JwRkbysuC
LTGGMnAz0pVY6hippT+M/DYcufYJQkJwo0it93qU5fVGUPs2HWC1BWhEsd5j9SwU
KSaAD5wVjo5hULQB7f/XqdJPye4fxd3ih4RqvBdxg4fs6rlNQATBkqYoNLczb3AY
qjODyPWz+JrhCoqqJY5SKCqeHHXTtupSKoncIprVQSIN5fj5cDoKI8CL4QW0PFnl
1XfJbLwWd7iW1Juot1Irk/PoSV3PZiJ5hhSyQrTkPwFHSwdvnssVIwjipolgjfmb
5Qj4yp2sWZneoWzdZiyNeBWW6ikcMHbY8HTb/1Ib62FIM40E45SYwweDTRkIOPdA
gN5zKzZz31O66a6M7PFrxikRFnJV3czqzILKgZDiuPH36df6clAM0PdKX+hrZfbz
aBqDFcqNj30oA2GRz/pkwQ6FRHQGIfbmg2kQJ/zh3nPSMmP54Ew3xpeMbu8eBXDt
uLB4rkQv3qGgZBtMV4hjxCXIQl/dRQ3q+JVgygVdgF04//oTdkHmOLQwF7JD0/xt
7aYujqtGieVfCIQqEnIP6cxx/Ka1g4Z8cdx2ayat1/PPZudZ7VRz2+w5N/litu0l
ByOaXtDQoqLx+1VibDW261jbs7grmtjAZIFuZ9Pglv1wqwzT1IaU7Pw9d4awgO6s
TSidXY8F7xCbKrULyfyv8Z6MhF83l32bxRA3DO2vjzl9G5R8CUqDcOrFqHXAJVZF
r74XWAl1VreNmBitFTv0/y/iyX66OW4Ysu0+x82TddXxJcsuxUDoXmhcD3doIOwj
MNS2UAcaGrfb+oRXok4Gc65AY9PYoyds8JICKV61O/r0NXfSEf7ACMvcZZXxL4Z/
byDU8eFXeq5xPpiftzuM8VoGlXWD2IUgjxD3kXxtVmWDjX3QR/yuPdpnJ7I8D+6V
GL25tRNh4DGJlWcF9RwAmHTOBvsWj+xaSE2pNQ1TMVPaj4BAkOy6RLpmFuL1a5tM
dqzSYtBmKuzh9mdX1jfjg1qGEwaM+wR2kZCtC0eBdQXGOYdb8gbza5jVu9BsUphK
Ol2jIy0EeQdnGGlypdLe6/k+ll2R5cZHfbXSIEc8XYySAcmEGfDvofyEGlpkA/h1
3baSKHfGT8Lu4RVAP3nvR89wTm2h7pdHLxvIc7GUdRrkz0L3YKkvFfkBcpryAH4c
NXmL5hl8i67K+yo5uRgW5joHmaAtb5mEkMAP+AL1lcSFB/YuTwu46OKx044yDDlP
H3DouGZxTjm5mCND0r9ncusJ8kSVdBiSEKQAWxdCTKOJEnWtZ2XsIAajXiUDoUL7
t8u6V85cXw4NfEPkUrPK1qq/MMFH2jExAEim1+pjTjkk1hRUlVylZCXotCFhMWFv
dl6zEun/5X7eaoBB0geRQVqzOP/dGmCr5K3nXrUNq50OOlNx3zAHGpxmbcMtC1ba
Sg+/3qmGA/z2r3d7ZYK9RbQYbivlD0ZIpukY79y3qKUNh44e/K9kDQCe81N/teud
kt1e075uQLsWbwDqs2fHNiFfDMLXJl59qzmGE9qFza+OhmtYjV8Bt9r4yNfz9yRm
D6ar3fWDmej7kHPVlncohJqiWxUYZ4uO5+NBNds+tW/zM34nzlWmG7o7f5zT+FMO
ydMQV0n/Y+pZDUdbhMGZdsrKYlvSF1sonSlNA2D9BIy+PCbh/nAKylAqeh6CEwBS
awztZjt0ZbrTIdkWd7scrBiTzwLGlzcbyAYhMBk7++qPsHYQ2ct7W0T1pgsZHvMW
s4gVEBh/W/d8S64vuObnh+y9NTnqMGd66ju1/szMzsqxqHc+Ltl9+mz6xAkK2r1y
ZDq4FUd2FS35G2K8bf7mjI720sPQQCvRe6UpVtCoXnBuv7kOm9cB7PKUttzOVAN3
NjCiCEI8YBvEE5J/gpQA12EqDRdgmZm+KW+5ngQPsPCW1ncWo9x4cEfibU5dgqoS
lXAAanHCeVvZo3LRm1IpPqvNFhNy1zfS6hRmzY9HqabZvdDtqvf0HRM8rCsBilph
YLBkIaIr7NBDbzepSTt9U4gr3kKV2sEdSFasEaF9lpAoiycRcUUIsLjEGgcKW3gv
AjIsMgDmjzvKXI5uRVAiKtTi4MUEwWnPnLlq5sKAL5AlWF/Lk7E0BTrW9ZLEncUn
NOzZKlqy7MdBRxTK1RXD06Pg0sHaPeV19SOEeU+QRAjWDdizbcCDGROEnIAbsf+A
n9gv6ph80LXMat7flq0R8qWkTXqGiXRq30mKF/j6gNTwUhVs6/J6kwzm0sANI6KC
pPXQz3j83HPF5P6OfYBLHHwxugj/nLz2x3j8t0tM6GiQfe03dN1z1AmpD/6R9OfT
5YvJv3Fo6wYE4MRHnisSR3cl0zHsZU3ThbpFOFL/qdB9C0EoOwEmw7B90l5WtujH
pXqhjsQlXOl+KZy/MCM+4Ka1trWtjAr/TV1x72NqSjyqbq/UliDy0nx/rr57WZBq
KZsnyARJlT3SyLDy2HxkX/BmzqByDHPhoDkc4kaifx5+SKOWKp0fvpFDLOkXJcVX
w99IWPcFoMRE8esYJ2atBGx9O7LH5bYA91yXNavX7TbMK/5VLTcpBLPt8nU3pWnL
FgzqpYKopjAb7+RnK5UjGECur4SakJcvVKouaPdHOkOMKk9EeS87PZeegbvgMg8C
bQqR95gybWi7P6+UyB4HIRh0ULRXBRm0QsX3DF/6gN+UNlmD84V4CmFVmItGvCWu
oSqMRzFLbejLmuCiFFWk+GTuBjBt47uhSn31fDIDPhlWucGMDpOsq1WheWtj+a53
UjhT4X24J7xhoky8dGnu7SsB79pDqWMTm1L2Jzc4bQIO370RgXF78ve9kqZeEq1k
hrGGfwpkUL0iK+wSKQLvYyxpNmvytxSaTFlJ+aawVCsY4shNLOzLFNuVg1Y5Azv4
nCCJMm9ufDYl8L4LOu0BCex1MdTgjBTOujq0OQPqKtTdxdWDC1QeEW+7Pe715dyl
DZ+F4Ithi+qneSMsA4jI15tPq5gFwpRTtlz4hiKwVQPdPcZsanG+uxeN0AJSmdXu
WcMjtMxGzPkqJH2lenBno+2ZeMANsIOj0pucvGXnMYC4mkgajiCmnP6+o+YrsIhO
88EKj6Zf7yu2MIF4usgDUP61Dpq4TWn+RSJt68m3gKWVpV1XqQFz5fNYaR0LvZUB
KYHP5xu12O95bd99FHEdltfaxDd3GwoqmGxmZmR85UL5uOTpz9FfwBTRrBOQdaz6
z8pO4uDJPWE66sZyVjJC0IgGAfz0/zw3zrpAB7Vnw92XZMXWL6gcg9LEYd/YYPAr
m/vJpHP/H7azaLDkxFlcrNs94Wzk5M/Ftt6NrO4xw8L8N17G6iBXJAR6WyPryGhS
ZRBnckDMYWBMK9DHqtArviHN6Ct2+6Vh/Qcx74Ey45Y/Thv1L28Wx3+0uIO7H7Yy
YO2RZbWpAZ1JwL8pW7+Az84iX5R8PxqYyhQ6lGPBB0h0E/0LGNAsdAE7yDNiUIeL
YNiIzXaCEMLt5QcGAh28kupumug9cFTSoVlcsnj1xkclrOBB8TKCHFRJklQ91b8k
02ZjYilXJ8JVtqBMJgGiDchdnoGBin2dQ7rFvArNHiDr6NFqYapUQsnIlfiid/iG
FvyiX25W4P2Y0aOjIOtElg88UX0swNf0dUykmjz3pwpE7YYQlA5LKqg7hgu4JrXy
70W41xH7hoauVcpo/CrPJlVrzBmwTx0Xk612PUMybIRHGh6H+w9gZ9Icsxw+j9VH
UPI95uTocLGYm1DEcbC6p+ebh1DqHxb7Ktsgx50RS6MuvjaomAmgmUQsmTyV+fLn
ym315tiL1RK3A9rn03ASffeZEArbg9819Pq9P7em4swLejSWO+00MfiYLe3uWPnO
kIdgvO3I+XEfMUZLGv6JQLBmKKsXlDvY6sJcToewSb0IO6Bhe81g0Trv02JYYMeQ
qRhgh/nfain2LaD7SiAS+8tmi8yMx4GCH7ibA0FExx5j8OOcPPHdj4zhsRCKG5Sb
sPNOoyucUczgTR5YQjO228YmyV498dYrTFwYlqffVokYiPjDS2SxEweSFVasMpzP
jzBobFRyEgxT1aCj25p5NG2VdMuw9MjablWiVG3LfxDUAwfxKCAqJppd3jzjYx8l
uR8FVL9z2YtVvRSnhKYqLeAZtXeq2N1CtldNumwaUvkiZINGEZsdeg4HlUZDwADu
awtkIgbs0mJnSG5MzwrZm+90zbe4X0Qa1zZk2ut2DmPQpWxO5mdfM2wu+KUr4+8G
lUS/z/2tIN7hRqroHx4jvYOUeIJuR+60rZS7SRaP4fJFYvHgQW/cmnE4nsWBgiRM
4glR3nIkrmsS96tvFgijFsPZba4hoGjrIfcVGMKgEqkN4qAyXgdxRLL+TE/rCmtt
lZE7yYNogvxiwu7h05tSRFNHYobVFNHFYNmx6Vyd5g0WjKANB+Av/RUGMZ02/Cg+
bsjurhh5KvgzHl7gsFndtwCQdGN8bDnObiJVcpPVhd7M5oOSXWpD3x+8MxILGiO7
2xjnVEBItP/MZeneFfZYKebSH7FHJjTvjjzGvKliGfW3MAVCjSifT2GOUrq/Cpps
sm7dPK/3PyrA+Aa+iHhug6iLKwsia25U8mCucfbAkZJe1BG1P0khuo3WzI5FNX1V
BFfu3Yg8EhFJza9xUhv90AjYRowxFhqNExYZAeq1/LwarpAWPiYLQ1PAD2skPbnC
bb1B5pG9yz/jbB+/I6EQGhMAT0mB6kErGFnbsXGo0Cwaipcyw9fE/DL1uCsTue7c
VFYXI48FLBrkvIOOTalwIQjQRy1nmBsmIjIFdyGqihdNJt95FLRvP/Xeh92+gbSM
/7IWsK2kSr4cNNbO9tnwX94OOAfAIpsFd7nBIqfRUD7/GNblGVg3Kxp5fCD6bfNb
kVfeicv754LLFkTlExRONuxVGBpcLsdkf1Uja8MNymUkmMBAPCRZucfcqJ28kFFo
gBF1Hp/Hvx9zMW5SImp79okvUFPABMo/2hDdFs09eYtUoqHP1fvh9LU/BlD2Ngue
68co5GTBaVZjKY1yNR9ZF92mQiTRevwyKbqSNoolkBUqb83ChZO1UC7wwlHjhf6z
XepptJb9YSWFZS9bgD3Nfnvbx45jGm7P6R1GBXUuXR91IK4D3sB2BbPR5bDj1z8I
+51OEwKgrQqCZf7riRGkpfwoM2nuIHCsdyFy/X4cGReRhsd5HvTcq2AB+J+iv2LI
hcUYYUabYXX1i+PbWUOTb6rkaxzaKJTbgaR0/Jvw/AqivsAxGZBQs4y1VPzKyyZL
1ENUJ3drRMD40ByriWz9MH8lIeMMOldr9/RJgurSz2LSDudyHvNMNjV5sWigQI77
qk82SMuF0wLutO7PaLLsI/4vxmJw5vNJoIOLP250WyGvBledxpu7idbToG2vOhSv
bQPd/qjj96AED5tcROY5bghkSp3SXpaAVtb1KayaSM5TXIUMoXMqR0XMHPdcXTzT
MnkCYzcFJlUQVZ92+OndD2J/uUjokskHiYrTmrKKDnmGsWK1c5G797TiGctYTKaZ
/7zCkgsPbfDRfxq4Ss2GsCqKwdQPoA8+ExcWfiTWJgz8dk/W8BsfSYr8ruzgJJfE
Io0iFHnxhuPqN0CYwVyfj7zWa//gfQktIZHnesVK7FNFz4A2XQnSwksFeWakzHOh
Bw9mZqqPWTHfy4Hjj8PU4sPykFgpx9ATC/DwAzU+ErrpjGu2GaFKglmpeN4DsZUQ
V3RoWbVivfBP3J8sV+oRGHfp/p380W/Dj7s1/PzDsXbvih05CNSPfYaZ5gtGFMLy
+L901gO0KoZuyhI8judR0Z1WtlgF8e3vrUeC5MGD4sCa6ktEq6yH42QwCvDCmYMf
gVVAPOmJnFE9dCKKxl85c6zOpEGVUnJ+u4DlI9t/BoZlLWP1p7EZHpLtZhnTyUnY
CN/C0844lkNqqFHLrvulSFzJDmrpLekbSQiiwZyuSbM2YF4NymDxD5dwwNBx3njB
FvmQTFPwjOe0pFFuxmC+UqxgMSVxstJ47cKb0Mr1itzswfsgqUOPzVC+KuiH+Ybs
T+ZlKcc0be0KRXLwWPW1dZrP+F5dEhMNfYI0sf3IZ2jq1IraGfNbOEIgiJZx1Zfy
oAPhsmTKDKL35DPD1vgx1xRrduTcraCK5utqrrJOTiN4naLNwl57SitN4YIx+id7
7xwfAOjvMlo2rgTB6U+I3i4r6t+cV0O/3iI3UEzqA/I7Zq/M9j1sm90EM1V0Sq2I
9LI9L3WVtJ9kcr9xrchGKIrgVxcCNxHVXa5cCNwZzHn4em0/DLm/MKV1BvWVxdXI
uHH+OUpCXi0GXHLj7svnUldlGuoiChWE34em/jKbg7wi/4bWeppBQdJxsKUtiDlN
WR3GmPL84eLvJSX8OY5L5nF/hziQHFFudcTqA8mCOQ0EHnKxNxGUAqpnLdZ9/R19
Vrc6B1kDPkn9XGmr9A7Osky5YQvV2CuMlAzccilrp6owK2gfEIpV3z51JDJcp2H6
6MeGxoI7e5JFAfO3sLANN1DvORmhuzD5UHXiVTCIN2tTtg24xEMDrkxjEUTk7Ccr
tvBvP/ErNAN9hPJfVtknBmmB77HK21dcaAcFEEQvDUn5uQdZutnfbk4xlYlowNXn
n8JVGmPnAN7Ely23B6apwRRQm1YvxEthrRqc8giaNY9O4FYt7oYGiCYFcaT7yBRR
lWDZ6W88xP1mNkOwrSs9WODrc/mTr1cDP829cuuauXidJaz5/l2Go9P1MD+jKkGb
CSaxESEqlyRjW2YxkXGCGs0tdCnEFIObGpzPaJ4aPcWXlh0+CwwGAN7rpiW0jak2
4XgzVzcJoTw9DYQm4PHSU1dznE0lr/smNVdlSCCd4X6R92NxRL9fLXiErdF5iRT8
stXFn5XrKNhd+goSoL3lDnVwdah13pUzU1yTKqIR1LBiq0EHRAJTp79IMbEF0zKC
Hjdf2EP1gUqXmpgZMcXCpSqXb7hqChZgXR0So9AUmNdCL98nKDMwY6pozjygoUy0
2X/MPpSS9va5ndQZILDgluKhLG3JWBTS/FXsrKEfV9awi+nXU4Tvlq5qTFlhDULE
ObB/t2boJJLEhqF6hELJPBjkU9gt7pUk/1SXVeiBJqiC/sX0K2mYreZ9CUAkOKVx
ZnwpWziuR9GHHsu/RgxSTBRyw77rLmFTp3ONLv62QFLD5FFiT6uaMeo36IlJg1gz
P0RAfmsnO9HkgXWJL4I1/FxnEtWHuo08cf7Jc7rluqpZ1DZYDjaOI+MwIG8Y/Do/
FCGVp8JOWhqw3VuvcIprqQJvcph95ojMde6J+IXbB51rPntMCL9vUxSddcP3Xztu
upheXnqNAIdhpy6jsIaVwEwaC594zeG7n9ZY+92CfDtzRGi/Q6F4AghXaRnslWt4
8+6OJAM8wfeodWcKGO7zPCD4q0nJRg1qiHEDXDQcWFFX8FptjHxZMdYOMfm8Jr3S
pcFKRARrXxx6DGzYOlPab+3mxvR4zLsYOlxCS9TT/4vvRhKbAqaGPqYccSPhCnLB
DxGjXeD2zeQwgOkOKGlGLijXzctIfzT1nm7ZVhpu2wHjr1XbqxosECxb/Kb5yVoc
WuN1aBv2mVHpjGXtTZ6ZXfCyyn2tP/alldeU2fSPG2RFAawOoCyKeEaAAgfyRdJF
ZWiRVISFSJ9hi1j+cCgNO2idKRkmZtnzVBH+akBHtZ2QXH9G8W5HTlxOffj9VURg
PfGuWPVFtJnGOgEgM78JuY2b5C8j5hJcBz2fC1Xcd/SlHlKPtHFfsg6ipEQjT+0a
EPsFgGeK9qaLJVsZ9IipEn+selc9wbj3XyXXHwgk4x0M4DZrZZlpZ70vvEzFCsMu
79MMlgsQai0/HypHmQJhXc2/NrRob99LPSecMPQop+Gq+WzZBGul3FHfZGM+hinC
rkA1e7F0fxeg+tongi0mvcwWZbBefsB/1m9gX/L3Jj1zfTq1FnIgFCTPNjTG+UH/
rMuEf4pa52AE1nFU3w9+NzGb01AwTpdm819cBK6wDNGajjkQZYHExBsWkNk1Eky9
8Wwh5dHhYoBzxnd5z1wgXQC6159vFPKBlquwZMPvuWb4UJt9w/QSkvkZBUn1B/Wf
G187qO3w2Qlr2wKR70DK9eN/IxrR0qUWzqNj0G4Jnh207WYPxySV1eM2Fq8MAnPQ
GmoQrsxIHH5LG7xKRw5sC9XV21NIk2RqJPxKFPHtUNvhQJBc2uk6rlq2gZkuwHHo
wGnTcDtiDTKOc56ogfXDvNKtDDNAxTDNJm+y1k40ViOtcnu328e8vRjP5wLdGsAC
6FAPvqN0di+dsVdHeF6lurm8OeZK1KcrWvi9m+CHc0eenVrzAn3QngedOpU7nqBN
IKlhp1ev1edT0H182NsU2QHNGw1SmZeplEfWjFTu7u8AvXPfIMGurMEp3i5wXwFt
bIhaPCXiWJGjHIKmXfs2EEGqoNo0eOA8F+CSLwOUNB4kH0pbHG2WoqINZ3z6GSYg
eCI4g2XdcgalymWu5f2GNqWebGf3kXQautF0g0MjeQKqaH9O6wyjmAdwbh4cjO2n
fflizY/ni1Yc2Espr6JtWFc1l7TPDSJR6L4I+ApJmlHjZeSG3zReqBKzTLgRytSx
ZMq4xkqtn4KjV+7b2uqqWT55lqOIV8SDre6IMpAVd4BjHWvxlRz7B/gBox64IecJ
Pq+K67olLuksgWy8PuVbKH/HavVUomHtp7nBiN2nKTnk6jQBAYNihftVWW1iEISn
GYF4bWJQPGkqJaH5nUXaZwxjZD7bgg91Rsfa79p6PaE/bfCy6Za76fKZJ4tPwoAt
AsJbz+Ud23AlJ1VRnWXGQQH5HFJ5rOblngOvipx38UOgxUA1+gA2s7Q8W9RW9c4K
Km096hzUy3qoVDaUbXHaCVMRl5bWx03yqg3CeOmB8dP06t2zLhiQHZHzDN5IXoOE
5js2czOkNCFTuF8TBfKE7po/Rieq6PMP3UhaoKRkSTsKTF25CihlIYE991nn6KrG
6iSoF/fuUoaJiSl611ua2zphFHFv8cuqNA/igzuClM4vHZaovPZ9wk+XkSHN7fTw
wsAXCB6OcD69VW76nomWELqMqX2IJfUCHzLTQMZPXMlsBiMn6UnNWlkVpU4gWgd9
Qqcysc6A/T284VAa3N0/U2IeNv2l9xjeTUOBKv7ovYika635Vu6z3RYHCB600ReT
AoZe5bpDaedyEtt54S/F38nxMMYwcBA4DXruYGHoquVVj2TkBNrYeIYWcDICzEd4
NBocxA+htlrl43kpV1pL9amsBuE46lTjFQUMPwbw8YNibG1ZQa+/imWPobB6VUV2
gm9B/ttuERz7Utfg5E/HZAtZt6cdlKJ1xuuqK74U2RFn1+Lodm0NxvXGPFpyG0lU
zpQvgUtnFXyDBVnwUiQQ8cmlmmNEyNbaOaaYZO9StPbPMmGZxPzOltjVLKmo2GoO
zVlFPXyibvDNhJsmp0IQrRIFzFUEh+jEWb12BPpeYuL0XZqG68t7Pn0KEhF7uX+z
ti2wt/dEOMZDDKBSFFdW7EYJ8+fuirjtlWIIpQzocS33XdOjV/0FEARtbdr/Rmeg
STKyfsN8GogUw32bKlaWlPkhyfHKQyYbXxVU/9Qop6RHYc4pWe0xVJgc/z1P+d7p
VzODTHqZ6KgKOe1eGceP/D6pseJR944lbU0IkhaCFLc/val0zOKqNZDZL//dfOct
/YIoLjL/m+lJ3ADmHanvspkneqeN7XYEFnq56Z+u529uincYYDizcPJ6b4J7dn+v
p8elb50oCUyef1oVDpB7QHucCwiDI0uyirfPKC/Br/IGg92hvmFqmTdu3PU0un1k
AHL9tXZ/frkzMuqdYQTixNyHGvEC+Zpeo4PiVMwnLZExmYBgIvKCzAuTWdXIMsHW
tK/N/E9SNvtc5XhkBX8jvxYiVqPghQT+z+fHUiiulBq59PLVWQRN45bgS5KvaFtt
d6wLXh9tp9VDpnTDSPIbJFeBFzLExzjJRsY+lv1OGowix2YS/N2I+/KApRDTiT1d
bPcx5kTwecLIgUSDZGxTwEIqUWESIOaQl3v6XEl49ITSxi4npjZd5cqHPrZMLRac
Kbc5Vp7cL1dRRSeUrOKK/tgaZlWC2H91S+WLrPk6bl7X/VQkqzycIOEp2WMYVH7X
DiHnJjgvhuHBxXnW3q7NnujaocLsFPVSeyKfylg315iXttm3ykhYC6zlvY8mTdQd
oXSTrpjBVpirmnpoSkeuAvaYTXI840TpZVmS8KcnpgDyxI3f7UEje0U+VfRTBTBo
MkZykdGHXVP8RuA+r3vqytoA4gU6zf6zXnLaElqp7px1QC3mhx4dKak5z0KLUX4a
VMzAh91U3CHhNFlG1napgttQ4xyIPF7+zeaIt/gIhm+kWwBj2og5kVkt10iUCfpL
EgkFs9uZ5F3MHcq/Fo+fOVbhVTiQtPDcrMXXQKCC5toG6kGM57+8F7oI8vsB5LHp
VRJieFCWgnW0hSV++Bi1OC48btSjvwcxoAth6D4WTX9ge5wKte62qFI0smvay1dv
DCI+1ZIyvLy0vob18YHfWtR7ZrN7PstAHUFvr9ZdoBuln+HkLMfr4b/OFRPQRvXw
IlptoiErOgst2u74yGqQVU5q0QjHOH56xt87C08absfLyGmtyTs7jNbIVfDRk7rT
VAhGyD/2YtE3sbLT63l/1ot8bwF9mDHrsLS91nTDOXKzi2/4ErHYfpLPWIIrPnuH
m+p21Vy63jziJF853VNTX36BnndhrrVNzT/t7fGA/5Nk9UYL7tg5Qw9JGMJyssn2
uEb3SB4Wad1hHd9ok/pb062LqtBEvpcLIx2OVPct/udYJKqCsf7H4zVXilhkBJ//
ntrpr4pSxkWh9sOng/ZuZ1qD7IINK6MZed6IDz6YhLTzUKFgRn+YnCnHiw3522/A
XySViY0p3OR2NcAZa+S59z8qjeeEKg5FK2/EiROXSUqVBho0TCofWwM09pR7zUXG
dgDRE7AO1T6E2qE/WFs0MLfEbaXbJ4LoXSZRfThKvkmXdUVGY+jtv4TVD8ly5Goo
w47fXi2yp8ksPbdlnj7muEXAauNm+CkAy1SyAiiymNUe7Hu3QfgdRUtAQv4ofK2k
BbxFOLHMaxRkd3DMI0O/VbLxQerz1x4TjIf6TbjjFrvqxHVA8hvWHQMDdelGoQcZ
ldfE64s0oad7Jdn+X2+u8xP3vhx4kUcbtvvkg9L7ud84qNlJPQvVsxsTeiajrNin
D3vSooAxkHvXMP9I7whVUJ68fUJA354Xsktdet+TfeoT6exnj7wr6EKcSqAIYazQ
e+U45LWENXg5JylTWCumzmcrF1JQR8lbFOm/VooZED2aDgc2Exye6dGq5IdsNyIH
yo6i5NR0Q/MCzIZXJ3Ulc+Xcxy8U8IKvIebfIXiOc1PaccQhSFUDKvNgj88E+nAW
hMkjoBBaI/QBqw1/MrOZaVn8A0i/pxpc25YBXybYTMO5AvIA2Lt24iGiASm4VL2z
06YgNT22N8SogKqE4mZf72KTiaPCG3F1KV3vPzsVFByvEq76oQO8jv+dMZVjbCdz
Je16eNN7QPJ8oAacxlzt167LcLhx+UDUgYgp6Bfqd2F71q1aLi6A2A2PZX+W5aD7
2+7PUQ23XhDuEGyQN+hgnCB/NcWzYa8xh+B8P528zqNUk10bzfo6FK7/Q2f9ZUy6
qcuKygDCxhkX2/mKTAHYkgdac88Rr0Lj9lyGryXixK2DPbqkXD1a4vyYYRMpwu8L
u+juK1xOjwrSp75QuA8AQ9uWk2WzBj90qUKwWmh4PG1GKJuCjo4w6hCYRFGlPcj6
u4VGss8f+CvwjTJQkWx5bq8X2AZS730dWfZJZYdJAAqaZexCZKCXkkilSLIGnFUr
LzsIKT2yseDMjQcrhaqmBv2oUQDpvAHhhGeaXs74lTZGlDNDL3atolWKOO76rlWq
HgXyvXOzdmFSCG1AyVOC05oEpYcuBQeqOatCj/ujI36aVCx9kvzPQZMEdu8HlqIA
aWzAKH5nY38+kf3KlXlBM86Ho+RlONVd4xHaVtgRnk4un1KuuTS9Ds+KLj9UMFPn
R87I11ps0I5IpYIbiUmFwP6mk+DQ7V8DiS1J87v1Ab3HHYE0DwkEkTciCQSp02gQ
v9vs0Xf9wcjQztPKHjt0Hvcy8DMZx7qWAZrGRds9eZrm/sB6f/jX81MNb+uWbLWy
0n4lxMwjwlHuBXwpI50gPAgBcDxawWworUaeXgo29pEH0MP5Uvi19kNx5AkLAHDy
jCzQtfS6m/tH2q11hVyDk8rKJzhfx8xEj0dcEUv3/SxNR4K/MFAEBTPgBlCzZhue
7Uf0gbaQvwPxXEG0JDgC6lsh345VsD8cvF4Krys0W/bw5QKDCAZjF9ev1aM5iVee
WDIar7d4TaRFAYALx+0TvjUb33KyP8mWgOGplUR7LRUpKQushWos/pvX0DpeygHf
RruS1ijqAZ8xIwNlMfISHvQXlU5RXncsQZR1vSfNP0jr7duN9Y1dZkBKo2mmLmN0
dP57/PzNqtQsW7uPY+syyd0AaUhJdzJT0wLVeOk6fmT9IqQ2L4uYn2y7KY3zgpxY
EpZOgnjg7dO3AgttxMYyPA4MRD2Mx99bMfjKALiwzvAQuXXnr0KX75nl+JRfGhmW
kf0iPMevCkycu83VTh4CBLFqpg5g8DjW3A60OpyPkxEM2Xu2VLJzi48uF9XvMAqL
MaXKztmsZDLsdfrbt8S/LdIp5vscr6S4sKalojzrZcjD+ffvy0UC7tckmX++lbhu
CWL1x9zg0UAUdk3yz3CA32hMb8pG0DFDMpDuRR/R+wnX4kL6HFXFWVZqAhJf8sL4
u1FY60JAVsu5URk8jpFafMqi8KoQ/jcgVdoJEEm8Z+3VYRG80K4Z42xLsm6CFa80
AaxpJ0vRSzC6fAS87Rb31EJQ9E/NkCtuPD0MBAEEZ6O93rhddcIdu5AIcTEo6Wxc
26lvcSEzM6G1S2egcstckEFPQeosMONtYGyeL0Q64DL4jhEx2bYrSZtks5VdTL9F
aisL1GdEfnKyPOzkxWAYe8pdHDNDFoTl+SeWIiSXhwSaCT/+MvCwa3TV7Y5bzsZs
z4y8n/xBHOARE0Rc4WzdVgZzxygxfI2He2mLirGBfOp5UuBtOdnghQQPH5PIux+W
G88G4n0bVsOAsphH1I4doy8m+hY6EOWLuaBO30xN1eiEsVfMECbKPbl5zAuIDQn1
lVIyC2dK/K30SSKOo2vlooKibxdHrdNwAW+76LkpRTrS7qeLqFmB2JcA6Rjb/8Ke
MIKc47ppjcg6jYH//d9IVGo497XgVHZseiPKBdn1Ni/Anp3Dtcyd4uB9Jt7hsTRQ
sEZ0Ay0VHTnjvr9HJwItkLEoMkM3oGnrX4nsUVenrfapi1tktXbFjlCAF/GE6JLr
rxY3AmiqXRr5BZC0kcyCGeQ0zvIrgwa1Mzer5IbLwHRFH+btLhotKaXZjV0bALXt
omdrOp4Dx62cE+yDGvd1JXC7WlG18kRgVI5osErJDkWj1WAhCHW4rSxueO3/+1mP
8e9Mlwk+JwfzhECS798E6BTEhjHzh6ZgtKkdBVONFfOD9NzhsQa/jPgq63Bvve7b
LITHeajJxsP9yQEXELCytltwc/wNrXJkljhmQVX7349P+ZocfVdEq6kvAJ7c4XFk
qb8kpUu/itmsF0BrtUEqzmaSVk7yGRXYtk/+kXq5dk3n/k3o6au2Hugkjqb/Rywg
L7bUArchn10WnTq/g3eA9AZJEScweEd2UzWN7GhhG4J+9T83e5sThB45KhOXzYeq
plF/Tr+28n9VTuNShnOVCuueAVWC1gKuewkQZNd/f3SkgfkdS1k21v0d0PNghTHS
7nS9P1FymBKuBGDIRc1lqu5b8NJD9Pk9GP2clY5jyGuTw1HBHKnhi4trTevqJFxz
T4yrxAtJ8za2x8SElBF5pqshddUDaIhEoe/tAnN/d6+I6UV9Qe+GgGKbumcepka5
Xj9RJzoYjWTssJx1vpq64BZv7S5gEIlUOnmIMr24RpEOKyR3MVs2n09NREgia2Yz
baYlcTxaZWFJy1QnZbpSNmpRLC2PrsMykbtIfTjE6l+/BHRzG23iMFOpMCcFp9nA
JbljK6Iz0Je77V2HiC2BKD25oyR32fHO00gDdYrUVw+/xKYqw96SF23ej8ggE1SB
qKgbK0jQGCOd94MXWWpA9YHrJFEXMbcC2WU/TDI3W+L3+E6xj2+jSe+u56TCCu1d
5Z86sBZ7599ZVMZZ/KNAbXTD2vzwmiitqW7+SrgviKZ5bZMsY5rAKrNkVzzlbA4X
PprF6n18rCoPMlAHKoKNdqh2a0zUTzuhzgPkVil9K8B97xFnCCK9qsMH2LEo3nLB
HWQr8R8K6dj6t8ISHwUe6JMgpOzy52ZcSctwOeZTcwtdwk+8v5iUmxup/j4iwVRE
DbyfP9FedJ39xl/S1xBRXUU+KAPVHxsDaPGgt8uNR4VDGt0WXAR+tvqmXHqAZLmX
f5q+BMORO1BMBT2oakDq5FZbxImlZ6NZr6JLqXaxtuD0eD44GADl/Bo2VeqcSs/+
EHiR/98C+61U/F/Tn+ZNvVgS7Ro1SbTZWkD2tcTOfrtUvyNfnKVlBUwcp+rZ0RsI
op7PA+RDie83nPlremIS3hG5eHbFqpmn7ERxmyeJlI0DxHQ01/1WOvewm98yaNyO
0N87pMPBMLCL0gaahTrwnQuvi11Q9MtKE9KDm5uPtHPJWZIAU0FE9R1gRodrbWJQ
7ZVtH8t91HJES6WU6IGRsOkozc2BA7gyjTKfuc9ruDqXQTzc9YAdVuYqH//msgTm
yzEb7+zbLhCC+fmiGolSJ5kvjfRv+yZ7Rw92PRItEYemnHflbCqmj1T4hNAzfA5n
WZ+W+9D9sI2Zm06ENgs4baG8bTn2ZSj/y4gnVqWQIn7L+y0n+OOtiEw9+3FQW008
HP0MKKy5crjgrzvOYrvC1m8Zd1z8Gx6SlOTUF+0WzU0FS+5SYRUvdtXMh+spnaa/
XTuFYuEyDf7c+XTqMDbYuy6bWp9JFhfoMToEjXoEIeOzic7N2YsxMFaP+Kg4x4EL
ok9duaHC10e7CyWTYShISUDOlKLLxDnqpRJahlc3T8Lb7azZCbDqs59+FltQo8hz
f7ngfCY388udag2mQzop9qtBXfQbAkL9a1MnusHbqivjqFy8oPVvvouFFkcoB8kM
OjwRAzqX7H55rxLFCx1wtNJP5xGNB/ZV2rfDEdtQZQ5yU9NFenenK9oDZZJ+QagO
vj5yvDzWIrAVgKMGEuNK3FP1RjHABj2EP4RD/ltnTzg+8lVayDt7oBdPO/a9WnDC
VHkV7gMA3WXuGaZZrePqx526FRnXQX7dyz7AhwN8iE5bUOjAq0x7w3lVGQ5aqs+d
hf4DGqYPtm5kUupxpNWO3IKYeiSamq3t5gGPyRkOIStHRjsjDyQdvuVVndxHGmjP
eI0eXGYjgzoGceWi+0AnmQaZvGPT8ozemx+5qyra8O9L46H4N/0IWLZuHQCqhnUa
NcQS47eZFh3831o7aNTrw2cZVtv8Qma7j2+C3oZaE6n9SmU6zy9hTE+cmXnIe2Ga
llQrjcbmXzzS0KvXjrmsCYdUeRSMToPoW6EgrtogfNulU6WIpq3Xfhgq0watWcyD
a1I5+pfoJReYSn/uMIWI81sujblC9mp0xkLZjfQmsblAPAaXpRvPs7P9KaevEYY6
CAuK2PbwrjDeyfU/G9R8Mbb7RkJLe/lhBaygcb6zLWLs9Bm/ZTb/YgJnyAvx95sy
1Bx4TYxz+IQXNP/5H037/d9Do8ch+ZwupJvRmsH5unqfaaHbX3u7rQ0F5npt/Xrx
ilH5lKLOtNvlK8Ji7f5P4+tW6nxsLbDpEt7/Ahqlfy239MRta99lpL0Da4SydVNQ
VRKR6h7TMHQpAhSuJLkBlxWncJ74m8U+A9SWl6XsFamIJt9BZdmTvahGsbg4e7Pc
kMDmXmfuGVVSvOFlSBu47JgO7/6YXfYtLpUrpQUBlO0vD6rfcb+PEUj1RcHk9BYG
LauIkaBxTMjY8w37BX5axpD/t3OaOV5P2c0yc1iznvaYb36pGSuUj88tf754Cj/7
ZiExT8U22CsDnUo8XtoJZchommCXXi0KwqhB43pZ13SSMlyJwMQm2bL3LCOKDWwj
3I26v1c4rWz78ohl9o5QgNWqFDnhUQI5deoswXnAR/ZiLU9FyycDORG3JTekn4VC
Jm92ivSI+r6YM1W5uGhJ9FANzYbwFcVwMmC+1EXCErTZ2B5wKPpBDPFYL/Qo8b+l
r8+wMBv93xnk4JN5BIsugrp6QHc+e6aS1QCGukE35byiIU9pmQ77W3fJcqvNu9Rz
xnkvS79XJxdxCXKV3ICUn+A4+33T5Im0L41xB8Ej9cVaKSr22uEQeL7UnLj+fHW5
/eGwny4acRzGZAWUX68N/GSmyEVIMDMcTjKATOhNlHKzCVW5hp4zA+JCalX+Ndkp
lp/asRr3496E0xJJYHZc+Il0p8oypy3gyUc6kaLtSi8hE8q/pWwkz7tTDkER93qw
AkG8st/SydozDEdr0Ral8Zj+jBHd7xQT9k14cKRb8QO+XWmeRXsZbVWj+zrXPq9Y
td1f+aLZewzLTK2kp0yRq8/P8dE6liESOux5U2ZgE1ZFtJPxcO5Us/v/lyu3VLVk
0ss4EzNH9UdLOIgr1WvNXEaqf7XseSPdDxRv2Ooj4rrRe7EZRrk0BkLGkLIh/RWp
X+UWaEZ6ErX552Own2jGEpt0MbD7FAtapluAcRY+pS255SU3vJGknppLsYTvLIR8
rt1TD8/71GnfplHAWzoxdqKXJYMTqbPfo0nOxYt8PIUY2s8lfxIorI7eIKXIMJib
eDA+HYM+8f5/4kwV8P4IOrIFQMEmou+tMSPH7d2qb7uBY92Mh3BjNnCc0n6V8Hwh
1g8KdNpXRZDDl/RdLw4Jy0D5EyYgd+ESGM1pwJd4tlSjZRZcWee9EpFD/A9xP2hs
Ns1IIyWnkwniBdwdasOBUWRLNWZ/DqCHTneg46NGSFOJf1IgjtmYwR4Tm8nzaPT0
Q9HPyJEFx3dG8Gtu//gvLXWKTTNufqX077V9L5jwXz11yFuuD4otJworGjCi48+e
o5bFwABz1YE7DD4ShxAW/0PcefXYAwkmr9txv4xlgdjquOQWbV8iz2WOMfCJGsSj
8xUVDUT2jOAxHbZM55iGVx5xSDwVWvg+J0A1WYdcz02FzBN3XaSkf0CYGOKzfgUH
U8EkEgAM5z3OCHqveonKhDOJ3LtJY2h+qfef3HAvUAubZyi7t+nJKQAIxRpifXDK
LoJqCG1Xb7bMwM4Zs4FHTgJXR8rQQOK5Qvj7Xc8LrXBtrz9I0J3WUYin6HGB0k5h
Dh+VeP2Ix0cF8V8oJj838xEBBWozQxpPNDydddCj94ZTeyUY1OIb6jIf4GiMv/oO
L5r6Li5XGMSYfJ4opu1xCvwXy9nbyaRpINAt5PuAmC3rTfWW4EGz3VvzNR0eDMSC
tJ4Sp5spbSB57RLI5prBTsWfzUvy67e6/0DL/k5XYVNoFMDGMEijMmJ1w7vQn7BC
ZgVm/hxaus/jZflp6C8Ej36Jb5ZWMm3UdZASMpx6WNxN8kZOck8Kvj2FT6GFm/Bd
yetUQCKi887G5904RsvIk1cINTwOE/dTNfl11l2QFMOk2hcqjOSI01nu5RX7aB8z
jbARiHwPFPXR5pw+hI5px/FO3s36BiH973QRibf6BFyklolUJY7hpjVCYUrX7fqd
Qsqqe3sZT9F8G2NsCMnPVwo392sH2U1MZkIlNZAJ3QvZwaKcRqBhUkopwqQjE1cq
z+O9zFamqU7/a2RGCOU+iec2x7yr9A+lLAYIuFm6RJIp1eWJp1u/4hFyUut+5SOF
LU/7aevLwPEbSO1Mm8WDiVPwhgH72/FV6ZdIFoDWevBxaTO49VXoaacKXDRJmbBK
FswDqJYaiTNZ1aQ5IP2uT39mEYBqxjwWfzkIogjbt2tuDjYHlTGs536NL4R6oEQn
h0hwf0WMl+2PDnTBZ+QRbgqaRntTMUAoweAvXNV6klvmUkqIavHhe9oGlSDq/cs6
VCHyPgwLp50ZpO23KyUF6+dIrdIqkMHTqWyNPwNh6cwividQzC7i9m5HmuPkK4ET
b5y/X+2QBUc15S1LLckbw+H+6ms+G/ZiJGeSv2lVAHLWkf/ubMDxkJD05dhDxwpl
tLYBSYy9eM57KRT5b6wDsHspenNyzmmgc1I4XiOJE4qsNMRGxsQncaLaCD0hcH8G
HsP+eT8+FAmkwuCu9K18Kd0V0j1YN6R704cuLhYFIzfH3oWYSjndPnXFvO2u7JFD
oJQVLF5xegBzpxhmmC8eQ9SZFuy4ycFQHW0mnJ+B6NqgqqMnJuP981lstJ1hnXBA
Zffcu8TEOsq+ZlELo1Qbvox7Ut7981RuVGH8/dC97TEzSikvclxzG45KP2SFF7yT
bzXln1rFho8yAjGzpxVIAPSmPyhPv+iBQEvYBF+ysMhHzqITCxj/z++A6i4pOiZu
tSJfI4qt4aZk9JTBk34Jv7CjkvMYhBu+fZKmNX0kUg2PD6pP3+Wp30CxYyTGFLBQ
i9kC1KU7ELI1P4CkwRl9E6bVmyn9SWbEsprjW5hI9bYzTA8DFRYBefk4Kk7Se0un
2SIHUKJ4nLyNC2ni0c3KBdUAVDRRerW33//TkbHfIcQv2gtJ8BUPralVCYquJFBN
9WOUUvqT2WbjGV0xEcwBA1iuA/aAl6Od23oHSE+5BqmT5gt1HGhE4pvTGL6HZahu
iL40Khx7ijFckuzw0g42mmSszMdqtmHlYUSUwwu8Q/0r1gs6s8Zfi6XfeTlyULR4
beaoYOqNskZWVKF7Ufrz9twR+GFUJXDaZsSfC/es6I3CLxmT6UVR0LRMRXhnx2SZ
zKYjJm1akSc9ogF9uwZOW4E8PtF/5IOAvr2n8kG8RmcxhXzk/aEF0f7mnnmlehXq
4/rT0lvEFv6/xft3J6cBsTIlJgF+mGmlKe5rbOjuNhl6TWTemjIR5KCNbWAYO5z5
wZ5BY5Alz0XymW4bNG1XOMGDHQ0CYhXCiupnLUo5zzXNCTqiY5QBDoX+NFF74kB+
MELwvr3KLJCVWsfjH3IPR1zcuBotTI9wSRjRFBxpH9lumZpXIjLJ4VRTn/gaLiTa
1SAJrDiQwsf5i//gkvxFUMQRFL6uvcki3UJylYG1x5/xb+4RhKxALoasFriMNxx2
cYRcIoKnPAQ3ByMhtz1dEo/qDeghKnrzSAM5wWXR4EsVfmE80UduHIErkkjh+Aqj
L1hoLhYbY2M2aBKqfn3ldABF9exvtDxv5sKzITr0CJPr/qckCoWosDnXRhvs63Uz
ptKEyvlyUhdRa5yO0sc2Ry84OYMqKsjHxpMeZy39V+ksglYqga/zShm4sDlFqV2v
SDHvusJremKQC/rPYNy+I6EbkjUjuSPqITJ4w+/kiJp/jcPwUAmmv5C8zm+cr4CJ
gl0Wg6eAkPZ/G0CqrxGExPPOcCfDn/ut/ZZM2NIPkG0ksvjDyc2vwHQ4t8Bt35BS
BlZecBkKhheKOVKBFt5Q8j7kdnbzvzuC1lXexWNnoJ7zcg/IIkcyrKGVtE3SRZ4A
BRhEauiYj9QmCrzutiY7Xf4rl9abH4zSMYiE8Refh2hIfKyLrXiX/gdsZNxTRaCz
jhv/uN8bVSSwFO0FzhtqKkZ2CymSlQU7Cl1tNfvRUES/TB6+yw3XI0Q4ohJZ7Afr
F4WL+4qDaTJTdQAoCHwleM0ndawUW9EtFIn1eHnDaZ5/SsvegFA+ldLhSNxjGZvX
emQLjg5JaBWdW64hCebk+vJGCchpl9o6mHKlmbjs1RL6wFQgtlN2rrC2sSFpoe9v
laN/CM8iZ3OencNUgUg1PRpYYGUJCUyu9lXSVV/lJvZEZfmBooJG+yDtSqRVXzH1
VIbK/CHXaENbHNE4yfTJulpYSXuVtimq2cFosjnp3uzlKYwAK0p4B5Y6LkafbsBi
QruDmJv3JX9St23nPDYRNtrgaMZyZKmck0MFBB9ndolSfoPeGWEhDHBaTavzLmt4
XXimvOde0mKr8pocdQ2U+JGmRKqMKwP3UQ8TND3j5kbLtdfmim81LIsivVwAO7+i
lkQb7y0ni9Bcn5pFO6k5mfgt9l21l3KPUWU9K9/2z65psecdjaWdNaVFmnmiaATZ
IK/Df2FielBVPo6+AEzB0lmi4MrmdX7Za0XTH/dRZRN2TKXT79RfuaXFikKu1DdC
ye6vGMzmAwZmgEcQEmtZERdOmpx30/6HA/pjPJLcSbCAHY3siSaOK3PUZO8S3Ccs
N2HcEF92kmlxDJQ1M8FvQctMDBGmJtxcdMaLRzv7lwJ2UVsNmk3grnPkxc8D+DW9
8TAYqDCXZpQ5ji87NX3HWbFHizmTYJNMQuB1N3u4FAxcnOXzLjlJA6igC3uTdlLX
SpaEdC6XGXoufYo79N/qLp5ZUO5J34iJwilrqRuE+rJ7HzxQuQ8oyFTS9FnqQFKj
iyVxt1jNSiGDB5ibZpRdCFIVy1V6CT/g2GjL7xxh9nGbMRqFHVIpFqI+Xn/F/K1o
ggxF5wO6JTJRT5M3AyiRbtG5/Lt8cIdhFltDRJNnitALrQNx9RFNj/PRsOHqOC2u
P28RKSRW2H1tACQ0uk3Br74BJuiWpzwte760ni/O71FdT0SURycP6T5elHnau22M
L/n1hT0luspEjja1oLdRWpsR9d2lUiFY2K8BArNgmw4q9pkDNtEZF89NLwXDYQgs
eyXAdCNi1OXeBcQRh5jPMkltJ8JxG4Kp2zl98KBosuIr9Oqzh6tXz8uMoLEZ6omP
oLPvMLvoh3s+UK3HCISu9aXhSP3GR6LHACBd25DbEBqnxMVmr5RoiwMIx7u/Uoc0
kvQTlN8cOPoJURP7rQcXvrpGNrLfjh4bS6RDS+6nY55GbBtIgbGYieJQYo0Dckrp
9sm63WLQieOcuFy1TdaqVK8vFFg3XGD/wP/jqU4sjrnQ+37j9Gr0nBo/vrIiy3yD
JjkBRFyC3NUXpAisqrpVi9/GgTVZdij0v4efAAVvy0BsLJ8rMi+YAWNHpMgc4wLu
TN/JvYBgWmTH+gQYFuu5ggcXy96GY7DDmQ8ZKXKjxk4OCZ1TFlck07s0BPESBNu2
5lr0/NBBi0Rq0JWODUd0TxV8YXOjW+JSMIGQpW7dVh5jfsOcl522hP0dsMy2g0MS
bSrSJ0UeOrDdkFdhCzA/3TSX1W78TQdHzHaZCQhv3YhQo2n3GPimpQzOwKD44lEv
ezV7cgfiXkFpuhcGH4ASh/CJAoxsXOafu6kww90gNQlj4wp8iucJuWq1RXVZxura
R2rX7Ku7fz/EaN/IHchzIZCUyZL/TE+wKnbVowdpGH7cFn9D5Pb+1eZdQn1Z2iPL
bfuqiI3RxBBzcMCxrP7jQeF4GFf+9d8bjDGMk/CVWucfe3dDOl2HsiNIjUihbM8n
B8gVJKj6CIgoY8umCAQqsVtUvGqaCxixwFid8AoKeuroBAwYFIb4IvLHKiXO28ig
lNDLINVGA9APGjCKJDfa7Ufy88ERZxmYk9bNca8Fq1mZmhNBlXAgsNQmI2qD4njM
gJ5RiDWE3Uy0gqrUFSNCAiCdGNe1G3IUWL+Ne4oC2y/oP/GgnC8gRCCHJ5GkrnuR
3PXA5j0y1Ywv4FVEIStsTdO764Q8+vy3wBxxpdFN8zC3sHKkb0B64nbJVqkjm3yp
3QHZv/pWcHlL5WmTEZYcpJzG72sf/hUN89YLKx8UWiZp9e30gTL9LVJxAtPcvHZo
xWmjeFER75O6OJHR44r7BbYtFY1R7uamMzsgYnTHIggnjzw62KZPvnkn+9Js/glO
3EdWIJ0B49FA5EmWyBXs0YU7MMheXUAefZwHnyYjy6QCAt6nsL9usUca9ylARVeq
rlRY3CdM/A0e+xiq+wSPqi8cNKb3e6HmYAimgYVnJOOhYedoXou1QXUGmeM/5hWY
omDl3TCm6TVj3gqNzFHFgNqWu00VNRPFQlkxvNwY17rkoJuEGx43ZKmFAclgX9NA
yk6SOxcOWBGnf7MIJ4MUQiSzoeUJuFCiV41bfyIjIf1GhAvne2LKq0j468uub+Sl
TFmHn2P9IfwMwweDD8afTxNw98kIB4CUohWZrw5iF5eVTnyhEZCRrB7SBQxrp++d
BMMIGoZ1KMszukkXmM7Xcg28Lk1E224ChOu1+C2aG9ZaWYxloM1nUgXnaqcoP03A
LxHISHaC00gI+7Qhv5LuQm1pKdmz6unxkAZlH0cHK0/jdWfew0V6sRq3eooFtc8r
QNAXuT+IPw/P4jmCUkBK+D4jcb9j5dCV/Qz8ERgA4uv1gyMUOTOzHS9ex170MdCK
N+Pz85XfnMuNVbRNfbgVVExfztoULfpPuQpzFq7aiUpWURlxDTEKH1F7gFVGCSM0
tKpwMp1PzvAVlhzkuG0uejd0lbvzP0JmtFWRL6t1hpfp8Xu+nFh35bI13CoOnCux
5kpZ3NuzCPKamfPEz8fjcjBda2oafU2rF6w1g0CbnAd25o/qc7xSZeFZKWtuKoFa
n6kEM2kuLlE43om9EVIOggPJDwKNotqtU7k/l3jLnvPq+0rj6T51kJZNtqqH9dnU
v9mPJenkStMEH+N+jrlOlObWfVx5bVSNrFigoi0HUbRHKCCr4hJICm3imtfGYorN
rDMzVWNq6x8ACVHb48WwAaMr3U7C3g3oSdf7QW7ERnpeZItevlYvWmNAWZJmTax5
Znpyq1bQYJpolE3wVY8VIMfAX4EGoBbqWwvMSHzhktN+xdD2+ZLvnIAvlHyRTso8
SxXwyaMm4fxjRybzv9LMgkSaofOyTBSzS4BnOsxCn9SSKYkbTFAsTOpyL5GYWJmT
l9z+TI8ByoTGGb83Lu2BbkXCmk8vITPuRq5EIMJ9bR7ZWT5nmSh1OH5S0IH+PjFD
9W+Gwn+UCngIri+AQbWE2Rgdm+mMq1/4GzPr4vTcqp7RHh6UCvEiuYZGISlUB8SC
Q9LyKPvnQgbw3fkVjDZ0EsQvVLc8wwhjxGnxVdfNl38OGZmv3MOM3hlG1+CrA0hx
trvNuR63KjVBObllLHNAiBEMGOXOEvw1jrElSp6KbiWdTuWIY9RXkNREOVnYmsX0
dMwOsCrj0ngQxpIYr2I0o1xtdSTfYI4yFF8ZYg7NgkhhX5gZGn7FD46ieezCdoQ/
56aIT6Zz0VtI/lXnlbZOs31G/Q8iiIn+xPOXl9rWxX2AjD4ph8tWI83GNRZ0RsCp
rz5Z/grH2B1pr4ebkkfh7bkYeXAEqdCh30OOe9+SnQtIVyXgBs1KpOb3tZe5fpMc
60OgMbSMSxOw5ybLWjRoRjdteOWJmyS8KSUqcl9wCeO+sUWMYUjKfAyxHa2ISsaw
ZfFicNPiBdktdOg4uNv577iv9KBKw6K8wMBujbRRXMfFShsyth6Dktjk6118Jbnn
KFU/y26SdHoi53jGS6LPu17REEr+MwrhFjL5DG1k9J2fBO4Z6gyYSM/vR8lKHzd2
0843KANGbdXRLNCYhkM3spbrDLwOa9Z4EMQjpCfSx5bs9waD1i68kYJs995c3SX8
h4nFCIE+eZaUVSTCzld59gh5j4fc1TqS6Jn6OvYHXd0akoFuCcrmSIV/OzCYXAHT
4gSvTn62RDl2bclJ5OcQpUIMym1knH+5mI0284cIPB9czAm+huJUsxQ51y6WAcQ1
wQ4YYOxmzKHrb78JGWkrsKPB3CWmTdrrOF7bbQPBTss3T/H1A0sQmmVazjJKBNOc
QDw1PxV2KywiNLET1Io1zFPUuLSm6xGF9rHIrYV3RBPVvxx+g6xLXHvcKRVOPSVi
GA/psaPjtN3fFqOaAHnDcOR3m0K97cCexWSSwD9DnwzLLCv38kqX+ZkeCi+dXs8d
N32C2Shbto6l/u2CCIe1VLEnAJHP89a7Ga8MgVEPaIMQGY0Vsd1eq0PlymqDwHz4
FW7jY04EoDX2TEirW4xqjb1ZEFF1SapYjZoymnbaTNz+ymYdqlwAL0R8aHHCF+Dc
LvuRJVZbUUxYc/jKxc+g0RQ40gqKKhw4ajbYS24bTJiBLwvrdnuuvdyN7jEmsv1h
hKxrY1+dJxKQIAK8aI5TsvJdAeDv5RHDU/vHiEVM/xjtn90PqS63BV65ZicVzVtf
A/mOk/v3ocQeEI1TWbDYq64TQ97yxk7m4sUA1ZU9hHd6R3xDJ43S0dZw7zTGvHn0
1fCubmc2AZ7aPAXZd3XeO6yAFKVAP/N1qb9PmEQUkAyCNIpo0uU/P9aSNpvUg0ti
/uGt6SRkrGyYfwbhu60BQc3kfyH/AfkNDoY1lldDQmjMjF8dMJ6n33vxfzKs/uhF
MkxB/y8i0oB1O39cPCNwV+IGQ7bpXd3duJECx68lfYq6HTQQ+gML13bV/hAv2Fqt
2KdgPKeu83oQ7Ydl2GWmEpTZvCTEPPZ+ghtz4CVwQ7/NIO2ci2I/SSEpQu/grHi4
R3wYwiIDPueLzbo9WOHx32DgZEimQvdJ74F7X0MO3GBSbPQFK3cWrZ4oKoGGwdht
ue2NBHtTNtWLM0TfjtMWgJT5FBmt0BFfhZZI7xId3vMAMWBJOlwJuiWRw7FYE/x9
XFnKPfyI09Mp7itwlsC4xeiQyjdHb7zvTH13PtgIQ6485ekp+NLOwEckEwOnLc6L
P4YWluA4B8CKCuFyi8aBIC+daS+/Ru62sICQnq7oO19+scqOzKBeCozoaNK1IA4H
W2lQ5rAkiJLY4BgCyFxxfnXuD7xmJrvJqUvUo7nlz41UHD47vJlKxRJPrntxg9QR
oOBR/2mQlrqHQfDndFjRvz8CBPfPRC63VD5104r4SZkI1YsWbFwxa8t2U6qwhr5h
4fIkcRovtWlTQjocz797fTDA1fPbVRgQjkCd2lwgwRQf1BYNRuu35FYaS0+4FO+j
Az/9/iUeFGiZZm0cncqaAQUadQgENIh1Vv6izON80VKN0g/VpS5aizJporo1y5mv
ZC0gtsOGswEe76ClXahaCuK4RG5BQO2Vb0HiE4E2pv2IOPNujX+LFA1n/XDvJpJT
77Na1BRAKsxLZ+PoiNnXOAdh75skkCACXkPrYW54a1CQ4qqvdTHC6oXtmGmwDdtS
JzCcfRlv66CM+BmKqsV38ngNLGTQjQQTmDtrgj+e6k5dtUF/SkZ0SZsIuIbhjwco
mJJvzcNQTWeYZ17jJD51WAJsYYmVireXy9dQI1OcOrxDup3E0EsGDKPLEN0HzD9L
cLBxEo0pm6YxOFIGGN4Nxhh1eoqwa1HbBfPucugF+m5OC1u3fAP+QSzUv/GOcKJY
calK2ijaQym51gmtHfOWQSezoTEvpQHETiYwLK+If1oZmOTSGd7UdWBXzL3fAoZj
kr52Q2rRNYJ+DLiC76k1edV9Bgwsn1+TwOYKrwjPVO0pToXt76oZq60w/3fpiQpZ
LmzLhVsmhl8aofJYvZtOqsljQKo96mXD8xSNw0n2R79UTx1W1x2UuC+TfQZpQTDt
aY0qXFQwrayfPZruqW/BeYUkI+8LBxF5Pwpf1ry43rWSzCRmsBz1UgcS6wm9bjNj
3hQNxsF+8RqgyYqc2tU5MgvIJLPtRo3UhCHbrj4ZmwwRCDQSG5Aim4a1zbZaGCA/
ABVCvORBNwmE12969S7VOwC6k5A/WZel/a7YME8Pgy8kVfkzJ1acLZpnAUva6RCx
HrGBFxQo8MnH681KYk0UG030qF5UqIuml4E64Dgf/LoaUtgqwQE6KwW0Jfv8QPEQ
J04OmFXA/zO3qnQo15y77rWdDpwS6qb0JL5ZxbhMWiX/G/ePWTV+j8dqMmaW2ZUZ
JGFEnDMl54eDR4ydY6zj/SgADR4OOTZFbicRVwzpsye8LBpv40nnr0vUWzhaxS4C
jqeirHwV9feFRTEjJUYngFXBloYkwm4v6whILPjjN0/5PvI6bZGGIghlMS4T5d3w
6oavtOSZ2mh4LNv926A8KnYPqIkUthfTm1DO2W9W4AWouMMxYM16dUlTpXTBZF3H
YmhShPgyJ8r+4i9UpFs1RrFFqbQO8qNoYreD1AXnSM7EB+o+kTZ3cwjB3iSLT4YL
TbGp9fRdxIzUW0xvV94eRItA/rheEcQGCmE3KgqwIv3NgQHNCmjGGgc4A73R25z9
6LqzslguRxNnJ14iouLJKitFkTKB4BqkdYKbx08kqaCTUYJZFJHDGMQN0MWvVKCo
+b0gYN0S3YB0VEOaU8xKZiAyn7WtwT2YnJGoSgFN6f07K2+EmQNvfn1MW7l9wSwF
+ydKg9p1McUuEWK8aMCw/75U+ubvQnUTNPRmjjBDHE8wHdMLrR+4ZYAKKHQiFuww
toLBuViJ2hn8vbKVyM+GZ7wcYPCnU9A7CBmrkr0ZDjAJYrLF1t2hsM50HlzTDExR
wAN9N2crXqKPEyU6ZmmwRQOovp11tjV4uzT2KjmgGpf/oOLG3KidGddn/lxxIqVV
WEKqSUaxJevEtkLqh6tHEXaBpCKRgG4gdpwpfMhdHj7G09QlZBhJsdZHgAQiXNgS
trZzmqPeDdXhevMnnxPD1MohtapO2BK7WOpOxMVdqzh0Q2b1Qf0lY8G2ZOx1s2Wy
Q+3YVXid2wSdf1dYrptaP/SMhoN5NNeGAM4CAO72BPG7ZACwpDW48sdOtxYpUMeL
Z4QFbcmhzKFIMeGshMPq7D/HMeWUKUreOcX/hchmICyDkssp2qiEVJSE/ZhgzLDu
A6ocw0F8nPwHfFaDmIZgJAM9noR9CbwalMf3tEvc14W7BLAKr82WOf1fE9tgmxTv
UOKLBWWHwwIvvPTqJmtRf9D9jt8nzPRJdSLuSuZ4hrlB6YgkRsMkunPVozUcuV6Q
xpHUgUO6xTeGe/0dHSaY/NUhCbJu2g0R6tzaRFNha2Vy0zm1V7D0EK2Do+2T0vnx
Jsrub0A63bRAQKu5GRNg8OeBtYJv+5GazCRTcAKgjDkrkvQIvdBiFy/S0X4gk4gZ
HA5sgybsdalhwz/oSi9CwyPJhXIMw2shNLXpzAkRpNSsWWQyQmGOEFNQJJs/bh+u
F0kWZs3RSQ4D1LFGsj/57O52E91dA6RXLNPsJi3mqcfrPpN+4rjWEPAmRWhaH61/
NgnGIIDloLT/dnrhv88s+CxAOr/AC8B8WbQaWgkV9y1SM9bfKHXOSgDeU6c+LW5f
cLD8TkH015xkMEmjFEjb9TNQFi93KCbXtJ1AmDyFSh26RZFdbWsDY8g7S5qbqWNu
yHFUocF2K1XMuyxVIDM6OzjzyJEaVqjZzs/C1RM2noHrPfMgaMvRHnfLuxb26u6O
SAANURXqUreYyCVmkoie2ebYDtHAVxj53IV+tnnJM/u00DlPLaMtbwzgLD0EOJSA
5A4XgX3CE60uJN0+OWTWOtkOI5q2Z9piuJtQ9Ck4NXVt1scQKPlEZF7kmqH/z/ov
dtGPsnkHUzOgejYlnDKsPQgwz6CpyyBbvRHJsASBxYXOZsRPa/v5kn+pVrv2hSRi
3y0+OLc0OfzblG5ix5JoypxKO/7U7jYDpnZ5mIFEbQcyN5IFe8NK4WA8ibYvMyjZ
GXfA9+vgvLTuzVDj57WJ6eWbpeLZGcyjYW+Xq/5gHcMX2+hBh8guQPzn8YfSo3hA
FTjyt8ZI2h/8KEfNSAOsYidnCREUvz7TRm8NoenTZtSgy404oBAUj2ByFu559dzl
9maZDUMpV2Gw4ttxq5Hoj1NJOqsIulmpUxWR/qC/6pMv+GatQjsamEvF7lFHkzlo
6cCXTIfl5Qj7Gtw0ZYhKE8+ioxHbv9HP8VOY4erteSaOmr+e5oq4/kr5J/X0eJns
e2m1wYIG3ZR/79xWHS2H2a+t7RTOlkTYDBzjqhXhq0bJ0w41oD3p3jtyWZa7rwIT
HASeL9DIv4kIn5dRsm3w18MDTbamvLmVwAtB6m06+hKuFh7NQrPv7a36cNnnapA8
xraM9b2uIq3TCJSZ2Qw0F0R/DE6gSxg8x+455s14MW+AW2bRZv8qY7+SWK4RHbfb
dUJGb+9MHBbAkfaSOU+03b2K+8ZZg+aqrK4Id/nZqloi8RoTERH329ujAMGFhIzF
J7QzVu0JPdLRdaheByB3tfTei3Q7n8Z9rdu4rA4zuCDVkywTiAMuuGUVLiNMHR3T
Iwd7AAeWsbAsNeeU82hqByItXOnNE3XY7KxmqZQ9x4Yw0ax/wl3rLf/eCmSikGLY
VVi2RqWBvbd8MI518iGS5qLqn2WzRa8yWKbJEgwtVSXTB7j+WJuW2i6F01a0Ghpj
xQvbrefTa9o1npZfqF1LRz5XyXpZ3BD9uB7rJFHrYJ23IW5QlBhJjowWeVwqpYIZ
GKXZ3gtUUZlcBP/IFe12iC12sibNqiFfmCUeohgiun6o6iDtbDUpWmg1YvT2v+VN
ro1bsLX3w04z9Lz4tJUDmeHO9D9SVBMljpeaEyTB1XUTq2XZ0xITps5gCnNRopV5
rujcgDlvcPukYrh/sqOd4oEKyA4yeWqQlNMYtEyPIruaCqLDUwTbjMtU72iw09UC
cuBHqpyM8INs4HOCMJUPubQHVhg1GE58wkzNT4OBqUTH/bbiiUa3jRS9WXnvl+Ee
WTQJE9jC+CXETA2pyatBU0FkcrCsDqUCOuMkcUrMDN/gZJ3upzyf54wVwnI9g9Xf
UZ4fpGl4OK41M0rcO1evws/xmHqK6m6YJUj29+U1rt69NmhYnq5UkdBr0lqV/0vu
X9NM1fTMPpH/PmxhijKGnAkMm9+pO3ZDBcMYlyaaKU6GysqD06PAJ2WGyYx06yKe
nTMZzI19uub224KZf6QbBCM4CNkDjYKySNESZDdkHd1jtq2U0bs4jH6Znjc5eLZY
DGKiJ0A7qokWFzqg/rzQRNwfgajt6vbTnGD/nFfZXXzk48SB4b2FWBEIQUKgyg+j
OKJaG7kItR89IBbpBmsCJ8F/y4h4kcN1YKo8SnXhJDJWmVeVAzKLuqSFbx3WqOSH
5YVbyw14gbauNKhBh5xMDUfQempqQsatshEaFFvJLVrEEe/1WfGnz1sAKlw+s8y0
v4XZ7gsir171XHwCkM0soOtK+zB3q2zMesuGBjeuCa9d8/jGKs6cQyTQpXSpubkM
RAtcPCauD7IG6u1ZJ/Wna5qkz5q21nIy5XK7No6VpovTgzhT3QtqAfxx62SYtscb
iNVKfUflIZTli3Q/HIDfRoQ1p7tO7HuwTLcep0jk2A1p0E/TjXRHjQ/s6Ozgf1ow
/BNC/6XOxjkIqp1f+KK9832WrjtyEXJIrfYs0gF/w3xEngfMhKmb68jDMmy/xhJU
yMMqNzX5mfdrj3ao45HfgX/VpKOqMYbi84q6k9woTz2Lao1uumcg1/ldOqjPFhsl
NUKw58Cnj2Oni9pT9HLZhcrhLj/5MDP11H6q8QjhVs5cLoDjxKMFE5saTPYnEHrM
S8yzfPkBrorIbHzG6PtVkaI/yyWCfuzfAN6qFUyk46ZQvE8riRvg8mgYdxXABazT
v8NVn1hltiEIauVCrYLVr0Khv4vcslmjm2cEzyJKtkTq+n3YyVWj0+Rf9cu0WnNK
bhw5T0aCykFh+t/07Tw2+uPLPm+Fiy3n/mIULVI9jfdRDu5yxkHlccKeT3Wz8vhD
sfymuRwUYRo0FCnrcCl3zEgJ7KiLeXKr/ECDJDwi9C7zsDuMY+kAQvIEOktnuqIk
ja6FiaPCc//6o6E2OgK878NCzgrs8oeaBe/3ZJW/aons/Uhn+93cLc2g0XdhYsSz
lllo4HM1kyOvwQe1YXQ/KAmHVqfLsUeTdmjn8dZnGOH0L65wcayiVp/xMLjexydu
r4untMJCJPAEYhGCKiRrkh1Y1QMObnYJcfYp3/6+Ba1XNU+BOaLlJorAJBU3CkCk
b9lQIa0FHHHHinEqrWTmRLMDpRnLFUOvhwxEJ9ZxV4/TrtIV7rI5uygHbuUBVHPK
FqhX4NIyZGT0DA4CYLJWEemcpiBdIL+hCd8829wR7snzsj7sLq72cNFUgo4oGXxh
y3KM+6UMwVG27jTMpek3g9J9kQ9w1RlYyh38FmV0Yfz09mrNUI903ktTYXYODD56
5YsY3eMxU12gzCGLOk+SkBcFUBu299xB61NJ/ic/XZC3IVFPTR/d70eZZMcnrF3c
TJOKUh0X8Xw53S3TbiEGtnGXPfWCJ+pyYCx+OE+0tniACB4op7Kapmhj6WaqDtGw
SZCkuH7noat2Fxbw3CwtBP5xoRVxujf3EMdnLi8UjOSYYpjiZY6uFDw9+h3X3xeb
4jz07/mMmQ/xiaepiA1F0Vyv9SzVN5ttdqrAKECm98SoVDjup7wLODO1pwgvRwPK
F9TEcasH7+ZsFSunteE3YVh7z7L7Y5gnE2loGbq3GfEyAQrY7KcoMajnh5Aohghf
pmcp3koVllX57pWGVoFhMdtwtBNoIeNw/PtFpZvi1tZms1VCKY1yqnBkna3LshUl
NbhkIuAvh7gf+Ys6x+/3eXQQvp7RBPtz7AU+wcnD5iaOsMgdJN4lCoUZwCrA7IBW
tX952VLPtaGAH3V5uRNnYKHztxCSLuFVIznJPZjtLiPtHcHT6hNicD0rxw/KkFC+
ktWqA1Wu8YAlwdClhQnZzwUkK3Q0hzPfhsxkjjy4ntVdbI5QexkDxMm8yrcMi/cb
2/3oKajoPbbKR54x6H2pTPMmg1AAgEbSS19OXMZ1cVrwUl4b3U5zAXGqnU/8yRmE
4e9/t++k2DScpgwvIleEceicEAxb0QTq6kZJ/83knkWc/O50XaWVF14In6kUj2Oc
w1oZ5pQHRjEuRiiqUFs67/phE/6QFhWPpdRd4McxxE+vp9qFxKbWNm1qyko0xvgv
aPzQ5Y/wi3wzutAW/4M+uGKd9p2yg4iAth4OOzyeyQXOjyY4bB8QmwMTK7TJpnGG
WjBq5FAIkYyeVDNZ9uADdXF3NYngEtVs7CEd3lFvKgQYICz1nbzIxbNqxIFIfZ08
la0sgbtZl8E/sImsRaqB1KDByF7wC+69f4JiUTv8CGdFgKRxpHodY08iTuNrc0iV
2ISCpEwrHnKfkTZV4vsorOR5I1d6SQeby4smOXW8DMU2HLSFJOMsfOi8/3lcFGoO
SVhS5uCnGdi4mAn93RWdgWNrccQo3zV0MfV9Rol/EKu1PocYTYWZyuzFnrLIr3ck
mKObuUITwtRV2ILy9lXR6ETOcR8L+kpVrMarkwjEUT979JnK0DSes5GV7aQTlBlU
ilENHTX+i3vgwfy+CsyPPKjKBcpiz3a1jACs7TB//JkzrNq1SHXigF+XZ2giM3q0
JJlP8TyavO+eRqLSoinh+P2XqlxaSXK2uYFvM39kkKsFnzpARJvNG5GVE8HNIHl6
9t1VRW5zmqiWdhzGx8f5x0yD3jtZgfOSkduyLNKdHjcxFiLyCE+WpqrSnkbcE68Q
rYAoo1nYg/C2/oPal6z1tXwWzLNwPEEi24rfrzfcmAfg2Sitx+4zAHHWJpk40xf4
UFnLfUYvnE3QOxOLFAg34crok/uTKwD22sL+2C7wzKk9utJhC3dpL+eie3BK+LjO
eWNrVE3xXvHy5kLJGi4FAAl5lwyXAwsFFRIwDUr0EImzmee/o28tyZjwyZRCXrHK
v84eZW6ADdyH66JDSXZhJrHi/YA2nae1WPBVgIsX7T7qDTERrzMMSYo4IzBPI8du
0ik5LzpGvLMds5hLDt5jmCqohmd7kTYA1wo9diBsPnm9AakVljay0ZMjtOkHYqFp
n07yvawu1g/QkjosOedoBQ5pAK945SC4rqZKjgKZ1PlO4bw/B9SN33miD6I10Va6
L64fP6WMSJktWtZnYiKVIgarxQ2rOgd4Qyc5zq8I07t7lBISgQUKJCdEPNNX37q1
EEcgQECryHrA2sqi7GJBNYjAtdnOZ4YC6BatQMf0Ugf+BDrMBc0CV7rDU8sUxcTP
J3ed2nSS8BGNnWdKKOe8bMKXHBK2yA+qu/kUEByiLap3j5yQnIn/vRtQfd/2ySKh
tRJSVB8qpnFIGiBi72576uH4RUDJpVM/3u1Yrj0fvp0bxh1Wwa47rPwmnWsJt+uQ
tptb9nnTE94X7zZafpxecApz7x5/n/L621lVsSd+qaGlT0h0gGI69u02OCL3u2Sa
ylw5uIn47j+rLqpC7NdvLm+4zIu564HVS0Z+fOgb+NsX/QbErPM4R/yNy0a48FCT
VKvJcx4k/YIhiAdDnbBZmBws8jNyAriAihegX9fzt3bqIzQgvLIJzVQnVVr5b8LY
Rt7pr9+nU0LJ8OCHNyaQtJFcBGfqzhLC/z7fKehNbIizhHQVgBGQC8QCtcTerlGH
f13A+k6Kt0zg+h5f6W+Pahd7DQ+S6wP1LH3Xv/hFrEG5caESpYX7KrR5fi5+SRpq
j1NJmWlc3bujUyLwEAw6q/9vQ9uFb2UfthZbQe9r0KLGdGVrXd7NR0021mm3KBMr
xdSXHjjYfOYafNFsZKc/5stF4ZpYLNg4YsmRBoDOMiRen/78433/qwqgeE1QUVO6
Qti/8y94Ak2DzWx+PXAu6vIa1C9NjiVk/HGAFgwvL9zKulnAAsSyVxWs9sAEX0u2
TY8UW8PvbKotBRnb1bHuynHg0zhjUd+I7RwKQ4itMHSfZ8hK4uxY7Tt4NUawoIEI
kC8q0O6XnDEF9oX/xcACvNdmSCJQPWhchRq1Oqm30bYYj9O00wChSwPDSW76KchM
uIB7EUDJ1ZGV0CxhcGwI5cVXAqmoN1htymidQ+tfr8BM8eMJPsZK0eZo6n9YUbm0
dDVvnoVkwyvBn19pVJiT9JeAXpxycRhDK1lViD6MihRt7dA15CeSpeovbMUL2gGP
5tXj3oyxOM3xmD2C9zOOQ2hq8U1AbjDQeyytzbFW/fBTbzfyeQiJJ8tIkZRYNZ6e
9bos3IrSLIOtCWtljuDACX+CkI+O6oPTuCwURjUddT7N6j3MTo20TjeUsoEatVXv
XanlAzl0hb3uGUDg5UxVqPVqhx/2GkjMD97kpI/7Glnba8Kfyv0t0KuwrMpuS1wX
6myVN1MmCE1awS09MkciI89M7pUQk3uSS/jGoyISrNS+oe5va80hFkyoShpwCeuV
LtPpmrl7o7S4k/y/UVK8md4cbWxc5qu6i5jc0R5GTlHtukW36DFNKAhs7D3K+jJV
cz/ipLbR4pQOP3yfiJgd2MkCVhXirXfzGO+FcXMj/S8duZ0ElgBle1AsGGWcR+j8
cWumQ7xFDBmJDzteJrKd0NfJMpkrnW11qcUbMdO6o+KUSZYbq8pF59QTUCmBDTpL
5WNTDX520kEJSY97XVEEIVeeCZboOzx/C1tSPrm2pYwGogiRUD5FxAsAzr9Rxpg/
HkyilKm2Q5gjUDVauanSnSZH6FIxNYmtVBk8vT4of6zR/oLossm69WSfUKA6c4Xt
AzecbrJ5SIDuVgvvKjdlGxcUt82AUTZ/dEg/yqgmwbPgJpjgf4T8SyNr4lX/3ye0
yHtIbjjb2/ucFGhGT6wwjfm/P/MTRAukmw+j/8AMkUp+6NmnSzw3CqMocb1UlpeD
Cj2MsBQsLSK/iYCHc8uEZFyL7DGYzgEZO1LcqNTeXfQybvbuDBVC4agzoGc9fa+r
znlAGa6hg05iHVf1oKoeuuEvM2NY3Er04qkrOSjTREKzC+EyUxfLY2YfvXRw4ZXh
9lPRJwP25n1mV2jixIBVOrDwesx1sZOkkZ+LPDFHz0gJTHgI8JNjZ6228/79nigj
pxMKek/SsOi2jCNZbDOhCSGaebJrZ5QaAZ56RUjRABB6CdV67NT2KzbwbSlAGVTX
ibA+jaaYnO87Z0sme2pHM2HCkQfuFrTz7/1zJOo9lArZQcUBD+Q0J5et4Ve18lUM
KtN2WviBI2mB80O1YPwn8asdZj/jsFHeZoQAUyrmPE4Lj8lKY3OP4qf8fgznaT5c
C7L4tm+D2wr0sEFh8e0oNb7kGgumk+HavHOtoae+Y2GxX7+9nLioYbcBM0mD5/vO
YsM8ekZJQFEMaw6/jY6l2diQF7Pd7FOsZkJlGLAWFXHukhGnZg73Kcyz3jwz0Rtn
6gfsHsmZsnN6ZlTGZrFec+uVjUQeMuybaU12mIQqGEp/oLZjqNP8b9KsFKpB3p1j
bXrABV0aEQCOLN1f2sRqxbs3Ih378hv3wbxqVmUqalyc1szFKoVgBVTJ7ONV5UhL
VxAmXX32PDA7V3XbJKgaVjrVTImTt6dFFThb4C99D8CBPAmyI7um4pe6IbSQbtHL
9xtqYdGhiQLpkKIEabLSxF5UsEJ/4QAiEklsRfPT/gvCyYKQEJ3jD7CMQIqlx/PZ
l8+3T1zhkujg1cNsnffACCg2hLQi00HO0OPzjzJuSC3HXfaGgeRuK0CxKjT4kpFO
QBmTvI9o1KiXu6sEj0uccuieDsxJd7UHlZaai9dxmIssJvvVli0jK49iUj/Dmf6S
wRfiqBnkqhYAuo7jfbaqC6LeE7G5fLHINhToIl1MyHzB6ZAtnRZ31VtaOmQyJ5SO
ryyjagxfAOssjk1MnSVQpJL8CmRl+LAPUTw8SOduDh8O85tX2g3vKFXdnK5oEHo1
lSFDOkru3jvNeWl9Ex8iiwHjT4/OoXc0Z+NWsGF/nqptjUVJVUxkSAn0Lw3Z0a6i
XtoR4OcFV0n0qdrTzo/j80y49piQyd6c046fodyq8HWZ+lYms5kO+5VKWGnIAZiJ
8fQPhXXBwvPXHcxLZF9cJ0C3UeX3jZTpbWQ5H0NPE6zGl6RUXwSTAbZMWBnQFiB6
AjYpMKYCwZNZQIS2zmOOmx7uWb8L0iJGIbKyLVSMe1pkUZ5he8tJEepsueSEPQOD
1tSkRE2MwXqYq872gNowYiyLqXMGPKKjAlKSE8Q5nOx66gACq1abpy5WNlngOqyC
TxD530SnmZMVZHpCR40H6keCdyQ9+iyjGNaCZu+3EBc3xBwTtmBcnEaZqMirrRer
JPpe0N51sgtsE28s6Iw/qjbJw65zx6p+i8RQyuIId7IFZP0buUGegMGV+RpfNcxU
Qkp0Tp5JOAM6EUB2q42yLcty7dZVwMOUXATfw1rL8+YaGH1d2XIaX1683xNuA7XK
gDx0N72jop2hmMYppnmG7/MG2WZMSMCjO8OCgKzJ72wZk7A9W87G2ZJUqXdWDRwt
bbkiJou3DNANKCUNhtVGZ5UXPrmsuC72OJB3A7xuKnkd2XGBHc6udKHDuJheToFv
u7tg2dl2BQeRiJIZBE8dVm20yjcexroogxPt0KUiurQjDnkS6su6btxdBTBADvZO
XUnF3PfcnmKG5+UjkB4SF/J0yD5BIKI2fFPTnMeFxMBajPc8DW3RcbZ7q3J0NwI2
sA5TZZNMf5nxOxsbChAg+4nDbGSdkf1XQtSRns/bJwLsuh3b/5biimraTDWjwL+d
r7Ers6KjSnrzPDpAXiHHzSOJYMJpnSxQzhQmyttO5Dc+u4GoKj2cOPQZaaClX0KC
D6a4QgfWtLINNGX7+Vu3rf7FSZLWN1Zj6mXLJjIOl36UaGsOKQjL7ce0AmWJyDf5
o/RYhCzXkPjOz2VMLNyF/4bvPUab+t6RtI95Lgl43r8dA5W3uaVIQgqaDR7GcgGn
zjFmhFtZr845NUSvatkschnbLZyQ9DKIwZHbOUmHSfHXx6Ii2ShPPUjPh5DcF8g1
5hmdLfPclg7KYNuk/EPz62k0dxR8Ie4MGDArItjfSFCT9tKO71MMNHKiN/h2DlGF
TGpk9kPTYgg+Socb6n7IZXZVtNIEEx0GGHzhb9DZmAk3i7DtErduftSO/OlAYfkx
7oS4r2+rOuFM8K2S+c5Nip4zEDJvtVo2R9iBIw6DLQqJlCsil1zKCaAJU/nIYqo7
OafhuqYTIthR3So1m+D5oz8tn9C6godXo7qqWkEYGhQJsRycRH96H/EjKjxXEyzv
fUdas1MPNYuPyGBDH9Q5MZiek4ljG2AfRlfU5CJPeati2xMJ1dntG+kua+4aC3ZS
cAYAFxZ6myxAuZ3z3ZuoY+gvi+YSORDOvLkm6UtdKzWRW7Nue0SzVwRzCfzc0Zdf
xJaIqw2k1IkwgXJwi+K55ImupP1BcFCz0DS+nGfBXaHPuG3QgEGOy7cTdZ5Ex5Lc
8Ig+uStZKOiQ1LaokOiREsDHOTVgHdlLlOzlz/o5T/iIgsbti2Q5ZxzYZAPLTiez
S+QV36B177zTK8mo183oOlU8CnUvDakfy0I2fsqvxi5Z29XJzz5mFDNy7fJ7yGu5
/H8fN6splF1lstBRmemcPWNac8J/0niiYZjzgksHXk0a22GiVQJ1y5PJIbKbub6Q
xCYRvehY8wlNBBkHrQ+cDAVMt58K6C1EGE/5XnuD+5+Df9crFbMHlbghoZCV08PS
vytPi2Rgm2UUdP3UPn6Y2feDaqHtqdbnCVQNdoF2v+dfVpNnyp4PR5gGeOTeUsiv
VFexS9M/o5ZSv3hKF6xV+ud+7cZp8tI5665SGpMSmSVj8vmU/pfuKL0KMGO5l5I7
5hdPDOCpbjg+84zRY9L5g1/tCY2OceaDpFQ1RPSQblbSLxOBuJX8k82tqvIJTbGq
/yqlkS47cWeluf2f9WFWZLMUDH2Ssz0GrpCqexVcGHSi88CVOalPeRfrZ/E8TwXf
G95vwN4MMsAnzObiH8c0iWT+sXjRGA9gQvwLt5+XdwH90Z4vz9y8INkoLl8KhL+P
A3+6gWOgsMswzy+x+Fd+n5B9yYzgB3OuHHrm9JMBjHgIe3Azj6PmeRj/BRdD2IAR
y99QAY4qiyAmCL+9UNcIlFiwd1tC+Vf1j16hm1Lww0CqlhEos42kyb303DbLkNLA
GopzRb5G5soXM/2nEdnu19HMSypPnkGydPP7KFLuzbCWibNOAHTwDPp+7V4SZLXU
bUzsGoFKN+APh2vJOkfQulv1KvwxE4L6xsbb4VMeaf66RVeWjCry2EZ9poxaa6M7
dIw6hVzDDZeCHgkkPo6mQX4XDp2UU0zs4h8lvpFnnCtQSFCPQToP42DFreKcNOVl
bl/5qhY86t5sOcIc7Fy2+n7fYShS8N0NiRrlgO6UyFdfMl13GoI0CLa3gm7/KuOd
k92iSi6zs8FNfS4ul9WEpTonQ0RAhgda1zEWjdqiOxxnlXrUaSsbKLuIllVNOe2e
oMOStgpZaT/7bZIm2Ax42vqkXehujCqrnlSUanzmSqat2iTO3NomAHKZiAqtKvvf
mJlAsiaZMzXIHX8EW451rJ9+2ITf/FxMjpKQYZSv4NFiWXviFd6wDKzhJ3Lo9FLN
bAxRyIZjw4YAfO0fxUErwYcVOfzORc3K1CkmX5WWVwfOH8sQsabNAeIw3U2zunM6
CCJiRiNEAxvO1Ue6NepMkv0McYMC35ONcSaRxYQNSL7WgdaiFq4NTuSKeUIthT+c
5IpGaH3EmS/CIHr9Tt2W3EwvEmXaAjr/8mL4nVY+TJLubi/3WkW6C7I4AmHP5Ecy
x88cEy4csv1NeZom+x4hBegd2lcAi8pz0lf6wUOCw+Tr37mTDmdd6wz/qOvtKJ0m
ihZv89w53JFfz/tklcnAgWmE1iBssrVKGk76wJexL5PkQlHQ8ZPzHnndjXjYEVqm
YzIfQ1S//t4iC6RgXeYbiz8PnFB8+g7QHgysSOHGRYjb/7KMqY2qHiPxkrxMbC7T
sziRw9hTJ/PUgyMjXEQ3lfw/NAoFEEtBEX//1o8oquZ/S2xstQpNExRk76tC/bY7
4IxcMYuRCcccLG+P4yW2zHXXd/N+Wa0F2/lLa8YppWHqR27jRSmvf2/SguHNcQNV
XkAb9h0mFOfqrfM8+L4CgoIRxbEVND/hA0pxUIPP+51oiNQYzg8+lY2gVDb4OAGF
/IvfmAKXZ2+n82Yil+e4ywECPowOwL3fhR+gNX9h7byVJEumZGmeBswZxCw0Emk1
dSQkjAiW4/H7yckioBkAUcGNHDLdX+cadkvc7gOZrA6kTswX42pvbzhm4tGqQ4Y6
/EZKhpNgr9fqa+6cfo2jbT5QpXFB7g3wxI2XtKYxOvvv92AQ/3tH6MregMJp4K6C
grx6vOwzm63lR4u5IUlzIiZzPNdpYQNSNw+ZLCl3xak37kYFJO4vucUACHaIwS2n
OhsyHu+kpKVZ6eKBqR0W4FB4Q3Xy+jza/dU/VDQAiB3MQKVgFLI8c/ahWgY1Val3
jZsPtZM4iY2fzsCLuH0EWaK+EG6QIrpZqRPlXfsZHE9uvU0eaTWLcJYTqTPJ15Av
7qpz0VS9tp4R4AHKf7nNronmy76K24ppOCd0cfwkAybtjQgyDYaEGbz1thPwSINn
XeeLKZoGR9FG/D6klsIiy9jePcZPL7J1s9En9NYvpsu11N5UEy1VcEbfOsmsCkgJ
hRY5a4ay/BQjY2zN4vlVjiYyZhxZd1w/hMRZfpmJO393qhVQop4/w3JgIhzjCJlM
n6ppwpCCrzKU7NZ88NE8jxrC1YrkRPKhJCsFcypPmnWqQFMC+yNK2WrBJVIZrm0W
TNDex5tI4NEXsYfIyGy0wU1RWgKONdHSulcCVDvQoxneQQDPR/szzwMRNnM9huBX
YXpLPVfay4NQ1uNJWMl8DKsq6+doty7KdEnVVrlOdToNugB2wIL6EmjEKosVuOkf
IH5fK2oqa9T4OvSjbi8G8jsF/Rp3BiGLTp32Tv7Wa9x6fF1hMnuGQzusrWXCsue0
BMOkNjGEQaWXN/QDhgL+eXWrWzSrdk7Hiq6B1dU/qxshNu7SPQxAiQFqdYeTEugK
ZclTjaZi6243PcEutETtsvnTrovhFmMSXg3xhfrssWysnlqLh4XnRsC4mIVsBgna
Nl8M/p3qQsAiPPpeT915uvtD6EJqHA2kw1FdOkyyYHmy7H3Lp0ZQknyvNnqawgoT
DD6LNV0MJmu/zFLBaX3wQeYc2jOu+lDAUTtTOlbPaE8OjKPpVvAvMT7DsWpYBqwq
Lb7WsycYFmeKz1VxtYDjsS4F9+vALF8gB5moAlHgGE3sJ0bBamb6fQBn0gmHEVcu
12JRyPHhXW4NspMn9QTJ7AOOPnm2qrTvuYCjZ3cKY5NcA0lX70L4W1pc1iIRfOtw
iLcexuc0/aJhW3RlW4Hel5aGFXYcMnf69x1oKrYrWGXosMbXGFQHEy9J8WrSsgfh
lhFQUj3p8wx6zdWDybg2tROMKJKud5WsXDE1hz2MePg/rDWX2HndaEAZXz0bIFQl
W86buEKKQjg8ye35omKW5dhkrO6OMrmHDp5m8NdnXsCsDtBIvr7TX1TaeZhNMIVY
BzbC1V/W01VhOPoO99USDPtCwzuVT8w/3KhVQrpuuIqrtHJ5Td3QR4kH+3wVAqrd
P7W8XH0Ki2TxijTeq7tAY672UJ8XBFM2lDEm6SFOju/ufMvLaMTGBJkllgKJJnOh
++FYFvs6d4DtGO742/ziEym106zs4ngFGTJ05nyORN5kFOoX8T31DjoNbmQ/xe0A
+/J9ZhPCbzmJPb3ulotZLaVjmzJ0fOSWcVOLniFAVfTKC5uG4SUCfDmQI5fxqzzR
miNKPhK6st61NE2diF/sj9PrCQnFoVr0TVE6XKDys0bsCZWpsStfN//7quAk23hs
uZsnWJrD1HF0EVGquVezqtTriO3BOqn8KKg1qJo4Dk34UPylLuxIEoikm/uFsVIv
NgCH7prfiZ7jgEehbkYyaPE5WxLdU9rfT8uHikC8TMdgK9kinVJ4VE4mdrmcxMJj
e/jkT2I41PsTOIh3uKtXXjxnHHLogMhOLcooGDEnA2W/79WykVhhk3ynj8JqlDZG
ALFyuuJ/voAEtaYItREo7CsJIow83Ng5KeqZIyw2ilyY5C+ALnNjaRyhV4sk9yU5
74nEH5jCcs7s/ug6GDeHf/cfDFdkoVDBq1Q9ciL475bDCacuSIrX4VYqoAt+WA3x
JUz3aEGQu0wHsJYU0mNtQGmjOwTEG0Oj/bJ56F90facvB+ShPvh96RplGErUDuKv
1/nrVVfYqj6WBKuhUH5+WvDf2vP4FT3KogEx32kPwPabBrwSEXmtVWwBc3KlAZR3
j7IoIUge0fwYIold3R6QC2TvyttwI0KhiCD102C9f/M0Fg9lzziMl8fH1L0B8HQR
aISblmfBOx0qHDwfeygDkbntzKH+3c7RU5l0bZNtDa4DybwPPU5fjWdKXMTUaZVf
I1vg3zz0ciSpZBLNjVJ+xtCldID4Y2QGZVCKZWyKWPcNIkAMQE6p43tpZKAIWh8q
mTU5iqCC1kxpBgPw4QAAVxVrmdY8ZXl9FrJMKK0mrqj8AGOrEVKxA1W90PO0SK+R
s2FvtOzr26SwZFHp8VWv8HAhq48Wxgm6JZk2KJzOuVzCTKLyZggERG9kJ/9ANXNP
R90ftmqLS/dS3DIwce2aQ93XMCNraBjxBk8+Ek+UuYCR9dIkiO+t/ZHzbV/Md4/h
t+eXg0ZLN+U/BDD/SNa4dRT1c0pRloQgCI0mT40JFMyTWN+NVligcCSYAaIzR9SE
1etSTR//PyTA8WsEGtvHyQT96xTJ9Q66Ngef0xsxrNgePpwLYe17EJJl2SQKuro6
sKrQj7+1Y36WIk2RZNG1HxDVs56IXbI3Zdi0CS8P3EF46JFQJllleMGIm8Rx1ldu
98krXfJD+1QGvVUaWhQnFCPHb8qp0p0alD8faBGr/dLNVmtPSL+F4VtatkJ93Mfj
B+G3VRjRd4blekWfpRFp6WpdNKE5DLbliCil37UWN660sffHjaIP62Q9iLuByUP6
fpHnkm9Ks2dnu4scE5NM2yiYgLS/irgH1XfnrXgAmWCF4umD/zksjNh0pZjDJTe/
0W8/N2HX8vysmk3QVIkJRAh+qHmswTwf5c2SdB/C2G3XI1v/OJLJ1Ri+PnszeXLD
p9zzGF/DxZzyP9VvZq1THffOn5uH07tkkTWJaV8W+UbSNOozUsZU/k8Ggumf6WoC
uCmnkQ9H5CO6mp0KeseTxVjKTZRpjM9wTCO0xkU1w/EW1VCAQ/tz5MaJ6xR4sbST
bF/f/ESY5gAuBbrv5QeY0dFCvWBZtcNSq0Id+Tk2WadxDTX5BsNUypo0yq854bku
uaxT6VQ8kYd4RaKPf1aCsdVionvAzzNCEbxDG9n1LFznj8Tc3bLUHfn9EBQbbSav
mJEweS590C0R77qGYgFauqXwo3Z+h/pH4cvJedRFLAezTQXuivre2mgWt9PFik8Z
K44nF26QEP5ux2gkIb820j0me38txqK206vBrkpbepLw5mVhcDVaA1hqq69HJIfd
mkL7Gi9Cg28Td2PBlZIEjQU8T4RTShuBMF9UyiPhJVDX2FT9zWo/KpujIuWK7l5h
i4Ye2968rzrT5ehPuH9cmPvQlB9/wxx4sXXOrBd56bJrVbepyHdpeScCV47wita5
s0jgnlVp8/1HBZBMPvUwsIRgfDpLhvZ3BsRc39lkf0CeHiTzjjIhPxSOLRnhrtcX
01bYpcwa1SuKs2X5xPWxmG7ntFkAfxd07Od9UBJKC+/czDkEKIJSbwPp1OsVoLdo
A8Zh8CYjKs8g98rwOcU+3jnk/mRKfBorLkJXm2jg++9llNXkC0go+RLJeY3z5XXJ
M+T3sZqusenPtGbZcsH2+elu2n1NSVUSJTn60TDnwusQhhz+FB8nWWNIcrb6j+p2
Uf9V/mzqgNYlNsG1NZUzbb5k4NeZlLbKaIyZKRhV4O7FLWmB8hV1fK5+WYVUC7ii
GnBirrePrwHvnqZPqREJ6nEA7e0wOHfALeAQFDu6bLWpIvjqHKxD7b8juOo74Wo1
3JSjBf70MLpqJeyhXJ8CIrAYGTwosb+a8VDqYgFtwWCM2ZpHBF3PXo3ssxY95AX7
xXewTY7gflsyPiJlEJ2QEE77gt+6w+X3U4yJJySGdSMlCp0X9xi31XZkbZ7IulTQ
PfkcZkJITvKhc/23Z24FczVlKqVFg+juWFhUw9N16ryp0x0cHOW2Jz1zJH88KBZ/
S8am7F0wKSTJUci9axoP69LvDNABm6oun0cr2CtKEzwJZl0R0oe3+EFoJW3kAryX
qGsT1CXmpEwB6YOKZKd9RwrI4cStM0V+eLcVE7WiSsk+vRnWpLMJ62snGFpizjAv
LEKPwf8hNiN1LAp4Vt/er/x/sH77L6hNweCWMqbA7vmWwOVmH3CG1n33CFc0b1gC
REwy8eYWs5GBw1R1ZivrOqVjI684VYe0JUb38JxY8v+4WLsEsgbYFaOomMWLm0td
GsOnyXF2xvJLX4681B7mF7M+K44oBdVVYcy1L4ATOALrSTFjihEU3UxGDCbEirUD
XfuPe9qFq5YJ4rG4N6SBiPBONUYpcCPJinm65+FfoCjFnlo0EhhZUBAvrpHs3vf9
xdJ+kl3XWPvT0tMpALcLgHVQAYdRdMW4ekFEZYrKLwmiV5uIxptJ7ywmX8vv86Mr
QjzOapLZ8S1wYE4CCiOqlVLVF8nNOhgor4Ch5EGUmxjpvY6Ufitv3E48keohS+TW
Gzey6b5Y95TILjDFE15n/PR25rWpgJq/TM4PF5bAPce/5ZXXR+AgOxutybTh1J5d
MwHr6nDjv3/xOAht3sT0FWPouIORsStJYFE2pRzXxuviNoq12MUAsIuqxNwblZp+
p0avCC6ef97TnTINKSFTVCwDXfqr+gEErJfqzyPwCIzCekOp9t+6KjKFZ46LAZqi
azN07CabvXut/9QhpC5tcPwN7F4M7DG1z/L8V1YKsm2zoIIjng0b8AVoaIP+ooi1
sAlMiYeLfMzSStUZUFTt2M2Fh7NcoYWc9ejE+ZuwDAajtCPZbRvrN0eC+obU0ANy
ZjBDqtVroq68lfg7mY0IiK+s2boqlJ3WnhExZXKmGBoDY9hJc4DcuQ/Dw7lu0nih
70XVA6z7bTY6M2nHiUDW1bmmDt7PTCxoMJJ7wiDCLS/Tp8GRDT08fuvxfJiJyKIj
wE9UEmwihqFxVMrJR4P38aBI+iKgoogzY4Fl4V50i5l+iNMsb8KGk2+VBiCExsY7
6xWmcBeADg0OtoY4PRAxVlyL7dcdX1bsRXYAwntFB24BbV6f3jq6ELgJJksoxjWv
uNWElM97hnJzrVpjW2RyNgC0fWiQFnc6Ce8Xot3ut+NMx3wHxCJ9VcacwQbrQ5rS
44GsUSkfFBey7UnaWhVf8yWpclA/bOjsQ9y9xPqBQWEr9Joek7Qy1O+BpiplObEO
WVmAJWRMe73TQZkOPqLnGI5vhDir/BxDdNsS1i4KyotpMzEOA6rOpfNFF42yAaaw
pjc2EiP5pepI/mD4LotktzaEggtOPRBtnQhs8BF5lXvpSVBSgZVEsSNjhzxHeA8J
OCGTWfifD29xk8cqdth+4li1+86DP83mrC+4RpENJj/jVoHOYELZfLPEhX/Q3Ulu
BNSJQwLPUV6zRGhZyJmHUJ2Jx5CYrts2RUYS24jqzKcc9dgHkfGHQClGhP2hqiHj
WJYlNXy2Gg+RbGnK0WEIk5EF2uL5N4OGR17y0EnGkBPdBpkfk2ClEEAyyJN4CvwG
E1mYbuUZJphElmE1wmOy3I6XrYCwVGuZB0tjOFByTfHEsuPj6011EM4FCksra9Hr
cuKIjQOxyjLhBCIubfhP4YZoXfpAC4y+X23RgJABJPQfll0MWG8yM2G3TjV4v8ZE
OqfvTElvkNYf2ZZ3QUcdnBfAhsjLk/7HEIGfBwfPhQ06EEV0g3CmHz1RfixjVWle
O1D7YZo2FO/1IXB+ZJhFErayRxPwL9NL6FyuG9bH1JXJhVkfGEkYL0VK6a/jAD8y
FQ0CHo9KcvraG4QbSYJnWCIQrfk3X2INIDf+bYdp+r3oMXRrsTbtS+H8yX7AE3jb
F8VJV7AGMWJ7Wa3mxrPdbbBel1XwHruJtHG6RD/tJz5WvYrK4E7XEHMv58eIrJLd
VQlPSfGUsCGW4Zun8fi8fg/3XsOkfWgQ9N/L4kJfIpBnaM4BG2yFHvs2zcDNNJvu
UWmAzpFFo3gCQtd3PFfSdLuuy5MnqKtL/Iwkx2ZFrxxeoE6SkY+j7cUK8ywIOsEl
npnm0ZwPALrq4bDsCNS2EU6WC9z0KxE2FDOBhQ1oNMwzTnKZF0a5vFXLuRARpDi2
H+sNlkBAGoiBNywWnhNCtyckmfTdHpQG5nPrmlQQTtu0jzSvEuCzUcmmjX6+aah6
3SC2qCVZal5XqHPqUpNevSEYef+dXPLGUjVP95anuJEA8tJhdpbnXqcTtMPQ9b/b
HC3a8b3PQH0nkkTjsNubLIu6C4RQzVcQrwnNIbGt3FUB7Awlu/AVSRcnaXPL1P8s
fn8DsRhUT7BznVfQTUnBwRwzo/ED4hpcj7eCzZmRthp2gLg9suFCuDQSoNTBSDTu
O/lf8jqdonlbge2YXeofdV20EbFZAjSSOFsSa0xHRuTRugSfJKKTkO3LndMuDUTn
ZzeR4EbdGMJjdwR5011jlRbl15GfZk7TSBGQW6LYopr8KmFjzWv/FuEKh9E9SJnr
1NtNZpPblt8Z6aZi7r54nBEPBDh/XN97VK5MFACdCrdaI6/1m95UoFiavOOds1nF
LnvIZwmv81y7ZOXOTih+oiPSzGYOiWvtL8pTZYJXul331pJZ0Kb9hzJ2hwXVSJQu
13Y8oY3YMbcjhIH9d1uufFHF1mN+x55mIm2+2a+8Vbo+er0noBX6fU5kkNRHuIhK
fog5tJpol8T8+3va2o3UFKaGTT6+wP/kIeT8XMdD8Fr4OxgmTylXDBmCix+dy0VG
3O8fiZxtUa2CSBDDbWRjTiAOccXNDzqX26Upjscw3hRLJIfULF32aEA6gBc5TtC2
15cWCLVBe5iWLxNUB12C7OwWfvjrKAW/dlooj9OZ2pRR2FsfIagYR0pD2MM6rllQ
3rLQPtkBXa8Y/NVzu+9NEzLI/AaQg85hVfGLWZfHaaHkxgRizx5Sz53lIqqljZma
+6vxeGx0s2ZmE/77KwnM8afbuPMmyQtIyTHWtiYgqTvyWOrhtF29zckEn38ATXzS
MVxNbSJ6OHEne+Y1gYGEfdex1dUBmccSIh9HAaPAOX9An1waCvT0Vp7hAFWrRJjV
8DIeW0goYYaLNnwhKzl8jXzB25N4RqcMUUCsvULHCcxQ0o9RQEYjspYi7X6CbUkI
YdnK/TrcU0bbV0xCIgtxMysSTyZA//RwmTYETi76eRM0B4dDCssO9C1vpn5QC60Y
cXu8UpNL4A7cmP8CGhx+gnOoRajTgfmhgXxSQ2hhQbryvSxRClWNy10Sr3EIb88J
k7RItMxH3tuWsqMicehAutwHynQnRKEYYnDIRsOfhKxD+KMqPWHiAVvyNC/LcUVQ
FGAHaauSy0Dq9Jxp1XVm6QagJFE5ryUMF1XEJuTpBowIZl/kVamiLPHTMorxE9xY
JDsUVEX3x1O9MQP4Hy4XfsJi6nbwsIS+PGKvUEWCaInk22rUO4tX8KvZ4GWptsQ4
0AUi6Odst4IQW56huL7qsVOH6OSpOg2Bj3z4mtKb1D/rS6KJj4uxQmJ4Kedl3fZ0
33tPNIZupUhqjR+ld00nBWXKS+++RuO6QKBoNWAjbkzWwihab7x529rklyi6RRbU
zH5Him8+cUHnkR2ISPb1X7nPr5VA1epXAUijBSUG2+6k3S7slct6gZ9Cc7PKCpHK
yGzhhZaAag3T8hI2tbjjfqUIQlS4t4MgYETSdDppcx+NFRPrZiWV4cziibM5+QD6
NR9PrFwEEH4AzyIp5rjF88MlzSJ+22jOdfkdr9abEIvkSS6JzfBkpwi89qSOJ3l+
UU0U51g7u+2EaD6y3ADOj5RcaU0ql8/MK02V0P8Uii1ndbW+WCcHJChdNpTpASnj
FtjttoPYRPyUrpK+WLaptjUFbxsFLocBcqAUWALTknoiMxzvahPHstRzC3+/Uvgc
ljAlb6EQkT8k2h+DejVV9qGHUgAXP7/WZ6yuS/moOjPaExM6MxGP9MYAHKmTOPZz
6BMP/LM1Ctc6/iizvLfOWWzQ6GMvA3fecxuMQbXgqfNK1M2MQXeEw0/1pZzMx3Op
5WPKKiwnrVtJ3hRF8mlFaBL9LWRkNTu1uZxiu4NjAP4Q9pg2yO6naO0scs68vfo+
oKctMAPgTQ+SfS2v5uNJoC1eIqh3lJycTdBGV85TdHPP/0OhJz1zvNfX3XBnha90
niIT5a5dQCkyZupXviNOVD7hhImnxO1EmajxZzzzQvSrPJPBz3WMt4lV0E5Prk4n
R5f+Y0i/7cnINySnuHUvSOD+0fOMC8aLii6yN277M8zEqi4kq3ZnivOvlPVOu2p5
1hL4TgOX3i9CmtH6dl2K6ScMGBoHJJTtNEvHlFpSIvG1HaLrLdqeWJr3F93VMIBa
DSe0vj+GyaSLpipYR4C2+34OobMNfvOXeW0vIhmqOCbskkIbr4nHsnGtfzWpw724
nNZtXBd813Ofw3cZEic32p7zaUcZHT2mLrvqdyVKsRiW31VZt0OhmamhhmchZeqU
oRODQTVScOMrHl36MOMBUqIXgJGtm1bLGuOIAz0psQmUDqGzuG20DpKkqpC8zYAu
ITcRXRwjU9zOVPUY/iqEg1LOzTjHAinqt8Uj8Lb8ce1zX0jM5LiRVr0UMKW+OFCP
sj2BWW+OXraxLLnA/JlvkHNQ1vJvEmltHqPy/2hpZOeTV4/fCvR+ZLoXg25eRXqt
Y90QYMJA7h3FVmVFn3Jkhxu+DpaRg2BpoYRYGUG2OJyhft4j1jIHJiKEVPFcGu3r
B17PtEysFAAaobubAjySAGHmvgV5F0/3PlUmUu5KykCWTv4jpQ0dmu21RWFr0Iy1
x1aqYlXeKfG7rty88D+GO3wRV79VOdI/8XfKIWevrc/7jbR72yo8c7W0vV2rICk4
ttpMbmCi+UziAc3Lc/o/vyn6aC0gGT+J5dnF2zGwXng/Z95rdPGHBT7+ErrrPwgz
Qo99ZopKQOkRKmveKa0UDcYdRctXRTcuMt2tgLsL7MnXLRjXcW4IZEvWGfHIfIOE
E4ndtR7AlcZAmlnASVZ6eUOLOBVWLXQF+Nw9c898NhG0ZbPG7sd8hFDMFTgrUsdM
VXbeHyfRXpckfve2MHA2tuapcBWrEhiK1xUvCjzZAilDZ0RO7Rw2H6Xz44Y3L3jQ
9FPBxXlnbLLgdQlfpowr8X40Dd1YVYhoYYBImQdU8HbEHJi9WYm+3XCcF1/nbauH
XsPbN24d61BXMUs6VE54jRS7kXu4Fh5pcG5b0V6RozpKh7eJfDy5C3dMztniM7u9
LQBs7qEnYkIADrufC9f1PGibgvVrnlMTiUjw+1ZFHXf0iJxOy6HX0VsFw0CutpWu
fhGBu1+EHm7SAZsdR6CmsJYTTkCirPui4RPkivBh427OvM8G0dkS3qK9OsZR1lK4
CU3byNAOVbra1pKnlJPHJ5StOw+QlldlpUto1yqLu2DxM27ehhHbZIDARrHhl3Ul
qky4BP+TNqSzz0JMZFTEWllx0nhwrPMcRnqne3oF78ngr/yIdNLsNkKCBkBSpnCC
BPsxaNV8urbo/58CplQkhRM+uAHa+eALc78FjikIoz0svVRS5z6qY5M1Ctmh/GZm
G1B37fuwJ7gUeYZN6q3QPSe+x5ssWrEdhg4UZfizUU2+feKa7xQtBPU6c2Y//WGA
A4rYJFksnR/vf/4H2EEkxgQ7pMwb6NVhqceH5w9nnzS7ESTB5CWHyNX9198Rtpuw
8/UX2/Lkbkl8RZ86p3S6QRzxj39Cb0DpLYOLsNfJDXGScZt4KdlK9tn87AduP+mG
/tkgoFOPC7GvR58wLX8qkuIhhQCxExiV3bzp7nfAm9Tf77W0vtdHIRZgXKKDGk35
aQDgAHHu2X3nVOKkjY0QVuzurCi2+Ezvo8EFlgl32toOMyUt4EYB9SBYlkOOpDeD
E+M8RN+gZ0geonhRwjC8aulO66c1ljL693klruW4H/KxO4Kr3WcD/4Z53E1zZvOP
dTTHeY66zkhyMumDL1KhSn24uRqS0m1q14WgbUJmRBaBOmAn9QPdbNfzSEHn/90P
RNdnAZnWze6b5glha4P+SUMmIhf5LZmiMhs7KL/5l8ibFFdt1rRzwi5Sc0D509LU
I+REWKJMkofzYgN5mFX9nw==
//pragma protect end_data_block
//pragma protect digest_block
RPkUUVv40JwJf5VC25b430iLbd8=
//pragma protect end_digest_block
//pragma protect end_protected

`endif

