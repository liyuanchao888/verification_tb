
`ifndef GUARD_SVT_AHB_SLAVE_ACTIVE_COMMON_SV
`define GUARD_SVT_AHB_SLAVE_ACTIVE_COMMON_SV

typedef class svt_ahb_slave;

/** @cond PRIVATE */
// Note:
// This macro makes sure that hrdata is not driven beyond cfg.data_width.
//vcs_lic_vip_protect
  `protected
MM?+1FBc#@C70;3^5-/BEW0/E0+N_[,X59MZO)W>[Y0XF.)?6K+.5(Q+TZV3M4E:
X4(V,CO_+H]XKASH<D)QfOZ/NGY(GHWX<^MD\1\3FJ6]UBB2>\1]L^3T9c-[_dS7
FYT;71I:.@KbQ;R7H5Ga):A\2W#cD0_4+a)fAe>4+-6#&M3CE]C\D0@g@@AU2]/?
#GgdRg^3A<GEPN0K[a8.2;=3+E<W;0<+=Ma-[](RD[3(T&D\F_2P4]BW;c3HE1IR
K0dUa2e?#&OUBZ2)B?4O940Id6KYL3R,OE3RJ1QP8N1?3aFY?g(;@XOY3YdQT@/f
TC)V?U]NBB8bOBB815cd:bNg^/K+B07F_c;RS^L?,JM:(XOdER:4cfNXc652(Nc4
?dL+=Gbc,<XNG_(G[[ZCV@Yb.T\94;+VL2)ceQ+bgXT8]:\-V.MdJ&:J^3KBR<(DU$
`endprotected
  
 
/**
 * Defines the AHB slave active common code, implemented as a shell assistant
 * which basically just converts requests into VIP Model requests.
 */
class svt_ahb_slave_active_common#(type DRIVER_MP = virtual svt_ahb_slave_if.svt_ahb_slave_modport,
                                   type MONITOR_MP = virtual svt_ahb_slave_if.svt_ahb_monitor_modport,
                                   type DEBUG_MP = virtual svt_ahb_slave_if.svt_ahb_debug_modport)
  extends svt_ahb_slave_common#(MONITOR_MP, DEBUG_MP);


//vcs_lic_vip_protect
  `protected
#&3^bL^FVa^gHBQVYXC4-_LRgM:(6F6RbG)@9R5]QdAb610M)=\N7(BgLA2BcL(e
9>I?\V9GY78E133L-8Z7YcWQI2451Z8eO2#/TgJ)3MS4bHJ0D@@U#<)3;IS[B#d<
3GaJa1<_>Q0IM)G2eMB)8JFV&[9;MKeXNPG@e,E,9bHd7AICJ^G4^<[_(33KH<)E
E><KB3Ub-b1>MKW#CHKVLW)^cFKT+.&;5Y)(TR&<QT@+=c+IHR6CO0^7SM)-3M5V
PXZ)3-@[.E_BOS3WYL,2-JIKO#MHL=7SQC.;=7W;[8F94PN<R5>9-2gCHd1e[f36
BcIHFM=8GMG.gOY\U9R46>L^DGd;\&H?NP++V#^]66ba,<,AaE&Se29DYH?AEY[T
b+ZcRW510IF(YSMB(Z>\)4Q-B<LE).PV@(/:\-7)UAaAPM([[:B^-B;V]+7O31CW
XDVY)83^;-.T=Q:1d9g;O_HGaI>1C6_RQ-T)EX1Z1&?+\FHXSN0XDZ;>E>/)aT;,
EFbBB1\T2f&HNQ<E;U]/69.:H;Q]be)^BP]b^R@O4J(\-<WbQ,WZa)<##eZ^SY](
CC/Z61.;)?+1TV_&J>RQ:\M_D7#XV:U1K3NYC@ZfPOI15)?MJH\VC>_\UHRKg(01
Je&+aO.KT1?W)Q9B9dPgN^ANQ9-HXNG_:4O3N\],>QHfd/RLD-b,9<5EY[+\^/O9
-X]#K.KN,.Y)V1VcBf:e,(8+&M3H<\[1+Nfg8aHCYKDa[LE^T?&+cZ304P08.VZY
b?0XS4W#R@\:U7&U\3^_B?f]>I?fY2G4.EHf(4DRY^(e&cFf,Y(IEbPg:KLOe;67
#LdDLXQc5SD-Y;P_dT_b2Ie1]IC^].PZ;[Q[J)F?ZYRC9#f7=JdO_EFcF[d17=a^
_1=(#/;BaRPDS.:JMIVM8SZ_>.WF@F@f<JAFGEND4KV.CY7V<fU>G3aMBN/?M#Wa
)EW<7DG2\8OcGAS@C.E0QSE7gIVK2DF)_Z>RHM;a9@g4]d^,]@X1e:#V;^&b=6A+
@aJ5f)Mc]9#&[c3c1Ge>RXAC/bW8CVD2INO@E;Z_5f;WWY,I&SLeLBZWG&B-:)^U
Z)>?=MC<HWfbUa1,/DAMF=E<?Q+#1+K3>C6DI\Ff-MLP98&3XKA^?M@:f(;79-#4
Z8=F;V_)YYJ<76G/a2e-?XX,cbH<NK0(]5:5YDM9C4XAW<TBJ/F?@,?+U]SZYX0X
^PG^X_C8VLYPHMV[gH3d.Qb3OIRF2CQefd_[\0fW70OK^QK0L9\:HB\V[YJf#Z[O
W_O[N8/D.;]_bI]_NGQL#6CUY6#]SP)US+9GPAM0UIY3HdCGI7NbLV3^eQO+MC([
QbP].?5[R(g7L31f8DH3K7PXJf[@Xc1G-W[d8Y>=D[4#[A[/F:M,_[WREX/g1fF:
7EKR&+I<MTE_.M[N(PfC.Y0\b)5RE;8W&e<Y-BMcM7P+Re1=TU7QSLRF)N?+6EI:
D,eY\=ed8TZ+X>I0=aZF8CX&8a[@.>AU9KGAFb)8#)F&a2Ue(2N&YN)TMNMB:/8e
0:Q+V]cY_O(bSP^DZ&YFA5O,J>]+BbF\E3EBNN<Cb4XFEV=TT,LU,aM&QH\(9YKS
a=#=WSd:Uc#3S@1T-A-I+IZ]6<be_4Y@Le8?>&DE5dXDCGT2L;_<U?&G:1\BZ7EQ
>-W&[&8C[02MZ9-^36X#=DA#DW/aAf5JC#V3;Vc;:Q\eSW#-Dg/[KDOXM1@[J@2B
]<KLRFcH#J,^T9/Ge-CVJ/WX#+X<TZHQW\4=F7BeAIf.X#R69:.;==8.=V)\#HFR
L9Q/@94H[?ZQEObWXU#N+0cQXGV6UgW:(N3eaAc129[]K-_=1FZCZ)U+:S<0Pg8H
K9Pc<c7=LDL4<-MbfbDIdIPMIJ7,N:gF-BLB+.gHOKHe;dQSb/3W&1;=BG<H@SMT
Z&89fTB;7<\Wd[BB_FM63ZMfEKA_;:cX,L8d&A&UXe?L6:?7Y;O#)4(,QY<g.P?1
J/1^;\=]c?+9KZ6-eTBNB3QW(=6eK@IAUb_7IB3I0[@DSRWeg;GfJ0=Q#fY[:<aD
,9YB(gR^[^_76^X2>eQ:dgZ4\[5(.+:Uf23\LAE?I&^#NP.0c)5RL2)BC\)5_O.Q
Y3,(TK96OW#5gg7G0X9I=,X&OB@JVTR/_UQ[c@L+_g[/&PD@J.LQVR==(59Nd;N#
bZ35[4W;N/]44dOg1;5BI_,L#.3c_?3/#8GE\=a5bfL0\Q1TJV^>K+]GIAa,CK3\
@4^9Q6PC0:PYZZ[J.6Q0K)5X((5>FXV^I<Q)YXbWc&[.f+GcH+2JIcO[IgW2&K)T
#?44\__X-Z&/9/cJ=L7PX;gOA/N57bC+E]UF/a4?)e^#<&G[EK\8Q52bJFQ;fN92
P^H(2-GA3:Z6D1_?0M^ZfU5HV0E)1b0W[Qf>+T(](T3-Sa1XL3=)P3Z)c6)Z(.9,
eK:4Z3LP2JI0&=J:0gU#J?1:+9gZa-,Q7O+]I1a4-#)V)Z\X_;f=?6BC3AS#_-&.
\_T=1F&Je:aQ4^5bOAG_J\T>Oc5Zg[7M[4-f#/@NH:7X/[KXTI,7V+XBCU)Vcg[<
9WfRGA.>;F+)N<KX+>^-T=H#A@ZcEY8#T1/8(7L)cdYU#Z90#3U>&:Te#YXO,A=e
P.?P=e6OcbIcV<CGbJ;d2=>c^)c1<;^WHeRE(AY>#7MD>HU0&>#@(g9R/JUP9(ga
ZT7186QfJ+K<6:5db([Sc^f08XbOI;2TUY#,683WR(.&LSCUO>,PZCLLMIQ++_I<
GFBB^NS--;M)PTcGWFG_R9U+O0I5N9CbcD#ecD,0G=[Vc\>dKUL5,McUO-W&\<U4
I;7cCPD=B9XQXLQM70E92:MVU<BbUU2]6&B<U4g].+^cG<3dA]N[SWJ79R\>+&XP
F9[f5350R][;3b]5MV_A+Ug();&;@\[<0C8G&\^0dBTN8_YAQKS5;RY9@I\M2R_b
4A,;U?:4aPg)6b9E9)G.[<#b0Z(Za)FN+2):O2WC0^dDX6BND[(B2J70dA0DRQB4
O7QY.OEZ6MFS+LQ)ADe,Q_c8^59Ze0L[<&BI5N?)(SdH2Q-:.3Yg4G(HQFN4R\a>
@CVW3cF^F_LUAWZTZ&JVdK]]GR2/[8Y8\7f1(AKV:RYI[87HR7LU/?2AK\N^7<V?
?K(fS1</c++GgedPK).1SERg_aG6H[=5F9I6GKBIK;K_BA(>97?@+_g-[W,.=LXJ
13e#_.X(\.a,SNO?UH_d.[c@fE&3=N,,5^c/-&;PU0SW9AN&U7_ENT9gA@2G\D@C
]M6g/.CV=8\-?(84AT57bN8UWaGSR5K]237FP,@J+\S?5ZQCLGR=PS@>B_c@;_2T
JNA]1Ff4;eV=_LeJ[9+^8;-O4Z>8QC-SHFZ><aRfFfTQTHT,V:^53(;S&AcH]=Q[
_Y2J@3(=_Ac_\E0MY^Tf(gVJ,C(<cHI[<7=&+;d^L^4.._/Pee[.U;,=b97f6=6:
,0Z]-R\TW+#-W02@4CK-,ZC-97dZeP]6MBZ;ce<W+-aLXNBGMG._?&&#@>FVJT>Y
a(N&0=SHdF-H4b[99[Igb;Of_@EO=TAHf5?88XbMd:Bd\9>KD9#^c=+cGGbe[&6=
_RUOC1cF=05>)E_]_?9780>cK:EaW#P4Q<E7ABbV^ZL7^=.,=?gL5/W.M?_d<fZ^
@K#DFQeV4A5FO0(FW^(;PLfD@+cP2cVN61&VXeEgNN+&43-6-?027[G@fQ;7,cOZ
\(\7\-K=fD>fJ0G=S356g+\<<R]UDF.KPXc=acYAQ>-[Q2Q^b<.gSRTJ9TJA#E21
TO8>,6.J4^#=g,VOVT3I;YJ3,;,U@HF7JXe?TSdX/+Q-Db4?PAF:^eB&R&@FY(2C
g=_@P[29C-S\]TaGIe]SaCRaa2TK]HDX&f@D]45@O(;IEe9NZ>]49D)5[:\(A.FG
EHUK^0<MGJM10QH^\\RE.g78EcVbUWZ[44IK\J.QK&baU:NP])6>I]#-SSY0O;b/
d;SHg04.Y^OKc1ee0MgaOdaJ2d\c.7\Q]U3_U.(?#V_b2cPJD;T<NK>1e?^@1K.1
bMO.N-LZ6>F],UGfaOUM163;+R/:U[Ye>SHZQ5dbO-SB0KWAMS.7;S)FZdS^HC1=
9V?dARFdCe^^SRZ#;fJYXa0FU2e(7V.PVH&502,3T/MEK?:?P6gEAO4[KgH),>H7
P(I.E_=KUP]]?<7gPXe,S@3&4K1>GJR(BBPX#]B_5&:dQaB]f=\-H9]<(-B3g,K=
4f8(\aIS@CgV9O]XB#_,58X>20@/#56;8A2V6bBa,eX\cVg/:EM@)K^ZG\]g^VVP
T/,_9JKDY81?3<[T&Q--5U5W1G0d5EgbXcHSEBb4YBc]Q;RB/\[Q+PNfRAQ,(eL0
c\C[Ld46==:APS@#3;R=/3gL3f;)N0;0/a>T:aH8&a63<dY>GXK/@TRKMQLERV^U
#NU,QdQ7YO4J+J?g<2QK>LJ/HZS4TB<ZA,NHQ+874[4?PK;SWdcDQG#11U?JC3Q9
E?Ta<K&T2Y#0/NM9R=RV;ON&NI_5I-9EV;8g<e(2M;C),L#J,bR4HF7JY[FSd8VQ
C)Tb8OD]T&Z7eT57ebYSe3<Q[)(PYKN=UC=EgIXSc.,31LLD6^_7@ECSYH+K:\ed
,9;HU.cfNFIM0c1=a=g4f(d;a(&1&CVc7VCR\U]9]1Zbd3FE\c5,gAV[MXKVX#D=
1=U;GeI-KI4-_9aS;P0ZTD0;\:+2bd11NZ\BRZ@[F>[&J/[.4?5=WaV[J$
`endprotected

endclass : svt_ahb_slave_active_common
/** @endcond */

`protected
81GGK@&[#76FF93R@-02dEAJ16,JfLWc#L0.DeS-DbUQJ3)]\))D4)7APV<H-#Z#
APeRe(?2---/K+JCH<+Z:EJ/(D?4L8YPT10]-b_Q_;UV5T6CX[]K>9JTPfYX&e\J
2+\beL8/3Hc2:]<51-Qb[H^EQNU6N5#T@RUX>QPXc=DO>QC:(?0:KC2.NQ#d9L/:
GPU9;L[Y(=W2[-B5c?64<NMF)[Ofe1&[2Tc>Q;>/5;[K=ZW&H[SMS.8O/M))_f5X
;=KU3_QG-41c1dT2JR[(@8J[(05d(X\0G;U7E+#FCLcbb^fH7B2#=ad@C97EP3J<
H6gRc/3_1QM0]SU3/\.[X]]5P6;&OKPN][KOJ@+1g&0:F15-C:a7/G2dR]e)IT2c
9+HPVJ8Og[W3VZ9P4AIWgU=T3-A?<g5P\DRGgdA4fQKIDfB)g^3:,e9_IN@QSUd]
?9M>f))HDUB<eE,/)F)c@;[PAK0\@-,)N1aJ[cLZDEd[/6N(I7YS[3VbHdF1V8-0
&]R(C1e]>U.&0bYA:R,BaZ1ZfZ.)I[0\DR/HVGCV5PE,e_g<GcP(OROJg/W2X9YV
/.F_0WUSRQD&/$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
,VfYB)f>I(,[=b,GZfe?;P.F_;SDLHWT2#EgD@<Z=83;S<_;I#W56(>D/0<A1GcF
39^HP3+&@9M\b;3+?C]3AT<YF+^3<O-EBdcU^PU-S9U-Rg4^I@IFNFS,Z+(@)SQT
TG6OI?27JMZ]3?=gb>8XU@+@[N9;GO[BV7+^X.?9F-GEeH\BSFOa2RdO[^U-JOIU
RQT1U7X3D3aZ0EO.O;S2:X8T./a+1V5@E(-<\#&.&YaMaFVI5?3[&;[g?b?2R-0)
6SgP@]+G+P_Q);>NQP]1Ae#L)KW5a\cUT:AH4Qf,CM\bb:9)J-._.g;ReKY8Yfg6
]Y9d,Q297L=67GA0a5d+J=Q-PddaQ@DJDHP#:1dY9-<4d_U3S\_c39R6e)O@#H_=
7f4KM>]KGb21LL+JfHZ5,B\IRA+&121[DDW>B[UD:bDT>.&g6Z8<WM.K5U#5.@b<
LWY5C5_#\eLG/#WY^0EI@.NB]MGGD[3(Z_cb6,H20N;fH2IZ>a4;J36P+VTVGGb,
S:fd/>@3-Z.)=YVJG4M<8c6],,2IW(CIW?PMKU8+b=/M.aG4IK69.[>E)a&2cCJg
:5-e.6G0\e;09&L(=&Q(+cHI,HLPRBUDARD/Y?]I+:OYQNCWY,)3XD<Uc8/V@;&E
R&:#TSFVTcC/R;0gVgU@/RBg>JJ=a?_g2?3EHEY)bL[+WF&GLXb66d;Ag.C_S5#+
gCZ4;b.Y?H=IK=5()#^988D:<f=:&[X1^e@WXR(XZG.2<fbH]GIRba2P2[dC75\^
1:]JE=OQ#WLZebJRH9f9?\>WgX#JY<XR2<X+O:O)[A]^ZBTWUJV:M3gB=JT0@O<)
gGWH7:[N8RcU8a^=4GaG-[d:9WAdAgH=B8A9FWB70PLSUWYe-K-L@:dZa5d?WDY=
g<M:>^I=AX70Y+=5HV&>JSd2O;4+0C/aOLK/#gf4#4]<E;VU(7YD[&5,YM?1g\V@
;850D=_A&49_/JWAS9/OO;b2_[\e<GT;]4G+DN+)G)-CSL^OfJMTTRWQ)(f.P#VQ
OdL#e=J56GE6#S1IdeUW/KSBB_)/XZQ.>FX]FX:<TRU^?ID4)[aT-=f[(@H</B?M
eTg3._(JZMX_)@P>cE8YB;b/6WD>AIRO:V);T2\Lf;,9_+bPE7^OGR8RCR8Y40J=
@fN]#SH/QgS0D+?9;^4X<FNSI8346U4(:MZGPM9_;cH9?IUg<LgP&J<:XP\e#[2Y
[26EH4)CQV0]Ra@AeS.FcFa+7:gOHHOYaAe0U+U@2LICN\gU?WXf0FFd3=#OKGMA
;VA7^@YQ\])\]O)173dFIUESMTQH[X3TC9dW4g1E[=dX?7bQ7a1H,cTD9Af\HB0J
(G@=AE=X@J=Tb;.FJ;/?VYUFII#8PL]Dc0WI?AVL&G:UM0E=AB0+O-ZYZ@\eeKg-
T4gU6PK#_VcdXJP8Q/G9M\K\UOO\LSaSZWdM]Xc&_.cXd@?1?ePBSZU@.M:&A?<^
:UcQLOT2?KM^eX4UY8LH18Hf<MGDIeOE46XY#gJSe2;P<)GD^A]&?2.e\f)XM?E>
a5<;#CaZ:8#]^TFKU+(QG_VLN4e@UFYS2b&BOVgS#[BcEUA)CJ&TYB#+0JeKV8+S
KdH0/KWDFC0Q)\1;O#1Q?\b.,LYf=1DO-(,+/;?QKE?_0_P;2K0A7B]=d492EQ.S
Rc@?5T>O;BQUZTJJ:LdRJ]RH&@?P584ebe#BQZ,OXgRQI2.D47N[(?1Pd.MPQUg]
.T0C6e?6(_Y/S?W3Z8=g]PA-/OWX_9@D@<)EbJW02<5<HKJ<AdCTQOgPT,W=B5HZ
J4GN)6b9dS&^KcNQ(UDeRD,DXHHX?PWV-YAK+0ZcK,8.:2<3IT.F^ITTX&a>]>J&
(YP&AgX1_W1aZSP=\&?bc0g#c4.dbb4Pa4)\>1K^GW1.F$
`endprotected

`protected
Z^;&X2SMM7=<b,ePA]4>LL@e&_7AK7aW-S(,M+GgXI[/XD?7#^]7/)eE=EZRIZ?)
\U6#A-UOeU?</$
`endprotected

//vcs_lic_vip_protect
  `protected
;TQ[\E5_C>Q/2b0NLaQ)X-:\W([T3IPQYe.C[N#XVOKXg)UFH&+]4(GLXR@5DREG
gG644bC_,)G850O-U;];.:J5)Cg?.UOR[E,W).4FW\H\6L0A4;&b0cF/1a4R2b&8
6^T4/QdeICg;ODCWf8PJ.IB<UP[H.FI6<IRGN@d2.;Ja6^,Z>c_U6H>g0dHPJ/X?
\21a7\H]Q8X<;@7E=C8ER6d+,fUPOO0+Mc^+-a[M6)-C)5L-@7fUSU[MFCDRQ[[.
DT<Y?21/6dX^7CKS<W82H(QN]e0:.Q7WH+caPQ7D+f&3Mc+YJgU&LcPIZb^C:Cea
7KW\Of)W^@;3UW(NF.BKXXZ(\F/+BZW49Rg1&EgIcd/20641d>AP&VU;8Tf@]7eC
,58].?^J5.,g=g,GKEa.,gZ31F(Bbb\2S^7f?[Z)#QK1:@U@8M2][7U9ALeB.R6&
+48RCBAAWRgSQE[:W6BC@f8FRcF0HLf_.[9M<0ECV@^ZZ5PM[B#g9&Da)(A,cfQC
[G60:XDW\CAG3\c@^05=Q8]F>^XaFZ4UgM3CM:1&C,CKa;SgKK)6;U,SKI:&b(Rc
b<&D4U>U@3Hd0Q@XH4f@78=-5]BD9g,]:1\B?RUQgg9=-].]d<K\Fg+-JWN:BQ\,
3H04a?a=2>[6UdPA-..X<3aO:,^VN:Q06_>RCdTYAGg+5N.0bT=X3N(<++A.0Yd5
HFa#f5<HKLJ]&08E+d8:P-K3856)0T(-9FZU+F]N/&MW.NbDFCZ4d@?I>64W-JTb
:e^DTW<(c8I4_/^4VVCPXI=5H=V(56BTTQCcg6MQ;MR#>QSXT@Sd^13)V]B:A)QZ
7>4HYCAJNaEXF-+:@7@0cO+[(WI,[1SN1Uf7X)G5DCZD4&KTP+5\f>[076G;_2^b
RUI(]H5gIN;D/)Ac<O&KX&/A_B#8HBO_E>f46=[PPLgaG.MBe3b88AY/T?aV<>g^
G/7-R,a=AUXe5&YO=W>1)8PXUL4#UT8g\LB2)F(K)B[;.?f?dPHR80IULMZg5?0d
Z93#C^>[FMVU?\H)[5#X0+FY0MB,FK0HN]@cX6)L=O.E6+LT@^[+LfVJ]+QD3B_S
KDF:;I?K4]N\R8/]6Q(X8HG#FcR@8>RT,gX8e<1MV>a9_RQ)=f#>(J&D@e3fJR_E
KYT0+_LeO[?aF;WU8WZ#G+W\eCUSN<ZNS9Q0.[D17MYU@T>2a==6=CMg_R=9::>/
Q\,)dS+C@3[3IMT?CA>]@.3X2aE^)WH^L03fg>>UHZOYFX^VCd5a4EWB.G&^X97f
B28I<;^8]f],>)N/Z6[WdM+.D,U4M\.g&,1)d4@#8^O-;-TY2dU1QKA_2+RdV8(3
dYYf>Va8WP&>D+XUQ.gRG5PULC,X1BQ^M09JEB8OWb->0V.UB1b5Z#EFG:PV(;bU
Q.e^g#PGfK7AFeaL&[8d44A8WeDWJU1YP0DEL/a#KF&:cX^O-E=(AUD5B-GYYFfO
L/2E=P9).^2/N:-]30MZEgUW\RI#I<(I@8(?NW[L+(?TXf4QOd0X]#WLIU4e]2Ia
2e:T:P)#T;\/3&680ECT#,JaHddUS_XQS^?/?CQ#J:=7_Eg)AfK8ZCUO:4RA3c2F
=XWB28@X)YH<[?Td)M>7;bWP=XZ&U6fHB\GSEb7#<]WTPJ__eXFgJdQ=#@<aF/5X
2UQ@Ce>R]4.HFUgTZ4GG>/ZF51/Cb=7U+W,]VU&6J(SL[Z0WS6B<KScV&ATOcK_;
>g,LK0cdP8fd?KIL&<V+aUU<JKB?2CPac7N^XZL#4V+IU=X,RC\OZg/Ta&4?/<LK
A3)&3#S:S64\_=YEJ,gZ2<C<92U[\PGEG.&CbGR]Nc<D;W3[^I(O<=YFZ.A+a;#(
0eK5cC#P>9.&#Oa=4Wd6Vd#A9;UXL_M48><<T^2:?RYL.N,,=c.61<F:;?@A.LO<
KHZ3bDQK:DR9G25<H_Z9c3b<HdO<.Nf@I.SfKEM99\ZCY_Dca,S?>V1Z?Da]6L,P
[@-F1K<Q4/N5\S1P,0I6POAO15BMX3SYTLOAV9d5aYbDQeGSEOc4FQaSe<9/6S?6
UPUEJ8bJ.3[f0/55=,(1VHML]a=TYXSEB551<^GaUF>,B@I41eSQ-1T&PT_IF-Ac
5HW5PFMdA-)SV1@\R&KK9^>:,ZWR;=D1>C37YGF:.RP.TaKF1CYg7&P2.TdFK<:T
NCAR0@L.)4VQ@f=TG.V[\;ZA(54[@C.5[SXU)d>fCQ-\\3.E&2A/>5B9SKBS<LK&
B_ZOPF5I[[cMK[51cYC1P&]&aJb-D-Y=#U>#LM#>KJXNK6CZE,0bV,?gW<B8YY[(
K35+5#^g#7fR@RO1TS_<H;;?GJZMc^(5@-)dQ>aJ(H0d4ID/2e<4+#1;5.>Bf@6M
)O?@S_HJ+)ARdObc#57P8:OX2#WSQU+J4.M.7/J020,[_7b2TUJS##B,\=XVg5>Y
QaQaA]-^gXe:C/6WMEO[9+^&>0W//@dKdUeD&OP/WX)&G0AVM8cgRVAgKLP^]>4d
+P:I,fK6&26=A3\a##c.ILPK3K[;5B+OG2CcD9ADW?RL4JLJVI7R/=U1Y70H6X\]
7GV_FFf)4(d@5Y:_JO(N9F@&,9e.#QV<9d\<KBJ)19:_TJeUQ&NRFEEB=W5dO)d[
/I)?-9KcC69,=X3\8TVD.K5ADd]EX(G?<JOfQ>Z+S2;J7fJSCbKDWFbDOKMMb(&@
Ie]Ke^0S2A]NP350c5]IFcb3J#7#<OF&:7X+J&J[_I[_6_/CcNHg<OEC]b2Sb(^>
:#acJ_V/)/XQD5_<#1<JI4^7&Z+\&X\EQ(gSX-g+RfKF0U.M&_gXc+E&bYI5:,>M
#cGFQdD+PaOHIU,(-I9ZaAU(7\LN:g64.^E-[?;]Q0#)(07\bAa6]F&gT_8I&O+_
EZ/GDYc4,A9)E67^MD>QA9D?KP>;97G+[gD8TZ\>P;6W10=B]2MD\,NJgcBg&^e<
>bKTC=-GKH5-W^K1_A4F0LQ7CAM+KaP#69IgfXFP8d4T/C4:(eIe>Z>-K60\dFaW
LJ;X7)=\E9[2a6B>T@XPfc0c95bg;9P46H4E\+[Te>0,d2_W^PR74g@B(AcCC5JT
1d7b9=E3febY;:F-:;/ZGX(B/XMUWEA-):/RQTLVdKaMXJYKA7=a-6^LE;A0D5(.
76GW=O2,U(#SC(9BDa1?QS^8/0LWF([9;T>aIB=-Of/gb+B.:X,fG(Fb4]F.YJDe
P0_c1cZD9GWQ;B-a&D^8D4JR;\6RGbcOF0geBC@_WK6A+7;SR>@VF\J:CXIKCJNM
gf<dDa>LTeUe+Ta&?c:,\KLEM8QAW;_8Ug+g]]C,bI2=d:Z\7\c/4V9-VAWO3.AY
T583UGE)+#0V+VMF4UWC&&4MHI4d9.5d;,g+KFJ_:,5f0:>1&.3OW4;Ub63Q),)e
SDVT=^dM)4,YGF:4fE3L-[H1F^D4_Q^B=N0)>PT,GKePV)QZZ&9>T2WA75g4964B
K+RWYPJX^T1,WFN2];7J=;]_Lf5_93c6RRS9AEgcYLT6.>>8T&CJ;;[8\e],I>#W
AV5WDFJB7EK)EO]99a-6a<CXUeSYcW<&-J3O^:5b2Sg6T5dIHdgU1?(\BSMLc/^J
ZgCS/9+BE_UYK,S)X2V.L8@AJVLf6UINQ/>a7?QGYQ:U>\2]8K>7/NIQPgC^^e(2
F.H1ZYHf3NO5G2\,P[He^82VN<2ZGa<cI))Bc-?9Uc]9DXMdIa-KP-&K]BXQ_a;M
8:WQ4SFFVK@1&UPJA6N@?O-0bNRIV66<>[6=_&\^GefTY^?HO,?cc6A9,9_+Dge<
OUP-b<9HLBN?aIg?<9]#/8PcUb;U-2_J_7D\ZDSWTVF1=7Y[;9GRPR?[D-XJFISG
XN1F28g2fF@>.OG+.DTU+<;E1H[M2&5;1:Ta>T58-C>YJHLNJ61^^W8Lb:U9:1NN
1HB)N>A,S?&6NYK4CPHb2c_#DP;)\Z]ITbdRe5:^.9M3.X&Z0GQ[-2Y0M=TTYZ<f
I7#dLf=]U&Wd;?1I]D#O:;_]4)B8(8D#8)HO0W@He9)e)7CXeKKAZbQgDALB8:Uf
_=Gd=0K-ZPC2TWC4HUf9K@]>4+AaeTB9>L1/fBFZaYE[-97KBGMMMGY4FD@D#c0-
cO893H;A=5=MD35bD\@b4(GB:<=(GMB)cXDgNId47GC74PF)U^&9Kd)<QSAUgT(1
Wa_N6K_^,R[\39P8I#8Rg.;#Y^4BFC9[NA@=b]ZPXV:b&]2NFce20G&=YAL1N-CR
H<M&g-HA3@E_5YOgRE=SL0P/0A[ISWagUTd6-RCZcG:PO28[e#+-)04VeG+R6THC
eUB=F@74(YWK[B77O(g,a25ZGC0eb6Bf3BF(TC1#/O;#bW_KS8.X_I#;(:&O];dI
H^TW>)1cddGgG^e9]Y1H&&1c>],(](F4BJ?-7be+(=5]cZFG)NZ+cO[-:/BC4fFc
;9A@3>54BQ,.bUc\cV^?M#CQ3^V1#OT202/\PG]B5X1X?6?PAE0eHRS<.VKXQ1^-
G;[@_PDD4Z93SSIM4F<[OeWHb&-84F8)A0<S5Z&c/)#@.RA7+JC=CEb)cZ7QT580
bR2PN]LB79#F]g#5#VNY1K>EEP?Z]OcD41X.=gO)Ab&1Y>0?6X>.ddX-@T,3f4@#
N8239,J\O1=&#YcZfA(\:M&>\VHRK8Ug3+QD0cgWK:g,?5=K&)R(g#?2V8EHcKZ,
4_^PS2CA7Dg8F/#A@8GJOXb#YVTG;]gTK7S^W20IJPF?3O.9CbV7F4JAWH?00g3d
/H?_9SgI9FWP?bP>AKPM1YPd(e::P1[_.ECI7_gV\KB3VbHUX?Te_^3aP(=AHT/Z
8gC[ZIE860);Kc)-J-+bd(C8):/,KXCb88SD4EGEfe;LPK+<;P_NA&Jc/P<KUWTR
]8]O54P]e/Q)6U->e1:3M(1R_KELM^-P0\PcQ(.c@Pc\]>;ObK.V&#e_&K/@4CQ9
AbT>SE;68eg:,be@S+6;gb78c\-b_5R(ELM[L3ggXF;)V]ULOGdY+0P5fNJAO<c:
Tgg-4^8H@>ZL;C(CeOXd4YD#?V>ITa<EDWQc3J\E-)bOFUWD@^D@41(dD7e65)XX
KUGU-P959HNJfZRVA;>EN,>X]WKMcJ\0cNGRP:/KI0>#=M)1GTP@R0#A(:W1gRCf
gM[N,O,WD^LS<d=Hf<MP?.GIJ,(Y<RHO-:,OV/3<d^Ca57NJ,#:3>[L4/)@6=V22
HC)R4eO(80U\V=#bO[9\f:3GK/[G///K2GPc)AHAHffbK0Z06.WA(HHJ5+0F+,&g
=[cdI5=T_g)f#8GKKR6U6Z><W?7ONO@&YT>LM>Y]L2.]9L_TFS#c;6CWGPW)A;ZW
K]d.3R]daS:XE(3bIU-93K=c4g/1MAPO(S>0N2KVeN<cSR#IZ/=6f&ZRL([e@DW;
WHPea#?NT6(_DFO7XVM_IOcP2P7Ed5+:_6g7]EO.D?1eCG].MQ+JRP8eCNR-</b2
^9d9DR2JM2]JQaQ3MCedg<T8MZbB7bBcQ3PWPEJKLYL0MH:B.M@.3UE..7?C9919
V&Od>;:[d)Z]BEDBM]<F6,_3b62Y]L.X5RAWFa<3440aM;1a2-&3fCBDLHI+Z:C(
f;]:4NVVUFUVJ1+H1.Y&d29MB=JBLADROCb\FSd)#[,gESHH-AH[^__QZ/_V<0Wa
gA8[Z(DW\EVNAY\/6<@.F4d#T;ATN79O(FaUdM<4)+]@<:>IaEQ<U@VL/O8W1Pc_
5PWCeS/K5HN/6R,gUV\BAQ0B8Gd&TFKY4UaRgB?)-F0E8#R?CVN:/XCd6[0X/,B+
e\CXa_U3^a_(9T\S,/C.AbS=fZ8?DUY8A9713?RaCb82I\be_6^GDES-XCAAE)&2
b?Ib3C@F?V[KE@:,L<NMO&LQ,#@6?^2DHdMP=+aLF.Y(B[VP=\cMK;FW)0A@ZGdC
</dZICP<P8E<,>_@f8L50Bf4-DaY1GcdHAeLQ^Y\T/;\Da6eCR_@eH15Z]1c1e:I
5eU/KJY/S5LOTB&KNN:#OG4&;S\HE/J([;9Vd:E@@C@\A6=Rc.Yf@.0QXcA._WKQ
-SYDG9,6H?KGb2GZD9V4&Aff1=d51_@VWCN2UHXV&:aN7S-X=ZBB??EAdgfIfLMI
RTV6VMF<LSZ[;;D:(PCQ1F6H(S/V,.)QTDGe-B4AE>#6&RC_gP@7CAOD>LWgV^)G
&YSd>J^eB76G<(BfGM,Ne,XdZ(+CYDd50,^[D,F&E,aZcU(]I<LJDP=,2GWab7Ze
[bX(DFOd#)MK\FaVFDEb&0A;^;S&+=#Xa6L=FRKcM#K(0eC67@Gcee/=2F),^,26
9DF1Z@gb\d)dGEDD#(/,3;QcO3YF5?+7FJN9?SBD0g0UGC,1BfgbB+g9R_R.)@R\
N&GgdVf&Z6BTaJcUFgD_b[_AHOBTSX6W0[=aL+JC7]TI#</J7Q\d,<=S[ad.B;b.
,)W@/,5-H5-XOWDFf-95dI50\1NR18LB>B#AJ5^ME#-3BTTQEAMYD/:Z=GMJ^=P9
=)HU3)Ac5JQ[0:VI[FILb^>OD>MQ:fd6;+#_f@b?2YOUefHHZ/EZM5^3+NZ:&LbC
\PeXOI#gVcT,]@LH3E9cN/Q0[F9;&.TD7V8f\2d)ER<8V-XUDSPc;X>045+a^NZ>
2QORB^@S\.+5].[2S@K)U048gb[\&YZJ([dP<Ce2I4(#JJK4b;)(B(I;IgH3SBgd
(8c,gY10C87,F;4+)#6V]&f-@+Z5LFJX57UM67fZK)#&^UL[6MW?8=?9=XJ-[S3,
\=-H/,:L+)9<P:,)1T[1f68cHcYEbD0<<WPV4&JQIKU6411Z.CS5=-D5@a.7?HJ(
>=L.U5GK(Z=YXb>NFX>4;[4?[46&IH<IDFe_^5B]&S4+9)+?B70)D2]a-#GG)UQ+
^g5E]C?@:85_XEIKY#MBf]0BBHF]&<>f-OB5+.5?7L1)@d2[Ge<5;N9)TITe-Z<\
XT)DBW^1M><A4@O]@4AgI;f[[8M-5P/G(ZV;gDL,P56MX2Q?ZWbKTRgIY80L30/_
decH2BaW59B1Z#&>;&QE@=C.TZ\0Qac[HG&YS2,6)4d.^dC=)FJ,)</2[8ZD.9VO
0QLU@Q<+=?>A:XWKXg0J@M&UR&#V[\,M@NgdeaO^FJNAO:6T:dK-Vd/U:AS=f>SP
AK1I\W)(/L.d6@DX2gQ-FN8FF^Fe0^:?_;.Hf4NYAU/@cNE./6>cAT#FLWYYFXG\
3UDF5Dd;3SI4I_G/?TU2WC@<47&5/dE5:,:ZeV/cd?F7HFYTU5/UV.d5eabV25@/
&-^[4\6GLAb;@YW9+eECN=]XT8F2T3bG[[&>DKUYg70E[[8BH&.A+0W])bM=Gb5=
::OD#^;8fKKAOg7F>\Sgc)ZW[D.Jb.:bW^II>XT)IE&g1=4Z./TF^2O./:M>KTZ8
NUF]Y\)9C&)5<H.gg8^U:\;8dFP,Y,XCZWFA<)I2MV:0?3#b>,EL-E47K>+304MH
aNAWNC099b[:2Waf.,3-3)c.X7N][ZA)<Q0/9gHLNU\(TZ>bD?QXEDXX3JG&^M:K
25)68Y0Q=,@ZY^FJ_8=TJN0(FTg]NP\X3ENLf0FK\YdLWOc]-N++P[7;&IS_<gFZ
[fO/dJV_HDFJb.0O:\,EI/ZLI7OfJRNTSRG,g-2XKI#(9fV[J<GdL>(MRGZTJ<PE
BTM4TTI#]ZF4C9cF-P=@MI#3LB^,(,]N=Q5&(/XJZG<7;RaeW)_6F@\+DI\F?M4U
VQ8O7cDM#QKDEL=.?6BE.DMQe:e\FV?4(G&@X7H1V0<_77fFc(<AgX@J]SS3NF#P
90D.4#><-1N9C&[3#)Q[6.7]^X,DLAP<_De2C0IOJ(?1W_eEYB&)d\YPdN86:Q:Q
4YIf_eGGYM<.)D,->LSR5A7Vg1]C]8&8D]#;/NSf]f,fP_/Q](:\aI\/+8DETX#J
R/UDI[DgF\AcI\f)Y44a\EaVY9-M?4Y#AW0#57-]7(dF_B8>BbD-P<R-..ARQ9V?
^b>ZW=_1Scc9&&bOX,3?>8#F/9,3M]67c9cQb][URb<7\7-bg6EEJOKPaFgA3])1
&;Sa(@WMUbVOX_FWR4fCIfAJXJQB(/,bD+Q&K+2fB_<#d_Xa[?F=:KY25;9;2&-U
[SK>JfOc/37de/1&A(SPN?af<WJJ=K:bCf\,Lg:^LU)W;TOd]b<6\+)N_Q/^_70b
M0/0A4OM[&AG[PYU5Z2&GEJ>WLUK(7YD??5&\REPQ2TARWb-.f6[fZI>#2XTPQcA
/;Da+Ag]9[Ze,]BX;2?A^&S>__-[d7Vf#[a<S+LLU16I[1F;^?2OPF<M/3?/WIa^
bNQCMfB:MIgLL,0),SONTfT\D30.\2YOQ;.Re)@Db/gbe-3#55];89W]gUKN/J[4
/>WB.cBY>dM,?.g[Q9,3E&<?<8=N05.DN=U:@g-7UD_+6Q>d:5GQ3QgZX,P-:TP7
:W,,7cA.e^5F_I6e-_5T:JBJ>4de1/GQC@a_FdS)#eYcg(CeSf@cKP>=O[--U^0Z
)&)cSW.[\[6&^1_XCA[1g.M[D>\J(2J[^.Ie?HSFV+0E742/C6-=:XO.3?c(M3O>
&PAD#=g>R6_I]32OYD;P_@<9OC&6^WaJ<S8+6Ic8>P:6J]LQAMg]?g4_:Y3=/M6?
-437dTP<_fcgTJH20@L=^7?49ELQ(^QQ98CG^3M)T#4CV-,]?RNJE;?Xa2@VYTOQ
0HO@#8Dda4Y<?^=P-fD/,)E<gU((]4#=SR#]MbI.32>^3b,=a,c9c5bX,2VISRPQ
\a)057.a<2U4,O=O@&=c=W/YW+3RQ?WU7+)LaQ\SbUD9<?8QCB&NZ,YKe+eITAS,
;UabIV+Q>I\cG,AC#C7:H2HIF1.Id?Cc;7S4KJf^c>S4D_fCW):1)W9KgZFS@Of,
#(I#>6b@YgOPDZN=gd9=WRgGe/-D9bP=f-c@O<:@:SWGM;E_7G.AE^50YDYcILR4
c@)=)[O9:9[]9fGUeXCe#)@]K_.EX47a#fZ9c:;9P?f?Le7+ILN(M;e;BEY06eM;
c,+_<K:VA.T#P^OO5G<7-GZN(M9FU7?E)?NRg]#S(5#WS5BPFIK+K-E&2Z+6Z6UX
FOL-87J7-a,aY/S9MHKW<=ZA_Ic)>(NY7IPb+8>S[LI4^#@Z0X5]a&(H,XS.K9B7
88E;:8O)\(ae#JAbDbZ&A@TebOHDgN@R@a@D>c_gKWM5M,YY55Z2.0+2S)06e)AZ
EgII]OTf3(C&;P@Wg7Q8],[Yae^XQC,D&VaIZg7a>=_O8XOD,).DUK981SMY4^,6
8K^BJfCf.HO/QC^7S.R;O>&5^]C(U>I7R\J9@E&b0VGSQQLES/<L8N<ENCJYLCTI
.8;ISP:+J1V1gR^WOb2ZILOJ@HJBd2WBe;I8H4O?VgA<85FYU<NZ:OaU)\Q,&E)J
WWKIVZYJOGYX3g[RfT?@A>#R0a?b^9=,NF92P/HI5&@2\1ER&P#R&Ga#V;M29de@
fZ+V]fZg-cESFC]@O[P]3_?gdWL?@gP[bRbBV:QX,WE<YX^1/4XB4>>M>W[WQX.,
WH>5]DLg):Y+#9g[BYP_gReX88)5HCWX@g)A@eC;e9V</:YR;3^EKPa\KPETU&SH
f978&3d714Rc_I6bETY<HZASgXO3dc67]J0L20#U:TQe2;53[T<.gWQ&I+RZNgR7
RSP.^,DP)W1D28#8SNI@3N_RBHea2X401&VK&A[E[<I)AE<?LPW7d0IF62c??5CM
DW1R+N8/aXE72Y-IUTS9T1&MUZ\D_3d,BLV=^..#4\K;e41(K[=?F6;45L:W:C:9
S)Gc7-Y++SY5T(g.5ZBGbSNQO>GN)B770BH1=3=+[e>KDA>e()CQ5VO.JJL9_Wg<
Q[\M(G:34,E=6)?LYPJ]>=&^?\fMC<5^d.c-BK0(Of[M_aa>7,PG_R(=;W]X_#+-
L@>0&<TTE:b28CM-2A[S6CC.1_P=c56g,)b493NPV\?U(I@?a/c.=b8WG^/[b1HA
Kg[]S-O,<LIEbEF[RR>Q^^_EO\U,X#;A)DgA5>;0.@@e#QDO;N]ca,)OfTKV@,f5
.BBI[,e:eL:-[++>UJ8S/.P>O9bELT\EOQ2B.KeXW(6(D+eASeD3Q]K4@7M_\]<:
85Md;P)T3PD<PK2]b#a;C?FKTdH8,Z3gKgSb.RI(-,31_)UHe7<9EAaM\HCE.Me6
-]V=H8[L[AUJI=^VE[Zd+YM697Z-3)=SN[4/P;6<37F58>:[(X)P/4(0Hc7<_SIX
SFB+SP&6X7O)6EBbT<LL&Xf1OQd4YPfb7[=gJQT:Y7FO[SIK2aWK35IbV]^]D2KS
?dZ0ZN_YBN/,K77eS&_EW#1ec30/A(G_b,M8fSPNZ,@7_e+33D0f^:R4O;MW8EOg
.S8H7)N8Q^b8_1DM7@;fg]_K)0;;a5>#cXcDOTOH-G+99:C-3-+2fP[;,DDc^(X-
6fO.6Qb=X9N4>YZV3YTWHN,=Z37/0cCeNTQ_HW-XGVWG7_RJ&E)9)4YF?);39Y6S
-=(FVXbZS0YJf?D_aY7@M5]d94OYf5d77SGU023c5B8HL0HSAQa5?>[84ab2)[/9
9Q^dMR,C8_J:G_gb^05ZZIO6U8:eB4Z)Z;OgdP8b;^<C+.:,\B\M/\Ta8b.PRSA8
\BE@C>:02UQ=JYbdJ]4\60e^9T6-B5GR=ESG8;36E9SPS8WV+.KM6bCDU\Mc52JL
0dB<-MdT4\UWgN=3)@./#ICdd;.8D+S;YDGG9.EgUEUKdg[TC3fG(IX&WF&1V^+I
][J.gc5CI=bXM_IEL88(#QQ&L[2##^S+,T6?E9[R)[bN#[>DfQ_:)5,J68#-_c-/
&B[2OQP:>U8)^Pf?];BA/+X=L([-#6/c9aQQXS7@c3A^BE0()6:G,:S&f0IZFU.Q
DXPT3cSaB^.[f)D/AD)RWVJ,KU-_>VZRU[<P^TQ^;4HYO.cHORCJW\?3A\13C-]T
1O-JXLAg4)#d?/T@[U54M+/[/,a8&1>3U1A(KW@V)H#(SgCd#9WZ\2>1<DIb(e^T
7DTM..FV0A@-ALYM+.SQ5Q2-gT,_?X(I0c/((T(1HJ<^<-B&>J2W&6+R;8O4U772
[Z;NaONC&-]FSMGJPPQgK[Ab>)EBNO\QD^,.Qa#\TS6L:]#^S)G:A,M,f?CM)K:[
A^E]PLT3^a&2B^XNU1Ka.(a35ScY#.DJJ:TdX?CGZ@W-E&1:5BOZa^/@XS]I5/L+
A/1P/L=1/<DP)S7+\Lca^,>-Zd_g++=Ie@O6Ff[0g>H>aJI&+KeYaG=M/VU#,;0X
UeX(g4?GE[@3]G4_0^#?3.;,HE;TY3N\==\;E^/?Xd\843K87P^cT#XVR?[SE@_F
af8:QAGNXNRcQ1#X/.2ZeZ[R/1GBACdLe[aA:>ad(/.PM?Jbb@?^O9-gH>f8+/1d
R.P,SF_9/35gce5GBW#<,55_#aBDg(YQGN-OE?TH=g_4g_A70WFH1L/K]6]]95#.
5[8ZM[1I2&3f/\H/Y+9<T5D-=R;QE87XA]PTSa;\WW/df1b:7J<>@<1L9C>]B/Z@
VL=L5^Jd<f@3N:Cc\4J1K1eGgU8AgK;HS5,gWX>V&ddK4:GE?Z600bRY^<#/0;c:
_LI;\83?D#f27(M;b-BI-8U6>G:_[X\&,>F(OX5MJ_#=<>GI&#(#e\4.gK?K+6gG
c^TQG+OEI5WdRLac;2I8BDPHcd2J@0JXDgN6&CZB;K1Fg3dCI@#g,6P&)(MZ,Y,R
@@S45S@dd40L@+_&M)^8QFOcBJFV<DWJacNdH<_1W^CU>UW_EO,dZ0,Mf2ROY7-b
J(IJ;7<@FJ.A2TYCa2PT<e4F3L3AZ.-::H]D6dJb>(E6J<<,eLU^B_+>,/4AXAV)
Rf21,7TC75d_5?,17P/ZF_>4VbF)QYPX?7AMgZ;RNQE#<-fFDT(gZO]X@DaW7C:Y
L=[([QH)K5LFRTG?V/_E2YTWPS]Pd;g;+^P3[U>A:N/?C7RJI^8Yd/0,@]I89PQ.
]TALgXO>VUdAgFa.A:eH;]-IFf:]H(3)-O>gFY)=>54=-d#&a>>57BW)V\G,Z70@
0PCMgI:C_8E4)b6\eZ(^5R1540S?)J10b.4UBQ>52\Xad<W1+B/\3BSVK&J>bC^@
=I6AJ>5[]FF-&Dc/R^TQ]&D.01f-VE)]U0dId_f[O]a2Tb@GZegA>0&fLga.EPI>
_1__)80NYL_1CPa35g?UHSFL8Z0O-H#ENJV^G<5GTEBD,E[OXG0Cg6E_H5+DBQ\E
1]_YCN7SBcWVg5JCP5P(g></([c=,1K:42d/_WVU=]NT;[=44^EFMG)U@U2fYbC(
FP3K\UVSTL_2)1RP5Ic\RQ04>Y#;B<E1dRB].L9eWH4dUT0/XVd/d@;]H43VLcGA
PQ3U+b)#L#=\MeK].eBX]+V0E;b;VSM;MGc0^[7aY^@HLg@=9X)BHK,-:9?YY/Y]
7ZfSY]b1dAWbFW1XJ\>CCd6)?9[#]+6?dbVP_/MV1&E_ZWF4J+7a3bM+B#@(WaJ3
S+.29=><Pa7U0;5[7LPF61CEc3E;aZ9fF>e;/b@Q&SSCg#,\4__Q=5>X=T@_6/-K
+a8c#&._TRU>cGJ38S9=UUWC-afD,\OJgXag\CTR]=&eG-J5AdD78BR.5>&<_]Y]
S;4Y#C@UE=+ZBT\W:)HY5Ke2Ye#,F<G#-?WZeE9&;2GPCB@326]2=VdQGLW]BYeR
+68?Kd(6UT;bM_:MO5d3#BN:L<3\6XLDH:O&WFSWXN46Kd85F0D?QOYUBBJW,?-2
F&N/-P_I\DK07G-(Y@bcK7@IbD#M5c,?N<g-^)Y&2X+^B#EG-BEgeT_edTD)\4cD
Y_FP@f_,MX-dY)7-g,]g:Cf4<U<A(9=7A9;S[=T?7N/:2NAV0H#&ECY>>\e4TNT\
YW-EJMS5bN^R)(d7Z^(E,]Y^2,#0J\UTdKN,9C:FSdF@g[W1A2SGVgCbBgaf=AC=
X-U3R0P05Wg2IO4#75^_JDBdV),4a[95GC.SP,.?Q16d+YDc-Y+IE[#OfT,86H\I
<TIc,LA9^/#c5.:e>f[^85]COV[E^bd)(<e3+0#6MS.6PRdONX[&)CIO;5O7fN.J
27LZCJ:4//6Lf:eKS@ZHO2f,<LV5ceE8T@I5UEB<LQUW<c)U[_89FL:E,bBWCTEQ
RO4]])^6-ALXE9X\V-Da8.BMO?2Vd@aHIR5HR1;FBdBB\\GT_W&TVP/?Q01=_E8.
dS)B@Hc>-90V8/^feYDe.;I+8GM92/Ac4aaKaMTX@gIV;dgD-/_ZTBW8GVLf+Fd:
((=C9H,NR-AR-ZN5^37J]RAX&^.&\T37ZCB.6K\X20I?E=S)FE5O#Kg\LeRJ<9.K
22LBLEUAVC>IQfZ[XE_N3]W\DQe4KBZ:)SI]AU8NS=g-B_:T>3__Q\_=AeeH&M6&
64.a#:A-&F7N/I.6XOE[f+YFA74.f7TYA0cNS8@fZT/J-4/gD@LaAMbC)3R;&Xa-
[VV1D?_6c)Lee[9162SR0JAX(,SQd>VG-57\6:QdI^aA:-#M>+f&Ec0H29:31:-0
&7F<ZF3M./eQ3>=5+C<C)1]@Ob\AHgd<C+\2;\1]e+).@b>:3PH547GBZ_\A?.8C
7]9T^:&D0W^B]33R)^MC4R4^>LF+#J.4KRf#XZ9ITg\0_XTM9[:^-M]KL/F4ZUgZ
6[#=UY/(2N.)AI7Z)?&?JW:\E1X2U(&^>&R6^SE8=YB,^+P>#:ggO:VB7F9e7LV+
9M@-BN1Ha<+-=R0bgK-F>Ta;1,2EMICIJ/C>[<^/bLKgLAgG)]N;SE_<)E0BHLB,
#)K3=+X7_1RBSde67ET]493b651A/4?LH[.g-bdTFVF)(XNL9b]@e;U9,,<g_+0L
c<6+_=4N[96FS-3C3d]MD1HcZ1;[7RX?:F-><BDK3PZK<P(&?/V)9KCBcEHQ4S^L
aZN&>IAJ]>VO<FHPg;3eN95)+>+PK<OU7=DM-b:F0aSBS7O8FT(Qd<#\Sf.U8ZP.
M+Ba:#G4IL<LN;?(9596a:UNLAQFaW+S#YC@W\?b,0U;Vf7PL9;U0FV-9O_ELf>C
+^+>#FGeddLKX_HF_@3R9)T-Cc=Q1AEJd(db;S7IDZ7.JGV9O;5QLECGH3L]b18M
C,OUZG=d<N3T@B[[7+L8/G7[T>86V7/fF.DI6_-=.:>:9=ALCK(TP=)\5L573WSI
aO&/@JEDQC<;5;g?V-1T.-;B7RKT7LNUGDQ:S=.E\T\c=K]S0\JK_AG#d.AY\9N8
EYM//D#feH/Ob>7=]\a#0;]/-\gO4X\LHC-[>HVA7;/Me@Od<(,3E:W8:Kb>62RW
fIKU4NJgFe+EU0VULS4HHDgK?Y@D5a=5]K7=.a3ZGQAALb/?QEG\bQ2OO(&@MMSP
]Na))3,M?5:,-M?1O#=SaC/OWdNbU\DZ1X8D6I;;:-gV:M=I?UQ\TQdG>)EVKJ0E
GECH)[STNO[4LCcceXAef/HBW/?KBRQb?f-\-#JNE<_8UgD+L^ULD,>:[S\.+IWY
:S&\_c24DJB,.DegCEgIHNUFN4@BLbBM(1D,&JXd):K]E<[V87<XN>f;D_B>ZGTJ
b\^1F(d6:UM;baaZd..Ded5Cc:CYG:BFgC#&\Dda;G)\;c2UN_KKRBKFNc1)ER\E
:\KA=0O2H8>b@JRO,cXF-3^0/dIN]-2\e7RdR/EDEMOK0\b/S7g&YLg>0&0K&[Y9
W[gNMG80K.S)&4b/]N&]WV/6gf?-PRL&(,T_-ABIMMK<40_gXaN\dDB<W=aSG@4(
HT0c2gIG2(>08c(;81<&,VMU?Uf-e[P<?AQ]EV\F;517LP6#5&Mg/@W,0Y?3Sf75
DUJ5@23c;I/O\I2UM+1X0+3-C[U&L39M\LC-&^1&34UP1Q<W8Z>;b>TM0)eBA;C9
;^QT&J0YX#3GU@4?.,0<7LOG2L31VbYFgVS9F[.fOS+:E.)^S?ZR-D(K91RH>4BG
QVUE@;gU47a028dZ\K/VE=9?J.]50FVT1IOXD9RP^d4QJF9/8,)e..6,e=\FgV2c
g.:63L(0NCZV:JfVAMGMgbWd5V0.&.07?<<EJ\@E]>Y+XGBaLUOa&O51-B(@HN8Y
_]NgAN<)\\=Y@^OSe/P8J&5^C1>O4IHE<>:B_f.TA_;RS.RN7d<YG@RACJD::>Gf
c8b^eWZJ_W0.6;07bf47@;;W_&eeP)G0f+U_3B\WdF)RW<7g28#W/1Hb6)B-3FJH
bO\]>K+2YAA@.RQ\UC>D^:dE<WRa;,7KfO)a/CLVW>9g,-]I.AMUgO)@?I_UKQ8&
::9gL<^+b=E:]1>E5;0[_Ad@5b=NTG)a<]5e[1QSGLIPLfb2KXdCWP>Jg(0gXXeD
UJc-d;IWQ:?39&)E(G/c43EbQO#)F3H2T+Jbg=1MKUd9=-,Q7(#=3A&H_3QaAZdf
2+97I8Q[]VK#76Gb2ZVP,(:b[3:\QbUHV7D6]>6TR2gC\_J7^e?,8EXX#-/3+PNU
#4N\Z?3M^L,[?T7I7gC0eSffS-0MDHWaTE1\][RY^.2TTJ2Pc.=]1N8Oe/(/PWQ?
&D+H2.Y5H,>-R1X6,O^2eZWVWAR^TX\#Z\<DJgS#dUNN.-+C0Y_gSfcgFWeMY&Y5
@M8YZ++>Fc6f)DKZ+YKJEZU]?DN8YB\/[FCLC+C,<IAa:TI1=/Z_:)^]Ge0BK,&[
3f&34ScVf68A3;VZ+&UE(N.(g]dbA>:<^OgOONT42:PSSLC4N;>O&&2Xge9;Rg&\
]/,fY+\fN9,2&a^/:H[MSAa,X47KdIU:M8\09+Z866d<SJHNFL<?e2Ig@ES4E45;
N]S51]H]?DG-_3BOQUFLSD\:6<3/)N\/^LgbY@Xd6A9Obg4U5)^X3=&Z][;bP,S@
9)2AG.:gPg+<#cA;KZB>M5,^S+T=fH?&?7b<F>I@)7B)<TJ[J3DDNePK5FgZ.,TT
PX;(a9e8,/UPIW;DfC,eT/M><g9CdRR33BO^?H8_R@[92YIPF/O98&eDHaVG0VF)
C#d4IId[=\@\4OCF].7Hd4DS[M&f)UVYT=1_G)M.Hd16bH[=O7d]1Q:CgPE#GB)C
LQMN<CWPP@34(;G_>,>P&aX?564fBd9Wd9DJ?T-5V;K0Ea2E#RLTC6>L[7;dA=[Z
IKXJ+8+X+;ERTP.FN8F5Q4d,G:CgI=.VgPKDg?#c7K9/^G^0G<O#YfI8>CA5T0OU
3F&D4,8VW_E#XS^<;WOE)aI,BDREE([B_BfT3Ag#L30,F2GG;NZ/QF5ITUM4?^34
B-=.f93]3@7I0QbBU>:;8(;Ib&JJMKaPd5\QIb[ReJM;N1SEI\&&00T.M)H(dd.,
9:c_N9aX+8Z/HTN6c>U<ff6bVN\3^WTN2#7;G_CLSbeE5V;B9Z0G]B(FB@G,>Q>F
0Za;QK^bLVH8V:.2+_E^^.8B^HWW[<0ZV#<-gEY<#JD10NBIeTU7/g8E4b\U[BeZ
VN3N.Z=.Yec0PP-.4C6&]EH@I_gg6_PBS2N-CO9/\OOHAfP,2ObBUM\,GER9XS-P
BQU(&,Y91))CY95YVTQ1AEL)T,,d[ATV?JK.J>E5dff2g&9X;35U9O9SW\6F]\d+
2RWH/6@>6,-d]d(\9724MYG8[O+,QA06Y\-fW#UWBYB_eOF<[,aVa=.Zda;<>:>F
/?bbK)H>A>]dH=M+XOD?aVbf[+/&^Kb0#(T-e0D__Tb;-;_=dg8CT;DZ.M;K@@(U
QUUZ:eB@IP[&12#C4+,,\0?0XcCf0]gDT,3X<_P@Z^?42Q:>?LU:5?2&0#R;_Q)6
b7[7+_1/GQaH^3N48QJ96K_X4[?c:7Q,Y^T#G<?,L=-g#/g@8KEN9IJB\]0^&6GL
KfR)2KJA)?3G=Z)VCRMKEB6A:&OeAM:?/HM\?BNF:@DE-D15NJ#P<X)N1c?Q4:>P
SeR-OAAAS?Q4V#_f/BTUdUCSB2beSCbGSQ2+-H]#A6+_a#<OPbC0dd:<\?gY[VU?
c;?H6,UZY@3B-gJ=HdYQJ=GVPU/c6-1a2)/(9>X)Zg\ZD:=ZO,C)A+Y9T,3cCFE9
GZT.J6cfNOd;Ye.34Jf6<D3Z2[Sd[966=5T<C\1V9DW102>NYe.O(N-8dV4(U&V;
,9@a>.T_edE<gKU5R[C&./222VJSPUdX@eOPUU38c)=7;>?+-SQdOa:d#QA4/bVT
)CMc&ATIJ9fNZ+\=f^L9[?\92F@c[B)4Z[(e1d0O:/ZQ/)&L+S@46(2^U5CC(e.2
VS.bY)7DZ_ERQ&.7??3:V_.Pc7bHKDaeN6>Sd<cgPKU)5K<Q9_<N6>YCT[a@49]S
bT=3fMbDG)<26&R7cNM&e08gQ1=WCVE.[U)8)X^D5DdG&-R0eaLF7^PQc5-#93NW
6cC1,14R07C=)5f\Y-5?fK6e,RZ&b>10,?0-:XTDaH4EJS,KbLC#/-2[F2^)SSK/
5Y51S^H/d](;=b_e7bN9]D=7#XaJV0O>2Ye64c_&;aINR>J.M1UKa3<VO<cI4R>\
8T11EgUOZDZT+?5ZZ)gEg\(@5ZAaWA^Y(,<#dPE2bf0F&EU_42H@,K5Z[87ZTV5;
3Uc6AQ\472FcC0Y#.a?37gPGU[Z[e[5\#_&73)O;b)8fV&6D2a:0I@D;W6(bD)4e
JZM/.NEKQB.HK87BDK+aIC0e</G6Qf7P2gcWEK)?g#21[660L>]4a-NTVI,C30-(
1=ED;9+U-ZUCCTc]:aD1(bX@N>?_L7[-7)<2L2.TS4=bQ7>W1_(:6D^,J(=8IAOa
VW&H0L7;\LDSUUO8&\N5gaVN(L32OSg6.)JJgU;@7B93LQ=NC((>CWa.+2SWUS1@
a.QO+NL>P5ZFQL49?;MEADG>@/Z&T750K3UC6d8R-5<:^M&ZgM-0YTZ]2E/O#[f7
V[Z)bRf?G[VGgJ9=>FgCMXC6ZYK2U(,9=E@eJDgEe]<O;e(-M.GLa9_:aKZ1C,9D
C0T5T\1@)&/#Pb,g#,??[L\Xbd[WR(X&GL-9?.>M]X>UZ]c[X9^aM&d,gALV1X#g
NGX=-J-<@Z9J4NB3](7_T:7Ud=G9/Oe_U/bP6&-2fYfeLYCPW=:IT-Hdf;3Z[D/C
aP2C-a/+dUWMEMZ(S(=dR)H02JW,VL@/P[&fZQF/Mg]YN/NY.R6G7?Z_0c@?VC:b
97bA]-VRR6M79D8aE\DI:.b/c1/c;LEcF^dCQ[N:7LZ.X1Zc9,MTZ=43YJAE;^&C
ec;[a/aBN;?&J:;.+Y8;dLIB60TF+WLaaBe11EN8AP&/X[VH,X]b-A::+4?6A(+.
19Fdd8G2S=I4X/ZG.agVM&LW95e/=K_+--=fQP+fD]X(QV8\3LJ>2X)EKRg@T7Q4
egCBH86N<C2EO6[1GCXHSDaU,BZ&cD\/33_5O0IKa0fTe5Q:P<W,D\+:W_7aFI5,
K[A>1O4c3N+QE]_I[VKZO:&UQ_<_AL.\+#a&_T@RUec)FV4)QV8g@.MWC7:@@T/0
=4^YXV/Y[cU__P6^c9I;W>H[9+=7e<X66:.FU-\L5]^#IKF;LBI/H.Y6OVFEgNU@
F=>:RKF[,2EB@9\^-__ZW]IZJNV^B+]JC?NEXJ@E+0N2G6;D<&M:55.SXIWL>agJ
\/C_LZ@@M1B_DS_CC,2e4R2]^P\gC_e57RWH^VDFK&EUbF-5&A0>>1V^U5R3HN<-
OGUI5Q#:U5F,W?;8W@#9>8cV77/1Kc(BQ_3AD<\Q(d2#8dcZfGK3YHT+Vd)Y#N8(
Q#01(C)D(Y04)gf)BNcG[K56)W:JK3BO<&O7M5+/eeG.=fB#YZRK3&\NK<cVKFgT
80XBW^:S:6[edaCEF(1+P@06]\D:[8)XH6(4KL0H\aMfT9&T+IMZ4:LMJ7=&H+3Q
1X@GL(OC<d9fJ9FMc6&103&b#FC[M6TK3LP>e;76=JVFe^SPT]-)eL9TX/)++-\_
WBVX2)eO@WCDZX.A/b9F\C9<-G4:>1-b:&,Q&L?BQaD<f\(B@Ta(I]6W\D_Z^ME;
+-6g-BABPOCPL8K[@6M3GfCb5M/)?S.2@WFfL6F[H<I/I4eN/MG@<+IcaOG#<0(+
f>YaZMZ#L_eZOGUWPO)@N1d[@V@LXH^^&>PB#I;aH\>BBICGb@E_M#3c?RT(e(A7
2)c<6&II1\KC2,0I-eg,C5&f5f\R8>^T&Xb&c]4.ffKA<KJ.Vf]U^U&&11)f1/A?
/1DUA=<[XXDX5W1,)GdUdR/bG9T&e@G6W+7@/(>eJ&QL87Se.Y;14P1&BIZW,M;Q
@Ve2&)LY>L59VEB(.NK)4S:V^A)MBNEJH>MB=](Q2c.(/B)8.66A46fVFa+YCXWc
JWIeD?(b\83(.EM9M5?(#32BIO2J#7]9b>ZKU/K4IW/dVI:4TO(I7MGZ(D/+UaYB
UVHI[@&WYUQ>ZDSgUBZ@O+PIR4>YE@(c0g@7N@?-G2?GFS^GA4WN)]W9U7FfHBHU
2J<J_RNUC,+_@?>99QI7gI>Oab^Q_HYKgF]E<Be_f6PfK-:A(6N&N]JPY+;\+KQ)
Z1b8:dGBX,7a,PeZ[P?W=>EGI)a;[OA&HY-FDdaBPS<,H3X=W\ERd/8;_fX5\G8=
C]FS^[bN+N1f2R8?@F7)?YcFQYVF+#:FT)a.]_<5DFXM4Y/E@\L(>Jc<4T<<=)<?
DM,b=a4?<-/TYZR_&V7dWT058<_VE_[OaJMAL[T57DQQ:[WdZ[<[?/=DRO.BFJK8
3MbgPe^Q^gOQ-V(eGd--Hf;C&]b1>:I^cI?XE43DC(])]<EZ<.Rc:)aD4GW(c74S
Mcfc&<NJ/,R4Z1:()Rd?LR[RZXEaLdS@L+;Y=f(9G1C6-e7X88O-)_.dZJB5X^A+
7^+&=R81T?)KPaW=U^]IXX\Z8G-HG&40Rf@FML1@f[ORFF[2.LVT#=J-f/ZR#d)b
:PU7T[Z+IVFD()\:3K8_]@)-MXe/0UZaN3>\9D(K?BWBbGfQbd;M6]I?WYU5P;3P
<&_f.B^L3MP_/c[[^]YW5A13&KZL-XG(J?QYH3[US@B?<R0+<J0<c,>.cSWUY7@/
M;.)_^:2Vd^DcK/38RgcHQKBU/0ILTLf,<80F5_Ua.&G1c0>;&MJ>&GfegXf])?O
I)^3)XW:LfAJ:P:?.M.P_gaOfH)8?.:ZJXZ2-SZ/JG9KB.K]<E91eGH,LA33)#76
cE?#)YPWe,7H_=4(4I#XMAA[Q0Ya(=@<YX,51FVg3aQ0JEVPA=[9[3d+EagFCZ:H
WFMCb+f>:R+&&1Ye+Q9N5,ONT,_L@5CNLUC.B4&:IbKMIDBa3NFfH2B;F6?A_)9O
Ge038A9(0S/TI@S7?X+L0c&Z-(K5:)C,#I?AIHL2N7X3+.ZR[6Q>](YYR2#HZ@&L
<:aTCXK0>Y^3LSaZbI)9_KT9fI@VcOA8Q.GZ:J;\7+9MYEJY0<82a)+P:+E_5)Fd
=Ydc?O3V-O+EWCJR/?,X75KP>7c?daJ=E6M_BY.Jg_A#=D[R/,1Lf#8C[(2G>2=_
2I82d):5E@HGZ>A6GSH3QBCdND@:GXY\XQ<B.aWR:Nd_BA+QNfaAF[/2MYKb&5cN
+)>,&3L0M@?4);dK\R[<.NRM6/NN@;2J[Xdc91#^PDaSB@P&gU,&RM-U:&F^A9R_
D5-Q>Y\Q.;(W1=#/F>#a7O(52]U5/2XW#Rg3_UbY:[];REOLUZa_bUaU>,OOV]+J
YI;NZA;9>]_SPU.#[3>NCRA[/3)KL.7)FT7dRN]3(.UI]XF-ea?(cKM)0TY;1V8R
#/DcaS.c2\74(&?[O_9JHM0<Ga&C-7\9?f81,1UH-Q.f?M2LZX7@6P6BVb_b8#=b
6(F5-d9+I-Y_g\.6Y7B10f3QMZ&3b_M-VU(+;R13<>AA2ZP#=/NOSIM<U/dQ19C+
]XD=C29)5)2HK=S0C@fUYIJ2D?>B__>GG[b7_2]KNUO1adLVd8BMG+?B]#UN8Y6W
@HBO:D5H3R8);=?5B++<^82gYQZ+#Sb.;L]>(2HG&<6X(ID.B4PDg,IQR@Z#WREL
P_H^WQT/T3/d#T)BBfVCHY2E3>]KVC2_@D7FJXHB_1[J92Y>NA;]MX9c<)FZ^gRS
:CeQ71a7]&\I\=IAOWRXc-_fe]2Y/W#G@5,C\R<3M4-?=SKSNXWc[B.2C1.1b(9T
e,4CXW6:<2]fYJ6PQUU[I7IL/P7LPSU0I460Dg3:+d3-0[WF66:-QX&?<^g])\#_
AP?Z?1MF9E)a:HC74?0A\WV\JRV3HJSNI>94SJ#=)e7c34EM?JUadad538Z]P^JG
]N_OCN,[4+\BcR353#0&+&fYEAfe\IZdI8U_?M#d,LSI-_bG,_);:\dB[7#3CE#]
YF-]2+Ff+];Q^W+=gI36cW)6HRcfLPa5SM>W<&[CBC)g+WKCNX]cAUOAc0KdA_]]
f][TRMO>3WOVDYL1\@R1X<8BNd#gZLP]N^Mg.6<OE3O;2JD>#+>.gT7U9N]YZ<Zg
T4Dc-_E8]L(\K:]a?O&=J81XAR3g#.NJP&H>@A)_4Zc,L[IEF1gXJ:Q7#ZJOfD0g
YF)b3/ZeP^,3RY;0HYDJQ5:J-4Me\DLDQJS[<L[;9:176F;6?;48MU9c<<b&444:
TG^b./CQ_QLgX>WV0Z?\F0b406JQ08_;TY]TRg+7@d?3^FGU2>]&@QJe,CJ=9aH6
O2.d+8K=GA/7>)SW#C0I6.J+&QG(O+Be2#=1.ZYENW3Z9gM83_NR[OPb5.88L:1b
&R\+cC-1#30b.GEFI<_S>(aO@^\YRU(-T;V8JMY8)[Q=;fLZ@adbHg[a1AdD[&We
Y/=DU9gD/]P0273G3a:GC,,V#UQ44T/E/X+;B8(^U<TPT^QZ,C\C>_+W<HMF+TA.
VW2_c:<2d@?21KR@K474HYg31#PVLBYI4C:a8@[\9/BA>7Hd3(K>E0H^/)C&-&5=
T6:QU;1a5T/>X1c2a,OgLT.V^BN+9d,RaT.,,/VQ#<-A5JeAM(/I-Kd=M:KGM32A
e-;-06,>:Y[#P7B]VC9E0fKDV-\I]1/U7Z[dFMbAH/A&>2/(1&:)V=.[Q,)0BX:H
MP[Y3NC]fF^]KF1If_Y]FK2.e8MVZ\EaY=6D:b\dQ6;5E6S\U4;RT?X<>1dV:=>N
L;WM#1OZ-I#:34b[[b,dW-9FaK@GGF(P[RB7RfS+F0cV\(eX5f6D>AM,Z,b&;IXO
&OK[E@+/2cb<0U[89T)134#b+.gC)@<g]TTfVO:6f<LAe]8Eb>7KA)Te]16Rf5=I
8.)E.HSE,72gd,1aOaB;IT-V8P>6<bY<6.@1?PZ1K?Zf:P7e,-;2geb2NIaCD9:<
Pa=6JGd05430;LNZ#-35bGGX/B9<b>W10(e;g3/Rf6eANQ>4?ef06H.N]J\3K6.H
8dL<W(ML9_cQE.W)acb/NP@QW#9,I:f.(-[c^BBV[5L:dJ76Q5)0dDa?4WFWf=Wa
@Y?AXP)YB?eT_(=VCHF)b=ZcdJe3W3[Xb-A8JD7:f]E)7(LY9(>d57C(bCG&XUHJ
SNG#.Hb^?;0Q.60PK\1=fY8<AKUW.,Vb9e;5X+7eQUf6MF9a#2RQB/02-Z#.N5?9
,]Df;DBCRJg\^EVV(N&/\GKJ\@)YJ1DbJ/2V+6,:F_g@1Z+#2][FKF+^1SX@)RgW
FQf8IN)H=6+=S;TQ_fJ]^)?Qcaf.2+_?C&=&,:@W362P==e1cdb_=A9NUbf]MEeK
>2G@]^.MaEO@X:fXRVA[+M+OeSQ[,P/7,+d)f#YD1LYUNAVc&cC-FV#K[Z^.IMJM
QAK+5Y.+Ra:?#RV@0MN^EM&-#2HC=??4XI=PAY#XY7X_0]Gf-+A<Vg<A]/Hb6^=X
\E@6c=e[&3X0gd/G^TFGc^T+:dH>0UN9BAKU5;/;.N^Ca5CDHc@)Ea=(+H2CJJ]F
>_?()T>R8eLOMAGR^0?<\9g@d)J8b(GVIdF+NIZc9R:5F:,RYgG;:RVZ.ec=5^Z9
Ha6(d72bS4RM7)U4U,JT]VOW@TR&9,/)edY(H+06PMeF/.H3M=O8/07PC6-T^OAP
ddK-(L]DE15AXHM+d.08XS0-@07gGW-)RSb_3M8[NbR.ZJ#@9G/PN/V)Q59Z-5OI
=2GO_?LI7a+XKH/-ROO?@^IIT:=g_,f,91BL7ed>EWR9LC-;)g9Xc<F.UQR+);]Y
5e5b,-YW72?<Ud#O3Kg]cfa-OCeZdaC5GIc8QGJKVZFLb(6?EGDf-d0YZQ+A:#Ud
d;9L3)(IX<Y.g[(/eKK\H@&?BLMQM49RGHHOQVFf8A/6&3aIF9C0=fZ.;O]JK=8G
AM0=M4;f>6g-JV/(-6bY&O2S1<X:\GWR#BXW6DSQOHF0G[6fD#CR9FZB#D28\0,?
J\JUMe>_\Z[)^3P71DHfHLJVfG+<1N).:3V^(W_]1;dUSe02)U7Z&A+.Y\2.Q>Z7
17=<=7:SG^-6G6H1OIGYWA=g08Y@]E?acae@-B7+^Hf=D?#6Yd2&=G2-f+/R[MH^
=NL>M>5R0)AFW(<7QTM7(g@S0YbMSRS:dT2+=9>;G34[f1F8/CK1B=M>0#eBJ#TM
d@+f:#>,C6>E3DVd-R\&46PG#-W[NUWfWfDQSARWXD@A@[Tg[0^;1(1:EJ\8(IA7
CQ4W/6.MHUQ_CN,F2Fc[1PXJ;9W1TF57W/RJVEL[a/--T972@TXTcfcZaP_7VZ\D
W1/f8C/+.F-AIA_bCM,8W4JE3(__U#g^=DO4KFU)1/Nd@QNTTA/d(Q_N@-&g-]B)
L#<TN7H:>feMSLOXWB6+BF/LGEHKYf_f+Y=Z+H&f2.aA?>V.DGZL+82C2L8\Z_b&
cTH6Z?/DOR>ZN9M347I:bCGM)[>0JeELVN;UE[:E;6HC91[^,_)6Jc(@Y8LZ?PD]
-:4aV,;TLZ^,ZF\T8>\09XNN9\T55fd/IL:KfM1?6;eac1^HadW5TE[KAO>[7-g]
=AgYI/LX@+[[d0=X1-VWAUg8+\^SC<9/6J0PU52@OF^CCdc-#CfY50Y<R.SXaO4I
]4JY(g(dL@dT>6P^MD-A[dF@F@_X=MNNGT#@4<-1Tdbc5dU\<HM^a1H5/0e>;K/K
>T6Q8SGJgDE&a?Z-^V0J<=KY/J77YB1;S?Z?Y8C\ZB929__0B]MAM8e/.]>I0LC8
He9Q=21<Y).;@[Y=?Qa7:/>&6&[U:g/YK9+W,Vg:P+9BQ&U[F?_.e4X\XUI,_EWF
&.YTQPO<dZg&OUSN;SaCT5N3(&.Ib0,cFQV]IY^DXA7TS&+.]4DYUJ9+M,:MDJC+
-A5J^[;Q2WTRd+-P@#3eS^F_3GQ(W?M3?[6C^3f5>3feZ]P?[IBQ<P;&gWe;#&.5
^FUIeUVK3V3#SX(\=[6P8T\-3XbZ7g3AK_7g7SEE[2XG7QCeZXZB8ZY5d5LJJ1^e
NO&Q\_TOIe_;0b:,7CX,fI674Ic-814^>&,^>E5SIQg.PN1J:9GN9GX,#8=_[;MU
R&V#JY<4R,O6GgVfd8SPZEN[?:g/5U=@Ue]Y6LPLS[_ZK01C(^aL+JUXSN#TE)?]
_@+.-8b/BIc4&bFKfcG_eYcJd^811d4OX7A/S6:Zb-HRe1\6f:Fe19;@9NfF.0cP
LE:cMWWL[R6/+NH8G)TG3XI,G_eT00Ac#TP>&dI947g+d\QA.)eJ>W7@cA>gVU#T
c/GGQ]g3#N6Z<V32Xc;e,5/01)RV@M7/]]4@R<)(66[g)\^5eI0RGePTV#]W)FGf
0+V\..95XW6PJX)OY4Ia)M/[,_ROHaf(D3bGO1?TfYOM1H?Fa,-)ENI9cMeSLDN]
d.9]258(1Ta+=(b=MfFE\+.BbK^)AK-5]\OK8V:YWfS[XZK]]3bf1eT[V;(@Eg/]
gZ5^;JZaZQ9R[L<f(J_<gIMP?.W(S1e<=0df8C.16LBP]:\F3Tb\dS)3Q6McaMIZ
?3QfX9;5-e,NJG>3#[P2PgV&96T96&4;BQZRGPTb\D\<_1XSGLfWgK2)Xf/2]QJ/
A]\(d#G0HgXd=HZ1R^=GB3L)8]MX@a<W^@T@X-/XFTW+M[M#-JOL_3T^T:F)<_S&
2.U&EI(49]S9/X-,cDB.L8&Qc^A_0B?UcRB/GVQ-NVTJ5-9b)aY6K0-KZ;gGZ\U;
d,d69]FS&TE=QBFV.=FF;RY9[P-?<LL7e?ERZ0e1(I2LDE=O24&47K2XO7G3VTED
@N/0ddcTET+R^,O62NEI:aK8G=I8K0K[0/U1S;Q_>9=5e2UMfe+//9OL)8NeVSHf
Xg;UN.fNgOQF^[D4_+Z6/8NU1A]\[AD(YZBJW#FR/d;<+F:;^H(10PF0/\<,<F8G
;S.dJG-WPMMQ23T;NGGO,5H8QTGCOb;NG=M5GW6>Kc=6K:W1/d_X480\DI_dM9\)
T^0N#?@J1<TF_P<[ae96G:<BT:_aI2QVcS4&^PHRGG&V-;9B]+G;E&K7,1)(?:8[
ZN-QX/;[+[7R#Qa14;NJCaAg@;_J+<c3<<TP0aG[?gS/-LRd7KN_MNLX+D02M>aA
LXP4XO9U5K1=/)ZO\V0+#HQCMBP5HXN<9ONL+BZI(,++5+a<=@N;^g;.,,N0Qd2a
C\;e2AaBSAdd(VYJ,3ULYf1A(g)W?b@X\#.<CY:F>^Cd2VJ++>3ZU_(X890aSTX,
MgQ0=C[;ZQGA).A5gB2MS1FFcF_T>;+Z#g;A95PDD#bfJ]Va&8K<8A)YgF>40<&Q
V?57A(54&1b+7SgdgP22ZZ\+fMM\R?C=SI2IDL[0&Ka@f9R<08CJWbJOB7^W6X@^
AY<K,.;gS=#+G+QO&\g,ZBaO5)+e_#Sc/DDA3b/#,(I#^g#fX3Y&6C8D/bQ:@DZ-
XGcZD,\?:@0&#4KX7]1g;_WbZ/G1]D?WT&=dCYV7W9+9U?-HKSSLPUA_ZfE&T@KJ
8eTdQ>2L/C4OLVX,EeFBH7IWg@5)_(^.;D9aRC>AWF)cfH4GHUJH:9ZX<+C(#>S?
8@^G(0c/4]TY0>C?R:(62_MbeY#1E30DW+1Te21<IG/EVD=?[DQ>&M0I9;MUXC>5
QMCQPfUXg-0_&bRORO?A\Fc#]#gg5M;<JLE(6:7YN]+Hac,Q3K2feS?O\@S7(ITG
)D:,G.EJ21==,JUa5,\c(WP<[:O2JN)?2V-Y1A:3FI#^_\DL>9R)3eSHH&U>VBc<
V>81[4)T?=3P\aMQNH)#9(M40SfMM?>48cL^NH=:3VE(R;d><dF4,/B3d3R7&)+2
U:d@VRfQXbZ1+AU5fS\RGYEWaN7X_SB<HIK>CNSO:],#20+TNMBPA,=Fbf_]KY@+
QD,M?VR5P#9ZZ_Q\H8S-DU4:Q\+B]^aK&8AXd=&NA&Z>c7-KOA5#1G+_V@dU/eM8
[6@-#VDU9KbD:eAWEJ-C?J@,I?,Y>A/T#.+#3RdZ).,5^a?]4G7H=CYbC7ZAd)GI
T-10(Z@d^g-GV&)M1DHF/YY8C]1VBU(J>LD?^6PBVTBEB1eA(f_cBc[I60+9SM8Q
CV>)cW&^)BH1(J-g8[@6>3@_91/>Y)S>Ye.X^^J4=[OZJ]HZX[<OT+KCgC=IZC[I
[RFgCSZ/0?S/WH)\A2Me_I3Y5PNIFTH2>4]0<<#]J5T?4.DRc2,TQEJ1]1D7<Q9J
JA2Ze4@d4^9Q+_O7WMNBXJ<5<V++K#8\,[Afg&=0JPIJ9N[gR:SX1>G9E>1Z0LX^
48QVS320cR8Z9C7[c).7?Cg^V(cP_FIN_DSOV_?3.4C0XgSX\[F2XNC/Cf5afC#b
JM>&YLIK8Q\MZFB<?TJ=IE&Dd[PY@DT:D&54G@I;;N7,DNO87W/KSbV#_fOU@RWZ
G<G#\)@H#b4;7K(V)Za1aWX&?QcPg1,BD.WLJ?C-<2d6OZ&?d]^DKVC?DS/\\]_f
c4)J)\]3.QP>97(F:[Y/F@U#1cN9bWdS:,BgP>-&0W:F#EE]UgT_K(B6W?8R1g/I
_G<&D9>E7F3)cX\\@.eYa=TV;:Hc:,N=cG?8?G3I7\1>d:E9SO]dHR=^LFJ0AKaF
_GEC&@8\&#>2F5.GR-<bfa\fX_2.M+DBfYV5J8ZAd/]L59(V;7JYVdK@F7F3W@9I
6/0-&N6HgEVR)D+EeMVTBg2KL0H(/05^:[-#F(NA\PRe;O2A04+N5<9^1C\4U.JJ
G,R+XZ=4eG9/MUP4J>7ZKY<AaXP+825daZDDH1?II5[1IL.?LU#\,Q^ANG:N=_9\
[:0[YA#Z<Q\9]?-NgWePS?CY;I2)5c\402[eMLNY]ODGIGg4LCaV4(#aD/HcZ][1
VfP;VCPM=M3<;+H.L93YJe#:FKMEQW;_2&\(Kf:#/8aE0Y]L=>7PH7@VC;U-P/fC
1:K_agF&eK(aEJ(IB<d>9PO-\#SVP4_5K]\]V@^Q?<Y]PFQb-fI@#d_5bL64G]>N
+KC)[e4PYH75:0MB]I777N<:A<Jb9EO@M+8,:FLT^S_1@c0^\#N9-Ub35FHLN?NL
>J/O4_^HGEQ6Sg#V)cJD?DeU\D@\(c,TU002&Q<g2)<Pf620bUZ5Q<?&-,.,<Z_Y
HB(R9gE?@^QP2DI]>/-Q4NdX/>Pf5>TEPP?4<dK<=T2O:^aG1T[N:3&dfJZ?(=9_
d+a._d#cTYWd5a0=bJRU?Ie[VJI/_J:PRHb9;L9=WC6E_5c9MJM\\BLUZBQ>E&/M
9T]?6F:?N,G9YI:#R5DK8B43I,.IL.f]=BfF-V5817@#4V\:DgfIO[9C#[3UT^,\
g5.A7QgP4)A>[.[d-4O9HO7^KAP4+?YJ6H8.3WKHd8#XdZ.FPP_WdZB&bCbHK4)<
D&6/&PcS#39<2/ZCE/XNYd38#eYGMX7Qf6CSH;;;(_B>Q/76Ea<#\B+G806\CSW?
Z8K8UMDC4fU-NT+8Da]/8g)+]]O<RO(\9<7VIW5+4_+1Fc8Ec6a9HKJde;)X?#KT
5;3c523<XTf)U>JEYN>F3/)]BORASB-WWg,2+=-]JRcMIb9S0=,-CHZIRP8Q4ab<
[ee.D]c\9@\ScU,Q;<[P9H68Sg(cF[\gD=.+8[=,PBB^X:KJJM@DIM2DLC_UHE+D
J^PaMQ=SGLHKb+N\U5fC9LBBdK-6dQb_1P&eLN@@:@0#S]6.dH=;fb)BG>8f5X=]
ZYgg\>8914,Bdb#_?9A#C2T9c_\SSa>-J[8f)&TeALMG8f@#ACHX;[6bXS21\U#,
eb^7_47fXS(dJT@Y\T;X4SJ75N7-bIX>dLH-STGc.&aOTV(3?FCbN9@R,R9-(Ca5
[(WL6OcW\adQI6Wa=K^B,?C74FbeSd:d.T)CJ:M@7d0RA4&M2XX+&cVH8#P:ZI8V
V2YD)a&^:=-X@FL^6,.TP9T&B63dc\[fc0+Z[UUag09/)C;SYSH#A55(#;[6HL7\
0OPM+Y2b\K(_+8>X/6]8T<\PAVI7dbV6>c#+FZX\_R\#U:Wg0Y_)=EAG#=,BSX^<
6&deGE,13g0OX1gEQF5gN+(HDZ#XBB,?WP:[XP.3Ma>U12I1a6&>,V]R7VfQN4eJ
W<c]L8MfA[WJ[)K8KF#3414O.bK<QR;(K<&<>bO>a,HY7d9_G#GeY\8DL24;G3H/
IeaO4aCNB[R8XZ]E\>B](AWZ]1/KV3?L3GHcQf.ZBa4[Of&0SL+dF7KVN\_493&Y
QY13E>dV9>VZ9+YFU/H8cHC1\C5&_N82X,BBQ7GJPc_OB<:\>P@OK3a82ARR]55O
IYU22/[<9bLY8FK#H&G#cJMV-a)[M[-c8(Q1WKVMBWaR]:&VI=<=4?S<.d]3c<;f
A2H)]a22bLO1@B]\.7J,QFOT1C/_gMUR#,4Z/7R62X4bc,b=H[QfB=Y&HPPJR5QN
dXe+5PG)<FKY&b)?A&;GE,BZAe<JR2bN[,-)+DEL]6]aSI;Bd.+:71XYIf;T/]+>
LP[a.1QRPR#5S9>E)87/G;]4VNZHSKb@O[.C,SY5;AIAD?XW7H1-CW1.F7_\Df,7
?-1N#V_K&fIH40-GaSbE69cU-)[FA\/X6f->:1e=DN[6QMKM3VF4&43DaC.E6.8c
>g\7W1V\(R<8-LTF?b.,f(Q69@/?OX0EYU=BU<55&3VD0(\FVIZYI[VV/IAd((HN
LG,CUD7;=RQN)Y;I-U]aL.&YK^DW1bW\#5dVKC&96)70PN#DY;785Y2IK#E_S(4Q
A8d^&05K<(0.^39C>bT\PgD[(V;,2F)DP0R3W2)M0Xg]c.(f:D9I<-:)(@U#]0QH
?d_WS0E_g5,dW<\;5DfGJ#Q7]3NPb=E,MD=L4M-;b8DIcHfSg,CP3]W.0,E2TUSB
P]MR2<&J27;;=3&8J>P@?feJSO7>:>2b8:(C[M>[NRa#MdMe<Wb]a:#FR,;2NJ)4
ZKeYTQ4=X#6:P/&.)1RDD2Dg_TI4H5&IGPdfd\0f]b43DFH,8/4[1@(LQP>YGSF1
8DY;f?7D2fY[_]:9WdJEF94>Z9N3Z:C1UL@)a[gZHZF&;.#+M&2M.4Q9<^[ME(DN
9,KO2M[B[(B6eTSHQgbMeL0@R3JYN&dK_10f3X&I<8))=SYf66)G6/4]BdJQR7gZ
[c<XQC&Z,]6I5?P/UK4Y7VOLPe#TX01-dDg0+>_Y01,]d5NB&dHFYNM^be2M7b4/
5BPV-GI<=SHg[#=.H&,\<+</BW)EH?B<QEPg5=+1;=c[-@Ka7#8>(dV&cKF<c3JL
0gM[WVJ[,PdFQ,PWV=\KM?AbWCBCUEG@K(17?SL,Tb#d2d:_I7[ZFL+IeM#^g++e
;[IcV>4\,g@.NT:RcUP,07:Y?e]fOSIAJW7W9EVe#ER)ZX-Db45.A2>=e0]1._:,
LC-0>O1:_2#LBGca4IO8L:]O-BYE/7FDOD\(&]2?670dBU)6KUOTTGf0R;:R#@X+
4._(Z3III]7=3.9d0f+_^Jf,WSc[f#5._;0@.2RfE1D[4QGT-[0b/\N5<_&VVK(&
GeB9CZ]O6GeG8>5GP<UfRH\[YgD7QGJBG0D2N1[62@e9ObBR\LRW8EMIJIFVI?Lc
4?g,X]#4McB^//:X&cGR70L?4KQLDaM(<OcZKRH7;1&AVN=<+?gS=KS5G?U:V<^\
RSUV?eU.RI;PVc-Z-G?J-Lb4/=6Y43RN/#[A3eA5CB3g6X5+aLA6\SD5_/9@&XA)
P,U&2/HHfN2DF50(U<N7#NA;_Ja>1ZNd<A/CQ4XR?3JF8C#6S(A&H9f2ERZ#-31:
5If0#IKS^T4T-U?N+L8_YXHJ/]A;/D_D_R2_McCKHgI8>P\MGVa;A]TXH_#WG[=C
>,];B:+XJ-Pc04S[+_BVLF4U,-YdCIMC54+,Y_-T6,5;Wge.QD4gaZ0CKa6SMPJ\
ZK=TF.=.GR]Dd0aKJ1#eNef93[XC\c(b.1SO_7P/WVNgL#&GbIG7bAc2fZ(1?PM^
KHcQC^N&b<U[bP/&)A?925+dXX@RPV,BS5W[5/C)E9AGGfW/ICAV38\]3&13PDKQ
1S(7YL0_bdS-.8\2FfLN;2W_8-d-GF]9dFWULY[T;4baNYYS(TTRWe3:+S)BZB9R
(,=cd\=ba+\0A8:5C&HPC?G?5R?XH;gHLfa=G;Yb548EGS9c^D4.-&-d>=/\A2D/
PG?SL/&W:aWURM8;[]1Y<<a>IfScK0<=T459].@9/CO8XC?F?Y84^d,eA<Saf<A5
-)=[1UK>RAa[+Zg,-0N&UV+aQ]d>F)1O/+@b\PF7^Ibb#E+OKZ0[Q5F-#IQ0I4P3
S@,<UcRF6\)HFE/:3IJ)gE5EKC,ZbE(8VK)3=O(/PHDU;E/N-9QT&;/9)KJa?cWf
0UNc=fO]A\c1[840P7/Z;M]E\5DJG3BBOcTXRb?Y,C8XI9T/H4,NJCJbABeQ6A\Z
d#cS[T9X.HQ[-PLPDN9K+)ED/Obf0cH[C6_>.7\T43?-ZY7a[F2Ue/aS^V<G[GX7
B_\4LH2MIDLOSVN<:Sae=<dN8<Me\fU>Nd._A(@[G8.?Z&M@)H9CE;;Y0K?;+R:f
53O)RDDg:RHK7gOgGIHJ84-KU8#PdDa]<@+1b6AQ^_a1@bMfMWeXPA.?M>HQ+GB[
S^Z&(N3K>eTT[fa@c?X5_TTd&04bHa1D?bOYBa,&BM.Z3L_?J?3WNeKfA4.D2,4]
G@2FL-c[+4NQB=9A9]\9G9E]9ATbOIQ@[2;8T&d-QHOKc=Ied5T-16R.JSbb]I\R
5=ZWZg@g=/B_KIgTTRG8fI9]Ne9=bXTbP,HR5^,()I8@XKGGRG7@NYb(O.([NM.H
(\5GVIZDYOFPYDK#(3BIa@H>aOV)NRN&>/W1=O=&OH_>_1L3@2FLTU?2K#RDO\NH
?4\HB@0PKC@=DNTEfQGbfP>1U32>Qe<5@RL-B/eGO\T<:7^M_M.JA\M58D^U#BQ<
B?O+8&:[,WS+gQR&@0\_24^AcWa>.,9:2GI\<6#FI_(BRdS<d(&[Q(g4WL\,A.6<
VHLOE(71Uf1SaY0IYJY7XD3YaB]BCd8>8cU-R2Ig#8,B7Tf94>FCM]&^/</d2);C
5PQB_3D]eO0eLZ7E-[FYWL^;ZfXY[MPG&4=UP84b5,/Mb_AgF.;T)e\6L=)IX^<3
^DBH25VF#+>_BW6^<P.70b0DZR:aQ-X=N,F&T]C,:5Ea(,78.)0XVOW5B:KTRSEW
PZH:VTWF6AE6F(97U<F1X^[=-?JQ;BZ>)?WF3(4c<OI7Zc0PcE.?YT7>f?aAc6MA
6JF_V0>+J>3KB,gGYN[AH,[=7$
`endprotected

`protected
gP9a5B;YVOSfg6H]2g/D?ce2-;cXQWg79:ROCG<+>eO8+D8HOAeQ/)e_;bcf1?^c
HEP7@=00YS1_3_C=(\HL6O3;_=),Wb#(?$
`endprotected


//vcs_lic_vip_protect
  `protected
4Z4^R4edEKIFI,PY:/LJcNYF.,_56Cc1W:],S84b,4G42aEJ0WKG4(DR3-K51O2f
[-YWA2X9Pg&^K)TgHH[gMWW<LEc6&OR^.1PHfg5^.[d/+,5YTSg:SO\576E^OR?C
+1=[]]#Z=ge:79U,B5N(0+V4CbJ#BWW6O3>Tf^E,CTO#0,^)[G\&2:48T>]&Oed/
d?[21(g&5?,E=D+g_WCP=B.T;\f=+fd<]Jc4AK7OKZ,e-?^dSLOUW_ELA:a1?].&
L>I6]QX<ceS9:ZV)&#b[#IHZ2PEZg.W=^JgN]\6]S:\+V7IRU=60\EJ2\VM&2#,J
L/>B.M4Y.S(f8fB<;O]N)P[=>UNGfaCQ&[b3gI]?4Z06;K;L5T+-GG@_[]g<&QE)
<8=L8b6I)GPd)gR7/HL.bPTAe0WG1fH<[=;gB@BMP++<X<0RT&3M7N(&.\V)gd>;
XSV4bU7=])P)@S?:(e+fc&QXS6\>c._ER<):Y2G<B:UIL7Q/7dVF7/#0f(2+A,bZ
fCH#.ceb=I&KfcB2-/HV546=eI[/ILF:C3SaY.fBdB.:a>Y/\8:VTW^Pf?/_JcU8
f9&P(I7W6YQd3CVC_7X2G-bM#5Qe-U&BU0dc/C9Q4F8cD;Z[F]NdJ@gcP=FZ._WR
.H,4;Z_4U0^X+e2_==d81GG)Cd+G-e;/,[@;(W8<)T;fOV5\63R219+\g?aBE@XU
RMbW-J&ZgG,.9(>(&)?]-VP[VRGW\)9+f<:e81OB0^KL#F)CSWKDJ&\42\XO6WU,
eBR.21ScN+&&C2)1@2^&,4>>Q6;69,J2d\//_?#\^Qe:PLM.WPJe-e[1>Y5D+F&5
6UaVPb0c,0ZCEM(Q<F:[KEH,#Z<]Z#M-J95OI-bQbZPA@a@edJWB7-NRD93];f=V
98e[8RB7R4cL37J:/:<gGNQYL1)V3Web:(cba4Q;&L96)UM,0Q#V:b,KIS&ebB>S
:KV#2GNXM(-^RHJdId8f&L)B3_JLW@>5ESFNLFJ@[a-CHZ;AC6L,I4_Rd&J\(HVQ
#[&Bf+VgaF(UGII+W>;8a1bV>DcHEZQVL;2,c\0JNIAXWXO#1;gB6:Y7[cR5O_\8
+^X/7)#BYC&]8B0IPM)+0+/YEY&RJ8>(/&7#O;O(9^):/;7RE(?>\R4).5EJ6L-T
ZY/52fC822XR=H7:I)L&>5V^-aZNGUeB)VLgHT+VJEeIL#Q=@9TdI:F);?F3aF9@
+@9#_;FQUGK&ORVJVX(@9N,IAWJ63K_SFV-QBL/Q_>^IZM:cVK&<S64LITNNLOe5
dVXOd:J2IW#a.-6#9H1M=Z\97\13)O#0dL>R@2Lb2Rc:]Jde:_I[Y[S(IA5&0QD+
8=.(M7eIE@Y;PgfQ5(T\(-;OKGE0g/ME(2;KFee726)XEPKP/,GMYW19[,Q(WgJ@
S,QK6#M:Zg3TE.WX@WF&]11[c9da1N5JP6Y1LaQeH+-KA\?>;9),D^6<-?C7b:A=
E2U7\52aJG=94g,--4^?dKQ,f:[CWRPFILSFRd(MRWW<Y?_H1Z?3C<g<VY]_ZH@O
3S;6(JZKeC]F7#4SQNQ:+,ZO0G\IS-3P4;=;&/TScAdBLXHYUA.PT]2dM=f?+_EW
NQ,b_0T3;?Q39\KgVO^M,H)W\FF],cRBVAUCB[2e@eA;Qe;>5L+ARD(<49/;c5>N
(2.N@<#K=JZ7:fc750ER]Qbd&Ic6XaK;)U2<02f<FA^C#_ZX&Z;I]_JDW)<ZPeg4
]/Q^EZ=9_6We)b_O]MODT7O9LdAVcY.(QPa>TXN,,5G/MK-@F;A+,30McCC28ceN
1;(WRYUJ6\.8CLRF[69_;8G.EONCEB4(O?\4?/>b6PgPSb7[>ZWc3W7>FPH0F<OY
VLK<9B,3AfeG998\P;D<g9ZPT0EN8;e#c3ONf#d<;bNDbMIge?6W<8@dCG8fXJ95
/dW]I&Bc((F2ZI^<f&>:K@R,_e]OfO,gU@NQ(>-JP_W9&0AeEe<EX:V+gJIY8@?_
EeZW?^f>D_BS+4P>fe0/9LVH=]UC<<)Z.>cEb&_G=TbgAXW&SK>]80?cWD/)Vg6S
^V;QM0BG-L1dda5J5,U::BO^c1Ad+B.L;dCW=F8QN-eN=SBE[;+a)\>G<ZB2AJ_S
2_-7LO_<X1,Wd[/J45Pa[M#D[+aBgALN@G[6.?Og5WK1GA0P8#3TMcR(PE_Jf5&,
_,0;2#/F\6#>?4BR4L1I/\.5^2JM:MB9VPfJWT/I2(aP[;K/;IMU20R0/c<)IW.Q
/TLg[eYJ0NA=Q?d;6a>7T&e3a:]9(>aI8_CH2O;,9dO>GG+(U<&=P#-^/BCQ[7G7
.gO1AR(F4GLQ5;S+R9OBE5B/.(C3U_JB;8\A:2e(#dgY,Y[eXD5?[g]87DIOJ@/[
&g5d8<PJI3_10[WKHR3<P0;#LM8XRc,1V2W,=53R?#[g>Lc;.caB_0&(K&,T\B&D
FaWeF:<b[/T+EU(,\VXZCQT]>a.++B)]adWQ-Z-OE-@O?G?9-DS<gW/dC=XLN-TK
<).Wf+@6F9BEOeeT4e@J/\6RdEZIaUF;9&>5c,A-T(:;XSFP\</0H0FE[7.5E-Da
TIecIb+=ES]FGD-38=9:DI5_^#gKa_0JJ\=8BbGYR]E^;^JNFXS1^P?;DCYa.5YE
06H)2F4S+)7K(fQ&W]&##0G_5d+=?)L7a2db5^/J[/2:1P.:_3/XW6b57O+55cS<
7_&HKcYG1<?g2;-9-S+IV/CD?UZ.A9TbTR^S<+6>04W(c8_LM2N595^8a14SR4K?
#CG@N^C6F3,WA2./&:TNd^_L0X1f3_4MaP5f>>:44>0f#H.C<-+Jde236cF6U7(g
8+24^0W<EeW-gT(,DZ1TKZJQ<-,?8?M8,NE:IX;JH/g-5U8.3M@G//fg4_cJbTeQ
7+17GU8P)0_<+KaPV\aK2A1ea(eE+U3^-C50AFZ[&\BJ;I4)D=3Nc<03We1@8T,F
Y(Pe5LBB7\(L?9DCaH8T-<,<+1NgBY_NP8-eXB0Fa?2\SF6ZH5R7O@FTO1/I.dfd
d=dIC]S8TCX:Mf,-#@0Nbg@eJC8>@Z].(E<(1EZ,;Bgd#@dCAHK/NK@;eYJSQ_db
G205V?C#0]-;O0EgX[6&gY)BcJLN<OCCT67BGU-dILRT9+>38Ze&8_>]5YWDc1G4
?d-AHV2Wa3?<=O&7-Bbf>+CJ8]=O_.P;]=_^?D^-O.#Lf/S;HfA@E_/>c/LbL,&X
41T=+W<2=bH(AQ4QW)gc1Z:Y6dG/]<HS=00GCOKA7(/\5ZJ]XYX&e^O6^(NH5B#U
35&148Qd2CaefO-[<[CdTP2Vd5g#5KJ:KLF-N\@>L.-MdG0Ec<A)fCE.^c34--L1
@^M-.B7=JMc99J4N=Cf.?W<+J@D-C6>.^e_+;Q?NfZN,2bTR/L[3J.HNQVcFHZa1
:cQ.bGf,IHS_,)QYU.Q1b@)@\:L+AQ0739^6f_F(MLUX2+fN1/]?]Q#6Z>>3BIdM
fAeJE0bB8;5T;e>Ic/KE,;Fe?bFR?>E^P>c_#H;bcEaCN4OfE_8SNd=5]P5^0VgL
=:>#^O<ZX71N+<:Ba)SYF1N[1U9\M.ZgBZ29_+9G,?&:^MRF)&0YGU;S\IQ8]P#O
U0A=;>>I-#7^gQH?-7V(XTF\?3H_-GBBFI9cZ1g3Me@_??WZ(::dL2T8G\Z#Gb]^
_IA=2T;]C@]>=(_@gedZ?2;O3<=cW5V96GJORfN4NfVN#P)<6-(WTBJTNd0MFGJB
NfJ4_-2cHS,X5A_/B1fHNc^V3?@8VV7XZQI?)d;[+Q;E7@c3J.P;+?LN8+:4KB:K
cJJDI>gF.DFeJ&Y\Z_a)FJTN5VPG[>I/&RO\-:NSB60XbXBH^8[QVR97#HLO/O\Z
g4]P4dFfH[JcQfFdb2K9,E]XL5VB6a#FA#gC#W+e>61GT&<Ie18Cb<WV69O7R\N:
d=3>;A&ND6S]NBXgJ](e]56ce?[Wc1><.aV3+ZQLB]83>4QV-dg0GfL5ZD=XYA08
6T/,>KecW@FNUU7+Ha>Og6I@MULN7Lf?8_;(44@=OebG=B8DGDG[--=H1+-#)]RB
.8OYLUTffRQDQ:V1^bX(=8JAA&#c4b;<_,YYI(F?9[>23Z-Hg=Z4RgM_K4EbU,7K
+gN-/a>/&bZ&cBL1T><RbJV6K2MSTTCFP+F-H_)CSS/V4PM,ESf6REUGB+>)T<S,
E0K#SeGUPX)Y8L4]aFeU&W]X4V2?;ZWB&AA@->,0Sd[,7GZ\1T/EQ)IF696]#OJe
Z_RR-8Jb]H1-g;(XLD.R&]37c5?,5UEf4(]SM-DJ2E@gYAEeR;<VZNG43&5>/FG8
;?W=PNf@NRU)J2#eI]N)f0c6&15G3S]Mc9FKV9B?1Z2:PJVBMB^2Z<7a;>#.<E]:
1LKM,<>?=#Ad,N^+R7=I30;fMN/=Q4WMga5]1c:R1]3ZR<UX-L/=Lg)Ac,CL<,1\
Ve7b0MX,W>T8LeT_\<_9g.<Q\[a>?e;R2ddc19IV]D_\]gX:(8QR?@VDDc?I<Z1+
2818)R4@YIS+gO6d6B?fD80GHB>[Kc7/=\[c>LH^I3<dZe0RB===VY4BE,Tc-/Z8
6aX5W/RRDIfXR(8?[[Y@:4<[A1d/1)^Q^_A3A9b3HV0\LG:@D^f\SSXKO?7T00&f
PWg/7C+G;JP-fQa>L4CR#+_6J5&<cK8^8FG#8/cKS2MQ7/YK-4Z^,EN_+GZ,KNM#
;CQ[3#5F&V5(R2VAD@@XMQ^^T48-fMJ.2:>\ZCSEJYV^)#<SJ]Z:2dZF41DJ:&4=
W+@D[+Td2ab+M[WU)b2]+NE4\4L:G];XFbNOJ:A@f\VI3G+ceTVcX1EJ&/A1-N:1
@_Eg9H;T6FUC73bSN:T<d:2<gGAC_bVb]#)I(JO):O:Bg)W9N(4,UV=03KUS/db5
6Y]#UDPJS58=8Oc7NW-gfIc2DVF4,Q=eIR&eXSSB1A+])9/9_?E+\fa:PX@G0W+d
d6K;D.SLL+<JW0&WT>,0;Y_6Z66JV/>/LUeF8.=0Q[#_(ZFfK7F6AV8KW[.QRHc#
N[f/^XX)07[efPU)FX(?VPU/c>g_-5eQE:LIY_P8Mf8TJ;fV2cHG33PGLd?/?b2=
8AG#RT.:#<D/GMM(^UfUT^1+SLNQ@4A^)b#@)640Z[:,[^ReWVV,,(IS:6>&EF6]
fMb+A@.EQ\N04(T8A^1g\[Z_#eL[ZY7R\O2>;+W3YNWEMRM9OaI@4#?BO1I53WaI
<02C;Q)]5T75LM?<XM8^LY)TCa4J2=1+47\A^I#JCLI77]DD+bP4)gOJ,67)#T6T
AF#9H2[L-ZZ\3<:?B^Ud:240a[R=&\XXGU4B4TF[VSI@O7HC4@//_W#XT)OFSgJ.
D/)8JKD>B)4@F\Z4IcRdYDE\2Bb@G@]=.-<_YAXXI(EQ&@A+B]daI,7X3^4E<.JB
W>>W-YTC3.5()@d6b@PUaATI2Z5BKf;OC9>SXY?c]DQZY?47L8<:HF,=IDgVDD7V
[2X74EVLddT5U6gbUCI<B#E].D3<2)WgY&>a0K@6#E;MU(<=?<c&K<6=N&=]J_LU
AVS?W()Z-.:=51<E?JTG7+K8?^Gff>(Dc9d13+C(VUDC;)4M[[F2e[,A0\UUJ^LR
^MB\U(E3E:62I[gZE<4HPKPL&YPW[OB537S2c3[9TE_@(=V]1QagKfXUQP=BE8=V
Wa;G<P5BZTH,]1.GLR?01&K[#\Z\N^A97-Q51:NIG.4d+Y[V>,Y:Y<G(E;-.E60>
e>05KeX[OP;]e5J_O^01E;(@6LYKbWfd>+>JfYbR9#0T8]FUa(b[PeA<__@b5?]7
P[1YOdIVH1>D;24F::A,9TFUQfU7,PTXBR+I2dK_^0I-0K0#RT\FWU);TO>R;acS
G9?AcY4O5B1D(gA^G3F4Z-#J:Nc).[/e8-CF?6-Y<S?eNbBM[6eI\^>[3)_1[5SR
aG2G(29[TPf<N0+IIMN@,\I[AgAE(c+b_QI5CD;G\7Aa\fTF1WX)@9>I];/MS7R[
ddJXLQaEGfP;-X6BO]Y-7W+S#.[&UEf.[Mg;37&dSY.\g:I#,5B<(QDeMRX-\CME
+bXYB-;GGX/N<_a(,c]+8)@]_A@I:FMg\_;U#gOS&2]5B\^I7#4JY<Y6_4S]^5+@
BYRE(Y]\VgEKPA24PG.KIA5(4=Rc71/X&)6+I60#^YaQQL-3KB-H&bJSGeAe&LPP
eS)T9AO,);D#VW=eLT36),;8fC[dPR3V;^c-2(I0;W;1AYQ>IfYa+HP)/,_X?9(Z
7V@3cR]VJ[/cBR]:1D_c_GdbdT9RYKZ)6OU,Ld\<KC/\9A;QTQMHLP3<Sc-P47H)
I2^CPFI\R]@;\U45NI[BL=J-8/\#;Aa(]@VQ2O8#DfI&&5X=[6U=U<IX>KQ^Hf],
\/7@-VQCHSVaY^aWB^=S#CC(>MUdc[F(4dT@.Z5G=P\XcLa_BA]5:9HKWX0Q&[;I
2F>4O/,>\;&T@=]@94g>&BXWbX<f?&DVRBb)JbXZKRO7gaR^F#aS6eN.KHE,+_<e
ZadYY9IFL-_9K=^9Q@^eTPgPcL[<C6+OKa^[N_HS=J><#,;O?OaHV?R4d\)aO>2P
Og+35g=H:5;.:\XcO60T-b1[LM@HUZUXF3=CWA4L&M<\.:J#-5,F0gZN:KaMONE/
,)Q)K<>WcWccaX^JIcIOA#>R\/KAMIAA\QB7cSP0:PbUf(TXK<D2++(+e\d5)UBX
E1M[Y@ecGOQS:9)11O=F\<K)QRTf[D]Q<^060]Q\N2We4S1\4H]:?]\C0Tf_XaJQ
>V3C9QN65@U8^a<LS-9^DTVf2Y9#HVab]0\=,d663518.O</=\]7@L^RTAGJN_8P
cAR)TH50G_H.3K^gQc,L?3RW1.+N)P/U=.X=WPW^3MD;==#4J+O_R:&)QFDK[3c+
&V06I#RAL,)R8bS[Ng[,-1M_RV=c(<[:f<AN/>VPBgQF@8?eSES^<X+9:1^S4>9D
bZ_4NR5;f+\)KZ(?RS_>5E-Q;2;,(7aCX=7@>((K>CG1UWOS7IM7IR8;bL,X^H1c
2dHU1:SM^(#D)I^[;QJM-ML+[=HSS0]:Maf)fDK.V_a@Rd;RTeYW&L\b__C>3EZ0
;F\Fg>C;6XK[f6G5:dP9[8eP>;=VUb-/8YH1.Ib9=33BP0K^DD7QWH@>.A9?9NTM
S-]=2fCQAY,\dYB;eSFMd(6PC1BE[>89)A>ETS0SS.Fa(XA3N,HW>,0F76FQ.&JD
ZP1:dNKEW3=R\b5<E^E3cdDGP,VbUCI/BL)fA\bM92&>1DO[K/H<QU3ACVN1KY1?
YMabcdI\7B+(N&>a:/c^0C>g9bc_([=?.CVZ926;78eK07<Je#M4TT^PIP:(MW#9
2W]]e8\.KfeJ3W]\SH/I),F[EZDPOX__7S#Z[S-L:[.9.cYZ;e03#==H+L[[B:Pd
W.ZRA(W?W)0X?@E.G+Y\UbS:EA#?KE2K&MW.2&6VW?X^AZ@Q81H_WY\6;JZ\\^<g
ANFEgcdU?X,_^eYb.(PHKQIM7<fV@&(\aRf;VKC@AD8,P139&I[Ze\d:fca=>RQX
d8aA#.QV>3:&OK&QOQ=@#:c:SH6KcSg8<fe:VI/V\fTdA-4[#4<?P@05#3\6R-?2
[gZ1gQ^b+6]3GP_1+ZDeOG?64S0AC56gK[BJIf))]/gPgdKT+0C(.B-68e19VQ)G
8<UY&a8ee=/S+V38<-C#=a?dR11>WO6JHW1MO8?9^NKA=B+C44&D;9.@68]0<#\[
/#LRV>IT@UG=ZeL;Ld.&UbAd[#bJ9)]2RV#YCbEaI5&dI^AMUd[E+c0TG]+IJOV4
#[(01;&Zcb1PBFXS>7e6UAB,TV/:=&X@FLPW<F6]X.>653?<V(50]6@aW]N)>H:=
2Ee[&?,##50F[C#8g?L5DL6B,>VW5_;J_HSI&X.Z)a1U2Ac-FQG;\cQ7\A,<TZ(H
QE?/UON;U:NH2)#L3OW]c>C5[=:P=(KYd5=ERS4BYRb=D(/I0U1P5R+Zb55?P:,P
LE>OJ4]/:<ES2VW-IFbC@b6TK9PM7AS#1K(85bM8W:N1^b,),\=3INMXB0-DUL)(
2)f\aS0VTD5YP##4JRabDQC4e(#R5E(][8OAb0V<LVP8(+bSR+>g^6#-BRL?_@NI
&]5>AA8NU4&-R0R],<.-?1bWb^;SJdB,2SW6MC2K.Sf0JM4C+c27NTOSR.3/4+N,
@F1eMc<H_=1]SQ\LQQMLK[Kb-0>^YF/N?V4:?]V]a4]@Q5[;.;#FRX=P;.-.INHI
-1cJGfD@T@=G?L,9Z7Q5)&bKWZC,6R:8&,GT^PIWg_<2TfN,QdQ;H0WU?6UO:egT
U6:\)HQW6=K5/()[JE3#[UTaG.(:/cQZJF#<7Bg:BeGY>3.&R#NWNNNI6f&XH>39
c7I08MU6T;C.)g4Q[#W]OALJV//R<<]9[3_.:>S9?fAQ(3Z6f@\<SabX-aZ-=_)2
6H(D,TLRA2MV--1A,01]Ng02LHR=Y.:+Y)?B7BKfCV[GJC&A.2cS:-_g31M@6KPZ
]OE<cH-9[PX[.IVa_/FF04]OHaS+^d:b0&@gbJ4>JE6d=F7C+.9<GJab#-4LWSDR
bMeV:F,]<T(f0^S(Y(_RG:P((WC9>^?e(2VC&M?8dD66/]1&8X:UIf]eGe<A9II5
<0[D_3b1-AC3\@<B:ZT--S=/&5]:)]DgE:0K?XO5MTVFbaae.bLGUX5>^a=]:Hec
cd1H)C980c79\E\3),_W/JaZP6@LD3c.;D^1O6V9CC5DAU,ec>?@]FWR(NH3_P/H
FN3)P+<07@+g4f4Z&gFXQe.#QW)YRVb=ERPb>-?ebO@99O^LR<G8Y26F/A<XGege
XSCPY?RKLf_I7(Ibe/9aT_=9TT,5e]B&;-VaNgDMc1F:(YQDdS1/+Z0DZOA:Qe1(
4aaa@B6FE4#Xd73E->1YK3Y3RX^:B/@V1&2[()V?C55RE<;<5MR#+KVS#8N3R60G
VXVZL)#9,ga?dP^P]d_TZ_:@3NE\O_4\c/eVIL8&88;e49cDO/<T?Z7N]>_5SIV@
.<7@:30:4;5:S[T3Ld5\@BXL=WC9aUYR>BOJC?ec9C-V\SY^0J6,a;0MTbO/#QMJ
1HMSGJ5c&^d9^I0^3-3XVaIedL/K0W.?fB>209C;S&X9gf0>1He@IJcK6aUZ&E=C
DJL1W==EM1g)<5K3^+,62#?-;IeI:)N7K?DJF>1d@@)FJX,KgLZ+=SeWI757@AST
ec[WZOb(:O4QV5EaOdV_#N(g]aC:d?WS1(4IUKMG685N;QKG-;R6#0EFGJ[H>?EF
?1@1R3;^3L,/K=AcagB6UNe(@\XWEH5]Zf]BRRO8A??2K;fB=+3=@SY&.T&g^Z;M
&;XMI\C1;C2?W1BMNZgTI0PXSV3K\3gEVdE+#I[eS)YF,KF6c51[Y@XRbEJB0a7c
GaJG>C@:SV3]]8e;,#HX_IET]1@4ZaFP6+PT>0R/gC^E&5NWDaBE2[O_W1cG?R9J
=64CAEJ:([-LAR?22T@6AY<?I7R#TP_eT1,?^N&BL3Z?D(XWFG-c]-\HGE(O&()+
@L/Kbg:<E&DSULJcPf8ING\FgTc09/dXAd;ZEO>VBW:>8J-+1)c@F<K0XL?N#Y30
CDN&CTVHS<JZH-^=7,U:D:EB_?8UR]Z/&U0^g6ZZe599OUWGJ4A:/fLePF;6PWXW
-6LEGg9T]U,C<^@__cdgV;41Tb7ecD-P1FVeH_G?YQ8<_;NUM/[b1J28[;,;,BY:
bZ]-a;_+Yf1A\R9X(___MQ=fM8I>TE3:63VT7_73ceg0c.b7f(<2-?1[6Od1F5X,
d2g83f[Lg?/G3_CB?M>93:_VFF2VY0SF?1OW22+cUC;[5ND-S\We&cWfKM.-]+V8
a1&4&DLI&T+/;\::gEH/cf:1R9)L1XUJ6,UEAO)7,;)>2ARV>G?+]@7?^M0HWT+T
GTBK9G+U4_BfP:Q,&9^KdWDT-@9-=_6b:&OM@#A09_gdcL\EcH5AVdd/MJ(KE#5K
>PGM>e(b(-_&-b/BCO(+LW+Ha^G/Q@<&(DMHT;c7^>I61[=ALHWeG?Ue8WB@ZNLd
@GON8,bV72dX13bI6BgF/>^_<g]f-&?T2@MLECJKY2d^\NN\,UF#g_WHX\#(7&A.
^Fd./Q]a/2RXdW7/fU?RP]W/cTT@IHIO;+,S0;X9.^I2@1\W-(I+X?Y=STRb=CA@
gN,)H035E)1#<eY00+H^M>3Y]L2YG7O@J6Ke7[]UW#7#PMD@8@YE+0&]GUNf)ag&
&9B3TW6/ILbAOdU^LX:S:R@#dJ3_5WdOT\P_PN<#7QVR,\(G,;-(9Q1SeU.g3aGQ
YS_5Fg-W#N#d6XdD5>.=;3<7PEg:&W59X2OgEIb89cF25:2NX/I:^^3L<UBF(AQJ
DM(6_??9a/670DDXI2:S,UNWdBR:#Q0X@M=WP(QDM:a//dD9DYJ=IHDgU/21##-9
)<DDF4O0([[U6F:aVHVR=U^_]De4SSN4\CT62)K\7=I8AHU69M>4THgdY+)SUJd>
<5EVUY(d@<0,We>>D,>.g(TX#1d,?P@F#[eGP8/MN2KRJ].;CH9BI0\>1>dOBOIE
bd;1U)JQS^/6PFANZBE)SD.QM4:Z#VVgO&_D;2&PK#b\f&V_OCX3Z5Q[/O3/dIV&
R>cgURDWOU78c:c4CG4I0=(<#53;B@4U[L]@Y\LAV<XQ8(]CgT[8=5HQd-UO0ZI<
CS/X+D@9S#WeLP5c?^+]QeU+&Ef5)Y<]9NDP35I.Uf]E)#g)EL,1W=WGVG>/170;
_W--HUL;I)^c036)1M6PZdTP7VH4g6U=_eVTR<Nf@8>196VVZ-E-,AC\QTG.]KZd
]@5,OA2:VD<@0<XM96(,]I]G>MKb2JQC#ZeJ>>DN=b+#EU?YT;Gg,gUe0,N4=IFT
@#^4SgIf=a3^GFAI//EB;4PXZ0>a8I)H=\TaNRC)[W#YYg&7D.6+b&K</^9)1-c4
9-6@<6A&Wfcd/T]C0F_Yf9,5>2I,7]N5(1Sa^;GE^1ePKN<U(<HfH98/_OGIA?0b
P=c5/@LG.Z0^:aE2?,=04.:aBE/4db4[E)Q_FU?]G]8Wg\X8cA?6(_a=F<:,V\<U
TVQ5+JD2.f2:2E36Se^#R)#/X45L&Z/6FOSE;HcFJ__gY.#P0KRf_fC\(XM92[07
cAa(J9E/YT);JcS8&C2f00/64fa.>#SKH3__=@OYRQYeJZ?71<P^cAG1[7D]0B6:
>KYS/-+7/)(TE?V:BL9JEL](J8KRV4:>[I\W8FU)1TTHPTZTI](Z^YS0LA50G].\
Dc4>Hb)/);+:V/gS;^8XD=ca:Z(J//YIG-\9;7=HHG<Ed1:L_Ngg7_[.6a#4Y61@
T32G;DU^^0eWbT-e2]PSHYI]=2+[GVJ>[@Fc/LaFZ5>Q30.#7I+:KN=XadUg;_0Y
c??O6+eTM=Y@J+97](X>1>ZMH#BM)RKa?XCWb-(O3>S7+:P;\F<:C66L>ROZI_;2
Qf:V;1&(SZ89(IC68?Af&Q0SUC2-Q?M#51VV0&OPe+?U)4_EXA>S,WS;)MJVXO6Z
D]V/Aa&/75Z@/:AgcYCJ0YCYQI<SM0VN9YgHR:^eS1a:C2>V#7Q+4b92YH:+#/:X
W>g)I+e/0I4]4C^2>6/5GeCD:)V.SGN:HRTeK)0?K/LdU=JY,Z.,IZSR+e.HI_N:
SDV8ZNVM1=FHH#V1B0O;F;GS@bXWC9]&UZ7;5TV_Bf?LZOA3:\/6BZ.OV(GCNH1F
N/DHg(e?C:c-=b41gWYRWUabCKSU0ZT&QM]1UcD(;DZX<(L\9Q_7IB@QO6EA@0JP
F8P6LV;<V;XIAgb5aTWY</UBN&X9b][c0?WVXG@OT3a/&:BO366J#BPeNcBDd?^M
]JC+.4.M/FUe&/ME+bT#_\:7-6\H>0ARW)T9?Y[,aVZ(>Sf_]b17Y9[5A8OZWegd
)0ae-SVHP[72KeBD,e7BG7TOX@3AK;Yd(c?,BaI-Ef,B7DJGa)G(5H2PN(&:ENBd
MU<EC22g(><J1&K^E.4YIG,3F:<2MKb#[;Qa@>Be;&7a?TL>+B<CP=V6O=^O.FZH
D_M[CcV+1<PO=#N>:3_+&@-J<2PP2d)H2J>EX#ge<+?8@]YLM.=-2?_bCCI9RRJI
:dI8)>]QLQ\<,K=RH5W,]#\VS0&AVO;5?HQF)cLbBbW1:JG,PQ;(_>3_^bL9SM^]
@J:8CL,:E>0d)f(7V&BP9./Ld?#B1e=be&\92^f8SE_f#OL>L8=@=0.IQbb&GI#S
3bZRS>3A[M/7VV4IfId)gHe[U0eaKTP;^3Sb5^KRP2H)#VFD&XQ^GKJERQ4.EI)0
OJ=UeF=C##.5N:5ES72&a[&bgcU>U(Z1X)85e&YV;b5LG1-ZQHbfPB_e3V-3HVPI
=fV(3V+\b0<-7Ha=&0&V_Ne51cc6:4&JB_[;)P/Wa#7dXHW6USF=N5E2>7@Q,0=,
HK/Z,3VFbG<D,<FKALB^;#C8-KWAEQ,8&.S>QaIO-S[QN4B3KH(HS()ABLZHTL-(
P&IE\=(#DWMg)CfL&K6XK9Kb:W,1M6d5)+P^1BVdS[I]QM]^3DU<NOW->_Y/e1FP
X+>CMZ_U5Na&E/e6V@;I+RLeM,O++[P6SS6>T3@D/NBbaZMM)c>a8f/C0&A09T8@
cNGP7HH)8-D9G0(e/)#2dKXRF>F7+J?<T;;6R3K^:,IJY+#DfMdS=1W-5gE(EH\-
-?f]#7O]6PHSE<947EY.A;B],SdC.1U1]AH/_dJ8RS-JD$
`endprotected

`protected
80K-QdGKO(.MEG1YGB<D,E>@9>4XA@G5+)LX]52b@3]RZ_b00b/D4)@Y&.Z-EJ5C
?=./)F[.)TbRB<NDRLB&NK4+K0c7_SdF)Gg@WRCbP.4-@R]=e7aY4+@YM$
`endprotected

//vcs_lic_vip_protect
  `protected
c[O-UIYQPN7QOO0Y1J;(6P:FB?)@If>X@WCJE\dWY6R4bO0AAIS(+(f5g:FGJ9/Y
?)>:)IJ^RI6Gd8NdWT-Z.(K)G7QWTKd=dec]QN7Xe]Lb.(XU;@fH-MAdaG/L--&(
aZTL,?_I]1,ZJA92FS#8/]G1L5CcC9^<Z8NFgdXR3SQDZGSU3.[7:GJ>ZRD__-gX
/,G1UT9XY^bU&<ULGe2(]D-F[CZ^<bS)e,>6WPD0;((FUaOaSR_-VZV<df+4&e2I
J112Ec_#97fJ)<N]M9bO4@Y-g4;632_3&b6FO#R37ZDUb\e@<ad+-N7cF+:@Z:G.
3OT6T)I2R-VTDc\E9MEA/:\2SEdG)G5CXZRRC(&e;5.UG$
`endprotected

`protected
X.,].X#IO@[Je@eFE/4<Z?)\YJa38PA1O\ROO<cUG.W)11Ig^^12-)gUFg-#@;E#
>9_>e)Z,S27I9LUJTFAc6#b0XNdOC8c0e22MC=eF0C9W4Pd7@-D]M&gUL$
`endprotected

//vcs_lic_vip_protect
  `protected
bPYH-DOcK=UZ;(VULU[@D#R18FRXf41W7b/\XYC9+RDJFfUV+W<@&(3b2&_U2AW@
):T>2^fUYd.[5Z4T+ZLC9d8U?9CVaNe-4eP;LP,Jd6QBW0@;O4.fFa,df>>BcWWZ
>9J?gg^?I/@gE/-)DHI69+8U8$
`endprotected


// =============================================================================

`endif // GUARD_SVT_AHB_SLAVE_ACTIVE_COMMON_SV


