
`ifndef GUARD_SVT_AHB_MASTER_ACTIVE_COMMON_SV
`define GUARD_SVT_AHB_MASTER_ACTIVE_COMMON_SV


typedef class svt_ahb_master;

/** @cond PRIVATE */
// Note:
// This macro makes sure that hwdata is not driven beyond cfg.data_width.
`define SVT_AHB_MASTER_ACTIVE_COMMON_WIDTH_BASED_HWDATA_ASSIGN(width) \
  width: begin \
    driver_mp.ahb_master_cb.hwdata[`SVT_AHB_COMMON_SHRINK_WIDTH_FOR_MAX(width)-1:0] <= beat_data[`SVT_AHB_COMMON_SHRINK_WIDTH_FOR_MAX(width)-1:0]; \
  end  

/**
 * Defines the AHB master active common code
 */
class svt_ahb_master_active_common#(type DRIVER_MP = virtual svt_ahb_master_if.svt_ahb_master_modport,
                                    type MONITOR_MP = virtual svt_ahb_master_if.svt_ahb_monitor_modport,
                                    type DEBUG_MP = virtual svt_ahb_master_if.svt_ahb_debug_modport)
  extends svt_ahb_master_common#(MONITOR_MP, DEBUG_MP);

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Virtual interface to use */
  typedef virtual svt_ahb_master_if.svt_ahb_master_async_modport AHB_MASTER_IF_ASYNC_MP;
  protected AHB_MASTER_IF_ASYNC_MP ahb_master_async_mp;

  /** Driver VIP modport */
  protected DRIVER_MP driver_mp;

  /** Flag used for handshaking between phases */
  protected bit drive_data_phase_active = 0;
  
`ifdef SVT_UVM_TECHNOLOGY
 /** Handle to the UVM Master driver */
`else
 /** Handle to the VMM Master transactor */
`endif
  protected svt_ahb_master driver;

  /**
   * Flag indicating status of tracking transaction.
   */
  protected bit has_active_data_phase_xact = 0;

  /**
   * Flag indicating if we have a preempted transaction in process.
   */
  protected bit has_preempted_xact = 0;

  /**
   * Flag indicating if IDLE_XACT is becoming preempted_xact due to
   * SPLIT/RETRY received for previous transaction.
   */
  protected bit is_idle_xact_preempted_xact = 0;

  /**
   * Handle to preempted transaction in address phase.
   * This is required as the preempted_xact is local to drive_address_phase
   * method.
   * This is needed to especially invoke start_transaction() for preempted 
   * transaction when the address phase of current single beat transaction starts.
   */
  protected svt_ahb_master_transaction global_preempted_xact;

  /**
   * Handle to preempted transaction in wait_for_bus_ownership() method.
   * This is required as the preempted_xact is local to drive_address_phase
   * method.
   * This is needed to hold the transaction of second INCR which starts at
   * WRAP boundary if the last beat of first INCR receives a Non-OKAY
   * response.
   */
  protected svt_ahb_master_transaction wait_for_grant_preempted_xact;  

  /**
   * Flag indicating if a rebuild is waiting for address phase.
   */
  protected bit has_rebuild = 0;
  
  /**
   * Stores the wrap boundary in case a rebuild is required on a WRAP type
   * transaction.
   */
  protected bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] wrap_boundary = 0;
  
  /**
   * Event signaling when the address phasde of a rebuild transaction completes.
   */
  protected event rebuild_addr_done;
  
  /**
   * Event signaling completion of transaction.
   */
  protected event data_transmission_complete;

  /** Event that indicates that its time to fetch next transaction during locked transfer. */
  event           fetch_next_xact;

  /** Event that unblocks nulling of global_preempted_xact after sampling is done in case 
   * rebuild happens with SINGLE burst type. */
  event           sampled_global_preempted_xact;  

  /** Semaphore to control access to driving hbusreq */
  protected semaphore hbusreq_update_sema;

  /** Assertion time of hbusreq */
  protected realtime hbusreq_assertion_time;

  /** Track if this is first drive to hbusreq */
  protected bit      is_first_drive_to_hbusreq_complete;

  /** Track if first assertion of hbusreq is done */
  protected bit      is_first_assertion_of_hbusreq_complete;

  /** Handle to next_req set from driver. */
  svt_ahb_master_transaction next_xact;

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param xactor transactor instance
   */
   extern function new (svt_ahb_master_configuration cfg, svt_ahb_master xactor);
`else
  /**
   * CONSTRUCTOR: Create a new common class instance
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   *
   * @param reporter UVM report object used for messaging
   */
   extern function new (svt_ahb_master_configuration cfg, `SVT_XVM(report_object) reporter, svt_ahb_master driver);
`endif


  // ****************************************************************************
  // Configuration Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ---------------------------------------------------------------------------
  /** Initializes signals to default values */
  extern virtual task async_init_signals();
  
  // ---------------------------------------------------------------------------
  /** Initializes signals to default values */
  extern virtual task initialize_signals();

  //---------------------------------------------------------------------------
  /** Drives hwdata during busy based on the configuration parameter
   * data_busy_value */
  extern virtual task drive_hwdata_during_busy();

  // ---------------------------------------------------------------------------
  /** Update flags and drive initial signal values when reset is detected */
  extern virtual task update_on_reset();

  // ---------------------------------------------------------------------------
  /** Accepts an incoming transaction for processing. */
  extern virtual task drive_xact(svt_ahb_master_transaction xact, bit invoke_start_transaction = `SVT_AHB_MASTER_INVOKE_START_TRANSACTION);

  // ---------------------------------------------------------------------------
  /** Internal method that accepts an incoming transaction for processing. */
  extern virtual task drive_xact_internal(svt_ahb_master_transaction xact, bit rebuild, bit invoke_start_transaction = `SVT_AHB_MASTER_INVOKE_START_TRANSACTION);

  /**
   * The methods asserts bus request and lock if enabled. 
   */
  extern virtual task start_transaction(svt_ahb_master_transaction xact);

  /**
   * The methods blocks until the arbiter grants this master the bus
   * This method is not called in AHB-Lite configuration
   */
  extern virtual task wait_for_bus_ownership(svt_ahb_master_transaction xact);

  //----------------------------------------------------------------------------
  /** 
   * This method is used to check whether transaction will cross the slave address boundary or not.
   * If it crosses the slave address boundary then transaction should be dropped before driving it to on the interface.
   * So this method is called before drive_address_phase method
   */
  extern virtual function void is_slave_boundary_crossed(svt_ahb_master_transaction xact, output bit drop_xact, output bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] min_byte_addr, output bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] max_byte_addr);

  // ---------------------------------------------------------------------------
  /**
   * Drives the address phase for the transaction.  This method will block until
   * the address phase is driven.
   */
  extern virtual task drive_address_phase(svt_ahb_master_transaction xact, bit rebuild, output bit is_aborted);

  // ---------------------------------------------------------------------------
  /**
   * Drives the data phase for the transaction.  This method is executed in a
   * thread and will release the drive_address_phase() method during the penultimate
   * cycle of the data phase.
   */
  extern virtual task drive_data_phase(svt_ahb_master_transaction xact);

`ifndef SVT_VMM_TECHNOLOGY
  /**
   * Transmit response to transaction.
   */
  extern virtual task send_response(svt_ahb_master_transaction xact);
`endif

  /**
   * Executes the steps necessary to complete the transaction:
   *   Completes the driver's seq_item_port handshake
   * 
   * @param xact Transaction which is ended
   * @param xact_rebuild_in_progress 
   */
  extern virtual task complete_transaction(svt_ahb_master_transaction xact, bit xact_rebuild_in_progress = 0);

  /** Drive the default values of the control signals */
  extern task drive_default_control_values();

  /** Drive the default values of the control signals */
  extern task drive_default_data_values();

  /** Drive a beat of data on the hwdata signal */
  extern task drive_write_beat_data(logic [1023:0] beat_data);

  /** Drive the address phase signals */
  extern task drive_address_phase_signals(svt_ahb_master_transaction xact, bit is_drive_along_with_busreq_assertion = 0);

  /** Ensure that the tranaction is valid and that the handle is not already being used */
  extern function void check_transaction_validity(svt_ahb_master_transaction xact);

  /** Drive hbusreq signal */
  extern task drive_hbusreq(logic hbusreq_val, svt_ahb_master_transaction xact = null);

endclass: svt_ahb_master_active_common
/** @endcond */

`protected
0U2U2[0FBd4?>\X\/^P42FU-#:-&P^YHBG77EQ9b#?-Z50)0K>&K&)VTFLJ;QX()
^(F<[Ke_IV<?F5aFM>?6.<76(Z#O2d)2Wc;OPD&4?E#<(LFKP398O^b=<K+MJEU;
c:\e>+A2&<dg4?)X?,8D-LLc^T6^T=>Q(76Y@3;][Eg4^A#D?Z^de8XQ3G6dK<f>
;IcR5+@-C@R):PX4GHQONDI>KeB+;WZ[[KFILa/5+\__SW6[;2eW+&SZPbdR6Z\g
#-PKU#[3X/(-RPDWW2g-V#;G2@K/BTL=FbKR1T1_[KJ20._)#;0[5&MS&C;GA4bM
K#)@+Yfc2Z#1)@GNOK74ebD>;c;a7DW\,gF]#O\#O)T-.^1JWU^IQNbL;fGe]AP6
(X0<]4PYH_&R#KR4E7_)dP,^6N#OeJgSYM&dWF1>5YMJ+<F5bP=;@E9&MeObWLM[
XPYU&_[E+U@1DCRX,34+O^[Qfb7/eBW&aMY2K)I-2B\C;VaI6_Ic\87M83ARg71)
7dd^0Q6[O[Fc1D>N@IP@4O&LbMfJcD^FQG:LaRD4;LG6L)5HbVK/&87<(KM#&N&9
8?03c04KQ77@=0XAQ>FHG^]+SHe7K,bR+S[:CEO__F&Agg-T<I#2Z=7<P$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
]/0_T#O#(=<,GM7<ZGOX3G[WD?4QO:e=NeI#899#79@HGS\Z-8\Y1(#.IH?T:9]G
/a;O(;NDgU;3-A/&P8[C.+GabW,DPET7APG:+#a&4d(9L^?XTTeBW#5&T_F;#.@d
JfTPe]A5N8YKX<eT_\1><9f\M1PeZH95OI3IK-XS<G-,NSJ=c#Nf/QUP?8aE_&4=
O,\6SLG#c?-Xb]KGTP8VSY.-\QGMegM\0eW&:dC8R=Eee.Cf2UQSU&?#VJaQ0>KY
7;J/^&R2(J=(W[.4,EAVdMeX.;_cQD:/EbcR.K66I^H+NQYfWA^5.GYa>&NJe@6g
7:691Y])ZB12_1E.5G=O^-A_H:YB,=,\cgSZ8\])B-;B_]);POGW^(.-VZ)ZIgNM
/eC&F/ILO;B8J>0_]A:_D0V4[KU_9^Pe>SRLFBce93)EM5,A26&M&F?(EV&_&3;T
/;IRKc&1(+)Ra=^Q23@RHBSbT4acUMFQSdgQLWAB1]?)N30KB\H_b(@Y:,EIIcXN
:6?1b+03;R\-X5U_,CT]<#J[)ZY^d0E19&],J5I^QY&PTG+5<OY_Z-,0>B94(A]/
?ZQ4USGdK,fQ-c(/2@1@b;_E<Z]59g/4RDa0f7XgU:.8O&]^WgPEHG@#(EMf&:e5
B99.]+Y:=L8C.V?;a2V45[/?+fP,.-O9b_1MYa8Ea4:.9Vf:BW?G@J22fO^7fBK4
_d0])6)1Od5LSP,__2BVR.P#^HJ+g.Hg4&/]7K?&X&cBVT/N>UCC\e931&,b]&7I
GJQ=cSRZ?38A/3QS)105a]_(?>N=^/,Z@bX/:OK7Ceg&+@CeH(eHCa[M(YNPX+,g
@Aa^WDeO26\\JEKdcc_)9?OD7fL#B-Y#[F#dd9X:S3^QJ5HLZ/dAB7ZD3#FC^:RN
FL;B>.^93g9)AT[G7SE29&LbHL<NS.CC>eY(3<,T&06>(HY#)6g6KLJgC&3cGe7K
Pd,#6SXf5W4/N:f)2@g/8X;>3-18b\MP].c?Of:E?PL7#cQNaS,V>W;P@ZTE3P?[
6@N=-5/:P#GSD/QD0X[gV@@^5T0\5@_GF;+C63#G5(/AB]-9]/Bc,baJbV=ALGe+
4#.CN7V0EMR48:79D3HKWR^7a45=5Yb9)O4]Z@4H+.8eHDI[RCae)L#?R<J6FSK@
c\Gfd\aM)LDWXF)ONPAN[C/fg(VG)#5O=E\0;0(L\)dPT=CN>IEKH[4C.S8.UcF(
.[LVDS&>?&CKQG>X)RD(11_CU^O.UF6I#aDVdW^;Db&J/QDQ9_X]0LE\f#0DRf1M
[#>]^8IQRJHY<@:SeRAVgF;W1D:Q0N?gY+2,UD5+CTZ]>g_b9\fc0E++9d&J#\<Y
SeZ>.Q+,C_=cY.N?BN.G/G<=<F=;\[?C]A(OG:c1]K.81LE&F/d]E;]63M/Q?B7e
(2<4(N3+b+Z0@@(P+[6fbW_4&[@].9gfK.FR^R@I]FM9=+ea)K>XNG7]cG=[-)(@
^-];DDA,1>@=b+B_77SXeH@1VH_+9=61\^.]@+F(DPNg;gXg^&9]#:>H[0OJF^&Q
(;D7L,IX\71,;O48E+@3FK[TXKE#NPHH4ZH4>]5)87:)eQfOZc1I8U@50>=bI5\3
:I.U+M=FP+(6S9>YB0>8=DQ>bc2@BJX18:RP;^U<K@YNbH33XG0UYa3eSE:8O1B\
K6HGJS(#e8?Z@(CNO34.SO)gOX^gR-(cU9AAfX(@Pd[#GDDKN-b=fRW@KDFV@=8.
-e(I[[2]MW-G.HaGT4Kc^HA6EN+;Cg)R)Z/)K029#8IY##/Y[Fc7Y177e6+74@>K
+T7BE=_G-1B@Gc/9]I2SL\OC][IJ9CEM,EaGA<8#N^A]8;OBDgN9PB6[D(-aH&.;
]H:cE)EQQee(2S^8BePEC5HRGFA63<.#0CRK:F&R;XEJ?&W],+cY^_R9RV+8-I)+
L^KCTVga,,WfO?UNC/TDO&XTb>PNH8D0>NJAb<8aHWOb=JI3Y^d<H^==^\aGBA/&
\e^SVcC?M,L(cF6?Q.aOPK]]2,UUWUIX(dXTL5eRVa9WYd1,4CM-&^&K7];a(&2A
c\</SfA.==LJ2Z,;e+EU0),.B;]5[Ld\]DR^S,We)Ae^B,U,YA9=UOd9cT(=E-GV
H,2:&EWbe:;E)L4TS;T547IG<>URZZ#d_GJ-^[V@\-D+4<>)?>OL8I^K2R.J?5e&
XG@,;c,1N8fc4XZV:KI/RJcGCF_?c55OgbL@faM7@@O8.]1VH_HgR&3WTXZ1D\(/
]QaVZ730f2)\#<9FYZVbOSY2I[6[/+@Oc-(,A;@3X>OS7[8JJ3XaFI,GGS2#CZ(N
I,9B1/]GE_));+dAK3bDJ=78L]LUDG^&W+(#YEZ(MAI311Qf:AdO_8EWEQ=OI7OD
MLFbP4b?=(HTH[24C_;S;E0f^=Y6=Q85R^^@1S&MW<P.VFF,E(?Eab;<GTD0#R\O
Y;?<9PRZ5aD+c+:bgZdaDYM[cTY_L,a.UF9E7Q^K\X]]7LZ[_5]Dd7SBDgESXUH4
D53:KFcf.RX0dB2;TdP(QaW9AKGVF,Q^5^(B2YV+P4M0Fe);1)WdLA&(1QfJbTQU
3QAK<7@=89T)T>>d7f36>;,AN73]F;=P#,9:VX5\=?@aTU0bTb0VQC(B?V?B#\VR
JVYK.&1aDG@X[P9b75AD2IQX[Tf^H[+.Fc[2FLHAKGRIfN;N-d#eP\>)F,Ed=C]_
W&KgB/f))VSF?M=d0Q.g(G9g80.)D49/Ee&4;C+K.<EV/a6A&+RWQfK<H&4DTS>d
egU6VIQf]U,;_)3619^a&S5@3C/;>3-F/Q6PJD?;D&-W3ST.eSO2(4;U:a:&5a-Q
TfKAEP8aM-7Pc<9W5-?I&VAFO+bgV-8(b)/K9(GFb^UEN4^-T6G_:;F+EaJcJ3b0
58NI(0<LNGK09(DLY,2gH2f#U8a2N;E@/a?I,T/TR0ZK\3dNNQW2^TH_G/_LIaZT
GISA?;=Y+V+aZ9aA6&VHN(W(QZf4X6E4Z+c.ecD(B/8RWK-KX,Z@>MS:P3a2>ZV5
8bQ=D/NQ/N\b>A@ZGfdYO++6c+<M.._E4?\5&D>,fV@KZbdc&JA\OfD^g>L(I#54
I],]fR,EMZ^V3eg<-K?L<[#aFCF:D&(?6BA\BD(5S=UM5bI-Cga33/bAI;^&=5d)
W(O:OSM3<e.J8Yf=cY26&NXM-W&>V;J.71YYNe\_4WHQ02MgAF27-^Q#_OO-DJ.:
05PR6@2VYV6YV81=,d8GXE>QUORNPA<@b\LPZgI-@)^C88OcLZJ,,dHAU&BXQC7b
7@BU][3E9\.;GW3.CQBQ0+7(>d2MdPJbE]b:MZ-]XBBUX++<]WT@W+9@>??9,Ec<
-<L6+.U(6-7E&c=U81Sd8I..Y\2U-Fe\\c\1d6+JcEdM+@R,^bD:(6RFV,GLRFWK
\UG7,1OZY6S(ATLD4P86HWPT=,-c&39d]8fcNKLf4O<<R.?N:GDUYW7,[edVD9OS
S)a/S5M)V8DZOP5&;6_N?(S(=^,D)^@-(d3L)XR/YH+CSC\?>bBID+#\gR+9\(5N
HL\]Q^DW9cC5;@a<<cYJFAO\J6)VTTCJZ3@BW0gQb[8IaH;)fLI:=JWT_I@).+,.
Pg7De=cT<C<.Q40ONQcd<;=1JH6\M&9,^D#)Y&\.SR<QNZ)R<__cG4#W+=/RLe5(
0Ng9T]7Bg?6B8Z8TG=JSVffXD6.6MQH,>N##P\:bIAEPYO0cO/1O0+YMbb+F3S9Y
S;UQB,0(1g+&S0VO0D/?WH1dE2.I4D0?>)F0e&6^,6b/5D<8<_Yf/EG[S]2:L#&K
3:.@Cg_45[OFPF5\HW>+/g2<bP0BL-a&PZ8O=+=B;bX#;/8M7WVU^H/BB\e):-J5
/L]?J6?88O]eCMH(K<5E,DE@b@7)ddc&+.KRGXb7B6JN0?<9g49\^\C=>=V<0@IE
O+WfLcg0)OKAMdAPFe9XBc,;462<:g9Xg#;4AQOMVNBY,^J0WEHg@GB3MT=G<^-]
:=La,A0:QR[;,##MVA,bZ#@MFcf>ILE9aV](F8[=b&6UYYIY?6L;/2ESO(La6M+\
CO5@=YcE(;R7A203O:GEf#F-ZWagH25I>A-Q(SCRAL]1c-bQ-SYX/B5:@@8;BeHE
2dD=WcDg&_>TQ^,:>90-E7eCPK>ME/V[\),Z0((8+B(6Ubf.JKR>0LX;Q/<1;=Zf
U8c7?b+gY:gU/0^3@[D+U;>(ea4g97/)<gEg(,A(LH76N>;MW(XVX]XHYAE1),=T
<-aE1@GGR4N6Fd=Na.I?gU0/0?1[7</DRf#dPTFeV,OHTBERW6Eg9_0?]f/]EIBJ
_g#^O;,D@9IHL:-[g>dUZ:a<:+7K:HPH^10=8We5BLLA:VGeL@V56D125M58eK8>
K]QNb>+/B/A/+E&M;RC-96fDdKeg>NC=O6aTL\W>]c2@TTg+C,(<,258B^QOCR,[
-P,DKb[9IA6EHYNC:SFAW.?aETAeIZ97_Q-Q8TeMK<C?G+)^;)__0Y6X\c.2WV@C
7=C3CHJW9E/fd]VcY[GM@NO<GIR0g:VW#aa3adPI(2YWKd[?D1[+G9OLDDaIQ+^f
B>54WGYDU/#\Ae<N#:fF21=;)@LWE66;3G5M^Y;caMVTXP1DW10\_4MeCeD;F5T;
/YW[BY\25Q@W0,g:55:O2WET\dJ1MCaAPAJX3d&b#+L&H=Q37W[4<?@A1.L4<SAU
b41W7f,JN)_Za+3;7?O_Zf.DOTB30[9XGf@P]&RVRBFcS_0;1c>?<_#TFJ<MdVd/
P[K2[Z2J[0PFf=:Q?DRS?/<A8F_N.-Q^^YU^P6QFH960aY?dX[WC-PCCT[;dFDd[
gLM?3-U7Rg>fQg]#JV_ND@e&>O=OF-+9cVHI#3HRLT0D5gVOU,UeR[96K7@H:8]T
GJP?P/Cf;]#@:X,T6.MJc>fQgD2e_gU@(Z^=\CC]:BBKUJINOSTJf+_3OR#=X;()
52aL:?5D3RH>T,<UP^afT^M24:(>F&K1dbVc+A8b<-eF)a[SS2:-5Yc(c8BZ3#&D
df.37O2O6OG7T3Of8<&UQWHJbVE;5Yc#/#GWZ#g.;0_+#9SO>#=+:#VQ#DVAB:R8
^N4\:b9)7LQ(JU&<@?A,Sd94L-OW0aFdg/6UQdc.\H5Y50U/1-O=UN?<1/<IV=9V
U=]Le,AL>3g(ELeBeH[/#;;PY4FY&eT6_d\MVDU&X=g>e4<JFOGceg#PGdQM+?MN
JN=5Z>0eZ=Y1Mc5G?Z[,3dd7JP;SF(E+-=c4M4TD23]_L\<G(QA[L67Pe7a]fI<K
^R@3P+<9Jd_;WfW@b),acY@===d-B9#WAB4L=I^TFCA3QB\;YV3<>dCY12Sd^NTd
8B+e;Rd+OPL7#X;UQH6;8R]:Yc5UN0M[2]7=SfTCVDRWaaFJ&M8F6,K],4^U_6<R
H;<L2HG[X24;OYFTM5?MF-a46+OeQ6d&S<3HPbB4fK0.fQVPMV&W[>GC-[1_?#SK
6H,+/_NOBGI-2I@2d/S0<IC>B6/JE,/M,R2GLc5aJ+U@-G)PA8.&DO(gTBQ/CN6^
F(+F_TcD9L8aB/)W^T>/NYeGg^9SO.PJa9@Q^#&@R3f#H>RQVVg#ZQNGa(DA7KWZ
2OVY?c7Q)C0E4X2Bc<<#WI<,]=F?.=P-^#g-MLC.^eaSTMgCTAN,8>3ISX=L>+F9
67Fd_.\H6X31I[(,WAG/-5gDBR9EV4:/&99#VNOHc>,dWW0HOcC(_2Z(/<Me<aMZ
dA1814&I;CX0G/E\KTaKJ4-L?1J_DS#5#g][@?(<3FfKX,\SF7aP^T,^e\)gAaV[
#IXacF(SB+6F31EKQ_K][)Y6-Q_D9[Q=bb6gDOJOOH;g[Ud<0:XP5I2)&4<+?229
)9S_e_2VY86SeX73@RR9[_A(0C>]J6E7:(?eSHG(/G,^P=7a5M^8b.;A^RYG;4f3
ZAO@TZ/9g4ZOJed<+4g]/DKZUU\UdH7:3ZABMIDR,6=a?>6bFdN(?B_-53ZD^<UI
4,S\7Ob@d6XC[2CFZ[=/JPaB7a[J1egdfIM53UaR,GQ(Sgf)&_bFE?3b=Ig0McTG
&F5W&FbH&-LR8>_1gQ&g,KTLP&F>aUT[,;[:R/(aI?I5LFIP+V.1BS<0dg7\_&?d
1>I@>+/5@cP[W:7c-XPO\20[;W91>XQ,JM@JK:O,cOTIOEOTX(_Y0e5L]58Q2-(L
)Q+6&e)XUV29H..?^S4RdFS)DY?Q8/a=3ZcJ(LEM+3NYYVZ3:O.D]W52#.)DI;LZ
I#NE:_)5Cf8fAJAH0/e3L8c99&(]W=R55eR9=3&@+><bD0^SUFZOb@-];gRF,IBe
[_7[4)0B8_9;K3?dUNW98@HBeL^eCC8S5.+\d2@-aGM&fdSb=TK894_6]6-dG0R8
C,0U-A7Bc\6FK?aWBa?+Q6G7e[ZWV@A[NfM>_FSH,L;9RX,.<](_b1f9fX9H8W;+
F@<-/,((SUUL-T>4Va-\,O[NcW-\Ie8_<EM:H0_HgfP5RRHO?:F57.YaLG<N\b:&
Q8GUZ:R+\36#IF-D#+9-^ZWBQZB:HD#BeDgIZ600]81N,37\]2B+YbcX>g:VK3Y6
@JbT]KLIHW0B=?5NP-O22UE7ZB,a)AUN#VAUBMOMQ7],aREb)&XK5BDM_)LbZe[e
ULc:/SE,8YdJd-7d.UUDIZ=/EQ&<LLEU2D1YXEUa8cgE\_#@5-daSRI@&E,+RU_.
4D:6..(7GEgUH(?WQ&[\PP,83&+eR-16Sc[Pe-32LP+VZLE>S6fT(H,eZZ(X:O8O
N+,2)+^-KDCIR5VOC#C>L/G7+gNJ7f5^d=V)B+]4Y8]0=aMe_Z#eLff+PgAM>IXQ
ST^;U.MdIDC\?bfT0BW=dXK:81RD8ZBE-V[VLd:Me;YCHOQ^9G(cLc<,JFbVcX.f
<=]_N>d.?CF+QF^_f)MYa=SXb76;[R8#(\KQY2H=XU:N[XSH;BbZ^>5&\a,a10Pe
VQ6PeAc\T5H4VNcT-KO#0eDLICRea/CL1P?7WGO.JCB7F)DD/CfR^L[GH?aN7?Ue
0Q;JCd7XT,gdeD;ET@__?KBe@Qg8E]F_AW;4^93=&[RZe&EX,P34P(Z:@GI8TdeL
(L9+9fNI/?1CXaQg;)1?,T9I5F_^&dG.U)T^XE6#NNX3H/fJ&FE\0I+P8#88ZGXZ
SgVBOU7e6/UWG[/99A3>.Db<:C>8FA&f/?]cAXZFMB&2TZ54cJ-P+c3g1RR5=Z7X
;(A^fGX9.>f10]GNDFGY1]UL61&#:?R&<AK2aeL@WOdC3Z3+FP@JR7bAfMX2F\dL
7CFTC:bSS0Bd\b^+eE\+,;=9+Z#cKaRb^W1AIYQ[9T]=Oe>C[7O>TJBd&e[OY@PN
fg3N,g-KMY][JQ.EP4[e)MGFQPc#@FZQB;.(#13K>J,_BMd4/]cIQ(;b=<Q8_5TM
3dDV3=WODS#6YPP/(=6?<BfbNY2R8cOc2L=9GU84_[Ba)L-\&GeJJ-Y>2/]??d^-
SI/37,[g8O]d6Q#,K&Db4ea5/AY,?,6fgN&+68EA\,=U3@X_19N)-BSd\T4C5dDU
]1J4\[QP(A^=:;BN4RK(Y8f>KQ+Lg-ORVO9Z1BQdaDY=3QdJ#E8>2]:aa;dCLU+(
IbM&34=7gg,EHZYH#aUTgg@RT5TBg110IF7S0MNc,S(:FLM<O>B^OXZ[=5KZ/BQf
A7Y5M&TSG?)YV[/:2f88GSOfMI/B2WNK.W)PXM\&NdgbDcUQ;cCRTMV]X(7):g]Q
b=\Ob#OHa49:<d.@Y,\87#/gU>=S@F_3+/H5D1\YMB;c74)=J>fYE@M4@@Cg\>EH
&Y\<Lf@0-F,ZR9>aA0P):KPMBIT:+H/UITI]#ROO(QV-W]ARL>(44;8^fb@0H\bg
@D>AbJ@Ye]Y5/PBS+7e2GO1Z,G89??=4M,3(/b2NLA0f\2Q^B8I(V6+E0f-=K0O-
Q<A4;/QMF\<c8f+c_[UB0T-7.:Cb2P(3aGLS,B-,KKeLa2R2-L=VZ9bI0=?5:TUT
a[e/QPX)<KZ]7,0G39[H#T21K+_55gJf2e[^O>.1g&Kb5)V7R2+#S(f(0F^We1\=
<6gT_T1d.?Df.QdPFV<W&<YZ6cQdCd]]#K/O\5V_4DLgRc_eK(R;0A7PW#d6,H&S
EKUbC)&;0c4&;-W&3JP_^/1);X],\.N2;8(1><W9);;H@Me)&/4gcLQc[I?Z\U>?
)<._(7UV(0T.NS<D<=-08XHO+4dccK5\YL8_I[05/>O,[#VG&\<Q)_MS5=7F_H]/
^+VDV[STX1LPMR0@/?BYeNUV[A4DL<WD2:#;:VRMU=DY8L4;J#:=D^3B6NOX-<,B
YAE#MdC7fR?LJ)97_Nb@C51,1?\^DA?(C\0.BPd]LDdWbg#:PLeGa)BeaaI&#G#>
Cd?8DQ-cX=VXQM-bI:[0=CZ--B]04&fI0#[9FU:X?aGf7]0,K)Dc@;W^3:d8M2[e
0&2XB\;K0&V5+H4K1=L_?0_WJ?W4?5Q+2ZQ@Bc)VWI:44AO>De?J[9-XZ73#Y7Pa
=3RO-Z10FMBc7[,NcA3fYf5UO#8;@S5]@L_S#L4):UCaAD]+d[Le+F(LNS\FTa/#
N-,4\+KcBg/bJ6YBY4D9La1E;Ha3D=C6ND+=N/-6dK-J7OZW/O-XA4B9TIWcFA5e
,KCJP#N)-??HQ@\(=OQP(.FfZ1,TO1XPQ/OOP/GB8-,d/H[4740KBF:Zf5/aNX1B
b1NdA8>&:8J:];HX65V8YX,/&_KRee&@-Jac.)MT:^Z4^fJPcd\MaA6=QJU]H5DV
&_&.^LVR?9G\Qg>\::1?T^8UN&0dUVHPGPIU^Cbd.VeDIXgP./-Y6Q>SBb8@CSb[
IGWOD,6)/?I6Y=BX_X5IG3)\,>VOG6:;+XW.PHg:e0+C>[Yd7XI&a><Y#=OZI?#)
c1?=e0M>/bQ.#>3/>)TR1;V8GaX/5gQTE)QN,f6>(WBDW4?_B/P0BacWcb3e0a?P
Sdc.JK05[/><X>FNW<@]&,aW=>4,3a=gdIbGd^dSDK7Fd#]T50#U,6CE2dH46aU=
;SYB5O#74UB-5-Ybg?I=PY7OCg\#L5[4dMf]9MeI?dOFf.\F@_<9GCc5EU17_.QT
^>\>=J\5KX#Sf(V0,X4UN:[6LS)M_V&0IR_Z(Q?25AR.]>R>R)^KDW)SY(^@fT)A
cIWLW6CQY4].O11bgdGVJZ.,_F7]N]/9WYPc>;X;gQY&#PI)4YEMaBUKQ5Ua)eBD
F#R2S#E.2cMQ+.UdG>ZfafNW8SgaM9XG=cI?gB@_4b.=7)cYZ85_;-W-BU#\FVG-
J@\f]8,&)GJEOCBR4[P]&#gf[T1(FI^;?]cRb-UM3d6)f>@DgU8&>M_/A0<39/;^
B?]@01G(TLC81JY6O^46DGP]f,/NDGK]Cbb8C:ad+:?a74(B9:8J?QMTR[7cW:]K
dMI=5e@:O(=2Z[A\L0QeL:96IcPPDTL-cbF/(2M@HcY&;ZKK)=@-GQ+7EK\LBV@;
/A0DeY=UD)BVW78@]44eZQ0SVXFNZgEdP?-.?VS[73AL[7MAU)GBfQ-H4?GTac>@
]9UUXULbEY19N3V4DQJOeES#7&8V-W8M_7_8bPMNV)?bLC0cJ_)28dbAgP2I2)CC
QTgOERG@@]6+.g87&J=@cMAZ;:^RVbYB&:WTO7Sa^fe/DBVH6-+\;[g\Td+?bUeX
:C6aU-O4CL^?,Y:#d&4:;H4H@BO]#58AY9gdeOUOR,83V6cLK#@VL_,#FX,N.f@E
:@KG0_-+CKXUgQg_M_/W&AJ;IV3Xg2H)_WJTA>Cf6JSNcfZ=UfMS2eK&&HOBB-\\
@Re:.ODfKAdc^@=#COJTC;.P^gJZ;?CO#Qd+ORHCR_dg)AZTd0[/M>+R@^8C7,4C
NT)R(G/@S\b9,;a9OLBM&-P\LD=;1ITLYY_,,E0&A5XHNJHL_+\EU6@DI,R4?\GW
I#_?Kd&3A9Cf1OH1JSb?Y=(7ReN_Pa+&fIG^CT=1\:QUTGL;JD;?<]Y7SAf.OCC8
FH-1[HO955@I#C3D<GHeYaGI+<f4_WAF,E/H1gK7\<[G4J>gO[Q]BV6J9f?H^V#=
A;2C2_718Z&7a?9@RWQKDc&,:#/1NVXW&:)](XT?]1+.\F[aT7RF3O&>-];ZbTb<
AH+7=.<=S5AcY9V0C@3JAQ9<_K3SbP,@&DFee/dH3Mb>f_]gDB5HZZ3fL@=YPU/N
?<e<.@&J1aCJLb>HIIYEIM4QODKcOYZdD;HD&#N,^Q2ZSNN:-2_H,,7Ob,Cf/NM4
[0gMYR[B)[ZSSO#:RDgPW)0(K2H7d@)Z_#]W9LY_6F7,Q))4;>H(43Q?SHOcO0L<
F.9^>ga](ZAf9AWf<;MBE_UV:>9<e1L-fHRA<6G.ZgPc4]\IDC36d:5W,-03[^2M
EB:G55RK<1aD=\585_++8L-cX#0@?O3>ZHMRUTU6f-M_a[G6XDe5;b&8TY<L):Bb
Q1X\HZHXU[>=ZeJ;I.>L9V;=IEa02a^1^-\TE+fL.:3QN].0QI6e,=A6\364,/SQ
b7PX-=+-F7,00I_&BG:C^RR473,-_XV,0&IVLV9EY3YRN/+S8-:JYYHMLGf@B5MQ
=O1502U#fXHgSAF[\0e3C(B=[F>c[UC3-/Zb(8gPKI#T<eTVWD_(Q&fNX_HO-N^2
PGaa\@eQ=0OcJ3d+Qb+H.7OUF@5,)YEO35YW4+__a4O2?Vc5GPCE92Z>#\TQFECf
G<0HC,=0,Je=I-QeG>UfYYg)L&+5?/3A\c7;B>5b/B=7^ALC#(K6S?Eee^0a\e[E
5/+;W]3NeG>HCR7A6J1gcOfJ(NCb3/AWG6a<QCR#SEZ](V6b9d?^^bV,7R,L]Ic#
cD/<Vfg7P[gRXU)=VF\<ZITW#Q,LJgQ4dEbDJ8+_-eS<0T\abfTb;M>Ag;-L;9^g
Mg83a<R?9afYccAae/IA5c:/_J^HO/>PR43<W7,gHQ]06fe2](_MHc0\V6D6,WV[
3JACN50J):59_ad:(KWB8(6c>^+H8c:KM;-BG2[;@O.HU]FQ8289cGK2HfG5cY?O
TY^^4](d=^b/N[_,_8SL:4V82PE8bIb&_QH=U-V1X8)GedP:=@L&TT&YD4FUDJ(\
dW<9X\7(:&X=.Tgd>DB4c[]41E/a0g@SB_[?P99gT8MAIZa7V_c[&VWTg^cC15bd
H=)HO+2;;^K6E?RVcQ35X6:C#PXfDg>=C]R#Y:;KfN?@QW-Q&ca^4Q9V.R\((YUL
=f7Q2)g@-LRR/K,V8C41DH&fB_OU.=L4QK;&bA+<#<I)864a6UJ1#K=640M1Ie&^
fO/dTNLS:6Na\fdZHZ4fT#A.6Q6BGO,T(NIK0aeJ&@[+U)[,bOe<NQZP/dcW2=c[
I@7RW<#7S&F14E=<R(,JXSHeP_c1CSB#2NF8\7DNW-g42,A4KF#CC<PW9JEE<Vc=
:fK,KE67>dSTV5fVA<<=F/\eS-@.7&)3Q;PW9:G;^:Y(=fEXEP35.IR3&1BNTC@L
OL-IP[U4;),\^/7;aR#>R+D25-\LC-\]:91N)T&/J0.3dWRcCC7f)K@0G+:cE8<c
2aQ@.;6L>&-cXGM[L0GATE0@T:5;Zd4[+(YF/:XS:PLTfadQQ4Z]X=L-\@fQ0#V/
X3Y5cMWe13]KT(:YQJIXSa/,C,c1#T8:ZJ,K]c50BOTf:G_I7+1/=C\)VUW:d5Ic
S?&N;3(9V-L5MgG\_ODXc-4A,/=EgC6]ELEA?0We?.\M4.+P>Q1MAd^JJOP^Y+?>
N3QIc?DO5;T#=9.P#Y2Dc:TPF.;#6a2B+-SS45.L38>aM23A#Q10U)0[[6PX1Db=
FLXQT&5>0Qc9XY^L+K_\a284g8b6e&2#9We&b/)HAPTa?US,YW^c39V_O7F;5P3+
[KM0.4a3]>0BC9J1]R>OT4X\Je7EB+TBQWF/?DE6gS(Z:QW#bD+Z=(>aZ1Y[d?e=
TJ0^WWd(cLS)[2E+A\F;616e/49c^BPb8/69YOK-WETUcW.2M]WV@&2[eUKR<QH9
Pf21Bd8P-Y,Zc?5IPa^\dAH-I1RaZL+,a7ELFJBUfX9E<<0(,1YdYDHESRO5eCR+
M)35[8CLWV^I+;9@C6-C[2R)eB3>I&G>Wb[MIe\2U+bR<)\5UJCXb2IAAKV<VC0Y
B-)fOFCR3DWYD38X6W1)ZXCgDF.D)1fZE?\d463.3YKEA<JZ4P41P-Nf\F#EJ02;
BI&>YS9a2]NP27?K--;T.0KIK51]YBJ=^?_aTA]J+6NR)#Ia)Rc<3f<UeHQ8,7^;
91H)1Xeb6&5_FP)KBO02?\4/gTf(WI>VC;Y.LaG\QHLLUZH&f@>=M@d3.]c&RDbL
X]aGH.fZ_GG^?4=:VgeKQT(I<#e?@.&@IJBcQ9HIbBBY[DOPBeK_B]f),(-Q0+_E
XC^c[9(<a8dUSS?SI/@ET_U^4-ePCb+(X]gZd;9SdQc7FWV2aLEgVX6>9B8U,-__
7M;,G]c=a(CH3@Fc-(A2gIgdOa]>5=L_P[&A4fU8V,=U:\\/<:,0</aF3gAB=22P
e^2,JMHN71WbMLg)+XQZaC;Q7_Ve;)Fd_8X\C12OSTQ@;)P-8]G4H?7E6455?+9_
]R/LA1=7/Y.-G)(,64O\1U#dP)5\HL(c:K_-ES(d2bQG/Zga<=&2+^,L?>/Oc9F3
T.4S3H;BEF/3<3AdNO?[\\+]5FS/UeBDS^GPAX#N6NCE]2(@(gONHcXSL+9<YU<&
J)V>SO6fMD#BLWF>d;1EN4P3?&V?)gWc>HL?ITH\MBBRGCW]=OK_Q=T&@.[BSDaE
4I130@A@UdD+:3(dgS^BQR&4]+CQ?T4-B2=Pf[VR1Ra#eXRU#YE9->@0Ra9M5e]#
AI3^&J<P+-4eJP[-<c\[e5.5(+[(3O&-^&/]EK+F;P4OU681IK]6^Na5g_>B8<<T
R<YeUd>LAOZ5AFU+I9741e[X<\WL;\=]5\XL)(^,>W-WSf]-[5ZM]TaL6RId).[K
&JcU.Jf-L2KO&Tg)+Ab,@6&3V=S/045E87ZR35C[Z1?X>Fg3DF(I9U/)\5gC)VN<
dTF+NG;dL[ANA(TG5Z(ND>baQdL&08K]HN3=PGc0eP,RP2_7g<DQ6+R35&+(P+Ob
3JNBMED,^1QA<UA?=VZ/F@V_@(_9J^FSM149-:4SW2f^0^Y:29N+^6Z.IS_WIQX^
g)GHaEWZS+DT]+[BJg48fSL,]T@?fCLP\&6H=HLK61O9_/<\gB10NW105DXaE7H(
/I38A45eeK8=Q.?_.bLHf/[O5>ANF;^8==C/>\OZ8(T4@KK[13V\]I#B>=S&J6H3
RW\cMK:J[+X=e?@00;NOE9f;UPF9RHQBUV<YdcdLaN76[/gY)@M0:TB64J/U:27T
&_GC8S]UINfg#S=VN\49XJ_0@975d-Z9\7LFMFeC-NFa:_+.R[KH>cLEa1fBEQ3O
<;H2Pd5]1D^LZdDDdAP@R_a(VQD,3S\&2.\>WCI5CVXENC[[dL>)+E[SFG-8:96c
(PWV9]g(c>BaLfG(c062S,=d8CKeYN4XBY-;8,e\K,@9U]8?:2)U4,,\G+KG0c[#
SI:[S#2]=EUQ=.>N3Re(R[CW[2)a=c/f1IA<ac(Q_;eQg8LFX80^F,D)3R.>gX[?
ZGdUB^H-Yd(Z0SV;Ed^R)<-L^Ja.NS8PDJV(Yb&W<P>9BP1BJP:AX\A>gA?3;1a]
N<;NJ(7+)]C619fK\3ae4N>)3]N;;.Z2H##ZDLTU#2&KRF8eB]]#C75OW#2DXZ_c
fA65Bd;1UGZO8F4If_#41EG7R/,2>YHH76MaF1)#VF,VCe)#eOEdc2VJT4a6RRZ,
O4F_RNca>U0UEa/?2OU]1d)#9[,eC,NQ34C\AQcF@B?0=dP,HEDK9KXe0<I7SB,:
/Q#>,JO79KN9aZQ8,c[Eg>VQD8C6,b[RIIAA@CIX=@XQIO2OR6/ed7ZU36S7U]XR
Ya<gW][?;AO4_4-TBIKH[L?cMES.,_5[&4[G^-G43X]L^T+.N<,\8^Db<SXZF&V0
Cg7@0JMH+AL?PZK83CIF3@?IH>c=b/5;HEP9gXa.e<R0&LOD#)^WB(;]7[@1@<RC
1,P,P,.?IW4/767-BY^DYgGO([e5-0(5a>VQZN,H\a&V?S9_D&,#O0EHZ]HF7b=(
&8H;<Me@N0GH@Dc4&JN;\b=T50g&A0]Q=[UF&BW>CJgJ89_dW.41@/L7UK^Gd-DJ
IALY>F+G-A\JIX-UgTAaQF?N&.O^:bdb_YLJ56D>_0BH1+bPGDA#c[HdaB5Y\dJb
-=E&.3aX.7@;?0O,N;.PK@&+7O_DJ92BROR09bHIe-[76Ue]Qdd1^Z:SWY,L#e3N
L1b[6)6@S.@7C;(>9gQ)I\JYbfT3eJ7+1WV(HB+E_OK;be1NG/f@If-0dB2OV?45
DaRVLgAT))H-&4H-=V2VDYDHB(;^(S0M_[=CJa/A0XcLWZT,;2I=0H+<AQU7d.M(
2U_d5@9Ne&?c[R<?c11U8L=)5Z0cS?bBR_UR+/F+IdAg6GHX#2NdA11[>2SR3M8;
KNE6gdKgO&GJ<-<8#aX:4bFb@/8594K:cA-X+4Y[f>LB@=>G5^]KQ1JUdO+2#:.I
WDPCc6+91U(Z^&:=1FFJ3EU)F1c,W.I[+fA^(5O.-1DY?E>]C:PTDKC3(&1cBL_(
+9>M0_5PD<O]+YJ8N@4g_O>6ZT,UHFE1KBXUI>SdIf:_fSG<-(C,Kd8:J0+GU@R.
A=Q)[+b(>[V3^4[Be+^57TcRK-U^7d[>Y@>&:Ia6OD3Q,3bS>aLNaX:Vc1L.(5fI
Ia>94_C4KL;Q<fMJ?Ke>SEER-]>XeI_<>,NB@)2e8\KR)PNN^UN/TVa7aX,R&P0Z
KIO@V,39a_C9Y>=,MfBHGL7FP^0fC&^COZZ4dbFP1&S<KYD]:3;40-]I<[CTC?I=
,F3FL6bX_c[Id1B7LNU1VO#8;P@5dVAK.F?3)3Y8X-WW&+-:3NA+@.5XLOGSO6Q9
a-@bS]3);]>M;OPO]dO)Q^Z3[TN^0NbG1<_S8/1?.^^gWd3DfS\0=5?8d+II+6RJ
4T0gV@?[&>>CLMVQRK4<#eAB(DW#aJ8H)2/_2\VX]6\1(A]LeZ.-4,5&XD:E>=#,
Q;Z#JB/aAW,/Q42VLPI4A==[H,]KK1+PI,aMQd1OD0_UB)S<^#+<)&Ybc(Ye4gFQ
\a_Qg[\aMS\H\7SfV(T6,@O8T3OY#UW&WJ()\O[O@>##@f@\_1#9-6I2G,7S?R:7
(3K.BGE<-C\MS?Kdc>=.;.7496/[M@BHRW93D()@d^OSL,DcT=M&93Y:<E18>YHA
3_36cVe+@),?bV<7/CN0VQgK\2+.D665G5[-C&?[L6X4:/T[#2\VV(b&8gf):0O9
0dT+gLI4OLSd^A9ZL.=\aMXGY_:520E-K7\H>dSPOZ2#H2/5:[XT,e95#a[HZ6^#
FQRY1XCf<egL#VM.gQfg<NB;RFIMUW;PO_U59IX/39EeJTId^W;_PL]A9ac&B0Q;
FJJ+Le-GD4_QV<3-IN6H2J\<8\PYDB(2b]O(<8PAY>M<P?2[]&>?-;???\D@+CH<
G&&Kd]&AJ;<Y+]JFLO<Q2?[05HK;K\8=<$
`endprotected

`protected
@bDNYe;+;W70a]SAPUcG&^8CE/@WReMN6,-daV=YP6TSP6DA+Ya-,)WF+&E@UH:P
1O76#>S<HF@XGBAQO5RH.>X8Q9=CAY2+H_1CRYY86.5A.=6[:B;fDC4&7b\>c@a?
0gL<Q,g=D5<_UGdJ(BVFZ(Ia_/7S6?QVTV7@5K)E>ZMK7Z@3)3@>6ZAZPdYMOZQM
Q>MJN.V#H;a_Q1K;+QZ8R,aNB0C[4&^+B@\;MD+\D\V;44e@,Hb0fgAZP$
`endprotected
      
//vcs_lic_vip_protect
  `protected
KQd/,4\EX[@Q.4/fFd=:__65K8W.6+?]/IA9D##KAHNKC8[=O,)L((#VbQ[&abS8
7^:b&C_KeD?Z4UH@13F;4_U=:CUM?a[/7@M8/3T)CaKVFb:K9>/V09\:c140eZBQ
K0,cFJ=+:3e;&;#U/6#E0(VH3?HIDSV<@:1-0LPK>3K4ZYI9?J(F/#4[4)>a2#d#
=NO4(.JcYKf\:S1V@,2>^4YX9[OAAR[[M,6Wf+cZ;b#,P^BT8#ec-=93IGCM&<(^
+dCUbL]&Y,RB]1MJdJ,:#RfYRNJ):cFQ)1VF+Oc#>0D?fA9,Sf69&f<NOQHaA,@K
AQJ)RT2gce-.@Q=ZO08bTJg_7U;0dGQe#LaSc6bYa(2Pa:1;@dH[^725YTHc&AL=
6<f,XVNCWN^=eJeQXfI[/I[+:;@I[?_Bg?gL,^QdR?@6\:#VC5:X6A+9)2G[VTXW
?4H+>FaZLgX&RFVWdad3M@I)aRHZ=#6[5<U[L5XNT</Zaf2RD3BLR/RS<T;dO)&K
/]VM7J8D7\SRgO9>D/OY<]Qc;8(A3+gF5#+Q[L+ae]=7I;/YIXC&&4Ma+RgQ31_^
Q3ZJPANQMg)(--5]34M60(XbU9/4;9<WATZGY4OgD5Ka9ZceU_7Bg=B]UPU<:.GH
IF;>4PO41,K?U4Y7L[]T5cg@MDG0?P-/B(JH32DL^Sc-M(2Z]cMKfUB#2B\-Z3O8
NP]>2.U?L[OCe/GaCK.0X@d^\R#YY<(P63V9P]I>5Ig/OQd7,INT,XcLPJ#AcLO4
C@Y_L1Wd27P1_5\gY);Za:7L1\]O?geH8YGWJTSS2gAb)(S539QS.;Hd,>>:M7D3
TE&DgGO-77CO&PH5)f]3SXM_afW..Bd4.V6:>OA25fN41LMc;MW+H.E/UU\<:W\/
Qg+X?RM^b[efME(4aWE/\P349GG(Y(BdY/#S8M+9#7^IBX5<HT=2XO;GW@&R2T4M
W.)A,4]4U<&g8_6GE;&M<VfP5QG=EbL.O?S1[0GJTaU+CLW]?>ST:S?EDIbWOSNG
T;=P&YV,5JE\G/U38a,@Y+,9EcdcE,IVH7XLJ2R.QMOdRHa-,R4W1(b_Y(EES16H
]gQcb>KC0>Pd13SSZK9[?OK7IK.2)K9R1VJ8X(&[+E8-5#CO4^WZPG87Q?(.E+UW
]N^-,L7BO,_84(GUWDd?CNN3&Sc:.3WLIbP&=GLL27KZZCT6@-c00,/3@UD_P@M.
,O9#WBADVA6-8cFE_-/<,d3T(Wg1@[-S#K-1K@/[@cWRSKQTVe2\J2M60(^L?6b/
]1[M.N7.SbBM2_<>&F\K5gX6K_@_Q]WcL]ZYC=@K2NP(Z\>FLNM)S&OgQ:5R(3JQ
aPS<&bVdXNHL,8VYOfN&(X84^=RM/.6,?7C6R&B@H9Ad_D/>A.\]7e@2IKbb;1&e
f-^+J,,VD4;W&PI?P:1-N)P9C665OF;DFL@:W<Q-BS(XE+cF(@;(AQ4TMaW?Da7I
U(e>2Q4P?;(-Fg/T\#4fbAJBaI4SCPO0aTRYZ.7HNYTS(bd_VW:EWa(J9f0Z2#6-
(UZ>25F=8WObLAM5<SU^-5G16P0]0E1([64\)7MU(ObTMUe,e;I0QT<Q7^;:P-5c
D]<6=+KE8cWV(+-+W^([UTgcfKLT\_1ZFTBL)7WK8B2YZBB_QNXYNX;J::L]M;EC
2+bX[J3[/\5/XCbAWB8PGQTP1a,\cE6X&B&/Z@T119S0_1b([^C\]9[+FD858HR<
?-9;D5?cXe7E=,B0BJO>,UG8N?<cJYFRSGAM/B;@<(H,Z-9BWaeed#.-R3(V\+#]
VcJ6[Z+4?:SE3L+\.#@[DF1Ha<3OC^GH9CDC?J_YRTCO<]cED)LMcU#,=4Ia&@gP
JYVIQ4,Z)Xe:g3H4,72C[H6/@C9:E+GDG8_M)RKQX[HB&?cSPb[L4;9VCbR#DD9)
a-:F?1LM-N_9HZd;9\Y8I;+,[GKXFE<3:JK3Z\IY6GD4RI;bT,WWL<86GU/VJD4G
.R_MfX)L7^:gd2E,+J>^cC-GfAO67(Ze_LE\(WPE5d(Z:A2Y:<&G@W\9IU_;RJ+d
0:MWU&B6).+d-9ON3<([2&+7XKMVc-YBVC(D+Z[+6463Gfb4HMdG5/fd@2cP^3d&
GJX6H3c94H>\KZ^=+-aEDWbSf[-88D<0a#BBZ?;;bcK6H.PZfS8,+R9@KC\g5@.7
/2EXCgbfO(?>\bRdJ#;X^0LJ0g/N_Re:8--beGY9RV_14539]NJg[7F3a;SPVA,0
)@H[.[SG;+SN;1H@EWG?^cV\e]\PJI9gAR2^)TJKeaG[P5SAZ3;VP72=[bc1Yf#X
>b_KZX[Pd6aUfF4e1/8R0g5C9gM(4P2AgS^+Y?7e[VfC\HaSH.?#R13EG\\[/-OD
=_E.<OK=/;USa?dI@2Y\LGY0HaNdAe3+/_4A.;]BFA9=-I(g,Y1)AOJH^PW<#d?(
ED&]\,K==<,A)E)\D-8^P9OReL1/B/?:HdI[aU1)<;Z5/]7AbRO.0<e=6HXHE_d&
fDWZD;f4a-F1]E[eR.:XCU\[S@]Eb_JX.58TOMK)a+XL;8597EJH#bE&ABdM2g6#
BKJGb?G1FeW4SM@>.9,/=eEC_QK0^8fCK93(f]&dU5S.^7-+UGT<D>:/A@?T2eIf
a_RAXT3;5CM2RY&)6=dVYGeD]d?WJ?[d[C)K61KUUBd,g1]KU34[9QgX.-4J=?5-
\9,\LCC@TRgUU@,MEQ:fNJ+eU1\,gT.X9/VN)1EX+eg[g16-+-TY>Ca0>cBCWOK0
dXSJO]+D,a>Dc5eJ<GeDgYL913cc,)<DHV6FNXY&W3)TEK?^9Gdcd05M?.FRV+..
IgVBZ\eU6\/<UVf12R(Y00;H\S:(9HR3U<R4OgN17@+.A3\WVg\B8^M60&VRQ#[&
?3A3WH]^Q7E@X.f]<.,HQQ\BD8[C/09/;?M/^/VfU6U[:c(1:bI0R>DB/FX>dH?8
)@<^J>)[:S<WTc?ORYN^W)>VdUU^;V8F,dO@27#RMJdD.7N48>/YS/<XAJIEK^c0
?WL3DfVZ\4f=VCaNYGNUB>E+W[I29H]5eaeHQ#VAIECW<,2/dZZ,TJ85>>-#a7(Z
K77C5=S(LR3>Cd5/NeZ@/K:&#ef]NT\B_KG4J=[\J43)/86D#f,QA?\)JHR,IK1[
5^(5CQDggN/ZdQ]/R<^8+>\.E<dPM+9:gNNY:V.QN8Hcb/&F02CLHB(W,1R\J^Q;
B&ScC)NaF@3NU;@ZIZ).NQ6.0HJS2d^9&[Ra0O#E[-@@PJ:ND58AE-;ED580<WLC
H3>7gWeAZ>T(>;D<Xg^3U?SI.#1-O_[DPI70AJHN,cY-&b)<B,dA83e4c53RS4WQ
?AV2GeVEJ/U2OW1#WQg3]1<I?7BXXO9]0+\;^bb<O\3dBM4?Z1[7UENFC7P;]N9@
D27U.NA-C[O@T,5=-g^4U33)AbRXQ?\fB7,W<^YSVQ5WOg^fZ47RVT5?b6)O4PO6
M-)^PXDSLPI+)L9G<-97<<AO[&ge?ECP8cHf[MN<EK:(cR#1JS.V^CZ+cA0(K+aT
5/9ZKee,Q;_A-XR,2[HOQ33g8Wf+1/0(<F^:/=G@#&dMff_ZF5R/7N-HU2_1f,2e
D)Qg=M]5R#P7E;Q1ZORQ9N,0=5.Edgc@H\+gUUB7EX+2T69@,F1_#8a6-eCcd\/C
K6U8[@<:Za+1?)S]&-;2>K,I+2g.-BB]3-3g<M^874]R2JTVf#2Q&1NCK[5>31A;
g7F;&0cDY8Q<8S;9gM,=V6b5#++(B(HX)Q>O<V#Kd.PZ:P[VD-6G@TJ15c=?W=\:
Y3(U[C,KZSU[Z^S?()a=O;A1B?]<V8WUV>Qae3Y4E/<]ECL?I\:I&U^K8\@_<H#<
a;L6?86(ZN^JN+Z3-Y[VN@B7RaDQ.SLX8Me&@;VD6M>]fc@B4IgI?b0ZDEXcUcR\
]3U,KY^VUOK^\fN#XPg^gU#NW>DMH6^.S/7+LP^_J&@,ZIB@:6ZN/X>.\gQDRHEW
,:W?X6X4ZDgA-3YQWNHe;Y_F=MP_=&-FA7efRFL#e;OCGKMg9799^R8e\MM&EAeU
>]BgB-b[C5NgC0fV^^11)O=ROg^/C-?_=[H,UbOPa&2[D_<[?J1.D<60M)FH,>92
YO.)M77/g&H0?E;5a>#94-HeKeUJ,+R9H3>g<R5L1TC3(-=aQ-]gb06>ag:91,#b
3bT;,e_eTDF@);M>b9T84(\c+MX9])?+/;_#,S+]P<@^^RD.+cNXC(-(FF9@Z>5N
?1a90QNO1?C4#O7FETQXg^Z_LK_T^aH0?@:LKCZ\#4P&Q6O#]8U;/32X=^P3M/#O
CeFcXD:+Of_C?/EW@]4Q]c][D()CQH[MJcP(+c93Jef=9GQPKG0Y?;359a+aL9F4
_^TXg7<X,?]]OSgO&3bOOg>,R@AcM):/V3b2cN<IA-PPg(dS<JR.O?^4NU@gH#XW
J2^VMZ(76KYcb_0d_D+4f/LG.SLXdgMf^6DU=@2IBdPM]FPKOLDMJN1=8DFYV?0]
aXa,^?HDd_#0=I7<JIRaQ+73C6=,,-0>bK,E=WWW2&,)O4XeOMSc_(/S4Rb(7+DX
\SD2].WL9;1.=7&>cA6KKY(+[</C91-9\YffQ\VSFaY9?/5XF;)C1-<JJVc8Ufe;
-]ObPS3Bg^EL=GAY#:.TdI&2]&J?R.IPU^5P5#G:Q_,/31R](Z.c;IS#F6LRTc[W
dU+gG]O24F8^KXgf-GWc4M_,M^=dMZY#7&)R,Y68I9_>_EEQOgL\/NM=://?\94.
I>EJPcM]5eGN<XY0b[_fO8DN-7)E1._J=>.9KEZWO)CR,aQU/EQ/0Db]Z\U7E]<O
8<f-GV_WDJKCV6c(7:4\A[79B)L8WI<NS_NIYX7N<3(P:JZ87<8]G[b:.47]+(0P
]SL&P<]:L&A8=0.0V]CZTY<>]YOcU+6LKFJC1TDPFL:Fb63L^/:\.1RY)TK0)<cC
fZ[-a&@()..+H0QdV_R9@fYFdTCF\>9WO003<0;W=(.REbEFEEZ^HZE7>V[+U8]a
e&9X.W6.-Z6UN,SBYN&95G?6BW+\&B^dK;?ZOS6&7F^@4&7e)eFQf4O9-4=4-,TO
ZcEPPKab?;I;5=8#5]D&ZZFZ_A@3Lg<L1H+@]1;H/<K\.KbWGRC@806&#8c+RW(S
FQGGd7TNHQT=fU+1.HPHO3(;b]YBeZQ03>-_6&a)1\@8C3(eDZeE]B)b)RVB>b_[
OW(4D\-eFZ>8g0VE?Y@-La#@Dgd/3EO_XYM<e^D/<1BdN98_HU]QNKe6=_I:.cQb
XQQ6FgROgbc)JXO2X+8[&C>SBCcfg31;^7[<K:OJ7LT]NVRW6QZ^[eS&PaY)?FHI
LKS6KWE1@WdRUH.OLM9I=QMbJ;C156Md=ER+_.(XXB//@K3;QJWKfSS-75AC53aG
L=-;:)dCKeZf97,[(Abg&bT=>]&FK;ERa\Y<+b;ba]9D[D:QLCBCAb0F:<HNI#:1
Lb8I.2SSa\-C1@8<cZ3a9OFU)@(51#eFJ\=]-LBGON>bJ:d2ObBd8-K\P_B08C1I
K7MU9cPS3CX^.R\.D&?2O:D=,LcE5eC2F@bCD[MVO@2G3F[g2SI-KfWVDF5W>91W
CFHT=X)1g^992O5WE_Ec,LBf@7B(ABL&=BUOe:AB/b-7BR1gKV61;c)cFN3K5/gR
JZ<4<S-,-R1ACdR)B(_:KGS738<6Uac^0;M?E3Pca+#GKc^6dK_+>#bIe<_?PEaO
:0=_Cd4YS/.&,+J<2S?CTcW<#I6ASE/\7e3HSbYBPa=D()8L4cDSJ,UXPdIE4RMa
6OTHc4@DYXT7G/>F^Ba?c^@2I;H7>1K=DEf<VHR3X,_X9)5Q40Y(87b(FT\G;DBG
,>6bJ6c+Kcc&FJfI?LDO\R?80K.B)_&UL6GQXYUIN)fC^]9YBVF.(API]CC5Y^3b
8\M)GK##N-UO)>29[J0533:T3\VQ7N>CW8PNV-):bf9bCcCV5QF/PLRD[XC/V_0E
0d8;f++]I8;3JQW6^\d:WZ>T>>FEY)d/_FC;6b1T#I&E&YVC/3L77eK/-bU);T8F
68TWaWEUd3:/;LD=J6[O1@?(EbOFNK@4CR54RZ>1#=)<KgR94TWX^2b[GEg2@?T_
#,SgL(MLN#\BR&X_b)?GYLNBd[-f2_KJOJ@aCW+BH\EN@<79:_+BUDb6(->T:5[K
Q&JFYaQf5HA^a<1(YfL3d(=C#9c6>^-A)-];b_0:&4Ib6K:,YdD7JL\CO56Y-#0>
16&+9G0[-PT_\I>9&Q.2TF0PN?8>,bRT>M0f-IV5\R)5)R;XZ21a9,[XVYC4A41@
/+6-.f^\RG__PZ,CYgW0g()-Gb,;Y3_&597UaIQ)?WdBL\77CHU]N;G>Z;A3=X\P
Z,=4IB+0c70G+@W,HARc;?7;fL[LMT\\>:17+aO,ENSdEc7I+(D/S)a&OSWf65L,
S=>,S3S&^,,Kf8^V[?bI\+&W-IZU<<LN,GIQ8X>/#)D;.e+3H2B=8?3[6:O,5@>.
cDE_6@V91;P>6F4VM8?I3^8[fSYMV8b;W/)=gR]N3,TbK8.^<^U+;Y4=cV;NcAD-
DBEf6aD2XLfOc[T4=Cd^g<^_BM[:6=4[3gK/;U>=d/c7\U\c?IY[2U;D<5-C6Fg]
+P05E1X.cRWFEG1J1fPa#SD-WabaMg=L[7TW+]G,d\K[:8\@KK@c=__7EZFHZ\XK
7a75K?g3a[>SC7+bLP+_XISO?OKY:3J1:-_V0;T5?]I5.fB^6-L5O(.YTa.@E?cI
]1]cKVX1cJP;.:RVLRf4XW;]8BO_)MPY,2S(;+(>0:ecc8X7>2\>I0,-Xf:gOc+\
OGC4AX:I^^#./X-B#S)UQ-W0\IAJDe7>C=@Y]:2PAY6<V:1O&ZR_7MNZ6,J189D#
WYbOJb0fN=LU,SWE>+:8./.WS5_O<<3T]]Y^Ye(Ze=@X^F<+H,JG&36e^O.7[GHf
_@)c1=7V/E_/S>8(@JE29(&0QBH:N6:Z/IRMMR[HAD8]W248<K;Q0+a-D>RJLQdS
;3&Ha^NFe=E]KF0]EYQ4NgAM1][R-M?X;WZ;?dCf,I3K2;I4/]W5/d31O(5^f5;(
#@Gcf<EBg;?;,DBI95R_HQgVPCW(^e@3M]:e)N-^CZcdFgJ&?[_a0W]Cf)FbI)B?
#N+c<c:9.X=D3TV9=fCSM=cLeeH&R_>)6X@JXUDN/;RGSVeb5A.W4#\Z?C1XbP@?
/3&d^;b[KY6#G6T.<9C@4QRDf4+aN++/:;.<)VA/Y^5:9_A5AgL=++F7U.0fKcbL
W-X@:+0)W):^IXEAO1^3Y)TS+#eUT+e48a[L#0Y]-TK]KR=2UFR)6Bf(\ab(6;7=
3ZF5aKR<?44TVU\;X,Q&T9W(>#R;b+TFG0.gZPZFAcVL,G>E)_ccMI5(_Y]3(.AM
Q#[M&Ae^6<+W8P)d]-3HHA.&>#b<g^2Xg61M.bTIU^1I1;X2H>HS;_M9T:Ab:C0[
#WYSXI7.CB]YPVB\O+-b4R0MfR),FdVR3(-20H#LcE,W#_@[<9YIETFS2C?Bb0,:
PL;^VT@e&#/1_M8#&,HgT1:^;9#]WD_Y8/4d;UM,\SP2;7TAcL>:Aa+CG>Q7b\;&
J1ENP3dD0YH3=\,C0T7Q_;E?)R0cTfU9?@Z_&<W:8V]#VG(>LWI2#=_2\HQV\)Rd
7+0ac/Rg4&QB6J&<eaD?9;5:IO5066U+3[&Zb]1_C8P2XX(a.VU22J=<4/29VD3[
K.,N2L<2V99BNcXCab;1[Q,^e21@e5C9e1@G?P)D\#K=3Je5CXPYCVE4.edb1KaD
?CXSJ1J,D/-Z)>;:KH.GN01)GE(M,-W+.#E.6&FR#9RL>K.g.dT6FA55)<8V&)E:
V0f3eK]NJF7/)GXc]Y9W[M->aG:-gH40YL=I-b_3WRLZ7&2,5^S]U8_E<EZ1E8_6
<N^VX&@.?e7L3G&f57XZ\&-3^eFQT3D)G:DX83VLD@8#6AWUaQAUEDE7R).>VZgJ
647QQgd\?_OC\:#T0C3;1ODfN&NYc?,g>7AD1L:G^6dMBgcT0LI[^<cS<+W(Q@51
B/J\Ra5^<)SI<H^(,W8UDUCQ[MQYd#^0K55:A-b=(P6Md,c?;(C5)(#B_G473IJ9
PE#D:KO;]Q[dZ=-OI8N?b97?@[+;+f,+M\\g,>T7Agf.&Z^>-F]JMgaaN?I[cL_,
G\=&-#G0<T28)T8SQ;.SI+7=N5b^WN+/SDcK##cN3=>5g?R_-3ed>A,MN]4DW\M(
?J37.4VDD#U@DI5N=0MOM1\[2H621^TPC2\+EXE9N=+gI&R9DSL?b_0AF2=7D5ZP
+HgSfIOa56?3.=Yb7ZaGbII_I(aA_E(@5SLUUe4-D6,M+4T2_MfVP)Z13E7J56;D
g,/D58\dIZJF-^=HB7EcU9J3\7\V&JCAA@TTBcKG-g[#,O/<:b/=,cTXZ<TFU>Aa
,=;4+<1M_S;E&bd2e;c?AAC)07(N@1QFB420?7e5(](FQa_e^J#bbWMI.6#PF@X5
Qe/CWQL-GO)c]]3EBK:(->/&SXUXSf;Hcb+FJ_79I[F#]OW-gbY3g9&F.bN?Ld)X
=OYb>KGN,IHAXKDENK,[g\FRf>Z)f,D8T544351K@(P&OP-(A:^Z(S6B?]>0Q<(f
efcZ5X@WP,G)GI9M-ANeZ[2Na5)dE8MgKN.Q>>>(AV3)(aV)b<Rb=DLCb&b3cVZ<
NM]beMNFXU:B/HdPP3e(Y[GD9,EFg\d+GcQcFHR+b<T<ZOQ+a[1T)9gCM&)\-ZKL
)I<79@96H2eWFZFKU4+g5#7.K4Qed[:G[^#LJ_Bf0F?]=cUT&L\K4-V0&cAGJFKU
7^F@P3-)BcDJ-24Ub?:U?[PbO.:5WeW).E_dg+_@aP;6gb6EA)HV[TEQ@^#-RASY
CZ./9VZ8+W<N&\6e0c7:a>LGQJ/d_8@d<8Ld,Gf6c@90..aS.?.@2=b6?Q(BABYG
fI+RF&6Y?1M6YdK?&)aKe?c45c._d[FAX4BPfcN&J@R<[I.4BTVBP[?)GY:3Z7YQ
FG>#UJH:6;/c=L2)cX38f@8B1.2^[9dAfYbDf[Ef#,/.=-NGD810_3=YEZDE/QU9
6Cf0-:TeVSV^D+Y@QVPYTZ,fDTGEd#^)F/L[6P7cO\E#^=TE;,6IUIM7AA895OOa
aE(4O&0=8<+a?b0g1Q>Q+;>56U_U55HKZg,).^.V?:0YYF4-Ua,L5fU,9)-:36b3
1R[>(=^g/M9P\?0=VRDDeMCU^6UJc7L<)Aa9AP;JIW+EM,</DL?;A6aS7e6G4[_H
4D1><&+g^fRgF.T)UIb<W1_(^=HZ)31Ga,K)gX,0?e4X]T3WO&A,^@]]1@C52S=P
5dJ/.#Y(AJWVBMGg+d\F=QfbCEMEYDFVPgPfaa82ER<>N<BGaa:J3M]VWa\&7L,M
dZE_dd:Q@)H,&]G\dJD\Ng55F6)=(VG2JN+dK&Jg+4C-74]/3]fg\:ED\]YI=X>Z
5T/;Cg77dE2eBE3>GTUDG_QDD&=#O?10ZX4O2K1UB1V\7RdALAbB3DaO=?Dc<J0N
#<[QZO>A7NIM=>E?V\UTJQa]EX:AO>;--IZPWdBHAfJ#e:HF4NRCP=a?&/GFTd>J
4@:[AN2EJb:bb.#3dN&Z-K05OUb(AQABc1^&Q0TUUc&V97QUZ&AJ23:a.^47JVP^
E[8TGS9OF2J5df-52;ARAfB?W?TMA7-c6\&[[=a_-4,HUL((]6L>/\8H@>6OEJ^(
SGa6Yf9^gc?f>[(ZE:.5U[+KAa^-<?Y4P#UILH\OYM7\]?4&4K?X]e2/Qg?)=P(2
aS]fYc2+@a8FFU<O9TRZ0AGW;?O#XC\53QNGRdeO->E(F>ESg9]\,->3K^JS/cc8
VXDAP.SKH-c/g(?KYP>V,2<C<cE554^\GP7GEZ&UX]H4VFQ-Y@+-#.WeI<\\YP7Q
5\c]_\bUJ0MabT1cc.afHS7_L,,a@3ca_[@-efC,ORML=aPL_2Ng0@XEFR2Y3aDD
[&fN<<7>YdE=gFXTY]RX=,g5e=3+&<\MLO41g?^L3Q?ZP1-HRTV&X>[[D=I1M=0)
-TQ@JNXI&2^)<WF1ggZ:J48JE3cC^T\NBD/0BUIRX+5<b(6CJ[8geP@:L;K?bC[8
:Q4L=6C/O^=QF6Y:)P71&JAC6<>FSTHJM3C=ec.e]8E=?XM#cP5M6WDd]P:5HI14
5cYg@NgZ_[<\+B3aA+eQfJ49c.ZJ:0f<@#B1WI:[2E)d(4\VBeU9e+R_a+]IQKL2
^E/KL7\9[(4MOf034eSce5G&F2KQZ71-b;?CG\GN7+77.Q(53_IaK=;3_(_3@5F_
2K4GV]8_&S2UcHDA/1JI5bCbLF&=?(f@#G\7CB@G6e,85dM0B\1cPdVN3KA-9/8?
e,b_LX_L_d2@_:[7WFJ(<1fDcQ2WNI?RM1N7OOcQ;?JGU,(AgIZK,I?80T2[5DTT
a3@;@Q^7ac8_TB>-)ATWMC2J77#@3_.58I]ff-T5.ABd)Red5.fBaOOL&DR#Da8@
UECdY_e-2L3]Y3(T5EWP3g9MbbT6Tf2EP\P_0X#I5A)QLVH-UQ(K3)ObB2a#Pc1.
@J4=eQ3MKP@Y)LCPBC=:;7Ib:#\J9F;bZJK(#7@=K[PK)D0>=_843,Bfg_29cG>2
3?5I?EE3g&C&TNb#/M;+<_FgGdW,R[?VeeDTf_6L7e7/fcK_F[c-^][F@IXWC4@2
aLQ&E7\dRFAaHe1T4TY]2Gg-Q7^2HYO.BP&)[Pg-&g2;g>MbY:7bP(JH)UZ\SREK
9a@<T(S:PZ];9X79]aE=:YI@85KV/C\X.-gC+MQ#LC)Z3[36U#B#5Lg<W-NXO6^H
AgM>#-5g0\[)Ra,8(??g[Z=(N:_28G0Dg+;G66][dFHD,;\b31LFG@&-M]L?^[b4
^+d0gDORa\>FW]?KO[8GFZfUT8JdS6f-gg9fQVP]B2aE.(2A^>WU:LgXa5HO_(aM
PO=-;<YM575E<DPY-e_W<(a/Z0H(#\2XRCZ2.[0Jf4490PCTF<:2L57YE@5Zc<)7
90QD/IPX3W855BAKbU0:05V=WgW&-NYa/,.YW]dd=baV>>I-PI1J?:d];/(]+H_O
E_._IV2PALB#A=;_0)XN+8WB\GUC5QA)K\:>J]SA84_g>1KC,9ea1_3L^E#QU#a7
A>RJf2SIF->1<;)Q:9aEMOM]Q2L978Wg5\H8)FRM.PCeEYgRXOHRYB5H_-@5DT4^
E4;KV@4I_P#K01E.+1;8VL0=BF7Z\W9Cd+5U4[c2FbW:6eK\EPag,QeJ@5IKbbM_
Q\@\c?8CUAKS:)C#6Z1bH?R\>DT/.CF(2(R#HUNUdCA7D5YeMY1e-1=1LS.;R=Ee
HP/K8Y.b,TG\0N7+7M2aFA8PPb=O[DaN3P8e2T34d6/QL5T9JTD>MRHMY+WM3Rdb
d2RKARR8-W\2CKT7Z:3AGZ?,U&[P>Y4(B02OWSTcMeE5SH=b<59V-#-DCJ]G(WV8
e+;J+VQKAO(&B0].5@MCS=18]AV833IPFE)N:R.7_>F0Eb9+,^)<X9J8da?Q25&J
0DVXfQDA59L>:7ZGY,@5SPQUT<6[NLSB&:C:T<[cTI.e[T@d3:Z\KAce781--S,:
0.]1X[&)N21FDK5cBfM#2:RA344/)=g&_6OXS/RRRYCZ.@NPb_?+)TR.\R+gfZ_9
2XV(gS#dWHSa>Z\HMg7:8Y7F^cRYWT[F6fa&0U-(^c<3.;4A\4)UIFOe[Q=QCOMZ
AH\f:3=)+E\;C[>8X;CHG?QCTcZ8YP\X5\LAce):5F42EV/d^;^CG)V4D20?NOH@
QB_./b80C(2PeVJVZe)CX:).H3/I>_#XV&W1([CJP5BW7BP2,<Q[7S,#H/357^TU
G7TN.WfV3Z6,^VA:gHXf7a4R>>,_A9db?D8.3FT>e0:G>?Y(J.#)#91]4_9YCHB:
RG>]50[@(e6[;L#Y[\7K<\@>@:OH,[gA<A\I;e,708P70W&:_f/9)Z6MW1-?9+7X
>;\(4O>Z9[<=a#[Fa05UT>,>Uba3,7TVWA=C]6]PcHdG^]QgWYR]WOg89T#SNYTV
KFD@MS?JAS6C>>ULJ0#V2d=,._(@QFaf6_II:V>BC43P;]UNP7c4\)4_\C3e>9MN
AK@<E<_S+Oa?SOBg3F:ZBZTZGLeFL2_@CJaK]D#907P=eP(5a;GePPY\+O>&Ec5O
d(E43cZ,fIYH[;TK;:cPV8>PJ89KH&BIe.?K;aLe:DBaW;6c70=Y?[?_:UO;K?8T
8_]1Z)Y(c^WBZMFNMJNa0F/&7YC@@OHJ(LWK:8HI)e&3K_LR8[&FeFU,T1N@b@&J
OMSOSCGL3f,\C.]<))RJ(^:28e&=>E7N-5N_:b_6HY[^M_f&6D+-IZbDF5c-BebN
7&);C(/1.;658?GKV-.e,(/-U7->:LHb(#2F5>aL:/Ue>F->&?M+2cR-EN[Hc7;<
\6ZS9DY4NBaU]@,)VOX]fOX#5c(f(]gP9FURX[Kb6@d_Wg3[ee)eEgK>N)0Z7?:K
TO/5Vc,<F:4;<OAD=^\UVI=d6b=>TD-<97f].HVKS8Wd7-H)3+\Z6T>EY:>-W?TM
Y#A0:8ATYga42N>^9.@5-)RW-9>&LVMfD[I;8X_I9c^b-=.?K\1&;PT-]/VW^R@]
[Ta>#-ERZ)a<6;K4D;C5UCVIZaCF6d(T9B/NP2DFODf7U#_X(eNT0O0JUP<cTKZS
?cH_M5=[,A,7Z=\7\b_O6[]=(6CA&)-O;8\VVZKL&g;E(_>_2R,^F^[2YMa(<e>I
+eJ4MC=4Y&d[Q.5-/Ed)IRUY>=1KQJXP.\]X.^H-<9>0dE;eNM4S3d6KC^7d^?0\
3J__&T0ERLJOE>@MZ;#1UJ]Wf[_)7D>BFS:7RLgR3;+T[dR/9)6F^)/ebF)BV2TS
H1UUG(b/#ZEb.5XA9B3;+[))7CF.31Cbfec1J\H(#G^R[XC]D.d\#O259FNPf:SQ
/SAJaQ[f/XH#=C^_HJ;YN0U0aDdC.9geGRVBS\W_=SgE/5&>A(5(D0VQgIT#,H5?
^\cYH]R=B1QL;VdKVF\?Q^M4/@59e\(/1]?:<UP(ZR4[Q3/HdOL(;.ec>=1^&96+
P#+:IIV.I[)[8.C#dA,gXX36@MH<I?,BDKOHL8CQJR^M8(XHZd+a;8MV]3_AI\Ab
<WRW4DK,@Ce^J)+KIQDLWIN4:;bZSF)[6&ARJ9:GTUSOUaWeXO;;5+bGG\>SNI,=
N/Ea9NLX6)PScIUbC?DE6H8S7C9d9-#8AC7P(=)MVeDGQ?Ba5_eUH[Y\S=>,T5:6
X/AaJM#_UQ^_.P)cHJ#KFT>V;OAESL5?_0#;cVF]O\g7b:C91E)ecMF\JdX@?Y+)
/EGCR<.UZQ-7J1>EM_43:/=W>.:fe>:AU,(RBW8G^56/_f&WP[QSE/d\_:+MUXDW
))2@M\OE9FU,OFA9M&>P0dSV,bL:3HVbdN6I=\bEQ91[7[g^1.,H7OTKKbXND7M9
#gbWP+O(HZZ?:C]:WQIK>FG7E_]M9L66#\RK)<,9a>b(5?H-H,YK67Nd(M,F6M@P
;E6<-2Dg9K573I,gTAT[:H-O7e;E2Vc#UA([=>8J.[#,_R;HPJV4F+RJY(\X/G52
R?G4T5760Q<cTPbNL(Xd11([N]O_F:WG>cVgVU<9gMVE9S_J);6-GB&JC?R3QP&K
<:KWI,(5^B/RESc(dP.+3I-7WQL\M[/V(54KVFY+V1ab8&ENIBSL09O3OKPNFTC#
=^:A>B3d>Wd)37A?,[3K-P1)eAaHW:NZJLJBVVb87PM_\/ZX;X+CbW@C=J?_KN2<
;>ZLK)-J,L<M=XfJXY5I\#6MML38MI7;DE(L2;:P(^2^dT.^0;1ICAJ+OSVP81GA
9A4^TKd/P1/a2-AATLJ.>?W)ML5Q==01R4WJB/Y#2=MHe<T47I5.<#Xa4NQY</:0
(R>]I9=#JTE-7R5E72N4fb=V2P=faXGYL748d((,-0=5=,9WQ&Y<_EHf<XW-?Y?V
^M-ZS4JJ26&:8e3Mf)Ha3A0;W.QE8#GfMJ)WJ\BZ4ZAHK<C0F5DABcN3aU<F?M,U
3d3ceR@fU8K^3D.,7aTcc@,Z\EDYCIA<[T7=?cB98RdC><<UIUa^g@];KLT/HH/N
]X&eK(IF-ABUd9MM.0FXeO@da.HaNAB]>GPE)DF/>0.U?OL+D0KM\<OC?Lf28B7Y
8]EV1C556L>=\&JZP;5\]c7EGB&(<HGXM7a&AO-OX:1gPWf)RBJd=CBR3>&FLLVK
Q?>AJ7B_WB;Ib?53(DI7_@6Kd_52C;A]XQ>b&2^JG-4-\K^?\Hd9+=C9\P+]7BDP
JML?]PbFbP/58be2,H-+GD<_aRAa1XJEb:QX(P]WBX-4,/?cJD/5/U?)95d2dPeH
O:1MKE8-?:f+?[,^&?I/P[2)aB/A0?L_La0]D@5FANS+QCKe4:P-/7)C/[LUBfe)
B.QJ3EYA;II0XW2)J?ZPR.c^=Eg8I&Obg]_?TbA3<a>\DT_A)1TA3Uf+,H9MbJ86
]@>HFBLPcJ:2X]:0B<G)NJIV4>L@Vf[KT\#@bSQ@+aMW(/M+b4aa6aNFN99C?D:]
JB4KH(W@\E#W]06GN&I+-NaQ=6AHKQ;b>7Vc\3DfaJ6,gL8M?b3b-XeQ=ZE4YbfX
2HaD]K\&_VW:_L8KE7/R?LCJ&Z7[KaY7Z,^^_DQMEO)H3bVE0?;5#[Y1]-;]:eZU
#&e:3ZY:g=SE?@6J_2?Z-Y:_0XaL>gTPTIReJ6A(GEEF;FPbe;aeW_;A0N@V6A7#
+5B0U@f[HOg0/F3/?XM]ATHS]<7[RPMYJ;O:IQV2+Sf-=-A<L&\T7M&PNBe]AcdN
T.O63PA2[^ESR@(?5BFM^S.02]QRK+^E+3G>HTTd+WOMV6@(fC/RIG7-9aO:KHU=
HC?Jf.7=[&<9M9IcX_?BZ.eUME<41PP.,37B:WZ;/>F:SSS31ag]G;S)(ef6N]I&
.WECPMIGNd.\>8)6@H/3SK#:R9gVL9)G[XFcQ]2&<fb+L[UC?<a@;81X4AA(9,]C
Wb96T[Na5GR[bO8Q5VB>70MM_VODZU>daB^#9?(_FLIREg,2cU]=U2(ac=#fLQ63
b?fNK^/S^b82_=fQ]Y])6QDEAR(YMOQ:;\([a]#T[KTQQ=?3[V^Q6:EH?CG]dM/M
AdE?VR=F97Q]/b<b/EY1_)=Q)5]7AR8)2e(GYa9P@8QA6S1I8QV@&U(T7LLJOFW<
I:<5TNEd45R204V0Z-U48(/bcQW5[?b9ddgAP&G:T/XCeYTGGT7\EfNBVHZ:V&3>
9DFP4_fS77X1_Y8:DWG8FU&f[S-11a0Nf:+217CLL=-JS:3KeF)c_T/f/PM7OTY(
[RD5;^1.QN?1O/4gd>L/&D4)WIB6A]#Of;IP9bQ<@,#H=>bCX6&^]PL(Be@9=0:O
DHIMT>&(_D#U:ecT1ENW5-Ba=+=IG4G[PL.0?^B:9J[^SPbNg8\.-4ITC/1,N(_E
1g6Iaf&RP09@XfJJC]U=-4<3QQZ7]STU:;#:34GB64N@/WE;Xa0#DP@]OUSdcHO^
-&2)HD&H.aZcPTTQcQYcIJ.,a)G<=:c:.X7e>fUH^_1MRH3#KG-]/?1E6@P)Pc_Y
H6YZ3^\M:RW<3=-;^]e,O0?_S=@PF5;L&G(4a9PcJ:P0TRO>2,^GY3c]O@:[&)C@
HJI@KAFD0CKI.6RW&1Df_Ae6f,Cc,5<+cUg_J],H\27TCbE[/^A<Bc)7F+?Oa=+Y
@03AW.KB.@<PP1_e;_=_g@A9:H#IcUKJ)W?M_BKf>>BR].-B&8B)GM_V>8^U]DAJ
bd0\g13-GKg05/;#<:bVBYI(N_>4X.dW?Hadf)dA&Q3KU_N@]W3JV]G+W_UA&1I;
TD\bbICfOc7F@U&F]DU\6<;9>))&AQ-&+<]89TI[N\7Lc?=dBC1CSY4T_\J,.PDb
TIDI:).UG/5,bDQQ^\[Y:7T;[<Ka(DDdU4S[75SI29gfCJ.\-6)+]Vf#X)T@^Y=G
D=cD;3GLD2NS];a<KPND\72BDP9M-7TYC#4R.R<=F\,1V5BCLVaT0dS5]aJ5YT>X
@cMBB>34T1@T9DE1=f#K@dDKTH2Y+9Dff9DKW/@ZK2R(GQIg5f,VL8(IJ<GPWY7A
H5K_N8??IGD9C-F8&H<+80d5?,2g:Z11(JZB[X39KX01;^(FV0WN@;LOCS;949>T
[U1E4AHgKK;C2#1TV5B9V<a?#f&G0D&IPJ2=W--D08A#J/f#]MeQ84<Q);OY8bEX
^4C@\-==)gDg@FA#-\HX.dNO-VSW?(6Y;FZMUQK06dPTBQI2MB-R0[BbA4)-Y=6:
PDM&Q[H^\Y=LNR@K5AbFfOEOM_[2-[&V=)J;IE6()AE_>+RS\J\[/0+UDM(Y;+1E
DM^&,V4Y@E?LUCKD8M_CKZ&IRT;d/F(7@,AY/gW3-_efTN=\D9\>b?=g;MN@EFGP
S)N=50MX\A1>@,-L<e#USRe^O[>7;72V1.9@/d+1\Acb-9Y8BL0ec.9RD-_7c_Fc
HR5\c(S7H:P@faT8g4YR7[TFP[9aCKb.;^e4^997/0#Y\]IDU2b)-\J7d0G>fDF=
B[<LK4P;9V]A9XWf5B;[URAfA]_dLZ(CX\B]GMaNJ5JUC]FeR)g1=f5DLVZ@KKNa
-f6DKQ_Ng1EK0WLFMPV\QbG6\GTD-JD9_&D@+@MQ3OSMd6W^Rf3fB<JHWH<^gB-a
<:XM@A,Ggc6H0G/S#8DY]+@=A#77c()TB?0f.#5H-0.7C4U9=egS)WP>)b?9IYT9
]A5>,dB?8/A@aP>W4f3>\>\6e_-5B<_C@e++@#=>LAb[I4?/.<](TYVTJ:JD.54K
1eMOb(U#P^8e0@TJb)Z27Ia.gF\[;-&/4,\<9LHaVTZ:-9N,+da9,9c<4#GE>DI2
W:_H3#Y;Q+AW,ETfISYaE1EGe;KDI<5D0PMLG:#@.6BEJL\/=3YHI6(D0aZM2;BL
CG<>-S>C8B_)[X&,5;[DO2B?5)NJI0J7;WS@&=g91M[f9@7CaRD,EX,eM#f9\IY<
O77e[=XOdK+F-XTR)(]:J7b>O>.T</6a-X,P0V3gFF]F)?X:FEUUDXWg;J1c6E-]
:HaM7S@.AR<9:1UW,>Y09A6HbbYBPNND62^9H_1UQJPa=ACc=_.gTd^7CD+#>P=Y
&&PW)TU2&Nd<^T/Z0[98[fB\;ULAgfQ;CW5]DUfTL-9@&c6V1aA;[@W4XA7(QGV^
H16RGZ@4)@6@V\,eLVD6Lb.54)J>f.)LH9B@HCA<7B<SNDdEG;&FH2f+b_bfcI8e
@K,R/UH#AVgcLIP;CVf2GNEBQ(&_+QW&PF[1)YAfV&3&4&UW:^c0[OZ17>5G;?X6
_NR0>gca==Y3[9OZJ\eT)?R^7=0I:@g:,M2\L[=9a=fW3VfgSD?L;@Y#N\<0a6R&
=d9gUB+A5N0-H-,<#N2-4@H_,fL\<Dg#K+L4DQg#MP=B&\7=We7(bgF3US]EZB0-
e^2-YE?#Gca9Y5a\)O6UA>+L>[T-=@WYF#I.=R:+7CJSPSJbF?[8)\RH?4)JYHgL
Hc\JMESd@KHV[##YS3dSY2<bNf815e<G@KO,HOffU8HJERC-2aFG:1092:,gZNg\
N&=WDYa/[Lc<gJD<G?@OJ:UM@-J34NAS0N#WC^gXF1WK.]2bdg#G+^-\bKNQ&Q7-
fd+M03.,4IMGaHdWX8R6\F.NQQ)+fMIR8KgZLN95[+4DZ[I.Kd<LJ,6XCd8YZ>[;
0YAVR]#_(ffC/fH]&30IgH0BL[7I/f0Bb:@J2f/<N_D\;>KROaeD#K@[SV\9;6SJ
N]BS_]HB6d^b#e#Dg97N/8C59CaK@6[DG\<<E^XFY1R.7MgfCAQG&Y=?<GKW^+C1
-8T=]K]A>+<c\PCS5ABRc_RZ,\LJ=cW(aYOA]BOW_03L5D].&0?7geg87.C/WMbd
5^0,g)0)6KR2H-a:77+/g&D(Dbf.ZTe6Eg5:bA6LINQU-S<1#faJ[<Pg/J./C0)#
:H7UR.eT.RF_C;&]V+CL:K2_1fPNJIN;?=JTIdBeX9)_RSJA7&.BF/P^D..<:,#D
DKN9:7;O@3@@K,JJRXVQc(;19_N&d=XYDY_MO1,M2XFPZ8ZR+34M-XNSdUD7V:MA
^AgP4R0>f5[6&dV4acYOQM#,5/@-)L9fDJO_R[&LU(4H(O:5,-4ZLdadUd4E\[C4
g[+PXO\XA3ED/f)(6<59A2d[4&D5N.J>U]8UAdT\?G>:.[-PS2BI\+V03,R=+&6X
B=M<b0MRF]Q6M9.Z0_@.WV#9b2S-^C.A8M(_&::-.Q@Z<BBS?-eQBRG[VS5L&K:-
_9g[dKeUc7\JR3RL0aPZb)CZG=[QY\+[8bdR2/GI7a1VVG5#CINHF;9.fU7?DBNa
\#^N?\EW8GN9.[PI?VNT5FF>^0[UKJCgAWf\M5TPDLRI]3E#aK.WL]QYa:O)BF=#
4<9H]?W5<<f(5;I3gVJL>]G07W_3D7\bO-;6O/<11UYK:=UO^PPdKJ0OC\R/BHd?
0U01IZ?(5=2E[<4dY#>U=cP/7,=S[_S>,73])Zbd[QE(E:]>^=^MW_cg0=8CTcCe
+SM&LLU>\PYU0eEg1b8/@eBIg>VafQXgD<8][PFM/77:(3L4-T<Sb@5VI1)U1T34
W^d8a;U7#P&;(SNQDYH5]\W7K\Bf#\[&+?V5dR]/9cQE(d7YQY0+/8#&eS5H)4(2
#dE;cE4Se\+TY7_a7e]6/?[Ff8OT0;R&AJ[+&.E]bN(/1IQ5?&&<T><PYAbWV8;8
]?Xa.;/^)Tf\Y@Fc>\JCfB+IbEcDVCX1FdP=@C>f3[8TS&&)?J\B28H>&6[6P(=O
Wa34b77-cI+f6CXc+UC=47:705W=C>DAI3NH=<Q=P)9@&RQ@G>XgKJ]MIUDB0(/,
-Z/cR-Kf#8\/VaW7+IZW:E)R3B9D)CN;#&&AIXA@MWQ8F7&[TUW,+,];GYf24XB1
03R7c#TN45RT)_Jg:;6E[14g(HGc6-HOYGPJEG?38UM#0EI:O22?:CX\;RV18gH?
W\N#Z:bRIT]1THMbdLB>/]AA/NQg4<_JO\O^RG8CP56gX1+fTABM&fW1]YE-aCIV
b59VGT@Fb:N4GdF7fdHR/)AdNc41g&VNDQ7.AW2S)&/#PW\=8^IV3VIaCM<<Y<()
C8JPL=3.TQ1^K^51]4AfN32-,7-S80K+Ga01ZQ,YXfe<5c4dL-g++b[=4@GUCW7K
f)#0ARgR@#L:f@R\SP>@#Ce38-fgIJ5KgX=VE3(HIG)Xc,,,LV7F7T)J6[5g_-W;
2FgNIa)(Lcaa^=)0(G/4ECRM@1O19SBbZc2/V0b3_O_UU/_(D+?0-\7JH,(6[e?3
1W3/+_a\V-gM_3JB<P;>&b^0=3Nf[aREcUE6S=3#.g[#?7bYeF6B/6)YYf^f]Hda
4V\)T4:@7HR.CWFAN6ad?+&O;07#bM;SH#_\)ZJd,g[B#d)5f_]<\OKX.4daU&dZ
=LHM3)(\1E],3#6dP7,2>1ZQ.L<D#JQD1L97Ra,2_NI8cRe5]IL>6+b:KKc61Cg[
85(R:e1^UK/?gA;Q0c_WL;_4&LeW3<<HNY=I<]AV:#5YB[ZOI@[C-ga-T]19&\-L
D@a-)>ZA_=5(fcW&:=3(XCX48P&UE?dQ(P?]1<,\GW1?T;8?BRc.I7O3+TD?>\;b
5YbbHU;bI?6Je#2KM/RaS(aL:WYTf:Q6#ST:C)/VZ,Y.d9-eMYa;P,dBTN<R1UIe
#W=Y;X]F_HFA&X&5493H.@A?[>.ceKgBaQI2U^SEGE]0Y^&c./F/<Af<,COF<:BZ
Lc:G41WJ9gfK1DBeg4F9SCAF8LbLKJS0f5#FH0BaR2e3^_f(X433?Z1TYg-V6a&f
SUEO&A:+S<@1>4e_5,O-JD8:d(JGSLST5?Cc3/6^9XZ0E68.fN+-B(VIV?)]fE5B
8#C4/QV,Y\0a[K=(cd\06[/^_2YRY/XaQMJI7BfH@JCR&W>;_Z>Ba?&_W5Y<@OZY
eA:d)\1HEF.[J=]N,U<g]d@ACDDVA:T/ZPf[&[[ZQ/T(.BANV313XcPEV86L5a/+
;c>JW.Wc7cZA-N&JN6L<?GS9.BR:Kd?3KE?gKKXRScb+C<=JS>J.<C\LEZ,6.PHe
=ff7+O[I:78<_gV?SgZ3LP:gMfD#C6@+5]P^FIZB=Z]F[CLXJ4ZKH=:4bBLI0V6K
.S-/ENJ8X0c@CL#J(>IS=AQMdIED\1V7A<5g902:7KNC07E88&d0Y+:T7eVg.K=@
@EI7I]&NOCONaTb-==:R(eG:YCA3MGX==Ua=S.PCfP]eVM+4),8<+2U+?[f#eF(/
U+Ea)g@H:N_E;T(BG(TA.:]f&G+e#]c]#^1Pb_[KX/?G2JN?\1gNMZ=^0LF.X\gV
KCaIWg(42E?J]db=aaDMUP0QP.U<#Ce/g.&Y6T6Z-MR/SHO=PEM<Rf5b,ZZX4:OP
dc:9.eHcY/R[N\V>GZ1Mg4g(_U[cDY;eAL@>#02_-;88.]AI^<fJRZ?@BT-e6>aN
G\?G5L<:,.c&I06cXf?&eYOfd>N)SJ3Ja+DGV9bU=^X//7[N6ggH1/97(X-gA.+?
HL@a>>UGEN^M&=P7ef\-LHYL]P:GGEB76GD;Aa&07G=VHP27/TbXD1T;+G8Y0]D8
.E/_-WHdYBXF73F.S/F,-CC2f7#2U_)(QU1^Y7/\BCLKC1>=6]6D^LL&-CG]g0.K
U)A#(Y]W_+_YLB5=<:V[S90431^VL@252>FGC:IfMT@C\P4DeDCfVX0ePT8\]Z@O
&;.U#eM[OKD&<f&<YB&[bgB3E0B2=:I-fRc5D68@/],g=bF=9<0dHSL?K28HH_;C
)?f)e]AcE4]X#WXEV9W3JbN&a-eR1b2Bf+DXC11QaeZ7:g,=>(@#-5eM=8ZRc-K_
#C=[F]<Y50M6AG_56:C]QT7I^bbMC(4fS]&2-6U;2AT67]>.1Oa:;MH/T=?#ENXH
<a[0Ya/UD^T0DM2cRG[=#L1JQR84G9^Z1[7R#H7?MHS+gbYZ;_5;;@#2HedE&V,H
#&Z>X6^=/W07:A84D?JO<_b5+S0Se:RO5IU8f8M0bK-YJ&7JZ--g95e/X\VdOP8A
fR40RPI(=d8PDf32Y@P7S:>-Id9XbOBIS?.RdS0a:KGGdP:[dUAG3(<]YPN(D6N#
>W@.J?fJBQW3KY7C?[M6WAfL:@HD96PC?.9<b;HRP(0<c--;W=fGa6Y-[bWFPT?N
#[-WSe0CREQ>7]3R7;(6#I>/E:\SA^K6Y_5OfL,<AE@[OHf4UTE)J&Wa\/d+;f<X
F5(#>PSS9=,DB5\T/,ZG<_[b?I[0F9C52DggL>H9IEUYdYg_fU8HZ;,FXMGeMTH.
4>0eJcEc#g?WJEQOLF@Y]>;^>DgaH::DF/bT;M7=:MZU<X>SVT#//@.]KN#2eeC,
HEGVF(3UV.ITbQQgD(8436V&?<5d3a[\N\W=8L-,J9<W=WQUYRQ>c#NHUV>=BM1#
Y(ZPB4TV&:;U2>ZQ.6G)834M48f\<?4O@JT5=1Ja)2F8B@,<(<6SDOV;F;.g6CH=
f]JYHF(0QWd:&U_Y0U60)SS]3Od^QcO0_I)?7I;HF:1W1Z=S?(8eUEPWc-Ze:DI&
1GSG,12d9F016M.+\ZAGT@=R^[ebMVCIH^8fKbf?M5L=U[f@f1>c^;ME94V_C2NT
AI\?Z@&Q=-ERG>H+/&ID[MF>2aSAJPYC_O_3E:LS0<JR8HgS>)<A7Ha/07-->5g1
TS+EGc)\:Kf_cI.T;:bLZHAbA3&+@15+<_F?DM(D_X8OT@c8YX@Y>EF[=GDD>E+2
.Z]NKC5)V4IT5HTLW\=?7dU.U8)8deU782;RYgT3E1Y-&3Q9T-G^IFY@SC;<1H\T
[0OGdSK/S4VKK]><NIZS]2KG&)B-6@WGN6M#V\<bCbeX0Q4e\c,UGE-8;00FOb^,
b(^-L2S/bNX01:(Z#d?I?,R^YDbT6E[=b<-N5\-:SCU]]QYDPefV.CT74NT2,BLF
N=,\S4()KcY/W]\Gc4<@]OEBV,WHFU;C6Z)K=FJ+dWO[eS8@O1RS8<,Jf@Y+)d.;
\DERD1+O:TPa4RP&c5C<eU(4Q04g<SV2?(d;aAcQa[N6\:.3_\)0U5I\aT-NaWe]
Rd3bM)O9[6W&#KfMH:1IaUNAE9,4D_6NH/@52@:[W-e-S6#:T^6C4KVeC(;B=F+K
2GU;f(XEbEcd7/4Ya,KTM,>f=5ZIMd<^TL=4LU83PSWgIBHQSAK16g9MCLA,a0e(
GX1PJW@PdfLdL7FP0OA:P^e5HDXAYUJ)9F5:G5@&Kg_bC9E(XNI&-<d<^,;aa@,.
/.R.]Z/3[,TDU_6\4\8],[#IZKZGV0B9Y8)f8J.OZH-DY_5cZg5=IT;60L1+5&)-
L)fSa[M/7JHaZ)8_d6eE=#G1ZEb3?SP>8(T)=71F+CF7Q]aObQW4P29-5Y73IQT(
5M_C;dC1^-1Z1AWGP@Lb1\P^KH_&[\cWDb.POO-?fM&e(d(4WT7Jga3G.KF0G61Q
ZHFUH-<fb9bUGC@7aD/,6I]\?8<W:_[5f910/^^^36X+4UO0EfQ\\B>(OAdWVQQA
3JS212Tc-[(3N@DE)G6UDKQH[Y<C.6SNbHR2Z(I>cP3^Y:K:Y),-MAG+YH8)DJ6a
)\a1KNd:2K#=G[=2O(/bGf/ZXTOC4-)eT[1,?0#\2ZI-IW3e1<9L]&K,-Td0gS.4
THJ\_2Z3L\QY/-HQQgN)d^ILBGJ^X7bSEG_NSFd8/79+_4)CAD?<75SS];)cUd:.
K6S>e@@BJE-B2^DL19c@d<e4PZH:K]F&,bNBf[1f_3.E3Y<DS)G:19AJE4La)S\J
ZIR82.:eM#OOc>KNPT:CM^\/eE(DK,95@<<-VHC0G::0(>4?RZ&\]@6Y(4KG]E,J
;<1R4WG8:.7SUE(U\7LOC@WZY^VLIQ4/CQJ1ge@/X2)VO.5[UBe-=Z>UXBbVQI#f
e3VVf9?.57#dZEW6dD,,E>DEgGL9VAH?[I4&]gAKcXASEN893R6)IdZ0K[B71.PE
-0?1;#=Ude54#@HdALSOIAdJ3>KX5f3M@4(-cg-OF?OL;6&49<Q/&cX<1N?gF12<
.gOBAQPZ19>7GTc-M&a7DKd)f>]RL.G=J#M/5RVaZe)K9X:_?b4.3CCMPQPLNg>E
2ZR>=LZ]=FP]>LaL#X:,5aL8\e(9Z0F]1=D_R@W-F4L@DI4[Bb_YF,YMHWA/:?B]
gG][,[?@JL,GY]DUJT@Z_3_MB2UbI\P2R@#T^91X<:Bb[M9N_R5ENP8WgfOL(IRe
-7F5TKc^H,UYH0TDebKUC-Q.cKGZXdcDKJ_77=R?[4YK[SaGW&[KG_5^X^_UI9=5
SQ>?J]Pd9Ge>./MMW<dFF#CR0fKQ&ga/T3RK5Rdg\#?e6[CUEgH4P.&\KR:CUcd.
,35HZMHXK\.fFI9H:A\LXD--:M<aRaP/MQ_T+OG&AUDO[Db16Ob@E5=)MfL/QRZ6
PAC2R?,A9M?Y7[bAC7\[g3,aa5/13gA)c^99>^SG@<I0U^U2)?dK6:V[S_6(S/^X
5^c>F4,Q.7)F7?b1;aIacW6G2ggf>2UGS,X)eJ5-#0<<,HOfTQK(D7-0XO9DC6G>
P/)YMAGd8O,NX\8.K>[W1gWV8AMT(JY)Q9UF/>4=&BUT^#d<_/>d->cRbfI-IZT_
9.gCH\T:_a1>-.=^dG2Y16&(1cF\Y57MgeL4ASbUFDfd7;O(gHW2C@(UC=E]Mc1g
B3WTPDEAB\\gVfeY)=,FGANH,OO9dNcX4c.5VR&0D;.6X[^158+75Z7R3BY/Ue.a
^XIaX5BCP8J8J)f(gK74fF9_O1MYI(.\-XE@UIe4PNZfL7+>_0)Eb&T<94E5E[ag
D<g0bgJY&?\dK)7N2(#B=MU:[_J#U,WQ5VGX=K&BM;Y-U9C:D-7g,JB+0Oe=JU@F
JJ#)1ffH6@bLf=d)[U;f=MVC@/)>S.D/HVS#Q^[4f4O#Qb15SA1/KAKC/[Y@S[fV
X5_;HPEFLHMN-D:\3I_1GD2077fKGCM3\QB9IOJEOdZUgK\&Vf.FM<B6X(e_YEI,
<96.-SM2)I+_27_WD7>Ga,S><3I\gC/5<E5=641b?GN?0IFA)B)XH@DN1FKe8/((
0MXO@7J[TZeLG/f8NCFK^MNSeHBG(cb+U&PfG=>a;dS64eE].+^]eV5_X2_9.5>T
KNI+21V+NCECS2W->IKgLJ&#SfSOF\8#(<FS?Q<<MbT+UPdE,]e^1W:T\H./?C^G
O;PZ#@S@F#E\E(X=]J5QgHVVcNC-COHc^<9+H2ZYU@UUM6;BL/B4_IKYgN-(KO[@
C>eF/d;S5;4L:.ePS_V;De8G>OA_JdcS@Of.,g-HWI(WS+LIFe;&(A=Fdd44BEeK
Qg9(G2E:36#NRU>,\&:B/EY3>feC#b\f<e1@(YOMJYH-deT:@J;7^T8AVKN(aM_2
Nf>U/=?L9V:>9XBPXbePW3QBD?gWR0)RaGHLX4OO17WZ48>Va;aZVC<)D#[Z/I.1
gRU3O>1MMfSDS+[,8&)?1Z=]fJ&9KH;P^<[T<#bNBb-#7Z\C(F)4?e&G2b=\JS;[
5L+>f3(E<_f)?#fIA)g&6K-8P,-U23I1(a&Z-0BP#PI=(:P.E6D419gIEcW_)WOf
V&N6C(g<0K&QFf>ZXFO8N44C)L\Xc=T:d-_9\Cd@4aAY)=KA/N_3B4#?9dN2>6YW
#AH\c#KA7HU([)VDO_]/+cJH1g4:CP;?](B+DU+(\SW3](R-?g2fA0Q@+OEHA@L0
<HD5gC&3UKI50Wg<+E/b[)CaK3ST=I7]b.]dP7fCL).TW;GbTPL-SLE,fW>g8D0L
:/HGQXgWS6//)F4d&#<N#I=bJeJ=Z4.^NF5M@e]<\):H#@+3I3-THCJ9ME+K1H6C
ZRFF3:J]g;.D;KK]QLT=V-)OR>=Kfc9POQO]b7NaV;;4\PN4g8GQN5b0D)EL\\2(
U2P/?Y17P(BJJTG>[A17,8_K=&Pce??FdJZWE@+&1B\a8V?5;/?NgRHJ7^[W3\:@
?C_6RW4&M_VJ]G]A:#4-#W0XZGZS:Sf8U.Z/+Ad/G<;4+f?AC=GXd]HX)7e?79+b
A@DQ2/.a=5MgKYR)[ES6):+c=J0b#(H8;Y^8?V.95NOTSbYP.e8@7\dS/C2QY?)b
5\&0aBV(TI_9_-6AYJC8-c_H29:g&2aIMXSNDGBcDYb;YI=V00N0dA0(>B(_)IJ^
6[(#2G[V3JH.f4CZ2W:#GM<DHa#JHRQSHe0M=Ec5Y@(W6VKFeW2OHUbN-MT#SGA[
-EOg836YNK35;2[[_UOX+#8gK<E<?+\^K_Z9aEg-[3Q2HdVe]6^BIMO0Y3RTd&@I
JWY13dVPVU(+IQ9N=N8g7:/,<@f2bfT?H);AN\K/a,4F6)7BGO-5Y(6MU=GGCZH_
R];6?Z^H:6cJ;7ND,+I77IQSY1d<;;S<^BS[>[81HRPYN-5:8STJ+E=82-I,V;9e
cM.Q,Q#KM\@W6&UE9+WPDQRC_&T)/e==\0Kf<+8DQ(WS&89DWU#ecS.6(82,:JCG
GNI2f/QR^ZeGVLP[G;5@ggFS/JE9:D8PW:8(:;>8G9J#_XI([EBVW(F1;;(:G-EJ
\J:U@aA4Vf#@.\3#V+@ZK@Ob44DD3,CFX?C^))C:T6@(:8&MJY&N.BAF?c=fM+G<
2U45O_9cJ(dOME+AS2XY]</KYC39-3N;:XfSC7aJRH(-+W?9AV8ae8UX2_dOYUZ:
E^/BD5;QE_RUI2R_6&JW7NT68bW8:4=[Y3JM.18R=[10FEYBME5@Z,<795OLAQ0A
<4g^/ACeHeKCLa>J9V^>5U7G3>;cW3D]^Q/4E,X:EHdRB5(2IIIGUE<Q<+W1ZR#[
G8Uf&f,6K+3W=aA[3V)25,a8.9_ccHKD3P-9&&fZS+<F/HYWZO0b]>[4?8RP62M.
YEgB\RF;93:(?1,S.\HbDX.(3B\-/aAA#7<7^F5W4[N8LFU;=\^Z[dT)1;F++;01
Ja3dJCe:O/0G(f[X?K9dTd=G>74,M9(d8>Q?F8>^42Z5^21Cc.&@-<9\?2E;OX25
2#Z70=NeK0]g(bDEX,?Zf.UB<dgGHL2&/dcGH_TZYKR3+9\cg)L>?BD;QXVg8IbO
\eP,G0+VdLMCYX3EM0E<<D\&eNCcB9JF\gY(W4C&QOY98(GMH9)Kg3O&&S6V1H-[
W(e)d)>?.]V[82DJ4X>T4geg>#KP/9.SVW>_\VFHM&ZLN5I#-LM:1JP0:Me2>/fR
<ccK1K6?cT8KVa87>af;a=;YgD_5##e5#]ec,.R8>NXe:A&#;<RecMgMa=B23/;4
[.45Dg+O4+RIX,;^9MY297gHZR)DS-<.K4WH.1=\d+#]dS;>2H_#gMLb#6?79?^D
T3D<X_^3A/\OH+4/>U)7PV;=[b^_[[.Y[e&VNd@YeeO#IRgRP?HR:_+7e_Nb:dNP
_gIbOU,V\/:fU&0P<22I(?.fEE0\YQ2cECA=_;<(bU3KHE>L?53IG?(,OH;Aa1C2
He;GUFTA9MTHfCcW_5TcgK/,R1.IeTF<X(_]fOD39_DgQ4fFL]?JH^J.(eRT)Q/+
@0#-&-LaPF4DOK9TE,G3=0P&?_9R^OV/8.^4P:VTTFRYY#b)>#..C5(Ib-5Q5O&9
EXcQ=;(_IMHDf0;S#IV4K\Z6U&AVI+d8><7\E0#9fCY&/IC:5-4Rd-TK0<+-bR3+
&:U0U\\c1RJ643C?TEPKG=7GYeLd\62;_;1,e8>J(JXN4U1R\IeGD2_1#HUBbS1d
1=#,.I;,X?LN=Ud@RN,J=/.F;/=K\e0@UPg^2UHW9E+:P3f@]18eS\OV_#c(Gg[Y
M,P6/P@e;8(8dQGQH5fHL-K=Cf<+]=MfE3@M,_ZT[Ae5LPc;OD1g[5[+fa@.M.=#
A2404P8_@^8_2CZ)+7-ZG<PH^MabKbXB19&+@7#V=]?@A74UTePDXBccM0a7Y+S=
2\38[a(5U0P?@.eee_O&O[4GFQ.Q9b#/MSHBegM3B]&+ZbE-1//[(5Y\@CfF2_;Y
2A+f\RQ=++_,RZYC(D6<H#CV#CN<V:HI<2M;\1PF/a<HEA-31)PC4INZDN[SK,7&
65T0YBAK0,UgR?M]D(6],Cc[++:TJ=PE86DR>B/QGQbKXS9Q-(Y7^T1aKJ_2)\Aa
()_0]X@-Yg4DIUV_RJg.XEE;\,E;WG^M5FLIX4R:f?57d&OT#M[-X=9,2g2\Nf9O
7@c#A<HPRIb6^b6?OQ4DV;V3Xc\LA2:]U<9?G;ZM5QF8<@9A4,&X[B7CZgJ-[2,#
_cYg5&7:L9EHb,@^E\>3P<@G^B3a8ZBD_;Ba[:T.<&\3)],ZZ-C-ASdDI?>9<ZQ]
V,b\9aF@4<&]OcV.I>U;3.;fGI2,QeLcbPYKf6R<)]7@a5N&&b=HV_e-cB-b\&Q)
9E63&TJPeDc_^XeM7W-V#)Z]^8ZJK6I1f1G=3>+Y\2GM^fbE&,O)d7==6e5IEP&.
L#X=)7IH4V/ab^#>7_>2dSESYc=E/(0Q@/U5D+DbL2Z?EZ1/=KW6S//0G;g^,U[C
[5VgfNC^ed?=4BYR(7T0<0@U3e>&A+14UT5?/WMIC7H0Y&.^NEQ1QcQ>Kc#/,.28
TYaD16Bg5;Xg[++f(G(.T.^.2_d>/bOMQT)5<?>GbcBMGU,OY(>g:NTc20dN;24@
93B@E1UP#A1&&;B2?]U1I\e2D-=5FXY<5JPHT,/eN(Q0H0.Y[<>IcMRd]5YcFHJM
@OS5DG9;I3@2\R)X+J6XJ\49_VFMNY6GKGF/3)ZIFO.ATKL<?-DP4.4V>-^/4:\\
7>A1-L@7X#_eJc^L25:CUV9]@J59gXd+E[^KX3,e_#cfQ8dC?(b6JE179LV27+9D
)(Y,Ge/:24L,/EGYHC<=H\9YC/E(77_.f[X5e3VR76Wf40RTC.&8.Ye+#6<:?9:9
7Fd.FNM<R10PSHME=OQHbKXa?)GWP5RLec2P,D[6Gg[Za?._];)P:\6@YeQQe>5Y
gZK4a2C9T2[ZQdA(N=;^-T<]bGUE9EQ5RRZXPgBc<.\0-K+X<R>M<+4JK86MFST&
FgB0WXK@OAb>Ke[/a+-&ENZA^3F0O1S,1T#d?3)4-2H=&<FBJ-]H7QBV1^H&0-;5
e71]I:)L3T_9500^:@)HX8L#KIcXab?W/TF5X5N/gU:a)ZH&J,D(fC;IgQ]]G^I?
)U^G1I/7e7I?KL5EBP@>)]/IA8OR8+@H;0cAa-[^?YQM1C9GM/c),I)]E)P6,1&N
SC<O(4N8(;g8bf-[1B:4J0:42ZLb8e=;Hb@4K.G93;0)Dg2UR;7,O:T_):]_JI@@
Wce\?3b89e&+)7MQBecbYfd+FAD<WUB#)=-1?U?DR<CY#+U[;C6P]\+]6>X<[b8O
\&\44N^Ed1,Y\=]9P91.9YY7aW\Z0^DDMMKQS^gPPP2+bK0GgPePGEW^6/;-//\&
CHe#Rb4+R_UZ;5)]<NYHI2].IB-;eT]K,;U/+:1)c/A-/J,L4F56g)MJ5@-,IK]4
.:&NKb^(:->VXeRLWHeTP8fI@\V3F^^c_I_^Q#9V2#\.0Q.88MO\XCK.-,(&/GS:
?cQ+6Q\e22HPZ]cH@gP9H/SJE]/G+0>H8101d8]6P1:4ND1a,)=GB67O(@ePMd8H
PJ3@9C.QB\\BbCHb.cFBSaBY.JHZ@(XTN+S3+Nd6=OCNc9W<Z?X5fK:<gQY73RG7
)/B-cM_(gb6fX0Q>:21>NG:2Td+F?Dc^8e4LcEDa)[(&2O5e5(a1MKL^5TO-[#:[
FQa:CG+^_<I3=Pb)5XA@KDKP8Af6/SZ61QVEH2KTfB]&G@0(LG-Rg_\PaZTSIa.@
\21(L49#AdJOBJ\c=TB7c-Z:eG.LX@<ge,(X3T?4/),A-)NQ_c1M<-f4D^Y]7ZUR
T6bR4]Bdf_[N-a-ZK0MD,]/NgW+VFM^F_O[__0N5PER/4K7T]#\>_Nf7_g7UKd:F
-a[TPHEc56d34>(C\Df3#\#eW3Hb;?cFG((HM8Y6<QF3[=7>Z(1gW-Y5U_IVP>cO
6O9F3OZ?F[5R4XG,M=BcKF;Q)C9a/]<S7R<W0,.V/d68[6X0[f:&X047==:@cRMg
R3&#Y&B#JZ/TDQ/d(7f@W:7.1R3WeIM8P7_<S9eZG_>GagAF\I\/,RaJ?Wg.DU</
TFA6,K97^3c_C-IV[ZeIf&fZPVR3HOG=T+\7BRXB5J<LNWFU<MQMP3)?A3#[]6@V
01;c5=b;a&:3JJbLa6Cc2DbWEfV>>R&.9FW>9OVGb)gT3+WCJ6A3g:N(8_X/V>],
b;X[NU&d#b;-7c48HHTX4&;Y@GQ-85/RC4W+9-T+@(ZG-&X(SYVHTTSJ_/RNJ^JY
8&(>+.2VGP[fM+e?I6g]]5f@B,1,@3HQ@]c:9&3&WTQEfgKTJ\a(?WF:.Z_MPT76
XDLaZ+HAG)cgRG4J6EM@_DKU[#N&.UEFAZI+=d_f8GYDK+K3Q35D&+GK;JGbY+Z<
Y7KP&M;B9EHVENNF;E)TdLFTZ8+fI/#RHgV<P&U@GF53K+aa/U1GAO@;)bR9aTD#
L1@)e(X(L>RA8EKW[IFT[)fg.L)4+S9KeD?KP_BeD-OZ\)]_93DPY6YZPH8e,10_
.RK:.I:DK[,b@DE[A:VYY3LC_(\#eY9EMc(PPW?gI9Y^252P#:YN#a@be23YLGUS
IH33Ag4gNG(T-W2-\5:16DZc15Z>_W^Z?7JS8KC;#94K_+<.^IHUe_]C-3-A3<FT
ZXcR-aAU<<+,dASWDQA=P11=Yc-67T^3?UZN>QEE<YCEC.V=;AYF81]+F8(M/0-+
c[+TeMA-LcDK4MFU&BZ3JbP-MgU9Ea0]8:V)3;1J4^XO^0+#6af@^=U[Y0dgU83)
.:D3(3KgYRT&M<DU/Y-YRVUBcJfAFY2ZIM4IB^]N4g,_>9G?.#CA+I/>-+>WdV-F
WDXSF>07aa=LPYd:YC^Sg5#2QI&5SJS5d0YS)gI,I.&-BP+=R2]POfYCHQ4/H2<N
=4YKcRKT3ME1AL4+BT(a=CHUE[+4H0WJ]6[M^d;g\GD+3;7@[,-cF[DU&WY=gTaL
>?1+U<.35?^S>FV3>NU5O;().YeR428YL;R]bUM]4W,>=?cK-4#cHQV-WQ8BGdUf
b?6b>EbW,;/K@PFW(\Q,4S.eIB/XfW0cZgM</,O/KCXeY;[SM.74I>]TOfLL&[ea
^9]<C[W&.GAT,Gg>N_M<<,^0/8.9>OP&c)0:K2B#F_^BW3;.U9Q.\IJe#d.+4EZ]
]1-6-7[0>&X=#:)KIPMBC]C8]E==;497cY)U[S^M,EaS6T?9RB;O^BbdMB<ZV<NJ
\-4B)]61596X5SN5IQ9^5,I;/be^\F4UEQ2Zb4-E/<Y8OB]d<^#L9-F(7L8&#L>F
/ST)e=558&/..PdR&<\Ce?@b<5@O5A#>36L1C[A\,PKc>a+SC880^/GB+2.X18W=
CUd5;K-Lb(1A]cYGGV6/#FD2GM.>;26QD]-8K)U15@I,FGUACaQ>4/DS9X0]b0/?
=-NbW)2O)FLDYfV7bQE4)NS5@E_(PL2^0[9NNYA=DEXRW7<e=#FU3=RDM@F/cOaC
7J4a&0&J>K:2f\gUH]b_<#Z5[](@C\6?+,NU,JbIGMY5,c?4a3K):])Q54(.Q=5T
Ze+^R[OBGN;,c?K/@,dH>[0..bb>W\J?LEVgd5//:TY7I?<#DH._/b4),b\<DRCJ
&87+-f#gX5AfP9]:eFTC8.J/(R(>J_BQa+KNb-J2fIee\?AO52&QB\7Yg;;VA??b
DS,0,C69-//fU3FJ5N8+/bECREW+65:#QR>9_<cb+-YY&9Q<2bJ52\U](Y&?+YK_
CT\).&5+(#UPf5HE,:.:Ic9KCO9_7\B&^K[8.NE=V=R165;40MdRE0-bHPDFIc#_
OaO/+YeDaR-G_HQd#Jf49H)32;/C73Qf;5Ae1c(VBGM/#QH_L3Wf^AJ2(+NVG209
g:F2JP)Q=K0e^\F_D>Z/VfC\2ZfUJ;)fMT;M_J^.@&0a<.Ca/#9gEcDBCdYRYJY)
SYCMeB3K/B\;PL2DF]J2\gQL_b,D#\F3E:e&_S<aC=6MHFN+JS^W9\7F667RFaaK
QD-3dPa#O2QPGVgMaXTG1@;W;MGcX.bb@/O(_g]7Q#ZC7_S3e:EWWaY,<(9Y;4g=
bee^>2^44];?LR5Wd#HYF)UO427D.G:C)Db&=S7QMJ94:d;4T?<+\0<]NGT8;-H]
H^FB2(GN\3RS+=bcbGU6K7I_;E,fUQ-;McAZU9&R[;<Q=X8\YX+;QNW5e<eHGJ_W
&H<44@AFX5:YPBLcb/U=_]\)LDML<WSFAeF#J?Y6)>-4aV?EcL[\/E4]#DU.5MBF
eTSO2L2eQZ+6NLR#G=]_X0Se)L^0KGT4C/42#_N9FP&QDA.-FV\9SOLOM^?RP31W
)H7Q5R>Mb^PcHf+dGF^P<Z5>TU8=Z:-a8C0.IaT[O>F0XKC-C4K-ecKHG6(W,-Ng
Rf[UWG:7QAB[@5;aUF7V>gN[f:R(4-FcBGF?Y-):a8WV_d@>Mf@6UN=4QfPa<Tg/
3+F@c_N<2_@7d3@(NR@0;5fBN>K,<T#\_QD8M96eZ]L&6O>SX&3R/@.H:RcdA0Id
09[=\dNBPg[0,I__VGOVg7IR9eR,GAQ^G(#ZYAJ@42X-CY@g3\a^T.4QU:c\W4P=
VMK3Q/8/DC5SbL:.gPE7LM,DaA=]DQ3)J>\N4M_S/aLcY-W,c@CWVO#Uc)=5c&W.
)g9FTPMbD7<gC8C+VK^e@@\]QLIJ9^a-42-/\5^MM&G_AD,=<;)c@8<B_>2RJ+e<
H]9\S,&RWQ,[MfM]IFH-I?CV4gWV=H[1fS6/W8^;VbOTTV?;#X37/,TXAD1H7e1?
-#?Y2?LU&e(G_X+QN=T66WDSLSBD@Q?5T^E/+AQG]1ML7f_2T(IE=>LP3L^NC__^
Af8U[a)]TDcg0RNRZ[+I?IgW.>G2Y7XRa#e]5+39#HEU8;EbU^_aRC@9WA1ScD..
Q=4>DTd>C4M;Qc:GE_&2D=@N([I,Z2O,8U2,f]Zc,4:eCPaFceB5+=0.35?g@&2d
R9c2K3f2PDNgB)8HNAS0YLYQ[edEZTHVX26]/Yc\E7^&,:RSYecR@=\6Y/@3B14D
](1Mb\?B)]cQ_/D:7VA;EFM[Ad;LD:9gH/U0<=SQ&K5g.?NK_I@#cMBV8K=1cXDE
<U]S<Q0Qf#MbKd?g42+3_E;7WB]e<+O1?f@M>d&CO4V#SARf@^6:2T+Yf@bI]KgN
;Y7L95-@_c@d=][8^T-MF;S\1+H#RC&7<VHO4#N>YbGX2@0T)?A];IH^,5/?YS4)
DC<>-3RbK^M::D1;_;2?B]N52UYH7)\dWP24bb<7MfgV^8^/gM=:KWQ:+C./.PM\
..,R([/LO_Sa>_+>BOU+gfB#W,(=[#B/_e:2@_TbTNb^6eGH3C((1&@_BH.,WZLf
I3a[5A.,#B\3FC@6BbM/2@;-ZRX&I#d\:OQ]8#1Hb0^]SIcMA?=af#]3,#]K(YJC
(X[?@MDRM)Je]N+Ff(3(S&fR0ANX)-7bWU4&5<<g6GVGP4.Va97MVZfN-7IP][bV
<Y6aD-9;95(YA1g]53bG3M4+)Cc^=&636FKYdBe,HYLO=5:eU7?]7U8aNb3UHW>F
X]91FZ76@YKb0COF/4=@A[#](2A1&a8U,VG8b5aG+HgSALC0.f49AJbF_.U5ZZ20
BaPda]X^<6YBG=VJG[X/@b?JBI^_@b^\Z+VBgS6[XJ;2T-X-9G?cSH^?:a<,-#9B
1]X:7YKZSff^@(bdEA5:H/02NH?(3T6&)R@CI+?d7N<_-QV?I]D1,WT;#3:XCe&:
;N5FO>H1S^[;YSe9\bXDAOKIJ8B0:9AUIHA/Q>N8/77]QTD?&gf=-dP\F-A6J7gS
Q.aOS^2f0D@@H/O&QN>O8D/egY<f1Y7V\GJ?O@OW4#5C,?@[WB-68-;Uge_5_IIJ
TQRJJ&4KTc?35AMA6^b+M@YF<D8MP(g4EJC]d[4VISDbJg25EY6O2YV8509.7?O?
,Z1<27XL&OaN6cU;7EL/B-31/J&OJ()_VY[XVFE^JIZP2B-.Q(PU10)6&)+1?L(;
9TG-7[6_3-4O,[.-=cW<I@90&/1WN)bcWJ-#9J&JA.RI3V<>TG2+dJ30cGc=4P5V
(<66ZQV#/>R/Da=@36OO5V:06a\A&ISZ+FP:WUDf^;2N#1,gZ++?^<G/CEXPLf([
O@^/GKVX/eA,6H&dQfL3/>RW_^E;a[@_O1b;E:1]IL_dQVQ.#b#BZB,ZVK-2[=02
1[K:Yc(&#@5=SFQ50T/E6/c@C<(=V@P-;FGZg[:6_RUC;G+F&C?X(<[_)OVN_<,\
(e(HB@[:ed<81V^2Q9V4744AcYAO]/OZKS2R5,7J+68aWD?LW,X;T9g(Z/3<J795
._6VHPe[bcGV->CC-K85@;(]4VH\b<Rf[)4].N&(4/>>aI9P3(UI]+LJU?9V-(/g
FRK+X]cfARG]Xg[62C;632QF;7Z-3=1,e+=F3QgS:Gb[=B((bP2L\D[E-X?c3W9&
ePBd[3/ab0J8:=+TZ.RdH>eLXH:&,U#c(#AQ0>OP(O0B<(>E(+=Oe&1OP<a=:APd
&\bBW_YX-Af6<K74cBAV[8IJfWS/WU.SQ6(RMH8:T=C4aPCV51_^;A+>J72O,1F3
]JSfU=S.Yd)W?:0?H3YS28MdBQ(?KO,N#a1]eL3.4BIbT&QYE2D<_;>GY]WX>EMU
e#:</;2\/,.CT\9<KLaDSXFc&c<[gPR?V-Y0>5J.)DK0^]+N(b<GQ3LT;Zd-KBG]
X6EDbQ8NK-];J5CJBOW#_V1-MA@G2bJYH8V=4_1MOBdGMHCZ-(UY3B)fa,IB0=?Y
BP:d==g_)WX,Y:U5gcRIJIb\[IaL1H;,V&_O&7a\)W(b5G1I,,<=Qc+1591,dF<[
#S0:/EUR0R:TY\^MfB8LU]RPK22aDUAX.8H\=?X_Lf676Y0=.=0RN3\[Q]QC2B?7
)R&@eO)C#E5VLAMS]\/8FeYE<??E6KH^B\:>5_UcYEg6/C?YZW<d-YdHH))NBNZF
#Mec=9+Y(_AFYVLG+_Zc+gfWNLN0^NN5fE5CCQ)@&..5U6;^&UVa-51>-EX??<(^
NP4->]_,&g(<PJ:H\-6\)(BXDP+H9K;LL;,UV#[-MY081[5Qg]gPcU3/cgX7UDG#
A-KT2YRXKF;,S@AU:W7MC?;Q3]8B@Q4)d(\F].Y7/?IXb\],M?PVQHZANVSW()51
ZY^&^043L43E79[aR<?>eb/4a,<=_ZNKdQ^e[^4C7IUg]ADW4XJD3V1BIPf2eI)g
YT/X604:+V#eYKLU/IWA3[6<M7f[6T+(+I;=QL;4e]bWJT:?C9c)54;6dc.X7DHO
bL,Mc]3f4E;f,B)Mg6?E>KT)1U#g4H.=bGT?KE0AHRM._-KdZ&/HTJdPaO;:7PfN
/-&:T07D+W@R.#@VX0SCC2e/ZMNYHW#2D@-0AM^Yc(T,Ha/8<YdKb:Ic.5R4G_@;
,N_[I?1OfL@^NHO?6V9\FB,+dF,P3XRIG;/4=AT8c>A-Y42YCCMOe-VH5#^B#a(&
4O:1./K&@Hf^:](-(J;9AZV;/\9,(](ZBCORPea&V9FRNO]7A0a=#[OfI>?S;5XE
Z9?CM).>eLI+PA3/ES)PZ0f1-[RRFfUa^UA>2F,U9Mf9@C+;e(?[T]+L?9P,46[c
^HTDXFFQ[b6GM>[69Ea>a(WKKHA@,.6Pdg@4RD,16QSH=VP/@f+DGD,35/_;KR=M
c]=F[U01BU:=P8,V7;9\=7@>H>(6,QEd,QPO_2Y(^9F4M61\S(W<VEPaO-Q;;Wb2
YXSQ1MMO6Qa&MUW)Q35-2I)[@#:A3&1XX+4+)3JaXU)&b=cT3\bYNVF;Y\YBSMc,
5;QE&WAJ-WUb1-Z=]=T)M3S_4F?4_/-HYZ9,0>WS>/W<Oce^d1TSP?)RSGV5_>\0
49/T1J\VUCe1>B:>Pc1c<8N?:QVLa+/):[9P9dUN=8RW\(g8V5dR]E(--:J[-U9+
H]UZXddbAJ=O&CQgNJgMT=edgegE1]T2<=^;8#84df9&.)BAUX_aSQJTe?[,;_W-
8^I(0(SIOb>UEf[+X?XNQ3Qg;7BDFHcf]TJe;2>>A^70/9D#6Y&T6N;6_Ig>G#8/
9aAe:[2_;dS>CIWW;^fRf1>E3CE?&K-&a1Wf1N4d)A+4E7HaJ^)SCDK,aIHP^Ke)
+.?3\9+>>aP6UEPPKBG7>M8:R_#+7TW)>H((AbU\Db>U-.VZR,+U.\R3cY/#Xd\&
<PWI2Kg#AZB&7.\I5N4TU59TF]ES6^0_L-d7I?I&MW4?\c/(;-911U?6VG/HC?.4
VfRZ3\:7cO.g],;&0gZc+M>Ne5JGcfKU2aS>>CPJ2/#S4;O#JgTVa.H<34R^7F;?
JQQZ-+/HVGbR(&:eEbD0#7f)3/8__aOP<+^VV]&W/2C5^6@7E^VTM]#.N\/?[?]O
JRFe.gRK8<?J@8)Q\VIIO5dF@+bSdA;bIN+SM\)H@[0#cOMM/_:N=HPCE6#cT9N7
Ob2ec&6]G._N)<+XU2_\LPWV+,FgMLO5c:_:2a<)dO>)7O2)cg@:U2:NPAGYK8/N
[:)L+[)aF4TJ9Pd+S.fVZI)PLGA4P[M\@,B]S>]d2G4WOY/A^aXcE,-0&XMffO7b
CD<03&:YXaF-KBaV1=[A-:96MLJC:;S4+4eO:C.K2B&9+^#L[KQ_)G=6JF3aNI6e
a4A3C(0\=W9I51:gfID:bMc&9,GU#?_YICU9M(J=8SQeZfK8B2A^P_b9O^7-95T/
/.61>W2/14Wbe5(V@.U&\UNRK50MC5LL6JCH=76W=41G1<fd70@)GIN-23AA7S.M
@OJX:g::U+/CEA4:7O\9N+.@:YMY._-9?)M470c#TSbGA3JHU5)b><6geHf.7J6G
6/VWgfC9ZMLX:J#;A?^9:Q>/B)<.88&KT[FMM-G\PgM+KX0A-aY?GXMTO)4<cY=6
4L]Z-\#dF+<fQgEWX6(45[7U4\#SE..(XfcWf;,-XU,.VC?5.0.WNH+W.B<:<Ndg
SJ(4gUJ)]S;bTKGV<dA7=:9USJGM^2eefD599ZVN,W.b\EZZ@JXd.Lf8,F7,B5-O
E6Z)G@]-9O=(c\W,2@fP;.84WOb@gb@>&.]gcO7c->BQfQ+X)BZV])LdL4<.8(^<
MDEf7MTY3-_AS@F=51cRAM.[2[JXK-MUC_IdZC)VB(a2/)\LXFU,489]3R?.TJ9>
c=X-:UTXXe5b?^-F2Eb(?BfGNYWY>Rb+Rg[f8.+&f/-Q.e#R0,UL6-5K^FB;8XSg
R-Od4IN^aUWSK6N7E8RKOP:4,1/[8eR60gK>@YG^F=:?-DObXJ-GC[MO#F]fPEII
&&DgBLg-0\a4)><YO,:-1HDJ8&KWU=BMO)LYgW0J71JCbgNTTB6caA[gV8caHMd7
#AP5:@3]2A?MPd?W.Sca#GcA[a<CA[g.>>CeC5O9TGF5aVUaN3JKY]T#NRLM9[Xf
/0<H.XN,&]/dWMR_D4V(2QH;,5]8.3^)-Mg8XCY@MaPG8^YM_[=/]+LC#FD6J[.[
,9K-0Q[#A41MG4AMc<,NddXGYB,A4JX>@[_0(eBK5-E[Y0c[+(c#Q2P2GX94O#M[
NXT5Y\IH1dUC<a2O?S=A\#S-<5]&+L/g>4#EUL1f._3=0U<PN^FPDWaP[6+3a]?_
DIA(fc:6#>d2bQX\OcZLHU=X,a,H+/T:GP&S9gQf)7\>H]6f@J&RUMJG1EE#5UWb
7:5:92(KNXB,^3NX64)(De83V_J4D9381I^SgJ;;Z1W.K\XY6S3AgSCCS_:4Y]>+
Q^OWJX9::;TCO#SPd2XFQ]WZ[6c@=>#?YKC_O#;XeDLT:3:@K(?T03?\9B[RUeYa
^Pg:N,bS_JcUSFc+b^eWdK@G7J26HE64cS\:+[1(eULNFK]#/&H@@>XO6HY88.1E
+;D7egSZ86T?UdZ_RWe.WP81Md)b+M2NacG4EW)V]X#S31NZae@b28L&+3W=<@.<
b:4d\VFETFb<\g/e\&6HJEf6#Cc&fSI>0=(.^S1=O8)LA]?JBdgW],I[@16KA34E
>Y210+1IOK1OC--5A-)21Xb?a\IDOX40?0/L=[,BOHD1;U=/\XDJ^X@e:/?YJXKM
[)]?+\30Ef(U3@J5<=c&D;>:8JPf02dI?=WA,4@GJ6=SJS7eOK[cZ\8BD.KAJbKF
Rb_W63[T2^0:HDdZ^S+WBCO-FP7Peg<R33bAb03fWP-KVSS61QMX:XC2RR?DfSF<
TM&FODfC;P\.-[06dZf4+/8SB:Ae,R:dE_LUI32a]dMe:bX_UCZSJYDK-3W1M5<U
QZYV>KGTc^,\cAT^Ee5:KJS?4;;>NdDfY0:S7U,fGU=\aeD\f5Y\PE:Q1F+74VdN
If_P.]2S/DcScY-d.2R.J+7SYE,IASRfXH4+GHR2-@]Q0COWgH)\:L]8(74.W[JU
U@;7cY=BgMR/1QHO(?aOPF9C?Xa=\H,a+92G040STFT1B.G/P=19@]UD2+K8(f5;
S^a1Z)a)CdD()/D0#I(a3;aT]IZZDbE^75KR)\6DX19,g1F7=aRH++M:W/_U9/T2
Fg+R:51I(N)R_4]>^&g]/eU[]EZeBC:4&^I?D2NSD#-G-f;1?9]ICUYBX]FNB8;W
(?9&_9MC_Ye,a]MLJLcHSE1&G0H2ad/5(b5/eQYG<XDZ#f8)=O(aeT-+^;gRIaO;
J-C#\[Ng/ad=@:\b,[_5e?\TD?G.Cc^NFT[B8@GDUHb^2bFa1A=f#5@B6Baa>S1-
(6)H,;S_1WKd2VRU&V81DE@92BE_]NPD];OS/(MOHRBA81J/fVN>cW-N>#X\#&NM
?1JP?>E@]?1+@c7O^OE-K:QG(;-Va6GOOQ?cea)dJ_2cU@-H+;c#,/9606O/T4AE
3<E2750:Pe(WV<OB40(QB>QB\VfUM]=EK5ZOa2NL7X7O^GL80Tc&J:+^F#ba@e:N
C_[,HX1bD^N.=dZ>U65=1ZV&@7/,;Y\FKV[_@Q71I0-8=S^XH28YR.H,bBO,](-R
D8/J?dF&ZLF^0=C&IeeZ?(J7K)[a-#N.Wg6^/Ve52AdV4\acaQ_,WB&D2KDMFK]S
HVOFH(aE_gGLFPVEOZEPB>dc\H[Bd&K=c<F6)?W=\NOF[2WLNdQ1:JCV>Q0X)Ecd
M?4A5KMCL[,ZXA>N@Z/OVRD338.>AE->#+186?9gMC_V5GU?8?H;)HV(I<FN_XIT
&MIBOabR@Ob^IBN(IV@W)N^5g_Q5FRbAeK8V6GRddg^WRW)#+[VfCOEOHAQEfG)V
gC(U](F^IR3>31>]1EEBC0/Z9R[I.XTX[61<FY0TQW3JeBSeVWaLFSK?Jdf4CBRY
8>QQ@0Y0&U5-b:)7_#]1UYR=6KQ[J1VH/XMM6dBI45SATbcg4:^2cAbX^#AK;/UG
INN5WeIL0+bR,5&39?J@edf=M_TL#0T()VUZJ+&=N>G=2C+F:g^\FS?RRd<?59&_
Rd&388Pgab#99E.\9GE9d]8Fgd1328AAXF2^>FPL(8V>SAeOIf?.gSXa99gK.UJc
C,Ba.5[_VNPSMP>]Q@.Y_-TMP9A#9AYNTSD0#V;W\KE&AL7JM1U#^U.+WP<L6fI7
WXL@R;>aUCMa7CfSD#D+0,;NBBT#E^S);E[+L<d##3cXZZa,8D)eKYHCM5J,fde-
agZ2X=\9WQdeZ:(S;,SDM;BK>/fZ#f1].:[AbW7T@OL&+/1<@N,XJOT&IDV8g;2H
UWDdI5-Q^XXW^[UX,A/-dZZ=HB@G6_(0<1/\9c1dCYSR2GO:I&^BTQ?W9N>EAM+f
5U<5b5EMP0U&Gd?M.BP1QAJM##P:R98>TBIC9T(88VVg/Q]O2C-\P@fFMc/L1B^[
X#68HeS0E0_R&5:B?(a0Z\M:E2HK@L,D_IXK,e8>-6BMGC]Nd4>aM-[R9H2L.>Z<
RGaag_#N4/=<1J1SR0e7eCH7M]M6-35>9fEI0fW@:Rc#TN>Zg<FV,[-<QD;fVW^E
,6Ac9RCQX.B\CM,&>eg^.XV)<1OW??2[.)L:5-M2,C;aC7bIOW:>;D3J4A-7H&(d
CKT3,eIBQ9/(UF)P-,5K_We236?N^)B+5K(<R7:R(VEO.F_U>)B^V#+7C2@g6g_P
e\9Jd9,GSAaBK?9<45#bYJG>A#V)[UR<8:S&V+38PQ<]6Lb#/[2V[ZaAA?+/)?N\
MVB1d@:#/d_P^U8/[JcgZ>P+:]J=#62N\WV6:Mb^4:TNTVEGDAF(QI)WYEZPJ1c@
_92U.403>WE\])CRAGDJJ8IF1^,b&<OBQRUa(Z/,A5>BcOOAQ+#C<)P<CPCeG11=
AaCW-9SQGGb1f_\#357K4X#;+MbV@_4b]]W22dR6X6L64/O;++FA+B[J_S&2+S,U
_?>:^Z7J(F))P1cK48)GT?faE#0Y+?OZb;@JM8>R1>;C_fG6B/P&J1gZ0FObSWef
(/&KTE7HWCXaX\B(1;?]HP,QZ[<>X+X4VZ/OOE2fT4_T@F>/,c_KU_\R1U9WHC7g
_F8DZd<NM8QgA?Z\_H]UJS,^F_2D0B#faHXUK.6V=O[LZZQ(KDJWP([;Ub+@fE9\
(]4J7QM.CB-,B,YeI.60[@:LLRK0BR4R]ag[f_5SI4CD(O+_+f&M@4&6V=CdOf#U
8F6UC1+RB^Yb_-U5J@F:?,C7OQ3Zf(#7SgdKZJ#KX<UI#3aV0Y<[[gS,Of4Q0]fb
eVASTMKZF5bg?5U;.)KX]Zb.bgWA[;J[Sae0_eaA2IW7]A+@bA;2aa@C>Z/aBN#g
44=,DLWFH_0Q#A6W84P[MBW6dPOAI,V+?afEbEI>VddMEcVNDDOgJARL6.<_\&1,
dLeSDIU4a-9FbSZ2c]W^IX)OFQ/)1X_4d37:\VWOK[OOZP@&,:EN+I&GR8\C8)15
W+,D1O(HPW+CK87BY1L&(Q@f8\2;4[:N=)#6R<:XX4\TBB.O+,^b>3#?T\C_ZT<J
efIU:L;IB[]L@9[>3aLaS&E9?XTEd;V5LSWO-GDY)<YAM1NH?&_;50/0573P7135
gIg,M51].)bAIcO9NI-QaZ5\.9=c.Qg>_A^#YS16Ub,7OIFL,5_68bd9e_@aIg_f
S>6TJ132+[5N&-,=?8WN8L[H=>;E]:2233[Fe^3/bQ+C;HZ=U:X).@FeXUXHX8Rc
B9aD,EB-<7/SSJ)A425PA+Fe)G9JXP1;UXA.-gaYIY)aU?PX,\GJ1>=X16a]P>RJ
HRHD&48-,T,FV?WL=1I(0.?b8-9)-)EdP\7/8((ULSDSX8..\JW(gM.QG\&&+6,]
5>1f@eQcR9./HELTY_17Z(SKR\^RKG=+707cK=/]+L)ED0::)H()69FRK0/gP^17
@6[@-)H+6:\//$
`endprotected


//vcs_lic_vip_protect
  `protected
WQV6fHI5P+[V6<=N)_^BfX<^W(>J8P+B7=S5W?N_]OfK7B[/7D.K&(;J/41?XMbS
a6EeN-SR&TW)3G&eONWI+VZd-8Y)HTYJ=(;5-JWf7Q)<CE,^S]=O2YJ?<B1RN&ZY
@Tg<Za3JM\TB20f#0;2_?T<cb#d?8+G-E=G4>AcH0/.a;S<2D]?,C6beE8[WF36+
TPG6@;Z81=-DBF(Y,[[H/f.U?VPF]fYKXS<U0#L/0G=ZIG?@I@ad3+[OUL][[H[Y
fY:.M&\.1eWK?YR8Z(gZ3)9MS2dQFN(+1B[P+MH))OAZ22E,@L[[Ic7B:QVNY#P_
?B&(;UOO_(aJ\CcE+RSg01GcZRBBYJC(g7YYRWH6f6M]FdSADZ#H,]AI.+30MCV^
VK\0&J<.B#0RI?F,^Y8OZ>XF3e(\4+-fJ;\+3A_NB4d^F1@g_XE;,5@T+,&I/aEN
5K4bRMH4GUd,C^.P.64TQY]9#XTDVda:_]-@Ze[2S1(7E(#S,.\ce7C_Bd.@VP3Z
T,N_D3C(d9HY>6.bf1#a\OX+f>Z/MCDXU.Y-J)\5MWV@CRZ]\cV&,-?JNE;S:H^W
#G,D5<)gD?c1^SDQZ0&CXI32ICWIA+\_^1YL.?TIK0\=>:AI,R>D-Dc,gFF,KB[Q
UFRH;Z;)d0^J]\Pa[?S,V)/U79WE2<1Rc59;6S?5H0&UM:574V5->1ACfHL&UZ2G
ZJ[]c]I?6YMfRXd]_Ke?+00^EWJY\[RZD=>S@JE?Q<J.=.a;L@<-RL@g<T@H8gX0
f=Q7G70/1[Y=D58LG_a&C<d^fY?DN)Zb/Ke5Ia>]SG);>:8,9:FJ=PZH@ag(0d+;
c1OJaF.=3b+-OY_/BKYdWd3K<WD.1/Lc+96F<S9XW.J[MVZgOeYP77.gcLR:?3,a
=LfKZHG;F.&>a(X_FZ(=ELGNA;;9@M+G(RN4<F5_O5UQdXI-(?-VbMBEL]6M\<]R
E8Q)aZ44X6Q@)Ze;0eT6739[S<MBd&\4FdE(.a(E#dD]7[)?)S0gR+NF3CG)#eMP
a27[=aPNT#Z4eZPEBAcNE-ZeP&^2SMC)SEK9_GcU>/A+-L[+0b&.E4L-@b;@1d^8
d3XK&3498:F7c=Y(F#5BX;d=/,1GcP-ARWeH?716BX0cCUSEK<HL^08)?5NSa+A(
LD_Z=;BaOAYJf[;KQBW.fe+Y9O9(<\ZP;ST2[81VYCO-/f007DOfNC\(.8XH)R3G
OFb[+J;-GY889R-5^:NT&PaKX@18[9X]D9(V(PN98IP:GFKZ3[=LMc-R[)UX\6R:
AU>I_R,=S/SPY2I+C^.c;5a]#VU=@Vge][2HWQWc>YAcWN]g-fOeG-f509017ZGb
cS.&bZ-8\TFcNWR\Pb_2;g&9?J5I,?@RDZR:/Ic1/d&2cSg+cd5UD0Je(9:(0M)H
MFTCQZK;+]bc+K>6=_g8ENR_?UKZ1XBK8BV.BVAIN,b4]\+_./\[OM2_:R_>=XbP
b0c=UGN6(f74A#5C2/+80[[^=\4(@&KM<PA]/N;T<\+EFMf60OXa_ZTcURPF2W94
]F#[1B04aDSbZ]5[:\Fd70@W_HX+7U#M@VK+OK?(.6H#;SS2Q2NT29d,#)D=CTHT
>CE<cT;=f?,))A@F,?WWJ^A71AL&?K+)DgMbg>DMaU1U\A@V?e,4G+V5^VYT7G82
f[C;[9aT=Q9RAaT,b8[=g?I7CMKNQIg=(2GMB16G?PKF^R]A9+BV?#8[4.YD5#9H
Gb4EBd8E#F&N7SK3U21Q1VEf,L<aLSKGEL.S4OX[C#g04\bgRR0=70273[E5ILUM
eVJLSO[O?.dE=1@Z>L-.UU:+V4Ef:)2]5;H1]g&3SI)b#YDB=<adE5fO?=aK?OK6
G_fYaIT?=[<7.B=LfaVeaI&g[S[eec5?c8f^C7)K.C&#U?;S]U<e\[_5)I^@#@B1
4A3[A[-36[.^gYQ.6FS:f3))W4bV9H20(OZ1c?]ScX<ALK?R=X-X<YfHC<RI0CSW
=aQ1a+]B&XAGgdK9JV]1VTF:aMbc3:.7S?]eHU)LA5>JTJE:0;P-HUZ;]W.,gRRE
46?<6YQI^bca,Q5.GX@;\1LT;LPH^1AMFSG7Sg0_#).EAJQ@LB^O:^7([^a(X5Td
e77)SG2ScM<,6YXD9[C3[00B((Z)eW@<Q?X.5eSX,T#EA$
`endprotected

`protected
;1Y@dCA8=<^W_L4<XD\+&6@e^e8dc1^7<S&@[&O9aT:(_fEIc]AH()cT+\?FS^L]
8_@CC,(ZJRL59.Q[&==:):C95.6dCWJ0W>.\MCPbT:faUYRdFf]54Q\:E8GU,I@7
J+I5@cLG/)LEPd\P0@7OU+((]\:NLU<Z)M(Z:TJ)7fMZJ16g>7@CY\0(E>P<SC8-
8S:?F^[=JY0aYFa\L<##d3XCW4]7Z^G+;$
`endprotected
                  
//vcs_lic_vip_protect
  `protected
#1PTS&,_R8Ge+??L#O+N=YYM6CIc?b)^TN\60,RY@aBTKP@#30?9.(JO^B1RH(aC
RR?O.5>&^EFD5#>2@[g<F,Vf4cG6C#O)T:]3HC^T,Cg9AXZ)Q4I^OBeZ<7@PMT>[
&Q#2M8#2M3[RAI@:Y45,[aIGB&FL7BJL_N>,0/gYaTWOG8<O\H=\FAUVGD=6&S+2
]5EKIb--6M2XKLc-H361I+F+5-8TI)N<)5VA1?>PRI<E,\]B^,Xd6([eIPcLR:.8
8g_ZfO.c#YKYXE=JGHKY]7]8fb-+=Sa[R@C7]L])a=Ie/UgPN5b;7K0c:5FD)1@f
8=MW5B;6?X)4bdZ3fF:Vf-KHR&;QIK0gMdR4VX7g)EL@fbB\RY@E@3DMHS3&W>.a
8E@[YLGZV1a-D2AP(&IUDL,P.UOET+>>Z9_5a;H3_cED-[JI2K[HO2GV5?NGTF[>
A3.018aCT0.=3773;T(>D2[AY^PN2Z(D]HXOc/Td3Z.QSX1;J6IV2/U:#48N_/9<
^[UT9.P[K=RB]M<ARE/4Z<=f<A&O6:_Z\LY7fcg_G>d6EUUHS>^/GNMG829/M1c9
,IbU06V@(eKQWf@MH90YL2N8?U;c,@R2(9RFFC?.a^W3G.?JL=C-a#Y#g#R;U=Se
\.gRU@Z)37;382&(^]/fBIT4cXA[XgY,aZ;&3M)3B2]FUIT<3CE]cMA9Z73X?P:K
_\Ag0-X3W).R,(aKA]F1,]^c77VWF<,eO=1900J2bI14S1&5fPO_&653SSW>a#W\
2G,6]#b/)U[><+:Q3BQ[ggOA+aRXZ3/<\c(F]SGESKcI:#C)U?G=T+FXgY[PW+/W
(C=?8f<INI<HN:7I8cM_3)S,39B:>CWO3a.dOgJJPS=<:-3KM>JOTDJ/U3::XF<7
S7A@8g3[@Y,CCKGZY)XV]S=;@ND2;-&8T20..Z:4L/Q)QKVaB7I4YN+ZOY=S=1--
8]OGGY=:YZ5)D_0#bH..+QE,bLV->IX-;E?,,^Uc3,\[O88QT&\a#&QH\SHL,Eb6
J)@K>Lg4/CdT#_gO8PYZ=@gFUX:>CU;,88HXBXgCaUc\@f3>_)^FGV[]N]-Bg4AR
>UGBZYH3,0CP6()UcKH_?:G(WHZ-<[+-G7+CDO_W=dL/5d<M[Q4(?b<+0a0<+3\9
UUOYDG&3(YE.83H5.NF=JZS<\JOO0[MUYY2Vcgb)6,YE\I-9N6@=UOJ82OLbfL<]
^Bd(210R+:gQeAA#FC1E\IA_Sg]R>+N>&Z08Y8JG8WP6@,aNKO69VM\fQ,9d=:X>
RS:^_:>R2@Z<6g5EP>LZ<A9/+J^ab(3QIK.:#+_f34=e_B0H1VUXUDTNCOBg^>G2
d/J+:=7.I11ESM69(NW1@2:6L3bLI/FD7(FWKfN@S\0&K;<-Z[S_gBUXPK^b[(5T
WTI;TG,]3SQI+)HOcYfH#(TZdI1G[A4f+=#ge5/?M2NR?<@f]gT#/^^g=&V-a2_V
_>B5P7Q4a,CETC9Q/(dJ&8?>84)-X9X4g9Bd5W<:;e=a&/e#XBd<CR:9F41NKa#f
:5fTZ[O45HS4G.(A(I,5I,><I\]#fAgN^P4F57^-#a[(<fG[YO8L;5[;O47:-47N
XYY,),R>F=<H)eGX&SCB0<7[YHG>QHL(:H2?8g)(B(<K>^;T):fbVLS[;ANRN2YM
6&?TZ)>BH,AED)^]0)AaK+_RBX/)Z[[V-&EWd+FS)6-4P&VEL1+\7UW:/^dPAEdE
BDFgME#b^B5bW1;X=PUZ@TV@(EWaP7ILg1[X>.a.B7[(OJA/F.M[G7.&\7DVR>\_
A;O#c^=HL-XHNGb@N?7UTECNG;X5,c0d5HARY]g171YgJXNTLWQf:@fA^,QA)T2+
6aM-]:W&X1TZ/5/;D7:-g+D9;d7LFQ@5=d6M3?d,V&9B-)KKc6CWTLN3:QU8/WR;
4V@9&)&E0ge>,0?3#M4YOUNc3-A;;SAHSC]Y,XYTJ[4F:a-GC_HG:eL[T#K/U59A
_YIeSc[W^B=Z0;aZe[4L&a420ae-S?P6AbO7Y#49CN4MPHE:5Ge)7D?&NE>Y5-^]
[K3ELSLCJTI91,U0L2[f.b)Hgg0:+)27ZcCSN21KV#[5BgR.NAgH[M=9]4VWdG24
;9CN-#SEQVC/ZU<J,54decGBGf:ORJf.^R4>Q27b@d_^bC4Q?R,D1ETVS/@WEAI6
YJXE3fUYfB(]:]E)<Ac<;2.QZF;c_7E(48H#T)0cC95_;ba7aQ.T-4<J5Ug\9(HE
DZ.(.>VJW37^_Y[2&[\Qbce7bcK_V5VBLIU4<VYMA]da-X[R2HH1).aMB^-gDRU;
MN<.]=gM<&;b-TU^T00H24@>\4(;8Hg@QRP8AaT\e1I[^AS)NaTf^73-PZ<T=Y>&
4./IW&&bDH:^R#76#ZXA)He\?_5(eQ/4IJ;.f5ALCFdaC^,+?5.F_dMZ)[1B\_.E
@;-SGR8V)QaMV-IB2G6c17KEC\B-ET>1@5LV>c&g#Ve^cGJLJN:\f0:5@SI49=9Y
6)=gbc5:R\@.eg6+RF(d7\]+XR+-TU,T)=\\O>6A_^2bF0A;bgAPg8VJ&fQ\BRPO
D;:,GEf^A\>Pc&CgGA#:NdE=_2U0)ERfH<BT6_O^00#I2Z-#=fM>@@_\--J#+<QM
+W4SFDW6[8C-aM<PaH)>=_&DWS[e?KZUHfB.LSS7N-@&R[-:_UU.M0.U-MHX[8g7
\GZO\TCYg-aG_@-Za_4g4;/JR&U&g[;V1/fW^=(T]g/2@;^MA82[0IV10\4KC2>P
G]K=He;^dNOA8X.0@;XM4:2-Y,DQ+29;.3=?N;>?Q589XYf_[[2A=I=cU=C4,LKJ
bTO5,+Y1=Y8=TdTF\8D.0d7gBG8M&[:&ISATaf\8&9;QIZ7O1;Y2Y=8R/dCbGKd5
BV3;MVdY#]?IROI#cW@^T]HUVMNU-3Q76NPc<ZJ:c/19ddb#S#\V>Bb:6BO/g]af
5/,/2<NgdCN(])Lg-R5FIC;6J#YU>(<4Y-fC4QM,K#;PD&c0\fIWX\;/8YQ&8S3?
I2S3#[T6\_LHB)?R?MK1-T>(KRAB;3WAJ8Y^,0<[[fccYIbHWYL,RA-BD#Z(FJ3a
\X>eEO.=/HgR0C4@.0E93]2NM[C65[I7I&Z&--@3M.cfJ>\E_d^\_YWWIXc4(5=Q
_@\JdGE7FBV=A(>#7Y_I5]e=K6I9)Bc5(E<c_Qb,T64Y27ZgC(W.HB4;VaC\:[g,
_VK=[@X(Z(Q(^&33-Y<=K57<W=>3QVL0T[#a7,Jg/b8XS).3gcG=)/^&f/]YE\V#
:@fg4DYW>AZFDbae8PESeeDD3+]KM=0E+EY@CfOY\);=^NcgK0U=L)(>[AS.;K6T
9GZMIFI+/]2g/N<C,<#fO<P<SJASe<f9]:c<3X^&Og[RSdT&34[D01FU9f[YCG_b
GaJ(0,5_])8+.9_+FBTS\^:Y#<Q@dMWT^)J0DR#\#]2+JDDCI-9MMUY<H)JfYESU
3,N^-J.E+a&4+X[+AUFTQ>bTKY8\0O(dQ:0e.AdaV?8T7Qe[RHN/#\-1)M\8,B)Z
T.S]Kc^MM.L.=HcL,B<ZEd-5]1TFDY4eQH,P;3/04a8PGTYJ.43I39ZH3K7Z+6TC
6MQa00J;e@]97,d_\()4>Tc5630WGb]b_dT02CbZ/f^PP]Dg<B.0&_1bZK0V^P0D
^.EIQ7_@;1FMbKa>5bAIF>-].I8MI#<d],NNf+M9X58#YXW7-)_=K.RRY,W4>I;;
S=,:-.M&0PW:0_&_a?\8gU&EUH:XO=(B10&G:PSW[VEN<;4bRSf5]1g^HF&ICf+6
ID520F;^IS_eH_dR5&cZ)b>Z-e;2+0.GdGe<]HT#5c@<cd03-\G&\K5U<<M6^IIF
XX,<Q#K[7U2^5+:AS:/><T-.EG=^\9&]H;KF+>8^8d>N[gCLB.>0Q.U>BYC20S=5
&6DDSE(OVJJ:;<SPY\\32&]D#:[L[I5U.+,#<VH9Ef@S1,VJQe66MNVHE29MU_\I
6,:4O02#<??P6@:=P><#RAOZ;5LAZ79T655-&,VTH4VfT&R:>cX5E41?99KHKVdL
cF7UO[;^1L@3)=-G,,B.F6g[42C6NT8F8^)+HUbVHT#_97@[a-bEDFG>,.&_b@X/
_#DUJ;.A,e_:QPG7.Z04K=U8:_7NUa-UHgaR,W?JL6C1g(B,_YM]&YT6]V5>ZfO4
S0=&R&e]O&3[a-,Ha[b]Y4E_NF3LbG^?-VF<O\VKF4^N>+AIL:):bR4=/Z>d[Bf[
Wf5;E1J1B85ObY&CI]7&G<EC0NI9=#f>)MF;&@KJ).JJ718_)\UW=?Lc2>F9P>eg
?4W0:]A+MCd^1\U;TOL?/L3=XC;QJdX8b7e)/1RSBSP+3;Z;]^[d]O</Y.#S?0YE
<FD\GPMTN.Z]W@XC>g@9V]]6;=:(??(,\U-7YV\MJY>7)I_Ta-aDc59]K8[d&H#>
(4N;K<?dDd;4D</X;T\NJ^aQ?>W\Qg?-W-PbN0+P<a>>dMCAH1?;P0B1:4UJgcJ-
^@62IBDe;U[/eaHK6+@IDd(AVC_QPg9NC:P^8Y\@SWW__XEFC@ED#1gEB/A^T?\F
2,_;/+)c^eTf(\:QPSGbY6L,)b4=:9@Z^#R3](?\J>5edDIb@Cc<O1YE^IZ81/aX
A<3N6JJ=RPC&0g,F[XRVe2@89Y^7CR1aZfM8:COQOg]=[U#0VO#13L7)H3N],7eE
R-<L/MLH)cIWG7.&KKG?F@P=g-/@dLA>;Z)9g)(<GRfRV6@;<@d()]>]GYOK;b?L
2;7e&T9I+Gd[S_Xa2D<?E[:A?[4f#eDJ=6g4D/(62YAKCFe&8L\Kg/.Y2V6eN1\C
/eYWgDH.c_[QEF#3AA9A8e_<[:#cN4#M(DAWe+9P_3D7JQ3g9IX#T#d?W]f3#fG]
(59eY\;<?,KM&=ZZH>(/5,cW,8]=a9(.[_)#;/=45D(F.-Zc^-7f;0e3f&bUO5#J
6f)1^1#^04VcF=GV.G0WP]84d;R&Y/d;IO2g73_AT.=-T9Lcd^0:Zd9_479&F<f7
]e-7>4-d7&\<a/5MMf1W,YJ[&DbB85K0TNPDGW>:-NJ]V]Ja.b2bGe4/R6@(a@/V
N(QBM3f2_Yg5]<3F&M+V;_LXHWA+I75M95YG_SQXLYYPD?3RCM1=[KJRQVPN=U@a
&e_f6/,_TM,,AR\.KJeT@WW?AAXWU3>KRNAFC,]#SMCP0RE^NBB\dMC-.6>-b/0R
gUAg5M9V?d[>RFIED^6@9U5LfOZ\Y@_..)e><\5JD7T.cTAB\M93>JHA5gQeVZ\<
<W=:d,0X)4][PNQ373>c(D+@?JPCfDLF_NT40:@O\OQQ]L:<aW6@D5T0.RdHAaK&
MV,M_5_bJ.X50E]R9Rb_]G]C=Je(;N^E#T7:7KK1QM@L&_R)TNFSQE^5;#Q]A#)T
1CK7PF;LT#FN?bNLUW/\SOW.,FDe(0@f\^EV#L1>BRXbNCY:9E^&cD.X?,Z6bC+W
IKT8c1NK:aN&P8a#6P&&ZbdW15/=2Qd78@2PONZaTYAB)GI&HJX3aa)OG0O12PUg
(M4XXQT-F/BP(ZBJd-RQ^LMTJA5F6H2?cGJ#5690WUfD9+)S9H4[EUJ.)AS,4/Z(
DTG])QA1eUIP9ID@6W-F.NAPK/@FRdd(CQd#]dV<&KaR7I79MR=PK\^.6K9-TV9E
dKQFc=__/<,YU:B_Ab[&DKa&Z1BQ@fMB4TQPgZC=F=I_6.VTb[-+@ROJ8&_@f3,L
/5g/<d.)H2LDK]L.J>6(3e_P1<Z574Qa-K)AO+&&G;-:?D57BDVF20I<+C=dT,>c
P?gb0;U&/fdEJOG-O1>&(DI#@UD3,QfQJ<<aagZ]I0UR_:0Q)+>2R]SCFVBDf(]?
1SU(:J9;<K/P7;5++I:KOLNUT-[OZ]Vb=M3]41AQHBAK7<UCXL(6Q.&RIOO-DKL3
#2bDDOLT^0d,dZW=cN4.E5>JbN626L.7P\&Y_6,^A<:@5ddY?CdS\,-2V,[0(]HT
bY0<GT4^?a7=/&UTCGA^8OVW;9J.P&5:HF\BdGgXJB16BIZ,;_=V\L(Od6Y:b0L4
BM]c88c;,+]<LSPVdM7Gc2.H.G<9Nc(=X&W@OX(1&LFQCcQ:2JEWRINM2=;PJRWH
DL/G)H6RULRCTP&,f/:SY_ZTYTWNRN]SU=WR7-aI<bPC+1aD.Lb)^PX)8BdY]QBJ
]&5VZ7VBG&a0T5?_FCJX+bKPY=3[DJc#YMg808=Sb@B:D)3/WALO2\J(O(JUMNAV
Z6@X=;-+9GR2^YCIAb#<(b98g1@ZAHD8VB]G@AXfK,1K.C.I@,dM&ZB1OaS+J2\M
\/T=W5fTc0\I[e?UGb\Y:/BEa7=MHT0LV;<</Sc0+;8<.=&A-+2ZLb0eg\LdeGOW
4R-.feYXD5McN:gS>VXNFDc7L;[:RQN;E5Z=+&<KM#2.a[D<UYR/Q<5;+Zd+:>4c
#OG?;K_O&=:1.L6Rg++c[Q:e=]].0,^/BLS0I77G=Xa)&Aeb^WY?J8,\XC=&g1GO
]_Z\O21Kd?&_Mfg;OY=^=^\T)7aML.)HO,A?[:XF)+,UgS=P=A.HPAO@K?bB\g_b
L;1\H931W9ffWPCf^#UR6M7^8QQ@)3)UN<I/afeBAd.VG,6B14fPT\KC[A#KAI3;
(#=dg@O+9M@\g3)ECJXLa0PQ.EVUL>3Q7N<.R#52e:Xc-M@A\,@GVY+_^9I\>M>I
#A.3:MOO016UW+Bg?\A:I5OAa4PdcO:9@I0cS=QBe9U@W/N:4T/gWMN@6Y?(XM3;
1F8^++17?/;-d1&]P+3fTZD\#]]3XM8X(:d;N<b7@cA6.@N43.A4c^72Y0Hga5M1
X\;Eg5fP-=U05Z+5(AGKTOR7<5JR<6RJ)X@E5(<1cA0A5XfR>HXg8=)GWGPX<JXN
5,Y0YAY.YV0K?1K^#9[J,_]R=@I&@=H52I4S1L_9.DLAS915O]_^KIB7AD^Mg)F,
(E_PQe0K4MNHTSR]CRb4&0]93SML=A=b&S@@5bKW,;4Q1OH03(a?J5V^HPe)B7^H
9H&7#Y17NOKP;8B4[?ad;_]8\IJM)D_XRJDc,U7[-SUVgYQ=&-5<P)WR=HJ;be.,
)?=16ZIf8a8^],S,5Xc7&&W#B#TS<^DQ.+RcVQ6L402)I95eDf778:Q&UBe\VOM1
<R>7@QLYUH-OL:dP2H+()&eX8(GVFRa,AY_&]NZ)6?[P0H:;2N.fFUdgD?(CLeg0
?1^:PJBb:KLHSZ&BI]RBV8\7N02A0Hcg2Nc0E_>N79R&+1[GCTHde3-2+WKA.aZ?
c2Z2.TI##\,)0[&8;c-O_9,B4c>U-_-=,>P,#BD6Vf722AMU,T^B:BI3J>Hf<VL^
?FNb[9[V,3<T5K\_9(]+D2#MWWLBTN53?QdPEBEL@<Xf^-.5<DLFfNI?.g_?Te?&
ge<bZa4aUc>=#M=,L,Xd\\_G]KITc\O6DP./Z(./RBNdbMb_>L<4+e(>e0]+34YL
Cc:fCOe\O6W__M4_--1U:M8^f[Y/G+<DKD2HdPMFdAcIb?I^G8DD=\2NO/Z]e,L9
M>[9-T#/1aDOEBWa99^[<g)5e[\>,I3Obb5fa;&83b@8GU7NQ18)I[WR=d9GEgC:
XXUAT.FPAABMK^P+P?Cfc6UD=/eX\e5W@C7K06&c2A4fbbG>AK_YSSI1.Xg:2-4N
Pc,EIF+-X-gYHX654XF\YJ)#@a1UP&1N@_0CFTQ7OR&>P:dH^YA/RY+9^Of.Hgb_
LJUS3IUZUPe]e?bM53Q\8J-Q/-d+H@/164OZ.g1@c(5<PTG8<[3NK>B^M=WYC^a-
RgYS[g7LIL)NW]O2B3^b:#bD@=+aU)3VCKK5_PTZdMHXIBF<@I(A?Be5c(^b_^3A
@Y_a<;9Z4bJ:P\ZH^fM5D8eVeb#92.>PEPf@ag\NW<R2S9TZ1F\R49C&]WORN)UW
X+5R_QQ6<bXaU,G.]&#/[TFd=X4)WNSQ,-9=KO3T@\?95Y?3EJ6Z71+Q)L(]]^6)
ZZ?8aN@1.:F9+(+LDP_0ZYQCaV.9@BN0cD8\K-d2I5QZ;R&f1;JHJDA;\_O9HT[]
41UAcEZQ(W2YXER\]Tg[=R9fYQG/<CS]+EA8a+2><V+<Ha,8N,_eN5fQ6-]5:52g
=[F6cD_,gg)X?V-894gK[N>N63e+Bc>bf>SBb5ff^3GR2^QL>W+P38NSb\DOYf2E
Q/LR>_2)_S5S6<F)X\FV?:<ATNYYKf_=LO8C:05D;MLJI5_WDGMR=)2\B6_7-#U[
8ZN^:LM4\_:CTdc]]TEC7/,YO0^IQ_&([6c)YgJQ:.\D-\O_UR4PYagG-[XVV0N)
fF.bUOZNPaYLY(b]Y2C)G1bLJUD4LPGQL.B:J3ZT^eL8IA;WKM[-&M]TDG79A]b[
P&bb1dd7^X:U]/aC?(#QG@8WLXU5g&HXYdGI/<gb;>EC]FP5ML-<PS)J&DD>:Q_G
/I06cGEK:Ue,_7+>^V<)[M1AF<(=6&H@R&8I7G.abS8&&1M]/M]+e4^4CIC/2/0:
;=<4J^SIV&48fD,J078N\5FM3\MU0N+>XfLP;UM_CL_6+QKG?-F99TG)7MM@7>,1
Ua;>WT5WN9f\>9Z<<=E>(&T6=C_&4NB3CHc3H_3#FTALfSD/P#?[fg]FC-0g]I/;
X<Z8=WII,aU>7F_,f7:6Q<0[_gXGA4MBB#2(9?3KC/)U<MA_-V:9]Wc=;6SL6AH:
&&&/adB=K;71=]W-@eSO]cE2FPYZF5L^[6IN-;VO#=5E@G\0,(dEc&P3X9WUB.4I
_IWaEKO0[9ZFT-bN<26==F<?FGMO\9KKe=B[U=TN8?Mf<EeZeKg,[V08L+T(#.\^
^\@faB>T[dV8GU)L5)41BMNfAf>=AS,0NOH)[[G7(Me;V6eGc#7b<XKXP^43Oc)I
+NaCWd8#Y7S:#:0H_bMGPacIQ\5Cdae-/&3]Z]M448bN[0_K)T^9/[D=.P@&#^J;
T/aCR66=-4R2FbdLZTCg3KS\.Geb[>/0&125-,@fD0=G&aZ.CeW>H1Pe]43dVXM#
&T4P5DdP3<WQ-@P1#fW^J#A:;S,4fO\/?09I##<JMS1BTPdK24SeI@;X<);g=.dN
OgKLU?O68@,-PDT9VZ1gbTX.\=@CP5@6V62/T>J#.7959IZ,R)O@fU;CQceV#G;I
^<V7+BcNd@.+D[S#/_2BV3F8g1eOB;XbMP\dCf02K\KGRC?5adD0SHGLD4DVX?R?
@#I\.:4\ZHUBD]a?&(7AJ8L4Q?P;8>Y.#7<c?#;TO;9C9P1:J#,W46;U<K:\X]G2
@gG+D0aBeB13G_&,3>^T6=A.eR0JNeO^Z=,6Y5Ea[0YM(=DC>JKY1V\2GY>)A-2B
]X:e((;TX/GFR+:dR8[M/WcW6;Q<\e92Z(US/Y6,-\=-;;2B]Q]^@dL/\C&.7KK:
dLd&5\Y7#H05+fE#^8_66d@fa9N/OH3>f18S=?V@@8K\B+R&ME18Yd;;dBDR/)W-
9LH(g])7;\=c+0R#VI<Z9=46_J.34^1+cS#JMSZ2f0:X\2fgLC593\)(P&T&2F.e
E]H76(\8HeG)HC\fXT-4b@5&C_VSLa<JP7]11ZOfHH)\G&72_WfSY_Y#<&-JFBbS
f,W@UU/Udf?)49.TD6H/(JZ7fd75-?.1dU8.d9@Q3c+>S@MJ?00D\(])G19_UH>\
YRaPT]9Z2YE1PY4^b.J6(]Z0CT^-1[A(Q7=-B7D0A&;4HI;1ODQ.,:(3?Og\_a,#
gE+]0/B1ZIK80aWc8/2TV5+=E@B#B?6ScC6I0B2H./U\SMSVJ)=09g.)XF[KW].+
&DT#W(\aE2)O78C?08.)S]NFAT<I/DRJN@_U?V&d9-eY?FX\B/1D>S]B5S@,_Tf)
K<@cS=G5Le)NB>98VbLb76:BT4,.A5EHA0gZ;d;>/34H/cG&Uae67]ICI@<)A@(>
WKHT825.\+>IVc<RC1@HQJBP7STVJUR>EFR@BRT2eP3I;B5ATJB=2cSA./[_B#4\
fcHc<V;BV)BNLD.W_])NRST>c<P6G4H33]C^YJ0WaG(\X>4_U&AMPQT6-;F#E3AV
OZ;)dZM]NfV8:SC+#^.bL+4,bJCCP@G/&L[T,.)ZEMM(J_9:+:4f^A@UFFH_JZQ#
5JJ)O-WF5A<7IB>JPI_fC3=NQ^E=;5OTV&H;Z5bb2PIJ&@EQCV-#W[=]f(YR1];3
&W\6dA1XI4NJ7E-)#BB^YeG@_:H4T;JIQ.+>aA\];M09M&Q?6dWQ:Fd2)[S(1HaM
M4?)/aB=)DeNb6#^0[A1AF[DGfd:4O:b7^IY#@<&>b>MXe#6VM[SRMg+(L-?O@:A
eJ/::QMc(2\K&AJ]-RF]G=ZWM,4G-A)N4-[@afPGR<_9O3VF=f6cYB:e,01X>g=C
)3bE1-/2GTOeBWCF81P^3fWZc-UYMd=-,O&PcDNF7FY+)Q^\fAQ8BG7AaHR-)Nfc
_Cg6+]5;(d89=W3)FbbW@)R0_QALb_1]5)XOS8>[cZSNS,B:_F#d#=Df]a,=1^JC
/e\[,2g#Hf/Cg]2OBY6VD#-g^:)]^[W=-=8J#&If6e#cCP7@XEaUYITF49a<0+A#
HBKN2_]+++[KP+e8+RA]2<LL_J<N)1YDVT;]@=c17287:\5<>c]G8+;X<)\c655a
PXK>LC3-JfVeA6<4Z@O@@6.LH3Z_9X4OTI3g@^&S4XeR_Q1Wf>8T2YWK06_f]YHR
J):KD83;N]]+T<KQL8LCY5f;FRTXC=MfDIT/C5ZM9H0.F-#2>;^/6]\:.+N1aQZ(
PB6Q-AWe5Md3Y-M#_Z+VK3#P?7@>)bPPNG.b-<aGQBB4-,2eB4YbN)FdU5LEDa?7
Cg_Q6aY_1--9+TfN#AWWA1W^5K8\&<TYe@ZS0f@ML.J.eP0g0LLa&>@U3HJ_QKQ1
-Y>(Va13?.>#>EU=^^5:0U[#://V>/?35W.IL9)_&(2D,/^GT.8ZB:?P>?GQ4<,d
CZB:Y@L([^PG[2FP7GX6[@bJ=Lg8[CA_O#:6N:(+B\QIb6D&T_5TJY35P7,d,+@-
SR_b//[#W\a&2EeO/++&_99^6L5LA4HA71^.A:XgC.I+\Y@Ac9VQ>6\CA1HfI7WX
4T]Z>bEX@Z,W<dR#0??MEcgaES1PFYg>c@](Wag?E25PT(TE6b,f)=8BSADALFf,
?S+U[&6a.+XSWKED>P.efU#HD9fL_1IMX>\U<@aB;HBXYg7>f45)0HBC@TVP8@)5
g]?.]gb<XQg<^3#_3#CTaP82FW.^27@WH41PFAR79_59^AR(1:K96AS:Y,fTN_5/
C6:NWb8IKDN2dRM?]cHJZ>[K,W#R3__A7+KOA6H94[RKgbN0,<#:819]<4=UIdI<
,#H-=GJ(@6C+YH5>JI(ZAbT(QgcP]LH(S9cUcD<.P-8Y-V(JZC^P^N+^_<c&_(E>
WEF,V+LGe)3O?8cecZSQ5YZS-H6W/SKN\90\OGLYUT6U:VNNOINP,YgV_Ug+[SS^
QCM6=/Lg6fJS642)^N?Yc<YTT&E8Z+2N(0S)c:I#CA]MF73e-.SO,>G6Igga/#9R
PPI39WMT\[QeJE989BV&&8MKgDg;3VYP<>>_[PIT66E13cc>CS[2QH4J@Z6A+:3>
T5?S4H2P)5_\19O6gUCB)2TaCS10\PK)SeEdc_7K+DI&@(Ib\Oe4.f?eda6D.^KG
N,;_\J>IaK[L8:]XAJ@FEYg5/4LX9ZFEd[c7)BQH(C/2V<=/Z;=@OGL?-),I?5:D
&UcBC.e:YXXHJDY^037edN9g;V^?K,)2[)M3WE:DF?Z7#A7aQ4Ab-;CS4:ePCP?Z
S6THTea)=\5^O\==>M/N<IDdA@RCY>cXE]WI=[]&6@U9Q;+H9Z<8QD,[DV^.#U+W
J]6_eQ)EF8M_XQV9#B\U5Da<-+(C#KKU2DL#,FO54Z5FW=@,ZWa(2(9Y/:#;J#?2
2-EV0KM;d-Ra(Q?>4?;7g_dKV06Vb/eaTW?LAaHb(AO\>OX9DCGL9f+;ZNRRbb&(
E4N3[.d#=S4(fe2;62;R@I.\+Id]:,4:,#UN]<PC=P,=g8c71+#8=,bN]9^L6RZf
=#1X_A>)W0C.CQ5[d+4_aS@&e?>9bb;)RR,59(I:g_N/@:K_Q:F2TJU]6UTVB]G1
0eH>a9)7a</1f#5E0H(JTPF1:+2:7=?eU&=.L#G8P.X;]AfZ8W<F.bGO_3&CE=[=
KDO<HV)O3DYE4]6Xf+U1P#.10ASJ&29R+fK0b#GEM]Ad=1Y=dC]V_6XGd7=BH8]T
_#(+X^@TS[gaO@LH<DLa.3g.TJ<g;g7ZN5eOVPgG/b2XF\/)_.[\SbL>LScV7CZW
Jc,g]OeO&a6+NI;^_;89_;VH1?B_/UaD_fa#>gb10)HK=<QD&L3?343T#0Z1eLdC
-5NJ&E6U80.>:O0CQ;X\GbXd5;/S]<b5b>+fYG-40b9g=37/)LB[I\fd-gb2LTHd
f=D#]E?>L.&D^DdHH=S42_G6X@g9De+=;)@=M6JOW:V8;=T-+S3NdOFaPCX.-L2V
E4daf=/Q_M,dD46=SU=9(:AEU-2RNB^H230^&Qac(82geRTXHT65H(Y=PdSG7VFE
Jd5@7E#.NcG34YOJ1O42TLYZff6P&GMH.K#T(.b#cQA]^B1VM)8f^PCCDb?G)5\?
]E_0f:Sg7GL>EVV&g3GDC>eSD,Z#A4PAN7^Pc3e0A@5P)E1WPIP2Y)K(P6;K5d?L
M&RAJ-&;_S(d/-V/H]<:=K.[:SG0/]W>>Ff=H:5-T</B@7@D]GadQ(E,0^W><Mfd
da9Z66RFP1RJ0UT)-N<)L5fWW;+e]Wdae<<_TON76WQ:+2c3DRM;A<aW@<3RR^TF
cH9/XO6;\.U[79H[E&+57Mc4b1]eKB8#6a87?[eFW7T6?JD=LBad2G61f6Q1VL.C
A-Z(gH_8)fgGeTH21FU3,RfZDJQgH=[V877ER6]bF;8-KPd1Z3DJb(@330/I+=5Q
?(H.C^9#aX>>@#0fb>CGEHMGWZNN(9T<bGW0Ae;:J/e8Nc0V.OUI^Q=F@D/_-2;R
AUFYbF-)GUA2HRMaI-/=:05M3ffeU(1;T1eNTf@4(OM4BWE/];<.MX4K.)5.#,(=
>8&gOQ7cLMD@UaHI/CeRb-aJR1d-=QdI?V0E=C:O<.B1Kg[7HRNDOIf3DIZAQ-@B
S#[3cLa#D&@QS#4I=\A0XM1OfK;CJUbMU)9^0[I6>=PV81^dRO<+&EI3=b#]OH4B
AZ4T7P8^B:6Hd+8\5B_:>Ie]4Oc(FGb4.Ze2#7-]_c4;\=MNQR<BH-S(992;DfB=
&);CUG4.(=5V&YM4+Og<)=<8C;_\S6>@W9<KSIGW36Y.f62#Gg\Dc=@AEJ)Z(&]-
]#a@#_A_H&ZS^3_YUTK>K+Oe5SV4D:.P:@&QSgQC_:c0D0L[.-,_9M.4?Of&Q:6W
;1.\?R89^7S/XBC]O7Fb)1c^DHFV^0JEfA.?QR,Q4a[Q9LN9E?Y4JK1<U?9Q-L+C
=+(@>)PHM&IKfEQZU4C7]D[RHF7Ia:G7JG;A/DfZ(QC_EGL(UYGYQ=7+Eg,#NJY@
4Je:;9&8GI&IgB]&C[f4e4M95314CeLPQB.-,[YJU)R6JH5[PD=/7G=.9.S\XVS-
D@4;b#OL)WZKG3g<UU(PL#F>>W:?\6(fG1G@cNDgB,<).1BDM2#XDBX.cDRgL=J=
>8\E:(Df1-I.Z08K_b+Q9SEN55G;9_85G5#(c#PM\5J-;BS#<WL(;&_+He/L=7/c
M<Rb&R=JSc1B]5b-39;28[6<4W<D579-d1:K^Be,>C44H6A&@,3#K\C819HP#6PW
e?(RL6e_T#=F^1W8W3694cbGIV2F+OH&a7fKEWD6F/K>4(6HU;ZC^UE6cM?UJ#Ue
R[A)eCGCbU>D>#dZ6K8Z&N?)/NN(dY-c>-13@T&ANSHC+VbMR\b&370\KO?aGA&8
KIT?P10FCS4BE:@_XH,CbI]2gALZOYO6L5#K@JEf71L>?;/W8;/R)PDMJ9YX9C0^
>e_A[M7Y5E>?^?6S_RJ(/Be^.5O>6cJ#^&CeB2^(eN4]/-W0_4<#J^5<ITfJ_cA]
_,5[-0)eEe09cAcc,VHHL<IMQeKU82Z,Z(c4+60Tb7I[7B@\D6B8-[XDAgQ()f-d
:RD7,:V^-H8OSU4>YbbNVa/.]=()D)]?-<34ZD,-4^g5+Q&1[RFeQAD;S08\3ODX
0):fBfJ71^.KHU<a=/#2cCYM9=\).E>,cdRD8f8J(ZgP;g[PHBTYE;7d9gYZNZ&3
)>ZP97c&@6gc?f4d_Z6L\e)HdE-<dcG&C^:#S[A>QV9L/YDYL^CF2NTL393aOOB/
BG]5?f,c).Y2^cFSE+5a^WZ;^?DF;Fgd&bCgXcTE4?6DIL^+Nc2:?^:G276([d_X
<a@KGM+C-#=dcTHV]P@R9]/>A<>b3J,PV=+aZJF+c?:-<Jf=@7V0+=f..Ca)@X)b
da(bM&E=N&:)Z.5.aWR(4^gVJ_0<GeOb_LTXb^:[?f(WX_Q1gP2&C?VfI>^/#[.1
9_\Y]HYfG2V@XVXQ;[2>NBX12J&=&=AT#Hc@Da&DLGB85@)O02LFeH?DQU\-6D22
#W;5@b,eNFZR90=>c[B@/Y]?c&Jb1UC.b1]:CH)?XI/M4LNU)+f/_)&e2>dKFWRA
ZDeAGf5=9<cVd<I(cL+C)Yf>5^J<BX-]3(EFg7BaUT=JDZ<bE-?;V6[D:+_WT9BN
:6O0ed4T[MI3g.V4PR2I6]+ZIFC)DDI&aOde-V)/[WD^KP+\Z>>2#A[A8@a#8cbX
SVM7AWa^JaP7=@V)EdgO3U7bfeO)f2?_cQZPOaE@4J/g2S=VfeZGHOY<DX;A3JY6
D(W43^FB1e3GS<,gb#62eNZ/&Ng=?QYKVeT)9WbMaG:CML:G_Z&Z,N3T+)M_OL;M
H.e(J&G1PZJ?fd^8M/PW<&IFa/-0/UT+HNXg8=9ce+@@-;_D#BT>O?=728<c<R&2
g2a5PcAD@^ECgF()1fgSR2B(aH;fb743-UOU7,>-WQY&VILAYVHTURdL=:>ec/E-
^(J=H)^AE:[U90\bZ]801O/P)e02>FV=LfRGE?f-cbVC?DP4/F^K2-DH:e2>;fMT
HU-fJ,L:+NURIAVDAPA,I:PS,@f^Z?H+L3gHV6g(^Ha&=<ON_.<NS_aV@Z6AY<1L
NT4G:Q3C#]@A+1bd(b7-U]WY1\A357/WeMA\Ed=a[N8f,bZJ;Y6fO\Ub1ODNH?=A
PgW;S5AO=K(+A4U6e2E#FeEKc&,11b.W-YcTCQZ+YcLK3E2+PPKJ/9:VWD2XL]Wg
M:-c0GJ442a6A-]AgMOSA8Z<a3_CI75cNe1;F:DC<&DBD93F@f7O\0#HI6S3cIOc
/6^b]fG:eQ7UN(PCY(1A]&Y<dZD0XN4)GS(.8+N=b81_NW7:eG9CD:P82^C5b-,&
HCF9A9)Sg(g.QD83:W@WeeV]8e@=:b0(-NB&K]B7P?cDN.PBI#CUbdNMNB&L#H#W
DX2Ra^?FV;=M_1@<P(]_GQ&TQ/D;?WHfP\3G@_M+L5_7RZ6e4Ae(a3Z>+YD?NFZ:
CaF5aQ#5gQ/458K4Z7=:d^gd8QRCCUQ.IT1;3+SK-E?OBJQ;2\&6E65c&1B-/fNE
V,@DZcf,/[1;]=5_dd,AF,Za:2>&aCUGUgM@[.ObO+(ERgRF<GJGXP^RNT^b3Hf_
:e<+CONQ>)=3/S.a.1?P#ZD5>?DFZ)GM\B+;09N:P1[.V>(HD:BB3fXK+B+6SPHA
,JPP)B=M=:d/Hb=GEL=8D;ZB(VZgJX/7S,dMXLN==42X_4/]P4=aM7#MB41:#C)E
JOY?36bJfW1T^eFQD<R;ReaQeZM[7g;:P>++O[ZbT26-#-d@)TUa:X<B(TL^;KA+
Td6H49.FAM8g^.<SJ6A??[TC9IFE?,AJ?B\6I53AY\_\HI_4H,V;CA,GbMN[gE0a
PT=,O:Z5[P;9=>R)ff_+^EMSSUdE9B=&^FL#A<fLBG2,5WQ9T44++#2DR3&FJ3gR
>Ce7_)^RIH11DM1gM+.GV-N:OHbR<Z)V0d3JE_3QTZ?\<bc>IWTZ;:=10=B6.Fec
/>c@H5EA#QgH4A]bQ#]X=2eYRT1bG.J5GD4K>=T-ET\CDdKN3#_CHNY8<G/I4M7W
d_QJK4238+6B@8@>4aML+S:ZW9(8PU1Lf?WG7X&KK/\;UdeC&c&&16\T-P.<P7<Z
J=f0YLT80CZ]&62)1Ta3^4CR#I\,^;JQ>XJg1E3KaW:T:^]3=QLKX>Z5?PENTfe\
Wgf7M698<c42FVfMW2XR,8OcY8UFPZ8+;K)-G3VLV.CJV/NKHT4G@Z[QX6e:&Q(-
G]BOLL;?2a:&6U]44\WYO.9a2M=6[]:\\LH,V+I+BEcM/3d0DB@LSH.e/2,.-HXZ
)5<<GA741Ac\(8UbA=+Y#/gFU\dI@f-Xb@e3H.dYOf37&),4IT;8gefb^,VEYbT_
bN;&JL35bXZ::BTcH(gR/e_V.G5U[EBdF=KdF:JN/.YWOV_4D@G(1#,Gf5T[#@R2
)5G]&\9RCdMZ]OV>e8+M1ICLc>PW=,HX5B&g#L4.N<d?0KZQ52N2YbPe0b#aY=-\
F2Bf6c:--=M:FJ&FP6SBELg76EG]7;/[.DM;&4fK4(4(R>-QQS=\=Hd>@,IZ-1cH
KRWWb4\=U&4bD/3fGU?B,S5RW.g-03O1>R7A1)Y_F;d>Y(28KPHZAN@^3Ad00<Y3
Z.51D-O/@(OX6acdH]I&0F/_-F+SKA)-?0B_39>U)<]AIXE_@+5f1+V^>Q[e<X[R
J?XTSN8ed&_+@+VP.e)+dd9AbdcDFIc0CG&^g#C/P)Ic\ab.&>TJdILZVF9_\/9E
HcefF;]3ORfB]^.gg9a.H0Z4V2;M45ZeL1W9,\(NgL^:Bb-;;d,C2FC8#/O)>Lb2
VFP8B][gZ=\54-A-W-L=YL5W3[4=+GB,0dDAB/Z(2+DP_0RH60V)C,b@1,D<:RLK
A+=(HPUG-:P2S6,LaERU1;0H>PP90)H0.fZBZ_#JRSeWQ-D72@T.@JB3d)TDR#aW
LO/4T1?HR>Q^[ECg.<1AA71SY(N9I6VeDI0D/TNR0YbG1N?BF?(SS.1eQUSW5UX>
\L@>R3gJFEMV/9[2+<D@@a=d3+R[=T;59gZ0F7e&:+<2/#cbB=<TK9+=YNBS5XYP
XW@QdGa_PWBOeR&W(L[-AN#?-F&1e(4NF?bg<e-9(FYS+gH_e2ZQ(;-N9.8J#5F2
G;9P]ZU&d@N?SBY;20VBW;bSP>X68a&27OT_O:QC+5b))#Z_==W-2LJgD^,J,+eN
AT,V/GF^Ka]3[gRDJc2g&/()6IECI&&HaCZIA&@;CTALbRB4Z1C61H)..3YJNE7V
Ta>\F2(5IF)Z,T@Q=C040]Bac((b+K(f.:#>+f3YV]WbWg9dXf;[WgT&_@BWX)d;
S(BBKI3&Y.\>#6.0NU02LH<=c[8,DZb,)Ngc&XSQD8I4B]B);3d5WgGeH,(5e=T&
;4)>/XgJ1DG5UNW].[I.<.GC?0QH;AAHBJaHSgZ0Rd[Ja2B5L4cOHIc4)W@#SM&O
5d/G:/Ye++b>_-K-S2)CWAF[[7.B+<9\b0_(50(?_2@7NJ6f71=K7&>S+c(g.Yf]
,UXOd1RfgC>I7+)eG0f1L>AbD;Pb^EHb3BZ0+#-P#K=;=OEP(E:6Q(R#-J52a#a4
TUHFKGN=/-f6\e+MS2M?)&YG6)V/PUU..+THHDS^KG6(TU^(L1NPZ>GCc_AQd67I
6R(1&Q(_:;W)^=E,(96MdQK5PfN(\V3f)<FH,CF1(77_X-Ve[2#HY.42eK[gP6;&
:87C(4^35X+)#Y0E,J0Ef)SN#;R3S[Rf_IJ870Y_5-.M;5FL,7Q]J@TB)P?V#W6G
g]B;HJOHQ+\:BCNBK#6&)X@R<UQ07;JW6Xf4a=/R/VZ2\D>EEe<O?7R0g6YG@MSF
)#QFgDg\g&#gb6aF/SUJ7R:BRTZ91P_VQ?[73,b]ga+2W1Sd(2/489a[>J4I[LgX
89AFM=H]TTZ])^/OG?Kf<&,.>X=)WI2g=^>F[O0JU\2&?\FG7_NIfVZ7W5-Ya5#N
7=E.&-WNLMZ&gCMF0dUS,d<##C?>3aMK.J_NYVOGMH[KGMg6Z^bZZINXLN7X@=7G
gcUGe;M#AXK+d(Jcf6PGBDfC2AZd??7MPRXL.1Y0MR]KFa\bcI@;7_^_LA_ZV77C
<6NISE:\.:^#OMC^T8H206C]DZbf)RA#5[,T,Ia-S^Q#S^(=W:9YH5b6:<g?@]ZF
PQf3#::DaGGTS70R]cZESU71MNI-9+&F&]LTL60\/F98]AY_cZAR0NU:&2fbc:LA
P:7_GB0J19Lb6::=X5DcUI8d5g0@B(IEd&^:P8fd7URHPea9&OE&cU,:R47OdcC-
F5g?E0?)TKQM]T<c7./c(2e[Q<a6[dED_X)UE-B42;3(V]+WQ4UWQG].JL(/e1ge
[^6ZNRK\G[.:R:(&^9gZ>J/R?-R,BKAVb1L2bg@fP]A@>H13I8cZ#(b25QGMR;V0
P#d-HVVT9@NW@W1SP]-=;]2^:ME^KK-cJ,bPC^f33EI1Q&456,B#33BE:>D0R\G3
L<HT[YG)2^,92?2bM^@]Q40c<A<H7THO+M)FF3M2BDZYD0Y6R:WK/SOTM&9Q.c2A
[R35X9cf,S[+RV8Y>GAdeK,9^;5B#/BE;..OJV&U8GV]NY3_.OG/#+W^,D_@@/]S
,OWb^?/XC?Tc(ceHO3D#-Y(:BV&18K>[L?_4K^]3#AO0;S+b:KJWg58Ue^#YL28I
83^<T)4Af8dPOCDQc7TD8-XBe9[J/^<BY3]=.<gc30YOAL:M5VSR.W>\]VV7&1QC
UW?:NI.L4W/L&FY7)bG>HHG96QG,^\WK=cL,R+Jad)RF:[SME6.X,.;R94RgO#Ag
b71F<_M<MP,..OG)RO\__[<_M^,F.NH[@bED.<R^85g:M(?S@J?H872QVS=c6U[V
T6OJAPT@ZE]b]XOd4,T^AM2YHM:#8d.[YE5XegXQ=d\cYC;OgS2&(3Pc2c\&+@9>
/[,CdI,W6@-V.L&7JPAP?7gf<8[b760-P;2<Ud#UBVJY<8^=/.JL)=[.NKT7ZZ?0
JFbOe=LAU-VAR><(bCF)/+2R.\)1(;J@F7])fS5d#Laa4\]7eK0):^LUAe9VC12V
)#.^R,aL=)a,_4<](K;59a&c;==fCYVIc2ZQ4cBE5@0L/050^6E.;B46]&)T4).W
.W8g[GcJ?K\C?EV#O65@,F7IWA\7T<]S1cJP7_F0XEBfcS4#3.HDO&,\SYKB1eFP
92=Y_a-POB&D,G]^9U5=??FeF54Z8#W)74:[ae55FG35SdOHe:3@YJW>aA;Va[f8
S^@Q@[G3[^3)cQ-2&XcUY1]S4X7=[..WUUKZ&36[g,6ag7V/-XS+)X4Fb_bgdB(;
6e#.OH(ddW>KY^/13gZ6F1X:?e?;&^;3PC8Oe-@6.U=eKa-@?9HfUD?a&CdRcBc3
.EMg_VQ+\O92>f@:9S2R9#a>Qg>7-\^BeO@X.Ta6U652&):;++C1,DL^2a1@.=23
Y+PBOU0Q\5?0Y:FaP(F(1EFLHZ:dNPe90TPGf#gMJaYXW:>V=7-fTR]BNU+\>_6J
Hg2]#gI,ZAN\N:QW@-(SBZJ\Nb8OUOWN_I;J_<>ePDC_@gX>6YN(>O1Z7;2@ZTPM
6HDdcZMU/G8(7_g;g33-QL^6/4CJA<4J-W+LEACe;bF77N.<3d@LK5UJ.-cDW,K4
CV>Zg?_(f)0=W?,#N+U6d+b0CGD.L;5>_Z[bgG8H/1C\85Ac>e.F7..-45LYQ+TT
;&DFWDEeGg7VG++\A(A5XUQ?3K,-L<1d64EB+&[_1#;D]b-R2\d]4GO^#d7E(K7I
JLSIb6L5@I/?NBH/^5G-85RH6TQ7\>3+?=QOJeD6[Z?OQg009/U&aJW;&NB47c31
N0+?P:>8bZe,YR-_M?\>,/YMf?K818^PbJD&d+\D(6?eL0Zc<^CU-bDTg7@>>X5K
d+=XD&(9N]+D81_Z7N>:S8&A_0=4aKCS(#WTaV.Y.R/W>.-</A)NA^f8[#P[HSQX
+BTXL/Q76QD;Ag=\EF]J-eU_f3=ae[1N]Wg\-@.LRbFEMAU/K#Nf5?#&5KG=W56\
Mc.U0(=/Gb1LEbae7[<e/V^VU(103Ef;+>V^71(>aU)+H\+)Ve\S\1-N-;Z:_K^-
=WgQg2Ye)AC0)65#C9X?7LgL;KDag_YVbOYIaVdRe@;412DK3JF=0,KaE:d-TW1.
Q?PCU<HbO82)+G:)K=GAUc6;A:VgaP,@7e7IfH&R1EB23NRBP3G8N+(E&e#Fe@[G
A7>?.]TZ9#Q0RB?;1_6&3&<J>bGQe0<H.b8CeJM-X3(-[9cC2TF#=.3VSA1Y=P^:
O2aTKM_4^f<=;-(ZK(?=)POO&g\)J;Ce=&0;4gbVKE^&ZCVY33/\^g)J^-EO^4(B
c[4c:#A-TNbWGPc<MTB_;e=eQR4C4ab5D7.,bRIYNd-<LIYS+R6YLXT\Q&20@=MV
@Q.9_G5ARYZdZ8DP?cS[<adTJbZC>NSV5&,E3^X(QS3?4,UK8R-E&D&I>E<OQfG7
X5K:(X^X6OQYcLL<eB[f),]/c&aQ0Agg9CdCV9A[FH_UD>0LAef\#e&4:9HS7#6,
Y_/IJOd:D)(57Vb#S>UYg/gS+YX#,/?756.d2>Y;#SF)S@_gJD4Q:.=MSWF^2[&O
M_9MVP([GUUGJDF1S#\Y5[gYS\-)3FSDFQ-/Og7A.AJ7Gfa4TZ@[;(e>c+LK)+;J
/=LXX<OK]QO89Bdf.=#J&25W1)[[LZ5?S=[?MTC8[#287?344VB\?Vdc,XNYf[^P
(9KAZ)\//bZd.F+,ASE@<D:_N8Z6A&.Faf1:_XITW8959E<#IP1Cf+\#81,-HBZF
fVM3/XK5]DAScc#(WDd1K=NQf0&1/aXH4GYYO6;)cKd-^\U1W/d3]G2469.Db+Q5
d&#I6-75[?[VKVe9MIY.f[)Ec2_>D=f-)NbL^c#bcR1J0AEQHPD>a5IWKQ7DW<gA
M/.,,Y.8G,R70DEf0CaX&[LCL1ZQ.KUA</g7=DE/[EJMD.3c)Ha4EF;+Nf:a?X:G
JY-P>WFE6g;9d>aM=fK4gdHd=_2ZZ?;.1>XebK7c(O/&@:[g6JW<Zf__(W64M;W2
C?,Ie?_41.M#(K+\G]WY#??eW#EOEQ[fXFZHU.@?I7T:U@TX6gSJE]B;:&2>FGHf
Wa^[4RBN:Kb2ZU25LKH8f6@Ed9<D502)gK3,<IPI=FEgFI(Q]?eb2M[1590B=Z1E
\/FE&H(P>H0AMMZUI&)D5KcJe,-?FFNf_&BP33:FOH.;39[/NBfL;RP)[+232R&^
2caf>dD#6JG2JgA7FcTUFATJVB5IA@2KO./+?Cf7=OYPgPA.I()0e&U/-BIB)Z=B
]9;6#+FQQ8W:g?,aP>S3O/E.XOL5IP3(eb3)T[eU[5MOTA_<HPUSGWD-IUW07SBO
_ZF.XO0M#I/H<50TdDPB7&LRI[-/LA3Y4@2[0=+4cCBgP[<P_K6G_DVS+DOFcN:f
I/=G\I2J.R;SPO@X+61M26?[DN]BW)TadYHM?X^K[b6R]J\9B/=X^I::>)3>_.IJ
CcMEe:\4^]X#L.)LCIGZF+=3=4?6_4G(_Ze.^b)PQg.^8<QX50bY@I]F7).>a;bP
[Bf;Y3f._,Ia?P(EHWPd3EQIQOb[Q2Xc;N1.P84LJZAfaJV,<g6;.GC#R8,HSd]P
E0V<NccT+-Q>LICV5c)/+De8a?P#eI-1QH;Q>N+BC+_(F=Ec/3;<K7T2A;C5[7_\
(7d6L9PF@T<WZf2P=>U,16Ef\R?)I08ea?f&)c@XB](F((7_8M#E8B,U&W108A.1
8Y1(>GU]W/D7N^81@1;Za?V3g4_:4+VY(GB7aV_dB.dbNXeIDJH.F#8ODgSTC<TF
\)EK;d3KcD47Y?Dc)CT93,GA#JCMPAH[Y0WgIRM8/AV_Bf>O+b3#D16FVK+6DK9@
F1=4;2[0=g@._FbM24-aT(H4PAg]TQK[;W6T(FE5cQ/>fKI?13c-O>)fSS0D?-91
#22^c7=6:dMKP#IJ-&;5a^4RdVL]Y:f5Vd1df/VC_-UGa(Sb^H-.I,=&@119YIKS
;_aK;K\];W-JCBG659;EE+8XJEK34Z:[;g4V?Uc<ZO0Of(;9aJ=<e9X_).0[JTK5
LdL=G[?UHf&d_\OGX.3A3JSa0f9f,P-W5:AM)W)DaeW6N@639@.UX^2O>09GcTGf
=b^O;^UdNXd1X5OW.da:NZ^#;VLR#V0;O[7J12]b?IG+XD43)==a)28F)(_T#OOY
043DJcK4/<4R)DcG3[C<DQLbZNeK2F:J,/<BXcb9Q/(ACe81[=aXZc7W&:ZU[D@Z
?@?5Q#UDF?XY:1+@BS=__6;\?0=<[O\GZJ1UJEX^D1_Sc>;L1>21G7S\@<EO(cBf
OF>XS_/,8gGLb@Y-89Zf93M:&&fI([RV2=QeN3B6R5.eYfX612_Lc_/Q)Wa3W#g<
]KYe/JXO9MUM5Qc]Y#XMO;R#ZO72PCXPE>XMS^K93a&DB\2N0L,]LGVN0O5CC>LP
DC2a4CYg2Q0_V<,f[0bBP)5V@)J,[SV=;QK1SOB4&:;RLFM[Z@VNK8Zdd=_bc_.A
c&3+LX-bT8X?5FJ(.K[QFX,^=T.cD[WO^NI(cAT7>MSUYTgESMMD^.^e.faebUN-
X4K5:HDRM3^4C&K?Jg/Z.(2g);C[8C?:(.U_NgP7+TIe,AG;3MLJT(IXCZ5O)V7Q
S0.B<Z#M>(g]RGN_a,[75YR33IL^feB2Ic+CO])PW^(b8^^T=7IKPM@f8/ZA-f.H
D^NaBO:\UE9GV(MFK8@T_OFg54DLS6VH0IRZJ7?BH;BZ;?52Vc.^4?8DMT+;4[cQ
eAbSIZ#N#1K6NG,G/&ScZ4?=7f^W.JZZMgT1473;S#E-/RgN^U7PR^(K6ZA9.8^C
S+/H-9]Hb?DJf9[)GDQ2X1.bg5A#S:;+1OV+?)[-+ZWg&bJV(2gN]\;dW/bS_d@2
=[\#[E^b+[(OEfK8M1fK:e.IQJL;^@#;;(92Y5b]E;#H98H[BHI6baJc/S8-U;ea
<VX;;C_;.^/@,C\4BX>\g0EQ2MA]VJO3-@e[6(.gXRcEIX_GQHDb/:F?Sa#fMc>Y
A]78>^-6g0,#T9^/MWV.VU[#U4&?AXS:3E37SU9-F^]KGDBGVdd0#eK6AK=@05bF
GAC7c.TRR3)M1&=J8f,3eQ(E@H+[P:O<O+:G7?dZ]JM3-;.-+FH(TYVXH=8LbHed
:3gDWaL2d;JZ-]8.aTOH(FgQK:KeV@1+C_f.#.12R58:[&73gf1.06H4F-b_DUS1
Q\I[5R3/F/NQf)6.-9)KV7/2;g?O21N0.;VS;e4^GR.[M)>3:Ma[115;WAFBGe5K
CU7=#HYMCDP@ART31V\#5a,)Od<Z@/?)CV3+K.Y?,NQ_8-@2\&4.6,-K/DL0],c;
W]@()&6ab57:V[?=9IdB_(5g1MLQV&KS:dGU7-R@U<ZLGV5QK3_b(OEGa7ce7V[6
Z(:dM217-AY;PLCGdXaP-L_0(Q+H)(^4?]c,Lg4f^2TXEF+#FKbLF:7&10UfbWB?
]]a(C>2Nc:OHg4Y4MS&]S:(X+=2Od[FN=@ODbI\(eN]L>If6e&0Y>cV4:N,037cI
RI60)F588HSM_HB2&J35Z0_0I>9:UQJFVDOY?(K_BePJZRA9ADZ6G)NS,eHPG5U(
9@8C-9=CVZYcKW3G6bf)+F7DT_KP([AG9]Q5gJOOW5NGNaM0JD5b8C<K-=1NVKe-
53^NA_UL6\Hb-[V#W<dU4B&CE;[IV-RQ5^Df@44gaODS>VgJ[D84:(-&8K<I-Jf0
J:+?^#LSYXBBA(-S[[8+eQ\EI8Y.J=Hf/L>AMH/M>>&ROQHVaaP\X6>C6?AN01Y.
dTSH_1-_dKQFZZ3L+_406V7W@0U]U>LVFYT<1]?L5EfP=9RYdaOY//HE=Se843AA
0,8deDd/)K<+=N:C@fgF6,Tc\<;1<PYK+XdAB3ETEAS#6CLcOUR[M+g\SW?\a>5W
@9(M=-@12=CRL[X2RRR>A9=[4@cf)+QK.ZOQdP:(dLQgb[R,QbH7Z/AM/60B/]DL
d=\.B_OV[9]R\+&[<^I4:48P[F6@Q&H\[F4<69gIM+//LR)K#MBENG99>_F9.aX&
9;gDZ66PGU;F[Lf2ZY:09R^e)R)eHOFcK]GJ]D]76<_#V>GXR7M\Yg^5CU6M]TI@
\4f4QYXYU9UN_4d4g3OY0+)#>bKM2G#3XCb0e@BeMLaW0(47IAe>YT8OY>^(U.D;
D1Ya0eMZZ:e^4)6;MJ3K=UN+BbJLKLD&TT0=GU22.NeORTD_M9U=gL4,4_ac5TID
BB#/I2CWW\7D44HeNB_<Ed?L/LD3#V6[>DMO[?\/[FLZZ[.H.P1<<ND@)\8a&<X9
JK:Na6/CXX/VbS.c,MMcFO[fV_U4[^;OG@K@0Cebb8PQDR1==9Q9X7-<8=40Na)c
OUH(M/@^3E[R6E=X7[K(>O^^Gf^;UO9,G/7g.OA11QT3cCb#6bC&JDMCYEX[]ceU
&JVOJG;0b6D5AVa<FNRQWN?SM3d@>609NEUUH[B0RLOfVOg?#a9Aa9L7fI,R;Q/R
Y@Y;:YaDPK^_EC]#a.+@Kb]_.VH[IBCMeA#F3A3<?00Q_]+O]OZW\A[IPNe+d?8+
[eg\9]8R2W5A#&687G?Ma/:^(e[&7LV<RSH@_d)IPY/HaFTHZOU3D4SAc1=,J4Q#
>,dfW7IVdYFUX,Af.(+_aEJ3AI4b6A^_d;eC]H3U/g<dSMD\CIQVR/D/;4,5A2:<
g-Xa^:.<&F>eB))e6)fd74ZU1fY>ZEc:\-6(=aD_eW0[^+L3=?8bS8OQc^)\7cF0
.5[bPd4d=Ha4W)89Y1^=,:DJ<ISc1&_1dBADN5(>W;8=>/;RB#(RWL#91a.M(L,@
?=7L<VZ:dM,P95_4+7#G=;N&SJ];FXDgbaK&XZQL<;6<N/^>8FYS4KPC4\,@\^I9
.V=8<@I>Fb7#Q5.2=MB3::ML.?Zcg4X7RKe3>SXE6NX1[.T#RJ,4ZVX^QTOIXb3K
>[aWFCMZ4@)JbF^A6A-YH+RKe&H7@A[gWOd]@RTM7-3ZTd8I\2=1]I?7L)4[28E:
HM\7\X_G+b\b9(V4&L18R,AR3Y>VPZA(g<8:P^,-Q?I:)M#IYd;ON2>^-bT_SF>#
Rf9<eC#?27=d6:\Ka^CZZV3G5BH;gO5?C4@)_.0LU1>C>+F)FCPcX,Z]OWA2e_K)
,503>+I\/9M^UgGV@X;GHXL2V4KQ>#dAT,<ZY6T(=:LZJdYWQCM^VYZd]b;IJJ=#
5gCAZ1aKVH#W;e53.J0?[U1+#_C215E^f]>85eT(JA=eRS@M7]NKGbd>d^C>8@Od
DI;1L6+X=cdLV)9R#AXP_b)+_3<aPDF#?^b\e]U;U0&Ofab_I+EXILN2KXNMbWPS
1@?Y.Wd<:RQ@+WfeZ,51)JLf_O+@&16V8)O,AB2^Dg9MI90D,ASR5F_^T4d#E@Af
dMJ;)9P_WWS33MC[#&UP.6ggU96J-fK^2CgPYME6.\Z.AH:b,8VU]Q#_/-5UH3>:
=\)#LT8+2(aB8S]^;dQW-_/aSY:PO^\D8ZdI8]ScfG7];e&g;eIR2M8:daL)FPC^
+;8R4E?<GH,5?&GDCGf/^.2#N<^QNFN1B(5FQ5R@2,Cd2:8D6fB8D0CH_\VSXSS#
0M83,(E3c^G_.2RV&PZ.D[/2SI?(b@)VPf8C58Z_bag7?HgF:-DX:K9+1TJA+.8=
ODWXe.ZU)MNcbSU-82\X3L2c@8KfdQUa38UIB.A9]<(YA55?e>K34/#9XG1e5RdK
\JZ_OZ<<FcSgD]BfdAbcAd]S[WcO)?V2J&Z/IR>+VF7.;TB]<eB2#bQZIAFJ/@:V
)gQGfP4&XL?e3&Y7ZPU[e[d^Fb3VaPTRcJ,FD<K_+a\eVS^K5&,5;4-:+J.@25(M
GP65=^03M?)#SGUb=114QI2dXa]^BJM0FRR&+6+P=@GN:E=(LS-A5)b&-JgU^W&f
FAFK#QJT4#1/GP<dIfUZN2>RX.KEHZ8--]>4f-FK;_HMP<(NS=Cb/d@gT(0eN?<0
2gX@10Y+1];]N#2Q97ZTR<L<;1bT7&)AT;)3.WQ93P<H@;a#0.9D=G4[Z(CF<cfd
1+.P10(F<UPE-gG<@(-[+aBL_9OW[1WN&4=b9G&W](O).QgL^2?NNVA4g+FE/T/O
:?B_=<DE:0FX-W)4ZaPFY+HFD.X5C?IOL0^PZXW:/HGRce24a=-U;>-2g7L34&c^
(aR31X81PSH:NdVLF]YD(_a4[9Kd^.;Kgc@[L#/8OJ.F)J+Y+(X1O^DN;.7E2S_4
O-R?fR_QgHUYMRD(PBHL-8PZBLaQ8JgQ4c1J8gaAX<^7LT8-Z<7F4F1/dRZK4>.]
6\7O]e<.d,(X9ES?35[Q,R;M1L6\LD7?JN[(R1U=S(>9VD1E\7WR[F5JGb>N540G
5IQIb+BH5C(SNB#G;A:436RL[KIX\N(:U=MZOW:2Q7a3&_/1Qf(UXLV_NIYBL<&W
?9^6(XEYC&CNLC-]F;?J.V^LaK<N^X@PQ_#EEWW.L,Kc/7(HHY:01)8JGOLg\a[e
#STc&9?,+T.A,,MT>?[>EC177P>f;:SNd;d20L;1WV7U+WISgKO83].K:8,RKKZ.
LgA.#K7KeVPKBRE)+C9XE2Z6<#O;RD8T+].>V#>YNIG>4ANYdYQ^8@Da3UE4[03)
ETQ7^(XX4K<_F)X6X1@BBaT6P9Ae>@19Y;bIN6B@KHNTAI-IUB<R5.F0^W;?L0f-
3gI&/f]5c/K)dZ^\6T,e]X\].7\GT_::bGBVU]=Q3/PVaEO]@7>=.J(Y:=+MHYEF
fC5GMJLe6J/>Hg?#fR\+_>=.3(K<ZY3?0;CEMN>#caHZEfPSbWJ^-GL]]DPV#5=.
-N34JYO7G>M_-(C&@OMc0&=#GT;4L<,9:[@P;:=4E>c]VZ+MaKUPY0514CXff<(f
&c10\:3\G9\7f\[96]>8CSX/[>6>RG+TKL?fg9A=:O_a=15NNe7H6bSYa16Sdd@c
_Pgf7<4K^VD\0?/\2JN4.cdLbJ+UY6OJ)X1c]V-Q+2I1ce[+\#d1Y=ETD.Ag,:DE
,_0H.BP0bMJN]P02fBa@aTY=DK7:(Q;XG/W(WM_#VSAY=?ARJMZ,fUR,6Z)ZI6d]
M27[P>/Te=)JZ1_ML_ST2[O.7PURB<-/5N&T?B;HT2TIS=/?:K[K8dNVB2A5#O\\
FB0JRS00?R[_^<0aI5B]^PS1)CJE8^;J:d1e0/>82CIC:a#[L;XWa19&8bZ(&H^R
>6VA7T371X.VfA-AVUGGHcS.L5cQ^O8#VOGJ9V(-AeZ1:^A<3&a1#K^EgIUfS0/&
2.R4[(@6C@2M@>B:dPWB^K>7,fQHO;aT8.A+ZRFYRG8-PM[HEdMPYbIaL.CbMU4>
aM<L4O;L<JW&W1>L<K]HV/2Jb<a\)3/X;<[dQA_fP-X)4bfMSg:.\NfUab:G#[1g
1J9NUVg64WX+X0QM.P=g?+I@JX[P/->7B=2.LGbU]7cW0QQZV4(@#\R@LG&&R#bO
NW^]c]X;Q>-24(5NAD/U_d.72F]/KT_P/:8=[V3ea].0<BZZ/#:I2.V9U)92\&F\
&fBC&#V=PQOI1E.U?6(Gf-@6-:G9Ue2<:5:VSBXFD6.#Q?1<3UX]Og2_O[QJ=57[
)#HYU:M<]&7<7WPUM2Y3Ig_EWGdX[OE\4_;d;@#b)da\(DTWQB.M_^VKQ2C-GNbb
A0;_8Za@\GD=F=M:K2A4IOT4:G0=04&25Y>WSa:KM18\ES<(69;b_<=YYVAd>RBC
6^NX\6ZQ+XM<E4ENH8\a9aE@D;>T)Ub@TAKRT)T=S=3])C1=>0:JOGc?cCe@,/+#
E,IU@3cFd2NR)7AQT-<1#ZHBKNLRb;&D)S/.6WJDdX6QM04VB2&TUM<&P.\bG)VM
Z^9FG3-Z,I3-Q(d^:)+C_^7LS/d7Le:+K_AL36cgE8V1Qd5#-AB/9A=>PDHT9Z1T
N^b]6^J>g)/59]/JH?PE^.:7f:4]>_:E<WV\9^#@Q.F#7X]@>,d;\-14\6X9P=G.
:^J#-)9])\E<]5d(;9>-G;/2+O[/+=->Z<F_2OacdDW,SHHfFg-_S34<\gGDMPOF
5g?dBI5\I^C)d8/U_H[(/ZPHXM/B)f)(JP;K)_EW6G1f[EVC]_85>:5^8\2<7BS8
;5b4dUN5,1^_^@V^gTb]S4A>G3_>^XfSW33WT@?fMQT:bPd6014L@-e1<;9U.L_M
AP=b[K\NHM-?DZgC.1WDQ-TE+HQ-bRCGW9NIL]#3D?b,DFKYLYf:9Q6Bf[5)DaNO
D)]B;)^9:S9/K][S\b>&aHU58S(5I74>#>e@Q82W5:Rf7-5VK&9C]/Y2g=#R0H6^
g#E&E1ZbBT?D5ZM5I9ERg\P]I]/;d5;WH44@f74&->]Y1<TS\>GWOfD3FP.XDd\e
WXSH+]8&>8+I1DGKOE/CDV9<B0_-DUS;4f-Y2TZ,;N^^[\Q&O:2F/E]6WM/NR3P7
@]#MJb;\I]:gY40-P;R(>L&dWN_PS0fRM6&<LF/e,T]Ab\1HWWE]GgBOe_>6<-71
LXb^cd5(]0dJP6[1g>NDgB-_]H&:8Z1#6,0QDS;2.UN;@XZ>U:bL;L@F&5;/ZT<6
8=-)d(+E\YZ[5/beOBB[79G#f;fH_0e-PP,35g?NVV[[g>Kabdf?=B]f2b7BI:3>
D?J?3K2&/?2EcOHX#(_L<.F84I5WG6?4_G9F)b2Z+@BU4JFZf.Se>.:V>]\8g8U=
NH^\U(A-B=5FbLZ[Ld<MW[cNM^>VRFU09fc:14:E9,3@)HZEZ@dYN#YH70+.1M3P
Ge,,&YK?6W6VBN]cU^-cc4B=d]2_[KS=.eM00<8E?NR#&TQ7)3S5I=4_^Fb^:4-g
66(,;)<G;.^VBfPG3W1C@N=SN<RUJ).HRg:;T3BVLHC\Y5R^YK@VNMZ_U#3,K6Xd
6);/)L0MWT^dFegI>(=KaYX_<4O@@M.LZLRE9/I/<#[(-)DM_07+-Ef6X7fBP4d=
E+W6,O\.3/B)3Ze9I\5+g&IbbRKXXUg+,1(/ONU-NN2Od5E9aO;/-)DD#2IM,0fX
gKWR_4PfaIK4TeB<_Z(W&.CWVL=V]JcaA9+bVd\fHHJR/@.#OcS3@.EDJAPC&W2b
NgVJY7eF5-0C\VI\1O?A1&d1;3=Q+\ZSIS4:S]A/YaaL12\TGE]f9AB7RS_/_)=V
PBcEL-MT9@Ud:T?BcaDWf7XYXH1A?HQEL4e>;VML^g\PLYeTH+?QbA=BW,E>8?V\
1Ad3eJ^\9c?PQDe-4WWBM&bA)#FPJQHK?OAbf#K;1H:UDF.F\cBC[E(I545+6;T&
#-[:;JH@T0+9],5099e53UJ[eQc[^RP#;b3e/dagF&6QPdGL@&@K-6^T3&(WZdTS
e-?Kb\R/K17^=?@Ee&,Bd,L-e3),#GMU_\\:/^HF#,\]JReT./Dbg8:Z:+F>8J7e
M8&g0b.51,X/-EHNaMR@#9MM8//F#=bK[\5Q+&[;5]DZCT-e]Ub.\GV&2]_#=P6,
10-WH37VG:T>gRO<A=.;4N=]7Td0KB.R@WX+f(N>_IS>MHc?K.N]IaC1/0(L#PdO
_6RYV^EXJ/YI?]S8=.P3gCJ#OaWN(=/;#bF,I8gZCT_[FbF?e8(&2f^_718\.)eC
=Y2cJ#II02f\fZ]FPDR_7X&cAdcD#H1cb+27aaIH1?_IX&e,QHNMdbDW\.-8GM(4
09KCC[L-N^#(+3g-OS5F<X:+]=N>-G3&G^MLLMM4W9K._#YdZ-RYD:Qc51,O5BG6
])2#6]9/]7Z.e(AD88&=YfZfMP@\<=NeVET=b<5V.;P]X2e]9^UVPZHd[_cXRH:Q
#Bb.2:&bTgETU2:c]ZF._a).^W3^gCd^1\@,Q/3]L604IHfKK]TM2W5@H1DIDXK[
RV&XP87^8QW,&8YaaO?248GVV^ZHI,Vc_+#.FbI:.Q=.I:U[DeR^F2\,.?GUf^29
c^d@SNM_^1<-2IbX;G[+BC3B&YF4<H5X6,]=1O?.TL;3NeFAVO2dEL7<E5;b,J=+
cT,2Xg/?FY&\IY_:Od<FRI:,:N9QSD6PaE&[-3+:S).Q:M(;KV,OgfLY-RKJ)bF>
fgg0RLMNN<973a2SB4Ya6F+?2,K=AWA:Na@+UEcHH_X;NFV/eS?3KS4gOXeN+ePd
9PX@1AEF?UC,fb#KKY-PH.<=TU1FNQP2bH2P@+;Q6;2;=A<7^M4UKGb)Cb\#QAL\
ICYCbJ[;_0R0^QbFYgXe.]6529,&g61F8>-)A]fWJB:+-JL^gGO(/MMe;Z62]Ue&
SCWg)fDOE)2RD_(6gdKX1eRGQ>Dd5/6I9=)95g;<PD\;RfQ=A93^5[OHE>X8ZGT7
1_=\?abLJ#?0+QCFI7-9dJD:b5DaU4.3K\E9dZJ83)NKJD55e]c2<(J4#7PeD<d9
6W23>Y]cS)3(X\5(.b>6:Ng2);+O2DU8)O_J;5^Bf@X7\^DH&BDC/\TWd1SQ+VOP
,J,I8d57):eX-4Be7^YS:egCAM2-PYIbMYMW>(O/<_UNPWf5Q7G.F^;K9^HM#,-a
,IXWF(INCgNA1U)f=0L&,cHIbfUS-aV0QdK(fYFWG;J8SD_##U9K\d5ceR8OU;Tf
<fc(MQ\,:Ke:EU-@^QN\OT/G4;MgOTTT7SVJGF^AJc/5QNCIZG,=c0\;R?[\T#:_
R9dK\a3#8T._G#MP9M^2X?.Q,\aU.I1f)8d9Q05fYdD02?4VfB6;)P@gDD67[](R
@c^bg<;?U32Af0BI#XLKJE-S(:@g+_fJ++/30dFJ7I-ag<,2[SZ03QFQ.L3K@[2>
-9ASe)Xg(5,_0D+QgPC9XXf3WK<CAd\QWJ;?&(EaEJ)#4MIQeY.D=Qe\9/<aNIQg
1gOJ6LP1D=NcADDbG(E#75XNcR[P@<4Tf7KS6-K=/[B(W7UY+dIF_e>+R:JG(Z,T
.3F]YYLB)M.U=G[MALE0;1TbICSF^RMbH;/dG6V;V/eYP)F@Z)D@I#]G#_/FfKa>
2MJ4EL)R\.:0P_aH1DY22^eccRACL0D1MUJ62cV9UE8Z.E7bTPd-f?L5^,LSG5,>
9#[#/aO\[+TB1)3f<Qg4(7HLE#NA_D+H3F,a9SG,T7Gb4_eS>_^.EQc;VH1BB7PA
a2O;NY.3^dZ/g)&A,N@1.BV8/Cc&;ARaaHGE9-31WXXQG4fE8d_2g[VOJK29g-DL
dCGVVf_FLbb-K0+-;;0ROHTR?+B<:/ZL0FF]Ze\-\UVLb7^J6fZIDJ6)7C]gIS_2
Q/,&X8([YcMb-@;\?@]#C>1@eNa1B&@eBee.5??We^6NSX+QV;O0/=T=<;_a2ZdS
@\;7N,97X0?&<I7\#>DZ_;P7\?>dZ=JE9/PD_?X\59CgF6+BIC^\M#_9b,:NGLY-
G7Xgc9VGXXBDE:7KQLYLYIad;Z[&>4H0FYR@)MJRe=<IHC)JcOB8)BCYb7T\K>\G
?BUM);VG-;5@PGZL.9X9c7R20?B[Gf(]VT[YH^c7C/GY<,3U&@52,N@A)YD8]K^I
E-N32A1\XG4Wb90VTJ::SeX6>L?ba)4T-Ab-OR,7C-AF=)Z7KYadAf,H6TUI/]Ra
,#3W&)R8NSZSZLe[3S#2C9CfL-+-W59>Ig<cCRRM#VVIb[D+;I/&cbM9-U)B2cA_
D>7WR#dIZC[3(=KgeS5/DAeeC6BC<d];[.5<eE.(C0/aBM=C/;.Xg<[B+1_Z,S;5
[6EYV1\D]X&YK55H[X#bTf?f4(7f41URA6+P(#QI,N[c6U<MSTf>X+4V2GbgBbUb
eP/cSM2a;>B2)b_[J)7bE0USQ.-f<K:Z)C#WY-C,HZae2V5#SKA]Ja+LXPN3\T98
]Nb3NPDK06S\bGF&MQf413RD@YLP7be)9^6650+HDR(:(J[U/<3[AG>6:DMW3EUU
;\S04AL7f4ONN4,#6YR)<79fe/R=[)g.Rg_)4B[)^VZ0N5E18e]/M&AOT+\?])TI
ggN=P/YO6BJeWU_Of3F+N5=&.F=JM/.I27IHFE96@J3COMCQ[H^9fR,0;V2XFV&2
;b(EB/TGPQQK&CM)=8H;6N[[;Ab)eeGXC9,b7U-@&QEfQK7bCS+QO?8<.TS<Qd,U
fg?+2O<bbZec/aBfO7;&_=VEe<5>E2_+_)]--b5#_2>&07HU5F16C1G&GbL1PCb3
Ec#+:087DLAL]44Xf6?IW5CF@)9FT^;1LUI7LQXP=)3&<(ccNZ/a+>R<>Ye5JNUQ
@Y)TS=3JaY>ASS6?#e,C\M3T0=B^^DMg8Y_G[g@YV?4H3@12_;LT9T40WcB]C/+e
Y\@Z=)C>;+Ic/_fEcSb1#>Ze6Z2a.7R8YS[,NKK4Rg:W(31B6I,=]463Xc[W[9A[
.bIDJ_KZ=S=Gg<40C=96B,#UAT,#CGa.1Y(#5QHTEZIaY^QQ;/gZcXWgRX]X89RA
cT);J^):QFYB?O4DR/58]g[d/W&5&FY_HR[Ed\f/:-N-d.,W.R.d+;3NUC-;[AE,
1fMG0IgDR;.gM8=]WG7,NcN]ASMX[Hc-9B;:B0GNA(_JJIZ<E<??0KM/<2M_6[Xc
F4cTFSR]R8=H>BJCP8;2CFB[PXBWWdEFSM)KMWg=O?<PUVLBP8eBU^]G@WGTd+:)
02FOOX1/\G\X^J+X.BfF05KEBVQ5R]<&=)c^CLXJEV@^L?72cX6_X&fUQKaU;/Z>
K4[See0(,,4UNTD.O6BQ?-T_RGBR>)(JO[f[)[a3&>NKB(=+Y#YESN^L2M)]AKT?
8&AeL1.aKZ/<0:@1HVC)+6;>B@UdWRFW-Cg@6O\[L1?E9OY3aIe>F9>:N]c&=O.7
b^G2,aP6JL3BQA3]Vb4;C]_b_?GX#P1#&cWg9.],58JGg&Fg24]\CL)1@b,03.[?
U>bH:9;D5E;5E9:-S]7?9E0]@XHP:N_J[Ma94P&MQA^ePYKU(FC_Cc^ZL=-PE(V-
:ZJTDT>79GZ+YH\<5XXg2X/P-93P#VBGX^/_<EMRYK<W\_ID;(NBTd_6GIIWa@-]
Bg7K&H8Y<4S(NbV6eO_?bgDYARP(GK:a#2(_gQP0[^?,@c;b--5C=JcWC:?5H#-?
GQ6LZM46&#]6BFIJ==U/IbU6._&FL4WNEVR_a3?_d2W+Eb4cRD9OTAaFBUg/b.R2
bZ[FD)OM.]33-2&IT2HH7<4baVc]+\UYg;AC=51^F[LC0:9bZ:KCEfX#a^+=2[Ag
-d9bA05dVOX?636/CedVIAYKQ8Sg7FZOd5?H[6/?#<<TW2)@LQ3B0@MUc804J//O
YD>d^S;VFNJ,+N;&&6,S^@\^6fK<O.g:LbC(OSc?7N_3,&+GJ?1STC>3cNfaEK\S
<[b[D[ZZR.36/>cQ)c?b=T]e;<@2@GSR.\8CG45JMRNN6J[^c.6#<-bH@JVeNZJ\
NNLCWP6=dL&NcTU<C1gUg?,A5K2,KT.?-GNY&X&Vg[1E\J.1.S85I7b?:)U[bSL1
;>?7@a[E21,<de-G.@b\JQ(4D4\UC?gXOU^E3A4C6e1TI+;0./=4R<W?N<4NKg:R
FZM<QKHPS<fce<gH/]#N-==Y>\Z]4=NdCMf(W1UN=6Z5BQ\TSH]>XE(F6;4PYV.<
]2UC1(/7>ZX#OR/O)>.L_X7HC1UJK-\+c#WWOJW-8F_&YY\f7_<ea/JAR+RcV-J(
NWG_W?ZceC1X3SC0=(P3[H;H6ZeYf(O/#CL7Z0;]ce4J3=^W]VMgC9K/aeB12,\N
W6@SPEI=Q4^2CbJF(bHB+&_,P,VS#330^,J3+G+)2fbPAL=0,;S)60^3>U/+d2a]
<TIg3D:2bK.<]S81^LP@cOA<Tc?,Y4U2CQ:fN,<OCc2,_P(,E4(_#UcFCg7]&Fab
TMK/>E54:ACOL2>d.U,U;S[3]e^7S3W)ZKJO_/ULaPR]G1F?cPOd>@T)G;/3N^6X
_N-/EVX4Uf-7cL+8QX56[_CaD?gHM4I-M[1BR+;N1Zg7Z(0d(@\K_)WMc<M(T&BG
Q3DMRIN-OBe5[=]:F@?@/,TOIRYDKgLN5SP#_[IFX[fW4?/E<P?G4K-@_)3_OR#L
JZ7XZ4O_;Z5B4@1^7d]2#We^9C0XKGCBH&EV8R,AZ7C6LdW/T+7X7SMILC+@[=G9
f(X86Le-N,LC@O.=>f\H/9@=N1]ES)?/?GXT,g)IQYZb)L#c_-=UM2SKXZeaST=>
FcC5a:Q&_0_&<6FYKKUc0(PMJ6;53]I]0gAOLeN^<ZH1#0Y-5&P-fS_WXKb0Y7\V
dYgK5ecYdWQaHHU8,<O2K)Q01cDON6=;+_=<Be)P;AM@M1(T5Y4aVD5/4#J.,eQ+
1?eDd&c-N]cF59W=[:KQ^=\RQ3e,5B1^LGO0<2+J#2Bc<:FY6d/-X<\f?8>c\:#+
b;f#?d0+A4OV&=a-\HfCSQN?,<Q(_WP8?_-1^+29]daW<?f]-gTA5bC<fL&bN;5E
I&71d/aPT9EA,-7dfXC0&&A9d^UVg9+HKcVL>Y5>D\@e2N+=6bMGQN,E)LR\?B3\
cQG_A[\B&Ba9&bg/.E5\PP0#FB]a-9dK>>+4g:@>e.(W/,<dG8[D7MP&0G-O+G&[
,(e8M4Hb?6DJ)c;c1VES/S8?9YVKA:]UK@Q#cZ_?;A]dJ-9dKc#a<LYG:P<82TY0
L2W/AQTRTYEX;N]d53<HPXL\SB.1V<5]QI/&G995Va?;Y307^6JB^Ye2cSCeQg8=
2ZTK==OLB(#2@SE^,Y5S@A2.D5R][G@HX_-.=@CE[b+L<Tc?f]GEK;ef;)&.[\AM
5aIA7)3/<W(<FHGJ2#.SD/cGUAEgK;g@:P()8C=ODK>ag0IWKHMTZ.-\6O4(SAU^
gD,e75:d)=H7>J8AH#@ES<aH20>-5]LcMB@P3Y1^bR\KXX,Q:TPW)@c1@V<OK1+V
Q\=/5^-L@HII^]?=Y]0c,NX,@bP.bX>);Y)Q>F.=+Q,AB_N0R3H]22;IE=C4MVSf
E3KX5K0c>Z4=(TX16PZ>c57/TKeKTM_L/Sf?720a6:A;J(RB5EP24MYeZb@ZSL=a
g5RP0@+daaFX3b,&7Cb>,gZcLCTM&UF+fFVMfP1O<WHR(GeF@8<1-<0WXF)Z9Q3^
9&NL+gfGL)\Jg4PB;1c&#L(eQQ&?)-#>S0WefJ51]?]V?8UZ#B<3^YBX+a]2PYL9
TYM:=@5V\=2f>?[(F05a@B=4B.LWB85[\YZW.)Z)@69/,Yg>/LLMB-]84,)f#.b(
[Hd:GN=O/[VJ,L-EM@bJO\<12]3#G5=\O];9gI7&[XX?eNH<fc\SX@/+5R&c@.+H
-7)f.,0B-ILH:=JE/T6S84(U(7TP.baH6M1PQ4/:9OTE2\L2g0AN,Ja4BNQ.FP3\
.W3J&THV-bA/_ZBbK7)HV5IU,2fNN]_NX63_/B8]-O,F(NGAMAL2<6P&\UN&77/)
\dYKEeBO(4dbMH/8&5b12WO_PbJXP+PRdI3/Z1A4\1-,f>]E&S7J.5,EKH#XGK\N
@(a?S2\7D2ccD3FOQ+gQ(Zcc>9c4\J7L2,;+L)Kf;9M07LJePGUdb-QB90&H;J0\
DI(1FHKSbGRMdK24D398bcLLUZ&\aZ=XZ(6GPFA/A,G9]1(aW3BO0adeeMY\.XLR
Vd&387NHZF4DfW#IcOOLTc[\&[^KR[NeZbQ>OVI^4J;Z1E+VQ3;23WTHO6SSX<@c
Z)UOdGD;gfeZ4bd-^\M>&MYY@aeDU?IVK.W;Q.U/M)&]PSc[8>;edN,e:e;f>/MV
@C.g=NF2/0Y\K@g7.I4I+FQ,LOfE91cPX#gL/-:19Z0CW^.0/O)JYA)@5Z+.fG#f
S4IG?Pc&680UO>>Z<O2W^HYBA8H1X(#B?)+\ee9B4S0bf)=,I<.H@@/DD3Yb3GK0
=?<b<.Kb;0,Ga\ERb#K,:fH^;;F,_gQbf=G:7-+HCQ/eF[b[ZLNP)Sb0S_/-.5O0
V(2/cEa@OW6N5c1@QQ\I#UM+3Y]c5@3,b=b[2PDaN=(JR,H]?1PX_.bWW-ZQ+@U-
dG+c<<Z/XH7(WG]H&?JU5/40fPGa,>71CVYBI+CfQ?EK)(H4fJP2R.Db2I-WOW=3
d3V7USHQG1F_M(ggE,+H]5C>HY:-5](RVRg09_W+ZE8\S)G(&-9LBNb.RM43c.+V
&>,PNUDC]\5<(Y1T@XAd8;AQBO1,GXH)E-W8#J(76_R<RM;eX_ANcMagF;+>2f=;
5g2KG,WTT(>_G)YW&aVTR^W2gg(L20dB\]bOeY=5X@dR;:JOJ#UD+B>SI/M]/@Ab
7C[b0I?>(R0YaW19:M4cAT0UFDRT(IK&9AUd02BX2Ia?QBWdEP]8+;-:4BT94BSE
=OWb#d)_7L6]ABecK-^b+d=S:+VFPLg[-B>\/ULO4;65A+;LPVfY>]4C1g2>OO<R
:eCdQWO=VC+@(GR,6QJ3D.UZ-EI?I2OC?^/=M9&XPM^e1:5-RN.Y/+-HSTIG^O<f
<C(KR5S7bPe6G<L]\NC3-F2Z5=D^1J0bZ^(7g;D9_HDC[aT]JSGeg;85^Z,Vf&>-
c6Z]_5B\f8OMDQ)\5&C_]&\^H>0JHR6g[I(S[XF=AHcJ,CQG@e+ED.@X&7[[O(J6
]I)\)gQ-e;fUX-?:<[U9.GcW(Ca&-c=LeC3e4Z<d9HIF<WY\J--K]4d@,]+_ZINf
e0-9_O>5[=49Je9/d55Z6\Mdf8O-,<e0YKQ+#L4AFI6>d=\DZ)ef^+[]1[1+5JbK
F^;>FQ3A4G?5Ra1D5eVd2edOH5gBOAb3&84B>/DM5bNR[[82&0@.:@#+R+JZ?J-2
.6/Ba@D^E&[-/Bc8;QUVAJ1@80c-eZSRUKSL1M[I?Wg(.?MKMFE]1OU=d2)+ZJZ.
eH;<E#[-6T=?3QIeb+PM6GFB:N@@I(:FC=G,eS6]/IKcK7>QKC3LTN.OT>6UTJE9
]#8Q=+S&e+3(:/#X1?=B]=]dJ?Zd63YEC=+Y8):;FX)^N7FKEY@PCP.77<7E/\2Y
N;6.[5M>158O,gB+GCcUCHD.[Mf1A/LR1H?Rc_SQL=BA&Z]N#C)1:@R_-[#QO.E#
OMO1-77c>##F3(TUW,Sg2,U1I#5-95@>W<<\/IZ^CB6FNVDdWKB>W5a#E)HMETM3
2A:9JZOf&+/2XDg]N/OTZ<I5F7F+>[0#UZVV338g;Oe&0>?_f)Q5UWF7\6bdB@@>
N)=AYdPBb2R:X>DU)?54-7gCUaEH>9.:(B,;KARNg,#^<bf+-1^4:MgaOTb-gX3?
,FK1YJ;9.-aNZ0:c1cg[M1<(LF/_FGVd=_C\MNUaAFd11^M=<58aJH.+dOPNaG1C
:(<.QK^5a74M=Z@aI;#_3UWeJA1RV>f(\&aQ1/WA4DF3fU,ZE&DY\;]P/M/+=:AP
Eg/JfDQ;e_\BDG.4C2Z\Q;ITVZ>[C4.1.Wf[VD4^F>Xf#V-O+eDGI/5)ZO=X?@#>
6(L@Y3d55d7U;>+,S&W_8GSN+&L:3B?G7;?BD0[a/]JeeTZ;E:KIaX\EQ.?R;B-D
<e]QNc,TK:@@1?31O29C8\CU]9]X=9Y?A?gVXI)=Na]bA/:L_Q,<B@N4d[8dV5-5
[6T8((1.aLeB68@4>?IeJW2X0fAe,2[IV^KXeG3/d,_eQ;;@a&7#[DF8MFc5c@7R
>JQ@U30E^EfHM+6K47aNAQOVbgSeDagE[6d]D8^I-?.\.&:[d4@1T=)gMf/g+RYE
,1ROEbf_TOdOX^;[,E&C-?(f2?]BG5>82G)2/[B@2/JRQN#XX&JeLJdBeHdGUJbG
aZg,K@@(6Q[f0ac&fT[2/K6L-2cEU6VfB6DQTb2D03W<?_7/Af68bJNEg?>)EJW-
2M4C@/25;CQ71Rb:_T64_;J1:_&9_RVg/Y+HIMN@C7:>@PGG6I@d756T[/9aAVE0
<A_1=&AW<?373;b/f[&2RNN?[0a09:6G>?e#V_S_7B9e1:2104,4(25AWJF4#5_C
K^\\5eO:Wa8HC/X4Z8?][@QgLdB</PD<L7+Xbe]AT,M>8=@Pdf/@aM#.2fHTa0g,
:_/Z&f2TLZ0JW_BA8@bSRXa]@MDL-NG(AAfF3@=V;5Dd\?3A]2K-/0L#\X6),/C=
9a1S<Se=SV&7Be2:3260OY5[6b:T=cc9;+>:I/NaU5J91JaYc:A6X0B--@?/a]P/
8e(I)#@Ub[>(4EAO3/E>=3[gZOK@M;YVgWDQ>R,WAW\K8dOLH5WH&DJeX.a)OC^S
3#EI+305ZG?[+Y9]9GI@YH6:RgJXD>GK-YCUaR-0M]4Mff6TFGHegUJX5bDNedOV
5@cN\=7Q2Cb96RB60A&bd3g#Q[(@Z8V=B)ZYf^LXRL+P)H3&X]IXd]DFdBcN4>c;
,,^)ZB9/eMgL&L(8d#S^a7\1e>^XDNb>?I_O=,]c6#1P,6K>Dd:K6FWb.6-?SVZc
<0]X6\b]9bg,9TB@\.-1:X9XJWb/g4;c.>=-4c;=2\JgSZVB1BdN[eWPV_V_IS9;
QTION@SfJ<WPZP4YE6J6N@KT+/\aJ2df^\]OR22?&0Q83JA5T=E84>ea0EaIRE1T
I2AF4(:RGB50/<a7]9\?g^0K#[eKbZ;.73<[HW;<;fA&7DgL]4)(gMdL=42[08#C
U,JF4(/_&UJRU+c_(6FY;aK@cRZCSE(S:5N>Pcf7(R.).,eIO;.</(aML<gX39f\
B5^46,5Z9DWCJef;S;3))D93&=O;fcU=8-M=VdAE<EKL=NFHaB6,(=g_-9?(b8=>
+SX#G/3DEa2PMC_a0_2VEc_:Q?;fVV41e-7UE6-A6LfJb3COf[Z+9EH2[-/68<B#
[PPE;RF4B;L]PB,V4\YKd9)QfUIHKR7Y]\7\VYQ-]>Ag/X)+A\R8#&WDCG_X>85]
YR3Q/&(:1,1AJ9;a&I=O2a_R,G)c)ODK,_\NGcFg/UYT<=^)\F#8_a(b^-bV&84-
/Bc4:aXMG5;1:gPT#8#;1MCH=bFX>ED:K6O03:1<AL2UUBCY4Z[@a6_b-^0gL:f<
5-O[;#3eS&3>4F;<9D8#BK5f+,GdW<ZBH&+;C@IGJWCHQa.I219YN(L1VC&M<X^[
M4:Y&C&1D+6M50O/1\,-KfP):G3If&78[<[;T7?N^C9RLf5)FTB@DZdZ4M@XXW:A
e-&]^Te7A33,PL>_H/1a[NJ2@f1P#R;>H[?-4c5J..C(9DYO0ZQB/7/-FZ27;+.6
S.ZESPJW9G3.8<YOM)^T1^M:[LdZgcNI+7/S9;C20A?9g[S)+PJ^Y);IeZSad.6^
F\g7D)KJCQ3KedTK=^C2P>]SB6^1B:SGQgb)2H+T=QUP:F1Ya\X30ND1Ze@<:C(e
-MLgd&Kb7,YQO8F9eK_GY>G-:3_<]^GJOLTG/-#_?-:&AD7U7Y0\)6U?2;^(Bg\T
4TQ6DAM@@4,(,[eAOW?058KEIY9.D^DL)BdD.XbYX@##9G37J3^E2JT(d,0F-6<G
Q&36_)cAb\Gc1H;EfQ(./)9N?HWIP1GU&bgXcZ2LR[,7^7:@W7,VCZ=d];=(5g0+
V3;FMA(;?2=6[MOe]A](HU3,83/5TB<eJSQO,b:R/0RYA_UG=YW<V9Y7/]T.(.+B
A^_dWdP0P-=aG7ff2agX;;WVX;Q2,ROJXB_:7D0&\,7D4g&M)MW^756:PcY/;.#.
8HCJOO&g05QLC0<5AB&S2WQ4Mfg)4Td5^[8\0bQ3VT:^.DLRg?bBTVI@YP,\42N]
FIcV66b-9Zdg_X1;XSf<C]P]IPV_PdI6QM#UFe<ZMW1^3&8S1P[JE_g2-O\+@9FE
/ce2=PXb]6Y\BfcG(f_GEECL;_-/:2/<4-?AOgL&&-A^7b)_Vc)L(CY\+XUXNDf@
QOSd3QOZ@POSdM(ZaW,LT3bXGa[4QG)\dA<f9_6:5XQ]M\V#?VeEd\@SbWB>9]#X
e2cZ]dV/UXBe@:?B.(;?\0&<\Pg^[_GfgN?>MJeU>Y9fNC5.8.0GEMZY6Wa+Lg<,
]&>54X73JY_a4A1?_T-AfDRc:1(3^>&?&F8(f#J&d9gPDZ99#NA@[2Y--aE0NNWb
I-:;BHbYdf14=BZ[d_P#[V25LUeL^;1L5>CdL.K33C@NRX5H_B7\QN_0faV2?\WB
X.WBRM=@Mf(YDVa;@33F6SKAK(T6N:\a)G6U<]_4CD-;3.J9HQ?ZI&V:g(d[CI[J
#@MBdU1/cFd<H<ICXeHK8,gOMgS\/F>&V8]f_3+>+]+(+_TOO/6d^Y-/W&K8Y/@J
1?9@DXK8gd^E<U/;>[HaD+Dg/O/K.be.X(0L<cdBNQ/),4^JX7]g+WI6Y8I61.dV
<Y7C\#M::&7)g-9E;<aH?]-I+@L<BH3P-B^_8N1SZ>f9Z+Bg>RQWD^_JK/#F4bO0
[&#^F.JH+C9gY>B.?(CJV-</cfaVg(Zf/aaPD/g>B:]b-g?49E>2(2J9G&CM(O+R
-RY7Aa<-WW0;<PcY44A(=Y3?<Y_OWQ2fdeS.MT-_+<4\eW#6L6Q189;5G4ASbK.d
PMNXf;BM_=XZV@&@)eEN,[][XD-WdQXJ#)#?^],aZ->cZMdbXb&,7bB@Y7UTS[0)
7@K=9KH,ODeL:XBb#:UNXbVOG3<Z[MJ>bg/0&?ZXQ4B?805.^.5=6OKaCg80P^:V
9W^1_gWg:NSJY[\1<&V40^]^1?#L<>^=T7?BfeYB6KC[WfVcXfKO\1M9:9(FbH\K
>^b@DVg(]3VB3<:-VJc3c)_QbAL3505RVc<VT0@E_6b>d&=dU_^+HA5NZE9>JXeI
geC\:R_7DHfRZ6RV.]W2S092V](G@(]-;Q;DS,3bL/2H[RO2=.IHd,,4gN;>Mbbc
8ZbE@9+:;AG)Y(HI9LA1c/5EQ4V+a#+9)-OeY4Xf0=1defEGK:Kc&/fC-/;b.0Q=
+L?\1V2dG8,+;T9H-,H/3-+((MJW._H>2-WES@F9IR-8-->EJ..[GJFgc)Y^88/M
4J9R?aCT=dg0)1FP./_-X96_CC@a=EeLT?CJ(T#(RU+L4&7+>S/A\&32FKe\<;fA
3eFcfQW29d8KJMM[N;=FUYVfR-;K&)N,QbHW8D(HMIgP\:DNEFIJS]f5cF@g+_6.
61&ZZ51<QUfG_]LEJ;0_OT5g2be20Z8Ne)@#-\]b7E>-Q73\(UGZXf>bPZbKVV@Y
^16X[+=S+^IV+A@<C>4dHX.00=J2OXM;OeK](/BA]aET8K4I0\UEZM0^MJ00T],V
A]LJ,?b&]eC+6>,fT:6U1a.Bg^,F<83T9=a73E.]Pc&0O6Z,IX#XK&)\WH7.C&A(
PHX8>XPPW::0_:Sg<-(AAR<&TKgKC=?OcaVC;IT,CYGX>UNL^RUA72-]<L/11[SG
(9d1_R)F3.d.f4S?3aZGW76ZZ8VeZ_bEfb_bP0NX<?U+0_,bKg5WK;TegDZe@F:d
USC5X53HH?<F7Z&,+V<_X:#9H#&LeIfQeZbNH+QM&HVE,Z#,[->Z7e)H6AR[L@)C
8Wb\L8<#DTXR__Ba7DULB(g]KV=L0=7ZNV4<.FK4Y1KUGQT0?AKG@AJ?8F./bgN5
&Mc&62bdDL\77g:I>C2@P,?ND@YANJ2.+S9FNZCEaN/TI]X8KK_NFOBK#P8K)+YE
+F/P:#;fOVQ13@Q,]/[\P4@@FUFX,H09\g43<2NXOQbd1OR8f6UPa^8PME(#RA4]
Y\PgXMfc:2Sc_LZI]35(RcHI(.aZU]U5ELV3<(Y;1D7Z+E\[AS=)3CD4D\d]b&_;
],L<]X):YP2,Jf/#U,0#>1+dWGd+4b99AS-dN^-.;Pfb@HGZ8?d0]ZdEC_RN,[C:
1F;Q^\KVK:IT>+D=[:[D;Y-5D;PK\VR^3V(T82Z+KA-0:XCgDZ?S91]M-?F)LF1<
^VDS_S6T&FK7B60H5#bUDT^W-@a93T=CZ#&#6fCH6YXEHT9dM[6@E4XI(f=;WA\0
FAKg]=]b=RcD@(+R:NbP]AQ+5IW&DR+=OWG3aM?M5?Z]M;1gb3F4HEgb4>QT>WCb
KD^P-++WbQOH61J@^AJ@19^Q1P1L\6A_H[)e.2\C-)&>/G3N4\_J<W9b^JZF5#J@
AHM6Ua<f#3[BN4a,5A9Vbg<13&M9.BX5OXAdLIJ^5ZQ/(2MFMB/YXD=23,f^CCPc
?FC;-^K+Hb#TP:4ZcCQ:IDe;X47g;(gJb<7CYC-FUR51#28WWJfKSQeLf09X\Sf\
^=LN<ZfcCXeI^^#S/bYcK?I,1B1KADBfWabgMAM<EJHM)B/PZQMU:K4bXd@Z1C1I
D-OQ,VVaM:G7A7B,?0EMO8K?F^X>+G/V3#8MG=@\WH-K\c;DUQ?5gZRW^@_(B4X+
?:#R/GKD3YW\MbDK)ZLHcY;/H\<9J<UXQf9CA@#BD.5b^@HGQ2_<[5\;b7AB6U5V
ZC/L;WP>=X6=-^KbU]\K:[3J&=V<9?>g714U<]L[.dC7JL.=4,6;UP?e&\>PWc23
<R&fWR(T7)IAC0&ZgOJF8E(#MNS-1>-+AOD],[dg+BMIKd)=QNJE=@L2^ZgbcK&F
=S5@IUg>\f1W@Z97^^EKG;S5R9a78S4D3^JNP.M)VT>fdgT,IK\&Ie:6-IBB1.Yc
EIaTL\B_ES6F7;Mffd;:aYe-W/4Z=FN0a2Ib?0E]?8I>b0NWW\-:J9&]&=7B],aV
J6/.YSFa_D-^c>^/S=<-gPc\QI59:cd&N&7gT=8KFF3G5F9KaRQQ/@5cC0()4SD+
CE0)#=,Q301-BdgON#@32&&B+]a8\L?d5H/Y3\b4#L;?eUK01U5@51)&HV+VaIET
&AH0[UKaBe?A1)Da1&EG_R_U[N-L<f)WU:#L+5e:IL^1Y4?Q?e&)cT+9\JI6L8XZ
cD,ADBN4\&>[YI]#JIT67T1Cd>-/,/^<cHd>CP@N.^#M2@Z791>+PPEeP+.0[B4>
ZU4MdT2M5<G[/H6?O39[]S-gBGF_Z]WL1P^],HK9J+e32,c(0/C1BKeY8PeWW\4e
2((X=T5/+>a-T=]S)TVGYLH<IL&.7WR^41:/eF&21Q[.ed9V(AI1[UM?Y_a91_QP
ZS7TT.+YS[Pd5&@C2WKc=&94OE0aBMQLL>YXHHW1\>-6bN-fSfUZaa[EEP#7g]3.
>(]@?_@LR3a3afI^N3L)eCU/?-;^.:G73RX#[_URQXd=gS#\-(GJ9cf?4#UUVB_)
Lg]B9gOFf].A-#g?I.<FZ0eYFH;c#TV0eGI\HG0J#Ca+?3afU:f59H;2,;9BE_eg
gg(M3gebd+B?:G;1g2Z/M.O6AR5L9O.76LC;#?P3V@;;H6<MK?@P]2;LA88,SfD3
)O605GC4S&b]aV=c=)O\M,Yc\5BJDHGL:dP_96TL.fa<A(C4(_9:<H2dKMQJVM-@
8FP+]PVOT:g8=e[e8V7UEcVHC27(dXS0)C<&da;-CY9S3XP7_4e/EI_Wf^)Ma2(Z
=gAMWC9MS-JOSS<FgQ-37+eZQ#YT>JbR5S)gMA-3O:Q7e3f#RV[E0C496UUf\JbS
T#AN\5939S+JD#(Dd:ACEQ:>H]ZVcWD5JM30XLLdAaKBDC3FE](SR/0\Y]K0:2BB
dHF6Z^d7YU<DDGGW),8.L8S.JL\?2=_;1LS1>)W(N6CbJKcZDRH3De:6?N]aWbAS
EZIgE:E&)SU?@O=NX#R,(@MeX0\W&2))QJ?Wa5c>\A1_f>#e?PSBgGXRGMV&d-f&
2A:06d@/RHfcR3>?1&BS?aINd>8<VX@I<006QUPL>eQL27U#S-b9#\VZ>(_FMRDd
V<J&&g_1?Xb&1?1Sf6++,<49I_fcVMb1-0g=(WHAd.87M?#=C?d=aL\VUK:cb25U
5\)Z5)07K[ZBJO1O9_72f:FfcdZ(>,1Y;5HQPY>YF5UE2JQC26]PfP=DcX;Aa<U)
O>X&gV-Te<ZDLf0AH-d4IB2SL3-S9F:e/(f;?XO.K1c:^U6d55W[?5117b(31XE#
+-4R;DIN]]\,_eBP0]QO2DQ&[DV\[GM]_5-(\M<(8H>K-Ec,#,;((1b>(3\AIA>\
<-CA&.)]FV6_D#7&?5>WTOYR>T;.(NI?J5^+dHK]8>c]:KQFe[VO6FST_a2T<LLI
^&]8,W;I.UWZ3>U8<4E6>...>4a^0RcdEH)69;WKL=MIUHb>M\KfGY_IC_\\3>=N
+XD:UYbTX5fGH&)[(;ZdZF1c#XB@eJAQM<OQP3+gL_^K8]9@f(K&a_KQ(&D;ST^J
EH#dY-U3d064N<GKL[Q=(N1PX@R,^eVbJ5K2=ZT/+-O3()gJD5QM4DCR@\I1Q9bU
LD2e2CJ-@R/P?3A-FD1@0^dX#;;N-HZe/Z4\U(1\:dNNUTIU8#Uc<MJ?4X\@7gK-
,P\U?+QNEHA:9L)P;E((<+dOI)+TO[S]7/Y-(L2f\5?-J(3C2):B6Id76KMPKc>3
(+#8aQ8L.fMBO^:48:e(;BOb@AaZKUL#<.5;1:)D24Oe9QP.L<fFV+-bM<A4S[5T
_:TFeAOYHTK_6EeUB0@,;99JA)95RUWfCbJMBJULJQ7&=&9K);P;Uc(0K50\M2Rc
3cMDGbCZX(7;Wg>4>S&:U0X[,9472^+--TZgcCb]XE8dA0^#30/+eI0EbOX4e&KG
e@2LXb0N1@JdGWdc7S8:3[DU475,3F?e)A68g-C4-SaeI]+D@(dNO]G8-;N>SU38
gY]c(H1X[_<\0U3gFE[+bC9<&fK\MKfP3XJ#;U6)e/VN=W2Yf[Fe&@IUNe=-)U)U
UIZVAF/723.D\gS[.;V)#A\\D5ege=H7Z,V?D,NGBORfFE5ac(K3?>BJ#L>L:c4?
/W.\>g&24WBN8Q8;5>WGa1aZ]Z,XHbE?O9GI.GaUfX27bQI)@_.@64CB2;)A>6bO
GALMA[ZJ_D<,OHb23YQ\&e-CdbB4c\Db_g;MQ6c.WJX>[_W4TOdHgSd9\;;_#[/#
:eG#g4#c9_;?GaD\AHKU.d19KUMNM]JGNaSGD],9)577B#B-d[_+4X0F\g4OaD[e
,N>P<=]9QH/XSEZQ<bBC_E#WEa.[gR276?)bfH3(#7\V[)]cf@W\a=&8U7fcS#@;
Pd[R&;d)VN@4=NaC<)<MLET;N\;dM6CSF0HCG&9T,++gK_Z)2fN)?>N/#XDF0RE:
a+[^:LG3TXcS#Cg<S0UDWV3ff:0-&fH7W:6(;625J4f^B4Y]dF-&P8]Z-Z08\O4Z
fV6>4X]J2WJ#bGcS1WSQN>VcCe((A&e8cRb2@8&Y01cU6cS?LS@I@F?&0-KFGAI5
T)Q)3a)e]^08#)B422)\gYD[&cED?EbIeRGZ9T6&f.#UIbg>dg:_KeVJB38-JE/@
[8/Ja@.3YVf#(6^M@5>L(.TR^c,c-&P(2Ec7=MIC67\7I?]RCd]QaL]RQ.N3CSJ-
A-SS0/&#0Yc<b3C@c/]EX2-d;[[/Tf<<GW5PN8+F(]EZ:JaQ4WSd>PUQ-?K4@I]b
BF2-D(0(B.>]eX?&SN;/3gb>5g/[@EA)H7#4A84T9TD@RGL9gV/C<Xb/b@0-SYe:
;Xa6GD<.G(=#NY0R>#POa?@>,3+)a62e8^2NFNKcDX]-9,EE8P5EVL&-_;BZA?8F
cF4fV:g,QKSHLZE01G3,7CA,-.(8WPX&^<+QP)MS9(La-&?\.65_:&X+3^MKD<((
5SeME8I^8:d1_[3JUU;G-FQVLC2TG7@7^>QG0ZL7;-RJ_]IPe>WYBXIF[c1>B?CO
E6#>_/+fQJG;Ef=,ce<S>A.eWGf)/^eKGUDO;bASC5/=R/_5_)(Yc/a/R.fA<S=P
dE?C<g=H&PT-3Q&_8>0dQ[)O[YCYN4,2WgaBX]53SZ<bMa,P[CZH.aT+.a>MG:FM
(aH9Z-BL=PZ7:-AD8X:3>b/RN6,8Q^419/#=6=;Q&TA2#FBHMIO4NJ0(NeMX&5]<
Bb0&@\XZGJf]2)O1a(UO2,B)4?D5Ya>1+6Z+S501,3K]D5=:PdfR,2Kd@6ET=0HZ
&H-E@;1dY,QA5NR-\OZPR^SHdT;fEF[;Zc?-fF9,/H_bP7->C81;b6ZB9:)N9Ndb
:]Ye^?9[ZSWV\fVAYT/:VD-2(SJM7GGC_))RLC.?@54YGb7?A09/@W=f0f\X-3Z[
ff9W4bFTJfN>04USN6/++<5:5&:M+D/+.gd)_W-W@eXEaS=SgM_Mb^B<SNOE3aJF
7,W1c3D0(M]:V?Y<a-B7>R3UHO5-eJMfE58,2_:cI.@fD&.F(:e0+6+])ee7L4P7
R\P?]25XDWV]\KVVPXLU_MW)?M_6Y&MbQG?-(:@I6HGaJ@10AW4:A4@V0VXU4Xd<
.-A)^49Na(4EE_J[3=B,#19ZeUWT1B=SR/b3&dW>TgD2R:VR_I=MeYfAc:)\8T</
@b.TCID3S^[2K-/+7I2;g.SH]5c\]DgN(48b5cG^.,]c<?)e1UW-gJCQT>)#MJ:T
^(57]3XO(53W(DEGF;.,aE@e\UIc3]6NLKabL7aU30=N[F8H68A&EJWWK0U5J,Og
G3+U_9G9/;JQ2KcZ=8((gO>5NeTZ1;:U(Z\AP.F9^NCA:XS[9,O4f.eV#G[dGbJU
>,X?IMWS5<??faJ75(>S&_#;=MS=KZ65EHX18C]RfK^Sd;ZP2&)\6e)\K_#XN3d>
^4I@D0VH(,3@_[<cSAd9\K28UAd_ZZZ@f)3HVDQ#Je5T_;\dR+ZfCd<KRO+OcZ+g
e#BP/@aF2X7P4ETME6A>5>775JO<f:-^<6K/#=TOa:(F))T;gfg-TePD2c5fSgTU
;.d)g+F.&VdZ4>P4DM=2;8QL==V(;^;IF.?C#AU[+d?L.QCV]GK,/gTS[-cH#-B8
WA3KJ59CEZ_e6KN7c@^3Y2)_KG.fSNRE2_^XG71K7CJ.4O/aRe_g;FI@UBcc]8.d
YSSaEU+Je^U.LPZ(:3HIX[?8(YJ>.E\B+])]CH:TXR)RTbC?\C+C.cQ=gKHY)GN8
/&2E&;RF[]=7O)L,HR1J3N@S-82:Z(>)L&G^YBGEP;2H3dC7(]BO/SLKHdOYLR(S
S@5Y&98AXXdVG=19R>P5?\NB7J3^KTK;?3QdS7]F1NH&I_1Q7[B)T0eW0^HTfFL=
)SZR0(Sb7BcUIJT^M<[^JS5YV]_RKP+;^MLJ)]:2W7^=:2@AG@NG[:[6gd#.a60@
2.],Y4/4cYUC[WBX#a@7D4BN#WUTRY,_UP_5DJ(W?Bg))3,0+g(f<#2E>1JA8&U1
_d>UWM<R(P8g;[]IT?RBC>J]\.;Ae;P>KcEK5>.-]QR6R(G#]C[]7GA262]+7<a3
(f]P3I#UDW1D:E=b<8IG^:ZO<V:9E1eGb\IUOK.2AT@GJW9)/G9C@gYN,MKQ.M/\
aIT,7P79O70GFZ_dJFSZ2O\VQ0[EX>L5f,4cgP-7PcB76KY3e6>dR-#<4T,O6gL?
-?AST,2N1/14\,VAgTM]5_5;_8,L<GMEAY,>B7H\6/D1[6VHO^+E\LLZc?8NO?b)
^K,a#3#5(O[/c#Bc[2[ND2e6,W=.Hd9T79H0S;#[V>5QOS(/>ODF-R.Nbc-M\X9-
XdO&WXfe:V#--<&>[A^]4(C#Z<7-Nc,\Y5bc7SJCVdg+^@/91Y)@b#NB>f]V>J@?
H3807QL)AM-?9>K)??Yb.@:([STXe15(_T3KI5]JQPNYT1g4D)L\X)>(W>QP)PF9
<Of=.ALD]?e1<R#D\;fQgb20)B(3C,bLSS/fILT;fU>F,</>RT;TY@Vf>V:Fd86D
f:-#7bGD)/M>G[PFNN95PNIBeBE(Z/O>ZdF9>=;Ld8](TJ,]eYSUUWQROF;L1)Hd
M7>4dg@16=.-?e#e>b<8GBXW.^0=cZ\<ERW59>&N+@g9>3L?XNKFQ^\,;GL=D8@?
;BCf]#VS])>E1F_@gbAPTL&0CHKF\M+ZAG&[T]M9)JLBfMXLS?JTg]+1>.6C)fDA
fQ.=)A22+E:&1+_<@XPY,#]Z28Cg<5CBPX7-3dd\XcE_A;b.2+M\CPNfR[8VDe;O
8JYQ0D^7Cb+-TX]+9?:+XD,_18C0(<V@e3)+W&<_f8ZW_#IUB9G=858I5_aBeKXL
[FM^+@a75R?,C@6_C30B.N/a6.36g0[M[?TK:eK02HV2)eE8DaCPFeIgB^d\SL.U
NMYMP:H06Q.)2J<#NR-f#@[V/VYH(]VGM?.M82bXCQc,PL[bdKa?JcI^RB,7GOB4
<+aXRCLeUNgbQJ;LU,G-K3R@6KLM^NKT=<5QELAYKMbU2#eA6N](,U-.Y.0&M80<
g:QBT0LM5S_>,E,X;MB2P?bVK_WgVKdd9#OaOb&Wg/=FHS1O)A;/[;cg\5eU@aOd
Qc^JQdA8VE&Z8]g,@2GDgDVNH89(>3&-A1aC)3#N<_e(Eb5J8]3:#4HD7W1X?5QQ
7JWfTEZXML28CX.&g+5+X&&N73UFNT\&D+c2:bg7?IQIaMU-2(KZ.<C=@&G:&WLE
b<1Abd9DU5-cX4]4HUfUO-,=T8Ed[E\UV@T2#]<92RR3NE^40>R.-]+M[X@?R9<R
A2TS7?#7],)#+3Jg0@(5R^<=<#f(M=(:_CW]GVE<R&Kdd7568)-H&(CgUTMdQ84f
M1@cR/_[6e/==TA\MSC327[SMMAO_@>ca_HW>1UL?D98-KbB1T>)a&(IP[_Q8V(P
&(+CFd+#3KRd]O[@U3KJF9Zg3EL6VY==(eCI@9TPP5>^)caN-3NHW9_8N;3SU-H_
/]-#Y_+G&TTbQ)B45#-C#eG_B-cKQQPK.F6O\D6MGAV/E-##)gWY@f8GK^N63?e/
(a90N3>L)]C:fV)>U3TeP(MK1-D?feVV(Z1Y=@:[\1_F7\BgEG7J74.FWXfIc6@9
(5(XCeB.aKQ;1]W[__K&/HJ?.\=>-D+R^T(e\a48G.D,B088[f;3TH&+6(HNKF[8
2V;)dJ\Q/0INcTd+C,+6gOCfSV0Tf-7dcY@F-#,3GK:Ug72ARHXcRT2K/^+8D[O1
QI@E@8_-B&9[7a:bKdML:Y0(FfA]H0Q)K,g_V[8YGI9>UW+IOK5)Yec;J9F_;c9,
9N]S,PSfS,-X4+B:LXg5Lf18GI5Y@O(5PbZ7^eVQ#>S^<B::SI>T-_fU9QVFF/e@
N72^6Z9.>5R0Pe^4cV\S6-1W4Nc94M]f2#S=gd]UC(#X4;<g:];LZ68(\&]gG>XM
fFEVT90FC+ce[ERZ[MTMHZY]J&Y&W_(4c#4:9HSJ?YW94Y/TU]C#04==1X-XQ?>&
X0V0=OTPaW:>+.VTD:[5Z/.D-<]+Ib^@PMXccKLDddF1W-O-5-N>N\_)Y/Kdb\T[
Y@<OC.O_65941&7U)\/6PM)cd)/dcOfY[&6bVC2/426O&4I;@dE^=,\#@dXSWU6d
1[D8?(Q6):O99S0QPXa]eIMY9HJCaO00e<5@PT:P3A&^^YZ;#Cf_>)@>RXL5NgP]
2\f5=:JMY#c4B-W#^NV,38aLVV;K3<GH^]8[/^,dYfU)N4.@XH;3:F0BHMHR6BDX
c[M9^>^8T,f[;O2:GWW4&7Z6]<U)+c39@B-I4\8]eY^d;U]EJ<R;Z6^,W^I#P,aO
KJN<7_Jc>Y]=B?7,6?_5R/1SJ9WfST)^fPCCJRWdKf^Ud,UfC@#X[Z@F8YE0.DHJ
aYa3>Hc1^[b&aT<,_W_^XTWWRCRd>\a3?3b+YC/8X8>S3a\1+)d?UF>JT4H6ffD0
+]B#gDeag]H;Q^Ke^Q:R1<_g_6YX0\a8FgDdPS>(?.4(E4.;e&HL=<G4[_f8aO]g
79G3/(Zd_=\b9-3N^.HF7L<18E6OSgZ[M])D_9b9UI\SIY,(Ce6;B[-CJ&R>AK=C
R7S-7[S:OLEF_7Y8Pb(PKK9\+AB-00c#].NJE[<K(OdB9.S[OC2Z/;A3@6F>4Dd/
1_[\@/,5==XO;aM;@]N?VM8f+@5I[GUSY(CPY3-_>]8\bFSga<1A;=ULI02&9,NL
YN>X./-,F.N1.9cC\FDg5.KB&+H3:(;KACX7/BBbVQD<eJ?gf.VKQHX86;e[_K07
#JFMAdC4Z=RJ6U=3C.aA:ZD8-:6C_++Web@LK\6E)V33<YaBaC0cK2U?6H54HS-^
2=0CIdB+M6AN>780(+J@MeB:UG9&#V?^K1#\P)711Ng=#fd&BI&,a]<X<0b&d;G\
9:@ST(9UZ;4OR3+JJS-1&OS0gEK?7_EUO(-=KIKP7(CH71JE@G8F-C2.0AZDJb=K
dIG@c\;g2_CU/Aa:R.VTHJ_e>Ed50_9I??JOTI#6#.N.a+HBO\U3Ff5beXZ/0ZC3
AS29T)V\CdT7Yb=Y3&N#YY\c019)IMTD+S:#=?PHC]aJcN3GNSYFRDOPP,EEKV?O
NdF[Dc,0bGC5#Z.88SIG^YC@0^3;RH(O8YWMa8042,(.&::9OW41/-#ZNUAFbYLV
Db@N-bd0e8,D^U2:@-C7LI0O0>Id)>F3)A28H1H<.H1Q?b.Z++;E)c>R(RCf4KTC
7=<]MZOG@,)C=0L984AMYEEOf#HNd-<+GVg6-S#1Q&>X>Bb\=A)Y<+HO45I^XObT
>,T<44B:,)\@IK;UMU(PX][CNb_N<8O@XHaQ5F:OC?TOC9dTa3SHFAf\DbZcGR]4
ZV(.gW:a#[-HcLF\.&F]YF=BS?\dWefLDPV64]3eB.^E?_=]=9H/aZ;AK.ce5fWY
5FIG&@\HFN7)KWSZ&\7RPfDT.8[#g+L=F)D.eFTM);.e&b\6^g-aB6^MODcQFF>:
)c6S+[f:.ZW5bT#SFRC@#-@@1X&+6JWOHdKH\g=3G-2MY92:\5(^-<c#gPVFWYK_
;c)?2H[Q.17S^:c&f>8\FR(c]\NIV+g#7G]##UB:Y6BdFFc3d9M>Gd1_[X&=[LBJ
aD+=<9WXNY#d9(7e1(4aXT#DY75@M;f#7Bg<Q:RD,_&LN,CcDY;LI6-gLg74CVBf
[cC>CX>V3WFRVW+0BRcfEHKNa0B-2dM6O6JW;9^8M9GDeXAB#_&ZK@)VA19X9.cI
,\U=X82NN?<eg-4M_dGT+-]-8_&_BC-H0=QXZ-\Q)=92\(X>^Ed@;LKaCU,7BYg_
J]c_:Ic.;F:8OR^D)W9QeI[98;J0/MgI,YYd\9fADT6TZVe\:G>]XCM#OeXJ+++]
e+[DX(aVXd?=feIE+eB,2EV^>]/E^3dJg.acH\J\,Bc;A0WLYc.8=dcbC.RFVTBW
a:>P/YHSfRd4TG):^=+fe(K=H;gU0[Y_Y4D)>AR?L/[<IQT=(Y5fT6@K:#-&VEZ&
TU5--D<7^^QYGObfC4=-^EX^WQ0B6eE6RM<,]R?O1Q_-f^<_+(NY/7O_#Z>H8?>G
Ma+X[2b@EWZYI5g##@B1K.:X,/T3Id;:BW]P4U;KM.P8MK\_JXQ)H.DKg#?M>f&(
TbSZ=Tg+ZX5Y[:+VTMQ;,-.1#4#H.aL=T7<[-4?XT(:#,OdOgW@8Be]W>d[V:MSX
XETL@dZD5G8#.JOeNXGgPb3)dN9Nd5DJ^[&a2LIbVAK6[RB-T5H+-QaHcN1E@RJe
OCRHR+ecY)[#e4<f+<.SeJ+TT2KS6d>/L]eOd+>LQAC84&((bCbVFTU?:[3=aGWF
ZIR&^331>H,YJ.F>K\\4;[=DR:;#H@TfOA&^B^&S3N&LF?J3G\IeE69]36O]+LVH
P#.J;]_ZR[Z]ZXEH@E1EY;]://Dd2QJa^EH2\[YA/1;ADSDT/_6D\Jeg&.aA7F;T
G3dgb01@PH??,4W8KZb.AE^0)GDH8Pd,N-7[ccK_UXYZYa)@627V?YCSZN=N]f64
XUd;U;BWWV>9H0(gLPU08/aVUX(\#9FD9+Me]\>_+(618H,?].d(B+8K5J#P5CTG
fO?QCOgM2>/(A5/X(,AW#^3W8d)AQX+fWM(30URFJ,J6MY0YXEC9:Oa=]\<TIKNM
L_a8(V(E:7G?;#./LO[eJ<_F\9SS5B>5TSM3d1=)g75SYA11.L5QP_QC<bL&P\(;
=CKEE3HN@d\>;W_DdS<bB&R?-^O7,-KY6Y,)R^3#R-:-bg:LXRV,JW42T+49Kba6
48GP@J0TI^>H&A<,e,[@5gCW4c.6_Q^X1AcJK)MRcX]F+^d#^HF87@<L\Ra29+Ta
YYc8DI-9\17UU9NC:DB,#I0a=M7&79c@V[BdD_XTU1PBWYQ&X1Q)^OQ.#06dZ#Z,
GP^D.IZdS:g(9YS5;1F,T;Y9,H#P?K.<a3A3e,U@914ID4X)4b__U<ID=WVKA6:@
#N&TSEZ]99->1#Y.&6=/;_PWOfeLZ6PW3K4F=S)@&Y5\,]\2WM7=Kb0R]+3eG?E]
7Lb)VHR]7\DGPG\@Q&FGB_NTHeUWC/LRLGM6\QC9ER(.N=OeY]HT0-]9G)0BA304
KV/@_.f@,/7R.;?V7GB+ND91WW4P/7Z7gbHEC8&,PA^C&(+@Q9M0OXQfI9<+WBdQ
&Q2.47#0_f4e5b<)&X&9FMbQ(HZP4@Tf?P6B:M]R=\R4Z#bWFSfQDL3.TL<&H,Xb
UX-;56=XG/+>6/AY9MT>034(8+6@=KPOX8)Cg:EV/+<6b;8b82Kb[_F3eG(OZbJD
_D]DJ;95(f@:)4]]&9b<gWCJa7;f)258:TTIXg5V85T)8\V[XB2Na\\@JC1ZX=U/
VdI_BI61O6f58@Z/[Ff6F1XEWUC#2(C#R9B/&=/fUNSZ9A]PW_Zf_DP1^_\BGHX-
d^f<C&P-=-);ZMX>OV;FYM,:\d=17#I.Z4<MX-1UL<?5>2LcN]QBJ59YKK6#f1U<
^d]#04+&)FU;Z4LZC[](?I5WHNPTY@DI2Gd&6abf^C]7@6.[P>44X5-^LF>E(6[)
K6GC?+Wf[_?:7F/aZ<?LQ&Q\/22D4,QOK.)?49.78V6#0cN9JQ>JO3I..1ECASZ=
Gc4E(ABX\PIC,516::IC<WCSUPC2B:0c>QX[e<eUd3#WT6IaCa>M69;M7S58&=CC
NeG6(KIe(OcY7P>XIQIOLaO_9+I40DR;JUGO@Cc4J.XcG^TXRBAF50FTBd7-RY?>
#1JI\ZIW+:?9N,_80;HMJ-2B_;R&-bE;e-:;]<a1)P+LR3F:Xg>+;;3N_<@QfE1L
1:&W06RRK^YYGD4bgJbg9.[KDPP__#RG-H+f<#CC[7&KJN[7d,^RfRKAM?05P_:X
^\AN83;[,O-78fENP<^R<V2LY:HFbDF<XaF4/JY9<#Q9YdcG04SWE?DJDB##]J9X
SEW\egK2+<(5R;#73B+&@81?\MK0_;),[)c27-C39Q4/42-b)^[Abe8S7ZJ?G=PD
J>WFZeC-aRW=4F>0Y-2\QTU,B[GTPfeBb)O\\8:C?CNN)E],:gDB0(=0E)G1.W:P
K@fOYdg,4:U[,>>1,)(TM_BU<MAdSL/LYf;5+b-J>&Z.a[fCP?Me&#_724J>X>Y,
4)YLG/5YIaVTQba\JNdLd78.UP)-Mge>#2Yf:.,NK>\R?244OZR1dQaZ]PY+SI;Z
d4M8[W]^3QY8,eD^Q_6G/f(_8a<RLMM&-a^4Q,Ad8(gE+f+dg:PF<6PGS8WF[FRQ
;_Q60LIO>#Y-]<Y[IGD@=-G#QCWKDJ>1d=FF1W3&eI6U+?BO<bC(2_Z;,[P/Fb?S
eGKNc1&6PBCDRZ6U76-#H9EcH6):Q+cN?OVX>U;]1C]:gW/F>:cWQdW0;,+7(F2R
AMP/5#g/NfPG[O[H56OI[dK?(/(3;aZUUG@ATC:WX?IV4Q_?1KR>H_]9T590b#0#
95#PA7=4+KgYHZ=&ZbeAB9M?&Y+E&I.24.>&8:;dfNV6G+40.Y-U;Kb7E05Aa=B8
CT&(LC9JH?KZA(cLNPKgBX&-5+[V8TD@4I7V;c0#G=[9d>14LLe&RQaBgcC+_/4M
(^),T2,fN\W@0TDOUIQDC/7;B@VdQeCZ++HKX.CBR\5U30C#DCXYY_dcYT.K(bfG
cT(ff;CbAaS9>F-I]5gSK:VA@^N_Z:^M1AUJ43.=LFBU_16>19=OC@egM@EZ;?8W
SL_J5,>-8)ZKZTNJ8g:K3N[\6cMMS1(29[+GSbP_bd9Ja.EUg@E7;6[YFd).15D@
2IVFCb9bZ2&bdF2]CbY<aI,e[5-9)J)1YYU.a&ZNO8)R[:S_Q]e9cb8^:7cDHA.<
GH#24MY1KG31Z#_,Z_U9][UIU(O0G(/\P0)+U>F_c24HCKf[06b^Ka@OIZGSZ?F9
KKIC.,eBA=TaK@f6:cT^533R@M493F^eeS(KaC3\K3CVe)PdL>3#>3/deRX)GF#8
DQD]V@.#=<DOfA0)LZO#ZMUOYA9:WO6..X.KQA=Ma8YYPH[/.9E+]dRRFD.BeKAG
d6C19Y9DDc/=]I07XT[4gdcD7DJTKaV<&+fbSe7I-&U=?aME^>c)32#SCVIYKKJZ
)@,e+I6KTE)3&)[Hb\;D1B#N&6W>RGSeDPMdJGaM\C_P7KN4:bF4O&&W6CR<1bb[
[JF55/Z<\M1cNCe?8?@5226SVPbGZI7EY;c:Y6<NR0cKC0DA\AbDTCFT;E9-6[>#
#UN(aSCV2^#(3G=RMP<O(.TXI##C:X3D?J27H6#NAE)+IdE;fS3fE1FAPW?VV@=6
c&d3GY32eMW,X89A_5d+P91WJe:,;7?dD4-QZ>JL_)O+)0]Z<;O5c]bg:BVOHeDD
[_cP-3Z.)9Q,\BU;L_Q.T1V42cL(4CGH/0J.&D6SLA\^aMZIb01.1RdBeNd3M(ID
fW>[d,=;_X[cO,+.CS+\/gN^BQYRV,S=e<E28UG;,cLe/DH)3PBS.(?+U+?fDKAI
IcY?)/OTKVN,==/V:NA4LacCP6fD->7]4g_=@\E^)8,T5Hd8aDUJLMdCdFJSQSb;
a]?0V3DDY)QMF/>V)?5FV-V-a_7@75/Y,-Q<FTd:HC<LJV^1_f<&=41T7J:PZaQ+
ed[<BP6bR=B^;SL8FG@+WD7\3\2G6309I<XRJ3ZdI\M4_#KO]5..aVZDVZXe;=3a
,5I3FNa-A_XVegKQaNKde/cKd.T-;54W8[a#bDK[gDPgL=>.a:N_Aa^CEB?6ZN)/
-TPLF)/L7NV6\;H,N0O&,7->fd3(FfYBAS(@]<CW.^4A&JSY=+@C#<9WQ#CO[_g@
LW/#gQ5D<V,)ca/P262@e?e>\Y8T3XU1J(<QO0M&,BQH.A>5c]1.>,\c?H)=Z(&,
IG1GQ-+a2?D[F)\3QD?OK^2]A9SW>df1SQY<,8G-O5#MJ\2XENH_C)1bAaJDEfIO
QV?F@d2Z[OA7NJEH/G5Mf9##\FTS&(KYO??N91Y:aegL.L6G+2#00^d9N;IW;e=B
^G0XNCZ5DGN.SE6?5=dE.,10@8M9UQH^)LF<R#Y@HNUEP#f]&NJ()+aN<;?>)S03
Lf&&==_\Y@SS.4KFB7;PYCAEL:RSFPe\;:-&:TI,<2FD0\#CR(U-(3R[4H-fE6.,
9aLB7FHD7\+#7KfaD@d#&_[V)_6OPJP0=W5V)/Kg)+=<X2HA^8[;0#aZ-)&/SH8_
,(3(1Z.NeH]QN[3P49KdHNXgecF<C26HD@Pb]?0?a)D?1;Lb8(6M[N)KL8H\D<H;
2[7aBaXYAYHReZNC\fLW&c>TKI+&^a^/cWN-]KLa?IZ\@VA9)c5,N)T)>PB62Y^a
8+(D/#e\<78GD\GS:fK^Db:28KW6X#)L4&A4P=M_+,W>PQT,aJb4E(PP3gB-;VCB
Af+?Q,)a-&dG\M?9E::Z+.8S<+=Da6JQ\V3)&Xd?.FZJ5T5H<)<Y:UMJO2dX</HZ
EL:cWU]RcL-Lg,V]8YFDRW4FVP;QGUQ6:V)9fS]E=gE^)D</_CY)W_&RT8-(aAeZ
J<?IaYAX1K3UAcS\L0P1ZL3g^2K#H#^BIFeTDFc-F8eGG40,_b9:?a]Z&^@g<1?@
VNIVU55SRbIeR/Z9HadPPN2.fPGf#B1c+0A<=cVK5f.B(Te<@KKd:,X77faD?W=;
ED3P?6Q/PRMCUf&\UF=WFUQf1()/<#.6CZNHbD&]aI9WA4V96[URg4?0=;T.\9S5
#WD(/66ONb6SRQM]e;e#.W-fgNN/R5VVGBH</cEaT?(?5,SaC>d7=89(Q1&S&5(9
#JI)(,df0[V:5c1WYEF]^[gB>LG4R\7[KcES+Qe#[=ST-V3@(5c77a=HD0QgYE]?
#6HgU]>#Ade?R20Q)8)bV0G-,6?,(;gHNNJ=B9cF/\O+OAN<EKJJ)\^WQ6^I\15S
fcN:P-L78XBM2JfRVCU-g]?5Rb/OYT/ZRYfbZF8W([@M;a]DJ.[+eE8XB+BH^-W^
(+HVYXB>MfI4f(Bg4BX-78.Y:2FLda\>:PPKSDbX7&.TfCSFcX_S+23MX4:\#PdG
@A8BVBGL0SJ20?dY^B.<Z;AO<(^E^:cWM7/KMDUA85VCEf<^-.7MKdU^BQ)93^>K
3A:[QK;OH+1Jd^42IOI(O[IbQX==23M10TV95&)0DTY#ICff6J)(O5S8]FCQL<;>
X5ZR#T_dJ0?T;SZ9fJ_5TK5F18>Y=.Z;Y+(6O)0UFgO1cR,ORPX&,]M/K#7(3f^X
dNV5S3=bDbT3/_.;X)1B1=A2Xe,g41[-A9\&&9:X2)/g_7]ALXRS;-?<R#79+RPW
U3Gd]ZQD(T/07ZVa<^gB_B1M;gM2[_PP#,b9a?<Ab_[2B-UB4D9<cL>ISD,&@=YY
C&CRKd;L4,@FQBeL6\2?d1ZOS1T2OY@W0,9e=[)FQT:0C>)VV87K4L4T>dMd)fM\
W@FdL-4_66TL[Fb9SK4LIfg2[S,_K,+K^]9?+0_C\fdg<R/X=(6?WMa+b\eT-4BV
CXB2f^<#0T.9]5agg=#LYG5HS@1a<3=O?KL?BEcS?>8bBf\\E)d7OX)d(0:cCBVA
J87)9_D^5J-I->2AZ9TE;7?XbJ0J(AQ)f4I;A)0B,@g,CKF_G+3K1#gd_?W(-g0M
_d8/6;1,+Z=JEE/84c+\3Y1[MPHW3b;E=g^SH8AV9bX;H;\YgBLNW?f,RJEaG&I,
BW<FfPN.3?gQS=LV76fC1HHM&XfK4G^(D_=0T,<#YLU@^AIBWT/.[&0Kae0]fL/[
eO;;gW:L/HaCO-9A+/P5@_fN-[]Z9dgV[##VE6]#,4T3;O7Z6:=1?&&4dfPR[[IM
YNDSg9aH88gR85.?KYFVK+62<A,RfHLWLXA0GD2D=B=_3;T_OU>bSB8:dD1,IE:U
(Q]#&6GDD-SCI[b,4g18;G7#JL+3^.Mg.?/8;Q6#bPL782[2NUEFM0/AKc1FI/(a
MT&d@^5P]I0]3OZ\:HA(VWRF80\W]F32cV>SV;B_bEU]C@7#TP&-]->]CM>UR\bc
<HMJ59^A]EcFcN@&V;;953abDYF59B>JIHbPcc[.f[OOS5)8de&eFGO?1D,UN]@Q
8>;Wf9O(>INaSe][K)Q?Y2aBf4B[c>N-d\64^Lf(SW5<f79:G]BVST?KfLF#&;F&
6a;NV2RZ.-gg>.C+]W0deLeAEXKY)JVa_,R:?7R42D_OF6?]8#IdP3WA[2E:I[L0
E(F(-Q]0J+HBQ/DQ/&=5^BDK)d_<SBNI+0/TKBYU6&;NYA(6G30^OOFe3;cARgBe
<X/d@>]W(gF6^<_-XdY[:-GBeX?dN@^ZP4&6U,^S>/>?JR2K@L0@KQIZ00WaRI?K
0@)O_5^GL]6RB<^Qf.80CgAOA;93@.Q70E\07XPX<83BECGbe3T?1<</@GgI5==I
):B6VDd0\-^W.P7:.)&8SYF6E4#,FBJVXJ+6EP,f3;V0S\Oc=_V:;5:_]\=P;5:N
EE;Y.5CgBbR0QCE2P]</1W?8.:UO]H+X@(VcKAbC2Q,5dGg(9^.dK/>H?#/Wa1JL
U9f#AcDX)ZX[c#a]a-[\?3^M&b5R?(3Ud79E[)XB,_OIK>OMc&-dZ5>&;G:C\I,>
GfKB7>C7#OO:#B07(8?d=gM-/0d&N72Y1?\4X9D]G97PRV)f9a0CeK^f=4N(1Zg.
5g9C_L],T-((+5>YB0UHGg@fQO4gIWNPGg/DGTcM[,.(D57..-WBW^11ES[H_5-<
DCef1gQeLT;6_5&[(<Wggc_JK1gdF]5Q>L/[Z1]G:A-)5d3VaW3Y[U3J5TYMa#9?
aQCf-KbbbGU,<S@2WHb?4/b.8KRIWF.;=.>X;c_RadNPeAP+M(8=dHacH&bf0A.K
M:7RTQU:g^ePc_dA>)e2cf?.Q:)4A<VLJN-)XZ#?U<^eR\H-F<O+>-_?U0-_SB_P
\_LK26ZH\KN8e>g6H\:[K]<Be#GS]N\<I]ROa1/-b?eY8VV#:G#d6:RO4(W\;-RZ
)MR]A@@SM:IM=5af@C0?7@/VSce-QaB=G/#aaRS-D#9NfFV/)XHYMVYR_(Y1_.O;
Yb\5\:WYKDNU67c00\568-HM]ZDD@=VX3AJ<S2.^]T[R(^c,E.KZ;ZdNWd)7K.H+
1I\ad1S0;+)eYV5F]a\;@6fAcH1U]cf(R#(T#22XO>cR]IS4g9KI/b?g,?W@:(WX
Gd(:6(E/S^34R1_3YL[;7<Z+,<+MVA,LFM>4=B3.A[5S1),7MA2&bA3U88ACPV@=
;_5(D:DYYMfVO+DbfJd?[14T?_\_:>c+=Z=@I>X;+OBJ:NKN50DXSPM>f#fTNCHC
9H&P;NJN/(#R3FB(OV.2<:8S&<C8\eF.TKEJaeL5.P(PH09gKbcS49@2WSJ6e3UM
e-[@G?\_GAB#GEcAS)aE@<LgLI1P66aFTX6E)da:9O]f+?.VLUc&2-gJZU_F9ecU
^,3[&06Ac9R+BQaX;g>\M9IQM2IEJ<3Z>E:=Se(.+Ya9?aQIZB,fIPB:/(R)d3d[
FaS9^MN;18FH>@GGZ1W[b02)<&M>4FVcRPZ^#/Ga^/0IeMTX5g86Ma[/T+E+>3CU
TGgJQ1^\gFC#JT<K6PR</;;CX.^MWa&F8T?d82Ca.YJUNDc9f@c_CYg4M2]b7\e\
4_P90]IdbQH12d/NKF(-)5:PY>^DQ2D7(4c@H]22F26]QC72NBbb8Z]VHG@WcZ_,
CAY+V1?S+:LE6\WE7K()f8W(J7+218X)bIBNR28?(K#:=QG#LWPKEJ>fZLfbcW^L
&>2TgZ0DA)#JBH@g#1#DB1?5JK2aL8H\d18,dCd<9<(ObaC0]8RL1eR-UD=MJ(H0
3fKDNN737I=#(4\QLY#5BOK_57]cI_:8AZ41f+/5#^gB4^E^869K#]](\e@(1QK2
PTC4W9R/2U4(d5&ObT][JU^M8L?N)EJXIJ_+[LfG-I31S]/J/2THCdQA/WY@\J<R
0@)K+9RJ3+ZA;-c\ER.B]M.aVSDUZe#7(>6ZP4&5VcfK(5RbfR7@>@cZQJ;dAZ=W
0aFZHR(+TfMN[)gDa\9eT^<dTe4:1ID,K&J>_A5<[Y13a\Z0a(F1gLc-dLTHT:+P
7R@3+cWF5.EaV\W>OY:Xb?+EUO-YA(OQZ[MQX:R(724,+HN0CL;,H?X^R?KWK\<1
,1?.C25XA/:X96(?#M]GP0CY5274a:@d6B<?B232F=Z][4>fe5\OF^4VF0f:__4a
B4R>?G756=MW-V?[GbZUOV;_8NW><Ze4JMV8UPZ)W71U-GgC3Q-E_gXE+IOX+)1V
HGb^D^YP>8@,&a\A.GA(8@&5AB)YSCF+fcbRXL:]U(bPGL=329]PB/D,b?=F]fIR
g7Y:g=5/Fc6OXRG=GJC0@7+,c5D8;KW=PEE62GMACB.eg\R9@RcPO]_SJU7S;_bg
Z@K<=H:W]2603cBFG1UA3bO>?K[X3[&O+b9CI4H).0)C6b4:Z_@8R\0JZ?_?>\[C
(RfMD,\M3Ya1IX4?RJU0VB0JW#/_N3J^.HOMM(LU2#@>&7-1[GU0>UMR@UDB-+=(
B6-7YA.LdYKg:F=RK)[:RAR2YLJ#Y-:M<^^\-N#JZX5T/f332FRL;BK4M\?gM?A2
3L=73U)HSLWX>M+K43I4Z)3ffLUF,ace&.@(P>KW8HO3&3ZHM#/)B3EXJZ9daG>3
-Yb:X?G1E-JC[3PRdD5<M&?B&H_4&9H\62c585&L;#B;@]6N&D1_@[,S&TXNUC#Z
^e6CV2)P9^ZU/TBF9aTfN5ceJ5bHI1)S0V8gD)aJ432YG?>/g(UVR.F1<;T\3V?)
eY78>J?@a1D:<&H<ea(DE7I5Q>gOR)R^cJL6/[<=YA3.75e9PS&c+A\J)O#FP54J
bLKSgZBX-gPCc#VQH_6.7-N@b:J5M0S[]+<VV=X^;g]YN=?[-ZUgX&WE6S^d)KL0
U:^fQ8FK.Zg,=ef1H=^25,E#V<c9Z7WYTI@\C2NaHYaP)Cc_Q2<7QQc[M:E_:F>9
IGWdN5Dc0[;&BF^fa1<<SV5H4Ff64<635.;YXG;C0V]b-/eJ.e+cWff(&cG(c/gM
>Y8-@3Q8J[<7V?2M[U96\@9>@I,,DO?O3Z^GAAR?2EB@,bBFa&]QZA:&XG6(92c.
WKL3L5Zd)JW?4A8M/T.@4+:\g2dY?[&_GLQD5#IKHQQSRJ:XKR)39N^,UW;:?#>-
&f4Eg\PPJKQL>3]TgMY.FH+AC6DSLH7Tf8T;H.QDMYHC?FS_SLBXIE=EZZE7d<gM
aNZZH;\bK@SY,(-UY[7c&W4f4BM)=D;bMdYI0;RFOQ#NCSW@LQU]+&CEGR@8N#G.
>^FGLN^f4?-0NG^OXbU4H(_I^:C#OSUN9&1EKT=Vc#/_eg]VY)CHcM?A&5IM:B&L
>W&/@.VF]OE[,eCfCe?/J);TdF\E5T-JF_&^43G-5edRXSeD6T,Ac\RQYY).SLD&
\SW<)BHF3=e8Sd4Y_@=[BV.6[TYd@/ea[5M3U#4e\0.PF[D_,?).2G8b\0JI\.1C
O4HI1]MUQ0BMOF]F1[<VV.Oe^6+e96=P=83T\;PcO1M+L&.CHN00MTS:EK;COC:N
B9EXMZX,Q,fD)8U1>:McQ=]-=,dKg[.+/N+=63aD9aV+8(&A=7-3dP;e>54N2=NC
cS-LKA#+\BQ.Tc;g.]Z60OM(-];I+6?/[^JdW[L>eY\fg:0KVAW45U#7K4M(773_
T6NP8NX2/DXS1bMIA9E26><&K(5CF5#@LJ#AB<fMT.dL;@/dH^@=L8>Q^.GL2=7^
ceX93X2\POV9U:aE<P(GT<UJc2b.479ARH>6VfNaF.Q[,Xg56f0YV>TVU,Ad\3?>
[W,55O[5FDO9NMEKRR2dIMdJ8_P)GC2K57,.g(6Ng>B]3[@./NY=(cV_;=+Y),]L
PdM;?MNPZ-1UQ7I9,4N)88XO_4.IUS>dK52H+&9>>G;c=c(P<0LC.PaK02;KC;8]
0+LL??gG[P0:df)CBW86O)_JBAZSV#6EN>Y6g7N&HM^=GXU?06ET87NLAA(G:B@+
,_X?EFd4H.4XB?MBCRMIZ-5fQT():/0/C-DZGc1A,&2HJD^bG:=5Z?Q)#E=QQ#a_
5U&?PCRPU1Q[Wfc0g>-L6;)4=\GW2/\fId46eI9B>I<e)@JPd^^976QK<]2:dXgE
3&NT\QcY?3gC9fJ-b46639+.G8SNI2GQN@^G([+QX&G=fgOf&V61eRV_A>1\OBe@
NY^WV5&A-U.V#<X5LWZ.G&@:K)UZcS;CL:FcHe89g@gWI5BIgHC);4]X9QaV/dWT
/7gbg4F]RgCV0@eYIZCR>]-NK#9V&UBWFWBC@6;6O6;ZaNDH<RR8&J]GgN.GPD]N
NH]&dY^cc&f(VZXB9O\QL?NceTR9d07&cA2\84;,e1;\_93_7RQ#/MSFY@^\,S+A
;965C)Z5T@J@FXY-c0EdO6Dac(RBA/8+,:K.8XW6QR.@__40Y189XOY2\34_FfS)
56OPQ,@;4FCU7YOO79e542YaE6dR\bA@L.K41Sb_\13@X)fJ687>>b;9,5A,cDCC
QaU8-M4[&.d7gO234JeHXI;<Z:WKZ)bVD.+b?aPIZ<@&3\b;+U=+JcUFQc=d49CW
_0[dXcM/J;F+)@@?eMZ)=;[(7UUS@65S@KF<T_[?7450X;3IO740.)IdSc,:b..2
-;V]DKYV=+RfJ\,:T(a#9^]-.a&>8#@PD@a<,O#Jg:#]2T4[AfJB:e;VJ0W[6W^D
1Y?XT3X&&H1R&W-DeaJU4^2?H)\fB^)Y5#6(Y_RTYMaXI,)g=,<F2GZ_LfVOf\fK
:V#-a1gG0C,W4)LeN(K8gRSB,8.KG3b-I:K,Y>5c&W+F##4EJ8\NIZ+,Te<V<Eb?
[B;H,V(AIUQ^aSc;[gf.W;Y2SBg_g8P(9R&F4caLH#D<@^1)NP58eaDD_X1=GQ9M
;V02OY-Fb1+Z[3O/NOXZIaYcf1SMI9[[,4PV?\J\L,M)V9<+S4?9eD<+NATWMa&S
:4\aWZA\7UZHH8&J[Z?LM0M_B.C1+[)@-^_(GW)LJ^8KK11d<T+F.O)=944[=WK;
_M_.c(DQV7Q<@[:3+@A^b?-,78/NWQGa:4;VGfD9KD9JZF7(3)V4d?5NTg\N3d&@
571QVVJK<](#D#UgRF9#>#^\b@gRVKdg0fVBW[JB6ZXJ3;a^^g(eNOR\TaGf(#F#
3.313&R?GDW,.]EI+XS\&A2a>_BRH_XcCTPOQS=G4C1.6V+CcB>/#\JQc3E6./5#
[IDOUfJ16^5d6(4TdbL)5?=cQ6=eHE1D@\d6=BO+DU]EW>&K:eLW3KIF&,H:FIQ+
f@&&#4dL)057CS;D7,FI/Td2]\J_JFF\6gVJ>=4a&NN5DfN)+X.0P_,A:_3P/J1T
Y]=d7L60cJ0+[c5:]\5<14^&@14FL&=O8\I8Z[9,06C,3\@0G29OF,C1^S=)5DOQ
B\8.J35TV(4^H#ISZJT<MW15\//&Zd04JC+AV?/g#(>dZO82g6MH]d5A\?9EgFd\
1e2RXN2+cfIdV[cO5M,=]4Wg8\T0+6=\?DfG-G6ZA,UJ)P#[<+8b):8a5&bDE,N9
#K,UWcaF#?;RBQ2K3_F/Yb11B6Yg7[+<5e(T7b5f=11V>#=GF[JU&d>QGI[gHM)R
[52AH]f5aQAF([RE[5cVS2KQcE770.0PGAZ@=VA:1?63/EaKa/&ZfKZEgU=-7\PR
=g=<]Y0)M4RH<bG)2Cb(:d7YKJ<Y^KZ/)\0)V(GKBdHcbf,BaW2<Wa@61)Pb(]CJ
QHS1]3b/D\XUE4HE,>J=:.,V8X59U6C4O;TC7dF[/K+gUUWS1bIY.cfKP\X;4gO+
FaSe_4GVFZU+If)6N;M6g-[^IZ]4YbEUZ:_9KQXHW^6d,;a?Ea2135PWSgd_T:;N
<-N<26g>_90NMH=?X+Fc;.Ta))L+ZFEECBV]+OcV@7BJI@6?DZF2=ggGg7#B,fGH
dH7;5P3Pg4e#/=?4D?)XfWdCMO8-BBBENJ,38W2OUJD5\P7)MV/GY)Fg[2BOR+WQ
eG2H#+Z;=9L7<Vg8VdCWDBAZ?>_9PJVW_BQ_92,TOJ/0<_X)<;b^[eIeg503UUP1
2MELM@b,8VQ\G3VCWgXB1PKeO2AJ<a\)?A8W2]F,c^5fG64aYUGGWY<_4=B;Q)(9
_4KM0fJ2P:U>T-.D#bI40^6db-FZZFW4+#=gK9/=<Y=98=G:J1<,Cd\aDQ;L^dT_
CPebTDS4DMN]M=A7bF(?@OA[^ZGXCG2DT),\O<)U,K1&bb]VHacR+J^:f]ZV^33F
HK,SZ5WO[Ue_g9P@c8<Ff80W^N7>1FR/85QPF1a;;XF:,^Ja#SXKgQN\OJ1N9=.5
ZKVOIcO-LaZLU5T6^3DPK;fGVA1OZdV\IF0]dCLaNA;UbT]f8&STaFLL#DDIGIOL
F4W9:R92Kd^+fV)cG4V9KXC>HU@aK#6047c_Jb_(1T-WU81ec\aX/caUWe8W97XE
1BCJ.I).Y=TM/DFUYF78dMN.FU;P<:V?)4FU\BdLR\??fHFW+ABdd3<4X0ceR&[d
[60]dU@]FR&,V9aMX_ZL2\;+]OKfeg.W;\McC6]g22;FfKd##K2c\GER1JY)M,W0
]Q<N6f@F/PJ[DbL6HQYCRg9:>:_[]df47Gga-2KKa>M507fEV76[CIfFKT-E&9JY
.UF0=#A9ENX1&-/=-21E>b/.RK&dRH^U/.]I#.M/R7X.0XdIcfD0^P2f3&58>50]
:)YCK>LBCQ]:WQKK0126,d<D//UQ=+T5S1/8b/B\gN&K(?ZLQ]5/(S4K#WfDXP4R
T?@/KH<,=UgPW/P5VF#77&9R^,NC&6IX^RbdSA3IDC?RBS?\1;;4S]\KL(&6+BE=
I9H<If\#]POG-eBP-=D#PVXN^bTX[M(Se4b(F=aLaZW:M9:5,@;Za>DS?@)7T^gI
^Z\bPZ(eL)FHXYE4DfGSGc=P=IefML+abB3A60T(T@cFGS_GD6WMg>/#UGN[DfNb
3R?ba8aJb4C:FHAQSF120YM/GS,11Z,7J58)D>##DV+LgV?;P<[=JJ6\]WO5V:\[
GfEbLW3#Zf6+f_O)\9^(OfH7HS23f)5^ZMNTgO?Mg.[G8<EG=[d0_PS\WF?-15A<
J)1?=?@,f2^cSRf<=Y2IE4_Q7d\E?\/M3fgCL3SUC1QGE$
`endprotected
 
`protected
;?HKP\+/&\GYWK]C_<W#1NU.FIN9gYEZ&A#bA+_[9EJSd:eJ@>O@/)\cMH0S6AU@
=GJB)29_[5GO<4FbWQ3cD[(8D@Y>IfbB^cF+?f&V)<BbOEH0^WaSWG4<OBP^]_=I
X.WN[RPWVL19?AJJ1A[EQ,M&<LJXEX.=.13g<E=b-P?3E0WFT]PZ5E[[[@>XD_:8
NQOeCAEMcBO+W_SOC+<?K1F<@;(C]X4K+0AEDIA[3bIFYNdW2=\ULZ;,KMF(Q)98
g=UO5.4[L.?UTaN/N#eCUcA?S&R(4^B,X];Y\]aaegH];c3=H\Gc1Yg>OE?M7:6E
P&1YGVCa\b\T[C26C>E^ER=e_+B-,W598&WZAe3#L@]6>1.>LO@(UP\gR/:_,NVD
_7?(X,a6GQ3@-&P]\=.4DI)#L#(0F#.&Q]R?-L@/(V:N@M0A=+6f/((&86:M,L3;
,X/_He#/F2;S4e+GE/X2#/5UDIES[-8,YO78I.TNDRg3]GE0IS9<e[)O6:f+bcVR
E/=J(;B=SXYPVGL1;WbePe5U1$
`endprotected
      
//vcs_lic_vip_  protect
  `protected
SbE,2c75Fc+;SBB2-6_Mf;7G_OLX[URK^Q2S^;J@CT.-RP;2P+c\&)N=RJZ4S/.C
<DdHI^5N#27Fe59(MF+,0F]K&Mg^b?d_4d[R8K8NM5035?IWV(M=>CX_0O<VJe_C
1QcS:B7+.LBL)INR+c:PESY<U4]_\YI:[<UM<-97Nc&RZ)=K983\/PL/2HH-Rd]B
QgF_\_4T8KMb0Md82(>GYDDCL<@,dB[eD)G0H6LX.W^A2/7:TJ;/N:_R2VI#0@[W
0=-2NH11#Z0WX+b.425/KbRL_]]WgEdLf-X)GF#.W7^c7YEZ[-dVOX\bP?U6?Scf
6Z5HPS7@=-L-dbR?Gf#/C:YPJ#@]1HR6K5[0^Z=]]BH8^,8_MFPBM,EG\FTTPHC,
&SKPQ=DT^9[Z)>.NGZ?PDXKZgOOAQKJfZ8?XOH]Q\@Sc6RCE(&V)]CJ?,2\>_^;K
F@K@^a8D#6-PO,4XALF&E6.5]A)H5A253O=K+cG&<5VZ#2#e9QSac4E@^2HU,eVU
AG1)CINB@2_>(&915:U.B^;]#XK8S08O^Y[5[WR;g7.TNTNa:LX+R=<YUNDXZ7<R
F3:e]->770Ed^4MT)1L7G\ZO3S3bU]^M__.ZZM[N4E:P1>\C9H9W_VT?JH3H4(8b
f\I0g0K#))?16]b>c?>d]GRG.83]DTXQ4APaV6RSAaM#IGK.e[AUD\MG(\1P/-Y)
?HbMX<<c^de(NZ^-.+)G-+b7fQT;aNY59f0dc2JO_.cVVYJ8b8W;=8SI@WTf#.C]
NG.Y-2c[K/P6671PC:gQ\bK1LO[B#PZ@]g]V\N[,\4:<@Q-9g?DFV-TG)8FB@H,4
f1OK^;ERb5@TV3.O@@&4A]X+WUF6M\c4C&Q9?aI-2/eRE4BZFF>IgKM(OB\e@JLQ
.L>:J>>X;M]O\>2T6/FJYU7-DY)ZVdX@^GKKON.W.JZ^6\4W\P@-SLF]_#3R.c84
^3G(2]K\FV\fF./=VMJMHT0E=([&?Z^7d#WT0Q9W_/\BSN;4)8d:dBe>EOOdGPcN
d]./(:I#TE7]IMK&H75Z^;M/BI?;3RCK6Bd&UP&#O\6B1[J^T<e7f8V9W/I]=7YS
?M)eUJJ>:]32>5@R6a1S9;,Y83B@MWLaHFPe@F2eg)f/,(cTeg;^P2U--C?=Db,9
;4\8IeK2B4:696bg38fIAT-QJKVCF9OBI0QVfK+K9;5+Ac\[K#F1g([P^M_+,V8?
Ead\>D>Q165(O?<=2:S6c+>\BHE1UXPg\XR#43&>UgI.-bH+1AeaYEbMD)?5LHOP
&?Z]TSBQJ,7+GG<#5bIB<UA>LK+E;SSEO1C3dAb?27EW>JG3G(^eaQ\BR8D^4>GF
^0#C^,.;NF\NVI?M84R^0_C>OCgc>YgZa.&R@CaL/3A.<ET6G>KL9^SINbEVHNG+
?HC8&:RYYQ[T>R,A^JK3Weg)NSX0CTHd],HV-F&J3XA;_a:c\:TLJbae.BfI:4UP
3b2#]=Zf1.Gf-g&I_/F^JB<E^89)XL:[Q=>M7NP0OcXW/,_IPR66<aVb=(#HCWN^
/G6\9GQ9c4V,-Q)<WL&[FZCU46ZKSc]CHD/1]If^bXaP?I]&)YR5.1>E^BGT[<LL
6@U5T^Y=GT(@U>=fcd8I-M?8P?XC[If61[AY#<fJ?DJLP4)1cZ][)@TO\WBL9cA-
LGC:&38RUReE8>d(Z(WC26CUT=YJQ#OVF^CAFK4JX:Wc<eGS#K6<H(4ZI;JAUANO
[/RcWQ/2#=9IBbQ5CFQ?T]\\>(Q64;G&2601NBKO_YG#NSUL_6NRT#SW4,8,_GgH
g2F94_+0,5CDQPXU_a)+OX28F2=NNRX#1=6NDI+VQJ2CgW^MW^ZeNC#:G;CDJSF#
RJ1.bccH^+N5WJ2e<J\&4bF\O6Pf;D61CJ+:>Q;EK85J:S\OY>7>:VAJ-&U9U&dI
J-g,6/UB=9F2=B-7@:\^)U-^^I70;V,fZ-IW4W4cE6BRdO)F>2<I2GF=EDe^/X-0
/2].,:gc&0)-4)\OE<#Nb+cGCO:;+ebPUf7#?GZ6>M1>4RZ[@X,VX9;QYVC>/\:O
g972T3D,J=fHDELA?)IKP[,K14V<gg;892AOT)a@(f1Ia3D10g&f23Z7Y:;^A\ZQ
A8+1#V=LD,QL#_,Hb7)FNG]H4>062\<edUJd^aU<(])5ICQ,RCPbY5d?K>2P#9.E
G]5cHG;Nf9I-:?Y&)Y>UKBBX7T,#JJ5,^0\gDHO(Q-<Y>44&(1^LZ4P[Va_<fPI1
1d0_A)HHfG^3GL^PKKWZAWa4OBBJ=^:EA\H?g0c1B>)-U,S]DC=&<QdL@=;bdL_,
?I;9?H7MO(-]_=EOAHLA1=H;bP)918RSeP+@^.(ES#/-[-[gB<O-CN9NW^^@HHX4
BfK0U:7\5QC,Y8QYYE#1?(MO^RT6,DT[Zf<\A2fW&4g43c:KGC4C(^&9cENgNaCN
W85a5A3CdM<A)7A#d7-&7S&G/LZ>(8O4UcBYD-TNeM3(C@(6=G3fJZDTS)I&K((2
X5==9)1HTFPdRGQR)Bc+U\aNV\G\5D[-:?1^9H5>HGV72f:.(OV.IeP(L=DI0aKJ
?000LQ.H0?Ic9@(ZGc]C8+&\]O6/8-.CCaG4###R?b_N5)1I+0+e?](QZLLe#MKC
M&I1X,0P34?;R?,EgDAcd,>e\R/CKXQ5f?)aPPVa4_CD,GA52;+_bBZS,96bED9>
X(Og)I,1=T&TL^N8F_;M-H</:F2ca.g//+c:gdS8C\e=&2PJaaQ<Gc9L/_993#FC
DfMZgd:\=DVM.eA&A.+[[Q@DCY2RCWUMT[e+0AH,]ZWZKPGe]>M]B7[UCeC:)b3>
ANf[U4V=W45bH<4]f)XJ:DJ7PEWF66>e_&EU\;)=7ZLYFTX80C?>+_&)O-/I)&(7
V-V/Z<J:MaB\X]UQ]&R40J&/bDCeQ#M>W6<?.IaJTS-Hb<S?<:)>3M2V#50a4BYW
E9QeYKVIWS#;&+9VP&Da9S3]gg_eV<QXAW\[?R36DbXd?QH[KSC)74IaINDE^++,
Nac48JJ(F(2]fMgUHG+bI\:]]?@BBbLMYeDS]8RD;431MTg]#_B/[>P-3-OB^ZX[
P]cC[KZ&/,BQ/G(Ddg^EWL)g5=7a@ZM8)1+2SeK?;[dQGT/T:76S3VYQM-UYB>)#
X,XdOa3PbFC&]5g(d7JF)Zba4dZV@,@0VK67]B@?^,@?Q1agBG+]gBNd13GWe-Tf
WTQL)YVab;fB28<_2C<_XB-8/R=LBKWU?0E#eYM<7U6J0K^.<O+-_F7/\2&RWKX=
8LHKJ4f1\a(]eDDfO:0U42_>,dT\<VbQQP0eJ-;D?7A.HT:9WOZ)1[U?^3eHbEP]
CO#AJYN1-T7_g/?>2HVK=+8U<YR7Z3:(<?ME&P<@UM:,H)W,_7-7G&=S66@S,La1
K<X445L9dLJPX/V>7c^T:6)V.?R,UY0Y>+A-e)N9]FG;0I9]_a,Pe]ZecOd9#[(7
1-3f#-9S,3@LKDWCd+AY1(d=b67fXRHNIE,(,_LV/Ib:/8[5:1RG7Y)?^e(L4Ta4
5f6U\88T+:CLI)FaEPLL4;ZWN<18=IA#2)TE-Wa\T>^HO.B+4DI>/=MI5.fK((<.
P&1U4OS:50CPP6+A_NWTC]A.>30SLABHB1W@&c5++R5_#^ZGA.OcFTG[5^H570Rb
&O5f+&YNf5SOeGVeAeLcN]N8AT450,[MdJRZg^-/8c&;aQ=A><POPO^:B@]E:<0?
847WTdME@WeZ=4&U=Z/fZ)-eN:SVfF<ef><;LVLg6(LAIWPIbJ>MH,^F(LMHgE/.
^Aa7OVUEC+MTE-BUZ1/6R#^dD]&H]-9gLAJ:UW@,,fL[KVYC@NY)OOI4M945\aNe
^ae]-RCB\R0FK#659UOL(7[9,L:;=[6EgAF<73?Ubd7UGc1[a;S_T_?e::8M]2Y;
14_40R;;ZS4M3->3:;76RQ<(g8c+MR:ZMJQ1V094\C?>,].-_aKEbdfMU574<]XE
;_<&7CdD+:WgfON?4DMS@/\X?HSWN^T2Q<?D++E#/d@LH+CGKTMZKQ.=#0H,YPIF
/4V1T>_7&U5<1PZd(1Z@8Ig]9@Q#HD7T;7F7ffcGDa&HPY4V.gUN,G];]0=HZO>.
5:^fA/T=#eC.@a4&/TU+@e?OTY-)b>55-:RL3I0/GP#O&LG1Md0Af4<1/-RV&ed-
)(\R(K^]3K)2JUTVU9=KS(U76_c+A87dBGL-M,:B7/WUO2,YbK9P9-?6e.I.^LUC
I<X;7D/c1cF^[5G^Ba+M>Hf)3X.&TJD.?F.:QVIZF3R)8b&Q=X^FECP?_L:58B0L
2Ygde+N>?.5\#TQe4&fdQe(FJQO784<e.ga_6-3U7=AA]T(HaOZVb#+B_a6^FY;V
>Rcf[b3]Eg>R<N<:(IY[60g:W2C)KRR<XW:)FE)fP9a;.)M&9Oa0E?]QGN4QD\_a
14B,(cSKNSE5W[4a4Z@=M&;<SX=BLKc;BEN7KZHM95FBUg;PEbN5U>MM2?9MUH/X
6+)C2W0.+F+CK;_?S_7aFdbL7)4BZ8Y7/[Vc_a[0W:\]CeK7F<8K?M>@B9R-E>1J
Eb36@BA&3#ILcRKIUBg=?d6R)A@bPQ^L^^^T:#.0G]9FUPK+<KG/VQ)9+1g;F)EY
4efWF(LY2NR=9@aY8_S.[,&:+NGSWgL8)b9)P;523^D-eTM<>_J&Xc]AO&PZUZ3L
-WUe9:H?SR3KQC/agL3@KW.cHQ/WYLT-YgPN@9-.1LD0Y;Wa,W6SYT)ed:-eNU-7
\W7O?WRY,2A:<CF[3<?2#D]a=]IF21MIUQ6FG2eFS_Uf+@?_27//C2\g7C75BZc<
YAZ:-+[07FA18fJ6;\:9e0GeO5-67)ZJ.<C[?V+>cLd_>=2PI#&[?3LYI_/)0,2V
eRVV392++G7BDDf>4dR(9CQVZU0b9]?-]ec7H260Z9g@)9PDV(HFcGC8Z>1_;LU0
YAdeg3I2\]a^BPM(G&#E?Y?3D^94FYKZ8GMe3PK=GF(aHbg2O4VVdPO-b2M057U.
K=DH0dc7DGf\ZQbQ?KLML::a[OR#4A?84VLgcTC1fe(&?UJA.Y&R3:NX\\=:<JBX
Be.Q-R#1-.SJ-Rd-&L4?^5C/_f9;fD?=UN+21<7?7]C6\D@<gA<]7ddQ0ggH,\J7
/<b985eb2@CY9BQSR2IMP.,5\D,BM8695BA&e)&]CNTIg-W#,,)/6-D\Q1Nd@Z0-
97[]4>4HeJNf8<(Q@a(G<WAD(0X_IP2;O:30bc82b1J^;bERe^@,:=[aCaa3dS&+
P.BTA:B>e.8&_4^R8TID-2EK.aJ.&A\gB+L0^41c[JQF-a>HSJ>,4-+KV0WVbG)=
&/N3XAW#TZGHB?(eX)5?IC-bd.4G(DbCb/bd\6P]NDTIP#X#SRgA:=&S6SV,1YC@
>XZZX1DHNc;M,OZ>LTFRK,ACDeaeT+G:3g&dL4)7A7+SBD0>&?U847[,;cB=4+<2
ITIc\5cfP]\2daJ\X67b(eE/4^N;P,70TY:?UYcBD5/[F:@eRQ7+Pa3=<46gXZg0
YTT)g=gI3Z[Z\WZ.;YSB8P&-96HXE82W82bO9L9N]JSR<a5&M?S6H7OaGRMLgCR-
4DWd.89D:H4:?/BaJCe0\c=@&R^>@6W^BBM6:?]f>A,9I:HeLQTW>,1#,^519>(,
EXU/0-YU^(cA>&3;F6BA;#7L\VeXB[)(&1)JQabTdcN^KOaN>Y;#B.3#3GQE]dFc
\BD&-(eD4eN[M&-+9QML+FYLA)9MC-MaI6X&BTU9d=WTUWHT]b&XF&^a@31WOHG@
3V<U\<4QS>GU2/F/[eLEJ\1[_ED2ZTE\b48T2f\>a13g_A-bR+&.1?U(a9AOfeE;
&/-?C>_^\Cde-AZG1OC<Rg+(af-+d&]_?OB>ScL,<>cY&ZH/??gRU-THIL+f\fTV
>0H=gDZ/Z5X&F>QPX8K-5(bI+g?-J<TP(DLD\,W+_7ALJ^6IQ8VfE+G<#S>,_C1Y
NUY-R:P93]?bI.Z<ee8LOA=C::TDTd\W<?a&LOJQ3S2QIXX+\.RF=Z@/O<\&#+MH
BO.CbA09F)X_H-XX15]K[V:<Z&e>//g+3P#]SE<@#e:/VM[JE\?fXOH:).,<d9bG
AO93V@F?E==Hf><O\TYL-/[b)3>E\e6H81=PH]CR^1EQL=f/4Xcc2-[HS^#=AU[F
c2;dW+fdHPJe9XACR&?0D0NbLM5Zb)MUWU(P]Ae7VN_U.+O>&L+/C6Kb1P>/P&JW
g^]L8efWDNANH.>bBcG-.2A)cU33Y<22N_eS91=)GHZS)2#99#9C,LZJ_A5JMY4g
+<KM]+1JW/@ANdfC&Y_M&O&@&b\1297]W^<LV0C/-Q6SUF6K?>XN],-2AST51<#[
(R=MQcRdC6)(AR1U6V-abP\:g_dODL_R[+/\@]VL[9(MDT+PJ-<KgV=W=K[ea;=1
FLFfg&fR.b,)^<&3W?@MRH]-9)2AE3b7VL)e;#EQ:&+(Sc_^JMQ_6Z/]H+QS7]KO
GMRX0Z.X10)XL>HC<G?cd7b[JFFX?\6WM_X+d&)6TAaa_A_TYgC+BUET)NFL2>&B
+C_U_QRP5E;ZP5/+TH#:E63=aK@KIcQN35NIOT3N^/]CKL#eKHG\Z4^b&PDP^_Qb
Z^D@_H8<<(9CM<_A?ZK9J6SOK/&Rc#+705Ab&Agf(_g&<CB[V38gW.4M#,cfYN&;
+/?L2@e2gJS]FeGN9@?1OHZ\T]bY]5+B\TAUf\)d_EU,bcS^T[=?L><Kb/BeOUX_
^a5I@=_Q7FN^NM\K/MDgH7T&bJIHN.S8[K(9L-SWY][:M(_a>FU76OQ93WK,C(YY
4=DRC,M#1F)fM32K:,>b]/^-8-97G52SL#T6HWOQ([3?YEc/Ne8?SD9@_^BP9?RF
Dd1_,)T5aIAE7M+77JTf>_L/)&[;cF;\aBWNbbY0J94;PEgLQD_>;BK_@Q@f,H]W
SX>2d(XL18fcSIP]e:,5E>/fUaSA+#JVL->9HfOOQ9YRa\-W)=OA80N)BdI<1_^L
C>T4D3BEW)#dCV_,KB,#g70HLOH)>=bU?2XV<MSW@3a#U;/E+ASL[_,BTgDQO\K^
Xd[<5143_M_PN2-e2c?CN5b/C<JW1G>ce>N>9BZ<KV^4/@&<3<P?OT[F5.(&[=N=
Y&8OZSf=).#AXb&.QGM/RU;-[eA-SO]P3^>^#8U@FR(U4;9#.H[EAdT8S#Q8AWd5
V+.&)C\16@],\-C,:(7gcZVRL5J=SKYA;>(_OSSPV(2<9KWJQMH4S32TQ6KRSWc.
VYaIGV5=<F7/G^MF@Zf./Z<>/Q\5PM+2#Y86b2Y3&G=-XcZ,C^)(-D^E);Od@<.(
T1^TD917YF\EZfM37RACf?&[)G.-+0S-6Ne\._]N&[SD3(b]MXJC\997T:WTQ#()
B<^afKCN4&7g3GN-PSJ1=L)(Z#F_X4QgBdXZ6AP(8:NS#Q6JW:H.g72@LO5BV7O0
ZcC1C14ZgZ@#PWJ.FJ8U5.\W?[Df2=1[Pc.UBM8\DHH0(N_F4dXK6fdeUA=Qe:2Q
)d1)E/=Tbb]T=83cM9:XDf>0:+7/\^7P)P^E]0:S>DXAQ?aSJcXZI#]X,P^T40Vd
#P5@V2HUWaK.0,<Tg1X>#8#59g3M7/3@6<6&>O?3.6dZDgFYH5ZJM0f^@QC_UCeU
)3F9=>0_>J_WQ0M3-dE5@NP<:-Y\F,T<]OO/T<_GPL2_^#<H2a[EN@V55ePF391O
.R6VRK.cfQ[:2@V/LM8?Z:GB8+cADC^FQQG.I?)DL(TNJT(YI_+G=S(.GRTRS?5U
0Ld63-/6QDg)5;,5KVfJXV&d^C)&W+F++D017;,5^cdPATe1V/88c+#RJ4\;=(76
Kc7g>M4bJcNATWJ9>JJLEH/c=]^68e\M()8#dP_f4&/_VYJS[.PePN=EI];4][F@
->32MEd7NTd8Uf1QK(=5BRO^MZ44?O^5#U:<?+ZWAERIWf;/M#c;3^)4N10JWTII
PXTRF6[=AT:H.I>G/.H.OF#QadLY38bV6T3[]?;:I;XCBJ)N4D)46/8cO;5P=2A?
7S8_.V^^9AeBWXd>X2QR346M/Db9W.;XHOT(\]&8N;YAE3AF+Lf^SVDZS#XB0e?H
E(@Fb^0(DbF+Ma(YPJdKP0J9V\<XBfX9ITeYf#:))5ba1Q0Zgc=IT@D#:K1+510L
L5S&+GZ>-f-d]ZJEJ82L/,R=[ILOQ=72X?DgLT7)Z/Ud5P78)P0a.]):62JU4U&C
cFL?d>HOHKa]KUdG0HU>ADG>=[Q0VOMS)&/J/ZK]R?Q<88<cA\4>3>.1.Ka(V2d#
d<)S,dI2VJOLQ:]P#FW@U=(,Q]5K4+6>?+SdD#3,44ZRg/.M;F4EH48]@=R&U#YF
ggAD,H_^>_(.O-4Ma5Y\8b7P<V6ID/1(CATd6CU]MRfeG14XaEPY-L=Y61I?UA9&
V<M1d)8LbAb([]GYA^E;9W\RLIP(RL>N3J04ZFbE=4O6A=1182]Q(4;:FI?]VAe;
1V>FBIUPd=.[Z>DC#=3C=9V4=+P1IK62UZfE+PCPTd<3@2VDHSVS(d>S=_W1,I81
S@07fUE&\>Re]NBdagQfE2CNL&bF)^Oa+].^Qb>E=T?b.8)5A?3;&eYT,E+.;I0=
N]L2D\8JEL2UMSZWRaZ)\=<WNCb:,.+/]LSg=XU[F[&>AW]HD6Df.G-gP]W8adRF
2CZKS<4&4\=\#8[=;d&D.NT17&8S/J+e#cVX@8B2Qgd+F#9V]UQE4-SL]+#(6#W=
_>(+_,P3aI:2IK7/#ICZg>4\?EYR(]GB5gKS;(J,FIBTgWXa]1#-PDK@[PaO9ZRX
9J[6SB=5#H3&0>+Sg<9I_c3d@]4N=7^:I7e1Y.?KZ-^(d@PUTOEOKfVOB^/9Q?@-
3=W3;+;DdT,Kc?2[7]/-&d^&\ML/e3WQfdGM,8QQ)3/FS)/<Y8^1(RP>NE-0&>dM
>TbJ5M49gU6-IK1XI-_VV4d6W;.7)^?)=-)Y+P?Ag65E^R\)B@II+BX_5@gRE4LH
,S6DMK&0b;ad5@R\U72[J<LVDea0S_YYHVT=TNBUMSH+[I11V(8Pfc@;f/QP7^O-
I-93+12^\G221b;B0,KJWCX@+N\GWE+OO?a5T;;14O?F+#Ta0bQH^a73HE@7<a67
P/K^.6QT&^J))5;()G,^^g],02W:LeFAM#;T>,PX20M[H5)ZM;S>LS9;JU@KJ;R-
H_0D0R61N(PM0K_MF<0]7)-B#,TH+7WC5a=7=:JX6MM,(ACf?3#fN\-f]BgZL^QG
0R.+cR82NZEV94f,].Y=>9Te0OM03aCQC;e)ea)I:\fD&=8/+KP]C.=gEDBZ7.9f
WH1>\48YTa@PK0:AWPcKW67?g)6f0V<6UIdecK3>>U6d>O4@#2183YUD>;MC=?L2
Hf<bKfAe_=Je)YFS5L[ECb\+DcDPD7X[7)FBQ:-Z3(OIb:1<DdcEe/CdVa,14TJU
_&VMB:YW;6LNYOQZfY<?9L+.5Kce11BY6KHJ>bTE/5+WWTT-8VW3gB<#<>Ra>^IN
SIG(3GP,?DQ(EdfZKRL)QX18N5NXRW2UR>d0Saf.Y+Q]:3)b(E&JF]V&a(SNE:)>
5/<OQ)G8-67_3[8[=;_(N_0HN67D0P6bYL[.OO^SdN96;XRQB?K[<F(eLE4[Xe&9
Cgg^#cEcVNV[4e?#[KO;IW/+_#:_?8SbRNIY+g#[OO<[AMTDR&5gQfP]NdfB5dCg
aK1NI-7TcIf6AZf?I46,B;?e_AD7Q)b=:)<1>H7^VQcHX67a/V69^W[[WRR^RWbf
8@f+;^b]eSA2@a#?JL5cH?F@WBF/MZLR-E54NP8_3GER+bMO\K2(SGEMf+=QfLLU
5#0&QY<O-FT8HbW?(,]]6Xdf#;;;MBB9D><1I:S2U6ZHZ@AW)67J-B2/>).[[&U1
/@\);GWYPHdD:SNA@X&17b3V\T&IN,L:GA^.af[PB7c5&B8e(d=Tg17?;.Ggad3g
O,6Vd6UZE=L8;V5B5HR7JG0AQ-f\;(\B[;=;XC8PYbX=]1N3:./W;<Gc1>#:7RYg
#\/P<.5?>/cBMSVbI8(KIKFPN\bSJQY^&AKgD6fH9#-cPI@#N_9-7>KPFM6C8U?U
WH<U+]/VSL@&QcQ/S(NaG51(^F0bUO0),4GY[aJD5LHUJS&)WOP^\RdK84CZO;?+
).2T=5Q@Uc^eA.eP.H\6&GFW@bKcCZ;ZXfB6UOG7P8(AKZ@4/>B#HD&18/_1<.XV
aZEQE209a@+Z3\[&CD.=6\RA>Y0FU02cOg0/S[<1H0>C2QXP-S2DJeO4.ebR:?g@
>8RS#QV=:H>SXQ2UdIK(:-&9\dTRcO,5]7gJ[W&REV;QQdIcFAI9)BUNV1J?DMF-
75LT.PaO8]N:I3(JW_4PH::KM;W<ZD>29Z+J:1/_-816adZ^f=2L@d>(MT&bVg_Z
a3fDUQ(T)M]6XU#7V@/N-#_3&/K;AP>+-Of^c4Z/?S_43.[A.X&:J\C:(Z5>f3fA
&NQII7@M<TA9QO_c8)0[8X;f-]751;70[AUdY6@T5)2FZDTM(.#50eL=0/@;1>bE
JL#EDE0VQdaIMVf2)Da2HO6S72:IZP@8LSFP.:6Z8]9V@3c^Q&a0@.<A\F9f_SEH
.2V_gEES;Dg\6HV\[2Y2B2XfVCWCGXAFBP;E,gRZe-UeCF:X2<;?[^[>[Gb_&eaf
cPOb2\DZC6+8Ebd<cc;:_>>0:\gc-L2NBLZfUZVB/;BA/gS][.9MJU5<7VAg@#W,
PG=V,e=_]FL#.H_AfI;T/Pe5Z/1@RF9Z@7JD9&B&.9Sf=I7dXBdL(g2.YOA6_X;R
WdAEbP3d#YAN3I>-MEDbQZ?)DYV,<Y,L_BJed.d>D^KQ>PK_>LP5JDH8E6C.__@\
&^JbV)#-O^73[R1-e?VVU_FJX5YdLGca?FLO+]QRI6Y[HV-G^LdB?#?>CX;Q4L;U
-5H(gQ)e,:03+FS;:&f3agZaCaEBUA(W:M^M+8;,0/D##?3W#cb@\69)O;SeL.S(
XF2_,[^/:UAON,ga2b(^3HdB>AHEQa-Q8?SIKACH>J.B5[?MQcf.<@XWd[SdX:(\
V:#6.W5CT?EfdK_4J8&>_;V&g?gE5B\R\FB5?:;W>[-a?&>F4XbLaDIBO/+dB+N/
d-D_E,#PdP.8<f]1^Hg([;]M?L]RHdMeU+aTGQ=(]Y?WOeWL/PB[fI<98BdVSX@[
U81g7(/8C3[Dd(1Rcg\\N-gIdc#d2/)0D.V=X4Hf7eIYO#7OB(T?BPO3MXFOG>Bb
#5B_\#:[(f9gM?\b9@^C.@_a<(4CXe6?I<Ue586U&-:#NE(N:-2<AWUP1<?f]W&d
6GR@O?MOPAMK4,\#a_(20+[#3],XHZ+<&#g066N]?>]V7@V8<V()(fX&:a0>MWU7
?;)(9V2f3V,WT&aG;?0^ODK6]KY6d[b#A#&N&XGX+D7eYCS8#fBU3EDUV9Qf<QJ6
d9>]WABF(eJ+cGWP,Pb1WR5@T3DKFFG5gNQIMN?gO4>4-S+\HI8cd(B&(RD#W<,F
0R.G>e9A&4U(S-]?5YSc\;,e@7>F7b7?eTJZ9fJ=c3Y4\R31MbG@;T)Z3,I:+>8b
b>J9fGRQ[G.9]aV_#1^\8&PZO92H0=@3#@N9<&<HAHU:-X-9;@ZCK>+,:M4CP(8f
d=K0_cFH[F>-11N>LD3=41;57b?bV;fQ/N/]L;^^\=0TPWA?D-B6WUG9W934ITO.
B49&N?7MNa@FN1I)#9bN=^1(V#8Y_3F=8dc-W_&K.aaa1b[R]^@2I]=9WR)(I(BM
A/<;/2KY/eJ:a,KTEeQGbRaTP70;.TH(0aX_&>4BAWV@XDOPN,;7F^\(39\f\T1X
GPO0/=gSCV0:FYP4NLMY(O#<)GM+H8PF-X\W8R\\N-OcaL?A=KdNH+68(f/3+3T^
0Xa0JD<(9:R<6EZ90?YF-3KU11DbCLZ)+00?83X&<>?K,F2D&0_][IZKJ43=Z#g4
TG0;[]=1Pa>ZGKUD)Z/&94&0f\e93BW<@E0&NPY?MVcg6@FW6R?VS+3&:,4DB3g@
Sa+PXP#N;;;=>M5TGQ&[baO_&P.,H+:.3c=@I9QXVf+I8[^UF9MCTAOUA45;699Y
63(CF.NN.UJ]U8aIgdX:IIbSMODOGVJJ-/,BM@ddQ7MB(CCU<6eBM.\2b5XUO,::
W-[?[@d7C\eaVZdaANf]P8F1+I<OHd#X&DVd-&?8Qg_3S6?.R@7FaL8JG->?8KE]
\PSDKV(VX:3GIY.XKZKMKHdG^8cIJ8B\^Dg+70-3Y>X+[.,//,D:F5CIc;A\HQCb
gU)DD,M+X.P?U^@UI8G_C2G9Ncf:bN)QRG<g11AYN]VRK(.G8DLBT-21g>J9&LaU
G(6^H+I=E=K&Be:Zg3;4Z\CZ:1FWEKH341R/9CE)\f<LaQ.NFGcg?RdTQS/>B;M0
K3[f<^[XK9g-Y3P7KB#(\g?31)K,MJNYeb/;(+BgE3E#F+<G-IV-:[D#D/IH5[^E
K+_>?OF/ADX?WNA-]9gQ@005RD>bRKJY1T;<N&8g52Z2)AV48S[]_e:F>5cM,A[N
RaMgDOa]0FJcQ+U4>5UGZ8WQFcVNIdaT?>C]P);bU&VT,c2S[ZU8UCdB+JB2dH1]
_;R/f2D&,;8.ZPg.&)F,W1=F?_>KcNM(DGC5P(Y7gK9Qf94Og,SRKZHbe5=38XPT
Q-)WS<_67EEg6;Y>VA@WSgBNBcN<Zg]G5?)f>[Na]^3f[J,]IV3G/[@bK/B;9FW#
ddMf,f3K6A8Z#a^RKSK#FCS1dO4de:YI\?TcW7,f?E-\D5;1bLXA)^=R4;aK+U:]
b.4G9[D;/\H>3f6+cO7W-QUKGS/?_2b.a?JO7VIacK<2Z910AUb>_QYA\?2E,5RM
/3;;+GE(&];:b5K])JWC;5(?g3?=A+BYFd35dCU&M:]TL[THNYP.)>.@6F\&34PS
+4#b\C>KZgY;T83aGY2dLO9P4O3d\[:8&.fce/ce&/U;^H>CCee2\V:^<(BU2Q>W
a,K[/M]P=X:bBg(e_IOCD-b\>;2>M[4\#5AN<<]XF08e]GTP-#AS8FM:,MXE/Q)V
+ODKO(<K1KJ2Ta,0EHSRE6ae0gdBFPX:f5(Z)L3eL?gC&#Y]X0[BgR^-QWBX=_T5
]b.<4@:X5DT-V_AM;GJS,]G:eB-=HZPH9$
`endprotected
                  
`protected
;4#S+4]R&A>Y0M>;+d&8/ISe@-X2B(1VA<SI9HZO3c<^Q@5K+c6A0)2/4L.1_\N[
5O-#cXJ]9UMcMY]KTS3P2g[C5JWgO>4>R>g;.(9P/P;90W?ZG))J[dO348D#Q0LE
R;76)(gG1=Z?_JX0FZ5/H?U;5BCG__FSHRND<BO97XOT4bf[?P-CYg1_J2Ic0I=W
cA#Z[R^6&gD@K2OD3\H(N;R#Sb0R6?=b;$
`endprotected
                  
//vcs_lic_vip_protect
  `protected
15_+T9SU[]L>01D0EX>G=+84ZXXY<I)d>OL)_VAO9I@gOIB18dU(/(\:,6KQcSN_
.HbDZZF8XdPT?<O7MfH]A.@eU+ZWVE?b^\BLHDB:Cg-(.ddE.K,?^\bIIWACE@M]
Z];SJ<(1]ETa0^DUVN,@RSf#_>Tg?#/+EY_b;CT7=D[LDV;;Y<]-^fTUfgNaX4PY
FB0DCDOD+<KL^5A5J^Ebf+)ZH17ZYR<U4cFK-X6JM?8H@B>K:MDTfI2=DY2>bXII
0K\f/M2@OA\dI6]I.)de,M[=g&/Y(eNR(W>D-RPJ\+FUc(M2+V-Z^+8[g:a2Cg-N
YHSBL)5?=AfIDV<Bg=DWU#ND0+I=/FKg/gFY/N5;^JA[VZ0_F3]IUV?(ND&Q\G+<
ZQ)_T<WCC&+ML#d8-<USI&ENf6gIWIW3=b2d/.?M4#58E3BcU@<O?LK0U@^c5RLY
\/52AaXA.9.^EB2JJ-fOVAC/Z13WNG?e)eF#YHL+G7#4EJ;U939?H\Q\A@]a^B7,
36PQ41U9T.WRK2:AN:,_dG5-IcZD/Z_<g_8B:LCO0.<_P:gG-7+a8-9\>XLBZFa[
S/.Y#=\58F-?;BfFE?aaY-bR-\MI1=9(f)<,?BS5?Q47_BY=\F_MA\FNcMd^WebD
&aF9WS4><CG4^MK7/X)HWaAWE>76bL,RU>@9W1c;0_C++[B2;X^\<F2#c6<_<4GK
Q1=L(60@S/f(B3J5JY+3:2N)#RIH^d&Mb@_Y4HggNe3?bS^CX+N?X39,L0Qbf\6P
1<L4Q)YD-L_3LC?2O->[>JT;(3OY,BR^F>PIIFF>L04aRa[a3PTOH(7fP75SD)(f
T9RB^J:_HHge8B7)fZT.Nb]DIb=H(VI]26)8b<2O.7f-L.8-T&.Xc)P.@R_&SG.g
;V#9/V,NNDTZ_?Vb&Nd-I(eV)7P[_@EK902IJIB5VJS]HK+eJ)(2GTUY=A84T?A\
E&V.W/3M<#.^e>7PU])Ec_=;0c8^BJ<Ve5O3bJ1LL4Q[8II2^94M+Y3)TZPO95M\
\86<U^bg=]eRdA048f@?W5RD+ZMcN[\/^?,Se@JEERZa\c6g.f\VeaV)0QA)e&cB
WT&^,SaCbaLQ+Q.0ZDB/U_&>D?eT/;1S]gQd._F8N9T00)@VSCE?>5:GAP&eZM?6
Gd7_9I^@V5S=PMHAYJ<>I+YMF;eB2:IRE:eK+OgN2ZIN(BN=6UOL@?d)g#1P00#Z
Z-6:X9_OE8W[:>9]>ZB3;<V3TDOA8GOW.3TOd#GISM61_K[3WaUa.f4=2XL&Y[DG
g558WCER9-(PNfJX5MZ:(>c;g8+4<<ac@\>:9E1E/G;G7N^0Id)PIE]Rc9VYCHe2
O:P#779L)I=/5IIb4R^/[gLM4@5OEdLJ__L6c3)YE6[K#EEAK#gM6FWTeN^F1>DO
D2WND2W1aC:YB2f;L7?.(N:BNABP?/RL[,Sc<:-W\_Y;d_e&>O=6d@2-Db+U6:5F
;Dg,bP+]L.-N>UY=Bd(@b9/NT9DHRc?Vdf\Ze,[QC>5a,9N?2e3<2_I>;+\2O(.>
UCM.@8^E@:&O:b21<D,c9/:IgfM:.3DV34F/>e]PS:&171&BPX@Z/[4I-G.)-NF+
#)(_3#)c8><S59Xe.NZY^0/<<.(&9cTE\023\bM),1/Q1&_?.8BW4&QbNOK6I<J4
A(^f)E[b0W.F^a]0DNH^:XI8G(;c7DZ,WN#47UI0=1MWU@f6ccFXMYUf+=ZO_5UW
J169>#cSMgDfDTfSfHQSRgaeN6,4C=0Ag#@J7:d@R4[VJA,</L567:XVS-\a?.@9
V+L6ZY(F-P&&NVa(4FE2SQOe7._N1I,F<+&(.6E)961BY#bJF,Rb/MKaa631L)Eb
_AcJ74F.E_AU&fTW7D)VR<>-caV-SM=eHNY-ZgT)0L[LI4b3TY@ISYL=V,&I.X,K
WgV)W.7VZTZ&E-XfA^<.R-[HW>@g2K.TE#TA=AMSg?QBEVG&\F4<d4P(F@-/+]]G
)ONH?-XdRT9@?];14dRWK?AG_0H7]CR:WOfaA2Za?RgGBGcc:+Q:,R,6RWbH1)=<
Xa\LDL&e3IZ<-\6a6+/H?HPW)-/d#R[UU1,)XS_BeJ2L)Rf:gcReS8;Y314R,[T9
<ec0a9[J5TgMWR\TQLM&SI/C4+fb/+4]/J+LV#3g+>8C^^LdEJ[R&Q+.4<(b&_5<
F<_OE\M]G0X4L]S;AW>DdW(\0g]bUePTZegHZdffc\e=:?G/<@4>Y&^Z9@GJV1L=
^/8^1eHB7D\IIUW>VPI_d:3+S7@@bada0_K/\+:Q]#@EVL+0MG8g=GTeAH2=6+E3
ZMHXP9,_BgQe?FV#?792#Df:FY]<7cT0:FK45AUGSB]LOT_N)A@5NW3[U-d))XRM
\,TeW#gM/#f9E<RRd#1Q<_(7(beI563-61RN[L7GEBcRKgd=/E?XM^6DNQ4E[2HW
1V>:VNVWO?V41e>FQP/FKdf[gZGDaafZ.2=G>I_Q5a-6=76#VPQ_9]6b;DVK;)(-
S3?ZLebKEBg]?IEb&4Q__>QJW?48GSYGVJG,bc63X,88.;D?<VFS7:KG<Z6,?_6#
A4Y>R(87OfgWO]PD5](3aOQ_d[6L^&Mc8WTZOX\G=QL4F<c&daBbRE?A^eKE5<GO
@Sbd/Lf#[&H-M[D1dVO;X5=WaWVJCWaQA17\/#VV\3/2HMT:ACfae\5f7B#<3A#?
N6UaO\2I?FcH9G\G?;6X+^Mf-4O]2O>,)UC#>gC)^L3aQ@F;+2_g=(9)B_7_04OI
FdP&S5FGK.&8GKV60=+#;^3\<SKfA\N\0K^MZ/+JS<+J]7G68:0)YDGV-]])I87H
&T9GW:4gc2[)GL^,fcPR[+Z>CbgRYRB1H(Y[#WQ@=]6J@\LJe[Zc:I2f35&YJ>b>
T44Q@J&TJ@Q??.+QN(+.0I(5XTD0gF4ACI:gZG/2M8_-KTPE@FXZ:[8L3&L\-H&4
0H:GN2dEeRN(=\P>?+II0?:\Ig:Wc,Lc1>IAOV[6G^)D-^0GL_7f004WGUZ.4g8,
R5RU)FT_JEDC/=:BgS4:F1(Ha]H<WK2&,MP-60/N;5J6d#?K-E/[,E_,S0EW94Ge
[A??#&O9&PYU7DLbN9e::b>Y]MA3FB#;HQ,/CO?2gW[_+SU](:^XE-b56>@@(AMN
=)=U\,1fIfK+gA.b-QIe\MK;WT=_eCPVR:[L4^?(JGEA&W\KLQg]0]C=<:2<gH6^
fZ+HOA4GY77#7O2^BYS&01fVV1O:\<W\[[RC^TA>/MA_4+/5+E42V,R\W0\#e_Gd
(3UO@2CH^N+:N.E\WJ:&)5V0O90[MC;[R7Y&ZW\VGP>Je0^WB8ISQFc]g;8g-Y;+
V>M=[?(9aD_)ILfe97H9:PJ@VZ_+J)^P2BIaab\[>,@d5PV2#O^]X8]XQ=6cGgg0
.;W[:b8NY[77g3FHb+1a3Cg59cNe@FG;V@Q&HO7Hb&A2;#K>@0IVZZ\2JGH&SJbQ
V#\cR0/ZV@DU^@<//_e;DdHN\X([8Ped35P<]6#MQ?PX/ef+0^+cU99@6\g+(QLB
P=4,g3OL:HRJ.Ca-a_LVW?)5K4WMdcfAE9:^9]9G@/#(JB)8U]2g/([dGB)<&N^)
D:Wd>_cL&NQVI[;>NgXNEUb&MJLBfU@ZWGMaKQ:<\@C9VB,#652C@(K?HWWR&;).
)(DGa-@YB7d8A^Sgeb0\;VVcL(:=>6Y?(7X@:#VFfcTd+[eA>3]S;fH\^;<?-]T@
(.bB&JDWY7EU9f(YdB9ZedMg@)N.PAA71Y-?bdQHcfOOR8QJXdg,B_78Ua5BB#KX
[Z\L]99M+deV,M/SBfOec(A.>QBQc03/7>30PN4_.?a;e;_fXY=A?R\16<NMg^Q)
Z7#R509[,,NFX4P@U]22?T3+.M:#29^Z+;9&P6[SXG[P/EDR(#B[W3CEY_ZL=Z^F
F]B7abZM6#-?Lc1C@MNP;;Vc)Z8OK,5f6YDID8:X3SVP7F[_4D(OII^Y&b@[V^=O
7B\McOYK6<C65_4GF)Bf^b3e:MbaT<3a&)[LEUUG-RAXCGF.#G1d=VI_7>SQIQ3e
.X1@FP?;c-2;426fZ=992+f,])C?3,G1c(VS@W;QZUAB_EJ1;EaF_<dT\KD9(IXf
9L,=/0N4X0D\W+<5DD6-5/:<-]T1(KU8PJ9NYFdgZX]8\=&cdOLQb,)]SM6/0[.X
S6AGP;(eaf7[,F1K](=KOT=PS^UeG@eC65f>_396f\f)WT4LC&/Fb-5G<:3\44SF
@;9@=\C?YS5-:<=)UQKKB4L#@^TSB8#4WI<R,+[bGSF(,(P#)#H0?HP::Z[L<VB4
JEgbaa6/J2ZC+HMgUfQQT,f+ENTNWG+Hg].WZbC;O<eRK/X^2Eb^A_C6..W:Gd/>
Bf_].<KR/4R:5Kb\TLL@MBPC-W_Y1aRF.\99O4e>YW^OHZMNI^S#_BX660M;271g
?W(+EQ6QE&E4+=f^Q0WO/)#)f90\:/1\^1UN,N1c/C][)c#E#_#KTGF0]6C.Jd7B
Z0M=4Q\)+V&EN6#X7WX/f)fJS.3?BVCF^>9GaX6,f9T7?Z0VOfOIYX4LTT.B[UKD
X=@e(/MD\F^?C\M>DW2P^Rb5N0@UGG=0^##)#S+H+DUX4+RFL1JcG@L:GRV)?Te/
a0KU^57[,YV4,:]N<RIARE2PNLF^YV5=dA;;#0+.[)60fd5+8^]^/B8OJ)]S0)(,
Ja?J)eZIDTC05=PH,&2][9NEU2.Z7R&5>6_QW\&MDW4Y-5?T&;T4<B9BX=MUQ7,Y
TZNSB]5[P:]_HWDZC1J\C>[[HUfa,.K4J&<M]VFEb:Q?1K2&_NFD>_84<^aB,HEY
cLCS3E2T]:V5KHa,=;4bPKI5HU@#_\1<-OYUYMGQGGF5,^9GcU7KfEA(MS2SgW_A
\Jc_K.6,RLH@GDg_OeDfJR_<2)Ude[A7W)?PR8G&Sb_.//XV5,0#94(=.)]##g7A
1c2bL1+FH=7SX#/(PHS#A)=OK07D&<<XP@_,gQ-aTQXX;/CZJdgV[&\[ZWJd7Yf[
?#d,4P=[Pd.0T;_2^-];9/N)G1]bgY;LNTFRbT0ZS7?SCAb#[PA:B5:dR4V0;>^F
>?PO)P+GeC3_VO0a5-^LgPb&e.ANUE]5RLUM?B(/Y(.fdA[-L]\Q0AgR7M/0<)OR
eBMa2VR[>R^<3F_KI,a7+P3A8<<K@+<N1FbRRaTKB=):.N?-X8BT6U:R_c/cP<-3
7TI_#S]K:V.X6KK+DFNCfZKIA@fQ5W[..UA]3<N_^7.F)BX.gA)QK,:#6]\g^5EJ
M)KaQ0g-A/ZLcH3IJ;D=&^K;c<c&/Ob1eG&QMd+\O2LgW,_gKY[#@I4(cO/>E/c0
33-_+cS+#C1>8GbcC_0a7C.)Q)M^aA_dQ,7N-9HJ09?@7>\9PgR;MgQP(<B_#E6#
#)aR7Kg4D3,3XN6<?WX97G[L=+H,C<Y1W8Z7L@cO00M#MHK,Z?-L-><-aL-2U[F(
1aW.&UT8S7a_+^^1e&&K;RUN6G?3S[b1?NGX;,M:&fC=&5gI8&3D4Y>#8W>P7RW7
P65M1:9YCEB;)Dg]F82K\<7RDKVBO^gL<&aP04?&[a5X2EPaFA0#X0&W;Gd=>(2@
aI/W>d_-c9&ZN1?X[K3YE@:[1R/GfG>Wc1O?7fMOP@bPAR1aH7c7)LX?Z)HBA,27
g/+@0La-7d,d<<Q1TDN#S0K=gR&a3HQ:gV6NZV4<L+101<RbG5C&@:W\-L_LRLU@
CdIZ2Y?PRd4\B3J(>+6g8:K\-.S.-4T>07c<1&G?@/BPaCa0?Y_:G4Y[]T.RW/bD
e^VA=\a<,5(#P7.TdbWE[@d+NA&U7O82FQ.Ad1G&gaga8Bd:3QJ-FEK++d<3>8:f
a7E#D6E#AN<3a.V7HK?M)N\B((<<TV>W4DCK22Q/0IV0.VFd0VXJD#ICSC-dET#H
@V/RI3ceR=<PFLf@GS,I@H,Q(-Q(BQ=g:e?.EfZK(@7S,O:ID@@YbI81a6]T2g\f
)cU11d]<R_^/TV[4&((]eQaHc(,E=GUeId?8V1dbC4TbZ9SNSPQ[RH/e+dc?8@^\
3e28XeG4G=@L^0VT#L-Z[X1T8B&CDXa44#_;NSf0.C?,/,HU0Q4LAMaT<S\>#Kb-
_1N7K4YRD(2-B?NaS/8/L4Og_<2+a[.>cY\TYJ8B/5gCR4W@W+QAS-cE@J.TY,f0
^MPCZG?[[F)=>?CaM8cIMg.V.fHFJ^9CU?;KJgfO<e(9X)C/G)Zd#Y=BfAVW4c=U
\G;7/3.8>\K[Ka4SgUD/U^A/J/U/@NZKY-=/N5e5)I9N^\_H7&CB;@deeM7AL)SA
.d,SdV?=C5;aJZSM_:NRcYf&LBE=aBIP,L_,Bg>+fP-]8A&-&b2AI1<\V_I83;#?
d?OJY_(EUf<8)84KUK_#;\EVPG/_Y(G\\@eS4).(]BWUMbYBR:Wf54JYIOZeR&V/
PO[JJCZ.gDFbMbEf<dYfcSe6HJP)2FRB-G2,fa///42d<QHDWeN@SY9B40H>QD?V
BROb=8Y7LB26aI5&U_?.R.4OcgKGH@W[/1UA4[\>#POAZ8[Q]AA,XYND:,^<0e;A
;0(\VYZ3<+JfeK0H_6f_8AgD5SR7+7<AR^AO>V^1<8Z)dDC_FfW[&0=A#D,cG5eK
e#36M<6[#M=1ZFAQA#dO6(6ZVa/e0Pg1G6(W=R,<UEcDO\H6)SEZ:J[:DeIXD^7[
a/,-KY.GX3MI_dZD4T]Rgf:4GCCb^[\,aU/)a_,XB8ff:GSYE:Y/A5d1cSC#NAc;
AX2<,WOB43N+MgEQ#>,ZT6Ud:e+8Q0F[+1^B115C>VRY0?M@<F^AUUUSVf+-:f-Y
;_&7.[I^R@^e?McDYG^Bbg6:ZZHP.3&0BfbdWOSUfd=4Pf0LV32]7)=VM6cJCAC4
^-#9@1]]P.dDE7INSC:0DKITRg;P_66Xe/ba[H)O0Y#0&[E^1J.#,B8[JPZaU)=S
?0\/.b10Y:K8Ag1GVZa3J43</BIP\(9?)Y.CJ/bF+U[)/R7S.;dW2WUZE-3T_OcO
0c<EUgP>Y]W;Z62OX3BDGaZ9,9[&V]3E4/fEERT@cY\=@1/d[@&:7MGN<P.SX-.W
>Yb0,6GU1V1TcTd=QbAF^<W6OCY,G2LaCPCAOUcPJL<LIM>TG,Hd&7ET2JQe08-1
;]6C63QGcM]NWg=TQQ=#,FHD?fG&VS5NXWSDM>dL0DT\X@_B?R2E5?K[a/E+MUbD
d)eH)ZZFD]Y?^G/_OP-CI??;,cUQ0IQL)(HE]?-eE&-0#,Pa(KOK<VBg<-&=_a=,
VX36_M1CY37#d5(@6#?:(V[O6a6&gKCe]1@^SNX[3Ya<e0@^YPUAN:L:W&:\6^P#
)L1@CSHf6FAB8P6,V&GfBQc2U-W5130KJAL^?\;[\F.XOc+P2RP-N<Y,a8Q<^M8)
W<V-L3[c,?@c.YH<&)ACUYBB4?JLea-?_:INHO,YKZY-R0(B]6b24]6XUF#6-d@-
_]V1ANL_Y>>;\+TP5XgSWaH;<)9E<PC5[Z3TAbRDH]88b/O6:,TFQQK>&H;GBCRQ
Ec3^+G1,8>5.5aAO?N6\7/d1He43.-J)AG4Tc<5&NM1]23(=gF;7F>8NS3(R4G1d
XbOZ4(42-2=BN(<H=O>I&C-7;0&]&3V(>DAaeM2:eUMS#>EFY,c;;a-7TGf&XXC7
):=@a^L>\O(;O#gBU(=>gDb@A1=4P.ca4&9db\[R7I9)@K#Q6X<(KLI,JDUF),[,
L47J](W]9aN8V>0&S\,98?dYOeE&&WV+O<M[dC)S(0I@3(/IDNc>:Re#2JPf?,_@
E(aFf5eSOeMNX+#W6OLXOXVX\8@S6JF=<.dWaURUHBXW#3SDG>643.EfdX@FNHCV
/GV:AJH[^GK]7,Z)E.5NYCWa/JUM1@2=ZOW1:6]TDUL]6c.@XQK&f-63Tb\)2C,H
5H3b6Q7C//>V_WXd@[P^@08fKU8GJ><>Z9L[F^&dHWMZ:0:>VDd^J-J3gaK<;W2W
c^V+540@=@_132G6(>MEA\D;]48V;M2PJfX(/@85W,7?5CE51gN+;8QJ-4R9+T<2
S3;e^cMNZ8;V#E>2Ff&5?Z4B6a8VMcD;Df&(CR2[W--4^[3JO3Za]57-JKJY?\]\
X^6KT[>298Z]WLP@(BU1+:M99GCM2gFE^c:cVC?efKDPMA6&J&JH;OC_0F5P+V(-
K+S-WSOO5U)D_?\:W#IA5O>@]U)PM>8d/?96J@?UB@^/L?FN:;WEN8C@42Y0CN@6
a6:KD1f^-^4LQ;J=?c-cbC[M^f1fOAEebCR@UEd)b3+g\#]/eVT&9CX:9-<_[<8I
0#aEQId_/]4.UISW7;F1X[fU#>FU3+LF<e2eWW=gVf@8_^#/c-R4XI^_,A9YVW[V
3f?g(T[C(a#.gHB3CXYda5Q@RH5TJ.IaPGZNaQGf3cM3/:XR9-KXc@G8/3NB53K.
[&La<+_MSUE>bXKV2LZ-dbe24d:85+/7=3D3XQ#BAW.>I/HZ0/Q5R,6a_e?U;KSX
9=IPWQdcSa]T\>0_4(MIE]fT_),fL)[8Ub9CI@-_g^1LD)-O3+E)@-\cB18cOUL1
.P=L<N0\?17^9WT>+XM2<>ZV>G(:W8#:7L9X-FcHCcaQ\FN\3LfWWMcaBC+XPJ.7
GAB\\c#E,<cIaOXW4\O7c2W)[(4C-1LMRDLO;445/_&#W2\FNG&fNE/EL9UC84LR
dXU.-)NXG?Ad[_>gO07&eO9O#5Zb2aNRIA#/KS,X\\>/e_5A7cSU.d]MTE8YZA;6
fQ?XM[V&;RF_UIV=\+XG;b>9.?5;2-A:e;33?Lf8/Bc9O.POVIJC.[=282aLIUKL
FPDG1CCZ_-N-50HF&fGOXHJ=<c?cR<R.(e:+GA=#WS/F@\L8EC;E(2^X?,H^PY0_
_#G>K>=cPAKgf.:H,#Z?)228TC)E=ZQSF7/KI#];?A42Y\e_SAd94M2#BQMV1UB1
UUD[DgBUQ)_4MXO5,K-\B1:PX8:D0PM(#YF-N/41</5+8GPT>[+?11W1ZK<9X^=[
dY;(NI?cLHCB9V:M&>CDW?P6b?UL?35/fV>^0C:(G/J-/63Z2dLd_;07g,.XS/:a
:5;Hc-X9V;?\MR,bRRBU(0=,54cE&=J1)&X#+HC>G9;I:_;:002STZ9+.L/LY#?f
ILRE,Ie/(PV.\+F)^bbN1G^0ceRB,:G@:BTU_U441K&6@RHRbDJQCS95LN>PGBJX
<DX@.BTeMJQ]0B1SY1_Ha.>dJO#HSWFR,c-9&2YbW)P;O>Z^Bge<7-FQ5<1H6OXa
)EDe45cg_Q\LHM(_g=c^<1Y1M[L7;QbB=?PVKBa;.LH7\<cC)f4OcVEF5F.]Q1Rb
a+_U+11=>/#D#V>-XbUG=:bQDK3#KOL6Z8@f2ZIa9#,YX&E<<TXPfNI=J.)5GQTO
A/E.1W1R&+N@8WbEcVaC)GN?G[YOTQ^M[>]LS6Q>V-_6]b5GO4VC3YH,0PU8#/eX
/R3],HE2^1J>?1&V.Ke;:f04C??+-/C6WU-8^U#fO;F=J9[90[(ege]?3AdP>(78
S07=?SDL\_AGP\T(0G93>#<5[_f5W7aH\)T0RN(99VQcXK)[K=f.Wa1.4MA-:AUf
MRf.M/2\;0,Sg+HI+:(T;=3[<(Y,aLb[^(,35UE9U>O1.Vc27fMg?c>T<G2S,@?9
4LE#-IbWdbfL-Y4]/ZTQI?+_c1fN.JA[@bTT_9:6#e\0S+7>g=,&A88/f1)II?/@
]P8)JVYAd-B+gMD]4=PMg/L5>?QTe7KVA=[,ILN.(KGTQac)AV5CQQ46gGgLdX7Z
P5PN1N+-;.Re>+f.g](g,C:N)9MLN:4P&V7TQDcA<;+W^1L1d2(0.G7Xe&Naf1JV
5Nf=>8.ec2&1)=fUd,.9?YO?eYTD\N,GS)9H2gSSdI]_K\_8)(-LKQSc6Lac6\#Z
+)c#L<,OVNH42d41B037B2OB)(<f;MH.Bg84N6MKU+Z]CcgQ;d>ZV&NEI:61).>1
UUJ-Bg.^>1aSY>+=KC=<AM@QBb8^SgJ=f<3JTdOFYEH64\:GRebd]R<VXCR3EdaL
Y@^SF-C@-P0=gB65cK8K<BAN+H7aJa>b6\4Y,DAbf-UcaCK3::)6;2P65Pa),M_C
D6FW(e,eE-Rb?;Q)f)ePYCT0,c\A3111F3KYJ.<0gDI]T@LH_;\@<0X0UJ[U]Od^
^E9JQI@a=@DBA&C=bKLL=1-V&(E#J\f(b-BGT5bBVMRF/.Dg8]W+/EbS(Jb6YW9/
_F.ee83)672Q]Le8]),_,]T4<G7DNN66XV]bD\CR<F7g/G)_N#Z_TWc842NMI&B/
PX02PQUA5,#MECc.7bW/AM+1&/S8)__)[+Q<\gF2g;Q@<,#&g\RA6Z(QX[ERD5#F
V\MB4N9_Z4LSE^0IBFc,KE:1+TZCf<+4G1)cPC#]cZZd[aI]aE:\2cAa:NY;7d/N
/@U9=XF_7()K1HVAU[Z34UgM6cU?ED6^HQ1@Gd@J([PS7.(?CNgJ@]17g1C\U]C_
:N7,ZAg7B:(/O+>=4Y77L)(?X(8d.[bNOSb?,1X-:Vb@0N^W3KBF,?/b69#AH]W:
B&BA-[V)Cg=V_+.>,AfVJHdJbf=TUA;.UdDc46XeJ#KE8]R7^3^:\AE.R[VVaXQg
UW[Z#[#QdfOc?.-FTN_K>[Z5Z44e.68T/)2;H5/>6-E7bG._^83R?^+d^ZScOHc\
+C[\<=Fc[CbIL\YTZ.(65CCa>ac9V71NW3)+8@Kc#=/0BV><fZ55#eJdCJGUJQf5
[52K1=HFdVa--S2L,AbFdJV4DAa=f)#8L;3e/f#^,&7;ZcXbH^.J\M2W&=eWFD:)
:2-I0/HUY[EB>TNg)9T5N=0-H?c,>HM\WQ;\]L(IU001IbGW3:.]A[HB6I>MZ(bS
AUN5ZWB^2H2aR/]AP=QU.VT;VgaW;_H.RO@D@<;(67/I>?.[_O0_4AN+cRT9d.&D
Ea51a\STQ08aEXW5\TJCN+[ag9:DN^]INR<JdWa.9bG(4XM0T.TS)/U7gI,8(Z1-
2:JXB+LEQGFS5ONYA\[bbN1Xb2WIN^G_MOLFH?8a&S=P@#>1COgZ>QV-12g]7cD7
&0T/I&)TgH)1;SH_M1TPE44KC?<Z[b]R[Le?Z#+.PaY1JQ#?TD>#3)JA4AHF<UN>
fGJ=ZE5d)2d;4;[cM[11(QfSWH&.AH3&[IcN&)e_Bab8YYJKfVZYURfGU(>?F6TC
YJP]^Ee=,4;AXL3c4G;.b?0GK18][6W4fBa)8HCCJbV#-KO2KLc4M,NB(LbD\&(Q
/bH:@>gC_1Jd@>J^-O#bPM2f/e[]_?SVV1@X34HTV;d3e(R&WLB/<A=WYHA.C3X0
GLbXNGO2,H_UGOE]O(ecCI@;4;e<#6&K=Hb)Z5+FPH-eX.CbTGO60@&A?-c#:]fM
e^U=\fd6AK+)>PZ7,g])0<b9[d#+UW+54CUK91/@I?3QO;75EZ^+&7_.M0XC\>(g
ZE<OKHIM/Ggfe50^YFDQ4,G@F;5)BUcA=BLJZ1:#=T(gdDMUC:a3&38,^Vg2e6^0
C1LZVIUaAE@NKe2<]]H8N2N#<6P]5F-Sf3+&bAaSeCALN&N6c/1MafVbAd3^;d6(
GCDaOLSdXJXIa/Q(e4K,CPOP[=^DW[;-7=+NJ9&JJ9][F^&DKV7Hd+XNE1L\1/:=
_W..VZGg8EV>Id.2@D#bf@?b@)]S#E/2+I.^KID:S4SSLWY0b9e#^JYeNDJ32E1f
Ve(E3?CJB):K4AcbX6_5=Eg8CXHfP]2Q.R@;e.TbOA#F-/;@H=5?4Ta.TZ6,A->W
TcDe6(N<#E\E1,P1Yf[g^L?AE4=c_LD=\Q=e[R1eC8L[O(9^W9&DS+TK-P2Q5D@M
e_6(d,B(5#fF(JN4_4I;BHD5=#UMDX)NFCV5NKU:E.1;Wf72;#^54@NL_\)aY:;A
]eP@Va,R9]\Y@3=OQK(\6fRV1U^4TO#.N:-3FEgU#N=N;b\&(>aGL6-ZR0H:F#0E
487(FTbKAUJK\(/5)[[BLVD4[M_\VKWJBS[a3GeBQHII[&ZgLVT1K^aAYA#;3HLX
Z6F]0RfI1HPVDRL[GU<LPbU#d;)96[^QY6COYJP#U&QB:.<H_;_eGH;.b@bB9QCM
]K+WT=E-ED9a)VGQBWT)Q#OO+AgOf01a0VL;JK(UU+)XIgb5(S:CL?+\3QR1feT^
]cIU@IeX.f2:75]=[2BQO7,R&N6WD3Z+b09#]B@7R4-Sb?&7V3&.U<3>T;DJH95=
Bg5OD1D,B2-\J&;aM@<7HN^U=+82:?cF6J]S3JH.-X_NEYRe-a>,?:GK=3GZOaJ(
QYH@[?/WBYV-:@&K3P4A\[USe:Zc4+bdD;&YU5LT2FV6Q:4_^Ue+5J](#P9c^D+(
,2+L+HV@I:P^/6OA.d4(aP^]3#465&X^JT45UI(F(:?#WN)(aG^3^IU@U@C9a?TZ
.XMERU1=OQ[f<6a)R+^E\eSOQ7W:F7MDc3YTV2X/EbRL6?cKB3BJ,gS+\,Zd=>-8
)084b;&II;^ZL7GMA0?>4a(J/4Sd.AeWBCHJP_aKBSf4A&EU,Z8KF,c3Jc>;?-<0
9X6:MAGI&1,a&<[dI8(WCTV&D\PK4^HRBM8G-#-U4X>9YJ8cK>TcAgY:[Ie,OeYI
W1G08>NbU523=[_?]NZ.gH?a-2X(WZfT/YN@@_@OJ@\K>Kd2)TR==8\=Z:LO53C-
X-a3TCH4YSEIQ_MTLAF^T6/D-Y&UQHU0MYV.^:0C9O:_^Y0?N7?>HIe<(>>CR/X+
DS6L#)QI7G#7].JNTW,I4IeDKPHA1U?H\,Q^Te]eU-.(GCJPH_ZRDb[AGATQXAV/
1?(SbBMTHXH9e4:8>:9NQ\4@/8_BO+fAaIRM^;;[>(],]]5,Y;gcR;IaeK>LFQPT
I3eTbUQB,f;2K-\EJC=g4I\ZB\.G:67)ETJJ7Z@8-)12;CLR:2[=Qa;^3XR1@58b
<.P0+dD(c&XSP/P/MGP5.RQZ(H++/873Q-@7Hg&MS(?OAF>ZT(EO[MB@.[LabTU+
]<+fIB8#QC,-KZNY89W(FTFO^JF6&N>B(8UO21Q.Y5+XbM2fb24:]8_Z,^#/[=.N
]07RZ[)QCW?W#&b9fe\I_LN(WM.MZ3EgI;LB?<#PaXYY:Cfa6E<6MGV7B0_,;?E@
(<g;E,VBL.=b136E):3VfYg]A1X1L/_KP8UZ[V@U)gECT6cR/-5_Kff&7?;C4Gg?
MG;#(ENZW@Ua4K&)F+5O[:E:6ffJ0b43<))-XHRGH2c,Ib92f[Q(gKKF]&EYMaV-
LFK-a^S=<fE7#_A+5QS>AQVe\3(E#MXg(>TBBS/KR^0T@b[BS]R\V_?ZSCK3O\?T
;2^g4@D?4g\RFQ]f4CfR3RDL<,KB^[[C@X(93JP[=Naed1(-Z]3]DVd1E4eKcJ,b
J.L=[9_)8PB+Z+;Xc@)3(F&=adg_7:c15=MRT0S^.RFAY3:bN[?9c)2QO_fM1ZIP
YFQaZ-R?3?)G_R9(>/BZ-^P)dNf1bGDTg1B758E6NReB&+b+_S-M\c6cSGA(\.9/
7He9#0C^Y5721&P064-[/TS=W51gQ?ZPRP5PE_TNVP?ZTX)+I@A=cKU[LCI]MPfA
)SPO;]WV2..1A0CO)\1ec,#2CdW9.FN0(,<2?Pe^,1^6Y6GL\8VKP^aM[ZdfAb_@
2Q?-DaHd?=-.,?-)_EQ9SGD87B^;?VVe#a3dg>NU--a2-U@=L-3G::GPFP#:]::E
]H+?+F)-7JL>7?W6W95,9<M674GQ3O7:4<VR7I&@bL6X81<(>Y(D;F]8./^W,BbF
ABJL\<_QG#gaK36a[IT(OJ9@aWQD3T_3[/-Z<JS>#a[P2&?-X]?Qg+Mg5GR1&(S#
HaKK&._^\:95-/d#.ebHZ:580Ogbf4aV3,F/\c2g(NO7XGH2&0,(_]99J+CUJbR?
B3GTEg4<#L7<RTM5YBa;9)_E[N9KZ+KL4KFJ=X0]WU09\)PbQ7)>6=SdS.BR5-Y]
M(adHU=XbFD=MMIafAEU)()ST3DdJ&F>Y8?M#fD1F6c<A@cW@TaGU?)OBRAUM&P@
\NKA<deO:(),Ba=E#JHUUBL?>E6TO>b)a,0UQK@1L\=SXW9.NYH;8Z0C62gMa=<@
EX7Q>;&VE\F[ec5BBK/.1Gg]QY(cVZ(E-E76J_1f(=#\d.E(aPJ>.gB;CXILPPPG
UA+JGK\9F#caY_EEWg)U5H_FQC4c;=B(<R]3]Ne_0D>A-PG:C)]PX(L0DZLJN(^b
d_,=]T#&;c.0H,C#9#H29+A14]YSeXS.I0K35)#eGO(b1\a[(PT52J0+-1XIH1)F
g6Yad3?7f:P4]gA>RSMD+0D:=P5LNJ\V=E7(-ePJMY@Ie_a@.J9)Kb\?ZDH1E3K2
ZTK/a_QIWWA^\&Vg+OD./eN+FQJ0=&&:3/O5EOSVYVcE9Fd6IQ#]=?J9D:DRBZ./
g.MR3g1YJCIP1VIZG<GU?[Le;+P5FJ#[<CJTaPEC?X;D/gJY^a]^<G@>/QE065[^
Z<1@g?].BGFUf_I[XDBX1aH69;dJK>K[5QDO&ZFYB[HAMU0&Ta<==La>g94ALY:K
1NWfGgc2?T6B<N<@Y@Sf46gUGGA2&UHR@e84#JeF7YGJ=EJ8X/&H.WY58EDC5EY9
/M_)0dKUA^#d7/^?d-D9D^Be:KHV6b\15bg2,\XS_.1FJKYAcWV9e)@e;=2]]b>^
PYG),b\g^KEJX=J6DdSH675BPB4g]_^Og>A7@0Cbc5QFGOfTA8@[g2P;E?_Ne]0T
JH2W<GeHggMR;^^cD]5@P(_Cb;cH106-Jg.f)8-T8S3PU=U_>XY1Y0#T2>Y3KeV-
_=_HCIBfV8]C:1;H8g&ZdcB&RNLB]25DJ)5gLCC_(A<G:=EI)7d3S;]OZfP_PTB8
&fZPGY4_9UPJWYcERd]KS,0Ag(3>_&U6?PbX]K(V5O&@NREQUM8P)Q-M&WD[))4;
48>UI7YELE399NcR2]H&W1E:1W;+#^NE.<)J)g^NH,;>D.(Z8<,Y7.Z(\/a<M_3(
?ZRLN<]bC6b;YLC9M;E6>:^T7:d=e54D)17I,aL^.(\5^A<ZP45/J17&#g,M0+d)
_/0#KHZ<5S]<JO/gQ20(\W&4>7RRgB/McXHa4dO>(7)/@/0SQ3;#K25_P@@AD(YX
?/C<=.CQUcd4Mg.PD#+aFIH?3BF?:KG=PV-gKc/:\1Q^61eH#5]118<ZAZ<Yb2>]
-_[HG@H98N1V?>W<R=_VW,c-7+4;5YGDFbWIN+ZUF>L^V3gb[ZGLK-OO?Va<7<f^
_B7?:2<T;W1f1ac,;0LfD8e_O<-B_@c;>Q?\ZOCA/dF+I8@VJ<a?4;=QBSLK8-;6
HWI2A?5Wd\QC:N/cQZcC1Y04I_Q6C/QUZ+?.g&#MPcTTac@c/3V[4b6R:1_2f/G]
f=F=fWc?=HF/4Vag8C5#;TV)6Y&\TIY,0BGIH;G>NO_KcF2I_QA8U+NR7]_:\-a3
).&7[=H56E4W:+I^V)J>O)-R;cB,?Fe.Z-_=1E&D\)T1M^DIP=YPYX)TV4&PY<?W
RRg-?)^)N@4QW#V4<9.ba&EVaeSS-<)[gg89#Z0UIR)E,Yf(\#G&0[)?.D8S4gbO
<[Z=^I-F#RLFW^_:@=7:TY773R+eb@dLaY)C>DeWJ:_5ZB5ce[]WMM[P=aNH>_M<
2\6F/@=QDG\@Fag8T()FIP90LWPc(ALCOH@V/L6@-E0_;g58FUeY#33623L<24Pg
d],/W#ea1Of,gd3H9Ob63LJb&&[;YM]8/-PW&BXC4M&NTbL\K@93B3E8K2UDf)#8
V3cYdA)+<BH^<RCH-6J(cNZN^O4,..\9XTV//;:K-26(L:AN]SM6dMJ-)2CZL2.8
b+-W>NQ-3+(QVFU97[71G,Wd&fXX8SMN(M1]I\A7GL3,b1]b7>?R,Q6fY-J5==W,
ZY/c#-K#3P;9aL(g-3:3a.TCOHJ^8)I6Pa>:@I6<-bBAV-V?IQ:8WZ(1.BYbag6[
7-(KV8O9b0?1B_YF_g[WX:fKT)[F2Y?T_:fA,9;BHF[f92:7LYXZP\.VPa>b(9W)
aY_N_a#g&@@9RK>:W3&S[\a@<LQ42TYXO_R]:0,F77(PcCg&F+H=X8)NZ2CK_7GX
&;eSZ>QAA;T1eJ5NU,F<<Q7P6+L4UBR&\CBY.VbS+eSgBVHegO/K:-[Q8PYEPCY/
.fg?-4XH(3M<_/YFg7.H/Bb_5O^#A_>bW;L&K0]DZ?I2:SEMaO]A@=8Yc4<?QT:1
&9c>^(I5&G8#XL0PCfWW1=0=\R;^J[X,=&Fb/>)\1@<65L0\7@:K:IQN?P:(U4\g
@LA1FJPXHXSKVM>,K:B?UeQW4c^YSUI2BO9=2cfD3g;VHY)VWE:BTU>LN^:@d;OU
-^NGbEfcKZKSX1YV#W(&aTVbAJDCb>8^;]PH]JLG]9OAU)A2-Lg_B[@^3af_b==S
eM1IeMI;gNS&VCe<JPT/@3>YdgAgK1E6Sa=EPf@VGQ&0G7g25P8O.QZ=QX8FR8Q5
[[.44X8^ZLB>Kf\0e^I/0#C(c,;fC6d2Z6_)(3PI8NdQ&Q^8+Q=OO:f>1BKDQ;de
OS7V2g/C3:]9V<=4RFDF@PW4VPY&^SKZK-7b-XCYFK..APR:L\@-c6HBJ@Y/BfQH
U:2e\g&?dZ&Bg6ZA@,[FfL+Z1QHEL>Cda^fE_&NK^=.MfE300X_;SQ&NVTHa2E3a
6:B;J^1EEKQ]6+d3/V>./7:I^C)7>\;WS]^a[X&^@PH?(IF5JX.[)+GEb1^0YJJH
LY5(Qg(7/PEcNQ8QT,5X1]W&G,(fN46^c=>KYT50c^\b0N<)^a2Mf8_S+)QRF#2E
[c,QXRRN-c\5/?0357)A7/0)..5b+O(6?O9W/ePQU-;LT#J_6MQ:R2XF0?UU8ILY
+a5IX]=J9B4-aVA]GH;LD)(93^PMe;3AYUIgbIf-P>6M9T<:NVcY;A=>;R7]\\E/
MO8/,)ENRfg+]LC,0GX7BUNP8@e9VG>g)TC[__6daM2Qgb>-91\1--J/cIWS0&CA
]aEPL,Q^ADHHR.\3TVT3B1>8#/@IQM1UOH,7,_\c.8;#C[+KYZ(Qc=Jb2R8D;Of@
XA6]=_,XeH=?3<88E8^P[8Z[,TI+\0C84-:TKgD7V\2YH4DD)<)SUC112I,GSM:5
>gU6)9[-&5O4.8aD,K#LK549&C5d7V@Agg\WM854PDNF86+LI;N>WI8O.U56T\[7
K15#0aX<:T<(:+,K,5VX;f7M\YUDOW9A.8]U#R3dd7F/.C:&M8d])/:D9I@6<-HN
@=.AXRK&&R]0g./Y<[YT_7bU#R-1H08[;][WaZGF6G)c_dcU9VJAK3[OZJ1ZN4A#
F+BR7I59L5H[e\Y\D:78)bSH8TeMfHcH[(4P\2Ib^5(]>-aVdOV</.K^GZPX)X/]
V.+80HAY<?1e(Occ2M4>Z2WR)[G9J@)8KZHSYW?b,ee\?&V4=2X@Gb/8K5bP:e7J
GMZN03P.BC,]\^D4b?Y?+56QcHZ(>2Z0N[NeVAMG-gYTDHdV3=#9e_fJ_NXKI4K0
fMM=cHU5U8HQUUdY0N^?<PMS59H0IIY_X.)RKW5^E\F8:0;4eI==[QF[+OU&P71G
2a3aSR1d=;@4H8KB\1\gH)3H&MYY.N(CLV,SCAT^EfHGC&]W8H64deK4AS_>U+T.
aKMDU^YM+@/4/A[)503K_V#+5)H<\,OD&+1Nd)M3d4\CZZL^]>^Z746_G((M41XF
)Yf;>-)=>PL9]EJ7_fD]O+1.<@+<6T[^)eS2.+M]C60OHDK-DSaGd^Q<fPAeg(NC
M_-S6[>b)H,.L28c8[AS[3XM4.T&GW1B=HD51ab4XX>;&SZM=P3(8]68BA+(?7Ta
fOM]MYQQ.<X_QY\,==^=/:.>=]G(SZ(N\W.\/cR^Tg75@S^gT6aMK,S;Xd=;UG@1
@gd1/81Z(>g\I]?-(YQ5EC>+DL[UP?^XA>Hgd^P<>fLHCK9\71GM]<5=.9QX1DUS
TZ_dVBL&&DJE54Z=O-=_/>_Q#)QJ=1RgNDd(X4bEL?EK_8?#>>UD)@KUTcA.G,E&
,A:]E[PUM=25>Y8-,XMRgI)>f[QF,GQ[a34R1[[-.b/eTK/+2JZP&Cf/-Q/XL<d0
4;:(60\Vag0eBS3a#>@Z,\>.YFg1HEZ2&F1Xf:E30JYYA;?E2,H0JZI9OE0.XC;a
Q>4PPQN[O8S#@8\(Y\c3)>H>=a4G28@b5\DG02[R9V=N7S<=3P)WV?(^6KC>L<g^
:Y^:II>9G\-eR[[2C])Z/eR[(06?\TNY;M:\LW#bA[8#/bR;?_@J(0\<eEMR<GGM
CU+E,GeA6cX7[+52,4?HSLfPb=53C9:(\P3<OF,[]O[:@<EXDO,H)B[7>X&TKW<;
(AZc=5f_aRFYUP4;=J)8XMN6Q7.bXUJWK/I9^G=N/C8@=U0b@CTQcd)3191dbP_c
dT5G\6X.Nc60?H0e&>Qd7E]U4K6bJXcTSOMbYeTa/I<JaMEDKG-D+WAW1RZJS[LL
E=CG2[-c(fCEKgM6.\HJUg7><8e\4DQeVC(]>bWAa+):@B#7\4WI\^CVWaSH.#a@
?U8eUW9N-:6[+7cCHVB1V-g+0,Pce9?IS#?\/4+21]cb=F,74G1I.+JMTZ.4g/@=
=fBK.?(ML3(44;.\&RHY10TD552(-S-G8V1)[FF#-3?dS4W#@Lg;_E5;E>&P^=W(
/Y,>Uf?A9\fdG:TQE:e)FP7>gAbIWXCa_)0:c1L/&XVa=_E59PF]5f_9,<TDYLBN
HK.9P4T<ES.M?I#F?B?B/AN7E1@gb_0>NC]GIbJM.#8RVO3g/N6/P8QL]/c,LDQ(
Ga6DQKaZ7C_YIS?1T0&CPc]_3Q&_&KK2MVQRe@5U/Tb#6<_-5)V:6RA7E]ML(=L3
FH?M)=2EKYB^KJE0c].0OI6QaDW1(TJXg7]F0.+.I&D\_+D)8ZTM/H=F9Ba7&3#E
M4F>^/6/R^/[JW+A=W[-[J6[BO8[B7_)DHcN83Z)9>T1_,=)WA@:=(gJV?.:</A_
[LdO5EfYaDROPH1SU^TAfJJ@6g]SK<EJR-H1Jc(&T)+_@..?#fFeN^MSSP5218/V
Ab?BY3gbX?KLG@c+a_TG:.V#SP6\A7NH:aUKC4I0U1TBXSbIf#W(MQH:Ee9)3450
=BWCc>fe(#]2S4EBd^-1;?\9DeSKPdT9VR5WID4DAIHe#9/,>A,79PJ/6^(CS:_.
5F>?V97(/AH1c3HfT0cO?V6.7M3]Bf?f,0O7TNA;A^d>UEd-[:]KED6GJH1,<ZZU
gZ,,/a[ed@CD_@?a52^15/VP:NB7TS?=J9.+W@75&@9QI0V(>A]gfL9\SA);L3+J
A^KRQe]bLLSN#4E\P5:;HU(7eOQ6:;[O8.#g7,EG<SP2dW(7.(4#2V;V);#E,a]>
D)X;)3O5W_cZKZ/g:JNMPM(Y;gU1[=CfZ.]3c5D[YX,Tfg14ZQ<IF(<>TPb@b>CV
/+M/P>-4^<g(GU7[(7P7c\;eE7GF&Ec4c?F(;&N06/L:@L[#(QZZ&[P7bVA<W#7Q
+^EW3FT.[BcZHPP5Ja.GB5?a-_[VN;>g4=QRMU7Y/>13U5d<TQ)V_,UEGBG\6(JZ
OTde13e<E3G60X5/KMX,X]R_E4cEI=2&CY,O[e\M=AZ.=HUC&^VF:6):WA:DR?/0
)OMIJ6Z//L@:eEZKK.;^E=#c;[M+gO+_CJ19(c[0[>;X)>5./&]/bJb+PBBMSOD@
F8fW#1fca/4RGeI7cE@/K^\b&QC?[/N5Pa1[[9FI,+-T\UXaO=OF=Dg0a>dFHX7V
9?#Ge?34&.S#I;+]S27FcD2_]MB_=R)>E/9Wa7ZdSR&7e@S8J/O?LX]4\5L\0\,&
Y@PC:BBODO]7G0M(d8)(8IR=&UMA(5H]\-P,,P/J/=_Z^I(^RgGYIY83;-K<E63<
:N\g@#)B4B09GTcEL,g2Sb07dcBW2(S.:eeRfA-a;ZD<IeXg&>\L>DVV>.RCaWf:
GK@X/b;]Z#)7T<7I@;2VTf#9TJ]Y\)@fB7e-#c6(KO9#9<K/PN[CH9U)#-P2=)5b
(V7V2L=Q46NF7Db\OGCY[B2F3E;edA:/d6Y2R^0(8bGLJ..GBK8NcNcEMdSKQXaA
WK;84-7LG60Z^D-<,^cO6&0J.+KLDQ77FEJXL9dPg=9?ULb)0O_V:3NM0C6BE/JD
.=YYRL>c\;@gL_)\d#.GXI@/0AWC@5\QNC/<Z->MMB(TTK;g[.=ba7^WDB94R2Ec
2(d?P#@5XLY26VRga8?a<UB31?3\bSA\f5E6YA\C)0N,/fA)[KZe-G.c[2K>UPV6
=UA]/EG;PTU\S_C]b.C9,^<c0gc@V?\Q\6MBX.Qd-JcV0I_0L&O+@M)S/@ABE\_U
a00BBX<VDZ65QY+Z3<(YWXJfcI28K_X1N3U=(VR>Kg29:-@QYfL+>44PAEU,1d:M
LC(2:LX87&d-[LY)bP,J&E/aG3d;]:K,UCIV^I0[Bce??Cff<)Y.^f\f5W2&)V=9
O]Wb05?1QQ]-bdZLY@3)5P6F];E+f2S#e=+TA:;#9Q,aV7PE&U2ZS-IdY?U<W30Z
T++ATZ\X-X0NSDY44@,-<^+CX^/9JK;?9;-QfV?^ebS;ePNb8aH0]Z2PBMD;MAc_
Z9Ref34(D:Q8#eZ32].WPJ<C1T;XZDN9HW)A2c+ZS;>YUV&I.>?K8U)_S.,AHVG0
J_[(Q/;8a2-CSEA?[Y4AGW+(E^ELb_95:DNP-YH0QZ<K^M2I@,YD4/?T:D15Rg5M
1f/]F[#R+B]^1^@?+ET(\8:JN)V,V?MP).Q<8eOeba4Id)b)EX])9RU@fOf3J):9
Y9LO[7GH1C<JfK7NW3Kg+J&GgTE^WH##W@>dU_?/A>@3;L#_V2[6/[C\T[=ZWZd)
E/a](8C\dZ=OZSQ[H<DL/MP?,/1@[7PSVIMNQ2DF/E,N.VW0_JYNdXU(]gE5MTT8
d1_e]4N^d_4#Ke?:5VWB/bEO^S&^Z9B&b5_(:#QJ9\fgaBDE@,cD_F^^HZe&.d8_
6Y<Gc+9O[T47TCWZ2MV/1/0,ZU1&+,8SPD?HfYJ>QOc]gQLfA47^4BCQNIbd7PAb
]?D3OZ;D+9BWg(A<D-GR_QaL>d>6K0GBK2+6P^QQRGK#W)GWYHgD2CD\4:?9\GW>
ZKT4e^][S#(WNE__/?+<3ONCA9+#RT3<V5OJOBY6QIgE0]1_dPf_JfI@Ve:2=V<1
JJF88>19+NL?\,Z]7UI^>ZZ=.A>G)AMc.4(^N?K(2fOT5,C25dE=:(#A./d&Gf&F
HQb1+^@?eHV[S/,0];YBCeAXf=D2\g09>SCA.@)VLG.;[a9<@<;g:fVV_4>P)PEH
E^C(fFUX50?8gHGMX7BI:FWZZ+&V\R83VWS7,3Y)Mf,6_;93>>.;<Q67DLMd0QJ&
3=H>:7ON?d5O98@75Ze#cJ4Mb>M\&YJ_MGK\EY#.&dBZU_aUI/\DM5X-S_T?>3K2
]O+ADL.,H:.Sc3>W4b5PLYcU1\V3@L(d0,gLZ5eYZ6U..,)NO87F=@A#G?N@7D)P
d_NbC1=T-eJNe4WZ-5><RIPDbB0[-H/+N<1(9<;fV>62PO.NWHK<;b2d&3?,,QG^
S\)FaC2E7B+7PHDV+b/6cFOHY_R8?,E&&bdSAB1&1>(:Ic-K0N=>RE<f\EcC]cbW
MT_WLZa8&UC8([<E]#6ED#^9Z/WGT1^.0=B7#PUC7<NNWX7.e?]@U&cEMLgbZJ2:
>7;^17F3b5][=J>d7_XRe;:_,+<DPSTe-]acC8+DW&Z+A-C<=E5.49<ELa<JIH\A
<[>=X[>Nb=FTB=8U2P425@W2UNaV2+=:^gEPF2+XgP_a/MPWZ[G<ID@7ZefA\5)7
I=;/J^?:cUDVFfCA3LPe_74bW-.HOS4OXQ&P,18YR,BL,,=WZJ_RVPGJI9\J/I,<
;.3OK.geLg\6&T)Q(-a)O7:G;T;9Y)I/H@BO\S(CG,U&?2Q.RT=Ud815,d64e&,C
-O1L)FL]1_VQ(;X]RD4V/8;ECPZf_BY>0Dd3ZF,aPYEZ^O+MYUJB-2)SW):fd10a
;cINR)VW;0^UQV[R@7#c33YASc.OLRQ_OPcfMKW1LG?N4MFWB&3?:e^MHS2>^,^3
D8+F2UaI39bFQb-^ae.<O\S-SHD+5\Zed-@Z74Qg63F4<?>YQ?4X7R5aNe:Ka5>L
6@4N+J]=\VZCJHNWF8)+S[-aG1#A^P[?,;A./PDC^^WRa__(De/E9F8@I96D=DYK
12^]c5?B,ZWd>QA?I8-0Ka(@Bb#5cK<]NdF)2Y8L45H5U:&:Y-TH\X42<A1O>8?&
8/5AFQ\GR1?ZU[-]@0adNd0R[C=Ha^S?D-KgEWD4FeBLA0g_2Q\&>:Q/U&LMVFcF
:S84>91I[@)6^+A7VPPg16I>BXa>69#PYQ7ANad8\2EXg.@a;,e(XYS1;7:)fA0X
e>3==dQd=:WY0<ec-NeSF\P=7@ITXGVE^/#b@BAA.1];c@12V]HaE]3aNJ0AVSd?
R_N/60.7UY=PNEG8)VPYEaUN1@5e7A2GZ\3C.+)RVGc5B@cCg&KC-ag)H&b[=YA2
6De1YJeA#HK7ec8,1CfG(U,Y4E#Fe@):_G82F>ZCCe;UXG;O5S;eI2_+YE(CS\[(
N;DJ4EZ<+=QI&UY=,6&@,AEQ(:f(4e1YQ_[7_I=1L,+U+<[1U5W_&ZfKEa#cP9&a
YdK1TK?(DTDR4O3JIW\=PN1^S-]C7T5V?-.bJ>PNWaXcA3<J9_C\O4PLFB??\UYZ
F&>>#T<HJGc[dTa1\+64N=N:PV<8,0^1+.2^Z>A#>]::@eZ^A8Pf:.Z]eBC6VGP0
PDK<@XC_CY,bN16N0YZ21U?bX/B2FA,g7NV-A:?1:=,.BbIY9#Ab(a3[&[/O:3[c
bCI@S@CJd,EQaT+;CU,_dB:NY0L21PR;_4R;4g547LS[)a;HSLPT1L[[6:UK,WUM
:XIaMaQ+VT5_2V:-S84H\?=a^[45,Q_:X-c^B.K\/=Dbb>:1&\dLWI0g,46/5bg+
E&LB?)X^gT>\N)JgE>1d/R/g(HCF,-1IQ4.6J)?.8#fIRU./>7<5W.N^=g(_d1+W
c<-A0Fb)gFdG5@<=#7]/dO2E+)E8IFGKL/.eM_bZ,7X4(T],PJ7E9Ic41U:;;_87
HcG(gUYaJFHX,O<CJA##&B(O2<,7;1(d,9#dJLN(\1cSFZTQY8K^D50?>+/PCQKR
7c]I8O:@]D_?TcH19&CBW&#:c2Aa5O;[-KKZ[82=Of8<S5Vca0e7;4d4P98)3&9S
+d7Y+.X_T()TU=GH\PUZ>JRTT;>3KR-6QB>=d#:G)+C-XMP>f](_JU9HFQ7^S=?c
?)=JDU=<F];[Z.^6_24>XZTcDJa4Y=Y;9f.dUSG(R0KKf(GM6bVP9WOdee9:#)JZ
/66WX6QGA.f=+OKM3J,/CFf2WQ0C>&,Q5<Sdd2QS4XKZCD=/<M4WC@)5@T5d[++Y
0I,fYG0K=T<dfF4[>V-JW]_SCd22;<7\JSa\E^)L9=MGLc;H72Q]+R=@I.NbRJ9O
H,2Q,S-VL(SB=faCL)INb_6=[?d>:#VHC?<XaN.Z5002QJBaUg>Z/C62&8Mbd=;T
F444OBH<#QW;SMa1W/<R+3?LXgQgMWI+;Lde>/#LH>._?47)D23Z5-1:;(5KId^?
8K(F+LMUY:GUZQ.]24=_f@cF9XE=>HY,)Z+U_#4<8gf^E^:GT(,#^+&]B;:N6,<X
c<.]PgV;X@cd(^H^LBgF@bW1]&T^bM,YXFD.?eY^51aXU6?2@II=Tcb-,f>)b?c\
bUM3YCP7G=0B1KS;ADP-fYQI^/TJA+OO,#F01NKe\c)7)2E+[cR?M4S9.@.D=a>B
Q8L/B47bg1T4Kc(ag<FAC3PY(97g+=/CGeF9Z++MK@Y6&=_XgB_GOFVf5U]=fTP3
d;_ZDCHUe8[Te+[@_Oc&-7VNBO3Y4g22HR,SbB1@c77(/gd?(K:b&3eKb&L2#/R7
b,gcGN7c?_5_OC2Q70^]5G]HI#N\\^LZ_cN)?E?_XWXLSV>XW?bG?/5aY:;OJb-[
F&eB)5+&_b[Y@2F+Vd3S7de(:(6Y(f?\9P#;@fEV#_KfQ?]W0_O0?0gZAg7^.9T.
5fZV@[-3XVQ;D(ORT\S_)5P?>]?9DRd5CF&.9,f2/XLBF#(4XJ]E_GYZ-,Da7B[)
RPfIXb/FX?].JU0:TOE;BZYON4;HQFMJZO<KE^4_)1X<gbIP[?HcIR(De)Nc@RIS
AGFJgM<M861H>83f/K.0BS3_Y4^LbaW=3.:GBLF+_bWT7SEORMTCP?=QB^8UfBM:
d-S>\5ad9I]UUCTegLY@M9@FD+;3V@Ud8&^@=[UTM13=ICbWd8;Bdb8<f/P_S(:X
OKZK=.@7V74>DNU:H2G+R2fJWUI^)G]_.5WSNQ_9SS,E4[/&,H(?a?fNaP[eQ,[(
R5Mf^<L7.Jb^[>/8M#2cI+/D6?_bOESgMRgdV&:=;O4ZeJLIR/AgF?UINOJGf-5V
YYSb8CaOWSV@UH=O70g(]O[5XEcBZ,_+e;#\T,AdMNL[K&XE91OfTR<7IJ22Z_<]
fD<PSg6>:,+XJ=#b<?XBJG9[G8M[AcdO/bJ/SB)@>;dJ^B-(<QO<MJUOP7GY+K_.
:Cea[)2K#DWW,+bFO2N;eVGPM:8,&+BdN+SgFD9KM6/f^?8Pb)OM^ETV_eaQXW(3
]=M/#Q_#U]HfLUGCXe/EfMc?4)7NL:N?ML9Hc;R.]A_:5,dBDA69VQ<M6<@1TZce
WW+RP<MI:K4923T8=EI+:CNL+a[K\7T,gIa>0S>VW(L1XZ47De&(aYP)M(fZT^YZ
(?Be]0L[)WUFQce^8I.?](DDf7Y2M6=5E93)QY:C30QZ@c/]ff8R[&@C:UEY?CT>
WLdaL\)B+cGc_KTSE7KKG0WFX&ga6,4^Md>^_e\]]LTJ[]XUO,c@](0>0\2GJY<@
8O0>#KY4I[2RLHfIDGPR6VN(3FLAbFEPT#-4fR0fMH@+W[K<K3#V+:P0-9F#,MC9
A_b;2,SEKBa6EFBAVID)dSe+LUddP7RBMM>eL:](Q2<52RP7_6BP&Y\FM@Wb^E,e
=dOeFT[eJW^-86L]#/?SfH](YNP)V(Cd:TWR_K)@YI&7#2CWH[YRI5B^&3VU(Q6L
9I=KeIIQcE;XO1+YK6._c-dNZfMUe#+_A[)EdEJd&Ke8B0-)OLBGZEdc,LGWGOVZ
/84X=2+YPQU&#K^MUI8XW^FX5^]Td43TF1g)Z=AZ69Xe@,#Y_I4^gH5#Y22E9b]:
&L,KG<7;U+-H@_465VecC6-UKM#.AGcVP5<4)XT=dVbONWfIcWD[01#4<VP\0+(+
5N@47cF\gZ49P\UOd&d=I?G5(DD&3K^IC]ES[[P)22&ARS:K1g^^L()D^dR31b[?
MQTMXQ)5[Z-J7O+GAV=?@\#O2VNK_WI;=A(9L\R,]F@Z9KC.c6T6YD8THbd5b:W(
_gJ-:9P^J.Uf,PFQ42A:N0WMA[+C5Se-;?KVd.:RCN7FK=AL/VJd_U)9K/;>/3V]
JdAICI;\(AYEYO@K[WT,XKA,f5gC93:f>;<05.229Mg]6G?U);UE\O^RbMJGB+SW
.\E^V&d9W_/6LEC>R]#@EK3=M^/RISKNRM6#:1CATS3>H9VY5C^:1UF/6?<9>DZc
KF&fZ)e1LeG^H>0,(2@\9HO@-THNI?+Vg@aA4LGED4gU.+Y\9E=C[6b5a\6/93RS
eFg;B^dBa1];1IL^1B\6KCb0FG6[U9&H109C[&IW//W>OZ9IPO[4QKf+DG+K/V/a
E6Oga7](O;Ie4M\TK>Y#AQ9D1IX#S51>83YPd3#C<=KQ&bW5\[;5?;/[=LE7(eQG
ZJc]ZH(\.GW5DSM9/^U]Xf3\_-@JgWQ3#;8FLMW5dI]];A69gcE8_c^#&>FZSN-b
L2M_>WI:ce7BI2Ra6N^0MMdPOQ+@e2Q(W)^EVC[GRXVM?L(CE72N()P:G7776fD>
.>JHV,EPgGb558IM&<V?-?Q1I;[<//3KZE6P8_DP]R8SB.f;=>IH5ag^]@^1BWf=
S?IO24ULQR+A8A7Ae-2Ef#4f,acO^Wcgg>5RJ_A3R22+:ON9QX/@1^cWJP3C.F>@
/<99,^M_>0;B2?F+4#7-Qcc]98WeW\W/a7N\(_gYX\/H?^_^;]b;K:6b/<NQ,DB9
N>/Yb8S=/E5TY\;3+P&7IFI/Ng?S7d:WHZVT>K1K.5#EXc6?b0HLb1--MV;[1<a7
N)KAP=PB=^?JSF<T/TP@YI[)NDJ.I190:?DN^U@AT(6(GR260126YgF6>7MfNYSQ
BUX6C6ONcDI]6:N8@Gc:6^+<KgC:I()Z7Z=[]K#P]):F2We4U.EH7SO>(=6?Y-2)
UF-HW&X,4Y1Q#?LJ?[TW?Z9P?Vd&G3C]@5&WE.RZ7[+]2[9RRe&QQbBMF3C>>0fD
+(b5EX[-3cX0QGEZL6XQag:c5eWb7:N,-.KS\H\;3ReWPU<-4NS@/KOWgK^Q#6G,
a22_?(G4X]2>11DU.BAUG_04R66O)1K8\Q?b>I/#+7-NK,8Z7@<H\]M?9a69\_7D
IY?]+EUbe5P9TEf.@@c\fe:ZgS^V;X;(]6+P4[>G)DT5(AT1D#:Z.;>QKDXZ#DK+
7.1&a;-gBdS1+(^(DMUW:S5-Cd8B[ZgRHXaW(_[6+I@]+8SH8E<Ld?Cf:U4[NMg+
1Q]?Z5g;3+G78a6G[g4Z#DH[cBNSfPc&QU@7fF#3MFF#)EYc<B=HS,O?\bV/e[/1
YgEIc+8N/^&52)&9-W0CMKR7RUW_+#7L8:YFEd1154>3VX&aRg3+)K3@-(>&>IRA
e9.+Xb)M)E)KW05<&L6X?g^0+f:I;Xe3C\2^-/>PP.4QaJM]Y3ZY@I9+T2FF?\g@
CFL^P)1QC]ZE[?,:A2+eWXcQEbQ(M@T?Q?#NFJ<d)H5bd(>\)G_1095-\B:J_\PD
PV;e&<gda.T-MJ[=LBH@;@1L+Z)Z<7WP&gfE^DQ:9118.#:b3\]&JT/G>U\G+a2O
MIX4d2YcMJ^WeA@VcX8=NM9>J)9=Vd&7[<[UNY=ZP/-^VSQ8bd:D+Q@b]Q_e1UVG
^.9NQaXE-B_QbNL2-bBefP(>4[WUZD)0(X/P7@95?)JOOJGO_0>C@.5(Se)P>MJZ
R7,c6?OIbR;M].5X<\=;cV(I&5SHT6:863&ZeTREdP+&QL+^G2:+a+B=FXZEN.D)
.8<Z)2g-\[Ec^d_.L/C2_A@DdCgO+/DgM8J+&@gK5];Ya9CR@+5XJ7;N5f(cXQ7f
>0BU]3ADcOAZ\/2A2?L823EB>L^Z>OKW4=b&B\B:76YK,K>0gEQg(B;-EQXe+L_Z
aO.HX8JB=b/QP=U]QISf2g?^5-DQUF143bXLQ8B162:-12S.1G5X[8.(N2,cd<2-
&I9:.gIQGBQJWS>X(8MQF)//V2aLY\IL5^Z:M=TCIUX4NTV^W_VFIV=Jc#.fOc<E
-;Y2N>SQ6KBV3[F,[M@U<PXa<e<3Q^XHc=Z@,07\6=;FR/V3V9E?K.)HN-WWOE&/
6Q(OTV6,Xd]E6,/G?/PCKY64SReRQ[H7^?B(C08.Nc8Bf/?MM020JD,b2<V:<eTH
0.CG_D<Z+L8;/JDS\d0<DJFXWfB(C[O7D4O0g#]874<5^_#AP-a=NG)=^WA6G4:^
M8P+LdEf;1De@>5TR4&PNU14\1Y?J&RZE#;EGH<,EG<>Re__>>HTC.W2bDbX0M&>
TJ_64_#&f9RXC<AH=EcP]5R<7GV0+,S+;T632^Z70)RE2D:F\L;HC8Y-#5B<S2=G
^96CDWF=5(0SW1V91V#-E@A0]3aZF60N<WE/gIcI18WE;Zg(-]EB3bCM:d71GMdY
J9X@eO^?VI_2F@UfX?H)O205/PgR<6^cdE+Y5DLN&Oef<E4/8[9+YTaPd,LeKTg>
_=eVDXb?8DPFXW?eD6T=2IJLWH8T9=W-.R&dba/W]Lc8@5[^+C^e(AEVf,NL4ba4
OYA_f8)>E8.RK<DQ<6@@8)a:F2A6NF.#^S:D:;71Lb#2T8(&;V4[S94f4gOc]_<S
T8E11J-6/@I;^RVgeX#8EHXKcQf\:eBM<-@0+M]+85D#>VfTd4MHH:gQOG;V/ZFY
CZ&^eYI4<BH@)H.\YZ:e1C(+(IO/<IMLdeGK8f;5@:@KA7H<C3\g?/,_a\-1J2WC
G.fO3[BP4N<<VPL6+\-AbV?7DU-Q\4GU4YD<0Ug4Dg:^(6U#U8NZ_E20UQ;:Tf^Y
f0M#89.QZ3_J;S)O@\a1AQ>.3dG1&-AMESYJ?[f87(NF7YC?5H,DOb^=TLF&^XI5
Cg)RFeS63,GB_B5/EHJ7@-OKJ5Yc/#ega3_b;d.6#P+TMB[+^X/-)XCI?fb@I4Mc
>UQ:>I#?Jf,f@&G\ODc\)@NLcR(9<1RN9DM-#aH#&]&2/c8J(@5GcV5+dZ@;9<IG
85@>V-e68;9NK9QX@-:e?NcHF?S0XYSW&76_S(_X#dD7,\W7D84.b81U)A&cWY?1
==b5W3U-C8/_L[3b4^ZURR/,HF=2FaF,2UY1@C94PV1DA)6+KQFMZ54X7[0I7/c=
=ceI[NaV3SA=I(UfVAFF,Z#<:9cc-5YSVS5&H@6Bb18IE49BTEaRecDV>&Ub7V6M
,QI?)@f(]7f)YS?6(>Q=gBCMX^D>UV.@(Z]?Iae>;;48M<8T)-a3#>;e^S0L@W?O
dR78(:,3^.f;8YbD#1<C-)DMSEZB#[QHcLGA(=[IMW2A?75KX-W232PCG)&gXYc]
3PC<eG/^M,DRg80J<N^CI6C]Q/[L->=TL0Pd\N[+[FdW/I^0ZY&cC1VDF3-,BR-&
aaYNNPde53OE]Mc=@#22CO8ccfL@E-XYNd[8=-[)(7PJN.(c]FCW<Q]>T_K6TBE>
[K9G=_G[^<_dC5IMe[F]@Ye,&a#a]&GfUB#\8Q.@<5:V4).a6S8DZ>,5)I]XO+-W
/F\6e,51<0P&^=6P;T./H&IVFVX;=(Yf(Da(4>1dA)HY>+O7+.)@B/>R^]EW#[ET
9c81N&VE(,\>g5_>dYFd@CK;gL.9B^b-?C+B^)HH<PNSYL98Q@NNc/:?197EDc[?
-d-98QX5FbF<ABdO:-7>f@>;/K3+Q<1AJ4ZbW/?,9eZ(EZ45(J#B-b(PZ8Db8V>T
5d5K;FF?XH_AQddR&YTDB6)E=Q^_6<bQTG-\WB:^08Lf@_P5:#1L/0Q.MJ<Xeb_c
]0gY;A(1XL=N1bUE@Wb\P=+)NfZ:ET:fM:;RK;J1&Z4>-eM(9-1^SHLf1\&CM,gM
IAGEZb,70Y,AO)^LYZ8F5OWAC(R+)PU5=gX/YFE6\+AGc[B&#?Z.N9+9>X<@35W]
8_C7aS&:S_AN[&782E]NAQCD;+V\F4a\RK);S2:?C9^gT47,<#.65B(14_QN<PLG
NI[Q4\Y^[:4-QBS;BND7B<]V>a_e/H=,;^G+W@,+BKIA.Xg3\,^&fBR7+_8Tcfc/
55,(7WUQe^N?#\9Oe1N7A?UK1;0LGR7]eJ:Y5&J8W3f?E2\BZ3+G/AI:]S:@C&g&
6W-,GJGH2H[(-I>B-2OV<AOLFSCU3XH??0UKB6IY-F<^5Pc-N@_I#1f^TF(LQ?.1
f+-Q-YE\JbJVWcG9WUKc7EK&OQAd78J&8_LKf5IdK6HTXS(GWL8G3;JE-NgW0ISc
&]9d;[fb_<)KT([gB&_>Q6SKY09YT?+3GO,)TAaOMWBXaIg;8+7-G=7VaZFG]g3J
L)R9JJN3b-F0P)^&IU\DKSV6FE+16[CMCVBMINWQV4VWV)PQ6@?J]bB2:cJ?/2,\
3&G2J:TIP@cf+BAHUGfZP,(Ac[2I;2#4DV5TeC^M=J-K,.T+F-7J1).1,MN1NNF6
A_/#1+cQ9=YZG/0UAQA0bgJJ?INX,4-F8_;UAF)Q]S]Hd+1-TH<bE@gfK1G/4e]g
f?=X[9ONeR,Q)cU@O>)Z.,&gE_^@1W=ZAX-8QU/F+YZA>9J?^^OgU/]>F_5\D=_F
,UG,Q2d2c/&J1.,^#f#,0d-&ZMd/TMMC=4K+03JbJ.Z]QdGM8<#XVEF9&N8@_25g
?f(^IW]C5/,09dL8^<OCfNNe-NEJDWG&@eM],^A;ARY7OKP.9+<gS>a5#fP0POBY
Dd,_dO+e:3_(McYO#9F=H,WJg+a:_&/BA92CE4P[<gJ#MMW8[;391/gC.^Y]f9;=
ODddC.bYW_.VC+-@M540FFbN^_1^PQX\5SdC/[+EP0SJLENdXHWcHF9Uc/)+LCa5
<VYP-dWN37_MA-ObBYQ;F[VFRH<73dQEC^_;L5c#Ic4eM6DA;0T8dTDK.)=P3YHH
e2UCI9W=QO?3NLcHLYE,5^N5271.@QP0#gedWK\P(.OA+Ia^.&<E,QS2=,4G:JU4
K0A#ba7N3?++=QZ+0IA3MBIP:QE/?:_OS@)TQM2)Vb9<cY#@/a6F^bXS1TcV[D2L
H_#0PX=]^0g5gBa6HSYK(I8#@\&e5LEN]c2>AG^H[+d(@VG-;6Zc+.6_G8E^1VD)
C&=[aa)726A[ZfD?ZL#^QB)(f7:<MT?Xfe=6#fE7=?)3DULDF^X/SgOD8[-NR\bW
.Bg(c3OT@/)IH>BE]-(f@L(T704)P?@;G=[<TC,]#\dMZP1aDJR3WA80O3bd\ZTZ
cKR&#?B-b?OdQF<A7)]P^+E=E]fb>]:XDX?g1Cc/^M]86I-,-G9dBRMQZ[dJ[Naf
deg\V(B5eZ\]GOfQ1TP)JWb4ITNS8bdaQL03P;);LB6HGGACL)];>(P8Q[;C]RGK
BHAdK>TJg7(AUB.-&]6g83<8L)E5SDaQR\P#5VgS3OLM&^Q:,fAUNK2+_RF#g7,;
EAg.#dY&Eg2>T[+G(\=)-6CW;?W7(BJTQLBFH;;CL.3VIA+3B2G+P(YUfP[-23)U
:MR4O[SCY:c5:SK9&U530c=MbJ#5f(G5+KI\1eIdAN;R_<U[1:CJ[G^8E)7[Xc07
I<3Qb.]QEdbe:0g-c5g_=>J]Y5UgT5XV1RcI&_GGI;M)(EPB@B#@ObFZ<((GP\^/
:L@.=eg;B7CW/WCX>gXS0UUUPF&g]23&d<L;YLG+IHBbX>&V?\3FB.-.YH?_9C6H
Z2?-KN5#+VFb,3g2&;(S&4C3IB0)8E,[^L^9O[R\3@AL/4XYIVW9=-?6?5249\+)
.PJ<gcY<TA6I4#Q3C&9X&/1K/HaCRF6BHD9[0Y72L:a7gQOR=0Q:UUe6Db0IC[3V
J((&<J\N;KS<(cCbX>L.(efVM1&5(;dgVV5R6Ec8-]\1cTe<b<^-\91V)5a.95PX
FGDE:L30V/J#aN&SNC+Z+<c]5f5-:&c>E(U.77g_gKf4VcVXCJPV,XU<CZ#Q#P@J
WJJ)1^6+(aBZ\GE+MG:W&7&dNG&U8@KcO\7G<X;+9=bg7[NBN]fEb12fQ1Q&V.6,
Lg9dTg7?Z[&\a0:9+SUVGO.DN>:QVa-GO@AJQIbPL.@gg8)dTM#&@?L[:a&->2+\
g,&-I/2RLS-S#U1->DI^bS+?HTGTB-&eJ@X#89)DeQ^c@PC8K/(-TX2AA-NUJ9-b
#=9/aC1<YXQ>VY;\beF<KCA@#BAC#T4)D5-BAI=]^-^)F>S@P+_QXPM+g,H)-@YK
a@D,W3EK[HG^5^F04CC4]61KY;5\@9X5GR?-(0HaLgR@Oa+RFT0X\M(d5DYAH42g
NNLV^cE]fWOND5NLM))-bH#;bO1/+13#F4Q+DQW^9;.KJYa77b)(b77W/3-Z3R(2
1SUR/6/d]dc2.2:=fTN&D_cK+7cNUVcP>PDZ5EZVfU#<>d?B(7c[43eJMM^.^T^G
LgbP2b_N;<YTB84+=(A0(BG+?W<NP7=\3QW&H2#CYcS8Ha)FFaDR2]DMFO:/)c=Y
1g/YWF3\J<&Ba-(<g6D@_7FWJe&e#3R?)US?Vf-7A.6^?.WV>JIL0+J3f_>.2eN0
>b=Y8DO7>)7J;d_8H<Rd#8[&#TffJ_c82VN#DaXJDX?.\5<MF-K9_VJeI0:IU\1J
2b9W91g:^d2^+AQ:L<;/W)?03B-0E1&6-R4e=06_&;/G^INS5W5<:_H5\egf7#,.
]=^:0/(4_\6KH3L>O>+&IOaL)S2MK^ZAM9BEVgY>-Bd+EIQ.R/8=_#B0FFT76;cT
.S\&;_Z=,d<4>:I7[&e(CXB@c8O&/21;g3UId@@JbS;d2;2AeD,AWPLU.3#_UENO
Ta66&eZE8(D;I[I#@<ZA)&(LSUH,[#:SY#<UI_eD9<82;;J_XQ^WJGa-:]YR4d]J
N&Z2L6?^,\Y>)@<?Y^cT03N=&K7KLgQ\5W1aO?-IC.O4BO+Ra>f5\,g;L/aT>QbK
93>/\MUO6^A&e-c)K80G9C4HYJU#6fD0J2(@TSCN-HRa&5SPY4f(I6?L^]67=(L&
27;.@</#f5]T=Ngf7J;:CM00[TQPfIT-O.T?5HAU\>H<WEMYEY?bSJGc1E]BM#@/
<f.ZS3+1[GZTBD<TU#;9dE[JKE@=&8RA4T?ITQf9AU8;Xd<bI.:3VN5#.^0T]_(F
VV#;)L[U=@+.=KW<O5V107P+D,MN<C(Sc7,+OFD?@aWE=C]1AI-EAX:1bS:I=d@/
-^G20?;2eSZ)=G+aYA;b->3^JN[7aA,P<RBJ@[X@?DVP?24Z+V?K/F>_dAA[(+eU
/a0)Odc\84G<X9?N;L:c0M0R,S?RN)+(bcb3;^9Q3>EGf,DVOZ)1Z5>/HX3:YXEL
.#.MYdG37W?#VJA2R8_Oe\NCPF]G\bJ4Z4R0-eS57e4eU>EGdcBGa.CE62M2e.@\
)1?&AYPQI69Na&>bN;d+8Y::EQe#P=.MDHYM>\;g:SKFJc.;3f57]6e4HFeNI@M5
P8c1?Ma)S>>FdcZJ:8dK:?/J]<9U9P6S6&PG8V0V:5IJNF/XM8a:0Jb7c<UI=I>N
d_K8(GP=^0HUMQ7V&AXB(+BJHX,:GZR__e^Lg-?fKQcJ3GB;O:VV57TbbH-EELC]
21J9U0JDJFf@g9R;L^>FRS+]Z=R@eJW#T43J3fSRb(XO2[UN;H3J<dKY4gf_=SS:
\O9MgbcLPY.=1<C-Z(8XG,JXfKX5ZPO[[ZA=CEddK2D<266,/Z]9U[AReW8SaQ7<
WE3-35:3N6W2VM\ba,V6d.F_CZc>f;>+L0-155/MeLMGFZFSeB@->Lc91>P28XKY
f3_YIP?+6-<7WTV2ND1L_3fF:/OOVe/G[(;H=f@1>)f&CLH,Z^>g.E9aMeFU.b,L
V\;Y1LP)f[S3,Yb>JOD4&T>^9V+T377NQ)YML#-c^7fJDcJcRV4?>ZN7/Z7T7_@0
6PM^)ZL86K1D9+8ND;N9.TU-B&I<+KIbGQR+BQ:&fKgg+2B(0Y[g.(N+>:#\HG3d
fEAHR2+M(0_=g(a<@];UQ5f-<_Dd-0bM2X,7eD5CgF-\UQ;S8PFMNJNL7G&9>g8=
4@^8K&_:^T8,GMcG4\\AGFS5E_MYAPPS5B0\E&e2UM:ANPE9;b)/U_B3G#PCde&^
]1H?a&_K/bgBK-_Q(bA&)=c2[Oe6H74Mc<D.S_,<Z>5cR(O]:Jc\W--.6g]81^H8
Qd9Q8W,[6FC8c_SS5[9;?Z#JL,LECQQ;-Q1VTLdBL]bK>d)Y4HN?B:4G?>G@8D&]
e1MT1;R^A/5bgIEOF:]CM]SF4K5;-DQ((HOYc^FB8]J[0c3b53:QeO2EBc97T;F?
5&MKN:#B]]>,>>]#fX6SL78[UX;K[R.^#R98#GZ<#7:Te[Q&,ZT^JaZ2YYE@T48W
42MdX5Q@?Y]6N-TW]=RYH,;27WFYgI24;R>^Qg8bM/R;8OgSgX_(U,#U#T4W)HP3
YKBI3S^<cUFU5;3PENZadFSe6_KaU@6J0710K+Qac\g@+Mfe&Eb51;g;?A0X]BZ0
gA\)JC0^]:1#7#&D#?1.EV@@@KgNNB8GY5_Kd+cETW,09^#,@8_HeaAQ&=c2)OXD
EbCHeK3]eIRcHH^3\XP(8PSgFgQ>4e]N+,TL;LC;9UZ@=(^52BNG\GINPU3S77SA
W\Pc4<09:E@)^@?X2DS2VN@Ya\1AIGTg?MaYLVSQ#2a6EK;c&Q/H1H[Z\-e]ebPB
4d#P4J@[:BV4M]5WI&[c/:.=T0_9(QTD7c]d3Wd+]bIHI))=LPa:BbE8I_0bY(BQ
(9AV?aNQR^Qf-:T@GEcTF&BGW?TM?WMJXf-H47_E=0T8.\5;<Y=P3BX.=7Za\G1Z
:\;^JfgBO8#I,5,C<3He/,+#[DF#OR2]MRO1EK5Z\O6LXBSG4d8fZ7Y@/?DHcaML
HE6\Ad]CgF3RR(&O0@T=d(ZRQ/W^:ee>EE_.8T+TD8aN_/:4R?d@:O=K#a)d-,aE
V4\RLCLeRBCYD];H]=<=.\OeT261Y\6<>6b)S?cKg:F?5S^a=dL.Eg13DDQB6[WQ
97AQSSOIGUaUZ>JEgHE9feOB.WF/E0YM8TW3Ce6,RX/5HT_#APSXG__-]<^,TYLC
]aNR02C;fKGOG1g&6)7CF5@d(_.(+W(MZ3a^=I:@JbL#X:MbZLf,8[e@AgN5LR(J
8I<4:YIM)&NC\ND98DB(Y#SLVMA8faO)>ONeQ/@cVO>ZH\FYLIS=Ze]RaJ#L4+HE
XLB+V5aIaODO6Z0-aE^>dWT-g(P@)KdUd+@2F-[>cZ+\\J?)X.H3Q.(Re>#=?IXV
]JN9bI70K7CRW:0P^SL..^((W5F/\HNPN#,C/C?=BSfHfN#91g9UaDdF/.dSMf1&
^[N(ZME0]_@Z7;79\[XM[XP</QG2(QBW8(/<V]V8[1=0f/SLI0S/V^P.O<EO_d:S
X?QK(FM\OgX8a+9Md8?\;Yf90]?NL@5/_Ng&?O^+W,9X3#Ab<IAD_?\W\_=Y<7)Q
?C3_D<7L1XATL6&Z,LBXcI+[LKP)0X_7Z/L@dFa\B#MA2S/<]0/:0gf0S.\YKG0]
0Q?e?@ZV;M;]WeSVAQMO,O[,4;POa]H[KBW\W_-61.LONC3GZ=c1;.Y6IW1HY)4\
8RXVUV6?HF<,d+5L2U_?Y8AFa:GcTfX/:R;=L>M[LL6?\6A9=RAT<-TX#T&&W5+.
Q&_:8)U3YK0?X2I-N5C\Jb[UA0c8PRI8MPAH?/_M[ON?IS;3R]4eUC<Ff5UTd=EQ
@WgH+8?<C1HJb69HN,gGQDf8WC<YHD9McKg[40:,=_(6PE_F]>^:eB7C7U^R<T,Z
UY;8F8NZ,e5\UYMII7S#ee)V>@&4-QLKAOf>+g231/Q[;_@B+e1/U)M\FWUC,-+A
]VLXG<@_]-6;A,,5<g]P^7EZb3QW4aR=6U+e6d,1.U/@#-=W2^6bI3K>T1NJQ8GK
aOA=a)dae[P9A1CJM3@U)^D)4=R2fKYO]f8V:\:1fAF-X:aD9Ma,4W74C27T-;+5
-&f,H0L7J515NgdZcG;+I1B1^/IWM53+62G;dX:Ea=::E.43RL?VU@(KX?3I4=30
/e9bCTF5B9&4:^6+=M\\^bK)E]CNNK5^S.U7:_8\QH2(_I-KJLLfe+1[bQa:_]D8
e1:ZE^?.R7J\/f<P]H+9-R12)NQg3_L+\SE^N/3,8E2FFR1dCR^e(4,9Y(E#HEC=
QAaW3SS@,JR6L1)gc.5g69/eCF:JI9GaRX5_IW(ca@3Sf(MX&(aD0P439-KLC,aJ
;Uc^,PLJLG>Pc3SNdKFWC14Z(4]5d1gcGeQ;EK)U=(Z2B=U[BT;VF0OG:=U>IQ1X
RWLG@[U+b-QF)]gaC)=T/S,_R#7C:MH74SIZb>7LB&GIW9&G1UQ&1,7\EM,(Vg#(
J<C)56(b),J;G@9)/>-D(a@^cL2=b^<J+U(H/0Dag&Y;Y>X)6DBK-#4,^X8Wb:3e
6fH)68Agdc+AgM[M51A@+T5A.MGX85I\]Y0:+cX>0^UB9QBN?>Of#)OYBJ1H8F)3
U\^-^ZD\97aPbG,BH9,3WfR56\<3gA4\/d(W1NI+ef79O?@+\IK^c8_QHLV^(Sfd
5OX14Ue#0gd/N?)aA/V&NOBU4Md1RgFe?3OdO_c+RQW(-2E_5R7fK#=U:P32)E[_
JfFZ05I9Wa16b.Ua)2aKPRX93cP^fe^aYERJB257N@;5&M8bbTJ4,?6VF^E(YP[@
5)g0ggO:V(g&^[(WJgf/8VQN\Z;dE[fgDXZ^[#UJKL.J:]\@?DO&g2]a6P]/Gd4=
YBD<L#.>]C[&+c<aN^[.XIaS/9DYA>ab=d0X(;3H@eTQP7=PWT]XaIg6&SIfMG8+
=UH1,g#S:?[O,T3]?5&?A1;W@X4LSUZ^0?9.D2>d;\,9<O-cJ77]eJ8)),SXMO,S
=PNbe+=Pbg1aa69b>-R3?_JNO,3O5&#G9V_cR,&]5VC[7DaNH/6(bP)CU9V#,UR7
J3ebPcLU[Uf?&[EVdSCAUHQ+.-P:WRP4R;&&T&U@P,6fIA_VC63/.F\T09;>B08?
2fJ_EIb9d16cM#\J,0aCUAOcH;&<EV\Y&gWTT7R:D)G[@>@[Q1H>MKJNd>Lf#a:.
OK3e>Z5e+AS:LbV/3KQ#R#3RMfUN5ge9(QF=GUTLa:-4O(0^(=IW<JDPV>91:B,6
L2CObNd.-HcH0805D8I\L,f;1Pc)Tb/S;Dge:10-I=?S,11[?WS8aB^9.a(?a+EF
?2\O)TK+.J[CDI6.N7c+DQaG,QDf>8+Qd(UCVd\TL74<X=[BJ5[YO#OS4&2I@?4f
V2D2[@Z6)UCP&UC?EUeZ&((L6XQBM7=Ff>b86@V<J#2Pa4_S.-<b3e;6+V]TY[DA
aQ9;87?\-EVZ1_H]H#LH6_;M:]PU>)N&NH[M&VKa<P)36F_@U,X-&1AX3LC1\fbe
M^1DO9GIO_JYOAY[,_L,aC+W]S-;WQQaCTN,R_P4;/,YA/5[;Y6=:dc]EDJA<fW=
=)51,DfC+C=HX7+Z8cFUYEC:^Cd?9-KX5C&../LP4@>N(0=e.-\5eS#(MTVU:aPc
TBB]LA=7X#2A4D-\R9B^1a=IZdHU\ZV[ILA?9b(T?<aU&b92KCN;MLdgbDYJ+Q_\
XE-f,/+O/cN;P1.EH(H#dFg#(G&^XUVM^L)2G8EA^g@GFO,L;9(6UGa^J<GP/f8Z
fR32H^B3@EW(42RQg6>?DF+C1U.5W<MS>,76VG+M(K42cYf(?@/:^D:fT_QZ1Z1(
AM+-P-DQHCAbTY1A(-]KBEPY_Md=3>fSfcJZCUE/aR03E(\N]1f5>YJ.&EDXXXQW
()SZ&OYA(g;&C;W:Eab?W3Re-4;d7R#[Ae,[/3#2R/OT.FALRGN/g_+a#IdbUQR[
gHa<92NK95@:BF\NAU7CW@?P_/Mb]5dTgY#=_8(JYYffP^C:]2dRZK6eUfc=,+L4
b14EfLS+H_^bO+Yb\8Xb(\QcdX&Y=T>I<b?.b6F]U)#UYe\,c6X];/g.<?2cNAVJ
:&.JeY6.X?M&G(KPTbI:&d;4.PNV9-:0\aULD9H)dLG.#eX.,cOaa6FT,5T4fI8+
,E650(K;c_)C-d/1AT\?AY/XB+OQ)AP&E02d0)7DI[_0,6f3Nf8H;ALPAY7RR98\
I8FN&Vd5HSL>L14CI6)2BaE=Z-(JH&_8-Q?0#?N[;?C(]D,ec0BQZ<2Q@;WXcXbA
&.4C@C#B&b&/9Ze?\S@9#++JU4>+9Q\UDeM-B<Og7(EUGI;dQ@:(XG#L[\dU-EC(
IBA3gRN485AE>+.._f+QBDb:2LNAF:60RAJ?ZUePZSU49UY7f_gSW)YU>6bTUF6M
9fbe^?8?bONOaZg.TQDJV1V&8fI#]:e\Wf6[7RQE8D/V+9<fdf.W,JbAe,XSVHe2
<]=a[QP8P6M5\BaAJAM7)ZPIaeG^;[TLPZ3<cZ2.0R[R#1_)EC-&)H]#>Ca>VH=:
^\Rdbg.TL]>?W)4^;^g3.U8)g\gAe@515-(J>Q_#KC@;Q)I:)3MM6WD^^LgRZG5A
PD\B]_P01Y:aQH4TD<gH8<e@URR=;Jc+HHE82Y2C=9@0=cB;I/YF(5.=+:H)+4T7
;7Y(L=E(^R;&5S/KA8S+E]_AH+b4^F;>49S(B(bYJ0ZPf0]ScdMZI4aDc#1:YN,e
U<OYb9C6F&.AL+1Q,::[<#YZF0(2e1?3K3PS7f7R_ZEECEdgB+[-I>dA2;0&#[fL
WD,+3N^)84@B^3DJ=)BQKd983OJ:,b)TS]=W2M>6DQ5gd0ZQ9AFT_=)6=##QV34\
e>/-4b,RL69ZV?aYXcGVOWR5P]R5\15g[5,B)PX#_=WZ>09@LVVF>4FYFV#;cO-0
+;N3?_ccgY@5-.RYMK9BBB2bXJ1\M0+_fQ0L2957.,5-Q>1ZN^gY@OEW.7OgXGGd
b-FWV99BQ&E.FO=c7N4LUB@e&Y7:F6Y(_-M3,EgWe)Z_:D)D86G8d/QJ_]W-B=e7
8,H?2S1&S[-G5TdQ4aWBYd:H:18UQR^0O89b9BcXNPBAfOWHcD0I3HO#I40X5b>V
0cW\>UYMO121ZZF^SgLg>[?f[4cIS\+bI)30e7;ME>O]2AB<OD7W&A&@ZMT2<McT
5A+3)2\#+^a^3]eBe+,ZAaAWU(QIbJg+O4BC#V&W>?Z8c@fV_<bZMZ5[TJB;NA7F
Q[]O)894(1f<_3^@F[]K+KEYBN=f+A#D9)F@:5?:A<TUM3L0/]2Ya3+:(<+2#-;E
O,?0#4^X1:1E<KVLc-8NPO(BdH^39F:JZY?5(Cf8aYKcXRA&gZgN4f]F>]Z[-=H7
f?T>OU9(_+L3,__1XVa0f:A,8TdLB,JF.c<7((2E:75GV7OFC<J243RQZAT9.._R
RdU(]8-U4)@B_2&feaZE)9#N,DI#49S[:WX#U]A1(DVcR#^=(,TfV0f5RgFG[(&a
1cVG/8-ER0?\B8cHFL]2ZS5X.aKTOdORVP3[.3f0OKH<YV3Pg<]gg(SMS<R=E>H.
,O1+^,88,>4K^e?J-YVTff>[MMaF,VW225B8=[K(3(b4&gGKeZ9,)XQ+W)N6Na?>
;^E2<RLOJ(W_;5P8A-&.f-RO\&AeLYBeB@<^Ja#_&Y(T<G>\G/V)>D[5]f\EeZT_
NA;\C#&JL,UYVVENW<5G1P(:Z<VH-7.Y1Z(OKV>0_D9-9CU1<&QY/T1&AFdT=QF&
0IE6H-(Y])G>=+I0>58Q8,aT-A5/4HXJ#faZA8Ge1U+5NRR>9gIRfTcGBP^(>+c/
4H?K/V8JY7-QWB76Vebag6&BDbILJRfFQ);[f7X3>.gQV=-.&430FQ2K.TfOW_NN
F].#3P4>MI1R^R^22+FHDLD79(42HX+;\_?#HT.9)(F9-L)SS>b6[TO&E:<g^@&0
g3>TK<]]LS,C)1Md&8;I2_9L5T7de;Xb/^>3DHW1)N21<Zc@B0G^1<(:MBUCJ7,c
(X[0aIUWJ?W[XBY01[P[F(1?PBBYWB(;&YASB@97C:05Qa._JZ\6K_>1,)_?WAM_
/E-EH57YfO^E&F[eQ?GZ,-XM;#-[\,3e]-(W^28(I=P#,89=36&TV1@D_4,O)Kf/
)c=PI[b.H#3E08N]fD90aN1bGLEgPSd\TF,_8E5ZJD;:J49dFQ8UXUKLe.Vf&7]+
#>eO5<SYIAY20__+4@3K\-3GKE:U&#86#VOcgB:BXGFWRCS;\BXcdF=AFfA5EGC;
3Bc35)51\dWF)(&FSgRa7aUHSH5fF</?NI7GV9AggTF7>)JY]4dJ=_]^4/gc7FEU
f#-9=N(Q60ZJ)O8)Y@Q@U7P=3b;)]5(@?8Y[(.<&2I5>&EFIcSaPYS(b(-[IS.03
/A=N_&279EA(,+3S^F-PXWPceABKc,La-6J#001@Ke4=MBW)R(_?(#=eVO7WHRTL
80KMWN-eJTaYe2MDA>R#2=;9;RC#aa3](&X8a7>YHB,7CH)#K>E3_6^#&866770Y
M0E.-;7#@T^[37<SfA_G08#GK0aL?bB<5&J1N=#]WU+LMea[_?-30)K5E+Yc_&U&
\M#>(_d=^P/3]WVCKH[_c14IZ]7?.,BMbBON-/&/]:K+4[PG7]:Ra-8b7_H\0d)/
QFHec2M.<E;I>^./dLX(dQCK17>HcEZYN).8Da+V[g]#QO^KKH7BOZTAHQZ0Y>-4
RQ#?_@7eMTe2R;/,;TLFQ@HC#CUIgH8HG&d/-5gX3#_>5MG<A]/Y)g&f9_IcKC3W
b(+BPU[VS/<fV@>P.c/LEN+Z]b-:K.5.<E8=,LM=.4SQRIEfEII&.N.-WY14WB]T
a-;:3(9a&L/eD]G@==QD8G9#V9T?DDKH7G,J-[1Gc.F?WJ7/WIFLeA+(M)E,H&B4
cg-GX+6S0Q@VPfY?RBR#,2LFe#K@4TS8@KOG+14>#7)<9;LU;@&LN2W_BK8^a781
,eS4G0L5cZg.7)F,dcG;ZUWb?3]:T-HaE-8:T.[[g-f7IdKAHX.c/C=#I<NfBJ48
T2aA]L+2EI0a6ad628ZT5EERbR0Id>M:,\a(G-W//aKgSKO)dWVT<@EcB9:6:632
]X/5+Ig9(R_-?26&d]I.J:=UIbZdcFU8fJ><5A<0,3A<8VC)ac,2_d=ZK[8WePfV
U?&a(T.TY2S0Gd[G5f)^b<4YKO;=e_M2:Q865)<LE_3:FaP82^N2>@MeF^V<GCf5
._6dZDHM_.H_E8C6U.&4KF(QJT^O2TZ8a1cL72AQ.?[D2]NF7[FLB/K-JTZaM-0Z
MX-+#5#?^OJ-ZJ=eAPHQ+(.AB0,V3(f+MT.:F.c_dS?.7H1bb\UB>Ug#S9b+0(Yd
P6#1A).f)&:L//aPUD#DJR1<0EBf6b,0R(4<bYYJc8FQT;YYC0,F[B8?9YZ9G7OO
f4&gBN]A<5@^.9QRcJ8@c+fOBIV^3dF(BI]CX5I@5A^RddV1:D&-B>?LE)a5AD?X
JNf8[cK?0Y@IZ>fD4GRc,f2#KI?T;^Z<Z]dP+2NC:Oe4.<]R3gV?fOgGY69N1?Wd
@Odg4ac-_GR>7:^96Xb_B;aFWD-3@W-5LLP76SD<N>C2G<7]e8#g?[J^]b<PK8G;
78#?dCFI_6\E(#TI4\J<QXO/>MGe+fZ))5I)Y(,D6\VaWMADUdU-Cdb.feX__QE2
FSG-I/4Y.G3=K9>FSRBRGd]E--9A\=\LY^1U,^FTP#EF[O-04->==??&3&<\aYQT
O[cV_;8IVXTgJ)ZRHQH0^NBcZDI5[Aa8OF9cG^0EXBMaU7GP)S81[JX8)0b2]3[K
>0A-SQ:A>Gf_ZD@R#J(N.-PT(@HC,5<CB9M8^g??Mb)bGe&WZg86aBR_F/1fbP_-
ZJYPaP3;J?KHZQ-X9#WMdR\KX_dB.2U[I2EZPJ<f86D5_;ZG/02dIZ=dV5.EVNU1
[<>gaZLBB_:(YWI+-dFWK#K+HD>G3_\QTMd0O3^P??#]c@PB)c;9E#@WIMCf1T83
(PT0]1&GYO9ZbQAUJg3E=HbYIdTHcMS1CD1J;AeC6X@UQD&_,S7(><;H4>A3]@AW
Tb]@N.HX5,6#U[4@+(P#^@1[/R]>Kf.PG/EUd(Mc;KT?]>(OLKEagD^[B9A+WR8/
\&LXd+eH03^R1Y38])I&21.US0Vg=.U6\L463Qgb4Sg:R59/PRNCM,&Td^YUG]Q=
.c0eWVC</ZZ,;8e4OB@.7=&.[1A=Q,?V9HUW9.I,]NT[dc3Z5;10AZ@e(K&&:#fU
?XZ1Q1LZN#QT(IDF/>._^6cM;,/b.Q0F40@Y4WQP0M9\\)8?_E(Bd/;<fG(1,D;&
PaP&S2=&I9RbAXLFR7#H4JHe]Q((f(UM92KVdJ+BI+fKg57^6[]g&ZVO\bA@VbK8
E]SR-MM@Tc;>[6<^ORD,(aU/)/]OfZ5fMF+DP6]d<9-I8SM;/D8H,C<+KfIfG9BU
a5A/bIU.\_^Q/Z>c\(20:::)4g&G8K=Tg+13=QdJFZ:H4SJEAZ/Y/GM,SaZ0XHM+
<:><ABfFE;Q.DHa]:RT7W1?Ve_\B,O0;8UCH588=^f5<VG^,XL3&YYZ[D[L98PeQ
\SL?&5ZF6X\M3CRK\NX2MN507?G=6/[VLKU[QE6baD+(/[?=b028G:?eM:dd/C?3
+H=)T.RBcbc-I5F1VXfUCX//DaH@=dT0M4LF.&XgF,<EZ>\V&FB&L)E6;#dF@5-7
[XgHeEbFcTg0bHJ/ab/e^1ESYC&e#LgH86Tb&25PBM=:1D7Q58,[\.V3AA8,@(Zb
&(ZU+](4P9)CCFR[:YYX../9V)dg0X.NWacZ48HZ.@1aJ)@ALYW3WO@TP7Z)1<SA
L,D3Z^:A7#3CESH76Y.STeWW4L#J8XW)74L\Ac&?OUJPJeI&+ea1Q&Td2JKR;4O^
G#0Ed?K>;5aa=GRNX1TGWAXPTKVg^=c\O#BL+R<;)V2:[^+99M.B0KOg3P7RVNFf
fB3T-B\O=LIZ3#[5?=IV+PSOKe.RD+c4Ig4^NS@-;.Z<:M.OL8c2Dg=X^-V)Cc0c
bSDLE/]U/;>#X+?3_aMB(Z1/[f-+LSg(gD7G2OJ_A#XCbXIG+2P36HAODB?;]JO-
YG9NV(Jd=ZS/C.VXQ(SP2V];_/PT1YaYR>C;(=DQ4g;+1;B_]UdT3:K^QDQJgKM/
4V=MP/>15La)>O\23+H7\EA&AZ1)Ve^8.fZZHfGSQN)L9I[fADd9D4:^<^JH8_66
=EQT(,V1Qe2P)U;O7=3?HJ+S4,F9b](OaG;_98@SPA35^.-gZ]I,\4f2T7570/M;
:3O7O6T>+UPO,@?L?KXdIg-[5T:)VYeZCe[[2-YdBC8WW7\c94CR(ELA38gT[XZD
K=c/WJ-.H-F(H.V#<^6RbKW(=/QX_=I8a;+d]Q0aMB3O3DGR3MGYQf<]OL<7=.26
S_HVRB8H^^R(A_H;M)8Q0EIf+4VJ/AG&8c9\cBIJC=feXMF9F2EKH^a^2(9a7e7X
aA:cL,ORcXJR0=[.F@;N[>g#2HEU6F9_Y1f1?Wf94/cYdN9^L2Q?.VZGcGO5P\E_
RPU_[DQ>P^/CRZ..LUd1T<+GdHI-11g/aE^<a._af=P66\?Xeb-V4A)I/c)>+#g_
+=<;95?W&Yb9?Zc,RWc:VR/FEQ^YW:G)H4Z3)5f\U7A\=V:3-,OUSBEQNIcXA?[B
M5c-/dBBV++UC#XHDg/&dGER6?QWD-4G1]Z.;VaU\79V7+314#ZI4Kd8TMB^231H
1.13-<&5.0XWU.9@:2;A#+7<DX\cC/>X;dXaf&c7NV@>7U)0BA6BDfZ;R5^2\N+4
I;7]RY2g;[R,d;SP40-[&KeLA]L&SEI_?@2;B:e;:K;6U:#,FT5435X)]_.>gPA6
PS>dK^ZMKZaO0J?1b8]-8;X#A3Zf6[I-@/A1_;G?,7@ZCCgD9E:RK,]A)+MPZaAc
\g;Oa/QS?OgW7PgMHb_1E,[&aMRf=UX<@Y+X\23a+\^^XUFENKXF?H81C3P1FA)5
de+6eZ<W4DFW9399-KL1E\e+AK#YfFHg?>7[[Y.7QA<&&;H0VT.ECQ:VA:5FE,0F
7T2:\DK@Y0PMYaR,2(IU?B:M:KIZ1-Xe6H#;0WJXL@,?OIEY,=ag9V2#H^D.]/D0
(,0JHWe\W[/UUeB-eDaY;7WKeC.W(E<T\KQY2JQU^EVRdY<ZJ,+6ZI4Q.P;9+e=S
W+cI>OgfW+Wf7()-c4@0+)6FARPba#g=;^Y]f88/3bB:)[,GeP)N;eP.CBH=\SEQ
cH>69GYSQ^H-H8F]>J6X]?.>e.@0E5U70_QdYI<A,1<J]_e-48@@+^Y@R/\10X6;
L-8d5d\S1B2P4K@BS(D+^P=;YCT\VMOZ<GQVd8gORCZS4518]#TN5Y8&8H@Lb6(=
Y2I/;a-JH=VeZKN@ZeFDW.?(<_/#>\Y[H:(DdV/Tf]J,+S89L=?650VDDOec^E)(
(c)3_L=RdLX8X,a3@<Y>C@EG81I+>,JLXX>&bKL85gMO8V/BYP^>.G7+Q[V51cG\
;0_N]a0;5Ea/APDCZ@-]@I5Pc1Y79.^PEUcdd]HAeT4//3@.>^d0#WDJRV5(V#@[
.VYXX897035_\5DHg:=J[?2&?;\GY6LB2A1UBL5c7,aYBe,-dRe:cb@dZQPGef]E
VQQAP[+0e;V,1CX2dE\2@Q8]RHRZ=gG\U68fQE&N@G#=\cXZ.D.6#II)BK7Y@C&a
:TG@<-OE5XO[Y[,Sd8,YYDf:HbEDC9-P)C;0^Vgd@bEGS1.f@;9^DT.W;1;^aY;5
6Xc[U(8Z2/ACT0]VWc?0VLd<+UTMF=fD1XZHW_9XXKW]?YUFQIdG^FLd:=?_7\+=
@J^(;=#0^Y[\/<<O1_:(J,Q?:NRL?.=LXg93_Wb/FQ2RZH;V:)8C@0:EIZcRKA,A
>6&^F+=Y.6)Q4c-;9Y[8RJ(;G<SRF:G7C1DA#,2Y+C-6bCdH1T+3HA#NBd0S8B@]
3+ER^9]^_D/EgL1/dG))<P@07YQ8+A)SX,LV.:8gKf_HKE51b4I7g(SaRDE^>aV-
75L/C8Y8c;3(Y.X.,P,c9DbC&]BTHHPX\(^>XaDP-FRP+<?OgfSX4DeQd[>4[@MX
9LI.HZaUG(U^@ZBY4?2\Z/L1/bWBIR(S=\Q.99[H\.6(Hba8(T:c@:710O=3X6D^
XQQ63[L6>Y,YN6cTM.U0KUW<=b-2^&:GY.;]J)8Z^0_Q[+(30g&5\1^@^[DP^dag
LV[<[ILS0+2-;IC?4);10e?1P7A2[3^1.(QJ/>;Ta6NB)U+WIQ,ZF2)SNdY7SBg2
a\KdL2He/S+++8:&ZL,Z.81d0a-QS\+d]GS&M4+MGE#Y][P(4([NR0dQ^[2(.,G=
01ZTcbe[Y@(113;45XW)<ZdFeWY/0:I9,EE5T/@-+Y#TI8=,E];^.G2S,R(RJCGA
gC4edV#O;>[YZ-@EMSN#Z3NZJ=MJ]5cVT1&@]#19XEWH4J62[R4A6YN&1SK^1L5,
He.A>0GO4ADI4/L2];g0W^Je\aGAZLLX>bSRB<LL(-\egXa]1.KCI^+\V;N>B#+d
JO\-D.KbXJS&0:Q&2K,+D79ePbdS76)==UTC8M+P29W#T[IGPIFP4OLfPFN@]J):
63:+-,Q@W4CJb?4&5f(X,C^2_J1cMQ.CZ45>WT3TQY3V<J;BQ=,8YLR1[)//Ya[/
6b;):PQS[EA06[ACWDC:f+/ZPb)9^WO=W@^A-d[[9Z=PWbVBT\EUJf@L(b#T>8[=
VOc&-:\da?>8M-M_Vb1eYe:,39DWV?GD0TQ--A,VX??aRC4&:6]I3d;P5XVPeLI&
Zba;A</AO<geU70^N3FK6a<T),.F_RZXHV@e(e3WC,E(4L/AIH_H-Q,8\BUd5,/#
^<P3)I2Ac1#6\;#S-d(9?_b-_[^AFSMEQc2Af9(@P1\ZJgc[>c]HJ@1S,)X>FPa9
3Z-_9,0^eQTG:C@/SYWg?A=>aT-L+_cHNNO+_)AS,FBSLggM2N8gQ9MeM317<<,K
H&2d9]d^A7HgK@[A<[SdON(4.S2?\S0+TDDWR4M=7PV26JZC?9e]c3[Q5WY,7#,6
)X0O_f\8IJ/]fe[^U2/#JY#:#HB)cd88g2ecX)-=ZUHUF6>S8RHcX.E[PM]=O]4K
=BABBO9T5eP.e;XD(;WR\\GUDggU\/b49bf;MJ0/a1<TG7^?M>D9@]-fg)B@7866
8.(8-7HM::NZ7AZ6#dg3/5+ZQ[.AQ6/M6]Y#c?eVE>&)-gDXZ<N5ZM>Q5edW4MM@
NeB9d06a6YT&6XK>D165^--(T]1-Pc_)I\;<M+;2DK^gW3WY(8=5>Y1,Y(7;M.)/
HO6AN=cCaH+86b(YKUgg_55_G-8]NRNa7,F)6_7/\]f3cZ>c<V\XX<&;gDIbLA[d
?^I5==)0A>[Cd[^cE#/-=V8MT1Mb8JV:cM9VGV(W]\+<#H)T@A=g2a>:SC;=5f)^
HDeWSg9HWS&<a3,g(-6Y=]1Eb)T9GT5[^G]J3G^;fP0I>UaXe2-8AcTg:;VS9&X?
U<;O;F2Ic;YVU#)95dEDfbV]BGO(;Y0F,#P(L2QTC7:dZWU69E--,[OeQ?T(Of.g
Z4SGFd>S\IcbK4)G.\&ATfSL<-?IbFR.TBa7:c_AgIAE2[EQB8;W\5&d_7T80,d)
,d9HVe=Z916CIN#F^WF\>T:,)(CfBB+RZOE4c504751<KKFYAKfZF96J==,)27H:
FJGbU(ZO^FK5/2D:N=?:Z+LeS,2;^4EE#N>JaTDF@(8E<5?5=TLQ9#+c_@9;A:1U
3SPaA6g)-)<3U/VcWZ2MKRC.BD=(WNNI_0ZM?U3ZM3\>FJ,=1_B30,@7KC^eCW@T
D?[56SD+Q.e(UO06b_DJV#V]WbMNK^AgfG#Z6IaAO3/CNJEa3,f5386;=/=dVJZ]
BaZQ#cAPQg0KM8-JP\fT.8X4bM)(K43PJSb(VQ(#B#S@I(^750_&17a.2]F1g2cW
5S@fTL<WeS+GQ1.O+d8^L_^3X_.[Od&/geZ/:Mfg[\[^^e_ALCBN&cD>Y.^dIEFD
Xf_PgC?>,8_C1X@OA324,SLGXce&C^XB_.W(;;;+9gOS//N^BZgYC-gYNY[C/:>K
304N28\W9VId7Ue<E_C3IDX2_SICYEYZ;V0^F;?>8UY<;0L.BTFN(;+R^9E+UQ7e
W?A;(OYBQH<1fL1cM0=4g/YfZ[L3AaXe.RA]->B&Y>MLIN.FD4@O,;5V&/KgT8O_
&^OB/9<H\&3VDPYaE\a\b>c?.J0=?[\_^3&E0Bcg<9F61VdVC7:I(Hf-MQ&1_EYD
fX)0gSB)/40g\+cLTQA\fZf1P]#E:R0>6L9],V9Z:X<&WDg/]E]6K-WCbd+(K0KK
0^C)O[<IDfWAO;[=]Y.R]c-;MMB+@=NQ<CN&7a3f9#ZEUROV4;J\Fe+e8?Fa?7Ec
1?,HGJSXgAIP)gC,Q&,)U]b&O(IE5--_8?H3:K:2)=^UN?23UP==[N9X=9B4#_:)
[9L#,I,bb3V3-YUT2HIX9=WW@_])C_GbH?<_8bBV7]]V;7@V^/+>d),RO[1^7R-X
\_@[3]E-Je7^4?+_XC6>9gJW&R(;cQ9NSdWH8HTA\(00:ZM1,.MRGf?BM2B?):0(
63OO+.I2IV];\,0Q&\>Yb@-d=..HbK(Ge#T;>6cQEfP)K(OXG#LS.HYY[EQPFEG7
WJee6+B/1_(,BI.3ZWRaKc9ZE<67I^[bPT+2b=W))[J6^&JHa]UV7JA(70).EaQF
,6@W?VX&CNE4Y^I88YggG7JMIBI#e3;g<=.R2H],QL@9]6EcMW0R1A^4I[TQWdTU
2bcJ^gGC-Y9UcRZ7#8gL?7;K+Z8032FQLS;^f(C,L+DOJeCFA>TDdN604-Z3^4_:
#(TY>MgbI<eLM@7gO(KKEb;<5fLa0L5P@90P5VC[;NgS_MX7-OKbA@=6JUFcH[G&
fKaDMDS19^T&1:RN/cQH,Q_?8X/A;Z_IWPK^L/c99GVM:4QC)EDD5&=&SM,K]LJM
T0Pc>)33Te[b)>L[OHc<;N2G,\L78M>Pg3RKgPSKN.aKS6V,(BPKCFM5dbJP@=WB
D[<?,;[&P:[>4c31#/@\^J:;H;_.MGI6_RJ;)K]7&B3+1RFbER+-dS7NXWTd^^0N
-]F<X;SAFT2NJZQ6]-#<@B>fS0U6?VEE<XUT79bcF<U&ea;NQV<?@ZS>&O)ZeN\0
O\S[bQ4e[d=)&e1K)T?Ig/SdU\W[87cK=bH>_eb6M7O_</LCP(E>)eVd99E:bX5-
RTg4MCC[Re/G/;U-AP5VO0LL;W+)12#\T[\<\-2=WRM78Pe+5N9BW-G2Pe<SRQ(^
61[S=F3/6f8SdN/+YP2TYJ0ILDUQNMD>FPU+g]-VRKWS[ZP@XV49B6-CW;dcdG88
R]S=;C8P#E3Tg5_/.1_@Wb98L1FN@bM0EH3EbeM8[LW[U@fbaD^ST3NOZNXC]2f[
FK&7;1>?Hba6#TGVI[11EG;Q-T,#-gP]?-1YGaUQ;72:.YMeT)J^C.-B(2Z?dY1H
1aHHXVAee.[_,V>S3d]bg<I1D)OCXZ)?cXL@HJcIG,8aBa0QDX&g#AK1AA<d?6(<
d:d+BW@Y,D;V8d,]KW<0f)3P4d6_.-4\F<We<1_dV.BSYUaX.CMO7EYJSGf>(VQO
>DJSMLQ>4bGdH\TRX-f^036ER5;/f3((>/6+C1V\H5aI;4]QTWJ.&M,]LN0/a+gg
Zb3=R,.[>SA1&X#=P^8L)G=Q2,KfYUISYUZE3I^IRWL3F34D7UGNgd)D0&bBI#((
-TIZNK&bRU3:#E;BS3+g]g@T#FPVXZON_&eK&aK5/>^I<g/K^d-a1QMPKgL1LYI(
f::4O97>QeXG8CI+\XNcF0E\:)O.cQ\bB1dN3><P94;N^dX/]3S<YdLR;dYI:CDf
QV9DY[FbDLg^Q:I[VU@O-B/Ge;AG1VF@2F3?NRTO=@@e2-6YdE>Z9XIOKVJWX>;\
&@/IH^SH?ZF1TOB2N2Q:#:4#>1G7.[IB_]_Y@c]7;)-46)F8ID-.>3JO(PB62AX3
1gC6>?CJ0IPH:[VNWZ+N3<[cR0\X#YP3VU&7O_T>E,&=@JKPH82VJ+L1]TBPDHZ_
Zf3U961D\L(-d3W+64HE0>b#.U>Y[.HZ+?+d/ZYc+N)3B+5Q43ATF\04>-c5/YQ>
O/IG(3+1Q\PgX[Ff;<f;/a&TMa2#FY:AC,/X?Q3V?U9Dc,]K8.JQV[c28UJaS4V8
)e.&\B;:CLOA/KRAfK<HdS)6^;@1R:GHa<GPJ?]Q(8CQc>Rgg:=GQY4cO#?BP=2+
K-?B^F&)H40HV<@AfJ[_AO:[c&C1N#f;?Rf;e_]:RX3Lb#]W[9KHPHAHAb7eL]JZ
#UH>5Xa9Jcdb=S].Z?/:)<T3PF5KV+a1aS)XgGP]M:Ef4PB#].5adAEgaK]RR>8=
-K>fW?aVUgWCA:\(NA)fS>?,e6L<)]J-+8_+SO_LT/KD(cQ]SH#?Z&-([/B5V5UP
e0(855aS2MFHH8cDG,cc^8=@&IK+WR0&NQYB^(,a.S[;NN[NC7(RH1?;K6>.BX1?
g9-+@bXC,CO^B/]7bCI8T7VaH\SH74@0:./+/Cd,L5;XQ6B<47Y\&e+M+Z<DV,,J
TG<QU;]?@^Y&D/<gU/#Y:NPaX[AK9]5CB(3T]8bRAgDWIXZfWIa[TVXN&+(bSL?0
ALf]W5Y^&9]=;=WHVc\T)]<ScK+=_02:Q7+>S.+9==,>4WE+#@Vg9W+A\?NK<9eb
,9?248^c=:J5QA)A&f@LCPb>B-V6g:00>=8E?ecBX_<)cA)T^gNbN5;D(J=b0.12
a>P[@RMY=<T7d1^?IV0?-e[((6,N^AaZ&622fQ/<V9Ed#P2LNd\8HH;FcgFaED5I
2MV+,Y:;cV>MJaH[=&eW,.G_Y=HXZSIR4S&3GF=G,:V8MdDW3W.)?_c0LaC2_\dD
:1O4_4X:2S2a1bC<AbIJAWc3C)U<245_7=JPZ@AN8>ML,FE^)Y6^7<>]]:1dOU^f
_PL&)e4WU1>eLEdX&.7[8:X]E=Z/E6;D;6L&[CUfSUa_&.2UQLU,#)gVT^32_fdg
]QY[3YQQ+ea&ega/LI0dM,909?FDRUW]++[V+?Yg..f8>3_d99RY.OQV>4-+Ua@X
DISQ>/F_LLPC5/I=>2<8JF6^FaT-5Q(^I786ASA,8B=_+V<W//JVL]T8]^04,e7C
_R+^?),^eM>][&-YPN7dDRB?.@FBDcR)^?J:L06VC7R+NI:Ze/+RS9T4:0B-CL+-
JPb<#0AgIY6)P[P6T::RBd-25Mc4:,a7,f6Q5L1UB_DYWd]>S2+<]RK<)^F]L82J
\/30c720;/U?V;X99fIZB2BOH<fC?[+O;B>&_;+4L-;9^GF&Z0+5R5PR(5&9TR/g
+N;QMb.\&-S+D\\P-YRT5&e-=CB(69PVG4;<FD0>;&\&0?H,_.P#1@+Y_@a3DR08
RP_#QSe)RJ_eESG),F9\Z8&V^P_6P,W2@)91eFN4<@4bK\E-c:?6?+3aJOdWgKQ.
@[TBYaSbaG8V\2.N8f>>2e)b>aJgX,-G/?c0f\e7UDS7,A-;=.U<_]Y=C9VeReJ6
WZV+gUO-_cf=Q;5VA^(,&aH.951L9CAT]/W0HXV.97bfgCdRV>UEH8GHBZS^Kc?Z
-6Kd07b6+[#PG/,,5J5U>Cd)1;+b?Y7C1KJ8]e8\K=>]=GTL[eW9#^/=_TK3;BS[
>YMI=D,3gX.I@d9]#K&AZ7A@)3Y>Y<1eM[A\PAE9O([;7,7<K>g=\38T=7?LF=L/
bBXH(7U+OTYC)adNM&X>.F_Q]@b;5<(RG>]XTI6]BaT1XM,/_4/F&37E3d>cB]DD
P3=\b@/N]e-\P.EP5(fT&E4Ob51O<D_C:Q9&YM7a^-AcWB=fQ2CX0S\,17g8Wd8P
:cG0>^0HbABMKcUAA5+.OcUKH20f0?EdN#&/Y,HUB)T84A;CL]?AfQC)_/TL7+cX
16/TN^5J.S2c)8?4SgSBC-#63)&9,Q:FGA5EED^AB/b9_4g\dYO8BTJ/E+:MdYV3
(O7U7@0>Q1HQ@?e0WAaD1C&1aeS87+g1?N@VU/PC;0JWG1YdO:WWNC;35;<CT#M-
g;2UW_WK/UCSO0:/E8Pg+:=F4<.)0c,WUX#5KgQX3;eU=7[QT:4\0T:2BE5+f,A;
,MR;8#Yf/+fA[(-&H>6Zg_8X=>#^^^@,LK>08L)1\^6S/7F^/&DL?KXa;bGM]4:4
^O+S:]Wc=.D>7HMZC.3WRb(gX-P#T3UR:-:DNcLT7/Y-^Q8(Y<a_/(^XbT3LBJ3c
,-_HYc(U9@-(QbD?OY4BD\A/G_6PCc5[8g9#>R[cS;d4bWGH>c1_0E0;3d(QU:L=
#+/T2FGL0^gX<S+Cb8@GQ<eJ7=>6bX]M7LOT(+fIMWbI?@S1Mc9\;9YNO_8#@\>E
)_V[e@Q[7bWQG5fdV#).d3:F<PP+NKgRTH#->R:ENg)Z;TGZ5d-bNBc(C^GZ<\#0
IH(a.@eX>DGRa=J@H4A@DMNc>M67\VUe70-6_I[_2a#c-S1>W#c<G0X=>LX=JBeW
DZ,bBAC#<2#VZL75B=HN/9S6L,FI:_W-0=3JM4R\@E9U+@?S><>=-5P7M=RQCeML
.Y=P31^<GNUd6gDO/GHM8ZD9U7F6?>CQMF<^8;F(bdHAS&IHc/K;&Ja-#L>FMMC1
ZO._JgaE[?b)]_HQ3X)&G##\D>-eDW.4&#E9dYI#RK9FcSW9W(9&0:2?a.X,1KE&
Y:?P659=PPW.:^6O;5U@S\4X_^7<?>,B.T\@+J?UVDDdQ?eMJaGO_9=A11B^2S]F
HJXHVBK:XLDWg/5ZVL,(RPe/#gaG?Ub)N:TKS-L/GKRfc7Y1>,HB1e75e+X)AUFS
8NNVPbQf#9:V86f#=L9_Rdc01e(>b1cS>/DPLg)&+)O97U<N(BL:?_GSTVNGXUDF
=1:/W0>#D[=QJ?T&3(82B;BdE>d))dT=R^.1UA:QcSZR]#/U(I@fX3648Z&AB)8@
@3M>H1<QaQGG1W[Q:/SW#?7:SU2;]A-MQP:PY-I=S,>E08=T.,8&fATH<2)59._J
g(9a>CMVOFa3=.f(YFM^19SP.NX,0dYZIO-O5FYQ,TL]dReC4FICeK]d<Xc.ETYT
XW1J4_HDM6Ie\#c0V3g/EB,H>AI?NNGVL\L^.=UC#ZZAGM(IF,GS68H7>M=^UNE,
\EOfXU@.-b^C.X[A^72^>2HSZG?OeY9U#O5^??Waba>P5U4d4)JOE_CPXA4[b,b(
/a_25J<U(g&L,#KKg.(bY_<B2K:G__WRP1R\4VIRHEHMd\^Q<L?eC+bMcTVK^2C^
(PAZ3URY7P;ATJ&b[^YN2-F=V[\=[WF8;Xd8H8WXM>F(4_/K??GDNPd#-#-=TQ+,
0CB.G3c6PAF9KY1YRO&AC+[D@0>KIQ+>1?FLF.7([@>aQf]YH>4A@=^W.@M2f;AL
^2I>(OA:BKdAg+A.cI95?<[MIb6;[6DX6#A?O=G_+/[2MM(f415V84#;d<(5(#QQ
M_P\-6WXY2BY66DG9HV4&=R>E&=7.W7(,E9M#1c2CcP?##<#F&J?2(4Eb@5R1#UU
8);#d:-Z:MD)1:=59Yc.>_B=R^&F11<W7+0>D4g\DZ(_;e?V0V)[H\>aX#U^F3(.
C7U1E)a<5<5@+Ze[;N0-:;Me8QBEH=+0KDIUP@V49dVDJW81UL&c/c6d+WeB#\N[
JM_T_d>G;5K(Rf0T,B=f#P3()BafBMI+ZE^LO/T:4Z].BX^((ZU[Q[XN#YBGPYIZ
e^F<8-;G.HAN>JBYf,5D&b8B1BM/10,NQ2.O/1XNBeRBJ(\:/Cd>V?SC90c\F5<I
XgcPOL7e_9g9+Hd^7BNLM9JGX=e?W@P>)fc<e[]X\FL46ATH7^<9g8EgM38A8BP=
B>4I2\_22>=4=^>UL+F0B:>:&U26^_;R_9[@BQJHdg:MX1]WJYZ0#4^SH^,EV9LE
D_\dWV.P]79beLPJ#UV)/58g2cK[H^6Z5<bP)<XQ4C-TB1,7V[fGD+8&:4g40N;D
=+7>,N1@=4BT]L61.Sd^E=Ia?[ZO;#VFUeODT>@X4T14,QBCGOUE8)WFC^CFBO]?
=V>[1=b[0FIcVWI^=#E&\CGNc:L(YZg(H2:f?.Sc5/B#H#5cO9IB()5((&ebS/Bf
7ROTUARZU;eV^D@>>B0YcKMLKD@FWJS]/,J\VMM+/&VR_/[KTf;(5dX1L(1^H);Z
dSG).PBN^P50gaM.a,.2]X]@Ob:5VIQ2.<9dP)WARXV(B\1bdWGL49/43#cgSf)K
_00F2]B/S)__M1^./XJ)?=g?T-^C/3Rf9ZLM]Z,88bN<ER=WL@UIg:f>Y_CKR9RA
F4@OR?([O,NS1B38,S\\GXI##JG2+V:3Xd0A:=&Cd(25>6Q])F/+67]c-UACfVb\
R(V]))[V8&gC[;J\VQNC:4e.E:9RXWJc^LR)T^==4#FRE(G_S+ZB=UGd;7>d)W,4
Wa?>6?Y)?OT4&-QL5@,?_0U^__ENO5,)>R:;Y2:EM9#XFY82\OW4XP<A-)E3IgLS
=PI0YN)&3C+AYK>:XH:Y1C7B]4^VES3G9\AQg]AU\^\c.<\<Q6_R.b,U?@AR&_W@
Eg).]]:@fL\[dYKg2aFNYc/+Kf,d>GQGNOS2]4)_@X&GN95Ta2].5f4X)87\<QW^
S#1D:/([a>ZZV0M+HaOKPL)d[ZM65/5EPA3\6?#OWVV(0<PaYMR977^/ECA<^JcJ
F=JPQ8_F&2.,-]8A[fa9L7B&ILR/K8gQV&,],QJ@EI<[)N9cL_IJJZg407PZSQ\9
XGUM09RJ).)GaNMC_>25^#8CdJ_>;bW1-J8Q<)_BJ45JfLIQRf?c6Y6(T#<GR7#d
./:QF[e;5-d,9W6H<VW?X:@4,JPcf(IR#A(9KDfcWf0+4X:G@JXgEE-8:^,((R,F
JcZJHY2bVBg^IdXT23/8GNV5<F(dADeC\LZAX-;YfaY7?dNM<McdOT\5BO5ageS,
GP.]<Q<Xb7YE3aGA;M;XV[UcU)#,G;#-0/_9(1bQT,UF=P33>FM-I-_R?22H,aK^
^2^Q5RC[bb/MG\g/:S86VR#.HZa_/\M6Z.ACM@=c5YHM,6.DaS(^c@DcWGEWLQ83
JPPG>Wg2NJcQg[\DX[4>HG?GGBd0P1g\C#(^c/dfF_1A902]Wa#:-;1IV<W@L@&b
eQI?)@^XG0#BJ1@FaAJg4^VQ.WagN&M:Hf).RbJdPR2b+,K.X[Na]&T>:89WJ>S9
QRSC]/L?9M9</0GdRVBB>)R6H-,O1GJ/9G1(Rg?5ETDd:B6CV#DLGbR)WRNT-I23
g6UIWV#HJA+:[@K/D=a#YHK^PH<+MDO7[C5<;LgfD31e1C\[+#A-;>://O4UE[fD
Za[e+<XYETUOUAZB[3)NeJN2LE:N/L\[U[):D;R3Q)+:G/.GR0A8Q#3PEeBI&GWf
@=D8UWSP.f5Lc;NS(;QX#\,M16E@/KgRS>EFF^V18UcJAP80LNUe3bMIGM\aTO4:
PE&Z/JAER,CYdS^^<_[;(F42WL4)XS&J9;&,4^K7^d79OH79Z>^7AREEA+-H5Gc5
09]\QfA[/###OE&GGbY0K,::NV)_&&;CE4.MDETO^7^<aMAU@V[P6b+eXaZC3P/b
SFZ>?=E:E44LDZA,XSeZ,;/OTLZ)=H2&N-4F@aC#1f<V8CbFLe;1J,2F3L6=#AF>
0O3gGDbdF4F.G6KJL:B,Z6Ne]_XJ#dWL)WI18+g?P/Acb7\&d;#9VF;QcaE\.3O,
L3KZM_9bI?<2.2Q+;J8HfP/@7O;B.d07N0>SI@d4&daIdZc2fEB6D;R8;3W&A5dH
:b@C46Ae\I,UWcA5LK]e_E[>ZGGQXfX0EZP(U=8:<Xb>1dM]AA_V3@=L=4GHEY8-
(:/(d:c#/>2?3J@Q(X-DFe?6>eYd1dOVb&W591R]--0cH\E307K04\MF:VC&gPQ7
#WG?eA@bPX<#OK(QBO)b)D+@&.fIC=#f)>b1&GPD;c]5VJ=H\0^F@>cB@O./VWB<
<+TIcV\]69>cOS##8KZ.^fF-;6S,H<HeP=&9706fM0GA:>VF<E(1,;Ua)WQACFK8
,R\8<VYePKOEBPfOWZ3Y::RB5O<MZI168,O7:S<AA+YUURM8^C6/<.71,@MG_80S
MdL.P9#/79d]2BQ]aAI35I@D.&MTHRV[>&\50Y9<];LS4D7NI]#N8;,\I&;<&aTO
RcAePV@Qg@d3Z/4gdD?HD[KUVI=X)940NGA@1c&e07_[Z1JVNdYcbJ[L/J3?B4G/
fY??NM3ML-d\P3EEIJ[6Lb/VD]2Ncb3C_SHIPE:eC0&[G=E^a(.A60ZdP<N1?N-G
Yf/^&Y;eKV1+B[X]/T#TGU(ZSdb,1?.GM=/TIJ)>]=gN;-LaF)CFJ,QeM/HW\bZ/
>65#WBRZASIOA_ADJB8&W=cBMC6I;1DWOJff3+Q]205bDW]\d@GCVUG9/eY@abUa
H)EgXBPOSI1B8PEJKgWJ2S<>U-;N<1>W/2(4K;-0>D+Eb2B?NW^-?6<ZC:)]M1Z\
BGP.0P&O)1MQb<@=2CSX;3eR__.[IA3U@A<[a6P]JC==PW-6DQW4?g,.U+5&DX=Q
g04gL@<3+I66O8;eP[g96PK:XSYfeR&9HXK\[P/PWT3(dZP\/WCH4X@[gg+IRgJQ
MF&NdJR-<EB85Z<C0Vg#2,JQ-[QE^D-55058S+;O03\.W,-1W>2O.J_G&I(B.Ea]
5@@R=.KH1;MN7I<6@+TH<[a^Y(JC(gUBF8#KD;J24]\R=Z5g>/3Z)@1_FJ\GLJ16
GGKb)67-1Z@d57Fc?+f@MW[UDS@Z0TdVeW63Y)8F](0PRc2Q5Q[Y/=?:YH32SP<c
DYFT2118/0[^,EIJd>)1K6>@DeFU.DPYcee2@E)OB=JcVgP@ZN,W,W-@Q9PJCVN7
^ZL+XNN_.D&ZU\A@]aJJ&VY?>79:I1JI)>ZQeHYK/.Cfa]\#WOUcUJ8__<2M\1-1
5&c5GXMd:[56P>.=,W5R9R,=ad8#g\5AXZ=P294GOC6[PUW-Y^W>AXZ[TQ?C0@Gc
)^,((XMe&:Z.A>]YKN9MGdOG?\])T1NddX&LdWY&;\bWb&:+=gX+GLBAX/M=9_e2
]B-;W=,@(E_JYRA<A-(28fBGSS+&C:.SKS[GV55d)NCY[4DQDeO1^@D[6M^QWf^g
bF,J-Pc9&JQ;5Fd37<=YdI3H=?G4SWUA-7:RbI+O5.3)U^\9UWT))4QOA6_U.:4^
.=+X2(]]>HT=_QKWFG7TEcK?^6G7CO#d#R?J.E>1V8]C(;fgb#DbRC8O.6Jdf1^T
3F.3_4b_VV;#/4_-aGa.8\H\/&:_BM<&<]-[0D3-e5Z6,>]PT8\#(g22TPO9BTBf
/9G#>0.NEJ]92&8\^QE_B#63SI1ROA<_d/?3O#YC#Q<#QXF\T\4)QI+\ggCF5/P&
d>MEK+H&fC?g++49O^(bVJ;#&M-BP2_f_@CFPfMQ::PE7c:dY=fO?K?4DYb;VCWg
^GN+8]1Y#Y6+f.^73cAM1W:0]EGe[QN5XA6IUUJ3X<:D5CV08XL)e:,<9d6VK+=,
8KCS]W4B83I[N;251bX#GV79ZeIWQ\N;_4+JBX]+f/K0&T0V3f>3#dN_@-QYU@R7
BZAc=dOf/PE[/O;ZA0PfcC9>#V1b\@(@f1#Q7<84@aM,Rg,(>(GP.4.;H@QG/=-5
+Y_#c/.XHVKFN57<2M4Ig?aO/X_fTK-[PfT(1RDB3IJ2?b;(Y]6[We2d2.)8D@2I
bN+YeQL4L,WJU=:,UYOgC1VT2I(RD)UVZ^&<X5bZT..aT/.^.J)Q27@052G0a#3A
R@-CKbKc2RfO\9DU8gZ@4#DG40))fgJS+fKJ)(UY3db^d3b7C=P(2U73\L3ZZ77S
0<[BD[(</Y4,JANM;L2HTc1#?^I7LASK7_D84)ISVTOMK]Cb[Ab1J+3H@fAfU4<R
CBHFA2FPF/-DfGK9@:#f+CC3#MBfG4:8C)cgN.,bfB0]#MRK9J1P7V(B1aM((7Zd
-5Q//-F@Y9UZ6H,OR^MT+?#Y33IaS0GW/5c<W14R>X+-a1/RC;,RaO310;b(G\79
g.W=e\9#_cA;8;8,\A7)Vfb@J)a;9d:R5K^3\QLQX:;c3ZQQ/HHU34F-b[0Y&#_H
EEFJL9,YTbC)I=TOV4-eK,Nc.P14aFK3e@f&+^9>,a/I\X/918I8AGHFR],R2A4X
g9ZCg8G+JZ&9+.O:N<:?2dAc@0WM#BYJ6&ZQY-P;(fEg6gA.Ta?;]4=768_S]&AU
-4RC\;YWdC-EI6HL-A^<BZ^7G#^:]?N>4N&?@aB#_EOe],DI8BGTW#5,;,3OQ=\B
6=ST;gF9XG=QZ+ERdJX];?#^MIXU(b^>#(MP0Xd_BZ-Ba22\;H9]2F4W8L#Z=@Ff
_/@;Sf<#@.VZ[F]f45EG/Id4M]eJ3#\XR=R:8?<5@eS09H&A>\Ndd.EgCSS;X1c7
R10g@S[Fa/)..Y1HDC[^gMZ,cS.f@/;eeT+YU&Q]53FEVWKaA0ZaL>60Fg@-5Sc/
K;ASeSP\3.T4PD(L1)T>IFf,VO)(C@gc>0Y-Xd8-a2[dPdV,&@,[XD^<UdVG;Z3S
@;/4WD;/GEGU6Na.K:d?=(bPaW;RQ)A)^T).8;\ISKLcM<X2(&6gXR2A</db]##e
Q<P.,F6+A4QG[_<JWJYAI.OTe/B@UL\9O])bRP]=;FFUeWPW+SYFc]D\#1dO(A^@
JYbI46R9]ZHF,gF/BQeP3gB2ddJ#Z[I18Q+EZ:TT?0U2CJ9=JZD=NLV9+fC)--fA
g0BAB2F=fC#aSZTFe<E;]^EHM.+:QfS)[ZRB7.2&Q9].4b_<8AU8DbOR[_;W[)SQ
9Y)IUEaBL-MK)gPQ>Cd<bX?RB9H25dUHVY;FYD^b2P.=F+ZWR?@Lf:MJ)Q=9L&=Y
.)4)[QcM1O:Yf=2^CcGY)Ef3C&8gf/X4K3[_Ef)J64IMKDL7)7A4[\=9d.T.M[-/
\[4TJ0Q^(;;F@^1E5E8,RM:W9=T2<L;>+H[@a)IGaKMgHTDIXQ@43[VZ[G30>c5=
#G^:fa+&=79MbTWA]d67]FRb=f-3G/QV.W),H93>0e(ge(E>IBDRL\NLbBOb)e@6
Z@Qd#4QgV&/FIc1c7YfP.UYRPGSIW_,]M&(HBI,CJ>UFKg8a-[EA569+-<SS<[X;
@6]>NXJ1=;I;Va:)_@7,9AX+-\DVO=_2/26B?a0W_5U:a-06d8?#,@0K6Q@D-0-5
a<R4a0D?-Y<1?[KV@JY>P(R2ZF.6_YH)1C1V5-U-X+>-GfSQ0XL4X@cW^#FO;48L
N3,QGMN/<&X)b->f9(F#784(Q3YG7Y4KR5VVWIY,H7CCHL8..;@<?)VF=EQNa;3S
J]V[Ee7T?].;JKE;N+EOf]);5XBZ\QQ;S)ef+GZ=P=<2aA-?CVcE-cT+YQTOE9]/
CY9gZ=,J0J+D2HWe3aB[NGV]2VZ-BG:#WMC.EO<f6,KX9]^W>b8X@(?M#b]J:A@g
.&V-d\UI\-&2_R:WA8]LHa_7g\J7K@G^UacYTGX9WB[7[<M?#.<9SJPGY>;O1g:<
9e)N@75P\AN/\90O@;EITVFILe=ZU\8d=-P^gB9=<X7.[fW)&1F)KY10ab-J-Q+^
S<eYOACAIWaZfWPTP]H)\4V^a1ZP4TR0^#N7K3gd1;L=HG:HY&&3dE,bNDPL6L9-
@NX/4a:GB&A;TUd#-XU8+Rg=5TQZ2=M]g5B7Ja,LS:A03Z)OcX+.1g&BZT#=]B11
b+&MBWa<MWWKeKR#d:(NO.?T[S4HeIW<VaV97+HaF\B:/L#]H4;03<(J8+<+dYa[
b4&UP3G3PFEEJ/P3CEO@OQGQ-gG(UQg63baDOEPd_V#<(caKJLbE8)-G7;&0F/[\
D(M]Pe^#WGV(K=&Z=-H6X8g?84,M5&HO<G>7RNe\A/Vea<@J=(>/>(/Vc?;IZ=G:
LJTc1<,=d7=FS9-&.]\6_I.Da<&HK7)d#()O87?TM,SWeKdgO53EV0FQ^&e?@GC^
0bJLSfFQc:.].Q,#2MEa;6dG5J5J:,0ZWT?_GUC\\E:P6]dT4D4a.C&bcSV&QULa
Z#@((I/,@[7\R3=#&2?QKUG^_FW.0U9IRV5KS0+K?e<G-W_[\fdA5?HRYB3O0KXV
I(^AB7U&?Q,1HDPX>_4W:Z<MQEXDYa(dH&=Xc?6EJ+K[eZZYM[6E7JK^/SAX?Hf(
=;-L[Y8.KGUdC[7[U0e&C\R50bJc1=>(-??^UeL<<a7LD)SI.,:3Nb8<T:VQ/[WC
@^\R]/1d[&/=_3<EgeT2a;#ZR\](d/=eA;]3MAfZOg@CbH;_(-Lb8#3U90AXHUaN
KQHU:)K7(\Ce1^YF:GBS\?;eDC^KYNJg;YIa4M=;#U-X,4W^QHbe@J,1T7dBP1-3
c[B/LH1M-Ie://[fCbYaQ3\Z4E@UWd?Z@4)Yb<LaQH;PSa0MfeIAdg+.H:J7UKK/
JJXQ^V6=.c2E+fK&XAQHf7eYee(B(dKdO]Z]HXA136>.\0M>O32;&dYP6G\BG6Vf
[.F/@bR0TI)2OSKB1-gA+;I?-@Z#S#b&E^]8)EP]&+1^f;V[?\ZU6SXDIBR:EC/E
V0F+-HBAW:Kb<[KB>7,3#QCLDD;#(MOB24S,?2bAZM2C=52)/58S7#-YDC.\P.=c
5a_\Of0/K#7@RXO,FH3DUJOL>V-Z^fV\_Sc20]3c()g&Ib9?U.CQ]S85174[0b-L
UCE4X]D20c+1?-.<Q;F;0^AK5aGQg@LIE68b^H9)[(9Q#3;.#4^7Y@-?L]Fe^BOB
K379XO4]&/BdJ.FE^eGC=2FZbU+HCTQWI@9RDO0M:(U2_5D1]f_3]QY6[@Ha\e3L
LafWd(F\XRGL[X6,<@A&,=_7Q,Q:^FA.dC)4G(7+9a0G;]3XY5];3;JdF_H0fAg+
C]fEW83b200E.PCN,1/V-2.fAU?0P3V8A):\<NeFLME&gBWQ/27^X)E:6^S1g;5M
^KaJeP6A3)Z/e.=[-8P.9S23PdEICK^>9R<5T#I=6/6?aM5>Tb#==OL4.303ZJ<+
8Z_L=GX#9JYf56CfHSX\f6W@X>]R9:W:K66YPFdU212A^J-.=RH<0BR3PgMFFdMC
2.)X3Y.5[=^74>>DV2JK#>\W@=+Te5P-5Y#W^dWb6fY1dY1@UGB&O-dCA\X/W9d<
a/-#=bIC2\7Z^f+7McLXGgNLSI?3_KL;a+Q.e:BC5WOaBS)ZD9P/5M[4Q;-:8[DQ
Xa0QAUY)>OgOUR]_W:X\([3bc,9V@RXHHL++<b\FGVg:)N[eLR@2\gdO1fa]e_6P
6Y20-+4BN]_VXWK)HI0T;FW&23@eD81D+9eTH\g]^\-+<_C<C0A>D@A?PPT##<KI
67+#9Z@?QMH+]M31BS4_+773g;C\,.YRSKCX#d4\Q,dZ/AZ1Fe9WMK:+[T6&0NA;
/7T7.\4YK0cM6E:L;W[LEN/(b<@KWDIDLRg9#8<6P@/He_K,J[5^QXC:;C>J8;W-
TfNe\F)Z2-.BH+:6#/e,C>e(dFdYZ3K[&fE2.5f?HFD9ERO32>EPCL]QEX3XZgE0
>Z+;&-TXMSQF3V1AIL<6F9#3]-4YIgT_b?)YPc0G[K>V:8LfST:26+>;>2>V>cUZ
-4NT#Ub92ZHSfHeZ7/&e#RD946+F#TY>,86>e=aI7X@FK:3NWP.V:7#NV^Md01g)
7Q.9BC.->CefQZH[LRG[:2eA7ZQfT1XK9_JF.,51TG:?)2)]MCRG[P/1]DcCTR=X
N0783TP05:L((K/K(CC2=BI_]0W66IU>R_fUc;1c3dd?6cV_c6/R@R.4X,,5=+6^
GE8=+0=/,&:N:<.\Y;+dA++DU/HJU,5(9T(RdGGHH1TYAFY^=5cV:I=GJdUL/g@A
-HEI.VY8bPbgXA@(=bW=7GO>1cC.G6#(]C(Qe4e&OD2E]7e_CPZXU)RdFX3H/MPI
Ff.,BVLV^EfLfCA335TSeb<YQZKXZXG-bV+cZNS9)e+DJJ6V.#8W97_^OPf/gS^Q
MJ4<CMf&KR8],2Z+=2FNd3Y0<Gg3Db44&SQ1SADX<=&;<@eY2H>P#L0d?1g:1cAF
S+2>ZLLd@#YM7VEAI_6_ALCSab=.Z#E<=BOH./5UbM0JL(1VF-e]>P#AfYP(ff2_
Tc5SW73(H:+,CI86)CRF1<@D<:OS_15\XL@TN2\/,O:Q7+RZVGAa#PL=,ZIZ>2I]
]R2^f>#QecZNU[)&@XA9I,3@]H(0@7_E[bf?_35bb]>0K:A<O^3g2.UO=deZJ4RL
[MY&9^_Lf[AM-D?1g/7EbfP\8UGOGK058;a>,<c;@28H07Vb4dLY@0Z\cc&B=5#U
COF,UR.5M<?.fHPMg@P9@)N-3dW#:b5ZLMZ?)4GNX&Q9]&=eW]8I6&Hc9)P6\D(Q
9XAfI);,T-[)dQg^I:=-O(>O/[TN)PJ,La2O&9Q&aIaSVA_e.+ADXVBd;f,,]3G;
Y&QL<7<CIA5WHZ2KGb^7>:J^5L<d4\.KUX3bZ;6Zg1.:T[IXF)19(J\ODd()D>7P
I;83^LKf0?f#;8CPR@83.L&<RVTQ4a6WR6(L/d938,H.6OV:MI?A?LWQW;7_+UaC
)4GH:N9@NL(M]U&XZ(,aR?,E[\F^X.?NY=]YWT&?)KPbJ=5451UNf_.XHHWXNQ/b
,_=.NEa\VT(Y_6Rd#FGNUGRB?C8P.]=&7:^RMTc]@1,L,JT#GZbD[/fBYMJ+Xa1e
([a02=ReAP?Zg1eb>e\g(HK6]HYG2R-)NPF?),e67SSa20XR0aW]bPNJgB9CE8/&
5-HOQ.<(5A5\G)C3@3E_b9J#EYa_:4I>IDKND^/E+a#Q-\3S;abf-ec+gI,X6]1P
=3I)b:\R<#g<H\<CC]A:HYf5#MVFGQYNBAHW,Ad=NgDBU,>S?.MUVea;#[a;Z,<(
/K9BN4b#[B7\9V7FM,D4@C)4FY@IF/g_6@-B4Bc^Ef(1PM4a0RCOOFa;D\=8VfT[
GeIH3)U/eP_?e]:8+aXTC):@caG-HIbC:2TM\<NBOfaQcU9<dWD9g@4&:?E:]-/J
JI-=d3O?/R.Ka<Pg(_YMf_S^.T4XPMY9-J)D2^S273Pf1X7B=aXM.5,TYQ4/N72g
>M;U>KII?J36.=/0+/CGb<&KNBd;PKK,Ga6=YG#MbZKNXUWO54g56b==F_92T#CZ
8^<Uf,Mgb,W4]?\H7IV:=S:Ic3]D[2N4(\8.-:FWf5A.^NW<9gb.D?KY:#:7U:2L
N+JM5e@UbP)LMabR<K]W=2H0B39[(E)+#-QAU.G>&9IS#LS-R_SBP9<U<]2XPT+_
(bCEgW__5SMH^SM56Ba(Y02=;.=[Q0QHZ5#.HI;;I8AA5R/<E;X=6G^(C144U:fZ
<AIA41[\ZeAF&.\D\YE6)5@ac^3[P#C9M:#2A;3_(fO/,)J16<T&DO:V8FJNN43\
RXd;&\7_dEc5JHU0=Tc>OTVCI&:#ac8V@7\2S:8#7GO],N1I>COX[HZ@S/-X]EX1
,]3b(I@Hf=@5\PPg?M3:g<J(M0OXD?G\IBELE1YWL1)94c7Ycg^#S-e)WPF>MLTX
R)9P,:WQ0<(d7)#C&^(R9,1-D:GOdIaR0[-DE&GEVK,:b+:VB;ZPcA0&+K1:F2+W
CZGF5U>.Y?\:E1;DB31dF7]PAL.4L4DYAHYX?&TV>O?-f)Ng.IP]OTV>3S=:00VK
CKE6PgaAFPR-&]b\(YD\+A<C;7K>EBPb)E/[NX0E@(c44OV4JfJOdT@SQE3Tb@,E
L6HN-R6DB@?M5GHf(2\+gZ-52d]PeP1?d5B0?C(I<3WNAP+2:[LV/(JPg:[bEW5U
ICVV,1E@#+5P-N2&(&H,g=?7TC3N0dPU_K@?1OS0d:IQBTE,>Y7;^A0KK??DXa\Y
+Gg#d54bOE+g)g^M?OS?3b,XA5HOFL#;Y+.7f<Rd]Q1aA/E4J=5N=>5[^HbZ@IUW
R//3579[5XK0?X)Jac\FFOAPJH6f&2-e\=cdD[DOW46]D]2\EZOUEE??7fNXROL;
aBC/1:@&K<T8\d?dPK[5#LZ\)3<V1MHV]WJ>@[&c]PK^g>bL)KZFF<L+]NREE<ML
Nb:ZKPeI0O-NVQL4+U8O9#6C6<c^Z30F^<-g-QB0QcLYV)aVC9CM5+\f+4Q0),WC
3;+>J/A0/F66O^?>8.5G&]GFcP6B&[;;A6&95UXL&C;bWS_]0XSV33R3ZC,R9[:(
\K+\gY9#(K54_c+F377YbLR_OD:2KbC?E?^1N9g.<QE6bc3HT#RN;\?@/gF#K^:U
4PVc-Z5_&bAU\.04T0<W#YF_17DTUI@3R[^UOd\a;7dORJV7,=,PBL4KK7,O);;Q
_e-FMgT2=USTS02KQ,6VN:3L4:(7S_K5&R^R\Q?NDV\>X<E(4A=c;-U/9H-Z=cJY
2+.L2ZAO;e\L3K[P0L^@;>D[?E>K6Z^9SKF9+/J,G\ZAC+F]_(;3(6X,XgbD^+MY
b2:HcJ2]C[eJ+#WC4Kf9g/1&AM/=GA\9U?=Y]2,_A[&G,N\4\E?0.6QWMa?>F(]S
6bDJAH-^P#>;)CY;]TH)X#Y#,;M):IYQ(bYeUC]U(1;W.,.P=;EV)gb=:[Fg[0Lb
:KFDG7VGX7DLf7Ua1BC,9OXc3;)AH1,[HU&S02Z\H@N7J[SZe>DG7.SadX:UDBGg
:>/cdd;3SRS:+4BFFG>aNN,#6R4>QX-PJ9@?U^cE6D8gO[A]+;bA]>gF/c:DF(5)
eN04c00WG_Xd1GDXR.94T/RQ]UF&G(Le,:17fCf=E1>2A5#N)+KX+/Ge&:(6[^AQ
W1P/,R\W<H6]g=H[[8AMZ&8b2_&<:L+SdZ&gf>b;?OFQ#+\I[JQ7K<d0ZVb08?HD
K8gD:\efKP]Mc,VA;G5L6Lg>5GC-/\dW1V:]IQG/@4[S6N_\0#+HH^.c+T=))#,e
T-Cf-Xg;2+cSIgDHB71?&>YPc(Wd.VOX+efSJ2S5g\#IGH1],@/O;W7#7D#:ENgT
ODggG7C&Z94V0QddSbeWTQHJ(fKB)HKUAGAS942B8TB2G?/P0(a^OZ-O.NfYZU10
IH?SdJgSMB?9W1C=#[_@-9=G6Ra^1@+OaVb-7MM?V;_T)<C00g--ITPNZeeXJC)/
gZZG0L]1A?)+1KGBF2M4-VEC(Y]:6./PDV>dU)\21,LX+LeF@NWR:FHd](@Ye@7+
bW:IL[T4B7>;KDb[JL>D?I,dN--c6PXYf8gW:&4CK@7DDR?BNP?[f;cB\O9gLG#-
eD+N)#4+Ze1)+==?326_Oc6+b3L&=,STNS^6V#fNSZ^:#)RJ/JSIJfQGPC+G<L<6
0W9f@7g-0DG/NE2Q=4C9:V#?/EQ]Y@J]g2F:G6W=[UFONC(7O5R[V0L3WVM&#c)/
83VQc-9aUV:=7Y6[,K/=g/6f@bL?V-UZ8A]VH<P\G?S,D=Oa^ZI6Y>aEc9U=K?c2
DV&,S1U<P7R,A>9>WS<]9?f<9U\8D_P;5be7([5-aRB-,OILEBNOJT],KfL@1E,Y
;.H2dB:7S7Z_;cU\G96YENCf7XW_E#C&S[E8<+<SQ/W2_DGW<TPX4G&FX)D3(C-9
U>S:Fe8TS+JHH5ZU+ZFVBJ7K/fW[cHSAM,QZd8A#AaIaB0[M#@QDQZ;VD6<-HB&F
^SSO2WAg6gX,=Y+PE^9a7YWUeB4S6>Be_OE)8f4-2Y<A:NXW5KR?cS>e19.5>Jf2
OX2SKGb[fd^3Ee;4R/Ib5A[QOJF/Q,+HU;9HF:_b(F)V5Hd?IEHc(.@8(=6=4K?=
:d>e2_MK825LV#JLbg85IZ^UJB5/=;/b1.]eIOU?0C1.10,^9>IOID>#]^J4M&B7
\#S+_U^CJTMGKfGAP,_]M86EcCABc+F7^\R;>=\L-bb#DWG:-:K5U[5<0<06HBaP
1UISXXD6J3/6E[5@\6b&6Y4_A+c1H)1=--N=4<^U@C90?#+LWWBage^?gdMZM)C,
=:R/5K/DT<\@-X3D_#_;b5G,d59^=F(7Z2;,L^>AI@&WP=YH(.H]Yc&f8fD#9FC\
^[Y[+1a4e93LKVeZQa.3AQ1]:A\?F]02SRH<V6MF@;TMC]4FQY\KS-.#>Hb?]fFa
(B.^=3ZEY+:7=34+?E4TP)_2L&W1I.#EQ;Ed985A-(<Sa+X<KD7&9=^7/I1H0[;9
dMMKa8EJ6Y:PK5<(cF#[fS;NEfcIbFO#Bd:/.GRGD>DWHY1fO(bVf,+-9g=CFF^Y
AQA46D],H\BEPgA-Z234a170X,MK,^(#<HQ7O[P:7S_HabaeB\&#M8EPdV88W6LI
DdSFG:V:Y\]ZQYF\GSfE4U3DO7?RQ-_8de9g?28EG^2)PP#DcTOH7)b0C_GBF@NS
6KWQdC;<@<_0V(GJPdaRW)>3H3c[Y7756SPEX?8H4\f0P;3HcdYR0-1F4LbJW#Jc
+0FI1.&Q^AfT98VG609SO.dAA;NHXT6fWY/UB=\\b:#2I6[L,+3T:)&(E]HVJUaR
#09//?@P5T@+QD>RT7V0TA)I7B,#d=#Yf26CJF,^21LHN7)_ZM,^DVMbdIY?fc^Q
SZc.1+0UQ^ZL3@,5Y/-DQ/U<Uc:G;,6DJCW:.P(.VXZ9F2WT;ET6C:]b^8UFEETZ
0(,X@4_QDQ1IRL>;.d1Z/<eWYA5&Z2F&(6K\FaTZFP=4gC:2c,3^-2)b+XV]<,Q4
;9^H/[#CFEV)5#6V/=7?NcSP<&W[/Q]+=\2:5E9NC\gW+[YHVX-KbPG;.;@^P_31
+R?7;/,_>RF9WM<]C2.(b#bJQ):_O&EN3LQ=GcSLR:Z^BKLI90B-+-,P>W0&81)f
@?NOcd,/c=L4Qe5WFEZ-3XNC9U?W6O#eH;f(91b)Xc9,WFPQ]D0A\4,QM)+)3a5K
F@;[(Q#cCg?4P9&dGNM#IcT9eG18OFdddXg[>Q@N,3T>:N[cQ9Y>@+R?QD=0[857
f\G/g@Q05AC+I.V8EgW>GPW@HT)F6K@/][T4QV6?5eC-K?FEEDGfB/N>3/]C+JX;
FV>e<5I.T-;DE@/J5V@>ALc)Cc2U\X<G.RQ+FC@Of3UUDP,K2\(g5@L+@ZC1D#;L
ed7BQ[4@=C#GX&<H0b<DGfS#Y5gR[,W6DgfIe+@aABQQ7?(bD@M;0Ub>RIAR6QYJ
VI,QBW1dE:)PX(PW1RdZ&?K.f(\VCIcg3L2X9gUJ1?_PNZ.?HC1JdZGc.fU+4R?O
3dND)Nb<KJA7(N+ZW:L.;8:3-#H6B3L<U[4GCgYgg<MO_XOC6g(R+^4DbTBZ<;=4
-JT3+R-Nc)LRA6fY);P@VW#Yb\fBH_W4][d.PXSM[8@_#>MLe;c?ON];JN0,G#3B
;?-(L6=c<[_QCZ(fL_^]LD;Q>bNe?C#/RFO<2X4&L;1RGYNPN[N(65)[0LIPXN)J
_/O8fM87F,CX1XQae&d3VU9.,O<6]]bKIJcPd1.JSRUCC=A,L4f]@=PKf=6a/cUE
#=M]5:,=.7)4]EG4AX]I<&=NFgQDC:^/&Z1QU)U/(7+BK>XGXfLW.P9EZUB=4H4e
VggfaL6CQ@R]HS?EYTc=HEMB?^0/^^SFX?^0MM.?&XAd-[1CTWJGdPR?c4I#W@WG
b9I+dZB=_(-_)-&IHG3(,b-X@(e>Q4+:U,/\MGf7ZR+g4BD>]Td#_4=&cNPL_9aX
Z15+1@BUT,5ZY(Y;N@:=\@VOXULX5]W=MMPCJ=U:+Z;g:e]WBefGAA.=7N+]J&^>
R[;OG_<1(XW0XG?P-T2/dBR>E0d::]Z^[f47D9.MY>0b;G90QKEH98;\:>8I4HAZ
_.=H2K<LMYa=KFU/]3P-.]f:@a^3^:RN2E0J\;WA(O<_4M3NU6<X?2_=:bdN.97P
dOH4D@(H+Yg#a)_[a1a3I;6]R-fMYWM#+&PY_?CAUN-ae5<5<L;19fZIEf-)9_F)
IV@&KD;?YDUX@,]8dN-5]JUf98;J&B=0f:Sb^g4QN6LHC9.DS2MMB\S<F?gNE021
a?\eEZ=gI.?FNNV^JYEB\13T+gYG;#R?[[--gIC[fWU.I9J7BP;HS56Q6@=BRT<=
1.ffCWC1EJVIM@e0\;CFJ+Z#>2BJI[d/&RKZb:AcNFP5&3XSIgXE9T=Hd.;Ha]8b
f,NDF2991c:ENI8Mg=4X/H>9@Ze/UPX_A=+Y,I&<&>:448&S&aN28VQ?=)5,T/L9
aU<KBK:b-a_,-NQ]e=J<T&1JJf(QCeD)MB#NbO..H<[Eb(JN80GdVD_;09BPL6+f
M;cTcG_Sb.YQ09NOCBCD#.?8]fBQfDVUP^B)1+fRPTNf1>cS60a7(3Ic7-f6ggN;
8eM-BZb8@YEQ++AP1JPBQ^\^U3XW,AT1L4Q[UI#ae8R9JAYR6L?)>B-GQ>&+FG:a
#D;JT>KdNGNGZFA&.(.0F0O;D^V2IKdVKCN:GUK38<2QX-<?T+N(]W4UFT(eVVPd
HU>b5K-587Y,.(51ULY>1/H+_Gf89bS#5SK#e_)U2P[;V;bM1J+T<7aD]THOZIfA
S=fI@H(0(U<fWPdPK_X)AWC(DST=HES<_<P2BOaKU#[^HUT1d6EXMGAFdQ.WT,c+
J2)Af#;=UKM[MJV<H^>;#>6T,U7#-4=F26,H..OD=O),GI(Q(J^,5]SFDb<D#K;Y
R+SXa/<@66]]c[JaN//eA>7S=P;JE/9cec&GDSZ5>bC6\_H8@AEY^_ZN(&BX75e^
4/V<1<7C)WR^^;c(ZD6M17GA\428<(&&dAa-Z&G@<d&>[ZdOb@R2(H#_5L<<X<WT
;1NJSE=Jc4X>>SX^._;(=fK.1f@_23(5TWe@c>c(1^+&da\8>\?KXKXZ&Gd[I=+6
<1U\?TQ[8W2Z>]GA_U&2(gdX60_/cf)7LG^e@O-c23&#G/L?UV+P?)b<_AJA;Aa>
&dKT8F)Z>gU4M/=90W;=1^&O52K]U0<HFIgLY:9O-LL?1fOdK(JF4/8P[15HOd4R
_.Q/6@g3,ZROeAb/c/0L:f82;(JcP1G=\=a<R;KK8g>I<Y,U:);4FFId[<36O32I
<He<:Ag-L_S_T]NNFJ0ZaKc&2:0:YEOdXA&WgLTIg8:fP?gIagf5O+FOD:_A&;7C
d]_g7M1B2;dHdL7\J+aRN_fCT(OD_<_WI&=MUR>c]\^#[B5#_Sda[TP7[f7<AXPP
&=f_U9C/g0KYTd+A<4)KA[FH-PRV>E]Y;]BMdMf<1.^G@L[cPU-cF]#VDR#H10aO
d:F#]W4V6,?:D7COT,:>XSI4bg<2+3OOKMAf?ZG-ESI7#R7@A9DM8c4]f/2g@Y,4
2/RS@fb=]05egE.-@Va&K=f&D1>:+GKf#bKYBN.7OFEQJId-LX=E3C#[,AP<\b;[
71(@P/d=&.F4.4/b)EDM@/D@L9A_[K>6H/,cHWNN4G.Y^H0_A(@9bFJ6-72a@TQ8
[gV?a1<8)QG1N=LfO2;]K-LN4>g4KM><gHN=^=5?AL:CYgV86QW(86CTHFg?cJ0\
Qa=X,O68f/a?SOE/B?2HS^g@761e^4YUVETcQTb@5W]Vb20M755)<a15&+S6S0Lg
I[RI:G=\I46N>WV4M-QYYVT.WX]L\GN0bI)W80.LH3A@c(T.Q8:FR\V/AJ.,QVTA
AcK#;1FKX>MD4MK_.VW/+1VK97RL18R<7;Y/LLQBc=[#\VcfNZM(/.#LZP0H/Ib/
8[[7)5a4/LbDYa#-ITQ^.IB1THFM9\=fW9?08GP7a)SS2F_21KE?R8d&I-Y:(2A#
YbMFVPa&S2)fF/QgW_6<JcG6eB0(I2TC125QHU/27VAeV1:cKQ\dZ3.ZHM3bRV:/
@8W4WeO?1KTH:XG?;)fKZ<7Z6GG4JTBU9,N3PKH/YH,,-@FA?T=WAc;4]V_V4+c,
7B(5F80cc8Ra<&D2L:S-\0e_>f7I4F06?Q^54ANe>UeJWKW=XRb]aN2HN,ME8a?R
Kd_Mfe32G]Wda)A]T07HLZZ_\a^Pd26QY].bM4ZAI8eP1\OAC47LOX<RCSb&9V7N
]ASCUO3,=7LP5?0c_M-61679d-f?d4.E0DT3bZ\ZGeV5K+=EN,bB3/<e..P-8AT3
2T+))7-a-=/YT@3aCFV.F)BR>#_/GX5M@3E-ff[2<N?6TY?0N3aE3-OWU-0TbD-b
AD(C[f;(NcXfBZMfa+VA]dV]Ig)\2A&259CQ\R5d^&-5N/ZaR@IQ\)<1^6/UIP=H
(<J,)Z\8Tcc?G6RBZL1TA_g4##AF>bZ9)3K9+P/U4.)e1CbUO=62+WeTIQE.B6C8
7MT/G@.M9<;:,;Z[\0a)\cF[10H[b2-PB4fg&+(?;;aY],Fg&OcKOa>9?=?.+2=<
G\7(E+Q(WB]afaX&CcHA^G@KKX+IeW)c1H);C0d\/]][V3A?I>U\M+Y@8,c6VQ\C
gRJbC@QVEQ9_6R.,C#SEGIG?N.gK_(F^5DK;Bbec#&>6Ba;L.3;ec4;:<PG1AMX^
c]ZZ)AN.Q]_:.OHU,ZXe(&.2=DE8O>A/>a=b6<0eF5]L0C.?Eb]4.F-^&cT@1B>0
bBDa4:.G;TY2Lb2OR,OLS,?039RY_BFB@#a<Lg9&Z+Zd:RP?H+dN5eBV?.Fd>NZ_
g7WfV-^;3;AGC.C^.+X@CQSTJ,3RgMN9D0aeAS4\>^+JV\RYHE2O34ZE3GbS[e22
9[T\,@=DM8\J[7/4T?(BA[HP)_+b+<^A5gW2REA:)J8-.4^@VMZ_@[7NWCYLL&I2
Q(beFS/-C42Ffb/ZD9^0S.:B?6K3cf:7J0+bcFY3HU(V66YJ7G#D\ZPR/4T8Fa#3
M4];_c@#61F@P(DM/ebMa\;X8(W-cFZIY:M#I,eO->-1WJEHOR5;)RG0O003J(Ve
^Z(^Mg39XO0-7eOR]d^E0;PdA<>G7(),9IY\IF/2(Ed?748F(_fe/38DV97EOG/C
CH7.-1J(V</NZDMcSF411:O0-C5ITJaY=(aeJP&b)BC@;DS^Pa@W&.D;=)gOgH[2
/S(B#8&>&8VZAT2aN3A166>OJ07/K#(Z-dGV5_I_DDKc9BT_?9eJBbgY\<M7@WQJ
M4SJ\Y&+3?+5XE^BJ19TgdF_W#K4O(8=RD)8:8;e;+4;+\&YS]fcLBN^I<409_UT
f/\c,KX#;Hba>aGE,aKGP#VD_\AUPBgY&/5C@FBQA5B^V1:[PN?Q^AU1_/K;D=2b
(2/6^&?0<0DcYPa)1C#&PG((9HQ_4cf-<ZR3I1;:)M=)4_g:?XaEZcLYE0VVdfD]
1S1/)NCK+.^=ZG_/T<eTFF1FKfE(Rgd?8g&DcO2URg00QNX[WW#Je@-A0+9?@@8/
6@O=>Ud[F;UbN[\6TETA>SHNQYVZ5G5-3W;/cZ^EOYUeF3<F&4bW.C5gES3(#9Ha
HYY\NQC?2;ADCI)cS;:eEII]72>6E>HFBF+.A=@CZ4b=0W3+-57:[\+W;[8V[2RW
RRfW^Hgd(D>:KWR=9E]6aYU;3Lcg9Vb?7He6&D3,1ZY>9HgLBbaeS\G#CeU99+Je
[B(55JCUPFM3UQ-\V_@c/c#.LL1A7bNZ8<LbCV-bcAN4Q.A,<c1PR#++6=]^L-.6
[DXHUQ1GQd7(BPP&7&Q0#=\2L8Q]+8UC&KH]aGHXR\#L[V59Z<<^O.(H9KPB1_&3
?bN9fVZ.1#DGB,FZDV,K23Z1<<(dXKJ7&5HV0GT-7O=9U)<GW6/6C+D#H8MFB;YW
\KF&SP22D/\ENa-_;Y@6;\3LP4;:d@Y]>T?cO3FO+5E.+XdX04OF,P/3M+^Ub?<P
]TJP;gSaMfP&b3;E)(5IEbf]\H4#.6/d3<8#bEGcf>Va-ON3&GaS>5K<,JMO&T2.
_TK\KKN-P:+&>&Ddd=&0b5DX7BS/HbV3PEgaR05ZZEZ@Df7#;_VHL#E:)6JW)MOB
5S]JJfeQ:K0Jd[Q348cDRN]S\5XX8A2AB\f:c#:)^,^DY0G.M-3@JLU[e84c2XN+
b&?Q)##>2dQM?JYEXH/?-:0e?fB6.<U2T<_Zd=XO#A.]1KRVGe;=QacETcNA<bF4
N1#-OfJd@69>dS81P[_(--Sa7(B>bC:bI^Ud0<P_/SA)c\X;YO^WTc=#FF3LHN33
PNX<>(QTNeQRE4Jg7IVRP^+12\XZ886cX5]]MLJ[:W098J9aDSV#c<DEF7IYCRGd
EQ5,feS/PeTWRRg(:CdOBCcG-X_ZTX6CFHBBA+05O-:D)GA<JLf4P06b:(380FdN
9E>,=L\_YUDJ_I&:2#43Uf1D=,WA6X_McJN(B4M1C^D--A38A^:e0<;HQM6:ad34
e7gg^;JQ6#\,7:<E/IfAP+GWUeFSN\X2]II_T>##_9b0X5S5a-:Qb+P?X5N3ed[\
c9J2F(<7>B4Q(1P+^C(^AgGb;PRf<:::CT?^2g8#(]@@[FK&3ga)aTH\#--:X4fG
IX+\[GM:HUJ)(Id:ecLd/<,VfYFUbYRd+JYGdDRB.S8^,1Q8ZS^X4&W<OSGFcH03
^3#,58EfDgIaD6Q)[D.g-.1_ZGE>ZJN>RB<V0S/NR_;;cTFd3FN\,YWZ=X6_LaRN
^_5Ae1Te6XAQ,4TfV?7Rb<1HU5Y&+?N=&L?+D=O?;XO0R2+]4SfYBf>3Ea2/\H?R
\1O;WU>H^_Vf6eBc==IOSTJ;-&@Ef-T75/-:T#E:1W)6)1B/7_6V<ZPZ:<CVSSY(
JM7KU\39G2P\^J<UXI0@(6HIgI31-:9MS3P<+P[:aG,F1_5UaTHD^2U7O.Q0a[R8
;C8_WG=@&+_5D)C&)Mg=.O(8FD&2UWNZR7\#>F;eBXZU,S>+;?&.W1-4H/[1OJ8c
CFH-9I7Z^9C))H0eQADT42V?_]:772a?Fd2X[H+bZ=BOKI[aA]\,#N9;DD,J2J9L
2E+?N0#VQ40J;,Dc56FRF<U>/2fX6>\T0XI6P]8Vd\UQa\=W0fb\]@8P;H-80)9<
DKZF3PdR-W+IfeAbWN&I.EgVFQM8DNaW,R=Hf-0cC-/fZNg-9681XE/f6WPf-6a<
\U#+?#8S,YU<Z@6O;^WKgKDWFc-D>8KQX9-/BB6^&1U3NC/M;JP0BV[Y.L\FLC+I
eXV,FfT6F):/1?e)37O,&F9828]J0gRA.WA^I4cKAdYcbg-KMV?),[0XDZB]\R6E
LI-4WbbT@P2D)ZdWDcSB+.+0,_8>.\H+Md-3MTc7[@-:QI7/21dSN+8RN.08f]+:
F+CC)5_\5f@Z)BAB/1H)19,/JQXB>bWI?,QH(W.?E\Q6[g<2_:;=bZ];9@R0#1MV
[Q]1?4+86Q(=0_@1f8>\d+^-P<a0UB[CBG[6L3]eU84g0#KW8E;3MOa@#fPe-2eC
.<d&)2=VP]Qae\E6L(9EcBPJL^XG@HCMUB)GZP>R<(U4A[aDW-SAgYG[#VY6YB:+
g#9)[2.HS588eM78#D,.bBM3INJ#YNO@:G>]N#2&N<b@Lg@fHKWgBfMLe0g,J3M.
,N1,]R<HFIa=0+Xd<E2Z7.S^2_SZ_,G9b@C9>bHVF[1;2))(;bgB/OQCPNcPP/..
MQO-=D_K)BI:[=^/WDcbN];cd@[B-ZO^JTS11MH_[ETZ.B_OVO.1RC1g+X[b1<K>
L4HK^4M,<2W,Y6A=:bc;c;B08]&B&D3#&.X@&AVG);+6(P1(7/f8fF>GeK-6=7@U
P.g,fJKc[5R:FDF<X;)G2RC=<UEG:>+M(;EY.Y\H+efP&Ibd)&+FX\>HSQ14&+f[
GDOAZgN56@GKLMX9_;[=A91=Re)W]B@aL\?d\[FK>YD+)/5\E)Bd05O)gMe(9OB\
2+O_-O\>P-8ICWEX^cWcN::TECN5X^-0VBJGGHL&.-^DILR19V+SZV//P)9Qe5E&
K]+Ga_+cMT<3C\1gQ</9-_PAbLBHWOCa^NffNN(S3egf4##TXaET0#9;9fXggeM@
O=X+g?_8;2B6=V3GQT4/\.Z07=ee[X0#MKE_8\N2^<17=dTc_e?Z\-ML0a+^G>AK
Ze(1Q47DENTIQC:Q52(I6U_^.(c=(0;@HLf@9I\.2WJYbQQ9O;+?EM\,87ZKH1K:
&@.gG4>#a[8-)7cD6fKZ2..\#;,9b;EK+W3TP4HAg8K[CEMA5V)_<:.OfXD2-Q4g
BXY(P+401GSg7L6+K:V]F^+f,K9PUTW,.]Ug]8S?)O+deKf63bDH+FN&;a#LH6fA
V-]R>-C6Z=[Lf=Q<A#b2Sg,:1=M0E&57a5_ZX[.RUY#b\MME(<M.6>R09YZdQFcA
HGYYZN<.FL^?#,#<f\7_6?>REM5cVCEfZLQ^ZOSJMT-(@E3GPZ1T\=_cf__Z),2G
OO^\Ma+4R0K0[8..(Va3e7-W7@L6a45;S<gPVgL)2BJ0^;XY94MU7RYIafg(M;OU
^3[[L+X4d/K-\Q>S(3?eC_1L(dH3V\GZVL::]1K.CJ?cIa3bR;AI.GAObNcHGT_F
>QGaGKR:gD7YS845MB[a:X:RWL+B5d>e<&X>:f><2Z\1<-)0L(fN-cV+L+fgCf_+
SIW4QbY^6Q\@0ND-1S8McIVQFGbJe(BHTR3X&R(IW\d=T[.4^=DX,<E\,G3]#]Ga
.]Z\@e9-TJSW(8?((OaE>9I<Y<K7U&B+8?VYX6_L(&TSVE3]Ee;?TfD6Fe6S97F6
RLbG9g[aVgS5UNUE6J&29_WA(=Z&->,Ie(JWEQ?42FUSFQZ6+LUYV+QJEYYZ(J5)
eIARHHdfY4910B^FZS#beZ0)(9><WdYV@e.?c?BCFVQNeYLVQ.]B-6H4LPW]=CA]
TQUGEZ1E:PEC5FZ7#28V+:812-2,TVbL0EU7b3ABb_P7YA6H+I\ObN]MF_NPOZ.D
;:Ge4dfO(TfFPMg0b.4fKeV8@+.OU2CNH(_VBS[FL4<3c(]bfV[SW(91<]S-TZIH
&(d2@Ed#8-Q:PcK12O-Y6X5;&A-H<>JaTH_3;R7I.]U2QY\N<Z/O5L)eGH?(f@\)
.MZ7XDQLGURU1eMS?9T<,H8-?A6?SCObM?QT3aC=CLIM@6?Zb>,B=GfbfGg?^Z8]
>JEUV;N\cY_&\2dA1;7LV@#YbHeb)X@cB[f[eYETWYFB;Tfe.N]J_PX?5I^C&dR:
;GS6PeHEFgL?T14+#9VIa].eI1J@>L(Lce[_I)W=QS\PZ7?c7bX@2E3<6d22WYXA
T1cWEF0A?#Wc?-a1<CBZ:^(=Z+&2WMP,^X?YT]1<1-V[Tc+S8UL_I0bPc-:a6ZF+
C7,6X(dK)/UAUd,3ME@A?I.CITb(1ZFgPU0Of[BO#F>7B<<,RgGA+fPJM)Z0HZ1g
[@Ddc1\c7b/?6LVP^&#^VC)<I#>7WSO>c(M,W&G?eT1V6BN=3WS4c7Ua9;(&Z-&H
cg2/c89ZI3AcfQRcf/]AON<bcQeY-I,OA[=Y_WLR@[3ec<UZ,a-1e/J,N]:/^_2)
QGI&/I116eFU\TJ;g;_/,L8#+/-I&;,S;^1)X.43b8,UWCRDVe4=?V]YMMVb.MLS
TW>]AJUUHMfRL#[6J,#?IBE>_dO70bJU<20DW2IHXC?EW<D0Qee@4(2VW/(C1_:-
V9QX)\1.5@LJ1T?TZb.G)YHGc9Y>,U_OAO2K@6e#D9A@SNW[JBgD_\<EQAYeA#S\
:+BFR1HZ<-J,(&O;5XI;4Q@ACf-;G-S(6O^#REaRd--gc0E(+^af8^81NHQ^@-)_
K2ISUD6AIYI^J@V).NC_dg;-SF@>ID4U\gc38Q2d?DMNU[L^8PbA8S6:;cXcGH:A
E#f:IJ/,TB53JV@RX>6TbLGM/:X+eW,(Aa_)(ZHZTIN7L(afgOd+@/YTUcM-U&^>
+J@(:I7JA9ARH?/2f[6T,@CS8&.\QM1##a16>ggJWVMF^9O\,;J6b0PK?]2HOH#R
=+N3)8[+Y,IW,P;[T)\+E4H[.f@E;@2UZ8aT-ZSW\88A\UJJJ\OM8fILbZ7D..8+
2;)06.X08/ZOOS78f70(^+;;S&C+?X^O_N:.K?f.])eYFM,b]V0[;TFUbFbNS^Gd
O0f\L/CA?FD.T(>VU-=.<9M-NMM.Y#./JGL3=RRPE^.-D;1bQP_)8T0VZXW>LRM&
O2+fb>(MO3\0ScP<GRg]^PcDB.#N@OK(=KLTXcB89b)f6Y4E,]O>-HE,4JC-W:<#
e;SR=(G];)Ze]E\6A<+=QYJb/=72Q]&;A-CP940LW)c>;,I/LS-I>0VNY32)\\G]
Rb/@Q8)c\H/58Ng5K[,9Q6fD/4@S?cWaF=B8c);4cF>aC&,CdX^GZ&a:f.Fa\RF@
aY[4WF8YZYC<+0)6D6RP=aBZMLL#W,aQBQB.>9L[.M,f9>:gb.4e3_R3,5(G2dgV
/Q@8<V2TY_f8OC,\R]C25b&_TQZH[8\V.0K06^QQOX+GY,?&C^cH=<FNZ-(9>995
;-(JZ@B[CTZ9f^f&&J;AD1@GR3J(83eYWG\B-)4e^O?PPL)c@VR)X.):f[PQO&<Z
[VcL()CaW=Vg97_F-_B,7?LN0TG?@CD<,@48T^[HFP^.G7MN3;HfV6[2Y<3fG,LU
I;M&J7NZ,[4KC5Fg9JB7(e5UY8)T3B>GOGD96L<bc966gE(KfPYEKRS-G+>9G:VU
Q@)L50?&..H]_UeNE.f4K.OSFD3A]QHC6aV>W.[4Ua/Y\gB=[E9QAX&PAfNb>;DT
g\0Qc@RdPZT>f&41^5[;gVG@b)J\)K39H?7.6,0<RgD3FL3dNBMI^PHRQ7NKVX#/
.VS\9-P@Z_@-KBD6D/d-5IS>G>>@#B9Ccf2IW8]IUTC#Ta7UDXF#S[WPSJHcWFMJ
JC^;(SZ6_6Q>;O2CLEF[);-;V8\H(#K(QaY5EH:&R;C9L@.0&^NG3^68\+4[=NaB
.cWYdFIR&Q6B^&YDV;\IT@(L1V7YaSWIZ&7ab871?I+R]L6,4A1?A+-c#TQXKRCE
,RX&=];Cg@]87G-BAOV;L3VKOdRZ3O<fCKaOO+1I.I2R6dF0SJ03)W]URXKA1b;X
fcE]/>Id=;C2.MKZ=:K++-9,3\<,O?YKJM2bb/CEQ]>QXf\bTd4?2T-dC5E.<b&;
J65JH+H^7[KMg+1Gga9-.MDPg90ae6Z+H9J.OLA&+&bRYd)QUT]J3OG#F/F82MJ4
JL_[R>>&#P7F<A]Z<d:LN/MdZN,(US[Q-3/V1E4[<546CCQQE.U64YH2?)a(],>O
ZK18EOJ8(OfcH+S-4@R^D;dWEL321Td/T_1WP@U5(OW,OWRU0c&g\Q/Q+UJ,MCJD
6\<4\0.3WKJMeG#]N-+J6Z_\:5.SYA,\63:)eE_^Ff@cB8HH3-F7,6.E]AagBVQ6
.PU05#VS5]9^<I8-OJ[G#>0FT>#^5VJ^ZZ<Y\N=a.eNJS+Lf8N8(@0.3YZd=3[GU
@>L>A&)MA@[QX6ZL#D\KHgb/M491\TA4W]Df)2^HM>/(M;=+(;U6YE>B9,)\N#+&
FT(/TX,,dH2(aSRTA=6c>Y_0&[24Eec4E^5Z,05E&Dc6U6]b/@e#BS>0;V+IJ[0-
Q029B=_IQ6R+ZSE]>L(YYZ\XDG_Y#aQ8/UF;d_&SE8X?;\&[L+LV];b@+-&QJ;7G
4WTQ9FJSFbf15K.DZA#R=f8ML,a,\UQN11.=JFMBM:/25.D\\4g?@-;0CI.5UOUg
R8BW(^Ee8[O;9=7F839ZC06+#Pb#5&9X,UCITO1N#1/b7ZNX:>S4eHL+-F8H[;Z0
QKBP&^W\KUdZ#8dD=)#NX,eFAX<NP,;g><gAKUUSON9@,RI9&TW-CO(K39O@(#6Q
(-^0IH<1/>9c06SS86LA(4;4cS1D4=2+(C:cSI.PY&d6DW9<-30>1b^I_>WB.G?a
c-32YQ2Z@Vf-ebW8<\9&I2+<Z(>F#/50567g0A-Q\:.=Q4&a<YY<^d\g_-,E+2QO
VL>VRf;6WE=L3D:]@?3cZ63<fCRRF6D9U0SNS.[&@If7237a<#T:0YbR.O1LP1O4
E&d[)K7.(g#FL78H[#JX&La@H&Fa015MQFcgJU5)d#-G?<b:,.OI-:JQScYcRD[B
7E4>,eAUD;bdH>N8ALfP8C4aa]0J2W)DCLC_caHAYLTB&b[?cVLWC;Q^PPO;L:,+
c0J<JY@)F8@X2^N7:[EXBOU8C@&gU^XCO#WHV<8K&:XdN0.g(4F/W]SAd2P27]M1
-_Y@#P..D)9e:bZQF)U2VVZW0I&VR+>ePU+J:3=WbQRgZ>1.e6QB&U]fP6L<+2Q?
+4-:\.Jg95E6W[YM;4;F>cY<UMZ=-7;2:=3OK<g&F</IgU+OETTgTfCc#D[D[8L>
f/N0J>G;a/,=1KKKL^c+1b?5S8U#gWR1[/a(aV2G#BG0V?/S(3[623@H6MO0TA99
>c?g2&e]S9A@=1G[R4d0a\A?4M>&4R9.B@[?7:ZIe+Y1]C)?B2PP)g-+[V9/FK,Q
9K\I/;B1L;-P^++,=OSHDMO1](g;3?EN#_TN\N)9-DY8NN@/0TNUR9RE5]7Xa.Q,
0K=E(U(E[NHf@Q-C6]YT0@ZJ8ZH_(I4T3cc\^IKOHJ=B,5WcUS#b=VADJE;&2-@4
RJSYOH.&3/^9K(?G08cX?=B549@FG8HBPF-YRB(/<ge8X\U7/OP&LHb0R6,[9AdS
NE4)#R0cOINa8[?;J#Q>B0N#AD3VS[+Oa-&-=1A2YOVDDL@RUJ(S7:51/4S\&D;3
U7ABX1LL9)\[:)cZWUZE&<66Z6gY3-O^b&@^=KdA_PE^B38e7IB:[2CbMHUX#_H5
.R9EE?:M3ABQBE</,<F#[=H<>XKe&^)aAb]S]<1:_F/G?gZ[W?DU9GgZKJQMB.[A
;=X3&9baMG;6WN=1RRA<Bc(\<-P2=egHBE4dOZ7U4=_X=T88XMPfYJ9gFG6Q>I9.
cT3?G88Jg6^3+S2SKN([;(bf1Efb;7<<(5XQ]LU1;b-TIgE(83O_9F?-:Y,PQ/#F
LG5=8A\fb^JW.:6_@:+a)GdN[).8(DSS5H,HC@>W0=P?T)GIORf(9&6(e9QWX??e
>=g83gdS00=XZP^Id(RbJ5E>.=_GEP[9XEa/bAPbE&@D8(4(PU7bM540bC&14QJa
9Z4Y2@-UeC(SMcX6,UAB:H+/9fg4.UE>bT90>]<67,6E^83=9ZB079ZSYX:]/5Ug
HFK4e(+R6I<9PI/E5:\:YI(@:,#SdHQc;>0XD+JU;8IF/fFfg5f#7;P0SYND4,MG
Ve(4L0?2U(L&_W):#bY=#4N,M)D<W__,cBH;:2RcK@R+[F-UcTK5E>#RF,Dd2-bQ
2)P=-YQGX)2a^9)9a=J.cJ6a)@=&0<0/)R;M7_NeWgEb^\WS69+=[U6cJIRfQ.Yg
@<FQ?5?R_1XUOf4H1DY>>RbN=(?P6;/c5EZDdG,)(9=J?LM6EFN:3)fMCS3V(C)G
SAPW\8\5VTMLVe[KOZgZb;9QF]Pe(R.#AbK\)b&+GOK,>YdI8)RSL)_MSfK8;cXN
^/dd;.b]Qe8W)1N^:aO4fKH4J0[(QLfE,>RA/VZP4\0<=&e@&\0O266.1/&R>T]2
<2+<eKeRT3g@9U5;dDg9cb=Y^)<?F.H>7aAV?PJ2Nb6JZ-^I5_GG/39BG:>Q-:0c
)9K8&,.A^N2N0aNV\5F)d^^c)5H;YF6L8JUg)CSZGNX73\TLUAF.#Y,g_>ce?d/G
@2Eg\]-gV7e0W_H6+@UN\MCQ<0+YVB<:>1Tf\dP4/DNJ+[GXWMcDI:&I@RfC,>gU
Od4\Xd8^#NcMcKM;EK0CGLb7<)7f2J;6_VBSF@))JWI)GCV7)\T,NL&YT3e7<0gW
98,e[A-g+HXG#](/RZMf&e6HbO93G=+cO>9>NC,?3Hb#OE4TO(/5VMgMJLb]EDb^
^3aQ5B\I#eY.9Rf+(7GCaK#&IRE3UASeUA=?efIVaM51/CZ5AeMG@&;LM9B7K&:K
=@T5-E6aJ3:BP,0#(CK[/#.R8PNH(@5_c10IVOfEBb-cL5#5>_bPQYad=\JJ.@=d
S4S2VH9g<LJGd6=^dba-G5>/=:2-@LZba:8KS7-ZK:aE_Ed71F8(_U-^Z=GJQWB(
dJFgCAW4B:cAGXZZ0:-?\GG0dDO_#+(XL2Ge_?U8Tc<fb[eO4dBQ8I]54P@,?CNE
&XeUS(KO\N01g-/58CQ^M(CK?e)cVJa&76(;+gYe.)1-:_^a:S5]]VNe/X\G)T5b
+f/?d@D:\IZ.08]?.<FfLXWE]Y7Qea^W>7<#NbS?+1OdTb9H?F8<<XVDABWEE^d?
C0_#Of9C:C1J[XH;;-]Ca?Wg]]7-]VA9JX&Y\gZ2ef(@,\I5g18OSSgQUNHVLN)T
ZFBU+PG]BA#,X1LK3/9VZGE/[@9_@:[G5f?^TTMS]J\Qb-Pb;51?&9G(H+PT0E;Q
-V^6SVLOQ#C.[)S\M-<XC-N=Xc6-fNe?=FgVIPEZP]?#_eD1SN=KI,YW@OCe([e_
VcMPdf507H2)@JN=CX[?J7L?fWK#[#c7CgD(JQK>9ae);0-JKSD=F+N1&+H+V8K9
&C1AVV-CARJ)=IAa39^b-VLB(+-FcVNd&T379M:7(c/BXY=(9DeA;gZ^[,We[.##
bK?)WP]NKEX=Nf74Qd)d[9SIc[VeOLfO>>_cHV67NFXdVQIXB7@db.+/92e-g3B;
;1Xa0,3][D4C^>YE>N#WaaeI>S6]1E@H53a&-8M)<N09VQefP7,?fT#/bf83E291
f1T(6P@==;DA59E0\RdA_#EKX\E5[6bS/.cB-]GQV(cW5V_DHEIN^O]Eb\^YHB>7
6S0;E1Z&FC@ad9[EWC4Q4#RW=Gec9#D;8-;XaM+5L+/L\cH].0#S#B//7L,6\_d_
e2JIVEG(d=g1G@T:L4NLS069D>?9V0]B<(\UH>dM5F^N_a:.eUH:R6-&Ve)bFI5P
=;R0,Xfd)HEFW+-G]-N(&fZBQa:T8BbA1JEb[d/J2.?/T58b&(^)L4)_fHT>9+;Q
:C_A;36>8cELgUW_K?[PL&LG3)I>8JcY&J&PJ.4F.\g&ZX#1e3&^PdOY.cI]Gd\5
\#])e-69H@cK+>3E?+MHX<J,S-gV]5ESbNgBbQ=6\c4\LbCHLcRIM@48BF@LF>#0
S9e[R=J7+cAV0Y&H05O<[(gIbT8S\+eB]F1/\d.6=L&^?],-3SaJ108(dI/;O[WV
MKWDR]MB&\e5KCb-=3V9GBV^a@f<P3?B5(+Q_(\.IV2+=[@MGf&=g.5b8KOV#[e;
,_=71f42-GN\,&HMOU^-cU;VDRa_<1KG#V2M?D/6C)5(W6=f;LLN)&f)ZVT7O];2
U:(-aVG9c\;]WP[.g/XW9<Q\cX<E9EIHUNNSg>fD@>O&N+#8V=6?OQ+M_N3&VeK,
C.R&gF01=DOLT=01(,C(e9BT]TO,<I;#C,=VVOWEUYTDPP)fHV-].QF_Y.EW4Pe,
-DR.@aD,7J38C@7ECa#\a-2D5(=RY^<0cSHI6A6>>6bd)JX^T1Vc464P4aZ\KcBe
V7[R<YNM^V&.F.SR^eK58[A27P1/C-Y._0M(Ye.,8YT^>L)70_gf:MDD\>L_X(IA
aDDMK3>OC-,Dff,7Kda((5d=b+3SGVNP\:2U9Y\Q>^7?AAS/fZW2[f?.M6e9/d;C
@X]&H,P6/=Z08\>;b;7a4062O[]6HM)QD=?S7Aa]_WfF_@G3(3K^fe5#ONHb5X)/
1L;_cY5K7&gK@PD0fAV^7?FN_4f[CZ,a88Cb-PCJ=^99&GA+AUEIJP&aN5)DZ0-5
V-4CeVATEZ^6_KeL2>ccSg3AF1Bg.=_L3b0Iggf;IOgO6d]NOM]-PV.TQ?\^Nc6Z
T#e9Y9Z7)7]=a.WMLeCV;P_aaC\7CQ1g,G9f3I4@+>49FJ1[5:Eb?H.9^/+dX.(,
E(BfcKHJgSgUF;:5cN5g>UJ2_=NKba2;@M=&_+R>7Wb?MFMdC-C4GQ:G]c,AE0A:
N^]g07?_;-2]US:dH\1.4]D+E]+XMg^.JP09RD7BS_^7@.]10.HbX9.R#AT#OA2R
TNY(/;gGVP_4F/LcJS8:LQgd/[KKCA[.FC<B-\RF@[&?6EcLaY@X9<H>;,^;fINU
QCZ,8Nc_eGBNJG=5,ZX.V5CIYbea)F<cg4\e3&JR#PIV0T9.#<C)Z,36^[<@&-VS
aW:7/6-6GW9QMF[XgHNRO,,@Z))f<7RKAW/.,a@dU[/_B)^(TR,XS&H0,Bg3@9]T
@2K9J1.6cXJX2KJCU.Ra+PKL#;WF>D,YC):[7U>;>GZQLF#PN+1V05H;]9Jc>,NX
gW-9@d.V>0\Z.75<Qda.^EZ;VGY^Z5a9&:ASU6U-W7]eHc.VaKGRCBUFPKIR(0ZT
fJIJZ<c>fTc;@Qf2)@gLNYB0W<A&CCDDPdg>XQcL4MWbPSGX)e-3A@HH8-[#@E-c
U/&ccCaGI3U@=JE;4A(1aHcO=M&]X@NSWW\,7N.Re.VB(LD?)FWPG,BaKI0E)>c^
ZNNdcWV6eBL5+1.X.>;ZS^2IaT.M?X>/\bA<CA5;PK\gQUE>+9JC[g-B^<T_--I-
PG]7Y[Z/=4&8f5&8.BF&@;cVZ254A_-(\Zb]U=M+0H\VMALQ.NMT<8O0eDe>-2E5
MA9=)M?g6D=@eMGab]Q#9(>a;:<PI2Rb7A&SQNV@P5+-aF:?O[7&PL#T0)>1gBI1
)Z5]_]A0>0KC5)ccX#;9W63Tba>FFQ?SXQ^M.O_M,Y.37_c8@ZbJ98=-?)O)/>Jd
MT31]gQUSP--8R9NFK2+2<FXf9=f6EK_<_bM6QEC#&RD3E,N+b,VNIULH?7/(bW&
a/@:L&7C2D7f8:+9d3cY)EHaZ&=AT#23S=LZZ=N4-g5WP>=e:Zb@f)dGGcOV)WBe
Y>8c.AP(/cT8L8]YFLYY;@3CI:_L_2.\d#W,7ZGDJ.\6OQ;CdI/5P;L:Wd&G5D^+
fLf(D88IT)ZBX0]?&A,3If4:P2T7]5T1Q=5;(6S@M\T.C=G(HPT6\^ZZ/dCEV:.Z
CN\3g0E]\;;5]]I:a[8+EV368QL1;9GP0T)5?#J#56&SY>I^Fb[YI]PPVcWJP<_d
1^_F.E)T)PaW+IUVd3:Z\5T9@JJ<6T@:d_RR1e@<L4^bKW6CB&F4E\g926U\BddR
,O_f+U55:T)1f5J<AQWfM<c=BAOd9=1QP:H-0AXaQLO;\E4daLMC8g7)e8;(L8P5
Eg8CT)&@0V][b+ePc>QTeePU/JF<4K@0OO>24FKFE1Q6_7ee\F2[E=?ea&NE<NBL
JP35e(+0EaMV;PRVHJO(b&KP),I-A8F\:(JK<?CV7L5UTHY.-gN._YOAf_@7,g4_
6#FbO^XU/9^PA1^g9V/YOHD<-fDSS[L:Ta,LDf;/3;IA[I3dPB/[:_9_Z,a&KBFG
X,1V@ND7ON;;XURS8)YQP__+f(ZI;63#K>9KA/8F/P()0F,#WICB)RcO/QXE9-2X
]HXcSENcE@JF_E>KdS2eB7N/gTd0BB<d=AgG2G72E=H;3W;f?CLBWX]C#4QK6QUT
B<:1WKA+\URTFKCU^g#1IeP[B,ML1/XGF;@f--gP:N04EH#YO1Z23g/EX85aE[SF
0Ldg^S^8f5gT_DK[b]KR<]9TJE-4VeWH7[QD&UaeU>>=<B\NQ??&[WLV\KMZ7e_)
DM0&CSCc[?/A2/(7);[JTcFaE-.RO92UPT2L;E+<H33.[G/6#RLVO;?5NGTVK(NL
L5=[:I67):95@L>b8IgZ7ga#N2UZR)YSHCO[9=?48DP=&&ELURb1^P4?^2?O.Y44
@2YE)->#?0GDRH5;C:4YS4+GA^HfVeT;^Sb^D#[XQ.EA5-?,QeYK^[G&GI+a[5OH
4J<D5d+OV:+f9M&=dM>J<8.eV@POI4fc9R5aVIK.:f0)SV8?IH=^0GL9<_L;MUUJ
;(LM;S8BUABMeLK7+bPJ@=Q<H72E_bBABEQ@[4QeRWBc[CI76+2e36#Ja+FH8&Rg
;5Z.EOJSK-15&b/.^Z_8c9GZ<::29R)_;#5fVYd(E^:>#]eEJFP&-RaW^F6\:8QM
K2_8&D=QMWbc;1eA^+O5fWg()E-bf(dBI7Md/eD?.6L5/]_C&JK6dNODL/Q2)-\a
^E4JGMcc6XC<9&&6\RB=^gEZaAO^ZW#-/aU26:I(@4C02&36dg#W-6O#I-8VZ_ga
cdVH8IG?_ZUMdJ,2,e\\Q6O^0SaT05N>-;(AX&7R/CY7W?WP1&@+2W6Z)]]-&.1)
H>O.2N\Y>92LX7LLR#RYD&NO(4UHTI3a2K]8VFg1LAc4S+O4>CAgFbRY+.-&Q(Dd
<(5QS#<<<DB=GKV+.J1TDA@?Y>3L.+eGC\b/f@?AX\He21O?3FKEE25SKUBDGfN#
e]:3gI+=UQ7bX3+):/M^3)RL206:Ied+\BJ(]0g0<C7S^4CX<A4B+5=I?A(98H[7
/Y#L3aP3;<Z8:(fgI,WP(45)K^+G#P-/b96([SC7A[Vg.D@HP@E4@Z6(cK@,Z<NZ
HM2I<<?[_VW;Sb.TXeT+Z7XUa4Zf^gc><$
`endprotected
              
`protected
aX/e4Z[IeUC46N5L+5VUREZX4>ID^3P75F\Zd-H@Le>VC4eV+91&5)28/c?e,Q[X
A+;3PA5FYW5Y6)#.4Z>9N\OU2?G3IbP5_\L]\(.1T4-VG$
`endprotected
              
//vcs_lic_vip_protect
  `protected
RB-W9PYdG:eUC\_674[N/b@OZFK4AJa?4Z[UJWDHgGdUG[0W-O@,.(FKLMQ?)3JV
_;bP55ccGdL[C]/2RCN3dY7=UB10-D^[N2AG-EHD]K7MEI7[0cXJ@]G=5^-T+/+O
M:7a7,60:W5e)dKS8^#d.Peg(1+N:M2/,_M=]acCA9K+)?F:Q=]>3A9<XM3<X,6g
;>5(FQU>YPE=+42<LKFI@>9K:GWa):&D+Y/.-_gP<WHCfK<c=ZHU\QW[HOd<7ED4
FJJ5LD<6ICF/g^_:4c:.fWELOO0I?C1TaP5WDQ+IF1R4egF_M:AdS.edUeae6HGe
U9)\W+^,Hg7Mg,MBZET(13=/2DOF6<O^VU<(3B+.#P9>PP0N/Z/+?&Q.Q02a&2W@
@PL;9KE#S1Z9A?8fg=I+[aFO5<#HM0MS:1U^CHT]3AaL?,+Ld(/?)O5:-fYQY4;0
.QCPV0/D(IN9<FZ/M8YN>g<?:M+f)X>e9+Tc]dL?29bQZ6<>3]\aXO?H#PdY>a0a
,PCWS0_.5MVFeUKGYUR[/-\QS0?#XN:D^\D6JML/Tca?^fXO/1/;4F?WA09RZ^1U
;3J5E73T)-K]:C3XBG91<Cc^<@ONQMeK2,d194)Af\AG781SY=PL:.<:P)D[L(FM
09VM73>?fPVD<,PJ(Fe;?S&?;FRC\E88IV4\4=EGfcV9[H_[gc_BO9WEgQI:3a5a
:a7PTQ9CCG3;:;?_B<.8H2T&KG6>C;0XAd.U+(^ALOO#@@^&N^_]AMVP=^gH<)R/
LdVUDbW6/#EbY:G<&IW-RJ)[Z>=e_OW2JK<;P>#+P)F173YM.0[JD,;+d@_<CO\]
F#-H1NNP0>/:3A,c>7&+INY4_&/]^a_)VYY7N_bKFF)]J+UU_#=JJKT?YI4&3Q-9
8&<9XLegO=PWNQ?78N6@&\KTXZ[;P.AYTXK\2A-59/#1ET++P^N[b@@J(;I_/PVO
dJ=4DU([)c8LZg&5LeZWBBUe^f)]EL1,Ac/L)R4:BdNN1.2.CE,[+e+@J/QW&Y0F
Y81LQM.L.U_^>g&;.-/6PUA5;FS^C>VgT_,eRT;TU2QNTD&(Y&NX.[YPKFCYEV+(
F&\XH@c[17GKG/[W2SZ>,VGU&EBaA^GD58_OL=.d;]B,H\d>SE@7TdWU=#a6g/Y-
3P@P,V-KAYHCE<([,JTd7ZVWg2S;V3-M(@@Bfc-DZFNI:_NARJA>RE\RYJ:9SI,G
&AZ+DNLdRc+8bTZ>g5ca<[c<\1dY+df(fF=]2?:NcebR9L[9)WAfM/H3QQed+8NF
@046IF0M9HWX&Z6=1c4DeD3@\WZM(6@Y_T.EM>6R;Y.LgZ7fVLaPN@b^RddU[\^F
+@INI9DWPc1fT\2[f#(QU72AdU&L4]L\9O(0&P0NC9W?f=cQ7(KG4F3.9S8L7EcL
/,MHI]S^OQ,SS2WSa\^VT?UZGO6b/6EEZgT[RePELdbG,Gf26d4O&ZI2Ag?K&-1]
RYJ,2<[NEHRQRG+A\b_8,)W_KA9MN>Gd^EPRgA9]\_aXT.T:5[d(?#<eC=JHS@>=
LPBOU\VfdAYO5BY<5/dfYOM/>^JZVYWKNJDL\Q[3&IBHG&1/IY[g(LW4(]S71^60
PI>^EYf,_>5OcG8-OfFLcO1?@VYF@/>@?AIg_MA8:DdE^,C;M63]GceEcV.+L#Kf
_7LU4,-Q18aMc7:[PJ?g7>Z-aFJ>E<JM6YC-e/M-R0#?gIc7&I>BYJFQ?g#UFN]R
?Q&YUE/36-(X28RVF8SY<[0Ag)U_RI&;:2?b)#c_>3@McJ7T3E[>;CbFcS\\f]#X
XUC5^G)7LP,W._=21<@^QMEJ^#PZaeEB8SEHe(aD7YOR5SDPZ:A6;=YK@S7T[18;
B6C/^Y\>RP[]2,DG^D=K[G\CaH01.fXePX^&.\VV:N?NCDdD-/,^dG??\T2Y=9[4
R(MN+cA9(Z#=aAFZ@#9V;[gG?=;6=Bd@#/UJ&+]VD=ATBSXJ-&+3]H,R4B\..@S)
S9aYJN0c=5N^SH,Ob976a3SBSKA7TPF-0_?\=9C_R@V=>E)O7TYP1LE+]8-a7PC]
?B@DI?/6;);=/6-d&YQMK&1CP??^CX>B4&Z45LQ.c#^9PK4SNbgSAT]5<^_3+MPe
CS-X1_P\d#,^CP-B?a-,fbBD-,[LO8\NfVV#B&>8#0\4&=.4)H>WR@6.>Y7?(bEB
_:6=YP)G((1@_-36,B84[a5=)0;8]L51M31=9dM99(,ESIE]0O8F3NN#[PI(@C28
O_bd#OBdKNNga.+/-B9):&Zb,6KSTf\4>bWMK@V3d30LPIVI<:##,[QJ_adGA):f
d^?V1KSZf^3S<#[;OPB)QeX>N]3[(eB5<A=KE^bDMd[G?Y:6,:?P#@4MD?TWXLW]
^Wg,-WZ/KQ6V2g5gfJ3f0-^&T?0ZRBF>fb:5K^,<2G-&C?753cf(:0P6,VgBdF=6
SZd]ca=&F(;2U1YT#eC(3gNKG,T2dYdYF&G2^+2)=e+8S,2R\2af+QaH;a?aYdH3
JJ(W;YS2V2Mff_5^-Y;+9dbLWb7D-5]C:5BS;^@NdeN#0U6K>1H8694[dBJ[L,1N
HYV@&V+UO/80L0^6>^.aV(NB2\,>eXJ\RR-P56DO9SA/0gAE]ZaBPX)gDS6[T2LK
5=NbA6=>T<7N7ZHWIJNT(P[6?)HM,?5[-\g/2Y;T_--==\5LfYb5RIQ^b:fLAQ8F
b8S:6Y9e4UI<.AKLTDHT[fa4_@^a=7LR--XaJ)\V3I;b)9.MVXCPfbdX&Yf=[^+Z
8P+ZM+AcH\P]6A2]Je0(7T+W[72ZWQ4&YdJDK=I&J_BcKZb-15g5Z\(C8;@#_4F.
+7;Zcga0G4c[KDc.DS6,,?<_\#2\,fCKA#09HB886UGT>a,4M1^df7/FaZ7Ocb1D
a,_FC2b:_Z2V&]eR8\3OJTebDL4IQ^[+U:HNcU1/4>3M\(T],G&bDEE9SOfcGQfN
]:Tf/N\X:-X]HPPda-RR[2QH<9PS2V26N9.U>Z5MT^M2SF?3RQVDPf&CFVH#(^TL
TYG9Z^=+YJ+586c)#W,,OM_&4Y9-P1BW7X=@,8F?;NA/6G<[VP)_b<3UfVF;8\B3
M/>c1Ua_L-[Nc]B_S:UUHQ&Ld,LS8DR[gF5]&F5c4+5PH/HW5-]aN4-:7&FBD^Ea
=X2LST^PV-=L2LQA<dLQKeCA3M_AORF#1)ST(/0AHHc[,+fAC7(<,V[Zd=g^W]+1
93,eD686L5HP=QB/70IYV-V=,>#98W:U/(=ADcd7U5/,Ac1.IMfbY=dK4@8YXf>7
4&eWQ..g;IJC+-^S.d5]_#8b>gPF];@a[^A\,S7=Y)beRQ_WJI?8;IW0EZTdUO&C
_OQ>MT]Z6:NM@RL_3EWQeF)N+;4ZK??ER8@+cA<0\UAT-P@4eeZM[b9KY5LS2I1L
2A8aW72#8OP-WD2bP2:55C31IIeDR>?J.70\F=X2W0.9aI#8FVA)._R2QQUXcI2V
VQ1dQN0]O-5H487)]>YISZ/;)79d_2B0O;eWJ3F.0G\,+?V\b2=bT\)7dZ6\H#V9
W[B));.S6EF+)T=0;Qa9^L0dd_<U?:T@QM;Q\1BZC\,B7E/<]4Z?G2CVX4dC<3O<
WI:d<158a-gXE+OU-FE5<=S#@3__KBC5d,T6-3/\U0+HgBe.&0.W@XB33Q>M>aYT
@W6A-IA.\gOZX08;5P=;6bQ#O#-74BV&.=USIP-S8g??P72??@\CeH-_28\M.>6^
a#RE^5=@4=^BG#D\#ePI3IDVVG:)H^/CB?28@,WI]3X-IcS31]#L77]S\EJR;Afe
#;_&KMU62db[KHITe0Z[_+LHO94;-5P66W(W_)>?L?12S_g0ddIQgAJ=7W.HV?1B
?^ePJ;#ZGE[U2g7-2VN5.SRY(1RZH?.54[CUeZ6FAD&^J?Y9./+;F],VBbJ=BQ;7
Z86[#1F@[3Cc^T.V,V2GY]56=E>(R)@DNWQ&3QffaY?5WT3FN9;<O2cfKVCR2IB0
V2bHU5SI4DRB)RbSa#O1\[5>=.D7a]YJO#_I?C,4Y;2I/b[deF@b_GQ@-PY__VY?
@Y=L_:];]CB]/4KMUW9/Fa??f&AAGXVaa1E/f<1^M:OW&(a^cXM_b[@CXA<2]4D2
PRR)Z6E<?<(.F9_G.Oa7,.SIYe&fNI+d2P2PaKB(>RAK</]VT3=_b#HRFPa):R4c
5c:4(#ZgS;g9.)A<5N^61+H=DcUAE[d3cNLK30Z<^M3AO]L9aFOE==bIf#R<f/Be
a#_d(U1:V@.G7Z91(^N?fS7I_Dg62&D.,K6ITJQIHff=Y>ddCaA+DDa+L=+e7#G+
IAGLa1.CS(?=Eb)X4aIO==L)#E[d?0BQ\ed9^AVUMS1ddJM9(&#B\\(K_d^A2Z0Q
YXHW(VWd4#I(^R?G>.\IHM4\(&,2]6<JA55(c,WH6Z5QE2EV9PJ\1FQ/:5Kg>K6)
J_P/@X26)/5S37/4)3T70dbF[c?8F+^A6B9+M0ER^Y0M=c^Q;^VIC:7PS#&67BCH
KD?T8[6Zg9^?1+\.X2047(GGMD<LQOEHaf=^2_+ee=bd,[&N?WFU@0TEHgbb9H]3
?+89;Kc:WK@RZY0V+./]Xd,J8,E6P7NP=7P9C\<7b5AE)X_)?HUH]@5OfW^7(9@T
,/<25FRU-N2KQ#([(eU9Nc?ZZUdA-DI:0=df..6AX/H[O;]2RZV\(OD7Y8?A2YU-
Fea1A^;X4\TUP+-:B.gN[TGb_PL0TN9?X\B(G-FEZM/<QPSP+3IdXVH(=+J3[11M
BgS3]XCT_cfL\a>R[D#FI0-AeGSB+X<aM0,8dXD=bbMY&\aP)MBWZdV/XFNcC(gK
,eB+(EFR2#86YKaN8Fb:b).^JRcf?3eHQ1gH9,D35IL]XV,_A1<O/SWKG7EK@,dK
5X-HL.4H=1F^KYIdIK0+^cFSc128TgTVJ8_e2Q&gCg0E:VKJO[CQJE:#-0:X25Z5
W:,G6?W2-;0=93GS=GOadTAS3<]W59,&B7Mgg]g_IBdM[c0-aJS2(S2-:a9N[d^Y
HN>I.M\QN-d6J;#713TC=CfL5U1YALZRJ+\e+,O^(6eLATBf9T7Yf\dc;7:UeKOM
D/A---SU,7/:HXD9XGCXZ;?FggI2?22^&:#D#C8PTY.6-V>c4a31FdRKfNVQ5.2F
GWOX_6E3YJbD;0KY-cUTIDQ[V]c.D<JO2E;_6V0=GZ01Sb83>fOfG##cR45RUe6[
9/62MeI(K+:0fP<cCU^76YQS(WCS2BP+-R/B>GBQ19#FHMOd=^Z#W#6L&<9R7I(A
@#9&&LQ6bP+d.9_0F/YWT]Ad.6RXJX=]1,^1\P]bTg,S,NW_&A+e154.1&U/Yaa8
O?2gDNILKg,YX+M@3RQH3?;[I<2>YRB\YUL_9e+]U/,Z4O3[ZJfUg[)gUW<E5dM4
JfF<^fA=1e:(>Q[+\=WU9[O\HBHD#EORJ6(aVg,<(c/\g1W=:.Aed>,T579C(VB_
6Q<B;KU@6F_Qf]PUeX>e/I(TdCYB__)fC_9[>G[+5B67KG8==gD-E\_=@dY_:Z6B
f0;,.IGU,D7\6GF.D#)<PR&^4[dS?TA,V+^e/^cV<HBPG0)GT<Q@&4>TVD3+WW;7
)#?&RI06c?RagL#[=8BY=d1]Xf9-WS4AT:ag_N6O8ZIge>6003<XC(BDG?g0C91:
M^[+^?5W;OE8[JPbMT<K5F784M@H:Z,c^JQ/Y(]fSCOQ.YAb1\cgJ_b]DI\Q(QT=
HC+GN[,^QVe-UGG<U\C]B5S7:0S[PQS9YU.GP34H.&CAcLXaZ>:-L@.TC)>[AN/0
/JJC[F;E6--VQ@CW?DV\I0V;U0BDBK\)835efRNa?TGP-^[U,((^BQB47KR(1,-:
dMg8@WPF@Z0T/C:V7IJ#)e6Hc=O9&80,)T_LYG,;QB-D<AOP_X3HNd:>b4?2WNB,
:K1;]dY>>Lb5SA;RGaB1a#,I_HFRgMYE?Aa0SB[S(Q.]Wa?W?DBR?V&[[FOf)AgK
<bE/GPcU:dEZ#O<We(-4B[HCP8T:.[&D#E0c<8ZF5#-3BB1TXa4DA_W62\YT8_#:
(MIXYCH98PC6-?5+1+<0GMN4EMbK9e8L4Z98SR]J)1TD]gI&Y9)@Og5PL_R,<P0T
D2KU0/R+PG^5[,V0XEKVM7P8c;f5;GXSSJG\c6_.UEKKW(:aX7Ta^eLV@A>9/H..
d]H<KM@+2cQTF23?dH2ZHJ[5/Y_R8YN/N4D4e<ag7\U(N:GV]_A9MNUV=DeI?C6D
>EWUbYQ/RL9HX?I+#N_Te&@@KN/(#Z,d[ZSdeWB5;N,@756RA\<g\UP\(@U5^0W/
aRX#Ve/??1+JcYC7#ZY?^?X9d+2[KN/dbc94):KDXXLQBE4.57PgZd3XUK:GdP]N
QR=#H;&b>NV9QD)fU]:((c8P5L5VI^Z77TQ(bXDQTJf6@[G6eM.cD[RL[GeQ,_@4
BM[:T<1fKa35O>1EUbLSaY[8.B(d=6:.N:1\8+MIX#J-KK&W9:4+656Z9TG_[.UZ
T&XK^-RYJf]M]SKU9PFK2,-:]e0_>PTSY:A7RAN,SdD^I>c6^#B?)bPfdK+_2abM
2/5ZIDLSEP[71.EA=X7+I1Ud>&ebPQF8^,:?Na)I2gY;UbL&/16G?/E6]fY25_G\
9(PU4e-X\29[FUD_,NPXVE3JR7(\DK=3,T_c--<W92K:[R+35[B4_Pg,H=C^dP#N
8&D=#fV@Q.1<_DF.G?.bBO^6\IBY^#f(4#5-8&Yc)B,\[67&gb\G9ZbA)-_1WE],
#4/,T_10/OVI0T+B5b8b(EZ6W4I]IIOU\^J^N+Rg:RQ66+9XNTM9;STDZS-cQP,F
_Z.^<0>VGR7R8Z_9+KEa##B)P3CS.V6:A+FW-L?]-Q;M-0+e3X.AX]dS]#AY7.+:
1I9TN_MACL+7CSHegB8BR8?ZZa)2Z85\0_XWFfOP[5:L:M,D]<)ESYeP4M@c8,>6
b4O9?,Y^^eY>B=VKM,_MA^Z)OTE4[c+]V\9d45R3/K05^2DZL<,8REY>c4S]L@^D
FN^I2:U:0BaVZNX?SLWbXJQ/T,EG>(A_1&f&Y09\,Tc^ZNZW+E:_f+VSUNg;4;RN
XTW>O:6WNg/f0UVB7XYNUZJF@TBVS_N)K/O;#W+][,=[./->L2fJ#<#><DDYY>aQ
(0:aN<P?I_;.=X#dG.]LU9.B?^X6F\J43&Z0VZCKc56?b>):G17c7gALOH(W@]^&
TBF\DF6H<FD^&@WNgYc9-MWg8e>YG00b-b54P&2Y^>YIQg&JK\XMLfH=d7YbII1^
7>JPQH1&;BZP0XaW)]aV=A^Db6+KTU@5b=AK3(eG0c84Bc;D&2.949=WLQ^>\OHV
E>V;eAP(=95Pf7TEZW/92b0,GTfgKI+_9FDe7N(/:4aa#gd&g#-E=X[.,[;Z<32V
NWW;(\f6<DASYfDJ_?4YZK=AXLCL^:D_-\b6cf2]Q-H>Q0A&;]U-[F^[=1Y,,Mc8
1:+9D#_X6caE<QS99C-Vb45OHLdXXG-L47Q:GKKA[DJg&:?LH;KFdd?;4__>.2P,
3>;F,?U\A<<ac.(J5537YTR/;TT6=JTUVagPV-H?1/BTgA8=U#,Sf+OP7.1O[&bg
.YT33Qf/HMRL@9XKWL0N999^51#e8]fIDZg?.cC,58<YKZa])-SK&-0\Dcg6d(=&
(+eFOI@OA.<H2;SA:2;-GP<Ie&\.[fWgdg)26K\f\RNG;=7\Z8A_Fb5K<,Lc>&>,
=7g(bTP<Z00N?\#I>O=OW\[8AQc7.=aVCbcc+B>\2S1)N_&e0CM;&T:5OFY0X50<
4N1SA@S3_eKfLP[)0+d]acagH.6^XL#3JJ&ONB;;JLI@K+PLc3Z5Yc(7I+dgB&TJ
DQIG8R+\+E^-JC9T7aYD4E&]J,ACa3>E@fTIaO4c,=[;ZE+T[LF=#B:N6TQE;#RF
AbAf,A?=#fc.N\;7JLa^:S/g0&<ZRWQW@YV>M3/:5EHEUI^SU3FV]>:5gS@;N>3R
XZ_=N6,EF(Xf0,bcQ@\_[/<JSCQI,1R5)EQDA)&93ac:R-8<<;<LT#-YfB97<D30
IZ_1?c<9C(/0aC1O64J;C.QO6O,ZR9B;GI&XI-/RZ@9CeQC:I/;<gfX6f/S](8af
0B\;NT<a,D_Q92NIAUYW35R2GH8?8F-49W_XLCUJ)I.f?JO6fKWMbgEMB^T6_)-C
M(XN)eBYafc&\1CbCY&<_bgDF\cOg&=H0(M5V/]9:@WS&aO5R&/MY<2SVV(1e,T4
KRE&W7JU147=S7&f<Ic9g<JV&g=_>YdfVd1+CR,T85Da,3G:cY<BS4RC^I=N31Z?
FV.V0(VMQ/_-.GA^d]O-c^T+V6.1]Cb:;-0_f4d^M6C,8d7CB3>2EaA,gIX,?PY_
?G4#1NXcLTW6V&G/5MOFK&^=]?[aIU4):95W)3#c2Y09-X_Nc>AB8^I>;WV=fVZZ
7\b2ea11F3_O.8Q2Q-^?a#+LIP,3?E]O+E\-2X>.+Og/1;Bd@=&/1CD]N4CBOCaP
NZO][QbU#VVKO<2_EdgV_NH0Ic+^+_XS?[Bc06(9.9WQc@#6L6bBIc<LJ9N?X2BG
F4-RSE^:e.A0c?6F7\18@f.e:P.90VV0bEW6KL3_&D[[@7g-Q;CQL?Hf5O0?=[][
YVYR;DD@-7fJ9SXH?GJOO0,\4b5\&=2;X2+7)1)NLA.U.Ba8WROOdP,3:)^QXf^S
cb8:29--@\H<F+D9_(,[dY2JJeI,+)<2\edA2T_9U1H^R6Dac/gIY5+E1AI-)MP3
LIaG6D6<Q.EU@08A<7O=K=AReV_fA3QJ-Z)].AU\^>g.?acd-b=)Df20U<<(4U<M
GcKF#J,&4C]:5F5KMV_SV<@^,=]UTNP7B\ed=#K\<@a])&X;+,8fHB0AP#._-?0<
DU/[4b>O5Pe#S&-I,P.T3d(DX8Id^+&fD&-UTGF/)Pb\MS7Ab)/=G#=D6_.?]V+J
TSbF;#8X^g#YfVQG_7<^g7;9BgRDXE52]ZB5[P1ZQI3G>1M.4R6c>9OZ[7c(e,E<
;\VgL&N6;^O)R^59QA,\B48D[^cDKH\D;b2_cB?c6>[E<OMea5g,g:,eYPS5A+5>
93V6>1@Y__D7bG9=.P]D//)+B3b\D3g\EQc-eQ.KG3=J1Ld<eU_6d_]XY,&R-C2T
?[GO.P-(gg^RXOD+:K@QTe\UV#8WFSI8a1&A=e+.<,Xbe\Z[[>CYg.(:60)6L_6J
WN>72FWK4@d4CB1.2AXA(0O=P79\25K8H2M1G_bS5d6X[e_<7Y03E3THPZ1Z&_10
VC=OZgIBZ]g@2YPJZO(>5:O^[N],4dTUR[:W.+B+8JAQFA90&B6J4G_8=e72,3aP
:cH<Y5M2ZJ=E?eH@R>DYc(NM28=7bM0GeWM_D[<0fcD:],)?;J2;[)1_P;M@/L4]
\,VOQf@EEVS_O+HgKQP?\,PRG;dGO95U.X\T-Z:::<6I95@F]1JXHKA^c[LX/I90
W2NJ-;]+?a7b[+HQ;&EZg=W\bZL7?KOfT6FARBWDN=H1,c1V&4S0>,,9O,\+FW@>
OIf<-R]6._ATKBH^]75aK;RM+a&G>M]gC^39F23N++IVX/aCdfbR--N@K2/\D5Z>
B2FGL,=&P>GB)JMU&:+.ObLY:.Q3MJ;67Xe)F3bFdN)bBO._BNI/a#;.aPgN@>E/
bK.SUd,7=MK.#RDRN8BHG5b;,LXZW^M-MLcc+?Pab&#-=Cb8bQG:6fHT6[>&eaWR
+afH79cC>9-V^2=;g\^##1C_#FK6.,&3H2EW.\c+c1b1Ja_->J5f.55=/Zg-<7Lc
fL@<;A]fJUY9;6VGQC;Z<a)I-^1_B>YEDa=bLR;[3f]PQ(Tb,B]>UBTB6.J^NNPd
MAA(Q2IOeL@a=E+BJIcLI^(LM=OCP+EO[YHYgcZ#Z?I+Q:Y09-OCMGA;V_4UE3G]
MM6P;[S0AbRK,]^@RIUT3N]AM?GMCXIfaH#-FWBWJ@Ca[L,NS;.[+?P,W#6a2Y&:
7G,YB0+6F,<]Z=:@+:2+Od#[MXd)?Q=&5Tg\M:5)?G1KKd,G2A)97H5LTY6[1QVc
;aPe[RN[_/8T//0,V+,7&c5[cXH-/5ZO6Y^N&7b4YG#L\3]f,9#4KUVRg<))/=S8
>a\<,IfK:D\&VG.<.(Sd#DTL[H#0K/A02W56QfD@Pd;E682c/5BW>QI02_:(.NFS
U1=Bg38G\(#])7aD?M?Fb-?9D(/bX[EHfT><XL7<g8YB55E@f)D)S3.:^1X9d_WY
+7#3M;:AI[cgHSIA42b=Z/-b40Y(?=>gQ\2PX(OMIOD6\1-__:d]ZMDc>2UH/O.8
b(;eOIA6e/;Ge>O)LIaYe_T?A<QUd#T2I7[980,+X\egaK^A^]:20&UcJ[=WP0,H
DNcV6=?\<LRE+-Tb7GW@7=&YUFSLE^(1/dB,O)SI,[M).U^?]VY7IGD2U=5X)42G
YS@NC+S>:cI?A-O[AHK,e?3X)2:aFYHM/Z_afBB^ESER.CWT_\HEH]FM.>H^)OXa
(e[g,M0d2940CV:/3f9.D>QE+G,N2MD:R><&4OfeK55US\/9<gI-56QGQ(FE2MfM
fIVebe65E2RRFF)@BQI>Y0e)W.\)c#K<b^7:&O#V)Q]KSL=T:@738[gI-)II2&28
4D(>-K^2:9MID.Y]=/R8#-@#E,XG8&I#KLP5V0V-3?F?;;3LK_9-6Yc+?(YM-DR4
a9ZYNJf57Z\M1Ob9XH:=K&R:-fSEG&-]?gL/5>;_1I;DO;f(X7<&M[U>224EQf:/
E@N3+>K4W\9&:?RaD_HQf+g^eZ_MU1XBV5,\SI&d4W)M2f[,_35\F/B[JDIDVfa:
W(]Y_,THSd37E1#BB\P^&TSL_4_Xe(^TGB,)67N,N^.T5MB:2E:6]URWJN[^Sg1M
/g+E]c2=\J&fOa6,eX8CD<cJWF.1Y/CGF&eMH9LOA<WLNJR[Y:\FO^F-e.._=BgQ
Mef9ZF=XLPZJ:\gc@Lf3B&[E\#7UE3X5.WD89P(caP6M?c.27P+7[GKTU]Z,SBUV
L\(FF]3.1=Y5edY><KF>H3AGbCZP8JBdNU@=E6VN_PE=?[ZCR@KJX(-^>-BR3.;2
[?+M?OYEH+bUVI^[14d\,EG?4H0S#D9cM_Z&LV[_.TIL8]/\JPSCJ;6c@P(X\Me[
Of-gSHZ]5+,3cM0Z4O]O;;\C3)J1:^DQYKE;Pf&;O]T=[;4+OR3<\P)J-_L8OFLL
58SC^/HWa]e4:c_6Ue>BadA@_2Zg[4CHFG^eJ:QII7+^9c7,LV;^M/GDQSPT?7_A
6//)F]d=g[.351aTfZ_S]WF1&C#RW>3</1\P<>1BaAT9X(I[7QUZQ1dTRY=f21\&
FT/@E=D]CJ92;=cSg?:9N=HM:_?d1[0+eTHFd(NZEHBEL13?C^79[Y=gPGN_:CCg
4:Kd@_-R6CQSO5fA70=f=ZQ<FaXY.N>/#<6UX,.42O-QOEP>_aI7cL<dbIKB)bZO
L/Wa/W(R]>2g/9YNX^7PW>N@C@)_cZBI]&ccZ,XQ\?Y+.F]+H\-M]W6#HVZD#,YO
NJ1NW_S1L65b;?VJE539c&_H_ZeL\2=LYb[=B?88?N@JF?#.eZ6?F)aaMH5I?:12
_.bW7125&Tc73gQO8#F-8P@Od&J:9d?/I<;OdS(90c58EF6;/D0Y^NM-K+c:KW1F
b>/fR[_4Ya;54HYaRPP<dcbP.P5EXg1SV2cIZOC5KP-Y+SO<).LKf&J28H>SI8MC
E8WE&6bX9]&gK&N0)W5II:=HcJDX_[ddd]ZS<]TdV/K9Hd1C.5CCBK\dH-;)X3]@
TQSW,S]DbL>>X>^WE54aADE:NV6TG3+W/-&WaQ/Z^ZA=KF:dHN]Ze-[&CdL1Q.fC
a[A(X.M_Y4]6@6[[bZ@14;ae1BBMU8:ZRgf&YXd7.H<09-d-1@C>He8B/@GVBdOV
+U7(bE;Ig)cbM-FRCb]R[.KVF,&\C2@O8G&IXTQBgEBV9JfFT_-#EM-U&e;5Fe,5
U:<eaD+WP(Z#UBGKRO6(N;2+>[[.g?eX4a3K;PK8KR0=MZ2A0L=83)],)VKZAMI>
-7C;+OUESTYHg<:0>aZIPaMd/;S9./+G[fJ;bVd\V9e<@a\9KM1021(A(:S?_63&
f@V&^gZH_Za30:-[QC^Cc#+FXf31a7N]JDdc0LK6?Zc;=@&4^XS;>\&BX^PFUD]F
2N-_I)]G)+);Y]gN\1U=,?()A=H^#,M-6^JN9P7+<,.P<DO<c;:9(VTc=/]9<4QA
;3R9XK^CI,AJ84XS)KHH=c0830gCaI?_K8RPNJFO55?dUIN[92)RZP]2eN+.,BcM
X>>9GF&4AKV;&.=]^FYHYQAGQT<&(8G^X:dU?Q@CE:VR#@-SLEV7FI,8^<M=X?0C
16g-dTX+GFX[b&gT4SAQ>;17>YH+#.<25-VITFU2gecW#?;M(,CF,ag:]@/c6S+2
91NB)PUS&B=I\[.3_ePd3,g/7ECQOXEJgM#J83,L3N+HFXPSbUT^6/G[b+@2(/e[
&H9\^_fcAbQ^O4;J\(#4-Q))LJ[)91NQY4?BR_A2bN.da?1UECRSLUe&bV4-Y0<E
AII_ZXMb=_XSIY3=YT>RSHU0D/J+H81GR700:1<D7-9dER(gWg;.;-QLLYbSF/-^
;?b^?Z&R8\8?36V#b\<4MJ@XCEd[=5YFcB1g/PEU:@UO6&cMJ\a3e8^IfO.EO#a/
KI_NQ=:J44A(K0a\g]7,5;+/[UV2,Me,\A9VACeHdHcFJ=?FTEJRZ2I=SgTD@3)-
@UGFQHB178SB8L(g.+06>12[3S(W2,Sb-Z^bR5/M+RZBN@NSW2:;2>gT94f).4:5
E>2R]OZA1\a2HQ&3)ABI,)BfT^ZBQPH<:1RgQdSET\Q65\.VUVJa0?RgG,K2c@_&
UbAg?=gBLf+3Z;]5WYeS-S3WUT2LeL^W1L0S\D-HR#A.H>bNNT_YW2+DJKN,99\5
bC.(B8Y-7F@5.6>6I73>AcZFWA2&+e6e:Ug+R.KA0)UV,9[D:JWfU>,(\C11/NaC
HD^9b+OGI1X;HLGTAYBP;f+YKdM?B@PfV2:O(4P0<0UH38HCPGfBS6>O6135_Z2P
?RT4P@].WM_\d_K+28FF7Zb3;)6LSK_;WYGY0@b_N7,W@7[8Bd5eDLR582]gX#<2
O(,L-L+D5?@(#-&VON:f86.2V>?#AVK:JO.2:P_;PSOU,;KBc:6_WDceN]RXWI>R
EI^Ra4R[A>C/DfFf244+WO:+?/OdV/I7IS6Q3&b&L1e=Xe)HgP<@9OJ&(M3cUW.@
E^<WXW^?4]SY=_6E)E@5YAD/C79=DI(fC_T8f42:H0ZXH4]>M;897N1?8M39UaJD
DA)6dB0?5F?)B_,3YY47.>SE>gZ)E_7=E+FCU^YX5(:<AN\]L@MS1aK+GM-AcV5d
=I:eCT)A:UF.;D?H@MEVZK3d0^:;TW^.e6ag&f(->f&\JSd,292>;a@02<P4K7EL
+Ea\[^K16ZAZ]-g_TSO-XM#^PZ&(&C1QWXOPN7CK?#S:XebAIL0?U-VTdfR4H/7f
Z)>C#I29.ZH\U_T)P1W8JMSG9?@3g0,B1\[1&K74a<:Fa0.8ND&/.F0f(]:PD;@K
@6@6QTbI,g;c;=->>eO@1b^4gIG87HZ;AaX2TVS7M>YR4dXfCH69Ig?Y;dOd<GX0
M[SW5RFKWd>I^e\O7.597JUSZBGeLI3@\^0C\CPB?;,RHRW926&6\TKV[N@9f;G]
1>WDSXeaQRXa:H9DYO7P/fT&U@J)d/T31Z[22eU:bd:2RRTECBQ\+Bf\E5\=B/3?
W,(#e.F1PLbTbOCGd[QZ+<:T8FGD3W5G0V;@99_[GI?C1R]c6Ef-V]<O#C=Oe0Q#
@)4<]GaEb9Yg[b-\9OTE;[L&fY_52e[&d9a&8-<^b8UV.301K/MB<7S3S)HD5>D5
(&UgJ=07bAT/U0PgZ,\3;D[e[JUQM=eE/B+1L6@[@E7#O\?\+)ATA_7T14JT.2fY
A0/2fI-9<J/5D)VOgXY10W_&#;#2A)M)6_<9;]LNNaU)Ke-&a,a=_Q;85VB)&W-P
IAeS@-&Yd:+4SZ2Xb3^.;8E@6PTWUBa_C\@gZ,5G3K+@7UXB]O_9V6N,[(2(1K@<
bgK)+U-F_\>J+1EG^DgUP<NgI7d4X:9H^cHBG44X]D.=Q^bL8X??3.9N=[E0+0g=
FF\)X@.Q?M0CQYKF&@/b:(8A2TEcSMF2=C-23[H;92QXKOAJ[Z5W_Y7.3Y9+_4^O
&<M6O;I3OB9WQ3;(bD66I((V<4Wc:4DS3e<SfW0]+=15Nc6gX7e/N.#>3<\E]QM.
gH3OR(#/-A<&/6S(Z;Z=Q(WC\8FdF6O<<f(a+c+[06.[PESY8IbIgZccC-8?Qg4-
@SN?FB:2cR@4M,ag@R9fQ4&cQVWSO=DFP2^H8?>R;^.3A8#gSD(b?M(]fbLbSDQB
2LQBK-X/GO9+\#ge:/E)Le&U3>(+-8:Md&SA?FSWX<?U^YI[^g(>K?HKJ-Z05G6Q
7e5T/a:.aC<5aX/^R2gX87FY1gNP[1196bXP#.:GGF.5NYcJ-ba1?g)cf5&-8/Q]
71]33PFf16_g38-Y0^3(RSAIU5Y&0ZW>[_(RS:N)LR[3^&7]D&^fMJ^R[K;g<1;g
U-1DQ9/T:B,eF\J7L3VQX?FH4U#/Y4^[2Q3I;EQaFLW0A>#Z-L\9bI=.1P9,WA26
FN2&UUa[Da#Ka.V^)f]1O0K<CYf2GNX:aDY+1GZ((N?LJYP3Xfa)eI]W1Q@)dZ9V
/>SC-O3)Xa4gK9aL@P&.Id?NB[c27N,Ee65HQZIZV]5F8[TLT5Z@9W.D?MC]K/@a
=MUPRGY92La4^I@&+Q\3YceB\#QOJ?\[\GE+VPMgNSFIWfQ+<BAF,57.=#>V0J^)
SQN@^bg&NBJBE6fIL-eIQW&N6_=F)#^bM1UH8g=)1>b(VAbNcd:5Hf\U0._DR)VN
.gSYUTUPTc,gE.J389MU]0]c_/=F&<?KAS>MfAe\BQT<P;eSFQ7[7[GWOW)^fB4X
]-4A#L6\+2V3:Y4_QI3Ga-:GVPG+DK@cDM[fQ#>-C4T)I?Ba3H9YAP7)(I?14PM1
4M5&U?/)aP_YbS7ZNC>?JGb?:D-1F-77XO<bNeJ,VeSXQA11K,aHU62GI-J7T9^Y
>J45N?EY0XQONAKD@BHMAGS<Y-<2d/PaM@G1M,WcG)@f];6?.aWWEc+:f)^)f00,
T#KM99@#7[,MCTbN_;8YWc+f15EGKM#WZ>^\P#SF^&<fc9IDN8F11(gU9SA1]8>[
J\QUg\70,fYLP:0ZSb),L@a_8d@8EL_Re\2\CM8@LK^3e=.LMD_U5XE=T3[),VgD
(&4AZ?7<<Xd50E#3]&g6C8IZ8NQfEB3EI\cCS-Q&fT<<G=5(6+]=KgY5,Gg]He5)
MdV1+JJJ];2@EZbfDJBA@+:DGXO)^4J?PS8Y6#.PdJ9X,5Q:7IN+6L:)29e;bNT.
S?KR1@4BM,6IcVYP6K(8SY1V]QNFceH&UTK,aRH8N+#O5-LU(6IHV>10EB(:BUE<
g3:IJ=]IL45GHb@b?,3GP:UE&0g039P<^[X(aC]O[Rcb@K<RYaW8W0#ET>_EYVA_
+#EPD,;bcMQO7>Q)J6,L)eX\HL5>4)7>@HeUaP6?77?HDaJ?83N1P4)TOeB;VE?a
9+<OE+.bU\)#4A9>#?be2^\5X-=>&+0;9<^Y.A2XDOe-^bP&=Y]dF&5&IRD/SO\7
D_8-<7NY&eQS51BeQbfV;.[;Zd95MBDcXGOYT71@1MD:9d8H?3dX8f_+2c)T3HN=
<DO3(O&0MDdP?0C^Q8>24\&L>)&<7OcD>Df,#5c]TZ12^EGbI[@GEU^O[6&AL(=4
8I:ID&-f#RcF)6dN>>[:LFJR&B#&WeE0N_?(NPPe8T1[?TR<U>R9NC;9b2>[FFI:
H_K3#5L;Q8KNP1QL.2&J3K32JZ@=d9E<Oa7VC,+Z)b3WTL2&X8BL#JFd/L=[@GKg
SQ1)O>3A4PU3YHcFWTfI>/2?#D2#BN+Td?d.#<#JT/7U[P&.]9;\PRc:)T-^K)(A
81Jf(5F1OCPJXgS)&\WBYNdEYSXQ+7OAH2,JA/8>#GY,>_?R8ePQ@K9bV:):=#dX
>VWb]Yc8R\KA.3(4-(=<HZg.LMU^?\Z]HeSTBYRWYXVYGC\9]@?BOg,U;L\-V]A,
g89LceI_Udd:4-@/b3]>M,4_=fa2Z@_WD.[?0LL/_BU>)>,CH_3L<ABg+G-?&YAA
I6/W<N]bOLKOQW_KEHg7M#.@</G<L;A<FPLW&;DG<:aU/@]OSJ@fP7LK=cYCA)\N
f[fQ_VR6Oe7)QLI/aCH\;b:1^LH68C37ITUFU5(fQgc]=&JNEYY6M^YR[IZMXNWT
^BDVZ^ab(3=CPF5PFAM>I[JF@+HIbX&c&F[bKJe2:9La]a#J7gE@_/-PCDAXU->I
Q:(9(4WN1eX@YgFS_W_)J+CPaYOLB1][_E5M:O[J;]gD)IdZJNGHQ/Y6JLS6=([P
E[,0ef\9.X]KQPI:V&aRNcaVD)C,bB.3(I\GFN5c]5L+\9N89:dG;#LcOBZ2JGKE
Pee^E;\UD2U=,2]PWUUc5<^?O]IRa1Q=YfN4QQUYBI<T]Sc1RF@dZ?Ec.\R)A29E
f^f&DSJA4G91\X+0B);-WTVVK=/0VE.5SW(<^ZdR8e1,J],B3)37>X.&B+NX.BQ&
6OY)Q?BRG>27e6e@(f)_;gacg5.>SO&2O+^cZ93d<<\XX.)9HLV@B(FUb>[/;G]?
>F8P60734./g;7c^??&[d]g_Wbf,^cF18<3IK1=1#dY5B\US,WFW@G/U=&+9gTIB
/+4L81dEW9/7g0V(Z5\9Z8:eeJ0HZN3:U,#8#Qf-Y]HAOPXAPN)J;KR#TFI,D(gF
R(LZ^:ZS]?+@SE3KE@J;1f>9K0<?-((.O5WK_ecN0UaQQI6^\e(ZW\)Z>K>KI[GT
\[cH]X0W.,a@@/].T]I/bDVZ]XZ2>LG:WM@GG0Kg69>08JRcGYV4Y_+b\=JRE/X3
TH.8PLGe99a;EV6C@Y0/7ZZC]F3Q>OFT#4X=+a1^OcP0gNSQ</-B<]f+[WEg.L#T
f?R>c86-JSJ6LH5.MV3\YB5cMAfC-/7FX.3<S=GeScbN#O7,E20C<OM(V5A(EAV7
e3]^N)5I#3eP-QZ7_&fH?ZUNXKfFQIB=WH<WU?83^1@788CAA(;X]fc8+G+V^BMa
e@=;,(d4.K^G=IW<:]O?G\\5&;S]EYD80-dDC;F>>4QN7\._fb-9)>-A0gSAAD3/
+Q\V(#8(@[4S6[T3>1HU-H\CEOL8)-G_F(O7;4G[-]:fG#A]M]9TXR_gK0JZX6Fe
62E)dX@&\\S;4L1a1\)+98A]QJB&M)#I?+=MYCI59R0b;b7NTC4WURc7CJWgcHGZ
4bfa@Pc_7T)/EF4V\)8(94MC2U:YWEGa&9&VLe07(A\3)WWWXBdO6eaU8E[G@a]5
>C;4VYC?ISM+-6Y\b)@K84&A?3JQ?1X>:@ONY.@d,TOZDURb-(\W+23\;.V[Hd#K
aYNLCd\T3AXPaZfVNgC]#Y.A(&15.MgL_c75);/Y#9^]&&>b9<=V4c+@WU]>b2^K
\(][UK6U,2U.8-@9N0+WP3[221230Q/G9:<FLg?<@?Y9\BY&F\UIJ>H2RH,W9IGQ
SAR+@fVc:-Z?\XU&ZXRDb[KL/RX+?5HLTc30QOA&]eZFb>G@I__;caCT6EU5_?.6
V6M:Y:FgJ]X);&OBK?L_b/1&#<D+]B^18;OI+gI+U4[(&CPI^db#7@e+7SAG?^FH
RSL;c;22O0?4C4AX0VY;cMbfVRf98N-?G74LM6XEGAUP?df:&cCE3W;N8-@?1X2A
A10K=0<>e0&^_+/5.B>7Y+fFKZF7[RC1IV:TgWR:U6#)YISPcKc,-VDVJ\QeV0X-
]H1SB8[eGA.KV5G:6ND9/Y\](PO9VKg,\fZ80Z^/WSd@Y+KaM09b]d41L@?F#bcD
^W-TQ[L,G&a)U9f-^)/)2,J=(HaYEX;WRMWQY:<BPb,HD9\dS[<MQffEe^)fHDWL
C9/<9-()<1=YXFP+7CCR6FMOe+L9KDF>.4eBZ^ELZBBSTG0dK([5.a7,9RD9KFd\
,L>\1KVM3_9K/PCJ+Pf;IaIYf/=G5b^Y&7cD7U1TEW5EJReBZ@:48+RN\FQ.GV@N
Oa:9Sb.ASNEKNS,32g1M5[.(X5UJBf7J9ZOOU&;&ORV#Gg\(B(7.MZZ#?L=.\R)6
eA/8EU4A,fgYCZZ&g.1XAf3Tc#IV\)B]d59V&##&8WFdC1ZW2P;?\fSU:1Q>DQW\
bfUBMKB.<S<ZL0aK:];#.Z[],B5]Bg+d7>2((B(HO+bfU+98MCgL(&cZIU6[<4bC
(3I,F72W^]Z\<S_aY(Ag[IB&XN1//f9LS_8dK.ZaK2U(Zb3UfCCb+Z<d5&A_c@T\
,MP440GE_MXd3NFM,b>6[TLaCX/&e,;O6X<,K@2_H@NU63N_E]SV_=Q;HC[72L&8
I^S?16HELB_fX6IK_+=QG?OGJ54IaHP-6WEg>SYK^#]C)-WVMf75:=E^4Ce;d#OE
b7aU4#>D?Q?-b#6#;e2g,\YWKTdO,E2+D]53T5OIbga\?4&QZ:Z[]7/MQZBd801[
CS0+TRHWP?G\e+QTY#9]^:83H/5Y)FFAN,R&#c4T4NaGZR\-602E[9/VNV_GD)d.
A\GKMV65>1_Q6N;Y)8#21M??gG=-AQLX@\>=P;(I&BfF1PKZGK3Q8<ZdK/])9O(0
C@G.,2W&/L\).]N1G@gMJ+H@#Jca5LV:4V4>S7dBCFJ#(XQ+)bHF@@fV@Mg8N3gH
;F+?MJ>K0=1NW2-MeF]5,5R(;57X5)f&5<-<E#7WQRV^&U@4N7?TF>0YP\-^+>SI
QI,-VFd)6aA3Ja4Z=CGfK9\TFg&Q>OV:OMYSbE_46e(TT578S,APWg<d)#;=IF1T
>]JT]^M3c3)KAVC6V\.g3=01;02W]AG?558]@gP;RRf#PeJ;]<E/O#f-47ALcFba
LE/Z9X6.@H38:9H,6(^WCbSS-+X-bG#@f9OVSM13^+M8ZXZCdLD-;.Tf_IX>2A47
D5e/3gYX:cKOU_].1MA;:eZ9e#6ADK?[5D>6;ENKN<CMWI?_W.C_].:T0Q.VE-B\
#5&>^4FR6N+^ZcN8_6./JO7HTTU7;CE=@f924.@1:DZA;URQR;&9[QU^YH)<+9\7
c-<:_c12aGIY&@J#5ER>g5#6W&:EULgFEE_\@(\B?0)a0fJ?6.KbNT>-gZbfIP(#
X?gX>H-D(X+0<(,@)1XPX5;BWHRO_^7XZYZ=(4Veec<5_KAg9]eYL-T5Z<UbO<?(
NBNX/6g;[Md8WCU4Ig7IBI^8P(/01Wf?d/:6X_UTRL<1GMbfFJ/23D9;)B1FF@X9
aT6XXX#Xd5[BN#,#[#&e^[VY?+eYQZ53L;P13OABJV=5/Y.f&f=K@Sb7QgN)e341
See,CS@W-ZId7Z#W;b8gD\_?>f2e2[C;c65/]\WMddG0.D#02a^[_9W/>aaUdLgU
QJ2.4I<BZAMTDfY,EE7ZFM@9OH7K^3TH3TR<7&Tb4.dAJQ1Wc(Kg2Q,@2V5;/4fN
WK/&#GA/];P27>RgE#cH5J]^FB[eC+/cdANRP6eQX-HbT#QPSZLW#XR:;):-M^;M
H=MJB:UY/^^4#,8VNKc>Mc<49Hf\Z<&/1=?X5BOYC=+E_cT=fW);^GIPL[OFdGV0
H&E9AA.Q4U(gHA0;^^AG5g3_H8R<9X_][N3VQ0^M:\U/CZ@-A6:FZDB2NG^Z.9/H
fN/3<_/.62Q<,S]#0A5@2KFMBHb)&M];M-a@&X;:g^,]JK;6c0860697D8CG7<\:
/&RaP42P(4JA,:[J+C6bMcH6f542:]Y14,0IV+WWL+0geW2(+3L)5:9I8^VdO>>R
e2O[OIXGJ1g/YabC1]F(D05P46ZSFWOR<ObC/:[H4&NS+NB0V4IW>Q06/2+8NW@I
^L3PZQ-Q:=>LXJUY\RN1XgGb&:7J_EaSU-gaR)IR4RcGRD<1#=L>6R<T\=UJ2d;M
0#A[RRe^LY-:UZ#UK=0T]8[UV7RV\-&0Mb&]W?SX.NfS>C(P11]/C>3DE<1--=a,
>5?>Vd_[;=dd^^_GVR#gDA/M#M:(R,U0?<&-V_;9.<;:af+I^+[9#_\@XS-6SfZ9
C?[+bN52N&=&47;+0\_K&>R(f7][1g2A6dFI07BY[XG)-g1_YOTRc#>=S(d3\abe
=KG@,^/EfQ7]ZQGA?_\9G[\NO[M&-g?37&;K[K,5-#&IQ]SY/<(?+1343IYY.1@9
=;a3E37H)H@0.b2</gZFJ^/&S+;.B@PYe:[,3.V0=^&9Y(R8N+3C_VZ00_F@8YNA
e/>R,0fY\QC#B@Q\]2JZIA?M\;82EgY]G<eI@>H0gA&ES:-a7?#9VR6L4?;;[&TA
c?XN4+5Y^/5:X=DeZI])SRf7[ZegOQB5LEcRF]-IE1a?X0G:_DJ1a727)]W@5(Z<
U4EBAb03GP9C>4HE:CHfD6?E)MEJ0PVOT.UCG-?+QCQJ)>E-SQ&5I.\eBMY1]CZf
)gGe#OT6X8TYOcR?-Eac[g3:b)Cc-,?:P25D^5A1/@faX,V-4F#ga2WJ3ZI.7&g.
(ND2?)RJ;.Xdc\+IFaXeLHM4f0@?D3=>/4WY+=6=E7<(H)H3cWWe5N\22?B?/84&
2CcZc,Z<Jdb^4RIJ1Oe:PDE,(<EDNW@0gW2/78cYJ.._]YbN>EV<O=Y^0XV50(.J
M7:Nf@0#HfXbBJOG\GaHd/10bBZa9W.dZAA7G1@APAY4F9dTX:,a._\K-])=^>]7
+EC3[5R,bM_LJKgN9Va(d@MM/0Jb1GUJ;Xa31/@1+-CHLIS8]a(-A;ZYUA?OZe59
Xa\@a)6+SL7?<5B58;E6RG3>?YGCR]Z;eJ.cMIZeW[@#TIRGO-<4:dTJg,7@D9bO
6,Y15=3NVYE:LRYSH;&U3/RL:[AF?8GMP9G\LAJWS_TD+=KJ1=d)JaJOXLPdX2<P
+g_2\S]09K,Qc&^3B635Od5\e7=\3#MHa;R)?LB&P2X4/#Ab6abaF+[g\]WM=0[e
SC0HNGN<YS\3)1XM6e.:1MPEWNP1->Acc+L0)ePHZObP,cM^aHO#@L2VbVP]aGI]
M7g4^BF5&dH_R;XdL?&M#g^2(#A<-4</2;S6T?FT:c&GGMS?+&-JSZ6P<=JG0VOI
>JeC&cP+MIMO9]7eX>@c,]DP<gFf0MIfVTEZH1-gE+?=J<A6R?=Ta456X\,;LH[N
>X&/f5Hcef-09?M08>g[dHUYS]3Pf&^Q\@cV0K[O5WC9V.@84\894KQ:g_PeO6.D
OUQ>T9KTEFJOC#XF,TTdXAaZM@SG[GLA+[_=94.(M:CA5Z/._b9AS>gdS#AgJ6>;
OC:e#_N2L)MCM&Te7F^NI6DdHHPIBb(?&(1B@Z-[WF85.-WcK(gB:_CU:0NP,5TR
)3(RA0HeZ2^g^_5S>ZRQHgI^0HfX7:=OWg3OPe+0+F.cM[MBKJ3=Zf0dW)OaNW0X
IEP6gDI9S6Q4?fH4P.A+=\3_,N+ZPQc[<ML^b4PN7:1c9GH1ebIZ_56WdbZ78(10
LLO>3;a\25de?B1QKT@:?O]_[M)?V1gfAT;LLSU4EN\&P8>gO@)<4A\MQY7+BFTc
bQ6D>EBW\bPDBgYe9IG\J_24Y#/K49SVb9eU]XPW,bgCBO_@-(Bb#]QH3F=_DYG[
RIRe]&C<Lcfa;,M)U:#Eb81X7NZbZ20A/e=J:SDWT@F55[KM:>1<;^GL:TJ>/Y46
55\KdAM^66.f44b6;ad>H<>]-TH]3aSVPKZdUGEP),CcQCE)ZZC9WZgIK7J-a+(Y
5a&DI\LBc05bMHeS@HDCWJG?[QNS481F8#TP7?B,]@R1<4B2VV3[38B9+ZI2Ra@@
5WaC([B+,&<N\>c1Q#cVEJYQESXB)3?\@QZ-]0a8A@9ODI-@V,9C51Va/7DL_K1(
@9JKKD90B.Rc:>XGb\;1F;QFbe7<+1eg5H&?3@BgT_J9HcA8K,YY5ERg:RB>5CUC
:9Z)Wa9F@:67HX^LeS)=N=3P<4)^ND4d;[&UFV5:CB50Dc8?]TBLKMbaXAc;_9Og
P>GDQ.X/gRX13A-O)B/H6=dR&PMKI+b+b[U=R0H3N#7XAU6.&eD,<dWTa1[f[X.H
b6#>1Z4DfW2V=?=DX=)TG@]_5DH5/d?8)9^U></3IU^b->O\HO8+;3T0Y,9UR^7c
K?@/;@(VF6X5E?B4MLPYWM#M>\QH@7TEb@QPO[>KVU@a\Gf8[@QfA=<IeM,LLKSJ
e17GCD^@V??<NM8YEP3DF=Fg_,-G#)[4[\+(T[^;^[PT0a#6H(e&=e\]dJ?G>@<5
-LeV+Dc8e.B&5/06S208Ef[_<:,VQZ0CJ9PT:QK+)e[VYCY/<GK@,#af-4Mc,^Y1
B/I_&+L/D?,E_]5-3bXA2AM=RVa(NXK&Y\cBcXC?^ZOB&bVI5^&gc?#IU<L=THd8
<=I@65_b(O[3RfFVd4?8ZR]8g)>A)9a70Nb?bFCZ5Ng[@PY[W\)PKHM3(cT2[C1.
>_P(5.eN5A[;5CDBKN,[4\4>AX1[Z(&^<6IS@^6P64V,LXTJ(.DFXL3T>)&>BfP:
CXT?eAeL\+aK51A:Zg)(-[]aLI.d]e-_4A+TBK-HG/\MI,_LCKd=8+:1H?BQaK?&
+/b786XVTC.57f;3NT21Z22Y+6NbCY=L\NM.aZ.+)M@Ke/d&FJ1/AXU0QXS&_H4:
T][A)?AC5aaB93&G<PPVJT\ONcBdT=_?K(.+-^B^eV:B?7fgLe,2,_a8TRX79;)I
<?DSI5d2=]:,+7fU+@?G3\3WRQEE5[aMSRfS,2EdN:a+P#[9.\7S7#Q#&A7G)2RH
TgE1U6(0^YQ0_?T+QgPV\2-aJ?-Z]OUbFgSJ3_VL>b@?=eD_HXW)&H<RI1ND>K7T
B):(38?8/<@.BJN/P[I1/:WQJ:E69[]5+>=C=?U<QY-@D5/bXW(6b.Gb?DID(FIa
Ge)a7V9eOb[:B;RPCBD;JLD0@&,K94#UO16-=458c5/.Le0Ucc02W:-FWSVIDG6e
H9.Jb&^1W+H8)L@+HRPJ/#W2f74^5dI]c4K>0a#bW]/Z2<Y.HTTKg9TJ:;^2YB_T
2<:-ALNV4/,E8K=4=aK?FLNKO9(OSJYAN9OS\0^HcWEB9@6R[0P</6[ASfATKb0U
SFECK+:PB4@g/O@_-^PQPU;^?8DOf56/(04O7HD8?I59]6#.]O-5X67[;[IJZGG0
;eN]f0/ed4e+UUEWaHCagBPW_0PX_K+PR2-Z/<^^[K]-W\GG4JX8(ZQ:)@H0[:@N
;/f27P-=f&D\e0_1:U^>PNP,/L&XE-+?/D&cF)gUMcK;26@1I&+O5gb?KQP9J9<3
_YGJT?caSPS&^+A]Eg:GaDV=dST8f5bY2IB(1>;c:eVbXKANLGIWee6O[CcXBC<8
2<S]1T2@&^/S@=E&;0dCUU_E,IMc->5;O[>G2Q+FR,R+?&R6agTK=T+PNcMUNHGe
]><Q?VgW;PccTBHI#5+A40,BZ;^e\cK&QfDOUc;]_L@QIQb&P&Q8+1\;<.dSbDVJ
<DIZdQSM?TIMgCc.9C9c>,#W8aX#9K=VY)IE@O5fZH-c2+^]:7Q>P/>DT8^1F_3,
1AZf:0cg>T0ZLB_GO8>U]BK.2>3Yg)0,0CTYEHTGFK^25QH2OWD\E4\NJeS/^a9a
A\2D853D07#:[10c./RJ[Y5#J-WF,ZeBO)874,=[aE(GIF3ZWf7=/@a]J>=7K3L;
J</Y[O:fH?dH11AaWP@T8<D43B0<QU9NWgB?X3<d_&Q\F9bVAa_D__1-dZ7CYb4P
A?:BP94T71H.VIMUV;MC9>1;336/cU]fIAGYV.=Sb\=[Y;?H+TJ^THUA]]07OeXU
=3GNV_NbI+E96C/bN06Q[P4&/-P)HM=#S).Yd71(DCffW4GY_>)DCN_#?Ha8IBJG
e:a3;-f-MRJ7\;U)BR<-K#a2>8gK5ETKKWQ)A#768#dA505BX^GC0.[\]aBUg1?[
@I1PU>71Q9QHaDFcCG&aAMB20HLU+3>^g:&DVRc4)_3B?AadL#]23O?63d=P\.TX
]X@Kf?^@(gGe8VcEK0E4ec.:B^V@fFZ)4ecQ93ZP&eHd^f9]3XQJH5Lfeaa(R\(X
5YMbO]077)J-d@X,T1]I3D.GBCJP69J0&3#3@U,KN&,K1/85^f_b-+1.dE&8045N
_Ig:H6LNXS8SMaIHD;9/LGZ7I;U&D6aA3Z.,I#VJ1^R9FTSf5e#IfSI;S8\Tf^MY
=ICD-;&\RV0gg[4<3MI)(WReXIEXV2S5P3X:\H8T:K8dI7(V5EH1-SG<#EDM.0LT
Y6S+#02P,W1BRX#EH[6=.?ME74OPXFVb^=WY@D_<__#M65g5/_5_Q(Be<&bN.XBM
(?UR4c]gZ/9\=?=f<;\-6@QJd^WLX^BR]2ZR:A9R#ceTV2K#7.3GH1>X40fX\\D<
f;.U;<CWGE23I-D,c?>PfPVaZ6PGS;/3C.MK&fV&-g7>7D5BYHB6W)-X-AK_M+Jg
U@[V,#<d/U=YIT86:#U6NCFgc5b+15c@I=Yg,C-]L;<AMNHJM7JB@f3#80SbO/f/
.N8D<[Z2@e].V&PQ_-P>#0,?7F3edfJJR7,/C\CKA76Y/=QD)e=GT#IE<>-1aVCg
;=e8Mdc\ENg)L5+Q[YWC9e&LV5+:7S=Q,/J@TE[IC(3PI)+#<?5I34gTKO.:NI]a
POHS\[C,,9NOFd&-a95O@:=#5CU<HRHEV^+fUg_[:H>2?WSU?g]3f?Y/G@&W8g4+
B?/f\WB/]RLSHAKV&&K?fFHMRWET[1QZG+<\\HY\-/FFU7/8a1F]_GQ^K=ZI>fDS
[b-RCL+GZ]AdMcC2O9O6_R9T#&VW>:DAL6+BBDKPU&2?Df3g6?JLP&)O36R,)bL_
PKDC7IAPD44VCIc(dSQ7aY[);f_KQ]XeUT3Oa/,+\2(4TF?V-(=+0P[C+2W5c-<Y
-R)A9/I2gH((72PK>(0B3UXV<VZH@QFJ+c@80#bDV26J,A;Y1:4Q7ZSOIZTg6N_E
Y6(/H^6BI^XaDdQ)g/7TNP;59OFR<RfHc-+,LDd[OdJGX\#c0K:@<:<:OE>TBE,M
[b&6-^;fVGgV(W5dS>5F+U=PPNY2ORUc:OX1QMUJSb.aX=b01GNVZK34ZTcE:0Y_
6a7#bFRgc,D=K6D(.cN1W=MAVABb;HD.134)RI[=d:#[#L,(K1QfTD+SKI3>44B3
g03c6^W&_3<e#1,=FEM_H\=,fAM/IcR/4RD[3T3\MXC_XJU7f2#ag1=&CG9T-X,T
^L#-WX,YW,//S#<1JH3Y1O(MeVaY-eg/AWQJ9B?@E-T.dHEc?#_AdgIPW&O&2>-O
5JZ[Rb:f#H^R-)<@+&2/^7JBL[fS.Ua7117T<_+#5&Qd?&45=(2/(7T[;\DI0=;O
cY?S>5N4YIARX&<7CJAJ?0T?9cJT\X8D0b@5DU</_G/fJO+c>LOaY-Q8_fU,cOOA
fU?I^_0?WNKJf(,L#_S^&JHKSC9T7BUDXBXID5Y++&bb;34_VfMRg3A:Nf@0L\+L
S]d7(=S[=+Z8K^5XK-9FeD-76?2TGHeS)E.#]<g&DHVa?^#P-X@_E39=5\XMWF^C
L+XeR33;f#;3:BdI0ZbgaV3YZA?GVW:]#d=;Z2Q+8?+)_dW\GU#QI=^Z3(A[&YKK
aZPeKF(F8A[FT-d_6Q\(J\OPXQ0;(XTcdG\I92S<H<cYQWePUc-/(1L&L)^L+c0<
+#G,JV-,3B[^;UWM>7I6Ub8J306;[<Q@4G7(^,gBXb@31=U:DBBaY,J/>]HY\6X+
5VOfB[JNDGFY(=Td#WeIA&-LeeR(e7gP.&P&_0&RNQH#HW8FG5?C+L?>GXZHO;H+
g)8@U-f@F84E?2N-PV1e4_BKDQ@:V[0I88L(_):5IB:9cC4M?24R>#2Xf/(&./M+
8\>9<0Obe2()P3g>NcGH/U5E(;^I\dSfD)bbb8LPB9BeSE)dc/-TZ/3+;YVC#@?V
11Q0KeUce/<O.&g-d+@bKO+9W?d8bd2?@\4ab]cbIXV[_\P1GM23#8;deQV>a\Id
^-)6GIG3+aMG>ZbR)OUR;(S&Y8b)<SG\Z-JfD.K1bG4=T1>)_JC9gX]=74.^Q0OW
d@RF(6VM(L>cV>e&[8[aQXM>L,\G:H4d\UJQR_a&fXE&>E?[3=VDgLZ-47X.Za/a
?FQU2NXf27H;gS[a9<@Z[O@S2KX(Ha<LVS7\S+;-cc^R#7QbeI7A9YR#A&8Y-cC(
M9_U2<)[OIV7_4_1_+[=IJRI(Kd>Q-DF[HY.&6SVV8@M:QO=g9HIWM/SSU39LHI_
c/P1Z,DM@13<MKA(6.6O3)SQ^@2B,+egM;D74gb,<R(N#V@aY=\cB94f8+;93GBS
&MS][FAQ5T)#a<:\N-b@Sg7b@=8-MA8EU;bL&JKWc8&bQ?+CP+F0gQ#AcPgO2bb0
+[R.aHb]U@)K1GY#AO,CEH3WcaU&5&@cCb<AW)LH&+8YLJI@(g:QC[T:4?P7DYI4
+(dVLH1QQD]Z0Eg;\KBLR\0TZM0gU:c>cdDV_e7F,V\ZN2DT.?R&>W6K:H#-SeUF
3J3>Z[.f]XZ4c.PEU5aQ(G2/C<C7,db@)ef(&d.T9H;4-0g\]:d0);?EZH27K/TC
]d]7V__]e.\L.4D?Sg<T1&R?758&W;0LaOZ&^127YK1WS7[g]\0e4b9^A3K)GJQb
6HMK1>.g<[CP+Gf^Bdg4Ie2E>EMAG(7JZ8M^^,2ITD(?f<1;_D=gK9(I8SELPUR\
=7K>YU6\8EFNK#<5)NWU,KH;9Y1+DK66J8@&MV,;/g^f?=dE8-YC]P\-3cWg+J&U
>VD8XN:F+5XU-U66KYbUEKKc].=#9=WTHc;LX94R6YY#WUGM8^_BIC#GLdK#X?@G
O+T.IRU+:>GKUEC@0EV6b.gfG(WLBG/-[AFASSPJ(@<>K18/8]P<g5eB5[E=YHY[
TFDKR)^8<FCG,aNf)MI7,dCW>Ad:GK[ebeIbG=7Q=]J66BH[\,P#4>-HR19R=TBV
M=@POb;(=]/AO=/P=Ad7\\e(4.CaFd9MX7;0gJIF=2dW;DL?=RAO8>:SK,1/1CQB
:3/NUDeFI)CN6G1D@57B6]+Uc5#93Z02XWN>:Q5a4ZIER]\XI[Fa_<M/V[:8(CNc
@,G7a3GC4dDB7>f^;/JT]1LB?WDOQI\2HJLg2M1/PU/AdUGA>aH+WD)/-310c7U+
_F>34F@1N(/gO1B2?@AW:;M5aY2:_?Xffc0]NBcC^Q8aD(GZJ[LI&W]&VJ&D.\a5
=YSZIYTI=356P]W-g>/K9\SOBW<F/UfBgL_RRb7TU,FZM2e16;\1WI336D,?+FK&
A<V+-(U2:+5/U=#GD=aD#0<a83(&+Qeae;eV-EN,>I0/CR29CJ2K4NW@37EYK0.7
;\8S5dNeMBU&(]15a6]Q?2X.]/<gW)B#WQM.CIP44>[:IT<F/@:0T53LCL<+2;GC
6EN5C&RN<3M[?\AQcc19\^6/AOKgIM\c3FOP>cQfFNS#cQ@-]503A7DD^\9S.A>L
E0eKYWAN/(.\D-QELS=\FK8AMDg:DQ=4RAPKN6;I#&d&E[@(Tdf)TJ]3>8X42Uc/
I54&S-a-1\)HA^>5:Hb&O#M-+,(Q+3=^(-;Wa5UBFMJ)\UYFd)5.g][fDJ<KV/J+
91b76g,TUWO,<0[8=K,3<d@ZL#B<\E&,/(BVX9P9OTH=bT5\TedeeDPT]P.bc3c.
MI_]8&<M0\C]^5?=\a;GA.XMIa5C+==IdS(GW61?0EcOIOFVU_=&g=d-QGQL9F1<
KePT84,(.B9H:?33;+LZF,.C1YROa3K\\L7](ggNE.<f24>,-c/SE(TS;U+OD/(Z
_R5Za/<&a>?eCHA)?AS6U4.]_\1.X[W(/S]#=T.1B0L89G7S]EE6UCd-f_?bZfCB
e@Z-XC>bDUGe>)Y9cN75F>=b0YB@<3>7,ZQ1YV@IEBCD/LZLT&=RJ\c5=PK:b+@O
g(I^LJUB?BJbM?QKYK^Re>0R;W-;NU9>M/-FTLY:A_HE&F?e-9a\_\[;&,A.;c,0
1_0e/XTW<5GTG?HOOA3_K?<JaQgEZ=.ZA?N:OgB?=.UfK(I2e+[T5:IM5cHV5X;^
LS]\+?]5ee;DP26VALMVAQbU.8;2QRMHED4[15#aa;<N05)#5cT&OT6PA&IQ]?e1
9Ve_C#UIa(gC?,<d18Va4#<dfJ.<DDfGEIT3/(N4D?V1G2JWHB40X7VMG\YeB,SD
0<ccYO]R<a&X@\^95I+)D1g&IK<KUHFKWb.KXSHFWJ&/_cH5ED;LJB?CSe,V]EFK
/>S5?6eQTS=S4H01@[P&PG.)PQ:8,E9:L>ONQGbbV.?BOZ]dg)U&G>RUR2/3_8RT
SW\b6?g(2a]aU^,He(]T++S38C8V#LVe4#<5Y[W4<P2&<>38e>865Db4YW1Vg7e_
VM(&JT8)&?+AaP46]4GD-1H8109e2NVfP?S0C@S;[8X[dQL5RN:adN_WQJ;5]DEF
VF]^C+>0)\2Q>bKaNB=S@)#[/RUC]bWGB6:VS^da&_>&1@dS>]b9X^9QfU_=35g(
RD9eUSZGd5[MK3P(agW8(DdLQD7G)JaMe?7LE(>RPLB3R74ES,A=H30M##_-CI;H
J1E&10Za+XU,Hb;HZJG(9]0+(NOfM>-5OU][E&,(=&(HD:+X<2\?CYGP&)ZEGJ8g
113355E6LLYQM>C&H<K<d8=/f2S^d1gNcLT3\gTB=?+W9Q;]#^fU[+D+a3gX8=3;
86.cW#M3Dee]Y8.8KC?WJ2bHd2>#bG<MMc6]HEK_P92N>AJKfVRVH:^,[XF+f_da
/0@E]C4]ZWPKb8TRNdB18T?b-\MJ4CJ.?)=0C\\fS+29a;KJE:<I7CdJ.@WME=fR
PfX?-Y4^I3eY,a[>_Tg80H(GYCQH-g)b..;?(:7+K,@KJcT_@^@,OSY-B1PSR\1\
bIZa4L6aG8gZVGOfdg9DR2F<F[@7&U1=g(b6I<f48O?@HB##;VVR0</N[1KUON&X
JJVEf3UeR#X>@4IcM.EY?HM^Yg387S48(7\^/4NNYf5c0#;PMEA^df2J1,PM[]B)
D\b/UFFaVAGKDS;7f15?YJ#M0<WYgZUK3E>16fS#;F;810&[)0^]^P^,K8WP&.dX
6XAG4V20#=Q,&9Iba<L_0SB9V(^T:=9UEFD7\T@ReCc.+:E3H;SRLIaL3[2&]CB_
3M#B=?:JRXW1a3&(GQe\cHd_=d(RP1W>)25WJ<H&C1>2=@1Y2#C9+5L^FaRJN#/5
^B:[3751P-:<d>8_.18;TU^JD:C>5>RBFGX>;H9WIR77<CY-M<WV[#C)D:#fX_=S
.g8\:5?1.OAK9\?KVES@CGLX@Y]N_?-X^a=FP;ILTI>>0^7I36CC)8\G-1]PSLT8
XO_bfB]/JfA4)7bdJ&07C@DFbVdSI>-LAcXE:_>ZFMA)cW8,L:a:TG>X/#;(U\4O
B>bQG,RE_T)M[&f--)\X16T_/2MOR-+<>da8Nbe-V)W&cT8K9+79TR?/d,/?7)KQ
dM[3V_0_,52CCbE@[NPFVI5a7B\F2><LM8Cc-^F:VX7eg+Ogf19VIC?-H+da6@B\
Wda_>+ef&ae::8B:;HU])cA,Z:A+FZ<HV^L=6eT[9J1\M3S.c.]f((M&C3R=;](d
RZ&3-G3X1g);AT9^Dc6H^L?MOKDe^W:gD[JCKD3(/#&?7a8MSg1+GfQ7g5[M=64N
^g6#;b-<3DJ2R7UMW9[?L-4b3OJ#.5^X1&a17Y[V;ceYP4a_J(+K1GX3Z]WWdOE,
cMJ8/,3&c7c6#:0TJOOSgYd[eL>ZU;Ib5.eg/T]cQ6:JF.Z_9AB0\LPdfE-__Y#+
J4Y9-[+X+J(0>,E2c/N;H<06\f\R9-dM#-a#f1IHQ(5QGEJFe-cCe+#THNC40A;_
aHe/X1MNWCMOWA3]PRL8.9WU5RH.<GZEd=(GY2a[BB0Z#@NRNR6.=B??KQ2=]PDQ
.@P:+f)_DU,SUD&NK+&:fe.b-6EJRB/a3PL@GG#[?f:?Y2-^UIgQAU(1Od>f)b=a
:+]I<B<d7LQ5,,c-L&=RE6F5UC(U2]^8B(5T8T]8<c>TYP060<\gV;0PL#b0ILEQ
Oe5a<1.HX^4La/+)JX9A0;3MU2QG2?;3R/[+K74772.N(e/NTX^JaG(P]g/1?F:D
0.8DFRdeSc.g[3@H:,>C1P9b5P2,E9P:@BFgV\I,09Te_?<X;Ng;?X6W=Q1f&X/9
Ld37_M5HACRTZbX<5PGQ/.@Ng+Y9fF1;,O:#C-@<PPA[#])\R=A@N3Y;07VX[Y&V
6U8271@:bfbIJ_NPa:=KV0I^DNO23P@cW\aKP230NVL6R\W:_(+a6d)Y+O,T\@R#
c#2M6C4Y+_]HQ<ORL=_<14BF\+dK>3&EB=CCF;S5HJ:G:1CO98edFc>X:C]YUP)@
@FdQFI>&LA?NU5HEV:^1[S@ATg7&dA(^HSEKH_H32b2_Ic<PHHgg#1J[[bf[6\8I
=M9B#ER.>@L)g@L,ZOT;LNeR[<V=WWB^D]+c<gZ?67HTa5,<6>#:<R\+f_]#06<b
,=Sg0IN<ZO+c69OdX_8K,/bA=AIW-4e[+;,[15FRd8J\(9_XX<LZ?>L&]BRBWL6b
@;X7(<+U>f<L^)[Nbd0A[eT\a\87J7KH8DU/709+VK^BJOG;],]PK3W3b<-5/(H_
X_K6.KD/JIf,@M</D;_D>7f66O/B\@AN?#SX_HC<KXV4G4>887gf.>2V4N0,HC#2
f,(&^+E(Uf.[Z+SFP\UVNg&X\3cbO>D_OHSC,^97?A<A7bBd/V=UCLK=>WbY@84]
8FT;SSY8UNB>(SA4Iea=M6Bf,I(46L.M4]3I?\.EYWFQS#_/IY5_BDgX_PEgaBe@
e\?Q>T9B^5)H,UDEaK@+F-&3XF)9Ldbad(Yd>UFAZM:c]Saf37B-\MG;:L#;eSH&
8[5X6a+E/ZGLBUG]=<Ad,PF0=\P0L6,WD2,DT2f?KIN]=\^8Ja8d_L3-93f7eRF@
RR1PeAA[?R9;]..NL.N:9,U]1TM?C-W6[b,@1\[XbHAPP\J@GR>>?3g.4K0S7U#a
MT&_G5Q51S8QNI7#E.<#-\NB-FF8aH5ZKLZN7FR.,(4\4M,g55-O(FFRM6T&fF;L
]:QbDEbHOIW>=KA+?V2,9gM)=K_I1F=N7SMMML2G^M[Fd,(g<K(@[1#13>f9b+.R
H@5dY<gY1?-XE#VB[M56D([19M:/A?cY,aR/2.EXG&]LN1C3O4Mg,dT7]]1fKG0)
:H)a+,XR9HLF0W,LZ^:+CKR6^>/?:WeVDYM[ZR3B<#gPYc>#&WR,Y>TU3D/94UH1
;=1<0CGB(V9GYYcK-X#2Z:/fL-e1Y6UOIV6Z^E.2O+e3bbI(A7YB1VDBbSM7EAXL
8V3F>Sg-R350^_1>Z/,(dKf;1O,L@G/V67JD_\BQ)3MRHDdaHLFD/5b92X]:.BH6
6GYcVX4L?S.00>?0THVP2Z?&5H@5:JM]@bS(=Qd?T1R3A9BCf,Q7G=^&:/MIH,4B
gg/bZEdDS,1^_@5A1&\a3aZ3962;JP@COFJF\FH5aY<,EHM.#ZW@:I5,R1(b;6I)
C-:.3VU]EN_3-W<<28LZ?8;)Q.(bg=A5a/Z5=cAKdeS:6bM,=+-dQ<8UbL\aAQS0
8&]G8BbL6UQ4H?8[#_703]3@Kc\[^2287>4RYb93+X[6C4=K@CVE]B47MFAa4Gbf
Db8>\X8:&,VXTPBG32]2M);?6-1Ne/A3QMQEGLMK^JPa4/\F2P1EHQ\?7>[43W8&
D,dScE9BL@T/Z8fE25_=b0J]:fEP+7X;I2EN-2?9:FJ_P5,;;:K(NCYTFA2(Y)NV
[#K<3\(cIQ9995T#2OI,2]H[]TOaG&G]b[A:X(g._c4GDJ)RQ&YQ7Y)W3EaPCWUQ
WNJ7gCX+SGK?QP(30_T)96U2\K;-<T\7<9^6M4GWF#,LV5eP7;;N2L@#4^_<]GC.
<2O-1Y#UM5c7>704YUGgMT)QD5+Q5#^(S]+G8MQd2^g@^]<#GS^WIK=8d)-&5D?B
M>e0S-B0[0,_T=QW5d,GV.B,0LBS_N7QFJ4+J5-LQJZZ3YU]f]^\c^BV31W]E;]O
PeJM;O6BU.EX7;[4d0dfXX3J<2M>0+24>\cO[O_3F#.cJ\[0&<cN+6.1eg1>a72f
IMIBR4gQGS#C8#_60?Re?VYT4?F-T[-P::Qa2c:L8PFCZcF@</aLbW08Y.^JTQgW
E8L[fH14_cV4=B#d<6GNaHQMJIXDR3TJ>)B4&T(JLb#JB#:_)HZ^=8TV)-b\K>7W
_bF[_.9H9_4S,=L]3GZ&TCK&.9fIgQRE@,YED4W]#USa:MQ[MYcVRIf8;DH@4MG5
9AX:aZZ5E3;0>K=#]4Mc+AFVWKJPF8\0-M#[?45H:C;8:Oc8DH/AQ#[bD33T\9d=
R<Gg/<OP5^&[DY<XX(67I78?:FBTK0H1=g^;#eR<Q9EN6AW_:2I^\K@C@^A:VKU/
,X=QSKZ94eWf</DK7X79e5^4T=K.92G\Ac.;IC-2=9QM;H>3#WO6d<@J;J=(1SIf
<6FKb??^U;.eWVH(,eaBNSR<]Udd4N/SK-0^3]SH@@)PK4VabJ(17YM33<9[G1cR
VeOHS80DWJZObW:<A(L))<YJPL-R6ESMGENN.?c8_g[Ef04gJLf>8<^[gU5V60;g
47BJZ][?<GC:FBFPGP=-=)gQVB;e&d3f\MeW+e\_PA7?0>O/_.;\#@ZD@<6L^OCI
DD;7JR<OFIX]N#DUH1J4[D8>W?;@O=,HLRESU7D=>^NWbNC4^V&UTE^_JPMSdN8@
1ULN@/T-3ZNFE[]5)@b5G3(SU.deUK)XECB=CIR7S(A46.c4gc,-@4>#MYCH..^a
X>,A/B@SKb_GH4C\M--K0\MKKOdLD)9]]&\X_(#CXUY;0)<U^9eBB?E(dG&_S&1b
F61YZf)HPb(+\,Y5f-5R(8F>.5SF&;M4L;J^,e]0#Z^:)ER7,,J5f<7G3N)\(RZV
4KS[@g3FPAFZJ+eNAEZK?+I2Z7Ac=aW7FgV:2-2X]4[Q,[]E/HF]:e,Y[C@3gaP:
C8;E&OR?C>W\UbNF0WFA=/SDPMN:(+77=?L\L-X+E>HY1e>0RHf6S&0.f:X\0dAE
/Zb+D]4Q?bLOZO4LM]R,4]L9IC1#E?e>FP68DD@^a@c\<0aX.W5g>(EUF_([Yde.
<STYG_@^-&BYP,\:g4.(.]f,b_P4WMCF7;[WWg4R]f)3A4;NfZ@1&UPdbHOg]9RO
P9/8F<Y\4M=dZUc=eM?dcJ&HgOdeMO=8A+1#8R3b9V,1=[X;@a.(d=8Hg.(N[fDD
?^B]J(K?LO#HRagOKC>ZXgL1eM-2&K@Z#fa:V(fIAH[):,4<,SAaIC_S);(7R@I@
R1U_ad>B?a4Xc7Y6?V6_[O<RV(Bg+#WW5-9D[gGY(d1eH7R5]U:fJ0>9K;_I2KA?
/[J>PET38(Q,f7ESL\@aII3KHEXSU+Q;;K7@Z83UZ:P]@)T9.G4eQ&:^&dfSLF>e
[)2&>X_.D)Z.^Q_d,/MBR#09>K8fKEP#d0eKJ_HKeXMZHcR-AML6>XHD2J]O\XdT
TOQF.R4=^fF3#7JT_<G2=_g]?P,=dV#WMS8?;B8_T2[3W\<eWGZaOWI1:/<dRF8C
[ZG)6ZJT\WVb7VV]..Q0b0G0Yd4=Q46+Ub_4RX08:eKB\X5gb=ZDQ_KP9=VM:<Ba
MV0=Q<L-P_5)]#IWSKEK#/+V8Mc1/8Q5QGJION5:J,6<F/MI==N5(1;#R>>L(Q))
K6&O3W_BM48AcX6NIZ=U(&aCFR@<O:M.=S847FK+Gg2Y^8[IF]IR-BL[@==&Uge7
eT&>a4b1I3D7;T0VSK.?ge..AQ&RPJQ0[HaF)f9MD(B[419VQB)G8B?V&4,Af^KA
D=KX2P0OgN<)A/D?eN1YD]5e)<])YGd5NFI#JOW<]P^[5HT@b#G2]0>&C6-90_A5
YGLFH9^_<@bGZ\TBM_VXgVH534YVf^+6G&CR2UNE(O?1BFNdA2TU(X_2RRE#LR.=
7FE,)&e26bgUgV,:4+3BG2Nf#-EY^0VF+:U3:]E,YEU7;gB6]cX0]?[RBO#C?_Ab
V8);WZ@X0T=D@E#a/23+8X#I5g1d[IEP6e^,E:Z/QM=d<dgKG9KdfA@E2)/8.F+I
[QDf8/F3Ja]XQ05E&Hd[C(D>53(#R#F5;F18Y[U2;f-&&WY486dS6L3dMAGHc\J2
<fJ#]VbWa;_ad<[&CMO9VbDJdYQY_Q03B/M(aH\6TMQ>3;E#9Y-b+))2FH\VV;HW
G)WaH71W:N-W3efZW(7JCU-C,Dfb=JAdZB4SJ&9@20K5AA^?T]e\@VQ5GJS6c9Ne
FN8&K=7_QfWKI(D5e2]TI>D?+DK^&dH30F?<C;K#;O/=6\_:P6fFb#])@\19^3b@
CY;BE>O;KM:;dV3+QKZXb51f;V2ZNDAXNS<.+9_g0g4IVcPS4;AF@;_+?2V3#QG/
[:ggb[MIEVCCM/E071Aa6V(P]/eVg,2]@c8(RG[@XTeU47Mg3GOYY_(&ZZB75KP8
V)NRVc0E]8M\b=D6dbWXTH+\+&P,-#T]J;?0eEC-\H3O#UI9e-82dd.MONGH]R>D
4Y9)dHK==7/=>FFD)PIa[9MW=]D80?1_a&gOVJ3F[.LU(+71VEJ^;MQHSe<b)CaU
R,DcFRe2[:U^H[UT48J(4eHNP(#S<aEP+/O-I(c)Q1XXNA,MV51HD/G/_^eV(E1e
ANg5KI1-D.K+50UPXUg2aV9?BY2H()\B969e#Mg<]+_@JL>#-e:M-GT6+6RaE@Zg
>24?:Q&D-UXYY7OIA<AH>]DIZeLb@8>TX\e^@WNd6N7@F<6ZfSKVD</]FM_C75Jf
I.)Wd>31&I:dW&TNC9/>QGXIS/+fOR+-N1;PU/J1K]]6SY9,_16f@>fP_&)QHIGY
cK58:4^@EBQ]<\UGX#94a,FZV@;VY9,&\>V?4J^R)U@Rbc-T&=_:HB=>.g>J&Bg1
gB7FZR24//\2_]?T\&)QbUeS;DF1?Z-.P4E6)^:?W,_:ZQ2_MZ]CQSYXE[5Sf2a1
[C0SF[Z_W=I=&eGX>;cg@82KXYDBe4LYad-RAM/aT]JS.F?2HDJ6VWB-<_N6)=BC
1VbHNPO7#b[a_O0XC_[YLgUG]cdDYC-0\83&R@02E#O2<H@&CC9YObK#S\^cUW23
:@LJ.cZc/0/.ZGX13CEFWN]C-F[b\IY/8JLgIaK.5T?0DP(VI/-UC<e?PWM>^eGe
E+g?K-3&L\B9]Tb_<7FUJ7D,[JC4@(96V9:77/f)&\WWb9ZU]?d3fJ3[d79^4Q&]
MQ9))9EA<]PPNbR-7F;W\AYHH8\+09Y1^0+91R5Zg26=D3cJQ&XEA+:fN(a\7BD/
f.7+5YGBgHN3e_6NeGIIXB)G\(H?^5N2IRYP>-^D(c02#(5ZWf]YL8Z]]C@2]Z,a
:SAdX>LE5ST&E)d9+N[2RW^.NH>H9d6U\=<HB:@gCc3\E-+Ea0g85Uf4O_/E+RWM
+1_0/E/039cIE&,.C1HD0,F^T26aeI1=d<[HHTOK(;)ZW-#DE:EOMR[?><..2#F@
.4>Wa4:2-_8e:,5Qa#Q?GDYJ@9;#WO&;7E1:@5Td4@8NOBZf>^0=5-O7eI510EWR
(\f7)LE?8_=[:3LM)9W;TE?E2);+AHB4>-_B;1CMX=U.E:-+CUK<4G:2[C4.PNRP
fVJDAYb@:-?WREA0@;Y=:2B[^_&;AY4.+ReAI?Td3/1:fG#UKC5R1E@e3GbH,0Z>
JRXI]Oc^YY6d(/+(FC&#Z6B.UbRD8AfJegG,b]5W_&d]L:4+bP_97^?C_B^C3ER9
Cg9.dLHV:],D(T5@_dAGIcSb&DT_1AcV58^#(S^??6BY3P./,(bO69BfUfKe>L&K
]CZJP&E]K:>GGMgT0@3:CM=T@:/#PV.Q3;0b\\<+6_UgHL2IZH9#/Z;I6W5b#.20
3/[eGY:@8RBI4=2TW,+N.](W4T[.#LW_FO<<;ZV=B)_\NZ&V]C_aY6b]]N?,A7Q]
Z7_&>E9ZK:LKdc8DIO9_S>PBeeb;Lg=CSW-R]]2[[bYQ3_#QG,eLANU;I&(GLE33
U9&:7-QaYY9^d+gc(+GRUN?U<.4IfYY3]fF@@?>G4O>2\_U3T+F(LL(HGH(0Rd7Y
Ca)RFa0GfF79#f4d)5H(.-CDa3W+,;/#^<;@E<VTI;^+/WCAI<^#BYQ6^8U3;\I[
]:<DgQ0?QRW.K9SUVE3?IU1YD(BQK=U[687cWT]1eVcBXbgcOGfP>A?L4YV;cc-W
2^/++<PJ[0GC-B^F^_]G-fa2W[_:=@HUP3N<(E_C.+dLR3eG<0NK2WO;eH;e]#ce
F-d</33LFZ(]8.46aQOS_5Q(8&RgO3gKgV&C9f]4_d/VAHJ,Z(24R2PE1f[Z+<D5
-T\MWS2XN9Te6EV2_JN9Q>.\0;2F@aM=QY[gAX_K)D)::P@]J/.dU&gM5Ab4]+FF
?1/gYOeB0<.V+]:1JIUX?M0&(fLG/S.H5XS1a5fUb7LH[?GNf^g=9TM>5[F,YAgZ
7Og#?Y7P/F3NHH(gcFGAI\E#V+0R)b2=/EK>I)WTgM&0=2>R&5@\e#NC85N8.Z=G
:g[B^7?.dfYXfE/I_)?\W]fE<BG3:XM:Yf_N:-@fVY>35gTE+NKVJg,4FNCW,3FX
g/Ya&1,N+:OOQSaQ4?^Ka(CERdC9_bYa/(Wb&d(Q@P\&0VM.,U&:C4K(4ZKZba4O
+H+W=:I=1gE?Y&CGab#C+--^YSYbKYf07G\eXPXO<(G#Xb5_T\?8I74&5_B;3E3.
&HbE)+W=D-<[c50T&NOXO>,:/7NL2T^0,]&Y9CUcb6#^_]FU+aS6,[b^A:;55J,f
F04Y-;d]\1S]Sb5FFD6ZL&#GTb+K3/fBZW71f[LA(Ed(;?8f0gQ4WC90EBU1H#c)
?G(--UI<_PLJ7dbBG;EDDIc);eQ<gB>.U=7/Af1ae@Sa>;.(1M2b7S:dEK4^VdgO
fZ15S?b_RN;4Fbe\fa8)&3&JM@Z@;W?&H<;C4^aC)Ug->DX3P.O=:O4Ka)>_OK:K
,e-)NL[J=+gM<#W5D&Cc2e__;2).7Vf6O6PUZW,RD@X+a#Y6g-XT+0gGO0.ZR,J)
1EObN#:G43(Q5ZfcP\^7GW8YEedf)QU&@IdaH;H01^V#G,#2EQ]&1.ZIPUE<B7ce
d5).PZL:O=VZM+NaQO47a4HeH.K#MODGO?YB;XL]^(?fg9RM3,[@@,SFGX-Wd8\V
M3T>b7bKg?[2U1^a_:@(_a,cBQKKDAY08;b\gfa>U2BOS6UC1RJaI<bK?)a,;]Ye
SYaaAP).=#Q[P<W9H3)=]XaTHN4C)RgUbP^-.bN3;e-/(d=99.>[S&.-E4.W<+&K
Re?TaNF_&MAce7942cMTPc[g#1]+W[RE@]_43^0IJcUSC2^-PV#_37W2IB),fD8K
@<=#J;8(d+?YJLZd9eV.OeTJgcKc8LCf=2Q=BNB#@F-1G5=<@6==4+3Z&C[W+5OO
PW?BMa:eP+A(ZV8M.0=8:C(Vbd<I-/d@MDV>7K6=)1<&1=C+@93@;Pg0gHQ5B=Zb
_W&bC8T<P+OYe&(@E)GJ?8^g_@P4.I:(.48^<[6PD>4+:E^LG_)MX>2YH;\[P>J>
3E@QL.g3P#UJ]:KTB,Gc93]55>UVC[D3EI1&=GEJUP=\(XC1R4W(A&E@Z@2?\=Hd
I9VVeI&Y^9@N\OP+>bLc8CQ?_Bg)dH5\dL@TX(C@,bSD7@YT>;C-a:9]6f<BW(=g
5PY>\]O].N1@BJd:XJ.W;;YDG-5>W>?10c\;KRe2]VfUD29:a2\-8Y_dc3abH/?U
S6=9Q6E[4=/H[fC7.+1NLC8K#IX1B0\TP6ZM)T+;[K?TC5d[O+)D?IR@Y5b<I_9P
B?OHJ08Ce/,-4/]<:W60b-?H-5[2DBGL/SO+)_9c0=WZe?#S64Wg-L#edZ?&(G=\
#R18UJJ>([QCVW+IMV5=Ff;UF+HFTR?X>]6984MV.1P/6C[&,KeaEB77TSf.X@4Q
eW-2DM8RM.8a#dda#4#^?5&^Y^/e8WZD[R_]gOCcOJfI]Z\5.[PaIY.#f4WP@f-]
Z59D@M#SXUZA^/#ddc)K;O0&CTA;Q._-V4XP5+3?+=)RLXRS6KJ;=_Q>H5#<4a4F
MdXY3Z-KUJ/U8)f9<b)?XHTg:_F:_^B?]LgQA_4^-8SA3d54.PHTA8)CdSH#2AgY
06ODg90g1LI1GMBQ5AI>MVQA_dD1MMI/#Pc9GMUA_-R5<d8[:U<RXOb;00E.&5c7
#E@K;=4X5VLO6&KF)^-B@Y,eb7^CUU\g,LWW?M#:RMY3D_^]O-W@M7ZgFRVUN-/P
MHQRX8FQV>eMB?V/6:b4EU;g=3TNg&QS0,.G_W-AL4H5YDaYX6T@,8+69/UB?\cL
J(X-<<0E/HO^Q\A/2cf0(JGM.NB,(cLB^2:58EPd1CD^LS0\(eD</99&TD.aZdf5
(.c1WF.>]QH5N-86/LJIc2&RT?9IV?5WJ6BOSX2,MYWS<3#A6@7D&c3-SgbKL(7.
[6\.C(J,S:JD)4gd2HcRZ[\)#,N@/&d_VM/9?2f80:4,_\[54ebd4<_<<93^<TI6
9U][#?F#&dNLd,b)@G5REV/\bD4#g[>CA>YYY&bJ(ge4GY9\+#0eF_.Q\ZLMZSPa
-g>.NKQ8aI3;?.^=5CR/J:[Y;<bKTORfPF4BdV2-7#@JfES3X6C&OM+;\[SH4_g,
<M)#6g:.IXJTK6]5UM-R[FY(-K?OFg/?B767/Ub)Wf[cA:;Z7JXWPQUSRD8:W4fR
=R@3a&<0OXgAg^XfJ5cdd&00Y\bRJ_FK\[Je\f,-LOHgeU,(A>4<3b8d>:aFW6O&
,ZaU5f\@X99Le>Q2T(5<C<f)\+I4_O^5VJXGfM5;(+UbA6_05^S@.HK8g(aTI.cM
[,KW>.YS::d@^EI0UCYX&G]JKX&_WfLH.gT5#EYT>dg]dRR]E\3U,J.N1\@5Bc>V
dDbVAB4V.gde6ND8_MZ3)W?G?)bV5]HILQ6D;b,)DY72]\MDX-I_:V#BdEf4>FI@
E6IU.3&N]aV3RG0FW5OOZH0+M/+H16E>V^9YUB1^I:Ke)M1CFPNO#?93&64\Pa4,
(EJ?0J)13CY4\TNc#H_dG@X\<&egKcJ,D&XEPJfHQYGK@3B8=Se4+)&O)N@??DF9
AaPH=?:XT?[OED39^?&gb@E)+N1+8]=8;PLL/X#F]6FL;7aZDB_Nd5^QMHU0\L+b
KQ]R@KB=^STb9]1;:9I;_DOe,<5Efc6QgAVgU9Z#d+1(f+F].11&WE_9,\@WE(_U
&SN1R<\^U2T4UOZ#H(8ER/-e\f5e(,:ce5W+;Ae8Y-[:A6.FSD7C/F0\7Qe]Ha\]
Z&g#F=eWF#->R=-b.O43\O\Q/].3&L>R&P_N6=b&1RT8b\).bN1]0G=.;3HYJZ(]
-+&:eN-ZU(e3TeSdVA-QP09Yd8NN3W5gQ7-/SV94]V:]FKOg7B;TAKV61#g)f;^G
LE;07dV<cIe)8=K8EPe09Z+9:7[D(,]cY]?T5=-(Y0be_eR9f.>_N3>adX+G1?0R
f>2f.7O3R]H#/,4=QVWH,:;Z#E9522@^79MBMM9e-717O+/Qa7)8;QC.gLW?Tb(:
b?#:U26=\#X4_B6I2?(Oe#=<YR-C=;IQ_R_[=9:L8?O]UNWXaR9O2U_,0K3/c2:4
-7>;>Le?@7#86_\H&=/4O\ef[O&,=RV<T,RdOTa-Zd9Kc\a=1QKK?_Z<UAY<ZPH9
ML(d>Q;1DXcbX/3=Pa,U\fK/J1&5?OedMVf+J.a?B5/=^eYAV^[]/QSB2Tf(:ZbP
+<D>4K3T\Z)f7/2__1Z7#=^X//>+K9JI:e)UXR-F=bZ]+6]dgC3fGaK8bL&Q3Q#c
b_)AYCEC/eZ2bRGWL@BWRL=/+K=-T;g_O;9(/(PaIGYG-]F2:TfJSbWRRJgW/eLd
E)f^&OfFKcZ[-T/;T2c&e]RZA2@:.MS#[]M#(O)>C\\7_aXf3-U8a]?1ULL+N)9&
Q7?Xe[O9S=g&b_3^0TBI^[G@9QWg&@+,b+D:C_->27;a;-77S6+B<G@@a8[94P?_
fdG]a,NL0,/GL#L?Y?TeV-W0C5M&M7_<P?5U04E<7CggG79@:AZ,R9R;D]Q^HZYR
H.f&UET7Ib8T?#OgHMUHAbfDBRg5A-bTJN1?D>=g-a&8WLX-0J;&[^#8/\[+I7W.
(C=OdcFd,_4/ATXXM/G0\ZfPR^?__0=8O/>Za1ZJ[R6A\S2/P+eETH[5SWcMO@U=
2MUCZ2CcL<g3dP]-48f[2U\.8D.Ub]N]abDb/U1)-+NP6,7C-@FgW>UL1\g&K7H3
K=c3?^#+<@1NW3.9YN<[^E6<MW0B<C4,+(70c__XMRHae.BSU8>W)9?D>PCLHJVU
<F7D9M_g:)B6VXXB&DQJVbfUH?N#P?GI1Sf][V3[IGgE;N_8OTF-5&7]JTe,0^SG
(]2cZOX#?+&<,A5QE8_(XgBTO?g=,N)-4aF#Wf:E5_Z4DdRN\[UULU185Yb-6-^_
?T4N0_ffBV3?d/7K&\N1,QMM\4GPU8CA6O]\L+LG353]SgUP\4\ER[?9:)E6a&OL
afWT4#Ve.E:Q[W](Kd(@V;/5(2.@+Qf9_F5VDC5B9R38P[ca\5Q(Q)>=+(N-/UZa
YM/_6WT2Q.64UcXFEC&#L35#ZGe=+9)2;Sag+EPOFGPJ\F[3AG&9R4(64b30=4#H
+W=I\Y\S2GO9f43cE8_a8R<T8c1V;6B73[8)?cUS,EE./]@3_ZfR1/BN3<F5cZ8@
c4aI,]5/N]A5Lg_:8gCIQ7.<JVQ@Y6M]IIRd3Dd6Z-A]F-RY0-O=W>ZG.<FKA#9B
^;E9^(:D0-3;f;=J^.g]adGO;(e:>GY<77:GaY4M<=g8;XIZT8=);VN/dL&,S,#\
TD<EAdS><dG-WWY-G8TIfB;_Z1b&bS9AL]2<T(^bTJS#:>_^Y83aBBVTX2\CA9ZJ
9KO0cXb>>#F)+g^Z_#,PC1K+\aIJUK?F.R?J2H:d-\W>.7H]JXSXU7@:A@aGaSSL
cB3LUZX)BQ&,ZE>aB25N+)OW+eUU[2TB;&@>+ECULNX3XH7b,]X:=5G@:;&7d7c8
I#Jc#RUbD\([3T&P)W6Y[6(-<XcIWMLX^6R42>#O2\Pg-:H\P^eecUbcZ2?,.65(
9X;GQD4>CZ=@-a@8P+_WZ]d?\[1eE;OR/V+0M+eO;FJYSI+KHH6@,T7fL1Z[\L7:
XRSVbP3>5#a^_E&6K<gFaL)PX8@66-Z#De@R?@W@RR1<)dBGK2.f=WTcIZWFRU>c
X)CBH3[g7T(#.[a4R6.<=21)\5ZP7OC-XR@MM#:.e9d)MTQL+LH3L2,7CT#fa?9Q
V.;1[D1#7,\J301C0&\cf=dL@BEZ]OYc(DN62^+&D]-2W30&?(ZJ4SE)J41e8Ua]
[JWOR7X]=963KMQaS0M8+@UYdM\Q+f>1<.-.7(:JgB:60K,Na-,@+E;-XM<Z<@H;
AG91MOCE/L7;^C/bUd8WYZ;YFbZDSS3?NXSEM-7S&d-A2LWaV,^FVcc8H]5/gf)9
HO,.4UQg:JF9-fN<XFTP+53UXR^)>_9VJB1&:)Q]3(bNb0aUGP4UeI=YcD-?P2=>
WC:NA(=_7.ffC7aA^J(g3&6?c6Ge(F+4>LcW5[B]NeHYH/I_KBXUIF7U+C&&6cg0
G2QM87D)92(;bR-<.H.Ma&18\X=NX?OP8_XG)+.3275N3YAfD1@51L57[8A.Fd?L
<VAX^\D?W4[\:;d;B)F]?++=76e(X>b3WD,g)BEfE6&03MH\4DUJR4a8V_LI^9dX
WQTfS&Jb2JV;6bWZZdYJF8DU)1+;g38?Y7]E_&Z_[cdAC-aFb4J+(&Hbb4\IOO&B
]Cd642NWUWH;;Ide85UX+2E7)dX5(JF-[.]:_),6ZVA_#Zg]S<4_>fUH44+1g8JK
P&L?LBS[g;E4AUWLX:9[L=NI4<=U\XC]^9W7Y?@?H=--Z2AbcR[5c9L4O_>=>?8R
F=&-]9CP)^Y:^HAFG_ILW?,_,T+75PR@.MaL8<O9^PN;EJ@P:]7@e=eHF=]e,,Z/
Gb@CH/02V(\Oa5^)78Oe7OX^&X]=X>6R4CSY2680f[ZE6gDCS6Jg_,/1CUC,]0b9
\DAE;=aY#AK0;B3:4EB1/:<=f^HBc5T\UUYf5g_FeT1.O:dU_TcB4M65B#ZJEKD>
4ANAJLQdbLA7Ta3Ja^[-=VYSZXCYMQGX/[:N)eC0f?)F^eZC/\D6]<;dMIL7>^#;
B#a6H^T))XY^U/A]CKDbK;F8((2<O<(U9BLEg_LC<6Ad)K9e9?,=#WWcS9+=AI(R
)(CYJQ.AYGME:SAT98[Y2]#SRE@55Rf>dXBU_34&<)b/,U#7K-.B.CI0,c&Z\3Sd
9]&FHZT:U2(4T3FDefdG+b=66TC_1@1@5Ib#Y2WC@3<;N>T\a?C22OeO6D2YcX5-
>dITZ++dB_YeEIU8:BUOI+[#]5SOfCU2UPBT)EQD-fdVR^U3V&=_:;e4]/DF2eMf
=FF2KSK@#.N#A.)E7KQ.99[,OG>aSZ9)0@V#IS(SEFI#VE7dV3-.1a?(65Y+2HF;
LYR_/3Fg]b0@e5CeO4:ISK/X2Q@SX9>)\fEW+U6PfT]4EJ7W+DN:F<PCIG]Z7a?K
g\YdE@X5,IgEGA61)0V]Z\.3_/4_MaG>XQWI;Y,P>N-?.N6U2@YfN<7.91C)cY61
55+>CZ7Ra.?B0X=Z,_;M2@<8+8CRgC=LOGJJZ3IU/R49J@Icg>dH+6B-a[_^&LAN
>D[.HGNM84DXa-\:F=V^_=MCE2AIJUH,dYN/7f(XZB--gad284T3(](3]83B:=b/
QV7g,WDRDY,efb])2T;M9]L[8^=2b-AXE8@I&>W(5O;f@.:b8,IVB1CT-c^1&5B;
a(O,Lb6JK^C(73BN,EG.b]XVFa2a(.Y&VJ1)ecI=?(]b[[&Q8dfd5CLJ/7L&X2bK
K=5@/9R^OXgK->LRGaIKf7.H^GK;Y=RbPe110/C0MI@7P;_Y?.:W5VabNDRHcJRc
[JLBYHBD6NC^0R&g=d_^5W:1EGG0;:gI2gVZ@>W;)0L5=?GaT2fH-VW<\SeV]Z<M
-<2>cKC92KB@adI:W/E[16C2ET\cX(a,D\<dPDJe_M6Y=KZWA^#,\/GWF.G02JND
G.Z[H05G2..gbf78AG-)+BLCR#]K,W/3.A]3M_3R:_V?cP40#:2CQc9:G.Q=JPf>
@WAHWH;[\MO9F>-97^@bY2M^KM^f]^+Z7(#40O,J#8M3-4Mg16S[Y&9Q\g8.#K.H
S?T18a.<MW&QGIWQ8Z;VELaTCXccUK<a_;@0B+@-e<0DQAL@@7N9M64I/dZQ(IfC
#+^=D^>,\GALIANM:96(R^[T\>(a7R<=HJT4O[>+fFT6>#6]=-;D@eeKae&@+YQ+
B37V_5/2WQD,W(TPJ&O)N8J/a\NfGaQ-1Fbb?G;c^\+(#1.+:Se2]BEV:ZY#TD8Q
0U?H0ICd.G4)E?UPe]D:R#-;Oe>ac&:E[3,:HRR.Y&=QOe&Pf]=94gC]3H]]SOHZ
\\9=B<<2M0YNcYYI9)JE-H>/1T8a8E?Q1LLTcT(dJ[HEL2_S;S-NEdWBB)-Q)dF;
dXYZ7O4Bb,4<7HO193VS(C=Q<XM?4cA?LS.6.4[_,[I+FOP>&5WQZ\KKUM8&;)D-
??eIUc1H1AEa\ES\@0P3Y)6#Md>G7-?P_;DIReD9RON]5d&gIW>:<>dPd:?PM[,W
3W<+QBE#B&2Tc.5L7(/DWZ#E;@M@RW6IV/TAF]\\U+\bNFKN,\/Y1+J_5N.M1E1)
8d#J#V</E&)_-.c?[45]>^/C60#5f(/6bL/NSc?&>HINLQPO@->>K=[:3(\;W9)2
9d)7QUJ[R6UA@Y/:?#EJ:N_P>SHW(JZXUa\+D3)>O+&SZR\AGdC1;INT[2<M,YDO
,d66C+5.R5;&dZ4ZIA76&3[W]0^gd,8MIXbc2L].9Lc.1]:g9O52V.^._4B2MebV
/,:CF,.S6=/KP\A7JS]?M,S(GCgD:C2&e;94>?EHL#UdG-;_I0GRZg@I@d.e]Dgd
3KUE(=-],,W\HX,H0B&;c[/R-fV?3^H)?EZOFAddHUb3\>Q0D:)?/>aCLcac2]BN
K-bEW(_fVXJJdc(:OT9J:Kf..199dd0_(^QcEWJFL4S:=H^MW5f@dMR.PL/6T3&I
J?Sec4g#H0Z>ZOJB2g8I&=Q:dB./Q?XMc]R&[>KQ6UaSQ(ZDSLY\.1^(1M>K<Uc8
=c7W;HHIT6XXV3Ib&H+4GFCE^N2Q]^[bB;0_BaII:e(-,?&B3TOIRL)<f,3;7+M\
]MK&g@KKJ>-C;:/O.dFH\TN<26@_K46e)-S>:FX:Ic[E8)QYM92dAaJKMWHW9@g3
9LNdYRL&>Sb.M&A7XTJ\Y2-O<].)Nb@d4\U&P1<EbEEPZb:>;F1^C8eS;#9H,&)S
3>R:XOJLR7G.-$
`endprotected
              

`protected
.XH2X.f1,F,d5&&@SIJ3Z0:[f+bDUX9be:]JZP),\=IY1U;1MQ?+6).dg(NEQ4WW
W(HG5I8->0X/;+KEWD/<+2[^P/AV)ZC_;.+K-.gU0>9e+S8LOQIDdO3@aGVER65K
Nc(#IdAO0PDc>=-]4R]R-3FF&8QFEZ+((dOS[8^5=1VP(6IcXH^T[B,8=,U#)6>6
8R#f/M?]>U(><<9=9&f]4H17O>fM@#2E&F2(EI&U+9:ZOF7ZY<J&&8HaXf#7cFXU
WT>GN1E6FFWRcMQ7c&]Z#,=HTJ80R&EbZ<97YRKCC,P&0B^PVIdUB^DB],,B]GY7
CLCM:&e7ILaNHNL+7Ua2^F\R0A6?_A3M30(LV/=6(:GZI6DFYYbHGEYU&H;<2WZ<
M\G]e?#6MgNZJG]dKfU64\F<\.#P4Ha\ZB;b3WPf4Te(gdAUbc7KGRYUN$
`endprotected
                
//vcs_lic_vip_protect
  `protected
bK-]&Ie6DFIXN]EWR#ZJHd?:7K+>JCTDf>S&6\^YJJ;4D<8.M8AD2(?=MI8/c+4E
Q_ICfD+c-#Cd@=]]^SXP<&VBH2.RX6,K+fSfNgE]b,SZ,(a28T,cJ7Q\e_6b_6M(
6f3_9CV1X+N+bgAVAef#8O]HSGc@J0eC>3bNG7b/);_&&<K)2VcD1VJZZO1VS;E:
6SEF]\LHG\A]0<:?]P)H1H+0]Wa;)L=afYb8R,5-@8E7,gO>_[CR<bg0bYS/T,E\
Q:cWBUQF32TQH(&H>JNEeWK#KaCD.H8Z?dgXJ@eTc@)A[,H:RcF#Y>3^dST(LZK0
[&>TCP7RERVQ?8?I<cVRPK:3gY+b8F3:ML_Z;L5B68dK-?P_NA\D32#SAM.KTRLf
QTC5)a=.F06YQ?1FR==&-/-LeRb<EbVg94I2<TAfc.=NA&g6KXRYF4B#,Y>H].(F
(N@]K[HS7WHUR?McG;Z/e?\J:)1G(B&3dbZ8_d1a297.WS7+9#=b0/P&7=4X:Z\^
I/(U^d#@U?MfB7@AYdH+#.+gQU(Bb:VK[X61E?75L1D069#[FE/G0B]1LN3=,2J#
OHa1<cFP+,KR]Q_X[^;;gJWB88_ecWA^ZeXW;&58XL<[TRO=,HVZB_Fga<^+QUB5
0@=,2UY]J:(&,Of>DFZOLS(XY=5J[5(GG9a6g+1\S[(4,?O#)AJ[@:<16RdI,34f
J;1B.OT=4aD=-CQHfc5fON0bgN6378L_GPTLcVbJCQfOP5:TSK+INgR+AaF.&bR-
+6b5Pa5f149a/<bI?H5c\#C-#0Q.K[4S-3883SLL&6g:#B_6R_I@<Ba(O6\SO4#X
8>.3[@Y7Gdd=5P7.4G.C:UZZAf0AC^QcVgMUA3a3OK?#R+-c05NC@WW4E\U:&WfY
&>@8QMgdKg0E@@HfM=>NMRCE48/5H7M_bZ=Lbg)[<_P3)G@6,6Gg_XTcX\_D<(b<
Bb.dOX8[AFM>7ZW@MEBG+#0gKZXUd#?+<&T^V9Q5Qa([Xd?<AVOXdQW=;c;YQ9T;
D)X#0F9/;6f6O53?Z6)X?9ce&@Q]dBHJ;KdFG8)<BT+7&WM3TA2Q<bMNTN8/7Fa;
4D4bb@c&84Kc@+fN0OD]],CYDCe<P,/3F/=;BTV#/<K3+_:bMDc8.OV8Dde4Z7GE
?<B4bN[@V3&b1NWb4b4[aD+E[T=X/RS+&^Ef=L[2][aURc#&W4:UG+E3^.K+cUZ1
\S;TIMSbI_Q.gN;bGW]5>NS,BWRPZGDVcf]=f,3H@)((N.>&<+gVfNe5#DDG-Y@C
T>0\I1;&>1/K_a^M<_f7HXe]?gW0?4.Kcf-<^&=F+7\[VC=/Z^A7dW9N5UD7:a)6
&7KSZBg/6_9ga-Pb):B7M8M(X.PJ+C]0QQIOgI76YM,Pd?@3N,3F#JP#TX<^Z?]Z
:V];J1A8B>P@HY(MZIHNTM<E7\FX2GB&1#G1TX_4JZSQF6W]+BP;CbB;T&U>LX2N
]@+^KP(eaF1NQ8+;7:7+VZ@8b5DQ\eLG_93V@.=84XF87[N@bD/Mg^0dP:;D-1RV
NHLZD-&Y:_EKO7X3c03/:\eLFVe:1cdg-1PeL)gbdd_L[#BBLKC=6A<Je&,0)G,G
b[-+&/^3?<W^SH4YY6ZC&\XH@Hd5:W)1_/9KRM[5OM3RZ5XfD<gR@)0eg=G,;VV:
&XC99AR#;4_W8EfBFE<WB(^1O1#+;&:D&JP,N3,Gf(TNN/96ZW,#HHIP2>)L-?3F
=XB+;DC/eUE<fR5Y7e)F^O-O(#+(S#HV7I^C8?/P40O2X_,bOUDaQTGC<KcYMRdQ
_XNAWBd,<cNM\@D0f5L;#K19(Y&59F/9^N=e5:P]8909AeaAU?=5T16e&\baQQO9
.RN0IDaX2QeBY,]2U]_D3WCXd47<:8GJbI/LaK]f+/7@WIN7(T(9T7Tb49I>:,Df
J+Y\=_dRg<]/J^0X^NPS]LEL3\VV9Y\R[-H9P.E6LBN):LUfSdKB\<B2b2F,22XF
:E+L:Z,c=c1)L[31><@C?#PV0P&BVAI8^:(T6GDU.3eV(geg?80+R7053g(M<5KU
(P/?^G,Aeg4J<-\+HB;^..EFd(ODBCEQAO=_YKH;470d=/gI<B8<;-I\)VS)<)b+
X2FLBPD>7IU^TT0+9&CD+WJ]cE,66&AR,&CbY2JKDO^XMAWOML9cGUKPH16-EZ_4
Y/8e.1IY\\Ac0LTN=_](A73TabcGd709X#;V,KdDb_R_H6Ie7FCSd+f#S=.MA8,=
e\f8XL0]7/C1R&6;cU>@-CGX/,G\_7M/WX=J3^;a9,J.N.<;V64T9ef>YD:QT^M_
D(b:E&8_8bNVZFRQX/:YXMg^MFAd>PS8d?XDZ&.=UGWG?dL]6L(+:<Wb?=f-ZC.&
X(6KHKde,^MQ)T7eNN#;Y/+<:6Z#)ac=X5Ac&Md</,/XP:b?.A)2CUJH\Bb>2@?Q
<^WS^2,dD=c(DdWE?8H2E-NL:Y@U0bCC_4R_FI?e2JFU3YE<87f@Q[1bKQR=O.6L
]DH134D-D81?EU,@E&V2(P(PbDBc;d]:SEZ:68TV4#cX&3I)I8HgeG-U:G4McW0.
WPY]aWb43]0,T2&MR)Z1bZ3I7Z\UC]dSeFR)3SLa)P.daH7[g71f\GAU5\L<V:K8
#SX@N#[[0)0G+bL;-]UAIbRff#T9;B+L9?J>PX<]=H<GRE+^<+)8VD^HL;/gR92c
_gVNaY;,Y<D.1(:K11c<LC6;g^H>fdHAc6FFf__W;^L.YXQ&7c2+M4=?<aJ\=g[1
L:4ZW_U+-g)<C[@YOK6HbCG,C/>()9[:P,M?+O0a=F#U7Y+gAX;WZHMS]C@>ZNCK
9,Q^D<2\E<]cWb5>^DVAA)+P:IL/UgB[>c]VRK4BbY?.Yg(G>aYEd&S,QZ5Y:aRH
eU@&UCXKAf[AQAA#FSEEU)#VD9^@4.?Ea\6\MJ3?F+aTU#IZ.GTUE>Y-XXcF]?]R
g>7b\^bJI(]Z6F5SS>N):L,0:4JA7S:?@I:<HANBVIdNbECea.Z>I.Z<@gTD44Sb
=b:bGgA.J:.B?IbeI_7daBJ#f6Y69[(eZ^=V7#Me11]O#X)?.HYI,g5KdYDJeN3U
3T6.YbTa<>0^d1K?&)JF30,ZC5Sc,MA;]91QFeUA#IUCgT-&ZaTFX&GdG0K<FH(S
T^)f/Ee<A@2Md;B7FK?UG\0JV7M&X=/gSTTaQSQ.H4d0:7FN.g0OTF4Y/eU<FBO]
d?^HfSRQMLF?O&>Z1M+;>XOR?+,4V(+OI#La.f_<#N3e-KN?H7;RE#Bg2[e;@LJA
2U8.9]-W+UCN<VA0L6C5?\c2SLMJJYU8IJ-SFEV)8T2JU6_?.&fX[>\f<25F=6<L
#TDXUA.+LQ/FVg#d]VM@e^<;WY(W)gQ[UIac/E);LXb^a^UeXGQ)D;Jf[d.WOLg&
WD[JRa(\E?>-<?D;bRKNM1<_+9P70<Gg024fPWC;V55B,FBdJMCbA2FJA2)Ue<P5
,YE:b<KI<.RM.EAN6[D<b?:Dc))dcR66>,T[g=QU-DD[\@G;CLeB6I4[G[_D9<K?
3HR7R@T.WFa:<QWcX6X<R^G_.O_c\b<eL7a#a#)VZOWK1X^Yf)=:&BSY[b#.AZ&X
@4@12F>O;8)+NENKa)JQX=][@MfCO0=UT=,^+a^6+Nc>7I>30cEAC[,ZJ32?[eD>
8@160Z9JC<3<NZ8;+5R\8E)YIT721&O\Sgg>T7)49[JKbG=W]@-:HG[Z#R9b5SM:
HI-<8-/Jc67J]2Dd+)(8AKMTXR/+C,LS4K.)3e4aF412M:.PH]TEK:7EFG6C1+8_
Cd@bVNAa3R+4MN@\O_;W1R2aO1X2,:f?)P:&fJ@VE2+#bO?d_.M<;<+QZ080?S/]
;@T7NC3GCNR2C8D-AR7.eO-Q#O(I:eFG1&BI8&M?]_PHeD[bHM_/&Sdd3D9ZTLE&
:&OC_V/FO>>]0@78L@@XdF^.>CBV5SDaf]8>YdcZ>5bDc.bBH5)H5@6_eEIE8Uc_
g=P2&NA]3?UKg<,-X2c&1fFgBFeW/-[)7]ADMYGTWPa(DNg/&ISKggE?9:f3QVdA
\5#?e/]W63L[5fB7X[BeZ8#7>N[UVb]&MbZH@]RO@FR\M#S[4<LEg38WJJDR;08&
7C9M86?RFDag;--Z2a#g[O6&F\OeG),<M(Y/O,]48BO?FdPU<aYf_f1(B?O8W,D#
NI)F/2BF;WQ25gfe[&90Oe\a-Q@JEGO1^9+:6O0M):a8b@W<3@Y1:GS2S_;/<180
R9GN(-2R-XJ_=0?R@E2c5SfDBI<<YZf&W.PKXPaOdVQT<dYES<8&OD]7V<bBF\B,
W#,bgW.e^=R1KBY#@f:\6_;Y1Ia=8;OMN>M#:b:2BKSP81)&>87ZX4JFb0D/-UYA
MMV6FbdSMRdE6.)71;RZc.(PbT9eQL??_76PgSJ_FZL+GE6@)fd)D;[Ff3^;H&#_
_9D3\a<@+3c=2PU:Z03fFb\1<M-3[ZW2LE\\^\d(VTON)FAN\9Nd2UJW]?RSJd(=
XOZX1_^#@^ECAXVRIX_R:^=g,S\SEK,G0++BNTTFfRC0]61&_c&;?/N4W)eC/.@J
1eR7CFOf\bF2V5DYEddVYV,&?/+RR]#R;R<c)NaSeDP?[-B4a=18DZR]:60];.Re
8>+@0TOWbDSMEXG?0cY,;aGBJeE(ZSU?N593UKEZUa,J6P7cc:Q<.^]A0+EP?Q+A
2]H2.4E-LM?7C1#440=d]6KC4GG37T-+[)8ZaAJc0G3bVcC@^Va->G^7;X\RI/9X
b[<J..2ABJ>XZSNS<-D0W;d6^BE_FX/DFDSC.G,\M=0:V,)b?OfRE:6dXSD06-e4
a-#<)J;?)dL[+UI@3(^Q7/_gQ(]b0D&Q6?]^2SgHH>eID_5a;5R6M+<##6]YY4<W
gSXQ^K=@04NUQ1Xg9L>[2_3(+Fg\JS8O?&WgLTY0N4K7S.?,5BUT.c=C+7[XN7ML
IUebKU\[Z?GgIFCg&YecVa+Mc?J^Sg9;0g(6+-;>9RGD)8#-e5JOa,J(D6]G35<M
dV[YgQVV7HC8;HaA/OdLS:aXE6\aGAeASDC76OH)Ig(bNOU>=[^.V5.e3dX>Id[1
0)6XDPgYU,>78MgI32[R(8TU[5[2.EE\.IT:,ZS\O[WWV#MDK(6=[LB_b1XXe^dU
E8]QSWXU;?4A#FV^8SLYZR,@&V_E=TJa>2Ze);>fAQVeM1?CcQ=,g[N\71;5B>#A
CWe]6RX4dW(5a.dRQ&O:_QL+_\-UdbDXMCVH3JRF8]A+)2@OXSa>:De3\bW1(JWL
IHTY+<)\QP>QC?J&-D#H54HEJ=C:H(8WR^Z5<)E?H\G[XM[6(5,OGMDD,Gg=QCDG
V.<P#5E]YBdJ]#-GAg5e1a71.#^ZfEYfS.7\->_C.G0R4EU3Xg6QJM68>RXeg6N,
&0HL+VR_,W_H+1+d];VTZ0PBd1:LA0D,WEITKJ9I7-))9d[PE;W&3@((;<Q1R=^R
HBT_2W+Y#BE0ZL00=;VAg=LKS39#(-ERMS6?,[O:.ON@B0^MYX-N]TfJASK,[Y:.
DO0<3LW6Q6GYXe,.DF(O^_[^V5/,DT:.OK3D5^2Va4QNbG.d>ADB;KJ\e[f-8eJY
Q5aSVC(I987Q/<ID@RRcXGJ4g=MTTf5:R[8AN-.a6La#RPKB]3;XJ68c#]-DSIbS
RPXG,:;LF>OR#)]W.8)@@R\5G;c)T=X7X_6eHF^6,0XDBYaN\FS73)c@Mb?,.#L.
6Qa\M#;Y<\L9baeY8,SgW>_DZ&IX@H9SIOR,S[g]8311FJX;HB+QX8)WEEN(bN.C
2HRFU.].f\aJU7>b=2ICQ?3^5@Hf(64WeY>Bc]a+PCIe.Rgebf&HXf66QOJD<ZcZ
C\dReQ?3-GYOL\bH^cOAV01ET_W?@KJ(]N9_a=#/c[U\VYg2A8c:G]M-1<<&SR-W
9E21-R&+TQ7O0\Vg&RIMC3190,9GX2TS0<&fN2&4\[M\RFIGQ/Ad64B#M=)DUOe<
FbD5@=M?LcNQ1JI40e&^51;9V:)C,+8gURebKbQR,2]0,5L0@-J_-3TXF#AY=JfD
5X>J<DNI=>_7CgR:M4HPKbKa##DYIUdb1I)0J)B>[DIU9Y+9&[eB(4d]#85GXI4(
.g6,gKIU6-2NU@SAfaP#<LC9fXZ>g^PTE[>fD^?^+.?^&1BK,P.86)BL.efDI]+b
gNZ>5L-R#^@10fUA.&63:XUR+ZC&0<dRF7]BB1E\6cZ>Ld[KLD&<M?TWYPOYCHW<
F,#+(+<218ZffAZ]]9[aYdC?K4(DNf\9V>[a0P4TKaP_A]?#OS7aS6&SeU#9(dIW
_,B1PE5L<[d:19:LJ9bT;Hg-&ZWP[;=Y8RAd,)Bb&,]@fZ.L^<QS=)a,W8X,8db/
6(D[eARCF==)]R2MK^L,(DY4b5c0;38QO9&;A#e5#CK?S2O2NK;5761X/0W<USS,
=,f]c?GG4Gc14FL(0c4B8#^D&)J0ddQ2cU4(SHU:Jb2EBV,G3D^,9T5O5(R<-_3R
.I=@1U-/;gcHS]E;Q24_)?@NKaf(SYdJMSG/H]-b(H=Y2ZCgETJXS[Nda68_<<R0
OION74B;?N5Q&E,0V9FA^WD_U86N@&3g7/Nc_4.;<G&BL:DF5[.EX3,5cXZ_]I)H
O(A1NMX;GS(4Z<aP7I2D69KUN[d_/Dd3JYeS&YEgeU83BW][IVS&EDL3<ELgZ)83
eV\5#MJWGD5VO#EIY<K4.8J0Wd<@10UNA979L,Od27J&+BB+gTF>R=\+E/^);g]1
gLJ1.<JIeQ02\;_B1)g<2RG)01^=5-3C;+U2bT]Y-N@Ed:06FVF7;NH_&/(O@Z[#
;E,e[D/==YT1fNF<3@VJ,IJRfHd;#Ff>LT>=3b)^6?L+#cDLH8ZZGG^B8KR(1//E
=S)P8XB1[:=BO7MQ,:g93/d?-2L.76-<_GK&KaF.LKDZLd?g4&3=0&M78=QBIA3?
KT2b9/287:TPfXAAI8D?RBf[U.7^)4;@DNNG;[#3RLRcab)C_Q)^e^5&-0(@5G[V
eUggUeJ+IP?,5HAW]R7F0W<&Y;OadT0QS]QSN@fSG4EI=XQ^HM:Y[C3>V,c6R#M,
9XHS5eVXfbDA/U_ZTXd.+Q7>KNYeB4XdH?fTYF7d(,>DcQa:IYS_SGg=E]Q;DZLG
K9M(95#0aC5@XC.]ZcVRC_G5SX]g0<dSa3GRU&gU88D<C4=?4[#96d_3Id89[TbH
+QMX,-N,5R&>\QE9P0=&J._TYdb/bGKcM&YLLZ/AG1^5.5K[7RBc]U;RHO=0/Cc0
\f#Y;W=,_[\cKJMKK-Za]5CB]DTbREVe@@LeaDVaV4[0d)Mc[Q:D@;S+e5G<dSIC
gPHN9N:G>HAJZa^LN)4=Oe-b[6WTMV7J&.4@9a57P@FLO01>N+CA.VBK#U@69@CH
G;),D?Nb9G28P8YF#&c>dXSdDR@:A_Jc7)[?aVASQKJ@-CIYD817):;WGaK^B8^N
;,/V+a3f=J:?K<Za:)eVGFE98WK-YI6JEE,b6M39c60S^]<1ATS,6FcOT-=dfL_Q
4^-7bNEC)I8W1RG&^f4b#&E:;(5C&4.?;O,9#Y)U1]C^H(W\fO;[;b;C.(R;B5_@
3VEe;gD<C_5+&B<GR=bR(Y]D,ff[5A/;>>.9N[cd@CXeBSO+5^]AWKUI=B3>Q=fO
47e&>UM<PIEYHdI[KX-;=A@=O9KUX3gFE0PMNIBdI5>b].U9LIALUGPL(CCG->(4
9M,C::A6=^Z[(aEL?WOP8\g:E3BTb/9F:&<bET+eGdODWBONL7c7UT)\gO?\ZgH<
ZPVQSZI0X#OYZ#\[-T0gg:E09G)K]/>fT,;c@e12@<STaWGITAN#<<W^@OR3WNK.
V5FRed]-&;LS0ad07&g.N[gSCBfRaJC>;.]\LTXRJ)H;C/AI3G7L.5Y,TV+3LEX]
2P>Xb,Y,3G0SB6>4HM+[Z30>6@YLMV[LJ)-HOFNIbX/CKHAPd;J:aSK+_QQ,\eXR
JK#ZAU7.W<A+C2O)Z>3:OR96f-[a\0PAe40/3-4BM3d4QJW:L3SQ4OC1^?G43KD@
#]^gI2ZVgJ^8FYT(5>>.R4:N;O\PP/+3c9OHW5CSDGC)P<B)>\ZL)T+S0-\e+0NO
G()[3W(Ma1+8@Qb&(QI(;f;?(&eO,(UH(+TR1F)6B03;;SeS\ZPOEEF@7UA/+7;T
&-<+<B3ZO+b_dQ;LHM.5N9T::g+=8_AS+FZ@9Pc6>7EZGQ><.9-3LU?)WaB5LeH2
NQREd11O>b=MW,:1U<0;OB-&>92d->PZ]UCQP/^VgRV#>-9(Y<<@BL02855&)],A
@3ZFWK4G\IO;=#@0?FXJ@U[UN7?Y/#KLaREM?6b_4T8;QJ\,Dg?a<E@WWDZ2\&5g
+MR6:I4RTfA7E:YZbGN;,SRU>d.J3G#7\-O(NU-912J;>M-J>BU\;G#[[2Ff0fTF
WI2MQ;4_/40.8/^M/E1^/Aa8&CGHRUH:36PW4E0XeSNg@W84F5fV:NC_ebZJ3)=Q
0>\8PfD_PUDE[];4/QU,a4d=W@&-1]Tc<>G.f_6U)L=@[bX;QQ@#A#af1X0f@.I;
&V)Q6JICNZ+e-GSI=#I6f6e8:fM0WJF)5K7#C.QQ.Rc-1;Z=^<0P//>MY<Y24GFL
cH=4W\7NG,QPB;,M_7+cb5Z27DZ:\6S>W)+>H8W+FAS4#MG0_//F1MdN0@W</9+^
L#:deE(;D;J(WVE21\56#61?N:d[cBJP)JF&V@QCca1H=c-7(cgHA:S0]1P<:+FP
.AM4JN_ET,:Uf__\_f&,5VeC7;1YFXb&MUEVO,RGb&SW4G^aa5.Z?_VU(]UR,LUH
MaMQSWP&H9dH6OSEU+,&[\JDg1>H(P_(_+QcYd7AeM[\LX9Q:3:NDKOM\,gQ@ZDW
5_BXE\KTL=BgH)(?6K7Z/b]P_aNa;MaQFJT#.]>W5gTG_AI8LA1L7Hb8H>>4cgJ>
M9ca3#2QW,(Q@?ag-R+Rf:b[>PNFc;/dG4M)I#)#GJLJ=STY?G7NRD7YCI63+@H@
/?9P0K5b48L15XW;Td/^P/0&L;I8F&dgV]8PE9V[&Y1EJCRXWJ1bXbd2]ca-Bf>;
aB(P4;OQ.=N:J+MN-a]ce7_R>N7N5I,4M641L+T/C1g.g,Z9(eOAK8/161IdWY@T
]IOD=_0KTEG(T(^O:Q;:QNYg1;<GE5Qa4cK<<<N:3@.>_cH@1-OG>.[C\Qa5deV;
,W:O5bJbIN@AaS&DfKEb]gg<9)/)0/WW044STeEPaKE6V5e0@K9=4VVd;[#SJT:H
#Vf4M9gA,S;.\fa@^<dIX[9P]O[VW84ecOdJfOZK61/K92BG8dIeOedMf19II#X#
+XcH-bZge1,&La2]VEcF3[g[)70=CITK=GO<@+/T_B&3cP[J3H)645WVK4:OTRY@
UTY:1deZ,d])\IZ6If,>;O=0F=eYa]>BF3W<6;<3^/K+8-0M[Gb_fCOWJ+H_673>
-ACDg@Xef2KgCTU3;Z,;1gg\TN>Q;-8ZZ&M,^;c&:QSea^@3>(#Y,[#:NR@5b&#b
?)LOSNQF/)M.//gTYeJQ>BPWRO&7IfEfMgZ&C(742#-,18IXKE7:O4=?>+&;;9Q7
VLDH88>d_8L22IGbL#Ze/HH#a@YK3?dX;:<^Bd7A<]Ad2S>ED8>7&2[ZRE=Pd)_c
f;N]3F)bKKY7-UfOEe@6-4UK^/T/533)@0QdYcZ;;-B-881T9^=O7#>ET[08@c2B
,EeOTCTbJZ/D2eDa<B#B[LPa?+DKTJ5/[@b.YWOS+FO^;d=b)fb90DEa?@25E;(Z
;KDO]B>@5\=#LY)U?>e)bA?QU.+UZZC7T3DP@XFKHfH_R-B([[Rf3H>.SW[,KFR(
aIJH9FbW=NV23fHV&5F?(f35dZA].@V?+3CU5<[)bJ2W,E70#EZ6.eO6=#2_J:Aa
fCQaTVI67/P59ORbKYYDXWOfdD_A0KT8[],L5?XW>EG@=85K29Bf-Q]Te.0)MIE,
S+RB[cC:^MG>1U=\6JC,bQJ?,?E;]?g]5Wc+>[CQc2b\67A3YMH2KH,c=9,Pg=#M
.WJZ_(^,.d?#?KPB6NOS;W/\P-.@ZOaLN,&FecFVeUdT>F@b>AA6>4IE1Y^[HN.<
[EE5aaFfUK:RPUc&/S9e-M[XJY6MYd]2AE/,EF+Y<4d/+fg\Tf,X,A+,?Q5K0QP8
7G3F9N0)@7EPZR#.CN43>0Z\N>1JOYH@;+?R)N9<WU=2>7=T.X<F=N0^JP<Y]K6P
e+dd?=^)XOE+LF,RVag8FN3fNO+--e#8J-SBH[cFJFD+RaYeEB+9:7WKb?KD9e_T
\(DI_G(Z5SV>-N.?W_AX5W4&b(:GHX8S@(a-X[U[&<Pe0]2^Pb?Z&J&O^WK/B.H-
N74;?D8MHRDET)U[>bZ0OHTU>#)0D4MQG16W&aNNFe)bAfaA+&aB#Je>H0,]VXK0
bXGYV/TQ5(?,AE:9R=c?^PU&=eIb1aUR]f8V-^#D#be@g:.8eJM@36_(ZY#;R9R+
=29#1<=T7O886Bd+@VPG4WW.U[U#Tdfb.?DK98fKW?gR.6Jg2H_B(2E8c&M+,EJ<
RXTFg;,:G2>V[;:=cP[(\2U-@:_3>XVgL)WC?S_,E,])<+cAN?e@bI;C=NOF2C[J
B_VAZ:;XVP]Ff_40=g>CWAXQ&RN+7;1L&M49T-J97W[AC5]59ae/X?CB4+dGKfR_
5PB4G0KH=)e17Q1fL&1W>a,5X:[NK>_&>L;:L3JTI:05721+K4C>16W56eGf>K\E
fV3/\H<XQ;Mg;U4H2V9FS^V#>ZSA..V]IO[HR6P_T)b[/cPOT>6d,<-e]R]]^DCE
Y1be@O,KMR;.8):CA)4Jfg1._+.P-J7,F<dMUSN1-_O,=2AIK>F<\F9(=ER=.X)0
#[6fPUN;)aONf8:)M)&N98L,J>PDfPP^EZaAP;<4aEFSN2FdCW,TF.9Q3.XW9<bU
=GRQYX.MXU>8X?ST;=^d0+85;#2YBOL+4aCY/D.aP^S2EP7#).1.9d\X19)fa81P
,VX[bg\FF4K@cLOeS6H<NMF(:IQ]H9M#Q9SIWGfL9+WLGdZga0=TILHQOBX,dZ4D
-B4)A#dfNVA7cR?OH@G;\;56[7VbW7Y7aJ\DaHOE(RPPafMV^8W#?AZ]Kc&.=dFF
.52SN70RI&BSC0?99XFB=C0CP7+F5=E9DQD6MUEJa&3R_AE97O&<VYb[N?39W?^6
X314[VIU,R[3+<fI:=CDg]VUFQJEZ=C(:c7;fWG2e;--d=D[_cHATDcGb+)FDSBW
-2VGYQ;Xb@,+FG3gF;UM)V7URg:g&e-XfUVR(N54c7P4OFV)3S)]:&6AYdUK\afb
QZBVQJQL\Y_K/T4L1;KAc/^Xa-?9TN(+c5^+?[6,4\fPd4aPWW.UP.;]Y_S//H@T
A/UEa)BBgESI3gQU-3ggK]Re-GV=aTD/GSKBBO;/;152W#8cH>]P/-f;5&:.[G.g
\/NGdCaDIUV^NS@?+f3/Z.7<OZ\5b1b;<Ac/+?HQX,35?9K(JM[Z\E&A,fWX,K5N
R=GW8VOXc?P&CPH19LVe(YHa2)@DN7ZD\RH21>Ye]LLZ8Z++#JZ=R8(,WdX=P<JH
e1;Wce.=<;bIS8-B76Kg-SVN#:5?)KKG+^O@S(H3HHKGK2#P+9#WBJI,&\J)@d1/
XV&-/0KVWd8S5EEYOWD9f2H//<H,6Q=]AZP0#2Z3_0S]W2OOgG[aIJgbF,Bg(U97
0F-5P7A5bK.f@_L]ZY^3>A@X[dOdYL47(TXV._=^a9P?OXfY]VSKB9(UBf-d>V>A
Q\;+KeUQDAgTb;KS7:244RQ9M=,EI?[=ILTQ1)^&D3N(45g)aU.?W[OI?W4;;J(R
8cQ2;,-NM56.QX0#Z0:HM3^HEF7?^2:>&@86S+Y\ReS4aO]P0?CJE/bGY<\U0ALO
I\M5E0T23)g(S+.Ge6:#/=1bHbEC7>bA:8.-Zg4GQ.0TN2G<3U8Q,3YSC1e>)RB@
X+aP+8g_67/U9L_7_L@VSX=+C(YUJ87A6B=VA/(7=4XH/MJGOGWGTLf7fFd0XRX,
0DAIa@M35[3^&1]9^8e5.O3SUGYCc)</_ERFaS[QJHcWEU+=@&bTgZ&0B4YN?]UX
7ZVZR]R2JRUe4Hg?#ROS.0&T#[Z=4aQ]4DNL=]HK-:E:H+NAKGNU\F1EL6M&;+TX
?UH-b_HK6D,a#AN;cY+GU1@6K8;+MP2f8IV6c6=E(Ng6M<a.5ba&LBFSEFV,7;41
I:[-0-L5C:YDD<d@WQ8HPCKU/0]b+;C0</3=B#?6(<WGJgIZL46U3LX[XMc_&4I?
fg\J#4^LbGAg]d30OdIM/2gXW>.(O]HeJI:F,=JY=;J.4?Xe0AJQQJ<4F,1@?P.Z
FQ\:\7g(gK7bMScV53\<c]GIdU@I4Kb/I^3NH^B^]@B(XBVY=037S;8=eIW/10Ob
LSK^Lg7(b5f3NT9NL^3W)aAO1)=TDBVF5?^27Z.=DDOT]bT1T22_B[>c\4W1dEOU
FF=D(,P^Q10F9>:H2[S?JAQ<E#G:\KNU@gO8,K:a8=X6gWfV3e/B;e5eFO]D;,J#
gHY6dZ5SVdS]J4>c;ffJN7ZQBHUNFbIU1:;S);GO86V6@\d1I>&KQN13Ac:G<)6#
,#S7^;^7NPd)3=77bE6PKBCNd4dcg^Ta+)E9VVRg+[PQ4PfW3^>F,4B-X(TLO/;A
C@8J4aaGF^BdB6S^U\R@,\ZaQcQF?G,[22UY;VWJMM5WISW6G2e:dIKU6XO#YQOB
WXEW[S.YT.CX^c?6G.@5f_^C(,U^/F88J4SR++>^2\&(@E^8SHL,1fD&T=fCSVNJ
#KZ+/AXW_.98@cJHF:6C&W)=5G<0YU[;eP^8fW>ZQ]U,X5g[8PWRUfTfRYRZJK98
#5RRNN;;K9Md:g>Nd:28b_ANPEa\96/>b2U,2U7M3.LDCc.//J/6=:3=UfY19X+c
X-DHgY+6+PJL8GOO3TgEV08H+,SUfM\=./\7.b2.KJE6-U)]1V/7eZ[@gS<&f\/4
#eM23?CY=W1I4@)EGJ1M<47fVCa;AAb.^c/;\<:d0DUU)VQcdH29@a7_JD9U5^N-
6LK]OU4c,T2@7<<XM1R<^//XIM_LUUf=<TT19#U3F/T,8L/B:YWG/XD2BS6d<,1>
:+:J_-d9]d>4)9VJF#>1K&S;71bP:.0=XRdEebP3D2P/NA(]46[MLH=K9feYMV#@
b5V-L5ZF3@.W>b\#:4GeB9K_/d/+&E[\Ef2YNQ5(:TYWW]d/[)HC+8J6/]a=c0ZU
D>5#[Df&PA38AF,c4]:eJI]-#&WSJ6d](c#A3,R,3gGcKA?f(_=\7ecYc>_PV)T_
R45g,HR:?W9+MOXCXaZ).X([3KL@XLaFEgO.U)JCd&H?>VH83I,T&@dHBUJO)A6V
KWa1YJ7_TRR?X:?D:#e-T7@67)SgO+[Z;J;J2a2\/U_7=,+9e\_5L.B\=,_g9?BR
KFAc?NX:N)NEPL[UME-[8f-QQ9JIU1B3I&Y<83\[#W/NBD)0V_O4.>;3e&4QfX,g
F7Y\gU6O]M91>J]9I-MY?8O_+^G^-W[2#,<E=gP:Z@f7K&71d3_fN&Y_@g;,=PN(
Jc1S^YMc8AgUYdV<#^A1JH,3[<S7_E>(gE4&f([[C]Ve;PT3Lf,D<>DHM@GQ/,da
;;1,-Q\@1)OJ(T;a^=)<+D6()H)O1+8=Ad?IC-KCXC.bNT6H(LMZ+?NJdL<5(43X
X(6VV-.aY36?dQAY:O68UDfD\&e[[/Q>WZ\JF;b\cC=RNE1S\c<V\^UYKAHK^@91
)?CRF_)7)G;ZC^8[CUdSbY(XLNbH-9cX?C6_fc^55R0AT1PFHWM6\32=UD/CgKV+
][;T#]=F6\9_&FLV)T1+>gAfa+G/?ZU9XVY^D\,QM&<@HEb-1Q3Q7@;-&B/KZ@W;
1SS_IH/M;HXV?d34P@I&\1Z5]@P(DL@[P@daXY]gMJ.ZJ@.R>J;E@#\^PfWg6@d.
C6KAONHb>>:+8-eIP13b4W,c=d;]0Fgc-VNL5TDN17?U+?aYY-UD3TWG@aBa+N:(
N:_VDge=J9X&[IC>(_TfW[L<S56P>Q>=,dBRI,/AJB@OC9Y)>0\OS^1A>:Y>^)8N
D>0?fB(,S:EeENH-J]ESLg&P):-N5S]NR;aA=d6QXN36cX/+S<S,=]fGM#JSD73G
+JN8>X8MC-VG)bgO1H^4Z=FM@#<cS==RK,2^]XD=MU)=R==62c?eY175UYb9aJ6K
0g]FLRb/e]<@aK@8@,G3X\VSFHT(GB9OSYX#e9Y=4TZ1-,_EWFc>.JUPMY;L_]aJ
FLI(U3d@SFP@TR85d]YPJgScU@Oc@Wc0E3S\?4WgY4I1-JAS?NO^8Y-79a1eCQ@C
7N=JVN;I37TaV:Q(^1M(FD+WRC1IK-:H8K\(V7W4ZG:]TATf4Z;2e@Y;],25Z/(f
<?2Q);Bd.6<G5.@eG-V2\Ec,c4:]L=0Q5+cTBZb_N5@+,+aUbC,bD>2><OIC.N)e
])5,T27I1+a@SYLXA9EILEICgS7Lgb9NBL7EKG-cfZIR8K(]5\^4;dc8OYc:S_.@
Z<]>BC+#)&T=0[MH89W-bQY\00Q6_1XW39^2J>9??d8Pgg3H@>R8a5.HJ>Fcd&UQ
H5De/QEH+7aPSC#I_e-HVY\S:Kd,.A-HBUcMEScM]=()<(GEIaaX7Z@2MOCZ13Pd
SN39>O4J6+]+XE8aU-c4XEe_EK?^=Q4\e6?DM0&WE(gf0N&]b-26Y<59YU5^^[=5
@,?1b6I;CDKb0I#aPY,X[fWJVPX(Pf7,=c_,PL&ED4f>c11T0gXe0bM\\TH1?<ZU
#a7Y=QXRZ3OT(F#I)F^c/JeG_1aLW__-];25[]^+g>eaE/)FMdHeJ4&IJ<XVZE?G
+[1/(2d_AJ\KUI[1V,.OZ76\BCXO9Ec23H,[MGGe]Z:d_(dc>R;/H1V.9LXH7KN[
eX<+CWQ-89eWE-a7RcBA?/&-Yc+N<_d6IRJ<9AOSB@V+_8YI[2>bI\(bMHg)+2&M
;\c>BdCG[CT_dRM3O7](6?A-fH8YPSXa3Jd]U<7&Pb,^C[cZ&&UDV^(>2.D^GdA(
9a]]<+318Ud415H3>W-gdfL>H&59YLK39/3e,9ZK?2C;+K1Yf4/B68V>A/3)Q6]@
J=,R6c>?@,EMQW1C?)O)?JA)P@B:E.2I?+H\JNCYOb2YANb@WYR-1]g2=<IAP=Q+
N)8fX:K)L#e1XdT(A@U4EGIU12Ca6B0JRFE(f[[TEf>)G<O^DNB5KFQ1M>bYB=f3
(2-)VJ9#I-4K@S-96H]+B7d2K)<Zf-gG<W6A\TFfC),[eD/RM=VSc?-PDNUY1SH]
O<;L]bF;)1HbQe442#5a)B8eS_I(F??]8O2BCJ8-,)?D.GWF(K.[NI_N#++/VBcb
T@eJ(c6V66bCEWHf>]P3)]@gVU+HWCQ<B0DRgT6&845<,^d0>PD[9ZK3+90MROMH
DWSE]UOTbPNVY/L2]EbZeD2,&LY+(Egd1(NdIWK>\KYH/AYZJdN)9>dd>&Z<9NaH
Ye5^#4QTaSN-b@(_6QEN9-TgNQ,_c]<(+)]9DbMbOZPHWRCZeJRI\J\cB^aWMO4^
[<X]+)[P-dKU>a/3)9L\8_0/Q]OQMJ;Ig.)UA44,\M=C7EQKDZA\M4?+UeX8eRWK
aE(:gWXcb/J1Hfg,#P2L,J&;FB8-.?X]&FNZ5B-f^dWBCf>3_O^&/,,<X)ZV&Y?R
5b:X8WegS5fRL18NA1KM[0b6WR)6Y=O0]Bc)eH;CXBX+6G;B+32?cQ4MVC[LfW(9
PZ(^eVb#A\.2U1+JXLX4+E(PD8RU^-86eNG_^HS8ZRc>De#f@LCg;WKWZ7(E]c;]
]RIZU#4GOXQKCfT>/C@db5-:/Rc>J4PMP;V=Z^3_00]:eKWE4<]H0\N6K+cP1FPC
>T,AJ>?DNZ]14?B_LH_/2JNB+MMHb4VgbE:43fa.EFJ<&465gK4J7a+B9PWZ?(66
dSG-STb#(S61(?&_@P(OeT@?Y1^gHDE613.e)CDJ&2K50K@)QEF/KE+^S.bYTf+&
>&61.@cf+@6M(Na?TP6cA#e+3HP4X1>EYK60>\<]:\)f&ZaXAV?(d][==X<CNIDP
U8.6(a&IOU@)[8JPWF\MO8(OM[X\F99:IQO[+d;S(/5<Q\<Ve[3^IBTb04-e2F@0
dT7BO1/5[2(1:Xg(H+BE=1/0;U#M)D#_+FaB;+^KN4,&:?-#aH_,<>IOUEMW=aPd
J/F(Me314[??H<5(8[0aN&-IW]H13>0]T-5=#(gGV7Q^7R=7]:M&IO^bg+@FC;Ba
QB+&,)0/@>@4K\gH^;B2<VTV:Z\N7UMeAcDF05O1_@_)HHF;(/?&&=9<E.abSN1?
;>R]#RbK7cT22;#Z-DKgE,<L\_CR>42M-cZ3<g<+B[B)BO32C6(L^9W9:24][OP]
Kb=4dg2M>1J#:dV#B1)(eHd,2_@,YH0:92NG9Q&>a#\Y_1]U9B=eE>=Ag^g[K/2f
e,U8R?d<-_Z&8?&DQ?RU=6Y^Na+QF1/K+]=82YM#aXFC>FIVUeW2F2]F_7eF_2R/
AdS03K1c5dMNbRT/04YR17-&PB=aG0>[T=Y;EaXZ(bP,-g7QfB.4TO;=BQ1Y@@WA
=:bTaA/,AS@<@I_#NL+K/SHOC]X4F=Rb0bbQMRgKRDA)3fXA:4H<@(c.eB6AaA#Q
<:[Z68)[V<O@J)SS_&4QPN]b1:4XWb-H>,B8EV29:2/=TJO@N3+HW3SNUeR,SLDa
N?eSBPTW8;XeB[XDH^X^<U+N?BU\[XQHP>EU#ARY-GU->NNQJ)=2D[&[D9_.=b<]
B534(M:.P:42N?=#=F/EPM=EgNc,?9H\0<?ga.F\E4N8K>PS\4+J^9Q(>61D@:T1
6EJW]]D8b8_GII@&e]XI,I_RfM0K+T<X/.<MB>.\aPIANX4_AQdeE9Egb(bLJ@?F
5\FcDTf:GW+_YSaH+C9:?PDDbT&gT5T6cMX)aIFL#+NgQ?VF1X/)W7OfZ,g]LFd\
FQUHOC,CDUbFJO1a=bbQC?+,d98SJeXT)GgXMEJEU7b4:H\@(cT3b<<]Wg#dN0Gd
D<&<YdYLORJ4V37LUY]36\C_Z,8aF_8U1YBU(3[Xc3:V:6&(.T_67SL0X.08?,A-
)+_@Z:I^S,9cgaA?\M^(9/VW@FUVH@N^a/>2R4]X(\0U?FIX::EMM<>,4J2M.F^U
&0=CA-_EW7Gb3(a,ad90(&@R>YHe6^2e1Z.8<#]<XW@b?Lg;C6;E;+?8HA_N6K0E
I/J??#ReOQWK?KU7Y^+T8cV[C^R/5+7GMQ+,B&DD7,A+7VN&G#f7NX(IF4LR_,6-
NK8/L97R_.&=KZ^/;Z:W-LRFNVg#F1UK;Fe&S_8G>-1AT9La>Hd;N-LB4[Q5^\OY
d>#?,,D>(gF&@8-G)>8GJ#+_g=0FF-3:H/+4>PZNE&_1W&5]X)^IXddCVU8IWK@3
@].V^Ne_I]#GEJ-,RIIHBfBMQK3\IWZ/UK,PX6HZ#aTI-=cXZ9G;ZVg8T2c7a1W6
MMU:SGI/]g]43]LZ4e0W;^;82E@6(;PLIc&f/6D6DaIID$
`endprotected

`protected
=G5VCG)HJ_=#f0:WGa[K/DeZEH)=1A[TLV=d;]@0=:QX4I9EU@Rg0)KW(MDJ00^G
3e?fT>,a7P-W:dg=A/KJ?,eZ5$
`endprotected
  
//vcs_lic_vip_protect
  `protected
:=c=SDc<)VTOg]9fKeKQ)[=g=Y<Bg51eFcU@5E]7/cSf@PWTYX7+7(T)I8RKgaC_
JM#<M^IJ:c^aEM:=D)a.]8;ML#AR7AgB,R=WGC>IbM8^RaP.Z+OQ)+X-7L5LD=><
NA&+URFeB-Ga+$
`endprotected


// -----------------------------------------------------------------------------
`protected
7fg^V].O..3);PX^/^SMRC,K2WWB.G&.DG9W\&33Wb#@+43[7.>X4)3\(8&FX]DJ
J,L.57b<:@L)*$
`endprotected

//vcs_lic_vip_protect
  `protected
-9S\3?]DURgKZM1V=X&Yf...O^FQNa_]@U/^53c9,TV_RJGDaVYF/(G94G7<17=A
LI>T7bdfG(Y&;R-K\SVD[6H[G2\,90F>\#[RB,0gfG7K5)+4/9/8OIIG[R_HRU#Y
K1@RT2<\SZOU=3C:0B/EW@DZF,:(&-G#ZTJgN0-Y?<N/SVH#Ccb.:KW1S1[c?@5e
7JA?F,eM=3_?YVB5/6WLITG2-V6Q9.+W<W3A=--L&Z=MVJdd>e/5U8T_=APH8WU?
&IYOGA]dfG&XO,RTLFA;2-bMHEN(]4\IH/f/@M>7;#CWeG,S8V<&PDeY1U&JMIH4
fW^8FSSG6gJbYA?dFbM:)e1>F(;+^WWR]G@VXQe4>(LY<4&[QIA_5(C6VBf)fHMb
H=.5L;;a_(BMIAb\1(@8-Id\<SA67b5,@&Ba?,->68QM;7a]]AgbZ,5@G;YY>#2>
B[;V7DaOa4W+7POfR6AP/\L>c6RC,Ib9/8)FMA2cb^Q5.\Qc,eBC1,G?+fMN)MA=
5AHg-@dKbN44C3Q4b1>0;&aE/].E6-Nc(]X8g._3__9fce:YE.&;A7O?&fXIeJ^&
fKBM/fXQ)8;GEB2SV\WIIE((BXEb76TbRFOMU:_@+XDB><cRg4D+#>](P22=OE>f
T6N6/AZVN=^\@Ygg1)^#H_#3=4A,&d=##H1I]_(ecA>DN1ZHd[a@FD#]W),]e<d@
A9I?g;9Bc35F_4Z;=baL>?HF6+Ka=ZV2#c8Vd5BTOW(,P+.[U]#@5O#?</Og)bCS
W9>(^_.M8b)VP1#52+&(2)eec@IA7)&+7[?YgW#c?9eKfS>e=31aL25@MH]ICJIL
IP]J:QMT,_0(,SWP7O?U>L7+>S4,<JYGY3#ECY0?)6Wa1WZ6:J.0=Z-BCMVccG>#
^6#?GLV9#+.)_TTEg6#+^DPM4Y8E=f_82(EHK5aY5[gf<Y5QSTVTLOZCFC&,,Ie:
_aV7DZ]<O2cU7Q.UcZ5W\QU&]dc\3#Pc9KN^)gQ@AF5)b+\2E<cO?I:\^8FAaI5_
)+Qa)5&97LR+2f6L3?POLSdK,9Agf4L/2/,G][(:_bXPWMdaEA-W@2_WA9&OORg2
46A9(N9R],I^]7M(1fIJF8141X&?JA;FOcePOE;Q3c2YT7^A+1MfJ&P;DAML7ZSb
HJB(,_J(M_#\X@@#BO?J?_dAe\;L@RG,CRd4;87A,T^N7?)c:5TcVJ;LI5g&+N__
=8=W3IZ06AUY3@=,XDVB/\#<]JZe,2K674FfgE@EQ&;9e2TUQ)ca]>\54Z+1GV]?
[_7#HLCA/B/8D56Ba:8TC-ON?00=7GPHRgREEGFNYWWQIFXXV7C6MM@=0O5?K2D=
GYd:BK@K,0D.<:UfVLV]NB?4W;OHReE_a7,YXS3A<Qg9g.C8[LE_X.&Y[YDQa73T
H.Tda/2M@D4:(/>NY_[&YG5C^3?BZ-0GCcHV&SeO@U/e;@A=.:\>_^-aPXCSV[c-
H-dI19V27Q[O-8<1K]O-T/\G,9HHFJ&Gc5SN^XfPOeBQ:E<fc?e(9URHEI2_,=1F
d;1Wc\]JYXS[@>CW\&KJ@1NIKdJ/Y:1]F7/+(3I&01OaOTR((a<66]Hf+RB-,3gG
R^&VUc&f_WGN(E:.11H?Eg=H[X2YgR<K&7.)Ig)A_OX\8b;BE>ML_(>_\-;+NN)D
507BBE-(+aT?A^9AQX(MH2.Wb7]RT]-=-;e>ZNWaZ(#5I^<_FA-)(NEY-)K@7EX#
gJ;I=1P?;g\=T&&AP=TA]AOZ2-X95MO2HH=:fC@M(PLU??5eU+HM9:5OH\:7@H[[
:&B,51C^3>^fG#QEHM]7/g2-)9YS/YH)LQfGAQQT,GU1V^Z>I[F9GVNPb_/4WADU
-QH.0:8JSA_)d,9<K;C,g&RA;(GW>OG#[04g=_AXf#5>g-E(b\O&>I1NdZ@4YX_-
RQD7.^-A.+>BG1U4VgKe[ZAe;eN+CG?d?VA,7IIMY7C2fC9:SH98G]<(U;-YZ\CO
@01()4c2\I\LG=;S[4MH?;UK2eI]0I<8/6]cH=]U6+1Qf\H6b2G<LMZ:)D)GQZYV
7MEdY,X@>V;@_d/]Kg=CQ+W+<0E#:W.+=F6OV^(e2C=dI_=:Mc8N5T,XLeKCBS@<
SABSZ,M9:C]4H0SdY5[0D.Q9A/95?QbQ8#3_PBZV)T)bUJQ\Q5cHUJLaR#\_4Y-L
JZ&g<a/+caZfTAZg7/QNF#V<TV]SeU,,((,cZL5&1610V/KcKRM5_R@H+)3b3<+D
#g8EE[==C[gBP1X7#1W3#4e#S?V=2SS1DC6#=TY_#fICaDA\I7R8S-0_XKc2[8MV
;K@cJGX=ET^TIWMPVBJAW..ZH8)A?CH-B&[GC:+>GVF3OR-e@/cbS5M]VF2?J8.a
UHDUW29gK3g\,CLSHY#&UM0MVOeA8??dBY:CU-YYf2[HZAHK;5K:16eN-J8JVOCb
B1aGXL_,6>Xee1gdRQ5U-g4AAbR[bFNUU>\\D2TQ-aG&(H]]9F2T4F3-:,/NVZa-
W935QU^PNH&a7gB_D(EQ2[e2],VQH=>>DMT>&)-^P=6)(=09P^Qd8M.Y?&:14&6S
aLaI+U</DV^F:<GL(]b;:6G[F_Fc^?a]TVW0Q_)Fc.aY_2)=]20@4aA/R;,A<@U3
C7>[8c#ZD,EJaaLX^g1,=:e9@Y]/>B+MA/+B16gJXAFb=:cd1(6())=0F/R1PI2;
6_S1ODGLF<:aO&/d0X?S^_]?@&ac0.c\5X;34C@,@P7=.XT]]e(,DYCY3<CT]F[f
.)50/6>Q;6OHX?g;+PGVA?-e75eJ^6,@\-.fYFW.LL[T?@QD/.2_HdHT@R4Y[3RH
ZaS3;3Q?XYP/6T3g3@4=be;N\@+YI&XcHe,GVW]U&T#M[N^^(b_/#6B?e;ATCDAG
55BTWF@Z&J7Y@e^N_D.=f)Z-W4(YL_6dOVIBUK]Ae_d:G+8JZ41]=2:#c39JG-N?
3^c=4=K)e>LCb_e:@O@Ld04.A(9SeeE5HTF8#O\&ZKBN9]G7f6b^I)E<3E>E(7RV
7dZfPcS.18,+W7e)],U:BROQ\J9BZ,<3@77SXPC,J>9WXgI@\d7cFRE?K=?3JF_I
IL.Z67.9[2aQBd^ZW?XNNG.V?K&87>FH3a<Q-55WdG(]HAX,>_F>AE40L<)DR]IW
0g<48[&Se_:CJ,fL4,ZH]P=_4T,WVa(5RGG7:9Ja6&Xf9ELK_3Rb@DCC)C]@>EA[
]9[a?\U;I)8:Gg3:20DZd)AB,a:Y?P^2-g0_d-C>X)AOJD@e#;O-U@XMW.b_._[7
DEE>=GR:#YL/a);D,eN[\R=X6KUaARWHN(60Q)<P;>CScIfXd:>VS\@)3XOX19a@
O]gU7a232C9EMF2XO]C#5VdIX66\.D&\)Wb7:0-D7eAG6GfKD&)3VeH82>;-LbL7
G91/U#LVAaT@.F>L=^59aET[,eMDQDU8#EI_7F;]>+N:RU,g(+X<B.f+G2=T37eY
.&&NYW\0K<#.^EC0)?F2WDS64OVP<]V>GWOIW-UVGDV,/NYaI[@P<Wd8\7E>=PQ:
dZVFY(8dbI[R/#Q\&E,AG?7.LUPa\3Jd.:T;RBOR,:W7R2@&e1&IXa)A_;5^J)BV
H?7WdbC,bDbQ;)#O))?-X5,@6YU9(eTXYZI=N/D6/G<C1KTLgeF=07,G4@/WD.f.
4/^.140Wf6<L)30@E62g,_OYTLe1:),W+PFdY[Ie+WOaF67MXE&gSfY@4QUO7M5+
J;SCS)\-B.8)UG9H(\O/M-<5E]GJ:c_<T^,:6MK/Mf@LNKXJdF+cBG(gVY.YV@bU
0ZGHEIN5G)7(-MeVG?>[9?(J/^I(C)X=G>/X29V61E8_+=IB6Q^Yd\E&(J36_5Q4
5XL3[d25(@XE/4aaFG2b-W,cGK31LXR7bU015bBA>f&UI1YP+@f9gf<g#NEaK-fB
LJ1gf4Og&(8da+;=ZX4)<Wa6YGEa8N:CNf4MTB,C-bA@LRYe(&dCa>MgHOLS]_8K
,<+1gR5c75bG\0,abRd<^J_5cf[g+.6:WX>>QCVC9:UW#Z\+U4_[g7LMGI-[Z]FW
G:16/DaBL7(?H,N.^^.Tf[IFP;@&)bDC1:JQ_/C-Rc4H;EaaENQR]1IVg-3KMNVc
aC+b-<+S>Xc^JPbVZC:-CZM-MI#L>#BKH_^4O]Y:9,WY=P:(+&GE;cb\^:[YW+0X
;eDJLY:.NE[-A-P+SW^&c=<Z9fc?OIe[DYO^0++9-CX7>AZL#=7]T?,ZR2V0XL#0
Z1<P+O^?^OV4HSPaa_gGP9.9Uc;/EG#\Y/<5T&a]9[D=ZN;Fc6PAY[XWXP7>;8\M
6ZEfe1=^6Z:UI@[Ne5BI8&LTTV0e>+E5+-DKYbMS,XKUc/,>[>F\cZ.-KBQOa2<F
;e/-]JKPF.5=96/Y6H(\2#G5]NB/3K6@#;/CO_I+Q=^#EL[<JIfFg/L,7:bKaQgZ
Z:-=_P]=#^LN[@0Dc4?L068+E6d_LB^0:a>.M&0&650?a_[R98?IdCF/_X2cJ,2\
>TWYY:<\gCY,e=]DJ,N_e[WQJcULLZ==AMJ@&@IQWe]4\RW;8[9/00.8/(UIa(GR
Le=)_NgIZQ_CeRS6YNWO9JQ2T5+A<\aH8eU1N4ZC-eYB5.#/D[16S:.dNW1X/=I#
(]7/b&]ecTTZg1;6/YZ9#\I?G,RT.-;M=1EgT]#c71;<1X/WFIK04G\<TXC437.:
(FH_=b62-bT;>^T>d,J::+EVg?<3KSePLVf?3\RE/UVW9;]PU>fNEc3FGS)aWQOK
92e7?I+IA,CHSFW3J6eWUIOOFB5=H+(.9b&87#Ee\9+GeXf<&Sa@Db>)K4GTP]3)
WV<05ZG\ed4)X;3S,H\W=&+37OMNMF69F/.RY/>cBV#a6Q--f^W_-KA?P906e582
608<(_812^FCTZFG0DJ8K,4QV9]GX3E463@P[f=EI+LB-9b7/D9cO2&A[WUYEc<[
&aZSf#eDJ<29-9#WI50WXH;UZ6(^=45O:)#;)UgHLO4<XYTLDaM\/W:_LF44)&S[
5?]&]RX8Yc1e=8^9(aQV)d)EJI,<,BKd20M^K#0-;?-9QZ-S+800IEcXZ#b9XJM4
Bf3KKgE39&<.=gceYJ^B=9/?fI<TQJ>[,[W5>+GJ2aI/T-@=?_>U7BGUKbcAQKP<
QE2LDZ9_NMDHg_@?JD86NKLH1LGZU]c21+Sd@d9\;gX#JfIEbPC#Yc?Z3/65g>G)
J\d7(LBSf8EZ7;&YK-TL0A4BOTC;Pf>7\W8DIQJAB\Zc15+d6]NMCb\X7bcbX6+@
EM)9D>;;SY@aN+)EeSaSJVY3ecK0ee1+WCNb=0I:8#eWW#@/RIKSMMbNN==4@P37
W#2]C978=K7P9(S/FC683WF(TB7SFd;\7E[FVb6_A[_ZJXM.0]727\-5?Hg;[]P]
?2cK23He_,:&CID2a=G)a0G2,c<P\=Qe7?7<[70-SOO?-dfb4#dB&:J0[#E(04E4
I<=gRDdcP]X=K7672cF^LY3E8C\#_=PS8)D44\FG<7M,/@X/6W:+KKSXg)?gS_\F
3Xda.#8Mb+=\[6KRJUITVL_GQD492B7.5B&SLVZ#-b<Q@BKP8;@;<5MYe.K@20]U
VV@7V4b7N]L,:A<?7JW8g&+QRd8/5L-KT_URXLa\W#?a@HM^=J_5)BWTJR_0cE^.
Sg:/^#H&F2f2W+BO3S;P0Y:7N\F9Ba<DLXNXVI1OI[A^X)QcM9M/W\Y4c?S]e=K#
/?gbL83<0)^B[8<5K[LOb2[ZTG@0IAF^O.5PJ_b-\gfER6M3XGJF6\+[EAgN4+D.
4I11SaAZP@0.F&Q9L?@3FW=,\01Z5>)0<T,D7,3<8X[d5Q(];G)X24RW&^bW74cU
\N>0aV^@[,9R#aFgSXGT_e@YDg=N[7,B]\bR:IEL8)Z6#>RfQ2;gOBa=+[YP#_-\
(E89FAMSVTccCa#<b_1gMb^f-L5aJ?0]>_9Z=S9gA=3/0Y(K9ZX>TS6Q32]KVKe6
Icc_Zc_68)6)LeS+;5)->>F2CQCU/0^8\&D,2W4gF\94c\J3C]Ydd5<Y)c/]1KE_
g:a#6Q.FNUMZ<GbGC\Bf)(ITDTVd&90TCQaQ(J4R:2A67Y^;<@g?geOb03&6BQdY
-HDM:GMU67ROB1G>?8cbg2/TeOAX(R??1Td@^)O?KV[:/B3RLC>9Wc12+/8[_Y?(
0?A@H]C8<KL&ARZ/^c3G)TG0-O#U=K6L=,\W3FU17SX>/CO=#5\MI@U^20OP+MT/
OCegDJbF_2;46.G:0gRcA2=^(d?UD,ZJ_01^CN;Mg/UE9Ba=98bVDVO+a1N^9&^_
b\;/VL;B\MJ;3@(K.1,J<1AY#1SaNMW4NL>RPRSMNQWW6F;,>OJCE;:V.Hc/d^\)
QWU;DXQTT25\g&1Q3S1C)4Y^g>ZaBC8;E?^5+CW6;>DMZLCZ+3CEI?3M6L5NcE81
T2RK,:LMJOSP+dO#-P]0&JXHWS1S5[7[Oa?,V/#<U\L3,76G7VbW;(KH?&EV:&M]
+0L4MW2f0KK1PR^^)L+,bQZ9fCgECT^AFYfY#Lc-JWJb?eXO@cKN1F,V=[D<?]/#
50LBD5B656\H.Y/7?,1+:eT9#cJC^--V&JU@c+O4;DH05bScLa9+Pb0SMEVR1b2J
[N=J7V-E]b:(K:ZR8IfLSXW.]RX>gMf>]QL(4?YUd+bc^,g^/9KM8HS^L90Y>.8>
(Ib_QL7)VD#PPP.?RM<ZNB=66-HY85bU>C9[D<Q)K61^.B:aY5H^?L+fJR0FZ(=L
K;[eEg,,51K+N7/9WNC5-HMaDH;Kg91,Gd4TA1XRJc&9;QJc9BN^WPF#B::3P4)c
C9?Fa8OZZW3#?LGHY)^Eb:AK2GRPYd?;Z44T0Q;>#F<D]W./;)<Mf_[W&]]>7VL&
,A3=ADX9\-B6].CK)PYe1=2G^&\T:c<+Y^5_bZ&\6eR7d3S<;?NK-dDOMXTHCWML
3(M.WA;9=P8&9=SA#GSMZD]UXgE8Z6]KfXVAIVWA+MHT[)\(#9dJRFL6I19]-fg[
B#3?<1?]cWDLf.W+;:S),Zf#NI^X5OD:NZ,6TQU5[BQg>_I7L<Z9gVHS[3U[eE>e
4)#1BN5?@:0Tb4_-H/Ab/_WTPRb4D<#WE0#SR:0WI;,EN\B[D;eX&f+a/1Q^JBZV
1IAeD(UMe+.&,1\[D8;)(^U7OK]cK:=5)G8UbJ+V#4SZ?&6E#UF@;W^gLc/^Q9\F
)_+7:AMWM=K(]KR?g4FbI,VV(_7a3-E8ZSdS\\a?2OE)^)?c/KC<BD,,=>J6PK+Z
:ZG6T&2]/.a_d:T\44\5KQeO18]a&W(bc#.KVF03b?BYSSW&[6^,fZ-gV(.SGH7K
OD[W38XRZ8C7E9RR#32WT7GF1;94Z4-cB=fGYA;I^[=9XcOe[O4e4b-5AK#5BM_?
b,O4.d#96(gBZLL7-XA8M<S/]EDBPb@R_K3J]423-C7[_aAOa,H+50,LZ,K_,E(;
^eG7J_70eS8G.-(S?+X0+aKd:Of+E0GAf/XP^IB=4c)OC-fNWY:4<bFbAL.+=AM6
Ge<g8MA+2U\b]g?Q^L);Sb1g((\40^VD;DX1]INZ40Q8U&D?EX5#G47((N;c(@c8
07eL_.TcYS3Z6HbZ@[3Z.V_T25b7[bGH3\>P]N7-\e-\DFOUXdGg+<33)M13eL)L
6Y8_#(.@VY=eE&H=RD+[0?Z_UCB:B?Ae(afAB5f5D-S[C59;_I[:88Y)TX]RKD21
g-a^LBVOSQS6X[bE-QG)GES;:J[8RG\DP^ROZa[5?2W5PGECY4H.6-T2+a((4HWd
E0-5E^W?IaK3<^U[\Mg)ROFK6RMQe;SCI6:_]ES[&cMK4E9__M0#D\BYHJ<T]2a_
&D)&0gg7P<1)TX>a>LI2g@/+)OM[DZ./#e5B:J>4(cbfQVI4NZWgK[Qbd0,32<#7
[_;8Ded3Ge+LX^)ae\<[9FE7JXW5+QbWOBP0=c)U-S3AA@V8IX/O0=:W9RP1^_N8
MB&,1PZ5=T=PJQ<Xf12[3;4X,XI8@7V<+E#>cKPXe4b/S/QP_B\\X[bR[]VDC?S6
N+.16#De(9YOOdB?]M.,9GOI/\B(1>@>.Q(S]M4BQG9-dQ15VS-Q-JB^D_RH?YY]
15M^/Fb<Z<3IBGX5C,F1\T>8D9C-@:;]:641N;.B1gDIWVOUbHdG7W4NTV^S\?IK
WXaAM)7\ZVXZ6Y,#g?Gc_4&dG3Q.84;c7,07M+2F2KQ_^b&\\cER?^cUa]fe&6[8
,]=(A//GFL@6/RfWga43=9H2BJM[//T6L,I[-0[:<gPQ?V3^Q8\_XQT:5SI>YB[Y
ND@c&@dP(b;&<41dAf(#D[O4C[E+F_4K7OG9;#0=2@HQ/8]Vbd]#Vc2-E-;Le2+P
H1C=\YbU^N+dRdO-5T@FSTJWX?O,9DR+SJXX0]8K7XNXYXfX^C7bQ0cHR=E_dQ#]
cO.\FJZ9I.Oa(aT;^6PcEeY8>\<9@666J?-9XAQ>NLA#<L?9_H)<1&X,f)bbUGCY
6@-7Z&UKd;)\7-aIc&]X@b6[B?BJZa)+bD.MC:B1c)IB(Oc^[3/;^B(:\39^LN5V
,T>cLJ?P0>H87WMe_@1eb&P2O#AA-Q+2Sa)3(<bWXS,4=FJEMV/:,),D05g(MFZQ
4N9M6fZ+BBRG\#TL,RIB3G6-eO5bdg]7H,<ge>@;;B+7H^((CWQ5IWSPgQOa(Ad^
R,e@YD5WP5Z24#L-39]P?R8dE>TLcQgZCCd0a.b6fEG?TI+U)7>/E/OE6Ra(1JRP
(O1KgQU>Q^.A5Ag6+a>A?NC5[AP&?e@C;\7_ba@TG?[F(&M=GcFbbb4ee7e,e4C:
0JUdX(bJQTLg0K2F=,@X^GD.#9F&Q_.XD/EGHQ9;MC09@KOeb2,L+M,Y5[+AYKa<
e_#F^;7/ZO&=9R7aWSKQ^QK2FAE3+a7Z8M\b;V4Z/0#RfAYA9-/&-G1M>60a2P;+
a\Bfbc#PK54H-4:K0ab5MQd38V^?M3&7&/4E@D,6>@C;-/]LS4L5,31&e1^CT_M,
F[aHO,LD11,0d38LD[aHC<@7\^/3/L6)48PNUI.<c\Ud1gY443[+[XUH>=ME)g]_
F.g1_\MWa.Hf,\S)L_Q7:L,Nf-E;b3BdXCe1#,<VbD/K@)_LQKU5UC5Z,[<?PXe.
=-TR-,Z>HVIY<67Z^4_=4QM;;25,<,:CU280ed?;8H_dQT1f)E8+7>SJH=_DJ6)=
LOE>aXA&g<4329L>g3D\dNc1LC44KSZF;7@_LF/N-(FS9=YBC9IJ0dA8/b>S+3WR
:Y=I06<T;C8Y+Y-A\8CE&JYIU0TaR(MJRQCD&UQRaK.[7-0A2dC_5#Yd]\eb>.O<
M\2BC6\R&DbJLJ#AJ,<0S-NWWP#</b64S;T/8V505_VQ@3XIIAO1BD:GS-9N^O,3
[U5,Ige8]AaBTAVGMAa_ZXId/KcS<V.UBD^eVdG^,7e+>,;VM?cd3Q^.)?Z=&4-O
eU(6>>&:cdIdIQMT=H0OLG[P;d9^dR9bN/]<266g>AU^e3=(9(K6&P.VQ/04eJ_<
K)^[BQ+RL;=ae9gQXGbQ_YZM8agFVeS]PI7(>JP8TTYVg=S:GCQUK+3f7<L<LAfe
N+XKQEIXfERQa0LXV]fX_Ff_.eA2G&ZVgI81QbBf,CANO_a/]eWcgGg&&\^F:J#?
0-f:c+/9<?VG5&OLgYV7#<&A9Z^WFL@Z?EBZ(9Q>2-S\][e>6UNFL0=Bb(e2>T?(
(RZ.&dZ_JaODePA@4X(SZWUd]A?VgXQXf-^[9_N^S&B2T/5K6b0bL?XKc616EP(3
3(#F.J^@-5;78EC(&^K[Y-L-]GO+;7R7Y1T]?LL(R:g)?OA/_W6^2V<Z6IL/W0MV
86<QP9Z7g>84<YM6DZVO,K,d.6JGNMG+)</d<V^M:&XbQ36=0JCBG].)f)g>_D(F
8f#Y^59YI(JB@Pag)M_F_N(c3&+.69L[5g.P<R^,[1g[VX()0]CfV\5.=@)BWDGc
DXYJ@YAPdTf5[[gM2LK@]O=;Ea+6YSGdU:-c,Dd-fg199//F=AK;<IgZZ7&IePJ,
7JGU739:U_678]YU+::Sg0@gA213[FV/Q4b44<53X<\d,&da>#A1V9TdM)0HfLIS
A9B5g]ZK_R418R(b?05:W65_D])OT>=@LaCbb7VJXUfaS.X_bI#Q2dF5UEGO^/Z7
.]]Xb3D7=PV]f2?E?O=>BTda=<,X.>9</bZ-e-dI^eM;)=E8C1c[PU<2FU[00]H\
V-_DA;D+.]UcgF[\bKS,VN:4>G7A@^7FP;B1@XD=YU3+;b15F1H;Ic&[a<cVfOLC
Z;&5/]\LG+^[TLY-d([=>gT5[c2Ve)FD(K:+Y2c(PT#g;[F?^?eI--^-DP21,/AX
3L>3R/WEbD2+Vf8^d(WX,8<H7-.c:d7Ce_b=g[YK#4VSX#6b:&N+a@SbDW(LP+g?
Q)-TYE2(+c/GDR2QEYTI.)=4_)=6:,b;+]+#=&;Xc&WP=_?NE:Sd73Y_K=OG8SeE
#>1Y^6T8afg-4bb=\[L<Ob62Y8Saa5JP4D6f1=PL;&P&O-cC;=)7IUO(c&GN+J[_
9P.^G@gN/4,:Me2Nb[+,T/<d3HFX@f+]NS^B@>Wb0(RJB0TLJARV1.@UG71=0G4I
]c#Ya(0SZAXF9\4&XYLB3\S0EC7R,QO<@>?RZ8Og9G&PWDNbQdBUf9E)7/]aLF7b
PTM4T=+FbD:],2A:)K?>-Ye6GX<LU_GV,IU2#B0_B8EV#1),Z,.6&Y4g8D/]Dc^Y
0+a9@>JAbPKgLGSK;&[I?=T?HQEK9aS.Va&4FMEcC-4>6MTW9K/6<G=NdNV#LINa
9gGQ^2M-?G?]-c^5E)+&=_6MFgIXbBHN2I;MbC41NF/XRNEe/;A\/T<3CD]\UTO/
[ZL.2M5ZPF<^HQ)E(&b2e,^O6C0fJVE>>GS9Y.:X>A@dW]8;OD31g&e9f7g)_-9,
:QPgHX(>gN.TU>C)0-L([M[D(T@-TODe^eeIJPeRg2@QB+#MP^W,_F^SJ)@9[21e
GNbIXFBc2Q,4P1Tg/B#I24V5:cYMST&8WFYY_6=TG6N_+@?OMQ(B)DQ-MI7.BY+Z
+gEM(4Y8BNE_-_M+?gJ;5L<S81<DcQZfeWA^7K.)MWWB9-1&f36#GLR_Aa([dV#>
UW[UeBV,>WO:KXYI.]B8OPb[U;N13.AfgbQ96dJ6E^&7GJ[\/B=@E^Hg=@OV@6(:
=9g(WC/Va9Z6daHUVDD,11[TZQ3<0T?=f5\:WH6^@U/fgY02[Z](H_a&7R)G_L4Y
?HCNUXZ=<.#b[N7US<UR5TI1CW6LVC&V#_JL)WS93@V?A<0?FX6IM8O@b:[X)N>1
&1YfUBFJbIE]gDGM?VOI53-/@ELHTPEdfKFYG-F[YW3AJ.O>:HRWZDA_\-H7ZR6Z
Y=OP]<OX8U+b7GM.:0d45=R)MKHTDPg)_1aSDdZ\>ZI>;)bb0RKe)+@#J1I-XZd8
H?J4R,[EUNc?9/XRaNcS(FfI0@ANA447#3_&32NdH5>R0bT<;Z.KX<86O\?Vc<Ff
dATM@,FPZNA:A0TI/2UJ7gC0X;LJ=eWDc;S+2><dFc2RA\HEIK:dgZU038P?8g1g
&<169,AVMVeTJ4U0(4;LK0MV1Eb(dVUgX4.Q(A;@]O]MONA6SCG\NeED^;O-EE;X
caOE>2eU_,UY?YB6;W9.508aBSWOgW+IH=R&ASWJ55@XRRLX7=90,K5e8Ve(E//[
2NO_<R1X4<9UHLfDAY0^-A.L]e6@6WATGe5VIZ3IecLBLOYECSa5JA0FC0bTH?YN
EY6>N;MLbL#Sa=<&Y:d72@[4B99UVCP#.]F[7\0#D=92FeI_J5=D5<6\9C,W_EaY
QUbJPK<L]:1-Q@#ZIRKFEM(>U2IBQ?;NW6S>(^?\;C?Uc_cD7PA#H7\T/P<aN&4+
G95A=T3)Y[PC93,f\DC3X6<Z(60ZU55(W;X]FR3<^b(Ef<DZfeAa(RMMG;5M>g_B
IS4:AQDR-#J#0NLRMQ-0C?1,SL2;CW>^ORPePf2d-KP0S66C.3D7WH]KWZH@1YR=
^M6U&V;<9Y&=]9XB)OAKGT,5]Z;Mc/WCA9[B]JALXe3X=QVHS+ZQa=P)/998#QON
YW9c.K^FP@);\2J_;C&KLPU8MH?&58&T4cg5J@,db<Ed3AG1R#&@NUQMF3#NU?3D
[>bA&+9,-8?/cgfSg?[.(=>4@)#bdg.Wd&O<-d[6=M17/#H,S8Q1S#R&cKQ8.^YA
bQc5-_fAH+eV,ZWa1<>ONVdYQM;5CAV7,a)0/U&HQ0O.f-\?@MGfcS+@QK#&U:KV
S/D)VPQOL8E^/9)YVF-+:-P_H;B-+CfITNDIKQ8J]<&51WXN<g[/-O#(\MXE_25g
d;BHN[FCH1QT#DSCO_-.Tcg&Xd-3^8B(5KPMJ&JbGI)&_-7)Y1b.TcgR6JKbJE+;
:H[I:>cgU;+;GHa:g4F<QT<f>K.WCE[4XDE.&QDDDV2^g_VT>1:6WWC0b>EbZ;F3
E+..??AVP0&S->Ud#2_]XOWW[<M@S_Z\K/M.M/<503+N0\>RPR;(1c,f).Cg^7<A
#ZdLPef<8JL(Kg9YReS,LJa:G<P]IQAe-J1(TJN8=8FQ&>b.JgE+FLW;V66Sf)6W
0c3SC/=<,KSUdQ<M1K5WP^_NKP)#]\3<8T@7,,c9^,.K9O@+bB94Pb_],Nc=V9/<
71F3f-f=#8=\KgbD>GCB]?cN#3+@P.#O/ECd9B49LZ7N.6V#BB_49V_?eXU#Uf,4
LJ)3ZT[O(e\4:YKAZ73/_Y]#+b[FMbe1S&6Q+,b,LJf(H.Q9;.TMTJMb)BZ(Zf;L
b/6U8@NCce3JEKH,DJN&EIRNeZ,F][JaGF41;DAERb,5Y=2.b?@>Pe&TcJ#fQ^(e
R6::4,_S@\9R&VDVD[[#.a&=+?44T3=X7fL6ND4)7b+[[XK]ABF/:CF2>?:+]]<\
9+/=^\-<8C^ZTfH]</&a^><EAUP+VH:f\bCSZLb&NHac?:OgN1J,QL#&I0&QDdA(
L\W)CaD4]5;cGT=OFX3CSX2S\:7;535Ka]@A=7O7Z2f,I338S=E4eLB]8&BQXd2T
@/UZNR4[P,-=9LQ]3)M]VE,R@#V@,@SZ,;;TF1De?b5eW&PIMA5;T/GMO#Vg1;cb
WW\,Q58K4aMW44IBg^.C_SH?NW/4[4]bB3-Y)D9L;J(.<NedeDF?NME3P+V<L/?,
Q5E-^R5\QUNaVd\<1;QHX<FIC6[4P4YH=Xg[T>WR-f;XKMfFGNYAf-A\f#V\\_5_
Q(5E&Qdc95+8\3G7&SOL902(b51][7B(LWJZJR=0LT8bMGL):]gMEC1E^3a=[9S?
#B7[-BD-G2.NH@f@_LV<c8/GY1>UfIZFLa__&fQ9:A^,:)BbG=(ZY<[F^f]6?+HW
L.HE^TWEA^B_-]O;<JD36NEGDgeKXR:<;KVa_Fb<DVIFP7D80Q?f5C=.(XA;&T-F
X-Hd3P]LeIH]1G07L62Z+UDfFRcFIK=H#\WHAWEM6?0\gWg;B#&IY@<M\=EU]agX
eRM;FLR0DOa&4.<RaR39C8>8CA.->EVUeTZ6]]_gQ2Pc^D3e>g/QV7a4=K?C]dG#
]eN])JK,QW=JQ#FK:_f5_DX=,>02Ha])c#IZQ4e5,,VI5dW^dAK1g+6]2HHKd4:F
B7CHCaO&dV?T+&,3ZE4#FNF)\=1((^H^RE2N&#>GbM->K<,cHf\QO2f.^[QEQM>-
W)VDaMbFBA\NaVMW^a>dJ=cHf+@0U=g#2//>&PG?0OJ@LDA0]?GLd<WgUWG28L00
J^M.P#FWMd-,MEW&U?V8Xc<EVC;1?a^HL0]_[QZ/#H\CYQ?T+BUYMKdcFbBN94)7
MT@>a9Ge_0-a//FbOc7OVfRdfTI[DQ5a4)<eY8Te,:f1<-BC?EH)Y:@(.R0d0.I-
M2(,]9#.<OGd<PWJ&75XPTMR?WZ/ga_2;Xg77(].bBU[V]B)TB#e45EMfKc@e@2O
<?95I3YW2D[3I[SJV@)<0(8&UZ?(d4?+/NbZA5I1:EHR#_=.U_]O3Z0\?U_AK<C6
JT-d.S_6S6fENIL?U4Z/[)/7-E>Rg,\K3R&GdGBf#-g(Pg8W_GFJ7b)e1IG(/GfJ
2)eg+9,HgR,Df.+P+E:CS4/M/cFX36[TfR(GIUO<=AZ72^5FOWS:K]RK,;HJ&OF,
Rda9VCN8SB.+D;^3\3V/(-2Yd&fS+HY?O+K38L;3W]5fC/ER7:KZg3EH)M3)eVE\
aA5:I@=DDDA5@8I[KKT<1^7G1f)9_7Z5)]2WGD]G]S@+d?I#UMGXL\O9K1Sfa,#@
G2MS)P6d6fZaN4YY_X,&6g3_81.>M#[A)WVg[XE;AOWXXEfJZW:b+TgK8Ib.U.5Z
+K1MDMgHC/OCUZecFU0:7IGG8\(.2./Ae:(NdUO0&EUDF+2)V[UCDf+>0GNG9EgI
GYO3cJ6ZR(gK<g&I#.ZOI9SW1)7>aOgQ8.+=USDPZ<C:VfAWF4V&74NN9.#OaME9
G>OL9OTGE>2L5T/JGTN/4;)e)d<F5<G?c0ZHFEL;5ZY+Y,SFEQGdf:=4SSKB_.UO
#)O8;YE:#3dV,&&02fX,AQ#2GF+VfB[S3U3T8\0E=6()f&UZ[ESX_^EcKJe.M/AA
W[T4:Y963a3J<ZP_D/8?YS;9:Y2WZ?]CFQ3;ZQPF4]1c6EZCBWK4,Y;G.Z7^L@-F
fWHF8b2F<MX?XgO2Yc+,WQd.b/b<V4/J-9HX9(FRd-X,<9D?WV]XE635c[7f^2aP
+O4YYK>\E>PTS91TH]6JI6H;UEXLNTfa/^L\DGf\J?R3YBJ\N8@[PM]E3#^OF=;Q
@2V[X7?-Za<QA9VI9b<e[5UV-S89b^F<gI@0KRCT(;XK=GAKVR0Y+&>]&&P6N]c.
DBUK>6fK?DS?P,6LN/N[7K4f.5CZ+eSac0DW7fPL9KE1NF2W.e_8RcXDbaV[eZIL
9KMYXP:HZNSO@S>D2SKWFZc:7gG#F4\-))V+C-L(Q7[55&d40<]BO5;=418g8>@<
L8>,_WJ-@[].B.6SB-&RR[K7W-1SD@+95>SeI0cY/]Ye,1;VGURTQ\0J\)aIN\8J
=QA93M;LIe-D9?UC9ZE5eC(+/<8Xd&W_&)Ifd2aa?EA6U4>V<L4UdUFN&RcSHfOE
:2<F3JRV=@I/;I1dY=^bOABB,?,#^10Q&(Q0EdFM+85TVIMeNBWcaITXGdVK^WWb
&?K39&A&\\04B7Q1,]J#1:1?cEa1=?IIA.M2@R9GTg)-Q9XK<BO4^[AXaC0f[FLV
T8C(d)db;a3gJFc;LVI8,\(RS:R;ZW?#2=S-_4Y#HG4d;R4[(JD-J>^#=N0>[HDV
NJ-H6G9W_gMe;=.6?##24O(S^)db^IV;CVb>#;E-<MOPPecLW945]1O]0D40dRRe
VUa):@7\Gc(\E@]QdCM,ca&:@\]E)RL?Q6:N2BS<I1aT@Zb49MK[G+2IJcNKZUJ=
BD>a0Wc\5aC\@7SE/INI5,3Y[d3BO;K#3DT717fB088^BZAc,N.D7@K.A1[La>=P
,Zg?3,GN+BGa<b&,I\EJIWH<J808N&1\=J@@EL#1IPC/+R84DZ5E9a:Xfc07D4db
LO4>-?\+f_Q942H,GJRBS#RGaQ@UMeae1ANV:/YL0FIO&FO>(WC9H0L93G#?BWBX
S7eUN_0a@9//EQb3]O)Z(]X2SHOKO3d<6cW/BQ\G6&Vb[9DC5;0KQW7VM@QMJdJE
fX:?a_E?IW6B>=-,5O#Of>f+g.?O/a<86Ia@+QG^5K6gRE]R74JSW/g9CZDc=.21
HQT\O/NB]ZeDXdaZ;KQO?077#T.f#L#RIV])>;-&egTd7U@2[8SN0SDP,=e<5_43
JfTVVMX-V3?^[_P?&RUN+IVbV/=Y<9G70=3_(P)7\EPWN23LIKT2Od@NDBXbYOQ0
Z).\ISRC1a9K]f-0P\aH)=HH[G2cY^76<8T2Z1W)0T-Kg1E-H3TOH3(0D,KP7\L6
.\KFFCXd_Sg5TgKVV@;DPHA;M9&5;6-G=Z]5a&Ga?81:K-J[bOc2ef6&6_1eJd+O
51L)SfD<^]Vb#Q+dT>KUICUTGgBaF-2_fD3P4=;DQ&]NFQIGf<e#aN1_Ta8dL,1O
KM:D?M91^EZ)6:KE@1R824#=FL8[=&c57G37)N&)\cZ7;?cA(KV<Gf/dUW9fJ:@)
e4&BdZDa?0cOIFGdFUH09Ubg6LUJIJ,J\0=9&bH7g6]d(0M^SY_GV0B-g2ER-T^Y
?2FZG?Db8c+ZN)XYK:MUIK?W,?>9#3_#068^D1CTDX(7/^Gf?O3cMU4NJ4Z5XN,b
QN[cZ>?4_H1_WdW\a?;F#UFPf(R/V79.=[,#3\Aa[AgV:.R5;:(gM@>WRMF>cJ@D
J0>&A;W0TcG:#XAG3;[[??9+C=/NMX<_,3e.4?NI^O?^)8:MD<F:[H:/QUYW?bON
J3JG<7U3VgFc6;]Wa9SL9-e7Z^^WT&Z=[O)&5P=,N.WabO(9\<OO>/]@[FcWcUKN
TU^O6,5Rc5T_5,82ZWOJ;??68?>APG3A.6;3E\PX^T?L.7>085Ja5>f&\#S0[V)&
PVcfUDNX;acY4[e0<0X?R<T]1ON-7\L83G<-W\[[2Z[M390)KXbd,NTcMb7Hc-51
0.0b@#PLd\.L2EM.0GeH05C+5-5[f&NaIH?IU2Vb97ISI;d\5WY)4Q)JZC^AIJCW
A+YH;[^R+ZDF2+.>.bDX/RHI1>2dV72=Sf=VF<gN87[P]/C6;a;NE3TS>aFAES(O
;?O3H8NJ8_Pbag8HaW^8f(:E=e&7CDL-W^f^0BLJET1g896GM<G)&L,OS-JF#MU7
R.CeJRR5=V:[L2;.-URf_Z.KX(<gB,/WCX\a5[=IVB4@OKdKUSPb6_\Ae[fN[X0_
:f#@(CeD#<c8@(?@PFV4)>d]F\;.gI.WFZ(Cd44@Zf(85RG-Z#eBF]TX03)H?8WL
.CU=S?#\=PN,^((+IW3Tb=R#G/>1/X[_d6DE8K8+D@^S>N-UNUS^(#L+R(OLCGTb
e1X5(1690F[UE&-)Y\[Z/DJ0_N.Haa>?^H?;H\IP9.RN]&D]4L3/E[dNG?NUVYO>
e,K\LN=)+\gZ=?95-f]]KR]TA,_<-@@Y<KX,LR4DLFNd,/0gS#bP8?TSTX<f8]Ga
J(9\9(80RJf4>\QYI,ed#X8f@M19UVHfTg)4:3VB[O8-./_N#?+656Y9V@H\aLP)
,B,..UVX7HN9<Qc&[4>0dC&H19(]UYLVCf3A?gQJ6^W9&J4TJ;gLNO,L,0G&97)N
IA.gJ9ZcC</B_I73dMQ#FA=@b6.DE3G,O.V/K2(:5R6JPW7&1W1)>#c/Z5.Ne)>V
@>>3FD5BT0QdI>cK)b(7_/fLM\[>b@I59.\6-TON&DJ]BE_+gF1Kc=SB//AW+QF,
^&)g6^7T4K<TSW,WaIBC=3SDcVCXU[1?&ZW\&KB9f9Z1,@?\LNbE\R:5BWHP]XBg
.CU<W0@De(ABTU[&A5b4C;R?/g,H#R5Pc).XW<863-?LFMC-)&5Y:Y6a@Q>CLF6.
7\S_TeIMS+W5dF3a@\\RSCaPB^F0)^<7R;W5W/Gc5-Ceb<,?Ug>ZDBNYS8D_3.J4
PW<XZ-?HE6<Eg/PNS,Pe\JS;BdYAXaMfD8AZB#H\S<f\1TGb8Jeg<9]09SH.ANS,
5RcM4-W(_4C(b8HUD]0:f1FC&;<g?<D7HU5(4U[XP/PW^:Rf#3YRGNgXg5-9UeU0
#@HND0J-L6[K)]@E0UC2:@M;G;/0FFA60?bbG1AeYC]F=CF/E2C8PI+)82&J=+BW
8F9EH6\SY=;F8[(R^H^R=@\dYK=A3KdAX@.C;B3.]BJdHB/\\@M7190@JP:_fMg5
gB^#OU.f=QK^[:WWMEF,\O_eNT)g65VcBLZ(cIP4_97D7^V^<6=IX1=)^LFC(HK[
,8?/3D-HZDY=FW-=6#I]?B,14,PAO28gM9GM9MPV:UY6NFF,&6ZXRI(JZ:A@a&dI
ZM3X4ED93,UebI>=[F-W-@L@FNaW&3EWYbF[BT3Y6Cc@e458UBLg(EX;6>0SD2(A
VARJO0^?>?_-E#3H.gCOOCI]?fXVJ6J.CQD2/b(YId,H4K@f-VZd]#Pf(:]-)82.
($
`endprotected

`protected
@YV5KXP+82d\FPaWI#N&X;J.c=XgIFIF\V(UM)7&_BJ4G8WB\57d/)abPIYHcK-)
:dD@P&GZL4Kf09L7W(0W-(.fc8=]:#\:[.eJ=d19+1)fd-;d5eg2/&abM$
`endprotected
          
//vcs_lic_vip_protect
  `protected
O.C2e:E/cg&8>ZOGV\))e(9I;99Z99+S#2LE8R0I0S5=KIP4C4DV0(5gMC)gQC)9
eR2g;Pd_B?Lb.Wb-WfgH)f#48T&(29/QF:c+FP\fff4Y=G)V5RQB3BUSZAYC,@V^
(0<A(C+f7X=eK/aQE&2M[-:b1OdG[2>B)@)Kb9IEJ>?7INK3:M?BL4W/DS_;&)V6
5BA2CA?WPNd^\Q.DTP?WeYfde>?[BF25OK@TaTGB;I65(8XL\L:\E_&c?HQ)8:&S
d3Z\S5f7U7)Gf)IH_H,H+bA_N+,1)AQ.;-_WPf:aPYDY3Q=WD.LFMPO<T)#9)gRe
cR9[ESAcP.PAPS3/87Q[M.@a,@]Yg;+&Z?dH\GH].Oe;BC_AFMf:g&2&WB_WLEOH
Mg6c>MC_MX/72,g9/7(Fb8GZ#@_4/<RIRNIK;0S9/76<T3XeQ(PAWN?]c,N_FgQN
BVNP@AeE5Y1^=G7X+K]b[8#f9gRS=)\g9K7X+If#U,a+VB7CA]F1[[NO2#=KDUYD
McgS_VPfD+T]Kc(A:H+-#LEO(2NRH/5N&2;bJ<^gA7CLY=+ARE1DW/@>SU9R+cJC
V&1S:35#e:3CQ_Y5SD008S,Jg:C,-VgPE8<A@2OUKP4[3IJ^XT4GDO:2,[fS?/9V
_OYUEIR];5a)#&F+^6>+cV([V50MV1YL3Y/cX@b-,0c+9RL8J8J;@47GR-0.@TC.
C+W.H=Aaa_VPeJ]U@/RTJbg_)9^Ic];Ma;L1d/fdF_abNGSK[7B?3J49A=4B,G0F
TAI-6,=b;5Z^0CI+G1c;d8H23+9P\V>)[@@I:\VJ?S#aFIL@2#>b?e><:)SN7=&D
[#)S/YI#@Yd4.KffVD7b/[QaLA.)e\L\H9LU9[34KCQ^D1MS=FDSd>U?Y<MB9&;S
_=;\SOa8CgG=GcRMd?4HedII(&NR6V29<=/GH/=Z2R.f+<,Tb>N/(.H0--Bfa7\9
MX8:>;PbZCW,dSQJ@36^OI@,FT\7W4ENQ\1M_7,W&WC1](U;V0Y)4C]ZF^A4/X[0
+b02WXUZ\6NYZAY^-gQGE/2Z\ZXA6S>QAAafF&b_O2G:TdbYa8@,-NP2K9MN4,4_
W,4b/DBSE2B^3b-)fDY_f6^TVYQM4&1H[(c@-0;>F=KV=Z?g<+7cfV=ISGYaUB^>
A&a1^3ED0aUdJb))E6J8.MdSGLUSKUeXaX;7^]<2J(G#<]XY(0B[&DdTF+&^=c(4
PQ2@_g4cJV^3BJ),8[D[QQ+)FfHC(IU+GBY0]A]V4@3G)g+2XTH;5;RYTAP-g.9@
#3GS<g)YfQ[T#ZAD1NK8KAF+bF@&5@&#[N^J8\1C_STF\LW+dUJ4[2QPQ/V@B85Q
388K[cEFO?b.]0:ISO^DISA:]K+/UZ-7)ZC2BU6>3<AAAA;.@\G0.6H/9cDI>-&c
@Jf]/e7^gF1C6S1KE@FY#MBF]E&_FG7VNMOHgCR=f3,7CMLDQ]YN/&G,N?[d&?Q<
e)?,+HJ\ZXEO_/c-<)&J6>Mf8LUCKIUR[T-B8X^]ZPMD<]dM^)1UH^/854?g@N/(
a_2FQTUZ?:.MA1&_&3EL3J/<B]22G](_[&PY-L+1,?TOFP(5G;Q_IVg^CQ,=.V[.
_HfJDKbC<YRT0-[QIgAQO0LdC7Jd>V?B>I0LDPgc7fDO&EQALC^_eE1;P[4LAP5\
W)g(5[HQ#g_R,V:cYU4be62d,AU/;=d23M^cOSe5;P7a#97[FaEbgV],9:6XB9-g
d0]^GN5fR+S:MGdJTQ+g7S=,O#0./b6>13?7(QX;<0cU^Z(5b]K;:OO9^FC=cZ&3
4T>0LF?8H&8A)<8&E,Y<)5Q_W3=92JH.(/4dd>=]L#]?@C=4G=Z-_5#TL<+I&=IG
YZSdQRSQ>Md,)If-XB0APK<4H>)4ILNIT2ZB=Q)ONZ<^<^GC-[FK>3D7aNC,=HW5
NOPE-Tc]66YK/Z)gEg2WAfL[9P)M2PT..6(f]_;2XO<G9Z3>)4YVB<L?]a@/gN=,
AO\013@4WDFQHY8JQC0;[ECKf)Fe(O+(Q\QJBb95YYc++R<5])g(&LfaFU,f\eYe
N.0[\4(6D6,5,U#H8^F@R_K;:YDO7H&cCOF?dFRg)Ha-:b5_K0.DDg-WCYJ2I);<
_,G+#NI,V.?dAR?0DWbF4@Z@7V,^O[e1Wc?1VGGT,VfQAJNYLE-]@.f]+[D;0b.D
W@R_0M<Y,d2(<T)WR/1H18Q<d^+^U\1.&BfXP3):>W_)S&FY4DN;#M[+S<BJ@/[L
S9-9(6dHM2/-CQa6QA(+6R6X><\OT)V]RZgJ?55_TLD]4E?>C7(-^]P:dZ=N<I)(
40D<ZC?^1CV]YS206&\eNW;NQ#F14TJ,_^?+e9:0Z<cBFg?W))<BTGNGTAfZ)\YM
gZL2565?&dDD,W[g6b:8=/FA30<5LYcY??3?]/BR>Dg4dZ=O_GSU8[E4TRT0KcIQ
?Y9QVEJID>2^T?;VY0M<JJK>D].^ZHB]aKb0RZ:#Eg@e=FLGUW&9MZH3K.FPfLJ0
2&/,@9cDc90HNWAVQA?ZaMceT^\D>.T;ZQCME+CWN(0dC1,1;M-8M_Yb5)4[<HK#
^1TNT@JIJ9#Z)dVK&S/#32,#TM>f0BO=MZ(f&c@W4dFVHL352dA[[LHKRg)(EG,]
c=CV\K:F?7:N=OH2/8:ZWN786\K-Q;>F]/L>;86BcUZXLUV@ZIT#0@MV)1D)1Aa4
>[ZgRS]N&Of8CHE:-:X6&S@46gJYZ6[d1K6cg:HS,&:RR.f-F&TIAIMV:E:4K.D2
@Q:(_3f0+T]^6+=MQdA+C+(DC()gf3RPM1KS4(WQ5P=Td8D.?e&QQ:T@<Z3KIS\W
])>(dc0ES@+KKB#5GdaTeb-&5Wf:/<FJ3TE)P2ZF;_9XZA.K]HD33d6c\X4UVF76
OGAL80J1/WK((R^;,M^#(^64JTdZEEXW-54/U>Me#Ja?<5DaZNbS#60;2Ze)R\0T
S5L3SH@;[]?95R7X[a1;@S3?PY:Y9(>\?9]/G)GEf)A0YJ9#7HD+@#(R:JICFZAW
Mg]CAAD24-8g=/MB5J=;.+.N5#ZRJ:H5[aZO/_D]@ILd(GH-GU5EIZ<LG^:eVa1[
YS&SB0.Y]7cb]M(]cbac>&)1PJFd/40_a61I(_(PcdH^4-)dT.[g-KE@Y_EdJE?W
I0S5];:PXOJRcC_8OF)_0U&WcRZJ@aeMMXTLLeG@6TCaE)9G_7NY3A.,X.4MM/gJ
U62-K&D9)603]365NO0\F<@/NCGI0OU[(OQ?\.5S.O3b\CQL)ZF=g&#ASAf_@dQ-
5F1B#GbCNCLB+(N=\)-b;^+Pg7N>GDQ^0?8cFa1-U&X>VfWL:RB1)0?VXK<#0#TG
G2]MJPDDDHBVWJ6GbUX5_K_#>b&4Ogb#R0?Y8;K.W/7M\V_]AL8SX?gJ9dSfF://
\)N.]#M@[+E+T&5GV-/VYbO7(5KW5F^\PcJfEI<&,TR=PM9;(\(?^?e[(e5>Bd=;
0Y^4Z-^=OHbG0/_TSCXVJb?OP6J\EB90FPe<<FE5+?)0d\XgHH+D90CH0T;f)8(#
OP.CC(@bNgb^NOFC+5.A6aW<HfA\8,M5GQFAg9B0R@&/]]1JS7GdI?d526&#42U?
N&BS1WDUDT.O@,;=\2;B<0TBcK-9E;8=R0aC.eQ?#[NG@NGOGMCS\TH:0H:#1B6N
eB#HG-a2W#d[0UHfLO:UI8T4g)_D9Wg1cOP,0JdAI&b_0MUD3&^NK>33N.W8HIXY
=1gF/AeW\6Q9W+LM^BTb;^M;V>.ARZDRIXG:S/f/g;02/@VOJ&;WR3M+[;QTEg38
4T-L0cJIg-HPTSBH-+VeTZ#.C^aKWBE@+N5A#5J&ddO>?;0<DaYS0R5+CA^JIT>7
b7a;MP_LFE)9GgUWc/XSUVN6HD,\W@b+bSSe&2,a#X[c:I;M(_9M:+UOO9:A0\bB
I6[L6WEV[AZ2.gW9>]RDLQf,FQ=;cY)PF\(U_d9L&Mc<@.8NOY0fAI(29.(J-@<Q
T=V2&Z0\T[LaSFKgS?XGSGU8GaSBR0\K,]Q)R([[F7+cNUP0B4>?F]@eZ][f(S^0
ae5(Hg(5VK55T>#[(,L47L&]3Q8Y)F.=,O:DRdEXf5WNU^HR<0VFDELTE+4S;TII
<&_.@<Q->)d5EE-=_+N0U0&-T]_NeC<NgRU:7\:8AX1D/-d@+/Ia9f]gfSE&YNX0
C&4/eOSL^5^2cNe+Pe@LES9D:TPO;[LLGee8-6#](Q^+cS30L:PSD=e0EbTbb.]9
]019Q^UVM;P.PYg)?D_=TT@E?&+L:Ng:eefX,Y@(9ZNET;(EY.Rf.b/^-&YWc#W2
5[-W2;[_OVb)6+,eV.W=#O3dJ4G28Z3b.dc&</Ne5L:ED$
`endprotected


// =============================================================================

`endif // GUARD_SVT_AHB_MASTER_ACTIVE_COMMON_SV

