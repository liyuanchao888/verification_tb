
`ifdef CCI400_CHECKS_ENABLED

`ifndef GUARD_SVT_AXI_CCI400_VIP_CFG_SV
`define GUARD_SVT_AXI_CCI400_VIP_CFG_SV

//`include "svt_axi_defines.svi"
`include "svt_axi_cci400_vip_defines.svi"

/**
    System configuration class contains configuration information which is
    applicable across the entire AXI system. User can specify the system level
    configuration parameters through this class. User needs to provide the
    system configuration to the system subenv from the environment or the
    testcase. The system configuration mainly specifies: 
    - number of master & slave components in the system component
    - port configurations for master and slave components
    - virtual top level AXI interface 
    - address map 
    - timeout values
    .
 
  */
class svt_axi_cci400_vip_cfg extends svt_configuration;

`ifndef __SVDOC__
  typedef virtual svt_axi_cci400_config_if AXI_CCI400_CFG_IF;
`ifdef SVT_AXI_SVC_SINGLE_INTERFACE
  typedef virtual svt_axi_port_if        AXI_MASTER_IF;
  typedef virtual svt_axi_port_if        AXI_SLAVE_IF;
`else
  typedef virtual svt_axi_master_if        AXI_MASTER_IF;
  typedef virtual svt_axi_slave_if         AXI_SLAVE_IF;
`endif
`endif

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************


  // ****************************************************************************
  // Public Data
  // ****************************************************************************

   // Reset time Configuration Signals
   bit[4:0]   QOSOVERRIDE         ;// QOSOVERRIDE;
   bit[2:0]   BUFFERABLEOVERRIDE  ;// BUFFERABLEOVERRIDE;
   bit[2:0]   BARRIERTERMINATE    ;// BARRIERTERMINATE;
   bit[2:0]   BROADCASTCACHEMAINT ;// BROADCASTCACHEMAINT;
   bit[39:15] PERIPHBASE          ;// PERIPHBASE;
   bit[3:0]   ECOREVNUM           ;// ECOREVNUM;
   int        num_cycles_of_no_activity_after_reset = 3;

   // Common Control Registers
   bit[31:0] CCI400_REG_Control_Override	;
   bit[31:0] CCI400_REG_Speculation_Control	;
   bit[31:0] CCI400_REG_Secure_Access	        ;
   bit[31:0] CCI400_REG_Status       	        ;
   bit[31:0] CCI400_REG_Imprecise       	;
   bit[31:0] CCI400_REG_PerfMon_Control	        ;

   // Peripheral ID Registers;
   bit[31:0] CCI400_REG_Peripheral_ID0 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID1 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID2 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID3 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID4 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID5 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID6 	        ;
   bit[31:0] CCI400_REG_Peripheral_ID7 	        ;

   // Component ID Registers;
   bit[31:0] CCI400_REG_Component_ID0 	        ;
   bit[31:0] CCI400_REG_Component_ID1 	        ;
   bit[31:0] CCI400_REG_Component_ID2 	        ;
   bit[31:0] CCI400_REG_Component_ID3 	        ;

   // Slave Interface 0 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s0	;
   bit[31:0] CCI400_REG_Shareable_Override_s0	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s0  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s0  ;
   bit[31:0] CCI400_REG_QoS_Control_s0          ;
   bit[31:0] CCI400_REG_Max_OT_s0               ;
   bit[31:0] CCI400_REG_Target_Latency_s0       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s0   ;
   bit[31:0] CCI400_REG_QoS_Range_s0            ;

   // Slave Interface 1 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s1	;
   bit[31:0] CCI400_REG_Shareable_Override_s1	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s1  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s1  ;
   bit[31:0] CCI400_REG_QoS_Control_s1          ;
   bit[31:0] CCI400_REG_Max_OT_s1               ;
   bit[31:0] CCI400_REG_Target_Latency_s1       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s1   ;
   bit[31:0] CCI400_REG_QoS_Range_s1            ;

   // Slave Interface 2 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s2	;
   bit[31:0] CCI400_REG_Shareable_Override_s2	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s2  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s2  ;
   bit[31:0] CCI400_REG_QoS_Control_s2          ;
   bit[31:0] CCI400_REG_Max_OT_s2               ;
   bit[31:0] CCI400_REG_Target_Latency_s2       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s2   ;
   bit[31:0] CCI400_REG_QoS_Range_s2            ;

   // Slave Interface 3 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s3	;
   bit[31:0] CCI400_REG_Shareable_Override_s3	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s3  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s3  ;
   bit[31:0] CCI400_REG_QoS_Control_s3          ;
   bit[31:0] CCI400_REG_Max_OT_s3               ;
   bit[31:0] CCI400_REG_Target_Latency_s3       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s3   ;
   bit[31:0] CCI400_REG_QoS_Range_s3            ;

   // Slave Interface 4 Registers;
   bit[31:0] CCI400_REG_Snoop_Control_s4	;
   bit[31:0] CCI400_REG_Shareable_Override_s4	;
   bit[31:0] CCI400_REG_RdChnl_QoS_Override_s4  ;
   bit[31:0] CCI400_REG_WrChnl_QoS_Override_s4  ;
   bit[31:0] CCI400_REG_QoS_Control_s4          ;
   bit[31:0] CCI400_REG_Max_OT_s4               ;
   bit[31:0] CCI400_REG_Target_Latency_s4       ;
   bit[31:0] CCI400_REG_Latency_Regulation_s4   ;
   bit[31:0] CCI400_REG_QoS_Range_s4            ;


   // Cycle Counters;
   bit[31:0] CCI400_REG_Cycle_Counter	        ;
   bit[31:0] CCI400_REG_Cycle_Control	        ;
   bit[31:0] CCI400_REG_Cycle_Overflow	        ;

   // Performance Counter Registers ;
   bit[31:0] CCI400_REG_Event_Sel_pc0	        ;
   bit[31:0] CCI400_REG_Event_Count_pc0	        ;
   bit[31:0] CCI400_REG_Event_Control_pc0	;
   bit[31:0] CCI400_REG_Event_Overflow_pc0	;
   bit[31:0] CCI400_REG_Event_Sel_pc1	        ;
   bit[31:0] CCI400_REG_Event_Count_pc1	        ;
   bit[31:0] CCI400_REG_Event_Control_pc1	;
   bit[31:0] CCI400_REG_Event_Overflow_pc1	;
   bit[31:0] CCI400_REG_Event_Sel_pc2	        ;
   bit[31:0] CCI400_REG_Event_Count_pc2	        ;
   bit[31:0] CCI400_REG_Event_Control_pc2	;
   bit[31:0] CCI400_REG_Event_Overflow_pc2	;
   bit[31:0] CCI400_REG_Event_Sel_pc3	        ;
   bit[31:0] CCI400_REG_Event_Count_pc3	        ;
   bit[31:0] CCI400_REG_Event_Control_pc3	;
   bit[31:0] CCI400_REG_Event_Overflow_pc3	;


  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
TZ/s9c6W01roliQVzckuAIrBTRE0vcLCw/Ukw009oTX/NWA4B6FlANVMNDNoaZuA
Jeub+M7LlCAV+Dk1PY6RQoubmHtEtmdmMMscSqFAbrX5gqX4iU0AOhuysh1JGCyz
vM0WGUXul5MqhOlCGnINcczrmZIFss5EtYuWzR/XbkslMEbm527XEA==
//pragma protect end_key_block
//pragma protect digest_block
kEaOvNWXRvJd6sojG+KK2wev118=
//pragma protect end_digest_block
//pragma protect data_block
gisHHzPTrHgRAYQNais9CPpnpUEuKEJXASl7Z/hcMCzfOuCDqHfcjYno+j8sfXSO
AyOM56X98j9mSVYnHjx8n9YC0AmvhBiS0Kz673KlSAggHa6V7Vxz9HIvmuD6+Pln
fi614QI3RtoDgJmigNKogccwEGQvG58mtoa1oXpLipVhQqbidkFqt5tREEEcZDsK
H4QfXIS0vFG9dEgTT9rtV8DlaYi1upq6zMXC2tClw2mf9zgsWScXFOS+nuHmyg7P
njKao6UZsnUqo/Ad2FmZvLZd2HYyT51WjAYm1xwIpXY0MjA2WKgSf/cWGuPC2oX/
2UZcogzYh7WeNO/BRNRu381DkMrHwKrBxIIgwCs9N4j57p0s5c5MHRhOvh7NYBgt
XKb9HgdnYMzk/tBCBKYq6XovQPcPqCnBJ63+bPOmdMv2Djnz1MDI6cli5OhnNwD3
j6bQlHcdpqT0/hyhnyXnWKvhoJKkVdKd+I1c+QODRSAydFRY9BLH1eaFwjlF2WNc
UL1xOw5O6wGNrS05e5HftynWF+D3A//dLQ0smOgssFEz5NU+fAYcdiGyxru+triY
WHC/R4j767Tjafjtn5M9APY4mB80z8p18N5XpO1KL2xbTcZm+moDeT1y8kxSIJjh
hvAP8sxuWVYcTN+dJ31VoKZXMYVz7jz97pirM8HJuzfDf0ghc7+UCw4Ngug2SsSW
iru9eDIn8spLdxPgwnjOJcolSpggrqqFa+HgI3R+8S50Ox6ebnFf+rdF8xIS0dvH
W5pxFjTyixssOiku6hPyeSAuF73n8fxZYMxPxiZm72IbOCqxUxHS3kwIYpZba/e5
gsjqdTfvdPzct0d5YMlFX1f8X91uCsn/RXALCOvxsTVksOpZR9DwGJtQRoTVrEeT
Lqz07Sgjt7hW++ikkLzwsc7rFnv1ZS2PETDaAuJQlEhX9VVi+h7FT3KUpxz55yrA
Ua8g2hlaNR4OVbij0Ho/lTK0YFcwvJFbIWgVr36UMd5ePSiFrZoJNwo90bH6XmRW
UI6E2KqRqWmq2BH9IFC12UzfrmySWbKUp22Ruf9jCKW6H9ZOIk+b8A+IP5GvJaub
ncL/gRXx+3Dzg/uA69+BGef/YkCVi4KJXUx+VrbzTtF87e28DVYd5pbhHSwu7Wul
TKa7iUoc6KVEfSer0jEHN2SP6zOrymiY2bgcFnS7M+FN/iPowp0JrYAM9It+AcCz
4qY9oxHP20Pwjq6nD6PMucTMCOWZUh9MN/TwktwXtUx3H8mFzGRGSANqMc50sPC5
MRO7SpxUD/TO9wvA8v/UKOJSByAX7ja+RQUPDovlwioXQmpGLqF8XhmYMFyJljQG
ZWuZ1hlPHrsgJVvxNOsh61aMcxAJ2eCFGX9mO230HeeDC7oKukjyKYxcoFH45/lJ
Kw64P84mx1mCjYktTHoTvGX0jXkA/YJj3jk+djDjzTW6o4kgnoO04jXtGdkmESpe
GPWcX6Uf8WUGYIvIpiT405dPp+dgDfWVbnYM5JsDqsGtZ4g6xASTujzJroSkGUW/
VPkDD5rAKcUDDEmMxxJ0V6saTtQ4VtWGuC1NLEnFPfcofjBNVA7nJv3N/Hftr5Iy
htgLhB/aMohApzHBwUQz2C2MScJi24NF4utdldmNfAErOl5Q8p0pKXaNoq6SUpzL
Suhak1lTi5zbzTl8NHIGdNdRO8WXUzaPvESXTnTbeA92Iq2OFpfb5GdybsJBvZ82
zKCIyu0FGmu7MidOSdc/cOrNZFUHgZcsBDQ8PBwOMzR9iYfYlcn34JwTNlOFonyU
r5/hO87szLfkaNueD7pwPk0yOY4VBB3xJlCukBOd6d1u24kO76tgoTQE5BaEjk6t
JGVWGQv+7coRFQ5NwIoR51rZaMVIczGHEFS9YlFF81Lz+fEbC4eIW4klDkzKSst8
d1LadlSHat4yH3/xQawxS9A8LNxOaZDFumX1OgErQimkjnjUqdQqm5QXe8c44ouT
JrVmbqEt6a4bDuSn7+UvsR6+RWgRCu+TvKNf4iQaDdBHuJ2oMTIipsVsMl+Et0bv
Hu6yaCSxeGqXmya5bKnbPzHRVBFDqD33lFs//kiSU1zbps9g8nAOQjjS722VFoTD
q4hag0jsz85zmIFBWI78TZYjM14sL/Df7Iks+nEaP0Rnirx14GOxU7VUPe4mCT2H
+4MID6k6JZumY7ERujqt/pUaClS3EPft0PIak5PAIiQHPjWwIkbYJyDq8I/+PKbh
k3uDiySc1v0Hk5m5udveKq+jv+imvKRTXiN84Y4txM8qt9ty4J3y8dHN9ZO9b/Ly
wFq5SiqZ/AU8H53WNkvJFkHj0M642U9aa0ktuWuyROtihemnzhfjHQmyGZSkvFg4
qCMuZZI5vdyqmr/NXHwTDZDTS6+doMy6f1QWnTh1vPv/ox9SEFIU8+9VoQyIt0zb
PUAJ8QBJgnEWutCR3b5lb9QTJwwc92nzYASXn3RSXzHwnLjqGPeSEKGagWtTxelS
72HTlvWiNKOluoyYL9KpJZW+p2wrWHZgZ1w0377+cWgVXxI671OpbFTjgjwQOGgO
3VGHMHJnGG3VPWKhE3dM6RyR3jvp/wxtJpb82qYzk1Pr8M+gWsfXEXDF7Z5PCMy3
casZWNNEtRyQzV7DxnlN81NMDXoRam9DagvFKN8Z1/LrugBHtVsfnbCGfaLC/bCp
l+zBOKkr4GuQEvaOhE0t7yCphmlP4GbKgUvzUKiFejVzhJeCgt6ZtPMh8TowzHde
aW62b9DtZGjLUKrTQrWn3idX8zwnPwKAIo4tDAfZ+HJP3cEko860xOYYBFSbrg3e
y94QohzWxLcKnaxJWEAKJdWrc4SDjg4oKKQZ1TJLq4uRhpChGEbjYJjiPfLcgpQG
mSBRxVhYhnzda+tkZo+Y5IyKw+KDn5L/CFuiDcJsCAiWUdzA/FeZBqXS76Pyi3gw
eOh6dIqcHC3M9j3OfQ1wQsVFcK4PFyJUOSqymmNNWV33rPk31gL4TnApfRqkEys0
OURqhmArNhcfb8uwhhqBI5qo4Arw0A9REtD751YxjTc696iq8qKOsx6L1q3m0xMV
/Ciq+kMICZywyCumZi4sIhA3MO/GtSvuoD6ABgrpv+0JbPQQkQveoiWoMBMNZOM8
lNPkXncsUheki/Pwhh5gObyUCdFd0DkB4A/vIcOPhCvLvEXBR0gCfer0064GyTA1
9hpGZp7RNi09Brw7aXRm4FwrC6zzxnXZgOjxjl18kPnacQwQ2YSHT7VRcOTMKQQe
5XrWhlb9fzPv4+82KZFEyE1MN2HQiAg/eFXR3q1JFNxv4g2CDYVeA6Ia8c1/hHFU
oUw2w6UGQqMt4S0AlQPFUTSnvajtYJpkBNtpNklE7W60roArqkCtwr2Q3q5Fn7nf
PnJN2RsBysD89IRZ8fibcWWBKWgBFLPs6ynSJduufLVWd1lX1psIFg646lJhKDYZ
DJWnUKDpMlAQN+Ua0UdiTFEmg6NYoU/FgKIzaghSRaAgXDb1V5nSJDYuSLgCT7Lk
8jCLfiDvJ8AAgbR5/Ek6Ly6nRSxtVrDS7+5mvo1B62/4gOxzXnQpNzb2vQKzhbcI
FpB6SuszDsWrrF+WtjndUZDWCNIdaLzDt5duNhJVmOtiu7qXbZcYhV5+T22/nNMb
gttBRCji/PQ1P8SHVWMXMXNJmo5oq+W+1y49QG41dqyJR+Gt/niIMAlo8J5Z8grd
yNsUWE5ltMTezaF0W6WlhOEgDGAJmPq/5qGvWPAcdhP5hd3pm5IG8HsqqKMNG/er
qm8b6ZVpAv7o+/kATvyHp+tcMXUNyoee6DUT95u7oLAT/CZsplaJZcITB7f3L3Fp
fXZTNH6X6ScgM4r1co8SAtoMVVsNlKnOxqvZDEX5Q/BkbgTZpOQTDSr5AQKeeLvP
Hj+sj9ZNSkgClzKnOy3QusohKUaxQoZvKi7zYfs9Tf9hPMGXQfyhL2ocaIkTj7wh
TMaBLqm7Z/YHtGjVDxcvNR33vThaV7Vcjz3b/8aX30/999LVHdj/1mSTVYKLsIwO
JESqMrBeWWZ5mluCbo3k8nGpBRjK3y592uCsEnf6kcZJg/jkhBnBLwLxQ7yKgvr8
e9vIT37aFEWQz72GwegXYNSpP04Zyn++8g5Df6ZYGyj1kH6YiT56/9UC+2q6iX1G
Ski6hrIqDIu81cYdWVXDgYrlQyQZKjyf3Fv0iVLzyyM0i8yk1ksRJjiC421mAWqe
PLuzLnQKRbKjaaragPWaCTNgdM2waeUDUx8dUTxgNvqYoqVhh1EnPmyzUsq1xA/o
3vauscyuTdpzLSGnWBOgr/4/ITtNqpCtjJ4tB7L3FVYs4dqrp0Z9nGtIsxXb/vf3
3Ly9LQTY0vWBsxSMDCgILpBaAoNKGvzYCvgTfm4wfTnRMNW1Z+c23++dvtaqLwpi
YxP6k4bl6XpIQv1ICPPwOEDMtSrVBFh5KWt1YqFApZbCLTGZP9norxjSbry4sU6f
zhiCmH+bLW5GPTDWYQ1SEeY55GpKKP7InlKUvmhvZ6SnAwV9y0Wl2X5NidxFNvHU
DT9spWpJ2yxM+eMarVCzgS/kGscmogKiQwLle+iO6/ss0tLx02v3TG5M6fNIJddH
/HBC2YeOwJkfdHrYXm5hctK2/vvDpG+uTZfaEtYB1l4VDaLmMajMilnw1J0ABAAl
fJiRDr1wC0n4xbIKMi36zdZafc0snPeF5k3fhVGpvk1k0L/Uyty7mEPk/jwKyCuJ
16vb0eWK7QzDYLclDtfjuvPVDMRCqKpom30eoRKmhL7AO4gmC0/qiOIsBkhopF9o
bOLynZ0TNfvIKpG4QWoxE8DJlD0dDVbPyXIL6a3EDJFtGXY6fTO1RcwYiWRtqAq5
TO+u/WAiDVD8DlnyVwnDMplNWoKjEsDtO2FkP1uf1TZQUBBIcSiBocd0nXdx1EoB
ZAOqc3V+TX+0X7O7FVWpljwAKtBzUsT/FZi2hneRzBCT1vlm3T2hNglgw3YFrJBe
j1c9bInfklDjs3m8XHBhH/L/VfqvKIOc/Tw4dV65+yHdiffCUYmYsRHI9Rleowb8
WU9CyIHm6mBiVG50xxHj1mS6uFiOmoSf7EoUZBb2WqBDR6bCmxWmqqRosB9fnwox
ufzeJc6jz353dqBUxDJAGpP0mbeYKc6ujxGRmVx4zWR2pqoOUBZIsXJWWLqyZgIv
/L0bsWxM6lafxa4x3yxlqv27dfqJmPmnt5jpAaVI+4b3idq0PGB0KVed9/zSNpKL
rLdULfHyhuxHgi0NQh2lOF44EIe6dif/aRE0pCbOLQr+sa1blqIHSct8BTC7nCK9
mwA33od3DAaA+SQhbLgoZhGamNdXJ8JeUv0II5D2XiKYTyNRB8BY2AF3mJrgBp+D
1g7pQO1NjWsYN+Jmu5aooWT6ISQbd+25wp7bl2QbO5ABPH5gVsUhjOh7Rfn3Fy5R
gck2cInjctjx3GT02dxexDMEWne6Ez2Ob9l5uKSdRD1scYJhm5VVJk9kx+Kb7e8M
dVfZL+F7J17ZD8F3hRp3Bia1c03f5NkTY0zKHdHI1e3Ao6SaLlnw4m13uFnMieWs
4Sk9qvjkDaYkJuCWEyKjbNG2UGU6XnY0aY7dLIw/Aoo89I8rDKqdwohQXAKObRfV
scFDnKxJwZhh1hxHYMoUBV0mqDjCvBZ1HsiHHnPqbS9izbulTB/vQB1p2wd/Endb
dW98nsnHrB2z+srqXIiMQrV6/t8wIFu5ussnmRwcqnYjqdyvv2G4Ho9ja3oqfICo
EmJYyZhEr171zBIu3dNtJA4aQEr+B7JBQ20e59qC0OQu2XuaNlVCcFcEWT+jEs3u
+lMppo57mA4LH+TmwukzhQMHVDXrl82KINtDzp5XPEOKQ0CdOGWJYszbwao+OBEx
O2vauIvG8fcbyl3Sgskuwt//fzVUw7bercn8XS1e2iIytg8zY3o2VIewFclGdjMq
TMeed61A5aS3IQr4fwuYj/7QLEYr63X323oeC3GPjKDB6ioV7HK49x6i6620meHT
SgMLOV2x2fbhscxbHqGOqv4e9rczt8G3Ql8WaZvWpDTXpFD59nSlDu++4v8NR/nO
LRv4wcUXT6wxHlN+b3JJqqqRtMxFM+Pbt2cJ8fF1OmWDSaszCeph7k22vHX2C07u
/KMleYrnBLqbEaNNroneYNAIloxseCRcQe/sCUMfwreJdR0lHe1yHfMHKvbqD6t6
fH1+4kL4KiAbJDf8m6xEm3OenQE/G0GLW+VToJum35aUQsUrNYJCWckuG5GtGX7Z
WZ3DzXHjpNCdeGkQMFXEgDe/NdMx6tlJr9wUilL3w83h6EJaelROQPP22g9v51zz
9DcMHAU9DIGEbWxPHO4x9urXtr9/3TjpXOdUpU6HnrAWIV7VqqzBfoMOmgWeB3H4
4IPzrxamY07KYOlYtd7AWEFcpKwEwfLWJyrTwGbNVUxAItgPW57eeLX2xFwXfCR3
WtGkFJgw3N5FiVaWPw5V6NKg3tPadDUlC4aLT/el4f3cneVwTh1Ogiaeq5Djbc4/
qhKJTHx5qCCS/FBnxz0AwKcx+YnGjicJq+7NoH12vrmIp45ZzNUnkf10EJg0WMXy
cNr4IWzXL61q5xdfl3eG1JzFUwBFis0A3imt3eEcbi/eCmW3QO9T+dgLRmcEpCyx
PUwoABig+vov/pdJLPy7AWVLCoHLj5G3zi4J1lCNy9IrvhHE5zohy5tqwXrBrA77
Ao8TLwvuuYuCLuxYSZ8n1fnrTZr007Lk671xIKINDe0O40slydzIaOE5miKqZECd
xF7RLU+s606PibgF+3xz4n5WKm5hLbAhtvFrDcHNyyBgFhG7cxEiAdZdURoez3Vm
1ExWmVUUn2oVcWIhFu1qhIadjpfr61h4Ijkzco8gZ1ElIHcqU5RIya64QiOWbKoR
BhT1c5QSAFNcKAnQDAbjnnCAMro4DwyeW0TgM2IUy3l0cjdc6If9Z63mhOmy7IaI
OUbb9WdshXAvtaBkHnrOCloECXfNbNPH77EMx7Ivc7VvlmAcAbnjoPp+88lHDNjD
gO93evAktVQVKrpywQbyE03NxE4ebGX8vCG1HVzfA4VrIt5iYEg9+nc6K1CSoj4e
MNJjdIRR2hp+X7kUDMnU8jcWMSNgvfK+EM5/zS6lQZiWWkh5WLLICBulnRALqRiL
LNA9lW0maEuacKBG9j471pWfogtS3j0xg5aa2FBh3rtvVtsAAORQv2YvmHFravZ2
5MT+5AP4AwFzwYlXWcVsQotVqBa3Qw9NVU+k9JjL5tb/GyjiKuVogH4cRhE/8ai8
SJ8Eln+Sj0Og4KV8yMnTq8fOeJ8LQD89lXzHL6pfJZAQRcgiFFOsdUL+rIP702aB
/3ZprO9JDpwo37BeH40v9kEdvfXT3bbAB0znXz6I8pusUwe232vHcmaRp2OG4NgK
XW51XNcgE2ynht56pJhixJ8AjkcTvO75x691/8lQx1OaOw+XW2XqHib7qN5hzfgm
yKj9qXzvJJAMoZa40lkV7dyB89zhDX7dVF7YwMH2r6IX+cO2Wm+f+rabEDxBvB4U
y8i5SeRQbj8Sx4EZKn6iD+l9Rp1pZDvsZ517HBkUFiNe7VdkgGnRl/RYWg1sGZdz
9YmUCjpNCeGQZ/Y5ZOfFywGnzeRzZu74iJWojIF7sECk5sr4VvLnsriHxCkzqPFB
HlhxJ5QW74FKXSzOkxHTCVn1JM3PZpGxrRn+wbe19UL9qe/FuEshwE3NfSAa+aUw
wn9CcaeFjofcDvBGJYkqcQOt1hTO9zRiwaapR+9FVZI1od4ruaf3tVhjeKsxtk0b
jGAd/7tsnlYcJmBquJv9c9V6KEcYMO96Z6IilXerqBcFaRo3k3+PbFH8av6h1zdw
Htrx8gfNTKkPP++b5TtM3Px8P1qaJInLipm0Nr8a1YItBKbkCSvKYJ6XGEF/Aqox
gUq6cF//ivcKhbq56STKUFwFPc0wuAINhUBFSaAq88lwsNgQutLUu0TzTOW4oF2z
5arKo1oUEW3Bd7jRBW6k8x3fc6brcdywv4VyCF6V3UYQL/1Le3nSRngjXmBjgBEZ
hfo6y8EZFa39+kDV4kcWKVnpmkOcwCMRJF40J6LNoS0pnSS/9RBcmsOR8Oy04oWR
kr5ocE5YmuPtYna0yZZnt4ez9Kdg2Xl650vijugY7BCpGIP53BOCMMVKcf65u45c
DKI8RuzD+ZYnXeMOeGWEktJmUxEt06EkskT80iCc46TxD6ulZ2jrNEiz7SDIYU2X
gs0TcWP9lFkQFel08O6NYSmwGlp/xQz4Pw/Vz8u3zgn3RDG/DE0R67p/VBfs/9ym
yx0Bew7XlBdPmT1QSDQ9AyLC0ycHyBYSi218Eqhr25RKDEbh0vIGHElNz2W7hS1S
gvDf/HZYraLeCjrroBCorEwgNnTY0mwhEGegQ/wS6Z8uQeQ9QYQMRjz4bgWhBVTy
ENnvgmAb/GFjB7C27vLzW3cmezGTebrF2ZOPGrk2f84yfmfndGyjq+j+3ltR+qDj
g8PolAPyacbLF2uqCTNEeqJumAHl2RBII4zxV6+Wn5bIqz6FWuSq6DXH36Id5aFM
z91Lali66Ri5fOgdc8ee2IcYA2jU8WLVGTzpQncpBRiw8aSS7SG27ynNMPNOickO
BvhUa9C+D+iMwJn+bL74At11LTnxjvn2DhCzUSzdgEO6yYP1LBDgx22uNd44JZAP
5YAw3hPQ6kYmZBl1niHTMzPzmSyE/R96AaxOtZbdwDRrIm06IdBH6SdDV1CBO3ha
QdowzljD0ZjZ3L0tnRIVf9jc/PxykiKQ9QJiymyYN/JLgvKGvEHA12v38jHzAW9+
aZm2AmwECw2DUCco2UjjRTEnwiue4SKNZKXCroaLTaOHJkZxMbdDsHbAluPd+wpb
VsmFHjLjQUzWxEk0FLLkqcgBKcQzNbkGH+WJXaPOF4AjaYY6D+6xWA2h1q0roXcz
hMnkiQORNvFv116poGndPufAhfNPtBtB9khwu1+tnCqaUdNmW6mimoaAWEbZ3AgI
7COsslUMZpK4JImpotnHt4y4tjqiBpkzg945EWZalUaUGHffTfSIiyiCRNDBJTpj
MheSFK1L7Cn/M9rqu8YkbVbfy29hsb4Ma3m3HKH8fZ7iReR5kSHl8f9M77FW0ozP
JLh1V+7ZsHI59n9B+iXJXS5yv7wZ8w+LZhfcm/T7x7XgikidQ9dHSKj5Y3dAzx6W
yi5LXLcq487n/zHBB4qyR6ePiZmjTSgDfoOXXBAl4n9WdaDo5WmkXf/Lbt6ciTTp
oWdDMMcHOGIAIC+ycmn0F79IAvuBZqlyTJhOB4vRqw3APb8G+mCORIv5yiz46Wdj
XI2wTTfKv39DIUS8z2VU4SYtDcYexK6lpW+8jBRy0qx7Lu7lZDV2+KUf3tEEdUKY
Cigqg0bSFuBQ1MT7Sa0OPz89iWKn4cHr9XUxho5DDcssdXj8qENLTUQaL4ZaBpqD
AErOfMZMUOQrevpJTi40FSsRCoaM8vkEDVESVzeeLlXz1sleNCY4oP55oaaG9/vF
oWLRYEh/gcT1bPr/89u3tzW4f4qzPjgTapyPxGBx2wKk9S48XDuDNDyktO8ZR5Li
N+0FofpnvsvrBclKkqhzXaX6wCSA2o7iT1Ac7vQT84ibCP9UvpOAhQTjc+GSAkBw
e3g+PhAZp/S6HIyIqPccvPjaiVtBx5EC1x3u9Ya7y++sgmKUEo5t+UglqTKn5LBz
JWwkH0mmk8tBudrHGMGK1LzOBewx4bdjG1zCGV6o+Q9zSfGKZFgqDpLACMOoxFr1
Fv3z/TLN0N7uS0iD0izXMgBo8xl1ySEx4sDXu01ybqVx3x50eF9u12eZYp0H0yXm
j6hah9nxS18IAGOkKbY7BgksOI8uPWCsr6gVlT/n6LA1/TnCxattwrrU0GS/RcL9
M4xqN2r7eley8lhwkJx8HgHIIfIZPWGJUvWHTI94Pp+JhW1eYHIVfqX6cUjnQSpo
eoJtSjYM+tspA7sRyZQAnjqDfP5ZFPJPQAyhhlTQsYy+sEXN8QpQriPFFd+rEnXv
fu0JOxU586/+e0SLOpvRCFtbD7KZsuKQHlKTQOICwuM/5RzOG9VV3M8lfsjDb6JV
MzExXdIWyPRWRYsv2DiSgjbTPiePgVV2oV9A6iRGv2UxMpZYEgtxABRoTlVcMd4Z
VHsAGS/VdOVzp0UcLXUQCi/j3Hng95OWsg9UrKWT0hrAYqBAlTSERAyObq5mU/aC
bHYYnQmcrtLyQsWOywSecKewkh4DE05uaXMuGumy4EESGHzyKsnMfmO94wsV1C0d
qQiu4dMi9ywalDslSkT83LwKu8K9XlDMxtcKFmX/0gAAnmq6CV3vf9VLS8voLPlx
51cGXvaH4qaVrR0TajibXXl3ZJltr6ydniDkQycL85klpGwrMRhOfTMFJCD/4dVU
1l8pwA5hYLAM0HNBwma9aKqC3y1/uSjOeHX3ltVRpe6+KsPPhf4aq94Wu8QoFzLJ
7lcqZR8Jf90WFamU7Le4Ig8r9/IvuDzS8MHSQypNDvzLXI/F1pzPcS82Og8NsPli
qrZnUZn7wLkF/7By/12Elph05yRFRT9f74wK4jAI30wBPOT/Iho0+mIDox4lf3bV
ydU/zK9BH3dWqAM0cFUPtk78nK+E9JgoYluJyqHTTT8tjuHZKtECc2TGeabc7O2o
NIhq9RXTU9j2olZCcY6u2WsDvEyoPGUE5Ap/vSU8EE+f+yXVkv84vNgM2mQQGGhW
uroHwxQ0QRP6lCj9oBmdHcpIXlykt+TiiQpHlEibt2xkCa4eNXLtmc779fB9BtNp
aqxg+h6JPzwqSOu8tDrlzg1LvUTda+kMBQBM9z5CbVDWZSSVwWrYcoestBj8wZJ0
nx14JDXkn+ssriZhAUaH5OBOsb2aj70Qro0eEAvWYe7SbTn/CEijnS+5HUeGTmaL
/q8Q2RzVbaJaLRetm0CEjU5wzockRK0CsMB1s7Ct5wRNVymaWc5W2t5MfgwA4x/n
XkMZBfHZRGf41JWtF5q9qkxl2qtXCAcKqfU9XYEBthsDGNoIfceDJ713FVSJqYca
gsTid8W5H3RtHzLlgwfzSpFxH7ioBtQAm7NJ4/ilniavHQA/xa7YI9kaLpmqAerL
5jpPKLQcw5e1jb6lq6QuMqC2tMPONUfZEHB3R3RONO29YUvKGxtOMVrIkfn8fCl6
dtyOcWXhOuLvGInVbx7KhmnF5kIg+RmOtEI6QqiZpl/HWWjrIDd8QCNyVBCKexRo
2qvRtOImKnnBK1sMnmD2CKDHGbTS838I1S1h47d9MnWpBvRCBfH6L+VapecYn8L9
CkI22NZ78S9l6sVxTkbKUqg8NNItqB+VlPHC8UFqVdDw7G94opRHMrKwqBy5Eznv
iaXCuolftCG4iKFfsKilStuFnGA8qA+txXa8I/j39EwhVvSRR0wBhSc1uNevRZO9
Yx+DfMJtcBNnasZWGWCdDrBt1mq313G8FMKLYtlIZPjwLTQhGXcheFjRatv8K5eg
1LOYXN7OSNWisa+ET2kbomYu7aTDn4cELcmX+wyW85h2XeJQbdKWWT8wNfNO4pBV
6cQ2JgtvuEA2xOXpSuwQa1O05MGmyglWAiqQj2//Step5VwDmkU+7VBPAldsQc+4
+Lytf2AAvO3BBb06BFOV6CFSWG4lo1GptUBWqkMOKBQu46QGLOpScFGE04z18YtU
KHA9Fi9neNM7xLsaY2bJTPWOx+Kf0l7J8KkKRS3zYx0VxdSmmNdvXXKczjq2m9O+
43mkCT+f7UVMAUAvwhYVMU9RHwv0fmL3ikj+3szyHfKKW4Hhu8wQ5hxtWo9FRgzP
+IfVdz4DCqrsKEsxHR09hf7zEenQkeKRRuWSrCkGTQS0ITxdEmid3UckAqd5sOXj
RrwN2x26FBTIT9ByHbshfNboyqrXVU90k5r8ltxe6U/vHcd4qfZJquvHBC+Mbh+2
Sxkea7x9AVK5S/Ljap/Ohft/DnKR2fzhInWV4ULQr54socj83UtDGVggZRVY8qZ0
CyxkYKbhUYiQVrp06CRknEx0hG8qMacJ7ROKAd2OrbgyxSiMSA0jwE5QBJF6Bdhh
Z9uCPvti8s4Zc+TlT913lX76C7Uda3dFNWDjLXFZrNscL+FuETzkNfDI8tT0h0Pu
9bfD9YaeQ6WNcwdPYBWpnDi/wiF3XaQRrzVPcF+9Zt9GZCapPpPL9OZE5dqqAWLR
KAcw2YNpTPC1NdPNMYTnDAvtgUaKHmnaIQqaaAKNAa9c0hmaSmqBlmdqCko6lPsf
13L+6qP6M2RlsW7VjumzWh1F+DE2ou04pcOa/vUODPcX/u8ZKaUY+JoE/pz6v7bq
dTMlRAZmukGM5k7b8aS8OoyCV/ePyY1wOutaynmKmQVhgCTRXJFUqAg3kL1yJlsW
hjchxnwXtUxnbeECTSQ1BlnuoyPP2vSS8A3zahyl7B9NBvF9+r/7IAYq+tbGUQJQ
AFbWjtpoVZ+m04C5VOVwvJKF5JTIScdi5orms560nVvIl/qoJOGKXAxJMSvVvPvi
KgqT7pwq11GLjhXWIMgUSNLz5AaDPbeh+jE4PK2G1RM+dYBQ+gKFmXl3NHZqvKs2
bksC2GWTTyyVj73j604YzuZe7ULYC5tT2uOOJbhGP0WGS/HtsTgtcMt9Wk3MFxMm
bi/FVp+b5NlG3fVVBKkNvfzO3ZeTuBhlXCH6w4FFMsH8SdDepRSXJAEfweu73QL+
J0w0lvRMqVMJLsicuVnSXCjsIDUd/H9WfpApTjLfWJY2P/DjLHiyvIaslIUsCIHG
pgzBtLloLUVt/ZFrn14aHfLzNQlbYwzfNTsivYocGSeXSZ9kmCez9QTBi0v0wAEe
9FhzpHJ1Hinia7nH+qN54FlSW1TFkftWHtkXqGyBUO2InS+p0ZbOpVGnfjqMBUaF
pQGEgghsOC4qfkoPFxW57a33wEY6RR/48TW58heen/HKFNDdMPMsUu8plbQR1Uq+
RfKsvf0jxE9/ny0FHwzBWkumaLverl0mVaWWwBqzQM8wMNvR4TQXTwuSywBLyV6r
rgg6XicYjrHfteY9/7ZHva9Vto0qfoGH8bwQQ8w0tGqSRRBphOn1UVjpigIrKG6L
yBvYCnyCbzK582yJ1yB3Mx1p0L9QbFHZZiE/KVR+2sY0IseVBlSSxhvkTjoGSh+C
p0dsbs1ZSBFBcW+bNf170zkeBjOQNRqD9J43iPRpwtnLiFQ9L3moo/HF/sbvEvK5
alZvHhhVUiDsWITFtTsLzLYjyl6DeEz1t2bte4jWBd8yH0K/eFg+4B7FncLPxlyO
NLbL9ssxbpzBPfMi9VyuL26BZdm8XQfD5cAOddait0yBjhqI7mNsoQ7cSb41gDoV
Xvku/xkiC4e1y7uUiL+uPecP5+uyLOaetrYpKGbvjmVfzOxxj+dWF5Q1xf51C8mN
WuMlx0C5vBtUkHqbwdBiLuwIbuCH8EK0ByZQQr6kXQH+9mRihi8J2xPzIdje7sXd
aqKCalBFZdgeR8WrnMyOG880jNvbDRSJp/6PSSYVf9LNv7HebQ+bBqhlgJ++WKwT
5JOiCNVJOqX1S2Mkw8FG/2eyqPqU5Nk2v9ACq99gW871ylu2ies8Z7vNrj+RXSxU
i7QW4uxHBUQMTRVa8usSzZJXYsIIZ4Iske+5hHXxrc0DZ20KYYL3YW9pQ1eFpPTT
Ea9VZz12VBe737iWcCIeG2Q+glH0aLovv4daXeCTaFVb8BxaxHN+J0kJFZNEioMC
9o4qmWh4zbBmU0vQ1G65z0lICWSXTHrx00uLz5aXnEg4C4O/TLFna0JWPYqR3HXh
YZRDvMhEJbeDlb9g8bepSaJcfyM+wKf2V0/tCQxcg0DrnZRiIQXwc1M1hun8rJCh
2VKrR1/4d4LOeaj+aK+Wb4k8C/fcgDlHcz9kulwQVxSfvHPOW5NgdFAZa+2+Gb8V
JhaFuJCnK+y5HtpGigLmi1Srub8khUulUsHpIWUdnnd/v5l4uTVaNTGglIjplBkE
U9rAov7nK0Frx08GDsfj+ALWPbbNu8QW6AZZ2FSnCm8+cOCs15cxw9AnanzKBYzz
C5mwnMjTV83H7zM134QpIyp6M03vPVD8KaqF1PeL7ojbJpisUEhKS/gL08mdYqbm
7B/Z3vNgli6/x1Fx9ZBEnY7Cj/thmZn4C6s8Lo7Eau5ncQG78UQikVZqdSn9cc0Z
2904HQYVpU+L7GuvvFRww5//dLRPQ/c3KjS1VHDocAGZG+I5QDktNs17AuNFlDpP
d+shOLNBjZeprGGr2HroIiVTAXghA/rr4PrLpTmpdkCPtukXm9EKNC//YniC+0/i
Z4VV2zTjgcpeW8ClrUHJx7yPSX6Xi/mdwgHIoANN0WOnwgwPkh1EkG6xrvBX6c0A
Xwxu6wd6dbZ6dJK7C78XkjAdGNSR42lRnNJ0nCMZY5Cn3wv+Thh7PRdZI8CcC6Sc
43BgeOH7mrfAMtDQ/E3vf+R8Htgz7MBJ9QJK36cUukCB8U0+XjkhBDhVu3kmAH1s
WOa8xyWKCkiFsZ9VLK5kcMLlk7shTu0n7OY4fVP3Vx7f+u5e+ZPH49jzxbC+NR4r
m8LY2k51cidLh5cAfspI2Coz0YUH1fZm3w+ss3eO1NuAGzqePadhH0eWe6wzmM3E
jbx+13LufFHVhfXd1HrKUKR/qULaGOOe2A+clJrq2nbj7I5tVvu5FVNVTUthUh0X
G4+zZjDveAeaWjh8rIl2jaewdnuuEI8ebmHBqxC2kzrN9vBrI+bXWU57rFXZLLrk
pUxDEL4RDzep5HqVJlpp+vfnrtLfWSDge1GGLkUOelOlrlii9UTDiXimguLCOMWr
kz5ZEesU5P9CYBMwZlZN5ix2r1xboYf2KgblN+liauFumiyKqf21xYnDJwuPl7Lp
i2mZOe08DkuRyWhfCrIK1BGsajhEErZwcn8nup85FLXs4IH7AeUYPmX1syYXrD0Q
1kz5KokiFHhVuovH0EODyYF0K7PhUdBLeCDmsoVkyzdk8/V3/ElcouVUzOHa3IdP
U28lLCYKguIZ5F11mbbuozKt5fMIRFQAgaWl8KoR+1ru+EBDujSkBvmCRj+9L3a9
bS+Ez7R0aD9bObKW194H8iFBeioVx6hxvEJ3l57zoRRWBZUIfviJN4i9Vfz8QkC8
X+27pSzFRgITo8TTkRk4+NMAKZMSt3PZ1ORl+dIf1u1alNXHkd4Q2CQjbaqSfqnY
PnY6l3UbfvdG+ASNiP4POGjl+WRrL/O/A3PsSDOIME0C3f6bluLueDZluKTpRkMI
guitZ2Z0vChULDMmaFU2g5uPykkonaX+S4LygcS8rB2JYBIJtgapRWjyl4r97vv6
1r7IeZ1Z+vomFTGyJJo0GDeG3CYL5ZxH+mrrhxpNQM2gkLyfC7RyFCoD6fNp0ME8
9A5imW3+AJuDXT5bj1yriTG8hyaiC25y2NBM7OC4PKCbiHyTMHanGTHpbURYnhcN
EhISn4CyL8GhYR9pMaYLHVGfYQNzY8v52hsSB9oMpzsH+Tofek3D2Lf5IcanBirf
RFTJUf7D1wMWkP63Yt/1Anrqy+EBC3tcddQkbQsQ3f43VcaiapD3urjUvMuQ+CYl
LQcmsPAruIozD/zCzUtd550UPtWr4DXlf8FeLFx8hUCzg24tFiYVtI5nM9+DOjU+
U1Z5+aMC/SxGLtSinoY5Qs4TrUJ/rRlJC1ZYCz5gzetlW6cncVP3BUd0euANZd2B
+eIDC1PaoYaxPfA1SSZfMkSASJxfKWTTQEZsBE7Zcr7w+cb3eY0yIDO/XtGAqUzz
GZM38AIYtjRp9lCqg9U/N+1j2/LWzGFsd3lKi3vCR3oDL5f/zaTYAk+EGQ43pLB1
au+Q/gXDJVvvKr9bUDVzjGIKylKXPxaexw/Gc2xfuoKd9+AWD+p5h+awkzBbNA2U
fe4dHT66WMkcE4JJWeROgceonOOPmyCRkuGq5BXtpmdwrL8vUQWFgINdYzB+VQBZ
/FMHFE+yURAr1uFMzQphVVdTo4bujbOyy1uxldGKy/gtarftfELyKLfy1jMAjtKD
PcxnYCC0hZzxA7LVtXEx7WSxCMOJaoCGAs6IdMmCXKZuLWkF+pF1+s4MvGZaIE+A
L4lSDQTaTjvDODIllMlxhk+wovd9oawnAW7W2BidEq8tp+d5p5UUaqGy2abg944Q
dDLkWqYCp2lZEPpFUxlIQoa1+qSxYSt9ajBsqE5L2wwr0oumr0jiGMCRx8d6mo8r
T4n+syNAVZDyFZ7jvuhCvs5d9sG+guPTqexc0X7mow8MpqeCuclzdxwLLA05Oq4R
COmnRS2EVXGIAeY/xL7gieT+B9wHj98jkh6a/jmTwuv4kQ3R5RXicXfS5PyXHlsX
Wilc2MtcO+WKemUcD9zDyIspq1o6hqKBRb/0z0gkGieZsnV5DuFf1gfRneTVYfTm
ppN78SUmKoGrP+zY0vdjGRo3CyghWeeuEJnQ4ycg2RNPYHmo03mSaKXz1UHKOYNe
sck5fD107qXHpww/YNaZci4x/KchHVFwukLUvaMN+8enbCepJTLuXJbH6KbWO4DK
TqDiR8+mk5nn19MCxCGy6kfIaybxrZjz2q4QTH76ybKjSCOx/O7zlptqhqovGTcX
lxbwxsQCPSiKSCrvzW03RZZn12XPJcShn0tg0WQq6WAWVE4qWzEO9vuj1NJg04y0
68eCRhpAbAHx9czssM/gqfBC9B2Fh9WmCtvqPSokysWu0gdcv7c+0i/Iz4mVTUVt
8v2mb/UV0U5wr3eXgjzosjRWgYz+Aw7HrVtiV2y0mhTQFu3jLn9rx0ik6oS/sjIC
0JfiFZSdjtNxD57wEXSw9LQTJHD4HoV6TCIbVVvBggjYMtmVek0u6BgWxgJ2MFSv
wjOH/ctS5E8nhMriMH1wzRoer1XyktYEL7MYJD1OT6wYO6JP6s9E0yTDnbSmPKLd
TQqBridI+1R8XMWMJEqa3O5ShMvYfMkxZb7t1UEfzSX/IfBBDrzeX2wE0IWTP7XE
eRObEjqhVb8xVQyIMgNp9AjfEu3euSh3G6qj7l4za2qdXdcotPyyO15W76NvHp7x
eaQcT6WaaVxg6gAvtNAk/KcrSZ+1+Y0y7F/IYd2bBibto2OD0S/BK0Z9C24PlMus
MOL02pweLAl5SMIK7Gxd/wlu+G2Dz6CJ8UFb3uRo2NPsjB2tzN8Fl7lGa69laxhI
ZfBrz3qsPeKajzzOtVtpXhbrz/uk1/uW6nLWgLk2YjcAUcvR0Lc22PyMFeMfKrdP
Ws0siRUoiZomKvytbqUr4hGRD5dBIIxugr6zl0saA8boy+gynM1nJcAGD4OFjBzg
PLyDZ9QyAk0j+5js1ILghNFYIG7hvh0dY+WJR6FsttSvvZ9OC6rxQmVZMRlDgZRL
jhE2BmPw3QewTWBkEav2PLGm1gWm7PMDukWBOsGjLojuuZy4VZGeT8+RReWYK85/
dAcmQnpmXExbb/c9jGyrFgTGPXQNUFm6xzrMTWX4O+9hYngCTGgReOQRJa7aLXZv
mf3SFmqwwypBG/tNRpcPw+FqQ6Sm8qu9H9Zi1P/2/pU5xTnsiDvGgn0JLG9sh7yU
KD2vtUVb7VdmisaFvciUHnykCa2WqsiP7x6j9VocQVTGsS4PpDK4RblNy0n5/Ugm
DxeXXLmY7G+t7OXuWqHALcPC92X+eFJKnBkSTaFuw7JJFm//zaxXv1WiE/KNtq0M
DEs8dm22b/Rn4zyeLL/o4ZOPigf5W0VzQd+L1I/YkY2YISg1YyFP7aWEvTyAlUss
JiNfs0dwI9wb5CLl+qhHuJ0b3SYdqVqVdbHEHm5T8I4lXkf7un4S3t/znYQhzefP
w/nZsiHlzebaPaKwKo8bJVd9wC9o0oscr5ATjHANuGRXTRAOJnPQYzUN7cELSW1K
vupb+0F1Q0Tv2SsPVvCcoP++MdR+dAEWBOBCw06vUye3lEKwjTa9L4KMFt3Nxtcr
NXEUzBOzUqrfi8AY6RCHZFY7BVfAp7N7MmjkQ/q39RhCqDRv7TNv7kuF4l34JtI0
F1YIu2CFQTAikpRajQ19NegpAnpPSSfXxGRoVBt8klkH+It5CDFICiWNGcE57MzC
ns8EF4hUQH57iqj9KXoDrw==
//pragma protect end_data_block
//pragma protect digest_block
6VhZe4/GDtSGAJ45PBy5PEkK0Pg=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
xz24mmALZL1Q6FM+HQ96oA10icVrYDqCvD1HmXh7VdNYT6keetWyjTtIaTM7jgdD
p+yHo6UR/pUQcL82Am3Rb8USoTogARonr0wgJpGC0pgZFWXCzVmY8k+C+cFPjZPz
do7fvZoWuFNXz+ExE4SQ802h3D5EQv5KWX0qMSMCeijZ8CFwt8VQ4Q==
//pragma protect end_key_block
//pragma protect digest_block
DDcYBxP9bmu63zqmB1Se507FIrE=
//pragma protect end_digest_block
//pragma protect data_block
k9M9yxKiuPIFPuDp6G1/6IV7V8VpcdUfDzACp3pJ86eWtuOravP5EOCPNNK3uamY
rCm7K5FJajYYIpesb37CsOEfdBmKMm8y341TOmQmMU4DPsx86m2fR9lobIcDiqxU
+Po8OaJkPTzJpv2xR9tko2ON7XKBH+nadbmJGLmRzd6/GvT/B/hHoFD36n8MHhQ2
e2K9aau2BmlOD0aX7ddNcXeHs9hFCnrYiTP1DjfWPSRJPLz1nL6qjq2/dQ+Nbtn2
qCYiK6205rtwzOefYyEuwisu8TUQ3OIDsj/UPADADf2tCP6d1DdMaFuZxSpARNRr
TAcmGTR9wQHKbr80hE3LCV4yagGC2++Kd4WfbZIE4JH3wt26RAk+MhEIHuWk6uCg
GXqPR5+rhWI5w0yg3/9H8VJYmIVbUh6ySps1otMF3GHtGuY0kDzxAlpc2hXKzufA
q2rtycNIP7J9q2JvvdSmjqwMF7soWRYAMXN8DHCujKSNzWBpBcMcKvv95UALlJQh
iR9iKv5nzzcop1M5k4/3fuXkvBfRZHpJfFcjw7e0TrTnGTBBWfobNQLQZrwGRSmM
mFAsDcrChKekpYBZu5++jzHVEF49Z3BbnDfALilinkh3YH0udGovdhB28PzZSlRf
zAGywKTLiK82G8LVQAR6TxQrH058QXTbbZH7aMz3DipuyAbczDdL7e7/wrwyJghG
IU/QTerAEUUNpCrTnlNJ1KrHuyHvcbPAZ0ColM5E4h6+fuGsVNXRcC04A9w1ZnJE
4fPqUGLzyAPoZOJOZetspb621EVletXNr8uW3geYlPLaO9xMUpt5ZpIn0teYR5OG
UrG6L5+MhfzGBNZ3Qw8QyNOU7ZJJFBIXrEj6bs9XkBUw8HaaaK8vjppmyfm91Zvf

//pragma protect end_data_block
//pragma protect digest_block
xtFiaUx9gA6hrjcq/svGoDW8cVc=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
b/qZIDQSJdiSl3Sca2r/Q8tgo1IZNFGcbH5bWuI+/UX/cfEkUUea8FZwDvPD6in/
FpXH/dnLeplJq+ohZT8jNki53UFoYj6dKihsaHyr+kMQQL+EY4cC82RRgfwwoqn9
di9dGH+TOWpOtunL3f/uxMhVlGRE3HQuLCnyJddt+CeBPDY8345BpQ==
//pragma protect end_key_block
//pragma protect digest_block
q90jgPkYsOuJpPjdKgkYjTed7FU=
//pragma protect end_digest_block
//pragma protect data_block
nhruV2j0hsWvH2nDZVcGXJEcSRXJ9Niy5dJcwJzuPQvx70qn3XeYo59ZIM4bCsnn
zyZJ8g4fcK0virQ5Dbf5i+vJLhyGrMwY7smbCE9XQRVhcHjtpn4cj3Rr3f+1xiSq
2sFsccimtO1KpPcGK3rHxH8aOT+lJCKxGV8myqmeyqVhY13nHgzIwQsBREIL0mPd
BnbALXpTNDXz6gZCKtWckLltckC0D/EcjcMgP+oyZ1BLH7d2ciHi47dGHVfpDoXx
6hgWlgRhjWLtcfJXe+2eWp6fiboRZnxYW5Dpe6uuqp0VBDp/x59yg7JCcytIOD0w
NOHO2x1bY8A7HzigM9TyV58E7aKCnPpP6xuhiZiQjH/mVQRThwQ54/Arkmbu+eGA
ZpSj5a+SPI5cVkqwfimzDJmhwQvIH0T1id73W5ImedP/BI/Rbuvc0pxaP6m45QPP
m65uXKqFUMSn7SmstnN3aj0dpUh2Xr9FR3eQot/sza2E0+iKzk3HmUr2g7vEwDu7
k4xpIOrb5r6iwOlNo7Z3w3+EUGEFEgCQxZvkSGCm2BzDnw4XaC/M4UHspQ+mT2nC
+F6vEErYqurTGGl7UCMFOj0wEpf5piGS3XEQCZr0mZsc4IzCr1hGM8YCE2YH/Z1o
0ifyZjXS7zG6u3LzaOHFZEx5rDlzvADkZH7DumDHav+FmDwdPexx+WEfTaGccHWa
OHT7pC+4zww+C52JB04K67pG2TVafP9Gl1sSUyxMRFDdZ3kAojO1CcZaj7ljoM3q
5hO7t7m3+AOuARnHbdYQdX6eTJD1up/e/S/lXIId/u5NWPboxaQcPUlOs2UMdyTZ
911i+7G/FGbpK1rLfmBUra0zUMK2vY+ZkjIPxkEmErIgfvJqEImjPRw4JhXOOPzT
6o605GqC1Kax3kzmIW3OmobHUqZFbLxbkR7GVtuci35yiklEQl2HKUygnWV+gqyo
nca0VFoJ2Oy2u51ifp6ECylJRWnBGbY2Vnk1t4pdAjBVw9ez5sKmXF61ckEGBm7n
mJZUh8o9uQwLHRp3qhquvxEjmQNEAlSecwK7oTpHKnOZhe0Yv6RhzmS/1GAHOYaM
Yrzi2aWfRYGZcMDw35eky8XKSBcwDZ7uFoApHwJY6qYXCPKO55D8BBFS/xNKkG1a
etNBcg5UYrt8MX69a0WE84jda3kaXg+aEzX9mvhhOyjblRE7ZdzfW1Uul/DxRj8U
vPsF7vW0lySIFazHY7PCcVZotusFSETW74SsSq/2H82+2tebWzouLFfeV5zKkVgk
AwLIaicsTivRWhXlZKrZcSpHsxFxTQlSaIvIW7ZO8yQ2eKVjFu6cM1ZrKJEWZu+q
acPqAOphPzCt2HwORuh/FKAci1vFgEWROA9NA2oOXYWzLWdLUGun/gmT7g2IThwY
geh0gkNyKTgnzXw0GiCgcs7dOvhCKuayIljJaw0NawYe9Tm2FZknMCt4m5o6zeiu
hTjNBJ+MqjnKJNvU0bIOEOZTy7lP0O61qnzyhxWDP6l1S6m5t0cTcb/kg2E+n134
6uSpCCvN6mWHTVc521iemqKhAGFopUGkPyLaeJLdyB2YraShuWdmlvBbkB8wKISN
TdoKcq8rXzH5PpOZ7FsJT2tKkUlNbjY8Zrm0ab+Rpzw9glrSXV+QHG7Ff+7aoHl9
smI50iN4M2rHCHguL7LEURypWzt09XQ/ULxnuMuGHtafJ+4hjks5RdMIs9BU8ha5
zESl9pg1iFuiYVt/C6ChcLoWotX+GeHWFDcgNbOzws3w4ulsYwuTCtRcO/u7FFBk
NzKqUC+HT17Dmkb2tH8gPzhocGZzENrYv1w2BbTckqJ4KTbkuM5thMzH1wSHtObL
CY5Wwf+jpQiDI5mZU0r5BLuPntLc6V+VNbj7f4xCICabWUXnofz+4IO0plkNyRfB
QJKwEBNTu+itGeXPdxYWJJB60GkTrFxrG1uCkq+WkzfMHnlagYU+4WwFJERvxjP3
nDqgCVsktXk7l1pV1GjF/Vxe5zCWMCWgtX5Vh1jZ4+ZR09vAlQINLxp3xXuRUYRx
7ITxDCek6V8VvVHVN2GCrGDoh4BaFHrt4ZbVF3LUT7WnNxy2kk096VawtjCcYNhP
u8C2FUXm48ajaK6GE6+aO5dPxyNq4myH5or3RDM0PhJdVgDAT/7+lrMefXAmeXXb
bpoyjZhtzZDX3i8qH257VGYQ+nGVIWHZFCoHWWPFZh7mHpOMweKF/K330SnUj0LT
8CRcTr1om3WXUi5+o0Qk7EV2s7q/fSo9lcsos4femYptsROi3g8L9Sc2UivYJNan
x4oVSiaiKo+qcG07zPZFKaukeZedm6WyngP5X61DkEJz0cTUTqXkIxdgzKRIPaMr
fq2TIqJaLdpY22BCwUGvHs9O+xEcTjqInkJYZJYi628x58pCPVyVj4o0IRQlOsbe
H9Eh3RfcdAgXjV/Ll0Qr4TGdoUV9gSQ+0pNbbrge9LDBlKKB5C8q0W+DXgMCy1xw
olIcA/vWQOuJ/FwSh0ERBeiM38H+KG+6id3VTXYbHjfjn8s8XNdrwlQPiP44KXd/
TbfCLk3KZtExNC+zK2SzQcGzgUZIXJ9iezCglGYiaURaP4RHUMUFTj3HYa0e2Jhd
SiGxpBkQq7UhR2Gc87kjtzxNkloog1eKn9n8Go7BE9izhXHKzk/cLgnIbxrCXlVm
qT4+y5t4ypsraPoclnNv547J4E7BXRH34p9TTUqwD8d9xFQZzUh9NRGP3ovxlT4o
NWq9vnzneIsCUEcoI8iK8g3DYvPGB5c7Onv6EO7iPQStUTgoW1/+JIo3PQIU7r2G
dCwqTwAK2pa1cuOx9ztqIsqpDGcybH9svGsgaS6cSGZJ7ZLpO6QZmz48NWK2HEOM
HkssiIHlhXti6s+AxgkhQ8K19R6QrLnnv7o0lwlYDK0nhMia9dKWeu6xOsd7H7S4
CktDH8cVLIrRIoKxER7DlZfDboL2PivVNbxYhztRG+A09nMMT5nJVRcy30X5wdeo
ppkiojpU16wl2vlb0RBeORLTJ9jXXdNXoZj7wex1Ddd6m8VIrYIBz7/bZQcV899l
9Jty863SnB1PlSBOAQuKRYLvOVmUjA2WTaeOEx/rrnGqZzWuAYzhA+niAPQ2dPIW
njYfFwYliXTnjLCyTIrGkbKblwcoimEIaTf8AkrmolI/FHK3tt4t+V51hbHhdcgQ
NibbFPPyQ4S8wfyib6jGw+wSwMsPSEb92NOkhc7stBhclIAqHjLSctoi8QCfFXJl
x2Gy732yziJQvW1g2WGlczz+3pLmD9fqxM2iD0ZGieAqGtbNkp2eUwAcDpLgXBD0
0G1/AYq4wQOnYy7dp9PblUeULYMriqWPRETke9Bkhp8ccy35ggGuP2zaYEU4rzpT
/8H9Dip42HANJS7HzZ1Qm5NHYYnc6HwvF7bOMDaGk8iFMoPtNoZM/hwod1UAD5Zp
U1i3j2HWDVYuD0UkrQRgAgfLZ7d5eVHKAb+UQ/TQ5V9a4VmvmXi8di9IHjoKWnSC
1eS7SikwqTerD9Uuuf/yichB4iB+3NnQsPKVuBpmCy5ewXLdJI/c4adHbX7wkqK2
kByQgYJmB6ZAkiD8DXwBZjSDguEA5TmCIZO8RKHRtaJH41936Xi9IpQwtKlnMt8A
ZEOlXoYv0FF9o5K7YyX0unByDT4c2Gt5kXdO8BZctv9ykzEU+25MnHf4J5JcRio+
4MQCYeSyT0IEoernRRP3Kp9JgZfaGPpV40H/9pEg/sHNM/+L8BvgPajGxXQ43wNx
SrBaF2DmOi3mWHwAvswRKaYUyjDDpQbeifEN4q8ggzwkf1G3KWdHyRBW2p58XmZg
XLuMg+YO2rX1w2Xsz3pQNRAodbGhyAuzbKOEUssAstbfkNOgLqu6GSSaPge4f8kd
74yVaotFOEkyPNorQhZ2XMQfZMR/hwuKKcbEA2+WE7XDY2Nfqbg+ueC591+PxR01
OD7uVlx62W2nkJ6xGiTZ+VKtNH5aeYWCs9tVKJv4rDF4nhPL6G0GuTw4ubchaPvo
huDBEsRSIY2R4LZPO0k2EFb3H15vlJ8amAijsCe7Ux2rlQrJPUfMPdwndCuS482e
vQMo1L3IhR8l3xSqxJuZve6TI9CWWTocTkKA9ifDjpOVhLUa518UU2WzGbivq9zY
CojYC0VUNRMnRMMSDhHMHFt5esMPC208ptrMrHKTYRM1tCMhJuFvuqjAqENcFf72
hhnXb8MdaBUA9heH297ynW67zIW1McJeGR7InheN9uvtt1aXC+DRCiKFRp4L22bm
Gx666P64o46eL4fyQhKC7jo4eKiEzCtvdkXBETIiefThopQnaKw0Bc35OA3XLD3x
EGsTtoELbax48WwMzJvzdfULmDaXJ0sCg+c4IN/11QZxkhYpOvqFtljF27Mndbo9
K5lDs2jnGBGkr27uHbQHBYFyVC1rG5ccA4ta6K/qqS7nPNqOfLAt7Zoy6MX8l/lB
2/fBnjZ1JRNOiAnFhY3GvkAGWBiTeLRNTr1Egkrynks4OXqbOVWD5tK3XQr0VrpU
l3q0qIPxh+gfCjeuZJGKZ70g+35v3CRFLCP5h+PO+XjeVeM1px4M9nUA4pfVBWaP
7U0F6On6foyVp5qJk0y3eeY8TL32r6ksSWZ3bpINTupLL2dUksanO5x0Rk4q9mWL
Lt9VXBw6jfJtXxq4MUQt44xR0SIgmIvTU+bz9Rt8FO7hX74RG9K96ZQyaEdXsvTD
I+sxDwSqNhwv/sOcULQd9fNGo6mSvpjZ08516xNwZ+e4DLa/rId8bNRHyU2qVtrK
xpogdTiZngMU8CkfKpiIPAF/NbnaUiUm1gTKObPMzY9dghRdHZz0lKJ6C5Q8kkyV
OW9bBfrvyn9BtskzENYcuJq84KcJfpP4QxtO4ot/4wni42pMvkngnhyzCwbHuuCW
ofu3OCl+3N6xhHfPLDMEiuah2W8nH3Phgmdt/Pzc60ZVISW411TlsG8anv0+3CTV
W8/rqE73t7it4yhq+TTx5gwFyeFYZcZaT/X5HP8o+irvn7vrpbMHf0I4LSUg9ACH
yi9I3UuBe3DLDZ5GBXVtJlbsIP/8B9dftUMrEJXfZCYSnbgyll2WwuYzxqZhug/6
8PHoc+Jg8itVXwFbW0T37GN4EzvX4aFYoS806cwkhBKMlGz4RAz9nEb4HUAimYXv
hq6MNaMbGnYHgkXkLY7bqErI5Fs6z5XNW5bvL+jO9KbIMl/nP4WR11O1M7Biprq9
As1WgsT+iiTB7aE+aE1P0Ux8Ii3iry1pxuhokDD7RsX1dMutPaLOXIMonsX38tBE
EC7wJFuzlzkQrTfeL82d01OaZ0Qi9uuTNm11ao7b2gWgGNCcd5hQCuRBTLrAtU2X
VY/0AHEUiM+W+c24LzYeTBNEynInVdFvutT4mpLwUNXpiOa9V+FPbRWlKNTwKudc
NpazShgFAIjw4xiT+qH53G+IWP9TUtTtRVbXvYnateAShGlkFFrBOrO0LUBGU1Ub
+LRzRigijOgGUD2fX1mCywx2yBP3mZjev5qrxUfQWeRbBmjjRc/Sf0KFRgI7vkqc
sCOD24hgBFgYfPOTsVH+tRnKm/R9frt8zzvXf87KVbzQhzZD2jgrdp+PXeG2btIC
PnZGRkqB8a0mhopPL+6sRiyLYoo9/lzT0EHiuTdNZcXBHgXK60CScA4dBbaP3DEW
h4Qxcn7ZTU2LlIrzoqDBYb7wVAo1x7iUy67ZWqeXR0s2P+F7Yh2aGATGPA9UMO6f
bai+ZD61n1RaFAveY3MthDMc1PU+i4RlckP+ZcZ2+QZMbp/267p5E1SczfPbpMDH
d3uMHZM+hK8mLJNrvMRMcsMXZG3xeEQ4pIdyYQAVFjEmINC2n8GEXFQSJl8g/JAX
EiwHqtLD/kQ3SJ82sS/3d0JOI0YgrnAl2REhsJuE70sFuorbzDyaTAxXZ8LcDkOz
9Iq8twJpea7OKGzSSejsPwPBKrj7F/8KyR0kLI8oirOjoi9Nqe3Ic3U0QEBfFM3p
qhtavF2h/iD6dS8y9ScgyA7C5367NW1bVNAOiMSzjqwuM1ExML9gTDGwhGINelea
OefaRTEwnEuuduOubK2nkwZBaua0n8esHBW9HYT5TVCUe4dBEX0tRrOxbL5sHVms
9IyTijr+7TTKlaPBfhsWg8M3Qe5ABUBBm62i6hUzjjaya5jeam8LcqJ/ZejV6e1F
GtRFpnaWQP/2TvI0VkBS6vOp8O5DgOTgkl7J2I/Fp50nv44qkT2LQyfe7S1kB2JP
kYRT3NUAaRWtlRRUsIe20nRwy2enXwDyyi/+w4ogIzM6b1qxBT1L13QbrPwUz8SP
34WNfU/9QINEOuu9o/5HY+LuM2IIfhWtdgxEpqPh3IJHEuaLQR4oF5Sl4Od0x21l
K/Zt2H64NOSvUIQnjI6wX+WjlMMK87seRpay2tTMnHoqEKshzrx4lJvPQgDpE/N4
dGVvXVmH9TpEWyuevEvb1u8+eQsBmDPIiCX8q0atJk76U0x/MlEiMJvM/4JBg0DX
Zh2i9cu38ImNzPnwiyvCt1y/VP2HnwKj2tFvYJj3KeUAUe+clrLCVgGv6M9wq8WT
NIDCVTiK8k8Qc/oy8wQsq7NXA2giD2Kuh9+QfevKA/sPw7QFbKm9jvgthsCkVJAX
WK127oRTMBXi7CFunU6hiho5us9GkoTFBvtX8m5ghBbZ02+03QSakXWM0wZcZ4Yz
Qus83uxSpNh9/Mkhcr11B+9d3sMHbCH/cO6HBIvNONBh5HndpawnoRGzJQD1s8sC
3rvSTuuIAzTIRrBEeY7Vuek65tzLnM6UEzvBTthhYee2uSqGVp418eLmNS32opLo
JkuOgSgV9kY+O6LC+v4CCy91CBZ/u2qN1aO3Aqd4/cVi5G9MZ5+KcZozY2Lm1cYD
n2C/FLnyDJVm4pZWbBPe7XAOG6dUFDRn2NzZysf3KxQ9HtGORTUPVTEeXUGFR1wh
4lhDP2L7c3NVZ4FBQSexvohvTH/ei6QuFY3dIGhRW2Gd77aMM+6YWe+WjLef5tHa
HBYc5P7Ba8MBF0E0cVvorKBs+Y39BrmIqgNq6rRuqzARHDizabDfnxtRk+Xw4mor
X3yBtG73ql5+rP9xPPYHpr/i6cqe+IhuY5/GEzltH5c2vl1ZcJuF4DqunTXFRKjX
/eRrzRjupwdauaDukpex++x2rwmK5nQuB1qp4VValEMIGPIOVDp7G9NuK130l4p/
GQhgdJ+fRTH2ZkBF7h9EP+DXH6/nlwIMSwdJARGCiYDiFoxgD3G88P9LZHunHdey
418hUhQhOth5LPu9VxdUB1Bv0KtCQUTjrq9FHnwLsmE5T5qLliS8lJ5+Q0sp8OnV
Dt9AdMw4RBaeYVDll+yB7lg38qEdTvVT8bsY9ZhK9xkr342z7xnbA0Dp/rFIqgI+
PqQ3n1i9zbAJvs2kVAzqg7Ji5jXEzfDJ37Ubp+PSCvnPmJUVQ2Oc1qVeMNtQp19Z
RYxgPQ4sVgqZ/b9P7YA5XAGNckU5HlsmcZS4+LI9oiJWPBjWPW1aZHC+9oCtk0w0
M/qqeTawxbM8f5HjO8dfGjjLHA4JsvFimCpRL6yfbp6Br7iqFMnaq5X1P5OLB76c
/9O0ZjBcIjjPs0cIUeH+/qEWc/9LdG6IvfJauv52dgUNaqTVHY7saGBS+a6/OSzc
Yms3Ik0FsrdUfgz7xsZtfut3lEyo/1P1fE7fMYVUrcXx9ybwLRlxqvAkCoxFnR8/
dx/3dXrzKw/J7fT14uLWf/Zk8OfLHv0mrW/x1HM/X8/YL9MC+p6Ifhlj9TZ+WoG4
CYkcIX/1+g8vs4ZWuNk+j0sEoC21muoOYnpzJFvNr7VQ1RbukFb1zzbPYrVai24Q
rqUrnDrX/yfdMwVjqXdRNhzunz5qbL9UF0zHIvpAzmd+oAikbp3EOY5QBHFtPUlT
Jhzx1lfaLu4/I7qU/i0i569W/6FjFqI97bkC5XPNUYJmeybc/eoRN1+PfcKOgWNX
SdH811SQ+/KaH5O0rF1ggffCEVlHfptORWhreUtgqiWOJhocxU5gZ0BH8krIhFTT
QU0Q+UP0CvLRFefT5geYtlcrA7rLfPHMc1dc0Iw29oqy1UkdekdfUNgdssRzLXCU
KQ5jSKqh5GSSpdEKKqYCleiw/mo+4rKC3xT31BOoA7AcmpgWaua7/JtZFa5IGGHP
G2A+XImqaz185YVVJynrz0NxMKTVMozlJcOFfycBMuVAVgH01RAq0/tr/4sTZNbm
hGiJ1tz5cZOuZuoZOTPxiTJXbMYFkG6231z3uJLr7j/a9aHjUWawkIoWwyYaSDVj
7Pt6a1vN+W9Olt+Ic1VBlfLk8HS1Xuymt3U5To1gozwIUEn9p5Spi5Ub9KkU0eiz
n/ML7gGRMAqWMPI/ixMCZZI/f6Lolz479waHe/YCWkdwjSghXIFXKLwVVXzRe8og
86y3KSwEyvR3s/gvFTl9nFpnhwNHBQIdbvBdbq79IsnAQkmp2tI8SxRXBScEhNCP
DrHmzVlBduCOEmHjC8GEc5UGjQvUjQ+JrUsr+Wh49y6V9NLABDq5m4StdMj5zjkA
4Pm/YZFyXuzb+kCeP7bu8neEiTn31sAzvorDx1izbjQ5rSBr8Gs7uLmuZLlDpsDB
Fw/47XIajQ27Qhh2gmh6EQT111NQo9qmXd7n3dNyeUgmwpklk6sSqB2h4hn+0Zg+
RQXuFNz2p5Z+sYF5b/fEpwVj1rvoQunH5fEAhkqxOZG+kkV12N7K24enRHr03Mm7
RF6McWhEWEkRmivloAcL7nMKHqL+mX/U3rNRGgMrSriKPP8s7fKj/0ean+TQeN3l
3BT9akP97MkI87HAajzo+rSk471PbWIlp+xMjSCyLH6KRIKnT+ZLAJ8Am0DfSnCG
F/tznP5rQNAF4T1p2BhMN8IZd5DyOi9QTQnYZ3TPv+JSkerEFia5HwJO2xiJcvEu
AXfIMSvFbepdw4zMhsXgSfFMDbdkaVOMc3r+3lIPpNMqz1txF/3zgo0yYkjB9dfX
r4kaHC+ndPdcg1TpK5acOZF40wF+xuJJWVZEmqHtyWB2kL0EUnLK76Lcy20OFoTM
/LMeRCu2AA9ZdTZ8/mBKCU1I//oPWrFYxjxtIS34V5jLnbG5Okkr3NzjGSa+mQPp
7rVhlSLBRUvpCg3+mgPoHyVo1FqFkRF77kHdFF0dvoNvlnBSqP8vMNdZ73Qax4Lw
3Ty8cWU99ieMgxvSq2thapYzaFhwp6rC2h5Yd/ooUyTYQRJKcBMoA2lnO0hvvBzE
BPfMOWySMBOBwf1MLlE134eZAJ+E7vKWzxM7Er2WK3EgOiWh/5XpgQ2YUaZbIzwI
+JcgFGWUdG37JtWY/lGlIr8djBJVJCNn6QaEVVCFnGcch3y/GnrBI4h3eUUeeuAQ
tgwv5P1Hokz3oTu6DexpmCtpqkJmZw7iIf9lLcappsfLWC5gOTaYQrz5e7CukWxV
jzL2G+ntY0ADNyAK5nqmHH4Kstk4qG+ktUMGEXDHXvm5Mw2w1s1o1mncVczaPTnh
UiuVSMSm7RR5TJG9c2O5mj2D1Sl4CZYtqsg4/ii6VSwl2NM7tQx1MxCndRGO47j2
FEI20rHsqY9iljZ19KYvmWQYFzwGvUwvdZ80sLzaxAqaGc2G95bj23eON7uNssd3
UCI5XJvL3Q7zUUUIGVB0NO7s0JQnSayBSO8AVR8eZDSbIIGmpRwJ1uCkAgJE2iRm
2PN0ZXG9+i/noxIHokxOhW4l9DtQ+m34PfxuogHi10dIMBVMfWix8pMTzkZxDjrt
XXJHNDWs/uFtbSqgYibCjs1Be3ddvzIJ3bPEWgsIUzqAE124qeTuph+DBPZtd+Nq
DKfvukMa3a89JLNqTr6/EImE/vgxkaG5D5QCoziwqhyRiGgU/ClUI9j2V9mRryZ8
FYTswJvneHu8n9EIPK0af8Wg+HYJbuZLnR1XO1wzMAYN1A0CuaI9mVjMyiRu+7XN
Kbk6yycnedebVFEptbZ6npctwvUbiyFpgHwziBZr4faVVWpm5pmJMD6mGs8MA+Nk
+Sy0+oN9Af6OayAPZRY30wEMZFr0tSUTx5aqNhKGxQ6XD9yDwpPpUgsZ2YdfrV6j
hr1m/swHCLVt4ockbbl15M/dMq5Zyc6Rer1YsbGPt86bvtKQo38bbhvCkojzftb9
j1QqFXhLjCKM0WuKeHObkq22Ih0peyX7oJbIzIxpKuBby1yrFAP9W6fZ1E/vSg5w
SnWWu6e7dwP2E7vEfVWdI2LxhYGRMGFPKuogyKCHJyOPK+1AfvgXmfQ5SnacIk3X
lL1rjfFx0UHCnit2ZcsTPaaBY1Ujigc4Z5wXJihKCEGYWfNv0sN6WkbJTqWet1ck
2oFxfFXhXq4SpQ955tk35gWNuOUpT6b77g5mZChU98Xyy7gvrOBE7UBsw36EtarE
LrSE3ApcD/n4DCIvLeXQB92+gI/9NOs8Pji01TwgTG+GGeTtdUJ0lrOjlwEdkmar
Idv8/GI80htuQG1t7tMQXkawe3qEJQohMkgmBrKBww66yjBJLNGT19R89lLvYuFv
QDXLpQZAk6x/2yDRvYniuBVZNcyb1xliZk2eSmNBKz0DOUJXhj2vRb8UjayU2DNU
nzZSeHZfFl/6KCvptmbzIrpJosIlwSPLFSUGEOj93RjGCEV8PINlwiFsUOeNirx4
Qqi1UZaR1IuwzvgU2UjfxLeqYcFZVsFv2ZZn2hy6Pb23cVpZje26Kuzem+qZQZiM
5BGPO+f/cSM64qT5KrFt4Cwc7d+rqssV8355D6hbWNlFhy/gAoy1DWauOzPtcAT4
zm9WAl3IX+QHxrMGC+qHcEmJgp1LAqDwyi/9OYmVcP1tyhTf+ZfmnjlzRn+CBHKx
QV2g5jfqf4XlQ5THOPXF3yl1GVcYJbaspXdbUtSlY00jVTXVSkqTvFBWpiaSce2F
MF8o0XCkEkTumJhlhuUjCEsmvU2HdRrcfUb2+7hrf7o392Ucrsog09iM11QOr3Il
GOBK8wo3PYODXP4wUi8D6BvMUUpgq/lDtL2PKB3AU5+ce4gmTRrPqPYWl+97LJuI
Eav1rp4/Qku7+/a3JzLABx05FmsemYijHArIbJ84hElHKNWqpLVP1kW9VRmvKJBO
CWNK85vHSwTI3dmpMT33pl/opAK0PGbf0kXHhrwV531ZIO0OCOufVB/MY/ajmWaB
d8dXoYRy/kXVVFgPromtQ2UmCA5L9WQ1mnfjjeUYU78u/4RrFcSlzW2V2HqszLX6
/UvVMknwiWBo3wLtZKCJGxi3V8qAzTy0SXuZQ26voynSBBu4vvM0gli6QBJe2s9t
ZkRWTJK/7cGYnop7ZI/s8vjsSOVv9rLdXJcRE6bz4XciHetsMkQfaVj/n3ylDsJP
6Ga+oRHQBxwzYCgi5cWy+d43h4UXgnHlbhKi1CuxkBR6rKOtS3hq2RmmA+cJzj15
4xMTvxbUDuG7KxkWNbKpHu9lvp2k4DL2nxOmzJDgSK3gozcITBImks8vbBTR3H2Z
MJGFM5BNz0yxCYGF2RlXvbiw4N9qOOJ04POGc03n3ecnuAnObFZ3XWlD9ywWEQiD
S09TjwP/Oop/IfhejG2kN/3PrG8xy3ZjhMZ7x0/adq3kc7iGh2ITun1mqNevsK1D
LXUTbNEb0PplB0Jm7kyDtEwZeaC0P7x0KyxjwX7mhz631Z3/of2Rnrq/arbKDTcB
nDRFHzk7gvo5QRCDQ42NwdfAbiO+nc1wsqqsKPTtc2dcHwYLmtzC5uf1KV3WycJf
LgrTkIl69uF7tNf2Xf82LPKs8/a3jvR204ew1j+xmLcINGA7kM6lUXVGXEzDOrvL
YUHdufsr3OvMXzKMGGczPkRC/XExat5f1OW7b0/BaZYDNtRURzl427kqjGzEiX18
tpMvOPddys28bMGTLhJjepsh83PDs1GIfxYTdKnjtGhKYC6YRbVwWwSYmHzG+aIA
Cfn7X4C9RRbBr3JblaAlanSrBY0HA9+Zm3d/RVNdVqCC+de/bej0BjubueWwqcWc
XD76nSfFZeJd4SmcbKe0vr5hujJdJRnHoOZULfMOKnBxtslWf0oorCdIzPOcEo2Z
Ck06MqAuucPhTrt9Nz1Pxe+DWgJycxceH9ozy1R9+j0vSUk7tqUfxIveHQqjfNAJ
Rg8Heb+wg8JMLD97a1qeEkUprfaJVKFkCVGYcVw9FRCm9ZXoHhDcjv8v0HDxuDyp
en4Hle5CgDVD9uWhSsApqlxDjrOM+t3SKhFtPerfF82wQAn+RNv6b9bz0WBbGLdW
qkZjY+qNXy/X9Dn7Bed4z4XRq9n9AAY0MQGtAZ3SFJf6gOonw8pWhwuvimjcgWY8
+gKVQEJ2rGXw06GQmsGgT+5/yk7k1tTHT67DUpXwgQlRDCFAcmWtzJzqsfwLlPhD
9vIPz9Ljd6og9DbyJsdTyNGyluWEE/ee2/fm3025PbcPN5K8X9hC7RvpKXwheyYC
rA5O9qk2UTnfInVlMZXHvkfopODyoSxmH5vQOE4jZD6zv/qlCytfdN7/c1zEb/C4
/MOw3I5O3hjEvBb7+cuOqoMi2S3J7gYceyOjJ7ztOWY2HKMbajp/mTncCwdza6FB
OmPEb+SSEegDc7OnTz+jZ9k7cnmh4tDaRCrhrNN+m9y0BBpQnUyor++GXJAvh3p/
iolQNf8kYHS251tunpWIhMoGP5ru915Xl2ED7GBQgClvOBY0W+rJzjyimsWneuJn
+mLUgJVzKSVMECg9t/UrDf+92li/Coj6/dFvvGpWlizXriD3Xp4pJFcm15dRqZwP
6Yv6pOZWzU78hgnAaoDnNM/ve7oTQabL7A2F5pLS4jWnbtSuFeNqt2QcIsJv0RcM
qn7axkXh5fzyHTiuLtAuo1xGQZSo6H/em8SKpvTmtg3CnJmH7j6Yxp8ObIPUGBmk
52e8LLEEXSaIpOXrmm5befcnMFt+9u3KJ2rW2HUb9GezQ2jcSj2hpd4cToTNQHhl
jmZ34Khk2BGGxSjcwjZOeY+OasK16AMNwsnV8wgzpLG6bBUSjxI6Cj68MSHMjo4A
qZcQ2Z+Yclx774eOrP4ZTv1CeWLoBoHwviFZK0JgR606J3GecBl3RrAeldVccfn4
GZByuQSnpyG6/14wDtEZZ0iOpIddeebXMv5S6AQ3vxfR6IVuMG2yWfJd3GZjJ5to
GrGzuvUSdoRWRMbRRhimOlQTsGicybwLoddKGZoBKB73J/KiOy4oGWj/dcIyr6DW
gTfEmxWEBDsIJgYCAf2NtvWiVIqm5PjHk0L0DmqHpZfJyHTNVUAUxUwsFO5E6o0H
8Ngi72JvnMioAYswEVV8B0BAf1B/ysaP6IHNH5lGgQy7N2iYly0P1dsNA3mChDvS
oF7esTe56eqSWyYIZHf9rpAv+y6sQpaofta5OwdEBbp88+l82jvcV7Ut5aFYDUy7
tipCdp0QqD9b3cHWrRNioLNen0V+Mlqg6HpUO/zCyFKpTwTjrchFZDUGXEu0yGHL
wKrl3mHn0ji1jtVFTftb2RiTinByv2KLy6wsO05PKaWa6OzDFab4zwrMjpBLPz1e
wc2t2CkG1ADNqGHHsee7+ZfhOwzOyjd/KAiuSZKb3J8ZwGJ+ZIgvxmiw6rH/QYam
U/flsagx5ufitDyoMJQRPAM/zF955+3ndJZs/HpxOfFwQKxuPPgVj2CpGDQo5uEb
uPdT/JqQRQnER2M38Y/D2D/qD53W+vhMtkvLrde9Niub6BPnsHjI6m1YOJbFsxXx
JPwwLs5lkrFjr7WmD63A9Y0hUIr5e85NjvzG162Q1lVh1wQbNzSVcmnL04Tfsrqq
GtO/r4hSWFgiaQpWXtMJHnLhtxOK7Cs9bQ2VKI2vo5rRIPoguseg1JARYEGGnJGI
gNH/gnVMI92mXuzozgsxRgPsYcRzCB7Q1FmuQpqPUMghK46ddQzn9iKjPXdidJ+Q
fNwo9yNQO2MWCcH4NNtBbvUvv1Q7kT4WDWAE8qzPqiRQHPsAVz8/jtOrdCJ02iYM
UmFroWEpTrLfn3QNAQChZB8bS7b16dumHAriyO/i8/mCWblGyJrkZiCH1NXWUqIR
QAghWZu4HhzGug9EEkA5Qh+CaXbp5YDAlYItZMqSGZvmsOLo1OS+wocTVx6buUpK
Os7XZvzUmRYwZWgw8MSyCsBGNOz4iUpj6hZqLu5I2kc+U0ahtJeHxNY/5eRumIP3
wg22HhkXWnW7txFo9AlNvv4KbNqP6bxW9/Koa/6fO80eWMowYFmREIPVj2H+/yfr
cQMwfQuy2+FspRCKLzzUwqb6uOWpdib2T0wJJQKHZnjPEzIfzyCTB3TzMuy/LKDz
w43YwTf7DZxnOyPxtqglJyHoYZ/rHTX5IvLwBh51LNR7xb4OofVuB0/CUcFFf0mN
GniziaVv4o5OWaLpRFjrHChiBoZe9BYzWd/eg6yRqdHpd7qRyylzDgsXcq60Q/Gm
v12BiFtLbfTbf234MoEy2t6RFEFVOcBdpZQa1AJj8YHF/0mVGzRcU0DOJdUJ3UaU
khlzQdVIk8bZ+a54fFQIsVyfKQ+LxVetfu97CLOcwHETdpE7U+ERjIgdRLYKMWCl
+xxr5XZFu0lMjGX9dok8DAA2a+P20rj5Gzqsh1+fFR515jT8c0jAQPxu85PUFNHO
Ga/29uziUEoihdp8EJNXJfqteZxw7iQOIE3XMgFdZTl+Z0yx3xAhBVPWFpCJHBWy
MwNGCPB6mRrTwWUaTmQrjAhVIreqnrakVxh4RE3iYXpZO/teQFUquayvLp2IvmRo
IaiUWlQf4vCt6hkuHXaVe1YizJZkm0gNlmOC37uqbpx8ibFviv2uvq8JXbvluPdL
vy1z2NgW8JdxAeo7fvIiXnx0nP6uUWfBT6fOmebB45/aW98+n2zpC6mBJo7wOGAq
Ua37qGRCGxLkfXTRHG2GFosvQSm4iZAOonwNqMdDjjDt5NEjMgES8qHEFesf/NLe
uw1j4SkukWUHhcK7PABkEM/IOYYUkGb2J6dalIvFQfzLFk1HaGEHXcv91PLQ9xXK
wZ3YFOKH/moWzSYimHnk3xrysMeNlwwvHElM0kjuPwTLbbFwYIRUNym86CF6odOj
lxNVobKChxV0Wl2KiBIg4avIO3xPdFLIPp/ocu87bptwp0ddDjC6nvUS2p19CE+A
4AxHFLTRa1j1KCC9O6ESd1wzIXBRlvtGo0BAyN2s0BMYAq0mRfIH/B02GCKXLz3r
dMgazhT9Pobzz/m6IZJzWcZOkjT41GetUolrLoMeHmQHndCx8kv0mulJSwRVrLZY
AyJVcLlCF70Zvq5ifa3hBUKdxSP1ivB5ifq5HmabcY0e1NcaxwE31RFq9iujZC1l
gi79/nn/AF3tMT3ovXopoymJBqIACZ5/rBcd4Kj7kISSfHKH1GiwmMYKylRujmpi
8yXpR7M9HgWVIG4GpK1vqBasjaAGwTQw4esNg1kDCfur/OC3tRkFDb/pmhSxfYLA
xzs+Z/C9RDBIf2mmTL9c7qlxQjprYfm2SlGBU9atJdEu5PBZSeX1T6uXyYPnfhzq
RIjQfJ+2jlepX831DrV5N/FuPVP0nqYYkg9DC3gbXuEZ/N94aBXlod81EHfT9M2s
Il6FdRIiWD+IdRKr1eJkOeMVHiOISgFNaYtqvuAnm18IXIEEVjtnotZyqlcHIidr
BBhr6rj443AA5ULZSvq+3+fwe6nXproELboyJJ6Q4DQrowSXbGbDqdwWpsSkQzwm
RMheBNA0fnhEuRa9wiVLr2bNspwBuNSjQGQ7u6J6JRMUo5xXLf4sqtFSKfdq6m5Y
HIN95naHK8h2H1alQXH3CcvPnvabSP6D0zMyYWF12RdugmqwxtdM3V7mN3RlLw2u
Rcfl0ys1ow+pB6VyGIazFdR5HS046Mz7IySkrlUvBDVM4wAJy6+sY3Cse6uYRVmb
a6H1/xJ61MzSJ80pL1v0TCPU0SRjPMkkfY3UTlcN+/5Zr5JPZdLV0GJziJt8KrKB
tkMdNsmfWmF2R+wuF0/uFFuNM8mObLvMIyl41W/IdlBqnO3X4nHbemwGIaQhpl9a
bXgV2aTG0oCqmIpEK8pGOG46Zi3cAy8xzZPUY1uixalXfU06OsrhpJ6s8d3J44Gk
5mGVa356QkpHHN19A55fnsRROT4Bdha0Gu4YN11siEeN2IiaFA97SQZ1xVXSar4P
4uMavl10580RjH1l2Y7c9XYbapnp32Mo+sONIblMtGxUIuiwHNK2G9VBuieEfyDB
8L3hXqoIKO1pr7wnPbnbdWEURPdHXLPrdjqz6+G8mIC+/n5ry+0GrILz6bnsvR6S
Ht0gNUlIQTyF5lRICjjbbOsSofJXB+zjag8LsswmpOrdtU4dULOYt3vn16nRVGj9
9l7YJH4FUIGraLBOeN9j35vke8u9iFyY+mTUn1BN9ve92doFrhjXldqZ104B1e7y
MaRwy24wmFZGdO4HsjjNizxkhvgSIDk29tn0FLsHVZ4oZbXnTj6rs24zXtNtUSM+
qLDif0B2r2tOnwBVXdfWjXbansFjtf6LTc72xZdB83rlJLqYr9h7ASRGH48PDzFi
Y1qD3jbQcQULdPSM1BpxHZOkRfilNyEeXxQYZtDvr8JjXGz/wApBiC7YZWnLfrha
eJ8KiPTUz4ysdU4v5zYNHGrBDo/2VxIBaBxEXQZaQENMIQaCbLb1sXHv1nB7fI10
Jv7Vvjf1d6VLdp8y/z1mAPc7l+VWczybB8jzGoeEgUzo2+N0nNIZgeZC0VmgSJ1l
9+9+Ck+7F1pEi7A7wOzrzsrbF/+laLGFT+pod403yxzGV3P16/1ie5ArE6QK1C94
i8JANjWPbCqwRJvS0cs5AcEr/u6skwZ2VxEJ+7HvtNRr9Z56bzrXwvHmRd103v45
QIcY6mHsW/TNqBLHLL6AGUt/ix0/RObHK493sGV8u0hxqRIqgx0TS3G1WAtBUqIC
1xW7UA2vowsUV27/sgMYq7D1CRqYFpfT881W0deaPn81KoNgYjf3Eb/Vq8gfG9k2
NUu0QamHtpPK5UXy9a2i70yw+KQ4P3j2tUGVZ3TfILAKocpLykMKQFES3zDyD/P9
oZO0IhHCupH7tlDOrrVTrC5OzE6fSJpIH/DL782/nPEj6obkJw41h+hEoX2dwjdQ
v0ROlbkqyyex8rjuionvXhsRV+KgCQSFpbEkeVi6qxcRVxXIaKNfEY55X/IUxK0K
/OTS8eqGTbROnWIEajFsZU7p/wPKgMLDATtGgAG1oftTZsWir8uPuhPLba4LsaYS
auOyXbfjhRyC0V2t7KZxv9xaC5Q+cDNbH6UDl5OsebhjgyLWDROFVPOkYLPOZKo9
7g2soBp38qxXPciBRk4uW6FnhTMSp0T9JeX6wnF45I8+Yu9SWG9WUoJKQouVU2zE
9G6ZqWREoGQFe+uvsKJjUjQgIisr9kTzS8vV6bVLB+BkuwGHceo752OeYTvQHVTg
btzX1IotJdgLtxKjmRohqchWyPRGMI+5iZ8h1yCXqaq1n4UBfGzExTB7iBkKoUR0
5qoLNbVJ+eLeR48fiHTOULJrwk+4w4Y8+IudzBsWL26EBGgS8KwmWXsWFB7zX/KY
DzrO1gmT1egIcjVWNWo8Bp1dB5CS4C7kdYjTUCVk5Sg7vx+tSYAaqVbRM4BUiYaW
xMWnwfeSQ3BNjnhrVerxA+f7Dyth8A8SSDrA6V9U+7f9UL0IFC5biWzfHMT21p4C
LeXBZb9aUJ/f72fOGrDalRm3hWKFj7+6i4FOlDtjKCgDTiBn5U5MI5dMCh9a4vg4
RJOhuYt1se7mmv3iVPFrRl/N839ybsWYu7yGoom5FO6gEHtMLHZhgjN5O6UdNlEG
VJ7+oQkc5C58GeQ0YasTqXU1xLgdET+PFrcSyc47pV+edrE2hOM9mrMAxZTCXmJ/
eWyW0uxFpZP3Qd6PdEKqndtOO2j35UxJcTEjrEXnGMMhIInCjj8ClVpGeLt2Jk1K
5flRfLCABTS4P/df0SnEc/p0aBnqNXJXaJF3cGLRhD6UdJUVVXQWw9pb9yXfxDM1
ot73TvRtgIp+cbBmEMspWsQS737p+IH07p31HvqKkRJ8PRVF9taFDOhTm8sy8E9y
X0Wyh60VptrOxf1EhdxCVat1rpYE28QdKLv+a2Jqx3yOTztE/gynPuprzFmPsjnt
/hH/10w/ySjtGuZxhmvbpjDxBkWt4pCcK0bWtn3/tkcEVK4yxWSUDLj0u7nG7/+T
Is02kWznvc0SXkmslbvnP44MvPBtCljATF30c843f3PJyt8q/pzWxJkC4DhHNG8M
qYJUcEQXuAdI5HJxtdH6BDAAosRICs4qCI8TyN+B1aCPlGXdljUn5/patWwz+E3t
6ZQG1wTvjMJ18IQjO0voaJ8JmA1R6RP39kS+vlaHmfJmh7hKza/iCp8WztAoAbx8
yqe1eE+Ky1/eQ8z1sIolMblqOFSJ2uLHjm5w03YdHkHVwEiMFJz2JVjacuBK2UO0
U6xMbhEWQftSB8jJbmYgI0mkHHntKKUdiC15DUAVQDjgOiiePbzwWyfsQ02rUdcp
vlaHjNUiczo9+p3n/o98AQYz3kZ1k3Lr77PcE3xPuQpiqS71LGHRzNviRwuw4oZn
w+GXtJDgHTHd+WDxaylKuIyanEcEOudP7xEbwfykIJBKkMWzjH3zMwxWV49bCDM4
yDmY2GgGAaWdadDvgfGW+Yx7RPMC/ai86kz37nE54KTYIUyCssAZL4SGBOzXXjbH
JEEjVQXsL+Of4TqTgKZbDQbp6TDTaoKSdVybtQzz/4/0KCLOri5U5L80mCAvvl2C
CtQeOON+6i2syWXYavIfQw2hxaaD8d3sfTkWtHEsCDL0h/6wVZA7Rt8AuAG0nLLO
b1E+/fWAfwgi8MeFFDKxxHJskHXGu5U1lAWP80L9ICa6O8XoiCmMGH5MrUsQPaJd
237SDSqm4Xmx9xNF3Nd+3zWQlnu+vFdlsdzw1f8BZWKuUHZ+0O+iIvLLz3L91nXU
lYD/sKqRFlzSM9nbzcmOC6q9lhR5a7kys1r3AYhf0/LmTUrmyOhayL1X7jPXnH/u
Fe0UQqF2iGK2fYY2sneVjXoq+qUn67DtGiBXA9eDB/8mFsknGOM6+SEmMGZ+xcgu
hTgekbRiXN1OzT6zUtTkASRe89T/qdWTiHgh+XQsykRtnSX2xzCwnlQt5GkJn9vk
LekCGaG7yrUST02IO30csJVQ82SXRGvWNQcIqSzBe5LXJBwjjXDnuC55QUGanK6L
sqsE4P2rErAC4KYe7vsxHyts4eSKZFEQt460pYJ7Ti0i7utRR+o+D5tata5I/SOM
Qu3AFUu3R8ULD1+EmqlsKk8DjFxQCF9PWE300N+aZNC9tPAuvNs15ylMIIdE/ULJ
ySmaYsoXiGgsMMbmJ60eoNbZ3Kjcr+y7yOr1ZO3GlHRXWmQn1VGJWYhRvhMhvI+T
vrMPBDIQil2X7ML+agHZSkRjLsFuwnf4Aplm4q84tOzLuJksYpsz1w+9Vw+UPP6x
/L0f/NAqvgpKNSOZ8wdGcIVPrMPHQCRTODZUFDKNopthhbhVwnd/WJb4uMLUSiYy
6fgh/WmEWtmuMU0Tl25wWVSyy7xx1Pp0Si9z1Tjo8ksOpsgVmQ5PGXxwQhWu0krR
QhBsu8YFDE2Z055fcOsZZLxCkgvnwwoW09Drac2deQ1iNTuHcZzppQnRKkgvT+cz
tgDMgKvhjwIrktuvEwL7IlXevlbaVMCa533Gj4slZ4CveURIkWMXntvZOzsliSoS
cPu684TWbpXSrlvfRwC+2fst6glCJEsiB5I/B+J0GrPZtMI8okl1bcuSAzr9si8Q
1BjBRSKv15BmYJLHq6jTkynlMJXM2tM0UP7G1WvwEbzZwKaC5At/9LsVIXHFGReh
YW7EwthtCYhYX3C0Y8tGcwALEQGr6CvumHzGaNdNDKX+03QgXg4KI0ABhPQJSRy8
gEDx928hdOCDYh6T11o3e6y8TDNl6RIyWroWFRxgHkfTqDe7DkS+q3Gmuh4i4Zq+
AaXeqiypW2Y7fyv27swpugIlBLkX5k8EnnpSbJs/t4FECdaitxMz0gX8dx+p0nfx
jwxzpO0j7W309T6d0ZLmC0Uzb001Usu0lV2/1+cjrYguTsw5meEhWG+q43NixTkQ
fjAsrUluTNBuS0JR3sRzkwaprvOpnBF04kBMZLG4bLdioCIkPDcHN6k77mu9cRUe
XfnRk2DGIKzXdN873lopgTHs1ndgWK5+0EJpJe8k1GrYIQr9GWnSf4BbDOGUlrH7
9PnqwHPVq36+u8qzDqyIkFoFzy+0YjlhuzOC26iUE0N9R27+uUlfNHNsGjxIY3rr
NARsh+nwCikMmSP67yTEdP8y/fCGettOe9hyVBmX8J9DfhWzyqGJRh1kmpNXdzWt
nDWQ1QNznLIkrlns3dB0udK9/mbmVOI4fW+Jot7AX6rnb3WnRs9d9Nbm/F3OfLal
Ly1WC7MRn2yH/KNPeOIDbp6DtRs2Ng6VPlb+F5HE1NOeuaC44heP2ELNEywF2Mr5
I1Gti1bla8WzQH91pMFEThjVXqa+rohg2tc8Kst1HrbW6JYnvxSMt+k3481QQ2eR
jXh6hBuf5Ai0T/tPLFbCW3EYqYbnsbUgY4sHQf/zKMrYZVFgFl/MYoSUv/r9zupx
sOGd47Pq38Q5v0EGDoyxPm8hQv7uCiXRohO9PAJybjQ2jQcPF9sBVl1qwd9zxAxz
tmmm8ksaRICUveJaUXIoEHY+r9VyBD2rSk8dmjwcxkmOui90UKmt1+ZeCwtOEf02
F00bD/f/p1bc6/NpkCsM1jh86ofAt1pFIKUv1XuJotKwpPV6Txt/Xtm1KcpU3mpw
1g/wzN//3qHRnwhlK/Gp1c3D1ehzuMi/t/kAKQ90q6H4LlAqPKYCTbyysrZDBwI0
zK9niHmToLIJYVVchz6QrFxC8/q7kewmNPZGaLBFopnK4sXjV8ryTOnQhiLbiYnN
aHKf7VyJ+3/urNjMP3tyOynRHydW+GdTmJw844mUOV2ZV+JZoiw7V4l50UxB/P6u
Y7KRgiRSxYh0RJ0hs2r2w1C14YnVPcIU0wVBCrQ2nxX9uLAJOEftaYqoXmBXLJM6
gPPQByPz8hNlgcCiiH0BukuAxWx6Qq/2toha/Lwx15Lkk/Jd2WBBtH0g3iYtUJB4
V+tbRZ3K0y2jXkVOwKh9a2HV7VDQD6+8w7tOxDZur0SHRyZMLhI9aM0wxvLNZwmD
sKVn95hZrOswlnU/bz1ww+4+rUtt7YqHwtnkBKItRb+3nNShV3v4lEuyod2xEmdw
kXneAH0uOW/T5wqSCe2la17FbO5TgZcjVu7J+JqYfb0QwlVeAdwRP9eElo6+Ws9J
Cnhn4nugH0twaJOTwi8S5Z9BEC3mtMGcxkT/zCeKVjNWsYG888bgdFYMiYqztZSq
PrQUf2i6612z23oYTiUqwCWkZGrXIw6t1ZW/RtNvXRUOCjk8Uns58K+JB64ngXII
gZYKf6mvS64ZOzvCj/Nkouu8/OtUXeZML7uI7uD0LM2KRAc9vHvSDTzCFDnl7AwA
MPEkUdG9/N5QHE3cRZOymxuRtH3src5Af8lDPFP2asc/a4KqzOe1N7t8325pSnNf
DlCXzm3VgAl6fquXLOn3Y2w7XPP+s9kt7SKlkHRO8BiR2k5qYXxjBGvEFiYPQ0Eg
Ta1sE43P5vJyynyF5AESg4jQj0LTQY0X9ajSVzTOhKJxO1XRDg20XsJjxVLSEjwb
gyN/D6l6jhMkxxr8U4ECGgorsnlFO2yqMUL33u3xSvb2cv42TbSHh6vdzw+n+wXX
XWJHumCIN3nzmrJaJYGQmol4I8Rybp8LGRoF17bQydRAT94l95C21bFdh7bQVfSq
iWQIORBQRHeoymMGAnZRupA2wNlUDQ5jBF0QsiYRG683uw2kH6IOYRQhyxPJOAbA
EYOy7yUsRofJ+kppPvQVb5feVZL/h8D7VSMgdyQFxus6gzG90i9FtZ7EyakK6JOZ
c2GByuRYEb/wZVXS22TaSlxzG5PHlBYDguBxQA2NAAutPRa5y4t4Pv1tzko6bcDR
S8NsXP8Ty0b+UgJyHvLrtnFZNRKZ9rx+qNRhA7AUjyQpEkbQxaeAEQs7I2IKYEVJ
/+RmO75UUwYSfNcb7iViuaIyHCkwDOkinPA9zh+s5NUS7Q9ecs0UJBpRPDPflYp+
SeoiVNJ5SuN0CTjOfDpuOwl2cP9fr1WQE7geiqzntue8xHw6cv3OgS5fNIHdRkUH
kSath5GuxiB1cXFFXYRHTfg8mjaFNCZlnVsBlf7RwZGSujg18C4ttJQDKPBMkYxT
QNqs2nI1jsJ3ffUdwLOx2eqNvgW2LNqCSyFlUNAjRaVuXQyW8YOopkHSvOxJ4F2v
1+F14Jup16lJ83ZDGejF+p9dbVTwACgqXymO94tOszJG93Jj9+IqGmlQhqaUKgNZ
CpK0QIxjatBpZ0AbNynDrhSZpoYjdlvw0tz0cP9Ip0NbXGQS4j8dHVw9+Si5Cxj5
2Za/LEK/20r9fLQKgW+LwOwJbk37aMz4QcoYJDRCVZtIvu7I+23nCzue7dKnVehc
xlavBiawVvwzdGOGW2k1gl8HgDYLVHB441Ieo3hz3PFKymzj2FT2ka9X6Peu4Vvt
3ZKiWxPUlvT7c3q9Su7eiSq+YfjSg4KF1s0IJXODQ/kCXSLYpIjQDZtI35ql13j1
NS2c22YdfpBCF0sT3zPyaqzsc6yguP16ln7veiF4LNITFSnWRXJ4IBUgjF9uvNFS
13Bb67Tnt09ughUcMDWyf8lajtmVG9xpMWSH73/WJIznk5YajheY5ubbQzVG1rdc
NqElUFmu+PUanSGTCM+IP/Niarx1lD7b6T1BMODS23pPx30yJ2xI2+fzOXQYf5Bd
fqn0AHAAXT1rVJXu/Pu3y4UErM86DpdYb5ANMs1IebG4Coz1oDQlAJmHc30vZNG9
yrXhiiqSigNVi2xcH2zYbmiLowIbwAcNSeniIkW8hi4+KR0L/OAsiXRSu8GmQ/fA
GJmjjJwD/Yu93pK0o03TxSZom0YhaWkBJdjk0n4XgapbkhBTKPQUGlzQuhjTDtQY
mXuZJtWjagx+ojwRf2jhoNOc6+Avbcn+n6aoFtn+D1jafaQ8H/PXPWklAfikd713
1MFFeGzwEEYNdvXm3bwtue98g1whjAtK28WKX/As2fwa/lPnB582luQzjHn4nVmq
XuyYFERFHlaT2yhvrw7zo5FjHscwZ6BPVoF4nEhBVRdWDVlrIETGlKHt08wkg8G7
LRUeyuwX+6i9BcnkJE3U910cUnFG7RslGmCPtXLjLjeIWqD+CIbd0KFgiZGyGJq+
zOyDkASSUufDC9Pe96sSyZJ1DmHFJ0SljFiVC4zBGEER6V/eG64mgSF4FNRwjVMu
TH/XAVhy4JAlTBEBZqgOQhduXgTjVsgfeIFfpYTxINhu2Gqw4idWLYnICbmtMRzD
fTtHuKUSx2NP4UkAyNlDdHgLKBJkx7KiW5K5WpkQ8bHc8wbkIUCjEul8BiVC/D6b
gu1XopqF0lWGp+Ms8EbQwcicExE2vz0i5BjY8TkCoFrO4K5DonWApUrfkzF3ktv7
lqrHx6OxRYmscIRWYiYfpYshQlaAg0bwK4fhtLQ97IMsiQd2VmlXb5E9GIskERoS
ljMyz2R4fEMLRHiCMpdsMa2WZ05wITNJ5d+rGiZHCFidtwWb5KJ6kqgG9hmmt2R0
+pk6iIOgMOiLmZf+ELfM8cs6vGFmBv9cgMDJ1EA7TtKUXIMWtE+wlXhaJnDb+Ge1
55pMBipbr+QzQth7M5w+h5jxnVskccl7wWYZBeH/zylcFWjN5AY3Fh+nY3B2TPp5
KLVxuhryg80SeNMSLSaiHt8A3X9s4Bi1zSSTHpQr3IPYI7eIdc4uYWyYBs7LxHsZ
ZiLosTaYv763lIkaUpwAGxkM6v7/Dn/nfV188sshn2ewYk1XHYXPo2X33iUNIofw
PDzSmO9yqwKyJCzk3dCp22hXN9IoPVs0Cxtidhj2/jCYlYyVSfmeLh1McvfCAcZZ
Xq3Dbu3tbxjSoGtpr12RYb3HqM2TXSZeNwMGu8M25JMRm9Mtoq7I+lw0Nfo9X4NZ
DAC1jWOwsfOhfM+fhaCU64LlptwHh+2G7+RoInAss7xFEn9p9DBlPCdyyYmO+mmc
+drwmQXfdmzjG/c+iW6UJZPXC7bD5SxXHhsAllT98TPZNGi23FnsraBPfsIoS+xV
t26QhzETZgMoo82GLgx2IIci84LQsgMk/ckxabc1muwL7UuH0X1l7r2wXXiYvZo3
w79oSxrz9HrkKK/HROTKRjI2gK7o5gjHRYoZu9zPiNnLeN5Zcl9YJNFK+/Ye4tLI
+aapdK2EPxJMtzgkrXpxlKBu7uQ9VWwQnEecJp9lWuYlQn8+VsK4FoA6SAl2/ftE
ZWxsSomtpcTSFwMlPr1jOUZkh9H3R7iyKYgT+i72Ky6uYX2NDTszeEfVIfkplmM3
pktkChN5dJNkw23RE2kZuEYJRbEzLxw2LpTNi5Nc6mRxRxv2hdPTPKYlaCmBEZxR
cEyzLsFMyQ/YJfESgCI0Nk2bc64DQWSfvOYLVbYy+xFgZmbw7KesPhrpbWK/zIE7
6SIHdNvk3X+r9s02cNlNvOAKWTX3cWrB8ausbNLuf/KUMPlgjCEbO0bgUtZfcXCQ
jH9VW77yTpUk6TNOirQ4nc3BfF7JO3FNE//KzTZMEvUPGsOfa15t519XUe1RVsKA
2Sln8js2XbDamFetGbBRs8fYbbRpgBykb37sL0hKA1HqHY4HHAhu5JMeaIxCacCc
vkoYikOgTIJ1vdJLXqUqFnwMa5xBA7XdSK4A2HxMFcBBqeD7GpYpof5MtfRALc/K
B/DCpa3Nhlb4iet8C92YZbjTEqS9N2g5qa7DtYE5A4ELJpZRwF6uv/ji6nxNRGm6
UJaR86/HTyeZYft9RJrCQawmMtTBoGXrXBn8RRt+6tTuweJo7LTrzxdSD8Gqq8GX
bSm5x0U28Bvlxm9ZtIMdUvhOKAYFbqS2ag7mC1dbyNRL7fcxuWsSSruhiowOC4xE
s+KYm5apC3Zk6pJdvOg78h8rBle3iqtW/un8rML3wcrFDMZVDvvNdb7AiAOFsI29
m/Kv173vsKH+wb0OFmtMstko6Y5Nv9LJsQbq96Z3wHhd9LnI49OW/LVKqa8ncSY0
mOLvytIptrMQUderWcOFqghVdjBX7F9XIYsD0Hvm03UUYphPbfexLeI7C9DVudsf
ts1iwpbdp3HTNDmBS5VJSh5n49GLPSKBpSjT8hZsRHyuewYz/IgkD96IJexPBKH3
gOkpiShj2tmx7Qe31T7UTZQWDCCNl7fbweHsflNEziOM8qaQWnY5KoO8H+/K7Nyp
uqOWKUNKSJ6+noSGX2XoqV4fa8PvdLvrNyeXZJ3Sqlj9KJUnBZDRvJVNSZODP16T
wUCKefdopnEdWDPX2PeEKgX1JJudLbLCEfWE6RX6XEy9ax0VXOdSFg26Ukxo8TEw
QHfSzMclgtVuDqyfnH6iAxjW4nfxylU9SkzuuvQaclz+NqGWnr/FYKlHpi4YkUeX
u1usv1iW3t2msOyHOShVFmzgBO+H2LxEbMSDcjDIsGjhjDax7Sy36S23dylukWYJ
GeWRcYFkQmcs2XbxAHwHAWOvRTFAWZzr34p5GMeWz8gPnO8uRFXDPPKisN4bQ46Y
BCpdX00rh2vRGSt85dZJUYDtWIXQqUV13lwuaR470XrxDydwLgjtZu0buKXc/axv
4HJb9BiD7J9SKVfIjl3e1BsBQZZVwuyavrxZfORy/bz2f0EEmOpzKnXgdByEvF0Z
tUC9LxD/UmEjM7WCljjbmFRFcMQT4LY8JBsMGTkTg/mjzUNb+QSD2sUjfr+gkWVn
4jJLRg+n1u4kUaxFY22DjiB6f3cvV/yOcG7mHubUbdHL0KZQp0WbHySa/B/VZ9YB
619LcuakjXCStW3pVmEGkhBGoJG6a0qUPRfwr8ZHidPZBu/KF7fkSF+tqi9klRCG
wWcP6LqkeWW+Krj+czJjuJNLmOTHucSPiqeWExBU4kUdlFx7JKgV61Ez5m3O7h/o
T9Tcf6KGw2Bb3uCnmCum8zJk+3wcyLFRurk5oP1ID3gR+uXfTeOyNLwBI19NMVNH
Zq/IXVVFdZTjnYmMd6kgK00HADKj59rqNDM4vRmtW8zloyaeBRj4vOk9wbrUZ4B+
OsGMlzz8+4RnOzSmuKSrqNCdjLHtmHdrgFPFTtkRoH1wRGM9vxTkLJt/xPah0VpY
Fy6rkpAXjBhr/UKR8zd0YsZFMSomQdB6Qx0rPjt38qvddWFb5m4m1pPkdHZmZcSs
mfE3YG7jtWABKwmuxI2cO0P2V7aFsVtFNjCOwa5FIxw6GzF3Su1VtO4KLsZfSeqd
8Yxq2/pVP3PpqwX9q9m4FP7qM6E+4Qk2x6ODrf741Mfe45Ayl1preSsnYUkeYwuO
+fh02X6yQ7/Q8DRR0iN9utNYt1ZAe7yTRJea8gGLi+Q++FzUOimO6Zl4sogPMMQS
L22NEheBuYH9oBPvAWq9BNjNgR3PJn/BZgI3uqkpDitnaSB98BhQrrK81nL/4Mqp
OFXmXq9TAXGmNrTT02QeD1u1AJ3UP/jFLcilO11P7h2bBWng8kFWPahRQ9oxhtO4
PyYPTWS+SZSdlOiaiVWgG/UEhD5BVmofiHTDK2mO6TxmWS8ca3Y4NmL4NZ3LUEP/
E9v1v3HjtdxQ5flzZt0DsR59vmOal7h0sXjhtqHEWFmtKJFVEy/USxNiiHvBhhqF
zlSeGKqIO7f3N9HKro8lgHK7QkIjxLq7YhdI71QeDG3hCWtGBOftXT0rewjYJJcK
pu2X5vt4sXgU2N/bwogj8VDrtlP7d/Ch9NdxOZmkvdnsL/UcRuri3N2mEWl2zKBR
TmhGGEMdL7rBUQu+xadxhjTsopYnOevSdC0l7pNd8M3AHgPwSGT225lP3OL7oJbR
0fgcAzzEt0S6GEscFYwmYZtbGfpHm/0lZzS/03tBwTLrSqv3CAurkvE0OcHAYAG5
dev6DqJJQqMbVcI6aFQ4zxJX6qgFB6271pGtrt8og0usD8KJANRpLsms3Jp1qcXh
yxGKbgba+S9Z8dT7Wg7xQYoNAtpr75cd/QojQHrU7h1oHpjt08+yzPFgo5bgro0v
7ca0xyBD/3a5uUNqwClBir3EzZlzLc8xqjw3tKKgMQQOlz11cF3KcpEi4x4VWsGQ
qnD5rmXtS0pwmpEEFer/x5Q7mI8DbKYgJFA6O3JqWjZ/rsOmP3x3sYZj0HdUbeRc
aczl2aHHpLXhsIYX0vQm86xM8pTW6bPfXrmYBUeNPwjoaBpMz32fkPZHgFxmC6T5
l+gDygtBLBbXjMWVS6iy0z9CO1OP0zyWHlLp/pOQ6KtBdSSsnh1jRlreV8MDBJlv
U4UwLBJeYYJh6ZUha9yXDOt4LhxjNID3/DaYhytq8+oTh134YruSW7SVfJS9W5fF
AhbruBSUdzZqbQsEDkQ4ke+mdEbHXQHYIrwRJpIMj+LFyxRpnSEcI1qA842cCnrE
QIb3IdtFb81TxgXWXesIz/cQQ6fP3aPvVnHLuRI8118DGiOLPEseSSNWqDzDYlb/
KKGSBQD9N1w/znZxcpt4tjnjQqOo+5Uoe+S51vIbjOs5U3/zd1fUL6d8/OvtVofG
VfJUoSNX7WvJ/FFawVOtORVFWOUc/art2ZfVRlNA3lyuu+PuPSm4gL9QaiHcQo0U
fHvYAOG1B7YkNCQkFcKW/vj0Q0kN3RLRN9UMvUFhWaDZV5KzyWRW/07SgDSj4TCz
/yg7mUtNYLWz4PurfzkqrgvJE9m+JRyYuU30uhAODXms/PgrejXa+tNDSbsX9skR
stiueJG06XNcbe0wOrryJssZUCJsOz/Zn+lFXXqQ2w/ERb0OXqYKOnm1wiL8ykve
ZiDR3rth3tv+HBd9IYeDtQqV1xFi4AoEktPdhjYMH6u2ZFDtCTSRhlf/f/lees1I
E05thjy3Y1z20oFQfsLT9jY2ftFwX2XrBbDJesAWBcdhqkkRAPb572HiaUQtg5Mi
73FZrm5L8yKau1TSrR6u9EGxJTvRhL8teIudp7F+OWtDu0oGHXmjJSVKgfX9eymY
uTvs4jTicpgzCA31OKvSmyNyv2eoMSIeXOcocao4qSqdnF0M+EMS2zP3HXsnXAJR
gcuhUzeeBaIaCB+qZ5svwBGhdxaGjE93OWETH08bN7zlB+SCukXwAL70C/aGaN/X
/QHbDKG17v9cJvYgUnpiw2/lSjw92DaY/ZKYMdy4L9OhFtq5/lOiW46XJCy+3cKV
ZcOvTGDqNz8q/ODVSXA8yp7vT4mRNHBHJr8U8BhNefrGoeMBW0PEnYRcV7XLBt3m
QWwudLMVfLfxO9Oe/vO7yVrmXpLX5jkPysmqASvHoRO7szzBcl9wuCl1kI/ITliX
tJCffRfgW2+wgIobqW+/APEjB96+Vk7GvSp+OH3lXXk/da0JiJhlqYJ99k1fSceR
8FXKx2y2mZdZHHq9VVj5gDNg7AArmMa+PQ5UiOmf+cxff1hx5JG+pH/ebuBMWsVZ
BgpRkP53jf6Mqp4mbYUhhii/85ZOWQRngNGG5HpA9tqJgViZ+UFiuklCytKPHpVN
x7zZ0yCxCTYWUxxR5nRdKtFNn2sg1+7bQb7CNJdxT9SDQDKcFEcSQ9LvNWMYwcoo
SI7Yy8aJUwkZzpC3KFVNfQjdr8t2+51MXTb1nGlw6nixexx0N6bq4VtblgM+RsdH
zrrsI9rH2czYinqQwWBM6lV79GK0eKjqn/4PHnlhrhqKPEAk2JnULpixrDqwcFIk
/I2VfDWOVu5JO9DJSlPISwRIa/f0iE84BddwVrj88toL3ET9Yue7XaCJSMD19bqK
JzurPD6TgoNpWWMMFDF8K3TMWPz53ix6AndytiNG77yJD6IuCR8NbAlGvjFcvyW3
+PEDF8Isu6jPD/RCmnaDRd74PGqFhh11bDs1iX1o9M1KBM6Y3sDk/+wOYQQ6OId6
+jxpum/Gf05+uzjP0ZVIwZd11v6VsFmfefZXqyBcgrWhqk4NAzwLzaL6IpURXRGx
qdn0JpWz+ubjwhBg2ogx5ftojYtMbgXLqw6W0RY1NTBj0fhr+Db8QOvKFJncnhJf
T/co0SaB1OW0x9BmqQcujmCEFZxnhmI/X7NoV0/TKH6uiaxOXnkLwv2jC2C6RJmK
tiOiTq/vrsqS9MpW/vO2P6yuAwPy9Y2wNLfy/vFDaxVRvyH0ON7sidqwNRtrWqcF
wURQDzc99hpaSKo7YEhkFBsnJt6nQKHJR96YAvw3n+4sWfys/rjB0qfgGIb2QHkM
jqGP2cb1oe35rfG0wfGsVUVZR/Yf337/ddWLYz64SUOUqpXsIpe44RkE/0anYKm3
j58er8t8wb8v7aOMg0mbn5PXoZXfxQaxXKPsYugNe55y83POlexcp1L2lHmc2n7o
/A+oAQvsZZLrX3oe89oRPWp1iG2Z1giRptMdid7EYWbUWEt/rBEsZ17gnVRiX/B9
DH+j/1ezUT+mR/pGDQrYyifwqhH2hWsL4jVR8yHP+VzrdmLtP6IUyJN9On2CNL/b
Um29PTiDOh1aCXvQLQ1VGH4xjS8Fhw8hUpVfq0KL4MetyacSFzQDsHTQz/MNevFz
pI9B46tPHWlnNL8zmkpLdu8xWSJPM3A102YDG4MSsP03rEVJsv74UiuijV2xinSM
zBITTPZQAfDtp2vZkN4i2U8ACwY3cNxJFtG/CK9CxWk0/C2zl74q83E8u6zufceJ
tJB+LiucwxT9YUOtuCxGi3bAiUnd8UrB1NxSk1voJyTwBINtlM7XM8qg+w48nuX+
8V80A71olcAJ5yJz6qpAcdE4+IIgTp3W8mgkec3BcUFY13Gil4dxTJAx+mkukeIg
SS50ts3P/ZyiWn2QjuLfQ/5TPQ7XUyBPQgBEYlu8qrk8Q/IXUndklQBnm5fcWuSB
8Laj3WUuoE3uCq9kVb0jzph34cCApCeMAlWPneA4vk799VQzTvW69fTy3ByY8c42
lVHbvFd3brW7IlJQiKNTmD+Xavb52uetx/m+xgmMvCJu2mJGkC9t/CBnyrYQe+mg
9N0M/78pTn7GCXzbmITJ6zVmC9lw0dIsH8dBcA410zvbKMdv1uPk/ba5sgR/DI2e
b5Mtsvvy30SKriVt15Rv+EiAe/sCGivoKM02wzXrRDIC+lZaJf5E1p2ycuGgIcqT
5ost9qAMXCPfV0YwL0/A0BHZMttuplECbHekg2WL24tSC9HabuhCGEyhY9EZghGU
t9MV4TPDhXyvPYjdjj0Dk7ywO0OJn/loWkO0W3mr4664KuZDxLGVzfY5V8QYLNPb
z8RY8N2xHkNbVOLrJlxjdBrsFQq73SDH/t8EJh+9rZeYKXPfpeNiRtC+tFcPcec6
8AZG/Cp2sElJ/rdRaodrEA+0Dc578Fzsg+WcdZyLfCcUuYFWoOkxuUSI8SErqCk0
5jfx9bcgG22oJAGg9sF5Y6NG5Pc8IzWfWsOhv6yLFlDKwP72N2kdJns1PEyUgGzg
imL/MWW96OwIzHK+IA3Yn3ySQt9Iz9McWznkB2xzn7YDPxjrNvr3fUMvlrsGAK9d
9PJFRZqf6dmoyiHaiVNBjwYE+xqz/Vum0KV1r5I/b1PbUGW2GS+2rIoJomcE1DNz
N2wF0OPG2CbrW/5r8EChV+1R4seO6nu3G4s4wpVKRCeqbM2lG4otf62ZPeQ68GBB
TpeiWAuKHwW2/95rtCwoT4eiiEEFOPfcKpJUE5+/zkI9wdxmTHRNAR6zVRReRPlj
jlqM+nbb6KzNrSMR27LnFtil/bzdN0PPX7szouf3o21oHhseljepc5bsm8MADjs2
n9HTXBVrKXzYl9QG5KI8KuOnBkpboPvsUDoOOVhb1DKWPaOT0vKi7yT+wJxSdQHK
c4i/A2Ooau/4wi35hSKwmX8d59FhP5oFSrXSvg9J6LWVYM8Iljb2AoOSvd29q+/U
ueC3madF/hK1TWe/HVJqkjlXATe1DDT6kNLjKjfvTlya8JNUDemVV6N7G7S5KFw0
QzgfaotLfPQnPuV3zWCdZ38OpNQH0NQQFBwcsAOtWdjoXh9vERjcGZVM6K6RgPN1
jZMi9QFvoUgQOX/JpDldgqtnZZGetZ5X+q6PYPNfsP+BK9JWMjO/ru/LXCK7T9wJ
8XJ0bvNDPTnWRM5CLyE+QIrial7CSmYLY1Kptp+yNfi1W+NVbm4tY2AJ2RAsZuKe
q8trhs+GdCKDXJE+ct701S5A+Ad1bQPfQSoX21r510de1ouq3DIW9yjLN4PZoQ/C
ZpF8qgxMUng4gH1P5crIY6TgaX6B/j7esKwuBwTJE1R2QjWtkglu3EjR6GxQCkoZ
sEFjRro29Zc/BnwqykWJCf0jql2FaJc7F0rVaC0VWGzPtbxs2X5dsU65MjRyj78r
4j6qoqXsDVxx603FTPC8oBwny4hLVFygkCLGnjSKAbu/T00d4UAZLLjUOUmUBabi
99dkKX7qDcyW2zWgumTBrlD5gq/t5E5iXEY6hoSXKR+2l6w6QrNjaMNMrFl4nXsP
sjKd4bmHP3+TIDgH6NUOuGZGQqqA+lZ5QpeaoY0RBy7HLtETdRYtuF1VtYBlIzB9
YRbUqc26qWxj79yQFBSzGdRqI/HM5GQa0ClXoU9GSVvu/5NtSLXCWFAFzh+rqr+j
fYSdigHkOFdIVHCO6+vhCoxsRSPFoudDErOf3C4gUAk7OKhF30nldntrhPoEaPeQ
fJHV4QrgiIWgqOQTId9GiQpwap2m0o4P2OzmOYEYsvpmoi0dyXTt7dNV5fLSu+Lt
KIQ1UuhIsWzKa6W3zsgLnVK3k25Y7HSxhoxUgn84gudNtdpiLC9qqJPEdhg2rs7C
9GpHTMyeJycdtU2Or91Ppr+gmTZOs4qy+ruHIVQncmmiGSE21cJ0Q6NEGbV4mLVt
XoXStr1L9PwOJb8eWSFSPIYn1ue5eUL18rMhiMT4VoRr7NcgxZ4/COIrwxmaEf2e
JR/F6IXx9zKOLUbwRJit1NW0ZHvA9rj8nbW5MyraehO7afmHjrmUFNFDM930FPNT
tGazPQwTDvzWDVPXZ9c+z8XqiiJGBEiDX4HsyWeIQGAfvoJbotx9iowqGykrJIHS
29XitJw8SfJmVvEKlW9uWXUGnTQGHToOqZH+4OzjrF+S4nhEZxRN+fkOwKOLBQ4d
mzNQm4RYs8mVoHJ6Z4BYD7t3DcMegHGqqwwZ5Vx+6ikR0Z96Wqmx3YL/BM8Zf2g7
ZCzNshQsh1IV6ObJhTytB5dXoHtobCpmu4lb6n0iBYaYyNoX3yRj5KbeLzaY0zga
3HKNlwzTmfeMPDrKj0NZlqgXniXnEovha59udPJFE6xDQ9wbFDqsjd/2hl8R1WcC
swxumJtRSnfrnbHA9sfoiw8l45uUSBsNQ8qXwlC5Ai32lTQkf7AQrvIOryXrYLWa
R3K0RmFqZLn6hD5yc/YaLY8pTKcEPW8QBbbHhSnwtgotvB0FRKWiTX0QCb1RoZcQ
lQVXNyCDFM41vCqf31QYTlQkXnrC++vNpv0OYcEOmtJV5k2fT9vpbASnxl6ttf1x
oQPtqP/dP67FzdJDP5dLcnMe/s7tjjatcwZkfro+NFE/tgQhYIUzZmkRXGbcIjhv
x6umGqi2n8Of8lRZPma9MKS6OmiUdi3Dze/CfEZApdiz7mVTu2lk6vK7g0/eLKoN
ih5jhCfkEIVKEEZoTm4eSF8jX0brXkalyk6Ey9YimJLw9clva49qLjagsOM35Hau
Sd8/W9dXzRiGcWViO45Zg0ku1JRvSZFaEMd+KUxWuI+J4pQAIKFJyYtAQbdv+917
kng+7LU+ZAQD1/YqdEBwNa67DjDI+xrBBfzyaTc1ovTkDTD6c6nP5+FJ65/4k5JW
EQnJ+38pkQpJw0UVZ+udJ62BTTxd4ZRZb3nSU5n5edXkVwEFlGWVibbHZBezx8Hw
LCZP3JjOIFpVC+kBjHRO0XY2+9fFjkc42wkdXV/4ILEAb/rQUf0cIvYcCCVLmKkv
cKlSKYhK7NpZVIFC0OS45jhr/gOQfnGha98XzH0/zOiA1DsMzq68QTG+T6wEVm0s
necT4vDDMH0lagseX9CkpHLEh4c+WxT7HDzsaB2Gpi87ioN1YIYOaFmCQv1ktoVZ
pjJt9FLGqxHP12wYAh9VlWLq54X2dAlzBFlWtX1MirG7IPiCoMbYiwQtj+op8V9G
amlqwPGYwZt2QWalnh3XrSsPcmzNzYLk0fiU6FN6c5Imwv/25oK7VlPJxP85QrXM
hiUplEGCm9RpGT4cf6IxymCgiFUGuDEi6zffY/S88EwnaRBAUzcgAepywK8fLJjz
abnlaKSr0FucUijfairvUY6l3lHRGpQF0W6neWA+9zalAFpGIuxLlTR/uy7ksNR1
dRAXutYNRJfzrgYBNBXZCAGiHaISJIl/ADoACO/lxE+cxWScgsHmeXvHjeUS6jyZ
24C4Z0/a7D36jSFtTZPyTzlF1uucDXTUXD1ZzKJKXu9RXQWdYyGbGaCbxzBwrv9Z
XWFYx/CxgqMaUys0+Qo6TeyPb6iazYMAmT2lYP5xZkFn4TJ8JHfqdaxBegmXpdwl
62JxH8K54r/Zlfz1amNI7fiP1jn6WOa97AiHoPg3to8twJKYHI2cK1WkmJLTb2BE
jYZhcI92Y2e2pvlKdlbkJhC4F99ydw5XWunS4V3lJAsLxNu/07+teRmAaugIOQuw
0kWkpDBXMp8d+y4xHyEK0IfBVr3zDSXe9/HFcbUYHhuwCc/bwR4r0kvQtae219M2
2cchyh8X2yaWuFCr71BoVFYlmce01uU4diuc2tbCIxCzUvfXcyn2odoAnVNJm8Qx
83Girj7TAtpAiRDJRbogzBABji8C+rJBEiNhuHT2SQLzRKdkuguFGaEc7mlVmO8B
+90NN83HzQwGQKqXewSp/rb/a307PaNekfH3ZtKDL+K922Ou6kv7Brt0KG6gd1hG
FWqiPp2ajrL2iKX6ELoAY6cVkmpfEIjGHLjH13kaAjmns6jFFubytSLELU9L8ntY
W8F4J31inlTE135LrAJx2YWvTZWNBx/jt1BtYheGJXtooan+kWqXjH+11rSeia4p
Bf/u394EMJC6sitGpiiI8JmP5/KSBwOH/GXGEaVM3DaV/7VUwZMK9sGS3lXDGjM4
LqRcVpJftKM2bqB1860gSXTuTpjRN7qVH7/6daVHY/qgjAURQDJTQ8Jlm5LZiUly
r1oSMNYCfsJmyK/pU6cYGv5doTA+Xylh44FdPoigt4hY2Sq9KhYFdN/xvoE4mwPW
Ajs7YexxMsFqH7C+fTNAITblyEs99Y4XsZ89pLVzjzeTnoBWn1D/+1YYAS3BYi7i
51yz+qtEWnEgmMZcBY/61pAWEyhL0zZ6r26ruiFgfr75UoG2vS8IfbIzjBhDvHwK
zFTW2JYclQLMM4gf4Yx3HbWl1YoLN+4uiOtHhUImD6i5ws2GswoFQjmffF3uVbSO
D4kZVeyqF6LJqEGDANPm+U34fSyCcRhj+5sNP8fVM9/dNIjgWFrYfnKuXDZ4FaW1
uvOxlLtVIU/QFswjSjVjkLpk336GWq58fQX/hzX29ILHleoJyTdWWLZ9oTQNquDV
rLoendqwNkrAiDhr7zsXXHD2jT0XsSid9kuaRMHX9y8OyTwWt+v1GQMkp5tJ9zQO
Xh+PYDj52If/CZHklbCra5XBggBKfQzHniumXE1Mem3EQmvTzFDX8ga6BBdTjqZx
t6UWaLKM8MHzGRzEQVCGfPQasw7NhR3nt7zvGxiYk1+6f+hI9nKNKO+09bBin5GJ
Nu0w5ZkUz2bkgzAGI0C10NrePg1/6aydGABf84YDdxspBtq3HweifdIdFwxWIwPZ
mdTZoZkPF/jPhVl4L73J58+WicymEuw+l/3DpodUawCrZ+qiDx6yokTdZJE90CRC
OOVYXK1dr4CqBf9g6iAKjiwPL4VslxxqZPLiLFnF24ETM1o2z4vb1mX7Jeo1rDuO
1QImIxcEP8+3KT+4dybDU3ZA2f/hjAMgAffbSbOetz034j0LxaBeza7b4m6znXaB
1E0Qid01L+Bu/z2B2zlwINXN6Mdw/1D1TIpwYfwXYH8cO+09QX/SpxTgqzCeqK46
2fVVF9Zf/Y1+Tw9ChUOxGm/78/ld8aHbCKiebnotgwo9z3XkploBRcCk5hN9r4ss
zDiquYHmg1Lh2mI/mrzJ87GBgMBmggnCSh9WqNpfjmdncAysyUVA7WnmHgA8JVSg
7/m3upqyp0vKltMpGKx/o2RxAn9qRmlUCT7D8pysJsKig50tCKbadLaHdoWzttxg
5Vr+kanHCI2BObW31gKmwS7+AIojyQ2HMwF0vO0LytyVJ/QWo88dRsJQ/W9X12V0
svhZ2kH6UbMLCiD7z4b9qLjCCjMan9lpu4dx0cY3F4FQidm0/2CkVYDTpEwBujVz
ab4Sa9DMs6EL8PDIcoURGhPR75Sg1SLTmtN563zOyzq8JiHyQNjfcjeHWLvsR61o
4t9t8emlrldAo/Qf60X99djZnT/Q+w7NbpxZ/Rxl2Hbm0nsAv5zDUnpParDV/B3+
M4BY8BAcpS9PoghiHcP1vPtFvIbz0SFW7GeU1RMv0YDZdnqQDHFtcXVcItkAb7Qr
fLxQHmy5+yDAmkoiY7TXLLj83D1c92KzC3etVwnukmRUpeYyneH/bO/aX3Kz3hMG
VX54Xeqmj+sfM3mD9cCNcZH0KiFjxWrW/ORxYwA2fsCzG9e4FbwGJZyhbPyetcyZ
5/J5R/HDAE0GvY582koCWQiftH0UhPM7TOjD/wxIO4347afulc6vAuLdPiEbJj5F
/OO0OfXxkKsJv3efNVfoKoOMp6Myuq95G0tOFwDPDc55+FVkiJ3A1Z+821MZtze4
aMQehYi7oFN0z+wQ5RugFakRhSm35XxzcdF3u1FSuBOrhW1qvJT3TW5rTg8utPIA
pfyOQ3QmT0n6jSDuiB0n7xIRWEYxrO4Awzlw1crCDNAgs51svcjNY0WuOF9izHTy
QKoSYKrdyEmXKS2Rj01G20O5oEXffqHu5heTl5TigdLUbJ4ZNYjVgPaUwSCxooV9
1RbeE+NlHVVQ2GHEagN7pwfmVr1ZF6N0JcRBOCb/0y2JmAejeIzstlW2T3mxVkOR
V1yrSh+fO34RQ6H5lYgmNffzqY5ETcOo6tD1o5U+to9L3oGTxF/QI4iG1YLWrbB2
PKVPV1CyuDKWg4X7J9P4IdO4vmu0vIciCE/5ems1QaJrSXjrq3pHL1E9bEemJLZs
sBmapg/Nc7+U6KR2VCkunRHbnrH7T5WF/Wq0qa5V2pv2ef4P5+ZrBf2nwp4saxg2
oNjqOvuJVCFs64+sHowtR33poiw2z3FGqVwTFYo5pTDXMCZYj8ta1Zn2bUrFhAxt
MinP17IRoz33MLQryTbT7iuRuO5VNLR8+mij1zqY74/IB6B00Li3FxOVyhuOOaZX
XEcV3FBFHN8/utkqSTON6pHdsXjhQUibE1YcjE6GTYxfNvWRKbnvaocZl+8rLrU5
2ox3NnnuXLBmm4y3wG/RA18wvbkxYOyoLRek8XrNu6WV6JS/kRE1596KEd+/cEir
nIUiOgXYZg6sHQKyVEbyqevN5pcyzKMkk/5CcW/qHeel5Rtu76NimJRQT2+crXAH
7YgeZg16hNvcc9aC2zClST1pxAQwmoqC4GSXvpLbY5g8Ur4DIgVfRnMDUFhXJuHY
7Gb4vAHZSN7GG4SA1iW4MH46tMVoBaBJZLIZxA+MissDsBkZyXHmh9S53DMRFDfO
Ap787IQXpo2o/WmuXWtpeyuh1e41H2f2XDgP2KMaPxCQJb7ut9Kr0rkCS+VhHVh7
34MQLMUBzCQu/s2Z6QnLUbhTbnsxXFRRkenCns2BM236ErTpnotmF+Y8NErxgK+z
dB3LlimWCgFZi7KV2c2nmGs8/p11C72iNmReOfz77AjS1yIZDRylg9aXe8LHqVeo
u+P8CK4JBM/CHxlTiVf0qaYeG9MvKJ66ZOXmS38hTcKa5uE8Ya+etpHh28Smy6Kq
tlpXhis9OKJmyCluAqmKETIXJss21MTOj0gG7Ie0bdBRVCxBWQ27e6FM2WcLOL/u
0lBDi8IwG2Uki5U6BYx294LevKSG/YM0dBHxl24sCEg2LX/sQEzTVmY1m0NpYNqh
mOWmc7bInetUkzCKHAgvKQCEVzfPZyrWQ2EmuWv6fb8kBNZK8fCKUA9HwA75ljYQ
GNsM/vReDC2IdnEgvj1EJ2xT8SXweIOC7o2FREAHaIcnbN2n3EZqb8KxgGAqS5NS
TZUDI//pykDNGh0t8P9F3U9URPuDwdf4DnOju8W4BKudonE1pgjBvMtYYClLXR9L
1dUkCCSv/zLiE+aMaOGTaD6leecZxGhiW1S4SYjxljDPh2dfsT0r2naE77eZkxEh
qKNaX+q0g907b0+SucmzZ3EZOQXSizcr0p4lYoM4kXR/WbC7l+qkFe8V+6Neev/w
5zCGgKthBmD+O5AhKpLitFIFa5VucPTkCii8UGzGE4hebNI1DRYHUjxVqxwhTKUa
C5w2fgk/KCwAOpIsmus7wSAXgJRjhE8Zmnxc1j6RunL9BirlSRU/IfJm+DAj+gUy
ONeiVWV+hKHjQJhf0aX5lscrVlsDa0aFtcSBy0ETdNOr+hjrsKOJdpVQPkrRgBNS
jd1YlDgLT1+H8xeRExzRI4YHWy+nEFHMcUcdPcZyFnaBRsc2iy87wg0eExT0nUQn
y6tGNkJTO3+EFhXeBjMO1nZBcbIfgUgR7Nhwn1jPpALYMoWpJEG+xVODFzjdE1Ep
/M4W4xwafwVOPKNBIjgZNpDvdIhzEOm3NAXIWQZeF9ptYf2rVTKGpWn18q9iTHP4
9/ZF0y6XY7LB2++2AuHiLLiifo3RIMQyeRtvAL9/+RtvXc3nbmeRj1xsY00/rW/p
A0dwEhBChlI7FXgxdRYnzOizdv5aeC6Zojdf1UUvwzcQsYPfvgjNa5MfKUI4Vrqs
dpflUF28MQcWXiJqluonNoTUoBMG/qYiNQ7qyGXBmpXSddkI9eXe569lmU+H54Zi
tYy0EoDHR5ieBtVAkl0EZ8ACHw1QqjmZ2OIrknzFADq+oF23H9uxpXjlrxNRyGsk
8Pe21pRDG7LJ8JI/nwPNtJRR0OhRUf4ts6yYKedq2911znns8FDTy3qwvhMEPURK
wBAU7a50NTFIbgkqHiyGxGqmLWnrD7E4R6NGCUj3TPDAVAjtDoFbJjyw+Wq/KT01
VU2KdFM78Ku3VyrTkzNSLG/FLuweAq/PQmHQOR/QO6uzGOoXLgo+dH3S3TFUyjYI
sAWKVf88E3uHswGtzGq3aWASKwda2k9eGX0gsTWehUSrvSmHw4LPrwh0WK7Ar+/9
aOmlTxPHS1qvJizVlvdSS/Ou5FIY61BGYoAwBpaKahFggSM8jaRG0ARygr0vohYZ
umhPPb0PeRM+9jL4XKueVTHxV6m0vkwHnLM5nqAeytu5iWr4sfsgSl2V+FqMNECm
hCQyWKB1NgmHbtUcVqbgK/LfgNljuFTCzTAoQRPgysqzi9RpIaT335vlgHci1eYy
OoXuPd5K+bixKzifkjrPavMU3AQPUyH5mzsMI6PjMfXn1aoHdh8dUNru0n6Jwy5e
cYp6ouRHrCaVVJlqLMf9AAah7OaOvdGvbGERST4t5/2GQ5uIio3Hs0xN00emN/ck
pi4cohqbBcq/uAtjqvsZJaK8UqVcM8DrAL1mpXBnS3Ix7RzOq+VoWWpxScaaETsp
nONWkEvwr80xJPhcn2PVSiO1Xwv0CLzgB4HUy7dtUf1v0+5XFeKIoh8n3Eorb7y2
n5DDyBZO0RWJj8/0iGzUbpKnnK2mrpmGSJPYKcG+rZ1n1g0US9fKvm4pHbln/mir
E/SLUZIN+AOMRobKS1m+cqmBiKvgElAaITWZ6vZ8MAk6BvaY49iax3Rk4AZIdknu
nqgd2wO5/a2FsgWLCBSDHao4glavLdEVWrgN24d605bgd/IP+maowYTR0TlcrH7o
G6uf2BjStaquPLfssWuxXuUS/w6MUGerBAclD85d+7rS7HoPY+WwXWlAi4Ftwuo2
QZd2kNd4k0GZhqTNTluJj5YtELYPY/tNg0TWWKyK/52Efq2B6bpzNcoi9+JVOi5N
yGOHFSLrZGCktcEKS3jY17AfRmWiibtMAtDKKefJsIgP07JoumyGJJaLWwNNC1TZ
e+3ei/vt7w7Sh1X44DkYvTxImuVzpiPJcqEn6S10dsbQBx+I2LSLxoLAdda++bDm
KLo60kQYRF2YTZcm0TEoGEWmwuovujzH770e5IkP3PivYI4E2lveKUXTxA0XnY9j
hRUalNuCA9Xe93wu6TuUo/HIYsFgRD3z9T/pVCbKrLx0xuXMGNCKr3A8PlzkWmMe
GIxdww1jeOlhWYlZPRObECGJVQYJDisZFZbvIatqo/mOAqK+0OGKm2mdUrvsf1FA
VHkTTwgeFlNoSv07nTd6V1/DI1RKC0bgJeh6rn8Ly+HQyITVNnFlO1fvPDSHOADU
77LdClcoAwwM79rpzKUNiZMQGks6wEFzviaoZD2uf/41v2zR72MABBcT/YRxhBNa
zq08dyI+OLaxjYqewz9yz+Z84B81YSKIov1DPLQHj4LrCWT2YcoIBVwuaH6jM5uS
xS1/p+aNJlLOYrzklbdCF0JVLHSe8dU19n/kvSxLMEZKMJTwI7zD2i/hn+BH5boi
p4JtuptxKQuX/B+JDsc7t0MHarXzQ87IswZuhlQMLJzglu1ZI0uwViEQ+qE0MdBL
+cbfE1SAwTIlXMnrpANDFB57sMP/i8bJlg2N/kRkoOTgVkoksOX/Z5A6BNx2NTz1
5CPFUAJVlG4198oQ2tiv2I1SU1heqBbHVHM5Lz4WplcEnI6tXlbSGjjH3pmynsbi
oLC/jP0pyFXqekMSiixZ3K6crBK39Xo8MCPdkz/iCwTjRe1BLguO97p+wwkMS7hr
mOUqLgDeCHu+31RjeIcHaeKtCNytnp6OzLlMBF6JBgE6e1j3vh3pEHSkYJ5CrNdL
6TznXL5AZTyq5NAaQREKqYDy2E7oR+c/oETkQCfs5a40vp2DtPAUHKM8Vlegqpul
BIkbYSf1ivQjRKEmuHvItTkRoNcvExASKY1Y8xtlGawN+8HiPzYZ8513ObDw90v7
pOXHVEDsZ2pXrR+1atJPcDlOxacoZxFGcXiIZeUqN7QIJqS6DGKQpKIwt0fNSZXz
ORn8qAvyzxL/VRKtTKq71sUdBLurTD9G1WxmVe/5K946kPVsNExQKn0EEKJdMPeR
H1LnBiq7iObazP+5QRgoBPGvKGBogfu6GChQur3+7lwqSYRwBGZOWPPq7EgLJSfO
M3HyZJtqk0pV1oQq4MHGblZDCbjBT6AVr3ZAm5oYUjvWmKmEHTuJJ/pqtnDjnb2r
YIS+hFcDIG9dAeR6t8MTLNLvxZQan2HBJplQsTJCVXNhKwzHCaNqKyRltCpypwJh
isNlAUtt5Mo58zupVG4pj8dGjRciF1ECCfAATJWjcBFLSniN66l3M9aAWOBSGgUa
F5hZEafWHiohLaOFyX8HizAseJ+Sq9Cpbh18H1fZNzW8q+LR/G/OtUPJFq4KL+Az
OBv9LCh7YEuDohF7Wcm0eI8voCMRxNf8Nz6RJl2u/yrBripDnnI2peuulof7A3tI
uYbEN2YlT/T+91hLiVQBJUN7yShIekovRsdo4dUQ10XcyTsLu7EnEEv1khpq2gYt
+kk4Bc93awJ/Pt9OerfO+VAdUzSITh5hCQinVpRtIjZJ2oYE/dsYFcmHHYQoi4KD
nYmgP2JxYjaHSjb33I+t2KvbIfPDnv2w8kFNHiO0+3DDJ73wpOc6fj0Wju/kT0GJ
GeRlGywWeOZYADTqUYHnvHEux+CWOshhXKHzefTtO4Nwhzbi7fCDxeQGfLcvFMSV
kBUVjTCVC5T4W0oeI2s90dUnXc+FDoeJhvSsk5WgK/lNS80rdRORum4SRGZ7Z7jT
ook9YJDUaoIOhiyyek9UMxLTz7pLfGZbcghhVi7FUEVPCm8IyK7mfJHI1X8zQiDE
JjFZzUZqhAno+d0jB+8S5rZmBLgb9X0zmo+RHq1qeJenKCld3GdY/wo4KofJmcCJ
9PyfTpMQbCEQfzMQJ2uOOcNpxjBJoCQyOdjkDJZ2SrPR8MnbDjhr8ZGU5s76L0Dl
BSKYQf9eeKuTMcI3DWhCeX2iRhFdCHTWouiqIMhN5CKSgJ7G26GOwAa34zDwR9pd
tywsD8wE6l/ivzlfGurkPGHecgaZApPerEQlbwHhvjCg20g3BA4Lrqv4Mc+USzUw
Q8PiJmAclo7hBcrJ8i7nI79kjT+pfSkP+C6N2eRMWb+3sKy1HjKlBZazHdPtVjZL
aDlIYmUOz4y6MVYONFN1Ge9a4SFJcvtSaO6SB4A+Z7vZnkWsKRkmPQWy+0iyHbl8
J4kG4uH6l5ihOUuEsijMGxOuc3T4pA81C9iZe1vJrS4jGF6IF3+kaS/F2nqJUB2w
Vo5NrjkdBYkuMn3GT/f6zhIbSLOVHEeH31oE4ANt69SfyUo2Uq/2ifuDbcohuwJ9
6euaUoSd5rQtK/yKtsiUP2/DID5xl0Ksy+nvb0FDRm64w4HGeIYkV2dppvrJDX91
0kbnZ5kJpZIMOtwlg9GtW3Qt6Hh6wd+ii/SIiwZQH1jLDe0/KzLjyZ8OgFx3fLUc
T875GgC9/1EP572d/68kLGHzG8kGzVUJeP0RM8JvGqTmVSqsBVFR5BNTOzUNjQTS
LXK210MLKBq75SPeBA4K7zWvpQ8oHM9l+iFgO+2DsVkshbbYlxOOlc1yG8sm/t1v
DhR6GPAtMjTIdVNGPhUM8ZlP6Qmyzj8i7rL+qbW00tVSkgkNTY3SAxeAfQugcrUv
F1oKlLk/nn+7tNBDTiSxyd6U5Gmn1Afth41U1E1enEDHzhxVpWnZvIjuqkYKgeVf
xCB8M5CaNHl3lL3XB9qI37rAFubpjqSeesb0wSDp88XOaC+SUt/gEmZGNSddVAV3
aJWMMKcHLD5cbxORffD2XaW+OcC6ASWQE6jxD2N+ucOsf91ZrdagGmz+12cArppH
iiTgAobzzcJqHLQKqiB9H+0n8VphLFUNzGaEVwnjjUd+u+8f+r3BKoHrXTNiA4Te
Od3Yck8ie+mLDar39tUTPp6jKBCcBjxYh0z3Ka/Tq9tdpRYrt/OLH25t4UIj7bRU
ucc8fEN5TDyAyGsddgRqljy06rQRlMii/OYYTB2lJ0UYdTLLFLwtbVkTIkIH6OwR
5Ab26mEdrDe1nqgb3ndqMO/NCP2Zrpfur6NuIDqokzvW0PFpaAG1lKHbvrAFEjsO
B9w/+VXBsTLjWIduYW2DyBCeDpPZZ6bF7SWVSA5Cb0xjzwoUPm78ZATzCtyMZ3Sf
1ghBXCz99ksmt6bN5q9eveEePi5qicphG7c+n6pdEOpRMhK3rsowtHAiKnfQeb/G
0CGXQ7WpVbZBio/Msqt2YnL7oxWoBhEaY8b4MVtIGoX9QHwYLbZuhRK9xMW0Xdcs
LDlmbHv7LPYZz0DWfX9js16KxQ6dyKc/BXqlo7cPUtFxPG0TJahLHG1CO2bZnjEF
Boy8e5HfAnNmro2Oz/CbyyNDO0/l0CbfVvLbsrMxAFv8DsGM+IWSPyGmbw/MgbkW
TpH/ZmcdVBcY4JtdMjCbzKqkuBjspE3T42da38gLUfTk4kigNC4oMYUfoZ4A5x4T
l78UwB/F4s0zKG90lNPAWS4yywtcIjqVQ+AnTFGMNpE9vpph8lkwpZ6uH2rQlK8w
prFRaHgBubtBMCXG4s+F4FdLLC/CDGPf07JTnfaVWeZFNJTF6UCWFJo8cL3AS8fB
RzTZDqwkbzZBBeOrXS0/R5GV9swTDjuRmQpZ46+NNXYTDDT8CInQu0FGPmf/oXWp
wAfqXxsDJcNaeWCJ56gVQfGblNU2NjipM1gXecKHg919PTvbzyVxOpbsSvkgsBnP
Vp9H3sBCoLU2MqG1B5Q5n+V5GgAiSHspCqx79n5mzDQ/kZNosENklk3eglGAa02i
4Fejm7jRLms7Z23ukcImor7atX8oyMz4SPQOi4WtSjF6UVYl9fGlfaPoOx2IsOtX
i/vRUyMUijYCh8tD/2LMskgNUOcfdb+2FZsl+xqEfY53SGTCajTdpUsa7AyTXCnP
M/W710im75g641O+N91sM8aRADrS/E/LlAjFrKw5qRCBibjUCEC/5d4qX0Q0oxy1
kbR/aRFEHwPz5KRxxQbhWf3n3GT6V52/TWa5cEhwc/kYPG1TkcBx9J7aa4gjYvHd
JS0lladRuZYF+jPRbdmTjSjV7XJT1K+JDyjtw4AQ0IP6/fdy499QDcCH3jKGZoEK
qOy8LPcAMMM/1e9wWluxbJjvxjtgd2Lt4DGedUqH7QJWYayXFUK6iEWcoXq/9EpY
ur6Av5+MzXm+MR8bMTqP/4TFTBc7fq9+Bn+ZF4jN78joK02VPMqC4QKMwryWdoLd
ZjR6i6yede8N1BC9Y6HZ6NrKEX4UnAqYV49j+PX8MupzjRHYdC7KnEK4dJPxl9MV
+lwRHEvU4xEGAUeoifNj3aDCn2yEjZL+/uJIV9gVC3/nixIx3jI6wWAD/9VXYgRs
xIKa1ZeaI2nLQu2C44d55kT108/6JnaH0YEuMHXOZ4MdnA2Qt4fTN25nzL3UReVY
dZ/5LzsvPhokafB8o0nmkNmkBdrpofcBd1UZdxj2c2x383oFxcs2zaRE9EQXsGeq
InboEbqIoxOBISHlW8KLN/gt9b6qtEu7D41+8PNSPUe6D4NIxzhKZVL3bJ7hChn5
pJ5GxA2rMFinvX0kRxqQzZHwyOHGW+deafeD2MjuBYnhEcjlAzC6bu+FOmlEQ/GK
Oy5gezuLWP12BuXv8YFHJmICD3h88AFxFayRwvcX4leTFyA2b+y4qpXG3VuKF44w
UWDCbYL0VSajRkhXcinndvzqOc9GmHhj0pAyZRggZy+orIBdn/iHfVH6UwFYJe4m
NQ4IzwQSCjJywNdxWsUXpc2B/VyY4e1VI1quGgR+GR019a8+9m3lE4R3O3OIUVDB
Z/pXol4E+iG2Oz02nEtjRGwYVMs4bcND8otKOnoReXK0SpEzGaPyZBrEhqMZMiSO
nfFLK1UmfAYSu96zYC2lr+KMZ061YVjjTGbAs6/hznzMh6Sp4vS7n91Ofu1UUPJd
EfK0kLiiOmvWZ6q4XXKU9ps2XcjPf4NfJYiPr81EOys+sIbirUPBL75fPLhquTqG
JUlHQlPTBlaTZBiYrTh4aJAJHg9XJjSo8y8fOXu60JmPD72yddI4Po/Ux2bxNJ/l
iWLu9hTAzZ3VD0dYXu6f6jXqJnFFZpBKdxICmLkN8tZ0H6T1iPOFaMDawvx+afu6
W4FdfZGhA9ves6Z3NUlOsD3pylxWxdHKIlr08OL95QKeJpj3RZfQApozTk7xL1te
/ku8SzZzp0fb552r74z1sius1A4cima/oRko6Bhd0+0oG8cXKKmYnD2eZSqbnBgX
ZaMSaFSr0h438JuNcxRNG4U7MjWwytNxucm43T+inMAlocVjycp9CfCjvMSyHN5L
rN7BO07vgZyJ5IvtdrVUg9fQxq0vB2wcaIRwhKkJGHnei7nMntcrIwUXm3GQaj84
HXeGHfOZ5nWDdyXqCrNZQXJ9DH4axyItdowKqAbBFIQQEUh4R7c4UnogXkYzc7er
iMC+GkJ4i26eE+TxjH/JEIA/KZgBpV5ttMHiHOdysFuhtrt+3TKAFpBf4Vd6ujF/
RDllKRdlUqANi/WOdPjODto+T2ArGSnECLPlJAeV3tuBA9N/0cQqN0MvBgUrQGeQ
UeuZ71P43tBVfYXweDFo3zLZWG7LZU0PG7o9t8NPjBXTs5D1SWU2XYNBmTu0WacM
sHO/3EdKrBpN8B0/jNjkA4sa9y6raNi8ZapquXKFyp+RroiPzcOdpiUM9trwBn5s
8Mxgc3qhDbMgR96mo55IKB+Iu3wEHNANguFODU1idPmj432jOq/M6obiC5WqjevR
CUS1093ehq5KeolCpdk1g1F14//oTrBtxQwYRf927/C3Axqtc37m1B8QzHq8n0HK
WNnNnEm8PvS5h+GKInomKyzV7IjoTJ1UD6CFtfjvZn3ORx2TtVRiFZcvvKH+M2rH
NRXdMk0yvIpekmWqqgTFtd5cd1e2pCuUiZ2sW8ZQzYY0WMWP2fMjF30b1bHI4T5g
bKZIXZ1JtnnIDNC5x0f2SWJxAea92SNuMc1DVvlyhnrIYvs7LrUAKouELvy1cW5M
mcZfKFg6K2lsQxgFH745iB0Wd9a/GpNo3pRjexEGX6RmIM2cL1RY6fZ0rTsNbSpf
mbN+QemoI2hxgKNKWbA1sDlofeD6nWOlcHb9gfKgW7SBlvv23EGHgfzPi2xCELjJ
R1c2u+WWp4BaY1OueXSWopSFuISOpd4AUGYfFE8hAutAd+1jF346We7JV+vIL3Y/
56rc5GOZF83VT53Y27bByD6Lxx9xgVB9zsOWKGpbpEwSst7kSP6XJJwipK8SkHML
ozHOd/o0fAfCX7hkyyJ1P8P4ymUJKd507U0kjWEcNAX28xAd035ERKbsROmZZWSz
9RpD7k+ed1rLP0WF+SIx3HJki3brFVUo+eA4s9CBN0i+iLp7IgBY7d234avIkxJQ
dbiHJQvqMwDGHsySHkjSf5BATO741WuR8RzzLMJ81KJn96UavWqGet/XRoT56tDm
Qp3DDuuqmvf02iFI8LVBGlJpnVadhwlpBJgR/wPRoe7MISLehCLAXYX7zCt9pR7u
WAWPIh4bNvV3QXulEdK6l+5k66pmaCAM9vj6xtlAJyTH5qX/euVAuaYFpMS816Ad
l5g/y/F1Ws/pNuwUSv/tl2n4sMvh45T/fl63so1enflmmPn5ky/wEN5UmHEt0p7n
iLsSFAJbQZRghc4T5MbuLLur6PDn/aeSZj/56kIaAw6QregmDgJW+aNxh0yvtX6k
gbw19cFKudU8Jkz1Hz2v3Sppdq4RvmQ/O8mN8njNzPCNH/wrfgWptOzaZ3x0IxeZ
FDt9VWWSbPb42A460N1jdcLpNz4w/o+5gESbviJ6SJdUwv/dHBYc2nFqf9v42lPW
qyWAqknlx0qrtEw2kCIuxxoUtyTJZXtSKazhtH5BLgxAoz6TCx7x1GVx9z3e/7uu
aCGhuyHzcx5CBlXz8QH4ujcOi+0PzWF5F+GQUoqdvtkEGZDWrDhqxqNE6TQqjEIp
WQH4OcVC7sIxJVUOqXseF9WwYtDGSsG1lan24qxnMH4OFA6mi6pwjWR0m/zVLip6
3sdMOfm14y0jwuyEg8dl6E6e51LhR6rVw44F5ZlV0hlEC4LCyRAgdUaITktOjSKY
7VImjJCF9HYg28H+80ycvmD4Jwpj+ktu5GPFEM27VTc58V0W3rost+cTIPnYuGjT
xj3NHl9AY5DhhdQqnhQoyN1PISh5KeS2o9nDvp1Eg5L5Yb+fEB/5bsywJY/EM7KC
WpPdmyiDVNPU5mx/eK5fsq/lYADiy8jl35jWSOC6adPq379pSl3+q6wrvv+gU3By
dWkdpHCJzNnr963qf3UtgiRq1UpwJDdJPkmK7nbxD2sYWsb2vZaAl9AiZdSvF0VT
BDVHR7Bfds0H0vYBUIdsgylTuTktHFrmGFD4GZdqNEE5DMAW6CLHuT2Skd5tnNBt
KPxPXflh8dBmtg2GPDELY4Rxr976+nvmmrhMqt2wq4sW1M+R0TMExd+a1sp7xdmB
3EvDCghC5BhCFtgX6voiL/Y0WxfdD5hzYe7i7nvHtO9ZrE2nFmjsMxwtCq8OO2KN
JwEV2XB+hoAY2RMsk9PBhQ003XVXBXKO5Nkacm2b7gqxg900UhgNa6D3VNKFwywY
619jMNCc7UnP/NgxxR304i+JV5Z07ylQRVVWdu2E0/9xgC2aIYT45UovQ82pmDC2
uP8QbBJmxcwyhsMWLqsdPXmhmZ4d7rMCCFcUafIi+4VTonM+akDt4Zr5e6R7QHVT
BosrFHQLtnGxH+s5kVQOf+YW3sbQ23asS2YKg7epY79zRub7af3IEXS3Z1590uWs
0tMepFJ5aN8LV7XWnStWQV1a2PGvPzzqmjizf1bEdDqs3ZOVb7fZXq76p8f4Wj/P
/H0CX0GsWPIMaXeKr/KVmwA2D1UhNcvR6IHMYnVnZCKURB08yVn3XxdcTkmvIr2T
/dN/vfn3x7wDSVQ/HBGcLKaI2ijZSIXGK+95BJPVsVUKYrforn8ZBovT6HJlupXl
SGYtNLP22fMNXOkgmP/Jipa7Mb2GuChBAOtcRLIK30BkIc1kchWFCuW9CnkicaJG
wtvIybIIHV/Wq8F9O6rsRAtdpj6pJlNAMiqSr9kc5QG5aC7qD9a20h5ObIn8b1TQ
5Hk0btxlKy/86wm3FrjEaOhFPQ99PvldpS41tPzLUvPq62GKihXiG/hS9e9jqDyL
+cf32OVvZM2h2iwHjhjaUwZCSyF5u46WKl5lQ9/axlYygZ/Qcchw+zeZGdUkolcY
GCNLVyY7zxOrBtM01FU1Ig3EPqlgm5f1+Dq69V5jgVrphC0s3XvN2l/zm1vsDbvb
H7OboqFS43FZfdQ6pu67EDtezEz+0pDb7Gm0MMxsimlaiGnxsvaZiCBEqAc82+1N
ISJh8RxY0iPZ1LPfb3RH9nDAwjymVhJLqk9CIVp2KAslQ8yOdGuYoirH8Gl8d5ml
vNh06Ndtk/eco3i7GCbvsTQvVaHBytbGj6g8ajHlP4yhi1iHUQWGwMpCtatDmlPO
rtnifxSJCmE5+ihC0YXHbpsEq8Hre61HtdGMsk8yKmdw34MN9L+VR3wckmqhoJyI
m/ZlAi95w0kkz61p5URvazyafAOufBxCtetDzAW2YT6teiwdmO/dsLP8gobmYUOd
IhkXRRn+p20xzdWFommv+/yoQ2LlquSpOa2OrcG/xM2+zmkobHtR/qO+3QnBKUjq
NLLfBRohpEZALEiWoW1ej6YOlBFAiGEmKjr7JVFF1eU1WActYDEL1+CW2NLCzxoF
JLn46KSfimYabkVUGri2b6s4rBx1wYOsaKH90MVPj1PCuYdlF3Zzq1IYlrmuB66n
4FPN8zJuoAcx+qP7XdECT9UcugmorwBLe+05msnrkNUQKjqxLyuji9gcysu4o2Nx
jDnLX462h0OiuJx5eFge7ybolG7hNO2pi0Viiy0CFcJw7EhGCbc0nfe6NeMyTQuc
284DrzcskEkMvbfm84Hh4JtLUCCpE5SnuhbDdFBavVc0TyLwoUbZPms2zyG0LNnP
7txBP5eXBeeoyofQ8xj2AR85B77QF2YH0wHT/oapZyVXHOPMM9bLvzyY9takCosy
2NdMKHpPphpnD+szwdUIg0smWt37Mx2AiDosJC6epSGl3JYRWLUEzSkKbf1i+hDe
SM1DhZ0W+oxTaqz6XkEaXAoYq8brSQ8QBwG32OoHTGLB7oNtw47roIgOhKPZ/PZ8
HJ9UzpbHYrZFbd2sSo9QnqZ85s1ndDf3dTIKdUQHybGUa1xxlX94BMtrIXIX7WeY
S+BQDTs6ppdvCtftrz3l9r1+8OPD8QKLzXIa0Ja8GqOahYgh5A2NZ2J8n847hCqq
P5zdFeAhTK08WUUovzQusNo0VH2BM9ffMfztpw9ZN9XuRBQmoycX/Rxdqyupehfa
02K3/YgfyG50v5A/V93sE3RGJ3/0oZHOQqtB3joJEGmi14rrhtadqVmyeM55Ai1R
U8GK+YqqaSX75gLyew8tYZmAFgCVSkINY8yW8+hXB3nCsP4cpdqZQ+tjZRmu9ene
DfTvEvctVHv52L5BpTjSLX8qkZQGo7vG+/sOE/hs1gK10ME6XRNJXL+2DGzLAG1P
4OQmmkcxj6ZDlTiXZQETU96blFM6rP5Drr/UKLqJeKx3GFCf5OWg3ygOcE5u3j12
6tRCzgqXu+iztB9wT0KV0ROJ7lvaoVZtIJ8f7M0vL0qjfCmjvjVzc2EN8Ak6IBQK
RI6MhzMk8mJXhTQb/fmsmIkWGrjOC4K8uaoZZKRJByGdKBMyCfcbU9lBHeh4uB03
Mncyd0FjmTTVZMl7abnXXf1RIXMPiWpFxyCXJu6n4NrJTt5Skdo1vefvMyJdCMCv
Sp0NyP6J8tcO+1I45NiDDQ40c61xBW3Jk+ASDK/GF7aOXr20A2JdyvPWBC4XuO2e
NkA0rvao4QfOXYCIuVA2taw+Jrcnz3ygCeAfK2oyJSaWYIClhWxMK0v9pZ5uHFhf
15KxtDVufnQ94KCaZi6taFlmfyb62wq2k/3An/yq9EecDjPSIrUWySaWF1jkymhW
wH5aGLOGxmuoIXhky7s+mxwFBQevyIoED/vxlaVeYTalB4hAvcY48Ua+qU+if6HY
AisquYSaHJNJNTh0cqUwGha6MslBQB3v4eSik70+3ErJNqqvlj0hLE9Iw6b5+c0G
KQwlvV7Id5o/d6ktbtcb4NhBwO1l63OVtHAG1DqMB8/uvk7idG4oLyVPDAuoVJlK
s79stizF8Ee/vEug//QddFhm/NZVGizO5a7fvb5W0+hU1FKmnuJj/sJo1TK2Ld19
PZ+kz7Enq1KnnZTmSYH0GXqaNFamwmdoa5tjUXzxszFIoSPY2QkVIEcIq77x1zxN
vV37fmgA2uZJjx0AZ+GEUPai1i35UqrVU1FzunpK+q/Whx85nxghABCD4LXjpXxs
v/E9Gb+5UJO8WvRH/FNdsM2wqICf6dsqZ9dO0Z9+flmLDwDUc2u/Fh5SpwBLZKRC
p6xKacao/P+f1Sd4+cDdRNRvwwtOXX2/Ds8uWFvilBB12cjOC5sHDJYaSo+2z8PM
cdghwy7MRHcp/IfhR2iykg8kFamfFtsLozlohsfFwZsWR6rDrX8Q0Gdye7bMaGlP
1m+umbcu+dqzIr5WPa/ilYjWGNY3sH8X1GjyhHDg1UhORPix6UVRlgPPd9zJVb7Q
2RLZOx1qmLDiSKBvJ8F8jJHzyLET/ufKC5mNsTYT4CLUjAFnwDzmqcmmGGmxaSFc
oO97dfVORGnotYsv40yEQWRQWiaa8ztr52ESaBxADFuzad3M9rPXkMXuW0U55C3i
8sbne2CL+kKAm7PUEUXk3W77lvtAh12gO7WUJWWOr4gPk/rxVudfwdTcXlaX+0BA
Y2ZXsHW2H3b+iqouczXv51C5YeODzx/ZrsHJoYdlLY51wsssQecSCftwmsXwoOPy
PNdgypMQvfR14TsYW5UG+CQtmqQFmF7WoSkvEgRPqINvDS/xic6O3DGSK7+hjyfT
GbWVTwdi2ieAEWVzrfzOVfV2d7UG1e/zjXWwbT4SJupzxFwEHLPXxs/4Wam2ywND
nt/1V20WG/yc2w+TxMw4/h3mHPQ1yde6q1f53nx+MbUsOfgwBL7Gv25g2A5mP6TQ
MXN+xNFUQ572C8yRhIPo4hRHrVHYBb1karEjdRDRWFfnJOa+TYaY4EyiJnlAxhaz
TZkqREtZkb1dJyBxlMXNIcSBEr3EPbDezJ5cGGSYPBGP4kq0VgVC/H/AqjuIcw9I
z1Q8TXwr/8iHCgRlp9PMe2Y0/3peK+xPveXM31NO5bggYTZs4eyAXdV5j2kVLxZ4
zHHckA4EBdhXReu9ethreC5FC4iYiFKszMo18WRzyrNqA7uTbJdVVIQgY+zKjtp0
QhD5pZZG+YUDPLtR929K32h3RT+PpZp65a7BoRApLLbCFNo+8UIlyHn253kv9pyP
kh/tAlrPcoqNWc9dLWuUBpHXIlnx0xi3mAV8IWL/w9Vah6TAlN0yVoglXsLmMxMT
VfjKeFxBdgUnihJmK/KL6y3ozuAoLnp9pLBUAosH6L4KTwc1HnKxjp9T3GLGHjDR
mXEu2oYMqc9SuFPNnl4DXZl7I44LEo4LLzJPJtWLwGSuJgbW5u2tqe/+BOlNEVFR
h+JkYR/FAl2dWBQuBX5N4u74Wx6/+/XZWxFsOwFBndBj34Dyl7+cqmsbcl7csUxV
B7UuzbjWXLOWPKkKjDsJaoda6s1Iebpg6U43J8xC8KQ/K3fltDo20Rnos6JvYeKS
m2N9AB6afcrVkvdyRPWfkCpPPzW1uyFffWjCWyIZxLSaAhHbwh+TYBMNEle1voxk
J1YIoRvfRyvooOLluWQLtVJenpZiETeIW7Q4TJ22EHvEmZ0/ninBj/z2ztmzgAGn
H6tP2lbG00Ye4V3Xn3QYdir4qrXPMiLW9b8syK34WfoEIRuC/EwdD0vfFv/XAU61
Zb5Dkj8xDtcP45IDT3O6EOOEQ0fDdAMuviAYQWHIBaw5SSRZ/GWt7V9InuwlNj5+
if8ydGjsLGh4aLVW7RWzxSKdyqF2TAHNs+KjRtA7FRnR/KtBvF1TPRFTeDnzXRi0
9NSS4ae1EL3PBLgPboqUcUPFiTe7Gote27vWnkUlNxFi7c97UJUvEiacNbtBlWHC
OOw2mRRn4vAmzeoaobTiUFhNnzk/NBgphXvlyRNNa/tt3UEKt5kHONTHAGYX0sZ9
CLCI5S0pVSEnEMdPJFKvEdJg5xDMWFE3+l+l2eFWb/dO5aw7XVedc8snXUCzYAEl
qfCnwOKRhDxc6N3WLRAp9Of8hX56E/NTZDOtRIUYaHxvU/1vHhuop4yQRyLKljaO
34Rw/8t1rGqATIzF7OiltvqIpaQpJX3ZpJ71l1BO2UrSloOsZelwtcKUtANzuVum
lkQ+dC7DE2Vnr+QBqKETKhCTOxGTwnjKU49s1zgMvtPGSQrc6dDf/3gMJYXOrZXl
Aiy0aiABBVkdNfvelX4N+5nX9mAo4GvQXExJ8RVQwIGP6FgQJpG0zEAcmw1fzBPC
XMtSHFsWCrW4g3Vkn+PkB/FSi8yFwtxZhfFtfRJ7xvOdHhsvSI8/VRUz72dtKnIq
tHGIhLTt9u54QOmWdghKt9Mi0ewLlXd3V/XXBBbV3IEXVLEylza5J5MmA1a/+f1q
7QcM/XVCzqPTd9JTkLfUaXYan2F/inFNLgF2Fb/iro5lQG2iw8F70CdzOe6pQ51S
sxqfFiGXNfp12/aONNvYwv0MXWc2qv3+43PCHF5x1Ly8u9oORS6c/X1Fs49H8igr
OYMRQfw9FpuMOd5mSAMP+tIZMyRsFszftiuM+T+Hb3VOg2dB67N7F3yi8ThOfo8b
VQiddvt3t+KGRg2gcnUQtMWHshdRTdIkrWoVDLXmdvwum3GmItdnJl0g0m0bcFBX
rR/lkF92lait3bm4GhtOMz0fs91epXovVCo2pv28psZgHB2Orj2L26qF2QB0LFpy
P8IXBL+ybTfffGo+vpsn8e21ZQFXDx11I/WsYhM1BYLE2IYmxKU7Uy+ZTQs3bY8I
kWmN+ra2+2d4Ksz3+A+Jl1d0CLYBNhANdIdo+yXw8BhutMy5d22+Ltdld7CJN15o
KyWxJTt91XeSjdfr26+f/MPFXZH2k/i+PQn4kYxy1t+ZZN9zPK5q4hWpcZw6Lk7T
oSamJeH4YWVskuRMbztivpb6MoBdEaySrRcy5tzgttya56OOk59d9S3FM+M68Juv
zBEJUuqiW0n4p6Zri99icqJS4lWmVtgzsL7KbQ9GJGEvDT+LclBAfrGUGw8RBr5+
xpMHJ+MjUAh+cW41FP8Xj0hvoaO74ZCmV10dnABrAcdqqsHnP2tcFLs+zxGmojVa
rqB894WGkAYSr9jfiebWhKONuFx75xUotvlRpbIbQro8NqcCrcw8YgGIH8LDmxYt
VU16CusDz0whm5TWJAdfEvnHrhcCk5Pew9/+toFXBm08ZyVF+TOwB6A+2LxMnDNd
tbYMdGfABevAl80BHfFDzTpAlnyc6un/C9udUwPSg7SDuQj2SdQcncwk1USDI32J
OD9f9RnWTGVUafiEs71hr5dDTMUjbGe7AoAutp2CZHKlfiQJkZ437wNWv5YUhAKU
3rT8e2bozSOevSFFT91bKK2GvfvjhwGOBhmc8GrP/cYnXRRa6Zzdh3v3Zclok5T+
/ZKPIUbm8xXDFUAVmYHOxh8uuMql16KZcZCnJ2Lew7/WeekTpDMqHM6Rp5QOMZ42
ZWrp8jhVGTq6SqtG13lZSA1w4N92jBEDiVyYwIKP1nLGDQOGXz/eePM3rbfz9Obt
J5510ij4Y7NYHGrgfW2i76LP3DDGn0YIyQJ7hhgYEZjhuzQYgOs3Zfo9xy90Xn5U
84XEpoEDv4PPBNem/XrMx76xQyREQDpn7MbHvhiNx/bTUM9A/bEVMYBKZ3FvfhYs
tpCiRsBUXvBwLIUWWW6wvwgQEa0YQ6/0Skt8UWI+TxdhaUcCd5kB+g4ohUd8RY4P
EdWPDv1/uNrW17HI6Z+TwUQF8xuixmNaI5XY1L2ww8YkdyNfgP9tDTkF4keEg4kZ
fAddorozBSHcq0+yKaTx+SQlXcDkz8fPYQptNUgw8JIpOG1KkBZp/G19W4JP8Xgc
MUi/97gpBBLxONrLNy6nkaFmmjkV31g8rbEXABngwtSxTdoSLr1d4LYLNU1E8XWC
qiYrvMStJIcF5X75pFBNgqBmAkbN4zFX4BYE3ksRPYzRyuc0wLSl5RrC6UhMs7f1
xP8+RxFU4fTwnFXAV/G7ejwHuvMenlm4wEReYr6bVNuyLn8uW1SPurgR9EAcqEHL
jMzZaurBeiv+NsXeZ7RLj/icbEyiSsSAL8QD1jb3XFl9eYxos4ZXEI6GoL/SrDYi
JtlWuNysf4R1M+btpDYcvfBjr3asOpLF3aium95ZdZVI5SJ3vcr8atNpI2Oy8KJt
ncDAARNVhcMResFdsaoIqclIQIWfBSRWsmX9hKXwhW6DSf9kjDgmxt4izN7P4ZTT
BDSfsScMz3OIRaESMmqN4s3F1eHuX0/zpQb/NQnVWVnnPR4A8psForu8opJ+xiP0
nPkVBGQ5jdhfdD98/tg7aC/Q6EzyriRPsgjxuny/vA9P2quwgL/jlgIHq/ttPOSn
6RyhdN5bJDwlj3orBf/EKwmle52tmVrW5e9ZT71s7Xjh9mPYodZST3FNijmWPE8Z
WADzZBlAKbJnwa+jzjwYrrm3G2dNNGuHNm7lOEPuDRZgO4P65f05XRc9D+c07KBb
ePPICnoy/A6dJ5FfC4jYgNujcvVYW9A57pb66rm2JF4+LjRsXJJVUgJTwSzumyxV
c13GtZokpfXXjQn8694OLnoDk1tiZatHlXEYmi4S+BlMlEmR3OyeZpjMIF1ydH/h
C1eAnGdpgJPwaYVZP939e6CcZskGrpKcusOJn3tk5waJchU0s0Tb3EN0x6tyrkqV
rCuxfSyhF20FUKIb9JgE9b3YFelQSozQTz4Ss27e4LMIl+CNWKUJE/ylb/opknEs
2gTdXJm+xgQRLcbZ6zMjHWruqi/NhdlxrnEMwG1mXdqI2z/GHmgAzXmzdbyCVAYD
H38JiW6/ImEKwDBTRS4ggdtxj9Me3SUAt4h0C4+WZmSWgFUeOiKOrUMkAorrMWug
9j++aCOuTDKV9htFlqEoqix+Vvvvtf/pxLzAMB3D2bqVwIe8QKaSWbFlOkVFIlIo
TixpjHy7u1IRcWa9DN6CRUhTrJFHSxC/x4ceb/1gqCfeL98blxpsJREt5E8frFDJ
U+iqOvxZy0CfiR0I433TqoCzOBLB4W0fql+/fRpXyyKr9nKs5ngoA3FuydJ1vMz8
9sRSFPjXJkCizgRZIyUWOOxgbDKZ/cpA7MmmcTQUUF1dYqRQnUlR15GySRS8vz6M
AIw9vYWEG5DqFjEw6/GhwvjCzqjQ/BRr9xN0UdlSEwbVnfRZsAgNeeNFQeqkUuO2
2vIPekvO4pXF64OlBfmhBeadwheJRUvjpK2INx+AVwkYNAU7YBQBm4n3MnHlNlH5
jRyYGdeovbPg7AZ7AtyHtwGq3IsaJmu59v+Opi+NmmtDYcXr0dYUi/lD3CzqCd2q
R6zogFrK0dTUq3F+6/4ZqvJTjUbQwL760TZGU14eNTIraQU+S+KGY3p5coUgmTL8
6T1xQOZ/AoRztprX7jAC0OsQ90HYyL1+wJDfP+x0bL9SRAE1fCgIGm4PStCNeK/I
RHpzwR+9pfQP9q4JHqOFBHHp5s8U4nqCMyXj4MkXTYw3SNd9o2N40nX1Ep9xjXiQ
isIhqvWjcN657YBXN55uAHANASpG4yBMlMmFNVmW4dYqpkkUJeZeSfPibUP2UCcE
tt62EFdOeVvyV8D5ZlT2KZK+4d782fH4BFnLMjHkTGsaWxEIHAt/OSan9N1YibTt
2dWz4mPRwQ572nA2QC03eXOPQQb4iZ/N5kMl61/7pjsSQYFJpdegHeeLiyxdyCXC
OBnx6oKK98Nrq+GQRiTA2Qsk0gXBMHH17W2R5r92QKa//P9PppouDdFgjaV25fad
rQWSpgHG4zr/oWs+yOUpY/z2KhB/uqrUhtiiCQrFAKVmt4HeUB3FZqq6twsKcy5r
Y3apKcO2CRLhJUpMKwf+j7edPPOEFvOLpJfdOlYajUZgkhHI9oN9yxT/68TcGjNI
169mJH69XrEaH2GqYruyeKA7ZpqnBn2NBrpRYl7QlvqgQTdi6TZQOUvDdq58ZcFJ
1RohlBZ/kTXqIYO2x1WAF5JXLPMCdon1KflHBf8N0bSMAAJsNeMuNGHkE+PgWTyd
rrYsNyYttayNlYKmp/cQmRBIjYq9rSEv2V9TpyZ6vYNk5oXx2EnUX0l4kpx6nip8
IcSUtNTiWZQdDhndpX83nto1MaMdNrSY9mmjSrK9a4tO25t/BjmW9E/2JIgWr6WX
V/f6DXnbayor1IVe+QhgGmgjUPmNLl4G8BjCdyia37MeBeQFI8y4VRBNhLFQhuWl
NX7kswtXCiwzms69p/SqTaagEoKxH6g2vmBDRWCJYRC9uyfGVUSO5gDhb1uCIEOU
KDjOIYafsy8kH7MxRg4AlyNZ9UEyORrKoCiOKm4Q6NoMyuRWap80MhSwASTIwBXc
MRo3KVGD1qGdfUqaLSqUqSJ4xillLT61EC1XxS+x7HAXfs1NicrqCGfKKWCLXS5A
q8BiVZOAuErBb6F5YVAG3z0l+W8u9A0hqWls3/Viav2n1QPQEKTJnd86AA+egew8
2AGKgl0OwkeNJuGk2+5UmiuaMV5xDG3DtzaDq3qG/fI01vezlsWfbS9UIPTda+p1
08Zdk8bUSzJmkANBdtYdSnk+T/r9kAuptS+Urezi6tia6K6n5Lc+B4uvts7MFi7Y
d5CE/Nj8hlsodZ6UQmz8Ugo2eR+RXOZnGKmmjOl/i4wJnZdqeKOR0zSeSrHGvFv4
o2D2USVg+NIhF2DcKzRzF69XKd76EGiBuQ0RfNHG7YJyctzjYvthjlUELAZvf5wl
89n0u+2W3P3gy1HxMvgh0IctoyNNvlCGNbQ7rka4baOozxdA4qbtcT4ClnuJO7ie
R8WBR3gv0ChU47/SsxJ3Acf/B9Dq+zhWd/GAHzAOkLkirVov67eV6vh3m5M3z1Sk
HWPnz5wnVuY259gZf/+Xvy4qzan6eOcY0RjWZzq6XHYLYjSoQRhuB9urEY6scTQG
ruK62F/vEbp5Rep0tXEy+NmUwamXCAy+7MwAn0aMZ+l3DtsQ3aMaeIhlA539Nh6i
ML1FaDY2lCf3RJg24JzB+xrqxH+FReasyoT1DErcU3WfBX/Lu9luqM0duaV+X0zl
Zb6rYVdVTKgKDoXsvw02f2/T3aqGnvv2NMG92Q1O042BXfP43k5BiXej1zjrENU8
Qonfu0MuCb6ZjDfUFrSDGV95vuqORs43YYtOWCTtEW+z51phwwTqQ5K4q9yRwy3J
9P/JuIC2BGxNI8cZIJuQvga0gxc8WsCdHR2p7M/hVSR8CRP4ETDzxmMerAnb94Sv
t935EI8Rc7coJHPUrQtr3P/HFxC6W0H1opMKR9oPH/FZb7aSHzRvRNfba4Q9Xa2+
/djjBApGTXt17IQrYWjgdw8CVt1V+eh2TXP5sQm2gRszpDMfI8Vtvoo8w1PTsC9K
4n+3HNgdW/Z6W0/BbPvvqfhYawtvwTngJw4w2/3860dRRx+DXk25PfsMyKnePVPK
ZEjQ52QtRGB07RpWWBQPiTo7dZw3C+ADa/b+gOihGGW+O/Kj17IYZ9jTk1H/bQn1
mUdtE/k86cd0c90xyoGBuwKHkarIMVFTIej/3EWOhJmp9n6sx+s5B3rOVcvBxi79
PANNrWIG0XSzLnFfl9usr0X8Jl7gWFudbUCNoX8qZqqEzylIjZt61q0L+eOhSVwO
o+Nw/204E6utRVQ6ItmfW8CFZfOf/sdXi2IL6BrWmILttuqA115d7VnMYrfj0xYd
37AwuVPGei4kAXCW0oRcr4UOImPmnyCEsd0IsTWBwP9IGLUhEUdZJOKzMDuzHqBe
W2cepByAKnNCToSZ303gUGUmUJ84Qc4ZIb9UBHGXlAsFQFtvWnPUD8t+Fm5DtAtc
M09xe9AunL7TGVqoM9zW+2H/dE4s7tjWYM8iCwLXZZhlpXxR07/dw7oOnHkU4kLV
pZyFcMni45ZZvcHk6ahN5kkDp/QTY1GCHcnnYx8cIJ4SIzCF7mcaj0c3/9sXqt6G
p0TzfHvEHAI+nUEQk2m1ohyxN8vL14H1wf4k0UH19ltKXl7AW9UNfKctclFHzeuw
L88uHPHQOKloRmfEVsfYR86SzdAVy6cr8rKdc8Qyy8M58GO/FctZoqBln07D9w+p
r3lEkCMA15BdIIhZw13C84omzC50tWemSyuFa87OlkA/hi2f7yiMeB0XSuZN1DzS
/HXB50PYx3Z2uj2ymGURUMxPJpOXylcxQviPZYarJmqSjxhS6IFQWKMid4vL8ZbK
blfUMRO5gQlaFpS6JC0MUWzS+QuzDDH7zpXOwV+G1XLjZyzMYNysKa7EOg6hazeo
jmMZiyakbSi1smjlSRDG1RmL2mOAtDt0VAgyE59zPZMjmhP0c4fwYsufXI+PYLEF
RRaMRqw9pDM/xHJvPaUGGoqfzWsQjsPjIK4gwC95c0KLNCsyWkb37fy8qkGfxUrA
8cVD/oHYwrov2AGCMFNlFOwTxisgs80649SCy+hqUWbjwT87fhLJbcwpAXjex2Ma
xwKsoPlZ0NsTCsCn8nmfYSNLCIYHLSuDPeSiU6Ti3y7LbcsWyJWg9cr4DQUw62CC
dT85gHBQQxX5QIZpx/GtxI2e7Ngd7WkFhuginWQX6e1HoeS7eeS01nnxMcWZIANk
t9OS2x6Hf2GcFVvhe+MjK54KGtu7YfrNCNmKz7szjMDxpubqdlCLtpBuMpD+nYL7
0Acrob6rO9WNoFwHcIJdoTrF32UilceWEfln219TpL+uD54Ct+Xyfs44jAJe1sMI
EsKPJ3wSU5ZtK/fCIsqJyhqSbF/eMCY2QiSbPtSFFeCKNE15becbDeYYsMc4BeVx
l/3eGJLV22QINbtjd9d7GD1d9sQKDaZ/y21vexe7XWh3aNwyeFeiAHlxh+qBYapE
IAr8yDTOtQrcwhh3I5GTsymGWY/CCVywLddQ7jjqYKild4PF5pTaX5Rtj21BD+QR
FvN+jINRpGDel29VqGdhaWA9lU/jSSYINQS7ags4kLoABdxyrA1G9uBHuwLsCLgG
x7TTkZ1QLRtcyuZHUxwDr5eHa8TOSUe66eSHEoxs+jHTafVp2u8ZclNZas3IXHTW
DrmUPA1LcBte/0Ykl0A5Zevgp/VbNnWvufj1DPX+2yjaxe8J5MMjLKwa9UkQ+OVD
I7wR7w2HYSrUwVSOd/TZaEePVRmARbDAQI87u3Zz7UFql7FqJoPrD8yUNPqoneEk
0dkcNhxCp7tuQz/1NZGDL24rOkZmE72uIMrBRIDDpZl2TVeycdp4dpSzhtv9nhfu
396diWPbGzj/z4l/Y3TZigVzTByDS4ZSx2QMluaRojxg3zc/JnWTt9VpXrajeBHi
KwwvuS6F65nuUWg1xF68mjSuQ2WvfYUcODO5vfhmaxWYXfl0Pt5KcNXp7OPjcsEf
hsooT9wXPUoe9sH8BFuv9VorR/Hsox6U0Qkz5bXXYuHKEOjoX7hHBAX1zdTsDsLN
4IniC27nJHu0zythS8OsqNtSVN4ereMBM0nE4pHQYukWuW1twCI9nVjiDamj9VLt
G4GlQI765bytXmc3M5uqxLB+b/1I3mUIebeCNO50zYklkhL+mBEZh/JSQLnzCcVh
X8PEnnR33JuWcen2JKCw4Y4dIqZUoxYoRmNn2JtSDztqXbUMQfgaAWw2qe4QEPY8
5anufEhxRPdtWtyBZi12yjcxqBagR8KGc4FHiLim2bGgLMqSxBFa4Oq9wKWnZ0Ml
XsdDcj36CwoRg5IYsl2Qt8+eX5JFFLauf8dill1kH5dLnC5mAmxpuT28iGoDCFKY
yjiusnblKOOrPvKdg1kUYQEChKBeR/L02A5iY5F4xJ+hw2Yxdw6EqvBexiT0BBPF
BlUJb+wnhHD5SohAJXIE7zOcfhgr/hglxFRbqShW5J5tqGm9KvjrB6n5+Zana945
nsRlY2r4kBdZIpEjqfGO2YdboUOevwaAWqqA55ShEYp7fWE+CTbzw/E/bPhSVAna
6bkSVk3i7N6tKat28aITOnl0so9ZVHjA+qV/EJ02kKsokP18ER78/hUm5VDoRL4y
siGNFMVRoyeIHty3zql4gHMd399+z2XKghtO+pdiw55hGagw2adKUH1c4JXUnzcB
C8kZFa7jiBIzp74N2SluU2vGBN5I5ALTJ+eosQLfPkJEPnWSVoYhX2ms76mbT5X1
7DSnTl5VcHei9T3rNh3lMjaPfY2lq/B2ni4qCArIxkJFHOPe5QQ1uh26HKDDDJn9
5xKnrAMDbT0800v6h776Rim0hXl/HwJF3pCzrm53CCo1L8ocEcuULASCtPSehEiR
1zD9em0grU6v89hTdUuapnF30aYLvRFWVsrUNk5Cq6SV1uOWxoQPdhoLeQe8Ms7/
O6p+3iy5m4zA7ZkHOvSG926J/O4CkEJYLWajll+hSgBPVAE1CL7WIkqIIQa32YmU
muLPled9Z7mb5OBLwApADnilDQIBAJor5KY+nvYFMTdByBNMR55pKIQaCWMCdMfA
Jca5e/kHy/TPjfB8Y9kZlEGgUxKhrr4q4jvi8SmbYV6a4cfM7hcRvUQ1uiL7y2SD
O7VtzDrXy+gPan8B9EmrxlPjBPfVsK7t2LUIF8Q/4xVOPs4OksAAXapL6M90/d/Z
NoQkBPBzw2kjgWKtOzqd9FTsd4PJD48QCeX379jSjpJ/T7Uf1vlIz1FMslDYeboE
ylAboFEtqpADQRbBlZnkgCxWDmJnQwpnDIs3UBluCN7U7GGZSDB33E1/kkghAaqA
DeJQW/bOFqNu6lqg6dJM4wGEuwOhCqFcbvADgqBHAndgURtanWT7fBssuBSkKjq+
LoKTWcznM37D7YLTJoQvdl8ohkXdth4/l8KlLStRkRgsbJf5kKZtUg8hZ2ybr92P
MJolNwhc18iZwFiFljNo7GAVTqWKfS6qOuGvFMg1U/2A2ulyJ4NfowpJBYomvVDY
Swhwi8iG5KAK1zWj3KVyKsj98+VdEBUNH+xcf4Aqjf57Qy8teTYl4cOgQkl3hyJn
WLO0TdQjzoMLKVKJrfdk2iylJ1A/Hm7xtGe2U5MS3HLknFkjznwvdiUpc7gnNB+s
WlsU1jl8UY7d0+r8SVd7vTS6hRyxlIswWbfcBkO46wBLB5cN2XyuPssQIV8Qfnow
EZYwG9uGaGFa+PvIrAm6/HgerJZwTMUM+4Avtfs5ckwVtd3gV8Cn+0FW+GLsym16
ldAVE9afPVyHedtrc2YnKA8MI8uZttggPEnwWiGMKZge38rC4L3RjWEvqy6UPzoC
fHVe+Jz1AgxK844uZ63NPdY2RG3B4rU7Bao9T5oloIUh16MaCN0FroLfwdDSXnBy
f8q8iZBdFGH8WgydwBmsJ74lLtKwHYjqZaAJAoEdbvX756GmLoGYf0qWlu+GyKrC
wGFMHeodRF73B8EGPgwlwV2x1BmgTERxAXeA0kR+lAEA7zR7/zvioyuXI4UqzKnz
jTWzhFsL9mA03ZCUd1orqUEohYUGrwiU86quqk1QNMjP3pAIpLc7k0faOgVc81VU
VF4ucq2CmH3SQT0NeVCJHce/9h25wIqdqy8/3x/j3/rUCQdGBLyMjhx/d5qgntsz
tqDSREwrt2pMPaF57mOiz04WUApnTY+afwTn9rD68sMU//rpYFbGH47wxdjPaI+r
ZrOMqow6HNlnTSfRmjk2BlChfOj5OG9lGEiyk/n7CdlgoeZfylYBwqx7of9++oR7
25a/D7buYowY0I8WSaCQHC9DyRzQTfpet/A7ZxaaEVg4blnNysG9ik/y289HnTqX
3e/f3C2ptHa6Rb+5GiFhwd+Rernv1WzRIZ0mvZBuuRpe02Mf5LGbeoLYJf2wvGKr
zY9rQO31PVfZs+MS/WNlCwgfW37GtOYw1WQR5iS+wXu5VqZEEb8/eyHBw6VsGEqN
LmbUQMGDh5XMKhOaiLdc4BGLlKE29/s9nLrhi6cYy+ddGzIimcBYMVAmbPnK48ZJ
DfTQyvmmHbOfPEgdOm2VzTKoYGhdOvK/Nh9y3RZaI3ch449iq6t/12OHLB8mwdJK
2jcJivbLSPc810eYgbJzziTm4o1thDIDhf5rIYUx8RDH1nlczuDwCTutD9sMtOSB
uIEOvGdu+uadhlJxJCAbSYmnGXhr50kMMfhNgb/aZkm2qkgl2hQG0LS8VyQuQ7Qi
cZ2RozV9hQMEOjE6vf29jZK8Y8/9GLqNliXoraZA5HyBLdA5QKoRB4RgoYmIWGtz
cUWD5v9hLNZKdS6pEQki4CYqNVBPYqlG1xc1MYMfcJdvnPwrEFylLqqa4MLke6wg
saMCNCdlmvR2FsXXJmRvoRtD7C78cD0kNI0kuZhcK4od+hshXHXgD5WXWddJmoE1
8IXfdlFY3TfjUPru8JqpIJ3OxNgjS1q/8TGj59BOUqTx8kdFPDaa6/bEDsS6/CKS
OM7HfXNrjniXJ3CWf1dYD6rlM03EBsv7F1NRZhjZLbvYywFtppajIqSq9UVc/R2l
VG5Ga4nJllLxF5hnp/LM28djrCTUmmbOrd5Mu/VMCwn5oTsE6BbjBJwGtvthivRJ
2cyeuSW7VGMJ/JpGN1hd6JHvz3C3WOFoWH1zJbUTcN74NJBi3GKGGNrx5rioxaEC
98TGThIfkbjWTTR0vMenvt/M4zooibyUiv4WgPm34Nqz7nVbNmVhHE9nY5QDj1+7
7IficmXJusgFZQELfmavPew5oz54aYbLjE7930bkKao66QmpKIUcWtN3YkcF/rwu
4ecT655tNnmTg2hSZVODFdYwOjDB171uktRdTXBxrJWcvEEt25eqEyizHRzQBJPH
F4MLbgmwaYmuw9WZTlPpzCcwwOBS4TnGcgLsBZXCQ/nd3tHgDKSKlTUyMPQoLVWw
lyovcf0wfmlJNbjKe8jSqD+u7J8XGrIH3wk9V6f6SHEjOag74Be2V4HTsov+0jGu
2NsFmqbEQIT1BfK+KDk/STbqG2dBRSCg4crAqbaVreWr6jzblCKmat9A/F7nsC7q
PNS4a3AJglZ8I/TC+I5pfMeYavYDPNmARonR53eygKJ/twxkmkBhS1yIFH7S8Quk
ug1iU3w6ZbLPQdS4lf92T9OOBNjbIUD4wBFDm6i7JqMhILNsQA3B8rtJf8qIvOQB
uXVIg8TbpGInQ9D+1nr53Y5Wiyleazcphnb6uqTAFHlPQqbJCxP9Ne+H2zUSgVXT
Xxk5C31lzRzwvncBMAg4TUIZwhHJa50U9oo584HNsjnGhuVgkaj2b1pvaf4jpvKw
s2uXovRfmEdxMQTSdtD/nQbVkDNg5+wkoWUcxdYbQK2vSk5BihSRpKw+QFopUw6+
gJsE9O+GvB3OtYyQpW5q6lQg6+PnJ2sfL0ZA8dOjib9kuJ7LXesdwYuUvBsz5YOn
HGQ2okzRiV05w6XCilIy2nQuvbVWHmpkjeRNwe8XaRTZTyiG0UnXyIu+25CQY73m
9YmpzAvj4gODvckvl/kviRLuXrgQ3EPBo42BBcNbwPsHo4hnF+iGuj5+ePMmov4Y
k2pDgG5haJo896SSm5sxSMqtOVCN/3LCz8EaKl9El5OuusqYYnPvSqx6gZjwbRB3
QLocO5zdqhcT5SMOV80jDsxOWzd/X4S3B/uKOeyPFOZXu/ZxZBNYcA0+jnDmQGh8
ur6dq+tfRduAOSHBbYd/jMJ7RuorJryZ/p/Pv1AEZW8dlzTeiJNNxtmH+pDvuN1L
NErBkO3gbL+A27KEH4LBSmOMeiPA7lOSg/JkjMcSe8LFAa4rZjmr7uVUbX0mJ4px
rBJTiSO/drSyBpMKeSvGDxiLACtTftFH1d17jSume8paSEmEl82QUZ1AtANvZTN0
Xs1GT1eaKyj9BGlHWakjzRy9QkRGHDn7WaLFSNCxmC++MHTR2mC6yWtaWvav6WLW
5b/NLN+m0EOBa203ICOWANIPCIbBq6+99XQvJe7JyzMkTcEVhXDkgvOnMj5FxxyW
oHEtt0dqa9RGwwp/Rn/ognmKdssLaWf/u8ObMtWzFObLVWXRKYvK+UMHimt87Y3u
oD1+koVOTnorz32DG+20griNeMqQFETY9qO9EfaH35Kh9nup6XrrwKQQZNkk/x7S
HKswBMWm48bxMwVsP+MPghpRqJut9oB1mk6bFdvq/NDZ1rbUreB4zIYbZsjhtvSM
5z50sx3wU20ptEyjlFZrSSRIpP0VBf0kWB8mbLZ9+zNg6j/oMstEoXWEw/aS5V74
fhxK9aR1P/wp6lMw1rIGv3Up6wCpGi6djw9YxJLBzhGDMZiGPhnfM1yupGRWPS+p
j/2X/KjZq1Bl+LYZrHJfEVciHvKnGhQ8KilyMSnpktHOTwAezrcLNlf4Sx6h8kdR
gdcQE8SNt95svZ2mZ6hz5SkGLz7GytKrtBQwgKWNp8c8L4Ci+82n4Cpq0zSyExl8
ViAukS4YCvH42EAV5wI7RbXGOzrkUbdImzdiKb54busRxNzq3eRnz5qWpQzgghCi
VemjqxGjRCzmSnvH64cvfEe2zql8fe/3cx2us/wEy7LMmAr1lrjJPUps06vpUfQO
3VEF5LbAVpSSre0qkR3pddrWpCTF+dIeBQr/3qiwmSSaQueiNMpcyqUicfLvm0k4
0oljkDzbjMdjl20pic85OFk1/SywPZpaV50RQDw2K+O/uxLmZRdtt6e2RT9kI+5G
VxcytJ0Om18i+9JfiErq7G7pO11ej/kM09K/MnZ9xgYD3XD2mxYaUJ/KMGFFC3/U
IZRCWXgo2ps1rvjpVTIM/NuIwuBu/joruou3ZDYtBRkdDoVkOOR1YlWo9EkAKW/w
4byiTeI1nEfbTxrHWIDCDS+6cKpTuHlwmSRTdp5lAqG1lCTr7vl8oE7IuMCllMlC
uWgau4IOH/xZB5pA7TS6LJPbGupHsj3d7kT9Wyxu/ywtNhPiXhEVoF5tl9s05NI5
X/XfTngEFMBvwAsEWk0NTMH/YCysXpBOwA/5s9xWg41PLSykcK1nIFv2t+wFpUVr
sZHVX1uEGCG29NzIZXR/LxOu/X5xejeD7/IJbSw41K+eiesjbQbqE91TK6m4Lcma
SSLtoDFd+BfaqnLJQ0odokJSmIxaMPC5cmBGiRyfyCjc2qe+JK9KVUT41qulgIcd
NESC4y1ePk+TvzANXReQB3+iBOZJGMVNzYuKGEcukFmEcOGzdw5A/K4Q5KuJ37y+
/iOQ98vjfDrFzrg9hXa4d/t754SPNpeV8PyRNw7K7pH4L/i+8S+WgTwL766C9Wfk
/oX5eoz4aAO5BVfKD7WVbPG/kXl62OV4dVHb342f+9/RmfoUm7uJBkoO/n1j5NWc
yWI4joMmmqCUydo1QQ3YBSfrA3u6eW6kKhcN7o6jxqaLx3UakgmptJMRlUK5rpF/
UnDMJvHIgcfa9jFRP0bOH8lRr5hIw735L1+56obywPZnl8sPGGCSoL7gnyjXmAiB
shBKQq/FsXwYMCZvtIb0KNKPAHzhZfcejSLzU5ck83TBFsZP5tq5S0EQ6vr4sw7i
e/au6DgbcoyFiSgELDEX0hbjt+xMo8EQTqERWqNuEYvKMoPdpP7tozTxS1DWsUS5
uqw4eQ1I278Gl4jETr15oWX1PorEQKdAAM6vWlnnsoidgYOtVCaSJgHYIhD0ReFW
WU6sXUcoNrp4iHvZwMd7fblN8BUWftNZy3APHVFEHMk/EW0fdVpQSlUT5VKtuW0y
lKtd8KsM3xL1i1Fgqn84mBjwWcd6Dx11/Wy5K0TTJ40Grn2akd+boOaj7unPSVoT
LNv+RZiTjusHqGJJak2h9RLfeMQ/hiosAubNlMYzmuEsDAF6f1bSPzyRVaQXDj1N
suBC8YQ+9dZuY5ygB/jG7xiNJVZUxlsTeRtIDDr7RzlmnzxuFMnAjQEPDZikGdTC
YOwHo1EVg1wnmPkwqBYcNFAx8nm6Ixvx6dCcbWxESyn6V3cboiVHytssm06kgtTO
r5fljcDksSQRCCzT9/qZZV4ooM2rAyE0wAiM68Ly3OG/+DeWF5pWjAXUVYQ2v8i3
HDXo/CRVs9kNY9XY+Vw6FirEesfcmDmH+Le4XSs49a08Vk4d17F8ZXnYV/et3Ywq
oYPsIcJB+a7nLg/PRXzIbIBlBO4b1lhB1rgsqJ6MAD2vo4Q4dF9v8B9G/6QLmsYu
xvuB03QChFdeJej27FMpePtzkN051Sm1m3oL8mz3NHgMz8YacEat2qj2qjA1HC0P
olAvHVopCMpf9QW49toSSDlxCNiqF5yUcTea8nT2BGKEbIcrypnZWmlynwWiIYw8
GrdOk93NobBIrSyWqoNSvjszvnuYgVnSVbAzha+WI8asyCxwC8se9hIOtgbJb52u
IUqqHjalFzyi+8saeKbv4n6Pu+PLRLQoGs/vsTRJMxZXRz8R9jae8u+/4hkONZug
8Q9fJ/HwTmu7MJGgn/a+6/Z3Mry89DGAM1mM2NJ2YgV/AFibHpO8JKH1PJZttRIr
94AFr/juIT+VYgO9shYMaV/0JzhqmlD93qmea6/DLGvb2Fcj+Y7qRZdL1OfqBrbY
c/34h2I6aqJf6J1kR6/rOWY7DHW//+X+MDNsiQnyh9usJhHZtVDmfqISHiYTDkkp
Mb16iqIAxpAY7bOUDpqedK1vHtXRNydTvSx4hYY7r0LeRbnIhdnsuJhHGt2xk1qQ
1VZ4ZQ0iddSuNIlVxdxK7F2WGs16R5H24wCmpmzRS6UVwnNNnR797BEgFPwWFaCR
VWCD8y5NLG6EdjctA5qcpPh2GV6xqkAbiMY1tEtGBZQ4rAWTPOYkruXGOjXW6tBE
0gzDjIxZRvFqDV1pezV8iyUCcBa/H3rz0Q+qv/t5jwqqe1EOyoBXvluQCbtGkBQZ
X37IST4e/YEK6f2uT8u+SR32GPd3obxHtcILXuQhK7PH59zb318pwke6iRI0EnsP
j0Y3v7ASyguRv7Z1EL02Cqvb2NwtqGyaykmLOGVtGm8Y9oWQB2mVrkBRU16ZX+hB
znKi9MXv6NbbVZJk7AlE6HhDA9tF1Qp9GwEehwm4yJGHJHUzsbMA1sJEssXuCZ2K
fswVxDjjt/yZC0U21i/bNLKWDYcMMXv/+B0nAMcu2sSx5TzkCJgI5016r7K7yRLy
Sgd8qQFUZ6O5CF8e9Zx6PdpVnA4aqrusZne7ySAg9mtZFg3134X3bZE5KGkYoUN4
JMqHZdS2uW8SXtVL4r0Ev+QPHGjAl3PKY9X+hJVcG8GBhs3KUdr6V/MMMg2bXpMA
J/dzmaw0RiThlM5NzHbs6KJXEyAmvZHZvz3Fk83uLPslZaL3YhqBFUn6qA9Gl6N9
8/Z1beJ8N9elpJHz6nfzUDSf0JaiF1Su348/SEqtwRhIESdXWM5zswigWIqH6X99
fYigSPXZgYcAASSjqZz3+n8P1iqMt5dNTJwF2SoxByfEpxCbc/LneEp0yS3gLbqW
00fcGK660PlEuLMzcdbTjycH0I9mhKWhOQD3zY2RyY0ZP2elFF5CAjVF7nrBaG/1
0OWn44Q5LVFHCeV1Q5jOxm7HIGWTJRjCc3pcTAqGwmkCk1ScNc5/8+SAZg+Yj0Bd
2I5/x0bXyLWoZ46r2igGY5JvojkpBx71zWvRSYCcHxvVY+itL3VVGCnluVr1E9QQ
IUlzEBSPBO8zOoD7qFj5O6xlJlJ/a1qaT9rxL0+ygXnVcOYVb4qb6XSTA7/0rm4l
fGoPUmQCO09zftlajuY2kRgaM4ksD6v8inkpkAu8C7t4bkxE+/PlD1OfAFNXLV+T
kL+Yhi/diTlw6L0vJmrQZgnWPuUtN6OBnxjC0Ik+Euwm5E1SKlT2aeVW0woyCXsv
8QJUl3FOQCb7SZTGa2yGprchbffjomQpZh5YKL71iWwkVBuARPZ/s6hZlCowOJ5r
WBPlH35EcvRwJLepkthysIrYeoRfbZmBENJSkvwS5LrvojQjh4M3liQfHt+njzTt
TQRhDkLF9r/b/EBKREslJr6ddM4mbhTAZxVNURut2bFSehKTExRDFzWbn5B/P1+Q
BHScCjh7ZfVjnfbe3AF9Kkhq5lrIa3wuSkiKAEhy0G6gK1HimwSpdM88wxYtn/7Z
bMb+zjLadGCSJVdSKHJLTpE7ajnbfswyuUrja7Sh1m2NaB3nq1kZGit47u+GfSZ6
Qv2FHCma6DhSP3C+y7LjdPudL2yptQSvZ84/0MT3fc3vbL/Bcis7l8kyPiqRmgiY
qz2vfI1DcayQlIvuPXps1oOQ40YvJTS+85MSs62entueJto041BA7OK2OQOWIar0
tsxQQe2cK+PcD4qTzOpBK1Fkxd8+MOx6pmgKmTufr8kmZ3dnysfO5hWuClRZJbJU
2jjQNC4RRGUBwVjGHpoLkuku0uTL6H5zWmutZaw+ORXwZk/QHCeM+/rSlezH61IQ
iW7SYSKVX0fZnfJsHKYeqmdTWIkVhQ+M7YlSe8bAMHVQmWaOnFs7D8aMr9hHpz4u
6VIaNmzQ8Kw4Uw+/X2hvhDqVatbg2X+mmibtd4xvRJgCsB2Fb62HKtu2qHLkWcSP
ioHz6fGdAEoNqF1SdjcLj0HSdsmDL94BnqRVowdNyLAeTi3UahHUZ2SlRqLDa5oZ
hlFFFldMr7TEor8s5eTIASRjiADKcNkzCVefwX0NHhoazRsgqpxBKbxj0ugCHDkD
Gyd2HekejQAKfo55W9Y8xQe6af/D3eZ4RsbZiM2twzdEVy9rQbnawcc3bOvOXA/B
ees8oErnpVtNHtMh6UXKUDZq4sQ5ESJAcG8xgdpnI0TPi62lD+VCTUB+u6Jmp9Lu
lYb1wfXhkp5Wom9kY1L3JvTGKD1K1M7JKJTcMdV5eHLzAp6e/0g2FnBeRd9oeraq
JqiQdmB4dOWGl+uoAktuA2quGtMQfVHpEXqKbkb4jlYuV7YmmLX5YOrfF3o+08ya
BsiuDfixS5WKRdkpvOHquYAgB8hz6a8ZFTLg8QqgXsh0CbaICcneShgOsIXZ4Qdf
XStfey2uTQd7Tf2MXI4Ylp78vBzhLKWeSNib9dW/zFpyB84eGST4LyfVEMkpJceW
OhtZ8qH7VRaTErlB202EFVQyrVPSDJyDBlDbxNfyieQMEUUa6UQKHYKDOSauIGoK
zMmNDDmvQpWJgCBxAMWCtcvyiL5TytFalpHBKQ1g63Ucm5rG9THmuf39Gon2/3f0
BLBVBQLFVxTtGFJxrSc/p/s6NlfHmPoeU9UtHuq6AKV2mnyTVP5iySxTi0uqh190
uFv15UzQ5v6GMn7N7K9/6GbbSguzHd8EqK2py8BblOofLEvj2fynuThlToXdKx2a
gEEL4PweNpAiE1Ey9P+fL9PT8rTtRtH9c2rGP1eTLt6rzIwnOEbsW84larQcy60R
RBxI1W5EjNrjpQyjAbAN2sqZCkfY3SUropbzzIMk3awWqihMrwUmiV3TkdZ2O2hy
AIWnu7brpDrD93SWs5M2Lc45OoYFnvRTwlfW8S9paWSb4/0bSzRjR8+gLy6tXCpP
JFy2zNsKtwpRO7cMnnDDbkSDMvNw7EhXEbQjcQoAeMPz4tmrVmrPRdoOIn5RlTaW
b13MuHZXrKLV9pCWvh5KmECcJGlY3DhsDjA+n0n84gf5UIASz+4Jd8nOTYpnF622
go0dTAfg1wRY7F98m9f2O8yKgBG+n5IHhkr+ry8+w69Qa9YIp+a2idAXg6r3nA3V
5zPwinJyBy3xD4DuWtd0nmpvSUA355aZWTwZx6bs0CdAvsO/qKrt6LgRI6/1iQ+c
zU4eTC/eqMngrU/HUkLqCS2xq/vD/sro5QA7GK7c/PXOQosA5XevpeK6FG7yEI1H
1FqsQuF0yiIMLUSad6j7GA26MUX5mSFnMJ97W8HIzSChU4lnKkeHkc8Zp+fspM+p
Fdzbe4TqnjoktPPJJtnbQgXVgD/indrTdPmwp2hmR/hWHTcvNPb7BFc9AcjGUSRU
0xbbWsL0pB2tMkRplAUYRxMsxhWIuR8253FjTzXIrnGvRMiBncUQ6hIZGdJx8wLP
ErCGaHA1lahWT3buWE3u+5A2DuceBG1v5H4+BfnBd9ncgzHU32+UVeGy79HS8kxH
z4NJwQ46n0vIVPhyzYTQ0NHbHbCDED8KdDF3N2SFvVp+BDosezvphM2CHlce7Y2k
1fJc3oR83jzNUTxmGQRQWhjJ0tvKBucKbzg2B3fv4YOTOonp4EfQC3uIl9eCa3xa
T4ShDPLb5f7hzrVNiC2z0ae/d4Mf7pIG0OWZ+xF2LPMaffgNYbTyXSna+g9W9Qc1
t3ssx/QNaoT8Fqwmn3zYcnx162O7xtBachUmFiY2NNCrqh2vju4QcdsOfS2H8NsX
1wtpwi0MJ/dCaF6IteqdriM8QySaPij0jbobVyBaGalIhqPR6caowOyxjqb8/zUs
586za+pO6iBvBErtNVNXuXIMuWn6dQEXLgCzON1OhaCwF38ZB7/0bfQMlgu/RqfS
bdKPIHCKR6Y+y6Rzr69xmsivL82l9h9iiCO6tEhtGwtt0LWldvS/JzIi8I6tSJgx
QS2oBIqrO/8W2rK6CpUGXYQt0/+EoGnKQ0MgIAcF0ahTOZWNP0Ff/tZ+PG9pJ+P0
hSxEDm0AldlN2S9X8li0x4iPEwrCQPl+U/0z+RHIwx48pSSKF/Kfx4IF1Q9pI1/E
LCwtSSyPQrf6oPugpLtefosNqutqzjAD6yR1YaUpUPe+/zG+zbEmhh4XOK86gLu6
PLok2nD/VIR/7a2JQ0BAjk5UF1g+mPv/756/2rfpEYCdgV2EJBaLJgW/EJEiqcP3
iV4pwMR8k5UkvL+hXqtzikUGYXjzZgZSuoeL3WaW0caGz3nhA7+98J6p0Qn9KBSi
mgkrH764OZKycV+sZpFAcLCS91E5BCyK78jjGTUdzRTn5hbgBu438hZbGQZv9IB1
9dGmLumSC4h1f7hok4qlwCLGYcV0obIzPZ0XsIS/555/etwVUWsFYSuOKpu3Zv17
aVW9P9cw55EwKZunBwfDhQRau8SjYCqHf1NttIdA4N9CulkrdFf3hwGq5xxOqxdj
RcN2yGKvDolcpGRqvhaZ9Mxq8ynO5QpGUUNu8bksddSpeQfmlhFuhZae5vXiEiig
g2uS0uIp9Z/cm7WCTFYNeVwlczCbsMsmwbrIGRfRkUl9N67Bhn+8PX9NWYmV5a+z
SDW3ZUgfRSIJ50mqpKNlQjVWXHr3+qs5iNftRw9kTVpN1vwNUCXVFttso3xOXIex
c1SPgVWdAnPmcCD+haFzIX0nG1cW5gxpyiZwo3QIgKDxmxSWYVNRcQU7SmiuPMRQ
6pw/VjG46bZSAfb5mmWjLsdnsPgfEMhRnRDA2muUi3Ka0e0p2fYUjFQWy3aXVweG
5rpNe3+0qsfHzmlZckPtMgbh031uPeXxkJGD0Vmobjc6c/aN0lWvaQUM5BoYfMau
LQeY0Cbl4IreL5/yxbDHEhP/1PUnG/Cp9WOrn8s73LkfMLwJEcXUFrzc2czvDW1l
2+3ayf8L7+raiP3srl8UJuJfomAvRfz+7Smk0UmqSrkl4WY09mWxJPVAiRve4N93
Roh/Rc2pmpRtGLOIfgkWLmB9O+bfiG5GcELFnZ83Kr3WyUuizHPNzpc9H2N8saLX
3ssnq5jhB6dKJGG987WFbQThMfHScizIYFyfgt2UDrnz/WSohQegDn/PCPRlHcBY
QZPMDUMkE13SHT5Ho/Nq0cYMP11Z4xQRBqGoLpCyDsTLAF0p1b9JWI3xOCOrVFJo
edn94Fp/AMq+hFrwQ/vIB6/6qI3Alz/aBPTbeC8dB9OXlCPyDmMYhKwNyG0CI36d
efu0jLvuWfK2Hz5+CUFcjLKzlkOm0+qTBZWRYzdlNC86Hmh2yV5f6FlxjOfvBmMI
o0GmwtqKmEpl8GItteglAff2aCCa36bH3Lwpm8WsYffvnt/3OXLfGO/ZnKiGDg9H
1Ecgeyf/S6CzSTmQ3PqC/HG1QLflwAMgr8e6LaBRtxPZFxm+qbcaqmU0w9Koo2m5
ROzXO890k04a3oV19ym8JB3Q2Eujlozoehxh7pBSok7ugEwic/2QEWw9pRjMsp3T
m2eTDHSqkK98/RsGj6m2NULle+98xLuUP+tCMZTBCfwmoFZUs9oj80uRVXC7LChK
Y7aEC/ONnIaHhdyMu+khjXrAlc9nKGKx4aQMEILYTkI2BkHG0QWd6t7nyVWIC7H/
iDN7SvE1kf0rxxHNs+dSb/xKTVghvIkrpS7RPBwnIAOhf/9zvg3KcKR2geEjo+l0
EgFKgf17YNoY6bLQTBajQbA89clA7GcUQnykB+mMp/pYFg/bOf1xDXt0NWZoGU+L
wDJBIiUpjPqGDTfaB6nJqpixK/QYfVQ8BBMxLivzHzvEXvUed9AFKMfKuyArTdLQ
ywhiGv0tOM+owQIkEG0g1zY0s427S/Jejg80LoYnpKEaE00ZSQvOr+k8KPAwqt2H
8TtxOVG517uNXBOawyW0hF5M6TVAGRE70FOKnBMPanH5pcVvO5Z3OzNsa4b5st0T
ufmzqlf5yekjCB0rcvOmaAiQmWDvPtp9gOe3cDwzxkj4YoxtTGfBHBx/soAJbnBe
NOmrJQ7PWoFS3I/38zcMPTWgS/pCLHoFhSGO7ckeqHMH/2iwHt6iBIUX8ofhh3Zy
S3uk5hrK9D+T1jfEwWzOklE9IVvl9vjB/e99GBSe4ExZ+mXz5VdSVk2g5Ctkw3Hj
1RcOQElZ1+hsIIgb3LG8G3e6iyKQBY+CNYWPTnxKI5fMn6QwFSVKc6mx6QkpYxjf
p9XHoQv4PTW86VkD0tl8R44D1QZxxIU5iudQ599o2MoWh7EDBy+vuNv5lux3xY4Q
nA8OqcSQvZOCUkSobjrbZp9OLhT57JAx2ekWgzX+7IuO20q++V5tDny0qhIOZf72
bCsGddVwaQcJ8ij94dhEFBXwiRrjwvDDzWSv8/37OnJ2R6pEZ6igCN1m3mmLXN/L
s0d26YESzqgibYmv7DroIH/9VjzNH2h7V8QNyJlS/vxtGGq0vdYt6998elmZGUKp
ZcdSi0ZKQF9B3zpYbUBhsspEJPdLA3wgZSmCTEFgc5osxwGukqmrMKnWDtWkseTL
jcmvoSK1YlIuGFUdxqOyX6vBLuZxgONo3qXNqt5oy6uqos+5wBTYYd/ZYZ1mP2a2
J9hCpfiMcXod4EqQ/pdCp/4btqFz4fFdLtmVMJiL7yJ7riG99ltmStBqBR0ruvnK
I1qHkXxQk7Xwd0zXGg3SX2EGYl/A1fMGoTPcnqZKYYF5NYXFyZ3uvIHtwchzhrpN
2pFGs7rAsbMu4Rvup0puDT3OB6pHX5EK3Iu9Pkb49Yv5ygyYeYRkBYi7EQ1Tu6z/
L0Q8XFlcp03JnkvSi0dFwPbnFcKlme7CNzNW2pQzJB+qWuMo6QE+cVAwoW+ZRORA
fF1igxpEyoUe+wSo0fYoJAlX+auxwJP7+lRncVOkCd55YsahxLscSfvrCPXdxLXi
9CITFSCw/p+j5eSLcpD9vv5uhFcvqnqFNtICcX7J8Z3BDqHL73Oyda5+MiNDx4do
ldEVQb9ldiVwSHOpCL4vup+MuYFvKtXa3UcKcYMUCslK9kk7baKCwXKjH83zS6FZ
C7HG4OoOUBAeSf8t1l6ToLvOk4fWkNNpc+y5ng/YoAAK59NFSk5aYPhWTegb5Obk
QecKkooJgFZkD83zQNx7nqbXuM56yVtULcjqoGMFp39Dx2AWd6x+4aPrnpA0uZeK
NrkDuJhdlVkZrz4pHLfVa0m8forrdc8159ys3GHkRIGBd/HKwZxswP/FVhHYuEJ7
UPEkHeuko3mHtH4DHf81ezFg8iLyBW9zeLktDF3bo6voRMQJF2P1oZ13Fif7LvIZ
cKcBsBHCCMAWaeLtsrEWdu0Y1m4Rsei1wTIh8aGATXMT3IeBk1Ju/MHrDAqJw2XL
iNz9UgcaknSW5bkdHpXTjpJuWoBNx/mzK6GsndbidLyuYxGC6FP8vZBvNO9WO2H1
mCabkmwFXjiZSgGETL41YxjSV5Ea8uSeRJIN8Q+5aPy6MqWUupqtXpQqaE0vShjr
NbO1mjRdRFdVqJo9u1GHdUYDIj3RCBHGHcM6kyTt2Vvhv/GrAZbQMLidD8xsl3mM
ESzPkZhAC7V13cCVzwbMisrSeAIS7UZzPgEyq4lwun02KcFTi3OJyU4ukJijzSNh
Sc0WmNPWsYrM0BXQ6QK+7YUd8ZyDmdPiHvczusB6ZcPLg9PtzxoEDhqWD5iDwF4i
dhseas2q3q73Q31SDdZcdeNHv3S0PGarxvT+Zryliv/MZEXEy9Dp4OvQxV0YTq63
mp06GOyR74fZoVacKsOBPNkyfFBTgxuZi/0WYzBUDxQ6xarC95cCV2HbczNIFVrs
TsmcaxswiviIUS0ubqiADr4cER6Sh8hYvpbfqDJyCgKseR9iqtCgzgOh+mdcx0uJ
MapXUHjPTUZFHxabHWfW5T5zMm1tFqUjC2nya2DmzON1IcWICC1bWzt83tjz212T
NWmXXJL+XEmR9xDeELmwFppI+AOMz3D8FIsJPSQZ+Fg4ALUA7EMdiFiKczktNOlX
Z4I6mfzdcJ2hvd1wSC7zgHylSuf98cpoQNHA+xuBdYsJIxc2arRQc6q0ldENbIvd
BzoQG+m8pvuWt0hTIOofHq82EHhC3XN2gmzpaJzVbcfBreD/i3mKaV1YXHsfjucd
4OlyXSYj+k/ETWq3nYhZQIQ0pKp6BCo/6cn6R6rajMb+nSdRXUNBnd2uNDCJLUxi
x7XjlSeytAb/8uJJLoTgtFQ7e3X1suGkldUto1EHT9PORTKXKOFnIaMPD8CdaNBZ
L9sA1dFXKInTgLRIigJDNTMAd0iMaAbQHHWe1Q9emeIjOuk7mY0+hk1URyt1qSzw
rApcsRlZlQS6MoUUnJ6zmzQWe2LNOtYdeaztCB7SDiDOJ4qyhkhdL9GyjqNy3rIb
eBYOCtJX91CordcIi5uM53+CWXGbfo1ubaUUzgTN4GpWY6dYhHiVFE28qZ5G8+mB
hKK9z0yet5G/MO/w4GPObpAjleKhWwpTfuEEG0XTmBjGBvE58pA0Mk8KVePJ38eJ
HL3ZMd84E1AhsnoTa27Uu0De5+g1tIzxlbiivcyH2arHEF94nWP3eLwLm57tr/yk
Gh/hoboQNHG+HNHXZ1Q88xVmSza06WwTXVhEc2rbuf8gX2I7T8vxiFPzDG//prRy
njLTLO/ePjJkHPUiGT6Q7GjbBDf9CYVL6ZpI9NRNbSVCkdkw1CRnGZX3Y9ljbi9r
4nMa0z+FzFkQ+1Gf9LxUH7D9Rxl8oRDqMrEPlMWT5oVBYgfXhPEAx7hoCyiwU4J2
KuIF0tN3A3C3yorKPhhFxhVc27szEzEjs5yfWasUGTkfpCcgAEzSDpQ9N4/BG3gG
9Gmndbjcn5Imm2AqrJya8MuXF8WC2tdZjZGtwNBtS6NVfmvCOeyoMkvjBsWCgr7i
Ag3XrPNoXPg6qmENhiuN2VaXgWF2s4Jabbj43oJNpbaIwB2WFuOb4BhHKqKW6D66
D8xdxUGUORAGmsnQ0ipHpyd1FkrgAcjQ8Mr96Q1t4tW+zH8v8RFmeDXm7YTog+tK
zzOvVpFuvsU4FLiaD4JgmpgzHOUqCbMgsrHdgsS6Ie3oSPX8abXBE96QplZKQQwR
C3ltjN3qJfihZqfif4fUmTnngZ1YRrO0kBiInUlCp1iWZM/rqb0f3ffzZDwih1XJ
GR5q4pm1hHpvH0SFZkXNRBUjUvVi2azxkGznRiXxtsmUCtGf5bmip3zKaY/Xj6gD
MBxU5XUTOJ3Ys77hVif8hpBEE7PtdPW0iGh65ClvczEcBsBSRjt/4Vih5kJZKOVr
epTsC+lR8SK9rWkD5+PC58daq1peAFtcl38rljW8HHODfVZAfRWktDOjPJZCJM0d
zzbh7u6KzvfG9Qh062DyFtlzTVlZuSjQkuEiubTbYpHTD6e6XPaSEiN5lq4atbr7
3JQCUj4Dc79lVe3tess3CaHBkuQEqJ7l6m1hXGzUsw73L31iAb8lKGMIeBjdIKol
aQ8BR7hDjcVY2AF/NbHkcmOmNM7yTf38MbKdPKRzXib1rU2VYokxD9H2NeWKtMUM
RsyBjLenSidcQgkmhQkKGOCzqPEZSpJ1KTv8l9P+BgvLyALN+ntCnwSUK5DJQcw+
Q8DMJ69vxDwV6NGkybd+SjAsfN+3CIxew7/tG50HnCSCxv8K2RgvPGyGDGK+hi3G
I1c4Gii/vXZTs7KHDsWmRbt792bKRTrNfjMwvmCh/aHRAq2R03beKamX3OT3AD1u
4/g5iDMMcz9XqPD5fjZ5O/2I7pnAgp1+rOCP/Wq/Aogs+8MOSzjrjeONnkmzrJWP
LF0I9UYD8xmJRW7XwZjjlE8+FxUyyL1iexsWkFRYF4MfaUjcdqaoTWInI7FokVD8
LTDwKp0aXDrW/kEvUq74ddLRWMfhkx11yALT/Ssq4GZlLp3sb6HcI276hnY7fE34
4jdZ552D1qDcrDRJ2ZSBeCNhUhhPzoMhnVq/o8iw1wE+ff6y0CWLdvZRHVLsmOHy
9UsOnL2TaP+P2ekluZQigWPinRkvIc3rmHQRDuyRE/4bdVpXZkn3my5QR6sSorFx
v+ISo84bzyVASuozFPH8RgpE90Zl7F2A2NM7CzX7LDmfb7Qf6U+a2DFBC7dEM9qj
FUAqdMKgzkXCcBA4uoZlLbwKaBgHGZOMGwmI5G+NJBOFsNpTZmcrAupW9zk1U1RG
I0GDrbqjEXxo2qR3ql3dOF4jhcGiFJZqqgAO53klBCLNeoIf5hsAja5f/Ja+5Nbv
qjAuTOnBf9LoXicS9WK9LRvq2TKLiSC3eW0MxWmAeOpr9Plgxukl+tnJFSezyhgb
0AqAJQsBmGwLgB5XaGbmxR3lzfpz3mSwk4dVDiaq+0w7e40jwCPpGwnTx3UW8lYq
DuFkwITBXbiqe/mYgZHXVsX8jCmCMjKn7JtEXiPtqulSYb+sXL7S5TgU3Pk1Y8A+
Zj0LGo6q5LawjmPRWJUxEY9ZrVyYxMINBXlgo8gQNDVasXWWaFihDSiejV2hErEQ
WwxFTRztFgJ+i5njUyL9Sw9OcwwvooJ2278nBHMS4kATqroYUzZ50OrhGmWxwj6r
8GjSU/3I8HmP+PjMk3PF0s8vO6NY/nWE57/Q6LPTT19DtSrzdJx/PZtvLn+0NfQS
QffsvNKq9CoeXJJvfvCOQyoigAxECVuHAuLCYWr7PI3c1B3vTlbeqIaQwcyq6Ost
lY07xMk7IN/3HSfoCoWAsSWmUhPNLE+x/8FJqPx72QE6GtVSO150ClsATeBoggzV
LizVYccPz0wxBtk1XRKRWyvYgxLFrh4NQbc6TytYWQ4S8xsaOv3cfP5yIoSnEBoP
5YVLc5GPZRO2htd4UMnxQHN0LUR/kE1awpAEfwXo9Fai95KnCG1WrWGUyyk7qVeV
k/WboOSpdtQa1yoYGMBhRlG7txLCmiXYiNz9F7ZtMs1iIORMwBcYqoRmgPh1tMgg
sWIFUAoXd0yOkJwpwh44P12NhsHzVbif5SZGF85jC2Jdkby/ZmEnSi6l1eLcxods
/86wEXFse4hIOFP5mPh7ZKXX6RpoKOIaWfOaQD8YrD5Cv6XK9JbwEB+Dz38OXv1t
ZQNZu9PDSASh8MsIfPDXVy1C/HwuSSr/AaH1mt09WylXvLWl8d7qw9wRYD9HmrFn
JVMdCVBVWLP9mi7v83/EZHxpj8z42Yyww6BqAHGF5hO0/mwaEeEsVDQvYzzfF9eA
ReriePdGnBPMeD/+0b0ozFqGpEfznbcMxyjJpMWuW80seR5kSfxCru17dkQAv7iq
m4Ib0KEag8xWMB+pWyP+EnKRPlLWolUCU4ntU0QKUQe3BSpo6/UTqV+vChUoA4r7
P6aJHaG+Oy0hiMBZK3huEP0WMArvXX2ae7bcAl0CaNQUnktpBeFOjH8qQ3x9AlJ6
Flvc+Ie8sxisab6LXiFN6bl6A3q9P8Yrfwozk1CPgphq13ljH8fWfrSPYrPctl5Z
YCMWWnAJwWxbOwUTmrr/maa+4EwBSQq5iY7fqcMv76dghc4JMV+Hv582R9kIT2jw
uaFf0jHw+PnY0eQZbZIEt60fVJDqZNkv94LMkenm0jTNrq+oUVZoGPP6zw0VRXIt
BOUqFPn2wa5sCamQH5m0NYuIHoZ1SfC9t5Cu5wJMEo818AkObJHEDkKl94K58Iir
KeL2afTvftUSxkvwgNgeEWYte5typs5RfzhFQArpni6JSHcImmD6hPKVPe49Heyx
nWMUp16hKL27qPZeEBgypKZmuRhNlRHtHhdk0FNgX3DP9/74bipI11Sj4vTwBwYj
pxBZD9Sqtk2o0RyiFVdglQ0WXpEwFqOM/b3mMXOZJm1xOKF3PhKTJSaM5qBh8IvN
XtB8OH8eRjCP2yt40IXPNHEYpbXVNrdytWVR67QB7hCzi4vGxansoAV+ve+2rGiv
LBPm0ATEINx4r7H7t2a7L2CQL+2oTeV7FaJzWQDThm3tbn53x/BgV2XI2Ag01MpN
xtkS7t5QORM3VrYV4iKQ/cLQIVH3aTphQ7QcLMoZfstqUXLJ14NrQ4wBlk/2qsM1
IbL6agRAO0vv23q8vDPxapdPKprMo1hzXLLvYSiqty7EMJyydazIPnhI2U272TTB
JhfNRThmxhoVCHt8RoA6q8prYyZvD4OTZKkQBjE5DqMljnCd/y7VZPthaQKrZNUa
XG8aWdU37yLQg7fvQufchcD0LUu4zOogNLneB0U1e3XC40HN3OTnBurBF7LccQB6
5NsG8ojhXGKGRcR6NF3XEEeAka+67hzNmliJugbHumjClhXgabHjmfub1IMk3H70
TlVHEo33zs7CSzy9OCPoc0dv+Il3tRCaS3kA+F8RbtRKFwp7pQXNsOqZ3I++V9v3
xHtQXYYU8xxfTjZos3wV2ssKelZjNh9qDEBlduZKF6ryAWDXBRna100tbEe3Tr34
9InermRr7ppXa0trSt5K3FCt38vku+3Sux3ci47aw3pKI/9mHhEPDMTtvDtu7IUR
pE/ADey5toU/CChvMEaIJxk5sDdEmeI47zLaCX8ulvNnJQVcaF4TEI5eTH8SvRT0
9hz7V5Gr4PUrE1ADPRudacTjKUpCYvDVbHmR4dSFyWB/wyI9o0DUdWELL6fg0qdz
V3r3BnV8FswfUPn1Doykfa+vNgGmi1rToFPBFgGZS29IiyJvS5QQC/hwU9YnDqf6
dlNDaO7tkP57k67gIr+EQB5D4K22hRkWtaQpY3CBvWQz6UpiMGnHJRCK5+YTk1Ii
+40HgftA87RYlq7+oXrLswCHpXsmWWhHyDzkNvC3ZlNZdmJJuzFDmMgNlMm5lRDm
nNUeQ1y0YZiE74SivK7NOgwhZHUyYb/bqCk/vP5mYuOmwx4x+qxPdQkv8YynsI84
bvGLToK6woUKNA+9uKbxrjdh/cTDv2SeG4j5Iz1nHhMyjluq1lt6QTwcL9YSs+L9
fZGRS+UFKS9rqKxVb7fACVIqP3tb7ATStZOyFwldihml1OEmeMMOwgtcoFmjPGTp
h8c7VUNdsZ95VP2tJ+bRcD+djgnGSPnSOqOy/cWujrHl7GJrRpFoznC1vVNsA0xB
WPbLJpZvfljSWScTzF9RWK6KV9wbZsYINrCfztBR/0EdgWMtoTnehEbGJAw1cuKT
4PmiWDQPZ+UzhlitBvdN4yS0xqIty+Z79PlMUL+ktZPc5eoFXl++BKK6tBMLCQlb
d39l/i4Xs52zl++Q/iu7K8x5wfGx++UlyOFUEZgnZKHp1SQznLf/6+fO44cBqtPl
c4hOMxXJBvuMi5iVlG3XtRa5Yff6sorNuQBEILgy3JIg09QQWi18Twl6CJcy2IyY
7pghSIWNMSmFBGlowSpXjMB+2VNdIKaKW8EgCloxG7qGJf+S61tbYCk0H8H4bZGr
r+zMpCwtas9ywbaJVgaVfqf/VDUStovsUl+y/iXObwt7v6hy7d+2W+fWZicJZcTN
LI3NS+QmM1H+2atX9Xbqfl8ayExw+q8llij697XXeUpIqay28tEFbUodJqx8WAf6
Ng71aWvhrFM+9r4W4mJh13yHW0kD9ncHVCXiix49VsJtHNZh3NK1knrWEJwfcaTm
iX6G5ZD8ls94o+PXJnGMNPCOK36v9KE2ToJbMg3z5MUxChgJIIWlFZXMx+tFoMaR
GUlkJjJ1iO/iuqwGMS5h3cWtvKUdOOYf7JWo5I7eM/a4nAiwO2X9oDROR/ENvdFT
5y9HYwaR21bmr0C78isoU8TW1dVGq1WVl1MXQmimOmXxFz31ND6UlUQPscXkTVxn
q1zPqnjoeMUv6s6UHSmZI4WXnRwIGyuMvzYUzpoinsOb5NXO6Qg3zegONR4kpbxG
sWTM++5JSPfkVqCJ66u6CU2NWJlYrHZWnB96qErpzlbSFfLM8rp70Lun+hh/iEtK
1lD/WbH4jf+ufthIXQRYMSw6KhEHAvqtnCNfdaW0HsOKhtgiINcNI2mAItcTumUx
7/m2ys3c9BKcrHqkVgP1Hy8qfh7t49rX1oWb8VGD8v7cpqrERqeZFGK8G7raWem6
bHM18kT287o+KWbQfRzAuaouR33mjnnf0W0eSHCmV6Xkl5W6PduQ91r7MgO5RXsa
WkZDq3Jir6rBXn+mqsYMscNsSyTPweS/+426sA3JhsCp2lJQEJG4bmoBWuH36PBz
BzV7xNGwE31wM86HOqCH8V7+0Zehdlxeqyr4zOKf9cUkWmob6RjQZJG6ZjJZZhxD
yNQHkMLdNdQhKY4d+PmGZgW/afZkv75mowGInO19LUT1KgsBDbsKGojumnqcOWtt
cmd3AMNXCfTLEIzb1FzINQeUlkwme9YQxoh/QZkBoI8e/QefqFm/3w9jfD6268YF
OiNzW9VQr2Q06BdGO+H945GOS+FNXTvZUvZIB5ler6JYm1dpbSIB0gtmg3psNJmt
C6LvJ/JqRsL9u8S/n5XGHlA/Oc3ZaCdD7OXncUXMpwIccUduTGFaMba9N6t/k2Eg
/aKUI5Xshl531UVmPEhs7sPHt0YM+aborjlHRiVEtWl/h+X3n6ctuanKTHZnXIKy
N0SpPap8VUaEDt+M/tTLqIbq6BindtiGB6JJv8UN0YqAwVLhrjW2e7qnnq70fVK6
pFiIzoF6lceIsFH6bkED7asE7Bip7BjNClmBs/GennsiRNUf06xXD+2BeiDLdaBq
SBIewNMhKMYWXfJVUzhNC9h+5QEVqlTQ1K49CfEsenGYxmRzY2DQrli9w7BTZtMi
7wtFO5cPFgLP/JdDbh04IN1+AtTtYfX90gU1xHWFRAC9bRU1Apx7fRCdKQ+iuhfY
2HhVgEELdNhsFK6slTAJRo055pFXtbsNRHNEEC7K5a1FvGVGsL3j/IwAejxmF+R2
00xygadBTpKP6XQgF/OTKGzfVX6VIBH28GF/MZYOEVG+XBhtIANfp6CDVYNfwbPk
MHGieOfgLdnelJ6bJcUOq7XiQOwOCHVBsFSGII5/a4itv13RFW5FydqpfgfhxgRc
CTHiYtg4OsH495dVX9eGEXXfm7E/UV1Mm054zfT/bxFBYUxEBT/9DGkErIi1WrTW
kSWQcSLdWowvnUAodysNdf7k/UD4Y3BaoP3FvdeZgnTJN31/hzIwu/4zUHpFeiHV
Hwf00PCPb6wwlHZUYgcAv8hWSfXd6PNG9/DNzULg3ihjN7vpt+Ps06yG0sgTbN+8
1EuzxxZYwACO/KoIp/nwlZegDZoriNn+Umi/MF6yqXcvCM4k8uQ4TD/DReVjd7FV
uf+7bGZtpaLnI3u4dLrN2XetdZfpOHHCUtcFLlW+ey+/MizTmGKQGAZcFfEFlMoU
tz5NZW1Q2mIy2FmX39wjDGTp0iaHeUWUgQ94D8qsBipX75zEBtwcgMeuDN8j2NY3
o+INhs93OiFRrzR9s+9EYZU2e0lmIGsVUD5kZqdWtELcoSdpSA9Pc/gIp2gRbE8o
6+MLMRHLi5PMr+FerMzYAmxr4C9VaafI5cl0foTCd5PLJEJj072AMrZRzVCYsIiM
wk7U7dI+e+GxUtZH9APKqQHugdofDwq2nlqy8xsL3icA6JHQkoIcv81DIxvHl+nW
O+cY58gJpQWFNJs+q2xtcS96tcfq/jIBQfDImjPwWriTGipsgZput1kVi8KoM4go
jzMwnpZC5RKd0Hz7OJY8XD3IjOM/Yvpcty+a8B76MoJEuQ5Ny6aKRRJTJiEWhg+a
mjZx+MjEnILYI0TpFiMm7/ngNXHDLn65N5x1j4RBH9kK5AI6sBLtPa9sjTCkXPOK
lhosPbW4DH7CFzNGCS8+1UVdj5ZQPs/nOUJZ2iapJbUbVU6bULCztUwj/09y1HCX
3GSzfpVUx32F0E/GCKAfLy6jEuaaRFmSCH2c8TSkkLQf50Tfpzk/h+0nnYpG2Y1r
fzT3G04Z76netRxLkADuHdjEyw0xCrz5kskYXBzF0wIjpSHNmxCBH12XgYrq+8da
NqAZPW5bM8RFG321tXU0tBSDsJ6pQngBMKFcUZz/EYf11/jRVOpmF8NWrrRheBuM
IFvPvAKd5FkU1frRjyNBJHS6U3iAaM2cRg7SBZc9HpLMNlkVcPxNwQscWWO72HU/
oo6Pj5mMm2bTzOdf3qE1/qjD0PB8GLgDnCbMZ+0GajHNcZexPzFcXrkGCQ2KLPBp
pQwA6IeyqF+GnYVbuPpkHaUCy6DAF0PxyR2RCsPmp6ePr2jmrSFBm9QMstjgRfHZ
9d70SNP29rJY+cpBEuSsForhzuA/bRP0JG6wyBxIwcniGIGQ+J5tI4So3cMc9IeP
XUN+FzFX7orWtJtxRlTXsaZHrilIQ6Ag9fIz12ZUeOLrZcBksXXvx8MeWvPz/Ad5
p13A2vvCqVToSEg6xkaiKKrchemmNM61bxW9fr2Xdjd4zVNV2LlUCZILwXIfvLp3
2fqBa5Xtb1jvE6xouUTUd6WVtrBLYk6trc146BQCerXAJx0fv9mGguTJjLIKG5ND
fGW6dgvSXSEkG7qzHoi7vrv8CZ1XTO0W/0TC7s6eqKg2SfIepwWT5YinUa+JM8W2
O1OIaxM3gzMxKL1PLJjp/93xzsjx8/or4T36LdWN6cr5qemDwCCaHSdYTTptXCl7
w2aeHGGoOXEm+awpkZoy1nd1JFqfCjbm/T1/XfvIyST5W1Ppvbk/3thtAzIIvHxe
lZm0R+3dx9VIXAk+Qrun0iAYvjglwDHI52i46rLUmvNgsSwGgRy6kz5jNsnYCDWf
gDDuv/4C7hwHuDorSUX37w0WJJ9M+SHLlsS8N38xgAdRQPSckqBquZc71tdDfh5x
gK2G5FUhXwHNyl8/IJ/YcCDfGmODGby5kpehtehw3aG/nOC+GUzy7ZDFjz6KF+CA
gNrSYEzNZupwfAJYCWS36jeXaFqgbjVaGh/TUv0seIVNpVIggkPyPAsijDwGXWLX
liv66XcEXVP24j13/51tOkDGI3xpWPGMzqXozXZ0r3gz8DwlyE+1D/9WE0c8D2Ow
QjNdwD+uosEMpLY5WW0cVJhvDWcHWhS8qnS98PgOIUa3BJJAP8ieuiC33rbZ9aCE
VFArSt87oh4XXegWDiPD/U3wz7+seNvxjyxbZfQS2goyqagYqfJ34E1RU7cZpD1u
rZoNBAlHw2cOPOf80rmrN4Cb1gpuDGiMFqV8j9bxPP9QlggXUY8S9jnHDc6YVJ02
q+iOJaxWBiECfpQfHoo19hiZQt+o7eZo2RN/q67D/t0iRwln1QpLQHCY6VxRvkJq
Ug1eV918lOwcL3AmoN9aOC9+Q3HsZfPTEbUdqI9+60yqCyhxnr3r/0NUr/d7ke5r
T1Aq0PXjty502byhIZFv8M6OMZUVZR3vXSkNwY2H8JwQuSp3HC/wQf4at9Fwo1oB
8BB48XmJYbZAqKuWPpd23N2ZWWWPls03VPiQ2T5xurANDa/GB7wlR5EySlWzMITN
C88J9uXFsQQZUsHXWAY2SGnSbwVQqaS1o/ifp0Y7DTSitIoMJ4+4vMQghluULoIx
uSxj3VJeH6KYeIX/9Oc6GCBNv+r5RqAPLNy0KZED0ZQ5HCAAJ/8qANidqtuSNY3D
rGl9yE5usMKv4FZe+Tq2L7KMiFPR1/hFUQfBMA5wJ03DfsXiKqMetZF4HbTAlMmL
UokfiaxhMhEorZlIRKUNyPeNPXajo2cE6kmfNRqMYBE3w+SU5n5CUsqLx6ZbGkdI
fyVQlCHsdrqaUeCp/SEo0UEJedtAuOWw8g23ZDwjNlzBF2l0vBBnNIWSKJ1w7v+i
vK37IR3G/B6NoM+OiPhubIYBmSWyhxY1ksxU9iLB7IM/uxIYhYDULrgPhKoMxENc
/0SfUxRt3C7OsNH80qDnZ1YfQT7Vp3nHQkwwbl/A+CPzV0JHOADf2ssXoRliuzvz
uwQdcERbPE0ALOVbTkD9Kcep6L7t/laTvSHqCc8hXNOTXzSBKa6t07W6UiEmBEL/
vEr4WPys8WOQmesjdUMU+MOAhhOyID8kBtdabkDWnfMvWYatjFC+KgFHZHEERzZc
/EQvyejLnpzsXeBo/rimJBJB1bf7jSAX5kt7jKiwhFeIXTSFXHphdkNUaBqW8nCT
lfWi1Y/et0m6rtqSueNm2/AU4M+BptQZ/vCikv+SPkbMcXkjZZdlSxhmY1Nr1J5x
MZs7ULmhvvPxgCAm28dBlpzHPJI49trHbQlLoGn7NBG9P6bbkM9RonxY89ftqHaU
rqgXj2NtRiYuAhgy3sqatsypASeHEsUz4mRyraG+TCOEG2CKVUY4Q/38M6mMybpd
vIq/+h50PlJq22AP6SdldyTjKL1bOCRJujR45LZa7+jVnvvy9uKEkiWTrn6WvTxX
xzmpVIT3ryRkidSIjhnUuzVwe6V+q0gnJMbwc7bHMJO9PgExacXEwFpaGabMEfCL
OQtz+u/WSGAILckXHYSE9ZvAXsJGRzHbfQuZsgtieeddwmPGBVtMaXvKkBFa/vNL
ETkyvW7wzWpJpRCK1lWsgI7uU7JkjoPQ1y3zVSkPBN3HA0N/J6VVSziOphLyawZD
PzCtjqiRSXLVda3hGIEhq+Wtos0huci+sEDJXSAnplPvmQsp8gC/mrBUQ5cZGRq3
lI6HOY0ygOcyutZIl25vQXQkmpGt9ogCLbvYKMgeESxvArwJrcAmuoluTy08+3we
1KRg7Rq3bjflYZZhLyR6BcZ2jmsqtbnliYzSktzZ/KBcJTX89oRI0SjP1LzJBW4j
cMZPtIXaUB93V4dKT7pW5HuAW2pKa59hOznGfP8RJsyMRYEqD+PcYnLBwoyRFG2G
KBny052CRcOBnQ79EOCiWpaZ/l5zo11KdNcbg6VQSabQJqHzNHiuM8pYqURabq64
BibyDcKvtS4b3KmBryRKq3my0TB/4M4LPZ+jNCMU/Y85w6XLq5ZBk9hw+AV6QVCS
H2WfzJN1GiGgjAwjUdrMhRYntxuQO3S/nxb+vNYS3+a4YdOIJ4dp4WuU1+a3+7xG
pq8/1RbEV6JXxpz+4fmAGxiGLfqT4P2hUmWt9GMg5+zBDmQlGc2wXK7BCGrTXhzs
pE2MNQfv812HBH9WTn0AQ2++6QkFcIMgzkx/4lIH0nzkuBkILiXZaUuxeIkUse0l
7/j7L/TKB/etsjLGgv4nrTao9suH+fTrFHFDkSaZdycIVuSYRxX9lmJtTgqwOnyP
+ZWktuZsX5zMaKYWL1fDL6ovAVUeoWUX5q8kX6yjEM98WYxiw9bm7NjgXN+zTyAv
ba8f2pgb68rdAvwjn2ov1VL4rFVMSm8nYYXKTa1o3jbVjNcEl9wnZEPalKhe+AaI
tLZaA5WNWahU2rCXNJ6NgoCaf4+f5NfAR3Of9As/IqVppozWTSEnrEVKX70o4hKq
ObVOqemabsMX4aZ7nOp4+Dw2Ck2sr5iXMS9Uu8avFms+8NNFtCWlJBqC3PtdmbTx
AxzLIB8ZHqz7TIXPBouRdvJOkoIGItKAHjnDrrwi6v8OAIWwmTMecC21LppA9onJ
Lvvld5ll0Vu+KY4BPItrgVZONE8nCP5i+htz6YGI9tDq//t2B3CbjjY0fzSocVDI
4O53e2Sp65BzB4RcbYystm1SE34oaChlBJXIc9I0bhNl8SoBf56vhXja8LZqBbdz
bfI9YRGOUBvl2bDmC3Kn1uUumi9D0X/uJTIjI2hEmcgPsNA79Zhzxo/eHXscPX6y
4C/IbPqog2cnn2ZRsLComiUiNbEIcCRxUJhoghW92l85zrT+Ej27zbiiUmXTtHfH
3uW2w9Gw3WH1zZLYqgG9bSKa+v4q0YzAOfLaQoSLiXDwL3/bZQ5EMXU3RVM6PNsc
zV8soq9ThDii68mDDHP7MdO3Sqggwb5R80sg5OBcjfUh3owV74/Z95W4mj1zX6db
yQUrQRf5sxRfyLKG+7Ko02Snc7eEmT377lRqilOJNnnxwTgRjOQ0n1ih9kYMyZz4
9ekaSEJz/pvgARvszJlDxAe5d9g2E0wu4ysdA5bzyguhjbSPjUWhFZjj3CpRIOj9
3ZRi3ZfRvRavxRFwLIdBk9+QIJhSNYDpJqbhYYZnYyCfAnzhiHI5woHI7tQ+hM2F
zU4xYO1PeRmYRv6w+JGGEBtlWnQ06iGhJL4dvMTTc5iwJAlhllhvPG23THRok/ve
VZQBeMqrSLvRiayf4N5pxISv4mUzIoZ5AxR4rHEQonabj0dxMWG9zHvqvlwgSUcV
3XFeX7KuhpM8KWpBnGFeZRR56gaP9deC7q5BnOxOwwxN9Hm9D0Mip5Oe8Klo3ipL
qeHxZyWbNnW3AMPGsXFufyc69F7yyvmNCA1xuHF7v/+4OCxyA5l0BaX5EVnE9t4+
v9BTZlJxsVfWcPZWMv+g73AIgjdXI+4BRi3j9VuO7nIQyQ7xfSHGgLkTv8QbcIqv
LMNeBRqpA9cwmtpBk9ePgwBjMnAU0u1RIPpPnbH7HNeHn8B73BjinCmTVBwoixOJ
5qPeZsHzSZfL0t9pnSNJY1tBB0ekiVnZqCGmwpJYD4KsjvRZZciywmr+H/MREZNp
Qfkx2basbq8NdWSY/qlzxptK6aTCV90Zb7xG/NDgdvbEOV3YJGJbO+Xsps+0wKHl
qGvP97ojYk+1TAA/sOy7b256QnXQf0AEXzUbr4CeMO7M2BCLs1SP4ThB/0WKvzRJ
be/xAEmDe3zfHEfNJKFh7OJDXBx5CqT67jE29B7+UTb7sAEN8VxCiu01349ONYkT
qNGL7H9Xls4td3aYBM/48B7l21AaMF1jZM592bMHLsUo+fNgDDmbWYlCcQV/43I5
N1ZA36WOyTMdwLaa2eK9htDzS92WIO/G2s9/m5NhWdlODJecrQI16rqJcs8Lx8W+
DeKhVCyWKrd3JCqb2QqQoJgwLngvGMHEqX1LLBaMpTWFs+Ru3nt1yQ68mk0eV9Zi
JbD2TPrBhYUVApfCaSbBpduqmWT0c9p6bx7VwswWMwRWE1i3HX1S1aiT/c6ZIybu
GNCgPIsnCmmsceo94fOl7hcqHk7p9yMGOsZiWemeZG3b9NDN7f7tVoaxObhWq1S6
BpyVHqzzY18FnrIzx6Ia0w18JKmjeiF0KjPVVYA9+j06+/EB+fvpSM+0+OU8JEQr
89ly5p4XqV9+M/BIqjiRH7Ix+131m1s0iE6gESAKwYuv+SW3yI7IPdpMrV+DTVLu
2maZ82jsjKe+mNExRLvQ47Sp+g7kewGQqZHBxOW0awj7BT4UF+JgVNfJwm3BQFXR
nfuK8ZbCaCictXZUbqyimrzpsaBVuPk3hUxRc6GvhJQl5Xaz/ClnoBCrVbju4+k6
RwYeSCYt0rWGDJ+nYXVwfywfqrdbcpWGO/bIA/xrk3TvIHBrDN5uHJ3md70lQDue
OH37FmfMuY31veMgssBpXlhdJ4c43KdiWM51oxg9p3SLxv2uQLB56ZDzpUF89Caf
ttvxGOCGur7rgH/XZ0aZTLetPr7KR6FM5jkiA0K7cYHXbkh0Ey+tTjLxsAMetlCg
/p+oxssI5tsER3arHSjQUS5BVT7xNCjigkhW+xDHDmBxfDH/UiBKRIOXUtGrTdTF
z1/R4KHY7qL7Sm/IoNngykxi2vrCnSHaxyD4/L+Pn+VdmKmV6gwS3Jd0PuaEnK4C
6oke7v+QqiecTpJWnqeyUtC5O1OCJcYaLkJwB7Iwrp/o9QvEKUeUHpd5D9SoIyyf
sUQk8LzmDkGq/lL8jGWRqsKgPh5JVbHQvoH4pLW9RX/NuPo+fxj3mWWP9jLI+UaX
uQ1B7sSxueu/M73o1s9iyHujS7NlK1JgTb2IuxJpNBrLuynXf8mSBqu5N072+/Pk
YIvGRDUZ6/uazLBhj31YG5WC5caJ4XnCJrdn0Cn8xy2G43/v+rMGihlB6VwCrgH9
l2Ldx4I1UXc2y5sdYLtqHywsZj09daBTAq+j1hjzd6XMvHBmdWIYH5dY18wKzDHZ
rwNBBHrCEB3dxcy7IH9smtgqNHa+aHqzZgnKBOFDalTBBn79RQz87PHRCycejs6R
x31e+wO1MEFQc8Y1jCoE1dv/ZO3FS2b0udfW6+4JiZVUDlzl03KoBLDl091s3uKz
qLpMK9sdO4urHbjkJkrx/4NqoZIt8J9//WnnYT/X7fNV4SYHv0TQpgMjX3LUDDiw
Nlqgrxu/v7vYddukTvI/jRKhK4SDUl4Rea9v0ejPEUv11gljEGCU/uP8cHPn2rKc
sczjs7RB5UvTSLcioyKFq39vI9Lcz7ZFkQyoMJBML62ZmApeVEzJlTatAylPgQLj
WujN8DlZwofmr9v8YuhVlrMXHHs7AyNKix4eCKN/6V4lSO8aiS2Z3JXCyu5hK1pm
sNsiv6CbGxBiM8V/IPpYU21l/8WOGn+wte+S05KbQgsI2OBNLgdG7RrUYdZV5Aaf
dOL4f28RMtUzfDzzmjy78/oueXx8Rg9DygXyaeo0bsoQPO9h7MdjK/PbIEzeXnGZ
CH1xmmuARU6+kr/SBLL4YMVOTzRrd7dj72w6NuEsxAQ0hKsOw0JhtAMUKEiWmk6t
6lu9brveqhUf6kUfDyCfGyVrU5uCciDsblXPEZYnzxDqAeD1hvhgXHVJWJxjULib
8BFbmj9KsBiy7hSNPZnmcbFMJ5rRwQgGFzFnvFjHw6q+SO1DQkD9LoHrmwq48vU+
KzirRbbN4Vg+5OfUk7TtSR2oyGvJw1BBscS7Ch8FyF1zlZwwOFNnQK4fSrtETDI5
CGoPii4k8wFjeyqDzk3xEWWelgMvzqV6niMS4PAvOQxmm+1VvVoR0djXPFtq+FZ7
PfCw0YmwKro5nd947tSpsVTa0+WVB3O9ZmNsrzI73n0QQbsYItZ64NtXl/BpLyHl
QxI3TnZSB1gicr4HXE+P19ZFtBsMESYOEYzdCBvvTzOkhnElZdnoH2Y2hdcvqVx4
xodLi3WdTI3VAAK0rwyW9hDeehH+08FRUILWIajxEnAobILZFIBxaB898IiE6ciS
SCe+6OLWoRrwWBHVVQU85UzRs+h8rjVDMbEoIdvSQ4GuCM1gKnYLwmu+9y/xc1pN
rC4KHuq83GXlDXeA6A6GRDOilfYFMBdVHMGLHpz2dIaOh9AKFIbW1Tczg8pjOC/Q
NZqdJYB6gFv3MADucBaWRkcpBpQ/8FEwZeSgtIEr3TZQoog+tbMp6NitCU4AmdkK
s9axW85Nqb21qFV7VX4vWpmIxhFoQ9n7ogqybflQTVALYC1ScnYhlKEsQPFARJnh
Ddap1a0EETigDlvL+ENvcM9JjlBWEHkkD9nx+vOwur/lxJ4ZngaOCTO6fdGz9MvO
SmT+NiWyO8+1goCfVik09Ga0dqjiZcyv/t0DxHqs/RDdZRFPicgnOuBkCj9kCT4i
/M5FhvWJCZSr1e6OEv1s8gqVlp6GXWfFBwS0BzXZph4EXeHAw5B4yTV1O5SBu8Tt
04BtxHpZJu8uhw55XRYUbh3YUuKCB0sNSIrEy9ogCQ77NVyPrd5aPxUKk8QPdKNK
yB1BzlR3GdqbGhnPRwmEA6yxXsUO5Tl6wJ5S7BMFI5MARKjXgTSJ0o5RPRmcMA2+
THU9ibE1BOnHZXT8v4DlDrrBNjNp/3X7WYQmItFIEKe6dSM6+1QdkAidBBtzRQvv
ULhRDv/rhp1hLwwbrfTlZZffeHKBklGwWsDyKgK6m6+bD2Czqp0ahFiGI2aRAFKA
h0vGcGJAaSqlzpfqkEEQpFTrhwtv3HoxUFu3vw/VTHishVKX4S8a0WK0M4zs2Pyl
UGIDdbwb8GLpUpz7DG5cJmpUlCIQ6H07xX3PN0YvIyt0iXPzhOz42Q36BXnsqk39
Uue8ddZAMAZmBtyOfsRtj24zSMg86172QuDKCwXrkCnBi2n3ecFMaRlXCvz7NUX6
8r78Dm+1HMbARoJZQy/iVTDoa7GE6m7F9xGw3aJ6bIFeeigMxkqwF0mul5yzjQTc
1RleRph3yq/NJW1ws8DMjBUU5Bbv6hlJVvFSEIp1LkcK4oqPEZIFnuNvIzhapeaT
vbpT8k5kpmXiZP8Sql0P93xKfmAcvOq7Jt7YSa0/LgxSUvBwyO0ph/nVIF3DTWMx
TrZBlyZWtMR4CDIDxEK8qcmo3psL+Pq7O6bOSZd/ThvJLthEgE2fDT951MYhruKz
T3Go77O3PWrhpyGeZj80f5IdAbenZ8Yo9L0zsIvKhv4G97bqYrmi5lDuQMU44WX0
WnoGCc/seEixQGyQUpIkJZYKbUCHimjjpcm6c1JKywtQkeYckwWAY2qNEs5Gtn85
nu3pLxrJ1q5BlCl3ZiqSSpkau4EMYyl+Ruw55WYx979h9lM0p3xZqxjvguwhHbAp
dJqHWwPO+GXYViborBjHl0cinLOkyBJekQLZ/wLBt4oHC0RFuYNGMJ+qpWrsKTdc
ZJIugR3IQ1x+CuC9UztSoaNJvR8+aB3P7KdhFB5Q2RMB5g9+R0XdD4nBt6WcOPLc
o92FpjcsdXue3QNKMITDYLNNzkswUCqigkb1KLC2L5d0wwK/HxqmlQiwJ7rwM70r
DCCBzTfDrZrYE4ll0rP10zxyupUwrxkCA9hYHB9vjUiOuP7THl4R4VK/+2V4bs5g
QiRrB+KaLMi6N3SXRD7MBsSMejiJA6yb1JBiOrBdrVbjBB3AXeBvBxu4zmhwTlmx
/1gIw7PibpG6txWHv8By50iJ3SUcFX4qHeL2uscFTEfaKRecxsGH0fQ22og81oD4
KdNUFOvMlugJ5DY9xyLyWxBuyIsKIcA6Aro12ZtF0/LfF23m90SvTcwxCNcICKtl
1Kh10WmPGjxlduES2+ZqtxRjutzwS3VP4LeZ49XiTF4bM5C/pdFrnJBKpqNB5yWv
xh80DQAkQUET4PyvD1wjL+2q/6Bf+VMpBbLjHHTFgorElo/gBAiDNU0BFSzWXxNT
I66xox4XwGA9SqXM4SoAec5KCQGhTkb3oaAXdGSMWIHfxKfGWjveUat3Ffqz3Zlh
aWmMs1R0k8JFOegeZd+s43Xwn5+JB6BBZ0WD52hN0tWZoaEI3H/fREOwfyQ1s9OF
lP/141Bq+eWCcPlTbdlXPS6FWxfFludyA1qYKhPpHnEp3OEQLwVgHj54j+KZx1x8
mECh6yew6Z1ECqPNJsGxAoq8VSYrr1Mt1wM453t+OHp5MXQ/YsTku01anJvHfAhJ
ne6kcAJpig8z7+3zQlPjDXf4JL75WRriPRFOO6Gb08ZJAGPrF8JlKr4pFPFBNFD5
yd0hykgFe5WWUM9tcVglv33dG1helo0uS5cBtHWSa88ghZobPEymuuiPJm6wFYbz
G3ql0rODqPu7yOndGkLqT461X8BpjviXUxC2rtCXNK57sP17RJfMN3XH8JfQvoaR
faqbd65MjVHmwY3VOFbMqNcoSbqyvl0OTLQlq5Dyv/xk0bHoIVFry7NG19qFqvzX

//pragma protect end_data_block
//pragma protect digest_block
MpFot9LMub1q1CkxGidIUHWamnI=
//pragma protect end_digest_block
//pragma protect end_protected

`endif

`endif   // GUARD CCI400_CHECKS_ENABLED
