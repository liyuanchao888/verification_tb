
`ifndef GUARD_SVT_AXI_INTERCONNECT_COMMON_SV
`define GUARD_SVT_AXI_INTERCONNECT_COMMON_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif
`include "svt_axi_defines.svi"

//vcs_lic_vip_protect 
  `protected
<1g6<5<^;fN/OM087c6?W/=0ZCW6]bZ?I,07HRJ]YO0J,S\&IE\#6(JTa.DbKEL6
Pa[0-ZHF^&d773ILcR@LU1^a?WKa9<P<FRCV0_H=@eg4]Zff0#L9?QXb7cPA:3BL
?OD4&]?S,^NH]c7CcB4f]Ye@.K.DO?=WJ6SWOU-.;WY-(AD5K^L00OQc-Z#A^:X@
2c?^2M=Q21)R6+[.>8V/4g.=FR=52T8>cX=>;f^1&JN=..SaJ&J@&YP;(JFI8SHc
#):dH79KN>\@6X,+.W3#JYN&H4A0G0?/=)<_J.I-6ZSX?gCA#1,WVE_T>6KP2P85
_[T2LF/3bFO7L:NI[,:9(6>E]D:U6M-[;B<^)WH)(-46P-F>2+S;;=TNA]c7P?+F
G0>6F2,7L-Z-E[fXg5IIE2=3&:\J./&>:9^_S@?FNA&8bGNg99S0UZ(V>2H2/]M5
)BUVSLb.X7=PB<84K(?F1<J;<f.<L2GUf28AQG?BXZ#5Yc.UdZ.)]\d0L.BdP/\E
M(_O/Z-K#[RSL4:\aHGI2gK;B04<9X#FUH(VL(D+N?=;IbW&gXG6/.I2;XWJ&Q3-
A.DB<-6[M&c.c[@=MIaQ?EDgg1Ne@b>Q6?YDgVK+N=#7#P[7bS]:bS4HFb6^b,5c
L92cYP,6E<LL1TM^d\&-W,@:d7IM0A8#0)X\UTM@T@DUYO&BCMO5,f/>?1>DWCf0
#6g(G+M\>&S+6W:RXAWcI^>VRQENWA-Y[CT=9;RU=N.dQM=eN^N)HBN8UM]gPJQ0
:D)O-<#/LY]VJ0E0egJ4MMDJ[;\\[FHV;<^][SJ+EZ?>O@7f7V^+F0[HEfDfR7f6
\W/07f5EO_2Y57;?LV@D2=F]fYEU#LRL]:FGE-Ld2:Q.6N:R(H<UW=M08TW1MW/Y
bC-+/Q/e+YdeV.K90T&a\#D@>1UV13SD8YcR(a+b9.;Q[OC6B&f<CH3?M&OC@71Y
aMEN3\_F-EZ\=_:4OQ?V58DR0Ha=/-I>W2,CQDOC>0/dQMc=I_DdI2GH)0RB]H&:
ZI8[PD_K,;B)#?a0>:OQQ>0CX;ZUffE4YAQ#:,#G/JI#B)C@(&Z6P[Gg##b(eB,B
&G]O6/NDOb:6RS\c6R#C15,?C=ZCNeN+\d-=QVAe@PF]OP]E>/-P+a=R5MB-HH;#
e.^-Y&MeSI?.1aK>U4&/TJLDQ6?P03/QT(>_2E_<@S@^D04B,=fb(E5ZaZBdU)<,
14bDBI\#dAT;:1Ed:38+A4>U[(2)+0T5B2.)#UZ2&<FU^(<#U^K7ea7HLPbc7CCS
MQ:3/@2A[_5e[+F7][@+EM&ZY>@]@YRQ3R^#^<O[0gX?fF,C)DHY(,\R6fJOCFK;
S4^1dK?.227KII4T7WC\J[VY+eeXTR41]0<XZB7ZX6@[F3+\B8FY#O#\+28-KQ6Z
U5][:FV_)\RLV>3U-.UPKU=Nd+F)=e.fP7&)fb?3T./LQTCEU6+-/3;TP>L:1(KPR$
`endprotected


typedef class svt_axi_interconnect;
`ifdef SVT_UVM_TECHNOLOGY
typedef class svt_axi_interconnect_env;
`elsif SVT_OVM_TECHNOLOGY
typedef class svt_axi_interconnect_env;
`else
typedef class svt_axi_interconnect_group;
`endif

/** @cond PRIVATE */
class svt_axi_interconnect_common;

`ifndef __SVDOC__
  typedef virtual svt_axi_if AXI_IF;
  AXI_IF axi_if;
`endif

  /** Configuration of the interconnect driver */
  local svt_axi_interconnect_configuration ic_cfg;

  /** Queue from which transactions are popped out and processed */
  local svt_axi_ic_slave_transaction xacts_from_masters[$];

  /** Internal active queue of transactions. The difference between
    * this queue and xacts_from_masters is that the transactions in this
    * queue persist until the transaction ends.
    */
  local svt_axi_ic_slave_transaction active_xact_queue[$];

  // Snoop transaction channels/ports of the masters indexed by
  // the port ids. ie, snoop port corresponding to master[0]
  // will be in snoop_port_aa[0] and so on.
`ifdef SVT_UVM_TECHNOLOGY
  local svt_axi_ic_snoop_input_port_type snoop_port_aa[int];
  local svt_axi_master_input_port_type slave_port_aa[int];
`elsif SVT_OVM_TECHNOLOGY
  local svt_axi_ic_snoop_input_port_type snoop_port_aa[int];
  local svt_axi_master_input_port_type slave_port_aa[int];
`else
  local svt_axi_ic_snoop_input_port_type snoop_port_aa[int];
  local svt_axi_master_input_port_type slave_port_aa[int];
`endif

  /** Event triggered when a transaction ends */
  local event transaction_ended;

  /** Report/log object */
`ifdef SVT_UVM_TECHNOLOGY
  protected uvm_report_object reporter; 
//`ifndef __SVDOC__
  protected svt_axi_interconnect_env ic_env;
//`endif
`elsif SVT_OVM_TECHNOLOGY
  protected ovm_report_object reporter; 
//`ifndef __SVDOC__
  protected svt_axi_interconnect_env ic_env;
//`endif
`else
  protected vmm_log log;

  protected svt_axi_interconnect_group ic_env;
`endif

  /** VMM Notify Object passed from the driver */ 
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_notify notify;
`endif

  /** Pointer to interconnect driver */
  svt_axi_interconnect driver;

  /** Semaphore to control access to active_xact_queue */
  local semaphore active_xact_queue_sema;
  local semaphore multipart_dvm_id_in_progress_sema;
  local int       multipart_dvm_id_in_progress[int];
  local int       multipart_dvm_coherent_port_in_progress[int];
  // Transactions lined up behind a multi-part whose second part is 
  // not yet sent on the snoop interface.
  local svt_axi_transaction pending_xacts_post_multipart[$];

  local svt_axi_exclusive_monitor  ace_excl_mon[int];
  local svt_axi_checker            ic_chkr;
  local bit                        is_reset = 0;
  local bit                        clk_observed = 0;

  /** Semaphore to control access to queue into which masters put transactions */
  svt_axi_transaction dvm_xact_read_chan_queue[$];

  /** Internal queue where dvm transactions transmitted on snoop channel are stored */
  svt_axi_snoop_transaction dvm_xact_snoop_chan_queue[$];

  /** Internal queue where transactions from master are stored */
  svt_axi_system_transaction active_sys_xact_queue[$];

  /** Internal queue of write transactions generated by interconnect */
  svt_axi_master_transaction memory_update_xacts[$];

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   *
   * @param reporter UVM report object used for messaging
   * 
   * 
   */
  extern function new (svt_axi_interconnect_configuration cfg, uvm_report_object reporter, svt_axi_interconnect driver);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   *
   * @param reporter OVM report object used for messaging
   * 
   * 
   */
  extern function new (svt_axi_interconnect_configuration cfg, ovm_report_object reporter, svt_axi_interconnect driver);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_axi_interconnect_configuration cfg, svt_axi_interconnect xactor);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Sets the configuration */
  extern function void set_cfg(svt_axi_interconnect_configuration cfg);

  /** Takes transactions from the internal queue and routes to the
    * correct masters/slaves
    */
  extern task process_transaction(svt_axi_ic_slave_transaction xact,svt_axi_system_transaction sys_xact);
  
  /** Task to route coherent transactions to main memory */
  extern task route_transactions_to_main_mem(svt_axi_ic_slave_transaction xact,svt_axi_system_transaction sys_xact);

  /** Waits until a write transaction with overlapping address has been routed and completed at destination slave */
  extern task wait_for_prev_posted_slave_write_xacts_to_end(svt_axi_ic_slave_transaction xact,svt_axi_system_transaction sys_xact);
  
  /** Task to route snoop transactions to masters */
  extern task route_transactions_to_master_cache(svt_axi_ic_slave_transaction xact,svt_axi_system_transaction sys_xact);

  /** Polls the internal queue at every clock and processes transactions */
  extern task poll_internal_queue();

  /** Adds transactions to internal queue of interconnect */
  extern task add_to_active(svt_axi_ic_slave_transaction xact);

  /** Updates memory hazard flag for active READ transactions to overlapping address */
  extern task update_memory_hazard_flag_for_active_xacts(svt_axi_transaction xact);

  /** Removes transaction from internal queue of interconnect */
  extern task remove_from_interconnect_active(svt_axi_ic_slave_transaction xact);

  /** Sends snoop transaction to the specified channel */
  extern task send_snoop_transaction(svt_axi_ic_slave_transaction master_xact, 
                                     svt_axi_ic_snoop_input_port_type snoop_port, 
                                     int port_id,
                                     bit last_snoop,
                                     output svt_axi_ic_snoop_transaction output_snoop_xact);

  /** Gets the ports to which snoop transactions need to be sent */
  extern function void get_snoop_route_ports(svt_axi_ic_slave_transaction xact,
                                             ref int snoop_route_ports[$],
                                             ref svt_axi_system_transaction dvm_sync_sys_xact);

  /** Maps the given transaction to a snoop transaction that needs to be sent */
  extern function void map_tr_to_snoop_tr (svt_axi_ic_slave_transaction xact, 
                                           svt_axi_ic_snoop_transaction snoop_xact);

  /** Adds all snoop channels to an associative array indexed by the port_id */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void add_snoop_port(svt_axi_ic_snoop_input_port_type snoop_port, int i);
`elsif SVT_OVM_TECHNOLOGY
  extern function void add_snoop_port(svt_axi_ic_snoop_input_port_type snoop_port, int i);
  `else
  extern function void add_snoop_port(svt_axi_ic_snoop_input_port_type snoop_port, int i);
  `endif

  /** Adds all slave channels to an associative array indexed by the port_id */
  `ifdef SVT_UVM_TECHNOLOGY
  extern function void add_slave_port(svt_axi_master_input_port_type slave_port, int i);
  `elsif SVT_OVM_TECHNOLOGY
  extern function void add_slave_port(svt_axi_master_input_port_type slave_port, int i);
  `else
  extern function void add_slave_port(svt_axi_master_input_port_type slave_port, int i);
  `endif

  /** Populates response and data information in the original transaction
    * received from the master based on response/data received from
    * snoop transctions
    */
  extern task populate_resp_and_data_post_snoop_main_mem(svt_axi_ic_slave_transaction xact, output bit pass_shared, output bit pass_dirty, output int data_index);

  /** Gets the slave port to which a transaction is to be routed */
  extern function int get_slave_route_port(svt_axi_ic_slave_transaction xact, output bit is_register_addr_space, output bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] slave_addr);

  /** Sends a slave transaction */
  extern task send_slave_transaction(svt_axi_ic_slave_transaction master_xact, 
                                     svt_axi_master_input_port_type slave_port, 
                                     int port_id,
                                     svt_axi_master_transaction slave_xact);

  /** 
    * Populates data field of transaction received from master after
    * receiving data either from snooped masters or the slave.
    */
  extern function void populate_resp_and_data_post_slave_xact(svt_axi_ic_slave_transaction xact);

  /**
    * Maps a transaction received from master to the transaction that
    * is to be routed to the slave.
    */
  extern function void map_tr_to_slave_tr (svt_axi_ic_slave_transaction xact, 
                                           svt_axi_master_transaction slave_xact);

  /**
    * If dirty data is returned from a snoop transaction and the
    * initiating master cannot accept dirty data, this task writes
    * dirty data to memory.
    */
  extern task write_data_to_main_memory(svt_axi_snoop_transaction snoop_xact, svt_axi_ic_slave_transaction xact,
                                        bit pass_shared, bit pass_dirty);

  /**
    * If there are transactions initiated to same cache line around
    * the same time, this task takes care of sequencing them in 
    * a particular order
    */
  extern task sequence_xacts_to_same_cache_line(svt_axi_ic_slave_transaction xact,svt_axi_system_transaction sys_xact);

  /** Removes DVM related transactions */
  extern function void remove_from_dvm_active(svt_axi_snoop_transaction snoop_xact,svt_axi_system_transaction sys_xact);

  /** Waits for WRITEBACK/WRITECLEAN transactions to the same address to complete if there is
    * a hazard.
    */
  extern task check_and_wait_for_memory_update_hazard(svt_axi_ic_slave_transaction xact,output bit is_memory_update_hazard);

  /** Routes transactions to master caches and main memory */
  extern task route_to_master_cache_and_main_mem(svt_axi_ic_slave_transaction xact,svt_axi_system_transaction sys_xact);

  /** Process barrier transactions */
  extern task process_barrier_transactions(svt_axi_ic_slave_transaction xact,svt_axi_system_transaction sys_xact);

  /** Splits transactions targetted to multiple cache lines where each split transaction targets only one cache line */
  extern function void get_split_xacts_for_multi_cache_line_access(svt_axi_ic_slave_transaction xact, output svt_axi_ic_slave_transaction split_xacts[$]);

  /** Processes transactions that target multiple cachelines - READONCE and WRITEUNIQUE transactions */
  extern task process_cross_cache_line_access_xact(svt_axi_ic_slave_transaction xact,svt_axi_system_transaction sys_xact);

  /** Populates data and response information from split transactions into original transaction */
  extern function void populate_data_and_resp_from_split_xacts(svt_axi_ic_slave_transaction xact, svt_axi_ic_slave_transaction split_xacts[$]);

  /**
   * Returns the requester name for the supplied master transaction
   * 
   * @param xact Transaction for which to return the requester ID
   * @return The component name that generated the request
   */
  extern function string get_master_xact_requester_name(svt_axi_transaction xact);

  /**
    * Returns if at least one of the element in the input array contains non-negative value.
    *
    * @param ids Array of integer containing used transaction IDs. If the value is negative then
    *            it indicates that the corresponding entry should not be considered.
    */
  extern function bit is_used(int ids[int]);


  /** Samples interconnect reset asynchronously from axi_if interface */
  extern virtual task sample_reset_async();

endclass
/** @endcond */

// -----------------------------------------------------------------------------
`protected
UC?YFRaCE:_^RAN?@66e9L^.FDK&-gBMZRH)ZLeL)[M6&-(bK<>R,)#gMP-5ZMQ&
#@9[0-O#4AGF,M75eURLHd.Qd@;V5+3RY[D4MNN(/PaY8&eVT=OVTZ,<@\.R417,
MYC-HgJ;&EYY<B\Td;Y7K@ZFP3R&&fT/1^(YPA/G\#SZd]JXGV_<.R1VQGg=PMUa
f\8g5BW#20^BS7;BcLIBET786d/NUTc8IDRB\HJ>OTWJJb.aCe4:6#S8c0,GJ@(1
24OgI4[:[C-)YCaF1D3^<S8WLFR9Ne)Y:3d8Lf>I1e\),c3GL=e(f\7AK_MI2U@f
;Lfe3K=51G#_b1S5SVL+N(>DN2&[+S9W>b5/6D13-#L9-02+Y.0:d6VNO<=O,&83
CBI?=f(H;;K:-Df_;2]B-6[T,9-O4cg=WGHW165SV>G_gD^?P4gf<gTL-Z-R+].5
^4)@N=T<XU#0QQXL+I>()L,EI^8bdU+RN6@.>W\JFEg.bQH:UK(/I2d1()B5a2-+
^Q8>RU1c_]2>WQ@^WB8dT^EM<GHRFNcJI_fP?/^1Z)S1SF5@0&:]EFOf<gMCFB>>
#W+XB,cE]:7Ec?e01)JMDR\8N^2\9;)VS9??H6H-\4<2+cM+:0,2-<X.FLc]]&a4
>?9&1KB<FJdgMg@_O@_JBSIcM+>b#7Qf1P25[.e8HfF\-9g77>IdI_\[&6905GQC
#Da6Z-50:R.5A>2F4QAQ]XBEDYL+IV,BeO-R4I_OTc:ZFf+adc&)IBB@8e_V=Qd9
X05cWEOT)a^^/NB&2JK7#b>NNVVS.8TOD7SSTU\^Y]X]<6F)NN#;PQ-L:XS@GZH>
WK>#K.O/DgMSgKAVPI+FYST<0QX^.D]?.Te<Y]eX0KP72+5J_9KMT:BH52TaPeB.
+W;6L>CUX>]&]DOR_S[cb^M/J/+=X6,WTce-9=-RK\_a3VEa@RCEf(aK+Y0,D?IO
)db(;O>6R8;W&W4Y_W-+DDFfdF20JN67fF+^\Vf6Z7(1C;0D5ZYIO6;[_Z3OK?CS
c3NF2bVcH^UQC<gX#N^DQ8-AbYYLH?D1a+UEVG)K,HTO8Pd[WU-S\[N&1RLVW:SL
RFJI].0A_WL@HXLb=.5OWXVf+H:4+N=<UHeB=+X:?RJB#<ReP1DHd,@&J94UPL@1
e8N2&R\<DWeEQEaf=IB[60D.9\7G&479KM>e#aVf<\>(Z15G3NbC0(&GK2D[&VOB
K<@<.NVZB07F8U\+D:&?V8&7OY+<+1-Jf?;@)WV@5PZ(/,3R0NY4(=_#IbG9F^W\
^X_^da=GLI.@RN7@E<IPc#G__8?HdN.&TcfY5Qg91;0Q5<g0H(cN.?aU6,C@S;:,
[a?TV+aagfC[^N.:69?0_AOXK0?#D^f(2>_<O;FT3TCXT/,C/JL#Y8O0MF7JKH>0
EWC3,AT,&RN(?9.)]](LA3^M4?7\Ob&UaSH325,;T_]?c+JD?+;6<7IV>0MIAM#Y
&c=-<86H;BaX=)Ue(NYfKZ//-D#/d_;TJY)J4-g9-<0Y;UN/\QGJHQ8\,/KL?PF7
2+R@0DZMBJ#8#53(8SW-?QV<I#AX&,Z>eIQ9Jb91Fb(KTMB=+2cX])SaM6ed5aRY
J8:S21P>KeeCW.W,bX6PV<g(=2.d#F1fa9=I@c/SGAOf+0(#QI(@e[SBM7R(;EY/
c)[ISR,Id<XdO<W/:3a2G)MU>PcQ9TR\G=NFYW,<C,..@(8V^MX79S:,+PVZ^>MG
I[S++3-^T[([GG]EbJ85]9WHKU9J,A?/E>+5LB9-)3C((S(--[Q^G\3YQ80=&DS6
a1B#8?S;TQ89\[AHJRaE:b3UE3#I2&f6A]Z2]\>>.fEG,123eN>45B-7NcfUEV#a
e-<NWK39^2+[=F3&LJ@03#MWU;NHJ,L_-6ZC(]c6/)4/PR]&&S,BU.WDOG0<1.1-
B5G#5+1;6A]5MI-LJ08EH-YDbU)CY.7YJ@4Y;+_RHdZf-CUA?LB+>EcMS1:2;IYD
_7DFTLf;^XKG9XGLWI7<f>EPJ?8JE)F<)K]O)gD\>\QB#-R2<9SOQ[IQ)b>;_G30
Xg.QFTV[TY+cH[8#L,7L65?X1Mc->/IfF1XYJ,./(cXY#_?P3O428FSe-G,V#I7e
PWQ8+4?SXI,NXILOB13d(/>=1PeK<;/f>M;a]e,d:(T.BfLX>WI^_P),<f3<90OE
=BP?.^SI[SfHW3PPL;158]a9c4CW)b?RQ;Be(B4&3)K.,:<-^V3D_KX:]d(7\?-X
?(5TSSe>^1?63IJ[>1=NDg7a,1+LXHI,H_B60NI<80H_V1@I-<030)Y^a62DO>MP
U)S]1c^<?]Z@gDW.Xe(K<UMbO&\gcQRDQ:9Z.2/#B:6/GU(@@(9W6ER\5[:U(RLL
V-S/gQ6XEK4#3K4;KgP.;BV_.SJK,;4,KLU5LgV3^TFPeJGP@YQ7DS^31.ZNBRGf
VZ_XP1EVeZLER/,=USY0]6_ggU>&AS^[PgNY4)0<_HT<\G7)-;7RW7SIP7&=?1G@
0O-\2N##S^dD4_[c=M1.f/Uf.&fB>C2e8OZc]H>7+Df)bf_-^LY(EDd\X7TXH7.V
K5AUWXd]QDOg/[)0-ZX=]+H4=EQ64MFR2YB=&eC87TVe;K8=W#JZI(O#6D4>0f0:
BdSFHD=X;)526@aU5cJb7\BPeRL0@MHJAHF]b4^I/>O+^3[5RK59=c]gMH;&GJR=
EM;@7PCE:)43L?CB_WG?)73Oc;8;Y:bYd(O[a-L<#@=Ac7#Z.-RR4K630OOQ/9K_
-))5aa3G;5/M4S2a6LRCZ^N4P37#TFgDJQKE&4+=4,A;MecWC3FXVb[#^=bSKXUK
9V0N-fF?YJQ(,M?#>BC.J3>-A)W9ERbNS(,YP-W;<aF2g3DcC(;eY&[U?VdVd<IR
AX@HLYOeTX--?<M?MR3GCGDHQYY=[KCNgM2EFFIgaI;dF44A4C&/+6_,OAZTGb(J
0EQF#(C6+&Md_?fPWCJSaU#]9OV,(cbZe#a.Z+TfJ<&6Tc,a=+#M)8@].RI37&Dc
=YFabO]a=NI?98XgCRAW;BF\WQ&</&^cL<3YBfS5?=.Ee3LW_K@VbNHSF\O;f\_d
W&,?3]g&DLdC\C=ddd>@5eP:.G9=_3X<,X,Bd1[I_5+-+=g=.3_X:JAA\GCX7YF9T$
`endprotected


//vcs_lic_vip_protect 
  `protected
HR_SRLeBUPEFP99BV],c]@[9b\7W24HO?31T(?V=QA\Z34&VC\?82(NA-^DEAY[7
8F#@LFa&T(89C?_(_IOYM/#Cb8dRIN)&eIU1JYHYc9VNQGP.@)5=AE9&Qc+0)B27
+,I,^\#bH3d#8:;V<XRDb0Sa6:M2#KXA^,2NCd7Z+,bcGXVUb>Bb02G+&;a#Y35/
6&IdYM9[>.L34[V7/,@68RdWB4Xf#/MUc3Fd[WfDe.K;3K8BKGORW9UAR[RfBgPU
[d]f?=:)Vg@-BW1OC=IM#P#QC2N:HA\edX#WZGG/8<<2UE[=_g.BD(B2NcB9PJ)[
#R(4ZFFVdK5CEOWJL_3-QT>1T3<b]]=6)AS=KF0g^.EZ)MJUK5T.[])4Ve4_36Bd
=QLYY>HOV.QPCXCd9>Z82NIQ7A@U9J3Y_+Mb:RNAO3UC;Q]6a7E/L.ACaK\SK2g/
POVR8VIH_6>/HJ-4aa(@IS^9O(YfQ-Xg6Z.]&AffG5Y/AHZXKEE#U.)P@2Ve(e#;
2e.9N38ZQ;@HKUI#-dS#^AZ.f:N<SKY,O22KcaD8<)aN>a^.=e21_@@<;9B=^fA&
1abgX9A\//HUf#;=e.U6JMa=e+6/a4.2C#N5GGQ_3_A6:SXIcV;NE1IbI.3#BU@T
e=08+?aCH623GeOCL<_WG;a6^6;A/X>=5f\Y:Rc\/1TV,_J7P5(AO#]A&)XaF;M#
W-8(.AX]UaP=7dD3<cS<8XYeD(U]:RXa#^N+/f,,aOYTEY8cMNFcb3CGgRF8K8[\
EQ9.F3;KU\3CX6/0a:R51gGN?6WgX0fU3;68E2A,CLX]<I\SZbVgbg9SD9.E>D1V
WVW?^168)g7Meb?2eTTI&39W41U&R@1OX-2CYZ7A3]FJF04_;O6[C=C#VE+(EN79
OEf_I).T^K6A;-A-PT;R8&(ZC&_(g]Fd7\5Ub;]Q<,?R.VJ^&;5MZfIJ0^/6S>T1
^2M@[BNWFY^bgS8DHB):a-/B;,b2IX70H6)a)Nf15F\Q1LgX?\^6]Ybe2LY<cIA9
Q=R01EPR#-?AS/LVHF3dATFa7[&Ec+g9MAF>_2;06-WXL.6:;g8U-NTU+9(9a4f?
IX&edZP;=MQ=)5fU580[B_A.?<b\dW48RPd2YI;-=F9D#5LNFb(X(41#O&MOAXH)
,8Xd,Q_NJVY)d_eT]JT:YZ0E?fCg/g+d/O[Y3=aU1+GTR+/=3<VT)#C#_B;)=fef
1,A1(HSfE.fP^HBA>P5VV.GbC.+A[4[0<c?++HHJ>dDWRL#J[/2DA[IaY2KHG4c/
S[/ROaW<-W@>8&7VUM?M-dVXJJRb1<E.F:f^Q=f>08^[XVL;JaJdI.4WE;8Y<_N6
:V]fE-.U,(7abQB1<J#D&I&P#P]#d35Mf]fA12Y&)ME-1=d6ge,=-FV9a3S;?\3(
(9:[b5g)X#AB4]aK(aD(Rc<K5JM5?9N.\\)_/]T9WC/aZ>0BHFbEab@WCF+gP16J
SR@VABa[D5&SbUa(.A-0=F9KD98ZVA-VP?CM?F6@_+a[J3;XI-^;]1K)<1Z(?:(9
c+4XI1N^<:<(#ZP48S+PHd(+,S0KYf]>>1,@FaYIG4?H9XVHD0eEg#e-f(P./.QI
GZ>SQKWQ\:J;)?[PF8(Gb(^3=baP\b9Y.2D]/P:VJO,=]5<gXeZ0eUAPa1^J7TAL
7RKX0<bgeWZD,AY/0>.-YOGC<ESTMHG+>6dW&e]:5VGLM^Ld1@UCY-O8U33DOYR/
>3Q<GISW0DJ3M2B#EM&___B[aWb9B(5P85+XUcKYc\(Ib5A^g;F;g,SX,(8,+GM4
9,6\7+G^J4#Lg1d1gO:(JY^):Q+QM?g<2gaO<:PTa?@2#6,.WT^1H-Ed6H_\V#]Q
[D8-;E1YRJH;<K.LME1K(;I:a>P5dPXV7).ZeO;FbSZf+.Rc0^9K[9_fH3B-TBbU
[TEUTXZ0NHb+aYAQ^?@PXW2/3#G7D17SD.[>]NHGD2[SZJQSaHBCCC]EX9d<-R)S
J8-L7VUfQA(dd8PX]WUWDR:3(;&@U-\)WFGF8WYQU7A;B#OEU;D\]\M=)<:SCS5J
YD)OF/RYf1N4Q1MVO13NHJ>4BE/eN[Q29&D/@0f]K1A0399e(ZV@TV^F7cX&N\_K
=1#6Y8LNA>cL5FfT3&>4+,Nc<f;F-JK=X>&2cL>\7eSg]_>^a1]J_K(Y\S=ZU1M_
W]3dB:_e@;VS0](Z51F]b9@\D1\EAK62f.O\.4+0R:]&dYP:0:ZPA/Y<6D6g<4[S
[ea3RQKS:QOSfI^NeD2-3egR<,PafYPJX=(1b:=YKL/9+gUI]e]AF->XD>I;eUAK
ZeVRK(b0Ua&0@?C_V1O93f47:[L[@>Y8<cL8)c?PgW1YR4.c;W>M.L4KO:3LKMB8
FSF#2J/_d_Cgc+3fM,3\4MV^CfFH>]862:0(H+DK4Q9[PB<HD\OT1<6g)e13QN(9
<X5<<V)(5Vf88>[E?8]N]R0,3Da/C]E=W)?OePJ+<7UZA/aH0Z^OaI0DUNRWL-1&
CGe(JY[.4+bQ3=g]<LD3@cJ=0R4->[#ZWe;0J9(4&QdIU?4N>BQg&O4\39EC2g6g
AOT-Nb>TWF^4-+]A9TaTZGXVNc&Td>LC\+W?AL[+Y-YQN4Y?dEL/7]QN.fGZV\b7
L[EU2-+#.Ia.BJNA+4KMP)+PZNCF0@->V#H#E_2Q,VFWSZBN70Z8.bY-4RG45S?F
6:/(.84+0:?:fEP._R(IYZFE2=KH2dS4+/XRe7^SZ8)eDSIJLFVc;gb.]<.OJ&/.
]@.ReTN.SH>Z>9)9)<<#JNI3EZVQ:5ZAS>L;2(7f76<=LD<[[[0NQ^:]W;NEff+f
LA2YAGZYA0T=VW3f<6SRA39#=+d_M<?T>D?1:Aa0^B.;E5)=&4fR;K4W5&^M&;I?
1H>?/NT7_FXU;PA-YHY<]8]Ab_?.4_XKWC7-_\6<7PeX[H(@3Sf)0dgA_5G+Q4CK
2/#9[76P7649=W;e@BYg_R+&OTA2(.163/T_;3f.EP[11GNCI2N#eRc77H<.H,N/
1XJ>YLNG;0AZ2X_0f7VeD&OKd_X?I[Y@&6g(8N]BF@AW9GWC]C3->c/4=MNC+G:L
<d;N;ESX7+1LXeC@VR9BVPH)-)>d\gf+/)#T.gPNB.YK@/>P:GSdCN5YW\UL[e@C
cI11e,,R][,Q5Va@MR,^Y31PF._KE#<Bd_)\egUBHTRYDcZJDc_a@g^&C<D>@?(;
16FT:+KL^@./V626Q/L4,.-;8VC9Ebe8PZBEUX+PWWa8LY:VMW;.5R[P>)3:9f/;
AGU_AL/0W:J8DF0/OOP2.#R8S\.+FP@WL#Ce(D-<UCI-/_YJRRAfQBa6QIgIND[?
Ygb@K1-(C(YacD&.3NBIRM>7LcY+GM68N=H^2:TG??Q\ICZYJ7_<eL-O09&2JfS(
KGA?Hd5NaY;XV_V0C>WZdFG,>4)&^<bV13,A.2].)=XZ(cMdDg;V)8E:WLWSE7NL
3NUI;PYP+dF\)-.CU;@c<2JE/ScFIH\NR3CZXbQAHX&/F;\QW7bMcdNTf@.bcfQc
G,:H)3-MQYEW40F=XUG,>AbD:TJg8):<U.=fKD0HRQ8&#AbR<0E.WU-6VPC#-UY)
G-I^-/Q@Rd#6Z54FH><)=2eQ_D9(.9+MNZ:WT]R.-GR,&dJ(]T5K))TW.LJ4W6]B
bNO__SH=XH<c7.Pd\[]::.+[aF-J:bec_FCUV2<,+Pc_]F^UE4Q2;JF7+U;e8)a9
#@]VCYK#[7U-?3X96b3fY58+f^P;7-&S3#DC2(\g^RWGge8EENN;<Z77\4Y[OHO7
+:3Q,+82GdM43;;9]09+&IOY@cRZMPANc4>/7Ic]FXTO.^-)F8e1UE^=eEVb4DCA
_V^08g0GLA1J&N:>PET/f3dN6XW<#fYY_)CBP3_-C@4QO<#YQN&8HgfI5)g?cC0V
YdbN>HQMcGKS5KfeL21_Q5-DCW]5&3>BSTZfHLQ3Y1O#K-cBAJaDCHPKU&eSd[-_
_0(gH_EcYD];F4M\(9X&cb.,E&ed@eM](MV&(-Be5+_Jb8#E_B0+Ec4NQ&Z+E)S3
g&?[\M32,9/gQQ;b3L=W0cb@XA2QN8R\YX+fLbG1Q2X>+W\8;b#abSJ+d)Efaf:K
=A/KE)b7,g6)EB7=/E,-\9aCSaA.?0f+U=aCUNC]gDVNE5dONLRc<7&O:;Lf&egD
WD2U.gDg/g75YHVG-XFSebA=(36\46fHd;GK,^aY_&Z=_8XPF>.EXX#Z65JPgfO6
IPS_\BS?/XG6S?<a__1I(V_-dS4#@0Q[RENKER&:PLf^eC&.3c)8KHRT[eDbePZZ
I/OSfDZSOO)CbVPT1826XWT=^GLaR,(_45908D\a(1W&IgTEP6+gN,b\FVW-Y[dg
Xb4KH0;L?(:@V9H=\[LGEJ@\OX>DB/Ue2b@@e1NF>U4S\OT@_KJWgO6-]N)NWFQb
fTc1M\HQNN&cg/?R8b(C@JT?^Q1B^e6F134VZ,?HSO+d6G>faAF697/-:ffO_[b,
RHB<_YSeREEUcZPgACYRce#6[NW:<H3,WfP]GX:J6->/a2,+5.feQY.dI1gD]a3D
OG&P?XF1M#30(fCK<)].^@E[K2X^HP&5\])48GA[;13R<Q1,<8?&)F3U@23AH+?5
/91S,=\N0GC18e+N&SWdS,B8@22#/B[OK7^<Fc>:,5O+84\U.S>M[eO0&OE.JfT]
6gC?L7L\V+@QP;\<eXTG@\5@EX521Q_Y])/.]YTgY:e,.L23XCWN&:.:6^3eHNF0
Y\6HJ5R=[O??(4-..:8(f]FF.9(b2DUIFF,Q\8&&H=GV@/-9VG2MaFD4&O-CaEEd
59:=^VC6]A)7aQgYONg5=O^RAO5;;d8A/W.5A9.CXAQ,a=UY)/+MZY<e\Ze\43e^
_7&?5#XOcPY5+-)Rf[&D-_cf(9,MVERX)YG1N3.7d:FB+2?Tf=Q2:.#8H_VY++#]
/2QY);+IFH/8H\dAPKL_BZ8A,;^ZRY;42Tg6f-(Z7G\e@7?,FZc_:-7UR2@3+F3V
(U3/,C?TZdgTfWX.^0,,(HNY,a4ZKVda8OC]Wc7XC;TL)-Obc,4<8&Y4=H(SfR+F
:8AZ,FSSXbg5E0b:YYN85;H>DLg/,IeXbI:WFQ-;[.RWW)GN=d@()7Z_:bY-F8/\
bEA/N&;3U3DV4P-17Lc&C&>X,483JM>fASA2]=Pa=fbGRYK<EAI=]\dFdP(adK41
e&=:+LJTQT&AcR2K#Fc)Ye(A_0=\K141][3@bL@0;#c<[E0W>LeXBH+QFee+&9G(
-dSLF?FEd7\8gGV)+(2@V,7]Cg)+AHEPTBVPD)0NUgET6E<bR0@).->G/N3OT4a&
^5DP/:ONKc2^4[V2>0P/3N5O4+G2E0/).eOCQLN=V.=gNPBW;HCIS5&eWJ(E;W4b
DLLb2R_D8T(QW1)6MH9gOJ((2UX82Ba_VEL-VWW=6dW@KP_G\:d^1])KHZ0NT,8a
JfVd=[cd)c76)5+U.fRP.f(^>a#KR_/@OVd6;4E42B@;?J6(4>;M(-UJB;3D1:BQ
WH8G9GW2+T[R@5:=Eg,Nef^73Y)S(>11R50_RODg1F+Da[e2BGOIXgUJI$
`endprotected
        
`protected
Jde\>=eb3#W/K,;]1AS5)YR9M4PNJ<+3+VaN&2QB>AFG#]6YV0:P4)Z&XX3U1ec>
C[=0SBV6(+\TdK@OABEcb3M3&A&_\P7+>R7?,66CdOT(T:cM[FT)CA#Qc(86H=\8
eIWC4FHC[da6eSZW+7^GREM38$
`endprotected

//vcs_lic_vip_protect 
  `protected
bNVAUb\)7gg##K:J\eS21fIJ7Y=9/G9,5I(7<5d31KBN=-<-A1Ga7(B.La@Y9+=9
?;\/C=P[e8U+NY2_;T6\_/_K&&C#_O[01CP55#JA5#1:-VQeDVF;P3?MJN-[&6_B
Y+6WQ0GUb]ZJ8:D)A^eK_N9E4TKAf1@&F+-\X>fdTcC_7.+;&a>NI5.4&-D,_FO:
3ADgJS#?R3Oe9C<aZCF09dB550@3G66@>+=&G+1]d<.e5:B0ST/:J/g+4.A)O/aQ
_MFKI<^\)593TQM&[8?;T7LDggS18EPfDID8+<U9DGS^gIOc-bCcX^6&310I004P
\@d6U&>gHZ.5IV>PE0B30\GOD)?LbT5Tg=1?cC7A^A@J_RBDL>a=\F)ef=<8O3(<
9]cP4bB:INW0@L@](2\TaH><bM7SY#)<eALEVP#.5GdO\I>HXUIQE,<,8e8UfME;
dX327_188VIE_C@KE821,Sa+9cWa.J^@>53_&^U0@HRdX<6(GHGKB1>aT)]J\Ogb
#+NTR[a_>dB_RZ/8Xd(C,?2QSMB)OU5R-a5&2)c9/J:aE7=@?R&FY2;[#b>gLT1O
SE114,b;VALa\.BP[e+Q5A[)>0EE15^g<:L7Eb2^M<(5(aH]47cV888)E6X+)J,8
=)c3R0a[.7/(14P2dFdR\ZLDY,STSLDXG#/_#_>a4UO<Hg47<X&&\DP>5XYBHQ(J
aGRe.3WDMJ(R:]cIJeR/[OACV_FCcYV:NDD>g)7,CZf2K^-7YR25cAD-\L#IBUOE
,e@/8L&TJ93N)]TT7#S?V->-5,/d7[U\#3)Bdc9/)RX71]dG(?;XL)H.M2[Tbe#O
^,dEF<8&P).O1OeN2.[=4+-bOJRLL#YW6\YH22b.J_\QfVWX<VQ&N.Vg+8#?4b,L
X/67^=AE&D<_Teb[RP4\]A7N4K<bdJN@W9H^2#fOP;DCWP/:7;&Ca4[=XPRIK0T7
D]aQ]a:YF+e51,<@CDD5ZQ+g+TX[II^=JVO7):ZGPR/9[E0T37&/VV4(JTICT_#+
V)(Of&?W-bI5,/ED8<>8A9.beP#We2@Y,4>/a-A;)8A3V4>-2^U3FY,W)RGBL@Tf
3CZJ-QLdBdGF860[T^4F-5M97ge77eHF=QJB-Na^1I_g2(51=_#Q<EG)@LXY??H0
.g\gHV>]Ac&R[8Gg(&/3J.aCMB,:)fK1CFWQ<:)\^=/JdUH48ZfXa?V@aO[A&&R]
]7QS-QKfON>C8c0^V^CU>LbD(Y=_@f1DTgcUI8O8Vd?>&;:0@eKZ26ACKVDPdbfG
dYe\87Be0LF9/1/fQ?CT9](J+9&H946(@MIQf<40))=&O>1:)Z:Y-O[X,U7-cS<f
\N/),M_gY6GABD/8,M[fYUY:=dB=>_e3W0#PAR1a0IbSFYZJSH5^1Y\gZ\OBQ5-F
)KXU)Bdd]QBL3S827dUc8#<53-683[@;L&HONfI^aZ:ZT-,==<DJEbE.A0MRLX0K
;S<K7@[Bf<?J5R2^c8&)5J]<2C&P>E1)fJ&f>9H6B&9[H+Y;I#;GD.fETA.AKDHK
HR@cXAM:3&AMHQJN[URGLXA4U&6[CWQ/]VNG];F48dS8b<5fR/]:1/3MNO2?Y>SD
#;JQ-TQ2TPM03K+e:F:YM<HDVH\f_?T^+J+V_Y>I1GXHVTYYDQQ)dF)U2PSbTM7=
b[)K<=#VFCIa27SHKGR8H]cPF;)8LbIeNPL19O-Z<EU;HAVA_)ebAV\Z:=UaXAZO
T_WB5W14Ef?-8>2ZENb#?YP]&6O]_bII6Dc6(1+5C1,D\QC2W&\=PKgR+_3B>Q-:
==U4d@QFI;]PC-J<18f-F7g2?M1#V\X78Q7-4RS6gTfOUZNFZ5JDe>&g+f.0+8K7
cO\7a7TTac/GT0+&b)3BUJeBe80A6.MAa]X1\.#<g\J.g\bY.96f0N=6]3\<7;G@
0aR;(5eZebQCDDWN9cHBRa#)f9_\_a0WBFYG10RH5?FfHDD>b<4MS;]PFYX8@#a;
VV667\>\<aRA9-/.Q_KY?bQ&gaJX[?7;ZdJL..Ba)b?._UF8f)2/JaNHBPe43L97
;9Z^2#2gbc7Z=-bd6P4DdW:_&e=TR;;CVCNbU^4+fY?@Z=S:G8g#b<^QESNP+J^\
.0a2M[A=T^4D/(L]BfG0=M>\6;)M(BAX\-GYP6gXMb6/V92H690g\41M)R6ZMW#K
N[B+HJ(eOP[#J)WSA:gAAg0SbTJ)95<=<\EDe>,53>f(^.UHB)a#1CG1fO0IDD;b
2<R\TV]7IV7U[-L=2P7SgP6.1?NMaMTIW>8&HPKU5K14?#)5.UOIE2\]>ZL;40Tg
:;>[<dgMZ4ODY/93?:+X?b<C^_7T)9&QPY7\<1>@H:GH9Ug.XDM52:+V.G<BaBD]
G[Wba3A>7?NM:D4_G=aGGP:7]MbD>:9F:,XKe;g[cF:[OQD#X)=+<?D0c926HBO^
E_Z?J^Rc1GA3/[.0N6g&VH-RR4(#I?,XTDAV(&UE#1X(+_,K\@EN?,a#:L@1B2Ec
/>;];V3;H>Q5@\K;P]J-+WaR[F\MNZ?3Q?U/DPcb9SX;O/aCNAE+gBAQ^F909BcA
D9A^RW7U9SYHRLX7HY]W^MZTEVI#Sa)3f,_(ONU(HAQaHOdZ3-?Z(@/]YHW;.7@J
d,OE/eW3O_bG:bN\/W5BdO^+P/.0_a,0:)[)<6B3YZ]ASW0GBZ;TQJAgZ\91CJSd
7P7ZNKK9Oc)EVM7L4791DIgAc96f.g^X6N6#SH@BFJ9[=?A?C719HQ[H5ZJ)=T<V
eg-0Xc[.bP,WJ4W?]F^b[(&Oc&9CZ9,W+)-L2e&7)#;_3Q=gAI@+UIa+NKM[QX&5
CMAJ@fBL;#WI0[9?2e5:XS<GeSgUD:D+:RE95^>U+OOB_PSKI_8F_@>e1C;VFJ,1
^[<3?FcA:/@M-7DZ?KBM;L^35\a0#<=OeY#-a76#-8]E5d0eI>5.9RU6)da(aHSG
&YNMfEDZa<DG@>7W:665#db8g-8K:TL4R.E#V=8L9^\]7.6YXa.OJWgLfPE)F(1G
G\LN=L:OQVO8W\HJ[DW/\J6HENG@ZSQUW<&5FJNTBLI+?.a9f&G=g7F=55PVb7[D
2^)?K66A#U<aY?fFf5PP^\Le^fDU56GZd6\a:[30EU._cE1#+#EJeGUUK7SMIYI;
/eN)d26ge5g+Lc/G088gJQ^@;=8^6X6(C)eWeDb4<I;@P<DGJ^A\M&J5P6Q[I5DS
c@O.16gRYOU0g]?Jf/+Z96FG>Ib5D\#/95&eTRVO^QT7M#N5-6DGP6a:XI+3;&ZP
FLWEAW20^4>VUf=BacC_>+X:Id.8D/SCcHT.Mb&@GS<HOF]Y5YLU-g,C#X4_&e@C
@eKKL)7KS34I<^VWV5N5=[7JC8,5g/R_FEEAZcW=fSOD5gSS:<[Qg[K#.2IfXE9T
B,7BgW<2H7g^81H9a6+^&T^PeAE7NDZ_BB@fA0Y)AK2->,YTK?4L(BUQ_#eNW2E/
V,VWG>:(:5S6YU4\;8FPJ[Xdg;e\=N.,dR&LAZ8;Vd:-=0T,NaQ1/+5)d?9N]T)a
6CdZ.ZNW44\R1&-=AY(0,DEU>\]\3RJ.1;WVWRS5M6Z@ba1\@FT;CE=<b[5AF@H7
#Of025R^GC^X[)I2g@J_4U8:S)aM.;:5dIY30,QXC9471Q5dBW-eW)&KBcY13?0T
(I<E5-&\D#fK7Q]cQ?VBdCd>gVC2GZAQGf,fG(OeV;&g^:F?LD1Qgc5?H53UC8_G
?A#\-4)#KM+IZK[:/.g7;/<)Q?Q-bX,09OO7NW_MKdNU6:@S71&WcB9e;M45bJ\:
c_Hc1G/.MN(?Z#OW<,]?PYRPGSfe\9)U<LOVRKUS/NaF.-N(Z56P<3Y^I63#/::9
GX/FFXgJWYA>FE0\6LTKZf7D#BZZUMB,^5@c3<K5Q6D)3<e,Gac0aH27_;?&.O(8
(]FYPO5U=4N?&[R8WRD&Z\#=TTUL1O4U->NPC]bcV>]L#GQ<e.3+c-gbU=M:3\Q#
egRbU)SM4dLD;CgLIJ&-)eXb-VTV8HdZSB#4/RD-WJgSG(b[8a[LCZ=HM-c0F/(P
=KWLPOS\]g5^cQf;C+UJU<I_CZa@8NW@Y4A[Q;/J<<UQc6KQ&?=_,)G\0C3?[PAG
;7^EH;.>=<W68&d7Q@,8IVZBTaW2>>7H7.g62=\bRJMF2&#I5N/+F:X)#N0=?3Aa
9Y/W3g_5Q,aIG<[3gX_>2C\99gK]&#?+#9G_)?#M6(VI9Qf<RUAK)J\N=E3aM,89
H1N/5G.Ib_33[-/7ROWL-U3L1daT27DfdY;I0B/(?8_4T.J03/47)_?457dS-@>_
f0/X#B2@70U35]9:81,S:0RTAUcVW7(N8N+5^PCZ(DWF2.HJa)(:XH-f#IZ?L.6Y
.]3gW#4@J)@AK\^2^8R?c.P?H-eRJe2[5X5V\dK)LRGHYSSZ_BOH]DeVP//:<(/-
I_6KXX[>c5=]@.Qe(;MISSb,B(^5GS9D\=F:H(OP:OeQ;?DT,R+#N.8[YR(_/8KP
H_5W,FM-W1@JWXN12aA2,38/g3P618QBAMCU^fbbD@W72=2/6-)W[RP&ZZbBZMTE
,F9_eOPbB+^PdZg@D<A6(]V>DcY1Q,4cNg]g+0WS6ee)#U5NBE19I,<=:<.+FCGe
_MN:f>Q6gQNZ1HcFB7-?W/ZZGfHH>6@0YBHYD/38OgLYID-E0(8FFGXf)T2WRB1(
LVSe6R]9-eNF/O9[QA\=]#>afd9_7=ZUaUB\,&:C#/<-@Uc\gYS.C=VG_FgdKA&C
H]C5CdZUbA^]8fMH0=E724,FH>Z<RP,H(2<G&U]T3cRPb=H^P,<#O8(C6CIeT54/
afF?362bdK@)Xe:ceVIJ0JX[07b1R3/Q:;D^acE5Q.(_BQTU0U6)25YN^XQOFMWI
<3.c:WgND]cN0L8J;)e:SN&;(](._)DQ.#+e.P9FeeUVSBgDFCB+MGU9&?HS@W-V
^<ZO0&^SB\48P)AXV88^e^dQLS,S.?WD(V9L).Qf[K86R9DZd1N,HXP_=US+3=_7
PI8g:7XT_)OK1?#<:9]]MA6>P6Y,Hg@)DUV\J9&OCJWXY#E5E9f\G65@^aae&Nfa
=<cc,77HR;1_D)Xg\Be?XXB6T94N93>8<#8Z3-SZd:U6e.8GdO^8;[<,B_QA(1VR
]NdA1XK_86M[M)FF)C9eE.^?O=c(U6e@\:QS18<N1cdL[2,TW_Q^JOO,DFU\a\-(
-^YRa-3S_0<G[O74a5Re<1-f>OF3NIK2d0[Ua6>LZS?f^0+ZQP@\^88M-D&U+c88
_(=-PeX/P2D[FFP7V9]-T(;,SEC6(]GeMRG@T<F1Q6_6XD=P=@V\+<NJDbYe--Le
=X6a(=c+88);FC9Zg-ETcW9V[,_g&A=dVJDP4#M@<G\JB-TKdPc:+^TCM5@N,=Zb
W-)M9N=/4PCZT-<]a(^Z<;P(f2//fQAZVCA32CAQ[K<HXOGD,?#9P2221)dS@QC0
dYDB(@5M#YPX69@9CWeC=^,__<8BF&dXES7PM5]&4fcEg0e(g)5S4]&g\f2CBBVE
4bW-TVa=M:#(@<RHRYJNQ1=+Y:2ea:K199A[S;.+5\&EdVUM:4M+YF>XRJKS)dCf
]3XMMeP:8P_;-H4cM5fNMAI/<)J[RECXAMFW?0a2aTIT#V,EbU8H>QVWO\J[TdA,
:eY7c4?DQ[4;?2]]a;S79Y4+.0A9U2]RL],BA#?Leac5<LV&[;7.Q?FZW^+2W+TS
80+BI?+(9BIe&6g0-6F&23=/UW/[9\bY3dJZYF@FZKV&EJ5SOd^V?@CC5:Fd=HQ0
I=6L_[5<baM8WD#S>UKC<BUD:\P[KO6-bX20U[JGM6/_e]c/Te>@QJFMe92,72c^
/Y-3c,VJ62@aP)-36#A3ZZ;=\O#2^4ObK;48C1R-D2E_c08eA6G_f6[M<cX>,J&5
(<.66J>3<Ng;)J(JZ+.GgeUKE?TZZ4YQF.Sd\1E:BeO8Q,eB:9]U?<1YIeSS/YaO
f,0^Nf?Tdc#C:_,+M=6-JVgHW/A(E6)_1#5^ZX]P,gY]Bf,0D06T8Y8&X8f_]Rd5
f4bF;Z^6OJ46Q]D40(=519EEK^5Pa_CbF,EY+3OPc):0-W[:8HdXQ5H>._=5M:<)
\<](45J4X<X5Ic&D3G3V<A-5<:f1NbG&=4N+;UNGg1+)&e>J1+61X-,C17A]bO->
#>fUQ)f4A4&=a/f?62e[RFDLL<]PdT?+C^00\X-7A^e>;CCWN-UOXXT-P)M6\NQ9
ZK_>ILLN7bQBIQO8N.:,\&\:7gXb&RFC<10MeF4K]V/3fW+UfQ/)07;LU/fJ\^+;
/b@eQ9+J^0S0@&3B()fUPKD0L,[KMe.,Y&F^==JAP#=>M;^C?3[LdI8&BCe;NSa8
ff<Y=DLeBX?Oe?1>&0<37?VOe6P1J6(fRGB0]O<dR3A#=L:MeM@1J2(/.Hd=5BP.
a3;O^?5Y2F;6LSR1SM#d5R6@Qg4+W\M.X;D&eb48U:_?F,a[7fHY^-&SD+0La>ZA
M]1O[[IWa73/EaZ4\a.a5KW)R]@Y2\bgPQ,5)X(+2YQF:W?,WE)CQ:K\@K6WP?(6
S05>XK60D-G8JJRd2_NF2_XXM9CK18SVU7Jg/eBK[R@V2e)3Ce2P^74MYc(dRJ&(
g=UcYKHOa?&dF6T4Y4gEB7+7HRdA/X-R.V9OX.],^)Zd:Ce)cFI:S5J,,Y.[_V2T
R3bFcMZO&XC4UOa]-0XTBeb4&?R\6Y^Cc[[e8,[\Ie)(-O#5(+:Af=M2f/f]AZG=
+<EIXSYDaK_]2T=9)MHe1=;IPFI\BVT9L;^:N4;N(]c<ICCb6AFXBMY1&0X+0F[+
Ae/@SL8+W;K;Y95LO.6<-b(Vd?Pc=25PRW6TcLY)@HJ8<&Y(P?+6+)IN=\[X^@ea
\f\I8b)Q1[(KXO_,4b_W\T1cGENUT07GfG,S20->d;ZJ?#3aSAVZCMV&,cHD6F_X
UAM/_YB-4>VNA[0/]ObV#e#HIC\TZHeD7_[e?N(EXY1PZX-1]OEJ25W;I\]Cb&5f
B.CfBgIITFabJ,Ig3TQ;XegE(F5]4XPa0?V;HME</Va+WbH[WE3A1?94<S=5c4Ob
60edKg.aO-BB9S3b5H)0;_C1DU.M7C6#0(V\PMWN/CI+][aE_S#BTabZ8OGEV6aK
<g^;ZAUKK+X3GU7)=D8XOdI<A/^8A1a8:E:^PJOLO_T8>E.(dIOR7gIAQPTG?#DH
WD__Te]gTS,+HX=^6;fT.5R\-/S>_U791-,HcX-M_(R,XEMe_PO59MTHN5V\MX-O
7Fcc\AI+ZW?4+02BB[S<(?\ID^X=a4.I?4JZ.IRAfY=W@C&W/SLC7+#AB)PJNN0^
)^:)9A:NA3@=Z90CS@2AQ&[d2<Se+(?Y.e(9^KUT&Ke0BMQW>Z\<:Pb[7,[S1;,1
<6+N9Ma([,W.-c5b9D(&U6,,UJB/Sf.X14ZTKE>XE21^2\<54b=5WNU#ANZQ(2,H
]Y.acG1Z-DOaUXEA2ZG13@<6d>f9fe)2?((.\GJPBWR\P2;0D528E,c_TD;>T0)c
^/CX0#W,Q,:]3NWYb)U>)R2-)B&8>1T]DgKJ5A@KEX5#(]\F#8VK.,,DBfD+UYI+
,?VC<78I;6a:DA?+J2JH@5\U>57;/5R>)gJAT^&8(TaFc..0P1;-Gd5.eU7<F26S
A8TG:Y8/H@2&40A?.#E./F1]Z8>eBA+?)U4)TGDZ0fS73E9eV]V[faXgLf)G=#b2
5HR<H-G=/LSILP>Pb+OLD60#B3?C-7a)I,9CDG-e.C9gG.2JCVJWVaP:6Y=3b5]f
]:aV/T9gVe0d_4g5_7DYW/cO]DEMeD7C7E4[,LW#d(AE^QWSG/Q[Lg?K+[JZQ[ZV
a]4(>#cOTQ#[746Z+b0f@A5:1?=240@\@.1M]cL#E>)+:?Sc[EOIVPYAd]4;8#BF
2C3Y(-58#K,O9MY[#_5<-A-A,Z<&+DEKP=>H<_E>@F>WU2Rg4[dILe]&>BT[+2+#
P],ZNgb62+)YI[USIPHR/X[dL]K9J//#gQESb/=H]<4CT#X3A+<SGgf7?0]D5b6f
7^2(O=>b@3cJ5GE\3ZH(PYDBc@EgBV#gVe>^Fd9N]Z+^E]]c,RN.Z1R+DE8W7\ab
gZ,=cIRTVMQU_4HgDXQR5?_#a9DU1fU;cPRSZf[OJ>8\>,6F;52U;fcHSZ/d@7DD
.1NNTBA6afM<;R^H)B&GgM^7Q3/7Z2O>(cBMQ<W7T]\UHPPT93\2;W?MVCNAN+@D
^;.67aS=VZ6X-32K#MKgb8M>V?Y)aEbD:/+7A)e5MH:Ea,EW^XN84C<MTPXW9L]3
Za,[d+OW0_30G\P4NfWQWa#+3Rg=:=@S.2/S@ZPZ0O32R,[@Z<W:)H?G4&X>&#eC
UT8RC,A@Z_&;\_<I2],PSe5/&3=&AbT2&7O29^9f(_5&<,G,L3N/=_1g\G;AW2@I
]/)#Rd5YEXIAVA+JX<e0E\&^-4;#7#BcGT3+_b>BU\=8KV:HOFbQZ-(Pc&UR].&K
-E_^U)(UZaBD[@1&U(gVE,A<agBD#W6fPOaWdd4d-BdJ7WM+-O78.D]PM+gTd]C.
d:4DYdXF8&db8B5c2@+_?64>H)fWe0,HCPcCKcZVRYMNSG]UE]2Y:C;<A4cJ5dXQ
#EZcM42#d2A./;UaNaCBH-_&dc_-a5Q7?A[RPeV2VV)YMDE4\Y1Mg)R^OTgRV&RC
WCHegV4V6C\cS+Z^UF_6SWN)#?LS;#E4N)VDV:F4PI<,XW+N99<DKKOU).N>3QY1
U5\:W7OP8/1,cZ6B6:AK]L76^+Qgb()9+ZRU]WJ[5+(R12<@Xd6:E)SgC<O;#V4-
JT?e/+B[K+4L]6^(P##5LZHD(_Kb^f#>.TQ>WaS8ceeac.E5S<4^Q]87+BQfF>3C
F_K)[JTfa,<RSXF8CSE9S^C^/e7=AgOG#=&G3W?_G?b(&],NJ_^-;WPBS#]C-IC2
.?+ZO1&2#&>PV>/1Q-+&OCJ-aF^Q]4RRN&4-#1(2X:E#c/O38VGdV/,@^]M<Y1\^
C:f;G^-/J@gO1C@5#.5R.KA.6[:8<TVF0EI4,KV2BJ\&KO_2.aB@HO7B<O3X1P<-
5^F+>3[SNST\<FaHd[=J\ae9:I&VH9_6V8/O3M2?=>/U8]b3FB[-][]I</H7?).\
IWT2NMZf(TUgAf?2X+)bA^TI0M^bMQBX+4H4WdOff\/F5&MZcEF-<8e_U:[UaF?5
(G/X0(<PTN_&[0W^KQcBY5-J,JP&L/CgOK-8,-PVN5aEX-)9DZQ;+JAST;ab4>[F
dC[Gf_I:AFCYW(<)X9aMf6gAMO#N-X&\+&+0-]=@6KMQJO-5]bW\R,eb6?0?#f9]
eIAfEPN>[J&[WPaNH]RHdT&D)0)0Y^L[W.8c>91HC]&/<E,025QE\X:E,@TF=S6W
3M=e@9^DP=RZ9Jb<3TQ+]_GG<N[a@G_G^[cJ9RFa#H8/aKGGO@XW@G9Z.J,21(af
3;S]P7fY,B:&DbJO4G&cZ5.&aB+#a09g.0)g9(bD@7f.ZSe^G#ACTL@,<MNO&#;Q
a3+3.OD->eC2WKD/J\LF5?:L+e0M;B:a(+b7N6O.6;>6IPENcG079_=.-JE9)V2<
+gSdFP=aRV6F?KbVF.7OF5RJB9L#=]eN.3CJc^YCbg0,&@geH>64c];?H6=BK<W&
=SN.VXIW+V42^WLa;O@3#G:aY&-2b>ZDOEcQfOHR8./>ae<T97C+FBX5Lg3c80DY
/ASXPLRf=AWbL(LcY<-;4VW2_D]cXZ8<gZ35VQSV6<+1N_L4c?I>JA7GIT_QQ[c3
06L/^Ce1^1Eb2JF)35#MMXC5DI#B0[4NF#gVZW<,E6b.SD)V[/]J);7X7c?-+Z:7
@a18]>\X,R+#)MB[RDREW.^T0I1[XI.1U7C?aa[Hb+9ge9d@gYTX-XVXB._DQ7+)
e[;NPcFNY;5<I+dD,fV<03BBU(Ec=c@4Vd4BTZSb-RJA8:BM8g4]?NZLDaWA4BO#
F6/[LQY_:f:F8RJ)d+f7TgUc])+gN6dG;+?21R4EVWc@f9NBQe]eU2UYVIA8_BQ>
RP>5TSb/V2X<fUI@:DPH,#8d,5T4Z2(6gDE>I0T=TV(<[1Ee+bA-XP^F<;C6<?O(
dRb\/3^&MI51KC_3#+A2MM;Fa>SUGHFeU[&H^[Z1#H9Z&TR^a>S&I?S>5T\=0YIb
W4WI#1/(WH=[(b-_B)=WR]\2RZR.Xbg9F0S>41F1:-d#Y/afK>X:e?83bGX_9+DC
WfWLc_BD64D&_B6)d-&FcGY4XO=;<W#fK+C;7-6\bOPEQA/ObJRUdJ3IF6:/[\U[
)RXU#&=I/\3041/0:(VXNWd>MJ?X^GBPJA@C1b683VH-)LD1,>(3K-2,UI?.VH;<
[Y277)Y#LeB:S8\#abZ/-+P1V&Q->bV0(DdEfGc,X/\.K@;JJ)=Z4cLT4GBJf#e2
?,eaI-A47UYA/N]D.6DCS\-7YP=F>2YW:7HL2ebHaOQNL[D>5;b:<7)HNAfG(IEP
Gb82(0<IdY3=fU3A1WGRf:_GT;7T]ZC\A9D0O,KYGI8=dc6Fc9dW/a6&S)^05PO4
#)C2c#4b8fGO&SJ3QYB8[@@,HcRe-_A)/_&KZ09^aW,MTT7:_W3F.O@][F)Ga0D+
PdD0Fa6S7?&Q14?3/&;62RTS\_#gV4(K.>1,7RYH-b;[>7X,CT2LV:]NYG^8\XYQ
FfSI6FbDXeS95]5gbB2/F\;A+dEPc)?c-?>e=I8bV:Sg8=K;Ua6O3.&#gRL#a4W^
&&V^@&:Q>K<;0V6ACVQNa)(P,)c_-eA3\bP4DEGg+-a\f>:4;Lb1Y9QJQ9cE/A?V
7A-ac^RJZ+/@,ZJ]KA&BR,6I47M78@^09DM,CJA<f(?7F782BNaV\-f\[G=B../F
ReT7<)C<#BA\W1HRUJ]S_gMU;Z\1^F77K=)VY(M_]Dd;.MfR4QF\24e:_aLO@7[W
YDCae2T3Sd2d573O(5&3(2P>27K6C@eKG9Q/<7dCfZ#c54OOL/YNY+_/11E3NR^G
W[QSLGS9=S?6S.S^E:gUC<3=YGWCBQ@SJU[.TW@JD14Q\7L)+;_ZCS[&AE1HH)eV
+PFL?1&4M4F<[fd_dO@>>/X35d=Rb[4]MZ8B5H/FQDa@8Y?X<&1d9&b];d5B/dQN
adP.g+WC,ZT3@e/+]WYBU]cI<+@_B)EA52YeO8bL0)HVdRJ@?-fN8c@.SO4b_,(U
b@#,@>@QN3YRO)[NO:Y)d&HY3d9-d/>ffS1f2W9QYb6P.D\,UN@B3R/Vd73JD>U3
A,H:S\AP&D.ge[8eI494_433?S:)]=P(cg)2]]+IP+HG_;9@f_]YZGG1f31.,C>>
JcabAH(#V9:cW>b5Sc=^,e[X?KVZ+e_9_[LUVEMFSZ<)_aN2M)K60Mf<e8a4/6@R
@=7FD9a>C)-M7Z-f2ZFS7.CaW92eC>.@,]5M(6a2CBfS91C5HG\#^gC374^a.DdW
U;_5,64Gf,DbZGe?[f>H+)fH_L:)&[_:9_H4NAM?UB;ScX\d-9M-0A]c<[V/>Y_8
_<DMO.Y=-F)J-X64d1J\YY_W>;_>PBZMW1J56@EQ>\A0fdYK4(]GS2OG6ORQCaBa
=[ZCWNNFWS68G+XE&@(VW+PM>R1>SF@fd5FFgfPL^-d[@CZUHcfZ^CcB(&9X4_b7
AKJd-T[5\LO&][&ES@@HR/O]gbVZaIGVO2,H>^M@HZ3]F,O@g50E[N1^GY;9>fd[
IH>H+VEB.W-.X@@ffSNU;]/KQ:aZ8^g8KU,MOUKH?2d-?N&-F/<<Y?0WT/;N1B^]
0@I>G1?J]UPJ/IFFg[R/\;]]VNU(_^<U2PVUS5Ne+9(+d.,>>S7FX&C()^+Y_S&d
@><(7>=.HHNC45c@7EUO,cfPR8>RPP/>]TeTGUQPHD(R.bM7Y99RFE3/,CEa9_WZ
1HZ:\9V/H#@,fRBDCXO<=,c.ZgC,/B_;+HI,QYgGcGF5+#Tc:3(:OAd6T)RHM;e<
b;eN8#G4W&3cB&MQNL.Z\,c+B^MDSCeK74GNXRR<A0I77Y:B5a+<(Q]DD[[]5<K\
+KF[D@(JN7OH&_e]?)II+MKXDHf65JPa-EbfIJEd#aLVUWegc_/d4.V_2aIIT436
[0./^Q=f_R#<GRO8#I)IdV:MgC8CZN]>fLJ;b3:ID&DGNbU@W\Q(_TD9RVKA5LP6
?bcGC49dKAQcb\Tg[^XbR1HQ6FO=S^9_<:De:&E#35V3Hb_c#fRf@U6FFH3W5,YS
cQbSDKK8&1;&Cd<KS6_;O=;/&>1,@f#V3+b..ZN#I>aS]U,ZC8Eb4L+Q?_M69L-)
>X=XU^_D8.C7[S^N07^@E\=5C&CU\FV=g9GaYAdfZA9,S)A6&BNd#-P;[TL5SN4<
FNbB@3P(I3Y=0?bd2.d917?gM_Y3d4<X;B-Xa#A=aL6Z[[&c@38(2@WOSK1@QQ;4
0^0C(@^Zc4+4N5.a(;H&;ZF=MWfRX&Y0.<aN8fU/L&gG^J1Sc]D[8D3)Vb#:/PHU
/f2@Gf1Rb27R>H8&O>VQ/b5IIOf[<]_77#gcCP^S;UZ0S4TB7T14&0ZZ:gO0W0Jb
[BeN,\;7WYWO8C&RIH\=g;Z8OID),XaZ)BZc(=+#CSH;^>6J<8Uge98\/QXg#ZWC
aJ;-\>#D[6&cRc?&Ld)WG)VUHART>YC8-L7Y)Lbc\#MPMQf77KFVJgZ0/[Md,5\B
^AfKfH6W-0)a>eQ^@7R9,9aIaZK(gI0050+D.dC^?\C]G->E37C?W)0g&(E3T)3_
]S9;<B6++X7@?bJ^(9O^HB\GAdZV6BY+>4B/PT_>0#Z5V;LTN2U;;:(6]<cT)O3d
J<GRAZ.\E-_),,U4UPV@U@c:DP(UYI>d<]F;28R#47:SZY#R.GZ[LQ9P-[8T2LdG
CYG;#IT>YYZ:B>O(AA5))U[TC3VTI@7NLM=be0LHN/JR)EL#&/NK-?^X0EATRAW6
K)UbD6NFT4RQg>Le.fD&V<BF>O#c_BHg2&XZ/?D]f1_d6YHMMHS7CAYB0[7)[+1,
@1H;OPV^SRDa)-WPP-P#CKQe0T/^b^-L=9W.&(aM0Td-&E2cS:]#Z;X@#-bP8a9D
b37#ESdZ7J.fWX:(/?XTf@7R2ZWND&NbP2\eJ]gH:,<A)ZSYGaMG52d[@Tg_I8RQ
-0+=;O)2fKBE],<_>ZEBHSE&3g<bQbWV7cJed8S(EOHB16A\>f5[+&@W)8@=HMER
1\Ad?\OD)FN&a:ZMTIH6&,\@5S9C]KLL:B2X4?&1eBH);44#KT0fB-d98]88Y][E
:]#,>fM0+.6;3Q(a\:3N<<c_()W:cF-&Z^fVRaS.X@G8(BaO4M)K.V:[<.Rb.F^Q
ZZdHP\_:fSeK_8C^ZW@=1G8U\1eMZ/3\8M&b#M^E.S]<+L]896Q1fR/HFN@2bUgG
32f2/CIPR)C(YBR#.SAR+]C;=OB\=I,5(<J<LW9fQ_d;I=7WTP]NE.&fMPH.,)HA
15@#1I+>,aNIICJ>(,ZJ3,.:PFC;[/JW;BCX3bg>P(2>P5O0LWT/d?cL&ggDS8>5
VW9CWFbB-ba7/&NUb#S@^gCDLec6Y&a5G3<J8eK#ENf0N2f3b]C#GD77G3ZCc/@O
KF)V_.CG>P?W().S5baZAD-cVUF0V^>A:;g[E+51f4-),0KdY:aQRZ1Q9G0KB\,H
KbLC#Y&L3R/9H=;[17E@W]GFbG/?c690dCgb5?&E\0KC&G=bF-23E?a7^?M;QdCE
^8g33KQ3[P#[S&@FIM?#?bfJdcaXYBY:&__9178::>b7?F;N4YIa8fYQXI?R0MMR
>:>8W4\/A]N<#7fJB(7c(KMRWA)._<KTQ+-+.K-M>5?U=:ddA-[)IY#GOR1LWN0<
M#P?5g<a)RO4/Da+LdQ;T=J22-b/I,SDK>\2geL]+P[U55ZgbR+#LX?U0B/.KR=_
]YOEF/8NQQ5^aD@1Gd30))_\C0Y.C@3JOf??[ADQcRY>VOZd??b-WWD2]AD9O,/H
VdBgd;aZbb)U8D\@2;)K^0SEcJ=dGZJ8-@BaaRTNB)=5\4b/NVfRdEd5GgCbSa_T
I_HU#GWM,=T;EaP7.#g85eU\D;T8?5a6J=:E+CX)8@D&7.eaG[75b@VV?_Xeg]EL
EOFQC?/P4(]L;;XE+XOCMR\T1--]<1,Nf5/5>(.J0;4MFe=V7W(d]&V:_7E+G(e;
2#/2&G&E;-V?LXO@[\KK4HcDZ/8;6^IR-/d[JBDQ?)f;gRb^]K-B3ZZ0).1aUJMA
9Ced9XabCRY^]aEcLWJTNMTa@L_U:(D+MAA^#S&V&KgX)^gdIW=.5C@@W+BT1];O
SJ]R/]gKOIfa)Lc7@I_DAY6g.492[F&A5Ba,7&[AA=Rd1a+O?L^9_UA90L9b0R5F
VeQGdcU.=4SM-RM>V]<Q#05+U.L<YFKc7(N_/DV^(+L.6FXIGL(F)I&HL3+K;,^a
e&;I^@D0;+<U<\CNY5=9M,(P^PDR6>KO+I9H;46SL6[WM/7,@O@A99A3CABCR[L1
bg3A<bITF/S[QK932:U0H^_0,R<G=7Ac?GZ82CfVSN8S+HF44^6EVbBQUJLZ.+=<
[\T)dS.^@Q=1=L7F&O5P^-)-+f^:]8(EK(ddP?7JK_,-cQ&;@7+[L-SY;W>LP,6>
XA)?M>>JT/eZMgKO5I(g/7,5RBD5b52B;Q@_Y^aOeM=4?W9J44_5ff.H.LU8H9YD
1IYCP&Z)fNY05/YI0N,,#Y&C]&P+V]<Y_Q5NOW#JeY6^Lc.;TdR043^)+5R.Wf=U
-[H(bXJDY_cagT=&d#@YJ<9-UNME7^:<U=-_1ZgUH4f4]b7^QA]VI&O)JTReCB/f
FgEf;>GZ49Y+S>FV_DE6/ME@=Kd)2Ea(c-/#^ZF2L)YFTUeV(LHL@RV28H>fEFED
3\6A2U,BHB5NSJF14JLO&4DRQeU>c\0#b=bOLJ,,5M6]&KLK?HB/^LEDI^aP@=LP
D<TW@<e6=Q4LFE&L-D:3&TcbI=;6L>X3f^.LQaHRAK/:HDc(66-P5ZT#/:=N/0PC
&Ka>aO0L&3LW[#VSB&BCS>8W7L.eMWYNZ>UdHfM=1.Qf#ZNP_@4fLPT1c;+SV#FA
Sc+BBG^J>DW9WF@ICU)^_,(Gg-D;(CdV>I#+\a4;:N3?J5NO0D.&VaQbd2)fV#&C
SWdPEE0IZ6[]VEVFRUFGDR\AcY_21TTVY<8F@e[.[@aZLf0f?HcR62;2TUKgHbN:
Mg.=c<6T2(<)be>UBWO3ZPQQ]4E4CARdBF8e,3(:e037L_Y,QO.RSeO,=:E&(,18
SB.)#27fT<YJ587V&(DF0D9ZSW;O4USO-?G;(U>.gSP>QY:X;]>.\93L?>eP/&f0
_WgM-VIB4]gS;]6=EIJ9#7U-AV:37;gGaOHa:0</^DLY9ggf7Sf?IP5;f&:T1CU9
WX/ZX4V9T<,IH/6^K:JabBG;.bM[_,NIQ@PcC1JL;f(76[ag\f7Nf]fNCb81f11.
IZFQF&RPC,;Eb07I0GF4&AUP^G4ZDF/N1:4:a\e@:/[d(E++89L11)<\B^;E0gRZ
b(I#^b4AF\@6[;.F>8\EK2W[T]cgfAZSE^4.Af]]U>85a5U^3Z9/CRDA73dNR]S)
f^W_LgeIAQ(-&+1J::5WGCGGBFWM9^\\(4PCD>F8I^T^__I;gIe#KJ4(IXS;GN[H
=EC-4(5\#-X-(;8GKfEBB@LK9OH?&a@GKH(aS6.G1WdH)[W68a<0RAP</:RI;,gR
1OU8QJKSIQ3KKMgU?Y.Z,G#f]@2;P4FD)-)fc\8\b1/H3X5,KeLaeg112B@MZJ&M
AE&.H9C52]F5[8ePI^RMG#AK&9_@@A/E5WX8.6N>BZ#e(F_fW=ONQV9OMQ\K9G01
JK1E,eaW/)8X1HFGXg1FDL+ZP]?Ug6\7WQLJ[I@RUKU=[ZQ2UGX\aR^B9:c:_UbR
=4-U>JV6WOISRfJNcEg96_OaXXEM.W[3+F9IKNZg)0C>3IdGa>e[0;#=/F;RW_M+
YQGNO_YEJ\R.X3Bb-K;0B@+)2DUHMbad.\4SaLSAGE@ec+ZCbF,V<E[9YX8JY>OX
-e0HP-DWRNR&HD_DH,QLF[@]f:5XPID.:3B8ZA70VJ#).9;ef;<Pa#4E5P(V]/WE
aF=P869\SA=PQ3F]HeFaW70J[05bXZF,NdIbI-^X0K<WHWEa8U#I?,3EOd^f[5B;
#R/eHd;_@e\VWVUDbGZ0T9@.;4R1?H4Y/1Ub](FC&4d8>R=NGD6^H878XdcE0>_A
K=R0B_BTT2Y\/dX]PQ&e+d)0X@F,4LBJXf&B;PU=,91:\(WE@@EWcDZ^LDL^8;-M
Ed1+^Y910e.VHP4Z?HGe9\&bP,^a^/52QAIMD1bIe95_:e6.//9X\SORa\;KN:DS
H2B;S,3=3<D8=-5X:I7Nc:MT#UE0FIf\;c4a=,(8=,_\3@3G88]DI^BR)[.1Q2FN
@BVJ4DUb>-Z\?f7EBK,Z2SN6B[T7;(&08>KD>&#NY7K__Y8X9FIBJe,DPcf4:,7]
-U>\&;?K_;8G<8e#^0R_eP,&95eaR/D=a6_(;F/W983:)(8gR39IGDBD]-+3b)8.
/dI7X/K#T;JDB<AX#Qf9[@,R:@6?9AC&6XeS?9eM?T#:c7911P,dcEI^I-cb5g0f
C?KFM1d6BOMb8LA0GBJ3B-c#\SNA\&S#[;2W(O,Ha&P7UY-a>G]X^LeV0S/4-YP2
=W>IdT2W6/?<62OZX#I3@AE>VFDc0V\+?bGZ\52EJSGcK<G/Cf6G]/M]0Hd+ORZH
fXTWXOS.?1/W_E9)SHPMBg])=f[XDe?Y\M2@9Ia+=[.:9S(&g7=aGA+2=;XQ+g8+
4C<;@V8P^_Tf5^EWT9T0FFM.b-&5+;^A([&^M75eZRKP]>CEO:/XKb@B9;^XdCC.
(R;J4D\H8eI0/1-Ha,&Z>3GGd.AOP<g4?YbH-SKZWZL=N6[gAN)a5XcE>JMb4-7]
]9;;a8GJ-WEgU?0O-JR#cI7F4(T[=8g(cD7H)OR>d,)6T/fXHD4TKA[1GJL<Q(B1
Q&G;,c)>0,bD&MMO6PKT.[&J1He_3-,.LZX4b,Ig=G=;YZ;SSQ-1@B,T29e]M&FF
Pb03(;4H3+KLcad2&KA])(--KE:[7P[,>M]Q/105RfLV)K4XG7C4C_SU24HBR^X/
15\M[J)a_<DX;8KE1N2)<3U&HQX+RLM1UEFXGe8MNJ.5+/6KH2C2HA_F6>V@:U]S
/V?DSMe4cE8XE#+2/2bI=1O1@=8HY\c?<3.bSb_0OH(7?52g01+c4^UHXN@97;::
8=:(eJ?DNBO]D6U5:#YSFBgA;If8<0.APN2ETb#a\NJF?_Z9<MAJ#OKUE7/S,?L?
WQ@J?^TN-)XgH90MGF<5+Z^=(/1QQNQ9dSXP+BU)e#.d8QBbgE>._M--e?EffCZf
H4a+_fd.]_[3cN>@5)/f)#UQ^ZP&CAV]O:<.]WR1e\Z/CeFFN1U4WNUg.<Gg-)1-
FEIN#IA1F8]5P1S7;^IS[=]5RQ\?gP.BF[gES2&-QKVcT<I7^Q,(V)AW8R0#[2#+
+MQ/c3[K=[1-6M><gHMFU9[McI,HA2_]=KLA0D_KK)@Y6=58RG,>dM@2g\@4C(@-
V,L9PP;WB\&9BCJ)Pf85Z&M(f3@fW).AHFYH=Zf3E>UB]^b@BZ4VH-+LR.?>Y&(6
N9EaG(3\Kf(L[YG00Q7@:bIL0Gd)>KJM5Q_3^>^@GVd@]WSC9G0?9P4@D+G\f(SA
PGV^8EVP]D3;^HP,-d2W\Y@:K;Ufd:d:gfdTTg)S#2<KcFV0TT>+NXK02HGALY?d
@^4+PKd,6d-g4@74G^#LdJaC9KO_??8(5VGP_+fHX,H#H0R^5]>XFdK^U<MU[,U+
CcfYf.SX2U7P6eY<DaE=TE>R[@W#?&e(_Y(O?0AIaRPe:CHQMJ#MH#R/>#@\I2ae
R.;fT+]g@PY97P[TSMD,C@06OTKO)..:4WAbGKe8dKU7B62a5-d<&7>Z3d[(02>3
+P6?XM^<E_#OQMN\:aW^0NISN\;gd7VK.HB3R>g:WJ3\==f/eS4^FR.3-U&(1PJY
G+\_<)_Ue5a7M1?g=:>BFLd<E0?QTLK++>^bPYQX^CI#GMG\)U1@49U6YA2+?FH+
9I6R<9XNOM8M1Hg-U<A);.f+?_5Mbg);8H890MRB2eeL@<Y_X=4-V?;/45)PaeEY
>Q=7-.XXHeg\_7B,LU8KIeC&Q19,O)bL)F\/<]gbZAe<gO(31=4TGMG+UGdXMU9X
S)V^.W];6bN8VW,OXP,;^S,ZBT:,Va7a\KZ#GJ/UYd4Cgf-].>V]/fHI;)7:#F,X
fKbKNQ:O04#Y4NYH1cG_fO6cIaVAT[&PJ9Q-f(aN@TM:8aYLM]+7SL,==[97EM^7
PIBM,ITU=MVAQ6/O_T+fWH5=,HTA]/0,I_I<&9cSOA]E;e62cD:&UW\KYW-EA.@=
QfJ&d944BOV9MTIe:9Fc)6N.6AdX4J>Tc2Ja(_N@CY<ZAQ-<>G/+-8a<IE3g58]N
A70/HS,B04ZgeD8bUIF-d]M&2&.9Yf0d?K9+IGNFbfNe8LgU3J(:,N\39:[bYUST
+S;Yc50I:F#<6X.EK9NKRH=(a)6a@&Aa0SGT\JG1]++S<.C35)-=,BW_,.O:;6Y&
7(6[HUZ=U?#2Z2>F@0?O:T6L[La+-gZO-]7BAeN>E@\JSW+/8b/\01/V#7:599FU
2U;(,]I,EaDMW.f124L/9Da.6D10CTJ+/b;a_D/;]NZGQ;b(8L[-JcOBdPcEBB:F
TaaU#K^)E3Y@?__a=5>S[;3#&SLT;SSe5CS\A6+O<446O<cLWALAFf&f>H5#^D&[
-Cbg7VUg0M/NGH?L;YZX>1/(\,.NU7P@^DMS3::D[(0bG2OF\DKa;+]#QX/JF,R6
SM&;5e_5661[F.IR;gTVDeHc.;9e6BB;=5W3d99K05[gTPNVe9GQ(J.4=fDeBOX1
NU4?#:7]f,.;86)>CTbJ47AP_H^\Y=/4L(8EJCTE-()S)G,C;3:-DI?0EB\LR0dJ
;b)F=2?@T?R\EcAKcVJ2PdadI8/+QD/2]+@\Y_P;2[LAaJ,<OMPPcgeD_<<4F5^,
,I]);T9W[e6SdR\eTQJHQL0;_a=0@:VaA1(]1a8+?L_^G/7:aF]fa:d;K2H/<>)\
KbQY),M#0Z>dI;D>;eIK\>f\)I4.af?QK2M2?,GUf@BUJ.fI.dg@T]Jf:^PeB,0=
8WBdIVRgWa4>W#J^4g&e4#4^M-=[20Q#e/:fAQM9EU-S=S?)R5VG&K,VL+WR#=SG
g7#Y[YEMGDY1<d;aR<K/3+fGESS_CU3:MBGG.Yc&I[L+7O7geagOJ1&+#PA6-62M
+>#O@bYOPQ8+;1FFTEFcQB#Z)M8-2edF2I0I97D8A;6T)AVH/^9YG;.EH)gKgJXR
&GQL<bf).SAge;JU0<(#EX8b.#P89ZXb<L3gZN3O=:^8GK2dH=S;=2B^GWa2Hca+
SC2)#MFcCURZX5+@X?KeC67H[UbJA74=O:./Dc2V<FBWMO\Tf\3Y]QH2T?6YY;bL
A(W,^]T?fP<)>Q?NC\3:P7V)a8eDFI2B\#4EaOU?dJ5@?7OW3\<LUK9DKH<f;M/T
)@^&aQV_#ZEQQ7P=O#X7WPTIbT_bf.D/61WEZ;2PT+2FR^3DT4,9TBPM-Y+YdBDH
;68g_^>[S\J4Z\4K#D3Y)F?aZUAOdP)5O5(g-FUT[@G;>SL=?@^#.=-NR;/Y5D34
:Z0_cf=Q9?I404,XJCW1g_P/^-QBXI5,R,(M2aRf8.5Q]?7B.@ADX<Xf--S<=#:-
(2#8-,4aK+45.Qe_TPQL&.V+0A&4dS^1B5[Nc@PRb00T_#-HH6Y=-W<4MT(4(gT9
W\;SM-gU/-H,A.20^Ka)+][\edQ/P>E?J:d8_6cd0#1UaQB][_1gcI042(->f-1-
dM>PgQ&QH@?,E;AN=?b+f_ZR5ae)+PaX:.BHMeM1?Dd7F7dV[+\N[D[PFcN0R9gQ
]f/fL=R^9gNJ]=e<L_aU7XcUf/8c-eIfebBCdJ(aNS9M1a-1a/,@FL+M9.BMNP9[
;13Le]PK]B\8D:6#SE5V]?TDH:7N=.(8:ed^?10eCU;E<R;H8?C4VgaNSAW43U&+
YPP1<&M+.1Fb\QR.6&A@d3+f[aR;RRaX9d]_8/=2H<Z,B6cbIU)YbgW6@W#VG.)\
G?HB@5TRVX&?PES+QIC_=\3-\T7L(L[?Y0.(+QV0(=EDWX_.V9eYBg#L:,DPVe4O
5@<DF9dXSJY5^VDW@1HT\9]H(2Y.9LHD5bcX9YME2-?_T.6QS[=CK#2ZN,Y.S)a<
C@MQ(F.UR&2:9ZQ/T@E;B1>Dg)LCd_#CgT<9ED)?:)+=IJ7N,O=S.K7)ab+V0-YY
_afE8.R6Z4E4,5g@Sd>AT?D?g9^28D:NT0=UKZ:J7)G4+1Yb9Va0D5]U@:#Q/_8,
.,H__N4E@Y,=S\IS+@K@3X],)7KG2LQcB?3+U:?YJT-f5OS:[W&0Fe1F^#:6SSdB
59>>08cXggT<8BeO;?fQ+^&NF-eUYNRP:>E\LX\-aB:[2.#f,2]gU<ET8/,D3[;S
S#RU5>38/D926>4_BE@9.c55PAbf>+:B<(O,X&g0B&:cYeV3)eNXGRU(#<LT<g=M
,XDMD0#T6Ee4b-P^KN:OOQ^UB>)3P(ggH8&Mf_]1((7#+I=IcY<<F8]da+>/\.:f
_EX]3D34PI1G1L&Y@9E0=T4[TZ:4OAff^a[,f4QZ>3B(=V2DMDbA&&U]<-f._=C5
0W\N-;)C[34CIKG\18c7?a1I/LG@KSA)5=f(^DDHS_.FB#G(;6YE+eB1KB\)UC5S
VQ+<([Y29[M0a(8P4dB+GASWT=LL6ZW8S2J2@SZDJUT87286MW[9EJ&PX8e)/P1.
I-3d0fZ/]A2e2FX7B-Q:g1fI<=)IB\M=.(>S1b@F<Ag;c1Q/6a]:ISQ,(RQVQ41c
OZ\B@ZeTLeQ:>8gadCIcG#HX_CB^NQQ=454.KDQ,U0YU7YgR9)L1bKV+EdF4AXb/
\TY[(4Cf:L2f,ATg.eN<&B.XD,-)d]+D6H,U&QMO64I;)S=eVWUDVR1UC29(7e@2
.YU[-.(-I(;3=BEV[E\f\J&/3MWE,?dcM_.^I56+d#5;NeTJKR8CQRJ6B30FFE(R
8FDIQ/&&UH=P8bT5X#J(YLaBOMR8G73<Q,S=P9=NGbK&C5EPNVf,)Y76C->PQL0G
M7<O-fT)0=C@O,R6#VILX=CU42ZaeGQ\01I,b1FfGFOJb-Z<L;EfR/C&@6__1?IQ
PEP\_I2X=GG,gfE<32R6f\_BTI\2-3JF=_H):>1E(g2+]<+D1E0<S,QB8AcdEK:W
3TLVS\\ceff740fDW>c4LXV?K4:,FOVWCU1)GT]b&Q._29&ZZF6-R.DK(&)_AcM_
JZ\UCH-VA/#/-,F>;70>WIW8URaZ<U+5/A]RTC0FdCb:1OBN.Sf6511R#_.25L=M
@Y0bVEMS\VBAC/?-U[aM[]V&:Z:b78H<.LR+gJe=RC\g&YDJ0.)aD\0f-=e/JYE,
2ReRBB_&P>P:=-QDM_<_YL8==GU4#=5KC[ee<fMAUWN//:5>d#B&HS>K;Vf2<gCb
c)0KGSeJP6K<#&0@[eB3:c1>RHZ<2O573<4S(]g87g-dN_<KOJU>Nf9E6>2a/<3+
_Wf:Tg.afTMDIIG)\^/E7a\ICH9L4aL4G^MS,IJ+0F,\1_.5?GKL>@244W/4^,I4
F:f2Q&3^(O[QXe7_28;g,)cX=R]NH3)\B^Na^GZUDJOeYJF4&8X8U?\8_f(4-PSE
e;1ZSZ>M3KENPHUBB<^8g8S(e)\IV8#YY@D;1@N&^G^XTQ=LT:8?W<a&UP=S=0?(
(F;RTC+G(CF=7AI<CN<]VSO;adF-;P:A[Eca/d^a0MCIA8Nb9GHGN1>]C&#KI0@6
D?;HVI-D^5G2F?C-FCZ_,>_(2MDRRRb@fQ?e6._4B&eAT.<8018,>(MEF<1ZdBRa
:MCIW,DUR1U(YQ:\D/8?QD+A:H8.Q#>G:^-V:0eE7YKG<^#2D<-Cf(N_-KaCOd9\
U1+AQg)Y<<aOB3?-P8\]3/].?(15HgBa;P^B<@V)fAX3ZU5M).VHD+]OUEDC0-Q;
R1a)QP=H^)GOZ-]JQ>8,F\1bA2S:U.3ZE))EVH_f16_5H1d&WPB2(0)SY6@](4M5
=UQ1C?0]6LI+bQJ2.TKMdLF=4bT5N]O52Q=EML[,C#9aJ8UJGR04B_:\KaJ1X@YN
&J@OP)MD4(g##[U#7?I]TO/)-WP,Kg8B/)Pg\/QFQ41=WE\6M[g=Gg66BTa62#aL
D:7;+cHG/:.<<DZ@>@cG<:,23_-N;09Od;bX&Xg7CMBR6C^6(,<887Y[AN@69a2,
g^.?LZM_C&&R_&VG-Q-U_U10>Lg@J56XJND418MX325M1-5,b-,ZEcCL8&.WI?UU
C1[6WN1K1,FJB/V#f\^baIU->L=NC-,)+4JG#32eF4JVbW19:2M^DRMT2dP_;W^J
A;cOLZ7]/7&7>Q@_36#B_JV;&-g?)AfJ^5H7Z7&c_\08?.4BROYA4#0-Y:fc5dN?
/849)gZG1Y&[\Q?5<9fK?[1-=5]MMT1>ZA8\]CZTM(SL9_aa\]GFe.?L[D+@I;BY
6b-.V)I@Id?U,3+f/QF^)<a])De:4<KP_fT.M574c#V<>a3_?VX4e/ZSX(PcOP=.
H-T73<(d28IH?&N=/H/L_HfALO^J\]3S/GT3>@9.a;d_.(^#gGF;\;Z8O8TG)]=:
LX6&E1J]DCNSW@.Q,Z)KR0S.N1PCEMd).\;f[[V_68K5A,7IJR(^7.>HK^XaLe;/
91d@T)]FBJJb72QR8R;0G_ZBfDJ)c=E8<g/1:PP>X:8#5^-NAXR^gTVJ.CX=GG4E
)E4+(D(BO5dVJg_\,FF.H[4/#S5)SXeI1L[7RDKa))G^+eW)H.YL(GJ(2LO.,M>V
OT20gOK0Y3.I(JYe95I3EHDPMf>^-Z,_4.?>-P,Y3[]06TcYV7Z(_&\(XWWY9>?&
bLP;:P_HIJ\K2=7=3RebA2fZM2VJHccRI[9EfXJ2GZH-IX\7UA<3&5.P:]KdTe5C
eDKT0#1T@:_SR:GdPa/)/=];eC?3D8E\bVX.KJ>9Fff^,DKEff,T<^Q6L3b-^&<^
[GZ[0gTCB1MD;).87Y&</fH:gc)E_g&LZK5/C.?/-02TC&Y(T[0+8ST>^#3cP=R3
31=_5g2IJEFB<.]<3PD9#dU)367eC[Z56aBN^Y(Q3>DgAW,>ZUcTYEM]S2:B@1QK
_5]EK3d(RVLI+-0fH+MA>;W?72BXMJ=\ge\cB=#K3HS-Q?UDX[;dK&1XV/[WU2V?
\?3.[U4X][GSDE:&]^U1]]_Z:@cD(/N@\UOYba1&8&<0e/V&?,SaD=8.XcXUNaMV
KLO=bB(gaWR@J2(VA/cT<>=TP-U0V4RQYZ2)==gP8PVT=)EM0>4,dN1<#;4S73>1
>&UXEb,1.2&QS.QVQ0cL04XUWL#3cadgKHCaJ[NX<Pc1#4JFNY).4b->N)1B=/PH
91gJU;-F[01Y</(2.dRTJbJMACF+C]b9+(3,N0)0bfQT:eA\E]8[H7D#=08UGCAP
B9LH4RDYb.,U-b@(6)T5[KZ5e<C;afd^:dGEf^=+1P0I@[,5@GK=64A//X.RW>C&
K(e.>g&[\IX[LQ.NHMPB3HM&;+O?9/O8+GQA],\WQ.2/]\KL.2;&XRbV.=e3aTg[
@d\SJT4Y_a8UQPcZRVSMg,aHX[3T(0?.IXX#4O]^gAPG=ccZZOHU8X]Wd+g=Y@ef
=^NOeR1()aRYQL,EbUK^g(74F<POdZHXX:eL7Lf/46#YLS;]EJgOOZ;d4MQL<PXH
8<5O_B0gf76XKBTW#XLa@\&\ECEFU#aI5LC5B;>5[4f@K6>UMR@2X)RM(#0@V=Yc
Q@>1Ab_P[?>#]G79G\HO0801>OEaSd@Kf&/ZfcE.Vf>NA3Cg/L?C[UgJ_D7K.?.d
/+HWCga&;7FC\#(\Z2QgMC0D3e_U6[T_ZH(&.[bc4a_U6/;R>:4L)]7QMO;\_=>[
685c[N:@4,)Y&MUAdd1:H3KPXWbG/358g>\U99W2RI89>CGJ6-3.DJ>(0)_VgUU9
2AOe<RZ78R\+I,\BADA[c;=,^g_8/\=:N:OQ[P0OZI2ADW^(c-f,YIJ7HW^[QQ@X
99b16eP8F?1S[TV3aA0J]);-0?GG&49=?O]cJO[IWC0Gb45/e7424(DZ.7f7K9Yb
1H5@e&DFA&</LUYXV&d/BOTP:EK^4ZOQ8e+?(QH+L.,KPE:-54^0)A-;aBLVPQ59
F5AA1S(UG4OJa,1ZdbR4(e<XU_+-E;:D^gDI[N2@25-;ML[MMfLQW<7R3X.CK18O
09\a;Of/UH/E::GHT@e^=YBTE7Y(23S]Z:DPgMBQ5/@C#ePAP?;3T9Q-gBWB2>ID
#Ug1,bcAV4,Q]#SFLFN@XJ8b>c^:A1:^19/=N;90>N:N(Z.cQcW#P8UMV]b)5cM2
EZ:Q1OOAZ;(&A#4T7KDM.PW?N7_8caeCWeYE05)2</IGA/\Zc4G4_.[Tc61=.0Oe
2RV?@,V>-A-g08b98KJ#MK@(WQa(b(4OTd3+Xf8&H>HXIIE45//R>U<DT//caY1E
9c&(8V2fB7Z,\d#]B(#7K[0P=W0(.(dRGa]/QGcH1QC+ZFGZY6QB(/2P@GX8ASKc
K<D(G3E:6#eDbWf6BeS>((F#EN4-32-_&X\QRX-DcVHEAW.J5B]F/GAeQX&::9_B
:0-<O7KW^K\Ic-d8?IOT5QYN#^Q-=[+a(g2PVV1Y.>^HE+>4DP#J]cgH_:6KVWb4
b(2?[2SAQbc.>Wd#e(2<D]W&4ZC]X2Y0ETA:=dO8B70?fA+faa>2@-=PIWKYf>2P
Wa5Tcb-4IH-/_@>58OgE2;.N=7:4?=\U76/0PZS7KTA:D+3V#QGd1W>;L-JY6^bR
+&J=Ma@4S>WfD1?4>?[8]DOIY<4DVRcJMfU3#^)H;X-H0P:LPIR+Wcc)bfHL250Y
5#eUY0OX+IIEBgC+,33QOA1fIf7e[B;?3OFPL,d>J1X>>^,+)Y7O&O]GB&Rb0Pdc
B@E80WM(&[6cI-,)L0\OCgRAKU>M[M7:F(aUO7Fa5bQ#CP(A3?Q/T#0M8)g9>>Ef
AXPJCG=(W,WU5IF;+b^c@a[;@2+TTT,0_b@M18YLCU<3>W;P]E,_7]b65G[EH&e6
([:.>FVSOHa8D8)38d/B_Q6_A98DO8b73X@LNO=P;eb>[[]:X+d3?Be[E4g\A1_#
c:_M<@-;NCOG_Ac7Ac2&K\XPC3MZUC:ZU5c<9NFD+_<eK_7CCNCgV28SdZbPVO??
e8L^\9VLARZ3UWRX^df.P4LY>?<ROD<LXBZMZ/5<)-BGXBS67J4Y;&6f2=)U;>6K
XQcM+C1BBS,?->(We64#.EdDZ]c+EaI[_6;2RW>aZY?gU\SUe#\?K&0O/XQ@dVbG
R&0:A@G^91+6g]Fd+8e5[H0[QKgO,TNJND0@5f;(FfcPE#I2b,>=b?W9U^fK.>dO
&3LWA[HVNXW=d;eJCLdDgIXRNC&Y2@7P4@?e)G>b1&+QM^2]>>W\OBX2[7G0fa^)
dD,YM>c:4F\>J_EHf,)TO1001=9?eNSCDH#V<IX?/2S>1QMaTF8.<c/fVV:V_\2B
4HZV6HX[a,<DVV?dR-O^[XG>G]]05UZ5cPI3+0cgASgNR#>2K5^V;L32WD4UQKIY
H4?PB5POZMWEZ-664,U=.d65[(O7&CS39A<]YA_7ZYYE]B2TQGK>VT_7;@ZG#+#J
5g?#Rd)VSGfdTR]I0IG__]Ne6:CV@GBPPR7Xf@OB/EG?:gdL?gK,c>2ZB2(WI]@e
b&(D5M6?K;\S2+eTX3HadSU9f@24dD;I](AY10WSdaWNP4d\1bH)A_87;fV(),28
(1U,3G?6_Z7^WGW9.^-^gG0?A,0TGW++9+@KL(,]/a]&O=I]b?B=,f]@.HW9V,0^
Y#W?cKD+_J>@.7KIK]14bPISZafe0S3PKg1B6QH:Y<^a3?IXPY.a4LV9aI]2W5R&
9B1)Y2\Od@TK4XW5F>Qce))Ae+ZL);?D-;W0R?e[4dV&^N<>3,N<Vg-;D5=-OYZN
0E(][9+CD97PI3J8++0I8/>#(^8H?UZ3LAU/>eI]/=PG+A=J,@XTCd]QJCaY6e=b
3Z/3MPV,a(#&BJfLO-XbL;UV[?dV?:?..1T<&&H4L+7aa-MGIPH&0bD6_/QA6d+N
:=01BbO0Te)J/P13c>1.;9R]aRE,WDK@L\SeBR&F2/5K)[H#ZMB?/@:951B=.U<D
]>c6R:T6BH<[AF8P.Y]9<.:V].266\V>g.;-C\_W+(V,bOC4@aEBG1QGH+;\.T4\
d]4LP9):U+:31I_JR8+RTDB5PEdSgO4UPL0\=?11=DEM-D1Y_OS(X&Z3]9EbcTVI
T+G[GPgU>4HPFSVZ,g<17R@]P][=4A_:f@I#.HVKe/;6T8HKBBcS?SU;Z+D[KF)B
9NK8D8.>0TJ_QZT=?_QSZ4Ig_H1KXN&+<E5QQJ7YIQ;;S=V0/W?F,C3gJ&H]ggc;
7:\81G0+g@G=&BN=dQJ:^I9:f-@T;>9KN:09e,#N1X3G4/eUMK#a>CRKJcg[:Ca/
<BBG)@S>ecNBc^10;T7DFCEad1K_NM2O?aH:P2;S#.1_AF(8_[d?O>DDPb:,?TH3
@BH=,>)MILBY)P4<L9?cZD^9M(#OX\5PH9=\?cKKY7@=/=N1UB44PY5Y[+F1a,)-
TLZDc@WC9cDSL=.R(N-;XARILP;YZg>=Q/E9HTFGCgdIcPO?d?^<RHR8+a^SAK,E
ZZ5H9CI(IJP;HN12(AY3(WUOgD.ID#[aL>P+c-,N5KQIXaYD?a?3<?AU_>Q^<;0:
,\:S-<B>4MM6?Qb/;ZXebG:d)Sef-g=:LdKSe8VcD(K2@MS2gY:/=JG=]+J9R;^Q
^7#Kd;6\@3R/O2+N+>bUTe=OT<3(R5P,A+eV#JTf9MFD@S/LIG^1gJRYAc4[(;L:
LA5+#C&DR/fVI7=bD\V5<24KA.b<]e<@ecdSCdEB+:ZV:4&A2XXJ,4LY3a1QQ8Od
g#)>)[8=0-.HeM3HYL_^]7;7e5/Rd:dD0Acg[91e>Xg\<SAGc/(KH_bf.0)#YQ3\
Z9712;>);576=JBc]T0a@<D?SMW-)/=<aVK/Y4Wc5AeafMA;Z@)gU3L_2D<WE:5D
_g+9?#Qg[7\09Z1QZ9LV2c8fJQgT:_7QVAS:+)c\b[]L/-<-/3BU97X:H-(&NSDZ
3DTN[MD4E_cNfG-\KTLe4HWU1M:B14_gIBCcT:CD#Q<>VNe.SU?D_JZ[Q3:T[Z:5
gPcJ<\(J]2E,AD27d6.KB4=<CLD^4+_eMZZZ(K4BCM1XI^@^-&bU2PD=ZDE4Q@T.
A&2(Rf_\=-.2>Y3ZgHO8D\dDB8bNg0WG4>><=bGQU3YfHg71Z[_EfHPO.L_=c./g
+FR.74G=33JN(7L7863KUQ.:a0G9;ABZ^bZQ.)(?X8K3df_/U.g@K+6C\SUCL>f8
NMK0;GDYZ>LR>V_)_[d,V<6cU@92NdGaI0d]0?Kg4DDcY.A;8,L.IOa]Q:2RYOC+
0b2fQ#>aTdU+,GdSNEB<+D\#4DH<a#H,RC^R]S4?6>XL</,:Y/,Q@H(F4[]<=:H5
f=K;-1V-M8dTF:g2FS,#4(P.@7a)GfV-L\/@gS5VgX^7\I>0B5AQ3UTH([e][HD@
R:Z-D4/c2IL(F&V;=d([@0P;2U/\_(Y7+g=_GP4f64f=YWDH[=MRY&^3S>IQSC0Y
ZE;F@2R5(H_3d0=g(>KeXIR:a&Z9_P:L\Z)5:N\c4ED=T8T6>T+B6E2R<g&J]]0A
OD\Z+VC>W9S_B:?YXfQM.)M0bfe^,I1b1-/2.TaS7O/O?2QL/+6(@)#<L4AY9K(\
#W7]E<[ZT^Xe6I1>)1:<4],2917]4?\CY@\3;_EA/.(>K407;+DAS>79/965M3Ya
\.IW9X=eK_FC,&U>/d#?]:g_P6X-Y#GA^bD.D#UA1d780#NF+9NFR9cWX:aK1347
^IZgV#5S<I74\GL:D\@PR]c\#IG-SM,P-<a>+:9f^@Gd?\@_\^5]3A:)RPW+cc&S
fG3Dc96A#Y+\D-<1]?WRSK\gFd^V:4\U2ZVP0#bG2-79#fWag;C:O,VC_c]c9IVL
)_W1\ZCMV(J+be\]#T#[2.bEGT3P3LZ_UYP3@d]\9N3cNbXJ2\Q1+HSR<Cd>?JCH
6?aH]P-^gc@24?72KZ;&2/VSJ)GPRK.;&GEZ](&<_K;WFK^A38Ec<SHLOE)?a_C:
=K_9<dBd87H@TO-54X]dfd-E?aB+1O3\:X6NIP^-fG6/@T-ZdUa4#fgS2N=JET02
J4+E8??\FY..U8TJe=.^SUMR:_3;WTE7&Q1d4b@J@dF=eN&Z4JU/e)ZAd\QJOfC+
4^9cb3IBK:<(_@M>?(?E<QRc6L66X]Q)1CeUPFDPgSXQI2J;//QPDAW(J6QGT8;,
HgTc:,X[?Y[4<aES3e4BP;4:OD6BDCKE,eO-+]5[dVB0Q0a9eTa-CS-Qc67?G(K>
3D&/U&\-H6bI]Q7DF25b,+9U?Y]:O4A0@\afR@,BN4f8KG?V7&->g>]K:@2/JT.M
CUbBRFaKd^I;^YLS1WF4;[>f5Z?1J_\f8R;_U_dX6UO+8>^?b7&a=Ea?)ROOFMLT
?TP&0f2&bR>V#ACCdSbL/3/@:RXCb8Cc7]?CfQ[/:7>8VRAc#M)2ISJ[8B^GLaAd
,@I.+9c_#KB]+[J=)cZ;-[21\VUXSN(d(S+L-7#,Y=[K4eHa6U-W4f9F<=g1O02,
?^c\J=72?2CR]_LaD8?BDYBcUFH^CP(5&3Wf.cNd:XRS[,bb=RA&f</1P+DAVbEc
PfM40L2UC-JP^0;WQ3#Y;D#_dENT/.@KaV1)/U4<:b<KLBIMZf4e#f5=KKZ(,Q@Y
GR8Pce:CM^abcBV-XZSUB/XCE=3C/=9@;@,0aEE)9AK@Y4+LeERP2<9<FL=3)\UJ
AQ2eV@N2,29R:_/<@C:XB&ccGR_EFVQ++5ERE4RJ]K/2[MUHDQf<CL8Xd8a]B)cW
;:5a,GMG#UeI0L\N5-;K-f]WL.?V<,8XN#(ME;Y2(5P-S2LD&_8&gNK.LB,#:)[6
&_Y.^HO)RDN,VQ1ef?&<71c,dZ9_U(F#O>8BA^^L@D(R@69HT)]DNPa(\N@Z65-6
_BMRc;?0@eKD>KU8A=PaOIYF?RH,Z;VcP&R)O@-EcH)HQXg.?4c;)\bD;8IZW)?;
Z=@M+=1L0YP^Q[Y2U+FT#O/AXEUd-HQJY2\-W@YQJ6+a;HG8e(<3EC-VIV;JOR0<
(U8K:FaX6T5,A\8PC+M:[3EVe@9/3&W=aG@&BeW0P4f+.7I+5251FQBY-G)KMUTH
N<bQE[;DZTLJI;aZ3T]@^fJ<Z=9QCSDF5TNEg/f4g)S#\HL]5X&bXTEIQ=cL5]QQ
W_+dSO:)e2]_GIcMVYZ6BU:Mc^4H,c6IdOB>JRYO]fZ?089=2d?(V8YY;J)]gP?4
Y+1>L-+WEFbIW-]8[/Q-\CC-Fg&7:4&(Z)Q=>MFg-W26NPc[L2gg#2MZ\IPTM+MG
&V8LJ::LA\2ISTFV>9FWEMC-W[Q4R9-D<YLPg=Oe#dMM5R)+Z+=;gf:0HWAUf/7B
0IOMN52Y(6e],^Q(bG&),O-32^a^aPdX]CISDL)G&^-^Dd&e.4@FCPbC<>>PKY-?
(6.5\:(gKCe_bFdad0KYX\HEB]?I+AV,2e@B-d62&g#.Ue(T\KXPD.1e(0#=,C-9
PXd=g5I<R4LFdHP_YPEdM.U_2Q+;;f7+6RT4,2X+/DDRe#87_JGPf57877Z>Z#G_
=D)6L8.@LT1A.=b3M=]<GU2WWgFf^TEEE,6(6JaG;82)0.N)dQ51RC9Q7\U)#WUE
)0FIDe=T?5_/G<#g,OB^45c#Wc(+44N65K5MX4Q523eKa(]BF\[2EZ6@(268O-7=
#3SSaeJK0N@VNM_6GGaIbNTR@&WH57/E^]-/b92TC]deCTcUKD5GAE[RK71CKLIJ
_<.JE0g74@7Ic>#cHR#ARdJdgbN?^JgN5@5YTUYcD3RCHJ:37V4gf,65VEQb5AS[
.P@>-3ZP(>a2RS]@X;F5WE5SB]844/aM\_BbP=V-:@IIZM,/B#0\XdRI:M]^cgL)
eNF50,K@@BH\25g^#SE4U0QY#/@c)@?A)DANC+^]LbFV##<J#GBM9(&)PX.FT:.4
XFa\I78N)(1_P.97e+0CC.3,W)/QM6Vc^ITYeA^D<YRfM<\H1SOg/]\WF-_fODUb
a)e^A;T1Y0(Ld=-g83J;N9WCFc/N-0CD1]TEM,B2R,L#]b>d(E2NUGDff5.b6&@2
52;H94,8aUNL:?T#ca;&e#K+)0IF<S\Q\D(4P?2W;_Q9WY98#WO(&B(@39_\aKG8
K,eXfAJHcL^6]X)@4=RHTVOLO@8+Q])a=>&M1][#I[-@5RdYC#\JG5+RKJ)_1aUN
70W@(13/UT6B,<++C(:\-V1d7TF7/VK4D7?ac&1Pa7O/0WQ[F/fV8aRe(.V<&O>N
2eIUYQ[L[>_8;d--K&YfM.Lb@5ZN@M:aBM&,X9AgY4Z<G.L_)SSN5Bg1BPP)1dLQ
G2PL(H.Zc]NOb7/9=/+[>]OH^0,./K5[)TK(=P&LaE&=9?:;A+N5?=___Gd,[T=M
D&WSPf5@+Z]&&X,?MP(DIRZN3SIF=BNPG17HBJRN)_B(Y4+>_(+JI><L)dVcZZ13
d2^ObGTd/B1IJa(./:#>1&X6_AN#UCD4>7J&f_?g\3WU:?62,0?W98TBfE?A4J45
H<\e4)@5?#6N+aY8bTd-CE([KK(/;Dd7:]5Cb_SGb9?SOZNgG,=NU83\8YGQRRJU
&/0\F6P+<@><56E>ESMY+H^;>R+Ab?O0JUcPM?PAc@VQWH?EK?6^a-LX(?1[[-UH
1^OWLN^WVSQZFa:&=+R5HT3D0_OVR.GLYLSZ,/PEREP?98c(6@@PI^AS5(c+JHMS
bfNL-aM4]fLX56aY7E,E.DZfV>W^_NTZOJMZ:98_Z6;Ze(MF0BHSe[KZSc0NgO=C
0@B=^QdB.9-XZ.dKZF[3[8L&OdOC^XF&)Y04-0;aad(XG>?5.02L3EUR2/F.eYJ/
d)a^5-6U2:cZ?AB4ZG+(\48+XRg97;J<IGD4TL,E+1_M?EaXcgP&&/M8\0V>TGZ]
LI]f4?/64(P?&_6/HgLHOVA-egXFBSSE61+G2Y.?R5/#e@)DHRR6Q,O]_.XH8^FR
CfNT1JNebOJ:gdD)O4c-]Y3NU-TIb)GS\P@d.<AFJT1=,f3\UU9TZ7EY[a[D.H[L
)\DB&IcI8BX@-+a:NM6I5f-#gR8R]5Db_YJfS=O)K5BN2G/S]He3Y)10&5K>EW1N
?\Wd11_cfJ@8gHX+LD0cb;?7Y[KZD8RC7>9IX&C.TV;>[=5BLZ]f.(6CN6T6>B#O
P_eVJ.2J@g:BGX7V\U(bZ)e@)8>ICgW&bEgUU-KEC\CaRUJU9#?fBE;T:7)6Q#2M
.MbROMJ#FFMP7A7@8C/)cgF\VK,)CHRAKTecJ;K.=-He9N,AN##4C(=\Sb7eH=&X
<#&-NgBeeYWe]MOT(QF&Z4AZ:E=:6e^,1/QaUTY<X((AU2B01fG31DMDXMf8N:f+
9d9;a#-/^g4FM8[\Hg[Z9UW)D7BFF[H3;f1:E5aLWO&/;T)><^.9TCQ\\VU<LQZ;
3dP6E/0H9T9Cd9fE)fb-@+TS>),Q_]@H1_3]d3?4&6ZH=@-Y7U+B.(1V2V9Q/WQ6
(^C&g1SMDT(:-+^:S)ZF7;2KK-9L5UAF^:@M=9UE-0-K\D)BXg_Abfd_2N2J]=da
&P:+0-08e;C5MZ?bg>HVA-O2@,@Y1a9\V=1?<0a#Y:O\\PVLI\+?f+<N-G7RUJW0
GV5@JZ?(b)eIcZ:agWN,&JbfS;(QG3A__P:Y[WfVDd1QV(Z11G(0UcCNW=]J-dX?
T#cWY[3+P]DCPYFVBW.dNJT,M:g]ZJ?>>=\YYC:\V-HaSI(,g-YB6M1f9/ZM,(d1
,R5P1+:Db(4FJU4R2dNA+F8IB0<R=78LIE]J7>@BCS8ABcF+Q1H#]RI]g:19,]^G
V^3<,e3,=VZeU.(Eb^aZH5MT1KT_6MDB)MF=.OJUbGb[OX,;6LJP6/^A-,XadFSE
.]F4W63<-LLKF86JLD)dXDMC&?FYX:>U-(-V:R+7M,8[cSd=-[.M[&.,X-cKB(6c
<\:_VA5FEP<3Pc28R_69:[d5H+fKZbHbL4&85],a_cG2.#PFT]W;4f:3.K]D9g2V
I6aZRbUf2+b-U&bJ4Y0-J<aS6A<0[<CMRYD2d=@WD96/f_)0=6L-XRC?I2A-X>M+
K-#L(KDSf^^.f++e_0?098.bR?.g&88Wc_F5=>:&I64SB&SF-8R1aN[Q(H_cgXOU
I)@1I41H/FC#+PR.]+#4WV0P_O/dWTRMPfUZREY4BO2K]5Xb,8@P=eOU\.-1X;?I
CLQf\(2IaG/AY.gTOcVJN^K0SQ=[>?Bc8:35ALBL]:BA#B90EY+2.+ce5.dDRf\J
6:^^8@eOdTc>dCI&2/S-?@8B2^&SS07-Z?c-cTDU:d+#9.b2a4YgO/GW<,-[<bQ:
ZYP?GZ+/K#ZXf])R)V]J9Z@^gV&3J@KZGF&ZBa8<fB-c9HC;&^P6PK[DdA29SX5,
=9=g5)Gc)I-+?_gPRZO69c62?N7T#J@^0OM<R/B&/(1O2;EKaFF#d1K24>:+gSd4
Rc+:d7V+SL=[9ZT+)09(b&FeKBH9UF>NBa)g[Z-L1J7TWe3NKE7CLU^)L/YFQ[F>
]7SXUOdD#U9B>_.;;:?-g>&BX6dPQF>7Kg]7W=H=0<08=IEIQ/W,#C3<LF/2#4AB
Yc^fB8RM^G8BI#beB&R50I22aP4R4#:_-.^R/^/eDU>)B2Z3&PM+V:H(S(4eHHg2
UdU1&7@CD/a^gV@NEBdbaZ^7:a2.OgGVdD?S5b5#fI(9V,\47A-eM&/+D+VX<_U7
0Sc0&Z8O/7U)R.306R(GQ)X#fRGPg8^f3CK:e=JL,,V/RTSV_PQ])KQ=]L(<9T#\
X/1Q.@:QFa[\ag+),PT;P2+=@ee5JGVNO90>K0Hdf]EQSMd@)30W]CS>YUP2)[C=
4#PDdZRY;_UO_\)[_I+SHI],<H@NZOfP<I;XW-c2eZEJVg8)2_+\SXGOU:1+5XSA
W)9W6A0DX_c4VXZ+7(\6)c6F.QA\:75?-:;FYG:]Z#MU>.\cXWd]dVE9INc/2H2^
4HJd-7AWZ:&-(Q5[V5TTMI:SA7GAQ_M+C=JY5M4/38[94?VGXMAMMDB-#WM)aO:W
2OCU0RUPOO4@,:TG&;,7?b4?2aP[<K9<SW(M]^G>5-BW6EVK:=C4@W:T6DD.K\AR
X(U+E11T?I60Laf+98f_]Bd^2[c<2-gXU6dTG<NQ6gIU0.UJD54d=4TO#&Y,&V+W
_(7HgDRU@g&O#d=H>WHN7>.WD7e.VJ)B<;9-WX.Q:FZ_UW&V(fJbd/2@)&)[0<fP
+V@aH;?f=YO#V#Ze&0b6E\T)N97gP&+,0PLPA3__Q#+<XLdW.(A6egKZ2LU?U9/-
(B_)W@5II/3QKJ#&>,;G^2D-O\UJcI69ZaG[#S0CbAPc,S+(.YL7B&(^d4&W9POI
W;5X34OVV@CbK706dV6Z84&#\,OV\a5Og^US:VFf[B-g8a-A3P)37H8<S.fY)6/<
X6/+0Z(eWL&Fd^gE:GD6EMTD<bCBLBP,E][aP?DR4B.8&.TKF?LUH=cG\d-M.A)d
b<MeZ?4(4bR4C=d3V2)H/be,d<@>S)Z.=+f?Q,cg31N]AOWaH)c@P53<4.D8Y/T(
SbPF]fW7^1O@EdHUA&D6,SNOeTK/[6@Oc&D#g+e2O^J1,G_bZ:WAONX-\>EOH-8(
;D425b6[79.OF(,,a13ff;P(C/^40Z[L_Q,dZg5f+]#/ZdDMAZYA(D&I8ED&CG6Q
&8S.=\gPaZLGF/285dVRDBIQP5JQ4-;K_4O=[73>ME4L3@=Qf4-Jc):ZT9\J&,f0
PLX6<)1L0B-U\K&MaDb(cQ(f.^I;DeWUW1/fK-&8ab<dI5_fP^@<&H6+EDKgd:ba
<VVc:I>0T^5c8a.\CP<6C5C@a)b8];0C6Q8ggQf/R<5Y:JVPXCD:b);()fBD>6_(
C-g;/\,JcMcWP/0cXSScg0dgCLBI;4gd^dV]>J(d6J5dgH;#J4<57FIbbB;+A&+6
.]CR87JHTIN((2D87R5RNL=EdDd7_J7Wa+eG:/3=+Je7(Pc);UG,>^/g9a1b#+>:
74+DJ@9S(dS1bYRR8=QJ[V#C8Xe[-[?Y+0DGS7D^d1>:e.7Ad1&@ST&IK\A_O;4J
?<.>H.=@&#;+5P\@J@K3b/O?ODYXXf2,60=9YI=;FG6#1(I:ffEUOL(R<7/^0RT2
:K2bXfg0;^AM=P_&YZ<YE&ZV.11IP,3I@?HIBgZ/LL<#].K7U-?O)?T4ZFbMVY04
Sa[d8@d8U&,<,Pc2:EA6eTDX?H_O.))(16ICS40f@QDc1HOR0cb[EJ^[UT4FC5ab
fHKN1X+M,Tc;8FU6>P\FD1F\=Y:9H2dF?YTX?+-YAAc<S-H;#JQ=;VY5WJ6OFJBG
gJ\.dFT_:=9<.eO@B@&JA_511_028059:(3fLgKN2<dJf1WG(8be3T:>LbLM6[^M
WUOUS=T#gOB0bX7&Nfg6X-AES:AQa#/4[)VbODUd<IQ,:G6+6J\[9<Ha;;H\RW[@
VT<POb0?RHce.O,[S_P191.>>^<4()(CM@3MQg\7^L8DJ]O.KBCP)PS/aa+1O8W^
a3?bN0FDW[O\/U@=aPWd:IbVW>HGXaSXTC?d]]J,EYE:g-&CHBPR.;IB0BY]C_1f
,3R<6)]1DY<Z<UWPATEAE1:30U?5//&#<45\J?aIR1I,::8Q7;+A-VOOKSE)UK-]
Y6d@#\W]Y?3/0VSMP654+QMbA#?I?+Xb>U]H3-G4><SRH.\AQQX)b5LD<4/R0GOT
6H27/g:I@X7TT4;d@PHg<@IAT9V4RUQ=Je1]dF=<N\fE2&Y#O:@[QDXVR.U\\&:J
D9Q<P?R,b;5[&]DR@74f+=f4.^NH45(=Yc3bG>g(9=fa3^GGJ=D6f&Z?&7C8-eBI
+TFM^0\Q/fNT^B)?RXE;?MRS(g:?a;2VDUd-eY<M<21TdfYcQQSI[\3&C0+/;+Re
fcN(-I#@)O@[U/1<E8I7M(/A&3V+fK6JST=(JdN_U6eY8MB3c2RO2LH0TTLNXY9B
Z0\\ScU7KSG3BE.4JBScCW5U,B>XK5-:U6HKa7g39ZZU/HBFG0WF<:0LLVJX)Ra;
CZ87J8K5;=Jd7f&8=f\X^7+O17c79H]O07S?a00D9)YJF:4&YIWSV6G@63\b7fMB
PXDbeR?;0O7NaP<Q.F4g]d9BA6CQ=&F&QV4VCII:;\8,[,O(e;\96Z2AI.JLEL8A
.L/8354+gA-R=eLO@ON#C8-HBR10[>W9fW(bTF7A69-21?d9(Wf8G_^_.:?@N6/>
@e1T)F4bS-;&gRK/=LLAABJ=JQZX^5V[7362-E&-HX;aLC;\#A0C<\)#dJL7-WdN
?2BCS]6ReE5SJ;>f1<c4c>4)Ca_;(](9IJd_YBM<2.74=V7,5LP=U:>HDdV#SFR2
:QKC82MVV<eI5:_]]W2_cdaA1?^g1D0[N&Ka@K]RRQ.:-fGGJa4,7[8(eS2fTRMH
XKg:6Ma72HF=B7L?/JeU,6UgE0-=)Uag&[A5/^KZ&4.AMa4CJQQ/fHFY/gZ;<HO@
I(a=OUGdU8aC6OW[8SQd+)EBJb]V:S\14bE4JEdAQ^;(TH<PL072bN<Y^U3?-M3d
M_VZPNg\WE[Lc-E:S1TceN?X1b.AMWT0IagIW,fcSYfD6X+_Q7\DO81\VV1W)Hb;
RdaV9b@<X&K[Y:g7FT4&S?e8MHD02NZg-#b[IL;eI9gW7?d?HQ(L+[0a)_Dc>_cf
XW\6+[c,<EMbF@QG<?P76_WH5/Le;K_EA]c?)eN>&OEe#DN+fNad9XSAP3+27Vf,
g9MBc@TLU:5-4D;&]R/+(_ZW6eY<V>Y<#1gF_KN)Ea\EPJT4d4J5;LTVOcV^AR89
1D+Y#E/APLIEN/_0WKc#_78XP^MbKb9EM09+R?AWH_2)gZQH8##H775=^UL&5B\(
;^JY1V,&0J5RO+QPPaWHW+-:M>4&D+/RREagM8X64>bV+4EO3IG@::<HADZ2BR8b
(E#:KT[#99eY6U]<_^aNYK-[<MZQ(#bAUb^AMMZ(5a4;0GMGAY249W-5@2,3@M>a
\^I>M[?^+2<bL-ceYaN)KRNE&K&DF,F/3.XbJLLacIB33GPe]<RC#Z0NEfX>,O&Y
,+6E^()S3a=0>O1M8fTeK[>0I];fA_#2b?64c_7JZHdYQ-7=H]_,&KRK+I3QcC/G
2V_Ka/-#98&\cI6EbaIgOR+_8T.P.AK#<dKPSX[W-16L>@-[=Df.4[085K:UBVd(
/R>=K<B-J5H&)+M=T@+G@I)\4B8ORdL4F80J;Db#7SK2QPKLA9-DVY4P5WR2\5DP
/=,Y-EE[cb7<]TgF?[[?Y-W+.NT&H^JJ<,SBJFF,B(PbdS@5O(];_OAM#17/9C3J
CBb?0+U>NPJUJBEM]55cV)U8F#C.+>6S@UQ)H]LM6GYM\:5A_+fg,7C5P]\D3A@6
g/D_FO7M--0BQWAVcXT2aINbA:K66T9R3@=f:TEg,UHP?BBN=G:g[YEdK-),V[gK
WZ3Q2K7Y/-+77([eV32(OL4RX[S-Pa=-cMJ>(K^HL=<MG^U,B2Lc:8?15-/aIebW
EFF5_P9LDc-BW7NP6dYYT3IR-1RDCO4=?BA<RHKFX9+/a])=Y[X9ZV.aH3D1Y[d;
?OY/[D76EAaK8BK_?Ag]^^EQf-3fXY4ML@3T4-0C]FJ6f>OQ>@W.S#&:=&)Q>NgL
;@(9/YgFC<.GT7\>T#F1ac)a@#-4Ed_=a6V/<F,.GVH2:R&DVSGH.bJ=VKZdY7PD
KaW,S=C14Q_4>C7L6bOH2LbUcb@O39C8)?FU@+bBFSH_X#1.88O5]T3>6]:]0^R-
2&fR[AQR_Ge9([0>,KLaD<V=g\O\JE29-U^]7MZ:^H7G&0,XeBII/\=KHJ(L-/F2
;HMN^L_Db/[:X;E@SD+R_LA26G@-P::I]AD_?\=HO1RY+fb93bO.3N>&[0]-?/aI
FO\&\Pg<5^&?d3\/STE>SCEQJ\1U_6.PCTQG<)gCIMa-U7a.7gOOPP+H4d>&UF)c
)(;OIC/g5GS#W1Q@JRUe3NW9[O<?XgDTN36K26?(_+1_9cf16bd<Z>M&M_Qc?#&]
ZW0eQc=/;?4.W[?d]7UY@PYTf217GFIb0?8]@gS\dD;.LE/@T(X#R]Nf&F.2MdSM
ZN8dECdF0f6+VX)LAZ)]IL30?&Dc5e26M=-YHW0Y.&e3-JGA[RK+\IUe2,\2O5C(
($
`endprotected
  
`protected
9GMBCB(;P\S^V18ZV;ZbDK9],8YTZ&1.-0)EQ#,Z/2gJ6F9/Z8UK/)GUM4YHf.<X
Gg@5/[J^L9L^,$
`endprotected

//vcs_lic_vip_protect 
  `protected
gXaGXc:c?_9R71NU\aW=&YFZF3&1;QFOa>RA,^XV:NdN#2Ng:f\Y-(,2P/e#WDU=
PW+G?^6:WMKD]N=Z.7F(g\,:.?3/;]M[<]BY5Tf>R[DJ)A#F#+4,G_H>fCcM>[MC
1#LMKN/HX+=AU;&M9EUML^W7U^(f]WA6Z]7[Z50YR(4EI1D&MPb&AQ]KV,WM/;+.
G>S.T1GW/L3;WGeTLbJ6MOJS7-5PQa/b7YaK[][^Id&LLQ3O0RQ4:KCNTKF:<5I7
O08ecD_/34/8YKL?dH[Z03AJOQc)U;S?gVSCW6Sf34T[V^M#-AE:FFYKQ5Od4J(C
AC[<Y&fU7Q/-I1WRTH._G<KLPW=dU]MX+/ffY9UE99(0cPO#f7ea2^<dD5#.(>da
e5:KLW&TXU3.^?XEfK:V48.AE@1YH^2dc>;-@HS?[#R)?Zg7I5H5.HK6WcW[_J?,
TeO[HJGRH(\IX.fCgQAS+N5N.K3a=:g,1CP]C#&e6--^/TDJ.:/+-,Dca/O@M[dD
V<I+T+>H+4<&C6]+;S[PCMC7Q#aOR6(4YgWd:1&].3Z-MLfIQ0,_B1I8MHJ-ebH=
PK/G>,L.3fRX_S,41Y7I-+b&6X7J=3&3+I:d2>g)V_J2>HA9e^2TZA8@<.K3^A?&
0+3S[?eB>46Q94fER5J4_@d.M8aD>1SV#G94JV@+P-LJ>[^]L(C4QO.bMR^8_(I_
dR&D]<868]6(Va8HD30<)ZG7LB7HR/dW6^T.&J]5Y0(KOc.1K1JOdOHQX,G3_)),
S@Ob7:LIc.A7ScZJ<-Y=W2J=__26_AB:5V;7+](G_+SKA86;XXcZ:IX2..2D/e1M
c&+>eEXRcCFMcT[&F.&Z_bK)3cPOeUO7NY(>D+2H+][KG#R.-/RfTXDcPg]2Bb8/
d/Y.?P&8SK0:R>(=)@68Gf:.ACP+^V]aF88HI7QQ41/;AEEZ)I56Ce?+]#NZ+-B=
E(BNHPRdS;1>-<#T)KL4>:Z2[WZIQ#+d707C#O?gM0CgFR;Z[M]\QDa.IP1I<@4Z
J5<Xb2UX_eY/KQ#,;1@1&JTBW70I8Da\/TUU<=0dWQ,R]2G#FV<8ZXH.+?963cZQ
>>KaE<7N+=VW?8^C_(Fb/+)43/d5K>]6>$
`endprotected

`ifdef SVT_UVM_TECHNOLOGY
//vcs_lic_vip_protect 
  `protected
][<&N(:+W2@GK?S6B,8ac<?1L2.-EWG16#N-;X&Y?.9G(]Qe7--7-(bQ;(ea:a:8
CKePM\,;BH/R)NB-31a1(#6,O3:Oe;+fAO]?R>gWFIK\MIVWR,-RG1cQ17TQag(1
+Z[AN::TeSU/K-2?e&VUM)6D94QQ8J/Td49[?V[@\^O^8+>)1<c@4Y@ULDL&LEOC
W[N@&?7)V?&6AZWCLQYgOB:(3^E3J\/>6IC/LC?[c(ND^c<,I&/J]B63.]f7G6UB
Z4aB00ETPY6EIF[57FWL<S2fF1Q.19TI[Tf&&3N6LIZQMFc?M^@LTXK#/9:0OHJF
L-Mg69:[MITV3)C8@,:7,##27]WIXD83MV]Z5STJGCX0F25F6C9<DV:ZR10/G@<5
7gWfZ=/JCFgCg.YIEWF4^@07c]\:9Ha):$
`endprotected
  
`protected
@RA6PZ202?MCR<ZEO-_TTV<:_^O\/]@UPF?S&@9dJPg##d,ZKY=g+)e<_S)3d?WG
N5HZI6JONJUV2<c>G42dD4<:2$
`endprotected

//vcs_lic_vip_protect 
  `protected
RC0c@c&3SF:\>^8-OY#?M0^Y@QPBU4^>DHI?PRa.X1APWd@83)ZY4((4.LZ+ebba
-(0OgBKedW:27AGBB2WfVHTWf]Lg,C,1BM^VbM7^60321,c-c[(Y_:W5L0O0WB+6
5@OZS1X.&&/P9^\1]b0L6MB80BDO0&9&?LJ1+Z6&+La#+:Z;,TXbX#J)YHA-&TYT
BcDD1S02PRYZDR+1,X,NIH??c-\V3(Cf_Ig4VIDQe86K3YPBMf;C<e(f5HRE;@Q:
-ZIQ\7A0POa?(G_:egRf]X]L4^)UC-(6S2A9\eIdHRU&&DD@Da<@@SVeECf73)I,
4GNOQ^OB+e.NQ\;H[AQ:3_9?^UX_(<gXf)./(VN@R<Hc=IC@Ta@1?()KOXP8Rc0C
K?)_g,A:I0<fAbJdVaDbH=6(>Q+FJfODZ[4_X.4H<<]LU\P+R1#Z6IgQ9gZIfPOQ
D+<;]gJ)DSdZN\T@EgYGcAb8C-aW67,S5C&BF/#WK=:ODM<<QKTPI-9@DR?#876c
DAaIfd@T74:14:N=T[N3LG9g4a74Da(>b5Jacb^];;\b3&_a2E&C3&1#E6_:FDIV
8B\:YC6/K?3,050Td,85(6FT:YZJEG9@20+P+@<g;P9Q)I]X8+e^J#5;?YO@aOCL
K7Z8BN:^UXON<#;@N0-g8bD9+g=3FIg5GJX/[0I#H8-Z1ZWZQ_/[6g<AH>?CEF@S
DDH3-Hd\[X.R4@efacTY2KMPWc1N\,Q5@R@\1RY)(^TZaI(Gd(PSV-<AM$
`endprotected
  
`elsif SVT_OVM_TECHNOLOGY
//vcs_lic_vip_protect 
  `protected
f^NBESBG5#6#>WaYE]&;CG9:#KdE/HDE5Tg77Wb1KO/=S0N8^c?.+(YK(0MM:B,^
e\VM\V,6LE>Ff?F(9IK.Kdf]Qa@)TL3W5d_(GYb_48,>2LaJd,4MdO+,C)LJ(LKP
F1NQNEQ8/4;E.@7SG\,QSb&V,IFJbK@F+fK]9103A_AXC]M&[B3\]b_5LH2dYM=H
OV+D^U\f85#,JKR<6D;R,<fNXAYbfTLIYZ9X&eg8G<8=+cB&efQ4ADe6Z=H7K#Re
:5J(L;QS<0W(B,F#A@2M,X06^,<,/,NX]D=2We.:ZG.bG@D5ZRPg\dFV\.Je^fR]
.C<#b&H(8cIf@/[3=DKN,b>dJ[a]ObKXfPMA57J-(cL(84,2\M+(--0JWU@355QO
6N6S-6=c:R,J&X#cSGDdH3@JKQ,U=T8K=,O)+NUO4FW.,22-PZC=3IC_8]W99;GF
^[eAWTJ7RB<K/_NU[c[b-f0X^eePJT/MEGHQG_IP^<,<a0W\c;P\(V=BHC=(1S#X
SbA=d(gLSHBe88^Pb8\AI4.B/I=8DAF>V?)C7;9S-(I6BbXU8gBg2(;RaF)F>:_-
Q4^#WB>YSP,)c.Y20)>9[O:8(BCIDAX=HQC5eJGA[HD0/SSCL847CgEffTHS[0>a
D_LC9FbUfY&Sb]GOX)cZPL?C[DD29_HWdIP?+,-NTCS6P0S+01_F&FbbU4Z:]G@d
;<YOV(Be2P05)62UZ/X>>PH07##&F;eH26JJ)/D85#-P8MHd].GWGKQ9Z\ELbA#P
NePNK1R#+_]H^QX<G<RE]7GOLNT(]=A86dCDDYM2O=MW9PQ)7C)b<L3Qa<9/MY,F
CZ57H;6U#[1DVQd-3FS7F?9YdU_0S6eMZ;R>cB+>;8=E9/B\[+^6[/<EVE>[@GIV
AIeV=PC\UU#?^FM=(<N1aIOO^&UP(P\=<A:F<,D-CJICSS(9VfPF@70d<8.<O);B
DEBT,.<?=U+1[e;]2&6(BZ9cb7K?g\C<dUA?fa#gLNU0ZK+SZII2G^6>5(5G\Cb#
g/e0BJPIOF8a?G&+7C>b\A:/4O_JfKL29T#H\;9g/A@1I#1#RJ5gc9@IY8e_dDcN
9NePPO1,d>#b4]H]U=U9\Md-LR7K39>YYVX72H;@W<9/dE4;OZ^g(c/4=4Y4bLd<
RGOd/[-OVV2\N97.g^O0c;b.T+MQ0a^9<[=T>f?&b9TAA)W.1KCI(\4/II+e/K4@
LE@[g@?;1?]MKSa22fE]T5<H6;QR&KPYKA-5GJ>55bD8/d9V9S\/BG-g3N_G5VBE
UDP2E9RY=MYM.$
`endprotected
  
`else
//vcs_lic_vip_protect 
  `protected
8MAdQ8;\/_U5=[I02d0UfO7=)+W?@U-0X74U\\MY.R3/RB8H]N&?4(UWZgR^0U9.
+=5+^MB)S\<A@#4\<QcS7T5MLK.&XTC9Sd#@9&KJ6e6EJOdA3(N4W^VdPW5&N8a;
B7gbX.6XV8]>gG^.4K?Qc1,OOOUBSO@H]2V,7H-KeYN#NSKeO-WWF5eF92GR48@)
>6g.3VF<5a[-N]91g@g##;:KQ[<1E2UeS^VWE3[:d5D(PFfI&D=0J.gc(>#=8B,U
)Q0MG96VCWTH)X&G341fJ+7]bJMd8[6Z44;1=3.^+P?6X.g\P^N2CVBeF<9ZS?IW
cG0PB#4^eZGM>8be5e1N8eBSI=<ESZEH[A,U0E=fO088SRH<_CH1,dLVe1#GYGW5
IM0U3ad8Ga-aZT[?69Sa/;Q]Yf;;Wa3M=cYX3)ggQ;3NZ@4\PZ1F71?8Q9bN:+,6
Rf3\QEgF+AFA.3H^YKLD41V+5YPQ3gcQ5J=:2/VN0e0NF?aASF5E6gG#=fR9X#aC
b>f5SCR\9BO4/g\S&912]\^7e+B?O1+eIO<MM-/^-5Q+^&L65QQ\7Cg;VA^2,A43
=I7IJ=cU<68NWGD+20O)^Tb[BfVb5MD&cA3SZg(&-[8+C$
`endprotected
  
`endif
//vcs_lic_vip_protect 
  `protected
f-)cO)^Z3C<&F5&O\dS_J;/54XX0[eP]RTNFdI:W\O-NdS83d5O4)(A:Hb>eYXP,
V3VYVPeG=XE9D16gYZ3eS0RFg#b;A[]F4OE&5YV?65K<H+a955&;/79;D.b:<2=5
.(/>CG+PA0[G-+KQ40MA(SK9&I[V_B2>]g2ZB\1;<A0<4P(3c2a,3.;G<6RN,>.b
OC5c92.Yf?B3EQ&aNg_QIA/X57Y^^^T(CSbX5I/RPJUag_&MA9RPB9@D:@Lc/L\?
0/O10/BN5:<AEN0^MU#PP62;BI.I>E_S[-_WD-/Y@EOIPZ.=W:I/EWc_fNX6Z4g(
R>GII)S\QKD[fLW+a3eU=B+<:\c<5NP<@<8_.OG;af;#9d7?-=Y1>Y#A<LRf#0#E
C?.6F\,Z-dS4&Y:<4/F<CO3XgI]&[MAL7Z7bK2B;-1\EGAd7-[(&,YRQ+H6MM^b#
4WgM.T&2A;9^2)C,C;/]g&GMM(?MN<,1I,C5GKe8XE,UD,K=]cP^<5f7_/LDBZVG
0Cc)-95Bf266QQ\?_?^ATZ=566Z8d9,c+HeV(3]OWSfDfH#9T.cSGE=N\PESD/T)
#;3&=c^f@CeSE3>9WJM&8X>+R12RAF_2@\H#/,LbP;/=<bJUCS+KX>G1Q-1&IXbP
L4KM57Z::HcBcYcN&\8PP-;a^)W.0Ef_.WdPYJeeCeO7H9e]B76Ic@5TE.(PT\J=
P&Q7MGVa\W5G\g;ZdQPVB)SW#,6+UR_cc>eQ372:.^-73CDAU8RU&3I3^[d<N@JH
64A9&BNLI#UKd:C?7>[EZ753^CaHd+>NCFT[RfVTE^2Q()f:aINS5J+C-NVRDG;\
L^O<3dBWb0/Ud4?T,7RO7IML2I,OS,_350Q?7F9YT\e[A&TZ#G5R.WIY8a_/16K/
c+.=S].SMQMa/,a#VIBa7YbWX6AfE8T6J&4-7VTb586);c3:0bGCLgHa90W:bM2]
.BUU>(eW2H\[2[\g8?NR5EW<:O7T7T6?N_Q)34C6@4)(KY_N>ce\>2JSOLdKa3-C
F8@;]Zae]M2F/U0V/+#LLZ4:dAdY\OCJOcUMLNAZK=,@<REW\e=DeBAXE7(R/U^C
:ELNLcPf9X?Nc2a>GQ2?@_Lb3>3GY=_6gAH\)=SRNGa&J\>F5E-eJK#-)#QICGUe
OZ=+TI=APV:OJ:6cb#cK80SGL668]O619S3T\aF&Z]4aTYOa5DX@T9HJdb9)d,=g
+a1E#eWa#S3EX\O/@V?ETI;\6Q9b/5;9L8,)I+95UX:DW7#fD@F7^=?&+-?gG\]g
@1R8VQ/8Nd2(62XZL#9bFaT-)ZH,_bT#QU6.WD>90bO7NE,AH],b.[8ZD4TYX<Pc
.4V:BYQ],a50L[H[f8PI@:VD:\E6O0\#@b)8^aN@EfcQ8b3dGeIf-g6cTfU\2<^]
8ON#e6JcM0afDI;^[==026>.,6c.(2WIac/);X>8HRN7:BW3CD@#G8@]TSGN-@Z5
GVf<PNK&_]--CS_9I](MM\X8D69e25N?0fbCIcMb&?9V@2MZ-O7B6WcO@/^[Lg<-
L,E&b/?XB7LC+WZbcU>-4Jc4(Cb.XC/XedQZ(5Xe-8M+Z\?L^=aEbb7N>(];4VLR
WBWB9Q3=)VHdFVPbI)_]:-Pf]a(KB0<NBBc0&\<-ddT[DA6c,cCT2:@cAb4#8K;]
&WLZ:aH0GeR>_YJLL=3f-_U9N\A8Y7)_b<OI(QI+f-#-<dCZG3J-^@O0,LGW,\,6
gU=^6Ge7FbL)VW2=T<-B,f:0-=Yg^fJ@P=-RF3TaO&5R&W7;=H(J2_[<]EMCC(LT
;B&FO)BMAKL+cD-TSZEXYcNc_S8,)4cb0847G14)-bZ[9Q&S7JgQ2JI4LWTaV&D1
0-L>4Y#<^Z91aQCT;95+-fZ83ICE5cV2K)a_d^_Ag&ZN0[??1P,2MS1MNP<>FX;:
9Y),.\d8RLI:(d9)0+bIcL2_F2O-MBVDEN4C)>fX-NVASG5LXFN)0^WSBLCQC,b,
I<@A?_6)+0.VcWS8O[71[ZP>J)/c38_H+_HQ:R.:<_B0H(45=;4f3,Q&5Z\eNV_/
b7=WHP6,E^V4)Qa0RQA1+Rc:<c3_\S/)^;<VU\F;P7:aEaG&3EMGHEUM-BHg-Z@c
-)aR[RR/)[X72C#W3BGCfKVT5LfgB3M-YEP=+f_F314M?=XBD\^333(W8]-IVQIR
I?C5IB:&IMH(05[.EaDNfJd5Ie+CNI@g/ZgFYW)[X4777Je#Jf,BIe\8Kg_Yf[Q=
g#;\4YY/6?4/Z-6<>_<)LG<MCTPEdf>W78PaE081Ac\I[)XG48P4V/923Pe?E^g7
C0[+A@Ya4460K)3K3eX[0e1BcW.P:,FP;G_/\[1<a(L+/82A2_IO=8,7]EN(>:L:
gDW9//#K:g9IP#e#?RRXcLHW]D)K&f,#\Ng?]>H+H>NTI:6Q(6>fcPBG5:43bSD^
f[gCKD?LA,A^.BS\<d5J\26[^-S1[Af)MVa-0a?]>L8Aa7G4<8^:^cGMOZJJePRd
WP6C+d_X:J#-(D:Zc\ZD3PD^&611?D@(>R@V#f5C.B>#1:T_>P=G\/;TU<+g,IZ&
e,57)YP0RAP)7#-L)DMeaP0g6?)LFMdE\W9D;1TF@]-f#2=f&,KP;#NeN-2O,UK0
6XLBW<Xd#f9g-OU:5AH&HL\J&#J.Y1-_XYDL9K7;75ZLCXA@?cGQSZCL7ga/<.WY
:>=<;^.6PDQ)X@DNa-O3#ZQNAIHa+LL]\DLg)1ebfQT24IFd;86JX.UROgC4RG01
E6\9=54I2BL;(]J/&DfZ\UA<YQ3(^;8.T^K>1TAQ:-7[HTF4T_6:H\[Nd(W1IZ5A
5Qgb;._LS^UQ@F/:bZZfM6WcN5FReS[;b.4e[N<d9<KQD_d=DVLO@[5E84=g1?U3
g>Z9gR/=?E)UZ=[=AR5U?C<>0&6S06aYOZ&ECN2[)L(,e#LaZe6-P2UUZ.c/1d>B
aI:YAd5N+@2RU/Jd-cU#TeS=6HA4e_AP<WQb_EVS0+UbB-Y.U,X34G)(IF?()G=d
(1D2C@E<Z8?CRX\4W1c/G/X9RE#(]#>bD]PE-bGVdMM@)CY8)RJd=#OM4V#VI>D-
YP9e>&.#=&<SHC]+eb)eJSQ(DCZY,OWQ8B>aHJJa&c;6F;HOHR^XW6;QG:AJG>V4
ffM3J3XHBD:S)8Gb;CfZQTH\f&g8T8,US:Y>LEX@#Y+^KR+N@<@NP;PP>QL(gE.-
c/5Jc>#CUJYBH/MD.EeDX=462+PWN0HZ<f9T_\#A[dJf<Ze&TLa74I<4J\RFS45.
dd\Sd#+C102R15&:]X>Z4&+&TZ\[(.9@g:Y6EA3T0(ROF88TXAeH_Ug7431>5:Yb
K#f.aeM7\/C.YDD29YR8d_&,NeeGfU-,FTQ8,>+;BII@)=ga;TGH4<c7\^VRd/K@
d^9HMW,)a+Z&#R(SUdb6aR\&H#16XP]TG<<7;97JLW4+^4\AB8#<?L^WORIDA:\d
ALE5S\>CJ)FFgQf22&AHZRD)De3P.N_3BbHf6K;]UgcX;X;AHEBC5_I]P4X7B^F9
]+6)UKQG^bX(1[[,,JN&(Y,@0Z7/NK72D7I7>&Ea+de)Z[Y?YB8Q-A8:-]2/=ER&
>fcGD,@^7I/=7NRdI^SP0>I0VXQW>24IU_HC=g#S79\4Z6]/46f7/Pc#9MK8c7@4
YU1\b/9XY#5QEZ9R8;@R?.d6XN;&HD.6g(U&UTDAR+,8fNI?3G63&=:179587]Ng
?dE5D/J,U)E-[[gO56?<c[4A7D67S,;GII^gNHeG#4LZG14ZGG02OeB)KGdRXOYE
;3@ZV?FKM1@L:-;OI:>Z?OT\/#be0dN\^TFE55^QBf)2PZTOEIe?bY,]YDZ[ScMB
<LS7PA/Z_78KBRVc&FZcOKcMb-&X.6[K?=5S0YXW3IQ8=63.NM-f,#bS_ZB7ZdT9
KUIFQI=JDQPW+aZ;Q:1M]>_30BY+UKE<(6-9Yb\E#?OM:eV?=b\<?LZa(ZCDT&/M
JLa<(^+]K0Y,e6/=UHKY]D#0Q<:J//RA.=TD-Q?/R)4F#ZGN^L,G+G,)>6[=;+F&
.TDgDeB@c2ODf)X4@>2>?\I1VCYb[/GY2B(T^T]g-VXJWFU(M_WOeJLFVJ=G+@GF
-PcR48HOdO,1,gD627>5:3?XO,J;7FGUTRG2N@-DYU9H:9[/#B/5B0I/DS_KT,IS
,V_W8/gABSXI4=1g;dFg;]c>.=4M0FAeZC>,a8OT^#+NVGV,@^7:LE[@,&5&\:B6
IPZNTeYa\&gG(&Q;I)RI03dLRC]EC?SZ_MA32G,KQV1VY^N5\eVQO^,.D(U)@,<f
L1TbF^(-J>JQY-W]3#]/5GLcT0\@\N+cDNC+&F0P=@Z4b[(UXH.2E&cM.eKLDa5-
KL>)-Rdg&(6O1,UDS(.E,8[&a:H(cbBaR#<#\5H#K3?WTa7CJ1XUK[Hf@/AO+::J
5aV.;[67fR8R^3@02.YcIKgYE]0TC.QLE1G9B9BfHA7CZI?[OIJf_T1Z:IFH)0Yg
(1,5aW@37fHO;0+Z@;HL;=YSc7OM,dX:J>^^S>W_D._=UIbgL0\f..]d7JG19W\C
QM?22BUFOf86B#cZZbR-.>(]=_H1?42FK#>YUf1&XNF=DU:]SIVGgO_NI4FPgd5C
6[9SY[_BO;DE/WQ])KWZ2>7(O//.C\3d&JH[M=4bBG\M1Q34dXc:?F/B^1Xb/Y8a
0PNK+&P:4<QZ\GD=>CBGMPW4B[c[G\M7Q9c+aN&E-6P2\L=Af7UR4@]1H)DIGE5I
0=,RcebP;>e7Q>bT)^D6c-)_G2[X)2L:,&ee]J)eU.g#L&]+JG/ebT?CIG(3a/_>
Y4U>N?f6F.;aUM3XDeTBG[3Ca82aZ[W+>>_E#WG1/;(8/FcP<cRO#.E/200N7bE]
#C6.OLc(H2T61CK]Md0(+-_S\c3g1/_U=?0(H3X;IU5?:?FLUf@a=BUZ7J:<@MWF
.)M6EYF_X&N5W=e)FD3Vd?&MS>-GLOcL?dTCGLXLB7QW5.D=4ILRba=4>)1W1E:>
3S>Wc>X1^\CJ37)V8KE9S?N?7gPP90H999JgHNLP9Z__MQ92Y<^cdQ-&1bZ.8f/^
N8?Q(d<L95?X1@Y<;0[c749BR[b/DLQ>B.R-S6X^GR0eW3YPAeUW&-f851,KDW#4
0Vb]0?Q_3LIF99R9+Sfg5N1E1LUgQc/D2H(F/8>-EH#HeSJRNW@T:1JJV:V+K8//
d:H52YS-ZY;Ef+0O88+<6&4646:CRZEDEe=(OFOS:)49A]]a=C2a-#+<a>,9g>d-
]N]XXf],1DITWA2^ZG/YQD6A8QPBD4QTNBd:#YaO@bJSAU01MX]=(L8g#9f9IQ#\
]8A[1ERNGb^/&XN7RD/-+X/B8E+_Q>6bg@V#)89HYB_XLg1-/<UGCgK1SU5H\@PD
BT4+7VcB(bHC\^8(?2^J5K,N9JYd&2]NJAg4bGYa3LF6=bICcb-:-Z_DV^:10b0F
EL:19GZMZ2YM7V7RPX.C8MgAgIV1G2++Y>=d<7a3X4/P(_UU]9\>P90],V[_b>]\
\_C5A4f9GKaKWA8,<H)FN@TAe66#K.0Pe6cB?APQ9L259TTUY@DYAaG:=UG;:Y^1
=5Yd>O>2/TQI8UM9I=?0Ca6F(JCB8^)\9)@2S&.,[X/JL1\Y<FXW_&2W/)FX6DS@
O_;/W?IV#b#)f:)=JQbTEdBQ?a1-6B\H(=J:ONPcQ]]WANFM<>30F)-beT_,?CUR
/X2V?MTHZ2>+,7;fL1>fdSL[(e8cdE+XM[/B><5CKV2#Q5N3BG1CXc&DS7U;2W3J
XP9;d8,_N/2HEE8_FRS8aJLW;FC75f)A9,MII5#KU]B(Z.+BZNf4:>f)H:)@2@B3
?#2+-BE4TG9ggD6][SMIdX+KA]@P9/LM3O&EGWI6#J1LJ+WKc9J[S_USYR8QFB_R
e#9e?R+_#cK>E(RC0,A3]3[L#BDe&PbgcXS+N7:eDJ4LQ\@(RL&2X]JG(a_4.Bgc
J?(R>F\\R(B/GQc0XB\OI]df97A.2CK^0/@-=W)A-/:e@cYFc(RJGcJ<JN?3ZLEH
<3I:fbW>^?Y<g]]g/VJMR.8[,U32(..M1VK6(X(=687HD?IF0_#d2V8XP;U(KfC@
S89aH3C68Hg=VDAQ.V2J?&A^+-A(T;8)@Y1&],D+d/#-54BI@X\f9/MGD_ID=FWX
(5a+;CdFT5=TeQ<Iga61Z/Od=W5SBZTP@U-WINQ/HQ:-&d0Rg5Y-1Eb;ZERa5<DK
N=AHXU9@<bEV,;0].&V;CadJ>a<0\C4U)J^VO3Mf&@ZH8YdaG7V.cUeDYR]g/H\2
I[3bC3Z[L,^^Z:PG7b^NT-dYG)UG[JDAa:gf4XIeMT@SLSe1QWZ6:N-SeK-[A3#@
bKJNQ]XgeYef@ULZ&g#HEf6#NBR,]4I/M6][07D=^PLC.5deBF&V=3H.+W@\1U0#
6Y3gX3gb;2P;FQ_Q<,a][&3AV_TSVacR>B?d4ELS17KPQ29Og_#B89+^=?R+K>fM
IAd=;Zf-Pa7MbC,dOg>U+U(;WMOE6;YV>OKQ;_b0P>&Yd2:FC.B/JF7RZf98_TP7
X4=2>gf+AW.K@17O#aZA98W/H_:#>)Z+W#0?a(.K]45J1]f)bV0#G[0\S6P6EZ,S
^_ZfN;[,96Yab/,8eT]HMWLaIVKIad.\eeEe>V8eBFebLdK9J?C0PbGF9=@Y6B:^
(-WV8[T=(Xg/3JFT\)<6.2LK2]:1]?T:<e(Q#Wf]X12H(B.Ybd_FY4P4g,S#c/WD
SF,d9:.:BS#L1fH)F\4.X8M#_.@FQ/QHI/5Z03C?DCb,9L3?R8P5fbGgTZ/IN&J(
+ZS?PV[(K_#dG]1<])3;K9;Z<Y&((16K&(LIN6Z36d=RXd]PIW,:P_V#XbQM17PD
0W:d-Ne[]aTH@)W?L\16)XE>Wf\(BFFcJ0C5=0Z@(FdcFVLSWC^C/&([fHcK,14R
#R;_eI=MX2\04N\9UVXR2DSOS_MYFF0CA&5>N94e_])S.D=C[?18,/,IXK?X3.>5
9ACGWF\5bLa&QIb+4bT,<X4S58_<DUaM&SQ628A]WbK-L#Bb<XF(g]BH/aQ_(aAf
?-e=#&_0.=&:EB4LWHS6He8[+Z))22J=)[RR(;cS(X>(c^0B),2>CV\7(#8UfP9/
Q03?]4C7KKW5K06d.Oa40Bf9MJUV]^67UHgB[)OQK9,TQ3bS@<R=\KK(0T[8XQR4
KO]<RA-SDB/FZU^V./Ig1@NA4-=#E)2Sd@bfe2<4NRgQ;dcD#V4EbF&&J-\gOMR9
]S,\E\Ggg#-D_4FcTQ,^H4P@V>R7<FT4Q.CGQWT<S=24A^7OY(VJ410(@&JgQQ9W
eSPbJbN>f;AHX12&_Z<Le=^KD<3(N\LTaW1gD/\8.&;2b+&M=D,+>;;Z1OPYLfaN
&2bCVT-EDR(EEG0cIM9W-ZVL8OOR\<R9B2MJe4[\Ma[2;?;P]ED[1E,_aZeMR=\/
F(#WgO)1e6d@Gd,&A2ebT?4-gR0Eb\0b[:CF=]1RUA[F._0DW6;][CWBWdJCI4=,
.GWA[f=W:[aLKge(\/=/(E5CJ30F?L?Gbf\/#RPTML-J-J&IgM0e+(EG,BD;.5TW
6f3+6YNIdHTaX+LKY=ZPYQ;DJD?U).g820/3JM#=0)>&NOC3C.a4J]E\5De5GUC]
(L.#K.,@&4<<C1)W6=KA2F9X+Ic;c@NZA_<@+EY)/c?3SO,WX#QU,f.+TeH8JU[_
WN\33D:T#N4)N14BCcdGHAK?A,I&<L_S4R-g?#R0=:?SE8:9#ZU][@IHW]3SW^Mg
0AU^Ze,89MYdA>]R5cI&>aPK47SEWIC]V27=]TV@E_PX+??#;)1OW.I<JW8)G)/@
EX=5=_E2K[La^I9O3Qd@AD<MPF<QS)CVXY+d33&@GWT3<\BPRN&P,-5XGY8&f.=(
R^3L@Xg7;F>ZJMQ]g1?_3C8LcURR123b-H^OH75\(.A5#X/^[A4bfWX8\,GJNe(4
S^d:[+VP)7.Ag,(4_3UF#Uf0MG3?(;=JIb9E,:E0,HD561[JU^UOUBKXBNV9Z>:I
Z1\6F?P1cO7b<.+++)Rbgg><Be9)0KTNF:LX[[:VR#>//?V/-ddZbL]K5,T>TUBf
ggQP0[XX\aY+GW>/H/d204N6gfVN[;HdLKPB^WDV[/1NO[#X&Xe7EL5D]d&DTW@b
Y1D.+7QDD\JbV,gJc@UO<EZW8[,<G(GZ;/S<?UEQHC_.YcQTP=]WEY[a6=gOa[d/
O75(7GRb8(^7(^=EY769GQ05[J,P&@J5:fcPDW[B<9SWO\3(e31&fU[/)X&3X+3W
.)W?A^Y;+c;;U(.N]LX4#HVTT:Uce[+^A@]#?8g&acZ7I:fQ0EH5:ASK[4?SO@PQ
D\LEg)^>;_/S+g:X/R40Dg5/E\R_8Sa?>Y7D)Mf?:\KO>]&9@.\MWdCf=KOJ_QDc
d/(\E/#RGdG5UZTRKV=?0LZAf4/?fKF]O/-JJN8YV.CU>cDJ7Cd,UGFD\DbP_:3Y
>_1A/?N:O<TPKefc8g[ERW4TA[=b,d>)dM-gQ#Z7XNGF\M8R=FB;>-PL]>EV_,fR
4[?>)Ma46OIS(?;?-OILL1bN,OAdNMV>#@N^a_H&R<=9d>1@Q1)Z&?cG;9>6G2^]
ZA0bCebGaaWU;KZ\Y0H\NGfG[@c<-3#.84Z17<,S>VKWQPC<FZP:L<)X-W),;C(_
LKE.>,<G@H(H1O1-ZPSNcFCJ=JG7G_A(@cc=G7e9FSCKL8d^.YM,#BCV/C;BZCa:
^Q(P]a<5_2<D#-gWRAXH)63,TC#]Y/Cac>gE3b[=J]4(2UQ&fAAJX3TaZQHQ.OQL
7+H)YHZ=]R+=C]BERX<K4Q1f=OC5dTY?)PaY8,=gGVCD,dMQ?#P2S2HSCAbAL.eB
X?YRQ:PD>]V7QBV4/6+)W\QZ\PBW+UKCg:+F+IK80a<c=938@ZZ;P[?,=eV?E5LG
/CV9bQZ.JZ[Ib6L_UcVY7Y8(V&I5e(LD^HQ16RO7C9PZR6)+=>IXHN-5#/SE84<S
UCUNRb^Hc=AE\Hf]CI<5a\OJ4:\<gU5f5.:.+g4aDR)-I97D)C&ZRHe>BNaX)0Gd
36.3;IL.EI547W\:LO@Q:N0#MJPPF8\F&eQad\U5^WPG3IB0DY.b]VYXPUg0L.S5
DBGaDB(IRIN,Qgc>,^@1)+P8eN+\g2B;_:P./(J-ROCe2U8NP74D-]L.>(=OC-D]
T5(ETeYR(D=-OR])^[bS([#H+4YaV/62:PZRfF]Y&c.4L@Te<b)@:EY6,7YQD3U.
S>8M?LPF9,LP_9@),M;ZO&1I4R/D^^dQQ?5U5ADgMNPW_M7g]F?C-7,<JJfY2EA<
X5aBYR34DcYE0EA=X:dGWb?d8QJgBEV47f+@>b+F4E_8X9NCKfOL(,TL?PRZY&?e
[e==e14X6c=BFOb15O)&VW8O.W8bUAYFNH)AIHBB.3_\.Y)]:>.=;G4,<K]N7M62
6&_>[RN[&HLC\[]?+>),^YGIG?G@1bI\e0F@Cd\BF^)(4eDF<K/T0g=?fe3(.C(C
97S::?1C^+Z8JH^3/f\RaGN#QRQ/Z4d2JX11dH\2PeDH)LS-XD_7c7A82UO^d>7g
NM7NC>M#?^REf:-Y@QX;P9KWdIcVcPKKHCSN2@PaEP&b]YGYU.0,Y<6<eL-M;O]5
DQ.HY,)2/F.7f@G^7f5-^9J=H4,=8OcAe4Lc8CKHK>-N1cG1&Z3Q)X3N[A0S\6J)
<AZP<@2_OIA&,Z93IJ@)M2O.^a.XFdZ;,N,=\Oc)WE@d:G2WabY<#:#:e2IX/Cg)
_^RE[dR7S&[PYV(./fFLUb6KWXeg8<F[1Y3)I]GP6:FV>?b?N#K=bgLYb9HcN^9g
=J=24U?Z5cLcUd;c@0g(5NdH+B\,O88c60;4\\@3DId@-a0ZUCNfBDHfaZNZMSUE
,SHT(M^17?5T93@C+]0T^O&/#WS#b@e=2LEI6_]P<aGa5IFF\:McC1Y-QgJ?SMN^
@F6.a^WJBV[3aYGFIO_;+-+T#309BcLT2NP&a.7TW?U4-I_1g0-:R>O_[M/=f8Sa
HF[X#QLKM(;);QgC;6UCO9DBMBK^\2C2[T/;BAN^J+c41M#42ZM)S)gaeMKL<&01
bcNNX5RF]5XI&I4/#^5#AEeFUA#e2CEI<c_<(0O=F::MSGIa#S_ZR8G1B.POR2[C
1<R9f0,K3eJLCF,+FDg9gMEXA<JW/\SHGUa,8b:aWY7e=.Y.=^HfDf?BbR)[0_93
Ag64@VcCVSf=4eM>Rf(P&;X[.Z1;CRK;0-TP-/c\D@feB;Sa]1:\.;?Fg(4EG^0+
E707P>1(>#MH:]H9G?2QBW\?7LVVIeYFLUg+g#EU,WfNffPNLC?\LHMb0NR,(=N-
W]>K0&.a#g:[RL3P>Q4b46>(X7Y5RSLRQ^CW-WD<bP:d,Q@KSIdM]H/8IS?:9LJZ
b9Mf2^)R;8fI>2Y&Rb?GTL7/R[-#BHGDT+6QT\#D#+aHQ^9QVI6(,JJ&1-R-1[R1
J(2TA=:KN+g??dF<a3BPc4T9&:TbJTRQ>+RU&/8M+8=_D?YH?D9(5gbUE.D\,aKU
Zd^PUDS?(TATX\1^FS8V(;9;F4Pg\b[f&d53B>EH9F/LUE^-;FGY=E>aG9F?]H.0
EC+\\@J3[.]Y6G[Z6U)ag(EDCWP^]Y5#d1A.KJYVbXY[1aLNGW(\8]J/e6?(X65S
457M]3fLXYDLbUBL_W&AF-@,aV(;XO+Z^8I<UNR-4=f^Q0e2X\e-#bd8)Ib+]gC^
42/#Y\Y0&fGgJZcX+dHQDY;U=L\Dc33=^d?RM8Q9gEbWHL27gIAP,V>/OQ0E7/c[
bIRg2-K3H_I?-M\Hc+TEd+d_=gb4:44?XN-Ue;]gYaLe@BLaIPZ?BL@PKXVN,a@(
&#CLe\4XdJSATI^?.42H;.ZC),4XRY_VJ:d/99]=1R\IaD@@c=96GYe)_a.O;QE2
F>GZ0/ZAO^a^6Rc8+FXO=6e43FaNc82WU+)@;8W@bPK)FIFBXO:?8feaYD_2e/@(
G)Tf^S8&8#6?1E8P3QS0-Y7F6.e605B/gU;dbN6-A2f>b<,04d1,^@BD_ZXRS^B/
KcA:WgEKL-2R=5(7cdS,F^ULOFbW1EMIF7Zc=;.)T1=/4@A;aXVR\E,937FAZC=9
^[;]J?,UZXIGZ=::XVIZ<GC[9HffdM1)Y)+@P9aD#eFJCC+d-F&+NIXGLRU3EU:C
[O]+#b7I=cP#9+a;Jfd]Q8RC1F:E3UK-[<X44F;NG@@E)EQC31[6C#_?49aFaZ[=
)/g@S?<<-Df3b/Q9+KSV>7EIC_,:@K4,Q_<W6@3>5dY1F73.PXc7NLG3Vg_V1eX#
U=C/2gBR.\(eSE2DY<TM(1(aHK:5(dGK]Ic,,6b42\JGI.#_CWe;,P0=KF>N]9T.
A-K0=]9Vfc]1L#[\E,\/5?I0Q,[/5N0BENZ1P\M<#(b+NEc<[LGfPaZaQ#8:?^78
HVYU:gT]U&d<cF/L\ZVHgWM)G\^(=>/3>D#RD#P&@[I[[5VC3C6&;Xd^f[Y4@Z6_
aRQe&1=4cJB]bC&&>a_0K6V3R7-6M^O-Fd_X-L,]dc3eITad6_A^X);c5P/MfA<,
D]V.J-gL9RW)dLL:/5V)08/_J?KT==ZLIJTE3b>a@LW:JMHa:)d8.=J?=8RCOaWM
YT4d\/O;2)S-8f2=\(R2<=MMQ6);?cF5PURJL3)e,76@+M/cL-NQVLNc=@I,_O:a
4Cd,Y,+;#He)6;@WIa72@L4eL[D:2N]OeQ/H/@,NZ:Q,D/ULQ(B@cG93LN,=E;#@
9GC1Md;#>3@Y_#CC4EM/-A45JXAFHEO=:DS?P_^QVAP-L&(fY3H\J#F^TL1ba&]6
#FKdf?RB>d?/&\eYR?XVF.]MW/g3Z@DAcE2H/G7OA.BK_M?>2]d22\5)\R&c=K#)
]1U3GPUI@]U4ZE+-QFP#XF9&HYYfcMD@;S&)?.HFHCE5aIdF(/LC/#6DJ8V(^68/
YO;dMS8@aP]XOO&()K+@f>J4,K#QBNT2B?;9&SEF(]?g<+L/e3MeK.7MGe1ae;,e
9e:YB#9J1cSGQQ3#ee;C-;SE,+B^UF77INP2J_ZE>?1bGK7UD0Y3HUb&;E#^V-.F
5M>3J7d(2J5Ed]_QOb[,d1N?&db./\5&c,KLYP+VZPK?QM\Y/PRUP.Q\;d^,G9#4
>RCF6#g7.AZQ7JDD2M0_;Q^C4I;RT&bB_<CbAa3\]a[7[<G;:aS14dTCcU(YN/Fg
Te>Lgg[;IYBYA)LLD.3=YcGW;6dc9MX4WNLd)9FKLN/MXXdGCLSZ_@[98f(1268O
899Y\YT#TY;F(V6UV:HgHV4IY\)AZDX37KZ]4P=bAN6<W@K&dM@87]3/RbgAX)bS
NS0S2d?M:68/HUWN,SeKP8NI[dZ2Hg5NV.d7P^O+6(R<\WWfXX[#\4#T=@G0[102
V\;GY879TO,-QIfUHM7:WE@R_Zd,J>Qc@E[RMJS+C/I]B=,e<)RJ6)@)5Ac0,I];
aBH)fT0=OBg&L?]XQ>FO1]8AO0>J2_>?5I_GV.-:?_?I0GDOE0Yb[\,T)<9><Q7Q
R8UR.M&E0NX],F1(_>G2449gI+;L=H6Jg47^2KaaB@N#IgZB++5FV<P(>D\ZEUUV
>O>A&11@MDU&&^5LB@N&^#2J3>70)Q95f,2-[g,,5\Q[W6>@?G[=AMJ[2WI?I00R
dJ/P@NULK#XRYQ,:c#?BJL><D7Ed-KJ/Y0b7-JP4@Wg+_Z(9^-):?\/Y=YDZcN08
A-/K<-?GJ3(2<1g8-MWHUH5c8BV]91W?,L9&VPG5)78]5HUT+c98J4.[><X>I.K1
I-O0(c2-).f5B\<489<SU@g[dTBXZ#:ITfAQ^TF;Q)4&NfMD]&J(=^MC-I0A77WH
HP=A^58K/K4eMPB<TA-@bd7X988LKSM+Y0Lc[^eDe[A[;495W5T)=>IN<C?4U=^7
_1L,G@6>ITF]#e.94Od-R)I9YM/.=];Vb&:?a?K(LFE_+g5H(bGOLSd_;8cS8AcW
P)VD,\6Ga059#fDec912GQ^KBAX+(V8-&V(BTW,&29>2R2G8PIEb1a[Y-:[(7^)f
,f14<9eg\>gO)QTD715G&bB&5+NbWUQ8Qc\6I>;@9BCPd(-+Q0LW>):D.DAQaW0W
12\JS<()_;>A?K83^Y^ZH#+-#0(/DP\IX[LJA?YTCNMfL=^;@Uc[BKQ3^9[5I0HQ
6FD>2,@^a#\[f,0-)XS1aP8UB5S:g84:42\.P^S(\1IF;ZTN/=I2+g)X]/@98e.M
KY]aOV\__V;gFb2D0^14ZZ5-_T-OB@&EK[c.5I[-K]H83E361FbYP-Cb;MQE7gTb
^[\ef1^&)?]):XAe&W)3>1L7U7RU<^9,/GK@3B;3L^WR4aa>R7e>)@gM:,#K^4/7
K/2]G].fVS?5^+=SCaBefVB6Q6755<V\:6IOG:4F&?ET;;2=&/VVBT])T/e@=;.X
JCRM,P+M9/>NSO88P0g3,N.cHX^>9@67JM^1J_2.R4]GL;dd=W0ANAcTK&Yb7P.L
O:U4,6W8,0VDFJPTfgd+X8dG1Q.X9FCZT2=:BJPHJ;R;SfDU^TTS6#a9)P#ga(L-
R?b0M5Q6D(A7>J>TGO+>=^3)-,1cBI3XY-@ffd^G_]H/.)?ZY#4bPUMcNC[..?(:
W9I-W;U?2<=4;HH@:gUZ-?.?<?ON\@(,_]N;bBc8gZ?BfJd<98S_HX_]O1)Y#&F[
(/?,N^&VF_RN39\XO)P3CK/S.R-cg\]X?[0?+2?B&Qe1fF&><]K=a,WV@0K0AX_&
AK-Y<E+33DTdE&Ea4U+=aJP5)3F]3Yd#@>C.9@?7@L5=?LZa(_WaD@XD_+XYG1\7
#>cBc+6H,H_S:(9Y)V>?[Q^e:WM0:a>&0DSONMZN2GE+IJ@<DV9]>e<K,>c5Y.H@
AS&D+7I/-E.3gVY7.DA93]_>OBG=,I3D1.Q9XCFPXJDP5T-8M//ZQ3g0cOO/d(M3
GHP9Z&H;L5V&D>2ERcBY24cV;NYE&30K7^5B#[gYfP=^[H=GYfBgNdbZ-;#=GcQL
<@6IQ>V1Q^?a(2eXI-??6gAg<1D=GR?McZN5R&]fEJb7#C]FGT[[9OC;W(_;OJ>2
_T+bGSR64]5ZUZ]IcG(8Q\QZdSE2L?^(EUA_Q3J+ebTUIA9E&.EUS[Z;>>c=b[^g
X:B22abgc-IT7\E<,<@A#-H<bAWVZ78E#RgCR[C5N##EAX@@8GgJ]T(T)60EaPgO
-fYRPRJYF[YUIJ+Bf/f?a)L-<(g24)BE>P9BA&\6MD\1W)@S=:=@QX2AU-a@/6B>
@)J3+P83?Q(R&@TQI=VBK4FXM1@e]aR9^4TS(RaN/^+-POX4^8\J=&3Y=_\DD)+c
@0=&,NF>WX?Rg2TU0(TIbWFPRS+R2?(?N2^VK[YFTUD,-KAE1I2&JQ2S_]I(Cd_V
gd[.(\47Z6[0LUO>-2,af5M?U>&<Ze:KNO0]Y&?(V@23#5I>O0eB;aF#>[5CIII[
;d0IZ<5)XXEbfY;9eXT/5AAH_MS/[M9=PcTKDI.=]#,1a00KPRW+7@d9[?E=VX2&
CY-BPL5&-.;SIf5g:ZI_K@CW+eB+8H2Q4&BJJ2B=HAP3=_A\G2FRD\2D-[a4ARDS
EOa+&CdBc8EY_PF97V4I@=KfQ7_3=/8>0?RO/B,KQ^R:\Z,ZW3[TS#Kf/.ZZ<YY_
71#G#&MG9gNG7eEge#ZZC_=&AEO.94#;EP(a\2P5^A98NH:SBZQ:\0CZ)e?#d+[M
9\&fMeP@U#L8L0B4#bWY+3H.3D;<+OWBQQMgKXZX^J&4TP+-=DBZW@6eO=A4aIAJ
U[NbB4a<6@,62[3R4+Z)2BSSdMbBV[FZL&TeLC75PLMKORK.WUR67Xg0fWa>1)?R
&X<4PL6e9K-324ZIP)6;D/?Y>PK#K8O^aSY4RZAX6&TMB_T5T&Hf)^6.>0JPMf,0
;YE.d88?&fJUO-W43Y9L(3V[P@^])^XbGR/M.VHZNMeKOEW)#_P[5)C5;BA1>3)W
N<.Ra124#/RM>8G^e\TcKc\[RS,UYCX?2R)dZ<@NF8=GX(((#)B7]4;]@;E__ZM0
NZ=.^[G7/K)?@;-U,2gA.b3]F[9]^G(9E:b;a8)<>Ye++<&)AZ)DbZ#E@]Re]Rf:
U+7ff;LGPQ;7CB=#=cL>d&X1EEUEFI>2)KR;G9W@eS^@)XSfF?IK>D1.&N_I/UWM
XfU5#NC[b_+fQP)C)+B58?d#:8WA-7.EZVPV_:;L6JWB<)1)[XU+E38JaPXD)ROC
+5^)1+_RKN_9U3JVg];AYS(a,U.M609RLe+Be:ITWU@Eg<^,d\QYR6&fa\DcIfGG
J<<EXIW.@FfK2baI]EXSgP3CXe:+b@Y4VBV1)80,Y/ZA]XfB-4Oa50b:M1(f7FS2
V,<@/ZX\T.PQ3)]g.4)(;)9SZN]AS.X)W3,-[E&OZW(eYaQ6ZU#d-ID5]3IN6SFW
D#LRI[D[/(R46eV9SH_YQ#P98J?g2Z-&(c.#<@&2)=&XJY:<U,=4:R.1\47\W\84
OFLN.G<O0Yf=aQ/HGK2FKQg2/WNPUcEf2c_:PVCFEREB\/0.&[NY],1d#1YbB?Nf
+.f\E.)bX-b1Xe6:+\A-VKU)V?fd-E(M(3)753>I2Og07XXF#&;W,.7D<EL[81@P
=fZI:T[H(_/c[f647DIRZ[/a1D@J.[J6G4&U2-I&e-+J^I&Je\AdG&WYRSG\f0-c
))6T@HfX6)?V2/@W)LIAA0)B^]V47QG+RZJ-M_1E[;-R9@A1,F4#egV/[L,F@-BE
Fc8148AGCIb\?1C8)95;^P9O[26Bg#@/5@(fC,3[R.[+HFgQ-_F-2K-OA[^eHI38
BbTb1[MW7(,36b9FD@CaKD^3?07F?de@WTWGG+eG_SYcc^c/,H>=bLd/H?+7C(d)
>2P06E\?R]?&MI(+)?[.T]EW-2P2<Rf36/e;?c>8KLN8Ad0)&&P_VX19SST@]a<L
;;O2IL=cffJW^GGe8YBYNb<S9;R@.EOP,&<?\c&M9Ne60Zb]dLP(CWfS8RPP=g&T
G-(Y=ELQa8[NBeL#VHQeUcA[4B3g)Zb&f=\D(,CAY6Ib&Y&1c,6RBY<>I:U>@[/@
[<Ebdf5CA?QXJVTE]:E)MMfeKaGDJ8)><K50D_-Zc1.2HQ>[6T/^_8DZe\LV5J2?
@J26=Q?FJDFeG=8(D?E3Ta3=E2KYIfC+-5CXOQIE/\SSP_<eW-cgYE94#@0GDR5@
5fAMFJYN;:F/Pf\WZb1/.Ec(TA=FRT3,2NUJCaY_(3N1/0XKaZ^g\E-&(99g-3>&
fFZgRH,))B[H2>0]Ig,-5M<-8@M^3_/7Qb_BIef(^N@NcK?],U.3X[d8c^2/&g-I
[ca3:UCKa1IP1/Z6f+F?=#dfTJdLFU0Eg836.<ZJMLfUCeJ797Y(0S128V3;c_0&
LBA2_<^V0@6(IZQfZD_CdK,,D;-=c:55NJ[(&YVP&WVPTH=9GZgR&#H+M[J\.BN:
e8<;RW;JX0(?R@&Tc@IVYSg])eKHI/I0<TaWd_McWB59G@4B<@S/_XFKg5VYM<^U
CNJ[KUX92HY]gS/a]<^>P()U2Wf+G7)XBTaLC3DZe6;]A/Z.JCd1ZQTOAZ?-WM7Y
Fdeb2E-E+0#62P7g4^OV#eEZ7E4LD-\Y?5QE?I;cDJ9^XgE6_48G1cb5C(G-&dX#
Sb4+FZF@/BgB3R)F>Me.0X1[?YZOcAZfc+HFQdVG&<]ZTOU#=0f<I+M[.)Ie<1-=
1BgZ2UD(F;63</JVOOd(M=\83;0^f&f-fKF>Y0WV4Y/K9D=7JEI;Nd<daLZ[ZH4K
4&IR(dF0Ig\7aGTZ(5^^dYb\dNMS/<>M7./-cFDWJ:@b.W5V+e1J57IUg22_c_5(
^MNa\.5PBIdZ2A>TY^^6=GC:Y25=D#6:XPPRPe=MYd9Q74NT9(AS-(0&)QR1AV0M
,72>2])?]CYDNbdQdTW.Z+<e;JX2EJ[?:QA#Y=PCI(HLMZYbYF6K#d/V7+-\dLY\
TA<QUYT#9WV^[X#Pa?U<<>@[RL.X#S\/Z+d#B);C+>_Z>N3=2f=ORYJTK=Vb?7PA
V6-[(EVg3.PCd;M-I.A.If[0:UJ:Gf9+++5:H&TTb,BRN/dRK=Seg[ggP-6:/3#F
MMK]-:U46(;RANPe.]V6B<Pf7Q4a\+3=P-@)LJL\^6=>L^P@#-+)H:(JCO;.ZI;-
@YS]9f8ITRZB=V9(,>X.GQgNMDLW#PSGT2<@L+80B92W8R#K1NFK1K/TFI0:.E:N
^aS[BRI#0UNSd9b?9cAW0BSe,5VS[5P.U4-OQ0MF0UC4G4gbTa7@TTB?B7L6&NaA
FC^:b6b-2QJEE<c+gG&SG9:Y=8#3NIKE]4#XHJ;c8/)d\.K\@[gM(DM[HMd4]LCN
-0B)2gaQTHM@VTdQZHX6WE8@=UFP8#a3c8C@e2gABB>e>N+;c#?_a0?(42_]S7+2
M-d@TFE=E6YS#dL,#>0T2R(Ld9E\P)R?1/D,FSdJ<<:Sd\@Dg+&/SG)^IHQW(SEH
LVFd_^E.TG=@UELA2Kf;gW&14DTf+a<)Z^39O&=ISW>[C5AIT5&<X3[ZG1_eS8Oe
?fTE?W:PZe2<Q:(<>&I:4aR-L+4^Ka&6PIB,@A^TN6RYa=?#PFO2H.2ZBcEL;#BW
ZH9;[(I#0eTB#<7:b:_KD@97X11F1Sb(BDCaKa5^.-P-,0Q_be^Ac/#FdQ2YO<@S
C@;aXX86Y=DBf5Ee]_1O)QL?BcCBBQ??Pc].UT.gJ6cL,a@2>-_G43.CU_WRfcUK
PS:;/Je_1D?/-5;O57S/9bX,A]ERYY.3]^dS&)(Nf5^<??dT(YDEXZS/H:.+dX-b
;VWU&2>?&#bIAZ#T^0R9@FOYG7ZHZcZ2OFd,OD.?>ZB7<>E+S-1a[(2I<VJ/S2+U
ZL^aWd9c)KD62-2<c]RGOg+2\^J=4dbY^ZMY-^><2Q\6b3-;E^A_UXZB[aT-T^Eb
d_V&92I=7UBb-8#MM3>S:>[IXMFNROU?[N_L5<;6I[_5\L9RDQF_8Z1X36=VNV2A
;5>32aHGLe1;+C;?#T)EX-#HL5@KWH85=YYdN[X(I)=P[a/R&XF\)La6&UQ5cM]1
G][bQUFc85P<,;#df-<V&NeO[BAgKB246Kac#C-7Q75I;CORb6I&.CX6B@T8M/JQ
)C<RDVLXcFgeLJ<&K./b>&Y7@F,3I.K2BEW^)A9RPaW:P4WWOcT>b9++YXI]@f[a
<5#[S/GWgSK>CV:GYcK?9Sb,RN+#/1C5L^,U+PS9TP^T5I0\cMb>E+OPgT9?-;9L
-b0JUBe(cX\cd\ge1)X1:.-:_[S&5,4eaG.M+SAL]<V7A<\ARSe\f3CO4?6Uc]c/
2L.g-U,+(_:>1;)@+C9Y\K@VC1=gSfZ9D7Z-X;gG:CP?JJ[#X[3FJN.@NbI_#Vd1
gUNX4Gd.TSNOY#.IIK&Q6\d\HPL4eY1]?W;JA7c?QEU&-SN9]NA7FOQ:+L[(;c_Z
0L#EKI2)S]e&N6[8=a-X\<65eAbGE/&9PW=fCgEQ]FM][0A?@6U(e>22VfO>^@<2
A[HW.7=Kc,dWDgQ.U(?)Y3g<1QDcEBZ)8(/1bN0QY&EXE5&a:3f6&3=G<Vb:DcN=
_7SL+#2J?J(HY\MLT^WXPa:80c0L<f#6=EK:@(&<I\08U;Z5.99Z3/ZE?6ca.X:M
TO09P]I\+@7K>E):&eM1Z_01fVGRZ.7@_,@<g)S&YX:[^FUW)I/<O<BW(_1U(g&5
8]+/;.1>2G.A4((<Td>SK)M+gN=@b@OLNcJS6AZIgQC)Y3;XGM.N^2?BD[C>+We#
CPKS^QWVWE<KH_aGSeI23=YCARYV\eLGfW4Nb-1)9HYH08W,N;aJbHSG<.T(O54M
M2_dMa@=JH&U;d(d;-R[_>\F?W,SR)R?.28/9\WTLZ6Q.N/\9>]YcCeQD-Wcg,KM
b4PY](SdHT4?E@YPNR:)D.S>f;<FD<<=bU1>_,)bZFMa>NKW>3b+TZ1cV-fdUPC#
cV.c=;BaAT(S0eG1C(WG2,H6Q&B65H]gPSNJ@?6cM[3P6]2)PT6.T)IL>Vf?#X=W
//T@Md;K]?>]D3UR:f;WLA5EVM.Mbd[QfWbD8VB?-eO:AI-f4)5<XBF+8:18.cHF
+1&L=fbKQC)R.S2R76^YVc140d&_,O0^KU-_.VXE>bN=0P;H&c);\WZ4&/SSf0R-
?Z1\9L8gY-VJ9AXUVVb?8)<^=.69,]Y2:)I^G:B4)LW4[CR+)S2G[=)d<#Z;H]1g
QI]GI^QXMXF,2HX15H-BG9S>X]IO.+-?DKML7F.F^#K-G;DCWV\^JBa\F)dZe2M-
R><2c57<E47d3/:W#F@#C>57We2V)@dZ5XVW2NHXIP,G50&Ye^,@_&[_FH(.+\P0
X;H6@YC)a.FIIT\0cGVQbNQO3=8f3FJ]+8K_ff4T,Wgc.9VB2\[Hb1&V]Og;<8SZ
[)2#BO0/&IX(8?SEDcG0A_MC+BQ8V<D1\]gV.dfN-U8,0?;/RbWUeO0;F0fJ_0=.
DC#+M#IBR5F>\(R1CV:0/&?Q)5]4dV?[CU/Ne;F9MZ45E(/Lg18ONID@(<)aXR#5
^\d3>B2BJfJVP=\-T\2_CZUY8UUg=(XXA,E6_1AU[LHLQ8(cbBa;-G^[/0],adIE
T(IKU(YK:Z.ZOGM9M(&M4_@PH8QeYQ=::^=42);PGc9.4)#0.E+]BfeQ+d0<B,[H
/EY4c?17<-cd.3cHE,e76IAb_46/UPQVT]<_.a-5/cVTT,1QIc9=>6O=:1eAL^+)
W9.(70-:&Ed.C7N4[5[3;fdTR\+0>LF[&>QPMA[.7eVN)7e.19<;da-J3TS(9A+6
Cged8T,HX0J.e6J<TScS@IAdI^11[:^[eF/P6BNg5f=_N\>@7Rc_UQ-W>5=SMRSU
_07[aGE@?P0fS,:=ZG+eY+1#XRb7ZP-CKXD2O2[=(S>RHZEd,U1dRUK2(7b-\/>2
QYQ=Q^SX=DZV59>I;\b&97M(+G0cEDPLWeSbQWO=&URZ)KA>GO8EE7eZeWYN3f0Z
fEWSB16C-^#ObdP8.g+W5.cfBYYJfD@#CP<#9MGGV3KYNDL9c/920\GCD\OeDN-f
<T7I0W,/+)GKRAIWGG+8BTN<?+2C[[@2Wg]OR.OY^PT)H9SB0HD]P8>]&\LHZNG0
H3gEPGU7-KO5HO0_4L5@AY+M6>BKAO^S3Z9NWDc\[N,#NYdUKHUDV)GTdcbW_-U3
GUQ>+NUDG?aUWG94>Tb:eKFI75B3@5:>W>([FKD-:?O1g/(,7^ZfAdca-Gf85HX^
fd1E02-[&23bK?e&#QMdVS7:\>JQ<BUO6#(E?d=;Q)H#RSa[ZHEDgKD<b>S@TQ;8
L26L03AYJ&L]4:eKOaTDO3fgfcST27.e1D0R^BE==Yd47BD^M4MaG]La+aU_)g9<
>\1/MJGN1B,,5[#e[NW3eNF:KT212ZO@+g1&4VGfFEcT:NKB/W>FLYeEd;S1J\PL
Md&WPDD?9;0_JaH3EW<Nf+>5K#3<GKG^D6O+SeQ3_T1(VQK@4)bLS0+XV+Uc=&1V
V/Y@fCA650FEH9:>NG=#?(K1]M/]]^6K\F+SRf8&<IR-g5@ZA@f^2U9KS;L3Uc-:
MF]\H3^aJKeUI77]54fUFV[fc(V1EM7eFeT6Ec8#D6aT8Z1F)Yg=5914&9[/+f0c
a[B5LS]8-bIXH/NR/F39R5(EOAEa,_9gbL:Q.S2P-EbeT(bO:\,5f?KGJX^[;#La
;P0VY60bRG^XEC7&N4R9^AC3=V_+=\ZCKI]O:\K7AU=FJcMCd/=a-[3#eORH\?W8
+Ye=(A;#A29,5G43:;fNAMMbL[+4E9[(1Q.J5P<aC;Y?PXI2^:GLKM#bF;.NM)_1
K54\Qg8&/H2GSFT.#RQZ]e@DA8@cR-fX+bF)5_aKFGKU[3H^^fQBfTU3SB>Z-=af
?c5)XSB,]aX7bGK>b^_0,DK#,@?PT,d\2JEEYKX]S3O;0I5b^(VMZK1e^V?9C30V
4FP//3,.S0N&(52.UfP[CS96EYBFZU5@&S=9g5W.?JPE>D(-MOF&_<E>Q>-;S,.M
-K:d+1SN93CcJg)E>2V:=,Y)U+:/][8ICg5g4D]O]PdX@;SR]M&Y5&>DVX@ZF.=J
>f+:fdaBWe>fBHc7&6-DUR^M()Jf1[d2A?NLQ0&FQ1(ZZf(3XTKY]OZc0G-NEP1c
O>1&]\=<7(@END5_[Jcc+Z7P</8e)DM<W3dDL-LP03BGVODE>ZG0)^-TfQX+JZV/
/L_,[=M0?SK8_<I1X/#-B-\0&C19+<&^(#R?]\ZLWL(PO3JUO\4f4g-ZeZJa3d-X
9S38N@^U\QCUKL(7cSNUG\PU5X])^K9XN^#ZS5+IBO?LO+=a]@,KT(1U__Wf#e;I
<@3#g[.e#cIeJ>Q.F>O@_H/6#,_0Eg+2d[#9\J@\WBC\&QKfM5(A_:CgaG9Xb5G#
TR[G0\R&?I6Gc-MHCS<Jbf(>BK:8DWcf)T]_cSg4ILLVWA5YGN4P):c0S[dHAIO2
NEQ1SeaG48PA\NGS_<QLQ?7LU<3/fGL:Vef)>9=@W]P9.2_a&0B4G7[/7ILA/Zg9
eV.V^9/662JCLf^e5VLCaY0K8=/bHT7Re3>=L0Y5^&_22<(X?DX)&cbS\3HPFe;0
b)IJef#<U3^JJcVB/d5]VENEZYUCZV=VH5OX#LB;>LM>GGB4:@+;\5caM3Bd^;2)
KV@QN=QHZTM?HE1C/G1T:NNGabT2aMM:a-Y2J[dB.]N]Hd7UIa;G4Yc4Icce]/3U
-@@)0AT,J[U+b1V[KBK-Z4bH<WY1J<UZLYP+dH9cP_.]Wba[6<)fBZ=AY3@112@a
]-CUB9c7SZ#\U)>+UFEP@:5<@3I2PdT@<6KT_^+LM,\ZWa>A)AB#ff^IL><\OJLA
cMQ4g+ZDNHWZ92\_+4Fb2D-T4N;<FA-U.@U_QGf;3+J4-UKBK_&-6AdI_TDZ1H.#
7@eZ>8H6N_P]A4LO?;_CA[a:dc0Y)SJ77472bPJSQJMgF:XX\Z5bUF6\89,:2=Q#
D+BO@=ELKG,]XQYN558E]#/+?V,TV=:MY=;gZ],TEH/;MK]00Ec?aR2C,HAG)>IS
AI>cNK=GKZ5Wgc3GZ=(H#d0dXF=dbBLY99B2P1M)#EMDFI3gaJ8:QI=U<^=@E2XF
\^.RU7L4J>=c4N:L#<1DaQYYgR)<eXCSG:=:RT^Z^:(+R3Q3X\2cG)29)Cf.O<TO
[YV2=g3-Pe]Nf&\g#Y=N]#GNaUDF4-dJ&.^)&[@KYA>LJDD6eBdI_gf(A6&HZcOO
Sf;7b1+3X85EfL?J,<<<@>T9R.-OAZ.NWQgCbW]S_<N+UJe7@.9D1R\8DB\<b=@,
eQSeHSM&LC?R_QeMUE9ZE7PQ0dNRW:fcVBB8?<HY+\e4GYJeaU1KSY-T#^d&#6Q#
Q?7#JK]^@:]:4)AF?c6<3L#-,I2/W#2>)]EAHLI_d1K^396IZ<K.[UO.d.;]-AJO
^\ALYVZeJ#=+69,;aDFQAV-gaD^GE^T;M4N=N?+L;L4U2@)2Ge:)FY_FLKJWIgZ:
-KW9T+9JD>FDcaQ=[W-516&O^70T=d;^_#A6#X)P?0Xf^B.+?G\I0@6/K([N25bB
T>ZYS1eaeH.(+9Icg3.c=;0</0<5C>0Tfab\c\D&.Baf:R&R#VR9^^BE2&O=f23#
+66ed7].N7NeM#.eQ78L(b,BF8J^9MZDNNLV/OA-@S:7)BMcU<IHE+YPA,JDcE,]
+d5(C9GJ&L/\ZZD-&S+\&2.eI\M\P-E,\[4f_F5V[6I;f+g?ZPL?XMLK/#gDDGG3
I+MFQ95T\7;R7E\-59RFZ5.e8$
`endprotected

`protected
(GRQ-@;[N<P&O@J<e/0P62J<Y2\H_B/#JS&5^PZ]-TE1@be<[gBa1)/(N860G_>Q
AX<-/G<9X_CbED4KEG@f6&J<8$
`endprotected

//vcs_lic_vip_protect 
  `protected
]fLCOd@5KGPLcW6=QLb-RWA#V6<OBU8U1THbI[?9REUF6d,FSB\Z6(EG[=&@SAXY
AZN;QVBV+=PTWY617Y@1SY&6?W,][fa>TFQe-H-]/-CS.;73;7/8MMJR.68<aJH:
#gaNY<):7NDHG^ZE,=H-=QH?79>#,6[0MZ1>&gcL,J(O[];1J421EXS6:YcXTf^J
;cW#+JY/LKA<&]?9bIa2(Ug4&N0eb0fPLg&#H:TA6HED&Ue]N/3-gZcYCf9,7c]E
X=>e;KgJM^KPaO4ga?6:O;4e/UY(JU05NE>A@1H6Y6SU?e/a([<EY=FgONf[-:Q3
3GP@/=?2]2fW=SJ5J2=Z?d76TaLQ/#FAe;@S](YG6?K#51QV8GJFVb<P(X4K_OeF
B_O)U(CWW<F9T>D>_+J)@7cPJRY3VGP(g>&gJcD<-^>QWS><IZg&;W+8]58SUT6:
dBJe[DD22<\Db\#[X>,K#L)-g8gILU&#bUb5cFR?Q3@Cc:36\?PHRSOS;=QdVEWB
#\,:3+HfP(=@6X77B[eSHWT4[0\FTH=g>6X.S&N<=g@]Q=?1-5/D6E<=\g9^<C\T
K0d,<1YS_]H<-2^D<NTIGNd&g-L+-7N(9_5EZ.B.f._OOW&&-:BSfJ9#<D6-_+Z8
<I(=@.5?P-?SP?O7Ae[TSG71Uf.cAE#S@Y2)bS;@VNdgJ)?+YK&K-^T@TeG01?C]
eC(X;VHc9KVS1PR\)_1;\GM:H#GbN(\?Y-b)9ca7GI)<a.Z)cNA&X^0D]9Y+(0H7
C=^e4Y5+)NW@1WXg>6TL.JUC4K>,gL.X](.b+B-a/C5;SM_V?IN)@8c@]3Q+AR@=
0NTC?Z=838^C]D\Jc4Z7@@]8?P?KVHP2DZC@Y,@&K-I-RId8Q.Z1[KLDY]d.<UR\
@Z,;aV&MGdC:L39cNFg+e)K[=C7Dd7S#H8-=YDU_W_g&3g[HJH1Tb68dIfA-IWW[
<(R#TE1\X@/R\7>WD4UdB\D[SACR=&^F8-)5N?&TA9H]C/(M.:ZKSf),Y-KZQJeC
5T)G.]+\\;K@Q\-_AT8BXG&/&Pc30.B9F41LE=MF#SDK.]aX@(d/#DTZYT^O+7K6
KbYXXXdV;.6bBO#;a6TcGc+)F,S2KSFV,A)PNU>,5[+9dd@#?gFFDO5)9-#RDI.d
8EV43W0)L/#>CE\8?3)TS,b.egZOX\.c81-C#Rg.HTD+S1Vf,E:ET<BeWO,Q?<S#
LZ\449cF3?C[PP#7B=0eC[_1aIE;G?b9_R#?,^L^U;LQ^Uf_baNNUKH3b/^fHF(I
<=WdL3>2WYLD[AYF0.dcPQN]3PW?YI_G#8\e>C;_W5B6df@4g[+89[\48_0_T47-
NAE5/g+Y&_4I0f6c,(gPX-]a_N.GNd&JW:F0RG#B_=L<GdSEJF:^WgR-b]A/gST?
g-R1M\WNePfIP#K;1YA)&B)648Z3eXfJ]CM,=K-<X8>@K<4KIF(./cbK+D8Kc@df
1GZ.X0R8&VZBg>=6N6fGIVZacN5K5e@d17=Vb9WC]O^B,gDYQIKQO5(JHf+3\bTT
LY9E2Ad:;:CT@Q+W#[#+NOfd@+H?eH@0JV_SgOJ4BTJdKI.:XEQ)18=\&AUS/Z@E
UW;41W=\B)e66=X\@<LGReHUc8_I9IcV))P/g=],:10LF8(URPZ4_YXZDN?a#J3^
+DX<]cJXTJcR<J@KO(3P>F]+3@U_ZF@>==U.BL6b>=+CaYU(BM+JJ_1OUNe(^/J+
#O7Pd7ZVN<3RB@F>RgI8193^TQY_<=4\86dRQ8O:)B,\@_U1f;XOAB1cI(IXX547
d9CMaQ^=XKD3+=CB38c,>;U/._.;2b8A/cZ>e]OF3DaF.XcNSW>G;-)Y;5]L+C^;
]#OUaQ?@E:cH@c5X#^MR_V&-1&g2:9e+L+\_@1<A2,8AYH5d]8MQJ.NT;23SH8S:
#;PCa5dD1VTEe^)0#>M(E<SN<9JY_?a>UK1K@6Z>^LQ1:]G-cG6DM1DQTg+[Y+T\
5+D:^+RI/P7gc/cSJ1WZ5/9WIb.eQCKeFO2F/RWFE3:4>LCg.F_4/eWNSU^\FEf4
2\D>GY_;9GWPgecJS]9PP>J1X>+;QbS@II?6J#]&&6/cQgVY\bg.]O_PYPA.V(0=
Pg]b37XDT/-5IY,SDQM[)^ca1S6&KI1M[?EA9XP^E23MG(STCXZYLf=dY_8=fUe_
/PEN>N^2>P0LRKW_T#AMD+1M5A83P=0;;>b]HP?X2+<;)=NaD:TL<KaMP.I@fcS[
6RKAQ0/)c=Z6A@PgM]RU93.6D#dfELEA8Y#_\.#8&Qg5G\LH.Mb/W0GZ(OE=WI_I
&/aOWP#8aK0b,Z.eUaaeL5[[dcL0d<]d=+M0,7:L:a-<I2HdLB:JJI8dW[8cS)]<
MU<>5e>\b06+\]=B_W7B3@NUFP.dCG&YZ5HJ#SH;FcRgG2_D;?V&Q3POW-#;Y>-H
abS(KBQ:X@XK^(gb?;;<YSCaV-VC,e=5U.(?\R+D5<+>4I-P@NIG]ZW9G^g1>5NB
DY^-QJ66>I;6)1GLg#U;;Y4FKZ;(3FHGDBQ=R;D^I;^[6bUad@d+635[gdUQY;cH
>3)9cAY&8&&S3CH;?I.>)\UPH?J=.;65>453X.:9YUAFeB,Q1)2<W)gTUQeN.N\]
e;=Jb?(<5DCESN(G>386Z0aM&L9BJJDD(cB@?R)C6M?TLK;Xa.SO8=5_&K5X(ZB]
;+0gRJIMLLOH8;)\-]D=6#J:OL7#2a+I-bZc(VdNTO3U6E-eUR]]]&0D@V+&KdG,
<LC<MH,+8OV<-=E=Ug4QQ@]X/]Mf@<SB6JWe:VJ[05^\8V@Q9UUP4B#=//N&D@I?
FZ_^TH._F.B,XMU5>+98&7,9&#\gDEGAZQ<g-T(\>:S.g,Zd\SIJMA-e_)HSd_aG
=f]8&;H(E0gX&J@:-5SOWH[[.VUUNC92b-^^]PUVU.?D]D;4TC(7#;:?AOY0]4PC
/HOLU2:4)<Le+//F3;[g[[+VVadSO&Y]<T+Fa>[K_HYQ,,5EB@5PP+TF1_2.6NaA
7)D__L^@C?U5=XQ[NaKa.,[>O&/_PS[9QL@WL@21(P29Q1H_?Z7Q<UE>FY&4Wbd;
cTN]18QEH?)cXc@&L.8)6NJ;7^ASQ:WAER\FX\USB<Z]@,P;CRN9\(3K5/^MdT>N
>9ZVYd-bF<LR:#I7J3^fIAIV<YPQ-ISc,ga_ESbJUM9>cS^9WN9H9BVEb64&HUUS
@JbI>S>5(FZb,9CL?b5aRDbF>GNEg/+)4M(<,GP\;16,[))g+[9Dba_L^VD#\D9(
W[A5eOdF13_Sc<BLWEI)ITc@<PgO,:OA[b0=CJM-(0[N97P@4\g,FSVZ40=,^(SY
I>\c6363C6_;635Q0\>O9L=M_?dSeDcJJ8W?R?,MJGS7ceM<TBaA2dG4E&S+Y>8P
g)RggA]6e#a/E\)G;g;?W4c?,,g,]WE9@0D.P1T2eI[=7J[3eQ8IKL#KT_NBP<fW
=gXR<(5@4DHdX>A^7WE>(BKA3J#ceQ<&TY-Z4-=VE)/G17gQ:3f)PC&]e_f5E^>3
XKX/B/NR9(A.+I#OLQ#g)f?A8XTH>W@5?0SbE#H<Q(I>F84:8g:9GF2V2/N4gCXB
H2/\YZDD_R&#MdN3ANXBg&Y>5fQ(A)^/[6dTDC0@R<,8R2K^SZHI/.M-C2XO0a9E
(P3cae]Y<dGQONK\+)YZ+KH]e5cZ]0UR<#R<:63AHH[;<;OZfN==Y8,cPA6FI,1&
X^W9#beEHDNP>G7SQX+XVeO\2g@F^);54N_EF;7IC6c:cV=Lb+:J67@_Y\1KZORf
<7PHEf[aSJ6&Kc2bg07(7@&.@;>F2X85M98#];EZ<O\&]L-g&@Y\P([CT/aLg\NQ
MEWKQ2;3J.bL4e4)eg(B7RMJ]b;3&GV/K:2RG>\YVVF7LQ?1QdTK47D-aK-J,+YP
,[U+]I/Da9Q7K&c/_K;gY2f/Z_g(C,+LBbD<9SK>&YF-2A&2H3P+W\&;<Ge:B<IK
<e,]DG5UJ)e,\<)O>S/RC8E]^5893.R#7b5)_&2X(M&-gV7fb7V/ag:X;59NY67Z
EBR[F1+FdNJRg&ANB8[cX,IbZM@2IV2XcFL74;bC:9)Q(G6]DG6SabTJ0Nc0BI=J
(V41BK]bfZ,3+<K2^PK6KAKBQ7+X-Y+C--S2L3/<aFJ:WC2JG5b[&O98N5d17F3?
gCeO^Z)-8S,R<A6]0TAY?c<BV>@<-X3CARH)PRN^fJUQB=LSK14QW)?[7,))#b,^
F3LZ@+8B(55fVE8-,R0aR_<6YO>X9CY>D4,2A5S,W\/Ifc0)d,WUfPYVReR3aYVf
,NX=8R?D,,Sf7_3C3X#JNNTgLA,KbEbQ635D,6Ha:1?.0gVI/CNbD.J@9T\+5>(0
OVZ^PZeT,</991&e_KX+O]gaV@]BW17Lac_O+0#2b<cK#KE\_YTdEV?XB]NGO-1>
O:;?Yb89aBSO5YZ5VER(7QdD-6O7[?Y]MBI]^3)/[&)Sf(a7?#,I/]>;PBaM3IDe
6X&&R/WTHQE.f#KIKEQDHN>FVQ9&3>deISBe0QH3YT=R=ce/f5gN#MW?+SBJX23V
VWA0aOET7b),\FLJA^Rg175a)5:6I=V8gPcb+bZ]FISe9e6XVYg8AY4@1ZV5))._
&6dKQZY82a\GK3&2F\_eQ42_NUK\7E#/AfU5N96e/E=HXQ\4cV/2#W4I0#+.PR?_
@c2?>MC#GU;BW4??6)d\PgGd_bdI04J2M=,/gM8([^c2<@CcQO9bKPEY(C&BC.@5
CY)>2-JZ.7N1C.EU>IR\\ROZd8gKAFTX@:475&,af,YV/TT-+)()0_[gbeKJcYdH
Z//.He7M#IHb7X5H#B]VfRR1S&W4B^)@>@A24.LF)OKB-a><g3)ZEKWTBcOJ(QWT
Ic(;f=@O0(9A/e7RZ/(#0&gg8[^XGQ/g\P?QYbY^YVE2<UCM_P^>BcN^GO66LS&Q
D6]2C]KXV[9L:EKBPJ05db8KTfF,FO6H91[[CD(I.S&Pccd&>WeIS5I;,K/4PdQ2
9FCJ(HMQKG/86=5W+YCaZTGAHCM3PW+;HKR\9eHNEBU#Wag]D^F)WI(U_MA4>^K/
XR@fM;>geS\2:RE[COMBe>VRL;8g(WQ0S2Mc(/^X6@1A[V=&09/;YdgHVcN8ZUDf
&R=YNUGagIE84&L:0\9,]\>@I4WG(7[076J/XU0BNE0_S3X5g[AFJf:db/W1.T.K
e,Z2_-D)b5gH&;IZ&W+B4Id>99E;g=(&=.e1IFE;P[/A\VBP(3AYOcf0Xc?3W<=5
b?f?]f_LTAKD,:WUW^FgQ/X44BXXaFKRB6gJBU9&]KCTa\7G>f[C(G16;XE9#=16
T3>J8:&UANFSa5=)D447LD(YKJ=8WbHP7@f]0/a-)H,,E]F-,@QH8W?/2L,<WX]1
g99QIMSZ0Y.FYXS4#\+8+)/R-@X40967A?4NG_.JE,)H_b^<CJ14KedQ:8^@&PLf
PWN(gfD4<.@f-IZc6I,>eH#DS4E.:cbR<:=-2X82;VA<Fb/XX:6-a?:Y=+.3e\LC
O0H-?aO,/-/aYE[]J]=c/9P-WB>cdd34;R5D4;bT^;&0[9KJMATH?K,Z5.YA@)>-
d<I4/XEDIQ6c6-99GXU]QQW[\7c@\69d;3E_fP]bdRbf/HXbTR=c-K15A&DD^MP(
cB)8,#d#]:75DXL.AcVA]PU1F?6C]c=L_<D2Ee@_C1^f4MS<,(2C@bD4bJXY;HUc
@(0_W\AWcbS6L&+HBGf1a9bH[[XJ^IWP#PVSO?,Ra>C:[=)<F#1^&MI8:9T:MB9)
4HD5F];)8CQd?eA#7Zb^D)cB>&&Y5=@9f#\#8^19]KBU+(L=P7g/G/QNO):2?/+7
[OFX=KEgS7eG\PU@(/(HIC&Hd[D9EP5?LG4JJ)5:=_VaeNRfX(J:Nc^4XRZXPUU;
^P#BC@g09FCdS/;OU\gHYHf^LDd(X1+[&=?.ZK=<+)45@CC+g\RQYaJD_]R]W3UA
K.g4/6>76YfbZ2gR#=Ef78TB[Sae-=HP/fW]]?CI?/LF5S+cAK_?>=XSHAa@S<d(
]BZMd0UC)4BQB/3T/TPUPabC8RKN7b_eVcDH_@=bU(]e)FHG7Wc:F[Q#A\,CVU=7
2d3>5aX5><Wfa[^0PKSUB]-7,9>2VfF1=#-e2=J4^)<?(U+:edLCE>RSIVW8LMCN
Cf[4Ze)1JA9ffCX].R;W:M0VcXV_T/Y[>UZ^02J9Nd(PGN;8IQZ\CCZXe5EMU++(
L.A25JKB2^1fFd38eII>R\?J1DJ8G-DD<?K=X<<\?_4&e42#B=c]g.2>51@W\#KI
L@If(/Q]dT_K[\;d]9N3#;O,\ZPc@TLI/Q3USAGYg+75GHTZ2A@1X-]W11]U+=N5
=d2;\[10^B/ZFUEM16OXeA<-9I^=LO[/0e3H3d.]Z4YWgK3Q4U,fN\8eS&8R0^Dc
J6PK+I1MaRP^gg\658/0MN>+\5SF=Y;eLGc__(<7fN0eG8950E]LJ:J(COZT;N0]
T=H=8bZ9f_6C)B@M.f3=9P/Fe=#7=:cSX<8EaVO5@6W6T41g6?e:0K<FafGAVB2_
)cCTcGU[5PXBaLSHJW/<:e5TDI^;+)7+2Ea6,QTUR\)5\-5HQ1Xf(ON=7+N-&bUc
Ie1[6T]eSbJW0J,>OYBcV4L<-f+70KN6FL0<=;#e286-+G?f2Gg&CDb07[:JKR.^
OgANXUZDf2g:M]@..COX?a.4eXA]MEOe2^4GJ#=LKQW/3L9<HGPTCWdTgLTN/M/V
aU>,=:UFO#43CR@SIg+7:P<;f)[-Z5\-BC,G(7)cME4aH4?I8,Z^704e_2]\fT.J
5f.=^3.DPI9>F0BQ)b4-F^H[IARecRER38#/&=#EZFRUK#-/0Z4YfU\UDF&R=G>4
OGgg>]&JMNZ\cF,()JDBH1S:?eMVMPUUI_&,GE\9M2:YGAEF+&)V,.[SICSDQH1=
D6FM1],SWXXA#/AJV+@<R14QaT\^YO5(1(.A7M\eV4W0)WPXJ->WQfJM=Uc4,])F
G3^M\+>T>XG/@KA#;RG[DJ<5D;I,N<2#W>;8E#4F\LPWVZKBgK2N3Jg^:;K)AR=C
@FQK+<>RIXK^Fb7KSIE\M+6:e8=E8><?#N:g_;<O&V?D3DLJ&2c#143H9G\-:;2.
eJ4E]4.B,5X-1Z0Fgg\=Y&d>6^I>]4)H#^PP_46=Kgb5VA_9]O,.IA?8RXb#1&80
3JF59RL_8@\J6=WY#C]L&-9JOc=U?Q@?Ygc#S#[R6,J3;XBHB<e5Mf-JP4#fJAGI
egbZZ3X@Pe8=M7e@HO@FgP;UP&L_,9-TcM&b6#C8EM^^(b.YZbFc>@ENL3T-FC#Z
PU.87LSG@?&A8)^NSNP2&.:eBe1-YR+7=UI_IKU7=UPH,-L4JXA72X+B?f7MO_2g
_SJQ/C/D:7dMNa-_50g=(9=59B@QL4]DUaM[ME:aXQR5ab<C]+Af>_bBZZPPb+JG
C6:4GV:O\X+YeZaeT5K<3Ag,Q]EYAEJX_0I)b[Tcg06Qf4&:/RdUb.8eAYE,S4XB
^g@a,+P9M40bA-VN/;a^,SBA.[F:b-X;e(8A5CG@<X5CXdP#GZU[VZ@IVZbI^b9Z
X0f>]f@:>IOXd&=ca0;N6P=GL:XB5a#8]L/SPSNA]fUGf=bHV_98MIf,FSg&_6+T
_5e2<\^JL6bI(\M?K-.(Ca,SdC.<W@Bd[M(NY(N;D)8=-+YSC5,IVFFI45U]]7C>
/KX@FW[L+.9H6-AZQDF0U&,84X+OT/=ScfSB4HA,R/L?<4/5S4+/PT>D9-=GM,c+
CK_@bGAOL_\HE[>,&bN12Bb.)+eRW7:Q<BBY3g0b9^=DN)B:@[d)QOQ09ITCbJ1^
Q_,L_?>_&cKR0PCCB0D<]Z/8D/75IVR_;=5R_=5U.74_^)W96@P/@X2Nef.MR#74
=P&FU>71PL01LR9dcb3<0Q_d+U&5(J<+XDZ>LFb_ceM6FZ:RF,g1c#4JBAM,8aZ+
/[aIXHT]=WWR=<\?C3bd0eB35^P7AD0fd6CK7[Od2Ja9<eF?f[LLb]U4BbXgZRU)
MHEQSN&YU75fFE,5+UBU1MKAO^W5A]P)F]Ed-^cI.]b+.G-c\c?;5>7?HZOI0[B6
XXF5/&5BJC--K;)eN2?^:EXD,O:;=H:9JGd23d<+]07><IX#OEU9JSY=)?e:3<gL
6,E_dMM-:@1@QCT=WY)Z,(W[0<F<UAH..f4>8HX7g_bG7FUGX-/D\GC#fg4P0\T5
NAY)_TD@/A:[,\YVT62HT3)F)=1A)bFIAJ6CX;BW?c/PaL.?:H2VI_VGU\C@TV^+
M;F:&=R\-V3/L@ca@T#G>TS@/2,8,AN;=G\Y<V3\O4DG;3D0ZH[ZMW9U&<P>:_I#
1g,,(DFKS<E7RbPR\S^S+U6gCD]4E3LZYU(gIU?35T#H@]SOZ_LR5DU&O_a7TR+@
d5U.c3_?Ab_MSdV[G4(+QI?A>6=>[;MO]e,:>E8#-E2e1>);UDDL26gI[8.+K#/1
GL@)9Q6e\a:I#.UA&>:3=Z[(^,AMG?f]2N?,)@H]<2&V#,F4A_0;V->=caRSNf12
ZY<E.WcU0N.A&UER@R#4I\EL>7A5_#>F0^eN3I4eK4NC@2fKA?8KRD]MQY@G&C/b
YA.9d>_:JY6=,6Ag>dBWNASe+bYF1.2C2YAa)()(//+-,M.)_]4ROe]Y=2AEA\,B
-JV2Zb;4(Q<Kb@UH:?GeHFCEb,<LEH<Cd78ID+<:BYH#P^S/f36eH[B.+#=.\XEO
=,O.d1+.8WX,#.J#6H1MT8FP9J,+K:SV1IZF9ZZ+VSQHc&_Z^/S/2A4eK75V7D1,
f2P.97\DP_R,>M.ddeU:G6I<F,U2ELA&;A.1:WaN==DT.OO]HAXFODWO+US0F);T
XV9?F(6.)Abc\9MH&dfM+AZRKJ7bL:gK++CAE\Ya#FbaXaJ.AF9ECV72GgZH_6gH
/Q.fLUITFL&J96DVT_e+YK?6RgDUaT9Jge&Mf7SKWX<)#;N)0Q_V:4SV^gC(XWD>
[XfXbI/YTd,?3<P(a)OZPQU(g<L]:.]:/.KdNVa/-?E58UeGIXaI3dCYI<Zg:CW/
95[UT?b[&dK8YE7R5\_eH8ZG5;Q:KR)KF4=MXY=;#Z8?T4V?f0XYPH<27(/RfEQ8
F4.V/_/@_=)=^YP+#;^+RMX9+FbP5RDfE54[#V6/1,7\NT&>#&\X8BAV6YX](a/8
W5:MYfP>IHDgV#ZZU<>]=?9HgUdFI9c)f>N+BbCbX6ML^7B8Qdg5-1O<SLYU6)F0
G-RIUT6L<#P2e(0dX_.cC2)Ne[#4f&:^EJdD38;P-R+GUadIRKX)][VJX1PT_f2J
)ZP0\GTMF=?YG6A=,/=9=>e:OaHY_VI2gd;c3]#+2F>aQT\G?G)>)f>FfG-7H=<X
(?@;N\MAf\X)[b/SK^b((C=]V6YD>UZ&#LTTZV1F^F)MTdgMagcdE.678>d_G\P;
XR<A?ITWPb4\L>AZTD@#\.^>bCN:)Pd8bTg<]J8O2-8f;BZMTROF)\<fG?9)O7C=
5=93H/==#0Fd1b0dV(W/_R/UeeF(bg^d?<8C,AEIES1.HI(QT0<+90_B1dd:4ENF
74#-+(Q4>:L]<;8_^3TJ_36_fRW1[X4RDT2MaSUdgb)P;\<J#NJBD494F43>&P3a
?&Q@Z]WPe\>6KQ,@QI(&JG2L4@Da9SR+IBB[E1;d9=]9X_/B7cUPbN_OB5_K?<>-
Bf[BU43eT.)OO7Pa8gXE?MA?=70NZ2YIB5aG7J6O,LQ>Vc+:9fc7AAU2_&58DT1B
+A8aY[aFT])O,$
`endprotected
            
`protected
&Zg?+4X=152]HH24:XOUdIGa\3cP^Db,fc7.><Q]D-.1TY8>B?@.-)#ddFPJN31(
4dCbHMR>@)##R0VaeN=<aC67(,T8\?PFb\U<7N##LZ=(/BQCO4f,eU:>FJcB-7D(S$
`endprotected

//vcs_lic_vip_protect 
  `protected
WH<ba?gEaAR+:\gS+Q,M0D5@M#TX)SgP+OE7X/P@c/<\0c_L=-;e)(^-UMF072a=
YI_G[V(B#Z6_=M@g2.dR67Q5cBY#4N2S)NB1Q&DB6@e+7\+#A)B2d3<5.cK7#gMW
7I;,0(3[Yd:@#b<-(^RPCCYgC_OV5f93f=HY\a:)g^5KQ=&X3YgJ>E_g29#8>K&8
GN2MMCd1W90b+I7LgAa0:dN#(^SU4W:X@=Eb4C#>I/1@K;??>>>?H-KQb;S)9ae@
dNN^=Y7J2.(Y+B;gYRd0@e?+5FfRQ@LdC</_F7R06?9E[==g,J1_0M8PQ^;.W8f6
0JZ;5[[gg/>T3<=-1L6H-\SMP?VVV5^6M6RR.&26X1)gBVa3Q.BKIOKWZ6KQ&NS3
c[c6;RD,bfSBTM-Q:B9I_d=8C7+T(#RPHF(^AGXeUK=UTL@&g7#ZR5D@:VD<F\aE
^8>43FUcU]+M/A]TM;1e)\FNK(TadX_.^-,dW9X+1G9C/USB/7=Q1Dg/2,g-Q^8D
LV\\gK3VgL]91A@L+U>aTS&b_[H<B+OgG#g-b/e-_=Q6#-M+.FFLFT\6)HD5Hg^E
.5(bHS4X7QMe;;f(CcTN&W4e7;#>0\0+/W[K--7?<Q)^DO(9g6?[OHdc:7JeNG4S
7#/^M/a&Z<55QN+9/=^cX?SX6cce-56)EgI1a8D9#S/B&+@O?5\)::]Db[^IZTe8
e27T<#B(eE+b&a#2fE)_MW6Y5G\.^>11a5,@OI^+@RI+,&WOA^7K:-MM@+M<;F6U
-b7fFS-[H6?D(DO[N+7A<8D;7,GORXMCeNNW:,Va=&@Y54UaP3C7OJbE;ORVI);-
bW]B\Q_>JX?4a)6ZHMRgYJMBFc7L&Wbe0.Md8+F1ARc,8@-B,^cR8;N]9E=13T_X
@,2dF>D@9.&.LO6Yd@HP.g/M0Ae:Ue8JC_2../CJXXce[IP52)C2fQQPUCT0?>]F
>E9/39J\U&)gB.YV2XVObS0M.;aW9ddI6,e=N#0g:>5;=^AdTL=Hd;>F9N)IQ-TC
,.0^MH8P2GCa;begOGU]7KMb;)7YeMNIcC_8B@Z^B0<Xf=YGdL9ULYF1Z)fZ8VFO
7=fb>K37b\O.gZ#[A+NM6Hfe_-)=H1Bc.KM,B:EeD0&OK9>@ENC5Vd)M[;/?L^^S
2+U([[-H.JZS1;5/&N;2^#CVP+SLQP1d3J78gKG02UGX9_A3HX.5f,7/A4=@Ke5Z
e0](IA?S&5SF/_bMe?A8O_[P?<f;eJA;Y;+.8g;#V_U_18I<+Pb^21#MBGX9eR#e
YK<a[Pae-6._SZUR7E-Q\dEUGd.2\\5d7OFeFKEB2N[GTc,\_Q(@^LD]HT,deH0b
SES>QV3PLE:X/TODK\EAdK=[eKNB96a&\_-1(KbK&Xgg=3f6>F(XRTYCPI9d/#3Q
@UO,.1J<QCX^b:DHC)C:ODdf0HT(,Pe&8(C6cdV[83&?b^=\VP7QfbRb:SW_OLgd
UT_KM2[)JIYO\1:]@TcgCfC#,J_<J0g]b[G.-:+M3aI1-W(.98@2[e\A4cJ_H(7N
E:;5+70<V51/>ZaBQ(QQfC=f\D7NAcH\B8;,R29RNYXgO=(PKdD025<b/QW?3,9b
AfSIW4Fc51Lc?K1Z6cLC[>F/\@fTNJD?T:=40;2FXXeA&B@C\Kaac(GG-a6M-a\0
,JQHI72MCUb&7:9N\=_4ca\=.\V;X7E6&PC/5e([R)fMT9^W:^^9P?OB-W7?\8?F
UI;PK?&Y8>12ea5cd)0[/4=HBH<O@a.&Uag9.:EBc,=2G+XT:6+/T853YLRReOeT
V>M\XFcZ\[Dg=7a8[Q1d3N:G8\2?W45gV,7P=OJ@7F5PPZ]NZ9\1(O97Zd-HG\Vc
&L[,>F<>@-cNK3a.EXUJ?HJe1Q9-#,+,+P](W5feA:H??4(8M7V:OZ58MJE^__05
<VONbHQIST\3\Z7e=V7BL\LB/6cY5c\B6(b#C([^>P2;f.6J.G5dd]?;:)UKLQ1L
AfH2T4#fC=cd2BAEYUN#cOefWJfcI.?3/\7f8efHB5,VedS+^U0-V^\X:>=6\_9@
>\GFR\7L\3V^3#I877<1R78fUTFL/LU3F,I7N#1cAKZfEQR:\2K0_C)WMP-80Mc]
-9\SK;<+8c:edd_PKaKA)-[W6#-A4?b6bE]SB+LE>6\GP60IJ4<]6FP,>SA^OZ3K
C^DQ,@E(LBg128</fb,7]M.Xg869=eK^,EKZ3CM2GEOfN1,P;+9T-NJ4E<;9(QLU
+W3A0I<D?[#95B=fG0/[5<#<CcS^J/gCR69R.^[C(MJf7f+[ffHS@4@_>/<_[UU8
>Vc<LN38G\N(K\?DD5QQJ5ISdcNMf\0Y(bWWXDMH)RXab+E&cX<_b#M27@a(SI0)
UfFfP#bcHLRW]R-:?:aCP@552c=,aDVgW(ggK=8aK.f(d:ZW[YLT=+^_Ve+.EBG3
O-5Y3E<EeNK<BbM26A(R[^Da]+.eHOW).US:BWV<De7JRH:&,3PVb0FUHL=\H0RP
L\@b0@4U4XW1f,E^R997&Q:&7Z@7XB//?@g:@_ZFVg=,(ECXAS)a+OaG)5T3>V\T
NT@N@KTUFdO90S&]2#NMRK@W2L.&Y4AQ:>-(L+[f)_06f<-0Q71,T(+&S39@8@gH
608G12P?6(@;3EV[-QT>9<1R5VG):c@+UD)2bdGQWL7\>KD,CM_Hc.+?g(F;fI5;
JB\AU.CKS?8K.QRGE\&cIR#.X>3/dec,CES9/[]BIg<g^81PKa&E2;.&.c_H##c;
1BQI1+5@cVfX1<3>Hf@YD2AD4QgKE;57b2FfPcXZd3EU6.74Q>5P+C:]N)K0FUZ6
F_IXD63A.W15GZPO=VF]f,MD..;;L\0:a0L]LE00IQT[]0BVI+>.2L?,&aY43^^:
Z<S.44,3Jfbe34(2WVAc<=?3C&_AA\1/?I\9F\E_0eGB/=95VMb+#^152D9EEB7:
3PVC5COZb3LFJRI&=QP4#-dUgK-:9ON\PB&V.0/8b&Z(_PMb0DG7\b8:T?KORDO-
>49-#-MH]?8A?LA=._LB>7@+9?YBOCf\ZHHS0aO&+/MB=BCIT^,-SF74E@\:U_ec
O(YPXBD0_QKFDg]?0gJYM<FR:fd5QK-#8UNQ\b.7T>cf9a+@<2<BXP+&>MZ)L]7K
/E)=I,8AXD+/^+4E_[#RPBBZ745[?E)SgB;,G<RF2ZCg3.[&C-Fg;eLdaN;1<L.Y
Y]69e5&g^?[435GMfFg1Q>XF/,6?/LZTXOeTaW1+0NdFec)W#IM+dMLPBK9&XCM+
Y>@^#.+ge>,4Eg?a5@RFYH/57:91,.(>,Sf7WPeQ+#4P\7^?E9SHX[A4[4ZE>7-M
Z^=3WJ&VCPF7LN)Z=_Y]b5Z0;d_5];6Id;O_@QA-f0;U<T\K7@;RWN<DEJ;f0SR^
B#6PS@-5G/BNC\6LIJ3P)H<H])dG-g=_Y./0@3DG?EJ/c./BI>D^cbcP3TS^D:@[
K)7.OUW):<[_^U:/&AS)ZFAOX7&?AP@16d[fb7CV@RT5?-Z+Q+2(9<\T]-gQ?TO]
;MY:6[O0S>cI+S72S(QQ;E-L44T@8gD/^c3.O\&d5/M8H6)[ZG1AKf&a8#.:9&<e
5CT]5L_\WdX3c+6II)5^1_M81.5K14J2ZO;VY?X&IA,Z4MWb6>S62:WI53?WHCcb
5I2F&E?/?<[4M6ESO\fE\-SdF=(.UV#MMU&BL#6WEER8D\/4ZF-c\WPPVCZ>ceH7
IB)/5OZR2U(@9MEV&U:gdGO-;AN:DD=?MDb9@>[X+Z3/Z4^<IJGV(C5QMf33>K,F
LYcd>RODNJT/MD@O;c7]<P?<O[UbeJ#6PZL/44J^Y[-#EMCMg=T_:-b5P4TLANZ-
MLDYPS?;.B:fL8<E;3H^YcR_db0(O>^/)_\<A<8-I,eZ3K2TFSH6SdUcE2e#Qa1;
e55CJ=/NY=R:;P9PW?2Y\]VTeN^SDbE+?f.U/CI(0((9aC]dNZG.G-.G)/++RF],
525(KQF(FUS+\8@FB11;A]/,?3)aab>Z1#=&Q.WXeS)K;6#6aP=JJD\aN;.3:UKg
7K@Kd=\9c-0NT[O)2R.H2@=?NS__(a2B66;_,3g7B^)V?eI+f&^[4&=([F#-RBdY
W[)PM[KRSa62?)_6BLPA=F^O3:&Vd3D/2g=fDCZbZ\^R7eO#f]KQVB57ZTNN[W9T
7&]DJM]bC+\=\:5dPNf5^<F.ODY5SN7LJ9I2Lb>1XgVfa=1fg7c<Y]Y<#)3cH^M)
IC)FUGDKXUT&MH>TgQP)T.EZa^)aK.eMV15/WJKfXYGPTS2KJ^CbA6.KH/;C]PV]
EGDgSD(T-Y#H+?=#&:3:_#/P_Ff=D)II=L0;GPO9?_(SH?ac#@L@_IHBc=PGD:Y+
Y6--,N8Zc?X742+Xe4]FK;cVLI\66;4<&3ba3/#cZ1NND?<deUGg:(M#d6a/PS[(
U2.R_QCdK9aV<//#&48^<Gb03UBL+0YDE(4ZC[[M.7d;WfM3N>aCB2a&JFEcEH;@
@I-<+-f+EN4-Q[9dX0aGI8<O^O3LQ.P.bXWLX2.gEEKE,IYa4(UGMF9._//KVb3/
A<2cNWW6YJ4,Uc<.3P>5S3?YCCfFQXP6]:ANf>SF\^723,Z=CA]4EHa1&)L6N&5e
6H\Z?;B8JDVg2g.e\?+=6Q+262(L^T9YMVCVXUfB@,eQDDS?M3QV[ZKSJ=+7gLHH
&0/NA7V&LD9f>a0BI6MZTfV>YU.:e[91]b_b27C)bSaF,V?8@9+9U\J/6R/4U=#D
L;_;L70/B;BZ>T)aWH50YcYe/K:S6KG>0;^R-0YZ,<)]G;fP&De6J4)]QU31&3NJ
SFO_[G43g,ULQ.+8C+aC?RgGFHVf-<F/Z+3SQ/f4d@J^e/G&>7R4eN6^;WCW\\XP
#WAWHT=SUA:ADTR?+@FR]^4?8OYG)bA;6HR9;<=F9GJ5FC9a?KBg670GO7UN-YIS
TI)/Of]U\66Z(AUd-V[1>DE/P=RUOQ7D.bE<97VM4O[^YfWg>V).g<A_Z(8<-KHV
2be&A,5g5\QTN8M2<cT#7)SQN8,8)KFNHI(9T0LOeF@DGP.b62_,EU3?f)WDH[S&
?(JOAKRLRQ:L(O;F\:M(PZV8<V7:M>J;DU426(DUG;..Jb>R1N:W3SZ>eJRGI#Ab
Z:&E.U7[5.S],.L=eBgcb5MUdBW-c0?.HM.?>?C]VS4H#H_R>CDeSJ#&H5bR&3ZP
9b9YRD(Z6I)[F9O2X6KGPC/aQ()-KR&-TF/@f>1=f>^>6\9Z#eBC[.9YOI)JJA?1
AMfA65e6FW3U9CWQ(O[0e5@/A8CBYN+95bGQ#FKVT5Xb_EKST;GIPDYSX3?9?#\b
E8W[LcERBB]KHX^7ST:=TL/e)L4e7<QEHS.d4Ue8<,0_bMcW^d(KJ)<H[Z\4;(EG
LFO.dR\U.R/&JTN,\:C@P6BBb.;6=7MMC^F+Z^-,92CR2PU)\G3.-e9R7U/5cLeU
?ZBE=,3HSTG]Y5Y84aA^LHa-P0N6/_5O,PELdG&B#WKF<)SIWRLYK6\8?.Lg=55_
gZK)a/CL>^)-2#^J_ed(CER[HSMgVQTgI#0J0B(;)+T3[H5U9K21Gc&2J4&Y]aIZ
+W#4T?X7:4;a=L#L[CKYS>@B8Z7MaX]Eac_)fBC_&5&MIb,-UW0V0ME8e#)RAM_5
;Le@>J+5J@d+fD[^=,dU(EV\<L8b#[)N5YfE<06_;Z-Q3BJM6L8\-Sc\98G31J)^
14<(2Af\P#c?#faKA_R[f2Rg7X-;:R4#Dbe.Tg0/Pf+\V=[DBI3[EH\8_RLL:a=#
&X?a]]=CH0J&AZ.dXA63(F4JO(f0&ZBJ-K.=P,@TR0f1g7OJI)4=?\4I.9DL(gg9
eaXC6?a+e(=f##+@J)f+#G.\BV>?)<3HcEcb7-N\H>TXY>8C#91JPO&;9:1GX6IB
bdD&]5PHI:@:K+DC^OQ3\(UP+&0A5YUZ[R>YegE[[J&NR9J9ZUO>+KW8=b4Q_O\F
9/F:4QdFL(;Z4ST,=DYZb.91UTA?g]]&S],PJ8ELf^^W1NBc.X>SO5<A.8?fZQE9
W:F4-#5ZbPdeA#8OKTL0<Y]OC^Q>76@bP+fgQPbe7b?UCTf?e4M\]IIgW+)&OFf>
RXQa1TTYY>>,@S17f)J;e8P.R<P?FY1+](aKAR5\e3,6S22-,J)Pf2#ZX=Jb@E>3
HVT6)N==QgM=^:/(0[U_=a^PNQ1U2CVa9ULK-_34:&OC^,@,D466+PD(bJ>OO[_S
G\;,NF-9T6ff/1WBR;C9()F9HAAG5=.[L-]FJ/ST2#U@=#_2^.VT_B+1=_2+S3)W
;7;CHYI#A>6bD[7Ka>f2ANGbXBR3FUP;AG90)PJ1?G[;/X>;6^(?++@NS<X_fAZU
4Jd89^/=Eb[BULa<NNC-;KfJ/-ODHA_WbR6-.>K_PBRJ&XJ\S\QKUZ,SYT5b[U[C
1eZ/\2&#Q(?62Z151dY&HaLRS5:O8T_5@-W3OME1)0)UL&\@/E40:c5V;:aLW1VG
,/e#6fU/05?b4DfN8cYc2=8fgA5#OI5/M0;;S35aB=9MNULQaJdM_FH.X-eN4/[1
bL(H8,2(E1a6L1]b7XG9gV\L)VA@Ib;;dFE)LVOSK(98W3R0f-XH=Y:D@aAMJN5&
MOEL_BBRGLbOK[eX-V_T0b[\2E^g2Q(/cd^8,+?EA),gUCCO/R^+=D,F6OEg0&dZ
F+(4U=QU2dbAGQZ\B2YbAab#-;eR+.b3O5^F73_GN+Ng\8W+U?MR#_^A8E#+WN.@
G&>Z6(F:W3-&HBd)c[MeDaf&\;efW+0JABMA(77ARIF6Zd/&EB_SNV-.>&F:]E?H
ASAg)KQN?4,7b]e)X96M9\IAU:aFLSZ?N?@GKEU@QXcZ5-(?[UU<XUN--<Ic&OR6
7cgIG?+_79e59W[dE5/@LF;CS_N<e3\T#2HZc@(NR?@<aYG&O^Q38dBGQKG;L<EF
=<BNG<:^L]DeU;2GTS:5dV?)@,_45Q^]^a0-E(:7I):_gSKgZ?IM[MWU,3L\<KE\
:b=/FKC^CS;:;=.A-U8@XZHC;S<)KA9I+]P4VE7RM6)C,5f=6TE&-e>]>&Tb]6;)
0YPfeX2.WLLK+1?HQ=]/5WMdJ900g83@4+bA47;&^7aLSPEMMMWMQ9I2e>,SH@=U
5Zf\)4AS##B@&DQW-D(Qg4/K)_0H++0:TeY1gAQNd?60D;18C<Md/9(HTP4]^KgW
?O>J(IM;;P1&<K(F2R=+OX6bZeO47U5W5GF?84TRX2K74F-P;MdVT+RM.+AB63G5
=?OF(R,)@I/E]Sf+;+DW^5,f8BWFf:1D\eQgC+TEQ-?F)SfZCJP]c&XDIX],Me_f
22V7Nd4J+J5ZISGg#1f-(dVH3+,G/:cMAFB>cP4=;[Z\f:YX.]@-e(IXb2>R<[f(
K;[Q=I(eX(7?]^)F<af.I^1CBX]./Jc4KT<Kg-b;7XJAd\^_1N3F9;9FQNSABTU;
0O[X(O09dLcPEZEDX7KKUW/4YBU9NJO#:b:SQf0X[1g];LT(H>XPRS09_/La?&SL
a^Z60-)U\-b0]6^+F4@=/19FN6)2?211e>];^c+,L;+UER5Bfd;Ed02MFJ([SI)K
CBAZ-QF-R\Z&,Xb0c;HIB8O9/\e)C&b4(_cLcZ@QDFJ]HfcJWZcLPL4+H3&CB^AO
?+WR\#=A;<57OG<?f&P3WJS\ENI-;UdBD]_](H.IXY^F?T=g3d]45g3-8LFG8I3A
.9AVIPN(c5-X4Q:.DGZ1FGE>OBF<XYH[WRJ\KAaKLN_bf#@9Aeg0]dG[;308U<b7
,>/O(W>?Y:[+23RY7F.gd&Y147HG@5)9Z(6DVF@HYD_490-2TbKUEf4QYZV,#D80
/RL09=?F.4@:EGegBa/^;5JK30=WWbWMa\:UTC./NP?1bM]/.EO3eUNO:0,LX<>,
]V0,\UUdf,d\3^/M<]LH8GcZ?9U\ZSLMT#?eT9Qad5&-B1-GIT<U0F,=1KWCb[=/
72YTUH;2J1f&RAaKPWIa@TK=JNcZ\HPcHV#6\\_JdJWM_I4;R>WWI3NbR+J5&aQR
09YN?-V<9:.f.O4FR7Pa^&YFc^P;d34b\OLWgORe8J\<5X]:EC^(N52/=c1?EgfI
WDK7NXW3cV=LdS/OJ-fV?JMAf\G4UMI41OLMI5cUa+#-J5=ITWYO3gX4BNR2BF[4
B812:\MDMEFA\HL=XE:Z)MVBW>YHXA(dUUTQHcAF3Vc0[cGF<Y_8.[]STX1aG4OQ
CAL6f1^V(:06;MC>^6Ig5-BbHAI9+5bI=-#)+0M,42c()Yb45XW<;LRM6M=f37-e
R;,NL^&EA+A\:D/2J7#<AOSZ.E#M@H_O#?3d]=dZ,YJbaIgUYd\]<;\>gK)X4J=/
8>(8a[LMM1;Q;=.V\)WN@^Rf<aCF/=<W[TDFMK]bE#I0fX4ES-WA_:BFfCa=RQ;\
\[BI@4VdcF8Wg88[O&5VB@MI0=FKEQGER<&5@7]1MGCW>3E\X)YdI-Q/]gcfQced
>7.(\f^b0[X2CE_K-ITXHH@fZH^>:^&6]?AP4./_0D,+\HXH4X+67+,)LNb^KWWZ
U=eWK?CaQf95a4-\bVEgHag[W:=7QR(T^Yd6f]F:G)4,25O.]:)OcNceXG4Z]]8_
^EU,@O=OW8(XUTaF4R)[K7C&LZWRCD=H2./OG/1J#1e+&9:Qg<PVf3e7BW?3fB<=
Z^\_1c+Zd+HD.<5O?,J#g8KIa31<<a8V\Z0#aBGGaI2=;efU\;#JW?LT=:&4:EDI
b,]\\><5@,52[\&g2Z3AS]:7fHM)H-SS6PVW3=H\DB=];N)C83J&X\##E,gTgJ@.
YK.IX,NUO\_(]6+#<d8_<XL0b:X&ATTIdL]NQLIHMN_(0C20I244=T2F[SIEH2R/
JDHH013.dT_Fag,D)8RE4GbDUb0=NS7>,/C,Zg/L9:8+2);SPf6<-^M3@34CZ]5+
GQ0A3OSP//0Q@?e7CT22H-dJX-ACE]4f.^QP]0;]-FA7GB2aE=A&>,5e5PTCL[E)
FUWP:A_D?#J)?b;M3].(-XM(FG>VZOT#L=c-eZ&/DQ.6XZ6H?.CY)(>/&bGXK2a^
+&ZKF)<Y1Z5^>PX0dA]<&T2&<=3P0L>73/a_BH1GNc)H12Db-Kg,-AO]<O+.cd_U
[8V)PHO[ML_UJU4:88,&D_](,]A3^IW._6:;86<7+4L67^dLPL\9KP+:FY-Uf.@=
J7=4MH/Ed\ga>L3I/]SV7\9JQ&(g[dG^6c(^ZO11#SPe[KGRCY#T^O2P2D&2aQa/
?[5b)d)]g=:2QB2&TF]B^J]C+U_?X6TZcOPLV4U?AeDJ@?/E?02,9f?,)<7=:UZK
daNK20a3Ug]<VCO_XIdAR)Y?aF+>+J0WU00\/dN?;/7Z2:[19H6PfZ9RXOdWJOB]
Z(RR;7(UOF0)Q2AA))MX1><]L/a-,)fPV56:Dg[?1CMT<@((P+\>>7L=4H_ca;ZN
:J,L0dV.A@<Uf#WHY]FW#K^7&LDR1>EeOZZa]8+90^d/H:T>U1:O0V/>H,2Hc6DZ
GHb:-;1:T:LP3FB&:A]D,H]a:\+K_>NcI30.?UKC@Y)3X,_ZLIM_RaLPH=I6\668
5T]-a>8MD>L(4J_cAC2Pca.U-U+.9T.61,G21O=a@S=^UdWDb0V0(@=-;/[P<R<>
X^0aec)ePO-G))+&HIOY22K;+YbdH41H+&MU6,fVI2b=<_-VYf;:68#4fGWaO7KH
0E1H,#Y(gNNY7.7W/MUGQ0Q@)K\&XKL>=X^#[F3dNCA?-F\fbdIJ3GS9Q?LdB[:F
HJN(7@HQV&b8&b9.B6),8LQO9aa)>CIaXZNbJQOCcCA^,7)Ocgg2T2F6,F4-H&S-
(_<If2XaPc/IF9_<M\WWU+(e]19T(\UG[3;PELP\#5J=HRGE[GcfZ9?VFOQMI))@
X:<I5\KF_0M9P+S#/>IZ/B&/I<5\@ADM0Z/e1#+XEOYZDG+],QbUe1a2\aJH<W.2
EBZfX)YON[4N&T1\41/&X_;>V_])<@9f_ETWb.VdJUP&d8,RE<?RYYV+NC\,7.>S
._PTN\3#5@#NW0c]AHgEI;&JQYaEfCd?.MXG+_=K,(2:7BU/f[B)X9SF78^f.Y.X
\?R/JBgTTU&K#U@.9S7S5_=K=I?&[_ggRe),QgfG#)<TYKLKLN[V8]AceP8;R?8a
?^A^AX=E^1Q8&2a;-AfRYH9d_;c74VB_\Y=EG.G7[>Q#7#T6Hg0@WX.@^cF^_B2+
HV<eR]?e48Z.DQ^S-^>:TdMNCbSTC^9(>W1fKg;:O(-VV@Z0@1_/\=AP9[fOc;CG
T:/YQ;:+WUb(_4;Ef/03A.eVW3A2O-gZQ6g(O&?@J[[F\;/MSV-<M7LgXTc\0a&<
^I5FI<N-.L^V9\#I#XLL)4#8[&/eeaf@\[O.a0(Y3e#06fecEES3VK,5&\]_4H^e
cO\5+FIYR>-W9F?7(\O#E?A_-N>;6#WSdI/&D)0abF2Y2dU:+)?E)f9FZfL]g>F)
@g?SAW+LM+Pf.@4GF_fL#K]:T<YIgVdK.2(6&X8W:K+.5_QOOI7NMK7G;D:DFL=#
M-EAW1ZeDALDObaMH,#7.\+?O-N_fVa_2e;L1YEXedN1VO59:_Re<2[F2KE.Ff8\
H-1(@PU<0=/]N;F>/VGS-7<[IaJ/QSAd7QXIAe<12P1);@1+?#3G:PMaW58AM_gP
PX;#ITYRe^YQFEdFW=[+/3\2)f]d_@C/V4;a5)b[:+^W23U_g4@d4L-LM6Eb6STf
&eADKP:;&Rgc6D8cJ=>4A#W-8\^17eG@EG-Sc^[2Z3E>/Od\U4W104Y-IVaA8OO&
BOC-+T1g,Ye.,>6H-4((B/eBRf3VR>GO+_QUBY14D?e?8JQK0Q#e5+B>VO?WJf/H
@aJ3?<.2SFZ:-B@:Q&0egJWSL,8^Nd9).H#\e2g\5U,c0<X\WO=fU:.\@N,A\DHF
S<JTcD@GZJJ>2?0;U&F&aK,83>.>1GgTW@aHb>,>g3Q5P\JGNcH6B0JF?&2\\G7P
T5Ec[O\NbSE0)J,@83NAMg3<7=##68P[LL6dFaRWGN,N=UdJbQ7BX#CaG\^R#FGD
1#G/=F.85g)^EO,WA/e^?)].\S]1f\0UW&VM[-X/639f=F[XUFUMIdGX<&C[4#gV
)7TIUF.NFICV9^CXU-HOP[>0=SfKQ0^=4.CTTFAMM-(\(FFcYH&)^PZ,2Z,<2,I4
F6LQ)-_2_:ge7V-_G06Z?W((3(<a?aIE@4L#]5cLFEJN)cA&Ig[6XOXQ22ZCC<1>
\MOdbBX=;);F_YLX1#R;(&,QQU23]4]75ME3LTS.VP<:N>-a8H=#[(U85=.^1V1)
6d5[5OTZ:-ZP560_YK=b4&.E/N9U\^9C)S0eV[1\6AK/R\MW5);-\V>^Te:UY@2O
GJ)31eH:[]Y[,@<RDG.b)2QS0VRa&V9##+Y+,Ib_^^T<?RAXW4SP7X4<11Ze8>cA
^:=.0bfGEgGbTF)IeT>A4[S4c76D3G.NeZBcQB&99UbXG(KdR+AG#JUCeA0dT?BW
\#]D#YDX8(SXYBAY6/4B;.S)\+G8XW7#<G:(M#@Rb?fQ(]H=1YNE3B<N.W6@\9=J
S;5D\ENg8g>Q;UQ6_;Fg71A+Eg[(.+aG=(,(X/^E-_^(B[fgV(^0:_P1L=[9AKSP
3AA>OK4V9]>+S0>6CfJ)bg@fSOTgf8IDP)KN-5ab\UI5@Ha),S>OCU?GFUGR8040
1)F52ETDb2?-4W9f70a56BXH2X0gJ=13,NU<=1,d@J.5H9Ibg&A/=8g&H@U<@_/e
9RBf0.NZSM#BTa6MTC?NCK77NL@Q(=C1:RZ/#=f;BgEQ9PY;>c^I#;-536(RF03e
S^6<:=&QcV45ZSaLKbdg.C@J.OO:13O5=f>V=YZEM8UH_I#>+)(:)92^9:NW48..
^/CLY+-ABO]f<02B(<@-J82VEZ];G;5HY\EURcG2fE62BBRf=Y.Vf4e?VUAGJV,6
KLb3\45#_PF0[ZH(^Z.\)c1B,Bd2+,22V&2XW4=LO5Kg0)GK)4_LB:[JT];@G.N>
Tf83,2M4MZB.bBQaQZ)TBcg&=ZJLA6^(W.#^c_8,#bUc->RN>;V;R?+Y6H5/3Sb>
fI)+=ZTC^BcW\EYfMQAJf\JK^>G/8A;G)&aH#N58KNPb?UOe757^LNA.&(R)L\g_
3Id\N@JFeUa[Z(aK+3V3\X>^Bg61&\a</O6[B70bGBKf)H9F],NPR-a&HK:K:F49
^c?bJ__W(TT<9<K7>H?g]0aXUBcNIX]&Va41LG+N]eB96V4>dMEBg&32YcXb#>8(
E#/WBU]S\?FE(R_PH2cPCf?L-SGWH2@YG&0)fC1?+eF_b,SMS^c=)9Y/c9G^_UNA
=E:5_?HTdTO,KgJX]<[F>@W?=1c@T=#Qb/)&:5?ID(JV8:YLgUE;CJPc?QLd,M]G
a?7>64RLRHH5aVfTKT,)[8SO\P?\dUJ(EXV;P?>G4I0&&O73D+)QeY+N@0IOJeD]
/c4I8RHNCKdNK\VT+ZAHCBfY2OHPAbLA3I75,-/E<2=gIWS:Wd9fEUVTY+WK#G:K
D]^dXPFZ/A^ef/K[ZYf85[6^KQEbG9?MdL/O;OO>e]?a6GI\cDA[LfKMIFHb@=(-
Fb/a-6f6>4DHNd3./N)8A9Ka^b\@2I52S\M0Mfb;3Q<6HKL\A&8P8SD,Z4FJ.US)
gRAKOO)KE&#NKQ@#KTd5.HS?]/<aFI3,ZR?+EZ9dEF<&,A6Ie1?JC\8=Z2OW.07X
?0F,;PH27Q6WT)8,+a?98&G<W_BbGf.HXTYJ_-YEPZUH^IC8@]<eWD3R2F#d8/.I
T)[;38X?d[V>,-I4#&,7:MZ#;cU/fQQW)@2ANRNT^=D+3SdN8]Z1Y+9Z2J<d..T@
=>99(:;Z;f^>[U6P:>[GSF\UT4(CRRODHF9-C=@D-S5S7S68\b^YOWQAE[6)SP?6
/E8OZJQgKD0Q731+)bcC=#Q1<]Le\E[9+S>Q<<8,J[cda]L=R#&MAB2AR>Wb1)X.
-MG(eNE.=KZW]\D#.fgW6<3\@^2CX[+?4[TCBdc:YX+3G=.J(7ZCdeCQ[9aJML=U
JN_feV>Qbe^5\_D9?<0dFIN?.I[KAcCa\E>H3D3e(CKK3.Be/H:OT5TcSE_Y1JE:
[^=3gWF+49-[]?^^.,:WA5-^+W9<A?XDL+4dQ)ZZNURLB^T9X7B8S-_Te4D9-_,8
+M@dW&e^OQ<I=)#_.N(SE4-OL+4BEedgLD<W_c+a?W.@IYBcMcNYOMa\J520O6T4
.)9#c.cE4(=\WTgC_D))I:>&-#cESXe9]D-Y>&H)LQR<MBf:+/KWT\e1MAAILd#S
KQK&a49Q57^0RaH3\CVD3L)cWdI[\E#-=SAYgLT+ec0+13)46+N\].UP<Y_)eZgQ
UK]N)SK/f5T,[Mg7<)Qfa.L.C5?aNK:E=(bO>HD\S?]QMX6>:DbWH<VX<ReS;-_Y
B/N-d_W#WU6dEV+H+FS:G(W<\EEK;TH/:<\&(RPLXA_DQ8+F:YegG3[3g[W8)WOA
[I8)b:LMU.\XW\G=TTaeP,_Gg;]@QPT.NHVIW@KTFB=<fTXQN9^G2a.]Y2&dN9aN
4]HDEB@Z7dTXYPI4[Ig/<f8[=Ne]-@P]aPV[f\Y_]L?+BF]^[a+]9Hd8H@@7O;QA
H])1+S:E,M1LBK8^^I&/;fGLCOA9DCEaaY]RcGgCOb]BSQUQS6gHF51XFFYI)[<)
R(:dDc2cdEB5UaV1)d(:_RdBSg#Q.BX]<9F(,1cUEHH)3?7,XB@_\KARg3Z[=2B2
)L2WURN:HR/].f)T0?8e+/<e,F0TfQ5-((_GGV>C\+-8,?^aKVSeQg#9O7G@+@b(
JF_b^f_4\_.D4O0NN5\#1Ze5=,A\ce(-5@@B.?I5LV3Y+EbBe[We\/YL+@6D[TO9
CI-D/)AKaHN7.>A0^TSXf;0<_<\beUVTFBe5TPUV9=:2a3_I3>f?G1?PM_(8?=?-
@DSXJ&6K0Q>HD:g(2W>RH0=AP@?4b^eCERE79&P4bJ-XLBG4#C_]?@024cPa@J,Z
2/TI@_:OANOK:=,g+Ceac_@C2OCYZEH</E0OI^_]-\Q/NAUF9O5X+U-+R0RG3Ka]
g\#7)@8UGCWT6D6CMF-TYg]EfHT5cZg;b9->+@c_T/P=XS87B@V1Q^DWIC,?P[c0
KV>1cYTEA5?b@g>4bb-RKeWJ4U?_8/c@GL:JYNBLFS5MbLP/aJR:8;MXf<bYQ11^
=Z;-LePgUX#P5H^E[7b8/F[WZa46f/S9)((cb1Y.JT)7YQAH_FJSW9_1g[:f8UbS
(,GeY?UG;B(<=Z.QN&1S,,/ZS+[N59=>d(HdT+4,<bX.&R9F7\+N96F>cZ/E?c3A
+])&Y)1UM9H9beRaagRZ5KE1T95/8E+3Ob-^,75GD[#GPYLbAKAHJe^1I2=S\ZD(
A9;-__6-:87=Y0>B:=I0MI:1:6[UfVFUD\4O>N?1P)T#I3:@5=e[Qe)HAPd-afFK
XZOH)d&-dd+ZKT]NJNPM\ULI\YeAdP/;#G.(QF(@aA^Zaa,^3/9-g2X\3O:#&T2d
:AT=4&<[.>K0dMaU_K#gYW.@gg=I]a[G(aUb@IYIgP0Bc)J+AQ9E@RcVJ)XB6:d@
KHLR2=00g@a:>faU46@;37?V8ON+a(;6QC9f_?U7L16N3:0KYQe#.9_U4(T=,2M7
N[T>(@(R#eaXV1:?Fg4Kaf&XK1A4D<8T)FHIZ)eVfQ=?\?2NUSU?3K1f/d->a[>T
PE]V91=T3d1a^_0a822Z0=06I)c?6J7dQBH[8Vcb2V[+=ZJ-<4GX0[\)7\0L2XI+
Kg_Rg#?Wb,4.P3&,bT4K)B=3W+\G\6[/7K1;T+CVUaA7MXLO>E,LV<5eQB8MDUD+
H3/Y_J^31C;(QIY#)4S:X\V?<N-Wc--W>+F3]B3KaAD]F),eE>K.4HG:6Kc@:DGF
A[+J0dQ08.CO9IbO(A@2@?B4YDH4I@+aFB(;H0T3CLPLWGDZ&A3@N3IJY^^QY+eQ
cZ8+Tc\PcTV5]FB1J?I;Yb-^,gFPC3R&f@9;-53LYS[XHK_)d2XVZO2(D\(42Ta4
3cZa6_<5deH3)DUdMW>XUH/Q;5gHOK.2LM5,b<Y(fb-cJbN5RH=JT1PALP/cbX8Q
Hb9O5X.::HAX^T)W[;XTdKaF#_E:GFSD8,Y1VIV-#1J>G,0+ae,EG18d<A@>=N.K
C&,AC8AZG,fFL9Q)6aR)Y[=aY&CLbZ_BP_/B@NW5VcS6C/XaAbTdA^[==Ob7EBT>
8Re9(I[)JOTN2gZdRe&e++)g=-Q7FJJOW\Z52R=_Y/V5:bSC/^[&LcE27S7Uf>72
^_bUJDC[XYM8@+^QReQN#D((ID7PI1LBeBQRg/4=O)W,aFI3DbZBP(WF:QfU0O0a
P0<D_E0<<]>/cO#C@76+(]#V.a^[\S=OQ?e4DBF7?Gg[8=:#FTD&D\?YT,2=@D>P
M^D]7YL0f06_R0]H3^ZN98cdJMRY)X/;S4P/g44>9KN(,VR>/0a9V(B#J,Y-0.c4
VLgT7dRD5g<SRM^(f6^U7;AX5-2SN^C01eOBd&C[<X#,b(eQ@&-6K^W3d/XQK<U:
K<L7Y(6NVc=]7_#RIP=BPY5]\+=[NPABSD0R>\PcJ4JL;GM+VWT)[G[+SD;EC:30
&]Cga[ZHB_DFeg\EGNAAa1O?eL+Yg9I02_KK7Z.<UG+;:cfR<Qe/GL[A_#580C>[
^ON/(#+H@_9G0UCG1N/3f.7;J^8aPc[+6P9YLL7R/L8,)?=\H(:Z@&-@<T9\IKP/
=2&DaY<\>AH0aD\Q45gUFb8>:#AaE&bMb_PVKXY8#OA,&HY9_.65?Y8ULKHP7.M.
K/?.:/)dBH;61XEKAEaFZT1L@K:;_e)3MAG^2H@VV+SeX@[TPLTO?5&f?[1[9/^0
#Qb8,;c;>1+VRX@FT^Y^f@GW-2MZ_-,YQ2]&1VY+?>J?8>c:P0d]fQL.[eR]VTCT
=VX.T[OfK(7=)#a3DD_PIT/=aSPaa2NE4JWM<;f_<c9<GJ8f&Bb\MdIIPN[5L>I>
&eFM-Y4d7MY@8]J-S\?@X#)Hc1Sbg;fAQ)-^].4R:.N&:NN1Q7:Kf^J7&K3-5=E:
HG]W6]BX_a56&_A>Q6f0#8XKgO=,AbB)WJ.I(U19+.1f^PNE6FYF++(KH]P[/=-Q
5VQN;Ed#?B@Z5Gf_^D\Z+?f:U_dc8@fU>A@MQ6]YKVZ1MC9<.(HI0QGIM;L,-T/?
b.M<]Ff85OUZ(Hf6&KCW6MGIN@HgDc>F61;Q_;ZC\I+]>3VAc2_E80?7HNUgV:,?
5<+aZ/;(bM:70M)6[</&J6=U&\(6N??f=3GRd]\T)9465_VZT.Fad?5f:UH6J]O&
Z>H^N8J5aE89S9U=9&Z\>CJHOeI^,TW57-(D5SMBcaZVLN7Q8/JMadgNTg<+#QGG
T)0TZU##&a;2YRVQ(/;7d05_=6&KL@BTC-@67<:EdPfaI4F(94]g6&&ZGJ0#K48.
/]JGf6E82g(/U-/e&ee]3FG))daCc-_bAX:6=S+Og8Qa7L0+ff;=?6B-7C^S+SK/
8_f7\ZOEYb<?3^DN/bZZ&+fL<]E/Y]ZNWCRDfG](-5dR=/.KSMHd=(^9CFIe>@Rg
VFM_TI=g_>Ggb_6./>^59F1PbAAU/<X0DN6N\C_ZfC+C<3Aa3:A(SMOS.<cJ]5,(
M1(f);d\5f(1P?LE=:C,Y[M1<//<)aa:IM6EBbVS\181)@+_EXN_)O1<5H<MCRE[
[PHU_19L9M&aZ,Y<D>#/)Ff2WS06?b(D]Z/A7B:H<4#W4A_fcU\BH45deCM/VO=H
bV<b7+,TK?^.0&30,5#_IM/[,f3SB7A;;?EgQQGg(HaAZ[0T0.F,40(aBK.<Q]28
.R&2R0LBUJTQ;/P(aT+8e,7Ca_;Z#KB#1TNU<-8/Mb=N+;XG16=]]#=WJ[Q9.&BW
5FT>]b:GO:+KbbI1YBVAc16^<SLdcH0I^H#8E<cP:TI8USF[KAI8+d=aJ_NI)aa2
TE;,b8T+?_a==/ZO<HYMKfMc;:K2,Z-_DU#a2Z<SCO437aJb9H]&K/T?>D26d=6[
]=E04BH[X42-RYALKWTP,G;ZfLN:CI<,UI0\MB5PC1240UMKS;^YP6EOEc8)HCH^
#(?I/8=U@&--C<\-5+B:[&9]=RV_J+UP&;UfEM0H3\8-+XL2C#)9SOKWY#Mda[b8
TN[)]/;?Gf)9g0.+&5[67QfMCO;HQ.Z./?BV<Uc9VTe2Kbf6ACN:aL3@U1dEeE.8
.=#?UbZ_5QP7&DK51F9SQWFb/5,Q<)Z-])Se\UZ02,G-F(a4H=9eIe<YX?cDQS2b
2b^F0]K@=39KD>G6AA\]8cYO<04O@=Y23QW<2GS7.F_/,88#L4c\A8GX9f/fMGT1
ZD01-7dIKD1a[F+0+Yd9>d8?>G2XbY+0Ie@g<-H&D@NRbT=JLbCggID5?@=0TJ<)
U6aO]H#G@G0_P,YGP;I5XT.^:e=;Dc^K7RNc<FT^AI9UZDY#d0XeBJA_.A9d7JaR
>^VR\[1&=fESedgObTZ1YYGZ;aMO/KIBcJYB#SO>?f99CRP1]:Y4XMAEKB50-X,^
@YP+\T1QV5;QBc_BXF8P:86)Ta6^?I0C)QU.-2E8K3J#J/G2W=>&7+TNN9[;dE9:
EPXgH(4UdNJRYD[-4[>;f&)WK[^6G_>V;G+OSFHaNTE_8_a]<e>]eQOD(D#.B=YR
VR-MN_I<@C[I6X4LZKMVP6f^2d1OSDUYbO2UVEcUE&OUD(CNbW_gYY[^;.-]@gU4
fMW.Y?4,I]1AV5YHJ5M\,F5gP5\cf9>T@dbR=gXc<O1b02RD+Eb0CU<EL1e/CXLV
Yd3]7W/>c2M]Za)#b;[5S=<D6P@b>F)S#W;NNL+Z]WeXaIX5]dD>+(#LXYcT@&((
PE)(5g;XC27EESL3[HUD0NFTFbeg/CKdJ<KV2^-;IdH0;UA-WIH?10QJA?:??eHB
?X6[X,D/CJ,6(@09TNZW.)I5Y(a6?NFL1M_IXE@:B>;+,:O,Qb6Q;O._C2-6AJYe
S=Kf/HI6I;aAFYEVAI2[,<0PGID700CTceMC]gSD7TV<44RONJ.Be40fOP0b&0\:
<&=5GXJ[Mf1J+_6_(R,OR:#]0cAfL[;QVMdC+BAeG-b:]b/L6:FbbPPWQNfB;7c&
TNg&,<LM7B;JN[Y/94=?g&1&7d]<\V5O/JLfR/Oc>>PR5;/.KL(;W#MW\YGPaXQ=
^Q<=Y/L5S9X2]2EaWYc1W7R0OP\HfN:#H5&?#AO:T94HIH6LE45?f@J).5@&bO[,
0+DI5Fc32b,/6aLDI7/&2<7MX1PCD:G7RGA3[W7,8HV0I+FBWJ?<1SPO:#ef[gdY
ZeI&@6(R+c>[AQAGc>65_SP3WDBebdYKVa_5HF)6]Y&Xa[/R7[3_3YbbP8L=4/c8
TH1f?R:WO\PUBd&C8d2^UTd1,FfT23A][RKK<<\D#?OD)V=^5<_+>VOX?bE\:5e_
T5@d3baQSOD&;V)LJV;#YZA8H=:8CcB45,Y)08<6cc(dI4F)W@AC/CRHdXR#BR4Q
6Z21BY4Ne;AdG0DZ)?Ed?Sgg8X8&UKCJaD;H(S./@a5)LfL3Vb68EM-ce,3Cg;BR
6/aBMX_f__3([+&@0B&cM@CMb?V8Q1QS_FU_9N\2^OH<]8;K,.R+XE4;Ba>1:SZ6
WPQ?+USOVQ<4JU5E9&^5.7G[/0Tc-M,_97W[U,+KJ#BdXWH29D>R#17-W#YX82d#
+BI>RVeD,gTN5,NbT0-XU0P;[DRWK7,2GGL;:RJ>KO)Ab?RTB#?9ZT@@6-#SeA0g
@-L)U<2Q920d0UT_]WbZCYL,)8;JJLYD(;eGITRQXX5^FeYXdSe=c@.=I7a]RT>K
,c4B_V96#Z5;>V;Y(IEM5bLD6.e,c=:,d3K8I7J3/:H&+;OL:D;F3/:Q5_Lc=A+)
TOS,6T;X::C=4cJ:8Y]KaDCCBQTQC55(aH,M,cZEC],E@_>=^WRA<J=f:]OT4DPH
dG)&UFWC2eS94TeIU2WV[8eBL:K.c4[bAcN1\M:\[XNO?6]DH\Le)eeKBNT0\<MB
;8+7bT\=@6@S]LJ0:(K=BJ0Sc@?VCE?^G/.\cO7EVJ+<0@[,DF3gB_[PR5(d3Acc
=9NY+c[Y<dEGR1ON\<Yad&B)d;O(C@1YWYgF<HLP-&+/-9@.(-I)b6cgWNH^PYEY
3aNMP1-e@&?M5C8#R9TI0A4c;?=G=Re]OKX2Ma&A2gS)eN3@?2e<6#YCUR?g>4Y?
6Hg-a4>583f8OL0gB0\gM]37gIY87TX)-_#^,(XI;ES8>1e=]Z-<2#2>Nf8=C47+
;7H[a&0XLNZEQZOA_20d\65M.<QZ4-9GALF7+BP2ULDXWbSENO?[RNM+6;U@:/X&
.BP<c(HJM.(Z-@46]UKb2/@)G:8?PV?L42UZ9Ib;.#OY0L#dNH.FK+B>E\O3.;SC
^6S<5;.FBGM\ESI;WH7Q&P5O/bGKfFd-#]J855,04TAH9BZ[(O:7K10]aS(G7.-g
>[^@=^-D>0,0;\Baa=N<b(U<ZM/b@N8=I>=^GgM?_]2@YKB,-WSXe)-<b<V9DAFQ
.7:;]ZgDX]S7Y\G@+^).C)^(LHZ(/;M(6<-_a.c:aC&L0.AMDZU\dKb1^105aQT]
C1FUON]1B8d7;,UYa/I<S@X7f]]2-Zee0,RGG<J8g.^I^?6f,.F/fT3GLg<8G;f2
85&28UPbB?(K:#D)#K2A(f[cILEX3FFX+JHU0>]6DLJ-Jf[Y4g#@H<RC/]ZW#9TR
\V1=I,A^;g;84E#=VGL_[K3=B<c^Tb/CB8aZ5J.)WA[Xc1W_fJZ_QCD)g^3Q2?CO
G\_;@WVAFSfI^.W?,5G\,-3c5f7]:+M8J1..Q;1g,.(d_-&0a_?a)+JO<LfY(C_@
a36]aP11:7SQ<DBRf,LE(EgFaP=L>;0+W(,dd=>6Q.B&DG^?/@Zd358KOeE@+Re^
OdYcdFM?(gP^^L3:LB#d4TT=#4_b_:dg0AU?ZeB64.SA6<Xc&)QeS\=1GS.@b7H7
P_dSLa@J\Z\8c?FO+5dFe4cZ-dP-I,A67EbNLZ4)3M4-HU]S595?&)BAUC7f.TR=
G5U0ddIS3D9AUc8LOR?&T@@IC:==@R&2R[+6eV(5G=J3VD\6)B7bIb(9T7W)X1#C
GSF:0=)C_<dBbB^<++gKUWId??5[4P?JB6?96D/AD@9F<+U&fU-WW@DG&e0+)L>Y
#.Gf&7@5T1=2X0+YNTKe9AeG_.J5O8\^/f[f)aLFEMXZ^2MI4N1OG4-9GFd>ER--
P2+R+R,?E][K;JQBe?5.I+L(T+,AJWHB>=>^.DMfZea?5IW\1[M?VAd&8-=;S_>.
fD/KaX+2TNcbBM8?G;4(DGD=/,+TY:NFC&Bf.W@@WVf0E+LYMQ8XM:_##C+7a9(R
\>ZQK<QRK5D+_XVVgL9PFK@LcA.5=;HN9#]SN#XB&eIa;CV_2[R1M).J>P.0g(RY
0-UVa3(,0aIdF2Ze)+^?C(FBS4X^9#B[^3I?RT5X4_a:E];MAKPU+]_7OZ>W^GFX
HEB(UCRf,/F0/^I<[/W3^]].&YU@X17</LQ\R9.fX;+2&2+e7TKE3PTdI4H/2RSJ
@&IDcb/#dC3@dJX;f1&+WeK>0DYa[(R4G&O@<C(KIT4PU]0?5/W)181.]?CNSFJ2
DCfEB]YAXc;Q\e8R-H.\=LcC:-.e225DVW03Lg_@<>ceA6U(H1UJQDL9Z,LeP+F0
_T1=B@MDQV^/CV&Dc9f./HQYdeaJ]#GJ2c)QCB)82>#ICXYQ\5B:/g>gSD(gW.\d
Z<U)T7X6aO8;TgCE<]&W1:4N5?5L/RHR<2e+Z=+dC0^e,&+M2d?8g@N5M.>/ZE--
;RCf-8N6F_<V&TJ?6I637IPb?L/6M/U=Y-G^AGD7/U^?S1/_+aFV9&&Nb\XC=Y6E
e?e[3Q=6MC+DF[1\./Zb-73=?6MVgbI(UP5M;c,+=bZ/P/ROedA+_]+KM&698ZW<
Nf)-T7BW1LRI;;XP#T)9J+9PK-:[aZf9cN.[,)2H>:aZXX/,bC^Ka(4Ba-1LXDcb
;0cA3.ce>gc,TCRdCbT8Vg?e(AI&F#M5(R_eGf5@=OU\LbL7UR>>f]G3>1d11PM)
NL#MCXC;\(U[4UC:D>PfF/P16_N51&I3A7P<e?0,2A814aBfF261&.7E2EAUQV)d
5b<8bC(=A+bWX1eC_4DcKBDeC+IC.966#GeB;LQ[M^G4K@N)G9\8c_UXLf>GZE4Z
PgFaPDE+JNfa;PQ[F&a>Y(;g__NQcIU+a,e22AXQM^+dJ_M9#+Md=#IU-O(ZU>3&
cG0:>Y1ZZf18P)(F,5R3.5\@ALR5/L[L8Jf,IWCN#VMef.2F\(e?UTGUD\HaYBW<
<KeYLeP,g)=MEJeXMB1-NHC3W[cG?CT91/N+A3<fC:O;+Y#+<]]8b^eF)&XBM1Y&
SRN9#3(aTN>dN-d#f@_]Cb^A8@Ta.V=fJ5b]-?0Vbf8K/Z+)Q6]6;^@>4fQ-(C-\
+<@;RDXN=EU,0\SEV+LC2eZMLfM\O9<3(>B+bK&\&/P310f-MQLa?DAeDD)]NKc/
[,g0Gb4F&WbRJgUIdEPS-RMG5A>4M^WGe8\^R0d_X5E#^?ISB=Wc:#DGX?C@dDU<
^#9C]V8bNLCO_VTCCd)aeVSNN]98aS(RPR;ObYe,=Y5;Maf#dfVf9VB0C3[;O7?J
C-]8T;cd0fZ.?MK+6=+D1BDQPEdN,F40G_<:26@J-+[d=P]<+&37Q=Ed-/;IJ:<#
^b^R&O)F_WZ.2NNRX1[:@d#&43TLQE,X&-BX^ZXPRUgVEH?@PA1DW(Y&eb>:6aSY
,a^#(=CNSH\BP,/#@/0B>)BAR(\DC=V8a2;NFeOMT?LD:[cb)Hf]CM8fEMea(51K
[A^bdg)Tgd^<-(I)WQ7&X5_g6NL>]@#=2g#GBHfO4[(2)[JF4XQ>^^_@,1_QGQ0,
D@&+X5C_95Q\3UMgcC]JVXdHH\F6M364DUabAR-<Jd.a^(80,/@Q07gCI^V_?8Q2
[??SYF,bNI1(,gQ_#[.AV0Q9gPfUWb-^#,+7+ceJOe?TDKY+_4J8SFW5^JbcLgPI
e&&0/e8Y:5,G?7GP_a9\;\A):MQQW#,M#PFba)DQWa(bVR(V]M#?[PIWP?LD\QF5
Z=R3fZUDK&J37.MK/2YC6Z#Z_&+8#=;_70KBFHWNg7M?O:0Yff=#W6:3[T7H.8K1
O24b;g-XEbHR&,+e@(6C?aQ]E(]aV1-_OY0KQ3@/57ObBg@)79X14H,-,;@_63f=
GM+/Q_LEN>&eE?E_8/W2WcgA&<D,9cO9c@A.Ad2ZBR\3(TWW.\MeKQO0AT?eTXNY
\e3b>cXJ4HdI+B9EXH@L1LD0+3T^^.D5#EY&26K3gKOZeefGeE8UQ_GUFB/2d2-a
f.3_RYPgC]eIdSWbfV^a/.A/2N3(#cM,:<SZ4:LGfK=9#_80?.=\K:3=EB86RcH<
HOGV9-1#/LU:IdN/[IZY@B1V\)2?Mb\DL^W[+S\SXe0.:^HRBR<0Ng^0\a,^03):
?fEE964<Ng/X8:Ef0?DR:^9@49HX]118,3OJd12+)&E@IfFVH.?R#3eY>6d^T#&N
,.]92B+CQb6(beEZL.8BFJ:S^=AV-0-=A,d[d^W).H,G>1I,JgBa]He(Z@@\5=a6
D<<BA):UCaO4)5EU]g54E5RL5Q9;&fF9DL/DUN>>b]L\b-a2Y138c)MD\OG=NZF<
aLYMc91BEP<BM2_>_([=^cP;JN,6-@E@f&d7H^M]:C1^d=Bg0[0DdDb4TZ#4;1fQ
AZaXSTZQY5<52ffUP[#94V3(YF7=&OA6Q5PM)X(Ogd?;f-DU@H4gXW:Ia+&@N#2Y
#+^+L^.a#_8-Z:,CR3LLD#:)fXX#9d(10:ASZEdbOIG6>d#X0FY9UMe24<(MH9F7
ZD61:(RZP]Jg0,GACC9.H0O9]YEV7.U[J.ARP@gCR-F4<W@<g.S3dBF4YM=Q=dPW
XW/M+PW521@EJbZG0e.MgO.9I(VN7X:C_AG<#e@B,4Q@4I]/Z<ZP^T+K;0;T[g6:
G6bD#&#R3FCV3^C;3^D&d/gQGON)>2eD9<Z=@G4P](L=H9cM?bOH<9e:57PFISgT
Y9@Q)1(G9,:,[eZ[bJD@]FgGT3VSOXZLR:/^QT47.5.d_-ONL-[Q);T6e1cRLHI<
>8^T3[LMF&J7_R.c56[W[4G160c&_T-=(\ebXHH?.6D/0O-\bbb05KTfXHCJ5g\O
E=#&E>;6MK,O0OeY_f8BaWB-,^=RB99KOUALJFA_fCZ/IXeVT0,,2E]4c:ATL4c_
a#FP/HeM+1&He\^-G8Ub)6OQ:106dV-#FIeZVLH--fU&See4/J;WHPY;<A[3dXRY
d?2OX:UEc5F<&C/4FJ1^ZRWgR5HY?Y\eAAa=V2GDc&@,#TFB60GUSWAWTY\^LP4(
J+53?RWN);@KEPg.\SS^SgC2&d&P#0aLB)f@K8L[_860=&e&HB2\N?FIN99/FO1O
dV+a#E>CZG,.V.^Q7bBLONMW??,7K2c8@=_//[.BW4PaLbPf_GacUI(.&17OaVWZ
KD^>OR2+c5/a1(^J^E3Q:dXWC_fV)aX>(74_d0+9.O/@;]7^S5BcgF2b=3gV=R&&
JfcGV-W3L3c)U3B&>H4L?Nf4_eH(=BX^JV#IK+[3C7bKT#6#0_PHWMI_(/7bgdUJ
5BYaOX_&R.W7g<&Ig1<8I9F4dP-M1T_P[B?/aR8AMgTeOfNFWO8ga]3IA57:>EIP
RP)@8?F9J5fRdGXSdR9/L)2Kgd6YO)Q);_+6.4KN^&dP?_+_PKf(UO_fKI)-McPA
2#E/EW+:5.&F5^LdUMPI.cA1#&O.#PC0&>fec.)(<4J?.#W+A+6gOLIXG^@OCKC+
S??1_\V&U>D3L<)3,[5f43N/5;#EL<5e43CgATeSH4P,;9N2SG\V&O5FU[94YJ2g
CIMT2,[ZGU,.<5MP#.G,AJ<SI;aOGPO,;Sc8_79@cS02>1.4)eSeH0F=V8a\MP.S
FQO&LH7SOaVT[fASOA)W2Z#A5<3^K4fK4PRbQ[G2QVGTX\GeEH2b_RbHN2#WTfea
SQVU_SLXR<<2K4QZHY.aKFJKPYZ;@PSBGd5fZS(&E&PVDB+A]Z:Me4/&_9TO:2:3
1(f5GM89Z,I#1CZ\Dd-B)Y#S4Ue:5PBaM4F/&e<M;DX5Y-,;DI13M1D.[4U@.\Y\
Nc/D8a9WDUKQO,Z/F-JLL/]PSDeB>d\R68KY7aYR_4R[<Kg:[Mb2GeP4U-2cBG22
N?JPEAQP(9+[JUfT+aJJ1/K4E6E1R8=d]3(.5<_\YZe)g8??RBcLSMCU[/L2VHKI
dUTE/c=\VY#fYDVMGS\Y=-.Qc.U([eP=Nf8;?C--C5G?@<fP?)_PcM2VgfM.CO<d
2c1KF(6D>DL^2cBV-KdBDDKRW9N\H^_L?A?.)OXQ@aEB<G)=CII<d8T>Ca0F/9H(
^_->+K?=QJ([Uc<ba?>NLF63ee<\cTOX)a#36KGIIfEU\87XIQT&WZWY(\V\6Wc[
.\\1ZG<@E[8P@\(WbT],#@XRd3>N&?<XM.4A;3F,F\:Q#c<NK/b[=MTcW@17AJRS
1/D\aBR.=N=SLR_d=5H>+_XSK\H,@Z7>\VAMAESLc@9OO3?bES2XYe^NYZ)AfQf/
/U?6:)]16Xdd74:ZA3M0F6DS;UPfSE_U,QB/[G[Nbg8)KV]f_CQ;LaWAH8C9#E;L
#-[I6e+F<^_-K84S#/[cAfW8H+\Kf,2&>/T0Sc1?#6[HeVI?P5VbZ@H0F;MaK](2
HKRg-Y4)cJ-S)A]^/TC\[JMXGEY^HW]09a).dS1Z\CL<7<5IBT4IG,+_\f_+:7.P
([UfX^^:<I(JBc.#Ic+dfEWc@J.T,PFg^B-c+DcI-\A88BI1]E0IX1f(CDI=:Xc<
CFaQ+VK/=bWK\>UBQdKZP>L4IES2Xd2=0&ZK&KfbQ&Me^V\(3J8eQNAC5-O:8gM+
5Ya&7PHbYQVE1&PW3Ce]RB;BR]FI<S#.F-3)RPH()J]g:P#c-DB^G>4D<^GM0aB/
f_KA=d_ef4<A&fFO&:KB<GaM-X#I)V-P15X^bK+dXT5K)(B^_NOF6)IGfGFabHUM
SI1E(]dK)BNg:K^&EbBaSc9WS4,Q07_HZ]WYY8\L9]T,0_-5Z=BaCSK1TfI@J9R5
RXb/54J&@;;ST[cITR;F#c=>(L1K#2.DBM<I1UNa9Z;:&C3.&#)#1X\EJ&,_9BX)
WSE/D:ef]IO,IY7?0EQ64(FaL\1aTT[e:dUO_^:g96#<Td8d:1^EZIC4KXg9DQ2\
0CL.REF-&QH1CM<4XIGb2a4/a^26+Y6((NWUAG8]cePAeI-B&K&[ZMfAZNQO1dLa
9.VFd.,JN#81:>Y>EF0A8RK:M^aUWS\H<HAH-L0=;[e^Wb>X4Z)/&E_:?H8S4d&6
T.&R\bQU^CK&>4^PTEPYN@^#(HY+B+Yg^LY_6(O49+bB6d]GXcH.Q-@B)5BgeH:8
/c5aM;-[\gJJPOf.84IB9UJbN1:A+R9&9S-9.T#=KL_f/Y:DfBV4I82M[S>gG-).
RaA<gKAAa?cFW18\Q\GdSKb>g[W5F;\ACX-^UKJg8_UP3?(JcR3/cCLZc(.>H:@b
EK-;P+/&E)@g63LEVN#/W053:&g6[L./#HJ^O:fGAJ]>P)1YN7Y7W_2gTe(fOb8(
Sb&+=V]9E&f5RPVffX?=_R6aAc2KZ)5#TNNcFJR,_0YK;fOJ@W,UKLSNV4-,V_Y8
6TU0/?H=<4@Q&RQ(S@Vb3I,2-3MaV8NUMS2.M<fFS]MbU:WJKBW3@)DMg69&ER.U
,5U67>4U>dP-[6EKHZ=Q7[Yc&9@)D7F>ZOEM8@,A^.IL6Ua;>cFZ_Zf?fZcKT8-g
X081NF]412/4OG@6<8Z(Y<=#71)P)_UTG_U>)##0-K1;J80aRH<AXD#Q=0((\dU5
9N-[VdeU:C#Y0&]S];T?<1[U?J@,)M,Q?3Y,2DTDN6CECK9/M.g2?HBd]<.:#7/(
1ORR9DEVK-AX]/9.+f&RC9OAZ&K@,ROc99HE3OK5:8)(5Be8?#b79@=0Q8JJaWLQ
CLVg7e@9>Vf#F=H?H8#68GAdaK#FQ7[[.XfTV\B][D&6RaO-f_V6K0&O^M]X>IWM
Z4#_Y8,\#P9RPQ-aL,/.fLBa_#.44><+T6^K4,b5QgS/_]X##1QLJ2_\358&@T7P
C#.:=M0U[QGIW1+W/@_IIDR4SXDMUD#OfVJ&_X[#,L&D7f(RU&]V460K.WW7a\_@
E?P<^D]>/+S9W^R=[UQAW]gM.=]9)K]>f+[E6+<E.864L@4dd\U]UCfSB)74SB-C
N@=:d/c)E.e0CE,F6-A.)E<:TE-:B_/_&PdfcLL[.:A3SOP4Ne#\@XUTQ/VWTYd,
2&>\OR+BFe]IH931E4->WaO9242LU@ZJQWf,<+[)Ka+ZGZg:0>LR_9fKgNLf;b-c
fOD)Q8-.@.ZB/2a7eT3b8KOL[e@BKT.L6U4AfN#2/g[CVQ^#@NTX<0K<_Z5W+:SW
VaIPBGQ&1gYEVg=AA_LO22<d^^VcU5]ZaRTR]#^a=9>J?J&QF>.G,c61L/Yb\3Kf
Q=8c&REGZL1<EY_<U9+/P9b:>.O6-^0eVF3110J&94E466JLS[UB)W?8_[YOMP1D
^F7aH_fF&R\MF]KV5I[#BZPDM42-JOY>Y;Z5H)c3d4(g5ZT6VNS_]?<]L625JSF1
gR19^16(G7V-A^8T?1.QPf:FIcb.c0][(XUG[gV0A/eI^H^VD2aMV0Y;O6CNBDG]
+B]]_):>fOCBG08QKS&[#ND;W93^LZ6/-VIRW_Qa1KdD]\[_]8fg?A#gE;K[H4[W
4NY==6NT_Z3D(M&&_MV((/;UXHg,B5;d4GX0BWQDL;>)VD2/fEb4XWgaC?&))49_
M,&==3E6QR:I\8fJ[7)8<P_eb7-bA/\AF[P0S?Df]LAf\1DSQ_2YH_JdBY]KR1;S
<F;&T9YFZ\Q[&7Z];ACNO/LH](Z_4]9bRE4g?a7OY@\EWgUN@@(@BE9IRM#P][31
09)]=UfH>Egf57@Z9)Z:_<;_:4W/3KRB>_2:;fR[A\Ad8Z^FS?Sd\^\,d-\e)37]
/9KPE:/FB^^&F_-CfWW#YfKdCR.FN6JRb(a>\W?LGPTTTc[JfLI5@)5C39@6[a4P
dP88HJDVe(VQ)eWZfS+S+?_K+M?XWS6=06c2=3(EK>L^;9RHQS2CU:G<N2XJ9PLE
YecY@MV7I6>V&ZXP.)GG?9dYR#KDf6X[T9AXY4@W\W2M<da^[3^T.&.#]TTV(D9J
@X9=e(0]d+,G[25>d?;H[d?dacT<B-e7d?PEIRg_]E60H0A.KGZL3IEa7[<PI>2>
4=N,10]X=GV7_F7C0R)M>2.E&78(cD-JB_81bAZ2^C6DZI?:G\Y8bGLZP1COJ)_c
a-cYd2d<BJ]GA8J0Q2\#KBM3ML<>7CXdLY2bZ?T-B(QYKBaHf+73-X?)#G8M1#@V
aT,e#M:ZK8J,I8];FXTd1DY7?>Z\AA/e@eQO8MT.:8+6<YMDK8EPX9YdN7V32X&\
g(,W+]e=W=EEHZ6d/U.2CM=X@#0FAI\MWJ)1:^L]C1Ugd)UO_>4M4-TaP^PH>9TP
KI&MIT]/(_T@SbHMG6P>a6b49g,K4#Y@dG@H3Y>S/BU;4862dH#\JGfD&GGaNgBK
DgYD@R.Y._Z5HRT#0F.YU\T1KR5EW#Y-Y&,<J)Wc-c\TF/]4KD6b;J,>5<g93=)X
;,3LXA>RV(5QE4]Q#077VZ70JWBGV:=e27=a+?6HTU9<CL:96&TbY5T)V5)aSO3K
)V8J#DW_;J1UP=TDfB=4?QE-;K2#B6F8NI&U14A5&<4+Z_K]AW(T8/8:=1:\<RXc
3[=g@6#gK_BNMdEf]4TQJ/[RBg(R.NZL,+K/-0=5d;0K+]1NVC9#WTEVYf)O5ObV
aW#N6SULB;VHZGV\)<<P2C[L6Y7Gf3-MSTN:cdbe5e,S[_N91/QIX&>XL)P(gT<&
<Y#cK[X=9+KR8fDC)+Q]\;ZM^KL)PKGVV&fY>^+U)K/?U@]F#LFCHF)]fPTY9&4G
E:c,SUSb(./9#NX\C0+Y67\AJNUU4)/R+R3/S-9&UQ6F=EMeUXP@1J\01QLI^RY4
fIY15C/A13[6B:;7^_=P9/Z0cLN>,L/2P\DBFXe.C[dMO?O#Ba7VOQ+L3^=LN>M.
?/?C7;+U^Q;CgOWS]=V+1#_HK8[7PG[@^P>;Q&CR7\=]B,>;H7+;O0dQ)9J3V3^S
R6^[B(]V^Xb&]W:CHAgPARa>e@M_a0Z@-\_1=F6=RS#5c;f3GU99P1bH<+_JT.g:
/J]T(MbR/VgZ,<<(U=?1(,(;(7THSISWLC+H<C()<I4>CV]0^6aB6b-MX99b[&D^
/NQ=D(<5]aEC+0]31UJJg80G52,2PY/ZX80NGLB<UDEJ=CJN3J/UDaId?9-B/;7+
=cG:H>d2K3+e,Hb95IO:FU]:;@@E0,R;a8F=2^Rg?YDJ&:AJ3+gc;JEK[)3[5OTO
)_DO8^=Y[:0Z(11B&]M95d#d35Rd&<[25]F@AFWNdcJNH4a?LOK&e,45AN=FC7Pc
eSQ>@I25+W7#4L/dXM8@e>62I9&0(Z[&TD\7_F=B]?S)./)ZFCG#??)@LHbQ9E[1
MFE7gX&:7YU75g/P>25U_8a-V:A2O^C1Z60GXYO2<Xf2+(WA:H9ULVP/RKS2.4ES
6g)Z2PUg>=88UdVHG(DMdAHD;.34?07YBa5AgP7_3529_^b)3FdBW_\]0>N/;C]O
A#PHPH+d;PFIY8fPUaHKHfPGXe-VE4E9#dK^@A[De(e&(/MV,<;:JYN(gJT=W#U]
\:=;gNfETHgA-+1B85((dRGNA[[;J+4T:KPZI>T^9.?gbW-;aDLMKKP7D>G9AVY]
e5BEBJf#?RC^&W&F9F(G-<HK--@VHL7IXG7d)P33K#)V]J38]9gPTS7YQS55R09^
2RPR+Y.QXQ&ZI9Y>C8d^#99S^X,NUGT-8:f3CL?dX(3958]XfNX@-R3a7NN>^H^e
b3BGX0\=R+:Y^A6Z9RdT_K:+J-\9014CUZVe,,5.)fJ#dD:cSaV+W92IU?22&XbY
fQZW]Lb0fPZ(7=3BN_GDb&(GAED37CX1800WAggU80a63fJ1DO4JB(#<&V<(:H,#
US2RdP5<;^VM/IU/\-9a3/a.T@:7F[3:X_.<AA&+)gK)d3QTPgI(=1MY/2EQa3Ff
A00ON0cW,3PIK?6aRUR4;/^:+S/DdO5Z3O8ZNS9dg-_Q5G\:XN9V]AcMU7[a45UM
#D0#DcRC6Z7(E;3THR(^W8RH6YDa:P48If)g_F]2,^b1>,V&7EB^GaP+.#WG9@X8
X&&OYXS^SX>&1_B1YVDV&K3_f0:-Sge-/A(O[-:RPY_@H)a[AWAGUMa=NLM\)X>?
\B&S:Z\bb7T2&aW)U]Y0ENd+\S4#8MVe#gX_Cd.DXCPT]Q-=Kc+7[[3c^MgYbB<O
V&HIDaGPe4GQIKMKJ@X^GK049\.LV;ZJ-4e5;-UG/W,O6U1D#,4g9U\9eE;56(f7
3B)a-Q9_YaH#)A7&bORg->T1)Z]W>/QdeQ<H4A9EKB0XH6<9XUT)c^C8_AKIYf\E
.c:P@A@I>J.b.g2;a<RU78-RBL,.ADWJAD&__.A=<&B-];H&CA:<B0R]1^CY,c.G
9[fZL(VXg:::GD3dA:JYITg_gZAC5cM)AFN0=d3OL+V(EWb_gJaL;#4))EP.R?>N
G9S]\.g(?,9]S#K8.Eg.RN5##>fJ?5B,)^8&&7)Q\\5?a.;\e.N6N/R3?#]/:(-8
,(]<1O^#R)LQ>0OD27IOcJ_T5QDTUddI2L3KPe>fHG.NTP:E?We=JIRaT(BTZ14<
E?TX?2Z@4;I-)#^;,YG)75(>;O1H)=bb3.V>.3OZdVBKD_<HVRN)^TMROZ@K#<)>
A4b(OQN+M;.S,GbZWMMdBKbQX^EG8Y_e]73.)?Y=gM?3NAL^7eYR)cJ@b:,_^9(K
g[[9E?0cFgQ]aeG#9UYO3g?J460^BC#^T5;e@+RXOfA/<PA/-8Ldb_QI@47aXTa^
DLLAARf_]4+(2#-Vd9)6)[PJKGXM(;_6=2GXT>W#R<3cea9[2W3-QDXd&d5^EBP2
=aUZ8aH_G2RdfSNPTcW_32bC+9QS(5)/,aEf:<5/4PR@c6RIA,847(K^;f:/\YY,
IKf..@_g2YMQ5F5.[3YV4G-Hg3H^>f;\F@gbU#C,dY5^_DMH;gYME[LW]X0Ie]T:
M5f_J[NV<1R<G@AX6LU^2+9aRAKT7/-<FHbTUKH[g/RfIWc#=-S6.-T61c6Q8[Ee
YLCe>a)&D&XbHP#4]Uce0a3<LXL&=5EIB@QDaeWCJTB6>(b\eK\XeIEA&Q(+dI,H
CZL.eE.I,Xa^^V^gMAS5A6Q^#2cE&XN7F1/c(L/,;=a.-f+8XRQNV1ab-O)7<,^c
PB(@SM03H,1I@+TS6;&^GS@0e=S(W:d)P8L(>X^OSZVg:TNK;Kb0,NR5@CG<6[C#
Kg(fZDT98_+aW_A/15TN&Jg4aZ5SZNO@Y3dX--AIBaW-3M&S#L..#cY@;3S-+QQ<
>U5\IK9UdIFL<54M@fOJ3>R5P:)A+5THPF5_/@ZPJBQPR.dIb/0X;)/@45c\#9Ob
G0ORBY#a=_E1ZLLWK#L2(,ddJT[1:N[D3+;SbN.6Sd)UY&gG3_J.c_8WO\@#?_<N
gY0g+BN25VVPFK:W(7,<Q_Te9?FID/MgI^_PEcOX@]9JSGY5;)DcgBf]eODdO51M
_T->_gL,_.d[d&e,BXL/USPO]R>9.^<^K:([d_RPC<90[XE4BD7deY#UK4M<V0JX
C:7F--E#)32DQATN.->)\9)#XLAU[:25_)L?+AB#IORZ-dU#5[9\E]^7.=dR,AN\
V3M/EOW/9M-2:XFJQO_DTSXXec79?BN6HZg:1:;RI_;A<?D:V<b?V07#)?H<;MPW
a)U/VBT&M#H)2AB2Z=4=(XZ=g/AAL<12;F1d_f-3C=><=J_N#G.^P69-.+8_ec=F
:Ia,cHD]<6<XdO#eAU+M9_DU#_=^].<8KQG?DH0d6<L0(#.R969.I4S2,06_#>\C
X2gX=-K3M5G>\I0?.\</,X5gLF)8Qf]a];fUK&4.5=VZ^P8(P94=bH<I=K+F<d.K
](8XQWg16S>=M?6KN4;8PIZ>7=C>@QC/3JSG.:S1[fQB_/b4OPN)9]9?4XQH^;9a
I1ZL#SBBH-@2?[7ZG,=A[HL+@5J<N44d.QOZ+QJPZ+0^(1_EaMU_6E,T,CK;?5ZF
-gY)dR.&[\@R(#IR8D3b+]AaLAKR_6dD+2EV9_M6e:1H9)A5PFA@0<?e/@GUAQ,F
fG2?A<,^QF6gL0.ITfXN4]P?BDBDA#&=/Ib^W)B7@2fX[VGI@H:d2OD1O0Eb_ZF5
LHVP8Y6=46BZ-A)H:HA,4b\Oa5^ZgE:H5FO]ME;RJLca6J#[cRZ@bcXgOGd@2Vd]
?R)<c_fY\f2RBT-O?a8>LaU\?DCWAc.>QJbG[0XRP.QW]D:M)dRJ)OVdFd+##<a@
HcE^b><g1U>EXee>,I9+Sc>C]Kd8fVfY)JC=H29b4\61XG5CA/]YJFaI\I&e6]P4
-WEEPG-)A9Aded/UI1\Y2JUC6O42MCAOXfR2Y8]RA7]RSbW?;.C9:UFaa(ZI^EBL
MU2<.XZgXM6(BDBT2YeUBR+9?FX#-fH1B=a9fU^J-a+UdWU#4=TbQ\aU0T>^A@5b
Ia[?I04-8gX\FPcX_e:957P.1I@V3J+(WK1=<9BQ76>-QG3(ED34JA1(EZGfA(UI
7)SCJKHR#\SQK/)=<3H1^Kba+=HbGYS)&;G#6CWFb-MH?TC3a[=fHY+.;8e&XTMT
CeEWETFQZ46F+2XcdA+Vc>-TZA-T&PXgGZ)e>WJ=(1]0X&dC<8GbF]bH[R/Y1^LI
OC=,JKZ&PM]]bG)G_D]-/=>@/a795bQb<PgGAI\[6VH_M3C)9#)N/f8(I8A)G9.8
4?S:(1.#+[5S4cL(EV<3ad\&HQee6;ca;dP<>K4C)/b8Rg[X9\&)WQ@X;AR6^A5L
ZYYe2E+?RV>UJ.FLQF_Y6TK351N)OY(PPJN[;;N\<#0^_X2K0K5gYA99g&d5[>OE
H<78#,>e4(=BVb^5_ENGO2S>H6B48FS5QFMWVS;8g&UY/[7=@QaGdCLNZ5b-NUDS
F[KGf=/5V7E]^G_V<Vd9VSJK.R-M-E]eB^N_Bf6?>@GVbX?S?;(D9f5/b_#IVN..
7<21#9,Q?E.J>1O]N;[Y2,B2:+_3IV^[#0XAO.RfdXg^B1H>ULKD4.DMVBF0;=,f
N>/a7Q,W\>YERP@.1QE@;AI..3Z5[ef5Mb+S\CI[#51O&517H947)F;g\BM[gU;:
8[1@?6#G[F[18\(+/QMgLMP]TTPg^b-5]W3JB[10>9f_6<PNfC9=\>?37NJW_FCG
K;3f,c(EFSeaJYcY@RHFU_-#:Y1_JFE2fM&5?^BFCcI=b=(c#b)=ggR0JMcP7-(_
<Ka_W.9I27/B42=_PM59U<?EN8[bC:UN(YJ,UZAA#4OYBfF@^V7/J2M.dUUAYIYD
aU#9SL@@<ZS[Je,F_IY-WAV09PaPLWGP43LQN&L@M)TBf?OdTS_XZCR>G<9D:S[O
NM#f4EAaDF7IETI_#1HNG]NaOV;OaX\=I,Q>b14BO&V.]I,,DfQNGA1[)cK-Pa,W
d[L7#^51dNUY@5:56T9VG#?\K7,_4c>RIRNMVCVERL;XRY_3&CbPa+JZ3&V&N)&,
.U#HN)#6<fQegBVB/((RcIS8TJGX_]AfLf\#<SJcQdfKYX4d@4_TEXJ3SALNg8)E
.(.8?VB&dd6)>GPUEJa/]ZQTfZNL&-Kag]M?+SZD5,=>e^SOX@9-)3DfFZW[g;\3
\,-d/)DOfMM;_a8.e6b8,a5E)deCP\@E-+9M(0ON)L]02Pg2/#=9W]g(^/f+V#N4
U4R<@e&E<&&Qa#)@8Ub]N-\=E2Z-Y4HeLW)Nb+2aEG8;\Q>eZ@dTCc_UHd9C+R,-
b78;f;I&#Kc>RXY1),D4CXa/F8:)VYQGB6;DE(JeD\V<3K0&P6SgKJI@8<Zb5#dC
J=E9?3d(&e=ff1T#+Ee[L(H-5U9cGDHS8#,M9.9A[SOBSI,[E.AH]D]#A6AJe/@5
W8S33_AX(d-=P7Z,TJ@-HO/EfBB&EM(Heg21EGgJZf1b02DLLM8]MV2LV:?f]LPI
1L,_\2bAV&0G1TbO)K:MX,80@a+_B\>TM=WXCK#?5Z50?+E@6[#Ac].EFJN0DT@6
PT^;9QgTM+MI.8+6]\+(<NXH-(70QU66PZO[Z5]5IJ@8ZNCdNEOgIHHZ6g^2((b7
VH5X2VI9YM99XH)DE#U@-OG6D2=]Ie48OD[4(44ZP2Jd5H?/1bY76YC_K+]Z:]TP
N#V0:5^1NZ<^Z\21_#[BC1.Y6dPR?MSgZZ-;#C_HcS?P9=CFD/=R6.X+0U-0F]R@
X0Q+D?<,C7T_/C0Q<9/GLNaO89.)e-X/9RH-+QDJbP4Hd2:U@;Ca#<#F?ePB+?8+
ZRY_f<LQeK#)7GL6;J@M(R.4bXYNR\WK)Xa9+PYR8d;?1)_+6FNL[Na]H(&b-g#.
ZC@@GYO83SCA=a7eJa^K+8S,[[7ebf&,SVRW4V39R&]GMRQD?Va.@C2;E,;N\_P&
LYS5#1C6eAVBL2?5UU,3NCcHI9J-G#A@K(OS.4;;QBa_IQR+;](X^?a\\-#SWVYc
C-/MV^,CW8KS=VcDKadDDC(,(^e2=E5&GU)(;5D^[.O[e:&8ZFaQ=57FP>.V&<EG
75P+E;J^B&/_XRcQQ^a79-d:(XBc5:f6;aWR+WW60cIK6R:>:H==<5;6<T7Z+e:g
^_J0.3^#R)c>Z1Z8^4KSFRb)2I.:@U2_W)Z[RO19O>[_9SNFa=7(Q-g7T+WH:.LT
H,[e;Q5]W9X>[/MTbeU[DXV2H>fCGGc#S8W)VLAFfD7FN^?<&O\K9A5P_AJANf(=
AP0-IL80:Tc6;:+<O8e9NC&Z7gN=,agP/1J]UAL-^8E]4OUd79Igg[@H3L,7?(4)
WDU<]&;d)BE09>(#1Ha8R22=2\L)Ib+d/[FZJS-,4,VPANYIadC3gJEP.#UGb?LT
UF7A\^T#bST8#VC[66Jgc68aMcKcA3\cI7S0cICO5+T1SRK/N_O^:WML1c1G=PO.
\:TWF+_5JY_M(C:9&Ya[4F-]gC#&8#VTcc/Qe-2[(T3Y.\:WK;D?/geCF)@8cOZG
<@2gFaB5^3KOU1bSGJf52c>&[P?C^L0I)3#H870TX5D7J;BV03gX9MB>(Y)WM<(?
,G:2Gd:EWY-_a5<-WC5#AZ_AEKI,Sg[,4cVC\5QGX]d9f:WLI:A6Nd+FX#&.+#?;
X+G/B/^OE\DDa,a3DNRPd)10BCQ,>HPB-6&UNVb:@E-+cZ<4C811)\2-;G8K//a]
<P-^U?GH[]gX+,:ACfc>K10\M5VcdMfC,RBa)2fV(\CaFUN\CeZZBM/M6B&D8ZS>
/N_^46X5809<VU/Y?:IPUXG0CA9;@V(,QJ.8#3,L4,cOM(Zgf)D)(P+_(4>T)FH.
.X8d>?2OFX2WE8BdgbDH6>[ab(9:.0W?6N,=bIIQfX#W]<L</M?Cc]#EO&0g8U;,
UD1SH?E3Z97dX>He-fP-RV:3H@Kc=KCZMP#C)YM&<^efY+CR=ZX2fDVb\1(NQ8CH
&AK&Rc;BO-Y<X,0aKcLPO#C]W#E2C;fBSb4b6CYfL5K^YZU4P<5(4=QGIA33:[19
6R&;IK73TXT(=7S;3]?\<aY+KX8X.1;^)aCQ7C/cO_g,S/CS:#\)?=+d[]7]b9(R
[\;&6E=e)/g5[@\0BAaL.)J:0_)K9V1=PEBdX[O93=EM:e5MQ=&5=(f\_[S[L?UV
eS;OU(#f^dA.a+;5HM&@_4&K]+6[5A1S:/g8@Q^N?e;M>EK3X6[=B+D2aQ2fG,1H
eAP9HVQ7,;_T[4TgdZQI4A\?COE-2aC/9RdMTFg8ILU2-KJ&CAg3:SFM<P\[]Q=6
\[:YAg)W/YG,H@<&_WW2Q&=GA+FHGe_OZI1eA5@6YX_/_\I+GBaN:G/eEFgIabN+
#If4E7[FaIBDZ+@VKLV/S8-eM9XDXI&AY_,[=N[f)d-Ba(^YY:#J?DTC]eL<TZ1V
+G#^##F)1fb?7,5)[C\Q:/A.R+O9<2\]b2cABXDZG7P>65^gVI4cd)?08OHMRJU=
WL4;SG0F,.C)3U[69ACQ>:7VePT-6J)/-&YZ&Qd7UIW>\CSdO7dC>(^9>eS;b?TK
BKKENG+aXKH<655=4?L#2eO+,G1BT6E-235QA;549b1T=DFRZSRR]W.\QTKC:@cT
XC9f=?>gGN+30[]2M/8]D/2TCQU-TX]aY4a?HDT1D#19Y)8M==:aWC2JPVIW1gXe
gEd[fIPX:g5DQM_D8]1@PLHN2):LNH?3B38SQ6W?I6f5[MO3VXUX8=_>Vf7&^V(3
K+I]V[:\^Ra4V\5:8\A8a8IIL_:[+NC]GKQb2Q[?b1<9\W6E_NBX[LNY<<X2gE>G
PVcXWH&Bf\H\WB#R+g(:[>12IY#1g/:BTR@O0+KbJG2AVRF)B&?&b(OSD.b8B8S.
50aG&R-^MA.3:8/RT\Ef(.eY9Ud+6^KC4+IZfUPF;KI8;DIV1[GS:#XdE?EH]e=P
;2N_]M<^G5LKW,8[TEPBdRV?BL[@RI.T#E9DY^d>#g=#(:Q+@GeV_0c282?<N?9)
\D(&bg>3NB_b=0a#6Zf57R9P_Pe_ZIO41(+V8ONb_JX:aeYH(C,65E/(7G,DeNX0
\/30KT\J-36/Yd+I^I\c4_=DKeJgEF8IC8L)YeR:)@@_CZN-eccMbOXGbH2N?#=1
Zb4VG:I#<EY,?Y\Y-E?1,0gKa</U^)L@-7f_cZ\<;]a_HcdBLN9P9<<6W=0UW:)N
>[ZY_cN.@GG-B1aE(]HB+:fWe:@)Fc,LI.fLKS<BIH0A:V53a\)0YW1<VVU-fX6d
Y/&-?,3=3PFW-+CU,0BDa2Bb^5<K<&_f3(6fb2PNZAUM-?M6N:&gNMEc,G)XfeEX
SE27]E#;Cg:f<Ub>+_-/MF4Z7M@@.EF#BGR1KGf7S5@FH_GMc=;=R;^J5+I?8N)J
06:<?56Q#4:QeTAB:YDc<[eTKJT(G>3_+fQ.0]O)b-#(a=KNTf\9BDO1^(dJ?@J5
dPUQ?C3.F.9R2a-Z<OePW5;7SQ7=(b2-I3e9?+9\WCL,FHgB]\G2U:HG16-08c<e
aEcLRZ(E.TPDMV?:RQPD6IP+bXH1+0&NL948O1?96YbWULb)9/L39&<)\Bc3LS]?
.VM^@?P8Z]3_^Je,=VJSHZ&G#9b3c@dW#R7OfO#2G@^G1Z]NF8J^4HK2C/aUT4\O
4F-Pg/5ZY])1@(LESR@F8Ug/@.#RC[,Rg5-Q-E_;cLD]>NJ\a3O5ZbI/D.^]bEMF
KM/,Y5H+5TFaPTa^I-AON=9g#+GY_8g3MeUJA14eWFF:Qf02VU39C#_/LJU.)c]4
KZ9:9C;;G6We#Je=23TM86Nc--.Oe>/?eM81>JJNTVUI;RXM;g,]N(Xa6)FY6dAD
#<R6E#SEMD^MX/GP6]8@f,\42?eOI^R_0<=)V/Q8P9Z-LfbE6TJP::&\fQ;>_:7;
0F^X-85:O<I7VLA1<,J3deV26-.T43aC;.UK6cPY;dW,d4VHG3NU+Y,D.@>I]B>L
:fPHL,E7be)I9O4Ta7A]-\C?8I,C=KdX#fLcSf9:E,5fCP=+20(+LU=OH<6DS+<U
0)ZO(J/3UM29.5&=1H+3#G.9HR:3[b<_A5YLa:50?,EVU,7K^>VW.&ES_.,a3Q/A
L6fGXWIHAILF/e5a6ZY34GIKAMEcWK2d&;]cB[@.A7RQd8[Y4gdL:_XK9;HcKSND
^RH)/+MIPM;(FITUVX9_8,D2+be05-VT4W[^4-1]Kgg+CY>Bd8FS?bC)-LgX<@^/
K^+>RCN9e@-Z1?G^B7Bf75J)?41(08cRNdg>:;#R.H^cdT&W3#,&)Q/#Y\P:K+[G
Na/9RVXZ6ZGU4ae9/96I=80&7\?.A=cR^#O0f3ee.=&A7)Sd0CA?,[^b1gMN.C=/
@9;:+]UIZVf[43R?&ZUaSY;W8S]Q=31+9ICFTI3PFAEGRCKIN2A::))8b+E=<2>b
6RKM<I&0#R),,1,K_YAXUP=L_4RgGT+VYTbGY22R,K)B&T7I]2(-0+@I9F6))b_f
MK4[3]2M-&/?]0cT+Zg7/b(H3H#.Z-FIO87ANcI/HHQ[+[7,f1A;-ae#FXQE=ZDF
Vda5g8A]QcNN?P87_T^P=bB7dI7dXf?J3Ma0CVH5UQ4?B36#GZ/W9=Dc1Ic82YD?
a[[Me[^ONUI;^=E&&[^-JS3N;^&+05QS=HZ(M0f[0]>_JKd(]=-DYfDK,MZ[+0a=
?5ZfRK2CI7E=TYaEH,IMA0g,;1<X@965?UC#34X@HO62QKS31/7UEd+F\)3MSB^K
Y(XE764ZQ]YfM)(SS1H437BE&9(NU2JXR6T3V&@;AC(d6VgJScR1W5@DL-gM6fd]
4YNA:B;BK@Y,-(NP=#Ta0dQ,1-?Tg70@5;<-U40I<Z5f>XE3T3_SEM;M8J373\?C
<CX=FIDI;@/J5BJ<=XXd,FcbX(5RYZ&B(Pb+P@aTRRLUEb#;.U2-\RD9\_UZ\MFY
Me0LeZaP^8O>4TXf&:ZIS+1TE3.E?)W?:gCg2J\(+<T\.5QWG-7N2)FAIFgW&(MU
0F_a:eYBZN4gX[M1?F2MQg&)4F:N\7.:Oe&#8:QR^9FWOb&EUA>C4+NGXHE>8M+?
=K<R]dRB5.H,aF8OP]C?4aGWC.3Z7KJ:eNAC5fgg,]5YG>ISf@7L0=5EbCCPHe]S
Ae8;,/6BGbBc_@/NJ55M.CZFT@5L<9#2..VJ<YcPT09L,0Hd-E8=TX&FN-?AYCXT
NS4SK4.\T/L@=2AQXgX#)G860VBVdV^\cX1(>VP?>0(B.<N,9KY)UZQ.0bD3a6Ra
\c<N6gXb^8SJD71ETHJf[:E67-:C=DdfYVM-Q7cYKC/#A\]f:?M(1#;/2YgCLa^8
fSUeMcF95&[2@=_S7OO7cMNQ0&:5E^,-Teg6\#)P--?/@+97E3&Q[=[7?8:-7R]H
2X>SO:+P>Ca@@?1HGW/W[b&^6Y(e._4#c>@eURFUaAP2-<_:QfgZdS<bB2E1(@5G
++<_aYbL9?23=11?6Sc@g<?ga=d?NeEYN)Za,_N,B]bL#2gX)Ee[2FfSA<[Q963F
eAAV^4bd1NJP]f@]O?PRfU#Ub7bE(4D.@0OW982QCI8e.Wg.Ec3:?)0@+J,)CLC+
&M2E92QM2I_QS-TH]72RdFY[g4<UQa^aX-_P](UT5DTPFR\N&,baTB_#R1,B\8?7
_<//L<f-SbTTfged.)(BN0VSGF)M#0#eB4HbNX-gP0//H,C<R1c9&E87Z=GQ_?<H
B?#_;.SC/1aMF\0\Z?4+UI&J<#E&M>?V_]_5N\L6(H@[V^TF<,1313WfeN,QYCIc
91-JH#9\a4fAO/WN6S?f;PD./Ja;#gY>>&I+TB/>]@.g=+6/FP;LG_KfcX+D>4]C
b5d6ZCE^I-<HD46\2MUBU62/V.P9^0.EGPZGf:DY-?@?JAUcA?M/aB-LPW+>:/2A
6K3<SN=UeEUb?ZJ);R.KA+AM);86/JQ@Z1W4b#9[,?A4?f\@UFX+Sg0WNg(Q_4Z;
/Le;dP159M?&BEJ_<-&^c6VZe+5<c)a(a27B.V2LW=X=+3\:G>/Q4,+>,g019af0
AF=g8R5;a6Y0a+\3H.I]deVKGA.35:gM8QP?1.HR:L&Y,7WA2K67NG^Q_d_))R-^
CU)G4Fc</VQJ=(2GIg:KJGQDPS_ac?I=W+WOe8_G?TYN8F5-)(N88JX)NQR@#f5A
GGBYFMC#2;[T&aVF:BFH<-NSOUB^A<K4:E[;S0E6O5NV?I#f#)S4-+2ZW<ZRUM_Q
JTX/dCdFH;/0(,8>ObdKXDD@>U74HN:&E-a7?]@)XRY8)]-CBBHA7gIN528Ae>c_
Z9#g1]D,Y7JHdI&AFRADHgP,R](6\53SI+Uc@16ZW7_FJL=PM^YY0RU.2X:cdR+e
L@ZFabLUX3\7e\K[eB&a;AN0YA3G?7Y9?E-F.&ZZH^7FIB:_EI)T7gR4480H]ceR
H[#[0AGe)>eII6SVC3W)K:=Dfc<\^&EUWSR#./-KV,E]/Va\2+K>1;d@(gM^VJ;D
ZG1]VU[@Q+V033f53?Nf8P3=+a@K?acKTW^Q?3<eE(OATag@BEE6d:IVQ46d[F_B
&\b9Zf[d,2X6+V:Vg(SFG4?\_DVfA>873&1[(4c1bR(T0TZN;EK1@7.XgDa-XGgZ
L;MNK8=\2Z60fY>G=--C))5-45.LQ2^Y&1?QK;LIXB6^W36=]ATF.Q^NK\H2U,HW
,Y.B,G(XTUYXAC8,>UD?MaV[O.SfA3Ve(.1HHaGA4@d7E.ZAY?9U&?,5E\WdcG+;
^#[]]9gS\>D:#G3G^b(9MWL+V0,79bNI<(DBD\CDa\&E/XQ(>9J:EMa>/fHb9LSX
Q>OXBVKPGbC3@^BQQe:(N?&/C7I\6))#_UPAIFTN^eJfJ/aV-F@:cIN9JScW;5BF
PH4LadD(UCMJMZ=2\\fO-54Ma4;_RA]IDK+0F+A4RCTO@HMLa^[H>[?RB7Lf38ST
;_6N2<#7+Z^0&;R#gV5aTGR^b#+39g_b>MZ&PEbg?GM)L+)_3K(.6HgEK><[<Kc\
&:3ZK;&E;0L3DXb(?MLd<I^>B]X=VGf5#H[ccINCJ+63VLVY4RYD<F)FQ;1d&(G>
;K4Rd5Hg.MP[d-gAg=3f5L2Y^TH#0_[65\07&X2P5QO3N7@R-PC+T:<J7^4fdZYR
.@(#U)#f/,Z.;]@C3;IUY^/fMPFf@#=2?&bT#9:74[dJX?L_>S04EWd@IKIc?(+\
9&.S>,Z[cB@]U8XF?7@E6Q70SYDC2C-RR59S9>Hf<DB=H_FE\YZN[ZBYR,2)NLXB
+bI#8=P?DbbKT+-gX31-UN&1H0I.e#b\UY@UV7]&=Me10S0I9eM\-a]f^29(:50g
@N<A\#/.PQ2;SCb4Z9N+FQ_U,a82g^E]R9=a:fONY/#RF<;62PQI]^BE1Ve;0eJ?
/7S]4TGJY5CN8K,_,0#gX)CZf2M)gG+fOFU?]a,-V5a>/T-BEC@@]BZ^/.Eda2U;
FWA&\ZRM8d2g+WHGYDPf;IX6A#eDN#CEdK@A0)=dFLDJ2RgVSa[8ML+EV1UZ_U/A
8]#G>bgaFR]ELY8=\GDN[1J\;L2KT_Z:EcLRD6=X=:QGf3)?\9ABS0EN5EY4<,;b
bBQ&.H-c^A1BSQP_ZPb=@^>Uc3VfVcO;d.dP2ITR#<E&W.#>+C;f,a4Y\SRP8++d
O+F55:T,@=KJ0aaGZQg2>,&@[+^OMT+42]U\fH((^\4XgB16P74UADHY6BHg,W;L
@+[V0,4ad>DXQ936@B(X913TQ@L0+,_13\@cSaFY].JHQaHJ.>N2UUH:&##ZX9.L
:?]=N?YI:fO1C\WC[A^2+>WB&K:D/]6IJDV>EKTf?>LA:;NPXSD]TfC[b:>#Q6(D
8@[eR[GSg5]Y&U&Ee?TUDc]BMOU[F-ZeIADJV8#NRPO)@H#X2X-#Ad#f9FBX5f6c
#fR@GD[a2FOY@[Ja_fdGc7FBQaZQ&.RMZF<W)Ia(5G=O1:Z\TG6SI4?D8\WABHX@
,FTa19P\8/(R6ac#eHF4?N25Y&;K_M()/[GV-\[NU&J@5M]eBad:@8059G,4879M
e^NN:89aLdA8SF_[#-_[g?CSX@e.34b8_K&,SebgV#5B;T2PfPN=VE)5)3&HOddJ
@NZRd._KHYZ\092?BBA8eG-<X(@5]VD-\,])K.43LW2@8+)IP4TBNNb6<fI,0DbV
9(Y14]\.CWDQG0?gYeV2U4Z+&\,g2g.8A](KFE8#a.aM95>@U[/E]U98_M5R5Oe_
HYa_U?7&GZ+OS=;AeVCX>/ZaJ7+17a^6aGOLH[P/:.T4_ZX-J)[[^1aFWbdd:4YQ
A):7O-=P];KMNK_=L>1RcFVB/,e76P>T\S;TaOSNe/CYJ;P_#3[PGLbc[H/(9)Je
(<6)a:[@LbU]II<F)C/:=R)NQD.++U_.K[8]EXb--a<#@YfT#0,cY^)G8BOHOBX3
4UF>A6DW5V30EQf)4Q&@cHCJ.gA,U>)_@5\CfI\J=@S.Xa&/2CQQSa&BO)[IU6?<
;2cWX++(H02R(eI>L)]M21/_+F-HGJ04)dQJ]^4K2XIBEL)FD@CHPA0V;ORZbVDe
.X,.,9NN>=>>T5TMUUB_;G13/#^MY2.(ASgGF:;1E_S,g6F>A65\)U_[;fS+16H)
_20>I\#E(_T9?)O3(1?LfEQbT#L&C_#L3K(67/@&T5(+3+/_\<Y,P+X^18a2U=##
a4BBA0+]ON-/AUCW/?4[Nce,\9WOJ:RV,]=#9@B(b(JPeB]]4=J24R=V;;cf)??M
.g?dZ.WcJ3Y+ET#c?+TZ>^cXaKefUR6V1+6&dWT&AbM)N+egD(:5_9@Ze,RK0G@3
OUO=5AON?0eI<]:8_T\cP@&Y@H7]PZR,J)+41&\;eU@0+bHWDYES7._5>=8Jc1?+
KE=4V-+Ha+AT[f0HW^0=_LM87aPD1-C7A8?Q,a4MUD1P6XB;&7MCR-8R5Q<PM5>.
6&;cfE^CHPN+0AS<+Za0316@S/M5<g/6.d(9[DgR&[]GG0a0J7>Y]c6NKFY&eg@B
#b=4J?#<BZOIEaFIKV^fFMM/6A=5)O;.U=9,J,&SC0.F.a@-IF(_LVT-+-5dKf?/
<]68b9(U?#=)JJ1B;75SNL(a#Q&EC&b=/K@_S2?ESXeNOT#JM6Mad]K9L:0#[Vb&
-S0)Z=/UcK@e/Z2g;)IM\T5:faTD#9@Fd)ee+c4NL)dE:99^P(;XdfU>(OA2M)YE
eJ(^aH:b9.CZ94/fHT/<ZdF3S^,U=X:H/AH,678-,S)YXJ+5#gg7.:4(<7bV<./V
C60,PTD@b50G@F,1T502)[K6U6b73>S[I10^4#L]0f55U#\50eaOR<(POF4>4>Q4
PQ\U]U2O3O=+)?.)X=ZZ2,O<cNF\=;C(?DVa/GC)gN#EXS:I)/K@gT\cIAL@S@^@
9-IMTfBST)MIAU:]XSWc.SGda40_:C7Q#d^>#>WY)U_7D#MSc@]//4@b5DWA3[;=
_8@Wa4[2F,C#EAg#QP9]WZ,<:.OPXd1[S972[93Y;8P&J,Q#5AI[KUEPEXcN&-F)
69e9?];]4=2C.3TVK0a/6_ZS>gVK^5)=XL4WfIFB?L92QgT;fb>_=S#g<6f>-(,-
.X3[XX36\e#0[eIGKaD_?)c(?H<:(_A.fR7<Y+3c969VIe)UfX/#5Y,A@>N6AU]N
#\XJ@T<Ge_JCA?Z5^bd[X38<05dd]SQRDG,AV:)2aC<)fJ9>93XeU<>V5U345g^/
RYOH^2^[RM&EH#aO:S>CWB_57T?Zd:DAJXGZ8.ACd:T;/<,,bB?/2d:NeTQ=8NbR
3#?=7e6=;.c<LC0DM,TI/:J74d5/DPaO.R?;;7g6+fcXX>@3g&25><W3&4Id4d/g
?]O70aS6G0f:Z:SMT].Q[9JVd>&\4(;A;-_WI/V+C5a6cRY+I&9A-<#SLbb=T@LI
1UGb<^\Cb]AgG:DNMH0#PV8ag](:#)f]]edUE97dUSU-3L7e6)BQB_A?dJ+BN+D[
3&8)E9[9X2946Fc>ROFQMU^\70#]J_:ZWNMH>8\Z44FBR>_d=/DS#\3;X-\U5-9C
QN81+&[4QO5fLCLGA9-KA]13d/.TH<A&+ba&G-9U58LP66=?V_Uc]U3K(JFXKa\+
N:59+b2gJSZI8IaP\Ba2?BA<#d8//d0_TP.-FG=b83H?1c^d0&&M&;dRW86@922c
&L8DP.c79B(3\.G?\Q<>07&65J6ZbeTg9,6fb7^,#POfMaC/aRP]:b]fT0>/De1O
J7PW3-BCT^2K=PPU?gRIZd8=H.C:7B4CY^?7.FN/g@P<>1d4YRN9N:G_BHdUa4TF
a0KZ_6D>KB-P:+e)VeX.<@O]C>4^7P@9;f8PY\?I@\R/5:N5(N.-Z@#HEC8@c<44
RWSeJVIBD_+6d=,M,G_G^NbVBBVe0>GAA;Q8+P:4;]:4C4&fE<:MB2.(6E0Fe1.O
SAS)NdR7MN=TM9M@-Z#:1K7,;(H=(Q2C4IZaC=-S,=JAd0b#:\GE9>JRc68bQ-Gc
4_G(g0]gHKW3A>cV:;)=YF0,A[+Z^]Td+/3>E>7Hb/<Z<3CW<@6&0UC_A#H8I_N)
HQE>DNN(.YRFXS6fNDZM^9PP.?^<?#gB]@4K_<1_D@,JQ[ZFUI.;250Z:1]9HLAN
Ld<I11N0YI/]fP<aTH/TMM/5b8:#J/Xbf3Z/9WAF0Uf5C@.23ALK42B(C\gOZbf4
&=QB<:aMWRH<[GLFgINgXZ6a:.M)O;a^g1V@1?^MHAT]80Xe3O-TJUS<g+)H_/8@
]IOR?AIICLEZN)@aBQ5f_;XRKJ)gZU4WX2R4(O/^PXe0L5F\cV2fQ[Gd#JaBE4.J
f>T,8X-D\Q1e=V\PBYf06+=RBGaO3a92gEH)_e.Q(BXaacUO.EZ>,aX>A?2?gG_G
@?_KY=#6900[X6=U[GLM:AG^@2_=c?8e,-CR[/fTcb(S(>;<D+>d[-G/0&@M^Kf?
[;^+X6W@YWSFHVbY;-)+OT8?LCWOVOC0RE3CIJT)OS(d=:\NDQTd,UBO4S:(GBR@
HfN6<E74aF;cgFKe5JgNb[+ACT@,c?N,+ebd1AfYY>,Gg?7fMA]Ed&d-]RZCe3>&
;f_O-_XL9;0SOg&?Df81X3][L7HO#OT;>@T=HaM9BN;?_F9F(^_/CNHOFHeSWF6H
a(I[VQY7I?#DeM[d@fRba:<^UXeLU@]0X8X@O.:3_S(:I]V@7&=4\[_aQJZg6=ER
.3U>[WKDd;bT6VgcRMa)6)AOB7-C0VXR0.?V=&afafB/a[[:aB+G6^DNOU0bER0,
Mf6JU1A4e@X;=M#4L>==].ZK.bgCO6A#,V6Og,@gfW=RAS@15QILOH]?:#-<cG:B
X-&G)NSVQF<2;>S1D9CDF0aVeZReKVXM2Vb_K]3A^ffH9GEGP(_ef:c\MCFVTcJc
^7=;:D;B.3?Cb>e^0Ag^b)RAb4cHB/[c(4d\HA::DHG,R<@-NV4H<HB>;6g9-&>2
0J0JQH(&Q0TgL0cdb9RfIa=/3Rc2W@K0(ZPXMCO/96:CH8C=SW]N<PbB#^D)1Y>P
^RV]NA(N9&/E9Qd=GI_4Se,3HCTQS#HGTE[EB7N2MU5SbF5Je#K/_R;(D8>,=CWQ
SO5&Y5@87g7G5>1UPPQ>CMGa1f=7^K^Z@@cC>[7>4bEMe5?-:ZF3X51)SVQaG(?-
.f4&B&[KgIS4C]N-@(0>#T^PNT[27E5&7:QUHVaO],S7P8d.A[\/VO/KJE]=I-G-
bK_:d9L\a?;OdM>@V<aY]gEQ/;FJ0gV\(Kff(N+UIRdOXcJ_DJCL9]PEM+J7N,Y:
BPTJS#6NBHGgYeY@f@1HE71YQ3K+g=\Y;[WgAESHX4ag22U.?dV9Z-+V=&)1e,,H
OPca9X5)3MPe;B&X/D.UeRH7]f1&4P04H57:/>b#VAfK-02UY\Xa6R&<.=c2[&(+
C2YUPWDY1?48-_9Fb<Ag>I,Wg+0Hf<[</3]:7^#(QKU3S]BW>b9=EX=V1EI6:1H:
LNT]=9J.cRW]NR)ZJW6DF]CA.[CaC)7PZ[BFW&.-e9)I1WE-/TF(VZ;J=SK):KUJ
PcN0N]SP)?II/2?1^I7c\_K#TONY1J@#(C?,BEF/+N]5SXIDA5@_)Q4d7a6>f+GO
cVYZ[>,B@CdbX2_51(S/K)\IG<(M@Q7_#;AXEAbC\,R]AdG14f952/(,@75\1IP2
dbRU&1d]::@FWgg[;83:>eW-CM.&)N]Qg_IE@#8VY\WRQINQBb^6fLYIZN/SE@f0
aNE;Ug-@c>)1@/N1HA1Lf9ANaBX?O_L,@V(DGU_L;9H5ENbV&@]]0@CKTY@g5[3J
:2,,8C<c)Q)fV2RA+a>[ZJ#OM/)(E2+\fTNFG5F?R]6&9+DY7P:L;>2,-A[\H61,
FC#MZe2.NWJ-6T&G\25V3+Cg3O9IJ-<_X]W-TUd^?^9S-,+fGc\#F83ZfbgHFKB7
62#W<\[4JeHIVRTPOFe8NKf-:Eeg\:65YSGJ8X,/6b,Ac/,WS<(R;.O@:(6b0JN5
7B/B#RTF_CX^XC&.;.00<_)cT]>4DMMd<PED4SDVA4JBOK.4R.+U;O0Q)EaKIdP_
#6UJSJUAU#gT14U[CDc//YW4fMTH22W?T)5VXG23CW2NZRe9^(](38MF#c54=?>D
(?gNZZB))<13/J>0?Md56Y5FJVeCaB3-G1C=cgFL]:MX9Y_fUb>[e#93g0DGN=[Y
WdbORfK[(WINDe7SXZQ40eYT0=1&03XN8-)-]CHcLKDG_BT;+;.+9CA0gP0fRIEY
?MZ[G)/6?7/d];FIE-H#@D9:A>Tb)f1RbQ;::-gaQab>Qe_:Z-;BTHgaIK?\,e(f
_[ee<\X(H6=I49_6EJfKZ=U.d#KR844L<D>M^c:T&^IH.EXQ[/L+#fXCJL8.01\e
_3U9<SJeG3EG8:(Bb)(XIM0eb\HK_UUdN@ZeaCV6XfHH[7e6\<\?6K6W?eOa9ge]
=+AQ77+6Va^LQ,AH6G=#]Sb/BL])/BRLZ@CXF.OJ\XZ)&d8@;bX28@72Vb;T_6c=
=/0)7E_Y@cLGb57eXaaOS=CG@GQB.2/_,:AegZ??+D8bG?5/ca;7b.X2/BV]LGIF
gJMEJ^4f\L+A6QZ]FLB8Qg&V[65:,-)(GH)5B#H]KVT)OGc0\d?+KEf[><U>)fUA
^Wb9CC?F+c83d(9K1DP[KVYO_>HXdM/^Ie4ARb5^BW:>@O05@R63>IWQ4NN@AcUE
K<d)I?GH>\)?#^LOaC_OIM#B2)QOZ@WB@+Z.cT8V)47(40/3?dOLWdbQ12SP\YB+
[,2VO+1ONcbB8dOg>)C93_]8A6g^>S@Og,MOLQMW^;&UG5NMM^e1K)GZ2K?]30[B
g^M3G&12VWOE&A]_R,:>\Yc5C0)7DQbUfS5W#?5D?#Kg/;?D.QKJG<@A.@A@QLXF
DI#-U-6RIA8GaV<Pg7]BEd9J4G^1@GdP?N0]RIX65C.1cFC:##C=AJH4\E-=bc^G
+=70fD2I,;^_QEJ8:M+)@=[]G9eLL?#T03S;a.Ic6Bf^)C[O-[Vg8F-aDI@?YPF0
RB)6ZL==dDTI0U--<<F?ODe([R##KaS.^K9>033HeH8;-OK3MBC8+b36gA6;#&4E
f9<7=?3fSY-,JG1Q-M/SN(+gJ8c7J02QV_,K8.(cR;Lc6.E3-]]KU0Q)=[_==QcH
5NX/.G<-JPN_?Y7XNcINb+4H(&.W)3;GK6/gKD9AUBCOf;)(_DLJF6Kg->BB?9B\
bcde4M<+-cR?6++1\4N9d.3SA:V)f.H=/3L9TR2K(R#F(5]G-KX./1+.3:ZAI6V#
@)Y1.b28P[FN3Q5KKG@/5F.C\R>b[3CC;;_[K3Z&V,Q0^c)b=XR0F;ZGZ[5X0XHS
3V6Q?IS5O-LWd+VIf;^6WWTF;PO,Lf_:XY8;YFBX02XDY>+G[DI[;,[DZ9>)@K[L
]ZM=-aAfLc+/J&[aPG\BA?7>546?3_C]PC9Ag5HVJ;G44]7G6ec4+R_JJ057bTcI
\C<b4)]+DJ:M?@]L7559[JF-HZE\VEQ+Q52?K,J)>K.RTM/S1-Y-F44^,L5@\M)B
dJOC(-?ES6WU(4RA8>gY;2B<Ge?I0-/3AW87D2CJ/HXFM9K5TEDe+BR3HO2.2L7E
[_/5&LeS?(cX,EEN#,H#/?Tbd0cF=:T=B:>aL=V+8SE^1BL\3;d#^I35Y#)U6gb<
T\ZPg&D@?<)]LX]Y+17FRbZWbg>f>:V,d\Z^KHE&>:QWH8KOFXP/c>?:]UM<M/XK
VF(d4G+aC+=H_4TG^A=D.B(d.0_L)LD4fadC1@9NININBgTR^^U+1S<+LF3#Hd#\
J,<IQ:S]<X?)J18.g?95aXB5.JQOaKS0MP=AF\e_O_FNR&^Z41FJ,3N^36/HGUC<
U9FTdPE87NJOBP_WBOee0OTN,=g6]E>@E;>0a,M5\>#)2HeV>Z-]1OK6CaeTSbWY
WY2L@?Sa:Z:VT0V__+=fLMA,TT(1SSPI_@>L,ZFPg\Vb2+Z&JQ1,&f.9V(E2L,1#
f/\-&RU0NY[AVd>SgAZU9@ILO]6U?@[Y)KMP4Y+K4<e]]#C,UXR>];@6Y=g]+3ca
K:&HCBB(9]FITY7Q7N0a_g5A+1DE?Y77(ISV5TP6G^gC5<?fI/=]Me0-8c@1.#HO
EK>2?M-R&L<&gRA?L[gWO@XQ=U]YAg.S(CV0@XPcb(WbbgDP/,-U(P68Tgb3NCQE
RZ86=^b_6d4a5P_/g;?_5B3M79,7E;NE6XA32R,^E0I-3dL58,K(cO/Cf()QRO[#
P)bN7?U<_H1@<>V/Ve-9/B:g.F[&A,V3Q02#]]g?U#-EH76<gU]S-\WL?U-TWA;C
I)5=VZ3?H;f1:c>[8L?3CLP@dSTX-AJ]7Z12;ML\-dgcU)_?Kc5X-8JB&E/&UX_H
4cSD(^?AD;8Z:7O::V8DFZIUA:3c2Q-c[36==(b>6f<;_P\AGfa2F5^]ELW)cT>^
A_+(]&,SSE@M5_6GaWXbb).3(DT]U[Q3G\+I#AXIa\<4KL1Ud>K-d_ac/OJ>.?a[
71^dQ0P?6gP20CYa=Q(-b]X.7BB]Cde58LWF#)IQ0ZA/@.7W/CMd5;U8,+8-9^>7
7T/280+LA[@cLQHCOAMX[5VJ\57?(f+,O_FNG50db:(WEc(O+<8&HI/3F7[#ND8[
FF(VQ2N^SDY7^([43VXcWFDOSNJY:M;gEQK3DZcfT=d_4&C63S-6O;TQb\HUfBKO
SZ6_cKcR[60Eda0P@Q,4B]YDafP[+O=\Q,:KVS\IXX-4A#H9/EEb^?CF+@[Gc1V7
B/^#J#EA3,V79>=;DL)YL1>R2A5OD;L3EZ7Z-@;HNZX5FJ6O.2;ZgAGASTF-XbJI
8B/8[PZd[AEFVT&7T4eP177J0OY.(E&;1^XV#\NV^d>3fWG+bW]-c:f\T8SeFg>;
@@eZf7M,T9-CaP1UF]Z-XOQQX?UKNI2deI<FXM:W+,c@K7Q8,0BK7@]0+.:]29@]
MJ840S[#W.fS(UYMLGbSN4O-I[)\V:2=(/J)A0@I@^bW.Zcd=1W/Y187Sg.5-V3Q
0=#?HWKNT3/]WOX&W8U8WTXT&)Z>(1E(6P/;Ua/QUeVIe78VVEZEGMU43XRIIL2A
ZeHbK:RSHL5.G.F5]H/B-c5CVQ/MTR6IK+5T4,1A3f]=K+G1FUAE0d+_41\8@>7f
^a//74:0&b<c.Z.R6aA6+C+AU3CaP7G(-FOHZ4-P\TLe85V:ZHe-Z?7SCS@,_X-D
VQ1H.013Y1XFY_UddUH&W_-fSdSGB@&[A]B(.EXPD<.D[Y_Z>2WBNQIR=Q/9D<0]
8Y+Wf(d5HW&WZ>[;GBeQ:OZQZ_U1676S.X(b9:2fd0L5+=6/gU,OR6(8S3dU:[KF
:XERb(M@<6b(c)g418(d7H:JM-VGA4[?fI<ec7[PY_U4MO-;Red2HX<V&a/51)SN
HM[75eRN^LaZ)eJ^XQg,LU5+faH:cC/;0?.H4FQW-?26M[HG9ID5g9N?:SY[VLMZ
@66Zb)Q=:Db7>RMXe/Q-LL8.Dd(50VB@:Z8RdEd7DZSeHG+XN0J^&+S+RW^G9Xa,
G:C+5Tc5Q,CLe#_YgfW-b2dO0]#IV;=/Z[&:O.[4d,2L3YS;(3,U,d1ENGQ\BG1d
bZKX,AP+5@9I)g0H6Z.]]1:dJ5>4GJRaEL#LLJMJ)bW@:]0<XF[NQ5<PMcd-U^WI
0_?<\9d6U0TJRWeQ2e=:9b5@B.gY4^#@Z</;]g>YQ2c#7\BJL8JE7?EH]+-g#DO[
UAXS(T-IQN8E@Hc^CVRKFM&a6f5IJT/bI+NJd/I3UR62=9LS?A_-86B9b1GD=d3.
B5G22/:-ERVI7A;6Ke?6MF81L/Pd,0=HS6587ZYEH39LUVe1.HUZRc,b[8@S,/>b
Vd&?4N;S?_87OGL<D-;B>gE0Z].d^5<:TOM>Mg+#+QK-2:3dFcfV2KFLK<@L5U-#
5YaOeU&QTZdT>X,MK.29<JOMAF6,=O;5<SQW;[F)S=UT01f4^EK06A)&CPN-4b&Z
//P5J^J1XHZXFYQ&,E?;LY37dd51TMd39]1aX1,F;8ZI;Ub)5AG^O\Y4+#KH_bI,
3AeIgg(]9_H)K]1X-Q?f)L7JBfYDBb;:5S5R6BO([+#X6JOPQ;S?ZWf<:cb_:7#b
=Q9^<M,+NBU<>JW+UH4V^N@S+;Xd5R0ZNH9#;=@Ba7>aJXPZAgF8[?)TF[-MQSX@
]GDE-,E+69#Kc]UZK.J71.FLXMGKRS3((J-Zd(L;WV]b,CF^d;UT4EQKeVORXfJf
BUYa5^cc)-Me.^ScS/0L^.;gNK-2HVRZWf;A#eU40a>YYYXEe2;))JCfE3-S,,,7
7,e://<Md.P]d3P&a1Z1--4d--;DH9<aHG#-D:/2>TO1U#F0ZV@\)5KBEgD:7.Y(
R&F<OG+JCG<-^T/X<:BL=3?U1^gULfecXdCE?;/11-[>?-X0ECH2(WcQ4XBSgDCH
6ZG@WBF[TU8ARC-VSKZAGd)<RIT&f/5(3H(8RP<-<[P:=WaFdeA5T+_YSPe^O;<J
;ZOdQSLW(_>\<HGO2>QaVP4&_3bdFObBcb89EG\(8@U,O[JRTSI.R04UfY)dHDE]
#gDYGb^_8:[MdBf_W4MSV;VCC9Te)V-#QSK81+SCa>YcV_d-b9GGDK@,<NQOZ,BD
G>2Kc-/CB@&cLLLf-_fXPOYUeI?WZDO;OG:1=)<BdT#L4A9&E&a0RaP>W)gEeEZc
/b0ff=I=Y]?=V)0ET6Q4DNX@VD1[[BYM459-fR7.d(cH4=CBGf?:eZGd5\-&?V5@
G/+gLa6FU;>]O/C1I4LM_JLgSIE4--XWYT24AA)U^BP+&MH0H+47e+36e[&Gb(/5
1OTM@L-Fe33#e@Z>?<;f<G<ccbKCKI<03Z[33G9b_@B4T^/@3Q91:Rc^+K,D(L-N
d@Y,#eNS;cP6Tg-00f8)#=9Y6_C75M?N,L53;:>R(Jf(bH_T3c;>8..;8(5Z.0LE
;g1Y]ZGEQX_<5Fc^3#A]dPO<UcFQbVGd_VN?3SSQ<)-PM:g869#95SI7e0CSC(]f
2R)EaS\Q3XCWfD7>JD:ag=G3A&)RJ?V8,-b.A(c?Ua-cMWZdZ95J[J_+dF[,T>3D
DQM1/8;?V0WV_(Y+;E;A&^X73F\?)QUN8]H=]2:N1^X9f=EJ(CZ7,?M#Qd7TO>.U
\>cTVV4\:@e=@_S9[]ff0GV#35g^CVd2?A(;YY0DY5;\LAI2g5F3G5M1<e359)2T
/;RLQBX]d?0&g3+)YI:6\Jbdd,Xg[QR-Dg\b+OaNV/]]OT_\9H_9FXO6]@3IWAJ?
C:4GEDLf&<7PecSQ0gSMP-f5_;P.;eVF/FFITgabST//=T^(;S6+e4T[&c:Pd7NI
<N5/dOTF-9Yb&.E#+c+A<N@1)1:)&<-RW6(#EVLVK4/f\O:3f.>?RIcBT(d^H[CF
981;8;VCY_b:_FCN5301=J6Ve1&RWU)6)NCd)CV&c7c)3.1630+RM?KGN]8ga(IK
Zd0f7Z84^-N=#T/Hd[e&S]NOZ&1faGHNP0;SNZbWf9:#IAbI5EaE>K3JP>J=6?W;
TVW9c8F?f3;@4<[-g7D_c;X1V6QKN:8#,+P72B/=IgTH6HK^/DKB1U&dFgTb8EVU
OH&9<\C+P+3b>N_?[5I^Ua?AQZY6b,Z@D[+)85>7W,EKd9LCO.SdR[.e@ZP;<U+b
+b:Q+0DI,J50GcR9740)X:ZV>Y^K/H1EC03M6_be?/IH7Z;-T:.=:UIJ2+1CP-Sa
J34)f2&=<GU-JbH]Z=Ug?;@VN<M_:4[DZ.&:(5eK9T#R<_T@/T5ISa?f1gaCV1P#
R47]Ja@8N3(F;8K-7/UU-EKG/WA#VW+HS+JDC))IbC2aUQL\d78geDfV&b>[V@/B
;[3g^JK]6Lg,<eKJO?45527CST^MF+GI3g&PeZ8LcT>(=10;3;-1Z7d.PQ/@]2-.
Ie@-9=5XT&@AgGgB?R/gSH+QJV54g77Q\8)1@5O_RI8M,L;Vc@=K2dK8\VI].^6\
>&H>7d9H/81dg3KPa&aR_TFR_e8W4d0)bC879ZRTW8VLW9F:X=16[2Fcf)_/MO5(
g?[DO/QP8#JQB^cg)/CgeM@UB_cBZaQ-V#^T=7=CIBF;B0)[4T+d0dJg/Ob+:3&1
\Tce/?7Vg@QGOUaL)Zb9eIBeU9LT8DYd)E_MEgR1Xd)MB&;\Y9HfcMCK2T2316@9
SQ3+=0-^>@&d^dLM#M](G];-?XBIbMM9:.[9GTPgR8\8IgJM>Cd<5].96aB,R5aJ
PJ2e.\_eH-XJ)(R0f@9V@L6AUCY+_:25X:GV,;ObXQ6@[NHGM>DgB@FJ-+GEF2MM
N?=_9:KKW\XQ3DB5bc?CQR3/T:&,C6&B=ggedU;MI(>eR+AZSK&?[G#^@V/0--EH
TSSgFR6G2O(gEOFQP=f:#?e[J<;=<Efd@6D2T6:5I3WZJfSY;[/8Y(:)FZfS-U3c
#?,J5#gLYE0&#S):32J>9&QQ0eP5)dXJ=#d,,:Lb#,E08<E9E6O#UJT#Vc32.cR3
bI[.Z:54CFOW#;&Jf.\Z&TKX\1H0V8((f3CY-3&A6g-\EG--F3c@\_/JS?&cU;fF
>P]b1TN+THbHH165Y4gI+C\E[F9/SJOgV3c7&2.0YJ-R:].1dgB)]dc\9>OPda=;
8LUJC2ZUM/MaeMdB)Q[BU=\EB_c2RZcAcS<(JD/\XcDZ4R:K])9]?2e74-.d_-8@
T?e&N5<DfZDf]=P48?fYF&.L,a)K.PYZ/VR;4N.+?I73QM6X)Y^WR(R85Q.QUUL&
<<TC)KI0D1-I1&.,<7Z\0;7-S4E6d0S7)-@_B9^Xd8BUCUA8W0UF,YS@(&2Ga;O#
;)23ILMbL_#MO[>QCfOPTRO#<ROYLN;4G:OE#+d/&f[Z_J(]G>aM.\)2S)/B(FXd
T=<=W()fML<#PHd2VaQN,;ZSC>JP\7NCbbLc7a<WS>FM?[NQO((SRDd3ZR+(@&3<
ePNOSPYIL=f7?&\=PR#Vgf1P/NHE8RS=:;]Cf[JeL#/b&K=9H^\@Hd#@7..Q2?GO
U^I2+T+SBM;K.6R8WU+]>&B41_:CQ[P2.VV:TU5Zb@K=_/HIO/#-25.)M,U2^J>3
1[LXa8NTeY<0O/FfM<99R^)TgZ8Kc6dO#UVDb4F:&8fH>gO<IR-We&4)5@YJ:;JM
IM+<b-e\DF+3M8ECKF@X1^F_F@9PR/TK3X2a0@[Ya,Y@Z;2^.c(0HU7,:1^aV;,)
^BS),>L@T5G-6gO+@(^L7TLZE>I[X;ZRf/eK,_AXZR+=Q3+F3W&Zg7B)eLK@B:+_
TAZGKAH4g/FHWfN5X[CS8Ya__3<9R;\d.OHTO+YWGfNB@D@&U@[ZQ0S/d4Je@cJ)
W.6MEV2<(=R^(<8N:Aa1VaJ.\GP/TYK,=GASIRgd61^E]<6Z81&\8DfZQQ)4=X]I
/+\A0<C8\IXZeTRR^8(XZf[]BLS.-a?Ib?c?Ub@0.=g&QM@9X&.69e;R@188Qcb9
LOADKEaV\_90<[C5^QQ]gA=U3cFRNZ/-C+EMd#)cS&4/HKVfH^YdDI498WAW+A3A
F@b.MT<.[ZT24\C9=8?2OA;(&8LT1.4HATA767OZ&6/_^<N[\:7#NL5Q=-^,]Me.
65-F_)[Y5@X85<0>N5.KaJKL5SG>1K62b8?QL?1O:)4dNTa8D=P6(:>9_c+8&aCW
2@g7\3e(A?9ZA#eL[I<B]X1d;&9bM:?_+@&YCRMZJI+OI?a6Y60V\Mg1[+7RAK8]
/EJU-U,J\]YdfJ4aN1EQ>]DeC^-A04f4a/3Yd5Ag=BBX154CLQJCHd[&3X)Hc\@C
[#fL//#W#U24LE\/UO]I<JP-V>3Ncc.MI.g#;KP#NJ=b:)B68b71ZNJV/cca]e))
?)@<aZgJX4aGGbJf5AM58/FKOBOdc<CI,_/V_)[D7PCLA[2SX@B0L@WJ1E>4V?DT
^b)d1K@K&YS)X&CdRP0aA1Tg&]=3B=B7?)/45bKJPH?A/@&fAH,8XYOHV1Q;4WcW
^89JaX)>:PIGCMS8GT@BU:[d@.g^R[YT[S1>:_<RSMd.HM,:S&-dR1-[<^5V9KA=
]Td_+V2bN9F4+R&@&=7gB_VX3,;/S^fP7.JYeO1E6(@JI676fX[cYKfdFFZ7e+#7
IN\(M;\L@ZD\7+&_XWP;<3^,gXHNA#VVQNXa5eaK9<MP:-H=AJ3RA/>)\LXIZ8(&
Ta&#82:+eV^,[)8R##[LV_I8]5a[9IZ[DTO)LQD?a7cLQYOdFNKI(/JDI]V)&0&G
L&P8?FFS^SP>ONfYWC&<>HCLMN_\OJHe:=/Y\eQWLYMN3TYR^T(E-+7fMNA4Q>._
F0NIQDC@T>\g:ePQ\S4H328<P]D62aY5g93<g-YU)UU7N_SI;G2S+ES^3=;RX;=N
Q<Y;10G9Y&T)3)(QF,(9@SDNXV+T=A1@DUU4UR/I3@&B(ZgE__GKO6X]O[de.W^c
(OSNPQ__]<:61f.E1K)[&]R2^F6F1XJgdVHg9?)H=Y<7<gEH,T5e_<\NDN_85X08
>-\5P/gL.K)J&VPeIW>4_3BW3Z@E#@(a\(b;/>TCIE#SHPKbR@Ug[#f31WQ:.__1
ga_[/W6^7J/O@Q&#g&NX7D6cJS;UP-6-DH?QZdV2RC)F+=&S=_GF)f<G080_6YI6
;4/T>I0Q4Q[\;XdCcd,M^<b6IU(]d<#^:6b&6VbV^LYMJJV^0Oe9Og5474_f_Le.
O)QM8.fceXWP(M</KH;a;&M[_@;40NVCX<\@9KU:GA:7b^M]eGDc=\RKf,?P+KS^
^HWHQ=N@&2F\^0?b(16E<0gC2-TL;>^@fOS04e00^V&J9I.3K-@W3)c#J4R6G7b0
(3;AD9=5AW.JD,@G,Q;2#+a=G->Y5eD]>RD6FMF1Q)@X]/.7][cM5TaG#[D_>Y,0
fd103<?,:RJDAd&@eNDPRR.EWfJYcDSB[MR;W+.(D:CUVaeXK7JRf2P9/@QdL]FQ
U>M<]W]R>F]5((RaVZPD+UG\ZGA?O40e:LG@YbeV:K?3]a]_f+PL2OCB2N8XFe0>
>YU9GM>L&[.0e,e[T3-Y_?2WE0B7PMC9gf^G^/DHfL]YUf_O>3AJ\0Gg.93-?<K>
XTV:/O&/>D3;2\a72/E(FQZ,5.XWA7)^R&c,/8=f@4#=-(c-R#d<5WA6-7Ua]9I+
Y5:F?9Ef<:I(fce6E=)(>/dcXEf+=E^TU:,PCE8D7Y-0gBg6;2OJEaMAg3=]8N56
UdcELO1#-NU=1]88+c8,g(V]WXWK.Gf.13?Y:2&OJd9X^g&WGU7/J13]E)\D2X^[
X<NYF2Ed+\b8<g/d=Q]DeHZ(.)<]LYL?CV&GKF4F1HaFRZY;#;QCcUP4FV[ZVQ_c
Z/Q;>-[(0C4^8/([T=<5.LeTVNE5_QK?DP0HCOJ=8RE_IJg_EHH-V1=A&A@7##/G
W]PTQ.+;:YVf=3Q18./Nb<0e)UE:YLIX+X,dbd@f(f0PKJ1SK>#X)Zd]&?XI(;<&
Z:\9D:@P&K(0gTA4Pb:19&1N7?XAG[B[6U.8>fA4cOR34:g)0:W??YM]9L]0=.MS
;1H-B+Ta+FP9PWV7KIa+:B\NeI:8QE>/fB82#PT0/9B:ZVJIbR,((#U2PaH[7bOf
8Z@37N\cfU9J2^#S5OTNA<.4I)C/fe]g4MH\^\F]^Y@b.(8AT[9J<,b8P(]:AZOL
4[]S0ZF[fH,,+(\17d/W-d^:_1JN6HHIf?9g?DU\>4e4Z]f,\;(:J3WgR3;1Yd+R
SOgZ,f(+3aSC8;=Za6RV0^[N?:P2dIIM&:),CJfXPMgdZ<Gb3Qab_LBFR?MH1UIe
:O_&Dgf>\.e#1FVSR6GB:&DBC=Y_5B+9G=P\@=fd^M50:]L0Me]V.FG4:.a5Tg56
6NKeYF27f:2_ST5EeWG@Hc:0@\Ub#P80gN_:JCd=)Fb?E8@+Y5F]S/b786RHKB/C
\Y?0-gCLKP>gfPP]D]IU?T[RB/582g#BSXB,=@#AY,0@f]_N<UC@4d</0U=(ZSLR
0Q/-e?/Ce?/9<\&7O><2,,9X+0V/]_]+O)a3_@-AC]=_bEcfZ@4K4J+H,6VL//.C
=&?M3\/),N&P5>CZgg6eQ(#YS&^[#TD>2,^8U:b@/Xc8.65Z?364ZA.a&(Q4fIAY
D]dQ8A,T>FBBP-TS0R0.#^U4)#ZIX;HO&JO?.M/C)<fdMEEG+<.-D;B,@,#gX\>[
@1Ea7XRG#CG(AA.^ZFNW@CJ-3S?8V&e]KCG@dNNI]:.(^I.dVTAP\KD<E#UJF_&I
S8OIJg)Q33edJTdMSBHVDdG((+e72C(aC>X0b6dM3P2,K:1g]CSDcb:fZ_@3E8C#
cNQd79c(CD@6-+=Ta-?T<D(a1&D^L#g<b5E:XEN?L75413@L\_=SB.7Pa#a+<N)N
VX7]VB_0CR=?FGVP3H[V>9^EV];.LTN;VJP3/KM(L5G016aLL#2MW>>g[Q+eNdg.
,?S.b1QcV5BHS#?YI./O&K;3J=RX3Y10AC<OPQ8^S4Y1YbK=27#^6aV5LY\-8cdJ
/\5+Y&MI(ST0OKVEU88V-M+\J)7LC#:1PMQ=K4c\#N2#_(D4f+Y20OOT;ce>V-/Q
^HI5FR31CQec?<BJ4^KK@=DEg:T)8f-PObe8]JRH.ZS:+4HM1I4O4HT.?M7AfCA[
.,TUR+;0,A-;FK_K7+e6fVJRUUF/T>)f3YcTRdM-OOMFYNb1c_U=U4PNWAW9>YLH
,@cc(K3^Y1.+VX>aCOLdQe\1S@KL8QdbYN3O<J@F3UdUP2dNeB]KUV:[-(BAH/-c
N8_-Q1_4E(KHN[\S&0(;>fb7DHZRXQPU00,QU<PS\?HbG\g:A,0d_:#b.#_QOVcW
5Y-],gMB):H->?W6d_8#@S#KMF)A<7KVLT(];\>Q0Z4b/5VXSZ,/\KfL69)UE#19
/NOaSF_I4dQAY_]YDOEe^4N5]H2_X#7BcA3C@PaWU9O&5HSMM-JdN?N>:V?2U:HD
1c\<7^\FW/SJNGc)1fAGKeXY]cTCHGa8X(Y#6X,fRS6RX98a<F:L0L2BB3=A&_ZY
&QJc4<_?X4c/=]AKNSBHS>D034@._S(NKMP+SYDcZdA0?(U_ZVI]R3P?8b9/D^(/
IQYM7[77-3N1B69NceQ7SA48?Gc4-=[TK.HJ(U-b8aZOGHZ3/&60:f6@0+?O;FEQ
S\abD,Z5a4dFB[H:BAE&.:@+/a_[Rf4O./H6/d5:,7Q/.BJad>_X<2_dA.27LQ?(
H8B=4@.^0f]8&,gEB#5bQ;?gYeS[I>2(4[<=:J)1&5cS#e=NNU6VRRMc<=I^?&&N
Q,21?5?VQ9T8=f,RS3B;MA;.Ee>4,3:_=2ed^KGO;F>6ER<AZ5-UPP[;]R^Y+OF:
,<c@Q)(01Zed8R6\C\6eUI/5Be/AN/@gDZ0.7X6PQ:b\10R_.</)@0Y#8WH>aD#Z
9Be&H7>X@)CRB^SCd5AXd>M6)VLcB+:TX@Me5@4/3K/Na[CJIN>KWLT31:>9AUcU
N.:JIGRP-.1KTbeDL)=IT>:5_Oc>1)NZ+RL-+1(JRYUC-WWFCe;9;U1=dMO?\[VD
358]JS2CPV2+45P.(aUK79\\>UNFEG^g^N)O5^PR.?,[DgXQ6Fb:Oa-/BVJ#b]E0
27&5XF<bVD+?a>5LaP_RB\ZOVc-W4<U+R2M4FV#/9),&Ye&]Z50?R45?5XI)dO92
4D9/b683DJZ9@;0BSH,2JQC/._/TbQ/A]_RRRX[K4@<H1==([D(#Z/FG74b5=:=C
\2E0?].a#SW:fSI?_FQQD8:6]OXG0d4Ae3Q<[JQB[.7WaN7F:7##)[_bd80f>g+,
Q@;R>0;Cd+CUR_#.E;@b(8(DHHe:-Q:aE6G>Je/Xf?#4D9E8(b0]HK3-7IO=EW1&
baJ8FPLf&&M@NSQ(KSLT28?;\6QfS9?0YE&T20N=]YI?/U-B27XDb2-IO+MMcAT+
TE=YW7W7\1NKQ6S6:#WgFHOV3^e3LP(BdRVP1N3J+:9+7_#5@+bB(c@2/D6b@a7P
Ie7e#5UQJK-gF&?<5V-S5;L05ZUYg/&X9:b3H&c8KW0YL?Q0]1:32Z;0T?C:6[QO
/+2V5>Q:2.^0P3Y5O+^M;SDPQ0F)0f;aPGU(^97PaJ>?eaK[@M-#P[WV.HXdeOf>
[.Ccfd+A@B9M5(<E9/J<[/dIJ1[1A\X1eTdUK4[\Q,.)6,K2a6eUF2(3b9J0(?Nb
3-,3)I2,/B.=644KQ[);DLCTKgd^.aS67TQ2VU5:YH8@I[]aW:V04Gb@KH[XT=O4
[@Y<@d_]-3d&&V=U[_.:W1N.JaXKUR0F;XB(KdC(Z97e:8\)X.?XbKEQXF4c0c(_
J:SaUR&;Ja[B>P497#7OT9M[+S^+_9D19S\\[.F8,M5&VZ?M?>Pa:GDdgaOAWI#T
ce((Y_4/FGd&:_R..fT/EAVVKL=6e6RYTKL-^I3VBKKaMR-FOVWBUdF:+f]XUHU)
XRTN.)MN;-edRN#-7C.e-?M[ZA\P8+Z<9fX12Oc+WDa55CZb+.(+;LT]9DC:PfCN
?R+S<P[eI\L/,5VaaL/89Tg49f,M>4E]O^,c1GO^)^8[1dL9^KC=_K\G@&M/e8dW
S4R40:_/KaSa]VY><fN]E94;R.LUe;L_/HbDV\)A)=:97AMJ2V&@Jc9ReGfKP_NG
U.D]E:-X/SQ<],>PK-TM3W;@;bL.?R_[^Gd7MaGOfW4T#3LH>S[UYR;-:[)e&0+L
ZWY:#9KeQHZ>G<X16a\8K_@Qd6K)QYd@Z\?6M&0\Q7dA[OZ]UO=GMg[dK)L>@)T4
1cO,_+Q8b+&bIAB.1]^>&e)\5ZPG8=Z7+3Q/WUgd@K&HP9.R4SV?;IRHTB<^/9(-
BC\BS=+6Z;<g>-;=f^OLg@G;DL58X>R:^Q_)(G+4UbY#gHR-C=E4I^7)]M\9_>[Z
]1,:2_,dcIUUK49A^0A/G25>[8(P2TLR9GZ(_2MP-Q<G<<@F571<6J]^5Z4<[-](
,[OS<O(Q]\&#YS^,@<J2-T&K#[4W/>Bf?IgEYNZW;<.,-)OF?e_#/C(G/Y^gX/8?
><FWNJceZ8HU.^K1g56;]HQV;]_,J:)#;-AVP>QMc_&RNH(^<08((E0+?X6G@geG
e)H[#\-dX^ZR0TJg&WZ;BgbHd;:a+4YM7<1H71g=(,:XdFUSOY]]037G@f4II=9N
gIL\O:X?.e5RK=/S<78G:26_7P3=ZE0J.O97b1QcFb@KEK-ZCO0fSAS/TUI9]ONI
[W1.1&:[]K_cJ6RN2JaKO#8L\B645ZOU\MF3-/7SWNV?4\2<1;+@O6#@:(2SFIC\
>cd7-X-3J6d7BBS3I8.3-_PTK<cNC5T6ZE(&>0Ff(Y,gAS6XB-;d44M@e4ET\QR9
=Mc8^IU\09E]09S=NZ^GC6c5<QY5/f8\3HLG?L0[(LM;JLf_9WFfWOT,Q^W:./91
&-2R5GR_(U6W.0=US\Q(T\&S:H[J;)D]R-LOfI6<SJgaUgMMc^a,1WQE-Yb()@K5
0HWN+d#6EG0D&=Gd5Y(;IYZE0XM4WC&]d]X6JP3X8faX>IBe&5WWVQ\8F+R[.LBI
MD@S]9(K3IT_H6>42AS3V@\CM40I4PX#4M0_38b>@WeH2EBC,#?DXN?=V?E9VN?J
aO#9JSD?dOcf49G(GPa@[.Wa[5>W(G>2fQV[D35]+O/Bf93E:Wg>+(:Y^@-77-]D
;)eR5^;<,-37^YW=E]96DZ7JUN8RJXV6KY8[_^_IAPRP^CH2K1?WR=CReCdQ:5HI
W(B@3EQMO]2R,NSDWTRNI=:P.c\TNOQIeQ83.?I5TW&1<,BMAND4:g7F@c][\gYT
I+8BLDX)+;g>_A_Zf^fc#;+1FYF5?H134WeKFXR9U[MV6Q\_2+bLMGL3bUZP9gZA
0e7,Xc,FP)bY(bJ>KN,LB/#Gg-d.S.E(/_R#9.AG6/?]^[QF/KBUO];H#Q>NE@M5
WI.P<Q(:7#b3c#O<W)R_0CSIH_E9[;+F;=gVPYfW^P,ZeB.cGC(F+cG&ZUXN&5R7
X^A@9bAYU,06=f\<E)6JEB]g;X0f<>2D5-H1D_B]HbdB3JL#fedKf.+-^^BSVP][
^6^-)[_a0NKJP>9?2]?W(H1_IH#,Mf6e.T^XPe>J3?ANOF<+8/Lb>Y.MXZ/c.Kdb
#T;,[@A1U?(;SHJ+Dc]WPc\;SJAT+K3[SF?OPE+HN(G<GbV8B8HTQV0-b1UcU\O7
7PE(G^READEa89cGJR+\,0;c&.LGab3YEdUCa\B#7UId9@]/a^FJe.c?:c9FdPIT
]F=S6g4.I(7dNNHS,,QO(#V@/^8_8L\&).O8;^Dd:GQ\NdF3A)\A#8c/W7J./ZW_
N/K,^c(J4]W84>?<a]<L[/Lg47gG_2<MVJ[?6C\a,bdL14P2?A>NR22714-HY,5;
J@3de5?P]W&T9B:JH5<DfGJ^.B6P1&_\.<2RY#N/JI=bV]XdL(\Nb1VH[7+GM=b@
e(E:I;NKA#/_+Qe03)55(RY[+06ZG\@5&)EAYH,a@E]P_\0QKUaMXX+91RT<[0B2
HeXZOJ]OO,W3A<(/fV]_,?]5)WX1gPFeQ:_,?-793[Tg,Yc(+PcGJJc\IBgP&=H0
PR=H11I8eaKK92+0eAX1)d#Z7VLAEE6#:Ff\5-^BJ?<<P=H,2=92@9L[T+W^,ZP(
TX>3?-4JaA_8@P__TU9AJ)_OG0bF;2aIc_M.3P)9_NCE<=gcTC>DdcU>1WegX6&:
H]eY):DfGXXg)M+N48Zd;d^7cCAHf/g6eMKHHE.U2@S,+4R<1:(A@bb)e@3&;SP?
X+Hfg_g5^F-24e+MLWQVG0=AeL\AC8W2ZB-f+,CC5)AO?^e^Ug2+JHX+D=WHJe5/
_J5V:X8(dK.).^8<DcU;8U.82W_dCa/W]C<@(R:K+NM>TaMJNg2M6M6+(T^.90HH
bFb],Fcee.VV57P4PDN@O2b<FZbFIU0IQ,JCL3@[O@AOSCfQQ=AE8X/6&1R=N,7C
=PeO+-e(112+LUf:-#3dC)CA\U:FfF9BM>e4b)C]XL+#BBJJ,]USOR0&N\<D+RFR
(f(+c]gS+06.2XdE:6J_EfL8^/P7b,>,0bIa)EOT1gY4.&JME;\PY3]/fHf5Lf.Y
H]OMRD5VM&O1+QQ^a8JE=NQ+]@QB5bCY28J/[?LE;Yf<[_E(PO(G;1<WIcADCRC1
E^,Z)aRZ/>QSQ:a#H5P@5c/dW5PG7:#@.#c7^I_Ig?S1N3CU#)b_0[W)_ZYTGSE5
,;@(XU2b50[5<1Y9[ATQ]@DSD[-7-X@EVGd8-d3Q&8T^)T,)1#F-Y42G1Q:^<c:5
V8N270YLCOaSTaO1-0,=#dcX])_#>\.62<NG0f3L(PX?M<)JOR-=V[T9G^d#Lb+8
(#5gKP^\HV)RTNHgPJf#T\/M^\fTFNMDAb@+^?C5&gZUaSD8\)_P]=e(\_&D7I>C
^&]EE&MXX)W35_=A1W35?SIZgg#QYG3W>BRXSP-)D[6>C-R?.0>>[#>P]A+J3O?J
Wa//-D_QKTa:2,0)56&3SB:eTe;O8-EU+ScNg/PgL2P:AX_L>.)K=;5W0dAY1-MU
H5]U&@EZ.Ja]G8A.57U.Z[&&^&f;7(D+<37UO<Z>Q5L3^Q>a=J,R5#13A<caP+^D
\IO^O8SKF?#2T<\1,OcIXU<<CW81=a.]HU=?^1DP5#MeYN-4/B8-AUVb<U9?=,Ng
,?P/#c[P;&5JDIg6CQ/bN3JG1L=#?V4cO2L(a=OT.AFA,N:1)0?=AebUD4W?f@D&
.c/(/TT6gIZgd@/-A41JSfaP=([@Da]7PUQ^NVQ0VU&FLC]GQ+2O;6D&JSd]^=3g
_g)A/45R]W8c:5VG&_@=JX/=OJ6(\ED&7S0D=.=Y](P9L5M82c/W#^_UY:],[,:8
@C>-AO7>f2KY#EN97Tb-NY.BM_J6T13Nc[O01HUO&)c.1e(aGOCU.S4DNH>Fg6.(
.R+#K\-FNR<>F>A=0f-^3a(:>OA9Q8^0_gNWd--S-UNC2ABO9^C.^4L&e<>\6VcO
&_;bM(W2P:+MLg5919eZ5(6-V7V=K3f@dg58D9b/,Z^#6K]\?(,a;XLbYE<.^WK<
E]gQ--T6PE;:JNI0&OPN3R()EG7KTB=4(3PK:+>G?Sb#7bF1[P4[[2[^aA7gK53S
4[](^DQ(G-^aZI[^EG=Da>;JE4VDU5)GaST6Fb]6L:[U;<5]>&Xc=-P;T)KdUS++
@PAf[#6HBcL#1)3e9?V,KAOLQM#X1W(ZW1@1RCDd8SF/#NB3R2gV=\?^(T:&#L\c
1CeSVQAAC+NgBU,E=d]WOHT.1EKdG4J\f6H/<H1_].QV>QU;f,2dB1/B&D3P5X7g
=34+>@P[>b.bP0A>Rbe9ZcTC^X\X]D886;Y/6dFC31?Z?4g6[=Me?bMZdYKfSCfZ
<5B><I0_=?1:256cJDUA;[;c.g4ebCYW(g48ee75,Y4IOPB?QWZ61KBKZBG<<A]L
&YM21-)G0cDTXda:WgaK52]B7-ZEU[N[U8<[aW1c.BKcBZ<a[99^c--&<>SO9e^C
#1KQ(dAHTNDU8C18eXaAN-YJ_:g2?UD,GYa(bf00Fd;UJ9?Ze0//A/Uf.X(OR7H,
5/4LT\f8/.ZZP6WXMR/B,/YOC/Bf>=IAJAg5CR.g8J6&1+DW<EI5P7gX95_4G)J5
HVIR)A5d6DU_8RJ:bP_EBX4UTGGZFdB&D\143NV1_RWL??#>Z<:=+Oe#0TLN[HKD
Y9O&ZC)0E5APN3X#,^7PD7JfO8CO\SVKMOg;^6JO4O^1J>WEEDb]80b<1Y(1.CX&
6/Y/R[=FfbB(6-c.KDfSB2G<OP>L)@L?^E-6.1_4<:QQ?)49++f<H1I0Ac6TVa5#
+,@3f1Q<<DC6-^BEIQ<O2>YRZg>776BC.;W]8NEOQ-gNJ^b4.ae;>9H6;,/UY7Q+
dG_G/,c+b9C06e)[6M(A&T53f0+aXYYb28CV4Bg&9+a+)7I59[Rg84>/]XY;KPT.
&6aY&36e^6eBR]Y-Z@A-\(PC6FR8&-H1E\;#c81UR5fVG9&.U[\APNIZ,6N[#3CW
RcgJ_[\E?:_.(7QaUPH^a_g2Nf[<G(76?JY@O]7_5)c766,6;S98f=aU,B<KO\g.
_>=Y>S<ee5Z:_9-Ub<1M7\+^TR<I)P:+6W,F.+K=K);[a:7XR,@(?BQ9]XD7Z#d9
\Y1V&4N^-]KLQX/.]]>eL+e1C:0edCL_C8)b8[H;ERSd20.<6Sf[7[.^UD:4)N,1
[6VWXQa3.^+b8UMg^I.\+-=;W,W7<>)GYV6)\T;U5^NWOgR^\0#_IIS0fK0U(MV.
5]VN0<3:^JP8\d+SASC6gP3=;e.#J,N6L+0+SaO)?b1V6RB5W3([5;3ULQd3PcL=
/S[2XQ\De13-K>O-T;H2I&HGGZSON=Y4,dgdU+]#G7;Z#^D)/Q:d20dS4d4[K?6d
GAESB]g)B9FF+-:gU0X->d-B9;M@T(E9<IT2@gJN22f.5N?@R9WAG<eV<5<OCB,.
IMHaa653-QKV-R/93LV<#,&4.]2S-(>4EHTNCB@I?FBJ>F?Z#[=Z0BR5C@01I-Z^
(Gf=N9R=KY08\2FM^XNa_6Z66:5ReRL;T^\AR,#b0_FIL0d@f?eXT4HLeMbAD779
8\6:6f,X,_Y)cV,IHF0?EA5]cOaJF3_&>UOaZ],^11M\Kf:ZQHFfNN[cUDO3MSe5
VX248X^M(B@9@_3+:@3,eM:S/b9AO5M-0IWB:#G5+0CaFCB(6T3KQ9&J0KfYB:&;
[7_b#6QFT&>1eDJ&RZ+bDIL:6)8LQB1:d]J:f@JX9Pe[BE7<]:L]77.XDbGP(9UK
N.9+e@0\3&IN2c\OJ4-P+ORG<gUE1-J^WM@IFF-,YGN1)PSY@^4QJOOSU:/1.+b]
QEN<.b6AIG#IT8S4R0C9(98aDN@e7.eZF.d2W2AI@T56L[_Z(OY4MVf)<N4?f:L/
M]8>c_WUOT3?WW.1I_/f;MPRVW#N]Ma<+=-Z:S#Rc]P-L,;.6.)cfXVOA@>?=:=L
f2^I39LgG9eKe]Q]cB2N#VA_@HL47:a74<71I0.^T>M+0>D)L]DGZRObL,U,XMS6
e<KG1-EMPXaE6<&1f7X]a^@OAW.^X-?6[g^\V2Je3#caE0Ee5LPRGAWgX.5IG/1#
b;/>7,3@-_FaBX_#W_VB]40^4KGH6g@,eVE-+<(0^+72]8UY1U>:X8bL4a&Cf+7P
3FMW749MUW[#-Oe)L]^BS]5I^,OP@-^YHQO^VC8R-T)NU;W:-GZ0E7I^5/UGcM-C
1H\N)JKY.gQB2ASQgYJ496LS,I#cU<>^Pe9AA@WGTBb:2F[M?(C,Y-7Sg_4]cHK+
cAG8P49_H1S7g=Ng4F:0A/(-,/U151=]]QY=7aE8B=Fe&9DIZR4V0QHe,3EdAI>9
+CXGcE^DK=6A7_5.^ca2cE5,VbdTbeTb.Y6?@#=\EEaNK@:D>dBH[@<#M#>0W+WF
_#3bcV4+,CYF4\PC--#\?QZaQ#;>D=P<J>E6WG=[N#=QQKK>BE4>>S4,Y#&\6U9^
:G\9P@>>=#6&:,9cBTTOIId#7>,/&I;OVEaC_g]LYEE.&G8R/385f:ON[M^A=;IF
1XZ.:OT\G:?=F103U-)LT/g:OQ->/aLedSFI]]AA7-D?#Ob3(_=1KCI4UOWJ&9RG
]ZfG+[O1+)>dU#-0^7C7Fg[M#JFd8E8H7@>_XZBNJZLbM0EXa(W)QYZ:@HZT;OLA
E7EC);MBAM/2Le<>#<O[YI9fEb]F;NX[Wd5;X&F^RGX>8845CP[U,DMUc^:&5=FT
3Z^@@da)N3.Z&4^_WR.1d8.T,EL/R1_3C(<9=A&13d19>53FXW8T#d\d^&V&Z&KS
L1&KSZREAIHOII#@W2I#G9.825e_<df]S]UFaZXS^0LOeA0CL?#R[BU_5FRP6O>.
N-@f@aee]F2LQ[@CN-CYa\0=7DbH4/WF>b.)RZTQcAU?CM>7RF>b#N(e&PB1])D[
^SMRS^0Ce0I#_B_c2SMN72U6\(F_<K74a1P5AO=WLB)&;GV<0#gH.g:AH4e/4gQF
#_D,HPHWFFgJ2,60(TYK(6>g<D.B]EVQVKB-8gM,bOHfSQg)+I_:g.IG[V50J&;T
W;T8E5]D-NL-(F#4&2F;)C,eG&eRQBHM-3C4@SOE(d-Fa?DY.OJQ^]&=gXb@8D41
LNSWF+#b7O5BfATJULDB&8CMU<?90:8,g8,(1,/-XaGc8cO)9S@T^JQL_K\\?GKX
M]@NU9cHFF;O[I/Q/_6JZK27VEU3f8H=Z#2GE?b@=7Nb^^1gZP=c&>G571X0H#;C
d^,X^K2-L90,&W&QbS)(c1aNN&0N;A]Wf[\c;HY@40^U+FWH]6N39aDYLN0GLU/Z
<6\=47D&S:M[e[A.d/R&UaG@&:HT,C9]08+9Jfe4\(K@FOLD8g^Xg\29HK0OX5VD
_YPT4WGN7/NfJ=?U@[dR(]C1[_LU2bB/NdIVFK)3&0XN.\K]S_=1ROOC]9?AG?E\
607JbN2^7209E=EF&0RG,a:aZN/fT6NBR-SbXcK/KTfAE.VK(.)N,)08>,#&V4>J
\SaH>f];C]@JcT3YBCR=?0fI&6D5J\BPK1916UQV95-_&=3G^7bG(MDOL7D&_C</
Q9:U1R9SSgW?I:Z3ac6,g@KX4P9\,b9Kg#[P7(CaF=YB4HA.dQd,6<LH,[(]M>3.
ZM<;TKD.8-d\,+d6BA1-R(#UG.BBP-KAb-bL,2BVNG@E^K6SH6&:b\:2:RF64]WF
GLN33LF-cSTLX+T4C#ca5DfFN-^EJCe[\;?+XO2:,JD6PMG>XT@fTO9>=8_OA&b@
DA2a6O>E-M#IA#@WfO@37)LS(_c&9K_d&g@_,,I7A.&7Q,-BT+3]KeQL?&;.0?N_
@K?29T)E)Y6[WD8(f>+.WGF+G6FO+\6@[1[>HQ8C,[J;:6J_Z.^)a+:LQ8ZKgC)^
fQX//I\@@@7F-R?g(OX)QM4WZ9EDX:O_H#NELe)=20AZ&(f]>B+]DfJ35BU/>G8.
DA?B[^VC+JWT<DdF#C0#G1_B+MX]C@HH35He,b2/Qd?<ADbAJT1[U/;/.(D/WFMa
IH]+@ZN8c3a-I,J75.5EcN7):BBMI20,P4B]bb)d)AKGHZ-BD2dZCCa)d6ebg?>,
^(>Yg:3<MOD8J0Ce3OCXZB8Z@JLXHM\8@]Y:6WE.>YSaDNAf/MI#f@+e_>[g;CLI
a2>(9bPPX:N;W:<@P?I)JMSMbegeZ4263,UYKGEgfUd(Hb_HKCQM=MI3Ub^-=9TD
CKQ^^P4TRA.c^G]_KggO\Qa##2ZAZ,ZYL+6[_CO3D0R35JF_0O&D&-[QN,BI^g7:
_WQF&c8&];<40JIgSBHZJ3;K:;FL(>MGK.?0RCQMT0^WS_Q#ZSNJd>A(c<X[AM[2
,=)7O1^0N5cH_S0:I.3K\\RT6]6H^a_V>O+MZJ]T.,:64/.Q/=c>g1FfQ3eP4]WO
Q:aBa^)2C/#D)e1R#g/BORg7F7WXe-cd,8S>S][cPAOad3[W9>CDFQ,S8)9NEeID
,XIFc+=dPHSN-NeQQ;O[46ZGT6fC)/[HAN\,cT0W)S-DUba_+_5FW>gQ>BU.<6&c
U0F_5AT];<=6cBPJ[TBI+=g+^?Y<>I1d1>9K3KO07++/(+c^]8[SQ8&b;CXRVBZK
#FHgZ@eFEDaL@S6#]L?\]ba?:Mg8=CObXF5f+&/2Q/<J)7360J/6]^.e)#(O,Z2V
#3<.RMW]L9R?YAPA_b)3eMFc@=#ef6&36.^VcG334])[YU3N7INcCW7_O</(6CaV
aO-H9\FKfA>IdG,SM5?,R\I8(I.:V-VK:^DB[RW#44<g=a\@SH=O,X.@T;G1;7VE
::8ST.T#c<g^0-.KRX+7?&?UT0;&U0TaVc>F[2HQ7IGH(+_-VL[CLRFagR#R(36E
T:,UeaX/3g--4Q\NSQZU+^SAb2Y2]DA37+4]YBeI5N)Q7e?JGX3A<L5@_GLAL?G2
(bbLXgB)NF95d0\-YTPDE1FR&O(3N2:S8/Bf&fg,QX4cJWGI-+#EF1(6=4W#FSTE
DPJ>@8[5Gd6AH]VcHa<8d<JYAFFa\^J4]C_FV2-OU=dSHUW.KDS3SVY\<?S9+JMP
3F/=1BO)B_KJ47&Kg-)d7K3LBK4X^3T>_4PTe;acL@,P8GG=gPB^<CR4EV#50b,R
SNaI9C//17X:BY\E6H\D##OEJO6);6P3LN2/dAH8P:1GX(85?cNMRI)JOY.Rc4IZ
J.d>8KbfXTE[XE&Eb7g=5EMgcPE]<03bA>VM(;EeX6)G8MHF@E=^.9+(6dSO-_.L
>YDg:N_:K)))IYMf=97;KKCLK\ZRUF_K&Vc#3=f)Y15@7@bcM6O@OB>L;U31bS;5
R>J-334VY,<MMTO)18:;)_(:;8bOI:d=?42/9.9R@9?eKULC?[/;RD#=_Xe[U2HT
Sd\Ge<LgS._K<(G4a0.5_,?U^704K9GZJ[CYCOSE#/_?G+XIccLEMSTPIbJ-RK#3
P/C0.:WWS[aDB1#B^0FK6YcaD,T-:6;S1b;?:=P^X?&Qc?[G,(R4S/#TH,F,7^0B
JTEG@8C#F>X[Cg7d504#=DRNCEc):#P3+L?J)d\fBX2S55I_8c8Rfe95?7Vd?dN&
dfKS2;-=?K.Z<2Ua;M;LIE@:>L2LTda2329)=SW#7<5QF[eC+eELLS41bY&d=@b:
[#g)EK34-g8IHJ)GJCSU7Y<NLBMeTd@:CZXWRFHW2M]?BgE3L&B.e&V_B#LNWb[I
L#g\81c6.A57N#YeFG1I+Ee1F<)^FUSK#bLQSD@0#_b>9BV<5Mg5TFLI8A9/P?H[
3X6OBb^N6O2#\6Ief6UdJ3?E#1,Vaa(;Y[=ZFS#d0];[MF?e9e+KZ:./^YfBGT&#
dX4SQ]_L3)^fT=QR4S7]0b&G)e.JRZV8d_<)+@5eR#WJUbT00Ke7,LCf\<3+gf_T
@b:U4KB1.2Y8;IQ_7bRE<aLN&).&2W@MbPdL(H<K[G)E.\9;&c7;.]PRa5DCH^DM
+0[LM^JCKbaUa\-_d(2bX<eJYc(7XQT7-;V=?HX\J:4BK8Q33EYYc971>N#59S4&
\M-9P^c[T<:/\5?ZeZFC\;;_+fSb;NTG;\SA2f3:_gf&7H9R#T.K#d^5Rg:L(<6I
IN6d.B+aND+-D2Q/Ab,ea2=8=0405-+^CMf_VCZP^Z-Z=P#\C)B4Nc+()7+RaId)
Y,H2AE>-5ggeAF(cDREX@-6:TF,RRO4&SO>TeC/66LRVE@3ON;E(CHN\cXC]TRX1
_4GW1Ud&K5QcOO]+KE=IMa>#Kg2cJ^2T^]0VU-fB(>^7&<Z6F:0fP>,SXJ+/X,S^
[,HaX#N:,+f0QPeN>1)UbG9ePH,WF+b+4O+[4Nde+&5d_g;[6,N\/GA/E1D&S96C
<=8K:Z(PLWD:eB<]KJTBNZLG&###O_+HX<W:Ed/Zb<AMMUM/e3M\)eYL[WP-c:]b
_D2_?X1.e9cM)6AYQR6<1JYC6L7S)V)/:9H]P34_W+<:I9FK9GR,SWQS4;SH\gA4
=K_8_R=\X>3G,#Uca(</Me^[FHQg&Hg>\M,4]C?V^#FN_&/M.b/+&(;F@3LAAAWc
gdA78^UE8c+)X#TXa4+202]9FD#Rg2L05Wa&g4:^>OGLZC+;Z+:5-VN[AG@CL32f
:>^OPP5+a167,CNZ]a&RdMc-[\LcDY@#CHbH<)=;c/2NE7D19dA-(6U-PLU=NKPP
QD&7HL1L8?0;fc)P=_QCA5IN@@-WaBKX_URO>@-H33e66-K)UP@S^6XbXJ_7-4V0
VC5)>Z_(HTC>@-)99VM_WGP)U)VfVP6FL@FEd+E[MP;dTE95/R-(R#[\WP^0NgOQ
SN.KbCJL@-,RU-7b&(Z+CD;TMce1XP6]081UF:&86KOdFbO9W2<<Y,+:b=<#]H6^
Ob5HSTO#^GI0NK/7EJ&>d)2X&U^9J.V7PdVM\1S8G_<TTXLEW/DNV:7JH[YD?278
cMfS68f8P3[a>/9d@&]VX\8/Z(XR5e#41Ke_Q>?KY;K@0,W.N^-5Y(O1dBZW9W@B
<4V6e<7-HWZcRe7QY,NHbLgPJZZU55(dGP6@X#/9\P/T^dPHNUHRb5EM?T7F8W3<
,a,Y>Y<^=:N4UHPd0<3K3&g-9G)OI#V<)/?Q?#NEN2+Tca10+HNSC<<VM3;I]9PM
)?9T<MBMC98P;QFNb^T5]IFX&f=_Z@cS3WCI:(g)aTb@4J#\ZT?==A+45O@+T4GC
aE3;IF1RJD5TE3+aE2S-)WF8HHT_1)P;QR.fQfe7aHNQB7+=&C=/;8,U0>3+C@]F
9/LBMWS)6e9<M<]S&P>BI>HT0G:.2C;0,bRVPaTB)Zf-A_XO#,Fa2&HFc4c9?^S^
cL]_BeSf@)SNHO68R.&Y0\PA9e(6c(OY<>G:),0>6ef]-MIA[9:Sg(f/&3eT;F^7
U(f7/X1Pb/EA/G_QF.H89+].b<_EXF(K;\3O>ATWKX]#6:9d)cUW4V_S3GG:?JHO
&,17-WOe@GL?7KF>Y4M&.5GJ?[\KV2Z(<A9AF4eBQO(\N5F8e=G?S]827A&2@K+C
N33R-6Sg)b#)1J]JQX(<@?aAA:/:V6Y:=@7IQ;dHU>><&(Te8O6\=Sf:;J>O.XY_
J)Ia1X<dZW=>:/C4UKPWY#4@=>]I/05cJA7A/B4O7JUKUHIVf3&8[&#5I/<,0bV[
3[\=&0]D\V:-)Ng4@T(&462TCU3V<aGY;9TZ&M(J[]Sf?A>FUWK&S+@6<Y>W;=;I
c5TO[=8/0G,6AKS#IA2A?AK\?@[>E(FL9.H;Q6B]aQ<I);f3V2)J/Lc-<M?:11HR
OeMU=@?g(),E#Oe=gEc;KGKAN/_N\:.)9#ZQ1BD_,(9M,R/g++M-M3G+bD7IegP\
K?[KIP@Q:^AI?@=Qc_LYfa739E)9,)(dU(@.77[aA]1e[]LFE<e7T1L#3g@YXN<:
aJg_HOW)+??38e#>K5(WSYb0COWg;_;D)M6T^EE7GSY41Q+Y.0XEd=),RH#FG.3X
&@\OJ3g;T,b:(P>c&^>]4KAV]PD/4C2X]a1.J1,-aF50SZ0BB4/Rc^:e_\eSZEI[
C(;d=(2L2[S(gDY.I_#7.G6YD-+S85=a5#&R)0)U.(<##THfC-K,fg#ZAHgD[N4d
g())ZF1[/XSE&,C@5.&f[>@7WVg7A>3C6L-31T2#WbTc50;)D,/M_[4KJ+9/QV#2
YJCXL(V0b).GOUME+b_1_LgNA,O0[7CcYH.2.I4;2bK;+#,YS?aC(>UO8]L_]4=0
&4UIYIHCQ6aY\cVANX.SMA6RUMZP)YN\1VAMW2)/G3)#D+_cG3d24W0A9OVd#M^4
Ne>UL#28A-N@?eN=c)W[De-g8&X[/eT]eA0cEg)a;b3dS)/c#)L&I\aY9IOBRg]H
T9-&]R)K.,TK5TZ[MP<HML44P]<M+-C&aS4?G(:YRN-YM@;T(=dG:P&@5dG8\F_H
J.X\GSaN;NMg@\,e[@LLc@.=BP&;OB;3e?BLJ3R&3MTRY/ADR3D,c1P2VZO-+-ED
T8FG-;MB[6+7^\]5EWC#)>A1#/FQ6[L(\5&6Z^eULQM,TMW5;+4W.-<8]/U+[8MM
VPR1cMVWfd3(;-#BFDFCR-d-BQ[&TUX3X49\(BW]A9TFQ>eHEULX2<;.--a-OY)N
I,PN59=8gV[RQ[&Vb(4CSCHYQ[[&O^d0RF.]93[KdNFJgJD#/9#N1OABB1(d&AT[
V.B8M5A+?d7=[;3OdcaS?95]9N(e=:#DX]MI8RKH^<BR_a1JT;>2;(A43a?XZa0,
c46K&b<K_/B9UW7aX8C8V2_@E/&,NO#b\g(<EYQE?+X9(ZPUaI1UR>=,-YdWK\#[
c>&Z;5PAR)R]/36.8AFMWUG>FA=e&@XSfE)\D:]JW&G9_=Bg8+,R13Xbd/bdJ:R>
JbNZJ5c>&J1W-(eDO4b9b02Y^E9YXb@&M<GSS[g2V-T?+E@ZC9J3K,]]I6<A.CG)
EADRJD-d?H(L].0)/S=O.f16-2XDEG[I0?f.Q96[PMd9WBBg:4(8]WN1GOLQO<^7
g/.<g+<#Z1@aZFWLPecK@ZVY^EL\9DQMgfe01\gAI>TBFEg98.3e>WI:5Z7M8KC6
1RF@:NE^8:]3=e#Y+FK1HII8[QG[Wg(c8be[)g6>^K,b_6RGD6O^ESN>a,B-,)C/
SRGJJa#YU-]L_5-\:VfM.g^_0JMTdQQRdI(8C3BD7:RI=L>5c14#e[d>TN?70bIE
(((d5;/H]W_FfR[_UeLc_W)>K[/A\VWRNFH9Vd/R5W7+(=)T7_[C_>+1F&@a#Z]4
R=.?TP[]96P3/T9AU4O.E4/NHdGa<1a#U),S8?0g;7;)=Q&D#1<DLF^=MP)LPe)a
<EXUWSMDEaJKZDM^7.H]@UK=dGWC#e1g_<d)BH5F]VN8&7AGB&PUX1b^LUPS#++=
2N:PV-K#LZ5e6Ja;1,K;1D:+B.[;29/X^58S:O).>M)4Y^34eT(-+):N:IFaC-NU
-PUSDZ)<]OYC&+(B1.^+12_X61P8c2B)f:(E8Y42&VNgJ>@bda1#SN^-_G.9+4T&
+QB&RSGHSNdga.cI;^.KJ?7^7gYZ1B9Q[&EB47T&AJf.9d2_J^@2KN:G4YNH3->.
Bde#.WMQL;MK](?G648[1-R8eW(66W-X86d_+Q)#:&.3NdYb.O\547540ed(Ab4.
B+a6_3#a]OYCeCc2ENILJ(NFMAe.B^g0?>WA#-[:P<bX+@b6?+G,QG^B7>7Ed07;
CM,fX+59VcaW98bCOc9d;KCAQe/F,65S63V8N>D-26e,f,0K=(Lc+:,LTLaZd^^T
PK(L=L@\S>2?e1<@JR#TZc[cOBgQg&3:2T0O_>LA(E;<KW<MIFG-c:+@20dW1LQM
8Y@:8?-70AE@,,0_A<aB8:R6[c.N72bJQ[.2+U9B1/ETN1Y(;Y&8/aO6?[L#>?(:
H4<O;0d35YD=e[.<M36R#JBGK1JZW#U=FceO]df.LDJI=Z8:b<3g/B22NRfHBg\.
@61CPV@BRb/ARAW[.;Zf+cT(IGY,B,4ePBA<A^DG&TQDSMIQGLB5CB4YZHOLQL8C
6)9JaVWR#g91(B)@dS_f0;+L.ZVR_\F1BNg+d=NIUdD:;+Rg8/M+^M.N2W;Lg3c5
/03V.?ZI?=FDb5&2&Z?.23_+SDZ^J?7beg#eWP1:+Cd7#g?(eGRPeY=-)6L6YK[,
6XU]U]VXXS3.#<UZ-cW=U=LSe,#HQ06&FfAX4PP+X>US\;GWCVDB-._T:^K@9^^C
<TTcG@;:(:e5S@QRA136]fKT0a?3Z/XHW,E32=I[_T#^_,+K&\)1Y_43fZGTGT-3
LRWUL,UX7Y_?UX0@&\fFMX9L,R4T>YSW[UgZ8U7\4Ma^SX7H6(];/)VAF8(9VSQ1
bH7O_PJ<&&[\&&(F1PE;]]VBPgVYc,8X1bWNbL7fgLaeOf--#cT]?QgY^O??:5G3
;YJBDFc3b4?EJ,VbU<IgNbNe8H)OdA,:^@U,MAMGMUW)WG^fSBDEgB)[Z4Z;EC[d
GU)Fca?KP4RNA&T60Pf/0<]^/)60&7HXGKB+.3CB)3A_.=RD[2K9(T>I?b<.5_gN
..,38-0@Re;)C/[5=(K[O^8[ZQ]7)OG/a2^K5=TeKC?,F<T4L)^Rc30;GG5:\[^D
SeLQO/_DQ&Y+5PDZ6UD0EFE?&&#\8DJO>?MK&P^E\KQ&.Z(<Q[;@BS@4d@,^N:6I
1;_Fa;M].G@P^8DQO=e#,BWDb#4<RP-8Mc@X02:5KaL-8<I4e=_0e,UdR;fg/gZY
5&#7^2E.SIPD^^S:H9E9[>VVO\H++J./XgN\.\=@/S@NGPa9J&4CPAXY>)II7(IW
-ELT-RF)V<?=12YCVeTLeA]G=ICQ;H,FV0.16_6[U/[M3U=27UK)292S1.W0B)X7
[2O4Y1d8f9?ECJ22],?f:/8VR/bFC&-+cDCIg,>)3ZdM\&fJA0Z4==S\9@XB1W1J
/7QC:5R#=4cH3UX,>05N^\eQ5Q5d1(F@)464]09;_G:KU)UCC+0Ad<_e&;Y)D/]I
DeQD[&>P\-^EQcE:_I\<[RS8-VR5)C44QN,)^W@URAO-G+0<UGE>LEdcHSGc@PN5
51.AgTCUT7DO_JD0G7H5Z@4.:&FdY,]\JXO@9?)GCEZV\VETNQ::J@84+QNdFV<_
Xb^8W(/;V\;]3/73SQW<Ja[Y8d6A]T0Q_>34W-?T))#d1V\S^&&;U)[dMUEB3L&M
@4Z8#)NJG363aN]0?D:7bc/b[W9VU#P=-Sf.4)cR&N)71Y+b(6,0#:[CO:WT@-NF
ZQSd=IBG;;/Y).e2E.U(Yf=@W::.gWSX4JMRR##)ZN7edGc&bIKD]5cb=3;bZHOD
g#3J<R5gUG2C/JdcV:^EOY5W^cMZW,PZ64)\BH/KZ]E\gI&E3:4O)Q??U.Re3L@b
@Ef3V9(X[_S;@7S/6QRG+/Q=GcbdE;K9b,fdFbE4UU=W,d,0Sf4&SZJ^M#GARLL:
8.f]B_RX:61\;<)ZfGfg6b3:1/NZN;G58F8=aR&W(:TWE.Y5]8D2];^Aff]Ma/S]
C50A(+>V@SUY]:^4-\&Q_[KVM44>def>U,@E>EWF8b[4X6DQWN6V<\UJXb:LSIXD
Lf(;ed<OZ\^Z;>O3O]>ZZ2+b6[CURbG\4FdK_K:A\8_GAGT)=/JaU&V^RbVcA7Ae
.c9W=\00gef3@Z:aM+)G-LgWWC<d.aGc+2[NK^H@13=S9<?A4?2f<0N6R5.TPJ\[
10e,SEb6O/KC[<.PT_V0e^(8KFJ[)^#/&,WUc:de#0f(UU,D7:4E[YP=bEP5MBNB
UIA^H9bU/@LA=9:WP^a><J4:9>W_YOV@X7@RC:J2V.WA,_];Dc0M1Ec6TWMVIGM)
Q-88P.=SN;.<\@RABbZ<FIT^NI>-#1E9CYB)OI:FAceLTS33^9egI/KIQc6C(gc3
R2MB)@&5-5-5?/fT^HbP8X4F[TD6^DE2OJ\QCg,UG-B/SL+KJ\BGLI6Ia]cgCI7g
:]GC1:0]<4&YKbO90:)(Z_X4]84,+19V.;FEGeY_PAWP(Fea+d.JEFO=_f).A5gf
9NT)Y;:D[MaMGU<V@PNZJ>[\M[X_0(e6&/=)2B&:L3A]#A5;L<=5]ZU_?W(+55=R
J]?X=R4Zg_b4-K(N),Q0U51V+JDLa>X9[AES@GRFI:YI-J.Re#_UFDVUgJG>Z6fe
NKMcA4b2GN;M:/2=dMT@&fa)cA&[W2BTW4#QWFN@8L2NU=._+.8B>/9b6V?&UJEQ
-2ZCLP?SA+-a@P_)[(]\U08AC],aL2>G;GP]>g(GcH@V/bGd@S]4]W17Q8SI&D64
H.C9L-/e,&(a+4(RZ@-856]-Q7bWAcJ;;:59UbNWaf5AGE@J?44?+MJ9;:[FEW;b
+Z/I=(D&#9g?)<&cJ__SSXL67FB<4_,:Y;#f38PPSL-_DD?Y[)QgGIZ2BCKL=C]-
cOL0HOLN>\0Q,fd&LVMX+GVf@@4^G2A/V8@U]HI_V>J?S,8]\I12Q9(^c@,a348I
=dcB_:];IL:R+P3@Eg?/Z7e^FB04D8V[QO8T0Bd:e;QcHIEcHf,[E/U:SND_6c3R
@Q-bRb>CH.#W^5/+0.B-cZ7RfDS^_;E90?fDAX,>b&P[fJdMOVGe\J+]V+:<KV)S
g]F;LLGA.;[#,=JV;_&@@OQDGb<)NgMH&HU\4OP+;+4(1:-ZZ-&Q[(X8Z=I?NIVR
QNE0fB,UMCWaNJ@EAEbO?GSH5RgU^F,9Pega===?F8-5D[4Jf5Z@d_Z9OB@KH.T,
V_Z-L0GU0)NgKde7ANP[5[MN&6PHC9IH#0[9d@]\-YD+K533-.Z55I2I=2K[:_bZ
:WKbO&g0AHe4]eK(_.Y4A.Vb<OL#Y@.,Bg:c3,WdMD;NdJLU39),\3b?f5eFfIHc
0^S<S[Ec^_P,efB=K<V)Zc[_Y30O\g(=Z7d7D^a8NT[f-W>JR/P3GPG?cdEGA,C/
^Tc[?MDV,(059([6Y,I#.F(=4C,W0&0)QG6N.;@deD3]cNfFXLJ]-DDL:NC6@+P7
\9?gTdL(?/;6E>gKc,<(OdD]D/8LZUf,@&R#Q3FIL9YE=]dWUc8KIDaNU36dJ5SF
Tc7f5_7LT4T+N;^,N9CNC\#T2P[BK4UKES=]3\e:#C_C+41;_;U68.WLV4QC<Y]U
fUgTa>Z[_(5:K_(>]K-\.b2G+d.\I/@)RHc1c@F?EN)c+Z,e\[LBP_.,cT4+5>03
f5M8TU)M+5f8_@-?(WWCOV>2P)4+Z/>L--\a+)ea889A.BeB/2MKcHc3/BW6?<DA
EG;^eNFW&FJD6_Z[b[R^>V=[,,V;;I__#BU);SMg8+?1W5XK591eDSP]HZ8ea3TW
L^fNIC=9W(V:S)@G_WT34bJ+F>cS1T[EHQ1AR)Ud]+E3IH:_YP&;4I,SF&=B(2&c
1X>WdN^&]RHaEXc3M0^=5Ab]D/,4;J3<_7Z2;eY.S:B6X3P(=Q:#XgDCXPIU>BdZ
69^L_EU_<6D@Ya.G.:)8T_Z7]ACD[YJW/VgY1HYF5^-Z[07/0Y.Rg>?F<dYg1c<]
FPQ9O8&3550;O\7Ug?e>4DG.X187)d64C.&C3&/WbC@.Pb>)9AZM<?VMANGG0?7H
,8GG)_I@dU-<=P2Y5SU&_G0O?YLf)C/;a;I9YD0U;UCOb94J>&;WLR_gfO4#1,Ac
S3YFV?\_AMBCfSSH&LA)f(UQ8KEc1(NXYCY^e[)ZHUY&##7egTNcON;(>77P&X+W
Y_->@;aD0Eg:9[E07=+3VJ4FHb,2Ia>;WKIINVJ0_;;6f@DF,C4=g#JcbO\Qc2]^
YdWdMgc)SRS,,Z5d=7-Z_?bF5;L(:VNCT5,YT,^[PQE9GQ3[eO-g;<S;?1IIYS,V
P#(eD#&P5@OD?bU(3#g<;\BFgCNNF4f->\LGA1^<17TBOPEL,,AK-4e-D/\M@._1
6XMGW;O]LS-3;:DF)F<XI7T<-H#EF\T4MKB7)(G#Je@XbR4C:M.NXA2(R/K]I8AE
MD&TS4V[8RCQV6U_TYM-[5BBQ.9A-)9&]b2+,R8\2CKQON6--NgOV,ZJ.Sc(Z;]E
E<-1f;1edDNLS1a9MJ+QSI=Y/0fREM2.4ReYMR)fXDM,<FR20fW6+Z2EGdWT8:&T
Gc_b=O[(PBPW>?8Q=PCG@0KO_#,XZ]2X]9(TMZ)ABT6JeFRf1JUL-geMNfBROT1>
)J<cARbfb\C>bGH<[,O#8S<D7d+S?0OV&SF/VPQKTW/VL0@gf^L-\D0H&gAWT^&Q
9(=2(UXAeH8LTLXJgIRBa\VX&6\&-dCaMF>^,d,R-L<)8T0gWGZcSSad13A.E:YC
Gb,Bfe>6R41(;5W+0/@aQa^bKPO\0:=&@a)A#S?b9,T2AX<C,=2QdY7H&A1<R_1]
KOB733;99Y3<I7-,3Ma?AXW[^W63f:3+De8^?1C]J98E[#2(B?1K,;dF)@D)P6R(
RJF0?S@=1f791,82#AYDb01/Sd<7A7[dJ7PS>O::9F\N-Z_1YEf(dP++d-Cd8G[8
0>1G/JRTM2IK6>:]L^;^.5(JXM&8Y.Z:d995&]YZ?H[W-)Y[cELSe7OPeUe_18?Q
dAbAJb=b7.Y@6SWWd\=QZVVJfY3ZX\S>BM)1LWQf64J_d?#CbJDeX<@(c6_R1Z/1
bHX8T5?fc].;a@Z39SEYeOE_.SS18K4L)aV_&b,@Na_?ACTE<S/GN/MWDM>@_9H)
B8f,@S(YfL#:S:ZL/SbE3QBf85E.9bH+^_/[.,;4TM@R,M+^GCbf,UG>(W=N?d[3
#K&c6BY]V)1_5,C/CeG<+M2ZO:GBNTQTZ2>5=S11Y[=Jb2<b=Y3>+Y8&+.<5&4CA
U1fXEKV4fP-SRIcC]L.EBX8K31&UeNJN(\\[XS7WO#,KCZN#1EJJF=LKeWTG4IUO
SVGg@MKVQD?SaEg[ORd6;6T>>OfbBBBbN)9Ze?/c2R=00&W[f&U7+aXB\BV&^N._
6S^RG\IR2G9L4H8I^Y,M>L5,;\P.TcA)YX5SF&89;=RPQ,34g]:LI_GHO#eFDeWB
?HgaZJ(S.\I0_XFG0)f,+,0B3F^.,S^K+A\G<GK2?;Z&DaP:/S9PY^9ON.M]WZXD
)JIQ)^<1f;>VE@/??cOYVXG2.Ye:/5G&<<,J/a6C:A,cYUAJ[>\D59[PaJNPb\4G
<#SJ_3&?)5U/,#5X9VO[5+;OL[4=_JSf&6Z\0aB-cL0b#FTFda+:LPK]83]H>a^L
28P,=(1P]F6889=D-?UF.&=f-c^;4O@0O,/6B>G#ILW@1CBGPc<-?PDQ17>&80UD
.d@V8#XeD=:8-S[Cb5UOV<HK1a_TGa/1LV?gfL\U>:&;SO^ZV)[02LC@GYPT_8TN
?T&O<SIN,XZ6F:66fHXAJ4gVMYM3-2?[:.K2AKEA&9VPd98>[Ef?d6AN3(\.eWNO
e95^\F_1/;+JO=TWg4GA^+K4L(A,b=aeZcHT(,K=AGJ)S/[W[.+3#K\II4.HZXdD
LU.8eC(bCQ8Vd-[6Q2[0R&/=HeV)TYHFX1f4=VNZGdR2cGV(<?&9AJ)FUQWBc++R
WK^d4]T+8c@DZ(T,S<AN@JGOOVP8:_C/c1.F7OcB1UVc5O)M40.BVCZEQTN>T2Ef
82TH8NR:,gLa#L#B?^093T6_VKG;K:E62<,GB>;4VVcH[E</bM885PII?BQ3>TV.
M,.H#g3G+\0IQBfSI&-QS)bG,:6]ZDGUICR8Wg5+SWSf3V.,g2ZM109VF\SB\D_[
:[YAJ/9B\XS/MAb7N.Z].06<0f<g83:Y6=3=6L;35+@<g<EBcH/f?S?<g]?C17R<
[UCfLX7,Ea;2c9X1a5JNBZ?3b-(BcW[#bP]c?/dHFdP^]@GWf].Aeec@/_]b(d;K
):E^#<>5-]_4_C27B#1AVSa=?Y60gc#(fW<_F[cQ.U^]E?TU=[G>#:<8^c7dZ^=:
gg9>5G2D8NV1MU-6-IV8K2C8B/<PZF:H0V70KHBc0N)\RS\&,VGJLa=CKa3;6gbU
8M&dTF@/ObKYS<CU20_,H58L<NEN0c4[4=+61)?Q)ZdV/=Vaa0:Z:W\E:-:JR1?4
L&((EgCS5]^WP^0LF./;ORP396DABU8Z<+eTV(C5D;1a+P/E2/c46LbAK7DF3ZLE
O3/KI#+ZUP\@TE=-4?/(Y-4>TeU2:,I\e:KFeZ1a0#+e.EfJWM,K@K4K,P<X[eD;
N4<U(G]S+J)TQ1<DK49S/=E\[F:@/+D.>;D0&dfHa#dFAD=/-JTF-JZf.FN]PKRX
INecdNMV6O/SC>,=++=U3Z01<#RRXT/WQg33W(Q+[JKG;5(HbDKJU\)X#KLG4Sd2
M)b05KF=WeAQ=6YP<6O5_:N4Y.&:/F=]g]]1(ZX8S>P,P6JG3/EV4CZc/(P4ObCR
X0D\BR:)c68[S56EIV2a?=K>T;+9&HPadU=D;NefNF^D<4YNBZXOS-WW[g0-@Z)^
4MRJ=FA;(g?a^ZgDeCO+7WAGEP-33aC^6UR7eSFT:cW89gE?1S[U]BBNV>TG95]B
SQDEcMSF8R2+0R2]d[>A<]UXYVP.WSBN>/##=RH(I9V0DY@2BR:KDZEdBYf&.QA4
@.-#9gN?Mf6:RdfT0H[CVBG0U<]WC9>Bf,cZ=\d_ZaSa6M37(THW([N-C)bd.^bC
;TeJ<F]fU6@0@NS+V\S9&=IT7^gQU>(a\\_O3&:9W:HI(-^VWSA[bH[gJV);M4W;
YJ<FU8V+^.d>4>+O,9XLEMQG7D1NPXCM&4>J?<Ccb3WCc8QZ><NB+,>gK_432RM9
adYKH6((fFNcU7YFFf/RO-FPdC.[d]Pe^8W\<f[=a5D3B=Y^B8]V?X2I7K_#;;ba
]:QH#@GDQ-QHOY<CW:ISJUVIVY+(FH1/dTVBeI2=/V;HPe_:Ub1#;<123MQG(,HV
5-EN1>G3ALeE(6<5Z6(UU)5QeT3/^F?E5#SBX?W+P:c;g0_0acbO-W8[E\;)a4E6
MTDaMI&XZ;2&IGU).SORX?3cJOe&8C,QPff5-W&[#Q2;b-3ZI]V;(eB]BCBT.G\7
DX)3]C>eOKdF3<>8GG#e3Rg\eL5\7Za)N[^BTHA]_.4ZIOPXVcR47]CV-(T;;;I&
E5^N;c\KGC22W3QOP#PVT&BLIE:/?HD>OKB[>W6TI,0daO-HFe,XZ5Y?]_e=8Ye=
cY_+Ne&8.AS292=IWYW1]_RF-:ddRbW>]TW/gf[ec@#IYc8cZb#X9ddRcQ7^c43(
6W^&Tb7@/\>b+TVMKENP<5[Ob2EJGG@.VC@3<)#E\MI@Ma4BI(9KZHdMQ<c:G^<+
R[D(gABLQFO:3aC?:--,1+cYI=2)gW(E3aWS,XeT2K1f&f(233S]>/FJgV\M]8Q_
+-#H7139E^5PV:J,XE8,@#(O@de_WbLVa:3[+L[R49;:LV0?OAQNcL86GV3&2&4U
0+0U6;[S4_YEaP+.GL:b\UcbIL4fZS4PPW(G]45ZBB5/+<O^Y-dWa;<D)/]c)O_f
P_X/Id9;O/RBM9?@U(V_&S4/1BV_JSOZBN)VZ0dT/CefR^6b-76+-W:.d:&,JD]<
Hef2Kg\:dB#)XZP),Q+]?8DS>M00_\RGa^:M-[eAO)2XDS#91[ONJ3KO98)T#I\=
\d#f;([NF0YF<]D#6JZ4E]g.]+Fa7>?OHWgeISB77F)RM1@LIZ+74KYQ)I+C?:Tb
Bg>:YVJ[BT&8]WCba+)KM)=88=5H0\USQ-17:0@=X.MY4KbccF#R-#bNL58[gLOX
5C47//VH2.gCX2IcZW6+5(]J2&Q18V8_cK)Wfb2aBF=g67_4.ZU[JE_XAR;Hag^Q
F6Q8>ZW2QJ5AT<1F7]e;L#5g;QXbb-O+VD,^_f=ET0^39LVMJY1Q>396ba?IIWfE
e(cD<+2Y?D<QWKIF1^1GOT&ad+6GA7I.-SdO?<413+9U\7V;L7Z8a#VC:G)V&<LC
a#)LRQ(&9:d_KgIWL\+>f:daER/=MJ?9]4;21g1OP90@?<7K9e^WEQecZMDK^WSg
,:ZLVO4=6:5L_]][=5fF@gf#EP1TT1_Z[:E?W>&-FJ;-+&X/LY3[Y9QU+MWYMI::
AZN2aRG_&dF<F-&88YG7+G,&dI)AN^(S17&J:\(;bQ.3#=/](FO?DRW/aL\2dQ\6
b/M46)e8>D/HG4#00<05e#,4&>1_Q2g8\.V0@<#YO^)adW5aSQZE#XF_7K.?=.HPV$
`endprotected
  
`protected
_S4ZLU,QVN]DE00,#G8VT29&+N0+)S)aCXM>K_W7&5<YLa8H=LY<&)LLHU,\ZB5-
1CN??5D@=If8a.)\Q2<8DT9&2$
`endprotected

//vcs_lic_vip_protect 
  `protected
1OcF3W1,.6/XcU+G&e8W,dE:+?RU#Y::P>g=#1AJ;6PXJZ5W4JM<+(@ff[;5KK8R
A.<OW+#[9\JP4FSOD7^T\8MZQ?e2bJP[GL)_gbM&ZS,0;BKCW<+-N_F(8dAEJfRG
I?YP2Ff#6J=EQR#EPZgL-EQV_,50bcN&Q7K01G9)L9&RHHII1D^#1&SACCga.6RN
\R+DKYG9-TAD_>\E_QRc/c]=+RBH3[g)-D8ME3IeVbN2RBGY9Xc7ZYKBV&gaF2-M
/HNZ9C.Q\S9+a:PeNZOcU?)XP,+]V=808=_EBS,E:0.e5L#DfU+K,<Dc3VC]D_->
;)<\O8b#4fO&7)+UMOFA0f^FILDR[5@U.9cV5SIU@7,;3L#gCQIM0=e3W1Ac)T+@
ZgC,e^F:F@c(\GCB9??HME+V6Q4Z2->4adD4dI?UU0:U+FVc2^@PUg_KE+dF^2]5
TE<Re.WLZfb&gM3(,.#48-&(=>YH7&2<B-gH^?I8KKD6F\5.H4dTBCU.SV0I./KN
)JB<J1WA:HQbPXDJA8X1.HY#@#HM8Ve^YcGJ:CN.(=f2PW\2TNQPcN.\C2,TZTbT
W4N(>fbV/5,4CXaa.TWV^6DIGJb:eT-SXK;MJ(\=5\W^2^4>2G>\/(MdfZH\1UZ0
C&09-WKa5/Y->#b/B9M<>N--5M]Z8^^H=OD:NP/bJfKSK^H]>QZgNc/G)3KLG;.F
U,gN,9cK99]P\.Ea,=B\;:NYM;cXNCG.#dD91T3\?+1gW=77RU->P\1V?7<LZNNP
@b+&6;T6ZB)f^2eZ7\6UXeV6Xad;,)9^7G_CPf[e2aNF,)\/<IIK,:AKZU_2JK&M
]^TH?g_7WfeZ93I9ZTg+;=6NE\[^(Q\9dD:Ga4b(g4NCg(B&-B-6f=Yc,=b4aeJN
-AVa(.ZWBZ#H?)@6HCI,<=.Q3/-.5]/>1548T9.b2RCc+Z1B?NT@FUVU;&AC[b2G
[>cW,+g_1T-K?L9=WK=U5FD;f\H#RC.7X_1FKZJgVUYXNJ.,\[4T4@=#:bX)GCX0
R-M3^U>,SeJ80WG:2eECKANJcDg(0P&<\BA.Bf(16g>6&f?V>c>/=^7QRP31KAMa
>g1?E>@c;?O:\9H^_93E?B)]f>TfC>ZAg702C\=CT]-/B>Uf+3^J,JZM4a7.W+/8
6EW\N@eZV/N34bBg:,.\7P,T7DP.=DD2629/3SGaER[FS]1.NWCV0Q(Q6:9UI[Fd
U^#?G3<JT:dgT;0-RLJJI?fF&.BKc4eFG-,4L07/P.PW4Z2@EeY0-\:aS^_W8(Z9
1C]2F\Oaf_6I)Y\C:c\[,He(c=@3gY4T+A1b\H3#.[U7cgRZQaZa40]?5[SXEK;6
b]\P^B.2:R64Ic?Ug.NSU=V?\K@&fA&I+#2F2IA_U-FbbR;@F1Ddg;g@?b<<1\^=
&XG&G;X94S:(FT00_9_V^5RAb&gFJZ;A1L=(\_H>(U5LK5;BA^VeY3+5H&>X;gG#
OO9XCU)R_8[Xg7,MXUKaMAe1c1ITP1gWUU@&;@QaR>\>fIR0?:K?[5[#e_E9QMbR
=,EX(NN3d@NPV2dDGdH\7+_F:#A_;VEX65e2\\O+M9FfU<Wbg7e1;d0^;]D0dE1@
=+TUFCZ7Z>?:=KQ]7+Kf:HBZI=Sa#]bHK+@UDQMXCaQ>\MDaOMG8JaH)5INgA4]_
4TWE[MPP&SgI1=R,1DJ0OS;=LJ/&Z)UN9Xg)c#F8Z6AHScb@:_:3Y_>AfH>1fJ=&
W]B?+;gRL:fKCVdJ4ZC1_MWLdcaL[I5VNcC\b#c)Bb]82N\0S3)F\/6]>C?9PYdS
1PD=T0\?M?Y38@QCWb-]QLTF<O+[_3.)YK/g[[)03CYEUMK74(CN\[?7GS(QC\\c
>f\.ad37\WIHS-VgaV,aL770@G=fU&.;Xc(C2=:KA<CDRW>0B/S@g4<TTe-Ue^.>
MJOdSDGbSCFG3JcDS,8Z.RL6KOe9?K_94++I2fb94UeZ2Pg88T>&W(Nga4SL[f5:
?Cf8NN;Qd1T7@QfG)]5E&]=B4AFGPfE,PO.IH:DW9:9<B);=0M1>]+;Gf+gL.F<4
=/c>]Q+DKc/FMb2?Y?dW[)[>\fe<LE/dHVQ#VL#6<ee+K,b,RTV9a59Sc3OYS625
+J)#\=L-.gQMaR06+VX2.E2e48O?IfRI#@HXc-LRW8:OWd_O9,[R-:QJ/&)=b]@S
cA^I>M^[NA,fg])@GcG=HI1YOX@,0C2f)#CA5LDCM)E)X&A@JPW-AKLBK/?f:YNT
gb?01F11U>FPXBBMS@Raf-F54IGcSAFJ>c?aBg/XU,BKBNc9e&GEI^)KWI?(366\
-^90Y>2/^I&Q@W(G[GSeOS//+4<#F0>aI+348=ADVJcW8(=?UYYO6&)]+?FUbdbC
8JE;0;)cg)/UZ1\F/_(2AeE+5VeZJb@T\\LW]SS,BQ&.c?;DVUTKLBZ,QIg<^+d&
&90?@#:1X>6M:T<):WE1Z\)EIUW=L2[U22_TTbE>#=^Q-<CBfQQ^A9Z&YXLRTH3_
ZQ[=94ISV:E_W<9=24U@.3aMZ_35N9]N>-a7+7I:MbYbg(9Hd#K(<2eIEQ#DHFX<
K)3\_BS<GLdY#<\,QKd+94>1=-\ZZg[Gc:1F:;:?(9>9+TM7-+:7A<V)YH]L86W:
U,-+F(,^/^L,EKC]Vd5d/3Rd8BL(+L.1gM@Q/;[3UO#E(JRbfgdK+2B8Cc.RWA;S
Q_#a^eG&C+#PP:7[eNc3Kb8#e9&:BF@[+bUQPF>dNC;M/+Kda/[9g&DLaXM49g\V
86SKA\648E6Je7\J0_2fg98ACBQ]Cf(5I4).):48#XF]TN:=8Cfa>RPPB8P6C&a^
D]&dWDgSQR+&GV,UgTOUOI#P=MMNVCW,_-aD)POaOFYbg&PDD(DJ.J84NMD>G79/
K_&0<eN+OC:UY6FF9.E064NST=C9051)9HHSPd6@WR0YT>MRV/H==&L@aP.6+8[g
aMV)]X/^4^&[14=J2=J?N#XYd[d8#&28fX)AF3;g-5^,eCfdITeJ44[Ye_>3Q#OM
0^T#fg,Q_KHHY_VIe77+QZV3LG)DC9P?c53TWHYM:B_K1M6<eM-23#1N_=Y7P8@b
T;&:OXLZDW]fAXd\[L[6;#_L_aZ>9[/J,BVON&2Ib8SVWW^dE0QR5.#MW?,_KF,e
dGT<XW<T27_[Y5[4S\[aEOKNX_YN6=_1^eG:b;EVGL83b0H?5E<.YKGf5PSM6/L[
50E#>25bSHRbEePGZJf@2J]Pf?>Q5VZXBD@:D?]V_)8-3R-3B>V=7IJ(8V5)_Jb<
IK^H/94Z]/^;c;86-J>Vd?ceHDTCKQZa((3@f8]>;(T2HR&1I/#bN:V+XW95_^CX
DT<J]O)-?O\YB03PbXP:78dg_&-(>0@bD=0QWcK4<6I,/QH.dMD/9Z>VV_eHT#F=
AB,/@1;>U-F@37(SbDS):WaaT?6SJZ=AQ#/UP\:/;6@.=2XJ)>M#f3,H@T;2E.B,
0Q8EF._Y^1):(Z#@P46_d6dX4H?9WUggH=S5/G+;:P8X.fD#D5^He^b-aO\QB0FK
4E_&S7M;E>Wc-]<;2b73-_<dRBQ=+U_9?a[).9_1JP1Ra+M:8HNHLK?DL\aH_6\f
I#8V48(A^[5JN4AQPCf\WUDf2aC>^+T&@[eI7^2;b.&)@?3D\8-C<8-3N:/GW@[/
N+-Z7e/3Q(ON&S#F&X/X.7P2<5GIE]DEcCgbR8b>0?2QdNKe2)^08_aKI^6E]IgP
O/R?[9;/d-HH/1RVDBOaY)+:Q@H8FG8XYW&ZC,_O2af\RAO#;+Z:/&P@3+K\GK]#
<,J3,2KU.e-OQ.XcOGT4&)_QH-@1-]9GY#1,6/)QE//IW(4-@-SaUFdfCDL0M9[F
B[SYP1e=5M8MPdS&&dI5<AZWUJTSK@DbL&gKe-4^Y;/d#Y&YV:\1F2\a\;JQ&JP3
a4@[=O\O+9FLH^V/C(6A-(Q)L-U^P5+96?#8(T8&-:ZJO=c]<6Q;f(55,b+d@L?9
84I[?C)R;]MbU=\8)QT\H]F.Y&96E4)IQ<A9>#/W,S-=R0<ZU\]f0&+(EXR[Tb.W
SX(YS/-a.TC-gAfW3JgU+ZJTCY^T3ZEH>:YD+H1AA]CTO;dTSIE0c=PMTUDXU+9<
-KC2L5^b8/RCMPc;:Z#MF:XOF]?[B7M]g?9Y\I;6W9,@fU<VCG(KGDL;^8;5(QTD
84ZGUa,agg@D9N56BW_]@]dR9NR>AdFSe+OI+=.eGZg=33d-C_,^823XD^UM,RNd
B(7NGD3)+;+ZT07W)1(?=BRUee@DAC&+L.Y/WdVF\.-E0eT8d8R6.e7&+ISF+5_/
RHRPALJ^JJXUMcMOGDM;8(2-#=,c.1#UB4@D@d+@^QV.8WV#?b#P+I2c:IPZ@LO;
ac=H>QUeNY+\#<+cMbHO=DAD)(PZRFR+7E,g55SKb)-M;6C=OSa(;V4@OOaR45<<
>\d--LD_[2f83[@3Y@feD4WT;bD.Qb31VJ42aIP+09dO&UYKZPK5#OJHK-UY&109
:W[A[MK^7=N(==7)Y1L,Q20?J;72K#RFeV^9E=:WeCXc<#O+KG;T87gW2=WML>ab
aGFDB^R@AgP+?#\dO&gL1S2U&#5-.+Q2M2\ffKYeQHg9K]dCW3QPXC;D7Q9ES#KM
>:X]I356,(b@E<+5M\[7/B#7Z<I>JFT_bB?;?[)?4QG;VeE5_])T]cY>\/G]IHSL
Ra..feR>E+.LFJ8+8VCWcQ.&-eQ7@QB8I+Z,a=XLW7d.BQOge6^K_<\KQ/O/c+.A
e9DF?3,?#XS,(S44c?BK,IF#1-,;[^1]f[FBP=CG4[.RSI)_F<Q7]E3HN=+7O_Bg
[W@E(S=^Y43#bM572DU5XfbBGBE\4aW64aK7WRCTZLKP[>-b+:KDYSW<,&aH/4@B
^+81;8[f_dQg>]:1\e@=_YbF:X4aUbeUa,W#[F:>e8Wg=b1)_TbgZ=+PN:OSfLCH
P2LBPDa^QK8]fC?DR4AUWA<HQW:3Raaf1638G2e,N+.IbVHcQ6>=+6D\Z^]0S66J
=4ZXQ_S-;0I>P/KTVZ?d\^a<)7Q,b3[EAF.J?,CL6&E#Z/<MFL+4cF]Y\bL1,+?,
X>LL.\R(bKV(LR0TV&6>V#=7C/-]JC\=A.4\:8cS]VU<Jd2U[&L9;/CUAY380V/(
WTUbFN5#4Y]f3Uc5YXH]QY0G;gSG9V@#:)f.5++=Qed3[W?De[4#fBP5b,+X53V)
T:DJ6P-?LD)]]3+\Rd@&f+c]^IN,T]32XF:4.[LV(W0]S@INN?OBM[RD>9RTcB9/
CE;Y3dKQB\]X8L@fR];;4ebe\6F4RD4d4dZ:9WPC=#g9E9JR[/PbJE0#ULcS73A-
5YR3>N;PFP=e)+&R==>[DEV1[CJA+8V=g4addf1N+;J0J7IQ[1b).@OB/=V@<&J<
aR9@&J0aXLQU50^603[2g5C&+GD(41U;;JT^&SYY/J-aJ/(8CUbC+O4Bg=ed03+<
H8e/UR-#VH8g#AZ)Lg@b;^I6:F#J/NB1N)b2#gQOJY,P=]K1/+]O(#<ZTWJL5MR8
(F+H_cY?<>26ZAD.#cV6bT_+:G.OW;.d@C&e6#UeZQ0;V3XD@S.WGD2UO\.8c:R-
@U^@cI_GO2B2>P00_3:#:QTbAD(>FR+/95C=8Y\>Id<]<-P9/-U3.F54@&XWEg^G
OP<aP0_]S-#PLL2:3(P08[CE(];@0@D#\DR-;=(GHbWF(716gLZ14=fT332:/84/
W13@[S2@E#OO><Sd/dRRB05g=Q>?bb++U>dZ)e;[W5<]7,6-VV<.V\4P,Q/&HFJJ
)a-<8@Vc(Wg6H5@M1_EcLL@DLD)LRbb.09M\/E[37F4NbY;NcK&)gce7C_&1Q4@_
X30+D8V/MUK9f<?,A.>UVg44TVIdX\Le)#^S5B[7_3-S>.e7f5RKQ_3.?K(3Na4Z
bVD&XcJ/=?T2T4g19SJ<a#6HDV=J[E(5EaK@-NE>&F3=JbHE9AM-,M;O\UE[D(Te
J^H]H.]9V&UMc7.fT@Z>:^\HLC54_Q812(,V:@U7>?+?>A)GcTd[F4g,@7WgK5&2
;\d]P@1G+R-07&UXEZffCdH\4>^UTW9E^L:#?\#8gaG9bW:S9IJ\@E5Ne#=&@Cbd
SABZ??K_HC^dbQ-;d)0JfaJ5M4dV9Q9BRNY=K(]3H=BG3\X).3IaW6GE6^^6;/_(
F&,&P^GD]CLbV)+=4HI3:2PAU[2]L<8[JQ\Yb-56N2A&.EfD\@\8YETI0;A&LEQ.
49.+29&L3g[O:/LeI:T[[@#<BR(?,5[\UIB4bDIL3b>FdU\SU.A1=H[D?cg>SWRJ
cF+LC6BgbU1Y@Rbfd-fNQgT@X+B(b-61<Z(D2Rg[+TD75Q+>.S<dJ)7MCX-RRa^E
fV\=:?WVT2[D/\<5;18bR10;OFV#_^L=^U,?c^Pb3@LJ-X0\U2G;e=?OT0GLd:/g
3Dd;fcb[fBM58;d_Y?1KYSX6>GQU+]V;SJ&dBbQPU.#,gF(FHYLCEcc?LF_.)Z?L
UPK@4N+H4g;_C7VI0DE-OBMO9[K6,]9KFd/.&X[MW_BaFeB1VV\9V&6KPJGKcLMa
U<(1&?]7S<EbbZZ-(S9J+@1N[a+LM@CJELY/XV:afMJ6DI9CP4aL4b0DTc-CdJ98
g:4B/c.<RE:RBH]>\R2:R;b8/eX99&L<WZMJJNT@/_[SbDSB#Z],@a+.-7O-WBTV
F)f#YGUBRZ<IFK\d1(=?NVZ2egY?:M@@T-]Ee.dZ8eO)O6PX@[A,aFKP:gFg4/(?
\&T4M80HF(\^?F^>b<X@D:4&d+L4QA4:-8W&?R^JMP?@S(6U@-^OW0&=^a89K-g\
T^-[>(?g=Z.3N6Wd_Y0eJC+aHPQPQ(7NGc,<]0,?97B1VFJDbY:e;a)+EMI[5\^K
<Ub-=]MF9]De-MdE)DXA:78?725=(#7Ge7&@f4NXAf4a^RB_PUgT7[^9c;gXb^5R
eF=TfR.(K8)J1c_CA)\Q51;a@^W5@JSM-dU1S7T9VGX<aSYa;&B.dY.1<(524JFV
>/HY5IUI4eJL&6MA(V)@fBbN1#6,BHMT-N7b.JN)^P#f0-7G:P[F;4[=Oa1I<bCT
>+1,cUg-#IL)#c)O7ANdV0&KS>G#_I)1P1J#./WXS+:a+?O@Y@,M2b2I7G^/W0e6
,XPZB:TG0N/?g=K;,JY\^;Q4KU([e@6I]8g&4aa6T/9:VI839)+AgDGSTV(J,@44
[#AJ;I6QC):cYQ(,XHB]^4T/.JHPK934KZVJ.^P48BND4P=9I.R_/[@R<PQ<bg]_
/PWCfVU],7[ee2\14P>[C(O/:)a+3\6NA6b9;]R0(B(&DFLT&>2BI8FMYX]@c\G)
gbAP#]F8(,:76Q:ARU8A/4dbZ1eGZCZW]N9e1?;]#;L,R[N&47EAZ@];Y;8)Pd.a
=]?YTf0[@eF&9P=R1_GUdHLV\T?]NX1&SJbI<@_-RM1:8=6EdI.OW.B7^eAb8_&S
GKa;f1?R;:a@JTff\)50/=.<e>?KTP3XXE_E[6SaIGJF5CXR7AD&N7-W-@a>a&]\
9)TN9F#S1+,QgaFZ5;580ML>./^aPZ(P&Z.H>5bAGXL4)c0C&6BH&3U8.&6ef46(
Q_WV/d9YFO)f:McA5@&P;K>)]+XKULH&(\=8&AE][/=>N55^a)L.bMVIL]((L/=P
[&8=)^_N/+2P)G[cD_g_IeHS],<^(]c^?:NA<D7F_cUHd(TQ=PbF:[Y0/b)W@?c9
DVf?;)eR7e]?dH8:V\b/=QLBOf##1+ZBAKge+HCBC5E61EeI6f646G?H<X>c;B.P
g8V1MU#CU2C8LP_gGBBTBOBeM<fRCR+[(<>UL@0FY&_W>T+[OX))/#:,bdc>eb5+
)Tc)aL@6O-bR3[U=F;OQ8bbbA]2OZf9BDaKP-EZH<X1@8EL#Q+CaMZJ:YB1bY?@P
+HD_0eQ7ZWK:V6\?5^UKL=@;6NY&(+BeJ:5>Qf:BIKaH/8?LD;-;M[G63]A/-:EY
J/?@9FNNA)KB4+Lg>4eQ57?75,T\+HbQV1Cd<,[EB\)d5C0,c27A+0AHNB_S<CaB
J?HZFb+5541@T.))g#.[V;ZSJ5NNO0^T_>;W;D2[MfY-+A<e6P2:EHW2JF#HTSZ-
N6ZC^=,>?0[TD=TFCX_1Y-IRCD5A?^MR?[KT8UX<K081aJ[WCEaJGNbc;7GgP:)e
fVPW46(50Q_[g9fZ)L/_G\D#S&a[_@]4b&L.#L3C>cQA_)M7@9X_9C_eH&8g=POT
:TADY].2cE-e)0)5?T7#Q]UEL68<0b#NC9Z\;BTNXRdLT12NDQ/CZ:O>X?16/J@R
+Q9L?BR,:]B@+9\d3ERO]0=_#L2ga/B.8:@7CU;R+YPWPNH5;ARceeKU/C[=<.XD
Z^K_ReWOR5PL_@\]UYBdZ3WTdSHHB+.4QSG+BV)YM?3XaUPZK>c:TKS)H8UA,/R+
3HLGNO\&B9IdI)aFc\g2;d_>F#/#Y010W[G1C>[]D&18L[128U++P<f0MTIM.aYQ
3=@M5E)b>R@2^EHN^UJ0MfX/,52FJ3T]&X2X?QYdIU8O?OT)89=LW8/Ue9CA&K?V
&5;4HVGU[:U:SeK0GIRSO2_>]7A3Y=-5.:\dLTNca[@^gU6Je^?eg_LNZ)D&[XI?
SEbO5F.dK@TP^egfV27<REL6;Xf_&ZJOYRV-J=#dTW,7WDU<7A[)0NTOa]df1RgH
Vd8B.bPALf5\aIKERa?Y4X,K9H9CR\[?K(H]>eb[TT9E\E)&?b32-18+5(#PTNc,
^<5Z&?Qc:W92.G:)KL&eS?Ld615=>EaWA#NAGXOc>D2?gIF>f.+?<VHg5a,<(A=O
Z8LdCb#SVP5,YV&F7\Q=VQcM\L3\]-;L<4M4&OX784YWC0WOMa5XEL5^53T;K]P0
;C[\gCR4f;\4&#0>@TMa(]FO=\\c6KB;QaZa.]P8V))=eJEM5c.eCKK)#VfA1eVO
QV[5L4RWFLH/bYT7G[/fcCfM[XM^0Pf(.dI99?d^]E/\fEAXea3;7OP.)1A\I<0T
H)QcS)Y9L]e;XT-17EDO9:RE^3bWK+VO++&O&=>2S0L_.H^I)X]1Z<a79HP^TS^:
1[?@)&bIgFDXW.HdE,0V(aFVKbO(C)_;4R>NE3<NLYD7gWeI553RR&1<g_)e2^_R
\Pbd&+aZI&]0?JW?\DZBBPd/<DUX5?f<VEK9EQESg/8GOPW+->a3TKg]/LeU2NSg
a2RL+)eH0SL=ELUHXHH=ZGN1)QGM[BB=a6^(2_A0>/;+ZNg=,_-PFNX@S/@+^^cb
K-QWZP=CACf/YK&&-O2_a]:K&>6Q?-IQ^IF&7VbeA1XQS?a,Q9T=I3Z3CZ1+:-,&
_?e;)69g;B1TVP#dcJFJY.5^W)]e.U-C1Q/YD0gIT^+ZOE6W,I1P^gJ<-X0D>7CS
8;V/R38fM,ZZCQ0QR-1=+CPYa(@+1OKRP[QN921,]bSTW0=U7SW04D)0(SK6L=Ob
M4G[SXZf3=1VX<Q[?D&G[cgE0X5V9@7#b>]\?gBA23S@&]91XSG^3\aTc?Y3d6O(
D\GeIf;J0[HbTGeX;W_2D#EeQ[-8TbKfMQ=U9gL:R:,OXST=1&CBQ2>GF,adHBSD
MLC;f5#;:3B;G.E@K@M7A#^2B4aASYH18]Y[Md;W.:d:LUO.T30#JD1KW\A;=/A-
NL6d[IAHd_\6SMaNfEc.>VDKH,S#DF63E4(5b9cZb_6-2=4IPV1cQ6g[\K_[]^60
^))WP4#,PCZ7a>3H?R9-)DQ/>0,R;@)OS;WS@<AMB_gfQG63gA[ZgaNP-c@3._++
.-)c1Y\5O594YfUJ6AA]fW<,Z.OeJ2S-_L#HSgX]&RTVV-FBLV2&2Og&:;GAYdQ.
9e3?K>ag1f=:X2I+cVfQ70^=LEW&)V1B[:2YSD63b-Lb]#JRCF8T>Zc<&ZIKUNHe
Xg[S4#;Y(/M1SF)dfddg2FQ,@b16.@4X#1X8V;a=6T1eO.,VWF=29AK]L7Hf#gTN
W^24=&9Bb58IS;IW_(^M^c^gVXZ#]bJNR/1A\/MS0D(&>9^)Vd[b:DAZTRHNdZJ0
V-P^7YSNEL\[5N=I^SK^6\WSag-?a@8ML^XRW9PT]L?2Y_B+C@C0TaHDJWJR&4VX
@b3Y/<fKQLEHa8b1)[Dd;1\1:a(R6L,U3SS,H\f@-Oa69YSfQ#;b_KA\H(.PUMT7
c0,4WH/;V6#1B_IecY:\dH-<27)S9@Q]b9K1b:OA.K2fNaVe)U.XGf.d:44XQHMF
0GZ1-UTO9C];2bD[b4fL6c&Uf.A6R1ef>BQ,\C;fSI32.16<:-L;L3RZP9;:9ZfX
]cXWe?MD91=d5(##bc\.R;[;J,F@1&Y;-L3P@+SBBV;0HK,#)B&Le,Q]IcCCPP>S
SWT3]EF-A)C_>f1@1[H.1<g6U8QD(6>ELdXB\#],Wc@gVFZ<PFJb\8:(cZM+O<T3
6?[[OV_@4W49e0CD]]3Y<X0dNRTM^+=?CE^<;WQd;&c3ab5;&LK7GZJP\>L5g#;:
]I6YR4(.Pe=>[#OQabdDNABe-Y710ab@c@GKNNDEdWTQPQdQB-9WTga,M^K\K6RT
,VJ,T3fO2c^,8QCcZ/J^BLH#YPUad2fY-Sg:ggRa8B-:WVXZ\@T3Uc.>S@WPS=IA
O:R3JV<eOa)P09?8:.SC1Qe9LATL]#-7MUgK9QC85S>/<c>1A/e0WT>DUG?\9\<d
5-g_fRO8;O0gI<^<27Jf5<K&L09&04?ZS]HZNA+(EDRfZFUF1UT^X&1T<1P=6Z-W
4)<T4dF?L:&.b;^Q<Ee];)U)FX)>.=ETU\gO^eDbDQC+Rc6&:J9O7g(EM12T^Ff8
dY7MUM(O6EG[WK</&,435A>M6(1R9FF_6MN]N^0fFW_cA[Ia-HSLNK<CJ4&1C^3E
^^.?XD)1O&4W(cN0H_6#Y13J?/RF<1S4L7?6O?TI,0cZSIXeHLY^U\U;_2+e5]H@
L5=#/0D9VC<5+KcSN^I+K.R_E/@+/^@+;.SVCI/PRQOAgZ0).9&]UP2LDVIZWf0B
0V[Y^:X,UZ.M,f]b,X:Ne?0@#RgG:EUC&45=C;CcPP<gdW.H>/GP[<e2D3YeCR:6
+OAaW9JTMWO5QUd@U3dQ)(e@]Wa1WF@8,8I[WCXSgK^N(+e#/3]+6GGYII)Ef&V,
/NZ-J[_0\XGB(HeN@6L;FH[KL4(AT:B&(>Z7\B>=U2\Y0=f>D0BEF.[&AG?\8O#C
+5Vd8#<\J0H;+<[O(?)6d^7L;QS5[-G2)U,@K>L0;/:3R&DbE_DFcHQ<)+d&dQ[U
Z]Q<X2:2N.#Tg9444(efa^0a=OY(9T[228_15=9f7^?(:;7QZbA.,U]W?[CO=aK3
M0:B+)23,9WL+T/0N07#=D6).2E.I6P56/5,b^EU<JCLOYM@WBZHMAA5TOQ.[E?.
7QKX&RN\=(PW;aW(Z_VOE/4,g7)(-R_QF]PZ&g2RH>fTY(Rb6@&5Re[WG)F0?Mb,
:T?X=DG=PX5LCDVSQDG2)G3[f5Bc)F#CdH]9]Sb,UOT^M0)8FJ5QcMIcQXO#DK-\
K#?6WY\^=LIUMD>0WbLD2SSN73QfW:WFeX81>DQ<9:G5cH,Zg)_>P@JUAg0^G.U1
7XO7Y-3fC6O=V5#93404R4#\f?(8I^gN_b?@VZC@)(JFaPbQ]]L,7Z+:D0[MN;(c
S-C]7<7<DJ:,#LZa.+\>S-LM1.]9BJDI89LS/UW^BZ\I4ZFRPLNNATIRC()g&gRU
;9O-20a<8[aBJfL?.Rgc?8I#R)1:-Cc2-P:_S:Cg;E&OBO6/O8,O.81I(NgG?3+?
13MM0bVQW22+S+O()N(gU2EMV]KfH,gC(d0MY4I;4<(-6:[a:c:/YE?:])(BV?.Z
,(6NY5g#MGd_G)AS77=>#&JKBL3C28DO;U,AK+dO3F_SRb9O0dbELRDcBBV_=O2b
94f6J^f0#G2RJ?\,X2O9WUaA:_B)G#PNJO)-2C:(Vgb4fXJ],H]:e[^Be9I=Sf3A
C&](0HceLO\D7J>9[74f#NP4/XCOU49]Q0fP&IHYD[N@.e+72EMd?FMDUQM:<YQ-
CgV[:5HPVS0IG0ZJ/Yf<B]2Pf2)\.U:<B:>.V[G(f2.7)R6?@FBSK^aEC@geWAg0
K5Fb#_0@Sb^Z+bBFCd0\S&.FCHYba\7b6Ie5e6(V/0&<&E[/CbRC][K96(IVGDO+
:LdM3KWRe(==S+@(8Q96;aTS;HNF4cH)bY]A^CQF8fEd\,+0cdJF-;@Ka#7?Re50
=&-N_Lb#X@\a0-52L?+aDR]#W&HNKaW;Z<Q)HG8814YQ570U_L56c+^@YJdg2M(U
##4f4@>.FY8.=ZVZ\N\7:I/D&LN[eI-KAHU5Z9&,-49EcI,YMQH?5e_d+J:)CY8Y
Wg_JJ[&YH>JBZf4_DF)1/7X8Ld.=FTK3X+(eXB8_6aAZ6SXI+X-M3#HUYW[CFP7a
_K)c5dT[3EQOa;LW?0\7(S:EJXQWOQ5W@8?;>S1,>N;)0P9dAf<_EPc,e>BV=-&C
=c09A-XA/[C^cAg3/Jb9)HFE\b.(<e8>:NZg?&fUF;LB^e&N9_UAIIOJY_QP]@87
U0N6cQ<:KDV>L1O,b7?6BY;a^[46TNZ(@^c,>S7NB>:Qd&CAH5)?5?6(X(DB.=Rd
C#B[KTfgCg]AGVV4FL7Sg6bGW+eP)LWN+B-7T.SYJV7@[UYYdI0V^G2=_:&Wb=XI
DFF\T5e,J-LC#QF][14\2)FU0)LWX2a905]?YG>8S3/ZGFXXU2@)Ffa5&M+V&5LL
;b3V36Y=d7<-4E/MT]==MKE/J2W?K6&U>^[?4L&g=I[QEFe#733e@RN]KO27J93=
IAO:[aW<<O/,;1c:7EY5U#Fc?DZAINE]Ge3LS(/19PX6343cg+K2JaM#4QeQOACB
,YI]D\)8/gCGB0MEREg_<AL,<:^1[fQ)T@]^O8TD&EJ7[EF.CAF:BQ<&&HG1)(Cc
<.LD^9EIA??1TOHg2+[R_BUNg9P]-2L1:I@BOW1Y?E,;XgTKfR[Zb3]M+8RG4K/<
D]54cdK&TY#.NTWOSDcaR:#VDB65BIYg+K[OWb68EgYH:BJ1FDY@:CeT_YK<6FXF
V(.J@VQNRGG-JPB1;?2;\ZLHWQ6[bcTJ8DOV:UaNgRHR_Mf\1HGO(RISZ74>FM[/
Q_egT@Qd<6\QUcA0HLZ>;R)6@]#PS=1a-S\PV@+#ecC88[1DRK26PUNKG[1-88(;
-daLPZFATS#9g-6Na,WD?8gbbg7b[MB(,PBZP6/7N3b[ag8\LC_LZFCBWP@4Jb8N
##GZA#NJZ2N+C>5f_MU1TFAT7+3AWU2B&g,/17cA4-Ha#?0e5_28S9UBV140K9Jf
3)FVPI:5;\)2IIX&GMPM\0](aQ\?FE^09[b(]06BGKPf9</;2L.e1D7D;@e&9=\J
QNLF(98>NY=g+.B](]3,:_C;<OH:D]6-6UaeXNEMROP[:37C#Zg_CJb);<Vbd)TF
ZN:H-[L=fF]B_OH3.S#gbI=HOWfP#d>9gc5>ff4(F0?W,J_FS6OGOQFS/Ad1>#UP
\)UHV+#IDbVCaCWYBcgS4WJB??Eg[Hb0X,KMC[bXU2.)8HC7dT4L,IHBZ_e-@<)B
+[)4G3UF5)Q(UZeBW/@>B\@(9NX?<b9UYd6/9GG@gcW_;<PM33[[BC8EWFN]]R_5
=?VE36-Ja6_U8RF[J&(g:Q2McXL(4M,b3O&5DF&a5XeggH(b[>=ZFL7&J34-11/6
1Q08,P?bL9E))8c0IEXX7]_#DCRQYL3/4CWO,cU>aX9TN@(I;@6?3?aV5L\SNfY2
-2^N,EPTRS@Yb7.GX0DO-#bC0R?A4M=OK2+f>A@68OKA3CK@685LVAWT:Ia-,US=
ZA)(I=E0]bMEaF_VBF[IH\2<.7cg+J@HJZeX05VVe7Z2a4T@:Xf2;7g8ICXF0>GX
EU.9S\83441YK\1DI/1];9N)?8OF9bEFJ&-^9f>XN:3R/C29\K#L\Q\OIA#g(4Of
NRUXN;<b,@JfJ/]=OH<4#Y>/K;5<D1US69=7QJ4N<50P.YU<@;TO(Y\bPX\:7D9F
[^B5W7c26#:g_RK,cTOSFS65[YBD]Ac^O(Xb0H2IX-gGb5/C5a_LT\YK<,eA7+K(
.<]2B;)(?>9AT#aC5IE1B/g+G.6=SQT;Ab[J-YSZ1aFE)HQ,;=P3\J:dD7>=UR6S
Y7>7W]>:d.BbOEU/6X;F3BZOE#:_:.fb/\A45D8H1J^gM6+JH.=1Q8S&0>XT97(_
#b_gWe7B0-?MKAUG/4)gJ^YM;G9L6[H0&E<:T-:+H-?MKF(Ic2YRF-\0f4JcW@D,
38^8,a:2=?8eNMY[5Q;16^_8O?]d^(CJ@QNaX<cQKOC1(e(LOK\#3W[ASF?.1Z>:
2MQIA)Za1ASU#,MDI-EX_7MS+2I6C,JUaP0Q+],4Nb[^<R+^?/<Qe4ECV9R6cR(I
/)?&=8N0>D3GJbZZ#UF#d45IS@>8ESI+HbW5T+^TM)Ge00:]#G6B0?#?9&FC]:GL
6gY\HVFK_]K.]C]QVZI:N<OY<9X4cOX_<[B&dWgL;]#=G.8<[cabE/aB1WaCF(ce
RW+<#-J7ON0Y>;Ad6#e;\#/UM72\=1:f4K43#Ugb,)89BRcN&>-V+^TEN-SXbHS?
0K_a&]B,?ED<L#EM3;[_eSYL@+g?cPF(C9.g2cNNb[ID<a+6OI2U\eN\YKF#8gRD
HIMLe.0HJ0YeVYC^MEB4[X[DXGPFH2CcD]\N=XV0&TV/PR:Da;F8Xd/c;_(W0B,0
\gJE0PQ/XR<cJ[NaKQ+9?/;N]85I&=e8Ic8YF@_M\TZHAMEGM.Q5Y,2Rfe(GB698
[(H:XFeML.7W0;EK@Q<UN1X;0/8#AgJTTcSVU_MPed6EfT8);LbUZ\4@R2HC.b#0
>^J>]RWIZeIQF^]g>\M2^WK,/4K5gKF8XX/;67+Z2HgJgE#FcB>g339\S9.L_d4F
\cZ0C4/a@g5JdcH/8[F?)YE\4@EM&fNTUcJTJc36H<VJKQWT=26eM5=NZH]@0ZOO
(IAed1B0;W0F)b.LB0T47;c<Y,D2^@73SFP)R8]K.E(Z]4@d&#))FMOZ@Ic?2;Xc
>+WH>c0F34#gB&:[E;a]@#9G)=3._QAL=8[6fc?TXdUX@4Y?J\[S#-V)81TdgQQ:
Y1],2DUZN@]5DegO3c;#?=(J7fSc?:&e00>9,<2Pg8LJGW142_B\dR?]S_Q<a;[&
##GKQ9#2J1FcO\2;A/5W8bQ2Na5>LFZ.0dLZPT29;;eZRI-E.3aU;fFfTAg(A]4Y
e_=c_:?6W<?RG55#H;@#^NQH=SAJL.\,8Q5.^1^+ZN[^R(XYA-P6GZ[_#a9K-@V/
7:^=R9YR]E;A:Fg2\G_XTA]:#-OG+?0GU[\M.A>5:Rg)eV;QE_>&.:b2:b_EAMa<
Gb)aJf@TVc5W;Mf+/;eH:I>QTVP3R?34Q_e1UF;UXDb0-b.6aIda#d/LX&TQ]^B)
\AH7(gZAQUY[#aYPQ2aUC_(cG_MVNgA]/Ne@#Od@CJFC6@3JNS+cYJS+0+FG)NDQ
QZ<Ifea->@(,#FPZ-WOI:I;80Pe[XGE^URbG-\A<X7(;-#g,<XT>.>TTTRMc<U9E
T=JLHH&2USSJOSM])@Gd4-(_U=@@PLa8N:RPeBUT21S.:f46F4H4gf0F_>fYZ[+<
W53?1W8EQQgF6;aa=#(2J&OF3<&Y_;+A_V5ITUVX2eHOe5;IIF<6AK)VI08SHWP-
_(C+XBe98)X:>-7IP3JNgc_Ne7EGKGD_NA=[R^Y&bG+CKDBg&bc_9<,R^Y@)U&<Q
LA5Ib),bECF0:gIgXN=N-+,)H7.ENKYM1?9b;@]HZ6QIf8b0.DJ[2&T1N][/STA7
P:Z/9)]MPYPLMH74QE:bH=1DOYf+<_HE[\1I)c(XGL0E[(/3GX_d;EAL8-dTge,_
#)PL>2V-&@/@d(BY+@K<afB;LYF10K3ZNMRdF0]&68KO1G0U9(L./7+/[a:DG78K
0J-Ef:2LQR#Y#)G\(+de(_.SQ2c2M=(3V&A(0CN<c@gPC1A@d8@]--HWA=T5.C7Q
TOS^OO\=<E3cT8B12GUKANa726QT+BXag[/M]35LgPG88+<F:#[>#9^C<EL>0WeZ
#COc>[5>9&__TOg4./Z^8Y+<Y3Y?<HK<AEFC^?gH>DQW+B-P8?:FOCYb<^T3Y,N[
JKNegIHIfb:f,]3PDZ#ddS;;PUO2SL6&/7IF6\D&2UE3dLWbgH^,>g>WBf3/]A)Z
94]Y5fg296BEUIM@LU2S/I(7?#IS(QZ;^/=K),Z5GM2_H/6Z-_4.0;0:)N)>.#9\
bINFVE(=aV/A6\Le3:(3<M;f:=W#_F7@((^AcHG3N#F_;2a)>=L0SQ3BJ6ZH.RTX
I]+bd0+\/-K=Sg1f\=OOT=H42;^LZ^S0g6U47G(VW/F7I0#ODe+[C^PNKZb@>ZU7
Y8c8+[27^&_+VDKH,XWQ6cI8FK#?FTaIe<=6&F\15[6?f,R98(Hec_a8VBPO-)^X
@,WWFOaXdK0=#/6>DUW#M\#)77S,CZR#Gb;HZ?4YX@/cI?7+(R,5CF>DL_ROL/]M
TXGg+HX5MUPd4_GHC,S=ZcMA0VW^S#?fTdgc?@]@NW[I#6,&4-JfB2<bN]f;A>M6
,=-#;A_g#d.1)4L=KBLYA[3?e_#Eg?aFIL)002K5?=+.^dYG_gMZe771f1.#Od:g
A.]>13gR/L,c0]f@\=>gg(5a43\;-7QY?.BIHaAcU9fJZL8((D28K46)@eU<+F)K
[H0S:RM6W\DXCF-f]Fa(_eN?T.M-+f.8L49C=BVV26e68]KA>:LPg_872Z#aHcEP
.<MAC23]AD6CCc)XL_b=IVX,P\M5^K+O:CQKX\]a-RaY.d1Nb^;C\de-f?92V2^g
FCOQb/DY_NSOf2B29BF8@K/>ZC=DL+VX9EI2MO<.BOOUUP50F,dQ6<dKQC:fP_aU
eZF<VOA0g]/-Z4S_E22S>Mc(^.N)/.0_<44K&g>E&,@_a?8D+/=,8cf]<H<[0ELR
&NPAS@GQN;K[L-HZ\,4H=+W;/L=e/G(:5Ba80PE/QZR12@\XLOWRCA,[gH(SdOMG
=9=ceaA/87NEIAG=MWLQPHKOU:;d?2ZUDQ6T89OI,NI@.GF<dDXBJ.GBG7fWT)(4
f3Ra.Yd#<d>M+E&9QH@=6_aU#R:6e<(Z_4a-.2dQWaZS>_O/2XE,D?5E:b>=Td_8
5]@D6#.FM_<,g\3=))MG]3<NF[]>SO@KB\RGB94&.fMUHKY2D@QdQ)BXR9Z4[c1.
bO\NAL,R/CGc9db+OL@<A_)E[(=[W#B45(K#F)b)/Zg-aPfaW_dP3@L.PUe7B]Te
#>.2]PNXPe[O<JR]aX?<R-@fEGH#IW]L=$
`endprotected
    
`protected
G.SJ^-,QKCULG0]dgQ&Y(dD,@T(VaO<.@M/AXZRPDDS\8R\D1eA+4)c/G\M1YMJL
8e/]d5ZUg?S5#RI_0OSCgKe5SEM+D#Eg[2S/1cfMMCW)JE;MZ0NK8?;L<(PU8,FV
eA_bf9eHe[I2fW=_LM(:7(EHA1b0W^gN<Z[3].-QQGBXb2I<bHe-?feIMU=caE?4
:A@0SSaCd^1^7cL+2P&8><f3eK]d,T+U.\X5;9DGAL<<CBN\;4:J&#aTW7OABDFb
M2JZbUd+R,a:K>?:f-8AJIV@;H93KTWYH0P25,92cF.O\96_5b_^U4C-?=5cH>50
>^&&H>a7dQT]-G1B=6;9+\ST;.NHB4cP;Zb818SM_G_PZ7P4LD+d9&S;NbFOBcY^
3JcT;0FT8SW\=S/\TC7c6WUIJB7)LVKH\9K@DV-3<H1)UaEa8Tb59=2=#4NgB:gP
=:Z:63Qb)#<(J]S/e99fQ8AKI8^3T)7/PBIH-\.Z0GGYWP0+GZ2=6b.e<C&.0&d(
VFG6V7Xg:<f=6[=NE,<VYVEKI?L:ab3\;dZ>87ed02e6/ZF]RIR^6F/P@J@EGBX?
IXO@6J94UF>^[;02ZV<#ANaK(5C(Rd4,bN#B^#PKZNd,P^KG.eNR>TS6dX06[cdU
;?:_OU_+17D1,L>V42J-K08YOC3Ba0A330,QO[X&31YUHIb@Fa@5Kf+e;Q(FB4CU
WYKFPbU^(=[C]5YD/D50H6/IdH&Z><C:D35Y<6f?0/8I(2.K\C?,?=@:HaP)>d@a
FETO&\@F,=REV/VPP&<K7XL3,_Q^bG4,bU)aCCfN3B3JYN-\F(=S:(@2XfXQHagT
d[/eHYL3Vb-JF6JII^Ga[e#3M:0M:fM/-H<Me#E>L/8-+R8A#_QK[Pea5ac0BAD0
K/:Eg-4-HRSN=.7:b-dM5UY?cZ>=C)0#NHI0^?VYf]C4>SXeceC+_;KZRgdNG]ac
TT1cA=<F##?95aW?1)F3Yf;CGUb?81[W:K5[6&IIHM345)(Q+P/<RP@:XNCga7N_
H)I-D\=71UVZXKIR3QN[WP.,/<3fN<II]Fg?)KDTC5SH8gZOX+E?T<K9_HO4Y9O9
/8+3_Y].-1I01.b&^X6W&<-HeM8P&fMH><,67:4-K\VbTUc<>QgTW92;gJaZVgFR
/3:84CZ2LNU(@43X@@/eCA:;IWJ9&?W6:L46b#beX2f[-bFd.23RR]>>=Y#1KYQ6
F5fI?cW6#D4PAK:PDTdW8>K)/(2Q<MB_R,U674A(</e/<^#f^]T@4JX9UA#E2S@B
DLeD/gET4eA@9_D;]1\6U&Wf(_dOJT;T\^9P]=NU15Q_EWD#FcN^,-V#GSXZ3A#F
45[QXT0,Q/QY42R]4[].V-)KUT6bS_(bZ\),dM4PBU.:LY2K<V][.WS.D:=gf#ES
aVYKXD_RMc>@_(baBfL.6:2[X-,L_07X>]Q-W[.AHE)M_AHSa,8?=,D3&E\Y>D,,
#1Z#S501=F@?+ePML\Y#<0]MU7S@+:YZPE8W[@.Y197+9a.S=Q-VST5EHd_[g\cG
K=PA8Q7eH&Q\XT+<ef0XD0@+^UPJ[NX.&ULW0RIW\-6/EWZ0H314<,U3WJ<?79/U
,#=1AP>.0?f@<2Oa<-0.cXZMGI<3Q8C8N04UN<dB(\LcOAa2[d2IN=>KD/L/X;-g
GDTC.@TG+7d<Qc]F;;H8?:XT#dM&F]Uc5ECc;9O1B,7)@P#8GOYZ266X4SYS&bW_
:f[AMN4N<[X@THIL5)P-R)E6]CeM?0W?=M2;d:(TQU4ER#^4T:?FGXA9P7.&4UFb
TO#aG3A45-VS2:77WgCB75@gUDE6.E:dQ#7<NAgXPU2a\JaR4U82@X65GIH;Z;EJ
/;-J.Y(]-H3GeL=1@Q]J9:Pc&XA=>O(AL7;gKFIX(bZW38d[K0#_FJeM8T+#a-EJ
]-Z78#\4K2)D9FfdC:#8\EW(3&@HQca#\NFf;_@FPa-9G[IO]RO(>]P8MHPdeR<b
U_1dD8I3WW5?@;e0e25LA16g:3,<D+EXESX+Q.UD4E+Z5N&V7@bN=E.S,19Ee1=5
H^K0dLY4YJZLBa@Af6R]\J9JeDH-+c\)X>KdODeQ)FXe&N<.754M;F9<a:>7++RB
:?4?cg=6]Q2f7V(Vf/J>fP=aW9L6NMY?;)_.ONFZLR)EI+G#5DK#]K:--)789WVa
ZHQS3/YLgA>&I/CK#]6@QcCYc?FID_8B#J2_e35e-W+?PTaA=7,ZAHLJROUK[M0W
5ac@W_QU</\?L/[ZZW@b\d[3TJF,(>5WXX97Y1fRBL;(..IH@Kd_##&^a,CS>OW<
4=#eIaf7EB/W_/c&-(VAY=V@A?6GVG>d0)8M35OgRP-W/=6aVE9eGILA>PV3R-9.
Q[\4V-+##@a;4J>-dT]YQ[;-QP^3fL^@S(XD4P714CEU,cdY:]/M8#JK9Z]g^#(9
;=eG.#QU?.QG-7D)F9F1HXVcHcLeB4&_?&D@LfCM6JBdLVT/^-;3B+.SX8:\fJUC
^faB]B:^8:4\E9Z^bfba+/SfX.4=H;^2U1D]V8Iac>@cGH.-(a>OXB/E_aYe?JW]
aN,O05O@7O5.+MDD<#>^-7>F4T]KWJ9=8+2AQObUS:H0@BA6PS@D8[>6Y17-H4>>
J\,3=)eZ(T\K0[f];-a(=F@P7((N0;NVW5&F<FMZcYPIQEfH?.NH_05+-+^K4QL.
Pcg[&eJ]O7(]dTC+:HSQ\FKL=e<MDcYN]P\NR:d6X:a5SPdB+dPW7],<\eAI_9=T
)dZWd5?,0SI85]E1W5#Wg<=FFF(D.BSCIAaM/cK75/:S04@-XdF5g1IANcJ\1/N\
<f)N>S7Q++&d)5?-NN;6c0T<[X@][OeB0ccb4-@gBK]LL+N6KK()6BD7_&[\;#==
ZA._WMQIa_&[7OZ>9fbPZ^^B@aN#--9#,ZC@46V-8UOTc2)fZPHaHPf+BD7b;?2(
CW>d_K1&;JeWN(V>6cZ@FdgEIEQXL7_\&8;CRRKY:M/7<FRcY-KXBBYDA<N5H;cO
2O8_&bV?39gDF(Y5K3K4YgBK5^?-A^TK8_Sb1@X\9LQ;4AV23c+]7DX+OYPEFQ1J
TE7&=aYI<?B9)IScXH&\b2bCV^FZ<W)SU:X_&9WQ)7<P72F5NG]GFI5BYAD,1<aW
0g;KC&]B^EL39T[<L@SI5;XGKg-A;eK2DCYOY:Rc?9QA<Og]UaKTQ/[W)9<0#5.g
ACa:D>N\L\MG2<#gBX14F370=0Y7,PHZO-?95HL2&ISD(99CG3X[[=_d]eXc@BX1
E?O7-4:-)Z&0[.gZdcC5N-d,SK24:R;+M#AK-JUO2Z<8(B?6YRG[^4D[X#4,+N;>
0X(UbRVBg.KU7;-/1MWVe,9CXFaR__]:U-_f1LgdLF<a@fM5M&&&@NQW[a5YL9f6
C[XW:Tcc)SBc\>_ZA)VI_)SF5_I;<0S\063^O188=2C>QTV<YTM<BKB<ACOPEdd&
@Q55D([NQT5AINH\9Z]G6Y=V?O=@b7Pf1)F3#:5HZYKZD#EW(D^gQ3c?B7)CL+Ba
ROf#I@^VeLMR94>3D9eV:HA8.ND#QF/0f,/YWT8d&AIZD$
`endprotected
    
`protected
&I)[TY8Wa#FgF]3Q&DP0bQ=0@5RdXEJ#ZK>D6TbfR8^U-C:SM]687)1H6;M/,C6E
eRf?g(;@PF2^C.M-/DNJ:G-/(dcYb.X&>$
`endprotected

//vcs_lic_vip_protect 
`protected
X)<5D0S03Wbd1Z/_CW>A+a2;^^]P75FY]UY?B\3MK9H.@^7KdX5Q,(9@RYgUL3#_
b_g<SL.<_WG<6IWV],#gdJ=),4eaD1RdENYHHTFK(+^\2TV4WRMYBV/+):^\BVKG
47D-16=:QHfYAZG)\&#QEODOHW>Ye7HAc.BEJ:0\B-7CX5:<(_L+E^Q9e_2;+KM9
H07WT9]X?b)59]fcf+5/.TG/,B/_O)@MO)=,W1_Le(gM@,K8._.=J8<c2U7S:cCd
,2+40&<cMH7,^gDUUcX[d=)bQ>=g,eB5KRgH,J+d&NE[=g#2([30@(W<,E[&40,E
9)9HZFG&D7;492J]U^9@ZS_BEN;L6REBY&G8.bZ+Q<&B>ObIbEF8dR07<0+f0_2+
bgW?3?f>NJ_1NE2ODO:afP@LQ=\ENGHXWggM,FQOP9XL6-JP<3GZ44ZYSc+eU(1c
1O+\ECc2SR.NA7g#-(R8(</;0?<aKI8SdfPadLGc(S#ZHXHST-6a;QZ+3LH835B0
,9W926[_<eGb^X_-f4EXB8[Z(Ag;6+L5.;9gb[<MK)^/XBR+)^\EcdgF_N=OI#Q6
Yb58,JHXc3(a=6\:B2VQS=6/,]a<28D?UW3BYTUR)PSJ]=Ig.g>+Sf:>BK8cJ[XM
(MV=a7]&5G/Ue]5KW:>F,TH^F)#RP<-B9df(WF5.aG9eXb8&gg5eG,0N>9G?\NC9
8:A5UEQ5OQ[bTgKc(SPF,.3]H@f?(=Z\B5+Z3Aa:_9-FZ;KKY@N+F_77-c?)gW#.
I4Cb)-\F<\N8PD\g[12aU[aEZ5:cMUf+@VP4a3MI,N^OMJ><RcCc2RYg8#DL7dKX
=91UU3<+Q:HC=3>VBER=1757UBK&=UE2S,82@L9gUZMCc8UdB]BbBaEIF429:@4-
93.\Bg;VX6U-3HF?V4VM\S>5C\ND.)^g>=XAd]bbZZ_Z2Z=c6.CRRSZ3</LO?AR-
+(+__=9WWdQE^bS,ecYgN^8P8Og\S5ER[^]_fL3dTSZQ:A9#I?1NNNCgXH>KYD;R
FK39DS-OP=>A;P6RE^<4a1.fWVMeT_Ze/^C:22(aQ/EUG<#D)M^QY^=e+=bceUcB
2_@ZDZ2ZR=]PN2Y.&Qd4TL1WD@PQ[ALH=Q;(F3?;GTCM0#O0bB<BFI.867FJ0V5-
eRggM>=93_NU4Dfa]>IB+Q5/ZCO/QX_45c=X]S-D1Q5.MBA-/<1MO,GaeT5VH08,
6J.)fJ]9DgG0\9b37QQ9DRN-dK#IARJc<g2ZUQDK]d).GcJVDb/gc@XE_eEGTM+4
?97MdVdc8S>LYSPY[Rbb+.52F,SR<.ccJE^>8OBT/COS9?;F.J1),R#JPgU@Z&Zc
.GQ_G5UJPQ(]H2/IU_94gTJ4P]QcJW]D:@KD3/#7HQ=AfSdVAN0?)g[8GISJ\]PV
KR\/7AJ0;;Z,P<RG?C>c[YG\Yg22gAI4eA,NIe40SX\1Z]?a63](7+7VD9Z(\a9A
N/(+T[_^eQ1.4ZJg=,E7&8bXLFQaZKD[?CUZLVcQBX>BH_+-P6KCWc2E/1,TE_3U
OQ#?YR9G_/QD]NY[XJU3C@f<.a69e?FGY--3-LL^)/3Q8Q\T-E0TJ9c6B#G=KNDd
TVaZV#S<RdZ#\>+cYc4fM5#&85A9Yc/\XI_V&gcB2Xe?5>YI2^_9d=1M-V3+3[D-
:gcD_G)E#PgUN;/?Z7Za;e.b<.gVB[5O>/V:B4#.O([b\;;e-b8ddPc94#DAD+eI
YFXWU?dMSIZ)G(F30C44)?f:d;X=3]F[_X/Q-\(dNP/[WU4A.L>_fP(,MH/\EU+K
db[CZ&1:_4cA>:J,6Rfe4:F4B?8L5dZdO9C\fWC@?.2MgGP:=YI4T\a=JP@=ag#7
7_N@cWK[63+S>M@CLHVc>5CJfV5WgER;LdVZ\DCY;#gW(WgFf3THG,XcI)-fRR5(
\E(=9+cTSAL&.:1A0;Q8:P8WU2gPP.LV)TDG.0P0]]/CV),,.<_eB/?MQB<?4P=?
TDH((HDf]7I^e=1N=N(I-6b1HIY5bX-6IOa<\;@6OBN(5;O^YFZJ>I=1H8A>U,.E
&8aT?#+)R>VKA2^S>)@?9cTIZ(/)cPC<QT57;RF;XN.>=7gAgOBgK=<PO7)4OfQc
G(XSXF)#M+ab6+_\HL<,;PL:fg:^\_,7(?f,;T[\7PW77^_HZ&C>9Z.R#E(4f__C
]Q?#e#c&HZ3+SEcd<aC=9MSgS]>C11]O2:(]Lb/=N35g##P4UdPaJX9HP1KC7[f)
)78G0>JcFVIP(3EFMcQT&g=\U5_D,cAZM\].?)<6F?^H#],XV#OK9e-<VO/Q<@)d
-@SW29(@d<?^+R#V>ERg&,#cDKAc=0UXC;46e&U\I[DQ^/;Q:6>;1<M)DPG8=>MN
NgGbXL@V/9VY,E1VSa6V)>;Gag_:/K9&OO^;MEB-dWea2Z.,TPR<THbQe-FGR8O.
9,A;>Gd/[Ye+&ZORYD4g>O,1&B<&1>RJfPJ:;0C@QX&GR_-/bSUA+G:@b4&?8:1-
#3#QQE&EL(aQ3d_]+2ZPbR/PA(:68T;P3P1?Yg9UY\V[,b-.abKQWAOe#:f33I2C
NE&RFU8:Z28CdE@S?H=;d1a\<_311<V_+YA/2ef>XUGK])4IF/TZ[_f(c^UGY,c-
/JU:K7VQ-]NXe70-e/B]e+\]4D:60Ng>&5PXe,a<T[UNd_=Ag&&)<SUCPY_IeAfa
#/(aYIND_,12d?&+?+1ZSLSC\7I^>H244+\RWJ0&ACc;NK@X\Ka]Pc#^:8Y34H?^
5[e;UQK:+4#>\Ug4.G5?TJH20UV]M9f[g2PT853ML,eG+55_@PMJDO=&Y3H>=.&0
-;L2/_dJ,1.OO_UBa_N#,gN8TYFK4TW508-A>KZU7ID)N6a&?W12ZF#,RS8B6IVG
4=WX&B1&@M^O/$
`endprotected
    
//vcs_lic_vip_protect 
`protected
)O<IggNNOQ.a<6D,<ZUYVY,bAO+BZ_eR77VQ5daIeYLU;ac\N9&K2(J6+J<c^9,g
+L/fH-J+>RRX=Kg8&]9;0@adB#[A5BK>FZ-3(HC90?6=(DaG1IK#=c&;U-U->@VB
E=/4NRH</)O6MY7<Z6g?G=(;EZB&-U3H/d\a(PEM_,6+[=5AX:Oc>cH>Y]2PcV:;
PPZ3^N/H0?T-KH/R^-KB\-3QHXd-Q1PD/Y/7DG(.+91I<g<;EIRB?M/-39RX:TPF
_1f41MPgA?GR72c;XQ18F8LC5P\\E(ER+4E0ZV4[fX&dQ\e6E\]gWE(VG\-T;cZe
Q2)>KSWPS@S7D+X\DP@g>H)D3>8dD(.YcLRK7A)J=1dQJd,TVIC(+:5WR4eeg+GP
OSVaB.ALf4#=-+c?VFdM29]([b4Zg#^]9=K[#\1P3LNESE4L1?K:M,1:g15HN2I\
)X]1WM<>GSQP6WHa7Q3]W2Z^YN\)ZMR=GWdgOL?<eZ=OA1LGQ8GcD69I/@S&f2O=
I_JU^FKb1-^VSe2)#^724)CK)AfV]NVXP0HOMf^d?7<2OI5M3<Z#370+ddNM02)=
:2&)[^-5MX)=9IG47@4a^QWSd(fe\MW;ND20OebB[GLQ?a.CWBYPW=Q,0([M9XC3
QcY#,NEZZAJB(;OZ16H0FP@^eRcOWD>W.;NeOYSS&R0N.]^]@9&<+YCA;LF;b5(d
D58.TDX(7ILM)/63-ZTV7S?Qf6d9A7T,AQ+,<0,J..=I[EBB?R\P2@<0\3_97#_A
[)A4baJ,>3<3e^\aA<FDATYJ?fDB>0A/J_Be/Z.HHYJZ^eC\8,Q5=]/#AO[c>]:P
7MEX<K)dM943VLRE4@fA5eKI@3ed\FT]e;IO-P0b,WRKdTe[&/f#OA688[RY\SQW
3[1BZ8PE;e3\9R&=K9Ic7?#c(/5GF0LD+a69SBC>(XP9AX:XQ\^UIK:+-]\+-ePc
f^\15B<f<T^<NSg_GHPI;3g-(Ic5HaF5X>X(:fURF/[QC1d#U2WTL(Pd6@bC#6WC
g+TRLJ-=&6<@?CaKWBdc>=C#OV3SDIY]BXHV4(9NcGfDA+AXg/18BLaJ@U;cQL]U
TGXgX<,CZ0(Q9#:M3F[OJ3,6bWNQN-5C/GR+c4GBaP/B?3&?&ACYUR5W:eeO;XSI
ga;H3e;g29-?f3Y=07F-D/+TR4Ua<E@M[D]>b)NbL266+Wc7P80T8DKg?^9/@Qd>
NMKDTXTSGYL.5-H&b(K:8Q,=K,Bf:I5=:4;QYS>KR/=48fe&09[SI]>@cN-IBK^g
-?+aL94aG:XWT)5fdJRR_AY_)F=[8P,Ua)gF6KQaA,@P_2:>0\X5/?b?D]^<>EL^
4_W;W-_VS^;]]<INT9#@NZ+^WQ0Y53T5<$
`endprotected

`protected
C3Z5YX>_=\4U=_SN\@Ee4P#B9ZEVJLb74[CJ1VTN;T1]=:1\If5_))I5\eaQ0cII
L?ceUKgM\?J<L3T?CNS#f#c)fQ]H_L43=$
`endprotected

//vcs_lic_vip_protect 
  `protected
?/gK6U[=9f1:cY?eZ>+][NY8M@Cc>b[Cd.X<@VR]77Ve=U)E4M9c7(fdW9=gb-dW
=P7fZ[=RE.d\]BTW[V42fbDGL-a.CB:QaXgcGe(O]bUN,egJc-?QdS-AaaQXU?VL
,B/WHD\c\ZRJ^M-e@JW1F8I@4SdPc)D?0Ca[H73^&&d,8I?NK2]8^#B4^ADAQ\TZ
MgSSc,8I)06,ce_/)dd3JW5\3SJ/1DGW:=\BdNWO[UdFM2-/cA:,(d:W#.0[Y?9A
DP_eZD]e7,Ka9#4K._Lg5E1UTT4cO]V?5H[_We(_L2,-SLJC=&9=fCG\==_C[JA#
UCH8?K3W6T?G^N7a>CbM1Q)5_TY]-g5A27G71]WXgPfK0W=)M@>,-2QUR&(RR?7e
,fW@CCdR,[Cf&&/<7Jg.,ceH<XeULZ(KYM]b))ES:A9Y\57eW5J5]#S6&RQS8J4g
fN](IMg3=UgAVPTV5bO^gJ)YE4gdH(\6(6Ig^I85B)Y\Q0G;&#Dc?Y8,?+52K>P4
FB.RY5aL8]KR:[O0X^@3;:9R<fW7/<_BK..8TEFB;fXBAVd--?3TJVF89UNf2O>\
1TgcAJ/+27b-P3DYFVf>4M.W:QS+8M8R0UgS]QAS(#2f51ag_I;[IgVf@/NIKIB9
XX6+26QB:VE(4=ITE.G>1abH.=N-YLI]MXSXP5D?9D-))7=MIGCg(89aKG^77(W[
a8\UX7e]aI.DG]&:QVF(SFGbV.21Fd_LISUKa[c86O_4a(Nd&52;[)L-&\3bgT2/
g-66\Z..c,?V>/.?=fJR\@PZ@=?FJ(LfFZT2K>?I.2ObVYR[KQB9]UDd_;.If4E,
Pa<M4eM;Z/fHV(#03T40CA\/(7ZS6T-Y8B2-XB>_6-V.Hc:@&YQY8[&@&(VX+.B(
U]Uc>VWGZNLBS>^#J4ZPX:PUJaE\;/24a(8(Wf2NXB[QI11A7Z4J99<=OJ=C+UXO
K<=GJfa<4->:0f6aBEc:Q.-O88UVNM:O3geM+/CW6LD@T.f2\B2Oa_0#65AW>8H>
R&FCcUPA:(>AG]\5>^2^RX8L-9WC@LOH@D67UbU@7_D#XZ]d)IZ?UKSeO^X5U>L;
&3G@)[)aJf#Vb<FG5aN-GE@_,-+WK;SZ6ZT3(H;f#SG@bKgdK2Xa+3/9Z^2+[0bf
U;/Q#[]a3\)YcO)+bGa+3d\.Ff^/C;IHAgY:SU=&^[eI6Y)XFA-(7NWgJXJ9J(G3
2MK;#[&fN0@C9?g_69Y7C>MZ2_#00QCAfINedXLUUX/YVY0<;E&(-aXC1DBR&YMA
9VFX5dgaD@b7XHYV818bNY6d0FE2;EEg)g7U1G?-WV<31&[aDFK76:5U]#4B@K(d
Je-&<.PQ(-]M0WLLb)<\dYM=ZB+O[La&Fg]]9H+KQ6JDDGU.FT7gag]cH6P.UU4O
=V5T-\BA4G&-O&-TOHC+g94Q</5[W)F.8PQW#<<-L5841QY(bMT9[\aPG4?#4d(L
(HKR1RSf5TcfFAIgA0U6;&QS#fU&?I1XdEa\aYL^O1@D.+IYC#g+>?9QO2ARR#H=
YH0VHAU-=2Q&4FT-ef+,:RP&Ae1M4G\&UX)<FT)gYdI8]@#,@2DVaLD24+C\]=S[
a4]B4@J(d-g7JUgQ:Q6f26dX-T(H[SQI)/D1MF-(Q,M]&,U;60&S)+;.W;?N<>1\
cPG--^93R4gbECI:U;Z(NUD[+CE>J_U3XfHVVN-&8Y_e(>?<V-W+_B45MAQ;4V3#
g?dKHEEaS/#L,b-Yf^4_AdB)b#a08P&5\V?]O\87074e7BWaOU^^,MI]g51DSe-H
GEIT<TED2IHC9aXHaQVE3Q;R4UX:]3]PCDb]Y1J)OKXGF9\P-B)c]&f;;=U8JIZW
:Q_KF=AP6dadHc8<@V:e5;FL)H[AQJ8I6DX8R4\@=B0:Ca26D>ECd?22.[NVE?W.
ccS,c8X6Mf.EB=TZ#Ta[2MaD@^^O8+Bf(]b13e/R)PPb18RP/_9fEaJ^OS]1D1Rg
\FQd1^M=g(F@I@B)Z2b+@@^F&^&dbA1HGE,eH)WEeX\V&9d^.,(]Q@=-4)1UGgG>
/T7T;XK37@UWaX>PU?SY]DHFb4RPgU.K,0IO5F2^GbPAV3KG)=[_F)+#F)^+N)@M
NJbCFKc0WgZ.fVgf#YV+8PaNHgMF2RcU]WT\D?&_L5),J^E.YKa1FC;6NSQC:g^[
53P>T)eJd]0^aM;,fS/>;\^>^=C\^(KFRECUHY9.XA<d;#-bH\KfVM2Q[CcSJTV[
A95D7+Q?VG\cgcM@@Z(M0;[)ZEB5L,E;(5+T=B&XQQIH]cH,\U;=-U?5(NJbRR6f
9T.d7,S3HM;P1Q-;J&5YdNbgRMc-@10UG>+MJ;0C.0VT,\d7Vd=V:LTJF.B96EZ9
E^OO6V?L)F&M5,PX(_0eV_3@5#4gSde.aS8:=M-GI]Z#7V>YBe1DI?T8C+R(O0:+
H<cAVZ>9Z]315I9?24Ja:GP4T8WEY?-_MgXb8NM7[[(9NR=W8EQD742N+]7>8B#G
W=G]JR7^_Z6VRWgY\UN?ILS]P&aL).\9E;GUe/J.NFN2fM@b@C8GG:>.FeCO<fK/
=;61)H7_OB>OFbEKI/UbSH\)GDb+-B9degbVZFJcP9a8ZS;IgA,ED>)HM:4F[Ad[
M7CB3/C.dUFaW0Xeb)Nc8fa#6]Q-L+]&?<>0c6a&V0]9#^fL1&7_IQ-3D_E/HCcb
#K&Q3T/[\M\MQ>>NL;-@.:D79-]dWcUgU<I:YGJLBX58;eK/HaB-O[7&Y7-<9EAc
aLI,d)FY,fKWQGPHbT3=LZ6U@Y13[18<6;bRBDMbK21[S95M&V1W4)K@,\/\K5/E
WC3D-G>g2M-.J1e;g=P/O#R36;^HS-Y<73e7&cb\7^]CW^W8,\L.g@(BW#Gd4Kf<
4?J8NDP_)[NQT4D2R&MH#-]//2^4d[;D?[-KXL=Vb,TA^&?.6Xa969I8:?&;T+#6
BC6:^L<(UgO/R<HJI0cK@W[7g4:=?C8Ga2I@H)b\d#N;LJ9C?#@-RR8bTD[GKWXT
VO\[9HSc+LSS3J<\9[fPeKR_e(7QY[O4baGT@d]FHWN.<.feBYaPPSHSAL6<&IYg
18Z#/ZVG)CgXB@L.JfW4?G,JF+S?E1F1<^e^#78ZQ?;N,MYa/YOFU(@U_+CXR?MI
+U)32>ES,aVB:G<T:IB(fa(?F<G-A#)+&EDQ#8L0Z/WW15WPX6+U-.gZ4FHJ_8\/
Yb<<c7.+US\MfNF0E+Y^I#HV1APO0]^aM+,e;YW9&Rd4LM^-0:..EJ42(8GE-HA:
,b\ZV1S>I6N4KNXYBPH/RDOf]+L6G]MTTYO4/e+.)\/^&\FG33:#/A.+SM8=-ZXN
<BeO^,F,&[aR)-@HP:0T3Lf1C4##9HJJ6T./..JNVbVA+S^GSQN_<<DdF9:Oa=e?
BSYEEXR4Q^:;._]<>4aIZX+&b,[gPfAI]f+Q?B46:Jg[;WP.#^+AWJUcf]@(=RTR
3TRUN]CZ^VBXX9[;^J7cEe>_4W(>&=gc@f?@(T<&PE=T9Z?V33\HO;QW&\-a(8LM
N.Z[LOVVKB<<Q8L(.8SC>AaCT;<)]ND:?)GD\\]&>R4gM+f+7e078X+Z-TP9SK^Q
.bCU(F?M^I6^/#F]JZF+ZM>=66X\BeCT=:D6>0B^()[G;G2.?f\YGN//-J\JTMX^
ba4);JG,RYBU2>VbSf(Q)O]c.d&R(EJVBBYbGJg_HXaGF$
`endprotected
  
`protected
\bQ^:<3C+]#U(g&?ZZ9=M#D;Q]FH)DZG,A&\)@0Wa/8@=U45VZbe()=M:9/]#Mg9
;GaNRR\XW>N8XH/=U/X>Td<SMLXO74E@&E]@C^(JV:>2Zd@dH[X._CG)9CZ1</cCS$
`endprotected

//vcs_lic_vip_protect 
  `protected
9(@>VS[2Da&JRRfQIA..?D>Y9TK0/7ED3\UK8Q:JYaWKe<Zc29K+((&3Z:B7O?^L
MC/B\=A7&d0P1W+;,W>?-^T6C<ZX3)Y)44XN-(-@c\GeEYb?b>BI(\7=+b(O50N3
WVPbR>daEN6?L^b8+49S9];BgL^I@G?+N>7R-32GcJ:[YI8W;Cd3K72H29JCLN=R
9@FX:EV0)M>@0gEM>#>3H8GdO7a/;@aA_S8.AJHP@cKYS)+SN6b&RO9agTcS(1)C
1@eQ[[ecBUE10/T9>a<C9)_L/HOgQf5/N5[Y-Y3JgHA:._2ZDY,\egJ&3S2N,PSP
dHDIPa+CR/RMdH9-K:aO97)XJa@e7>b3[D=_-TXLGSOUM4K(I^A.W_[Y8HK9.L\7
G@CAfB+K/PEeGVKKg),/B\R>+T1I.=P/3JE1B]U,b=P&^>KRdE,Ra(7Z#,I)Ye;a
cTO]YQ7Wf3,QTI8D^M?SYVfJ<IfXd\=29E<-_/Rb_a]IYO5V6f=3#=V^:Q8,3\SG
L\K2KN?GQ,=+GY-[NE1&AHgPYQf]NJNDGW[#<>BUAd;M^;?3]g=E04NP-V81+.:3
=1\:L\\T?c[60TX(4-eG6^?;DR6K+MP+;B6J;Z(PB4,b:bDO^LFW8+;4<)+MbMG0
8YL\E4QbP>Oab),2d[;QBXVVKI-(KcWPF/WW?(JZ[YLCfe]IggECb&99\\8;9\EZ
\#T=;>B3IZbK+X=b/_5/1311?@[F]PJeF7(?/;97#YXMZ^MaH@WF/_,VdKfBMLgO
M;3IRX2-LYfJ45V-,VA[3Ld>IDOR-]-,6#cBa]WCKVJC+OA/QIK_Tf#4?\cE^5V/
RY7(E0E)P:\D-G(H(TZQA:X-2?8NeF_ALdeW:Ge0BLCEMae;E6@ARJE8NM59:bbU
1W1>(=G]WM8#b?4E6=>NW;OW?CSVHV[OaNfD<^U21QVE+)2W;X<CA6R0RSW50]M@
D_W>CNUZ)4_HP&DM=d7G]a>JdfZ&9ZQJR-Kb7Z&/1a\E=#G5IW;5/F_3g\FX5<7O
H>AY=EB(3f+SN?PPQKRfJ,3\,ZV#D>4(=d^LC7QAD25X5.>1Dc^;f0>?^OPIWc6G
=RY&F=])f(@)_=C2)H5@LC=U#[6+_97RDGa>ZKTYK,:5D7>?DZ/9MHO;WJfLd,FV
>:89Z).WD&&JWP2EOA]#/]:3L,N@:H<Ja]-RF6K[g7<T[,OCWDT/=_PK7gf_.<;:
&^b6M=-ON9e&,[#I#J\+D+bc3,X9?V-a?RC@_f8T,AAX\60U2949GCe.]K;=e-ea
SW<.4G20><&96Z(>9^CA&2bEV.eBAM6_LV\/Z[7KF;=:B<1;OXICc&TGd02:&bW-
dLg)9ZaJD+3?2_IO>7a=?4I@28&T;=#+8XKZQ+S/)=f8ZRd0UY\99fgI(RF?)4a6
I8HWAF^_16T]GFC-J.3;6OXX[C?]c=S/XgA32VGX&89V3@N.Ca1-,A)LSHJ4L04\
\dKATae5OU,A=N7X98:I(W^I7KMF&@Z^#8b[&)dbSR/aFA@<HR[E^QVWf:/L8G>>
X/(L\I8V<Z8D>.P?WCA>2O)9cLZ\M1HSK.&:0HS:^6]TE70C(DNN[^^HKSRIE@R^
X\R6:8JG\>G-,U7Tb&#::?NUR53BgO1/M#?AI3]/C8ZI>/6](+D((DM.Z2;YQT,6
;KZ/e5N+P&?L,>6HS1&)186J9V98&B-68>ZT5MJDE(>#eSQdT:bO-(?WT]5M,(#E
Ka&D,g3Ic0WfEg#d)D\+QU0DF&][1UdJK?2e.9YO38,BJ,]ACb[&XFfK5EaU]]C6
YM2c,/L(#g^DVe]JTXQ6d]869(2\D2+I<XE\X])>/MK49TD5,F?a7A_,0=QO6NN0
ONaQcNM)<d.PL>[74.JOLFC?Y&.143/3U9/=DQ&^_SCMd64S,:?2.1,?=b,/Mg9)
S0EM06;KKHJ7J87Y/XF98[AI^;-WM=aX(&agdN-7\&T9^UKFRHd.f9JCKId/g@-<
X<4F10-=1<V(3>3>WGC4Ob6E3g@NAOT18?6M]d2#(=<QI_Db[I8->@1=-Q)F\&#b
@0DcWOP/]f;Q&&fe2P?AR8:)P5PU.Vb>],S+3H[X@SfEa]83cI-e\(Nd>)(A\N)1
+O?E;08aQK,FXH@^FfO>J:f@>7#^_NaX.7/WLGLL#9(<BJ2XJKI&HEUWDU\TD1NP
_5CVJ5T?#^F<P@F^/1<[ecaS&J\5We]gR+9S#HV,<EY4K(JO0TS#J;@gD-Q@0e(Y
@>DK2XA\[0[dUF#)/a00RK8b8Rf9bcSBTX:O^+IA_+YP^E6d4BOG4WYf/=\@c0gS
2GIaSDg2IG+]G:QONZ6GbB-<SEV[#NL6V38#1JgSC7Q<C04_);c3[&&g;:D>=>&?
\dRV&5d9]]ac:bHe+J@#8RcASM]d5L&WcY@2QK#L6eN<SDQf.3b3M^)=J/cNVR.I
8L7)B_8E)2O@-<g6^WM&+3&&aO-CVC@a^?<,ZR7>B<PPJH67c3[ER#N+VIBT:WF,
gGPX+c(CTVK<O2-g>5Cfd/.,D_38&KVg;FHAN4C98[G)0WG.408/XH8NEbDG=b/N
^X.LU5SKFU^f#ON2WAHZb+_1dNd=;3;5Z[3OZ3PXQ[gFP+IQW-(]:<74;L<>]bA1
;AJeKCgV7.7bIeJNTEIDX^C1)IW?YQ]9IEc</)a/O).A_;,LeM/W?;?E.5>2+ZeR
\b2dJWPA4gA7C0c3Y=5SIX@0N\VdbT-a7T0gaEWfe03;8O+d^D\T7e:DK/M1>JB#
>K[OA;)[&)YWZ@e\AMF2S&/[D901[QJ/P1B0g[-#;@Ae8?T#Od;5:4TIf/M(ZWFb
7a,,\VaR5;bLa9I,B>#<SU&DY-HW(TZY3EYf?(EE5RY,QJE#+=(BX#5[E..b5;V_
NM304JaYHZe[6&7Cd4T+bMCRX0DJ#[[[0VL4+0SN?HT1BGW.@4aYc3R9+RJd=4=)
2R2DX):bAP-3H_c-?^.M6:(^AS2_IMa\/AEO5+7+SO5@VZQ6W/8Z)<W@L]eM-c0G
c51(I.>RKUZNDfc3FaV9XOSSX5WYB)Mc_]S(g;>PMI>PA..J08dGR<db\cg/CEJe
eCT2G9K.^5gd;2.4C;JE3VG2H9TSW[0.UU3Sd+98RA?O2Y6):bfTHXE/:Q8SU9Pd
V@gb/dD-??60+6?-\-8\A9@NeOJ.D-5C2L99V:5,;_?IAP@be&J(EW0JX3@c2Q9Q
_(@>eF4eS+CSG<P[4&&@9G2J8Z6VKAVdd,9,PM<,WB#a_cHP5/VM.c--\@:#J9GD
^E-9/IM-/EAb2:aC-&H4#_5/]_HX3+G8]:0RL<,7,6V6M^DO#c=UYLg3=8\9P,f?
)2<e^56+>17>d]CI\?VOM(SeO@Df,#fIWQNU2Z/^,,RPc8#(+dePBX)aV98\\HH_
:J=9X34K)V4R)P<8)ZC&e-/Q]3RT=_.JC<#UU46<11\;F<ND=I7914&?6S6/9K6L
LaaY]XRg@WJ2@;&[EJ0f5Zg3UH]^D9f6N#05b,9C>3)B/1<a(+S90fP_[CRG+;17
27O.g<R+4NQfX+N9@=W8:.53TOL?B>[J]aQ\\>FI)b;>87]/IdA:ZV_bfJf]ID9,
6W.Tc=fXKR[C#GE#(S;O;PWcB:GQJbe(8bb?K]D]NL3F[RIg7>5ATGJd,)4^2e>W
9+NOd1L#T.Z1?B6(3]@)GY421FOaY-4ZW=a5?9&dKXQ)IRQ7QL\Q9JU@,<>Z47;M
T-QVgH^@&#5)7RQCNS86_]C817BL[#@]YXYR>FcKYHZ[ATcaO=HA8JPX^gX6\PdD
W34]2A1^P89.\gISHF5&+^EM\Q23GO=TUa\/+Y1BeF>464D7N;?9]dH]GeMP/GL(
.fGF,)[>:D&OP3-\19LGNZOeNX7.]U-(DW-bT5N)_4fT:JTUV=9X\cGM]U6&<YfC
Y4,EgZLSOKcZ9UOb7NUJ>#V3M1?2N7c-+\K;E.U;S&Cf;2)D8LVXEX9ZRGLTd#IG
=C24McHM+ZIdUHP@:YF#Qb&;K&I?BfT.DG+c6V^g=7-UULCR\/Af]>=C/,I(gN1J
N&V0O(g^#aC2#LQ5M<208.>.25^Ic:Jg2-+KV\\1G/7(8DD57b?gc-c;(OYaQDAA
VDWP?^T4#]-?15+9ROD5:ZU-a:&6WJcYW8-M@<c7/4d8I&3>7.Tb0RKRee#Oa8XI
bO<>9<#c4==MC2@8)[:c)cL)^c,fT?RF>B:4.NQgCW284=[:e+/,=ZBdWDL5.d6_
e/WcbWI2515[^c_a#bWa:3&FUFbBIX/bW.F4ce_@:bU8P.W7:C+(-U:2]KXX84FL
^0fHD2g+,Ba[U2&<9</S_-UC?dU/H&L9Y/_a#-eQ)BA<65=D<>f[+OFKTT#QMB/a
G6\^W)VY,19?gc-e^BQ<2=D,Q:Z8Igc,0GJY+^W(KVJL_QW:_Z]Gac@T=U74P_9g
O1(OZ<P(gAW#D6bV\A9#2fZD6JQWEANa\#KX=:X6V6W,F:UU:<c1^Y.I):a+?da9
NJ55C4X,K6]I1^24Ed1c(:PG>:B26?ZHcgSUT4)PCZ8eXTGf(8#OMb@-#S[BUL9+
M?gGZCP/8;_//QBC+c;2Y.\+RNEA^DWGXWU6aLB7(a^#5)d[]T#.gUAcUZAe=0g.
(/M.PEH.,RVYIJ4;WXLd56J3OU&UeEDPIJ(Z5HRdX\:1\#3ce2e[(7FgH#[>aNHJ
0)fJJeB_@ZY;E\d3(/14:d>^;\HeP:fZ7XcD=BaV.>9^FdQ&F/]Q/T;>O4SW>.3B
[_]2K#F;e(6BVK3?aS(<=LKGb/>Xb<D^#Hc#:/=;E]FA7L)8A+T:2DR5//L:7DY-
g:.Z:dNJ6LBKYE:68:58)[G.L=YcWg#D:J[cOOe89VcdP1(@&Ib&N/fJ@#.OP(Pe
?H1J,L?,1#BNOS-,&<T(@<R:@d2][]0IL0g)A9X#>[S@GH[BJ&37c]I[#e+X62,e
@_O3,T;[(Fa4:@4_<KNU(bY&&9JW+Ge0g[;fE8)8PA.[L6T2,+N<Ne(g6=O8=K+4
3.1F?,4,=ZJN5Pb:[4)C9IAeA\^eYFZZ9d3K.[IXd]OJ/Ie>\8@/Ca5=<_+fXCA)
eQ4c=64Fb<X_JECZd&7Q=a,OS/bbHN?cQ+37agW/PI4f=SRU[T1RJTG.=ge97WJ0
WFVPL)C98&.f2<)c#^]\P0P9dFOB2Ce(5<]TE,&R?SXT3P?ZQ(7FagE01]>c)AE]
aU09?EASWC=UKDXCfQPa._F+-Y:Kaf5TfRRIK5cWV_V:K_2,Y:VCVZ(SBCZU4YSW
P8,Jf&WTEJRMK8;Q&IWbR&I(A]F;F.KI]PJ4UM\&>Sf^:d0LcQ095SN,d7;-DQe.
e5SVfEe@g#LDf?^6>HA)1BKIgZ2,)D(M,,QLN@TCb^^I0_.QWG1@8_@RDSS_,YN9
_RR2^&-=]Yf(Z1TR?CRP\Ld+?EZMTg1S)&K-BZB]K)b7-NR(Y(;8E4(-#g)E7)@0
g5T\:9OV)N,+WfFUN8L(bO&7UWaf52S0;3c5)eL28E6WR]G&X0Z=<U(=aF9+6S\E
_Pc0eLf1RPP,\(>-Df?^N[FS)]e9Z<b.+fB65=SK8RO;a05V;I.E:a)Hbg(K.#55
+.3E4F381eO_bIWPBFSL&@);F6<:b/P&9#L9,Z/1D9BM5T=b^O-PMG5N_/M+7U.U
/(TcBU2;DNS@e46bH\Dd;=69[_@C))+dQL=[a9\]E2C&#ddQ>::NfC4bW):>Y3DY
TMCd7ZHEeN#MK#EcJ>>K2MB&ebHa#XGaOM#(83OCS]]GA4AW[7UMR:R9.Y,_dR#c
]g#>HEW+a\Q=?F:K/R-MKD@eHLOBE6YHDb<YadUJ@EH;;Mag2,4,4-fK;A4=3T?a
S+9::f].?=aS1H,JNDSZPDT4))BPH\B0b^53_:AB5KgeV1ZK((^]0P;/L#Z:NJU>
NFG2SU::)UT4eW+DJ,T\J.RaV]/S>H?f9bge_Q11J2^#XDYG0&(^U=>+)R?+1/V(
EC>U#+C9X-\&RPB>YQZX\(d^@gM/A;>N_PP.HTQ[?_];>e3HJ2e+M<4gQU,92fM^
3d^9:Ma)W\UgeOb.)5P(BHL\DLE5X?Z+e2XWP<CUd=T]C#APdYVH-7a^aXfAKOB6
KRAdX^:R@):MUZQ-D/YTAGCPe>KY:4\]\>VO=;&MN9H[@XQP?+A\0+Adc#,_XOPg
acf_AL&RgC+V4PVQV&.(3QbK@2a(@4LV]L,ICScXQX0RYF1(>WS@AOe4[QH<e&R+
a-_DWAW_KHJL/=2>0/Y>.&CZZ[F\);+A+#CaK=f4(P1fWJR@(aEQ10P2[-22&YSX
0Zg[g1aW2>[)^bZ=QOaG-)f+f153QLA84S8I1C\8MLG4JAf-J8]]1fdD:N1HU&&N
9a;4(38,:)Jb=&WMIE]#AVB9.B0-VB23g\J@[3E)D[_PeQU2KTG>VL9#:8O;_Pa4
U.]V1DBHWeYfXCQFT?0/fYSYTQV[B6AAB\.,b/aXOM/O^G?g6A1&0<\0)^7I.KBH
PON;G/K&<AQXbC&PLX,G)=R##BCE1YV#LG(/X/JC@c]+>>&W__ON6@Z[d27]UO]^
<#bVM4EYKD^=A&O_;gQVELDe04BJd.S.@@:X6X?]Q(>eB22AF.VDM8XYV1SX5#eI
@^SJ11:>FZ)8Te@WO5:\Z0W1S+&AH;WY+PL//cR:bY8dYB/1\ND]5:;@Tc1+eSd/
;#GA78Y19^\&@5H@_[^R_G1@P+8&(7V,UD#AH@\\CEFV]C/de<aD:Xe7?)O=,0>8
M+YT3Y2X3?.:9#C#2(<0]Qg)3Lf1@EGb=3P0P,U>BbU9&C&QBA&/81-<[)Q:S5D=
DIEPe7=;&f6VWWPbP0+-)I.8PEc^G4XL0_(b^2Z>@GSZ?&<,Y2:V;(a)P6UTAM9V
)IF;&@.5Q</MCKJ.,f0-/)R7MaIDF0]0F-Hd1/=@9H)^c/PJS/74/W_?\EY,^[:3
CH528/bXMfG76/N-I=9e4b@(2]KZ-[TAQc/bc2#>7N85K//B>YBg.TV0eU\X#,Q&
Y>-I@Q39ZPc;1cK6)Xe_.LTcJPPPM/M4TDV_>3]&A_d2#5<&/<(+CbW4F/H8\)4A
+?3;7BdB<5^9e/#4AE[.PV1M)N2c:\c6>/U=GBb&7S.W6HJ#&)[)7LWY0-JW]:\T
G>BTK>1WY7XI+-Q1WRV&.aX<=]:[0&)3<QKUFKEWZ&&23O]\e4._Fa1](;TZJN_D
-&Gb2Q(+:_8ZK@bS=4bGN-)MRVWbCW..3-FVA)gBb]XJ9:_9]BT,]MJ]e2.SX,ZO
XDZcU1VK71&@.#OW=Q\G_81A?Y#Y#8URMM5)QgIY667D8<^)Y<CF#G9ZUUPGO[cK
2YJY=):#ZNNB\NQGX3bF2E+DHc@dSX8KOe^4eX3La,(fdI:#DF)KYSFOB&N-VY[&
-PWELaa>58YM:R5H\)XG[R<;IbO)2?(_\f0G<<INBK(VcR)a8T^&-3@#A4g^2R&G
aeRI@R)Le2\\H[V0G\3K6SDMe@GGVCP@X-+55=M#/AP)5K\baf@Ed7+:<-F,dK.C
0WI]@8VBW7Mg&d)&b:eGCd4BKPf^5B@2fga>8H>S^Q<\@V>#ST1;;F1<5D)C-:<O
HVQ?&.69,:BaIf/P)J]\R5O]L\23)+#dC3T&LE#DeC&IYZF82:f09\&F7H[cYS#J
8<<g;^_e8HD<B2_g4Bb2Q+A_[X&c+K=f-402ZFU)B5H4X1[f<EcY:X^-XM]>-RUH
,5SO=7PFa[6020dT]ce>@2&1ICS>_EaE<7dd,g>&)C/HN5Pg6]SH<;EJC5T,+.0]
1gL/Y^([Y^PL#X7Z_7VP0cC)RU6eOXS-g3::bb+024c+.\+4;E]Q,EUTKEUVUWF;
^gXcZg7:?.-b2RDLA]#FJX.IY-fGfe=Be@L1f,?R+X8G17(SRgVc]=5X:f[;,-D6
Ffc+IV@6JX30aT5SC\g.)bPJ\5fE8GZBSS]0KC:5HVC1LGL#ZLLEO7EGbeeKaA+7
SW.,]JT9@9>RD/[aNRSO9GEdL0>TESF7YFbfB0fdI8O+Q0.9SM?>#,+g<&b1UYMb
NZR/5f]062T=^^V92L4QC3,OB[M05LT(50L#=\-K>/?dT_7AU1C?<&RO#a#VLI<)
b,OS_be;:ZY[IX?42R3Q]1G585KKT+P0UAG@2^C8NE+V=9.H4FGJ]0N)D#Dc(W#L
GN0IS)F/D,];]a/A2><GIgUJGHP8VeO=GRGQI1:;87_FNS51PR[#Z>edfX=\@6,O
<X.=70f:geUKdJYXAERQ/L_,W.R&8[B-GX?ZC1GV4(dE45_LSf+_MdgaQQW]C,.4
#K0(Dc1/VE+TRLcMg4_#9@@D:-+C:5O:9N2U2F5.>=RI\6WD#Q5I/bR:4N#b6ML9
f?)U:Y.R/EfU/EDF_[3aS3[UT@aL[g0,WF&ANCeB;+IK@IYQVBWW+8=YTcRIVW=c
8UW6W9C[B_XX<4?YL6-(?,H\D2<Q;LC7+&Bf,0PYITQ#DXV-MBeBLX@c8JfT/7+-
1)G.:;H2#PeR?\Q,^6ZC.eU/OLGO6B^Cc^,7NA@/dC&XbdQMS9Be92?CI:FRU.1[
)OR309Wc;E&+b:M,R=:-V(_:YNSUP.e^X/WR]W+I@RR9e[C&ZU0J-HcI3[V.E#FT
^/_=E<bECDbZJ&&WDOW#EeU6D^;ALg14,)gI79PEKE:3G1X6YX7@Z-)93P@5fa7O
]VNK)SK4.4:XRbW^B-VQMgO0M1U)Ag=:-K,IWWE)5L+:US<TYGST2P8T>eU2O53@
Ce5=49gD6])=,;IX]9Pd5W85IJO_@(;P29efT=HEa2Y.aP&:6eIc<B-;=>Z.cVCV
]&S6^WB3\4U[?;B.6YE^(U(QSU#a@.GX1I\,W;X[9aL-4KPd#V52#Rf-9b9.9Q4[
6+Z=.^T?f7eMDT^OY9Wf8EV6;dE<S7Y9IZ[XP(76a[X(g[0X_F=^Bb+gDWKeQb8c
eVOdc5N+^?]W/?8?,TYEOU.+:aVZ(M_d2](?GS+0AB51GFdE58/Lb(>]Hd&ef+c9
GaNgd\Rb-YW<8.fT1ZU)Q-297&R(K<OC&GJ9/V#1eVEI0X(8dF:S.g_4)=#RLRVH
I/Z6P_Df6Q/&?2f#a1@SO_AC3K2B]FO,PKJA\+PS(:4.[0->?\;PE)NX169IdFR5
eG1WHO/M(^XG(0GY&-HaY8eWDI<^QP:+[R9d1E,Z>O/LcI0TdP469AYX+9Zb2CNe
8D>^WBH?0XI2fJ2S-0aNQM8&])SLEbcN:U(;-1FB8Q>:a/0O0d@WUR6]M&]RF+<1
MXQF[C\b5W=_:+@&_bMK/0+3bO<2EU;,.Re+B\B9f:P>2==a@F)-XQUSJ4FJ,5C+
f.>?0d7_>&(-]CYKZE5^V;>TAZfbBb\]31\#-=L>e0+1>A&-RO3NJ-Z.;Q4CX5#0
87_MQ/^B_?(QIQ=<Ff_N2S^)YaQB&K9)KH2+X]9aD5)O#^)H7e[6e^P6Za>P)]7P
Q9^[SD6+-@W1Re4HC7?:VKd,=X?g2+G2TW@X#@fS(6]&HV:S.<bf;OGWQU:1N&W@
+7\+d-.:ec+9^Df^CN.7^GeJ(4.A8Ff/7M2CW0O(Y9H-]eQT&YGI^=9Q>aC16?Zd
]?gDCg2P/M)>^F@c_S^[[CUGe](-4aL7HSG@egIAHT<UW&70fe0]52gXD,,K9S_V
6TPTD,1>gU>EH&LYY7g3]NLP^cZ&J<b9O6V]_W=Aa(dcE<F&36L?[&0KN(^#>HL7
OCOb<M\(]+7>(.\g\M&5CKY(V(OI\bBG980/daBDg1S-7,_(/@?3@^/O&gK;1GcK
?2/T=K-#.C;QH]9WZV/Ud(eRdU=9TO<5OFJT&Z))a3EdW<1]9]SC\AIfFJ>1WNU2
S7,VZ8dWfA0S]6O)J?\S1SYW,Y0g&,4G^+2AVLET/>-&-L0B[Q.CEeFV>3Qc?(R^
U[C2S&FC3#Bga;TJ)A[6(#0\,(VE>HgLUOXf42_RLQYF\G:=-8\Y1?O^gOd8SW0&
D\bW+,N4BS?6PB;gZ6&FDZeRKGG?E.fTSR(YbZIDB-;Z6VZe0[\4\89/WZ-BQePB
>TWVEbad=c68eP]G6CKJKVC0_L:K3Z(QW/>XXc-3L5a#.Y:eZ8=eTF6,\ER32X,D
4-CcGT&,TRM4;5=FgN#<fM)Q9Db();edDM^gc4c.SJXKVN7a,2FC]Xa]JN0-1I>L
GT0_PVV+:A\Z]gE7<7[7CUgAONTbg9NM?A96@Ra-Yg#O+aM=4CTLHH3<QWI4\[[R
)3^c&/a395>;M;Dg8eO9+Z7MTM&eVO8_05TU)ORS,fM:D5M?[Z/(9/g5=F,@CgW5
acSHI@:/ES4>-=bW\7>bW:J-)LQB.WM_7=b7_\b1L_dH9EDHaAX5VFIB&Xg\?W^U
S]RZ]6GH]NBG[9)I\c0XU.,+,CP[E=#W6II\,AV27:7Y?XN6Od0eP(FU57V+J#Id
)g\2QaO[eb>e,bL8ObWc_3#1,TdE_/O1WPaSG,,J0PK0@]AI6c^6eA?4)RP&;PZU
(P@a>WgIU2ZCM12ZP81+#R&K9ZE=I<bg/^W)8EO;@-]WT6_CZLF\4\K0cDUO8_;C
]_8+66I#1XT>+[7E9-=.ABTUfcQ)XEaB0W[OS<?+-Jdb):9dF8Gd\N^-#?YJGH_I
HK(V6RC=ga]&,2],<9Y<#A74W0>3-87)&1V__3<P.-&ReU7WV4=X>#TSRG<gMGbF
,b\7g4R>R6+5HSZA]@.WEba#UHR+FVA.a#6T/cGH7RQ>MXc_V;&eC4^8HB.@6R]E
;3<:fd=<-T?gYLd2bg83-O=J,0-.KN&JaW;>:d6d22Y&@)[]TPYRG4:R#fXWWF0B
^RP-V>)\.gSb=NML+E@-7ON@K+PE\ZF^88)S=7CF^JgXNO27BDeMJA-]a\I<8I=_
g?F[fX4f.\gJUJ;V#d;VTd,1+SGLd>#8J7RaT[_5Fd))CCU-0X;KB4T4Xc_JSaY<
-;gTG#EaVa;c4D;C+?8eG&a:/N=O4eggU^O,^DDTEW-FN^[CWU#,f4_<ELU]YNA^
\I?P]6+A@#J<9PZ449ZQ-:;=^Z]:+XCMP4CRA[f3c_/,0AbJ9L/;;N9U>L1JN)f6
B\Fe3\GU_A7eQb?>P83<MG.SGZ8PA3F;4<B=84&T.AX:^<-ca@@2^(S:CNV_:/Qg
Ed;2Rg91QC\[BJ\B[L7)AcTVZXWJ=_(\N3>E(3&FS([Je8))ZF3P^ZQ20M>+T,0E
ISXbgSaAV7DMA>ga>?GM<K:V_GJGDJ4,XKJWDfT+e(8Z6gNP<?W?EW(dbP;63-H3
/?JMZT(aA3K6)1WFfC,B_0R;8T;TC1BA#L^?<fa0R,HE94^(1DH2eW16IB],Y=V6
aTN]E=/O\&I869D)_NSF6a)6>(N^)4bcDNJ,:eQM=SeN3d6&NS8\XPf1aI=:_QR,
;A=b0[CK;bEWH>E>JIdY&^A)>>/fLAF1W:)99ZUT#32WW1L3b5(RO1<5BdJYIYXB
<+OBFa)W?[Q??b04K0=MENSXN2aC,;3ZDY09Q7Ta,8M2L).U_,K9A<;L[bd,64U/
dM,S?HQ=g<&P]:7I/&JBd^412H1<c[cU&/e<IFda:[8>A<HGbPHOV6Xg^5F\2)+d
AX:;HKb0:O[@E1HaQ8@N)fL;\-TQRGa#dK&EbQQX1P?-U@d+2O@J2FQMc]+XEgYX
QH>IBMW0T42<O3^6M1)A2C.<):Df+/IHZ_?QPC,1=>Hg_RDZ2+UO=<?4?Ia2TZ6+
QYW<&80A0S8/,NH9?YI;-6G0J?+M0_EgIaWC,^EfU-NX[A>BON333aLB(YYHZJV\
eW?-D99Y&3W<(39Q0J3]QaMc)c,7N6UKBK)Ta/:0#1_<:&O2fNXUI(Ff1D_,Dg]B
RE>ZI&=c[Sg8._A=@]]2@7=+3Q?98<K5BB3WBed=c4P[V28=C9-THM)UOCH\:b7W
+B(YI\\VBdIO.R]Hd9ZSF,2e]DS]N]_J1?b0KEbF2:F#RaeeORUOON.^;S8@W8)-
-58]3C^[fHbXgH&@98L_AF+F-VN\E37U5W]UM+H>2)#a8VIY>/K7-/d0=9bG_bJb
\_(0ZMKZV?KHgC;b(]CV4c\W(KXQa2d-4L(3RH,A0X.COWe9cR6:P^V2PdcBOCR,
7dUdDUbd9M+8.T5^0Sd<8NS@9b_G@f)VcEO5?f.AEcT>?Xad7,SLCR>VI(VZ4[.]
gFW3L:TW5c-=E6II8H&PX^(0<2\O7KHNHM8TMSGC;X_,9\8b6aT^1;dfEf?<Z;7;
f(6R^9QU,UIcBTJ6M?1B#]XCD,U.THWZF@/UK-e/C+Aa;)M?Vcc.8DZ0Ja+WN^FN
KN,3(K@M@(W2[P_F?<G@XMI4g8a_EQZaKP+JKF#7cNf9\EA(U=W?e&F0ccT\;Q;R
-Ba8<<[T?#ee,)Ab7,V9]g+8.[<g=]>;JB]NAZF:M]HBD>6?X:C)I;5)PX>GfDAE
(-)R)<HRRJ17Z&Mg,,GQf8T#(SQe4BAW>]QV[NG)eJ3gcHGG2/U-O<H^OF3d5C[5
feL=d?=CJRc0MO^0EWAT,P8<_N6<J1JJ1KfFcBI^T?LeTe-?G67KI.TfYTUKeggK
/8A[.b\E6f=3VA]b:?f>O_4eaBP>gX1_NDSZaHA1,5P:/.OUc^54fWffF)E8Pc?L
#33C](D&0SF_S1B4[9PAbS]MZ;C1H>ZH7P1<,FYG2/Rc?[M1?E:#1fLA[BN4J3&(
>\),VaEIfK6Y2AH^TI;&7g9D^-=+XZXS7&R@Z=a??H4+H8[]YFY;I<P8SZ--U3QX
D5;>>6f&Q62Y</EZRB6CY?LIPBHBDLTHG1QO=?e.X6OFO]2_2OM+31@aJ7@eg7I[
20VC[Sd.U65KC0=Mg#)(.]2@]RO7]G0,^cNaZ;g0d7P8A2X>,>CVZX<eYQ3;c@?)
UA0,&VD+Z@/2b-Z],,[UMX^JNHG@5DF]HdD(P[Hd[e8^61N=Z<^:fd?O8C._3:X/
QM3cM<8N6A;]bQ.F=QOcIdT6[.BOK@?R9[];0H5E3TC@I.K>;B7Y,?Y0,^,4dM,A
.[IGTd\a,:g;WdP@4PJH7g39Vb]gGQ#^7Ia?US;10e+fQ8g:0;BD=&dI#a,C=[S4
@KCY&=c-M-X@EY.?Ce3L/.QMT+:[aZKdH.R.^4LQ6gd(McAO<#<-0Ua&=@cgfeWT
9S?&(>FUdY&#:\F;8Q:HT[O8_#&E/APcRdFa)>LZ[>F6D\2b672P-J7?bIH4geVA
566(>+U@c<NB.7T[cTEU30WPDLQAJe2(dYP<^+_Q\RbR#AVe()e<#J\B/-:6TgWb
-,eg2/(W;:ZGOe(FONMQFN1ZN6,37D_W5XR=DCC3K,QJ_H_D8cFDYK8A#<WAaYL^
)_]D3XGPD2&B)?XD^GJef-@V+GT68@DL8],+,7(c1H<bTCPg@7;UY],46dH_2N>^
=?_.F]V.S/XOKFa;)UAO>VA(43V.^0NN=0eBY?])K0=X28(2/F-8]MPQI2PT=/a4
>&V8+YRb4GH3)5SLTI+>X+WJQNg]4X45O_0]>#\S[QK8BfFU_0(g):3,P<Ub;QFV
#;TDH<gc_M2^VV?A3H0dY-E<dYD_V#Je;7ACDTA[#4327<Sd...V500L6#9S@e.(
Y5:F/4/0CK(^7C<8\g1XJOJQB;M8Q6C+O6OYMV\][\3LeJC5(>NO\&77U],Z]S5;
/KLC>AV.A2V75CC8G4F3IFd))5D#W]]b^g2BX@NgeXRBVJabD1J=#7=6IPD?7@TL
E;>@dK:He-0RQJO:LM3d<3RecRBJC9C?1d+=S-+0#&c7VTCP-d_G,T#^)#aD09cC
\1dPQAb&L58H81/Y46M7SY=;-^X#fgf^CGC3F(CgE^7Y:Q\NDQHJHe0-W^57:)K.
RTR>^B6TCQ7GQaGYf#G5T@#dZKE282cUKI6S>A_:44?K,bGB#R:^0I]eT_EYeQQ6
5#;:2e8.[_K[KA[S?+)TDe4WGEGK8+&P;9G+O_<:\YTVF4WbG4R^KC-Lg^7=e2KC
XW3-<KCGM3b-]7Q,?c(E7NQ.AZ&Z<9>:G4cNaL3Vb.SbN<Q:)HDH(5_G&V_Hab(f
C9UUZ><c9bX=1bDY1\;D/V,#WA)cTRT&4)58_J1.\OaR)IT4D9?;OI-[ZZV#B20N
9]JbGY>P.eT.,/PHU;GNSL=OD9^R558:2-fM8BZIcWAMTcD<>cDYG#TS\_JS,]&f
1KVK^d_VV;,aZ8KWLD,0IRK7B/#FTC#Y,RcK_\XW944L1/_+(0F>MM[HDKJQJ9\L
Q_PW+IaCQ;0X4;9ZAJXb\P05(FV3^aAWNV2,4SAZUAbSf)2gRYWE_cA],?ZP6:4#
EG3a_#dPB<\1F8J7U>.Tg_D(BJUX&0:/D&;GX2B,K2cI>dV&YT.Sd1ADF?2WJ>Y_
bTcWfVVK6Y\MFLf#WTE\+G/XMH08b-G.[DI@,377-Z_O,GFQS46?BCY_Y#.IW6]C
P\Teb9_+,6A2<ZZaOMSZc7M/C,@?YcA8gI0eH8ZB/cMKP\6Ag944&Q&a3GD_/F)a
8N#OB(gER7S(6\8HV7I,=]D1U7&<LAWG:,dR?\<O@4VUI9H^5##+;FBZ_X+HC&;a
dd-<LMd)>S-6SUJ,P,(6<0e9C4(E=BKebGQX^GY6[;AZ]#-+P34Rg.8=XT05U>=f
(T#OLQ/?9K_T(9T.)GCM])=4NfcfFX@EX#fS]JN778Q8&a<.#;,fB;F\a4WV\#<?
S.GM)RC??PZ9J8Z1]a+Q/K;dUSQU=\[ZB,(RS^4Z3R&EL;6UBN[W6)1\UbI#)]=e
3,PYU)R<DCLQ^I)dL]7R[CUJaCGL6&O)Jc-FC\L]-F4[RQE9E?O+.Z@Ze2=aeQc3
Q-dK.W\3M#[_.4BdO:IQVBDS_SD]M?D#B,Kg1LQA^\8(N<>_7Q)WCP3LOG?HENS\
LE=X9D9]1T-[/CJ89QG>(We7F6CZQ#FA;K]f\7XZX+GHK>I?_.1AL@a_9Ef?:VM,
CUCfSObCP2<Ga537YZ7[S,HaGF[.#UWOgdP@?2N?E9J1)7V6?4.C&8+]VRg_G<4C
2JD>N28HCW[M:1&9/>PWP53L1#&D5P2(U+EV;2(gZ7]V==e,N5F16:-XKRfL5g:L
XJb]d^_NU@S8?]3-1Z,GEbZ9;C[e\(\_CR]7bJT[(G+A)I>7f1BbbYfR>B9QW2g5
)[\Z9]\48DWSAT#?OgfK1Gd2)+R?[<_dgO_;.:K:YNQA8V@OKI3COfK&E;4B:UHM
W,AbCOQ)V[@_\RU)K;NJ#NN)^b>X<.W<+PaE<;Fgg\<-d(4LBA^1W30LSXP;F9L?
EFY&(JP0N;@7FLQ7.?MVaQ0DJ+.@U5I=e)NJ,<@e(IN4&.36DJ)6JGD8J0]BQJ]U
])9G,@@X(e59<CY_f0:He#0NDcQ/&]S8GKfVLXH4[BJ6+F5fR1BW;/]RUeCEI_J.
3)Q;,&8J6;Y-DMS(P29-X(7f@DE+))DJFF;XAYD_RWU8(7A]^a#+(-Ncd_]YR1VC
;;bNO[_HPL207WZRUPD^;+Z54BRE4].>SXE\=@DKf?XSI4OU2M3=UL(cBd^Pb@Xf
_N&<b=.7W(9KI@08/gGAUU^A32N8.PXeSMW0NZgE6^0:C7Z/G=R_cb=>JHYd7(SZ
)\2M#N5?SST1]6Zg(Y]cQL9e+9<b2\)bJ<XQBOgVU2<+[cP&,FV9JE=NJ_5[?\;:
:C&M-AT;\9:DO9_GUO6O,d;94(&^\;TLX,BR&A(A#]3bMA2YCX#aHH4U;7LJW>H=
fR4Uc1YbFN2Q-V2f,Pd,5ba5<9G8)_DS5G(JSKc4QbEHdM&)G2-HA.&X+R=]G[5^
Ra3f@>Cd8IcUW+Y5FQD<&-><KDZV8]&XG>J-=^D<W(K06INRQ\>@&dTQ>TFfb\N&
8A?#F\Za_+EeU#g,gg(AS]QT80MDH1T@R967.#W8#Rc\+WZbdF/&ILfW+Ofd]J)\
E7Q\W<.7^f3MGSJd@#^FS\+[X:Zc8I&S60TX2&?]2.A).K\5&XcB8#cL+BC(\[;@
A-WbWUZ@g:?_CJ25-0U]@;P<GP1eb/DSZ<]O\)[fV4H3[<a-Lc[T2TS34M8@5DUZ
3?ag@I)a20FU:[b4Y^TEJY^T)4]FZX\)@@ag^D_b>(EL:LZA\IEScKJMgJ<5H4WS
4X(SID]W.:DOWT<g)6YU9bV&=]D5McDZ9e>GZ9PCL(F=,:P]::XW]-KKN?2g#e49
;D<gJFM/g/^eKJ<e6JNP8=/EY&2PfG_T#g]1d7]E+G^c4-&E80e8QceENaeN:PA(
3-)^L>X^/-4^BJ1IW:M\]DYUA):XJOZ?fP1Q5E,=9\J=(?J_3QJEXP-M<0JVNDgK
G>VagNZX6FL7b[MbH8d+2ZBCJV?Y>>T=AR)0/KY^S_#4+Cgc0<(,Md&L?G(XB#P_
b1b4dP(Xa3X6DL9055,?)RAG,NRP#-^LWK4][EVSWHY.K&?BSffg0.M&ED@fGIS]
fP;d47K7\L[V#eE5I;:JBFMBN1V#4B?:4[8?TFC7@/)B9+ZaggUY@CU?(S^8T2J<
8N[R4=RLFPGf>T:@g_B6\A]+^I>SQ<HGH>,1@Z):G-FPgFQ???JOgR2JT_Q4:WE:
[&CZJ\[>9;UUb5STID_;\:EH,)#S<)S7K^eDcK-HNPU_C<K/3NX)XU^QUL7NPVUX
NbQKYL=EZN@O_fg;TW1Z0PDbZER7JR6TU(6F&&MB,2FOc<;K@,X;\W?SIK_,dD>6
M?+?156f/-LPbd5^8MP=@]GTR]gH+:6A6[-LD4TA:_\LTR3-&4CX&T&(\BH,UG_6
gQ4If@D6/\Yc+UDEa;^?QA#e2LO:B-<31><MDdEaPL1=[Tf26bGfR[&H5B+:HGQ8
.EEgWe<<\07QcY)IL)=@A>SIFgAb4.-^_U>L=NIT^A7GH0eUU[67BgLQaZ5FS1O>
O1UJDf0RW=)D0YN->6HfaJ,C<\DB)>891W3EUd5G6#_4MD2R;>GE;EKT(4[eAX)0
+6^&\AM:^gGM?Z=K.W\<;cZ<DV:0AGM?XPfcQ8/Z68HRNZ<W(b873YDG\-Z64NNF
[QF5SAf]@UDPUZQ0TcWH-g=]B6/+CW.c@>J[(3+^NB]JFe2OQ?P<_?1da<EF4#()
\C=4(3RF.UfG8SfVVF79;YV;;7/0S/L:[QP,.G/_e+a=19eIA0b/[..ZV#C:Z/.R
W58FgK@J7PP-Ef\SFI-1T\8(-cNgB,L0K1YW>d-KS62f8/U/F<6_G6.DPT3-D#@P
fN1@\9(f(?@F;KN_395C--3TeR5g[2Q\dQI/8-dW3V/?]UQ.X@6Y--F)=&F0J52S
Xf<g^JY1La#b:WBFW+C1NPN1T^0?g2e^07FeG,IC3<I\e70BOE>LN28>95_@51)C
>09aJY5RK4DA./5F7ea;>[>[Gf5(6a:Y@:J-TY2G&>^EV]MR^\(15bG2FRI0R/BM
Z?NT)-](4=bIOXa^^.cA4;X^\A_d5<Sb1+[5H:V2M3H9R0=E&+8II5GeSQ.56f7X
<=d7@b3_]4@F+IZe3TgRS[fHY5[>L(62a/Me=3b:2_V2bWfU#fQf77J3_D:<2<Q[
CP:KQ&-3..>9XLOHRI6<./S+TQXEB;][6+<Saa4/D1N8QNYA::EXacF(M.1?QUS1
39QgM6WV6YF13bV5-@DXe@?&P6f^CM7NY;8E<_6\NNPK7fC>4N(D=4ZIZBddJf&@
0Q2(e8IP/>HT>EH6UcTBC+fPB14]VcSODU6PS?01.<;JgO)(\V/7[W@P<.D1>D49
9>dX?DX9>g@9)N2;dd-H7ZdNFN6W;fTfY>+I=@7V)Vd?QEA[D?4]-E^K>PD;_1)>
,O\])=,/QKJE4]-?ZC@ZAY.>2#)XLY=A[)2EN[)9]Ka+V+I)Z^235KT&;JG@77A<
\C.K_.E<:49ER(fY[,EJ5BI+?97S@=_OB&a^154F3>Z_\,TcCL3D8^bALb.2B9@)
:6.OP?EGTOecdVadb27b@PV=PQ/d]&M7;V[H\I^7N,&bOP,>#Ee6&N)O7S;^TI/W
@(CN==P:7?8@+5OBD#]&ZF@\+3.G4=?>\?g2Y)D_\EGO=;U3/1e#/:4&D)DE>&1(
?]D@6&#51DP<_DVgCcfD_^O_4^A/d63\XEAH\@T:7W@O>C,S,@;=I;ec8_<W65Ne
;JaH+HD>cF[AG??d8/;+5&+\7T.(Z-aD?f>OcW3-Y0D+HEI9SRRDSd/f]X[].Dd/
bC&;UD5a72@CFWg;[gfTdeG9aS[?7D8daWJ?BT2K>8(6ed6Y;ZW+58;c2PXU=&B@
RZR_9CgW?4NEVYUD@PMNSO)HZaN3AT)W+XCUC9.XVTfS;RfXF1CZAD5E&]K4/8]H
3_Ud_35Y(\SR<BG,IQ[#9D4G[UA9Z?4ZPZGa5g0;LID[XTT7SWbWH.ff.e1ReA1Y
I^/e4;dK-QVbREQ-OYe4\GBf-H#X(\YDU:GI7L>MKcC\69SY8dUB3.P\8TLA/@M/
DJ[aDOTZd[aJO:;A]3?@9+g1X>[cJe?)2?UbaUC__X)cV_-\)fB_?O82aDTX<#Yd
]:bHS9]NB->3CPQ_H&b>](W;)B3f]E)NPNE;4>\,YeR<J.8Wf63TV-5U.DSV>OXB
8-=UR8KHFYf2@-1FHe>gH3XY,]AFdLgAGVa<(?2?@@MdG;;K/W-NCF7,NGMQ5Q\B
(a7d+0[/ZaKH?P\KQYVBG5)ZZ@FI?<=N@\2JN/f&7O-C9UD[OLHE.N87G8GS)>aD
J.\f[B31KO)HX2VW=O.LF]X;Pf(4:QSa389d,N,FcW;3R4>X>Ke;SFYL[c826-\?
0GJEBW,?XE27^Y[3e.[5B81ZCNg+UI?CY=f@d,?7J)[15c]-8/NKJ44V\AFI)cG^
SB=SYH^+N(McB>/0fKX--gA>?\P0]/cPSX>C4-SgKg:DTY8Of#g:a:><A(K[gLYU
^^HI.7,F-EWCZHR:?J&>;\aXde&JgD(b&]-)Y;DF00Z]G[1bMeHYRUgDdRB,:BE/
.#cR+Za:P9CNS(G:e&OO:^QX^fW&NBMEQWUPEH_AE3FV7XB6OU<2\AU6,>/Wb;&^
,+T/I?49e9BReD3-T;@,DWC^+Q[#5Z7)5U<UZOVaH/?V27MTN13edW=2DYT=cEN[
GbN_+8K?7YIP@5LU2VcDA57]3PG#8Jf,5K>#KQ)DJgJWa#+Q[W5;3O3?;aQ_W)1\
I7])E3T8>@)f1N(UL+/HZeQT=D=V@7dTBd29PD?bQQH)FdT=E5,:0DWbXH[P.)D;
T5KTJ>3FeN?LTTgW9<+]Z9@15&c]P.T&W,/f>gY;W4Qb6^^N+Y,[C&5F-:#2&98&
Z.+UWNTO-AZ<5I7BE^GeLTcSd7fSCHIET]E:5]Y2.[CH(OcN>KD_DfQ6AFMQN[29
:(H.&FC#;<D)WL2(;aF<D,QHCH>Q1>AM#Y721?OD2;/0A/(+]fF_,D6_8A=-TTcB
4S_[4_SfEQ9E7<0>^2V](B8IPTY)^JQN305dTDaLb_<JX(1R?G-R5f-W95Y(9DTD
-D).CV<FRI4M-[PeCUgVI^VB/P#[JB96Z]I:HE=YMAE7a:ec.5A;.NL1L&cBL];f
)3.\fI3TCS-Z>fCOK_5#PSV1D^[L;AGHY#<K@P8IZZMF5@SA.NMKOdaEDU[]^b0-
ROa\DJO,e\FFV5?^TD+N#V-<O2FF2JE5(X+WgPYWUV,<Y6Q0PL:/\F[FKg(3Te8#
,&6ge=ReW3(gZKYQ#U6,\f+,V,@@EKJeSg@>R3H@6AICH#B;PQL[Z:#eBcZC+JK6
A5:IW1L6cTEL&E4==aN^)/6K9Ua5a4HIN:(3:ZfgJCcJG&a^JK&LXQ3aR?VS[8>(
VFTd)S<b?UV/C^W[EZ-4b_,^OQ;Yc4HI<b(cYd7<(CNe3NIMTScN7ff=DbNE<B]O
RaKf1ZUTZ:c0^TRcOCfGCGA70^OSO4c0.be=@=58&2bcRTM::&176#eQY44Xf::J
,:g=?V\,NJ+=c^E?3-Z#cD>>V@TOQ:BR4Y<Q3&L.6_PVRgVNd+=),43,HHSF6CL-
MXN0)6Q;93b)dS\40QC4QIfKd3^;8V0:^5;A,J=>S2NX2WS)_KF1M\L0#?Ngb(-A
L:7Egb>fJ7Fc1X+7>Wf,:+F6RZP#Oe<B_-&.PK/JCAR+>S]ABcW9NI;I@/?W]]44
5,[=W(O4g)CaW;bU._X3L3Wd4fQKYB>JC)+)^?7WgaK1ecW5Jd2?X4GOEZ[=eM0g
YXF7ab(.eQFCa1H\/WF\A/R3dFd/GD0DU\DOPOUKR7VgTQ\HWMKcE5GBF9J-d;_#
N9A;1R@<F=VYXTS2WOJBB_)Z/C:FBb#I6A(2dcd@FNM+@I)g>35-eKf<BdPR=_MF
UC=9IU))G=MUWe=^81a)[P:&c]^TG(.#WbHe#AIM(F#?1R2X[bg#;(J/[MOME_>C
;Z\.MA&A@NDFX3VOSP[T<MI-N,NP\2V)7^Y-5-\RYEc+]38,Q4)f6Q^XN0Y7a:UL
I9TRd^,8849aS8N?=[GE1G+e9-G4>7c1T&76b1D_]>J#d+11PF(H3AUa#CFRB>>?
[#2OTOB(NQd(HL;SZ42)R#Y0F9A+a\c29F8638fK=-3M<.@]=+3TEO(B+@XdQYYI
&,,+J2Y&Fg-^BfFV8c_@X6-MNJG]Rf(#XCbe+I(1HfZN85ae2,Xda[6:E\7\g-ZQ
\5)>1<d_2FA3+1R)-B8))^#<F^X.LR^?F3;@.FNC+^=5/[Z6(=^#D(2KWZeCeR8G
&Y8J0+HfI555U1aVB&D4a4f;18I,gg7Mf_@;&>G&[BL>U\5(\QX]FP0ZL+>16g7.
<.RTb_<-78[[8Y.&W1D[dN&OUgBL&aN5XI<@cUYSB2\\@AT.D0/4+95ZV:]=?@M&
bU@#E&e#\+eYCUf)4Q.O>F(/4?]B0\02:?:(7HW;GDWCaP#GL)M3f<45(D?RHVI=
-T/^J\:EG3VZ>X9/a._TCVY2^QO)#GPI57E8DR,4OG)E\/KO:=L^YP>9^>6.)a#O
5\Nc)6-L1L7<ZQSK1X5L--M)+:6(AL.GV8F\5fH?=6FR2H,0J&cK#RK>V0GB]QMZ
70C59e7QOH,bWN/#PXGFW+bbB3)eY<2E@_+e>K+H2&,+9Hb8,#,BPU+;:E(Wd4YZ
Q2=f=.98fS8^)+,Z(MAF#XFA0L1IVg9)[:aeWG&gNg>g@8cE#a:=C2J+(c(&S[Wg
EPS5M1R_YZ\@e\e8+8(LQbUT</8CBO&SgAba&FN(&3NcLdGEd(Z1Y?63M7Q<TTLP
#]H^<6]\?8HPI>)9F9UF+DW&Pe-RfeKR#6HSCN\GDM#?G./<c?NS;(@W.+HP@cM7
?3RJ@)5@+TbJGgYG-VLGWDQd?O:TPES.-NV(A:N+9BRIJ#X9FARIed6BYH>]T0)E
02PXDZXJ:SI,dNQ@0BLZ@>-PPEOeA0JKBL[D+4Q&9C0<S8F(/WSV.]<LDESTV)M?
B0;3GR;1AU#A@Q(8/d>B32#@I.U+e\W(XF.R0MK]W^B\=ST\BY5I@g8W08)M7C)Q
7L#-&-fLPeYVN2d3,9R5P,3\OM)TV2e(7gM+RC59E4D\;[KFH4b\EXK(9S<Wdb8P
[I-4,Pd?EY4ZC88\gT@eg:39bZB7.gT)#I2H1Q[Y98-P93Q/T\3>b@OT5b)K5,(-
7O_XCLW(ZI1EN\.L7\dP;QPAUSAcX+SZ(&c[Td6TbT@#d\KM\E,-d.+1;WK[7-:9
81+P4QK29D(a?d[BV1G&#IN-\=.8VO+E,/d3\#D8G?68;>eaI[H4H2V<6>+^6I-W
_CIDWCU;K[GAT;Na@WbSEJFECBaMb4O77WgeJDa6JRG^-cLMO[=&-8^R(TZ5Z<;C
S^^CeE.[33#WWO;2DTI\+V_#\V-0+H\]aI;KHZYc.=Vgd+WfW2a,QTIgZURb2,.P
.^ECP)dSP0):EGR@V1P4<&62B_0(&g;bFIG\+5K5:2[(988U480>4YFOTHL6V+Gc
gP(XT\8&b7EF<<,K-Xg&?cQ;^BYQHC[>37Y7\1:PLKE53f(LB-\<-Hf9M2\PO?Q[
?/4,Z,9B+(:/:2J5/=U=#aPUc,L&OXE,Wd@3H1(/c&\7Af@f6Ub#[c<K3;H2UBe5
1>/\f0?;+aYLRJ=;cU_C>V&6ANUcIe_RD.JY6R@7Y((,PM3,DAW>\T@WV]bAPOWN
.;eO_W7>-4VKKUMEfW?27MPL?TK=8I#&@)/5A1IW=<&-U+4@\<LXP23Se/+FdbcI
<eN.F7)Faeb,=U2H-JYY0;.G1N_b_]C3L5S<+&9STWGKg)02J22[C#Qa).(L/deN
CY0XA]e=;^;&D/4,:LFK)b(M:)2]=IdfcK.8G?=^Z#HGb;XU,;4H.3/5_31RX=D<
&N)B3^;X&D[P#F.g+Q;V)+-X4H&f7HU44F4CPPd3RZ43C6JR73GX+L&D;DFI_VFP
>FZ2e#EI8DdM[W+D]M@KH4=#Q4a=D4L>3T@N/KWU\RFX,Of5@7?7Zf9=bIQ3]\g^
]@]Bca8-\eI_O6J-f=I/&O1?0L@SD4)U11DQ+)-XcXPZW=/VH_-QgKG;1&ebSW?<
9WaDO&Z[VdD@,^_IC5XaO&EE[C3TKJf1[T,VQDT=I5\I2>1O\C]Y^6[J)[W#/VV-
B1ZB;[Y2HdY//C.:9F)A7(-=]_X:#GL]SQFR-R(:9=+44>gM/>f_e>7MG.GD[J.e
(S0f2;<eII1ZQ[D;KZA_:8S\DAbU\8)b@M4cVK=C4,>_M32?R>_=HgG26./BNA5,
J]V;,^M(O,2+@;BG1a2HY(d&5PRfFEeW_Te42BRX@8+N-O\787#f)P,+Cb@;9Z9[
e9?#T2c++9:Y3[H&L9ERX/<J--Cc[6ZMOJA#W[:TF+f[?V)80;W@4;[bNL@J52VB
YOSXXGW5P<V_;PP>[9&M-T4S]INGRLf<BP1R+cG-aYcXCcAM6V/(;cW4_5N1JPP:
Dg^\U,)RB,a<\[B:PYV+8e.QHe4=g3\f/a&0.8BZd^fafA=bRGGBODVEHLORMG_c
OD7+#DcLb:I8fQUKb12dLOe0J@<ET8cV?C0KecAebA4Fg\=cRZ\c1P^QR>)K:Ib?
&.S_MLZ4AEaEdD3C-^CfK<@1CPV7=/]HR=<4I.X_RGGK(Q/(X>C#e:_He6^K189/
F(Z46Z(U4SNfW3B<K;\0Q(+[@3Ng8J\&:/3ZVe>WUTCgC-Z/LTcH1KS_f^Y.P:.-
[VV:(cE;P9V)D+W0+EK74<AQY(W829WgK@QG\R8HC+3g5cL+VBc25V(G3C0/8#LP
.;BD__ECFNSEU:O4:_T<[8D-AB23\[:QJfU3C-bP/b>?@0K+K@GBS#X.0E,E[(^#
JZW1_7RS?PQ>2D:2D25;.AI]57BDN\N[[.>N1=^D0Mdde_IdGIPA=RXTSVMHAD@.
O^bcU]c?A^g14-+/I+HG699PGE>L/b0(;Fb[Y^U;QG,=#>YH6+:1/QdW1610P_:S
HFUbFR/>G;8C/K<52V];#NRJRPFN/[dX(La[](+;08B4.I-J;1P,A;&8980]YaI9
b[a(QIYgR:I4JSUa@>0<STbaWcYbOG+9gM;Q#O^g#6IS7SYIPTDa\df?.I<V,Z27
C2,5/MIW0/ECAC/BA3[=U[40MM0Ye<)4[ZT4J98W1JN<EZ:dY1d)8J&P,\5&30+A
dBZe2>T^e>BD4QB+6Lg#,#R^LT/YIT?>.8B>5N;H^_6aUW[f7MB@\P<8FIXcG+F.
YHT;XE#Ebf4g3^ef0.5;Ee<>ML1a;+>2>5B/W0eWSGf41LYEYI5GOOf3F]I/-c,Q
J\a7G)HKRb=Z6.)5(c:V,I3a>@:NdeMcK]--;/BX=WPa]^^+[Tf4\X@DA1K5NPZ^
]C=,0?-aU\6dH3XBJ6WNg)bW6WMFL>?LWTHDB\:_@SAA=c<#4./1TKB&/-94UR<M
f@4A,2ELf:b#WREXA72P4-YAWSZ]4G;0:L9Q7Sg;PVPW<BY;0)d5b?U>gK6DBBX7
eHR\SYgf5_4<A8&]9@LX=a1XZR?H=7Z^\KRbaT2&AOcASO=)GV8RQ/a:9,CUbC;_
NR6g\5eL[?e.QfW^F4#EDC33LcZ]a&g:(CNSF<-??R>A,WSdAH(SFaES+a0(>F7S
W-5K[M7+#TJ^UHC+fT#DHMPcYP.Y=V8XS&fg+V=M=XIL]W5(\NAYSKZFQNS@b5(E
&Z[<<&7][g>3+^XGec&+4X3VT,aCfa4^44gSH0g+G\HDXG_V&bERT;EFLc(HNHDT
Zf8#D2Xg.XVWeL]QOA1<@5#0bQ/Q7.[9,MR?Nd[#.#8G+7DQQ6BORH^.f<-fIF-:
VBe_K_[3NV4-KUf7FSA7ATLgBTBAP&G6bAPAINMXLXcfW;FB[\2C@#IUK_[04Mb0
faI#D7CPD/3:=+H\-LSe]8M3;G#R9[NfU9bR0]C>.1Y-:6H.HO6&^g-@6^#PZ+A@
LY>):NM-TR84CV.\a6X^(P<2O9+T9DT05OReFKcgV8-66-&YOafMHE.Hc6KM?V1W
?Y6]?_F._[4.IM)BJ1>7f3,&6-DM2/X:>U_Ba01Y10595-H\=QYD=K0_f^>]F:;M
BdP&X_e^Q:fBQ?FQ&?1^HJ6(,9;^,O>-PEg\Q0[-[8MY.IRJ=A1;?ZFSQS]B;^]X
T=97V#KW]WOb_;X8?d&Y\ITe@WGE07)CM98_WPV\0>@V+H?Jd3)BCU?d3&^&DcKJ
f71X?R_=I4>6?6.WEM_c4Q0X#1N6b+R]>LNX.VJ&]RT/2=c(PDdgQ&CSX.c>1/K<
#EGA_aXD^K/FeMPYT3]&gY16gbeOH0N=;a/K()b&cG_7EU^F(CXDT?A&)-Z9>8X4
[?c;M_6L,G9#E0J9X?eBS08@BD];Q@gJfBY17D54AZ&1=:#:P[OQ5VFJQ+G[+#12
\7MPBV&@2FO)O?0(0EAT67L;+e@6G@Q)3CRX-PH)bAMBAC=NGOe=?;U\f,cTCY91
>F>b^5L3(U)&L=c?:Ia:ZF)=WR+,Y9MW&B8[INNLK?:E)2<IL_/]4(P[D@M95O@d
C><?K9C\dfT]XgYESSBN.Z\@T\A-^-\bJ.8f[7\=E]YbaLOGWS2;#?,/=+gee9N1
1R_bY][gBQ=[R2F0H(3e<7Ze71.X9QeM4SRg6I12)],9LL]L7)1.bc\^^IT9#/]N
6_EHY8V0BM.M+\XDE>NF;0Mf;/X=.F3(T3_ZZ&V[/#1b^+FfG,JS(&CU^##HDbE7
SI+@A^;XaH=PB<M4eJW<]bb41T6IAEcg@.aA_=NZ#ce46W4E5#H,M)gF<MBGee7a
M,]VYU9JO8aAC)Y6\=17=ZCI^[,Zb7V6TMfY.>@B]O77fa0c/K-Eb]@?F?SA@XMJ
KK+&L?MgZ5Z-.\@XN-BU7ITPAb2@U6d,<Q&0X_+:#]9BE7@fQaM&ZMZ;4f1KOG:_
<84(B)]/PL9B><\6XJ_cb16_dWON6c\dG++)d?P)Qfc<f1-64D\G&M63I4-;LHB&
U&2IK09>&Pff\U).e2D_LJ6CC4RPac@c@DWAV6eEJNb4TE<H,4U=\A#F2\ERN_VV
#@/7C,ZFKL2&E>=H_d58#08WbACI+[f7GLeCLOR,6fV+.O;LX:\G&T(S88@[X@f7
MHG4_=\#>XHS^XS87IM_CIeK3#YZ;Eb(L05_gBUTE;H2BW?R&HWG/=BU<DK:(RO<
P)]C=,<X-B86D:X/[7/3NQ:G+96.A#7RB;2+5HB[?c?<aZ-=@WZGYcG?KKWg>4>D
O:?VI.Y3N44Wf]A_PcW-F-9dg[0_c_U3:MP+0SKb?cB<9?4OS&R859be;XV5e)(Y
TL0VZg<OLfA/d@V.cYaJ4_:UJRGXb5@J,gGXb&?XZ7g#A77-[#>..^Uge?JNJeME
C_UCb\A^DBRdJ##/f7/Pf38L,YY2,Gd^;7?X2_?^^VP>BBE,BOPeM]8S[?)V#TO@
?>Y8LETG(-T-5+=gM77=a9ZRfHUeQ[H79^;8Ue9,7#UTd)W^eeH,RadPZe^7GQF+
;#BHSb/X,_+Z+XB)Z8KHNHU]dLGf+TAPA44NVD^7U^U91f1WQ<3gJ?A7c;?P\3fP
W81bFc6G:U&3P#G0OOQT)@FYL3);>_7E<eU5;0_LU=a?N0<5U+#61,)QZLD3MMER
W]HTMcgbWb_>Uad8B7M9N+PbC/Rb[(3P?64Q;c/]AQe>/V/;_O33QB7;BDS&(<I>
:?XBU_V_XeX_,a9DVN8/U/0F5[[JO)Cb#g[2_D<^RZ8ZF^577J7)E#DbcZb:F<c4
f2P:F7YXN@e^:_6bF,VK^+cNZ@F2\dSMcE/fbRP9,W]/bX06XMD^NfD-0.,QV/F&
&gA[K#DLN&>ZLLITd0,,.gOK<4\ZN8d^1MZ\1A=^ETG[Re/<f?935N,#/N]5d(KF
ES&4C50UT]a9c5<(g;:AK_V1DZY7#2_V4bJebeK,SKe.C\9S)MALZ:&E(gY=0Hf4
E1=+Ce(Cd)JT&H/a:f45_=,(T1ef<eK;).Z)ROb:-c]a\UTff66:G;DYJaX2b-2G
F@aSD)ZTUV+0:_OLLFJV#0=5ZA366Gcf0f_9K.R8c#f[?(4-?R9Y+YYRNfF:5OK^
?Y8-J0K^X-R/](A3cT(:F+7V#41OU6.CQ-CfW+9I:,1\I=a.2ZLT__,_I>3Y(#,;
f3e+ZNI\69S@^J^gba=C1dF#g/a?^-UO:=+]UDAFHA>P1TEX=O&\FI=O9K(a1=0b
a#<:d@1gQZ0WP(P-2CQ\:GN>b<K^-WQ>OS&;b_XHeeDP7X#R+7H4O;QOM83,:_+5
HGUZGc\)7DU<J:Yd>3g>4OS=/,DZb=EY-&PVT)/Y#<b[Z-.WXb_=@)0g1a5-Q@gN
X/HYTP^M;RW2.-_:Kc=.NJY.SB;4eaDWJ:Nb@X1=FR[^Xf^]Td&6D;E&6/@#2;>M
d8K[:,d=1L&KIYJQ@O3<Me;>C/e;0GTe,?:[D.cUM<BP@,76RE.F1M5?^WZ5Y:9-
XZOWg;d5N20FZS78K&/;A76&=d;b5eT7K^]T]6V/M3.Q4OG+\]>(QP(4[dCaTS;N
M_.a)^/f#8;).)L6I/3g,f+UNSF(MUN6^W[MFBe2-BQd+T?A;KJO81g7G;Zd\>0E
Ea#RHQ=C.\4=dA3_M8J=VdJ:S(EARYc@]J=2^PN?d4=dG\V:Q]UZI=/K&H=X.IIN
@SF1f=85C:K:aDe4MGPK43KR11[M<6e5SPQ,#Y,Q[17;3M@;7[c6b@c@fK=aHf5N
HNR@Y&^IMR@g^;,EY#9U2KQ?&BCW]E@;.V&cgWB&BTV#;G5+dFFZBAD/L?J]1?<<
-IBf.A2K,D=cf7e=83bC]\RFB>f=S6K+QCfV#B/)1eA([T.PZG[72R-I#J4LNF__
JS>_cdD6]#&(1NBM[aRX,.,&_1@.8UQS0.K7YIK(e/Ud_3?:][d;dXAf5YFK=J0L
^NWbJ;L?C)e)/0cRd,NB;76UF##2M8AF1C\[,gPV87@J2F/a48P^3M^5COe@gZ#X
H2a^W+C0fU1V/:5R:YSYN,ZB]1X\GU6;4Y]CI\1^(=9U\f<\D=TOBe,NYU-U[VL7
1e5FD=EY[0,V]_I3NXaL./+)3?=W,a1aFJ4Hc9L/Eb_<LWX82KG[;K4M;AJ?OJ;_
c1faN&O1)M8W1[UeBRdKOR(G;G?8QSPgJ:XL4_J<e.&gR]>(/AYb9V:O.2Y,_FTD
ID<B=WWTBCJL=ZZ)2@]IRG4;T6Z&5eS?B;b<8e(:TS)b<g4[3M?&).,9_B]DI?,H
^>OH&\O\L#M3cW-BN.OEJ/7Td:Z?RZWBCZcf&IBPMV[H3=9,S]F3eZ.I089KQbN?
[?@.9PEPVQLb[S_MVC)ePG2b/c\#G[0E_O>:aP;PS&66R?37[8H1,,GT+3YW_0[)
BefTYV(/g8b>XT#0\;MQUd4&B+RR0^T>_1@<XSN4YeC>]HZ8GR\JP()KPEcG2/JG
?,.J=^C0P/e.1D+&[(fEdOO-cLT(JJH/7;[R;.gP:&+):.JS7=._8\2#.5DWC0??
eOGD]1[eMP83;&)6/0S)UTP_fT>LW]\60NBeYf,,EOZ@H\B-R61V,8_aS)YN\R-+
K0MAWI-GdRP\C50@a/P,)@<b[9g,JLdAd5#+7:<D^/e272OK7\E^ZXX+]XJ6g,\=
^WI-5K.\)@;98<FCB)MZN274D>1+0>VO.LMC@7/NZD444b]fHGbMEEG?,;ISZQOf
;ReKL^RQMf=9#<YH-4.WcUJ8e90#58.Z.S@Y;Dge2c#N)Xg8O1g\#N:R9<]cg8P8
9ED+cS9cM@\:=FCW<c^I[-EcC57T&G,.[W],)DW3^.bPJ)HVc@=2W\:XQ(:b716-
7<;TNb096I0,<X5\QPa9DdegaW?-c3GecF<97^I5.IL0AU>19A7b;AdgH+FB-<PE
W,XM8X2_d@.MTaD^0>4gf1AT8ZS7XWU<YF#((/(X^6-faJfIBC&-T@RN3:?>E>+\
LBP&@2/@GaN0Z8]gA&cZ67JdaG.GMVR[<U54=,Z71K]6NX01_;_aD4a1c33NX,KH
FC]Gc^AYQ3YI@YC+=M94d+;H0E>D3)6=9Cb/gXJe,F]O(EWQF:(-V)EXf.5X&V@9
4^Zdd\WZ[a+;GJaWfA(AB&R[6++5&\[a>5e.RS>=QaMYg&R]?^f@S7,;d/^B=g:T
gJ1g-.2))80Od2\IL)7NFK&L@7BB2=;E[G#4I)@#]XEN7<=IgBVK(+^B<e@Y(S.Q
.OIQ@\X3LH5Z)Z]C>9[O])Rg^aFXf=<N89N:M\N=W]]a<bA\RVXDLQ>aELd[H;7.
U48W<S\8P-?_]8(RgP_4F0X-d>C7JNL4QBQd87bSAY/d2S.PYc4?F74/9ML2ga;G
CBP5.M/(BQ6Q/b/QTaNX(b()I4B;GLMS)S-O0T^]c..b5&MI4\?RK)[...ES).Xc
UQ^0Ag:=0/6FZ#2K-a]3dXNSB@AeH(C2F#Wc15N/DCd2Y7W:5_P,0J(^GJ)CKZHI
-F<V@,IW.&ECB+dUJ:V&6g@>8.f:4a<>bG6GWD)fb3Q3;P<<c(AN@\B7WNL:U7]=
)#L#8T7;aR8PFMb,15TS<K?JeJGd=F5f^/4;+c(RD-CY+ZCeYR2QZELY][FZ3]Ec
DfQJYGPL.G70Yd<2I0?W9T_AB&,XaPb>Z[ceQd:]ZHUQW(C6K5g^74?X@#c<8#-<
eB\QebVaI?N)+IHf65J9ONe8d6g&Y6Z&?4(a9FcafFdG<Sf;/E&)BX#e.Q5>.WXP
^X-8^D_V7[>^Q_]ADb,Z)#1.]>S.QYIJ]>ZS8b]L[IGN<I,3VM&09W,]^;Ib)D51
)?Nf3OFC+e#2BQRJRWO+G^2(Od03;TUN?Je1R#cb2@^1-fPQ:VHD5W;/N>=6<C-A
9R3g+g.@b6[6B&;PWAKI(E-dUJ04HdY,C.EJ[V7_3ZECRM\#48[SW8cg2YFGM@ZH
42VP/3Q4=+b3&e81-T9@dC8G3);K[5ZTY5<2^[/1@]W+.XTPGP)ab6A@7S1K8;M2
eKS[6E#FO(=dMP&-I;NW:L8]+/SXfF97)IDYOI>9TS^D#VENbF;cIbUUaG+8]fO5
0G/CO[,V.4(V&dRK<b)XC]#^.^]9IPAEgcSMRgcffK57dIXM7E5CP.I3M>5LJC=B
_XBL]5S]&\8G1d\[<3/P[.B/O-ZeYP0S&Wa.6C@-2<5IJH<ZMF3GB&c[7AP\P6>]
[e0\[^K7)S(1=/TN4UZ[3V9gP;5+UCO33_3Oa_7^_f7P<cRD8HSAb^g/^d^0Z-CR
V78X,RBA-cgHZfR39,6F7H8WX.EXSX;0:MZJ4CGB_R[BL;6c;7/GAc-XJ-H\9fT1
TL1:]f/U]<Ac1,-J7=-)UD5[W0X82\KKW]e0D,Y_:R+Pe[AV4,b^5SO@S;82PcKJ
/E=6+EZ)+fV-e7G_)c^6@aEd-[8;FCaRWHX5WDS7V>\_;5A1f;.-/+06+\06ZTeX
P@HVc[@/02\gKU2FEIX((@@#g+bII,&B_&-8J(6BS,>Ig(B8\[15#\g0aaM#b^X2
793VfMRWS&<]g@YLAE#GI,NL#[A<]62bcIJ::OS0N66[W&U/=6T?ZR>W2HbPe\]]
f6X+:)a=5B7BB?(NESGEMTbQ>3W<Jad/d4@XAW5_Ac6O1BP19=\(,1P1J1NR1NF#
Wd+QJ+K64(Y5YN+L@+VJ#dPH)]_DbXCgW.:XAcfPVU9_748ZOITIK82N--?7-ce7
[@()H35_/,BCd)66[^A[GF642;>aKABNf66>3Qd.0RQdeE2-WB5gT,PC/QM(A]Pa
8630e?&O9NT.-2\c4[SeY&:9^P0X<7@2VQ90a7]ecSf5aXTK^QQ#K5]\Y4^fVSJB
IW[fdIQ4?-^@3[W49S.N>>;Sd-31,)\E8gL,RQbU)4&/2Dc:UJP\;-[DJ+(<0#X7
PR#2\/L_7fJBHWF(e8\TT_3&?IJ3F)^]bIWGZX#[VI#PMI>H]#)1BBT;3PG8@?&3
-6dSO;44<ZRBJ+.be\acB,E,fY\)^56PRH:=_^+RN@?:K0?8YGI51Icga5c:(@4.
VaVUUGVBE[<I?[W).03LLfK,<R,BPd-RJM1:0=3:Wd?[7@]JRbS:(;48P?@,PbfV
AW2/+V^W0S9Mc\HV,HW0eaE)S,##XD(?DT,fMUbDLa8);CQ=/PO1&.Mg/1DN^&S-
MR6S^VNDR>QVQJgb.Z1ZUXJ;WOE-O/4VRW+cCfQHgdQ-Q0a>aJNBO5QHCJGSUA-M
40=IL#)_QHQC\Xcc9Ag4g@HD1N2D7_V[:&[LQ[81PZf@db&S[U^/WgCL:Ye^Y+PN
<D]Q7G=.FPQ0Hc\Af91L]X+[&ca]=C?4.N1>g2S9c#NTQVCf2WR7]SCP<&9NE\+N
H//T3d&JJ=EG)27)9<0VKLAYf-?#P)>A&9TLdJ.9IE/(P#.T4MEJ-M6+N):\CZE_
20IfA)KdVV6e8)9NG5DbBJ96<b,L\:G(HG=d>Pc-K#YI<2g(_T1LB,3e=Z4@\9+a
JX4]F.eb3g9ECWK>;(_<;N&8:SWXgYQ,<g-:?<:<Y&G@;&T(4;eBAcGZ6:aPfMX@
NGWKR:(+6:a&C738Dg1W)5CFAKf\:aSAX9YJHB4Q)Y\TR(\NYg.g;]C5S3N0V&cY
BAN)L1?#FF?BQ5IK5A,V6B=9/+<BYFd2Z/;TcX,b0U35Ec22^[V.1dM=(WRHL41c
9PAS4gWTDTT@X_8U\gD@2:W4R1^aNNUO7=C>K8ggFg3>[W?gdVaFd78ACRGDZ_V+
=d@/fQKT#)b5LXLQW_(\0Af59A^H+7A81S^.:XE-V(E;cM2^6g7H0JYPVac/a#WR
+3?OC);,4_#LfKKP^L67A><O8\O<NW>^T8(b]ACFHQ]75@bHTMW>afL&.S&\N_HZ
(E+_#BEGa#V5EDZ]?C\bF4d^K4bNP/)be_8#1+VM7O>>a&<A?=@PCZZ<)aD#9Uf;
2]-TM.@3I/-8(/+eA8DS.P^XDDgO0eC+ETJg=D/X#144-F<#]:0GDHdFOgBH0,+@
SQ\O54VSV0OV13(S)&Q5bdX=JDA97/UUAB6M7)+-)W#OH<#08,YgIgMX9>6P4TV=
7WCUBAO<T[F-LYeZ.J[Mg>=?M482&RDV)_Id#L(PM3NVGSSaQUKYb_8g)ROW/C/E
(>.LfY6,XBJD)VHZ?Q:ZA4Yg;0P9)&BW:=QJCUC;OB#)c5@0ae[YD0Ee=L#9]8V@
H)#_4TD,OG<GaLD6/;,/[[TdJ=]EZHOKT7,.;SD9^:Ve,Q6X5g>VMMaPO:CEXAXQ
4f>eVOC\bb:66ePKVE+B7XC7[<7;@O+6K\T:Y0bT\\@-e_b5HWZ<4N?XQ?g2U/?,
aL_eQHTP6D?=(OF/1-&K\aK(AM\PY9.[95+SWMAVF9BF9JFTNKS2e4]IS^.;2Ab7
a--ALQ^1c=X.T55F>S#(/=PdD+]-R-e87X7\92d@B]\^H&YOb1WTADG(<_S39JJ[
+QAM0<IJM/Cd&O6S@<_G28AB9c5V(5XF&&HB<8E:2,:b8gH^_&+8Qc=adLCaV,G1
+(eZ4J,24LZbZ]0SG-RTF#=G\1b,9L,dAK=QS,X,c2>TB-&;X\VD:f9-K^P&E#<T
E+(>[<I6?J^HNXU.K_2BB=(I>a#>9bBR9f=63gC6Y</,=C6gaUR^d_J)3.LN9I(T
::-f3HfYQTdFN_G&AMQ951D8\&=\2]B?ff>N(4[d1fXP[defdJ@C@U/9H2/fDGU2
3MFc)X<b#a-SE^MC6Y=fC\b]bTJMYWB0.2Xg&fM[]@H7(,54Z.G=2S0>c;[Z:U5;
49B,OQRE76WG1#PF>Ydf,490/YgZdD?d,T=g#>IIJ+@986]@7T&_5FA#@Z2XWN&^
[K(X6/@==.;eU8S/F<_P2=>U,Ifg\JcX9&[&JZE9F?M.gE=R:Q=<WaYV>937PN7&
gHI510),NY#6#a.(_D@TURaSdH+WI@e,OE+(:X8Kc98+CBI]9gQB+R(\BI)WG^ZV
>B+&fF-d=?8G>#D_;OKJbUPZM>fXUeb-(,]AVg?((#\438aAKTO&O6)\A;)6L_K^
_<-Pc4GccW<3AFaf1X+Kf)_W1)&YSP?]ZZM4TRDd5NRZf)0\#BB0VPUEO/Xe2>bH
PdHHDGU#)c&O<VUTJ.#28;YZS-,BBT0J:TN/KG9X/TT9LQJSVALW:ENa5:U\:19^
W=[1\2]&@@>;Va(HbLI<OIDd83G#54KH..,Za_MLOgQ;SUYTAOc(?[RMd[IY+=E6
EbCYQ62PW<;7-;7H=)Q8=LLJ#3GO#2;:(>\g-\Nb8XP:V42,DD,W;FN&+>C3AK5F
#YLS77\gWH#(ZWL):e-\(cUE7L&5/,:^5PFYR8Ne9.O_]3:ST</_d12MVWGa>;Q=
56>JN3?[\U/cMLE_dOR;?DHZaEZd7-VH2?9P+55=.W@=+Z=C;+Z:/58NfAG\BAGg
5_J?:<@Q]#>Hb)?@gKbScGT1_cK^L\#C980#\OWQKXH6#TP-:8.P:dX?Rc-)=PBS
H<&f0WSTO9FU28E\_KY@D/3J?MdT.Y?73]Kf3^-;UZQg?+<.T&Nd?L97(>QEI.d5
gS=b/DJ:+DX7FU+CU4MU,2\.RKY.HHA?LPZ?B3cE95Cb-eW08S=\U:Z9WUOHHF@9
f3NAZ?a0/)BWXVeA)5K#[-cMIHAZeTBdccd#O/I&cU9-&4EaJKI5,Aa9UDU<P0DO
72>+6/2[&@R(7JOM=[?8,EAHY>H7ee20V?5@WEINB/O9\=DL.2E4#5N]4-N90S:=
9dVJ8NaI);c]g:X6N?E-:[;G#,ZB\@^gWTT;I5/_c,\egCfUagRG:I/YO_U[c>TO
&0C:cWa_#-fZ?7+T<WGf[=W+7Z&b@SJcDC&g2W0a,=^NR9R0.eJ=3.:NFN+WIO3)Q$
`endprotected


`endif
