
`ifndef GUARD_SVT_AHB_SLAVE_MONITOR_DEF_TOGGLE_COV_CALLBACK_SV
`define GUARD_SVT_AHB_SLAVE_MONITOR_DEF_TOGGLE_COV_CALLBACK_SV

`include "svt_ahb_defines.svi"
`include `SVT_SOURCE_MAP_SUITE_SRC_SVI(amba_svt,R-2020.12,svt_ahb_common_monitor_def_cov_util)
 
/** Toggle coverage is a signal level coverage. Toggle coverage provides
 * baseline information that a system is connected properly, and that higher
 * level coverage or compliance failures are not simply the result of
 * connectivity issues. Toggle coverage answers the question: Did a bit change
 * from a value of 0 to 1 and back from 1 to 0? This type of coverage does not
 * indicate that every value of a multi-bit vector was seen but measures that
 * all the individual bits of a multi-bit vector did toggle. This Coverage
 * Callback class consists covergroup definition and declaration.
 */
class svt_ahb_slave_monitor_def_toggle_cov_callback#(type MONITOR_MP=virtual svt_ahb_slave_if.svt_ahb_monitor_modport) extends svt_ahb_slave_monitor_def_toggle_cov_data_callbacks#(MONITOR_MP);

  /**
    * CONSTUCTOR: Create a new svt_ahb_slave_monitor_def_toggle_cov_callback instance.
    */
`ifdef SVT_UVM_TECHNOLOGY
  extern function new(svt_ahb_slave_configuration cfg, MONITOR_MP monitor_mp, string name = "svt_ahb_slave_monitor_def_toggle_cov_callback");
`elsif SVT_OVM_TECHNOLOGY
  extern function new(svt_ahb_slave_configuration cfg, MONITOR_MP monitor_mp, string name = "svt_ahb_slave_monitor_def_toggle_cov_callback");
`else
  extern function new(svt_ahb_slave_configuration cfg, MONITOR_MP monitor_mp);
`endif

endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3US7KmI3QKozxfjOziJ93QjmeHGK8TDvM4yG5vUDzvzdkzMRBQnpcb+xTbA7LJxr
Ouw4LWgbgFtAHUzwOihN7NsmaGYPLte+xLdUg6lDKGke9PW+TsmMlRdNVrxI6WjU
64ISKqzUDGv5C5UgKAKT7VAKQ6tVNammdHbCWVjccUHc3uYB5PtpUA==
//pragma protect end_key_block
//pragma protect digest_block
tIGBoOIv02fYF0UPBPXvB/+eJLY=
//pragma protect end_digest_block
//pragma protect data_block
R4hLtRZo9khUwShzy/auC5ZzawRikNsjMcsHhZEprlaK79RYJKoXtJqAw7dEmeSY
8kuiBlz76BZ47mfAJTpM3rygt+tt9Z85RIQAd6PYN5jyhc5bk8+pPDRntBPloqe2
zX7iWjKdj1xWbnmfWLcc6CpuLsU4dbBRtExMSHvdBaTrJnYDa4odoqP1soWDJJch
1OUoP/xlmr4VgncevILHMlL9aPC645vaSf8C1Zz0rWahm+DrZGmhOZHDdrlAeAT1
LzmJmJC/Al9CWONmLBvOuc2lWkwH0NFIVwmbfkNhHQ0Dfynh4VmAoShOKx8/XNMJ
lOVhfJ1ICbmhixLo0ORtBEcW+4hZty5/gFlSAgVrF5f9vavDGIfjMKj6CRCFNQiz
84j5GJMAtY90kz3d4KGx3WpLR3jzTRspm25NXdAN0fAx3k24UEEtSeP0k4Mb7sEC
Q+Zhhi4B/Ddb3r2kNDy/ZspCBgrhvRfDSpIDy23+3MJ+TxNm/RfM22fJyAQ+WjLd
prnl2JgNJPtB04kdlIw3G/8U3c4uLa/rxHM5AYeamntIW3WPPV73DQF6mlw3DE9+
T3yKthNg84Jto06ziNTkLJ6wpEV3G62zHfaqNQKHUp+oqFfoWRnD4vktUMbotAod
Ng/Dh0HbCC4M7ZqZCYW05dystnTXD9Y0faA3CkVEir0NRbQOT4o1QVT0MEgbEphi
HFwE/wjTAROPOPT+hBUCvyadV789NqYrqhWcFbeWZUcDRbt1rZdicedAav6uIx2v
DynJ2DqEAEHdzD1bSeiKg6+pKg6mCcWh71ZsLgEuUgPkbiMnL4uCcC9e7taiwRjI
DEZD6HksNWj9JG5EMMJPOzmOnKi6w+knGxm1IMGCkkuQ9TTx+0VXfoO8FOLvUn9G
+PpM8qet+TVqq2rgN1dLZ0NpEErwQrxssVPxlPI6eKgVL5naf63f4AkjGun6ufp2
1sbuTFWgGhnVbgUGT1gJQOiW0QPGobyR1NlNHZbmC+MBFyJgt4Yzsz7tG93DHDQX
A6crIukrQWtq6/dhye6uzoMT3zRbLfRnSyPEelUAi6kiSyJrWtVQ7YcArqjxLJWW
DcijLPIAgaN3Bgw4n/ZZcmgjKjJOBLtyRnF1/ifytDa1gaxK26E9C2jd24pXqyNt
nM9YI8apFTrd5r1zeYbvvMOTaZ66YcF/lIF7pvmVHHDosAGJnypZNgPsxuenLL9t
ZlptVuhIOlOgVbjOmHCiYS8NGJA6aC57JNOeie51NBCKTYFLDOarYrNXomIKS8g2
6qo5+qBmMNzpVf4FFK7pVFXSfe/CWayKSdAuMP2OfBTXaUc1yDddA0f8Egbeibj1
Aiuq2skq86+P5e/+utAMHrYvBFIQcpperMSOnWJaH1ZzM2txGsaJpWF/aXixwCZl
gSJyOFLAyt8xhz4x8e3BWKRi7HEMI3YjLluZU9BBWqebEj3fQS/ATM1iCwp3diKo
ecq6q2nhvtrcPPs0rtdmlc7NgQtRJgZwRt1lUwahJZ7GEMY5vqYJgnqMCWpYwGWU
Ar/ys6o5ptmXSnmlbsuJMpvnzJduJAtXpybViY80pCGxJIugBP0vcVLUnk4jlo9d
/n6ddoM3g8sRkca/U2WAsSdMk8MwwA3bCgFdNPrTLtpJWUAnc4oD7eundMkT2CnM
qt+RWgXeOq1gddxwYKTgibVgeohO0KPNpqayL/rA4rs8JosAEoOX1alDqiTnj/fK
fgYrBD/VYl9aRvuY9BHQQ0F1LoYfWcuri/6NIRc65uoZe3KznWcmMLM296D7RKXc
BACXPvd8q9qrKPM/U3pCngrfGn4LqVuYXxENPfWysxs9WY5nxjW2J53L14y2HJM8
OXqMyB6QuL8mGWfjdrrGwE+BseQ/wwljaZFRjcf+NxBM8JZYoFs2n7KdHv1y9jHK
cHWNWdXXxwGJ5vBYT0JyQiBHw7KCSa9TU1cAQkn0mOuF+CUb4U23EfCcoookyis0
dyQDUzJ8f2/SiRqFKF+7iQ4xN9tKkXQ8gSDJJuFqsV/eH4M7kdZNxqjOts2VfIrV
LyJmDeyvpw6AL7DA+qHHXHXR/BC8yGSm6Ecse7RL3pWOcPIr+2jnc/JFxuHvmML6
YHSI9KFUdQyBY0iJaBiwKwQv2gEmjX1bF17k7AmKz/MFL4RNhCnW7yZak22OpnvW
dZedhlDRp74iaW7lPnweU5z35WKAdqcUwDQOER7CyxsZK1hMqZbNQPp0qfRZSw8y
sEru/q1A6Pz0mi7RrtlxFcjhpS1ZlMUBo5r23KjQZs4799MoyXVVxmLIclIvGG1K
A+vtghXPAyj5U5geqAldHlCcO3TyuHA7BTtqKj+bHH+nvDx35KDK1QCuesiI2f0u
4iVywezQmlbxoqGhAEyF9w/Lze5Q1XEs3MM07gTpwMT8pXCFMkrcPqLqtvXff/JS
nFvH8MR7quglJriOG/WKRBgy967BOqdGukt3EsI1IQ4/HTHl5fOHM85DUfk9pL8o
NobSB3ZlmxtHanuuKqJ7kSlg5XY4dPoERigPsctfxa2weXLypzP5AzNIABsyuY6L
dgsLSZJBf+glFxZAFahT5zjUTWUr2zqXRAEEeZZg7gHiTRR5Sz/lZqEij1DdCaSS
epoLmlrf7xVCLoe/kmaBCnB+83J6yQoTIRXvTCPODy3sK/DOX7p952Vy2RDZFlEx
NEBLk2FFtUNxNyaIu93hXQzUTBgRYxo6Ryod9OjS8nSD8DsuoZbukskq7+UP0/xX
GAuXcIb6RcjItRKB4jhmpw4ebiTVRJIVSNaqiX8G6KxI9K6dRxj1EGTYHxVsI57i
vPlUt3JPZuWkZ5TMieoXLPCNSm56NspMYGmXdYHtVDgsjBwLo4i9if3SWh2mWAEg
uKKZndqaKqg7fN3l8bKZGA++4JvACqD6akew1GvorFA4Z0Zy1ZX462z/FN8lZfks
rb6Vp6uMIIrsMGm4XEAomUJS6DGYzRPc6Cokii2ar7ra+vdr87raBxy3PhJTmj1e
uJhQiz5kS/wlmU0BtfF9li0CASlFIiWi8lhaRV+L6Ux3SE90flufE959sSM67S+j
025vn88nS8fxKLnYmCz4NScvhFloti3OexWDYTBlwkvjpqhQiU3OfaCP9J2qMKUC
MchUDId7kCaarBV5aaa9TWMC2BbYg5x1kUALdc4UWgEsu9BnsBccqPv67lZKZ77a
szlFTuvuIc9s4wEFL6zbpYTE3iu3mBnEfkqjN8LrIZnYZB9dK/Lf36wJPlTcOtUy
y23NRgw+jan/tgwfTTYWi2Fg7W3hi/gzcsnXpnNEcZdB1vVQJRqSmukYlNkJ/ski
gqe/CkPqEiwqusIQpAPJfuhSbn3NYbW9sMTHdYqTdx4Qg+8+4nTzprSlXugMpAjO
rddxNJ20jK1emNc1nEbXukfktDSlNwsb5LzbJdhJcEt45SXlZAmeZPi799z6Tivs
pyCCBFuk7AhkawF2gEL3spb1DvUtYLo+Phwc2Vn12PvQCAp7rZ65ycZc0VfSymHP
6xiSVd/sWcRadjAvxxvRmywEmdlRqMwhiH/hvAJ7pVLHgu/0kObEfgTm2H6EzseU
JFCHCgcs7k7vaMah8VZB8NISv/5pMUbAcAGQP7mWNnP2zMd58ZK3tjpflrmWyJrh
Yjkq4CX3AjWySPtTq+xlE6nAFZ8/4JSm8UdAdD80ffzuObr4Z4T3jQ182CyTb6rk
cAmgMlRRBVpGMaPKdN9rdDWahEJkgQA03F4y89y3pbk=
//pragma protect end_data_block
//pragma protect digest_block
nxqz2POw7KoBuyuyCjzPN7Phv0k=
//pragma protect end_digest_block
//pragma protect end_protected

`endif
