
`ifndef GUARD_SVT_AHB_MASTER_UVM_SV
`define GUARD_SVT_AHB_MASTER_UVM_SV

typedef class svt_ahb_master_callback;

`ifdef SVT_UVM_TECHNOLOGY
typedef uvm_callbacks#(svt_ahb_master,svt_ahb_master_callback) svt_ahb_master_callback_pool;
`else
typedef svt_callbacks#(svt_ahb_master,svt_ahb_master_callback) svt_ahb_master_callback_pool;
`endif

// =============================================================================
/** This class is UVM Driver that implements an AHB MASTER component. */
class svt_ahb_master extends svt_driver#(svt_ahb_master_transaction);

`ifdef SVT_UVM_TECHNOLOGY
  `uvm_register_cb(svt_ahb_master, svt_ahb_master_callback)
`endif

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  //vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
qTZ8UhMKHRmsWPzNolMxURSfjP6tJfCGjEGQlLX4hY9TE7yLyBKH9G53bbMKOxt0
R54yyIcdpyCZ7Vql0heko41XCBIEzOLho5x8TlPB36ATcmuM+a9ab2gjtka3rrwL
XGz1COzqoq4m6YSIaQdttWKCK/75GERdjTjMuYo/H/DNpKZEOstBNA==
//pragma protect end_key_block
//pragma protect digest_block
cKmkEkIrI88Y+2YSTWRHVdlMcL8=
//pragma protect end_digest_block
//pragma protect data_block
0D3olT0gtOySV4wJIdwDVw8aDZiqGN8GZZqJXtY0Be8rH7AnNYChCKZHL4qYDyNg
fD6ssj68tFYwI90jzTT4hdtwT3VwFWI/Dvh2KKu+xWO3lCCLeug4joI8aXNTFsaV
ttpnmcM3bw7ig7WGJp5Nu+alZ9WeGiMHiFtJEMjl862dPQY21zc1GkxcicmOb257
+jOpFUUDDRUn9Z15Fk4C5VASM5HttXdSh+rnVqA6hunGo1FXOFekNxbyVqBlG23j
v0UVF0gOvTNfxoTAFsfKF29PMwsYdb26vbnJrP3K/G1S73YrjgQwXbIX2Vq8YJpm
38+WzClQQcIkpwkfYYOHCvR3MqowdoJUYNcLUwmvZxOFQ1pAev8bhYqQHtV+1Hqc
YcpCtkJP9KRlfW9xKaXpG8U4xyqK7Pn6iruEuQGrXYlv0hAA68z4xw9A/9Zje61I
OFOJvJvwXTAbNX1uVVcjlA5KxomMp7IOqpgKfNT4IIErwwJjnM7+eCX0JZlN9+Gh
pl/h0tiSpGKeyVc7lSjoQYwS0/O01sySdq6nq7Xss6JThJ0+2jeDDMuBSuRhWoJu
5XF2Of2rNLbhHaIWgBOyZLr6FwoQa/sTlo5spwOfM77rfNHj4WL+AEfY3dML6V/8
eI6rNzSpW+z4zz/tWWd7gN9D50LSkt+QQpbaJWeMGTz4dbASri9YkGPDuBj260B6
Ill80Qmn1/0f2BhqKgpdTtDqihcJ44ln8bGWN+8wAPc6+fVf5VVya7J/xTupRCFo
PqD7eEgBiomGOoWlEYvQw+4trnXwZ7tKO4gz14fAbreGaLikco3okCEHeo+24CTu
yAZnV5XTtRQPVHTLQG39GK7e24EFFjqGwdVzaDwSTdf4hiK1eJoa7C8vwOVhwEhT
nsNn5jJJXSkcqQbIQJpB/0jsBuAEFPL3zqWVeMvTOcqbBTVH8HEeX+NFRCPvIhAa

//pragma protect end_data_block
//pragma protect digest_block
OyynPNS4//m3eE6wJx8BhH3Z8oE=
//pragma protect end_digest_block
//pragma protect end_protected
  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  
  /** @cond PRIVATE */
  /** Common features of MASTER components */
  protected svt_ahb_master_active_common common;

  /** Configuration object copy to be used in set/get operations. */
  protected svt_ahb_master_configuration cfg_snapshot;
  
  /** @endcond */

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /** Configuration object for this transactor. */
  local svt_ahb_master_configuration cfg;

  /** Transaction counter */
  local int xact_count = 0;

  /** Indicates if item_done is invoked. */
  local bit is_item_done = 0;

  /** Indicates if drive_xact is complete. */
  local bit is_drive_xact_complete = 0;
  // ****************************************************************************
  // Field Macros
  // ****************************************************************************
  `svt_xvm_component_utils_begin(svt_ahb_master)
    `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE)
  `svt_xvm_component_utils_end


  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new driver instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, `SVT_XVM(component) parent);

  // ---------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the common class
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual function void build();
`endif

  // ---------------------------------------------------------------------------
`ifdef SVT_UVM_TECHNOLOGY
  /**
   * End of Elaboration Phase
   * Disables automatic item recording if the feature is available
   */
  extern virtual function void end_of_elaboration_phase (uvm_phase phase);
`endif
  
  // ---------------------------------------------------------------------------
  /**
   * Run phase
   * Starts persistent threads like consume_from_seq_item_port()
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif


  
/** @cond PRIVATE */
  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  //----------------------------------------------------------------------------
  /** PRIVATE METHODS */
  // ---------------------------------------------------------------------------
  /** Method which manages seq_item_port */
  extern protected task consume_from_seq_item_port();
  
  /** Method which fetches next transaction from sequencer and preprocess the same. */
  // This method drop the transaction if it crosses the slave address boundary.
  extern virtual task fetch_and_preprocess_xact(output svt_ahb_master_transaction xact, ref bit drop, output bit drop_xact);

  /** Method that is responsible to invoke the master_active_common methods to drive the transaction. */
  extern virtual task drive_transaction(svt_ahb_master_transaction xact, bit invoke_start_transaction);

  /** Method that waits for an event to prefetch next request and then prefetch the next request. */
  extern virtual task wait_to_fetch_next_req(output svt_ahb_master_transaction next_req, ref bit drop_next_req);
  
  // ---------------------------------------------------------------------------
  /** Method to set common */
  extern function void set_common(svt_ahb_master_active_common common);


  //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void post_input_port_get(svt_ahb_master_transaction xact, ref bit drop);

  //----------------------------------------------------------------------------
  /**
   * Callback issued to allow the testbench to collect functional coverage
   * information from a transaction received at the input channel which is connected
   * to the generator.
   *
   * @param xact A reference to the transaction descriptor object of interest.
   */
  extern virtual protected function void input_port_cov(svt_ahb_master_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>post_input_port_get</i> callback using the
   * callback macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task post_input_port_get_cb_exec(svt_ahb_master_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /**
   * Callback issued to allow the testbench to collect functional coverage
   * information from a transaction received at the input channel which is connected
   * to the generator.
   * 
   * This method issues the <i>input_port_cov</i> callback using the
   * `uvm_do_callbacks macro. Overriding implementations in extended classes must
   * ensure that the callbacks get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task input_port_cov_cb_exec(svt_ahb_master_transaction xact);

/** @endcond */

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
HrOmr9ER6g7ne0wI5GjHBzdp+lfEBRTG0RttAkjZw8c0LrjQ24GNDgGRmwfgGqqH
73dhBOqGn8SF5UlzlgWE4RKGBrCsS8uE2mSJQ4eheWxgK3MH5CAXl1SkgvAd7pM4
TZe1qvGyrlY8RLXSgsJcVrQ7my1MBgLG09PeT6wJyCq9I14NTpP9Dw==
//pragma protect end_key_block
//pragma protect digest_block
uRfUkHTqyFLZVvxNoJqYSmRtYSk=
//pragma protect end_digest_block
//pragma protect data_block
XOjvdeUyGQNaOZRR6bboglVnpQ4MMFo5ypsB9Gd2JiSoLXL2u0V+NIPnavooMIcl
6txGdzQ1TN5z5F8lZubZmBfDwRk8Cu2n5KYKm0iuiwSkHNGN6AQkutv0UQW4RDxB
jNbXZ2gD5KRph20CU5NK5ZjWFa5j5pzzK97IMLfycq5i4gM3quDTZMFfn7adjtZb
0tQsIsNnjQFQgwzygh9WiGXJB+er3lP+5QtbKhvanLdBvxs2/mSt8FWFXFx8ivAA
igdP+Es9BpQ8fVVF38n4KCRRj0rVq2Jcw89RKnBWCD3x5RVItqGiq8E/TYUVDW4o
hP+NpHhowLJWyTSbyLoU1kNVuiimLRyr305IJFQUPBOQcNvkRp80MrTS8s+TWKcS
LWnMQqQK0oPPvjpv+rMqLfN9yFGa4rMBBg5xinFsorxKGWbe9xVxUyPpOlA2HMwf
wIkXLS9ps2e+EeZlymsk6XPwOJma3zxQC0B/RqnTOxIG43+jroZRSXqfiQtm6Yof
NrolZ91cnzxon0xLW1Op7L8wbLgODBcmuXYc7wt+JqE=
//pragma protect end_data_block
//pragma protect digest_block
/pJInKc6HkB/u6m3C6cPSsrZArA=
//pragma protect end_digest_block
//pragma protect end_protected

endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Bd6NzW5018xupbJ/1ekvgYrCss/1SjSWlqFtsMdq0WzN1iJPcWYuJJDkUSwZLtZi
Hr9oVN12MXD8+13jSKIeQM3c9J5pMB2q3150Fi7gE09TYptEmEK7JNrCnmxDzBIy
TWOz/S0LORVwEA8nIOGQlLQDdos0xm7UDwxewXLt6fBrxKyDSv1U9A==
//pragma protect end_key_block
//pragma protect digest_block
nBsyoHHPNjZxYpr0Az2SywIHayQ=
//pragma protect end_digest_block
//pragma protect data_block
5Ul8k39c1/33di77VC23dhEzWfV2ij/nB/rLiArOIx37LEBci7Kmy5B5yKNg76tm
20rmEdGAG6VzAgdM1Lb3uEbtzyas+GYy5TiU1XUq/dsLZX/iek1bMdQu4EQkvrkR
yR1mhJYhItOYVYyDsKPrqpSC0DvlzbSwADt4xjYygFgYo43kcaN+6w5t5M3ZzT3p
d5sAyeDCitLJI9RYFtg0NlcCZ20xY8z0s6cKQLer1ENMsVAyb+ObZ9oc4qv5nBsc
FBQICbGnvQLhP0VMgNkH7BPJ4VFp2rLJnoNwDMOdtxOpqAqhPQ0yCr37C1COgvTD
vhbqjwdzygjvkSDYUV46g4UuLJn15VT1wG6zVYeoOSqNnWevwUrAW8l0w33ui9jc
1XIoQ0OserG09jBZNw7SnNBWPEnegktI7wy4LP1SdyRw+XWTKFoUpCKe5L1atARo
2/N+m3eBCb9ktHyiID8Mov/UlX55eQXXl7FPWeM7TD0ICrD15z+Tip1vHtjrW76g
vMg9QB8ATUe+gj+cS4nCJlnjCfye7hZ1jobXDrI1UCWVWBCaGfckySiq4C5udrDW
cR+PA3UGzjYWhzk3/geSFzyNHVf8C76vhXjfsB7GErOeexVelDkjFSXFVk01ybxa
UOmh1au9SakQkosjInLJBOfa3E0BDlan0Tz2fn25SrrLnYuvCNsAEe9NNubniEzZ
vFHUL7JZP+sdwYcTGTbslRV3mGQcn+QjlmexTm8APDmr/o+jdmewS2UAHYMdJos6
Ql03m7EK0HlZILxoJ5rk/OsMksPTANvVnL2I1Ds/o3CmSiKvh5+P/nm2/BGXx0ex
Sz8ovjGRCyTVR5BEz2lgUg==
//pragma protect end_data_block
//pragma protect digest_block
L4oI8wwee3/DOoJb20gjAZ24+WM=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
REECuRvO302o9o3SmngrfajbIgS/8graJ8SJEvQ7tF+YGHrrZDm6uzqckhdoFjL4
Yw9j5Z6EDkPaEy3eDaKRbZXAzT46kbUWwJmmqB2Nnsa2WFqhz0excxCMw31xsjZt
AlRCahYN+3GmnPN/dGJ0bqIiUE1E5WryQ33S+Kzqzy+syDLBT4uBCQ==
//pragma protect end_key_block
//pragma protect digest_block
IDhnhCOvHG8cQBZmJa1F/lI+2Hk=
//pragma protect end_digest_block
//pragma protect data_block
PoNAly/fjgB+5Tablf03aB2P9rfDe8yEu/fAxKsB44P0d4SZKffcI/6R83oMDWJr
A4bnK2ONO14qFrvMC3LEOaWf3W7d7R0DN5CsHbq2Fv2XMyDOXJGAh/I/WdupkMMD
k0zKOkMVfCfgKSIbYcEqa4OTcwuIDrR/vtV0zFAUMW/JE1bUzQ5a/W/t5wOX0C17
4N4IxSomMd3onQHD+S8qJ6qcI2dgcJ7IEaRELF7WIqiK1YNkrhqNiYTQHhygCte5
DIGZYk1j922MpbFGsAGxV+G7rKA9pu4522H+pCDcEQkGSNhESwyazN56vkyaRKjt
axmrngipkvSVrxkbpLFEY0nDdxv7dSOQyHWRMYxMyp5OP2pn8fOnFc7BK3HhZ0mz
8FNwaO/+9kHZtcXXiLLLyy1UkD+DD3mS7s436wD6WWxNlu00fzpvxjNQB/U9lHBh
gv30F1cRU63RTXZIj5HfXQyIaeIZksEMNJch/LaSOANpSR/HUdtLmjt3froM1p/o
bIvWlldFUfy68QioojaNFGJtMn19EyVlcJOKyuqC1UUeliO1SPNYUPJKYLHYLMbm
rkc2aO/WejWynD8WLC1oAcMhGVqNygspASv8KJyISTI+V4GER798hhHOKQ260sRw
Pr3Pd6eAW09hIsp1xuDStMiNVp/pl/lKdD6JsqHzl2ux5oqj0PmEnoA63+cYL51/
Os23ucogENS4w4Omy8PzVAAa77bGwfIJypnHj9t/8t49Ecdb4aiTjr0HYs9vwrVr
XDIbDE08W2R10sYBThaxlcQNj6FdYwa89LLZe9sGJMmqoQLn8RFMq2ZOsDi1csZg
uJuJvbxkNooZouEyleTbprYM6GcVFm4OE7OTYG3pUHPrgyFEun/utpRPZieiVjQ1
W7Dct5AuyA20OJs3firujkrK6N/9DcPGbPCXhoz0xnuy9u3T8l7aWH40J7UOZ1Yq
mVfkpFN4xom5AQLTjuYnJIaIPQ0uaRvabvVKnuSymdNVUU4F63njEq7fKVvyJL3Q
LyVpQ0yYM1DVUS+vinJ5jSAtBUTWBnuysL3qQve0QUmi3R9OZNMdnA3WBWswOxi2
cURk8Pvipo6hXCu1Yjm1mswVIwf9T4mzkC9kVysR98rjK4nHHuvHB555dkrcVI6U
UQuMmcpigLCDcVLchpINM0qNTpB4dMhq6jGdI1pNIplRZEoNR2H+scuaOX5YGQqY
zPEuavQ3KXmSZqeB/JsfOMxvuOM66Uv2wOPR5cFovtH+Us/auMx02G4/rAbGLZQs
01dekxja9Os9/mXLsvVYFFx/k2G2Urfnd2Y/cvwuzQLjSTBUvdfYyUYjn/bd19im
FFxXXoI3MVVhqv4Ea6+8YGCK0OFpMrcwuk1Y9i3zNw7Rh6sbsWzNYpwdKwJZgKzO
Z2oa7FpUiU7wpQ7i5QfP3dn5E9F+N6TjSUmbtSHiVVcR1onJO261U8H3jO4euXcp
WkQXCKJiEzj575jaNE4SaZBWHAa/v344eKt03diz8k+POarKjgn6ETjweXTFrVam
9Q1ifsApSftJjDWY4/t+yB6YMPlUq5FroU69imgnfLTl4MTxw+iek0qQIzNojS9c
ZfSsdnb36UbwukzvWOGfo2kt9ZZxCxSjwJIrK1XxNlk/JGKbGaQ2KlrcCTXhd4I+
EaaSaRnn0E9Ky8vKEAlW9pvFWHF/xYvNMJddvhDLE0LPAgVyshVjB8ZXcKyjwiW5
D7FFDEMXfOs/jzrcUtxO8FOhLxHLVrusbvbss+Fz/SUnr1g1mtEpfO5vYsbNfQdr
n8YcuppQ3qq8Xpu/tyCDfMjP7YvCTULXaeTRCswuPI2lmeuyqwEhDGWqAFOnkha4
f16N41+EvApOmHNsv07R3z+rpCaTkBj5GOVuDjvyBwTmD3PnqfpWmpAZpK6tQlxV
W0mlXG0unl5/NThz7p1QAhPAtHQzULvR6GnmxCNLheV78fIVXoD5kbBZ/qGnok0R
4ovg1GBmT6bJZL+ajcsdL3zDFlKzUXXplX0x+oMhn8ExU9dYiGkRF7uIe7nPj4u6
ezViu36wdQBu4E6Q+6tB01oqrPC+Gyh43k3Bu3QVjPPn5xXryxpzh0PRveuL8nTa
geD8RCqvAgoR110Mp64w99WwFnpG9JDqDSSzhYp0NPa6zm9KbCbrQ1B4XFcpro2b
t9XAJCVwzFLv7hS6j8xBAWVefWc9MS5yKrFedXI7rDR4W7x5nx9rWnr10yNHx/uB
AyBdw9zeqDUz1kk90eGNoSYZ7LZIMNEyE3QgxL6YGkjWZ8kfrdN/ncZSMqJb6XVD
3MsPDov9MlZC7bCzjslsI94RaC9/qpNB7EkW/l8ikHmAOxTr4agvNCxlaDFZDaa1
NvTYl6lpswLroMVhXFCmLAox3ospc5bNsLZVESiD9Or7Xi97EmGm1jBFG+qx+bUj
RyVQ2pri1pwFGme+TuNx9nTa0xFoSKVbK4nKjDVFYYg5PS0Wb4aJz4RwkmcENe61
GdfcC7dEZby5i7X1Jp0wXTMUMcst9gFmAEi8d9ZNzp5tn7y69mHBKrpjZMTZatGb
gOSDm07LPM7p7ffRLocdQUpnY7aZxj1o/bOMhb3j+g2dVRBCFPAnrFetwbHHcsZQ
r/cSwJq8SiO0vvHXbdJfaVRrTqpRce716YA2PEQn8uz8nFJY6+NkGltDQ5QAZMCR
v1JGLc5xfw6lDGIoFRSUXB5ASEthywGxSmDSdcK2vQxCcEVqleW8D8CTU3aVW5Rr
Lo4C28Uf70b+D5EHXh04GhufufzyjqRvJ9ESUzTkTbBZQ2BE2Y012ui21WbRQiuE
GtZXh3RKlbmWMpzR/hhLsLrrWi63sDMMY+DlHh1htnDOjoxaVDIWxTUjszaL1qjX
oah74mPidqPS0fq+RS4BABGLBwHEt3H2TCtoorrCUIf7nmgXE0IXDUoLVvQS/n7P
Z1u/SDx6M8yd/ekXbeCCdAxVw3XKWL+j8XLzPUPnsDN/CJtHh6WutOQm2pK2FE8w
kcF8uCzXBuh/RHay9ZQvgxJmSgCYVLtzE3SSU23quh4EHqGwp+tRxp6KYQeWD1LC
ZNQ9/5C4k/S6nyL0xMHyqxbg5al/br1Dkv9GOVNdQFuH+csptTMd9FMBmQZvioz+
DKw3hBrAr2V2Ou1iD/TcCVfsdcUqnV1W1SRv6CO5vHRtiXjJiskUgtcQO57Fb2MP
Tjkt4CuRDyAWHrJ1SdgfXRpazLZBe8zcDmQAIUmWov9zhMtqcBsmO6FOds9QTZ7+
POC/fSO1TB5NvJuIj2n3XtK1JpffctbQNJqXP+u5cgWTZLr+niw6ODix1Ymxm4yx
8dXq+hkx6bvnry3ujriLnN4DgqduO8WvszkAdMx8ZlefgwrQa1FsZ1yG40iI8ja9
/lJMjlRNaRz9ujV9PjhpCLvBeTy5wvS3mjz6vpzg+LD12qxuj28kFhx3PZSilvZw
QjpnQnSbCAbXYCWYsvmTYVCJLog5kzW9Q4rzr/4GkIxze5n/Pon8peOsD3b865jt
JxowxL5m/kE+MW+QxKKy9BR8cwSNvOlAM1yWwuAP2/rU+U6OIjbis8hS3o+mHA+7
kBR7WX2C23s6mOmFnlB1EvfKrbMtoIDE1FoLIzEr86rzzSYltP/riwDpMiefBGYY
vGcifO9qgetawZzDBvSjWWyIytXuNTmROY/DlC3hW/LEVh6pmIMKkdhp16urdyJC
Y23OK+u2/kbVloJU1xEZaRu9sYZIf5pqYdoUZjCRrGMM0JO2mzWePvifih4kFOSD
ivyDVsabCqWOsOY5z7N+3K4zgWZzAOUNfs1BcBrRCdQRls6WWFY3HdlmM1hcQn3B
3jabToHRaTAELcqPSbrPJWzLJlhVXrwQowNpaQ093KCj+szFLaj14bV4XCWOfXtq
J9iGXt/6HaiLDr/2PIT2YbUtE1bt6fNhgGbfVZbYeJuTXuSEidb/Ec7eIwBi7HB3
9XDAPQqCRm3bafttWpVyKMPUR2I6BbY9M2nNtZuLMD0AgvOVpmbRlvShR93lcK0p
d6wJyvcZAru5O19f2Qgq54fixV8LIRYVULg6TeJNBLiWd88pejEWBpTRrCRfSYIe
oLjhpDEgSkfeJpA3CzYN8wpsCeKEPVz/bejGbJzw/qEebe+k1noq2eLrUA8knigC
C2++Y3zZ1mC2ge/RJ2Uuh8P+GCSpdRB3Q7UdRlhGNO8ATVOEFtKw/jKfkwZXGTKE
vDqJggQNxZOANyg8pqS4JXuYWdCWkIPTDN1diy5Olk++WCWVmZzqqL8HK2tIL0rf
G1hrVAoARSCSetSuEFPugsQku8n8G3VWKJi1fXaIvN6L8SGQLfyrxWVA/ZSRi99T
1B1p+4noZ1KaxolzCy7M1becMWRMx26i/naLVvkxC60X3JoHilBM6PJatFmAvXAI
T0NloBddojPz8AIzycVNibeOV4oXhqR2jJtdEay5ihkIryEugPe/wzTzw7GkpRX+
VUCTxDgzL6fISAdyJ1KIYQPfR+8SfjBmqJYuCVYXAR1G5z83MU7miZfraM0KuW8D
KwrbfQyJdUEuFhF33pT5lL/7JXiCOmUDKkAkq4k1HtjAcHD5ceNT5xBstWDQh/xc
SGUeFLBVi1KCWgxDxilKTcDFXPtQPT8gDZJFAeRrwDsCm1o6q2KSPqmpaFTgUFFG
f7cZKwyeq1yUUNSXAnfhFUGOi48j00FCO/mc2LJm58n+sNaAVUMkMK7W0ASvqqoD
H+zFr3oB1+Fx4Eh/n6oUQl32r3BJoc30YPEnBVbH67FvxQ6Xycj01Q93wFhMOv6t
qU41iOkplP8Lcfz8UB9FWarsAY7rgAFiJUFiaDF+UfhKTfcsLpDIPEe4G21x5rOX
3hhxNX/tp9ilg+pAzh9GPU6lDN5tzhHu6NFhBD57HQ1Qp6stcDHGrX3CNunkjT3p
qLeihylWmsWWAunjIXYlLivDH19bVg/VZFuqyV9KICrUa1261G4/xG7VjdN80uhh
BDlOetJHX7/nq1pXBlauL9P52aS17XAXa5m0zrllnsbr+W4KKt+cGlR9nzIZawNJ
9QmBkpddVRK5WeNByCQ/UaWS7EoPeq3FGMHTrXHLKieUYpA/kAO4sWbBYU1PW1gJ
tZQKo17dlE5VI9nZGIebkzUlO9/sAb89X72mwtnOqyQtIfIV9L8ds2NOiTYvz9S3
qJOp3jSy9FhiqFuOvLOa+fEVleCBSlC60bhuVwkJEqvaUqvGOBLraCprDBpwcrXt
Sd6s2VSTlIOk2fUr7A+tEduOm+QPVf9Hv12zZIvqMyOdJ8z5xwK8b+V+VrznJKo2
Ges8pOg1NC5GKkvW/PP8o1ZsKNRNIVjD7X4qr8ssxWHYUjXy1W3CeiV9/WgaO+8z
csqnWt3VTTTlh3ApF45VUVOgGtJvhbdoP8qvG6QtguHvfL7DTJjM0EYqRjDuePl7
5w3iU9aZHy7MA8SeBeqcdY72rdgqLPsOE+m8hz6oQnQGbugj6tEb/AmFYD2Hdd0d
r21K88qNrYd8OJNpekHtP1Em9ZaYh87d9OdpGop7ip3lK88TsLnPvtww+Mq9oRrP
lIw+fhbnYL8rT/WKrZb9OyBPPlMTOEmX0vuu33//YSjhh5WfzHZDujJHJLGhG3Az
SyLAQmDZuK7so3IKeQwbKPm83K1DyMItAb0I9SW+rFmABBFNTp1I6RQsSCN3MFtj
jBudRAS++Z9MoHrZp+Bc3v9EehfUjx7rqi+9gL4RIp5Zlkj3jEll3wzjgd7x4SLk
W517QYk81BToP7fKghFspxbTo2QJJgRntqGdyHAZLo+8c5Sb11hVyuHrOzQWcE+g
Moj5FBulQZb5Yrf7bRKziR/iMh1ResGAElSV/wS6DqLDqw45gJP9A79uM4559B4g
ym/LWKmfxRcYWQQPWddQgwDzApL3eWy90FJcSRzQcWzXMmQZeydd5KGg4091UgyH
Zr8bhYLz4uH19C7r95T3lfNO7S6+pbZuQwRciLcFUIQlQ3zvuIBFndUxpP9VrIo9
TrW450hD3+RlSxEte3KLnvmvm5JosUX6vD0wAJwytcn9fSVEfo7/O/K8scty4NLu
Q+K/o/mhi+ypAotbQr+D6wFcw7pAbx61sw8fjM5wPW3x5Jrzes625uQecV/2dEiy
rNsCnXYvNv516gA7V2j2givqVodYBlNZx9KBSnBNmDkC3cG2TopGcw5t3ZlizyhY
EojaQcZOQ9Q8K0AcTJBWER+xiPyn6GV/bLtqF+7KhIVVC4OJT08jCDKdqdB2nChc
h0542d7TXahXRWdEwLjC1JX+ggBJIMPCN9Y2o4GYgDX+EwFC6w3IpxaK0JKjTi0E
7lnQ/Ydr037KOGK1XjZIRm+Takrf1p1jw8XzGms/JJhdbX2DyeIKsMbmu/4N2ih8
iqpW98UABZ8e1lDPB+RoGIE2FklRVuimDjzl1DV1VlaLh1Wt1I7kQkfe+Mvkj/9f
WnHcqnZXLtVjPYbywAFcPsjx+dj68QPGIHjHzs5nxlBntA1ihfiMWEkRaVuvmuLJ
SYSuHOGyEWO9hd/dfp7+x0i4nIZL90qCU+Q7xwTSKYFnKxPL+dL7PoFEToZd66lh
cA1CeKx84NJRT9DY1p7P5FqismsRXwCTS0CGbKl2J9i+pmNYhHXrq/wJd70w6WOp
0e5o9ufUZV/4X7QnG9lA3/HNcljLIwzoJMAiL9xhvlefseLJNfDbFGJS4+ucn7mx
kDsQmbacAY5Db3Vm1a04YEhmDqjyBvKT68o2icufUbLWzN+cxqH6HNstpGUd4mpZ
55mFoEZWWxkPph7ryPnUkRm+mgkp9nYxYovxVD6NevV0aSwcbC2tiCR2ut1V4DlI
Um3FcHScUtSkAWaiAnKueCNQtL9/Ds/v06GE35T28Ex+GYH9Wu0GoZ3+7qRl0+rp
2caM6TJL5RtZswyYvT4zK0svLxFBTIuBAC09xaqExz/WKlbdDb2ql6bXs3q1v9Tg
uBelskyFTjGTnTvaI8Pe0tGJ94TLj5+9kUlcqEgvHk7u/Ue27ehzTGouzgMDk3fP
kSpo8h2Mes98Q4CqmUeCDRL/rM+vhLuVkVX5j3RYPZNILQdMWdvRSAqaoiIiQhAS
7cuLl1iuBJG8KKwh9Cj+o2OXXLzPE/l6VC0oSOumtxzmqrEf3b6J7XnhwnLE9WDM
hYQqCg1cIfuy2nwkAmwMv/Vdn071K1YuF2pmWpw1TuyBNOK1rcPviySvUi1xORNm
fm4sFDc1EJzNZjZLPT+0iCybRF1yjw8tWdmNvz7WM5rgbPPB+I038NceNKou9MV0
PDhl6o9shzx7uR5yqZpRs7ybtWMh0AeelRfJrPJHW/iQ0xCOzLaCJ9w8EMJ8orzC
EBur3ZDa2H3+Jqeul3WJ/w+6vLeGMvBW2G9GZWi25xxCwIQ84fW+eZVxz0ID+qwo
GaZFFzWg+nVavz586D9TDZqAbyWnPXJ+AHgIsTLk0aFJD3+OEMFbH2qh4eHwZJxH
444k85MX5chJA4P/lhKMGJuC5yibUKjZZaXZKaVBnGsAFx+c2oO941Sm+nFV7zQm
6gk0ZhicoGJ5UiQbYgCiIoymrfkUxcuGIbeAFDeuGRmS5RDJ0jwQbA5o+WtJWfsM
uIpWb/+gY/wp9AqF6Q7JzWyClF4qucwiDn1KR38X0Qi7FmftDosnkQLyrdY1ODCK
wc8OHZ9oSo/0BnZO4WzPjdWCi4e2QgvYk/KcNzReHNCqHw88N2mDAjp2lfCZC+++
1aOr+0BsrHKk8ynb2A/AHJ3eLPgnaJFDwuWlK78Uatm5x7bUVkKKzJkEH5VEVscX
FfVYh12K26Ryfog+/9SBwS3dXGe9XGTJegClpVGPydtmPap2+KB69DNFbbAr+yza
SDOXZaU6+hdi78/g7qJaMTBpqinBYOqoLoOz0mmMze5Prc8Rt30iyzvC+yVjajTA
DlIjt78/kP63Rsa79/Rr51BBfwWiG6dci6RiYWoj++2z9tkfuWLFlwfJXZqAlUSW
cRvSSfu7ZzabnB/7uIh53z8nZN3OAt4Q/tOLGiXJJY/ifEIQYH0+bl9NLI67h5pp
o7itF1FzNzjlP+7mfMDmwnHQA0Ws5ObKT8WJ+KwoMszGJ23Pe5GZSU45zZ16rlA8
4JfGLlmnC4wOVMxrhC1m96WlBgsapap03lOrtc1AMDMJLBSpTH3F6X5+I1LlNeGi
JFpuCYKNW03e2lISVkKeHwpp2FahZsY6EWfEuAqcF5BZVOQihbddTdicTGEyKzJd
0bzzoOaDw/cbpp43CNnFUytuv6UaUxktVr38rfxq2y6DcGgHtoS3np8gBhZ6R8X6
qBnHrLeHDoVeqHnrZgAuVjJFbd76LQeAoDBcgTVLKL49z/xIz8ONHKwqYYZcvrM1
DetlBmvE5OZAC212hKwSXcTnCX+Oxe+TQJPrquiCt5BVgYMZ9oimZm8H/1SnXPvf
LWy11VLjhXd5Dr48f1vFiIEK7Vb+sXExkQs88UNbGY2bd3VeH3IveF6GprzQjrN7
3td1sdwJPshKIsMVyT6B506Ld3Vtn/77VXWcdPeefu6rue1EaYVvlSvudrp2cpMA
uk6nuCwWKZMDezE4Aiyr9NsbYUUQy5u6fe7KNRlUWyRzx1V3RPIRm8JTHX6Ut5/y
24JqPoz8AXkOEPMOktKAd4ZApzQ0k38ZrEqnWegmH1gJIpA/nJSJYcMwKNJuwsKY
oYzUqIJNcTXWJuUoDDcTv+kaet3qvT9xF5vU/lFGHhrFCc1ZCxZ4mhS2a3nyS2nA
v9TUXoKPnwTgvhzsELa9q34sMfSq39dyFhWMfonVHcYxyF43zoVg+nNGJYEXEuq4
UJQ/rUx0kOYgywFQsKKyyWgzM7Dwz4aKiHaf8rvWAAd2EpO0OES/aDxWOnahPsiG
77yfvUklpxaKoq0X9jxlrZ14GdxI1ZdeqQcOCdLlRssD5E6fHgyyRxosdLtMqaQF
KsbbFQ0DNkyFj2ZBlQM+yB0ACFGIjzK3BtqTIvAWiX8RqsF2LauV3tPpnlEhMpNJ
NJabaDjWgcmTpRfs7yOZBvwiHeAD+/VHYsKe2DEiFtomJlKPD4vijK95aqMgMm21
DR4yL8lo37/H5sikZ1cR+Q167MzmGheX6hKKe6d67j1M0vhoO4turuxVRzlHPfAz
hZtVInEhbY8m8MXm+i9GsdKcrepLH9WarOUeaEDCWfjrkHz9Kds9Q52qN1dWGk+o
DjtiTeiD9fy+zlf6AKhSaWeagbnZJ2XQ1/qvyBs2sXQVCO+kcYSiLm/FJPxBuwgM
jZC+H+j1XzrHPWcZFVwkVMdvBkLgl72xe43kzvnTpLmQE5V+tCmnRlWp1tgcUzd5
s7sSUY64exxjazXY2r+GNjHHwUG+WBA8IfZQMiPYp9Abbv6WqeeZny2ZJOWVLp1k
u/4YV8abnum23QIWuMssFpISTGCaYOL1IdfuKiari/SePRsviSox7CdGRj/gAWG2
gIhz36ijUGUvooBn7ia7p6mH4YLZCN/8uO511xxJXjX/CeSCa5o/ZaXFUz+hvJEJ
eJYf3aEUPqbFzTvxnFqKKpSzGsje0M0LsehXw3i9FAiWiGT+CWZcNyx8wepg0o/d
ATzsnFouKUkPEhiU/bW74RYjI967PI4CqdQQvYrHTTSzH/sjtMW4zv9cMWA4iSPs
Gepp4fUHPei4Sc+yk24x7Zn1v6ABX/rG5SommzF8+uI5vb/HVc/RK9wxNGDqypM8
/i7EkzYM033vdUc8lUDo77Uu0hAtnC51jse5OiJ1E669LTboIOWwUUV2o/7AQ/WH
Jb3TIOqMV1z/y+4Nfs2K/kYQzyTKsYUjqfaFeyXw01BWCVbOMDU01k+IM2qrvNc1
cKDhajaREKY/k7vMvc8Z8ONZnQIiM/63DkSlRUHvcjcBUvh1u72x7HHY/lLeejPS
I2Z/oaxF74L+6awLSiK5zcxcByjpDafDrKFSF7GR5PFo7GPH8odkgwQwN45eBC3o
aVDxf+Qx+uS8kbkvnJqtcK+NERmn5zjkJtZfbH+txgMLpYIcVG+1xjvaKn9O8v+D
PvOr0ruvWBgK4UmAO8Y6ZwY6RKC/blbtJ6pgrsqBPqRMfw4VpYQhderYthTgTJ60
leqWz4k35u1qPepmF9EyvFQ95phkGAq1cpWgKPdWCDZL9yW5dFP6KpU1VxBel3dR
RPhVbXqDDIpBk9c5XrNY89RNPurKgBwJrTWzHCyHFhM9qEIwBEQXzBa9euP6lfc/
4GWZS3+6LsoH4ZHeFtqsr20n6phMifXv2amoEaYqu7qyxQP9y3uXNcNVm01VAeb3
NWBQHBiGbLQAWEeq3i+T3jJ8w6mv9mcf7vAO1+cl14K7CVphh7USE7gMEK7ieQl5
9b7AOahN5+MvzUQDRlYyE1lAZu74kbbDpOwpHc/FyEpSIeLUkTRrufYs4TweUocY
hBndn3vyMmGDJVlZQV4hQ9K0vB73ZWgIEZeIiP2ycBNl9d5+l2yEqh507YyrlYGG
ZXasRpCAoOnlz86SbLdw3qUx9JErwAMqGPQG+Ay1JfZKBGLubSxA9OVPw91qDGa5
m9zYfMkur/nzh6a/fyw/1QVQ4R/6YXqRKrGd9CCYtRjeBkovKQMxRnVy2/Bj+9Dn
qJgNpLDqqudDBk9iKu1Pr9V3salVeBm+6Fc4Gux6U9iKzUiFt9hvMKBDOzKYDcjF
SZ9IcwmgAoIIFBjUUlgQiNgRaDDOLm/MTrFXUWOIrpa9xUfEyClEHhqiGwD3jyfd
QwkVCToA8we/kNOLb2SlhsuOnjJZfWUwQPOopkIwsS4va5Kr+wZJ/eq15hThdx/6
mHriT/jjqN3aXcWL7d7EPBfYr99miE0IkXUn3QrwmrIHFIJLVPOtFIxInyW0g+iS
N/iRcHSf7HMhUp8adlSYdw8zCEI30us9FUumou1K7v87xHPMuVGcGPOc0ocPx31F
7lf2030XMR1DgGUGQ8p7UyDqATDP9Byyqct/y9JmcgA2eT0LmhGxqbkZSqpfSFlA
Qdd1sGrfLSvjrgCv/UpYlkK9rPdo+3URLaamNA44ipPIOwmYZShRMGrG5NEaiyIK
BKWkbktnLVu1cAif1IUP8CVLWq1ZmW87i1qy2pJOh0gt0+j8Y1SZDYm4THHZp3GG
4cLkFnNXVeoHB9ryl+1Ji4O2MfYnZJjWSpyUJ9oeD1WW3y8dSiJCDNeYv8C/8zig
SuvGbiwPrA3nDdkcgsbxZk0+QuwFibsven9RkH6iTMI7IeTe5xSIMJtZcyYnqWRS
yWWfWLxsczyrd1Asp6S/xI0QqO+DkdO/Yk1kiok8Ly8IEoVh1tqEiXPF2mHDWLkn
fYDJhtzLvMVWOZ9v0Y3wf8uDwFJJ8ElJFydWHCogtHVCcSsyh4sPGl5ki8cYBMSu
P5I3KtrZjaxfJ81TE/3VlutvbJfknnN+d4WDABmpRWjtJfyg/jFhNaI/uQl3UoPR
hu7N2X8+cdOV0GY1d+xXFq6CCiGWUYXZvHsYzHWX5rOQqLvN+tXG2d5SJy4AMk8u
vs1MWpU+d5mruAOq5j0eK3OuULOJg1CyvHpCGGcmoNIDLAXELvDHEsVPeunL/MxB
Qp8eHanz25DYG8+swUqszUT8ukmS+xKU97bMC0POqoocLEebFcWhWkHJehmotdGX
+LatPnp6QmozoXrFSzeot+BEnN9ZQfYvTkL6BrCuLWlJiJHenMG3Km3Y557Tkld5
X7HF1ZxCDTSxlskLfNREMqBSBpwJ54m/2yFfTuLDJB1ApFawae3bWhSvNbwJ+96F
ID4TULxfyXeyYKRnwmkE/fOe0lAaoghBaq/er1Lx4ycX1+Lmv64Db0v9mMz0UI0l
25IQ0aW41csHn1CM1kN88bOHo59bYbKFy/zjnUEsJmvNuVS9CW6RvS97rLOclxoW
FjKyddTQf8ogQxeJWVv6NqW5hu5QpeTDLc3dC/yP9mo/wLU81kfVb5pHdShfdPq+
auJQgZAH6iKjiaMVxoXFZpLaluEid5ZxBD9P356zBuJbCs3Fqxx7DWH2mVdVzl51
ryoWpqHSRWN9aH4l5u3nM4tL6OYYRVbLLEqq+wfU83iFMFqZ68a18vZ3FfL3cmPG
pPu5cW+9S7wxAqNi7J3EHYPIqTsnyOG3kIx9EwNxWQOwxZafK1C7PwSKjuKYIC/Z
aE8qIoL3ABc27u74rb9i6HwunOKwacdIM28n+kgFh6sHxjMEFFoduyMpV4q/1aCn
l6FHE8zBLw/rzkHIZY0Hg5LkEVeAMVN1fidZn4JkX5re4RYJZA3gfuB55pbEe/u8
9rCvaQ8q/+wGn1l4iwk8zBnRupIn3RSjOC2Bw0HaJcQipP7N2U7ql7wluSMJ7xMF
9+Ka/yiGTon9f+jwHoytWVTqHwJRIXCHvucSlE1m33TTby9zZgnlIV2X3wLqMApy
wOzRsZtVcnnV2rjxxJq0/04AB8b/mpmFzeBqRAn+nnynyRW35SPkXwm4nZxS/CSa
Sz+jEI2d45YSV3iLNMm/cI/okQqDAaHm49qIR8oP3O9n0s2uac7+i9ZrA/SPszKD
I41G512au4VSBJknimU6ikDuzSdwaHSlY3+i+vIEpKRFwZxBEAQkqlbdrWD5+eYc
ixTPlk0m/PL2aeF/VOXh5VjT7sj4zFQ3vl0eWXYV5fJEaCRD62UDH35MeVhkhyY3
ASqmDHXwscWi5hyVIWV029kKQn2vfgtDFOMT8g7OdWoDqmwpCEEhZhpo0t0GHrhV
sy94oDGFquiRcb6Ep+HU7WnF72ePLHY9RDLrkfsgEW2JN4/uglCqPXRgL5ZHQJta
Dl8nI3EfCyM/0l0IALijGs+yUvbm3NMaNWLx95Fnhx0x1RUdpF98EwhG0PGPNRIQ
jp+P+463K3rPjkVWFnz8T32iQsiRjSyhMhrB902nO/vWSarqszeYY0fvZ6LZS4i1
Ve10qkjacs+GZXaWdeSPFQW99WVZhX65S+sxTS7ewKaSeD0itfxfKCMtExLnGmAP
5+J2L6dBudGR9Ao0GLdnSmy1WbHZgldHM9qcYSP4Q5WjQ2vwFJxM0HyJpTux4r6S
ub/cpLVrGHF33ni1oqPm45ZUmBpDhL6ymLRub7Pu3m8Q1EjQJVt4c4RkOU5fcjDi
O7zVT15xczt4GJDdH+0V3HSv6gc7skSqsX88xXNDw7VLQGkzy/j2RpR1JxpKM1EO
UWUco4uVJ65L5GhkMA66hK1VXw2saRMSuDfU7+NDxrUxe3wnlPVQbdEOdhrf0UXW
0977Zz5e5140ZiWgdZc/fyUx4Wnx16GKjDeipPU2ul+HXS2PBUJdyEyYj+FVuugA
OG+S/LeLySepwo566rTcU1wbBhxk7wGV8TaZbcIv3YmP9o0bQMvDiJ1wZi44vOy/
SG1n9KbFG86oNWq9AXhwMaT6TZ4f/5zmuk32lCMRqiZLwQXZ905ODcbaRjn226gf
wtncIU6HmpxNvnv2Ymvm/JR23fPNSQAtoBj2kJPlVAZltbNkceVHo58SEclvErSq
sOXAKbxhO2HI9+bA06yUAjCuvpHGbGCeDfFPOQrfFEJfPrZImYqYniLSywWmINXb
ISOX30XTx6uGBhZV6Ph9VG5An704Iee20HbpAK5QkcAl+kWsNoTRs6uijXyUV3ZK
BFQYq0QvxCaA076OYn5SUMxaW31q1WRhiJXA1XFecH/e8cRzg1StM5f5vme+N2Pt
wb+JDd6cDT3MvqIZiUO1fVG3w3APpFOkfesa+wL/+G7/nT7lTyWWDbPS/cTY9nsY
xOZgD20i90GIEfvEvIdeiMUosl8IvLY6BIfDRwxurMOynjfRygIuuPX2tE5LWbT3
ca9xbOD7jnRFgyCpsa0V0TGR0m4X9w1dNzVqf0rp5TrFI0mJ17BuJSMzchj7H8NY
saPJu/bAxzSvD3obxUPUQ2DJsg8CwWA9uPYNjN/oma6awm9wsR1G9BbppQGoo67L
QyY5BSqEhpfYNn7UQDTG/pomwg824ml8AsiXw1TXRJD/LNikUuDXmp4oUn524kNk
FWEX2k4s1juha3jgfkaNRIEwi4Ehjx7SssIo9v506iD+S56NPkRKN92LccJrvJj7
iQoBbjbtxXF1Ze8vByirUYDIzrLi/BUWn/bAgMtvx9/h6FB5DXtTNo/X2+RgZVTQ
TZtY86WXYvGhGFdxxywNyAie2pwLTFvVVUaYSouU9SD9YAV/UxQiKx3GBUJcpOIS
kkYd6Z3EqN29jy9FD3HzToD7MI/4RaT0QpNliAEHM0bb5oPC6MOgpc7foKL/HC4L
cfqi1IWND0emYbZ8ZchBvxT6Gz2cTWM+XPGw6lUHXJNWk2GQrwdvWIKppKiTbfjU
E3lJPijnlcaS+7SuQ7H3XICeNP/z4e+4qPdCIXwUbaY9TvaNJq0/+M70OEB24Kh6
Mj7yAel/uak2WL3WBe/lMhxRSLYLtXuXPoyBga7SoxGhipX9NY2BzHMC8xnyjq8o
x+AKIt7Hs0VCiURzMWfNSblA7h1hPmC2ev0jF+1ENttIxPgZ2SEbp5n7941GmGiB
MTfRsH8AGhCrzg+clbE3CkQ9TaW2C2y6L44nx4ZRoRqemIldz9kTIjk+FC7PKaoR
uiycZ7CQL+/pRyUbwkyPNODh+5zBzDhGsSB/x+qtcxWEzDP17Lg7bwAVKhLRnAd+
WbIgjz6PfTCFoh3HcsfDwnrxyKIKYl+9U7euJgC4HcdcCb+FOcD5dE35JvZEOeba
kfgRnQmnigvrZ/vDsrAOqH+YieQE2/L2q+XwEXkN9OUWqxyh46r/vrkeqwgJ0s7C
MyjoKw0VbufN1JG6F6gOIHGpLs5gUy/V76CHxQa5LwC4utZvNoYbiO/RN2UB0Yan
baUDzVg3+xIw+CtMknfe1DsKoUoXiB24slDI8VLOxPmJ8ujXxJdHCzniTkHkokzw
cTP1g8jSFUdtopNjKZ2k8NAp5L1jb/FsJHvBZ6kETvx9g1HPj4NmqU9jdvN86ZGV
VQeE7HqhHW1Qs2vO7dk7omJ46OhpLOgKNvoyh/MrBKtTdSOchcZzgJC/OnNu7U1p
keZXRKvvwsFvzIvZqcZ9oZ+ylb4zgsuFMoL5rLQUINNPT9Jka3SKxZ9TjjFDa81U
3CKe5Hx9UyhVV4fyr0zY2SQc6QEAXiggO/F8H99NcfO2hb97DaCiRWLAswGOyfeP
ZZ3Ht1cQJZGDoZkNUyYgc8Gfoyh08PCO07/P3nnGWWZkBrIFzdfcZFWAB1+DuRAP
bJl88nQK8Sh7D5fhWOrbYVS+5oai8WVF9pNOJXcTkmPpUcUI6hJR5siVx8GrIQcd
EW1xcnf1Slf5dUwbOMWzcMpnZqc6VJaX5maX2s6PPG9G20Z3lzrlTegPH4vJIVzl
a7ZT29fVaNgNKuc7xORKMFBXXnufX6RedLERSh5TECq7GbzpDrMB2tIz+z7Bt6jq
GulMTgzc//VrR1FTsaaZ2unArUXM5bHpckaTJcq1QA6Lowrs17WouAfL1fYqpb04
YZj5GMT/PNqBcCd8/Rr6qqBcL5xIZhA+hcIM+QEgmkmJiS7rUWQBIguXn/B0eyYA
RtAUNytd4wJJOxbOMB+T9j7VB2Odoh/J43VUQkm/rK1U1AO3KOPnlpu2lyOnh+PE
RMbeLqSP6oANceQpvs9FvpQMclY7LTedRn77d8GT9/A89y0LSWHTixDe8mL5dDu0
Y49mo26vF682hDYIAR/bT1qIfL6p2VD4mRGo/jsfEyLRsvJlp6ox91WSxVvIJ/SO
KfU03Zi+nFR3aygjykbCSNUk7WYQrcTs+vyGbn5+pZGLD+YGfGTU/EUlvUXTwB4+
Y1yh29OfPEAeym7MBvvswFx+ycNT96TsCQhbLSXU3zqUb2AnGFm3rQt7hvtpwY+b
CaU/+YTW/WtBFfkHHgF425REA/qRufSN8JePxIe2QZzQPeG+L7ja+4YXzlEcWvrA
X5/mKZcoJ0IlXwAn2gJtP38/+tmxzWgjTQqqNs/qks8Wg6Mo1SbOG8vduKK++kee
5J1VoxI69rgj16yEpY/nA6f3CqpdMoppaQOasynDuPAyqYrtpgKJM4wcfx3jO+50
lrYqshbghI4/bnwPsNMx6mmTk5jho0KWw6ukhhldwmvtXzbYtiRFsKAeDuFypnVE
8Ij0iH9fX6I0SqSixGJtoulpZxkLcbzYkNmeymURotCL9DuxK4Xlvvta9S/lDfLF
ElRJCN0jGK1NvQZoJ8uOo7FsRwo1JEL0B7lHNDU2ZEp61Bnf3r0Ga85rv2B8geOd
qnmmZWRpmb+sXbMNNs7sp3nCpqbMD8+0BDLPtB5TbCmYP7dAj0UEIk76CDP3kEIT
3VFDMcpB2ByUpV/hgZFSC7qXp6Hg764pX+hMh0CeIa5op1XgLoEhodgRKuNl1LvV
mcM5EvE7dCEQPfVde7A5u9z3s80xbVAW+MhtGsgqo3DqxBmad8gzta8+1qwi6Y/o
uGd59prh63OEg7kdSLyDPWcnc7eirKAxmms97q2bkgHsW79E5HhNwErkMpwDrDeU
W87ADzgT6UVv66x7+oWkCSmUo7KK8fUzKWqGvOMzrSUca3ajgt/0IpGW3nwHDuZO
NPesqtbhhbcdXC3zlCZ0iJYXkAXdwF/MOmMX43UhvLsCmX9e9u314OerETS2jCIW
xsEc6OCOZGG0xYx+zakPVA4ETnEVMARAqj4ri4kC3nK3NIVZs1EQHA0qbjxgF+ri
xNlDx6iiUES3uEtWYDlTsuwXBEdyCH3zdULszl09hPXIy0RkZT1rnKENPlhXDI+K
gEeJBw4ty6XfcBMoS+dfXt5ybHfkQl8lz5qh/FuiP79405LNJJnn2diU+O4Osdig
zPb/RWPPKHZe+6B5ASw5GB9/zJFt6nyNzWBPCyCUNq05zz0wfOn/ytSw/RYcGzyM
uWCwWPRgM/3+5S2IHUKwhhqk2q6bDhFVwEJFRsg/GgOkpv+YByspACixoTX0Xr1i
jQOXH2A77gbGuo54Yy1/LPjL8ryoR3liHNeXcexcG+Num1N9FHEwb0AQss2BuHvU
Q0/FYKoW5hpTDJEDqHVpeLdm3LiQPqZ6bWuGWXpYmXPLjD1AUoWrTZotFYAvAOJF
YuO74gVNObpMi9UCKjYPOYUAIQsqsogaQJNP7vGbrLwDXsudwm7ld0V1C8lTrFW9
h3Ot5KfIi/vjZ2EB7D4SkD/WPgUamywy7T49jII9RC4JZz+UKI+7ofGwnSvDCCcZ
x7qQYGz3ZSDBnV20gXMMm4CLp4sqebdzIObn6broBY9eE3eUF+GndOAqKccgGehL
D1tdvrDVSX8DCha/I+/m0Pc2EovoMnzqihTlfgjODlf/sB/RpG1+GaI6lfr88Vu9
glM9cOYP5CMUhrPjOvJKAPV8ezP6juGCubK1nbV0t9A3jVtJo0jRRgdzbKVgNe/P
mhSeeCwMMDKn/cGApy/MSRexHVXZiR+lM1P/Qgj+bIqRkVNViKumlA4s21YWWouS
u8fhgjSKO69zmRgFAuJcohBtO8nYX2MB2F3NSVe6GUdatzsfFnpu3SuZ3KMRwvxf
tPpyTQs3ElQZDYWzQSnJ5ma2cNcGgwvE+Vxnq7MTcBCT1x4M99U41TyKtu9e2HgD
plDfxKZ+G6hKsS59WnXQJjfHxx1BC7HSYPpUHFqizKf8926kE3YcTVOwjg0IswJ5
dBENOd68ENUFCgkz6hb4Qph56wf3fg04D1YxZ2H+SeOltA0MVcPfOcgaoUycttLz
XUDK6hSO15naQO8O0x+Fc4EcSWEJFNAZc0WDCIhrdBQWVorNjUSHQg028H0Q04S7
JtTPtwLubPQVITbQ1coAxDukhpNGhgvFNn+RuAeaC3AoLMXcVb5yHqNpfmye0nAk
xnr1khMsvsezFzISCf2fB7ud2F528SPL7MgD9K8CS70gOrBVmY+mRSRRR4gNdsfx
yj1cMtD/jWt9gJ1I2/2f5SVWZ2IdFZJEmbv2473neUlusR98xTvlh96bGev9f8mL
uXEnPmycUciP4+u4v3FwGGqWhVLDK5cV8bR5IlipfQU+4fY0+mY8aATR750mJ0XY
CFGUAFyUvktJRtL8hGtqD6YBPsWG1kO+xa68t7PFdTZJfqDdRSrkOe9oQgTbq7iM
llGFdkjqvdOlXaGWAweDxXLaztSyi+lzHrDFlq/AYJXZiaCRuVC3tt5iskDDtmsM
IJkiYONOUSmrSl0m6+0Opf1JquAmnHRzaDUK1MfbUxuBVS9/b1iVrRZKkp4NSZhb
7BlwxYaqO42GAC8IaC9w72VmLJBdXCvueVpqzlEg6c5tO5d0b6GZ4bkGO0AitM49
kgLTEF0XxeiTQxDWD3Wma8ebTQrPKfpH1nt+KAH/hs7Ofy72Q/Kw8UBoBmX6wIOe
DKfHOgViPEdqQ0AFdV0QzET+lqjwnccKhxv7keF3LVTUOmgv2Af/hXBxk9714VoA
bNRa8t4NSR+8f2D7pXNoiF9nmQQxMxfUpuXzTTmub1BYd7Sse+/7mRKbqe5R9qis
eFXaDfcgmNxTP9SIiPGf4NUrZ1T2BZpNHkkDwLmoRl2R/HRjY0bLjQsF6t3E3T2D
B8qtPQrbdLhTBrmWxBuuEqii3BhEDJyC5hyZ2TPRNRDkILRWT6Fl5eOchUwn0FJC
5fD+k3CO52ta+3YvoS5BZ1UcE1oc4enaw5zDsSmryeAeq7QYexOzbLlXOyJFPBA8
De2d6W26kCHI5uSbO8uaZxtpoLEa954Gs9Z2pC0qMDtA5J+1sfTQYaPpgnSQYVID
n3BNH38GACFIFHGY00/MF7YcC+Kjj4nJmNkRUcsYw9rYe/Jga62/sxCASN4eyl2j
qUKvexD+/MCTTSUhNvRxjC+zdsxOYMtrFCXKQt653Aix5nfKGNbllQu+/97zKRoW
Ntw9+BxF+LvRqmuIRtskrMgV5mayzbFx2qmroDCJsof+FnHTSLamlGd2H6HIV1qr
cZ7yl/rX0lALvD1k8yhQK2nbhC6A/nwe8qpAVxH81cJ6UHe8PgpSMY9+ECZnNTLe
ALptDYNX04XJ/eazgQ28Ou7R4Kk3ZTuKGA5l/JApanZ91VIAToxYuhyWH+zwq5UH
4SmUxE+VDeCW0zaeGjCD7yslqOehskIkwVla3zOJoqAx4uAweFXVuFuN2BEEIIFe
FCXVQ0rHcrJR8eQouKC5DMlbTs08NdLD0eTKoS8EXl6SEcSEyAR/hkzVfmsZFHJf
ULlZSN06atYmomaKJ1reH+Z7yNgPJhayizzo7v/o13fTT3BryatZtvUe0QhMJsyX
Q3nl/g19vWZDV71roYlKfPIF/6EXIVpnaqDKXDrmb27+zsoZgsdkrq52btJ2/HRw
jRIVpfyM2DbAoYt8ZGFWHV61VXxVI8VHoGihzElqkWrBc6fa67ndZP7Kz19UZ2Tk
cMWsEUHQ30tigfcYJ/72fa7rZoubFOevMZ7RjbdVA8HvQdbBW7uZJ0IDknMDysTV
lGgUCa/OdGmeS3MTYKYV0Ky62bSyLgSAKQTAWnYGCaKcJtypZMJz6e1/WOcqiiKC
9Nl2zYS3LBSjf+vjvN1/rF45tILuykJURyGTNnfhbHwSwzYt0qTu6Nq7JotsaW0U
ThouFJeYoo0ZKxF72xhF2JojebM8/yUm05V8kdBsaeE/aDgO5AyKY2zmRfN4hrpN
jxGO+1he5SwlZHuMsW5bzaTFA16ShqIvdbss+3eu2qI4rBSfMXD1NBhQFErmaDCz
hb9e5dEKkPJgnLmBWYLQwaGvFamkZiuuXfBZ4O0zn7YlMap6i7+05hH2mBUe88tU
emR/I69SuijKLIDYKhxEb1r5bSl+JhLLCtJFH1AfbvRqVrjSqrf5XHcvTUObb1kQ
lJ+hiQeIfK2l/MKAR32nkSz4GIlb3WVFsc76vNCLHZJ/juxXruAt8Isvn0bD86jg
b2UN6SQDop6EioiotoOXbXYw4amrdg3WDiuDKB6MGUcV8MATnjY+KlNehpM1oiyN
O/5lso/+BzwdHiUi5irXbv62AT/CU/XcAMDk80rsRmaHJaPgFneIeSC8S1BTzwNJ
KzJUG75TPpr4Er/XbJX94Rc4m40nAzc+D9YFNHzHOfgwDoyIE6vxFOKLlYtLu0Y5
EC/hMhxlM8rLBnwwyo9zWNP0Jpbh34YRC2e+qGTB9fAzgHcdNv4cyrqvnHGGdjkL
PSvZCU0fNzWhIhHYCk7fXmYZ6xOlrlNTIClvQvEAMiC2zKmAr0XmzZMJB4TFfWZl
7x4Got9bZ7mSFA+Lvo+5bluxY7D7Ct3WwHfslNnp7s+f0Nz0qWLOJqrRCZIYWtlA
AGp+7/ZIPRcqVQESIzam+kpZUKqS+rijp6/8FwKqmAavuaze6bOQ/oa2gNPt8vC6
DdMfAx5OZdPyR1dYXPyUzPDTHw6UMiSDEMySlQpbA3BqaEFOFvw6Mf0pL2exHlmY
G8ON4AyKuBITg0hw+eCiklGoHDz7/y6xMFqj9kbRAzIjfMcqJpHvNnVJowuMWxwE
AGUYwz0L+KoVNWwlyP/Wg5GiNQCcOU5ggFcvICYRN6LUzKDeIGnIQ8wR3nwRT9mT
j3WiR9V0kvjl+q3rS/0H8hCYnRvLuQSn0rBE2YlgoHNO9UX7xkoLvBUdnrcQB2Ct
UIlcpFcb3ti8zyxrNZkqunQf7agxul0gzKA/wLeuGQ9jpo0UXFtCXFFwArXSkpJa
GNAopmSloiACTWtlTMFmfDWpJ8LPTvIt+M40PkF93JxBQtju5Sseb/AodlSUxAgc
bOy9UHM2Cp/DW6iAtQV1SHT7cnFChGTz1MxMAGY4zJNyNzpJgz4nWREhEHo9LNCO
BFTfNxY8cwYfDPH4Er7rsp17gFKnqcZjgdB7JlExGGFe0gLKHdi/OhmuAD4kqQY6
87oRlZUxXiRqSFsPgghQvKEGal3QJWQ2o2eOEDRN9Qi5U+Ir7e8dn7ZmAP4nSrQB
mcI0QUNzFZoxbKgzE+s/4bx1pJ86g2UekYUOsi6CjBXqGp6+cWrnGaPztb4FfG+0
CGnASMceSV4KBYgmWk7qV6qh8T7Fz4jspMcTipZUocpnncj+6vH97+8N+V0Eke+5
4E45YBa0A4Ro77fJUWQXjl5L/7FXw+4OdAbwyci82zoB8v+a3G3UzNpHqaEaw0vE
Bq+n0nolPyOW0VKkVHVkVq1wStxSPnlkowBAdkP6oynA+asGnvfU+Kxo9m65zrlS
CPB4ARsSg3H09/RO6s+jz0LkEd0xTRzCUBqcOcSmcUA//ivD/yw9wDPaTYqjAmM7
HdCjxh3vual5b8B6eOK5n0EpyoY2Hne4VLHHgun1sJp6W2c3e5lPm50TqVXVMMHc
+ZXOFS7TpBPiLMaNCYnY7RQO7dHPamvkNNr0CobwUBtcMpODK0tshHBJPDW8ei4v
pRETSixj/YEnexqlQgO+clVMjDsD1jtB8T5c+9cEMQvHwU0GP0ZiJiY16atjX60+
nifIf0NxYVufXvxlN/V2uoOFffyGErylmCfypOyDj9ku9cAODGekcCGRy9+QJ58N
BWbQm2Ha8weOoF/0+dFyigRvAvG5nOK7n27i7ven7NFL4x9/FA9ygf4IrwRkyaHQ
AMmmMhW8QOe5fXs5c+XBmYavs33Qhk+WZIJEMBRjV4J8Xo3MRWV53bu456TavGfp
AANoKykkrY15tQ9E17Lu3gLpxmNL/Zra2bNQLEkpL9MFintcgVJwYUbzQh+M2YeN
0X1AgXAQDJfMoWUiISJ2YhBEEd7bnimtQEzERWfuhomO5c7aAT4mkm12yFJQjOnd
bZLaroL93HKakevGC1Z9dm0NngMPgjjB2NA8bK8AD8qwalbFIj0a4iShoOxyAzmT
zhtieSQHqz0sbpwHdoO4Y55eFx0su1vI7apzagGSgn0fhJL97aw6B4vdaUhaUKG6
gEnymZmFO1SEiwwIUO8eoswcL10PtnnpPPbZ+BcdolVks+uS5lRBO0EQKkyUJc/S
lMdvuPA+5fb156HmsQEcxCxmMnSOtFcNQPONKlYB6kxHkH02HjHiKSBT440okkmB
5i35EA64lNkWdvDVUjmpmaDhN2p/RFv7uVp4Jj+rp8NcKUPXEtLrTIF7uz0n8g69
F6swoiP3fabeeoG06kDYfeNeYuQy6ry5DKm6FzURx0aHrLjmGPR+m6rvP7j6i1bC
C99ihp8LdzkXOVB5ZsgRfHElcCMS7l+d56SSy/oIMSk0EUAnHAJYYlxXbvkwun1B
3O39OXNry43xlwAtog9jga5LLoNzP7mz0le2MSOxID8hypTE17MJQWVj7f/OyLwu
EckOsuZCl0xk5XTQOLUPxM3OMQgoDcKThmjo4kmSNsf0ldYGU01GKzQPDAGFyZCL
je/J8nzntA0opYjTJQOl+PWcDch2LvzjPoK9r3nzHuPaWUcNjrifhVsOlhigWeOh
50JG3aahZA+geEtjVeIlc6NjYTW2e6/kQwD0tAQIhOHj6Oda/JVh0Lwihd6OYkj+
iRh2JTe5SFSnb8ipsH2g4ykEKZhAAkog3PvECbFjpXe9ZExUkmL6RQuTNGAugXn8
HzklIOXyGBoA3eXJ29oW0+CLWSbOQZr8hPs2OZb8KIkNYAKj7k39SSkQDIynv+NA
BR8EEArtstjajbW0VJTDM3nqQfq/bFamZc+9ojSSukefygaJHVe6qQiMGbC1U1MX
sNEEDeMJlnOzUy4swgtRaHy6BnCbytCSp9T5zw5/Z+2/PZ0fZA7B9FbwfEqBReY6
LZx4l75pFcc94M01ozjLTZXTf2hqW1AuoKquuQORss+stWyeqZ9weCSCqtGKJli5
9inB6Q0rZV4Z705ybdoUa4uwRD5XwA73EONOd7iAf5kuTZZGeULKIcxZeEdVbAPh
Ii8SCtm+aXaTOlDT8eIKxtFD5NdTMwAa101+RPqOalikKTVJX0Cv7P6mus35e0Dd
Me9ak+o5B91q+J84B2e6FK9pWesArzKGboQ2y2dVt+PsDIhGL9d4U/kjvYntM+AM
/SmQVnsnNYtP3mOwY+jIjCAtoVM4ZWmKZI0JqLQadBl5O8X82Mpm0t+iOL3EsY/2
BYIs2F7KB1AQG1L+hAAQKGlJEFRq8VoQ1RG80PyrY/a1FGQEtYHIcsg5BBIAaBFC
iH6dksOU25pyHStIbKGHCgJBFc4DDQYgbqXsPYhIPxRmKFKWmzuDc+Ubvdg9OA+7
Qo9tv4GJuuKjj0akeQARf2ygVqjl8TxvZhILDBeASaY8io35wfVdhdWGXft+xXOd
fmDNUL73Aqtl3XfTSavM4BJKLKEqdjnne7+8Aqxuz8vm3rcwsaqquY9NiiSUCDt3
ZsKL2In5mcOL2qiGR1Y/CRS005C2zxTBugIWyXTbAXqVJk8gnUcJJIfHAgUEolhj
AwqbxeGfSCygqqJ9n9WPtIC2AK/D25XtGnWrSNB0v5makMmm3xajgy3kgA9M08Z8
w93rZxqfn06YvHI8tDQN36NWAc8hOlW2jtR3tuarr95jUoWkr3b6YCXWDV1ls9VH
YD23TyZnb6pw9AkG8oAv+193Th468GINOG1CryQ0mzWyLTf9aNq33p+q0slSQQ1T
6De2RGair0GtJavNxluhU3zgC7RN8a3KBWKsbvcG13lgq2tJdo4Zo6bqkEKGJ8XA
DWYLy0usAmNC8SQBmQsb5mP55cSZkQRzLYdtzjCtFkw38GnhpNIuljZO70F3KcBq
5iLOGFuaKXQm36FWxl7uuDG2TYAkASaYoltA17n7ALK4KDmui5zwiWcoOuEWOrTf
lzVm7AtKuTP80EH4mVrneolH4LzwndwotOUqJq3ZFLeSSNlY5NYs3xKMkBocSKhY
rUACUw2jgoSfcMLFdEaOvD/EGLF88U27IW7Iq06MhREGqcUTtputQpvVujoFS9pI
wBXpq+At0bxqVpi83gCep5YHEpbQnTK9ueGUclp4VA9QpivXB1IYpHYeKOQ4Mrcv
fzh5G15XJ792FdpurKVdRb/rjxUM1qFLLrSfQ8ZI7xDvpxoHJGAlTB8KgAesf4eM
d3vtN7thHfFtfjSC0fvfs+w3TAAMo4dPkKWQoEe0E4WI06/Z8J1s1VcGZ2orindu
333+bhnFH7BcTN0XLrVQZvOUYdY6IFf97FKe4DyQg0hXbTP0oZlYukGXqwH+v6jH
oiad1R3Rh/4B84gBAsyaZ0iCngNmTcEaHXLdE6ux0ZpFqnyPs+CAyI4SPh7xYQJt
hlOeLzfXAhmzeURcpSwqEKqaPw9A6fN4adezeydqVOjOLLTa5PIKTO3TyganSMt8
s/vPg17hnY7LLa+aNNGAxQtzQ00FyRUfA4Bwy4H7mDzX71hKttEnNStiAY1Pd35X
zZfRttmm4/D9kKvkpo2elTKco1JuVPkfObwSLfx4DNqnNgBNmQuvIl2WhnPWAnur
uGYmA9g2KTIfpqCoctQPFp7WF0g9UT2xfZS2n09dqcUtUAzDaN7xHGaUTE7IIRbs
a5ztor/sq0SZQYdNt7LHiO1MpUGITpHeNOgb5Po9IrS1Pd/Z4xaqwgHtb2vwvQVv
xXnYg6fpsAKFiviUboWarnbX/WeEoMdzEyMKB9iESgG0k3+LoQuVDjazOejVItzo
Z/n/erTXIB2Avry28rEV1F2aRDq8lvJJ083oXE6ANlY9KnvOLLfxmxAD0xq9WuLO
AKXaO7qNSncjYLyYIs3Ce9IRUEuUdmYkd1Q8j0vYgmMVjP0zAiLP3e9ipyC5RfdH
dXDXSH8BxpNB/sk+N9Tv41II//rvFC15stuebrlq3+Dkp+1G3UQ4tY6nwn4WlzYk
t5G2O3wWfTY4cWwyYCLYztmWm4RVdQO5o9Q6IXp5h3AujS/CVFsfZco9O+gTSFwb
7tUJfgF9xYscXBnEbghDyvC1xX5M1NdN+FstCN3+QpJgufYkAEdxKgwDch2oyOIa
28Mnlg/ZyafiaIxNgV0vcf43C1O4HERuZXuuFksTVeUX9Gv/IG5cA066LQz/kI0V
cr4hRmXHAOiHxlzfvNCVV/G8MYa5Pxf1pWJLyJQhWtcyraEio/zQ9VLvV4B1IrOs
S6EN6S5zWrOABpiFDf8fM0Xcp1lPduDg+FlmCSvZnts9aE43Egme1HhCfJoMM5Io
uKorWICSyUnxv1cLNzo+jVXe5ZBFsPT5D/oaSS390NHycdHzAXcMdmHuRj8wkQZ8
NXNSQlAS5mRhNF64212geFm1X2XMhWIe290/I5ORA/kT5PXaqTE0+AL8uZ9LYl12
mYFL6AKawaPGo2v3PR7d0U1QqprSYHqGZdD74XmqlBtxKHDfasmjy+oYtjD1ubGT
bndtlBF3lMbJvsSKgwRrWwcc/P0B0Al3wtHe76mey83PY8arWC5yRBbLeFCyjt12
/uLWQDKLhGm+9Y9Ki1Zq4J5+eoCn5bY4x2dI2CtkeAtMpmsW9VTWyXalHyfcTpby
if3NK5y0Upjkuz+w2P9OG1hGlBfrEM0jd/PW+Coln/GI/pgDER9eY9dA6iZzeWn1
naiaZZbhecTq3LOaLcibV6jMddJmlLFbpcv+dgLJrZKEp50JVZZuPpdaOmj5jN3q
NO2061AqQ0I5l4PgIHGUj7qAjSEFEA5WZXhbLLO63H05gs/sEaQTkopzd07oDDaj
Gwox4Dc5SxkV+Eo5woTQTuRXB8wiQMrZPOlJXneBsFkrQyCPpH2IbnTWrBWrP6oK
X1YFLWgjTU9WQn8zTSJ11ES6TB1KLxEdnWi2WGay/P3VhQp7zaAbPj6VH/dxUxwA
N66uxZ1tSbXt314IjjmNkNbMVllWgwkipc3eMyRmY3BH3oOZLeVi/Nt+THYpyREN
MEy+t2BgNR3uRe22s7nw6FHxVCDOirGLxwT+FtwnGVIcCC9B3CeEtECiJftkAjlm
2GAw1GXxdQKoXJADyYITWmHJiEBqV60cAkWQ2YR28xBYycrEsGfLEssqe5frFBDA
9vJKbye9WBvEiD/9Hjg0wn6inMxsSwRzUWupfm5nt6coDPTSrGaKuIhYoS5G04Lp
9+8W9sqOFfTmmKhpKXlo5a+yKyLFqhQfm+YRgjRJbUycu+t9BKwtKJQVnM5RqQ7X
L+H5FoLJAnSW1UdfoW6RnKG8okQ6ZaSs//CdPocwr43uiQDtRdftddgyFT4KuHlX
xlWhOrH1abTXzwTmF7b6stRNHB/5yha4+B/xrXGL4gp4vLv50LWEO6aH+cT0Asqp
8Wur9TYmJtd6vtD4PLyUAQzSaQo2jJecQcbQ4DnbSzQw+oyLIj4u4DzVNF2wbIoj
NhovLKH0nCbtvICe3A324Xgikv/eQtoAnub3zwxa5XHh696cNRYTLFicVCkr42a9
N66qIZB7bVYaB/1IjoQn2mr9GbPjgWET5P6DE8vwL9TAuV+zV9SyEFIq6Upcb1VV
kYYy5/YYD9PT1tlGgh6iM2z1gyqZ39umjM8rwhtuaDXlsMObdrGZVk+ABtaZagKf
S095MxEqt5SEbO9qWZ/2Pf/OBR/0eSXQKrHbySOrn6IBkhcViyQ/J8bumHy4EwpG
mVb4b0ovkeEia0BMHot6h6FhgG6zoDz4SU/t4nVhh3IPia/wPmgNbTZm63ZOq89d
v7ypBtDwdTIefED++olctBfInCioNDn88Q4VhBpmW+MwiV+U7sJVxJ7Qg3uIq/Og
czXc3tLdbNirfnbMgyBgymCHLpVSj6XlJzAVxeAIpqhZoTbxT400m4E7hZ8mtQVF
C8PM3n23xXoB5C+3uBzkuYbM7h/ppCQXvkVZEJzth+2NRdokKJYO8/zkulUyaRdh
hQ3RnUdqBD0WJg1HxUGcmFxd4u1j19UkINZGLRcGf8KtfuiFA2vkQX/EtUSvUUCu
hx7nFXvv2bLWwtmgCGLcc8DACFKqEnDABYzloGskPybgwDX8YUrw8+WJ1N+wZ3S9
R/4USqw9HN3usOoLPuu5YTrQhOdHrI7AnCY6GDrGlf7I1rkW6ebMfjTRvMU8Vbs6
R+D/CtipCtuFyqaa/VwTDBs1dnOkOw94CyRggscR7smBu3PAsLLBcZx3P6zWelt0
o+8zNf4nZ/aHbkonWcGVUnZzP83ylOasOHzEvrgZorKlWwe3JllLasehmS/UHUIJ
w2xUGWK7hpZ2lhU8K61KjDUmktZ5/4LSs+VSpiIhdwfxAf8wzjJuXSKwYuuQeWvH
44IQlsYoj20Dr/qvt3oJDbFfUXu/em8n1k3WfSI+HBI81fySWwCv17PbypnOu5sx
fjPS/+EEjdog/w9iOTXztiaOgeKzi6omkx5tYwrGK9hLyWXR0kHbqDZoMOJfc0G0
UEdSsxe1ni8KQnBiXieAqGY47N9Nf8oRUnKUImM5svKXi7dcMi+8KtkTKRwzf+Ki
TjUzyW1K562ci8Hf88Gu3VMBnblFRUN6ljy5HqIfjZMH7QOO3b3OG8G6S/FxGn4c
LObd3ySFgApEQnZ+94KFp8xZIWcmA2aP8Pn+2ZhnFb/3kHO/KwQ2XF6/NGQcx0NN
rSS92jpq7g4DpLdrNw846aBqElK3pPvcFjFuitu5ysF5lCxWZFQjC6g1Xy66JVIc
TsettDD3BOBJBTddd+xhQPUo9LE2s+EiowCvowymdEJDiDKOBgTTNf8j4eSgfAeb
POk0vMBHooUdlnbKWZQgYOJMfaXDvFxbzmGHKeVelsOfPHQYdskNQYDPwYoq6Vmj
BW18tN7IqZepBIGU1nDZjeTivZF3+t4r5ca9QxLRaFm2l1xYBXGwZIG1zu1Dz+Cc
SzgshjNVLPdioAxXUXpV22U1ChveWgBt0esQNiO14sDjk7DV/qKPFyml1JgQ0n2u
gj/mvE71eRZHSJd3IeEVzsAX4cNcr+i/SgAWuZKXI3IwePpatYMqrMgjhJ8DIOV4
hkK8zkuQx/0OO1V3kxBeXfvPnuIzDR0WdBPFlBHgGmKObqZY/82Uf51RrC91Dpuz
DZkAooAA2VFlI8ZkaDf9sPcLPAmoTU4b9rKlNusIkilj0DyW4aG1wrjnQ9v1sUIz
Nkf+P4MkcNaJ90QJSvejiQeu/skhGefzb1XJ3pjDMwdJlBP1ba6vWJf+vioozJJO
L0ccBf0E3iHVI82Jl59yA7E4hjutzdmrUNWTmwAP18qunpsnmCE1fMPPGHYufEga
GCPukbSC7VL7vAMx+Er/lrOkdn0jUeTDI+BdtGEQZ9ecv4RSJ095nvSmje1976+c
vKBTInITrQv8cHQi2sHkt9YN+jdc2v+l+1r02gn/HOxJ5fx2vW+c2+mue4EI2B+h
WUvtkvmmeNjEDJEVDArxK/5pRAynbKIGqskq79t1gVqiYTdq0HaWlz7lUDWZpZt4
7YbZ94+by/Xus3umNFhbnMDrFZO1H6MCqcpb37qo5XfMgLj0utLiB5rY1ncmayDM
Sx4HcGn9RkGabXLdnqnFFljXGwWtWvi9s10oSY8v0SChKG9m+OuP+l8/EzaK51CJ
wHs/G3RT1UYXBQi24AHRcy8y2jydzfhbOcmqyL8YSXF3Y6zFEcIkv+l4fGOVWUYR
MOG6rTIF0YtPWpG0PVLbiaBCIxGB8fBZzlp45/hJcYRyKnCM49WwLJYmWWTy5DrG
QTHn6rHGQ/deD4mit506EZ6dXrB0T7rK7BqxuSFuB7uxN/9LmrPRCQW9AggUSJWX
sfGc7IYBxLNi05xrhXXWASYnB2OsjGpSun1rnJUVPvcJEwJhM4RK9wXEM1Rn5fvw
MQs2PkA6RFSM6DTUiJIklttk0I8sA3sGkUg2opN58JhtnrFQJmzkXNkGL78/68/t
rV1zWDwRtng7AmwRnXLD+yfh86Rh7zekxunehMRJ/eVAXC+uDn9d3v5uGKcoYMx0
gg6+Bj8XHRa/Prjg03rvGhVHhoij6UqEArI2IaKPxKsyu/1us/uD3xBk8cIFq1nY
YbHp815UfIvebZ87bymq46vayfgwzmsc8tDV0shamCJwRaxP9lQyk2JdHZ0pPztL
0YSlJqEcYGYOK+whmZOHa26KKERJvzelEE6Rw8JtPGAQcYGRLN56P+AMGYHOlgHu
T/kmdHtAFku2d/dB2B0xmBmr73n7Oeml7MK8Ef0uR572eDtrWdJqNoLDHsVmlaUg
U5LwM0iJUme6vrO3di+ZiOR6jVN3hWqLoQQrR0WWEAq1a8xRAtHX/M/xK6Qjvrt9
cAFp2vi6T2xYRo7HDUDbqQPjkwipyNyoz2ESRX04zt2QNOOPCrveAdFLr9QRtyY2
7UaXM49GqVBkH/VGCeOHfslCC8fgXXN3+Pj+u3Px7i0SIRSjJPnGewQpMz1NO4hO
sIYGZjSb9BC8kpECA1uMLL52fYNKKRMX1R+lGnhDzszKyjGO2Vhc7ZcxuMCWxNhp
xN2AbZqGHrtlU9fSA+m53rvypdA/YJQqZ6eENKPvYjMjIAkB7XgOl+sCMUVzxs3f
Vk1sS3R9RTx9e6FC4TYRY/4cD6sOJULK/p994eoIffffuu9i/zAqNnfHKAKyNPtL
QhyMDnRT+OanhcWNdiZ17DQlYsfYgtPC5oNMQxV8amFxRZZJPZYL6HYAoHxw+r9V
dLbYIHuMqt33XEdjBodARa+wU3c6trNo7tWgT952eCO5efq1zk21cFIjTXIWvdUF
8c3K7Ot4aZTVnjOOOplicVbdRmqxOnpnzQOFCxFaaloLc9zyiSHXZgknWmTorJdA
UvpFLelM+IW/587REmGUE9H83kzGTeUqwCQpCu99wsNwgkwGIY7krC1aaiyVeNdh
V+jsghXpC2y+ZJeZFF/j5jkyMKVG616LbF0d+bV4wOngMeltk7orykFOp/ZTFQ7d
iyzPrWnx7QVSRm/sHd7GJ27px6BZRVmpXbkiV+fzLurlRk5TJIQUS/XUqzJiMsc0
j1YgUrWW2z2VwSjpYR2mMZZlLUDC2CEz/XNuo9CYmjvYcYQjh4soe0n8zKcG5aLH
sl4IwJRwl+jrQE/FN1VAqsvBWcW6EMldxdOPNAtZvKcvh98LbCKal6c2TkJ/7VdY
kwrosXEcBVyFIZ2jQ8IHCVBrw5pVwrBrCDnTvI2SLHKMt9ePxZE4UUa5viIyVsmB
BISpL6zAWvo+52lL46PGrk3a70YBnWNGGaVT8y+jgTnw2+78XWpcqsqKtIL9RLXd
o3agOf7f/ZOT0qc2o2JE0JhxKyF2T8CMby/HfvqrErri6MK1wp5iEsVuAVccy/si
JjEq66Td0dv9FnSM7YRj7TYq1c5dtD0xJCXqPE0rMKK3EmbMuQlf9siwrqdpuUms
rKkgu4A27bP4nUVguS4SORTfv87UrlGgM6qgIZ3jns2g1PBZC3eVxjxvvAOcT17X
3+YWUPWKjm5ox+DGWhvvG9ZdFWPnDo94lH2n4catxmd4BpkGM7S2Jo/hSx9QmkwU
+ljyh2v+IE5Et19BM7DnXJvIcQkWM1BIvqtEJOwcDoF+5Vvk1ErOncFFXk3m/12Y
JEzfaZyhiPu6ZkVIx5lt6DIEK2b6L3HoB4b9hi0WXLUNfVc1ivz+J+rNFVIeLtoy
gku6wzKn8SN6j0uVtp3zkOl8lOzXOPsmev/003xi9jvLU/7EgTahonPM2vETAR+J
J1bxSp7cINtuA2m0TsLQoD5z6KATlEnherrSTtzmlzg8sDCgn3860W3XGmCt1wwi
oiPlwv9J8DBLclYVfKZ71qi7M7sHsVeSSzFqzefCpds/tyUsreHphZJxx5neiRIr
nO9BrqlJp/QZT/ClwJA1CZzTeSVdiZhwL0TeeDbbjnZDQG4y9GMi2nJsdEKKmRrf
w7Grxf5dljdHNCv1/vyvkLgy47nZiqXkCK8ga75sBYDPmyCSaphYrzpkCnd5JJOt
loZh65rEq1fLVriLq/Ik5BbNXXJz9XiLbiPQaAREVLc6ngXRmBzDD4Eo4aEiHjmt
aiiM0Hsnx24Czo3bnbgqmH7zenKbMjDa92fOiNaEhgf+J7qSH53GmPSsDrIjyKvA
rmPfKSaKbyaKHrF5K1p7Wryz+KAK7Xl0V44i5UnL7+wPUXTP9ysqunILeTr5aSa/
R6ZO1gicjb1mADieefu4jPR9JAYsUx0YvYng8R9Jn9bhvEjJjCeU40rueDXJYmaQ
+EHnSUSwjOHI080RnfSFwluD1xhO2yCHiQ8MCgc0H3k5d+y8Xcs6QUploOmUsOFF
ZdY9Mr/2D4ID734P+sQf1AqKyMvQrwlfHnGvMzcQr8apPBJJ2MP2NgOCDMCicnYk
pz7IjleSHXPUs1VZpjMMIjPuvxXcBTtqRJRNrlK6UC6px/RGySTir5MsVqcbS9Dw
5J+2qa8zYH3uYMkwohstTZ91srmQP4kyd8Lw6jdAFu21A93ZwXAD1Qe0y3uNVSdW
yXTebMuJ1bh1OAqU8eInfQak+HcMnkBfAuasDE2wec6+whX1OPZv+IMnibJOXU83
v8etCeExnIbfJ4Kw+DJr5/sfGilHI68VMeyxnfJhN0JNpg+s24ngR8sgE5ePk4D/
/G29jNkirRT4BKNrazmfSOEIU97LI7hdEK/EAT4sxXTMLq+rYYvSzKOHdgP/ygOA
BTPwDB08YV4OQ9BzUpJb4IB32FjY6t8GdMfqFx4A2eqCaJ5G+O7u8X/5FNxF5H2T
vRMHQkpdzqzJ7HPQHx7MBUYTuBkMigqFA10mFZe1WdFvxkwMIGlfXFzFGlZI3w6x
k554EEibqsN5WWfhWvn1aXUoD4fRqNfFgNtOFpVHAtHRqctJEt2ADT7HPoEJ8rP1
7uBkTxivG2t9Ox4gUntgbxiPg7upP96tLHV7NgrKG/QLKP6qhzMBfSEsNoXRe7sL
gHZhxBREMYIFso+Sk9qXZrHjk866ZHt8ZgP8KoVvNJvXB3aaLX4EPsDhqp/Hhb/3
VgvnWlYBwJkz2YxFT3ggfUtFcYx061TMdUsil2f6coiFZxVwWWpOwSXpgeAB6A2z
zsjISGxOjCme8I5F9G3qO9JTkDZFh3KNvNIruDou2ojDVw+RPJNvUhjLlzYH1Zsx
uYNw7Lcbq2fM1JGKcJ4rY3eJis9tihDyW7xlK7NOZRdXfP+h03epzOb+EUQ20wPD
yFiYyEEBvPNyYMfiETQGG6F3LRoA0I1Sq/53IJmOhDSQZgA3WGgEzr94U+Wo/pv7
0F4zToXvpL1/T5fe17ZHCKPp3bT9i/AKmiaOe5v7W0bnbJysOMFaCm/NOFu2t9Sp
PEfq+3Us/3NWcT5k0dJwJSk8kyNe2Glj4oXybGd3kJY5XRLSaN7OsoHb7veliTpa
yFKo2//R6AaG1bxOyL5hcf2h8A1XhHZtE3Ko7nkTg+UHZYkUpZIWwEkUJuOm6qEa

//pragma protect end_data_block
//pragma protect digest_block
77/VBKBz6BIDLuJntxZBUS8vQzk=
//pragma protect end_digest_block
//pragma protect end_protected

`endif // GUARD_SVT_AHB_MASTER_UVM_SV





